BZh91AY&SYkEJ��>_�`q����� ����bG��     >��V�
"�YV�j�5I(��SZ�Hن�
U+&lVake`� h[U)A�$(�M��"����͵"�� �W��^Q����5���I�l�[-*�0�ehڭ6Fj��[2�$�%�0)��f�h�eSjh)��Ʀ���"�[4$ �x�{j��m����mCl���2�L�cmXۑ��i�R�]um,��F�m�dmX�ٶ�ҁ��$h֙e��ճV��6�V�kj،�F6��,w�eפ6�b�Tܪ�   �θ��B{� v��k����Nٶw2�[�ӆ��iѠ���Z(u]��S���:�wt���]V��6����-iI�  t .{ER�=���t�Pl�n� �h)@��l�Gvn�h(Pˉ� t�X;��.Ű1�B�J��o� ���)�m�V���m��mUN   5���I׏xt�4)K�k�:� )z�{ި��Ow%P�J3{{΀u�(�/sRR�}��}�m�!m����� B���t��y�G�f�m�ki��*T��o   ,�:Um�w]�=hY��*�׮��*z7�o<=�)���������P;T� �Jq�qף@{N���K���XRMi���fڨQl� �  �by@
]';�*Us��*zʙ���<�yx�)��T��z�����[����T�n=h R{��iTPmy�J�ֵf�ժ�[m����V�  �����k��z{ z^��P�{��GG!&�QRw6���U��m
J
m����4-�8҉(:�ˮ )T;l�vj�U&ڕ�����
���  e�� �4��9P�֮�����Ln� iSW8:V�MhwunХ
T� 5�52�M9�  ;�� �՚����T�mB�hi[Vm��  ��r��ֆ�5�5�4v�� �ܷ �4��P+;��(���gP�ۉ� ��e@*�v�F���X�5E���*�x   nw;�t���
;��݂�N:���� \�� �0 u[ K�[� e�L ��wZ�V��ՙ%�e�kM
�<   � P '��ցF��s� ��� ݳn@6.q@ۣ�
W[� �x  �   �*R�� # #&&� ��{C
R��04�00���{Ԥ�R0      ��	*����&0   �{��)*z��H �#L �hh I�T�z�i�Dd�F��A� �ښ;z�����~u�ڮ�懺��ݝ�7o�~*2��Ϸ߯{����HI<����`$�HBIH~� �O鐒I	'�&'�����a������I� �I	"着��N�$�O����d������������< �4`O��bђt@:0���D���I� �t@:2N��$����td��'D��I� ��:$�N��'F�	�I�$�����$���!� ��tI:$�'FIђtH�F@b@��:0���$�tI:$��tI:2N����#��I�$��!: N���I� ��:2D!�ćD�$��:2N���	ђtI:2N�'D&���,H�рtd�'FIфчFc$��:$����:2�:0��C� ��@��@:0��!��,d�N�	!�! h�萐:2HFB@� tH:0�N�$�	$:2bIt@tB:0!�F!� @�$��B$D!�B�р@� ta$��HtB:2HFA� D��ђ@:0�$�@� td$�C��!: :0!FB@��@:$��FH@萀tHI:2@� @I'FI ����@�!'DN���I$�@��Ic	!ђ:$$� tHta @����I �� �$�$�$��X�I�$�tB�$��:$�N�N�N����$�`�'D�ǣ$�h�:2N��ђte�N���$ђtI:$�D��	ф��tI:1��D'D��	�	ѐ���tHtHtHtBtBtd,C�Iђh�tI:$�'F�$�td�N����:2*�B�sPa�?��Q�n|�/)+�ڳo3���������[;ڱ�L���b-#�e���U�SY����f��Ɏ�9i���^4f���<��-�F��F��4��VU�+r���� ga[��t�>,c�8�Q���dݘ��K�ȱӺ&��q�^G������c�8#x�x�4���ד��p����a�W^��r���n��M�v�v]��]j�[:��7ǏJf�A��O��p�_^�Չ����`Do�c$�YXs]� ӽ��Z�lv�ڙ��s�bo���I;N[:��{����X��6u��4M٥Ȱ�1n�h���H���%)C5 ����(�R�EY%�Y���Tq�z.Pו�DvY������+S�s�;W3�
�[�a�s8�2X;R��R��LZ�a�=����&����n���y�n�ڬȶ��G%n��f�"�X*��1n�pRt�ûg7�5�؄�o˘E��桐㹽�.�4����˻�ލp�c%�9�)WʻM�T8�Ӈ��R����$8�J��q�Pק.�̹UF�`�hT���ܲ�wX�l(��͘Su���w+	6F&�n��r�^u��%�q�N&2lO�y����2��[8u�����"����[��[\� ]��x@�&��zhm'��ki�#`��#b�Lx���ã��;v'����jv&8��2�.�)=���ٲ"bi�j��&���^��㳦7�r�8�Б-p{��kqԏN�sv�Y�j�MJt�ỡ^�G0�$]��E>��qwM��z��[��ʤ�U�����ǤLՁ
n�d;����R����{+%�Hͬ�M������pN���çV�+��A��)S��{w{����Ք�|��7����T5��s7t���Ԉ���G;�sF�$X�t��ތ��W[��eѰ6�8���^L���"*T�Xt�F�Sc\�%�^wv���d�����K.��� r\��U���Ъy�h�����5+T�A㖦ݼbk;�H�MgQ�ԝd}��nM����p_w�[���Lf���S`f����2���o��x3C�s�
vV0��qVj����m���OU���sq�Sv>�%��^#Rg&� �*�]+��UZ!�U����L��:��n��V�������ӮJh�E���X鋚�U�k#	2Gi@��k�}\�9{�*�ڗP�Ɠ[�l��U�w@�!�v�$�����w�)���)��ߦ����!qGF!�J�#ǏE�i@#p<Дj�Zv��`U� d�G]�{փ�1C���=��GP����7��P�wiX��dU�V�Mz5��I٦�������s;I�/ۮC���i�.7:2����d>�!��薔Ov��0����6�5��͔�m����V6��2mdn"���;��rMpj�nƪ���݆X1#˻�1";.M.�yD7���X�4��8eƓ��s��DE��/l��
�6������,A|ogЖ�4�����k��S:�b��T��pn�,�������hQ���Qtt}p1������
�*����53�v]�Ʊ����_]��r7�j��;�&����#�r�h�Ku����T�#{p�[b�H�����8nk�1�k�V��%��=�����{8��S�2!nX��z�4�(����Z8�����g+�,3ҷ�uM�wie��2أ&�M� n�͔Av���ܛ's�1GyYb:�x(��A2˹z�]��iR_=�O]ZD,w�۱�0�V�E�}�~xwg*�B�o!��M�l|+�tG�Uu��â<,m����i���<A� wRƫ�!�B{��ĥIF�2����w4Jkjz��Y���!�1��a�;�aW-'S\����I}�Hi'������Fn��l�v6�u�����ĜE�\3y���k^]�#�_ٷ��ϝۯ���IhCNn�1ͱ��NI�ܒ�hδ$-�q\G&�y�1k�ӜN��Ib�7�x'�֫C�j��L<�X��^,�܌�%$P$,�Q�/�ms���R{R�=�21��E]�ӭ�_���k��@�M�+l� b���-P������c3:��8��*��%}��;z�V�\�W&pX�&�5dL_�nf�'u^mխA�inY�f+��P�|���O&ɴe{�i�TSنlD�(L�~u���^�bSsqQ����\4D�G���=H���U�ŭ����)llO���C�kYB���f��ʩ���O{ab�'�i��	�r�8b�e�:s�(i.��4k�9E�Q'�­��`���6��{1�:�m��6�V�V���,9f�4�p�#9	&�GU	@�x*����P�ʹ�����#�v�;��w&�g+W���N�׶X(Q�&k&V���x���p�3.om$���teg-I���r����C�A�;���X0,�nQD�j�6��)��Z��b�9lG�ss�� ���cL�Ta�wwʵ6�tm2�ʂe��9P�sf�f��GH�вwa�r-ݭ��sEk���4���Q�Ơ/F�%ͫ��֋v	om}I\���1���@藹�77ys�!�B6tRnZ�k�l�@�	��'�k5�W5j�[7ח݁ޕ�X�-����&&�!�p���nf3�'T��l����*���n�p�ek_ L5�;KԹ�ק��.hh�,Z6oM�&���A�0槠t�Cc���m�7��i�3&4��:A/mè`���;O�U�V���Ti��z��X#q�8^&�)�x
�W�lMYάno1����ץz0���
+�[��Њ���o4����@�FK�0��_����ȃw+�u�<�B�
����������L���M����6=��n)��H�*H�D�F7.	�=�⏎T��~�tK�0��{U�̈́�c6dGuuN�R��,v��T���b��+��4!S����bos�Ѱ��v!�˖bwC�nË��a�m&��we߶'�9☡4�+=ַiDV��� ���Y�*�6Y��.�k�ԴJIt7@%٠�oӒ��$�Q<cuaP��m�0�^+#J�ڳr�;
�gq��Ş�����Z����0+��%�+kt�w�i�F�l׍��6�A�%���k�4�-��x.��4����˻�]�Z���M���7X17{��w*�I�ĺV�Gx]h�g�l��GT����&ꃛ�v�&sm�-SNǗ�Z�\�[�v�޹xvս�)��2�w{��D!�W�칰�HjӘ��R:��ۗ0 K��p��y�޲`$�ر��,K�
nZ�'{�uy�lK+hsGrn��cs�`��5�>8<�>J�Ia���Sfiy[��N	aL�t��{
9J���*�`��-�{r��xQ�.|&VO�9�\`�sfv�ܘMUp않Pd��ZXźH(��bݽy�O�a�`6���q˲[6��L�<q.V5q�*�׫����[�H�޶�O��R��'��I�Z�V�E���k���ᖨ��>�8h[?Mp��J����#t�A$8���<y���Z3,Ve��G�X�@x���v�n�y�Ó��Ƶn�T*��B�����v[�V蚦�=�-��ޭ�ńvI���cRz�X���;6n^|�è�z)�r�eՋ��%�x�o'9��l+���|.�$�K��N�$:֮:xq��&����<�v�41g:İ��՜u�ܛ�$��j�,�t+h&d�Nf6��u"F�ޖ�t��DF5Źw�EY��H�b�[8�Ě&5.T���Ƃf���$�̙�m�Ҡ���Ae�ڌ�"q��߶dc�d�͝���W`@N�a��js2�a��F^�-o)�gw������+M��I��\z�S��$ۡJ8l$��:Ҽ]�Y���݊~�����g�.��%�Ƚ��n�NkD��sQ�8�%�p�6b��c��I�ynL4_��Z�.��������S�r
g�����,���%��wo�e�.�\��)��-f�����L�p�WoL��wzA�PCت�=�M�s1t@}����i[;V`RS1�t��gz=e��&��S��~���*���Y3�W�d���f���Ol�&���.�gjꞧ�}ħz*��45-�T���2%���^c�P��N�i�kx�ۄ�Ǒ� ���͋l��8ѻVS�v�F�:��!�3�L��	�a��cd���yYw\�Ŵ�∬t�l:"�ͺ̢�Ȕn�[��P��k'l�G^���-]�7ڣ�ea,��@�ԙ��n��")6��F�h!fV~�{Ρ�n�[oa�ё�����n�nP�j��$Ob��h���Cr9IC�J�؆�����K���;�b�&�� ��Z{���L3�k�R��	�z&\T��+A
&1���ܰ�O�q���2���#5#{yV�i$-,uE1F��e�Lj�I�0��e�G�9(��:�49~4.��T�r�Bۇ��0��}�Ρ6e�7�ƺ=���>v�c�f��U�*�eT+�y��-Z	<f�ߥ`dͽ��j�d�ٵ�{�7�6L�+ڷ�x�6���5�"�ֵy�� 
饶�km�O�{X����p����v���2����+#�g��=�;,���#Z���=?=;{9E1G�f���y�w7�S��V�qnE��)��ȧ9.�L&,;t�N�D׫�;Б��UҳP+sV�J��d����A��ءI���F�9�3l ��%ƻ�n�V�ۼ6gt�����j��8���G��K����8p�v^��w,����~p��݁�MяmYk���$�8k^L�;!!mdǄ�7.�vsKOnC�[�s��'����;6r�ӂs㦻�25b<�r��4�*���~[���кoj�y+��Æ��w�އ�X���me�g��zr��EQ�[{�&O]i�.�|�m�j��(�ɥF�
����pCFU�!X���kh@�	��\��0��F�`)���*4r�.����ty���V��ӊ�&=���s��HsE�Ȏ�ls��o�%���Kh�b��9f�3��i��ḿ�j��v0�EƂ�3�9}��6����Cm��,�hɢ�5�s�E��ԣ��ѭ��1Ƽt�����!�ӗ�A֨
%�{��be5��K�,7x�I�yfLllC6�z3\644�ٲF�{[$�mk�6��1��M�ܥxR��r�<{��j�'	@iظ��M�ň�ߴ�9�+�yW3��"x�2ot�uh�;�a�7f��-Va�'u+.S�U5kI�L���I�0�]�@�8�Wd��� ���Ocrm�nU���vn�����hq�������̸rs��)P�^;����-�@�.���V�u1�ˡ����X�x�kɺ�T�K���ɕ�ib��9K�:�!Z6�D��9��t��Z���kK7-L�`v'��+p�3c�!	�0�Em#Ҋ8��)�ûu?�;�N�OnP���Ҝ�1���7/7�O(�,����(n�%��vuփ�i<�"t-_NB�%gU�9��`�A�̃�(�z�n=��kߴ���0go-�� �K�K^PYĴ�ީ���f쏣���:��e�@�����nE�&���1{V� _0��x�%u5�Z��M�me<]�rL��+�κ��c07F.�>kn�jy�	��*7va]����BA�A
3�Ut�^G��8��F��f�6��Z6I�Ze =6� �'�Ga���,�G"׵�`�l������Y���� t�vϑ��+S���)ܢ�ڸ�w�.j_�2/2�+/h��8܈�bJe��0�J�{S�K˷�O�s0�0���Γjż�C]�j��mr?;�p����̭�K���C]I�T�1��Z�s�H!C7 �ܸ|x�{�4iYz.�O@���u�ެ�
�}�c�U�9q�1�Փ�9��amۘM�&d�e�ݬu+Y
��"v0��/Z2�tĨ0��?S%��k0Q�4Ӡ�0����`$�A�z�q����n��2�r��`U�%Yܸ32�!qV��n��KҤm�k戚�B�1%X��}2�n��ŧc���&e�9[�+oC6i��[�"���L��u�n��ҵRD�c�ʕZ�����9L������
�tݷ!�S͝ƭ�5�6Uh�\��_���4�}��Q��#r���`�ef\T"�!j~��l{x($eMzoov��s�j�w�&�F0*����u�f:Nj(]��ࡻR��l|]�9����$rVw5>ۥ��QAJ!�֍�{'0�[hy� ���F+kuݱ#��x!��;�mdQ�R���n�F��J'��|
4!�YHy,tC���'!,�D���� ��W%�t\ee�&I�a����1�Бl� D��Yl�Ϙd%� 谩l�@����\툢��)EI�>�YX:��		F@��6���YREψ�NA �DixT� �t`-6Eش�9��1E��(VC=А��.Ȳ��#ID`a�$K=�97L���.�
�֒
06U���N�֎�Š�$H�]����+���	���b����Evz�t�}Da:ZEP�L���0�9�A��<S�1 �h`����X�ie�	�(L��EI��������9eo�~�?��=���[~���O����]ϷB�g0`$ -�j�hSg�D]��g-����v{�TtF�#,��@�I�X9Ӯ޸ռn@5��T��������i�9�`;�������f�Yis��ݦ�]��]��\�Nݟ��6aO���Y�B^�U�f��?&�����(��d^�R2����T=����l��SiV-��䖃�i��{�ݻ!O����_��۬.g��#C-�$�1ے����8P�U��f�� ����t��~���W]G��g���\�/���cZoB=l�n����V�Ye�^��y��4.ݙ�Vr�c��H!���(���[u���3;����HX(�c��EǍ<�ɡ�1<Y�<m��+}��[�i.�u��)Q�JW�zS���|� ��/_<n;h�ѣ��;�7��l����|Őo�5�GG�4��A��j\As��yB��pv��.�s���Ez�ǲ�f񌰜y�}�؎��:�4�f��q-��hܓ7Ht���A�Y����9;�:A�	�������f�9#ͮ�-�(�u���e��OmA�ŋ������m�Nt���tkk+a;֩�����})8�Ə=���it�z3�P"�̺��|�ZͿ=�cp�����.U5��a��*���w\嵌f��a~��nj��Ɩ7\���{'����LW�xe0z>���p��<Bhi"�M��8˾��vh�>ǢRN�|&��׸wR����5�}3�,^�0��{�����;Ѡ������5.��pT��L��<=v�vƳ
;�`��{����/�	�=Yb�V�%|�E�p�^c+�;�Vtb�rQ`�	�[�Zf�_6|go�k�ȓ��M�<���w|���Թ�K��]Z�W^\��w3ٯ�����v�{V"0ʵϯ��Z.�/���:�o{�r���1��V�-Lu�7���>���Lƹz��$��n��T0��7�@�r@Tz�W
ƒ&�J
�sr����ܹ�a��C�V�?,u,P�����f����2R=+$sl�֣��}�p=�<�����}J��5\���D˒��4v
��t�|Г7��7	�Ϲu��i\�;�ܛp��8��'ޞ�w��;��d)^�+�,�̲�;���sw_�l��ُP�L���8z����{�z\���ϭj�z�Z���M�j��{�J�q�9F�q��T	�ܕbYwƸsZ��3������������9Wṻ�1
=��3�9�v��!&���ݍ3(�k��D��=@���<M،�6��w��N�M��N�9�z�V��Օ��f2�]u���[�[-��3��nV I�R��97/����3zuiY���Gg���Y�ZF���+;zqu�Ο�p(�<w��5-���#5�^�6�K��|sb�r\Q�n8:��S�Nt�����dw�cȴ���Q��Z�N?N;�+�I��<�-:��!n�]N�w^k�9��#�x�
���:� a����_l �+�x~yջ9.D�ޒn���]����I���#B!귭k�o�
Ô�x����+؎��WVg����x�O,�i�]�~����~�͛_�L>qz�t�c>X�����b^�Ϥ�&��wG\�O5��/�w1��F�O�' m���p
c�}����!d"}�Z#{��'��S4�+B���L�Z+�V���N�G�,蔀�HA]Y���:�ٶ8��KY����٫gTwh��A�Ӕ�)�y�u�k� {H���]~�2���<�?{<٨5�O��Y16�c
�r�7��m���,��ֽ�C�ǧ��U��d 9�aGT��Ϯ�4)��]f�hh�\'R����}��)n'�r��
�Vn�1\�۴�M���ھ�viSm�+�cɜXy�����DW*�g�dLj L��[��)�c6�Bs�%ڠJ��^��zf�;�։�0,P���kγ�q�X9���z 0s�Fq�'�9��^�����.�3#�:-L=s�����\+�DgNR�bpl�u�?D�԰v�,>�m��s��C�˕!Ü{΢�S5u�a�&۳0�f�g�J�����Z��v�5N�I��؊�^Yֳ[Z]�5�&��*�ŗ���o�1H�Da	[����eּ�et�Wnc��JyyPQWu+�ʻN�����xf���j��
ú�,����MՒ�A�GxX<F�Z��n�����VF_��GOn���aO9	�@�"��E�_���)�*P%ѝU�a�uY8�]�؈������_�~�2eJ����:�4�6������Ӄ����%�:�S:���f^(Fd$�"ypá�E�7�n��{���4�L�!�$�֍�&CF����MޛC�;�#�nų��d�[uu&�7)pda����1�2p0����2�SƠ���b�X����V���:�ww�4���p=9c���+��ĩg��S�7�=c7@BW�Ko�>�|z�+}\He�X�>u\����[1i����v0}� g�\�Ŋ�ج���y:��KrglUf�3# zPtJzog���q:����禿,<��U�|uj�R�+h��� 绻�f\�����a$� ���T�m��:�Qi���eM�{�tj,���W;�����s��.=�
+"��pL���u�'<p��AJl8�uNW۳��[�����5f�B�����1+�)@��(����y\H+�U,�w�HI)��i��p\�S����w� /1������Xyǰ�:J����vf)���uÐ:���*|�J	R���f���}xeZ�f��:K2���+Ol�z���<�}͗},O0�f;�9�>�+��Wua�^GϼW���^�8�b4�"b��ɧ�ie��3����ɿ�;�FWt�]w/q�n�<u.Q�͵�n�b&߯�|'�䤫��<���*ɀ�������ȽR���֣���pݽX�
J[hnhkw�r����2P���E��^��B�k-z�\�˻�(�[s��*�C�^t+��v�(�uG��A����J�5L��e,�|N��"5���xُn]-���J����j�t�����*%)կ�v�����[Ag�'�<^^�j�.�֨�!L#��y֪��	��Xp=�b�a�6��)6����+��ݭ}����Y�x��ȶ�����.�M���,�*�v�g��>����	w����n�'_nA]%��@w/������u;~<���x7���R��1���-ل���ʳl�S}��	'm<�Gx;Q�]uܷ įP�_u�aD���W\^uL��i�ڄk>�X�L`(��q����[�.>��B�y�q�]Ar�gt�Ք����g�'َ�o]�cL�vF'�h���0<��3=� �0�~s��}�w	�ȸ�A�쾌MJ�6^Ѡ��G}̸H޺}�_���N%|��S�����2K���ޥ�v��UG�T��m�YĠ�&���sUeT��L=�W�.edī�7Ml:����@R��-��	�6��u	��p��vQr����9�:����cf�w$���E33#����r��VۢDĸ�ASP�W��S���q�j^�I�cAKhY;׫{��B�ܼi�;!���EIՐ < +c�l{˝$(+�Bv��E(��e�0�/���+"5�_�W/0�'ܖ�&��*�x�B����1�;qu�a{9u��79�=u=4�5��s&t�%"�i�c
���Y�;��e n�1��b6f����m-�AH��*�o-6���ɗdNW@m�[}���@:Qu��goM[/]bWh��>�)�er��nŸGb�.��貋�Nv��ۥ�$��o\�_a�R�t�׃;%�����-��{����Oy�4���F����,���1�æ�v���C�݌�pK�6����R��h���缋��[z���O�|qG���E�{��O{x�4�ӥ���r�X���u�E���MΡ�9�Zל�A^c58���}H�Ɂ=���cޏ)a$�л	�^�/�:���z�hl���;�[a���t�����L�0���Aٚ���u1�=��8����/�,vn�����s,Ir�u�2�J�ڏ�v�`�$Y�;���M ��b����my�ЖܭWb�>�̣0t��c��ʷ�{jÌ����/�ז� V@����18�t�y��o��h\�J;*��N�IY�C)�����Я#�jv��J�E��5���f[��Ct�|�
nގ� ��K|�C�he��3k_(�����$1kyV�s�7c_|�$QF|�˟h§��ܞ�x�� #O�����i�U��e9w�a�Wm�t��=wg�M&�i��ζ^!YCZ��Lf�M��P
R�y����o���Y�*�6�y4�_�p�|�qjK�:�n�&��I�q�u�9L�G��lǶK�ҳwF�!8ܼ��6�ݑ�]�5=rwQ���7��h��\�U�W)�+�lfvڴ�����[�R�8�*q=�(E}����f�:�p���	��X6�z�ʪθ4�@�,�v��*�N�;<u$��a걘��F��*^���ʓ�%��c�f��դ���eI�O0Vi�m�ʄ��tg=0�}ׯ��X�۱�A�ɗ�nV���1���}*���R�L����M<��[z_2|��=�'��<,��.���T*]�p �y�	lŷ��s_5�K��x<��G��o5î�������fg+Р�`Y!Q����'l��n�3����LV��HmO�-()շImeDk\`|���Z���i�8F�ͫ�1���s@E<�p-rᲅ]�)gi���!C}�*����+�γ��ف�1K�~�K�8:)�M#C��g�W^�+m�).ޞ]h+F����-������|���`�;TQ.��D!2����S�@�[�9��Zyn��L��hFRMB��wM�K�}�{��H"�HG��է����z6r��d��6Q�B�n�t�Mh�ݿ�Gil��{N�ss���0��*����#\�q�ѺAC���;|$ݲ-�+yR?��+ZU��s���V�S�`����m�;��xP�u����Qy����������˅篗�7���8�ළ���PF��.�hW�n�;�ɗ��k�Y�V�}�9�YC�?R��ሖ�5��;V1��^g!��*xL�C�h	@�q�3���1oB'B]iWM5�Ë(�ns���`K�B�d&�<ܽ%=F�]�F�ݱ�3{Iϓ�m�̗����&�;	�zq�7y>ɚ�ƚ�pZ:I������㺽�l����QB��n��,��zx���Q�x��o	�t��>xw�W��;#�3v�T^�3@�@D�ܪ(-�L���V�js�̱�V:a�Ѱ�M�puaG$]��QlY3x��d7P�+�N����E))S�չ��n�x R�aE��W�n����Ҽ�xG�d3=���|JE��[�c4��V�x�5�/���%�U�?�=�w��/Sj�̓�wCP��8:^mWz�B�L=��fױd�ٓ���ū�6�e��R�z��Ƹzy�.�bL�k_������nB�sH��v�!�v�7Z���9+�N'�4�Ir{x-�ج]�1�y�F� Z_{�;�ޑ�í��oZ8gMN��Eޑ�([�@f�G�����F��yu��bR���t�� �u=f(������9v�&U��b�t��B�U)yu�{��~��<�3���'��O3A��{-���*��X��2s�G�����)ca����U����ho$Ҭ��W*��@+-G�Y�;[zev���'y9��H�T���~��_>�2v�a�o��=׹����W6^|�=r�˹ڹrŻč�rwK�	ˑ>�.�֡X�����}��{W�����g����WT�v��l�l����^ҹ���vy`���,���=�t���5Z����NZ6W֌�칻S��>\թ����fC.�5��aA��#�m�AC��.��e���t=2��T햟me�9��otJL�i�a;޻���Ũ �ަ�c�c�5��Kx�sǖ�2M�wQ�!mҳ9|����|zg��*x3[��z�c۞�s��8D�ܡa>�A��]bq%A�),<+hc�L� sz��/̤)D�+Aש�3�a����nv�º���'xވ���oM�����,���57��v��o�%�g�i�/��V����7�H�v{]�]u��v��R�ܬ����q�>E	�h�F���Y���c�j�Q�;�T��9G�w��V��=�!f��71G޹���)����E��t�S�ɛOz¹R%������R�9V왪�Dnؖ����%<����3|̾�n佣�[Y�;��e�oI�b���?�!�l��N�n������.�:l�¶��[I�$�+��3o b &U�N��8�k��^I&E���s�(���0��(���&�s�`��^��o3���4�rl�$�2I)�-�"�&��9Z;�br��ܣ�ݥ�V7QNP�mM��=�[�՚6m���f�����r!��}��>[�s=�}�s�{�C�9�9�����%d�$
��!�a�	�&H�!�~`�O��H�����?��]	I >�?�������$?����!I���?� �����������u��ݱ�;���1��(�)Zx�w0��ݯ�4��ETʒ���+�x] LޱC3�yك�H�X�2�cO�wV���f�i��2rV
ŅΩ���fm���v��f�	�n�x�ڰCv�Z$o�ک��`T� �ї�ZJ���b\��޵g3�*�|'n'o���w;��6�>Xa׫��ܼ�-<���O6��ε��=VKz�A�a_�P��m:5|�I����T����?*Iч�CfهO"�����wOa���T�j��ֲ���rs�;r�5x���@�Mk�!ƚ���އ�75Z�p�X��c��N�z����L�E�8MΚ�=� �s[�N2�ՃN�ї��..{�Ϲs�q��0��WG��H��gg��h���h��<�]պ�a���E�t�G�d��%G���R�wy�O'����C��^OK�Q�ڃ�c�b����|����H�<��L	��x�Q}y�|�}��eW&5F������/Bz�����+V�R�T�]mj��4]�r}U}��b��.~�g^���#p<��^��{�x�zz�a�֥D㾖h)�0aù�LT+u�!�G\�6�����v�{n�WS�z3��GsY�{{�3�j��u�N�1ɞ^A&C�{5�}��z	�{����;���n��Z&] #Ƕi�}/��w.C-�l����:7o7xD��啜�+��yv���/����w��������{��{=��g���='����=��c=��g����{>���g����{='��{=��=���{�}���h����X��ܕ���ܴa1k���N��l�aث�+�GW{���q#��Y�ز*�PG��L����\��x��|@���-䗆E�{�b����\f�u��f.}r��"�c�@��o$�ʹ�vv�n��j��Ryٷ(����:��W)y�>-�/N.���>����zi��$e69T�:���LK]�ݔb�.&�����Bɇ1�������8z�6����� �vq��'����\�lC��yL��e���U�5��V6v�MZ��s�Qt�;A�p����A���ێX�������C��44x=�n;��C��E,KXX��Ԭ�f���zM��6��)>��]Ħc�]��-k{칗wf�˝jt��w��:h�Z��\G'Ρl��Va;/��4g�}y�T۹��X�N��	��*�n�Ǡ����oXX��}���9�ώ����b᧊���|q��Q��oZ��}{Tt�"��M�#O��"ŞH��wAX�rNvX]����ܫ��
�T�j��{��sz�ή��,ٯ��B�-���Y����b�����٘���͕i�CC.�%H�tGs� �<�w3_;B��+p��������A�xڀŧ�46�S��i�ub+�:訅� �ʾv��]7=��Ϗ���ˠ�K(>Fz�����>��'9m!ʝ�#��~������z{>Og������{>����i��{=�'���٦�{=��g������{=�'����{:{=��>�w����}>�w�����nS�$ƌ��z)Nuр�}��c��)�w�����S��
��el7o*�������%����W�%��R�g�D���|�(V�"���{ۿ�j>���,�)�^�z�!mɭcW�QT;�L)��}�O�v�W�}n��̺U>�{
�ٲ%e��f��l�%A��x����7�O�+�[2ӲbSP@�z���TzdEETX�t!�pdj�f���j���R�]�l]lc����7���A����9]�c6�S��/M	q��0��p�o7���y��Þ]5}�6�b���|�w����i���𽮚c���s��2��3��ԑ}-��-�g
Y0}��X���p�*in��˫��]�z���j� kj��1�mO�a���U7fm��~b�د����4�9�;�����xd���2�їx�a�1��pr�'&E�����&a�ə�xy��C�|��>(��ܚ��R�k��K�.�˷�YV���WX�6����iN�y�"�D�fۃ����gi���e��3��/� �FXkc���Ŧ��9�8/P�y+r������gpz9P`���~�䇙�����2P)Z��:`��-�~��|z�MQ��8�+6h�����{bȋ%7D��;����G	�W�z^B�#����2�E���ݹ�f���#�Ӑ���_g������?O���}~�{>���g����{=��'�������{4��ӥ��g����{<��g�Og����{=�Og���������{�}���i�����ڹ���>���t�;��tJ^勻���|�ݝlϨ�|Bϊ�V���]���ifI�uJg�ۼ�|.>.�.�b;��V���T�:��X����\ƅwJL+hśVv@�;!�fm�����k���m����X6�%]�����S���ٜ����ME2ΑhX-h�+um1:a^W�v��b<�ËǗz��ټ�c�<vt���e��a+�Z�&]��յ��.aD�m��@�8ݻ͇������5u�RuL!O��=�t��P�7Y�F��{j�J����p�}i�U�c�`����@��(������D~��Ӿ���n�RٽL!|�N.U��s�S$ �@��Re
e�t3_	y�`hm!$���9���3N���*�8"�;@�[���.mn���te]����}EJ���.�2�P�4H�R����h�`6�IR�ѕ��!+MꮆE�������9�U�vmј�>���|Ig�v���A�=�SW�p����};3��C�1z��畿W��+��9{K�u�eA#�����E��7klW�S�
g�l���y�E��2{8o���|Q#z[q�-���N����7��)1w�B�:�y���y��O?n_0��>3��&���E���ù��ߎ�1m�A`7'{~}τ��>����Ϲ��{='����{=��g��{��{=�i������{=��g���=��{=��g����{='����{=��g��ן'�����r.j�i_�����ڝ
ͷ�.� 6)�����(�m���>ɷs��U�3���6��4��b&���E��cH �k���4&O�5�vo�O}A���J�9�!H�
6�*ri��[O� ����piFo��t�0l�]��� �Z:K=�a�}��~�q�[��qT�q�ҟ�i�8���(k�鈍�e �m�ۏ:L�(�q<n�|x\�-�#/�p�P�'�I�2���U�Gأ{�I��FrC���dT u�r�d����܋Tޛ���y���Of&�R&ꫛ�n�H��Q�_����w�����a�#�ʱg)÷��u��"��ؖQ4�ȿ��}�ub�{~�=��'R���ٛ���k������ހ3.���E����/N�D;��T�%zj�}3v�1ʵ+��U��.�etQ8���Ow2P��\�9���ɯyI���7J�aB��{����,#2�"cxE�Y�'_g8T=��e��c��4��aF����+Tp�
�{���������._X�4;��{��F�qײ']kYz���xv»�V̔F�G�//t�3T�&�&m���;,}�5M��f뻎�Lo glvn�]6��/��m���GiyB�\yV�1��Qs�r��BM�Ȇ�2���;î���%m��	;�ڶ�۱_�Z(�ն����z��A����9U	BsG#����^�!�I���Y���O�}���:)Ļ@ʝ�)�-7w:fe�t�]R*�\�T�
�qu�QΫ71�xE���FG����L����5�.L�Ł���л{�X���2�寄�U�Opg���q?&h��j�87��f	���K�D3,�B�扃N�ߧ-Ж��V���S���u�����lT�pw�כ[#p�|x��~&/;껮���=h;�}��r��3c>"m�;��죌��+F7iEGH�S�����v���KtG}�'(vI�Ki1��+r4B/��xt ���>t?�L��&㜦���%]|sP�n�ef�ͨ��MT�ځ�@gb���I�tw��"#� 0Gs`f���+SyWO�.k8��kc{���㽳j*����pK���W��KU�T ���=�i' �5h����ы�~�NY����:��xDgi������yl��
!��6d�*�I{�re��ᤖ� ���B��c�����:2���I�֨!P��íb�3�.�ԍ\�m�o����x�94p�sJ{�݊��]�U�3x��WK|����D$&6s����G*lMp���sRh�Y=O���c���K9[G�����W{���y{�'e:��R=C����[�ɇ���g#�ί/�_NV��j3�{�ZH���h-�ு�|+z��k 4��9�����I�{�'�[C�nL�?p�n�o)���̣8���{����/��q���ֈ�`ǷIVQ}Yu�@�`t��O�{�}��i���砹���$��;\���7�����,�&j��r�q�޼w�Ds�hp�{Wg|����wv�,���Yv�"�ʹ}��a=$��ٲ��,�\���mQ�<��B�n�M�_���N=�y�za&qc�ރ/C��7r�g�V"�p�����`M.`�K��}4��ykk�tû�=�k��Sg��������33�^��t��*�"Z���i��� }��M	�Z��Ĳ�$�M�ڳq�D9�Ҙ�=�]���/��v��,��q\�X^o/u��+s�5�GV�<F� �{spn`��f�K��{�k��:�Į�*��es�4B
���7��k4&&�\����t�	��g�K^������8�6��b<�C������4��@A���$�)�.�k�11;��K��Q�m`Z��l��1����ٵ�\Yr��lQ\��B���	'u�0�|�%�X{�vB�[�N��J3; S.�*r�8�� u��;>|�WX0X����g�`T$�N=�c���*낊��ί3zou�ݫ`B1e�ܹѼ9YӤ�
˜b���s�?3�����@M���l��}F�[���(�e�.Nޒ#u�%��Yqn3����"�r�̗`b�歫td<[���A�=��F7�ԥ�)�Q���DD�G\ԛ�rZ5nߡO��8���.z��1�O<{�qs��t��v��ڥ�}8�Aو�9��,U��ٮ�m�-$��,I��a����x��1٨wi�Ԟ��n�k(<?�f�����ʻ0��&����-j�%ΆA�(kK����lY�_��>�B�]���A���;�>�n;2f�3���W=p��xR��ٸU��S��v������]�~����]殮L�b	��FH��ᴽ��|MRy7��h��;#kra� m�Mx����"��H��+�㮬��i6x(V���#��E����w�f�Y@U���,��B�<Y[k���˸ﵐ/���JE1�*��gv����!�Q���o���CaC�J
�%� �`�5�K�������ذ��(�3��0��q>���~|�:4:�'�3�+��O�.�J'8�yɐ�kP٧���/��unUX�����PL���M���}��;m~<ϔ��q.����$	4��{V�u��Q@��Bp��y´h����5v��y'!~(���!ǯ/w��O1^�{��C��q{��gE,gF�u�����7�l�����Z�g�lx@˔ �_3 ��P>hJ|#
���"�����wZB'�0w���U.���r$Ԣ.KˣX��d�:�v�Om�-�ԑP�5��^7㤫�����s���E���+k�w���Qi��}��]g^%�kz��[ۇ)v�޾u����&�I�������+G^nX�C��t@	�4wG�**��ߧ<��Ǿ�r�6�����!��nD,�r��Y<9�]\3���Y�Lr��pە�u�p�_U��O���a��X�B�=�6R',}�L���
����q�Z�J������E�a �y��"L�=�9��Uޚw$�;���[3�{�Sd�dz��N��]n+�I���a���Z��x	aԃ�ɀT',�c@�;�a��Ј�M1����5�}[B&]������3�ug�l"��3�uCBB;�(\SP�3xl)v#۸@��p�8�f�G9�hX2��o%��e�/�6�,���ô���v>�I��uL�"�Lu���8Uf4��Fem�ד�&����h����]��1��w��x����D�l�&l�d��2��x^�շ�wC*)�9�ykP���C�TՁh�w��<:2�|�#}�����d����{���f�	/���c� "V10��h�9���l�eA76mD�F덆���J�.�C�x��āH�)<4:�7�JEI󥫎�G}�.���^��d*P&��Ɛ-ov<�ZE�LwV>����%4�ҙ*�4�k�D��yݷ������J�+� �A+{MDG'�Q��|t��op�X<(�pެ�!S�z�!�'S��`�
�/^Y�6�������y������m"��]j�Lu�sE*v2.ݕ8�L�Oͩ���txW��x�a��Û�ǳ��#�|��\.8�v�z��3Y��|�}y�u���þ�f�k���q���1�AL�	l���*�B�mѹ-��9�a����
��
�\Φ%h6Аmݗۡ��3vT�}tDHm�6��C�Y���u�p�|�$ ՞�@�)�|�5p�gZz�\U>We.���+��U��@p�nȴ���.�q(���ȝ�'Ozyc�����c���n
>ѭ�bܤE�;/iQ<�1��LR��S呝˧[2�u��tw-(�/Xt"�}�C�!33N3P(U�)q�s(T��|j�/+by�x�/5�\4�{Q1�;�,!���\�,���~|��i�%Z���C¸9�rC���@Jq{���j����8m0B���7�8��Ut�Z��>1���n��UD�C�sP�����h|��=7�7����z�ݽ��w ��4PK/�D�=�-���￯�|������HI$$���c����-�q�V��o{���Ok�9��Be�Al0Pm�s���!�Mf�q�\��� �Yj"�%��Em�A*F�I����i%{�֨��\R�kv�Qm��)��Wm�k�/�7§ta�w��Ί�}1���l�v3�,*�Wh16��z��G�t+����Ҳw0�P]=Ǟ}�>��D�`�PC4�,������p&�����T��������������3s��)��u��rm����Hnd� ��x��ٰn��]\�S�Z���MAH��ɸt�}mV�L�Vju�=2��'�ۻ�=y�-�w	d'��7k�H.��*�oM�E�L�[�C��-!g��8��:�u��{:��;xDj�C�sdB�\�FӬ��f�FB�Eܳ��m����˭N�ĽR*�-&aS�3%�Ҥ�!`�����I]rv�t�P�h�wW�O}��4�u����Su��8�|�z��8��1\eG�T�
���(�h�Ug{݊"�����5�t5�����VN�I�>̄,lԗ���<����oF���R����r�&:t7碴^�8d�2i�U)[�U�)�YZ�l��
�.�q���ݦ/���K
�������Em��D�:���x�wu۶���	�Rv��י�IC�ve��hA$y�t��7�y�	W�A���r4d��L]��D�-��9ëk�=�f康�??CݒG)�s����x�Y�6�ƚߞ�ѻ]\{��}ٛ�8�KSK��$���r��ʚ�ݍt�\�o^�_���+�7���שڍ�k��5I���#����Q@ԍ�\OӮ�j9��%2��T�hi��%�p�ڐ��d8�NF�}�[L^��c�Lw^{�֫��7(�J(�P2�m�SG��Lww/k�t�)�iN�v7e�[���۝F�uG�i��uڲ!RȦ��M*n���F�}i�c�[lF+�hR�6(�!�b��K���٫�u5���Z���l��~'O�ȩ-��AU���m�����]��˶�����Z%]�h�0�]�5�PA4�y<�O'���|u�U�m��Z:�ȡD��ű�|j1�*���S���qR�������|�J�g�+��Z-�Z]h������Z��桕�n0���f�cj�(��7%r�:y<�O'��1�L�E�h�ݳ�њ���&��*�n�K[Q-J7&Lԩ��:�U�m3]�ȹ�����V�ݳ��[Z���a�.�R֗jl��m�b��Z#lZR���\UQL��[����ʍ*4l����X�ӵ��R�*��)][��)QkcaF�l�����)KV׷n0��-���6�E�f�+��ŋj��1�*�Z9K�Q�T��JR���%����A-�#�W%klV�X�T�T^✖u(��֚)B˟�C�oha��·�Fu��(�V��iL�*�YZ�ح���W�s��%m��>=­[4���a�-�ֵ���|��^o8�s����nA�/��
�
&=����,H�S������'Fp#&v��9�����uqw��%m�T��f��O�!��fp��-��!��i��M��lԦ^J^�F���(/V�$�{�S�&�?�z%���_��7C���I�Řhaʫ�7^��һ���(����v�2z�����xoܽ����t����m��~1�t[�T����Q>#��L��b�ݽ̓u��u�q�Y=ӗGCf�7` ���?��7�*�MC��'��3�����;�9�2C�꫻�c�τw o[\��3-b����g�����t�0ǽ��l���H]j���z�<�^���{����>�i#gnX�=h:��{���z�J���.�����'��v��O���y�m{�U���ܲ��+0�9�����Ҟ8��F��0o�y���OB=�ux����U�D�
яp�a�U�~�&{�e;�+}�rŷ;qaKЕ�M�,�UO7�hze�M�w}��{(GAm�Xa{I�;�m�A����|"3-����Om��p����dX?@�5�!Ή��{5��S&��Ҵ�k8�<�����[;]�1�>��>� ѯ�ZAL	S��s絷�7g('�j��We��j�+�Uۤ\q��S��7��g��4�3]Y��ft�	v^�2͍'B��$��e�b+$ݚ��Q����o�T�~ʠ�[��k�S1%޶�8ߒɂcw1�wb�6}K6�!�{��W�]~�A+�/�{	txs�!�3ȘU̜��@Z������:mͫ�B��EU��<g{�{P~~l\��u�D��c=H�w������+��w�D���<��	�q��z��y�T$�#�]�}�"&�й�q3��,�8�C���5��s{x=w��is�ܚ<ɺ#}��pt���zi���jr�#���IS�o�b�w��Nc҂�U	�c�o��&�6�Vi�;ٰ��|}^s{�����ө۩`���������"]�5am��'>���1Q�xWyx��9l�����z��Nq�����`��fNо��M�Q9�~�>����Oϼr��P��/=��K�w�-u������~�Y"����6Q�DQ��(�.�"��I.ŉ���iB���]�7�Ī,��Ur��莻��F��O^�����P�ÿ��p{��$ɯ�y[/��'6�����yh�⟩8>3��b�'��>X5%�ٱ(V+��	5e�X�u�e�Ƶc��N�͝�{���`��j�ݝ����`V�@�<8��2s,I���|�3��'%�#/���/$3�v�~��wZ���F��^c�+�)�Xs��3�G��O�}�|\^�7c��S.�ʡ�0.�����������zu{>�7�ź��O�Ͻ���;L��>޿�ﺄ���S������"��'��}.��/	��o�k�2��� ���;��Y�6�U�~�u�n����������5�N��j�b�:�l��h�YP�S�j���<�О��sW�y�Q�A
f��n2�M�V����P?xx��ت�{���G���z�,Pߚ�VV��;6��o�LR�q����g{m��+N�]�g��W����̰�|E���4�81'U-��x��W�Te����ך$M3F�1�h���F{�£ߗ���G�?��o�w$w"ǵ0W�/���~[�n��$4�<�,�9�j�V��x��n{zb{I]�[絭�/K�N�E����*����!=�P���D:��;�)�m�{H\������u>s_3����E�!xN��SC�{�+��lO1����L�u�\��c�Ȕ�L&��U�)H8���������5Ҟ�=�n?��ܻ��|�u���{�S��^F�S��jk�}=+���w��NB��v}Fl��n�I�'j���9�>m�U���T����*���^�z?h�
��tǼW��8����X��ko�X+M��s�<�;ܫ�d�=���Iz'n8�c't�4f9�'w���ah��N_V��I׷*�*����v[��^�w���6��!��Asٴd8�W�;§�5=��Wo�Zw��=��q���ܴ�����\s�?{�f���OI��cϨ����Wb��O�'�	����{�sGI�ݧ�"u���7|Oe r��NV���WZ�'�Znιtk��M�{JpͯU���[�>x�ԑy��a��s&��������$�9�s���A����8�9N�i��Xl�uv�U㘰�c�_W";�wZ˓��f�k1�&�GN�/�D+R�J��k���im��~ա�/2����'&�����}��Kt���֙�p(��Ųn�	ޒ��^�0�������嫭2']��dEm6Q#"��")M=���t�U
\��M{�G��^�\��'��<<�t�}����������g��&_O�{�k`��{_���hs�K9y���Gپ.Gq��}�k>��@���=P��7��Sߟg)�P���KF���t��;�@�kg6��a;�W��������o��}�SDM�r^��<[a㏅�@̼��g�@�FiW��7O߼��>d���\ếG�r���D�h�'&p���@��br}B����/ޢrA&�6�0�|g�r*��T�q�/ф��^��}o�׻~o��y��Ǹ����-�>$Bˈz�{�gv��MC��~v������$.66����(w��#c�+�a�y�k�y�p�Co�i�T>�쿟'�~� X������؏��O`�_��$�����:�������Ͻ�k�餍�O�m�>�Gμ�P�b����Q�鶨��KfYp{mn{��>��}N)�:��	φ�
<��|n���ܢ��W������t����.����b�����i��\�^�8���I���#��`N��O.M}�9���O���;d�����g�w�=;�ZonVv����zN����瓯6����mz��
�]���]w�h�/H�OVKN<�`�d��'���OC����{���;����GY&OkW��ܮ|y�����8vm�c e�Wa0j߈%�#C��b*/rz�J�=�R)ƺ��W���;ڸ��c��մ���<�y�c�NO_w��hm=��푼���������߷����{�co���[�z�~u�*�~����+|��W�ћ�X[Y7$ڸ�R误�>���%���5�����~��][�UN��M�^�#Usa��yHYz(��	���FӋ|��W裞���%���J��-�����hN�o�-7�M��]��Å�/�3��xg����3��_o�e���R����]�j�{,_��)9/N�^�����gps���'�ݮr�7��R*}�g��Rd���[u�g�H/OӉ��y/K�{��t����ų6�и�,V���Ah������3%�)�v�f�*kj�:��RYEJj��mf�6�ܗf������x�w�+��N�x��e.�z@�K�Q5ՠbgɡ<�ˑ����~�9�zZ����1}U|;���U�M��k��+�J��>x���}�;߻������u�|�si��~�ep���Si3�9�'�y����/o�W�d�n��`�cR����.�����/�%E�7�߾�@��UV�y{���w�V?ӯ���I�OM�i[��y�4d�߫j]W|3����k������A���{{�Nlǹ��-S3��k;G�8�X0[g%<���[���O�;����~G=2{Q�tOA����ْ~���;_U�7{���Ǉ��A���{��n4N�����F��Y�Oǟ_�Ȗ;I�۟:��?p㘠7�ao�m:�{�س�"/�O�⇡CW��L�x�O(>r���A�H�x65Y��7�\�QՌ�����{�=���sj;��捃�/�L̈ms%�JZ��8�pj<͑s�n���A�;}��^n���E�5%g����E���0%�����4d�@��)�BZo�xr?D��k�6+���ё�B]���&�,��-�Ӑ��黀�R�E�kM��*��˼���7�l:�S��&e���V�/)��S5P.��7N��#�*��z(M��Q����g�(���>��I�4fU4��2�@e���]�~����f-��D�L�6��Xg/�	��ƚ�N������{�\�)�ۣ��5�7�yRu�i�y���߽��� �4r�'�}×�Ix�$��$�%��W�ߦ��f�X�z�:qId	oh!yܩP�@��e�rr�}p׆��b������o�X/o�~�n��w�3<�g�W���>��i�]�����'{�d�7YC�eR��$��*��u����}���g�=��5�Y��Α����[Ǻ�մ���s�y֯c��|��Ҧ/O$4��W�8�|=�ૂ��h���;��%2�|���z;�m�p��>/;�y�����ݖ�]ƨ䍞�S>U^5�o���nP�ه�hfԮ���� c:Sڍuu;��J^n�I���q:1BT���۷�lc���^�8�f��철��fG����-v�Wg�oU�F��c�}-��WDU��]
�I.�L�.Zd����/B�D��>v(L5��ם�5�g'�ڙ뼵�l���s�/�bg���v��W�c�z��޶F����7������񯯭u����_f��>��{��H�f���\�=�3ɏmx�{އն���O}oc��W��&�=��½i�Oܻ���I�>�gōUY5	Aq�Dۨ<���⤋����Ѩ��k�TV�S��l����+i�����䞹ͱ��=�~��siҙB��A��ܯ,��/6ߏt⒍�q���{�Q�Md<�|I���>n��F�gH|{2�<f�i��>B�L[6.��)z�Qc3|6�p�7��;��������7ç#�����WU�x�g��j �HJH/���w^�@,�+6sC���>�=d����:�����i�.�a�~}���A�%��DtD������7����mq�8�Vy�!�g��'A����2�wM-F�ݐ�G�m淠��P�`ٲ�E��A!��Z:�k����n�ԾF�-���dRK�����Z�|�Rudݼ�{�!�F�˛kЮ��Y�3��)T!�3�����=��Z�%C�jᤸ̙�BU�''�B���Hs-R7�@՛�if��^G*��uw�&�7�㍾��J�q������ʙ=g��
���*g�����돴�TgR�l��^V�����Hu.]�G�u����}[)Z�U=ZO3����
{W2{�M����{]�M$Mΰ��߷�#M���4S�zz����z���ގ���מs�ؼ���^~�w�Qwܞ�9�«���{�* �%Rb�z��&������e���;شU�}�E��]U��%���v�>�Gi.͠&22�U{�	�8�9�z�l�
kެ���E/ �8��ִ���/��;G2��1g�����ՙ�̰���l�>UO^�z�+�)ut��˭˧�~�fo�|�=�#Z9z����]�P�ts������url�W?�B�}PR�W��}^���C�I��5�S�؜����aR����G��}�3��q�O���Щa|�t�C&��{g$[_��3�m��9,@���5X��y�����7y��D�.]�cNG�N���{�7����k��w��t-Wώ&O8�I��y&&��Þ���-��\�4�:��]�8_t�{�<��n����%��35l</r�N��qq��p��ùg��V�̿�i�/�blg�t��;(�l����\(�y/M(��\Xd!e��\��i�JvcĸZ�u�!��-i�L�O��w�0�[m��R+�v��n�{�)ڎV��7|���0��9�S��f��S%���I�T���)Y�Yx'H�\�!5�����PD������o�=���k^�I)��eFm�Ϳ��Z\۔a�Hó��e��k����a���.��n'%r�>�z�e��l�wu��U��w�51���v���Ǉ�#Ie���byw�+G.�%wݔ���G%��t��W���]�Z�x"�ƭ����룗��S��'0,�J�t;J�)��K�U���}W�(�9ǻ�sh��'����Zeزv�]�ӥ������2��HP�� ���y�{�䦯p��r��0�ѝV�Ξ�I5"qvG�(Ñ@WY����
�~�&��/i����v+��|qUn��p�4Ȝ*������Ϻ�o�
;�Ծh�6�Y�����w���/�
o ^���oq�t1b�\�i�̥H�S�K,ګ�PoY����M��DA��H�Z|�_���^l8���~��'��[�i�^�vsB��K\�
!��|5-�Z2�Ӫo2@�̟��=�3���zIV��^�"�OF���P��Kwr�ǎ}D�c5�i�TvP�2vыsl�衂�}�E�7��]L�0���0�8�IPk}֓��&��j�g/7���A��H���u6-mv��V�.-����U���-��e	]w��rο�*�D�T��'p��Ӫ�"��1���c@����@��x��d������w�gX�`y��L������M,�M��Y�������m��W6�
��<��.l1wN��0���C��z��
vH��W�.���Б�჏���J^�g��osF�Z����ޅ"�f�[���#�r���S-ɼ�����U��ùo�5.��uoi;�q�33\�}�y�A��0<��g6=2�w��K���Hɞ�r�ܩ��ʌM�{[,�VF�����t��伡g!aJ�����B<���=X�)�qg_��լ��|kV�x5���DQ\Za��h3&��iL���Ǵ7�M�-0 ��}�v�[�}aml���t�6�1˾.��zv�ə�
�z����s�6�p�MWR%�h��K��<Ysa�g���ܵ|(�C�e1&Bm���_P���z�Ӗa�;�]�S"�M<�b~�q�/�,�4�R�Q�ʾ�w]�jW��:ҋq�:��-kM��q��j\m��h�������:�S��>Og����������L֨}�Y��{^���_�ϟ6M��(�ȯm[��(�P�|i�2g��단���'�u/j+-�C���}O'��k|��ѣX�B��|�9w�b��Lm�Ui���<�	D�����K+�9�B�W��luׯχϜA������y<��C��f�1��_.���n�!��y45��ߔ�t;�����k�j��NZ֜k6;v�iu��~+���>b��t�<�O����f�~3�R�|�w��aͽ6o��y�;��|o=>g��pd���M_��+��/[���f�w׾!yz|�p�Dq��d�L|�Lֽ��^M������7\�o|�┭�PAEM%(�N�K!$�~l�>Zj�i9ɘ��o�n�Y��'j�j���+P̺�m��v�s�1ek��2�b�-��l����󮵶��f�v�:����WQbv�7q�6�e
5�=�Y\��xB��3Q��W	X���ͨZ+m+my�䦵��j	e�4�A�\Ҵ�nlVҖ�ZT��ǚ��*k�Y����b�)nM��l�����L�����.i���Lܴ���j�v+��S��f���(�!"�t�$^�W�F(I���I���y�1=�^��S-��!�s�V�,���.K�o�7��-����_�{-<E睦ܳ�Α��F�>J����CE?]x�|�(�[G:�f��k�P&v'(��ޝ�<��h�j���f�=�a�}�v���ǁm�q0ISiù�t�m�@��Zp,v�]����%�����֦g >�<X}x2~㙒6��4�
�kܥ��1�K@�؞^���_�|���q�.�EkK8��|1Fq���	��]���D�o��x�����9I=T��vQ�1����ٵ�[o@od ��M�į�Y�/}��D]	^}sS~n�N�a�)b��<le�l��U��0�&�]4ɻɖ�+(�ߗ@5&l��<J��}s��o�#m����ϰ�/�����>���_�tS�U��:��QI��M��1��|`76����b���H�p�xY�}�ʝ嗧�]��841��ڠ�~�K_�NN{U�7N�O-X�|�?��+����~_�'��������������^Me�*)�R}�	P%����8V7�~�9����r���#Lx_SDc�^��K����xd�+�]�9L��eH^�嫄�����k3*�q49�X#�刱���3����@��K�%���#�3�}@Hbr{�����r���՟���iЙpv^�����a�X���k�<AK�x�0�x"���=�"��KX���She=gz��b���m5�d%'��y�M�5�9�1q��ÖP4&;�3�`%��4%��K�~7R'��T�b�5� �m�[L�l��j�o�*�'��?� OO7����Į��1������@P�:�Y��{l3��U�Y=���dV��F�]yfϮk����50��������M����奅p���Ga��0��)q����]�@���q�2-�]�k�U�5\�Ňr�]�sHM��t�u����]�r����9#?.���u��H�b`�X��mހ�<�Pfˍq�
fو��Z��wyW�����^O.�h&���#�S�����NA۵�~���.���L��j��r���y�Lt��4�P�Y��K~����=?��5���r|�SG�s"m�n�DRۙ���m��ݓ}f� ��`���3IWNμ�/���8��
����~�Mbu[�u�Y����m*&H�dͽy���-�kN�l�,hj�wyFm�z���z�?�O�{b��m�d2��7]�۫9EL^��y*m�nk� ��f(��YB���	l� ;�f�åED�¥g߿�3K�5���0�{`��Q���쉘9��k�*��x��s~מ�����ѓd�X��%Qm!f�3���׳�jx�'�|�������*8�\gΪ�֯<_`ï�*��꯷=�L�m���|��@	��_m�'e�w������7h#�_��r�W2e}�����+ͭ�閳31�O)��,�{c�n���͘��07�����z���{T08��h��{z�q�K��-�2�\�c'����} >\���9=;w/�2�{{)�vi]�(k��|}w��0���
�Ǒ.C.�5s�m��>cv�	⒆�
3��s}����y�S~�$���P�1[�����&���|~�B/ܫ�)��6k(s4����w�u���PJ�0>yEJe��6w���?3�����Ѐ��t/�Xgux�׆���w9�_,n�Y�j����VsȪ8h��1�U��`�%��9�a8���X��;0�g�\�`s��x�l�ǲ6�0��s��3	9��`��b�J\m�l���~��),'؅����9�>[����q���8�@�ޏ:�`�Cr{S���S�$���%&.?5L�z��.�Նy]>c�Zۋ�xO �)�3{Z���郆֮�.i�J������:CP�3���v��m�ה�>����Дz�y�w����@��&��d����aY����}�:��ʐ�������g��Y��p�c�򤪯	���\1jt���\�PلT�3�N�aF�f�����dt٩��c%�m�~�(��c��Y��5��upt*��1�V�nu�Ѵ33�?1��tZn��6����&bꔫ+Qx�dNЭ&ß��᠃XK�IΣ��@�g��u#K9al�G��7L3�AD�� {a��y��Nۆ��q!\d�a����u%Ю����C`�n���0U�P�TS�f���KW�3�	������Y�h�.��R����\�z��&�Y����ݪhj�X��B��BD�j�w�y�;�fNw5^�liD�t혞%�C>���# �ץ�57�T�7P�*����$TM%t+�p�G�Ͳ�ff�oF:�u�{[�g���"jr�����3�����QW�?�&<ZF��Ʊ��,�ųф����=�=���n��������2�E�%�*k1O�Q�����<�g�K���;���7VҪ�'X+`��פ̲��Q��ՋkX.{^ɟ�l=�S�4{M˶P��L��lv��~`�f�+���a���ޘΞ�^�j�0��Sw`	U�բ=M��b��,)�|��x�ym�S�������Н� ��eY ���`�;�ڇ�JJ{���.~m�T�~`-T��Ա~�[�z��9il�"�g�Κ��m~��e>�T7�ð���Ur{
 ��#�Q#��w*��Tnʕ}���͐��ؿ
ܫ�]���x�d�]z�yĶ�fҋ��e]ު�WsU(w�\(¾"x`�7h���n�R�`��y)�]�,����ѿwEK^�S/w��ft����Z��ݖ�-P��>���ޤ\��U�s�=3}��e�l`O��n��C:��/�DD&޹T�Y����5),��;�i�:� �Gj�8?]�i�!Bi�.Q��	މ�?�=�!��-���e�67\�v��1����7�b��܅Q��bSN(�43m�����ݸ�� ��3�`�axf���Y
I��k^W[�f2�ϡ��V�<��Ǻ���;�&+��3�n���͝�PX"NC-�R�X;Vo/���S�ʇ���i��dckWD_;�=CE�Y/E�3��CCG^�˔���.�Q88�����fN���󡈐2�ٶ	���\GO����D�T�p�"�Ss��ٚ���4�������8g��9
��0Ni=	��󜼟s@������m�T��謾x���y�_�3^���FS�wE�V��K���`K��?����{��uи�a��Mz�ꎨz�hoQgh��e�q'z�s�9%�^�J���n�N��������`���3��&�����9r&��-���*�������j�����d��Q,�l�����ֻ���xi�DO��xZFԤgM�9���إ��~�:<+�˚�0�P��/B�ϕy��4:���U�ʌvo�ol~���o@=4����}{U�!�:M�T" F���M{�z������Ko�+��Y�*^�/K_m�{Dd��Թ�w����l�[4n7��J�4mn_RJ_M��p��_4��`��y���_�>/�utĜ~��͉�,R)����=�SN�Y�R����|��}5&�oط��0�;�T�m����T�qo�h��E�'5P��-V0�}֧���-���E��-�5��}���F=�^g0�Ś=.��j9�/g�۹),�'QH�/��cN]<���xD퓂sP���A��S"{��}E�C���E�x�I��y��K��t�4�e�S�nN�ڸ���Z�7�nLce�e�b`s�Xc2�C?k�hOƅH�th�`ъ��A�����NGK���4����[�ďE��P�$��ނ�ψ_.�}i|�}�����=R�0��Ր�qe�*EQ*�L6���>�Y���&h��lg���1�޹3�Y����Ї��3h�Υl�'a�яI�t��\Χ�Գ��6���r^�9w�z�ѥ�8�������1�v^s��BW���]_�=����#��w�	��c�C���TC)���{��T%��^]����lXs�}2��6���5��ݯO���0�E%�(#ȫE���̞ay�YuO�B���(pv
9�P|�O��ݥ�������xz�s{��
��-�S��:����v�l���O�2����u�@Ṗ9 �R�ے��ӧ$��c')��+�����=[��ׄ���L�b�7��꯽ت�̩����b��)DQ!�a.L�cK���t����U�r�o���,������73��c�??><Dw߹oT7��߲7�Ȗ''`�v^�;���:fǞB �⮝�Q�wM���y�Ezu�φE�AO�6�L�b���jSe8噵M�j��(z�P�mR%�T[����P��cQ��/���	E�up���^���uop����X�9�A�<Ҋ�6��*��1d�=���jl�X��5�m]��.�Bl�}��?D��<�&5��bScX�Ƚ�O׋+��5�XxR%��0��1�����Zިa"����z���}Z�%�g�{`.�C�����*�i����f�v�۶���>��%`��b]L���󷃩]Y�ߴ!գ��VH!��l�6����R�n�V�,��e'A<���JG�E#�4�]�g?6Z�����ɟ����������Yb39chY7�Л2F�-l�a1O~QR���<sm�cy��s�g�b���1���gg����՝��l�^Ǟy�e�v8ɇ�7Ju��,��p��ax�,�lw�E|/��.�*meڼ����*o�-�AJ�lNo �̀��e?U�g{XIV&Nd��v�<ԅ�.�|����f���\��i�)~���o�g�	{}��4����֍�����-��g7���W4oeλ��˱�f���,e�*
��tF-i��	������np/��N��|#���_[ ���2��y�
Y6�9����_%%����[�X ka���d�^ݴ->9f|�����49�������S)쮲ްN�iOFGB1<�K�wr���F�悀�Tɨ�[:z=̍�$���LM�H5g�����r��vT�;N����[��W��ַ��W���x�^��~�	�(�����G;8^�.����ǚ�v�88�ڙ�l@o*֮�����0��ށ�ږU� 椥�v�-�P����?-�Ͼn����k�2gᢽ����$�Y��~�Clq0���t���mx��������+	3o�������!֨騳q~�Ʈ�7jY�o`�������$J��K���{�~8�jUy	�rS?N��=v��_�}��Xf��2<b�R���lk�"SEZ��M	�jep(uM����V3_�%�}�"��S���|iw��|��ڄ8�g�
X���{����tڷ)�n������~�̜�ڞ����3Lz�����
̱vݧ���u��v���L8��Pou)��+��ʗ7��~c͍^+�ـ)�D5eu��X�}��*-�6��ZPx>����1e{�RӞ{� �0ne�=��M!)	Yx��^�f�yT`��o�o'���ב����fmu.�d�u�E!vo(D=h�nU�.��u�j���֔���������=�8jep�ÓJ�P��Ė�d���UL����X��'JQ}+א�⃯F��Y.ۍ��7bS��h����n�A��[�h��Di��x#���7U�bw�i�iOc���q��\M���a����5�[{�z��?=M/�q߰>.�4"��\[�TS�[�ő,�?6�Rq���&�3%.�.s�����C?��#_Z��6�VD���W��v�Q*�=�K�͵[:^b�H�Ѹ��3zo��@|7�L0�<��0h �j���m�����[_��R�G_>���_6�>����E�J�����.�C��]�(~}������N���w��4��+���ٸ��ݐm��ԓ���d��������D=����]�a�m�6���S��n,�T�ӎ�ҋ
݆gm��[>���ړ5�Գ�j���'z��(��	�Ǿ��]��t�`�=o@�$�z�;c��w+��b8��=CEA�/A�Pga%
�].���M�,n�Nݬ�֙G44�9%�\aQ^�f�۴�� ����x���f{�_g@���Y|����~K������x���Y��p���m�Ƚ~�����l]]��Zt�P �<�V��e��+��ڳ^n�c�4��HXt�,ʒ�����L����Y/�&��ٌ��+{�>ck��(Vn�Kd���U_��H1��1��{�������w�?^�^�	���*TKL&r�����=�;��#˾��n��2爼����,%�Y8�����Y�i��@&���=;꧁:�%�.zQ����VwkҧӖ�^����q��:e���fש�ˍ�Q�_��j �v��=�h�d�k�V^ã�7hV�9Tz�1�:`d�l�c�:���Z�U6�[Z�at�L�@��~J�c1�!/VߘϾ���]ԅ!莧v�Z��A�އtRt�5��\Cf�7�veV�����S;���,^�#i�)k��zh·l���U�����7A�\����U�Y#��Ǡ���A��c{3V��@�����˯3�0�E�� �'�~fʾ�gj�J�X�q�1GdM�]xsK��ں���[.uK���,�nqԶ�5o@{v��/^��nkgd�+�]��RP�4�;ww?b��r\�������K��過��XcK��j^;�����nʶ�J�Ք�
��z�H����4��P�ׂ]=���{��u�^}�sm~�������Hi�O���ߘ���O�p����ּOu�{��;��r��j�ʂ��C>1˂�o���������s�C�$����.X��cEs��9����A<x �<룂%n+�;ƙɸ��̨ua]H�Fq�2n�9nLJ�.���e/%&��b]8�Ʈfd�zpE5쪘�d��7���K�?l:��o�ḯ����`W5�0q+NK���L�����aG㧢[�idډ��e�z�=.��u���K(�n��&�]��?/3�\�s��zȖ����W��l]�|�;ǎ� cSN��Jկ��h{���(�ZݥW�7�P��nސ�P�zx<TY�Ӓ)�l��~y�8m�������4�Єn���G2W_i�M�����m�-�L���:XR=1�$��k�;��(:�Tَ�)��ueǌ�����wv�Ge�1�5������ڹ-�)}� ªo�޷��0]�u7X�0�\�� ����	�rU2�n���|U/oLs\�O��e�<�>�x�G����y���fn8��q�%��䝗������OGOG���n���猼T7J�j��nJ��랮|�o(�-��<�P�Gl��j��A1��>�l
k�e��/�M�4�/E��2�M�s�VN�qv[x(0�33c}Yϖ�)�K�Xj��\)�֨ͭO�"��y��xnS��ޑgNZ���̾N��!���,ރG�q�{Ý��h�%!Y�����S~sܞ�w;R�w���`���>秩���O�
X�,��9�`�mV��".bQo:_#���9H�����(���n!�\�mՂ'�q ��}s�|`%M�W�B�}t7��9F��W&Z��W3�h�9LFo�=u��.��0]�8��fѤt	�����F��UtSUb������y-ǒ�b1�֏j�VB�V�fՂYE�[k9���8p�|����L�����O������'%�=n}�s�YV�84�P��Pr�sβ�1�M؜{I�����d�kR�Er�^���No��"|�c����y-1�)�����q��̾y'O<��\���.�����=�=,�iO.��C��ǏK�P�ח]Y<1X���}�d���.;)�[�Q�ClL��I���.���*E9�N��0� ��X������<�#أ�;]!o�E��.\�����6Y`gh��<��ϔ˷6��NU�ҥ���:H�eot�f��oOB�Ry)��K�ql7Cj�Fn�{��~�����g�>q�ǆ��P	8�'��P
wKf� ���7mY�[� ������]aL>�C�O܂�r&�|��R�6�Cq�)�D-;c��v!L��K`W��Fs�w��4f�`T���ݔ�cL�h�3�ee�)/��>UL�r�tsg8�{�<��µ"J�l-9j�k�K��d_uLV���S����d�~y"nU��l�^Y]k�*0EYF[UJ���eTLU)Sm�-�����嗑����#MMX][�O���<�KT��%�(��KJ��mT�h�&G-��k4�1j��U���V�[e��3���\����y<��ꭱ���r�>J�Fִ�%ԩAR�Zڶ��kh�Z+~ZkU�cm���1���\YF�O����y<�Rڣj1kjڪT��WR�Z�h�X���E
��̭��n��Vh�*%Z�m�jTkmӧ������ݢ�dfK���Z�a�ͫQ�����AAb)啜����SYaG4]B�q��{+T5Z�|�
�iF��m+F�|����Es,^L������Cb�l(���hrn��[nr��PQKnkR��kX�L-KN���-��V�EL�h[m�J�iYjTjҌh��T��[mQ�(�J� �Z����ky���:�sT��T�ؖ�J�ɦLʈ���sdj�����j�m�%e-{h�Uk"[+DQ�Q�0mmU,Z�T�B��������{�}��i�绲D�)/�D!%�AG�bzW��މ�n�r�>c3\/�R�ܶ-푇��"�%�'\�@&�K7w�(u��GΜ��΁�΀� �Aq�ѐ�5���;wX�{f%��y�oq��T��'�2A� � �	��rB�K�o���a:b�#P�a�4%T�я���S�<��ƅ�%Ra�c��l�,��ma�����_���3&*���0+c�#�ы��Ly�5K�1X��}�ƇX.gS��$hcW�t��j�͝��&�[�O٫�M��3��0me�fx�P�ݣ��X�G��j��Fmכ��M��q�|c0Rs}��Kj	|Ťyy֠q~��--,�Q�`z�Ht�VK_������R*X���5J��C+�ٞݵ��Y�����/%r���/���t�}��Z6>zCv���\�f�S@�Ȳ�ed?@^�\�5����3c��c4�t��ۺ��6��yח�"�8)�e�虛�l]��ᤸ��pSΊ������_�)A��`Cf��w��n��]��b���Q�g��!Dti��n^�Ԋ��JK�|1L$ꕯ~΄CнSe�<�D�r�aM�+��3�%�u�{�/D���_�������xp��%����%ީAN�,��驯�.{�(���j��k�h��0���p�m!6�U���}�ȗ��+?���)gf�~��@b�X��46N�5��p�a9���F�{��ر���i��lq��\k����=Q��n���a�{�����,��^Jfyi&K�d\j����x�}?y2�v2i�ܵ�&�}/�{ĸ�w{�X�B�oNxiU0e.�;�%�훻��;}}�~{��ﾯc��_��߾���C��� � �o0��͵}�0��j���%>D�+�j�F�;[X��)��aR��.B~��C0�L�p<ӂq�DK�:��bݛ�����[(�\��J}�H印js!���.�)�(�~�7��o�h|ꫳ~{+u8m�^��y����;&f�)�`�T[�B�
���y�)���@��e;�hS������zܩsé<�ϳ�=��O8�r�s,���P�ϭ�����X�	��wV�vtĳG�E��1�&:*=�����*����������6�90�c�%�>��f����|.-U�QzƆWI��V$z�Llmת�?Aoh;���^�l=3�S �;<5V�"cZ.���Z��g/^.����mv�ƺ`ᵛ��2�9FX�M�l�F�sSf����1s|��=6�>���[=S��g���ѷ�FDHvp�x6Mwd�A�C�F&w,�>2�;��n��?W��%��̀}����2���s�j�7�t\7ЖΫ���Wu�a^i���/�O����̋i��ߞ��������~Fm�>�"���6�ne�ֲ��k>�����U2yp�cZ���_V���{��o0�P�fc�d��jv̝ټ�6Z��Y�qt�NM��X�H.���R:f`��ݠ��x��p�=��ǋy���U�ݪ�k�2]H���o�~��q�}W�ף�>���O�I ā����   ^"��Vb
5>�}�l	���%��YȌ{n̈kj���o���o�M�OH�J�Rl|P�LoB���ﮑ�9♰~���TC�A��Y ��Bm����,�9՚Ż�#/�xg]
�}��j�l��k�E���;��f��saꃻ��~���<NTlws�'�: �d�ıʽ���~Kv��n�jk��9�Tlƻ�X�Ň���~���w3f�^k,At�Ge�<]^������6�B�V0N���c�Z��}m��웴I�<�H���ۈ�Ⱦ6��}�Dj��a�$�a`޺LJ�V�FA��56����7�=���Y'[Pv�"�| �v֡(An�d�,�=Ƒp�T��΢��X]�DHjvv��T��x^��̼�vy��V�<a���H.��}q,��x�1"%W'{���%�x1���&�R��(��C|�����o�����F�;������6���}!�ґ�wx��E��
W����d(-8�˶׺6�cAap������;h?��e~��yfT�˩�R�/���g��lܩ��ٱL3�*%2V�B�=�fԒ�ڲ�&J�&���#g}6s��W"����\ȫ�;nPݱ	%`pےv7����U��xS�C�{_���񓟇&y����ɕ�,������$�$b 
I}~�����)�����4�䨷`]%��,�a�K?*V'��_��">�2FƓ�a"�q�9f��ș��Z5�Qn��'���z���i�}3�0{�~�+܂��?{�)i$;k��e�<E$�����r�WdH���fc,Sl&��n�$�����W��%̌nk�w=���ϔ�xD����wH�\��1˙ٰM�� ��n�P�{�;h�9N�|�i���*���ν�E��8z�@:z�ZIG(|��O��U)��X?qc3*��si��F��E���Q]�i�2Ci5�v����:���zw�C�Es����Z{��3�	��~��2zb��/۬t=�h���������2x�%)�=%sQ��մ�%t[�kK��v�|r�]auf�Y�����i�S���΄6/L�"��S��:d���M��۶�l�Uyl�4��7(�ՑV��fZ�Ǚ�G��5O���"']�ӄ�3�49���tRuϩ�?�E6�Js��ٵN!��.��3�T��t���h��E;�W�)v��GS�a�I���4���bGU��yv��&������M3��/���0�1����{��K�/Vf�v�/��V�j~W+�s�y�β��(���*�eڕͻ����?� i�N:����I��;�u��X͛]+�����ZcA�qk�l%H��R�c��C:8�+f5�b��<�;�������o~�������@�G��{���� ����0]Z�u�:-��[�&��!Q�2X���>�#ƿw�*���@�"�~�������&����ڕ�<-�;��K���\-�	�):�&�/id��YB@=��#��/�L�T�����5_�-��8���={�����"nIu�O��c�5��t<�qc�@�h���Wrb�
�
���������蝳p�R'�wh��m�z9r�S�H�e���-�|���D;mDhbp�;���s��mi���\�>U�[ا�y<h]�UrqغKF=,��]]z��l|⸏���5�׸��f���߃tK�~|T>~?Gg��U�t�P��3H���2)�+�
y��Y��\��4=�π�O���@Wʇ"'+y&l0[$:�42���CP�9�8���wU	���^��y��܉���q�S�6���"�yv��� ����"��|��LVC6K���b���"�G&D�s�c���s��x�w��Z|�+���)�*�o�15E�����}3މ��!�V������a��C{Ve�W����*6=��>*��ъwY�>gQ kӼ�t����]����M�޹4m�궞�2E��G�q���
B��H���w;�5��kFz;���y�a���xK�P���]eN�l�����U�]�K킹�yl��T1��}p�&�=��jS#J���9��i�rXI�W������HA�I�ߟ�~|�???����57�R��-�]��1L���peS���5�wp3n���3���7_�Өr�{��(�ل���ca3���>�I�a+T�{�(2��QZ�~K(V�.����Rf�iȘӒ4�.aL7خe���g�����<��r�2c[��%67s�\����u`V]d۽��٨f,�),�{h�닽[P�E�;jg���M�5ä[n�8��e͸a,FiS-O˯6��wR,�K�	O�7���д��c�Q��z��禀��%&�ǟ1�w0���X��Ͷ�<���¿ ))���T$�,��BS�R9cl�|�nk�)Y���z+�OW�[�罢�{{:��um\�]���)�ɐ�;&	�LS⊔���6qR��1�������m�1��Q��>ڋt �����^p���G=�'�Tpї㖯��0��%�g�Ui'���Ӆ�:-�f2�U�l{d];;!����#z�Ԍ�^��@��
�J�.4�L'�����Dx[M��V��9�5.-x)��y��^��7c8�A��32}�&cS�)��-�<m�a�����RG��l����������z���VK�32���6�x�;1��|��#9�3*�n7�Gܒ;��χ����.��F?�<�e�G� 1�xiz�����.ɵ��K{^���^;,�O+���2<K�g/0Tw���g�����~������` �BG�=�y���f��h��&�n͡�#*2?4V�5M���_}`�=/���@���@�=y�E������{�����gVV�vq� L��Msl�	3%�����s����~�Gަ�y����ؾi�K��s���Dqi³�s�M{���~�^�����i	]�Գ��}s ��������8˪rfQl�_��~{�%d�)�꣣+ogy.X�m� TSId�!�Fen��F��7�)c>�S��-�0�|*	�����ۻTY�^>k�����pϯx��FbT{o4!T��wz��_L;ag���=6��6�%�5O�f��1+��xL*%�[!�L��b:o̭��*J�V=�Zg�T>ܤ��,$ٳk��k�C�_�{��U899�:Vn�OM�C!�Mc_���sx��u�om��av�<<�|�H]��^�T���Qj/����ã-��w�{W#Fay���Gt�e��S"�5M�W�ec�� e�E'>t^�j8�]���ˆ�k5܄�Ly�l���I�nx.�"�Sw`��G��-I���X}>Br��U?v�^�2��H�UC	m��l]rc�����AN�q)�=� ��z�ҏ=9��@�'7�%��]L�G(���ݕ#�8��{ۋ���G��~=�G��^����?fS_�eu�,oet�h]��D�|���������H~��A�!�� ���ݜ�YRKz�v.j��8���l���[D���Y5����mC�4����;��G�2�u���z���{����`�@���?ށ���Bs:��D���Wa\KȌ�i�32�3;|'>%��˫��>�?G���z�B%/�oM��I&5���=B'�O���ލ��q�&�';���6�ۦ!���������q�>��	މ�����qr�鷁���m\D���^��;����i�7��y>��z�u�j]3���2#��D
>��?O�X�L�k�&˷U%l��4jb��,�P�\��ys�+ >�s�3d�z|	�g~j1����~�	�V���8�xs�lx���u�	
0�3c��T:����azu;�H���pGq�:&L���ێ.F��t<�(3�?}�2�@d�>����Ά"s�[^lн�<�\Z�?�{�!M��^�!|�)���������(���˿5�vv~+<����>4%<>�������+m��w�b��-��Pw��(�!��K0�7�a����T�}\ধ�Qv��&[>�
�ʻXG�+��g���6�㫒	c�n��n��NEt��y~۞�=�}����؋��n��{�q�x_V�1��)�|�lR������q��}����g,ɹ˥*�ʄ��,6��T����?8���o�����k�ϯ���������}��}����F$ b���  N,vm�h"E�+y���+o�E2Qί�l�2Y�s��^��(�L����6Xմ��<E�zw����r����T����@���@H�ݾ��U�\�>�0C&�V=4ɷڦ����tc�3��	�$��3��p��'{k��i�.�E�j[ ����}�I�|����n�
��0�]�Xvޙ����7T��q��mRT�mdph����5D)<���&��
�E��Se�k�քt��0'�ս���0�cՌ��䦟O��'�>�O3_G3����l��\�ť�H^�Z,��	��6��B�y���6ࣴ!�k��:��sԹ�	S8��G����_����ٗk�`7�:,��1��n�9@ؘ��Ϭ1�ζA8��E���/�;9wB��	y�ݺ�<�;�j�L�ʄҝ.�c���!��׶1��A/ �X�2�b��]ܫ{�a/p?,tD���O/�[J�.�	 �V�v�mOK6}@��m������]m^j���䃵�������ϙ�r�.;P��zx���s8�g$hc�ؚ-Ŝ�!)�6"�����"�$�u���Vm;>ZYe�ˈf���5IJh�ʾu4���omuj���ƶj.��ԟ�{��l^v����*B=�s��n����ˠ<����<�&\��׼j9ٵ"ĩ�L��b=����� ?Q	�� @c$�<i'�UۨFA������0nffk��������d���場Q�-�0�s�-����^Q�xV�D�0���S�ǃ��?��d_��������ؾz���LSZ|�*ZV�O!�8fӞ��3c_uϗv*f���0�a�+����Q-���zη�j��H�j��ې��À[1�����v��Dq��6<�"1U.�hͻ���j�5��oed�K�������+���EX���ڗy��a�!��k�j�wy�k��l�ded�U�s���� j(Dz�7^��p2�:��\S�T���eiEs�'���1�ڣl����oD ҆L�a�3�Pu4~���W�~<�R��߁[���������W�u1�aտ�xgO��Z!7����=�
�Տ�9t���y�f�e�������1A�Q��:m!1�A�K�e?��]�&��!Ij�Oα)�'c���Y����t��P���߿��!�*Z1��\[)��}x�.���@}!�v̮{x��7��Sr�{:��z�2#a��|(xGg�ct�	�X��ݻ��,�ctC-��M��J�yq,'��
YQ��u #8���M����,�j�v
�v�u�Nv��U��3	�s�vu/�
��L�ԟ���Me��+BӽW�ᶌ+&(�XD�+n���)J�&M;)�]/���t��)��qج�5��	�y�A(x����ᑝR�}�z�8�o�+p��K��1w����\��!ƙ9��G�s��ۼX�����\��I�`-�ı�pP�}9�蚭s=8pHPL�v�Jn���s34�E	�S�I�&Z����F�س����ζ��W�'b%��U��:���{d���b��Vj#$��S)�B��]r�-�]&�Z�\�&�.�"��̲�}*�������y���xy���njwG�GnQ�j.7��*�e+�f���fuoc��x2���3j`6f����l��C�D��ꍣ݇^:���;jcڦy�<���n���Ĥݩ��M��ڋ+��N{堣��[��8v5M���7���r� F�P�����Y��Z�uXV� NR�ӏc�Y�$/RGB�Dc��Y��.�7V��GC-��di��X쏆��!�Ug�㾏�~����{�X��Fެ����&F/	7�%++&]�	P���[���y���zk������q��v���ĕEP"�%���f1�4�;�F{N�I�ZDf���F��T�� &u�u�ۅI�kr���T�[�"#��ه.�+%��<A��B�GKcr7�d�ߟ���2��g.��o������R<"*if��ý�1)��Ʈq�-��5�C5�}[�A�+:���%�T���M�>Um�s}��e,?&�"h*�ʻ/t\۴E�)C��sB������u���\K�)u��� @����?]>7��w��^eg{���������ou�����>j0a#o�X��>��}Ci�Eg,�"x��5|�U3dS�}�v;i�t��x�Ё& 6�C�Wu&+�t3�,]��[�g��G�9wq���7b90�ѐ4��Ja�����ݛԟ!�����&i���k�()�.keBl/�{�����x�!����I���o����s8>��?�>r"2�O3���F�k.SV/s��J���jA*s�d���ϧeK��E`6+$G2���N4�>,�伆[2=��"{7����ؐF��{'��(�p�U�NV%�n����X2����_1�tQF�!�T��D�F�Bf�W��y���8$~��+��x�=|xx=������#|�{%�T���;�T��.�֠�M̢�Ev����q���z㙨c���g�������	���/��n�֡�z��0VP�q4L�w��r�+9C������!ϫ;���H
�mF�L~h�?[j�akN���7H����u-Եh�ZYKh湵���|����<�L��j��(�
�6��Z�֔m-aXTj1�T�X��eMo�أk:t�|�O'��e�e|�ȱT�e��J(ʥ�*�J%6Ѫ%�Z�j�2�B[E�:y:y<�Ug>&-�SĨ���[�t�n�V
s�Ί�jņ+t�Ν<�<�O֥-�2
(V6�VZ�b�%�yNUC�5(�m-���-��mKmcv�DX�E�%aZ������z̊��ͦqV�TȵR��ȦV
��K�֯9r�+[j5��S]�ڭ-(�iKVڶ�-֚R�PԱtkYR��eKh=Cj4�
��kQ+ljZX*;a�6�֖�z�ԤTR�E�m�F�Z�J���Cj+�TB�r]kF���F��	����Ҳ�Q�ֲ/4N"[W�p�Ѷ��Y�u�[3TL�ǚ&����Z��kZҵ��}Euz�X�=;qT�`��C���I��x�,�V�=C /9G�d�,0����XÑ�-�k��X��?W�>�{�w�~���@�F�@��$�I$P�)I�_^�~������������6��y/"ɐ�ن�3	�{
*S.�tO6�R���D;�����ɴ�oU���z��&U�x-�0qzǞy��U|4iŚS�
��ө#ܙ��r:�~�9��9�~7I�� �U݈�~z��w綑39���gd�R�mwG1�Z�Ops�v�9�QN�0S�����3Mr �Oɍ� ��yT�~^��ʹM���+���ݶbƃ<�Ü8�t�eM�
��/v�5��9��MSk�W��� ���p�0���#�lPִЧ7�5.�Kf�YQ�\��_��z��U=߮�mJW0N�"u0�͆*�&ND���!xM8��x�_XXkc��U���������́+��楝҆�p͚�p�J楒��:�)9\���c?g��%yfM�X��H1���;�K�=��I�D�F�s�2�au��7����K+�j�n����!���O��IaA\�l��ol���`�D
n0-S�r�U��ϻj�jU"r����7H���G=IÀ��Ed~,�/�IG�?V����a����rӶu��}O�!���%�m����V�%	(�=��t���uֲK��A\�����D�\���*��%!����rIs�7P�۹��k����������g2������-���Ĺ�q���Gf���Q��_������	�Ą{������������[�ǈ��iHM�H�z���"�[���ʒ�-�l���f�J���Y��X���Ǡ��"Y��6�E5�)d�c�.�U��*�`[���o�랃�c�H��t�M&a��pr����/ʘ
e�������#�K��8%Tȹ�Sm�k+$�q	����z<{Z"m_2ӛ���3� ��:c��gd;�BaF_y�aX�Sw`J����1�~�Ufj�-]퓗���U8�^�� 4E��2�S�v8M�ɐ��io5�������D˽���6{t̽2K�1��k�W祐$�U��z��K�uv�����֫:CI�up�-�mi���B�I�D���Z�ۚ���}��e�zW�{q�I������h+��~�1;��v��r�[_jU-K l(I�<���Bi��@��1���td��1�M���.�u�^S�VTSsW�L�U�*)��9Aeyڤ��bEñ�������)�X���G2y�,���	v����zO�05�tt�}Ƕ߁Α'�B3���ê�c;����\�W-�wN�÷N<���_lK~^ɹő�N�˧����p+��[7��c������I�O�5�X:]ތ6����;�`=NJs���>�8>!���z2��%jَ{��T�6�w�g��c�����)���<����}_��׿_[ޟ�$�a$c	���>����=�~{���r��Bh2d=(�Y�K��#�ѲL1��}�`W�(���w�{�P ���>1]��Ў0V>�6�����u�~Z�D�9ԙ8ϟ�0O�x�C
��v��"�Vm�ɂj�@�j��Ei=�wT������ǁͨY�$����?]/�r�i�3��&_��.����ߥ���"n�Mv��S 1L�W�7Y�7,f�Qa�yK0-��-��O~�}T�'T���)�s�K'%/���������})������3C�j>QRY��+�ǿ[��:�j�?.��vg��o�r�2�f���:�
��8�sR:��f�>t4�J%�e��m�����lfC�D<�&��x8����V��p�b]���B�v��d&U� ɜ��|�<�E�R~����̐h�����}7�Cb�c�Z��Z�cM{gũ�ڀ���k#�Z}ac��I�����a{<��K;$�Tq���F?s�~��J�8�Zx��>z�ǲ�D���.��.9��8�P`U�j}}��E���ޢ�@EE��R}�J�/B��r��6�s�#`��2s��yX�r���2G^\d0�X�t��Ѯ�4L��7����7���]�_�E9s���BӝC��:�^'D�;�so77w|��U���.<���]Ӑԓ�x6�i�K�5Hͧ����)��!��3zq�zvf;��x >���xx1���2I$FH���󯟏�y��K�������[���r�j�r����[æ5��9`���;�y�Xc>\�+ڱ�n>���_�Е/�/<�lT���P%�v2�r�4��2Yn�E��xC't��lE�b���Tޮwv�z�t5���΋�=k���B�I������g�~��dK��FܗÙ�k~g�<͕�~��"l�q��W���/�~���z�]3�o{�$�3�
��Y�^��}�,{%�����\kȃŤN0V�K�RZ�סc�jF��V���D�V:�:���F2�����;�1��n�=.�>��Y�g�$�I�������g5��Dy{��߅g��o>͢y�v=�b��^�ߺ�1J�?���3���6��15}G�p�!��3�����k~��
&-�>�nd�@����9?3c��b�]��3n�b!�5�xlL;�̾��oC�B��5����|2k�xw6_�0�⠆T9H�ɝ�lԄ���\]�����Sn�ӕ�]�v�Ȫn_�:�nb�HZ�k߳�P�z.�S��<j�Q��l���:����Z{zC��U�,�`$m:Y�g�*6�N앫z��d%f���O�`��k^r�0��&Hy,w{��/��=L�M�����7���y�0�nr{
�.�t-�s˭��<O4�ua+��G0P�ny��������׾�� C�BHH1! �!E�BO����߯��ǟ\�?'�������yN���Z��yP���1������iAO�0���6�Y��Sl�WɎv�jdls{�����YB�ʭ�z�����v]Mލ78�!�g"�5������ez��k��٤�}�������')X�z��Cl�����q��;F�����4gE�h�]��^]	t�`3@z���邝Zx�\��J}��H即S�cCI��0��n�t����8Վ�#Za�xd��c�yL��vL	�LS�(�L�<sa��&���Ö��U�^{����>G�%?.u����'���^�9�;Sм0u����t��x�U�.^A��AԦ��Z��ǃ��he�S���9ڏv{�����@�l��
m3f��٫%ů5	�dw8�JK�SZ���!��\A'弛[�����L�\��m����v-m�2Y��{��87T��,�k�3��&-��f�C�mLށ���\�ڑO�J���?�,z�[�vٸj�k�^ڟ<MsO����RW��vZ�Ν�9f*[R�uuA��wW;ȡ��·IW]I�z���f�����JCybX�x6�Ύg�-�I{��w��N�#yc�GO��7����/����Q+.s��nwm�[���]%65�;.�cUL,�w�_E�3�w�~�������!�@RI�@c	#$P A�y��޿�<[l��9"$NO����Ϭ'׾h���޷i�pq����g�01�@J趚��m�%���W:�{���_ￊ���'�~��XO�)|j���࠸+)r\/���fz�Y5ʪT�ɻ��3Fs�n�30p��3���_,�_P�E?��a���T�~�`b���vHX���n����p�+N�os�q��t�!��"D橷p��v텛��-��)�ѐm�K�j�sc92�A��h�kh��T�ݓ-��q�*Ԅ�^J�V=�V����@<<��4��ЋE�P�
|\p8�O��܄;Ը�B�}�>�*���2~8����S��,]�|0m|B�G�S�~'�~6_��b79��:w��v:�V� ֶ���L�UL������Yᕌ6sv;7,��؎uo_Z��	t:��}l�hv���1]��j��a�$�a`R��5�A`�M��r�؝�9��L�s~58����d�A�q58?�W�c����)���߾(|ޮ9��}�T�4Zo\�q��u��tEs�~m�+^}�h\���x3����������kʶns
��ID�ܺxl��cW���������^^۷X R�����؉�އUW����s���\�-:�OC��Ź��f��H]�ܷ`�SL�gqA�)�_��-\�d����w<���r@N�����i�U��[��g]��>������D� 2H,�bBF0@"�����Ǚ&��������d�孂�$`.`s�L?�#�������r{D觩���.���6�"C>k�R����]�F�C�������0�P۪n�2���%R�r	G7-���؅˶�0N�Lh6�f�q�{w�4��Q�hhmk�ޫk�y?b�-Aeyڤ��j��c��f��T�R͵8�75 آ~��� �r�+��?v�P��Z�`���#dV�����,����r�guN�hv�2"�,+���>y�C����t�Q6�z
<s�!j�{<�6�wVS�+�t;CE3e�ˠQ�[��.��8���f�� TC
���t�vX'�T�/&��^p��~���3v��y�&���Tzm8{����sĸę�U�f	����6��A���M�a���|Z32���V�T�m�R�1�S@{F���=;꧁:��Ū{S�V�6��Q����/�QL;2J���OT�d�W4�cVӰ��o�\V>Δk���4�w�u�~ǐ��^z��S]z`ry5#�j�Z��2j�ɵ+ݵ�����/�=��r��,�h1��.��h���e�ɣ30`�)����F(w���Yj#������n��Mc��r��./d�럳:���	�%>ب�j��wsn��̐ns�x���1��y�����N�񦭗��M���)���/��������OЄc	� �!�! ?o��������V��S����n�{k
�f��v��6��{�?s�u��c�D�gɂE�:Cue> ��m�g1������DS�#Ϧ)��mR��md�x5��c�n��y��UÃ��z��9���Z��ӓ�EoU�5�q��z���]y�IM�d�2�����y�$4�tƚ�Ẋ)�v�n�I�h�.Q^u�w<�^��Ҳ��������nbq�<k�'e��km'�R�4�o�"+�;P�3#���8(���F}k�We��jC��G+��]D�a�+^#��K�p��q�����|��.�Ή��QNO�z�|��M���0�n�4��I��p��ݔ����3�_I��uu�I>�g�;I%���� ���t_E=s�O�ԦaF���U�xl�
��j�f��fA�Z*��5��_Rٌ�����_|�v!��@b��5#��,(�B��H�p�����EPƥ�"6���z�1a��f͎���e���g�ƿ@�����jJ��#����e��h�4���?�hu��t�L�(�.hK��بx;� ��!:��k;��B9�u�G�R)��ݜ���j�����u�+�=��@��X����4(�Ǽ������D*�.�s����:�Y�¬�8������Q��fFF���t�γ2�g#���{,N�I��'�����=�H~��b!#bF$��������xz��:L�.t��H{m�,��=�^��:��^0�׉�l>J�5y�z)�?4;�M�4>O37��x�4٪��e0��N"8������Q/u����9�^��#�WP�
��.r�j7m��SϻǼ� ;����G��3��^�������څ�#1UC��C(z*m�}�m���v�-Uo2;���^R3n�#�ۼ7K�9ȏ\*EP��p2�G[��S�=���ݽ/9~.�8-d������&��7[��I͕�+o�k
j�bz��uy�&�?�s˽')�u\���@��{V��wZ杇�ke��{���ؖ߆vx)�qT1eC	�dh4[z4�	����Ej���c1=��KS2�l�slB�f�R�N��%�Z�J��������,BB��O[���ٷ.^=pj.���o�%:�Q6ȹ�(�Jꡚ�/s5V�펦�ӷ�z�LB	�e�<F4æ�z�7s�ǔ���h=2�0���Χ��Z�������j�zk77��a��}7�"qk�E,=�'��0qzǞy�O"��їfkRv��j��Y�#b�q���C�:��
U�U��0I�(,7p31v��vu���J��&�,�o{��α�r)9�.��]�6�y0!���1�9�-�t��x��K�1KsR^�f�c R��~�Oz|>���5׎�ji��}������?Q$"��E�0�H�HE��D!"	d/����ߟǿ[����-a�]%�cÆ(k}j7��g�q,��Q��1���)͍��Nnȇ�<�&���9~��CW��N;z58dw8�}<D�W�D�\A'弖:wԳ�Ic��}�6��j���:�z�I�cq)1�K#�.����%霾���8mv'���je
�gt�̐�	 @r״.i�޵e��^��@�����D�O^����ާI��L��_�=k捣�0ߞr؏��,+=�j�D/�^r\[4�����&.��e`�>���uO��ݶ�m�<Η�
,�3Y%=�V�k�2��8��lY���*�2m��|�Wkp�r�؏	O�YzY_*�ѭ_$Ό^#CY��T�f���ϼD����MY��jn�,�܎c@�!��!"r�V;�<�n�th�'@W�Vh�ֳ�I}����\u���,���^�dj۟�j��9M��$�D��iKr��]�����X����ò��C&V��qg��L��pz�'����8���,�_��G�7�AVl]��: X�q(.wte��_�~>�]��������Z�����)�-����[��ӜfC�aw������xޚ�j�)���[B�QzT*�xO/
�w\.�-�Ĭ�g,/a<ϊV�Go w�C�,�pG��%q��8�?,~�b�}>�e{�Mc��t!�q"��+;�Gn�b�oAK����0^-(�8��o5�r�Fn�Ԕ̍��pd�{w���B�]�6�:-��+8~��W5��+���������Ǝ3vx޷ͨ��k��L?:*��ﱍ��u|Ԓ���,����Lm%�y���v�l�];�&ã(����zrx;&����f:��>
��[�ɼ����Y51�F,;VyzP~]
N�_;��m�"��uH_S�0m�r*�1�p�
_f^Î�kn���a��
��Y�N��\�5��ܲx4�>��*l�*ayu���2������ֽ�2���D2<�G5���u��p�.��c�q���2��Խ+�|�k3I:ʧ���"���9��Zrt%\&�K�l�Q��T�)�ITׄ�:l`$�煨��REO��7�Y�n�'�:��ͩX�n�f��T�=(�P�ޝ���Y����������3�I�Uy���p��}r��tZt®#����;�BP�oc�����V;cKҭ��b
�ϡBP�p��O��J��{*���w{G��6U[�h���9!-6T�$R���;�r��n���Y��X�:v�U_�gyd͞�^:�h��+��fv)ϰS�l�Y5-�Y߁�n��NWm���[m��l���S.kV�WҬ�bYg>NУٷ�{��ח��Hf�V�b�\�#��n*e)��ƨ͐g _m^�Aȿra�!��Tǳ�-��4(�}�V1NO$�>C�d�J;6u�Ně�L�ɜWz�.6٘�/�%\-ݸ�Δ�#J��W���O�g�����Ӽ$p��[v�PC��o��P��Q*�-."��;w�^�d��P*P�z�!)l�\�ԕi[��Q�	Lr�Pf*6��x9n�K�O
��;�^c�cʊ�>�r{�i�C��b"E���6:��Ry�����a&k�C��K=��=kp�K�/�ν\dE:ũ'Ŷsn�}�»�Co��4��/SA���\>���Y��9��j�4y�Hk#LJfM�:έ����^�6�H�5��Yq��k/�tj��djF� ��X"Mٚ㏍iܺn�aň�4�־n����KdeH`ɝZ;)9₡q�W�dق�[WƳ�uZ�gQ�����`����h-Xy�)��E�:���Ӊ��y[��=/��R�/�M���IT�r;_�z�ci�6 %L�x������2[�F�N��j����;��U�@FU��ǔ/p��&��Y���֍ܺа��K�k�g�t��꺴[�")<#��n�	�Q^�J�l�`Ʒ"�2N�NNCܪĺ۫�����"ֵ�Ύ^�-*��j��T�*��5iu���TD�m�Z�M>O���D
��e�T�VT����fd0D[Z%�(���%J���N�O���>3[D�aQ�M�'�]T��E�Z�ŀ�ʕ-���3N�O���7ƋR�[h�QQB��F�V��+-��*E5���k#J#my�%�'���yKKah�5�X����V|��~heגi`6%�!j٭R
*���*���l��J��mJ�Z���Q�D�b��vr��e��V�U�WU�+b�Z�΢Uj����J5��Dh�Db�PPm�����j҅�̕��&�Qml�P��jŊ1X����u�7Z����ʍ��^��rR�){eum)l��m�ҭ�V:�.J%��)�+Zʕ�YU�Ym�u��F�[X�ƈ*�B�,UFVʖܚ+�R�y���-6YY*��H��+zʂ���<�O���NE���P�k�p�h��߄����
�����+3��Qo��1u��P{��z%��R@U��"�Ֆ�����4R��D9�d��/z���Kv��m��9�U�C���\���ۻ�x�r#� ���HF2I�bII �H b�0�8��x��^fE�&���b6�H�:�;_�%��Tl��qW_��!�]���x,$���UL����X����	hwd�H%�oN�ǧ=�j�w��c�x�۠����Tc��*��]Yڦ��Z��a���
�v���*��Rש*��d���7Z�p��;�D.����ېY0�cFB�M�=�Gz���g8^y2��t�6�atsu%+_���w�#�V�g�wO���i\[0݉���j�#��� NT7�na3b,<�;�>./#��Qm�@i�wh�l����	�h��7'VF;���y��wyj�*e�}��Z�ΥR�l(䣛�ç-؅˶�@fދ�D0e�EV��g��W�K���ܪ)�Ŗt�ޔ�;��~���/;kk��!*�e[�s+(��xk�E��8�e�NԌ0lc�ڂ�t\C����Ǥ�ӳ>�������ϻF�^�ԧsEfgl��B-zT��7��x���:���@�� �瞱ٽ�gݪ�KW��N5$��bUO��cs/(�.�OP��A�/�b�;wv�ǟK�O�-+`�ˋ*�<K.��0pݐ]�߻���Q��{�'n�.t�ۂ�4���zX̏��D`G�hr��
��h�6����Y��ߧ���T��Eޕ�\���������o	��D#ks9c�5��fY��<	�7AgA����T3Sn��20���Ha# 20�H �!$��������?p��_����Nf�/ ���$`��Ӈ�A�t��%�~I�����Te�֠3��汮�Ns�l+�^��m�'ɣ3*��ۨӴPA��Si��i(�:z�}M���霓�uj{���OP)�Р��55qL�Q^��,�$�>��o��[kز��G{�I�~���gt���*K1Pk1@��]�Q��w�̦;⾥���ƭD�mZ]rX�U���6�,�V֒�ֻ�3-�2nկ\�2�o��]�1�G�l�^�8�QY�â.�����;V��/%�{�m�$�u�-����vV�^]頨v����;��ZI���:���u3��>.`�A�4��I��a(���P��U�5��NC�;ˠ1�zJi��j�5<�St�@k�ѝ'q�[��Ƴ@�<���Ins�S�h	+	=��J�[I�!�T���Zͩ�����z��D��Qp<g�L�˾�F���hw�|]&r��|k��C�gs�4���)�߸�w�տI�C����"}ɗ���PO<�ؤSW��z9r��<$d㭧fJc*	�]o-tNB�h'ly�����珆u�gG�hk7�3:�z�8�iT��x*m�:Ŭ��U?H�a��Y�/�����Z-!}�u$�%+. �[�r�Bͬkn�Uz�v	����G=���vu�J>������Kc����w�y�����!������Y ā� �
 �!�����
�����}�lv`;}������$��y��^���B'�~4U����Ӷz���uݨ��Zq���E �q�g���N���ξ(|�s�C�α�?O6��ς�M⸊�[��vyyGW��hc,��$�k����.���NB��0,�x�#�}槏���w���/Z�'�z�2shu��n�L�Kk�ߐ>��.-,�@�[x��M�����ڿ���F ��8��������@�3������1m���M�9�gN�wQ��F��Y]iu�������G��g�Z�m���H:�g��6����Pf��g4I�<d�nwW5��]-�%�EL�?m�XB�g����<��^Ey��k�?:�
}�2:t���O��6!���?QIOzZL�뉯�g�At��b�R�D��ӗ�~RU�h�wt�t\�Z��K��,�[c�k
e���~Ь��k��J��k��U{��8��K��6�l��66s�E�<��Ô/m*�qw�շ7^�N��zU���S�qFoE������p=��E8��w��S�z��]�� �����q��oZ1�[��Ln�0�a���q:)�LV�UGnj�qj u��L��L��@٥��~p�{H���,F�~�<��������7�6zt��޾������o�h�FA� � $đ� ��"�BH�����~����,���l�@��h��d�훦|��	?S�M�K͜��r6��0�s:�t*WnlEfR"ջ���_)|z� �V@!��f�7T�p,��P�=2��J}�	��Rn��V�6l@n�
���D��-��}ř�|�Xn�yO"��s�Sfqt��:�z�|)\�b�c��X�x-�%+(~gwm{��DF7P��Jn�	���s�by7B.��cG�n35d������Qa~,��1CZ�C�QM!��~QGW��>�}�QD�R���i�N�h���@�V.����q�oT'��;�',8b/�C��oK����3)�X��O^6��Q��c5Լ���M��N��I�NB��R$�@�;+�����ߓ��,��n|3���]�`:m�$C�Z��d�Y���pI�ko?�}x2����D�ǅϏ꩹���[ݕa;Qp�x�͎���&yP��3��3�l{�<,�����@���+qTa��)��SI��]��
��o���=<�[�˵A���1DP<'���?����|���XB��Ҝ�]K#'S6t���E�A���[�{xُ.��/.�Z�bZ�':k��,����"vM{��%�/�C@z���M�{J�k��6�v�n����8��++!��k����˖���_����~�D?,�	 ��H�d�A���$����9??��^9}�%F,�(����}\�_��l�BF��5�6Ξ�a��DKl�Aa>�T��q�:��T��^`⃝C�ڼgr�_�LÂ�U�H��6��]C
0�gb[g��=��ڴ��S�b�������4���U��T����%4U�	�%t+��O-�xy�|f��u~�q�fwp�-l��ga�~P8����t*�&��ɶ�K-X��U�������}_�w��jΏ{�G���/���HQ`������p�=O��vd��3-��85צI��t�v�_8�̨=���%��+�c��4;�G�ܻeL˞��k;�Ѹ�ü	��}��/jf�\-#��?�z#[&i��v:�jp�T<����+�4t����z����yD&힗�"y��ڍu��ʼІ��.-�*)��R~k����Z�֪w~q:�pDB}n5=�3R����o��|γ�Blx=�sg�ۄ��Ur{�%����[�Ƽ�$�:Ǝ���
�Ľ�w�6��
4�'����3-���E���U-^K�:"%(�ӱ�`؅C��W��}�):�8�yi�w�OO㋓Bm%��wl��%�v�0�Ty�w:U�TO:N�K�`>;3����a���>g?z>��P}��+Hܠ�?.����(��:qܲ���@(�{����V�`���K���ٰ��5W�޾]���<����H~�F$"� � �	 �'��������o��}�A���Cϛ���/<�K�kHgz��;���z����F+���uc�2�ӹ�NU��n"�دt3���H����t_e۟�='��]B��=��=�[�b5ݴi���y-�'����ie/DΏ��Gs�o���^yV#����W[�k�����ͽ[փu������J����#�DjH�o��2q�PZAm�zONU� M�3n+�9���͈��n9�K�-���M�oA��|���L�eS��{�[�W����㪵���azj1�^O����3[�]�����)fӥcPz7.�9^Ȑ��
jY�����z[�D>�q���nK���uй�#
���,�(�3k�Q-n�%oU:�yT�h���#ND�;��n}���Jt������ӝ�ȇ�8�\܎��*��t4�ޖ�k�Џ^r���\�bGkZ�F;�o��j����C�����I�m��
#k��@E�nv����g��vz/��ۤb����)9�b�M�E���[e�6���Aww���u�t9���Fo&)ٕg���ٙlm���~Sw��no��T9�����3��:<�h%���:�U��B5a���*Mu�j�eA{@�vnS<�s�3��l'�x��"�>TenN\��V��0<]���5�2���|rL�,�����졣�M��eT4Ev����}��`y��b	�X)#�,�����eB�T~�F �����?J��������j���9/�@�������#L{��~釔,��Ɔ^zv��.9���C��G��k�T�+_u)����k$[1.��f;���]#��(E ��g)�o��v�vMU�.��ʥ�q�E�g�-��<�z�;-��Rx�yW[��}���Ť��<h/�P��*�?ۡ\�V(�f�]BiOY�4tD��hS+UW"2n����<��"R���:��_�ψ�ϼ���)��+��zxе��2B٪'0��n�X���]fǢ�\�]���8;c��zY���&���ƀ�vyט��篛/�<��|M��q���c��.q��P���#c�z��v
�"�8�[����&9��Cރ��!ֲ5����������f���@�y�����+���xt>��`l���=,�>ڬ���������X�^V���M��#�����*π��.����_&�:fG$bwF�',��}�j���%��ɉ��@��D;=�UGI.؞�^�%�����5��U��=/��,����!iY��sWG�M�O*<��ojf;)����!��Y�h7z�tqо����z��7�d�_����t��� ��:7��#K�	��+E����er��#�����������>Y���u��E���U���N��Q&Ü3n%�\�>�����$H���D�ȐX{ߏǼ��دt*f�%t���ٷu����z=Tٿ&f!F����=v�p���<��q��L=R���a��~���x��C~���zZL�K�����
����_�}oWm�Bn��Z�v�l5Y�U�@^ܝ{΂Cը��a,�[�q��ˇ���˫��>��Ǜ�W: .m�����%K��F'͘v���t&\��)?^*�X}�
��~յ$^C����_,t̵+yr�9���׵��C�-�4
S�Z���sX~�I��"qS5cһ��u�4_)�W.�L����W^����Ї	ru�F��f��9/��9A<S.~�+"���^R�Xcy{��ۀ��Ǹ����I�05���>�n)�߽AWzSv;�3�T�!15��s��¶���G|�͓��*����^��<F7P��x���Ǽ�S��{�iXdʨ~�p��Gz�ӑ���Z��,�9�a|ͭ4<��K?<<���w�J��%qRp�ݥ�z��ׅX�.�K���/����}��8g���Ŷ�ln��=��۔��+3ɟ^'j�6�eu�5|	o����_Eu���/s[�8rM�wT7VN*�LΣ�z�b����^</ ��|��+��/y$����v-�==�ˈ}n���싾|ϯty�ö��d�Һ�'���O{�����{���ߗ�v���ԟ��`1 ����R
����wu;��>�����uݖ����	H?a�G�*�� ���n��-�$걹��D���j��1l��
a,�-�FWSb|��]g��O��]!�r��>��ıc���V��l�u<��{e��~5��'�u&�s3�x�����c"�{vF���&<1��<�?+#~������\�����Y�B�χo1p�"���1�ug��Xsr��3����n�_MkM
S�⦶@)�k��6��%Sg��3l������̉��}{1k�����`�b�����U�4�8 ���TK:�ax2N��MW�O?J�����7v�����z*+�>߹	�����WN�@�l4%�M=���<Z�z0"ѽU��b�}d"�m�K�j��n�*���8�MjBm�%t+ƭiKr�f����K���w�N������/X�U�
b��2��C'�1M2��X�ݭ�{���a��-�73�F~��ϿW�I�-b]ʂ���Q� o����@<#�K
�e2��ʟ^o�c��Pgx_f������4n���b�������ʌ|~�C�b��#��U�}�z������y#���r^g,JӋ�'��z#�6��Jux�|����y�9�nk5��<,�11o�}�}r�bKNY���R��J=����k0O��8��󱐴S��X���I�9��%KG\�^��@�y��{�~�?1 d`1�bH#��2U��+/��R���M6H������q�F����;����d᫴��ŶU�ð�9e}����$���qv/)��ˣ���Z���P��s�S����0aQ�u#�x�������ܲ�����Ț��z���������D{��`��ګ���<k˒C\͕-��O����*�X;�m�˪m�2Z��wR�k�8�QIG7-����U�6?>������·�bvĠ3a�����HP���L�_C���w�;�������gwh��:+56����wc�1y��*�5�%�W�0h�9����||!�.��^�='�;k�sd�[ȍ�J��T�w덫=M[�����J}��t�����0������Ckۨ,����f��:ih^��{}y�.�s�����s:Ú�b0��=CC����=���m����5�cu��k[�����[}./>��c��!؂{�ݻ�m�!�r���DP�Ǉ����H{U������M����p��;��0M��|i�Y���̈v��Ɲ��!�}�Y�4궐��e���
����e�?h�5�U+ɗ;<7�l��-�%���I���[ۗ���[���ȏ޾dl��@�N����B�̆s�r��r\��H,�.��R�z�e՝:���y�X@���kf]�aku�/t�f�1�9�  ��Z�l��N3�yr[WiZ����X5��F͊CYm�8�Ҵ��<�v��%B�o��t����>����y꺟Zɻ��+4-���0���z�ti��j�J ����K���{���%��B�������[�/�/hkZ�l�a�m3:렰�s���*d�I�Q�)�V��nՁd�xqi���1�CI��/������m:��y�4�9}�^�o`*������˘�s{n��c&��I�o ��w�٢=b)<���Z�����ʸ�����`��r������%Y�٠A���(��;^^;t�K��O1�����mm)�Y�Y}�M��T���LםI�����U�`8�8Y^C�-a[�c.����f�ڵ�|ӈ���2N�� ��'u+]����D9Fe�:�����j~�MJ�k#�m��\&ڪ&�jD'���T�Ξ�öx�T��f��n'-�;�!�Ko�\L��콳ܩ'9,54���#lU��xI�YeV���ŝv
TUf��.	m��[�
Me�pi��N��;G����id.e��N_Uؠ�TKH��A��t��5��s�&o���I��r��#�eEp�ܿ��݂b�c��88B=���7�~}��y����ͬ���{5�k���p���TN���2�^xV�R
nC
ܺ
���h��3����Fff>7���-h���-��[,|��r��uLO�]��,�^�{�j��܎x�>�	�J�Oa�u)׆�ؕ@�W##S�3�!�;� F�3���6���'�7�Xf��DL�sl�%�nu���'��x�M��#��T�8�Ypựb"Tx��q�� W�+�};x�C��ڽy� Q��Q�y|"���ą��;�ǚ˝u�떦C�X��X�;�֮�(x�B��J`�&�f���D(0�3E^]9�K[�٤�&� �����M��wF�C�(:�ƃ�R�6Sl��Т��{��%T�7vQW<�|�F�#�ov���]'
䁱��5���d0��O���,�O̦��u-�X�<p��2��^r����8،�Z^����5�opΝ�F�G��\��ŵ���6��T�x"ȴі���d��jaڊ�ۏI�GN;���b���)e����@���=������C,<�1�{/Z*��r�Won��c��vy��|JF�D��_.B�(�6�m��4L��)��$�}/��r��Y���œ��E$e�,U�6�R�ҋQ+iQT�`�_�f|fr��m3Y�I�d���t�>��*�1�Z��4_�Y��Zն�6���+b�(5����J6�-��h���R�����|�L�5�Ͳ�UEDUh�hV)R���VE�S	�j[V���*���j����g�����y��1�3DA���Vі�Qb��T*���QV��me�f����|�O'�#:��Vص�%��l*7��j��[W��S6%m�UH�[
6�dTee�Z����Q���p�K�m���[AR����5�,�v���)[R�h��QX��Kk
ʕm�҅*�-�p��Uv�iXQ��@X�b����lb9�Q؈�)z��[\U*���6[d�̙�)KE�XT����lPDqK:מp�
ӭ�^{c[B���R7YDEAX�"�2DA@�A%�C@�Tb�os�2�S����}�Gڕ�����z���{��)��71'��r�l��(	��|��~��U_���`y��o0f 3�-���5U���|���qP�qǨ��?��r~�����pݠ��ӧ��)�;���r�P�]�Ԣk2�N�k�jIm;	�ط��zw��!�C�"�2E5�����t��ǃ���+!n�cF����p�6��u���vz�;�xֿ��&h+�p%f�>�1!S@��+���D��ӊ+���!6�!����]'���"�i%[������N#��?���&��w�0����ߺ�!��ξ��\�b����%�Z��;�R{�J-?,����-U�֭㵰���uf�oo��l*��A��U����gi�¬�0EA	�>���������.�Zi��T�n����!�F�4F/@V)���.��xmj�ly�錺.�x������pQ3�.xɻ���X�%�`������X;G��Yw("�.�a����v��&�x�1��cY�u�4뤔�[�'�-�|�����1��G��*�0+��X)U�����O���u��V���]E��[<О�ٳ��q�<͕�~��-�"'B⼏��*^�~�^��΢5�N�}|�^sJr�4����k�F�F��>v��gu�B/��\0�0>�����;󦻰�>]��7�C[�T,���hf8c�y�&���s�����#h�O�K��Y�&|9!���{�y���}��~?Db�1��Id�ܺ\��T�d����7�v��u8�	z���}�A�OJ��*yh� �i��k*
�v7�bڶ{��Í�5uW��ʩݐY<����{��c����c���z&y�Ѓ6\1�^JlxSny��1�����1�g~�c�t ;@	�d9b� �����~��=D��<�Oބ�.�+��(�C�(}3�/6������X�j�o�15@���>�Bj�|���vfDpn��A'�t>-8�m�����ݯQ8���u� /y�_g?�~q��~��d��?�|1����~l��V#�77~���^,�*������n��
W�A��v����B3n�ҪЈ���MDY��VQR����:g���˾lS�oB�eV��퀖Wz��D����?K�.mtF���	���8x����j�����4���Lk�LIln�L��<��7"�����l���QR1E�/q�Ќ��"�;^hM��q��3��Y����ڮ�k鄟��O�7�����E�Mi�ǧc
��&��vvJ�=�����%����=	rud�=�0�T}�%:�YŇC?bp�r��!6��U��N,d�`����t/9��)�>SNTą���E|�|Xx�ܫYL��ᆔS��������8bnlv���ǎY�&�
ֽ��,�������S:cn��|;ON)ff����_>������#1#1!;����d��ɞ��o8w�y�_~Kk��_}�:�n\k�K
?�t^�Pǔ�M?��p�"�ͯ]4�Zݾ��6�x��Ĺy�ˈ~�m*8�
������Z�7��"hx����{�?}���O�}oWv�qG/|��`�!Ѥ|3�mi��GBi$~xy�A|i�r\�^�m�P��L�'�r=��D�­S������;�e����Q��[��oWf�D�q��B0Md��7��{�^��o:��X:z�z�I�cR3��K�����OE�%��ގ��Lr��}eR�D��0u0��
Zo����wZ���1�≂��r�]-�&usW�羭߸�O���m����	�(:�FDF��vO�.�5N��vo�Cr]Ʃ�P�}^	�F�r�ْ�,\Գ��ϮhD{`6"T��NAO�J~��6�êk����)��cN��'b���O���"T�J)�>t�몈���d;c�]�V��;��ڦ�Q��Ǽ���͐�ы��W�����`��~�J����Q����-��!cV�ڴn"������8�:ߘm��h�y޹�b��5�H6�ɞJ��f" �5�8Z� p1E���=�ܻ�����A�,]���g���v�u��e��\/O5 d`j�Jh�9ˤv�QW��L�ܶ�Z��<���￀[��0o0��"�Q)���r�zIj��jf��鹴�Mt�sa*�V>�hj�*+��ͳ�]j������Ӿ4��[K�g`��)�\��{{)^6r�NhZ�e��q9��t5�v�ef[uo��=���#����l<���A��׳F�w� ��[ �tIa1�y2`�>�ʾ��;qSn�䪙:��q̜`��D�^�{����7.�B`&\��r���+ߓy)�7W��k��D�P�Rb��=t�U)��%V�W��9���w.1���hI��Y�.�D)�d��I�+mU/�CϏEŹ�E>y�R~k�������U�OϘۯ�d����|�Gv"ͼ���\-��?������E�<���=?ga1B	S��
 �GH�zT[soUQ�����-��Mj�glq!y�785��1ܴu��l��SM���T�,����P�\��l1�h�j�OoT�4�_m�|5�w��Ƃ�t
>�/�E�6oU����.���]{�P�ձ�@)�4��e��ۋ�mbD@�n0ht_X	����I�1q1ϐ�kަ�k��i���F�~o��Ϸ픟#K��yJ"��/YS��+��q�Pl�=�+h-��N#E����X�+�*W't����qp��8�����ߪ�,��:�K��<�sC]�D&?^� �+��������s~��oy���B���eo!����I<{m�al���ތ����^���~~!�1�+�P����e�w�7ӯ�0��P�#�y�:y+�^�P�_���iy�(�5�s�ٳa�AR�L���ۻ�=�������CF-��p����v���^m�"F		M�BS�y�ˑO��]CNڭ���K�(��}��'?�?�	O��~㻻U�L�D��!�{��m����1�,إ��{���5���0�!/�>	����$�~LMP,b��|�~�r��}+�^�d�M�"e���<�{s��)qS6�F���vط���N�^��@r�]FM7�����3*�wiR��b��L��]��{�M�1�C,�wM��U1���w��T� ���`C���`��+&NɄg;�UI]z#5!�UY=|�4�vF�1=oc�):/�j�No�m�%9�v<T�>�k�)֏$$I�eEڇ��ܦv�m��4m�,w�^���k���.5Q��ek�Qi��"��o�X;W���q�E>*mc����4��bh,#�Ri��}ˎf���v�w%E�9���	�>�C�G�ﳉ*��K�0T�������Э�Ŗh5���aLɇ���<���p�0�'9=��)]�Y���n]�;;�~���ݩ�)\n�ת-�����eR97�W;{u�9�sV��ó`Q�P\���l��! ���]�x������#�g���ߟ��9�~���4�~�H�������B\�)��M�q��iQ����.��f��P��l��#��׫�n
`�W�9`���wH�_�?��hz�}ʄS�ތ>Y���(��Y�P�l�F�J����r]nSI{H�d���Љw��������1-��,f��zĲek*;����@�*~��i�f�G6���g�4	�ig�VW��ѽ$j�]���������w)��R�5Ec�~��BI�N1�q�-�k_����󰗯�s@����!���k�'C�<k�H}�-R��d{�Ͱ�u1���%����Y�������⚴w��zu���^x�ؒ���&*�؞����5߫��˹�N�g�\��.p�>�L�x�^���E|�{�4����ϗ��OL"��`?�FfS�[O�]O�Y�+��7��#�^���
�vy�-l�����6��y�k0)��˄U�Y��d���V}r�%����7��a��pe^*i� �j�t��KI��m�e��}���~ɵ���N2���ʅo+vi�l���][�|��³=�:��%����^x6a=]� ��|�ձ�����
O����]K����(��Q�ru��s���2��u�Uwhk|���4��ȁ�Sh�*L�s;Em�l aN�_�7/�|>��`�`��'��<]]�%�͖��5	L�
�n?�B�ڟ�:"}�Oj��A�=z�R}��P��U�)��<>uC�ڦ������3��n���Ô5�so�|�i�c��>�gLJlk�t&E�lR~Œ+4��qo�9�)���T�Փء�Z��va�\V?|P�x~�\��=��f脟
���]����sP�rn�ؽ�i��]Ĵ��{
�ǆ!�o�A�h���$^Q�D8��<����W�Rx�<��O�E#�6��̈�\r�~M�F�ܾ�A_��:���\����ű�V� ��a@���:y���w��|��}�|RQc�ToP��z.�����r�:�9�V��]^Ek�Ò*�q@��%,���a�?���M!�������;�ٽe��5e���ZҦ#]5zf	ub�����%J�|���~��),$b/�b�s�W<U57a���:q0�"�:`���y=��)9��]��[���ZS�q@�s\����L�w��ȳ��+�sS/{�e|��ȃ�@�:��������}W4ɍ�\�`�k��2[o�}b�z�ʛv��!�A9xa���A���Eu�S�TZs��߾�(n��R���͌6$e�:L��c6�����yK�' ����#s�����3;�>z�'�~��;��~��Rmi">�/x�Gs�:{owi>�W���ָiد뚽�|��E�e�}{����8�����w�߿[���1�(>�X�4N�ʚ��%Zѯ^��M^sBQ���H�T����,��i0<?(E�/�[÷7�UN۱5��/H�g���HJ� 楝�tK>���l6
0��ICeS(����v9�u���a�.ۯ�ߟ�A��
4HY6���t�:a��DKje�ՙ�. �se�Tw/�e$�z�������l��;�m����*e^�$NP�X�Q�v/)�n���@���73e�K��xje闣 �Ը檈��USkg	���MH�um|���O`�=�&�/������7~��Fm����8*�'Ÿt)Ưw)d�
{�]o�+n_e�j������8��dx���X!d����{5������h��L�7������z�o{��A�-Je�?5N{���a�J3x׭�XX�\G+�h�~����N�*����r`�++òDȌζ����Sw`J���I��1n��\[L�E��c���"�;�W�833���;S�5��Z��eҮ/��3e��?6���Zw����j��&V4����Hsթa�z�w��e�?6�QI�R{rpk�*�1�s�[@R���^���z&��Ҟ95�檽�K,ն��� |1q�\��Α_k\�%��p�1S|����[�|<&V�u�e���7�y�y��y�y��X]���B?3ǋ����mu��-QoW�"x���b	u��v=T��WF��\���i���LcD+�C�� m�w�
��F�+-�����c���s���,Ii�"���F�U=�.;1KO\!
H�.#��+��w0�˼��SWƿE�6w�ۢ<H}��S*�WgB��W���=%u�j=3����v40nb�5�?!�z�υ�cKӧ��U2�6�U�����\[R����*5��ڳ�?u��=�ʞu�{�
\k�����S�Aa:�f{�b�kޫ�*�ܡ��/�����j�"��6�#�^���h^t
"~���}>^���-����Y�i�hi��M^�8�{�(׻l3w�n,�[4�IV;�9�ͳ�q��R�=�4��;� b%�n<�������9y>�̪���.��*Pm�lGn�E��Ҕu�aL�V��K��zw�^x�|8�Ն������y�������Ɖ��h	�ƞ:j+z�c��3��{�(��i?}��s�%~T�b��C S\8��z�X��L��1'rϙ}���a`��!�0��m�ǯr������s��p�//�W��b�m{'��'9�EԧݹZ�����5�DV�la�A4F�؞�m���e�eչ�X@xB�/=��GT�u˓��L����mN�7D�>��u̷��6�c5cnm5Gl5Xx������3y��`�`� 5e�䙥u��މ:��2j�ŵ%�M�#H[8�"�2�f��j�M�ꭽ6g^r�>i�U�t��; �<+|�N���Si�l	m��b|�)N���͇�TM4����f�ra��կ.��v�d �-F�����~�K_R�NJ"�@�V���vLX=�i�)���u�j�t�=�<���}"2}�q��3.y�5�KrP�?@�0ZS�ch�}�a�z��klo!��.�
��S"s�,C����� ���Wt�;��Z�t6Q3�^���
�)<{�GC�^�r��Lwp�����hD���˽cn�rh��I���>[>�CY;F����=�d�� ��-�|�x�;�Oˈ��}忝��W��OQt���5d?B��礪~�L6��4'��>��k�p�[?���>Ϣ1�	��WOc�l�Gf���YjY�M>�\,Q^Ǣ�mp��1��%�-��H��&�^��V<3���K��G�����`��l�$Le{R0�ύ�z�?������1�#��2��,7|7Ǜ��ʛ��	�xu�X�oP����6��0�:�lF:<F�ms�o79�/���4e����N'��8�}���[�r��K����b��5Tx<�g�{�����hM橻�������r�)����oG�wy�^�89��Hu�=�C�5�7�M�[��2���o�m��F�ΨW��ԣ��<��퀬�);�ȷ(���H�do��1ױ_�嘰d���W���ܳ~-�/�G�2����'�9��ؚ�p�;5]]F �.�`�T���d�sV�;��r�w�*,�Ԥ;�_�))��qr�z�̖��AXo]e���㫻�0��Ne]�h%�-}�4;�����໒*xٸ`P�8�}�j=�_�i�bY��v�-F��aܔz�=}��Ź5!�'�ۼ�_x�=�p#�o���;��H��z�_�����3T)��Q�B�����!��.�צ�����Esۉ�ɫ�6Mm�k���Y���Ǜ�GS���������=nU�c��%���83�u`Tֽ~-�4*y�ðK\t����:jX�Gw���Ǻ��{�F��l[:٦`�K��M��,�438�V1���}&r03���~�����L)*i�Cf�.m�*t�{���͒M2�fYa�Ӄ*�VZSH����^�l��ù# � �o,	��=qW:d�ZT�ov��ҥ2��䨚�*%����F3EF�wp�t�H�uƱ�Qge�$��3��������/?=���,��#���ߪ�wJ먖ev.�Z�N$�p�vH����x)O}�������K�N��s�v�!�H:�l-����8��v�����>z��(��;6ge�k�G�k�5�i�]:g�p����p���m�:w��a�;�9���b��;��ژڦ#�ړ]N��l���Ng�2"�+
J�Ħ�Fȸ�v�w�� D�e�X;���ӎ論؏�M�6�\p��d<�Y[s|��W�v��~n�h[��p�wQW�w�p5�aCyH�;������>�ػ��F�{�+�ń��=�^C��c��!~ڇ��t�0{˓J%u1�v6X���oj�%��3�"���o>b��r_yj��c��t��.���n���;�>�Ť��P��2ќ{F�X�vA+R r��+B	�Q*; ��&wP�[�^�nDպ�w�K3#�J@^�㉳3-ű�m�K*������p���S��U��	6j��[ő�m&%��i�1�v-c˳�����M�`w�M�Iw���u�"W�7�2�[|���5��He�S0-��ѥ�Uׁ����D�z�=�����؝a��т�eq��;�G�������~��I�<F��|�w�����$4B�L���j��H�r��f/����jn!�E�G�hv�|���]�z�+>�q�w	�4�H5�t���H�u����R*$#���؏I6@C�ۊ��.�X�y��X(]�����K5l,PTm�n���hگk�`����]�O��?��1����km�D��K:�Ң[Aj6KQmj�T�h�m�<�0�#z���Kkݎ-��,K:y>O'�ȬUSġFKւ�
1rڥ�em�R������3U+�������O����1�񺰥�GYu��X0G"�ƶ�U�6�-ʭ��c�m5U�b�렙�g���|�CP����F۝3Gm�U�im3W�0���m.b1�Z;V��j���s�6�A�]Z��tZ2�ݻ�AJ���ks�D�Q��]�m�%J�+���&����E��2+�,׵H�c̠�F�YKJ+Z��0j֨�mb����Z�Z̕m���D�Fұ�[

֨�jQ
�i[b�*��Qc^��m�E�UQ���V�m���sU�����iR���eX��T��TD]mJX#l-�B�B����ٻ��Rޭ�'m��Ҥ���b���Cw���n�P	y��!�2��e^�r�]�Ya���>h�q��%T)��ukE�a�x��9�h'J88��,�O�qkk�ܫ۵����WU/|�;��7|�w��#��f�|��ƻw���1ן���vP%����`&	�����/�\�r�o�Q�`z���v�����<=�u�w�EKfsÝ4}4W�]�T�������!��C��)��S:z�[��|�T����g�V0/Ӡ�C�T�Pg�&�m�7�2�1��(�s6� �ͅ];<��u^��j��<��{ H�YE:�{�Pjy�O�2��2wy��8�Yp�mT>k��APC.Q>ik��jK�:I��5���c�g��d�F��Eh��ٗdZ���.S�*m�P���A�=�/��D�S��[0��Wu<?Vs[��d��T��a�4��d����!�%ީ����*u���Sgt&I�lR~��h^�m��q4�<�Lm�7,����[N��ݻ�4[z=����gŚ�Ҭb��=\��P��i���M����i��X���׫��p����>��	��¡����2��4Y�͋3K��Y�U�t�P����gy.W�E2�)G��}챷ꙍ�.9`"�@��ɟ��[E���k�L�[��B�On�Y���3	�{EJ�X��^JV���,�ʹ^U�åY�����F�a>���mf`�of\$���Qȭ_l�A�AUu�ئk$;�tpU�ͭ�3�X�5��!�@�m�w_UI�c�f�����itz���5ܦm�N䠙����� O�goo�?]�<��u�S2��Eiý� 3w��AI}*OH}���}��y�o7�y�<*sR\��Êk���s|�'o�����U�,�%��9��	��[<_]���J�wkc/�#f�/�S2�Ls}2\��f���g�8ػ�R�o�z�= �;�e���E�&qŪ�O�T+��ݴ->:	�6ؐ�3g!��D>�4E2���ޢN��)1��f�mO5�S�f��Olt�.h���j����w�	����
��'��� ��W�~>����۟-��n|�-�����uV8A(ַ&y�dԖ��~��(��s�M|=�C� �XD=�6��%K����cZ�ks����/9.-��M@9�gu]ϮhD{F�4��>4���AD��0���w_T8�M�����32]�۰��=��I�`X?E0n�c:s��R� �os|�c4Q���W���O�֨5n/�����K;^�c��(7X5"r����>s����Gg^ݨ��Z����I�#12^'yf�~_Ǐ��g��#������O~Ě*Ԅ��?^j79k��4�©�Ɓ?�����٨{�MxFy��>����9��gl��S�����e׆�q���֜�6>�=`X��)�W k�A��oZ��Z7�h���J�̄�o{����{vx�����4�qU�w6���x=]u$�g�LF
�6Rz��_yN��3q��_fᾃ��"~�����>�7�����x��g�;�6=�?{z�����ߛT���`���Hhl��x�_1�U�]�}}x������BP����Ae��b���6�V���y(̈��z�h�|m7ً9ߜ�M(��c1��E��|��CE��y4��y�$�0®m��$���:O9���|.'_),g�=�y51�b2��C�1T�G7P��	��as�Ү.��>����B�Ʊݘ�O8�[;]�ǹ��-���-B���}oV��ug�L�} ���r�\Ur{
#��h|��������x�}��C��XX�^�=Q>"6��^]Q�Ϡ��3>�ѽsc]��Ys'/!j��BJ����Ш�V�NlLh,/�����/�E�^�=p������Ù;�+Y%�[l-�hTW��|MV� H�v�v��"���Я�6���R��-�r����~c���uK�1~�Ϻ�3G׋�o}$e.8u0�9$������r�����u+`�=o@�H1��_��#�21�ߞ�����^G��X~�0����3����ʟVש;�=z�U���,o��ڹH�����LۥNz���zE��Ĥ���9LZi����+��\k�t�u�ڵ�}fVw�{bw�^�Q�}Y���VȂ��S��yR�JV���t�9�-�n��N��[|�t�����xz�W��發����{�^��﨔��c;6~Q��ny�I�*+*��o}#^�*�K{��[R����M�<�<ߺ��߻��>�*TKL��'�O���ub��f�����~��͟_~Ck�Lз*MT�>ݝ���Cb],�G�@<�=�?���h��&@7�i��s�j*y�a�8�ۼg��uJ��s�%�^�Q-��]�/OÞ��z��"�EȦ�D<TɊRޛ�]�su�3��Èyg�p��k��]M"�K�G*�R��WV��P��)���'[�كb4�	�4�dJ2�.��끭�g���8�Ιs�b�O׉P��Q��@�ƆW��y�D��@�4�o
��q4y�,�;�T�kn%�0|S��ߥR�įC��5H�"z���#������[�ך�����A���xC�%����e>%����߾����(~j,C���GU�U�C{t�j	P�'(m�9B��^���P������ۡ�:(�>�Ï�N�n#g�wb
�JN�<y.�1��Q��`�"��uܡ����/�,�����X�̤l���W�F�Q��:V�a��i4U���i�]Y�=������n�35��q�Qݦ�u�kn೾���S����<��z̃N
���y�34�����ѧ4��q8Ų�w��M��ff��g��}Ǎe��2.,<N�o~ >�`�f�7� ��И�Mht��0V8�[o�e� 9r�1F:E���hD����ff���5��.�g ���զ�^w�n�u�^q�^�?4vq�vJ��ml�Bu��V�zq���l��pG��|�x��R�F:	P�kk֣�_� ���_��4[�~�2�I�N5'2-��|���O��2�����7&��7��.�oW�U/��H���W���V�Y��kUi	��Pր�o-�{�mk��S��#��W���yW"w��`�a|�+���_�Dp��Uzj$�6��2��f!����wmc���0���bW)��S:z�}4��s�:�L"��}��O�uEϚe���^�ʗe��8��9���͞]F)�gFy�ꊇ�y�����][�ڿ��rF�ݐ�y���B��NR���=��rT �\�KeS�� #6��/P�omR�/U��/�N��$�I^�暑U��(K�����
ac������J�Q�U�)��H��A�s�]�Y��^xmC���g���1-�j�`����>�ӽ���.r��󭤵�X�g9~�sڄ;��ч{9����f��X.�t�T��+U��ҮU���ǘ���c׃�ѳ�^�b�Ē����e&��sTCq5Y����������T)f%GY�C\�O����WO�^���쯟cʉJ��������0$�*Z(�Ί�/�1��n�"Ə�����;(��P���.��|k&�X���L�GY�S\j/�e)��	�qB��Z̠����[����3��=z]'� ��{�a�����뮜~5؃2���3%=���s�%>��#�6����rJݘ�������Ս}�}+u8m�V��3Pz���jSq|��at�m+\(~gw��nź���u�o��>��ӕ�ܫ��I����t�2�6��X(�d����	���0��,L��oi�gN㙂}c��ߠ��G�7�gJ�Nljz�J;������Ml�Q��M�ME��w�b��'��ƆWK�yP������,�m��7���&GC[�Ib�L?2�u۴F���I@z��T���g/@�@�@Ɣ<��M�\��ʞ*#s��n�SɊ�Wͭv�; n,�����qx���P���'|��������&��Zǃ�߫>�%W|�gwx�CC�#y��f�m�����ų`F�y�K;Ϸ"Z!��G�x�=,&[KS��QgK�;auf����Iikh7k���3���Ɓ<�6�������7�ԥB�	��Q�BٹC�e�)�r_t8V�ve���شV�R�łg_]�U�FUj}�vU��Vg[n2;Y�v�o}����� �=�%nj6q-�C�Ry��S��ջc���K���'~r�[4q0ISlQ�gN�hG���ּ�v����O���5����9JME��aۙ�M��=x�A��	1ѝ���5�dK��z�p��];	�eL4ɦ~^��4��¢�u)�ZBv�z�f�z�ss6�벉�Q�vJ�݌rY��-F|�p�o�FUʳǥ���2��*��/�������׏d
1�@�ZB��n3����z⡮Ɩ� ىx����29�i�����Ñ��-*ы@��A,l��S>k�F2;�wj�d���hhuY���Ec����4�gA�7�����}揯`&馫2��g�}��a@�GeΘ��ܑ�ܸ�8�.�L�\7�"_�{<Lp����������k.�_�w��	[�79C���.U���ċF%��.�Fv��Q�ܫpqf���5�oP�^���
��I�7�Y�Pނ��f�)?#GE�睡��iv[ ]�gj�����]��m�ʴ��[��SZ�J�&�݋(�V�i�-�����H�����R�.�j�3zn�̾e�@ʙ`���P�VD�ϩZ�L�&5���F:y�C^�!���0H���&����Aԉ�-^v�fk��ݲC�]��Է���sS9��L���ֿvIp4}���⇶Q ���h��~��o1���ʬ����Y_�M���=���5����~GއkŅ�dյ'U͟>�،?�յ��/85_��Y"5�p�f%Cu�#���ׯ>�~�l���rG�}5j�����.l1>�k��2g��īv��q��9:^���){�]LZ�{��vo�`,������=f����']��1��I�uߙ�E�����i��g�,*�����Z���A�^��yVY2a9Y�w�W8��ceʫ�	�B�(���4��M��/߷{�*�LY����H?b@I����iW S�Y�+�U�e��mO�1�a�e3��9��7T �bg�FE����ڗPdǶ�
�W���{����B;e�ӱT��PW���BNOY|�r�.�2�'�Ư�v�H^�uiCǷ`ݹҝ���Ԇ�k��g��c���]���W�Z89�o�8n-����H]N���,�p�s���(��&Ќ�=��r+M�\���~�n�9'*b��{�@KYDK�4q^h�����\�d���\�M�E_5���J�(�p�ؠӹcL�NmT��9�k�q���ݙk�z[7~�|5.���
F�U��Ͷ������������Bں��EGW�K3�F���=;{�e�Ui�lt�wy�9�	�Q��ޱѹ �lu���ɹe��/��[˳t2����F>D�^��l�66\�bc���ܷW_B�!��`f�ѡ����w��J'�w�q����S���� �v�{�ȦΉ}��;Ԥs5�����3��/!�v����g׵~Rd�%e�<��v��bK]F\LcX�1���+sd�;�[�h�|.�WO�r3ں@.oֹ��r2�c��skwk�o8�ff��N���P߇0��w���B����{��O�:i���f�D�6��dj6��T띴��0��
:�=ug���:����v�"V@sc�M���9�<Ȉ���B���v�}�zsݤ=~��1vr̹�V֚E�Xl��iX�iK�W4��;�·rcBK�>�f�鵳!X�\.ehb���zl���PMB:�'&wsx�������(v<O�>{�h��x��ET#˩��M��y�S��?��x��esj�_w+���)�G����P����Dd�S�5c4#M}�_�2�rzG�"�TIz^'����/���GL	���q	�R�fv�d�h�.K�s��Ci�mȎ=E��V�3����#��ӞEE�f��җk���*��o\�U�d";wkH9�M���*���=�UÒ.Q��59��`�;ݮ�ڜݣ��}��+�;Ur5Ob��K[�&�Ց0�'���}'&�0P7��E�����zO�rU�H�׌�_Kי���ռS��^�ܕÉ��U��E��Z�$L��y[Kw'܎*�f�p��]F=Y�O��U���a��|�s��]�^���8���O���]�1�͍Fg�5f���WG���8�� 2Θ}f(�� n#TJQ~���>k�S7T;X��_����n���Wу3(�����0����[K��	�Z�NK��o��4����Դ:yW���s.}f�<ܥ���{�����\��9ޥ>�-q�tT��1RXw�L��f^Ճ|�([?��y�-��+�ket�ѷ<���w�A�f�E�t�JR�ݙ���i��Ψ����k�O]!��ة��z3���c��M9%^���Bn�I���Ĕ�Gv�zA�۸��Lt����%�������.�z�.חd�.i[%�q����y���xǚ��-�2�L�ku��2������E��U�8��G��Xk�kU$y�,��R{"��&�� �Q�5�r��E��v�8�Զ��ڎ���F�I�z�ꁼy��jtVX�taW4�2)Q�y���x�ci#s�0w���k��h��\��nDVcfv^캗ײ��n�X|��H��?\cq❝�7OJ�1ܒxz_�dc![If�Nx��3��"P�ue���GmP�����#~�h�<�{d���n����7yr\J�tخ����NfK��7��=��A�x7�&JN�w����[f���7��5RmN� ����w[�[��Jۮ<p��/jv+�c'����$�U2�j��K9�L3�S�(;�����luҰ�BwM�\�b�d�t£�]C��.���GsI)ߥЋh�k{B�\�u���\/e�T��Y��N�t)-��H�������N��^��Z����dwN��De�^�W�x��**h�{�.��k;�I�L�q�yy��7��d�C������'$U�X��D�"P�1���l�^Ș)xw���Ƿ<������� .}��A��~Zl^
��h����^��ň�{@��Ln�`�Ӳq���5�(�MukJ}�S{w7ݲ`������8m�Y�6{oT}QKhE	��`�D��;L�,U�ۘq愕�XS*J���L�y�����Q��5�e��e�;M�����g�߽�ۓp2�O}������~]��=���16��Ɛ�#�nl����m�^��
���^��y����	�hy�Q��U�ұ���=���x��o�w2��͑�I~o.�f����\���8���Gg+��|=�׌͝\pzy��K�|�uݢN:k�<]��θ�����j�C�������k�T����Nܛ�H�/��+��pi��`L�u>2b2�F�p���j𞏺u�ljw�� �$�5B|C�(��9�{�0��
t4#�ɛ{ۅC�]�/�2�7����v��SYع�
���U:ȩ#eE��xK��%͡wOk���V�ݫ�������7��a�#�p|˃&ӹJ�-�uq���ߚ�#��<�Y/yw�=>��t��У��Mvu�M�̰��Y��+e�%(�쮲��;F��k1M�L6��=3�&���s=���m���k�h���\r��"P��e4{���(j�1D��6G$�&��W���]���ڙ�[YUUQ�F**��"��-�)Qb%�t�O'���`��+E��$U�U�\�Z��QZ��U��F �ҫaf�O'���|J*���p�AO��F�U""�J"V�)W�֨���#��<�O���T���A��(�O-��U��E�mDE��DU�"�R�UEA�O'����Uc��m�e-F"5J�chVڨ�++U�"�����
k��m�E�AU̢������։|��T�� Ԣ#R����Tk~%U�D����Z��((���ը6�J�X"2�"�.��R,UR�i���V���[hV#-9�1���X ��F�+�W�AU��	Z
��KJ�n�fIU�b��'j((�"�Qj[Ev����1C#eT�^n�`#�R(��T��re`�)�ъ*F<�	 AK��R@�NmԺ�W`��2���O���Qw��ţ�,aU
�;�ɻt�d�	�a����������}C�g2����U����g�xH���"�xf��m�y�V�!G��;���eY�IV�y����m,�i���|��V����@lJ`m�9hMl��������{p�U����K�%�{a��2�k��ӊvF��i�#<�5T���*K�����W�=�G��2�R�F�0���lsMؖǺ��L�m=����hǁ���S�=�/w�ux��� r��hg�a�k5�d�U����:��ELqS�7W�/3)�4���W-�;�R�^�n�we�$�4�e#e��|��~�����S�~����4���ŧ�S�����oի�Q�5[#��b&����7*���\`qk�6���>=m�.��V���`)�����VeW��=��]�j��wvG�:�>��k�~=��Rm�5��nV�$�)[f/7j�,ǯ,��ھ��x�>�37EE5��́-�����[ȋ	��A�-�].�ʯ<�
��� &��u�`��q��M%�/��g^5/'-��~j��UI�^�	c۞��S[�l畋��ESw:��К�ْ��S��y�]P�w�uɴ��ˋ����Y�����7�/v~��KE�b��bJ}�-��**��J�E+�yk~�N#�f龭��R��C�Y5�=}��i��6���G��/)SRǣ2��f�z!��3q��oRiΧ�� � G�S���s�<��ptjg��/���L��e��3g8���P�;�U���3�ΆX]��!9ո绽Bɛ�����W�8߽�3֓z`	?,���	f��͟l0t5���q�?���߼�/zt���\�%�loVz��yҤ򉝒E�{5���xX�9	�s*�{:e���z���ռ�j�'�|o_'�ӝ���曬��ว�x�ӏ���1��� ٛ�طz��}�R��ǯ��s	S�Vǻ�>sA��nc��k��U��c����h��p�6��\�g��W�zU��R6�`�z���B��:��Uu��U���~%�{:�~�N�7�����HF{2�z�[Zu�͇�<xWת��[��o`�z��7M,'G#�
����x��i�D�X�,�d�K�z����p@)�R�ڌ��5n��[�kQ"#��|���+Gܛ�͡�yS�q�ֽ�>6��?�l�P��̓�߽=�~�w����O�V̌���y���Go�VZq�d�P���+K��Q�g66kPO>�HJ;�Z����<_SY���aJ]�mVc7j�5��U�vTL�e^�U�9�\�~�����ݫ\��`�d�w���UÖ�a�q�Zޑ�2��Զ�q�*��f���T,��a��V�M�:/no��;�Zi�2Jh�2=���j�t%��NKv��YYëE�M�㷴.֣\�t�kq�5Ϡ��/���+�� ���^f{o�lH�����/�t�"z��V퀖����Q����ϐ�l���<:]�˽�1���ͱ��F�6_v����j�ϸQ��Am�8�x��גa1v���mʓ^��陂��đ���۵����JA[�o�@�%����zf��b/b��&Bs1vx�H����Ϣ
1�6��w"�o:>W�tO_1$݉^ix�~]�w���?]C��E�T-x��yy��|�[x�xA{!��䮆�:�����Ud�VҚ��uy��ܫ��o���y���N��^#�]�u�6�Y��;Ƥ�^�3�}���,h;�q����\G'3�õ�����������s���܍;��ub���":)e�����׵L�v���1�y�&
{+��\�ζb�f��;�:_��;�͟�mC{�TU`7X# �2O2�`$.��X��fzfi!�����Q�؇Xk�'��Dr�Q���ͅ�;/{�=��a�X��{a�7ې�1�.��<y�x��8�*S-���Gmc]C6ƫ]�X�&�t�Ҫ�=���-�ˆN�9CV3Kc�s��=55��fu��O[d���9�^��~�B��X�a
�#�������.z��?6l����y��R�OC<����?�st5R*�G���?d�����w��:	6/>�R~(�Gj���&}Wl��Hk�WŭHc,U}v'2�.�|;�ݛ?G�zUbV[��دiUXF�����"͑7(�SP��hŝ�S�ϱ*���[䧮�{�bF/^Y�.�����>쩚�oP�s�e1�9��DέC����A۴��g��tJ���]���A<��,�|.n�b��HY�/h�d�#5KU�︁ҙ�|�u��!�n�}2Y�vb&����6u�c�G�	İW|Ե}���?PFN풺i�񛷞���]�T�n��ν<6����#�E�K@����)4,ջ���a֞lAw�/٧Uws1�S�q�̥��pc�<g�Gu-VQ%C6�"��y��]Ӷ��f�fݥ��F�l� 7gL>ù]S� n#T	J;5��;��m��5��i�=�"xbv�`@��z �侯H<����l�픂[����C�M�r���q��ŧ���[�*�b�8��v�'y�4�ݭ�s$liD�1%���=!�t��7^�$��{��Q���n醋��8�(���ټ�͝ہ8�fzL�p�k����k͵Wy��K.x���hNB�tf&����mx8�u*h�����:���mؘ�l�mV�H�T�&������f�
��¸���@w��^ҝ����iu���p��A�/�7��We\x:t��T�~좆v�mږ�"�UIϦ]����Q$�Q�4+d����>˼k���][��a��k�~��3�K���'(����3�e+^�#NM[��*���P���3Gu2���!��H�t]��(e.�M�R۸滵�����h*��oV�-�x�j���Ǜ�K�֦R�Y���%S_l�gW�� ��j�펾�R��	��
̪q�=Ah��=����;�_�;������k��7�w�-������샷i+���*�|e�oF!�1a�u�����e��[���l�v�c��U.�J�������N�Yp�}�'�{���Y�+�Z�3��ܕ��].E݌�LZ�l�:0�dJ^H�J�a��r�-�6����k��U.S3r��۴;������+ܶ�n�	u���v,2!���yN�Ij���]������\����KUy.�V���!�q6l��e�/~m_�XO�!�y�m��RH�a_�g��MrTM�i���h�m̂�'����%�G���,=�}l��Ցw��=��]��KL�
�9���8��b(�H
���FГ�/�n�Ul���7	ڕ}/.��M9�-H��S��Ճ���3�pU�g������@Q7���f�q�𳫰�lE����u)�E��y�ȃ%�)�E�.�^mݟ�W3r��u��z�޾9�$c�ƨ�ԓ��r��j�z��4���-�ǔ�F0f6�<���{-������5���M����s߭m_���!�o�WLr*�a��-[(mL���֧��Xsz�wn�	tv�"��R�!����jX]V`ϳ������p�D�t��d�������/����IDd�!d�lЍ2��̣�,��
�(����c�����ys�|*�^����R���R���C~���o3��;��6u�_:b�c���z�U�Rv�W9@��v�US`�2���w��6�ɻ���K'i��f�xtB��j]f4;���C&c':u���/��o���Mn�V�LsC4�~ST���e��~���,�̊�5���rj_�I�f�� Q���s�8֧k�B����no5�G����KFJ�cZ�1^;��r�넭�!6�Sy<YM�+6�6�<YY���W���hU�2����r�R�Gx[k�*v�dܞq����ؼ�>^�c���wT�����ڂ㙸�x�iOd:<��f3��83 3N����!9+;�]�[�V�v�y�܊W�R�lv�\��0ޕ���}�����}�<�I$�o����;�1*��]>א6yN��7&]�����]��o��G(��>�Yo�/{Y��>c��\lm�E���t�A]��|�Z�m�E��'%����/7/H�r�G���ST��>F�7t���Y@,�2��(��)M��m�c�V���g�`|���z������*E��ٟT�|ݝ��*�q	k��N�-�{Ly��� 8U�w�#�u�Nf�Ev�m���w1�0>��k�Z ��k�l�c!������>��@�ig���a�Lj�e�5�/Ÿ��^Ρ^����T��Н]]�ٲU��D�������z'�Š;�����7�l�����dX�U��;^tS�ݗ�]��ۙ�:e��-c�[	Ț7W}�^ky�:~�0�8Q|��w��ۓ���
��7ږ�ֵ{�&p��W�0
�JןS�GWuޞ�6 �Th�[}�%��OS�Ax�ގ����g^�=�z!�&�����þ{��������Y<67�m������ᇞ��-oeK��ռ{��n��O�;��c~��1�����}/�@dj@{51�S[@$�m�����q]I���7��Q�;�PW�o��⣶σ���<ܺ@x�RQqςt��6@�M/sY�N����Q<��갳'�wU������u�v�Z�ˆ�$���g�+'hގ�'��\l�k��sثdR�F��U��w���f���˶�q�/6gz�p�C��"�O.��-�Uz�Ww%�+�+�k1�Y��U���ܖ���=��!� :\������Z��D������rX��u��20�qg�;qu��ם�)�hӒ9�v|����=�*$G�Y�ҵp=�뙧����?^Dm/9�&fk�\�٬3��@w+�{cqj|z\Z"m���ά#��$�[��W�D��3��^��}��͉����]���w�K2�*\�ܳ�eP�K�"�����r�5������Y�e��0��?3r��/�e�72���]��SW70z����ĝ6�T˵��Ӂ}��K�������m)�r�*�O�-�Ik��k\C���f�%Xp�������A�.x{��t\������� ����~+ƛ��������gw;%���@Pr}�Z�&�N�I<�0fHn�im;���<X�(��n�WH�O׏sr���F���������ӍV��yg����[�Y���ZQ��H����D�^ۧ!>�p�b����s�;���fv�,���׫��R�� �I�i����-]��@"&�оqwr�6)4vC5�N���Q[�2$l�.1S4�R6cφ�2	���F�T��&�e��s�wdϫx%,I\��YL�햣>{��U�Zi�7����B˱;���Q���,�ޅ��.�-����V+����'c��;�H�~{�7���k�RPu��'��F�q��)u�iw�����?��zԟ�������ZN��ჳ�T�a�-R!���n6#�_�!*RT5����͝�ُ�4o�+���:��t�4y�,�V�����0��UmL\ہN��⬔w��0�24�ś��8_��#B]=Z�U!e�oiN���)e�:�t뻦��4�hF��j{�*�Z�Υa�2�p�Ǐ��?W
�\�5��.���T-Qz���i7>�2k�>���\��q�y���;���[�;�#��4�Q��-����ܜ9�=&���QV�f�ʇALG���ǂ�i^�%�w&x��3_x{n�ۭ��(}=1�����z�#�N�8>���I�_��f�s��	>p���G Z�x��p���[J卫;Sc����'�)n=��<{7O<�F�;�^��A[s��FQ��+����Nc2�0�L�=�����Rr�Ja���;�jwfj�[s�\#E��".�\H�D;B��YAے�m�"Z�M��幄��T�i���]������zrb8[��}��V��ǫ����)P����uQ��U�wRs6p����]�	�P�]�'I`9������U+ڲL[
�t��Θ}<d2 w�۫�T=^��7p��=����kK���_%�xq���yV1F3{T�jE]fn��IWgy��{/��h��XU�T�5�t�t�)�����Ww8�+h)�Y���c��+��; ܙle/{V��+%�Dm1�I]����P��:�`Ϧh�y���{w��x��M}��P��-�p����S]�U/�D�s_�1�J�n�o�:��o����Ƿ;�w�5G�d@��=tE��uA�i��|QݶN�h,�:���rT����aC]G��!5U�����%�� ����R�5Y�2��(��/�&%ڨ���΋���m�Z��eN��AjqX ٴ��\m5�*FJ����g�rH-�H���͗�����krt%�O��ս��<�����F]�q9]R�G�[���gX�t]����wpw��Tt�
�;�Α��V7�doA#������=���cV%i�9��2�Q�/a"�򫚦�z�K3���ܭ��gs�|�>n�/��Q1���9w�{tJ��ڼw�0��>�ўu0۹�)=�����*����2�L�5�"wְ����i����<٤�D�z���3\7��a
�{��+Wٹ~�nD��Т�ZY}�L����ч*U�U�gZ7��,�X�+8
�<TDkZZy�b�ز�����@�*bNo"L�4Na�o.0t�WUwNB�KC&]r�
W���+���vh%˷F��h����"�|Y�K�e�Q�(b8�x��	�����r�Tuے�%٘Ŷ.�`nc��E�;�^�q�٤� ������0U�,�K�X�Yf�B$e�Nӭ;QŻn��A���ㆮ�٪2�u�����̛���%"��pY�$�&��F�� �}F��uV]
1eJ,V�J�}J�"
9�T`�hQ)��*�*���:�:~'�<�'�+���Q|j"��^h�J�T��X�ZT�j�+)iF"
*Y����y<�U"�|�cR�Ԩ�<e�]M\aUT�0ҫmUQ��0X�*�i��y>O��J4jPL�V�
��D�ʜ1�D�+Q͏0�UK�5�����t�<��(���[Nj>5yцAM�0��֓�DVڍR�kET�X���Qv��R�VQVTR�6�DR�S/]��6�mk�J�39QUy���R�5DSj(��U�e�Q��5S2�Tݰ�6ŋvq�*ۮ���+x)Z��YV�9�J1�����3[hE͈��S����N��L:��e�*�W5(��XTۓv�2S9ŴUU���է[&h�f�MKlDÒ�ˬȃmu
��g���P��)5�s(<^��e"�y(�h�V
*��hUee�K�)֪*��0��ߏ�xlmgJ��A���,�Zh6���ν���,*�2�����&��ܵ}�g��29N�Ĳ{���)!�ih�M�_{ת���P�m���MJj������m^١D��rb�U�R�KsRޣ��^�Qkyf�s۝ɫ�m-Z���
�%2�#[����VwIK:�o@=Z���8lN����{���b ��?��'��%�|�	�:3'ī���6�2�0��o��`$(x�;��U���n����^�I���ZP��w,�:�C\�M�!�Lƶ=*˗�z��&����W��$�պ��9q�,9�M'��$ShVѰ�5MLVv�M綏�XE��/�s�+_N���`��{q�[�ۡ�6.&�:��4�ڂ��an��фϠ,3ᙆ}�c�8�Kj��w��ʔz�;�X�v�b��fX�l���a�3�U���`�>����r8S7p�}�������]���*R�)�sⲁ�M��L�*Wd��txK���������mV}��wi�iM �HW�[4ye p�x�ǰ�5I���E�`��ْ���z&�vb��[���Dm'�P�`}�U�����S"��D(���[��}]hWp��x��^Q���|EȨ��g�i$O�o����iy�L����z���n���b��8����D��6��w9*}e���o��R�H�T���5{&�!�h�q|�oK�e'Y!�Ż+4�eo"ᱹ%�}C�6jSV'Q��R���
�`섮L]w�iu+�	��9Ƿ��gl��YO~=��7pT�i�� �[�n�9#'��� �љS�ó7��J��%5��ePr��)� t�]BB��+ԧ���OV�hu��Q�޾�>g'+ĝ5f�@�kQ�s�:��S\�!it��v�Ȱ�wMg���!�m����TJh�ו��U��x-�k��-�����st��ss�<�J�k�^�ޕ��]%�:j5�1�ǚ�b�z�w�{>;��+w�3�fA�W���4q�r����9�L�����X��c�Qq��CJ�95E��ek&ٜ[��G��q����u�^�܊�y�'�vW����܇Y���z�y���[����p�(2]b;��J��)�F8ڗ�9Ow@4��7]����"�2����q�G6A�vD�:��8df��V��qZ��.}�L�����`�B��|R��FR��a�2�)�7��/lG><"0�<�36�����߮�ܿ�-L:�-jl����r�1yL�M&�=|Lš9��zl�٧���_x����.��,��7��Ϝ���o2n�Z��.��95R�� �I�
��(�Kwi̓fCdp����OZa��X.|��6a��|P/#�+#�/T�n�_p��a2�:����i�OJ���B��)Z߯4g�����R߭q��r�$���P��xL.'��n�fkgg/F\�y֦�g��ґ]m��a�N���Dc��a�-fOFU�;Bo�Y�C<#���<��5�s����Rt�����[/.���U8�bwf��?]��StUKq�=�� 5P����QRZs�ި�Q��P���t�_���Q����#~���;��6C���p���1�5�w&�q���v�?}V����~Z��v�R&�+��ݼ#Z�V�K���\.Zr��3!�j"h�C(��c0{l���&Q��t@��dחZ9^��a��h1��:ӛ��/�!�`��%���u��Z=��Q4���V��e2q����ce��
i�h9���ي0�u�Xy�����y��;�|���LW���i�^�	v=wc��nς���󽩫�R�r�P�3�#����7�d��+��cs<�ޙ���kVي�툖^MU�c!H(��O��s�I���mJϭ�߯>�lr��Y���2-_f�����Ԟ��Nq����#��W˻�+�Y��Y�!�<�WGlS�e+3+Y�g��^�/�ےs;4.^�I؜�~�N��	�6ϸf�	m�[ڎ[JJy�.��l��|1s��:��K��m1�ޭ�m��-�Sͱ�S�t!�5z�t�������z6km"N�<�ǏM[�q�^=N�HC�^_���0xͬ�o�h���!R�������Fm�M���>�3���&��x{�p	��~Ŀ�������U��ٛT��;z�_zmx���Q�Q�.����j�I_��Pjߢ�Sҽ}���j[;��.yweH��!q�
f=,��-�����)ysz�s6mw$VV����R�:�s��s�)m%s��X��MU�H�m���~ϠX�L;2��"��]�\jx"C�'�k�kW��v�bަ���G`MkÆλgi]')ޙ�/56��1��!�<f�_��TB{��qך�����S�Z�����S����wR�{Z�),}�d.	���}��;H���j��8�7}�����B��PX�YA}wV���SN'��ٗ��!�Z,2O�Oy}=7���߰������R(9@���fJ�g_U�Z2�g.nnĸ��nκ[�F�j<ʮC�5�b�u
�L��oz��a��v`U䋞�n9�I��x��Y�}�l��=.��~JVS��HsJ����O��XI��]����ǟr��8��9M�,�Z��b�5ST��&�³��^o_$� �N+	wH)gP����gd0[���T��mcW��z�����S�L<�+�2�5�|�Uv�88m��,3t��ڰ���罉�qg;����S��cm���W�]��!s��D�4�pq�1F;2���@����n�}�"gu����#`�4�N͙}\�ʡ�33���4m`�v`��o����w��dfRm;���{ӿw���;΋����J<�շ��/1��d@Xn�Ŭ��6�/�uۚey��ہt}�����t�o3+�Uw�"�2N�{;�V���ؙug��Ԩ��x��6���{^;%���k(���;��jO/���Cx��{S+�{�N��G�Ъ뛲����gW,��u*:{�n-*D�j����{�y�'�C�����l�^l�3+��V5o\p/����7p�@vvO��� s�kČ�Ke;�|����^:�feYA��4�Ð�Y���3%�Qb�YB©��\8Rّ��k���~�}]ս��T�)72"�u�{��$2
����\O0����_M��/��,�k�zpze��Z��M�R�rWCר^�'rbޝ�nZ��77֥��m�n�Ԓrg���ڙt���Ϙ��h��+Zs��'��8�{'�����	�2+H�U�
̪+[-�.�k�5p�c�d����\�U����]��1���
Ԏ�z�dѵ�ݾ wjZ�
k�CDF8�	/;���Nk
�+�]��g�ڊ6�ݴ�WV?R�ݙ�R�`���+(�� ��5�O���:����ޅĲ'WF��m��p��t3b�NL�2�7=Ε�~��C�1F�z,8U�����Z�W-2N�[�MgJo)m�3�n�-�,5z�/�,c���gE�rF�:����XFp��o7,��Z�ص}�ƞǐ� u�O���b���&fY���+	��o����4�.K�������]����_�z}�0yyP���S���f��RV�17l��3����;
����q�#a�sf���u�j��%��ǡ[V��f`X�{_;xf��w*=�Y�{>�4	����e�"#Y(d5:hx�;�]�i�ah2v�k��:���}ud�w{N8���3c�br���\��D�y��X�i} ���-c�Nנِ�C�co^~�&ٚ-��6i5]6לz!�0E
1�����_}��͈�&�yS�|򭞂6%�Wgktsn/=�c��j�|�`�v�3;�׹���X�r���wXF��w��W�e�;A�Mr3'�#�������~B����O藟���̴A�C�ً�v�r���4�:be���C���+�$˲1n������b���j�����<Ay����8���g��� K�Ͽz�T��׈����� �<�s�;E[P#�i0D/��v_����Rg�w�Y�?Y���gf��r"��I�~d c�_�r��� ���MK�"�IS�����#���ʽ�O�TbovӞ;�l���F[��5��'g.���ӊ�g����<1v��wR\B�]^��UT�sP�e����L�uD�S��{j�Z�̈l�K١���t��XJ]�l���5Nء3��=��:[�33[�M���8�z�q\Zj=^n���%K��Ie6��g�ʜ�9�*��N�S��q�ළ��ۼ���E �s%'���gWFN�k8��ޮ���HL�۔���Ljެ�֟[��Ÿ�,M<����<��Qw�V��3��gH��ܮ3˺Fq�v�KV�/���u]�K��'v��#�6���;o1���+�l���V��f����w�E䈍����w-W���|���3�x�������Ŏ~���k��F��V u����ۍ�}>}c�A2�٫�ۃ�b��ſE�4�k�k�0�f| +3��7�?f����R�+����<�/�a�ua�v�q�F�j�`��v�Q��'ۏ+���*�fF�������|�!ާ{s��X����X%=�JV���w�|L���(^v��*��*�uف$�<��ǣ�g�M�&�DY��^��K�kl.d-�we!�Z5����pㄋ���nD�06���A� ���?��X5��[�ؗ�B��Vz��{7u���Q���)��힩�4�|�wƓH�)�m����?��MY�R)ߡߴ2|�@�ۆ��^s(�R#���*f�C���<VP?E���s<�5��s{�*#Wm�����М��ʣ�a����
Z���۽L��kSeP����o� 6�.��/Q}cL,�����M���[D۸�����p���)q��rA�UL��&��J���q�ЗW���)�^*g��㛓j�/*4�/Fwk�6O�L�{�Lr[^�&��wo��_�mŌ��n�ӽ�;nq 0�$�Sq�Ur;{1��g��r��Y"�g�,݇PjП�����U�.عE:�EV�������=���lnW��/��j�hgb(��v�"���qV�(y��ekϧ�z	[�Ĝ�����z��w��l}�Yt��2��Ql8�ѽL)x	��ȭ=��S�B��y��:=�ALkh;���|9�NƉk���'�#tR�c(�ɯ��X��B�o��)i؋ �J8FN�T��ޥ�>�]�%�ZSGwU�ʺΜC �����X�,�х�=[�R�ޡ1�6�ν��)�%�r���!��%��`λDA���8�m���o,c�"-*;��=Ε��cƕG>�͸���5�����tp���i��4s8L���7
��5����A΅
s�Z��+��h��h%��������aawTb3a�K�{�c�ݼ�Wluf���o��G-�mt�2 l6t������4��)yg���M���8,���q������)c,��<ezo
Z�8u��}̘y󿨼�3�8��K�n(���e�i�:u���/ٝ�{عc��s7����~����t������¼`��(�OW(��a���}ޒ�#l�|���&�=�\i�Q1�,�@��W$KD�f�u�܍;�˪2Gq��i)�p{���~*=�E��qF��(w��#mN3�Uj�Řo�4�d(��yn��6|����S1Vx�|p�}\�q��5���y��p%�Iq^�K��0^�QJ�{1,��:���\�l4�,�ݝ����z
�-��LFЭ�e��:lR�����Ċvrmr^�?(�����^i�yx�UvÇ�=�'�>�l�:/��/AP�&#��G����b^܏��3p��]j�?<=#G%<�fF��c~8J�ݺ�G��P�%�\�殍��Μf�7��� a�v5���yo;9��Ô��ݽ=�\���]�0q�"�o���It}�wCIն�u�����C0�����-q����ƫZ���]^�b³���B��7���*�,֜}����F�ʥ,^t�j����߱nQv_y�K�XrofuҌ�4w`�
 1:�q�Du|9@�p;n?��#���<+�Viܱk͓�^^6�[�}�)��1��:���L�2AbQCC�����CWA�j�YPT�������B�i�GcT��/��+�\��u��k�=(2b���I�j��s�Vm��R�\* �!Mr��vF���K^��k�o���Mla�N����\/�؃�M��ؖ��Ǆ>��])dBû�$��1�����;t\cL*�b���&�ǂ��p:=�Bӧ[����;3�{�66h�w3<,�P�_8ў�������5����ps2�̔aU���6����/~�X��f���n���P�9��|rL� Y$Ҟ(!���,��^b��k��@Dy�������kOv!����U9����tt����3xd7v�D��{�z	Ť���*���LϙK���������;x�z���dg}]w^��YƧu��pȥVL<+�9M�B�[��CB2���E�=7,7b�qu�j���a�e��LdC�\kϙ��v^pd���"�de���f�X)ܬ$�۾���Ŏ�vl�3!(N����[2�[�un��H�N�u<b\�;�c�q��t,�A��,K��p�ݾ�'1�J�U 	9��f���1��N�u�)k��m]''*�3rM�.f�<�L�M�w��37'�7)V1
�1�t�˹zw�xL\㭫�2��3��fй�ֽJ�#�7��Z��}y���0�>��~~�{��DT����OP��g�9�L�6�t]���R����vѣ�!�D�� �[�dɭa�~R�`+��U���Q�
-|��q��w"��S�뻺x����]�x�&�֞��s�i�8|���]�:��^\���i�k�`��UNY���v����8��z�q�� �LC��ԗ�i=A�5*�2��G���gx�-�3�W.vG�����VU���Y��fi|���ѭ��aw�z�H���䆑�)���.I!���X�,��֥��ܨǹ�c���7Kk��ǫv�D�NV��cZ��=����y�3���)ɶn�j" ��#B��J�gJ���v�[E�8��ԾR�=�J�[��t�y>O'�Z�Q��G�WY��T�v[\ʈ3D������9;R���9�Z�:y<�>O"��ys"��:�δ�h��W++���6��`�mڶTU�kR���<�O'�ȃ�x���S�~Y��j|ݥJ��d�*��b�atmF� �����Ko[��K��.�#-(���b�++�YZ�r��UNK�:���cT<�C�uڱm��b���֕E-�j�3p����QmX�(1�ih����T��n�9Ѵ��3]3y+��u7:.*�v�"�.�=j�e����b�����2|V��G�5��;�ݭ2੆��B�aX��������Q3X�ErWP���7K*ڈ�e:ţ�|�JDŮ�l�(�ʍ����Ka�m(�f�m��D(���qJDk*�nZ�EQ�hW#�{�r�]k6��ckF�_o���?�z�H����3z*kdl�]�J��vX4�.�al��ʔ���m ���X�{\�rԗ��\�I��;����������z���3��_Ux�x�e��Ms6��V�������u�5�������K,{
p�����[Al�P=�-�m��a����������dខd>�]M�R�R�m-�+�*:�	�X��u��~v�wօrwZ��4��.F�
w4m�*�d�=�"��M.-��j���oG�
�f����Y��sΉ�\l��P�&$�����j̿E?�j�9�#h�Q|%�{�5�fׄ-�(ק�z�4�C�F��xln�S3�����)G���ݺ'��l�^���i�������{y��v|�����c���;�	�k;#D��4���y�;o0�j{��d�K���</��C�8�7h�i��;��h��j�c���b�V�9v�Y������Q1»�>�F�hQ87wn���ƅ�>��#"���^u̚�/ݙ���B�O�z�xf��@N��z�]C.�q��������F��wun��׳��덜Y}1�qv+�<i���������!�fG�e4k�-QR��M�ǏI�9��j�XČY�}>��n���Y��鹽����_c��P�d>�O1E�dD�*�����r��OҼ{�=�s�Â~�:P�[DCrXަoj��Yk*�k��s{#w���Y�d�hHܟ�98),�n��~�#U�G�S@0�e�@b���Ϻ{sd�����3��:�h�&v�u��~!=x�B5=XqU���&��5P9ۺ{gY��k������=��F� U�N��jIPY+l�璻�s��v�l�]�r��]X��#t�̐<����Q��q�5�����+��Y�F�ip��7�����7z����T��jl�+fȮ-Y��[9H�_��[�7i�m�����oDm�^K0�M��S8q/�d��o<���wυ��SФu�$�vgsOa~��y�<�^�=���<� 6OK?3,}[ݐL���DCB�:<��2X�uos�{6�����:�|u��HC:l�$f��c���k_At���,wGE�[R�d�O;"�B�`�����i4*B&�Z��J-F��5�g`@n�-9��|f9�΋�=�r�j�Jzs�y�i+I���a�S(���Jՙ���pu���'-X���׳MUK���ȠK+꧕��pā��K�0f�vgv{m�%tx�5D���'ue�c؅6ϸf�n�2�l��3S]���L�ӊb;�D|��;���/r���j��J_�W�q`������~6�=t@ykO�r�}73� l���g|Nу�����%����8o��d'��w�Z��Ǥ6�&�!Ƃd>�פ#�i��1؞���M���\�RܿJ\\7I�/�5�7��.���<ȼXg�eM���Ú&	���̦�8Y�9��e5�m�����<��"KI͵��N�����ӛ���&o�]�ǳ1\�����Lǥ��|}�2���d�m�fN4U���z�+HO$����PՍ�~]aӨk9d���A�Hz3�%���/i:��Zצ�����P�y��kb0RU:�$6�������"\�u�8�7`5/\�z���i8��F�q�wO��6��>{��C$��%7Z��DƈG�5�h�'s�y�~<z퀍(��Ww���+/}�]��s��jM�M�)��8Gw�U%�����~]¿	�M횁�0��ٺ�sK����k"o�[)�F=�f���:�Xn6��g�x8\
���2�-9M��W������E\�|2�C��mg���Ӕg�S�]��+}�����W�7�]�Np����v�8���h~l��t7���s��r�����7I4ܸט�ėox��P��'���.Nu��/՜6厷����O}��W�=�}��e��,'�︫����u\X�&��11G�6]�0��D�kӳ�f�th�*%ܲ���Ȃ.��^�C�M��S.�<f#R����޻�����ƍ�w�1�%5��+wu��5�ٙ��	��ɲE5�f�e�hd���+_N�6�v*i��4Q��mݛ�B����:o�Cnx���̻�1
*L]��#.o�_y����^��:����I2�2�!��6t�� 2a�-�$8�/�>�w�0�����:�=��'\�W��V��,�^�:w�WS�Mkzf�b3&vpC�ZT����I���>�'"$��BƣӫF;��˫A��CM65�z���X�Άp�|Kµ��;��s�ծ�QT���!'98��������X��2������������x�w��I�t:���r僯��{g��w��(V���=#3%�o&�O�#$j���.5�^���ɟW���|�ZtO�*���g�4����Vko��䔆Xy��#�M��bv�8�n̟l�����̊
���Nz�V�yݗW�8Ov>�6z��ЯZD�i*��t��wj��r%�ڰn5�Oլ6O�#����2v��[@�ʠV<e�(�.$�W��*YO�(�~�f"(M�yX����	m�#�fo=�6��ûY�#.v��m��(��4sxu�d�ۂ�q\f��JV�V턶%u�7KL���m��l�<ם��y!�d� �*
�h����uǀ.��
ؤ��ꅑU�/^�+0��o�.�vtÞ�\m�h:wfM�z6������$�����͍qG'������5�e�0��(�(Ss�α�Y���	�w�Wg�<a��ˏ������.txx���i�3�yc��¶��}��q"M�m-���������\Dw
ˊW��������{S�ەǜǥ��5rn���5��ze#a��}�*ŧ�m^����{�]�)R1a�;��x�w�Τ+ݺ ��8���{z�6���g��s׌����Ӝ�e{�����{�^��X��њ$��4�A���PM�MUvv�͵Z��a\ud�'�qcV}��Mݧ��:�C�4�Mt 9���62��1N���q��y���	��- c_�ީa0�;xj�6���/hl6�}�aY���X1�.�ٛͽQN�[F4�=ʹV_$ِ(�Џ�:�S>
<�O�M��Y�kuY�;����F�o;���CH�*j�`����d9������vg`(MO�r�(k?_\Gwtt�b������'�H�Su�R�g��}5R���+hDF���e�$�-R/�=p`Vl��)u�UZ̐U�Q�eW]�.q���*_�L�,�"��%�q��Z�"R�/�ۮ��)co٤�^�>[��#j,�v��%(�Y����5Ά%0�Ҥsk�\�#DT��şj��Ŝd�/�R��՝f2����\�h�UB�M/�fG1��oH��E��s��LO5@m��{=�o���wfG�ZtG7J���㾉k��x���|��"=�w/w�w�|``H�& �Dɬ�zf*��L7��XVϬ�|Z}����
H��|�a��e����w"��l�^ f����R��8.�OD�`��P��꨺=����h�$���H�*S���9>g���ս��n���P�|~zi�<E׭'�עF�/^+zA]�[.��g�hv��:�@�Y�.�5)�{�Os��]ׄ��6󍔞��^9�׺��01
m�|��b��~5,U�4\z�^���?��Ɉ͑c�S���Z���m��;o�<���F�N�"��}vE�6:N m�ܨr�}�h�'-���^T������4���m���{"�@n���d�"�f�+6/��C�72y�7�t�ҬI���pHF̱�Ѯ����x�,/eKKJ�U�'�1����1� M�n�^/�;��T�Q�[��w̆P�f`�k��þ�\��>�䖩Zf�?��3��+��[����
Vv�L�s}�<���S`�e��2�������p�#�3�\�;)�YOe�oOv=��K�|ONz7�V��N�g�����i}�fE�έH��j�6����[�OF�&w��Q�9��"o�M�͌�Hk�2�=Qחg=wr���F/r�Y�K,��D��*gr�:�]u���"y��Fg�����V��IGhs���#3⛉&����1�4�{g�������׀U�{�+�Mz���>d��z�&#s�cNm�C�ev�>P;T:��SZW�XdlGY9�QsQ�9��ܝ��'���n��ّC)�O���p	n��5���	Tٰ�K�u���⬪]���]��ןq��{��x偛�!�ؚ�oZ�ξt���Zilz�4�7.8�N.]�
7�y�e٭Ia�7�/�(��~�C���i�����n�m��P�Zz�.z��'$�È��>Mb�5��Cdǘ�;j�w�Ll�UV�$u�	.�^x��vgE\C�'w�;{�f��!������;w@s�b5*�����P�_gT=���+ A�rx��{��/��IZ��.ӊ��6�乖n�����F�{!��~8�=����}���Y^���:�Lb��
�woN,j��(;�i9-����[�ᴚK�fI&a��]�J���UoR�s	!�L���}�3m蒞����"�}���Ӄx��ގBH��O��dj��Oe_�݋W��#���c�� wPn���aawW�Ɍ��~�,��n�߈!���ݿ-=���,���	��@n�^sCa��8����lLV8�}�w�{e����E�}���卲�I0%JCe4h�Qb#� �#+ހ�����Y$�	Zw���˞ ���B�fd>� ����H��I.�ڨ�G�6��4�#l<`�5�az��E�N�{����0�R�1q�h�w5���g۶��D�<��/Nڦ@z��[Mz=sA��t6S�ۡWwwNU�8�E��g�-�52��]�hr/�8��OҪ@Gչ{�s:��76������FxՕ[^+2��
בxײǳ���0׈�d��s�����:��IXZ�7ᓒeg#��ަ�|�}�����3l!���Q�
�G��-�=�z��Mq+Hp�ka����a�ss��.=�c��Eb�ۖ���+��Ͱ�/���2�e��x5w.�P,��#�;�^��!O�]9ڮ��t�wu	G;/����l�[���\U���	�:c2I������W?�w��\Up��l����1��~Ke���b�z�=}Z
'I]"���x��,�� �2.Ws^�)xEv�}��3�l]
�-���6k�`��^�9>�n@;,���tC�uƏ���]/bv;���$���}���x��X�P-	l��a�,�dB����w�k�c�#+m��?٤wY��J�\���=�dSe�pg�Ͼءv_D�'�mг{��¼9�Q��Z��<�g>9��i�G{On�_&�F�;33�9�Z/�k����Ѭ3h8���Tt5te4����O��mf�=;w���6x4q����	E
�{�������J��qv��u�K;��^�w�[C�ߢ�C�&�G/��0b��#��1�
	�ûL�P���������6X��/C��EV������������$�a?�	$��_��B���O���������HBBB_�`�>y��x4�F �F! 1��a!��B HF !	Ϙ&	�Y!cFpM  ��b �H��&� -	d�H�@�!	(D� �H D� �` X�I� � <�J  �d "  �@�F b�d ,R0 � X� ŋc$���D�����B 1�R0�"A#	 ��D��1"�B 1����$���a �$d @+$ �X� D� b�b `,H X@"$B F@ H�a #  D� �d "  �d " B! # A#ԖI� �d�2H���	B2@B I��,�b_HS����$�"��H1H������������l�E7��}Ϥo�����7���7��f�����z�{���O���$�BI��g������$��$����I!$D���O���`�?�'�P���?���I$���/���Ӧ�K���y�0��L���/��hXCE��) $����  A$ "� @  ` ��I �H 1  $I$��  0d D�I I H2I$d�� �� !�ARA�I"! �� 2$ I$�d  @� �  �@ D� Ā �� �    )!( )��(�/�����	B(�Hd$���?r~ ���7����?���=�������� I$�����g����)�?F�!���Y����Ȟ�����3��HI8�����������XI$��~@�I	'���?�$��>�?%�@�w�ě�0�I!$������]'�`g�
?��_!��V~'��$�BH��O����_����	$��|�Ih_��'������G����?�����p�%�$�O?��O���$�BI��������R}8S��h}C�(��������~�=�}��$�O��b��s��0�����}I������??�?� �������I$$	'������������C���e5�s�YPޭ� ?�s2}p$����DUURT��]b�֕)5�UP�T��U%
�QP��T�E*��R��R�E��R��I
�UD*r��kJڦ��P�6���ʍl����q�v�*��Yҷ`�V����j�۝m*4�L�Yk[i6�c��d6���h�TT�:�:�4�&-	���)�ae��m)6R��i�6ҶZ�j�jkZ�Z����.(����m���U,b�jXf�Fcfm�f��IJҴik+"�j�{��|   �{+���g[�[��+�k+�حpmvS�]�]-��i��[O�tg����QW��n���e۹5�5�Wm���9Y���6km���:��V�jv��ʥ�e��K3�[j6�  �ǐ�hP��ocC��;8C��
7��P�y�ǡB���˰�"Eޕ�B����^�n�Zۧr�Jv�q[�6�ݻp�8�s*�6]��w`b��wj�t�whk�u�[3mnU���l���v.�ie��O�u6jo�   N���t�n��m�m�v��L�۩��\��h�w1�Ki���N«W;4�tꮙ��5Ɨ��SM�mgs���΀s��r���vun.�ۥ:�2�)��U�Im�٥�  �{{���kev�t��a�]V��9��ww:���[��wZ�]�r��&��m�h*��+��e�)����z��8
�S4�f6��Si��$�����   3=��s:��*+�l�[:)�L��Vs��*��U;�6�Us�q���n�v���ݭ��æ��6�:��6�f�t�I֥S+h��o  k�A��X*���㸣jwn"���s2��.b�J�����GNv:��ᶒ��W&�AV�gm��8iA}����Z��5-�I��   -���F�u��q�\�����nH��[�t:κ��쫺�;j�  ��-�˫��
����V���GTl�EY_   > 
 {S�  ��8
 ���  [m۩@ RQ  ;�� �1ݧ ��ˠh ��  ݬV�-Z�4��P�3M�  �� =;��P�  �p  6��q� ��u4̘ �Y��t  �vp �]�� ݁Im�,�[dTҙ���m[�  ��/k��  ۥ�� ��hU 7.t� �V  ���( u�t  lM  &T�  <���R�  E=�	)*(��S�=I��d�  E?��   ��T�SS�F@	2��U  zjO���?v?��U_��˯�7�?x���)��M�P�5yդf�5���W��{���������m�oF6���m�m��m�m��6�1�@�ll��������,�T��?�3SaX>wX^cٹ�	�2%v,�(�k[�J��(9V�6�+i<�B��(�]�x�(����ʋpR2�{���2����
�X���bR���9{z�7x���
���Z��l9���v�`9���Y��h	�&�V:ժ�-�uf�ܽ�%����wOo�j�B��v�Ʃ�,�d�����PZ�U�������j��p̱L�+3L[���=;��Z�	Kx03XnKxqj��Um2,�70�F���uضh��Y����/1�Wb80����+�h`�Y��1t��ZU�b�"�~��To)�1���آ2a5�fנ�h�l��qfbGtU�a�۩Zj*�[i�՗.��VV�X.�V}3\�f��Z�:�T.�$G�.؄�d:v�=�)u�7V�ƛ��1�n���E[2�d�\-�B�2�lŮ�Խl(�nX�J�V�C6[��5���F�GGU��H͓�
�3�YRm�A��fj���/#w�dV���C72=T�Ŋ�5sa/2�d�)�tt3�S�]LEʱ�\)�-]���^U�cf�z�:��C����[����Z���#6âMmcR���
���(ݍ����uc����6�����ח,�{�)Q�Yt���Q����f�� ��3vm�V"X6��#VpK+
ލ�$��N7�E��q��P�Zf!��Z�sRMY)*1
�$��B�$y����FPl+ن�32̹KF��Xۻת�3�/1Ђ���'v��@M"nt�^֍�����S�M�נ ��ͩ�-L�Q��iz�ʍ^�]����x�Ex��7n�`�K�RԹ�̒e,{�\K���%9N;�)2�m9IQp����JϮ���`�-�9�6���CH�;�4*�Ŋ�Xm	GM]Ӽ��ok]K�P�a�{�^��Rw!�ïVָFe0���i�����֞���S4�!7uv�U����O�:���̳*m
$-�kV̧�^�St�*m"V�e�2�ݧ��AM�����*e��@��ͼ�R�K/oV��\"(e54���0���I��	e[4��6R�x���赔�.�sK�8Ŵ#ȵ��h��Ԕ-��(n���V��hwC
M��a�m�����:��n��,��Z֭i'MJ7a�S�e\ZV����V���6�3���m��+rR��P3�C�R�1ځ�67*�f��m�A��S�QDIT{�(6��Gy��t����V�k)S`����D�����P�Z5�
.�'`yQ�y�(�F;n��j*U��c%%mYi�g/ul��V��rRP�;ˀe��LǹV2杫h!�Y��$��奝[j��mb�	-���sV-k�A�Zd�"������,�Zv#n�ͺ�QJ�Wd	M���_µ��Tv�vF`���ŭQ5@��]�`̻9e�����Īe	�VK����qEH)�mG6���ɂ�Tc��tN��n",$�S�j���&M��U�f�$�X"��)�<�XY�$�^VW���YT6����aLSi0eU����%A��
޺�X�(�"3�]J���R�D[V��_ک��ՆoA���JA*�V^SS�7����� ����^�@��	�LLdj9J^�u�ј7,ACq�t1�i;4�L��@� x����/r�w;���ַ�X���7�\1����0�r�$��]\�V�̐cqˬ`�`FU��C���N��Y��[@[˅�Ek!�hYsd�I��E�p�	��p*K���V�#��m��m��!nU�� Q}�z�oy��"*`ZN:�EӏEތ���P��
��\�SF��4&mڔ6�7
{{ғ2����� �J���#(�Э/I�ˬ�+`�)�8���<td/�*=,��M�)��Њ٫��S#E�
)�33Cw����MYh[ʦĻ�P�1ZŰJnh�2�S4�
�L��n�.��5#1�T�x�!�n::QH�V���P=zS�P���H�(�S�)S�Z�l��i�M:�.S�Z�}��P0�V;tz�c���o=Y�\ ��0��q+"�ܘ�P��/
�����
�[ԍj�Wd���M���v�ݛ�n���@�Y!Ͳ K���r�42�Z5��ѷ��J�Ŧ�f���iwf�5$H�n]�j^R��1V	q}��ĊN�R����*^��u`�-A�sU��t>�8�8 z!%X�^12/J�W�:g^T��E�K2�ĥ�#%3t��b	`L�͵4&�&k��B�㘦#pj۵�a�A�m�n�h] .�7Z� f��Ge��k��T���f�۵xu���pW@�e�8�F��"'L%Gs0����Z���e����5l��V�	Y@��銡��@��n˥����ͺb�,5�ջ�����`*)��(i*\Ѡ�l���y�`�����R8ۋ$�h�(]�� �ȭ���4!c�CK��81���&�E`��n�J��&#w���Ÿ́[�?����W�#���ݼ�E`��RS%*
��T�r/��m@�Ѽ����NV�]m�:-҂�|�z��F��h�,�Q�<O~up_�R��eh	K*�<���썆pA⛵�����橘k.ր��$�,#+5�T�A�7)c+������6"�����/Mio��2�0�%�E�n�L��r�����p@�eӸ˸��"n���lTצ��w�2���٨��1���\Û��z�N'F�Ќ���^ +�qۉ�� ���w "��ņ��[[V�OS�U��bŻ��x�3|�ܨ�G��{Rr�Z,VL�q����U��� �ҏu#iaW1�:.�V�6b�&�wkh���SR�DEk��a=x�nԧ����l;X�֧�U��Q�"ɷp���b�]�M;q�u�5��H�P ����ifjm)ʂ�\�tq�x��2�Xt�Y�7���6L�nvt�p�:�GJ	kIe8S�%㖁˟eA�l���ln+ 5,�i�v�G%��EHI˓b�oU�ADZZ,��`�b�V[.�͍അy�+@0V���X��C&��c�,V��Ci�)L�ᢑ�)�%w[4��: ��U��m6՚^4��c	WVE�t9��-ea٘���J��v��7�B2��]�\�[��b����*�dӑ��f�(��LZ�A���)�k�
��'6S�	l���V���RĨ/��
C�-$[;mM-�3rk�Mcg�պ���1�/Kǎf��V������^�%c�nش32)D,܀dk3�^�me���Ow�-���+9HTWSotIb�`.�Yn�2�R �����^|̸]��Ne���(��k��x�Xԝ�o*g6���XDͶ�db�Y��Kt5�;TnɏZ���×��!�k\{W Z�{�e;Դ3�=�KV��tk����x*]���z+vV�a�6���%�Ԭ���Y���(�aܠc/qL�//]5v���:��v,�:�H���V ��PA�:?hQ��nc�@-��M�rD��VYGiZ��N�����ѹH��-Zc�0����[p�n(L�N�(<�3]��D�͹T2�a�DZ����L(����X �{[q����>hR˫ݤޙ�f��8[��	�\��Ay)��9�(
�w���m�GR�Ky��4�-P�72J8�k�":��̶����'��w�Z��#$��*Zd�MT�YuCf����۬�X>�Ww,&��K ���
.��1�V*AspV�ƯkiGi��[H�6��fl�f�*�HT�/off��¤�Qhz~x-�®��n�r����A��Ŗ-�/+�X��؆<��eA6۬�R� k8��2�F)��䩒-h�3Inl���
�����q9�֚ݺ�0�dd�����P�ܱgk �#�u6��7~�J��&*J����o�H��ɋ$jS��c���ywya�r@�5����"�R�j�nIF2�30 �Su�9NJ���D*O)V^����fB�*��͌lO6�Z�J�]�z�B�A2���X;$n&(Xˬ8�����0�8՗s*�767lm���ś[%䗷7��5D�E!
�5x@(�ܔ�*�wiRq��檙y1�lF�dI��N1.��N�AK�i^�[��Z;�5uu5,z�E��J��޻�^�O.���KNW�+H�����^�����,�Z��;I���T��4��4*�_�Y��&v�*z��4vIԪS)Z�*[W��G,c�ͱ�(���zT���;��W�1���[k(2�X�2ܙ�ya��W����i䌚W���w1h�E(���b�eh�i��5a�����0�76�B(�`'��Yֲ�6w{f!v��(|�͍��M�f�-;۳X��nh���u�V��4%�/Aܩ���äܻn�e
	(�J��F۸������%��\7G"�T��"^�7��l�K1�Fv��6��6�>��e�iނݰ�j��[��Zq�J���Ѷ� �Nm8�7V�IX�3h�y�7j����R��=�YFc�	�47w->`�)U�BLϲ�7��n�D�!F���}��-D��iS��ǁS���M�f�K0Q�j
9�����є���̣y��t��{�e�մX�yLF�L�����j4KU�^i��g+�leB�Sd��+�W��μ$����[F�eC���
r�)U��!��YH�� �.�X��d4��/�;t�,7)l`��6�elq�� -kG�m �e���K�Sm�)����.EVʐi�M�bHKC�f�VR��
�]�[�z*�U��7��gS��#�ʉ B��2��U� �ÂaZ�[�*U��i�O\���TX�J'j�1�9v���SB[���*��b�ܬygU���b;�\��z`��C�bX�`i�ն��-F�XYQ(��RC^݊*�*7gq�ķ!�6���Ƶ��ԫd#F�'���"'{��4�2KqX�2O�{Idd,A���tM:KV�����F�bU�q�nM�;�ud�b�J����	��V�����Maֹ��3GD����ľ9wF��4�tuc����L��,�6���q��%��m0�$����d�e$.HƲڂs��@)����*P�b2f�bz	�w����-�e ��ҼH��eK�K[�&։X6Jϵm�nӽ�zE,�g!boF	�4��,���>�I.�U���DXE�9�����Lc5�X��*㘕�{O�j����5�\�N���T�������Ս]���6��ۗ�.�6��jՋ�tӸ��0��4͚�2Q�Ij�
;�GYq|�WL�go8��0���Ǎ����
��u5L������*Ճ�˦@ƃ�V��Tȝ��"��u�A�9v�&��n:kMMõ��*:�fx�2������T�"�ˆ�[9�񑚬{�JJb*Ӗ��p$�D�өt�V!ǌ���)��`W4�x:���S�xl�rQ*Km>��.��'�b�a������+h���Ƕ�j�´l�:�+Z�[oql�B_חX�r���5c�1=���3t��Z2���&���l��b(�kŶ�-�+�7NVe�A�Fƞa�w��B�.b(� ���k$�#����'���,juu�
1���)�0fJzOd��okhV�[z�u�D�۪:�ʳkr�7F�+�t�i�����4��P�-f��pȎ���u#'.�͛�u�nc�a��	���،!�-�7Cɲ�˹�U2���T&�1{���AAN�z"�b����MǙY�DZ�Liu�w�*Zu�elѹ�w5& ��)���ĥ���X��%�TB�TZPn�i��!���i�V�j&���V{OA��:��Z�5��n���0�5�jk�T��n�4N��IӚ�����;���	n�*Q.�(����w�vR�1�䴪[�)P��)��,Pۘ.�]k��1�56סE�ɨ<��2m�k�;��nLi�J%Y.����e<f�T+�n��B2�Cc���Q�5��3E��i�hT`�(i�̲��X�­.�:�N��N�Q�XP�V
ݥ�i"qe+���vI��x+a��qe��[Ff+v�>�k$�XM ^��oA���;aM�0Fwdǚek��Y��3Rb�z銟7D���H�,j#r�[��#v<{��I�x�m*yf��am�.��m�k�2��P���-蕪�n݃��1�U�<�#gA��uL:�x���5VB۠�ͽ���E�P�:he�R�	Qɹ�ݵ�m�ӆ�WYYc#	$��)�I7��p'wW5d��b쵐�x�Z��\���b��� ��b%P��ܨ#ajB؎�l�n�i�E�RP����F[yl+pn˷�e��w�Z��jfY��p��9�mՉcS-AZH&Z��f�X�� �Yg-��5����\[�,IH���W!3.�㈢��x�#*E[Z���$�J��VuٌXcSZK�cr� jm]�d:ĥ�;��;)D�r�j�� �}���/f%*9on��`ҥ��Ы�Ki땴�hcZ"t��5�mI�u��*���)�q-�a]��u1n32Yz(�c{�J�b�YF���F�.;�;*�ft���x�hE��F䒐 TյOq�U���"��������兺k��X����-GF^]];Q9�R��蹃	� <ϥ�!�۸�ʛ P�ri܆-���D*<�b�0P�T�Vݿ�����%��T�@�귻L�]��q郘\�WK���oZ��sx4�f��Sn70�`ٯ�"�b�wY�*%�yw��%���)�`g4��]��\�l�s+h>M�d�˫u��,�0���;���ڻ0�����2�mQ%n�M���U��S'R���̓d���V��uSn\���ܰ,㦎�9H�`��u�^�JpeR�E5nc��x�#���oX�����W�V�d���T���>|ӵ�͹d�j����O�l��%k9Ԣm#/]�o�N�'�
5��	��e��+_Y��fce�]*�R�f]tG*tܢ��J��X;���h8^(N<]�&E�q��<SZ4�fK-��PZ�;.ms7#T�Q��45�2�P�ܭ��;|~`�)hC�r�Ys2��0:uY��B��of�+F��ِ���ӵʹ�3�.]8�V=]u�����P
�-�s��7�t��`Y���\M�s=�����8�]ݛw�Fs���gb���5�f��G�/�v:�g�V1�RJe4ko[�|&P	�v����͠��O�m�ڷp�wrAn���r�J�X��M��D���c���Ev����G:깔���EWNb.���R���YHJdQn��0T$G�W𵵷�f��ޖ�����^�U�BȮ�l#�t ���ܙ�w�d�V��㤆�YLN'F��W�']���͡��0�2��b\2��ҫ�+��V�͹�i e������h�� �7�TӦ���X����,��n�YKr����J�R�]>:�*�f]�Y���k��u�}�Y��G6٘7�M�x�fn�]]=Gy�MW�:C����3�[���9�q��V"�����y�s�aQP���R�.g yu����9wif��λܙ9��4T���u��֫����'C�����,�2���ou),�ݕh�������]Yn+4O<N��A���-�w�cC:�K؋���{�f�����Ղ��
i�sњݫƦ�t9�/������pB��f�����+y٫&��w��a�¦<�q�'|
�X]���`u�Aheٻ��D��TS��p��ODuso2�:�����z�-�O�����q�H�qYG��	��7I���uC\�)I���'����w�3pV̶w���U��{ʕ�׷P��� �L��X��n�ϥ��Wk~�G!�K��b����R��_KˑKn������l.��	s~-���v��٬peBR��։Î��(vI�L-5+펲t�Vm)Nw@�4�����Me>��ĻÍ��_�f�:��O�}5�Efs�]�ҋ�[��Xģ]��)*B.�t��	\�ob�A�ȭE�m- �ͧnT��ߞ�瞓�5�ﶽW���߶pv��­��:H�iG�n�w���{R�3b�i˻$���h6�N�}I���u\�j:��H!���΀@�K��LZ�vS��o��@j1.(�޶�j��ev�s����d[��I����@Y�x1b�eX��k&��/nvGс�
��b�Q�ǵ��:`�.�YY=�|1J<=��׸�\:��8�tN�ˡ8�]�k#B���s��+��Ry���սR����6=*$x.�	b�Iҩ��¶+�{�J�"��=�;�&�@�u���e
�>:�#4���wZ=8�y�f`�-or�\�:n��P��:h��w˟<O3$5
,x�r"!����)U���_��jaf��؅VB�T�q�R�u.��������sN!ë6,qo0�<�ml�Nv*�כ"�It���V6}������ �V�0fu�)�����Jf�GS.�	>Λq��WHY��wt6�#����sv�!td��@N�tլ���4D7Cژ����]bB���E��(Kc#wt�	�8�ϐ��j�ԫ[������m_R�%tpL>K��ɥ	g���J�g�i�t��`�OV�����m�+h��aW�.�49�A8"� ��o�V����ݢ����,�%a�SBYX6r�u|��XX�b�	,�퉵"�)���BGyr���vb��:��A�8�2P֍�pB1�f��C)"��4�P�w3�C=|ҁ���5��gj]e6w��>چ�i�z�&�Z�5kM�7�s8��-jʚ�F-�9����d�^��T;�P���n�7l�6�e�"ҦV,��k�A���;e0�6���dnT�j\��t�B��9��Ũ�OZ��6mn.F�PY��%�\[ʻ3lF8pBY��}��8���ܤ����	Zi����fc��\�7��Kmas���V٥�3�Hq�Nm��
�^$�EpUG�h/m�ي�;�|��=L�>fr�9�}���#�y
��LW�t�R���b]�q_2��8LΔXx5*wS̓��-s�U��jpf���@�{un�*�K�ŗ)0�Wh��8iY|M���iQ�����d�孕o�'��S�.vr�x�ű���2��|7��X��1���v�6ԑ�n(�lsձ&X��k��6*�@�|kp�Hp���Wo=z�wm�F�B�rQ�)�!��q	Y�oQWF`��z��w��V(
"��>ѕ�a�c9Ҩ�R�.vjwi-6_Ix�/�L��V�:�u�J��@��T#h9(n2F�#��pwֵ�1n�;pQ��X��K������5]�s��i�E������Z�p�=�Ӝ�P��$r�� TS5(�y\yU�ߵ�J۵b��� e)�i��嗻�l���C ��4k1��C�.:&��&o�F/������s�]{V/��N�L`���s��ߜÍ���l�����n�Y/�Uk����|F����)�*������9�
�4�U��Vֲ.��na�h�D��]�{���������@�.��TS�2W�,
w���6����r�(:�(��)Vj������ە�'��8��k-TB�o�������c�����l��2_6|�mx�U���(Atƫ0l�2lݪ��.`.R����˱�;}�>�/�M���^kYH��^�rP�HT'^w��� �}����pZr�������t���h������ؘL��Z�e��S:�"k(v�͗#�p<�r`:�E�γ��:wY\�l�jNӀԮ�,7I�WI�r���u�p&,p�9��\��u�z�+��J+P�w�#{j�aJ�
8��N�_Xv\���]�ʧp2h�u�/C\�2���Z6�}�Q*0(r�qV�e�W��7�:�	NHT��5ѺFܽv�d�-8w&r��/���*7K�Y���
.���#v5���z���]�x�8�X�9u^�hTS�ͺi2��6.��v���a�����Q���,����ov G`���pd�BɄ��Q�L�¯ 诓�J	c.b���&4ta�s�Tf�Y�9��⌑[��kr��<K)��IE[wdʑ���wA6�u�岘�� {��:���8dєk����eu=Q��1Yإ�ΫO:�&��n<��II�p];H���J7��$��N�u�@�ssjc���qq�cE��*����P펡1ǇS]�dְ�dZ����r�z"��GXJ����Hv�Ud]C��(� �m*C�f�o�X	t�#��@����e�+{��NY�3@���jj���$�r��8�0�������ʕky�)s��ғ���9�د�J�x`&�����{����\#��\��"j��ؒ�p
e�iU�k`�䫡���A���+e�"Lc+$Y�eV�G��'w��;TT��=���g�>�.) /f��,9vpf�9��aJ���Y��+i�w����fT=۷�E��ֹo���1m���C��Sj�F�2��3X����C�!�{�n�_\ά@�����E��!^���⺭A��3U,��&ه"�����+쬫l���U5о��n#us����H��[x�<�(s���Y�Ua���V���uN"��͜�t� ]�RV�;�L
�[��W�����VJK5ג��,�I�7G��1l	�����2Z 5qz�Ӽژ����i]��S���L�e �r���'w��AF*A���Ǯ���;+2�F�Ǭ`�(�{Tw��N�%�q����I�,��Xn�C��,��@��w�e1���u��Y�Et��6������ݪJ�eҳ0��)�(Q�+-����Z�oHJw�R�w�.:D��,�^"�|雒��m��)\����]+���{y���s���ک%zڞޭd�|�WB�T��,�#��;-N�8,V��C���N;9㯖yyا�ulH���7}�nYЯ��q�����8*YQ�RUЛ��癔o���F�Y��Ii��-ʺYY�e+>`�D ����d�,d����1�>�u�HP0R�{mgb��{����>H�V���^�wGj����3��vC�2T
���"͢�brF.� jY��ݺ��8�Z3�aF�/b�Jf����8��vcx*�p����U��4�s,;x����D��}·ha--��|�h8[�招m��k�*��X�]�v�֢�O��E��:����瓂��w�j2Lޝ�����8N[�S�[aY$���<�s��T���FV�u�.Rţ��7��Ʒ�Xk)�лsmo�m�<�r��L������}cP�i��S��y�Tژ��Ewm:$�7�L�'Z%S��ˋG �b���S�mf]L 1�޽_\�w����sU�m�O���髝�*�R��tp�a-aB��AWrKE��r�-��ռ�d���uq�oZ�����ަ_9w>ީ��w��,+��ݽ��{����BtTƪ�}��Fǘ�;����:��̡X�:�+�]�X�*�d��X��*�"�$.���kv��K}`Ԗ�VZ�%f�f��G7�����m�q��J��n��z�ohg�m�`H^�Ȝ\"��:T��uV�9�Ȼ��-.�pWu�ITҢ��c�0w���ej1[5����s�f,��jWN��j;��'	���5
��V��dAM��vr���`uo��O3W�*��f�Yd��(m�yg���|]�Rv 'Sv����tC�ˣ���{M釰��U:�_U�EPqa�El���fڹ��.[���w�^m�)�s+��$��'�ms��8��%���kW�#u��T0󙦟�ŝ��IDޚ��I�+���%�j�\*l�����[�mծ�tVή�@��[{���Wo��J���+�8���"S��L���t�WM�L����x��Ӟ�1�-��"^�'�����P�jhK��Gj�=���Bq�ȅ]
8a۵8��^Ö��6�S���5����8�%;^Y��Au�fu���Ó@��<���$4᧪,�)����]�˭���n6���:���u�J��MS�躍����t�*p�g]��a�[���1U�֌虳�x5�ɛ­�a#����L=�j>��7�70w��0�;Qa5����^H_��t|oZ�Ӆj2���ju�Lڼ����24�0�{��--S��B�����$Ⴉ�9]/�-�<���)�zbvs2���eb��d&J1�֮9q��,cw�����#�%�:oUd7b�}Nsf�Vf^Ns6j�6���y��l�`�JY�o-\�ʹs3M�=oK�>�hD
�0DYcP�o�ae'5WU���X��n��6ȗi�vJ���`D:��B�kz�3kH��Q�I1���4��כK��虶S��.���X��	&Җv�ڍ���w8X�v��X��4(Y�4��);wqλҴ�:�C������܂j�&DN��7*�\�A{,���}�J#x>f�� �lq�|��+��1Zܗ7_V�{o-����x���K����a��<�-7��9];O9�������z^7�lg}������ʉ��ɷC>uȨ�.eWu�ں�8(���)ֵ78�V�Qt�[�Ӭq��Wfi|lsV+ma����K�,b�+��gA��(�
q�v�0Q�����K��V�>�r��{sn�E��F�.#{��(m�������������Z�����+U�v�����܏`h��z����j2�έX�J&�=�.?�b_ݼ�5��6��*$�4���P�ZO��pb��n�U����0Gp��֏9�T-��;������-�z�ܙ��m�Z� �ֺ�� �aވ��m�؀g��i�̕b�/�0�f���ċ��M��"�M��ܷ l�/{C���r�Ԡ�H(U�~/�ʸ�q��C�;�)2q2�nwe���ɬ'U�F��դo�7&b�Ǳ,�ޔ�u�o�w�W�l�X���ywSU��}]�oow��J͊B�C���q����>.�2��OqX����]t�֛t��U�*�"�yx��.��Čy����o4k5�!��u�n��w4e2�1齻ze��-�N>ś[�Z��b��7r�N�-q���a����ܪ�|�Q��C'��g{��4���v��1�"�YR��H�]�H)D��Hc���u�-ӹ��ڊZ.�ebH}�Ve�)2]��'�.��K5�j�ٴ���b�0ձ�K]����Eԥ�ץ���\TKr�0٣�����
喝��n�)��Loa���c�Lv<����������-��9Փ �n�1����'��5�����H����I�St�o���!�^���4�q f�G�8�6���kj�a\L{�gF/�iws6{�.S�^���6�h��U�r斧0O2:����:P�l΅����I]��M,9�M��ҡ������m*K�t$1eXKk[�.�n��׎�s�j��6];�S��� ~�n��p�ʋwWHgN�踐���;�>�z�wvwl8�݀��#;_3�ֹ($�^�88�⩳�LJ���/r�$l,ʵ����P�o|7E[{�Y�|�;��԰�#60����A���������6N��=�{��  =� ����>��>���wZ��_����h��qN�u���[���G�NH۫�Ď7Zo�'�vC��g�E-���#x��k���wbm
#�'���-�|�\΀�z���������Wp�����N\t���3m䔝���[�h��WUСe5fbB(��R�CB/flܑ�$�ق>N^�ى���V|ذ����q�.�l���tGeC����ND蝙��C�N�.kܔiK��d_d���Ą��ٜ�қ�h�-�Ɯ�ЌoZ�W:��NH�X��KjQ=x����b�e�*v�;Z�g�z�t	m����59�Yy`���<W5OZ���4��-J��]�Gwt�kc���g_'��*�:�3�g+#g�C3��SQ�)V�g�=�t��I	P��#�Si.5t�>�Ɨ3RJS[�۝�M5X��������Y2�xkR�ծ27h�pp����a��ݸw`ν�tR��T0a�,�c�o"u*r�b��*�0ǧ�nA�ߣ9o�˭8X��ɃWvpg^1�RӰ����%��R���2��V�q��v�jn.=9���E�U���$�����6�nA�ü�i3x��Zn�8[�cti_w;����c�IX�fr�R�N�s)LK_B�<�#�RYu��5kVV+v��������4�ܡ7*���2�f�m(��n+b���YK1�Z}���6�Sb���\˙va�5�+���|P�ʔ:Y��.�֖�.�;�-�k�ms�'VU��������W2=���J�Mh�LFYf�:���8bL��YcF\]؄��&��Ň8���\"�5+&0F_)�tA���&���rv���u3(Rl��5�k��o[A��E<���Nҙ�l�i"�}y��Ӡ��s�·Q��$*8޳����c
wX��L�`"�0�v�;��m��₲�X&��ĭipR��ur�g׫*�]�6���MT��ҮoEu��)���s+.x�
�>�7[F��fB�]��{n���T�u�� �E���tg[ʈ���w�e�kx$�t��$k���M�u�${�vLi��zK���Q|����Su|I�B���th�%����N� �,�4���vB�e�$b)Q�EƷr�]����i�غ��O
vF����T�\WD:m@a�^�-e��
E�WeU��ζ6��(U�7�޹sI�u\Y�-�2��va]�@�gv����E۬��X��vt���xL�"�[�}.��h��ms��*�Y�"ƙ�Q"U2�۽�[�`}��g>�gU�k��Xbj�����S+W����o�*�ǽJ���`�Z1���r�u�N�Q�H�,ih(_P���!��;.�s�-�yB����H�bn�2�����}��p�q�j�u��C	L�ӕ-t��f�W��Cll�:�ә�աq�L�h�WN��$hx�Țv0m��֌�y�kb �НkZƺ�#5�Z]�`��)u�*�°���ul�Fm��ax�[iGQ��*�J�ٜ�\Yz����l7t��4�6��"�fD���1e�uv.��WDC�N�.�M֦��K�;wo���j��&6��:i�A
	<C����ur�YZ����ټ�n�ޱ�K[�%��k։�
�L�☻`�ä�鰂w��M^�l�1GW8I��a�vd7����x���nJ�3t�0��qAv���<2����h�@��3~�a��qTY���]��F�vR�֨	g�ع,�\�/-�����jV����5�]{[�V�k��y�(�o�-��ާ��\"Qh�RDc��}z�N���f�ʖ�iA�E�4u��kyxF*X+{)���*mI�1�@���t�yq���RR�P�nvM�gܷY�9����=��z@7i�J*�N���c�Qc�;�wc�j�'Iz�ҪU@���oGxh%6��4Fp�x�뭇h�-J�YaXٌU��-��Z����R5�k�}I�\4�5z3u�hi�(�;fW+�c������l	��G'�S9eY��X^����o�`���K�e�.n��2Fv�CrI����t���:�y�o���9�_s�Y�f�k��|6>���pdpX�rxi�@�yp�5R�:Y�b� �.�.�v>]WG)'R�0���Z�q ��£�o�2>BΗ��i)293-���:�ع����Fn]�L���76�����tY]Z�W��:�0'2�eK�c�B�XF�[�h����H=m͛X��	Gm�q\�r���X��m[�]��}}ˉ1��eɲY8��j{�s�w��ٮ�FԹ��e��Vӭ���Tf�3��E��0�V.±�A����X�yC"(Aiw=�m@X������)��+�NjQ@�ˬ����D���0
T*o�]C�(|Φ��O���.�$�����]Y��e�2[hL5Ns�E���7֛��̂����h��+��O2V �Һ�g~kl����\��%)a�Ӧa��I�y5�.��6C���X �Qi��ྏ\Δ(�jjtT80��2�u�,�Lc���a����ղj�{]�p�g
!S�*Gm�^�qȞl���`�	ݘ�9�:����s 2�+T�w3�j&��R�j�q�	��s!�x��W#�ƭ@֭�)��_�jV��H2��Ά�.Es��7�WQܠ�T�9}ӎ�GZ@�A%���L�lɨRM�s�Yb���<�
�A�,Y�bΝ�M�����S�i[#/:�ۤ��K�3t��-�(F*� ����i��y�7d�#��\Vq����˵����T����Cjڣ�7k��_�w;z�����j��Tz��
̹�J�
�e-��a���4����;���¢U۔�-U� q�0m��Mw]�f�3[+T�2����&�˭iH���-Q�Ӂ7��=!v�/��,�����o��+�P�\I'W*��n�[�]�����3�\���Q<C���/�51ƴn�QR�&ދ�f�<N�[u��r�,Z�)���Oe$�$�v�(��*�[���ʊ�o-�\9(�km!uaXܵ�8��;�2S1LEǻt�'!�0\E��0]��L�_^�ͧ������'d�7\��8���&Q���`��+ESn�2���.Ɗ�x,��j��W?�)�un�i�j���XU��]N�o�*�qGP9�,���TۏPX�jH�.�Ln���f3�K�Z�*�=R�(Mw�k�$-�5��!Dg��2Ț~.��[����1*r��F�*.�yk�su�ǷLZ�� �h7��T�ˎ�����o5��ʼ����1p�����r��ֆ�G}ԚmYM�h)n��H@�Q��|�t��Y��M�ik��A<:��Nջ���8��R7��6>����xC�F:S1l��Zn�>�H@�j١M&(�NS��U���ٲhuFkPT�iSc0>�ϥ��z�Jw"�>)=�1���Ⱥ�ay��a������$6�Zo�0���\Ɇ��-YԖcX)ث<U`�;��'�
c�{mkս�I����9F��bp)�q?;7om�u���$G�J���n��ƈ��W4�<"h�r�L�|�v�H��3�5�������u�R���]f�E�EY9��gg+
�큦�����׎���j<sJ�T�m�u��iqb-�]�.��:O�k�Pv�щ�:�\|4ƈ�����.�O%��Wz�.��@��ٌ�acl}S -�a.��T"u�%#�ma����]YO;��n�u�SxAseG����Tffa���(��X���U��1���b�J儼����әN���-����M�d�Q*���6��H!��G,JN���E+��Up��1Y�sr�fm����D�=�l{���M�u�cD��;!�&��#h��ަo�m�!Z1hs��i�y�W\��4�(*M�Q�vV�Q�u��ܦ��"��7�մZɓ�;<ge6��n8졽���l�*�g�w��Y7׍�25,uaZz[��Gv�j��1�G��ʆ�nӃ\�6<J�⩇W�Kfx:ꉺ���Vȧl�e�b렃�ҽ\�֐f��p�\"��w-����?s��4�P��Ӓ��E=d��]�x����w"�E�dɅ �h��>
\��3rj�HԦ~$ �v YΥ�zfRia�����[͍֔�$���PN��q�P�wj��Ҷ���6_;��7�˲k�ɨ7�Y�U"9:�4*���(���˼:i8gWb�M���Zv�p4��ݚ������׬�T*��W���Y�6��9��c:7F���ԙ�EfW*�]=#4��<u��;����a���S��c�5�9�M��v��2^֜�b�{R84U�u\��Lˋd��i(li���)�ЙZ�웦�Sǩ�-��hb�Z�(I��;eL��:Pn�Z����*0���K���r�󺱯j�s0JU�`�������N��mJ�=6����eC�M�5/bw�%�����+�'P�n�*���7I�q2��2[�����Ƙ������A�5,�)��ŵ��a8:�shδ���m��|y�	�K% I�_M;YWLŒ\ەp�7����ɤ��<8N�&X;U	v�c��M�V���#V%&�W��H�R��+�:�c�����9���6;m�[Y��0���	�f�e��+���oX6/�����޶i^����r'S-*؋�\/j��D��u�3H�z�����9}Т���h�����FT��q)un�Щ��\' �X*?���#w�8��}G���Ս�Q���A��D�vu\����nQ�E�>�v,P��L�F*��WgE���=�6�wI%��I𻧱h|B���D�vGk6��&e�V�ʗ�C:jk���B˺SE��6�:]�q�s)ԁ4]r��w�Uvi�k��5��=Qj�Z�d���F!F�-jh��-�ɳ���wpYZ��m��2�N�a���vFP��7��H��2�f%�\2�PK�5�h
��<�ƈ����r�A=
j0�8�RHS�^�9��:Mv�$.�J����	�2���j�.����ʺ�t�*�esXS/ml⬵ܑr�!	3�p�Xlb��+�*�9B�7�s�<��z��ᕙ�����y-�ءZ���{������Y&܆�Ųc����H+����՞ŷnj�)���3��h�Kz�Xұ���8��3��Eۢ����0E���;�:�A���� ���u�TƄ�VS�汝�F]���Ьԛ�5�giѭpb�8�@�{)�4�3��IoD [���C�㌣����-I��j텪X��WY��p���2]^At֍�;�[n�v3P�p �-VR�N������7+��Yc5'��n��lJyM���Zc�4f�ں��v_% B���f*�s,|���b����N���Zc���	r^��Ɋ��$�ʜ�%��4��`yi+��*���b���u�B���q�SgiK�lB�*�Ȱ�����.!CZϷE�83(Z�2�e��K5�Pq��AݷL�4H��!�![[t��m�P�b���/�(e!aU�c�y��3����¡�Aּ�8�]:�P�}{8T:�\�q���)W��rL��۾��%
aǴ�l!^Z�*>r-O^�+F"%)WC�Q�fg=���tR᫽3kA�}��h�
�ޤh;ʡ&��3h�bDZ���,�	�q�F	�2s���1�:�ǂ�.XQ��g	�k�"��\�rIaI|*n��QN!�`r�]���d͝ճ�fL�ғcq������o��hX�D�J�`��F�Ve�M�L�� Y��c���xr�b�����otB��:���V��n��6W\�,ky����؜�&/���5ѡ�����G�-n\�4*����/U��ݮd��K}4���:��ŭ��K�]�Y����+ճ�Q7 ��*ʜ+�m�]v���Br=��-	���R��I/�G���9$��wwT�ø����X����򣊴mc�m��sB�/2���[��P�@�C,�gfO�������ô��=�vVb�6�w(�&��id����}|��m\�x��ΓUHnK<7�չ׭��&{Y�n�U;ERI��R�^5Zz��>�>���ܩMȶ�h�p�aƮ��wIR�k ���o&^]�����|�#42T{�wt�Cv��J4�������՘�F�z���w�!��,�	��U���^�vX(���s�܁�EX���.ܷA"�Y.������U��	Q��[V�cحڢ�`�ԷB��&��l��v��h,;�n��πH�}T%��G�Mf��a���{�+Ѕ]kZ�Xڸ-o<]���-���:\۵Y*+��(�5ʁ��yśQ��s�K�&;Pj��Y��ʡ�wn�i4����g8(x$e�,ᡛ�R�28�G�G��.�LR�{v��8����;�λ+��gN��\��;�M@w�>z��u.���Ѓ+iWZ	@Z�s+ �9���Hއs�Y���]�S�o]X@�����늂mj)"����I8*c�Z�C/q�)��8������AW�:g��L�zиZs�e�U}Z�+.�}��^Ӛ�F���;*s�-�k�S�9,�+�+���}��2uvd����ea�D�Kr�F��)֡����8f�NE�����ԉ�r�����J�XE�չ��9�	��y��1�֡�BpD(p�J�Gx�>[!H#2�D]�s2�>3��s[x�j�mD���؝Z��k�+k�˴oԋT���0ώh�ڝ�����'f��Mڜ�VH�	j��:)�Xi���)�
�Y�����%%�Ck&C���%�V_.k'K�]��G�7;�nX�Y��#Κ�=q�Mq?�=�{�x{�~�7�r���{}+%cas�}Yd�K"b��Xn�B�6&��;�օ˨�۩A.�r���1���d��ﳓS�o#đ}5stՖɸ�kR4���R�a��x�X䖛޻��zbF`�ɛm��IM�L
߭����r�j�����kF���Is��U�V5��
���Pۜ�oF��K�/)֫& ��L�W�L_l��Y؍�"z���C]��ڼ�C�D��Uv������˖�6�in�sJ-4�Ν����6R�cn�'�Nce1�G�h�WW)��H\�b�{76�FdE���J�Lk]���*�a�c8s���-���y��|9��S����_Z�����*�5��I]���qFR�?Ã�z�Fc�n��^�v�Jڮd�:�e�EW$�vgN*M,��p�շ\��a�7AF���:cl��- ��]�U�{���x�EoX\���$b�YoQ�|m�޷���K�wU����4��������^�y�5S@���a�Cm<y/�L<T�-Zuqc��!�/_o��S'D��8U���y�R�Lв�%=�5�m`�2a����;�i]��)�]�q���'Z��oTh���nj�^�8�fm��B���G��U�)�Lmj��Z�.2&ӧ@+�/0�gLT��U��{�:v��`�3e��Wƃ8���_d04�);������(Y�ܮJ��$pV����]�ml͝w��ۓ
B�SJ�ZBUE=r����sB��e�.���T͖����.�r��$�OA+�����֧���{�����/U*
$%	R)n��;�^���RF�Ԉ�T�a�B��JH�7q�����)���v^���Gt9fI��;�V�������wst�)�=�N�A���X�V��ĝZX�4����Ts���eͦZNB�=$�F]Gu�V��.Jy��qqeV�9�y���t-Ww%��^V�W=�r=*��rvjDUD���̪8����S�^QQU�R��J�\'P�
���AKSBrO�0�x�#ԫ�%��J9�(�7%�V�Kt�
���$�ԉ�uHse�U��j���\=�;��GL���DT���".Su9�Ӭ��9\�B�ꈇ"������M�QJ!d{��� �!��+�nn4r,)���ҩ�j�wA�*h�IC�==��S	�<WE��:Wo9�
�bøC�;�zd�Z/x�.�_�꛼�M,�0��*�h�{���׶�j����pر6��e#"��$��o���<�fw �w�$P�5�5��r���x���|̭�Xq�;�M.ț�w8��jz���*�����
�%�d�a\+!�\_vE~*�)-��q*x����rH�=��|��e_�j��{��]K�c6X�@l-�B�
��B*���|�r�ŵ�)ݾ�k��!)@�eT��*����f���'��M���d1G�u�F�*Z�mv�F�y�k#e�N�Q����p0Ndyr���Ӓ/�om�u�w���h����k=�N��ꐂ�/�;��EW�,`��n��BNN�}c:\K8�vɌ��mv�>	���[;k�<]Vv���r��U3����T5~/��t7�[��|zܒ����.�kleB�Σ��9cF�<s�	��ٔ^��y2�0j����w����z���F�5<�K���l����Gm�p�]1y��#��HŬ@W�%�3��xG=S��ԬR�t��**ef����nm���Y�MF��/8nH�)Szv�i��U�;�j�+�A��T���{����������-��Ø^��gvV�����_A�[���R<ɼxr8�r֞��)����%�v��T�������R!�!kN��/�����n������f���� oD�e*����F�u�`d�&�ԧs�TLRu�E�6��|'��C�&!;ydt�7�M�O��f�������_#U�4V�'��TLpwb�j����qP�P"�y$1�*j���*��Ž�W��)d�L���F!����n�ߔ��V�"��/�M+���Ts1�vu8�1v�W��{�3�{�
q��˙�S�z&P�
�>U+�h3废�Bj�۷K�'M��Vݻ�y4g�����U��&��&�<�/⫰ܥ
sȎtkl�GpW�c<r�ףt��9˞D'�ĵ�=�c��jca9��S��ej�Jӟ#Z1�I��%�
�	�J�����R9波BnPrh!��qa�*�X���t��e�O����V�X���Ȃ�EV��C����C�֜�ˋ|�*{��k��3S�P���)��$0o��P"J���3ZN'�7����s�60���տ:�6���>]X;�oVDM�A��2�8=YX�%:�����g���4h)�L���@71Z����iVX.�Q�whCa����ɷ]C��g�"�b���4��>;�+���v��2�\%U�7|�󛷷Zr�rVf��ۮN��Sam`��ͤ�W�ӓ��Z*>֠�e[�m.��\4�wy�E�|�cQR�I�ؖv���֌̽�@X~�g��V�\�y+eZ�E��x:}��{�u��B=~'��w��"��n*�	�]��ۜ���F�Ȝ�T���VN9�����&�+6�r�ۓ���a�*�ƕ0m�GtЋ����p�h�#��J�n*��.a�mۻ]}��ǘ��
Χ9S�\uTPV3���&%�����L^B{e��# �*�1��sn�Q�Բ6��� �x�Qf8u]TjfW�0^8����%\�B�Ջ��,�Q�;���8npd���tH�W�
��Y���o\>��^�����/�z��{M��v�+�0�]F�;'����1����%���A���DH>
�1<��$����U���m_f�+x��a�N�Fꠅp	l�-���%K�!�j�΋�:��m]M.ur�ԛ�f4V�\�՞��dO��Mp��[踟�<ѐ��^��5IwrQAea�1��'hvC�V��g�˓�<���4�4�R�>e^���)l!���`�s��X�"����kab�KjH�]a:ɖ5l��
�aY�(]�<�̎렑Wn��$L8�U�v������{���N���q� b�B�s�,���Zrv�?pڼ�5��#���/e��3ޟ	Z��t(��_��j#���ˡ=? f����;P�#t�1�U81��tH��2�w�M�w^V����;�!�F�cE���b��R�Z�ƬJ�]�N�ka�/��A���t�����t�'�,7�/1�K��0�_�0��K2�}`��yZ��k���Dh��˸��6w��0�\L��ܘb��a���)Xx~ԯb�8����߈W(�˸��j�r9�j(��グ������D��^%�+|.Zb�(�|����|�aN��p�o
ӈ��}[HSG}NK�{�|�/�(*W���]I�9��?b
�۹��v�q�Xp_�3V)Ƨ�;#U1 [r��E)���̸��B8}:��3�Y�����c8z��+�U�5��]D�����]U�U��k��0�]:a�-�Vn�W�kzj�D�=7��y�(v�zHcT���W�E^UG3}K����X�Րi�u��%����NR1Ε!���C��p���<�S<|�C�xp@�͕}�M٭���(�{<:�V�Wbŧɷi�kA�%^msC�*)bb��p���<�,���Y.�{�.6�ҩ��RS�4\9E���	W=sz�v�_=b�q�}7�S�/��X���jj%퇳����͎��-B�K��]�)�Ln���.�p�:tC1E���Ɨ���g!����-;c>��(�@a5y��yp�ofܡt_�j�}���_m����w䝤c!��3���P���e�J���i����!d�M̹�z�R nd#S�L,j�<�7�Ok��g��.�&)J&:��7˶�:u��S��SoWG$S����L��:���H<�|���hE3a��פʴq�!v�>��n���V=O��Z(�- =���T�k�ea��C�����}V��b��Z�k���[�U`u[�0�S�Ƞ�xm�+��5�<E��>fo*�[��V�x,�.`]WA(;��ܔ��G[1��{����°:p����8��5j�ցΤsz�z�w[c
^��僧=���9�b�Ƣ����p�� u��+�Q�A���L t���Q�����-i�#ᮾ*�lB[y���/�2>d��顖��� {
X��s��p�ka���ۥ­W,1���C{O�l�b�!�۔��<-9"ὤ _:�����s5P/�ҳ��[�͢����
м��.�l�\y�9˴�[#;���)�|�|+u��]��&��U�	��iq=U�'�<�if(���6�x�g`���B���o׺P�'g0��%X�Q�È�sO��h`��+���]'Ǘr7.(4�t���ƣuE����q�~Ų��X��`g�ذ�����_K�aֶ&�����u�)ښ���5�
����z������)��E�x(����Y
v�.0uo�4M�R�C���[���/T�r"X���O|��O}�MJWg��9�X��P�y=Sn�+��j��k�l��w��E�P�eqϯ]G�q�|qq��du2�N�"�mfU�2��W%�n��q����-���S/O}+{<֑��-�}<��L��]�J}X�����I1��_#̭��`D�Ru�E��o>�:;N㑆i<ya�y@A�UIn���[5mwC!iH��>g��L�v�����BA�� ـ�&Q�N��B}H>��`b��|�Mla#C�;}TnK��~C��ڢgWؘ;����^}]�by��Z�ś�M>Lm�$\-��Ü GCRD�%Nɹ���8}q*w@L�	�a�;�gm���n��k���T1p�q'��7k��<�,��7)GO";P��'ۏ���V6������zvg6V�*�o)����[��7�(TFv��	S�!ڒkQ�� lLŚ�جX���*��.����ε��N�L-u�sCYY��1���,\�pz��U�#LX��ʶ�>1*�Y�05���H��G������G,�����)�D�;n�/�����@�S��뢸��m���S	�����`<�<�:�>�N�;}E������/����y�Fg��І3�c�Y,Xr:a5 ��s�aeD��Gd��{���|�|�	�F�U,t7t4��k�k鰀},1�d��e��h�ݳd�Wc:��ބb�_TC�'I?ft���
�ߊm!�޻�H &��k���~��]3��]��T,�zbA�����@x8o�k�ʷ��}y�8~b�xg��2»Iew����&y �t���u����Ƈ}
ϫH�c�k#0ڵ`�H����nho���9>w�U��r]0��l��5:`�tِ2)1�Wyq��=}�R����:)���W�W��i���)�^��^�T� w�QAX�l�i�h��vQ��2�o���l
S��n{6[��I>zM.W>�6�M�
��5�]L�����8J:��x�_�NX��^TvTXxܛ���Z���N�����:��� ;��
����<�ݘ�I��Ȁ�Bl�[�9��n�����yqJ]3��6v���E^4q��8i���=��J-Վ�X����K���:�b�$�b�_;ݝ��湚��ֽZjg�'9�d�n�O0��/�[��>e�*���2޾=L��X����|K�
W���W�Y��r�9�4�'����0Z�8�m���\SAFJ%�_/w���`eF���CW������ȽQi>kgjaC�P���ϙ4�N
�w�!9�!p %�q0PU��H�0�/��j�5�����u�ʓ7�������Y1�8rrt�{�"�ʒ�1�jbc��@tSݼ�*�m<(��a�����F�aW�O+|ҟx�j�������ϰ���3��*x��zL�;Շ~[��o�VZ�)cw u!�U�$��r�58$`֞�o�+���:��^�`�.ӑG^�Y��;'4��:��Q	Y�9���WK�q�y-]6��UH��P�Ɗ���o�u�ha��S{\S�@`�tg.�3O��IlQ�ތQ�s2�)U�����4�XϹ��,�v��/	�2�XXn$�^��N�on��������y2���ח�88=�pm?(~>{[��c|�9Hd���I�y��{�:���Z��t��/P5K�na���|k�Z}�aw��g���h+Z�7N35�=�Će���.ة�7�Fԡb��J{��ّ�̢Sꪷ����������n�o+p�8+EւS8� I�r�Eۥ��MR^���k��Y\��(Ԓ�����)�E[�o�����' sUk[*es��Vi��ZU�� /��޸6�9?
�릌g�pu}��pn����ݡ�f�U����Dч�_�1b4�L�چ�b�mW�����#]���������]Z��!�*<!6�;��,��KK�xw(��ig�t�F��m��?M�~�̱��JZ�wގp�c��W��?up��l�����<�3�OԪ��p����Ps-�����rr������	�g�C���e����TW� B�N�N8�wR����2�����a�����F$�#悤��4S�b��%�qB��f��[��籟n�����¦���L+Ư��o��8�Od؈�Q�S	�g2��o��8`��D��A+�e���'m�6Vm��u����%l����)Fz���R5��D�ND��3����^3��.�᮸S��b����H�&޳�H�M��Ů��8z@�jc _'�ȵ�E^4��d�F���^��E����M�ůc��%p��6�I<��r�n��H�dt�&Z�e�fY��L"�tt`������D0��j�y�\VS�ģ)��w6	�r�Jq��c<72�X�˄��W���J�����Sk[W}�É<-;�۴*�c�f	{�BÂ�(.1pt�,�vh9+�H�M*v)F�O���~�_{��<۪�	�q;�W
��5�uںqJ�l�J�[8�=Ӵg�u��l����3����F1���a=�����~,�^+�hQ?��-�n�Ss���=˻p!eQ�")`�}�	���Cζ�t�]�����?��Z������^R5��+u�����³g��8����� \s��seW$G�I�fo����_r��L���41i�ϯ�`vX�}�*%�ʕ��{>컧�����lS�F�p���nߤߎ�UY�h<:%�W�^��r4��s�}�'��ޱ9i^]��8����0�˖!i�jP�o�W϶@��u�3��~5�F#�C��C֧��c�1��ҫ �9l�v��
�3������4��H����=�����9{ܲt�j�q<�S$=�����pd�=�zjU���ӂ8F���hD�oe���:�q�da��T�!�&�enj�"b��9�_'�{N�]}_;[��<�آ�y`��ջ�����[f�gk&���ֳ��������ӻ����{f�B��p\���|�^���&
Z�[�IoWO2�0�8B��<b�S-�lۋ49*i�3c��*�P��_uPC.&T4��k�������0�1>	��Q͉ܰ�<�����S�]�]M�/	��bkFU5t9�M��@�(��T5�-�]���a�φy�����UnOR.�]goD)�*jn��z�d�+�(�"��C�:�sU��%o*/zX��]N���������V�R|��SfSXi��G��fq_\����7Kk�n��;��\4����d�m+�:������l�t�	/�n�Q�F7[+W}˹ڬ�()�yI*fu�鹦4w���aݮǍ�0�͇���W��-�ٜ�vZ�B�p�1�"q�C�L��It�=f�K��͙���n�P��V*d^�}4:���N�S�
���q�"tm̭I�Y���ݜ)t΋A�[�fY`R�h���޳M>�M�Y�K��cAˣ��j�:��Dㆪ�k\��T�fu�a*�o�d��z]��5%gks�M�޻��.T�v�[��Tո�0sV"����݃�Mn��Kf��5{V�M"����~�y�a���W��IdOw�����;��G6�ٔqɶ�S*�h�i���N��<��]`��L���*��V�*3ͻ���f���^Uo83"�onV�/K��B�hy
�=���H
��l��vgQލ��>>��v9Ƈ�Uo��+EŊ�x8:�������P;6Y�կ6��v�Ǹ��SV�t��q�-N}��7���]Zd/r���kT�=����F�J�@�Sn�m]�	}pж^+݆`t��z��	�L�"
��Nً+�:n�J��N�n�*�1t'8���d�k)�Һ7�j�7�7#}ǲ�,�"���x��7H;J�y8�x��h�2"0S�r7>ʹ"UV̬�����Xs��u�u9��Λb2:��CV�̮�����TY���-*��q���v�\ꋤ�tE��%��C5�6����eʣōޚm���C��F���`�S�ַS�d��*��sw*�q��v���`2�Zk�����l��l�y�R%4%�W7lG�lWK��>Ů���/���R�+�""��&��5ԑ�e]u�op��Ѩz�<șA��F~�gRED�Y�3,�Q�:�yx�.=�v��2��޹����m��hހ�lBq���b��ۂ�c�����e����u�*Z=/I�L(f�e�΂m�HS\{]rF>{r.olvhq�A>�v�)4���%z�PӲ��=]��{C q�t����6�ԩ�V"�[O�
.U����KH49�}��lթ6���v��.=�F��]
C�90���ܦ3"�=�l�7%k\ud���-�B�ᦅ&���k9���k0�vi�O����y���8չ.� Hм���^>$
INZ�.�
�B=YUQ�Vz��̡	"����9Ңu3��q؞��NeU(��eV��:�.�^���TyFU�wS�V\J�+��s�PH�!�(������r����C,��bW)�]��=��H#�sK�]t3m��:��LP�C��S��W%N���e"!U(f�EQ���T�Ӆ!�e!�J��I��P3T���L�1"T�NZ��GS�FRX�2�=\<�L�0"��y$d����;��:�W���HĢ*5.�4U�kB:5
J�TT��V�L���"l��'7j�Zi�����+2�����P�e���-"��I2<��IhGi��^�H��As��dTs�S����Q�������\���-v�^��r]Q	"��p�ɪ�JB�.��s��ԫ$�ڔ�]�;S����^�^���y��g�[�s��]ƅ�7ݱ����1I��m�dI�wy�B�]��!������������O5�&��w&��s�d>����Ǆ���:>;�S���/�ܨ|q'�=}?�<�����8 �����E�u�!���7IFƺʬ������'Ѣ!�"$����oHN��x���;���ό~y��]�=��$��r��O'B�7������.	�C��'���97������?�����a[��_������d�<£zyg�7J�&~?����������㽧���I������I�!:v�����7�'�<c��-�'�9ޏ���'㴏��ro�_�'����<[{~���	�����,�-�Dp��b|N��0N����z߾v��yL*��'&������Ϗ>�?'!���a��m�<�N��z�xM!;{߭��5�7;�^�=�w�z�zv��$]r��!K�h�t�.�:�Vz!�>������)����p>=�!�����'���xC�i�C��{y���8���F�Ӽ&�}���M���w���@Y��}��<��rs��~���܇#"$B�r_�z�����a���z"-P��O���yC�a�����]�4��?���O�xv��A�	i��=��ɾ�?���x�7�!�5���ˉ��L.�~��xI�r��~����U_AY�֫�qOV��K��,N_��w�ӹ�y�?��v��Ï�{NC׈��~w!����©�'������_���.��m�y���xM����C�ZM�	����|����&��#>^��}%��B(DHok�2f�����A-����>��}�	�y� /���w�p.����{Mϗ�!���ɽ����S�����ݏ� �U�w�=���Гy�?\~C��|!�����|Dvw���v{�mzF�ܚBC����yW&��s���ޓ'�n�?8?�r������>v���ӏ_ohxNv�y]�������s�Ǿ�����{q��<�|w��?F��1�V�10,(Ji�.��?(�׿O� �7�˹�|��!��������~q����.��r{Cۿ���I�P��O??{���_z?x����4�������94�'�{<q���i���-{�G�~���_1�*ɭ@��i��67,��6C���M$	��Z� ��ϲlێ5|��˽lI�V���,�'{C}���g��t)�*��ɻ�It<9N�������$��(���
�Y�<m��vk�3�wK�Yj!r���`�ʥ�d���_oNC���ǈ���0���}v��Wy���<&���<�ӏ�'�=��!����7�s���ǌ����C��|~C�av�|��O�s��R�q ���7"c}�x�^���:�w���~�{�����&���Ń�C�6>&�P���޾[}q��������po�����So�����>�|w�{<��_���ư�K�����ߦ{�"L���{�ߏ�����Hraov�ro�$<Q����|O	�ͼ�}I�w�ώ���ܚBO>�9���<����0���ǭ��σ��>��I{��;~g{v����|S��!_Z�V�d
/��_���S����?{��D#�����}�	��ϣ�
xM���M!&7��=�%0�PN�S�]��'!�4���}����粘\|qx<��~H��>�</��?;ۤ�>S{u�����U�SN?o�����?�}�Sr�_1���&<����_<{���9��������G;㴒]���,~C�aAO��9���=�Q>c�B$}p
��$@Ov�6�_w�&Hyw'�8?!�0��?����S����[��$|~��_��'��Гϯ޼}v�����~�����y��N'��oi����n@���<�~��>�����<I��|fڣ;^�ؼ>[{w8?�����۹��=����~y��~O)����8�y7��s����x@�I7�$�����o��>����4�,�}��_���dz�� -�V]W]| �,�3O�V�x����������>��<�Aɹ�y�Ǆ]����O��?!�>;{yޯ�����ǟ�x����	�{�{������_s��}L��>��F>� @�ξ�@" �n�fM˚ҹwgZ��B�|!�<!��㓓�@s�;����zC�aq��w�x�������P��ʻ�i�w�}���ɧ�|O�Ǆ�P�������1&������y�89ޒ�}C�>�(G�C���;�^g:�w��~~���';I!�߽��
nBL/���c�I�����x���|Nq�����yL.���z=���O�90��Տ����xC�{q?\H/�xC���Ǥ���Dn����xD�~\&{F������~�>L-�-���)�3�TN��k��������n麗B:���q��9+psGbj�����{��Q�N�Gt�4g�WWTi��w�%�4ww`�n5:�ĮN��X�t�2�v��Mj����7����P���������?E�wُ4�" �!����i��$<u��r��&���m�=x}8$>8��z��'��ﯷτ߿��o�-����nC/�H}(L��刓+;g'3����� �?����?�N<�|I���<;ý�Sri=o�)�]�5���דzC�a~�����I�i�ޏ��"���ǐ�}BO���}o��P�N������AE��N����{Ȯ۵}�z �6��<8?o�;��7�ü'��W!�������_ɿ~�|!�>���㓾���ǇN��'����?��¨y��ߌyNC���~�ǎ��r��5�� ��#�4EL�Lg�����ԕ�\�{����
o������כۃ�G�����>������]������J���z���&��S�|q<��d |E�~�i��O��@�"$G�"g1,��t[��s��.���&�!�>!��x������_[Ņ�I�'�Q�<�ݹ7�'�=��ǅ N�{��<8�O��=�xhzM |}�����"��|���������:>��n�wT ����C�x����y���&:���O�D|::�=D|E�Hө��|�8�,r�zI7������w�`��q�Rw���o���?r���I>�tC�@�<	��q�����}#�ٱ}=Yw}W��^��}�'�\{t�.�~���7�$������7�'��]����ϛ��᝼|��O�}v����O[��0����?���_�z:d>'�9�\z��">�>C��6w�$�Ʒ���d�ĳ���P�L*����9>!�M�������9]�~q��H&�^>��|v������O*�S}��;]|@�:���iӏ���=`9�]�EY�>�}�@��w�|�,x�Y����#��$}>�O������9=v���0��{��!�>���~<��:C�?�￸�3��?�~��&�����&��h�N����*O��E����G�\�>p��(������n�=�C�!������4}�]&������r����<&��A���������Ϥ�S�ra���&��M���������N<y��DE�� c�ӕ"<(}"!�>�~\jc�W��P�OU���������M�Z�ua#6ި�V@h�m���b���W�ᖺ�gM���jz��MVhy[n�0�&^kx����s����1�:�Ԕ��\�J�\�6㴳�+�2�w�&+a�	����3�ңW���RS�ISVq̙x�F�OxSe���=�}g��7;��(raWzO�>F� y:9������sﭾ��]�3�>�x�S~BO�>�~��zW����t�v���pI�?G�����<8�~���]���1��+�mS{E
٣~�.���]*�����ߙ�S�=j2�����x���;�yޣ�}C������q'�=!Ν��r��|���!�ǣ����O�ܛ��=s���#�"�n�#mg�����ۧ�x��{Bw�k���}���ɧN??������z��]��T=u�M�>'8�O^-�P�N�z�~t��y����P�O(s�����i�:
��@}D>��J��oƸ���9��">� ��ʾ���<>�D}�~��q+����xM�	$	�����ۓ��C�����iHx�e7�/�o�<�7�/���=��т C��dy�dQ��~g5�E>�����hyg��������,�O���(�� ������ǟ�~ON���=}�yv�;��7>�y�yC�aWy���n�܇&�~������� �q<��$]��#����G�DC��y9��ro��W�٩羆(�@��f�h��{�QG�!��f(F#>c�/�s¶���D
�̚��Іܺ��^������nG_l
;��h}�����ws��c,�ʄ�[�c#�m��F��-7�� �Ϳ=~(j�yk]/�CT@�����*��������ppT�"%{��P�t~����e󛷑i�Ĳ瞶�{͗k��`_��
���S�!�8|�:1T�:��>������;7��z�Y��S�]o��e���9�r��g�ty�I�~7�n�d���nf�=O'��&v�#۪�p^�6�+�՛�0]Dj��Vw0E�A�C����CzP��Q�(Ò����A��F4d��!T���W�'mH����	�n�V�Iȫ�t�wt�%f��-}-	�g,��$��D����B�꧱��g8PUJ�w���R�ԫ:�p%T�\G9V��u��#��C�ϭ4���$�����%Ӽ�K�����_��%�#��3�z���)ҫ>��N[)�1���S� �����W����=�n��nY�S���d�B-L��#�������!�>e�I�˞Tw,��u 5SW����3�����;V���T�$�����k���k��=�?�/#E(�ׅ��;0��:r��]�Ui1S��J���%�ɞ�v�T��~�ـ��E��O)�����u�/5���E��@����/�(�nY�\f6�BFb�hW�m<8JGv�6��c��j����ÄШ��*�^Q�;�x ���@?�:�K��8Dm\5�Fnr�g=���*�5,�%����Gt�0��&k�o��s7���<`l���<�i.���l[���F��\W:S��.�I
�,?N<�7 t��Ҭ�J��ų�f�T�p9h�V�0���ݼ�?%��_1�Y�R5᎓u�-Տ:��������UrX���t�Bj�?"�g\nb�hi�׀l�K}X��ۥ��$9W�u#$���@�3%`���Cz���z�`[�	�f
��7�����-�͚�G��RWR�[�_klZ��ˡO����QT+����Bnj��E�K8����TC�e��Rh����=%eG�iL|y�º�w��mh�~�bC����X����O�W����S� '���\�W:	no^��U2ql��F��^����.Ӈt9W�m���xv�}���Z�6Y�P2��� z�� =�g՞�0��LH:�������R��	f|�p�X�a�����v��}��"�K��#Y���Y��&��^?�����򆰇t�'�C�b�mB�or�TiU�f�qs�c���3�b�5HF4���:`��M�Ƅ^^\~�X գũ)�]����C{��Ϫ�P��ׇ�į���kGO���q�M���壙,>)ݎG��E�.H���������~Й�>���*k4���u�+���O���y t�$[=�gV���)�-:�_�i�;�.�$}u�
%��ڟ�v�mDp+6�{�UH���5;��iNግ��;v�~���7'��B�P�g�	:n�r�O^!n��t���Mk���f���K��"5�N
�j!=�莀�݊R�ù�� ��6��l�g�i?rQu[9��:�J����А�����hmz�s(��H���2U�͵���f���ة����+��y�9�oC�F�+�d��^��M!P`s���!ڧv�F�@�bv����P�uZ��	'm��w�N�~��__0�<�-+��:[7�UQ����+�J�I����s�Cp%k�8���t���0� �Y��N��2��/���f�LG;����M���h��	�퉇�`~��Շ~dx
ΙYqvz�W!�i
�wy�����&���^�^Zy������^.�|���/aأ��ot�QnvMF!�Dj�4u�-�ȶk���췗g|dG
���dB��a6(���<2�Po���]x��l�)2�b�*��j�Zɍƪ�F�_n1�䏈v��*�I+���6g�F�F��q&���yKS�El7�����_�Ui�����i���P�sZ�'~NB5oO��yG�RI���� d�[�C��}dX�-x.U�+^�����)���gJ��|t�+���ғQ���kku��SV��+�d�0�$�C}�\��aC	�61H�S��������oГ[t��Ե�盞�2�g�*�l<jU�]�#Pc���]g����i}��V�VoZ��4�LZҺ�^��uo��c����4͛��^�b���O��2�J\����������*h�W�U	�X����&�){]�*n7ǜ&DkNc�3r��B��`����o2��9��u���	��%������QDz._f�B�������1���%��)2����"�����츩ѧV)C%e_��� H���>�o;���u���n���}P5��1��~~%.��'$^}���<�}������H��Ng��
)�[��X���,P<y>�h'M�!�qe��ݎ�(�Cu�@2�2Ju�\�ζ�Qr�
��1q�@��H�N�1�:[60F
}0�(�a�x�qT���=P�n�b��@�,��LB�Q�=�#WF*acU�f3N���=<�O���3��hh��:wnJ�F�LUy��kg��T�|��i���Shj��]���������J� �l�:���R���]�� �!�dH�+Ƽ(�y�@v</�k�g�k�2����t6Tu����:�W��*$C��5���[8��֦0�	�-9"�b-��u���fF*�~�NzG����9�Y#&9D��N͞�j�l��?eG����}n�3*K�%ju�Or�(&����f��ZL�ޔ���]Oe_
�^����2k�倌�$�*=^[�6pgE�5�V8s���x�qg�q���<��|]�7y�]�¥�eQU�Ǻ�5�+gT�8"��j&]�}���Ȕ�DkBZO�wP��J�uw\]�6�x��0�Y}AD-���x�d��5X6��s�!�Q�8���������t�f;���Ȁ2�	��C��c�V�|�
^J�۷�厐�nN��8n`��IyJ�[�ݽhc�3�_r	��,�:��;��P�:'F)�4��B��\#D��j��WV�����^��T=�X����9�M��j��<�����Έ�E7N��3����P����ؠ�+�
_v�����7�ggG�����e2-	D޼_=���nt��E �n��˅���0�ܖ#4�R��}��۪��O+���f�|��.o55��\;ɞ0��f�iU��
�u,�v9�!C��֪�����zN����p�Zh��2���(�Rl�B+�Ho���qh��G�p��&�;u)n�s�J��A�=_S��#k����7�H���MC<��԰��s�?v�'r�{7/T���B�+-��t��-��c �5.8J���WQ��Ζ����>��5��[�([o�}o�_Y��C��Z�'ԁI4:S"��f�`(��$[n��S��G�v�E4x��ї��r�9�2��U����4%�v�xҖ����3�ʎW�^�j�]��Qf�%ڢ��5�`��F����=�F�j����+N��\JD�t�0gi/t�ʅL����e���u��c���`��7?�V�t�k����x�)U������n��<�\�M�t�����o"rf9�T�=Н�*eH�
J��ip�N��wyjJ�q]�77J����C�g̀y�ӐL,5ɚ���b���#������T���J�*��lLp�t�t�\�{�:���*!��qXT@��bV�Lc?=5�Pt�r])·��ԡr)�K��D���1�ɺ����X�Qxb.�^���q	C�j�ͯ)�o�׸n��E��sX��,
�&����X�K��)�~��Xaa��c\�2l \�<B�
@�{�o$��^�wQ�^ k�*@�h����\s~��Xn1�}_^N
kҡ�{a���Z\�|x,�v��򈸉�yt�uq��FĔN�M��g������<o�!�c{�6p�ᶻf�O{��*���i���
`mP�g�g�t+��l	6��Q�/���k�������_��.i�CƖc�F5HF*7������Z/NY��P�+�se�Y�B��mǾ������
���Z�9�
���W�W�h�J�����{����9ة;��t ���z���������Q��v#R��`��`EHQ�aۚtI�R����:sj�z��:��fF��uZ�C#2���ǔ��p@�c�&� �u'�mt��w�N����b˥8��P�טDp�4��v��XS�W�%i9N5�0,���Yg���x�ѯZ����mv��Hˡ-��֡�w��#NoN���D����5}����c�����6z;w9Aٺ��	?d�]�t򨫸a<Xᨀ^n�&�OVZ]һ�e1�0��h�h��ʸs�8�X��9`C�х�1Z���9W��e��l�dE��z�ś��UCӨlunʹ����_a�f�޺�rM<�-�}�A�����`𳹰��w���jۈ��V�a01u�6�dk�'vً���B�imŽ7��b�\J���ɸ����V���bZ6�rF���A�XZ�	; 尧�r�W{�֮���
�E��0�pɎ/�i�5� �Fj�����k� �Bps�}=8���w�1��,�|{,aJ�AjtQ�'hPc�Ij��C���X�=������uZ[2���H�R���8z�kM�w[O�d��t����V񾙊�ZLa��w^4LW�Lk �k3s�6/�p�_n;7�N=;��2wf���E����,,�VQ�3K��>t�D_i����enS�Ys�:�î��]�����m���:��4�*����x;)������޽�"à���L�U�xNsE0]�a���s6m^�\�i�����[�s���Զ����яgk��&��$��.��I��y����}� ��N��up�Ge���j�5�C���l��V�s�I�ӗ� ���ƻ9t�[�'M��yM��]�`��Y�_2C����a��Q�f&5�o&h�Kv3i){ۯ���xۧ;M;"��y��E,}��=�K/%�J�Or����N��\ʳT6��{�ɻ�K����.��V6�[� H��D�T���1.e�R��cm�f�h9�L&�-޸��
��y�\�2b��f�*�v1��W���b<,�S�Pmmʜ�)ƹ�0���Xƍ���՛���`U`wr#��3�c 4�i�\��
��F6D���=��T�{�M,���q�2ê����q�[�(Ⱦ�7���=����L4�'��={ٖ"�yˬgN�r�V�2!�"��%�bG��p�qԖj���}��B��bhW@E6v��Uu��m��3Eoc�yY�ix����t��S'�PU��5A�⿇�7��>��d����XpKʿ����iJ4�t�5��h�r�3�c��������O\��̞IG�6�+���Dn�1��[r`�kp����$Ӯ̭.J���c��Y.�+8(2^�D�m�[���k�x��֫ddw�P�Lң�i1��8������=<݄f&����!r���M�Br�ݖ V�'}$�ٜ ܜo#� 'Ə�A$�� E(Xs%&�,������½")	�j�(��L6�I�%EbEzМ���۱wq�i��5L�E���R-T����� �5-���]2L�NI.���G�#d��W�;�^.�9�Q�Um
I$��^b�'u�Z���#��N�z$&eWJB�C�(��u����ft�i�3����aqWKH�R�`�dA�lD�SI��5*Y�ӝ�&MDVA���U7:씍��S��GQQ1�J�Xn�X���'qT�N��<�OQ�Z9�l""�(��.�J���M@-�Nn�i"�����9B�r��3rpt��3��;��E��A�(�E�DFd��3
T�!�R�\��F�Y�tpӚ�b%�,�)8jwnV#(���G�.�Q9i�"UZ$��D͘eFF�f(��wn�^�x��{�*�a��Hsshb�'��D�sY%0�W$"�Y��\�2B�x�z�h�����AE$@��Q��y��;Ycz#g���u����,����yQԇG��[�r�C{�l<�!,����_�q�ֹh���ٯGA�����x��N�g�!�}��Hף#�ƕ
��+�u6��Y�P���vy>�ýe1�M3g_<�_S���y]��f!�VJ�>/�ߪfq�.���.���_�z>��Bxs܋�u}���_�;��w!��Y��.�C�Y*�^kc�O���8t����-�+��o���i�_mo������)�qm����X��ߓ��: �w�����%.w�S���У@'O�0�yҙQ����:y�s1�8&N��.E���t�&;�7�yи6m7)�������ȟ�L1������������ܺ����sڝT��;}�+5��]��RYZ���#�z(��Qx�}�Qݕ�.�]Cء�0�4ک�$���|qQ�e�����H�C5}-1\ �<;]-l||Hu׳�2��)�i�Zx�C>fD ���Bu������ƓB�P��U���{�FwljnQV�:��׹�a���/��[�)e�	�E����������L!d�t)$w�-���|��Ū��\!�iGҗ�(�C��:re3���]���8OR�/fǟ!�-����^��Q#2�9��Y���w��E<���S`]���ce=�ͻ�v�s�z�Gz�@(ۮ��7��ծ��u���f�-�g��Z%^�\�b�@G�G�Xm���Ϛ�л���N����3�{LF����-�b<K4�ŵ�}=����l;�xh�6���4L �`C*&߅ʶ����|E�n��6Vt�
s�i�q:�02'�!�����R�)D��O�:���|��^�U�(���*�����1����P�[���Y����WVUF�����琽r�B��ܘ�_L�f�E
��q'�}��a*��E�Fr��(����'�mu�������'������T��*���,��T��gC%��٬�8���v����]_\j����)�Lh���,b١Y9 ��Xy5^��t,���e�Yz���@=���;��@�^뇟鳃D!�o粄N��Q��3����U���D*�|PA��뮀E�Ph� uD�D�N�0�\�3�D`<P�n��k�{>��m��ġ�D@�\t��y�ÅL1w��W�5)�-�a��7]����=�c=T��mY��~!F�ݗk�ڳ�{M\�����w�q�X�S���OTN��3�˗VTYv(�����9j��~���N؃��V&�Z:�w�S=w�$�7l�v~=���^;�[��A&�ξ�WGb�;/9��ƭ>U��b,�#Z/���Ȼ�ݤ��u\"S����U��4X��{��v�7f�O~��{�v-W.��J�6=���_)ЁY���Hd+ƴT'��H�<]>ց2���K��o7/;�͎��-3L[}V�|�����Rxl���|^߂�C���3�Ve���[:k�du)i)���H�:]�9J�@岉ښ�&,���Xj�5�b81A�ߊ߻N(3Vz���jox*��?�Q�*1����=�����fn�rku����2�A;k�Q�amC�7TŦ�Ѳ�+5muܛ�^�S��K�C=��Ҷ�yq۞vƟ^ہ{m�5� ��kE�����#�u��x��w^G:�0�9�h���E�<��*j#�֊�Pu�?��A��`{��C}���lW9琉t�c��n녛q��� &�j�U��M�/�v�1�a������e&�(qup���j Z�ۧ�g�{<�߽86���"b�w<h��,{P��(h�{�t��t�J��mҚӚ�t����Ϋ ����0���9���V@(<7	�g�}NcE�������qۆe��N�kw>9�+��ea���&Y�P�b�9�4�i��.�`VAw=Cc\�>��tr�|:����$=�aރ7���|뜆�0�y����﬈�ϯ+�:�V�5�\� ������*s�FTH<N�a����}���Uc�����]��=���� +]%�5��e�"�+�>V��`�6-�\�Ӳ:B��<�:{Ui8�����-��D"�� G'��jw#U�'Z$K�n�5���G7�)s�}뙽�z��F�0L'o!���o�$f	�	\Uu�Y�&8;p-Vcc6�H�n��p�]���$s��+�p��uH	�b2��iE����Nӝ������U[|�o�r� f����TBi\Mê�g�,v��@��m9Z��.)v��{�.h���';���|�+��,�[;�Vv93_TF��d�5'�)�3��mf��Ͳ�r��_>�.��%ja�R�9ȏ:�[g�|��/᫆C�����U;��i�#Q�����N�tcr�5��D�9c��MT.����������IU�b�'o�׹�@��{i��)�
a�oX&.!�����b���"�t�߽�q!\�y���w+m�)y^>��j��`U�ნ�['���u���W��I�w2�䥎�̿k�.��=��)��n%����v��yO��o3�����Z-��͉���ouP�L���m|�����1^{����̊
Yj��>-�E�J+/��N�Ye��3G��=����w��E��ͺ2=3Q�V��ꝥ�jl�Υ_�_U}�TD�?q<\�q���k�Wc$�DMIC�Y��~=5ԋNth�Y'LQ,_�!eu>�q��p�k�Gt�Bd�si��kT���<7}ޟh{��JyX�\/��I�W��Z<Q=�f�98����氻ɝs�B1Q����탐岴��c8�͠�e#k��|{6:�s��O�R�GtEn���8�qW����twkt�J-���7%�R�v�bj�t���/_q��5s�{!��]Ѕ{N�M�	����\:[u���WP�-¯�����;f۸���)�8�����%3hS�S:LF����q,�/L�[}9�4��[����|��I�Ä�OD�����Н�1}9E� ������r�[�o
��T�u�Ԣ2��.S_v�������_Si�}H�x}�W��hnfAD���E�֔*
�v��ԁ�xe
4��������|�LTm��C���ӓ�!�-Q� D	�̿m�SZ��@�ѭ�*ދ��S`������Trv�gΩ[��kW��>�k��DӮ	J�U�[����Dե���/O���nrX�糰�zX�]�����kw�� 
j����۩婣��
kH���*��(��q�<kc�OJ�`�x�}���,ھު��Ik���}q�K��o�JW諭���,%wo;��K	f~��Uη�)9��&��;d>&����A���̱��]�	�ޚw�y�7�.X�"���������`:��#�}��}��G]��a��,E���${*q*�uf�η��.\r�-�4��2#�j@{�v�1����Pܳ69��h�k��}�v�K�g�B�����K��3���0�h�n�+�e��N&�*o����z�E[�yR3��^�f�cׇ�=~��<��0�ו{ٯ�%28�7�"NN��*�)829��Wt�f Ǔ�+�\��o�!�Q������������Wʱ���i�O[}\:��ۇ}���VV~OC�����$~7*�p��vxJ������;�m�7ެ�Ad�T�6Euw��)}��o��[��p���p8(�=��L���E��7S��o
=moڦ�a���	�,Ggr��"5L1����u��ɟz���G���(.;+�3W�{h��7���ŲB��#*���]Q����c�"�1����h#�Df�z,d/Yͫ�~����T�qʖގ�q����6�8dm�-��YY�m\0��욊s��p]�^��k2�{��s�ƟfNHm����iB�<��.����ݸ*�Ȃ�u��!��DN�|	Z���<,�M��t[�L���#Q_���舂�%b�r�&���>���4����2��ƣ�뇐
e��F���>e��v� o$궭�si�r�qfцz��#��O��˅Qp��� uA\tMD$�#�ARf&��L�[�իZ�t荿��rP�" p��KYuD�ٳ�����9�!v�]sӓ������T�D�G�ԯ��qo���*$;�E�B����B��jR
Y�+��0j���sڞY�WN>�nTЎ�pp=iހ��ā�,G��\r$auS�}+q���X��,+�f�tt[1�v�n��18)��g>r��,�=w��Ek�45`q0��ڽ����yp�B�9�j�MF��ѾS+���Ѣ�H�uU�.�I���:�}Ik�H��`�iow+�&�׆z���t꼯�\�3Y(i���A�b}����}QD�|�5���+%�KJ�CRQ~��͘4PG�i�\<*�쨬1W��1����C�^�Z ��	�h�������R���q�yV&��:b�{M�Z-�u���< ����@W��'��铏OUcHv:����2^ʰ��/XxgV���z}�)Ζ��3�*~�δ��ط�n/&*6�v�}F��ǂ��z}����!��Q��]����	WF�/]��L��Z����h��co���﯇^�X����`8��II�:4N�g���ü�_�{��N�MR':;�}};in���VX:-l�W=� g�le}���؛�Z+��Ix_*�������{��x�wZ�����T�#c9�&���7|#�����r��� s�Pw�~z����J��ֶ�cJ����YP9�*f/>\���s-�L��P�Oz��]�4T�N<�U�IQÈ&���t�w	F�0_j�
Χ)��Ź�'f��"������x���<�!Yw�o՛ C���&�"�d������h�����X|��D����<V������o��{B�)K��'�R?mP������V%s�\NY�չ%=�ɝBCT��p��8�9�v�Ϻu�����vtoY�wϬ��ᜌ5VV��U��'5+1¹���:���)S�㐟R=$`؀�L��雅��cDBDF�5����֮�ծ�����Wa��
~a�֍��:�͹��V|� "b�H��zT��c"������
��v��8C��Ѵx|b%���3�@�gy3_T7�[��\��[@uC��z�;l�6/nŘ��za�5FɨTI3p�[�ђA��YK��q��|��V,��Uܷ�=^��.�vs�+��o��*�yJT�c�;���N�yp�Y���flQ�[�d�OZa.̖���z�׹w�+��L��*����"wy�n8|�Z���4ј�9M�l���a�c1V���<��}�<�P�f�/
�J�g�5��������	���*���Oa����M�m�Fe���09҃R5K�N����ʭtNç��%6GLTsT	�w?8W$��T��N��b�0��	���^��=ݩ��M��}(1p�o���{�\����W�%�?���3�=�Af��*�˻cN�߷�Lſx̥{H�;;�����u�Ϲ�0�fF}�eڽ�r��{bT�;��{uTzR�����u�KY���rU1T�5�z����l�b��s��vD�n��\���,����L�L'h���V�F�eCЛ�R�.~��;`�c���Uٙ�@��<��Kؽ<�{M=E.?��Ѻ�Z���QW��J���5�c��M�x3F'���y�]ȶ�}��opv�⧺�-����8|���U '��Q�W_7�F������gTv߼`�}��l!�zX�x�{�Zr�ܬ�
�F1*�H���奧N�V�ח2�������
/gT�K<1�o$[��v�L�]�{���i��̺K�S��1�<��+�b���K#H����h�|mbwۜl�=1�qx���8>�ki��A�aYÉ��<���"2f��D�sl�؃"�}��U��O�׽�����[��]���܍�>B���8Nc�|�K�+����C����B�U�v����d���绠a�9?O�q`�Tk�ޘV16�`J��[��"Y�����/���z���O=^�=\�N�o�ON����D��C@"�3]ϖ@��D�N�3p�cDp�S�����4�������t�m�;��9zf�]��R��축\��Ӌ�z�x�ߜ�!u����j����"�_PӋ&���3|�V���uS��:I�6�c��ҧ�Q"�K�<ʻ�V=/����^'7�1�����j�*C����>���R^Ӓ�u�k,�{��j (b���d����u%��9��hh���6T��N݆ � cBO��Cr�51�{�ä �t�k�2O@/x{�چ�ހ� ��u	�Kr���"����ؾ�T���r?eco����.���v�AY��B��X��l�({ftDuu;��Mk(���#��� �=ަvo����{l�2#��j�p�-[�r���(n���)���6gJ��W�]B���N^Z�ʽBD=��VT5���k f-b��h���K��\�w�0�1|����w���ܝf�=nsc�J����(�h�7��Y��u'c�z�!���I�8�[[��$n6f�2�m�L�]�KJ(R����D�cݼd	\��4w&���c85w��j��S��l�Bѽ�̙`.��Â��{��*�I5i���Z��8鳹 ]�í���A���{k ˡ��.XD����/��s2�c�bJ{�C��s��q֕�WI�Od�� 2Γr�0�n�l �G����οe�%��n��/s�K�ţ�ࡂ�<Ë'I�lut;��7a.<�{`�ޭP�t�3�F�f��wR���T�6�����N��W�6KWQP��0Vp|�hcj��e��8ApӜ;VOvQ����ޘ�Dt�[�n�ON�ݶ����d�ɬ��#p���!��x2ЦK���}�3��gD�T�:�,��K(�C{�KۭǑ'�Q�Zow���w-m�,��|�q�e]���B*���,�v�U��M�R޲uU�`�w#{Ӻ\k\��q�������]����� f$��2��[��G��Ztw����y��d6�L���s�v�� \�h�N�\p�����讘_}�H��u�n�Q��ȩ H����<�q�}r�oX%���P�
��y��B��!�P�>[H��\*cL��޽���"�Ë2���8̩�f#�	�R�Ȯ]O�X��Wsnh�u��4G9.N��\�]��u�O����{���挥嬫U	X�y��(�u�������v��O:��b�F"�[ q��\l�-=�����){�G��6���<ו�W��ײ��3ƪ��6�l��ff��,cu�J���x��r��1�,µ����X�X��[�%V��>y�ܺ�QW[�ck@V,�hL]��bW<�I^�IU��l�r��[7Q
2��sE�)����Xܫ���� �uJBl�cC&��5�s�h�#dѪ��D�*�����';�Ws	�7�7�b��|�i���R"�t&T�5q�̩����CEe��Q�z�a���8)m����J1��ջr��O8�+�ol��65�T�sF��Ցq�\��C�dp/D@95n��6sJUZ=vm>�����9SH�u3�7Ӣ���/
sw6J��Z��Ϯ���&2�8c㴣 �i0�i�-����l|Ӭ��U{
�Uݕ�r/�kcc��@��e�NR��e�v�SaZ���B���y�@T5��Ɍ��������Ӯ�ǛO�7�v��{�J��5΅��f�'�[)�� �6����*_?�_����U=S @� �� ���a*)f.a^l������Ԥ��5J���W9�FJF'D%4�u٘�b�H�Dm	%JD�: x�i�U����\+�\�B��šf!IF��f��衅J�,*жBjH��9A��湛��B�J�4B�VD�bdl͒I΅F��Y����;����lȌ�%PM��X���Q˙Y��J�B'Zt0�1J:�r�FI任��B����ȐӨUA���a.��ɑ�)+3��G,ȽhN��"ʊ+u�쨼��*�N�����Lr\K+M+YF�iP�w��7=0�T�Jf��QE"�7:�P��4$����T��Pe�̲�*�fH�J縂(�b�wqu���G6�J"���-�e���swGJL�,S�j!${�̛�:��Q3]Ȭ-,ܗR����6$���9���F� U
MJ�v۵��h�"��,�N"a��6�;�"�;5>�؟RZ�B��ټ��%pW2�.[�V�³�F-����׼����x���G���&?����_i�گv]� 𩸫�Q;<%ZU���@_�Yגp��I�*V�f]h�Θ�+�r��G���݌��<Q��
C�B|�E0��"(k�������o��/�2�;�f�Ξ��B��*��^��o)--�%�"ln}��|�v����@e\�k;=���^��-������.�8]j�Eg�g���HUM[�u�g+��.��7%�b�CQg�VP�x�}P�N�84B��{(E�����VXn���1�tl���mP��d-�y��D�,f�?D8�l(��&|��en�U�#V7��5������+�!�����;���	�,U;V��=8T��XFP���2�(��]5^_�9C>�jT:M}�X@��A�!t�VT�����
4�yw��d���k�EM�O඘y���M��cw�8˨���E��� -2���M���ǥ�s�>�^��^��z�7*�I��p�U��]�X�<6E}}�E�pR�����,�1�sU��ȧ��E�oTȵV�c�*�j,�F,�M�2�!���ce��P;F#|�Rj35^��PgYחނ@޷�a�����]+C���U��_

��h�����,��Lk��]$����DR`�m���3�juca�ع`�-�KN%K��W��}V;�h\���*�z�'�l�s�a�>fV���2㓳e������3M�n�ő�ʓۼm�4�}O�ep��5�s��S��):�\=;�w���ƳY؄�e�/��%ϫڶ�c�8ɮW�V��%��R�[P�F�2����SQ��;�qu�W�nڪwn]a����j�Ӫ��A��6��z!.W��X)�[B?j��5��T_C�W˃g��oJڽN�@�z�PX��oiΰmƽ����+�Z+��D��VU}b��k��ˊ��5h�v;��R�p5�5_T�"��'�!ogr;���27B�=GM��ۥ���$�wk�?=�_Xҥ�AV;��,�#V\FĪ��\���a��,Fi���4@f��ͦd�˸��ޫ=���4L����o�� ڔa��s5֯��N[)�=Ua�x��}#�ŵ/l���^�|!�e�CS�2PS����<���Q������Vo6��%�1os%b�-]���9|n%c���8!�Q*����U!�4�b)��0n]�%}��ztrΞ��9V�j��]n��:7�,7�Y�#zq?N��n�B>�,Y�j� ���6t��P������M��`�WMb�����ZN�=��S�F�Q��۝׃jY�Q1H%�S���;����y�FӑJuU������.g���GE�b~x{�&ۂ>���w G�[Ԅ��m��;g��9�2S����S��2N@J꺌����E�5�g[os=cS����C]N����ϸ�����H�P)�ܳP�ƫW.���$�b�̞uZ�#/�M�}�)}_0�U��9�s����@�L�9�����o]>�S�B��N�s,1�	�~L�z�v�O��a)���_�/�3��%ʄ������V�5�>܀M��ӅW��k�?<+!�q�7Xe�|;lQ�r�p�$�7��a{����:�j;��v�/��)��A��Wb<ڌ
�X�0�B�����5Yx�e�p�\� WLgɺ�s���YDO�[f#�rR���Wf�= ��ctp�<��wk^��iE#�xq68�Pc���G�����������.ә�#��ڣ6H�I,|�tj-����cF���� TgN"�u#���|�Ȩ��lQ�0~����o6y�"@�xe ����k5�=��U/����vɼ1|wS��W�ol9U؁�{vJ��Z͆�������\3��=ePN��N]����vn�	A�ռ��્MF�_����̫��I��z7���}8�v�m��w*-�X��:5�Wi�`��k�ՊR�_=�t�^q��tk�'E�<< �e\�5��;��Պ���df�Z�CGG�D�����1q�#�l��-w<`�{s�W��EB�ڻ�U�ٳ�P���U�=�8e
��K����E^J����kB�
'�Fmh��O+ދ��Q�_�:W�7M߭�D�����g댃
��N���� ��{i���:����\v�m�L�N�Ӄ]F����a����;�4b_hR^(�=�㼥]s��[6��|�8���2��ڈ�1I��ςu=ǴF��1GNQE:�A��9�+��۹��`
e�K	�^�gɕ�5��Z�jE��&@��9�X,�)U7p��'f�\�V���ΰK���@�P�@)_4\#])��~^��a��O��R�V׳NOOf��N������~ˈ9�� N�Z1ҥ[����*�>��jP���^�K==Aے�M�:Ӗ �u�yc攪���7Jq^D���G�?��4�k�1�\�"GZ��ۼ�Y��9�t��$E��[9�A��,����LWq3�8Z���(�+]�)�a�\�gi��u�=s�Aq,�j��fL�*#��͓`��mt�N�ܙ8��6~Z.�����������mn*��l��fd�2���\�Gj�����,7��t���z�Գ}ٜwN�2vB���9��5tW�By��2;�=�c#���λ�������3��]��Oކ�ɨ͞����Q	Y�.8ȆN�@=���H�E }�4���c�b�.�r�WM���͇��7j����4A�	��e��d��!*˸m��Ctf��Nk3��R鑜g�0�\ς�)����c��<S�<?jS^:�[<����pp��t���B����D�ۃ�Ib��^���Y���\�u��ͺ���/��)U��Tc�K��[~�����y��j]yL0;
{\y�?��N���G�M�\"�'g����_�wxFt���ƌ��*�������n_��8:�����]e���H���x=���O�|��c��p�߾�Ǝ�.��Tcms��>���r�����\7��vl��-�KM��n�*�֠�"�Q[��(��z[u�3_l��>�ks�q������]�8	�J�,�����>q+rlg��H�΁�2�����VA�ƣ��	�e��v�`���dѝH.ˌ3�&�-v�]z��߆IE/�@��w@"��A��@�+����[��ȝ:�Ҷ,:��������O�R��t5Wz����启M-|��S(8�gW���*g:����ʝ�P^�R'���C�����D�t3�.�]Ð�]��w^�B����VV�Y��ܫ�5d�V��p�V��� ��u�=����Č{�T���h���	��%qFU3�@�z��L18s�ŧL{�u3�d���g�ο��8%��u�+}�_�6��\����]���Q1�$Ud�X��V]�I.HWN#aK�:H��J�E����\=܉e���;��q$�.�]̴��Z��V���i�7nT!�7�Urm�B�������H�y��۞ְ-248-�|kv��
i�Ŏj7��r�z��MC�s�T5�/�t�-�c5[��>A^�}�i�D^b���\�)ޝ�@GPS's�F�'����rU��&v��k���X��*�+�b{y��'+���)�
�]69m�fWc�8�g��:q���c�6�����-��R9lr�dt��E��;�E�l:�lkX�(�yQ���h���n�y�u������-������G��g����E�[�����>�ϖ]��iL��6�L-�\���� ��*Zo���ۤNVCגh��Q���:P�٢��*�2T�� 䭒߽V�UƝ1����R���G{��x���j�]N�N�c��ܩ�DfJ���з��ú����zS��ɔ4fݜ]��8m�z#��#���s6S]
��)_K�8�-�*����sx�9<�kk��˲^�
T��L�rsx���<ȕ"����'y<�6U+�by<�ۣL<�Y9ö�w��v��:q�AgF���W6+����ų�F'Mg>�kT�cy��שvCy5*��c��)����� ��۞�z�Ή��ʵ����N�o\r�I�߹���|;u�N��㌫���=G�rh�z�5�{v�� �t�&�7:iw�/�'�676��0ܳ������L{\�)�n�n���|�z�]�N�4�9�w3�:�OaFnR����AC���Ϧ�Ê�4Q�ʃ�W	[��̎��c�rʋ���-y';ɽ��S��\�%��9�y�_�������H�}���{�T�d�:�Ļ�+����7X1׿�Q�^g�Z3�;�I�|��M�{�d���P>SX��mn&����z���;�[{�R��6o#$��`�]sg
��K�W}g�C������֞{9e{C/ݺ^���E��Fb�����b��"!N�B����3A*4F^�s�2���Tz"#��>�}�
�/S��}�U}mYw�������&!�tV�|s�^�փ�7��Ƥ|��ӆ�֭r�Lw[w�9����;�Ջ|R��7��s�Ϣ�����6y=A���9�b��0�S��ս����Nsr3 �K�p�w;Γ2߾)\f�x�^�Gڣ麺�������Q��b��\Cuy����=�BK��[�r��vڬ�!r!{~]S��>T���*n]�F%��1��.�|�����<x�9sh��hq���5���އ�4s�m�m�#�=-���>��=���M5�M�U�Y���=0^�T^ͱ6�G%����W��SK��.=�;��Q��\@����ڛΎ���Y��Wfl��0_π����5I���*/�ˌQ�i�w�4�����t�`J{կ*�<���d��p#T�_��#7����;����y>-�h\T#$��b^d�S�p�JV��pqAD�2RLT_%�9r��x�MMl1��XA���ݍ��v�u9`��ǆ-�[���8�I����94�Y�s�F��siA+�{��-`Z�v.��j��5t��Q���h���h$�>��꯫���3�QS���cj�1b�	J鐟]�]�}���D�ܜΙ�k;�/v�@�g�1��)B�1θ\�yq�bB;f������=	�4�3���v�s,�v��)1�J�4���Yղ�oP)^q�o̿�uwg���	Q䓣��CW� ��@i�_evDުs�զ'6���/���n*��1��j{Qʃ��#���>D��|n�m�V�~K������1��wg|=�g��]�y��>v�>���յJ68gبs���t.3c�5��m̿�ߕ���l��{~+���u:0�زK�uN�ԆWR��5GO��M|���ܢ�m�N)�}�iu/Q�$�5(<� ǰ�6�3��o��������x�G��m���fC�{E��n�{�b�m�m��:9(��}�K�^��8��Q��w7م�S�Ϭv�}��d�ȡ9{����a(r�W��R��2+�	i��T�jҷp-�� #X.�i��ma��o�83�+x%�L�����#�7�am^�y����٥� ��y&ݺXԨIx6��}��9��wt{��a;9�B��ySw�⢟���>��"'��8.�5���T�c߬�w*��7����"5�_�o��+b�����ui+����S�gZ��vO=+WO.1��)�s��N�::�9�!i�˧�Ln��9�%A����"Ҳ�>u_v�{CJ{�y��ۙ�խ����FrV��hK��F�I#�o��'��xT=Fm뢗���"��m ������ܮ����W�*���}�Y2����MED�~D����O?���u��ٳ�ԛ��Un��JQ��h�>�����u�u����Թ�XO2�ru	����3�:�=�O0�,�q��c�m,����v����nLW	{����YI3�ڦ���
Twk���������l.G�(u�h�+r���Wo�ϗ/f��v^����b�iy�K�[�׃g�V�_a6��Zae��F�T^b����`3ɘ�prщW;g^c��@���71,�%4���P*�o���a�:�{�BL���-4M`.�M�� f��n&O/���ғ�C�u�P��gR/U���jDw	����P��뛤!�%���Mb�tUw��)r6j��tںR��ꋲ0��hwփ/y��!�b��Y0�F��t�oZ��N�]�#3MFyr�:�|�J�ӨV�E[T/V5-��b:Y{+�d�x��̏�����r�n��G�U.a3���ˁʔ�YvCWz,�톴t���=����*�\�*At�#H�Ef�祽�4�zұ��9mǅv�e8	td�r,�Zd�b�ާ�R�]+���?wP\��g��#{6>М3f��^8�YXdy���Q8�3!�[;���Q#r@i�Ʋ�}�.\�0TY��e�W�1���2�jS[�|�lu��FDl���Jܽm�X6�Z+Kr�(����-�]m�S����qu�����cǻnofi�N�W
�u��}3�)w�!��'%b޺�����������2�3/U��W,��-�hĶ���S���k;R���omh3h�����x�K�uō�af����|�qhĨ�ݮ̀J))�>�`�U�t�v��M?�tՒ�V�*�@�eȭ�$�>�Zw�QͻK�S�t̭���O�wjl	��Z��j�q:�!�6���@��1�(��T�3,���4�t�@Jde��c��K6�ݪ��]���\��i��*����Ua��6�Eŉ��Z0M�yW���eC�hLS����p�$�A��6 �n�R�R��m�%��4�/8��nn���X��j$�<�a�~�hhbJ�-'��#�(�;o��K:e�z&o!�{&�Pr��K�u�+�s@EVr����,NSU�egk�D����u9�˴�9;D�:m�Mc�"���u�C�X�mm�f��E�����$���"@�;��ōw�v_q�:#w���IS��u�m��m���]����f���uc8[�DbNq�y6E�Ds�vx����lڜ�v�r�@e�dH��:���Wl,�oiLBc��b�8ͽ�9o���_�S��}�Z]�z8�~+7t�	zDڣ���ei�M��Z��4��oN�_>�I�;al+y�U�-�[l�>�Z�՗W}y��PZ�(�V�y�WjGpHd����V�Y�c f���!��s��l
Ǒ.��LY[а�-�ۛ뾢�!p�^w);	ۦ�г��Hȷ0U�p���4���t�$�Vm\�N�
�����0��Qp���z#���c�4o�V���.��gJ�6��_:{�\�-\�p_=�qk�z�s}�f�͢�xVaK���L�[�f��*7����T�����\�ket��l��p��w��f=��gU��#+
n�ܫ(�[�����'�|�lc���h�v�˳X�#���e�U����w���|Ƨ�c���a�2�S}\���<��翞����JYU�)t",�1Gw+��*�LÙ�Es/"�S��jqS2Us��H��B��ᲉNE��*�S<�
)Ԍ��yy:�I%���d^��S+��;����!�^��{.N��w
�tI �K�d��P�B�g9�R���M-#�)Z���:';�Ni�]Ք��t)*����i�T��N`�!2�����8��jS�D^)!I��q;�aUIԊ�G���'��8�&�.!f!(����g�$��B�NS����z�a�E�)�I�<��R��qu��y���1'\qNF�uJ�f�i��#�qa��Yb��Nl�u�,����"�aYQE��2K��<�yR�U9�ZBT��z���y�J�=�M!7w�+�Vt�dV�9�N��^Z�$����\����]��hG����3D4$un&�$�$�:x�L�'"�'r/0t��+�!&�L4d�P>(�kx�鞝�D�K�#mvn�t���u�B�.�*�-�cf�f�O�4Px��2�N�8nnF�;��Fi��8C������w7���{P=�K�uF�P:�˅��vTN��AX�/=%_��m�h�<^��T���/�zZ��ۃ�6|�Ѿg�.)+�L/i�������r(|{y@}K�M���7�}�c�����(rKkܭ�~�>W4W�����'�Q�Ϟ��O;|ԍ��W����y�FE��֪E(��>o���g��A�6z�A���UM|�?�z�[�*�{��/w��f���ua������$��w!�B`����C�~�|�FO:��KN��,>Jr��4����y��y�&���աv@�;�%A�ݥT�uMW1������}]�'�7��kW�Gv��*j�L-P���X��z�MtV��l������s�)=5ΚY	��{��:����G!w}�L�T�Z�q�G}
s�o}[Tc�^A���jħܞpJ���t�GE��<v]��t��͐s����T��bg&�K��]��OE�Mm�P��U:p���L+H�L[�urF\h=�R�i,�Qk��tp�u���9�D�w�d��L*qC�=�4�.�Du4��)��t��U������=����gFE�_������k��kc���ߠGvюS]0��@]�p;���!���f�&�6�Yo�m^��nz�l&.�F�ϓި0��\J��N�G,�L�WW�L����k��Ĝ}�9S���J�t�'�[~��?bǩZ� MΦ�\��y��J�����h��T>��:�=@Zlv_�_h��y�T���#+7�ڧ]�������$��뜎M@���,�YnQ���*C��*�t~�S�ϝ�.�_^=נ�Z���n�y�Qp�d�����*l��;�w;�Ըe��hP��ϊ.�Mu�K���㜉ý�q�.q�Қ���-�譳C�ڠ��SO��}Oƪz�Q����н�ļzi��[�y���>J[��i�m�d�]�/m.��3��ka[�Bi^nк���m�$*-�۔�i5����o�ܚ8��Ρ�k�G���H��U�ԚF�1K�o��FϬz�K�/d"��b�\�T��Ws��ʹR���^�:e&:9���e���l^Õ}�Vھ����NN	d�C����jn9K�}Vجt!$0�����Ir��U��<�PR�����-���oL�rS�꯾���>�{�9�w�I����]ux�T&��ox�Źu���z`��4����gd�~%zsu��Y��ƖG[+U�����qݩ�
��q��^&��;7�z��/U����bS�W�e⎘���qM���]��b�4B��;�[77Z��ӣie8ɍUjFBU.h���nl��ڋ���W�`���+{oɵ61��2b�����J~��T<g�3�=��ҏ�9��u���T(�f�D]���/���"3{8V���W9��bV�n�iM�Om���M�c�kU�u8i�=N��f��u|���,��t_d���z��U$�-�>�.����-�5�v��J��N��*%9�]�i�����f�[Z�2���[Y���^gU�3��ڵ�R_B7�	�|��Z��[>��Q�6�7�q`y��{r��:��U�uh7I����9
	���ź'H�6�D��c�F-⾅��\p�<z��b�k�7>����;�P�U(N��,��+l'g�#H
�3R6�gS��t�_k�j9-��׊�cK����'6C��UÎі1�09N!�\�J�G��:��ss�+K�vժܗD��<�ZfLݛG���u~�ꪯ��[:��n~�Mo�U�e�	X�Z���/���s���FP�<rՄ��Q���#�;7��Hgj��zj��k}�mh�[Aq!G��(cfP޺S�^n�yꞎ�T��N�||c�]�����V�ܭ����8�.߰�)u�n��:�w��q�Q���R�.�����eG���ܓ����,�����ڎ��.ݪugY|�eV�˛یm�Ȧ��*�+�3�XR�r��4��^�'m�:(>�R�εVy+�:��Z�jy�&���S/$���[��9(�c��ݱ��|���z5Ԩ1)1W�Z���6�&or�-��˙�Ğ1ݫVMh���tdf���.k����=��f���w���6�p�Z�p�D9�,��#�ؖOO��b�#;���W=T�v��c9��&��F���_��=�݉�R�\�����t��`;�m�i �/>|�/cT����2'��R�0��3�ܸ����.Ypz�Ö�(^��ieˌNK��m��4�%٦<(nk��nl����.��Ա�K%Ytf>{���;p�V�.�2�݄L�u�ʋ ކ,9[����%^>2fF/�< D�K6]-�y�`���mߢ'P�ZԪlgJ:Q�*s���e����B&���c�~�ҷ'̎W�Ͷ�|kë�4O&��`|�d�䟃u��_2ͩ�b�P�.�ջ���ͯ9fn\`v�;&���[��h'�Ж|�rj Zae�}���y���X�������]����Mz^���xzU�����g���:-�I���2�,�&�Ʈ�sn���T�BH��޴���rz�)�A���fk~_K3e���=
��k������c�u�'��Qݱ[|���A�sV�v�Co;��]7��Y���9�Go��uu.|<��cbݭ�oT�]L�ssUs\�K泦��v�O0-�7cO<��Vq��n9W�Ue��P�=�c}�;�-s^�X��g���k���A邸mJ�Z�Y��'�Ɏ|��Z�u�c�qN�M,e8Aya]��'5
;1�6��Y�dd�2����>��ۋ�W�b�F�Ugxp�b��
��5�mp�\hΆ�����t�W��*P	A�[l���v;�힢@�B:=PΘ)�%�5q�]�`�x�?�}_W�k'>�i>��o�ΊO�Ϡ��AF�����Bu�þ�*\��7�k'!�mpM��*��֯+q�ڨi�j����M�AV�5B��ޮ�K�+t�	9�z^!'��U����F�tt�zk�m+�÷m�:�{ǙX�ĥ�^ɞ+35��6����vf s뿂�x�J/xb}��y�_�F�UF��JW�@��և���I����u@��0�p��{�x'��Iw�&��7Є���}���ï��f��˶���\�̸��e�9g���aFb��SY��hdѧ�ѯ�L�B����'�V���h�ڋa�vK�g��L�?Z$�{���i���[�����>�9�+�:���4�屻o��=h^�e����'�ᔢ����$�]�8���H�
������NgN{������CMgr;=A��K���k�g-D��m�9
1��;�p��uL��U���\�v��ܶ���,�$�����6������s��!�(�WZ�<�v��0X^xI���zJ����u�͙��1s�Z�n3Sz����yYϳe>'-jؔ�9��pn+���T��Ȱ��Dko
�9�դ��ԴK1B�}�N8���J��ȟC�6�ʃ��-���	���Ң�o=hZ��خM�+�����#]�m�]���|V�\t�G�uu/m>�:�rX����s�6��h>����}��7��^���,��nDO9��Uq�l�<Ň��r���F���c��b��yt��8���r_m��\�xH��ӻ��&�S�Cꌞ���e�m�Ȧ��*�-��!�3�ю�׏��T��}���Y%��+���j����Ի!���z��P�]֫eJ�x��<���N����:yR�dK�)p�j�F����M+����]���ctؔ����W��m��+����6�W���nt��*P`�ݙ��(NT�k��S���h���2�D7,���Ϯ����e��5}9���ًO�6��|����)�v�h�ƪ��bb)!�m��+IF����0�|����8L��{�[>/˵�'n�D��U
������m7�Ew<R�{'r�֣��N�2&fN���=Y���V[Y>���bm�n���Ў4�e���5���	u��ݫݛѤ��+�L�w��[��p27�p��d���9��\�'��R�ՙas�Mm9�w�f��Ve|�<�鸇6$�ʯ�v�z���;ˆ��N�M���%F�'M�yNC�����Z��!�{W�2V�����ෂwr�[�8��Dj{W�ødt��CdMA0���֤��8�z���+���ѻ��vΎj�r���W��`�5�YlNU��%�if���=|��w�Nr���6��;��+�>YG�_���^�]K��;�jmd��yU3mi�6�t8�kN7�o~/��+����FO�ŋ����Μg��K��5;��vk����V����?۸m��TV�!X|F�/S�����4�˨���-�/���tj�s�����11G�I`\;}�[���M��nmgL�3x�[{,��;K��i�(��ؾM�P���k�7!t���ͅ���5*N��αvt޴��|"�w�\���$w}�]=&�4PbQl�Tx������T��3n�����ΰz��ހ� 5�P뵦0�S#�ӛ@����M^�O�����]+*��
�o��M�r�FY��0]�`�C8%�è:.�����6��!N]ZV�ۋ;�}U�Գ\�g�5��~��3˴���to�T�'��92Q}�uӄ�EYN�֜̓��.�3ϛ���;h�Nゾ���v[�7�#�߽mG�"x���TRӵ�МR�)4���w'���t���)�%:@빸�~;rC�y����w�M�����։�|��zÄ������W�8�ʫr��T��
��*�����2��ٗ�N�KY�|�p��W�(���Kx��^Az7�w���SL?���^[?S"V��'���$˨m�3�2��̻ʩ���2UR��
rtd�4Qk*-���O,s����k���&����'��oP��C�M�����W���Ɵ^Zؼd^��s٭�ɷ����Y:vg6������n[����j��P�.����d���F= �}}x�Jr��`�Z����Z5ƨ�ti�P����y7�15�tn�G$'63��z��uй̜vfv�9u
>g�*c1�i
e��XxU`M]�@��!1�����6�vhN(њ��IY�R���v�yN��};���J��wy�.�2�GuQзev-y��zK�j�	��3��lrq�5.�t�&n�K�W���kg^�l�
Z���m�u?�����58�����q8fBy)�"5�����K�FMp�p|T9�o��uu.�}�j{׾ؕ�9J6��P�$�)k��7;���^��ו������U��=[�9KR���`�|�z��y%�ԟ�?9����<Н(�X����y�d�sv����hӚݬ���ᜲ�M��M�|U�Uƨ]Y�F��)�ǩ��NRy��Td��VzI�[�)�hk�zm�Lm�n�����ȷ�Zqߖ[ǒڦ�j�rrJ�*���)�si>��FO��dΙ��"����-��q��	d��/�f���"��n��36R����~��筟r���}D���p�W^�0��L-u�ٖ9:�4�`W�IK����qV��}#mc�0��B�ic"9v�N~��~�[�a<��8��SI�M.ʱ���1X��۫��B�����wx�2��Z�W�j�S�f��ιxpwP*�J֨[�8t�����SQu������*������,�*�Ř�2��aÔ#�d����e���ܗ�����L
j�J��l����R���2C9��u�o"�wQg^�*�g|@�9]�<�Nb�����L�R���NGo:Ж9$�WV�@[o]wGE.��دY�E�.U�Ńbc$��5/Тֻ.�[�B����'���9�Ր��7�P�������ށ&{����I�l���W����T���c��D�r�C�s&�=��ˌ�f���B��ᚄ]�©�v��0�%��X�q����e�-�=�=z;���pUû�U4��h��Q�c1�Q��!��U�+\-
vV=�
�L�K�֭��/���vj����c!Ĭ�}���Pڀ�O(�[�Q7�Y�|z������ig,��3L�*�Yilxsy[��#ɫ*";m����S�|c�W�C{��򩃅挠]��1�PONe�偭��;oqkC���ID�]�VRZ� f�aZ����Vr�X��_�$��|+ٯVgbe��m�f���KWݝ�9.�@�+�sL ��o1�-�����y̢�[�*Ou�P��ۘ���o-�_,���ۭlc�x�k��*g �m��ZVR"��h�����1*Y�(%���kpD�H�؄�c4�j��;��A}y[t���橕��WJX��}�$e�n��L�nK�)�k7��-��)���2��+q��O�2���K���U�� ��,�Y*0^2u���n7��q�f]<7}](u���}��<$=}RrI�#`v>�&ӗ�)��ohk#8�ХwS�`mbs�%�}�L%���s	��b-we��+��c����,9Q����[rRH���ur�x�>�s��ҵ*w^IW�x�<Gݬ\.��D�v���4m��������`�*��<r�0K祉������-t�Ѽ�$Ik{���K���$�Ҫ�u�N��*ׁ���W|uX"��%KĄg�S.��u�I�S�[�'V������.�av;=o�B�G��f�5�g�A�c�UW;�ށ�6˼'��-Vj'JhY�N �p�\t
�t��~ӏcj���I09Ln�uF6
�V��ƾ�h�wB�ůl�n�7�� T��������Q�2��>f>3/e9W1,ț�s�9����-���la;!�of�v/�� ���-�q�u�1�Ք9�H��t�S[�s��-;�A���9��[I%6��A�db��V㳹;,ؤ�E؍�)<k��.�������8yӒ+Cn�w�.�hU��*�`z�҇k�u�:���  't��\z�?f�q���I�T��u�ݗ��qjݡƗ|��G��=Lۺ�M6J����j��%o]��!�p��
��j�6��s�d���f�dډ%
>�H��G8Y T�G5��4K���⦲D��	ڛ2N%�E9�� �������$D\�U#�b,����su"�VD&�Qډ�"���IPT\
%T�fu@�qn���DD%e	�W�#��*L"��T�rI
��0��A���"��-�Q!�)#A$�ub��&FHɜ�q(���fEԫ
���*-�b�ʣ�9U�
��.p�T���5��ȍC�Tk@�2e��L���G(�:E��L�Ȣ��,)R��TMB�,XEJ��9Q��č"�Ζc"�*HY\�L(*��T\.G)Aj�]:�E�*���D�՜�,A�I��+��:��Y��p�N���5}��];8�n���@U�i�G��=��A2�2�k��������w6�����ʴ�:����}Z��7K�������k���)Q�	�Lpһ��a�8Z;ϫ��3�d�<ȹ� �O��r��f�b�5�NC�@[Lvو\u��L���)�|55��i�ŀ�g'IQu�uZj:.�/,���y\v�r�X����W�k�A�P~��T��ToD�	-��\�;��yN��a���o�E����V%�A�Քa�G���ǣ]��}��ǻ���LS�^Im{��j��и��4�n��^2�1����T���$h�����\F��'��ս��m��Y=�q.o��wgJy9�']By$������sb��}��6Ŷ�G]���:�2�ud��^�=�W�sH]���,���q�or)���z�oC�=Z��f/xN��yq����Z��y�{��X�Gzw!=s�o���H�{��F�rڋ��o�M�!�{���*ew��#R�U;Ѧĺ[*X��q�%�O6-�f�w�GC4tt�A�)3+�*u�.gsx����=	KZ���t ە��� ���K�Ij�ٯ5�|�u�f:M�̼h[<��zA����(�����������Gӂ\:T�d�s��9���L��u��\*/9��Τ��)���J.�7����MB���jS�A-�6,�K�}k�\b��_ .�X���.iL�iw+Rc�<��4ܲ�BS!)]2��f/�ly�1=��������U��t���־WQx���oW�9�>�#صS��v{�Ǯ=���5���DrʎMm�穱|�D9����1JY�{Rw#uI��6���ut�r����E�1/�kݸ��+9p����U�N��}8���w2��!�r�/6�:ޝŎu<��A�#�i��p�޹���z���}p���:#Z6{h��W��cr�E�^��K�9��u]wҫ�{#a�lm5.�x2�g<��W�����5ˣ�5��K������?{غZ��t�5�x2�r���9�;�kDb'n��w��s�Z�:�,�u�R�҇���zzw�C��pB�d��t�Q��C��[8�Q�w�}�o_:�[�/���Q�L�Rֶ�4;˝���J���<�Һ�|�������uY컼��*S�n7�z�r�n�1;u �YB�����>	�:��B��/�Tm�b�<	S;z�p�t��N��:x��h;�kyپ�<���	ʈS~]K��/���ty�w�S�Jg�ܮd�Gd����7ݴ!��ޘ��Qg�˻�_g7�����Sl��C����2-�|�s�k�I��B`�~ΡX��TD�4�y�}!%L�N��k�j��>%���9���G�|�uK�}u������j�!X���k��cN�WH[����I���v/��n�:X"J����*۔s#�VR������U���s��4�M$ҿ��oFO��+�q�b�T|2�d��]k�殶sQ�������.wq�����;�p��}�����<7�˅�/se'��x���jxlJב��8')�&z_C9í�"k���(�e�]�ib	n�z:0�i�+rk�Ov�,�����M���J
������K��}���{D��%,;��DD��(��ta�JNG�蚔��L�.�n0t����}s�*P�Umk�հ1t���ڬ�5�w-s7O������>L�\�T�h&H�EU�*����U��M}���k��QɊ���A�Ɗ���=�x:i�Ŏh���7�C�kh��=W��q�F�U|��֦q��`�L,��j>��Q�ж*�v-�)E�
�G�;K������e�j'r�X.���u��Wg4!��]ٺ�=u������q^����Q]��Bs�������������vv6�,�����K615@N��*ȷ���r�c��֡*���ݎ�j5��&{��A-e�����j8�~>{���oϱ�w6;Zn�2��n��F��n=O��mC�K0-Cs��7Ԫ�:��r��(�v
��A���qܖ�����y�Z͇�;�2I\6�TV�D�T�f�8d�뭚��q�eY��1<��7�.7=�Η�Wƃ��]������
�My��Z��<�p�D�>���Q�v5�>w#=�=�Ƿ�Ŝϐ�'(+p$[K���K� %]Z�U�� k;�ݨ
Yz���
j���/������)B���l� � �qz���Žy���o����K�:�J��dŦ�����X�ݬ����J�3X�u�7�`��hI^����# �`���4�����c;�+d:�q�g})�j�t�'�4��X��54l�^��D��1�7����C��)uL���zG�}CQ[��YJow����u#M�*�vI��٘��]�ɵ��7�ٓ�gi�#f���\�弚��isb�%�wG�K4CN��򅻆* Ҋ���}E-���yկ��SO*�v�s,�v����nq�����:/36��#�u�#1w�t:�T9';����9b a�;Z��U���V��,��{���֔��[3��Е_s�Ԛ��r�m�x�����3��.����ߨOg�O�X�&������\���َ��+�C�d{�UM�w��h�7�趂�Q�g�p��0ԫ���0�}�񛐟gj���OT���׼�o��߇�и���캦4\ԫ�T`�Q5FP0�j	�������u��uܕ�쀠s�X�a�ޫO+�53hm���z	��r���U8@���̩ay�mYvu�N�0֙�!��k�U�y�)|�ƴݪ�s�b�����|�UPԾ��D;hi��oo^�&��I�i�K�g#&�����#��H���w�5�5(�1λjŮ��-����5{Q�ՠYV�j�w`�V��N��}��U�Lbu�����Y����Qv7E�3
�s�L�TiNi��ow��\m�&H���L����ݕ=�s�=&�7�����.N��%q<�ej����c��e�S���w�;�͜d��-�u'�[(& dc=��1W�TE������Տ����O��{����:G��%ˋxCZ9*���c:MԖ����/�7���;�;y�:-��)1��FM:F�m�B��	w�f�b����zD9&�z��K�����ޤ�G\&5TE�JQ�]�t(<ek���]j�զ�'�f/�F�d缛�Z�Mp��:��:�M��+�b�������G���k�7ST�{�;��P�4��:\�]��U�գq�/�g;�3LH�Y�")7Pm���͗�1Ԭ�#�j��������r�֩��-MtFKN���!u���\j��$�{wZ�#�ٜ���{2��-�B��P���s$x�*ԟC+w�
J�0��q�g��O'������fF����W��G#X��f:��(E�\���o=��V���ٮs��v@�F:,�d�&\�&{*���Ԡj���Y�z�]�~__X+�||FK�{r��k4�=��V^�s�����yN��o�J����ׯ��xu>�������'*�m��䕦�B���Ro���/��>�_q�2wl(���dh�Upu�z_%���Qnr��:�Q1|���Zy��8��p9YQ!p9ԥ;�9S�=�Y��5�$#�^�Ի^v��u�p�{�)�j�i9�#ۚ��{��^IM0rb��*��\7�S��;���gpQ�7��]C��j{oo�<�9+m�]��;��w\d��LAPgX�vu��NZ�Bp�g1wr�WieVFgm��m�SsU3�	���Ԙ���|�/���/w����z�i�C��x;r�[E�w�L���5N|8�:��=��Y��[٫&��%#,i�u(��]e�D�kab�7�wV��@m�ՈC`iPecj�a��6��N^���]��>�@�Ai�GM����a�sّQۓ��Ӳ��vPz�/;�%P�ۚ��ȭX�T�D}�k�][������5�[<�I��F=�r�|Ͳ�4n���t�q��I�
p����qwn�P������׮6�J���fg���K+��tpfi��W����Z�́�Pc��]+]`]�p;����9�fݛfQ�]x�}�,�o�L�.����NJ�Eow���������]�]�Z�k8.����o_*v�)�њ�)��Z��N�")1�e�Lw}O7ڂ�n����7Ť��2�>s����y�ޕ��q -�;,��:��VH�Z�)Ok�$��YԼ�3��n��N�������y�w77�N%���Ԏu%�:V&u�}y�}y�3��~���K�D8��j�dd]T���m]��kfB�\��G�mQX������0�oq��l��zĸ`�1?'؎{T�$`�Ek}�f9i��{����d�]jh�t=��6�n�nj�}ehS��;2kv���{ d�|�U�P�t�7bT�"V�5YWh�e�YmZ��ۄ�De�&'������l��R�}�K �h��������wRn1�pk]��[:N����`��/ꪫ�ؙ�w���1�P���2��[��|�m�Oe�'�Mԕ�ĵ�-��ZÛ�{Bn�擶�_Rͯ�ŷ��Qq�ȉP�"�NoqԼ���'�㚲l5k�G��q�y�<�5��T'���8l7���{�ia�N�MouG�Ԫ5����#^�����1�9�*M����R?���ќ�:dloTK2�
�k.1GM'�ͥoB�4�Z��faXp�v�/�께�x+�u&}V�M�=�=ǧ�]S5.&�RՈ>S'����od[B��8�f�([��F�jQu���n�.�@o6�B�g1n�s�8[�ҝ�p�h�OS�1�RB'�]�a�Ю����4O$�MS[ܔ�;��@w1ɪ����=L�C�]�z��vGs���b��$k}6��SX��m��9e}ʅ�BN�5�5�W�v�9F�_����4�慭�w1z��6S3һ��ݯ�@0���4d�m:�=֫ܔ��ݪ.�bb��4
���~�m�v&�eئ(�B�zy#��׶yN���ˡ���K��`����ڨ�iWۆޥ�*��DE�qe��v"����5����E+�ٴ�QBX�3�MvP�O,O�_1�������^c�zg-���M)-
Ԛq�n[��	�/
�ׯzo����`����<��d^=ՠ�=�o��Y���ёq�5�g�y�[}^N�?�7��p�B��ܾqGS���������]��W;���fn$ݾ�|�K����ʂ�Q�u��q}�y�Ooc��=8�ꊏm.���\.�o�O6��[�Z���j��5�UM�gL��\��k�8�B�N��\�X���ަ�^X���t2�Vs�ǭ�}��c}KS�y�|����oo��m��o�O>�r�cNk1�|zsj�1�h<����kf�w)����վ�h�0�=��nz��{G�q�|������]0����K��|K�f�!N	��y%�ܒ��|��]�r~N۾8�D�x:_Ux��{��uw=�Jp�]���>�B�,ޭ�j�.��Z&��];�R�n�]��]l��>�{	P
y6��vp޴&P�� [���3�7��t ��U��XXڹ(�)�z��c�N����|	�]'qQ����Aٶ�9٫+F��mo����j7��BUe�ub�Q��Q����`��ƍɍ��ʱ�p�[���0��-x4��Ɔ.%w�WU��֙hz*<�hZL��n�bF6iDk���q����/�K��o)���o0��[(@m�u���Ե�;e[�\62��=�"��}ra��t��2�NO%U��ೝ�w"�'�h�{p����U�G]�˹���*ʳm���7�<�_Ju{&�
g�!�ܻ��X#:�	R��ɆKkM���[T����]�y�&�Ap����B�sp&~�WA�Xx�t��E1�d�4�e��,�i;)�����9>9�Ʊ�!`
XƶV8atO
�L�iM�-Ga��t������肫+�ԫt��}T��H"å(v�V�EW-cc8�3���0Tv�9�_)w��$;O��Yc�hǗ�rV��C��W��w�P��gHY�p�b��oC}��Hwۮ��kw�=�=܋��~����7��Dݗ�OS)��u	���Cr�K�Sr�O�@��v��l�x�XZ�Ak��ѫ�����Y�ua�@ G*�/�%ˏTȴR�v����7O 77*'�b]�n
�
E�/�Zxfq'ׂ�"Vb}Y�Vb�v���JqQ����*��� K8��}�ysn��=V�X���H���9Z-�[���hשv:L��qJ����X���Gk�y�A��,Vv6n���J���\�����+Y}Ŷ���|�2*]
�朳��W^K�M��̔�Q�-���G�u�����%��U'7�C�A����|�]��b��t�ka\��§2`r�U���(ˬ�$ë��Hv��];ċu��	>cw4J���C�tb�Z���ެʉ3���8�����Y�v�(VT��ՆS9�y���HՖ.���o��F#0���X��5��kw;��c�������}d�d�Y(
�F�X��<7-�ɜ�\����g�\�J�vN[$u��&�,ڊx�Hެ�7���l�����������Z���_g_�zhEwyI�2vk��j��:�Uˮ�M$�F^�v�3�p�{�
�-���ř)퉨I����n9;7��Q��)Wm٫�ͧ��U˨�f�qn{�8TwF�m��{gXQ��JQu0c��V�Q��n�,��bɔq%v��VE�6����%Ȯ������$�o�T���pl��2�N��m�Uh�hȟSKV.���o��$K�ᖔ�҅���[�*�ڜo�#/�W\ͺ�|3�Ρr�a����J���f]f��r�H��1�xH�mD�\i3��J��k���V-���ɉX�w�$BS,�̎%ek߶^템r���{�$w��P�ѵ���c�_h�s$�m�>Q
Ր<�'*�2"j�rւ�aj&uXP�5e]��DPN�Ad$J��t�Q�v�ѥ�b�(
r�ֲ$YgeP�N뜨�")1�dҠ��ERg�É$Y�)T�J�͕]2��fHUU\�A�X�˔I�I"�͕�Uz��2�
r2Т���j�&�J�,�"�I˔��j!!�6h���juYj�2�������**�&Pj�p����0օI�EuB�9�\(�eX����EVM%J���3"�G
��r�PT�EU^�֕UE)* ��"�թ��TE�l�9�)��3�S#��A:�4�W(�*��.܅���Ъ��t�����%�B�(hTAi��p��'9FK.��\����(�<�*2ID��Ց&A2�M���TO6��E�Ni\R�a��'I�RE�.w9�XS7�j�гs���I�2�Y2��qX���/c�ۻJ��>���v�um�,w.q_�T��C�z�u|�֮!�ɧJ��W�h��^�Xɬ*x�\��Z�	���N�G��TBy���ƪ�݉�R���YI�l�������K�B�pal�H��,m�@�uɭ�t������gN�2۞���u�8TA�����bV��'�c�{���'M����c-D�xμ��v���X�E���\��j���*f����m9�J�c�u��r�eW]��,^!���s%�\���݆��ٻ/7��`N5�{,]9�I5�h�N8��Y��\Gb�wn�Hu�45;����%��~6��j]l
�(M�y�;���i��ܧ}9_g!��;��nqp�������$�ޗmP�[A��e�t��{��g*�7mNTc�u��(���C���͈ל@�n4�[�Y7���f��:����f�������]���s�ѫ��ex�����n��j��׌U�ݗ����Xn탻N��4z3�K�{���Y'p���Cۤn�z��F޻[~���J���݆a�Q��ӜL�̪�#M�{X��U�`.���{`�f)o5n�j�o��sEUsU���.�ѡ��\������GsI��_h�K|�=u����R��j�9�
[������5��>���cz;� ���J�8���9���Pe����WT�v�K�)��7ƵB�Pz`�k�PI���H��R̍x͸��,=��<l?�?�{��N����k�È����N%�rR����I�����/�f�餚V�wS�s�t��}�s2�ڠc�t�yj�vyb5F���?}ws�ĸ�z��o�<��69yza׺2ݭ�s��]}x��xG9�Z�]�&�4��ӕ&��:͞��6�?��q	�'�e�OnQ�sL�����j�L�zz�g�wl�����;�㭩/Z'Y>ЅO�O
{,d꼱�8�ս.Ufk����u�eG*P�����|��a�\���2w��Tب哇��ᳳmv�A�CPɚ*�o�X�f<=`���Cz�28�f6,82��L��p�C�����P��t�K����M2v^^ۅ�r5yE.�U����r�ì�ʹS+��=$�b�(H'e�땖��սJ�M�g�q�8��X�'Qʝw:	7y�t���fk��Ew_e�6�!c-��8�}y��Z�L��u�̭�7"�jf��N4�[5U}���ȿ�`��l=�J��꼜�/���QZmq��b����]o�r�*=��`�z���#�m�*>{�R�������oW�Ƕt���J;���S��5o~�V�����M�<ɖ���gt����O�S'�{ו��淓ڮ�.k��&������Eu{^z�Ul�k[��-V1��'�l�Q��iv8�o�
���=�φi�7��*�n�;3n�EK5zk蝃�뉭}����������y����n���D�^Y���8<̧1�_t9��eF�\*���Q�I���Ӵ��6�We�5t�g�z�Jt��֙0�(���#62?�`|n�*R�l�FɚU��tY��낤��&�H���'J�t��ئ'Հf?,!��J@;j�ɝ/f�4���e��	WVܚꯂz�gL�N�pޑ�n�f��>`��Y��7L�$z��;WY{�����:�s5,���g�B$���j��K���%�rj��g>5;���M���:E����ф��a>�9ڞ�8Y	3N�Kr�Z�i������:���ww����Fog
�=F���ܴ;w��ɇ���)~�ҩĻ���{���S�s�jr<�E���5�l�A5��o�m�pkr��һ&�ݸ�o�T2��Pˇ�n]�`��p�S�ֺ�����-_�E�|��SO��\�5����̎�Y�j��x澑�b�3��o��U�w�kj��m��-�V�9i����7�bsx�\u*��M�_Rا����K�o�Aq�>]�V,Ke>�ڍgxv�VQ}�nӿ��\9��;�M���7(��8���Q&�oWF�B�uk]9X�;qFnw&��Л�r=����V�P1��8z|��OA�8꜁s�U^�!M�u.�}�eOz�-��*�S���<-p��j�	�����RkBt4T(L�e�g�U�ݑQ.|c�<�qь5tqG�N�D�R��AU���+���57�t���f���SK&k��W�%�ρU��ܧz���ۑ�yB���y6�4��u�gS�,[�y�]o*m�:ܮ���#}�6���Q���2���ܹz&�Q�\�6��f��J�c_��Wp�냳�k�D�3�TY����Z��t�+��gq�x���.%���9�3�Pq�j��[p����u*JLW��`�}P��ݍU�-��wh[�����Å�_<q�������ts�_Q�FK��!�ů*��A�g<�Q��M$Ҹ|;��?S���eX���[���VR�=ծylV��&:���i[H�s�K#�󂸇E:���f����m�u�9�#��:0��	Z� .̸���im�穟.w�q?A�����'��w�o�l��e�х�L��9���@W0�+�R��j��s5�n+�gik�vz�s���JcE|Z�+r�t�<3�Ή�L��B����W���{=��u���P��˨
���v�%o}y�`ɕN'<�N�5�,e�[1���d�_K��e�V^�qEK�w`L��G+�%k����nL
���`����Z�+Ǚ�!j�V�">��u��v
���r�O�<Y|��1�M��Z�R� ��GsN7��ZPd���� �׷�����%/���rI�m�~nGV7ik�y����ծ]�����ް��v'��w��r�Ou�q�qp�ю��x2(����9w�EY]�gL�m�ǃe�W��E��
��1��p�k+���6��;br��W�E�`ʈKf�qË��:]K��b�/��y�S^���~�IE4�<;Ц��׫���n+�'����}S���[L��m+�����k-<��qܖ�-e�Ǜ0�Z���Q���拉Ʒ�gi���"uGn79ڥ��Ul�W����mvSz�u�� ���֧�C�[8�c�5bY�K����o�����:��C����e��wjLg+n�������V�.i�U�t�Ҙي��OÞ�\�_ؐU���J����N����~�o}��8�eL�徥�*�H�J��G>�\��l��J_p��r�ɷb�w��⎲mr׌���Q�	/�|3NT�z��E#��:��$\M�־~�[��-ү��עG���թj��=5�v,���mA����/����G;lv-a�y�}܈���>�]iA�����mTw��ԭ��㻕b?v��t�U���;��5u��iM]z��u"�etkD%�[����8����Y�����u]����%��<�O0�ԥWh��Jܱ�r�Mb�׭)��'�3�eWȵ�����W���ωG�3���:�GB~1����_�:�b�ޗ�"�T�=�O��kF�s�vLg����=��~s�^�:��:�k��Ն�����F�7=��V��8�Vǭ:�|-z����@��/mX��F�4|b_	�MkCT��> ��Y#��v�z�L;�6���}\_�L)_��>��Ϝ����B�^l\�{�����ɸ�`�T$8�a�����#U�k�5K�k�{�c���޻�_��Vq�L����b�U?�6��9f��z���=E����o%t����ӥs�����ARS������
��R�;�׉a�+q�dy�u�����H�7��C�^����9^��˛�kt��x��Ny̧1�!9Sޫ�s����Ң��~�q���Q�8JGͫw}�>���U�Q�zH�A���WE�R�}�5��?���/�y^mHG���wo���3W�	�O���e�¶�rRM✲�}�7��k��Q�u�[��ơä������[K�u��lV�ssuv�)���V]���]8aJ�Z�vLNr^�T��υ�L���mJ�݇�7��<6<�^����G�ز�����h���uz�
�W�^�F��*n*��T� TY�U⻄�g��8��w�7�)u �Yq^Ձ����c�Z3��w/���w� h�P�LSt��+���F�����J(o �7��]�k��S��Ϛb�kc�hp��z�-NQe��'�nn+�@7(-`X##=Ώ��.q��}���(��Q>�Ӵ�?IE3��:+����/ޯ��@of�&�-U�e�@�\�̬ڙ�y�j�YP0,7�j���b��u����(�~�Gѵ85̹  ��g���3�k�X��l���c��}�3�x�9�Ki���U+��zv��s�;[��LS���z��..D����Oi�d�'�IL���.��MVѿ�χv|1���:1�k�������ve͛�WNz{;���/�YT>B�72�ۈ��}y[�竤�z}]�Å�f�exa}p7Y��{׻Nr�Y���;v<2�DW�bJ8K�f��ݨw��7_ 7.����;RWzF�Q����1�֬����b�P jո��<�t�*r�2�ՍL�fWU����L�e�Z7{��K��O��Nk9ڻ�3D�a'!2�3�h��@Ò}��	�8kq����ڕ����07��(p3��Du�w�.-�R�0ɋ�;��?Nh�U����k��V��򻇐��m	(�̰��,^�Cq9�#�5�;<��Ͼe��=�ыG��zkYD�/HG}}Q;���h��迢}(o��es&�ϏWGf�(�����k���8w}#}7�,��<�7�����\��گ>"
"
+���]�s���4z���;�VESQ�ZX��g|oy��z�u����E��ב�s�o5{��]�J�V�5*t��fx����G�;�G������|׆}ig���zV'��]w;|O����蘶du���3gՅz-�
�U��8l{z�Y�%MIa)����z��L�ڨ^(�g�w���T��]��f�E�W�i�e���Lh蕊�3�;E��r�x��`w�����$,�4�|r��oU򖴿}ά���@^��G�K+�G�_�g��>S�Yp l���q���T�wmV��懠��'
��W׭b����0;:�#�z�����r|.���O����g�]\eqW��a��Ԩ�į�2�mk�q�lMǪ�1��9�#���.3CKZu��~񬠭tp��c3�� �����	�������mߚ�%-3��.���nBL�U,�D� {���2\S5ݡ���L���*,K�\jI���vd�n"�s]/�F���e�-Gi�J�����.�����H��jz�["\KuM{�#������c� �t������� �{��,z��"�z��$�Li�c��k����MWo�'}��ٰ�+�'�u�|	-��@|o��E>��z_�v@UL�ǜ�]߲���VMC�gz����ր�i�*ߨ�ng�m���\f�
�;$���)�Қ��ZNyy��~���ྯ޳Q��[f���	G��_�Vq���e�F���pD:�/s+6$�]��?}�^[,i���O��!=̏b�Qs���6��q�y&�������%�������r�c�(�߲wJâp��|�n[�b�lxk�o����������7;�\W!^fHÞ��O��'�LU�w	��ӵ.#+�X�͚�q�@�\v�������D���qٗ��gs�j�W>��!���^Y���]���{ U����ݯ!�^Ӽ�u�d}��F�����{�]U�v]����yӜ{��4_�Ep�̒���,a�(z��;ɝ��P��P~C=3�}�#o_����UQ���~�����\o��]���[�8���膮|( ��e��y��͹hf%�9�� B�I�ƽ#F��J�ߝK�3�v�d�~e����Cb������k/����퇻}ei[��T�=Ff��%��DkA͢>
ٰ&�a�-t�6��q��-P�hS)ʢYϠ�+-RM�cC�����]#ʗ�7��xvT�Vf�C(�31 o� f�?Q.�uӞa�X%�WS���-���v�C���J�O+�2��㑩�yq�EՆ�l.��\���3F�,�ht�8�r�U�*���l`Y�Ւfɼnؓ=�a�ۙQp�+��`�L�q�{;3�>�sK�cil]i{.�R�0&��;T�gi62����^u���-�!��V�-K�'+#�ѫh�ǹ�Ѷ
��d�Mn!��F�n�aw]|�Ĵ�_`�y<�c��h3�0v�G�N���W���i��m*ɖ�O��}6k曛B���'+/&��ù3�`�*����Q�t&�u�տ�k���&���i˒��v܄,�vF�B��1鮊��3w�t8�\���s	��V�{�o��Բ�
�L�j[��`��7�x�	�0���յb��:��.���vv�%�#M��"���H��rf���w��X �-O���C��Oh�ˏm_PR� �n,�e=���d��	v�>�e)x�X8�i�Z��v��/z��{��1P�VGm�N�S� K�L���yc'!dS:�㇬�&ɾ�y��3PoV�S{Pz�5y���❵�g7����zYI�R�D�Վ���x�=鯬��� �;}+j��GWO�\��D�Qe]�kh��5Ɏ���(* ��_��=����`S�zpٶa��*`ٺ.uk���kC�s۩a��̎�TH�*��m����'��*�Ҷe���p����IS �e��A��6�� s^�х=F]�x� �E�2��@M}�^�t��u�+轶H��˲��6{�m��PgAò&�� �h�l���A^J��lh�)���:Lh��&��];i����]�7Ȟ����n�f-��Xң�˺�y�m��y5q�]oA�6����K�A�LSu@{�w�`¸��/7Ʃ7t�7a�ݜm	Ne���J�����tQ�@��d@�NUܬͤ�q�r��(B�O���*����Qi���	�f)Y�GT����EƑ�ݦ�uw@�y�2�N���k��v���T޸��:T\;�K(Q��\�q�՛׏��3B�72D�`;U%�]��|2�B��{;{�c�6�b�ֺ�� 4@_�/rju��3��4��(Y�aw\� �� ��q��p����ov��m�:�Ep�f��1���:j�0��QI`��-��J��L<���y�t��NH=j��/+mmA����}(���@h�z�^Ʋ���hyJvD(��Xț���N*���s\���t����?Bբ�s���Ȯ�;��+%9�EJT\)�IĊ�*�3�	�3ZȽγ<��C�Q�5�*��E��`PA	Ċ��sS�2�̣�W/8�Q.��NA��TTE�.�F-<�I�(�A.U�\��,5@�W9DNeYF�TG(��=1	�J�"�����d��E�<�����U����%���!ܖU9�w� ��"	RʥH�L�(��rL���LN�
9«�Pŗ�aU��\�(�+�̎VX�PADB*��\����� ����1�M�r(L�=J%xNr��ˑ�%H��
2��[�
D$)*KP���;ù��IʔxN�!Ri!/ZW
=B��f�4�#�
���ҳ!2��2
\�jdk�]�tӇV�2(�r/�<=�����eɕ�\�"�E˔s�Bt�wwD �� ��K{x̣/��}Y��g��K���u�X�����@�9��ݗs6���&U��v�>Q{��N��?�Ġ��b���_��[�U%�惿�����z_�Gm���z�;!�,�jŘ�r]m��������6�uzM���f��tG��h{"�3�#�.9����w�n�>t�/ն�k]����@��[���J�_�9]T�%#��/��k�	�Xq��=4�5�QO�=���ލ��Y}��>s��<[4O@n�*����RÄ�}����i�^^�UZNd����k���gں�/#�dp�S��W���G��̀ٯ�M
/��r ���w&c�n9ej���[ެ�M�C��N��rxp�~ ;�ّ 矏#>Kð��"ӻ��t˦}z�MVu��W$��������n����ߎG�u�Is���s��L��<}�8�/���dOMn�Q����]D;+L��O����6ӱq��u�s��ǜ�I��Q$����ɫ�|��7��2�V=��Il���G��m������ky�WLz�:�|/�\\?:�B�g��GUΜ�Q��ۼѱ㑈jlg��A@J�r}�n'j���6}���<��%���"��f����S�yѺiG�]o��U�K�<����:S�mvu��y[������d�����֞��Ղ�v�%׹��V���f�L^m�Ӝ�2���F �Z�'JԺ��z �yذ��S}��}c�I����,ܛu�bÊ�+鍳v�-W����a��~�۹�?4�-W���q�$�˙h�هg~�uC͙Á�셗>���@�����5�C{�� {���.�(�םr�8<�N�'���c/+n<x�V��)�Ys�绲}|��\�^�y��{���F�{U���D��ÿb�bk���^�q55��&���o�o��y3���R���X܎s��;�~=���j�\<�.���{�(��&b�zW�k��#�',�6
�W?\����οNmJ���g�:1���{~�W��u�9b��'�֦�uj��;9��͡�; �>��*fX�O"^O"�j�?�g��ES�E�B���y�ӠǻKjP�D�C���w!�u5�<z�����q�x��P9,�=��J8g�=�y��+ѾԼr#�%������O����S�Yxnj	����Я��H�l�ϳ�}�Z��W�_����Md��*6���6��<y���诽��юe��� 4���,9�����A�z������\����9�ә������&��ּs�;ģ��x���ȷ2�Q�ll�yn}9Q�X��X�����s��aIY���ɍ���В٨O�v"9��]Љ�� ��QI՚�|zӕj�`l�k�����KIҫ.�k���|�ނc�f��Ex>YN�u��XR����x�q1���8L�:��N<�����W��|�7�К+L�f�J��������w�ba�}tɯ���Ҵ�@R��'��[>�s1~r�3G�u�1�1G����g�o��5\�c���cմ��o�<���G��LLSU�o\�wdLm�ud�o�~>�s�j.�������(��U���S�z�� ��?
@�ϑۉ���[��z�MF���|�Ç����n�V7U벞]�1��vQ�� M����E�o$��9��7߁��׍'���t"�7�i�x���g���G;�f�^ܿ^�,��T5�wI��	(��2��s��X������~Y�tuO{g����V�ٔ=�9Ł1j�����k|Q;J|�����*8|�%�����mx�-�~�LOc��~w߫;xe�֞���7�o��e�ڝ��z��sO}��q9=� ���#�[2�ۍS���p��	ZHvs�X�FMib�g|o\���_�o�}�E}~�?�D�WlY�ח�#ޑ������W#�R7'�O\ET?�1]1q3��1˶iY��{�a�����=�Y޻��G��6{b�^
�塣��(vzT����w��L�vO�s�}/mƜ�o�1�vɛ1��Ғ��$�s|5`q"N��W�zQ��
��8�ǍpԀ�����3��rͪ�wn5,������)M�e�	�T���b5���]�kkY���}�����[2��,Iǀmh��.��:����g5ʎ��3�4?Wo�\8I״�H�q~�<.^+b�Uz܁*�΁ޛ�,�UPH]��<�/f�"�h6k�V�|����U��~U�l�{������|n'���G$�� 6C�h[��ӻ�{��π��V�
��x��c��F�U�|&���c#�e��؎=��N���|%y}ޤ��;�&ǌ#F/T5t+�W�Ç]/ߺ|�Rު��Qs��^z�5>��̫K�U������EE�F�|<��}10�_]"bb�W�����,y|�M����0wk��b�>]]�No��F�����nT`�>5���h�̀����14����~=��~��4��[ca.�qX}��p���^7���ϔրǽ�ȫ~�����[fl1ٲB[��Ա�=�����7���Ì���)�N�F_?Y���qP�=pQ&�<��N�����Ǚ��ۉ����p���ա^N�5/I�_j�=p���{_���5��z��=���Z�zz��\���v^\���S���I����ׇ�3kG�'Ei�s���-����þ^�x��^���Z�U��Y~Q�_���Ra,��h��]�KUo;{��3.�ؠ�W��pl����Ԯ�ZKw��k`^G
Jf�ɒ�������}73~�#\s���D��o����U��G�I��>��)�9cB�1��An5�9W4���*̚�c��U}ːPwS�%�Nwi���;|��5�1q���<�oӵ-o�=e<�?e��j3뽥п~�`�RA�f����>h�w�ï�!��ݢ�_���9}�VET<5���=]f���r��.^���KD��:g#�td�~�=8�v�|�R;˅!y�Q��e�=7P�*�~���5��r6���S���U��|�JҠ}�o�~㑾T�|����#�c��x��z�����:�L�a�l����po���zXͩ^7���ȁ���#ޟx�k��K���Ϭ����h�a"��ws�K�l����g���rl�hک#����U�tg�J����ק_�W�N����mL�EW��L;��5��9L�pJG�����5�
߫����:�=1�n.���ko��(��/���^�dxb��ynk�zwJ�W�z��%���w_���O�&�ڿb�M����#v�r>>�@��P�~��9f���s 6j-M
/��K~y�®������Rq��_�mw�~���&��u��/�����r-̹R{��L۪���<.�ި��0Lmvq;H�rn�lV���#���=��Ak5Ȍ&�a��l�U)�2�����@�de*s�>j3w�W��Yg��Z]N��!�Ln]��V[y��)�����t��J��jhx�f�}�7o`Xx����]=���\��Ec�wi��1�S���ϧ���L����'�Q���W~9���}'Ӓ�E9�<o2��ʁuS�����]���>/�M��TC���E}�wǡ���Q�ύLw�·����ϵ��w\�z�L�Ӓ��:��>�ԲV���z�n����������5���f�V��4O�|�A\Wv^��#.���䧗�S������ǫ��7_;0��[��׸��=�n[ >�tcyy5u�U[w���3�Ot�w�����H���V� O%��;P��g���f�iE���c�!�������;�#s�v���`1\t��ww�#a�����<{&|3M�챎1�s�^��=ٛ�Uz��zΏ�{��_ڽ~'<mއ�F��\Mǻl�oh���6{^K��y��P�3�
�R
�kO�#&uLk!9_Oz�ns��[�����6,T9�ۙ����Ъ�(��8JF����W���{ŋɝ~���A�S� l��FC������d!8�>�M_�{b��S��};�q���Y��(ԟ"��SȁVy)�WP�zk��/P�ʱ���_Bz�E���&�Ԙ��l�m�cī��}QV�owP�:8��K�k����%9�T�Fͺ�WMmh���)�j�7�:��l]��1D�Vo�Q�#њ�kB�s��}l>�egn�ޣ�r��nWK��Н�[�z���}�N`ّ�`���i^�f���l�RtF�RZ��!�u5�뚇b)�D�^/)z���L`=N=3��=������y?\{ zR>�|7zY*=���^*�˸75�:su��	�(��-�Yյ��3��[>܍wiTO|�֑�~��g=�tTE��ȿ��Ix���F��:~�z���zy�z�z�
��x�@,-9�����{��|�ɿ�_��8_{r�_En�X^����j�C�������_��E�"���a�Ki�����J�1����X�}�=��:g�1~I�߿H�f���$y麇ו�bb���q�}ǳ्���$� �%�s��V�~�����`Ϟ�)T'f�@z=TA~����;M�zZخ5K��Ly��\�~����i�w��<�CVi钏C�<�!�ݏ �I�$��,v��l/�ڇ�k�y�L{u��u]>�iz����d���6i������ψȄ�7��e�U������r�XZy=`�j��������q���h~������ٿ�K��=��س����<JG���:�n=�G�~�}���j�Hݭ�zY�`ӹ�� �b��|�N��\�s�@���=��R@\Ì���^eI3�	�j�l32+����{�,�������;vAs8�H�Im��3l9�m�*�m��Z�עk�\U�%e<l%��\�2�]��%��R�V�}Ρ��"�<�rgX�*Z~���+o4��!�? ��nv�2�&��>�c\���V��'��'8�n��^���K�EUM��Qǹ,��C����c#�'���)L�j2kK�;�z�|�t7�U{ĎǏ�l��n��'��N��4s֫G\/m����Q��R$05F�?���L�8Lr�U΍�*��,5��)��BR���������z����P� 쨒�SsP����\3��?�:$�1㸿$��x�����~�S뇐9״�es���p�x���S�Y�c�P�w?fJ�~�3eb�先.sր�{��9��-���o���<�-�����v;��7��W�7%��TɆ�������(��z��+>��ۥt>D�c���@*�j�M�~��g�T��3�|lI����_�oj*u���W�៩�S%��$������<͋���n1*a�2�V���Tְ}���6�o����s#�U?D9f�X�����_�"�O��p���L{����z��'��z��/�>�6=�ӫ��;H�ZQ�܉�Ɛ=-��@|j�&)������Y��w���K��o{t��p)���Iz���5��;;�2��]�c�V����S�l뎊�$��V�3"1�����=�s��#����J����Pk������Y�}S.'�!ұ?��+4�*N_�~���^`����G�׍�U�38 ]�l��~������
��d�)y3�;/���������rR��#J���r�q��Te�?Y�o΀�9:��\@yD��)�+o���	�ZWS�pO5���}�M�fև�Q����3Q�_����ǲ��˘�8�����ǋ�UR�O�Qe�v(�e>�����[;s��~����:'�k���}�l
\�*�}����@�8�Ņ����&��x�>�ܫ��8c~�{M�h���<��Fl֛�r��� ����gzd�(�m� ��=�G�״�9
�z;=����N�=�r$�����ڇ}���~:�d$#�	��+��wx�B��~Vɸ�8�v��p�����H\fIGIb�N�Exm��NB�� ��C�[��E��g����	��wq�ׯ�r7���~��'�����6@����.\ڙ�J�ҧ7�{F�Z�Q��&S���^7���z�{K�x�9~�q�X�6ǲ=P�9u5�n�͉[�~:_
'H����O�<�&�Pl�F;�=q޴=�O�ё�
��x\�����*/6sU�r����Ҿ����!S.�G��!����������o������2x9Jn��B��Ժ��yσ��7��ܙ�#���	���,�y�%�E�3bc���mU�wyZΫt�Ž�;I1��h��VLaWȭs�=����^+��YZ7ҏ���q�;G�9�rx�����0JG���^s���U���H7�Ԍz�Ӧ�Vj��biy�9;�}
@����:�ǲ����F+�K^+�oJ��Mw�:�mr��
��-Ӥ�|�ԁy{���w _��p��;q2f�M���uf��s��n�5��w-��8�;��L{ơ�+��SY�9��R�V�Ǖ?S�s�Ia�1�S�_����+U�g�G�?C�"~�+N�@>��9Kҟ��w���s�:Ϥ�:�\?m����C�-�޷[�������0��S÷���ZdW��|{ j�;9ظˈs����HS�e���5���-�b|�[6O��/�|U��5en��ä�Ѯt�VǓ�'���c�V�Y'����y��(/G���p��c��Ey+	�l�B��V�q��=���c��J\�z�%:x�Ncy^��3{^!��T|���:7��1�@�7�-�;0�߶a�����m*�o��y$�C-���@V�����םr/�oEh���<x��?}ٳ"w�v��ׁ��ї\����e'�����Hb8LVYw4K�9�	tN�I����ppo+���"�Vq�r�Bug>�ԭ�э��=�I(�ۘ�+&�!�M�F�]�P6�Ԟ��֘�����K�Lk8���e�e��jֹB�k��:;�ޅp�6���~�f�Y�^D�v�Fuhf��}*�eB��hK�@����%�ec#�M�<��n_�$Y�
���x-�8�瀷A�u,W���1���c�ʵ�op�s��9�5r,&�<o��9̃��ݚ$����v˳"�R��s��ӡ8=i��5�V�νt8IcYU�銥�z����&h5�=�1<���"N�=HQ�$���i&�n���5���|85Ȇ�b
�כƎ�P[��iH��TvT�����#t��^2{���g=��Ѿ[mr��'M�WF����M.��E����k���kH4�Uz5�{hDB[��
��e�4����Iq�rtN�ʛ��c�7����X��2Pݏ������g�-L���{������:�㐒ufAe;G{�X�Yt�[	�BU�%�b jm�rWkM���n�v�Z�7#�X铇'�; ��Y�1G�,������dJnqY!�;NU��DFѿ�d흊�.KB	��3�-O��W��Z��;�n��&�o̘кeJ4�l��q�]��s�S�6�V�n�9AK�y�L�WO�B
���a�ؘ�i��r>XvS/��b��>f\�˧�7��֌W���9����	��kz�7]p�Ñbl�����D�z�vW,�:���D�������kJ[X����{;�;���y�K&u���=�KqzRG�G�:�Ѭ�s��4�*X%� d�IL��m)&�ouҦ�j��kG�efI0����BYJ��˅�R�M��>�fsn��Fps �m��!��k7���P��:f�Ǝ�/>Vom�0���F�*7��M��y݆�T�5DT�^��4�9�i��·������u�g��]�2��s0���Z��B�͕;�#�]�}�>��*��F�6vf�]��>�����Rr�����e�d��jY��[��4�(�1S�9�<��~Uz8�^S%�wH�܁���7_���+5|`���0�k��K7��p��e�wz��ᤐ�cf	� ��s���=�D͋.�Fꍫ��J:��l,\4|�b�b�20v]X�3�w �;.��*�.[����S{ټ�fA��8m�]�b�T�Vq�mi��;r�-.�NϢ2�|qb蝥B��W�9S���siE�>yy��zXJ�K�v���ֺѾ-m��D�~�-�;]-�tA'{��n������������*�2�Yb��DR�S��e��G�T�
�" ����A"O<���9Dk��Qʓ� �ҩV��a��B(�:M᲏&��YI%UQG�*�Zx��AȾ(W9���¢̠����JN�D�DvMͪȈ��U�E"8y'��fEAÜ�͑QDs����Y�U��
<�5p��)�"�";;)6N�<�f�qx����.*W��;O��EP�\��dP]ၦӜ8Qs%AdEUS8AED�*��E9�żqu�QQ��	Ύ�Q�^Y���*��8��*xeTG<�g��Z䔭3�H���T|P�l��\�V�L):W�]K��e�S�DY$��ʸYEp��� �DEW
�H��c�kJ�v����M�m�sr���x�ˤ��z�{��t��F�|��\�Ed�@ܵ�f����Ԛ�v�fl$�IKb�-�ԗ~�C���*��K��7�}�z�J�[��R�~��o��G_�k��U�{.�� ��oya�C��ӳ�����t�rg}1���uz�ns���=^��;nw��P{7���{��z�<alu��;�^�_YG�����=U0'��b�g_�>�tC�2�x���}V�e��'׮{z�6���}iYF�~�q�R|cVD���T�ES�"E�Ed�s��V��"t�c[�o��L���z3\JG���Ļ�G��C��'���"��O�hH��_K͚ܼ�;����Н���c�ȷ�l�AC���#E}���G$���'�n_l-�;eY�R��Ywӻu+W/p��y>��滀�E��&�u�H���S9�������~�W����������xl���nx��R��U@3�oAai�R�o�TO��c���W��|Y��K��4��Po��	}��Fq��m"@���v�&�D�=�x��(c�?[�^�u����o�O�G]Y.�}�3���e����%�Ih��^&)��;�|;�K��!��d߯eG��F��|/FO!���U�j�ֱt�Ceg���VZ�v"6��{����kl��[���c���;09��nWp���cb]2����oMHJ�f�q�u[vs\b�v��5l3PcYʑ�9y��h��m.��#�D�"MO��mESfu�h7c��u-u����h{���}Nǜ�I�=P<��*<�)q3�t�����0�3��r�z��M�A��#ϻ܎ߣ�Hh���ׇ9�����<�ʡ��^�"��Qˉ�;n�^7��5j�����v��S�|W5�p�m�������L;��nd=�;��Q��#z������U��g�j'K�V�y;[:<=�=9.Dv�\{#�uNGzG��uĶ��q�>rVd1�y�L��Ԟ 9��~ζk��if�W>����M����O<zm���D�·��,��ً�5�\��J>�wU�ё��{ X? �V�o�5�Y�f?�r�~����ˏi[s��Ͻ��SʷJ�}���JG}s�S�_�yu�b��nK�z���b�b�gY������U��t��Z�nyK����;�O��~�r���9�D��6D��,r���`)�ņIUU���n���矰��h��mT&n:�\<����x�Ӯ7����^
r�/"�)
�2�U)�C�j��Nl��ew-���20Sw�o%x��u`�q	�\{ /Sg#�%��=���O���2�+�ފs㱕��8 �(��;�ll֝�}s٪��,绞��<4V�^�z�&��yS��1�Ճ�`FS>9Ԇ�z�Mԭ\�]ÏJ���MlJ0�ݚ����O#6�Z!y��[;�=Q��eV�����Y��͝�,^�7mJi���<��ܮ�����Y��= r���B�����X�;����Z�-�q��ȫ�əG�*O�=�^�K; 2���}q��I�P`�h���*5�+�a��x�F��w�lLx@�~*��f=�m��K5����=��9�9����t�����/T�c����9�w|}L�����k'yU�kz����y�\3��G���1�/�%�� >7�b�qK>�Y��O����K�G�<�v@u�q�֏yMx��K�<�ր���"���&���[������{r+:��>�����u�k�>��7�񿓱Q���p�C��	�p�c���$�Uzy���]ٮ�M,ˤ�=$���y�����Z=y;�5,i���,z�Os#��%�(�8���^-n�W�9����7�Vn!ʽ�l�ߤ����3�g��FN�������l��^�~J���cBݠw��ՙ�Z���O���j�7��Չ��u1_y;����w�e{��5��\��JF�;��W��W��c-+�p�kd�|���8�Z;������+E�碻�D�a�3��mC�x�t�K/*4��!|U1\v�,a�S{d���5ښ6���*M��&�c0A��y�;G�m��wۺ��SYy����Z�J�B�bz�ר���צ�=��b��lW��0��N���I��iv1�w�v��.��+��L��u����p�^c�n��T�����9�su����!�}�H_قP�X�Ҕ��}@��S�[SG��4sN��?]ü��M���^7N�7������k�\o��|<�J=���//ʽaƻ�V+�\���	�����>�w�e9��ڕ�q�������c��/�}������0�A~�S�Au��6kї�A����N��*�<�&�%��c�#ֽ�C����cZ��:3Gx̭;����1�+����K�q>�\{�,�c�tjH�"�D���o�x���`.�h���s��sf�w9�V�$z3�w��Ĵy�t��~�\xb��y�!��zwJ�Q^�����]��P<��i����G�F���i})�H��8U�����ơ�G��̀�^����ϭ���Ë���z ��Ñ�waL??7q7������V|߱ =��Z*-�9Rm�o����g�^�T��.��G�0xmZ�&�=�p�p�O�5�Q���3�>����W��H1�.�������׀�(�>3���u���!�\�2+\�g�KBv.2W���ZJ�	~�=�>�W�;&�F�t
3/;nST�%kZ��ƕ��n���;�]���i��`=�2���C5�Y�J�sFW6$`�
�WЅ��1p:�	:�a��]�:�����{\J���O�L��+T94�Ze�{�g�`��a
�����Wz�J�e���Q�V�y?���k(~��IyωZrO�뉺��+t��'ä�k�k�Vǽ�d�W��,����s�wjP���RG���o����A����I|t������{��[~�~+
u�D�]�w>�g�����߆B�QjNw���<�N�!'�\�Gn"v��.�u�<U�ǛGT�9��r�>�Ox��� Z�v����9�'P8��V���V��=�ǳO��rQ8�n�饵�=#Q��ᗕ�q>W7���o�s�q���o���=��q���ڮ&�������"&w]�>�s�dzǳv�|r''�CՓZ]�L�/��@�����ۈ���7�o���|����̔u�Q��n�MO�}<}��z��G*(ՔJF�Ӏ��0&"�X�����(5N�9�{Ũ�{���Kr��/}���j�=�~�#q/����Y�(��|���`LEO"E�Ed#�J��ﲞt-���F�U{<,d��������[#�V�F�T������q5vRW:�ކ���su�T��c�d��Ϸ#}p��ߺ���-��-��Q)��~�h��ܾ���$L���$O~�͉�CL��h�5m)ߺmu�f���6.�r�f����
�CC�G�r�^�7��J�a'ym�]���O��v�7�dy�jK>�wj���8�Z��Maާ9A3�i2��T_vH%�s^	�Y�vwS,Vkr��9p
V�9�(����c`.�2s����կ6��U�o%���P_[J�o��;�Ȧ?U��x�_�Z���yߓ�;��fs��}�Z{�N�9O�&������|Nf�~7�n�o�WZ��L���UoӞ�����2Y��d��<}�r��7�-�\LL/U�&��wԸ���'�A����L�����^�N;��c�WZs;�ߝ��s^����[<ja��x����h���ú��xl�
3D������W�M�1tԛ^u~9�C�rN������	>G6&�\en�O��TRRT��Z�.��z��ɱOI�p~�A�g����	�ꢍ���&�nǂ���d;%ؙc�)�*'���߸��E���˶�_ٴ��q|L�ۗ��/�zd�}���lo~D׫�&SG��w��qM^CPf�{�I҅�F:��2v�n4�����^����2���HdWQ��ҽ=ᚯ<y�Z�O��:n�Oi�r���1��ZU�d�V���#}7�,�O<�H��5���9q޾꼟U��P>���5S��Y�-T��{ X? �Un�֩�,\d��� c���ZG��M_�Ӓk���t�q����]�_�֐{^�X�!�ە�����y(D�߰��or���oW,C�<�{�[-�.l���qς:*���,�aи�iu��0_�.�r�Z�ЉB�SE��Z=^y}veA)�]jƤ���=�E��#��އ�hvyu�b�0JF�'�*���خ�U�T~�:n׽�4g�M��s1���Vcr!s��#}��=���W���4{�%�'��K	O�Q���{gP��K\hKn��y��U���\<��s}-���~�8\<T�������5�O��󽛜D�V����pٸ��LS��)����;��JF��'Ǹ�������{yr�X��]�5΍��_��qw ��F�9mz�W��D�Kgr5�
�ھߩ�ڤ�]�������lo�DᮥP�9^��-�r���V�񵮼���,�v����䫬G&��}>�#��\���t���\W�f�g�G�baz���>�i�wu�ܻ]7ۙ��_��@� �ަ���*��
P�|���D�s�H�h준��Q�?a\LbxZ���,�����=�T}���݁T=7���|2�_�z]:� {�l���,��^����F�]������}�a�m<��?���=��n9K�iب���6n��rUG���ǵgG�s�z�n(徐���i���u�|i�h���ڱ���u�!
[�Ӵ��*Gsq�]}ta���jtp ��d�H�!��fŹ�Kn����8�v�u=�u�.���k�aM�Ů�u��$�2��}|��XOM5YЗ)H����ۆX\n&�q���d��Kj{��O3#�����]ٝ ��W�Y=/<3]f�܏�<��*�*8kߤ����|Ν��;��:)����3Z>��>7���}�������U��{�U�;���eX���Θ�����rZ;q;P��ŋ͚ӭC+yg���M{�;�x�����t�`_����#=��7���,U�������C�=��YK���[���q3��z�ţH�^;��w��f�} k��wB6�q�[;��k�hpϣ˅!�J8���3=,7����N9��՞��O���1�ǯ&u��@L�GS��h���ǔ���S�|��y��U�e��~�m�>Hup���F������}�q�)φDmJ��sA��^Ӑ�>�h�S�:#�aoU\�f�w�r{�:�b>��q���Yef��D�ޙ`g�<�&�ͤ9S��޴=뮡%zgs~���n{���T���>�q�Q�G(�K�G�WU"`���^6��z��U�Kv��߀�>Vċ��������H���ó�U�P��CsD��*�Ϫ������*����8���S���d��t�V�紎*V����r�ʽER�*�NUst�W|����P�E�,�`s�.\��I��m��d��%����ʵ�19�]V����WaNr�cEg��[�">��m�_=X&q�ݍ����@>�F��]�����ґ_?u ^}�,��Ƕ�|3�O�C�G����S~�x�{[U7s������١E*x@b�:a���TO��WZ��N�����۷#]G���=��ģ�&���$�e���(:�TE3�sA~;�
���?��*��Ϥ��uy��S��36�_[˿ ������J7a���n�����.V��wǲ�6ӱq���}z-?\�ZȯmdR��Y�*cݪ���:���(�Q�>%i�>G�&����/�I��:｜���ٓ�2d�-����ud�K�FDy�=4��ǲ� �� %a�,gl���a����Nd�fg"�syFg�z�H�gѹh_%��2��R{����v$_���y	<p��h�R?�E�������\?Wt���=�o�>��� �n�p��<r��7�ChN���Q-��f���N���h�s�I�����T}�:�\��.���h�8��ieh&���<���G���D�;l�~���"rp��CՓZ]���b��Nn#��cs�����x�~n��F���)���u*v���en6�*��..)l�y�e�����]aA\`��-�^ƨ�
�Rq��u��m�d�k)��h�)8�u�ށ�p����Ya.��v�T$�{��L���72],P�*"�bZ��p�2�'�+3.�ym���D�D��S��L��jw�¯k���W#��H��.l�߀Qo��-,��x�Kk��O��<�xj�˿p�B�y��O�܋�{�ĬW���|adlL�_D�"�e�'�Pc[��[��Ofbĺ�3w��\s�U�e�a~��+��~�����
t;�����w��)m��v�_�m��{��7��{��"�q�d{Y�{�NJ��:�^���(��vy᱗~��r�n��s�'@ݛ��_�y-nk���Ҹ�u�H�?IE3��:���Xz�ښ��g�Fu2]�����a�Z��#{e��v:_�_�����5����� 9B_�.V{;_Y��'�q,�7������~�r@��-������.�3N{�FA��;�K��}q�33w��n��M=���c�/L�v�~ۉ�s^��Ȓ�뛨}��cb�����#�庅啓�M�Ŕ�%�Z����\S������|��'g�������"�~����qu��{I@Yo�,a���u%�ta�.O�4�.���pn��t/Uo��@yg�v�xd����y����
�J}y�:S�c4K*�vI�Y�Q��SQs���f���fH����R�v�5�ܲ�^�[!r79"Z�v�-���F�bg�V	-��+V<y�z(��\��s��ۤ�8* ⸱�w��"����8�pZG�	V�8��UT�2�4�Y�x���Vؤ%�,�2��-�P��)���t�&9neI��v�a\t=�yW�αP���
#'
ۭfr���;���pPl�D�v(����W
��K�=%�G��9o���s&B�"r$z ���ݪ�p�U�+N�8�Ȩ���L7�lʻ����wnf �^a���U�'/��$�r{o���=ӆ
.�(F��wI��,J��p��t��|��z��᳖��J��v�sA(�6�U���	|��2��W�K����
{{�����
"MN�."Nu�9Ё�oX����=ƇmC3��`���s�S"LC���}�f'Ύ�,v�"\ݝT�%AV�m^nvfl�I�!:�ق���Ϋd< �D�����-=X�����0�����;�
��*^��
����c���|��]f��2Im]�_S6����f���i�s�;��M�Jwt�D7:����[o`�Am�^ջ��$�N��<(�%������Tj�C���m�zvN,��J���&��;U���F�v�`$��+�Vt��2��Mk�VTm�տJ0
�Gw���u�A�E�n��ʻ��)����*�),��ʴ��AV��T5y�mLx��tn�>r�z�+U�\����%nd��:	!D:���,�x77d���{���JW#rI�k{��X�o�v-��<�������-�ʀ?�M٘
��A�����R�t�.i�Uk%;�jtӮ��@v[�G����W�A<�-Ĳ,c�whǂ�|��Y1/i�ᅷѨ�ss�Vތ�%o7�k.��)��*����RoaK��+	���]�W�v��Z����8�ڡ�e��pء�Xu.�j$�pa��n��5:P��۶�e���[�Z�ҐYoF�0sR�ʘ�+����:��]�$�N I
�Ԍ�j�㪏n䚜2��(����u4pN��G7#�*��������yLEaʬ�&��@�o�$���[}�e�/U�(�C��� ��^>�i])t�f��{�����;��*���3v%9�.�cyzs0�r:�M^��+�
d��N�R���ɤdݾ���P�א�ݞ�����P�R\�|�L���O���W���3��H�MB���s8��Kā<ٖ�5&VK5��_"y-�Rd��3��ŪJ�t�V�'D��>8Pp;��9��G���&uv�&�f��=Y�!J�^�
U;�3i|D�b�;9d���{�	4huJ$cޮÁ,�·�������Ǡ���/o)��V��[y�;a3�&�����bmq[��V��fG\�ki���i���	���Πj�D�/	�7��6Ǉ9o��u		s���2,XX�t��&�t	���YްtĲ�-|���j�S��:�+[�v�DQPV�!1!�!�D�g�9��:�T^dG8G*��TR��I��Qy�*5#S�QQ�C�9YTU��I$Es�f�99r�"�*����A*���z*9.�%QntPX\�.:�Us��wB��Z�T�\*"���AUU�Q��A(���sWv��h�Q�G'
���p��"����"=AP)ED,�Twq9J5�(rV��5�ys�*\�u��r5��"��\��]O$�5̽*��ȧ]�z�y��:Q��ft�$��$��t9˫�8g���uĤ9T�J��N� ��$%�ED^g1J�^eW#�Y���"T
u�,�6VN{#�9$�C�q-=�zj ��*��Ȫ�$%�q��]-)�t�r�I�A�P  B!T՘��ڏ)K�ˈ���2�'����k���z�Ň��j�M��r}l��-��,G��������n%K@�ȯN�,�cP4ٻP���\n#����ˇ�p�����Q�1��r��E��z�Yj�f��>D�p��Xx}��_����鿴���,�Y�g��ֲ�Y��|���BW�r���]���F���}�t�y�=:.'҆�N��t�>�}�F�o�X���{o��%U�� o����~��rUo˰��Oi���)eS_d֖/��]��1j����U�
�Dryc�}Oċ�����9���hvyu�b��HvOo�P�n��Xlg��o�J��:����N�ﳪ���iQ�\���)�;�~���lp���a��a_�q�6~�^R�g2��/���1`z"����L�ڨ^=/��:�����Zؿ_����Y���)Q({���ޞ�F�̛и�_���G������S�u`�q���Z��\{���ѕ%ʺ�޿o.�M�Q����l�/�Pz@�u�h���<��k�D[W�|�5:p��(�m�i񘼔go͘�˂��{��S�}9^��A�٨0a�*N�V��� \{mV�΃�gk�[3F�s.Hdҕ��f[��5cz���x�NxF����3�d�f��b�F�i�>��k����N}� �/�V�]��3��m���5�˺���N��������3@z��V��;���E�y�R�ь�$ͫlL|��u1��G^GZS~���_��wi�7�(����w�̃��Ah��(�ʪ)�W5�A洺��s� n��@u�����<3Ԫ�sӴ�X�|����"�׍�s閏CP/i�'ת���Q�=^u�t{�w��zo��kE�{ʯ��.��ft ���#���mK��Ss[땩`Ze�'�3�����D_�d�n���8��P���q��l��<��Y����r=P����n�f���\e�'��Q+r ���7,+ͭ6|'�e�35��Z{�����E߬����V��ק=e�f�I���������7�%��"O�۝��;���N�Ӭ�Ectz��O��j�3}�r�˿`���!�Ϋ`��i��eX���.<���Ih���C̟qag>Q2�pCW�nzsϫyr�3�} k��@V*��#"=��^�G{m	�N<�W�}�V8Ǿ��� x�hۭ��{��ʲ���:�7�|�Df�gK�K���\w��1�\)"�T%<�����pﾙх��Q�u����L����	���w�5���7���������d���W���ݾ���	k?L� �gk�)mԣ�_�RZ~�x艪ι��Zr��Pԑ�����l��zs!�ۮ�<�w!%i�8������o�E�N���x�"�'�=��V�!T����ǽ�\s`�6d�<2N�B�m�_ ���j�WIJzs�=�E�� J�>���}뇄�>jW��S� jw�3-ӒY������y:,�>�ĥQ��{l��Q螐;�L	��^�y(6qԑ��{>�V/d�x���o������|./��W����v�1��]���7�͠��:Ox6����֥�{nbV�w.��}hp���1�=�z���W�<�1���%�o|�1�B�Y[Rvk՝�;�V����O�}���+t���:�$_�P-�{���u#cޯ��{�8�x2��C��{���^�i�da�W��-܀����{"s��&��[>� <K}w�;���s��=�����$�Xw���DM9�;� �ӅK�p��F�ʫ�Ev�q4"��V36f��GE)��읜�<�)zI0��C}����F�����)cg֊������3�Ϝ�E^m3s���@��.���d�gļ7'�U��CW�z�O�It��>/�s']�:�/yd���s��z����
����/mX�D�A��7���N�/,'}�u��d���)�)]J�{����&�*��*��Zs��M��Y ���A��-u^:�a䦏�M)<y�ˡ7��z]���ו9ul*M�ːܸ�	6"un�ψlV�; M;J�}������մo&;cZ.�9w�+��@��&�]9�������u���0�~��T|��%�[�]����BN������c�%n�Țfm��r�=�{�M���k�{��i��M�m�}��ٴt�q�ԉ�x4�@xcY77"�����1�ݢ�dL�f������X|�{K}7�S�@�^�~7�lc�xI�H���z��x����Yę��U������1X��޿�Η�3���r���XՐ<K.�Lo�d��S�>�ė�c�G����c�׿?�<��8,��K����7=���L��Ż��;W4#�{Χ�'���?C�v�L��z|��_��7/��G�c����5'�T�S��}�
�_[ެ�!�O=\@�ah�&c�C�|X�<�z2#}�����:�%��)��;�R���hLŸ��=ԧ�[����n�M���5�j"ߺ������W�[��E?_���/Y��!�oՓ����=��`S����M
��Hͦ��z�Q�i\M��֑~%fT�ϟ�B^��U�~y�<��̾�S.K@��M�0Xu��As�sai�R�_���%%�w��{wn�*[Y�:zԳ��m��n"�R�S�������j\���hky_����Y�\]��J������Gh���E[h��_��茔��Y���XU\x�4)�(KO�G*��#2VI�Y�1��̜��bv�X��A%Ds��cN�1�Kin�=~z}�;���y��f�h�uNH�-����D�S��ѐ}+N��+;���h1�§��G.��;����м莸��W�.=9^��z�@V���ĢnKGML>��0߱���i�2ח;S�+�%��҇t9c9��8�׏���C��=q� ����ϑ�oy/I�Bk��|��];ˇ�����x��i��U�;��q��~�,�yH��˱�V�!ϐ��yTnϽ;{�u�,!���������i7���{���~-�ׇ/UE���u����4�g������^���l��D�M�;,e�p;ɞ;��t���,
���\�8�7V���,l٫fr���p���.����{�gO�$���JN�q�ZU��V��r7�k}��z�O�~�Գh]�Y~�/��7��x~��}�Wo���=�rO��ʦ2�&��(%�Ñ���j���>t{�x��$_٭ߙ]n�+~�C�����nK�yb�fB̲���z�7������&w��f;���+1���㑾�y�߯��^Z=��Sl��L����Gw��oxu	)!�le����,Z��'����/���^f��Ҷ�C�mŠO�3��Śo��68�G���.t�K+%�\ާt��J}�e�Z�"�óU�;1W,&,���ft\w�P^�jʤj;|r�A��ǜ*�����%���#_�/U��p]�a��϶������y<��r<[/�/}� ���xs)�k#�37�fp���*����i��7��w��F�?+�`^��벡��}SYٵ���,��f�3��>�g��!N�e���٣�+����N��w5��w���^^K[�|���K��caO+L��.����Qr|�Ѩ�j�a+�a�"�+^eM�/W]��s�g��1��%z��C!��9�#��g� �r�B���10��Ϫ�ez"�9xgk{��dǟm=9e���c�ԑc=J��!z��/G�@~uK��k�w�u0f��{qב^k���@�>�И�t��v:a�K�p{�yU��G��L� ޅ�������Ӻ�>ќ|G����ne���y�B��ղkK��<�_�1��f����xi����p�+�gGu��c'	�|T�����r¼���#'|f�^�&�K��zbpe������n�ڭ��U^�9�~�z�����<m�n����q��Yzs�>gnv�?^mh��N��#y���J��V�1��Y��󥎸����m�%�k��o2��^�t��O��񻬒v��e��!��i@h3o�54�#G��3�#%�Q-�}V,rŗ\�oM���s�l�*�5I,(f�����joI)DTM����{MtJ�V�γ�T�����Y٠�Z̔�dϛ�,����N;@��2��V&��{l1_��D%`�W�s�ʲ/-���Uw�܍��8}��5\v���X�$g���D�/V����.!���~z+����ˋ��8�';\��afT ��g����e޾u"3c9�&�Z�YK�h��8^:�y*5�ۚۻ��Q���X�nIgng������1]ÿ�g}7��7���Z�{K��O�_E=�쓁�x�5[�욕9�9����yuVl�*�g��L	����S���/�Շ���s�H2R���Ʋ�<��y���E�x�6��,��d	F�z@�\U0&����A���m��g�M����;��CN�WWޑ�W���@>GǴz��?O�ܼ�ǯ�f:�K�GdWR&���L!�j�H�~�u۪�Q�}�-�nF��U�|$/y�>���G��ڇ��G�B��y�!�}뙀��򬼯��O{}�3�rLx�^�Gֵ�K6dd�Sg=�@���+�����pl��U��7mz9�ܞG����O_� y�FF|_W����ς�~6���߫�x�k�B�zG��Ş��[c�g�u��u?xp��p��kVV㬬�p�>JJu��&jR7�u�U�=7N#��w+��_��{�J3x�lI>���J������VX�#��}:��%數b��M�Q�]�v�̳6�DS`_}xHᖤ���6��3�5|6�*Y���o���3"k~\��_�i����S�	�n��~;�
���?M�=���#~>{�Y���ȿ=>��Q�6����,gĳ�f5,v稇Qr�Ȩ�s�<kuw��%�U��v�<�<��9ب��S70��{�C�����$�����#Ʀ��/����n�"��_��w.�'�r�0j㩇P�Y>�\(�:�>~ڱV�D���$>8��x�?�am�VOt�{�яޥ���^��<�ۖ��z�1z��'>�P_?eؑ~z+AV�N�9�!Ȟ��g�b�:s�L�;q;P��g���mV��gNS (]��b����9�`;���q{�ggW �.����kGa:s�,b'K���
�=J��`o������=SL��Z7���S�A�Nz���9�D�r���H�.rp�C�5��d��b�\��r|��Zs��Ƽ���3�r�l��Ǵ�8�'�y�[E�(��˜�*�=����q�󩛜9�����^K�Χ��]P}g�:2�^g��^F��܏{���϶&Q�>EK�؁��q�N�E���'cη��ˏe��)Z��9Kpq�*��<�1Y���/}��d�R�e^F�V)�-��G���	/�m�amިa3����I�W���_aL��*�Z�՗�Z�t�
�p۳��و�-J��A_M9��)�= ���n�r�p�K�E��ʘ�zi�c?^�މh��W�_��-Nu���k�������~��+��%��<�g��@�zQ;�x��w����@~��{���"=�F�=���lM��^E���x3��{E�#j� y��:sW��nP;�KGۑ��n1*��^���n� �y����Ǩ:�8��;���_�L�K�@i��0Xuj�T>G3�XZs#U?�\����=�V'�T�����Y��gx�q�Oq�ˑV꜐h���dLS���9�/��qL�� ��3>�_���n#���~�U鋏K�霏T�
�~܉�g�Q=%�Ʀ#��p$�<�|�����&=IVѽR��}O������ߦ�Tz])�S�z��ːE}��HYc^{�S9w�뤕�p���;n2�L;��t��/O���~-�5���E�����.�xNʶkcۻ'+=�y�FC#��N�%�3ax�f�C������ˇ�7�~�E���m@�5n��tn�^��e��߆�6e~���%��b��s���S����Q�[��c���8�V�;����I����M�OMj���5��0��.�_M�*�wսg]c�{Ma����d'_b#I����akc�q״�b����B�9��G���^	�e�M��}�0���{�9G�e��p��ݜ�q�a�e�]n��̉nBGa꟪����2�#��_TMG���9$��������d΅�d�V�~��c���k<�ڼ^������g�xs~:G�ռ{ت'����碻�����ʞ�S�k��@��Z�;K�i��2��1�?e���^�#=��V�G?VZ���b��{n�yc�m�oMz����%z�u>3���3���a�߻޿q��/�r�^r��Ѷ���C��W�}�C�t������$���D�x	��\;�2���P�n:�\<��s���Z� q�y����g,���6�s�7{Z=���c�%Q��2M߁�����4
=�'��ױ�N��ͅ�̺�u��Ey��&���i��[����(��Pz@�q^�\�M��v��ޚ�S3=SN|�َ�,�^��ؗ�Sf�T��t�5~�p��|K
�0ڕ'�ރؼ=�>�NG�u���Z�}:o���R�ݎ�Q~V��]/<�Qs�;85z���3q� �����5��6��{'{�i�Մ��wRӐJGv�N{��i�nx��H��}��D|m����m��cm�o��m�kl��m�cm���`���8�`����m�o�cm�o�cm�o��m�o���6�q������m��`���cm�o�m��6�1��\m�cm�q�����cm�ox�`����(+$�k:��@L~k�
B �������-s�}_ �$ )@����@�PP*�@	 *@
�R�H�

	�5R���$����ETEQH�Q*�ѪP  ��nUJ�ER�E$!"��J�
��IJDJ�"EB�HU�*'�� %�M ���*e�$�d�f5Z6�K5Cf	T�"�T12H�  #p q�lhU���h�AN�
R� wҀ
 7L( (՝)@
Ύ�	�E�*  �  �D]���Kfm��&ͱ�b�%S3l2�"RVڨ����	
" �� vUT]���U2h͵��[X�Ɠ!)��f�BV3*6�iZ��*)@�$�� ��!LmJ��4L�Ҫk͆���i���l��"Z�l��aU�6��mTcT�H�����(	�j�@��ѥ͠�4�!�F�J�Mm�R*٪R��»XDh
�MB�  �  ��J�kd�0ʅ#0iif�ګe��mU�d�c[*QE��j��Z5T,��J�TN  ��JQ���*j̤6j�ճMdmӪU,QCD1��
���m5*�0���� p t��`�h����b#Jԍ���ԍT���V�� ���� ��[&�J��
�5hZ�*��m�����ؐҭ��}�O�4   ��T�	�ɦ������&"���$@�����&�a��0���z���j?Pfj�jB)� �$�2�h A�� ��J����      i�*��`�� �0&��h���/j&EtGĔ�/0�"�I-���^��UHI�EPg�! UG`��!5>D"�"%w����~��#��.��a����Ɓ��	�@�0�CX��!X���XR�'ϯ�e5Z(��["g�. �fO�k?��W��Y,�}��7�"���P����Y��C�́|s@�5�i>��zO�&T�4�i��V[��A9��[�0�/[{��8ۣ��;A�ӳ��.�T�`
�e�i�۳��i�.��j-뼦N8p�T���1A�U���Y``Ш�R��R�"�r8a�Y�Q�	-�i�j\w��z��ihg!l�	��S���SfB(��UƏe��vz�5���4�[$�n"�*�Y�2�����]�sQ:��9��U 0*���;�3Lۭ�ъ|��K�W�tV��"Sm��
�gx^Q��+�)*f�ڥ�HwC[�fe�@�{��Kj�[�O��='2�`t��gP�DS��;����]J!諬��e�\�n��2�f�"�<!XE�3s4̉ր�&1k�kp�AJP5o6���)�W��B�ԭtS�hn�a� ؤ���F@%@v��/fYȑ,^nP�,
d��&X.ɠ�Ypl2�r�6���OPՑ�m�fMq1���k1�1-�Z� �j�4ml�سV�b��i�ݦ�n�i�����a%��dx��Z�l�v��+06fh�ة���V	�j&�m���s�lڬ�K]<C�+h���X.�l�X,���J
��ͭ�nT�F!Z6�=˫fk_:X�;s/r��7�y�&�����7����i��]��*��(V+DcZ���+j�\���Vn̠U� 2�]�v�ɔ���oP���1[�(|o�����-��kpS�\r��e^%b��5F����I�o�F�l{4���(C��ȳV��U�c�*ˬ{z���D��Q"��[1V)�\��y�:�v�s��V��;,%}�{aiˬ8��5�M9!�ú�9��������­TN�Ѻt�1#��^��ZU��4]�����}��1x��kk;*�V���R�
�wU��*ՓD'��Yl�d+*�]��x&˹rQІ���rai�b��)�^�ݸ6�ϊ;y/��޺d������2���T=;�`g&��������v�w�S2��Ҹ����W&=1���
�YYVv��8�p_"�2۹�W
�yt��9�ʼ��ĥ[�!T�,M�j3��&F�&�ɗ�Vvb�Ir�����D����\R�\�C2�/�� �ئ^ ����Ȗ^*�ʆ�n�GA��sϘ6/Y��8��k��uL�[vk�p	>X��(��<aK��
w���<Wɣv�;���s��l'�CghwǷV�c2��vh�T�\:��owd7���;�Ps$xRˢ�+����9�q�)�T_	]9�<�\���_�]%Xmq�y͢6���W�Z��F�"�2iF��+Y�).�t��fnn���	WI��}!wS5	@%��J���X�;W
��ȯ���H*�: {JlJ��:��4>��f�d�@��hTL?�]�"���#��Hڂ!��s@��62D6��	�v�~7�T)h��ԉW*��7��Q���R���U�3wP��f��n����G+�[R�����=�n�����wn�[��I����ꂃv��� o�*ő@uA�ʼ��Լ֚����^�4�WC2���wN��ُl��[�ȴ]���-\p�so6J��#�|h�L��urj똫1n;�r���*�	�A�)�2V��:U�[��e���)n�H����.�T�ʆ�	�*�y�51��/�I�9XFU���7���wa:5���*#����8�ط�j
!KsDN="���Rw�o6�I'Vc��K��Om5n��C�Ygz�RO�4�ؔY���㥂��Ŭ�e��2`wLc9�T�{v)��+$7�c��E����ej��Vt�����(�k�Ij �2�6�+V r�AQ4[ʂ��qȨ$X��<Ì1&i˰�Ӓ�Ӕ� M��R�HKo�%�v�����C�|�g�k�u.�Jf�N�#X/mG�{�S5�����p����f�FLޮ$�k+v����˫5����l1F�*m�+j2�^�;{Wy�Y#8�O^�t4F�T��3�.���b-��(�>���6�?��F��m�5r�ujfA��wW��\�Z�5��E�^��n���S�4*�{1T.V�Yub���(j�Ӝ���r�����醕�ͷ-�n�ڲ��A���u��0��kK�t�uun�F�8^2��36��$ӫJ�h��&�F�`�E��2�M1Y��:��,�S��'kZY��I���33r���1R���eՕ-KsTٵ���cB
&q��h��m�bm57"{o6�J�nKR�Ł����y��+]�4wn@���^�����̣'
i
�4���6��9J��Jw-�(ʁ��pKY��wyYY1��N}`-34�+�襨�Vv��A�tQ��(:������9�W
�`��x�e�Y���a�A45����5�E����� ��t�[��HQ�*V���D�!��/��c!�n��ÀN��x.+"9�< ��,�U�a��H�3/y�N�<��wp5���ҷ���.�s�l����x��w����[W�<Ƥ�d�Y*� 9�*Pѕ�1I���`����Z��rc�5�Xh90��Zh�~�YGr1�wp��XRRЬ�O�`?�E�a3*Rn��r\�e�J��ر�V�a�-�B�Y�`0��C��aSx�ᰰ�*�v+��c����m4��%�iȱ��&]1k"���B�XzM�6�M�w45}5ZaΚM#�ѳ+	*�S��*ʔ�Yօj�\�:���ל�[L{yS��a
/Nr�� f�v�:%n��vɧF�Ui��.�9�t+E��]�wY�Pt���thE��ݴ�2v�[�]��q��@L!`f�Z7ٻz9�!��\�bC�ie[�F�]w�{Zo5�:�`�A�$I솄X����#�4��x���wm��sn���4VJmM�v�wo �in�"��8��ޚ?2
2:�F�L���o/j��c�%=��m�����;ky�BK�wI�2�e�x��o)��b�+ݫ$�m��T廳��(���f�����ŵ�M�_n�D��-^�e�l�
�v���3YA�Y�@�;��b�7N���В�kC9t_m<~��YW�j�BJx����B��Mzi���ֺږ�e�ѥF����2�*���x�K=��������qW���'�aJ��JIr�ŀ����7��D�G5��#}UxS:�'��]������T�N�+Z��WMLX�8�����V��Zp�.�ɧC��r��k���+��e�Y�w��ʻ�:f��wh�"*Ef��.�2�f��d�jq�@���)�f�E`��x�m�K0h�M�7��2��Ѧ�`3`�^�,�z�;'/Q�T�=�	k����"��FF�5F�R��gi짱R��i���SVf�m��Z6k��jr9z�6�jY�ON����f�yJ�m�0$��9e�Ãw��/i�,#2�]"1m�JK��Cxr�/~������/,�8���:G�/���i�M/����#B���/,�@1�r31�9h�d�hly���-�jh9G�p�]սu,fn3�/�;��4�G�j���Z�--���]OS9Cv��+$6��أ �����p��W��O�)�o�s��F���Ʀ^��wO������#��B��U���^��"�h���[{ch�b��WW�=�5�L�5چ���m��>B����y�th��f�J2���kW�V�^�݉����N�ѭ��j�@tZ�A{����V�rȥU���V4��9�e^�褎�3Y��4�I ��sn�&v���ݸ�:']J�(����vn`�ǪeM6�ի�e�3�HZ�����/!iYhK[�t�'B�ڊ_��Wi���e�D@�-cԎ�ڳ�72�e0�[���軠�)�&��m1�wt��^h�"�X{��nk�v���4�3���r�b��.��n��x�N�n����
m�N�Gk.�[#���$�nd��B�/�&�v�d�əyn��yt� ��'s�Nu�n
wO�X�tJ�׬�,�ź��^�|Y��7��|m�W�s�ǯs�"�=�p+4��*�s��Z�%�I(�;%ͽa<��E	F��tn��6�c�u�ܶ6� cЩV�5hZ���){��u@6%���Nh����f�0�1*���b&ƥ���<m��8� �XB�{I"�DA�p f]�
�Xi�]�x�S껱��'����،�n^�������GM�����s0#'�u����x�%*	 yu�/ �"|vv'+e��`Z��B5a�[w��L�t�;��0��|�V���{Y68���䉕�6�	�^��԰b����EŌc���f�Zz��O))౎_�%��=���7�#���o�^��/�[֦c�*�3u{��FyTn����o��$n�|��%s��z@��L��,��6�Y�(.0�Ǔ�s���VIyx����g�P.��r�>8fW,��n>�7W$y,�<Ε���b�w=}%u��ӹ�Rpr��ύ:I#[�u�Q��z���[����º52�v�&n<�6���&��+�D���}`���P��!\+hv����R<g}��mW|�څ����aʥ+��)X�iV��W5����V!���_��ܾa߁7W��+
�5�7wW�י��
�,b��u!�ћ�}��oi'�ml�-���cG�h�3�C�,����S�Dx:��H���|���Z�����u]<��Pgm����a���4̓����
B�M%���
�ǣ��<��Oh㙦ժ��N9�b1��ڨ�[���-�^ɤwi9}�h��-�U���tM5���*=��{I�4���)@�$�phO�j)��9�Pv^�0�@�qg,�Γ�z
�Y�rc�"9�ٹ�o"�N&�\��q����Q�+.�ۺ-w]���J��p>��F�y��U&b�Ҙ�%���읙��+�;�m8!;}Z�࣯hNo��"c�{Նra�$����)�'Y�Pn���y�eM"�zM�b��lO��0��4��殏]vE����+&&1pl�w0[��3H�\�\�㢝婣hN�h�[A+o���rpEevr0-c��)�n��(VR��t{9! {@��M2x��B�X.��n��s�-2#7����m]^�e��>[�T��>e���	��iK*�v�5utLy(��Q��:�`y��5�+]��ׇ�nYNֺH\Z���ٶ�=��ȱ+�+��y�M8��m���e��*0��4��P���>�4!]�L�[�w	�HTI=��8���l�[ �7���7��pϠ���w9���/-vP
�bY�P�-�;��o�g&�4:�7�3����YJ��-%J�N�7+�$��r�N����"#�ʼJ���Z����s	{Q�w��Wc����׶�V���귂U�/�W�wBY>�O#N��ӊJԁ�{Xcvnfva�pdv�̾X�fJPڶ�92\鷯k. �P(�So{!��7�sV���:���aSZ�o:U���Z$഻͸��n�x��֧�tG�I��F)�-��nu2t�;�A5�����oS�␾�,b��iu:5[$�ۍ���2w���c�v·:��ٓR�K<֝r���e���D�zV�p
��V��{ϙ���Wf��qO$�OA�֬%��R����֐��5�fJ�ˢn̺\2��Ngm�*��8��LoGZɼ2�Xe�<��=�K��}{]Y���.��L'!�3�LRNbRiZ1-h�X1lw��)R��mb}�L��+��X�,��rW^@S��-U�bO��]��d����x����y����zηI��K]�6����K�`ïonv^��o�PI�Ob�u���F�D�׈mx%��]��wkk��5��^�M ���q���r���ZT�	�sȦ��v�+)��ڤ#`�]x
��Gq�Q3��g��M��v�}��y[��N�t��+hN�\EXU�f�J@JVc�)�pkʕ7�;O[4#N�Tz`P�kxr��-d�=`d��м=��5rRM������
��g]���ӛ7o�_��M�v��yB,�����T��j]��7SPln.��
�ڹr)���k�L��LJqTP�\��;
�z�9� ;�ңP=�&Z�\���M�g2�*�N
���e����npD�1d�Ue�����P%$��e��{+U�\����pri�t@��$ L��G�r��YX��ֺ8/+��p���D��y>_IF���2�� ��ⷭhv����)s�Mcˮ���%��:��$v�+ʘf�LK��2�t�Z�vة��aL����/��B���jF��S���=׍��!�����gW ��^B�b#�wF���^�̎__&�r����v٘�,�;��Tdh��h�o7�f�Ь�E�^hR�E_PE�]���������$��F�;�[�hs��^uw'3��ӂ4�K��#�IԜK��jol�D�<���fݝ!�1k;1�\���RȞj����<��^�Y��Y���j����/h�7��e��$�V������o��|��H�O,�%\�c��u�Owca��_����؆��5��o|�L�=����8�ҙ�2�w�\q(���?�}c0X�y��� C��ӵ�2�+�Vk�|��N�f/���gs2���%���h
1�*�)7v�r�v>�h��,ιY�;'����qB��t�ƍ��w$bVP1�T��F��Li�ٹGEM��m��PG�*4�5�%�:�k����o[�V �:�'0t�gH�t�wc�L$�ޒK�4�}1����3^+�0cو�XwW���F��yu7�C�Y8�Ĭ^+��3yo�u�ʑ�EbyӠV�ř9r�����Ȧ"�2$�Q��%�v��tm|��>�ca�p��ͫ��m;��K�!���P�2k ����:C{���!��+woP|A�J�,�.D+�7Qt�+w���gK���@i �ㆣ��F͉�>{�Vfg�#8N��fD.��d�w ˎ9/aɭŝ�W�4[��!�.r��7#(neaJ�$%�V71�V�5\�	V�6����|�7� ��"�g�u��kU����7D��e�mI�X3������H�.��2�HRX�G,u[��7��4�uƂ]�
�X\'�r�صƮ�u
+<��x�ι��W��u�n�"��4[��t�齍��0�����ׅ.�����xxf�e�'���6��t��E�B������m�ʁ�`��2ܳ7N����8e�k�0��;9�cw�:wU��%�mۺ���8S��鳄'鹭��%�g���)om���5&�sd�APW�WYxv�j�KDXxiB�j��N6E�j �˽�V�כU|^�Mf��c�n�d-Npp��\''VjEJO�
b�š���K�����b|�>�e�µ�)e��N�q�������!�Y��X]��\k��"�ݤ+5Q�j�'9#P��W:B�_�2F6��u�C�y���y�9�z�2����v�G���w0$�Q���E�tR(ng_.=�[�"=����3�@a���ť���g`48�&ʣ�RΫ�'*5���$�����r��F��V ���K���h�Ӷ�;gAu��r�*�oq����!z:o"��_�0m���8jU���oaç6��wQ+dt�y�91Q�2�Ć�Ý\��m:�+��@�]�Q��%��ݜ�2�7R��A�}W��8u8�'��M{��Ȍ����J���-,٩R,�I;a��t%Z��f�-��;X%V�&��x��K��U�J��9�Ao4�t6��}�l�#��ݻFD�	���N�>�0��[ئ��.���l��6�k|�2)�vNҦu�|�ӢٗpZ�c`���E[�%8�q2�vK3_D�΍��i�ܡ���8�6�ɶ�l�F�#�㛏l�#s.��ۑ	+t�=�'#ک��#&�Ӭ�&��RI$�I$�I$�I
Qʘ��䠸d�[q�!ql[*Th}�Vd�{j��e���Dk�v;"��el.����$Rl�D�NmA6(�݆9;s�f��:�x��;0-4˹��h:�b�s
���+^vd�K�	2I$�D��I	�Ibf�a9�����rqh8�o_�"s&���=@�G�aC!<��7�rIV]{�]�S�bm�t�N>�6���+mFm�2K���ܣuۭf%,�Z�k�Q;���ne���P˒�J��@���Up���r��ĉ��U���n��j��s�]���W>00s�6����`�>��8T�[���l-�D�e!GS5���17凕���m�W�q+6�P�R�Сe,��1��9�X���R]�ɖ4�m˹�h�f����2�O����Y�A}'m�I�RZr.�
!�{�n-7`�0��V���0��1�X�0T,�����x�#���Yj�Vv�;��J���z�P�]���Λ���-��Ʋ	w"��i�����N]%@^�$*��f� �i���!U�Aj��e�ES�n��i�#hu�l#Bb�>}�*�k]Y����#Z����S���up��n��wC�vG���D�[��k00�.u,���]6Z�*75��ֳ�黡�8�� �3�MN-�'j���4��_ӖG�Fb���X�7��)�[�t��N{��%�����ǆ��tZ�7 ]:��q|�]�e໹���r	k3
�m�Ꝏc$�(��.V���|M0
�=�;�c:�m�����q/�qI��p�L|s:$f��')����V�E�˱{�MbC����e�ʺSx�T}j)�m�7��8��{�e��C��u�|���P�%��m��A�ѣ��	�
T'��[��dǱX��x�1�~K��F&������]m�}5cra�U�6�2k��'Ȭ2>�GE���R����wm��P981]���U�[��>�o-LHL���m]�b��[����g��=�fM��U������N�-�y��Ω��9���**���V���b����#3l�i�����,������cX<�,�P�Ȯ�&��i����AZ�����v������R��1ա�`(Q����q�b,J�ێ�m��(��Qzx氨���/2]��O�y'��VPNp�y��
oLtu���3:��{�T�B[�}�DKyw����-�2��-�vȾx��:��R�Wug]��FP�i� ��rH��q�\��T�u�t�Y��� ��f�d�7��\v�c��5	���N�4^�,f��N� Sǝ�)�iՋw�	�Y�Q��d��[QP����cXƅi��\:�o2\�Ԇ����U�=��<Lp'���*�XZ�op�i�K�V���3��T�h���-��[�N��כ}�\)w hj�g:��)�v�p��Ėf���B�Θ�t���J� ,���~`�b�A�.먫|�c�K�Xy�r�V*�ֻ�:�8���)s�j���4ٹ�Ü ��3u�����6eY����c��nY�)^�p�2�`*�Y�����d�����a�-�	G4��Y�0�.q3R���[�%a'Yz�u,���w�M�k��[�3����TLd����f�{�v�g�f�ȑᚨ����Ϟ���͓/e3��q��]��I�=�S;��dq���h�ۑʗ��s��J�b�i⣳v�W�r6v���r�sz������a[�1Z��:�y��)��ݦK�Շ�!긱 ��>��`��'w`͍;�I�I�(����2ڲ��7�m�D�Sƹ�L��6.5#\P&Q_^ nQ4��P���*�ѳ�@\���7okn�M͐�.���/�K<7��"�N��2��ey�Z����#3n�y�p꾣�Z�Ք���$�E��%\��r}�ݫ
i>�\�k�^�<�kB�t��Z3^���
�n1�;鼎�#��u_Giⱼd������-��c/s��W�N�c$��GS�֜8݇�[�.[k-���1]Y#왜T3�Y�#:�v�u�doU
g�ޘ�����]�Y�AR�iB��d�V)��c$���� ��q�@��Z��Y�/��2,5�hС�m�0����,X.d!A>��î�`�V�˭a�8+���ֈ��y|U����	��^���4!EI-9�`��6o�s�'�sf,��Էa[rg%��0�Yb��'�^�p��ݩ�%�l�rː�<����H���*��[��Z��݃-�1�<����ޜE���3\X��B����B���>�H�iu�}���-X�9k¾9Vj[�pͰk9�<2�1�u��'�=�1g;i;���y�B}9L���7r�c��lV)�L]��v�۱f*f����9V��[o����n�H��^�'��ʹ�U�.tG-�ӊ�C}&��,,"�j�v&�K ��kze.�!������{a%�]�Θ����~�Bli7wc�4Vk��%�5�4"@];��.�ؑLP�E��2�^+OZ���B��du|s �:��uWmL�\�ͭ)%�*����nbWN1հ7�e��ڜ��d���y��B:�J�ƪ�JW���49��gq�N�sR���h�ԡ�w*�4��i���ԗj3��+%p/Osü^m��� r��ֱ�d�c���Z{��5� �{��e�P���RS���>Ocg,O��l]긷P�1[�u9�{][�NY� B-��֑��`$v����2o(�d����[j���R�����r�����K��\��iÃ�����nhv��r.inX���Vtᷖ�5&j���5�,�k��E'#C�E��w0f�2D�d�}Se�,bOh�0��m��n����<	�H�4wnDS��	��^�F�%P结sz��\L�cU�q>�ĸ�M䍱Ճ��S�D�5,x��5*�d�̕�V�c� T�f�j��}3C�;Z����B(�^�Q���ƞT�8w�z��"��$�V>]�'V�.E3:�A��gUns6YMl��Gh���c��N�Ӯ���n�������K���=H�7�I�r����Xɗ��ҋ}� �&V&�ׂ��*�]��x���:ՅK�j�9��.���d+8�����홛��'�[5)��v���;T���2W�Y$��rY3	F�@�N9�{�7��T����wK�	�7�-Z�n8f�Tw�(Y�R��"����-�_+�^38�}��8�w��;���J�,�uW,�����BK�G�������[���{�>����n����BI�ف[,��Jy�ۙ��e��n��r�P�F�_Z{����D7�����4w�"�n�/wQ[�\Z����o+��.���_;g�-��DDasA��,���jܐ^�q�
����/_I��_�2<����ݹ}���/,XJ�'���&l�єUn�Rj��t�g�:�����G>�2�{8f�Ѱ,m=8��,��Gy��8�b����kxo3�M|����{�)�����[W�֣Y&��[p�MҬ����.QgV�On��*T�n��lHEx:P��C�,�8Ҡ)�'fK���ؾ�|�a����,�R�ފ&��֤�f-M+�^>�u*F���Q��K}�Pon����Idr']]�0|�^C/u;���p�JȒKĞ��FK뷲V6�����N��H欬�ј��7uE� �M���ki��ֈ�
Ʒj�t�_u �VNBQh���p����U�E�=}e�F�`s��.
�:�U�-Kؤ�z��5�w�r�hl��OS�̽2RA�W�]���'l�X�j�Q�ӻ�M;3����_3\B]u��Qδ�V=s.L�Or��g	L𹗉�tͲ��I5ۼq��=���az�f��V��}��ԄU�1�{4V�3s�C�����}��3K��&�<�tC��
�СS��l���ӎ�U1��'�?]cԂƁU���o�B��?-g
��(Z�w0�t����E�d���ҙ8�{��YEē�I�}���3)� ܝ���ȑ`�kV�M�D�}ʺj��x��7x��kY�м�2�&\����j.��B]i�U���طv`����I�0��]�\�zZ�l����f�[��YB��5R\��(äS!c��)����'���#���v��)u�,���V�3y�k:�3�Ú5�`#?m�^�*�U���sU��o�,	3��%�n���l�?K�+w�ne�m�B�]�ejzI$��b{Yt�w2	�1Չ�"l�it��*_GZM�%R�,g�6���p�����=-RoD���g�l!ɳs�"�˸�����������fK5�Țc�e�Y�Q� w`��N֪�X�o�jZTUx�Nv�S%�:�>R�T��8�o��Y�\��X'1��0�Hg	ʄ��'r<;�ؾۗԐ��B��;G�I�4��+j���btd+$9�	��N⋘qn��h&W$�|��i|S)1*C��Z�;8g�#Y�e�;t�0f�|�Ù�٦�[�]��Uz�L*:(�+�}\m��Z7�+m������t����l��b:Q"#�Fh�"�K�uu}�[������I.۶Q�u�uvRcvQkRWmN}���<��)�;�jMK/�&1����];O:-l��e�:�5��w;/Vi��Sy|<�S$����8�j}���L�O(u[�.�c\j�܂��b������D�/1_�m�wه07���i.D#a��Vp�[���F�:8X:˙�G��Aye�]��h�H��L��q�/��(4I�`˶/�,4E݊3�[m:��oB��Ǝ1'w�*�[ۖ���inb�d$�b\�,�۵X��l��
�2�F3�l���GS����|��Z�v�wGm"�9;w�^���R]V]�
�X݊H��m%ݵ�Q����({U��T���&�VJ��}�̙��@��+]F�[����%^��P�{��,�@���>��vu����)���Mպ㮸��-�G�����#�D��6�J
3eC�Iad*\�5��N��ޕ8����d�Bk܇��w�lO,�/��3*�m�K[\ʮY�b�5�Uv�T�h�eżpC7
����mUr�[�s1Tm�1\\���/0v�TQmi]F�[[�W(��E�Z񟍤�3+YbJ�r�%�,a�����Т��P�6�a���&\LeCkm��Q��bu��k��Ԭ-
��*T�AEL�e�U1lY.st��n����ǚ]cJ(�Sp��T��e�s.6�e�Y1-�b�"�]e�1Kb�ULh�p5�USsqMv�R����̉����M�n�Aq�ڮ�C]��2������m��q��e)po,��qp��wM�Q�jURe�1ۗ3uۚc��JDҖ�AL�W]ʺ�-`�w����Ħ.v�u� �Ko!�]��&v�xc��xb������u�#�E�9�"����ߘ��5y��k}Y�"i��G���r������7�y��7ϕ���c���+�O?zYY�_���/+��&_�C�lc��mP�g�|K�s��O��n��eQ���)�l��3Ճ�q ژ��ca��mE^�q��G31g$��y¿v@��(��u	���`�J6v��鳌��N*��r9�/�rA�<�{��T���I�t�����J���ק�<�䷧�ٲ4V^4���P���z4:�����a�2:WVGC��q�S���&��l3��{t����)n���9��нx-ԑE{/$mVD� ':�v��Ϝ�O]�[2��M6Lm��ǯ�� o-3Np>���E/->i9�y��Jr7�qۚ9��׃p�}�e	��=6�;�=»|C	Y�04�ɮ���Wi]��ۚ�<�1V�����o��U���V�wo��o���W���T�t��Qu]�/h.{z��=��{(���9�]���n�cp���+,��aGG;*�&�
��K{�Oo���{��$k.4�N��<>1؁t��-��O�<��S>��a����z�(lxR�z����F���2����{�}~s�v׉��r���ށ������0zr跾1ܻ-�kW�nl;D�N���m����+Z�l��Z*$K0k4�'n�Q�����p�
ڛ'a�N��Z�K���ru�|HePW�R���Q��덞03�'<k�K��uJy�R�y�N��(��qN�6.���p[�V��X��FQ��W6�*_��
Z�������ܹ��1�oRm���Rgvj�<@Vc{��T�>/5M�;��l�w���r��P]��F��'U���ik��uC��Ʌ`�_I��Y�T�e8zk{�͘m�ui{�s�\*t[��{t�j����W�x�Ͻ�,�Y�x!�Q�f��83���9��{���ӭ��Ů�ۣ]�q����6�G������oݧy�ɫ���<D�%�Ǜ~R/\#Υ����~v�T��㾮�Sua�[y����N��>0���s�l=�A򵔦s���3wP��[�G�kZ���B��ҍ�;y�{�*�qt/μ���þ�cѿPnm`6��m�~v��pq��y�`�E��b`�V��=I)޻�N�tX�q\y���Z���n[��M�i���٘�cz��Pmt*ތ�7˫�(���*Ag\���
�<|��68�B��M�Qä�tԱ���-̭֯潱y�۽��i�9�S5 {���-���c^��=UE�;ӷu��K��'v)�@w�Uތ���5��8�ݫؼ�7�1RY�Z׳�3y[��hPyC7J��G���|9ѽ��m\Z�e0[ �-��W�~9T���r ���A9)j�T7���]��rz�ۀ��k5��S��f�� ���t4�m#6o}�7
�%��C����ʛ&)�k�r��tLZ����ɰ�ų�ո�4�r�{�e+O��2�-��QO§�~�����X���Z�;�p2�̽��Fw���ܓ�s��	�ˉ����3�b�U������3���"��޽I�?i7��	m��e��δ˄:�ߣ�M�i��݁}�\��~uo{(3�:��ek:����;�)�Ż�l��z`aȥ'�1[��Qvy���L<��w_��zp�P���<T�=�z,8�H<�&���g�"��f`3��v��'{Օ+5��b�K�b9���]'=�1q���I����Ǘzw�\z�əƖ�Hqh2G��Gʿ}��ߕ7yQ	�:F�dg. T�Kz��j��1/&6�]�����qiv[7��ߋ3�������f�?1U���m���}[^7yrJ��66��W׳�*��u)��drH�⧩�F�y���)���l�K��F�y����ٛ�hDsY�����}#��#'�=5��/��j�����5NN|�O4Q����z��s\bo�}f�[�U�9��>Xymپ�=���λ�|��?P���˶|�ʭEx^�����K�t�㻽��1X�¤vxnZ�e���"�*%u��Z8���6V��dZ���&+��&髻t�=��5�v��9p9W��]z��:�F�P�<w��W\M�+5���
�L�#N-��c�G�a���ɡ�{��C5T�h=���po�{iژs]z'��e��t����1������bØ�1��]f�B�o�D��`��N.���(��ooW��d�Q��{�?tj���/Oo:YY��\�Z����u�^��\�Tͥ��ew��a��ml}��q�+�g�{�#z8L٫��r{-���s���LS������f��soX�Q��)r��9>V_5`���.�Eo<�Ӗ�CK6V�ެ�:�5Z�l�\�z��7HyJ�)�����;�h�ԝ]�=A�0ԣ��Rg.L�$V��{��[��1t^,ɏ��C�.q�L\~�2�+�"ܪzu���]�	��ͯJ�۳/�5Jٷx;'���\�;��c��M�3Y\���ü��#r;7<#�jS�����L�i=�%�;xN��\HΘ[�J���GV��SK�r[\�Uer�{)��s�^��;=�V��Q�-�q��}4�z�b�}{xk�<%ķ1Xbb���X$�J���u���m�,u�W���=���C��К-��o��͕x.q�9"�^��f��;��wWU��������!�B�ք^�[��dT�������7V��w��U1�����:۽/}���nGn�˭Df�l��(���܇ّX-�d�N}$���P�/�\�:��C6t�$��׬�^���.g��OEF�J9-�A�Ih�V�	5]>��Koj�o8���~�1�?O�R^[5R�d�=��e�Ed4����۝� R�o��节��߽�����C���3�f�?^S#6_D���JU���y�J���:dgա<�8�}y�A%��xg�If����w�qYj`c�^�h{dsݹ�ݫ����&��cӥ���u�9��=�<�w����v�5�����~�t��0��V�c�tw�n:����5�o_�Ҡ5��z;1���)��@/�w��u�DHJ�m�W}&�\���K���F�*M��<˅�#�;�pz�j�������S}�noM��7��V=�\N�߭��يeژ=���*���_6�|x���p)�/j]C�	[r\��Ѹq��qP��Td�/88�t���I�[��!�S��Sw�5�E��gi^�Iy��9��}g3SUQ:O�xӬ�Q*���#�x!GdyD,��y���4��Pb�Vn���P�7Q]xC�O�tx�ꋇ���|��|�'�T�ѩ�s�u&�V�Aݾ^�$���kO�3�m��hTG5��{�c���OY�@wo8��r��k7�SPi$;�>������ЭZ���Ծ�vV�guȫQf�U���x��\����@�4�0(U�Z)��j�Lq����D[H�F���鎗���{M��AͪKs�V���n��
(٨�44r�sr���������8�ꭥ��H�W$��Z�ƻ�mD�Ψ	Ն��p�N�8'�A�$��{G	Qv�eաLa:�;�y[���m1��r�;qǔe�f�����w#)��SBŁ���v����ų3[�%ֽ�=
we<�Bʱ��X��qN�ذ:��<�t�!
� @FsW#�y^��\�Yo-2@uCz�6�=����(�M��_�z��ts2�Z�5��j�:�tC��k�[W���	N�\X!i��n^f\�4���u���N�q�c��*-AQ��h����#���pF]�ro6��Iv�x�5R��u:Ge�vX��ůen��a���8#���?C�ǿ���#�qx�F�H�F���I�l�rcU�01�s�r�xND)سJ��B�LQ�a�[�P`�q���y�2���:�
$�6$%IC6�'h�Lҧ-T��"�ܕv��A�f�ガ�Hb�xT7d�t�2b�x8Tq Di��%�U�1cQI��b��aĘ+Ʊ��6> ;�.����;`�q��$���5xEg�ko3�+l�K�n6���D��^0)�7WVvK�Ӥ/�=��,�]�X� G'I��=sdb��ڟ) s%����7�h�OI�?�av�K����R�×��v��]oF,�*���:j���wA*��x��ӂ�e���GW�b2�㵅m
�	ݻ�G�U��	
]�`|�����o��)R�pM�P��+B���R���[�y��"��ʅ#�#�J8V�����;H�p"��I��2 θ�[6+��i�Ȫ6��̔A٩p*֙j��Y�sw2Ҋ�k�f1�v�rѶ�"��sscl��7]��6��bn3Q�nf"�,bb.n�
�]5ř�m��S���h��X�*�)Z�h�m��a��GnQMh��-���kT����8ScV�6�i�]�k�2�]�3(Ҋ��*����b1X�
��T2�]�ݦA�U*U��k�c�&�m�5�
jݦ2��0S2���6���X�[R�ar�Q�`��e������3��`��Qf�M�.�Y�̩��Z[q����f��mK����Kh������@�����J�I��Do���05#՚u�/�:��oT�'Pn�o�\�&�cPg	C�|r�u�D5��L��4��Ў��Q��jM�<��^O�>/k��i�k�1^Q���t�x��NoU;��ڌJa}��?�jjWӦ~��Gu ��}'��ﾯ�}޴c5�܍�m��?���:�jg�e�ex����U椹�N)�Ss�7"`q{���͍鍇�,#;ϵ�\OJ�C�[�l��Oz�lkB���$^�4v�ٞH0�u���#�%i�C���
�L�o��zj�����Zv�y�P6cb�*u�H�%��OG��<�:��8��6�l,}#>�y�q=��z^�k2��������f�W;�\���E�|��������y�Ri�Q��&�N!ԙ[���&�x2e-���=��� ��뎓���j�Z+�+�<�m%�<%'�~���Ӭ���� �\��<���9�Z�-�7R����$�������D��z��<=�v:�u�Q�'���R���Os��qgX���c���ԣm�i"�:���F����z��m_��ݲ�~'&�#j`^Lvl��~�<*�R�\�[;��)xڤ{����2��-���;��c{{n'T��ݻٷ���\�n��Я���`Vt�ZW]}�Cֆ˽�@ik�*�B+�	y�{種����+0�ؚ�>���݌��b��qx��H���ӑ�t�&�������6��vD����no���haܸ�S�M��S�ӣ,M�ݵɑ,����`�V��\緪��K9]q�3r?
��}qf�ТUNnQ��u���Q�u���kSn!�R7xβs[O�LS��ʑ�9�jK�M*.��ِ�e-|�+C�n�Z��ө�X�{E3|*]%�h�>�S],~�{�F$��s{ѓ��r���w�n��{w}���.d�WY�V���e��~O��7�+���d:���l�QՐv��vj�K��JGu?�j�ŷ�+��l���mv1H�8���������5�L����b1�̹j�{fZ+9H�w��8%Dmݸ���q����%�I�S]�jО��ݗ�㽗���;�{F'�g��������g�y�2�n�ܹ�����Z\j5��9����'��5�+M�yd�!S��y=Ef{�->rI8y����g��{;e��R���ܽ�2ig��M�����Z}cӦM�N�:@�˞��g�o,�̆��S�����?}�2����<I�!�Rl3�c$톝X���w�d�W�M�Hg(N��G�U�����η˥� �=��>��wa�%�̇���C�C�O~2�!�ņ'��@>d�Շ�����[��>��>���!��d�H|�5
���$Rx��z�8}��!P<d���}@<d����z��yE����]�����|_��P�G�G��z"b�c��O��b�'�=wI��HAg�<dY�:C�,�����2��&�9mk���h�Y*�:������B�rp2i�\~�^�}�k��:t\�>Y3�)�8<���7�KՒ˺q��;��K�u��X�`�z>�1D{�rb"��H�a�aP�0��l���`�|�O��Vv�ğ��wÆw��y����_N����� �O�J���>g�&��2t������s	��N~�;`)�XMd��ϗo�~��v�$�z��!����x��Md�~���l$;Cr�qd��䟼���1b"!��y䜺�w��K�`���V�wB�៟O�o�x����l�Y��l��9ՄԆa�5$P���{�#��ܸ��י�ڮ�{ѣ��X��5$�����!��iݟ���X��!����<�Ɍ�!��D��9�h-�߾S�ܝ}��菺�:޶E�t��N��lk�|���'L� xϙ��~C����Du��_>�Z����"==�=����(L���N�/�N����S��<@>N$<a:}0�l�����3�O����~��_~C��Y�N�2`q$P? t��{�$i1�$�7l��|��c?&R����s����믿}��?$8����!�Bx��hv�>CS�!�v��"�@<d��	��ΰ�~@8e��~`}�������3���/�����I
{�Cć�6�c�z�z���C��q�R~d�,��<Iǅ�$��識=�����w:�����z�e���׶yv�R�ĉO�4��ж�B$�D�ke��fғj*t�$A\���Va=GJ� G�֍��r�I-,:�}��˯�wU�C�v���
����b@釉<`xΎ��I�	�'E�`����_]��ڽ��g��u	�!�8�8r�����$��f�;r�z��vC�&R x�G���F�u��S�ߪ��g�=<�́�'�4�Y��<d9�ԇ�?$+���=L�'��bz�/t7�o�����da�����Rc�H���d�[��$4Ma�CԜa+��I�~d���G�[�w��q�d>A@���0O>=�|B�:Bx����s�@�7��	�%@9�MI����y��<�~��_�'�XbIP�����C�OXbx��$�<BT�,���	��|Ɂ��'�Y!�߹�o]������u��r����C�X���1肬'h��a�����'P��2z�RC\������Ձ�!�*���3���Τ���I?��=@4�I��
ot!�gV��a��;I��'<�$���MH����s����ξ���<������P
��t�t��Y!���,��	�䝳��v��0�R�d:BwՒx�P����u߽s�?g}�߾o����XMHa���Ht��NwOC7̑d�o2O�;`~I=a��|�t������?o�s�8.q��tp/;9�[D��U�P`� �Ü'k���2SƏ*�0���\�i�7Vv*\���N�X3+!Q�N͊���]solP��Re���Uɞ��=d>9H�Ϭ:d��SB��ğ�;IXO�䓤��ՠ�'�8���öl�'����޳M�s}�Ht���$�hOR�$�!�?RB���gi8�r�? t�椑~*}��p�<�3q�����}���n�=H�S��MOP�L��v��� V��$���X�@"#DD!�af�X����s�#@|�~`^Y�$��':�B���C�2��	��p�!�"�^go����g���_N�;d�'�Pjl�d'l2z���Y�r�=N�<d�uC���'��H����������=��y�ğy`yl&e�ĕ�ɻd��&��	Ax�v�����;}d�!S2�
}a�����Y�g_��z���'���!��fSC?Qd��{��?$���6�g(N�2z�u9`)�>����߼=���}�읲O_���'�C�E�}Hx����$�Rc�I��'2��v�+ꏏ��0�`��{Ї�Oe��?S����IX�u��'�ԝ ;���v���'l?~��5�x�zɳ��'��P��i���u�������zCO�P��$���t!�;d��a�'��x�z�_u퀲x�=��!���g�'��w������ϳ�nĒ�U�?�yA\h����:���ZF[@�Ƈ�KR�{���V��hJ~���n���`޽�#�/a��ȓ&�e��0�E��D�'����'���!��P�9�4�x��'�hI�Ol'<M뼆�a�'��yN�Dp�XC���z(
Uf�gS}/;���`�����d8��'�x�ndOP��:?XN�ά&�x�~��{�=�#���cg��n3�y�k����a���=~��a�̇l�3��&o�ēsܓ�E�~a��p�z�Wv�}9}�������'ޏ{d��VM����$2wa�5$�Ht��OS�!�o�Ht�,��wl3�߽�:����פ���ɧ���8�̇���$�~O2�Ձ��T�i<d��$������:�<�����E�|ɬ��7��=I����g�'i9Ր�	�V�!Г�R�8����N�O<y���w9�y�~s}$��Y'��N�O�ORk��C�q��	�xϒ��!�!�� Q���Dn���?�G`�ڮq8��B}l��Z�~����{�3�9￺�#�1�]	3^�L�W�2�>>Ѷ����݂���H�~7��<��U9��n�����~ʦ-�	��w�=�����Z]�E��x�X36���B��T�Jg;!��R��zo�e�_�݆��]8m��T]�L���Ck�9��Y�%�~��Iշ̼��g:z����сܝM��s����}�{(�J��*oS�7n�V�w[��fU����'��KXHv��wR�1*�hE�f3�.��m�C^uɨ�;6�r�>I�mh������)`۪R�ƐzN�)���pg���ru��!���[��r��b�7��R���.��r�Ή9�sے;6+n�juMr#n�9S{8njdnH4�u<�.�bru�5�ޜYkX�	�<���9n�\�<���֊2_����y�.�
�TlB�	iW���Z��i
  ��{@,�*5���pؽ�ۣ����;�M�X�u�]���xL��1�/��S9�Jtb��T��f�O�#�V�>}K� 
uc�NL�ܾ}]�\n��x�����.OW�>H^��)���9�vRX�=�7������yjx��5�~��b���#1��K6)�����|ų�$l��ӢڌS�g;Į\��f�uB"�l.�R��,�$��߁���2�;\�f��M������7���u�h+(Pվ�Π+�tyW;�]S�8�SS�9��]x)j��J*9o|��Y��>���E����=l���Q����<��r�;S�Ǟ���2���d`˘i� ��2�*VI���sG���,&9�ۭ�����r�a��
���t'�����dXw�#&1܃��Vݫ�ғS�*�ք·��6��pݨ�$�J��n��n�	N��.vV7\ճ2�F5_����x"�<�$ז�rl�u�;��`�ɋ�����L���q�՚�'M�95���d5m���e�2�d�6H�ڟ"�Hػ��Y�x�)�����2q��]�����As#:�6�
K)lt�{���oPY�?t7�-��:���Pĸ��nl��������V(�uw��r�Wdsz�����:�z廛�h�1ު�f�%���Z��͆b���0��m�<�Y��#wrJyu|���e��rp*^�xwǤP��ݖFv,�OVuǚ�i��ʳ03���4r�*+���+/��Xo)��o��B�fvML��&�ب`Q�&C�f'ras%��1Һ&���6,S��	�(^L,YUv�%!%<U�̲1�1�8��)X�ک�c���B���S��8+(}s����Y�(���')J�m<�x]�0۔ B��xIB<w���M�C�LT�̅ɆVTP2��"�+�G%���1��&)Lj�c��WyX �Jx�Q dY�k)`Qe*yE�M� ���rI�e��*�,a�r�.���Va*��0��q�@�Ѿs@�{6]�F�b�HN��s�P������Vq;�:vuo.��k-:/6����R�Y51g%��J�䳙ʺ�9î�i�f]!y@P�k�F�-1;�����^�����[Q�ٝc M.�ޮwY
��JT��6T:��ǰ��9"�*�ͅ��q�X�� �&�*���Ώ;9|��?��:>��>�P��J#j���[�1-ۂ�T[�g6��bdb0[x�*&Q�2�.�e����+�.�mf�*�]��EQm��-m���M±��W-b�Xe.;�2��30�UZ�Dq�7.DkdJ%\F�2��DDA��5��h�ʹYˑ.\�ʅ��(T�ıTR�PU1ԥ��F�k�R����̵V��0�\Ld�cr�Uc+Qr�V)mUV�QPmS���̪�m�f%AEE�DA[J����q�6�R��j��J����+Z+҆Y�F(V������8��C�[�{�u������t+�{2�ǎU��V�+u`|�nQ����)n�����Һ�N���r^i��K���ƿ��:٪o*�Ѽf;5w����yt�T�+6-���{]Փt�]������\�}L���짚�c���|�j���D�R������Vy�o�b�s[���h��"/oh�3��e���{~�@�[ŝЖ��_^)�aW��6r�K�=�st���Z�����t{��Ǻ=����o�v��ǿg���g�}�'�^M-*{��Fl�E�v`m���/<o+T,�x`�.�6�y=�1[N��*�9��8~�i��K��t��W�n���6ε�(���EȲ�����S�O�F>c�T|��q����s�U��^��K��!���!p�N��T�]�/����G�/��k��7���U�r�)؃�*v��שљ�W����t�ʉ�iV��=���=�9�W�����LWx}
TߟMq�c�E�T��r9ޥ�챉��΄v׵)	.z�1f3�=m r\�5&�j[��{����@��K~���.BL��`��\K㻔1�k��/;�d^�lv�
�oyt��>^�o�xZ�N�=�9Y;�e����^��I�/Z�R}��F��3&u�h.n{�g��ԶCK�Ou&k�ML�ݿ{i\��n��S��I�l̾�rT���0+b:O�!GW!q��b$bH�ȫ���n�)��`��[�J2����$�J�˒����W<sh��'yܗ��G��Oy1��xtpo7���WܻV����'r�c���r�*~ϒ�<�xWHtD��qW�MޏÜղ�a�Hv����4�ZR��y}ۣz����}0��:2�nL3��p�ؙ���cr�_��;�{�p3�K��3�&��>�p=^���f:-��@��{�yb[���N�Vs��hLs�Sv���}�T}P���ϻ�w�f����Ϊ�<ꔛ�Y�'vͨ���~�<���J^�'�;� �ݹs؂�u\�x���<g��Kk^�����<M<Be:�iuw�A�#*a����d(Y=�k��i��ȰM�nOL��ދB�q{�h˹]8����iݾ,�.�kk%�I�8�弿=�z9Us|�G�}/7rkG���'��^���!�	S'����9��=��m�|�M��L���=5)C�>�9ҷ�܎�^emRb��G��5aoO&��a�/&(%��R�gbA>Ը"#��r�n��n���fy)w�o��K���0T[|����;2��ی�R�o<���-�l�a�W��2A�������{Y�Ƚ��O�;7�γ�-��ȫ�M�65��{V�UX:��<�ޘ-O��wuN�:�v:�ִ��(\���ȦՁ�����L7&���UṖzJ�,��1�^���XZ��e�v�}a37M�t�Ԧ$P����䥈��jew\�j�r���
�b�Րd�˛�;���F��,�K��G���m�i��Tq/���}th�����N�^��e�8�s�y9�\7���|��<�zo�ںz��މK��zڠ�,�HS׈�X<ōâ��N��ۓ�-�qOf��u\1��ȵ�*��s�:N[uh?�d�燪u�Xґ6i>��>�3-���؝���/iWVF�}9��-�T_���j�j��yE=��峏!n�Q?	�o�
�3�*��ߢ2�Ą�1?;�?{�1�;(r�l��Q�p�=�����z�XN3�V����p��:2z͡L���;�RTLG�2嫹y���� Z�m:< ��b�uݥY�0FO)v���D}u�Y�}	}��z�R����G���׉��8��"�b�M�byK� �كA��|���YD�Z�_v�5a������^t(Σ�c����G���yQ��̞���8�z��
�Wm{`U��;�� ��;��m��3.�$���.�|l3����A��Jy���U����:��F��<U�0(��WY�퉺��ۚsEC��ժ��9�3
FJ^�1P�<�G�b^(�%�9Cus�����-��7\�H��;�ӽ��͂�7/syխה�c��iG:sʇ|{.�o���.Lml
&�fF�Z��V�S=.�]�zU���SY�:�(N{�u*�N���6�-r�����qgf���Y8��)`9ܷ_G�"=!�)�9��W�:���G�Bs �-��H���pnUř5�������/���1�w���<��bM����7��O>~[ϒh�:���Jd�ߠ��Z�5�U�8�LWrd�^�˻�����Yuځ�ʓ=݇��.��0b�+f�������^_��(��bҼ���x���9x������;���O����,S
���i�ޯ_���z2���T;D��S^�wV>��.\ڣ)�+���7����3t��N<�jm=~�ʛ��W�σZ���Y�Ʋ��M@՟jnΜ���[�r�V�!Vo��H�D����̵��aLG�ƃ���i2�p5	��'i�.�#��@v��J[6_�ݺ�p�:Rt�6�+7&��,}��Vts�NO�����"�ֶ�,_>�Ŏ}1Pr�^��:6�A�̫ƛ�+��F���+�L��q����P�����T7�T#
�o:�x>���ٱ��������W���N��e��I�HHK��g�ΐek)yZr���ɩޫך�ֻme��1_:3����C�ȑWS�q�=�h�A��(��j��Y�CU�-;�������������B��غ�������/���@��ʽzvu��0��J]_6KIr����ϣ��{��A��"/E��D����\̼8fw[�������U�,��hV�JD�4�f�G�z����4[���2E
FG'����e6��?{�s���Ƕe�����9�1�+��_*�2.�u��:rB׼�-�����R�����P٧:�.��ci�Αa�'�F�o�Y3Ͼ�!5@m���':�+���9�T*L�&�S��Ge�[t�Av���4������D���2ϔ�0��ټ|�a�I�t�����zj{2t���,	���a7~x�g�a�q� �7h���b���˕�;Ό�e�=��K�vg���8�O����8���
�<�8.� $�Jݬ�Ϥ��;���D�m۸��KOu��v�NR��vXaFomm��ژs�%:���R�ir�"�ձC9I������KnOx�~�ct� 85�ڡ��yFkvys��y����蹅��<�1���[��1��A_o�ug��u��LttҶȤ6\���Nڗ�/���5���d�Z���a#���������T���5�V�Z��d�q�cZ|��Wę�Y����N=�]�IvW�nW=��]�ʏ�}3������\���o������)�ܚ,V�0ul�����a�ίw1��N������V{��z��]�zG^��y�	������"_��+wF����_��yS	Е�N�L�R�	S�,�piTP�5/3y��@��&�q�]�j��z�����K���m�N�+/8Yؓ��(�(�L��k���޸ӷ˯U��=\,�`�3���%Z��19y+y��vZ+r"�'S݋l+����OvIEbՇ��J9�Bd��j�DHũգ��7�Φ	��mØ�y��q���zR�S0���e�{&��S[��G��� /�w�f�����6mE����r�\�����D�֌��
o*�j���
��Kg�'f�Ew��NޖxV�t�C"���a��N���݂�
�I ՝�v�#	1a��lJk�=�H
j�˶�%�������c.�Ki�7K���umR���q/ue!{�#ڛ1�!��]��r4b���	�6��OF�F<7O{r���ϝ�C�p��@��E>�rث�-6v�����ϲ���ˬ_g%�J]��w��fa��X���4I�e�o�����)˷s"5hS"�aɑ]�Ɋۗ�p�a�Ð��_�I�WtM.:3���4�YXq��ϋJ�f:̧F���&���Zl+�M+.:͜4h��jb���5y�� nSy6�r�hᆮ�I7�����3 {�4ˀ~D�P�)kqZ��G�T�5�	n���6�>���.tz\+���$K%�~1߽Y�OR�tR��$�,Uxi�#*����ɝ	�w�>+�kh>u�G1�\�m�;��t��F�._�,!,d̮Gs�ʕ+c&����{z��93y5�9���I
ɝP��J\�������Wb�F���U+J���0hVU�SXTƥ����UkeV�c��"�e��h�*R�ѥ����*6������W��4�mX�m��b����+F��5���mJ��QD6�r��-������2�+E�*	n���șw0rT�\0Q�lu�`�5ɖ�ij��V��W.GY�ptk-jj\�̸�ee+Z���km��򒉖ݸ���E0e�m��q�v��7*�w*a[Jє��.%�
�[&Rڍ���L�VQ�1� 0f  ���=��x�U�Nj�<�kT�aO2:�Y6�Ky{�f���Gr®,H˒z����4c����#V߆Ø�0�`.}���R0ī[�1c��[�[�_�
R>�F;	�]8lr�����x��TmQ<cL%��8{<�t�~�����`S��U�n�.�-Lm��Z�����ڂL;���ǲMpR��H羆o����p�@��!�w��U�K�OT�O7�zy���vl�䑭�D��q�[��
}5�N����[1?��bVM�iRb�QՇ3��g��Irj���p���
OWO�\�J��]�j�>��}��:��JG�C��zm�{�kL�|��'�s4qf����t�^���f	{+q�ͲL�W�i+�ُ[�1،�r�Urt�7�MC�F�;F� X��<4��	�����wW;�]	���?=�z#�݉�YZ��>���l��㻷��O;׳Mm�H����G��GM��p���o�?W�ڧ�(����z�ȭ�dpeZ��f��L��Mf¯Tr�\��<N��	Hs��r�g�z��Vp�mOk��E��؜�c�^�"�t��5��k@��A݄�r4I�¥zyeJ!��\]��Y�B�B[�����=ڄ��=�;/��^rIM�э���Qj�z�/aIL�������&{�7.5��k�1g*��k�X�X�񻠻#�]���r���� �Sb�����I�-ӻa6�f��\��-4���}U����s�ݢ����Ü�N�J[;�fY�(��=%$}L��&|�U�"��6w�����p�^�.�_v8/��ؑ���n\);9��4��n_=�=��>�M�.��<޽���#����Y�z�+(�����ʗ콓Xz���1v��Z�8JkWf��ihkv�׫ױ<m��C��xS��4���N:�eV�]���E��ژ�ZK$ u2������U���>�A�)�_H�mת"��Xr�y���ہ����O�n��Gq^�~T��%Y	P2�3���g�b��&P��ޡ�.�d�p�k�]$�wL��Sr�J�Ǳ��(�L�R�N\)%�r��R�ַ}x�}��GB�2]<j�;����x��w��my�`9�+��y��U�o����9׋{�n�oO	�q��9�9�񏍋�cj��y3��&��Q��O�ө�к��Y-w������y���J'����'�N^V�Y{�s�����m-�������:")^����L,d��#/�ɃZl*´I�쏺��g�M�ux���U4�N��"��C�%��)��«ݔ��5�=1��L�3Tt�u4����)yV���G��R���I�q��P���p&�F{o���m:qe�=�$�4�$6t����x.�z9F�V�u�s�XB����s2��-�-LvR��S�[KVr��z"#�Ս�m�m}�bsoGkU��R��Э3�/�=ޮ$�sY��#K-?O
�ͤc������޴�{����0��������I9ڽCݕ�r����u���[J�z�������>�У���O��GJ��7˲�;z��<߻�<����vF�ϩZ��jy@�����#	��T^��kv�9�r��7y+�V��_�v
�>��F�R��-/syȇ^��r���Y��Ltz��;:7ꉥ�VӦ��gh�%�\����j��b�Y����WJ3��,�m���Ek�1rP�؋N�|g]3W$�벖[��$� �2jOf�>�4�@�>����)v��V� &�R�ʐ�G-֛����k�50���_TG���Su��c����������b!������K(x朕��+R��K�OmcK�!��u��^��դ_�G�p�ҕ;�׻����sM���K̨����=��\�;�h�X����Ag�aB�h���L`� ����="omlv�;�ӯW����U�]�V#��Ŏ
�p�fN�S����i����6K�0b��Us�x�"Q��2�z8�H����C��D��e� �Pc`p�����2c���������0�劕mg"U�g**��HxhN�
���֏��z�ztE�p���e��Di�&h�1�c��Tb��n1�
�@[���4mv��]������� ��YwtX��էrl���˕���kV��\�ޏG�=�ҞN�8q�3 }�@Ti�H�<#���XH�S�#�Ʀ&s���<v���#ћs���,�5�`vE�=ۭڡL<��*�1��uM"�L>��zXU5E�����0��a��b,M\�P<�5;�~<�b��&3t��jo��"D�&(�1��Q��	��s�k۔�a�)V9�;j��E��x��D`#4ʉV ,Or���p�4w��	��ŏ�0�Kr�B:�Ab�c�F�c2z�A�b�oO����m6{Mt:+:�{���V�U�F	D������^�zp��C%e���JKz)N� ��|C��y�����~1�"�x�WkZ<A�X4:�]��]2�8s.�[�pT��a["D��Ķ����sy5�g<G��+:�k��r5fΧ�Y�9mn��S'ζ�r�38��#�o6oB��tǎ�:؜)�?}���n�>��ٱ����C��g��13��65���>*��;�d )�|+MiU�
F�Ҵ�~\qj!
�ȣ9YJ���Nc"�u���du��s�
TZ)x֌���v��ھ]4	c�X����gO�&6��ĳ���^�L����uy��`�ϵP゘�Pђ��a�S��#Z9V�&̪/�X��b �4#��g��DҞ!	�P��v�=r5������#�C"�a�c�2a$=3KN_m0Afg6�{�`���`��bWDNp��+���
��ej�;2e�r��ΊX|0`���j(**��򪘀BW�������4�&F3�78=,���A_*Ū��@*w/�wb4|�q1���˳��R�j�[�9{x`E�.���G��pY�'q�up�Ý������Ȧ)ֱ�<Y}��3w�M+rE�j���������F:�gJ�x!)�3O#���D_��b�n�,Ñ�;�`�WJ��o(4o����o���+Ul��F�:�����b��у��&�gg��&F�:�X3N���{5:�2*�w&�Xu�Q�N $�����3B$��\x-����A]s�
�\�#�~� �nV�8N(^��재1�A��au���U�Մ+�F�5V*�X��3�����gR�*r�0�{�Ő}����	�<:�dz(dJ�Q�2��������1hyʠm9�'c� 6�����;Y�sV&�R�{NJM9���g�j(P��)�:G�8T���|ڡB��ɉ�c�FEٱ�m�)逕��%׸%��''�v���^�Y[��#ѕ{R�������. �٫��+лp��.�r:':ojnVI��
}�r�D��w���!zDɷ�e$�"=��`Tbҟ���j��C�G�gm*0��ৣ�\-�x�3=��8$p�
NQ�b��A�10M��D�: �B.�<��z�1��|��Ư�C���M���˱sɋ͈a@"+��d����"������W�29���x��3� ��t��w=l�No�4t��F�Ý���;oӒ%�9�W{2��@V��W���ϴV�����:M��21W� �р0q8��̱B,E�F�E[X�nx箶ջdP�L�����HV3,���Ra��Mg#9"�LZ0B�a�X9��G2���:;�;m��w7=ڊ�5�����������>ѠU]^^��:��+&X�:}�&*�/%��H��S|ؗ�գضf���5a���C"5���J �ĔpH�;��]z�#����ҕ����a(v��Q��>��;&X��w�Q3���/٣kU*�xK��Tl^ zF�Ga+әF�Xk����7v�q�}����=��,�b��w-����"�b�fj���3"��[��沕	ז&�@$F�^��2+Tܰ#Ϸ{i�)1C/�r��g�*��F��!d��w왓��γG%l_c���ޣSx��� ����̎��KB���N��S$��"�vgJ�g��T�JWN+���ĕ��ov�u�ޅ�5U�X���U�����z��Å�*d�0_MU��,����u&�i�m�Q
��]����m�jz�W�:"�+�oH�w�)X�r�J[R4�v�T�f�4Q�.�5��oeӼ5�]��5Qo=h:IT��i�b`q�|^�I3rB/z]Ŵ��˕�R��x�y��oTXU5݅��v�YM���JwFPB�mѹS
�r�V�lS��{B冐�z���7���QwW��9���u�ݽ�Dkw�T3GY�.}�뺒 r.mYZ�p�t9��7yt����h�#>G�
�jG���E�^x%��|�a�ز�>!��}��������\W
 �˂�Q�b\��r+��J�O��ܨ�c�Ce�/m��(i�K����|�;(R��Gk�+�`��:���Ay+*S��f�"���H�m����a�j-� Ttn��+v�)�����}�x��f��QJ+�1][>ض-AaC+cc��y���K���c9�ڰ�*T�RfM�!Nn	�)�I"�Xs��!R�1a0[�����.�R����*H��x��G��@����1r��☶�p*�"R�m).�r�
�eYeb�F��a�F`�����Š�b�������ŊcDp��Lj�V-�mZ%�Qmb�[L����R�L[�0ƩU����9�0��j+-��X�[F����m)JX�m�3JZ��"�Z%�Z�4J�ܙ6�K�V���Ƞ���-��S1��0�Qkk\W2ڜwjm����LF�Gp��R��i��TJ����h��mj��ʴ�ֈ���+TK�+�x�w
a�@�Nk������9٬���Pf���*K�w���^vZ���[���Dz"�Y���O��5�9QQ&è��,�"[��%��-�#�73<����J��j�A�����0E��	j`Ld�H1ß�%��sxY�oI�&*�Լ�eg�+r��T&�46P^� t�U��kv�}: ��p�rj��!��)���3Z�g�35{�,ן&����L�@��} o\������PB&��%�]�ͻ��Έ�L��l�#x��r��<��:��Ӓ�`ɗ��6M�]����ҭ�����O��+8�=���+��-j+i�)(�bޭ<.A���:�k|Z͞�҃)9پ�JϤT� QlӢl.X�h�g@}�pn<��X�\�v��CG%baP�0�X��a��Z'�[G�\wz �ye���1��ɂq˒���7�Meoub��*�����7���N�}��"X�Im\=3i�"'9�F���Q�{�W`�v#�E�ꪯ���;óOh�nE��>1<ph�PC�d�Z����ئ��^�/;�u���nXw��,ل���T��:'��K���JǏ�_ap�7����z4�emp��1�c���´�b�.�y���V�ꁪ9���g��h��z�p@��S�Θs��Ԥ�Q� �409k���~E�f�x���N9%��a��!
�R�A1�l@�Q���p�E��,iv�ԭ��Apc�`����:8�WC��ĳ��#AE���]N���v��ȓ�2��1Q�x}\phu�Հ�'��˼�t�=�Ο-�hx�t�k(�� `���#���<穅�\����4�
�"hЎgݚfS�!<f:98����G;TS�YS�dK+d�V�5�zw�Q�Le޴OR�O�B��>���L����juk]y��p"�t��ٷ"���b�B�SBe.Y���=�*��su�Ԥ�U�!
�Cb�`,�;`�pzd�s�:�ܺ�p}��,g��$8G�$Eɛ0g�Bnl�������S��P����|�U���舡X*���5`�#N�m�X	���M�K8&�+��O�D��.��X��XW���J�����\��3K��`�*D��5S��e�$�Ӄ_�c��1n|���w�o�'GnFLe̭�m�J�W��@Ma5cyd>��-}	�m��$��I�p��Pxd[0��l �.��#�"���V��7�Hg�+D�Wa�>���Z.O
�P��a�p���\�e�"�b0��ܥ��WF�L��)!��w�\�É��3��Ɓyz���t}.MR�Ԍځf�l,ݥ���#z�e�η�z�&�:vs�@�Q[0]���.��.�Y���J]��}�z=�z޷u�z����Z�i�(��r��PІ�T��z�^��]�j�ŊUY��'��0��������f �s
��Âu�.*���Cz�S���R��[f�����0Y�m
����ՋS8�8.:2���T���dL8`ѓʻ�ݹ�D�-���p�%�� )n�a���8�e
��fqUg2f�|.,�:��`�[͇C�md;u�Qn:!m�Dw����NR��E�����g��|S����
|j�P�����貏%=��h���E���X�gj#f��X5�a#�
����k�%Sa�M
�X�Q�bb�ƛ��9B0t��xc����Ec�??$j�����{pr����	Ôy����"��X�-Fb�u�x#�GEZk6�lnt�=x�5��C��99�̻;)��m×.�Xr��WRQŝ��$�;re,-�K���=V7��5��s��`Oi�O�:&%N�e���61E����3����=���`��p�P* ���N��7��]��P�jU2V�cÄ����TZ)a�0@vR���U=��*��G�Sf������0G�9Ap��x����v�u�Ǣ��LW(!�$�E	ґ�>W6?b��ܼ���aP���(�A�;�
4`^Lp��f�ֶr~�<7���������*.�W��tP\�ء]u-c�`ZrĢ�J��֚�w�� 4j5LLQ�1�fp��;k;�s�E]�yv�������k�D+`xzӰwCo��
̋�Y<zj�Չ7��۞.�Gj
˨w�G5��n��-7+�5�q�����_��Mmq�BV����1������Բ���|����䠤*�
t��3���D��<�|���}UQEb{Ƀ8>%��X�#<�c�E�ؗ>�kL�4���;5K���檤E�34�c�z�p�b������PW1�p�h��7ʧ3OK�
@�-��W65�A����cZ�o�Ǥ�ߔ��cF
w��(�f�*R��Sp1�'��t��0cN�P�Gnm
V,]s�o>�EğN���i���V�"���u����P냂eL!1ǆ�Xc6f��]8�gc� ��U'8�1YQ��&�p�;F��
WVԖ�hu��N��:%g�B�B���\{�'¯-ǜ~_.�Pz�����!���!C�&�W�k0E�;ɘ=��!|��>G�!Rcf8�n��$�<td[�f�rZ�ʼS��]�"���xy���ΧZ�K�Y�@=>Czj����4���uj]����0��<2���Vi\���M��t�����oR�Ze�e��'��i�0�
��La&:�gY"7�s��CK��8P���1Q�x}�G��N��\aeWu���*/���\��P窇��V4 �GFiL�IoVǧ�g�I����PɊ�|tZ���B�T���jxVP�@GK���N��P8r$1f`�b�и��xP�Ʉ��}4F0���C�\06o�$��&,��
��GN��_�d��������i��q�^הO�E���W�)3[�����w U�7���NO��,��%A��1�9�,̫��1y#=38C�8=�#%N��<)=�(e�/��Z�}rvn�-�&��V��*oí��t��W�1�=W�7Ǎ�@�wxii�䓼}�B�o��F]J�7a#��[�-�ԩW,pF�����R�=�o\|¥=�v9[��"�due�ە.ΫF*&�[&5?}U��1���݌���:plY84T9��*cG���^��Vn��O�0��Uz��������6 G�\�Pzl\`̾��W:t'1!}�@��GU�{�~�}h����WQ�(��Δ0s�<X���PSh��kj�B���˗�F������c��c�jP��<8�!ݛ�Ԏ�i!��l��0��;�.���aC1��ƹۥ��t�W�� 	J

T>fւ=T���D^�(�U6�+�a��5�A���������W2:�&�0|g�����#�q���F�� BE�6�0�D�xX#תb�k�n�P�7����uz-�0n�%i�F���<Հ���Q3�d��4���zp�=Q�rf���3��h���d���e�����3\t]g�N��b�F&v�)oo��QoѾ���BDܓ��_U[*=�H������V�f�#�Msr�F�e�>�����RT�*�ǅh�>7�0��ڬK�Z�F���`"�� c=�bi�m\��9��b�B�Y�y�>gm��F�̙�4���`<@c�l��<^f��y�/HC��"p�U�� k5(�
����E�{a�O{3.큂�6aLUք�F�7�ba��j
�an�x<�6L�\n���8��*�5�8N�áZ6>�W+�=���U���U��|�R#H�y�q�LƎ1P\|�w��p��S1��g�"�:�t����*�<qX.j��&h���'F��Fɂ(h�����4`r����`"��3]q67�P�L���e���YV�A0`[�N��#�1Zy3���\+�y��(��<�z�8���?�������,o������
w����3����ʘ3YQ0!�'$gQY�S��P|tpb:���MT4F��&hףT����|�]��&L��36@S0] h�&k\Z)}�X�::zg~�;܀�J��C�Y�cnA"F��h�����j�ok7�$8�<+���(FT�K��}t�ײ��WJ���Z=�y��+xg�X��SlJ���\+��!��u�R�rf�c\X���cH1%�L��`sUc�ր
3�w6fwH�/9A���G	�1s4<�7M�5ӗr<8[z���h��Â�����Ф���4�V�sC]r�f(<��7,Fk�GA�b,ڊ�X��N
�0�g��[mJ����FfP�0ws�M,��ng�;���!��.iU��:��:�/����9.,�:�kbf�^e�X���V�E�f�pٗ�R:H�25dd�+]��T�u�G�)GM��ɥ��]s����4�eY��0�u�3h_Nm<�i�g��3
�o\�h�5y��V%3�/��k)�Vc[��WeF.�E�C�ˤ �sM��:- \ծCn*V1Ar�J��PӉ�J�p`+ͼfi�m�z��(&�+E44��;��U�%�����
U�؝�3���w!�ՆslG-�t���Ү�_b�yQ����,J�D�%n�RG(0qA f��o���d�_*ר*�|[�2�etZ��L�L��<�{SC1�.�����Fzִ76YÛ�ܣ���iQڳ��U��)���+lD1	9�`M�WZ���';^6��n�zA�RT���zV�����u֧s4��{�fб�U�qȦ8yZ�.|Ĺ�)k�k	��sj�wRu�86��כ�l���� �r�ں�����	g]�ᓸĮ���NY��ц�r�̴3%^s�{/����ov��ų��*9����4uk�OkM�xQ�X���M�ղ�X�p�__��P� �7wյ'I�zR۽�F�M�G��t�A�����v����X���Ը�X�1s5.�]�%G���U��h�ߎ��wU�9{�����"��.Ë�F�t0$^z�a��q�6)o.����2��4u-�KF�f��*UؾV��K�=]��ӧO�9<j��DA�vɻ-����u�b�o	�[1N,��[�^�"��{��X��/�m�D���7����Z��:��]7����c�)�n��곤��;��Ƭ��n�G�{M��]����5y���%ީ3&�d�����I�����@ǳ�����ǣ"���:�����ȑD|@�X�[�mTM��naV��	Pv���+m�1�(3-­[�]n��F����e�E�0Ȳ�YV�*�G)\Lc���m�eC��ME�c���n�妥2�a�j���W�3[S�,�2�4�\1��R�-�䲖���2VQPI&��J(2��H � ��ݻj�KKD��cm*.�%�2R�L�n[̸�F����m�Yf4q-��W��vk�S0�7p���9�F����.5��&�]˻h㘱�U��r��:�F������TB�5̮��*�Q�\#��-�m-J��(!"��D���w�?7��>�su��ΦqY�o6��n��|]R�M��Il^F_g,��_DDB-�&�͏�	�e���9:�,���+�Z)�SDG�>�&V��m������ DR��C(�B%�F
O�D��p��=L��c��fq8�ѓ҅�b$v��(X�e�z��P���Ef�Y��R6�UӢ�Be'c:����-gtУ�%YC�F8o"�U�֫g�g��Z��m·z�����vc�@�<!�V�6���g��n�f"������u����`͆M��E9��t���� lhX[>�82��(��2&͈Cݑ�`�"b�ZC��z.V-B���Ŗ$\�2L17�b��%��a��:�\��������.���&0����6"��C�ٝ��B��fY���D�_`��J��;jU=3��eq���pXáue��+5 -�f���\�t
��"\OoyӮV���*c�W�E˗��%J�v��k=\!��>Y^�)g��<X��mh�P���<��jv��9��݈����py�����xP�j�ϱ&��޿�H��W\u�#�Zr��Y��p�0 ջI.J�C�84�Y1�+���>sQg�3�3�+FP"����i�W�LT��u@ɱ��T�����d>��/�����vKŬe���ȡ��0�:`�� ҅��B�͈TF�rs5�Uq!����yVF�7U!�(�[����.ö�W9�����zoO��"���ï���p��14��'�>�FpԸ5(u���T�^��j`���@��;7K;�=9�f�ʩ���nb�E� [0�����o�F�x�ZSUʸZ���=vu�8�=��aM�^^��(!t�B�oP��n[ �}�E��VP�����
�̱��w-�w3S�e<!(��V��}yL�����#s���⳧9r���Bw���B���.A
�>f,'�t���E]i�Q\��`t�Z�Ɇ�g�3�E"�@жf*�@g�ё�N�� ;6�9��#9��
N����@M�!VX؉>�bum�1��w;�
�$1�t:����$l��S�A�1c�6)Gbƛ�>��J�^��A�KLm�]w("��sA�׊�m;�kpFQ�n&bf:ck�
h���6�ph�i���l������/�O���D��MLM9����1XL؍�bWq��pm�$��U��V�J��1���X4��
��-C�?t61��J������
��{�A����g�O\��)՚�����k1@*�B��=���c6�VLm̤=�.�����]�ޫ��@al�=�����C�����W�gI�ģm��ꪓ+u�u=g�ݘ�(��X�b�f7nXCAhݨ�V&�m��7�u'3܆q�p� S�P�3ΝYvN��h�ZTF�֬cE3�0{*p�4zbj�Y,l�J1z8b�ʹг�"0�3£N�'Ar`�6� 1�%\WRZ�70�`�	���l�L�`�NT8v2���/o���b������[!���*�����0�ʍо����Fg(�д����}�����f�)HS�Ԛ`�s<'�b��p�'Cƫe��8f-��^�;��H�68�2]F�":5�R1��΂㉹z�
�����lE<�,`Dؑ��#��4(�7y�#V��$�p�[3���n]�q�$ŇW	Y;@%(�V-7� rv.{%J�ɡ���+Z���.��{i�bTF�ۥ��;�-O�#����23�>�q�c�O��٭�E��R(*�X�Xq�P�[���p �9�8䱱��P4$P��#D�d�.��$���Ն�<�8Z,M>x`�c��8g�`�v3SA'�Y�͡�"::�u��G9�n2� ��'�"í���O�i����a�<b[q�S��DV�ep�S�kٻz�6��R(h��:x����Xȉ5f�OEc�[2��n�^=��cQ���U
a�P�� j64g˗��� �w�R�9����\"�q2����b8��tF�	F�B���Κ���N.F�!@�@��{�%#S3���asKxn��+�=5� K��@W��tu�}���Z<r��Ƿ��pz�Q60P[���`��n��{p�h1XJ�řݐ��m��v��t��΁ a���;&IW�o�.��@iی����ܗ��z!kW7jč�6 �Vp��Ν1q�4��g��� �!�U�w���'��W�4��@�t^�P![<��jn��Qu�G��>�d��1\T	8EYD�T��I���{U�/w;��l&�Ŏ�0�R9��|�.�1E��y��W_�7^+=wƄ\a�t笡p���sa�첆{˚��M42B�b	��"���q�GT%_X��5ep�=�.�RZ�;5ξQc��ɉ���8y[ZM{
�θ �ca�2'�WU��^LU��p"PtcGR���0�Lwf�8�a��74m��_s�V�Y�M�q@���RcG3�^*��`�³�g�-)bn�ӭ;��}�SUs�X6 Gi�/�Jr?-�=*v���yd���!:Y�[�![M����T�.1��h�e�#~
��Zm��#⧺�o���&�˛w�Õe��:�$��凘���f[�����wf�p���x��U���\T�й"�������*�T��LF�>�(p�9(t�2%���P����-r����,��a�_s�Č ����#�"��ky�.m��L�N�TY�|a��!���!#5����ΑD�b"����T��2�K1�C3�8��o.y�o��08<2��}g'�f-T�ג��G]�Z�����(O����Bi���%N8Q�^\-�pn��L���b�PAҐ��e@���@R��T#�X#�F��4F�	���记��P�u"����Rj�B��}��l#9�V����/�3S>������ GJţ��:��;�˪k��ȷ�>4�'�8G2�H���\2�A[������whY�U�ݽ�A�4j���jK�a�^��'i{P&�m�ХK��Mw.��ܾ�G���|�7H}jbӛ�hM\Тt ʞ�tܨ!����|Cˤ�a���xK;��kqU���FD�hC�S��Z�,���B��YhƋ�[)�9��ڨ��xDtPX�j��ޞ�^���n�
'�](Ѥ%�8ti�����:��H��i̙��Q��X�b�z������T0�E#��7m����*&�X�ZL�)"l���*� �C������-ptp�
� ��
ш��ʕ:0l9�#W�4��Q�P�x���Ng3̻��%̡Q����x�3��.Bk�;k �����k�
����Z�,���K�������޶��|����Ȟ )�c�"c���	MT;R+�6;��JW���x�*�V��0�'$��r[�ckH��oy%Ay��o@yS�;h;���}�^��\�Z�<�=�an�^K0��-����
~�wO��=uܾ:%{ì_0����3� ^��\��%���8+�壢S�
q��S�K���~�o-�)�"'/6��`vHz� l��rb༨�~s���̉8��L(i�i��¯9B/�8zg�Q���X��v\��t͉��'�J�,�k�jYyQ4pD�Ń$ە�m�
�ǋ'/oN����)d�\>������tXW�ۺW��2�;��������z�A+�BӃC�僆�4���od�gx������+�"��H!�ml��G:���o�ۤ�|��c����@f�;���mGI�s�b��+��ns�4.(?3�v�ĉ��+�`�N�@���@�,"ݾ��/�ShR�q��ޥ[�_iB��PV��[A��e�Gwj ��b��SYכJÝen��9�ۊ^�G:�eoU�V͞V1%�R���y'v�3z7O��aKL�G!��d�pp(�Z �nZ񺽶�(����2luD��4V�*�J�x��_+G�w��*4�_$�+�!�l�VF+
�s1�B�TJ��I�-��5�u�&,-�D��t`��!��;�aT�@�٠r��[ٽ���EN $^}��.X�B�0�|�P�65��]�� (pp*]D!b�q���5dq�p�١Qf�t�P���2���0�����`��D!NiW��bF�����Sk�73c����OܱaS���T:/��U�`ҕ�^�Qy��L��A�<)T��ab��h�u���/�Ϫ�<���917��d�:B3�-xlգ�r�V�U��b���F҇�6s*�h^���+͚�R���EVasKN;���	�n]U����`	��:9C�P�n�ڙ�Z�4�mNA�%����~�n�`��Σ걩�!��e��W�]�Yt�3���̔ѓ+�n�jٗ�"�J��2���v2~��Il ���noNef�~�w���J��}ɧ�$�4P��U}]պ3M&�Su�h�e�� ���*����yݪ�?i��"y��,�J�ΤoO:ͦ���%C�Pm��+*�g3S��RV#Ys�Q�h����U�JsN�������y% ��*Q�H�������NSa�*$�yո)U�˼P����*lڔFw�����jY׺v�Tǩ�vp�w��o�x�ehR��r.����3��}.�Z�*ğ�P�����K��p���ݤ�%4��E�3	���ٍ��̨���s�[C%�]S�|H�yF�MPm "O:��[Ԯ�=�3b�aVd�<7B�.X7S#̢�_e5Q�je㻒�Y_d��Xm��1�!���X�B��G*�w�v-�g)����ʼ�_)1���X�\r��V*1�#2�-�*4*��&ʹ���Ze٬�|�Ŋ!�2[�ű��#I�)��2�*�j�Z^bv	B�:��F�d��Ô��)ieZ��9rؠ-�J�ĭ��M+�h�8��h�y�9h��7[I�ER���C
v�P��Ŕ��BA�)��E�v�;�t�1�Hd��J�]�yՎ�x�[ͫ��5͢����퀳��#�:ȴ2�f!v;�b�7.�kh����[6�Z*
�b����w��p�r�:i��j��k6�MHg^[��'7X��Zn�7*VNŒ*���3�����fI��9��9q`y�����n	;GR5�|���]��V\�2���al�8��r�dŪQmZTq�mܦ\TS%��V�.�V*�ۮ�Tq��b�u-
�F뙙Ef�Ph�aq)Ej��1j�iSL,q�zҏ-\��Uf`���
m��U��6��`q�q1ƨ���J�L̘�G+���h�g3c�p���n%+k��1�]�L�E˅j�4�53Z����ɔ���;�&�*�0���+�u��5t�Ԭ����.%��)nfa�*.nb�0�ۂŋ+SS0��u�[�1�f\0M�M�����Q�u��̫��*"���F��74�X�̙��F�L��(�8[��0�yIE���M��U���C����fhf+͝9�nfuC����e;�w
���j�cZ��J��ݥ�T՛�>�Ѣ"�I\���_�{ޕ+��b�O9��"�Ϥ(����BS�5��TO`l��rD]��)s���[2����1J&'��<:�îJ}� 9(�x6X�P鉶�>�Ɍ��c	�'f�gG�<&Lh��
�FT�4̈���iy�ӜxG���`�p 0�!�^_<o����Z��%VN^(���B��|b����.���mܲ@�''C҃��a�L1:dAE%�6�;�F���mt5��Pt�i��$�N��ӹU�tT�\����ڠQ�צdh���'d�s��)�̷0���/6�n�\�mÎS�� ��������k��5kA	�K���]~�R�X�[� ��w&'T�:G%3�i��h��IS�����>ܻT@���4*�*k��1���6��n����Ƽ�r�/�S�k��؟<.��t�P��W����_{��od�ڌyS!ёZl!�x�|`W���[s��0���ʞ�w�����(ų#EEܰ��Aޟp�;G��_t[U����y�q�T�o<�4�)�����V[��7�r�N��4������n��l�a��2��������/�o�8�?^�`����Λ�G�sB�ЅCS�َ�*�,���^�P՟;��a��Ȫ(��I�ei`����{=A�k~�{�$������.�g�,f��1�x��0 ��ϑ�L���凳:*rXV��*��dZ3�
����F�/�R�w���U� l�J�G������<i��Bb�R�li�M��I-��R�����t]�c��OJ!Y:~ʳ��y�F=ᛲ�i6�8,+���,Q���=�@�k��Ť쟶Ôqol�R�E98ܣ��	��ru]]{�{s��S���D�T���d�e��α=l<�z��pZc��t�`G����c��Y���]��u&_@���S(T"�wSK�C��:���8l�J��c�n�z p�8D�tᢶ���-ku��&ǂ�1،s7}��V41�B�EZ@���3m�,�L&�]�V�6v���1�l��4��*Lׇ�(�X��V��@-��*ٰ��'ʬqN��ܝ
�m�F.��=T�K,ya �u=srn��þAŞ*9�N3�������2�w������\�((�0��	M�����Q��U�t��Y��-;��p�n���6,t!j�\�s���,I�: ��))�8�y��f5���k�u���|��`�/�^�&z�Q�>O��:#�ܱ�y3O���	b��nqL��ٛ�t����J=���Z٭�v#�<RC��������)����r����}��z���UU�򑘱���F�>� h���X���ᣄ���|`.m\e
�U[�ϭ��p=�$�eN���7�PzX�y:8f׹�s�{��Q�O ox���6\���@]�/*{^k��!G9��#���HK:.���Xv�1�����{�5�Z�b\L��o��HH!3�8DG������K{h<b_\�g�P*D�z�j�Ҷ"N�^��G!ސ�n�;��!�`���Tǆ#õ��LJ^��u�P�5��,:���z)�օP�W�]^P��(L��e��	���'�J]�v�Bv*pTB���|V:b���q77����|-À�9�8*1�t��P��T
���[w�ԕ+(�P���Ky�`u��&�ݪ�5��$�zkq�<�ܫ5u�i��oU�ԬO����S�8_JV����w�{R$�ِ�a��$[�H�s��8���x4F}O�#0n�3�5
�D��NiW��Pp�'U���}9��V����q��-��p+s9(��>�38��j���񨏲*d�d<*Y�7TcE\b�
.x9�n˽��j��Y6(**������]j��lTケ�r�3cjx��\)x;��sn��t�P�F\V֓Q�W�!uM�淅�/��L��2c��(1
��$.��n��������]N8敖�����ڠ,,J&��Z����&wtt����\8$�:ѼxmaA}5W:Ղ|N 3�����F��i�u�{i��IT�ʢ���Q����ʚ����fM;[�����tU)boe�.4�-r�=^
�`B��ì�b��x�Y��=��6�;@�,U��3��7������bΤ���hOp���F�r�5C:�3{ʏ�bt{5^j�3*Mu.Y��}�yx�Nw�ь��k8���d�9����ET�*�f���BS�ϑI�fF����=�8&W�(G����^�>��־�b�0F9��b�`LA	��*6�����N*2���m>�G[�@!����B=Y(�vW6LM�w�����i�2�.hTY������r�G԰t�n��c��5˟!s��>��M��YCg���ƀ��f��<�܆_����ym��٣長�'@_�[M.�O΁���X��*P���W���z��lQ�ڱ��<*��.�ʱu� ډ�ť�Z�k�4۾�j�z���,*q0�������ZD�w�/-K�/�6x��)B�j�ҟ�o�UKqU���(cK��ս�h��fL�4z��:�䮜nu#G됓P&c97
�]����V:[��	�{X�*���̅%2��.=�J՝��+l�I��8�ꪪ�C�yU��uP��:�'��p�-�P���H�qXc�N��a����������M.���� �|�!�u��S8m�h>��K��J1b � 4wf`#,�Q],Vk��(m��h.'^w6l��LhtX��N������^*ЦOJ��-j��Աu�\mUp�BE�����q���t���*>�7�f�RTI��zu�T�˓s�B��D�".zc������E�ϟ
�X6���:�F�Q5����%J�����	g������EE��=(�����c
#�xV���R3�r�`v��ޒe?V���.Y�F8HB�� v�{& |@Uݒ�ٚ���8�+�#l�i�xE*t�Tt�m�<��{��1�������A�O�Q���x��a��vt���\M�"��Y)_���q����"�;́K����(��j�]���q{Vd6r�I}舎u�`�CF�ϲ��!Y"���ŢÍR���M�G]8]��k��^4�P�iVr�3mh��b�����N	��bpbSN�޺�	�����3�5��:�k_�
vo"�B�(�puӰ�=�M����F�(7��������CBF���+E�n/u�f�5�X�>��'�9hw��3N�F��0�
����Z([1cA8���1&c�i1��5jPw��q�\�z�Ŝ���{k��N
�0��:8 ���u��m�S�z�S�:�b��<Lf9�� ���`����\cx�K�AZ�U�v�E��lL�c4�X��4�h�s��(EV�4�S�kCh��������L:GEhhRv)cZ��x����Q�����%,��ݫXZn�ӈؕ�t�б��Zڹ�W$[�)1��V���;�������<zmCz�����bX�»�������ܗ����������rp���p��20�0-���!Q�	�U���/�[���9eN,(��Y>K�f��EOС��k���z�J׾���
�YMXC*�>�w�e��!k���K�Y}�2�h� =�|5�GC\/Ni1b����tv�3���^C!i�`0\%\O��9�tw �:J�(P�)WS�f��:%^�{{���˞	���q��-��S����Gd��.�y��y���cY�tPwi�]W�D�Pu�ž��|��@�j}O%��"��(E���e�wκw��s�5�wNv����Kn� �Ƙ<8OdШ'�4b���&�0�i��|���hM^�9�Z0O9X�:��>�W��]���n��%�W13�:�f����a�X.�C����x�wb�s4��A@�H;�8�VmǆJ��6�����Z罧H��\�/��{�W'ΨT�8u)�zb�����U��v� ��Q60�Q�7-]�oX���S���E�	�U9f��#�w�B5�]߂�it�DŅjP�>��xGo{)�.m;*8�8K%
�(LE��D�؉S�X�Bt�k9>H�B���P+8���2|<�N�����j���k�ͺ+1�����đ���l��.�� iE�+Ƣ"�j�^�y�g�4ܘ�X���=(l	�ՙ<-;�w�/{qJ�,w��h�NT�v��ǉ����+��V��m�7��r9
�"�M
�a��T�\��ڛ�@\p�ѱ�]a.޶�c�>�bj �Bc�E�lwp�ҝ�oV�S�W���!�C�;��6Z���5�S��8��EQ�pr�w�-Sꬃ.��nۭ��'�ؠձL��۽V�x��WV�f�9.�3h\���t�;�P��ǬQ÷��p�ݺ�U[͘��2�AX�l9����r6\�v�޺�-g1�H�U�+mSb��M�d�!���9OH:ɳ�K�Fw)�}s���ǌk�z��WbK�
�7y�o~�֬_T��կ��w���䱻C�D5�]kM�/4�|.�{W�5�Eg]#r�Xp/%���2�dFe�t�#�h�F�SI�ͻ�s&LLu3��-�m�B[��<|�Tn�mvnx� ;�o3��F���cv��τ�Q����՛��:��yr��-�A=�T��Hh[RQ����͍�e�,�b���r��8M�(�V���u�s-�:�-�����ɺ��Z2�v��y��,Z��uM�o�ռ�v�6��ɉ�V��]�sw�,�q�n��&��_X�Ax�,
�.<30�Pf_�1L
6e�fB�(�F}d�i�#f��yW��
��A<�������43�@�-1*1R&��h�E�,�9r�ˣB�]�2FV���_~�ۋ"d�<�31VJf*.œ�t�/mX�r������\��J�n�Xn��1Z�*�6V �1d��WX�,c����^���OQ��/^uY=wH.��G׈6�B�,E֛(�t��+��$�wˋ������(l�3�WYkjvS������;��f4l^튌�+p^Y �xh�kS�@�y���9��d�S� ,8 �lzh�G��Ry�up'"S�}�6��}rspZ�6�Z�2�AO�1�a��n��<y�{�aAb���Ufs&X�����8�$ǌ�AUd�o)k(�����XۙU��eT.ىS��Յ�L�˖V�q��J �bQD��f9�\pU�p�A�b��-E��Q����6�a�ũq�Z�lQf��#i]J8����WU��cXU+(&���`����h���sV�+�jdX�m������Q��v���0�8�Q5�EH�11��"/-�+1�L冫n���b��-Llƕ�)�f�Q2��2�l��J5ڸ�fq\��m�L�k�&6Jf;�λ������^(�۫U�̘w�����K�Sa,�!m
�Z����z��ͺ�Zw�f-_=��q�f0T�"�����٠�!+�!e��3:,!"=�ʅ0y�]�M�u�X:)}Ǩ^j5s��S�4�i:T�u`����V���a����-W_�z�W���:���XՓҞj�:*��<I�XP�X�+y��=m����
���
ӴRs�7JF:4��<�Ԍ�}���	�:%$�:'\�l�/*�*���ε��+j�q�u�n6lX�B9 ��f2�	�Ís�HLJ�
�6���VQhᢠ�t5���\6\�F�ˮ���v���N��X�G"�#��3��F8m�s�_�[O���ks�Ԙ�j"\�%���w0�������t����d��t�84}����B�Ӄ�-����A��Ь喡��ѝ]'n�I�ӯcj�jx��v9��c�ݒi��h� ����K��DB*i@�����Ё�4"p�����&�YU��<wKX�
ŕ��a��S�Ά*\���<�pdO���2P�P��*�]�1�v�}�[�+�;X���S5��#����T��ݞ����e��U���.X�%m�5�쩶�S�mS�$Y�CظA8�F��
���TM�a�ƫ+;�58jO��k�HxVW�|��5�/��Z���+�,u�a�ؔ��2�Wn�KC�87K9;�a�U�:���h�*����k�{��:��~�#��c7'��ێtu5�Ō$`\P�9�G�����\P�
"��sU
�C+JCF�5�k���/x1x�TP�z�C�V���k�O��<o�o��˽�wS�G�L�y[X��d�VM���fR����Ҍxm��I��u[Wv�n��ϧ���M�3*hU�-�i,%�3{�Á�Xx[�9ܹo/��syx�B>� 谆�0�	*p����Rێ���Zï-�;�o�ۇ��R���9+ʐS�3V ����V���g����M��<#+U! ���,B �׻����Ǌ���Z3��h�tt{
h��m���Ϸ��9�jQ13�t�:)�((,,C�������njDJ`�&c ��*w�`J���HfZ� ���y���8f,xE�:8V�N
&.c'A�?L�Kb��R[�B%ռ���E��an�T< �7ƴgE\��&#�_enL�����ʥ��HUߗ�f��-KW��F.U�ܱ���;}�����#SOE^0v�R��k�Լ��/7�� A��.�lef��n�u���ot5�L���vy��ڼ}�k��:C����K��1�P�Vt�Ўs�Q����[r~����oz�"�|������u�� N��t�Y@���wrV�r)�>q��d,>����2�Юz)�jT��t�*�_z�5�CF{/M��6̀4F#��FN�J]��H���z|�ܹu�7��V�Z0O�0kKGCX>9������]^��g��U�U��D�?AS�WD�lFMLL�r�v�\�D`�:g�uLhC�a���u/zT�o����bv��M�6�� �b{�>(V�^9p�G삛��;,� �'c��̬�W@øL�x:���/
jѲ��/�p����"�]���%N4v�)�%@�/MĞp��Qs�Ǫ}j�m����pG�V:Ԇ
�2Ҳ|��ҋy��r�JG��0�� �V�C|�3iD����Ug$o�z�K2I�Y۝ty���H>�|��@)�T�{Z	p�P��u�Q��Ե~{�W[|�'!���w�蝞����Q{y�?N��T�ř�����i����	�� A���_��<M2�_ 3������(=D��Z*.\5�$5�P����p\ZU�&E��ԫ@��ƌ��D���iǅ����~5�� bgA݃˖bb����<���sN3�ē(��:ł6�!K/��!�4#"�r���b�0cJ���(co�=�ܛ�0�E�0�ۛ԰�NduX�**&Z:Y6�K���u�CY��<8T@�;j��i����8m����ejԄ��&ph�DΟ`���� E����W��&�
�O�{yҨ�f�.�X�V�U�t^r�Wk���#Zk�g"ecѵ��+����$���}��y!�A�)
�;9յ00��w�8*��"�3;����!&;)Ul)譥�9r�����l���,1�BI�!i��(������7+q�K���T4J��SÅi���v:��OJ�G_�e�%�"ќ������u����P[�4�b�}�4t�Ԉ�ͺ���M��"��S��(s*Lp�3�+�+�S��RD�"��`U�`UhUܬk`5�V��Xt�;jq��r�8PkK'G�nxy��&��:׌dP:���J�:R�2�{�uH���j�q��FYC�v�2Jڍ�� l+r�u�ѣ��WxK�E]�l�w_�1�^�� "|��(PH�$b68�xxPd\U_D���\�zcEN�3CdƣH�<>�rƌ
�A�NdqȞ��.�+�J�*�T�c��$�'��=�2�@x�
.����e>����7&JF��ݣS#r|���9ڽ���0v\��[��Y���@�19?}�{�t�}��K~q���A�,Wu�Q�|��jY~��������`|X ��XNT�����`�U��xVb9A׶��ͭ�Z]��١�"I�)� `؛U��%�}��y�W&����N��
�"�^*��ڍ[��ɧ�S�d�'����M����l������ÂyO�`��b�6����Ciüd��맱tł�,wL|��9)����Zh��)���%l^y��U�<<$m*M�5��Z��2��!)�����cH����q'E@�$0��&�![3p�Y8P;��ٸ�1og	�d�,袧Ǝ��,O�����-j�c0pm�
��/�+"��V|�4[�>?� ��L��[!�˻��[��B�y&>�'W��U"W�{+;�u+�K~��yP*�ۇma]k��&�`ܼ���m�Z�˖C*�K�"د���d�×S"������oo8�,6P�Y�lW+�rԾ��:���p!�nϐB��8 �à�:��|�Mj�w����8�F�mhc`��)٩�R��p��COy-/;���~6Pq�4,P���\'�Z��ˊ�
��rϨ���k�w��K?h�q{�+i4��D�n�@�7�N�y�rzc�S��kď��q@��;��*n:Zb���&*������p��X;�e�F2��,��;v/.R��*
[��h����D�ϽC;:P���c�%�*��L�Ӿ�[C��;+W'�/[{(x���F�EƣD+>��} V�+7]�&ӏ�-�,7���fk�È3}H��v=WVd8�w�4��&왦��8�RN��'��4�=�����!��2���Ȅ�Jݾ�[ȋst��Y�炳&5!�w�]��S�֭�2�'Ҹ���w%�LV���s/Rr<�닝jcg�i���8=5dM��ڧ��ׇ�P�M�t#x�����L�N:���U��r_��Ym��v��iSw�\���J@���^e+��cU8םo^�\�x��f�����\z�1�e�9;Q(��o�1��6�`�c	��W{�{c��s�t���O��B�.cpƩt�9wbkd�˺S��M��k��u��ǬPزV��b�ޏ���J��B�H6T�;�f��f��1Â���܏':���r�-Ap�G�!1�!vm�Q�w�4��΋��"R(�-��ݚ3a�r(�9���ܾ���������NWJ�W�]=���\�=<!ݥ�)Ǉfɡ�孽R���8�K� ���[w6��t�ؑ��)u�m]��1�$�ݭḡ�L]�;�1�Ŧ�K�u�d!
�7I��y���!��*�<��O����)�x�+�uE��}Ry�Y�y��oJ�F���ի�Ef��N����mR��7��[�}�1�P��>��~VՀ���U�uc/E�������g�P��5��@ƌZ�
�ୗ[�/�	=�Y�B�t� Ms��R���gEա��+�����Z0W!��ɶ��-Nű��؁���F����|j�#ZWQ�'%��β��E��7 �a�vRt�fI+�HNX��%]��"�g׺FV$a�����n�Gi��V�[��(�V�TE>��C��jk�'j�z"���H�)ܱ�F�X|��>��;�0W�1�b�<!�vn��ˆv����e𐷏hm�`�:b��Q�ϸ�JE�{7U��/6dN�dǉVQ�J��Y7r�;� �a�潽o5*O�ܩ-�g�X~�u�����[mϫ9���]�8x��6��ٻ�S�������yD��)ٗ���-�a��y��y>��h$���}��!�#)wYǃeۣ��W�N���s2���i�N�d�82�nn:V�x��,�w-,���l%7N<��n�&4X='�RaSGQ�!�&�ood�c�G�p=���sdj�*�Q��
��˩f�k�h'd`V��[��ʵ3(�0,4�Kx �0��rS�ҵE��Vk1�4LwPہ�vr�u�A�n�0����V,�b}2X�N��jͳ�M�5�IO6ԫ����VU���H1�8
�G-���˷���%�,A �T���̰HC^�su��B&�R/F��3��w�m\��n���i�I�F�^��B�PTY͗ X����ȨS
�8��*��*���\��a[�%�鷻t���۸l�Icn���,m,M�66�w�V��FUI�5˵:�h��:����sP]@J��Qr�{F67��J�;�eՖ���%�L��۸ל.US[p�����(��V���?��8�KkZ�c��(�Uq�Yu��:Yyq�F���KJ�h�Uܯ0�r�B�r��a�ȹZ��b*cn7F6�R�mLˍDJ��.f �q�\s(��Z�-q��M�P�T�DUr��(�G��u�w1����XRرB���̢�l��Ɋ+�Q�\0�1�VV�ʧ�.�E̗.\��n<p���3(��69q�1�1Qu(�F���,V(�Z�ER��e�DQQpJ64��J�A�\�9m�-��X�%ʥc����K�ƲX���[F�S*�V�_Ȫ3�r�H��Íg��ce�[��ll���Er+9��컏ɳo:(̑M��!y��.���7jk�mU���=�������5B�C���ȼ�g�h�<ۄ�G�sȃ#��ZJaO��o�+��]1�z��ƫ�]78��N�{��m�"�^l�)R��9*���Ы��昼\G��D^lo^m=��X�	�)Uk䨿"��q�u�ؚ�x�6��M�	�ȭ��o�Ӏ�Jk�����p��e�Y]29�O,��+�Ч�k��˕��`��1������Q�O�5���۵Q��/� 	[ɻl]n){Y{q\csq���A�!u"�U��N�y�Xȃ�j6�����1����t��ul���E�p�N��˚4tGλ/�B�L�[�aI����,��M�8������숫�	��I4)��N�=z%�Fwj�����{ѱny�M�����Y�J/={�İ�/��J#��q�Bxޛ���Ⱦ��9���o2U�&�d*:�N�:�r���a�	ݠ/��=W�_k!�D���6��n�&V+z����sf;�awL탗��	 �u귫e��[�1<m>���
yTo"�ѝk[�EK�jM�v�G`5�yWJk.����;�F���:Y�����ܝ�5�����{��;2k�Z9�UhN�����Rw>�$���5o���c�=ۍ�O}/��l���m޺������1!Guv��0^��|=�K���xX�^=I�\�(s���H�H��O28�dO_O39;4w2�ʨ����l��{�z�ت�k�?
[�L���gWZk.�l�����{�҉j[<W��L��L�Π���3�������;�o>���s>I.�H���v?RfB/�T�}r�,ұ��J��p�d����t@�o���ͧ�e���j+����q�Q�æ���x+M�q��zGo�p��	��h��q�(u�ֲaUX�m0�#{M�����K ���+L��Qg�MA;}P����8��J[h�W䷷b�]t�a#b`�ϝw�A��j�[�ఞmO���*b��t�M���`E��̼k�7�P�,[���[��R����q�T��>n9�#�t�����ٛ�Pu8t�����v��կ�*	��j�<�,�ٖJ�0Oi"�|�k���}�őT�'s���˗o�uf�)�eʉ�{s3�7o�[�q���g�Q�WP�ʛ���s�P9���.7���)��c�+�+b��%�m����Ҕ�D��,79b�ٽT�F�'1 �-��4�Z��h!XL�/ؽF��F���ktm6�ފ�1
c��Q�$�ʜ���>���Oګq/iy�����&��u6]:O���;��8�G5��>�y�x�\��8�=; 6i�\��;���QWz�����u����n�k6o�ʜ늖��Hӎ+kzI��^:v�/��t}���t��(�I<�o(�7٪`�ok���b��(+�4��Fko��y�:��j��p�7Bh 0���)��Ldy�ҟ\
�B���r�N�v�>���C��� �iz�����M=��-��j�;g�:�o��T�?B3}34󝺖yZ�i.�S��xZY�}�Q���-����?�̤�N�<1y�׽<Ir�%��z���ʋ��U��}��j#I!����7m�kr���{~Ϋ9�(��lཿY�h�@RÑ��f��ʆof.��&%��]Zh���A���˻؝q�줺��2�SsK<�u�K�ҫ6Lg��S�)��^�2�l�t`V�������U�8���rՓ���,(b2H�2^���}�>���H>�G6%]k����{ ����u�DL�4�T!89X�Z�f�dh���[�SXNc=K9N=�4��9���}��[ؚ,���Mͯ%��_����/�ي�U�����r^��j�^�5�9h�Q��UL�s�ˬ�\�9M@h����a��Mw.����w;N�yc ��W!�pI���a��5�w�{1�5�N�ޤ��W�|�>n��U�/w�$(�{���십W��ǝ*o����<�����>���gO< �]�^`X���tݬG��q�HY��MG��H�N�y� C[���x�K{�y-�j������l��c^������oU��mp���}��4g�S}�=�n��1\�e+�E`ۉUتz�h��g9Hr����z��R��-T���r�hD-5mf��P�N�;N�ՙ�T�g6�L='����}3���xR|t��`Tc�O=�§���,���S���K���r�$�������Y���[A�Q���p�"��꼍�����vd;]�- �}�{�6-�=��9���r�5�ȮWLTy޺�����x=����L�y3Zr��Н�e&i�Gn�*�>�����I�9eȶ�>�K���(enmǆA`o.*��o�$3ď[��In qL��C}�{���S�����t=����<�w���փE!0�r����Z^��{�S)�S��o]y��~}�����ʇ;<U�T�V�O���F��;o¦߶	ޚ�U�3��j)v��wg_4!�s����x���g���[O���1oǨ���y`:�-�w_=����T++�t҇��nu�uJ�jaӳ;���Mm��Eɓۥ�F.����ط!4v��r'����P��ʱ�����s�z�'�c �w��Y���为9D��6̖M���a\����t�:+��v��)J�/t�:�eP�z��+q��%��Y��J����X��MFI�>�F-L��(�L���{g��R��y���w�Z�$@��rrOd�.f�W/D��}^g�$�DU��%�{3�P��ݾ���{����ӼMm$h#LZ�yͺ��~����65�z.#��9�,;P�uw��w�7�=ta>�f�]Z�B��wv�>���ɍsӻ�J�V,�X���<H_7���hr ���X�����@�(xK�G���2�R��Eb�9y�\�d��r�yÒ3��ϼ&:���B�5���Fz���"'�c�7h{J�����7�5��ǻ��m�)� �F�q6O7\W���	*��Դ�i�̔���)o/t<��Fal�T�6���\\��ϭd`�1�r�vk���I�$�9�T�����+4�Я��5lr��S�<�ln�+sW��(�^��A>���o����� ����C5��&M51"T��{�=^,���jӔ��TА૥��E�/�v!�V����r�lvgt Z��=��(���P��x���txn������Kk�i�
�iӜ��E������Zى?p^���!���(<��r��]=8��:�m����J����y碮f�}�m�ee�/�A�x���V��$�ڡ��Q�Zm�3�ڜY�%p��IXj���1���l��ymsI6�㙕�K�1U:���J�v\��n��{G)Lɢ�%�b�%�D�xE���\�y�SVt�iV4+��T�;��}oy��p�'�>}i\#��U6�WbsY����c�Lee��.��3l31ly����ty��gE��57k��4�����etޫN`sW!)��%s*.Cj��[g�)�����D�^���T���oV��Rq*�b���5����뗐�/G%A�����nL��&H�<Ʃ�tpX=�΍x,�JO:ע��<�о�(2LxQ�B����U�.F�{����ɉ���4�(a�)S�T�٩�]�6]���E����h���]������� On�v)���u�D�ٍ��]j-C&[�$a돲.�ͣS���F�^��Шyp�\2KC6*��6u�ӵp�RtM5u�'/J���.2�0�x���\���±N��ƶ�J��HA.�hK�b���U���c=;ݭ����s���A�z|���E���s�A�!n�N�ٙU��-�/w�&��.�v.�7R�����o'f��\��6c�h�jQ�72��MrY�Esg>�F��#��,�'�T5c���S� �8@�?k�Eh�ډ��Ym%}|��
���
agڷ�"��%X�����h5�ѳ�9�ӥ�-L�Ž�(�
J��z2�i�鹛H�����U��p3~S���C��ވM�e1g���9[5��`ś��ZC�;\Y�p4,�V��+h�8署�gK�.��㙹�TFDj�y=8��P1	���\p����!j��?*�e���ܴݲ�0���?~�X��+Km0Ecl��G0��v��Vv�Q�����TQT�js
eWK�TL�.U2�W�ۋR�kv��e��53-b��j5���s��1&ff2��q�t�ݹi�0Y�c��c2��\�3�q;�ya�eI�F��n.R�`�%J�f�똎��53(m��nn`�����˛g���ETTwn+im�\���ֳZ-KYm,+M�T��Q1+m[�vSR��YciG����4�^P�0n�LS-�i�1p��e1��2�+Zب5*2������R��E�QE\�Lv�U��k,E�QV(����j��(��R��V�<�yi��,R#iW�Y+(�QkT�X��X%���F
��(�2�a�7��}\���ér���V$�ڏ�X��mܮz�8����-�!���L�R$Ф������+W���{��֗��VF�8�Ot�b�M�3�$CYn;�Uj1e�v}Pϓ�]z;��O��	1��fW�^�:�[N:�Mezn{�:f:}�����~�Rf�D�&��i-��`o2�����^rl=����ޗ�37!��LF^�o:�l��%�U��]~U�+%?9��Ν�c-�v���s����Z)w- {�)
�bs�K��({�>�%{{�(q�A�R����3����F��M]~��LqV�n^�4���Z���^�sjab��],K��8s���r%d���]"�F��f���Q�=z�@z7��W:�	Lc���Ż����l$^F�^�g�p��lAoz�ů N��C����4�i��B:�S��hcP^jR��+wNi�[���p�z�	��P*�����yFr 	v�3���fL�ٌ��C�C�!	tp���it�Ym�8�����n�.<�|v?9���YZ���`b���!s��j&��W�!����D�ݎȨe���Ru�x��E�O�>t8����v�OT_de-Yɡm��R
�VV�R���i���HF�����\�h�=WMPQ:O�w��g��v���(��31SDVO�Ź�qˡ�p��d����.��?.�0Ϋͯj��ғ.�yћ([7�.7��np��8�eac�eG�.�C��H�q�Ŭ��=�XJ��ݞ��4c��v�sf6�.y��T;���8��n��'-E�p�i��շۭ���������_h��a�<��n��{��i�EĹ�q��ع�}�J�lν\s���l���('��}
�5FOov�t���X۾V�ޮ��$����2p{���$�wk��|SF���F��׺^�r�^�5o��gep���+���P��Mq"�$���^�����3�j�X��|��0����ϕ��ʱ�:8���*3��fw���S��,LY��/wb��J��0̄��kFp�	S�2�N��#o7nާH.����`e9بs9w��:���o�A�i��]:E$4/0�V�8�1ݾՎ�L!��ZZfPp��aw9�(g¬j�w������2�j�^M5J����r�l��B�k��W�J�*c�YB,��^"�q4 k�/��߽���+;��x`���?F�fV���S�"������}Qn�*K���Y��U+�䟽�ج9�Z�$�%�3*c���:F���nq��l]6�\�yVɪ�+�"���j��Ro2��sRB�7� ^P.�z��-V��=P���P�;H��җ��Z�v+.����Y�'/RE�ټ�7�Kz�%m��ӫ;P#�CX��������"�mv�yS4�=rj��\�Ł�|%aKtNJO*A��N�_�ĽҊ�!ݘ���'=�gW/Y*��[�[�:s��Y��}�z��E$X���YQ3�}���7����{{�ߎ�=TP�mRZ���>���8�[�[��n�M}S��lT�K%������n�wLN'ǯ���-#��`��	�F�������O~~�o��}��&.�L�zDЅlv!R�t��'c��ѱ�b��؛�-4��#�K�3V��tf���r�b\�m>�d��]V���jLZي����k����>U�df
�5�R�Dx�>�P��qiZ(��K4Y��z$�Zs��t�R���:����[��Ȼ&��W.PyjY��t��y�\�m���q�"boI-t�S�j�1���S�_I�������:_sJ�GgW�/����˘�7{D��-F�[KB��^.2��
�U�҅l����T����U��̐�ڕ�>�&���鏕�{z���mOS!Ռ�̉�0��V�'�y�I{Sg����E8�R��#jFG�ԥ�����:Y�P�a���s�e���?�O,c͍����:,�Y�6y���^ռ� �=�Vp�2��-__��.t��:��&\�9mew���k�t�xL�&�;�Yh� ~z���\��yV6Y��u�4��Z�[��td�3,"�tɶz�����Sc��ᙧ'n\{(ۈ���m��ރ�8{���H7j�R�jָQ�`ۉkga��p�z�⧒�ӝ��`���<�&ϓꁱي�]�$�c�Ӆ���|��`Lg\>/'!��S9+3]�Q�r�5�ݽk5�o=Ϳ�Tԗ����=c{gk����Uޮ}���|���r�k�b��7�<T�N[ޗWU����������\1��o5j];;��i��;u<�uG�&jda[�]�oc�%�,v.�t�^w��OPV��y�Wz/gn���kvC�Ҽ���d.*��в˱(2-> ��H(F��V�SK#:p�-�(�����"6s4ی��]Z���t�2b���%|$ON��r�$JEds�f��$f��l�j�7L>�;���Kӹ��Y���죜WV���Z��
���]��\��gtH��N�^����xuu���e�{���j�����s^c����c�Ne(�}��3k�|�,*����t��M^V�iW��l8<t�:���G�S��
/��${���x�@(tyW���5@��	xt^3ลV��^7ꋂ[p���I[{Z��)�2Wt<}��RsѤ,z,���}����n?^w:<�!Ʀ4�Oe�>\��O*��n�9��^��F��쩯df�N.�.��X򳟚��W��tx�@q������Z��i�B�M`�a�h`���G���q���'�L{}�NrD�(d�����xf͎܅jb�b��"�`&�2x-n��~ӕ4R�����{R͊XW�Z���̌����K�[ϗ��Zcq{�T�N�]�U��a��]��̻�ع��~=��o��\ߴ�-㩬���S�SbmuQP��OΡ�%�HY��3s����o������Ud�/U{5S��#�����O�T�{}�`Fm��WSC�us\C���t��\���ɒ�kk�G���6�������t�m�;�$���m�V�}D���̽�{��^G{��/rd��3]Ү��:�i�,D?��J�a�S�6w:�����-g�6��y�Q��ɼ7xi�lX�%�*�j��A%�����U�\�}�Ĕ	�%��7���*�~��Ov�*έ�"y�v:��A�swv��W�%0�y�j�T����l�OkAl�:w/��#���^�SI7�
n���~˒޽���O���V�[��[f9�_d֭w/"p�s�ڹ��&.�Ye�Mh]5{
���R���`��3jcT����+�l��:����6<3}�3����CַƗ�<W�'��E��hedᙑ�^�H����\�Q�����L1��f��\|g4�
!te�;�i]q�106�$^�
b""#�%)�"!#��Q��K<$ ����O𔱗����&R:i���/,��E��A����oF�DzC9�������?�o?��Q�����I�"!�@�cl�Dj��_J���w8^�Ju
Se�Lذ��7X���΃�~�Lb�����x\LG�/�{��(��|R�3��l����h�(�"�@� A��b1	%����E��d�`��i�BG����&}NE�<P"F��DB�%��վ�(3�.�Ss2�E~q��Q#By��Y~vX�d�4լ����Eѕ�f�e>$��Ԙ�!)ǌ4��ga*�E�����QDg�� yU���zd����:e����!�P+-�y&m5��1{��A��M�`e�@`%��W�^Y��}�#���qo{_�F;B* "�d�&&���2�������2��>�4�9M�d�A��.[x���wLր|]�)�"�;��{i��(��iv���;��!��1�]sF�ܒ/�s!�!�A�x
 "O�E�P�$J$��l����J�0(>%O�4AB�SL�"`}�6dj�Gȸr�QD!hHhZ@�́P����N��+9D��A��Q�&�k#�C8II4ZR��L$�CC0��p9�Zl@D"Ά�=X4�4����b?~����^k��sI�q߬1�Lzp@L���׆��	�������KBϿ�HQ�99�Q�f�ޒ�%x�����DBK�@�c3?�d�4g���|oM)��32}��h���Y��R, �k8�.9@Ӽx��@R�@�C������]2�E�L��(��o�l(7��6$O)n��\A�Б�Y�{��d[���q@�Y�P^�T	
(����H:���imٷ%Ch�7&���Y�C��CV�b������7��B��@=a�!xa�8f���w$S�		gi��