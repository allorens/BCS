BZh91AY&SY��&��߀pp���"� ����bE��           ;��
J�*@ (kQT�1T�*� 
%*T�"���P)[%Z�P�AQ
*U�R+Y
EUZ��Ƞ�vh����Km�DPP[����[I"�EIUQ�h(�V؀�Z�@��!6��A@ʢRU*� 1�� � ���-��J\ ZR�Ԕ� T*EDMXD����V�յM�T)*R!F�5�T)�*AU� 7
U�   ��Q  1�:�|��ݻ6�ImK��;m${g��mKe:�0^���J*-K*��6�m���j8擲5%�ݒ�JۓX�jJi�����J�}� ��嶩()^�=��4���r���!n���AH�^�^��H�U.��y�H��+�����Q��;^y��R��J�]��u&��瞩QOMS����a��ER��U �����UKo��@R�������^{�l��={<�B�*+�o^P�������3��x���m�ok{�sY�E�����F𤊩�V��-�	{�T �;�O�+Z���j����B�y��R�M�p���ܒ���P4��s���TG��qNت*���2�Y�U�=P�){Խ�]�%T#�E ���U*�B�� ��|5AI.u�Mi���U��-ei���I]4(�.�����u;��I�1��iCc����Μ;����]L4R�u�%�A[eY*��A �O�R��nn�j�ke�>ǀ�ٷ��(HMvGu�n��i�;�uS@�an�p)�BS���Q
�/ok:�f�l��  wG���TYb��*_>JH �� � :9�g (�O�=��W��{ɜ ��N��:j�Mӏ[�@]YT
��	eR(�[mA �}(� s�+����r�x�ע�I� G=ٽ�Ӡ�;w�}���{ϯ�{Q� �@	��z��h�R"F���%))P�}$� <x��� ��zܠ 6� k�{�B���=� th�p v���A�Ǽhz4<�{� �4y�pSN����LҊZҡ'Ϥ� |��ۀ 8u����`�Sw  �׼==5A�/y� ��]u h�=�U{PwY�C@<�  �JP$  ��R�! ���&L�C�����     T���I       jxBjjR�&И �&�L ��(�2�@&M  i� $ƤRI��"yH���=CF'�M������_�G������������:�R�ɻ'ͭ�y�C���B�<�sw�~B��靤��5ވ *�D@EO�  *�`����N�_��?� *���I$��� U���?􊨢/���������1?kؖŶ�bSbS�6Ŷ-�m�lb��lb�ضĶl`��6��1�lb�ض�-�[��-�6�-�[ضĶ-�m�[���`� �l[`��6ű�l��m�lBضŶS؅1`Ŷ!lB�6�ر�[ �-�`�-�[#��b�-�[�	l�%�#؅�`�-�[ �lcl��b���m�[ �0�L�6�-�[؅��m�[ �!l[`�-�L�-1b� �l[`�-�lal��Ŷl��b���-���m�[ �l[b�-�L-�S�l�6�-�[�I�Ŷ-�`�-�[�-�-�`�-�[�-�b��ĶL؅�m�[�4��Lb�ضŶ-�bF�m�l[`�-�lb��F�m�lb�`�%�m�l��-�m�[�6��-�m�l[bF�-�lb��6Ŷ�m�b[��m�l[`��-��1�l[`� �%�b��%0�-1m�l[b�ؖ�-�li��i�lض��-�m�[ �m�l[b� �%�b�ض�0-�l[b�ضŶlF���m�l`� �-�m�l`��b�؅�m�lض��%�m���-0b[�LK`��6��-��1�lKb��6Ŷ�`Ķ�lb�ض�-�l[b[ ��m�cض��-�m�l[`���m�[`��b�؅�`�0�l[`���m�l[b[��-�m�l`�-�l[cl��-�m�lBض��-�m�l��6Ŷ-�b� �l��1m�[�-�K`�Ke0m�S�-��!lB��Kb�-�[��0b�Ŷ)lB��`�Ħ6�)���[�!l)�lB���Kb�-�[���i��-�lc��6Ķ-�-�lK`�R����
6���"%� m��lUKb�[؀�"�Rؠ��P��@-��lT`�L-��LQ`�[� ��V��@�*F
��(��U�(�@-���U��� -���B�(��A�
� -�l@b�lE����l`+lPb [R�"� ���[` S � ��V�
�[`�lQm�l)�����V� �ت�[b�lDb+lTm��b�Vآ�[`+lb�[[`lm�!lb)l � `�lm���-�lb�l)�6� � ���(�� �
��V� � � �Kb+��(�-��lb [�m�lUm�l`([؀�� � ��Ŷ-�m�l[b�ضĶ!lH��6Ŷ�m�lb�ضŶ��1m�l[b��-�-�b���`��l`�-�Lb��6Ŷ-�m�[cl��m�l[`�-�l[i��-1`��-�[ �-�b�6�-�[ض�-�[ �0m�LB��m�[ �-�m���-�m�lإ�b�bFlb� ��m�l[`Sb� �%�`�m�l[c�ضŶ-�m�l[`� �Fl`Ŷ�b�ض��al`Ķ�m�l[`��6Ħ6��4��4G�ժCEV[� �����O,�-
��x���rd��KsV	l9�h��3L8�5��2�-�@�;������9�L��r*�5��Zoё�f&XE�f՝窑s\�3H誆.ӫ��I�F�t��}��dx��';�"�f��[cE	T�z�vh�4B]�U�k�ehb�$t��J�&��.��r��KM'��:���8��S���Iu���4�ہ�a�-��4�h+�x]���&mݻE����-eJ�&��˹Y@���x4L�6e؊�`ƨ�ÛK0��t��or��Z�݉�T�i*��`�5w���N�,^yU�h��B�:i�2R��%�i�˫(h��*\�LeѮQ�{�vű�BlM���x��[ap^
�1Ҳ�ǻ���PPRը��'Mh�
m�=1R��fKyn�;W��[�%��k.VL*m�Cn��ey�+�u!�h!odې
Y�u���Md4�]jZ�,L7��䅺�0�S�؜`��QZF�uO�lV�v�-ˈ�,-��<T�e�)-.��V��a�xʊJkj�3S�k����SEh�2�$�ojP�ӏ�|1��.��&����̹cq֜���)�;YQ�K\޲FM��L.��ʗ��m#SE	-O���S<��^ѻwEj,Z/k1)�բ�-�Q�h�*,�2� �Ƽ���zl���(sh��ePhR�����t�;��ieɹ��z��
�U�؂8�YDK�1
���HJ������)MW�Rb\.���,t��mf�R��Vj�n �]^EJXI���NX�
8�.�ڷ�F^(�YL!L,ͪ̓jA.���c]�
�{m��z�en۱Wsa��F�<۷�W-㯯�r��7xӺt�F�/��S۸��+݌8��p� n��kj�V���t��jSn�V�f��v`I�f��&u
��A���.�(�i Q>���!F 'i��\Wr�6	�u"���G]����$X��+��(a��[ V���.�h�c2�ujN�,�P];ywM�Y�&������µhБ��[Zbֶ�j�F�I��V��U2ZB�5�l�Z�t �Ěq(+o�wD�%ϓ�Lڪ�H�feD�wu��#ѹ.�X3^\VQJ��j��(��*wp�d�`�N\�%�ۡ����v涡ŏ*&-�M����p��t�\�K#LNr5z���VNf��2�*�F��ö�a�,- ��K��j;�y���eY*�).�.�T�V74-uF�0R8C
�,�4��SY+*]7$���7�'�@7�؎i�.nPl@1�ͬ��]h�Xj�2���{��Ͷ㻛7U0��Q��e��	J-�)yN#d�nI�ʀ[8�e��u����JT���ad�m�;-�U((�t��雁���{r�i蠄��Eb��{\l9�;2�#�t���ҵV�UNk�7E�,�@���o*�e������7i�x�k�cj=��bH՛h@M���.����КLI���x�ǓC.iXMLg�)Pm��њ겑̴������iH���	n�4�ö����B��ȶf�h��*��	��.�ܼ�(f�ߨ*>��'��(�'6��m��K������D�����$2��oUfՋk
��U��h;�Y�M�L�w�M�w����7cS�wQ�j�Z:t��*��jիh"������6U������Z�Mm���R؉�R�`�.V��f��d�%S��cCrVr�KܨM��A�%���0?	r���+b��^�eR�X!܌�ȘUF��w�b�zp���T�`xe�ͦ�u�����-���ލjE{R:S4��R���DA-#�+t}��$�T^V�͙+/5�7b���/L�T����B��h��H-�5�*�wkKs	fG�ED���P�/7R2��y�%�����*��լ�]�Y�E�qڠ�j*�b�����=Ì\t�� OM<4���;��:�۫"�����B̖�M���W�`x��/R��t�C1�`4�&�Ҩ7uOYa�ض�.�7L���k�N�m�Û�|��`�L��S����[�v,×���۴sMj,�7��+�q��OY�p$�D,���n���BY�3[2�R��c��;�(
�¦,�.K�D[Ŋ:��V�R��'�q�Wb]H���8q�6�ѽ��Q�ֆb��ĢUr� ,�n�tC�3e�͚�e�н�Y@�,p̎íj�˶�Ѫ˻�`Ņy���n"#�jF@���\]��`�K4䬹�]���w)��R5m^�f�Y��%d�	��[ib���Yr̇̑��V�Y,8��c�ku�*7��7�l��Mب]X�pͣ���7B��Q9B�&�mX�S�&��sPBΩB�Ԏ��v�4�昙^�dО�5��leJ��*擻N�[�)��Ѿ2j��X�7r^�;F��9wpm�UڵH1�!���f�*���6��#!�u3Q���N��L�d�T��V/5�D�5d��(��X��4�jG	�4�Y���f�Q
M��X�㷣m��
=����]f��cfd���"�e��e�CFe�ld2����:z�Z�֗�^�7ʭ欲�&��K&�řX����(�m�ь�����݁e���XCy"/"�Eb�5)QP��V�pb�4`�6����Ѭ+��Lݐk:l6��p֛F�Ia�Nꦪ�%ݸ$9���h�Ӧ�
��ka�{d^��zc`���ɼ�JzN�:8H��b��R�5���ǣlL(�$`��U 5gέm����8��Q�y<}0��v�˵�*���ebV�7���N�ޘ�+ҭDt�
���ݫ&�������BЬ�I��#HV�)��i��R�*��Sǹ(ݺsK�4Ɵ81f���mZ"Y52�*���l��He]Ӽ��檵��w�W2�Sr%��'��g�Ɯ,Q*ǹ*��=V�P˽�F"Y�7�BEd���a^�L�X�XuP�HY�D��]���fGN��d`ϲ��R�Q'5`$v�d�
MɆ��x"�g���+kbg��I�"�8�\ԴZv��{��M>�3@j���o8��1,�Ԅ,��[��_!�mb�0K�Y�R��74AlZ�n\�{�V�j����^Q��C$�Cs2����b�:�F[.��0�9{����n2�5L�Np��'��M�cu�k*QN����"k1xk�*MG3{��;)�7Q��4��p(*l[<�L��N��w[r�!F�(�p�R���2v�n�{5m�2����B*Q��t�-t#u��q�[��]�̔2P2����V-�`��#�Rk��e3vb�-��6.���QJ$ �7��3/7��l�ڥ<2)�������q���1q8b����V�L5 4v�]<y�Cb���Y;i �*ۨ�א�m�m��nA�n�FZ�sLLZ��U�Uf=X�5�� D]�#/�,�c���y`���[O*�j�ԁ�A"�2_�V.����,A�:�����Z$�G4�r`���D1�EZ��Gz����RL�Pv\[V,a�tn҄�Fl!�x�j:�5j躧�A�CKI-h���x��#�w��;��J���ګp
t�:��&�Ȉ�ˡ���[�ob�œr�E�=�y�֛��V�L%��"Q\�A�/^^$2�A�8�l���$��$̕�<�H���o\��9u&��R�ҽ�e��Cb��F�kP�*�b<��K�Tyh++^ %<�@��-D ņ�^��Zn)m9��݋�@X�nj����VG����j��/M���vn�� e�C�<�Ѯhy�@�V�n�v�5�8bz���ø������:�gX���nʶ2�E�4�C0�R�M��E�	e�AF�Y�/m��3T%�&�m	P��1w{�Gtn������{%I<�C����w��B�Xj�YA7LI���i̸$(n��5�z��n�"S[.��V��J�i`U�ڦ0Űf`��%��KJb�B�fj���k4!v+R�w�K"ץ�p�і�nMP;yT��
iWVP���V���4�bm��,Uiw	�J�ˠ��I���c���t`��
ԇ!S~�A¥��&
#6�ѫ.`&خ��@=F�8�������+T��\Mb�17{Ma�&�1�)S�B���e�X��K�AJbVe�Dѧo) ��V.�ą�0aơ-Ũb�m����&��uo��u<ss�N�Fd
!�3NFp㭴!5��9 2˦u�@�ur){p^@&ɤ�O��葨^.�=p��vġw�힃v��廕&	�r��n1۰I{.	0:����,��̦/��t�l-A�̀��2�H�3VFy�1-*�Q7z5��1+,U��nX����¢z��j.�n˧�Ѡ2�f���n�ƔY��܌iu�uceXkv��Y��Kٌb(\x�9`\k�v��fH�Vo5	RJ4��١A�\[�U����@�Z4���Q,7�S���{�5v�.M���-�St�w������{&��.-q��f�mM��,^��>(f%�m�
t�ј�7u�]��f���
3�q�7$.y������ld��zi�v9��V��Y��ف�ol�T��)e�1����T����1$%�D9�a�;��R�t�6��Bd�5j��Xʼ&;��*a�eYY6ցZ�(B:#*�+�2V�˩(=�.em��0]���� �`n���k1`Ӹh�I���&�k��*��w�ee����k�K4ZE�Cj^�!Dt��2xnm�4+P��*�٧���72'F��*�c�E@���*�,M������O��ݻ=J���H�+D�q��Cq'�1U��o�SpM��e)n2\�/\U���M��fզ�v@K�շ�lka�=��6�F���V���b1i�n����̡�9�Fiu��x8����c�GT�ڈ���71�\*����^�]�gJCM����dX��VFaH�rػtq�2P��q�t"����`Smm�8����s���Ұ�Z��w6��[V�va����G�sB��4�Н����t�Z;{�%4�Wrވ%��x�#DK&��q��x�4�ȍb�v��"�MĂci�j	������,T�jUn���K��^�V�a��Cm�۴�ul���@�P&շ��kmҸ��>�7XyP�łM׸IvtS��Ѳ��;��pU仠��@������Y�3N�1����AN�j[��5��63�-�Ө̪sY�ۗQ�u��AUb��eӁ�.����е�/2�f�U-OY��6�e�����iZ��l˳Z��޶��W�[b���yu���H*���n��dG����R9r�mL�JQ��b���E�N�Y	d��n˱�,fE-���wl����l���8ʛ���J���X�o�":�����ڶ�R7fh���3�C�3ssh�R>4�[�g��J�ʴr�NP
��t���
~cy[�I%�-�ё�95X����Zjf��ܘ�AŬ�f�$ym���GSD�W�̬�F�*m�[�M�,���ZTԩ��b��(\�0YcY�Q%��5()�ւiku��QQX�du��ZV�{E���BT�β��
�ǹ��*�T�Z ���1�`��ѩ6cٚ�(HPO�nY�26�&f�r i�uv��>��%��m�n�cN�}2�{F�Kሺ��ݭDf$i������j!�dk�5��e�Q�ʍf�Se%���
�r��`k�0^<�y%��2�&KVX�,� 2���hOP��js��/Vq*�n�z/f�.#���(:̔���p�6���IZ
ڹt�]J���r�5�Ɗ U�Z1M)L�5�n�T�Ka�Ȝ�,Jڭ��5-SJ҉F�8�u�����s�sR�%Ѷ�Z�m.{8���	�=�p��$3�^̈́N�;�uq�,��f�;gY"�Y�K%����"���fX2���7���T��"�J,�����tU�a�ҹ�7��l�csY�7ȥ@�y��'v�ۀ�l�`���/641݄�9'R��(��z�i|B"��(n�1i)ÿ�I�o�^�����ZMzԥX�,iĩ(�T��\M�'(/'p�f���\�4�;g-LSjt�Ra������-P*���1�AC	0�v��l�=3!�ëAqd^�Z�Q��%1V�D��^�Y\~F����[;�"hY6��t�f��h6����ւ��q�ӊ����ʜ����t2��C:��!�n�������,�/�di���±JY�R<�P�]�H�؊X�Z�s.X�e��7f)�b�y%r@��v�x���@e'K���Ԑ5iZ��$�z�~'�$C�s�����zS7��T	I%t����ȵ+H��(�$ԝ�-�$sO��o���r"��?(�������y���m6[9�B��.ˡ�U��2�[�s#6��x�$�&,�b;fa�&�4�r�r�EGrS�GfF�F%���}��*F�ո���\�<�q%i��,j�SR���}�M&�Qn��Q��:��s��'���.V�%ܲ*�d�sM�r��Ν��Ҩr8�Eb0�u�҉F�դm4�\KmlD��ũ+KR��ITX��1��Ӑ�"�g�UZ�<f�BP�"�Д:"�*��R�	'g(J���7I&�D�g��,�g3(m>��M��#ȶ����R���P:m�ˌ���1�W�֧7�C���0�e�i�/	��4��C����L^:�h��jW��p���zZ6��'J�(]�U}���)�
�պ�ʵ6�Q-ٻ9ۮ;ovrW-Ea7t�Z�o�E#�E�g�R���4�5`���Rbt�[ă�
9�LUK�0sT��k�]gx��~�A�S�C����Myw��G[t���x�,ŽD���׵~�imAs�O��M�][E�I��}F����l��;�8�*I��?Y�T�v��h-���=�������7�{������}?xT��ߥ�f�}�5}���Nwwt�7��pt���J�nf_'�n��c���A��z���%Mӗ�ܡ�X�-]��U��ηIT��������_k����Q�XF��,tqڜhŝ4�x�:��5� �+�w�*%A$S�5������J�EA\���|0�.U �W��ӥ�7�a	%%�Fu1L%R�n���H��9���N�q��T�Ԭ/^�3�P��=v*1�L=�%N�Ȧ��Nt�)n�㙹ٔޛ=9�L�5����kؗ��4:�~!s�Wk$��7E>=F�b �P�9��s��W���6��r=w�o��V�����N[��q�Q�qw*�1�9��qe�ʃZ*c��I��)r��u[e���#�\����,U�_��e����-�Eox���ww�����]�Yۨ2Ly.C� �ǉ�م2Z��;Ka�O����,G�PjRn��T[O{m���/+�.����w&���8c;�);���7�2�3��u�6�jv[!�dH�u��d:o!-؏1���y��E��@�mK��.uʤ��s	�8���"�*�;B��{q���+�vmM�6�2�o2uș'l��][8[Z2V�a7o�.��iMz��X����z�p��oگeO��TT�|�5TwB�4zle'h���'%G���&v�@���k`�!�6q-oN}�]��Wt��au�/�u4I���uɚ��G6W���}�,��4����ͭ�R�EP�g%*�\�(��Kx6+BadP>�d��[�8���-��ͅ:��[��:�����a�2m��G��Z�R���ݧ7-nE�^���8��'��������s2\��Û���#�4��K#T���N\NSZ��z��5|9༤��qci�{����káʴ�{""����Y���/gV���v-]֊�f��E���|��{�י��6vؖ[���"�,�=�����ih���Ņ���{-d�j�H���A�|��R	u���=��*�P�����=�sX���CE� O);m��.�E	���-n��\�^�ܒ�Y<f�1�����GMn=ܠ�]�����A0K+���c*�]em;�P'��>x�E�vo��λ*�[dr�0��Q+5�t%��MgKPEՒ0���.�ȼ��؈wf�/6�!������*�L�{C�g(+���q�P��	�*Y������fF����:4Tv�nM��pև�:��ěkj�D췷���Gm��54G=�1 s����͎�sK�x�N��OA]$2�fd7��Q-c:�;89�H�;����^�v�i�{ٯy��^�J�N�:v�J��O�Q=�ے*���o�ID��U!'e^2�\��)�����&V�����Qfa���p�<V;n�_2�j[��Q�׵v1ڷ2�H�f�*޴y޵)��oB"���53^v$�i<ZK�[�x����u��΀�y�M�{ͺ�S�'6������!�Z�q���uůɷcy���Q�K��(�����ؖ��Y�w��"v�Ȼn�0F	=��(�q���x�#����X��/����`1�M��v����\ᏸU�:3Uy|�D�u�N�;���`�pbs.�r��3��1������bXo�X�-�����N�-G�K��)����N,�A��J�t��w}
�Ԇ�{�v��yK�VR�2���!�--��j��n��������b��##xd'�v`�fFEH|��s+�By��jt�s7������}�@���)ar��7� p\S��$���F��s7J�;�i�"��9���c�Q����/d)�u�y�q�ٗ����Kfv�R�66Z�ONm�.L�%s#!r��²wg7���6�3`J,=O�l��ݵ��k,��+�G�4d�n&ⱀ%�g1bM��M���3��4����j^5��G6v]䗅U����ռU����ekS�:�v��Y�u^��j�Ϊ} c�m�Tv���t�{/h�̳�hUk]�lj��x�t��L�[�ژ�-o6�;!�7�����qҦp�l���J�w|������Sn���}��k�A��If�7�z鶍�&&���X�o�\�ju	�.X��R����#����m�oLa�QOv͵��uBF������u�ʷ/R�2Qc�Kvɳ�K#f챢��yBz��z�X�� NJ*��kv��I9^��3)�w�9]fo���o����6L^�WicFZ�v#�ۏ�e7.��X� �摔�d�U�}ʋ�,l%փ*-��Q�{,+y��|�����\�Q���H�:�cp��f��]c�x.v�u-�skg�V	BÕ�̺A�Wa����8��C��C��Ny/���ui���}]�]�;n�ӂXB�09�a�9^Rxv�Ǖ�s�����}}ڄŽI��+*v��΄���A�J�l�U��o�өR9��7�fT�r��m�el�oج���v����]�G@�=�W�c\+���ëS�e�9��f����3��ڽԉ�j⤉�̉�on�
��9��}Z�e;ê	B���%�^P�c6����h7��/�tu.��V��T�Ӝk����ϝU���aU�Nq�)V	ǆ���pcE��v�e�xpL�jSV{^���$���r��i�p�;���P�����oj��5^Ź���#A��%+$�Nn����,ʾU���|�u*k�������l�ͪim���c���B�לe�I�W[݈�7q!P��)_v"B�Mc�9�j��4���x�c�}�;؉9���c�˒�Bi�tk5LА���W ŧ��9�O�%�Z���U�J��֠n�SC|�ݔMWF���@��o��K�f��'��H_X|��s��Wb�j՝�}֯���VE�������)��ܣg�vmH�:�q�וl�)ƺ�C��&@�^��ՊX�&���Wς�hǼĺ7�Nː7{������@�잎�:CVyw�S�T���Y�]p3��Twۮಯ��]ko�u�>���eV��
��!�}2�t{��(V-$^�[/�[@=&T��V���y��=��\+�vr{����#[c��o�9,|�r������(&y��OLD���@�%
�����oY�|�/�w7/8bb�v>�7&lxU`��q2��qP�_Eo���s�g,���z2u_��9Mg>PN���\�W����+�XƱg'[N֫{-&/V�X��D����o�-uui�����"�m=}}Zn�G�N�jv6o1���+C��oy���ur�RHc�j�M�ƺ=:fv^sJ�q��gYM���ܬ�J�j9�,�<*��TJft��&�p/p&$�=����{����רK6��vf��`�Fh���cu�z/�Lm"�؍��y{]'-�h�R싱�֬c�K���O�sޣh�I	���-�A3=`
́�E*2�P{Л}z::u�����ca^�w5[�Gp���P��o�Gz��l���L��(S����b�ʎK�IR�H(�c)�C%NOV'�<,��B��+z�mhx[Ym���Q�T��gu��f�,�
��h���
��2����u��W�o���Ğ�V�jJ]���mN��[��ײ�Z��if��]��vX�v�<em��s�N�ŗZ U֔ؼ��@��]�/�F�T�#ܸE�Qp�zR�as�Q��ve�w\B��v�)S/��l���r=�1Z�v�0,�رx��-���T_{Vv`*c����V9���t\�k��E�eS�S�Os��
T���]��i�o	�� X��̃vfEO���\��lv.�f�x&���s�[��Mnv��"�Xm짢AT)��z�]� V�Y��b���u�}��7u�SO��ܴ�H�Z]oe���n7���T�EyE��h[:U�gn�i@�T5LWV��T0���Y�1�\�����NMSi����Vwk��b��6�8����x���t�2������x;L��婔q���G�s�i��A��uՓP�=�n՜k����oK����.}�P"�+;[-����������*��
�;H$3�P5˻�;���U�;�e��C�e�a����P���ޜ6�JI@�3�;�S��=8E�f�4$�g3�}G{x���t�d�/&�)#Ջe�ԍ�s��\�ע�X��W�L�k�^�D�紵�店���F�����2nRSa�����F��v�;!��+2늭]NI���Έ��3(f���LO�.�7|w�4��lJƩ�'�����8C=�܊w�D�h�o�њ���(�F��U��Op ��,rTh1�Gz��H�K�)��)h;��#��4�<6_@Bݮ���:���)g(��]�{���Eٗb�K9�=E��3Pu}��\˕uk����x{/���8���V�B����,���z� M����,�:�2V�.��m�m�9f��Ld�>��6+j��r�wU���	�}�R��=T���MSi�/',�v�e,In �v��\��w�e��(�Jap�J���3�6:�AF��N�2	:��n�;��b�CcAޣ��#O>ҍ(XlgJ�Vj�Ml!���dC�<��� ��܉la�<n�.q̂��,��J��'Sb/�������7��Ε;�S������-A*�QY=�r�Xk�4/'us�7t���j��G7b���p#������X��|u�W�6�����\�ޥԀ1旎�m�%�twӢ�.֊�[�NP�T��}S:zuxX������Go#UJ��[.�Xk|$W��k��0��%v"'ٹ�EB�ж�܊��<��e9{Q�mԱ>�V�%��}�P-�����׻���DLh������s',�y�k��IG��gscA퇙R��G�]g	w$;`�{�M��rA@�N
7]�e?wo��"Ĉ��d
��κQ��%_3��_�i�:Ź��>�]��ږ��q��֘]�m�z'Al{qھ�UvF˖guG|Q:!����2���;�(�1�x�[�^m+:�bfT]v�͹X�$uY�'lf�p�ND�Pom��+iYםͷ����f�i��GY�OF>��N,��o<�u�������k]���ue��f�4��:J���[)��^��x2X}E�U,R)�5l�ކ%��v�u)����^�)+�%K�Ddeb�.�ek㻀��[�[o%9ϟK�8�*5���Z��驖�`5T٫GP���s�q*˄���Η��	i�`�n:�.V`�<��<�S�|DW����)u,�qa��wcr�C׵=4�p�Gm�V�K�6/A^b��}��q4J]jV֧�}�>�+�nTy��+��E�y�Hnލ� �����78�K:9�0j^鹙������7���rg/^eZϏL��૨�� {si$�ǯso�Ǹ�'��o�#�J�p��ՠ{.<�:���᳨&H䳫��-S|o���W8��IVF[͖\���)��/C��Rx�
�drn�*�#���ͦ	ᒥ*�j�Ӗ���u�C���b�E�����A�<��X�\�8㥈��+}���d֕�X(17�]�K0ƫ]-3�2�1��֘S��wPv����tr��9k��n�s���Jj@��ܸ�_w+[H�]/ru����SMf
k`*�L��y����qJ���Z2��"�ֱ��qʶ�垶��6������:�C�y���eK���Eܕ�9:4Z�y�7���xfwj��������)�f>"�L<:�6�-.�xkV�N�����m��nF5�{vbf�f�9�:�q��Ϫ�d]:���]:��Γ�^c��H�Nwm=[����N�2�]����R��e�S��p���{�A	=����µ9�1j�}������9��Dr�9�\��ގ�����=�t.\�s8Oq$ӻ���;��t�ӻ���wwrO���9�g5�ʞZ*%�o�)�Peн�y\��������kT��s
 ��
  �X|h�o�� `����n�f�˔,���$�'����/��붧�9J�H�!!�P^���_�SP�#��%l�9�R�n���C�~q������-�`�@j-̃���MOI�r� 
 �R2�$^Ða�����Gް�">��V�p�O2�� �9�P�r��J�����4�;�@�S����j=�`�;;A�tdE�FJ��R�&Es^YqL�k|�5:E>�wtH/{��)d�ԭ��#�ЅyZ�{5��ȮC%ND/�Ѻ��eMr�3�U@G������J����>3�߻�QU������s���Z=%��_�כٿ���&*=�_͢�����
�.N�
�3���r*!l��&Fww��rg:�CV\P�W��ch�T�0�F�ݽ^���O8l�w0��rI�d{w�Z;��\��밹�S,��2����3>�T	ܽj�
��^r�gl"�s�8��>BH:�fsAj9G����e` V�2��'72�޽�3)����:^��!Զ�m��5�(�q7}8���z�"�G�����2+X3�@���W'T��3�4��i/6�E(���S;Q<�W�ڪ��˜����Sx�������f��]q{������,dlҼ��|r�B9w��}�w�LK��.ڧQ�Z-2�kL�2gi琧��[��n�n��N����A0���w(V퐃I��W#t�
HgL�*ɳQ5�,��Z>�p94��WT�oea$C�q>�q�#uw��B�E�T3:�q�����%1��Q�Yw�=��yq���WH*���M�0�U�cH����hj�l�me�}:z���5x�Qe���1�hȇW;�6����;�6�>�u�#�h���kЦ �O4��V��h�맵6�ɽT���H�ϓ�[��|d�`7*֘��i�X4��}��<q�q�qێ8ێ8㎜q�|q�q�q�88�8�8ノ8�8��i�q�N8��;q��t�8��8ӎ8�8���8�8���q�q�q�8�8�\q�q�q��q�v�6�4���m�q�N8�>8�8�8�qƜq�qǎ�8���ێ8�>8�:q�m�q���q�q��8�8�8��8�Osz���;��V����;6ٹK0q�.��\2�u{On��KQ'4�a���"e@���J��tڭ֚a�в8��"�a1��F+#E�p�\q%u���-�%�doa�f��R��q���k:��#�
�Ǣ������u"�]�c4���!�^^k��%Jx��Y$��qc!*!)��W�Bl��:<�Ί5����]��K��w\�iC�}v�'ywN��JnJʹօ����Y�:����,�$v<�8հ���.�;[�51Z���$3l.d7:����g��.�g������S W��`�Qw4�{B�p1�ˋ0ޣ�)�:{�h��g���1W���8.��kz����Oxq:ih�>�[�{�R�]5b��x�*� j��8B-���C	�]i�T�t�ݸ��wX�X���p�n��
<˹��3h�fn7��D1 ��j�-v�`����X :�w+���%K�9�ͼ��2��ݼj-={}��IF�аKx�7��G���S�w�e5�:KP�Ǳ�Ϸ3]1*�k�p`sOY��1>T#q�QW�q����Y�X�wG� \q[�Ʋ��T�q��n��w�j^����<�u���v�ǎ8�8�8��8�8��q�q��q�N8㍸�8�q�q�qノ8�8�\c�8�8��m�q�q�8�8��q���q�N8�>8�8��q��q��q�qێ1�q�q��4�N88�8��q��q�q��qӎ8�>8�:t�ӧ�8�8��q�q��㍸�8��q��q�q�q~�w��ݍ5��^-^�9ƕ��]�j�g���ۼ�'lʐ6%�uP��1'�#����X���ٙ��^h���9�Ao��'��ɄJDHLU�LU�͆ಇ
8�؜�\ܫ��v;�Q�ȺZ���I3���Q��� ���z΍ub�����o�H�̋V�%S`H���fR�Zt7�����=ER��P�f���58�>�u¶��a�6�m<9�αQ�ٙD�鑧Ǻ�sst|^<x�Q'�x�7�v�8͇�е�vXu��h�d׽�B���������H�g+��4�5(�7�;�uo.ʒ��vm�n���X���2�+�ں%�IR� ��.�vZYJ��N�lB#�Q��zngM�.�tzx3�ɡI�8U�嚹|�����qzC�i ���IJ�Vƌ��kn`��-`�ܛJ���{Μ�,x��M\N�:��t�ӊf�i�[���̵'1.�I���o3ۙ�-�6Y�i��e��p�ҁB�$��U^u_wk�v����H��5~�˕ү{�d�|ɭ��m�n�B��ac��QU�Ϝ����w|+��$J�h�%�\V����Wn}�em�g6���M9$�(n�l�b�(����\Ε�U�l���s���ER��%X�L�dfi|O�,W�`o���^=|q�m�q���8�8�q�q�z�q�q�n8�n8�:q�q��i�q�x�q�q�z��8�8���8�8��q�q�q�q�q��㍸�8��8ӎ�q�t��q���i��q�8�8�=pq�q�q�q�q���N�:t�4�8�<pq�q�q�q�qێ8ێ8㎜q�|q�s�Y�Bzr� �I.^M�H�${GY�(>�]; [9�x�.=��>g�U�e�(�!���;*ô�FP�Qڬ뜱�����*r�5UH�:�9���Gh�w��lϡ��U�
F����q������의YA�{n��&��9x��
��}lv�b�7�h+M�m|�R�=[�T��0>��T�����Glw��f-�u���žvt�)����i��UX�s	����(�R\Ub��o|ߥ��[�n��K��b��nufF���}��Ӹa�T�-dB�x�p}�'*�n]a7����}��3w0�G9s16��B6%�1�8!3��p�j�7��r�$�.d�2H�1�y��v��[;���\�W�<�g¹�u0�ru}�q���Yu����-��*=�,��Le��tnN�clJ�-��ь�kS3�Hu㨘J�Y6��M]k*`�[@��VZ�*��ǹ�����3Y�`���{UAq�z5M{؟<;��Dc���ckKlԧq�u�V�ZW�0^CWӸ����k�[Vo�{m�.	pv��*�
id�xps�O.�b�]{�9�wS=��m�[��)=�mt��c\�|_f�b�Iv��;ݶҽK���|3������J�G�)��m�u^l���8�^l#��x|�t�/�;���*��)�-��:#pv[�s��庀��D��جa8�GF�
�QeR��,v�����( �z��5S��Ay
B�Ok�Mwe�!P��^m�x��ݥxt�7P!w�֖�H"�����Z���-��<n���xV�)г-���8�c�YL�)��a��<����s�uu�VK�n���� �Ү�(��l�iC�r��b�7�������3�Vyظ�-Ҹ��rR�t�v��H�dE���'[�{)�e�Rwv��5�C6�qr���pb���P��{2��sH�ɘ�T��̽����nu^�k�K#s�F.�J��ɶu��� M��iŤe�#��.� q�w}a9iPh��{nr��O%�]F�"Wl*� SY��^F��b�t�幅ۛ�q�t�Ԥ�p+���+���I��\z�V����*��yrWL�D:Rb�w{e*��F�j�8+!�nt��/�ϡ�8(<�iV����M�1G[L}׎�6Ooavq���!��ܽw%��Vr���D]R�64�^Y�h�w�c{�"���ɌҴ�#k�\�ǌ��i.{��S[���|a����v��\����y/�ٱ��7t���뎦2%7�Fe� o�P��eK��U��1;$��O@���wai�W���X�Ȅh>����1��(jm��)�@��&��C���w�-ͫsE-Up��P��v�����"� �Tc�T�
�4`}˸���ށ�!׬���sU���`�����Pc&S��b �\��\O3r�tv��*p�]x��ϽV^:W���py�v�H�5q'2��:Y�m���Nct��x�
�o���vX�k129am4,��m`R�v�j]� ����d|3~�OuB���c�jd0�ͫ��ݝ0֑wa���"�`�;�� �����Y���8���j��R�A��J����U��bx��[�<����)��+Y���W7��m���G�f��{R�Rl�0eU���<��FW)f�c}�ePy�f�KZq���`��4�5��kX7C]�R�vHZ]�T��0@�+1�fM�{'.���X,Y�I����k��Â�2�rcY��ױ[gj���\���*^���>J��N��BI[�����N�������
U�j�M ��]�X��|ξ�͘_�۰���|��
��w[�xi���p�DgW#اuγ�V�)�ޕӕ��,��Q�ٜ[˥D����HXݏm������FqL��nm�{raꜨI�(��_g_D;� �!��y��O�V�oF$�x�4^fn!�[�J(��=h!f�Yg�	UW���:��HXR�qɚ(��\A��UwHqP�V-BM�d����x(�y�p�������ڑNI�����6�ˡ�q��H���0��� ʸڝ(p�R���J+9D�IO����v�yR�W���6=w��rzhnof4�#��R��J˛��jBSk)��
���yj�,�(Q��7�����;E0�{������+���mV^V�mt�cU�2��,�{�-
d&����暨�3{^C}� �7���>}�$LPq��(]v��˃Ix�7Gf�m�kwN�������a�9���]�9W��<pT0t�.�����)��:������)���S[{X>�$�gj^=�(��I�O[mi�v�U�5��b�b��e��[m�`�� ���7��࢒�˛�wr�j��x�՛��.���ɶ�n�)i�2�폥��[2�GM��� ��3T�p��qꝼ�c]��ff�h�]vJE��X9:QqQ���ڤi����mX�\=挕�}*��NR+r`��*mq�2�й�X�d��m����_s�\8Ș���H�; ��n��E�B�^�7,�;�bJ����.IF[Kf����tޚ��8���>D���Cf�����e�ϮJfї���|�fXyg��* [��ޅq��ҙQnr�_-+E-�R.�/:��@hl����ݒG����b�	:*���;z�y��u̇��Q��%1�%������G�'R��t����v-��ְ��M�����*j�y·u�9���*���T
�]<7m������K:jFi �P�	B4����K�ҥ��e+e������_j�}�+r\����i}w���d����*�W˹�kx�.<����-y�7}���fx�68����S��V(y7���jiM�k^�Eڴ�7�����T��O�Q�ɾ��^����ޮX�V����Jtyq`���;hl_	3{���p��=����jT+s@SH�6���ZNF���F���Xt�å�%{�O&N�[3�;Y�e�wVT�o>�҆+"��hn�AV]2��Z��2�)�bW]��^!}�M�o1�֝F�zb⫱��tз8ĳ+���"���l���;w��uC֡��Z�����i�t�u�-B����RJf��B�ڈ����q�CW��{j;��1�_'N$�B�l�n<�s1h�*�q�U����6��NK[f����n��i���l�GH2�e����o�ť���kE����� ݩUk�뻐��`]����̠���Q���6ld�G�	��\���g\�^�S��.3�jj��,)�gf�q�8����EY�: 
h:+sk�7w���b��8�^�۫4Z\�ݣ�N�e�0@���)�p"VN�>�};L����U�[[��K*ާK�[�1c��xn��b�D��E��@3շ�V�����g��:c7������+K(cv�nv���Ŏ,1�j�xc��M}@�l��V;����ம=̂���	M.�6:9�*����C��:��L�*�����8ٽ����ج�r[�:��Z���MY1H�9Ɖ�1�D�w��hj�[g㾵h���͠�#�*�B���3����I���I��@��K�/��4wb�&���,Au�M�%�O��'��[�yq\,mk:��ĵ�p��|ub��t�b!a��]�н�5���>�#
��IB�!��6�Q��E�x��aY�ȩgoQ�F�{�Uu\�c=,$���[�Ps�D!.���>ͫw{](��V�t�r\��|�ApT�N���)�����r&3eE�p������j���R3m-.��^}�*-��W^=�AYi#yu7e�ҩަ�0ǧA/��̗E3�2���=E�|�j}7twe8��ou�D;;H��ƣ�V�/ۋ�F��:��qv����:MUn23�y���Y��*�\����H9���AwB��f�ת��xl�m�RW=p�!��9��x-u�³q�k!�K;��+i��'7P`<�����n���_oFFS�pK�j���1�7�Ľ��#�{[K$kx.%�!�#����Z�u����M ���
��J66��Ӧ�]]�Z^V$ޥݺ���S{L�h��ң5�������t�)����8��C��Vlf��|�#[+m���Aث
F��t0u�(�ۛ����f�b�<� �7Z�U��f��P:���t���k���#�)��Vn,�n�MeZ�;����80n���[�@�:u�ˉ��"���IxP-�흳���9ޯu�l��\�wy*3f��}AA�R��V�gv�ϒi�4gQ���٠�>�g�.�斤m�zt�W��56u2~w����%]����C�D��6�z�f����S��B��9���U	*��;$��S��d�ce�_9ʑU��^ty��]�Ϻ��2����n���;ǆ���ѕ����1ų������i�g<��Y�վeH�l_x�)�c�I�ι�&�<����O��`��� ?���s�/����ć��3@�$A��8���\%6�)
��#��A�K��bm��H4�(�Q)�0�$8�8�
�I�&"I�"?�NDXj�#�$�Q��!j.Hp7��H1l��Dq"�Bd$��aq0�j�$A� ���䪕��<6�D-�8��P�H�L����6�H��I�""7�h0�pF���4�1D$��ID��#)H	�B�N4�I4g0H!�MX��TM��M�Q(!`�ʂJD�2�*�H2*���2"EW̷�u��5�L����&w;��Ƿ���b�)]b�=��������c���{S�c�b�nqo����|�e���/E��!����;�B���}�U�%�s��kl(^옐O�;�]�uչ;�7��j��5MQ���5��w\����7rv�Xۨ�;i�-k*�\P�s��0�v�XB�o����U��k]x0�:�қ�T˝K��Z�J9��}�m&u��D!�og:x�84n�A�,$![������3�,F�����@mYn��+mŴoEƯ��Ȉ�qҲq�6��D��$V�6fM���-�]��

8zb眝ޚ�
�yJ˾]Ճ���Fd3a���p���i��A�<��G��f���w�����t7���	l*��9;�~�ȅ�F��4 �h�C���;y�z�"˾l�L֚
Gu�ԍ��ʉ����wA���W�R4�K&1�t��$�]���0T��#gzT�V�R��03Gv����+�Mn�D�����3*�-m7��$*���CF�l@�q]� �IY7Z�[��݂=�n�\��v��}��úwr��v�T��`�[D'
H�	h5`�T���$D�HSB
E�H�D��g�'e0�.2�b1��R�n L�4�Q�b1HBh�e�`TJJDԅ��	���I�N	Q2FF�E����ЁBFx�|M����E&I��3P�'��HD��H��#/�B�M!��<ED����U�C�f	�W��@���|%�)�䅒(	�Q@���8	h �i��1FB Rq�lƉ-'	(����E��K�C6��*�%%"h��6Ta�R�p"�CI���A"�@�A1)�D"��@�PUm#i�E�
e�L
��I@����#	"RE�B�-�m��HBB,���8K�4�qP�����r0��(�Pd��%�T|*(q8Q$H,�� (Ym����8��A�ċM�
�HxBqȑ|���TA5�=nH�Q�b56�B	��D]����MCL�D8�-���m4�@�
	I��8 ��_$%��!-�A�0Zy�xO8N�W��79S��y��]DX��7�W�1����^�x�\q�q��z��Ɵ7��ck�|�h*7�x���F���sh�w��~o������8�=z�ӏ���:]I(ڍ\4Do�<��r��dK��P�*���QTr��AJb��ׯ]�c�q�qǯ^�q���I�HH��'a���\��.���`���g:����EF���y�1�W�W ��깷*��6�]�|�q[����n���\�;Me��uB�9�����s���x�/mGwr����R}t��h��O�|�V���\��%͵�r��]ծ�{��j5���s�h����Z�r��YK��;�ˮ窮x7^w_<�
��]��wv�8 j������$+��u�q��v���v��Ӎ����%&I�m���|�x[#cMA��}�^wu-z݋�׭�����v�l뺥;���s+�\0�T��>7�~yy<�0mԸ��닫�����:���<v�q���P�]PXn�Wn�.n�.˳�.ڌ�Q+S�K�4Oks˱|^-��u;�65�9Nb<\�S�y㓸۹�bu�`ƈ�5/�����@���	�A�2����,��1I*a�%RB���A���G!M�H]�Q���s���my��E����b��J�c�Y�m���(��ƺ���%U�<]Q��@��B��TR&�$�F ���J6$���mNH[bIJ\�9!p��h�Qě��$��!�D%`�X1���Ȥ6ц)$$$�a�MH�(���'������*UB��o\�Y��)%h�i�JD�Qm&�2(I;������ w;@��]����9q��j1�4�Dw�f��G�NzZ����_=�zs��<��S*s2�E3oԞ�H���/�}�w��0����W����w��5��5�^�c�Cmw�z��7K�;��:I�K���{�$�;Oi����N�)*
�g�9d���q/�i�������=XH��G���0>ϱ�Ϯ�?owI�f�^��
�����o��D��t�c��b����<������{��'����^-^���j����}�5��	���.r��ap}]71&۸�ƛfdx�����^w���oz�[������:�nc�k�zXT��	 �Z�2}���G�b},sdm�2Ӗ"� �T�V�H��Hٜ_�zT̞��+���:��'�fp�N�ޘ�/N���^A��1�*MUc�v�}%��jY8,��B��ѓ7�&A]HF���]U%�W/�c��R�h؃�i+�\���if�9E��0�Lic��|���ȶ�V#�X^��NY��գPS�	�}r����ܝ;���=`��ɳk;9�:�
D��~ ���ٗ;��/x�Nz��ݰ�$��O��F��=��,Ăx��Ϛ;��4�=WfO���9��a��Խ�� �O��6�{T'*�sp��=����@boƘ�����=#����F��6~[l��57��v�vΌכD�� ���|�Y�`m
[Ł�:��:�u��.�5�n�m���q�s�ۏ<U������c���w�}r=�ɮ�}�{����蕍��7<ef_X�׷�����;7��,s�����=�+���]�zX��i��y�Ԛ��70L�t]�n��7�{| v��i�s�&g8�nr�7�dfw�cm�|c+�����ڎ���`�o�k��?�������z\��T��`����^yr�vs���>5%��Ͱ@4s3������"���AZ%�ɝ�W�k�;���n���ݎ�8���x��l;��x���z6;+l�f
�f�z�ڑ=��A�޲�yZ�F��;�Zyp
�ɮ�=��x��J�}�qh|��4��)Z](v.�ݫ�4��O����sZ-�c������s��O�O:Q��,f���9������6}bjݽnj0�3���[���|����]xm�3瑺w���N���lImQ&�K���ڻ���7�-��>	��߻g��J��z�}/�Y�m�{�w�VJ��3Y�;y��o��e��m���>�ٮ�����|θ/�#��wN��P��EO��4��_��Ԛ�����b���L�Xq��������������m�7LΞ���n'�+���؀"�_ڬS�[W/S�ݒ�ӇoƏ�-΋���f^��;e��L,|/��D�����w5�{k�#<r�U𫀃�H Q�({eo6��X����G�΀����M���s�U���� z7|����9k�]*�<߆���n-�h��AW����w�ʶ���,�����p]��eW���I?7T�N��r뷔{����{Om����gI�ƞBA.�M����^� xs�5�wU�c+�:��v&��ߝ�tT�m:=��O*]v:�.qe��5���7S�̾�it;o6vv�W�c�9G/��zt�޷���};�}V���#��|n����[�h��t
�vs��*����e�L�g��]ۋi��}����Ur�����}��k?B/��vvfw�%��o61����&���j��~��>�xŤD:��k^g{��f��O��9���Cw����[���ezױR�ַͥ���9Pۯ�ƾ �(���WQ���m;��wg�-��w��[���z�L��m�ܰAx*+����%F�����/_}��ަ�u<x���v�Hm~���0��r�U ��:�{�a�	;g�Y^����P�9M�kK�Oq��8���r���Q�z���"A�o�ϖ^�i���p�;ϔ�o����H:��?~ۿ������df��d���H:�(���h��<�~�뿂�^������&�՗�g=һ�T��B7N�Do�0�(�mb.��:��q��w�{=�Ԑ��2���~AdrZR!`��s�1P���Z�.iˇ�n��WR��3ڬL0��Y�������uEm#5��ğU����7�뭖V��ޯ�����$bF*����E� �TjkӉ�ޮ���a-:_i�H�N8Ta����`��2���?-�{Ә��h��_�ך�Z����j��Ҝ�Q� �����@x
�*�Fk�*�[i�K�W���Z�[;�{�+}q1����>�9/�{C��b�	�KͫSӯ�˨x|! �^Y�v�� ���
�i�z�\�8�j;^���R�B�Gn�%�Bk��~�}�X;뭩�����`��t����g���h���g������9L�Lv#�2�^#K�ci�M<L����D���WEj�ؙf�̖�n��[x�����O���A�q�1��w���C���F6���<$�ŗ]�o�.����$�w�����?y]9e��3�az�� ����w�3һs��T�ս�XA2wI��7��Q|Lz�K8`<4z�{�����9�si�����Y���ᳯ�gk��*T�&�e0N�+-��a�*��z�]7OOGۯ<�!�D����|@[�@�D�3��j�'|ոm��B����_	y��al�ˠ��d]�.ZR�pm�;�uo5�d�\�����85��y.��/
���`��ѧ�=O��M�s��&��X�`��l	옍n��]z�z��or�㦋��(GN]{�d��������V����w�p���80�6;���O���瀃wS��Y^��@��:���ܻ���6�������� 3��fɽ�^�u`a%v��Di�l��0g>������[��J�[9�w����Ae����y�7��b^*䝨q�b}� ��o�Z���_��C���2��Uݷ:z�3؂�x�E�j�~�����v�������,!���,g�J��ʄҿs0��j�H��B3zE�뽼7��ظ�o5
������о�`�ޫ�~�����^#z�B�hH��<��e�w�C����6v�m�1ވ���<d���^"D�<���4�Su���ē@����rv�b�&�9F��B���K���;�A�u�u1�@�|�ٜ�g#ׄ�$I������e���-����y��f��a�U�*�L��7�±msw�N�^*�rm;������R�ͽ�����އ9�5��ɇ�y���Vt
�TM�Q��2�k��[j��u��DX�$פ���������w�h;U�}����~���᣻Ǿu��ϕg���ے+����zsD���8��>v�#K����� p/W�w�|-xz��{w;w_��'t��\Qfi����ݵ�1���}pU;ϪW�}�W#���	L	����|7f��G�����=-�s	͓��ͬ��w�t�i7�9r�S�MfЯ�Ci�n��w��f���$�Ř�-$���vN�Ͻ>�ex�4�ptW�|�^��t>�青�]7�$�.>����"���9��z�.�K��{��{�K�>�i�������NY+���o��+�Z��S�RC'��N�}�,��!]�FvY�ﯷ=���]�w���o@�<��vnу/�W�����7D����ʝ���Xj �śAt�Y�c��;^~��p"��ӽ^�u׳c�F����H�K�Y����OG[�쉪��y���*\5K�P�2Hf,|��8;�&m��`�����T�ɔEr�x�rfj���^��q�`F*n�櫗���ύL���:�_}~�T�v󝳦����0]v�t�����͓��H{ܯ��C����P�M�묹�x��������������6��׃]1"%I'Y����+X�E��Lʻ�v��_>ٙ����� P�{COl=�X�Ѓ��=��Y���
�Y�1N7�ܽ��$��o/��w��C�F��z��3_m�2� ��b�y]� �{��,y_��/��*{�}���cb�iP�q|d��+�v������pZ9W�����
\��c�k������z}d�/ػ���T|v��rvK�W�fzk�"K���;:q�1ɺ���r�����:�f����x���[��W!�F��].��9��<�ۣ�m}�a��p���g��E�����7b6�>uC�Y���h��o����X=�CL�F�c���&A�y7��Y:B&��C�r���S��=z�}��g������l�lG>N�(kkv G;��^�ד3)%1�O�5N�/wSy�u<"S¯z��|�]E�Ӟ�;Y�8xxx �P��*A ,��:�+�wIޚ��C�Gl�Da8"䄷 j)! ��"F�4J���W��'f����W���a�נ׷����������w���݄�l�@
{�B�C��0�����$w���ź���P��̌;��ǎe�q�'�+ٸ_�[*�8������sh���/�u�_M���~>+�)�5]"ޫ�9$,j�3%oŹ��Cq��%���?�!�\|}c��`�}�{�$9�Φ���2L5�i:��g�E�8�b[@���W]u��U\M�v�s5·``��}��({����:�w>g���#|´��^������)S�^Y�Z��.�᝖�.��lP�A�g����*��<�U���-�ӟJ*]�ٰl� ;O�����8���vù̑ڃ]��4a7��<�ǋ��fI�~[6�m��>��lﾝ������1�Ȣ�½U�|�
�ӧv]��x��U ��%�p�Ϊ{�#��.K��XC��+��J�n��Й2c�7�w�wW�[�/-ҝJ��vj��Q}`��]�)ꐺY
_C%,�D��O�OPhu�jK�\�\�4H[��u_�,��]e�M�8@< *8���ַ�|;�UCa� v��b�f���I3y/E��\�{/=Has6G.��;D�蜥������ʫǜ^>T*e��s�*f���%�y5�ϛ��P��a�5.n�La��� [C>n՝��zO�'�;s|L��;���tb����+q9��^~�P��5XZh��v�A�NV�i&�c�ZK����Y�������3�I y�3�-wS��������_���F��ڏ5{�8A$�>�� �=��޺]�:ʞ���پ>w����
�jܨ���oL=^.��;Y�1ޡW�D>K,,��dcw��A�IuIײ�q&�I�4�x����n9��2#o��tgT���r,���Q Yn��7����Z�ls]�c~��	O|A0 ��${�ߠXoj&�4Y[Ji{}t�G9�X��c{�[�YO��v{���.oLT�N	S�KI�\^;��oO5+�>s)�uq�6ٴ�e�$�3��c8-!�z�-�O^2b.��S[�yGq^VĶ��g9��t��>�t8�`��uQ�cr�A.�l9Zm�Ɛ{�~]�G����P3�n�.����4i��w�l3q�ڸz\*ڠ�W-�����5�l��jT�ɔ9u��#�k�#����o/FnTt�c�X`4�Ǔ��p�+<�9���1�v\2��i��Ṓ(M0����IR���G���hM���Q�!�f�V�wu�Φ�\� �bbѪ˛YXb��֙}X�C{��/^^u�>�]y�Y�)��Y�ijW��[r����Y�a���#d<r���wAlIU��j�v�M��ժy��d�뽾}0]v��7ae������u�)�v�$ѥ/��go5 HuYg܎I����x���F;vU�`��.SUa�ݒ�&v��EL��2-�f^�d��+p��v �4w6�XC���AXWf�û7�n�r���,�+�l�rr&��>��{�]o�P�cz[����-r�UC\�ꄺt�ꪓD٠r���8sr�y�l7S�8�m�5��ř��[��G�1����r�[;o���2Y�&�A�*�<O*x͆v_U�6��Gq�ǽ2����R
3�K�,Ћ�km��y	�hit�5Ԛ�˟3rf�S� �N!]T4��E���� j�l��񋒀E!Uu)8�-.	�� ,�9�yu]�l�Q՜��+�ȫ�{؞��>ݜ�˽����ޘ�q�]�AQ�q��Pi��ƅj5�2��R{���쭽�gMh��.���bKZʺ�u�T	״�����uu,�}�s�z����4j��HlX�^�+���ݢ�Ie�wW!���u�N���[�\-:�<"��T��o���0�o�:�<���Lf���׻�u*`���"nܹ8��g`����a�+�o��2e��������v�"~�Y%H$�|�{Rr`����͇.�8T'9���lM(]t�+ʭ�g�:G:�^u	cj�t%׆�:������[ֻ"�N9�Ż����;�=*�f\t�$N�F���7ALV���)��̗�wH�+;/E��0*�>₱W12#���WK&���T���e����d,�������Ԫ�DΦ����}�!�n�K�3{�+�V�v��ҙv����ѭ�{v��J�֦vlM��O\��q�����U�q\WB����ot�{u��Ғ�ؖ�R� {�����v������Z9��u��]|Z����%��8���w�Oz�g\��a�a��[L�0!��֫W=D5����Hu��-�m7$�evR�V]�B�y����Ľ]��:��.t]־��HSrBI9���		��><q�ׯ��������z�㏯�ݶ펯��e��ǋ��W�������@$dY���^=v����____\q�ׯ��ݻt��a0�Ir~���.sY1c_��� ӎ���|v�Ɯq�}}qǯw���w��}�m�feb ��X�@�2chآ+�w�܀�v�j4`ƍ�l���Xŉ4h��ͯ�u���4W�����F(�0������r�j�$�r����r�_ܨ���7����u��_6����\�o�מ��Cy��JLi&�F3�{�c!bg��[
b��� �B��W�YE�u5n5�욈EP�j)QAIt�Y��]۳s�����\=�R���Uog2�~p�]�}i��Jhh��3g ��f��{y�,c�!��ͯ��ķ�FQ��z/c�fp����L��n�����hAs���{��>.i��~u�@�̞��d�	�O�4��������l={L���ߞ���*�J�ߤ�̫	���,���h�/'4�v����B�����O0�8��P�Rz�r����h�_]?9`	ﺘ�β�*��D|�����yC�^i��a����}k��ɓ0;#5c�� �y����N�A�O���;Y��(���~T��5d���N�x-��K�:Z✎.j��G;/x|�.�� ����M�����s-�YE��N�����ᖲm�Y寤�lB�����<��90���-{��'�����#玷�2}EQ�[B��T�=�S��E� �y���=��,�����gD�[��o�k��]"@���*1�'�c��(tߕ(p,�LN)z-V7��+��7Ya�Ɩ[X�g�w~�@�#\���C��NE���з�ްZ��)Z���b����xԧ�Z�<og2��|�d�oS�����\d_��P�����{@�!����}�t����/T�<��\�n�5�ѕ��a���n���m����T��5�'ju��Ɲ�s�,��,L8W{���t�:�[����86ε�ԛ޻�J���$��	�͂�985*�$W0�E؏��oDp;���#��8L��dYk؋3��zb���1�u�o�W���a��R�����w��u��#޾���;S����,�ԛ�<<h+�A��?Z��7���&������-�����N�_Z�k�{��nc1�pq���(s�Yp�Q"�
Z��y�|<�k��TS7=M���x�{��\F@my���-�� ��>	��"�}������Z���q֓_wqk��O��<���ǀ5�2�o$<��X�/^m/�miO��H�{��?��H���4�W@[�� N�����ާ�Wbw{��{�C���+u#~�
���_�s߽��:X]|6ⷠ�篌�xeA��*[���1�%.��U��l&�k��^��0�S�x��� Y����Y΂B�7�g8�;�f��2KZ\�a ѐd���Q^_�ߝ%�P�9��}�~�D;:��=L6ն�������+�|-��e�L��|���i?]�Lۺ�����EkמL�� ���qLz/��*l��O?^>:r��{��m9 ����E�&0�77�ף�[�)�w��K�b=���i�w��b��O7H ͸�R�iE����� �뜷R&Ϊ���MA�v�͙�_'�>����l�V�n�����],9��.���׈�w9��i�/�XV����ic����|��}��Z�E��K�����s�%���Qrh��ː���(*!�Xi��5�����V�ʍM�Ow.c�&���?.xxx�D��~)��LF$��w�}~��i�2Sl�-�ɍ�J$�-{�X(���?��#}��^�F8蝉-l}��o&W�(my)�qhe<�����RP���q�d����Z���!�_�U��}?/�
�^�)�K ����t�U�̼u�|��:��\��x��f.fc|�Ƽ@�ƃ]@�����F���_M?Q:5I����:+=6ȼ�H:fp�c����|��xgՉj_g�H��t�K�@X��gvt&�!^�M����ᗶP�����7���-���Jn�S��T�����{Xֆ��0��ߞ�xǾn�t��*g�c�C/xKV��y��/��S�FK"��9����>���x�o0ͭ�Ж����6�D� ��ض�L����]]@���hV��〳�����%%�֨��#i*���J�d�s��,�+ sy�cðf �$�}/2�K).y�>ĕ�g��.%�/�{�?��P;�����/���R2[�k�_<:t�A��La|[�=`x��齠.Q����[����^�����+Ԗn���pq���}*�������p�_��˻6>�S����iڟM���ۓ��&���D>�9k����jwy��#��$R�b��*�l���쇋��!&�֤Ө�[�����(���{�̕޲ ""�����O�NgFW[ݮz�e]��ٛM����GU<��k�P�P�v�U�/3~^�3��vL�>8�}���#�!���ǽ9Oì��x; [�pX���y^�%�}U�uK�&@X�K����a�a~-�ғ�6�f��>[�t�8w`4@bY|�������/�cO
�}�k����y��K9;U����ꈵx��/���&��"��]ǃ�=�c�;b~{�</����^�im;'W}��"����%݀:��V���?0Ϯ��K�j���*G���(�ʼMׅc�'�v�]u�j��K��Ǹ=뉩�
J�J͘��yX�D)��00ȹ�4(SLW�r��Q\G��B���a�O8�z���]Ȝ���I�X�S�Q�\�ڹ̯1���������^3���%��TYRe�����/�<go���+��Y�����
{��������`T@M�]��\��u�n^�t�����"|�.�E��t�	Lkv�J���N0D�C�Qq6�^g��zvFd�󆇁�[ܼ[���>L��6U���2�Ɓ�9��Nb���`���Jǿs�(�v��C6�"�ޟj�0�+�D8��R��o&-R���=�w�N4#��NTC��;]���5/���4^�/;�$�U�[^NA�����{��"R����T��*]�/޴ݭ�O����8�+$��U�A�}�^�>RP�k/�7����e��J�ˎ���Ҽr���jU'2pz�����>ڒ����('$� ��ѻ՘�Z�蜋��4,i�(F�Ѐ< f��]����*׀�}io��y� ��p��y=<��ݾT��_�2��&��
8Zy��s*��.�4Ml�exǆ�azx@�e�������ߐ<��B(zc͔r��D��������{��K�����7��⾿N� �9߼��R9b��A��o�K_}��'�]@�]��/k��TҴ �ǽL@Ɵ\)��fИSM�`̏,��F�q4�'��>�=�x����r�{�� n�)|��Ǡ\���>�1��F�X��k��r ���G��o\UCI�S��wF�u�J�����9�{�Q^�f(���ӌ�x�->�,O)�q;�w~�O�%mn�>g`��(��ę�!W�0O���-��d�s@��v��S��׸T_"�\Usl��}�x�f��S�u�9N��� ;9Ѐ`�T�(�l���O�v길;_z<e�emƉ�{�
׀�v����uo�����,�O|�6� �I_ʚ�J�	�#<�,c?���'�j1�I�5�/@>�����F?֚�Y1�r��8'��3�Ay����N_�[=�q�#�۳�	��9��mP���C�w���j�'��+�0��ˉ;{a_Ap�y .���o��{lu����G�N��m\��	����'�i�%[9ز�.X˼���Cޅ]��C�V��R�έqmDU��$��PN*�M\���}i�(Ƙ҄i� �P� ��d��{�0M�V��>Y�^�hg���r��8%E-�-�T�{{��
$�4��r���e
��o+����pG<>�f��b{�L@|ř�0S!Os��J�=�	��"�s�H|�v�M�Ateu�ɞ�߸��-��QxoϕS��=���>Ybޒ��_3ހkV��b������Vi�g����q����8|S�he�[��eC	�tx_Ph�y�ґBE���L��[�{�����7`��w��}W�ܝ߸J�篅s�람3��@���k���A�Jq���>γZs9�35>��;���^i�2B.�\�Me,���t{���� N/<!ywQ��uӵӥ���u�O�-:�/-�2��O�V��� kB~vCy���r�zG.z�.��o}Y�}~uo{k��{�=^i闥�]1�8��+���\^�z�0g�>��l�ŕԡ͵[yS����"�d�s����_}y��|���N7_D\�ЯoA����aq�Ƀ�k"�k˕���}`� ���ٳk��mr&���T _Y&����a�`0�6��&Oy�P�U[Z�o�zhh��r����nF�f��f;�]�wt�Vk�8�yW۶nV�mΌ�	ɚT7����3/5l��/��m�$i��zZS1g6(N]^f��)LPK�j
�z�ے�������| �1�@�1�@�1��� ����
��(��]��VQ��/ٟw�L��(��`�$��e�����E�-�����_1`��|@��vW�j�w���9����:�z7�>t���e��Mfck�8���˔cy0�_����f,�
�^`�S��]^�>�v5��)��ӶzS����o��	ή|=ll��Ę��,w��}7�g �<H�TH_:X�*��@��J��/[wVC�vo8^�r�;q�R}O"��B04��y���9c���
�S�%��r^��0�%]\�X���|��Cm�fh���ǥ�%�9O^�3�gM-l��辀):�YCqS�4���ڋw#xW�k}���90�^C���@ܾ��5�C�
%�پ|��{8 ~�9t�N��K�
ބ\XF�g��/6�����g�^*���
�>aȨ\����r�68Ҡb!����W8fYyPA�����̹�TB��&�0�]ɽ�ؔ����~�9���(s���zh���t��@ej��!{Î�7�O�w��r�����0�/[!�
�L&�ߜԤ�5G7QR��������wj�(C�mP��p�)ox�m+�	��c�<��k�lϦK�6��g���`׎a"��C7����%ecT��q�m�ڴs�l��]�;�M�yY��+h1ڈ�X�;��r�[sr�7�f�t`Wu��B��	k����l�K����16&�&:-�jFȚ4����;ӇH�oh��/bIJɸ�d^��H4�����u�ܮ��>����4*��4��4	PFAA;�w���ϙ�❓��y7�X�|�&a�q��]�b�GG$O^��1(-��Y˶f��n�\mx��y��L��`B	ay��7��TP�VM#����Ϯ�F��LG{�L����'��ُ�w�m3�Y �)�@�����o�C�_5~!�t������
3��n�0�)�+r��1_��L���"��Ϝ����LxG�:9��^���ʄG�"Y�5����4R��^CCb�<��)����*�Β�li9�zs���2�/�
<g����x}�ì�<`���hVi����D�>��������v�u��Z��	�X��YsvY|�yմ�N�G��doT�����<�j�,R��I?s~sǤF��b��{l�&˞�E�P��y� }_i�'~��V^-���q=c*��w���@��v�VLQg�a�-{�D4�PS��ރ8b��@��!2���nv���m�+uG�x��z�߻8��ۉ�1+7Ā�d��F��Rqƣ��G�Vy�C���f�.>��^�� q��[�j�,^,�"|-�S�]�%6����ǟ�w{�?k=�N���1������^y��M�F��J���A��vn���48�L�I�����F%�������~�!U���W�4}����a�@F��c�
ˬו�����Lv�x�[�ZwZ�%�fκ�R]�	�8 ��_�D$�Zi�"44��Ad D@Eo>w�５UD/���O�6 �e�T�:� Q���O��c/<���$�';�A��Z����Yw	�/����xC[%ނ�`g� �\�{ИZ��L*%�TS��-�\a�L�͔֣V�H��^���@���Z.��ٺ���j�_��{�ͧ�����J��也T�H<UjU�Ͼ���#��[E���]8%�������)��ª�|K����];�͑�v�*����u��x��x�w��>Vz~'P�P��o�i�ߏv�_��k�KR�֗�ժ�Y���x��o�>�^���3Pa�Oz���������L
=3~Էs�Yu��/=�8\� �1M�`�[������y�}�_B"Ha-�����g��zrv�>��@�s�_ft��}7?  ���;������(��A'�<'8�ͯ�\�K�{�����p�y��
4����x`��������^�'��&"�CxF�~k�{)������p	i���ƺ�-�sƄ�EEp��ez=�ey��c�i$@�]�m|5W�����޾��R`�P5L�m?��=<��>�T:"*����]���7.]U{�u":��}��<õ{R�,_M��)ƍ�G7-*�۝@jy��x�k��d�ot-7���+v�U��2y�\>�/�ѡ���V�QE���) ��w~r��?���{��w_དyW�%���oɜ�
�z����~��sK�g� �W�P��n7"��:�x�=��%HÚWY�
}t������t+b�v��)�M<��j�Gnڧݭ��n�GU�̒2���}�z��O���s�s����|�7�	|m|��-}�)[���-�4|���,����Ӡ�< �Mm��ek�o��.���WVzcL�O�{Y [z�͵@�f7�;R��9��,(�檸6��;���tǞ��u��%M����Xn��)�%�֔�z��� ��,qs�`����>��j�����{�O�aM)=�	�&�P�;צ%�������K�P^�����Y d� v=R
�����?��]��7���>L��
�x�I��i����V/T�N�iNP�����4]z%�~x`kA��|en�k;��Y�����M�6�sP>�z|;�c��7�r [/W��"W��8YRG�lo����%�q�g��Ɩ�O]���!�ˮQ�,�����& ��;\��7������S���(!+�W���H*�{5Wݕ;ZDB���<�R��/5xػ��;my�;"$��G;���љz(u0${"�Z��6]�����7�r�_�:�u;��x�����;�Pr�"�p���Bj$�!�׹H��&e�Ө3]�V���8^i�N����4޼�|�UA@q<�emw;�5��k��PX^�X��u�
H��R����r��]J����^���9��)햧N���%��oiK1�]377u�|7�_n�N́���_uc���!)��ٹJYU��wL�[�x�k.���&���w��e®2l$7w��̩sE�jZ�!��FA{36I��g^\�)���eu\=Ƭ,[ݰ`�N%h�tk˭�!Y7OM����[�=ӭL�y�t9.�l0>���m11��w1ٳؕ�vE��n=���Ig����ރ��5o�mնL����U�>]UC��!�5�zč�f#��r��$jƉ��OaD�����Ej=�垴(�3�	�Vf
�Aan�}w.��j��S](M��g.����=7�fkXsnrW苸iJ�8 ���eFB[J��[մ��-�7��V�Z�;C�[�Kv���K���R�T���Z�0�e��)���3*��du��q���N�R�=�N�=�X�&2�mm�NэKe<��@e�GC1�]�Wq����_��zOE ������q��IH�,X���i����x�¥�[�>��o�����jś�b� )=�;�\1vT�����iIKv.��^�y�}�!�u�"y]����5���s>�uc�Df+빍,�ܱ��C� �Re�vg;[��8�@���ܞ�:��p1��uךvT���$R/���c�u^�@�%}�����mR|pCN��ֵ,�wӕ١���g
���]�#΢ݤҗJя{�:�m�I�Y�z�wj�w��ҹ�c&&�N�	�C�%��[�صB�3[�}7w�R.��Q8�r�0�����v��$������S����\ɾX���Asyƭ�jt���)�gp��Gm����m>ڢ8Y���{���e�1��T�D93��ΆVZ�.@+���iָ���Rž�fC�L�2�s���%�D�M��\yH��5X�n�ɶ�`�f{;/�Q� 1Q���G26����R�?e�ֺ��ڞ�˜�baZ@������bt֮G��+0uYa�o��iS�M�]�5}%,գMp:Ng�M*�bHD���}z��}�̂����NoP}��Z�;g�-##�훻k�k�F���W�\�/��4�&��J�l�[�����P}��ˤ�c{/M^H��>ZZ"�ժе83�P����Q};\��5�U$�gf�i���f�E�7M8�ϟ=����7�/�$�֮[F4�����&�:ov�nz��.q�<v�����n8�>��]>��v��DE�	D�5�ni1l!$[��߻�m�ӷ�8ێ8㏮8��O��ݻm���V1��;��(@$�BBA6�����oq�q������_]�v�qI�L�P�6/��'�^6�+��34h��s_�r�E�<�>-r�+�揪��_z�V�1��|�����4��^y��z�5E^����[,[Ƽ\9k���z�s%�E�J��Xѱa(��m�5�c[�׫�R��Bߪ���~˕!7�R� � b@r�4@tU$�- g!1��(��!p��s���D(��� �A��IFq9h�a�HC_�Z�	���uM�Y��h=5u��Nة���L��G���\U͹���"q�G�^��h�悪��Ɓ%�Ri�8bmI#nF�0Bp�Zl' �5"q�ϊ�(��+��H@RE����I�����
0�URDK�	 m�Ss��#E�Ze��i��G$�"���Qm�4 ��҂�� ����%SvQr]I���I���N��ɴQ"D�f4� K��,'_p
�H"�?J��U�X�_/��G���� ��s�/�����﯄��Κ� W�;k�T�<fd��i�p���/�ɺ<<�i���8I@�zO";�H݂��,�1��H}3 k�+�ɇ�ι��͝5��U?6��v4\C3�;�`1��ߨ�>�@i}9B��ۀ�|oz2�&����u��
_���#l@��O~���^<`�ǎ�0~ z�5W��������u�����	okk1�=�$�y���~�xOʊ�Ѫ#�RcY�A��a1qm���t���N���NUN�|�<��\��͂�1z�##��UPdb��� ��j��/f|6$no8�W�a���i��-�2��\y�]ǆ�lE���r�ܸ�٬3ٿKIL���}s�C���-�ն�E���nw�s5
�7���E�yѳ���]�X٩t5V0���3��P�m$���Σ�GUN4j!��9�}^���f� Kup�2��Ǟ1��dT��)�8����b��ޣ.VsI��hK»UԟZGտ����#�Q�^�m�P��k���%�L?z����e��4�u�w�	��J���6|}�.�����,;R��j��ngW{�"z�4<3�UY�X�\ֳ���L*�?s`���c^}�Wd���67q�q侜W>3��1�2Ұ�ٰ�x��*ʺ�ħ�Y���;Lf�Q�����;��w��	oѥ���R�U*��������K��x��}����Em?������U����!���'�o�k���'0a�C!d��'Bs��4��z%�2J
p8K0i�\��\�Lj�O챷&s&+���k��^8PѦ+��W�Y���|��5K��^�RT �wL�v���CJ��n!�--�6 ����� ��%�Q�����O3�cyK��=f�(�*�c��WU��`�%���y���`5�s�}�U�f�����&�݆�pZ���D@K�*=�hЪ����׋��z��	|g��U((���\jaCx S\�V�wVp��em ��n,r�TP�q���5�*�������6��F�d͵0��r���j�45�ū��f�6�Cy�|O�A�����Zs���>\�W���m��uZՁQ�̀,����PZ�����]T����ΞP��G>TFz�C�>������w)�����=�8|mx�x/�/蹊p$(���|����3I5E��485��G�z��7�����#'3sH��[��z@�K���`��g|��[���lX��B��
Ѥ</�������eS�Rq�/]C.�y��Żח\F�{6��"{<J)�H9թ}�\&���bd]�E�a	��Һ��	]�!�\��X�ᖒ�V�ч��O���jĥn�|��6��c�h��eVɅ2��Oq����Y���aV��LƧv\����Thhi��T�����}�~Z�$�a��#Zy�!R��ō�
ۏ	hpY�,ff�p4�*G"a�x=;^}��{Oȅ�C�$e$o�*g+�q�����4��թ�5t�~�9B��C�n�v����&�V>����&����4��f
A�����j+�ȩ~��
:�xU��9����NRg}�<G3޻����M����D�,��[H���0nk<�"��(�m�4C�fgB��]<��X�"⩎��_@�Am�0�aNN@�>F)�`5���c�U��l�Xk.�������s����%Rn�[u��fۥ���7!z��md�Q�Uμ1�~iF=~t �Ձ����+� /U�z1�O��An�ë���-��7��v�ud��0�O0��w����|�$��MN|�T��h�0��#B(qU����Я�E܌Ykz�����j���������9��k�Hq��9!���=:=]����|��ϵ[Yw��@j�9�l:q�cT��(t`6�������qX�����9ʹ�}S>���=z��^&�M����h�R%�ܪ�=E\̂�oɃ��q�O�;8��oM��>���e\�P�R�l���yַ��t3�{��aOg5ӄ0T���t�pr쵒�x;�#.��w��K2���������4���Р�C@�P	=��g��ϞL�x_�g����P�dcz�#s�%��}��1�#�T������Iߘ]&��C�=f�S����MX��v�z.�q���ؒ�a���{PSH8��2����N-�=4�])~���Y]�����j��K,�=F��X>�#��_�>2T6F�l
g�826x�\Q�,��ۻ�%�(Un�)K�%�``!��vY^xf��c� ��C��*;F�6;�z;�FPׁ�cB�Y��>\㺛Xǚ-�2���yW5D�`I�<&�g"�_?��Þ�fW� �ֲ]�����+`�W���V���s��b �H���ojcHt�@~}-	Y�ũs���O�=��t�M�N��V�v�ޏ+a��z�y���s�0�*�ŝ��GG�v���I^�=��*E�-��?L'ɱ����逓Ϯ�@*)�܆�W@ō��۶�q�-M��sx7(����I�ގ��W��\�[��>
i�Q��/�c�uOc�^������|)�����D����Z���$�u�i�𹀆@��C��)E0� �-��ʟ^(��0�t�Z���	�	��S�Y.LGUd	����1��o�h�t���L�Q�U��Bup��ܑ�u�~��z���Ԇ�J�/�:w~^L��8�K�Q!�P��<|1hrYS[붱�O>�gf�b4��8��.2��(��6�QL��՜����%�%k{��f����AM�F�B�U
hhQ�"�{ӓ+�i	$Mʭ�Uw��Z<�F���q3L�*�&G�H���,���@B��1V�-D��?�@��Uy<k
U��>׮9��hħX��-Z�MJv�14�a�^s��4����$�`�b���� �>����\���7���ڨ��X��v �.��s��y#���@��)����[S���?U��{�A鷟����jޓL������j�1E��)���%���})���H<�2��]ºt���y{Cs̏r6<4')�����7�Q�2�1�9v}u�8���A��ze�@�K���h�����Zސ���a�������I��V�Φ����*��}�Y���:ڍ]�Ԫ��Ѻ�M�(d�nj�Zٮ<ϩݧφC�V��&E�#NH���Y.�4hw���kh���i��0��%�ȟ@֩��_FS�"��z��/��3Zs!�mo)��w��ㅢ$C3�xĔ�\���<5?j���	�����¼�����:ZϠrza��9[�^��+�7K����K��5��=4��x=�h+033XjFq�P=>wQ>קy�K]g�9ēE�_������k�G]KYѯܫ�����grJ�z��ʎ5�z߭������K�{�F��|�2i���5��\�{�H'�"	����ؖ�u�̶2<H��{Z�g��)�q���7bd±\�F�M%��M�v�d���4"��(SCB����Y�߾�~��UZn���؋�Q|�1ށy�q�[0h&-�)�kSd��OJ��OO'/��0�H�����%��}OM�	E4�	��A��F2J�M�s��Qj������2	d�<�v��E�ǟ˼b�hsU��~TF��P��d�N �9�f���J2r%N9=r1y�qw�j^;����{gbO�rt�uő]�ꚔD�:�^Q�,>H���B�yy\7�2*��
0y��0��j�تs����؉��� �:��\��\��{U#��T�dYqr���~�6��!c����+ ����b_�{Ϭ�#!�zS
=r����JdptO7P*V8t��~v븋��6���2�K:�t�6���>�6��ǒ�kd_?�6��YF@,��N��v���Fb��=?%慒Ϟ�7�#o�-�O�b��
�\u��O�����$u���kQN9#)����a�ǡ۹Ƌg���4�B���Y�֞!��}��'�T�!Y�:П������#hS�*٧/1��#ߣ9����%K���Տ-<�j�`���Lg3���g9k6�0X��4ZV"��po��"�:f%� �>��unS����IQ��W��Q��pT�}�s|+�z�@
hi)��{Õq�D�5�E}᪔lP��}���7�G��� �;���¯�S���8X=9كGs�x���n�����`����z!�4��4�j�y����q�0�w8�;�}����_M<�G9�ыxq�_�G��KG��<$�n�*�y'	�-@�KC�;>9�pٍ�욦�W2�&�"$N��' ��������zq��ܴ�ÔSMu
�����W=������^�֨�;��#{��ҧc���n�F�|Q|�=��s�;�m]	T�qt��LS�u���N�;gP	Ó�xю��BcP���z~�����w���r����Ru#t+�� �n&�Ĭ�J͘���4!�>��
B*����c��k�������M5{j|��;�۟T7�ʵՍ�,]�[Q->%�T�D�g>�g5�?��s���mpE�)z] �V@3����Z5LS�[�I]c
*�9��Yy��ՙ��F��rbN�AW#(�[E���!(<��%�
J�7v	v��Ypb�n�v�WC��~���~ݖ��P����S2mcc���j��w-o=')ռ���4>ʙv���-��J�%u7J�.�Ȋ#�ŕ�����ܜ��< ���յz\�e�)�$.S��e�G_=�%N��5�n�n�A\�+yɼ�� �J44��Ђ5����y?t�/èY�U�&�r|�O��s!5�@|�+�W���)>��V�g6������4���R��X���zm4x˺}k���Օ�T&n��b�tMt�����7���[��Yum��h�]����Uδ�?�tc��t��X�g~�M����)�;�m9�f��ǜ���GN�D�M��{,�Z�\�
�(Q@r�m�Z��Pe�{����O����7n���zh��<�.��B^[��ms��Ǣ1��O����u�Z�Od8(� Ol�#������Vΰ~������	1�Cy@X���|U���ް�9�C��������e,)zm�勺��yݵ���;�@/e��R6Cl[1o|�k�}��4�>�.�U_瘌��7�^����|P���E������dFK�Tc3a��_Tx)ʞ�ǩ���<;{��!� ��~��(94������}�h*�ܲ=�ju8�&��UoMZ�	�xR$��ƀ�,�@ �
�������jb5��r��{2x}�J�#�.�|��Y���0�sX"p����ۡ����Zq�:�Mز��w�N.5;Fb��,�ې��B#M��'ݶjLy�I͊���ѻ�zU��ea��W���u����i�%��I�-�[��}ݔV�.j���*��A��h���JhiQ]��C�`��e��q���k�=�KFӂ##��gl��Q�QĊ1�E��(�/r�xF�l��v'C�L'ʽ�%�Tz��"���N�^�=���9bD	����Kם�|;�y�n:���?z�v�8�@�e����l�[��L��]P�p��^�ϻ�l~~�g�+;��L3���5�F�jj�b�׏�KQEխT-�nt2�/n��To5�:l>���:ȇb��q�)���o��Ta�纆�0=��&�[�Fnwӣ���1�a�f�������l|ڢ=na��z㙠_Hf׬�d�{s��)�zFƚdz�-1y V'��"=�!���Xw7(3��[��!�<�cZI������&�uQۣ/���7��W���`^��Ry��O�(�b;^��)��^�0�k�Ő
-�9{���nW.�/�v�D�ț2)��Ѽ�e�d�Q��7ϝ�G5bC�/~��p#��-{w���~�`��_<%�9/b���Pj����������_���g+�Ss*�9cI~$��b1��8r\��q��W�����I�N/Q��	����Ǯ	�Bퟢ��c��3����;���L���z�4��Cuh�:rO��m�Ċn�SטE��(Ѡ������F�s�b�f��.��ԥt�鵮�wx�gR禷4-�M�����b[6j��{���+3�����M ���x{�;(Cv�❮�~35��=:Ŭut�L�/u"k� }Kz-���P��=��-�rfNNb�3xB]~�����׫�x��"s��/���*�O�r�Z�UC1��m\��S4g��2��|o�o3�S���J�3S�:|�}U���jy2"�c�s�G���}QCw�٦&o>�h��i�%z�r̞x�,�T�&)�wG�=�n&rY�䛨QK�m{�(OL���Խ[�k���g坠j>�h^��F-��	�C��#�u\��v�����}~�\��d��|U2�A��u�o2/Mx�6��9cm{b1�ZaF֩�>D��p��B�%D�5�r&��Ȍ�l݀V�rqk�����́����c�D�)�3[z"l��s��g]�	��6�iQE�g��0Ʀ\,cfi�����v���ϓ��`L�O�:v碑Ǖ��?G�{�	s~&|Q[B���yB��2+8��8����L?ol�~�3̄Ibh��
���@7K�٬CL╏އ7�ދeϸ������[�8j|���{�{H��J�q���y�2r���\�D.�6���V�7�ߡ�'�v��N�M^E����>��7wYgjf�nt���=�A�3T#��st͔�_�w<�윀�e`l�'-r�-�yo�ܣ�|���o�:8�LZ�fN5$���Z�c�avV���[��V.Ꜳ*d�ͽFP�a�U��n�Nl����..4�1Ս[�����ݙ�*�����"6}Ơ���K�UI�1��͙���ս�N\v�*��zכ��7����%8y�I�q�iC�a�N9��ȥiV_��U_5��we��!t����2�����OUUV�zgMX��Xr8�T��G��N�*qoVѥh���n�˭�7��	�U�h�z��VW}.�|��?[�����]D4�uG�v�T�(O!F��a40���d�i�zc�¹���ޓgk����Vvb��I�iQ�%Y���/c|%�kݣ]>�eM�]ͭ
�v]	|�y�j*x���0f\�]�%��Fd�M԰�5w�3o�+oIһ�b��q�1��'S�{Pn�㢐{��r�6N�7[�`m���a��MLw��2��[à�x�� w4E�ie&���櫓�(:�0���z��$����g� ��k�4-6��nh�.��b��A�Ϸ�Twq��e�;@�}3�1
�.�엺e�]N���MJ�r�Zަm�b���Υrgh�G��<1u��:&B�/����`�tе����&�!�桜���a��(����C ��;v���@Q�k���ڹ (@ZM ,��u���H��n�wi�0X$����1o�9��;�#���-�;�8�{Dމᇚ��η�3�)�������N��i{wt���ڤ�bRs��C��wW硩j�3�=�$yQQqt����.�'�����#�Z��v���73���dW�])ƸU�4�f�e��L�c�zw(Q��������®$�5��;��r�u�,���4���I�@�ӽ�+gQ�#5;#;OnZ�A�X}w�V��35�E����.�$݇��hK�=R���ʛ1�U�pq!H�Ol?V;ɸTnՇ��F K�}"�n���{E�Ր�����.��n�Dl��8}�i�So+^u^�����/_[��t�a;�]wlGW2���GS��/�_
ɉi7y����;i��g+�{��O��
6h0�F�l�dW�;zwT��ׯ�Ϲv���#K'
"��w���[�U�Z�i�4<Vjc}X��>���-��@]�ٝ�W�Wb����³�+�"X�L�yH��G��j$��;J]Ǥix{+�=��%LEU��*:���S��;�Q	���,]� o"�M��-�i�n+ﲇ\�ѧ� �wݳ�X�ճ�>�ܓd���s��+{��|��"H0���ȱE���52ŲW-�꿛�׎�];x���qǯ�8�o��ݻn⺅Cp��Ũ��j�@bDJ��>>�����8��q��8���n�.���"L�Q��~6�ʕx�޵�~o�o�^���8��q��8���{��xѷֶ���+M�;����*6Mx�5���|[x�oٹ�Gw��s�z׏m5�u}j�xB��\�-�^^u��+�^���VƜ�˖?����x�r�-x���X�\����ŹF�ws�����ur�4�}�<���Z�h�������w�X�������w_�h��U�/���ݨ�R#���5��d���H]Qk��r��D]`��O�{�}�PLU���j#�"mY`�ژ�������Wwz��f���ďѠJhiR����s[������3����2n��!�L�� ��1�d�zg��ҥ�4�WL&bxf�7b��͡'̳�N��$=
���ͼ��)��ѱ�c���
+���vk1A��і��;UT�n�!�����$�Zr%�$��u�'��b�z	������3ݞ�׹9q�+��Sۡ�98Ġ���{�%� N�� <:B�In���U�3��ԻC��ǩ݋ȗ�+A�ty���ݞշ�Y��Z]Q�B��z�q��#~tt��{��h���C���ϣ�6����m^� u�LKs(1�!�B���|V(�4EL�G�A�u��0��/-���J�x�CÛD�O��³�@0�N(����1�Q�-@�KCʋhF�tQn]ݪ[GE�V.��k�ô%|��$��*��fR5�9a�~^8;�&��6�|�h=�˃�`��M��-T?<�����,�׽��s<#i�����(�O��hɘt�:����Ь1@܌]�z4F����@�q�W��;���+�q��z�v��2,)��c.�[�voD��e��̖�SY�h�[����~m�^!�؍u2�U%R��TN���dս�ִƇ	'R"��<a@D�~�W��9y���{��+Ԓ�䠦��=W�֩���/u��c�n'�[rv�3\���2�g��k�?
����
hi�p<�;���k
�/~{P�h��C��>�%Y�|y���MA��۳f��6��r1�˸=	m6�e��zB>ƁѳMVa��/�Y.c{J��Y�j!�ݙs�w�{���3owv�ch��lg>���G����>/��}9��"Fe�r�S��������ڑ�}1�ԥ^������w֏q�2T�Ǧb�X��>�1j��>^aKjSw`J���r:^Eq�����|#�@��0�T55VX���м{Hx���!�T�qC�qxak@�:����[Y��L��^:���,��Ƽ5�P�6�x�1	��z^��aG7��-tp]�f�K���ߙg7�Qm��԰>����xF����A�v�cGv�o���׸��R�"Z@�`M&��ᐢ��^s�������`hhu�3C��!����<�j�<C<��ydϊ%���m�ok��Y�3W��9h�I�}���~���2:�i{4�a��۴�B/R�؞��>צ7ͬ���t��˞���������3�?%@���i܂���J*�՛�>�Ҳ�J%�&�.�s7-�[o;E/���^���'w�����U�5b+ ���+9�9���^ք���\��G@w��Y����ʵ��A���;�4.����s��o+�����W���ҥ44�M�|��W�T��]BYmk�KW���P����M6�h9!�jM7�D��0�|i��f�ff�Ϭ?!�$(���|c>�#F������Ʃԕ�:�c�u\��^k�E߇���`��GRF��'�ᆙ\�W��*2]���tJ�vAq;t����f�ب:7��� sd��N�C��ʇ>P��Q�*�3'��JےI-��1�d�m/[�-���u��2�2�IV�Q�t�;6�u�=��Bo���wd��j�:��z�b�f
��H�n񋡊m��Q8��]�b�g)�$���vg^d��=�U�QF��6�q�Yx:�Q�M�u03^��ISmA�nh��b����M�ⲅ&�-˞��|�ǯ���i�j��(Vn��w�Z}���6�ӚI>נ��?&'�r�%?*���Ͱ����!-�i�ǳo���}������Q��> h3ʈ�˵y��r�}|�+����b�V�n9a15\��	��%q�͵�*�s��|;���
�_i4�κf��3)���<]U���/	�����s�A����H��G(l�`�B�wH�|ahgNpq_Y����.�����Q�q�`�)o�b���\���q�%TB�K�c�S��/�k߯�غ�\J�K�lK�(e��l�m�5
M;n���'f`�[���I�ڴQ��m*���=:�;�B4ov�܇N��S����@:T}{~��i�4��Ҵ��A�|;}Ϟ��T��'�-5�]�Z3�j�(�`/Q�lֺs�v��@#dQ�ލ��[����{��:,=��(����`z-��'�E��[s��;rS&����`s>�,h��?e�5�'�){�ݨ�1sޕn�C�h�h,%I�: =S�@�2*�O0ʾ>�hOcO������Q��^th�����Q|���*+ ��a^��3��W�9}~��|i|9��.e�2�~�φ{�,�L=�QӼ��hXH�et����)!տP��I�:�jĜ��ړ�+���b���+~/��m�&i�}]_s=G�#�z���^�>�+>+����M�	�D��W+�*�f�+�(�5�>�0,4�*���)�={�]�Px����֔b�i�Դgv����<㳛��^�7��8g��W�,�f�R�3}�=�L�2�p&��!�,v��܅:�6k��_e�[]8̳.юY�=�9��"X]|3|�<�}\׳(��]ܘ�p��S�m���U7{lT[JR���-h?5M��~�~���2�	�;��r�%�Ǹ�K��T��rv�2�f���z�GVE_�j���b������;vd��F3+F�UYU��y7��Yη���.6����p��u��ݮ��\�n����s	�w�6����s����q��8�y��3�`�zV����b��3�e��Mj�+���V�p���<�y�R1ݱ�G$�ja�"]vq��':�J):�r0��qG�0���p{c�Om�C�p�p1Ǆܻeb�cL�`� �(R$lAO��4=^(�]b��Z��Ed�=[㸖kpz�?
0��Rg,$�/8���Lf�ph��':���&)�?`J}��H千s�I<�Jcq��/b�׸g��!L��߆�����Zx�C߸>��r�L�i�|�ɩ������cT�{}[�v����E���]��n���0(i��*	8�ǵ�ywW{��.�x�\h�j��Oy��b�ƽ����Ҷ��0�v-������[0O�go�@���n�;~�	�G��^��[���stTn�.LX��q�䤰�M>�"u�X��I��ɵ�#�w��s�qGO:��<�Z]E7��M@�u�,V0A�7�`��}�h�'�CJ�A8/F/tT��~���oq�Y��e �ް�nk�ɘi��q#z -u�y�����D�uvHvr�Ph���v���V LR��P+���pa�Y�n��C�l9�զ*�:�`a��g�	��V]M���?�<@�����:+��T.HQ���*��Hc{k��sk2x�xBzkaim�q�²��W��_s~O9E�����MM
7=I+��|�,�#��O��cO	$<?��)��׌�y���(Ǫ�Z��*[%�P�.�'{lERht����G�"$I>�w�S�;c���v_6 ���-��#�q�."C;��8���@�gҊ����js)�z����_���aȊ��R���U�w때�B��-7�f��(��:�q.8sJ�x��\�i���'����f�6�Ly!���8�L��o���y�jr8�Mvx�9d,,�/}K���u)&p����MJy��� �;�;�&���j����J-���b��Cͻ6��S�ێT�*k4޺�����8M��^n�x��X�S,���i�%��/�7]ڈL�s�5m�����&;��1!��,\x�v���:O��o�L.�pJ�[�y����Mrr�yvd)l^�8w�;j��_A�;2���мw9lx��cL�p�����T��kW����Z:��R~k��T+~n���@���i�O�\�L�wyZ
�9�����|����\�zT�x�b�E�9h6���ɒ��KZ�>�]�ܹt�מz֎�q̫����x���h�#b1�d�5��m��G�w���It徇��U'>97�Rےޛ��PY&�/���ki�s���6n'�Y��-���o?%�8����}�i�0�B�H��w�v�΁$u4�p�����dEĒd���Zi�,�a��������ڈ�Z]H�~A�z	�� ���|������ֽ��۴�;m��*k3܆c�M@Z�Ʈ��ܲ[S��I<=Ӑek��:�"r�}���x[��t���w���'-�q�4Նe�օf|�8'�kW����0���bNX���3�P�oI���}R��-9��*z�I��Un�C�������@FQ��;�7� �j�gt���ٰk�>k��0*B�/C��a^��\[K Ć�qo���s9�u�;#)L�.�W:�7�p&N3�|�7�V)z�b'(��ee=솙e4Ӛ�p^�}#�8�n�4No�%����W5D�IG(z�:m5D8�ܫ�y���6�Z�W5ُw��d;A�"F�!�2�1����Mӧ�;6�u�m1����l�])h��x�)���!0;���|�S�Jg	��3����R��񨖽W.ÖżJ��4����^���+�����^t����w"����箢|�
�zq��ii�,H����y�m�=^����ug99��R9��Ƴp�y.a��]Ԃݞ�p�V��-̢�=]�S�w���*Ҋy�O]��F>� o��}b��)S��n���QN���:�\ot��-t������.!kihݸ�I�ݗ�uU�=~�45M =�9��=���k����g?u��^� 2��	ֽ�W�Ǎc���ކ9c�����!|e�t�D��:`Kb���X+f��]h���LS[:P0[��E(�.2�6:)����l���C{`�p�g$��P���*�j��{^�d����=��*}~s��ۆ�c(ݤ,��Ff��r���:ծ9�1I�q*ԍ����h��"�=�Z���l1x1�����q�&�vֺ���\`oL-s<��������]��fqmŪ������bo�ܪ��}~yg�y�G<9��M�rD��(�s�<���ɯ���c��|���Lq����Ŝs4K6ù�p@Km��E����� QA�]�'H��}�B)��+�����]���ȭ{gO2z�����D�S�jT��5K��N&���(�P}妄C=�T���c ؍dӵ�T�&�W��KR���u������U���ăD�fnӯ$N�S�y��V�s���'yע�H¼'�Y��ݴ&���"��|D8#�C��_N��!��]���9��ޅ�p'������d����wX�S�w���|�^�W�ˎN���u�Cr{*j�y�2�3��#Khl�\=� A㼵9Kch�+t�w���Ժ�cqɟI�-����^24��h�g�L�W�:��E�̂p2qW'Q�~�hh)���3������������+�ȸf��g؞�5�����%RZ�����Z�[�݈�%�M̼��qd1�W��OO��;?|�`\���T��L��1z��><����R+��ND����7�^�o��w�Β�5�6�
�{��s�j�������;@�1��e�cc�2����	�?%Ӯ�<��ă0���*EW�,�q�R�O4���l�7RuY�!l�&�gP�������o���PKϦ�܉����>Z<�>�%�0�J
x*�@��Ut���T!�����6c�Y�.������w8���vn�y���Q�4�{�X�r��u��l�Q�|X�P�,���*�MC�"v��,a5�>K<6��ҭ���NKз�z`����/���3il��,� ���-��O8fĠ���rz'��:��n��U���ѹn��[9�����c�*/���q��&87k׋���!��e0��Hfl�`�9�\��[�M\��VE#�7/o������� ]u����cǺ��S��p�Wy���M�x�x]�Pv8��m�8�a|���n����̙�CMBona�a���U9����vCY����ip���#6�&^)@sY�����:��s��l�J��i�z;:�X��oG;P�ѩeZ�P��!�^g;��ge�J�c�c�hi�;U�Wԗ3��a��X�����M�����ad��Z]B�o�-�|��׮t��i���U�\^>EGs���IoR�:ŉ߻UWM|�V�O�{�6��'���S3�{�$�(��|���E��Ǘ����3ёB�����1LX��g��#��#eR�<�=���AƷ�0R5��z]3�����⽽���|d��Нa�~�3������^hW���M��g�/d���Uȏ��XO���z��DS^���׷�c5�6v��ڂ`�SnS�����QR��x{=~�j�t;����HrzW3�,U?����E�V��=>����h���dn��7x�.���/�q�A{(���"7��/r-�z�D�W�b���\���q<d�6�[�5]UMYu�A�}�]+x��_A����}) ���t��H��3g�ļh���e/��׻_}t��G���<=,��g�zqM�m��H%�>��v�j���/u�j�����9)U��BZ�s^:[�C���f5�@�Y>-��KM�m��4�b�oiThS�ʈt=�++yL���m��5e���[Nˑё=�m$Ȁ��BCgI�_���G��R���.m��ᣙQ0S0݇�Ad���i�y����Ӡ�*�[����KE��+a��<n�=�N�e�P�n�aY�Z��+p�L�x�Ϙ�ʭ������s�κ�M#;7���)_^��is-�*�8ʲ��C�^i�$ŀ}S��u��O(o��u�vZ�%��Z&�O2����^q���|������yt�`�WX;x��Y��W'�\�y�6��ŗw�	����(m˼�I�o����շ�{Z��j�W�Z�p�G�E1l@��Ol;����\��}�q��c왚�t�e$�;�E�v�����QEi޻R�,���'���m8u�����;�qu�b��	Vo(���_LklV3)XVd���G�0�Un]����α�,2��޾�c�IRƦ+��ֹm�y[�!e;���N#����Y7!�Q���F+�������;�������l3��(<M��':t��0Y��o1���iU%�ں����bþ+Bel�-	c2	K{��V7���uUm��u���],#��rO'���NЙ�i���2Jy呆#��΢x����&�*
�-Ԏ[�O}!��}����rl<��Z[�4��a���չ����5��N����dh+�0\F�#����;L����\���z�P��#ZjV��˳����
�m$��yR� Y��;f�'�!�f''�keU�ucSD$W5��k�n�V��-M]|�w)������L�T����K���X�=�d�+(v\�y/��5sP��.f��Y�������H��;{.��׈�@�Q\��d{wCT�}C�]Eŧ�}bL��v`��֩�w�`����Ӈ.�6���*Hdc�!5%hYsE�nN� (:><��vMɒ�ުG����N�ν���e�On]O���8$Q͹��pi���;��]I]z�۫�vfd��nMU%��P9bзoh��vjXӿZx�k���O_]����K��gF�{}ņ!�MU��"�b��7���?�.�G�|/�;ܪ*T�j�����_7��MZ��!���ut(wc0��侑�y��b�٠Sػ+M۝6�w!rE�<�3s&2�F�`l1'+�{]/&��ﻆ�J���&�5�A�j�'Kz�!U>�'f����9M�kcK�p�)6�T,U7i���Ǯɒ����"�f�F���Ү��je��SWi���d�����:ܩ7��^�rc �󯕼ig;����k����ͬ�9��YUw��'U�n��z.4[��&��]�ѝϹ��k6���r}���R]��L1�T���8�<�<D H��W#��J+�ݳ޹N�Մ�'h�n�<q��\q�qǯ_�8��ݴU��$�eQQI*$�9�T���j�:�������=q�|q��}qƟ\v�䝪5ET�l�DnLj4E�U��!*�HjL��6��׍<z�8��=z��>���v�ʉR�Q
e�k��O;��'��?��>wx�Uݮ�Ə+�ywuqr�����x�����|A(��ơM"�)4�m��<�G�$b��^7��:h�z����ӫ��Ǿ�r�ϽWdk޺|�]79����\�߾\���Zr���{�����.��ys��|��}��z��ݻ��tם������P"O|�z޲�?��s���lǫ����y|������ /U׽�7Ν��x����μ��Q��K�k��!ZE�&��+�`�L�
R>DBP����H����$> �	B��D�ɦ�a&����6�{�.�aU�T��� ���S|&XYe��l� "U��ɱ���R׀�7(�F�����ε��)��L	p�d6�@�L��%�!1��.Hو����L��S�0��l������1�dQ��I�Q��RH"nAID`I�H�K"�O���Aq ������\��&E֧��V(cB�)�qd��BF�l'0��>%qBw���	;�`��}�3%�X��1Okc-��5�d���%�t�X��"�[/w0�9��;��n�?��E���+[B��"����*�]v�r͞똕ly�۫�gkI�m���4���ޜ�X������n�hꉬڼ��˺�	:.�}�[h��\���i�O0�c��`}����oǋ�����'�a�ڙV2�����F6���4�E����}k;�7��zJ-���;��ȉ
5���R�N���G� -���c�S,dY�- Wl�Wd

~nY�00�݌sijjv��BwX�F�z�G��ΚO/���I�J�{~~9�F�k��<gZc���5�4lE�]�ZZ^	�76�L�h!@t'�_}oK8�F��|���Lov';�k�~����<R.%����U�t�R�z��m��	��HQ��|c�<4��^�jO��9'�1�'���8�3��(#�#_bd���A@ϭiȇ�y���u�z��Aw��g��9�C{�>��\�\�O?9���:1�~Y���������63Ə��l��ܜ�QvI��T��+:�t+�v�<_��u�)��Slb��x�{o����	�v��a����K<�n�]lA�&�K#m<��Us�n��<�a�� 6jq����,щ�uk��P�ߪy��)ɥ��G
�L��׼Ƒ���>WC���=�}�Tky^�sH��L4��#�@3�5�S@{ ��O�ͨ�Y�����9�e^��=G�C�={���B�?mx���ײX��g+L���$j�v7}h�4?���N���4�Z�]����FXF4�R.V1�C�1r�}��Cg��ߴ_8|n�#]�"��[�v�)��m��*��!᧐>��Q}p�pO!�-��C�b�?�C��v���oo�u���Rs~;"�h�5�����x��q��8�5�AR&߁N��]�g�e�s�z)�!I*)(��l�El�qY&V���Ҙ��^ׯkkW,��T_�G�|�l0���V��pQff.�@�י��v!>6������@�מ�n��S������fg�c���׻ ���F{3�]6t��'a������ɝ�!]��|�f�J�8ǒ辘��r�*pwI4�>�.]��RF���>�=?*��kǽ��NY�
9q~ʄɸ��������өڪ/�9�����=w�1S����V��Q�&�k*�B^e����	�֐xրxo�̆|9��h���Y6�v;\8��k6�[%�㉽<�3�uvʩV'44�����U�JU \��.�뵳�z`0!��7�{��=���V�{��G+Y��Z��#��s\3���E-7zC�I��������
bv���>e���~��[��9�5K�/�b�XK�B�%9k��:�j��zN�QȂ}�#�x���AQ��_���z��^�����u�ݚ�}.�>}R�3���AK�X';ʡ�xǒ�gP�>~|���0�P�����<D���Wz���Q�w�VY;?mE7�\��kuc{͜�W�TM@�q�&�"�v����x���@�QM�7"Jt��`J��?E3�h#-1*m�m,z��!�s@}����q�ߕ���|��P�-'�>��͜s����p���콞���q�w�^����ԟ&�u�����f[���~v�������Լ�¹��n�gxzr�Jq�M���G��	@�JxK�y�DV�)���F}7s�r������?Z�ʂV}b���	n]���e��6�>������&���-�5��MT��k���A8���ֶ��{��
OKP�	Nc��ŷ+v1���7�푌W������D@V�ӂ�wA܋}����̝p�)�˼�]�])�h�Z�E�����S�k+=.N�� �>�Ve<���Zke�F[�t��ūN�ؙܤ�,`���x,��ȹ�R�6{y��@�3F����o~C��o0��T7�IO+o�ָ-��b���SB���)�~!j��f�]@������4x#Z-����鹳��!��w|��t[�`�
��[1�蘦\��%>��r8�.C�e]��fl9�$HT�0��@��(��'{�������@(�ω,�A�^BpE��ИguIn.�!e�Ye��l��'��1��6X�9+??46F�Z����~�
��pF<~�@b�S��A=���LI���u���t�=Ǔ��_����vi~�E���D>���:7��gVz��>j�^��Zd�v9O�� ���u�3w8��3�n�t��/ʔ~���^/H�S,�pN׏�l�lL�dӤ���zMc�C���b��}:]dv|[&!�Z�sLS׀��4y�98�ޒ�`�{y�Գfo]"��:�~1٧cѡC_��	ި��?y�s�>Y̦|�³���5�ǁ������D�K������f\����hy׆s�b#�����caq�=�[��̗g���a�SR�j�dgw]���QwNS�u�uZC�]�Edd���/8R�зr�xV�F�V
�5p����mG-��K���r���U΢r��!����;wb�U.�cBV\��l���xj㜲eg9�:�Ç�p��ul�
m�Th�P����fs_A�9d8�(��E8c����P�_g� �K ��(�����&rzD}���N���c�]���ܜx��~�н�&���8h�t ʽ�XǾv�O���tD���8��apfz��)�.�(��K�&�}SO���>�i�'L��uc�Vؾ|9�'ݷ/\QJϔ�n���b:��������>�����N$�r�1��ac�ҍ�1}�,�Sm�ҳ,Y�ʹ�)�E���ooV窗�Ȟ$��h\���{s���1��W� �a�,�4��=b^�O�[W+�aG�# U�:��p�MH� &Ƒo���kdM�<����Q��f�4�_ zYN>�CUJmF%��["Nz��^�B�@U�n������v���W�a�T�㫴�0��:�4q����x���O�S�o+��l�����b�]�1hWC�m��" 8��e�� HX$����I�j��g��*�=��e�bF��?��w,x9񬖩����*�����U;�!ְ�ưwtڲ�X�fD����ƙ�4�e3
�m;�R2�3�����$/�wJ���0ݩ�q��s���]�d;��r���v_G��m�����z��a�^I�و��ɟ(ڤE+�p�!󂶒�����s�S0@�bӦ���]�*�䭕&}*ͅ�F�A�Jz�rvn������^a�z��c4��9�P�Լ�MM2��yÙ��e�9��ߐ�JU��SoT�͌��z�;ک��5ȑC�f�Ť!5�,��U��V +� �#�S�ј�[<V͖}��{�ש�Ւ(z��}�
Zk����G??��g�b�SS����k�{���حܽ��������A�zD���-"(�Xha���u� 2���4JI*gS4ձ|��]L$�ܤe���3�o��1!��)���7.�9�ע[Y�n.	��wƼˉ��������^�Û���z��7y�am��cX{5.��)Lp��-4��i_O�1�`�����ɉ��<�4��J|�)��}�����yH	�=0}O�	X)���]��a�j��|N����B�-��^<y���s���$7��Я������2~cz�0zԎ�yR��?)9T�a�T1NBf@��5f��ŀ��+�x���
�T��=;�J;�<�)�7���v:���["�J�����ݖ�y��v�)�I=�z��5�
y�P-�'VG+U������4%=V��>0l�a��{r���5�~�_�n9U)�邏2��bO_a�V팩�}���vq螢�M�J}%Ϻ^q�$;�`w��'���mڸ�z�o0�y��.]�2��4P�BP��t�Z���S��B�V0��q�ѡ��;��c�5<�t�m�Ȋ���2uW ?;=�хN����/�b��#[�H���l�7T�uf�Y������B]H�6<�����'z�<��ǒ�ʧ�U<��i4�ZL^��u���;�Xs5�6�<2n5���>�KV>���L�E��}��^_��j��?a�x'����=H#�����������˼���a�����f�u*b��X�A�o}%�[>���ؓ_p&���0�a%��k���|`o�fJdwZhfOQQw=;�k�s�.��#rq�L��[U���@�kH�Ũ"��(��������uz�e�ԮJ��u ��|����125����ſA���+�d�/#�Y��(^v�v�<�V��?b��Μ�܇M�p�e�dy��`47�`ҕIi|e�v�l��׼���u{�Q-�1��́���!5~W
�D�;ky����ԾW�+�H'^���A�mOua�>yO?V=߫WO\�7*sv�v����)Ʀa��3�OFk�p=��u��^�e�V�Ӳ91" )7t����Yۼ�B�f�'J�VQ�9�n��pZ8)]OV^!(D�w���û� ���<a��v���L51�d��iΛw\�m1��� �*�����!��������<�,k��WG+���b���D�W��I?y�A��}���@�Ug��k�nچ�1Xj����c�t��?�
� 3�%qm#��1�����[�u�)��M`�h��vn�[�͟^���<k�����̌y��ZU���t-�̤k�kj�Lu�S��}�:]��Y0�E�����aяŔW���"�&H������;�!ҿ@����-�``؄�8Ǌ�ݯ�fP:���&8�/n�Ŭ��.�X�=���N5z6��bl�f�Pu���&)�?:ǈV'T��ջ�Ⱃ�ۆ�,jnտO��N%gܔ���Vs��ݓA���7��dE�4�wu-W�x�c��c����n��>*N8t��Zmهp��ٳ7K�<���a�ϼڇR	�q%Z�a|L�G<�L�S�[kQ}wv�63Pe�S����&��[�"}���7}�)��������>`-ts�ε���6��쇈�i�^.L ��_�*��}ĹX�/-aI��4�ge㠕X�6�8u#3r��Ŋ;��q��6?z�b��F�}�����"�'�4����.%��#Si_6L��Y�b���.ʫK:�������v���:�e"��uu,E]7`[[���|���<#���x�)I8SR2�k_L��כ	g��16�H"�!��l6�D��d�i�Yr"8 ��	1w��<�_}Oϰ[�eH�	�����!��T9����3�zy{��g�:�A�ʆ_���~]7���(>+�Ox�M"�l��5Ͱ�����`[a�qع���
��`l�m����Q'c�>ug�� ����$(޸��R����=�i�	$xxH%�S���K�ixo�ai�@Rj �KC���1����Z�G[�oc���Wju�f.%�y���s`�̼������(Z�X���Y��:���wg��0/���n��t�g;e�w;U'�at!��P�ه��_�����~��C��Tq�S��s��7r�Z���73��(ipZ�TSJ}��#���ƤM�{V4����Pj�c�������DAܱi����3+�o�\I~~�s�3�~S�n2V�c{wwl�R��3|�c_�na����)�P< ���xO�#j�?uxk!�"l�G|�G���+���1����h�~Hv�7g�=T���hjA�aEFd�
�וq����c��}����)Xύysr)���~��bޫw��J!0��G���i�ؒ������J�,Wu�l�A������Q 򃥎�Χ1���[��-����	Yz�S�����vnoS���^	1n%oL�}���r�9S(��v����<�a���3���nv\��kQ�oc��M7R�l��l��QqA����?M��]O�����2��Vo:����&8��_��'�)���R���y�_>�p����n`�ە����{C�>��X3���� ��|��xe>��7��4"����ߙg���=71mwxC%�e&�\)�4�Ά?��C�	�D&ޘ�KD��2�Qk-QEG7-��$,�O/�m�g�
n��1mI�͏X�'�|�}6�p�^6"��f�lg�6Wd�B�'z)��ilsky�י�L��1�A�Z�6:Mk
���G���W='�F���{h���Ϫ3wLt����*Q�F����o��G�����r��B��Ў&��|�"�h��Py���t��$���6]�.��%#�1�a��>����b�����t"u�o�	����n�Dr�wg�~������	q��V;6��b��4w�)�qO�.D�0��w���l����=ˈp<1�����X���y��py��켜���J�A�/�����,אּ� �U���jmW�߶v���j�dh��ԏ]��0f��ͧ��٪,�,�n��25.�;�z�-�p��t�c�pvw��鰷%eX�}Ar�{]r2��0em��[ˮE(wب�|�2^^�u_>�ٜ�Q�xw��c��ۜ ����r� ��;�����,>�m�zq�i��l�?�n���U�mZK�CVL������ͣ�lM-d��̈́X]�{j��ш�����e�\ޙ ���LN3���2������t���;/ ޶��nes�\"Y�+�lZ�Ik�!�Mӗ�;Ǌ/.�]�3��0=vʑ��O�2���E��uz�Һ�!��s�]Y�5�U�wݻa;�c8��]�\y�ꎞm����̐��"��i�����K�5`PL���ƪ�������a���v�rێ����/B�.�~=���YsBԥ֛m��E�pY&��%�af��~���P;�^�2�m�}e���;;�iWgB���0e%zE��ḁ��"��ŧ����mΆ�����˩����Շ�:�v.��bN2�{�b�M*�ʮki^��X"�J0�������ͷ5��n���pt4o��h�Fk#wn˪��&�p�}��M98����w:�,pv�o-����n��md���aJ�W2���Q�����8˖��d\��	��40����v�Î��e �a�dt�]���)3F�2�"�Z�s%�	����J۠̓Q���!`�[:��02�i�q���?\C����yZ鸽H0ޅ�՚.�:����]k�܄�o`�;`���<x��ѽ�)(m��fU�8�]�)�}G~4h(�L���VNi��j��o����483ݧ/�o9*��W/�_��]�U��$�	�c���Cj��WXF�I5���q�S�шW:�H)h[a��̭��Jf;�����LGwr�Z�M�y+Mi���b��م�%�L�e��%1/!d��iB���h��w.��X��oI��v��b�\��Ձ��o-��Y��gp�9�3	���� +ag�<�W��O��P�aY��K_�,���\l�J����1��b���+�@1�җAߕ1/J���N㓰o9�m3]�L��� ���:M�ܸ7�Ry�luɢ���u�W#,%�m�;���g�-')P����әS/���3{e�h��f�A�6�c���z��-ŉ��*&-9O�So+*ڒf��!�:�Q�S�k�J*��4B��s'4�Vlj��8���0��>�f^2�ry�����;"Ʃ&��.ԩ�Jk�5�D��B�fwW���%f��s<��.��J��q��Ȼ}Ϻt�ʷ��Z=��	�)6�������(�;�vc}s.�]V�ð��;k%BG����i���q��z���}q۶��I���HƯZ�y2x��~��|k��u,�@���BBjR����Ǐ�<z�8�z���}z��w$ �%��.7T8.�(*	.\��j2�c���>���8��q�ׯ�1��mVj�D����,����������j�c����wO9wbܹbO�{���מW`M��F󮼗C`�t�WCg�����|��t]�o�]1yۧ�yݼ�i�M����A2�/{tLy�7���wv��#7�����W.�%�w/�[�^v�v��wu��/W`z��ћ������Iwv_��;���yw�]y�<��07wf��O9ܗ]�K�y�m����|n�y9�狆�(��o|ݛ�t/{�/\�
A� �H.�@�xAD�uO�i����FcT�P�z�i�,J�ʽ�3yK��z -=��cqvn�W���^#���^���.����o���Q�ߺ�˫��P����gzH;G�V �G�� ��W5$ݚ:��|Tܫ��݆�I���(���AtAF�>��"Bzl�5r3j97 �<�[z�`mi�ŵ+�K6r'��l�����!���1�'Yi�?j��L}y���'�=�(r�X�s혣�����1���Vk�y���V���|[�eL��056O��N���2&Yg/��^�פ`�=�)�z* M���Sl1�����^�dy�v�(��q�8�O]L�3539�O~�%�3�3m%:۞qĩw��| jT9���-���Rw���]Z��p/�4cϦ��>L��݈���6?j����i��fOst�뉵��rY~<ѽ���'kHF���=_�mW�]����@���ѽ@G4Q�͵ۙIos��8|7�>�/���8�f$k`k#��+Р��6=�K��Mq�����h�,�0yt&���Za���~z����i���4#��߰c9���3k㽫 í�˾�͙����\LU�b6��h�ٕ^�׏��]fm�lt"6D�(b"f4f�	LN���˳�D���m�+�4u�7�;u������Z.EW�+`����l�8�]W҂�,���>OX����L��
�|�u��!�g�߼���<�oz���5˓���EFo��������,��X���+Ѽݴ���-@�֏;�X����"�ᪧ���N���9!�+~��V�c6u�>ރ`?����C�0듺�^ΰ���B���`iH?3�����+�p@�?O��hS��22���\Xn�9��Qۜl�c]��:�gOA<��S�y��^ȝ��|����$�hD������w63���]�
ًא�x�i���H�%��������<~� IU�D�u�olL�0�vv͙~����3/c�w`=�W'A����j6�ݗ�lP��׺�b���^��p-a���gd���[�\�OL/Z�Be�ǡ2��W��N"�����H�9����׍��8��혷���z�k�`��q����pz�I���R���v]���b��/g�3��O�������1�vc}NhQl[F�H�o:O|c�jl^=�<������G���cƠ��c�;��\L���cE�Az�/���{䷪� �F}W(g���:���|E�f�v����c�)���M�S���,�ږ' 굽�u��س٬X���;cf��Mi��[�rլnc}�ڱ�r��U˂���_#j���x��ipO!�i��ξ3�銙�j���fe��~`�u/	U*n�F�,;�]�}�Ė�Xh$F��0���(�B�BB`i�����}���/~퍸סּ�>�j�x���h/�4'�&C�Ost--w8Ʈ&/�-c����I�|�Sv��Ҡۅ
9��E�f�a�t���p�y��n�Ц��u�4��u���8�6��YFd����	[��<���ٯ��]�qw7J��Kw���c$��"#S�ʅP�U�Ō���
���k]kX.��1E�_��9�.����C�B�L+���a�yc1����U�OTc՜�����p�fU�t�=;���Qح�ca�A�JO�a_w�0znS�O�����{z])Y]��K��Y�Pֱ��Tk�,���5��<���?)#cЗn�a�όt(�/�e��!�&�S$k+"F'�����L�C� <3���FDH�8\W� ��dn��,7��춷��̛�	�V���L�<z�?�Vr�uR;����,{�+�s�����NV��UU;U-b�hH�yp"_6�e@�W��([HnjmNC�}����"/�ڈ��G�E��Uq��{q���\�ii���Wy�ԙsw8`/��^=��Q:�%���[L	��\ZaѸs ��ti���r��_�/PLk�PX܇z�-4o,�cU2I�Z�m�m�Z���r�Ѣ�ip��cm����z�Cy{������²c������ ��Կ�r��pZf��ҁ�\X^�=��{�M6�d�ʒ��z��L���ٖ�}}��&�����;(��K5Ƅ5��8y��zz����f�}�;�H=��r��o�N��e[{8�Фg{m�V|ԥi0,5� .�ǋ�{� ���h�FbN�n���#	$����^F��{L�m�oN0)����r5n��TA��Z�7�w+>������U�F K�~h.Xq�-�N���F+��F6Cɘ�""�&.)!´���L�`�;��"9@{T�y�{�qzs�ZҎn�0�9�=�5��*�Gy�m{�>�]���\ ��M}���z����;B}4��/}�CJ�];�,�7�Qm>�=@�seC����M��q
�ע�d�x,�0f-��2�"�2g`�
j���n��	�%݊z�g��~/��^����R��Mt2�@'^��Z����ʹ��B(z`y��s<�rz�B�t��q�w����M~�}>�`�a�$��Ϊ�8Z�a?�W�z!����DW�
��#�3���\^ݨ)R(X���5�%	dk*���`佱1�QqK����n�"��֛k!�ݪE�rA���G,1����'�h�˞�
��(S=�e���Z�����u��/���g2��n+��a�����%�쩆�y��s=��U��7�	۫�XZ��/:�A��)��oXG��S��P���#��N3||��E����c���ۭ��5�����-���::��pŵߗ{�^����Tҙݐ�R|��S����g9\'�G�k7�??�"s�'iD����B���,O)�|k��r�7����m��w=P�f��ҳ�I���u ̟?���߯'4�w�dȝPC*e�c3�y3������*hA���g��A�Y	���.�
��@в�{��+�ĨF���3���@k�ֻ�P�HgD��ץl���Nbc�q=���+�#fº�~���'��g��Cv����]�w���6�� A��;z�׸�Se�cL��k&͏��Kb��ט���(���3w7
��|Bĸ���F�ױ�z�]-�-�T�=�S��׎�?�O�h���{���_�������ܮ�+���k�P��F*���kr��{õ��#N �᧙[E�x7��9m�IF}/P���q��i�t�h��k[`����%CI��ﾚ~�u�R����$}Ы����t��90�&&�r���K���ږ��Q/��_c�i���� �$�_R��!���Y�oaс�Y=tr.J<rTӢ�����ۭ�ʋ.��n����H��W��]�.Y�Rj�%�DI��,:�<+�¼<=��3�z���Pf�����&s��Q���]���e��9�}'��I`�:0#vwb	���=k���Y�L5�0 �mL��n9;}�P)�X��ZA����~�+pA�������jT`�滕ŏts��}+)�����hu�D(�z��,���zؔ�;�����:�8S�N����g�}|'�ΟgQ���3@m���O�i���C!�̺�z\glV3�x�^��S��N�ƫ=!��j���[��L�.E�f:mC��#>c�O��kH�͹���'��i��i����p�#��k��s�s��`�JUf-ʋ���(�,͸��;/FE�W��#��7��z��	��Wyo~/Ʋ�Kշ�Y���ᾩ���+ʳ]$��	���'���vw˽�vќ��f�ٷuѰ��OY�f���{TK7=rh�i ���=8����a�u��̏ �d�T�[�b:3�7&퉗=y�A)xvΚ�A�vj�^��w&)�Q�x~я�{�	����r���s�_u���-��Eո�4�JZ�T$Ǵi;��-rh���eel��S�b+�lC�(���p� N�YN�ye<��ٶ&'�E��ϱF/������wf�9���k���Nz����+���<<�Vb$�H�"Q̥sFo�BN�z��L&��������{TSM���]	�t+}�굅5 �%��uC��|S�[�<nͼ��˛S>s�^��^q�F�&���Bc�yp'W�(N�9��rr-m�`��#b'T0�wbQ�qZޠ-y��������n9���"|6 ��&k�
'��[��UE��y�,��\��y�b�k�l<�3���M�.��^ggNw"�TjZ�
�\d��SB��� r�e�0��u#s���N�ʫ.~�l���	
�c��48�uŹ�;��R��7��:�R�H]R[�㚔�zU)�8t����������r�+�Ao~s�c�!-\�<��P0Z��=�-�nabJ4Yx�ȦƯs�{��͛Y�&^I�!EM�,1uy�z�5Ĉ��"��=֔��\ge��Q��,%%��k�kDN�Ź��*��{�VNH
-��=G<#�d __&�
��U>�&�A���a1�Q�`S��a��T���C$GL�A��LQk}���GT3����ǡ��X��w֦��/�{vA��\���ُz��u��$�,N˲��4�قR�%��rb��
BOv�x�bo��[<��Mn1��6"��b��w4|T����ݧj������GWw��zo�5��v���Z��}/,�&��y���s*��������{�~�t�g:և)�|z
������u{�3iy�mvF���.����c*�G�nY��i��d6 r�} ���iv����e��M7���1�}����j�l�i�<��{��|͙M]��K�&p��H��+=�~3����A�p���$�V����ʭz��������N��9�G3𔝮�x���F�k��x���Ԥ34z;<jq�<�+�a{��Σ#9�f��g(���qӉۊ�C9jg���'}����T[��2h�q��Tqqv.�.d�}.�Z�ud5�7/8�+0$�Yaw�f�B��7��ic�M5P�bLm]k.�˫�f2�9ca�[�L�M�CU�,����o�fX���T���(�ڜJ��ƾ�(1�x����rzv��D��N��rЛ�ʪeJk�6�S�la@�̘��!��;�5��lǫ�$��o�_!J��6���J�Н0ЕJn�	U�թ��&r��i�3�Q�ơI�H�eo
���!2��Hf�v��х�8
1��?t�~lO��}���>���}9��
�m�i:uTʛ,J�~��{�"jSa�몪�J��Fc�&4|oG�rbZ�#t0f��m�yRO�.G�۶{��V��Vn�]�(��57�2[��J*��e� ׎^屒��=z\�t͹�;V������y���z��Ɣ-1�40ot��t�n��`������ )�sz�#"'��Of;�̶�H�|��������Hӕ����L?��p����	/�
��\�
j�j�:���q�5^�C�4�ykP�L!�\H�u�F�;!ۤj���`�y@���ѣ�gS,]�ڭS���ML��#r�U�M�I��7�:Ĵ���C@���K[�!�������Լ0����S�m��؝w�w#��p#�è�{�wJ�K[=���^5^�	�g~j�c���GO�Mι��c�鱜�7� [������llfێ/Ǡf2ZA����]ݬ�Y���˱e>T��;_����=1����a'�����MT<^�a���),z�[���c{^�{;�|�˫KK���*8��F�_��N1K���N����>-�f����Ȫv�w�7���Af��@{ڕ
9��L����
�ߓ�"����7����F�wJ�SK�4z+s��m}/kUӰ�=�ޘ����!w��R�n��,������7����4{�%�]rx�?��j��lp���C�5}Q�w�3:=��ަ��:�A,�^�Ǔ�D��H������.�#ް�}Y�ސ�⺊Go !F�W;L�K!��ɉy�����ӣ��ڢ|�P�J���q��\�r��O�0c13|߄�;^���{����!���bX��)����|W"dZ�������Ļ�\����B��ۤ�ӊ] �V��P�>;���daJ�+�?U�����9���&�)4b'tv<���ʹ���BK�b�:�+�7�reffыt��;Z���#�ۛ��o*����W :f�U�3�|Ku��������b��]s����ki8lGX��	k�a�o'���^7:�ˈ���i3ϙ�'��� c�9�']Ϲ^(�}k�b�S.�B�o��z��r�!�}�iIU�En�>��G˚�{]�Sv\����Jk&j���]R;/�U�ckջ8u^�k)��6ߏG�4�����Th�/��v
�ڨ�����H��PS33)�a��x;{�N��[g�x�7@�qm��D�Mc��$��.ڃ-�]"�܍j�3s�[�����ߨ��/Ϥ��d�^
?�}2��+�x�ֺ�wE(��L�I�:ͺ"[�؋�M��ra.��M���+X�5\�er�6`8���1YD���
���ք�y.Q9���[����8��-�
=ǻy}�k2g[ۮ�Ol���2��@d��D���!��!tm���@��$������B�>����7e&*��n���/�t�K�bX��SrxSx\����y|�o�6��Ƣ�U�*����UrN�E8�<X�]]����m����w7�C3������FK��Ǣ[��G3��+lѡn���ͣ\��(�,[�)5U���[�pG�ذ��JX����̧Q'5���y��\�5�5ü:��gN�[}����kIvU�Qn����г[���Q:�$;=KQ��s���p#I��;��N,4��J��t]Z�ڝx�̴j��l�Fd4sӦ�#&A��uf��hؙ��b��-(%!˜�����Q�kn�,u۸vme37	s�Ay2�*������F�ֱ�i�����5���^�xOdt]�}�tۚ*��ٗ�ݻfs�XΝӅe��(*�$��B(��{Q����R{*�r��N�r
R骆r;&���Whs8fGSp��b�f��
dZ@�dy��3�C�����kI��WēkF���,��L¸H�ز5��r7Ʃ>�?������Y6�ϥ���/"nM̙;�b%z��\�h��<mL��b�+�B�P���+s�$����U3n�9XuR[�<Ӛ��4n�Vz6�Ǣ����n��dK�u�6��-[�1�v؈��Z6Y��s�okz�B�|P�C�1��T���r��)V�G{�X��\1_
h��y��/*.
P��]A@���'e`�9�y�z̫0�@nۻ��}�ڢ��Ǥ�q5B�����=J��e1Uz��������5���W_K�3��ˤ����Atj�9}{��y�l��5F���<����`�M5U�ˮ�1�MU�</*�5r�w�N�+Yy��s�V��ج��#yǭ\��XK
���Z�u���i���;���w����<C�kj��ic�}�v���ӻbԄ����v%�{8��n�N;�8��FAMQz�<��>�{��*
��tƃ��+xц�z{)���5;�2�U�lE�$#wt�N�=��涡��:(F���Ԓ��k+v�z@74�;֕��{,̪}�R�d�;0��[V�݁���^<��3��aޱRG��>�Bv��)�j.\���I����k;$�I�������%JUG�~ �H�.�d��2���jH�1�o^BR��k����	$`c�O�=cǮ8�;qǯ^�G׏��!$!;
HIBz�n�����u�]�/=�F���v��]#�����;x�����8���z�>�||i�!D4�]~;$ш�����{�%	y��	��d*�#�ղ3�׏��1��q�x�ׯ_G�o��/D##HBI%�2�~us?8��\�.�d��b�fO���$�1�/=�̔�H������a����ή�14�\RL�p-Bd�$b��k��˄.\����O�"��""J��TR�H�K��z�6��o�E�����e@5�O~y�����y׋�i�w�\ē��{��W�"��޹��rf��=�W`���^:]��Ƌ�w]��J��t5����t=���o���J�%#��xQ�4
�N)-qB�q�xLm.D��6�1S� AJ#B���
8��YO�F�00��i�����Ŝ���5Y�)@d�4����n�1��m�H�۶�8I��S�E�/Fnl���RBD��%NF�"�b(�q��dA%����N8$d6�1C�3)�F I �ґă��e��(A$�h�"�e������IN6�� �1� �b�� �����p��AR�	PA�K���J q���mA�(&�	D�HȔl�)�¾��P,�3�d|����QB�#��(<��y;[�~۞��/�Fgm�����r�U�ڛh5��
���*��Lx�g�>�.�M ��>G�x X��G�I�Z��>�Yk)�KhW(�͛緈�R��9��e6:�K�r��4Mf\�#n^U�=�&Lkf�{]�5����zfdʳOs�.����ݝ��.Eᷥ��jkۃ�9f�'Y��H��-�5rpX�f�E����V�ނ�u�9o6X���r0��Sxˤ5�x�%ج�"�d��@d��ݾ���#���n��g�W��굠�]��~�a��]lW��v3�ճ�.���M����A�J;g�u���&|��9�s�̜s^f~Y��v���,��2����/ǭ�w�WI�Le�����n6����{/^x�qf{�ּ��ee���­	׽�ߖ=6��ޅ�9شcꎡ�q��9�0K�a���뺯'S�ƽx��xi��ո{GCū���wy��H=�$<& �$!2N�{l�vZ4�l��F�j�P߆�[��:?�[�kR��~��dNR���)��ql�M��忦�:��]������y��$�n	K������D�ӽ(�pQ(ۚ�U��������}�˙}�.� ��>�fwg�|�k�z����Go�X���Kb���s4e�v�5336�7��<d0p@1w=�D({��)��}��{�qS���\3�`�8{��h�N�5����ۋ@lF`m�rYM��w��v:���f�n�����y�L��~��L8�dzta�H�C�n��5$6�`�0��5x�C�f�on	F����C뵖�Ⱦ������C6ƺS��;ډ ��������X�1vP�� ��;U��������ká��v��~�oo�v�5N��S� dM��"�H0)A����PU�5x�7u��U[��n�Ѭ��y���o��垒�m�h]	a	��]�&���QC�ﶳ����v�L�:Z�k�.�3�"1��.0*��S��O6/}�XX���6]s����X���h�aZۆ瘖3�F�s�G��j���&s�i���e��χw#��iJL����nt�*_/[u�ڼ�W��~�|D�x�o=������gw��9���+��`�'�f�o��{}�����)n��5����a��{����&��Zu�{)]��W<��P�ve��R��&�P+2&�ʧ��a��*���b*�����|�6u�(��N�\���y+VwXI^��l�u=�w�*;^ǋ�i�s3��L�rE%}�^�x*d\�x�^�꧲��RΧ���̓X=�jz�՝�5��MلZ�~���:��\��*��4Q�����v�Ɖ��Jz}��}\hM�����(�q1��QT�p���Q�\3��'�Os%u����乒���|#u���pq��J#K���=���"繦'{��7�d����>��KOz��spb�+�22�f5x_~�U���6��h/m�ݶ��!�g=���w؈�t�� {�m��a%��3a��J�l4��V�ƎT�����zB��a{~���D�q�U��B����������鍇
��c;�)�r����B�ڦ�w�I��&��%]T�ϥH�z�f�4��l�Yy��+NѼa:����u��TF��4����ce��s�Z�u�v�}c0c��Q|<ť�>3a����dE�1U���Mɺ�i��8n'�(��5/���K^uFj}�h����B���7Qq�����K�w����z/}�OW\JRN4j.4Krr�|�������X�)yq�Q�8���UCQ*�K�KD�z���뤂P9h2Kž*d�3�!�|T}�l�{���x��h�z�C3ip�Fcrh9G��Ԟ����W3dDb�=Hc��w�Z���}�����d��Y|5�j�Y�<�[�^7��yB�Q&X����S�]��$��}Pg�Jɱ���+)�5s�b��ݱ�:�N�Ӫ�Y�;�9�9��.���ZYy܊���@�Ǹ�G"*�O�����Q#��|C�~ã6���[��+	ܑ�~uq�|lrc����7��.�tnh`1���M$���v��﷡��7oX!�G�QR����W���R����J5r�l��$ef`��$4`�` ���3�;�-�Ǯ�TKo��ߔ֕]��u��CnO�I�ջW�*z�[��9�ڲ�Ӯ�B���g�8�/��ӗ�k`������4��'��8xy����'Ǿncc��u}��GB�$rG�#�y���8�h�n��QW��8����{������tq�ޚa!������9-�oʳ�w�ۮ{�9��o����w^��0`����^a���LqWvs��4gO��j'�"�G�fu��ӖW�$�CE#��O[�m-��X�T��30p���2���ŶM��g���|�"��Mv�?]��,���\0ÍvZ�}Y�nfY�xhx��������|��f����!�� i��4�*s�f[�|�,��x ����PБ�����r��^E�iˑ�A�N��IV #M���/f�]�d���i���l��18�����_3�#�n����f�j�@_?������Ĝ߬;5d�ɲM����~b�VE���H��g`"����~'��t�?m��>�"n�Ux�2�2,@}T�U7D�*(��ְ�� �hg��fQ��-]x ��� ���,�ʵ�{�dX��t�����cOp��GDk/�[!Y|���9��K�f�/޼Mq��wB	^(�՜����շ�)ûN�Z��݈liu�Kl`J�V��G�ݙ����<+�¨�,R�&���^c��c�����ߖ`D?R�C�����:����$oL;{/	䑵��J�y\\���=�5��'β�7<�b'�'d����7�A.S�L�<�V�Q�If����h�1^��3.k�ͽ����6A��v��3�����&�=��Ҽ[�����r��M4�*�-��Ē	f����W�j���߫���o��Qӽ+WJ,{�mϷ`k���ӷ�hV��N���	��rz�� �bZ�q�/1O�YX��h�O^)�]���$�l�$ty�`v���w�q
o�A�rx0d�8�[E������ ��#yY�:��=�;;�lj]0.�@�*�⥰L�]��QdչK���*|Wyey"�>S>�Tdjm2k�-�Y5]�s�_XW;[�k6��N���s���hnLk����d�-�<=����zB�Z'v���z;h5T:��[�?x"��騮α�G��ٓnz�B����9�Lٜô/G��9�-*���/���.p�e��N�ډ���������ה�>�d����jKvֽN��ed�)=
<{F
Cv.��;d{���<<oTvȌ��O���n)��"�x5��>��l�)�,A9�]�b�d��*fk}q}�]���Όl-���6j{��F���L��ߛ�M�k�j��a`��B<��o#8�̼8�)�L�rX8B�9<pR*�q|�2�w�bH��83D��̲��F��O,�M![�ig͖�/wʥ�g��1����c��y6����Y�����&8�&��M�T1c�P[��<מ��*����[�"�Ww>' �>�'+ܤ��x	�TV>^2��XE)(�g��tV�޾�\�>��vx��������"sw��*�M:��6�˅s���6S�� r�}�� ��Pӽ 7K�bK��l����ŀ�(���S�c�dAuz�]&�f8l
_Owr�i@��t��Ol��ٖ'k3b��7]x�������H�p�+�!��y�i���tz���|�e������� y��[�����tOe�#�{�>�_�x&��,�w-����f�֩<�LCˡ��R�B�����1�(����h��BY��S�)*_�\%�l*�# Ur,T�9�w2_U�`��V;�Y���j`c0�߸�xxy��=�Y7�(��Ͻ�o�M�qIv�v
��3E^���0��狿h[8�����+&�u�J{�I�������3�\����Uz�{9���_5���Wl�mm���g��K��"N��_7:����_�g'x����z��^tײGu��b+��+���ёy���S�ŷ��z�)�{|7�q&��1��;���o#vZ����:� 8�k�p�X�%P����W���:ݲ��QF�.�K��D6�t�l6)|�9L���E�@l��Y1Pہ��=�dfs�FϏ�
�h�)��CQ�� =���6R�2���F�e�D�lv=��I1�%x�OW��HF��å��f^�Q��z']�+�� ��YFi�Д��ҙ�T���8�1]8nMq-j��SjνB�N�ɘ�d��k����0/6=��E���yA�[@��勫��?!}���HC��cwL���!�p����_%>Н�-/�3���{��4{�f#��,����4c�ܤ��a��GS$Y �H"��c	��aQ��t�L{@�B�[�pg���3�7kݛ��1<梁��'.��\��[Y���ͤj��y�9�󜒾��0#�;&�(�h�A:j��v��a���a A40� m�����fDШ���AI��y���L�d���ʊ�M�b�%�f�#o��\�1��=xkaM��1���۳>k­�Y��8��|�ϯ�_�>g �2è{�j�v��&6���GN�kp!=��5:N�_]P.���{ii���,A:l``�+���&�����}�T���܆���𘣏p--��Xe���"w���*�oH�*G���V5g`k��I�}l˫���N�d�����U<��F-W���I̺�8��&6:ϻ-_|<�����_�>/�B�9x�^�K"�>��t;��=����P�Gzu�>�V�����3����W/X������i��3���\�}z��y��QimFx�9��Xe2s�� ��H�4f.�c'������BD���Dǀ�ҍD��:�v�0fwR��@Vb��Sku>S5ɔ��}�S�M�}հfB��WC7�-Y��(Q�6����'@w�����+Ώ�&x[�EU�EAA�Z�5D3]oM��O4�����šuRWs�Ru&�k����l�ظ��g^�7�ߏ���یإ$3&x�V��|�Q	��Gl�CSj�a�Ǖ�$�쟫q)�Y��vMoy=�M ��ُYg���:F�r��4C��C~�"TG��zw�x��~�=���TGLL�Qz$Ċ����%���.t�p���j�]r-b�9�x��Q檆���5(������D]�yr="����OM����<l݁��(��������J�"Rñ�n��)��%�7��.�9�l�	U�9]찼c[��ŀ[����oj�sj�����1	d�����y�5'9���[���R ��`��uD5#7�`�⭦�[s�H]<{Ty�"�Q;zC;����x�u����M�`�N&���zC5�9���d��:tt�TWrV纱Wk�m����r����o�x�!���ހ�.�=�h���"�2�ޮ7|�6Aڗ�m�fq�p�.u���O^�q�Z���jZ�p�r�o�öL�j���d�W4�^��\����(g
Ӏ;1�5���࢛ؤӮ�����+Z�cm�3�u�MFa(J`5��X�*B��&���+u�ܼ�y�m�f�`�תOo��.�<�0��Vn���(]B�H���b�¨��c�JSSFx"�i���.�l�M�壕���خXw(�i�0H�N�yK{�6q��0]Y$�1�F�͹͘&Z]\�EVN�^Ve�FntP-����X���@v�n��ҝ���8c���Ys�+6����2����&[5�\��W>�o���U����(S�\���*��+C]ʴ���Z�-�M%&��ö�8M�Z����<h�Q��e�|����fD�$�\wF28'�C����no.�)Gjӂ@e��o' �L��Ջe�8l�M�Bɗ���s�&j4A)k�n�znS�NAs�.#OJ&�W�ړWqgf���b�j�N[M�RH�ݬ2��;� �(R۟�}4�ٜ�_(6�&��'/��KY����7!ڔS���n�0����3�����%m���,dw���<����:�r�%AǰSĵ��m,���!FJ�q��6�ׅ����G�O)v���E/*�t�W�wm���X}�Z�k9��ayi�4�����Ӛ��2�Ku�1ej�][���&G�L�ފ>�[#��ViΌ�z����}�:|�ݢI{�䂕���!;�9[G9�ܸ��)]nt��w����45CP̭�hҝ��7N#�"�Vpь��L��i�:��+'tx�u�*vެ.��탪�9D�Z��y��mQ��a
����}�ͷ�3�t����K�'���n�fT<��J�@��qwS%2p��p�ʭ�\�ej=KL�J��}�A��w7k��w��Ew�:e�97���V1�5�o���&0�7v������س)���to2�}Rʽͣ��SJ^c���Zʜ$�mZ�%�Wl�}6�`����-��;��aYvU9;b��mr��8nhU�*��1R�q��%�>�h9Sj	��N�����Q5V�}w�O$�)�/�W�dTݍ�0kw��(d��G��ro��X�rE|�<��nvX�����U�G2s6�.¨�iǳ��4�^,�zճ<j&p�[o�&��u��2�[�7qq(Z��I�x^�_>����3�;)����K8qR.Vs��M[B�r�]uv�;E�`�٨�M�*���U��ޙ�I<�U;�,��9�s6��oR8l���qѾפ�:�T�pG;�����)�e`�G���#}|�,8r�v����v9�ኺ^3z��v�e���zK����I��n���]����!I$�A'������L�Dɕ�qݺ
4����~n�Ί��X����qǎ=z��}v���p�1��ޮ�;�$ba�z��%�q㤦?�vx�@�	T��_Zx�����8�<q������~�����!")J�c��h��>u\�%�A�('�w�T#$�a$��G�]�x����8�8��ׯ��|||kA�)��ԩ�����د���&��;��Wn4�n�Jb�:�`��WEFS���M3&�;���%F��H�{�y#���u�ۘ�.�2H2QssO{�x���E�t�,E��/<\�"F>��#!�$�θ�_\J3�PB�:�ȓ<���B�P�Ƽ�ݸr!r���xi��+��^;��W�ܼ�>�םr��☗w"s����q��<��w%)�\�S�r�PY��ݍ��W4������]�(D���5�R/{��%�	�QB�A�/������ʧ	�ąz�][��v���k��u�N��K4)�L\ڜ���]�!����v}U�������2G=��K絴��֭�F��v�he�s�+��f.ړ_%���Xu�E�ŭ�3[$Y��"0vd�d�{_���\mu*� ���N�v��O��� 1Ҩo*���΃N�4�L����MG{]�r��G��k\V�,_Ye��N;oG����C�Ԁ^�����?W~��.����jՁd�6,�C�.�+3�l\��a|p	�9�B����hp�=3}��f�xu�x����S)��uu�]���x����V3i��I4�},��_KTk�)p�r}�>�eM�H�a38��n����9��K��`���m��4� X�e��)k���\m�gs;]Ƥd��.K������!�JPF�׊̚ob�z�[~j���m�&�oZ�ܾ�j�� U_M?)OO.U���f�x�̚������35ĵ�X�o�Α���x��g�rN��}���]��
��`��TŲ�����eԎ�:��L��a.�dН�-VޡF�Gt�����{��ڶ�(��R��,�U�3-�6�^ń�K]G(���ʒT{�n�L���y��o��+:�'�����d�&�FG�����r�J��Ҭ�J�⹷s����9�cs�3 ���O淎P��n)�Ѵ�Q�
���[��ꆥI{��4�$�I[ý{W�f�A�@,��`2�cb�Į�E��]M��ɵb6�������y��{���f���_&�����v����#�7��n_D�OH6�"���J�n@�ϭ��C_�q�U�śr�g���s�v�!;�f/�@��?,�L���c���/����ʼ�T&Z�e��>�3mS������"6r[9_v����M��v{�����8^��;�f\����j�TA�"���~��ف����i�ث�H�����kK`c������ G�<��c�}��%b���9�1c�+�e�E���B�5b3h�u1���ϔ<���JDM�9L4�s��wៅW-z{.p�p�	«p]l��k�z����Vv���3�I[8�mN��[3-;�˃#��/+aܲ�m�����5j4r�`�{�qXg7|f�.��h�}8�mE��!�:Wb]�6��Z����A�2V�֧L��U��ew+7{�h��e����c��%�h\ ��뭕�f��zL�lą#�#m�#0�"-��E�MS���'+/&�n��}�s�y[\���3��/\��4�����z�A�����7�ǀ�{Y��s��U����]+�^��)~�߹/�M�r#��r7��t�*�zK�0(���I�q�����$�/�DJH���q����SW<���r�5Aq�f�o0���riO*k
o\^��i��mZƷ�orǫc��M]���M�xY��S8l�w:V����Nxiծ=0�7;螥�g~]y���g��(�9�D�k��G�{a�P:���n�[��u��;���P~�*�ٕ��D14�k����j��f�i���u_��۔
9�6�dܰ� �.�2�@��j+�b���G�[莱[߳=w��������kNX8��\4>�����wSC��s�-���;�cH�z�����;;�Dǳ��0��m���ְ�A�N�Z��-�C�B�k��!E��#|M,����P4_d�k�V�_�4<�)d�5yd�R <��$ЪP�� ��4�{!���g9Ey�v������Z�K����
��Һ<��/�C^GO
�#i>�s�����c�*1 ���s;�>n	l_��~`�5>��k%@}0aW^�q�HZ�w�)���*���Wm���Ow�0���&
{q21nl�o\^Ɲ��m�(���阼 Qݶ��X�s�o����>d^#}����/�^�hB�-jv7��3J����=Ǆy2ܩ����T�z��u�D���ڍ�FRB'7�0MT�fb�8���ʅ��Q��Ч3h_3e�t�f��-�<��14��t�y�o��>�A�]��i�4i�����M>�-9�����9-�.�i��/��%+�¼Z�4�n�a	���n���ɪ��R�{^'f�&��.��DO)��jŜ�A��n�����.�5�z���j��N��e��6���;GD��/.�S�����Ej.`0���^���Q+i���WS�0�y�p�w���j�s�~_�;��	w'"u��'n��H7f��d�zm��5��6�o����muOQ|twN[�I��x������ ��~��$K�2EX}�]�V������A�qF��Kp ����.�`�<�TdJ�Or�GwU�6h�T)V��k�u]4��?�4�M4�@$F@����s�O�*��8	�ƀI�~XzV���ԍ��T�E�T��L���ٌ|5�Y�W/:����lf�d�1������)_a��N�x���6����-�;�#q��ns�c�ϗ�tt�J��(�W��^�ne�r��kM��{ �v���nΑ��m�텍�3���4f?ۑ(Z��]�~�գ�
Y��F��+g�Hל������"!8��,�����昿$
մ�y�D8��7��~a�!�ۋJ����櫮�9�B�^���!�3)��v��Z�a�����gt�-Ʀ��-��n�֪����\�����~�m#U~�c����w�'vRy�9ۻwq&�Pv�foeGCX�]�]�]��� ��y�S��v�d�s�$VnnN��uL�;;�^J���m��t�E<Y���j��]���s3��G��C�.�p����}��u��O!Z:��_��>@�w��\���7�j�ӄK��6����a|~�]/.�wvg�痑'��^w'���G��g�|	̘�N�N�娑k<姇.���-��҇P�_t����]�H�AM4� G9��L���Lw�/rv�u4;#Y�.6���m���.�ԧ�Y�ý��摯 �R���[�)�a��P�:�4�5«Sqچ����3��334/��5�@���|���+2�bΆ3ap��=56��U�\ͷ��� !eH�gkWX�G(r^���r@&�QY���=h4;}!��8�V�b�a���T!,���VAGg�c��U.�	V^�u4n���\������}Ǔ�~�tQ$��A�ͧ��l`�9�i]:w�����?@]$�fr^D����B/��z�
u�GX���Cnv�|�1Z�����Ɵe�7^�6_�׌e�{�W�y���l0����:y�^���X*�6?.��y�ޣ�P+}>��+i�����-�g�mrP�����@���a��U3��QYL6�~s�D}��/�������S�S�L�VM;�FYջ\任��
9�)1g!��6h_��V󣵉nwowm�JM>�s(t�4$�E�j�E�7j�d'6�P�J�&����#�W+3�l3T�V��9*���{�����ꮻ��Z�o�9p��Ɗi�i�����!�.T�2Ȋ1!$-�4�>��l���rq5.BEl�YJ:�H�{�=�A�?���)���w2?_��d�>3�L�uvЭ��͙Vt�z:f�黱�r;1:;ϤC0��7>�%�Â��Zxo%�Ǹ��;+�]�ϲ��w��~ׯT��V��W���l��ey��wk�<�U�%\ny�9��3��)]l��|ܨ���v���!�� �x��%�WY�ݭ�eTn2rt��o�]P��
��di���e���-�o�;��Ve�b�:&��J���F7v������\�R���KY��ۋj�k?�ꭱV�/`���Wo��̚Fb�� Q�k��P*缪�23��V�Fcf��O��>�R��ӪA����R)��5}&g�zo�N��i��a�o�mڠ��QE/��M瞵��g���WnT�Ta����v���s���}�`�f<�ό����\f�d��p�=ψ[{���������9/7��w@)��Q�k4r ��+ٖ��sdy�vj����m��A�	�&<|�ޫ���U�բ�R+\�5Qyv����ٌ+����۸�Y��a�����=O9�ƞ͎�����p���gb�ٸ��\���@�p�k��������$Φ�&�[��d��YZ[г���E�����˝�k�vټ JAA�l؈fu:1(���^Iv�l��Bh|��K>�ax��D��\�~9:�dA�"�h����I����@o�cVFm5*j��B�":�_t�9�~nܦ��Bo#B:��bՔ/���;��3��|���cV#1�VyPb���6�����J�ӘU\��)7��c��f؍n�w�������p�1~��Z��
�<�_V����0��k�n]5pU�+!���r�����נ��`�t���؍�>�>3�R��B���I�u��y���N.:�N�=>�m4��
~��p�|��������}�bN0���g�����:KP�Uw�A6ɶ<��$-��v ��͇�3]u�w�Z���1k����6K��G췮�����΁[[W�[�,��r��we_Z�_I�V(r4�m���w����w��9$�`���=��@@�&,��g��H�f�s�)V{��CqcV:���襏��o#M�(�u�ZB�4��R���˭���������o; &�74U����x��a��e��T��gtǦu-��\���||����?!��ɳ\|z�h���Al��6�G���˧�R�@�M��x��L�e�"Z�yGhZ����SF�+�]-w mG�Dq�q^�n����K��$�x�G�ɺȣkk&�\��X�"��Zp�����XKKT��]��`�<�85��~zFcc���؅݁.�k09���^-�!u�M��-�z@r;Q��Z}�@�t���u�%�7rY����HE�?�)�����y[�t=,���Z��$,��wKK��0}w��3�V0ptC�2)e�0}�z;v�w�����I�u�Y��㘲�0�l��nm�	{�Lu	8E��dѳ�\'u?C��:��,�Ǟ�Q����G��y��Q��܉��6�D��M@�.��,I��X���E�+�B�c�6t����[���m<��#�w��2�m���SU�����Q�hV�QDd�}�������ԪW�-a+��r��:k�Ug����M4@$e뵾���>|�=�j��&���&���k���CX�n67z�������{�`�j�B�>�s�k�#'��5�g�pr4˘�����Ul��Ǟެ�x�,�hP�����w����p�QR,_@�f���߲���d�]��j�|����<ƍ����C�0:��WFwL� y�9���[ls.�ء�z�{l�9�V=39��Y��:6;L
�-�4m�E?u���U2/}d���C5�	~#�rJ����u�d�S<l���ܯ�lӽ�8�V)|�v]�ӣ5pb���0��M�`]��`Y>)b��`P�)3KF�E�unUB����j�*�-z����>�';T��	�U��tm)��2^Vz��wq��r�K.��z�Y	.��uPJ�v���@�p���3;2j�^DW7��n���}�M�"U�_�ٻW�Ϭ�=­�ا��0e�L��:������{n���-JZ"��"|��p������˾Sq��"�3����uv#�͡[LVg@�ѥ�^B�-���u�j��2#���a<�����P���0�젷8^
�X�=���P�J#�(���xbW׸DHk�]4I���r7�;^�E��[�Qm�2�]1��ez�-���˜X�FS�DxcJT��!�"���I�.V�*=�5h��׳����2���[�`��e>�܍�ފ����#:ݘ��RD�h(T[V*�Y���m�q�5e�[�%js��;�Ze�Mv퉽N�,b#:�*P�ѣ��c�V�vN*�{�t�g����ޱʺV/lȵm��}�t�K3�$��%[��u9c���1���uЖ,຺c�h��L�>�������g$�^k�N�Z��(��ì�#(���!W^_��
��ս3_�������d��5>][����m�U���;	�U�Q7y׼�iѷǸj��%ہ�3.�u#ݩma�H�f�o*��F�]}�* t�qUj��!�/���{jWo�7ĚB������j-*:��V6�lӨ���_�i�2�<���u��N}�qQ�1�S���y����5RF��ֶDd��4��YW��.���wvJ�ބ��:�����u4+���J���]��Q[+(оHQ�qv��)R�H�m �P����']���H� �"�Ý5�.���ʂ�v�M��nS4!�q�a���uʜ0��P��%;vq;�:�X'�q|�.�����j �����6e^f5�[%�Z����3.���� ��k&�y̪E��]%�[�#��a�[9x(�(��#un��'���U�y�6�_+�����];L�9lr�\�rW��J�U�sA������&�{��q���jM�f�Ʈ��/�w��y$��s�n�]��()ok@���Q�#2�\7wA���Q�;�5U{��u2������a����t���;J��E���B��ͳ23���@���r�r��I�Y�޵�O	(f�y@<�ܯ5�Ӊ���.��ҍ�W�qvֆ�9�XR��;�	xo}�Q����i�e��d�慳F��T%2�ڈ���0e��n�'�U��+$��R�o�=�+7��=����j���ٖM�'܍w��se\!4�m�z�b��{1��NU>��f����%��Iz�� p]�����Gu��ؕӳ{��S����l��,p��x��E��0�!ni���F8�̢؝ut��YY��;��ڲ��8K�/2)\Ѣ�l8�X�7���v����wKՃ&�ڎ@���I�e�{�+F�D[�ʗ�`L���h�O���H$��$d"���#I��q
MF���5��L����w�ǎǎ>��8�ׯ^�_X��������i"X��e$C	@�;+tT�V��������8�8��ׯ��|||kD��k%�{�!e�\����(����iy�6O�����)Q�*D�޻|v����8�8��ׯ���o�����Wa��M�����4I��PE�\�fX��Q~���v��)?j͹h����v�db>87�P�
5��h�(�ؤ��4N��6���ŸFѴ@d��&�-LZ/](��A���)$VMc;�μ�y�b+L�4II��oڦ��%Io6(#E��b�����m�7��k�����ۖ�����Rh#����@ I �C��Z1�Ӎ�Ҝf0Q"BH�ۅ�CnDq�aD�%�mA@�
H������2?״�e��[��y0���[���6���J�7%���}+f�]C��W�ɂgG� �PSA���H�L��Q��J""D�b�⇊aaB�i�r6JH،�H���FE#	��B8�R!��l�HNH�'��d0�P�
$D��R?���EH�M-4)P<�n�rT�T5ș��%H��O�~��],�m�JJ����l�
��O��F��3��D��(�Y-ߘ�￿��۰}��y��LM٣Nˣ0F��^Q8ӻS�L��r7U�mgD�CR��0\�'��c�s
��y�>���6�ڣ�Sl�	6����w���G�n̊;�=ֶ��_�:���M��/�4q�T�Le��}ŷW�v�Lǥ�3�}0�������q�n{�V���X3��9��Iu�1�$�Y�g��<���n���u}���qi�%�[W�\�/+xG�>w��zKzu)��7f��o�5`�|�36�k��]���<sf����x��K��]�;����t�l.�yW[e��F����7mG1��k�y����t�ә�C祡���ں��d��{�-B1�Ӝ���y����V��H*ى�\-3粹�{jq�r�g�^�ڹGn�MԊVN\��؁ffC���*k��v�U�Zۢ!��vu̶��A-�����*u+8r��]�&�otM,0n���`��#{����)��b�l���4�]��軚�I� )�r��Э:���s]�#y�P���hQ(T}��2��YGQ�p�}�ُ��\\Hfr��Qͺ��O�wO�>�Q�
_�DoWA�ܞ������ڙ��ǽ�'3�I^2A��|�9L�{|��}mT��g`�\�8������"b��U���+Fe���7>����.0��ʏG*��g���<'x.��.k�ĝ<r�@�Kk�dIݩk*�9s7.�X�<��wt�:{���2��lZ[+�0d�:�o[��-�KF��x������k �+ܐ:,��G�6V����)�wXSPa���f67C�u%�X��K�
���ݟ�<�l��:<��`�ؤ�k��C3vZ\��l?)��։̋Y٦�Sdu�W�ċPF�9]3�ff���}~�L����xV��#�X�GL=�䊅�Y>�f�{Evb���$v�y�7�r��Lәb��B��3W$a+-ޙ�3��:�ݴ��O��GK��C_ ��Am5�]%`�(��0Ƿ�M�Fj��F|r������1�2nR�=j�ߎ�	À����}z�7NU���\˅���囧w]�+���K��M_S��2n�k�{!��]v���K��{rO7DwT��;�@w����{��������;eP��oi��a���f|���E��fZa�)�)�D���@�i�s~��a��~:h:3�ګ�
�ts7f^��;����sY��&x�œ�(33�Ԇ��^" n�R)�FVN����p���&�14��a���⺯�{Z�N";Y�s�gN�p؎r"�̋�g���S!���be�J���f=-FԹ�U5�~��Ԫ�s��Bn��!t�('�NI��h	�[����Uk��i�N���o8���P�9�ч���;�fJ�W����8�E�.����h�1i�n�2��s��ѯ�kX�t���1�ƿk%\Q\���W�bE[I��͸���+rr.wT�r<j��>���u2G7��D�������wB�B�Y]���>�|���2��X�;J��Fr[�����2�0۶[��K	�-�Uf��S�����󺂧5��J�UIzpPjgn^�S퇖�/:��i��c��g}���.ښ{lu2�~w{�N�����!�I�J�&� (Y�7hn�Ӌ�.Φ��x��'�=��\���(�C���w�ؾ��Oe��"ƞ�!����ܹN�̈́�~<<��\<@��&�w�Қ���}�=:�g$4{�K�}Y���c�gK�,h��޹�֮=ztƮ^�	+��-�����u�'�����w�%���s�����]�oO��|�;�I",�/��� ����1�՘+Zv���o0:V��.f&�K.�i���6�����p��O=Ȣ'� ��8�O��a��S���fc,5�Ǜ��O��r�qW����eo�M��9C�ey��%���7���?��7Q��`��16d9�0��<�Ա��ѽ�:�٤�:�*bD����s>��8p�����XKb��F�������{o���e?��oi=�" �� �=i�u2�},�}��N%18��pi���FKz�VL��p,6F��P�<E�}D������y��}�Cݗ�U��c�݁�I��Ą���q��ێ�dJ���yG%Y����Z��+��3��w�,1�&-y4����y���^Эh'�t�7x�L5����v���'}3�G�Ph��&
��2xq���.��fܒ�6k8��r�h�Sdy�.��V�OZGSlS���Yf��u<�3�]�s����Lc����!"��{�ZEېdM!�����|�F� t�D��<��RG��Af"���K�,�$���N�mЬ30V'Q�u�M�w��Hui�sov9�q���G=�}�zg�<����z9��Y8ݱͦbu�6���gz�R+2-��f7�����"�I�)#��I�3R�?=-iUo[��i&�}]�>޳C2$��fX%lD�֫�e��qD�� �mkˍ�/�ݺ::�K�AK9�|�d;ٟ0[���O�_��q�h�'����J�O>%r������Y�~]�?���E0�t�,K����;\�IDa�=F&�{so�*w7�2��������ͺws/Su��(�v��@��);}21+��x�G,u�����s��	�� �Y�s�=!�a�{^Y*�#��ʇÃ �X;���f�u�Qh7n�6��m �;!��{�Lw�<��"����F\Z���=��A�-�=���y��]Ѽ�9�ի����;껽V�L�9�g��<���yg���BHu�]v��ڜ�U�ڻ�.g>,&]�cc��\�1=�^m>����+;Gw��s��[�>�񪑦*1���3�F����ǫ�s@s��q��WLq*R1���hx���Ud_����,��^��
x��&��qp�p��/��D��Eu��*����~< 0�>x�����mxhj!N�����h���w�p�yH����{ū�Q��y$��mU>��s5G�X��^B@�fg�*�S!}�'�?>�՟��������n"jSW��/䦈ޜ����L��3- `�����3=V}��gS�&����<�5!Z���3cL�L�8u�8#�cØe�d�����m�ǣ[-�Ǎ]�*�"�)^SE�E�/s�T��I$��YE.�9WFV�r�n̓�S�Ү���^�S�bZ��E)G�8�'����}���2�m-�Խ�'*'�݊WVP��X�ܙ�<�A���ʽл�7�|�aokqK�����^��3Ks����DPƝ����^곓c���8r������N�����;l%�U�x1�}8��wVoA��Q����D5$�@��f�A��J?"^��)�Lу���1pҍ�Wj��Rh���Cw:l��W9n�PJ͓d�rb!��Z.�Y�Yv(�y�i�eW^0�K��}���y����+x�4���Uh��{���n6%3w��t=I�w-�O9���h�䇫���j~��j���|۔�y������M��z�ץ���P|�G7������O@��=����7kFDv#C%0�΢hv�>����·�fI�R{P{�WF����w��B���~*jM~7�YV��5���T@b���7`0e��jw��q��1�ݶ�s���#]jh���y��������I�B���&��<��F�@�j'ܩ��K��#�Ov�w~:��a��~�_��#ki������k�4��J�q��H#&0��Ѡ����`�� ��l
itEW]���P��d^��`�'��1�w<P�J�]L��p�k2-�2���3��L��^�vn�~�eP/gHד�;�o�'}�+Y�pE[�<�뢎�x�����%/Rn����5}��+^Km�z)pk�xG��Q���x�˘��q������A_i��d^V��G+Չ��Uv�d]�mӓ$�`��K��#��7z�L��ػ���h�'CK1��Y�룵�\]p��?�e,W�73�{�>P}y]�jE"v��ԕ�^IW^��r]�x˩������`��W: �9�u6��y8g_�+�Eq���SW��*o~�h9��Z���0�I% �!%w����ŞӞˮ讆+�=��OJ�$��)ASf TˁL=�ᗢ��h��Sp@ڑS�жBTKP��$MP�yLi�;�L�X;�����wnz�ANۓO��}��c�׾��~g/w��RBp�H �	s��p��yP���fb���_�eO��4P�X����ǝ��V�[��w2s�̡nd���2�;��IZ�9@�}Q.Β� 9��$�r8�>��9��e�������dQ=���5"`��4p�k�3 ��2p.x�f�\�c�hk��,[sEW��o���]����%���^���^�8�lF��
n�4!�˅g=t��f��y��^_a�O��6Iy�(S�Q���Se�I�-�XU�Ĳ�U�!�qW�JB5��ժV`|�Ut���_  �W@Iv �;uk(��J)�J�2�h�ur�QVH��՝��^�]���39�#-�˛���GE��o�y�ᙜ�<���bF55�	.�MD�UJ����]�/0�Bp�a�08���1��|?s�fy�<�|ݖĻ�9�*pf@�k[��&�ny��A��1�x�M&�9���h�\�w_��J��p�fqQ�~Y�c��ti%�ړ�΄o�4����-�C��1��d2p���KWFp:X5�BU>���o�^�*-)����tΡ��Z������e���E�Eo{=dJ��~;7���'�*ǭm��i�{Da�QKܟ���X������-O�}�*�����>�s|��76�^$���q���}� i��z��F�>k�K�ɷ��T�B=���/y�EowKF�7�v���*�F�fESS�P��b���O|B>-�'뫫�����"�DDq��ogO�@�D�hNo��&\����/�rs�2��s�ۤ@�f:j,������Z�z���^����<���=��%^J%F�q�Ayi�	//q}���#(r�lFtss�>g�pX�q�z��\���/t��VE����4�nͮW����H����\�
�oc�/Gv>�lM���ZA�06�8��m
жB�GZ�=����^�\<<�������|�)d�>)�[�������~�d�Ӗ�4��`n��s�=�КP����<��Rz�	�WH}��m��=��9ӎ�zJ	/�[��q|	i�m�m�i�hL�0	F٨X���*,��l����cn�b����Zr4�~�^��$y�3�q�5�PRdf-p������33P+k7F�oh���z���C�>�oְ��N1���8��}��+��ή��\���j����������M7=�����<�#��]2C3GY�uC�^и�7B�ƨ�x 3BM�f�4�)����5N̻�oS�C��>����AU�ó�όq��A�X�u�f�wW6�y�x*V��#l�}a�ی��UН1�Jh��|�T���@mhs�b͟��_w���o��Bx����ܪ������jn���T�]b�����U~���jR-e�k�i9n��3$b ��-e1�W.�d3�h��jͥ3{A1�X�s�b��,�K��Q���X��(��m��,��W�*ݼ��l���ȍZr�],��j=!,�r�E��Sy���3BU���䫑�M��ɘ�*�6�3�r�o;��գ$ƨ=�i��n;$�{�=�-Qy�uuK��}h����kz�c��Vޭ}�fp�AT�=V��fit@���YX���$�*��gQ�*����jR��r��^Fީ~ιz����TLw�օ6o��{9n_e�N�l�j�E+���\y�������%އᢊ�*#������Poe�*���Ӡ�3)*8x��M��V!�����ʗ{��b�R���NU�oZZ��8��������dp�<�`��;�;�R-Zu��7��߹�ܶ��CvADt�9U�ݓ@��6��J�Օ�{jr����M÷����]0��:��q�n�,��\�sv��^K1Hn�pY4ѥ�.Kk�;sH&�TkyO�:�r��q��*S��>��
�6�]u��ٱRC�T�����We\���Z�yP��6!Ԧs���:��j��q��^�����C��-E\��V����)��f�x�w��#�8ܣ�2������W
'R�սr�;����!�O�hm&AX�n��� ��WG]<���OL�ؒ�f�Iǫ�٭�L��Qr}�WII!��`��/5IiZ�]��t�j��g#\�a�ޑ��ؑ��.�1Sۥ�%�ח��nzV���Y;u��yz�w���v�^�o,6nH[��z8Y}��}}­���Z6U�9f���s�YE��-[o;u�xz�t�ڙ��qXڗ:�cO_^��b;tc���"rه6	�kIʥA�/N0��m}AM�+ư�I����^^f��G`x���Y��ڕ��7�5m皖K���g:u,���:軩C6v+��Ւ.�#=VkZs*r^M��uDTږ]�lf�/,2������u��J�]���Y����[���c-m�PYr?v���9�C�'6�hQ�,��3u��v�SVQ�06�ۇbu��WvpT�b������IT_`�i�5ɇc�R�4�I�}����z�*,�'�X�����~ ��3Qe;��m)}�]dد���ui��.��QYS-ͣ�{��l8���{�2�<�h�}&��&��5��5l��v&�J��ab����,ή��J]m0�E����w��7�U�(�p�c�}�++%�hK�̸��6�N��TZ�\�B�t���ū�E�ȃ��5X0��QM�D��v"(�H�Q^��=\���J(m۷o^�=q�q��z����ݾo��TIa4m�k�_�t"#�i(1�lH��!���׏�q�q��z������I�*�$rII�VT/����o��s�����XF�n@�d�����Ǐ]�xǮ8�8�^�}}|i���k�QSq�,��1i��-x��;msƂ��]�&��W䫟[slb1b����W���m�-��ԝN�����FH��#[��F(1h����F���lz�4ck�si�h�o;���A�E�6��h�ֹ�o��6*��;��|j�6;U�fbر^+{�_V��6J�5��X�b�jW/��s4hwW-?��c�]E���\�}^5r�Mx���#w�k�+u�[6�iQ���&�α\.���I�J�#�V�ZX��y��-�c)�����V�[Ϯ*
���������Rэ��!��ܐ+���_�N�Vj�X�V�e��w�m�l��g�5t�6��a�?rb��듉,��95��-�X� �ȶd�q�R�,.�GK3v�p�-`�/��A�Du�:��?R�+!m_�1��ʤ�n�x��Iޭ5������!o�M�4�R6� �Q\����%�tgM�;��3k��yk$5�N�`�\l
Jf�oH�����sd0���3��i�)�9�a��6����9`�-��L�U)�f�p���ٯ9Xz�剎z�j6����q�$w�a�;h1Fc��Vy5niU�p� 8sx�=g�����c�����qo��gꌺ���z�@���a;F��ð1��z���&�W�9!������ϯ��{\��Q�!���vuA��fE�5���I>���&	��1w�K��tO4
���m���U|z�}B�.�xs��>��X��\�/<�{0����l��+9���~��*e��7��(&��&Z�g�܏1��9P'�(�c��5Ǚ�pl��D���3?��Wo�H�98xxxxB!���z'~~��~�[P��T��k���&�`�Lⷮqp1����s�w���E������ �8�y����d<h��V��]\��hFS�>�6���q��$er�h���O[@0�[r�e0��c�ق��[OOZ���tI�oT�X��ff�ffʽ[�����u �����4��XW��֓��[��3�П7���S��[(;�>z1����2��f(+l��U��/jv:O�C���$V����Trm)�����f�Zi�5�vs��X��e��4��ۊ���R;^d���+:�v�܌닶ث:�kbV����v>W�Y�}ޠ�p�����
Qx1��q&6�2��Z}u��!�@9D���4�{��]>kC��ճn[�H��U�y�E��wS�'Ux�Z_t��@�^{֡#;�w�(��`��ز�]̇�Ow�%�8	q�HuJKɋ*ɔ�QR�]n�ɪ��Z��YA��TYu)�rb�3r���:t��W;��l9�!����dv��̜�����o6�*X��B@�WX;�6���jÙ|-gr�|��gN�ʯ7�_+5�8��?i�D��y��1j:��U_{v�%���H�))(\1ClF���m�<D3��t�5qf gi�\YH㺲Ʒ/0�g`�p��p0�Y�����V��6C�{ImK��s�dD({�*/�@u$F����s1<��[�;�J;��-�5�h#Tm�T�V-͈�nS�?3�H��W�8iڷT�v��#��^a�ݐ�Mz�(3w��m��W��BC����� �����z��v[&q�W��.z-1�-YE�6t���\�e��mP��c���CnzC��:jvf��OO3-��3$	'�����=����Y���ϴa��E��{�VUu�Cgg&�/َ�[�=�_��[�2uSB4΀�3�L�
C�ۋwW���A H!"I$�lL�Z�h>�i���Sh(�Uml�=�gm����8ۼc��Ϛ�*��0`�,�[՗�:hM>@��k�v������A��A��=U֬���ݞ�R�I���ܩ�f�>75�5���Bx�����6���0 4��&d���x�L��2�߭�}�2�u÷�	kOW^F�`s%u��]��Y�.,`�r�N��,�h�g��HT�3}��o7��3��'7t�BU����v��jԕoVܚ�Kr���uv<79L�Ҳ8F��2H0yV��礪�檨���
�ʑڦ��Qb���$�2�	;>�<:-�[�<�֙��u��bɏLk�`C���p���a Wj��- r� ��*����Wd��7\>V�A���T�h����x��E_H��fj{/~��;|�]ˈuνG4�^������.X'���Ý��Y:��8�mZ�x:i�,�q��fǼ�{Գ�"y"�d"� �f�`��g���}FEʇ���q��|;1�ar�ʐZ�7�!��{�y��������"��8�5�]͒ټ�D���ȵ^�iD���C�.�eV�SJ���W����HZ���#�����ٶ�5�d0f5�`}����y�2������J�_�/e����V��m����q�7"��E��B�.g�&4��䜰-�a��̕��o}����?M����M���'�R��Z�9@e�du��F�����m��گ�f���U�wW��o���xxx@<!��=w
��Ʋ�O�j2h^�h���06U��m1R)��"i�,1�}�z<��kJ�MT�d(�z��H,ek(�j�g'_���=��ʶ�WK9�r<�?��{�}�y���Қ�cl8h��\N�:1�����Sy���V�ߓ3~l$4ħ�,mXK�)�k˜�wP�n�f�8w$V竎��*IX���0gH�]�3�F9�+��Q��z�� ��ٮ��/�J+50ff��fJ���'1�l�|��h+8jg��4���!냋KӇ���v�KbW^z_5�NM����1Z�����;�|�8;���i�mY��F������^�ۄ�nv1K�4�w��B��l6M����+����RSL;{���S�\u�����k��=a���|��j6�._W�o��l��X�:>sx�Y}�&��/YgJ�T=�TOh���[�j5s��G��Yoh������ݷ Aye�sjE�=VO���2k�ռ+����-V��Ү�ѝ7��Y]�����Ȧ��OR��v���������0#���s}4B�y��6�5��Q�%���۠O猅�py�oc�o0���C"O���E�\==��󷂩����8�]�9@Y�2�g��t=ι�MV�[�z�w��&�00BbAK��������|���7������#\q��Sc���v7( �lyƸkS�jDb��q�.�;�d���v����.
�a∼�u��C��������]�d>;$��V^�`�oTսmʼ�^�	h�;�������K3�V���� ,|5�/{��˿�7�؃_-�ER��^�����ӪY���F���Z�Y$����.��:�߾G�7K�>2�v8�x��3�Su�X�m��6W����`8���JoY��R>�z�9�R�r�%`d�wVm�0��b�f�f�ʲ�[)�p���ֹ�ƭ�R.)j�7�|�YҊ+&�x�kdђ�#Z��ER��U��z�`ٱ��G���J�Xv���<�[w6�62��wZC;c�.�Ԫe,}ؖ_]�e�΀���ga��K֞����GTY3c7�j�.q��}���9m*v1�.�>��U���!�Ry�!s
��kZ�A�ޱ~ˬ��}mE����\F�pƁnCNH�(% )�͝-��l�O��n\�z�<����~S\촶ҟ�ѷ̜�r"k��WQ��M�b�=N:�4�
p+����h�෤O�fo\�6wk�O&R��[��ڨL�puxC��գFZ�g���b�v��>��d��p���d�"jT_@ҧp^����2�
�X�3�1<l`�N�^B#QJ��\pZ_�'�-=���8X���q�vڶ������C��g�'����e��G4�v%]��Ly�F�=vC[��S{S�kcB��y�����SCm&6��p��0�ޚ�ݜ�y��0�3���/6�icљA�q;�6\>#!�_ӝ���O�}b��s���ə��A�$�I��E7��g+�ܯ���:��8��gω�^���xMd%GN
���Y��cH�ӳ���!�N������r����D����
߱�<��l�yC�룶���%���23.g{����e�����ށ��*������њ�s��'`F>'qUY���rAE�u���Y���c)��6ihl�R`ʪ�em�|���Pmv�ov����#������� �{��7N�����Ux��O㩄~O�|&��$�r����d��܅]���|��F�M��˅�=)��x�A����K�NGR����o��9�{�g#e�H�g�\�QT��IM�yҸ��0j��ٻX"�a�ȥ��"�����l���5*��o`c��$�͊m���NЌ=e��;'8�,/mzj�d3��롩D����9*a�m�:����S��{�+ʾ�蝋dQ�t]�BaS-J�\R�Od39#iXI�C-��)1C'�}�w�f����Cv�Ձk�j���粙c���jg��nM-L�W}0��S�w��ɻ�ZtY�z����^c2�p�1ER����C��C_��;��b�D�ݾK����8oU����M�5S|нk��^��-��G�!L�*�YӉQ���^	���X����O��:�O.>\km��eZ�2{Z�]MhĨOK��0���8��7+O����XB�}�+���̘o��f8sgo%X���:��1;�k8o�ާW�b�mY�!u�/��fw;Td�1���ksߝ��(G;��j����Oz��׷%�?��v�fmG �Sq��-^n?u���Rұe���a�w�3���oԄovP?7bL��7�_3g��/[�:��}v3P�i'�����ؾ�{3߮�7����D$�Z��j���fw��=(Ë�U:�m'��[=�~���邊�0�Q�i��'��i��ؖ��u��/j���b�gx��%�u�g\ ��/�@��o�њӜ�W����R����/x Ek=�x{�^�)'��;9蝦R��j��|v*e�nD^��}
�l�1wTe�R~�;��*,�#T��$�QW-[���U�tL5K�JMGt��Wm��,~|�{$QoJT,���꠬y��ש��l�^n�
��f��������΢u�5Į���Hw,�C��۱�G�wԤ��ݾ`M�Vn.LZ�/ά���5�Еq�M��W�M�^nnʩN�a�Y���5}��ކ�6��<C]� ���I�������k�����U�Q%t�h\��ܭ���F����to�Ң��Տzѧ+#�NՒ�Dh�����o{��;�4$�E�ǮWlz��&�%���{�n�	k�6=�ux�1�����|�0mD���BT�'�7�1�$�[�5�}~�F�Qt3n��ۣ߄r�6�j�bZ&[Ɋĳ���.�+)�k�$[���#���mI�9�ۤG^�}X_�����H�y�j���gu��\k30�[ܬ7f�;��r�5�Kg{�_r�����[�s`��
g@:߻��ws���/�p��I;W2���'Ҥ>疁�^߂'ж��v8�O���5´�[�Dnѱ�6�>k03H�f?�9Nq��7#g�]hUCV�hfF���^�g{�fpBq�_�t��k�o k�����F�vRY�����������>~�{e��B�"/�ط��?g9���*X���Ӳ�)Gvg5Ƅ�1��4	����/��������R?�� �_�*��G����
��H
���GZպ�7��{�YJ�j,�j�1�jjV�S[fLe�MJ�X�ZXʪY3mf,����jf�,f��2ژʙkMM�55i��MM�f�kSSV�Yj����֦�ښ���Z��SR�56����Q��MMT�ڦ��Z�KT�֦��55SR��*ݩj�Yj����֦��55��j��������5+Sk5��mMM�jU���5-SRښ����MMjmf�5+SRښ��ԭMMZj[SSZ�����M�����jU���55���MKTԫMKjjU��j���55���MKT�զ��jmSSV������Զ���5*�SZ��jjZ�SZ���B ����5�TB
D�i��MMjjkSSZ��T��SRڛYV�[V�WȢ�BA<b	�mj�R�T�6���V�Z��RԭUwkWZ�KRڪZ�j�jj�KR�T�6�R�֪��mT�E@! .��!j���T�-j��[U-J�R���KRڪZ�j!@*�
A �	*�K�j�������T�Y����ڪVK*�B*݂A�A&�+5iX�V�++S)f�,�Z��j�Sm]�W,f֖L�SSkL�f֚�i��Zj[R�2�,f�����k^2�kL�Z�R��mf��Lf�V�[,ֳ&2՘ɛm�L���֬��ً-l���XͶ�Y[L�1�m,�����m�c&mU������@�s���ED�PRDERH@�}
�����s���p�?��
����������?�G���ٯ�7�'� �����E�X� *�����  �����@���p}�����-z����?�?�'t~����J$���
��D�եY�KT֦kR�֦��J�ږj���R��3Z�����&ڛ-�YZ�+TͭI�EjŰ2"���(B �*B(?�" ��U $T �@@$��I�U%Z�+j��)�L�I�JkRʴٵI�J�Ԧ�4���Z��M���TٵM�U*kRͪV��֖��U�e�k-STեl�J��6٭J��mKjZ�jmJ� EX(DHEB"F�_�
%��ߩ?�� # ��H
 ������
���u~>�����!�0��ﯢ��������y�������������~"�
�C������_�;_� U�(~�����@DQ�?`�� 
�O�����h|	�

���O�~G�A`h"�
���Ho���܊ *���1$�������\��B'�?h���PW�?��@_���,$O�ZC��(6�ʃ������������ U�6A��t��������}~&z���(��L
�hAE������~Ф?D���d�Mf���
�	f�A@��̟\���7�����V�[��4dm�T�I*�X��i��������D"�%P�iA$�l�¡Dm�$i)5-�!�a�h��R�!��hm��KLA�fS�J��e��[f���f�Km�UrkYTS��6��i��36�j�s��Z�ګ�wi�����"I]��Y�I��3m�-����i�d��j
�նŰ�i�d�L����mY7��X�Z5�l���vԝ�%��H%EKd��fc45j&����Y4Y|   sv��lT�wi�N�"M�Zɪ[gt�	
��h4ګkM�.:��v���+[eiFӭ´�h��us���K�[r�:�
9���jl���ڤd�mCb��  �=
(P��;a��ks�(H�҅${軅	;bD�
�;�ݬ��R����6©TYl���6����vb�U]�p�6ճ4)r�n�4�5�ڪtK'ٝ�+ �mjEkl|  ���"�j�YMh4���+���w��j�mEV^��Cm &n����j�ecv�t�[m]nU(���t֌�S\���gY�"�Z��5��Fز;� �uW�����ڨ*�U,
�ҵ[dPj.�:5-;�h*I���9�]P�]à��N������a��ܵF�؎�U%vհ��  �z�oDѳpP:Viw}�h�C�݇��ց��ݺ� :6�s�U%u�d�4
u�CQ�h�ִ�A�5������Z�m�>  ����[U����ӳ�� �S4�Fe0 T�u�  ��Z;p:��&;8$U;T�>�P(s�ݹʬ�6�+K��ZR����  ���tiZ��@�)[�sӥd=g:�%J��wU((){�� ���^�+zU��l S޼��@ oW���<h�*��]u4ڶ6�J�8�   '>>� ϓ���
V�N�=��z(�\�N�@n{׃U!"�����9��
z�z(ν�x�C�E����`V�X�)jjV�   ��E W��۞��{o zW�UW�X�Ѫ����RJ�����ǯ]�T�.9
k@�*� t���H�9�4,RM��ql�XV�23>   ;��>�����àR]��ؠ =o{���� ��=��ݚ*à�uyn�� �S�=$,ƻ�@
�z^z���S�)J�L���$�� S�S�T��4�4ddO��T�@h2d1�CD�U"=@  ��*FUI� hf��o���eD���ʣ���\vF�Pjv�֏a��]��0S�Z��b�𪯾��m�<x����kZ�z�UU��έ�km�������յ�m��U[k��O߃��Y��f�iUX�0)�q(+�M�̥k��S,f��-��u*��VыR��V�̷ZN�@� �����
:ЃP
�L�m�Bѽ˽��+k�
��-��H���7Vk��u���r�o\̠Ł�4	�	+���x�Z�u�G�P;V Gwq=\w�LE���Iç�􀬏p�6��z⹴0+�/m��V�!�NIIԩa��Pa�v�6 �K,��o.º+t
f�����P��q���1���r���b`�l\[���.�BHV�x����:���˳A��|Z���`�,�	UL�p�O6!�wt��{{0
�b�ȵ@H.ąTgЭ;e���8�h;��gHW�oV\�o�Z���װ�l+߉�ݺ��[Z�l�G*e+7v�^�
/���Xۀ�Qڼ8��%�m3N�ݎA�E%n[�Ƒ��ɲm3��VM�bڏ1��4ni�DL�[�l�5V������n!��)U�j~c�w}�v'���2��7�x�&eD�FƼ#oAJ,����Wu��%XY"���!��츬�U��RI�j���K�IF�m��n�к��Iݹ,�W����[Hhպ
�����܀L�P���R��b�5Q�ib��\_�im�߆s�rBjŞ��P�Vhm;�I(f�{&�u�l���xX�F�(�ʕ,vp*E����H:�ml���
�e��n�mjقX5oK ��h��=�{4X��]�D����`t�`f^L�ń�����7G��bN7�-�F}�{��v�@h2��wZlu����]϶�A�(6`�̰�(fee���:4�5j�Z��wD�V�]�
��{���
p�A��^���*�r&@��Xw��a�д[6�As��m=C	5T�+J�:�6k\�n�\hᔲ�����DQ��f[����1b4e�Ӻ8Ӏ%Gv�0�i� j�t��Z�P�G#�m�
@�<�L,��F\����`r���?��"�ݔ�e��ݫBËc��-�cV��V޷�bm��7T���x��.�(#4Ʋjr?��"�?d`�c:0n�đy0Q�l��'lJ��LZ!�Q��4&��UIP�xH)U�l���	oBV�-èL�d�7�u���qd#�@��K�t��)�A�٬��L��0�]4��/Dx������r��iaB���5�ʥ�I�Qem,��Z$�yKq�VcF�(l�z �m�eu��۫Xl�S&�@(1�mn|������Dа�ɔ�rk����U��������j�#B7�uj02���H% 7]�I��	�c�PmS����[O1�[�R��g2���d��a廳\� �@�~Y� _0ٳp�H�	R\v���׈�c45���x�K.Hf�Ѳ�����z����̓����c��Q�Jh	�w*��Oq+ƀ�5��˶v��&�A�H�7{#8ԥ�Av�Y� ܙ�ڒ�֎k�wOBb�r��V
؋��ì���lq�$a�f<�݋�!͍d7Y	;�
ǐc͂i�t����W�w ���<a`���<t�$��!��&����k��D�:-Ʃ��t���l�O=O����qhPf$H^R:�%Y���죃^����Z��6��qMLm�5PQ-�dYt�J�!�/i�n�*� A���W�t	��_'zF���b�t��bɵp:�;�7u��b�W$�v$BF�-�F�Ԭ��%[�mn�d�ō^AyZ����Y����Xc��*�]՛�̎T�K�r�Q�a�ݻ�ŧ�0ҫJ�zŒ��eM��3�Zi�25w�x�%7c B�]��Z��v\+-��L�Gv����c��hhF`�BЧ[q� 8�wuva�S��wK\6@���G5k�������E��Y��y{��A4*�У�/&	��Dǭ������sc�SL3s,7�-�A\��_��\�{I5�Ӭ���>1j���[e�巈'��߶�nSz��0���)V\�(Gv�c+V��S�����B�YY������S&)DSwz���2�h�XI�+��\���(�E�;�S����\J�ϴV�1���ܙ-W)��̍iL��$M�!��V�a�dAkK1UӲ���;�&�
���۳Ȍ��C�`�ui7w/[4 �J�Txe�Z
Y�X��۰727��=�F�kޜFy�B���삥F�L&�,�w�������6�4�'p��m��l������֙�.�����MS�h�9����^�nTcH10�U� �1aBƇR")]�Aup+RKb�>zh���F���6�ܙ[e}�i�gl6�6T�`%O0�
%5��F�R^�1f	u���j�2i�6�@�Qp�}��lH �0������-�繁w��1CX�d�n����J`� �E�`��Xxy�c���Xf�f�R��@[����Ug^mZ���Y1��)iɁŌaU5��Fd`ֵ��.n�ұ5^���c�Nn �����ҫ&�-d�.]�UvUEvV�BL[��%���(aɻ*�����۠;G\V�2	�L�u�.���e^�Q��YS.©����I[$�;z�<v�֦J)֭ܠT�Bm#y	� i���W��t~�Y!(�,��Kַ+e��^�©5��֤������,VD��e:Hk�u��{OLz.M��3Ef��|!%�t�"�ْS�V趶TB�(N��A�]�K��������IV;�Lb�R�N�:O*k5e�B̼-[R�H��fa���*��規�\�Wfm��Kf�����S�X��k�a=d��ռ�u�P�a��M.�c,}��Im9���K"�� F
*�H�.�0�(h؜���	�]��C���&k����l�DD�����7����I�޶1���5�䆶�5f�GCpYL<�^��NUm��*�j-[.���+CM;�V�Sr�ad�.��z��0���*/C�.�(��g���-׈l�zeM�r%��� ��bh�ѡ�&�40hA]���@�.�^�,Ɖ���-�h���m`�wnVL�
�	� �a�.Xڽr����'��u�;�In�ʃh�(R�`H�WR�+5��upV�ʹ�4�-K��&K)�5eǆ���V2Rv����v�I&LՂ ��Jm*�G��<�@�����Qxt�������6���kH[����q���������e��#px��Q��A8�,C$��z�
��b��ؐ��^��xN\�u�0���^Uੌ����P�^=VlڷO��_��L��B.�a�"���ym^L�P�����++%j�0+G�p�9���НIRB�*�g)�ؼ�u�ژtTˊ�3&*&^�N闖�IkЄtct���o\���UKf���-��X�F|�yi)6�Vr��
#P�Ú�.Ř����[�Z�0+��|B�KA���+N�P��+mn����Y)n�S�E]�AFuf2ҕw$˕�V���υ��c@�Utӡ���6���cYb��I�̡Ws3��q� �y5%Nm�����֕���5鈬�31�+��X�%2�r�F��[�iM����0�5��;�E!�b9�d���-ʴ.��+�o#g1����KMCb���KGl,Q�³E5���T�p]��)�ꗆ"ɇ"ؕ�:K������6.0oXX�2ܧ��7@+01���ՕP7cf�{fJ�[EP���T�3Y�m+f]'����.i�]�6 %LBc�42/j�7G#sEX��>@+���Ê��!V���fiS���p]jK;q��H���6GA
�P�����eu�Vm�WF�;oSS(PV���wo�g[F�at�'`��x���V���]i�d��'R֘��X�)dڱ�$Z�#���Z�	S��l��r� ��bQDq���YP]ٱ�P�t�� i�St5���:U,g\�DYP6Υ�%�AњůPe�f��)�&7t1J31F�p&�򘭻��7r�*�ɿ�"��$�k�Q�B�:��e�͆�V��� ��jLơ3,i��6�6�۹(�2�k1�&	��҆�� h�lӉGi���r�%����fZ�ɚ)8�fɦ�}�	�Ib����M���
c޼��q�AR�70;�m�f�b���-�]Ҁ:�yv���D�u!5g%+[h�	��I�*�ҭ�+wqX��&�/)M\�%6�C��,,\�%K%:�[{Fխ׋1�B�����J�{�-͵R���`�����*a�ׅfH�����j[B����5�w����$vB-��H�t ��k��jV�Sc�˰����4�ZU^���F��
U�N	A٫��D2>(����-��,k7pڰ��1��ER���ܐQ�G6�z�j�U���i�^ce����:���؈��O|}�k� 9�d��"�m�bS�.��#��Kfܘ4���v�� ���u�nI/.�:7�VȴjǄL-�]ȕLݚ�ՄTz�
�ΡO,����ѳ��Px�Yy{���e�Fh�+(V����rh�q8��j��0	evw7�8>���JAX�N���,�qe����"e��۷�mĔd�r�غn��&fT�$EY!v�Zr������Q��v�&�X2��ӆB=�O纝�{�Y�֙2},;`���ݠ.�������m�ӷ!������i���ej6��IV`	fi�7b@���S�*��.�L^|f9�j���Y��T����j(�vD��[̱wi�Mjv%� ���!|�E���WΖ��=���)�v)�4�l/�Ҫ�l%�ɤ�E��0h�rҹaTQ���[�X�gSa�k�)��l���q����J�RtolC��xi�Ҏj+9�GC'ʹ�)wH�E�1���n&љ��]��f�AY�ٌ�c��%:;��{{�1���(�T����wR�X�q�Ja���<��q1nK��$[���0��R���n���6��fLPA%;�JA�ka��h�7�r"G����H"مG�+)��dݤX���jR�d�à1{�7nFѠ~���0`���Α�*f�K��a�Lё�:�ы&�|%�m����ٌ�s%<5��;�!��ZmekT�e����"
�V�!x�Y������RÛ&��Y�7h����@Ѩ�i��;�6�r�q�Wemj��+4�-�%)`3GEQ�("VSī1MДVj]�w�J7�v�6p雮�JoN�慗2�+m:��	u�J;��BPȡ���`���+W��և���*z
W7���*J�����-��L�QnV�Ҽ;���Ŭ���y��RU��;Yf՚�S,��Γfk:u7cHXsA{lkբ=M�1M�`S�f�j�x���δb7B;
��0�a$�ʅfɓ2�"��E�
M�LyL%�s!��f��Ze����jS5�.�ʹɫa��(�'qn�(��Lۨ�f���Q;��u�T�+���`n�h�[*��,�yhd{ZVmi��nHn�E*�6�`X�ʳtZJ�ꢅ1����7I�s�����b+ON�,��K���=X�nU*���M2�}�B��CY%�_u�Hˆ��%�*`bjX�Ve7�(hn�p�yOQp��LcXk�u��p:v
�4}��ʽڃc�J�,`G֨]G5b�v�t�6�9���z�� i�.��<�b��$��"FS�֊�sV�Ѥ�%���ZT
�"���u���Uw��.�H�T�n����g�oN�K]+ll�i�l �:�X2=taKI,֭Jkt�Y�F.e�R�G@PZ��ֱ�Ҏ�r��2�u������܇KP\xܬۦ��u�F�-'/S�-�woq �uw��cvEX�Zd����(�fX�U�i��#Q����9�\Xз��2�,�8��h|hj-P2�W,��LY6-ۘ]Ӊ��!q�L��-Rl���*04�k,\P���%����Y����c�b�Ygq;�v7X�)W�Z�i�!��Ԅ���+iX��4�/jC@T���wHV�����lв�`�{SX����r�Fy���1�Ũ$�1��MJAf㨭�A��o,�k�LT�d�*����\�G.�o&�0̖kz"XD���E�Ƣ�u��ѫ��J�kV
�dG.񨒼�Sf���'&�p��Fj�p,GW�ܴ�����f�n��_��0����-�*��A�#uEKK3)FH�zl�pe �G����&w*�����c������5�
W�5�Q�%ǰJ��E�޴vn��+�7�`��\x�v�I] d���Vi1B��`bfV���e����W�#2Qx-��W�p��ǼјBj��H��Fk��v�*K�����t�`R�1SH=%f���D��YK^�ZuM�$��������G�D����2���wX����ݵk�(�e�6�U����yz�n"ֶN������IecX�����j=:lrl8��Kr۽{��hC�"�@X����J�@E	��x�"�B��5��3D,w���rX��dU5Z�37T���AV�HViaV��Q�n,�ZJ���7v,��^�F��/N��`A�׻IZ�F����MӣB̌TN���A�(Z����r�+"} H���~��	Z`Q�4~�j�0��aU�E[����AV��#�Pi@K�?���Oe'�Kq�z2�	%�	��2IoN��K�c�`x�1��,��0�W�h�X��M�q@aRh�BĂ,������Q-�HH��;�O/Z2�_�eYp��m��r��ó�����Lu@��Cn��殫ݢ�q/�r�L�3)�u܀�$0R���;&��[��ix�f�T�*PCbH3J^G��u�\>���������_�ʽ����P�X}�>k�Ǐr`B���Q��:�1�[E��<Y=����o�r�>n��,�g�꟝�\C#�l^���^)+ �5�Hی��}|�\�<����[�u�ܷ�!jm��*����
��Vr�ٳˮ�<%��tR��^�}m$�"TUg*���K����J�wہ���m���T�8���\՜�a��β���
UbK��3F҆�ّj�4�e�_!l�u*�!�32�M�}74MgC%w�yk��x�C˳����Gk�p��Qj����<��Eཀྵ�Z�U�j��6o)��5T�󗾵Ͻ�����I�ilwR�u��*��珸�6��J�5z02�*0u���t�4��a���{�ݪ�GM�D����|���S��vVV�wh� �kah�G�Y$5��KKAY3�3Wc"�;8ĵ��Y�]�9���s/`�B
 7A_�.etY
O7Ĳ;|ڢ1>˫������V�Ҥ�M�2��+@�lFd�!�5�̝��U���]ŕn��q���p�<i^@��J�k+���t><�#_2�}{.�eg��R�rk��t���j_�VTx`�5b��O]�q�h��q_s��#�Z]>p���*��#�������T�'EmN�XzPF{��֍�^�^��Sf-�n8�%��a���s�S}}_�/�
Wv�J2h�>^ڇa�mws����&];w��$Vvq��{��%�v��&�o��ع��鴂5�i���m^Y�|�Nx:ڇo�T������i\�ʙw9��L���f�6�W�oLHc�����)���1��ejGʅG�_��h��=����t#�����u^���v�������M#2cn���F7}Z�D7!�#9�c�f`��$�}�Bj��=r�k�.���ڎ7�>A�D��vྌ[�
]4��	}��G�%<<p���Z�r�#�K����_[X�����%M3@����Z'���+hM��W����F������aż8��DHkhmхd�fXI�=.Ze��o���&�O�x���1�o+X<��}+n�ߞ�X`�0^iiuMD,)�o���w�IK�Y�w@�b�+��N��I]I��K�̿�b�vV[���HhL'O-i��Z5&��fJ��K�שּ�ZC�x�^'|����wP�����N]m�M���F��5���1pZ��2y����-%�E���׾O�e�dwk�~���]ۡ���U��4�i���wPٔ9xA /�m�RYf�n`�>��h�Ǜ4����i�6��/_*5�q�x����9]��#����f��uύ�D\���P�b�����h��ڶ�9�.j�1I</_`i$��g�D�B�+�����,*��搙�U�},�)��b�BZ$#�0>#4&;�6S�
S�Y�6��5/���q��Z�a�"�%�{u�T��tI��\�6�E��k��ĥ�`v���Ff4&m[��Ҟf�܂j�q�H#�ëU�7\6w,۬J���S
�{`ޚ�AFq���M��ol[.O������`��E85\0��6�g"
]�b�Ʈ�l8x���X�c�=*/���CV���~�n?N�L%a��C/C�zf,��˽�.86Kg_h,�� Õ�z��Or�Eb3�G=#�Gq%��䋽�N����8��b�v�ƭ�C@�g���9t�Rڻ��!����b{�����H��t#��U�,���/IX��q��!�a����nCn�(�wR�g��&�r��i;�ĻƐ��+����Xȯ!����yiT������v��"�sى�y�/T�I'�[ڄ���}I���x��u�$|���S7+wu}h~�7��ZP�<�ӳ/W`�`�ү�	��{��QL`���x����	S����;'�ǽ��f��4i�\��;�O�/�"ĆmIZʱl�N������R�,%fy�b�}z.�l�MvZB2��d;�N����fBk��y��EkE]�[�����-Y���.껹�$S�c�d7�jc�g]u
�\&��o���-y;���R� �zcb�b]Z8¾�$n>��
ZJ����=Q�e���nY���*�n.v�w�]�UNNG0Z������D��n7AnVZH�>n�R�ֹ�n�ka8�|G1��6n>Ѿ03����`�heb��U
��8��K��y������29��1������޵��^��&z=��sD����Y�K�k�?|��z�p�ZCo	���4G{���]�u�f��elC
�pF�13[�U<B��Yy9�u8�`����l�ꋵZ<�CJ����w�4e��C����i����}�/�/}c����	xe3w�k��<���d)�a�[��K�/���SHR�Y���{h��.�%���0	g�Zt�ҡ��Q��6��V�%rǠ.�nJ<�<1.�ۏ�tُ��/�-�/�u9��ԏd�q��F+�ufn�����!��'Xl�)9Q+��W`�3Z��۹g �	MҪjpn4Fj�<���q�o7"
�WH�R� �Z,�a-a˨��p�tHf�WU�1�X�{5���Jᮺ�_> �v#x9�Q-xx8t��%��3���dK�^v#���Q>��U��;ܣ�ݻк�E��z�:��Χ���w�1p�n\�t/���r��I^b4�b�!^+�39k���L��z�+,t�Z��/�«Wզi��%�gp0��;����OC��ɗO��#A��˻�	�]��c�|���rj�{�I��8Y�W�a��oebc�⹾d7ٓtM�yV�q��1�m,3'j *�*��v�d}��U����O;8��;���w�����87k�����'a\�6z
}�����.�ek���jo�L�Hy�l'�QK
�ې�lJ\�j��e��7z�n^���-2��oR=hmA0f
��d�\��:�]ѧw���ĕ��Ŵ�T�!�j���ᶑ�5nof@�Z=� T�4��}�3��Ûα�.���'����p�(�O�������/�$���LKoUh��&�B�:�d�j�:;ث����&iv�@dj�r�<���O%ö����HvX\�����	Y�B�sr��JP�*�0����)�&vL�w�N�-b�p/��'��?[@�FU���Y�X� Z��n>�����Sh�,f�|�kW�����7"��&���L1�,���Fv�o��T[��.�}z�2�47�s�tR�8��vϰ��ɠ\�g�+/Z�n�v`��J%�@��rk��������OrN#�仕�3���f�IB��s�u�_+�ZՎ��"�y���BB��u��,U��ꇹT�.���h5-��	P��N���E J�ˬ5A%@�d�ށ��^ ��*f$�+xң�<꛼p�7�V|�Lu�����K��{U�^ہ�SN��kOP�)^�wV_.~(���{�H�,546`&U���kk�wV3u�����T�����r�:�/k��R2��<�+vt`uK�n��g�K9A�ʶ��e��3�Y:�F
9Y3�ֺ�T�G,0-C&��1���Q<��5�����@W��Ѵ p���x���9�����T�Y��٫η���eX�'���Ρ{����|�<����*����3L
a3`�C�$2�{g�bL��4φ���p�!et�ռ�;V[��Y�	F�v��*&��$v�7^c��T���M��=�Q����ָ��ȫoܬ�s��{�b�N���]#1�r���k���l��b;[�0	��:�7�<'V%w]'�V�V�Z�DQS���͓l8���.���1����m3�Ў�)p��[}�>F�O,[��3d�GO<Ot�S@q�C+P�+8�J�sN�xm�L�Ub��V$8
Ol�b3�F�T���ί,�~���.�s��XC�[��3j��qU��J�a-(�]�V��*�Ŧ�u�B^�����7�
�V�E,3�@�����r���0�Pj�����ٯc;
��ν
�:5[��ˮ]맡���1,]c��j�su����ܷ9u�js,��	��S�뾹�Wl}ˑ-�+����ՐJ/���� a�V�F����(7�.�����p6�~o��U�{�ԟ"����v��\���c��r����X.��F��a���"� �9.q� ��s*��W�@`����V_^�]Z��U�z/h�l5�[�,��2���CX`�{�����,���6�]b�4G��fm��a�Ӂ�;C,��y�m�R�*{tH*@�R�
����o1ĻzЎЕ�u�Łv&!���'����(�[���K���F��dj��z�v�odl�a~��a�9J��9�zE��N�s7�O�?kF��j�x�ˤ>���P��Q[e�w�2���RՍ�:��u�zY 8��<�#t0pN���SyI'z�ƳOm:�a�� 3����	�����a��9�Ѐ�����v� ���/S�K8���_��^Q*��w���4OH�|�8��kv�)���dB<�_�v?U;(���}7C6�د��J�[\��/�,��&�BQ:ͱ�I8u.E���[R��v"bY��'&��zZڵ���ʶ�H��ޱ��w^��tᙨj��-�����y��ssP�)^7�d2��V)�=C&^�u^62�s��t�F�t�b��w�7l��xeGts�ќ����:�����w�;}�X��꓾���r44�\�����Y]��>*�v��ԬK���og[��}�8���|6� ���=�$]v�@��-�>'p������sm���T��S@#�LUg���ي������������12S˖��"k(��&��G4�۵����Dn
*u6�P��S�����&�R��������͵̜y��Ͻ{Ԛy�����C��;�M��MVBd�Hj����!��r�f�Τ�{�}*x��g��v�V�y�gdS���n�B����!�ţ�s���X8�vc������x�'"�������|W�K���7Y#i#��X��^h��b�/��<
�*pX��⮝x�)xC��H��Ό|�Ļ0��:�-X.j%4�W� �#)\��#ޛ��,y#g�x�i/�t!�o��ڲ���C���P^��)JS7|�¢��X�L!S����{�. ��Cn�X{��'Afc�a�,nvڽ$U���[�>�PtMe9t�]
2����٬��Fա��y�k������'l�̦�"c���Ļ��)���W�厹v.��`����E�+��-���l�w��,Z5��0+s�k�����t�`edb�%�$q)|���}V�)�.�Хoo�{�.��\^&��Rg{6�T���߽|뛛O�Fpf�4-�}<�����
�Ԋ®��yV柂+8�6Ⱥ�Qz��I;*Mϖf�@U��0�	[�文CFXZ������c_��3���M:nl7�l�簊=)n��}|�����-;:�(ʼe�7�D�pq��r)60�ҋ1�&���]`�	|������@�ڂ�����v^���fЗQ��B7k��,Q+�XN��^'�jބ����wr�8�,��K�Ϩ`ܽ��f̼���n�=	�� �2��nRYh�Mv�qŵԥ@���(8i��e���V�{�t�u������.95�:�*J���ĝ����T�F�^WN���K&J+��z�L	D�R\�a��R+̕���xꁺr������5��� ��4e^2������d�m�e�dv��1Y<��gk��
�����j�vsRlѢȩ82{��D��X>!�D���k�����Tl�x�|C4��4�-�1��C8tb�o]�޲��w.��z}g��{ާ��Cn=<���xվcM��sM��8*R��yo4l�,�ӄݜ$8�eՃ��y�&e;]3}��Z՘��_8^�U��f���O���N
D�j��ެ���;�X//�h�D����aU��o[n�4�B#�y.�˳�;q���;��[iS���݋��Tq�7GI�H��t�qsˮ[{c-q줄oQZ�dꔣ�w��|�u���@Sl;9�]e;--�7^��k��Cٖ��\�ydi�O�"
i����݊J	^��t�naN¹���;FJQCϯ���M�9���D�kX��/2S��9-��wM�K��ut���K6V��������Ҧ��`��U �`]�NybQ��ul�ݽҭ�x�ҽ� !�5<�����	���{3{h7"wcD�H��������]��"��^�{x�͍}|WůP߫�[�oj�%��8�/a�O��(]�O�����#d%{��&�9�^���D����Wjw�'�P(�rxE�W�w�*;}�ed���O\>�}��ڒp�ұ�vu���*+�����>��;��ZB˿<�uި��g;�!�U�h�MCE3�~3Ax�45Rg.<qG7(N���od���ރC��_����� �|�Em;�Ҥt��AR�m�N͋�?a\.�Am��;�{[��sx"02x��G;�k��T����ןei�k�{�5�����编Bc�[��h��̉n0Ws �f��x�(�o��N�4.��m������a�J��[�G����sb΂9����,�t�1�B����3�i� ԝ�Y�]A�1�u�'� |  �� #���>����o�y�A'�"�F+:wIT�I���T�����bT_g[�v%�������紛�4��3���/^����<��n���qO�p~��T��
v��}��wvEԜ�Z&wD��3�)�K9n�d�a��X�Un ���mw����p�Y�n�u����>ֈ�`�{O��<��5�]{�2��	i��:A���*���H�0��Χ4��^˞�%�W}<.gQ�{�M�;80�T�XR�:��\����ʲp���/�D�2�)c��a&L�Q�=i7�]�a��nݾ����+^�G.
�7�m�Cm����ѥ;(g8�|���e���J��xl�h*�"h��>���|n����f���g�� iWR�Ei����2�oI�X�+������2=�֝`2��Q\/N�S^l������>θ�s����}��3�J���>���pc�W�/s^*���41���ٰn⇝q.]�&�ǯv���"�<_B/�D�\���h|Z'FR�1V�W*��l_���^���D9���O�v��;�@or��5������v[\��k�t����ۍ.U	^��$���C����0��m�#��/H��ݞ�e�>}h�Km�N������:�7�*�nW[�Z��(��D����h���y�M��E+�evkJ�4�X��E�i��Қ?M�໫���#��\u��'�|����k�ɤ���8�d�_H�Q��*�wW��Ӭ
��^)���oL���5��y*��0Q ^���z�F臇hw����z缒E<8z%�������
����c�S��o7�:��xwu>$y�e�<��G���m3+۵M��=ܒ�(��/>Ʃ��K+�	Æ xM}�|]�8�K��k�n�@Жs{R�)�y#,��t�!���8����n�ͳ6���RƉahz���i6��!s"H�R�8�u[����*���]����<OssGuqv�����G�T�KS��j��b�H-�k=v
}Ʒ�ji���mՆ)Vɦ��4��C�AP���u�rr����̀f�%�V�)o������,���p��������~b�Kw�Xj��N�.�X�ZD�����Ա�ٌ����mjT�U�f� ��x_�b,S�sɩLBѢm]ƔtU��p}�5-���3�0~����l>Fe#�{Z���cGn���wt̮�2G��a����=O���pTh�0N�!�vmMѝ���?*���v���_-���=��(�� ��Aϯ-faw:��̏R��l.�g�჉����BpȎ�]&�G�;���#K�o�Ac�7B'�}��ͺFG���*' �/+�����b�2Qo:ӱv��X��#g-�Q���H�s:}qM�aX�P#s.�)E��L3P�W�C))�L@,�s7�N gY�4ys��^ۄ��Of%rqϘ���`)��^nup=ȤwgjV�{@S9ٻ�So�.݆�<g&�r=��T֒�A<���,�*/N�EZ`T�:<���*�0�I�k��<{�,"���;܊�Ud��)WZN��Z.�Щ˭�kmW4�a)S�I��U�#��$�{-L�y�3q��8��y�[�z�z��;���ی��X�'1�,�Š�n���)�N���qCj��Emk��iY�����c�&���Q�b份C.���*{���6T��<2'ʒ-�r��V������>O"����Ђs��h`�낥�&�G��3���U�q\.����֑� �����K�wlO9$���P=��<���P��|�%����V_"��*��^u��%<�S�2��iW�^�w�d���cz����'0�=�մb[WOZ���Ĉ�c�f�"y��XF���G��K,���������jY)��>�5ao\� ��C��<�&�{]�b�M;ǒ4VFaz&d��
�|�<w��H����WFk���E�J��/=Z�L��QwdҺ�0�זϢ��{/�#o$G`�YŒ�M)����R}Ұf�����/5�9z���`[�m-Ah��>b�)��GpK���$轶������'ml�$���9J�)(7�eb,��E��nv٭�q��P�P*l���Vr���]:�p�l � ,��=ڵ�l�i[����	�)��r���Ay"2IWC��8����Z�;q���q���N�:>�GV����I������,�\9�r�2�SD\�f���1�jj�auoR�XWމM�ع�;������Y$l1��?E�B���1t�J��u��b>j�W�i��eXq�2�<5�Ѹ��[c&�wu��wn
��t����$ Q�]�o�ՅQ�@b�ݮ�x�Xm� �u��|us4�-��6�������.�>�����=�Y��xӌ�]�oed�qv��;h�V@���
\4�i�ne����f�\��}N!�j�=T{�wʟ=��8�xa��(���%�[�%��j;�e(��l	�����rF�b�֜��ŧ���g.�P
�,�̼��HQZ�׃+{�͡�^2���(l,Qu�j�ۺ�8˅���H5N*<����e�=�(*N�G�X�Pkkg,�Vb�l��'6M]�k.�ܶ��a�0)�O#�!���=Ȯ6����|0Ox�}(X��k_b�sy]����d>}�{:yz�
�(�,�t��Nɹ6�[�v^�N7��F��[Yg_��O)�՗�\��㸟���S�;+��\�7z�e��|1]���4^��NTnZ�+��-�|:N�>��r��H�d7.Zr���0�A��=Tޙ5+�H{�r� <c����̛��ûe�l�ҁe�8�־���6�t�݃�ri3i�BV���ǻ_^
�uЬ�'v��{1JZe��K�ژ`'Q�Z��-t�H�-�v�?X�w5��v��8��=��ܨg#�c�Fz�W%M!�ά|�i�F�d�9��á����&_��w�̟7;��}<8��$�l������w86M�fN���<��D�gf	�[�������O}8��̛��49�t�ryN�c�
ټ�����0��]��5�+�%qӾ�j�=����N�եԾ������x��g�I���+���db�����a�}>�� �.�����]d�o�>�+Z�����5�7tz��SB������=/,K�|k����.���;z�$���l���f,���؁�F�=Vjj��\�3�mJ�>�LŨ��8-�;iZ��|�/>��OgJ�ɧs�����K�X+��*j�㨙����T>��xX|����g|a��Ԇ:���P�g�&)�uwk��Gr�^#�:�"S�̠�~Y�c4�bB�?��#��]I�Y��&3��G� t�W�pW�^f�5��vd󙵊�7�ݖu��Ҧ�7 �*����=mv�G,�^��b�Uw�g�3�z�� ��{}���R�ɷL�C��՜8V��հ"�YTҮ�{��.��u��FZʚ�=ì1,(9ֺҼ#��)bdS����y���ttR��(�-�Zj�AXh^� �+��+����u;�J�^�����d�jڒ]tG@��T��!�����U����-��tH�b�,�-8=�D�]�ї�2N�qo_1ۧa�{
�j���z��Rw%�Z�m��I�p��"7P����)L����>ռ�k�)�������sn�S�뷘��Y�!bQ�si�!L�c�3bҙ���qm�D~�{dvQ��z*/��1�NŃj��>�i|� )���S��
�E����$G,���$����j�%z���+5�����]v�b@������dc�*�`�;��m:s.-�R��jE�FA�'U�1�5]�2�kv�]
%�R&�_`��M�kGn�,�#�%cDC��s�辑�!j�����`vka��S�ݬ{�0����֡(;"n9� !U�]��V�;�bZ��;��K�������*��w3��+���������'Z���'j�7�3��	3��-©N�vz�ͫ�̽���1�Y� ؤ%6��8��	گ1�'�
o�pU��1��/�.�t-D9���Z������!��^J��e�2i���-ִ�j;���`��������5ك8#��0��[���`t��~C�J\��,
�(��d	:���pG{v>��&鼴�ɘ��G�N��Ð�󊍣�wy����#��Sc�u�+� M��)�__u�J���\_S[T�)�����L.�J\a��㬋,���t�͔��}��᧓�����TQs!�#�����N��N\jtȋt�Ɯ�y&�:���=Wo��y�k!7�<w(��oy�hg�|��2.s��:������S���A%�n�ut�Q���ob.��qχM�VJ=�b�}�+Y�8\��*X�f�@B�u:�\�jj�I'�Qq�8�]��1��6�������������l�Jє��pe)Ǝ;V�PԌ��b��k�b��(����f��䷶�+��B���ҏ��wg�`D:�+_���	f���R�u��r�z0�\�Ep�9��t;�����=y�bvʱ�Ӷd�&r�jB����(��ZVE�`͝Q��f��}�mc%��Pڊ^2ɸb�g��d\��iו�_$Ds؇�2�Ɯ���rQ�:�{�uꓨel
 t+�ig�Ѿ*�X#M�D�"Ey+��mݹ��<6\���4&^�Op�a�n�%��Cʂ��0���S���ژʼ�LT).|�,Ôrp
s����F>���ǟp�M+B��6�mn��D��؅$�mH8Z쓪ܲ���WD����*db��5k6�Ν9��+[\ڊ]��o8��t��Y���27+u��$��9�N���QvK��n�-}bb��2-�C��|��|V$���y�N�u�����b���b�^�)�O �v)�2�#E%��|Bmڛ�\��#wK-|�6��,+n��h;��j<���]-�/������1[��Y8����P�.Z�k��╌���qx rX�u�Gt	`Si��G�Z;��]Z�<�k��!��][�7�^k�żv���[�e�;-�܇	��y��^䮶����=*���z���[K�uEMX�z�0d���h _Bx��d��HY/ES�3���b�Ո�ϻ{"�%���7gZ1h�����g��_�0uqy���/,��h"�JL�N�������H!�+�۷ݏ:�~mȚ
��Q8<R�.�,L'��r�ǹn����c�]��,�av�>�kv�+�
yeanr�j�k�9%Y�\y�zY��u֦��Mܹ�5���r+I:G��pZ��ӍƱ�:Tg���� ��*�c��nA��|�1���fF��X��[���"����P�����x3kz�հ��Fݧ7z�����ܙ�7X���jU�)8�EHw]�G"]ҝG��Az�=�0_VĞ_�%��)�2�Ғ:�䆣J �����SC��[���7����4`u�����ݗ#.N��ջ7�$�EԴc�&oN����}yc3��70�T�(�r�t1xn���.�ʺRww{WEk��m�Q��xn��G�ہfa�@�O�u򡚎7���vo�����e: �6�����6���k<pc[�(坋���w-L�)6����n�WRVv]�Q6����5�e|�LB*�w�:�)!�M�N�<INˮg2U�=g�R�J��IB7�I�`��p؉������WY�L`��ع>rp���rД7}��q�Թq�ys�q��X�-����U=,��sGv��̼�MOb�'���j����^D���5��|��vvz�7.Pѵ<�Ad�"�8]Zpm����Gt2�K��JPd����V�қx�G�SF��>���;YSޓ�NT�ϯv�F�A��|�[���w�< ���4���T5qi*X�ź亮��̗�hv���)�����6�v�Ɖ���z���Pٞ�VPw*��yz���xKm@���|�5�9ssG���kI����H��	��eoV����)����]ۖA��vm2��3�x�s�mUt4���W�E2�Y@D�]*]`��J�=ɏ ���T�ЩYm�7Vċ�0uHP����5�n.,��[��b�q�n(������=�v:�L(ޖ1{s�b♒{�>���&�����y���eG/x1�8/1�I5���%��>�?�2��l��`���y�;,Ōp�Ҋ�$�` ޫ������c��Io�+a��E��dV����jxWh+m'���1��S�����k�W��F<����O(���˾�dK���_�%�M��ώ6f�O!��`l�/L�`���n�O��n����g"0
.4�{BT]
��ʬ�k�뗘PS���hg	�r>�N��>����C�0�9��2{��`$�*�lvT�8Qg���^�M���y��p)�U��K[w��W!Jn�dk*'�`�̴y��� �����糯�{��+w�ݰ���J��8�U�Y��w]�A.�[T��6�Mڥ��v�-噈�D�	��3+1��>u�YԵ�MPOgB.�e�1�p�˴��j�C�A�'���F?�À����Ct	r:t�-�y�S�V,�E�ʹ&]	��rIZ#��W(6�m<h���cE9sQ4�,�?^޻��[����w9�J}2vWφTG�8���=����mZU�HL4�u���&�Ηw��Q��z�)�u�J�0�j"�;�mM�L<�H0\�s5c����ه<�}���������|�����e/�������U�:��2��U�H�9|n�	1��<֭�+�Yv��h�N��gk���N<�*�y�Y��b���ԝk
e�kY�ޫ��?�<S��S�4��}V\"w�ݺ�z�:�4?p�z�����ү��چ��}�6"K9v��1��|o9,�����?�&�=��0L��;��B�
�IZJ'
BP��sJսDN���r�Z����1�Ůu˞h�Vi=��q�ݱ
�9(�D9n���Q{ԓY�B��#" ��}�J;�f��ꩪR�$''PZ����{�����aQ��ۙ�T6Q�ҵ��g	�Y[}�n��sМ�Ftj?�티(N�txz��}�p�+m�e�(R�\d�yudrF��3�� yh}M�u�����,�Y:����ږvg0o����VI���9������j��vA&r�3ސw������r���TKDa�k�6|.�m��T��40�-T��Ǵ��J�E��!���p�3��.���ږm�V�sM�"k�qXZy�sh�<B	�tl���o�e�STƲ�^����\�X4<��a�D�B�h�R�,Cpq�O��V�x�D�B\*:۳���uxu�uL[�1�l�������pb��$~�m6k��t�[Qq�PlU,4��QNs캯����ܦP�`f4Q�
v�D`A��	EbLD$m�tCd� �I�\hr�E.\1��c�Ƥ�!�h�"CQ%���t�E.�sF�r�6f�$TT �m�̌gwM]�P�';$hJ)�Rc5"&�Ѡ�\Ѵ@DE� �DȣiI����9��6$�QD�F�1���b5&e����6F����I��I�")��b5�wWM�A"���APE�RY����w:&Q�D�0�@hfō3%2 �L�M�cXf �fN�6" �h�1�P�c)���o����~�z{w�ꎴ��7�6�R-�[]AF�8f��k����p��b����fܸ�s��92km�|`��ε�U2�D�Q~X��9g vdz�����t\�ς��������xQ6|�\u�G
�K���� Z*@-u TL��ps���D:���MDiZ_&,p'Xŋ���L�=�\���1�ǋ��-Dg�`Uo��:���X ���o�ur��}�����t%���Q�[9�^;5�BS��pW4���(	����୬ž����%sg����v�k<l�+՚����b�^�˪uW���Nhl���'_��Oa#�49A�@i�r����Z쪡K#���,X�8q ��(	��D
�������_`�����}����+W9�k��UbޓdY����#�Nф ��6�5,r3����M뛁��-0�+�}���4�@���蕛<�Y��g��y>uP�����!/5���.z�i�x���&5E���cx���7���bU� (P=�� �zWKK��k�ʽ��q{Z�[4⎎�Ұ�39G_��Vm�L�:�VMK��㲯̇��\(�LM9�=�՗���r(�4t�z.ge��Il� ѫ��1�Z�5n��L�=�s'�HA*]��ӿ'��'|��<�igiv܆����"}|��.Ė��*\��4�:Y)��P5�@�o	{8%:s��Di^qWv����=�A���4X����x�~�'����*N��L�yWǣe3�������V�����b;!ĺ4WP��g��z^��x��`I� 8����l��6:W_ִKӹ`n������Rs�2b���שƈ�,���UH�R�QcCw��.�Bs�������&�t�lU�ͨ����&ѐ�Y�w��ǍAU�i���]�n��9w���jʨl��?��w����^��R(�h+��Q캑H�RE5A�/�a[ ����V=aP����o,g2��q��՝M+�v��ؔ�ț g�ޒ)�TH��l��#(�u����n��4R��4�U��p4[�B��r�nc ���Sp cYNH
Lp͙�ڥwQ�W_R�2�w��@�	�Cd��TF�3���\�BN�1F����B:o�����V��Wީ����j��9>�V���V���倧J�x-��ħ��د��Yd^�*(���]0o�;bK7q�q�����6��Ɍ9;H"Yb�*�`(t�����1�6P��CJ�}���X�[q�.���z���fQ�����t@BaEWP��_;z{Q0�ކWz�a�\������{�3^��U�e�L����^�R���c�z��Qҩu[�g %"�M��X��9'k�=��Y�������&��Zv8�������YӮ�=�c��܁���6�;	[$^�V�u�K���K�X�\h��S���by��a��zxc"���&ݻ����*ʑ�q��`���vzZY�O���������(�!qg���p+�s�EE��5���d��W]���Z�E[��=.����b|���/0S��,�0ifz_L�Z��?.��Ƨ��.۞?\F!0��ȷ������F�������S^âɮᾼ}g��R�=���r��ʮ� ��W�ze�,X�{�g�o��e�J^U]�|��s�S�Q�ɟ�VSw��P�1��h�F�4���m�g�eCvJ, NÙ`q��?D{�Moys�u�]T� 4�����]��5&T~4%�,z��t�S�8*-ڴ2ʉ
��	#�H���CY��@ڛ�q�g���ԗ�q�q/����B�yU8{!�%��E��4k�6;r��z��v�E��x6I��]H�7�c;;�.pS�mheOR��Kf!s˸���N���L0�f�h 8�Ӻ�"9Ps(� �W��Nu��b[p^BE��7�Yc���9Й_�2�zV��#ěx�xl]w�]��� �ښ���6��ٗ��+A��{e�Ӝ��]���h;;0�}E����Z�Jo�a������gd_��͓�Q"����P�C�j�J]	����e��A��@����M�j;C�V�#��G]��xOʟ����
��c�8k1B�t�)J����0�3J�8u��V�8@�X�cbK�f�û�P�3iɭ1���g����+�MÙ;��⒳�ՠ
�+��*�Y��]��:�ˤ�Y���ãPy�of���3��jZ�p����&R����" ���	Mo3���Ad7tx޹�p8YyLgF�P�w_�Ӄy"��$�@2�o͗ŀ�b;��01Kޓ��)x��a��2�^@V�\�JrC:��O ����/U1|@����O���Jl6c!����5�ó��(�T%�SՋ3�uӵ���9��L`�q3|:�3��9F̄3C�g�)�2��u��4�=�����v�T7��gQў�-�!�:WՏ<�#x���3�t�Ӈ�df��Dn`�}s�T�86�kFW�ق���[*��}+��L�"��'�/�؂rJމ�z�j��<�4$6g�v6�;ud(Wnvj�Eg7X��L��d�*�ؠH���w]�&�_��M�m�pm-��P�q�-�С٭�|��׮#N�9a�X���Y�u���|fG3v����PK0���Q�v%咕�O�6�$Ҿ�K{tuV�?��zs���,1�zxY�k��k"�g��쿩�#�s�N�)�O�o�P�7�҉f
�(`|�$aCAWq��0L7,C��N���):��(���K�ү�-�:��"{�xr�*atE�|�
����*_#:.��Rr��Q��h�e��Q����YJ�����J�w����Pu�d ��P�uCw�)ӥ��q����9�m����� _�� g�];
��y�ꉯ�Tp��g��u9����i���[Q/zʺ gt`{�z0"_p܇���\dzj��s�F��Ք-�n��}�^ẃY����@�<��Z`�k���1��٬�Ѥ��Ӟcז�#��ǡ��$Y�YѵB��0Q��⎖�l{k��O�m�^k�h�^b��)b�QWp��A��)CDV��f���m��Z�f�Tgg����y"�OU�Cѝ�3�x#Sr��`�J�C�7���`�8�p�4� f���u mF<�����#�5g47��w;��v�m���Z�:)ӯ��Lhw�<�W�wކ����י��.왈xh�Hc���wo)[����fB����=�r�ͮ�3ye�YWư�Y����+(Ū�37+yVO�A���e���&��.��<�tAwޜ��UNZ�~|��|r%�çg�,GS��� �Q��1��Sl����T��j]��j�`j� n���!"�4OҚ5�K�zz��n���
��=Cxρ�U�� �_kND��)W �&ב(Fi���=mi�U�480@w>n �g�u���c`@��vM\�J�/j_)���.�2�Zr5�Gf���u��l�(�D�HA��f��3���K6�[���3s�?�gQ�q�1�_ګ�_i���C;�ۗ��Uj���a��]kb��f�,i��A5; y&� 	��<�p�~V8J��쁶^�ȇ#7nቼȐLe5�A�{�P ��)��q����<��
RY��T.���t���vS9:����y�%�QP�/J���+�ƶ��U��2�.�� w�X��M���F��}�&.��{;�,����-����.I��tE��2�q���_�HOt̓=l����a`!�3*����v�!�f�rr%���H�0x ��wLF�\���pq���� E�N_���$�x�t��aֹ��	�З��:�t�V�:�V�g�8ìäi�0%����֞�ϙ�R��o(��k�tC�ކ��w���|�
X$�����.�.ŗ�gY������^^i��u≂���Sv�z�֛6�ޗ\w�(J`os-(ڄ�M��{N�<2��T>R��~x^�wC����j� >,V�B���CG{���S���#j0+(l��`b��,e}4J�K��I�f-LŇh�@��랋�[xӌ�{����x�W���,ץ��〬U��V���H�
���=���L�ОjT&+,E���g�[�<���+>��W��x9�@�c�쥆2����3��"������]������R8i� 6̬��Z�CK=�K�A5\��~r3��F?�h	�+%�3�?h��s���/h��#t�����(>�1F��1�1%��޾�)�hW����\	��\��س��ο�^T�\ey۰w<��.e<���R�o�P�d�;�+�Ȏ�����=T���v8����R}s��O;c��,�d�gs=�a��< �|���5�xY5�*�HsȍW��0_�z��w,uM�k��z�㧳�r��H*$1���Ғ�B͉��J���<����1���UG��u�ö��X�K���_P����x�����][+�z���1�r՟vz�;��aaAa#�}�z|c��ڔ=k뒆�[�X��:E¦������1�=p��/>瞺���5X�gtћ��8����Ft���X�ݻ��'^�.8��n.O*K� ��]���.�njYY*zql���Sۊ�4�ω)d���������V}P��h���0_M�=(�S�󌞤�2$^b�u0�/*$+� $n����L�_!�C�����#��Y��7\+����71��{'
��rL�(3��A�\��l�ڼ���ۃ =�1����.0�l�q
c�LZ��T���)wwQ�4�s�.�|��������b�Y��_[��BiS�t����̰��,|��-�G��$��c��:�M��7M�{SHJ�.YT=��>Ֆ��켬'�g$�}�s�����Gf,UK�w�x��S�%sK3��k�s�P���h �rģjX��5X���]�NMF��ra2��ӆ/�����ڋ���Z}�U(ޔ ��V�L�ߣމ��/��u5_�Jj8�����������TE��A쮸��L� _ڥ���7~�x��@R���U�[�g��:M��5tߐٙ�7�'/Ub��ϯ�j�3�����O��s���?�Ȍ�[.B�̬隮�C��g�k�̈ਃ��b��wSEo��c�PHb/؍˫�%��"�������x�g�l�I�T�!I��(���\+ֲ�C���3���7Ț�ڝ��d�$�P�[�)��{�fCX���\��.���=����C�p���@�q�!��Ɛ�N�d3�T&�8<��� [sx�.�y�Cډ_a2a�Γ�6�AZүiuCY��W�*���x�����wmz�x.���f>Wl�̿8���:7ٹ>�>��z6��M� �?���:�H�/藆��j_f��F����kyi�x_>�f;5�鰛ڡ	��Ώ=y ����_3�优~�`���/B=��tM1r/U��ϰ��D1�m�b)M;b���(���"�A}@v[hL��F�=%���`���,��Z�9���0=�n�1��U�pj1����l�(I�+����'mFӮ �kP	<[�fG��:\�q��^��J�ok�����t�"g���!=��J5l��W���UH��t> .1pj;������TC<4�0'C��q&�Ѕ(5j�����5�*�uB��.${�Ӱ�S�y�ɯ�AW
Y�,ạѵ=����}	��[v_��)! sw@uӪ���m�_1����a�>ӵ:���Z3=cmE �s�����ڞ�!Y�����]IV�\�vU���Yt[Ԯ���8W_iݐ��Y�\2�..���eCʊ�0�wk��Ny�B��v�-.g��˃Os8p�J�_h	@���3��`龄{P�_�4�+��VyA�wb�c���N������3��}L��R�p�ЈPjv@���y8q9�������T���n��,!�V��F�m�'�C����O'��u�̽�fk�<�?\v�b�8��������.K�
�V\�(�/�����U��3W�8�GA��@NӸb�Q���T�N38f��p���:\�CP<�c�[V��Џk�� t����J:i+y�3�@�9�'�q���]�m�LVW�8y���Y[���o�?�Cb��O=� _���`��H�O(���l^�{���l�Ղ��<~�׏�����.�y�é+d5~6:��Z�#���O�iIă�A�#-m ��pN�X��_7(h�eh��hp�G��o��
g�s^�r�Dú�j7]8�j���Z~q�59�CD2��2��1���1�	�z��DR7+)1n��wA�l#Y�ٱ�NX��*�Qb�왎�U��8�gB:�q���/�sg҆CZ+��Ԯ��猤���	0�,�dUXS5�̪ȍ�"b��B�W_�D�;�� ����}�ӭ�]����@&�ά�9R���'��Hǅ�{3�[�x9�����3oA���i�V�MG-әH�a��:�u�n،JDkhզ�[8
�m��p~���ׅs�u����<��P� �J��C���eX�t��Ϲd�]�)4e'���Ĩ�s�.�#7�)4]N���N��N�Z�A�.b���ж� /84x����$�]�ﳷP�r�Z*���]��Ք��_%�\��'�7�e�S��z��,Jcq��~�����o�~�2&x�z<�*w@ 8�U�y�{����ą�N����D�}�K����z��3a�h�L+��o%
��܉G{�WO�H�;/j��+;V�,���e�S\���=:�k�Ft@���,� �;Vچ��xz?��/y�x�Z�H̹��Z���%���r$�_>�XV��oTs�n���ا����*�[�v֬�b��f�#_�uos�c>am�(3�_�uJ3�G�N1��5�-�t\w�~SKΜ���.�1?�놾iw�i�g�ZZۗK�
�_ L\-�ض��e�s�wo�q`�BΕZTԦ�n��h��ovF5,|NRB��@�9��78q[��R��q��k���g[̭|g�8�������'GT��8VBi�4���D����d	{�T�L�tp��sF�U�p=�g�4��}K��^[�Es�3wxӤi��R�^���o����1�m]���Uz���� YƏf�1��3T��q��ڵ�#P���OP�v�h�N�F�F�}7%b�]/P��N�o��i,��Uh0��т��N�Uv_2:��ġ�\yU�xC�m�q �r�͕���m���]R
�Θ���n\Vɮ�o+�����7�{��h�;��Y��>JGN;����__;��K:�u��؍i}d)��z07J���Dm^��w�i�u�z�o�@��g�����c���b��ư�	���Z[;'q-�{0ϳ|U�I
�9[�g��7��<_
[~�/����C��j���R돀��$]�{k�K���‐�8�
r�m}�FZ_=Թ+"�}9H�7`N�sf�A�XNM��`d�,��w�vPd�8[���@r�m��:{s��G�'���9���z�g�ϧ�V�Q�O���w��ξ�C9Z�,��ۦ�K��*������qa�:{\ߓCM&�d��u������ ���N�:�Z�!�a����<��\�>Q���w���`+���:�-��{�}s���B�M���v��Lz��]�np���7`�Ҡ��P�v��N�U&sBE{ڰWe�Fa�б�v�ק�EH3[��IX�f�=u�W�e6�S�3�4so���􈫎Ȓ���x;cp4n��t�;$��76�6������;���8*���/q�G��Wӆhc�=�}�8��r�D��"e�Y}���;����a��(�<.ڝSsi�U�Ï���Ko8�Jf^�7:b��UA�'��H�%Ih�*&ar�4a*@��JHA�.��F"w]�d�M T]�)��#9Ѩ����0����wr2iH��HXa�1b�L�˘�JlQL�&2np���Hr�(1��L&Q�aE&�@�#h�M�L�
"2JH�C&��4�&�e&LE1`�i�f&(�#5��1��B�&�%��H
R)�,�`�*Lh�Q�FW-��I�Wa�I`�1�H�V�܍��wRDi#h؍��r(�JB�V)�(�"� >� 
����P���L]Ks��� jƨ=!���+��+���X�*��{֫賽��L>�Y3���A/`�YӇ����=���LϮ|���n/KAz�~6�o���o^>��/�G+��^�]zU�sW㞵篍�^�r�~-¿Z��_���KO���z�;�߫r��������ߏ��o
*����zv���� :a=�o��T8� /��W��[����s{mޯ���5zo-��}��_^^���_�<k��<
�{��G�_����ڼ<�s�z�{⾯ƿ�����|W���{{�6#� ���V��W~�5����ńg���xW���W�μ���xm�����ߪ��������\��[p�}���KyW5��>uϞ{W�s}��ʹ_W�Ʈ��?|�m�E|]�ۗ��j5�E"+��x}#G�Nطޙ��u��5s�<MB>�#��H���$}�>�#�����r����W��+��w��^}{꾯
�yk���m�������w��6����ߚ����7��no;���[���ϫӣ�DG� |+=��78�ۛ��?=�}���_��6?W/m���ߋ~���_���Fܯ�s�_�ݽw^���Z�������}^V�w�>|�K}~�������^������ߚ���4E��c��DH�� �RΘ�i�����|�/ϵx��/k�y���W-�{o#~-ʿW�_�s���������^��������s�o�<���
��{����Mx}~-�����W-��}n�Q � D�q�ҥ8��&i��CJ;�D�z$G�"G�7�� �M}ok½�z��7�~�z��-����yW���G�����F���xW��������^U��ث�澵��xzU�}W/_߾7��<��^�3��c���=4��r,/����"���/�߿�yo-�E|]�}������}7��
��W
�U�����#���}��y����Z7տ^�{^��������y[ڹo^��>5�^����ޕ|A|G�G^FH�E|;���^�wkR�p��*�\���~w�~�n[����-�\�6����_�xU�r�������߭����o��xm��6��/+r���w���q��߂�=���ϼ�|~����CMlo�Йɯx����\HￃR[��x}ߝ���Q�����}W�\���׏�7�}W�\���<zZ
�k����+�-U��}��^�[�z��|{^��n~���>��W/
�[��
ߙ��+�
�>�F���ڏ]x���z�������&�g������t�M/)u��8�P���>[Ӱ�S���|/ޤ$U�T�w%�+��b!K�Y���]�0:a�!��@�Z��0���Ëtt�Uծ�N��.�˴+��/&�`��/��N���:37.�9�^T�_�����*��߯��3�; ��]�U���h����o+��x���-Z����|_�G*���ǧ��W��}[Љ���>���"3�#} }�G/ʼ/�xj����<��(�_V𖲟cc�ޘ��{5@����DX��B��m�^;^V�����oϝ[���_������6�����|m�m���W�߭�}�����\M�p��G�tNj�[�������Z��-w�y[�^�����m�xo����Uz\ۛώ߯�xU�r������|[���;ʼ��\�_Z����ίkxU�w�x�6���ۛ��|Ĉ�z\Nv��m�cH��qG�D��{ݛq���DF����}����ѿ�����_��W��+��[��~y���Q�Ǟ�/����+���������h��]ﯪ�11�L�o�S��g7!�5
)$�T�������?|n^U�n~�ֽ�?�_��b�B>9^ۏ��}�G�+kﮜ��"�/u�Ǌ��><���ϋ�|m˖��?5�xZ?ώ�/����zW���>���1���n�]&Rكc�>�Q_V��^[�������-�����+�����v���(߯�x����^V��^����?~*���/{^W�\���^�x���s�����[����������>���D�6zŞ@@�;�s�����~|�����w����=}��W�}k��^�ο����o�����~�o��xj��~���r����U�����a}���0DE#���C�,G�"!�+�_|�"���kY����>��������⼭�\�^ז��ux[¯>����\ߍ��^;o���m��7vž+�Z�_������߾~x��m��+G���y�{m��m��yW����Q����Ʊ@""|�n��KS(]�5�������J��+®\���lyo��^��y��ѯk���:��i�׏��k��V����yWչ��W��^U|\�j�x���r�U�7���o_���k����|G����Fz�{({��O�}z2��u㛯D�|D!��P�@�=y���~-ߗ���|W������/KF��m�~��_��-��k�yW��^�^�^�[ʿW�__X�9\�>����>:i���srz7�����t|�j�4�1�5���:1�w�k5�P��>`y�[�+yV��(�,�q��H��*ס��}3G:�,Zo�h.�X���jfU���E#/�����K����`��U�
+o�~���a_6����>� h������W���|�����כ��nW�}^��j��ە�}�澮��|o]���U�ݷ��{����oڿ��h�7�����W�ᷭ������DnШؕC�ĭ��ք��!^���kʼ/���^���U�s^�yo-��o
�/�|�ۛ��[�o�|�ҽ-�\��w���ܷ�\��\ޚ�����W���oׇ���ϝE�������F���"�����`WR}��s�p���}�3>��G�}�G�P���������-V��߾//J�_�W.�|���xo�x_��<[�堯?~�yץ�_������v�+��b>7=1�|F���uX�N/��t�R){�DB�"p��@�{;�{m޻�W�羾���W��ʿ7�[�|m˚�|����������׵�yZ9�~�^_[�_��~��KF�~-|ERV)
������9R���ڟ�0��m�b}�>��!�z+g礼�����_���W��~/?�y^��xU�s��}k�����{��^Z���k�^U�nW�{~�w�Ʈnm�7��7�~>?}��>�zc�����ng�c6��UݓK(�����~��D���.����xZ/�~<{[��������^5�m�r���=��>u^׏Y���ׅ_7��׆�����o}��-��o��^�#�"�����g�}#�5R��řݤ����"��p���}��^�|\��|��F�ߊ����ߝ�z~�r����m�ͽ|��o���s~6����ޖ�R^=u~�����7�� ��!��eLP�#�����"];�s%ġ1�o<�$i�DG�P� �ϋ��_��~_>��/��ׁ�����ү����>y���m�W����ߊ�E�~^���M�z7��=+��������z�7�n\����z��Ū�q��̌<�P��Fb�U�1�`����w��{o�|^W�~~���~-1�P�b#DH�����%׫���x������mV�۱#���er�P�Gq7X}s6b�
PX��9�H�CAWqφ��0ۨw:��AL#m��3��m.=�w��w���Ú�G�Fr7O5��V�q�ׇz�;ַJ(>Y��;Nq\����r��w��"�s*�|%W3w;}z��f!�F	Y��u�Q3ƒ��.>M�ǟ=�v�i��#R��磌�i�都�!��D�_�n���tyW���m_u����B�jx�{3#r�Xz�VBi�r|�R�K����kʮ���}�U#I�����_����:WSǚ=u�C�=t�R���8稽z�� ����t"�T��{�����jP��[
�
��B��w����Eܣ��m��f ��x��s��2 ,ù,}�^���3^�[�jc[�����W�$���P-�\�zgw�u�T#`	�������1/�6͚ru��t�EfL��.Qfw�N1W	��4��ѧ�ҡ_Ol�f*;�<S��]�T�SbRk�ㅱp�v�j`昞zue��^x:����U��8
�|��p��3�b�vo��ˋ�Ň$��ŉ�ͩ���7~��C+
�w����-O�7�< �ʚe��QT(��w�fƗn|E�y����e/!g���Z��Z�p{��W�Y�٤n. �JxI�B�9(/����ޚ)���b}���މa��y�éc+o��?���p%�erSУ&�P8�tu
[;-21�^]v=���*j�=�yv����u[�pڱ�tFƤ��Ev-.d��+�hy��yYt�rق'͸n=�p�z,u
Û~�[��᳼����?{��^lz\}.x[t�
��җ.ob�on���}U_y\Œ51�,���G�*���L ���/�yp�3�֙_^v�8]g��r2FN���[w6�"d��?�e���>Szd$C.��')��~��*�1�	�i{E���4J�wL�>� QݗCԓS^�E�xJ��G�s����K;����J��%�q�*����(GgD�*vEU�Fx�*�m!Np!t���h��TO-�Q����H��j���1Ҿ�C����`��|\�r�5��s�h���`��0Y�^������'m�p�K/�n��bQ����v�C�;5[أ(F��l��n�^S��ry�k�_W�a?��f�����4EC˩D����gD�s��/s�,�±U�G�~7Ԧ�ï�_ӄ�5ϫ�PD�.K�����:��HG@��@f�uuz��]��=�'�?������cu�rC+��¸J���6zT��H��r-c��c���CnX� 8�6�hGd��ՎE��X|-֦OZQ���߇���e�Z�;2�PN�����L��.6�fܧs��>�����h�5,�J�R1��� �o��DF�A���D�ǖ�&�4ŷf�r�b�:,vQ�j�7�	�0K���V��5RerƜ���(���i�xBI�rg*R�7yi-z>�������ݚ�����\Q���q.Z=�'s�Z�k���U���W[���uR��Ȟ�fL�{nݨ1�f�����HW�W��H�y�9){e{���~+���.�V+�%nw`�=wU$ ��c��p���a�L��9�T˸����ǵ+��.$F殴B�(D_T��P[,c#>ULG��.&����:2	����U<WB�J\(m�ÖN)��i�;ȍWk�s�F�^����^T��E����8�SJ�*B�f�������d�*�qɗ�g*�q�u6~�[6�X|q�۽�������*.G-��^پ?J�<+���>k<xJ����u�/��g��WZ�&'u����
�W+*�A����C��p@
*ctiL\��%/���yoV�
Ю�Y�������z�\1�w)��(`V�.�5'��s 5 0�>���U`�.͢�1�)�5�vv��P���������>�#Qz��v������#���j����y����9�s�W�HOy��W1'o&	n��"�:��Ι��^�o!L�S]�{��m��{8w���6��([�O!����!��RQ��2��K3mD��s*�3]b<^6M^��-�ϲ�絃�3l9S�ƪ�(�'�o��L*>��S_�&��}�}�}+w�oL�P�',�h�5�_��s:na0���!�1	�۳ᶚN��|�'��C�Pz���6�a5���Oa���:Ī�S �gT���WV&��1KqG}���t�"�@J�H��f��14��Eb�7`�bׯ�s���ܼ�I�q#:���Qz�*�:W���_���_�:��u�*���h��¼�>%3�v+��,QÝ{v�C�2&�,1#�H\)���e�F�7;�5X��څq�NM�D˙����y����WG8���7Oe�њ����Zy��8�3��R�)K	�r�Je���A:+���skxg�xx����yץn'�@��3�Ti���4s�r	��15<_l�8Ҟ@F@��m�����	���F���U\�P�^�T8��w��d�nhA�s�5w^t=��t����T�����(K�������O��Ӹ�@��,Xj����s嶇dG=�F%Y�{�5V6U%]e�g�&�s����6d!�P=�!�+X�cV9;��Q ����g�"��sZ�v&י6�&"Ū�-�?3���ԡ�9��W��.��ݝ�ر��Q������	ð&�w>��P��+n��a}�i�Kg&)�|�[�����B %����uJƭIV�>Y����ꯧe���*]N�n�>un}Iގŵ�
{¸v.�JlH��\M}+]B r;�(0"Y�auӐ�Qw�:ˍ�B+K��7)��RƎ�U���*";�+`��L� ���6.w�,L[���7%i�ss��qT���D1�m�b+�[��4�d.�"���h�{B���[=���s ��~�Ѝk�!�ƶ���Tw��Щ�F2t�7`mL:G�*�f����w��R���<�� FD��3�r ��.�P���QA��C{\T�ӓ��a��P�d�!?��LE'.L+�4��V*Z;n�BêG������<=0:��k�D0�yj�F�w�u�m�
�RW�3"E|.zb+��572>��K�t�0�cYӔ��S��w�+�{�^�y�0���Bh��-�g!NSl�����5��r "����6���*9���wis*jK������Ŏ��{�V�N�l��gl�)�9鬛�#E���$��:�@Iѣ,��\�3Q���5���?v�,Ƨp��c��l��v����Wm0��&7(э�j�Τ%,Y����˺���Sv��I���GwC]E������jp��!��3jc5b�c�x�d�D2�Lł�ק5���-̗�s�M�ȇ�]2Ž��%�ZC�Y�o��Ղ��]\y��n��I2�4)�T�!��������k"��|]�'�E��'e�80;8�g��@M&|�֪cڭ�;|&f��a+�gͯ^([����+��۝�2!��G�,�u�f`�u|�(�� �> `w@�z��خ��3�Ԇ�jW~sh[��~�w��f�y��*�e��϶��4�aVƃ�D�N���f�7 b��1��"�aֈ��_
����n�l�:�3ÝU��+؃z��5W~���J�(�.4�͂��@Mr�A�D����CEƼ��&Q���f�EEv�w���a�%p��_ѓ:~�(r7d%rYvm5A��c���1X��K.4��ݶ�!owUL7�%Kr�_�{\ �$�UMf���<%�Z=+9�ΰ��x�wM�/� �.ޒ˛�ʯ�\_K�88F�'���쪰(� OeR�B)�oJ��w�V��!�ᜭ]�Y.	�8�1Żya��g4l�P�����w0T�Z<���9~���#jZ]�F$Hr���ġ��� `bQ��'Nn����f�Ⱥ�����,��u�+!^�yv����̝�l�^�F`V�<�E���K�٪�na�V�V��ݼ��譧=��r�t��4��]���4˄XO��Qǖ�D���	oc�+������v���$����������tw���y��e V�C�n�*�$�;�}_}UUU�N�[S��3!y��=ݕ��U�}�܈n��.�W��DZ����0��z�V��f�}��
����J����_��s����AL�=����;���r�jq�\��y�WwzC�$}tj��C��l�9�
�Q�&v�x�6	�ᨕ=��gg�q��pT�T��_ׯI׋&�\��z�[��#�8Xb���d�3��0*�i�94�޹q�7+�gF�~�᜸��=Gb\�{>���ʵ,�J�^��9`)Үsw�hh���NP���O��N�C��{ ߟ�5��g=y�M=�~��Z��>$f_h�ѹ��o8�6T����e�a��.�'��d�l�c9ĝ1E�6�]����:��~����{7�oPR�V���#�Ҡer�&(�l��LGY�~kk�ӽ�[���H����� ����j���lG�N��K9T��0ƈb�#u\
�\��Ϭ�in��W�I��Sku9���=�+4{�v�����@��~�SJ�ʫK�z�R���O>�@����U�^11�L�9�l��
,�	͹�,[��_�l\�8�Q�,���2�B�>��Պ.�D��+�T�۳��q�C����v�gc-��b��$���_�,Xm�t:K�Q��]GԪekxbs3��*f�MZd����ɽ�T�\��^���/�����εk�c�ʱö `� ��͔��*W-vA�/���T����ר�c�wS�vu-t�Rz��9"�]��X�tK�ޡ��K�����#�5��tU+^'=�s�SywP���;�m�w�%��T�w���zh�Cж�xR�P�9ԣå�o�Ec�|�H�wp
�%^��8^��*KWN�����k��c���=x5��B:.l���#k<�2�yOrh�Une��D�aT�Hfl�GP�@�OqG.ه�D�Sz����U��G�X�FN���M��i��!�s�*�qm�/;)pX�ęyK�k:�V�`�ۮU���G1�(���֔9Y�"�&j����)��ug���ߨT�3'B�f�0�q޿�˚������W	!�D&-�-���foc8���4��Ó|Y�Y�3����Ot�݌Y�:;���G�Jc�#�
O�	�p����ꜽdZ}Q�N��g+��t<���6�7Nb�ݥ	���zi�@�
cpq�巄[�l��U�i��yNi�r�����G]+��#�!�Hq�H�U�����Y�P0.��d��.�>]��rљ�[}5Ĥ�x�����N.�J��м�'��ё���˭��e�����د_T�L�����Y2�K��uv O��������٦z�����]b��Mmϊ�Q�Kw5iT"�_]I���7ċ�����nt�%4�Yȸ�s�((w��b�ݴh����w���j��D�����')贼i���1�ٚ6��e�t�pV7K6^��q�8W%�����4���,�r�u��]�]��y�fb�;�7_�V=��)�
�a�o�p������Z�6�����z��i���\��B��٨G�m=�Vt�=i��������+ҭ��'���t2𥳐��f�2z�� ,G��l�|ybos;]���i��x�Yt&���g��%���3M巸�2��WrU`�9�bb5gp@���z�V.��L���{�|3���t���T�[�y��1T���=Kv�8�]���.r.F��C�ݜ����p�_u��-���u�w|��a� R�Th<��%%F�X�V����D���]vG(�^^�ʵ�u���&h�([��x1"��ו�#�LgJ�nq��57�f��6��]�1� UL�)���y��Xx��)���v�=}FV��a�T��uZ]!�)!��4=�/X��n���o��8,���fƩwXҡǵ7Ɛ��A�P��"8u���˽,��VF�w�q4!��F ݧ��X4\�s�����~�TY- ��F1Y3��ŀɊ a�
IKF��J�
�h�(�!RREL�6�&(�I���c�L͠("�PA���S#!%�]ݓd�ƍwv+1sr*#����!4lh�b��ƍH%�J
 �E���J���wr`�H�l��K�	����#	6Lr�u�1HDd)cQ)`��(��QFJ2b��3%&h�j#T�2k˙�(�Ɉ�`��F�h6DB�0w���ioc��D��w�Z�&	Đ�Г�Z�ڮ䙳^��4�y;�ۓęz=�]�:J`Yr�1:�R�
?G���G�7���}.*&wO�7�=�Oү�W8N<�pMg�	V�u��s:��y�:��x��cU�zg:r7�h���T�ĆB��0�=1��Sq*b��PJT[�E�O��pnۋHbCz�����A�g]B��8w�D������:ʆ&稢���� �lI��꬜��-s��)�`m�a�{P����yS���ܑ͜��p멋��G^��E�c%���en� ـ�멑T�1c�������D·ų!����ܹ��D�)�=I��K���8?�bx=��2)L1�#�cj�p���G�r�ʧ%cǔR�^q��n�l�4�d�W�@q.%q�1,F�L�1Kf$db��r 2�1��iv؜穭�Z����We\�ڵ��E@7>��Ժ?)BV�}�o���Ǆ���Z.�
��fQ�Թ��=��������*������b��1R� �Ln��������|�=���η}�=q}��QUj�N��_ۭ�< ��uL<�Gjl�G�D�z���jUÍ|O�7��j�(�U����~t8c���-��E��j��L��H�·K��]4����2кwu�rg����N�B�Jڽ��D��Z%h�﷔�)`��e�V��vpU�n�Y�K�V���ts	�G�P�����@��.-fB�fz��}��}��%Ǻ{�������u\4�����7�*��W�ѭ/����j̗[�y�C��<��SƢ�U�v��u�֏	��ȱ�x��lM��#\�q@L*����^9����)a�T	ˡ�X�iw%*�_�p1\��t����\����i	�	ݍf� J�no�@�cM��4/5�Z;"�Ag*(Ų�=&,GTL��C��_Q�^���
֞I��7y�[�g E��ia�j���63~�����
�����>A�bS�*����p��
=��qʜ���3�3��#�K��LƧt�Uj�t7��,��%<){��]�������<��q虠=�1G��S7�*+@�n��別4���T��C�eˢ�u�N�D�pD���T܊�Q.�c�F:0����{���O�l�[�W�9�a��G��N3y���j�~G�5����@U��CR[�l�	-p�1�����t>nd۞�f���nӡGsJ��F�MS�/#]>�K�a��v�͡a���ω�5t8y}U�rC��蘬��K�%��8���')�;J���I�F�����	A��� ��^���ס�c��o�8`ʙ��,�,l�QJ���n����3�i��&z���0�V��jJ�]wy�ɻbs����V2�|t��!�0iB�?(`�*�{���| !I-�j����C�K�b/���V}�~��A�"�U�#ܶ� 7ڔ���dj暡���T�c���5,C��G-�E� �0�倲�PD!�_1��5���	��f�W@;D(�V��5�t�# ����i��l
a�j�su����n�`o����P��U�#�o�u�N�):�=�고V��b���:m��L9��Cf�m�g1F��b�2��i�qp�����Q`b+\�3YH	�i�1k��F�:nh����U�n)r I���t��O.l�8��?h����%Y�xJ�|�(��p`��Ê�9]�i͚G����b��Wڼ�������1�Y���l?d䩎�U
/j�*ݴ�jyJ/dW{k����Z �� L@�m�Y�w�+�r�{f����9n0���	�G[��}u����ʛ�������s6c+u�-A��w���
�1�N�Y2�<�v_O��t���D]�U -�C�p��a��(��%�f�9L�t(ۃX�r�n1܏�	��J��U��̲}c{�J|$�ޥ��$.�����sE�l*�B�v��%Mf+�����]Fr���C�ڢ���xR��`gp�V������3�5�-��ѹ|o�X�չ�nCo_[*K#)��M}x4�ԍ��q��ά*�>S+���}��G�Q/U��K�n
=��]DS7/)7��5;�U��V��X)��gX���
�Q���XoD��Ǘ.y&j��;�y�Q�0;m�j� �z�ܝ��J��X�+/5�k>Yh�u���W�;���8��yd¯�!#P\�˪m�`9ʴyje�r��+��V�:��q{q���Jt�p8 ��0
oZ�����G_CU}�U2��
3��Kw��k	m,���;����OջP��U��t�n����EB2�P�Pȸ����p�z��HN��1���Ub�V:������{]}]��7�j]q��6p��$��T.��y��! 3|@|VM�Q{$B��E�����\����_�K�aE�tw���~���Z�Х�3tW.H�1�nf�,ɋ~��6M|�b�K�IC�t�N�:L�HgbX�rb���0��[(�@_3���JNO�Z�k�֫�]Vt�2�����'B���+d�(1`�e����O���͊�����2}.��}p����@/��1�͸#f���r�*�����=�I6��4nL@�y��m��T��.	�����"�p�TT�qm*��u� BI��v�ɈV{Tt.k7�7<q��x�dᬹ������ܩ�۷�Z~�G��#uݙ�ҾW$�
�,@�G@2JSm��Z5/��G�}׽����*��{���m X����p���7^��lر��4����|�n��/I�Ǻ9��c-k���<S��U~/�=B�����,F���ˉ���#�s�l�V�2]�osӼɥ9������s��
4��J�ҹˣ�c8�غ�:RV%E�*�]o��S��cD6rnl��c�옠����d�⸑����	�ˎ���u�B�z��qs=7�vD�����̤~�3�|iu�u��q�)�9��-*��\7��S{0{�#�luN⎰�jQ��fX�q��.5~>�����ɇ�d�2�Eʫ�R��4���m�o��f��_�ԓ�Va6#��uB���-��k�89��7�=u(��@JC(`���\b���N�*�O8���X�0T�)U��	ퟷ�N�/����֋��H_�_TH\V�y�]���S)�4H��0��?+�B�vK�[�j��f4B�N�b�(��_e&�n1�&��&�@j�#�||pv�`�n�O�xX�ym���yV���K��U�Y:k�x�xAKų
�I���;�Υ��|��r�������ez&r��J�N���ʤ��ٰ޾�p���V�k�u�Nʈ�FgOS7�佮2��s8H����R�O��;�f�X1���G�g������4�L�זJ�Yt�蝙 ���[�{��#��q1��+dY�g�q���z���� O���3ʗ
�Y���.�[j�z����A�%6T����F��(F�UɸjCsrb��n�����Vjn�L��I�j��>��U\.�v�`����#��;���G���hJQ�	:�B�����	���(���`������9s��X���cɆ�Fve���=�h�s,;�����a�� ����*���]M~y:�_e�?VnT�iW������a���^���q�{��P�XÂ�i��z���Z��k���`R���P�m{'�^+�+̫�3�i�9*���-����n(���_[������˘�}�GW��$n��_lL!ssXP�s+���jCѨ�d(���t��Pg�( �M��87�����_a�V�����aY�E
��q���]�9�Jܗ��W�K��2�]�9�a��=8m��ϭ����AravRT�f�E{�[~�]u��/1I��<H�52�#�t�ZPv[)���c����]�Э��C�^��	]�)��Y��_!N�@(�^Z�=r.;���:�'5��
Y<�����;�8����Ͷ-m��S}b��v�]t.�QH�*�
���p��z7�WQ�7����v�uC�MŃ���t�]}�	TF�nd.��"���Ǐ��Zڋ2o!���U}���Yz�uӕT\���O��"b�s��I�+ʌ"]2�r^�����֕=��Q`�Ov���%qˬ��eH&HܕH
��84b�
E���n�0�S�s(E�}8�W+����B08�<!C���ӁwG9�Y>IN��8yW���꽯���=��9���NTl=��˝�q�b&�ta|<pN����Q=��Z�WG���2f���B_�������1CA�� �� �/�U׹r�@�bP�GϷ�#�%sҗR8�gf�#�D��rڴqNSo� +���)k���%Af�+��Yfo��p������N���(��<@�;��ͤ����#B�c��|�Z�[���G�x+�4\�s�/aN�p��κ�:�Cƕoz������~����%��{ޣV+�c�r��npA
I�lL�1�c,�ǅ:�,:��/��W�M������=w�Rq���f�U^�<3ٶ��58b����r~����'"�}l���Wz�].�f.�V3%�p>08q��m�~>�+6���A	`�ޖK�mc;3$�Z�03�(���'���P76�L{�H�}6>�lE�`P�A���Ll��@�Pޕ�͉��3;`M`P��Us/�д�]��1Ь.p�&p�XE#۝�;�}���u�|9�	�(��k���a����#!<5���=Xt��B���ns�cKג�8{Mu>��*U�4���5.#l�N�GGzބ%{0?�oYx2��:�b�ގ{g��b�>�ܖS�Mq[TY�f����c+]5ʡ9э�l�����<t�n�.�:%��j���)�
ˑ��ɱ`��n �l��ia��^�X��G���r�\u�ƌ��2'm�%c�HNP�5���GNϯ̇��\(�LMf��'�&8>�U|�L�pTS0�����Ӵ]�b�"��q�W�W�sF�a�G��ړڮ '�|y�>Z�(J�aX׺��R'fА���[���Ø[�P���*����5ʀ�"�E���������)�ˆ��8�&�#ˌ��WQ�����ġ�ƳH�N\�.�L�cG,�sn�1)�zT���W^�3��_11Y��\.�l�9ǀ��y�zF��҆� �6�z�_�D���ݻ!_�+�v���%@�;�	Xj#�W�V�!p�m�'%��s��ë�����\��,|�8�/�{�u�� *�S�[�ǁ^��ۍ��޶bU��U��]e�Q��T���٫���a�~<��!.DȜ/n�L�d�������{�۹o��žʹ{��~���_�����<�{�Md�Nd��0@�`��؋��"`+�}�K��:�����l�|�)�til��=�/5��ј�}|_Χ K�!;�"�hȓ�*�X�Qxb/��ǃ��VO�ѧ�T���*�Q6;1P���"b�؄r�
�xu�\�yf��4��\�y�6�ryH��:�ݮ5y��_�h�48g�3h�<�'���b�%K�L��z�o�OE�}��t�:r-6�(�3�O6r�=5�t�P�㋅��}�0�7�+�p7
���r� +fk�rt���B��v�ڋ}O�K�5Jyz�w�o?6%<�E����@�Oܖ���~�"�u.�/*#T���r�%�e�݅�n�q$$����O���&��ό�6���,,����e�P���D��t�tVc��_nF������g�l?�75���NfRW�Ç��.O�J{�;n��>�v���)�����Et-3O>�U�yá��t�m�V_m	si���="����.�z�PUۡB�[�]�(L'�����wcyr;]�1�VNp^E�2���e�U����n���Q�^a���x�d�5��똅R�C�΂f.��m����y����=�+��}��}�Ϸ�!^�����ڋ)��Q�wZ��q�ηm�	T<�j&�e�>�&�3��
Pi�ك�\ڛ��[��94��=NR*���r�����?�d��oV�P���s���]ܬ�����s�t$��ӼQвhw7�g��/���M���ٗ�N{u볚��Eͣ��[/a�6*��l;���_<�0�\�A�]L�=4.V��'�efs����֮Y]��.
/�����k 8xGo��	�V�Ls�v���X�3��:?M�BԘ����Qy��[�1�k2����3n���}���o��=��b�O�l>�܀�4ʽ^#1���}�]F�jn�6���>�X�>�/��Pp���yx�/'+�^c��qE�cy�zwAַ�٨]��*b��x.��ʈ.9h��(��+��^��&uJ�'��z�+�`��NY���-�ގ�l ��,�ɵ����Yuj�L���=��/}Չ��`ם_�PZ9�.� ��{�.���9m�z��h�ݐ����3D"�Y�W���K��&�`}��fL+�ر��ظ�7Cp��ߨۋi���Z��.=$��^�u�5�Y�l�j>�ƭ���wS{y��w)�ur���z���:SoҘ{R���N�Ļ���)�S���jM@�9+}$�W�Y������Cbl�t�}y���B�>�Y�Л����K	\�I�`3#�����}kC�@;4�D.�W1�[�l�䘬f����\�����8ێ� ���n�A�����/�����;h���V��uc��DM�rW�N�R-�X/j`�7ِ�U6�?`s�[�g1r�p�t.����E;�,f������2n풎+��;��m����ō(7h��Ŷ��ڂ���X��R
�#��7C����ͮ�ܶ�s�kd2���@q��%wm���@­�.ɔS�xSݵO@+�.x/@�:�k�\�BB�ŉ�B�ٷ.���Yؒ�ʗ;E5�����Mh�tX4㓦T0́*�Z��;��2<-����(��A< ��a���N���PG�fe��'�K�<��enjV�Qw�p.�o���\}ՊM=��̒�Fn:�d�9���B{z�z�r�7d�H^d��)m�������w-�_'��� �=�[�Q��l2�x��k��0���!��.bs�����H0�>�N�����S�\ȜM��_Un�!��̒WV�AH��4"��{����I��T��B��۷�P��n���P�,\I�(4fw���nM����e�7Ke�]�_g[q�>Ή͠ �]�G���A֤��$\�r#c�s��d������݊��J�N��@���A��Z��҈�`�J>bL��S�v,����ԽBҰ�� `��gS��>^R����͜C�b\���]c�n������͚�-����������)��씈�L��i�F�R�C�;�x8�*�2RK�T���d�Wj��[Xk:Vʺ����C]��v��l�p�n�|�+GjV2�f�S}f�/����`*���-_�z+c�Wq�Q�U�����w����3@-h �ۛ���T��2�k�m�t���C��Os���&��Y���[o���"¤Lt-Nhm
Tot�)n�;KJ�b����������D�o	{�V��Y�X=O�5�%M�Mg�fh+�����V��vW���E������[Yv乛ekbs[�F��Q���#ٕ�C���"�-&�q�6�)�wn��͒�Di���d���$ЈQ���n��ܰ�$dLj+������Z��	
	H	1F��T�X�r���\�a��Rb#W7f��F�Ls��Hb��"�u�Ě4j4��̓��DLJ8]�lRLRbH�0���D4F�m��q���
5˗v�7w"X��r��滻Ɲ�,:l���;�t�nn��`�@S(ƹq �]�4r��ZI�ݺ\޹��w��#螜i�7&,���F��S:�£󊜇��4r6B��̔u�
�ѻ+��V�s�.W�<2�_3ݗ�Q}�N:L�W�ooY׸n�O����8��=�Ը�.�Π&\�rT�X�J�p���4�9��]Q�Y~Boǐ�}�\U|f�ӝr�w���!�ڂ&��d$���֮�r{��{ӯ>�����\�XЁt�,z>,���דk~#�����s��+��]71
kR�+s;�z0��qj�Tnvy~.b��h�|l�-��:�{g���ͽo0�է�Z��[IL܎Ζtn�
v >��M�R���tS��ZLٴM�Vl�n���Ёc{��i�u�ʿ�`�гbML}ws���ֺG��=*.�Ը8���p_.��z/]Қ��ʼ0�`�V�k����;���;5˚�ٷ6~���kt�慉�:�]_1�|�>��0������W	GL�L�q۹cVe����岐��*�_��K����0�\cn�#8�;l�P�����yɻ���h�V��ݮ�b->���)g��^vy���	�q#�^[�T[6��F�$�� ԃ<����z����tF,/WR	BV��tc®7J�[Y)�4ۓ�':�*�ܫ�,<ވ�&I�T۝c2�V�^���>�භ��.���m��X��1�¬��
����8n���.au�^ڭ�xE��w���VG1�~����K����r����_�����D&� S��kQ�\B��C9��r�o���i%�y?���]MeO-������΄��w*ga���+*9=����_Al-��w�iX��[�D<GZf�^���"��q[�\.gj1���Dsûe��)�t�U�m�ǥ9V.޸	@��q���c��:���ۜ�[޴��<۞� w�j��V��W��ȉ���1s�Qg(�ѥ�F�3˓���k��?e�x}�Y [:�;�F{���+0u���Z���ԣzQ��n���Z�jeXK�#��n�?g��7�=-��lw5w�b)򨲹ޫW�<��+"Vl�R��s;�i��S\�u������ury�3��Ovp�F�MNS��&��@�Nvf�v�����P�.թ�lW�k2Օ9Vϯ!#;C7ʿ
�óO��[�	�mp{�ͧ�!���2*��fw5�( �Y#o��َ,�Yr=���1s�2��V��G]�N�#���d���V�S/Q�cJ�<�Ǉ{&�����_]#����k��7��F�ݿ���n��<���ݎ��t,0�d^�$L_^�a`����ޛ�V��)�Zc�_��%�)L�]a(��������.����Y�}���պ�
��#��	宇�Q�9�����a�F�r�������,j�`�+^X}�
�5�+iZ6�n��zc��]Z��^|�OW���߄�M����`����n�!!/+FvM��Ll��t��{q+a�	�ֳ!�ٚY�km�Ŏ[B��S�"���C�E\�Ѿ��>�S6��3�.m��?�a�(�����u���f��9=��V����r���u�l�����^<ݧ�w���ť�[�Ru׳Nn5��c��+�)�k��~��i�c�4������e���$�@���vHQ��[K�{~}K'P���5;�m}�����y 8�X�%u�(�3J����!��za�seY'��s�K�r�n�|�}�2�6����$����d���n�����F�nu�;˅�2�ي	��c��g�9u����2�!�^�>�">:�ħ��T�mDy �i���*�qv�B����o�y=Qt��q�Ľ�}C�F[��/e����W�{��;��+���ʣ7��tO��')��Y�7Z��=��e+W���S�ϩ��*���؄���H�NЬ~믴�Ҙ��^��(��Y��P�br1ΑoP����m���s���u{�8��׀��تC:�5ȑ�p�+�֨�v��+�hy��m9����R&&�5o�R�6֤:�O���j`�VV��a]2�GƨzN�$��=]�X~ܔ1�ŝ�\٣S|���r�CscW�]�;��[���|�j%��[��g?p�	�1{(���OXa�������!u��L�H��9Aj7]�FGZ贰8�<�N�D3�+��Sݚ��IN\P��?�`4�-r��r��$|�����1E^M?�\�pS������VGSw
ߕ:�=�}z)����|�c�{t�s�U׍Q*�R6��zw)L[{�fR�.l��{Mp�0�{%�tμ������0+޵��*�Gle�����U��(��%�ŏ2�.>���h��?��c�x���{��mg�:�9Y��mē���6��&A�M�S�l[롋M�-$�vf���M�9q�D}��:���S�t/.�9���VOHS��B�������<��R
S#oN�.ƹ[�=�('�)�K��_}`�����Wl�����9��!���!:��1>�T ���a{�����o/}�����ؠ��u�8���%��7R��ʌ�|�������Mm����!���j�Ĕ[�P7A}p�^�ʪlb�\�6m�{�(�E��4���^Al�����8qv�=Y�϶���S
������].�eDqqʛ��5���T[{/�ݍk��;�#�'���@�n�OW=
�5��\����j9�ۇ�;�!lJ
��u�ļ����Ü�z�s�/���-	֦��c{*{���t��gu�!	b�������Sr�m�7�މ�|��)=T�J쿖��2��:��q�Q�Ϯ�l��ݣ;���օU�j�I��\WsSq��"�<��s׆*�������mX�^��B^g�Iuz�+U:'J��S���E��d}�t8ې��&�룝�u�.UI���OA�`ʷ���a�jW]˱��~+d���%�u����C�N7�߳�uAx�ҏb�72�+9p�ذ:oI���@�4i�t4UZ��<��-�k��0%_�[rw�&�x���7y�k�M:�x���5%�����sw�<�Ҙ��eTa���"����w+�e}ݸ/��Lڼ�˷�J{uT��Z;��Un���T�5^��yb(9��$�B�4��o]��+��Yu	u\٨*㓨��<�M�.�Ց竾32����3C�5���١\�HS��T$����c���F��[He[]��v�L��a�i%�G�eR�c{)M�����}�;~�jzZ�B����N�F�c������g^�f+Ǜ�A6u�ydSYۘI�V�	��Dd�:3�Nz��/�o]T[C�Ȣ�`�qf>�!o�M{��{�#�B�tns�^bO0��ώ��qxШ��.yۙ�B�h�0R�8�N��U}�1ָ��ʛ�����q����`�7��5[߳7�Q��[��͎��J1&����=lako�_Ģ�ۄ`�Z1lc:���V��v���p��_&V.|DK�Fd����P��6��{��b��%%b&�X�4�,&:�㎉�4��$�ږ�噛��N�D=�N+ٴ�����7�|�*dn�7az%d��8�r���u�.NU>�gǳo���i�d�x���o痓�I_�hw+�6��v������v�1��c�
cz9��a�3�6#]�=�t{�����/���AT٥���]�'��+���o��d7�����;*��8Y_D�JQ(��ҕ�]�3Jn��ԱTq]��=�z1�o`u��`I�:�d,�P��{ɿ���@�)���}���s�Ϻ�90���w*�0�ӥ3���[��]՜6aS��R�#�х��M�K����>��U��z:��M��U�N��j�����0�#�p�@��n"lJ�p��z�ⶕE�C7:���l%:�Sy�����yl+��fP�	x�A�]�X��ge���"뒣:�e���q21��L(y��隉jي��>�e^e�>`�Y���:o=t�<Y���<k.�sE3L�`�B���"�fs[I6.�hU-��,�n��u�<j�����7;�wݗ��x���x��=��t͂�dP��ޝ��
����gR�B���K�G��E>��d�9�VL��'��p!'ڙ�h�L$�7�}����%w���4� �&��k�q���J��LmBs���U�]�DbBQ��1{����3�r���V��Ӫ3��J�d&:m��˻yfj��7��%q�صq��7�Qz�'N)�ت1F:�Td�������ڧ�}ǲ�d~���^A���6~�YP�Y�*�qW�q�أDix4L�7�W�U�U��\W-�}{�>=Qk
Lݎ�y7Ԫ�)����e��aC�yIH�C]f���Q��z�䵏⯲�1�QbPU��MEu�����ncz�y���M�����/�ƫUW���>�����V���ߓ�A8B�Hm]����Y���tvNڢ;��<��ΐ�z->����v.ڰ�Gݱ�M�I[�~b���-�5%(����.��\�J!��PT�yf`�eNNNJeb�������}� �hvΗ�*�wk/�Ui�C��t�;0���E�}=�r��>>�&�hFu��	V�R�A���-jj��xOxm���s���\R��gv}+��*����/:������7�Z�z�6٨��	�I �菾��ň�V�b�z�r���*��0��P紾����ң�2~BE�Q�Hp�Pb�����J]��=+~5Xc���+_B��q��߯Nrgir��]�<��koD{ǁ��y�yf��o}ƽ4��9{B��W�mt��]�p�G ��K��p�C���˘�CZ�$
�"�_׼�-��KDŕ��9�R�8��DjɈ�
c��I��S6����F�]��y�抄����>F�^+���aw����Y���gl�B;�����3V�9q�]l;��Ԛ�O�ٝ��^;�y�/8���qY�����+w�1&���xmc�4��l8��/^\e꯯'1E�bd3fX��PƇK�=��S���]��R��ι��~fϻݑʠ����\�2��i�[��k��*V�d_=++�Pby[r�k��Q�u}k
ۇ9���}6�n^�7];!��j�����N�+���Pp�a$HӺ�E֎z���9M�����C�}]wf��睸�j����(�kY�/�˖u�[��Y|�/*��v�+#����K�I���}�v	��,�V�Qp�4�m�p�����Ǹ��gf��gw��W��u��z�2~N��㨷�Jʍu�ǛQ���ies��YW�v iY��{��F���R�rϬ�/���Jw&�v}��f �
C�1��j�Fr�����bU)�Zj.w�i򨲓��j�J�]��n�fm�Yw�m`P$^�j6�7�4,��;�T���WsSظ@���9ǵ>�iH����5p�v��{�w���}�jW3X6����x⛘yJr):&��_ڔ�]�����=0���]:Y���J�>�^��Շ�Φd�=�w9f\�;uT��7���U��
ʘ^B/�Eˌ�<e�5�#U���������o2f��;WZ�l�ҤL	]�}�t�T�')/	�����Co7,��i�^�5�g=���zB��jR���>�r�pU{���Qz��:��3ݾf�07�'�0�X=�USqbǘ7�����Ax�L|�]|�����^N;B��b)��3��\;���YF y�X�ޑ[��3k(_�a�7t��ƥ�q˛�Z�eK���Q�\\L�۹V"�%���*�]����ON�G�7n���S��ʻ	]�K`�MQ�>�f��u[�^*G�'+���4�����Wk�>37�*��$�j�a��,�l G��i$co�ZF�Vօyd�i�7hZ�j�OOc�r$���C�e�:�5X�Y��	l��ܷ�踃O�:�E�]�%p�G�E)�K]�Ϋ޺Jʾ�:��w��k�2nK0�y&ё�cT��=4�۫����AG�2�|�*�s֙a`�D��n����m2&���dr�f��Œ-���l�8^@��������"�j]��$�5�9ago{;f���ʐZ�v�Fs�.�V�<�r��*� jΘ�e�bƅEJlq��d62�-ԣ���Xμk/:�/�R���rrܾ�9;�OMkFA�����"���dW3o�>�)�y��iSZrAy˭��Ĭ��.Da+��Ӵ�\�b�x9�WC��A��V\{W%[��_+רD��"%�9��6�_����sA���-�C�N*qŔ5u���=륆]�]&ǺoV<TJ��{�+�ym��������p"�׸�<NP,d���2� �h���b1Ԗ��n!��M���J�-��@fۀej��ɫY&���`�:�h����,�,=�5����K��{j,����&&;o�o2�.�.��n��v������*sǲ\��'/v���)6Q�B9|Q��ޮٌDB$���y������]Uؑ�&�|�vaڏ7qN�c����h5`v�cw�I�B����Z�R�Q���Z涺��J�(A�:&0Q���Yz0͙}�m1z.��7�T�.�#��������R����؍�I+���&�3����.�wك�S��0I�daTrU��w�&�!te�Z���������k;7(�7gI�tsJ�^�vWpt���wa��u^���b�+6�+�=�iwI	���c����
��q�X���-��w]��x��f9n� l�r�<"���dA�YE���,	� �Gr���yj�q��#`5��t��T��)�]�{m5۝v��_V;�}�$�(J�mR����]��-����-�L�48_ 9�͹��>��
�U�w�jH i�/hO=��G�;l9%�����y���J���=��%�W<G8��M^=���d�Qd{�/'Z��N�� j�A�I��MP�8��nN:����b˩�G�(�^�|�+c��3�5�췽����4�����;���8bw.X��EY��V�Rʉf��D�λt�a��}����7��0F�<8S� �fl��b�Z�v�t*�}/um��\b;�4��.��]�)>D�2�nWfWA>���b:SU���Fj<s�`W[���z�ݱO-(o)�_il�x�IG�뿯�>=���߫��r�\��9Q����;�.s��'9�wq˲�w;Gcl��w:����]��sb���˘�D���s����(��6��n�AF�GJ9\3��r��Kt-���F���tp�v��r�q.b�]�	����]2n�"R�˻���˖��ة��I�半���Ec;�]��N��s\�7wwu���\�t�;�5�#���wr�st�C��wݮ���s2�.]wwv�ʋs]�s���]v��n�[�9Evw'k���pb�Wv��WwZ��Ի�����]݋����{��רq�z+b|�٦'R%�2n=����H������^x0�~�$�̚Sˊ�хt�+ x���h��
9\�N���}�KW-J��_�-�ڴ�b����ؙ��Fs���o�W��ϖz<c������ڎQb�VA���**#_'8k��p6���/^ ����0�wj��w#HPԳ�'�T��L��s��zx=�?6=���A�-�B=��{fw��͸ػ��;�U�U�k�������Z����q���@��AL�ZP�\b^��9��%�T-ڍJ4��pbyrs(pu���������I�t��&���M>C����6�k�m�H��ҕH=�WD�o6Y�Ep��{ɭ�naMo_��}c����ߧz'�|�E�Yd%�����6�n)ƛͻ��[ǡ�soQ�S�x-����[qQ��t��u��o���w2�<����&���섃�{��:��R���˻�S���3�𰖰��T�c�M��tOԟ9�Ә�=���X���)���̞6�3���eU�^�!�Gکٮ�|Y��E�\��wש*���4�m�;��}S����PS7�� �����(���tS7��+t��K���J ��emMe����1�վ��ɨβ��`ړbf���m�Nu����]R�4�kц7�G,ؓs�O��컌Nk4*Z�|��s�*$HM\�lT�έ̮Cfcj�����B���.�ˏ���z�uB0�9Ã*��rY5Tٶ��Y_'fU˘��B�r�!X2�&��f���o�94W>�T
./(�Dw:5�p�9yN��d�C�o3�"��{���*Ӿ���p��^vt��Lt�?v�t����q�Ls�zk��k��=I�Al�v�n�ZH=W�z��[Z�O:���ʍ�Lk	�/&���_b�zfv�&(�/�S�����J\P+��c~}P{�v/Q��Ҳ;~�؆��z����3:��Q�m���+�=�~]K���Y:���KO� ��Wo���^���z!�R��� ��8�]�B����s��j^W��p�7�gA8q�ķ��E<چ�]��XRf�v|�j��]z�SRE)W��ތ>�aۊV5{΀��U�7i�ዄ�W�N1匫xi�KF��c��_(��IJmc�Y������j�)����KE�e�ms�IC(��II���e�?���!ݳ��_���J���e�{�B�mX8 ��S"ʜ�Rӊ�7aQ4�ޝN�ޗ���<M췝+�G=�`���GaLc�ύk�w��F�Q7��ʲ�Y|�k�0�v��v;|�򎢳��h��S�o7`6��l��ۚ���O�}e.�K���,�{��>k�p���ײ����ܸ�{�����7c�eI����rjoLV���V�qYz��y׫d�7S|2~�IXv�\a��`������밹���x��:vsj�'����L�/����qT<�0�T����~�k��ı��f�u�4uF(��5��UA[I
c����ª�/*tv�_�5���W�L�CeBZS��q]�9�3C���-�p����尭�X�� ����e�sN.��ۗc��*�~O��U��?���wz\)�vzq_F��1��Q��^�do�5�y�i^�X]�Sw���{����mU�{|S��Y���S���iМ��/{g�(�|lZ��62��j�Ů�����8���K)��j���1��ɸ4lސ��\fU�Ն�9;[Iq�Zˁp��l����b���\�2�<a�ܣq��V���W���qz�g>[�u�AGX{$Z� ���5N;����Î�_���ʿ+Õ��ΌQ����X��[;�(r����>���ڽ�m}�+;��[[C����E��V$����	�;�JΦv���=Y'/Q}�?46��[<�g�����YX	�)���wY�6����TN���!7ܺ��{�'C֗�nj�t�Q���[o<�J��V9��M�V1���iYQ��+���i�.sR���[Lc^k��3����n��spkZ��ʾ���F��4�w�&�N;a����\�M�q��w��-שּ��P���ߩ�);�i��7%Q4�sO���oZ��o�ޣ-��+o�ZW���&�Qu���T*(M_�h�cz5�IqKR�-+�q�3��9�3�U��0/!u�&�TO�LN��sx7�άp3;�LV�	�7z9��d��5	˔j��q����!B���[���v�B�[��f,�"K�-f�jbDa
��O%�G!�-߽��j��6���6t�Z�����zeYsdM]5�;�ʘyВY�k�2�o(i�7 z^UqԂ޵9�r��+D�Ò�8��`��=.����Rt{�ũ(���*�&I|.��!{�	�o�#WޏPŭ�f�+j�v��un��׵�3W|�8-0���Wʉ�+r�'�
���m+�m��M<{0y��[��е���\K�s!�۷�v�a�ŏaVt�v��V��]�:���k�Vq޾����p۲Ms�&Wdfb���}����TMf#��!KM��=A�����<~w�T��	��~��D��T0��HKCov]��?���Pb6S�풢����s�S�α��[d�s�s�BS��72���ඨ+�����bzj5A�Q1��Ůgj1�Oj�%_������xZB�
�ژ�!G����^�~��o�*v�N3��厽�[�S�R�Ϻ�k^�Q�o{��E@��Y�>8�}q�(�Q��C�^ܗ��FR�9��M�U츊��k����efshUk�\���C����I[Q��l�GXa�%����T�j��p4uTt³; �Y����8���V\B�)�itÜ��ܠV�2��˱n$�	Ht��U����i�W�^~�֬�/KPN� y�!�,�1�O[�e:͹�q�;�]J�H��\�#�{�Տ����2�ur�R��x����6���7�
{��</�1�UZF�j%���:gc[��yku��z�7���/�����Cݸm�}
k���+o�ê	Gf��[w�*��m�uv��鷺N�5}����+��h{�Qڇ-��)4(�<ɢvM�����˓�Dus8j.+�9��]5�D'ܘ�]�0ʚ�v��5�y�����S�.��U�շnb
}wv]���n������<�m��<7}�mH����~�*ʘȆ��9m̓��ya�d*�4*�uM<�˫[��-	ɩ�%�L�q�	ٕr�+���^^�]]���N��SS�{j.�s*�)�t�?o*H8y�d:�:��t�+�>�3K"�؝ѪQ��i�w�k��c�ד�ATFl㴜�E:F�c��ӷY���92�7(�i{pNE
�犙s뙵y�Z��Nc��i*7�����ݞ�uu.���&c{��6*V]����M�,{hG�4�wȌc��jC,n=��dI�#^:�F�	����p��kh{�zPͤ����ǘC�b�0[K�i�js�캋�혬\�e��(oe�F��N5�����fA�)�̫�c���y�-�Xo_�����B�~F�]��~]�R�g�:b�:U���ήU~>�3_������e�Y9���أj��V��
���Mq��:�qm��ygq���v�ȼ�vqdYǔ�t��gJCVB�g��������]e�e�<޼��*�w[ph���g�P���M��L��^՗���+u7|�>܊oB�����\-�Xz�:�H{)LN+��`FWYsQ/z�*[�����y�]�����xۋ��Tf�)�x�D��.��((�q;R��)�)v�Xꅡ�r�L�59*�@���cr{�s����W�vZ��*��-!C�J���J��O/�ډ��Y3�`�V���_8ܽr�|�]�9H��\��Ϯ��j�/L���̬P�k�E��+W[y�[ъ�Y�h��a��6kmi����K9��t �˖-��}�+���AvZ@��y̅]l�V�S��zg8�E+5��yd��a�xlb��4���o�Ө���싘�Um=�/�t�M���}7�]+�`�T���>����f�r��FI��m�:��]����b�3��♏�����7s,%=��ⶕ�#lu���C����,�*Q�&�'�$֋�a8,�:'7'#9n��\�b9m$<
�T7pw^�^�D�:���C��f4��s5�f?S�8��F�뒳���7�\�pҝ[��]u�g"c��*n��?$�h���]웽�e����^��N��6	�6�S�
���.��>{qw̢��bߗ~��7qM��@��_W��qS���΄�u��Q�p6�ai��v�}6]\���%gIz�����Si�	�Y'��������-��?�f(\Y\�,����o/�L
�s����b���A�Vܺy����Z��	8;=;zu�
M��"�3}�/o��F������_S�\�T���n�H&�s:���	�3�����s�4lR��C�E����Q�;�q�%��.^�VQ=�,n�[6E"��hdX��վ繊�>��#�+�����/Q��4&�tH��z��1��_u��y<")�3�n\��)m#�o�6,�	4���3'J�B_,;]Zɖ��@�Ơ{b��Ɗr������b
%���񝰙r�����U�?
�W�3��ʅ�q;�q�XI�Ov�
��
�3v��Ih^O<�����4���+n�U�ZD�J�C�a};
9>�j*U�ˈ�S�,|�J!��ۇ�&��u�Q�.ж�bfo'z��-T���.������@������
�4�ޅ��:�<ʗ���F�s#I]:2��~�udV�U�������w�o���nٽm�#���N-��@��'N'�Bb1-�U���o�ene�O2½a�%�c�j5�%Q �ZV��ը=ل+�p�K�����O62Ø��1�ª�p�}%�۽���[���#���
n*������6f�\Ff*���P�v�kMe���ە=[f�$^[���9��S��;��*r��u�ߊWd��l��jbz7\q��[���Pb6[������w����g�dQz��{�qF1�n�H�UX���QE����)L�ߦ4��z�J��m�q� �_PҘ�,�r`3��ۏr<PqS��p���ׯ�'f�����<E��鋩&f�c��3�ź3�,x Ńz%�z��J��owY�OC�2�E�m.��I��r����T��D��QX�����P���j??S��U�͇KQ�g�]^�MM�mҹ���D[����qM��j�>^�)��|E=۞)8�O�)��݁��{{oK�������%p�,8�h���:SC>�a[��qp%f��U=1��Vˆ�����l���V;f�ֵVq9��>�ت*��Bh㋬�xyW�[���_;{_){jWx{_�~��g����W��P����A��=�Ŷ;�j�ZSǡ�6�+�y�бc.���`��=����
��`����w#Q�4�໻���щ�q�J�=�8�T�w"M��'A}|V8��UB*��n~)Er�=�����e�Rv��b�z�)��wo�����vf�c�K%6cR�6��V���R1�3�i�!;3B�!�8NN
�a�یO(���LSP�`冁X�@}��"���oD嘪��*t�U�W�e�k|�!�!�X���O���"ｚ�q/rʰ��A�G5R��-�o����Mw"|O��O�(m:�V��E��]��6B1�!�B�7	]9X�d��3�Q�����.�\��#]��,J��6��(�63fV%[����5N堳1嫙�WyG��H�(���28ǘ��)˼�y�{}ē���aߤ�I�xMKN��F2��޷�</�֫�q��3v�����4cXO���#lpSb�'��9ʀ|��v�����˦F�d"������������-�
�n�ڇ1����sx����cr�ů������m�.�j�IN�&V��St��ns���t����+�9F�}5V9!SgX�֛�K��º�^3m8&�]f��g`��7(Ȫ�v���T����\�#ۻ���OC#y����ޜ�CR�����~m�x���[�l�b�O�W��E�PDՂV\�D�PQ'V+yG���(T-:��B��ݦ�{{��!0���U"Q�7=�	�Z;��3z���V�w��O���G\��/b��4a��7�d���yṊ���NChn�{S��D���.Yl�!i���Wk�ZcC��B�t�2Sc���<��:K��ڽ��S�n���B(��QΜ��W ������Wy]';����Cr�^���!I}6�rH�[��xꮪ�D{t����R���s���+T�G jw8���g��������ygz9�U1l%����y}c��	̕�[���; (.՜_��Q-Z��E!w���X;Et����<r�/m]�kq8��:[�n��cln;���լ��n��8"����y"�K��7H�dEym�ڝusH��B�"��o�Eo.��\\�eC���ۙ����WOD�밢u�j�����}h;��=�m'c�C�,��U��v9�:��4F�G��|��ܮV�o�9c/�R�W��ξ"��ի�c�'♱�Q�ӝ�M�}���Z70.Jq�%���m����)c�cj4p�UЎ�N�$��9s��������ױ��,C��[||K��_]�1��Feɽ9ݫ1���VQ�Yt�ȭ&k��ӽ��.f�rP�f�$��Vw��s�Y9�4����]�^v\�c
TZK��Q+���.�B���o 2�f�v}�T<��z��@����9oj@$$7��#:�rS3�B���#!�e4

�B�Ԑ,�ޮ�}R����L������X�2��[���R�q��%gIpЏ���5�Rhq'/�)4؀ٓjp]L>.Wy��ݝ�wHb�ny���K=VeF5���E�o�����dq�̢�i�s4��h�Z�ԝH�Jħ�m��nV�g�P$kMaE�0��ԮQEb�Ki��NR�ON��x��5����;�bR�s��T/i�w�v�Ѕ%��(�x7�*u��0,����]�Ǿ�����'��9�v���t��4�����1�N�t�s�s\�N]��wWt\���I`�뜮S��tA�\����$�sI��"���q��Ε��N�J�����.n�5˒B��wC�nEΐS�S��gwl�����k����5�\���.nDQ]˺���'us�1�#g:+�.����B��ݗu��#s\��Gr�w\"
\�(�\���.s$��9�7uu1&��g;;�8��6��;pȡrv�����wu�r&ԛ��ܸ��
��9w:\w0��fB�s�]û��%���9K��'u���k���՚���=qMC��U�r!�o���#�-���}}�W��Tz:.�'J2r[�+�/^�n�=�͵K�4q9�u�K���gŷrM���xh�GRvba[10Z������Rܵ�{�t�v[�ڹz�v�s��:H8x�pG9s�h�=u�N��e�L���vfU��\y�T�����e�Tx]%��&�D#�Z�b*�ma�Cx<߽E�y�Sda�~E{h�=|�.����**11�il�4+E[*�����1u��<Q�]|\vT�.2�U��'�inI�v��݈���+ή`P5p�qq�����=V���E�vt�T}�~]X�%����nEU��޾��5$R�J��S��i���/ ���l�,��W1s��`�S�R�uw1��
x%m�̌Z�1<��ȧ�P�v��k
Lrw�w����C�+�k���<���1�|�,�-[|�܊nJ��OOw;4)�[�U��j菝jO|d������TGO��B{��zE^>�����P,�{��1I��K;�`�VclS��.��鯕!�.��n��ީ����0׬�D �$�Z���@{F�6��=���l�t��7�K�W���-o8K֥�L߲��#�]����a�_[l��O8���?����;(�qu�\[��S�;�䳃u0V�]L��Q1O�����v�L��!�s�*�N�ZJ��Ep��K�p:�V0r�BۓS�J'����.Zꅕ����-<���Fn\E�N�|;S�{S��;r�]-�71�]�w��F(�tM]ο�zr��Z����^��~��_��
�g�B*a����2L>ܾ�Wp���Em+F�����O,�#�� ��?���\�υ��>"���2�&���
絗_%�S����X�zs���䆧Y��jj�	�����n�~�Y�O�S�1��j��
b3���dӌ��kf�W�
5�ͻg"yە7i�9�����+�+��:��u�4�]n�����T�ڷ��z�p6�N�yw��\z}lﶯ1��������1N�PX�f���Tv�(����9�_7��\�.;*ׂ��0L��3�;{�5�)�pL':k�\br��{����j��L�-��~��ڐa�[��G�f��%E�U�(��*"F���[/z�*B�V��lI�}�v"����p�,�`�zB��M�,��nDv��+W+�k�,�͌�+��c=	or*7�A�Y�0��r�HR�.}JgVI���NUw�
^����-$\�W���g�g��f{ώb�[U�1hw���O+nrޯ����':�j�T;w�9��W<����hy�M��Kɾ�cŸ�ZVV����ok	rb��a���j�s��7r�K#`�R�pkZ��ʢ��zR\�8����bN��x��^�H��=�͈�C�^�����o88|%�V]f�{�����ԍJ5��]?�mW����ۏv�z��#���w
�N�7��I2��9sx{�cL��T�c�x����۶�d�tݎ�*�`Kk���V�GL�]wF@��c�At�z����TS�A��;�7�ݱsu�lQ[ԟ8���5Xc��I���ٖ��uT��3z9�\El��}�;B�Q�5ؗr���პ��`�J�ˀ�e�W:�5̺ほw��h�RŊm����kE ��vf�-�`)��Q�]���CǪ�uXФ^�1��o&�{�]�N=c��|�\���� �����Ϥ�Ėh�2n>�gY�d�D�TRpH;�u�A�������S�?*�1�.�.���]�b1c�HPw�<������=R1��M8|�C�(*�x7Z��))�ru»W3z:��W7Y�g/g��*���g7�:B���.���m}�q�q���_f�]��
ǋZW�Q=�+��v2�u��0u/�؃�Y�{Yo���*u�{]�Y�^��~�(�(��1�>�S:��/Q��l���:^=��C?_�W���E�[ߐl��EpcUSh����{_�7���&NVa��{��w��.��6�<��NA���+�9����w{�>���k2k*�V�櫧ٱ)�s��i�[q�ߏ!�G%p���_�mg:D�a�Y�,���.&�����Q���O�]�N5:寃ꈶ'�ZE��%L�+�]�1�q۱?V'V_;�j����=����U��O���[��|�h�AYF�ը�D [_Dsp��Ϯ�<ڐ߭�����j�"����!mI+�묈z{|�'G/��~���-���Sj�X4̹�x���S=��z�����j��:���,�@G�X�},[���!�w�GiՓ�]���c�Q���}n&�ĵ��vwխ��]�
c�s��*�,d��3��yܕMF�K�3��!)����M�J&"�s�]9�AO������m���gr\	�댘�t�2�vJ�rۓa>�����x��e���^gXj��3,���g8'	C�:4�-���BYQ:�xQ������Yz�4v�q�&�i�2�;�T����w�;3
��T��<��16EFN�1��z\��v���
�:B�r�p�>s�f�������Y�N�tgص���X3�uy[���5�8�q�%�$�����(Ur�ܸ�wB�&�Q��^�_�hOFha�i�y7��.����<S-N�J�.d��
-� L�|�k�6�Cp�|=��h?)v�V-�w�ڧ���.���&�+Z��ǧԽ�Q������u}���h��ζl�Gt��=��D9:r����>�rWN:)�zl������:Է`��X��党36f�����'Z�8j�rM# ��[�S t�7P;s���ou�]��:F�Rm�g���.Qr!�1q����W' \Td���g��^�ώ,����ɖ����wFr�}K�Mv~��g�z�q�mT�>4��ߗ�{��<�|P��@}(V�"�yl�+��0��c���c�/+T���Sͦ��^��aK���|���z�ou��d�M��;��[�Vq՗��JڍM�>/q��s���G���[v��6e8ΉU�V����:�E�UW;������=�ܭ�}(183�u֑٩�U;��XvV�bUAJ�MA�J&)�w���0���1\c�ŋfڼ%��r��VА�Z��Ң��$�s�[��!LMobs���7N��%�f�\&�ѹ�FM:JneP��@��o�70>�wU�CA�;�!�H���u^8�w�c��Uk돛�
���O,���O1dUUX���K&c�7���ˀ��ws�+���:��U,��1���+Y�y0�ϥL���5P�rۛV��b{��W<Ø崯�\=�=�.�j`#}��L	83�)ʲ4�:���>7��=o�7�3��&��Bw� Ug-r��&B�Zd�mfŹC�Z�����׎�c���{x��5�n:=]y�h��]�����q'c(v�j�yj�E�@O�՗֖s�/]�ێ�,�;4P��ΗWׁ"�RYݽ]�L��R����f�?%}��/c��>So�����@�V.�;�S��:����;r�K�ؙ�����XGM�4ge=.k6����sF�S]'�8ٶ����.����;�ܼk!q��Ύ�f�#h/����lv��q�]F�w�9Z�s�4�T��eAp���sf����t˩�r�q���1֨1*'��O7Y�f��k���y#��4I�����^2�����X�iy[�&)[sm6�X���j.�o*箎v�\2����j��[��+���3{h��Ꝭr�����c�d�����׶��ͯ�ŷ�w^!)C�&��V�Qg�}e�q��u={�3�Z"ru���]-�J�޼f��Y_N���*Ud@�����Pv�8n�L�6��r��Z�һ.����e�:���*�B�w�g�ǁ,��uk����Wu�C|aX�;X�!�.����vsr�i��!h+Nٽ6r��^Z�Z+���Q��^�,,����]��e:zI5�\˾��R��X�>�}��;�.�%锝��R�{a�Oj�X��u�}�n=�rB���ኺN�o;Y�кǨ����'����.����K�n��_m9n��t���m̛���Q��	�PDv�J;�$�jl-oun���sw�/�����"P��y2Ni��KWuja�Yu�J�jۓak��.̸	�v�+[\73s��<ζ@���O������7�u�[X�g4�U��7ǪӤ�!��I*v�S�qR2�O?����Y�FG�/�c��m���y�=�#I�a���݉n5��M8s�}�JN�R��J_{ބ���t��W]iޫ�����K4�Ðywax��9��
c�K��f�w�k�zu�������lD��x��C4�3Ѣc��������>�n�n�E�	����];Sz��k���L:�`;�)��]�檋�ʌOMj�Ңcy�x���S��z�8��p&��ϧ�l�Q[]���Lt�����'+�h��n��!y�����Oki	#�j,�|M�����@��z�my��Wzn�=��|պx=���u�c�g_H��r:�<�U�Ǒ�&Uצ�9�W�����\����wuvhY^�����^^R��A�n?��]�D/3���ovƵ�Q�K��6hm��yrs��i�[q��Gְ��:棆־��0Nl�
������tF��4�v�}���r�[��__�Ħ�1�V�-�ZӋ����/bb��Y\�yaҝ��_?y�L��� �w��{)���~�:Go*J�՛C;�>�d�1����w��⛺s��!�^e�fvP٩�����*��nM�J+�9���Y�kX����&f�m��f�U[kV(��S̩r�
�ڤ*s?`8;��C��Z+�.�"���EjwގLZwF�b~j�����F1=�ͯt��G�s��
�_<�U���Y�m��9��aT��Д�$C�p����p���;w�q���ʳ|�q�{!�W�m
�Em8@Ē�����ޭd�*�i�Х�ݎ���إΠy�kV_qYݱ!!��Gi}�YBt�7y���Yq���T�b�bA������u5�/i�t�=�&3w�%ZT���%ept�p
���o��̑�郀��ڹ�w�Wي�ǻ�t�G$�p�N�+ <�w[c�|�.uw�fW��j23b4���g?)�Vi��p6(��K+B�\/0y�Y�+��3q1�W�����	�ÿnmC��i踍�B��wN|�ԡ=HT���;x��H�=����V�d�l�}�ၙ���/i�Ŕ��U#p���;��K�R�6g��kb�h��
�څ�@ϻӬ�>����EO�$�e�/h��8V���&�O�$��Q���[>n8�6�N�LR�g�D'^�9�\�՝q�
���hp{�!V=��+�BO�w�f���u�� k���ޖ ��No�4�:;�xc�^�bO3n-l^驷��������'�P��crgY�|Q�!��~�i�9�w����!�F�����;^���V����XW���9��8�1@ew����L��s�P�Saх��ˋ��xY�~����Ou����C�zK<��"��,�#���s���QC�*/r��uD��^�*��G�O�q��z���̲��7΀}�U"�%�~�C��Q���GiQ;?8M�3�cf�":����ܫM 7�����]%����Я�����ܟ
�=��_�b��;@��A���l�����;>I�]̑��]�Ash��j��Tק���j�`��\^���,�ީ,��P j��q[�Wpr;ۼ���,4-Q��`᷸����.V���Ds����Zgpn�/ާE�%��	�{�)��޽R��� ����U%����(Z����d��C/
(�5���j݃���ٗ����i5�Ha����y澵T��Y�{|�{P����j�3%.��*!��s��JkL���ـ�˦w��Na��/�g�uL��E���r���fn�Wmuk����� κ�V���������0�o�c�j��n]���VK���M$̵���%��-73:Ꙋ.����L�^��'�����|��m�z9Nȇ\�G)p�7�Nb�Z�̈�����{��ǽ�Sﳩ��5�4�ѷݝK���2�o�KkE��W6l�����L`Tg(���ڭ҉F6NVgY:�-Xo��&e�S+Q�z��}�K{��K��L�RW���Ys�]&5���{�:���}�-5a�j��5i�NfjN��+.��(*l�o������hL�$=�S9��<df��f�n�k}�
�"֪eL�ٌ�[I�i>���䅷��/�L�u��)�L�%���T�A�;�݆�܂.:�Cp-e�i���LxfF;qhI�����J�k{\�,�\��߱lvir�un��
�{r���i����N=lN9Ƽ�y��y��U��S�e�a��+�)�j��ܩK-(�HM�c�P��6��W�Ǖ3pl��(%jܜ��9?_dT+}d�Q�ܜ��7�><�p"�X�{��Uը^ ��v�f�̤��u��On�h1-�x�>T5].Z97F�,b��0 ������:��w^S}V��W��n�!e�[��r����1�2�[�_u@��ة��k���R�����މlЛ�-4�F"�'&�r%p*]�9C3ҧoݢ�)v��ኦ�:��f�f���u�c@�Ʊ���e5]x4
j[F�;�WhZ��E�I�2N�K�V�D7��Ҡ��.������Mbg-Q�U(]������nY�P[���9X0е�@I�[#T����}y#K#9.5ٴ�u>Èc:�oj�]��V���i�r!����(�>8�t@��U����)���[�vgU�soZ��tHp3��=��a��v��.�G�ҾR]q�Z�H�:Ж5+w�ཻ��Y[+6�ÅR�����͔����^d�I�q���O����3�6p���=pf���e��i:Jұ�(�#��m�\�逐��M]��e�5!x�S/�9mqf3J� �_�����j��ֆ�;�aYG�Υ�Y%�7�q^:;R�eaz�O��`q`=-�$ؽ\D�1k��{�Wp��N�܊��W@}�� A чuw.Ļ��ˎ�rG72
`����.F.r�wwwd�6��!C1$�;�wn]݀�%��79��;��;�
� i�SwpEwN�d+���b��1����#���D��r�,Fe�vs�r�"a$�1�hɊ$�]�3��s����D�˻��!�\�wCt��wpR��Gw2��:��pf��M\� ����1\�)wWWw'wK�v���wv20s�wn��;9�bwvn���̒Wu�LPM�p��Ĩ$�u��QL����].C�\�p�Y��N�����$ܮ 2wvcC*HΗ\7svFi��S,�w]��Nq"���"�]��w+������w$�wrU�ꛙ�Z��R.�x�xP�顣��V����fe��=��Xȭ�S9V�Q�����Q~�5���5��E�|=��ً��ϸ�=~�p��>���6 �l��q5让��>�=����=3�wAR��>	_Wr�P����s��#]��̉)��7�7!`�����r�����`h���Ȋ� ��h�-�ǫ������j�����S��y�R�n������I��#p*z�s�H��c"�Vѿ��	U�y�ן�~�M>)�a�@�2�e� *�w����������-U�SV�ݢ_�d֗��o��+����o�w�*�\-!�{�oY��΀�$���6�y�t=SEΠM�9�J���
`��TqRF�v\Oy�Q1~#Ϭ��UP�L˘�蓥����U��?He������a�������J�Fk٦j�k���zkN��g�����կ ds���w��b��B���^F��c��7E5��)-�g��6�;=Y���f�� g�:�j�{'�c�#�;�z$`I7I�����qn=���M�p�B�5�%�gET{FV�<���r��<3c�4�c�NN�����Z~Xl�n#�:��=�O'^�+}���c��{��˖�]�^Jx�U"4���p�}J�c �d���#`L����l���]�>8�ec�4R]x��n|^Z�6L#6���6sL�����1^
���NS;Y�jUu��F���C��6�w�g=�~��hp�a�F{M1��T�1�I^��~S�?�w��R��6�J�)�b�6sj��T�b�����_�.�Y^�Lw��Ef�"��u�������\;�&S��ɒb��I/^ﮞ��^�oy��H�}��*���j�*�7�E3n� �*��f��lN���g҈��:�%x�G:��8�4to�R����N�Юe�]�)��'��}kb��R�Ib��d��L� TZ�ˬ�a_�G�B����
ӫ�u5�����U�=q\#��ۋ7j}�n	Ģ7��z슩
��Ϡ���ن�^�ſJF���|�<��*.[P���*z�Y+�!�e����Ǭ�l���R��� ���	��P��V��}�>�ޡ��ێ���v}��W��{נ��*��#ńtJ���"��9���7�eOo��z~ӑ�goa*ro��o�Wrm�� 7�3�wS �yd��3>�W��rG���U��W����R�������Q�P�"c�ʽ717�S�� z�(
~�d����f�.Z&0��a������,�tE���C�����q���#6�+�?t�Ky�W���\��}��h\/p���*闝�T��<��#�K�vC��w��H��ʉ}���f����L�K�]�t�=,^V��2N�;}�t��c�ֹ�f���D)�X[�>���@��3,�����|��&&�c�=�}�����ۡ�F��ܤ�;�T�����f��`	��W����Y��On�"?_�5�΄�z��{�lz�<Q�?m�g?C_�T����X?1��a���&:c,v�ՙ�v������}VG�y���2�w��ߝ�+ftf�u�!�k5�~������&~5u]��i�>�|`e��α�N�x�G=��߹M��w���R��^�Qi���3�Zk���vj�M?nz��o�Z�w~�M9���N�{^Gly�s�:Kf��Sq�ڄ{w3�vW��p΅����:.2g|o&Z/#�Cwƽ��ϸ�e{����ƿeO�rJG�����w˶�{���������t�5�@u<��d����1�_�B�q���û�*��2��r����w�tO��G��>�ȂPn&��M7@TZ��7��_�P�t�e)�S�����K*�_��&^hNP��~����e����ze�#u"�5>�چ��_\J��11�;:&8A.�\�����
�A��ӨHC7tm���+o���E��Ґܖ<U�n�?���5�k�=|mz0��+ٌ�Y����.���oGVrJ�8A��g]q�2=_-�V>7��V5�7�2�%���vhmM��b�A&wGNgF}�u�s�?T��w���Q�w"�~�����_lĦ{"�F>F׏��M^_�����I�G�<�_uC����� �s�G��w�ˑP���<�|�Ƙ=>�IF�u����R����:�:�ʎ�p�ĺ�s���'�:y��W�ӡ3p�r7n�%��,]�a���n}���j���û���*�X���n���s�S�;�;B��.$��$͸�抉�uA�Y���V!��ZEBA֗9*:��j;j����׼��*�,�L59��g9f�*�yܓN{pUd�2*�_ة���&kj�x{Μ��&��J����s�W+o�=ު�F�1~�������D�r�.�y/i�ϖR�\aT�u�
�|_���r�L�S64�P������z��ﲠSyc�����\�Y�؜�k�b`i�$��'zd��H)8fW�Ϧsas�����Ȇ��S�sʍ�eO�^B�B�n�3�pV�g���h�qT�*2kJ3�� c����`���ƶ/Ճg߿d�~�a�z��9������aM]���։`
CE[�2��˵�����Kr�>0_�.��+8���܈���JF��'�����Ce<�J����g<¹ ���1� �<�Vjӻ�%B����^
��9̮$X���n�4f-����۷���w��;�lЄ�pq�)�PЬ�M��0��uHc����s|���,����Ѫ^�P���Ng\CYjv_H�\�Up�<p79Q`LWz��a���L��sn�=�saO$��ȋ���\eIi������B�Z�0��g����p��"(��7p*���Y���x�:��f�F�-ܬ�׹\.���X�#��!�;��SL��@L��P�T�>���u�6lTNmiXh��0=��y͖_V�'�l�y\�G�N��[�x=��,g�D�V_��������X�fH�Wg�Ҽs6|}}\ĵkō>�E�G�c�/2�κpѱ^����!�F���=�T���s�%���@�=J{����Y��+��V��k��1��{~�hy^`/yfD�d�jQ/��L��ӟV	��}[GC���B�`d�K�îr�;�0S�>�ҕ���zk��ʀ�o0�L�i�=�j�Ӹ�	�D[�E!�=G6�^݇>��Cwà�����Q��l�7��㪬�v���������\2�)��J��<VǑn�2&�|Oj�սg��=���u���vv�ʍ�p��@3��	�e������]�7;�\M_w7nu;�%���ʊ;j�Ң��1�E�K�E�4��Y�p��*��KG0�v���)9��zd�vS	\srө#W �+6-T��+�R��.H�H���J���.��L_��x���]���eX���L�~��<{ÑҨT�푵�}���H^����.�tV��,���z��t�ަ4�Bf�6ڱ�=��Ѝ
�����݆N���gӲ��W\=پ,^µ���`L.�d�{k�\F����	�{�{��g=BC�3�П�m#�w��vv2��秨�k�5�T�� OF,�x��E�J����(˼ٯ5\�R:#����{R�zg=E��U~ɝ����t�:ůW{�DqT�tu"����F�Q~��F񯗛�X%Q���p]``���&���x��^�tw�}	� My�L{fu�x����a~/Ǹ�d����q�m�+#}DS6���c��'�7}�_Z�4̝�`�����.y��	�>_G:�������s�{�8ۿTz��c���^�y�,m��$|q��*�]L��-��%�q�����=ǲ!���3�7wާ��zlTO*�]�P&w\z���*Ģ��؟nU��%����j縰_������YH2�X8��i���y�]�93��ƶ32�:0�TI<�5Ԡ�[���/j� ����Z��3���O+��}\�]^ޞ��,u|������U���Iw��e�z����Ԛ88�l+�N:}�u���M�2���<u�s.���H���V9E�� ZTF}�t.��p�4��ِ�ȣ#����%��������#n� ��S�9���<��W����ܹ&]��Cŋ:%x�EeL��~�ݚ
1c�ûy�n�~�jω�5�L:�mR7�~>��K�_��`T<��q��d�/ÞC���ͷ�sH_R�w�?9ZdV��=�����õ��Ɍ��P*m�=A�Q�u�2'����;�0αV�7m(�p���,��[��%�_k�ki�R�%��]G����^���99ʲ�^��%���B8����_�E�ܪۏn*HG�=ޞki�'���q��2�jѾ�y���*S��0�ÿ���#4���R6Y��Ľ�zss���U������( O�9^�����q��m�*�;^ўU��)rP�ҳ7��7����!~��9y[p��+�9s�Tw�	�ʺ}��� u>�O]�m�x����h����y��8�H�7�:
����vQ��D����v�<:y��4��7���TR����ߧx���7���(�9%���Q{�]��}Cbx�^���7K�v�cL�Z-hU|�dl��hc7!��V������-�Q�f0J�ض��q�JR�S/����f@�hQ�r�X�&�k=�S�+Y\HN1Y�ypX�@�a?X®ք��[]1U���n��r�ф�o.�kqfM�7��owp�#)�W��	��/&w��gȼ���qW�������ƽ�Ő��=Tqjk�㇋:��h����������.n*�
<�~����,/du<,\GK���p�q�g�ę�������52*���De]�c�����^�e��}5��)�*2c�T[u�ܤ�8�d_-g�T����K{և�z�,�˦^�!9�L�=�ekޔ]�_�鱝zSE_���Z�֩��N(�iTu�w�<��=������?W���� 6of'��$]�F�՟�Ş#��7�}�<;Ndl���}���<o�E�L�q�8<�\�*|⼊LT����˳q{㜃 G�Y3�����ӸQ����]u��s��L�����bu�pdY�}f�w�VH_buDDN������:�bi��7�|;�����K���7�9�zY�P�~z��e_o:��^����d���Q-���}�Y����5���\GW�� �뎃�����)�=�y�c8lO�K�{S/�ƪq��U3Q�&�
��*�{NnmC������^��aWzD]Ed�@��{��T�����3,�}�f���T��8�͉����+�{{���Ս��+�lM���b짙����I��27����Bg�o-a�D��e�nt���S��|{@��_v�}5�C6���$�e��,�ݸ��r�J�{�Ž:B�ђ}�t�����#�5��S��U���IG."}�!�ϧ��.3kC�o�.,��0$�c9��O$w%D��<s��lϸ�%S��fs��k�<nʁM���*l�=+1U>ٲ�W��v��ix���4ϰ�8s�g�q`mBw���07�N��}�1=�W<b��b={Ǯ�}
Ǘ��Ȫ��FA����� k����`	���ƶ�Z9����LU�����Q���_�rܩ���E��'�U�Q���&u�'�5R�~�ao�y�6Z���tҁ��G+g�z�q�����D�R�rf(��ü2��X^3�Po�+�pG�qe���s��nv�C)���
iW�W2η�"����(�M��xU=����{�
|��do9�yP�8�H�>���w��^���g�eK/>$6l����՞��_�@>'�{������\��dl��z�5���ӝ|�ǈ�5�w {)���xmw����!{/&SPE.>8%��U#*g̬8\����W���;����m"�#�$k��mf�5�<�FdP�3�&C��e��
(�}����++�>�3�{��#�k{��V'�վ;���k��&��H��\�I�'�*	�7+���K8k�F-��ڽu4h��â�ޡ�7�Fk��g�K���*�Ji����`]d���u~���z�C������}�@A�}^G	h��cܧ��_�ڼ��?t�P<���_b�G���� �����צ�\��Ǧ@^�Ȭ�v�����`�xe�Cw�1D(:4��6��\L�h���V�z]�Ϡ���{,
���.U�SV�ݢ_�d�b��a'����d��8�^���=��U��qζͶ�`q��-�����=V.�����+�-���2d.�l4� ��	��|4��i��B��w�����G���Z=��X���Z>�E��T�F�����l�9���ٳ�;¦��ːQ���;�;�z�}Z�w��K9�'������rP+�H�sg�q�ͬ����i�r�㩁0��/ex#�����^��"��l��}z$_��Mh��Mw��0�ʨxk+j�z����@�}R<7'��B�%�^��y�C�9>���|U?V�'Hh���Cl�s��HiS!���w�g}-<
ޙ#�Y#��(��:��&P�N�Z<�����׵�
�*��tE0��L�
>��!��6�gߪ�W��_	|�)Ji ��I��gr�u��7���RAI�aJF<�+�zj�3j���������X��u���&��̙���G����\���[Y,��bOY"[�Ȱqv��Ԃޗ=�;��|Gz;2{�x8��}�X��������}X���u��.sM�"B����W�a]i��F��4�,"���2U��a%n��ι��/���#��+��b�z�]��ˏ'FWf�e��Qo�	�R�9r�N;t�k����}x�/]��"ʸ���ֽjY��,R�����+lW^�薴)b�ۤ���k=b�7����#����wƂ!�wz��ʿ��R�צ���8 -�j����*3mȊ
��ww/l��[��*^�� %jY�`B��4�w�H��T��ǻ]ıM�b�}�W4��m�`�7[����)W�XY�Ǝ&9S�v���c��zio��S���iN�����)�5X���c,b��y��ϱy_���t]S�hR���1𵝀sՋ���X�%o��������ܩ��z�U�˃�����a���7oi:�r�ۇv[��R6��/�,�*-Of�4r@+�`w�Еcoc���vk�Y3&.>����%�y6�5˥N�6�f�2� 7Q����m��K��;�ۃ%�u��N�
�a�ҝg)�(�=܅Ō��<dЙ=dCm-G7z�;�{��H+kV�m��ۗOӨ9q';���ڮ)���!�m���\�^��bV��Fy�c���K�
+W*��feK�]����#�����+n�u�{�oI~{����+|�l$�o(�8l$o�<g!VlF9u��G�R��z�L�gy���V��[�)��,�������g��~ul����cf�c���޶�3bC8����}p�9rcn���ZkQ䴚�ӷ[��[��bϯ9�$%c�(*�l|Բ1[:�k�H^��K�lv4Dk��+�g.�}��f.��9�vD�l��Q���1��v6|Y�"�`��4G�]�z�_J��F��mN|�V�K@)�D$�ع��N�f����z+�t1v8܇r�!����.����1�U���۬�G/8L��a��A���"����.�Y�ZW5g˗f��|���6t��V�����Gk*m�f%̔����SG�d�]�{s��8Y�[�w��B��7�Һ���9�:R�i9Bc��'���zPK��+W�=�����(�;�i�)�]��dM���Y��4EM&! $l��m��F�bxٱ�vd��!�\�]����϶�^�{\�rG3(�c�=�A���YǕ~�䔢H�g+h��T��p��IG9�%Y2�N(\ݷ
�Ln$\5���:C۽v�Nh�n����K�oK�k����:v���5C4��M!J�>�3�T��"�	�J�=���^����Sv�����a��w�S����c���:Ԭ	_v<:��K��P�>� |��n��u�gv��S:Q�ˮ�1(�wN� #ۧr�J��9�e�r��.�!3�������9u�NvWw&�ݺ���nK.��	c\݊WC\��]ێ��g�&(��������u�RI��awN�s���q����N�쳛�Y,�&����w]�2	��Й$�A@a�Fgw1bF'wS�]@Nv��#�L� Q�9�Ý��3��\��˝�	��u�s����,�7]�2I$�]��0˕���w!�9\������)۳Lb��C��S�ws�5�wb�4�����wws���wu�\ӻhW.C�\؜�1]�r�9tN�(�K9�w\�]�wG]�ݤM��ݸ}DU I�\�S�B���-�q2��;T��]8`��,-� �%�>Be܋<�*�{P-罨�ϡ	�g�{R�z�d�72�wk����2Ӝ�!��.��!�_�G��^_Tkj�*�7�"�fA����gv���4A��s:���Qr�b�ɖϲ#�`w�_9�[�����[�nk��=��C�Y�P��r�/.�Vl�@>Ȫ�u-�*ԯ[,%k����1~�<���:>��Y����:�z �h���*�X+�C ���϶�������;�ul�V�|FMz�?�T�<��%K��P����<�#�t���22���� 4s8�2.n糆kЧƳXW���wTx����9<
�z�߷.@�yNH>t<X��v⺈Ƭ`��>ܗ�s�<�����ð���^�&=I��9g<}'>���~��y�� ����|ȋܫǰ��'	���Pi{�m��r�Ȩ��ׇg����T>S驍���<䊁���|.�կ���b�僝I��sN��.�Vѓ��j5΃5Lz��,W˨���O�O����P����Q�~��~
�g��=AC��nEV�=�T��\b�����iW�d�ӧ= �(̑���z� ���2�����	�ک���X�<���=���M�2�^ڽ���]������4�xi}���[MQ�[KW@q�rq56�u�����I�l=�Y."��<�1��-����)^�-~e�{�7�:�H�ADuJve�9ڲ���t�����ؾ\��HǊ�o\�. ��
ླྀhd,�q�U�����>�B�=6w��>H�d�v���Q��x���ې��U��� ���ݦg��Ek5ۋ:�����X�m7>yӣ@Οqp6���g��'Q�n9�&�7�s��ڞ<=98
LG�l���\fJ)@.�a�;茙�Lk!9Q�G����*iϨ��q�{�����c�+��9ʬ+����)�	*R�G�b��l�qZHK�ƽ�!�ב�W���9�f
2�{|���^�u�a_��T��.q34�D��)���a{:�/���C��:9{��cWu�q�Z=����JVp����,�5��)�+&�=�����/X�o�W�{J�3��u{���~� �e��%�����9FFT�p,��r�W�StgU�j�c�T�"���;¯xTzߩ#e��g}�:*=��ёe����lĶz}�/���}����d��q��C2GO�̄[�c�ʛ��Qϟ��w�ˑP�� mqy��}v^��n�V ��X�WÊ����L��:1_q�K�K�58�$]���G(�x���Lk2{����=M�gJ�L�WQIX�6��%�s;4��[�wl�:��a��\��3'�Rtyr�;0����Sۑ�M��bQ��!��SO�p�u��啝r-��(3�,�����WY1q�-�9!Ǯu��A�b}�|QV鶮�/�c�rۙ z"=Sޛ&%���|;�KP��b�z�������>���3Ol��m�5nsK��]Ļ����l�M�U�p��=ټ0�3��j4�>����5��9v]�W��R��dzǱ���� rB�nr�Us<h�@v��8=��v��ћ^���=�Fޠ��^��[wQ�+��2��ׁ�p�U���7މ(����Zn}��m�(g�l���-xj�~B�����ٟG������ޟiO�Pj#ʊ5�~�'���W��qs������6��FMiw��i��#}7Ł��w���05:�)��v�M;��q)��1t4zhA�lC�R�g��F�Lf���L���@�q�#�}L1I���]-���=�9f�J�AY|7�?m�c7�n=R���Q�5�鋌��p���R��T��ڧÝؼw�L�n�{�y��x+�Yhh~�(r��)�Ĺ����Q`Mw���D׃
x��٫2��7��A��H��z�HAm���Um&�q(pP�z�,u���+Ζ�m�ӚV���E��vQM/)m
������|��n{���=Z�J��~�[k�	5��f�����M� ���^�S�W�8d(��W�3�����"���ˎ(�z:϶���?������n�[�J��k�M@=�ݩ���ER�_&�5��=�O���s����H�>���r#}/�����VT��l�ٚ���etX�|<�!9>�d����*.W����aU�hv�������(ѨU��ǔ��,�D�a��ָ�죃�tO#��/&W�ßAr�sO�W���D��3��E�#VTv��ztNf{v��C�5��ϳ"E}�7>��7����������,y��F�=Q����-���ZX)�ٯ]�}9^����n�E<�M��T��L���"�LW��
���=M
����v5Њ��\9>����M3n}@{�� .�~� ��H*��܊����۴C�V���ͩ��Z��|y�����.4rRcի�l�~�<�|������S�ɺ�\]�m-��f���h�{�1d��FN�5���d�c����*�����'Q�z�G��r�'窡%�.&���G��~y�R��=^�nV�\d�7�5�����\xZ�א9ώ�D�o\zH�P	U�Z�0sp��;X���.�γf�syu�z�E8V٥zW(�y�f���b?�4r��}4�P�ݬ��������e�*{6��K(tf���S|��5��Ymr�d�3O�%��::
��0��(̎S
�:%�S=#����b��/�k��I�.3�n'�q����,^l֛� o���+j�R���d��>�f�`p5���l��Y*nB����
�Y��*��+)Tz��[b�x̯S
�nhs����n��Li�%葾ޠ+�m�WD{��_�{hp�a�cږ{>�Uhҧ(������eћ0]��ھ�Gpi�p�ؽ%��jU���W�7�����r��\c�)\X+3�weU�M%W���ཙqv�^�b�}Kǁ�.��"���v=��.iTf��,�]'���Oyt�������R��2����t݀���E�>�/3�N�J��h�qⰯ��#y{�NT�t{D
����8�n��u8�R�B7!ĺ#� 7�ET���[ Z+�҈�a_�K�o�����p5�����=R󎾒1�wz
�M���[��@{�UH�_D�U�%���6�����Sy�z�da���J5�q^�4=>�3�}��y��~��P�r�G��hyN{7�R����?;�P�g ���Uk�E�DW�g�ơwT;�����{Հ��r)�S�/�:,_�D�V�����&*@�@�i��S��E/٪�h����\R�QE��(C�;���]"����-nm?�x���H�����1ê`ha�,\W�����^�=�����B�h�;DT�H�9Ss�aΥT�pZ��Oa�3ލB\���M6�H��s�x�%=�r�wN|O����lB}v�|��|}'b}���&=�˪"g�mq�Q/ˌ��h1�*�{�̶}�D++L��N���)���o�<�>u9��8�.uWQ��;�;�D���gWc��Ue�X�!�t����jz]q�X��Q�Ǽ*帺�@31{�|�Kg��Uε���wX��m���{yIw�^��<�� *�:�Ú*��M^��ϮNS�BuG��|��E�sB�u�/~.����ۆ��1�UHs��D�]㘐c.�vGvE3EO��p~}~�-9��|%��ۑ~���m��Q[3�4ܾ�1B��#�ۿlxL
�q^ާf�4���G@ڎt'7�;	�o�z�����*3�*���8��F�55k�D��G?��UFC�0���{����@��n����i������jP���T�ZIFw���)K��T��=���γ�����	����>���,
����F��Tğf�
�\,mY��ϗ�S7.q�9�U�G��S*2e��e�J���KO��r!�,��F���"`io����T�mw�����v���Ĩ
��bKG�������^�Au�1|o8���GL�ա�T�XN���J��9�>�n/,yޫ'B���M*����u�b�`ظs�{�$��*us��0���YN��RU���{��j�:����n���n��C�A�+����>��.X�j.7 e�^3�X�i����*����C���;��χ�#oD�wg���^���/"U]��-��e##�2�tJ��=���jgW�{]oYPѨ��K��_�GYq�����E��W���L�ټ�1cEL�Q���ߒ ُ4w�22�'k���i��~5��y-_���+�F�~����ܹ��e���#N�c���J�Qѝ�of%t��S��ѐ}+N��Tw���]u��s��L���}�=Y2���>��ce�ZW�	��O��5� ���Q��u���U�u�i����U�����&iEC�����`B}�}z���"��@�����J�6rۤ�e�;�^���/�/O�F��<�#�"�M$�ؑﲄ��3(�~�<����H�z(�g���*�Z�Tz��ֻ�]�{�sJ��^�}�q3[P���w^�]�##�xr9�U®�f��%�U���LOE���S���#��Vry�H��F��W�=p�����w��n7�Pk��(�������N�9�hz��y�U,��^V'u�jtFtZ��,��#x������h���$�9��I[[ɣN,Y
��͗9]e�\���b]�6mG��*v_eC6������
�[{,E��!���SyY��6�4�ݸ�8v��{,՝�h����<�J�D�؋�ԷkfaYӸ[��|?R�\2.�E�OK^�<�~R��w<�_\�=0-7~�>�
<<'��os�EJN7��F2��7>��,����ɭ,^L�ƹ]��#�u0r��̹c��%V��s�,���z/�G_���ʔb�H��S�.��U,,��o&|�g�/? 6��֘�dO�P��԰�<�{Ƿ����Wh1���\=�6�>���D�@OJ�S�p���V�ZI��V��^�8NϢ:�}U{��W�s��~\C�V�W2���N�sLҫ;�Z�8�݃��kw�ts.;��^g~�ţ޹���F�S������ĿW��Yt��8���9�3}�<��>�n�k*�Y��2�3�k>�a_N�П��AW3��6>u�{�G�{����M	��������?�����mu�[�<��Y��8;)s���I9G�Q������s�T���Dw����,�)��"Pe�y�9�%�J�A��,���;��7aE�h�����Ͻ9L����w5�zn�J�����z�LS��=�73r{�;}[U���4�Ei�U�o��"�v������T�Ʈ,U4�9<�=���?N�$r���1FI�tl�eķ�ñ)7_��V�S/^�.��|��P�c�c�;�hҍ;-�c��E�3�
R�2d����v*��}�j��Y��(y��,�@��u�~�X���)+�*j�c��O�L6��\4�	��:rO���G�ê�í^�f���rU`�3�|���.�W���;��d?tv�1��z}T�[T޻�>>y�c3k�=�o�N׻f�za�	��ުcν�7�6	=sw�Ĝn���l�|�|��=?��d�\d�7�k���m0:}Q�q�{措>끸�utU3�z�f$�\w�nX0E�k���q>���O��۳|X�3�=ﺘ���Z5�/�y�
9Bj���[~'�o��M��y�/i��>��VET<Q�,u�pLnJ�6��q�:s�;��R�^�&):�V���\y��;�i�Գ�>�T�1R�������oR"���/�������,m���}jy{~����^ל6#�<��tE7�2(�E��E=�Dg� W��	�u��W�;&|�9�i��u�+��������V�7j+k�gx	�ȩ�x���ܲ�Q�z� �*�	��EEϑc	l�G:���2�ё����cR�c��ξ0fC%��
N�L[��ǂ�la�{ݫ�l�슦��:�� #�_Թ�d�[ܕ�=�*n�[Sv:A��|��6�"��[�S�0=�L����.�y��4�w
��\�8��ZG�f�r��rÕJU�-���"WNJ��u�X�#��a�.�ynd&˗B�Pc�f���f������nB�W�\���U������^sY,*�s���pN3�㩎����~�
��\�;� d���!������6Ksge@}�UH�R�V.	||���/&���sT�{н�ed쿥z�9�m ^{���w@?x�5��s{2>��������<[��/8�����{��	�3P��m_���� >�&�:"��·�����nn��p�ѪD�K�	�YBLE#�,��	�5�Oj�ng<}$����	ϲ6�޸���ʅ��U�@y�ȉylvܑ���i�Z�|z���õ>ۘm�����ݜ�N�Q&�O�V��3����*Ϥ������r�����}k��]g��c��2K}ʤ&��gb�#�Ĝ�,�K�jS��W5�EuCණn⤄z�=��4��<�J�q����2 �__[�K"�6}�_���t���lW��<w>��v��q�9��|��9��y�t��d�[:;�ϣ��%S�+��br=���O2���r{�j���.�q_V��x==�0��49Q/�gP�b�^��jOey�$8w9�u��xe�G�+{�s���@�S��1Z��k�WG�_C�o\�Zt�9��֨9xά�V�v�D^�q^Ϲ��
���`���w���'0M�
6�ԳGu'��T;�˩ZG<|��ē��+�^��Y�Ĕ%<�Z��F��[��'QÜgzO!Ne�銈	��D�ŉ]AD򥌥����ڴ�(�vEK�'a��{�Q��l�AI����Dئ[�_d<��MDR���+�vv�DT�.��䷃�:�v�}���g9G\ٲ��F�4\�H\S6���RLq\�I��($.��4�v
�Н�{S��$�.��Uu��ܴ����v�SzFPq
��Ա�k>CC�Y,���m+�Z.�cz]KW\�������m% ��J��)]7̅�Ns�N������~mYs9^*���:�k8	Bgi����@:��1|-^	�{�[� 6�3�<o0t�e�)H���$nL��6&�v�3�/�J4�Ŕ�+Ɩh�sQ��L�8��V�n�.����- h�p�}Z�bH֙2�L��~}�g2�)�'Qp�x�.L�J�Μ��\+0�>�1eq�}�����l�k�Lf�Ω���UeɝN�!�be�tl�l�R�*˜e�:�c��\��Y� �`���h��|���:���}���Z2��Ƹ>�krHr�2��L4����~��w�̯�[��siاxB{�mi��L�b�[��r�)�-���Y�aXbb�5o�~j3��\{�x�����k�M��r�iUe���Õ�!�R;)�	�:�k��7���DmLyn'f�Xb�� `�/.T�YWZ�Z��0G�"+�9ڻI
�͖��i	�� �����c����;V��(-n�h�o�N�K�7k6�Iԋ�N�|��|�c{��R�%g`��D0VkU���X����4Y-M��^�;�9�����2�7���Uo;+�qm���ڻU��.ac�rSy����
h� �9W�.fd�r��M�����z9����b�h�R�;���&�3��/�i���
�0����{�:�.�P>��{v�A!���%��pJ�PY��
�U�$�:e��s�A	�2u�Vʈ�%��}4p(F�ӳ5uZ��V��X�jp=s��F����fGi�u�.up���r\ĳ\�J�
�{��o�[�e�tzd�����\ݔr�ӥx�Ɯ�=a
m^����wI�Y}���Ï�4�J?�9֎+�\�Ұ�3.��0��	���L
�N^Ԋ��XV�/�}�<vD�Y<v���w\z�$y���8����t��T�z6��a֋�Ra��y�)��a=����.�urD=��7��Ax<�	=v�U�N�`��n��;ws�u�i�F��w]�]�$�'3�L�3�rk�ܒF	����p�E�] &D�u˒����Fw\�)�#H�(��
Ks��ĳ"Fr����ġ.�!]ۮ��2��BKr���L�#�Q�ȑ 1�����]��S�E"n�l��r�P�h0�4f�wut����]8Iλ�	�]��F�4��1wu �LYΤ�䰒a#;�2)�wt� �B�s��9�srb�d�;p�.�2�t�D��]��)���\K0���B+�����E�%" �n��Y)F3!��AAJHw#!�I�۴�@�5+�� �����47.�1�:�d�#s���D��dċ�I2R�H�Ww%+�)�ܰf �\��&E�I�wq�u���t�,��32v9z�8	����7�Z�����!�b�+�T���R��~x�q7��KՓ��TA���J�tR�2"Ψ�p�Hξܽ��qgm{��Y�sz}|o��m}�:b+���3���1���R'�Q��ǯ���c�TL_��VҐ�*�*� ��lB��Z�����M9�����y��t���'9��{�h�c7м�nY��N�l������,��N3d��}2��׼p_�o��9ݦ��o��v�WmJ�z�rPb7=Ʃ'sqU�LT� U�S8Kۋ�^.$���<�]��},��]`z
Ӿ���n] �V]F���}se��D�\
n@m��(���0o_��'Xg�1���wp�$m���#�z��L��75�@{�`ë��Pq=�O�O�S\H��ہQs�ˬ��h�_uC�~���(�.=�tU���~���xf/T�9Xf�������}�LKg�"�FTD�h�@,-9����e�~�pNq(�C��_ )��m�Q��kЗ�|�* ��2 @�� �x�
r<�Ȑ�W�ޮ��]n`�:��Y;�Q��k�j*�gH��L�Ǟd�a�D�TKDz�=��	����h޹������u�,GcD�l��f3r�vF:��%Z�)׆y5)NP���o!��V���جQE#�!d}��W2�f02��l�M(��-Q|��R�K�-d��ʊ���a-���wb�U��6u[37�~'�*�v�e���H�R���&���̄��U���i�Q�v�_n�	�
\^m_g}r��!L���<隉Q�A��5wY
���:�>����)l���N��{+�� ����Y��@yd9���H�����x.���`�����o���q�w�9އ����=���xZ�d\F��<o_��{bNپ�IG���)�Y��n�88�d,�.�
�nr����N�:����B��ʁda�b�L�.�\u�H�c��� 4,�JhM�4�^5��\����XP���U�����ˀ+�/sk6+*t�|�m�ﲧ�r���9�udU1��ZX��g|n5��G�cG��s��@��ly�^��u;�5F��{/���m�1c�M��T�=��]1��+b��&bO�G��섐�^����jB�]��j��l_��[��6�|�%>�Nm��Nrj0�d�����S�O�f�&��&J���3�73�s�aTi��w�'�{>�W��xYYR�~�%��^#YWD_�"����Q�&�\
�I��ڜ�eC��"�}'Ǹ�o��U�r�V�{�aU.�g�vf h+�Μ2{��1O�u�G�)�Xr"j���.�ū)n�G9��Yhq��'��}��M!8�f&�uu%W�<mt��:
h˫��K�VU�\0�q�a���R��H
4m��},�[+s�!LQ�9o^�a�oq�V���M��}ڢ���Y�|:H�l�@>Ϫ�Yr�˔ϙ��aT^��x�M��I��fc�Er�cs��vթ�X^<}�q�*O��pKF�:%��$^}2�V.W�fς��e�QR���^�9���ݕ�8=vtc�eϣ} k�ndH�yNnG�O����dEPe�y9���f]Ȩ�f���'�M�W�j�M����X��\&#��n)�G�@�)��1g��,���{;���|�F8'9�_�0��b|*!>�g>s�ݟZ W�e��TĪ+�Z�"nƏY��V�a�ޙ#�*S��O�/ԈR�t6>���*�W{'C~�
6�X�ǽ;`v7��҄H���~�����GXx��?��*��J^��}(Hz_UT{#����x��K�x��Ą߱4�@��3��*���#ţ��x��{g4��'Ei��*�ɍ�p���%�骪��w��Ԋ��-Z=8�46n#�͘�k�+���q�e��HޏODb4���|GW�[��bо�#�H�� S綀ϹבY�&S�rW��
�Y����
�U�T=М�&����ɨ��˟JW�A��}�a�O�,ͮ�yY�^|�Gd!�{���%�/�("�����Y�|s�֌����5;C�;�q����x�O��ķ	+��������yzȂ�=.0�>�^��8���SdV��;�C�t����3y�I�x��=�����C���3tKs�CJ��XS�}���Xv�o�Yh@���k���w��}3q�,m�k�����Q�lG5���ʇ��o9��y#�w�&1�|��������s4E�xJs3���Ck�)���\r=��c�6̵0��������^��e���L��Hn*�	��DT\�/&[>��X��Z:'�)g�W`���깼|d_�N���=W�`YR�vF��f����*�]L�@��J�u�L+[��9[5n��_o�����0z3y߆{��EoOi����VznD����e@��h@�w�l�j�.X��w){u�(�0���P�E�q�/ґ^���G���Q�t/����<�#�t��Ĩ��{��u+�ޏp��Yg�Jgw>��P�_[c <��������t���U���)#Q�Y��>�ϖ��pz ��6�n���+�d��C `��=��U��-�F���L���7=�"��M\�Nz'ж����g�,/-���b(n5�[�=9QSQ���F��uñW!f���/��a���w1w%O�#:�<A�Qԛ��W��������dh�F[�\�!͔]�Iu�u�q8��x|�.o��X��X=�Y��>� ��w�P{φ)t��"��ݵ���i��Fl�iC�\�(ФM��`I؆c9��Y3Dy���.��.��s9R��]#�k�~����_��G�S"8��lˏ$o��"��f�z}V��MSȝu��:�į\���E\_��|+��>�&i��]B��r������E�H��,���Es��y �躍�R���z�����T4_��j�z	FϤq�>�ir�P�X�5�ӛá���|����x��u ��qq
�[��	�VV���W������w��2W�N>��g��>���[p���tp0/ӱ\�T��g�Bs���$��412g����K���_.����{�GQ�]�NUFC�Jf.��R^_��~���e��9��c��*�Q���@g�>�-�W��7⤤TK��VUE��x�q�:��^�YY�����Fk�\Y*]���'�|6�hw�:�dy�3cH�J�ENUXS�1__�2o3�:9����]�G_�[�:}���x�����G�튣q�~�y��I��@K"j.^ ���/}5W^��[��^t�>�1�:�0��]$r	��L`��=~d�-@�-�qf�GMN{�L�vE�� ������� ��(�1�-�s�wx��������u�t��|iZ=�(, ���b�p�Yj���2Jְ�fM�a�$z�%\�w����T}w���iv�Ea�Qd�
�Ҷ_nI���ʥ��ޠ��tȰ�3��,��\�z}[0�W��^�����<��	w��@#����<l���8�{��Nz�hG#�3�H�}Ơ!�6��~5}��__�ǽ9ģ�ܢ���2����'�6���U_�/˲�W�ʧF.<�|��Ġ�"*��g�pi=� !���\= ũ�hM���^.u.�4�["<ʐ�����5T@P#�=��ՓO�h���úu��v6;8�����&Ư��]K�<2eCwq W�ب����Y�ך�z�����������m.� �r}���U�R�����PY��o��v�h�d����is�z�%�UP�7&;�Fm1_izL�����b�UO�ƹ�<_�p{��6y�]��{Q0&�@��ly��ǎ���UI�7.p5���q��Q�b7;��gY�_��u1��R����z���������C6_\e�ޕ��p�鿸�&�B>��h�MˏV�Db�7�˩r9�U��MY��x)!����*�r�!��w�Yz�ӵbV{���@tJ���"�7&�I'��5X>}�V!�l�Uio����ϯ�ݰ�w��!�5����q���T ���Ŭ��pʳo�1��[5*m��K4�Փ�R��h�R]7��n�"�n��,u1yN��g<��]����oE�z�G��UԷ��r;�ϩ������^O�=�b6߭��ǧ�ΐގ�ܣ�M1q�Wd��u�/꽏�r�c6׊������)X�����~��qާ��Ʃ���_�:�{-�eO���u8�|��{yn���GѠn:���e��dς��0�4���D{ҼR��{ B�ڨ�k�Y�X�mu9�sˎW�n����L�T���J���9}�x�O$��3�)B
�Ӫ�A�f��SR;<�zz���Cfϕ �*�]K�E�Fo%�N��'�lC���;^r��%�}R�ˇ�`���<����Ge�$Q+�YE��̄cC�D�}��#��R�}���v�,dy�.n=�t��˨�Q�S�����of%�U���"ql��xLy�����u�3��(�n�@��q����8�+�����w�̉(�
�hߦ@^�g��{���9u*78������ѣ�̃�{�>�i|�|'n �{,��2=�i/M��a{����3��dՆ7>ݢ:�Vɭ>�����Ba�%�6m�PG��s����)k%Fi�W�U��m�c.eC,���V�{r���~�j��sv���6m��ɻk��
�.�}��"����M��8�Y��_���6١�&kD��%�t��C��]��έ�%e�}'WM�k�?ô�K�v:U�~)�/)<>�7^���1]9��u�./7N9��1�G��U®#ʢc���9���=�]�i�;g�7��3_m04g_��Ua{<P��W#�c�')�KN��m:�F�� m�c^���A���j�U�:o�F��P���G���Ѡ��Hc��^��^���i�x���ymX�����xa>"�)�vF�W��26��8���+��N�������r}I�{�[��pW{hE�o��M�yQ�ֻ#�hU\)4�3�tqqCFTeT*��q���������>��]F"��w��͎�t�ϸ��^(�K��e�C��������M�+ҭ/q/s��L�����_��ᛵu�ǡW�Fn��OB�uLa��W<՟��MxX{�U`LT�"��ȱy2ǯUXY�M�};;7�+c��W-t��Cl��;�>�r�,�fÉth�P	�ET\�-�*ԯY�𪄴�$�4��5Ez��O������q�u���#�r%	�_�����d�F��?ۘU����'�V�b� ��S����̵%����.]X��v-�=�ׯkL���)�=�W5����=@SԸ�fr9���R�y���%��]�V�xne��
�ہl���;wDrwƳm�Z+8V>!pJ�s�7�ɭڀ�F�q�t�O�vr�ܤ�ۣx,:�G�;�,��j���/ԑ�+�z���T�'Yb���a�ѭս�KbgM�r��J�>V̂4��Y��	�Go�}^�G�\
���4?mԋ����p�n�H&y�WУ"S�#��<X��P��n��S���wNA/wz�ϦY��I�{��<��a�����kiR�	��z�n��RG���nQ;���ǰ2�P�k���cӵ�����s7��aw�/�G�T�����Ϥ�©�=�Me����/�I���j�}N�5�\�!��^�>���k�y�4�4�!��k���߫�����0�;�q]$*����3��X+����gѵOS�]U,��^'���h��{MX��IG.}A�v��5<SW�w�y�^���ܘU�Xn0���@>��Kվ#>���xd<�3P�M)�} ����3G��W�n�K����*�.��!�n�q7P�.�D�Bڙ?V���;���m��3N�;�b�8/�Y��	�A�s��^�Y5��;�d2�L�e�
����=�g|q1ttm�TI�u�޸����M0i��x5��DN<蒨H�;�tj�M��S�i,փ�}c(O�j��b�p�K:S&g=�=�����q�qt�
��t����ѩ�|_�;��.	�Xp����;%����JDr��U� �J��?��x���	������LU�M��a/��u�1��5;���=�
����7Լrr�ae�z.:��6��m�zj�\9ÎU\������I������|d�3��Ώ{":�.:_�F{��{=��Nj�c���9�L����
3O1{�mU�P�}гh��{.5��t���]FKt�҆�<C�ɌW�p]ړ��D���(>�2.��+�g��Rچ�}}0�?ZG!�J<�}���ߪ;eEM�јWw�IUT��D��%�4�gLgz�F�5�/ƾ��r��
��gH2T��O�~�r8�H�}��+#����F/�'�7����g�s�:2	�9p
UjQ���c�*ϼ�8�>��>�[��d����o�q4�k�@��TK�p���`E{J�MYh:�ϡ̮��f�1E_�U�L\ڤK��7׬ONG���]�|j:�VD��=����1�Q��
�E(�!��d�a�.�X�������� {��j�x㝠�g��������'_� �����۸��.���ћw�>�
�v�Tn%�ۅ�WT�dv@v�CG���0��q���ǉ������y;፡6�`�TCN�Ք�Sk�з����fnɀ-�&��tĎop�5=N�)�`�p@�L����j#S�';�47q��^���N�m���h�H�p t��`�0<��r��"��j_�u]�xK�L]�{ʶⷈjn�y�v��gr���Hht"�}&+�e굗����u+n���9�%K	����k��|&���v��KM<���k�גPA��㥬v_ݹ���onSf����7t�a��CR�v*�����NCKQ�zXM�����g�Q޻���=ٚ�W�f!m}�s7~�q�i*���S�B9�U����,�[#e�If�*�iʹt�&5��*���J�9ocC8��/r��������Ϫہ쨭���y�D��2��=Di��� �0���S��*YRV�(&����xK����{u��Nu�F��B����%.ti��3ZoE���ռo�W�pi�󳹌��{E̐�w�n�ahԘ�(ѽ�uY���0r�F���O}u������ޯ�o"0�}�gbᗟ\��	��8{�ÑS�1�w��]�Q(@{�V���'M���qh����Xs[cG\��Q�+z�PYp�r�`���t��jb
�xE�T_]��
���}n���*K����n��{�\��i*��:̂�vy����uЬc_�n	��ǫ���
��)GYY&�uE�\C���+�p��v�����'�yj�΁-kck��5CWu7F,�yq�c ��,C��y���1}uӻa�\	��qH�Jgt�CiU�����
\�^�2vG$�e�^Q��Y�UB�q�;���4�`�E0"��Y�h%*��ٶ	�vpk.=KED�hk�N�+)�tu�5�����g�Y�k�:V�A����u3A�2��+��ǡˮX����z8��nbh>�ۘK��d��^*
�y�n�'W-�u�� ��͙r9F��β���':�BXn�� ]ɮ�S�7θ����E�,� +�9�c&d<Z˰�X\9�w�cpu&DTN�8�86�������G#}N�M�bv�s��&�k9u�5rƪ���u�S��J�k-���l����6zM꾪����68�4�
���w�!e���9PΫ.c��Ulv�' e�G=t+��P�W|��6Er}\��%{��o�����)0\�u#\�n��;;�[����l�R6� W0�s�EeLa�л��}ٌ��c�é]W�>�`�>ȶx�돱R������ЫQm)݋sO,5�T�B!R��<�{ӻ<}��,<ڸ��Y��0�w6�w�J>M{x&���(��.�*�M�I�I��G5b�V�I�8�N��v�w�9�.�ݫ.¬g)�rی9}�S�5����r�m]AQ읂L�J�\@!{&��T����<�]6EXS���E���"�2ͷ
�D�T��*�AQ.�'��k�{�\~�]�`
3�}�ك7@� 4b`w]�wn�2@�2ur s�"�LR�a)Ι�)�wS�A9�#�����':���aBJ��Nq��HMJR)����2J��"�N�ٰ�����$�i(
.�r���s�����e0�.ɔ�a+�Έ�f��A2�� ̤��2)���3,4Bnn�I4Đ��)&%���`�Le����!Q#H�˄�4���#
(QA��P�`�)K��E�.\`�2s�cJE��I���Ewtb��(d��1s��[��#d�1&n놃b&
�9Ɉ1�F�Z���� 
���ј%�]]K�M��NV������kSQGV O*�9=s3=Y=.|j�=�Z�Fn���;��	W�G4y4f�>��_�i
��o&:�XZ^�5P�j;3-��g��qp���\W�|�Sgui���}B0{��IEO����O�(���"�+��K����w�x��Ȯw-�GHN85t㡛}� ���`7Tx�;�N���JO��.2oJ��
Ӭ���`[윎�N��F<��yy��L�z��r9�F�&�*b�=�V ���'��!������a���.|_�Vx^ʐ��W�ަ�ϡ�S��t����!^����<���Lnɡ
�7�;طg�I�Z%��༢:�1��xo����Q�=�4dy	C��S��ړ}[qY�d.�!س����c�7�,/�0�J�x��x�?���������b�d���2/X��Q5���Q�`=��8)�'ܧ��!/O/eD�	��6�<��u�env������<�}s^=�ٯ�� ����? �.��V�l��{=΃�]�V��AdfS�:�%M;�!��p�N�z��χ��E���W�e�S7_�v�x�j�|�*`Ѓcxr\2�KY���H�SFo��[��κ&� �;m�Ck8� �|e���`zRW�sS��H��#�Q�j��t�2��3˼Y�P���|�fu��8uy�(��k�s��w$�j̠�\�4�Fa�~�i��k�..+�J����uĮ�2��e>�Cｗq0)y��W�+��<���]�K�^{l�B�7��>�{��	a��cJ��9�+���޾�n�F��5��}�8�8T��z���[���|�VL�oN��+�w>GxO�'�l������t �=�`<�qN���H>8��__K�=*���sX�ݢ=V�d֗��r	xT�!/Y�q���)ߠ���%uxߧ��|��_x��9@R�W���7L.9�VS��ZzxOl��f���B���9�(W?xѭ3m�&Ǧvc�z(����He3����=�5��vF�iw�?���Y�B�q}QE�(O��d��=�U��u���dd�����@��q>���D��=���X.����<��)�h�+�ϹJ=,�4���~|XVI�G����lgOz)w��6�����*����i�z��J����7�^ mqtF�[���V�_G�_
��Э�������k������9�T�L�me+�q��n�Ox^��o����>����$G��gq���ޤ0�W�y���:�;/EX�v��b��[�'F���_=�+�J��G/�m���nI�(Ɛ����Q�b�=�����tq�1�qB]խ�W��ۿ\Ӟ�O_E��:{��l���U�K�s�[��C�6��r��^e͹�KzMT�{.!5C��3�`�)R8�]�d㘲}�}�Cw{��;v�f�]w��.��W�;���>��2��n|^o��f�%�0�*�	���>E��O�2�E)�+٩*�]etN�:��>az4��ў�����S�W>*Y�ȏz+�nt�>�l����>nv9�Pf��9^���q�3��!9�^���Dm��p�
��0KF��}ܶ��P�����H�����e��mCU]ŋ�~��G��<��Y+�e��?W���]��/�ѵ�l��Yat�2d�s�22�[���^L?i+����M�S��x�)�bq�Y�wv1^���������"�!����'�s�;���^������lˮL�z�Cէ�#��c/\H�Ǥ�{h?eȨyU� ����O��;nH�V_��`,c��edmuuO��!�y�ֳ�ސvW̨�������H�tx��ʯ3�eߊ��0~��`~!xC�ڴ�u����OUΌ�%�]F��S���{ӕ*9����mU�5Ta�=��"�WBP�.��s���[�Q�/����F0\7w׳�̌��82��!��8����s4�v�Y���^h�lD��@���)�����%�4.�.�ͫ���D�U꣓b��XD�8��1�ktH�^E����MUE��Ev�j��F�������f����USዪ��q��Ĭ�꡴Z���T��љ���\�tM�?2��{p�}p���ǯ&p�����`	U����d5NO�(�V[��F�':�����oQ9/��V}S<�zDڌ�q�¡H�M�qp6��&)z��T���v5�L#Yy}�m��s>�[Ց9�m�9d��q��,��2�&��'}1��r㌏k��k=w*�W�����z���q>���+� ����Y�g�#�Z�#���W�*��:����ޞ�f�8qs��~���#�߼ty�q�~�x��Q���Q���W�q7\��xj�שl�J��@ץ��|n2e��b���g�W�[���ë�°��~�.]����q�[֘�0/}5b�P�g�&aq�za���#��^	oS*|�~��yO�4���������'T����Q����O��>چ�E��;O����3��	t�E���MdyOkQ6({�:�@;�E{�2f�����eL���^G2 �i�*��˰�zwv��}9Y<��ws��V�PEd*���pXC/_#�����E��)=}��&0���ʻ�u:�X4�M&���l6�a�zEu�܏�Z}���xɳن_.�_r�%�_aƛ/B�N�Y��,�]]�Rg+�����H�S��k���|���4��L3箎���&�=�^��>�������eV4�td+Nح�ڻG�t��`Q-��f��
z��Ü�>����&<�I�D�l�L{na1]\�Q=q�Т��鶱d����GQѻ�)d�T'�l�9�t�K�~�%�^��J�����jx�uzG��\�ָI��#��H4_�^�5�f���4y�@�����S���7R���If;�����l7����0����2) *�1]w^�����kΦF�Q���?a���c�#�{�sQt�㖨Y���J9z���Ț���6��Wx��zdƫyT͏m.�\"��`�E�«zf4;�2��<x�XcX�7�pzU�{nV#�=q�M!/L�0��2#e1>�s�7��' ���ہQ������{�Zʃ��(E�B�Fg슯NTd֖�[�<N{s2�i�^(�O���@�}R�u0�X��k���\C����E���>9��wIC��3�3�G��){��}�mN�FL��z@N��1��z��j��W��e!��h�Ũ��/�_!m�:k�k|6���m�{�+i3}2��6��U/�[D���N�����n'�+���s�����~�%��>ԁ�n�ǒ��1�SR�mA�
�w۷t� U�I�E��Ѱ���͸���y�^��YD]Z�\��Y��sQJ*��d�*pqyQ�M�x
f����r�����+���"7۞=�lNJ�V���dY�Kܦs�/!O�x�}��g�nz�5��_�3цC~��yQ��AbնD=Fv��&���c���/�����VT����vl���*�]}�W)3ZX^�/<��!8�޵'�+�w��x����f}�����'��pSG��ET�����oG�D���3��g��/Ή��Q�}�ë���^E�{i>�Fz��P?W����W�1(>���fn����^��fO�G�=��������|���q/��9�/V��xր�������9 ��@��o��:��}� &�>��>�ӄ��v;;�>�U��r�=8]h{,
6�eX����nd>ͳ3_SÖ3Y.w>��#�j�MDiz}�	xj	�Iz͚�~I-�Ƴq mjK�+�g'{`{<r��}>�5q7����csg��2�^�B�K��i1}U�6,���ۙ���G�����&�N�y�h�C9@T~�!��#�O�{"k�����8?i��N$<z�7\�y�s2����g�{5�����WlpƆ�5��măSx��&�š�R�ƛ,�w^���P��>�����y8���q,<�s�9E����]Fb����:�'�dw}�W;׋��o2�cK����h����N�u,��]���BP({��]h�~�A�Dc�8ߙ�G�Y���k��#8 ������N+������鶌��}�tz7���j���`J�d
�9{o�g:�=o��H���5��{Mw/d{y)��7�i���Fxi�D���q����Jβ{����t����=Z:��v����铙������7.�,'�984���0���3���K����g�n;�#���DJ[*E�ڣT/!��>���^����mJ7�e�K�
��2/�p���1d��9d7����L�u`Q<�{�L�n�o���;��6�Tm���Y����K�a�}U`Q�F\�;���Ϧ*~����5E��7��z����9{��.iT:⨳q�W��j�}�U`?cʡ���u�/cL�Y���.�|zp ��hd>�=��6�=��G�AX]�ȁ�[�����4jfn��>�@"��-�ET�-Pg�_�a���,8��l��g��WC����A���eG����}dr��ِ�Ϩ�ʉ~���^L?�P�%��� �+�Sd�m~��0�5�K'���չE�9�yz!�����mI�����4tY�ႅ].K{vݾ�4��j2�ݙڣ�]�}=����Q����c���[�z,�G�hMaƅ����ύv*�<P��s��Kz����<.�ޥ[����Wu�7�����)��RWL��r=�.���:%3��DӞ��G0�/o�ǥ�=o�b��H��S��§vx�f���?eȧ�^�.%���_�dnQNV��}ǻ�o�C��8a���u�q.�yRc*;iߌd���S�=q��P^u�@R|�lMe�܍���m{a7޺1����}9��.A�C��OV��_q��GwYy��_��S���e��v�!�Y����C���{/�s�I�E纷L+�6��s��}�ǅ|����uT�.5׉�~����t�do�;.���"*<t�r8�W\=9���j���_�M�0����c��o��R:�^=ϼ�7WH���(m=�oM�GNE���b��.W��WJ�����3�������7i���?{|iZ�}1��g<���f��*��{�}q7��獯mH�7��c:���Zx}-,��Vy���ͻʼ�]{0���j�R�K�O�]3�7�p�;(p��:d6Ò8�<���߰Ƶ�����Q�Ӊ��ä�/�2=����=μ�m�����+�~ʔc�kL�K�e�]�^��n`Ҷ#jA���ZU���v����7�z�h�c��n��C ��*�OP�[�k�{�%Ym#:1J4�2����<�[��G�K���Z�i��R�ʵe�{;��9\�D� ��š٬NH��֚�yg!7��-[�rg����{��vG�D� �)�:0��d�w�U�K����#^EyO�=<=�d?aG*+6״V[��q6|*g�s�%�D�\	�:�ҙ����}釡�qo��wd{��owt7�4L�(֯?4Oc�ۂ�hw��[��L�N}FFT�p-K�t���W�P��6}�h���W����m1�:y�G��p��߯�q����h�-���R������>F�VCҩ]#=���1��Q3�O��q�uϸ�-{r�SʧE����ىA�Ee�?E9�w�=�}�7�,�ԁ3�Q���T�'e�8s��=����̉��{j�
G�{��p�϶.�`c�(�d�u���ǭuu��;��e|���R}V�>�������f@��7f����q=8׽��`�L��5�*�#j��4_�^�
��P��u�!�@�_�j���A��������.�<�;z��2o��8��ݨw��5��3[P�i]���|^㾽y�M�N9�`	� x��R��45�-��pki��Y��Y��z_��Q����d;R�z������hf�J� K�V�Zvᢐ�2vN���=5��,d��u��ri϶�ڎm�-�E�y+��Kx���M��Du|�>qG
�A�r�+apҫ���i�\&IICNİ�giUv/��>ݙ_��qs��r��I�W��F4�)��~���|�X�ź�YpzU���b�����M!�w�����Nu����������<�TJ��`g��{�5�6���_4+tdg���ӕQ��p����C�wB*�0��wK�� g��G���6)<�x��{��\O����\Fy
��Ӊ��u�琮I�'%��U��=t���;�g��Hc7��[ӑ�_�ץ���~�'��~u��.��Xt�P�6�p2�&� ��\;�(W�n|�}�0�4���G�/�!��`{U����Mp��ڽ���Բ�7�E6e��z(�\��'=e��|����6�2��r3�=�n�	�i�q��ϴ��^�e��
����@>Ȫ3c��9g�?
�c�.;f�[�Z�Ѫ+�'�{\�~��g�U�s�t�5���՟^����-�� =瘝]V�n��[���ްg��i���s>�aU�pw-ߙc_����F��ۏR��_G�^������5��\��q�q�
'�v?��D�ͮㄴwrØ��(\J��Û����|�����*�����U��m��U��m��Vֵ�궵���յ�m��[Z���umk[o�յ�m��Vֵ���[Z���mk[o��kZ�|�kZ�u[Z���U��m�֭�km�*�ֶ��Vֵ��j������kZ����km�Vֵ����
�2��S��(I�� ���9�>�>���Vն���SJ�5�k&��f�T�T���&KiZ��̩ijiV�4(�L�X�lj�����5��L�bfm�-i����f�35kbU�m�kC$�Ѿ��0gMr+	�lZ��۱���d��Rg[�P���ͫR�M��ܮ��Mj���mm��fUkm�)��l���[SkQYm�os.m�(�M6�Il�)Mi��ڱ�Օmm��E��J����k*���������D�3[&ŭ6m&,e���kA-%�ֵe�m�m��,���ڴR[%��   P�� ����kT�-�5�Q&� �m�����p��ɵ0((�1����N�)U�q�U����6����   U@v׶��R��`Q��ܐ (QEXLQEP�F�PQ�^��B�(��(�{qEQE .zp袊(��(�^�(��(��'^�-���V�Z��eP�G� �@P�g��ցe�R�E�n�ԥP��h(�;Q�h1YuԠWlHhm4	U�,�F���mց�Ķ��e���  ��W�N�AM��8K���-�J�IP�Sq�ںi�am
i�f�t�kV�4���P�j��Vж+lѴ0�T-�۩�])N�l6�l�Y��d��Ѳբ&�#�  Z�Mm�^�ΩJt��w.ƋfI��m�M�#-gw
��R:w)l�ִF���t�����n����:UR�MU��hU����VVPR�T��t6j�6��-�/  ��m�l36��@�U��d�6SJ��1���j���t�䪋f����ڥ-Z�mu��(���\�mWn塛�.��ZRTU[V�-��d<   mq묡�*�V;e4����*���mr��h�Ӝ4���j7-N�lʙ�T`ִHi��l����7��lK i-�Wmfֵ4�3m��b��bW�  �� z��( ,mS��괶�i(
l�uNUs3T��!1CmFٛm`�Z�����";Y�vnԦ����`:t W:uA���j�]TN�j�<   ���a��v�-J����裫�i�s;�m�6��NVR����]m�m��$Rj͙��#u��-���Uwt��m�u���톃Eu���6��Z�բ*�i�KG�  �MkMl6J��4
��ԡTi���wnֶ�Z�t.Ƶhڐ�ZеE�J�iX��UwP5�;un�x��T��� "�ф����@��Hh�  "��	R�  �~#)�U&�0@&�&����4d�T�b1+B�t�H
`$�o�ɦ�E'!����_�~��l���o����$���$�	%��BC�@�$��H@�xB�!������=��~�δ}����OiBk%���c0*����C�D�tE�p���Q`�qTY[`�T�s�jI�����d(6��ʚ���u���y�Y2=���[R�f�jj���FՑcJa6��*��⫛Ie�J�4m۸��J<�M6wHP����ݩ��sm����*��yL�M8�ϰ*	�U�:��j��P�I���[�}*[9@V��H=�:�w�8�`.X��������-Z�4xv���-���TW�,P�Oa�'貹�|X^D���"�87f��oMST�k�hdlh�uzڮG��e=zU�3O�x�[Q
7I
^�4�,����2ʕy05�3e�V&���Bnm�,�;��@������Ǘzfj�����*���V��ۓ/]�����V�Vi>ܞZ�:�Fܐ��nl��Bm�
Qޠ~��R�r��!���7ZQv-0�co^�V�p;��DY���h�����+^��n�d�Y�*M����${���x6�B����r�r� +r�!ch�{�KB�D��PV��b����n��I�\�DY�t����T��y�"t\b�ꄉ�����)��U��/d E4R�b��+̽Ν���R��ͭ��T�,J��;�-�\IL�SM����K�6h�cNa;��X)lhB�1_�C4�-�ͩ�3kYC-5WY�ګ���R�5b�tf�SCE�Ym\�Dn��˭�����`��/�V���1\ ��bk�3A�Z�bZp����wZEm��-;{�� ى,Q� ĭٛw��O
Xn�J�Z>��"sj+z���{��L�u�"tJ��gf�(�Hp<5�Z�3ʽ��b3�X��W@���w����B2I�JcV'��Iz�޷}l"�Fr�o���i���3�(m; A���%�� �)um�e��}�{��~1��F��#ϳ-ǹ#:h!t\9�"l�*���P2��k6���ĭة�7�{#��:i�sf�e,��vI!�Q֚�/%e�b�������+�bIY�p��poջ������؋^.��[Z�-*.�Ӕoe�ܸ�r9��t� �['^zX�%T"p�1���B}��$����Ϭ��cE�z{n��)Z��,��s6�Ô�f��>Lz[/�� �2��z�ɻ�F�n ��Z�i�{tsώ��s�Z�8�c˖\S`�XVī%��h�f�{*�EM9�Jie�:72dN��4I��R��5I�/�rܗK!c�-�p4^])*���;T���(�Z�-l.��{Xع����x���b��9�	I0lwt!�7�S4�wQB`�rMAyF�K�.Ƈ�tӨ�Y��I�;*2��5�"�g��)�c�(^O�<�fXQKwA;V������qeJ�۬D8�ހ���D��8��q��G,�iE&!iʽQ�2��L.�w5�HmZVv^�bcY6V�M��Z���'�{����Q�p��_\��	b ��
ў� Yiʦk��B(3�1H^�^��U�{v��5� ����~�J��i���W�E��V�d�9x�L*z�%�8���"�Ȭ�!Em����ȷl,��yWT)�2�E�i��&��7r�;�^�7MjZʐ�m���kUh���9�c�L��V(!
<uz)���S�i��X��L/=�/o�S��k;��^�B	Q`oeѽ�3kY��8I�E2Nn���Ħ��{���S9L*41[(6��۽���"��F�}&�*��s��A�hVm�����kZS(;�Q2њN�"���'��b�AR� q��,�GB����\����;�o1�g�kwlT�����5���&Lr���Y��cE8&Cn����P�z��x�l��+Dõz�f�$C�1|�8��<ϲ��1��t�DNF�"/ԄV�br̓�f��^����o<�V�A�C�a.��
�|����V�ХĊ�BX"�iT�=Nɢ�h8�q�׳��ͥWä��6Mp��wE^5(��,���b����(%N�K���C��r��ac���ћ��q��f�ֶ*��3Mȶ�{�.�"�2��l���,	��o)�*��e�h�"������S�`�ȷASh��.]!ʄUyy�n�N��OYjEFo�����B��v����P���vMP�tf�ц�W�e�(Cq�ض�=%�OF����9saM�ư`��7&�l�kM�֘�O�Pֆkaw��Ҽ�u�ٶ@uF��/��In��B1�����PGm��m&I>�5�k[�e�7��Z7R�F� i����0ؽ�rUl��X��7�ٔ�Yv ����R�8�l+������X`��̭��C �YYw6��Ww��D��jS�`!i`Z��k!]���[�0��|FB�ɐR�@uV.�-(5�W/D��y	�j�ƣ��j�Ti\�������Ǝ��h�3;'p�1mvp��Eg2���0�����9����rV�Ո<Q�l�v�Bk@f�{$�
���uZ���ʹU��0g��ː����f*�U���f ���t��f�uL�؋YQ����8���B�Æ0�Y
ð�ZN��RX&�Km��u浖I-����];��.
��Eby�i�4�X��B��,e㷊u��2d��c��bK*%(��&�f��\�o�����k�"���6�&����Ӛ���y�h�eP�J�=��g�o�������3/kUK�4�r�Jq,���5
�35ʆ�b�w��a�q�y.�;3�"Հ�����}�{��o����T8�G�����0��˃�0�+Tn�0+RWEH���e`t8�qؙL܇^F��0H���u1٬��'>��\�4�^� ¨N�r+����Z�'�X5�7Oo�˃ #PlQ�#w%d_`(��/!y���š�l3|ǯ�%��ٍ��66���J�Q��sSq0Hۏ*��I�����A�Ӕ]���E��BM�*��
���"�Vȟ­Ez���"�l��i�hS�Z�YZr�&��/Q�������c����ҭ;+^�ʟc��<�JzI�[�&U�%j���5�aUX��41�3[Uf���^AXַ}�Ю��b��L롌I�ش�)����ܦk�5,z�c�6Jh��nͧ���}U��}ZƱ�@���<�EK�&�}���a���G�m)�we1�}Sm8Q,EQ���yz�|�8jngŶl�gc٪�ͣA�5R���ӗu"�JX��O~�V��`����Ӷ��z��2�ʉڽ�+�Kɕj��5�&m^��X�h�2C��+nS{��%�%Fn��,�$�fV`��@���E:��yiMQ��n��M�Zu��F��@��Q1J̶��Z�3W����	3+Q���۬O)��ZԲ�J�����$,D0�.h�fMa*g6��3D.���q���7�gZܴ۬�ƪpȤݹj�o����v��حڍ�����a�7.'z�E�`��G��B�_]�9u��˦�1z��7JI"����43 � hH��7��fEeY����3��;�J�X0a�F:@����˫��i|��tc ]4i�v�F3v&M���d;j˭��jf�ʍ]���(�6Uf��cZ���"�*��ΌRx�i��ڽqV^V�^��2��j�nH@R��1@�h��a��-����6��S�]>zD�$^�!E\xZ�r ���I��F�L���"1ӻD=I�����ڼfي��"鍭��2H+t9)��!�ܻL��߲5j��۔�b��*��4I{HJ��[�()�R�:��Lx�n�j�+j�4f�	��^l�V�G/L��a���WR��y���ovR�����%��d��*�\�r�n�m��n�]�$������.���~�	�¬�,$��{���T��*z�S�abZ[*\"G]��Xp�v�n�d����LvÙ&<�u�Y?X��v�;�ŧ0kPX-gB{�q�����a`������5d�*H:5���6sEj�E�8S��byЅk1n��+�ޛ���f�~�:�fW��R��m�14���C	�0Һ#��j,<�Ж��/ ��t�$,��d�ķZ�Gpd���#��!Ae��l���k�m9�a�$2�ch&(w(�909L�V�T�fEe̳(�#����P�ѹj�͂jڰ)[���OEl�&> �O�	n� ���vp��Wq��rs��䃶�vp5!eB���{�]� X�"����+*�K���	�h��j̨�溫���&1����P��R#u�1,Y��W�̡J
\�g�!����4������̠2�0�f�nd�A�
gyZ���{Kvkl!M�����Qg�Q��r�ԃa��S�C.�u��X��i�t�2Zռ�����Z"ks.� �fS��^hV溒�)z VMhE$��D�&��b�1S]�/���-Jb�d7���̀��WV޸��u�ě�QML��|wd>R��?,cr�S/nd�t�(K��n� *��CZswjة��-��N^�3m҅��d���)u�b���������Xf�d�v�i��v�ۗ �gU�����������S�lz�JR���̇E��	��Ge�ّ�O@ų-_\Y�e�I��`�B��������7.�T4h�ڢ�x~6P������ZB�-��1�dd���E%�VL�u��b�d�)ӽX�Ł�NјP��$���%�pӰS�����X�7|%��r�a"�T2�I�LzMjڼD2��K�����ݸf��q;t�ۡnl{��t�D�uja�WG4��Ւ�Ξċ� @sմF���i�2��mmӡmV�C�jP�J�eJ22��׿m�oX�!&5�i�ӗ���y�H8�RxޫӅj���k�h�Z�)��]���Xv4�Nlh�VF.�Z]���:#VAJ�=�)0�<�\
��%Y��v�2èo.j��t�i�V!�����߷d�7��+e�5�P�D95��ۦA� �6^�ֈ̷��L�Z
�N���Re�рˤI��h�Bٔ���o����
p��yX���P�5��ZxUAf]��#�B�Or�Ơ���`;�`i�2����Soh�O6��3U��妜�p���29�ֲi�@l͕�M��f�ް��h90:�����wEw�S�DQ�V��AEl�M�<���㐼�w�Q��8r�0'��dI���yg$�.���X�6�7X�̱����fVt��L���ՆPI��7`���� �.ʟ"�D�F\se! n��������+��KrHU�5�,��xUiI�����>IZK7�S2���N�(�йQ�0Y�2�9%̬��̸���4�J���"4Rx$���7d�כ��w�v3^`i%�����&m �Y�i;h+$:�p�i�
������\R��+*k�e�p������l��
��l��5��Q���	-[w��&�m)_�7!�h
o ��������6C��R<�T�f5-�ЫԲ�B�L�#��k(�P=�����N�9Z�k�I�y�0�x��¦��FZǊ���*���K��L9֪э�kr;[qe��½�I[`�M<;F�V�K]ih#��y�
h6,p2�6�Ї�m.� @�d̫�����-۰��em�aii���xu���^��eP���|�h٫1�`GYw�Z{M�T
i��ժ���Z��6L�F2�e˻���4��2D*$T����Q�)�i��bO@�>�J�w2At�u��2�VZEX*������;7�"G3jݹ<���cxY�E(ZEÑW����V�֬�a��:�d����=r[]�_.�q;��"��6�2�t"qb8�����՜pRP�76n��/K�e����ޖ��F�����b�H����·K�e*��RJ4�(�'HE[guň�Q�T�ɛJ���d^�ч4V�ͱ��{J�Mq�ݒ�~�*'&Oi��^�[��wI�L;e�{@	X�-� *�@�͔��I������m���h�K`
3fԧ������N�
�X���t��Q;a���ހyv���تZ���{��L�5�E2A����ֶP���Dkjn����WrQܸ2��$:��e�h�VdU˶0�*�
��Q\mr'gq�E̕V�x�]�u��j���%��ŷ�%M�P�Q��j{j�&�Ц�:�`��Kj�0/wM�$k.�y"�z(�2�f�e؞9Ax騞�j�nm���l�*���&�Q[�\j��"���'���۫Y6�*mХSkK	h!��#F7[��Z�6�\fS�C�F�=TL��f(�j���6��l\1J��
��7^��M5���b��m���qh�rJjr̿��!R��ʥ�����k2��@SF!"-�ԙ���n�����;fˎ�X��a~f����M����4w^�vp�e�%=�L�`�mi�m�"d����Zp�(ZՓh���v����\;�3�� ��f�RǢ���)��J^���}.%�)2���n�j�ϯpIN�Lh@F������KkY��m幈ȣ`�m�.��I�ͻ�G5kn��6����3Z�{��dVQ���(BN=4@�S���b��0�Tm~����R���.MCXw'�A�wb�S�N
x�B��:P�������;�%a���*G�ۯ'MSzW���)�7-K��`U�H�\9,�}k�[�Y���\�� ]r�)9�j�U_t�dS��z��ycho�n�x`�gcĄE�n%���]nl��ϒ������Ve�z������7O~���Sl�u����HmAˡ��{�ad�֙��%<�uOm�_|������|�C��K�iк��Q�]�QƩ�W0M�	J�-v՗-
oB��rW][jZ����ԑ��f�}RNXC��J۾��� �p�{,��+�Hxb��p�N
����آ��\�]m��N���e�2����,���X��{��bkW-U��;0K��n��u0ϹB���M��k���l�1T���t��;��e�����1���NG�F'l� 4x�3U�ܞͮ���jƙ��RC3�<G'�ϩ��^�\\֐l�2)�[4#�u�F�_Jy��i�y��JH�� �:KCs�v�'k����d�A����N��	hL���wUw�HsS��_tH��hnjJ�
wF|�d<�㚆$]Xt�W�1�㦃&�t{��2���ސ�#�Z�]}�<���2_a���,�,�wf�R�'y�tEX���{zn�DW��A�;��ݻi�`�5�bW��0��T�-�	��x�������@Cy�9{�i>��+�%��2�8��]Y�����TP�8�YG�)�}����:ž�0���b��kp9�gwby�{�6�R�o���"���d�rs�{җJ}��ⴖ�=�ɓ_	�a�����.��|/����f��N=�J����p�.pZ1EY]��`U��)Û�F�I�����a�Zo�iq������)����9��X'+F54V��Ӱ���;��7�t�{z+�<�1;wnz۹�$���զ�If���Ž������Q�AA�G��l��#s���6�6s�c6�n�2m������f{e�;���y�LF��g,�c���=̌��u�Wt޾9�s$�Շ� ���!gv[�ضѐ�|�,�W�@�O0�Û���f}h<�(8<�l���;�9X�3E���W�]���o{��H2|������;n�,��Hm�b:�s�%V�[xg*B���7X��0q#�u��)�.o�v�!\gYWnn86��減�7�7q�2i�I�WF��Z.�NAXw6�m(�%�K>7�$hʘ�b�7~�a(�LR6���|~�6_m�F��n,UvmP�-�ѣ�����U������U���WЅ�0�L�@^��]YZ.�1X���:AW��	����{�!+��e�;�]9�aN�ս�Ccu�G'j��iK�QRs�δ��Dl����juJ���n�%�O�E���;ً}g��n���q�j�\(���ʖv5���ve�Km�Ft��M\P.�1n#dc3H��CЎ|�m8sy�҅R�q�./-�9��5F���^tgs��As����oU\�|q�-ۙ��e�}z�#�&9u�T*[�)ԓ�e����q�4�&����2��Ԇ>�0��Y�F�2iS}+"绱J��Q0j���8!�j���]z��h�c��}��%Mt��#i�r=֪_BS�4TG�.���m��Jb�o8��ݲ�N��]]u����N��e�!��p�/;��\��R�8��%�Vp��nr���@L��ܟx��V�/p��c�n�MS�>�)��"���ڵBi�*뻙�~�2-���Bk�{F��t�}J6���Z��2�
g�����[�%MΩ�R>}���=o-��{���U���b�5Ķh��w������H裲]q�u�+R�}u�V�Oj&����3@�[�.����hU�H�9�i���RL�F�)�C�1J(�h���F1�bXA��a�)0�nG� p���݋��ms���d��]kzyW*nP0b#����ؐ$gx�nEE�(yo{fi-q�k�pM���F��x�*[V��'T����>6gg|/��\M�� 6�M:�V:�������X��*�p���L4ޔ���P���<�u��̒}�3Nh"G!��n.��\�����ɯ_����Ʊ��K��[�X�2⮆�ɴB�c�*7ָU�7XM�^v�޻��*W����[�+����u�<
h������L�0v���̄*�za�^�~�ۇ��,�G�`�����\�]9���j�ic�Ćs`uz^oVm��t٬ciC ��T<�s!���)c�x����ʟ8��"��SCq��]ѕa�0���:��X�gi�B]��란j�������8@����Eofiһ���|J��>����R�z��ID�Xxf޼�X������Š&Y�t�Ί�:�W]�t���7md��jS�w��Wh�Ȥ
��v�,� Ǧ�-Mh �!w��׊���E�(�R�R
5�ҫ�V��ɜ.Q��>����o�CV����̾2i5�U�8L;q;�銝��4�}�m���(�;4u�3¾R��׻��Ê｜���-T�6������hU�y��n����f�s��[�nwx�$�����Tm��{�-�	�\�e���_$C]��"\��i�؍�N���UDƚ)p9�Iw���Vrp��72�*�@�w�-��-ֳ2�r]P֯�f&��.t��}�,��.���z�m����?'Q�a^�P��\��d�YM)q��ig1�k���rE���Z�R7KP�����u��攅3vM$����;c_9�����9cdWKSXVIc�{�N�zx5Q�7o��6�G���*t�wP�jY�St �M��͊ɳY��Џ-�`2d��VgS���%�����Ijl���SE�ٰ�fsXU�{7����k�����+��t�`�n��X���R<k��P�z��m� ut�#���8��dW��ͺ�P �yaj'����ݱV)�+��n��fARކ]m@�9:��+��7�-w�.�$
�JH�qȫ&��N�jM�S��Ηj�m3�n��jҮ��{��i��Y��������ڨj�=*R��p�׋TG3'��F�gwԥ#�5��
mn7DX�-=���.T�ޗ���=��9��ñ;��x<D�-�����[��x�����C%~��rn ��q�i-	-"2�Q�R������!޽b��W+�l����ͪ�ǘ�k�����f�fq٣��&�c�Z�V�����S N�֚�,�y��b�"��\�����ћ��(e^`${]��{���r��̫��H*t��C}���F"����T7r�+48gB��U�a,{��;D=N��d{a �W���O�U��g\��rv�����M6�*eԐ���Z��w(�i�:��7Զi�4�y-�ڜXw�wW{ʱ�QA8�����k4e9�g3H�:m�+q�*Y��x�f/�ɽ���ջa�Χ���y]����f�J:���U����O6�N��_��F�a��VJ��["�K�VgNï�m��0���GG&�@^��=$l�]�ݯ%L1�+�r!�U�K�47��V:_O���d/q!nE��'�0^��\܇�����Gw0�(�h�ubww'<�!O<���0�wӲ�=�t�S䏨��r.���Ε�5�K�d��f�:�\�&�L\A�0�Ƞ�;�P�I,�9hxj�zq�I!V֘����b�B�J������y��i�(6�d��t��]w}�`H�{|��w�]���˧D�����7W-���Biϒ����[R��m�uo;�v�h�x���F�w7����Ր�4x��b��\{���}j�!2��%��W^C�]ō��Ϯ,��P���7G�+�� ���{���gn����ȋ6G�s�+)I�֯{������9�0t�>�.[RHe#�˥Ƕڱ��`�]��՗{K+�m� �k5��KU��t����J��o��pq����_1�*P�t���UD��uKMERk3p
v�1�TZӵ%��I9�oz��NLS4�f��J�5���]v�\{{V�n��m�be�P�	o�Jj<FZ[.���y�˥pTԏ�k�����������⨷�r�D��O��=���<�Q���ٍ����̏���f���o�^�ϖHWM��3݃ZHa|�Y�C�e��2�4>ǳ8A�Tv����÷�	g��\ޗЌ��;�벋��K���HB�\��[%G���Q��[�M񪮝�Ҭ���8�1S���sy��4#5�vM��7�5\��LY��`Zӻ!`�
��4+�JqU�O�t9�݌w���<qr�=;y�����8�$��-p�6o���5�VJ͘�)T�zxM���ɽ�]\6h7�W�m�.�B�2���Z�6Ģ��T���S��n�32���5���i��1�)bk��e\�@�����9x�J��ap����l�M��g����rQ�'.<6�1�E�7�O�J�H���}�ފ)���7�|�o� �j���|��F�1��YY�v��������4���%gp�a��K=fͨ92yۏ�a�®ݼ���^i��f{bX��Ƴ젙\�.�V�M�{��i���7M��Fl��ǹf|�掠��>D`١��s�����A��3�g�v0�A�&�,!�{0�?Z)�W�ۛ�&��k�To�س�C�Nb�uw��|�g�"'8����g��%�|�iN��Z����.�\�"�ޅm�8y�F����Wۃ2��j]���-%���|��ʷ*A(Ps�,y*��ocma�/�l;2C<?v&��[�D3��[�j�WtRm�	YX��W�7.��L�U��F��-+y:�+5��©\�����ѕ�Z^V�O�#3�6z�4,p׌2��zL�1p㕳��Խ5g{y�nA��L�����.h��3I���t}{�,�]N��K����h�7����,���3�S"7�w�����#�=*���-ȍ~�w�hŠ��6�����X6Kj�����aR���<�{���.�4�oL�~�@ys��ؐ��ph��E+�������͡ufR�EQ|v�@.�;��\��Wb�&ּ��T�
��+GeN�n�:���4wˎ���==z�l���L?;�z>	:8�N�p���W|�^c�h�d�֦P��`�:^�o��Ɏ�ᒓ�^���**��x#6zx���e�2��Ker7�_���9W�@��1���L0�G��,�gonu�L�	󑲕��̅R���ʺTU����xn;h][� ��<�r6ͦ�=�Ca���q�Y�n$������{.��!YB�A�w]�m
��V�_\^�"홢Fї�v^!u�ԑū`"(C�qe���D��]�[g+�.�\�b]�ub{{G��6�gf^�LF�s��[Ӷw3t3.�,Q����6�«��7�x᳓�^�f,�ޣ}�n�ω���q<�$��C(��*�eu/l���x�Wy�/N��:�n�ɷ;�f[�\N9m�Ko!1����;=���O��Y���.?N߬a�_^�4���6�L����=��U����F���I�-�9��1�H��{���" ��Ӹʘ]�9V����M�1�{��̨�ל�Ǉ�e'�L7�wT�L��7L�Y�����8�����'H�(�9��ܖ��$ȥ�E��M�����:2��IK8�X�{o$k
b�1��Nj��<tm&r��4���lY��L:Ӫ=�-W�iˏ6�8���>�K{���o����ɋ3K�$am�)�5��&�j��R+�)�FKάt��U�4���vm��JJ
s�-�}�0h�,P�钩�k�y�'����˘ܑ��S��^��r�h���X��/�wF�}�w�[ݬ:�RҮnP��t�ڂ��e9�ɲ]�&�2Y6#o��*	����K��c��f;�(�쇪6�����t�J\F��獖�\��H��E���/.Aym�� ���ٙ��j����`�-� �6̐0T{Q�jv�޶�&Y���K��6������^���^������w~P�JL%$Mp�FXږ��oH5�8��L[X�T�twj�]��q�=�uG�1� aC�Įw�s�q��F�K8���v�sx���l�4.�f�g8���X�n��p7���.(czt�1QK���s��:�[��h��[�0�A[�U��!�Y�����=+Ƴ���a�� �2Ñ�ٽI�E�8,6��ec�b��y�M���/\����E��{���Ӷ�J���c컌ή�l]�c�	f_8��30�྆��T��A��@���M¾U�2�NN�����X��gxuk=����K�N����3��\�6������P����hs�_b�+:R��2���e�f������&��J�����Vm��Z��.��8I]]�"@}�Dײ��jG�}
Y2�'��v�^�-K�fbނ�%%h����E�'�c��T�;������>��g5j�\2��5��a�z����D��Z.���K7��Pb�����7R��)L}��ejk�U��_[MLn��9��D�
����&�*��B�m�}tjR�Ʉ��{�is�p̕��Vj���긻��{�v�������pS:�l�}�W�NVV��ڦ7��5rf*2��un��MҾ�y6ƶ��T�jU3Z���"�1�%ũ��Va�Xp_7�}��9t�?ws�}	&�#;�plN�`�7�j�>A���7Ü�Ľͼ%��rw\R��锇t���M��$��.�~�8}��u�.����B		���$�}��K�xq�[AA��";�4ʶ*���D���CWM@>wyk\��W�7u>�﻾\l���Ͱ�W
y6v�x|U��z���ȋQf֜���c�[+����B��|��P�	ָ����C%��w��|2�T�/��/��c�ę+W�,C�d���N�c̰ �ͮ�c�����姦����N�/��֩��ȗe>O��0s<8�^�w�9���4�>�l~�ܥ���{N�\[�$��-�2�f��Mz&��7M�\�t����ȇ܏d"�֞�p-�%�>�R���R������	9����}��uy�2''�h�7c�0g]5�����ݤ�����^7#9,l�u����r�n.ã���ec�fd��LoR��P��n�Z��k{W7qкV�N�-��&�{9ە�Z���ڕ��mPص�ba`t�V���1ҹ�O��D��C�u����I�dڵU���9S:��c�/��j
'@z���o iqE:��k� (m�_jt���m,\�uY���1����P����6ܬ�{Q�&�+H�뎺�-�vZ�5nӝ�ibJ]�q��,�W�h��(��I{r���bm_ӟps�eGu�Cy��b�
�͚f�繂�oa�թ{F�����kg�æǷB0�n�k��u:b�UצZIAz֣��'V�7X2�s�7;8��N1lr���1mY��6C˧Y�Ò��5b���\!*�'�Za�7
����^���lj�y��6��e�vԣ�r'S�����7s���0����S�y� ��G Ǧ=��n��2W����`u�'Z���Ǘ�EVw+W4��Y.
ل����&A������:�S��R�1s+�p�@�il��0Vn��FB�G��B�+!Z�&b�_u�@M� a^�E:�͊�X�r��p��ˋ�k���v�-_wi��q�Z��zZ�7�A\m�ɩ�Z�FǓv��˙��73m �;�H���A��<F h<P}�V.=�����P1\gVH����Z2���]����q�C���sWjwK�ɽ�P��ZC�S|��]����ӮMt�B6��/_pT�����f7���m�@��-���b�tE1%u��h��'�Ҹ�.�S6���x��A�ڸz���tS��=�*t�5��')�	fh9�\B�'Ұ���j|�E�Ww��4�x���W�}���/6#��yJ�P�	�1�!ŉ}Z�u,�gQT���v}�Bwbh�'�g,��ŔA®���%j�!��*M/��>رjU��):g�[N
�Ɋ��伇�D[α]�O`���Dߎ��]�8z�s��d��Ѩ[��Ɖ�m�����o2�NෝZ���}���cV�C\�N����/j��ᦓE(�f[�x�L 8��d��;��c���Ef������;4�{G��g�J����0*{�.�d��\����[��U��P5����-�9���G��v�ᛷ#�S^����js&*���ƨa1ʔyЮ3�8�np�#kg'LR����%��n*�@�q��m��D�Ko�*MEϖ�+��Wۛn�w�B����C�-8�0���zQ�<��a=�M�ܫ�D�<��x�7����3ݍU���eY7���c[�Ahv=`C�ymb�a��Kmh��2^.�*R�%�E��c�=�>���]�+N)w,�M��ie`����A�n�1HC5,m���1o	k���˽n=�7(�H�e��E�En��x����J�mj�ŌP�'ou�{�8X��)wNeg�ނ�Ѹi�]��@��ش|c�Bf�G���3����bf�����i�ÂWQ��!���&�OS�I)�K�Zo�����Z�F��r�	br���V�@b��jTL.b�P���_�Y���wa>X.wg��C�xA`����j����pߋ����-8h�8�����y�
.,��:��������K!v~�t����u�ч��u�ot��DP
�9K(�)Bz�'v�U�ǒ��O#א�����E�^Ӯ���K���!�Dبmš���I��$����T���B��ɔ
���	W�볶Ѩ�2�8m�oT�
W`���k�lO��U��U-�s#2v7�7I
+�-�7�Y�1�w���ejc��I��H��r�V�i#c�Q�0R�+q����!�J�ِp��8�[]/:f�mk,̦��S�J����;o�7��Sܒ�']��6��R8�[ͺ��*��+4V��γ�Ga�6Q��m�]�6���ZO��۶���AG5�y�ʽN򘓰a���\Ŵ��F���׹7��[]��i�q�RU�H*}.��z����3p6����M-�i�̧F �.��y��*����d�R+A|�^��V $��9������G���(ݧ�H+768*�Y�"�cm�f[�T]u�Y�)�G7{K��C����'�N�`U��ۘ��ڻ���pj��I3	yV�ɨ:���q�x��)�7�2�����f��K���(�A�PW?o)�Aӫ>�q��L/��FL뛅țf;���B[�W�X�q��}@`zB!�K���{M�5�I�V��=6$
��+�vD�����X�0#CIҋeY9��c����1���J�p������غ�p}�V�x�
|���H�֎�Lٶi�$ё�Sg�8�q��]ڬ����	�gJ'u��n�����'�єnc�Y�g�+�U`��sY��V�& �&��^�S��3I���z�2f#|�=��֒�>��'Q��3�h�y�\RH�yt��c��`�x����u�a����F�>�%�KE������?��OW���eg`�`E�sP���#�Jq"�8.LƮ^�/�66��l��T�t���v�Щ}Z���Q=�L�4^�7�N�q+@�V{��6)36�@�q�m�~�e3�w�g:<Ioaѓ�yկU�X�<��1�RnJ��ad���+U�vy���޸�,�	�/�@B �t+u4bShU�{�*3�o�y?+B924�1��� �����n���i��E��Uw��v�f�;X�-ӻv������)DΙ�C�
[���k-��m�FR�r�o�F���f�d���`0T��=R^�o�W:>�1<h���喛o��n�����,Q�鿎���Dv��C�R��Fwb:\#9\�+E��hK-�x�����i?\;H��:��X�w/��}��R����]��Y1��7�����Y��V={�_g�|�'�:vU��H�BS�=
���i��@���aՃ�h�������rhN���o>ɡ�2)�̑��luک\Eh`2V�t%�\3M���}��'ƅ GS��1��Mވ<R��S�ܲ�:hfo�5�Mf���T���&�{��(^i]sr��u���p@%��r�dɨpɹoH�89Z8t��Y�g;s��Ӟ�4+���x`�#����p����"y.���gt��`�u�M���p��l�la�٭<"j�uݡh�5���v���s��SN�,����R���9f��ܷ7��\���P1���y
Y]�l�%���/s�q�áqy<��3���vBl�mn��&d���̞��I\Y�&1h�
�l}��$�o�q�0RQ��jc}y�o�:u)���{�qr���Mt6�.9v�>	����3uر�Ҏ��m��&���p�bu���]U�7����܃ךY[1M����]���@��#V�^�}[�:gTnV�t���&J�܎�D���N_bvPu6��Ա)��W"8�z���/+�T-��%��b�ki_�x��٤���֖�%2����]vghO_Ŝ��홎��Ym�M*�E�[��Iβ/#1ح�`�*�d}�hc~��%��9��U��b�mp&���x�\�h��%��dǛ�'��}CKX;7�!gL�᫵,pfڢ2���Yre6�iC����݋c�v����r�݀\�ػ{tX���&-�l��<�m+�3�)XQ	#�5&�f��D֮���~�ɛ�a�=���N��Pΰ�S�H�5]m[����J5��2uA�8[��wj�ݝOX��}�=�;j��<�a���]^�����mٓ����E���'{h�#�Ҳ/8� o�M�B[�aTXD��
&t'�yK2���/:����)]��V>^������*�4 B��ڎ��v��}r�q53�>ܷ0J��B7�G �O�Ɠ�5�o3�:{�Ǯ1�R�].��A&�
�Z\v��T�u��7q*W/� �9[8�ꡰef��i�c�Feyw�:
��1X�Bt5.��q7����6���R}tK�d�W��GP���Ӧ���H����,�HNhjA�g�T�c����i<�R�gr�c첄���@��ӳ�����`��#^WϦ`�|�.�yW����m��5�[���]=]��R9�cv@@��[6],@�|�56��RP4F�l�����y�L5�6��L��TEv���I��Wj�kGШ}�������
�5Ĳҵ�͖G?�8R3I��e�8	V��C'���4+l�ftneμь�l�j�:�
��=�}�qTw�R+�.|.��8�(��3h�]5G���X����=���5�Nh'fSf��Vb�f�e4�u��ʲ`u��������H��#�����T���ق4fh,�N�$];��g*ȅ�x�ξ'��z1y��V�E=�˧r��-�}���c�;�:tt�v1eO|�o ���EĆ!�;���dti+owy(n���]53���˴.�h.��Vo�6QR����@�{D��m�|���{��%;��q�d�cy�!�;v#�'���ǝ�G�L�����;k�z�Ý���CX��o��Ly^E��������r����aPc}yo���EXa=nf�=��O��u�Y�FSD_P��!2�J�u���׹���{#�5-�N������/$�j�p�Z�Aɚȥ*aY�1c�f:�{�
�u| �����gN�@iP�SǙN�"��m��GgPbĽJ�Ǿs����3�]Ry���c<��^�s�Bq�Q��<��E�n���^�u>��E��k뤪+��v�j��!1�H���P��|0���5+2����v}JO���4�h�η���wz}�XQ���9�4�샕&vWkt�Hh�z�gV��dqu���)t[ėCb:�D�(F����y�dԩ���򙘫$�r@�RgtG��>���MQ�X�[�1.�}�^�:�Ҥ��o̬�"U�JT�n�a����䴆f���,ܮJ�08su-l��a��{�̰M�a&�SD�p����:�6�b��%�C��)�ʗ�٦���5�NV�:��4+i���w׮'sgb�R�J�oZ�͍�]>�uZ���b�7��y������צ�-�.��|�hp�����n��WYH��W.;F�~u9��s�ᙤ<�i�O�����x��z"�g��ыo��/�n\bE{<8a0��Їm"nf�qV�.�{ܒ�=���C}��8��FV��~���.�ߴ����樇래w3������|y.[�U�9z*T���y�
P���gӿ@��\�h�􌥪R��4���-ң�[��X���a+E��E�a�g��pf�!�o�qm�eu��/h�Ԗ�B�t��8���B6RL��`����o���ѻr�EK11��;%UY� ���n�w24(���;�JX�]7�z�A=.���cW������kr����:ы�_���/�U�=jS8�n�+���@=�e��E�����@,��vn�GY�X8�Jh��:���=|2�<˙���v��۸]�TZ�1A:=��RG�lm���K3PZ�#��� ����=y���Z^r�^:�7nRۆq\�vӸ5LA�l��(m+�[��<'gTE�B�J�)���6��L�C�eTu��P���gqW�dw;���)Р�uѐ&�hP����;mM�.�Q3*��L�:��3
��v�ӭƶ�v�'R��'����Y��Ro�L|��᝕"�4O�]
`�{���bneBX�G��_eZ�<~GK��+����렠ʘo�}?�+ m��ȹ�\2�q��*������|V)�)Օ����-Ev�_x��e�3.�S��O�𕏰���Wr�cq�C2�Jd�i�A��UCn���}��w3��8r�a��Nפ��	���e|���6�x�k�d[Rm��ѩ;wZ�Y��1�&�@�&ݾ��vt����ެUb2[��x�.�Y%;J�K�T5����X+���g,l��ѮZj氳Nc�����k���˽]�0x�"_fy�̕�xk���z/��aV$�e��9��+�jaS�U%������s9���t�&���stޚz
<R��]�gD=�4����AX�G����W��LFl:�$u�
3�� ���դ�������>>����W��FqWG�Y�$ި �v�Ә\>��I�p�-�I��3��J���o)Q�U�vަ�«�;�q�f��s���ǋ�ҷ�r�sg8�C c���Yu3�L��3n�d��*ˎ _�x[�T��pq8%��.{ײաoB�k�f�3.ga���'�&��[���Gp捭�ֶn���(]kW;�w��^��I͛�Ğ��}eʜ��I;c�w*��7
�v����aə���I�2rU����0��D+����8���������vᰑ�*&7tM��ͻ�vӆ����W)޺~������G ԅf���)yX�i�eZ�S�ЌkQH�le�(�b
]�	/u��7��B��㪵J�9N�n�*��A�.3i�V{7e�To?z}���=CA������,p�jn�]*N=��P�ʯ{F��"&㴈�f9L߸۞���Q�HU������hv���ͅncX!m���萈�UGsܾq>���ñt����:���aeђ-�Ӯ��s;�V.�o��c�Y}ʃ���$MjlwJ�3i��ӂ�#�Ư+-�����i���aN6F�nf�a�7���fR]#ҋ���#�|�φ��R�����JO
�oK��}��W<��0+�i���yS��*����j��$����d*�-Wq����v���{7��ʐw��ћ������֧����,�ݹ0_40@V����nu�*cN�r�ޔ������Uk�M��fLPr�گ{�3��N�Y��0����A�j�+��j5�!b�Q.�v��.�fr��	s����K��q����v���]*��]�@Z�pS��0ޫ(�S������-��x�#ڸ�����:g����˴�`��f"��aA�8�>Q����)�{���ս{�"�;6�)�0N>���L�X���{�Ƽu*��gLy�n�7�o��6�v$�S�:޼���`'a�F�+��ZO�M�W7&*�N<�X�J<�ֶQ�|�<�Ǩr�>��U��c_��o?}o�~��+R�R)Y*֪ƴiJ�$R�X�*
�V"�j�P��(���Em(�(,UD�"�aX��"���-����J��`(F+E�� ���`�UV1Q�aP*,A���"B(�mH���b ��U��R�TH�V)Y*AAV��Z�*5��E-�Q��E*TX���#DAb�iY�A��X���H�(�E
�e��X��0D� ��QJ�(��TH��Y6b�)��EPQAEU"�Ŋ,Dd�QUYD�Pm��V,E�(�bDTTPU�AQb�"�*�ŋU�EQ�1�UA�l�E��`�$DUc`� ����Q�dF"(�(�cEDX��J"�Z�c#���`1U,DchXĕ�a`��q�R�pJP8����׎�s�MSM�+#,��H��#0l�`��Knc�<nE��m���ژm�����\R�}#��>�ǜE}݃���;����e󬸱�ǶP�QH�=t�V�۫Q�þ�	�Z�����EN$=!M��D-�׷��9T'�t���
�uv��}N�ؗ{B��)�M�T�	Lˍ���w�cE]���G��B��Rq�U�ޞ�����HKQ�w�v��:U�'��Բ��Ө��j]�b�l�,���,+��/�h�{�]�3�r����� ]����o�U�xj�r�*:�ۼH�u���w*)tv��i�'����pe0c��{�Ϋ���VS��Ot��R�����b�
��_�zZ5S����!�ɺ�3��[&I�1�����%�RW�������
�sܷ\�Y�뱻,}�ɽ��g.5�Nvf�˄0^4+٩�Ou�<��\��4����_c�!�h�xt�G;t�96�r:���ǯc��^v��u�ܩ{�V�ny�M��7�o�ca4�;;�PEk�W0�O�t԰�}D�?M��Jܖap)��=@�D7��ש��!��uM��XzD�Ư�h�O�������\r;�WgC����~�������!�Mx�����k����r��{�8zw(���.�L��>��zi�L�bF}z�z]w`��Z�X���N>�b;sl��`&�jY\Q�P�`�Du��%q�.e�Җ��wdj�������\^�����au,�W��AmI�f�S�m��	���j�%�aqo7�8{�;�=�6�r�c#���ko"�+RUz_���C*�r���by�qԝMz�Tm��M!�nG]X�=6k��S�Ԓ��'�lu@�+i����Yn�X���G�K��g1E�ηu��nԇ�������il�+*�Z�T�bu�����ݥ��uv�s��o.U/ͱZ/�d.,)3�ܝ.8�,���[:�@�
t1^ѭƥ1�i�$��a�g�y��ą&]���m	W���F	�;u�v7й�V1��p��<��VK����G��&�N]0���H�Eo��uPꊹP3��!�YD�ө*�!��w����+���JI�'��ru��Ş�`ː!�P���<I��-�]V�K�h���u�ڗ�vJN��L�]�m��J{�U6r���s���j3�9{�M���q?�]���{��l���P�V�D�t�6�R�|��u:�D�
��*<4q�h&`)�ttO.�1M�9ͅj�%G1nD-KrS��V��r��Jz��>I�4n浃�bf�x������v"��D��b��!G��[��z��ޭ��Vy\�XA���q��B[+���$K}=��"�u��A����B���i��We�{<�ɬ�8�ŵ�㍗�����+�p�b̭���ά��3Y��%^:��'�,9M)�,;�K���ڷ��ޚ؂���N�ҲfV�8Z&�ABj�y��C�i��K�],��N��V��|���*Y�^�V�bf�Ut�ӛ}�\����5E��W�X��cF����H������(�ee�maѓ���1����Gg��U�j�S԰��>p���Ό���w���7��i��p�˰�*�����(�v���8/\��K֜8�y+�fG8���L����y�tۺ@e ����ohu.��w�W������;�һ�񎼣X ��E��\=@����j=]%ՄЛ.�A}z�8��WN|N�{۞ �9���Y�>-�$��][MX�����C<7��/g�A�e����~�B����Y6��E6�^�����")n]Qh����j���r���mz�K��V�ކ�������<;��8J�Rw����WS7�*�Xϱ�wSu~r���-Wo�v^p����8ib3�J:����(������M�t�9Y=�,���m{��+��?
�U7��{p�:�������W�:��/�}��U�t��8;\�׌T�h��W4�zk_M[+,�Ϥ��C�O�
9�+}�ڨs�Q�
.����;Yii���N*��XX噕z��-�9��`DnP�Y^�m����z��S��S���_(\��0�D����ѧ���{�"�Y�^�=k�AŰ,�M�:&��&����<�,�ʢ�R֏+rׯ�oc�ڰ��P�o8�xfx�q��W�x|�H*�#
â�X�WvӘTD�k�&�i�?�v�m�+{ެr�����WV�����K'�f#}l��=eL�ϡRk4ggn��]��
1Ge�:p{����ێ��:�y�<�nL��sBO�;����ٶ��s�Vu/�M�gF��T#�M�^7�O'�E�&�l�o���J��hMH��X���6}I��bF}i۵�a_"zқ�YѐN����Q~�w�N��=|�������>���9�\yʤ��\�{�8,����YY��i$i�ɾC�e#��̷^���nWO<����h�����G�������{�����[��C�萴�!��A��l�"f;������[�t��Yo�Ժ����h$b�;�󴮅�2��~��gV�t����;vo�T<7ڒ��6���յ�Ļ��Қu�V��[�(t�Ee���}��Y�~|4�o%�Qjk�*���S�>��qB�r=wًN=������Z��!�H^��^2�+3��`�>ק�?lvQ����3ے���N���B`��A�3�ĩ2�����WZ�]:rqe��<Z���9�n<Q	3^�]O�1^���76)����F˜�a�s��d�ح�à�%�uu���E�`܉N�fe��2)�mb��?pv#1���}��ֻm8%b]�Z
�h躻�m�ÞVY͗]J(\�k!:�����A�N��QC����ɉ���F���ɝ���R�{�tF�Y��tҼ�S��pJ��P	=47s^�r���s]lϏ'4b�C��?tOP��и۝��YB�uf�M���)�����f�׹�t�[���J��ٛ�U��+J�z�^�453˜��Ya�Μ&"c���'35���ܗnu0�c(k&-w\؜��!��Ew�i>�����jǥ�-���1���[{�կ.��Y�4�VLtJ)�C4���VY����.�6.��b�k�tz65v�o��S+�*�sc���RJ+���F�,Y^���:������r_��꫐s��AR��r���k�b��њ���KSv�ENu��:����{ʃ����v%���'.B��+V��y)�6U�9T!�(����gh��m{Q�}��q@�c#!C�8p�R�<7a�ۏT��qR�i+ȁ��ͧFuEp]&��vlG���U~U.�c�;[���/_x��cμG<��_U��Sm_(��̋�X��s��2��1:F�ݓ�wc�A͖��ܒIJzwQ.��!��L�׵̚��4�,ж��m���$�u%���-8F���uWV���K���p{�W^��a���ǔ��-�{"۵��{.mj��3�w`oNl@c�D��VƜ�R�����5��6ވk�����mSg55\r->j�X��yS����R`[�q�Ǿ>�����
l��I��$���U<0�s����S8�ˣ�g��M� ��7t���;���<�L�s'gF��7�������V���̽�u)�'������n��(P�}�\�����&�i2wiNJx�Q�i-B30�b#�,M<�r��B�[c�fs��s�&��KY����콴�rM�]��7��f��c>[Gw�W���]+1h�3�:2�T���L��j��z{�����yJMC#)�����i�)wvz��\�p��ƃ� k׶��߱�ڕqx��/��'�d�}�RԨ,5��A�W��9о�޳�5|���F�e"`g�Y�q3,��qRK�b���]:����Y5�����;��Fg\F;��_|��8��/�v	��^éε�O�Ϩz�����#Z�R�":�X|�y��k��ڎ+2j4�#�B�q;�vs��6\���"�SM��Hͥmr�[�'ڷ�qr��5>�uVjkM������\�S���v��)_b��w�ٹ�.s�'�Y��*�f��9�8K��uC��X����R[Bg����«ؑ��ǋ���9��X��]�p�a�%��e]W�)��ќ3tňDNa�n�m=P��I���\�S!j�!�J�6
�j�uM��{�s&%J�]/V,yM�,���SN�*�r�@�*Q!3.�����#��ނ�I��i���OV#���mv2<26[vu���28�̻��Qyy)v��\�%&��q�����b�s��`�s�d��aP)�O�c�݋�6_zK�~�k�>�Bm\�|G�g��[j��-��p{p�ȳ	٘�������Ō�1ڛ:���`�?q����Q�{�_yZa[��yzg5��	�-�AX�b!����=���2?=�\�AP=�R�q��e���'�ɓjK�o]��k{0Psn��hhI��9�h)�l[,b�2fgL�a�qD����j�j�XK0�|�$��1�y�j����J�r��Cc#!C�S�j��KV��~f��Z��Z�ǽ�{��jy%���W3c*z������Z�Q�+�Mnv>�-����ʢ���}ɝ5;���Z{��~�1���š��Ѵ���[b8Ebb��5��)뽱�wi����h���r��(�՚¶nX���6��3��\�Gc�6��ċW�ݳ�,�ިX^˘�o�Z�n/,GN
�٤6jS<��Rv�+�����`~�<ſk��ty����.-�=���B���v�B�5R*�e8�q�-�ӯY�o��8��XtH	����r�
�WOJl����1�o:�^��RX�N���PZ\���U��ܼ<aa	��}��G{v�j�nFic��W	æ�z��	�ߒ4���}R(rq!�
��(�y�g��)hj���k��%�)=�I$�e34��
�Va�B���.vәFb���W./��k:�7Gj���ն6�Je��%K	tXb���N���33�B�fu1_�V�'6[=ܡٗ������P{Y2X��ON�Td��ݜ���yr�@;�j=[X�K��2T:
��rU�a[�*pރϙ����yPY�N�l����X+�*���v%��ڸ������tdˈw#���Cv�b���"���y�7��SW�X�.�����%��Cl�����kDׂx%#py�nL����nU��թ+�������rZ|�3����yM�õ�*)�Ѹ9��X�C���T*5�K�2��}��ý��WI��bx(�u����h`��q	W�&,�[�x�ėt^g�+~��h��c���V��Nѿ�g��n�S��礋ɴ����i/1����X�"��z�	�hW�53v�Ju���?G���)�M��'���}�ez���s~�4��C=x��f�A�8�F3�����H��m�O�x���7�ž���C�ɹ�R"�<��R�a�ٽ}ZĹ����Z�wB ���GR6;et��˫�]{pO�V4u�(A0�k�����n�Kw؆+U��6'ӆ�䛆Ydw��h��M�4�ʜ7��HI�*���Ax�������y�R0���g�9`�݃������G1*�c��s���4��{I��-�<�4�j#t_ohw��͝���(�w\�_@|Pn�o���>-G��W1�4���;=�߭�{-��/w (�[��k	w��K-��7%��{T�e��;+o�a�Kϑ��{x�ыNp�s��2�5��Q+�����T�f�)���E=ǫ� �w�H^j��n�pehh�����EQsH̸h��>ܪ�\����ji����_t�}r/��6�m�����k��:��,S�䢇I=7
���N�I��j�N�x7{.�{X%,�;�K�+�I� ��g��-Z��GO�d�9B���\ݣ;���8釰!]�R�{��A���N6Wଲ�J"�v�}J���NWmK����y����%_z6�u�����ǃ�������__cr9�[ێL�&$J}4��KK|{���3�$�-�Jpϛ��� g�����kx�w]�2w]+�kN����u����E�]�}�D��-u�na��&��Ù�m���V�H�����>S2����/D��r榆�]rL]a�p;�9P��.$;�C]��V�����f�7�f�#�`&��.ڈo1}Ɖ_n�uj��j�-R��Hr�rD攌�4��r��`�m	OUvVJ&�^�������[�FiS���Z2=��$�E�w��k9�Lq���ī�}�C�nD��L�7>�@�p���霖Ɣ��ܸ+Vp׌Y�-�u�+X5�xT�-��+�	 +�ab[+5�b�L4(ӬU ƍ^��A�}��	+�h��i����6�T����)yLmrF�ά�%
U����ٞ��p~�3�p�Y�WM��5�³`�彻8֕mJ�M�V��:��������ɂ��#����Sn>G� &��o."�1%w#U�l�׵���^��	ȳ��wQd�l��#���%�!�`��]�0�$�:�־�O,�4�K�z��Ѩy�7W�����M+��i�<tx�n��y�I� ��DX�A�u+sM�.H���KU�`����=;+q��!c��E#��1?:
�S�_��|y����?�K���x���Hg���;�4���$�=Wr9|�ZZ"*��dp���qa��I&��,�nj��r�F�e[!!l=Q�N�s�Ҽ;��wyJ%�����S��n
�0��4!� (7-�8��V��e��j�ʏp�hi���x�0��f�.j5)>�oSH��*y�)Ѭ���M�3m!E��a�v{�����t�s�n��T��fO�O١
5͛�NL@��b�ec�q���X�~�αp�ZQPYTDU�UE*�A�**�(* �"F"��QdUEd��1-*�EcR
#X��P,��TEb�`�mX��EJ��H�Ub�`��,"����T��X��Ub1EAb��R"0�*�YmDV�EPU�� �Tb�b*�E�DF
����EQ"
,EEUTV1X�AF(�X*��k",X�")T�AT���Q���UR*�UQ�-�X�X��cj"�*F,E-�,�QET*Q��0*�D`�QAQb��ȋX��,F*/�ETX$F�¡U�X��,A��TEb*��mDV*
DT�E"�"*eUUPJь�T(�����R�T�`(����ŊA�b�P�EEJ�UPUA`��,X�"�R�#E]�>(��D(F�>q��m�.]�JTt� ���x�m.���Ũ7��R����Z�;��Wr&�+�̫dѕ7�u�|/���/�%�q!�'h�v�|�Xj�]�뮎�fS��]�ڜqr�*���W�-����}�cm��T�������=]��oqW�\��s1us�eO���.�y�}yXP��g�tHL���W�[|`ԝu�J�D�]��Lf�+�
s��[�o���Ϟ>O�td-U�m��Z�xe��Ǥ65i�@��E��J�"Y�`t��by��´��r0���	s���Ӻ��Qc��!O�2!��~*�<�V�v'�k�[�U3��.�멝�M+�u�jЩ0!͠������YTZ�㊠[zU�M!Kc��8!����&�E�y����I�M.��2�\8���+�
�3U��V�3�xge�@���y:1�r
ē��̣3�"
˻��2��q��\PNc�x!�X��L �|n��D�~�ݙ����n�d�NFi�����<��yr�'ԭeC{�(W�8�	<3�-e�΅�:��A%`[k}����g��ӌ�J��3QCyC{nj��u��M����%���%�9i}�Ǎ��x6F@2��!�On^��Z�Blț������>e�Zw�p�����o��W׺�z��~�h05,��!��#�"U��|.���oo�e6���R�qn��'���BsWP��]/�Q�����-�/���Z�{f�.��^i�I^"���u���XŻui�e����lNM7�+CP�3��c[��֛��g�9ׯ_'z��ɡJ�޲�zj�HO!�E2��~˧z���hƌ�V)���+��jY\[vBL�xfw"Mv�s�oU����[é3�1#x����U�ϸG�iq�\��w�=<�5��VTw����ThC����V;T1*�Z^�v�oj�v5�I+��������n{���|*8�׶v��: j�Ŵ�Y�}��P�r��sA7R�Q>s�!�ox�*��(�A5y�-��[˻X���P��o�c��'C�Rq��E���a�zR�g�.We���Q�X��u�G3�7<�j1���i���p��ǯ�z�׮���|����5�r����Ȩܸ��fR��s׹+�RO]J�F�So�;��� ���&�V/xC��KW�Y̖f%��-�}LR|�:g�Ǭ��{[.G3��_���Jz�7�=j�>\�����D,u�u�
Н�ЩBf�2rg�ۅQ��S��勎~�rD��8�Ł�c�#�-��
i��..���g->d�w.�I��j��Fh�qX�˕ׂ]f;�X^0��x�5������y��a5�0��Ƚ��	w+mV\�cD!�':�MD��Vg[�/��s�A#pgX09�:��z��:j����;uZ.ݴ�����a�9���-.z�}L���O���F�
�P�xY&iNd��Z�Yn��B��5��;A���������ߚ`v��ǣi]�G�Ʊ�o���Ȥ����b�R4�ֹ�u�mnЋ�g�<἖5��wlfߡ�����
���{��u���XN u�����'�O2v�G,���ȩS�#���>��2������־��߿x6���!�|�!��C>�|�~g��ଚg�=�q2m�8��v�I�&{d��O�̝d�:P��>|������~���kN�xw��V�Y�(���s������sk�0(�=<��bN�K�n�*�L뗧{���|}pU�K��W�wCE<�u/l:��,��h��Sp,\,�a�:�`�O7�36��;[m��A�������m��>����'ӎ_N>���
"{H��>���:β��	�C&}���I��c�
��m�ю`�&�m!Ědϱ��" R�y#�G���B�.w���x:���-ϼ(��B>� ��}ofd<���=I<����q3��gSw���!��bVy���N"��^bu'm�d��g}������u��>���vI����O��6N$�����'Rm�g��bd<�o�q�l�ǽ�<��0����f��N�VI�6{�Oȡ.���]��^}���/<<�y�ml��'����4{��C&?bO0�L2~CL���o8�d<����a?�s2|� };�$���2�4�y&�4�>�;ϯ��]��k�q�����Ң�e{���&;� q�vȤ�I2���`d��CI�C�>�'�������'�M́d���M�}�>� �~S�U ����{�}����?}xs��4�(�y�>I���2]Y'�}����`1�u��>���&�4��N�9CL�!�7I�6���}3|�?0��}�s���[�&�v���7�g���3��#�}�"�����>I�Y�� a�C��sd�a���,>$�����0�d�i:���fMo:�}���2Τ��ݿ<��h�Ov.����{�8�u�N����:�/py��X=�@���N{d��8.l'�5y������{a�@�3�&�l:�qu໘����9w�ӿ����}����d�6�4�d�/�I�N����:����y���>����1hg����`籷	'�5�`�2���~;��3�u�>��S�G��ӑږ��8�E�ٰ�	��pM!�&�,��y�I��&�2�Ⱥ9I�L}�CڲL3���M���l�a����@X����	�`������3S�7RguWbW���O{��W�m��IC���aή��0N��TZerWO�t`�+����,Ђ�51�4�s(�`�Rر脝2̰���^&E�N��̫���(77g�=s��f�LG��܎/���޺Wѩ���H��?fG��<ߡ�b���d�l�$����Ğg�����XE�[� �O$�/��'ܰ�l��l<��hLs4��u�>����+iFn���������=�(�G�Ϝ��*�0�
�����i�C4&��&�C�'�7�q'U�g���d�,��'�`z�]��2y�����x~�z��[_]r9�Q�r��������#��������wؓ�!�7���+!Xz�q�L�͐�d��;�d��h�������N�z����A勶��~a^�9<���@}�/�C���o�M!����'����~�d?!��a�׽�?0�O�P�C8�!�4���C���I�]��O�;���T�I�;�u/�������{̏(�Gԟ�:���}�!�Y�w��O$���g��y!�?3L>��
βN&��J��m!���M2m�}�[�̈�7��m/��>g�}�A>�&����d�~d�=Hd>��Ri�|n�u!����q	�N���?2e�_ԓ�a�s�*I8�׿|���\d�����u�����d�P��y'6��u�&f���8ɬ{r�N�F�q��[��P�8�w�!Y'�<I:��c�̘g��{������wyם�_�ޒ��H�	����Qd�,���'Rq�v���u�L��s	���ON���$����|�{�H����tls����gW+�K�W-��{@z���|@��S<�Z�VL�
�$�;����d1�@�M�"��0�l��'X��O��C�CL�����������^R��3[_zH���a���>���[��2~fP>}�y&�2�;�!�L!��E��LϺb�I.�P?0��&��:��M:�Bu!��=��c���i�]�����Ù��:z[
�x@N(��1�u��+k{DAn�4�%�M��;��_BO��u�|�]��]�c��M�q����!�X�>`� tCԊӶ�9�k�q<R.Q�6��u�1���)�xN����ٔ�����y�J�Z���_�����8���ɤ��d�B�'(y$����2mRg���m��^��!P0�{c�$��w���O:�؁�F��yB��Di�wG��f�����ȏK=���!�wY�C�h7`,�)��2M�Y��pE�u��!�M��׻�y&�1l5;���s�sa<�D�W����3��}j��P���`��v�}y�a��L0��i3Ʒ��d2}M0�M!��0�����	Y*c}�CȲL�����!�ШI��߾�}n=�{��g��!�0��{�,&Y=��L���M� ~C�m��6H|��gٓ�u�i�d�<��쟒e���sE'��P�,%C_k�2�)��쫩߷7���i��#� 
��r���b�Y0�>p�y�]�%f��	���!��u��I�5�q'��i�d�ovO�y��l���=��Ţ�>:{k;���}�������b�$�>�2d�i�Cl>L�����P�ɾ�J��6M��!���!���3��O2M����N���r�fL5�zriU9��o�}��ܮ߶����e&�?Zq�����bՄ����x���p~`~a�i�ɶC|�����+w�I�g�4&��&��k����}�~�a?2w�pN"�|�'�O[�O�:��S]�>@�d?{�y����s�?��M��ԇ��M�Y6�T>s�`��3��>�8_���N|�>�bu�� φ�y�S=�C�2ɓ^��O�35����tn��N�3{�? y�޳l�K�|�u�繃�:Ρ>߽�!��A����1_?V�K��u��wރ�>��zc� u�51�i�j¤8�L�����Mwz�'5�I�N�3�Hu�����C��!���8��_~�B�;O�m�����a��S\��Xf5@�"ۧ�}���`bVir_�=���p㾒�D����kG�S�FӄY�<hZ�hĔ�#L(�I�}Q]ا0!(��2�C��涷3)�Cc�Z�!�]Io���'SF�����q��[ʌ�����| Y���·wNj,�xq�����9:���4o^�Y�I��b�'Bb��?2qRV�zǜ�8���9l'Y��y'�X7a�i8���v����{w���}��������<��M�$���~/�~C2{�
�0�C^�"���YԜd��6���d�1�=�@�xQ�y�b������o(�7��?}w�s�P>0=�<�u����`�Hm�;�~|��4��}�<�L�g���y&{�*,���w~��N"�_ q��dݠu�<�5�n�1���nT�[i1�Y�yR��,�y`>�3�~`Vu��f�}�!�y�h7�2~C(���aY���O!�O~�E��M��`Y?[	��o���}�����Q���:Z�NE���}�>����Dx|�I���'X��fНC[�y��X�XO�<���!�y�s��e�h�?g���m�����L0�v����N�>�jJ��7�|��1�{H��!>�Bsba���`i�Q��q��`+���gv��2͏�&Щ��8�����{�e&�Hs������_m�o�2�*��ܝ�k���$zϽ1 }�� T1�๲O$�{�a�u����$���Fl:��&�[�N�3���d�:���
a!��~�a*J��7� l's�__
��<�?
 �{��|4�j)Os�|ɋa�w<��3;�m�I�M^`Re��u�c؁�m��Xy��f��&��'��d�a���8�����WX�����I}�	���Y'�w�'�<�	�}��y��d=��L���� �0�{v���'-*3hN���>I�6a6�����)��h�W:��������{�}}8�&�t�u���)<����d�f��C̟���=�l�ۦ�`,�'wt����=���~By3���ۯ�����R�����9{傳f�BQL�C�I,��8ַz��R�T��%�zł�c�hf����]]��כ���̩�)M׺��|dw�H�uA�T��W�� w��yAV������c�����e𛙩�I�}34����Ph�5�pwV!��  �6��̭�5��e:���d�!�ϵ���u��~�a'�d�i:��Oܰ� y2�̇_�L3�va�~d9�u���t�����q���4�R���+��[�sљF��s�BTM��3��f��6Cl2ɝ{�'k��O"�g��<��(݇��v�Gl'�L�����I���@��aG�7��+*O�k��������$��a��Jɦ|�َ�CL�C,�6Cl2ɝw$��0ױ'Qa8�3�I�O[I?0��yǼ8�B�r�|���=�֫��.��?'�'�����Y�C��̇�l�5�I��5�ଚg��!�4ɴX|b��O�3��RO�35�I�d�t����#��#���Ż��{�v�7'�烬$˴���&q�O���YS�8�̇'}�0�a�5�`�u�~Mc� q�d4c�<ɤ�E���!Ę}��g�� �6rP�;���Q��o|�I�RO�OY:���F���>|�0C��{�q	䝴8���,�>�!8�({�,�	�3��Y?! x�y��G��|75���u#��B&~����{���'X?cO��q=I:��~I����Y�q�� VCɓ����d�4���bO!�L!���!���*�N��t<�ػ��{_z��������~9�_�7�d�#��>��� |ɝw9��CS�'�N�ٰ�O����bβC�~K��a?N��3(�ؓ�i�(��˾�/s�������O�a�?fa�hqO֒_^�m���r�y��M:��I:����)�C�4��3l��'�"é�{�=Bc��|>��r��������L��~�<ɤ�E���a�!�`��O0���R~k	�k@���0���e�_`'Yr�f����M��y��޺^�����f�o�6DW�],un.ԉģ��;*qm}�i'�Ӕ;C��gEL/����m,Zr���][�]����K��[�H�QW`��q*��e}p��I����ڽߴ���Mf�3��y}7aus 6�KOn�]�݆t�=^�?�����޿o>=���߿�2N0����!�y��}}܆�?"��O$�&gsHy;�๲N0׽� |�I=��ĕ�ɒf��3��N��y����?c;���Vo}�A굿'��Gȏ|�A�Oɓ�<�~aS'3�yY'SR��M��׻��2b�笇�0�gs���y�W��&�N��`q��%��f������_g?	 >��=S���d��a��L�O�`)�Qrv�)<�;�C��:���7hMO{٘@�&-N�0+s�ۄ�̟��k�_<�	͏���=F��>Fx">g:���'�l?0�a�w�Bh�!�O3�>7�~d�O"�$�$�c�bՒa�;�`~k!���T�|� N�DA蹳3�U���%��'�A��}��L02s�*g�'_��b���d�α<�6�G�Ğg��7$�'Qd�n��O$�.�P� y7����>�����LH/�'ze�Xپ��T�0�����?$���d�M��Bi���pT6�̟3L�4&�,��y$��Y:���	�N�ɣ�Ȁ���ab1�a��Q7o5xz̛g7Cٰ�0���a���}�`�����i��}�?2C��Y
����a�O��>3d6�Y5�,��M��$�=ﾪs&�5*�8����|��(����Rm�'-<�u��^Y���:�!�'���C���k��l'����3	>Ci�a�2��6��lz����I����}4~�dFw��KW��L$���2v�'�8����j��O2|�O�d:��2c��m��6[!�q��}��?!��'ƻ��̓��w�y�i	hɏ��ۑSv�˾���d��)�>I�w�q:�$�N:ݓ�>z��`u&_'7d8��g��q	�O��`�N3��g]�`��	>��>����NDl��6oT������+n��:*^�O#K";L��=K�2�TZ����7��f�7��L#K1֟gQzr�՘�;�\���p����r`�z�(uY�����7,0�3�q7Ɩ���.d�G*T����=�6zҜ����  +Wȝ������>I6���@�3}��d�,*�4ɟcN2rc����u��q'|�`|�XC�q;������]���|}��a��8+���Ky�Y��o�����,�ഓ�V;�I�2{�O"�<��8���n�:����Bu��c�&�$�O�d�'����A�O���Rt��u�N�$�|Os��?$� |k���i���^�'�0�a��*,��wt�����ǰy�6ԟ� ��2�XN�15�G��@��B񟈤>*�:���ڮ?o=�=$�8����y!�6�3g�|�2LϽ�Hm�@�:�,�E���!�L���Qa<���dݤ�Ʊ�>t���y��z�p�����r�syϱ���!�Ĭ��hݓ�m��>L=d������<��Mw��4��Rg���m��]�y&g�Ĺ�F|,|��tG��3�_)��fݽ�ܯ��s�6�	Ğ͓��0��g�	�CG�i�����̘M��d�B�3��CȲL�;a�M��ϻ�y&�&#�ù�6m|C�&o�[��}����ޘ̈́�'�P4�$��w08�	�&�a�C�0��x	�C��y��:�st��<�|�VJ��"�:� ��#�5Y�T�{��z�q�?n8Q�+���P�|yf����S|�z�MEm���rs�����wsCP1��ׂ��b:��\7�.Ps�j\Q#��=�Y1i����F'QB��C��U��b&<9��v��o�R�r��7������)��.����lf8���,���o$����e3��vJ[S�r�p�o�;S*�VHygNzʌY_o.��G�֠k�q]ޅ�|&�_�b�}��I8�ϥߏ�Ƿ��7�aH�z���)ra�|7ǋ-�<y�κ��/����բ�%H�)�0��=����>�z.��3�y������Tg#dq����<D��r��ow�6/�G��N����d��x�6�sa	�Gve��"��w:�]x��A٫�#ٯa�
no�Kt)�gv��3�{�PRƾ?�"����[�7��Ѿ�[�o|�P4ӳ��L[>I�:�6s/�܇�Z�J�l���p�9���ӹ�����D��Q��K����9Gm����g����L�p\vE5�{��6�N��ߕ�rR`2z���:�iF��9̭�f�Ov6�ќ����.����(ݷ��|\���ASJA�8V��3�����E$�I��z����U8������3f�-fm_�霺����u��2c���ϲ1Ӻȶ� k����<Y�V�N��������9���Ã�w%l��k���=�N�$��zZ���Y:ݕ��K���/w�%��VǴȂ�:��L����Rd2;��cr*�[Pѝ��Z��,Y�e�Ґ�DFo4�3%Cj��.���5�\�ӱ��תc�0�.��t�Ӗ�X�
��.��1�:��I���{dC��Sg, `������֤�K5^ؒ�bڙ��:��]"�n&�����q>d-�.���V4�ҷ@��CM\�k�z�-�z �%�$ݥ ��MKA����<s/n��O�:�N���3T�k�c���V:�C\yt;I:�/~�=�f�c���Ʃ)r҉�j᧺�7K,�;Sa�VF�ӫ�;г�=��W�{���G�GWl
��Oc�1��g`�]�̧���Kؖ�v,w�KH��j"sv+t����d�}���:V%�ЉJ��s�>a�5�w���>�Ҍ�^ �J�0w��j
�$��*	@	oa��������Ϸ*>X{Z�Z�^��.&�Fmn�O^�9��,V�)��gW	Out=GMѻ����5�8��C��ȱ![���\s^���t�m���{P2�HZT��Z���Ӹ�hY/;.�]-`�a걮��H;8�vL�eA�718RHA����8��J�l�U��[+�����{R��C^.���6����E_���,�5����Coib*���<B�Q�Ўճ,�FLiG�0�[l�������m��$���X���ۇ�Nf��n���;���e!�̶�((��#6irY�nCR�m# �PkZ%�XMO�i��FV=��Ȭ��b��V1����y��|]M�G�ͤl#V&V��uĝ���Q�$q��2ע�O�M��u�ZNzx�r��^��	$�~ �H V*�"�E�����"A�����RF*��cUX���B� �
�X0X��c�*�U��R"�AUcUER&XƴQdPQT�T"��E"$UX(�QQYX��22*(�UUE�#"�U���X��QQE���""E`�	R�,�TTV*E"�X�Pb�(���[J(��ATb1b��"�*��)�*������b"+�V.Q�T�����EEEQA��X1EQ��+DUŋ"��"(��b,`��J#�+��(�EJ�T�H� ���j��8f�"����1m�+(�� �(a( �L5DZ��k�A$�_p���B0wR�u��p>�YZ� 3'u'+5P#y5�3ח�+�[^�ٖm�es�n�\������+gR��]1���  �����t��԰~򷢽����|��kμo�-٭�2mj��wj��y���;�C�P�j�<&�3^�Hׂ�#^�����5�R�,��՝ցT1[Y�S�e��6.���VM�;4��&:�#>�v�b����e��3��KWlS����]�p���=tP�3��H�����un���Jm����kk��wV�K����q�s��E9����;Yyhd\�)evtV댅��.�z�O�>O�u����:;�v+g���&:_k�y�a��α#���nT�o6���yI���<�^��a�%����B5��윅{�]W�6l���}����l۶����D*�"�$�sq\�.,6wTSZqW�m�D��.���:�7JŒ��y.�w�r��4�}^�uG:@�qV3����ws-����	P�Yf�;D��qslbUл��vdcj8���v�9jk�M�}�v��j>&�ǧ�#�ӵX�i��Cd��3��ge�h�맺����C�bg��/��g�6����;\zQ�tC�%��_.�=��s;������dp�� < y{��Zp�燂�{�d	Y�
���Ftm�o���J�>xE�Y�t�u�������=%��� �X����Mĩ�t	�`z&s�f����Av��Е[}�y��I�j7�Ўk�7��A�`�{2�'�sV?Q�qco]*|�s�������:��zg�̭`��q*��z�>]�Å�6����F�Բ��y���k�n}��*�Ϳrͺ�zcd]W��^k�ݶ_�8��y�i|����1x�ԏ���x�S�H$f��n��&��#��F�mW{���+G��8�>ާ������o	�����X:z�����}x�%�����,o��my#WBV�"�٤�<[�i�cܚ�̮gZ8[�����C^�>mՁ!l��B9��2�56Ua�mm���2�:�{�a�r���+ =�!2�y����Do�����A
�y���)��u����S1���.0���ZZ�u£K���\�%��JS�o�p�o`�>����SJ��-a��<Ý[����Ös�������}�5$�%G+�ʻ�L.}�d�`c��'2�C��R*1^dWj˄�� �t�Lr%kJ�G�W"��s�D�:�:�qt��nap=�h�Fஶ�M	3Y3���K���U�B�MX���	���������/�mj��4���f�tB����	Kl�]W�)�N�Va�K�'�gc��w3�m%t������J%3*طlts��_�6Z�S���U��mN�k�.��,)mYs����ĩ2������E�3Gǁ���r������}��Vkt��x+ɸ�40�ˡ���4Πw狲���t[尪}��x!�aP)�Ѹ20eVJ��P�����B�}A.��9�A��ڸw��P��rX���X	=::0%�����h,�`秴��2���R��O�g=�R�z����Q[����ؠ!w�=T��k����k�bu�v��Ȧ���h5GB�37����E8}�	g���޺�����q�����SoCS���Z�(�#�o-��y�Ag�%���R��ɂ��ً'v�Fgs��3 ��T�)c�(7��X짇KI�;�	�v��J�=.5O���d��<��+�G�&u#����<<"Sҭ��)��?y��N�F���sz{�-���ª�f}�MB|t��8�'�����ԵA��t1kM�gG'";[n��ڕz��/f�P�(�JE��k�������������q������&������D�W��P�%F��Cu��n��Ǫ1ڴ������;W%>�{{� CQ~~1�ϣ�n�ҏ<�U�S�����t%�`t��[�rW�a�U��y�Ec��Jq̄����<���g=��:�u���m��Vfm�h���=�����4��Պ[P������6
����F���-W�\b�}֒�bU�YOBX�cu�`;u"�(�L�A0"VN���s=J��,`�1kW�%7�mؗ�:[��Jy�S�L��]r��Ύwԇb1X�!g����:�`s8���a1޺�z�l�EfG��dH�
^t[\e\V]3b �P��*mw<�pO`Y[~��؊y�d�jd�1F����#2������n3��nl��`��>.��Bޜ�n��� �}��,�*�0����pO�{{�x��Rk� ��"��d^u��V_R��x <*�WiAgs����;G�y��+�}X��4�`�i�k�Uج�/�o�����yN{~���ྮ�=�r���Q��&��˖�nJ=�;�u�{q:�	~ǀ�\�ג7sZ����҃��#�/�K(\��!��'^��`���}Z���y��q��QV����_Y���g5؍�̧]�(���Mt�+Zմ�P�ąa��~��Jv���͝� W���<V�+vi��k�R�;3���!X��g$j�:z���߱�ڜ��z�fߜ�o2:75��z&��ut؞���6:�$df�G�e>M?R�YV��rw��"WOH�����2���>��!�Jg��#K�ݛs����x�${�o�N��M�}����}���}Nz�.(��Y\���];���/�5b�����_���M�����i���><�T�n��3��T�o7�{�_/]�|��C�ͧ�Vċ�aD��f �K����(Q}QQ�[ۡ>!;���4ʛxZՙ�����Fr�G2��w�-�|Ol��Ӆ�j�ɧ2�>�9�A΍��ש��<��-��'t�[H�n�������m9�M�����k�[W�M��yM۪h�Sh s�'^n:��^%�_��m�#�?]Q�V�[={P�����t�Bn0U���k���l�"��zH�����=�`��-Mi�X�h��9�D��:,��݋wb�nh1E!���^W5��g`s8���w*\G2n�۸����e0T�|��S�H]�zq��|�K}�|�"l���7���7۳v��iɉ��	h��Ju�5�uT>Ϳ	w�\�j��z���W{�u�h��N�c4(\�I�h���y�<�9��jE�LNӚ�|�j��R��-�C���QI'�]�溼�qU��3��9�Ya���=K�'a��3ȏy�b{՝�r{>S�i�'�(��t�����-�-���U9�V'&i���/jES}���5{�z�v�q'�<w�E�^z)��F��:iUuXz75�]�M�9Z��Dd�G!�=W�B��KcF�kn�k=�y�����#��^�Æe��=�U�f���p额:��K�=]H��}J9VD���S���[���/U@��Y��h��nQ�����k��n�uP�]�6wM����t�f_�/�z�E4:�&Mm�y"�N�U���κ�,Pu���W�o����i#WBV�+z��Lu�5��2)��m�2;�V�.���Ϻ�mM{)��uds��>{�f!I+S��*:q�{,�.�o��Ӎݞ��L��""�B�Z�#�(Pe>�Ue9�\���W�qr�{*�ux�1E�<��\�>Wy��u�?-!�����[�Ҫ'K][���1ԑ�+^�ƶ�Z�T�L		���li�C}��wU��kk:�,E2`]�:�.��Ԕu��t9�ٰ�ԅ*0ա�b�NX��E�2r�Z�5"3Ge���;��m�o���ޞ��8(��*&�'�3�t��=�U�V`)fߩz������{�{)��IaW�x+��<�J�/�u\�T���S �����x�n=}k�J
�f�&�hb�&��V2!�H�_�Ӱ�L�����>��]Jv�^��zzmu֓� ���§>�v����p��X�'%�V�Q�67��]9uf��f_�˦�փc:���8z��mE
u0A"��_+ke��B;�Iw^��Z�ʊ�(m���'.�֣�g:���F�rE��xx�k9T�cz��|!,�z↨�t��!!ar�A:/�A�1�P:n�u�kȶ�)k��03J��⸎��YNVu�w�,pY|�3�j'�5�S}R����Y'��K�1��9�� E�[Gw�4�Q^��ک��+7�9���M�9�A^/gs:g��~�UԞ����\!Z֪�[s��.Y���3��f�nCN�뽵���{@k&�uN	ə��f�BC.ڛ���ַ�?^�#�y��֊�F��M<X5nMR��^�tI�I~&7�I�z��v���Z�?V'���ڰ"���u&�k'����f�c�n�v�bV���E�Cu��}Lu.=��%+|�B�W��dfp�=ۚ�Z���sA��u,+��B�6�k;[�^Ys�e+���\i���ó�;Hr��'�a��Et��S��1����P�Ĉp�C���o�1y-�|���,��g����[�:P��D`d ��AB2��8�8�]�XЖȯ����)׽l�p��J���Ѵ��J�����]����-�|ԨͶ�j]k�!q����}Q�S�v}X��,ti�;qC��{�Ώp��S�l���O^��,t1�ٰ��^T�S!ȴ4ƻэ���B)7�EM�%eQJ��y]/L���6+E��$*qu���+��������J=`O�+bEgH�q��nq���L`�gA$:���"8`�L����K��XR̩1#��LUּ�j^0'�¶�*|g�d#�]�A��%��~��zן�e���؍$D�ň{Y}�+Lŉ��,��v���_�p�����n�	�
�g�^��{Z�B1��1Ph�")�8r����k��!o��Em��q��;o6�U��b�֯u,�U�����1C�Yt3�X���B4l�Fo1Rw�Y�Y��.O��Yܻ"��˝h�E��91�����g$�t�W�he�T��5Ξ˜4�̄�;Uј���N15g ��x���2bi���l��/��ˋ�������qf�5�".�i�G6P0E��@�S�������9�r����-�k�B�(S���ĜMm�f�K�Gk�ko���^���n����t����uN�n�qΉ�&9!���n���(�}��RD���<����#�ɗ
�nt��:���  ;b����Q�:�^/��"�&e_V���"���*"���T���R
u71ے��[�om�5گH����o=خ��җ���>GC�1��*�@�`uxb�n�԰{��\й1Z�R�rZJ��7L�B_+g!��\��)��D��uT{φU�\-����f�Kq�v�Zku,('2����֙���Y�7L�xdlD���3n��j�vRf�7w7�}q�w����~M�g�~�;���W�����{�9��T.�3b:\�="Bi�2�Y;�J�s*������\,�u@�U��4�\N�cL�y�e3@cwzk�F�E`���)hNw�z��`W^�
Y��ڱ[Xz8n˖h_Ll3�^�ʝ.ª���Tbf0ѼR(�գ:�^�X�0�/ԝi��Y�̐�Z���++�f�B9w�ci�e���2g��i������I�2Ӿ0{�eC�l"��N��(|,S<�Q�;�h��b�P|�W��:��-���u���)p�}YS���VCfp�R��
�)��D+�{#p ��"<*��/�����d��*�Gm��Ǆ��!��	G��D���D���0��z�䯛^C�o��@�3i����0�(��y�0��&�.|է�ՆƇ��n��9�,⇶���74̲rSȕ*r��(���&���Jm].�&��,f�.op-6v����c{(�,�;w��z#�3�s���\�X�X�kR�����s�b�]0��޲�|��FJd[�h#�[ܚ);�憥���3��FR��Zk{cSY��%�٪7��i�������M�;����I��lF�r��N�fL�Ŗ�M~zF���T?Y�N82x��U\�u�]��eѶ%�y���d��oLq��3Z������o�f\��$;!ږ>��Y	��=a��
��{B�st��I�SV��w:��S�x�j
��i�k`e��n4D�B��"�F��)[@Bl�n�*�5c�K-�(s`&��.��6�j���Չ��︻S����z;��9R�vk����.".��zN]:�PP�R�hvwtWF�Bk��1�;eެ��MU��fB&���"��ze�w@b�))ۗ�q�[��亯3W1����/ e��m��ڶ�c�__r-��
�'�߰ǹ�"��9���ʠ@���d�;���J���o��ѽ�r�\�M��<���ٴ�)�E�&����ۀ�7����T�9!;尹^�4�JCt��]����HL���Yf�lU�uR�ܩd�Yw�F��z���B�;y�ѕ�?!x��5Mlиd���(a>o6
`Q��;S�=�PC3sZG:	Q�Щ��^���l���
@I�#��E ��y��ln֭U���vU�`��ooe˃�DelL��Z��:1؂1���SD�@hR��F�կ���=�w��WȖz9τ����d���
d�v��Q�,���k{%*��^DNs��6��؅:���Z��hO�l���e�T���l�WM\��.����[˱iRGZ۲�ۃ9���ڗcd-+�w�t�g_q��[�_ڝ	[��T�%)`(z��U^�F�j�*�{�#�:W9#�|Ƚ���;|�/z��I�Ӵ�����������=��z���+Ø��)o{Z�Q�u�]c���T_�3��|����%%��� ��U1�w�+�w%�m]�Ϛ�*o�4����t��s]6�m�<T�K�v�\��0�xek�(�ʻԎBi�j�K!��+�IL��}5�g��Vy��5R[}p: �>��h ���p��;��&݇�Q�<ߛ0���guS4�D�E�i���i�[��ϱ=AZ��$�����K��x�1a�,�+Y[h"�b�UFD�!�c��DV
)��11aD�R,T�"**��c �
���E\5b�T�S�ő����H1Q-�`���b*��(�����*��VV
�DDEU�Uq[�"�Ƣ�E,��-�T�TR�jZ�[(TiUR�E�Z�V#����UR(�Z��1���b%e��j�b�Z%)QV�mqJ(���f�DTJ�QR�[J��R����TEcZ(�m"�F1DU�"�-����
1�"*U+�"�R��1�,�Eb����

 ���QF3
�(�QT��(�mQж�Dk%Ke���*Q%e�QB��� (���7�����2Ɠ�m:�Ft�lvإW�;Yֳ��(7&��2]r�e(�����Gv���]���ɝ%X�]*o4~ S֥�W4t���_e#~�ʾ����D.b�R�o�`Q�^�&
9ʀt�<N'�3Dq��N^b^�n��/ԗ�� O��sE�����ت���N� _=�ۙ��T�e]kٯ�'X���=K\ �7Lg�2�>�F\��hL���L�4[s������L��GY���Qz�1��X[��-zߴ��CѤz�i�@�8�Y�����w�)ewk�՛��4x�F��`c�݋��q��ކ�	T��av�=J�1�+'�sJ]f��I�x̝y��+��^�9��,A��1�l��v�������5%����.3�����"w���1��mɮ����GM�#��`#��*���iN�E,�sƻcr��tTXUzҮ|��&Q�je�p�9�e�*���.������٥#��H1�u1wC��Lb�IY�%���`��0\�NK�^G���*i�o�v�<�ٳ��d�N�OD[z�����;��(��`�fiq>�D��]�0D,���F��>������o���������PHjvݫ���̈́���)q���D���I��̋��#�q]�[��ׇ1�&��˔:���P�,�ׅVK�4�B��P�..�	�ݭ%��3�h���k3;<<��%���ݱ�����;wS�|�������xH�ڰ�����S�GXʾW��k�z�Bl]+�zg/N)��E�3����'8�\�MDK��m\A�su�.0�͚��{0
9�BIq�b�C9vPF����x^:�U�^m�r����S4�M�Y��í�G�h�����)ΐ�Tk��|���ܓ9�.��,�n�̧C�(*�Bf��"�O.�"=u�z�����
Gl��{�ϻ��!����PP��3��2⽜�LW�"�j Ԙ����BC{,�����~�1gv@����R�vҭ�S������̸��$�AI.}X((d����/yb����,$.ǪOLU��/fxvb��Y1S�L�x����֠;,*!�;���W�܍�Y��}~��3޵P+� �{� ���ǣ��+/��Y-�dPͪ@ձX&�&�u��Y1����_?B����7���J�� �~��k!��X��������jo-�KW#y�'��/9��!Rd�����oע���֦�"�)^.����]%/��r��f�$�ґ�x�%k���[<1��9khud]F�c+����F�ۤ*)���,�����[R��
���#��O��z���2�_2a�n�W�(YzD'�y������Iֱ+p�kk�����!����Hzk3mmI���b4o��g���� �e0��{��;?��a�m�a�:��9x���<b�z�x�UL�zR�n���\��Kڮ헴��mdb�~��*��A,����.z��9q<%g����/%��l�kmm�T�o���ZI+å��V��������gy�Ђ�EL�:��-�GT[��2؋w.�Vt8Q���<o\s�>����Ze`���s�f���SĜ�耏$�¡W8���ǵ{/Z[�,��K����V��񺌯emr�C��K���]R>,�Z�m���81���i\d�!�ef��s��9���%�1#|�S	�x/z�8�z߆N�?u���}��a���I@����^���债���)è�l
RȀ_f��i.�l}nY3oX�3Ն�,@��ާ��G|�O����#^�a$�8�ڦ
���E��z�TY�X��p�^�q
L�c��H].��ˁs���E�"�_��=/�"�����;No=����xЄ�",$�O��]r����KrG�O�q� n	�(�яbc���d�7fe"оG���/�+�%n�'��*8��zkE��_dZr3rd�=�c��4��؂ �ۥn>�dKصpR�9���E����ޮ��2V��*��;�H����g^�qȺv��bz�&P��k�����]ڝ��n�z(�eG�:�k��S���3�*Ƨ�ɠl�d)7X^	����]A�3��(N,{�wf��ֺ�uܨ�r�Κb4�h�U�V&�w����#7�z��"����R�t��X�H܋be4ui��`׳e�,l�d�4^�*��s�豎Y칀�4#�Z��#)j��"���[�ȿ`g:p}��E��e\yy��N��>��O������؋��50o���ޝu�U�:&�K�&�:��P#g0z�9���j糇�L?{��z�O�7{Of���j���"����3��lU�/�O#�c�tR�}J�1���r�Z���&qf�+��\��ʑ�s
8�e@Bt��(�\bc������<��u,9yO��C顐�_F.2|��e��m����,ӡ<T�[�s�5�����0�:%p�<�H����d>�W2j-�y�YU���0k[��88��R{W%On6��ފ`�'H�Fz�K4/��W鞸�
�(�����(��)�/ɗ�|'�����G*�>ַ�穚w�cL-�w/
�j}f_���z��G2TU�Ud�7��q��Ӹ5�]�Kt,,̖Q���Y�u�r��x27�>�:�X(J��M`�6�6��W�.vJ8Jڀo�[�ځ;N�)�]J��<  ;���ҝ�����)V�4�ҹ���M$q��9e{�����%N�YC�.*�^��ݴ�(ˇ�掂�N�����0U��L�n��E[;L�72#��>��}�O�楤�~J��SM�9�|�P�;��/��\�G���ZZN(G�2��O)�gj���n�.�Ӱ��ف:�DD��(+��N�
�"����n��o���2fF9��܎L'S�&(Z�F�ܚp�t�,E�\�J^���D�W10mUQkx��3=⸩�{�Bpz��x���xXM͸��4P��ZYcYr1U��j�x��n{n�x���:Mz��j�בrQ6Y��6T��"KqC6h�v;\�{�͉�C��c��sǯL=ݼ�+՜���W��вo�+�͈���ә�U��ׇ���"�����2y��9��V k�/\�1�n��m�5��8k��Z��S���r������{og���Kܮ1^#T8���5=���n�����R�Δ�U��t{�t�7����Wd���tN��t�:�6�gr㧏���L
48U4c�Y��ߴ����Vo�\�O3�؛�FL;�>Wm���v*t ؼ�ܧ��"q�u�N��a��Z�VFx���:�77��35N<�A�YP�=�b$��k3�st�:�X紵ŋL{}˯+��b�0��2z�UmPХt�1��� ����_9������?�ӢG�QEۖB*f�v��!�6Z��T��o�z,��ه���ώL>���Q:4eO7�R��zb�8<R��]y�(�OwM(F��5mþ_1��ilH��ė��UY���ֺ{@i�7C)r��s|���q�S���_�n5�vy�dx`7���tu�դHT��"9�a�"�e��q�_ob�\���:�Y�,���>��,j�2*g.��C���O���!Տx��wC]p�8r&��B�#���Z��Ib�%_KiГ^QN{�����a��:�N��>��9Js�/�I�p�R���5�ɻ�Z�ǵcfƛF4���7��tB�d-�`6Խ����^tj��Bj3�uj�w��S}���S��H�OM�(�1� �p�9����X<�7&7�w`�7sANj+�Z��	�ɐNٔ9�-0iO��J9P�8�`�(W���8�VC�n-�4�Xk�eV�'���a$,1Ra�@�[�]zUA��$쵔��!��CG�=B���6F��i o�\´w���ˮ�px�熓�~R�ZsX��P,��efY׮��>�X��{��Cǡ�p�p��/M�T�P���8�s��vr���]5Z|/#3P	̸UK"TO�� xg�J�f�C��/h����'j��etUy�[�A���g%��_�\J�)�q}�����[���oa�8�Ԯ$�'[��;�@0߁"귆=�-�"0.�l��~y���Ul�Z��6_�������-P����������$a��3PeN�R�om�uJN��_S:d�bx׭�6&�0�a\�ǁg����^�+η-ݕr|�x��iWz�
p��yl6ͽL9�Z��z}���+:E�jx����=t���\�wj��)��l�~�%ǸZ��YYF��~�(ؘ��⊈F�[�5�6Y�62i���	�|�v��n��D��u���k��4��p��:ع�<#�yxo���<c��oxtA�u����u�P}�<޴qˮ2��3K�f��v���@�����%\�W��{"Y�\U�===�R��5pD��P��zb{��d�"צz"ެɨ�o3y�.�v����~2ȣP����Odṃ��t:��߽%!=�u�W"޷=�t����Մ��A��tzU5��
�(��;�ڷ��k�7�ѹ�yg�5s�� ��pԝiZ����m�j��.��Qɯ�t\ҙ���PÜ����Q�$D�L���Y�s��BUe޿������������l�k6ia��:�Nwۦ�~�� lީJ��[�"p��J��6�l`�:n����ª�ڍ4����,�8!��T����G�O&�ym�A|
�XN��K��SR����uSf�B5������9U����ܪ��N�a�8I�R�ң4�5�K�=&\���G^ȥ	��|J��s���ڳ�l9FJ�
5	�DXh��N ������x:�Em�G�C�z�}�23/zv�ݫ�q̩~ah��|1OV�E8Ȇ�Y��vL�w�
NV�N��&𼉢��Dc��Aj[;J]\����j�̉b+#Hb�E��άOk����kC�gί�ۿU�r�ՙ�V@��+� V�0&p�έ6T�h�e��� �<������~�J�(oj[%/$�Kt������B[G=����Z�����#&)��ʔzsi���L�����,X����}/���򷰎���j}<�,�y�,�^�)5�B�S�T��4Y��zvD��Ǳ�ڞ�X�t��%�����G5�]��2�K4Λ��X"���&���i�)k��ڱS�e%!�;��9�ymܮ{�}���tg{9
����S�4�`R����y A���1����B��u`C�/:+����<�]f�H����!�:�&g%��t/�MR���)��o�����޷+N�`s��Ymj�����*��OwR���b>��G^�,�����v�y�v��J�4%@�s�t'���ឩ��n!ڥA����#K٠����C*�p�C/���y-���Q}��(B�֝��]Q�|0�\,9��!�l>��:Ξ�E�o��>f�:8^��Nyr_����O�ra��(6#��Bu�Dd9�p.~�Ķr����s��%��WXf�<畚�v]�?vR7B,�z)W�T�0t�l�l�%/	���܁�����:s|v,���Oc�Un,�"��iΙ��������cc�J;\�"�lE�Y�!�WVjˇL���#!��n��A	ř�Wl�L��}�P`��N5�ϴ=��A��;����3�~N�O���� '�'��	��F�
��*�)��;�{#��i���Qۥr�ے�����5���I2�
!ys"�������D�B���vV8��H�6��A~�؄iI��X&'ב`��i͸�vM/�8YbԒ�_6(�h���sk-׻�ٛ�=׹:��.1�te��R�8}�\~· v.�	=�u'���8s�q���.��r-y:�	7� �5w>���0��g�p�`�&�A�|��}H̹�����qꂴ�D�~���p�.�mM��u�eW`�s����������ԩm��F�.�ݩ��Y�\89+�t6�CK�bk�)S<�J.3sp��炢��bZ��Ri+��ǡ�eV�-h=���h�o��p���F�W�s((�h�R�FV��n�<�L��v�.�!q��:�1�v;��N��%���A��w�t�����{���KP�%��@���bA�E�Q�)s�:YJ-��VҼ:Z1Wk`�r��{d�����nW�̖�m��Bܒ:�R1Y�s�#��*���IF�Q�����,����GVo%�*�R��	��X��p�^\OE��F��T;,��(�Geq�ⲝ.�י����v�oa�(��B��S�uv��.V'%����x1S�C���J�Nwp�ی[mwA���س����ա?��S�~_m
�Iu�'�ɇ�֟/	Ch�X	ݷ>�]�k�c�Z�r�Ϋ4-�f��Q�hI"Kp�ň�r�/���-����r�V���l�Y�4��m����T`x��wL�9a���D�&��R�|��u|�N;Ȓ��7y:ଞ��R���=h����-�:R�Z�n�w#2KcCe��间xE�E���(x��e#*j���sj��-4N[����7kUk�g��]uv䒦�~����{{��Ӭ)�\�$ώܝX�Rȧ&���<�7��U؞N�����O�a�HZ�,�#		.�"�mtE�����:��ٜ<v�ٌ��ch�V���6Fa�A�i(4.^ŗ%�������w���O�ϯ���X����o���\~�u6�P���81�1И��X�",4�����=tX�o��ʗ������«���n��Ö(�>���xR�RIB��-�wu�5��٧��u��t��Bc(]3ټP��y9@Lw����D�y٤��)�˻�E듳OP�!�o���#Uz¥7�G�܎q3o���KNp�������<�=��n�!�S�(L���[�cQ����#��8My��u	����`B��cS�=��~���aK+~w#c���):b���9 u���pl?���
[P��M���k��wI��ڕ(r'���V-��ޙ>�Gj�P�Qͪ�*f�5:n^�G	�������S?3��h�E`$1��ŠΔx���/�tsp����{�D�D��J�G�zˣn\�+;x����9�}W�Ƕ�P�$�{��eA��X�g3GY���y���ǖ\�ih���\�,�ȗ���6���2<�;����cܧP�}��N)w�2����P�l��q��3�z��$��.Y���]Cq�}(���t���"$}�^��:�$�E�i��.�b}f,��ͺ�J��م<�{v��2�κ��n���3��t��&ӵ���V�o�jp,zU���s(���|ڠ�;9�t��i>�,EK*(���0�1M��-B�ˤ�,`�p��fA��'%��xB��w�����SH�8�������oG3dz� �[ ����Pu�j�#-�Sjvz��Rx���%��+MgzvA,�e��Z�K�v���3�x�!b��Χu+�#��S�\N�Ө��	���z��j�u6��n٥�p������͎G[��b�<1 �<���^��{&�����R�Z�~�)\��_M��c��YG���]�b�Vۺ�s�_j0���zF(��Gu��k,�#��˩$ԩ��Q>:sm)�d�͂n�����B�[��Lp��9R�r�<�JFu��d���.�/Mc�A˹�!X}�Vӭ�{���+{t5tw��:��A��!m��j�	�\r�*�H��*���X{��s���,�����A7{���;w�J�c����1S��h���{��^ss�V�R%�C~ߺ�V5����bE���;U���ݸQbo�Ō�(�����Juf���<5�l���٥ %9w_]Xr�km����KF�U%�6�E�ն�X��+ʭ�����*(���UU��"��ZT������*�#+,X,dQ���*���TQ�mU�Q�ڵb5b*�)eQ�m)F�ZQbZ[ec���,Q�Dh��*��Z֭-�R�Ա��+b�֥�X�mciim�EYmh�j6��Kh"�*��Z�J�EFVZª*�R�V��k+UV(�B1�h5�È���%X�[��+V�PU�Z�h�łRԨ���(�RұDJ�UU*
PU�Qk�e�1HR����eѵ���KUV����XVU�#[e-Eb1H�JT[-���-�F�D����Uh�U%-
��J��F��4����\lN��bo	���h����b�hG@�Hњ����74rRd��	�:{��u}��WQ�}�r�����i�>w�kZY�O~��*)g\�[�n\��Z��~uXP�$h
�:ȜuWw{�'!W`�Z��3:_�E��Jބ)�Q���8:� �w�A�~�^�Cʮ�������/O�<lfY�O����۫Q~a��)���U�����x�?�g�x��e��`�{pC��Ν:��d���7&+�䘞zez�3�l��ʳ%[��՘ϼkyz���y�Ȓѷ:�[��}\����P��d�*�<� �� ���]"�6r��Ќ�w��i����4�u,�s:����Ys�J�M�N�� -���U�X#~^��:���L��~�6�.��3J�nD�̎8nxHc6C�4�mP���a����f��=p�]t�ȶ��m�`�=�����ÝKC��C6Y&��ґ��`N�bw��K~ܢ������^��z?F�>9���k�
���6�0�3��\|J��ˈ��E�����'o����{����y.T���P�y�=�6-�C�ҍ4Yu�c�([ƽjTB7�s�n��������|�Z�4WN
�+��>�u:����C�Ϳ�R�M���5E�l�Bm��ǆrx{�]겮�<3��'<<�=5�n�;�9�������h��b��,��֢e�5S�d�3����Ĕ�=�}WvJ�³���\Ak,c�}[]���W[���[ۮ����w�i�ň��8g�]=�(�5]P���T�l���E�R0�b~N�^��N��k����lw�f��Y�j���mq^r댼=\f�T��m�� ��}槣��V������ـ�:t����T� �A^]���n�E=2�H�OJ�!ȷ;�ݕw�S�ħ��6�"��S���C.�w]1�!�6V9�]�6�w9��o��/+���6u%�t�H�ӎ�������x�y@����^����+��1o��k�'�����s�<\r�}JY��b�!SB�!��b�ر���z����w�~{�}�L�*����������,�6��$����*3Aߏ	���K�=7�r2oi����&׹큄����pU�'��E��
4!:ȋh���"S��4lp�Ҏ�=��a���]&,�:�I��s=K!�=�!�#j�:Aq'9���\F4gU�`�pW<u���SI*񵡸7Ԋ�9n>'���O���W�+UA׾N��<'CFNiCrl��$�6�2*�WD�U�:�&I���Xw�VvCz��.�V��h��/9�ُ�ٔX� ��S��%p$�wP=�;�k��=�(E]Kz��B������ˣ�fGK5����������ⳉ�ؘ2�J��K����{qVwB+�C ��Q�2
#6:�Μ5��M�*P1�,���Yd�<]�yP�Pz�����M�O�fns��޵�865<xy����t�fU
�U6�L w6Qq�ˉ����د��Wc|�65�52C��� ��G��/=n�,���M{d�%#����+??P����i�K�`Úuu��]8b��{�T"ЗVB7���G����B]C�nc�`�E��Nm.kxh�������e3Vu8��(��H�R�[9U�go>S�<tO��fE7��>�U�'�/R��<�t�\I#�yq��@v����_N$������D�=C�X�c�6|�ZnvFm����^No��4tka��^ggݬ��s�L��!��vt�]��z��f��iPj�Y`GN�P�"B�'���;�ᰡ����;*^F��!�C00�{�}cE��v_j��<<){*�U<��j.ׄϏ-�|2j8|(;�ّ����z�.�.x��(��2(+�d�,�0�WN̦x\��u[�-4ɏ������2�F�yO�{ԯAL�շy8Cz=����Pd	}�%��gr޾Ur���P|8�u�u��!t7n�9yboQ�4f)x�5�<\�k�Z�:��e�K�L��E�s�n�ڎ��[j/L@=Ԓ��D���x����R��]����7��؁v�lH4�#�B��l�c�*f'�UEB6�YE��ǂ�n,יL�&��;󫜀X'�����^s�����L��S���h7��ᘥA�6G�z�O]\���^;I��Ѱ�S\-�p��o�ר�W��)�A*zb*E뽛om�7�H��`�U�Ϲ^Kڙx���z�,D#��S��E8Yb^V��:z�����g��VT����iWi��N[Y�@��|h^/	I+�Er�ex�2��ڧ�7�������FQgx��bFZ�W6��>C<�n��v�
�{e�3�ߩӚX_hz6���w�;�:���}��B�A��,��X]G\;5��WK��ݲ��h![�v�5��Y����~����p�YN�WS!3F�QCʸ�^��zs��p�k�\˭8J���]E��*���wZTz��VtDq����-�#�qZ��Qv��9-�|,��rVq3�� <8������nY��y��[�b�pe]%���\6\���(���\<,��E�ˍ-Nx.��C�����(N8���S�¼�s,Hw��v.�S
;+�')\n����·��P��cl7ծ��T��;�q �m��	���{s�0��#��Wq`\B[�<{<m�e��eq�-�A��6�յ3qw4C���M��/q�9�m$��8��q��:�!��:����0�ʈ⇥ͨy�6Gf�N��O���mJ�֥+#�	�;س�)EL;���"B�>�D�V�m��^>�G�������Ѿ��X�_�ϯo�\3��ѡ�C1"^�����љ��d��齱=�hL^$��cr�6��n���ˑ��m���ڋx��
����o�;X:��7"� �{��Ww��'��8㥎\X�\>�]���<�v?���j��g!��?4��wn�����;��C��v%@�>��G�Q��W!0�s�)SU�X�%*�_iu��-<Ղ��F���9S
L�8!7���#�lJ�F[HѢ�8�`�(aB]�L�v���IgA�Kl�(�<ʖI(�����a��T:���i-�Kƥ庵	�5U
��^[K�WFG\?2xT2����P���	�x���o\A[�Kɉ�ٹ�n܇H��6�h弹g
{T�T���p���#:�ě�oF�8 �9W���^@h�R`�.��A��t�f��P��ш!���nr��;ۓ� ��3X�[���p�uc�_l�!�3�fh�݇[(��
�w#/hM�ֶD屮��i�SV��w�����b�ڕ�O�P��]�%>{�)xz0�K�j�@=�9SBe�qԷ�{���
�1�Ɩ�_ީ�V\��D�"E�dqLؔF8��V��[�ٞ^�.����/G�]4�a��ϣO�DY~���VUi�^�'��`�C$��ґ�
p���Z��`�J޽����z���8�e6syf[���@xFc+JU:��?����*j�;���΋����hM��V�B6�ڛ���%8���sLv�z؞5�R��]{��fT��?>	1�3��B_�Ҷ���Z�P��*Q���%Tp�Qʆd#|��0��]Q;<��r����`LzU8�oiV8��V�����3�ͻ�LGY0,�7�Z���]�ڇ:���oYY� 4?#\��eu��ӪĚ�#k�]���)ʸ��.����ldxm(���������� U�\�,�"��F��2�T�F��#��M��t�0��U�-!���{���o�/!u�ǖ:�x���'b*m�5��E:�D#��3�_�<ٳb�����E[�P�)E������ʺ��kD])D@4�Y�&$+�S�|#�k��XNc�������~���:=ǙJSݩz�@���u����ث���֚vY�gYR5��$wv�v*�tsx�1ltb6N�
{�F�/t�U����*��	�m�K[ʼ���Kr�K��=�-�	w��V��uՋݖ:��3�XOd7�8�;��0�|=�۶���������o��O�]�iC8��%L38��X��[#�y�Լj#�!��fw��b��S�dLuk�1*C��"/��8f!�F9RY��U�Du���k����5E'����,T#�n��˙��T!} ����@c{�	�`����o��7������"E;C��{�ȃ5Z����g�V��`����Vs�~��Ec���[E�s�����r���7DA��PdFl;�Μ5��M�J�e�,l�d�X��L��:x=�y��\�pk��μ�_�>�����u漆��D��Su��T�k6Qq%9\V'K,��Ô�U\r���S+ }O#�ku�s�� 5k�% F�c�V,�jet�IзV��=i�jQ��mODV����\9�,���s[��}l�-̗hLq�N�I�8�lV��MN�I�.8���ʈ��6ߵ�,؞T́F�w)F��tiXmݐ�WcX����Tv�<��&x�z�H�R��Wڌ(��Z`7�|��g�	s4U�I7h����t��DO'ݗ�'�N�'�ʊC�QU�n
��A6N��h��x�㼥Jܛq���ѷ
5�\�S/���YNれŻ8�P��#��m0�L3w�r/�WJ�:ND�863�aǫ��p�@�1���J�K���iu��������}�&c����>�@�9Gb��ƽj��'�=0�g�1�.���rј��=I��⼤���r�]{ 3Q��)�:�1\Ct��d9�vT��3�4;M���������HF>�,�7W�N��,���$:�l@��ױ
p���d&���R�`��r��]ildib܈�]Un,��:�'L�R�`�~�E�+�f�
�3�NY����ԕ��J"���o�*���3�� �f+�]�4TT#�`ޙ��#Guޖ��7�I���Q��Z88d��<piߕs���N��1ү��g�x�ܽQ��s�� �����LW�g#^����d2��B�D ����Һz��IF�V�T�򹒸Ca��$�/����WA�O�A�?d���&xg���������+)_���]�U���;����� �9�)]F��O�W��&�eĖ�Q�zR(�-7<�S�b���,w������{i[�9k@���x��/>^�
!}�螎3�[���dY��(_:s���n&�f�����̚&ѭWK�/�V�S2v���f�1]�u��U�[�8;gU-3U�啼�ʭ�4�/y4��m�,���<��.ͫmɉ����^�6''7��l���Jn��3ңoF�����:h-k{H��U E�(��H��u�ٯN�wMF����~�!b?:��tl@i[-�ۛ��7��Uj�~��T-�j�:�Jf(5U���zq�)E�{~z��]��̂A1�F�o�T����Ό�G�i�#xd�cE۞<T�q����h,�&<�ߑEΓI9]$�P$(��k�_��Y�D#gC�F(
ۗ>]�G�������B�������}���t����Q����e��:���р<��n\چ�T8*<�,�s��C��Y&�نw^�UX����~-�L+���h���{\��B�fL��S.r�z�p<�S���턮�T�\`x���׵ �C�E��[�$Te��vo�$��=T�M_mu��z�h�<)�*�͸�ػ�nhȠf8�7&�⽋�̶k�M�������Q���^ˣ��-8���%?:�u ���be�Q+���Wg�d�o>躊#�Aְ߄Ba��oB�(�X�uQ�ۅ�&a��<cC��f�=���wa��s+C0`u1�����8�*�τ�^��_���>��P�c�|V���T�Hԋ��B���sȁ��YɆF��_+���S�è�w�E�oR���M�%h�|áE�f켻8ެ<���-l)曈�:�I��;��u(�F?xzm�&�+]��"B�T���慰g�|J��o��8��*�xe>^��m#F�4�ZA�=�s�:hg7�n����YR!

$4b��s�b@�a�Rk��3ٳ��f�d�u�)�#y'y�ۑ�tڼ�(a��r�8d������P�q��]{��o�+��f�3�Ż����w��῾|q!|���|��+	��^��o��>�V;#���+�+�s�v��a���z{>���p_���ȹ�3JQ½��
�5��2�[�\Ŕ���kۮw��ƳV�^�}'tm�>�n�[T��d��ۮ���EӦ�I�q�E�"���S�b�y�-���wE�=]�^�ڐ���l���K-yl6ͽLN����;ؼ\E,7��'����Oc%�:$�x�	Yl�KP���ضU�F��e�`71��qU<�o�u��y�����dF%����5q�P��� ���p�F'�Igjz����C3W�UC�����y#ۅ����#�J!�8�ƹgVy���7�]q�:x�.����������x �CN��얺�9s�������og
���U���%�Yy��wȗ=V��l��Zi��wm{vC�{�N�������_�͌�CQ���߇X:��n�>�pL�֬}7��e3�E�>�8��}�]�F�q��%2諘-h��Y1����l��c&�k��+{*�ik�Z��W��pDqʊ?���rL���@��}��,�o%sՐ��S��f^TN5-��&'�:!]O�]b%as� �R��:�[���ޑ%�X+�H�t�V2��ͥW��삅��p�6���tB�m����w��wX��0da�wA�����ɏe�d��{_@S�雱�I��}��Z->�&58�}�^�}���0���@d���m�NN�<R�VЍ�����9çM���B�J����%P��X�oL��N��] hfӤ�Wxn��|U����4������'�������v#�τ�*��d+�£����I�z;=��L-�L��X�>z�kX�a$wJ��M��\x阹��s����S��;
���2�+^�9G��	pd�a.{��A��S�n�LWgf\�$:u���p9��� uc�nN�|��o3��_Ȉ0ĕĺ�\�m�2���t�{��)�Z�z>�J���3i�Kia�r��������\8�^�N�.�iv�E����Q�"��fn���9Vi���w>|̡��^��8�Ο8�n!���L��8˼_h�^�}���|Gn�cs_T���v��/0n#qܳ7U�j�R�Qz��,����^��Β�媃G�g2
tފ�)�ִ�=f���)}t+L���cq�ȫvtkMZQ�D��5]����Ro�oݧ�7�n.� ��R��{c�}�����?�^��;7Vi�[�תWobϒ�G)h�7�-t�� �ڻ'4oy��g�؅ͤ�njV����<�_N�NA<}�c7Cެ�l�&�35ei�um��E�6u����'w�{)�c�U��(�ޕ��Ʊ96%/��x����f�j��t
e��o�L���y�M9��s����cwz�W�_F�N�1J��xn�z�d')V��YM')[v��hxLs_b⠋���a�����1��6qWz]-�ݟ�P�^>��|Fq�����^�(��WӮ��l����9"%������N�Fێ�X���j}�˨G��ih�-��먐�+�L�l���j�������!�ǣ�ht+�k�I��qj=4�t���	�e�$�g!%�>��s�F���o�w�H77��b�*#&W�i��~Uvc����pEz�c��2�/���5rE��g=�H��0&h�[Б��LE��|��T�iݻ���<��&�\�"[Ε��#c_��@��uL�l4�y�-
��/���9TU�����,����^���F�ޝ�$�;V�*���֏��Q�c��zcU�k��
�y'.:�t6�I�F���Է���g a!Ha��c(j�qua�-N>��Ν�"��}o\�������ť*ZR4��Qm�1�V"-T��ږ����D�T[VҔ+iQT-�T�E�QJ�E�EeKZ��U`��J!Qb�j(�6�E�*��`�Z�X֣0�ť�TV1DQE��5dPQ�0�J"ZUJ�Z(��������E+UUeJ¬KZ+l
��
��ED*Tj���+(������1SР�ֱ��-�[�(�ڣV��[Z�1AE�e-,��U�
6��,Z�"ԬV�amZŠŶ�j��-�k8���V3��5�U+��ԣZƖ�JQQ�R4l�[�*F%�j4�l�ZЭV��2��-Jc�Dh����KU-*�����ikD���m���[kJQ����щ[b2����+iFմ�m���BEJpz�������������YwwR����~^�'-����e7��ɏ{{��I�p���+N���=�s�m����f��W��?N�&�n�q!�}aeu_E�uPz��#��з��N����8�⼵�MX����3/�DQ��(�4#���=��&Q�s�c��E%=Q{ؤ��<�O�ξu�y�vX��w=qB��sxR�w�ZKS�C�uO��*��֬t�^A��.�t;�5{���Q�.�`�~�,��T�4�V ��C4*��E��XN�>�i���ұ5�o?u���ƫ����@�K:���MUs^	�	ץBb��^|�C}X���B�s���uOxI�̼3%׫�^@}�u$)j9;،Y8f(K,�S�#���GԶ�G���M�L���x��9щΗ�Y���C�}{�d?�x�.��X���r�r���|@"��AdEc���8��c*���d+�r�
�CF��f�]93�;ה�2fDY�(���c�;dr���r��I� �ڦ����q^͖X��,�5�\%�+blG4�M�5�F�׵cpj��u����"2��!U�Z*3��o�z%��33gU��o������%�׳�e������=�W/�����"�]ܽ�@�vp���y"aM��T�֯�H�bV��۬�3�B�v���W�3�#���P74�F`��}����j��+CZGFӯ%�x�o:���nQ@����=�Ǆ�v�B���d�8�����*,w�W��9a�<�9��t]C8g41W�!�P����F;Hds�|�X#9N���q5K8�:EԺ�0����K�s�̲�	u4��YZ���Y���e5��bc��bB4l��R�7إx�jq��I��z���Lꋓ�3�/�5��cTJÔtX�G�\�jaq���:2WӁq��)dܤ�NWE��vM�̬�[ӊ�*�����Fĳ(�����8mL��b������kì�S��-W���e��cֲs�W���n�u�\C��B�5�n�؂���_M��꛼��8�n;kW1[����k��Y甍Ћ,�'�H���0(M����B�6�g
}v�M�����R�;�����K���ł�(�6�֚�[5p �?om��ƻ3�_o q^����rK��9V��"��gN�	Ѹ�DP�n����w��_��E��;e�0����'<�de�ƠᲕ�G%5�h����sN;`�p"#��	�A�HT�f�4Tj�z>�������qxD�	Z���V҈M�$�Z�Q��=˨�Ln�*Ƿ	HD���]�q�䟩�f��@9���]JY���{W��u�����[E-�����-֕ �/[�x���q�h�3�o/���`�X�m>�/�t�T���^��)eqP�� ڏE;�S��D��X�
]��鸞�:Kݼ����t/ٔX�����F,��}ex�b���$Z+8���8����j��S�a�0�o=H���������E},���nm�\IB��,�R��q[ɩi,<t('X�TDRN� [[[�9�s�c^EI�����LDo?��WB1�q�k��7�].{����U�=p��T������{�;���c#M}=�x�X��nE��f�g�<Q�c�,��C��̕t��p`�͔TZ�.�#�4ߟ:�/��^y*�;5��팖zZ����]8ԕ�Tak��m`o���C�}B��|�K�c<x؞(�c�t8e(���S�&��JV���v�����<i36�ĵVt`�Gz؞6���JF(d'��Ven��8@��1N�cё\�R��Wq~�-)�[����t:���ʬ��L���E����_;YM�{q��#���Eۉ��)Su�!܉�f:V���Z�G^��%E=�]U�wY�J�N��"��/#�L�޵�gqS�O���
��p"c�v��Cvv�c�'PA���$y[�<O��O���1�+��ܖ���yы�� ��i!�p�\N��f�7�����Y�J�b���]m����9����n�\�7e�JuC�mS74�3�(Ί�����|�
g.054d(� ��/��9��\�sϖ8h�ڼJ�Z��ܳ!���F�����D8��Lۀ��ڎY�վƽ��9�7�Nř���9�������-�|�9�`����s���
a��l����RA�ڼM�k��:;-�0eѪd iC�oB�r��8*�!���~v���ҡ�c����{)}Z,u�#�Ȉ�u�^G�K���)�֕h�1���νu\� 5�}����[%���͝�`1tW��CaR�"��1K��O�:����t��ő�%>�w|���������Y�02y���P��d�{���0��
��nxuI{ݡ�7�"��[��%�^���F8b�Yr3z�D��:,�M� ��ph�m�kq��|��b���PP��ڝ5V��9T�!��Jf�P�Ǵ+��B������-���&�I�����k��������7��:��S��/�gp4����[��{�7��>w�&0�>g�X�ux�;�K��F��&���|<}���he��e��mP��M�¯�����]ս(���5aRfi���ʘ�����WSYG�_,�n��҃�3S[XNj��Ἇ �j�M�q�bv�.��]�����s���5��ec��]��t*����z�^���U�v02�%���G�tv"ȓ��t��_-B83����[�.�W���-�����R`�b��_-�BQiK�F�N8�ѳ�!+o�*��lELP��PUG��5k2�M�q3=˒��@fـ�]tB7�8��]3�|�;ͮ:�Wj����U�K��v>�S�X\��<*𳠰KSĜ�B7^��Ի�*z�l>���qK��GG;'pQK0)�L��;YӸ��W���%O@�u����:x��0����5��T��)�<2���f�B<{==�1�9�#����k/x��au���
^�:I~X���O��	�XR��n37(5��m�BwC��Nٷ�A�RȀh*�eI�Rk��\���#yn��31B���oW��1�:�C�l\#U�ڦ
�yS<f�:K����`&�B���n(ι��������=Ui���N�-��"a��PbT�
5	�D[Fp�P�Y=�iB}2T�SmP��,54�b���^�=�-��㇯�����"Є���^��bsO�I���W���ZyQ�Vf��B�C()'�{Gv2�܄�6��|C������)���aJ� �������b���]@���t�h��1�X�Vtg�Cx���쑡�]%�|��9tׅ�=/Ơܪ��T!�8�b`�8ȀXxl�2���K�*-gN��{��-�ui�>.���-�����_�>%�?	Yk��`�S�Pv��?8�_���Iu�7�O#YbR�؆aÕ�L�F��dfô�X�L�P_K^��׽�M��yKb*�v����/��j�c���k�;q]W��R��Ӱ���Q�B�O�z����8Ë�s�ԫo%����(��XD�{L�>���=��t]9�9����A�P�cՁS;e۾����"\���:J�\.j�Δ���]��K��F��~�s�LG=��V��X�8\i�8S0:�*Q�QǞt�0�S<!�����dm<.qt�:"຃��|2��2$+C��t!ڐ�OG�C=�b�ʨڮz�[���I\�QS��GDJ«��fX4!y���a�o�E��|�:�|�X9��Ӫ��q��v��*���y�Yu���5��W@Ct��d9�%^pk��<�⒜�B�[�aj�Qӛm��m�>Y��gC��=���Ry-��b�D8)e��Q3�u̖�[@6�[�M�E�������!��g�v�(}�Z�����͹��V�����n"Ѳj=^����6����0�����{O%��.���Z�����Mo1�#Or����ϗP�L<�a�v��8�j]pQ�B�q�e3��dV���Ћ4�O�<�|ŃO�;f����b����$x}�ҽ}1���{�KS4�<WES�43����B���8�v������k�N̖n��2([;L�ݘ"�k��Cz������4S�3<,nlԫw�L��n��ΑC��0{Tx�ƸZ.�ƎӚq�`k��HQ����T���z���o���8f�`�dS#h�\<2�k��u2��x��q��lʖ-����yw^~U�9��8]�K��"q�|�/4�K�e�*�a��b�Cӓ�L��t/��r�A[�N	y�TDW:z`5��S�	�5�\��i� ����a��-�|J��-�y�>��JQC6h�oےˋ
����M�ҷfw��'�,-�~"Ŷ���E��6ؚќ���*:��WT��5�ͤTg��G#~|�Ǔ�{�c���R����V���ir�8��æ媽���:=lP�W�2S1@�p�������9(�G1N֫�v]���=��j����Ѕ���yW��33j������p#�]z�j���3Y,��J����=2�=7J'��z�v: �3����,1}��A�St�G��+[s���s�Ώ)7祟'r��4l�VP�2��b�ۂG\$cB/�Wv��-��=U֧6WN=ᦜ�^��/�Cp5@Tˡ�(�ع�Vtd�8ṃ�ˉ�6#艌*����޳��5���Qt�n'���h�*b�e������9BR�T[�bG��\�N;km,�\Ҩp��$b���ຠ���[p�������	ǸYe@�F�o#�s��^�����|%-Vᜥ9�r�׶�2*g.3��4,)Ś�3����4��;ou�� �o��'�8�0K7XPF�}{h໗=6�o�%<k���>�ϯ�R�Lj^�/���o��t��Z�#��u.$�T��\-�p�_Ҷ7�
t:#!�PeJ0f���f��x��Q2B
f�~�+b���d?0߄Ba�V�!��џYূ�xQɌ����|����s&!A�������(����Q�S����>_Yo��s���Nv^�v��,,���IG�`*Y$SFnLW�Ɉ�+ί��g�t3�--�E����i�Egܛn�����d.ca�_�g���B�|���U�
���T�Y�Lg�v�)���O��gu!����w���ʜ8��3���L��V�p��;pf�1�kGN��xg���q�����xi��i���o{�{�=�ږ�Җ)Hͱ�B�Y�����%�$�w��I��DKFE��c�a=��ygF���W�j�����kT�,!�˹��S�n��UEڤ��pň\қ�e����b�ߚq���q�lwb ��!V�c�2������-���:��u�v�n52b&��n���sZ比h�;P�>�f`���9Y�4jО5nX4l�Lu�Y��Ec�Я�����a:­x4�����j������R��yl6�҆T�Z��n/-S��\����.I�Pޠ������Y�U2��J�8N\కk���<<��[J��K�y,n8v���+\���f��#��+o�*��o�J3NIg��6�b���m*t�_>R�Ѐ���`6F�S�r���3��5p|��r�L�ڮs�iDd��,\M5u�񮾓,)� �^b8�Uě!��0�}AX={:��I��L�$�ӛ�����Np����g+t̚|D���Dl�<r,DQ=��z���~�׵�k"���A����^�EqNị��� ���:7-��>±���<���j
%�8κ��7؞���CCΔ���[{E؝���ub��GoFs�x&�۔s�[�H�d�Sg��w�{(:��Ǽ�m�t�O8%uh�3:����i+���N�K+�ػl8u
���n�������a�?-P5�R���䛏�vovN�&��]ceR-�5�/ԥ� �U,�x*3A5Y �ᙈ^�Ƽ�>��4C[F��'ݻ�XΤp�����h��3�T�VT��ߛ�p��1���r[:�d�`ٌz�4]bz�������Mґ�B���"�m욇a��)j������)��J���Ōn�F��ZƇ	��o�+l�<"ʞ��Y����5P�W��B���}s&��q��ː�=\��5'��4�ʃs�蘞͜WH��	r��"�0��^=�(�9Y��nk�R,��l�ծ�!6n��6ƣPgő���~V2��9��4a�{���G�)�:�<I��ˠ3�X��OT�7u��ʐ���#�!�h"5Lbe��h�^N�45��/.������\5XD�>�{GK��x�w\�:goΉ��Ў��������omS��.Z��;0#:@�R�(oK8ܢ�͑ej��ƷK��wN�(ѓ�QѓYB����v��#�D���A]�|}����.�:��}���gE�i�\�>h�p�$M� <����rOE�/�b���m�dGR�H>��2c�@f6(��q���m��qZ2���U�����&�P�]����J�]q|�7n���;���!��~1m��}s=YP_��-�/ku��!��wR�d/�S5�>:�y}zZ9ǐd�݋�f�G65�[у�w$7�����ه{4�! 6o�����4�ʷ����q�ݴ�̅��m%��,�W��s�ў�g3�o�w�uv4)��ʴ�
4��)	Y�,��q�܂��J٫M�6�N)�8v���I�̞�|[�s>�Ԕ�J'i�
�o�պ�?h��֭��H6Ed��p��ę�L���C�������!r��Ey{t���A�muwn<�8GR=�,��|�-�E�S�j���� ��>�K�5��Y��S5���h85��B�`YR�wN6۫���7Z͏�o<��d���E۶�u@ɏ:���b�Xtҥ��{��&�U��ϗ;������9CZ�V��͇V�;�#���M��.��U�銹��VM��G	�U:կ��o�u��:⡷/%�]Fd,n	��L�hu:�ڍI���vP��,8;���˛�n[�95��d9ׂ��{��
��5`���Z����m]�}9��W���y��1���Ɖ�$Œ�3�V���eu���+}7>���i1F��T��r
��o�Ɨwec�@�#X2����B��p�B��w��^��=Z�&}�Dm�,�*gv���e�'�)[�(��#�{cUE���:^nR��J�u;"De�Oq3���ɬ�
�:�@�f
r��l� �x̶����̮=rg�a����K�̿���&����b�K���B�h�a�.}�^:$=�5+0�\F���8\}Sea��9�WM�#L�c��rJ�eW]�ӳ`%�fҨ���ݺ�ƥ�l�+9�>M��p�8#Lb:tk�`�ɀ�e0.C�o"�o���B�S� G!���.�3�����W�r��ǰ����\����e�v��c�B����6��"��\�ћ��O�ޑ�[L0�G�{蕉����!II���Ƽ�U�0sa3A��h�j
C7Z���0e���lJ3�vgw ��M1�1k2@�3_��r˔�ҝ���+�X�`�d����t�ݓ5�`�0Q�������;a�ygV�=3,Em���T�*����Pˡ{�埱�8�5��
�H��EF��Q��^U�!��䫰i���@��n"��ʕA��]�����!QPD�k?:a�=H���n��B�~�������!����khe�tNA�B�l�*�1Nڹ%)!�n�R)(7I�6�v�i�ʔ�Y����v�;[�nИi� �*v7i즮�sp��Ų�����kKlQK[+iE+e*
�kQikYZ5iD�K�.(,R%��Ym��YT�km�J�,�mmh�XTE�b�h�*VV���h�S��2[�-�X�D���ZT*�R�QQ�Km�--m�*5R��m���	FaUiT�(���e-�VQE�b�X�����U�1�Q)kP��[R�������-�R%��AFЭ�*6��U[V)cU[��qT-j��cDT)m�e��b+���V�5�m�1L���1��(�UEK�EE�Klm�1���ګk�WhŬ�h����J��l��*8K)mB�Ub£j���m����WPm�UR�UE

��jQ���[T��QX�D�TmkKRḥ�Z�"%E��-��V*E��UFV��Um��(�6��DcZ���jḠ�����b��PPm�5,c�������T�5��Q�-b�$�@'�O�/=u��=��W�H�/v�e��+GcY$�1�O�G�||i��)ʘ�n�/�%�}�KF�o4�ѝ���%�Nn��ʧi����F���g���QGi]��st�0�Bu����+�՝{�v.^X�D�8�L����E�F۞,������赹�)�}��#�g^n��8"к�������[�$+A�
�x�m!��`O ��:��pўq�[�wE>*�p����^ z�LPZU#~̠hBt��0͕�:z�wX#�w{�V=��SC�ʖ��˵���*`2geT/�Z���3�!���׆.u �0�ON��K�����tJ����f�7W�N���CzD�@Z���e�R"���l�[֖bQL�/?Zf	Xj�8=���3�1�9�Xu�p@vӏ�"��.������Ԧa(V{iq5��x�Fx\�C
q��lll@�r67���pC��MzQ�5%�ܛ��$�G�VI�>l��x�=>V��p�]L\�>��1�$�V��p��=��w��圷��J���'�yPf
��g#��!���׆�2.
����A�RL;5�wL��IY;b�DɊI;؋LdLEs9D��.U�4�ط��]�3�*4' ��R�
��TD�E��,���{s_�py��WDe���"�5�����B�<
/�v>�r�*�Oc�w?<���!ۋ��;�J�N��B�?I��{�!ו��h)vN(`<�(^�iE��.F*�"�����_u�9�^EI��,펚��(�UW&��@`Mu0ue��k���cΫ9�~U����/���A���=ڳ�sء`���0X�q^\eF�U��.��(��(��j�.�k�4��������uLt֪k�'te@}���ث��W���<7#L�6�6P#��)��p�|��6��v��|����{_.[y����ϝ{j��;�p��82���S�
�V��}�7%��:�KN䶹[,�L���tC���P7�_�C�Jص�
$��Ip���j�؏���VA����˶#\
<f�U���ʠ�.É���R�(Y�
�hGJ��p�-!�ri݅��ķ�y�\n\ۇ�(��R�;T@=�[C�5Pю1+H���;�xx�����.a��m]xr�W��j����Z��gթT೩��Ǌ��I{rƽO�[{�w+Z�cq'Q���rUu��ٓ������Jxנ�+��t+O.�,(RDCQ�nj��ѽ��մ7R{���|uj��Z�G=}��O��6��1E�v֊�3(Z��;e>���x;v%�7�غ �Zͩ�x{���Yέi��:{��_�L,|ĹQOH˼��]j墎�Ls��ֵ�w"���������O�MgG����ѯG^	אG�Υ��ʐ�p�_�	��Z6w\��!,؝����VsS޺�����.�������2\��p���B�˔F�p�����;ы5c��q#s�rL��s��A�r0jH�[��]w����fD�E�������k���k{��r�(ˌ�X�)%϶x�f��H��ܘ�s�bG=��]3�Z
�+w�7�j�Y<X2�fz挡n+�P�0XޒVt��(���
3#���͜ݛ׊����PL<[rd�Qԍ)�͛����dl�ݠE8`�-gR��x�g��XdmF�S�{mv��٨,!���/�1�5������LP��!�Jfv��ۻ�=����_-׼��z�V�Z���p>Ń!����B��ע����ZG,]R"0v��j��IK�f0��V<��'�>Vɬ��Y���댨��+��_@�1��'�����oK�W�\EgH��qP��L�j� �ڛʡ�%a�����"7��F�5����nĖ�68==.�eJ��W{y���m��.���u�ڏM��|�Wy�I�r[KH��Z�̙d�ѓ:6��h�i���⺬���S�K�_q�;��^}�%�����;:�]阺6w�YM�C��dS��;�X����r(\�\QQۋp��6wc�S��
__T-J2P�@�Qo��t/1pP{6 ��"X"a���q#�N�q΋q��m\Hy�h�����r���>�H�3�̾�����ʸ�J��z`#ƺ�:�:�U�ѓ;����)4�h�P����[8�QSر���A�2X|D�@8؎��n"$��QچZy��^�Ф��-W��L��&Yx�x�V7v$��QC|����Ȗhbz"-��{�vMx�x�H;N���i���U��e߮GDmŅbz��~p�h�� \B�24)D2�"$[ݼz��NC�׭W�a���gg�����gAe�$�U,ʟVӾ�<�Y�n��ً	��P:�ٗ��df܊Q��>,��
X(���"��nUc����r��4_�K[x=Y��r�r�J�w���ԣ���A�70����̝0K��1a������_��Ȋ�b�΀�z��-`����98�a��L�ܚb��G1�_����� +[�c���m&���Z��:$���`pK�m������P�3|��Zy�tٛ�z�U��M��Q���nS���&���ZQ�V�!8���ވ��ju�!Hq�T�<��ʅ
pnwp�n���q�`��!�)�_VW�u�A����Ɋ��gk5;�85�DPP���b`�>f��>͇^�æ�i�e����l�t��j���t<�,�@tYu����S�9�t�\�8��x2�:j2x��h�X���L�s��5���V�ӓ��E�^����a5�3��[�G}�{b��#;3~�>(��^b����f�ct��mE�"�0xحT�/��w�\]J��V~���ձm#�� ������k	�â�>8":ш�O�V�;��W�R���Qǁ�,��}lQ��N��5��m��kK��������훘*8��@�r�3(���eq��@w�vf�����3���wG�ǲU��9����D��6ax-*��fP4!:Gc�pժ�JmA�/�[�[Ӻ��I)�R�:�"�:�ꃴ�y�.�3~��1H��	�dCu�Dk��}�7ǆcKs�3;LߜQ
�z��R�;��̀��E;�j�h�C� 8x"����5M��ߺ��z���+yx*�1���`f�	S���q��tNp��O��l �1�%=Y���c�l��{8e�V�zsi�m���C5P��<���kc��X�?8�;ޑ3�o�'W���{�o��%%W���5N<�xn��}���a�i=ul�<���^���^����rk���ϐ��o��-���]g5Gc��焼�Zy3�ב�k)��c�N?�3<�L�xz�f��Àw�r;�)��_m�Cx���N	�͖xO�����<"71pux<���J���c�!��3ջ��}�F�S��fp�R��!W;/���t>g����|/N�[77I.�Zmj�i��dB�(E%OI����ֈ\l��+�֊�YEx�v���=Ǔ�)S�w;���}V6p���)%��TDRT�����jps�
�Y�x�3����|*Q���]mI}ݴZ=�Kt�W*��x��Lu	��x��ߌ�hf����3��	�ww�����u�gkVn�`z�9/O���w��¡�q��k��P�/��/;�ǟǃ�wZ��X�9���UF��UWv��}[�l����awMc.z�h��
ܣ�
�%(}�-�\��������_r�E�K�8�,��j}������*h�	�xձ<k��ٛv�Uo1����>�Ӄ`{��]��_�8��p{�w�p9@�e��FVF��Vt`�G���j�Nz^-sӂ���5W��{��ݛ�<9Lɛ�H+E+(V�G�(�{���M�o	�{Z��]֎�bu)0��v,����Ff=�v�u��rdN��VK�X�f?��^�28�9�W;�&����������Jjս���e�c�tz�N;�Tޜ�����8�m(��d��<CFgw&�:!�Ie��P�
�qnx��;KZz�0ز�j����<(��\w{e@=�[p�Tó��gD��E��5=�D�ލ��cwq�dX���&�����H�E3��&����`��?�^u�UrkƦ��e)��u�R0�� � ZH��9X x�S+�>0�֫G�Þ�p'Rs�n���Ng^'S;��Y��6���=�~p:�z?��#��R�L�HK�\-�p�_��u
f$^⳪ޮ��:tE{]�"�:����"�WLɯF��l>��2EJ��@y�;�9���k�jY��Mz5�'ր\^j�uu:��R���/9r-%�m��뮨s�=r�{p�cHY�����H�LѢ�8�%
�\�
�ʙ$Z��1�	�wK�e)�zy���	���E��ٺr7o�B�P�P�Y�Ǝ�Vt��9��@�F�����}��[y���d�9rhr;AߔN��
�ClePdVmR�1��[G�f)�jMԨ�,�������SO~�/A�m֠��5���d����Z1�=�^d:�Fbs�k�Y;�x��QBs:gq0�Ǖ�u��)w�8��9��g^�f�˧-[{�f��JƩɳ.髼o���0-�8`��U@1��ԝG׹�;�NNP��4�_��5�^��f�͍�x/'[؁US��[�t�LP�����}B�L�������w�p���������b����"�趖Q�d¼�)+ޞ��f��繩N�8����3��ʵ��˽�jF��<}rVG��D�뎣&1�#�1�x=�s�u���6�	��D*�K."�Ȳ�b�*�)�eK���i�r����u2<���ϳ}�:��,���1��q�
#��k�h��ts��4p���ϕGNm�خ�(��^�b��re��iV�p�`B���!�; �W��[�p�w��fWޱ!]L��WN$�,�/�猱��V��,c�q&�B7Q�u���f=l��x��7&���H��x�<�6��Qt�\J�]3&�,�Ҵ�H�h�>�0���ּ���������9���9��ȡ�]�7�n��DjdK41�qۮ5�/Gl�٩��)P��bԮ��!L�plٺs�(u;f�3Z"�K"�R̩1!v/x���p_`�y��.wpꝗIMe��1�8�ߋK.| �iM*%/k��%i�ɍf�,P��O}�&�Mܨ�Z��<Z���={k�p���-�2ӭ3�f������vL�|�l�O>{2������nL����݄�\���P +��n3�/<]�/
��9�R��6I`On�wQ��|�X�ޫ�Cv��05����y*��ا#&�m�C7(Z�a�1�C|��p&;�o\�'�0+��ܭ��>;M���N�#�W.����͜�Bc��opk�[�:��>�jע`��"+�Õ����<�&��N�:�v���c)�3H��^�����y�b7:Q�p��Yy�hN���DZ�8r�Ʊ0r��PdFl;�ӆ^�yQ�c�������yY������BsiI㥡���������865<xQ��xB,�T���焴���"����el�-`�[�O:��eÛ!��gq�<�85��㹕�yA����r��ۘ���T�d�'��, FȧL7�R�+w��z%"]Y� �Zw�.�we����j3E�eW��8f�8���"}HH�0;qR��b�W�A8��8��׽����;��g��pr;�r�i
u
8�0��N�ѓ(�$V��uI0o�#N��k�%P��9z�:���d�n\4�����Wf��w�50�1�vHGj�y�J.�ۦ���ZvG�Y��q�'+,��,��.�=�Қo��Pv9�����K���V��]����sT��V���u�r��������|�Ya�ƞ�8J(;���u�������C�`�N���,��򳏞T������V���h��O\+��du�uA���y�.�3`GK���!b���wO>'L�*�=KW�R��^����v���Q
#�0q�)��lU�Vy�5"(Y���g���]ԧ���f�Q�}[p��r̋��,爭��8]�UnQ'hB�s
(��w��ۏ3�w.^��g�
���1��Qb���Ȼ�"��g�4��t60[F*R׮�S�Y�S��rڨE�V�~��2�����g��1�ڭ�8�2e;Z�y��������FR�w��d��0׸�rb�����R��Q�k��h�}l������+���K\g�r3�ez���]��($@��IK���D�PP��+��cJ�]=:ܥu�lݰ�Kwҡ�#�
)Ev�{8Yb�Q.�;���r�J}�@mj#�<ڷ]N�5%w
Nsc�����]�[.�1�2o+�^eO*�����l����2Y5F����N�ji#��Ɓ���9�]5�f���*�m���=����O��.�Հ��Sb�[fL)�F��,)C�ѽ�����O+D��96�X���^1mi����IST��X;S��-�r��wM�H����ȴ$�E��y�����+��;�ފ�|�t���zR�#��#��ق.S�l�Y]\���3��YB�d	!Roc�`�ﲉ��W��T�v�lv�^qt���)z_Q������й�!89"V�ܻ>����'��x5�w��^n�RXx`��W���ִ#35��g`u`�w>��[*d�l��nkx�(��������c��9�=� �0�ŀ�Œ����^fC��8�5�>Ւ(1�����)���}s~N�Ġ�+^X�ɼ'|���U�gR��z�㝸�M����}.K�<c<qT����m=.{:H���1������9q��@V��`[=j�ͻ��ϲ��+kc;���X�⬽�p�piy�m�ȍ���b�fu�}6�Oh�%���P�ck$K�����On���'���H��^�^ �I�d������u�v�]v�\�To"]8��;!�G�S:�#�2-V𕹛x�@j�MQ\.^5:��6�E�Rd]�ӎ�H�C�u�C�.��@�� �͓J.�:�B8K��PuV%4.�N`��H���[��"տb�V\pW�����X�i}�>��\97���Mt4(i�F�&��0�X�h���W��my�ц*d�3+�|Q�c���|-�Y\�p�hȡŴ����K��nێ�S�d,��jp�62wxf�ũҍ��76��ɜ���ׄQ9���#��N�9
Bd뛡o7�;B')[ݥO�@��V������73n){���A���a����tw����4�Av;���f�/P�.}*q=Y7��J�T�]3�>�>���1Fܕ�"ً��"��Jh����m����]J��t�t�z�l�o6�o�p�Jӫ����1�C�{�`3_E�W_rz:��D�fu�3!�
aݹ��#]u8=3�w�һ���J���t(A�xn
\q�N�0�7�ˮ�㫵�1a�%k>�.�c�u�������I��_7Epy�{���md��.Q����?+2<���F��τLg�}�pXs�����r׏��9<�}s� z��S�ĸ�	��(3�9KNf!�)�;�������w��p����=��Nymj�
�Prgj�F����[�m�g�38���g��Lu�S�Ò����X�',BYeJy�j��i������xb��5��V�� ����Ѻ��)!��ӟa�o�Ͳ	�S�ʲ�w%�̰���0,(<����`
;������:�OqY.YPE2Phn�ds�i�Qaf��K���ef�Rm+Z�t0�aP��бJʨ�*,R��U�KP��-����+6T�e(����mQAml�T��ŗF����-�B� ��
�DER�KKiZ�[(�P�Z�2������(�0�bU�RڪZ��E�Ƶkb��-lQ�Ҋ��K[Pam��Z�*�֠�FՊV�ZĬ(��YZ������1J�DDbĶ��hՌDm���Dk������"1DZ�DX"E�QF"FX����m�jZ�8��Q"�F",qe0ؤT������5V�F"���EYm(�ֶ�D1PU�eF�H��Q�Ũ���.E������QEbJآ�b(�)Z�"(���*�,b����QekU1%��KIZ�Z�b[-�b�*����R,�`)PQ�
/�RҤu	�3�ۘ�n�B�p�v�^Ӈ(��+-ϫ���-���!@���r�*��oKΤ�Cd���z��D�}��I#`ɔ���X��9����Y`�F۔{6x�Se��f!ۯjD�	���S�[�}&�>��3��3]E�P�-���;lP�W>�Lđ��,w�6�y�slm�.�,U
�j��Z�N8g�[U쫥xt��f�,KUgs�(�bx�.��c�]�H��-1�*}g�N��O)mK �8�eH�����UgE���f#�n��Q��,[���e�*���
B�<U����h�*b�e�9Nw�l�n*�xE����K��pD��~e�(���"�c��ڤ�/7�H�
Q��R]�έ����̇w��1�;F��#��_[����ރ��|��Wt#g'Q�R��)�]J7
�Ac�5jC1>x�����{�lMF��Z'���"�eYJ0��DJ����7������X�`n�j-�4-]#5.�,�B6")*Cp����J������ׯ�w7ݑ#v1�Z�3�S�N�jD�R̖�l�Su�H�pN���n�H)w�.NĆ��e��1lY3�p(���J�M�x��&^A�q��^���9�Գ\w���S�w�1��K�N�2���f�J�P����]�կ�ל�D�X�eա�G�D,����w*pz�	M#��Iه8�vk��pԎgQR�K�����k�b��p��N\3��s��A�N��a@�1 s�1J�S0A�W�ҕt�Rs����{�Ν5.}YL�,ʌ�])%�q`�K$�h�Ɍ�T�(H�F�ؗj��Xw���K93=�9NFUȮ/�c>�8�`�~VK�TOT�n��x��CX��8bye����qpa^N����T��.-��q�SGz��75˅c]eě�'\G3�@]_B�|1�G:�y�`�b}�k��E�b�|�F���BY�)�8���`��ƬBq��cD�]\r��M7N6��m�.���5���,t d^�$�G8Q�9��2�g��sֶ�ІE\v���l�ƒYS�k��WP�tѶ#�ۖV�.#��"ʰ���'�,�W�#�Sn���TE�e1�k55��s��Ɵ@ؘ܊�'M]u8�Yg��6lt"�mqF��*�fc�Z�̽�r���f���W��< Tr���e̍��؎7�s�/\���<���$-�J󬉚IУP�\�;u��͇N.��Ш�Y��ӫ%g62{,�\ޛ��"�O���:9;�*Wu�1XK�M����0%�V^k�X������\v�Tb�ӏ4��yk��*��֋��&6b�\�6_m�5u&xs{��Ϛ��m�{�<al�g ,��	�<#:���h��%�ŵww��v�QY���,vd����Rr�%g���R�u�C'�E�
`��{f��\홗��%���g��Lm�X(�s�c���	:��Nè��ȶ'b�X[�U�~qo�wKO����3L�W�#n/.`��p�`�PȀt:�0kVybU)�������َ��^'�w�a���9�������6|,�e`*Y�^f���Q�YR͵�����0���O��\�ZC�]��R������X(�ʄ#����E�#�_lζ�k��ѧ:�r��p�|g�"�Qs%��p��p�7J95�w��ʠ��$ӳ����E�'�5��ۗ���"G&*�"+��5��� ���vpf^�̈3Z���q�^o�_�7��E�^U���8tyؽubo�3��p��2��!
�}iWG붮��C_��Nu�ܫM�*x�l�ō�,�]]�V,b��8s��� q�Fe9�
��G��G0u�.6��c"���ޡ,0����3���t����FW��R]�WqGk��X�U�����q3����Z�\���Y<�9���-Y���RJ�����TI�Lx�6!W��t�p�x���q�O5�[ˀ����l��7��Y���E�14����Fl����2�=8G<�V�~�����<�x1���Q��7�m�|g��o�	��R풐���P�~]CN��q����p�B��}�z���"��Z85�]s�̎�7P�M��5� h�g�|��V9�I\����oʧj��nO$��c�oҥ��#25�F�n�B9"�Bu�(�\�_
�x��P�;gg�!�5���NKU�\`4!�l9�"��6b��U#r̠Jr�X��ޡ��L�O� M�{�ta��Ig��6&��Q鏶=��0Z��7!��50ea4(���m<���j���%\0�Tyhs����v%����z�Yi;�XR7B&T�=���5��ݭK����P���]YTY��5s��:���]�|.ִ�ý�G|���x�M��6ށXu����B����FQ[:.W�
���a�Mw��ne7<��}0:5�8��U��N0��se�Ơ���+z�Jj�)��q08�xe���ӔIIqⷵ*{�{�՘;�~��сr������{�[/�x����	��ѫNwK�:u��Z`eR��t�A��nd /�X���aW����t3G���ٽÚ�$�5��șz��R#%Z���c��y�P�P��h���8�w��/_l��#y����z�\ą^)�m�1A����2xD��C=��fg"� ���f�����^ru�w0=館�<��f4������-���������jf�t������m�=�ڸ,}�<p�R�q~�.�p�Ņ$��WdBs��{��W�!�\��������v���"�p�$�S+Τ-�x�(m�����W�}�#/���&��7��Y�H��ߩ�ց]��X�޷
!V��߮�V̠}n:3g��UtUGv��9�;Zu�5�i�8pז�#r2ⷝ#;c��@��}��X��Z �w9l�-��������Ll@���qf��ޜp����Q���V�)fR�82�..��{�6��8&��c���E��$ud�1Yڋi鞷��������!HR68�tv�CH�Q��3K�g�+V�׻ˡ��Μ6�p�;vE�5��d2yN+�>٧
���-7%��X����ii��P4!���sҧ��v\��e5�����h�o�p����֩r�V��J�N��7N槲��Uӑ��.�u�a�Zך7���T��y����>�����|�
�|������'��5rMM�����u�%-�x�!��+�w�X&�[�PcĘ�]7}(�W�E�S���W���}��o�y�䦷8����=y�N�R�(��(i�Q;��+�x�.82��阦�Ug��m�٭b�vw"=�X%E���Վ��H{P
41	'��Y���h^۴Dڴ��iwዣ�]�r�L-Q�3}����A9��w}Q�������N��9���ʈ�k�3�D��[�A�sO(!�����v9��lE�d&�
ąR̜�R6X:]�*��7����iv�!�ٹ�fٝ���KqC��TņR.W���֢�Euv��/p3�7�����S��Z,b���o�x>3r��="8�PP� ����V'��в{&�_�>. }Zh�+�A���+�\
QWP�`8d�]$����;A.����w�Gq�Fs]�.H�s;\^	�Y��V�l@dh��JB�{\/%�X��@�
6���hVW{e���؃7���lo�-�)<�,N��U=�h���S�԰ ��F�Y3C�[�P�0�Z�z3ں��fϫ=�����kI���G��M�6��6�����C�ے�]A�{SKGc����1�$�/SG/�]X6��f��Ҡ��h*�A�#v�9�1؁!O%X�&"�\ʊGy��!�f�q��f��R}�A�W(�h��##��+8��r�[S37���]F�����Xw n.WWr���]��(ج΢�li~�t��6&@�ґ�Ȏz�n.�o���s�Z�ou��"�ZwK�@ݎ�ʋ��)����2�q�(�S�T��m�j·q�&�y|�^�g.�8�]�U])x:�ǂ��r:����xJY��,�УJ��f��N�U��֗%zt�����DH	gk��*9P�@���m3�X��/i�!�1��>x ��<u�>���]q���q�]PY��AQ�z ����?-�5ө^�z������ԖPN��Lj��:$[(\���%�lѷ�f|�Κ�e���"r:�F�T�Ap�jWi^C3�P���^9±Ƞ1��&��h��!Lh	�,����vb9]�bi�Cr";'���vkLaZ <���Tat��g��kԥ� �z����[��]B+6%����i>�k�~VX�J��wG8c6��cv�|���V��c)1�ib�4P�kʥLR�T)���%Ҟ��dн�E���A�q�1��^m�	��W1ISݽ��iRĒ�s9�οS*�E����R2�^��6����Q����|v� 
q���v��C*ž�������˛�=�[�Hwr�.�T��Ol���=$m�,�u�-�;HIm��jmə��)�G��%��Mg`���|wO��3wE�����h��̫p:��)8{No-�2���*����1R�!FL�F�7�~'a�T�Nz_�.��
[�ֺ��[�����Ĺ��&��~�,� ����o]"��u�ܧPѽ��BM�^��cca���M󔻼���82��B���y�^���}5�Bx��*㟦t��Zra��7kK$�6\��^�t�1���s���Ѻ��uuX��\�aO���������[[A�/����z���1)(؊�vp�$��s;{5�=�r�.W/'ާ,�^�)�
�#)�M�q�Yx��۾P���a�k{�+�ti��"�����K���0t͈��:B}%3c�MnJ�������7�=pB���f���s�����ס����)v����S�5��C���q%u����N͹"�!��C���Y��B��2b���f;�E�}ˡMX��m�D���0�<,?���cG#���=�G�f���e�n:`�f�<a�Vv)nF��4�+�;��v<�Z@o��D�I��`R�TsH*�{�C��m�� 
�g����G�ȵ0K�Ֆk�n�3	�� /(��ݣX�v7���eu���E	oE0hCt��iC*�l�~����jGZ�"}k��S��JHW4˒r���XRf����+F����WB�N�4׻fV$�yx:��xJ�S	㥍��ЖF���R�P7"N��M
�ꏂ�U9����Z�ny��̡Ԅ�7z�fۍ�h��V&(*n.f��S�3A��3JL�4:]���rSU	�#ݠ��W�#��R��~��u���L@�R	��(+)փm��1J�0eQ�k��h�rkl���e��T�\t�_�\�-`�}�-`Ӽ�'���&X�$��.bŨxa������Lg�����wS}������?(`�E)�;&���,�jIs�����=��{��)N���' ${��܏����@����x�"J�ʜ����mʶG��:�\G+�������#�NFz�xӹ~!h��y�����Q
��\>�]B��=C�T���{��*�d��4�7Xz�p�sdZ�̋�θ���o�CT�+N��b��*Z�y��ny����ߛ#T5~����C�eݮ�R}N��D�����=�Q'�n�t\8[$X��	N)����v��,�V�`�9j�X��g1 �*jq%tU�?����˭湬����w�Y�9]u̗b����/��BRw�eb[��p����t�fg��8�6�W��Ua���(�-U�y�t\�kw2�8�N�\m�\Qc8N��$����V@v��zg��8#��8[��P�Uˠ���"�w�p��Gkj��C�Yў�ㆅ�F�ʈ[�;�U��F��-�
�K�Q\�'͈�YU������m~=��g�*�W�PW��_�E�)��l��=�غ����4�ueNm��Ӊ.K2=�6a0zzb���
��p�����'aLoA�~>�h=�v�>j�iV�)���}W�PXX�3��ѕ��� �l�"�g��D��8�̸JZt��\>��Z�qq`�SR�a�.�p,&���:�B��2��!�I��}�&�3��j����Zz��H��d�s��t:"�K"�N����
���S2����Ԛ�2�cf+��~�H����8Y�h��]��3�7ʘ��y9�Ġ�ˢ�k-;�tt�F�M�{�㦄��VJ9�E�Q~�Z�^��Oޒ�/2b�W�<.yT
�U�ь!�K�9��,�z��+�T�
��	R�@�h2u�5�:�T�ζ	�9�;u����Z���N�ec^��,c;��o7eV��ϥJ�P�Y%w�H�k4^H�o�C�:�X]ZGd�Ve!�e9��zl(�-Ԅ�m�1��ig�s�0N�;y���y����=H�n�\�w�d�\2�O*Gݓ�d�K�ø�b&����|�֜98��S�ʃ\8�KaVCOUg��u�*��E������a���E�����KlJQ,��V�}��uR��_65[��P](^�p���[��=U.��欻b�>5��\��/A�����b�,>�؂ ��e�S	���5�����ْ%��F���ypm�v1X��0���\�LH3��Ψ�1@M�1.���ڲBy�^a"ݶ����:�����8:�ӈT6�!Q;�.�,Dr���"r�Vq])@��F,���R�.�Y��+�K9s�����+�F��>�k�sR܋B�}N���ob���B��r�#��N�h��Z�g]2�.�VV�v�;P�wmq�����aV��e�i'9n[�I12.. �J
zs��Rj�X�z�.�!P����,B2|U�xٖ�q�g�n�7��s���h��Fۡ"�˓q�<��a�S�Dp��(!�Lɒ������,l�͒��ST!�����'��=����6��O&Ut�y��}��o��Cf�!c�y/�x�?{�f�����2�(�<Ge+6a'�X��W�r�G��=&�yMՌ�)���u�!V����N��v�r6���Xڵ&8i�iXքX�ܣJ]R!��z��H�.��u��0+N9d�ל����S��ҧ��;��05��]������y������A��k��Ya`C,�@ �}#Ǫ�p�\޹kGx��3-���1������% ��8�VQ�ݺ��j�������Wf��.��uCp[G�g��Me�*叮���FT��(CW�p�9/!~��ܨ���6��$s��^�xR��2�U�ԓk	P�+��e��ѥc<_f��L��1"�$�m�f5d8�o5�*`�yQ�5>Yݐ�=��S�eU�ԡfN�Q�z��
�S���5���N�`�F�7���L1��c�
2Ȧ�U�E:v
wF��u�g5�hN��S#5���e
����[xN�ƨ�yv����zHV�J`cT3q�F�AE��/��V�����6K�v�7b��v����7�2uV$�x��N�,nx3f�\�����:��jVf�{pkYo�w��78��*�-�"�(����h�+jQk`�,F���R�PUU"#+QB�QkTX�+X�l����E�+���������6�VEkA��X�V(�Fe*b�UX�X��Ŋ�QcE��"��VQYV�cҠ�l,T�B�V,`�"�)Y+a(��dUX�"�V!R�ʬF�����FB�Kh(�E�UV-�!�V(�d+(�Qb�� �F*��Ҡ��.)��U�m����,R[V"",Db���T�ʬ�X���Ա
��X���ibȖ�R�Q��ʅJa�DEEDETQ	YKZ�V�
�V,bV�-�[��RUZ֖-E*Pcl��UDTEkm���V�h"��0ʸJ���m��T��X�+*(��%*ʋEX���mXŭ�E�k,Fڂ(��ijU�@cB�
�	U����mU���%D-Z�>�ٓ�m�\f��:���+g��^��;���c^�����$zTl���$0tA/��yDA�9�}��ɽ�涌��o7!���`
��7|��=�Rke����9�e��}Q��x���l)*R�nC(��z1{��젬߫����*�<� ���)�o�= ���n��TT^l��2�Y�u��X&�F;���T����DQ�e)�#,���?Cb	Y���<Xu� �������1���,��|,_�E�.+h[��\i�s�1*�W����Aݷp��r�N2��):��h�u\hչ�V�^��424�b��]�-�d/cUR^�Sݘ�
���Y��Ht�d6�����u-�������HwR�*;)���O��S����w�n�i���B�Qe�S�Sb�T:ģCfj)à_K�Fƹg3Dn����Lv�]z��t�x▭T5�rK=\��4�;ή�'�UcZ�	�����V�9JuJ�x�����R/�} 7�h�S�Z=�Ɣ΂��f5R$�B7o�4/[�\��l��_{'u��-u~k&��,��5pF�h\�p�)p.����g^��:�숪�d��+A�2�]4O?�P����w7Z�ȇy�"F�1Gown�j�@��b����b�X�e���w�L�ta��=�*U8�i�R�m,�����:��\���$<��L����.���~�ƙ�]X�yFG�q7�L�ъ{�	��:B�2b˓v^pGp�8Zpu	Ԛ�I�g��r��y�`���9@`�Z�Ɵ�tO���Ƽ9Ĵz��L,r-��&���0vU�]Vw2�n��+��u%'���B�k�����6�N���ֈދ�M-��_3��7����R"F�4��q>�5�x�T���j��<,7��8q�W�n��+���U��uǁ .k�>a:u�y��^ϒ㩿*��������oZ�U�xWrݛ���gt���
5�N��b�Ɖe�!NT�lJ�vG� �۝k=�oL5���qv�%Y�V(�PF�f� Z��L�l�����r�X!C^�B�4���sqJ�+x^��l�)��e�J���4�X����)�Չ�$�,(Æٙ�Dx�YY��fE�m�+_��9�t�|<*���V&���W���1X�ޫ���9�׉#�7�t����;�ov�qg�մ�*�DSG�Lk���� ^�,ީeź��(�	�$��
e�B�w<V�]��KT�����L�D�@�}v$��`�FH�H;��:��[�S���� b,:G����p�ժ�FoF~�����h��÷��?�汔պ�%H�pq��nor���6��o��i�y3~�KUr�z��{w0�=zS��b)��,��%���w�i��#~ƫ�/-M�t������|h+ہ��s��6���m����=>��q�e�}(�R7c��j\�F��_�:GD'v�9�YU����J���#L$da�l��sˌ�_)e�:C�*Oߏg���zZ�\ ���������_�:Gs�(�2���<T��GTgv�Ao<ی�P����e&�a�v�c�O�`��Hi��wН#�T|�N>5A]*��pE��v�X�.O)���p��U��Vk��w�Q�"�8f��4V����l�I��/U5`�`��(����wȮ��Bs�f�U<>5�(Au���5�a�B��S�hÊ+��-W����8k��ѓi�<�3�f��-�"�]�4�#��)���w�P�X�0xň�̨T���{�\B�Ӥlu�Z�& o�����,U�'Z�ᘥA�*L2��H�txk<K��Wy�-�^�|�;����[[�2�<�&X�
	��u�D\L@=��EH6N�	&�]*]H�@Q9o7qt;m��l�.v�l�	JwZJt�ٞ��r#7e���f: Ȍ��j1�P7h�b����M��<��?��~�K�����k��\�����{v�%�*9�k����eGy{9�,������T��|8d�f}�m*��8͖��ѱ��|����jWHd�)Cr���	��}��i,0FD��	������x�'�+�u������[1��)�);��V�w�K�ѝT�ҷs��m��ů���n��f
�iu
�N�>�/J|�p��g�)��XOk����r!Q���+ކ@����-~!
��cUn;�0vmgGD�^Ft��j$��C�Q㢺��B{]�e�<-��UҼ:y���I�&zFy��ztzR��8���W �e��+����r��!�N� i�nѸ�]р�q��݃{���-�g��R�.�󃨞eO.yq=1TԻ8�1]�[�x�t7^�6a�I�8�kȿ����..��W�0?8s�uH�ӤYFH�
�9{��f����[���m:G��s��zx�."�q�p#}
{Xb����.mC1�Ъ,�(�Wq��v�*3m�w��z�mAk3�-��(@f7�jF�	$O�q�b�h�#���A�K==zhA�ד�.W.���Gè�r�>�q���s.om��V�+�)�;�cS�`�a���f�G\w����M���q9�*�G���::�������1(B皫�w�rΧr�F�W�=]��M��8[��{;G�����[�;�h۶x�9�N�Km)wk��w*zY�gR�p,cW}P��C��bC�Af}hJ�Rk�����2��L�y��*˞�T���#\c
���0
t:"��YwzW/aU:?G�X���4��Ǟ�����q�B��4)��@y���Rb�"�FQR`کCZͭ��݂ }Y�e�K�=Ja�5�����]�X�|e�Cϼ�0�V�jYU�V��t�u֪���<ʜ$��*Lg�K)��+��-^���oʭEO�ٌ��ě��[��E[+��jy�:p5$��`��F4dY��D��{�hߐ����3�ŧ�M���i���������h�P����.�Nbu���0ᱞ@]_F�b�|��yk�ס�Rf���QZ�ʇ��GNJ4f�`ᢙު^��Y�s�prd������i����9�EG-����#���[KQ�F�T�hNm2M�)���>x;#���Od�6����[�x��GѧY�<�J��*Yk��l�=L9Դ?���t���^j�:}�G9��V9:Ej�}�b�{Xf�"&e̱��wI�f%�e+܎?�*��Zޤk�^1:3���Բ;�pd��ґ�XGJ�пN�8Ojc��.�f��Fh��:cN���v�}�a��pS��vdjq�4ff��\o�H{�;&q>�1�ޡZ=቞��NX$7[
n�p�qV�)�����tr���������8�4�U�Yy��jy.X��N��pl'�h(����<5��)��R��/�<|I�3+�MyN�1�-��������$K�ҏCU��:f���z�
�Ez9P�l�7 S�����/�w�]G_^"�Wf��+�Ȏ,78�Ʃf�>�>��[8��c���S�3 �8#�q'U�����w��v��k�����kg��*�Y�k ��P��N]�,�4��etL��pf�qu[/�f'Z{qQ��I�B�h�C*�Odm��^t�nGn�I��U��XW��gV���֗!���0��T��a2���B�[8M���v��)N�~
��31��"��������������8-,G�q�@2K����>��='�;���bA��������ξ�ay��Ǘb�����i��jcA�3��U,ʓ4+:�'iOL�8�$��`�uvI��}���Ԏ�~�&�_���kН`-��3ZC�]%�}���;D�j-wx�ox�Z4v�jt������Pf�� �\��E8Ȇ�Y��k�`�/ 3�V���]����1��G�D%c�����u��wn��u�rv֙IgS�V�δ�Or��,��r���Z��(��g�{|r^�(����K��c�i�Lut;w��Ls��eqל,�s��7=Qu�N �Y��4�i�ѝ@�C��I�D_�aÕ�̻Z	����Bh0ux})�������P�o�����7�S��DD���ֽ�5='8q�V��}��Z~��`b����c<2�:Y`��.4�<gr�L']�67��!�%|{��i@cu��n���=FT�`jb�+�8���#$'���\ɛ+�z�N��yc���ץV����V����٭<��F��X"���Y�q�6�`s���(�FP��Q�O�qf�b�sН��Fe�tabx���6��Cz����^���x9�9B�H������B*ܾ0{Ҋ��"y��:`�r0�h�V�݀s3=���r�tO=���JF�~��W����{6�U���8g��������dʕPנ6��w��	���NK��b��,�Z�g�EV�1��ŵ֕���m+0_�u�P̱YdHzD�B�0+�ڽ�.,�����S�y�}��]F'Z�WS�L:����Z=|b��:��^��Q�փD<�45�9�B�Q��N���[���\��w�����3H\F�|�|�A���¹�K����ʓ]��%�(���ݓH��a��MM��q�ڌ��[�S�w�7������݇q�q��x��fq�w&1��L:Ώ�%��zr*O�=WL�ɭ��^d��]K86���>\�׾g��,6(���M�%��:3�E+�f�UQP�"�1,�qK�~�}��1�5��qK41��q�l�:�lEu1A_�'|}�V�^4�A}�O �!��f��d8Р��^���o����c�l�AA"1A+N�u;�yS�SZ�~s���+��,c>p��a?)�m�=�x�q׃^\�� �vz7�7�}��I�X�{���\)]�,f�_㡷"	�?�,����ހ#�^ME������ͿRT�'�8[�ˋ�$ű�؃)��ˉ/�=t�T˩�JXN�AX'�rS�+qh!�ۍ�l��¬.�"�0�z�K�y�wy�y��8�>���/^m���Wf^B,PDp"n1��P���E���ߜ3{�׶����u�h��<�ֳ�X��s0��ſ7��=KC�I�TF�ix�T+v��:ZS~�uvV��g�k@���0�B�I����{	$�9�r;C���d��\,0V����}���j��mљH���.{�}=�1�0�K��A�힜x��ʾg:Λ����^�@V���3:D��,�3�2�Eؗ��\0cZ�%�Bf��d{�Х½��T�-ž�掋(�lJ5t�D"$��ԫ��(���L�}146$�=n�,y�n�dʮ�t��i�z:zb�e��(�QҺ4T�[�F(��l��lI�s�T;�[���TO�d3��8�J�/hU���Фw��7D��S]"�/��̘�p���kkR�Գ�un�F���Vu3�-�6ef7�jF�	$In;K�Qzڄ�œ���YŎ�y���Hf�nݳ�:n\�Ȱ�き�mG �՚�3A� ���O&IQ�sH����JES���g'H\�k��~<ML^�Wy=)�"Swx
R�$\ekg�3s
j�od�!���:C	��(��pXЪx,��l��9�R�=�se�H��ô�]%}bA~�rL*�1��S6!	��Mh6q������������ʤ��5Ư��^�����Segן����+�=4�'%�O�MS�ts9cS�ouOvZo�WFG\0p��A�.s����r"�2,�tLH��~R^���g�Xw�S�eZfT&�E��.x0cpQ�p�-�!v��:���,q����2���%Nu�Z9YS�Mi��M0U��/�`�>�XU�{a-�&�9��f��A�/g�FI8К�(;Q���|��3�@{+�V��W��I�v뵎�N�9Ӕ�cj�"�.��6�#:�ě��MЂ�����f��*S�w[��L�l��/yA�%�|��ݚ[��ߓ���E3�-��Ul-u��]\r��*_j�:�Uޡk���ƣPfҮ9Y�4hZt��K��,�Y��#p���d�9ں�u�,���x�T�bn�Y:&"-�|*ik�a�m�bu_O/P��K."��YL���|':�ǹ=׋�9�;��7��g���l�ȳ����nc�(ZƭK�Fv�)�ĸoV*��k���g��<]��⊇յ��j�]ʰ&O��C���ぎ��7��x�ޜ�]f�_���/��e>�>��+g��/W�.�P͙����UI!�飆b��c�����p��B7P����
c��k��g��#^�i>����<��k�n�m&�p��TvV�j��/a�0K�7v:Q�:a�z�bw��{��ؓ{�V;�=;���V�>�W�C�(."Y�bz"�6��kA����8U�y�fTic��
����`X���k���ɊH������_X�ƣ��N�]0����"�<�9��{B���Kb`��}E�8�vZ}m�jba���U��n���C��%��d�m�����q�
7��M��t�Ȃ�\S��_$}I$'^�Ǒ�-38]��t�{�/\�۾7�p%�ݓyt�[}ꦯv��B�l�Γ�1k����:�&�|�4�k�,�ĝH��v���롻"�NN4�im-���ܸ�-�c��/(��gM�B#���=��e����Q�'�UwY�y���:1��՚띷 �2�=��o�y�D2�\��]&�*�'�Z[2�6��/�&s�\̟u^��.������<�M�
��\d����ۅ��p��n���ɻ��K����A>��S�Uѧʝ������t_u>��þ~F�\�Fudݻ�js'�����"N�ͮ��P�d���}8�am� ��v�O��:n�n�mB��*�{H�+\�rX��,?wR�p�=��XXcd���ֲ�!Yy!��ΒY%V>�\)��ߌ%��Q�]��b�b+1j?S{f�[<:ms*�q�Hmp���4Њ�~��n��d|�8p�{M먻\a=S9,w���/�
��%���u8:M��>Zt�Vu�Cٻ��3�ǈ��Q�9ͽI��{>cG�Ǫ�o�+V�{�qJ{r���!M �5ܘ;T�T4:��-�S�Zyf�;\� $T�C���8�+���a����EYKF��?k1I�b�P-o�O��{���電I���Җ(����1[ov%����3ո��n��/F��-������{O�L�.��������+���7n������Af)��L���7��	FiRl沘��w�&���U�o2þ�+d�n��Q5�y�NH�)R���J��
�8��HA�P;�Ypuݨ ��2q�KY�jr!�@$�]XE����EU�]�be�(������WD��KI���w*؇Z9����V����*�i�I�֞_`ַ�Wiβ�v�k3E}�e��yso�Ѽp$h�%˶Ɩ��j�=F��X���+�.�@�]%M��O�
7�k�刎2�.�pل��x��U��G����/rt|�}�.�4��F�������i��u76���(1�⑍z���*ꋪ��ܸ,�Q���LW�g-���yv��;�&V��F>x�0��{�����'B�V@��������Q�ώ����������e�=�+��3uQ�G����/��j�E���d.U�f꣗8�z�������v{��\^��g���-N�(�wB��v���WlR)7�F4�jhڼ�}l�2]�u����hs���L��iyKkM<�v:fa�}�:�l��x�,����L�.�Y݄���|��4�nʋE�����i�ښ8QZU:��*�t�%@�����~�.����TYUW��ň�D�l�����F1D�DZ�AթEF,��eKePQ-��mkc"�+EAT��(��"��E�UTA,mmQF������TQ���
����QQ�P�AAT�2�ڈ��X�DU�jX�b
1b1F )Qk���-Z,Yqf@Rک��EUU��T+*1DFTѭA�T*�X�+�Q���A��#+Q-���e0ʊ��"#�Q+*1ZZTU"���H���*�(�X�Z�E�
�� "����b�,cX�`�,+
8J�(�d��*���Q��EQ�����h��i[lX4m�P�*��Ŷ����B⍣�T[hVk-��Q�J5��K�,��jڸl��Ơ��B���Z��`�kB�QYF~�q�Fnu��iю�拉{��Q�N�*�Z;�G��B�KG7��[� ��X��Į;�q��}}�,���fv�.U�~�)I"�Ą��x�q>
jVy�X�b�<(e�@��a�Q�ؚ��6��'���S-�$�<3��U,�Fh+j�t�������ɦ���s1Z���:�#�V���9^j�5D5�ElX�3�T���F�:�Z1fb�#� ��V�y��s�N���R�qS�%M8�!�&!�BW���w����XE�;
���BH�N��Ň<���������5�}n׷=pnU0o�C �\��I�D���>&y�#������Z����E{�������h���	r?x�V�=N� �~��J�x1�
��ǭ�
�vny���Y��a����\�Z�d^.���#&$Su�&;�,�e��kSw�$�;�]d�z���!֩�l��{e�kt��l��+�h�C�PT�잶�5(�l��؇Ћ��.��im��3��lU3(�7Qq��1ưEOF�Z�0�z�}Ԝ��H�@�`uc�X��x"�<T�P7a&��0��mN]< ���Z6�^O:������Rn������k��m	�[V(�خ��x�i����k��oX!XQk�U�.�R�=*g�s��i-� sw�s#���J�sՕ|��\��3Y��ḅȱ*'��>}��C�%+��NճDT��G"��騼��֭�Y�.�*�	h�H�	v�6�謩Ec�b�{�ͩ���"Fuk�'u����'�:�X�g��錫��,9��9g�k�Y�U����Xi�k
����5&/wN-���@f�t�� ��
�b�4'H�Fs���4��Y
��\a�o��]-Sو�iGu�F͘,%.��5B7ŔC��!g����o�Dd9�w⥗KTc�a�D�sۭ.��lqb�_EzT�vU��W1����k��>W��0t�=x����F��F�K��Q�iZ�g�WN6���
�##�7�9��ߓ�2(+�f����J��M��z�1l��\&�\h��&TFתY��Y���[�`N�]LPW�h6ٜ3�p��EI�}�s��k�L�r�`�2�V��X�g�F���Fd\2�ס��k��Q1AL�Pˇ���s��U۹��'l�J�'�u�'��ڂxz�_K3�2)ͨ�vM�p�b��anR�V��{�MN7�L�����.�����R�z�q��D�٨�:�P���sZ,��xw�Y_��Ȍ�<�3�Up�L��&�۞�|���y�-+>���<+E��:�:<a�ڷ%���@���اt.��ŧ����A�������)�otJ\͂t�5�ǪTzy��"��WS�e�W'vY��g�}ֳ�=�гR�K:��z_V�y5a�]˧����</��K�t������f���
��w�eٵU޷
!hz+=Ymì�7�U�����E�L�D��9�˅6[�"�0��ZE���^댳<B`8.�rQ�0��̷;�)�_�x�[8��H���X#T(��T�w��f�([���Ҷz�J�P�v�IvC���l�GR���%Mٔd���t��!#q��"�J���ALT�[&� Nyk����4�������Ty�KugDB6vؔk��D+�Ȳ�R��n�]]���,'���Gdf׸�tڂTB�Fק�0hGJ��rT�n�p�Ao��9�r����i8瑶��:Cc�����xY��!��Z�w��B�������  �� ��Tw��Pe���K��������ٷ�)�����u��+�w�ў@�f�䂌����I^5F�r�?%�W6ᙷ���:lm:��E��VT+SF��FN�]��*o�������q��A��GI�)�H\5�l����ю�b�j���m@;��{ĺ�ϰY�"�T:Պ�|��uc��9*��W(�iU݆I�p��kó8s�7��ki\hDo 9���i5k��$�{L�,^S�v�7~<,R�F�'�4�#p��3���a��y5p�Bʞ�F��g��ɔ�f\�TY�T[�{Sv�mL���l��pB��m'��Ѕ5�"�
·�t��a�=2GN����+�z&�c���%j�)�#ބnA��/"���Qx}��h8]>_N�
C�q�z2��w���gS�=U��#犖Iћ���*ذ�Qjh����r6y�(Z����9:L��,���$1C���Q�dIb�I*s����v"�ȳ45�1<�䲠��v; �:��?��[���S�Z����˪`������ׯС>���`�6,J� >�7"+_hb\��3v���*�Ac��)�����f~3�X�pH���'���,�?k�6���6��gr�qp��� g�oe���F��H��Fl�c8�;\ly��Y2t]Y�d��KW����R��Y��ڐ�<����].���l����KFx��;^&������팔��o�"�	�g���VƦ_�J�T�<5���/�Զ�]�>�ɜtN�f��}܀W����ъY�`(�	[|Q���G i�5u$xc�[F��:���N��v�vy����������iojΚ�i��9V
[�U��r����l�]�n�n둻�@��.�a�V�Cd8�R�;��,b��[-��{�+q.�>ZN��Ɲ�{�����FIrW8A��.�3ɮ�q��C��ڒG�IuM�on�-ć(b��lJ��8�1�7������l�e?�3C��C"+U1�ݜ'�z�tf���9d��GhC�j]����n/\��Ym�c*-<��D�z鲹hy�h����
��=�h:'�E�Ap��W1��#��~S_/e$ev�r��燉NZ���'iJ���rD��K5�K���^5(���,e.Ї��H����v�u�l椣x��f�#Z"T2 ��'�	ץ�='�|�¼`w���GB���ng�V�;k�� b8��0c6R�I�q�8I�7uh"BjM�*v\�v�!���{��t ���V�}(��2)Ō�0�u$t�
%5(]{����xxR�m	���I����<�A^�՚m	����Y��G�C66� ���('9M�1Gf|�_l,���4���#{dIa�*���F�GM�g�%���!���_:�����c����֤�y�&N���M� �s@]���Fl>��8omV�R�.fߨ��~��4wPe�aԞ�-�{U��;*^.ڨ=)�pKuS����zN����E��-]���Yd7}��x�~X�%s�vUܰ���T�P�p�<���^�Z�A��4��n�m��G�T�u��W9�l�m�+x��&1�`��:�lN��ӝ���tm�{V&�%o���j���De��|
��V���=�k�yEk{'9^:weZG�r�����Х�%a�<��{^��=&�%�k�%!)f�*<z?���ͻR�����d3r�,khacT���e�:EЕZF�mZ9�;k'Eƞ�7Qp�4��w�s�y��j�!1�H�4�<��T�({5S:�J,ȗ}l���ۤk8A��N����R[&����'�L]b\-�HV�K�:�iښ�s����)g� d)g��i�[6�3/Sޛ�oǨ)��2�Ba:�C6t\�H�<V���w���� �P]��A3����B׺B�X,����OLS�$*�@ס:Gb0CV��"�r@�#��ySBÒO\��⧧r�N�I�w<j�qE��	���v�d�T�5Κ�{.��YN\��R�/�j3���s���q��v���ѐ�Q��3$+rt�	ohBY�k���μ�z����uv�dW���Ν��]���V�j�5�wי��Z�4�ֶ=���U�p��lW���V��+��N%u��I�G.LӦ��	���&wvf�/�AՓ��L!�ڽ�/\�BB���=��#��b:�&�,���9�/*��ىYO�a����v�ܚ]<\�:�n����&բ�*�Z]��c1�=Jޣ���h����s���B�P�H�b���==���sWr�$pG���#�K��p��o�h�/e˗p�l���F5�-8����}ks�#?;�-����L/����PO]"��e���|w
gg'w�fkTG���jy����RO?l�A'{/�̩�N��a� �	�J��O�Y�cm���a��{�e�#�ɣ���/uS��:o�k@�e�2���y޷
"��׋�Yc_�M�q:�J�2q'��X43e
l�(��85�@ZU��:�;3H�����1wM'��T�SK*L3g�7 ��V��:."�K��F�QAR,�k�,�[)��:�]'��Wk���������K2�����o�z��<��+}�î-E��*q�UP�9�f�ƴ�Vn��RR�#�
eP��4�.[�:2ez�	���������w1��Zo�+�nYU3����PJ8&_W�����fzym@�����e�&�
��f�dd���(P��5��t��n���L�8IJ���%`�A�˧Oo�r�:&v]/���ۻ�n��ɉ
�0�H.cGa�/a�i]������f�_L��:�)�Wˈ�e�y҆>�y*����]rl�NJ���ݕ��jVy�}Q���7���vv�k���N��"�ؒ˲�n!�gO�Ej{D:j��mg<�q�i�X��e8��!�n-؋�*#n9,QM�X�����R��n�hB�w�K�9;�x�s�m5A+�9@v����D��A����˥��U�������ɬ󼩞���Bgo[kR��Zg�K�����)R����Л�ʕq"���o��{�X�0�#�쒡��<��x�hOE�peS�
L�)�ׂ8���)we^],���l���@���L�s
�Oy�pg��S���W��(;�O�^JX����uz�F8=[v��s���,P��_0d$��N3*�{���"^�K�9��k�ybkr�Rʄ33-@�u�n�*���oX1]����%�H�%�9�q�>�y^�BoK�+g��;�a���>��*?:s��m�6�yo�$�St�^�ll��h�O�p�N����|r�WUXp�[I��a=BN�H�u �]wVWC[&���k�p�3wэ��qm�W�>��f�u�#^��pV6i7yK�(�����%�&��s���wV�����k����Ȩo��L�$nZkg1�k�5���-M�;�Pf��ֻ���j�de��}Y1є�Ȧ�:ٳ�@�I��Y�k^��ݎ� B����1�ںeqN������S����� ��ʾf�����.V����L2�zG�v��0�q�>]7��](⸥�v�����|��aߨf��c��^r�/fs��sv���rX�O�]��W"�z�:�`Mu����\�r~;�ro:��Eb36�]l���aB|[�7⮨�[M_���Bw����EaV�����i]0u��̍	���6��Kp�B���Zq'��L'[�$쭷�06\*T�J�X�@����!�צ�2�]tv�[P��(9�:�0��mUt�J��-�Q���6�8)��h*q!I�M�@v��z�����3�2JI?��N���r]X9�g	��Z��"�y#�6�����[��ūD뙮}%vu�큧SX;f:����웛��P�XՏ�w9��% k���+Wa%v�����LE{:v���E���I��B�Xk�W*�9ؒ��چ*S��O{����&��-�<�Y˩�NTw:���fL��{hB��u���r��D!<ysRxi���ٺQ��\�wk�7��c��:�A�v":��ӯu]!M��t�r�ntY�X�a�U��&�������b|���#r}����y����λ�}�^���E��ɛ�����i�r��\�2��mڨ��S|x�쓊��3'{2m%��`a��Y���p������g���^�4zj�_�Üw�[�zyt=Ύu�$R���L�t.Rv<��W�o���j+!�yx���V2�֕�>�#ni��n$dZv�#|�{�R*��K�'v���ɖ�+��:�)�:�����g�u;z] �z����Z�L=��-���A��"��;�+���U�+��xx{����$���IO�@�$���$���$����$��B��!	�I'��IO��$ I?�H@��B�P$�	%�$ I>�IO�H@�P$�	'��$ I?�	!I�@�$��	!I�$�	'��PVI��Sb� �u7��@���y�d���fw���ʪAR��
�(E$�����B�#McI"P��T���D��*�Yw�Oy�f�cl�ʵZ��@��3fҤ6�)mͲM��[+lձ�Yi�wiuke�j��x��m�*٦E�Z��3Zj��f���j�&���d���,h�m�1R52�h��T�mU��[,��{Չ��x  ��������;v���ݹ�T�Y�m��n�V��k]Uf�ۙ��׵OS��U{��,޻�mKuWuP��]ܹWM[�^��V*���V�� w���k��m����Y4k�*��I�����ڍ�k�v�[u�4�m6�]�gkn��:���w{��]����=�ʗ hn��ib�=b媶�7x  ��P 
@,X P   ]�^�@ (�޸z@ (�� ��mݴ5Ulj�*v�a����Cml]�Y��m�]3��+63[vs��m-�x ��Y[L�:ڥ�۳T�U���i�s]]5ڭ����+�n=�{۝�iR���;�6ܜ��c�5Z��V+kN�b����clm��� ��Ayj�j붷Xu��{W�m���F��jI�ݩ3:+�]ut��]1M��u�2������ f�(ڔP�կu�P�BuZk]՝�u�@5�΀6���wn� �r35��ci���� �QMݸ��]0$]ͮ���e��8 ���:Քi�vC�Y��WQ�FNv�H��  ��$�v06�1CM�ܶ�a�nE+��;6t9�Ϊm�����6�6��1�k�jRe��F��[� ��D��)Jڙ&�m�a�7v�+�N�s�R��0�m��[�� :�ݵi�wwp⭖�iQ�  ��e���,����1���7f�c]��w]�+KZ���jB�Ӻ�suw:�ۯ{����    &%*A	��bdd�E=��)R�`C L ��& �)�i�IT�i� 20  14�S�����       DH��4	�CC4��R	4�)M114��&� ��Ӛy�8�9���J1��eJe�k|�Z��1�/$RKoD /�y�(��P�UA8����U Uy�PJ#�!U�N�������'�P�0�b !�܁$� �	?Ɓ C�I��*��@5�@�}��:�f��gW_f�UA1 b�&��}���&�	����$�DucWm6L��Y�{����mX�rn�Y#w��t��K���/n����C�d�x�����S?��P�ޚ�����th�D�uo,=ge�^��V��o�iD	D��ܴ��tZ�#�r�v)kushw7F��7 �<y���;��p�6�ҭ�k�	٬�l��Zq�owZ��5))t�P�Gm����7M*��m&��fT"� Q����j"/�i�`��Z����Te�3V�5�MQ��=��iMEj�3���@�7�L刉Q�2c;h��/h�����ow�T�3l�̳�&���9q��Wlx�1Ts7mc�r�ˏP؆�D��{RC*[��J�K�����tAb�X��wA���.�ݧ���%�' ���MЌ�H�f�fa[���x�j;����2`Z��[ԃ_n\z,�FJ
å�
��XZ�Rb��uH�2cQ��b�5�y�v`A�݉��)�'j;�A�У{c0���x��ɢ�Ѱ���7� )R�bzr�x�$��b�@Y�mc5�:B!j��ؤT�®�y�PDf�2����J乙 9Y���Z�)A�l�2�RZȬ���1�p���"ɒCp�bwcjI��\W�.�M,�V��h�c�h��Mj7bD�6]���6�D�ii]F� ,U�E&e��P�� �l���bt]a��T�Re�n����f�Q��5�Vif����N��hc�Cl׺㹤`��K&	0�Uu����Ko�!�YG��VŶL��D�	��r�´��ʖ�]�u����`��&������%�R�a��蛨�ʌ��W)�R��*�m0ёh���+14�K�L�y���٦�nQ�CYWL�#�RL=e��"������,bd����[�.�m��Y�K����v��e�&&eLTF�Ȯ"YYzn�(�Z��l�(�x���6��9	��L� �f+w1E�@�ӵ�M��5��x�S* (�ї"��l�Ǹ~{x-;*&�̤�y+1]fMRfg�LP��^����\�O핧j]�h�vV&�t)��jf͘�;B�T�D��k+D��kd�N�x�{9��v½�n��C�1a���Ѧ���w�m�2�57h �5(hr��Yn�#@8w�Y��	̥�]�]8!�Y��"��&��q]�1�:̻Z�Sl�[BH[��fioI;�J��-�F�yme���¨�B�=;�r��6M�Ыȷ+�[�*�
�զ������iۭ���W����Qh0d,�Si,5D8孼�m;�b�si�.)�AoB��܇�"
C"Z�gE[��m��7�Fgۆ
�F�X�W�@0�$��&�����fIr�:l���@�Uj��֌E�c��0]K�S��2�����^@[NhzY�FKAQ�y	)Sאj��f[���թ��@"v�n��VlU�,EPu��&�Yb21�WS.�gUJ�(]�0[��&�@�1��fVf�˰ћ��*b���E�q^;f��;���%�5�$�m�`����JP�%�y�(�2��;\�w���w �q]<Eޕ6�reh[�ީ�+�fm.��h10C�Q��I�sh E��DC��e���⡺,�BV��������3dz`���Af�*X�8��f�i�4�>�q�)��8��+nZN���a����Q�m3[g]� ŚJ��o���2Fu])n�O�,YJ�
�5�)uKe�8�M^�t˫���z��I8뺯4�n���-iq=T��4V�Q���y2���5���3M\��3&�GNF�&�V�4Y�ڱ��%A��b`e:t�Px�Ͳ�D�$V�hZ^������.��W{1��[+M�E
l���X4��}�E��� ��s\4��*F,L���蛈�WS~ŕ�n�Cl%�^�x�YC1|+���n�0�r��҉�Ŋ]֦l�(��@��DʘAX�:fDҫ�����Xb����#4R��$�ɑФ�J�r�������)f��r ����L�ي曻 �PʹOUc�v���v�J�a�h-2�Z�Wb �fc9B��)^��Gll����Xc�VY�Gq��2#J�`���Yx�WL3��Âvn���XT:&�M���6}�K#�M'kb�+wp��a�n�#1����-��r�iͪW(����gYU�pԴA䂲��ot͚؎�&����r��.�(UֱJJ�y��
�S�1�ET�,�O�\���ݡ�7n��24�@��E&��v�ٯR�2�����z��x���6��9�2�����KYa̙�5Ή��,���lSYGku�Wǈ��5	8��2��Z)�D�s2"^�cЊ̴���F���b�V6�bY�����Asecz�a��lG{{�B2����Ӈ�cKU`�mn3r���+��q ̠4Ә�|��vڽj���Î���{YV�I!�	"\79 ��:j`{�dY�nm؃�C,˗��ܣn�U��%�e=ˮ���, V��i�+�]�;��6�^P����9p��-��+3�M��Q߱۸h=�n��X���Ԕع���8�V���݅ɒ�Gr�y�
�sA���wX�[ڳ��bۤj7L#)���3�h\� ��ww���Dۦ��p��ZA^��Sji:b;qQ4�s �[H1��;��;0��,0�b��ॵ���k"+__+��.���Β��GTPnO�Wt��,%��4R�b�B�^�ʠ��o6�L���Z3"R�m�U3
�q�b`�YQ�X��%�4`�M�Rͯ�Boʷ�s.�(G�&��A�&'J@q�2���sM@��H��r��N�Ŭ4I�L�j���=o�򒅛0Gj-$���oC�A�����ך2��������%����ec��fV�,�yM�n�QO4˗����9�5E���݉��v��y��dG(�E,BZ����(#4��m����^����D�Ew�.���ܤ��ݪ�4/S;���R.���c)�qwe�y����I:@֋]���f��sj饂���SV�K���bn<Y�]�۸$�%/�v��pC����x�u��'�6��r����b�a����	-q©��ࣴj�$ 3/N�X��b�u+L�{�^m��
JE��w����'d�.^^���%��v�Osu�;[#��.%v����IBP���+kE��[+ Zc��0-w��lW�ܬ�I����K`���h��z��p�εt���$�(C5�m���*0����̦n ج���F��:)+��[��Z7-����_�^iq�������ѭp�(G��ՏM%N�e��镙wnfc
}X�&�6�ִ0��aT(e,�dv�M��u&i�a�F@XBɺ�����0R{*]�$���Cu�lz��,h�Uv�7����Ǌl�r���CV���n\�Ѷv,B��-�7��r�5��5��"/c��[	@:��'ti
;���;2`�36T[Z��Ą0SbޫءN��N�U�RHŹ�H�C��)%yfX Xk4]HE��1c4��1fn4����b:�ü8�KD��ɟB�2�R���Y����ˬ��B�]��c#,`q:�v���E9jL�H�3d��^��R���k5{�+�E��d�qFDR��)�6���U�5�5�`F�`�w8�͵%0�Q�īK�+�C�А`ս���#BaP��b��R�Z&��Am���jn�XX�C W�����L�����5r�f��P\���[�y���8Nˉ�6�:.��m�2��^fh��v��ҽ͔ӠMl*Xt��r��H�����kct �Dr���F��Ӌk�g2�H�L'��v���Z��"s�1���K-�G�m�P[b��1�fl!ة��E�%j�I�����A-���a��"��n���4.��+e�N�8���U�?��2�4�� ���x�t���FҔ ��ۏif�B ��du��0+JҞ�YU�L��أ�v�1}B쇌m%k�4,к�X����U�7�[N�l��m5t��Eeŭ���/n���Uk`B�(յ�vQ�"�4��*w2�6l�3��Y���c-� j;�,1�к/.�41�ʅQ��JQV�϶�=Vq���7]G�w��CI���A�
�[�2�f�"���Է�@��l����Y-Q0�y�Q���ջ�V=�f�XW��Z�d.F|\��z���q8�0�7*X�M��MG��09R��:��K�sS5�wn�5.���E1m\�gd�5$�0h�L/(�`�T����$�(c��
�Y���;�̻0�2={�_DB�Z�$[u�#=��V�Ĵy��*�"�l�t��߅�hʙN;�V]*9W�%)W�[�MDF<��X�ș��H����pN�r�o7K�0^26��+���q��: ��gTwy�? 5\�(j���STov�7�Wļ��qZq�8�$��2�ö-�ݦpS̔����M�
�D�<�s"H֬��j�Mk�V)���I:�Jv�-��0V�2�Pd]�+�ݙ,1mj�P{X�h=�Z51��n�O�Ԫ��D=���Wttg622������4�Gv�����V���}�Lg{֕�X�y���m�)��m�Q��m�۶1́l�A$%(D�I%($�I)B$�I)A$�IJ$�IJ	$�JP�$�JPI$�R�I$�R�I$��"I$��6�m�*6�m�)��m�Q�ɴ7�FV�%��U� Ui��N�];P-��*|*��aB9P�h|N��V��[���LI���q�u��e�w+��95X�'1�*1$-�޸sl��/,��w��^�K�����=�e�}cb�3���jV
�k�6��nE�q��-���,Ι�ͰJ{1
x2p�b��MN�<���T-l��1�ٽ�0p��<�h57��Y���k�����I��9$��>��&��i�\��@8xf�����B�7dq'��I;j�V;��XA����(�EE\n�q5}%]�������l]�������aA9���ә/��[*�\�|u���a]qΦ���9]yV�胕���4�t�I�d���q`_G\WL0�3Qɜ:�ܳ9�E=n�YꙎ��`��)�5
 ����P��U�������:�؎��o����y�70<�Sl�E�����Y��e�R%�WÒi�y��Pd)ƯU�p$��l/��[�Z�#ذՖ78�\��]8�-P�c�1�G�j�ڦ���2��U����AYY}���Un�Z�B�����F�w����[�G���麾���m�7����ܤ���鳰�8����SX�ti>Q���ԥp��������c^&�c�B�[���W�W�R��pT�u��rPf�JC���*ޑ�t�@��b�c��W.�~���haՂ�ۤʹ��E��Yr�z�����=La=Ҩ�W��ܟ3;t�"��ɶYͅ���E�T{rJ���v�Y�f��p�� �s��B�żݾ��+�sN<�oeH[���F���\{q�q�2����2�,w�Y3��Sb�!�v�����́W[��뫦��>Rs���:C@��0���v��J�a�
�⻎?�����ӊ+�W�b]nk�5�`J�I����֩��ߍf`Jv;��:��<���,gXQV�#t��L�O�5��>���V	����e�U�\Q��n��ZV�|�q}�ؾ�qK���bΡ.�����`v�O��a;{�`M\
U&�e���f�dS2*+��(��MTf3JR{.^SZ鋗זw��-�-�;��z�P���k��f��F!�������<ҳZ2D֡������o7����νT�8��
�ҟR���f�T��x�~b�{���ӓ������16@�eAWw2�9�]f�5�;�D*NQy �o�x�)�boM�-l�)�.U��U,\�����α�wXX�Β��ÅN��!7p�)���\5([�vʾ2_Q�("������������Ϛ7X�P��E��u|1m�!�9XRW@�n<�2&Zm�L�3�d/n�W����F��+��i��w�Di��Ad��uՀe0������N�J��rc�K�{�Gûy�>��]R�kN­�Dҁ��ܷ�IB�K3dHEW2E��gh�A�L�)���-���::7�wRQ�u���b<���ۀ1���V񒕝��#��c�p�*�KD�<P�36�L�
�Lֻr���p�G>ٚc�;;^q�0@���!X���V�ҁ�?R"���}^}���
��+d�!8Ϗ+�I�%����Ɯ�,��_gv�X�k��q�V����)-:��MU���U���'�b��٫wq=��x�]
O^�f��cn^nˆK�TV�u�����0˜�]w��BqɄ+&��(s�K�a0UayMR�U�"**�lYPf���i��*Gtbwp�[��R�L=i��� "�n��ؘuy�� �z�qofW6��KevU�R��Ѭ܁����&�|���8):�!]��f��
6�^E�v�%0�;{B��u�K���!�j��WɬIO�փ��Th`�[�@��V���C����
�˳R=��nD^WUr����1VF���yYj����L�M;�m4՞�8���q{�z�:cJ�:�*Su@�u`w88���n�.��]���Gs��wR�]fC)5����صf� �����v3u5^��IbT�*�Td�^ԙyh`�%���QR[���X�1v[r�	H�)�{��ft�X:���΁.��.����c�`S�X�9akm�Puh}��A����:ӉXt�%�n-k��i����3d��w�p�mJ	�O&�ODޣ��K��i�/^�y��:�M�`��q-f�K���2�M�0�*)͉`�%oj���x�;O{�s��({t'5M`���j/���
��_U�`�m[sK�*]sэ��	�5oG|�u�����+�,�|��nƞ�ۓp8��["4e��7γS���m�pe�6$�j�9����a�9a�6�TU����Ohi9�:��x��f���ƈ�/�:{�h����[�9��WH���d!Y�M+�Զ�0��[rr ��ìo�1�F�k�x� �eȬ�.-��6�f�@��D����GΣ��O�'i}qkr�\�g�f�wyآ�%�YlN�J��O�$�47E�Eȕ�P����*B�8Ɏ�]�E���t�s_s��u3�>bcB�ǋ���7y��Y4��%+��� �h�K�(�	�y΃��ĴAD��gE��x��};���ڡ�+�cK�K�2�2l������Ʒa�+�p7���H�S;)U�ΌM����FI9�v����æ���9@5]�v)���\U�D�x�w2~�u������\ĳrƢi�֖���;��P�
���h�-��&�.�-LfY{3�m��aD:��^�2i,�ܒ�<Guy��g�4ʰ�v�[�l�d��YN��t��$: �;U!��� c��
��T��&5�]hҬ:v@�����s2��X�N�g�k��������Pt���������.��[�q����Օ}�T�U{�x�X"�;��o��-x��'I��rs�[������V�b��wi;' ��65��{��$��*1�3_p�w5��O7�LyQ`��}�� |,��Ӏ�����ݎl�m����p܎�r���e�5*yb�IX/���SI���A��2�f��׬V	|M�m��lJ��IH�؟3������qi�UAs�	����l�F��XԌʽ.����]������'s����YZ�Y��h�uj(e�㱶3$ ��-jv��Һ�*�� ^K���`��8՛�rdH�v�Z�bΐmbX�s�:d��D`Pf�U�Z�M�,�u�w;}��p��w)s�N�#��L��;.=yj��5.�-�i>�>�*M�O��'�;IƷ��T��2k%.���V��gq�n;�n��i�-�-��yn���`�ѣ�m�Śۥ�����@��q��2�=�O�o��\�j�m�I��{�����b��].=R�`��hb�9X͡+����u|�m�����tU+���3Ao0�_L���w����H��bѫ�KHuN��j:��f��8�1Г���ʳa��Y�AQS[�eeF�M�bc5��ԝڑ�Ζ.�7V�o2�rt��˽��"\k�{K��OWt%+�[��v�2����k16;">_��y�Ь�YBŕ(�[ �#
��@rR�8�8��8^�z�cb�w��kB�?/�fr5���W�Ba�|���J���.�wZ5���^�}�C@땗ٚ���r�X��Z�9�4,�J� ��ϱ��V().�W0�Vo�pTZ����8�q@�SbA�L�͊���hrZ��h ���6Z�X�|_�̚��f�fLӫ`y��vs+�ǩ(��� x�N4+�����8�K,��	�s�+��y3<��g�B�k��}	�qKꏦf�_Ȏ1�ӝ�
��ݷI�)�p[S�;�)�Kr��:��6�n��W*�j@ꚸʄ��>��{:�X�m�;i�u)�
�JPإnS.	���dS{��N����.���-|p��k����ңk1��!��H�@�WQf�SYl�.�;��u���]̛S����1VҎìB4������{b㘮�e�F��*].\F��d�%$١X�8I�x������>G+{U�r@�V6p���7f������dgnTwM���E/�^%F�_c/6���F|�]�1���H���Fd�r��J���s�lWO�*�xF	�-q��e,�Sv�\�Y�LW�����U���QZ�@��Cr�Y���]e�0��2�z�/3�%X��}pb�� zݺ�JR�o��5p31���Z�5U=�����惸%�dR�y�Ԕ�Sۤ��t	*֐�BJ�b�맲^7E�}�,XJ�z&�v=��r8�p�$I�R��oz�VunV�&Z�Lz
�����^^�EL�U9GVFO,�w5S���q��R�Ko�$��v˓&]d`��J�M2�,�<Ӻ6I$��m���m�%FJ��i@I�	ILI��HF]�_ ��l������n��Y՘�Q�o&�a��®�Z��WH�se�s��z���{���_B�+r�%�u>����M��pE˧]�f�X$G�����fH��0�S~�8zqslU�q�/&X&\m���;F�m��um��f1�c�;�v�q�m�F���X�����u$�1`Ae�DP�\�(���s�8�4��v�L[m�+�Jc��FWұ�}�)���x�2vAe��*�U8��)���AAٟr�U�Y�]�&c�[�h1.��.T�%^"M����}�v��\�a��]m>�S)}��q���.Ä�)���	T3F��ku��2=���%X	�ºˢ���&G�������]�Q�'3���뚨nr���<<�Z�"��j��W��N�ڣ�Wh�i��r��i�F��w�P����m
5�x��(K�f��g�fjˡ0��c��[�W^��vV7�:T����G���m��\f���R�6- ��G�=��wR�*��\K�%��lt�ɜ�e�A���GY{#�I���)1EGX*�.|����라����E;�8I�ǀ�*�c�ʮ.���q�Iy���#6mK�[�-���˲�E�1�V3X-�Wek)-�p�r��U�8+����WJN{��ѽ]B\]��k�W�E^���h�62�ܵ̑������]�I���o������8������+���B
�v9��F�R�:+�I���eC��r���H�\�LbP�z����M��3f�g�E��->nԛ�h�EŘ_d���G�.�!�]*�eM��н��3��b��ٻ;�f�ZP�+�y��JH�l_C�C�H_0젫&P�ͬXJ�xe�P�c!k"UYi�֥��tJ�;�J{�Y��iF�3%�mdo���d*�j�����,\��j��Ǜ�	j�
p�n���J��ȶ�v�V��LN�3Ln�w�ʂ�l)�R{[@�90�%�C�FB�â�-#2i ��lQy\���/6ov�j�spӸ�]�Cը,8x���s�m|@�j�R\� 	PW:���[�����Fl�Z���6{�P�DV$E�pY�mfZ�gش��>�&���� 7"���8�owy|Z��u^�Ԫd �Z��P�X�K��s�#+x�G�7�1Lī�P��;]�b���';�ELpp�l��Fn.�0�d[Rt����u��B(�=z�c8pɽ4�a�ե��V\��TL>�>)x�Ũ򽻫�F%ok�Uu�fMa����c���8i�����
#��b�;a����o>�^����4hӧ����᪎�f� /�OQ\�sqQ6+�K�ړ����Y��s;
}��bG�cP+�����y��&0�'.�₃��`��;�9���Ɛ��{��)鴔�(�K�uٛ��+w]����v�T�(��fWSI�u] ��]���7m�dJ����aܸٟ��ث7@41�.r3:��m��.c`v9-��ʹh�͸2b�2p�n��૤F�9}Vằ;va�D)pm����k*{�ݫ�j�c�є������ۓƠ��ʔ��t8Q֪�p�6����N�k�����o��j+�C�Gt�q+ع�{�c�wh�Rd����:�G*��R0u�X�Z�.�P+-��g�{�_s=J�YՉwK"�)����L�+�ZB��ud���yZ\]D�;�{�M� �����.�'�[Kr1�vLm+׼�`���wI���n��U�NqX�+f`��3H��`����4�j�V�z1d�����	tb\Mw|�������@�z�v'����ǂ���I�V�#��Ĵ�!�A;݌
�ŮֵDɃ���S���+	ٔR#xm���e�BՕ�Ϩe0��k)��rC�yn\�ޭ/N8T����j�d�*)��[̝
��N��&h�ie@��ӣ9Җe�R4OY��YLiU��E�̼c�S�n��[A�w����D{*�X5;�y�7�X������4M�r(��"���M�G��N^R��+��1�=���^!Ao*%e�d��:�W
��T8mk9��ޱ@�.�k���rMw'R�f�e��R@
J�v�ˤ�o(X2�;yG�؆_,��Nvu���q:q�����Em����a1,kל�樾��%f�.n�������	֭�WV�˘T��l��%�Ku���e�&��T��^��ĊubC��Ք5R��@ge�g'L٢�=j9Y��R��i�Wf.�`��[�n���0vZ��D�ƕuX�X�ߞv8���|"��xI��u��(�4�|/�_=�Ҝّ'Th���X�1�{f�D�g+���J;�2e���Kov*s�;�v&��dC+�}�����t٘Y2	W]v���-�;W>rV��Wp��F�R�J��e�n�V���S9� ����K,b�N�Zl-������J�Ж�h��YbK~ݬ���b/Ɍ
�M����VoRђT����@��v��MA�@,2f�'j�͎�W]cb�i�볏`N�t�[��*���c@�֥���t�pb�r޳*Y�Ǘ},}zn��{}��<)�O��x�
�r�.�E.v,ŕ	�+���Nj�p���<����vp1P�V�����2Q��I0v5���M�B���b����2��R�7��˱0���X~�>�B�;{����Q��� ��������tݘ.��e�ut�98��e�݌�C]vہQܔ_`�i��9�ZJFju�n��͎Ivŝ�V4l��0��8��d���ˋ�Gvp|5�f>[�ss"ȯ���p��9B'���&��N�C�[�H��
����^��Q4,�w{��u�/�*c�X�8cw��NIpΨ��e�?L� �N�dTe��n-����\;y�e+Y�3��	�3��d�o!���K�SV,�,P�G�n�@Q��C�]���m��?���C,����h�������.�Tq�K`�pt-V}xOc)���u;7���<x0�u��L��rM�97j��R,VF�BLD�OmW2�Ùj�;�K���ۚ;������A�ؐ�j���)$��97f����{k*��0asktost���J']gP��i)]��)Û|[&�NN��g*t��]�n�}�"p�4�ٌ5)̀Zu����n�8��	�RÐ
,HSP�s��ҦJ��u�b���1M��C-�]�hu��}�Qde.eL�
�˚�r�TeR����+#풣�y�K6+��s.༵)p���h`��2.��Խ夶M�8	���K����ć�Gb��h*��}uA�]��l���-G�'o�i�Ce)F�C��MY̫�314ڮس#��Bu��ޡV{j�M�m�_M�wY7���ZΗ��F�2��"a���VfV*�k;�`$�Y��6�/W;���U�e�����.���&�w�zƚ�MbxP�����*���4�yN7B�+~�ȱݹI���Y*T��_l��f
p����i��{	���Vq�\�=�9CNIEq��&�r<`�������Մ�޳��(����$�Ri&@̺G�g\�wB��}�uո�X�~{�7OQ'Nq)3��XØ������z�Xj�P;hmn�����7�h����(���T�V�.��</��*�D�cr*��;�V����2�P�0:��ЙIm[�[�4����"�b��O�[n�к�C&9<ݝ��vM+����4�	FH�H^�ҥ$�]�n#�h	e���9k��K���c�`'ui��]I҇�K�Q�{��rW�6ɫǕ+l�#���K��2l��k1),��q�;��E�jw�0h�bή+a�Z(1��Wk�oA�k�i��wA��I�����_t]���_n7W$�<��pC]^"�_^Cz{%��m�juJ��g��WR�<�x:h���!���V��>J���|�E�6n�wukF�Q�yVV^�4#��r|)g|B��+3E:�{����*�O��bZ"�O1�y�ǘ�,�ќVV���y�@�9�7c�i�O[����jZ �l[��@���y+Mk������x_-U.��K���U�HV)�.�]i�*�k�-x�QKj�=X��fI�0��cL�t���8S�M�����;&���OٜM���=�k1�-��v�:��="s*�چ�|u�6�ً된i�#xA�\�ŽA���r��L�oص�Cv>f0r�q�bA���	6pܷ��i���n�+n�0d	�9[N���oE,m���T���f��?I��vt��YC��st���k��\�s��9|�[#[k8�
+[,pݮ']cMX�v����t9.�Y��L��w5JO�h*��-��жž�Bu��Ћ)n��NU�A�b�-#j@�`�hgmnD�/V"G^v�2�`��u^��Nk=���{7/T�4xC��b���fph��r�q�U���$���}�󚶊�v��NU��Q�;Y��̇3-7�R
o�\V�}!AЊ�7֦�CE��Mb��)��=ą7{��Շ�*pCYtt��(l'��Ȗ1s�i�9u�*+��̳���:��)�)�$%Cx���.�S�j˜�7zΒ�j��k��R�L�nnozȷw�`3V��rs��DD1�5��Y{�����L�5��%8x��,�R������������K^'S��������$�H��Y�)���!ݯ���H5���';�ֶ��Oq�9��vw�-^*m;ǜ�tp`x�T���7�u��+wpA$i�[�圱����`���,
���@�HAE��Hd����O{ށS�L����̮iZ䕮IZ�ֻ� �[�w-�'Hl%���y�����>�:�w�=m�-���4ĺź�+GY*jZ��eM�z'Ջgm������W�FKfJOs��:쳩��+�.��tM2h���8Gk�zC ����Y$D��U��M��/*梁;M��
��'�V�1u�zn�r�{�%A[��������D6� +4��bX:z��/^�����iK9�/e��f�n�u�K{ɻ�����꺗����y��Vs�إp�z��t��m����3���l<��^v^qܸgi����{���
~�#
7t�72��k�ȓ=����ͤ�#����� f����؃�B�ҫ�2�qH_�}>��ڈ�to���`�|��vf�ᨺv�Y���!�������S�B+P�km��Jr�s��-pn����T��ہꡐ�5!@�6`w�="RU�'$Z�7���ED
ʥ��Z�%�|,G����4�{}21H0Ј��O9����$�:��,����Z�+Z�P�a���U}����%���
�^6*����+V,��+tZ�cIW֌�8�"*��Lh�,UU�Ux� �"D^�+EUc�I�Qbe�DLL�*"��QX��4ժ���-�)V��0\��(��Ń�P�^���8�UF(�b��E�h֨[V0F%J�����Y��UVX���U��Qݢ�F%�NڱG-v�1#V1����1(1m̬Lj��"��X�����X�D���n�EbQdU·H�-QU4�]Z�j±UX��,P�F("�A� ���8
(��X�ҌTDݦU��"�t�{�G�,rڕ�����TEAv�b�G�(�����������%җ�'9�@�{��{1�dR�b֚\FZ�k9]6�>��ou^�jx�sB�k�r:��Q'��T��%�v�껭�ȡ��.����{ʖ'�({*���~�xR�Z�b�9��a�mm��_"���oZ���5�h�L��PX����@]��N+V�4W	Zxs��N� �1[
f��X'6����5',�m66|f�y&{���׹x|��Uؠ�J��#�Za��I�9:7�J���G>5;$�B�������bF�O����*�LM'}s%�C��>��fc"�eYm��!;q9>EڟH��+���L^z��Z��
���
5�{ԫ�=�o}´XI�=���VU ��}���U`����3�@��Q�KMh^����!Im.v�V�( |���n�02:�����n�B��R6�Gt&/���]d�i���h�5���D��:rV'��,���f]k��w29�ʪ5�\U�m{]d�o�Fm�,�踄w+1����Z��3)ԏ͑���01E������-L���|��z�
c���o�vX=r�DυҖ����c�Xsa{��ž�{Y���F��sO�S��W4��u�Y�9A.�a�����=�����7��Q�k��ȯUy��4�6)�g�=V�Rҁ]Ϩ�V??�y6��Ŧ=WG|�`���+�ڹu��Q�Xh;P���d�A=U�LnW�U�NP�^A��~^�|;��f�N]v4r_#���@]@g=�ex�ѣ����K.��F�ū_k��(^^�4��N���:ͻ�}< �,��K�ë��������hKf�BfD��.�s��׃=yV�3ʔ�Ȏ�����pm���S�+�Gy�d�6%0z����9��g��tn�?0~]9V�Z�s
T{LO8@'���=Ni�G�Ϗ�~5�k�q��cF��P?
�2�� �ٴ�z��׮���Z�EKc]�L�
�׌��.N�K�ಯ;�XڨRGb���(ow+���*�˦� z`u(˂[I���tu��ތ{��*8�ň�m�*��<c�:Q�i������E@w1W��_!�YtD�{��]iʻ�Fъ)���L�=L������$3J�")T5�y��*,w�I�{r��p!=�+�'Ø?h]ƶ���1�vF
`	�>;�.��M������;�f''�Y��4�)ت���0�e��>'�o�1{���ތI!��9ݎb��
co���0��@�o#-=`�J�5�����z��K�>�8�u�x�0N5G"�Q1�i�O��|������h�J��ף;�;Em�r��#:����y�^��x�)I�|S�@��pb�<6x��M�ˮ�;4����6�+�ꓼ�j�[��ZPζ1����'�����);��5�Gk���W�ny�_{��0R�^�CV�pk�
b]��y�`cb��+n��֨�_���bW��yw������z��=j��B]y��M�m s�
�5�b�*hQ��m��>组Ӭ�EM�����k��.�V��&o��˧0�fH��:�<�YG�lA�M{*
U58o�i���d�����Z�۾6�^��W�P@i����]���^G2�J`>|Z�ᷕ��~V��̶�>���)���`s�,��`�nB��0��Sj����p�mV�e�Z�����v�<*:N�����P�ip
����.[��� a�.���br*�+�4�b��&e���PE,�2�9`�=�5�r���N�٬�����d�'p{4"]��j��iϷ&�w��%��˗��n��J`F��rEd֭����8z��ް�,q�^X��io=Rя��C	مlc���`�Lu�?]�:Ƽ��� S����������S;T$MuC������g#��8�B��#�}p��1]+�/H�׀nt�V}$�S�qlQ����&��:��)�Y�Μ޵ȣ��*V(���N:��/fd�y��EjHL.6��t��4��أ�m�ˊ���VT3�X��,�J�i��/V<2��pb�N��@1��E�_�$���&�^7Cv��z���ւ�N��@d5�T�W����+��g^������Ղ�Q���k�f�|ĳ{LQ�u��<�
�[��X�����v�
�C���[O��i���U�~s-��{��}�OƁ��AZ�w:Q���_x�9�ןM�ok�(����0���v�BK�Z��o��*�AxkD~U�"���Ҫ�I�
Z6�Q�U��=<:���>'�Ml9B��uͪ۾l4xl�Cn�]CU�j��Av(:҂äT-���t��	��e�^F�L�y��3��P#�z]G��
! 9�u^�Z)Y�-�����eX��k�1���GcŽ���Ĉ�"�^L��d�t�gz0����VK��vE�D�u]�Nl%*"��oy�X���[�a�m5�G��rW8��Y�ŷ!{H7}E���C.�kwu�����;�l�vN��"��=T>#Mi���C�y=�Ht&%��n2|[T{)¯%�T�k���ި���;��=�f�^A@xW��f����0� 0�~T�|~K�pA
�h_���]�y�%}1jW�d��ܳW�B����[��l��>�13Ss�ecs�����Q	��͇O�u}|ә纮�|N�64ߕA7Ӳ���&�'{�'�6b�Gma:3�xһ�&iW��;�t���$ש¬�������	/�k"/��E�������b�\)���E$�J-X��C^�[��`��8j����NR2+<�j��A�Ll���):��,V�,��>U䧆���u��t����L\X��.�(��-�g�H��!޺^�:%���EL�����fM8 |9	2"Zm�J0V=�Z�����.�-Y�)��)�4�w#�J-��ޮ�F]ॵ|. Q�[�ˮ|VV�2�U�erq@�2G�W��=|����Urķ�b��1Ri��4�sO3�� �͐��O�ɕp�+=;��ַM������ `N)��}���ҥ�FH�W�e��~�8�Xn���K�*T��
^���w��q���L���O����TC�Sʠs�ht�T9�6�ٝ���/E���]�����c�Hgp׆_/�K��Ҷ޽�JŜM$��Tѭ���,�6ST�c�(��/�")CG��w��nr<S9�
�1r�\j�̩Q>2!+��=i`�p�R,��۔v{�^nǗ�����8:z���}�Vs��3�o��"�n�h�8R����Q�N��E�G¨����ב;����+�=���Z�>�E�9�!3
��¨N,ۗ��I�~�ܩ�o|l)V�:Gؠ��6#�h�=���U�.�N�5�X�Xʇ�e���a o��\JMV��3LR�lU��>���v7���ͬ�} U���D�M8{6���-���U���"����߆:��� ���B2��jzM�̮�G�ƴ?�p�J�xo��ư�Ch}�X5*�	�sД�6*��}��[�|}����t�F`UE�t�J+@XAŊh7}H��\��Hg��YJtX6xzݞU2�u�,Ժ�;=��Uz�.�5�
?b��eq�S+ʠ���,�4�E���`��4]J5��bzjn^�_��T��=~�����r v�۾2k]��O����N��e�_1��>���OL��`�I�6�纄�}p��z��[Y)}uB�T�..�T��\7�0�rE�0�팝���`����u9��B\�5Ҫ�+�4�#��rަ����XVtK7���G��^��\����]��lpm稸W�F7�ok.� ML=4y�+W��:��5cMf۷oI�XR�����[_���.	^+Ԯ��B=Gyc��K�����nu���p*������}۪.��c�=˭�����Te����LF�&\�l;�{g6�b\�bIv]d�5~�r�b�5Y߷�z��6��'��(3�AOT@e�wLtL9Pje��Y���I@���sZ/*Cꆗ�~����4���]C��^���jf.�������/��R�ݩzV��a��]��1L.q����:���8ڨr����*#��"4p7ɍ���V�((��R�}��[s7މ���z��9��PR��F�N��e�
W�LI�m��>nz�W_�C���k�~u���s�������9)s��H��ydVK����b}��� >�/6�/����>��2t��e���䫓����<5��>���6A�y/"Ýف<� �?:���,L\8;7=t�2����Eo��)}f�U��O:3��$�SS���ɓW��l���s9�+�s)K ��Q���V1k�1����s]����ٶ.-z_�T���V��FN��rދ�݃/�T	�7�ڭʜ�0�)Q��V4Юé~��q�NY��!�c�mS;��-)�r���Ĺ�
����
K�a�3�U7z�tӺ��싌�*H��1��kx��C�/j���\'n���n�X!�1μ�Gק�_��Q�űp��O��"�0��L��mh�q�<)�(��Zᡘ���x���pgoo&U�'x�Y����U�������6�
��N��в=�JhaI3�eL?A�ٺ�/&���qb����T]m���3���11Ec�z�)���>�c�m�$?��`�@��B8f3�W9>;m�n�] �#er�ǨR��� �Ϸ̅����]V�ܝ��]���lp�.��Yb�(�gޔ�s��9�2w�sX���n����?#�ҿ|U˯ʽD���K����B��wQ �)�vp���䶍A��5���c*J��xlJOP|qT�� �`�=�+����)V��/tk�*NAԸ�=�@�3��ȓ�����L�����q���\��]'��i��;jV)�M�Ͷ�s�v"�Tخ����+����R
��r �7j'X�0��q飗����0�N&P�]�h����r*Kk��Ц�5ӛ�eǜ�����Zܨ�jZ`u��Vw�]5���cZ��l}��_l;��\y��_+������h�b9�kb=�����<f^�2��V�K���+3uty�J{S�E�]�ɪ@3�yB^,�i\��.%�ɮ̬/w�������@+�鬂���謪e�R��3��b���%�m^�0�v��7����E�t
�!M�u��Ձ]�u�jzǞ�R�B��s��J�VJ���Ô�J`y�G�I�M`���]��z��t��3���/��#�H��q���
�2I�;�?O��?2    pt��_v���ʸ�ɯ_�!�Yy�VKד�8n�Eڂ��T��]M+R�7+�	�������t��r��S{h;�)�ߜgڨnQ�&�^a�f�T�,��­qd92�����!Љ�}����n�)5�PǗ�B�ЀL]is�\�P���㘳�ݴzMZ5���z3��*�q)q <�L��ܓr��X���j�;�j�N.9hr01#��418�xe��\��P�|�vS�Z����;�B�ӫ;����u6�7�D��%�R SF�\�D�(i"�^��[�֞[/M�E�s��E`-����M,��.��J�[���m�7� S.�#�Ͱ&f�د`��re$iM�R夋��3a{�v�ژɵt���ݛe�d�U�#�¯V�y�tՇ�a���4��Ԑ�ںRI%�R�̘I�I'���X�J)Z"���1UEDY�Tc)���
�Xm��c���墋>��|��,T����D����+�*ŌDU�V*�St�6�6�E��e�`��3"�/�0X�TGM<�"��Z
�*+�B�,�mF����Duh��/��/�\�Q���M5D��LJ����%b��.�(��填Pr؂�"�L�̈(���<�q*�¤�ڂ�Q�mX��*�DTX��1��7M�U��*j�(#db)�U���(�DzJ��(�
.��,Ac6Ղ�QES�QV-��]3fȟSj�4ݥ��AAr�*fU����DV�hf�y��̶=�)��-TM5j�b���R�V,��
ܱ�P�Jҽ����>boo|`|��"c�8{n���E�p�q�A�H����Z\ ���;Q�_e�nu��Ύ����	���ߎʯ^�X�/��޸_W���������}1q���3��\}p���~оC�A"~�1�V
U�|8w�7k��H�	��Uu��	Bv�2���7t���}�^S����X���j����5�,�$W~���q%����[_�x+4�����P�2�m�qZ����!F�`�w����֩>_[+�p�Rb��ո~�����۟=�pXyb�S'�~�W�=p~#Ly�������
uH��~��_r��P�A�l�HD�Pe¯��5>&:�ј}Jw��݌��<��rh@ ����a���9��o��Џ��������^���T�{E�Ta�ɽn0`������5����J$3X ��~������r5�j�t@W�BØh�����Tn���ơu��!���6A�P���Hev�+L'nٴ��$X����,O:���f�T�s� �g[y�53���u����:]�EI4���`�'Ø?h�5�%��K��M�d�wwJ����$�C����4�U>55�T60V��k�0��Y?W[�;y{;ղ���q��u|��>�1��G*r�4,�ĥ}]Z桚��CӋ�6Ve�����UETUʢc��zV��=3�{���_�!��߅z�<(6w8v���P��6��%l�&�x���Ϛu�⳯f����p�����km�8%+�??v-BK�I�~�;@�k��@�^ɞ�����������]�L"�.q� ������-J
��Ϻ����Jc��)Y�-���tz�K�ʣZ�������»:�+��5�*i���N�^l�9�5�z"9GN?�E���'�蜒�/���h_
�F#����փ�j�?�����уn���鶲
��9%V��^�j�4m<�s�C�+���?��f=��z~1�cf�KC�٧]�"�hr�$a��7h���rg{�2��=}��
'�)������Y*3��f☌��G�`�{��*�Ӵ���y��}3�eۜ�j`��K�-��g�{j��f)Uŋ�D=�F(�0��J\
�+k�X=�r<��nb0�v��U����c�"�z�HS��,���+��à��ja�8���W�vf]Q�/�a!�����=̮�g��5����;��z�1�
��:�VC����r��y�l������r���> 5�H������އ�v���
�Ɣ~|(-cw���+&�F�>��7W^]�0��D+���C���U��9:����!9u� �Y�̉���_���M��W�Uor�@X}�O�3�z�"31�{ (_ϮP��N���h�4T�,�0?[I������t(���H�)��l�3Z&V>
T�|����Se�%+�Ws˔��9������קV�m�Ft�ܪ �J�4B9�ے�c�t���s��pײ*Wo��{п�C@��h��0��#+�=����n��Hј��Y�eNɘ٫�yF���l����_�οG
x�|��ƴe	&m՚��G,�0*��u�%��
]a�w����Rt�Z ��8;���[�;����v1����)p��e��7�`(�2�=���u����^�Y ��a\Yi���JT�*�\�^�U�N3M�x��G����X�ŉ��-׺P=�R��W���?9���0w�~P(t�w�ŎEa#��|�R:5�*�[��:�W�V�n�
����|͊����X�����z}zmLT�1l[�q>��K���5�yB�7կ�*�^!��g�����PR�yИ�ӈ�/��6�Shmd	��p�N|�DHg�N�l����ùݾ�Sǌ�i�2W��b�z7bP\ͻ�LܛB"�Z]��F]��5 �U��c&`��T��Ħ�/h�odT�^�N�+�O��[��SXWk�M�H[	TM�b����?�dǢ=�l�A6{.{+�����@��ʔ.����hYB���ӂ��gZo����ۡ7&$�5<�Zk���jt
�ʷ�h��z$\���b�&��4W�؎��N�B�Pp�/�̅��:j�WS٣=n;�u�ӡv����z��
�Y�-=f�\���;�I�g&���֛��^f��c(r��2���w���6��5���`�iX�1B��)�uw����mY�e�N�
��P��,��ul��o��`��Z��)�EB��p�V����/�������� �1���Z�F��n��xu�V���ъ�0�	�e��tO�+H�,�l0����_z�4��T C_.��r��v�{�2��~��.�0x�׏
�2�G�c���?Ϣ�=�t�y�ˌX��
��c��/�-���XI��*�ՊVVC�����gK���"`�"~c�~X��U�_�rX;-�nA�Rk�,���U�����鹻��~�Vp�v�����1�G�)�:� ���T	�BLФ6�kC~^�ତts������[�h.� �8�0�Ç~75�f��c�Ɋ�\D����������0�Ds�|�W��Es��Qvk��O�+�ҢB:��]F�y_��V�7�=؄WZ�c˗|���vS\8m�T�v�����$��Y��Mŷcj6b�sw��;�%ͪ�� ���x���!3ɻ�.nrb�L��N+-�o�Z��r�\Y��Lϕ��YX2�V�]F}G��E������QW��ޢ�Mp��}==/VtI�ls(mh�8���g��b꺭���r���Hu]�Zȭe4ù��͐�cռ�P0��V�
�Y�h��Vm�c}x�xU�,9~��l��sO�\��Ɋ�/Z��Ä�/�r�m:e���ug�;B{v��GϽ-�GT�v�"��O3edwgV!�4G�����Q0�nO5��zDK�O�kL�3����ܑ�`�1��/l6�e�J8Ő���3�L�T�����zf=����{�o�o+ ����4�Q��B�'\xhJ��5^0V��{⨕�'�w\+���Vj+����i¸��T����h���0���ܜ6��_b��*�jU��S1|�
�b�+ʠ�kc2���������n/����1rz���;t�ç"v6x;3��i�%p�r�\]�W�����#�N�l�k�"|�w����s&��E��b̩�P<��[��xp�Q�i������"�z�����J�m9��Q���������L�U�jg����n�4gk��{8C�+hWY�oƘ�¼��I\k��?OG�天vb��ėA�TH�g�C�����x���<=B�(����h���ӈ6W$huy�u�����l�,q�B��԰=��ƻ��Qm�����*wa%�Xy�kB �t��f�a�n�0d��G�4�)-�Y0@��Βs�F:x0�RT)��0r&0�v�e	w���$��_`�ǻ�gj
e����䫭S��n�ɒh��wUWF���������̰�M���~�1<|(�.�H�qWL�бl�g��>Kh�<���ԅ�
�񼗬c�>8W�j�����1��1x7s��M�yXN�^��B�}8�zt��Ѫ����٣��{z/g�[�xQB�]}A�����۬n����拦/z�s����lY��fV�c�@�;��(�=�i��x��E��=�RٗX-EW�3�ɫE��gg�CF������aʽby9��|��@߹��N�wZ����C�e)�=@^LŦx����I���+���b��Gn�!v��Q��?���v��͛i�\��[~�)�B��B�b.�,K�-];�1.m_�m]�r72��~��Qa�Sǎr6��^�'n�J��UCT��p���iw��<��G�f�5��v�JYb��V�8��7��wW�CdK�@X�w9�ѷ��6R�J-;3�WW�y���N�ꯝ�UT�E$ >�ל��뮫ǎ����#��Η��P:GF���Y�5(!�#�<���rs���i�� to�������f�S;(��F��"gC&:����t�y���)����y�n�8��v�X�/�� /��O�B�]z��7���r�^j�%��59(�F�a܁NirG�<V�z�c��+Eh�<�X<7�s����ġS�0[���o�wY����5<n�c�m
�H�\'P5�Ṗpv���f��>�$�nlÊ���s�����:������=��-�K�ĩ�k��uj�[x�c��lR\i8���0�\
�<���绐�`۟i�T__Z$��,�,t�Pp���UyFM�2hF���4�D{\��2���U�o�)&m�%;X)_���2�^�e��5'�&v,��dۧm�986E�Z�����N��+�D(7�g�2vt�yw�e1G"{�X�s�68���/
�ӵ��x7��V�G=8(�u�z4o�>!!� ��H����"�E� ��AB,X�b�(�do�����z�O;�>;:0`���Ŋ���{QEB��âFN��n0^Z��s�+�L�b�AHZ4N�(��]lt�}�>�T�*�s��a�}u�ώ}p#��	���Ȧ6Έ��''�o���k��ʫ��u��4P1|������f�=�+h�yM�@�ʷ���Q��ˑ(gԍ1����O�>X(�a`T8¹���,mz�� �lvZ��P�C���I����'P�:T�&vT\��T���1�kKUA�ºZ����]�������ߠ�|��9ïr����Ǭ��(��Zx�g{�c'l�=B�zd�۶aXt¦}@�z�X_��U���p��$���=`V�����4�Y���n���κ�wgz�y�o�]}�~��_eI��v5�0�:a�����1���TJ�'�1��Y4�����M0�
�YY�%g�;-�q������S�g_o�3⪺�҉�gގڏEO�&>��sR�޵6�^�*)�d��w�4�Ak&�^�z�3I���ެ����g��s04�X�����z£!5�����3z��[�{�טY�qa"�
+�h���%m�aDF���1c)8��নr�ۅK�z��i!�(�^d_Ib�(VmӶm};9WE�A�d�#8��+%��OT)nE�ˢ�b��{E�Vjv����y����Lŧ��+ ��bG:ftz���
<h>�Z���rDJ�[a���5�΀����W�D]r�ECqi���4ݾâW[�(."��b]��4z�R�z�D7��RsZ<�м�R�i��#Z�8��;����$�$q�xz���˿*d�Z�Mm56�&�B"7b���W=�G�P�z�����˺έy�y��t�@��j�Ү� �N$�8Ŵ�����hZ��3�ˇxW*�,t�!�XC�Xe��3o��;���N�� ����rtZ7�����]���[��D��*"on� K= N�#[Ů�� k��~ϧ&d�u�oe��N�s����� ���:@VH�!Ԓ�c��ةV�e]�[@+)��̬�M�`��|��[}Z䕮I\2L������:b��{p��/W_9�d7���b�un�8���Q����Y1͍8du��G�R��K��w�7;7�pCE ��VU�.��W|��ݐ��ZhZ�,�ܥg2�����}�v�Jo��q
�"{5�c�.�^:U�ŷ(4�m�{WIv�
D*彮Wf�L
T�e�������*�1PX������B.̱�U�G��e��:�U�.�P�r9���S\��K]�W0gn��QWM���������%��w.rQs�.�����ZEjR�b�R������p����P��V�.��u�¢�ͬ�1���s��cevws�عZ�Xw�R�L�Nj�Z��Un�pL*0;�C����
[`����﹪��2����+m  g�3��\x����E\�۳2&�P��Wݒq6n�X�fX�c��ԩ���v�YY�>{��Jc��ZH~�eE;���m%����<���rHaF���9z��7�9�s�s_�?�s�R�b#v�m�?��Qc������za�Eb(*��P]%kPuj���h�)�m�QU,�ETX�*����QA��EH��r��V��u�wJ��k�Q�����EF"*�"����)F(m��`�aE�ZX�\d�1��Ŋ�U��UQV*����^e�UYݯ�TMR��kl�W,_2�U
*0UQV
����EH�B���L�1Kh�JT`��0�F	U�5JW�X��SV��AT�EQ�Z���'t��A;h�Tg�Y�T��X��媪��T
��rآ�d�F(���(�*�TD��`�AV(��]�V*��Z"%W��w��n��M[�TM�;�V*(��`$U}��}R�.�J��>k�T��;�d˂��a��t��%��Gv��BJ�CM��K�"=��E��W~H$x�KI�
,6���>d�gy�;I^0*u�6�Ht��a�vgl��I�����c'�E����&��|��M����������F����W�E ��N�t�H(o�Lt���� �x����PS�y��g��1$�:Cy}I��ɶ��:a�S�
Ι*k�>fLL��"g�0�}K6dmŌ������
A|d�1�����!���{����i'@�*A}@���¤<��i�i:a�4�%g�<;�H,�ex�}vg:�����^����<������}�Lg̕���1E�d�ɶJ�SG��z`VՆ'��E��W�J����Y+���"�^�w=��'L��|��s��u�_{��R[<Aex�Q`v�q����H,�e��Y1�hx�AH)��& (���d4Ι+&�f!�K�!�����Cė�+"��+<M��m�g�˯:��9���Ki�d��i�y`T靠�ͲT��Y��=M�(�;k8É�����I=f!��H,�{f3�J��9q�	������`%U�������٥��I���<a�;aXi>2�<@���F���`,�Y1 ���X/�
Ì�3�B���i���Y���$�ě�PĂ��5�9��w�uמs����T����c8�a�|yC@�Vv�'_Y��ɴ}���%a�3�3l��O��Ϙm1�d�N W�
ΓL1=@�;�#�m}��&�knx��2}��T���Ҥv�_��I�R�7�&���z�$�{C�z��9t����SY�x��6e&=0����vi �7l�(��u���}�~k�����:�|��m���%a�l>I_�4}M0�
�i.�;�3�J͝���tR8Ύ�iOZ��W�O��� �ǅ����M�gL6�>��'~�y#:r]lI�5Q��$N�xo]��T���~b�㧟^��wXRk)�7+ȷ,����fgo`1L��9nVw[D*Cy}�N��(���a*��NBK�OL�/��G���ȷy�f=l�f0�
�P�{g��8�Y;j);B���xh���_]s�l<aXl�����
�Xv���UT���q�I�o�&�X��}��޺�k���sw���B�T�������3I>q��Ă�&�1Xx°5��R���N���P6��K�H,�o&����8�ܤz�Y|���y׻��;�����E�O�a�q��h9�O+�q�M�Vu�Y+�:��H,ĝG�*)�M���q=f���LHn���b�>��!љ���/��~M$z���L�T�S��=���Ϭ1 �w���=d�
o3!�
�2VoVLCi+�<a�+
�hvS]R��]Oi��E ������R7��y�>V��{�y��ư*z�P��ͤ��xÉ��>a�c'Y��O]���H)m�l�����Vb)6�g:��4�Rz���=|@�aY�=��Ͻ�޾��y�k�M�Vi����QVMO)��� ��YHT8��=�*N!Y����� �v�k�$P��!�����T�g����]�|묾��}�뿀Q@�*|y~Om ��4�~b���;�H,���f�1E��ܓL�J�\���
�'Ɍ4§+�큌���3s((�q����׿��ٮu�zs�}/}�>2TXq��z��EH[gϝY���&��Ι�*C�H/|�'�,醒ya��%@י�Ì+1��t������g��߆w�����0�z����+=a�k
�T����a�&�d���S�z��`T��ή3�& (�h�a��aR�8y�M��Ho�O�{p�_5�>�Ϲ�]_��+=d��E'��S�H);O���oh���4�h��|ʊ���2V����l
�8�򐩈Ϫ=s�y]{��G����������A".�h�%VA�f��$�ʲ�q¶��IG��;�"P���M\Zk��#s*�{�u#�f�ԫ=6be�6�9���^�5,�yf�9��I�UUW������9�}�4�Y���9�H)���Jæ��*�i��4�P4�e�N�bAg�P�4�J�z�!���Xo���8�R��2c8�Y�"{��_q>d}�t�LDV�z*}>��d��� �����={9I��J�&�����~ޒ
CV��y��H,6!ӌ�+&2��>C$&m�޴wG>�]{�� |n��=�q�My@:d�T��9�l'L񓌜`y� f�,2G�33����sO(z;�_g޹�O��\��k0��0�bo�$Hh�=f�x l���+8ɹ��+9���M����W״a�:=��t§��=d�0���{���۾o�����;d�5�}`W���awHT��<���b���H)��V0��P1�Y���y�u����LH&���^u�Y�7���W����W�)+>9O�i ��nyCL���=R��J�2W4�^3���L*z�5CI�I��{`T���4��QCz�Ǧ�É�u�Ϸ~Ͼ�ϼ�ߧi!�y��T��yI�|�+� �I��4�� �}�@�>d�ݲ,6³�y�H(t��HVaZ��f�
��jQܻ;#�r�>?�<��>����^�v�Qd�s4�_X/�|�� ���g�=Ld���H,����T��\L������1�d�+=aٖ&c�3鈩6�4���a}����C�yI�{g���0�ݡ�6§����ed�>a]s2�2T*J���ul����6{t�Y�O2��T��K��H,��{~�|��ν���<}@�Ì>�XA@�+~öH(�=~d�S4���%|AaR:�ܓL�J��Vz�YċR
x�^*a�*t��u�ϻ�;��w�u��ʔ0�V�pRg�����+�m��,�p�L�d؏+ŋ�ufۇ��}\v0M��q
&���ŉMrE��>Ⱥ�eJ��_�˜<^s��	!:��{�~s�k�v�Y��Y*)l�%t�QO�tz`_�:�>f�
�l��Nw���(Vo�&$���a�*�TǢg�>�K�]��,����{�CJ���aa�
ͿZLH(|�<���+!�.��%ꐩޯ��gl*{hu�&3�J�uO�$������Ă�����1��f"�Y��]p����}����};H)��;f�i�g��1��Vc5>���&�i�^���]sz�!�OH�C�a�e&Ψc<d�=ew��`,钦��c��"����k~Ƣ�~�6�w�%k����_,��Aed��7�R
kۤ�v�Xo�}@���Ă��W�����Y̰�i�M�ĝ���e|b�gWL;aR�{��^�~����}��g��!Qg̕�!�bAO<q�Xi�O��H,�=a�l�O�Y�%}d��s/l�M���ü�֬�*ٝ=���W_]�}���߅��Y�(W����3vq��I� �ĝ�] (���u�;d�AC_y�����V(v���q��Vq�NZu��J�<�����\�}�����o��Ă�'ڳI�:Aq!�Y�xÉ��V�Ag��8�H(�$�����y`c'���L@QI��1��d���<�"��LD\����U�}ZP���#�+�k(}�&3�J���~�"��2Q ����^P4���݆�4ä�T�MfM$�Ă͟Y3��;���A@���˳���{�{�{�fӌ1E��ɴ�>OXbOi1�l��S~ka����3�J�Y*oT��6�YƤR
ví٧�
�l>�|�R
i���*L�Z����r�s��z��ީs�|��R��j'�� ���՞������X���M�M$���Xq�C�T��Y�jwCH
,=B�8�R
g��������x�ϯ��u��hT����^;��mݲ��U-b;жӬS�R��Z0�R*1FZ�2��p�3-���p�եm��ӄ�f�5`������9�{���<��=�~��7�<I�������H|��d�ݚgl��������<d���!�*A}C}Xi>g�. t� ��L��H,��5M��Ԛf0�]�ߞ��{�=ϽH,���{O�4����>B���c'l�8�~zd��VaS�� �=d�7�d�*�Y�6{f��!�y��+X^Y��\Ǣg�0G�K�nۜb�R��@�Q@�YRiĂ���@�ϵN�i ��)��>N�b���Y���>XɶW�o���0��2�g����ݸ���2T�󮵏�s�u��}��oݲ|�S�}�}HVM��&Ӵ
���M2Wl�u+6�_���RY3������Az<�7�=Aef킋��r�Ă���Rm@��>߇��g'�f"��g�S�נĂ��ZL@Qa����zxܺu��.�1W�q��u7}�^��]�]	uC���bu�Y�˿�98�n�ܼ<\ce�������UGK(A羚���x�<+�g@�n"����^����w���U��q}�S�ײn����T��;�F�VH0�z"���TD�}�m��
77�sk~��>(}�
0����Os#]��V/Շ�y���ޣ�k����i���墽촰��Ln�J��f�پ���r���)���ahw��C�Ls�a,u��#9�����'�(^SE�F�fr�&�j��R�IЂ�ִNZ�`�\8F�w^��ӊ�͊��u�ʆL�V�ѺW�����HSn�*lP��L�
�.Ъu��D><(���S�������w�VuW�h�[�ႈ�5�C�f��X�93�&r6���4�e8�!�WR���Cӊ���/���ˮ˂f �s�E:�>`X���w�nzpu��V�T)t����Po��=9t�#pm��7���b�����Ș�9޿)'�K�r�[���p[W#�GB��w̜��a\Z5P*�<6ʘ�"���q&�f�٭o�+�:_u�dZЫ�A��b 5����{y_�,x��q��u��X�rg�b�����&TŘ��Ll�V��|*M�(}��e�SfPB�K�S-�ko=�U���LL��E!��r=����PC~ּ��|��F�r!o.��Y���\7�k�t猁��QL��Y��U)gv�\�30Պ،:t*�r�X����ƥN�H�!&�ӏ�"J�l���ԮS͕��`��Ң��K��V�HB�'~���ލ���)��Nw޿\�wtbl@�s~|�r#F�↎3�^z��o{�Ϊ<Z+��~���K+����k|u��X��c�/	��8tw��FP��5¶��w��o�F5��N����o83o{�,���`-��\�
,z�\��՚�n�ӳEɟyHz&�./��U��E���¡����pי���g���t����\I�~��q�n�n�
���޺aQ����ˡ�i��d�"�Ƈ�ʝ�!Tt�Pf�������2!Q�ReJY�;+xT81��x�t���4ѭ���I=pX�?X���R��W���LW��V&�O����%�(���W�����3��t��s��^����Y��e����}c��X�P�D�?c��[w�M�㬪�ص�	�f�f����#oe"b^>>��g��nP�����X�#�2�_��.5����.$��)8:������J�EV��Y�:f��N���~���z<9�Lvl������n�LB.�����O�U�fF�)3�'�vI�zb��K6�LJ�"zbM@�J.�Mך�X�]��S�Y+%U5u=� S��;��nkp�|�P��Y<5��_*P����\5w�'�%`�_n�L��5p��_?���u�h�D-5�hT��N�����5=��C����_��:�e��^�1�E�+�ǰKpOx�fPT�.���Oޙ��t��;b����7�9���Ug��˜tf����B�?B�6�8Eh�/^{�{K	��Źy^�k",���+���{~��ڲ��y�z����&I�Ø�f(<+�~5:0`�\x�^]1�QEJ�*�J��8<�{��B�h�n����E�/�L5}f�5^X4h�Z�<�bg��Xt߇,�ץ�w\�y��j3ׯ�e��{v	�(B\�Q���.ӳ�T�WvKU�R74sP�'w�R�9��ĆF,��/z
^�J�����)A�D��{��RI6�g&>�w�,�-�.�������ޅ���g{�����I�l�n�An	]uS�~CUE�]b��0x�׏
��XrjV0����^і�9�Q0d>��*"c7��3+�³*���^�o�yF��pvi��JO*T����\:���A�,T3�!�'l�y7u�B��(en��J��Wr9����W��\5YW��.|}*���L��<C�YU�<:����Gǆ_�T�xxp�g�%�q&���(�3��$3KW�/r�5t)���c��ԉ��g�p���5��G�B�q�������Pc�9S||��ݮ�A�u�^��8R�NؘυY�^k�@�T�'�oC׆���
ꄞږ�tT˿�Fvr���
���ެ�c]X[�B��tF�a�/��9]M9�y-{LM�W��b��of�=��s��X8܁m�.�kc��㭥���k�#�Hy��G/�*S`[$D^_7��@s�j��D�`�k4A���F����T�74k�^ĺ�Pؤ���\��ޠ;�#1�U�T�{
��ã!��P�qc��pb�pެ�3�Q�{$�i�yu/	*�W^��'�M?n��/#F����0cxt���p�:*g�|�Af�U����R����r����=⟙�\0X��߼�j'S���n}�!�Xg�Z筲�s�3P@���И������4���?�΄O�N���ۨ�5��Xk��~��Wo+�,u9���*D�37V ����n���,|��R��A�6j��f	t�T��/ޡ��:���"�$����v�8�yYu�[��Jo£dϔ����}NY��1��烉w�:�=T?,+KF�
��Ѷo�1�𮯿kd�\���_�v���]�p&��>�E�r�寑�C1����n<8�3+�tJLd��qy9��e��k�}*�Y1�K��{�;�K��:�s6��6��\ҧ�Xu�&��Yz�&&\�z�s�k�/m�ҭ�wd�kO׽Ó&kMhg��Ӣ��q�� ��"�ל�tA���Yy��7L��k��v��܍m� Hv>D�:kn�a�چ�PL��@�:Y�Gr�vu� 7�9w]��i��ven�"�������Z�tI�g ��=�MTt��j����v;�-�6֌�AбV���5P�T�*:|zQG:U�y���Cp��w_+@�*c[�\ƴ��F,[;��7ڶ0�YgFT����zS����6��lRy������	�3��Ui��&Ҽ�|zHuT���I��l�M�q;�o�VZu����,���^'�Q�4e�f���IFx��@�b���*���u_�$���oM�MI��(��v[��<Ń+i�Gp��M%�1�8̤U��
��Jč_N�C����x 9z��<��	�V��o����Ol��Y�"�,��z�J8�\�
������L췹-���ts�ɵ��)�|�5�h���"�ei���Q+�bb�@<|+5�6�XW+U�P�ДO\9Z�mN�mN��f��r�Հ����i� �i�]*&@��	sJ&��x�V�2s{k��bf܍��}&�K�{u"�(�ٓbBگj�]���F$�/3�Ü�>ܷ�g�n7*U!�
/x�]Uj�f枒��͑H"���0�TO#Yn�U�����0īj]1��=�Ysx�Cr�v��Ҩ��ʠ�tX�zU�߂&WZθ�D2�Q}�XɊ�P��T��>�s^�)S���Z[/��4W ۡ�&���*fP�K�E)���'Q=Z+m��r2+�f����^�h+�L#]���+�M�P����fm"dq�"rE��̘o-G$W�/�$�kX�V��aEV,��L�E�"'�m�\�5;LQU�ЮR�1!TE�閗DR���ikKl��f��o���b8�QF*��&�@q+��S0�����3LW<ޱ]-�*0q�T��+��Z#=��/m�j"�+���J�����Ԩ�i�إ"�iO.���n�eq��E�F�D��k�iXf��ձ۴�5\/�QfZ����ъ(��ы�cmY�5������4[v�T]5�i��Ut�Z�4�E�*�,��ch�[im�j[E*J�(��F#n���&���S�� �'�~�E�t^%�HV��M|��qu#�6(Ȣ�5ݞl���5%�.*ƕ]�d����G��"��ܒ,��U��'���KB��8_ʍ�� [?M�S�E_r�]�]�^Uq.&5׺��?��F�J[� !m"������e��	�C�2V�Yo=��j��iO.�cpcߓ�$g��;����P��x'Qp�V�(�Do���u[�1��{���zo�ce�c&�C�����#��
5��F�W�,�_�+�����ER�X�U�
q��`��;q"`�n��H��s�M�d	��Х��dhB��\c���J����H�虫�u͞�����A�~�b���62���X�ف3�ѮE)��y��r@ǫJ�x~K#�a�8hNk�K;t.�Y�8
��w�{�ђ�����j�|o� ۘ�]'�ȹ�"���k>�)g�d�D�57l��k�V��L����Q�b��K����6j���ڔFP&>�Y� �wkJ�)��0C�N�3w-U�j������q��zF�-F:d���z" �gH)��1?Mw5�Wf�Xk�|�f�z�����);����i�A��M��Q��]�f��6����k�/�n���� ���rE]iE��H���O�ҕ�%��UR+g���ɘ�td�����Q����~��4Մ:������
_4?�caC�5(1����N������^�hv����O�v�s��n!☶���%
���*�}^q�<��z��<�~p�N�kC>�:|}���t��{<���<62
}�D�t�닂����̹�5l	n�[3+�Xm���LFO}�xW��Z�W:�˚��X�B�&��Dm:Śn@(���u�^_gm�L �`�}��TLoS�����r;�CC�0�=�X��O�n�0Z�<k���q�m�@��[�q��HB�8nC�X!;�;�Z���h������	м���g��ᠹ[�gSZ�r��s�`���&�"V�#wM"�T�Pb��F�+�nM����"=�����#�����Ⱦ���㠯�}|@��I��_f��P�7�G)�3j��QF��\
B��l?�ꖮu
9��^v�Ғgr-��&���"D5nb�]��
�=�f��*+�إ��Ç
cM��=H��yLRgw�ͯQI�"�JmW�( �a��f�v�]1�9�	��從[�^a_�t+ƨ��`����5�h؁Y��xk��5a������)�bX0`�|01�^ǕW�ۋ���I�����Gm�;i�h�0Ӹ�G���j��WP\������<�Wu�6g��-�0�ژ�x_�u%��J%�0���1��5��
nz��I���}WX+�z8��pk�@��¹����5�]x��ŞE	�밵�{��*���X{+��$�ҕ��䈵jr)�AU	G�*�2�ZJ�
Eʺ�̏��z\v�:���p3�A���[; ͨ�!���_t��:�hA��93P�k��K	����O�M3he���T͂К���Ǵfܕ���%Cu:V��oe�`����z#��	4�����qa��z�r���b�\'K*"��>u���q���Mp-�('��*�*�.�� B�\�!7p�ډ8��%k_Ã��)?���_N����3�,� tQA*�X��*��5l�=�d>���L!AEgT	3UGx��0���y6�s�8M�>�����pU+�;�������K�u*�L�;)�S��؝���DMŔG��;ಫO�~�qB��pb���w�"��9�/M���;�[y���vaJ�t������?�aC~�����Ƈ�X'����1H�=�~�����ӕj������n�T��Hh�`ژ����A�,B�6Uyp�s���
D ���4����1���HL�k��r�E�,l?yz�Q��#yW�+�D�P[]q>�k#�,5Ұ:Z)î-��2&�4�K�!9�a5�CH��tN�Ffݲh,q����*�/@JA���_�ވ�t#��O.jcǰ����*�������OO�;�F��I;�z#N��Y��n��}eٜ���p�ON@���L�.T��ݲ���q(���m�g.�E�Z�UU��Q�r+�U�Μ�>y̨֎ۼ391b�|�k����~�|H���4k9]Q�k���@��S�(T9�ƨ�Ӄ��6 Zk����q�S�Ξh�m������*\L\*j��L���ɂ|Yb����;��s�*ƻ�N�	f�S3~��z�1\)���0�T�n,�NB$X�
�KW�m�\�Ցx-��i����"�줡�/���R��du��c�7�[�J5���\�����kq�vT�5��a;����/()���
C��Ǩ`����0h%ov�>דӸ��O���#�5�D��xRAr��g��T���V7��긷X�E�gn5Ü��ι�ֲhK��y��z'��3���iĔ�d]�]�=�%}����4�qS�U@B�`���pIE,SX��՜֎
ʹ�UtY���~�ȓ1.�9��Z�L\����UثU-��e�m�!V�Zcy�ll	s�f�Y�>��8.6X�ޯ�TN��o�jԹ��OQ��(OH�c��7~5�������B���gd]/o��=ܯ)}���tR�����Ab�nW�`��Z���Z�p�OZ2��M�[�H`���t�'��5�أm���R]{������i�H��6(��h{���:�'>G��^�tT
�)��hp3����j�R�X�
)ʚ4��2������ԥQ�&v��+i�F|�٘˭���t=��N�LB.��5_��+TUG;'R��Bj1�����=m�>�=���<_}0���s�L��Y�g˅ʦoa�lW5XD��C`��-Kõz�kc����5�������[�a��wٙ��NB1����r�PZl5֋s'��U���蔀�2���Cr
�[�T���#'#!��|�h���AP*���|&��C<���_�*�<��~"����N�^��x6�[�� �U�c��NLӧ���POPe2�ʼ��E3��b�>�����NTK��zj
�Ĵ��u/��´r�t� l�B���KƖ�s���b3��a��^Vz��h:�:
�����5f���ǊG��;[���$�EˁFGQ�"�M\Fx���+���{~S�s����c�Ih�M�6�U���@�Ʒ5@�+�,p�ʛ/��Ef�(�7!�]�*��l���}E���W��\~�/��V,p��;h�tH��c��V�H�'Owm�8Fky�ns�3`"O�xsU\>#a��*I���'�^�^q3�#붤�璑ܽ�b�s��U9^�ZX���,�̏x��O�ء���L��*���uMj�:j��P�V���u�:E�%�*N�Y��U��lb����z=��<�g�mW�%״�k���Lw�ܭ�N߂�f�}��R�pu$A�BT��ߞ;���n��b��5����\ߌOI��6�P����8��87�0&2[�t'_J�<kFW�»*���Ю��"�i�t�+��Hg�p~?�E�y���K�
���'�Ҥq�L��Qγs�V���B4��*��j��>{3�ˆ>U7d]�v,��&��=ơ:�TJS��/�����}x�d#}C��3,�����q�է� Yj�Nw��h�4��<A߇
wC�sΆ֚�|*����������|���VU��y"oXΝη=9\E\�*�N�~�^sF�B�����il�';�J��5eH{�ʐ�e`��p�۩�^�a�k\=�U�c�m�8������$�<�F�2ed]������3]��|�^��]^+��!	�֘���YU�f[�|&��ʳv���t�r�C�6Ďcio۷'�����1wy�W���g�Ci�2��vk�<*����Q _���T�F�Kci)�3�K7��F���2��W%��7��":��4�SI��i�'qqY�3ӳ��˺���I�U��΍A�z����]�Q����Zq}`��5�ʠ�5K71��ӯCAoВ)����z`�\43p*��hb�.?<�{���:����F�}^�N{'���+�C�������Z�4�����tgϏ
��k�F������,����!���E9J*^�����Õm� #M��{ד}����P���xT�#g�T�E@��;#i��*��{���u�)��e����Nq�s�*�Pp�F¨@��Ҳ�\(�%��Smft�ĮV��J�W�.&�]U�/��B4b64�2l�}Re�"l:p�����q3���I�����%ecB�9`h��];�`z�X|����XUi�WL�I�WY���s��Z;��J���w9��!y$�G��wWޏy	[i��Ȝ���Lw�P���foŻ�#M�XǊc:]�.h.>�eذE!�k��P�����@>����I�5�݊D���S�@�S�P�U�)�q|�~�:��\:5�W@罸UΞ��}Z��z`���q�������({j�~�j$LUE���^�\}�ɵ�4Ŋ���Uyh�\�@DU��s�])m�š�ZA���6���u�K��p*����t�˭^8��ثR��W�M�c��G�ÈA<<8x\���|~��4����?Zsn��~RM�\�ͣ���K�jv':���r�C��z_�=�#����W��v����v�R�u�)���p�\��}-�A�*���L�A>�S��� қ�e*'��l6(���+��u\M{�U���i�˭jw]���u%���˧j�D8�V��l^\�jP�H����
v�^jjiw��.��ԑ;�3��: ������1B2˕Pl��V>N;��c�^�rn�|b���ݘj�3j�"��#��K��_I�"֢�*�s��W�;�ci���k�A��pn��mq�7���ǘ,���^�3lcJ��ّV�J�Vn�W+@�\&kw��9��Ԇef����mS�a�yą���e/!�܋�R��!���S7��S�1u<�����m�=}Ne��ut�&�o�K��OG�B�pT���5�ګ�v�CVz�r
F�16�g%�:eV��]I��C.���o���� lww[�Am�K�ue��e�������N���2f��K��1���V�\�N.�W,������s$���
�V�=vS��ב�����>�TveC���>:i<�Ӵ�܊�K�6W=\��gVPsd�|Էj�a;*,��+��/Q|�v@��c��8�&)��%�$�L�Y�|�d��|��eGæ/0Y�+;E%;!����cZ�0��]��ZSb���]�����_���p���q��үp�ʮL��*\�)����.��Adu�Y���=��c����g!6�"X���̭�7�U.�������FZ�B��&)B��K���6�t��3�?�o��*��/Lu�����]3f�/n�І�	8��%��j|U�A^�ug@|��<���yU�fCm�������G�ۅf�"�����3�͚��qs��+%��&Na��ZU[�78��^�|-��Ѥ�K i&�t."�#^)�M5��$|�g�b<�_hO&�
�7o{��*PwP&h[�<=[�����a�졁 ҥ�M�z�-qc�W,I�O�,��U�p��X.�:t7u��[��$�$&K�.ݹ&N�����wlR��k{�5�[A+b�<�46U�
+�\f9�U1����)�Hf�Ո�.=��1j��2ʪ��Tk%m���R�&	1�ʓl��4�T�P\�+V�(ؖ�9�����f��Pv�j��EQm���:K����i�(.[*QE����5�)�J�9�C��Z��.SY�.9��a�bf�Lը��Wg0�2�/M�*8֍�%r"#Z�Ԫ�,̰����J���k�ѵ��.V��ܸc"�ŹCZ��Rѥ�QZ�e+V�UV����S�0C���.8��j�亂q>�a�an�;H���,��e�#��7�i|���FP[�\�o/��j}(�M�=����cv��8>gG"t!��ߍ�W��IW@2�s��DXCި��Q�H�z�^<>ީ�=9&��i����+f����[>��NI&1l\=��N�LB=ŵp��ڮ�#a�^)���n�J����4e�C�1.���q����u�q��l�8qO"'0����3��qm���x=��APK�QS��Kp�^���4����fD�Q��~�k�n:�Щ�J>��m����X�\=@����AYvF
�e]�@��R/f��.���O�d���P����^��5N@�G�@���ǂ�lS�i�f�m4��9��0��
�i]�Tf�_ˬ
���Imi�懼�냂W�S����k��ʠ�Fj����~��Ww�Ǯ�f��*R���@Z��QZ�>��	�h
zWQ�X�A�ujʶ�M�ٔ�&�N�4��6G_ZH9/j.x7��oVW�`�c�\�i!�49|�������Z{�o�uY_e`u��j���\x�5�¹�(����fm�Oy��a����):aʉ�7�x'x
���
 ��87�S�X����K��FU�]�5��9�j��҂P{���}�'�Tp��|%����ˇW�Wa�Ux�]K�ǽ�7{	���܏���1���Ӕ)�?^�4�!�*�h;��i�Bo���A*D��ߋ��T�60�Leӗ��Edm҉.�J�^1�˪��Ӄ��堥]�&���ߜØ}JG+�쾕9��s)����5v���۬BSܺ��>L3@}�k��_������M:S�EɂP�gU޵O"9T7��ɰ�ez?�� (�]�i�q���כ�ۙ�}�`Q0y����U	ЭG����� j��������pN�4]%"���s�eD�$�c!`G1��Hq�%��'ćbd�c�gB�cpʚ_`�ݐ�%0���Ah�2\�.q�񪙄,����U���צ���pS��]A�����  ��_|�9$���N��{��Cǝˆ_}�v[9����x姖 Yhbܥl)��=���C_������9�}B��tq�^vӾU�8�Zu�h�����8=F�^��.�����^}r������Ϸ�a.<����(��̜�XM`�f���e��}=�/���5Y:Tr]0�谑d���>�`�{�ث�Ci�,mVk�`5xwŭ5A^��]�t�Vɏ�N(ha?/.�5�x詔�1��K5��/�rN��}Ms��ޢ���R�r�ON��(� ����C^��s<c�Z�Ԏ
��|p�e{&�l0xS���`�7D'�+�鉴*�ɯ���������Ƽx�A��e_/�֮�\�^ؾъdNN���U����F_*��Q��hN�96�ON@�Գ�)d*��y��N{=�R�q&N�9����*�>�ַd�Y�`iB�M�f��b2�7��̒��[!�-Z��GV�dՖ�q��U�y�����|���%��<3Ή�Z4��QR��`�}�s5��理�k�G�J�UCS<xLvt G�ݪ����wa�Oԋl�����R2����}B.5�ګ������*^b�\���;/���hO�%�jnyה�q1j�����U�B�Lƚ�K �Ӹ����]�ΘƯ�=5o�e�5�*���F�T_CӼ�4�#&$�8���P���'Z�p�}�
u��U9p�*�ϱN+[�lßS�ጅ91�}^S��@��5�j��?�_m�6N��d`�}��ƱU�~��#�ܥ
!�����*5��}�ƩC�Տ��{��ہ�(�(׆R�:6�;Yנ,~ޝ�y_m��S؆K�PR��|q[�C��Ȼ۪ܴ���b����b��LL=��:-��cs����V���-:�X�P�[�F]��Y�\)��(���X��5��O�YU��y)J�N��&0��oVz��q�}vv}�v���5�b��S���ͺ2'՜�� �l�C�9�o���}N������^����G�w�5�C���Nu	�����^�_�S^�O�A.�iʠ�R{[ع�'=;f�7S��f��
WP/]p�::�U�'���p��b�h_{Uh^!�)�z5 �ɾx򲑄7��Ր�5Qy2��oև؎Y��),��p�Nl���i�&'4s-_��n�
I�9	��y����n���	���=���^;��.Jʌ�w�5ւ�[w���\:�g2,T&��&ն��j0,eC�hor��}�����Վ=�){���\�(�	Ѝ9]8%�Di؄��m�JцT[��`�S�d=K��5fuv,L;�`�v1t-܎�������"ef7��[�V�]��ꥑ��5Y��r7���H)2���>+x>��{!Ϗqʼ̭Ӆ���
7�)oU�7�@RH����qVZ�!��ㅔ��n2�)�P(�)`�	������w��}����dhw��8#�0͚[��j�+X�w^�����謗{X�C�b���eE�jL��=�3u�{^U��}+k��|��3Ɯ����0v3���Wd\Ӿ��bqU�wf�e�9��F�ݾfxvjv/�zTu��Cl*��e�b3��|{o�4�d�L?!;n��;���	�>k���>�u2��G��uA๬Dz������s�e��x�-φb}ČKxv&�ֵ���#���ڨ�[���[ӥzS���{[Y�m 3p ��G�':dS�j��m�Zq��x�Sq������7J�\��\�7D%*a��wRHa�(���FbU:4���Q��n���ci�!`u�ȹ؃Ѣ��bgf*ϸZd�\}<�h��Be�8�D<���4��=�Jx�{�u	e��kЫ�؞�E7x��喵�HZu������
n
FA��1�5�`i�K"��xnk�䢹lu�
��+T�Wi�Tw!���,��n�]f(F�|1h�����+����L\-�B�n�楞�/X�����@�� 4�|���֏�����[](.�mX��Cݞ:�_/8`|(���ܥ�eTKӶ�����S��u6 1l���דm��
�b*ĳ;�
�n�؍�ȴnf��d����ueL����}�t���լ�Ys:��h�f��(�gF�z{. ���T�j�^\�wox�r}=��s۫a?5�T(�'�;.�{3�I��[����7�\=�o��@��V�?v��C�:����5�n�f�����<�VXe7}�8n�֢�*��u��Ö��ĂVubP�ddꉱuү�N��gH$����{Rk!y�Y� ��-���-%e����r$4�C0�l&�7U�:��jќ��&3S��n6�m�ldۿt6g
7�F�y�z���ĲU�o�/VaR�%��|_��>ї����ȝ��wiB��Yz
;ϋ~X�㗶�&Q�a;�t�D��m��n��s/ʲmu^����<s@�����9{��#�er��3���t�$�W�c�HZS%~��h'HI��;zk���˾�q��JFb�`��u03�$�\��\���V܍ �vأ��3ި�����k������V�M4�;=�6w��1	�+���^��ҵ&��p�g��H�%��ϥ�f���T��Ox��l�ߙ��v�u�`��O1��ń�P�e����W��ϨP�Y�;��`ߓ��X��
�83�̝|�T�h��SL����"�4�Y��#'mܳ�V�ޣ��i��
x'	�ӆ�P�ag��.+�U�<My`\�����Tvm�Edm�d��'yX�N�*�eÁǛz֫�q인hR�"�����f��}���߸����^�� ��u��Bq�o�:�\4%�[HG_gʑ��\�5-a�n�G��v�ّ���=	�'�o4��c�o+I�킔<F���ӫ7�oC�����Q��V��Z�3r�V���uO2	�����r;�}z4U��RL�n'he�|E��8!�}^F�(lM7s�'�����D��WC���K0���,��{vƘ2Ow�<)T�ʼ�~�Rھ�g%{8��v��Ͷ����z������"Mc4��Ô�Q�����fX����f����j�ڋ�:���U֦sUtVm��zk��ܧ�x�������^�E�hG;�޿��j#����R���'~�ɱf� 5ul,chR�|�=�['
���7�,��]�O�d�u�6M�����rR�Յ�3�����2:���UR����� _g;
�Ta����^aͱУ)�Xa�5-7��Vf�5
�Xǖ�΍���Fܮ%��ИT ������2��
�����PV�#L�����:�A�:ހ����A���f|a��#w]�U|��P:!�Q�K5�
2�ۙ�4hJ��[�vj��qFT�	��MZ�w������d�u�m+1h�%�={6�Ic�v��)."��dH2��N��b�d7�{Y�����nu�ۮ{��	���@MIh�@^���m�r�s��BbaD�GJ� ���,�{���^n�&����[�9;a�]Ҟ[D�ڵ�B�3C���05.�Qxu�� ��2Sv�o�hݜG� ��od�kiW<yȴ���0�Ђ�ϐ��&�c͜]�"��8&�Y��gJ�;&�;��Aq;�w��Ywn+��%�q�j�����l(����+E`���1cv���!�d2q��a�7Pm� �(b��ݵ�@Y|��;{�������BlgCg�,��c��[�0H�(t��	��*J5��vY�`*��;c`�$���d�7�^+��U.,k�z(.l8�;���sM�e��[&좸:���!��{1+8�0���9���{xz�Cgb�m�ê�]GeE'�2u����\�Gl+�e�.�:�s/�[����L�8���֖�45h��R�Պ�z+���02���ޔQ�X����oa��#�.���Nڐ���<����Ȯ�S7�Jm��e!�)�L�.����|,'b�6�!cE��H�j��n�(�%X��]{�kG���D�Vt.a�yӛGS�4M��(S�Q��R�gm��4�w��u<o-����kҥ�˧���s���Pfҷ'Y��˱l�>�x �����@t��:��ov�b���ǒ�_�Ԫ[�,U��2��bM����|�g�\\�ɉ�Rq�=��l��X�� ����i_2�Z��֗)�y�j�jS��V�ڥ�[n�U���Uj�Lp1-��.QimZ�:�2�"2��,k-�-k_rU��+mTTwh)�����J�R��2""+���maF�)S)�F��Z�t�y�ꆰ��n1UDE�[�a2�J-��*/��j�A�㊖���Ʊ+b��Շy*8����=kV[b[V,EjwK��(�Z*�'�#U�Uƹk<j�e��[�J�("����/9r������;Cp�(��TW�#�,���֙���P��gʉ]G���s��sj����7�� Zw�}_|���[��B���p�rA�싚w;����Ќw�'[����yS�^�;\h��}���@�^ظO�GN�Irax��-�]�k\Z:�tU��4��78G;lz�^d�0��=Wƞ�ɸ�M��ٞ�l!=C_9�WY��P�އ��
{bb��*�Q:.4�p$hp�N� �]��R�T�70���ۼ���ڦp�N�0�9�_��iq�r�;		5#"�A�3�LoT�]Bc����-�&�r6D]�xA+�^fz��w���Pp)����]UԱky��f���{�#t���]x+o3�Q-ۻ�3S��wP�%7�f�B��74�쓹mf�X�H5"��ht;����R���@�s�q\�+�Z�Q0������]��eq.x��t�g��J��;����J��=��m� ��e��c��ڧ��gT�o�^f�2��_� �O�2����:��:����~m9c{���p���:Q���[�Iy�c9�[����|i�`�h��.,@|N�����nE]kW��"wӎr^�nX�;r�=�4�I��OKq;c.��g�C��7݈`�*�Z�Ӊ���v�.�]
o8b�w�ص��nk��p7��J2m�{]:����I�u��,,��������n�G�=�N�7F��
5}7r%N���R���lD�$(�C�nF{�{+�"ѷ Uf#e��5�[�1������2jf�}��������M��il<pr�5q���3��M�	}���~�{�K�v�n.W���b8��l��\n�6tF�e$�؛w�TQ�յGJeh�^�424��X�9�2�P���M�N����}�ӛ�W���BP����ԍ�S����E[3�ŝ����.C����+�5���I�S���c)��g����sx8ScXe�Ur��.5xU�q�޹x�oE��ɽ���O�@������#�=��r��;mrA'�[��ٚ��6��ޙ&W�\����%�~�N�����֯$о�
�v�=&u�##j��LB�%8r%��U��;f�Ѭ�aS�41�*���FR�[�qUB�+.4�D.������&.�5^k�z�:e/��2JE1�����2�ȭȺ.�`�;�mp�ᰳ������Tq�L,#$�'��EeP�J�ü�ih�A\�l�M<~��^.�ׁ���m����vX�]�tdZ��h�����T�i�`.�3gU^��qM�Y��姌��p�����9+��Z��,�s�#��z�b��xڞ�����a#�!�Q��p
�.�~5�#ʂ��5�2�s}��l�,��{,�>��2�2�q��{��NҜ\�H�p�ň�A�� ��\z��f<#S|E�D�U�1$��^6��'4�D'L��6o'ωUk8Za��l�W9B�%I�ԷdC�`��S��&�]��bnJ�9�D������H�zޝ����Zîاv����aR9C�J��`��֝N�h� L�_�� G�LoJ�\f�������4YSo�w�Yr��w��8ؘ<�0�����^�r/x��"�#ؘ�Z�5i<i�6��lUݛu<��ARŹVz���t:g;՝!��鉫�J;MF1���6(Z���&��Էz$����ߢ̶����<��	P���yu��.��)w/�`�f����s*�J�y&�~�N�j���o:��s�� <f+�'�;����+�n�����W{RFH��o$�s��lU��-o��,���.,���H������
d)��ŋ�X#F�V
ؕ�ɷ���i��U���;�(wPV,��/ۙ����5Ĥjt������k"׫�w\N�]��c%���2zFB�:�0��BrP�Å���w���rINZxP�G_ԛpR6��4���� �7J��=$�=�	���u8����������Tv�(��i��,�,�n�QmA�]�S��&�;aL���^d�������E�
h��f�6�$�x���N㈗C��򺵃/u�s1W˨��MT���Ke�l���ԡ����ޥx�F��E�r~�Os��n&rD�|����;� ]��a-͇���M�ˈZ��)��y6�'�����w_�ʣ�'���D�˻<�YȔxSr\Ug>��Lz
���3�ܽk-x�[r�m��	z�}�y�&�7+�1�6F�P�	XOo�@}�V�r�8�w(!�듕��f�c�D����갱u18�#��c��ʬ�]�꽙(��A6���D��7�sn�t�3�+d���aB�����_�7,E���絈Zv�0 ��KCd�xQ��`5��~�˪R:hZ�d�i��l�e\�Z��O4v{f��7�!0y���8C4]��ik��"������Z��տX7&�B�a��Mr�jkY)��uAoM����"�n�%��Q�'D� �+������f�S����|�B�;Q�_Ca�ȝY��)�72�+��u��_t�:Ceۊ��T$ˠ�[u#YmOT<7ċ��;<��+�s2���i/%u�;P��Ȣ �u�;+�-�_��.͋���A���t����WJ��YLnK̔.A��ܔ\����jń�{��}�*{O�yK+����\x�h��'n¤�TP]��@������Y�N���,U5�Q�f�/�e�^�~��0�����;-��L�E�C�V�ĥ�S
﷮ٚ��87͎���a�O�.�>��� ��o�WR����.�	�$z�͎�� ��zs�|��m�Ad$����GX̸���8 ��E��1��i��h����O�Eop@��⺢��Z:�f�VQ��nkr�=�k)���_Mv�\�Ӆ]b4�����{�p��.����I��Q�\�ޢ���LX��N�=��U�F��AI0ǥ��R��E䖯c�|&���\��=���6�"�l�M�!����h��G�j�}�r�Wjiuӕ�����r!�&!cY������!��2�$������sq�.��X}��E���Z:��ɳ/�܅ތ��=\�*q�"<Ѕ�h��/=7i��+���y<b�s�	���q��H�5'��r��Z�j�������cpΛa�k]ʣ�1�X^V�.�j�ck�Ŧf�'�Nnz�{]y�Y�:5\7+��ELb<f�ٳ�E���35�&�<#�U��r��gb�[��<w�V�F���y(�i��T�<Hz<KɂQ�Oɳ�ϞŹVӳ���YWӷ�Ԟ����!�0s�=I��qg�??z���Yzگ����J�o|���+e,����EX����q���WZ��������Ƕf�4�Ȥ;�BbuJ��o��w�l'i�]vzQ��{�1�͙���xs�(�ʇ�M��.���e�=5�H���<���{��!u�IC1�r�D���]���7oL�Q�K̫��kq|
{bb��*�e�J���v;S\Y��1��Rn.�9s���jh��/��˾��q!�H�1(���f�ׂs� 2�Cu͋P�3&�o [0ْ�ruB\�&ycE;T�j�t�%r�sPB��V�qɡ��s����qV�e��f*�lU�VTJ��hD�@�\p�vZ�PO^En��G��m9�w�
b��,a~���Xq+\�=�2�'r��N�o�zic�wʘ仵�`��]�ܗ�Z3��v�%���C)�{*d;��b�"�ph7g��#{mϚ��j�k��� �4by4����+J�Tэ	O���_��N]q{g(b�c|�6`�����"bY�8�f5�*��%\�&v�fp+��j�YX�pht幖ќ7�H7���6:��Oh�+N7;�%�Hatp:�g�̮�]l%<a���Ž����%��R������CM��E��o&�<�1۸�%�oU��(pg�T��sP��FnE��Z�Lb˺ꙉ����R[b֧4��F+�ڛ��X����NEJJ��&�ޮ��x�\��]�D��{М����ikG�諒�d��I��(�U/xoQ
��1*դ��#M*Np�Q��-��C�n9Mm]k��sV�Ҳ��o�J�Gp�rXq_�Dw[/	P�v3�����)=h峿p��k9���m��I%zӰ�WSޑ۝�j�%}�k����X'v[췯	qS���9:q��|�;�}J������
|���*��Y�)��7h�#tp�JY�
��u�b��ʽ��a��\ӯ��2
��w#��u� �z���ػ"�]��3Lp��Cm�1�o7�b�=����ȭ܇z�G8Dr���t�Վ�W��|gP�Y�"7�uL�2�@��;q�F8��,�����/+&zӗ1E����]H
����T��	t��M��ҴMu���X���M��������ob�� ���[�0r�x�b�3])����w�073���R�kc2M��fh��:��b}��Ac�L�����F|ٹ�*Vp�Cö\��'L�)u�ъ��\��R�a[5:�r�Q�)ōʗu\j���Yin ��a`I$�Qܙe9$�&E��Ɗ*��QX���KJ#"5�(�[ѩ��F���Q��JPV[Tը��U`����z�Ȋ�#[�v�vTFn��.eYDE�*�^\������(<����1�������-�cݕQ4�:\Ʌj0�ݸ���U,Q��-t��"�Am*�*���{M��0��ݣ:���1�=�ň�J#�
+��陔Q9J#(���֩���K��X�c��YZt�Qi*ժ"F�vw�κ�K�5 ��r+�y�:�W�Db'wt�m��;R�譗�[\_�U��a��m~��#y�f��#ao_��4��Y���*��x/M�(|�/Sض��I���x5�� �qk�5�J�W���lnf,�ө��/
M�S�q��c�Y�o�_Dż.+j�V*��5�!3�E�-��9�#��z�i�!@��}��G\*@��=�+�P�.�{���=��Wᵄ�����b"CӮ�^*VN��xj�r,����bP�dd�Y74��^A§9_GT����DN�T�IドY~ǖ�
}��!�N�R�!a�ge�s��=`ٯ)�kX+8I|���q>�Fk�x����'U�b_q���`Kn^5�wn�{9���CEe��$�l�7�t�znUƙ�s�Iuݺ��������ɒ�� ��|9�U1�"����cI��p!�8�]��:���ćp��V2���x�q�FM�CZ˯VФ���6P~��w��x� �G�~�E'���E����k؟:J�=��c�-;���^c̈́��b�
5dI;7��eZ��7�f݌�uTsˍ"�SYe';'&�YWO���W�X"�6������GUL�T�gC��'�4c��xX٨��b�1�M�h�s�q���(;��Uޔ�ğ�mYpr���Ύ�ts��HiA�0�J�Y��	�h_�{GVh�,�Zѹ�U���h��=���{��=Qׯ��n��G���[���	ho�b�^SNA)��h�XLj�'rY3G=�n�T����_��;�&��}3I\`�O@�G{NiE��[=\@e�jqO.�E���Ό�Qٶ�Y��
͜$�������qΧ4M-�.�4�WX�(��M鲔��(up8E�6¸b�(�:�B:�5��5��
=�N8�"ᚩ#�"�h5��J�L�㺳�W���,���<��G�q�1�XGpgw�U4��nj
 [�1�$DD�~��|�F_G1oev�z�J�����	���;��tN�Bw/���ܪ�;�a>�aQt�'����)	�=R_�#�T�g
�]0�G��ů�C�f�cփc�S�9���i3�X�;�kv7�K.��.�5Gr�>���ę�#S	P�F*0mh��ӆ]m��ŅE���0����I��w��Ny�Ԟf�� ����*#{)����x���(
���4p����d���twd
�/�$Ĭ�@D�ց��l��2��0K3�z�q���A��{��h��x��Mn�#���1����H�!�n&�,�w��v��Qi��'�y�Q~�B��5W���7���z����T���W��iu�6���yw]r,�{s��E�ֵ�)���C��B��u��V��#\�ۂ�$�"vB��$�)5�_G�[~�[��h�(�$����1�u� +gyg��wr���\��n���A�ڟ@c��R��3.-vI��'b�'[�+Uw)\V�!g%e�Y	�(aށn�����܏����'�ne�J�4:�JE�f�4[N�v��;��4�k�|㴈���х��c�j
stԧyr��������/�Pq�m��j*h:;�����=��M+6�(�l���/�1`� K�E,��=s���-�|����q`����%�������ᅳ��nDp|r�ߚ��-T�Ѫ~��:{&�U�7�i*1�Mz�"c[���}��d��7B<=���^W�=�YG;&���y TR)�O"���Ӓ��S���~�թee�x�w�륹��?.y�A\\ru�V-F��u�M! �k�w�lz3�1J�Vvח(h/���+7v�-j[XM��wF���y�7a�MC��=ٗd�	̀�x�:�\��I�*�Pdv�j������A]B͜�����Tm�F>� l�� ���wd��0s�]�Zb���jіM�o-V�M�D�Q���:u ��׿M���]���ڈ�Qc����0L�:�Ƥ�m>E�;9�>�!��J׃7Ն�E�fT���P�8�z�=XDn�eBM���������-�e�D�hp���#bhNwvFOT�a�s�L���n,D�)lnk��AMQ����8x':�-ۊ�Ƽ�9�bΘ�2�aؾ���tpJ�{��n��ޠ������nq�9�;{ޖ�n��F�*n��vyٝ�������������6�Q�Ӟn����5�{v�S&9��F���Ǭ���A �ڙZ�ߊ����+��R�ϊAu���YΡ����ĵH��2W���S���~�y�
�r�Fm���"��6
M�H���`��͝�.k�	O���4HV�-�����L>H+zGP��܋��3�d]K�r��Ɛۂ��#
J�R��v2Bo�L�!H%�n������s!�A8�z���j��5gE٭Hb�����ծ�C>�dƫyuXl��ӥ]b1}��4��J7QG]��INQq��U���籈�T32��B����p4r����7Hq���·���8�����;bl\$�ѹF�ڍߪY�S_��F�Y5�u��
י�iB=L�ڴh7��Ø��%�q�╕t2_t�wS^5F�*zypqj��k��:��XK-Z��-����X�m=.��ok�5����ʪ4)~���Arm��~�1w)�$����#���K��֚yxC����Z��X���ć���8咊�ޚV�7V����9��T,���nQ�ǨX�q�թ��|GVg�q�j7���r��'oSk��fФ�.��7|o�q)I�vṂ���+w�n���CY���F��g&i���N����A�7������_�ӈbܳ���:Z)<ђn\/��]��of���e�>s��(��]
r����m\3Ä�K����`���O�4�G@%��팾��ml^rշ2fFˉ`�ʰhȪ��c&Gw�2�F����V<�TB��,M�}��f�7269���-�̝&�m)9^��T�i[�z�hm�:O����m�e(�cx�d��
c�Ț��v�ZЙיe�b޵��`��mw�YJ�tK�p7�%�!A��o˲VCnBV���Y*:��Xr�r��b�X�pknQX�٣~�E��YE�W��嚧��3'O��!�i�v��N���Ë�Ff�)��ª�����E��k;\�����o)7��yOb�ۯc���Ԧ� ��m�p~�x��vn�OfEn�%���cn�9��&�V��g�Oz�ʯ3<M'��w���^'ʃ�X�3f/s��}z)U�h���鷞T�����״�Bg��R��G��X�Ÿ�$p��U�$�x�h=;�/(�8Uu�r}6�v�o0��Ӝ&�O+�`�䂒�W&e��I&����i�^Qn3f�^�n���u�p��9���S�/�a,z|�wm��G�Z�Ⳏ���%?7���op���Η�s�U� _��YW�t��AE'�S�/β�iv��H��w�������{�0�[M��,�33j��7˂{���z���Z2,��������=�]��y��ʱp-I�N�*���P����β�+�7C�4�S�^�WҊ�1��g�4�X-����/�����,�W6��oD�����=���qM5�BW�F������1o��_���0Ĩ��}�5�Fv�Uh߬��}��m\�!�\L�#NR��}����muy�0m��DOU:pa��ڝW�.��̀�юΉt�%S�pj�i�?�^c�V�K�X�N뽋z��̬d���(�c��:�*�]��F��#��	7lǽv���;r��X�,9wR�#�L&v�r�!Ի�9���B��N�u��<1�6��a���vTP��:ѹ��&�H���_E���6;�ŇA]�	�b��N@�k��mݘޫR���p�mW�;�CJ��4�Bw)n�艮�J>�^���ޤ���ɵ��Y���X�ȳ�ړ���Vku��@�:+`�!�]L�tq�ޥ6pB�о���p�z���+qc�}b�9b_Y��.�H����Ӯ�r���#���G��;�n�eak! N���)d��7�eT�.Z�&�m��[���U��	E"-C�����H�
�B�ҡ%�{K&2�� �B���6�P�]��%��v4b���| ����P��f��#3:��\{Vd��!�d2�T�9b��ۛ�7S]G�Ӑ���]��6��o80i V\�2\l5N�#�W/--Ν�W�F��@�8�c�x���^vh�Q��9ц��id��Vwq�D�q��s.F��(l3C�a�;�9utL���r�Ϯ`��⨘�B�8n�#%��A��]�Iڏ>܊+'��GMy�FH�h�^�kAj�mr7U�C�Su��!�*��Z�&�-q�k{	Z�7{,d��ͫ ��fq����v8ME��A-B�V:Qέ�[�H5���ww5Xq(Y�"��:�[s�T���"�ʭ5G6v3Ν�P��d���If���z�(��6YV;�Ӥ���OhH�)D��b�%��Ҽ�V<0��w(�lJ����Й����1a�����p�fN�rW6�����Pܮ���Jj-E!�f�.�\��t�Ă}ظhY!���v�
ܽS{6��w¨��r���u�.l�;&8n-�����2L�As�.[���t��;�a����b���i�j�g���D`�.�]��T�b*���S�бr��ǌ��ӊ�b��{��1m)R�^�ŭE^�(�#T��n��N�ݳ��{��f\�m1D���f\M4W)D�*"�"w�o{�+y�P;�b*(�7h�b*�ݪ"��c"(�TP`�iiE�Κ*"�
�Wz�"��%feTPX���*&�h+
�)���31D�f�f��T-�c0�wJ��%��ь]Z��cZ=R��A�Z���uZY�[B�[h'��������G�V ���x����[�2,6�1+���r�㸦�h8���j��Űd��)*̪����.���(u��d]J��8է�`��3�l��÷d�g����P�2�ũm߁n��;�K>ݢ�,d��q�5���׼����W8�I�<l�wr�S����#m\F�>�ۦ�*��e&�����q�g��`�-�8W�B��̇��ݣ�=���&�pMzx�7S����Z��lk�.���kd����i;�G�A�x¸�K��WCl�Qc�qVArKb�߳����P\���M`r�I�#�	��8	�r�U�`s�ݪP��A�/;ج6��Ί+����/��V���(*�[ӉCZjuŰ�Y���X�Z�<\�%ˣ����\���idB_%�(]1�K��zP�g��	f����Ke�<ݙZ�Ҕ��Ȭ�Ul^	��G��<BLTm����!�hw�̜\�u��
��,�ڵ�cJ��F#m#bvp��f`��s��Z(��F���t�7#i��8�FV(M^8��X.�[�6�;fN�0�\(�)�\э��v&��(w��E��j!! �A�1U՗���+T�*�|�37MƥB�spJ�7��mM��)�Wmh�OW�:�3˶�n��=�5�v�\����Z��n��v@���^[����	jz��.�'�	��[��/��&��bu8FH���C��x�����!s*n�Yks�T@΄�0�^{0��Q��{:��i�v90�p��߃�-I�� �6�M;I�쭃��<-�eI�]]��9�b�E�+���3w2�@C�&�k]%]zj�8��;#�v�?�U�Jx�N{���_���Ʈ4LL�{~�=�P� ��E�u�@�`)o��ε��45nk�	w.���� �U��/ �9���of�`hC�$�&J8Y�J10����:���`np輔���9��i,����N�ȭɕz462X�2�vF2�� �=k5���o�)�ovӋ0�A�kgJU�ں�#Ẏ�r�C���2֋���s�R+�sYP�S^�C�����ʴ��c�Y�x5�X�ÝӼ�F�E�̚��O��{��#�m������j)���ʶpþ��4{�C��B�]��s���B����uv�u�/�J�����\T#W,ɵk^ȩn��Y\��(�Ôv�<�@���`��P����[sq��>�G��i�m�tf��nc	탞q�h��vuzk�>������%��)K��9:S�阎L����n�f�n�k/Lp{)��4b�#W�;.�ה�xZw�//K��qz�n�M�8����`��2=�}�y<Ln�Cc�rwî:�͚����Z�a�:^гA�c���*L>�#�k��nx�^�E��n"ˀ��O~�^غTd`V�aRgF8�+ p�t��EqaJ嘹������00�ipj�,=�F��Z7S;�uU-�ڮ����<��{4�+iE���ہw��Z/��:�R��\�N�r���Ƿô��TF�=�!P9Z�bȹ�J���2)X9⏯G��1L�d��)ˁ��g��1���mЙH��{�Bm�Wܜo��b�����y�h��H��ėx��U���VE�c�54V��p]�X��;���,0�Ap'\D���me��|���;G*��V���٣q(ܣp���A>���Q�ul���[M�b�s���
GI��s���h�٧��zL<9��}U�Q\�����L�&��x��s���:�{��V�sqa;8�d��Ÿ7��h����%~��Wsn����о{|L��P��>�	cx[�渭���Z��IJ_;/�<�:ѽ��<�ؙu�,˵�}��Q<a�Β�yB�E��	��5�vd�w9�"�9ǔ�5u�+���u�:l!tZB����7%[�I�hԨ����YG/5!-\۳;�-j��#qo,T�w��<��L�|��[�����'u,ꪩW�{�ʤ�N�5z���_�:�k;��.�
9���km��ֺ�br�
#�hŅ�$u��ֶ.�|_��R�`�t`�z��vG���j�FS[��M.[�F8?r�;Ō5��Yёe>"�"���T��v�t2b�FhUVt��ǖW�>ȺwG��WnU���n"��t.vp�zp1=&c�}K���hd��-�K�i���8�
��:rP���
�.::�����>4nQ�F��6�syC�{�P뉫9��Y[�O��NAH���3q����+�������p:��ޢ�f�ľ�G���)*����7�ב��X�O,F����]w���06�]={ǯ�*�B
��Go��}���=�����G����c��)��C�^G�m�-�����v]������IO������U�E��+v��*E�%���ێoɛO#�����`%x���W����W��u����k��%N����sZ����+��&"(����G�pT]�*y��#¡w�^
ejy����������j���g��J��(Aʱq��V��z�6;na�̮:�,���|L�A+�~T/qnv��i��O,Nv�Y`���ԑ޴�p	��3����Wr� ��nǎ�%px=k��q� މr��Y5�*e;:�j�:����N��v%�*�Y�,.���&G}s)$�"��#�q;�R�e^rx+�X�;`d�x�VF�K�譼VcDt"�t����ܢ�&󲾛˅n�N��q��j�ゕ�1�6
l7y�A�EFWFW��u�(�O�щ˳b�cS(����J�=��I6"X'7wÝ�����Tj����~�^=�4f�1t#��^U�S9�L� )-�f���i,]~�5p���Y�� �`L!N+^��&	�;�ꚼ/��x_�y"����Nu�g��ZUm�U�\�x���Ȟ{ˎ���8i"g#SX4�1K�Qjmo�)�U�sܞ�Ȯf24TcK�����v�X�;�;}|f��T�*�l$t���w�=����~���X����ݘ*Ǌݑ^�d^�K��ۈ�J���95�x������	�̕���,1��4��� �w�3�rPQ"2g��F���l��L����@,���q!L.�kr,��-1ѣ0��Iu/w]!Ǉ�7����
W,�O��y���œ{U��2)L�����==�Du�I��EΡ�ūB R�\��֦|��f��MIZ���_��๕ZxL��S�(���ߺ8<�ci�&E�5��2�.���ei4�������s*��W�YuQ�ҵ��Ji�]?;�&A�kں����a�UǗT1���z��$�Z�<��i�}�J.O)R3iՑ�X!����=����A��u��Z��1� )�eQ��ZѨ�PY�a���a�)�M��9R�-���+�f*��3�ra���u��L6��i΢�����b��\կ�͠T{@�Y�{U͉����$�:�&J_DCE;�ϥЃL��aC�5�7&m�5�>S���Lu=����4�ߔmx�Ve�<��vr��7���oP��{˱g��r5�WӰ�����3m)K5#y�g>�=oJ5a��؍a���ھ���p�M\L����S�u�� ���|��q�;��
$Ḵ����oE�,�0=/�q�4��(��j�
�ٓ�QoN�jq,�ʳaګ)k\:�$�؂ ��`�ҥ �adWF�n۫Zdةz� ��<���҆D#4mX��tn�rbe��噸i`L�̽/-��ֳ��\b-���Ve:��U�7Y	>c)���h$��Fk�I鯧f���+z�t��(T���7^�m8o���,�]�:�>��"�0f���\�)LV}cy�wA�]�虽BЛ&�m�6p��3.2���Ef��迈�G���q	�ѷZ�J�f�A��Q�U4)����utË(�{��e`�OM�Å�u�e@�9���:�p긕txȧ��u�g��֎-�s�.��U���GE\�JdQ����S��-�d������!����#�L8���h��q���u)�ᥝ�1oGK[�$�+���˄��,<xɱL�9u]m�$2��XX�g&���v��]G���庢�PC�pA���ң�F]�|�]B�A)_"P��y��t����Z�廸�P�$s>sO���5xT'1�0J������ Q�^��������H�A� ��NE]dD�|!���v��U�[7�V��-�xUnC��^�V�һ4�zn�/^�Д�vh;@}1����n��������2�� $�i�2��V�[]W��i��ȫ��V������d46�.��VU�?\�G=��[��:$��dz���i�<��-�p�u�*]j#6D�H)�ꕫ��)�u��R���^ʚ��h#v��+�/8��r�Nj=QJ��>�N�gu�ѕ���4��={�Wk��ca7:MB�����}�������m�Tl���=�㛲�C���!�{����>�Q^k�H�6�m��T�&��Do�Z��앷M.�º��,��[�9�G�0��YI3��4��7l,�9w�Wx�mm����˫:�Z����UJ��+TN#w�Qrwm��h���h�LLu�wcMu�Bjrlʋ���S˖����N��%�U�w�0��v%]��ӌj6�n��[i%fɣL���ث��5>�8&tx�I�'��WSAjE&Q�R�rD������Y��﷽w�y��g�|ʂ����lX���Ʊdw���ƪj֥k*�YEb=YV1m�(���U��J�"������mD`���(��AP@b�("�;���mE�mA���.�����.���U�-���o%bԩݮ���UADDQX��A#�QN�q��mI�I�U-�m�ma�W9���`,UU��,Ek
ȺkmX��-;pdb�(��\�((��ZTDQt�4(n�(�#"�r٫F.5DU@�h���,:J���G���Q�mlC���,�*;oT*1E��AE��X"��V��uf9h�EL�(6�*0b������Z�b��UUV,EUb��{�O���N���wu��y���y42J�#�U�V��{i�v���-�9�u*Zzrg�~��)��jx�^�+��A�����L�!*��r�c�gWv�(��Pc*-2��ec�f�#�.�������S���m�Ռ�@õ�;�B�
:_ue=E6z�r:�ޫ�3��RP��w=e���5b<K�p��}����,q^�Y����6i�������8Ϥ�{(�y1L1���9*��36����Av$ʓn:����M�5��c�eH��Oa�Y���T�܈��<�{Z�  �p�5�1VD��EӀGc�=W�(��)���B�!ܸ����2�=�ޱ�d����"C��BZrOz��_U�j%�)��Y��4\M����Y�\�R�5*~8�����Ns�aֺ�*R�tU����t�b���\���:������x�BB���Gwf���Vj�gY���}�.����S�I�3��tʊ�P�_����V���=9��ε�R�,{hm�M��j�����>��;����W��ZۥP��)����J��n/�L�*2����7��S���RNB�vN���^G:��L�>����F���F�cUTq�{<]��7i��A��F���7qCLّٍ&vi3Ǖ�,!`B/Ʃ��Z���HΡ���ւE9���	3�0c�)\&��D+ ����bre<>����V?&a�񇹷����	v�꼏=�:���ADr�-�l6�b��9�״/q+6fYE�6�GJ&k����z��C�Z���])e� �j|x����_"wPd�2����,���}�Yq1���q��b�+L�5|#Ƹ����V\������Xvmq���1�ad	fyͲ�~�\��0��z�b1�}�|�cT�g�x2���Gp���W���GY٭�ńB��O���t�G���q�ڂ��f+�XG�J����c�XY�qp�,oqIb6�GTX�j]�);FhA��ym�Ց��\DԸ�X��I��c���ɞ�vq�Q��E����W;�a�洢�Շ�X'����L�����7�]VZE�|\���}�Q�Ok҆5��M�[1vǻ	�y"_�Ec�S�U�ގ��ڷ�"A��E���g�l�&�����1��'n]�{�yT�˧���F�6c�iK������rIR��P5�&&�5�� �j�\6�PΚƆs�2�۫��|�6� ����$����P����a��ն�E�3K�]v���2����*��6pE#�F�(ܣq
���{��ގE�݉�i�����(��$D�]lD��#y8t�'����=X��;��9���2=�d����T�#�=���F��nnej�Q�ӶBL����+�kTn��̽Ǒ[������m��Gl�LSW���]VE<��s�BL=�PR�h�4�z�\�v��p�̅����Quѱe�w��y�h�Ψ8��p�=}q����dtM�Y;�meI��sDF%�~\�wN�{ь�$���1���� ��A}���H�cr�m^�T se�4��fIB��ْAu�:Q�{�5�>�	�����Dz�Jo�w} �)K0��Gm�%��=
�]�w�kK�DO���(K"�Eظ4ܟf>"���-�-=���U���X�Ql��*sD�޲��ج��Fa�"��-�Z�F�y�F��STwt6�s�pӞ���3��,�c%���֑��뫮���=����G)�:�k�;�>�V�S���L���9�S���42:fM5i���br��儧�K��\�U���8r��t�iup1�H�5��̐_m�0�c��P9FS��L��ݡ>��*
���8�2]&>YvǂrZ��4�YN8+/SWn���K�ڋU%S����M�tgu@~��u��d䏆�P�N1���]�pِC.�53[��ڨ)U�u)���Ĩ�S�ewٞ��B���l'y��G�]�683ye�Eu$5�܃[hC��X�L��Kԩܰ��[�Iכ�����K	��3{���[C6ץ�<�|D�Uy�.�n�(�gy�z�܀�r�� �\dPw��5]@n��T�OE�re����������_�=���Ws,j�<Q)��9ֽ�(�V���Ƕ�KZ�����W�KTz���q�->ݩ�rzzRWy!�:Ւ�n��z��i_.;����f���-lP;�yC�e{��P������W��-���,#f�ޥ�Ϳ[g,�!eFTuhƪ�9;�e�%��Ev�(�tZ��[���J���;*I*�li?��Ki����v:YBҝ��!�uK7]����'_V��C�
'��ۀ�9�CA n����US�o��2�ƶ:3͖�E�����ܼ%Р�t�[�ׄ��j������KV�\>W<�+0�]rk�gOS�R�*�㫎*,��%-4Ms:�.��ݍ��-jH~�Ȕ�e_V>L�����}�Ξ�0x���*��s��EN���q��ؓ�s�M�`�%�ۅ�~�{k����O��B��j�@��OM^�{�z�֌�;C7,��]�k�˄w&�acX �i_����V�p0D�O7�:I��3o8�&Š��J�x�� ���]RO��7X�꜡x_���{���\ε�����|6�@(�r�ק0 )��J�5@T�Sbj���WL�i�ZyG`��RQ�7��n୥�!��m��7�b�\Κ���RՒ�̢~�-"�n3��QS���ڨ�/�ŵ�V�@K�.};<աĮ\��-�k�g��.�::,��f*�;�4���a�Z1�Y�j���������2�fs��ec��P�!uF!���o;���l5Ժ:��%�f�M6�Jg��V���Y��=3fyq �j�ϬyW�Xyq�\y�,�����[���J�ڷ��P`r���]AP��vs2^n�fߤ�E6�_w��;}Y=tNU�R�=��{]�}�Z=��dX����[^G��MB7\�qq�q.ń�(1��*�����W-�Z>��U,���ϗVSp��%qg;*!i��z��r��u���:����WlUx��V��|cF�wƷA����N����9�]gՕ2����`{$Df_r��`�./���"�棟G2%�j��O2w ����h�ݻ���θ�{!��F�m�4��2�ѡ�z87�8���F/8����Y���VڞI&��H@cJ�$��ёi׬;ԆrT3�ro�w:+S��0���
h�Gg,��pX�l�jo���n�;ڰV���Wa�h@�|gM�m���n��KeG2c������콨l���qY^h\q���iz�kq��4\E��~sn�gg�����e��Rnc��uk���i�ge��X��v͕�ٓNu�e�R�3HD�Q.,��ac(�T�݉n�7�B��+�c�3蚃�+��ɝ�&�,.���e���[m��7���j�ёN��c�����'f+۱��Ö�۟�\�e�>�%T�����5��bT[wF�=\��\�z:�=��P�A�zXns{���_=wR���F�ӎ��)�TVDOR��-�յ1,�@�/�Gx]x�)(e/�>a��c���Z���m��OGS������{����\W⺣�R<����~��
ʧ�n6�C�b��S1�[�a����6�E��M�W��v���7ӻP�@u�;e�"\Hw��9y�e���|�W�����bkQ�S�*z1dqbkS�!"�{�E��c�j���i@�V��ǽ��\���+~���FlX���lP��f�&�sn[���yJ�tl&�[���]M�Ek[,v��/�9	"��V�|E���v|C�JE��������y�(aʉ[�L��EVo�3�AbV�� {��r����ek��3Ӻ*���I<@۳n�goM���yn��rYtf�JvvM�\8T0��@���`�Jb�e	� ;7F���ch�c8k&FJ�2�^����0J:��X��d�Ó^��oM�.<r���2D��| �Z�����e�<0�ΔT�e��F���t�8m��7b�D�(*HS�[u;â�JۛLi����N�$�J�J��nLޙ�9f�M�F@Hf�v���ژX���ʰ�X@�t*��id������_-�
���+�9��l��ig��̿�;��Ҏ�}oj<�N=o�ci��.j��>���'2bJ��H'hi`�����:W[�V��R�Ώn�1��ɤ_�����x�8v0�}h����Ix�^�Y��
�w��e��a��m���t�p��� �*�{53�kp�HM}��k�y�6�WcTvg�/Gm��I$���ۭ:p����+2+<esu�;�. )��<�={8��9�oᡴ��9K�r�:�e��K��b��8��aR�s+ l֒[��](uP���f���*�,:�A���[��Xy^���+r��y�J�m���k��ZQ���̪��nc��F�i�+rL�p1��Ь�V.n����s2>'^Й0$�e����)P�m�{Z"��Ȱl�[[U����$��2�nB��]-��	�q@��ID���	T1���{�7��XQt:� ��̘��o�<�/"�\J�;nkbv�ޛBY����s�W �׋���gT��Aʰ�L��6tGS
�z�0U�W]~��L��ۋ7;4�K;�;�X�q�r��3	9Јj�SUA��W�[ϗ�w.Wcj
.ޤG[��b��n�+yO������$�Hb�y0��$�$��π�U�(��EDU���Օ1���F/"��Rڪ֊=��DS��*.�SMQDG����\e7h�+VĬVe�d�̥Q��ESvT^5�T�\[6��(*�ʈ#�Y��E.8EQX�qU��1]Ң�ōK*9h"��"� �*"1dV
��F(�
�*("5�`����
�(�)j�����t�٬�`��"���3%��Ģ�uh."���#Z�`�F�%]���U�"�c����8ы�i�e���ڬtʣmTb-J����EF!��Z��Aa�E�Pmff��R��*��m���R[b���|/��{�y��^r��T#Y#�i]���x�Z���!q���v.F:d��B�M��;ݎ��E�=��et��o��z��tb#ʖy�󫏴v�(!=/Ul��^�D"M��d�0ѓ�����p�����j�
E*����X�z,�!eFWFY�` �� U��G��,�[_�8�F��\���{�LE�G��2l�L�)�k�и|�yr�t��T�M��5���lsQf&���=5ޚWëx��͵i�o%6�F��v-E\r��p׉��ޝ+�.;��ற�{�e5��G�+�K�����S��!��1���ʜXCA�.2mg����r�z�#5dX��^ܨ{.؈1D�l�O{/r�b����q�7�@��[���jJ<l���<|��ތ�;W�����Y�'�0պ䁥I��`�ɷ�C�6�/B�"��e^D�1��M<�v�&�y��6nձ���g,��5q!ͮ����i'2i�qdʥ��aE��S8X��GZ�O�hx*��"�9�E�.;N9ᵴ"Щ�M���P�����4�bq���^-��4��O�^9�V�9
������ѽ���X�mw��0�m�3�E*��ݼ	�l6x'Ne�ym�ДTY�B!eF'����Kv�oN�.�$��S0�&�md]=��%�)4��N��z�m��$��&�����Q�r���Z����}�T�V�E�BA�C�Y]J͋�y[�7Ɠ�Y������5x���;=�Xq;T��2C��3p6�qS�+muuKDf��&�[���뜩�B�R��''h6�.��F��.��.�w	��V~�]Sn�}��\՜�5�j���-E�������v��^�;�i�������*�3�n�=J2�yPn�=�����^;ԕF4ǆ�NT�^RY�x&�@��e��g:��j�b��*P.�z�����n��=�'����h�q7��4�.�^J}S�3x�t�g�����mRd=�{�~�'��ѥ)�x<5�76.#���Z��s�vE�aK�ܷ@���eevzS�km#�K����D��	��@xH�W�fU����U�7ؗ������
}�N��ҀC⫰и��N�ͼ���%�����'��]�\�E���T�z~�x��y��:�Yb���|��`6J)�n��!bMhh׭N���)H�i����f<�$��>�G�v7��J�Q̥�id%ũ�.*�l��e�(W?P\���!K�#�C�\Nh|z8�l���q���v3s�3�܆2�L�Kpdd�t�����RDǗ�=pk��5�ʇ��]���u���;��8����ifZ�TuYZ[���d����S]���Y%]X9Q�.�7{��]Z��R>�#�x�Ώ�
�����Ҙ��>�ˉ�V����^�7.5�#�@�4�K��1��ry�)%��*��h_b�����j�*�s:Y�<4����;�����&Q��§<���M-t�]Zk/*����6�B�eң��7�A�h�R���B���P��s_e���Ϲ�W�9����u��܋$��&�:���tz �s��.�:@J�Ρ�a���r~����\��(û^*cF�n%mWM�;Ȥ뭚�<�$�o�����wq�UѪ٫��O6�^S�
��'\���rWӂ�xD��[��L�ʞ�Hׇ�@��1�i��2�ǖ���v�|������ 퇭�[��*�*��RF󹮰�]:'�@��D�2t�{�[4���Zɓ!��F(Ĭ���T�u�1�4�P��a<��혱Զ�V��i9�M���즟�k����j�G�^E0VZ1�[b�<d�7�8�v�,3H�2�Zj�7�W#OVu��gm9ʽ�K�=��E#�T[PӞ�VQ�b��8�z���q��'����-�7_g�r�(S�Q׵�,�r�&������⓷2���ߟ��󢃴�9PR��g(l�ä�<9�9ۊZ���v��Pܒ�!8;��t~��mlv*�jdb�������ER�������˃f�T���P��ql��/���f���=��Cr*�S�U���\�l\��I����};
;~AW�5ɘvճ��ig���y�W2�"lwae�9aX9���8m���D�eYI��^�v]�m_�|O�gs<{�/M��86�L:�q�Zf�6-XT�E_<wEދ7f��y.Lm��b�M\`��\/�y��H\:��+: @8+HK>��FNšx�\U$�{m�<]��i�+�pY]�U�.�k[��}�i����
=)C�ˆ,���n}$�e��
�g7%�щ�
̛9�*�cՊb�KKC�4'4�✧x����KaU����&��u�-Vp�����6IA&{s~�B���/#mE�\f���^��n�,�'�����VHjJ,��CA��떆���		tȬ�q={�Kb�n&���V�J���ГEd�Կ���&;~��ﷶo�ѓȫZ�&�'%�C؏�hз��k�-1JxƗ���&e���ږOvJtz_n�Y�Ƹ��G�QFb�s5��m�0��&��6n��GL�v��u�I�ٜ�e�X3��8�*�HΥ��\�yz���Y�I�e;E�rA�=�P����T9-?)�k4`�U�&��3�u���K`�+�qb�jI�0�)ݨ�%��8��fö��#S��I;(Lnk���Y�z]�d���)>c� �F���LK�<�n.b�c�aP35[�򣊷j�FH�&��λr����{?���e��3�u�����D
��_����Qx�k�;��O�b�`^��p���tz���uY��ߞQ�����.蓟�b��}��o����9�O�Up�����T�������h��>�5"`��Zk���~,u:5��-c}/j\�>��:�p/')�5����~�Elo�-D�R���Y��P23xarAsgbT��q�Y�
����pp�K�@��¹�����]�:Zex��U��5�/��`�^�Z�ˆ@�x��շ'w{pʥ�����j������l��j�>1�%R�f�w8i;�6{���WӕB^P?h���G�D��< jk�s5*��J��Z��G'V�+�$�W�Mҕw�>�[,@�����ږQ�I8�jXɠ\�/�UҬ
�ۖ�s�65�e��=��a��^���@Z9��/�QGi�s]�gU��6�Pa�Z��TQ��C[��l]��*����=+�3n��WRq]�K��M�l��K&]�n���g�'6V��ᰲ�p��r�0�\Lp�k(?/�E˓�G8�'{�E^Uus�dQ�O+ʦ�0�t�ƴ�^�	hۧmA��CA�t����Q��,{+$���Q�]j�4��yi�b��^�/��M`��EF�1HA�E՚�~Y�����_wt��j�^�2���h�l��/���A�c�T5��~�("Ls®���{&�l0k�<�J�0�=���5�t ܭ����Xb�wc��ߎӟ92#�ܹr$uA��~�h��*�^��[�ƍ;�4[��K�Q��Z�]&�|��Cc<x`�pL�i�8G�[g/�r���NK���G��nVR4��/yp��k?p��Y<Z�I~8W�w~�N��̭��+���%3r�1%�%��-�,w�J���V��ij���~����n�H0�I�s�#�u�K2ܑv�F���v�LQ3�91U���瀔��W?%j^����k|xK ���&�+I�nOO3ymu�|Ѓ�n
�kf|�2\-��$ ]��Z&��g����=�{5�C�kѾ��o�O�4=}��^O}ɖ�Q�(A+xg������P�=��=5nL�f����L5V�,��&;|����{3�Ui�ƺю��ix(|>���ND/���mT������ٳ^��������1��1}�YP0�G㕫y�j������Fؘ��Ǆ[ܰT'��
#�}/��/��3�/*����w��R���,4��^h\���dhB��x5lwY��oi�;U�:(��믈��Da���_1,����]E���i��5ޚgP9�W5��0}u#Z0p��>������QkZ�<�a�w��""2LLu��"�	H�����yx���*�����E�q2�5%��f+x��SΥ�k��8�$?��$$!����!
C����Ђ�;a<2톶�ElegT��:RTPO#le�i1m���������O���kq�8�4������,������5/����-@�z�9[&�f���~���粼�,} ̂��~�tUT�*�$��_�����C����z�ؓ��LT���Y���P�:|APL|��n�b u�i���(n����K���쳚�j@�U�L���Cm��Ѓ��*=�`�ӑ��W(��Fv�PΓ���� �*(� AP�dT*)���G;�&�g(Y�;�ld&�a��UA67��Ŀjhہ����}B�'H"=����D�[Y����G�U�ø� ����)�7�$���"�	nL��"��=m���8v��j+'���4u,�.B�uOoG"��oId�l���;�;i���^'���䠪�nzc|y�!�y,��g"�$�ߒ�D�� D�{PO��~�`�-�Br�bW����vT<��	�X2��( ���C�hЍ��0;c!P[62 ��.��SV���b`���YԴB���!�	2��Z�q@����*����'aߘ⠪�E}�P�&��f�8�z�v��u��6�5��:- yup��><#C�y��=���<�<�O��A_��%AU�;]-��4E��Y�P9x{�	�
�$��`�[h>��g���y{u&������odȆ��.ڔ (����� r�טZ��̇�����������ж޷m�PO���9�����72E7OUK�4��P�MN����y�2���`���f��B
�	�0/�=���c���7�st�AUA:G�ԛ��]�����epBʝ�{�K��A/@A�$��#�G'���"�(H8Lꭀ