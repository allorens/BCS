BZh91AY&SY����_�@qc���"� ����bB�>    ��,�5ISZ�5�Q)�Z�USH�5FIKL�D��U��(ҳQ��B�����h5kl�$�Tٵ����lҵlVL��]B��5�P���mhi�f�J �l��,ض�hK3e�T��kMMm�M�%��LbֳPeDCCZւ٬�F�f�U�xyޘ[b��kj�6���m�l��ڐ�����L�m�$��$�h�څV�e�6�+1�)�4�������[#e�m�#f����V�6m�#.M����k�@   �r�h�f����mY;�:��ft��(�-�d��j�r�Tm�j��R*���k�Z�¶�f��|�QOP�M6lg�tu�Ձ��   ��J ov.P�A���m�nt�݅A�V(h����
�t� 7aJsus�BTs�: H
��hPk>oz&�m�Z�lX�j6b�e�   ���hJ���v ���M:h:XT 5���@I��iT(P睽���Ox=Ǯڞ��U�W�����&��R�R��Ҙ��V�[(H-�   �����@�[m>x�m5JPx�����_>��/@
��}� �x;�zS���Q���ހ(�}�z�Ae���Gl�
�==�z���a������mKF�l��   n�|k��y�����F����#q�N��]�k���@^nP�)I�8�æ���wvҀ�Q�U��.ک
'vۺh^��[A�mYMY��i��T�� �����ݛpҀ۵\t �g�tҀ�u]�Q%���`���9��A[J�T����(t:����v����i-�Y���P4��o� '*�(E/:�@�j��F��Nt�:h*�ú@� �:�(R����u:5l��PP��n G��X�Uj�[f���U2,,)_  ��4=U�kp��8PA� 9�n �tw  Z�8 e

�EԱր��M[6��[a��"@ kQ�  :}T�u�P�X j��4����j�U1@�r�4��pZ��E6��P��=klYV�&fͦY6�٭�  k���@�.�]�\ �0��q�t �� � �W  .��P
|   R 50T�T`F  &��� ��i�RU( �h  �@ S�2�)  �    ��
j�P d     "�2$AS���FCCF�I꒨M?�Q$���4  ���y�_��1����=-����ͦ�;�d��W����3X�D��n؝�@ ~ (�( �� U�~����� _h~�_��%�_�������UUm������UU��e4�_�-�ֶߟ�w�?����m~m��m��ʷ����˖��/�ͩ�W����k���-��k�ھ��ٵ~sk��}���Z�V����Z�+_ek�ھ�k��n�}�����k_��}�����m_f��V���f��}��ٵ}�W�6��j�-��Z�-_�����6�ٵ_ek��-_�Z��W�U�W���ھ�Wٵ}���U�m_f��ʯ����/e��U�m��Wٶ�6���o�5���j�~�ڭ��Z�Ͷ߼�V߼�V��յ��Z�٪��mU���o����r�m}�m[�֫}��km}�ڷ�U[��V�6�k�m}�ڷ�j��涭�m��[o����6���km}���٪��6ַ�V�}���ٶվͭ[��i�k_em��Z��f���-Z�ekm�Z���mm�kmo����j־ʪ��Z�쭵�ʭWٶ��ej��[}����6��j���m��+j�f����[k��m}�mk�֭}�Z�٫�}���m�U}�_e��5_f��}�o����}�߬��־͵�Z����5_f��U}�Wٵ}�ߜ�춾�k��_e��U�Ym}�����-{5}�����j��W�j�5_e�����m}�ݛ}�o�o�����5���??�/¾�m��mq��ټݤT���-�5ܬ-Q�wr����R��Gd��L��O>J�ڳ�ơ��y�[շEb[�����q��[��p��b�ں/�1��#��x�/0g���l�.�k�yk��ʵ["#mu�V����@@L�Tb�eH�0�w�`m�@����Нd�hfv�q1N��--�"��&�y���XY
̚�oa5�l��	d�I��@E��`Sq5�Z�a�6�-���`4#vz��׹�qyx���*��ז��b��m�CC��c�θ� ���!_��y�nC�k$��4��T.�juv��uHf���{i��Ե�nS$FQ�6ą�V�����M�z��֚���e12��`�	b�[�5]hǋ/2ҺPR�1�\m�[��ʆ�a�ߐ�Z�:b0��$֠ݗۺ��2o.'��V�F���!�HR2�L�����uyWM���e �<{[r,kXƪ��n�^T:e�滅��@���c	��ú������%�&�u5�b"�%��"��Ԅ�)G��m0�ֻǙ����������uld�a��?��a�.�U��e-dLJ*=��*1�X3$@d������F��,ҕ�ݻ����>2�KRG���92�ܲ���3M�J�&��n�L��*l�n7BÇ$�fiq�Z�5�emu�Ϊ!����fb�����"�5eM!�6X���C�e;}I �F���������e'��s]�[�&�֍L���(��¶F����]R�*F
�'-�r��2�R�R�k�F�C�V�A�Cu S+j���"�h�˗��@�5�s5��#�������
��E^3�S@Hj˔�`��A�U��k5��n�̴�g/(@ؽpT��Nd����͉�3���V��ɺ�i��Y��7�)�;��N�Y�ך��z�jnz�yn`�	\`��\�@�-��H�1'5�t�GHce"�����O���2�V[Bؤ(��lïn����8���a�3�$L�[ihYx�<%�G*�㗔��X���6&HU���Mk��4Hٔ�G�^�-AS"?�]��ֈ�R�cY��Uǃ7qǴ�*Le*W{�u��_|��0���O�t��׹x�:�q���M-�C�cͥ0#a2��}Ċ߅�n����y�u�p��H�������6+�
X2 cYۚ�V��6�;T�VУ.��ڬM̳+iS�U7�Ȗ�x#9��Q��}�v���2�Xǂ�-�A�*�Y�j��9��ZmlIҥ#1��Q�S眎$ ;,�8Q����mNn�F����KP�� x�m^a���X�Dn�5�Hʳ�C$�v&�(\P�ջ5�cefڷ6��~t�Z򛥗u���Rf#5��ذ|��k6:3r�4�fǕ(�����1�i�5�V�����S*� ��T¥��J�`ې+��T�d�&Sp�(�AVA ��?;�/K�1��C�&����:�0���u�$�f��1)-C#��[ V�``Ji�d|�'���1ӬKo�r�� 8�	�9�i[{�=��beA��f�����$�g~jw��`l4�+x�;y�bL�V�����ݬ$f�d�h�X�u�cv~O�� ��c{11��%�&֊�i BK-��N�j�7�!���u����퓁�@k�pa��b^�e����U�R�2jRŬK#���nFn�C(f���n�\w+�����;ڊ5F�ݦ��]2 ђ�ז�ۘ�"f����iږ��l�4��`׹l�j�2���E������";%Y�Ѹ�Vn�fd)U�0=+�t�F�.I�t�65�, ����Р���ǗER:�:�9Y���6i�bbw��i�mbI�Drᦞ�K)�b�3,�2S�*9�0S�I�M�hCH-z�@n��DGy.f�b�_;gK�j�%����z��m�g&��Mն��*��L<��6�����(�T�8q�R�V�궛���� DѐM�Vҽ˱X�{�hVb�٫Z]@�=��F,3�2�l��&�q�#�:�HA�%6�x�M))lŁV�L�a�ْh�1�6��e#1�)E]؎�Z����#��P�9V�u%���/�å�t��nQ)��K2暶saX�k�O�[͠�5�6�'�r�q����)�&�ݺB�[�����ԇ���q3X؛9�m�E�W�����K�F��ِ�5��:�,����ͽ��oU�bUn&F�^[�+]����یV�8*��6�Ӷ6��V���Yn��uQ�i�q�Y���H�[�3������W"�tYz�m�آ�*�u.^54XAS�5J
;�:��/$k-�u�|Jn	[X�VڣO&�!�	/.���S�QiO	�+_�7hXU�41��-T;�/Em=o"س`op6��4�E{�.�షdiJ�����=���w���	1�^d ��9�X��|�e�7�ԏ�դ��[�%d���ݗ�F�M�9��b)�6L�D�j��^��4
5���z��cN��h���&�1^��	s&fU�C���K�S4�ࢨSh�l�vo�d��]�ˆ=ɴlA�h��T%�6��n�[m<D�K:��Y��F�u�^���-6�.�5��b�|�v�'�7�7&�a44��c7LYl�6�����N�1�=���� �m�KQI�ê��h�w,ēƪL׃V�VV�Dj�*X2���Ty�x�.�b�c���Y�d3]�w	�Ӑ)���,�0T#��9�^���*�;0n�>=���r|9�s��Ü���k	n�q�f�I�y�*�-�xF��2��}};�O��{L*�o7���H��	yp��{z�%
H��� ��9��d'n�L��,c�>�y�ٺ�ђ��Y�܂�ƈ���C.�dݷw��ͣ�kLD��f���$x��>x8����:�U`Z��5=a�3As5�j!�#m�ÔV*���E���Zn잫=xFf&^���|���ը�/#al�OR�#�ᧈ+��±j�X��ʛTi�6���D;�.��:ډKAm���F�m�WG,�7m��/�9���4��IF[x���5�2�ѬVY��tv�^�����y[cs6��7`l�KE����L�ʷ��X�3*�]$.!d�oH
����P<QnX�!��;n��lՒ�/B�fk(�4ȫw`����w�Xئn,Kk"�Chڇis�۩mGf-�|�-&���5w� ����o;'V(��"7:���Vf��e-�o5�`g[��	t�n�γ�GuXN�E�+o�/�4)
��Z�mY�y��v�׶���\N���]N�V^پ�X�_�k,�kk��Yr��/1-۱{��]�Н͵�c0��kR�-�գ���:X�g+-�p�9��ֱ�5�Xvʤ564�,���x��H�Q���t�tCRᱦi�Y�3c#Qj
\NM�ju	���Y�bb��3yuq����{�5�l��B�J�ݢ㔞�b?m^fU���Z*�������x�ڶ�����*����{�+��GN��@�WMi����'�����n�����U�K�/�x�\i�w+c��]CZ�������,i�v�,���Fd��{Qh7Y�kQ$��1eɕ���[hw-��5#�b�6�Zv�L�P�cZ���(�}��Aˡ�Z�f\��
�)0����� ��<
 �&S�E���Gj�X4+"y�o.l��̰Kj嫘V�2H��T��m L�`<['ί��VHm����dK�A�Y�hV�٥V��p�Ź��[�1(����yJ���)b �6IhI����'{e�M�h4^��jE1
��
jSb��pDwT�wU��\J,8�7
Ř����&}��0n2���b�7�Zuy������ͩ{yeZL�,z��y�S��qC���I,�#7�Ʌ�vE�2����YȽ�Z���o5D%�fUϮ�C���T��&�e�i8s,��C.���B���+ac�b�f��Q�l� 	)��-z�9q�m7�H��6�-�L�n���F����[M�5xa4��+	?_k���[CS����I�*T��7A(E�l��B:�.nY�66�V��R�j�Z!<ۦ̩�%`Fbm�I�A����n�
�'��0t�N+�Q!O.9�(�_��V˕��Õ� D�b���@XCe�Cc��.�Ak�}6���oE��F!��5�n�"��ͥ�XR��-���7ss~��Қ�^ F����1�Tn�MB��m��^��ow��m�!�dcnk��9z����&dY���v���rCx��s��((cz��(e�.�bN��L(�j�1-�hm��*�[�
��>��.m]TJ|�I{["ۍlX6�h�䤤ܨ�a4����M#u�F�¥<z4��s�8�b�5�C̋rY�z�:%�S&�⩎����P�R<$J�Up������J�V��5p�Ki,xԄ50\���V��3�*]���n9u��Kt�fJ�%�VBh��n3&Y1HkV���J�Ҵ^~JK(�xC	;�/J�7�[u�f��D��2�`L��(��ǳd��zcZ`��:�"UՍk]K�*j��:th�IWj�I����,^	�^#C3b��M�Gd��CkvN?�I�x���ts8�%�х��+e��X�W��4�j�ɓ 1a�YXY������Dd�L�ֳ�^Vm��^:57��(XSqL[��,��eE%�nk��Fn^D�	z�x�Vr{�4��`�N�G�%|1��D���T/�!���Tue��9��/*�XW�vsoM�S�̃P��L�X�k[6�S�t�Z�4;�*ʬ<U?�5Zq��:̂�J�
!m��-��c�H� Cx�bk�
�IM�+7wX������v���p�����Tn��7DPJ�ݏ�2��m��u3f�$�;��D,+�ڧ�f�S�LnR�͚�<aU��[-һw{�5�h�͛j��1�{F2v�36�B��x�oC�u*۲G��E�h�������5G4;oq�՛�%mhl�CQri����a�R݊JmeobBh�r���:lh�����	K�r��
W��Kh�����&�%��,��S��aذA
��=e�R\r+:eBj�Â�ǲ��l�������2`f�ed;o)5
��
��1�P��v�7�a�l�d)NAB���Qo0BB�w�4����$����Z2�խ���?2-N���D�M�'������+�v��JduE+�Q=d�XYǲ~�Y�"���5[5m˨e*a��P^��E^ix.�6��d�ѦH�Ę�L��q�!k^�T̙H����R'!c)f�®�.��D�=�6�יp�	���طt�8P���k��Vɰv�,&2�AZ��^��$�4NꢈRʬݎܙ�Z����Nl��������`[&^�3`�a�uW1�d�I�#|��C�����]�aepڷC�>oT��Ku�*c�AY�٠"��k�nPm����uj����P���Ђ�(�^\ڵrne��d��MX�[Vs�sޣkuWv�K����]
y,�Vf��U�sr�����CS$�Hf�:vԔn{��׻!�
�ie��,�jR��Tl�TœAض^�#Ʊ7����m�ݱ[i�:N�A������%���ɏ.WSg$̦�22hm�R|D�;I�v�bJ)���1m�%hbb��Mm1��\�n�ڡ��vV��VQ�2�͵��`PƝb�!x�7����j�<���Ŷ�EXhfZQÊ��r�')`�vZ�Lsr��E�D2�6�l�i��h�k^��{��5x�^���[؝lߕ\B�e�N6�+�0�b��<)�ѻ�5M��t�m�Mט�7 #*�c�{�"�.��Mn-jD'�1����
��wpgTe-�.��j"��ܨ�SJѭ�Ak�t�-��f;�E*{`��aҀǚ�偎�ZA�{v���d3(b���-�U-����V+\�Ja�N��ɰj՛-��]��[ݷ�L�V&�հ�m�3J�;��&�f���*HpӢ�T�;��ֻT��L�Z��Wځ�Z���O����ޭU��W��^�(�S�_n��kd��w���B�P����䬱���uR�V(��A%I��̼,��h�Th��u����X����5���-�@���� ˬ5tH��E
2
B#0n���]�.�����~�ù��K�K�t��d�T���F*�2��I��Y���Z�TM]sj�wV>�3�z�ǻx�
�4edF��2���n[[D�#�m`����wZ1�+s>�'����pv���tU��I�������b�J�M��:�Wp�9[Z�~d�TR�Ar�'J�PAz&���hkZ[C�������3;uC-�E<��9��n��r���	o��M��V[�}���9m�5�	E}�k�ʑ��;�k�v%�Z{��`���r����d�v("4���F��5[��ӒV�H�8�dЍ!��'�U��X�4��.l�kH�-��]�B5{aB�.� �P��X���J102��%=@ȰB�����HZn��X7L�QDb9)����1��T�F�M�pI��ܽLLm�M%�=~��(ʲ��7K�Y]$q�"O��WGZ��W�(2�p��;!U��`(Z��ssC`�G����O�嶐:��z�/Uˡ7t7_FI6(����+	�|l��д�ӑ��Xǃ�)��Z0*^���<t����8*V�GWH:�ti�i�SE��][ �4e[b��74�v�34�=��.�[N*٢)j�@cj��a�VP�C�T�L�h8��6>I����J�L4h !��"?�Ͽ����O�����㮜i1xj��z�^��{�3;��"��J��vi����v:Z�0DO�����ؚZa��sN᜖bhͻ�m�3[{.�����y �!ƇM�U����3Nʺ}�E�澆����@��1��Ê�RkalX�4bv�@�ce��J�4ػ쬊��X��H�Q�}4���B99`r����ٝ>��Ff��"�ri�}|����v^ʭ�0m��U�|NG�Av��[y��J�;:vc�M�.�f��b(� ŋ1���ǟ"f�ᰟ��C���a������o\C����O�:�éT�� wm
�q_i�OU�J�IyR1c,��<�����M2�L��,?���fV�!U�~�q@x���F���U1YE��/i`�fzN�!�[]�}!'#oM�9���5y�=�5W�N�c�B�h�f��1�t�� ����pA��.��x���;�R�$��sE*E�ӚR�с�݁A�kT�F,Ӵlr�s)8ƕ�xѺ��7&��Mf�O2���(^n}}�V�M��_ؠZyf\��%ӒTS�g��C2����_n�0�W�ST����ګ7�ۂ]g&ցHM7Î�ۂV�;�5<�	�����ݍ&*��l��%�q9b��&��W�4�ZE�\���*AB�m`%B�vH��UqWq�Xj��6���)�ݮ�z]`SQ�ޞ��,��lSX4��v�<'���5)n=7����L���ܹ��>�m�ѱ�������b�j���
���z�u܁G��d�:Ak2����;lfW��PC�1و�Z���'u�1�PUvu���O���J�o����\ͥCz�V�W$���w�c+NJr�,WWFR�̖���Z�&Y�x�BM���ú^L"�2M��e#�$�Xј*�c�z���	�9�u�H��7�DSB��"TR��Jǈ����G��X�lϫ���a�eZ��hm���D6����h��(�-ź*u�0��]��^l]�"\0L�3d#tt��>3�79%X��t�MQ	�pSp������ɽ2��f^ �(�.��n�m�/�`�%dNP���V�X���s{��h�r$�r�J
� P���&[��X��]��խ%�fV� ���I�83\o�T��q��0�5y��͆`�/��!�{���$��ڵg���G�T���6QP^�mk���,�m�N��K �݊Xoi]���k޽0蠓"�np�:P�R��FV,�􋲝�K�����+GBh=�P�Zx�:��O��GGe��i�t���tg�=��:�$:�*#-�uބ\��>d�x�s��N�� �.�Tݛu5�֭�9�w>����nl=�45�3%����Ąn�+a��� ��%x��W�km���N��2^�#��+^LdӍ`}�+6̇�m�����b{z6�Y��ޤ%��eԤ�[�囧�I�7\6o�`%�j�{;�e�m̹7�6�j��;������6�9[7S�2L]@�(��V����s�rMR��<{0ꖫ.dZ���k%���wtf�M"s^-q{�w� �_J�a������]�,bQ̃���ZM۶Ļ��Pg��̳c�; �4����g-�1:�]��@>�R9.\=4����4�v>��:�4%�f�8�,Wpmt,��{t��[
Nm�9��U�(���\��P��7{�٦7�n�Z���U�L�wWZu6
)�́�Yo���;���:�;:�7�tvD^����ee���1�ލd�b[�%/�]:Ӑe.�z�v�W)e��XӼ:!�M[�h#�_1��MM����,,��K*����͜�
�9bk��gQO�.3k�wJ�&o�Sb�]�����^a�����)�� �{Ce�M�L�"����G��+.��p]J�t�2:wC1"o�+GUw�[W{�}��T��	�՘
YN�- ��%#w��]o�[���.�H0��{�kP�.��:8���˳�,�[xgN
L��Cm����y��o@�ۧj�?D����_X.���W�0lޫ��'B�r�n��q���3����j�@(��!��A�t"��6V[�/���F����{r��Ji�o6�c�x�9��
�WE�I�����۸��|�� ]M)/�"���H��Fػ�nI�yB^�^ջ�s�2�;iL���nKui��K�U5	�'7�.(ݚ).�p>;ى��M]�-�P�;�)����wX��<3�k�Q����K�-�Tk�k ��P=�W�J��Cl�ٖȎ
����i��M��5WV�l����V��t:�����v���C(�N�喘`�R�T��r�C��3n
k�.+Cd���*>����.���%V	��Z?`�Y����t�76�V&A�:��=��em��v�j�/�r��5:b�Ɛw>�������Z-�K�-�l=�i0l���2bPA�����!
���w�j�5%�wX�/�p�#�����6�������ϑ@��ʚ��\����\��f�NmT<0�p�R��"���?u'Q]�m�j#��Vw=�ZrR��5
i�8{�G0f�V�3��tAF bz#�
���j��ɚ9�%Z���;�B�b�A����&[�KY}�;���׉&f��^<ݕ���V��1�u�kf� �ݧx��Z���;���#��k��S�J׻V�&���)��Ю�����ܘ���t��I�}�q�`uoN����o���P���)LKW�ToY<{�Փ[J�ur���#���/ �+�����I�'C`r�����F����e8�ʽj+���Y�w᱖v��`��S��	�k�}tu��UGKke,�Ie�6E�\�Y05�+L�7@˹ǣ��sc�gNJ��E��omn��R��+�kj�*�d%�E���&�RD1��ccn���v�u�/;ERY)i�!ˬ���w���v��#.�����W\��I���K�+�l���w�`'�+�݅N�eF��5���y�9�bê
{Yk�a�'����V��oup�Ýy���Cr��#�%Kk9�����ܒ4L=�:��!�]|nH�qvfH�%���{���]�3���«���F<��h�!&]�YE^`%\���\��7�c<���"�S��$nv��#�L��m.@��1�+*�?̊5�BiקHm�{R$�v��Zym�S"��qV�0o�	���Ǫt�\Y�� ��˄��g�.���.S���3�K	�N`��z�m��$�3�ν�|C<������}*�n]!ooGI2��F��v��i���G�sl�/����`y�}�){M��bk(*�w9]�Iq��"�%v3���خUl��5f�,�yOۮ�Cv1+z�ˮ`����1��U�Ӄ!�	 ��8k�arڳe_Ŏ��һM�K�y���܉� �n���{I,�.��V��YśWB�.��ݒ��b��W�p[��J��1V�gMG�goV�	�d�}̓�y��jN]Xv�ó){�g0��>�t�hU�G$4YF�f��B2q3'J.��;&��v�.�ZR
�8>{-wm�͸M�'��$R��9Ԣ��M\�i������>���of�S@��~s�̠�pJ��������m�ؓe)Yx�lKA5��I���A*���۰��pr!'���/`{Y��/]��pk�)y#&CyR��#���왪c�t��ޣm�����a�)@��9��f@*��0�ս�������SB#;�������å�I���:����FtkqV�K@w^�f�!�Ş�-7����"&3��x��}b&wD��&Rwc�P�;�+aWl5�G{�!����b!�de�n\.�}�F�m$�Y��ZX>α�T<`ɲ��6�����&q���I�e�
wb���������XBʦw����Fv�O��vMlUU��� �K�K�wt#7�I��ۢʚ��D�ʓ0�/Y���:��/1Vк�o���>����.\�X��涮]�aҗ�F��)�y���
n��rr�Fs#oV:oUe�0�3:���z���2f[�%	�u�UL����ý��2�8zk�fE�赹\e�n^�c��{�3����FM{|�/�ˢ1�09�#n.�;fn���t�CGc)��}p>���� ��V-F8���q<id��@�ξ�2���F�ක�Y7���,@�-VP�S/X���v�L$b�]ǎ�7uO��eL��'Y.�'a�v�8�m:��������b�T�W!�zpW]=��=N����X3E�j��C�l-�c���бR���̻��sf�zƭ�C���PXy��%�J�&e�(\[X��8㬘��/21/:��P��V]L��s�epw��[	���⭊̾ʖ��jglvw��Hˌ���m^���Z��̭Y�u<X�Cf"!��2���8��<�O�$o���T��9Z-���Y�������wj�J<لT�*���F�J��f*m�eqR|4�L<[Z�W�����"<;�1ˆT��+w���9K���� H�Y�,͝e���|�<F��׉��ᘀ��tZF3�k%�F��~a!��?=Dj"5ń��u��%G���olOn���#�$� y���b�N�.�YrZ)�����4��EL����d��$-�-�\��u��!����ʒe��w:���1
=$:p���#^uʦHxU`:����_5�P�uÓ���\��3l�ېET%RDҶ�7U�d�,ڜ'v\W��2�SĢ��ZuVX��'p�:�W��qa��λ�Mj�%.�Hf�n[J�I�;�0��R#����1΂E�����M�|�U�mޝX���K���*���S�:�I���e<�NQ���X���u�Z|n^*{tU����L���J�1���ro�*�e�af���Ԭ�����噄CYw��G]qX�Е��^	��Rj�lS���!� r�arX�̬�po@����AC��H�V/j����c��6h��_:{SaToM����87��{1��"���̜Pd�AC�Ϋ'�0�����9�Ț;m��y��,��efjtۺ�p�QSKaK��\��7iI���rqur�����e�($��f�Lj0�����c�1�.!R7���i���Ƀgf�ϣUw��4�]'@�"�B�b<�*�WH�_��]&��ٻ	|iGe7O�V��>q�L�o,��m�f�(����-�<�Ɋ�m�ŷ8]X�W_@���B�*s�#(���6nݛY�cJd3-����@qb>Ua�g��A\�k�M�9"���:��=%P���ę����NA:n"�"0��罄���4�pk�%��a뜯04�%�J�r�+����ו��,m�ȥsH.g�����NU`���T�>���g+�`��Z�+ŷK����vv��yi*6jUnG�mA)�����;�}��.�n��N}�ԥD��[En��|+d��EAջ�=�w3�l�H;��DO�{|���7OD,1^$	t�s��*i(S��<lt�gXo7A}�3�l�4���Goj��r�E2[�<z�pM�V��iq���sDA�}�I��*�݇i��Rk��]�m��VkP��\f�O��42��ƶs�a	bEw��:Km�%�u�)�->C��na��m̙�F]�;�؃�m��	�$�y�Bu�eT��cu�vV�1�4��C�eqQ3G�b�q��liSw��-=M4;>��Y����Cρ:vR�<��͎�w����$\�5ӷ*�X��Sp+<�
	4�κ�t	֗)X���-�.��pH�Y\�ݴz\�LZЮ>s;�����G��Qn��+�h��ڊ��"D:��*��Z�+�t�ul�2��d'�}�W�pF�9��xVM�pɸk���]\��֓�.�}�34|{ �A�Rf�j��;T��>�ޜ�.Y��cӴu>˱}/qz��街Dn@7�"Jx������b��ol�7��6����͈�ۓ�U;s���w��CՑ޴]���j>�Y�	�@�6�'|Ôa��8���U�60���v��;U�6������5�2����2�YZ�2�GWu=0�"���v��1��%�6�Wj��:��Ҁw�~+i3l`������_=�Օ*gA�黷�����TJ�+_ ��"t�Y�yU#}ٝ��0s�I�0�I撝űţD�S%��n@�"��/
�,������ۦü[�Gx�D&Ҿ�;���������2�#rI���м�ut���-�Jk@6x�X$�t�hK�gR��L��+I�4u�V���Y6JYY��KI�����uJ����!���$����2om3�gv��g�^a�}0�5DpȻy*�A��v;u��9ّҵd���Ϗ1D�\�hCR��}���!���]ƞX9�l�b�m@�q���.���λ5�>:ɹ�Z�*Wd����Q�%�Խ����	V����q}w����u�݂�Ͱ@�/Nkm'4Vj��əSV��W1G��7���Uq�y��f3Ov�6��rn�{F��>c�0�XvG�"8����W�s�XM���X�ϰ&㫉�Hٱ������j���Yx�w#�*��{zT��jʸ^�v���
� ��f�#��+�Eř{�Z��2P�;�n�	ֆ�Z�㽮�by�3��\�������M�%�w#��aU�w:[Ĳ1۳�Cx]�zn\E�bt�3�8đ���m��M��<��u&�DB�)�N+���	�+����o��K��[��y��;~������*�j*�J+��d����כcm�_�9������b[�j�oe�q�&��
�LF�cz�p��T_/���Q @4s�u��B���}~M�������������<{b<����D��F�N�x��N�9���X�����q���w�7W���l�h�3	�S�H�Y�E�&r�
�+j�� ��Gb%N�XNo'M��X����������\ޔ�sm����m-n����q�-��{")�d,���CO�3���V�[O�+b���fJ|�f�9R�|`�r-���>�H���յ�+��%�.r�t�=��-ˇEmK&r�Ю�r��3���Z~�ۊ�M��B��`5�}
��m��6�J�8�@����ᒘ�h�Vet6_,�������J��Wbt�o �FM�:p^��ʒ���9�`ܧ�Q�줱	�'\��ٻ���XO��l(�ĳj�Ը�؅t��]����ʾ)�@_fܩ3�*<��뢤_
˽��$���-����6�����J^����02�F�7���W��?#X��t��qB��|�:쪁I2�ڱ��.7/�k�1��c,�G6D_�Jb�Wu$��(b�^S2��������Tn�\��7��(����r\�G�:��rRZ�{�F�k��K��ud���JQ��5�R�&��3s���;RS�|_u�g�<:��)lw*h8F����v|NZ��P�!��b;�����tV��B*��b���c2kKIb��0�4_���Xqe���b�B�9(*s9��c�_i/r7Na���ʹ�c�jf�b_�䥪�r�0�*8�zQt�x���d�:�B�=:���`�/��w_Z�@�m�4���z��*:��j�U�F��ҍc���߲���M�{*�ךWu[]�l�R�3od�I憷&U�������Π���t��7�8qz�f�;��<r�ހ�,U�xU}(�M�&����Wz���p�� ;哫J?Q>6�|V2ɑz�K���N�o)��E�\b�cc&���ײm*�Ah4����k�rĆ��<�r�)\��l�\-���i^۩/�T,�K��-��4$�bO���-3/���'	gC|���|��Y����[�ײ�@vf��ed#
��Cq�3n�7�e����p%Ψ!������2oJ���jf�v�N�O��ћ���p�v�1=`���弽zw��SX��:%��;WG{��l��s�aM��v����C8b�u����H�=��&��(񮗂��16	YC�;�f;�Kco�䶛��/J�#.�|�1��2�໺���^>�r�*�]�r[��v��E�q�I3����Sv��S�f��*DMnX��f��P7�z���h%�lE[�$�c���J��|@�rk:���P��˷���Q<���C{����ǅD���߻k_^�mΣD0�`�P�'p0^~��J5Q铔c�}r�tuت}�.޹a�H^;w��/6�V �4���ŪL�侔oe�ۓo���-=K��`��6�dj�Ƌ�Z��Xz�����DeX�ӈɳh��_,�[dBXʱ3�L��Ħ������;�Z�W�r�c3{[�f�)l;�� ����֐n�8��a[;$���-��[������� y*�X�[��t2�	�0"F��@�S���f����.�Q��ඹ��Ǳ�A8q8�X�o�]�6�f<�XSI5ƔxL7(p��0dR���p��*��h]ÑҀU��I��twg)�T��F��W,��5;ܜ;p5_��'���Qe.y�����:��{�{�"wqZ��ܴ�%O!�#��2:�ܽSBL�*�p8��a�Vͣ)�7�3"Zֲa�o�� �Uά������Oz��&�n��SJ�Yxʕ��)����L<�3�[��2/j밚kv�@ш`Z���i��G�YM-�g��I�u#{�(ਭ+��G{���D3j�=�c�ɺ�P�:�x-���ά�o!�>�S�	�q���"�dP50��9��K��R�[#}w:����um�l�muis���,���P��wqahlLa��ˣ5H0��|��]�Y�roj��	��N��a}�ռ#�,m�jq�u$�o�d����x!��ړ�$
���6��;l�W���6y���ɒ���.���7����D�P�Ϸz�w]f�h�/NT� ɯh�][q^$�[.��Y�\��a��.�l�J�cō�4֍�5;��-���ڌ�X����f
G���L%,%��q����h���uuW΄FNfN�9�{��2�f�y��I'�kc}N�������v��Ğ6�=����X/@S�l����5���ggNk�YA�\RـK5����X�+��gvj�	��h���v�ַ`0�3ף���. N5��i`� 4����NZU��m�sA��-�k�!jgĭʑ���0vA��n�a2�w_Rg$ŧf4��Ո}�ܛ�g�q�qS�ݝ&�i�6���-ͫ/�49��Kl�m�s.Dk�|���k��VF;.*�����}����UtuS^:ͤ�މ1&�J�Xv7j̛��"f>������Ӛ���4�{��(h�oR|D�+;��f���'u�e	� @r6h��ъ�)�v�a	dZV�Mb������;m!��Ef�C���ks_M���EnŁi�O�oB�ia�)�9�r��A˕�1�`M@
��Te�PM�(��|� �&,�]���L��pE;ޫw"FS�eeNծ�z���b۴0A7S�� D��yϕ�1A�%��HhT�ѱ$s�*ݎ���Za��j�^�;���d�!���_,-/���T*
�l��JI����k�Yy���JCt�.�1�E��![]���44L�\��W��S�q����n}x��[��*y�{��,�UFq@_2��_�(�W� (�z���}X+�
������K`V��2sF�h���,�O�
��k�TG�l��:U��z���w4�&�>"�k��削;�T}�����r�gL�w�`od<����.ۅ�]S(��"ԇ�h����̠�)ǹڭ����g88�%��$���(F�;�hj�#�0I#���6#�8��	�n��ڢV�Ք�T�[���s9CK0�t����2d�7.Ѿ�,Qtg^�{w�>�@���ݻ����o������4�ʭ=2�p���dl9!�oYɽ[������l����zHW��J�4s�a-�����?���9&48bm��P�ǧl��fT�l;��֗��gȩ��ˢ�f���z:��gu�su��ʁ�[�|�����^5ojy��Z�{u�.��B���8>.u�!�s��K����{R�0�%����n�$��8�w(:#�K��a�g�����{[H�Qux�%F[�a��1�ǔOC}���f��Ƴˣq�6"�����b$ݰ������6�K��2��#RU��\��`�lb4$m���P��u(�Ld�`�d2r^6a����Sw6����(�]�L���k�#��d{��m�wQ��3�jN��]6���+�\���XKq�N��b�;81ױ��r�F�����wp����3U#�!ޕr"��Y�"ݣofn�'�����t���-i�*���*9���l}�b��s�qs��N�]vQ\��z��I6���~XN��J�]Vi�x�:�=s6LruCͷ����Z��� �:8:v�m�4�BR�����>�t/��e���+����:ɤva��(�Vl�C�I�L�u��zrA�CW�Y�S�<C�:���kJؒ���l�U��rKL���P�.�6�� �.���ry��6�[V_��#��ۻ/B0)hQ��0�c�����{}le��NG[��[�c]G��T�r����x7�cikm���a�'"/l�֟K�ˣ��%hkZ�Ŵ�b�	���*���7Kz��B�N��V�n�X6/����e��UP���:�ڙ�Cw-˩�*f٤	"�<f��Xy�뷈c�7�Ӕ�s�3/�q�Ӏ� �w+���Q��s/F�9\�@j{R�V����ǏZ��ټ\-������÷ �P)�.���л�g4�gm�[�"���J��_!��9���a�ש�h�B��E*;�=i�
��gEa�#���H�q�3�T]ж���l�km���]M���ǈK}&�Nm�G��Yy�ܬ-�<�������m�'�Z6�H*��V��<��ҵ����j�X���AīA7U�|�T��4B%���\��QaՄ��,K[��{7����]�)��T���7F��}p�۹�/j�x c�;�Y\19�����l�gI���P�2��
�C��m����u,�@���W����eǭ�_XV�'G0�[Q��ڢ��O��/LM���9�@g_f��A͋�����6+W-�v 1��gx�h��/s�ҷ�g��w��e>A �����G Ӌ��Ձ�ݩ��f�JN�Y]Ȋ#��'@���Gr|.�#���&J3�^���C��Qz��k�S��=��E�+K���Ͷ��k��1|���/�_qru��պ��PU�t)���XC��K���N�`Ī�� y��{�ʹ�#אaդ������gK��an�:���\l��ƙ碢ĩB$���+C:&��x��v�ӥu�G�ݟ>Y����
;���3d�R�6�@�����ZU��w����n�}��w�$M�{�����Bo:��Y�������M��:�0!g,g�y�2��)/�D�cb�W�C�fY,�6����:Wm��5׽\c������ɷ�q�A�8��c ��gYވ�xs���r�Ų��8�ьݦ��w��JS��Ν"��i$�2wc�1���+2��*�]�J.[�~�ݪt�x���������;��h[	����J��?F��.b�&��u냨���H�y��V;�\�6␙�kn��8�0wJ�d��&݌��]�s�q@d!@�[G�.�KG/
�m��Ǭ:��1��ܑ�g�xd�zF��2�TιN ���H}�c�5�2��`J�;�[��'w<H��[�u�p���9ˏ.�Cq��=$����b�0F�l1µ~�ERW��oG��)�:�����������dK�e��ڼf�k�}�3��̶��z䚤�C ��������&��;�NVG�}�r�,�`,|dX�qz0Lw���9�:rs�;���6�P4�)
,[�j6�7۪4ޠ*$i�2�jΧ������`|	#�|�K�^H��LuD�,�yHء[�3{��W�D&�۠����ِ�K4ԋC	�F��kZ���qy|�'[]c{:��Eb諛k��M�c���ݼj4y,˨d��$�EO.�G��6����N���~�q����M�T퇮�l���B�+FΦ��Dͽ������W&]ϒ�\�/�LJ�C�ɪ}}Ne�SZ2G(w<�'ju�/�β��:m�S�˙���yZsr�b�ᕮl�9Y)v�%׳B-f��ֈ6Cы��Y*e�f�Ӫ�� ���n�ƒcLÇ��-�U���X%ǰX83���f����ڔ�*���ww֨�aMl�o^	�&oq�j#75W��黽u�V#�`��ݩ��bS���? ���'�*\f���wq�C$�O��8�x�&���q�w�!s���-��*n����Fum�
9���l�3�f̬M�2s� ��۳t@�����1^���wK�;ܲ���)c�]���hJ�2�\+��v�Ϸz�So'	:������:�x�ݚH���虶����e��{���`9�-G��N,<��Yz6�"U�x�bۗIfdP����j�ޙl��U�Xٽ�h
���5'�h�[}[*��we\���+Ĵ���(�Ӥ�x��K�n��wV��+���0��j���Z�W�ibDov��:��h8�wҹ�@ئ�snJ�J4�L�U��Q޺{�ƪ��s�媐4�s4ڈA��������a�2���޹[/�\��N�eܨI�9��� j�w]7O;�/6=�	�KN�1�z,dGGFv�V�sc�u�Ҙ����33n������8њ�cވ��0�u�󥽇n�7G�۸A� �nP��܈u��0�KR��{�b�)�{j3N�b��_h����umwD��l�&n�7��N��x��N�}+%��^`�k�䑲7�Kjе�SY�y�nY٬X@�MY���R��vu�&���g���W��[#��QH��W	����|�F�L��/�d�v�8��	�Xl�E�{��ɪ�t��i��5��Y$\���(Bh�7:���҂9Ӗ�Luچ�є�p�1b�F��!�9��ݘ�HHC����X��M^�#t��V�b���Gs�Zj���]6��QG-#˧n;�r��ҭ	�)�����a#z��t��cz��#]��ą�I�ѵ��F{2	�h}��FW@�[��Ȭ<)�C3�;y'J��A��Ӕ[������ok�!$wBv�j!����sK�S�;Ց�ҷ��n��Y�F��I���cJ��[`�jn8�:��xE�sc��lG���ZN�C�w����l�t�Nt���<�<5�K�*�8�9����P
D����֦wݣN,Β�b��X�U�/OSఆ��H��9��Fn͸���0���,u�ڹ!;Z��!:�Z:�Z�IU�IU҆�-��@Nu_@�|�%�v�38�n��eX���P�G;0�FPz�+�W`��S($k�dPu���c3�k����L�q,�hfD4�p\xM����/rVr���j	�b�N��8{Q�����5K����u�9[l��_;�]��djMXԳc�זٵ�fD�r�Z1�.t۠��Vu��q7��Q�1��g���=�%UTWɈ>?n>�?���U�/w��|�W��e�Ye�Z}G���/�#�O�)r)���H	�Ҏ(�m��M�� �[N����K!��LB�d�%�
!Kmsa�e @4���>��L��;�I`A���)�M���ts�N
��PJ2�2�c�3heV^n���-��"�%�:��Ў `e⮭�Q�S;����9Mf�o�[�kV�4�r��qnk�(>���wѫ�ﬦ��$��5�.;�G�8έ��yN`�z�d��@�qn]�i���:�Q�2�6KI>�{�2�\�N��q�x�WC�B�{4f���ۑ�Ȇ=%�XǩGy�}֪vJJN烔����u%���n�*ˋPO���/��F޹�$%9��el��n޵6��Q�n�,B�"Wv���Ũ9uf���)j�j�,7&���j�6:�I�i3�l)q*o{q�X���{���S�	T"��&�hh<��y�w7^FU���)K5�ʱ��ٲx�R�42�S���`�/����	�_ %�(�_.n�V5��y��,��g><JK�
`rW�G:ͱb��<��46���]ۥc�H�*䤗+:�ފ�ai �]L�Ƴw�;��]_t�͎T4nG��l�]�楝L�gI��ۡr���l���\ڂd�us�W�o~�Mm:75::̙U�;0�� ��-̏i�Ht�G�ˋ V;�diZ��.�8i�$�I��m��8�ng������<�k�{���]ґ\����c�Ч[��)!������|�ۻ�nD!�eN�Jۑ�s��8��]�'��w�Ǯ��������Ҙ�5N&X`�ALF��"
151��F!Q�
*�r�$�f@SNB҅$��،��H���*K����q$�~�(�d�I"5p�lM�4�$�#N7~?�\t�]�o%띺�.�3y����zn���]��iמ^]wn�ӹ�;�;{��]݆�lr���g;anWw��.n�rG�tu��wI���8pˮ�tAwE�v���^�]Ύgs����-r�1t���swN:�8��y��Gi˻����s�,����%���ӥ�(���ػ�"�uws:�$9]�uѹ����]��Ю��Www$�M(��]ˎW$�\	��r뻙�ú��ݮ����]�ήq�N�'��t��q�6�C��w#�w	Ӯq�e�+������:����a���ws�;���8w9wv�7K9t��:
�s��ru�`	���d�tn�b�q�����뮌�]�ݹ�)�s'cv����)�qԗwۦst��;����N��;��&6s�s���ɀ$�c4���7s�%
w]8�v����ο{��~W��LX7H�IY��������u��3��U}E�N�܃)�1K����
`��q���ok�E�����m��h�vK�ܲ��j��a��h'-~b(KP�dJ0�1�H6�[��U��6򺮆X����q*?�e����Vz���k��@�'�:]_>��_���o3P#��ײcdk�9@�3�fM�t�3ʻH�%��	�x谵��ʳ���Q�>�D
�r���k�I/�D��5���}6ۓ[��Fݹ��xp�Eȇ�dV盄��gA&��O*���ˑ���W{��yiܑI�9z�k�${i!�+�{�~�*t���:�b���w��w|���['��z[��W����z��(:����#�x�����晱��\������a3&��=�|��t>��]1j��t�^��њ^o->�K��G���HuT�����5[���^�t��f�mee������]p�aa����NmF�4�=���S^���O��cum�{�R_�=T����0�lGs-Mu��F��<�f����>e�%a�
�k��ݵJs���.�}�����A절�x�_u��RVȵ���ͬ�j٦L��u�rTGM<b��̋,C�z^o�0h�(k�Ǯ���j��N�
w:�Kcks�@��0�,A�^�5�c�l�{ۑ�齛�ⓑ%�9G�N56���K�^�CC�+��UV��FL�/���5@��\���OM�T����d̨�f�W��@��U��m��~��""�PڼbF�uN\$���G�rc�S���Y
"E��f�J$尺��Uxb�s�C���yy�.���?y����*q��3���'��X���
�I�ޕ��[��%�ҵ���7�]�Fо �7]<{o(�f�v'����,�ִ	2���i��8�~���inbr���A�l�-���c.�ZOgkl5wovɬ�]S�u�O�]җ��z��V}�����1~ %��o�x^z9����^��g�c��`�*輺��>����Z���y!�F;}ru�C3l>��}1���o�q��%�`q���/3�p� 5���8g;�N4q�H�����$�A�@ד=���>T:�۟6�ik���+��*�.��[v���g����IGS����=a�'ϡ�6�Wa\s2���4f���y8(A�n�Tm�� ����qX��x3+o�vw�(omm�B�y��襢~�k�{	4�;</i�S![��b��(c4���G��Blӧvj�q�"T9oJqu���V�=������==yF{c�>=gIc��'e���9視ȥO�}����������y����l������Է��W�M{����%$jߩeШ�ԡ���W��z�rl�j?y��q��[wCm��*���6�k=ʹ�a����#y���ے/z�!�CC?���ί-�bo3ؼ����������#X�����N�e�zm���>,Ϋ���g���x���$�=��x�I�FxՆ-S�;=�i�x�k��p�g�/3�zN�Ny&:N��H"����\�n��~��$�Z��]�PRg���|��0*�H��4D��g�ӆN����/1C��i���w�gy��/Tt�5n���//z���(xᱮ�ӽ����t��`�f4���L`�qC��-UM�?�-J�����)�
�y(�&�tEΘޡ�.����/u�I�P���Ծ\�f,��/��W���Ɠ߃�9��/����F��)?u�x�#��|7�"�&І�	�$a���4�P�F{��q�R�I�V<	��u�Z�ʘ��7 ��I���M�vI���)t������:|4H>ߤ�-�6�힇�|�ngǤ��d�2fN�궼~��U��+�;f����3\���H�8N���O3��w���<j��ψ�z_�M���ULފK�:�w�D)^��S�:=���zx���!�:V^xv�a���I0/Y#%p�:�}��/�ϫ�Et�������&��m!�۹�[�_�p��M���U�y�]U+�����v���*�8�=��=v?;gG�b���vH߫�]���
��W�Q�����p���׵�e��G��&}O3g������>na�Y�ik7C���)<�����c���(�>��a7f,���,Mn�ӕǺ�	�7=����<A�Ͷ��Su�-���K���ż����CW�_�;\���ƍ�==WwVZR/�5������T��~�u�T����p���t�E��]�d��e��A\I��<�w;�W�ܳe�D挩�w$BLV���*v���r\0�ͫgB4�)���[���Z� n��Z5�Hƕت��W:�����s.nv��S��9��y��X6Rv���p�W��^u�x�v�t�V�R���u����s�Ы:y���ћ�_��]0g�h��Y�������%xa��txP�#=4�?R��ѭJ�R1:�������ϽO�=���\���x�*e8������#���{�z�N����{�	���-�����7O�N�P���{�==^�q�jz;��Q�V�E��Ք)Q�aV��a���	�tE�w�,�d����r�_�8b��eP��2�%���Du�r�^컝�hʏ�r �[��Nι�9�=�n�)��}=�a�4��B+�ov���֯�-u 4������.�;�3��>�N0]���=O�ێ���y��mT�Fc�.�^aʝ({2�^�����������kɮbԞ� I�z�l�n��Ha��\E�^y�Vz����] ��z�h�X*hw�R�ɩ�cHgNh����Q$��im���"�^T�0m�	�X�l�zVb>�Ӗr<a{�,{��а6�\v�����-҇X����9��2ų��7��JS��*�O-r�%q�qIˤ���G�Es\�}�;�]<� u��rwx�HK�`����ɇ���A��Ŝ���^����/ݐ���s����6���~�7��/~��g��KG�,&��Σ٬���6�d�F�Oz?s����mO3*��jI�k��G�0�6��0#Y��a�p2�h��=__��9�8���U��T�ˌMn�~�h׶������ԱJ�0b�k��G�RyG7���۝޵����}�fUEW�����}d�]VT�W�<c�Rz��6W+1�Q���o����I2F�,D}�EG����ީ��Pi^�̾� �»A���������D���&�{��r}<�Bm�KN罊-jߠ�3�ݭ���=��k�& ٬���$f��n�x�3\k�:�1���A��6c��>�5��P�>3d�L@��r��[��Sc���C�J�ݴ�`�R�tlܞ�(w!:X����S���B&��2��d�$`�c���S�F=|��{P;"�	��>�%�Z;x�6�ǈnU�d�2�ǼZ�Sբu���<��.>���o7��]>:e^���sR��hu!2��gC�a# e���hݻ�x}��;�sSNdU�����$�*���D]����䍐��'9H���	�&���T������=�m#2�p�����{�慠�~��T�l+�f�rO3�8{��Ǎ6N�k�3��(;9�ola����MV�ݜ�Z�A� ރ�W��$�A�}�&��d� ���*��O{��a>^��^�B�M�)��v���<�ס��xI�޶T׈f����7o29�x��w�]_���xy��u��k��3h�A/ν��§&>6��#����t)u�O��z�k&�wO.W���d,���n.�t�9��]����_]T�%9�
^��PևZTľ7^�ʂ�%�S��Ʊ����1mFk>{V��j��^�����MD��/ݻ"r��;6y����=&�$vq~��Ϭ��b�Ɉ] �q��ګ�YV��4Nڊ��(��إNΐ��/�\�^��m�M�h�_��qk�}[��`�Cq�ʘ¡�g>V�*V�w�d>�u]}���-:5��L�Ӎd���A��Cōj�陆mu�v��f8OV����$W����÷�(<6o!�p�$�Z�3��B�R���o��mCI�ʮ��~�ek�2��**2�u
lm[�g������S��*��/{�8�Ԙ��VG{�)x��J�Gvh%�,�d��J�XG�m�xmz�Y>�4�5��{�#	p�b5�����J\w�|ڭ���"�[�U��juX%��ߢl�1�Y���8���3��n�v�x�t��cOm\�柨Q�5�wJP�� vi�{ؒ���%���=��r��&Ƀ�ɓ�W�Ng�l�2�5��E�������]Y��=K~�N��J��:��<�&�x��*��k㸍x����J�=#��1Y^��ՁJ���p�6��I7�v��`F1�&ܜ�u��I���Wh*�T�Wg�W�r��r����>�ys�f�ѣw:A����vs�&������v���S{�=�5��uB�c���^�=����ԃ����8���T�gù�khf���a�t���L�G#YƢRQ���~|���T����K(�X/8��Ҍ�s�6�����cTW�{{R���T��r�����9�V�\��Ř%fU�L�����K���ob(�\ݕ������l�-Jj3ܢ��]n�U/����5�z+�{��<`��k����^�^�{ӓ���ncS�b'�Oq�w�;�s �����`Ft��i;��2f�/GE���>��,Mie����{��i����{EmnLh��k'{s�}�܇zc���k_��;7��ռ�$Λ�?	V;���_^6������ �g��Cem
�bM�����\�W�-��cr��=������o�z��j=���@׫��N�4�vu�>N��9e�,��<zVy���U���8� ��u�26)�F��"���7���C*�����vE�5��#��� �
�6�9��p,p����8����H��.7/�C����5s>;�o�^��;'���Ϩ���C`u�����i��n0A�r �k&6F��&��ׯ���ĽA_QZ=���� �陇��@�`RقYҐ��W��/X�^4�Wӛۋ��]+����ϷҰ^U�����iGD��L�+�G;��Wޓݲ�B�+��#z�S��}����qM�t(����-�vy�S[��htD���t��Ѕ�;�4�4��Pr �[��i��{`�i�=�e%��rcnnǷ�v����1��r�̇���^�������Ԟ�}]Y^�N��x?=�^4���Hd�w��q����U9���F���p��v9�����-rM2x�ד Y���l�Ь4*���5'��*�0Nv����"���T�_��;�tv��a-��+C��o��7Q9�'��yzS����)ضx�3j�N&OL��>nfy����D��wL��㘼��3�\���~a�x�k���{�����;;�,d�l ��wA�T���~�6�go���Jg�=����X��?(�ԵΎ�>�{�jM��*�K
�,.��+����W`"����ġ�ܪ�U1���V�vѹ1�w%�V��5�B�gn�x��Ye�Yzx;x�	��֨�|��N_P�MC�� r��-	Lݙt������X��$�[l%}q���P�����G	O�o���vt�4���<k�sjv��ֹrm�+��!�OR�E�u��K�®Z ��g�eJ���!��*�YuaM\�wmHK�j��}��-�_2�ԩd���4�{V�;n�K{n�ٖ^��^�YP$�o)R���t:;��+���;�����՘9��++J�7�G�j�`�!3ێ��	*�#p�<ıݮ��� s7�����0��7ܲ��J���T�:)�zq�7r��5v�C�Ō�s8s?isf!�3Gfl�f��Q�X���s��wy��b�3Ftʅ�Q(K�P��ԑ�!����Ǜ�}�c-HX���M��Q�eJ�s\)@���?%��`R1n�g��W8�\��wB���}".�Cr��<�讆��Ë2�&R���B�-`>ҭ�f[��ס�R�3��E�9	�^��62�^Z[8|Paݏ�b�iF>��Z�33�'����$��R�ݐ"���s6␌U�3]��?n��N�ˬn��ՑK�cv+)��V��XT�k�k�]��*-����qh�3�� ��t���RS��������-H�e��q'�?N�z�����.���Va��ۆRMA/V7�5�Y��A�q�5���*��
��Pf���(vT�˻��(t�2�Ȧ��q���cF�����V0X��ڇ%�x�<�]H��hI�ENR��`�9�&���hE-�&��9Axo���v�+.���9�}����,!6J��Ei�6͵A�	�ɓAX�oT�b��h�t��v�P�k��9�&��d�r7�w�޻!�Z��T�յ;����U�b�&����S�<��t|L�m��_l�]���S��`Z�o�cY�c�mN�.��S�pùp��%�L���;y.�\LX��iX�b�|�\䭮
�^i��dÇ:XB�P��(Qy�LVC�z�,�u�oNwf��vۈ��wy��L�kf��\��lC�km��
X�,�B��}�+-To�Ʃ�=/���!]�����^8oH���s�+�w�E(=�꾉P�����X��9�n��, ��g|�(��$t�f�]J�GD�j3-��fvVOJu!�q�Y����Œ�m8E������;>��qg�0:�<F�Oj�J����n���ܹ��m���dWL�^��$T�u�|�(�kR�S��Y	�+�#mv��ښ��}{��w�	ƝJR�eL=t;OZ��R�����{�w�vap��;oQ���H�������G(���ݩ�,�f��� *۴��z�64vB�һ���k��Dg4��}q�@�xKh���l�tfß���U�R<!۫�cfvA���ms[m�XC+vb,�ߏ-{)f<�֣�X�Ј�Y"�i����-�Q�p`�����$�R�,`,�]�t� ��&�Wv�2��ݺ�K�wu�D�����P9���]!����wn�E(2�t�D�L�Đ�tc�t�v�a�3&M� e\��Ȓ139�
��37s�z���$���D��c���o;������N���yw��8޻���0F��We�4�{���멦$nq"W:�yw����2t��v�\u��݃.\&]]�����%wq���;��w7u�2#&��L��w!ۮ�<�<��<�q�"n�u���].�;�u�q����4#ˎứDMȒ�u��;��Wk��w�r�]wuΛ��;����u�h��u�]�����^���p	;u�뻌���H�C=�(�Q%�ܑ����Oz�JKίv����{�+۸�NnPF5s�Sv]&�,�㐥''p,zt�������.�t�.qv��r���{������?_~=������cnv�go�%��:�u-��p�D�]c�����e��8�Y�(���5�Z��=����pM��������q��|3k)z�A�g�C|���r�-�����goa�j�~~�Nj��Y��f�GB֦Ꮼ�=�'�O/Nk����͛�Y�}�%�W��R2a����p�>
i��Kr��ɬ��ƲwwT��KC:Aii�	��##)�Lz9��g�䩛�a�PY6��Z^F�2�{�%G&�������N�Ŵa�w��p����W���"Skz��p�;�8���*�^�����Ms�f�ir�Te'��-b^C,`p�e	�y���!�������M�u�5���B���D�.���XTi5؈�|j�;/ʅ+I�>c'�9�'�b��m��9q����C�O�/�7�WDJt����ƩƼQ���#ny���.WG��j0�j��P�̈́�J���&겸�����mzzx1�a�`�̧q>=J�|1���I����1׮p6�P⬌;1��6\����#G�!��!6Н�՝6�R{¥���t^��I�����ݸ�U�������,!	L�u0�o>`��}G?���.x�nᜫZˢ�@��Wn���Z�;U�M��kk���V�[����7���!6��3�&]�љ�6�
�
��WF��U6�!��a���9����M�Ȫ�j%�9)��i��[�i�[��0.�:R@������lk38>k6��g�e:֍gO�{٩���������7�_,Hwɤho�M,� �,����=B���0��7�wr[�e�۫��;��q����z:�hQ�u6NXTF01�@\��p[�4u|@��¡C`�v�oOll�(,��̦E�Yc߹t�W_��sP/��P�n�������.��q�ko:^�t��Yz��� b�YʄvI�,��~HN��<S�n�?t��;�Bۆ�C�cb�WM�vu��;@С4���W;#Y-��f�D�f��z��ŉs�h����R.�ߔ��	׭��6�H�x8�����I�z�m��?���4��������u˫�?{�0��H�˙����cgְ�ˋ��6
I����c{�d^�}]c6*��v��j\U[��������xf���Y$5��*͖}Xŕ�*I������9�G�ԡ?N%k�KDe]�ѫs��%xmEc"�'��N��1�Q�g/��|ȋoC��P-�5�Lmj��{fo����◄�봓:ū�0���:e\��)��-R%T�SP
�۹�O��-E?y~�?ۛ�5�7{���H�#��O�^�R�Y�����G��D={�s�f&N���r7ILY�Z�X��Bm).�&T����;���qI��[΢5�ӈe�0�9���:�LhKep�l.7���u1��S�b<�{����A�`O�KY�o���t���5I�v'���Xt?�Bl4��O�}%��tBd��b%9�R�j�UE8��3O�LN�y"U�d�lz��C6�޶�Jq���1�����e��Y�i�3'�RdY�b�ό��'1'w"��_�����Z���������!��'8���UeS���X�8SV\�j�y�X5��)����H-@=���rԸ�D,��C��[?9d���s�ä��S�C�ػ��a��9"8�7h��9+�[1\��qH�#���$K��ը�ó�Ǐ�=���¢��Q.v�2ծ�9��J������*�
���f�ְ��a��{p�0�h����wN3���)�6��:����@@PYT�m��B�(V���V���%���N!�����5�NwT�;:�kT}B�0q�<��,�9o`��e��E�6��]5�|��q�el.y��]�]�����l�@������������{k�dG�^���p��g�G�m���3��t�t��,ݏ^ǥ���c�)��yw�	��_=)��s���}�r6�.��j��Վ������%�bՓ!k�9\��]<�%3qE�$�s >���^b�øV^��o���+��D����XkKV8�����ê��6��3��c�¦�s�����/n)���2�NCz2��Z���������d4�m�?����ξt�����\V�&A!�p�hG��zd��w��c[��0��
�]u/X��F���.�Bj-=��^�^���yj �Y!
��ME���D>L��>�zz	�լ�����<>1~��e\N,3teT8h�!s�aT��Q�Up�7�� گ�_+�Z����N䨇%���9���&H��ˣ.j����t)�	�X�Rp[�t��K<������׫pw*�}��3_�Rf�YE�����'�eL��W�k��Ѕz�&�b�fs.�}��y�{t�a-JR��7�C_q�=[�zC��" �^��Bz��:{���tn�D��Ɲ�9���]̦���Ĳ.��)������~�.(=�z��[[$f���0\�9�pf&l�k���:H�$ٔ�"��9T��9�g�#�-��ߒP ����(���(t�)Ǧ,�����ͬ� �T��a�la��*��]/AdZ~b������p�^[��V枮۷)w^��0��M��[�vi:�3la7"��Sz��z�w9�R;���j�;E�3�Y�T������]�;<X&]�����fN��^���?���m��O*���Z�]"ѢsPQoTG��\�Ƅ�f�ɕ� �-秕oZ�ɤ�d�JP�\�e�f\��J��Z�Ik��i�:V����E�ũ]�����=��3�#&��/�>�yN�<Z_��"9�Ƿc��!��a��p�_�ӳM��=E���U�)���R[������ ����Քxo)��uF+�f�B�:ăÐP|������^��&�fb�1-�-����/:�w�6&��|J=���g�
=r�k�,3�.�������E�ϐ��ע�w(��m�U�Ү7d��-��wVa�c��ŠvW�I�Ũu��Ϻ%�r���ŝA"��O<���N�<�^;+�����xq��Fmcx)z�O�j4'Ț�z0 �ϫO�N#���F�'k���������ֈ�Zp(- C�"�'����H�ᛆ���$��|�dÇo�0�We\[�S��P]y���^Y�X���B��##)�75>�z���5 �*f�eM�����9��C�"�B����}�ʘc 0��|آ�=7��WH�x��a�y��O3��6��~e]6�S.�!�LS�6��w�ൻ:872X���UӬ(�T-U��X���d#�@H=���=w*�Y��5��t���F!�(�E� S+
���fz#�����Ξi����H��{��oUV�Jn KQ�)7���T�*'�.�_pچ�Z�>J��u��f�%�o@�F�fv�Ei��������G�G��9]2+����R��mJ�[���t74���sz��ƅ�97m�rM����)�NC��4�Tt�o��{3�0NNk������
�	_B/�?D�Iz5LU9�R)�i5��G0"��{��;Auuӗ��7���#!��at�uN���f N�<z�$�b)9Y�"�{p�CV���}�U��Ə`����Hf�<�@��r!6���n�gM���K�Bn���Z~O��=�q��OQG\���3{{ZA�zi�����8|``y񁯇!��\�{;��<E\h��,��hͩs��WH��~/��<�!��,k�?���B�Q���P��\�&],��:��C�
b������)�����ɷ���je�+b�ٶv}.���ǁ~��ŷ�E�GV5l<�.K&��v��>�F��P�wx�k,{����b��x��O�P�n�`��\b�)����gA�}M���M���Ϲ�Dwa��df�$��
�-^O�����n��K����;׵�a!�"e�Ds;B<:�9;#Y+ޠ��s�N��O�����35���{x].��X��r�p�����O`C��C@�q�>���\��m��oO�זi�[���|I��w� �s����˒��4�!��! �ol���s3�4�&���/7�<�e����K���Ce�Ӆ�Fd߽�8P�z�3�M�40���wyO�u�ukSBGOf����Zx����8�Xӽo)�ҦZ:2M�>����g�[.�#������%��N�$2q`yfqm�c��zm��Ę��o�i�m��ȧ|�R� =Ų/~���s�ԇ�΅���B�1ҁb�ۑ�8X�1nd���}͛eY���=;��`d���v��[̃8��\F`�ޮ������p��jЂ~ka�Cb�k=��|jʋ�6�����]�o�8�C"'m	��~F��Xٌ��_�!Z�ǢS�IQ�ZɪL)� ��ڼ���!,�G(�l�
S/��!��J�]4�N���f�}	���2.�����J���tk���ܠ�ne�/{{��j~�����}]0�p|�5�#��>�}	!�݆a�ǩRdޝ�â�O[)�ۤk^,y�D�n:l�y�-ᄍF4�C����_Fɽ5��ɹ�rm�79;+��^lr�d]g��敥�m���Iq\�AYc�j��=����\��������~��[�T�P�c&f<7W(��RX��;P�3��P�kAa�����#�=%2��z|yz s,zb���E��M��	U�-ts*�XI{���9�Á��~�3P�kpj��N�QJ8��%�j�j�zm�o �mj�N��O*�Vi7M��{��&�~qUf��6�tdK�cA�L�n�#ع�K�,��ɢ���N��8�a���v8����:�s���R�gE9XgV��v�s����/f^�g.�7���ɋ_�t&5=#�s��L�[�^Oҵ�%�	P��>�`��ߟjI�>f�G�
v+��R�>`�����Q~�Y��M��k:�jR�l2�p;-�q|1-s��u�&��53�}���/ʇ��_A�&�Z�)m.ɑyz��<1��gz��sJ�%��w{�#�u�F��Ob��F~Ш��ŕ�O��$|�jya�"��\܄6<��!=�{4��#�� ^E��CL�C�J�D6l��m�lg�`K{Ќ�O����f�˅�ޒ����]k�9A��@�S�4y^i��t���y�'9?[�rS͵�&o�������#hd\X���{��j�ʩlj\�.{�2��B��G�;{v��[Z�z�ߝh�}>ي�� �3����?���?��}�ڨx�?����L��v�Q��\�O[�λw��ul̂�;�j�Ui�6Q���ώ~3�@�		k�o��}/��R�-4�KU䧎��[SlO?ZR�&P���FM���ܯD��j5�h8Z�> �^��Bp#�=3U�U��)�W�8�^B-�Z�n��C4J�+��6��:a��w��'YGepR�����������#ASM��X-�yܖ,�Ǝ�$�ն�&#�ɦ�<�n9M��9�kW��+���=E���V�'V^�m�[p����b;�o;6dw~{� ��P�O��)��x���^�b���x�E�x�4Q�uNC�~T5ip|���������F^�7Oc.el2]M����ك=�Yj����tÔ��+�)�b�v�1���6�m��q��k45R��k F�5���4�uOH,k�n��N�⮗X����PX֩N��5)S�BDkM�J���w�]԰�(�-�0���;4]\���jSB���~�t��e�Y<��mB5�w6��Q���f:9��/nl�#�:=í~�٦�byz�cC�6��x�XU����X�Of��~�<�O�^|gﮡ;C���tØO���:�fFN���Ϗ�
P������U�<�gW2�2���ϧ�G6��f%�3�.-�>�08B���uP3X�n�����+��]Nç9��o��_�C�k����W��lZ�X�c#�]���;KqM��a�Vmi1���	�q1*o^��f�<d9#6�������)�!(���_Cz�z�NoGK5��J$�{G�kaKU���)�g�?�6}哝⿷��yfY���%�%ro/MͶ�<N�D�iz�ߗҹ-[�!��I��D�V�ǫ��Y�!���ܐm��]<�nk��ȫ�T�Y�Ҏ�������֗�Jvk;��\�j���Mm�s���b|�p���N��T8!���;k�:��N`%�L�����Q��S�����y��|������o,Y�<�e�C�� ���_*�-3��_�?|<�q��_8�G>z�grRͭ�w��#ǥ��c���Ů��J�m�5N�z6m=cո�t�w�-��{GUX�'��LZ�:�85n��U���X#[4�Y�W��<#}��P�V�ʅ�I�1�`q����M��jM��DK����8�W�!
�U���'�s���+U������Gk��� ��p;�'�\o4�_y�Tf2�ؔ!����ð_	M�����'�b%9��E2�Q���#ny�k�������,�OsgZ�4�҈|@Ǣ���gj�X�����3]	�vɒ_��9����@�^�T��I��<�D\����������W��'��D����nΊi/�
�i!7K��h��~���6�v1f���Z�}E�wyt���]�<#�h��ƃ_B�|����\��x�OV��������u�MF�y\���N
�y���ܫ��$Xׅ�6K�y�d�i�h�<�\���f_��B�P��L�
�k�zR~lF<�R�A��D��jֈ�U��-�!�.�t�馚i��i����<�k�M���m��3ɋ1v	g6��c0`�j?M�͹��cg���:غ��t���`�n'Xm9��u����^s85Ϻַ�u�Y*�
��Aj[��L�Ƿ�FPq6�z�s�����J�C=f�ÀC�`�Y"%�\s�N�^�p�R�^0�J'�J�N֣��Y�wa_K���7p]g۳��G��Rw;;Q�iޡ��Gh���@C�foM�WM�df��(F�J��[��iu���o)Վ��t�Y�SqK�|B�m���S-���iT�+�v����8���uk�ѲZY��P��+!���]���n)Z���0Z�Ȥ�.G�Y�m�n��=۳D����F����ӊ9;�˅ԭq����ivm�W}�iexԲ
{�΍˓����H*�<ֹ�������	h���	Ȱ^1i-&fe�d�72Bvqڹ�;mN�U�kI5|�ꀰ�pC�7W���5V�����h����9�����6��¬t�:������X��9�\0-���[Pe-;1G+6�0��i�ѮT�Ȩ"奣�br ��:u�s!T�õ�wEۚ�5�&���#p�KykkoE��d��3��u���Uf���*i�25U�M������n1�s2������D�g*Pȇ4����;���31�JC��o'�Yֆm豴a(�</�X�J�f S+5c�����(o�󶱒�(t[+�Mz��vL�������s.�G�R�Ѐ���6(����~�z�z�y���(t�.ã����ѧe5y�Sf�v��n����j�܌G'RM&Iu��X��� fdY�8w5tt.[�Q�L�2;'8U���q�u&t�cĠ����&�u�X�fm4�a�c�,^�Z���k�z��[��"D,7�,��Wb�{��Jĥ�wf8ݜ��dDյ�����vtr�}n��h�(�wб�+z)���/7i��{s�̂
=�b��(�/E]��a�J?	��ﲋ���ngD�!;x�i�̥��E��X����u��"�]4oaUbZ�)kN���{�'����G�N���JgϞ�c��g\�[�]�lb��ٸ�^ܵ1�����XW �es���;��J��"CD��J��v�F;CZ�ގ��Y�uob��*��)�g�X�We��Xvr���L�<���9��v������۽;��%���=j���ݧ�;�����B:'��kaJ��Hl�w1�R�]��+Uo@�v�>G5�h�.����ע����k@�[��V"��cVi�^T��j�n�V�r������x�ǯP���c��7WR`q�ӻ���\ܹ/�}�{| 2R��3E�Q)v�r�mM��5�����`!F^�tdo$�C�e��[�Dc�*��2�wL��7#=���6ol�`���\�/]X�RIt��ڻHD����L���]ӷ^����Q�r�ݣKӤ�v���w���˴��s����n��d��u޺�<�ǜY�J������������,s�&yrh�"7�7s���&$��t�g�n�5�W#Dd���W+�wQ%E=ې&�I�I����ݒ4�Õۺ��F�!$���#F�F2I����b1e!-y� k���������3 ��)%��삋�6�
�О�TƤ�uHQ�`��X�(�w] `!@��$�Ѳ.r�]h��wF0 �уL�RY�(ە̉�
a�����AL��E;�I�Jdwt�(T�1����Fd���hb&�$"��Y4Y1R3��k��a�3��������{�'{���^���	����R��W}6&6֠��mhmt�Ǌol���aW������	�B�p��gNԢ�ܺ�q9�}.G�1��0ZX�`�I��%F	 B׋E��^<K�r&-����r�h��2:����=zT?>�r�i�&Y�z�NǧT��j���}�!۠�C(�.]ݗ�{10d89g�p�����_=����q�fQqɑ�`�! ���e�\�\�Aj�c]Z��9�=�ø�s�:�퀹m0��ld���Ý"I��e�f����\�Fr�4�j�N��WF4&�w�R����"LcE�3����\��m�����e�w�{�l� �vk�#�ku�jf�{�K����C"b�ړ�����N�Ϥ2�,=Ų/�t����Eb�lU���+v+Z��A��A�pd��Fu��W���dgO<��8����ڨ�p��!�H����g<��&��W�j������[�nE�r�Om�Qp����b��<�k�U��A�
ϴD�BbS���b����e�~�'W�P�~
�0����g*"k�+���+ﳫ�o�}��U�*��R�u�'j��n})����'.��kk��
aGT���8����xuV�a�;�����5�\�X/����1��Fy�>%W4ff~[��oZK����lqn�@A�*1F~4�\u�a��Dn�:����ɑ��x�.�W*���F���O�E�5�H��h��5�yWek�/J7�{ �oN\FV�j��q�[,��H����e���aN�?�}_}U_{;�{s�s���׀X��E'���/�E�;� �F8� �cL9	����G`}ۦM�b����C�����E���m�[�ޅ�4���A�>�\�%�r�e�����y?x�,��nO�oD��P�]���B�L'��熵P�����#�%<;�F�>;{"�vCO���]m�
���Ԅ@M��y��M�a�3X��E���3`+�a ��}nΫ�Zϊ^UI��w��
����C���N���q�i�+qܟ�k�PK�6�R#��r�f���)�C��YN����;�0p3@Cc�a�͉�l;-�gQa�C
T\rx4�붫Ӽ�d��W����h%R��@���g3�"]�p04Ba�6ߣ!�'U3Y^;�������9ӱC/+�$�x.��6�30�C���μ��\E{DauR-�$)W;�t�0Q��I��K��yC��HzJ��l8"Ϩr�?P�	�Y��W+ᮅ�~8�v�B�";�>dr}��Ƕ��<���yn � ^��PDךE�S�� ޏW!�Z�����3V�S���G-�y�ӓEÞ�P�q,�7��n����ٌ�Kx�4��07z��_jR��G����f�t_bO�fZu�i9c����A�&�tX�[�r�<��w� y��%�ss�/�^ x����r�+ӻ鉗?(�|XP���H���ľ4���[j�!s�B�Ut(����dK�N�ԣ�����u8~�Dz���P����p��?���l�%�0��:��<n�j�
Ӽ��[e��g���Sn�K�}���S��ϋ;Y��0(������Bh����(؞M���Y�>1@2�O�8�`�z{�.�K�j�Oʅ�J=����ˌ7�����FUdp���#m�`�f�W��$�Ĳ.��L��V�F�
�0Q�����_�v|%�~����g�93B��^9�1�"D�2�ͼ�L�R��g�V�]���r�Z0��o�m����ux�2x��?��x��t(�N�)�~Y���T6�0<�1��X�)��<y�����ȸ��>���&�~���٢�Sۄ����V4�oE�ԫ�1kuF��䃮�@�z/n;`8A���0eё-��d�2 ���u�O�sN�v�R����Y��@���~cS�â�?t^�����!�]0���xhŢ*�u.��A�������^SU�\�O\4y�d�(�!�ر�~=7W|��۪�ʋy���c��υֵ�m\�/����Ճn�awlT�sIs��9�����;h��LhQ��iݎ<��͛��kK���V�+��W�U~��� <v����V�jf���6�ʔĲ���F}8�b9���1����@0��3'�Lk��j���r���Cκ/r���lx;n��%��Ǥ��-�����`��Vs��U+Wc?���_J1�Զ��O�:a���DJ�/~���Kdf�0R���׊hJ&���n_2`�B5*6���T!��"���D��BC�?�Y��	��_��i�7&m�#Er:�[mW7��Zs��
��8y���z�-35B��r�xy�Ǐ)|���g��1�֪Jh��-��ۻ7��r��+"��Q�Y�i�q+A�N�[O�X����K�Җ��wTuc��Gr��w�0~C�+�e	�'⢃&>X���UӬ(�ǡoV�^�o��P1I~y�w�K+�.mss��:���2p��; ��J��=��	��~[�ܥȅJ�]�m�5�l��I�dU;۹4�)���N� �D�e	x,|$>��_=q�I�|�s���i5�f�J牅:Z�=[��d�������`�fڝ���0Ta;�R�����?�ի"�7?<�`v���6�~�ǸE�ɚ��V3��s�r㦷�����,�3�l_�ha�#7�9�j���&������IqluX�^��3����xu�����y��M��6�F�|vk6�|��KO�J[�o�c/F��ʻ$�8���[�I6�tjپ��"=�X�P;E�~�d���5�ۓA���9\Ú�=^��y�XE�A�yȄ����K�(vmZΰ�Jz�Ή�Y��K�1z�q<�^���:��>=!�|�1��0Q�>�#�k;.~�s2�Zn:}�m���t�WdyBԍcA #��bC���$X���Ѕܖ]y}E�0hu�)�z���bʣ:@��I�	e�M[]����،y R�G�L�e{b�ٶF���6���
Eݽ^�����m���t!�9O����9P�n��qg�V��]>��&+����y_E$���0��FVUh����@0�N����DW���!���uC'�&Dwa��df�+! ��9]]��ub99Va�;�G6+d�,Z���s�<{Ds;G�(-10�͏Nφ�V7�?<�u	�M���n������|���Ք�[��`É:"���x5�%�q�ߙ��u�zq��ܫ�8'ۉ����;�h�p��]�S4��$�PJm�jG�̵���������x>bA�����Ǌ&�d��膊��#r$��-��5��y�^[	-����Fu��f�V@���{��_vqT��b%�疾ະ�=�̹a�5�h"N�d��5�h�O�^�Ck:�Yݱ����ؼ8f�5�,L_�}kgn-��Ra�:GS�jcX#��h��MRV�{�rT��WV�Q'�����v��`ԃJ[��D���jl�S�\�~*��T5ѭUu�^�δWEw�z�`��^�u�����EcPނ�_��	�d	bQ�g�c�����ی6�q���3_rWM���� O�Ø�a�!��g�i�ƽϣ�e�h�'X��R��v�\�ҹ�����XG.q��.�������(2�^�r��~�Ǎ~��}�?�������d�_Oj<�{�+��)ž�0�ȶ�WL?��5� z��/�?V��\^j��mf2�~��0�Rg�O	��y��W�(���0�4dAƑB~����l����g�C�~�ܬ�v�r�'�Fm�u��e��n���f�~Y� ��{e�D{�%,\ͫ^��x~y�Ƣ����(�L*�J疯Z�E��M%�#�%<;�F��G�9�C�ei��O΃��2:m�"n/S�\��&�Y�2q��%Qak���]k5��/�a��~�L��w�e��ݾ�.>�h<�?�}c!��sO�(Lk�zG6��4-Xu+u��Z�t���rV�E��Tk�)���X�j�{�a���~Cc�D��6��Ia��o#y��Z݅H��i-����W~�v������s0��r�T��H�\��"Эq����&hM�[q�bf�vb�����g�?`Gpţ'�\������],��Kj�;1�R�̐!!}���g��'T��:�ԆL=��DAcWS��M��e�������h@"땽�q��n�U[�����3NW���z���g&;�����~�{��0x4����������b�,�¸ėj&Y��8��Ls�[ ���^]�����L��s������"��ހ�]Cκ`�woS�����5��	A(4�L�I�ʇD��G(��}|�y��ey��C2�p&pBN$Fd��&���6>k�[��@�x���y^eI��En��6w;]�/���#�&}��[_:)�~!�������&���UKcP\�.{�A�8�%�*z�=�mA�m��҅�k�­�d-���^�tS�~8`#���vq�����!֊��^9�1�����ߺ����zAc^X�R{
�л���zǫve+(���<��,�яxd5���H��[�����l�5(BS+c��R�&��*��g�}Ǆ�o��!����K����{��;�67�pzB^�h@"E�O�̤�<^%�u�s�1(�a�-u�R���;�nJ�3��{�d{٬���X��l3��L	x�A��"D�2���ri:g�g)�]`�eX���<�VK�=㵕<���f~�=��FxK��m^)׍��4��9�Z�]�역(03͵-��t��W�[ۍa�ݾ�`wuӴ���5N����>���oWV�sC\z�X��c���_Q�cC��k��s&š��UV��ٚg5k��U�fu�����TS�
(� ��մ�ŋ��-�mo��b��Mt3c9��OHLha�o'qT*�u�I��q>�;�u�Fo6ѝ���w,lCzj_��������B��?>OFė[�3lW���nj��.�<���Ȝ��`�Q�j@~�����
SXA��|GЎ�A{W=p�]}5���"�m@��lݮبά`WB�I��R�>?\d�s�@:
��'�}�mʗ,�M�<Q�c�MO�P�ݎ���c~��1�Q���z-��k�f4
���>� ��zᡯ������n�oN�A�",��'�|����l��E���a�zHz���\b� L[1f�D[OS�c��f޸N�/�p~aA�xQe�^��#�2=�X�K��)�[Z��Y���M�;�T�d9=��J ط�"��{"Y�9hjd�C�$���w��ꗿ&������ ����{�m��qn�ah_e�����O\�o~�
b������q}������>c��<�WGO"�nj�n�2+&��}��Y���b�O��RO]���?��<��p�1d@�ksC�y���I������b���Oy�:Gl'KNZ��ɉ��^���ҲMN���!�b��Ap��;VXR���)D��rZ����z���a#�{�����b�ʅ��wT�l��,��w7{�1��O���J�$��w��W��]U[%Z�j̫kk[~?���F┕��ᡗ����ol��7���c��ɩb�O`J��Fcս[�{lw���y�`F̎|���g	�g�����`!�d���'�K"�R�e~U�V�0����I��s�#"ou��v�����i1h_��&��'�=?U���:}�^~�N��1��,��X� =kL��y���{{���?U,���Q|�?*��҆m����3�e;�=J�~����|x�gUjodƍ;���W��WP�\Ú�E���}��l  �z�	����~Szσ��6���z����MD��/�\&2�Z~Y���K�-�t�����k��㧆��u��Ey\��ٖ$k�m>19q,PҫZ��/4�ct:I�/Hv��H���v��[#>��+���0�@C�:�hW:�2)�A5mv4����"�yU��f��ͷ �g���K���ͮ���pn`�{/0�΋���~Ӓ)w�Ja����O��I��(�&8*�����Lp_�.�G`��W�����`kN|�i�-��hGW��N���`����7�2�o��t��Ј>9R<�8����p�u��K���� [���\��>����Hl���׽�;�]�qj�^�ߧ��ƥ��6�Ǫ�ܥ:r��H]a����Ή����*����&��程����Ƀ��gl��9�gG�����Z�[m���lm�E��<=����F�fqf���B_��E�r�kƾV�+�<�)�b��5��oP~y7�i��a�;����Z��5�Ԕ��`É:"�ׇ<����h8��o�q0��$Xg���'��#8���z�Uϟ��זe�p�yڂSl�PD�5�5'�y���%����m�1so�tܘ��,}�b���ϩ_�b�����Ÿ���3��3f�W����mO�8��6r�F-�8���n-��>c�`Mev^m���B~ka��%��k;���2�s&��=!����kNEMg�[�|�Շ>C(G9=�Y5�\��2״b��z�'�yݰ��ޟ�v���ɄC��k��_U�)��?��?�7F?y���ǊFAw����&�h�Q)ɒ�ݚ�n���O?_�T-Z�)�ߣf�H�h]��F4�t����A
Δwo���v���������L4�����o@LU�y��&�������F8���$f;�ޓ�ULѕk��NA�X-���Bz΁,hYT�ra'�Ͳ.���+K��;5�^w�~}�3wN^��x˶�i��zx���Dg9����jC:�޵�I��mT쵂���q�:��T�k;e�q��i�9�R�R�b�E�;I1R�^_j����T�l�*v�n���VQ���k�]3��-nI[ַ-7ıH����GF\K(��+\;MN+�:AP�����DL�ʖ�R7��ͮ,b��ζ-T+U�e֍Ґ���B�b�GmD��p���58@�^��v�%�B�A�	�o��g��(>c�̲�k7O��a��h.O4g��ݽ�e� ��v,_of�V3Z�
ħtҝ@���R�U����w�4�S�������i��7��+�(2�ô��f�I�u6�V�o,�*Д�IL]�c\+���Y�K7�F+��@NU7.ީ�)�lԂ�VQU�N�[�j\e�Ǜo�tp��.h6�����oPն5'��q��F�d�g��0^k�YԞY	lCE���+˃�l+���R7fȃ9�~���& ��Yxpkb�ӥe&`+bx�����L=�r��m�W-O��t4�Z�v��i�Y-^ipȃ6HG������))ZPk��j�C���-st^+�F��5�e�1)GXZw
�Mޗ�J����ss�-Pw;���3�#+�d��X�N����ֆd���j{�Jf�QuI����779������C��zt����A##������t�W����ӹ�T*�D�c9{p�S��w�͔D�oI��U=kT�cN�{3�N)>�P�]�^��Ż�ԂÕkb�u���\��N%�=��r=���.�@wf�z��vY 8�BH��	
�SJ�&i1�ҭ����Z��y(��[b��u����iX�]���3*4��*���>gf�Kr<��p���Q�pͫ���k�3��N�2�J�mm��b�[t��ss��i�Qf��z�)V4O�T����;���ށz��L`_+����d�82O5y��0P�ll~��9#����u�K&��)ܮ綁(R����h� ��[
W fo8���C��f�<e܀��`<R᭓&�l��K��n,{̖�̽��J�H�}���7%H�s`.�p>�GuMd�O��n.Y�Zg+h��E�Ůű<�EI��%���ںp�.؜TFg�cK�6A�ޫ���#!�ΉR�Fe-�V��+��e��t�!��l��\��3@�3���X�8i#�L��m���Y��'����}�3��[Z"�4�����82p�A��8XoZWӣBTxS,t}R���u� ���
.Wb�y�%�i�.]�E`{B�:�V�����]��6"1�����w6���i��/Y=j�ѧ
�6�Hj�b�}�;p�c0**l�au:\��.��U-�K
��3��s��z��û_H݉�B#8�q��u�m��E�﩮aB)�糺�����M�,i(.��:I�j4����!�bM��n���di6��U!$G�$�!cݻa���2Ɛ�P�".v!H1��2IC&q�$��H1�66';��4h�Yv��ܨb$2�#��PS9p؎n2������&W5��r��"�D�n��@0h�+�,I����]�m�H�ˢl�7Hӻ�����9���BWv�f�ٙ��f#���;��"�H�n\��r�Ous�2dŮpcr�"���$���wA�wv�t��Ʉ�v�yrw]@I�^q��J��˄���Lwu��u�e#1� Q!*(�˦�ƈ���~���-p�~�]<+�j�Z֚R�6N	�Xu���Ct�]3J�-Q��a�,l�^v��0��{둭[3�f��c�va!"bi*��V�h��6�mk���(5�����k~v��<�:�����(߰�aTJ疯Z�E�(,O��ˣ=�N�	�{�~f~�.��v�kb�-�"n/S�\���6�N8� �E���c&p�n.�Qg���Hm���ƨ/��A{P �8-=O���:6�r�`:��:ͻ��7Bɱ�lԭ�[�����ʂ\.�Ũ;��|�p�^��Y��	�miGR�\�0��1�77�0�Y���]5�af��5-�@�,���dȗx��1[��<��RgUsꝗd]^��t��,(q�.�L�v?�l:"��t�g/<��#N�[1��o�Ǯ�D�}(W�)�z:�VoS��Ȳh�Hz�PiD�4���d��;���UH�����S/J�3?�(E���ߦ���f���H<���r�ר�j��=r�ժ����v�u�2��u��<�0VR�)J?��:�˞3�OMnH6p{��L:�f�G�8yT�۳��?��q���>���n����`x?8��#�{fx�=�׽��칵.����ss�����n�[��vzRw��F����b��%]�	��i>$�r�[�M����S]v��&��}P�R��oMBu/�*���+�\7�r�T���Ď޼w����f�=�5�7�5x-�<CR��;�vݲX��y*��/v!E @` b"�������u�߮F#�j�Ͷ��PX�R{Tv�����z���
{gd�&C��'U"At�2��,�)iC�����O5�%2��%9�T�	�~�ߍwb�@�0����@L�=5�?ũ�e{��D��5�CG� �x@/�zF���g�Ĳ.��)�FS}�����wzFmWf~�Tu����B�v���ư�H�fS�x�Rt��T���H0��g�������.�KК�@� ٞ����z��<~���Я�a��*�qWK���b[w�:ƣcj�X|3��վ�K�!O�al!��B��"8F�P��.�I�`Zya�&^Q�i�Q;j۸n���B��=z�w9��C��k����C�h.��\G�h����]���ݻ��C�궑xru�6�'+Z�\X����(%����W�T�uvB��xr	]��i���?UOI3����t!�=����1׫�m��%]��Q��hϧ��j��cF,3���sTn��T'!�GZ��Ә�2��ݣ��a���^hn�a�/��1�!����7����	�w��ݧ���b�ݖ���7�%���9��ܛ�uc�2�,(b�v��R�^�����oZ���=De
n����|�*�D/8�)���t��2C�e��ϯ¢�Y7V�,��F���Xи*�݆�6��� �|��pt7|3_-����_kU�IlZ���Jֈ�bB!�A"g;9���juj�u`��K�l��PH���$ǂ��4>"T�{��f�Y�q��sk)z��_)J�[�nJw�vog���Â��lEC�dK< �����l��E��﷨s�{��EuMy�'�w���+6y�W��#>�y6����F�����҂��Nf�a������%��W�u�3�A�����Y6��G$>�ͧ�c�V�S��j��Hźm�ɝ֍������FǧB��v�W�y	M��PdԱM'�ь7ǣ1�[ռa=��/{w*�5r�|��թ����"XnT�H<��dC%W5{�N+�Ĳ/`�4�J��fq��%�"�M��m��1�ܬ�(,���C�6��A��'�'DN_	M������>�N^3�..�]�c�f�8�nr�{V�5��۞j|��T:<��a��a)f����f
�'p�p'�[k��x����:E��sȥCsj=^�#ϲE����	����n���Lre%WrE�d>���R�]�.�㐛��Z~X�y�z���:�M0�=!�Z1���G5�_��O2�d�p�M�19B���#�xA3�UHӾeK�R�j�$k���l�b�>�/Y��t�L)��|���vm�Z7oS��0�Nԡ}��-0��i���aWl�NK"�ʊ'gjm-̥vk�(�aq6uͽ���Zܳ�-�S�����m�ڣj�I�ѣ[�jѣmi5m2�EF]��V�)��q�\K.{ni���Z�`��j��I�] ��H%ݣc�4�r�T���5��R��u��P�+�\��ɚj=~��b2m�Tg�T�fJ�kH��k�U�����;�j�C���Pr^D;k��'���8ȥ�ԦY����]>����hmi�mv��.�3�j4��~�P��e��
���+=r��t�����T>�9����i�d��6��k�(�ԟ��j�$�ɔ�>(�����ؾzƟz�o޶Yc���Ý.�^�	����v-��0�A�^��6�h�.�!��.9�J�p��pᓏ��BΘ�*��j�zS�����{�Q�m��yڼSl�P���[�Z~h��{dS�V�,���V��ˍ�E��aqm��j�ݚ�m����!,U���z͛dD�b+e�蝝�U��[�;9tӼ A���9;�c��YA+ڊ��r�vA=yd	c�v�m�J�{��M�ݪ��F[��N���?~�.��>C(~�r0{��j�L.z�D �]�ޚb�'�3�X�*I%<�X���S�nރl=��L�n3y���y���Iw����\{0+&���������1��D�����T�Y{�df�{'k���6��9�k�B�����F/W�?��P&���1��5�؝�d�vTf�mLN7��{B�XՈ�m&���Ei*SUL���6����z�S�����{����U&�\�P�v׭aX����M����^�xf�jˊ�s��y���]H����ڞ���i:�j��
������iQ}XފE��t���Y�yn�*���0_.��ָ1C�Y�i�R�>�J�,�&*��"��\h�t�zw�xa�^������F��ޡ�C/C�O�=#�|.!��*��L$��Fm�tY�7x-/#N���v�w�:T֡j�L���8~h8I���7s�TQsrr��I�P9(yj�r�ͥ%�WEN���.�κ2p�6e��P��%��� �����=��~���+(Z�:��-%�]�T�U;^���߷W���ۯ>Wai�H+�+����`��� �c@OH��:^����뮮˻�:�(N�f�٘Û�ۋ^lS��oA/m	�q�F����p�`�#���69������)TV^�[��<����a�g��re�X�4^�5-�^=��/a���\"�̈́t&��s6F� ���KzY�9��v���¸ėj&Y����H:"����_���uG}g��ۊЗ���8�Hq�i�֩�2*�+��O7e�m�'���{�Y�f1��#I�j�ne���ր�VM��ԙ�M)�۩����z�'Z̫=mn���"�_b�;�g�Z������ ����̔���J�90�=9i�v�?��fZ��ѣZ�Z-C �
�B�;���Y姝j���',_��	;�����˰�z!���C�IzC���k�ǋ7�h����w��������z�O����I���'�)=�5�my�y�f�A�� ]ԇn�1tܥk2�9҆�,�y�\e9n������|E��!��W�+����P�W/ڴ����ѳOt���ۺ����LƖe
6Up��6�nb���g�!6Z��t �j�MnR���C�����G�
���KsQ�%6�2!b�IԜ�[���3K�.������~���v}6�*ַ9��	���Y�W�k��2���c��*S��^q�x����w�i���J�w����N�GI}��Ixpq��:��B^	4_��I�x�K"�9��F����K���$on��3��1�{��鵲GC6LA`�㜆:0���w��N�_*�R.��]ڶ$n�:���I�a���-�r]��&�Q���'�~=Bt?W���W�e;�����������'���������I�5Jw栜K���}��=�M�>�5�6$��?���m=l�r�B�U-'�Q�� 9��WSVk��H�FJ��9kfĚõ[[���ũsX{�Cf����<�i�,�u�V���8�=�R咶,�+�N����q�S�����9�%:v�����j�<Eɥ�F{DrA�\�_��F�mfq��U��w�"H���Tuة��yn֞ݵ���b;&aM�����J��Q��n�砲@|8Pϣ���%׾��Q���@[-��Tj��
m�NM2�G��52�J��=�ͰeA/t�J9��f����nb����5aUEI�����!�?6C�n>^�c�T��(�|�#>�z��5x��1��ٌ5Ok��ʦ��{Z�3��Tx3?��B/>��|/`Nç�6C�����lc�C�$@��f|s�G��m�4Z�����S4�g�%�r����@�Se�ӱ��q���m���S��²��/�Ѣ8n�ՔM�H�@��35h��n���O��a�������=cщ��ء�ws�3!=��]j��f�Ia��PE�%�<��m=�ZgK*���?�G2��X+�͜��R�y�&=��g���f��A�,�`X��sf���o
�E;�����c�9��6#PCp|ǘ���38�ڊ��%6��MK��FR��L/nϧR��!!Tn��ޭ�P�]�� ���0D�9S! ���"�UsWD �PF%�r�K'��&isk���K���f�4s,��&��+�z�]�_E�0��RZ��a�On	Խ�)��<M5EWL�\����%`kD��E��ߘ�j_	Ht ᛗ'ۤI�A��*.�wh���G
�ĭl��qH�T�uH��+����\q�ٖ��F:	WL#b��������b��5�k~?��jqow.n��o��Z����x2<2B�.͔%�0T/��$�7���������h��b�y,K�Z��nG�@���ԗx�ll�%���G�f��,�������BG��7^�uTKk=��/ٸ��Ut���Q���<�T1W0�z,� �}��l#�#��Bmu0��7W��q���96�^�
�c����1i�g���$�:���E.�azC�|`x�O[1R��p�gU�u:�C�N&Kr{z曬gֳ��Ȥ�7K��v�'�*o�@������2�>:b���Z��\������wf/�'�W:�&E1� ���Г�FM��
��'������]Ֆ��������������x7��� �^}�����~}�g�Ba�^5�=�H)�Bz6AsK��{�OE&��a��$z�2��O��<~4���u3��*�sC�>+ө�D.}���#��wQ�3bX ���\b���-���/��Ds;`(-b*9%��+5=Z�]l���ݔ-� z���Y�&�3Eڀ�.Ť�0������6�k�"]�`�oi��C�5����P�\�>ɗ3'Z7]��s�y�����v��[�VDwRH'�s�Z���/-'�iWoq�ݒ�b ]�>��Mf�N�
�ԳzÇ�D�6�F���{؏W#���t6�u+�y�m����Z�G���,��v&ع��-����'`�Q� ���`���Z��[�'�ʛ���[m9���z��3Mx��vJ)�dz!���>�S����nX�=���9��x����u��o'��c�_+�*��������x8�rb�VI^(γ�-x��M	�6�����ݭ]�
ۊg�@�;�N2�IݳX\M�'%���!?6A>��/��#�#���M��֔Z�~�:�+9N��~�	��V�i�6=�O�d~��ʾ���r��F�c�.�Q��Ǣ���%B��L%��[w�����g�[���&���x�r��k����|�<o�/!�-��'�)���Bҙ)�w�ȕ�d�=c�����~~�w_yL�3i�25hu|/FB�},�5�lM*L���&*�<�.W�M��|���Çdl���c�߄���AyZD:�xOH@��E�N�T��~Fm�u��01 �.O#�$�ݢ���V�h���y���\P(����Tx�_�S�#rr��L(�.yn�Qy~L�������zt�U�V.�s�{�sݻL���H���><���l�t��������Q��N8�����|�����_F6L샑l+65���w�zkf�A��-�Q��G�"%���n;wF����]~"�{x*!�����|qu;�=�}�ƭ%��M݃W��l�b�`��+�F �}��*.�qU�̊}f�!��v��Y���}vn���D�O'S�6@��#`.��j�s��h"�B! :���o���'�{�Ew�OO�ZQ"|��� ��
��Zz��|�~��q��<��_ѓ�1~�#����'�±�]+^�oA/m~��l���{�#�0p8_���k�#���2��ѧ�5y����j�L���b�Ú�~e�X��a�r�ƥ���k/�3��.�k�̣�J�8�4OA�"-��V�s��S�ޗ`;I�+��W�`v]��;���y�f�Ү����՝z�3��C���&P�/>�Tm�287��^=���C��Pb�K�lC�Wtuv�I�@؋m׊xe���2�Yq>��I��Qx��3cZ}yH�i��v�2�ڌ+	bZ��uh�^��(k�7N��������������5��1�`9V�1�g F;�:Qb�fl��ka���eТT�p��Dp�鯨k���~8p5��N"�gW���K4�]U�m��8�!y8�׵R���%6�2*X�Rr�m�g5��=��4)�Zm�vS�N%B2.%5��H�� �|���Є�V�%9�)�e	`�^q��Kݻ���;v�.�i��z}���$T8���U�kB���Ѡ���)2q�ͭ��a�sq�0ҙ��E�|�:3\=��ҫ ���W�XI�L�{J��G�2do�i"��=�K�9��ۻ[���T�d�uhFȰ�ۢ�N2�e�2�ù�hf�/Z�N����+t�͆ri���M��.��̗�l��"�a��.�W�7z�20Qx%����b�Yq.�o%�ED��w2��Rm�V�ݩ�x�LwbtW[�9�-ѽ`՚Ү �(\n��թԭP��*EϕѭEُve"�v���9;�r��+F8^	|�i	�{��:u%�I j��#w6��sO`7O]N	TPo�a�3s�7hfƚ��YD���s����ٻ�r\��V�����`�&��T#c(N�R!j�ef÷�>;Vz�[W k�Ǩ..�U�]H�di<nIK�.9�c���˽�kS����;IL�v[~gB�V�g����S2Ш�.��u���X������jY��nJq��9*�k���Ҳ������ҡu���nZ|�&��;��g�0��S��dP��/����u�'�Wi7Cs��ɾ��2=$���-����+����q��݋ة��0"�q"�=N��ѝd����������{%4�����Դ/�\�#L�Ȟ--J=��*�(�hwb��3��,uׁFF�����X-Y:͙�DF�,bXƬ��̒g��Ԧw29n]J�5�����^�5�9d�=ǽ!�;%��O���e�"�K��\ټ/rKZpN�V���\��}.�1�e�6�r�;��>�o�')?������ή��4�۽2!�[�y���9\�5�^P�:�W�ȧ[xd*j&+���82^r���[]�BZ1�7G9����h<�xPSE��H���@# �����
v��wy���d���*�DY����YVE\@i=��egJ���ђ��Wk���Y���i����Eݔܢ6�M%����0S�,��K�'/%���v��i^2Dl1}��	�޳x��=�+����t`�=B���t1s�˽�����؜N�B�/���Tl��f�ۉ� ;�������q��J�P�5���8b|WR��������]�i�y����i�s;%n>���*Ѭ�嗭� D��<�I�*V�#s`��PHTgV��2�5�e�0�g��p���in�;y�F�ӌ�B^��dhgaD�}\2ڏ]zq�?�{�{��^���DiKqB�X�2S��IB�Z��:����`���C���%z�-�@l����eо�R���'NN����fʹ(h��!�S*\Ø�mmd0��E�m���)b.\��h1�ǷI����]�wp�]���j�|�9�7���+:-N�N`^&Q]3iV���2�N���x�d/^u5��(��ΰB�F*M����ޭ'g^G�'*K]�h�*��s�B�'�l������Н�g��A �ƹw]��ݙ��`�wW"I,��L�1(f���BFBI$��1��a���K�BFLFH����m�6 ��a��Q�G���	5{��ȑ&0Q��.�GNb�ݔcY);�i���@&W�҆t�2MC����L�2 ��Xę/.h��&	��I�k����Ι3����둚E�9'v�s���ur�`�wX���"%�&�-�!���̛��I��̠�<����1��0E��s]��1&�˥͸n�\����L5���3c^�y�f�ؐ�E��UЍcn[��"$�7(�m���,F��T3RF"��/o�������ۯ=�y����ⲳ�+�x������&nJ�q���%�p�>=�z�njm��P��o0��H3��eI{��4�ci��lu���ֿH�eD�H5����K)���_���j��5��5lmV�{���}��gFL�ژ���u]�K�x�;����~A����8H"��zF���a{��"�@��c�7aV8��4��y>Ov�i�
�r�����ե�C�N����|�Nd1��H�B�'y"����z*C�+�[��m�U!�������G��
��8Bn��	�{УN`���;~������2e�ȴ��T5�R����8�`>��y�kW��kv��Q��+&V]���o6��*vm�jVP��2�j;��ҡ��sh/N; 8�!æ,�����޻���p���OM6��-L��`�B�䠗�{��|n��k��?f����ES�CO*D������vx}��0��@���?dd�=ޛd�Jb|�:�/�Ȇ�x�3��v���}�w���皗��~�`��|�+�ƈE�Cξ�Nç�͐�Ћ� �=$;�o253=+�W�ջ}^�p�=+�I�m�X�;)�w�X@��\LJ�/bv3].2�Cq����v�c{�Key��$��I�b�)�{P�Y�-^���Ai'�7�`Й�����g,~G%�������&}���m���^cX,���gw�Xn`����
v\�t��UKw�����d=&VY�U�mJy�gh��R�;���n�;ˬE�I#
��!
Ȫ>mYz�`鼧+���Ddx���h !b	�9�ߛ#��VN�x绤k}��4�=�Xw������_�r���T*���h�l�%}=�	v������y���N�j})�^��.*Y�� � �m�j(�͊N�z��_��:�|�72r�T�oN�#!׈q�k�\zPS8�,��w���yB�Y�.����U�0�ş����XfG���zF'B��'�"X\��Hy]��S���'#ȿV��<��ZR�n\]���p�����p:��~��7Vj~+Ś�0K��A/��;���.����T�ƭ����{b$���E2��&�}��mS^��2l��Bv���k��P�4+ٕ�m>v�t؞����p�R��E?��WU�9��Yz���a���s�g�xٗr^�쥕Q����AP�6�^�.�7K�(���<�^���]���0��1S�*r"���mI^wS�������_�[;M��O��w�e�ԍl�%�y>;��F�����=�������C�}0��BH`�D;'�Bz�s���Ơ���=)?5�2m�/�_��l����"�m�8�j���d�r�65�1c�J[;�=�����$��©0qZ��E�yHœ�����_]d�g��(Y��jG�~�;l�m锶���j�]���8tX�W(.�]�3.�Hن�;�橶]����e4���g����?�������d�m]�}����wP6-ݙH�`�83������z�����"�yԦ"�z�5�t+���[[��
�WX��\!����:Du��P;G�^��x�<3��4��)�(K&��	W��Pw�<��[��Fi� vW�b�)�h/aޗ�P+���Y_���P���r�������Us�������������w��]�H&8:��<����%ު�IuʠOIk���zy�!M�Y�%Չ���s�z}��L�G��%6�5 ��i��5�=�m��Tt��jl����2�T�KG �<ջ>�\����f��^֐q@� Ŋ�!���h����j�'�����+���b��?r���1���(!��P���TV5.��=/&b;zb����X��W=�tS�_@��$ֳ�1ְ��m}V�+�����Xs�2����M)�L�h���5�.g�t.#�n��b��ĨR�T�SR�j�NVì���Ċ���Y�`��ƩN�_^rf�\]��!}	��� L�ߌD�7�Jd�
��Yv;/������a��q�Ɣ�����fү0Ok�V�f����wM��y�B��8���l�jG|.puo��ȺYs�������3~��	�ߌ�[���%<�+:�`����i���tsz/��0��n�R�W�<�A�5��*H��Yc��3���c�gNlTqǿ����a��T�MɳCAM���Hx���陵�0�T�<�q^�E�4�cq�e�wf�{��O(�y�s{U��npB1��?� ���!���N�ʔ���E�g�����{�OMT�H����Z|�(u�ޡ_��r��)9�9B��B��eʓ�L�7,Wl�v�ǔ;e1GfhO��n5� ��!x���T�\�b}t/��N��-/{r�ݶ��;��8嚩53_�q�OM#~WAi���Lj�Zz�������7h��_�w����_���B�V�2�Z���П�h����D��ʅ�������hy?c�bw�u��?'4%K��ΤÚ��@�.��E٢�q�nj=�׋�g,�g�c�Cv\Cr��Y�y�I{�������G7���K�N�z]�p׳���������'�2�p���{B�dx��� ��'�X�7HQX���I����?hy��Tm�287��@��!����6v���|�ٖ�ի9�G&[���D����f�\D�\H��I�ME��^lkW���0k0�f���9�[B����w�v�=R���*;�D��6����W��Iu���!X�lj�)
�e��q/�1�S��N:�ί�ٸ+��0�K8�`��n!ۄٶ�(���B��Ym�8Z�jblwˈ[�����Cl��ԓS��(��f9��,�tB�v������4����p.U�CQ5�q�髦.P�x���I����sR�j�j=�1jđ���G��[U-������R̡D�:��zm�����`�Կ�I�f��eo�f��2w1qȲ��4�x��+fa�oA�m	���'������ƚxk�e/��C��P+� �5�ə2[O���|�L����|��z����%>��*��jR�^�zጙ��ʇ��W=��-�y���ÖbfP
�`�:{୔8|���[�����nc;�݉�U������8�s��"���(+���j�����x�r�r7�O�D��+l�r�(͇pc��◕���.:���<1�Y�vE�\��SAQc�̜1�~=S�����_3}�N6��|*Sۓ��� W�h���U���-?1NX��S�5x'����!�{��6�X�{kn~m�[3}U����Vܕm\���6�a9B�Ī2�-Gs��#��,��%���d��mH�`�tv�ң�[L6=:��n]&�[+L�#е�~�sJ9��3ly������U	���b�ئ
6��Xы�����=)�� Q�&�T�&�2Ut�T/#�hS���*ܨ��Őx`)X�?{����=�=�>��b)`Z�nm�Q�����[�պ��κ��*��3���ܤ�D�v�8Q^G��)�
RA�ME��U���]#��_��C��� ��XO���kW�����_t�+��1L�/hǣ5��{�S��ʼ�|���m�9r�h�������c���55g��	�yuf���?|�L'f�[ɷ{�`�}cu���}��m�DS���|:%�r�Caqb%M����t�_E񁕙ջ�Db���9C.��4���C�go�5 �o���T?V8S��a��/�&��}-X��e���0ݎ�b���#Z�̳I�Xu�����ɴ��6������#7����o�pVF�[:5�%�5>�z�8ǒ�m�Pd�)�b�$9�l�z���P����̍3�X�e=]�AŴzâ���U����w1�l�r�5yb�NM�\fl��l�8����xq�Q��6?Z�O�ZĘ��09ar ��� �����D �G&kun�=N�����QW96�a3LT�M\���Ɗ��J҃���"r�S��
��FM�J���L��Sg��:��A�$�G;�D�7�E2>�F�[>�sk�\/W?�1�&���Q<�/�*׌y@�Ɣ>���p���`�6���x�'.k�Y�m�'JPF�k(jŚ-J2�p��mԥsZ��v>�����v�p�R���^��#�@V{�7Li��X^0a��m� tS��k�� Ž�&k��I�#��9ܤ�W�U[��S�ؼ������d(q��RO�"����"����1��#Ͼ{a=��V�CI�x��48/'��@OOY�M)�aR�'!7K����h��R:��i��Gn�t��df��\��P~L#X���r8���z曳��W���jF����w>\i`�Y�:�n�3d���jC�5ċ������]���}S�+�X�"��V�z I��l�o�jb�W@{O�x�R��͟��`���~�NݢݤN����ˈ��ԉ��	�r�ƅ��]P�]�,�=q��9��
V�[���t����sW����v�v�jC�<x�LZa����<����SC��$��{��ɼ�a����
 ����px�C��e\7[K�~������YZ�܌�g3u���R�&1?X�#Yޠ��s��դ͗l0�[I�'�DYz����,��7�	`���V]}�=��I{C�hx~NpON6ۜ���2�'���Sl�R&a�y�7n;���lg��3q��7U4��x�O�\>��,!�u�c�Q|j����حj[	-�o^�k�}��8q�i�������o��R��}g��\�:��͙BdI��f�v�E1Y��3�7��tE� �ћ��\Xv�nVXZO�ţ��a�G�Cy`Xc+���D�_1jnI{�ʽ��ֻ���qmZ]
o�e;�r/�9��N{6ճw�*T{x�:��X)��/~y8^�9�ޜ��}ggY�fͱ��Y^Pr����0?yO�f*"�9?]���*��6f�~��q��_w����7�@�^�@�4Q�g/���T\9�����]Xs�2�s����p�g�	�t�b�ނ�k:�*b˦,�w��B1I�%"Q
�0�]Ql{�.U�3� ���i�3�{�%�����ǖo�����̳O������F"S�)P�~UE8�ئ=�І�B]��DmCbo��v�0G4��8}rWC1��˴���&X^b�sȢ�Wök�l�=K*8'��Q�����	 @C�cO��O�= ��0��VT��I�#6Ⱥ��Տl���;ɂ�qi���{ye�A�ٮT����jG�{�u:����B��a�¸��n��h:�]��`��,���o)`{���{�D�i�cX��!��Ş�����9z��b��#懻�{;�� �)�w]�TXW�t�9��*�^�-49Z	��?�����f��+cq��xvr�y��}���NHM��F��jéV�2�Z�䠗��Q�%u	����E��?����[�s&����Tɛ[m?��WQ�|v,��=|osy��鶊��Z4v�φ�]��@�w6bo3w2�ņK��-��4�Ml��ӭE�lk&��Ok�=�Y�Ue��� U�*�-��5�Z�r��p*�|�T��ڬظ�8�ɿ�Z�eԯ�V|-Ϳ�]2�bi��x�W���,��!۳�E�5)P6t�=�� /y���ʧ�P0��߬��=W��^�����I���ǃ�&��\ȊN�y��9E���,ݎsx�B���w._D^���6"ؗΟ5����4<�@��~zE���O�7�������R�w�8|�7oW��O�~����0��U�6��\3X�`Je�Fd����Q�'��n}��P�-go=q�\f���r礲B��o��S��z�X:)���!�a{�n�s<���2������К�j왆���H\����2�}��ڂ��d1q�_V�*rԨ��ߟV��O;���G���g�a��6�[����h�L�,T)=�Gh]�����6�^	��}���3��oxr�xd�;A��$����HM�x��Qͣ�	L��Js`�LJ���N��ͼ����ݻ��<���n'ʅ�J,�}�D��=� �ƽ:fRtbK#R*�p�׌�n�-�ڋv>���IL+ϱ\ᮢ�ch�a�$D&�����k�*=��}���3�O�a�����rq[Y�u��K嵖�cp�T���T��A�Y�	xDӷ�N;��>N@�	�9]s)��]_�z���=������r�����tu�SCD;��I�b�~Ȳ��^�s�{_S<�ѱ�&r!r�ȶ�5���R�s���kɯ���\Rr��]/s�2�b�uCu��r���*/���8`|�ze4F��?eN�n�Nq�P�+�.�+�I�U qWK�ȴ��T45Jw��\9����S��ܙ�nr�deט��hd �M�%M7&m�l&�V�Uz����*�AfT����
��Y�Ɯ_�M��B�	u`�����Bvi�\��N����t��7q�����N�9��H����tOZ��}ÐS�����f�&b�ޛe~��S�OO�v�v��<�0�E��'uz��B3%�uC2���0���軴k�x�t�ٲ������m��t>�^��=: �G�,[=�!�Ϻ%�r�=���˫�����ztԳh�]F?;���������y��լ!����8�$j��^�T?VD��Aih����u$U������^��}�#[�nf��d�Ie(#&<�M��y��8��-nB��y��{����� � �|V���	S��_�fq�rT����2Y���v���|��i香v�M4���F�|��w$���W�J��yܿ��¯p@��3WN�.��)YZn%�)u�c����� M�u����X2�y� Vg[�|��w'.w':�u=�l�eX�	l��w�煗�2�y��GB�Lܼ�rH:5)Y݅�&4���5S�䫛�/rgt[t]�,�8�5
�g~+07�]M��"��Z�7c&r����!.L��P]6k;�_.ս�.�P��Q�����}�f�ota�
m��.X����z�̱�E^s,E�Œ��o,F�2$���C��Ff�a�������Hn�a���T��W)�%#��yۂ�v�hRV�r�qfn �vUj��E(��^�쏸R�?a�)S�P����9�����DP�h� �k]��zУ4�t��H�+n��ߢ�v���P�X���l<�o�������>t=P�J��5w3��������f���1�b@���eH����҇-"�mޛ�y�D�uoQ]�ۂG����+�%e�\c����Q2��O;�e��C�Cj�R��E��֜� ��1}R�3�
f�ݳ�����Փ+�5I]X�n�b�u���uTq�%:*ͫ
�p�dO�C����.ڙ���F��F�f��]r!`�{�e{ժ%Y����mG�ѷ�(�Y�����3��������}�wZ',N.쮫;o)E��b�vL�wl{�@��59:7��aZ�-]7r
.�!�5̩M�{�cV�*n�C-=�(��8�g>����Ռ�f�9�<�U �����xz�Ng+]��"���e؇(���z��E�#wO]�&gV=o:�5�Z�l6���Z.ULR�peQ����-jɸF�7 U�,�3�.=˾z��霴�������kl��m�<�kF���i2��KHU�:�E�=nd���e9Lo�V`�^��2�\#L�Ae�,mGA��ly�n�Eڈ��m�vn �t2�&��nJK�c�����:,&hv���Uv�w%�~�)�C_][�	��ལ��ز�ּ��/Vz���j	���m%�ٻ��H�����޵Z�uWD1�33�����zOWL�,m��E�w\����M]�Gk�t&EȜ@Z�jY�����`޹ϓ�`��L��2�\�T��K�6C1�/���BŻ1Ys�&w*2�b�vŋ�͸�h��q�f�C�v��ͦ�o$uk݄E�I-X��qd�j�6��wR����T,r� W��V��gueN$���vz�LUVX|e�򒮂.��[���gj�f�Go^R��tc������S����\���8������;B^P�\��wz�я��H�P�|][b�2`�{0 .YF��ohN�X�*n��+��e�Q׈͒8�`�OBs�.�l��.���rKΆYØwn���pm�2پL����n���0j/	:��(ѱ�+�ْb��ƍ�W4SJ�Q&+D���cf��I����X��[ʹ�
�&��Q���D���uwv�"��@b��D�ƃ���0k�y�����F��Qj"6LFLh���	&h�h�����Th�k��"�cJd�X�(��RQb)6wn[(4`5��*�owF�d�����H���M���D&�d1Es# Cx;`0��q�ހ{r�荎͎�8�x�����8��k$�[;e�u��+][����'�c�o;��io;��:R�76�¾�W�	�*<wR�����^2)�08��a�y��O
��	l��7���`r�5Cxmmվ��)?cVg�z7'���=wG�1 x��o������,.b!�.�o1�����������6���ks��sר�p�b[���)�JT����|j�Ξ����<�Ȝ��ow:Ӹ"k�G�o�7��!m��d�'�b%9�5H�EA��h�#���ү  w�3�_ �%���O����F�z��	��ʼ3��)9*�)9w��P�J�W0��M��;��Jވ�6b)?�I����$4G��띒�:m���R�"�6�����hν������D���l�J&�gp��v��#��/�!�����|9z�\�=sM�3�k]���ͨ��j�M�T���o6������t�S��Ѣ1��x���n�vOƄ�
�V$Ȧ.L�T�P��0ɞ���2t;k�u�ҧmK�?}Q���k���5�P�?����@������>by�p��?v�Þ���@FO0TƲǿr��uɊ�-��:�;w;��π�L[<��L�1˗�W�s!x�ࡴ��~'}5�]{��V�ꕬE��)r���M�١�Z8
���]�\#��Z�����xgd����"ٶ�p�M\]ݭs-��-p����9��"�)%���U�-���t2�nv^tK��%�ɳJ)�\���h<�M�m��V���O����)8%��aD���1\��_��j�;�F%���]�&�Vc�_.
ۅ>�0���dk#~ޠ��:��]����I�_/�wXM־�W1���޽�/H�ڙ��I�2�xX�������m�<7�זe�sǤ� �� ݷ�皓ő7;}�Q���{kס�6��b%c��x<!�V����?ӳ5֟jX�48����SO�_���+YsU��Z�z�'�Q&u��l�*��Ϲ���q��y��z`�p	չ8q�TL9-d'�k����@e��^A=�%�kY��[�Pʋ�6��P.E���-v��/.֋�UNs(������sVL.~w!�>�ފN��J�QaL���T\:��{�n���Lhu[|ձYʂ���h��v�{,�M���tBd��D�6R�j����#f�V`�#*:U�MS��������z=!�v�.F��_K1 _v�4�2��|�(�d�`��.W��o�������
�d�vl���!ƑB~�= ���0%�*���H���t��EYq�Tb�$u�ߏ�������B3���V+��_uv�2��ԷZt�)��We�y�g�>�Gk�b����@�q�1��]�ga��e	+u�	��f!Ya��0>���bTe���:Vc��
ܣ�m��Z�8�LRx
�����K�&㉸��42��r�x	��b-#N��s>���-y�!����9�'(Q�����nK�=�]�t7�"Ð���Z�B/%E�����~�i��Xv�@����v�(ͅL�ޅ��⇫d��,����%QaB�O1��Z�|^�>�{p�3�����rY�:����#��l�a6T��C8еn�c����k�PK�B~`vDW��s�w���R�"�,]�����8��f\sH��zv]���u�R�O�t�=�a�r��澊�a.۳R��ɮMo�}��[��a�ɑ.������3����K�N�z]�}�(���$�L���3'h�ջ+t4��ڙ��_L�7C��ŕ�O���CCϒ/��گ���T�X��e?tu��{��:P͑��PiD�4��-����Kp̓A�Hi�z�DfJO�r�&|��D�>gom���U�[��7���<�vA�Y!
�&��q�髦.W�)�0A`�g�v1I�BsF�Z��v�|���Q�J�ʩle��8�1^Y���?q���
�������̅ܼ���}��ԉY_��Lѭ����ۏnp8^5�X@�nڱ�j�}���5��ɣ�;J&^�W��
���5�d�ޮ�����Ř��Է�:q��'�i6�	�۬ڕ��H��YR�JV�Ӽ+�9M�w��1\G'��S �;\���ڕ������~8t5�D/#�م+کnj�E&�d&T*�����]g��y]��Ő���к��~z��V��Ol��,!�p�����O5�%2��%9�ۢ/�v\Te2.��m��^�dz�̫����ƻ�o |���Hqm �A����D�����Y��f�̨�Y��?c<7s��ģ<A�5Wq�V���>d��߈�*����՗�*&�V������@C�����RtÔ�.��X�]N�_�λy�6�8T_��8m���*sd�����>�yu8�w穸�MЮ�����t��i���xj���Iĸs�NG[��sp���U١��;��&�L�>���.���s���Uz���إC��dg���\&SD�F�Zm���8
T>0V�ǘ2�����j����қ`��Jװ��O�K�LDI��X���vyS#�	�vB���Ø_�+h��<i����tI���cK�е
�d��m��=��k \��ؗ���x���y���'a���bQ����U��IW�����nsf��=���k^�)���ۇ�w݉A6�X���Z�'X�v��ʫEqwOw{�E�b�R�{�5ڒ3�wL}�l�z)wPC4<]$}%p,�<~43�Ǔ�C�����4��1��4��C.������Vk'_A�����'��>���2�y�'��H��\b�t<�l�v	v4*%�,+C�pT��(�Qޚ�D��Ѱ�zv19Yƃ�ͬay���@"I5[E?���~��,�{�[�ꩂ�GCd�h:���Za�<s筞���ٸe�tvIa�\�50�דi��Nx�H��{���{w7�&}J���a��g�)}`J��=z�g�\�3u�W�M�-���4�X�(���7�6)�{�%G&����t�w��ڀ���.=<+ʫ%{Q^�"���'��F���9���w�������C�y�����Uk~c ��e�"A�;dv�{z�0�UB�52~���*hw�F'��ܥ K"��v�7ش���򂕤�c���`�8pM�Sis����.�0+�H"E������>�Nlj�L��Mmb6皃�\:�tzs���©]�[Q���&he��,�S����Y��rT8�z�$��S��<�U���5�.�m(��q���t�m�ۗ��K��{`�#��!6Н�՝6Ԟ�.��tڞ�(���<�]����;��U�zy[]XwV�c�G�{�jE��?<�s�Ֆ@ʷ��m3e�~n�ksm�������R�H�,���]��2P�S��;+zC�뤘RfN�1v����vg$��]�/��z�R��V���:���&�t6v\�m������L'Ǡ?O�E�2�F���� ئ\�=sMל�Z��/+2�{�E�R����:2h�߿U�Z7�����ċ��c��"|���W%���-��'^�'H��������f�O�cxɷ�Q�5R͔Ż�n��C�?�v�E�˦V.NU^E�w�=�5k�'�+�fеa̦Y���-�N�	1\�_l?�uv�vCC�8�+U�+ �̽����Y�X�*��r�Xi'���{�1\�_��b�8B��X�.f��=�Z�b4A(��|o�}s`��f��A}�8;�r���w/`�R�gN��@{_�@��!����b{L>O����-�i:�ON6ۜޟ@��L�G��-��M�ڬv5�9Sh�=��2��^�ͼu��``�AU��ǇڮU��٪c(V�滞��/*A��?v�x8�~̒�!���z͛eY���K�X02FI�1�Ϙ���x��yc�;��%��j�	���a6�1�
5��c��*.и��>�����+�|�&?Ld�&V���NTș��FO�+�¼��ə��v�}*�	�Ў���Z����.W;�Բ����-�e� m<|2�jn�o����/�Y���OT��Ŵ��7;NB�fU�\��d����V_vTű$HiR�B<�0����٧�=�-������{��!��
%z|�z9�����ƾ��^�C�b��ĨR���
j�@u�7EM{/o�}<��q*W�w�r�w��]�ѱ��p�S��f�}	�oD&I˼'<R�jª)Ś*mC_E(x��o����o���Yzh()��zG�{�dLʯ�����.Ӧ�&X�LS4�i����P�5E�swvr�z�����[�� ��!�O�'�^���UeS�G3 ��u�&�������K�Ȧ�r���E�m��~g�`��0Z�5�=ʺ�y}��"�2�}���|'s��u�D�n�aTJ疡j����>�i��(yD�c��D u��{�/���~Q��J�&�h��!-Z�ӑI�*�KC�8��E���c2� �֮�E�y����uy��'�>� ��:��G��0}niT'�sm��Ze
�w��贠�ƹPXJ��\pv=t+���Gj�n�����w�p��g-0���e�3���)P6�|J�GM�3��M&yޭ�w�=ܵ���W:X+�>�%����
[K�dG�^���ÔX7��[ ��Q�	<[D�d�D�K{��9� Bm�
��̧���l����UMc�iA��_�ėy%:�Z*�^��M�;C��Gf�0�;���S 2����q�[��kE']:���m�eV�G���4�e��s:S<��H���g��h�+��Wsg7j��ۿ\�}�,ݏD��Ls�[9y�����?hy�O,"����\��e/��fY�����]�K凝���Pi�Jep���x��9��(E�F��n�j���YW�1�̧���ؽ)ߕ��ch��yj�9�,��My��)�P�k�Ί�����k�P.�����oEc߬{���-�۞X%<5�#6{�ǵ ��,�lG�>�S	����HC�w`�q��QR�g�#�F	����ڂ��J��KsW���m�d&T�P��s�ە�����������=L,�m<�53����d�I�&B}}^!��so��Ȭ��+E(Yw�4���;��1{Xd�-JJ�W7������C�d��g'�_l��%c��n������w2���,���cEL(>�s�tߖZ\2q/�O������lʝsM��p�\�pK�����N�r):a|jQu��)�b�v��-N��8zc�5����g�`�&ì��z�&ne �T��6A�N�{�t��i����N�ܜK��7���9[�*c?+3	�%����������)H��!�RP�(�Y�[���Ӥ���	�P�B��n|�-��c���
��Heq�7J����5-:6�����]�in�ȩZ�G>19���4���`���g���z�e�s�	ہn2��&��F�EM�s�O�Y���֬�J�p��N�	3la7"���ը�s7J�s���DEN��ԋ4��ۈs[K�G`8�!���G�:�ꝚmV'����	V0��J׈�|�+;6���j�YG5F�Ӫ��]Bv�;!t�(p��H�I��2��zm��潊I���2�Dlgf�,kX���c�O�^��j��b^�#��I!����O���MY�l� �#g��/�k+�.[���e'�_�C�"eq���LZ�X�c��1aO�7�͜9+^�;�^�`�!l�B'esؒf�9�4��0���Hz�Z�����?i6�1���*}f=�3�����^�����{d^9���z�4��i��,9+���dÇ��P�{�kE��s�*�E<2�yg�顈N�c#)��O���fq��S7X�(27(��	I��}��;��7~���4)��@�����\�1���o��m�Y/>��Lj�����f���൹2C���~��
ј�oV�^�o����,.b!���J�:��[ߊ��ѻ}�t���9�(��\�b���d�ﱄ�i)�%��@�<wvV���Ev��I~:����q]�l&H�u�a�y�U��C'.�u�%D��&��G �EdE���l�$FU���18��-�o��:��z2LE��ԙVgu��7:y�.:u��A8�bY���+T��	�`���n������"��y�dWX�����7��J^BАD��E�?D��(|"S��S*(�kk;\��ظu0�d'�T�h�X����6��Y��d�Xa�- �q �*I��Rr��J�b�a�l5�@�iUC�k�=ǜ�����Bm����Y�mE�aR�6�=W'��.��ֱ�2�Z��1�Cv�����y��z���[�#�Lk��@�}��	�(�w����Wb�\�Hɕ��j\��*̍n��Tw=y>;��b]�;�Y�J �`伈vOʽ=B�ԓ|MWC��f;�GB���k�R��X��yU�U,�Cb�'f�����~�'�Y�줱y��ϼũ�NC���V�S�^5�=�O�~3<6[������ �����L��pz������)���B�*:|��OR/��hGVI��23L( vP��[�9ez̋��uR̕����@w��� h�gh@�i���nvF�W�A���H���v�s1�!w�Ӗ^�4�M;w��~߿}�br�,�6ծc®��GaBE��.)*y�z�i�RR44�nq�{���$Tڱqӭp��؈�!�C;��á��E�5����K��+�Tó��Z-#�U�ԗh��;��!��g�A�VP���nhh��ۆy�s�����s{��5�+�A:yg��˱,u�s��lީ���:u���N�J&2�x���ۻ��R�M���r�,f]z9�,�8ƌ�]9�2�7���z#D4������J�ω'_v�5}�U�37�
�j�ry-��+�{�YƸ�w���V�61�׹{�R.S!!��[2�N�"�*��a:��C��U��Ɯ���g;��c���:�IW-���Q�8j��f����7��R&N�(�bչ7^�o��lֻ�^��"ِ�DS5�Fإ����~܍�-[K��[�M�r�p���F9�q�}�4�����m��֭0��_a��*̢T��&��r��Z�ۙ�j�(e�����s:�t�jN53fM9��魏F����P����wk�7����0��f�j��`����l���)�sD�md�DA��kG�O�CJż��>����s
\�>��:��i.���j}��YV�rpn)��/���,�(7 ۂ�`*[n�ŷW��}���"��K9�mN<��V�Ж�S�$�S��M�����6�vM
��F�<�F��i}�-���3Z6N����Z�k�/ASS�:�$Ӭzz��xzn��n�fZ>^{��9���Ra|U�&�|f��߷vptƋa��#��������+
22��cz�c$z���(.�K$Ҷ�X�k��'5X�p�I���UiJ$���6�mA��K��Ά(���ܔ�];uq'��9ݍ�-l����c/��UsH�N˯�ڷ��ͻSV��Xhn3��j��P���)v<�e��9�E�Px�[�weކ�-"�-�J��]���Y�Z����.�շT�EVV�0"�&ؒrE���s��s��z���+k��Z#�����e�(���:��a�WFt��d�5.i�l�����2�]�m����Q_M��aSw$�WQp����'c�cw�ڦ�U���=�vI���SCU�&� ��7w��9�a�`���q0(i�ۓnB�+�FY5u��L���J{]�s�0kq*̳�	4�33�w[�:�pǛN�F�Qو��t�����ŭ�w)�Y���R;�Xc���6�?�S5־�t�Vrok�����۽Z�'&��Wf%��G�S+�j�����;|�5])�h�_h������D�Z;a��+a�q�.��Ä*������f�խAc�d�a%��RTe���d-o;wf���q5Т�Ī��RW��ޫ ��~\�QCi���LP���;0<4��`��u������?�ٺ��K[s�W����E�e��ƅ���� ��;��5e$(��w#+3X�E���QDb�.\艍�E�u�#4�(�r��Ph9r� �IE�1`��M�Ѳ*2j��=��֙2��0Y���Hɢ��`�b�F5h��39��Q�$�)�6�1��4E`���&1�DHQ�#�t؍/<�3�hCb6-˘�X�N�Ȃ���X�uswUʹ�h�L�M�����捨ы�1�����qL�µ���de�Pǲ���H:t�v_NP��ӢdW2�L��x7t��X����]��)��ce'���:#�������6�D�D ��8�H��d����3�M������7=��@�U��=�6��[�?8����:a�_`ޟ^Y�i���f\�ڷ̷*&����ն�޾�NCY1��ִ�^m�6��.#B� =Ų/Q���|ST!v�S4,E��#H
Y1b�m�(ζ�5�n@�t��N�,��w~�=)�P� �؜�=��Qq����c)�r����a�C�q��o�@eEÛp̞�̚����7o&��a/L���P��v��u�VL.~wA���N�ؕ
VRaMK�q���c�r��j��������Z�G�vTC�=��H�o'0�v%�'j��n/�1j��=�)͔�Z8�K�o�)��nw����/�%�ب�Θ8>�" ���e���CM�m2�2�QM�K�3a�Ww�r?��օ�~5Ɓ~�.�t��w @AƑB~��A}`K'�˂e7�t�Ŵn�܈f�-s0Jg��Z���Z�;5Ȟ+� ��=���O��G�Cby�)�ޕ��N�
Xe0�9+�Z�\��T$#�%<;�Gd><�|m�?��T6��=g�E��M�M�WZ<�x�d�*��\I>\ǳ./o\xcd�#�\����)��Y��ޡX�]��3���(p��r�H6��װ8���Clboh�b���W^��VVvF�@C�b��c��wX`�ZI�2��M�t��Yn>�7�bΔ��[U�[�kׄ�W:�R(�8���E���c;J�ׯ���
�5���=1�KW��S����-̠t&5=#�s��\�V8�	�V������*9�b�&��s1��*�,��-d1�;�����50if�(tSL���-��E�6�t�=����*�f����ʹ��K�;�Zr�Ɂ���x�	�;�X��d�^��u���j+3"��}�{��!��Ԕ�v=�O�Z�=�q�����ևzdh�/"S�
��jfb�S�\����٥�{�]���!�H$=� Ȗ��p�-3��M���&�F��]�#<?j��I��h��O�x��P�C���B��o�2�7C�:��m3bGZ�sw��:��4:.'�w5�bj1��eT� ���B籆eAeУ`�<��c
N�Q/r�����o����|6b��U��?0`����5���j�����ټ�&X��3Ц1EUd�[�s���Cuxunо�x�b�L�VQc����fL����C_(�^oLe4am�ɊPbcO)�s!�^�E�U�Aq>�����o��3/Ø���m�z�)
�yGwwC'u�bYz���,�X
�4(�(��;U8+�wg
&jݙfdwա~P�L:mY&��$��֪=�p�h�/6,�],Jr�1�}\ګ��wIN�i=�$�+�c��]z���G��[�V����ZĠ"Ϗ��L|<��glA���-Fy�-�^F!'\^%�u��Lh�I�>�s����'�}hA�l}�������jn�������.��ʆp�*��w�E'L9L"�x�U��ۋ��m��e�۾�`WT�"*�w���f��B9�:cf�I���%��]�鼛����5Jw�hL1�m�gM�6�v�-���'�l/o�]�0_1�F�FħZ$Ͱ-XNP�T�r-Gs�$��T1͵�N�r���܆c���KӇ�p��:Xtz<:�ꝚmW=E����t�[���9�;dhD=#���~����d.�� ���(���4wg�g��C_�Ӆ��i�p�_Q�<��Vx�|��N�{��5�f4b�; �fq��x����8Ys�9<p��/7L����x�r��l�m��E�����H��C�W�LZ��;xwk�B%C�zج����˽x}<0��\<�u;��4�ͬa'���Š$���C�?��?z�I�{Ғ��ٰ=��d���\έ��FX�B�h�\��[�����RR);>�2��g.v�ˮH�tf��M���&��ղ_z��x{��vev ѥ�ԭf��X#ef	mXy���`�Q>"r�ޥu�f8X�Ǧ_��y�Li�FN|���%��ZZP�->��I�z/��ӛ����$��K(!p�4�Mv����Z����[A{�/V�I��
�?�?/22�Ǭ���ׯf@ƥ�S7��MΓ���{1���f�Z�b�k I�C6_�b�O��J�,���/�:�
�V0K����qy.nz��'�������6$eMK�{TgXz��/���Xũ/c/�d���D|��B�a���wS��:��P*���Nxd_�Ji��T��Dm�5�F4'�|s2��_�K6�`[��_�O�u�q^ b�:��D��%���)�|��Ʃȣ)��ѷ<�QWw1M�'u�t�X�wmy���߈b2p���N�鳃�,��0�I>�NW4	P,��7�U���s�2�wr���E������P!�9�k�c�f�y���*]���/~�y�iv�٬ny�Ś�9{^B/K����,0����X(֑G8���X�r�/�������}��8�R�7�۷���f�O-�X��Q��ćO�H��
!���:��'˾���uP,Tƴ�����4���ſa�Tb�l���gQS�Ȑ���;�[(��P+]��u�2wA/Xۈ��vY�~�KY̽op/,��ys��Wz�Qqp��D��~ׯ���}q��)pO�Օ�Z�[}f�ݻ��uv��yW6�geh5�q.Z���������3���gKC����_9��-��4ԁ�I��b3�R�s�UBr��D������.!zw���ɲ��mv�T�h�v�X�$����BՀ�S,��ߖǧc�u�/��!ݹu��PE�$],��s��΀�	��C�az��O��hGW��N���`Hqף�W4"���/���������ø�9��gl�\L,sY#��� aΡ4L�v����Z�Ҧ�����ڇ��Z�����ߕR�����!���^����{��r�}?Lز��
�w�3J͞�b����hD�4�|kOC�m�׶E;�e��Ⱦ$]@т)�D��X 龚>%n�kP;	㐃�
� ��Q�g�3f�P�Ξ}�N�,s[�
_bMI˄u�>���YA,j+���^A=�%�kY��[�VT\9�y<�ꐒr�dUvi��
ϰD�@LJv�zu�VL.z�kߑ�N�bT)X
�0�S�o�-|[��Wu�;�d6����g��XeS6C:N�},�H�X�;�I˼'���z��+	7�[���Z'.g�n�I˨s��YB�6x�`v�R����U��v�:b"�r�Wl|��FP�@X�c
Z\n�Nb�FK�Ը:�]ǚK�W-r��2��zu����-�lwJ��ԗ�#����J����
��=�A�����ѳl'�-�P8ސC�X�H8�F��_K17�]�f�ݥ6ǻ/U�ᘌ9�ȷc8���Qz+�q�e�;�0�qh!�!�O���ڼ�zs�]X��5�ݪߡb������OZ��"����Z�ٮvng��=�y_&�ȁ7jj�4���.�®m:�7B���L(�.yn��E��RX��5<;�Gd>>A�h��:׵u��5ٳ�Sr`���q|���W&�Y���J���]<�n�k�!����\�g�wRngnn�&N�(p�K���)�`����9=#�hg(Ze
�w'�Z�9/M�(.0T��Z��]-�ov���O�%�s/��P����_?�Ӳ��,9��R�VM?H��9���޽�W���r<�KsW��^��g&;���B���]bdG�^Ǜ�}Zqp�N�M�qa��\9ӱ����K�e����4��c�)���;�/�Z�&q�St�0�8�N�������An+z��^E��G��PiD�4�l����:�<��	;o;#"x�M��m�ǩ\�u{bK�5ԴG~�[�?n_֫1�[ǒ�zfّvϦ���K��=Y��kHڳd�Je���-::4�KHE���d�����:��8s@�NX�5EJ�'V��U��wHLݿ����b����^��*p�M��/
���!d�+������ �~�(k��J�!�"k�"�)�_ev

����e�-հ�K�:B�ň��/sQ�]~ʩlj\�.{�2���Q�L�v��՜we�wr�p�����~��g���p��cA�3�0�׵P���w׏�����oq�*���J��W=�k��ߏNk׽�V��Ol�@Ŵ��K�	���}^!�&���cr����z����ؘ��q��\:��^%9��0L���o�V�~Wk��>>�W���M}*R߆���l�.�&�W��$�^%�u��c@�I�>�s�{������(廦g��J�u.gX��o�UN|�}��7�7��E������~)�8���Jvێe+�����l�t{W�s�8{n	ٹ����zBc��Iц���8���='�⠱ɫ����X��t��X�!|����!x��zy�%�f��a9B���F^_%dƚuycks�ً[�1�Um�q�6����[��k�����'f�U�Qke^H���@�u/���[��V�	��5�V����t�r�L"N���)�:4�T:].7��7A�T�؃K��\v_M�ޯ�U`��з�?�k��k��M��Ĥӈ�K�0���@ݐ�*`Y�o�.�w��9�n�Ў9N�j��μ�5i5I��MI��m��~�}�2u������A��m��`�#���}*eP����x��*�!ޝ?f�;	�˛Ȧ(*��������fy���1�b�;7���c��&'����c����^�k�՛k_��%������D�b�t<�l��r&�����>M����jwt4:a��p�b��=��Q�l9����7��C�y�{�m߲jB��׌�j~�NN���oh%QO�C?�
!;0�!ͥQהo�v=k�Y���A*�'��G�-W�l��.)������c]/M��9���0����ׯ{�b��U=ڧ��Nǫq�h�x� m�4Q�k�m+�ua���X5�� �s�6�JEt�D�à{q�Lw�	�(-E�Y�F{���s>�gf9�c��s#�_b�{��nq�\����dk�U#(�JU)&�&�ڭ�'H��a�Z&����d��ƈ�����ϛa#�笩(���2���~�����kx��9ds{(Nn����s�\Ѥ3��^h�l�ƴ��/԰Q�V��]�\9ڼ�F*)�r�[�ق�ɽN��Ž�aA��0��wR܄�� �D�[��>�w�ʱ�=��r���B��ŹL���ٻ��{K<�Lń�K��뽕�7�ɻA#w� N�}�� ��H��ȍ�Y�O ������t9�^-��N�q����0�T�#1�[��3�[��&�7�-1��o:�x�L�f��]9�[t�#����t`a�ޘ�]Q��q1�ظA������FgeP� tM�)'�u��Z��Neԉ����SX��{�D�5���N=Ga��PM�KhZ�p׏�����n��l��x������������*}ݓz�S�����]ӽ&:N�ؘNȖ��T+r*��nLM%]�Z3:�ָl3�����xF�پ/�Q�vs���8�m	6KK]]*���{��X����:G/=h��Y��Z�!.N�L�s��m���3�����K�:(�E9�d��	*הi�L��8'�&v�i�'��@Un�1����,�O���j����oQ�Az�"�"TS�?���8����$�J9��Ϫ���6�϶��E��W�����5lv#�~f� ,R�K��g��]����NMG��Aih�vi|���ճ	�fi��G$<@������3pO��2�n�v��&=�w�Tq"⩪�3���}�J�9�V�	�dO��i��>�n���mrb-�v/�V�Db67+�p|����k����[W�6��(�H=V�M�t����CLv\�gc��JguǬB�#�-�k%w2
�FɃ]���3D��M��{���Ev^H����g�*�r:B@�#ի�ӰRWێmٶ�z����nof09�]^3Ʃ����vfH# H[�=|�A��p����i�c��ƪNu�H��>+�6�s��s�h!��.	8��yyx���z5�zp��zԛ)�ܥ4�\lsߗV�ݿ'�j���o��a'�s�ꧬ���H����A��5=B�*�])R0Wt�D?~~�=#9�/���~�8����96����G�GO*j�9��r�k��	[�����eS��8�M���@�`��?������OGmgT�^�V��	-7r�L�i��i馚zx�dU���xm��&u��z���Dԥ+:MwE����p͊3�.�T�L�~'(�<��3xj�NF,�l�ƮI[�	��v�|cn�������;~�zA�L��1�Z�$Kٻ;v7ʎwcƺ:U�������QԶ.q]MᲳ����#K2k�7:|�>p�9^r�����5��[B��d�3��cІ�"�����l@v�v1�!�'<�KA��Lע��ٓ�t*�v��eM�f�r}0�)�5� �q���#7�Ц"yS���-�e��Z��
"�	����!8M���u�v6|���6P%]oL�e�܁9"۰\z�~��U٩3-��K�6��]@�cG�N��_v����ϰ���U��,(t�����6:�v�x2d���q��O�VP����ϞM������	�h�C���a[�lb�hL�.���w��I��j�ݹ�ׅ]c�Tz�]�Rǵ"���xY0�~g<B����]%-f�`��i^�K�k�G�ɓT����ݗt�>҆�Ռ�q��Գ!犋� �;�c�����]���)A�;n��j�ب;7B��8Pg�'/�ɛF�����ݍ�p�3����c��˄��N�b��)h���Y���>����_�2���ۗ�͙۱'w���x��.��4O�(&]m�iʎ#2���Gn��]�ʔ�w �ͭ���f���͙*��˝��&�{v�R|z���Cٶ)�e$�.��8���TV�.Ky�������m�c:}�n8:�c�4K���ڒ�9z�8�y�]��k�Wm��%�R�8��=uޑR+�����r'��V"�Ǣ��绎B{�
:�o=�88݉���\p�и��N�)'W:(c�{(7e��vx����*X}�T�IQ\���ޫ䨡�H�*�V��z�_f幑���[ֺ�`���DiF�n��GC_fKĲC5x��hp<.4���{70D�E�*��S������x��DZ�Z3�Z���]SE�4>����(����3�;1+R:�s3q;-���B���LR�������"ͫ�� �t��0��6n��_ɿ���%`����C>u7j���pW�T�yb�K�r-ޑ�.P�1� j6ED�ȭÍ�}��7r��,pܫZa��4]�n�&�����{���zծ͋���6�/%�ܣJ,NM�Ԕ�;NAtt��i�p��ޭ%�JGM
�L�ǜP�8V_<Zm��c����B�5�&��i�5�P3��,�t���o�A��PZ�3�@@\����jA��& [��Q쎝����<�X�~Gx�0U��]f�3 ��t���q�b�\sv<�ie,R�͗��j�xN)*�u��S�GXx��,5z)�Jocέ1�=�=�Y�GVp*�R�~,^7ϥ��}��Y�ŷt��/��TYv�Yڞ-�NcN!Ju�yoP���	��N�#c&����i��t�3e*�}�??��݌kDX-��L�wZ��(�T�m�Œ����CDEݻu�5��9�b*��r��.Q.I�7U���s��sW9.�	ݻ����,9\;��F�C)6#&�F�7.i�!��\��F7N\湷"+s�N뛆���}�F�8[�9�j]�s\���q�7��771n�N�s�Xڝ��˻��vh���ӻ]��M�:�s�wut�s�9\�h��4[�2s\5wu�S��DZ���4�W1\�7w6���n�h9[��G+��\�;�Q_��Vp�]���?d����$z�8ļ�ARW��;�S.��)Km�������F����a���aލ�j�q��.$U9g�L%��{=6��K�4G�G3�����G�e^��x(��%/	���-�_�wz�ٳt	{Ϲڬ�6ǌ3��g����ndrzT�����|����{|>:�=f�W�"|H�q���]:m̍�t���2{//��"h�ށ�@x¨z�����D$h	$.lJ��Nqx����d<N7�{{#�'CFDPF<�;�����^>�#Q�0�&B�2�J������-����=���W�)_�*2_���}2�Z�S{�
��-o���mq���n���9��fґsN�Y�`?G	q*Ɏ���u�;����Z�t��^��9ȕ�)����4歯���FT/���m�?�N�v|�4�M}�!�y2��W�OAIUO�s��u5lᎵJ�!�������ϔ�>|>�G�*}�RV^W�=Ǌ���t��'���y�k:���5]R��1��pS/3��XUZ�u�ݘk�Twۋ�@t�#��K�ip,6���{� ��oR[6���j�3��7O-�/�����4�{�����R�b�ZY���x�5u��6��Z��PZЅ�AC��nF}���Y�Sy8�v�(S���^�Ol��w��7��g�����dB�E7\��"�ÞT�Z�4v6;�j�~-�w��&�S��!�["7��0ܚ��d��7+˞K����\g2rrf����w!��ه��D�N�/�ָo>�X#��&�7�<M�F֪���H����EIݐmO�����z p��6up"��na`=Ⱥ�bMp������'�sr�j^�~��{�1Z��v��\Z���5��\N%�f�Qb�w�}���v��:|z��A�;��Ƿ�n��_waS��HÄ�7��f�>Ⱦ'��#A#�x�I�E��af�[�V3+�6��Qa�j��xVh�Ĭo7^Y��8�%�-w�U;����8w����R���,v �!f�OՒw;`^Y:�����~���-��8wqZ��@$�@��>�vY�t@A({�/ޏH��P��k~t�I��!��?ٗop;���(�k�����Ȉ9�^h����^9�f��إ�e�gE	v�sF��ΥJ�ESG��:Je�h�
���3H����+es��2̭�+�P��c�o3r�vs:.���1o8vՔ��7��LU��s6��P�'�JڲA�t�x���+=sN�e��ńCIyW�8���$�C�!��Փ���oPR�&:փג.i�ղ��kګ*���&sz�Y!t�ކeڄ�-���T��@�)A2�5@��In��MO{fζWWn�|�d e�"ݑ]|��̀�	�z��YL�KE�랅������;���S~�<�@C!�؆Ѝ���%~�������
c�ȱ_&S��)�ۼ>ǝ��]@�����0�A�!l����������@�)�Nr�5�Կi���4�Z~�y��,���Y�����oV�˝e*gCP�ȵQا_�����eI�7:;D�+LR]һ�a�؆�v��L��8^cJ�ˆ{��;W�i�3��I�97Uܖծ��x�����K\^��e��]��4j��q�ϣ�����9+����˺��%�����&�k������p��x/3��W�k�V-
�m+qVܫ������K;b;Y�C	�bk���	sE=��(#+7�G�����geI;_$VB�Ǚ.�K�&����b�oM
WFe9@�S��,�N��Z�mL,���td�f�f�[�Ӳ�(Ѽm��
��4� �h���9�u���=e�=)�fl��)d*W�q�z��I����
&�"a��`%�Y|8�޿?�!OJ���}�{��
�p9h��tQ��s8��@�h�������GVAǯ������DH���=� R�U�s>�g�cY����m��mM��|�D���|8P�q �"B��y+-[���n�����xW�*0��c�>��ϙ*�l����[W�6��q��s��:�'ce�k�]Ӭ&0�f�&�8@�X�n�(-�rh�Ae#(�;Et���1����f��b��ݹ��8���:i�ճ� �("���	�o
��yM�u78%\sft����wV�z[�$���w�˭�u�z$,�H[�
�5�8�P)���x��y���<y����*���Cd솪s9���/��޿�3����|�6��4�����i5k���/s����C�txL oݵaJ��3w,�[�[�k��{p4W��"���Zm��0��r�ZP�^�';b}}Z����`�9c�
�;1^�Ze�A��6�'\���/��
��Zy��"��:H�3�[���e{j����e1�KJ�`k�8�l����Yeh���;�1��C]vw>܇C�c��1�/��DҤJ���,4�L�:�Vs������v��0.ò t��6J�4f�]Wr�k��|غˈ�97-Pϱe�t6�oY@�>�`�q��ހk�K�Fv��4�:WR�!L��S�Cpl��ָp��}�z�����>�n���?�;�@;6(l�H��0��6��M��s��gr�˦�=f�l��4l;�!�8|�E��}kF0(�����&�ml�F1���dV�U�H$u`��'�Ӝ�0�Q�Z�#-�0��̪�����Fl�J�e�W�����!$|D� pSq�����L"��pn_u��$�ʓ�Ç͏��I>��`��$D��������\�8w^M7owZ>t���^���	h{�4"c�VE��WG����Uo0�p�"��ebd݇&�v�[D�\�����STZ8���i;�Éۦᴫ%�wBCB�e�=��R]ՂVΒ��_-F�wM�f��}M��+�[5��de�̵�쌅w�U�b��G=��#�#s�C�֜/��b��:�f񫝛�L���j��)}?l(xS�d[���-ă�7�0�|���ux��]EV��)")Y�=�z�ji�p�Y1P����K�ʈO��`�K�}x�H�]<�)�ޔoƊT�T�W>�eM/n�`WSf�v�2��N�!��s�5d!�j��x�#X���O��m�ب����-㻶��?8"�ϩmzw���ږ�W)\P�ӊ�����n�ܽ���������S&�T����,��]�Pt,O�ml4{�z��2M劭��nz����6���:�t�/:�/�0[�o���*��;I�
��y@���1]��7����G9��k����t7�0�`��vpxغB�m+�3.N�F�=G�J�䶂D�Е���S���L3%������T�L�h=h�S���^�T��9�ޕ�c������p�ޜa_����wm�����Vm�0�3(���B�Յ&���z�7���F�vD���ƌ8M���#`i������Y�¯�[6�yk�r;91�q�y*��l֔L�4&��Cv�A����U��`��\lϦv�;Ɩn�Qn�u�ӫ�Mi��8�M�떁3WVY
σ/�0qH�c�}ϳ|��wĎ�/�xV='���j��X�㇤.�?���5@�L<+5�f�辳x�[Vϧ=�9�i9���};o�������x:��T�גo��w��c�3�8�$��`�/5u��(7���WK^\߲Y�t@A?����9L��I�87M��P̌�R\�OF�:ٲ�Yn�=�t���Ş_�X������NוbU���!j(.��دǯ.%��55ҽv'7W>�Z�����`�n���n�=��T��R��Lǝ�2!��\w������t>Z�*��,�P�EP�/��x=�G_	��s5�����������G]:�i�E׃�#ϙ�
��)��.�J2�-�psN�n�&�+�w�O����㫏Q��x�n��[1�8����1��.?�[9�]�W(���E�5���i���KcfcUӹو���p�/MӂF�&=���ܧU���� ��V�c̐���������j��W���`��FgV>E'��Į=Qd�y�����PAS@4��Y����M��Wة��*s�1�"uf����Ѽ@�-�IM+M� �O�J���-�R�a�s�Fi��W\k�.4��J.Q�5&���Q헢��J��K���m�qg�ӦY06n�d_wj�|���Ha�p�ٝ/�N�7T;��Kw���jFqiˑC�+���C���v7��$;��Fc�'צ�%u���.�Y���{���Rӑ�>�ƿmCW ��x����Ѝe���(�fL��n�cm�[v�l:ow�!��$����`p�}ρ8gU�"�%��yq]�;*άQ#�'���0f�/7�豺
�\�����2�`�^k��w|�a]�u��v� J�_��Y�J���}�M���ط��C�
�X]�i{#�s���^���r����xw�@R	����e\�nf�k�w|��fNv[���R�^hr������{%-���ړ���[��9��ִ�j��`���ݡ�s�;;�t�>�3�O%<�:C��l�dݎ��?�g���p��za��}�݈%}R�Һ��d���a���*��#�j��S��:+5�Y[X���71�z�����8��j�(h��Z���a�7FE��$�1���,}�QQ/�������'��R��C%w1
��kVZIsqٻ'�{;]<��y�OsL��Ȼ�]�)�g{����k��Yv���Iq�5Ot�n[���!e�Y\㚸bֹ�b�n�����+M�A&�:EX� �25��T��fI�R.�1v��tt�c��������J�e4xܤ�/%�xR1/'���"�C�F19y�/��v�cN�,-Ƅ�|�?#�jz��UGDҤhݱTl\L�:�n�f̢{xt��a��A�8`�V�z6J���=u^˖T]��֮��ͤ�&��p�ۯ�p�7[#��?�:��]�u���՜ec	�4W�$7��6��tƜo}������s��|����#y�!j�\i���~���ll�q�J��"Eg�E��l��f��1��O�Чu���7|�d�u���,�g_*��Ox��5}�6��l��&]0������W�پ�S�R�{
��y�3I�C�b�N�4��}N���ڗ�`����������� �M�9����eln���"��<�梐MNoF
�p- ms���xwo��H<b�ܤ^6Ei�\d��#�����4۞�tT_l�}�Y��=;��լ�����Y;�M�n��1 �"RHA�^ơ�$�~��zr���,���	���B��⋎���Vn��$A��0�4��S%����t��/�_�mH�����H$�po�1�2�똲�~1��^Eqٸ{�v=��J<A�����ג���5y
PF���3]M��Q��;}/�rb;�9�$V7��S�'j-�wV����pkʫ7P�Bio8aLjq�M�nu�JG���9�Z�v�)W��M�V6�WN���nI�3�����F�0�Mp"+xΙI_��8��q�4<�X�%�Nb��M\��{-T�Ag*<����>B���d�|�n/M��ٱ���fIm�s���p��6{<��aO�����]Y�&���9{|�||�i�Ye�Ze�Ǎ�i�DK��X��'W�Ml]e��邒��W/��Jk��x���j����u�%�Y�2�d�=�����#�b�QP�����0V�t�@t;	��üh��W=Ѯ�AuΊ�br�	÷x�6&Vm���,X�Vv�G����ԩ�Ɔn�����@޿gNٛ�7��pg�y�a �lX^v��Z��U�Untcc�*f��9`�T���R�~�n�f�2�d�v�Ew]ibX��of�Ƃ��(�q��XƝu��x%9���[�ov��Q
c ��
�S:2�B�1z��8����iw��a5i��gm�|eCr�L�jQ�iS��[�N�P��n��*ަA��:���!��Xݱ[�R�95�ʺ5nѐ�m�Y&�N�|��A%e�#B;�x���#wS�#W[#0�屨*ι�(��[O�E4�m��-��*z������֮�c��ĖM
I�wa�������ݤ��m��Of>f�%�.���9`C��R��*=r�ݑd�E����%��u��6.�Ӂ'CdT��ҥ�k�̪N��}���^d�.���r���Ҝ��K�M���8.��'/����ݝ����}J�*V�1�͌@E+6b�&8��'!��`ث���Wm��\�	m�(��HInfU�ɼ��������|`�˾ʈ�h�yI�wS��-PѢS=�ׂ��v �Xc}����4�uu̻;%�a�����L��u�}�����N�
��ɑ��4�A�b+�kL��ֽ��2�8s�4õ�P�2-J�4tL�`�#�����TK��;�<MӱN�ٵӀ�㭨��uy��{x����ۙÒ��S�ʐළ&��ĕu�d��]ʔ^����2a�r7#�R����&wi�7g9�����P�;Yz.t48q�n����`�v�r�q[c6l��l��A4e_V1Koz���d@�[�8>9!�M���p�rx("���m�V�oC����ZF��q3Yp�O��`>�q�#tD��jftG�g���jө��[�r��si+���{I�X^���u^�J$��K2�9T�O9�&DN�� 8/�]L˳�U�yL��0�uge���ݺ�Kҫ��5m9A��َ6�R���*v��ɭv7D��:�[j�e���p�K�ܲ t�Yy�j���["���wZ��71O��
f���%|`��u>��V:1�t��cWG���timoR��	�[V�R��yݬ���ﲶ� �@�{LS���j��᠏9�2��r��ivSVT�v��Y����*�Ǒ�O4����a�b����1�e�҃�������`������dV�%�T�ݻ���U9��;�ˁ#&u��@"����s��`�l��D����8���̕��Ι�����)9�b�\�r���9T��㑳�4�,[q^T갚c�4%>�^]�dK�����*3O���6
h�W��w�~?�_���s�ܮh���WW.�\�5�sr�M˔nk��	��ή��\�]ݴ����eI�ɋwu��t�bw2�����\�),nlE�];���d�b���nm�:�ws�;��cF��[��W-ˇ1�%��n��r�n��+���)�.\�������")	5ssp��������ȫ�G�
1
鱋��Iӎ�Mwu;�����sA���͍�i�E���\��\�κ�F���n껎��\-�F�9�`��`�s���똝�\4n����.�۷W"�ls���.㻑�v�;��z%�ݻ.t��.:��%;�t.s.p���n�J��ܺ]ۢ�#7�o����7)���EN��A���s� aK��ϴ�:��n��)�sL�q��mhkHLLV`����y1J��-�L&nҵE������e$p�Q$�Q8�G�o�H������^��tF�ûy���K�����~H�ԛ�bi�߽��k���I�9����lӧ�6��3���1 R�y�;��i��+�y�7��q�m}�j���XD\�s��y-����O��e'��SAL��v��sR/UEOtfÃ�DknO�MV�a�ҧk�c���eث�kK��nS��h�޽�p�l��8p�0�f@�e�/K��z����͙��u��ŧZ7�0��0t�E������_�u`F³B7��ڰ��7�<JC�nJჷ)f܂+[{��݂���c�
���K���e=Ƶq�ֻ�}ΰ�'7H׈�{�u�	D�\�ا3��,t �������ou�Ǿ��5�L"wms�D�>�B9�F�Q֑�Jn�F�=4��\"��lFAf��绝3��ɍ��B�E!\w���;����̶:�]��R���
�M���c���l��;�7���ˁ9� ���\����)�b�	��7��b-�~�.�����3�&Y㣹�r�&Ĥ�A�C-=��أW��I\77/%t�)��z�#5�r��v^i�G��kJ=�H�Q��ޝ�w�C{��P�n�_�j�����T2�x�*8[�gcn≊�ƍ�ýݧ�ur5[􊶀�'"��@^����ڑv���ų��n�	�;R��8k8�g5V�I)�R:ޡG��"����
�r���"�5�\��m���ﱅ�:���`��C^O\���e��E�!p������43û��T�S�;&ў��QC�.V�yf�H������QJ�U�bv�3��z�a}L�^����ֶ$
)���c�aJ�{#vw@hU�72�u��]"8�@01;3��q����$�-ރ),�pv�㥦�^�O�u�q�]0w��@#z|���������̝�3��/8n��v�z(�2m�u���0Aty���o���n����Ƶ�_�1׻�v[6U�����>�xi��g���W_��	S�\j�6����]B�B6yh�	R<+�y[w�yXf4k,����~e}��D��5���2}�C�x�RŒ����c��b���+["G��m�L<�.>��t��d����y}4e�9�QR��L�t��H���`#u�S��wݶ�|ۚ:�si��O5�j�F��>�x�ǳ�E��c��{a���;3B��%`�a�곷���ȉ ��){��e�zs\�ja�S���m�]�,K�7���WUxvV�x�J�'�p�"ނx�}�=O۲�m[�e�XOA(ꧨD��ɋ�.Kj��s$[0����Ք���}���;�=��p���� w�e�Y+��̺�m����E�|Zu��k����ݽ�LyU�藉�d@
�HOL��K�I����m{��g�����%~/�Y����=ҝ�u>�Ȑ�p|��c=>r�����с!��!�Q���"�sɒ�����sSyGE��;A����J;7�z�X��!>����B�h�J�L.05��[z�f�ׄ<��h���z=��m9���f����*���iR/���uj�٢�0^�;��db5�E-�.xz��+�V\��&����]^�ߊB�Mcڗ��Oi��o4-a�WZưkR&��w0nY�����*��vЧG\�1�N �2��8�aQ�e��[��9�����{���Wk�z�H�';�в���l�L��$�K���.��Z˗u1��ˍ�F����]B�ȧ�z��c�����=�z�;w� ,�1BV웭����B�o25�� ���jH<H��D�P���z�gK��>|쓺r����6|:��o�s@oN�q�crt+�ɑ{����'���EF��"E`]���h�Hۢ�E���s�{7���5��؏p^���*1��x�_?w�x#I�=�l;���R1�}�9��߰��J���Ψ�U���WF;{�I!ڭ�a;'{.�C�]���"M���i����eޒ������?KϾpE���6%����\��Ѵu:����y�T�2�X�5���a]ϩ��7R�y�S0}���}���x��Ă�td�Ƽ��l)��5!N("+r���{f���Y;�z��y�Փ3�Y�$V)T�H;W"��մz>m��0�x�C��o�z����A����N+K�v��ސn]q���a�Y�H�x��=����=�������	�_�Ѯ��r��ɧj��O�E�:���ZQ�EY�Ҷ�LJ�P�Y�Hv��z��j���k4�A�%M�j��`�{RI٦���u��O�9ݍ�ς��R�AB����΂�5B�JU�%Sd�Tau4�s[J쌩=��g݌�@WHɇJk�j�U��i+�xF�O�q�^�5�H8�wc��ov�^{���O��gT:+jw��!G����%M,�/����)�6[N���ǝ�/�dv�Hd��:;pY Fj�ι0��^c�]�v��Ǖ�kɩ~�}��EF��!s���ǃ����զ���<�F�w��r[������VU�H���	�6������!�42�㦥�2�e��*�s�!޸M�sM�$��mMEzS��䀟v��SQϕ���KY��'��F�Í)��+zQr�y�ޕ��Gq�ۘ5��N_[F���<�LF�!�f1�H�/�/����ל��9,�,���j��*��]!�]��w@����^�����`t�5ө\f �H���k:\2��:�u�R�#�����̍�]mlYΧxf�x;�D�m��v{���j�]N��w��5�s	tX���15:V�z+��W3q�Pv�0)�O���ٽ]&#m;s��|�p�u�Xj�5I��.o���(B�tO�Lcǹ�݂��S�p��������`ﱍq4�i�[������j�w&�ӢO�ymx%hHD�
��*ٷ3���R�~�҇�w:@�[�v�v����Q*v�{!qB��8�4GZsi\�Bn�B�i��u\���^T���.�Ƅa��|�j�ɍ�!f����=�ojD?d9F�7Zv���|>ɧɠ�uEW0xB��,���-AGK�s��ϒ��c����ȸ;�s�V�}V�
b&�Uz80/���g?���aQ�ݚ���f���-�v�*�UW�j:���x[$�HW��ɾj�
������my�%c�q�y2]@��l��u���(��-$��ɽʨ\�*����ŧ�P�R�t,���>�n�$�xj:]�r�5����F��z��z���[R0����p�-�JUu��뉍��4�آe��,��o�:E��nLt�������Z�T��I�C�@��wy��@��G=x�Џ���*�f4��/f<�SM���3�n��h=��C��j��(���/.��oB]Y�&M�a��q���b�X|����{FL��dD���n���o��b���\v#VG4���ww����E�11/�͝�n��m������k
p��ћo0H�wd��J���t��r��B�)�Y��[�\��H�:�w{}^.����k-�Qoe��}�{�aGi���t��ɟ�z��ɠ�:�s?�&��7Wl�;4Ji1��ӳ�c*����`�d��J~��3Ώ��o�K/�ޭ���F9;���я;���^x=/�iX�1��"$<#<{�<9e�l�w��(حiɻ-���6!��R��F�M]U���ԁ�q%Y�[2��?A�������S��ߧ��XOA(z��,,�{&*|�-摻9n�-�^kaj���kT�'A�TK����ň0�,�^k�XcwR�C^�f�=�����x��d׌�=y>5^�v� z PE�_�!W*����9K�r�νk�1�Z�:�;��v������m�\�=�'S$�͝�oPxG�y�\]�/Q�FSn�q<��1N�-3*m��ܹ�]�n�Wh�J=�:���0h�yM �%�w
2�����6�D�7+�q��K���ۉ'2��&W�+�X��:<RRc�P{��N���R�E�e��#�o���)�\��d_#¸�t"o�"�y3��d��;1UƲ{_�o�7�i�#n8!���cs���j�U���r�yt�65�3Y��潊��҃�i��n=s��l0�	e���煚��J{�������l�TA�1�wnϯOI�u*?W��Cp�l妄l�@A�>3�X���j�g��}zE�*�k��zV���zXh������Jחw��g|��x~<��1��}I�R�VI�~�2�6��q����k��J�\?^~��oLN��,�`9m���)�&�uJ^�ۮ�O?J�'����O�,��&�6����x0k��x�4#)�l�Z��"A#�GZͺi�w��\����՚��J�g����f£Q���7p�� ���kL��k��m�z�ڡ3�d����Z��N�Ω�:��K�^�K&��	�f[��!p�'���z7+���4]�(�g��޾�P=-�)1��Tw �iXʉ�m�E�����v`�ao^Uʍ3Ŗd9�aV��g`�#g��և�f�fby�!)��ח��1Y�=%1�ם���	�SC����߯�:�ۊ�ܛ�6D�����R:)�k�� wB	C�����f=5s����Н�}=�VE��[xPRђ�o)H��3�t+�3�wR�Í�c��4�8� :�aU영�B�)f�=���EM9[O�
� D��E�5}�ky�wz�N�B<l�	���dj���%S4�0�g5M�YJ6��w��=4��
���"s}�L%�}៼ 7�]�c]5����Yo�)	�Ú�g�K����*��7���!@��8T>=[C�9p&I���%X������鰂��#5w {EB�T����1��w;.0�+����o�����W`a�5�N3����W3�uѩ�Qz��ү�ud�.�����6�M0q����/�E��d�3A��}(��l}h�\R���s�տ��[gsR�xM�-t����yu3v�v`��]�\�
8cP7x�V(��Zb����e�CbT�][ڙh�,����v��N�uT����Vh�y�S�(�Sұ.���u�O}=]�Mm��0Ϙ.W���Q�[�NKh��76)9�s�\D�W�(;MG]zw�y��7�@�1���ޤ�n��ҧI��p�U���Nտ�zEo8�NvX&C6�i[l�2��޸1�<�C�e��Nu�N���5<"��f���RH�³Q��څi��xX~�F�q��"7�X��x�`�#b��d3���rmq�-U��)�noftʍ�#-Q�/z�Ȍ�<��/t�lS��fI�n󓂆��֬��|wfw�8h��q*z�c$�B��+�(�O�i]�
�Ԏ���=Vfud[��A�q�\���ҬJ��;�-�PS�q���CZw�Fh�=_��h�=��+n��~�����.�n�Y��G|���Q�Y�z�*�{�_t�xə9W:�Ԋ�q ��r*|Њ����v�Ç�oOL��,��ӷ������M"J��O���x�2�]��ş����C=��7�{�gk*�5*� ]�g�ݖ�d�9�^��J2rl�R�ѡ�k�0]�4B��,�������`$w���j��P:�$Z��&�]j��qJ�l�ŕ�o ��
}� �k��@En^:�öv\��=z����J��$��0Cc^�r���uumY��V9H�8�i��Y5$�R��[z����kU��]ĥ���w
6�oǅgj���+u鮋K�{�� �;:C)Ǆ� ���=F�l2��D��2�ٍM僦�Pn��k����c���A�S��9���۔l�G���=�r��i�]Dڗ��i�]��+;U�ݱ�t ���)�V�RY������؇���`�&L�4f���Z"G��Ӎ�Y���w6s�U2T���L,N�p��8�Y]�-��3�.(q>�"�IR�# �iTSV��8W;L��b3
� �Z�LQ����;ޭk�z\��=|�i����)ro4wLʊvp��][�B�X5d��:����y �
݊�XbJ�a,9���4+v�:�H��)%S�<���U��D@�]6�"s(���Ŷ*����c�4q�nl�p&vd.��"9�.���{wV]���ڳt��T�S��:����[�.��۬�#-�����n���m�'�j���
�Sb��s�'K7���ztN-���[!��;ב77:�[�K"g\�6���}c�	���4L����o/���#�S=�L����y��:6�@�*��P�̝uTE��X�<f��ȑ���I �{.S ������R�qa�&��+���P<�5<��\�(oܞ7��nYְk��aG�b&�З��>���"�%ى��Ɔ_K�)=z�*�鉷��֬#�2��w���6R��E�*΢�Y�����xl����-˫�dF���EkzN�y��[ܷ�b����|�xt���yb��7�ko����K�����6�>Ո%��r=�W"����6q�9F�Ij��<�q��|L4.�S	V���M�롧��ڊ����k���J�Zڕ6�k�V�릗T���g�X�6�$u]t�}`��j� 	�>�E��V2�^�7m�9x���[���@X5�^�\a�n��§`��R8��l]��ͻ|�(N�65<�è����v����M61��h� �l���Wr��t*N�輊��	]t�
Gr�p��x������KшmZ��$a��{iت�w3!���&�e�5���b�4��ޤ��/��)bӮ�yXq�e�/(I��|�-B��	�u�J���y/3l��0����A�`�o��v:k�l�2<��\HBT����c��I�A��ϖ�U,��#����Z�l^2�pɐWR�%&Z�2rq���
`Yi\��\��ۉ��M��ۜ�\���ú���K��"��I]+��Z�vut�0\�Cw8a���S+�;�Wu���;w]$]�\mӢ��F�I���nW4snn�ѷ9t����9�n����{/ur]��w']��us���Ӻ�.��/{F˻��+���u��Y�]f�r��F�ws���{��/7�1ܷu�7M�v�r��9��]�ђK˽��m��:n�.I���u���\WSnjs��9ȗw{��7u����{מ9wrt�νw]���wJt�{q^�+�=ttL�yw�����s��<S^����������5�wF���w]t��Oqݝ��r{��D�er%��\��Ǻ���?��߾�ۦ���3ju+��-;a��V)���~D��3�B���,�N[���6֬ϥi#���<�P_���i�]���]]5v��q����}��u`i�Eӥ��^��WefAd�ף�a�O ����q��'��;\[1��E�aY�n�'�(��'�����)�M�%�rM�֛������V3$nȷ̝*���v�]!U+�(:���d;WE3"�F(%��Ѕ�6ӹ���Xq�2���q^�B]��n�@C6�q؍Y��F���Wr>O���݆����Wۯ�)@ꡒ6�g�ʹ7��Fc�/L�7�R_!�]�=�_F�a��T���K�{�	�7Pn���b˥�lxg�qr�ν�ll�=�嚤YK��vW&���1���w�1.�8�c��kU[��/��f�?OV�Y����H��=f�K��;��<�tQ�cl�f�s����e�-�oY��������1ydA��BD��/2<ό���.�C�髆m���\���wl���2N��nf��j[�70��"	5J��6#�D�S����F���z#�5���W�T��:���`��N8�M-�1�|����c`�zdj^�7\�1u�g*cFd��s"�=�nrµ3�>���Z�[�Q�ٹ�q�\������"�xB�y��x���;+R��
5�q*�w`�����m��������oݶ�zZ��	CӾj��-�]Ҷ*����w�����z����xt�jIG|z�TK����+�a���_Hd˫��+^�1[���m��Y�p6�(��4l�*��ΉzL�8�[F���U^��z*���4Ix`H~�u�g]$������U�S�s�]]��ϕv�\Nb3{��W�g@u��HY|�7���H�h:
�H�قNE��]4_1��d5S�!����:o��SA�J��W��3McO�:��ݽ��{1��=,1�K�
��s�4f:�)�̮�[\Q���u<��k{�����/���3K��Ü0Y�oP���1}�r�Qy�L8훽m�}w�U��]�*V���o,(n0pޏ0����;�b��m�mF����6Ͻ7ǳ>x��O͚��<({Ȣ���u���������^�^��}V�
E�[Y���][N��ڙȞ��+�*r��ɸ�P� rÕp�����;`ڥrn��Q�*(�x/��&s䭟�����JG�T���vqɈ1�9c��N�Ȟ�[	:�S׾�W����{���X�R�+����錌S/�=}Yn�j��&\3���ln���)e�z��z7�іZ���q�y	�={Zᴉ���S}B1��/ V�5�H�G\�]uWr��A�.�om>��w��P��V�z�/��oJ��{���n��0�vޞ���}����9� ֮�����7���1�a���6��dH̗�NaxקP_��_Ɯ?Q<�6t~��/H�E�.yz�g��$�'��h۲��y��Ү7Ld���:R�

@WQ��+��%e�U :Y�"��|̄��{A��hY�v�Eyn#���+#JJ�)T����[������u��&��.����nIʄ�Wa|���T.�q)���ʄ�).���E���w<c���;
��Q0�H����M���9SC��[ы뫁����/�e�bR�0m�<!>�^�%T��I���>��鵭R=�����˵)�i��C�I��;{7�*D�w�f1	�Ք��i��0]�Q�����q2k�qN �d�WωY�b�K���
Z���n����ovڽ�$��ϵ<<�N�Y��[�o���"��mm�ޥ�����c�<�EX�kw{k��[`0� ��b�ukcUF��������8�+�.M)��|=GQD�-��������c%��Y�3K�Fuc���8���B6�VqʢQ�������i��y�|
������5��wG�÷�4	�B:T���׏*��.����dKOE4[Um���7�]�4��?PC�!�b3����p�#ߜ��p���L�w�}��T֟g�\-�2��{hgHn��}�E���+�/�/s��|Ӭa��vi�&����صH��}^:(���Їt`E�Yq2�]��+5i��U�=yg7�G���8�����F@ا��-Az&��e���2影Գ^lΊ�4���C���
�:jH���ԕ�>D�U�ח9��%���R�fM�N��4¯v~�;�6��:��z�lR�u�gO�k60z��R~x�6����|'������I\��d1_���V����y��K��\��Ӎ^��6���i��S��h=���[}��v���Mx_���6�k�W�������.0j��?O^���r���J8�;�)�N>�`Twa��)�KPW^�L��^U�W�cdo��������r��v�ۇ����������B�P~�xB���\�fat���m}�w����RfNUϵ[�l�
b*�D�3�m\i���-kK�?rk��.wwv���8�E-�î�N��)2�u��4I���Ӏ�gա)�O ���5�y2\z����GK6q��10�j����h�G��#�z�rl�IET�&���|�t��l�F�]C��-Ź��:[�}r�����������d��E#nv[9k���{Is��̡[�N�?�dB�_o�.���j��F�����U<U�O��_cmL�oa�qރ)L��m0q�#6@!�������o��>7��O]q�����ؘR$O�*벤Lw��s�[���.�k�2���t��R�3f�a\�YȨ�Y��P�"�l݀�{`㕺�8�0�')��~r����u�jw���˓U�m,�)�ԓs]�IݷDZ������Y�qm��gY[H�촺��W��O{�'՜��� ���6��v�p�x��P���6�'�7D�g0���2��Ϭ���Mף�t��>�_2,�*{UJ;���݉��w���)����7���}#Lt�{�i�8���F����b�!�]׷��D�?�(���y�&ٴtf���#N���$Dv�x��b��Y�}������hl[�CXQQk�^&�/�Z�3V*��PL��벓n�]-�Em�����5J�OK?��P�z�l�4$��a@�6F���t�]����	�AGY��w�\ә��?�0e��+���U���UьγѼ]��=���,�Q�fM<���O�i�i�m�K-�7g8�tVq�	l�7�V��; k�����Iq�4׾�8�͈i{����;ݸ�ݪ&,nC3Ѥ+�D���d�֎�_�w�[a�5�ӗ��u'[�P���v02"+qk5c�[%̉��'P�u���D�P����wt��������.w��_]�l�
I�*3��q�5�nf�g���ի5ٹk�e�:s.o����[%��B�]㥰b��\,93!e�v3`��z�,��%������d5S�����GH�2���nR�~Դ��������ms�!�j�����1�	p�Y/�t�#6j{y���ԭ�W��s�s�U��k�wH:]O�0@vdj#���y�-,��ҽusa�����|n���]�(	[��q��lm�pF�?3T������Ī��,�1�0�S���4�ҹ]�+��R�] 􍞦��5�����P�g$��`��L�C�Qp�gq�)e�z��z7XF�|z��������k���ڈ`�g�`<e�F2S��ȭ\x�w�
Ǩ{��٣�]�ݣ%
��uV�/�t�4��e�7�ݾ����$�!�Y�X�>k+���=�'6�qHhD���k���3���zKu����ެ�c�}5|�1�DH�;! �&�yJ|:)�a�P��7�4�֐b>��|-\���*�Y�NOk:�����2e1����C���+���n�̪�r�㣍isq-��:"x�r!��[oG�%K2�Nٱ�W��[Ree���r��B!�X��W�?��{�p��kb�f���6gl;S�+�̾N�U�x�PL��U7�&�E�kܗiB��,� �� ^WH��>m
���G�x�ڕ�sV��1)��B帖C�g�JJ�)T�5D�b�A�&n�o���|94�j�tcyeBB+����9�S�X&�}mݱ�gWKi�s�ڭl��d��v�4��H��t�W"��>��[{Q��{��fS��n��ǎ��=Ǌ��]-t�u��*<譍���l�sX:T�{���q��i��+!R*��*Ս{k�1m�0�A-ܪ��w5+��4�*Q(a�4,��+\��Ew-I�B2���s��5O]:���cp�i���P�kc�����O�g<�wd���Fѕ�*���D|�(p��w�ހ=��}= ]�hKJ&`r/EES@ۭ���n}=�GL����7!�k �F�b-�d_T��oO������n��
���\@��5\ԉ�V�C�o��J�g�\��k˲4M���eezy�R�5�d����]7�vJ{ձ.����lR!&]�zc}܃�.]�����7[���a��XΘ�H]M�r�u�vwhJ�VM{R�hk��ѓ����󾛞��+�{7������Ȱ:Clo3��B0l���_m�̿t}���s���ߨ2�5�Gd��t�tQ�Z��w@���s��)����힍�Ǿ޼l7֢A�D����v
26)�����fg���E�O���^���y�tD_o愭K�]&�y�Z����ݍ|wsbL2�9��HЉ��׼�\�H�H�l+��,iY<c�����X��H�m�i��,z���
�,���!kKL��Ja�v{��:*�pI���ب�䋚s4E���@�e.����pn������>�ъ�2�J&N�_�[��[<�9Y�
.���9����iƢ��� aFCw#@s�J6UүU6��ӭ/3�7"���YZ;�[Y6M�|�D>��tք���t$��q�y<uw�P�yo0t)�k�]��Ö��q���_��w����{�j^�FN�gt�*h=�{��\:�l���[dO9�tz-�"��y�QnL�|a}D���$0�h�ʆ�����I�r�f�\���9�����oa<�k璵Y��������1U�U�ڏsx�ʟh���n9�?�#xt���&��W�*\�hN��W���0�;���i��~=r��t0� ���oO�es��`�Q��ӿ<��L�fzl���Yr��;��>Yr�WH=��8�k�3`0]��ٝO�N^�Nϭ=�/��7xף+��^��g�wz(҅T��[����o@pQ35�E4n�!{_b���4�WR}Y^��NO��:�t{��ɉjb���p\eSr�|@�e��&;7�d(�sԬ�9 'h���1�L$���׊����[�S[�Gh��a�v��Ky��i�7���� o�b�~<r�������#�'���z�k;�(��������#`gu�N�0%�*f��&�����=o���s:��B�=�4"}꺯^#��\F]L��;Q:w�n�XD^h��|��6jܶܛ��f��+�|�����6�>h ���u������w��8��m�������~��M��ߚծ�k2�f�el�ٕ�-S+fkf[e����+fmS+fmfkfUL�̭�V̪��̭���m������̵K5�6�*�V̭�[2�e�f�f��m�[2�eTͶf�3k3U2�f�Y���̵L��U3m��Z�ՙ�3VY����vZ�ՙVe��Y��*̵�Z̫3Ve��Y��5fj̵��,�2�f��ٖ�5fU�k3[2��j���ՙ�3VeY�Y��6��ͧo~m������m�ٿ��n�US6��UU3m���UL���������n�j�Z�L�j�mj�UjekT͵T�ک�j��UW��Z�ej���S6��~UWf�m���f��3m�̵U7��UL��fZ��m�̪�f�m���fm�ٛm�f�m�����U2���m�f���m�eUS-UL�lʩ�lܮ�������fV̶̪�����������elͶf�2�f�el�ٕ�6ٹ��eTͶelͶf�el�lͶeU����ԯ��O��n�[Zf�UիU����������?���'���O��_���?g��?_�����%���������m����w������e�m[j����ʪ�l� }�(�����{�~�����:��+�g��/S�st�-�5󤇽���������k����G�sj֫lյ��j�UJ��j��UTm��5��5������[m�l�U-*��R�m�Ҫ�m�����U*m�٩�U5-��M��4�m�M��6mUI��5o�ҭU��u'[���/����U���6��Z�����-����(" �;�O��  �`��=.z��;��B�$O��!��������t�<_i�  *�4>	�����k��U[m���mm��W�����V�V���k�m��5��m�U*��/�q`�0�C���V������a��\� V<�<~>@ ��JD�f��=C���a��x��`��}�󄍐 ]z�x�� �����0Y=�z��@"���6�z~����
���>V  r����,���`2d?)^=&����PE|�,�������?��y�/������O�b��L��.��7�� � ���fO� �{w�}�*�*�$Q)"������U!�
DT�U@�T�"QT��D*"��D���"H�I�J$��()T��vjRP�"�!�d��AR@�B�RRJ��EUIB�R��H�@�$�IUQ$�(�R�]�JIT�U%�%
EQPJ�� ���B�TR�P�TJ"JT�*��� �CD�H(�BJ (�(M�J$�x  j���v��r\
m�u΢�����[�6�m�i�ʬtn멭�Y�kN�í5ñ]e�Pv�+sU�iT��u�tk\�n�҅t��%JB�Q"��J�  ޱ��ђ�]�t��w^��66��[kl�6{�m�E
��hj�cF�N�L=�ѵ�����������-s�wnҭ���V���[l��p7]���t�`���P[V�;�G\�w%�i[2P��B��"�  p���
s��@�[�[�7F�s��mN�V���mb��Ғ�@N�ٺ�nE;�lt�n��gv�v�j���f�m�CWv��[�����R"�R�	�Qx  Á�=v�V���Ѣ� �wwl�b[�.�un�gq��;���]5ݻ�,�t v�J�������� �J��"%$A 
UQ� '(���,PR�V��T�A�j���R(-JƂAH�i�@,��T�(Q5V�@�P�*P@��R
 gz�3`f& ����
@�T5C6� �[j�M���SY� h���kt .S4k@U�TH*U$	%H(�x �ʪ�Px�ƊQ��cMh(�0���%�4�V�h�U*3 
��@�� ӢjUT!$IH)O  6p��u�� 
]I���çР���  J�� 8��4�Vt �`���  J������
�II�  #� r��S�.6� ��E�  چ:i���X( (Ό  b�t �3  hl��  ��B�E*�N��	
*��  ���J 1�� @K�� ���J  � :��  �n�� �U��l (pwP  �S�)J�1 ��a%%J�� E<���   �~%*(  2 �)�h4 I�Bf�� A��B���	Ȇ/��UĀ��b2z�
��B�t�R�I�U��|��|�f�3T������ն�m�������ݫmZ��Vڵ��M[j�ٵ�m�����~�gB������Q� 0�ܺE�6?���x�h��@ّh�"����]]���Kj
.Sx�7w�(5�w��a3j�&�@nٌw<a��F�e��(%%nQ��G*����+sH�u%�P��-�%[�i�بʛX����3H��.��{r�Q��۽�*��)��Z��S���bgcGt���t���k�I̼8��	[Ϸ��t��Y���;N�8R�k���;�[� ׺Rz�w�]h����h��WV)�3Y����Z/ZZC�g!�� �IEp�f�&�Tw^�ݺ7����j̏aW���umiT��¤̠$����.(�ىV�mcߢm�P�ib��7��nA���BUw(�t]�V����jFrI-X��31A>ģ�V*e`T۵B��%Z1b'qG�c������,��W��Jnt����\y5d@�;��T�b� Q�eKfk�n4�����K^�������{�n*,c���S�`���a��f��*5���F�5��/C{�� �$2�&�� H�_Zd@�1�<�#wY�ea��Ԧeء�-У7e�5�>z��*KFrjM��%�mڷ%�I��Z�sB��� w�%w7$�i]H��B���E�jV�Ӧ�`�43�<���3�ȱ�XM��V]J�M��@�t,����U�MTiP;b��U��N]���N��B�%@b�a�*GY�є�z ۖ�5�����XVK+�ln#Ej��&+R64��ootю����f1�l7Kh�i+!��0��-���⫁xeU��U���,CsH��F(�d�����V\{�T�]���ݷwH���B�PӤ��@Lw���'�e�fB+1��"Z�-��� ��(��fe��N-��^���,7Pf��ZM#{E�M��j�A�HL,��1A[�H���\���J�̠�@�tH݋N��v�?Kc&�� [��`�yRͳ�S7z�*�nB���43�$��V7A+�k�K6�(e��������M��p�A�;��q1%�M�\�j��m�Nc�^͂rKYc+r4�黻l(I�%u����AG7��ޖ�����f��۵��-T�w�k��	R�ut�ԫX�(��x�h�3(��|B��+j
�oon�V��n]DQ��I��r]Q�HF����Wi�Ui\�)�n��(�cn��V0�#5�trj�7.�f1(��́��Mm'Hʂ�Ւ'�fm����z�X&�:��6�v^���}6���\�Ck6}߶��J`���L�a�)eG�U+�5�
���V�^�wI(��O#Y�t�cl�w1��cb��MhZ��2ܕz*�N�i%#eI��F�n`���	ͦ�,�V�э�4ýod=�`ZɈ��a���7w�hG�3B�WG�?dk2�ݧ���d��f,r�;qm�4T�7�i��E�$2ęW�γ��SL�c�4�K RƋE�j��n�:D��"�|��3�ŻG"455u1Ĕ������R;yS�Z�An�"�6��M@� �h�i�ښ�	tV�-����)b
MnZP�:���u{@�
Msk��]*Km�//5zXx�n�{*ܤ�^������M����$��,3Ed�Y���]!�-K ]
7�93.�ɶ,U��	UF+�f��ٜP����+��X x��TX/5L����%d�B���F�?AX�n�@�t�����1]�dH�Қ%hI1EٙD3rf ���j�R*7�X��B`�������"F�N��n�*����X^˺ҫ^��ax�f#x��db9��5�WKh��͌����:9ݶ�zm9CD���4#mG����Q���4�bW���R��@Y�%x�2[u+��;7o
Q$K��h�{z�:�)7+ ��	���J���f��3&�U�NZ�F*Vj�J[�j�Nk7�T&jrT��I7��O�3�ѧ�H^��Xv�ƬMq�8�:ܗYF�f��&�����vJ�H�Q�Y��P�U���j��CiZg2�L���$(O\9��Ҭ��8��@{�E�m�"5weس���Ҏ�����m1��VؼND/T+kQ�̆	���Z?m��P�aiYq�r��6F=7x0E@�̛��v�K,Kƀ�PL����ۡ����b�ګ%�N�ѯkYм�D�5�����u�jE��كH��ͫ j+���I6�Sfڴ���oa��Ln�!�j� ���Q�ޅt�rMY�.�;���!GE[�4�)4�T]�0)n�i8�%���4���;�w#V�@n0&��,�\@���X8��^`K�t�O�B���e)��yo
A:��n�r&�WxV�#C �n�u���he(q}���vhkVk2��v2�� R���6�;F�D[��Po�EַQ��"�[�v�ݼ��2&�*!fB&u��� ��k�"�ҽ�czM*�	�a����-:�N�����a��+u|�
�6�m�u^&��G얕/��3Ŗ.����Ԧ0�;�`�%Wl�l��(���B�,���\@d�V����J&��!�9������ze���7c�f��'�t*1Aa��InX��ڹg�� f���h�3	��ͤ�[Kvح-�t�U�.�<�V5+m���n̄]�tQ�N�+��e����Y�m�+[�e���/��@Epح�fd��ѣ1�N����J'a�� nٿ���t^��3DX�(<dŰl)^�M	c*�϶��K6�l0b�3a���Am@��h<��r�L*��fP[ܻF��T5Bm���{�`�c���nɚ��X�nK� Yi$6KXl�V�an�,F�͘.��M%�������* 7nBq#3h���Ư xv��r��ձj �z�;�ҏ�)�M吪ݻk��y�H�U���p��V����K ����0����y�i&Zەu����в��DbR �����lX1eKq��F0[k/ �w%���'j��׃S�;�B��8��0:sR�(P�����d1:.�nM��NB�~��6�mK���8 �$�*�`��5�!́���T�V	D�B�+K�N	��L鐙[��m�Ljͻc���j
�κy�=C�@�$��Fd`�^�e;�y[�����i�ɰ[؎Ӹ�M�Z_զ.�B�z�
ܳz(] 
�V�;F�7�+���)��h��;A�L<��ƶl�n6��>K�%n�D͛ġ��ӱ��ʷ��2,wz�
M?�㡫.�i\tFm�5s[�y����;��7#�V:6�S�*�u�L��0A����r)���ii���d�l`	l��5-j.
l�m)	�&^���!)��F.|K����Hq1^Z�Nkf��1pѷ�.K2ۭ�wa�妁2@_cv6�A������l�b�4�fB���Z1�G[�	z6��6����TԎ�r �i���ŕ��q=�j�H����V��;�3y�)
a�J=�P�h���u�M�x�Ɋh�R�^�/�<YH]س-�USq�!yy�-9��c��5���pܓa6v�\B�KWX��[�E��)�Lt�,�L`�w�Q�a!�z쁴*�5�����n����C�I��%� �ѩE�Wp�D�;�*)���"P�r�䡇C`R�x�+AѨ[e�'י�+$���fI���gFk�i�z�n9{
ǖ(�8�T�^�7��n<�|���.S�n�c-�s�����S0�I���V5?�`g�p4�6�&�����X�a�#h���@fn�C��6�f��]��Xd��SL� X25{�F+I���U�����N�Z�~��-cQ5��c���.;o&�F0cxae@���Um��]�-���Z't�����n����R4DQe�&Q�OVhm�J�ȕ5e�ڗ��5��K4�+q�l�e;�@�$�w��S�%R�>;y �A�B�$ZM;!���l�����ܺ�C#4Lv��sa۠�m�� 3j@��0���'f,-�*���Q��Ό�&�JT��R(䫷4T�����Y���-�Q���R[u �n^����e"bS�l��'c-����J�3+Z�s�1�[�!Ϛ�N��J��j�3�=�V��˸�^���D��,*�YV��KYBd�r\҃���	�&^!w��D��X1D�<��,�yZv�fZ���(oB'1�A����
b�z�.��Q��)4�{X��i��ݩ�v��j�'S�ol��
�r���N6l��U����a�	} y�X�0������7$İ�3$��b�Gh�ӂ�m�E^:8傯4��X*�#ֱ9M�F����gn�
�n�nT̩�̺1����jUC�V��� 0&P����u�V��õci���#hiMa�K����Ծ�yV�S��J�ڠK�+i������Wv��� 5�p͙2-T�li_%tv�
��a�u�5����`o-��A�B�i�uf�����Xp�.�3�R���ٺ,	���&5)ōC� p���H��u3F�z�-�T�^���ɰ��{�5��9��SUl��r�z\�74l
Ԭ�� ڰ��m�ʰdwW��ڎ���%�a�Z~��%)M�w��)����[Wb�d��[u���f���#�Ӱ�Q�F��@�����\��1;�����y�������Ф�F�ݍ^劋7]1�5tun�ǔ�yQ��=���3Uİi�3YL�B��܃&a� Ш�E��[LF�B�+D�	������ۋ*�cB�i'
yJ�%�	R]���wk&�MM���!�eR����e8�@d�Zi3�Q��B`x#Kpo٥Y��	d�;A�rM����S�3����Wv����۩YWn*�V6VTӓT�33 �a:���Ê�p��{-���s�� �R ��@e�56����L��n\�75K*�\H�B�]$)�oL"R�K(��í��i̻J�暗k��#����t)��*�Y�m�2�:i�P�Z5�ֹ4�d�	{����*ǖ)�`��F� �)/X�0�����;�+Mз��1��T��T1��Xtwm 	Vp��	��j���-={Y2;��ig(�e(�Yp)���8�8S0U�`���@a_B.��2+6��i�|ȃY��s
�Y�S���':� ��{�5fӒK�����jle	�
Z�a{N����fcݲ)���1
w����U�p�M� +*ٴ��b�K��R'P.,��N�O
z�ⱒ�R�9R�ϩ��@+u7Ai��^5�è��A��(�U]"�RV�[�3Ptm�	�?��ԨyA��i��Dl�Y��6'��U늝5[��4jj�3.�a1����4�T+a��%v�T������vm��q�2��.ER�v薘و�Bi�O�{�������4Ӷ`
�Ee2f�Ӧ"Љ{wePWR�U�\�^�R��/Z�G"9I�U�ϋL��X��z�=ۢpc��V��J�7�]'8�WB��rBr��G�i��H0Ѥn3 rMn�������F�v�iko~Ln�0��V!a�����h��!X��a�
͘hCv�`�ţ��wW�
�m�
�1V�,�5o\��X̺=�	U��]e$r�gCm,ҹ�Z��.��x�4�mm�1��ܩ�Wj�M�3 ��B�L�'[�YE�Y��1K-��6U��C�����6�#L1���_6��L�f�r�����D.�j���ۉ-k!J�ԣ���Tx���io&��a׻W���;�pe��z�˙�E��;�2^)C����m��1�՚��oOh��,^�Ԯ욵m�q�
�36Y�;Kx�K`�74^=S����hlN��X�FN��B��{P��2c�kn�y���7o��Vԡ��1�"��*CR�TC2D�%j#I�+e�֪c�E��ޭ�e�bUn}V�ʩqb8�÷�m�S!{*@���k�d]e,X�v�敩|!�B�EH��j�7LY���ne*Y�ϵ�cV^�R����0��hDV'��x�ni��
�5� ���N�{h��t#���P�h3b�c(�f۲�FS�U�x�0Z�5��Ek�[��
�i�Ch]ae��Z,K��PQX�kj'�$��6&ʖ6ޝiX&���1ƔHj5 ז�`�Ć������1`9&��էzF��O�bY6�;�e,�P����Z���>����&��Q�n����:X���}#1�vc��72A��ui�J��x�Ksn҄��(�el��P`W�XKQ)iTVFnX�F��6�x��ӕ��r��
Iȍ{��1����HՌݰꦂ��kݚ�o"��*b���Cw���*S�mK��JЎPy�X�9�օ�I��6����)Hը��(#b�^Vn��/	�R͉Ԑ\�����[�5i�L� �i�n�^B��Y�������'(��SE(h�KH!�Zf�U{����I�&*a��ƀ�Y�{�ܨ��S��A0�x�oVR��8�$ܴM��*aӸBGkd&v���2���MɤZ�-��P���Zk`��J�J��/d��/rӘ$ܩK9 �*���R
)ռ�n��4���L�)S��p��Y�J��{��>�4bcrQ5�5������7KB{yt�J�Pc5��R��z� i]8	5�� ���Ҙ�b�2I�ZZ][Nj3�z���wS�e7����yx��!�O7X�h�EEv҃5�f�*�U+p[�z����R� ��L��lyV@m
�Ҧ(P�
�wD��:9Km��$2�)��o�f���q�6�A%c�oC^yۼD���wg���ë2�Ws",��D�mGX��6�����|+�� VǸ����&�w���e�5N��Gm��Ux"�P�!}K(C򮽬G��B�ck:��s����7�	�x��9���}���bc��Yvw��K�����@^o���60w��9n�e��Tx��ǒ�{3���-�txѠ�S�`��0k��,Ȧ+�ώ�Lt�V���]X���a>xY�֪"�ٻ.�k����!�q�ҝ��[ ��8���b��\&�e���0�^��sm<*Zz��*e��*7"99X˭��QƠm�e1�Ǯ�bd����kr������tԇ':���Y���+��,�p@2�+r���3���ͮU�[�+��`c��8ַIb6�y���];�X��2*7������m�$��e�˵��}�[��S�Ƚ����j�%=���7I�L�S!�,�L����t��[��0e�{�X��v��R�j'�]OU���.V���(�Z�h��wYIs;�!�:� Gi����.Pݳ�J��)�ێ��2���wh .Wq$<��[ٛԲ-������`��gy/�7]IU�X���㶊�)���ɠK�+p]���WS5��j�m*�]P�a�=q��r|�L��!�n�Cm�uv�g3z�jԠ$;�򞺙�wx�l���}��A�ݐ�3�5�*��6�0{کI7rW^���f�g**��}��mqI�R|��ǟI��JL�]�}R��J�P������6�\�#Q������P�zJ/hݶ,����Lwf��(�ȭ�$�+x�W0�=<�5˳VnĠ�\��,��an��ϒe� -W]�L��[�+�����!��w9�Nd�-�l�� ɰ�xNp}��������o��b՛hf�'e�]�M��긵쾠�X���Q_P�p+L;�C�->s�."IÆQ⠫�',%6ͽ'*m�iJ֒/-���.�\խ�8U���ϰ�7��;;h
p���ppj�g3�k��oJ>Y���Ԅ��7�w����O6'�N���ެ:�efe�[N�dWj���澦�Z(܉=�f����ܮ���]�	���=��R�_!Y`��W�]>P[|���u�ǻy��)[� ��.�R��
ӊ��]Co��z?�S�s-�����8i�t�Ǵ3w��b��'���R�d��n���t�j�U2 �qrP�$L�К��Nw��ش��28��a�k9�W�e�bu��ܽ�ݐަ�<L���r��]�j�Z�j�����v�VV;K�3���ZQ;�[d��z�n�2�N������]k�vN�K���d��ya'*O
�aǊҀ��t%e�n�[�_GA�TN����"�j[�Q����6ˀ授􆹼y$��\�?��Y��^�g�}(�:�Nsz�|p�=m 5���;'l�g%>����ʴ��pob9Y�XcI�㦎�`�>Q��1�^�MWa먚�H�5a!�(���nU���b�`	B�՞T��|t�����N\�9����XG��ɫ67+Z׽He�j?;or����m��i<9�����d4�Ʈ�`wrExo��b;c5�(Һ5nMjЄM{�*X(b=y�X�ꒃ����%�p_^��]1{ъm�ܬ�D�v����&��0Ǹ>Ppq55CBu-X���s ���Q�+��ׁ̣�B��!�35l�U�h�Jx��yh�aq�j��ڃ�5���뻹+��mg0c=���w�eK]���iV�Y�R$l��ƵR��2��CǷl\ف�e'�g"��NY4Ҏpz趞�}]xm��e��8�WjJYF���k������KoSn�sv�\��K ����#�*��`[��.Q��v�yD��S�%>��%�!G}�}�QK��.�q�����R����cW>yA�ƟJ�2���x���m�c�=��>F^�Huᨸ��ݺ�6��Ys7������Aj�-��V��.̼5��R �[�T��d���w��;6�̺�w($W�%�
�m�f�2�J�2HS0.&��]
ɵc'�R���[w��8#M�ܶ�'u`�t|�˧����l�5h����;5wq�r�DǇ+*�)�GQ�\�	�q�wF��w6N��ι�b���}���=��v�yt�9��T���]�G��1G�I�,�}������:���]b�f`�I�G4T7W+���i)�b�}�*�P�ݩ[��%��bʷ|�C������rqv�'>��]���.d=���9�k����S��X\`Z����-���ԛ�n(�;=�uϟ3(v]Th�WWX%�F(Y-&��=[�).� [V�C��`��0���Y�	�*��
����ƪo����ҩ�+�f�qk=W��BN�Ԅe��e����W��W���;HRYQ	�v�%kN:[���᳕�B`Mn����V[�s�l�n�]��ɚ�1ԋ�4�Q�ojXU��H��
p��1'�5���M�ƈ�Sg1s�����L���	��yW}�
N�E�o�3�T�O�y��<R�W,WI��SFq&8Q��d8�|cz�H���`F�}�fu�z�HƮ�8��F�O&:�h$;ǫkr�l���Pv�����XY���)ܫz١�5�_`��>���'�<oێ�?w{��I+c��s�G�VYƅͧ\:� �[`u���t�v�I��Y(��Y�z6�u�+�R�/;��{�/iE�6崒���k��cr��9\l���KW���mu��1u�yWz�N�;�`+�.`��`rr"������5��}W�WMc:�J��b�[��Dp���c�EfkH�pT2�a����-�F����K�<�tuhV�7�����n����p,��t1\v�JWR����Z�7�3 �hKao0�U۩�,�,���H�k�sF'Ө3[x���[�U�e���ڥ�s�1u�;��ʺ�ݝ#^f���*�r�pN�+x�F�>ʣ��Q:��Gf�vf�94�-�(*��]
雼
��2;�peu�MYz�WSPPZs]�[܇����kM���R�G6[�HM����ٚढ़���2�
��t�ثY���+gR�71�sU�ە����s��,��rV��շ!嗇�A�W8�K3�Pkq�a��u@�70`�pv�e�(	nb-�݆r�[ZS�,g�l�vJ�}�o/�sfS�v���P������C�mByqŊ��헽�A����0d��1'�r����s#N����v3��`wRG
��U���W��OQ���gc<���k���8���N�iz��~���K�Z׼.%�Np${��loZ9xhk�LJ*�\�LX��&�К+w�:�E��y����T(@^$Q�W�X�y������9�o��#��)s0
<����up�T4b���O,��	Ҙ��a����o&��Q�g�]��s�Jc�M8�;�I�N쳫��
.kwi���t�<�wVR{�� �>V��xl�̭9�k��Y�z�eڈ���O'2��u�w��V�	g "�t;���;]�b{��O��Dݽ5�g�k3p��&Y�����묆��4�Ĺ*�J�I�(+��sV���Y�:�<tuA2�el��@O&ei��l��r��zhnm	p�P��m��O|(t$��h�	��;:-�.��b��J�hܫ�R��y�ޭh�<sRu�O�_:�T�O@� �Ҝs���YWC�NC�wY7�Z�V�omҭ�g&{d]�n���#|��{�]���ڳ%�F�x�ɲ����^��V��*!����z��9Hmh"���lE��o-e_u¤���ɳX��S���zzY��"S�C�E�D��j	Ѕ5pw�[��G��a��L!8���Eذ��%�ȫ���M�vh��æt� �C+���l����I	���c����|� �v�1oi��e"ܺSF¢9*g�Ļ����A��z�Z���q�0f�Qˉ"�32�PT�]"�9��=q+O���	�GԢ�h���=!�{�ŴƪƯBK���G>/��(��vZ��I�q^$9�`m���,��y9���ƹ[�hV�#�~��u{��-s�Q[���ݢ�w�;�|M6�#�!w]� V̧�!=|�s(wph�锳��\��]��y�Q�"�f�O�N7���b}�����=��MK+4���m]c����=Ҷ�����ƫ�`��мmr�ȺU�����;8o8�e����̼��
��Ms���� O��:�����%EB�vạ��M��f�����ۡZo���N����|�ɏre����Ѥ#�u� ��2��Ĭ���T�VT���s2�yI�Q��J�`=���*�h���v��;.�H���B��ޖN	����� :��F�v��.�Y"�5��G��h�ܛǸ����,�Tuxb��#���5�a�cz��U�kz��p��L�rp4ӄE��/��*ݽ�u����=ZL���DƸ��R�޺��}M�0m;��U��{��h�LWr1�{P��ᔣ�E���f&Kk<��ޫ�i��[aZ�;H�Ax�c{�X�4��H��y�9�S ��j���˭0 eh=ص�hq���[N[_X:(�����`��m⇹ﺤ��,�TX�Y�5���O���s_M��Pg#��v���M�*Ռ��V��a��R/:�N��9���7��]���-���d���u�vԥ�ܵ�j;�7Y:P:���Ձ���d�����Ct��ϵ^K�<�K���c:D6�yJ.^؉�����!vǉ��&,[YkbP��۠�Ӯ��}7QGcY�}t��N���� +I=�{j��gR�<�r�v�eIr���޺�s1�V�;��%�eu!P�����{$�3�J���7v��=�9��6�9&�:
]k�AX�7=̀6�4�x�iIګ���w�2���O�{�o|����)˨e^r�Gq�\�Q�ł���Nw	a��e+�"s5
[D��+M�oL��f�㾈X��9�m�d�u�{9������u"`,jx�*k����}�A�c��t5��U��κ(u^�N9 O�%�tw��5GC���
m)�E'sv�c��qS2��a��k���ke�4W
�N�J�]kz>��j��4�`�r
7�^�Έ�,elû�@t�}�̼����4�I�5cK�����٘�.��ӹ*�S2WU�n�vm���V���l\���$�
�m���*mB���Y1V��b��N�f��>O����K�&=�۾��Z^.�',��Z3�G��Ⱦ˼�a[����
�s�K�B�L�^O��Iha侵x0�;D�ɋ�ouʗh2�p�v�e���R��Ɔ0�w+�!�8	G�E��U��E����i�W�[5�e�\�,�t�}i-]�sb�hQ���إ�q�|���m뮴7���7�Ž!��c�7�_C��2,�xg!�iV��x�h��.��a���R�7M9�s&�՞�M�\�Ե�/+��������2FU�R�^s�x&�r�E=|�ܽ((Lno]7M�4Iv*\�X�!�:+���E�FR�oe[�V�Fkl�&�7a|-���"V���|���ۆ֗)��@L%D�Ę�$�5���%�	������8Pu#������t��h�J%B[ޭȵ��!l���|�1Y(R������܁�g�[8�3��
�C�G�������fy�+d�4��w,�ը�I
��*5�Wc��]id�Z���;*5L�]-�pe�6�m��(:�;�s�O��.�s[��	I	3�P���-M�^ �H���ZY�^Y)��eu����C+��:6��2�K�ҥ�K)��ɹt�j.sky"��_<n��!Tn�Ιi9khX�onve�e=����B�'z�P��I���BŝK��q�s-;�]%��+�c5���]W�;��#Ѽ�ǵ� �0J�t�_Ʀ�K�ۍ� ��Z���]����%��W�*2�nK�1b5%^hZ��[Y�u�;���v�����m�\��7'sgՎ�y�UdN8;"�$v���.��z�\Xfԭ$���٥�O&^�<����t*�I�Ruc1�;��L`��.{ln��3�f�y�n��q��d�S;/Sw�U�Fn�pm�4�E�,
o����}P�n�_gE׶w���;X;�k���HXN���~�O�3�t���u����J4����:{�yʕ"��mn.��°v��쩧�]،E�w���V���
�k��dl�7��]y���� �uPC�P���c���]�/&4p��TI��z�`�uݺ�nJ5�D.���nlҠ�w�n>U��Õ)���;+���qU�*�ʿ_��V�]ŧGVZC���"�@1Z��n�|螝��㘝�����a�R��@��\b��r�jo4�n�V�[�ܴ���ش�Ȓ���vaqZ��h����5����M�����֬�u�w�὏��j�8ĺ�q[�Y;��Զ��C�W�v�+���k��Wft#��AO���(�k�#
�>(%Γ&S.n��������B�W���LL�#���Z:�T�`����ڊ�^��ʜ�;��z�R'p���㽺�3RggN��FYͼ�z�+��ڐJ�{�Xn(r�c�6�Ԁ� ���������P��6��a��w2_s�m�b�����f�J��J��Q��ݬ�l�]{��:��S��t\��@�u "�.�w>�zP��զ��Wf�h�-^173d��w�w�]�͹B��>��D�Y"k�o�A��i@r/�1��8���;�o�w��>��e�B�L��v�0��w*��Qmْ޵+�أ;�M9���P&㢶��,�}�i2�eAa��"���\����iӥ��@b�b�͜�1&n�l��f`�>L3 ���ff��D=AT��8|؁���e��A�9ֹ�ό���>$���`��#1S2���L��M�+���.W#8�œ�� ���i�[�XQ{7��s��JZc6Nh��m��]��q�MGj>�i�`u��y��p%�h�ܫ���>S��g����WS���7�&R&j��M.��XHk;��ٝ��֥/2��V�E;\�y/��u0�p���(ɼR��vkw*�ú���j�Y;�m�jT��ֵID5��/��Ĝ���f�l��\�<�HT�)Ih�P:&h����Ƶ�[����ۆ�ٳF�r�t��0���4mo@�(��zº���!7Vti�(X0R�6"�R�pz���pb��u�*<U�Wz��=���Ѐ�W5=�4l�HU���i�]ݔd#r�7(�u�Ɇ��b�36���X�b8dTE<�n\�q��R ��o3w29 ��U%]�����S����Z�Ӫf
k2iQ�f�b^ں6���U�ojLAi���MtO���3 �L7��4s��rP�p���``B/pd$�Ë����>��k{I�*�7�w�|V�ee,ȩ^���Z���q�G�`X���ʓ"�˅j���Wv.�/����˱�y�i��9Ҿ�'
cN^��ҡ3�	�!�٦�.V���S\y#�\HLww2��p5�+0R�Go����VZ���lܮ������ I���H����w]����N�Cbu�:_.ٍۖ�]�K.�x�'����c����i\�o29�_D�4�<)HV+����*N�6e�՗8arX��>vAș��ͫ
	1J�5�w(v9�ƾ��+)�b��;��s�V���嘻(�O���̾fbj�{dۻ��GS`�=�P}��O�n��=w��a�m}�@�,'$��2R���Ug/��>�li�[�ҲJ���(��㹶�[��z�v�v�[�o6����A� ��JQ���u֭aRHU�=�Wʍm�<ũ�J��L�<k\Y��T�/������4�% ,q����&d�ky��Bv��:��
�8
�E���I�����ҏ���$�{�+.��w����;@��>u��'au�/,ѝ@��ݠ4�&�խ�4���ù��^ŋNK�g%+{.�'27HP,L���S���;7x�m=ھ�<-�ջ�	�75�O�w]w1[����M��M!Y��nL��ɧN)�l:/�jJ*����=� ԭ�>5���5�
��/6�h�M!��eh|�ț/���e�m�p&�8T�ӡ������'E-��S7a|tH��R0`�C���Yu��>��3��v��{^��2^"�kZ��n����5͔��fv��Ov����G)U���,���t32���d�k�b���Evqލ����U�v��ux֡�d�216�d�6O.V�.1uz6���|�,!j�X�u�;kr�I�4�׵ƕYcrv΢w+;��f��K2�W������p:1i�k�}o��֋�L���Y�M�H�y�DX��0t)��2	ً6KL�j��fZ�]b�����ӥbcEk�n-���ɉ��]J�ֻY�h��*_-U�e����u��3NN})D�t0��vd�d�V.��c��u���ʉ[O�b��Z@Ǫ�t��&�1E� �(Von��*�	�i�[ˊ��Re(��	ĚY5#6�1XԠ��0NϤCn.�G#}�3���ul���I�(�6��0Wn],��ZV��v�VS���T��^����nU�	tӻW�y��@(����*�NQ���q����0�f��\��'Ko�Zbҫf�u˚�s�v�%�o 
����k�2¸�H^ AeX5��>�-�����3-!e<�SU/�F�=��Ӭ�0��D�L	�8MeX���ɰR�u����hl����\�\�ۇ,�f���S]�Ud5�M�p���S��+���Q�n�=�v���tYB�YW���֕',�*�ֵ�^k8��-�T�yo�J����3Ie ���Ԕ�2� A9�b�G$����{�X�����v�Ӣ$�dV�!�F��<w-.��&l+�L�*np�*�0.�����6��!:�ܧGb�[áx���6o`Z�b'����#k.��5
Hk��� �d�Wgt��
b:�n�yC��\�1in�TP�F�v�_'͒�-���H�޹����ۥF
�>\�I������Rǖ��ؤWT��O�, o� ����#9���X����.ur�)�fAY0.��Aī��4W��͊)Ύ���Ҥw2��1��z��.���WAFm	�|́��nl�j�fN��#o��n���m82Nh�u8\Vw�C&꠱L���D�xi!�xf���t� �6���a@��קN���V����m��{Z%(�w�4�n�8)`p\ݽ��[(K�X�N��[6j�3w�u�)�L\,Td�l�J�a�fPڽx��w7�����a>g�O���#r����뀋��=�o��Jf%��4��.1D�P���pe\��"��
�!�p֖A|���ӗh�j.��ahWf��\�̳ʮh��f��[E��ۡ��v��K��4����+2�P�l�� �uj���K�f��=X"�+�)�+)t7�Y�8K�b��%�e�ފ���hՙ�V<k�%A�w��"���b8I锢�^#V_>d�s&�/���7�pY�`�v���Z�������6�
�Z��N�]��qs��ŷaʇb�9���׽�^��ꏇrǵ��"z=ԡ�kl��P�T�ɘo������~ɔ��@m�/��� ^��7U�r����G����-֮�q�p��&�n�Ar�ʾ����eI������P�����&�����3q
m�{�Y�����I�6(>Q�!�l.5�7Koi#�1m��څBۂ�U�1��(��c��R�2��ww(�'s����)5ge	�͌���&>�̍�=���,Q�0m�~Ѡ|�ud�d�n��-Hp9��dŋ��7�N��8��{��U$��f졲�Ǽ{p,��UW]�z��=�O�:��>�z�iZ��&�ӆ3:�j@�7���V��Uܾe��~&L�d��վw��/���R6�N�V��ܺΈ�t4����&KT{Ŝ)���M�!�X�)�f9ՄM��R	X)g[�5֙�/T�y�!�ұ���Q��9\F�p�;3Ͷv��\1�c`Hܷ�t��|�f<�x�w1�d�Ƈ:��x�S:��Lb�mY�
��n��F��חFo\؉{��9�"���]>��dpa{����,�dI��=�Uݚ�m)������wik��Ĳ�K�<X�wX�2oy��]�W��[]\2���"�k{ו��ӄȄc4�S���o+v���c��\��J�p��9��$���a��b�]�a��AqU� �p!�}fr=�Ee��b��;���wwl����IlҾ�c��C*��cx\�&����xj��J��6ct$v�A\@�Xv�G@��k��wu���,��*u��e����2��R�i�Ã:��98�7�t��Fe������Z�
�a�����R�%�#�"ˬ�NjW|�4q��Sj������G�w���{�̠�Y Y���	� Z;��͙��-��#���o�
OyF�S��������63�WƊbst4�I=�+��v��o�hPT��Β;n��Y8��:�Q��
Y��K+��3���)�ڨ���g�;2���	Nd��:�yWJMh�d�A��'Uw�O}jTa�۝��ˬ���j�VR`D�L�)�;I������,�K���҅�Mu�ǖm�*_Q۫�ޙ;�̨�p+i2�3��W%e��+|�i���ƈ�G�آǪrU��t/8�+���7]�s/ÆN]�<0�ౄ퀘H�{�����:2��+��ٮ{.@�[��?�^��O`�ˇ#Q���u�:[N�%ö�<2�,�
�|�\�D�Ҋ����/�z�g3�ȝ����W�x�V�r��xMҳ�T�O;Z�0�2w[ucaL(7�΀��-���kEL�j�s�}Z�{�]�������q�d�/&u��uݖ�"�^h�1V^_�˺a�f�v�{���`� *ͥ�\B�oy,��`6�8�X ���LaH��Ho/�[�׷2���K;����]�h�P�	]�;��ֺ�j�%+�,��c ���F��L��G�[�v;r�R	o�Ѯ]�^�µMk3���t:�L���G�f5BKr�ஒ�jQ�X�H�3mh8r�uH��Mƛ��5���M��P:�ۭGu��i�1��%a&�N�#o!Z����K�Ol���n��:	Q�u���=U��V����z�{�`l]j�SY��J��n9�P:XmDM�1R�Ú�����TnVָ�Ȳ�nM�B��4�� yD3a�}V {Z��;n�Tt�U��j�77(4����Z�01�3s*ͣr9M�����A�̴�0�i6�ں��E'n����R�\U�'DbOpg�!��e��f�N�YVc�u�F2��L�^�}Nu�sqw�*u+�ǔ�P��(��p�O/.�T��� �/3�t�����2��r�hAAN�2��]��dJp-�̲̎ݠ/n����X��X��'[�GemT{��4,e/��]Ėi����
T^�X̬���5o1�(��q���H6�.�v�nʬ���ZDssU��9Ľ04�L�[�:%�����7���ե���Kb2YT�-V�ѧׅX�{z���>��&/�\�R�t	�s���e�4h�un��P�����G���m*1
��֮�2�@��o39�@��N�;�L�(��4�T��=O�y҂�s;��r����
kW�O/`-YZL�-�)�ی��1h"��
���f��#��U�U�K�Ւ䜍�o��6�bެ���ͣé�RL㳪'O�+{~P|�mh�a��'V;�eN�U4d�6u�oz�š�^VIt2�=�P��|�\�Г��
�K�v��jw�f��i`n���%�+�Z�X�c�"-���Ur��d�2/�f�^F��T��t�]4�]&^%B��YƬe�V�Ċ�2�'�r4�֢�ua��,�݌i���|��K���8H��mEFA�=��7��H��W5Xe��bvE���xdn�	��F���F�Ob�cF:J`2��YS��l��[�	���)k����J|�v�U��ec��8�{��r=�]yu�2�ò�[�����Xup�$۫ǌ1�k`���-�m�I����B�#�z{ ��QYhb�bƍ}�C7o~{�D�m;���� -:�1�班�R�۪�Q����Ux���0ob)'Gc\oF�%u
�<hv4/I�;�\޸q�"�ԯ�S�\*;y���՚nWB�,�t����/MA�N�\� >�l�;2�
ܻuՋnܣ�M�*A9Nޝ�F�F��8&�^V%�S���X�{;��\�b�Œ	�����IU���뿂�u${s��#����r7���Z��]�	�Kjj��k1m��Z�iŻ�;�$��/r���WPa����A����nM�S�6��
���ޢ�N��4Y���}]����eK�Q��I��ۦ×ƃ���V0��mn17��R}ti>���W;�\q"��w�2r����o�������FvEwݖ���f��ܷzAL�go]h!v�aV�ky��%�p�n���X�L��S/;RY$D}�V��f���Zks����(�bk��]c�eu@�up�v�Iݽo�4�h���a]J�^X��R�f������8j-�M���n��*U�]�i�3�[&^�*`W��?,]J��`0Q6>�8p��T�&����e�g7�>ϝs1uf�����͠�ޘ���3��]tȮ<<��
���oBӒ��-^����z҉^v���� 4�&w�d>��ë�R�rL8��/�v���uU�zv��d쇶�q�YB�����`!�q�3�'���§S��nk��wZj$e�X���݋�J��Y7+3�	8q�T��7�A;i-�sK�� UgU���u������M�,i:l�
'���ӲGنI�ͬ0�J��v
]��yا[2�ZΈd�)�fY0+вo=�dTyB3�E����3U&ɘe��n�wtZ�
��[e�Y "�8S�i��T��w�G�n��~Ϻ5��K���I�wl����II1ܹ��v,}��ꑜc$���ѩ�(ˮ����8�E��S�md��j�Ƭn�v��K:��խlwOMt�L�`'\��0���+WN]V^Cޫޥ���60^�x��'-\U��-�e�I)�`���0*������6�eɸӊ<y�X�6���\�y��h��m��!ƨKcqWZ]C�mu읚݃vĽ�hj���m�X��p*�����BR1v���(�*�|
�����ؗJ*��eں<sy�t�[vΆ�w} �rV�X�YN��q��L(S4/r�F��VPK�����e�0*�H�wV��ح��b�4��PrZ�Z��c��:�9˶�ur����8��7n�^JZ���m��V�Q�&VGi�:z.��n�M�t\���	b��l���T&��2�(���J�sך���Ʉ��@n���>���k�WV��q�xz�x��O�/��B�|�����g ��Lu.�r�/Dޙܴĉf��	���o�ǥJ�^�T���Y�t2Q��g9ϭ���ݰq�lө�A��9��j�@ʐ&��L����}{)-�OS|�g>aC�|��Ni[���R���*�'Eӻ��W��^.�e+}Je����}�3 ���4�e��=Ƿg����>�Ӳ�`�A��#v��K5lIk���t�,������`}��u�����M��sI]�N�y��Hu�ꕓywL'�lW[<�>�}��a{]Z����r	��	�a���ڰ2�V�[+���L�Ȼ�!/I����lr�_��Җ�?3��%OW��ՙ���:h
�mnH)Z�5t8�õ!�I�.�2n�]ә�v]a�8*�4V�{L�	�`P,\��o���6*52�������J��Yc_6v�soR������g��N���TeJ��7���\K�q��D3aٍ఩����չ����R�P��os[4�J�ʇ����%R��jұ!��,4����B��<�3A�.���_]�i��Rt㙋�b�i�FfV�]�=�9H�9�/�xMM�E7z��`]��g-�vF;9	���u��	���͸i1�y�;��yٱU��FGX֌7$k���H
�� �О��XMԠoM�CMNs5
Q�mS��sug;.�;��\'h����S��r�3� ��j��glK� 3�q�hf��h7�(�����\��slݱ���S%9���a�ԷxcGm�蒤�\��Uܕ{��f�/�5�M�W[IJG����֎;������} G�k�[`᳦�k�w��"�D�f��-�Ϙ�=B� [� &�վ��o�����G�N�]����3$lX��S,�6$���A�P�c$j�%3c�le-&Ia�cRb�blQ�i���RX�!c����,&��PP���ԛD�fƣ�"0b��6�TAh�cAiJ�(,%�bCcA`�h�(�6#b"
 1F3)cd5(Ƃ�fQ�����UL1�&�h%#T4�� (�m��J1bjR�E�2�Pi
))1cRI�cE�,�Ԕ� �E%�A�#" $�X�1d$4�JƢ1B1�Q�-�$��P�B�
�(�U�	f���GO:�\cJ���^vd�Ŝ&gSNV��������� ��r��C4e�M:B�I��/F�7N��Y5wX��`">`j��v��%e�Rr4�ؚ��@�Yq%�"� !΃F���ؔ�F�� hr���?(��~Zh�����n���ţ��	����yG�B{��ͽjjp�V��Jr��i<�=��
Ш��e_q��[��N�[�9v6Fd;�T����ڿ������v�R�X�
`�0�5n�p��p�(�I������dejKiQ���x��c��T!�S��Cuc��8�cʝ6��
Ü�F3�u�QwIr�D�����^�<%��(]S���y.�����ְ1�y�1//�������K��K2Bv��Y +�������DcrGB���S�@�&{*ݱz�T���4��{�;�=̴�@Pg(O���rPֆ�\ef��::Ԋ];y���8Ǳ�(n��w	���\�2���&�p$��!�u�������^U�'p���w����0��˹�Tݮ�v*�����d�V�*A�궈�xCV����3��c�O>R����AܘY�j�tUt��rLmxl��\.����.�-�v�B�}ը=�elV�]��ώh�yF:n�^�(v� �3��KꔮWwr��u�p�}\s�����_K}��;�&r�]J��Y;��mK�Nv������¦��l�z��W���o����B��i���*��?eD9�!P�(���/��h��;�Jڤ�wir��rc��Pzy��FtE-uÆD���oK�7]��uO@�~T@dut���nf�E�4F+���[ -����=G��8=ϑ��p����9t��`D��g�5=J��lI��o��;����
*U��r����F�#׉_�Wϐ�ۈ�Pɭ{֕.�=}�hq� 8O��s|�u���;ŝ_#��0��-L�9�r�������^]e#���PE,�ɣi��@yv8Es��P���{�d7.�Oa��j22���ټఴ��˅����s�&��:�-!�*�eY��{�O��5�gut\�f�+��M�{���G�O:�C�m�j�dgڝ0��|z�*�w3ei=�^��y�KhEv�L�����T�H�j�p���@
�uZ2�39�s1o��:�᝹��//��[��?��	>�.'0�G�}�(��)w�۠��
��嗜+�Ph��v�YI��ح��$��j_�q���BC)Ku�:5��D��fwaޤ����s�Xx�w�j��3�*�L��z��m��'����\Ww�lÐa�~ݩ�3;L똭>RG��ϰ-���= �V�Y��
�)W�\�첱oA!����?�+��z*m�F��>R�/�+l��������fŉM�Ӝ�\��f���"�^_�+s�7\�������$�G��txߒ��n5��e��ڛ��bL;�_u�T����e�NS+��DN���$�(��nkX��	����'�T�Y�F�;[rʻ�g�\�	��폵Ô,08����3l�B�p�&�/��f�w�)2������	��,MS"�=0�[S�;�A��0[[M�AP��g�:0��+ֽ�"j��"��]b�,7\'\-ش�$3��1�l��)ϗ�+D��?iͅT+�N�}��Jk�>ݛK��0T*�&�L�5@���%:��\^�I�io
�si���ù�%�ѻ�_��pCg��n!7z��T�+����� ���Ҹ��,�[�m�	��s����F�������ܛ���ŗ8�x�`�S(>40�k}>�
R��1�r����M�Z�r�#x��=��tC���Rb�])Ԏ��u@��IҌZ�m����VEr�^@���/s�"C�_v7w��<��|].*ո�;J�V�$}�X[���ݫI9���E\�����m�Xq����_M_I�&r7�S*'-̣t�7ʱ����Aۤ���Q�h���[�������������1g�n�l!��O���90�����'wB!��r�%�c�������R�ۼ�����+����J��u҄>Ϸ�����p�Sp��f�@TVf�V�4��ֲ�E��H��r%�rU '9J����Qڤ(qDU��&a���إ����ziCC\�Sdj�2����wPr����`�����W���;ڱ��6wI�n,��[�ۈ�ͨ�*��N@�l��ڿ��sG��J����[W�����9}�Q!���3]ˬr��N�].�ޚ�!#ܸ���Ỵ���X�R��C�vJ.;�6�8��⯩�!0g��!���TX5Յ�u��:b.��c���a��mÝ�iO*�G'����[�z���QZ�%<oW����H+���ތ��a���@=6ka�r�aUN6&�B��]���,.jx;%���$��?A��)�H��Q,��~K��{��V���g��f�1n1�M����S?(Ow� �RPL1�БX��q���Ug�n�\u�iѬ���nVSh���e0���2�j�]!]�yJ�Q�M�u�AZ8��;��N�wWh;+M��l�}C�[��@�!{6�dT�l���J5f1=�nuozT�3 ЏH魰c��ȷ{�3[��̴Cۡ��[v�u���~��>7
f�9	��H��4��A��tAJ~�_X�#U��^�!kh��5�oW�N�?�h��0�p�ۢ99���u�;j�x��(�Y6�]���w�ɡu�PƠXk�<>�����rՖs�&1��:�&��۹u|��En�poLޖVYK��LL�m�'�����|b���w�Y[=G䔲ZX�Z��m��'U9��P�X�U������]�0�dU�^HB)s�c!�WE�n�u�ݹ���ޙ�B��G�î ,����K'�|�PT�rY���\-�د��q�Q#�7�-QL������I]Oq,.�ۿob��>�޹�O�+��+B���j�݊?T�_��{��s�9h.���>?�e<1|�k)���Q��j�΄LX��M�y&:n�d�7��y �Gm0*���3�T�����=�Վ쎭��N�/*v�;���K� ��UhB�O���>/�,p
�o���t������e*�t�j21ލ�;V�c얪�Թ+�a*��B���M���M)���ca�o��ݫ7y�ћ/�r�b��*b�p����6��3���&i"�6� )�,�k[��£U�Ïf(�M�1c��W��^є
��^��L�J<�f�-$�nN���S%jw����c�%��'��}�tB���5&�� �s�w��*O7<����[�"�-���"��pcrn�˘sR%�%j�r��a���P�4�.�:J䔂��Oyf%������6�츀� ���f-Ҧ7&�GX6LLqҒ���=�5��P�m�ՋJ�y�e�asQ[��<(Mw+|Z%��Ɵ��z��/�O���m<����u������oZĖ�qN����s�n��X�cZ�i���*��?e9�!P�<,�������V��՗}<���"��jwQ�_-uÁmW��,n|�H^��Ӈ�K�Ջ;2�c%6��Չ�rS�"s�����ѐ�1���Q��\���MZ��&0u��<5��x�U5�F��յ�_�j�h�f:��#_�&%m:7�t�z�!+����Tn�&+[%��%>���_���Ö ��ŀ��E:�����,��Q�v,o�3pEӲ�+̎Q�îc{ݧ�����O��-�ro��L�lBRX��z%�Ņ��ݰM�XM��*����d&n:^swY!�17���Ϋ�8n�i��mT�����}^{{�XD5`���-}ê^�4����s�|2�n_;�i�3J}R��d��qf�T9#ʍFMU��ڷ踇y:��ʾ����[hޅf�3�N�.�'�j�ػ��z�t=f��	У\���&!]���S�{�ޛ�#RzR؁9�vҫo(G �fН��1�8k��Â��u���l��ɠƵO�25:ac���eX�E��]ű�Q�{�r�)[3se��]�'l��q֠�TUKeΒf����q��뙄b�Kf�c���z�%ba�~x�ڸ��k������Ua����|�܌'�θ=�Ά��[��hzK�����u�)��M�:!j\jX;�(d�$Ft˩.j2���=2��nܾ���v�pN�M}	O2�������̞u�LQ�"M��N_
��ƫ+_ܥ�~q�]���W����;U|��`ۘ�6��V;w��A��-����ql�^J�5x����<��Ќ��Q�̩f��P�N���ä3 ��M\>ό�?.޺Q5��؍޹�`�%b08gI<�̋��	��Q.�v��R�ki���y%�9.!���o�뵚8/�u�����c�q��݋JY!����6��������jGFd��&`{����$��FcH���]Ct�8@���y"t�����+{��.���gk�W��/- s7Xײ�� �qX\�8�^�y�l������|v`�[�Vp��Nw��b���3���8�%%�A����,����MԹ���/��8�R���gN���٦�&q�'��|��<�1u<Y�T�o��탢+x'R7V,YuX��c��-����l�{X��@�sb��W5) ���Yo��Ѓc\Y�W��e�6;�>��m5���s!���-	��3!}ƆTR���^
=�Q��̾�ޛ 8bć-��/�^�\�p_��I����eS��u��9V2�_7�V�����]�JaO�P
����8���fڅ�!$��XL�3_Cr�$r\1�e.�L�ۼ{G�uԃNY=_�]bwO�.s�B�����ca��#Z�V5Q_l��T�+h�k���t�&thS����1�Go�B5b�gݲ�����d-�؆��$��s9�|��S�u�|`������?�����ږ�����:�F�7u��kgn��ੈ��J��*�e���3�ڟl��xX�CV�7+�\J�gb9Rd��1#G��ϩ��e�iPJF�Zj�Jy��l�1��Vq�����Z9�-��V�i����K,���zZ8���p�F7E,W���kӰmX�;�,�ى����fޫ���n]X/�Gz���Z�J#�q����"�\���Z(t������usV��c���@�	<6�3	P]X�WC*��S�E�r�M�/�����"��P2��!��A�]XY]|��L�:��p}b�ܜ*�2� H���V�f��t;���H�	�o'	�4����g�J�؅�`_>fKR��t���"s~���?����ug(�%���Cf.7V���~A�ݯ� 7\�Y�1;+.�f唺J1���Xoڈ��o�Z���U�L`H��,9ޖ�6^�#�h��J�e��nf�8��O��eD�#���=R� �z��J�5�[��
4cx�ޮ�)�f0�h�b�lBn�度dW�d�7T7�rƥK�������϶0���)�qʡ�@����>}l!�9j�9�"U�_F�8��S����>2��ooU�*�\9D�	`��hrr*�q���A��d1p�Q�%,�5�l̗�m=�b�g�ˠ�
`^*$p��\�mJꀷ�]ˎ6�*�i]���j=�����3˔ё��@r���ʱg�1,���a����ȻO��ن�%���+�|�?���A����C;4y�֟y#KF�����&�t�Y��ޫ�W�a(�.��Xֲ��d����5V�������{Px��z8����Wo�gWQj���G�=�����M�:�R�ݐ��yzқ�kj08�sb'U��\�Jr#M���<�O�+�Z0��`��]�^���}B�m��� N��ٗ��{�
��xP��~Z�	��[c�d>[ͫ��*Τ'8U��%�s�B.��\��Pu3�Q��Ĳ������\0�R�b2\�=��XqMp|�`k�|g��y�Ng;}�n��`ʃ1��Ō���7� Ō	��|̌��w�uI���W5�{8������[���Y�2�=O�*���ԷJh2�+��5&��TY����7$l��w��S@F�i\���ܭO?�)�V�1�������J�Y��4 �㒋CJF�-Ż*�.ءz��|�MOF1�KLh����&b�*cs���(��(v�P�}P�P[8.>�1��A\���HƇ�0YA����8Ԗ_�-��	쑦BQ�e���FOˋPP���UP��]��@8;�lt�?\b��]9�z!�0_�k����F�1��a�!
�OLN��[�[�[��6�kJ����:��2a�"��5:����\8d���+K��#��ȁ�ٳ��YND2,��7eͮ��K2[Y���3�u�˟]��<����lMn�s���a��b��|�;�+��1��[;��}8<�|i�5�n2��+��S
�`�Mڢ^]�EcW}1(��Y�b:v�(�Y��R�;V��0�<��M;�r��
A|�9]fB���=U;h�ǚ��}{qm��A�p����E�}�"%��0�0�Q�O�Z`�e�/l�!R�p|1"�G�A3	�R��Va�!Y���k'R2��V��]�l�,o:uu�d�!L�iI��3]A�HQQ�j�I�ٷҊ�nE+K$�����|TTX�.3O�{V2�s��Y1˘��1Ǳ^d�m���L��Y:���vt׸�CQ��v,m��G��늆mr޻��dv8��?]��`�]�4�Sʃ�D���v3�	;�f����.��Y�
-��W�C�H�U��2Pyx+AU"���K/�2��[�|���T�؅t�T�ԫƪMˠ�thp�}>�0yB�_[�(:�V;O�u��O��y�<.(��i�8�7E�H��Uil�G�j�]'Zw�]����T����a��b���K���։�Wu�OD�KZ�����A3���LA@���ܕ�yҳ3�μ�	L���j�@=�V����+��]I ����[R�,hg��7����2�Q�v�kE�����/�^�A���.<���,ڎ���H�Bn�ć;Cc)S��-繎�#{<��Hհ�xsT��.��S�+9)w^��h�-��%EK�prCá�sWPcÜZ}��<V��)uO�%dgG\�V��>E�ʚp�K�ej�./N�{��s;Z��i�e�dL'�0x5�����e�UՖ������3�`+:�X1�	;泷��L�\�d>��ʸ�W[x!bJBe�yc��6,b�W9 ���!7L_먋~�i 5W�#3%o�=�5�ӆ�S��aZ���L-�U�AI���ZՇl����׻ڻ��<�m �J�\.ى��6C3/M_YU�	9:�ѻ��H��j{Ǹu:1G���:��Ki��Լ,r�{)�f��1ER�B��Wf�t�3,RN���L��.�� 4+�v�]_�݃EFoe��"�kX�Ћ[]�MsF�����Q�t�(�b�HT��b�C�e�%[�a�}��Yգ>�\�;�+)�A��]է x��Tn�����,h���t6+V�;H�֫�����p]j���f��[���F��up���-�r[oڙ���
��4���u.[ٸ�^a�C��=^��8�\�r��{�ҍrʚ���OP�{U�����t�vn�J�H�k���S�ՙ�7i\�[���z��b:MM�8����[�(7��1;i��x����Q�2���Iǚ.k�%�ҧ�A�����m�ʙו�wa��3�2�n����)�9��T�� U_%��DFM�F��D+FD�ő�D�H�TQX+2�b�+�1!�S4h�h����!!�CF�����Q�h؊��I� �I&��6����h�6�"�c��Z(��53d��Q��F1X���b�(�%3`���Qh2F�aM&ЖJ1�&��$*HƄ��b4Ah�hJ(�,lH*,i(�ƒ�%��#"�@�D����f%��,T��"L�30�H�X�L�M�A�؄�Vf(�*5	1���A�#RldI�AI����e)�����y]��/K,�o����ˉ/����ԛ��;�yղ����[�o�.N��bt��2��l�B��k �O���>i����w�_�.���5��t�w��H�/��nＮ��\o���.�ͺ]-/�sn��ވ@�����y���I�Ś�r����""8Ap�����|DF=�Ѿ���̊��3��,�fr�̼�o���n�^����k�6�9��r��^֍��Nr�:c}h�5�����\��w�-q���W�^��z]-��ޫ����$B>l؏� >�����q��"m�ukEϹ�}D`��#�;��"Gۦ�y�m��:��o�<���+�����=���qq��r�=~�WMڽ_y�U�Ӧ�&�n-�x�ov��I`	a��"HC)@�e�q��_�O%���k Ag YHs�~vm⾷M���;��������ץ�W�_�u��[�t�zm���ζ�zk�q}x�sε��oj�oy�=�n�Kt��y���:m�v��ۥ_�&�?��~y��r�q7�"�{�U^�>#�|D|��O��t5<��wo��o�|�7_�m����}����-�_�y��o��h��]lEx�WM�m��Z�v���y�{8Y��,N[֙�k 9���ϲdN�Y�w�ݣSY{| �HE�r� v��ֽ����qW�����o���n/W��W���m��W���Z�o��Ś���zA�-�̩��,�:E�������9o�Lo��y���5��/�.���Ә<�|�*�X{����e0GH�(��v��Ҽ��.��+�����x���t���t����z��ǋ��HHN�qZ�2t�@�M$7dY���=zj-⸽������[�tݯ]����:/~��e�=#Ȏ��g�~���Q�yQ���uvޛqo�������ƻ��K�v�=r�U�x���|W�뮮֍�_���xߕ�h7Kں[⸷��}W�o���o�;���\h"3s ����sџOew`{7�#�V�\W������x�[��;�������ߟ�ߛzU�r^����q�U����6�z�˥�7N��\��{�j�-��z���/KF���}��{k۱#�=�<A���^|Ź }�^׵t�u��]��7׻��wn�6�t�Gs��&g���zވ`I#řrt�qi�����z�n6������۷M�=rߕӦ�.��m��UǊ5�}��u
^z�A4Qh�u��A-㣭�����6��ž״3_9%bV��[YJest����Q<1ٮMM��`�]�3/��K��y	�����s]&�*����Ǜ�N�w{�H�@��MII,����UՃ��5�)�B<�Tk+%]s�|��yc��M�;���Դ"�Xzq��f�A	�CŚ��߿��oKE�{��w^���뚽�wѸ�k���Ow�:��~^5���y��{Z+����zk�]5}s��Ŏ��g ���J�\����5jj�3�ia��nםsW�ō�U�^��uv��K6L�39�e�X3�{��� 2�u���ս��ܴW���ܾ�ߕ���o(u;�.��&����}��#�/79^�ſ��}[��n����_.��U��\i�__V��ݫ��_z���ߗM{�u�^�����z��}m�^�[�xf�dZ�2-^�l O�7r�^R8�Y���ν�j��E���H��G��r���:z�r�7��ѿ=��{]���[��QQ�������-p�uǈi8Y�� S��%�ə��k�����e#��HC(<iU�ޛ���i)���`�|G���b(B|ď�k��uz[��ۥ׿�wk���>/W�ץ��-q�o[�+���O˵^��.����[�;����Z+��_�r�7�nu���-�i`�x��z6�!2���܏B5�	N%��#��#�"=�UDE����[��+�߼���W<^6�uW��{mι_������W���5߾Z��.�ܻ]����[�{�r�۰�-@:Xȳ"9��R��u�=��/�o���P��#Ԧ�}�"D!�,�vqŜ�Ll �rدW������ںj�y�]��\[�qs�U׾[�t�x�ߺ�^�|\k���n�`���p��,�C��5�W���z63���Dp��i��~�>���U�w�Wso��n=\�ּW_y��t����Cql.CP��%�`�x����rצ�t�z�~��׋�];WJ�y�V� @#�!��b>���Ґ�ى���j﮳g�Z��`�9G-���������^W9���{WKO]������q���~^����7�����[��,ݲ�H`Hn #�ކj"��3.�7�O�xP���g����*t�.�y(N#�{m�r�:^o�:�6�������zn�s�W���vߗMt�����Z7���w;��W�Z/W|�[�ƾ+��Ӯ�9 �b|F����"�Y�S`����A{.��n�{�~�ֽ�;��Z��^��1J�lTP�ތ&74rfm4���(�]�UX#YŖ��l�e"����H�F��|�s��o^���Ǜ[@��%"V٩���U��]ϲ=�l�\B��S�����*���n�c�;S3�ẓU&�նt���ʮF�}�Y#�#�F�Q �����-�|�=u�n*����Ѻm�{�����5�\��-�t�W��s�{�7�x�./�.֍��z��ޛ����{��[������瞿}��ߟ��ik���C=Dُ�DH�o�������]��/��ݯ�r�hy;��_|����i�>/m{^��n-��/sn���_ܻ[��6����WK~obDA�:c�#�>�xZ^z+'b�׻�~y�?���M^W���5�t�O��|����_~y��^��so��v�����K�'��q�yͺ����Ϋ��{��w��WJ��/M��n|���"G�h����h��<�+��{�F�\~k��]�Ƣ�7��u������&�yqŚRf�� �a��Aod�o���x�6���t��9]7���/�{�M����z��qh���~n׵} �01t�׾��dK�I����C"�+��s�?r�������k�^.7�� �3��@FY��,-y.�@����ܳ�Ϋ��ۊ�?\��M7q��ε���׍po{��[��/B!�����Y6�
����;]���}�+��u���_WKE��Ϫ�ޛ��������-����-?r�+�������_��z���ץ���;k��}{WKC�6�~������ŧ�>���/Me��0���tՍ���D�͍��o/�:�Kq\�/w�:�5񰹠!0�bm4aF-�9f���5�鮟��\�h6"��/�t���z�u�M��n��|���w��w������'�W���&�}�"�} �{!�u���=�:,�Il,)��$�����󧿞u}m�n���~Wk�����+���.��W�M���6��v���WM��9���/���6೯~����N@�s���5�=��#�}��_�V����]/���;���hޗ���q}W�t�ߝ�v7�q���u����,}^���{{U��|o~r�����Kv�rZ2t� Lj`HB,�_P����
��r��,�p�D��}����[F�Ž_z뵿����k���i@���:�[H#�D<n��u����o�_.��ƾ+�~�+��\����/K���*�s�����Ζ(L'��.�v�85��u�L��u�4��K��Yc�����:XJ�<��- f��9j�R�ܨwk2 ��<<����*�Mcm�\���H9<VF@�N�N�7u��d�b��i��eaQrřV��}�	i��p6XRU�#2C����}X)�����և�4_WKt�*�w˯����zmǿ_z���6�����[�s�m�_�nE�7�����������^w׋~{k��t�κ�F����]�W�@+�oe�k�Kv���}B>� ���Wk�-;��yͻoΖ���W9�]����u�����������s�[�t޵��[w������߽W�_����>���tۋx�=ם}�oK�����>#+�~�3����+���>�H|L�^v��Y�L�x�H���d��/��m�_o��K~��+�9�ߗ�]{�ž/KF��z_��WMz�Ÿ��k�������+��=9�تc=��{��h�������~��6�o|��q�۟��^_�뵼W:�9��|W��ۊ��W�n�4n+��ݭ��t��z��CQo��t�B�h�"�D��@���:5��O�f[�^���Z�3�����H��� ?�o�Ia�Z�4� ��l���(��ͺU���;�5Ƹ�z[����Z��-�o_��/k{W��y�m�]�����W��o���\�۵�+�y_�w�)���Ã��V�]&:��h�#���$5����q��-�93^���^.�����W����_��+��]-=���z�鿞-�����Z����� &�l 9 H��(�'A����F����Y�������!�} �����y�o���n-��t�۵��#MLB<>�DN��Sgy�xg���^�Y�~W��܎<��3�K�b�hNo��Uم�3��0e|f���UsXn*���1د��):�|�JUp������nul~�r|��+(��Yd�f~�'f�fNm�,�s�0{�ش�I�w]z�;�$7���;�
�%���G�܍g�8q�es���^'�z^��=�V�]L�[��<��vu��-,���~n�p�B��_	}�}Y*Sp�Y2Q&��T2KqnG/���!@���&�J�陒�`]L���b�{,��ɪCm�U�ұ�Ap�xt��zr���Z<­ڋ��t�<���0�5KEwv	�^�20f��!�o�f.*cr"n�u�d���߳:�𒡩b��E����R�3�t�5�Bk�|��Ƥ���i�����\H���R����o^��[���` �#�6S?^*�eӟ��4Xmk���\d��r;���"�=�љKh�WZ!?�I� ]�]D-$_�g���FtEB�\8d}-�����T����pP:U��׫��I�ꝲ �5jS�"w`���|�@F8��������}�JO,3aq*QQlS[�r�7.�?1a���/�n�i�d۪�E���H�}Ւ�/���/���3,M����Ǿ���'s�MCn��� pB(UJL�J'�/u}�mbM��^zbɾ{��v�g۲��$�����K%2h�&�x]��MBJ�U�U[E��У�q^!�}�4W�A��k���W�< ��{u�[ޓMc��ɯ�K���Ja�[�U���fUl�ܨOK� M�C��qG��F3bɋ��A��a����Fjt8�QA�F�*��6��f>��4z��ݍ�yfMחL4�˺��9N`�֕����S-���\7�H��@��!�Y���wx`/�ܕ�ݕ�TK#1�u1�5�\8֋�r^��;|'P���R��.��BAq�WƵ+���N*����U�#��}	��%|;�vɃ�JE�J�S�9UHl�q֠�TV\v� W׮���0�!_ts�s����]��{ݛm�G���Y53�l�]e�s��b�]�vL�^�X���{M�gb ,ԲFE)�ɸs�����Z*}��9�ѧ�<O��K��+n��D\Mʹ�?X>�샣F٪�"΍�%���/���¿����u'�ٹ8)Mjd���U�U��=}�F�%c%S�Nf/�Г]|�k�0vy9L�w��4+X�َ��(,l�è�~�<(��A�p	@�W���b��3��	�N���5ä00Â�h�9�NgWoll��ξ��Xa�����I�Ps�za#p��%�C��([�c��oj�[�����u��E�8P66�2�T Xv:q�I�Gw�e�(]�y<v�%8�u�J�}�������w�&U�P���O�<�i #��J��p��W;,jX��8��Db5xW��$Y6!�����s �PQU��gŮ�g���<������]�=r�/�N��n(�8*ű-���E�N�=�).�M��v�g+�G�r}���3�ٔu�򱃣����}�4d���_R.���*�<�}���4Gfd������V*��.��ou��������$:�ݲΌF���wb�#�;�70.�8s��y�ck�ܛnc��d�
��S�C�w��Ԟv���2x�+�}�C�&�xc��j��wM��{|�j�Rb�N̛nb5�����f�o],��y���q\5��R���](C>�F�^�b�]��N��06c�p�e�Q�-.��Db^�j�	u��|�Θr���,�i���i�*�Q��vP�ƈ�YV�ml͎��X��8L������ʘ6sƐ_g�B�q2��stv���9O�%P�Y���q�H1|w����`���N�h�{X'�s]l�p�
�\V8'�;��q�7�i`��Zo�L�F���Ʈ��Y,P�v�u�Ӛk��`��w<�Ŭ⚝���F���3󨝥gFt���ƚ�"�)�X9�+*xF��v��Cbn�'��ݪ�]��j�Q�.҆EEm*�������LE�}Z��<j�,��Gc�*͸����eM4�m�2��1�������򿄇�s�p�뫕�dt��S�ǹ�D���V�*W���wR�*�0&�|uQ��O�4�3���ʛc��d�- ���K�)���kt#z�yӯVǑ�M�r��V+��E��Q&h]|oN��w�:\�&����SS���v�+cʜ(����9r���U_}V�:�"�n�r�ǚe���{i��M�N��'bԖ�N�1�C^�ul��j�,G.�r�sQ[�6X����*xq�,��c�~�FNo�u@�u֠�4xG�gfNSir�g��ܗR���Px��nū���X�6�a�Ӊ��ݑ�摚�2���������R=���^5��D��W�A�P��cx�ޮ���c�~�L����
���RS.m'��j�4���y#��k�1�����1�7!a��x}�ϭ�3�-Yf�O��|��el�H�Og�vҲo����/�s��2v	�y{�ɚ+�WwR��a�L-�x����%>��??��J�X��uD�D�!i��un��^��M�Y�&���w��ʡ�u�^�|1�W&���Rr���ಬC��ΖO@�iÓc�Œ:���f�Ӟ��n�f��A�8)^�ʞ���X]=�~��LX�i<��؆#F���J�E�����l��z�g�~ýh��@ Ngx�:��eL<1|�k+a������"���M�/�6��ꂻ��b�m!�#�nν�O����cC�XnT��:k7�IP�[Z���\��S�=~��Mm9�OΧ����e_dT����V���@�V���P(����p<w�e"[��R�������U@��eh�aՃ�$�i$���R��Ӷ������w���P4C(��1æN'$��	����^���C�WFD��{^\�%�p]��Ttmjx3\:�b�T�F��eWB���q;!r�>�c�U��xe��{;_�S�Ӛ���R�c��[�<���=	q+,q>ޢ��Q�\��5&�� �mM}l��E�l=�+��,V]���$R���S��pcMOٹ"�N7��������r�W��tj�ED��Ƃ�v��Y��ON��u	�P�S�7Z:�&8 I�}��#b�MnG��e߭��oJ*�S���J`3L�Bi��!�,�:>c)�GM"���%ۋ���E��N�6�X8\8 p�t	
y������Uc8���NXၬt��r4����_�c.Mm���Ջ7��s�@�<j:��B�D��}�3��O��=-{�>�[�uyh,����WsC��M��Ƅ����G�	`�&&y�Q��r�η�>#=��n�.gI�����~��P�r�����h��т�u@?w��ؼ͇� bj�ͬ����m�g������ei
��[�%��8��_Z�{kv�p�p�=u�]����]A�`�}ë5M� ��^ۑ��ʹ��Ћe��Շ{w�;HB5J�}wh��}o�l��ɀ���өqK(ZR�L���<\�k���2�טf ��}�Qݝ+2�l6�7f�|�5ۮ�@t�-�'�T��L@	�Uu���D�ns���\�u|��`�4;F����{&��Y)�F�7@s�uCxŒm�jQSۚ+�1õ�ǂ�lŕ.KP�꧰�_N-�-|��У\�x�)Uzg���Y��$���Q|gq�+o�f�p��8o�`�s��1�TxpUr�&/6Pvv����	Y݅Ӣ�P��{T��SZ,Ƹ�_����j����J+� n�t���X<p� Y��!h��&*t���Q��>*���ќ����L�N���g�Ua8�Pl2�ED�	�kq��D���[��98[ܮC�S�p��[6Ү|��`ା�gٜ��L�}C�������Z'�?2�����aʮ�C�_Xe����/���rs�7m�p�5'm�yH��.��j�*{����k��`�L�ӳ*f7�Г]|�k�0vz!9L��n��D
���ȫ*X�+S�-�VB�Ί�	��+���/ʛ+*QTbD�t��Hc�#�n��q��Vz���Jv��+k��hgqF�2�`�^L��<v�]�r8�:����Cl��seZ��P����5y����܀K��(*OV�_N)��)�j"�4e�Iy;���W^�mG7��w��t֊�ȑ+m�qV�� ��f�B�#S�\e���R�Z~\3��TF}��i筽/v��1��F���J��y
����R�z8�.,}�I֪�aղ^`]h��--;Lk�:��Cq���Ve{W��������[Q�J<e�h�ؕmsww|�j.�E]�J���5(�X��7xZ�uwLe�K�#rq�d�'^�J��9����vÔqqb�k�l&�i-����eu6�v�o���>�0Ҝ�P��l0����r�p�q|r��VB����$��:��r*�9��!n�@��[�n%U�R�wˎu��8��X��$� �(�.���z�:5�AS���bQ��P]��+��PT��\n�F�2���A��yѤf�����T�ԈetԠ�Uӛ�F��Fx�0A)��m��8�c2�����Gd��&ਂ'Τ6ۃ�΂T�*s1�'q���쳧�u���$��K�T�[���5\AE^�)�Yrb���)��s�B�,p]��� Q���x/�e�a#���o�u��Σ�H�y��`'+��z밠u8++d�&�R�fJx�jm6��#Q&����N�u�ohE�9^(*�����]FqX�Q)�q0,o<}BW.�s.u��F�\������0�Xcj�/N��L&�w�ͻZh���O�7�V�H#��ySM�7Y�b��['K��lC�}X�͎����]T��i뼵N��Pf�'[����x�q����_s�S��S7��ɡ�������/^�o�gM���#d�hbp�ڨL�S�2^+qo|�x��o
y�$��i� jq�V_K{���SU��P�u���g7��T8ky��}M����O��(��Ww���N�waV��F'N*�s��9(ڴR�[tb9\�����qX�{yp�s�;'B�RU��C�:��2`�^�V(
��5a�:<���%�4k���$�4����A�v�%C.﹁:�պj��G�YGC<�9#�xJ`19Q�k.��v��ԭ��l�4��&w�jpݫRF�ְ�"����S�]��w�Axu�(i62��p���h�M���k��d;B�m�W�uXV	c�#�FM��Q�q�K��t������FM=&��ȅ*J�;�����!��[�W��lwt�^E���(�9Q�Dr��%�4���o�=W�;�]���x���N׋\��C)�k+J�z&��v�͝����C���wV�ٰg˖G|�o/��;P��WZ�hIC������L/���v�����3�vۢ��&�\k�5�;�A�~��'��"wv*f\�hAG]�s��C6N�5�¥���9�8.��cne6����G��
	�Ţ#Db�-�&
�,j(���,	Q��5j�"�ZF�F�Ţō��QA��QPh�h�hd� F�QI���53�D�����Kb#Z1cF4�+F�Z�4F�!���lI��V��m���5*�Q"[Z1���1��Eh�h�536@4lF�`��V#R�FL&�Qd!6��X+
�Ab��J�
ɦT2�X�(6�i�6��Z�1��i(��Ѩ�h���^���u��}��rƃ�7z���ŴFH)���#l.|m=�4)�I�+ޙY�Ԍ�ܖ� �;�4�f�wh-EQge�>������:�ڙ��κ�,��j�v�~�#��I�2����s"�L$V�ľv�
����ˎQ��9+�y�(8}����r0��84�T+�rQ����L�*ԥ!���4R���cU��Yփ��rb�%;�n���&��N�	D�9� �O���،c$1y]��iv�XB����DV(a��oF���Gr��X
n��6 ʙ%q�Y����.;��%Uz_���b."zW�e3p7���k��l�a�h�ѭ�Ý�dN^`o��/W[����ف����}*a�-��+J�$0�̘i'fJګ�)aPי����{T׸m�yt�b�Rk�
�An8�O[jh[�7P���2�ķݎg�fv�t�z6z����3_',j�V���e��2au��?W��0�!�8N_g�yRx���h�4x?��b-k��,u��aˋ�"RԨ9����4��'�}�wd�^��"Lp��"�6��ρ��'_4o�wPr��^����Q,4���
�	5x���\�u���<r���sc�������ŋJ�qV3�N)h	ԑ4�U��n^�4��y�c/6��~�
����v�x�zK6��H��}` ��]_	G�C�-t�<,���:��$�����Ƌ{�*3oL5���.lL�y1����C�F�?�3a�%�/�t��h���W�eV���l�r���#���\�5�延[1M�
m��|7r��v\j}�Xqd�˙c*�Χi��%HjW�e��L1	e�R=Q��Wbɬ��ŏ0��t��n��@��B�P�t� �#eHG��Vk��{���	d��U�(��¯�?��g�O�֘K��� F��3&z�Jxޯ+�!����*8�w��;;s�ꨚT#�W�!�c/ ��N�zn&��KIn��7b��"xv�T��Eņ��m���q,�½��|Z���|j����2�������d�� ��vj���nɶ��^���7��W2��-�zRUcx�+j�c��;Jd޶�e�:)E�N�-��4�DV�ݔG�ŒE�:�WѦS(F}��\;%;l�)�_���W�-�>���c|�$h_���A�#ܧů��1F�S��xe�2�g�ټ��AL8I5��bFdn:�6Tj��
İk��}��1�+	�/��3�<�D��9���0���iP�]�op�#l�����&r'y<6`����n�k��RE~\[�����!޻ZT�B�%Wp�cR�R�R>�຿�.�={�
���V+�0����s��gs�e�(�������Jwn���r#tmF[����J���7�`�}�Gǭŧ�6���"��z��)d��9��DX�uGN�!i�򢾕Ճ����8ܷ�hs�[�p>��HZ��CP�屑	��7�������U�И��M������&�<F�>f?7�7/�$
9Q�_9��o.�s����>�[͇��^�a�7-ngt�;i��0��P��5�ǯ�N��ԙ�η_�L<1q�k+a�����ON�����Ǜ�e����L`�N'$��	��ˈ��W(uJ�?`��O���`�⎳d�	ݛi�LTج{�4����<�'d.@xe��g@�Ϭ�t�.���,2W7ldtF����jF�٫�{W+R�)��X+��h�=%�OfG]��w������S$W�'���yLB���pcs���i���8]|���̬��A�)����-J/�����'&0��C	����t���D0���f�c;����d�$��'J|3m�+}�'��� >�Wq�1��uS0�R��,P����>jK8%Y������o��bU��.8����y=��u�)wsЎ!���
	k<D̽Ce�_<P,�,�WB�]�d��:�c7�_VS�m�S���W+�����*V7p��.q��3C�)l▀�v��1:At\L,����9c�^�a�^�>P��_}U�U}�j�#e���~��Q�@B~%�#���)�V3�;u��C�8`�k]�bL��|jٝ���R�n!gΏ��L1
$�n:����ZHy��FtE|��&��eb6�j��R�J{�s>3h���3�I~M�R؉݀^�9��ٕ/ΦL��{���S��zSU��?\��5hd9t����Mցn�����M�w���M���0M�@Iܞ�z���R���%1P�
���Pɦ�p/"� ��P������Oϙ�Br�+b�{d�R��wE���+�=Ҹ��=��5PB4SR�]�7W�&���g�93�� {�P,�=t���܈}�b�}ePw�oB�r��`�A����nЉ�����bo9�GhO?��ّ�i=)�	�2�p!Gl:�h͋HJ�\=*�3��/�4:�N�@k����j�P�Z��>���eX�\��kR���;T��8�PV�*��X&�b̶i_bx x���e�fq:����a��_)�Г�\Nd*���/��-�7Y� ���A\�g@�g$��-f�
ӿ���|���\l%��GS�v��ӳ�>/�O]�w<1&(a�=�u6��v�^��I�87�սy�7�9�y򋫣9��`g��!��V���+�r����C�2��ZeZ�v���Vf���062�E�����=eq=�a &/�<��Ja�Y��N��=+m`LV�6x�f�[~�ۜB[����50���ܛ���h��e�d��H�/]��s�<#v�G�z�[@ef��F{�3$}��у��&���%��̹�ߺ�	1P���ƺ`ۘ�6��V?�*�<Vtfv>k7�����#,���"�J¸?�=����3��w���/Jީ�����=����tE�_ŀ��ɫ��f���#��I�2�ʱ'�,���3��5�����**'�G9���Aé�᭦�g��a��g9�"<X����T{���,Ӧ��T�Զ�+{��8�@��
�k늹nㅹ�|u9᤬s e:�&��SQ@�lu��c-Ṗ��Z�MZ\>p_U�cgY{�Dg[¾�N�8�pCg��o�MށnlA�9���A�a��}:N��J�a3�+��\tn����5��%�!g.�����zz��׼ ��Η�s����rH:��}�r�	�pԪ�]�Wo��ء��}��E@��rI���ڐ�r�aW�W�$:G�wD��,�J7v5>��ᏳEƣ}�3������W�v �Ľ��}�kk��Yq�X�bε��s�K<��Ӆ��:R��L|oje7|��6������m7��z��Ir�0>����y��������7w��p�qI���ڠL~��@ũdN� ���4�:��jW_n�憞�x�P���7��v�-��Cr�&��W���d�@Ʌ��c��bA������9=X����CF	���5T�Z�A�X�,4�H��F�?��6��|}p^�
�m*�=�=�[<�OV�p�J�Y��&a���N~h��wPr������]��3|ϴ�oiԌ�k��nV�̖J�oGdEDZ�w�KUn�v��w�\� `�+�ڿ��Ż������e7v��Ɗ�.e��?uGӴ���4�5#K���1�S̰I���b���T��;rWX��˝�\>w-�X�
RU(`G}FP�Jd1��"�\�[=-� 5Mˌ���+oXGn��1�r���z=�T�N�m�,P�~�V��n��m�^��Z���X����b;>��|1k�t�N�zo���D���m��N����f���'����,H����Mu�K6)��_��Ƥ�_��_��������Fs�<���ז��>��K��eB��W_�����Uo�<[�����<$f�ˤ������x��E^��i�4�5�	�&'�!�;���(Z�%�J��[�k�U������븸,�z;c��(Եa�Y�V�wE��HP/�Ù6�d5�R���  3�ʭW}����:�F��Be_ъ�o�V��\L��m�ǆ�� +g�Ȝ�8�&���B�j/fV�Ws�Q �d�$�ᱦS(FB�m�����
`T������s&V3�<��uwTh��j\B�FB$�"O�F";�LG���.��J���a��իYd�I�SpФ�F��E�"U�<��˝'����J�҂�4���_��\b��:pjr�ʅJ{*r���iя��z�Ԓ�K���(���"/��X��-�_�ik�^�֡x�{y*���!�q�p�R��Bj�M�`,/�ʱg�=,��ϩ1yD�ެ������٭��A�:vS�/�q����\�Js�6>��GwKM������Ҟ����J�TkE`Tbѳ�s�c'�q:z7�3�N���N����z��;
Q�w�5h���V�O}�V���@��
�4�Gj�4��*���@^�p��e�)쵅��7�w3S����'gQ��ouo�yS��F �eWB����Y�>�F���d�z�V�r��^�ٜE���MN$e��
��2@�0�-fEm�V�5�h����=j�Fum��̩��m>Wg'Al�+\e�
�{kEY�p�w`﯀��qu�W �5�5ݥ�Ȩݨظ�u��a-ט�8�5��<�0�U���=�4hŷ��ϩ'2�ފO��:�W��P�>�TW�"pW�6�#���pR��J6=��� ��^�Ƞr�\al�_,�nyܱ�u\܉��*3�h����ި�|{ص��HmG?l-\�4=��CJ�{26�ΎӃD0���&b��J��S��B�;��u�����tT	Ca�䀯x+ -�`H}P�Q�:��f�b��>V��CRY|sO�i�T1�a���Ҕ�����5��`�Q�@b~%?�fn�G�S6˧?K�r�ݙSP8#�Y��o*�9ӝ��_�,}��BI(���̀B.����o��v5=��ene���������=88��lޖ7�Ħ��,R�g��$��/i`�ѐx��2u�Z�����+����H���b�� h�MZ�D�Ŏ%��@�v�&�
�c��o���W`^zrj2r�" ���q]<�ZU�
!Q��5��\9`ŀ�T��#g�b"]��.]%H�[\�?8<4v~��m`�#��;�+�O+��A�S&�n@�wq�0�Y+fgI.����E-��C�k;�ԭ�WN�{�q�V�x����[����hm�t�W���ȶ��S=��M͊��w=�>�*qRfі�qRO_
N��G{7_2�W�&p��f.�0���cy��z�8#��X9���}X�	�X���u}���}�}�}\���vmm�̡��$�9�zF#>XU=���������v���)=�7쳓�l,��ᳺ���_>��a�7*F.����U��V8W��oy�5*�p��#*2$̗��C�X�鱁t��8\�q]���TI�:��KZԮ�'nr���0�ͮ�#_2Wsz�^vky4dx� *�T1h�8��u���SCt�nO��dU�҉ݸ3D`��E�ϴ�/��u��T�U�E-�v�
� ��膾U�*����{��������G�a�i���7�Qwݘ�i�w�P}���roh���,�j�e����V�n��,r�r�u���e�v�������I�8zPKO��~J�l�����\t��0xc�].��,Lˆ�^�Uә���a������CF�*�'�\ |+��cؼon��>詅촍�VƔ���%�=2�h���|1����j��A�g�#�I�2��{�ȿ�L$P��}y��Y����1ϥk���.��J����F3\�=pX�p�*U
(�r*��L�eu���js�
�[z�8$=ܠ'KϺ��V`6�>ϴ�6=�:������n��Z�mk�:��O_sP%1G�jv� ��vum
��*'.��癑QHj�Y۳��ٜA��ɺ���Wm��W�&��N7ɮ�n��$�E]����Y�EZ�Ұ:�{C���O�`��c�u�Y���[v���j���*����nㅹ�|w~N��o�s g�ณ�������ӱ�,f�w 4���l�cOqx��#8���rt�d؆ʂ��Mހ�FS��W6Pw���JDd��I�t� ��<W�e3q��6���%�!����[��fŪ�ݒW^k��V���SnfE|�E!�'"��8��)l��R�s�~�������zsU�g`�T�p�ҝH�p/���])��1jY���� >�
2�:ԻG5d�[������f�qу;���N�s-�;�S����x�����6>1�2-������&��+9bɣ8tGk޶4^��S,B�!�1@�lĉ�u"*0�pWn_3��7���B���:������`��)����b v�S���;�9���M׽����E13Zs���B�P��ʅ�G�EDZ���j�n�v���Y,P�w1.읓7�$�{N0�i�no�����"��N�����Ϡy�:4Ҡԍ,��1";u�ݷm-G�0K�4m,�t��S�vP=�#��{����|<�q�g$S�3v�S���*髵���o0�E̩�B˻f�@�umD3u^��{�	%+��v�Ʀ�ye���km�l�N>���
��@�б�R�m:�f��j1ga��)�P�HFef	+����X��Neu��ޫ�̭��J�a$�5�A�_[fc;P�C��5�:���w6�V�u�CJ��ZۂH��������j��YΖ1�.s�rSR�놧*}s-� ��q�G5i_j����1��(Q�y�Q;��1���ES�kf>��J���*ofї�������7��`/�{��ʸkk�Z �os��w�Y�(.+M�ڔ�*ðh�۷�: ��
����6q*}|ۮ��T4�x*Փ ܲo-��u�n�۳r��¸�VX�+�\��|��c�q�r�L��mE��G�*�����/n3/ ���m[�棝A� KeJd9�ʉW�.���ް�v�I�^��v	]���v�wXiMSF�#^�KUǅ�,����K�YS���x+�l�/��T�V�4��5�:���|&���-�8q�Χ�*K'J�󖝘lUÌ��yL�d����� Z�%�����ɋ�C/1<l!�9�����
��.���Q��BU3�_7wgp��E���0��4�J��[VI
}qV%�M�2�O�@�]\��缛H�<�sٴ0��eb�w����y�JsK��+B���{E��j��鑙�k)��̬S5L���_�
�N�y0�X]�:g9�n^^�� �]��;2���r�)P�>�F#y��n2ĵT�c���7R���_n���ǰ���9^p��Xk���֒����S�Wy���2���Le����G�N^
F�9Xz��v^c����J��C-\r�v����)���:�
��
�3���_3ݤQ�t���G4�Cm��B>t�̳qn�O9Aо*l hv]���U6��d���ftR�Q�ʭg2�ǌ �{�+���:������<��:Ҕ�:@�8�y/��'jeL�i&s}n��u}�uS��
�9%{����0v�˻r�Iq�
غ���O�r
S[K��ъ(V !4��2G�l�*ڵ��㵌��7�0xmv�X����[0T�Qp��wP��ٺM;�	D6�|��=;��D�H�N�upKl�!�pl���{fo�F,�f��}�*�o�GX�BN���s�V�%��'7�s���	�]5\�^�~�a��z����A�U˕e��?����2��4�'M7��3̀T����Y�mw������.�p�Pf�"M���̍-h+Moufʂ�G!��:6�==V����*7̛�:S$a�� �Z�:�]�A��*�l>R���@�"���iO��Z6���4��B�%#�3�.���ڻm�d
��P�����KF(**h�(�d�(���&-�j(э����AX�V#E����a"�"���F��m���h�(��cDF�E���bѲj#Xɍ��4cTh�,h�m�Pm-���j4�h�X��F�b���Y5	��#Qh��lh�$��!�ёb�*#QF�b�lYh�4&�F�J��6���L�F��LV�65��
�F+Eh,`Ѷ���ߝ����߯�λ���QcQu��w���z�e
�.��WW�frL��+G[�z���B	.�Z��nS}���w�z<��_�}�}��{�>͞��R���ܜ&t���U l!��b�u�3�	1�Ҡ�����f8c�����%����C���i�g��p}�o�R�F���~L��C��K8FwKh,��p.�ʺ�؅����L1�����MN��'�G�Q%j�[�ԩj�݅{\),�kW��D�P"��mnL��&:ݡ�lu*n�\��F:i�}Dmª�O�rS�}9��b���'Q oK���a��$R�X�8�����c��a������F�T�F1����Ǹ�f䑈�jd�G.H�J��S(B�Vl��Β1�)-�uOlN�Y[쾯J�j�5f�9.(8S%)�S�$L�}4.�T1����1�V��uV��#{dcL,���}�9���9j�8Lb%Xu�J�Q5҉ڈ1��m�#����پ�c��Wt����1V��+!�����$������*��)i�q�
�H�ýA��ޚ�����ْ��kaS9^���5�\��MMIQ����9`ip�hhv~vgo�i�0%�d>5ɯW��D�����H�j\�U۳IT�vzr�I��	������̺�f�<������腐I�����&�O9�k�d�;v�.psA��W�eet��ƲS�D��؊ۻN�Ծ���9q���������-�@�?4@��>��ߕo��iܮ-�9Lh������ӟ.t�86��N����uؚ�ۀ/���xyf#���'�St�\WR�x�ˌ�w�F� 4*��U�5
�-�8������J[1��fa�jٮBՎF��^A��z��I8`c/��`��׸�05T���:�cuc{:��Tcʝ(@xf��W5��}���[����<֎�د���I;�\:��_����eu��,,q>�~a{��Qv7ؕ>ǡ_t��V�E�2\m�,����[$W�'��ה�+u\ܛ����F*�SU
5�� ��s�-*9���I�MR�����%��ofF�Ύ�@نc�L��Ҧ4\h.`!���,��WmPL&40I��e��EuR0�R��ĉ|��mIe�ޝΪ�γSԪ6�����L�@�W�J�	~=��}& �q�g�G�UX�C�_M��yNS�_7U�qu<�<�7E��ڭ���F�y,}�aU��]�.�H�a!�qo�d�c����_���(���i�џa���scM�MT(�ֶ9;^-�s_L�GF6.�Eu�w( �M�@�U�]��no!�����5�.��4jqת��ԗ�:t��Gg(�8x�ʶ����[(ݣ6;�ŝ��v�Q���;E��mv�#��U羏�#�qwv��v�6P�F�\8d���f����q7�7pxؖ~�F< K>�:L;��F��u��A���5���S�5�u�+�MZ�H��`D�&�@�v�&��f;%��
��c�ܤgv��_^�� �.��H�+�����a��ۮÖ ��#�Éuod�dt��Z�zL�<O��!���ۊ1,��+�9���w�Z[{`#�S&�['��&-��<�y����!T^���i�$�U�Y�WC�uMm��\Ϭ�����k������uׁ���"��P�z�Ρ�����Mʜ]I�N L�]	�
�<8*�V��K��\���V�A˼|�11~>f��+~��8���W`�K����]�N���y�t2�`����4���T.E��hW���FY�g�f/榆�_5�a�ܲjg ٯ<�k|&!���)qs�+��&o�<���&��ӱOw=����ݔG��h���s^���M��e���)�FlU^�4��a�_BS̾w_1�a�mV���R�kz�l��������wh�p��WSX��i�	����j��\�f����)W�����ހ���Hz���:��*�_��v~�A]1g�	�0^�{B65�Zw��ػ���n�Un�K�|�����ǅ]�:�p�ը������1�:����tOe;�E���}5h�A,)�~J��9�k���Ѯ�3
��:�z����E���G����[]=-r�Zv�d,P#]p�>��]u�c�s�D�8i|��׼��W�\��O:���.7v�}.����u5P�f"Dh_qd�`�9�"!�ہUN�(6��O*t�<v�yK�5����v���?���u�DBWe] ^m�.��,�l����Z�
��P���_���st���t�x� �uHH]�oT�z'�/e������}AgE�!����DV(�7�uW;��,60��~o����p���$���^y!?;����R�%����qQ�ŝ�jܱO}���Օ:���R�o^\-u�
��(F\�؍`ҙ����	������ʼbq�5>�]��s����fc	�V���E�+�I��$�ɶ�#Z�/��6~�ي�]Q�
=���g��������?u�N��L�2�`�CS��u2l�z0��ܵ�w�.�U�:�-��:x.����$�1�E8��\m��K�'�;$�9��ߗ�J�u�ER�T��D&�D(�ֵ����(Z�����DH����
+�������[}�ܓ�k�ef��с�[����v��$��g]^�^�������βs�}U�Oޝ��:X�������Ֆ/檘�Z�3I�P8v��d|����3v'8���k�ƉN��n�B�����:;e3q�}lC�2���ꩃ{��t5�5zڎ��1�ͱ����=>
�'�H^z;"*"ӥ�KV+pev��̞�rn�|�P�Ra��Nc����{�}�U�
�j��#f��p��N/3��=��/���nZܳ'����<kٸ�q@�t�Y�Oݸ�Y�*��I���O�AV�Є�FU����l7p���֮B�q�N�,��+�X1	�Ψ�u��A���e�0l��3�qs��D��U'�ⲑi,]�WUl��v~t�]�Y�����@y�'=7S��\�7�t�fL5�����_u�I_��C".7��nL�� �[����jK1�������/6�}�P�]C1X�׿(Ni vˉ,	���*�X�8�����c�ۙ�;OC�ض��V��tN��N�"���������\�"�m�O��s�<+�z뮔�͗6�w���� z^�%�b���EU�&�O�̭B�Qx*��ٱ$��ܧV���gh|��4p��]���b^���W}�̤�J��fnLC�-rՖfvv���d�u���[�ˇh�|z���)�]M����y\��DD2�d��
��ո~ґ���`���A�2̍�2R�'�d��O9�f�v׭��~��aHj�������e��u��9j� E�W@u�"�&�>�pw��&��1�3b�ʝ=�)�D�U�L��)zb���w�Y\3�~��2^,y�Q`L'PDO�Q;,��H�O��Ւ�]�Qt�wa�œ���ӛsl�m���1ɪ�7����^�u��ٌl1T���8k}�f�ٹΤ�7=%PM֍(9B6.���/��
>���9;�8����s�gg����a\�݈}=<�������.(Z��^j�'����Ύ�"�Z%�ܠW6ڡ|�l���#���َ��P_�x��\=V:5l������'wDf��CE����q���>YgΩ\1.u�Ȇ���uo�Ǖ:P�.��4C��<��3إ�HK��Ue�������ê^V���?r�z��`��{�K�`f�����p� $Beq�5j�k;���l�K'��w,G(u\ܛ�����v�6�9N[ӫ2���˖�;AJT:�c�c���Ks�71,�.�\��{%�����S����J3<��HM�+�U�9-��&׫��v�tԯ~���k+:�\I(����	1�Į�4ei�֍x�!x��Q]#F�f�RcN�"">�%ul�i_H�\�'T:�P�4��CJ�{26�Ύ��4C.1�&b�^�Ί5.��m����n�v��&����,v�e1�B��a��S�e�_>V����:d@=��b:b2�()��8{�4���,� �V�`�� 1?���O31�#�]��Y�7��0�7��*vV#�z��8`���i�9�ү%������RQ�� wW��&��2!���#�Ӣ�9o�Yέ���:"�k�2%�1ZX��t��7ptؖ~B<W'L�jJd�ك�G��]|�b����w[܄qT-��V�����
��E|�
�^]����o��`��|V���]�}��>Ck�2����\7�5��}�n�bm;���y0�"f?�u�;\�n;����T~q��v,�;XM7p��}՛8���B��N������ڟ/&c�����o/ZH����Ú���'�Q���k0-u@�U/0��b/S�^N�Y9a�Z�XO[W+��H����	�3���i'�T9ݮ{v;H�Q�Ex�/,�^1�	Y��l�>���\����C�����)����Pd��c������Ǌ�M����[���n`�h!�
<��<dV;��5f���ܗ	���ư�ﾯ�����yw"��b�W�nڗ��ƴ�Nv\���ޮ�����L��~^�X���gc<g�搰_c����je�9�|�S��F�ۣN���:��M�\q����)g�F�ʁ)��Q\����l[�[m.��37.��*{�lb��#w/���W�]��Q:��҆�Z�l8K���I�l:��u����yzN%cK��eBλhOeX}�;,�+~Z�0$M�W`���m��P4�M>��'�kg��TRd�0-ǐx=yC,�w��q�MC}���E��ٝ�X���z��q���:c�0T�U��="bR��y��Ĭ��g5�_:{5���k�#\g[�z�*˼�S��{mu�^{�79���i�ڽMd+�e�o�ٷۉ��l^1���ڌ��
sFS{Z����dt�}�`0JZ(j��R�_ri\3z�U$FB�٣���|�3�Hd3O���|�d�qE
"����J�G"q-��t*�T�sH��x����=���(E��[��z̖tAw�@\6�F�ɕ���T�X=�sy�ǹ�uS�̈́�v]�Dk9B˧��c�um��.����������M��&�gt�7g�}�}KI.e��i�N���f��. ��yvg�=ᶪ2B��Y�ꋞ��Itn�o���
Q=�l� �\�~����,޽���ך鮝��h6�J\�m��B7�Ș�6-nk;8%�]����(����}������j�u6�2ځ��_���:�̝�;��S�*Њo�$^�s�g��������j/j�E�B�S�8謃Ժ���ȹ�r�����ٓN?�ű6����*;S���/O�q��us�h
�I*�����7_s��w#ت&�*0O��������c�kgqrR�;U�������O>>!l��}��9�c��W*i}��:q}Y�:���mB��Ö���۷:b��U ��*�j�-@�_T�9�����������lTB��&��\����ݶz���۵"�Nf�q��@xp��Z!~���^�(��`���7CAm���]>dve�ai�{��:2������O?X��K*g�{^ܻT�U���//�E����K�n���Q�����:��=�]�|)�4����&����R����o��z�KAxʝ�U��e�*T�7��7���&��ޚ����hGOt��u�c<�A���줱]P���ŧ��ko�p���Fo�=�=?����n�����:��>�*I����M��-�.Jbi���V�����q�=n5�r�oa�2�S�wO�Z/�)��Gx�jWK�;YWv1���;��昭i|��ʈr̢P��h�d�v/S�<'�����X���in����&_�]�w��(��x����k��W�{u��-�pwrM����� �!>�P�a��]�7��ZzxF�b�S��k�	�/+��?�ˈ�糚��<w	�6�3ɸ�Ƥ8lBw�w{�u���g�y�\ʳ�jћY�s�s����z��ڮ�,�������{S��O_�:��m.�>Bs��O�>�ߓ�����x=����{��r$n�������!Z�0�bLf�[�U�9�El�I�WP%7:-9��9b�Ѧ\wP�eht��Iwi��󞛎��WN���Y�e�d=�/iи�Y�Δ��A��V��sq��!b!��o@d�ޖ�Jpu�a<B.�k:��Fe���[)��st��oj�Ya�����Ȗ��
�l�*�>����t�:𛿞-���0���
�A����E0�7@u�5�WZ�V�'XY@���ы;�݆�guf�8�I����k;%䡗�t���Gi��m"�d���k t_&7�� I�xe�q[˵��� �����;N��)s��2��vR	:���;�=F�;��2����)�yr����;��CNp�v�)���ٲ�.�<�w�M:�K4����gzT��Ϸ'*�(0�J\����+��n����u_�,��Z/�r)l�Q�e�$GjR��!�k� �HSW%f��.�U8+v��9M�@UyBX�D�z�Hhѿ*G6�U���}�2�3nޭ-��)X*��a������	�Z�X3�#6(�N�Z�Iq^"�U�qg�6�ޱ E#�j��V�*_ow:}K�E����܃<R��4 �jd�Ԣ�n�	��������;@��f�f�nSƮ�]�m7���s�D���Ay�b�$�2��%	ޝ��;޻,����P�x�c:��� ��J��i��t�n�>�+RB�SFڼ��8�7�+h"	N���7�(9���7��ݽ�I�5�68��5ci,}� &�t�pG7�M�c�͡�ٽ��vXۤ�Օ��$]�R�T�iy.�i����I�3/Q~Eg� #R1�s�:���f%;R%N�LXsSFM|�(�v`F�zy#�(ܮ�!&����4a���S�4��|�D�N�w��P��mNC�>���0�y������:�}p������,�F-}1w1\�R��X3J��΅�`�>��ň<�{��q�w]�J��[L������z�U�mpr�o���*�ӄ�'e��pnv9��*��0��W��oj���[t�;ǳ�.ΦnXwr���e�f�ި�z�(n9��p���e�tG\�0>ʖ����@:
�M�H�}!<�Bo%,j��;C��{[K/H���N�;�*:�Έ�&	P_f�@�$�wGڅ�\b�#.-��2�q�v`�˚i�6�V���&���j�[m�R�P��`�r�O���>L8�n�n�艒ڊ�Q��:0�7�p��W\+��wpѦ��������B4[5w].��R�<�A�W��=m-��.�G�
D����;L�К���8����֝�U/(�1+��ޛ\��P��݅wZu-�Wۼ��w�%Gtv�X*�J�(T��uk�5Մ"���_�i��_u>Y$�-F
��OQwZ�Z!�>yL�K�H:��M�E���$����H�w�]�ZXŤDQQ��f&lF�1�m�j5�E�F6��
EF�h�lɐ����cd�ZE��Q$cQ�آ5l&�c�Qi6�1Xԁ�h�+%��X�����Q��X�b��b�lQ���5c|q�b��5��ڊ#E��E��6�*��	�أqW5c`�d�EW��i,Q�j2�`�9�3���j,cFƬl��V�￷����&�^4�3�t�$zkTi�ǔo��j'oZ\"��K���n^n��^ի�<��u�Ұ*�Nv8�/k�md��w.�����z���:d����w�.U����gQ��i�͸��{�N1���;S<�/�u�����!w�[�:;�E�kG>4����F��v��2.����g�oz���A,h�!�\�:G^�>!X�`�_N�5��+������o;m\:�V�!��T5rG���v���9�N�5J
Z�t�#�~�)!}�T�:���v�G�gm��������|���}J��N����u���ʨ���3�#w)����8{Q9m�J�P���Q����dl��p�fm�-����R鯔�ˆ����W�{�ߗs��/���G�k����EvƧJ��z��V�;�f|�uB��e���׸�h�leC�P
�vl�I��Z���5j_o8�5;��>G-ἚJ|��Ro ��I���od��5XK�H���5���U���2Ǎ��c/����]M<-��),�r��2oP���	S�e�� r�0�\�9���S���\}�V�2p�����υt�p���Sz,���u�uR�wz����X�VV5&���i;�+lȋ�735�<xq�3|0+\��˶�;��|��.f����I�:L�L��Y�1��w5�����L� �C�-ɩ瓺�B�Tdf\����eU}�F���5�օNk�9�Y���y8����S�x��8jގn'S�M�u��V��m�p�ホ	�TF�7�GVzR\�6� E{D��ü�y�g�Ć���M7�R��k�k"Qڌ��F�ZB�8IyE������{�����Z�o���4�L�e=|�s2��=����s�Ve�ܺhˈx3* ��Φ� �:-G_.f�%sb�Z�t.�nh<z�I��pޮq�^����YE\��Q:��҆���Tlr���)c5)��q�;"�3��dI�x���!g]��Ϭ>��J
Y�������O����&����P�7��}:Ol��v����0Wޝ;���b���Tk:�eo9ek�<���Y����IkU^{V���Ρ�wWg^J���3��[&Yӱ��s��qq�u�{��[wP�/x���&��&�us���'l�wd]��v��m�8%��|5�Y�tJDGx�K����+z�����Y�N(�
N=�+�L�.om�k����񦶯neO]�&�G3��V_�y�y�Sxhn�-��=�S�����o�R��_z-�&�%�&���g��s�m��_Ǡ�z(o5�r���[�b�g'�3oL����4|�j׻��r}ܪ�b
Z*�y��-�ɥ��xs�NUaj6�mC���௹<�,�!u@��᠔�jyv�G��VDq jt�]���5C��$k���|�ĪD�r ��C��m�15XXǽY���o�{ϣ�>�Q	&n1�P���ȵ����v���M���;fx6��]���jU��'SQi�5�n�YU�ȑ�0t��2�'u����V�Q�X�u/0���{E��vy�����|�f'5���H��|���k%�Vn�����@�U�a���V�}�/g��;<�3��sW����;h�ťdƺ�����$b�:TC6�v���3�����q-���4��ᶞ6���̮: �����̾x;�L�{�Tʖ�������"g�w�.�gU���t�k��W�$N�#�Ӱ�a��De��Т��]�}U�i)����g$iw�`uq؍��=��1E��5�Sкz�N���Cm[S)1��_6�{�g�vr���ΆnR�<8L�ٞЌa���R{/R8b��Q�S�\�rޕ���1�Y��}������RĪy�g��::�rp�m8J�k�c�7��|�q��DT*���Dk�Г�������f�Ӳ˸범�Q�ۇ���p��M=69��&k��5k �Gu��)�������#�%��/gKOd>��7p��l+��J�su�,��x���KT(t�|�~*@I���+�U�j�Hz�Nd��uKzz^���ͧ��gS�r�r��!w��X1�KEiMf@�3cU����Itq珣U?��낚LV���	�{�f��)F�p�Y0ἇ�BZ_-Ιq<��B-�=���������
F)G�;}�WF*�m�KK�tr�\�t�\���b}��ő��:dFQ��s
��[KNԴ��u��\� Z*k9�-���y�[M7B&���{	�؀dv�~���'MW��^3��l����f�m���f�7&����6�h��^�اBb����/�l�J�˟�Njmv�����}'RL;ƻ�F��v�#vQ��:OP.��*2C���o�J�̞y=�W;}	�5i�2���5�vxu�S�
��׵��~;����*�=��f�y-[��U9̼��)�iA*����N�t���9뇶v���F�5��k�b�|W�9�Ͼ�S���
���Q��̖�u.�Ƈa�:�E]4=EeN ��p�w�	�ũ�6��:Ws�i���/��X���g�/_[u�q��n�Tr���MO�F�'֢�7ak�.����Y��އ:6y7��ny�'���\����n��܃���tj6�%p5Ҽ-�����;m;���Wf[���ԗu�iO�l�W�y��*�'e��PU%*1���{�N�"�lc��ыc�n��'�kz����>U�����߅�U�nE���q�e<��)�PF����w<*���(����!�˧��YJ���_fԹ��0�{�IW�	�Z�F*����*���@�f�A
��/�e��S����.x�j�J��ӼhV�r��W��� �� ���kN�pS���b5�f�Hj�aT�G�\9v�G*�������X��ڇ��ͥ_
?wς���̱ƺ�e��Ԥ��N8�u�K��r�.ֻ5�uE�2��|g�/^��z{�$\�_�C{C��ϑί���-�l޽�O�T[c*!�7�|n�d��7n���e��Wݎy��N�{��%�3y4�|�x��4�M��;6��W��噙�3�(�D�CA+\�O.ڿ����mDr�j��M笍�����2�ԛo��N�k;x�u���o��vyᓝ���޵]x�>�x�
̷ңKP��w��k�'�C��kh;G����\�d�ٳ�R��{|�vr����B�|�m��k��'�_k�z�l\s�9�t$Nl���WU,�;�Q:�m�W�nڗ����/MQ̩��u�k�g��6����H�z���wfc��zB�yڢkh�l�'�\5[���)b*���`	�;�i���ԅ�I`�o�5��ᰰӝbC��&��n�ʹU���4M�z�^�q�S�;���_
T��g�ꙺ�v���6.Vz}/�1���%:��Zy�{��f��k�Z�Ɋ�Ó�:S;�h:��:���ls�N���źb��uCl��j�Sǻ]8���|�̢�`>U���@��X�|����z��u���ֱڹ����1�4���!��z���P7�uѯ��5c\&��e�U]�֥q�ݍ`Gn���Os�i��]�q�b�>�����Ɩ�m��G���1>�0m�*끩�x�M>r�q���l�E 6J�Y(%y�Rζ����c�vt�We�B�R��zZ���i��i��mΎ�_���c�&1���]�UBچ����u�첝�5�vk��|2"^-�w�����V�ަ(l�|��\	h���Y��K_M����id��&�X7Ӽ�{����FW�Y�D)��(b�Z*�y��T-�b�V<;ɨ](�ĵ�71�6��p&�63(��%*����O.̕9��>.J��v�Q�o�Hm%��6�;��F*D�!�:�XP�����n:�20f�5�J���0���w>�IJҾ�����ƴ=��
�u8��eH�ap|�%F�����L�1�D���]x���2t����yL�-���<�1�����v}�+'uu��^ue�[����Bș�޲#��j�.�䏱�Y�w=S.'�m\w-��4�N�	&Cn5�#q����4�L\T���	�L[�\��q�Ky�9�j�V�к�$�{�ᚄ���k���ʸ|�j��|�r/�V�[��[+2�'��ϣy�^ջ���p����y���%x�8L~�P�x�S�]}�d��P3D��+�'Y:��=P2u֘�;@��j��S�_����t2�ד�o��ϋ���F�d���n$������q�p����L�c>u����C�O(���֖�C�U���Ӭu/i���.���@���,����彙ѳ�gŐ�������=&M^��y[�]�H' �W���m(jƺW���,妟_ι��kvm1U�X��g��o$����/��y���}TV¥J�syoCy�iQ�ZZNģ����5�}ܱ��P(9��:R]
�t�h��t�%BI�C�q{iYZ�IJ��ۮq�voл�����㔁¸���i�;,�f�J�����\�b���D�N�ڈ��ڮ:����ۥ}����I2u��O) B��U��8¶v�[c
��Vy6�9��;�Ls���D;G���VS�(��=VY=\�zZ߻;��nO|�(���ԕ����⌧�;q�f{%�s�.��;܈N3�3z���;���AKDs�Ni2��t������ON����IC7�d�)62��(���nb��fzDZ ��e�K�w^��Ӻ��"�=�������q*Q�U���`�XYWg�g�[P:��96�j��N� �>��a��q�g}`��ytO�C���[^���u��Vë��̸��y�k��������C����}��_B�&6utf������t���2��^aůsV&#�6��0�v�f[�j�k�:�{gS���f��U��V�n!�]J���zbTR��W"�.U{I��K˄�kY�>��Y���j��ժ�v��qؑj�:�W.''*�q��b��3͌����͍͛v+����1� u`�+��3�#l ���F��'�0:jrR[n�������)鮷Pֳ���|��9]oe�	2��qBBj��Q�&�fp�����jb��,]�o2�����u��ħ�c�mCT�p�̢��L�� D:�.H��.팱�^r��=s��Ss���(����J��>��?Vtl`��Oy�_v貙t���ʗ�Vv���.�G\��iBQ�WR��)�?OAK�:9ʜ�W
��]'�k����� 4s��bvY��PU|�R�`��_%��H�z�S�O�yx��I����P���P`>U��qt~]�����f&h�q�k�����]Sܞt>m�8{_<墒�:{��F��'Sv�\�Ƶ�K�g;�mc�t�Y}ic�z�:�����(+�����ǳwF�WE������]��[�r_pSak��LV���E[c+�R���8�s�%�{�]-���<�h'��D�縎*[�k�J�|��,�T0[5ٳ3kwz��ѽ���Y�*����j'�m\w&��j}�\�.ϣw�|�w�w�L*D�G!�
t:�ɨ��{���p�4�;�P�������l�3�K%]̺G����G6e�]KF�UÀ���R�Q�-��=~�*ڇ�Y�(x���ry��o�'qOj
z��W�U�ю>ɶ��6�mn���z���5&Gn��t����m�lV�ʖ�QfN�qeq�Ӷ8�%�
]����� M:\H[\[�C�t�=��α� AƟV�X�1]M�;+0ueH�Õb�.&���X<4|�@�:�1�.W
�l�*꿛F��{n���M0��i ��G�h��}\�w@�¢����-��M��"�^ �z1�#�q���3W^�#�p�1	5ޚ�Y}[��~9���x�����%l��P�Ӗd]�l�t m��u�*ބv��%5����.�.�W<o�]��pObJv�-��V�g�*ű��=�f�N�AS�w���7�Z���f]&�A�r�펓вn&ۗvCt�u�'f����S�Ưx<���<����D
6w�3h��b{�;ҕ[NO��]�1�4�+Z�ܯ8IB��:�M��\�@],n� �;ѵ�l����;�uΝ�6AW���&���?`g_eަ���Jh��!x��v�U��@��>�q�`��p.��P�ܴ��n҉R��@V�)ejZ�i�O�V3:�8(�ڵ��AĲ�sE��[��4ft����2�T�ڢ���+8vJ���&U�4`YI6�+�V����kJ�ɝ]H�B|��ۺt�l��_8>�ϳohЬ賐�ӈg��{��i��;��{�)�\N��AĆV�� �=�aIR����Z���޷c�ٙ�{+6>��~�B�T=��Wܦ�V�G�*@I��&��V+�e�EF-�oq\z���HH���XZ��:,��t��ǏjoK"m���L��GO�ۣ���ˢ��}w�g]�]���Z�����]6�@�ݒ.��a�����B�ii�0<�tOm�M4D�/�������J룴K�خ��S&^����jv˳���Kr�d��z�qꃧE���=�
�2����'`�@(�չ�<�o-��^sSZL�7���Z�*,��N��H5XK/��+�prZ�_!��R�Ox���mVM�X�zL����\�[�Q5���m۩՚'NZ�hβ�g*k(����Vѥ�b�t�)}�P���	vj��
K(V}۪VƵZk����wC�wqrw�:���:�B9�w�����XŌkХ*��3
�]�0��-��+�����R�H����T��G�˻*��9k�g�����壔/�1�0���z'��M�F��ś��3��9��V�m�ܡol��e�����h"U�o�hN{���w>�M#���|�J��X�)�\�2E��۽����q[�vF����.]urL��b�ז���G9���@]g�:�g��N�6i��\%��Ƈ2�MD�@i���5ƏVF�8��t�]Y��b�(�M��شi66+���E�IH�Z�k���QDZ���*��5&�-6-�cj4fV-\nB1�Z-�&5%��+b���k���U�q��U�sV(�q��r�#��-g.k59�IQ�8�ql[��pE�q�-�j����q��sQ�W��b���X1I�b�b@z�!ԕ���j�3lW�V���t���ӯK��.᮳�:����ZRބ�`s!�����1�ԯP�y�4:T�s�͝.�w:�~Mc��Tj�`��D#3���7��}��sg+5�^I����V.���O����u�\9V��O+]ϵ��vn�E���c�;�o�Nֺ�ֿ`���z�i�^8Z�Z�}Gj2��7Ÿƾ����/,��ە�&�C2�t��m�
��j��iڙx�z�'��r�#z�Xgck+/_��o��G!�E\�ʢnr��!��gK!N��]�3��_�}N�b�-<�WwH~��d,��_5n���{�9[�:��1T5�o��7��������7����m�M휔��1 �KD���c��x��99�v�W[�7���y`�v��@j��3-f��l��;z��|�5g
<��T�k���e���4��Yǫd�����T��_5c=�E|���t]:{4�<k��K���:O��W�[����oxU�;-��_�cX��՘������7��ޱ��͠��v��|��S���Paj�7z�7d������H��\�}\6�N�h��ִ;F�5���#��6Yu,vZ�y�ˇ)ns�򺭾z����)pn-��񗜢˵կl6r�R�V��cs��P��I_%�7��r��ݩl�^��s�a)um�,���z�EDZc)�3�1�R?�F�v��c:u���M.���49�|����p���o"�2�]�%*	O�~�}C�PERs��j��������5�g�|;a�P�!1�l�5�2�i[�7����Y�3.\�{W�w=��0����|�`��#q���TIo:{rn�W�>���s�j��P�[�xi>t��$�{�N��λ���1�=��qu�x��_ˬ��d[C3�%�T������jݵ/L�e8Y�w+�u�j7��{\q��4���iv����V�}�2*a�0E\�	H�7��ծ
��q�u���������eAwşM�J����kٛ��٭���Q=��'�	־?{�$-����-�q����d4<<�=���W�u�ʳ�e�Â[��@�j �<�7�l]4���{x�StE�ь�n�}�KKhU��yq�Uޡ5y�;���W"&}ko�iZ{[��V��'5[.y��҂/IƸ�}s���ʬa@Z0�c�h�4�޽D-��g
z����|4s��}�k5W�]Խ
�a��6-�|Wfl,齳�gt�M�E�ޣ�l8�[M�A|l��Mǜ7i�W]+������M>�\���+qO.�`�G_4{����`l�S���g�DmQ��z�ȳ*-湻�u���]~��]���qz��Yp��}[~��e%�B�.�t�Z�u��sK�sQ*�@��7)�	�8YOE�)P���>�����������q��R�^-�`�o�t�O��f�nBq�O�r�����XN�w��Ἣ����j���y��T-�낚V��P�Ʀ�S�f	�׌B�i~ɄQv�k{�T�~��f��檑m����_̾����}uL*��%��B{���E��P)Pۘ+\�]��ɾA�}F�L<�����̺��omѹ�֕Tf0�'z��cf ��摥��'ϧ�������ӛ=7rAb����d*��R��±a�Kl��r�Z7��(_%F(���7�ok�.�dֺx�V��1��T\�E�76̥:�L/z�ɭ.�Q!tJ3;*�f�|����{�[h!�j̜V^臄�])n�X�R�U�jô��\}��p�H�sX�Z�vbؠ��7���^���O���y=s*���F"�s�s7 l)	�:n�kc�w�m�p�Q��Q�Aߟ\��U����F�z��Q s�Ɯ�Co���/i;�*^_�8ֱ������O�*ݫ�\�o��<G�{��
�Q79_	le�������62"^���/7����� �].�nә%��h^��̣�!󨛜�*\@��b�n%sa�z�'��_��O���w��9�������Q�'eB�g�,�5Ù��3�Ӑ���Mh��=�6�W������rt�Tw��x�}G���m�B��0�z�>MM��oe��7���)�W��[�`�oH�S�V9~�/u`P���_-��k���S��|��σ[q��C�[f҉�>��@��X᭫إ�7�֨c/@�n�[X�>�r�/䵮�q�Q��r��鐞ȓ�w$N@���o}.p��m��|�*��V�ޗ��̬+0	t{��	;�WOe�ƥ�wE����{Ӟ��6��J���/�����j��(��g��WGQ��i����{U���"�c)V��l���k ���*0����3L���oq���������|�P�<���uB��I�Ŝ�u�_'�FfA��W|ҷۋV�nY�GLw�H�9����⥼6���|\+IS�+����ynGea�
�O"�2�=��_�sS˶�;�mƩ��Ǘ�����%C�I�m�w��p�M� �W�[�7#����!☵&�L�K�����|��MI���n5�s]��n@���m�fX�&�E6�%T�s�����[P��ZN��8f����k�j���H���݃/���@O�f2���ی��ޟ��<�Oܽ4=4�&��������WF�ŵ��+6лϏ9�f*���V��Q5�;��xˬ�C#rb��N�s����b~���2� �Y*���Xqm�xu����~[��og��h?�$��������_����Ӽuzt��tr�y��:��Y�%��-����p�WL�j�'+�Yy2�l�亨� ����N�Y�y���51��YWRX\:���e��ۯ�w6d|�ѵC�����&��_"�w`楼-��=|����^j�(WU��q��)���܌�0n҇c�Q�9GTLT%��C�պ��]��r��y�U�ͪe�\��F㩴��Ӝ�5�८W|5�P�7��i��5��g�Q�mWK����7�@S�������ʾ�)J�\�8|�z�&��9��-w�4����Ю��w0z��%�!�躇Of���k]R� ����/�g]�[+V�U��n�B����QA-7��t:��{Q�+'3�	:�qRL�j&J֞�g>F��WdpS�L��4\�Y�ѐ&\��-D�H'+F���&��7���*y�D.��JU�"�<��#z��ՙ�x�ϝwt��C�P�3P��� <a�B7�	�CohA3Ud��'@��˴��ES�Ӛ�}�qܶ�0��4�`�Cn5�#d!
�qy�oi�+{s��!h�-�@뒻2�ٿ�V�.�V���N�NQ'��oHd�u���1���Y�R(Wu�v}�Y����	�T�]M�-��|lbʵ�rb��9Hv�ee����Nu;*>���xQ�	����A���C�B����;�����('w���D�/�`����\�⠱��U�Ct�&k�+
ڜ���.�'&�t*��i
���*�p�}qU�{iA�VN~���/7�U����1�hJ�N��g)7k���?D�����Bo���J{_�u�X��|�wSJ$N�;n��ǎ�\/��\.����&9�u�fTAw#س3=�ۅam�ٜ���Ij�	\:��c��S<����C�{�5Ϗ�[S֑� =����ð��w(��|S�}+�n�j�c�_alW�sb�t�\��W��|�el�-Q��	�s�0*���vY��	F�]������&�f��u��ܭwm+pk��Y��)�<�vx���������S.v��t�W��1lp����{I��kz$u� :J�*����/��7UQ]�pCarE:}��f=ގUW#sm���j��)D��t$�T]㟟Y�#�)�Im��=�V�������Мg<f��(��}݆�6 D�A�[k�i�[E�^����Ⱥ ���*₭|�9#��uL"���D���T�6Vk�].�Qo#��}V�J��:�5|冲�0��2�Yȯ�N�&Ae��ӳ�R�᢮��8�G�vg�2��x00%�X�R�k:�>U}�!�w��7�e���n�Ψ[��4��޵�௓cf���;���v�y�j�)����}5˞�"�|���s�!�����
%nul2�jN	}F��F�wv�ݭkr��)FYGh�j��5_a��ԝ�N�w�����Rʸ{��d+��5�ѽq1	����Y[�q��f��Z�C}��25�0���,b�-����Sq�J�]�?s"�����%^o��ջܢ߹����3�<x���j���9z��k�5�<���+U�6+����r�mۏw:����y���a}�1s�����F��Q�8�g�%Mׄ��M��|"�K��8����Q1X�ڙ��K���n��o�:�\N8<rE�w��!o���ƽ9}�IP�1F�bL�͍��f%L�
�&�Hnv���F�rxYk}~�8�X�u�ȍ�	X����i�ᛘ�����ݒɿlRq,����Η]؛���a'�����"��E�i�n9�eD�`𱷓��0����s�[+; f���E�X{X�P�r��`ɠ���*՚{��2�V���h�{�>V���q_AXX�N=��R��J�嚰-���yc��j��=�5��rP@,�f�����i�����t���I��0m��u�5<���ƞ�t��ި:y�T'Lf(��W��lJ��j�����בJ�r�q�{>m�8{Q9m�J��C���[�6��;�����n�s�jk��;t�Y}{	k]��:�۴�,��8�e����G���q/�-�����P7��:��ۂ�W޽���l S�J�������p��J3�!w�`�9����⯖��}��-;)kW1�x��tnc��øM�k�g�Y�*���Z槗m.��V)ڭB.rv��h��w/�gv��|�n5�7�L�!� �Q�h�"��h��p���)�˶��t.x������)���#3�Ș�5:ܹ�j=i�Å9EG_4{���jVeNv���Z�i$�؜3Qm@��<���Hz����i��5 T��3F�7ة�������	nG[@[�7J"����c��.\��Ã�U�q\l��P�Iv=��k���t��m�����[���+;{D�o.�wM��:�vX�V�*�h�/wwC�On�t� �kV��KD�p�l���3D���Z755{V�!){p�ƴ%�P蟫]�쀮���(w��c����-ԗ/���`�hƢ~�i�fz����`�s�vF��/^���lm��[�u�!�X|��ȁ)�5!]������B�8�x��k5
�=��'��ݻ>��2o����3]&<�u��[��4�����V���TlW�smx���x�,���v�)��V�H�nv�4
��JZ�t@��|�7����t����K��)��Tm*���\E`'`��g�ꢔ��ֱ�e����S��3�b��K|�m�r�k@���@t�P`w	�gws���Of�r�}E�9�O);�]k4�;Y����uE�JR��ς�����j���	�
�5�����|�"�?C��<O�T[c)�3�]�Y�`��?�R��~QZWOs�N��g|��������PǷ˚�������oWK��16��'گ�t3
ۭ��uďv�11�uc[���eY�v�{a>��i��oJ�\�U�np�noT�=�}�t<R
���N!䮷�[@Z�$����o`�:y��3�����,�s��듴�+j@+�z[Y7v�lt:�t�,tQ�-gX)�!l�WY��h�qU���:%����F�n^I�]��Zl��
��h��҃2j.��(T�=��e��=�ܛ/&>|����(��Tu�ohtu�T�f�-5�5����֠�՛��i�_R깫����$t��f%��T�ݿnm�ȅs�yp�Aԩ��Wc[5��c5���Չf>O�ɶ�I���k�(��%mˮ�����5�E,a8�Ĝ��}]�v�3����eI/���^a�*Ԝ[z��^o롴T]In�p�l�4r�rFH�8;#kT;�t�י{�����ƨ*#;w)�fhgJ%��J=�6K����/�,*��m�j	*艋��1��ަ�w�����}ծ�r�ð�P��B�
R�_Zn����ʾ�������$p���;ig4X�}�t�����h��I7�P���Πuc��o�Sn��Ѹ��B��x�����ģ�Z��J�m���-�b���r�l4��z�˖fJj���F>��'vE�9,�T��h���*����4��µ;#�5��3x����֨�Txr�u���ݨ�T~�O^�g��%��f+�K}���yJ��4�F9=�5�8�A<鋮oZ�r*�vWt�]0+X���PE��1v�L��:r�<�;�U��������.eœ��nd9����k?�ע��9�X�1���u��L��<KS�['w�g*C���]�Q��x�deQ	7��m��;�ஜp�����&�i��ة��v��ER&��"0=�`/��/���n�Љ��O;�0��.��hȒ:b�����xd����H_/�+�E�;�{)i����ה��8�6xs"-_E���t۷�;R@�V�oR��|f�#@�Qs��c��n)�0�e.b�v�*�v��A�"sd�6Qэ�]M����%�|}��M���pV��f+|�Nݹ����e����3��KU``�G�om�9���2f��ژ�"�*a���R�L"��Ѡ��m;�ގ�Ļ���P��.�޾��rT9�-	�]���T,_:�|2����f�y4�����U}�0������
�;'(	����y[����}5Ӧ���֍^Y�OgR�P�\�c��{Q��\�n�*7|�6Edj̃&E[�t�}�lV4�.�6�P�C��6���gp��C(��a��^$f�{]C9WL�IT<�EG�;m�k���J�9����R3�Z��v>0u�*1#���Iͼ˺z�Iǚ�(�6�@��2ލ�������{����	 ��	�" "+�Ŝ��j��j4`�[����lZ�(�\�qr\T��ʍƍŎ+��h��.��8ы��.'9��#n%�l�5�s�qQ9s\pW&��\q��9��Z���n"�Z.9+�qj�\%q����9n7��6���ƓI�r#.Nj�\�2n1ܹs\h� j&��s��9ȸ�|@�(ۻV^�ݯ̸к�s&,��.w-U��W��GONĆ��9]��*�8�rw2��q��-�9��i�oU�]˴,]����r��&��7��{��7�Q��D.����ž�sm��{�=�'I~�ڬo�x&�F8k���a����R��XR��p��?b9:K�UX�m���p�m\w-��4�N�I�Pۍ{��s�rE=�Q|R��_K^�<��s��#�����[Q�դ�\8z�\��.L��:��S^�k�UF�#X�khfuK�ܜ�����ǹ{�Q�Ӳ���fcjV�-p�\=���c]���2E󡘍��$;�����\[���\�q��E�s����kyu��y?sF��c2���j�8�����%�ݻ<�㠃A�tz�Q>w
g��_&�{G.hM�铲U��YVZ���|B�񻟠gT���X�ca.l_Λ�0aC8Ak���9#�_�Y���}E��:�'e��	p�J�6�fA.���^E����G���Z�<��rF�JZ0>�`wA��9N��b�d�C\�j�i���rm�e��WK��}A7p��3z�<�!`K�{���E�
n1J��퐧����u����uHή�osJ�t�����5���BDԗ���WPs\/�9����3�y~޻x;�cy�ť���u�^��HCVL��綷�;.�CA<�p��4��oP��� :`�!򨝔�L:�k]���t�\�V�q��5)��A��p�����)D�����ǣ*�y�g7a}��K����5�������f�nBq�Q���3���-�[C��K0�ľ\��15
��Y��u|������7�c;��67�ESw�$����A��K'���L��������|���%u�z���f[�ަ�pduC�G�;�|6�
�56�tԝ����b;i'��4s�"���қA��øƻ
�9"��6~m|�����e�|mS ��s����RC5,��q�;�����&�]�WU�Ȟc�Z�.mr�֋�y{���\�_t⼮N��������k<�^�,O-������2��B�����phOc�i#�¦���w�pޮ#���"�Qt��k�<X�y��p�V*y�S����u�_��:ت��=F���'�
 ��V?U��}(��l����[��%m9�b���n��|[)��l@ͽ1�WV�Tf8ؗy�A��9L!Xj^���HX���8�Q6��'���ME�&w�8ֳ��z�/#'$���&�nփs�s[4i�C2�t��u79Qy���TOՏ���n����D��֊to'��t�wZE���_Q�B�*P*��ʉ*_�Lv$�n\nlPڵ�j��={�69N���_�ۙ:�c7t�{_ǥ���2��wQT�3�%�sԖ�(���;5��vڿ���j2���τ�U��S�Ib�և��%�Bl&�,rT�[Wj�c[ˇ���Ɵ\:Oo�[��O܀�5�ٛۀܩv&�w*Z��s��J��ө��'��5���<��ø *ё�rV�/�����z\�IZ�������s�EOԧ�Vsݫ6��\�����~+77:�P����0>ih���B�X�m!��X�E3/%=�,�p�7�o�B�E�!O��SA<�j'W=BҪ� ނ������
0e�hM����7}���;�*�ǋ8��v�q����`b ���Y
"��:��:���k×+��x���ڬ�똘������gif��:4r�9l��)�w/:�q֍*�W�pO\u,0�eEn�H$n���V.���9�L>@x�|��r��@)W�@Z�7�PO"u9���ܬ��?��P�����6�8n1�P�T���Cd�Q�Ϯr�fL�g��W���MDM����<i�=����Mƴk�&�Y&E�Ԏs��e���Z��c�PV�{2���մ��\BN��8fځ��
��vBs5��OV�c���M��-�@�U/2�������ڷp���]vm!�	��*�+H�V�t��S�:���=�iv�a����Ѩ��b�p[�.����E�K�Z�
��q=jڭ���tk��ߊ��D��8�LA{Z���.vT;o5,��lr��HWǵ!p��m%�׵�nPv����B�	&I���"��WN'2�F҄��T1�IOy�{ӽ��ltY�r������1����&xT�
�{}P���}#[wɧ����'�[�gjWd�%.-է�u����׹J�b���}�ozx�c���PS!�s*��͌���fU�x$�@�e���l�Z}|�A�on*ʲ���X�cΨ�]�J����(2��t8V�-�����m� ��i�N�+nr�)2�r�{\��9��l^�ӄc���v�����O��]�P�T����|��V�r�yeqk��Ku�.�t���4�D
<��*�;����:{+�RP�+.r��q*q�R���q�>ȍq�Qo�T)J$.��|T�����Z �r���ِ��}�l��}�S�Op8��T9FQ
c�JC�Q�p����5��ׯ2!�3a&��9���	���f�fЊ@}��+㻵ؕf��������	�{�k湚�������
�5.��������F���tPp�ɏ�]Ak���]�}�is>��0v��5[��|p�����6������/*��ŭ�Am�e'�y�jU��h���y�<Lͥ�Tލ�p�C4ۃ�eV�!g��;��]/]�����e��V_!�1�WX�իJ^�-p�[�:���B�/���|�1Mb{1/�B�yr˃�Mf�Y�hS�B����꼛��jv�>k;�����B#�Գ˅N�_����ݵ)7س!�������f��|�Uȣ�1et����Ù<̳}���6L�yv�X �J�H�A\[c*���6�guvoxӑrwl"c�
 I�j.#%!���E�s��}������Fm7���Ӵ �J޸r��8/˽���Ss�%�]�'��3͌u��ݭvk7�y�M�	���v�o�{�L{]N�����acb�.l_Γ�qG^���غG�{�7��d���j�weǧ��A��ʄ���]<i�ö�u�F��Zx��GV�֚s��}�J,�w��vG,��},cM�}�󘚛�š�Q��&�٭�;��Pbކn��T�	�n_��}tUz�f'���,v�+�IT
=��_p5�2J�V���j�����q�άv������ې�gS�r��V�D�]�!�������o�/�X��ߡ����P��7���0��xo/D쵉_n=Y�1��dw5�4<�N�yȩ��2�6�О
��#_�{4l��oum��r�G�6�����.2Vewk��W%�:�]����7�?C��'�\|'NX=���l����i��LJ�ky'�Ö���3�Z�=xli̾��g4	��e��6=�S"��읺���Y�ϵuv�[j����\88m|:�B�5<�j��O�]ںG\��5T�4M�B�8}�jL;��k���r�\���ps@j����F���]�\���oj5گ��Q�Ny7���h�)��b>
�1����z�=Z��麊9vmby�)m_\ru��Ú�x2c��*5� 3R�TKV �%�b�;V�L-��v�Sʞz6�S��i�]�N5���c�}p��.�_��8��﫻F����k���&�A�/#�D�c�q
e��C�cgx�Lx�:��s�1���m%�����_8B�;2�c[Yu��N,S����V\N�ź{Mv��͘�����; ������ ��t������E꫏,��v���n�)���dRd�B���\ZT{��l�٭�Wk�q[�x����=��l�Rg��[k��@�OS�� �ݗ[4�ҏYg~Xq��/��ջ�x)U��`Ր�"!ƅ6�6��4�|J�Iw�oJ�;� FuD�v���G���uM�ě��͚&v]k*v'�d����
�����WV1U�<zӣ�-3M�#h�W��$
�3k��j�*T�j7��U��}�ڛԝm=�w�t��{���{���p(l�B�.ù������٨r�%�nк�Dbc�i������ܭ{�V����_T
1�.��!���o>J�N~��f2��������sv�������leC�x��߻�1�J��ϧ����_��ź���یѹ�Ѿ��Ѿb��!?[g>��x�d�z!�נ\zo�k�2O
3)��E��X��/Ľ��,���׸��J_���B���5~��"|_�����k �6�dT"�M�8�T�m�V��\^[j��s`������!*|o�Q���]Ɇߨ�P�>���j/a܃��"Y���}���nh�,q9�1���Oe`���^��c����~��}��=2�5:��$^=��|^��p����z�/���b�eH���U�\	�0�����������
?����g�8�D�����Ur5:��j����U��~ɡP�m��N0k�v��N��2�]���B�F�G�P~��-'���8�I
'"�g�1�RB`T
G���9�c��.����.�f�f�1���M�)�+�
V%%����2֬A�X��t{]МS;���;���B�����WX�uԳ�3t̷N|�-��Z]�X֑}�i0��ܣ���%���Z���/�[.���~��9�󺍽��Q��8�l��P}0�3L�dr�N1���e6��V%q<F���}O2�tm�w	gʷ�a�pTs��f����_���9�חx��6=.U�r<��� �o���+���S=���s�FtQq�>����F�w\�W����_�t�𿫪�&��m���φ�������O���\�̩>��sYݾ����ܩf���=Fc�O�1u�J}8�*%�;yb.��E߷��Ԭ����(u���b�l#�ޞ>�L��C��qrK )�`�TT�V/]���Ǔ���\z�������17n+���Zr<���F���7�yQ�X|�?G�j$�'��x�zNGo �޺�]�x�����+�>�$T9��\u�t+�z�ۈ��3P�Af�A��:N��O�rB��$�$�/���:���>�ʣ��[f2=;��w���&߽q�5�#�jM�p��>K|yύL>�$d�q�UʻǶ�={���j�!}�yY�9�Xy���;z'��`��z���ܜ�4Bz��v;n�r'�Y����=�7�l�|�r��p���uh1)�os^H쌴(�0�]��7Ìɲ&ip1�Ց�b���\��K�Mc��h�C��Fn�.E�Z9V�ɒ��sB3�خ�����on�չ��N���d�}f�Nኗ��7Y=��;�mz�𿟕܏Uн�]6*�z�\��z+��K��-����`r��"��ީr�k�YP�P���.�}�+ǫ#z�@�{�����{�h^c�]�~�=6�~�ǞU��̃��Ī��pvaTO�0�^a�|�=��s��Q�:���μ���~�q�}�ԧ�s�ˡ\l��Ӓ��4�f��ĮZ���4�:�c�{Gz��TuK�t��~9Ԫ<��{Ld':���q;�&��#�g�ۃ���~+����rz+#�u>�f}(e����:.*�6�X��#�R�x��x����z�g��F�g�~����(��{*x�������(Ozk�Dt��O}~\6�~��l<
��h�mz�>���X�[c���^� ��>�3|g�*w��7n�n;�Bnw��I�������;t��G���~�=����3�G���mω8Z=��+]r�>��vmǟ�L�J��}�8}�]��T{���r7��?:�웮
�%TB�	2K������z��VE\�f�f�k.���.�3� +r�t���ۗjZ�ȭd�%����!��+�e츟s]yƖ�8[���ǤI���Zט�Ї0ҫH�� �&�3��DHȡ�/"�u�ծ�-��9\�f>q-�a؎��K6̓RS�A-\u�����emH��7v'��aJ��벯�W�m�����9"�Hj�1�!�״���KR�U�@�c%���~������0`ngWV����a�{I�Q��ڔ�:�g5esJ��ʝ�n��ZSFX	��B�[5S�뎃��4���2D&*��SFS�6�z:�Z�[�(My��p�)���n��J��\�κssq��p�ԝ�v,�Z��ƀ���������f#��Җb����Cq��kW^���k��C�|��Pkf�K}{�n�Ld�8�9�m�7�F��B�٠'m�cq�sE#��b8:�w���ƚ+r�Z�0��cv��׶�G��HRݫ4F	���Z�B\u�ťv��Vw|�3����ݻ�]��S����u��|�Q�n�0�W�,d�u�YV�=Y �WnQ�+���'��Bq)�.����W�����W�j�J�u��m��M���hF�|-<�+|e�Gk��N ��FѺ[堻n�U ��͚���F��Q|��MgT9b��%�;��͛	��mV�n�:�<9��5��V䚃4��8Dg�����:�;�U'���s4>U�l��d5t쑚�MUs����qD�uz{��^�x�ΔK,\��h�7��/�B�"�}��T�J���@ݾ�u�o�1=���}#ZIu������%#nm�\
q�>3k����ܹ*K�Wa3�Ë�j0��ڬ���B���ֻ:ܳ[*RnJͅ�������,6�ju_PaJbU���$���=��i�<���;_ˢg����?�h��v�ˠ�uD���\sw���H)�]ˤ����͐JobԺ}x�m[y@	.�����l���N�����]���S�v�
�n���ͼ���ٶ�m;iܫ��ۡ$�[�o}ռ�Ε�Q�{�5p��k�BM�]%`*�_U��-��N�`睘�DpH5�J�[�`���黥���l���peʉ`��J��w��1I��C3X7H]�*�ع�ƒ/���څ��/�z�\�l>JL�Z�hX�0E[ ����i䛆$y)#����C��Z��+9�N
�U<rշv�*�]u�YQ�k��)�tJH/�se'A���[33�*��k{�E�G���Ϗf����6��/B2�1v'+��F]���"T:س-:dI4�1�n]}5H-��oH�+-��ݬ�X�h��@kvv'Ґ�7`�F�����\���Y읶Pe2�Ý\[�Ce��1�;s�͡Ѻ쥷L��8��)L��S����Q3��*T�{�ʕ1V��)M9YAu�]m}]@ (
�+����9�&���9�rk��*R8�68ܹ���ܑ��JW�-s�ƀأqW(�0Q�0��ӗ1�Nsn2Kc\n2c��\\����Ŝ�\�И��1e��+s�ѳ2IF�b���RX��qr[�����QE����n.-qpRi���×8F0I712����H��R&M"n.IDi��˜Y���@s�ː�H(�$��."dl�JI4$$��n.MX�^�w�>qs�O쾚��Wn�:RF+[��]�5+V9@�wy���o6@�|j�
&�ac��ȝ/V��]���(��۶�MYIb_��}J�T�;���TMG��i�����o�x��y\m��\
�q}��y��gWtmnn��<w��0:P5e������!ߩ
��zЋ�<��/�a�����_���N��9�S���~�1�\�j6Q�2[�"���@�微K�2=9����o��`�T�Ϧ[K���Ӊ{;$,\���ru���� ���g�G�٨t����Zy��V�z��\&+�����}��x�`��d�?N ��NB�s=p��g�&�����z��x�����?lϩp�MF�;O��QM�zKn|�W��� �TA��N�J�ȃ���;��T�̝��h�nw�^��Z9Gк_k�q��U%��t}����@yv/��dҘrd6���8:/�l��H��'Izpmj��ȍ�zm����O�|cz+�o�0uz������7�����ɛ�x��3��x�z0�`�����:���_��q�q�^܆�#}*GQ��	�KW��_+��Z�脮��Ɵ���;��i�4���.� ��|���'���z�S��T*����RaЬky�[{D�a;�@R׫��[����� ڮ�7�AkQZ86$tM�p,�=�{��]��f����7ك��c��/�$�t�&���q\�S�r|�h;qj��|0��(�}&���b3�}���-u�|uQwʣK�$���u�{�cx�vO
��T�E��;9�P��ʭ73������OH��}ۈk�-J�z��zO�c�|�tk���zus/�x�]*=��kBw��JJ�<vu���I�\���U}L����}�����*��]p��NI�L�x����+��Kg��>��M_�Z��d����Î��/l�a~/ǽJ��5���	���U_����Q;�Ϭi{����A�,#�q]J�%T�{�v��5��м����H��y�b6Fg���Q9�m__wzz ��X�>5��A��)zd_ǥ�9������~���t�{�a�g\v^�GNw��w�iW��t�����`����g�x���5n�,S5
I�6�<ױ=����n[;�~�8�������TIS� ����DįWp�|go�<v2Л����Y��G�G_��Q��>B��?[g#�<=�m0o��^�+�u����f�>)�jG��ѭ{k����G�WV
��gGBR�}�LoG��I���>,�|;�� �9�mf����/����ŗ��U�V�F<��RV=Jc��F��#{)Zd�N�_9�3�@u4����Fm]#�@y��9�ʆ�-��$��z�Oy}s�S(��9:Hիqq�c���^$:�	��"�[�#5%22��q�>�	5Lݼ�()/�W����q����6*zwƄ◦���k���w&-��2m�}�{�+�Q�͵���us}��Y)ҏ-J�Ӎ�/�B�EJ���oSp��1�]���܇�U��%I��+��S��>��X��.;�R*8��P.a��'tN�ߕΏv}�lx���潦�*�k��z�Z|��<_�hN�d�^��y����̘{�e{��[���t2hoN�_{w�'�D�������}.��靇�����6����_GzrM�^D�d��ÍOЪ�ifX�����ݹ��g��N��X�[���H�����Z;�6��U�k�6N���'¤�3�E�{0��n�q�f����2���F7��<�i�3��}�������Y��v�m��x_��\�����Ǽ���Ő=�e�T<X�����!���U��}^_�G��].]��UƳ_�����;�j���,�-l���,%jK '.���'���_��ۥ�^��*E۴3�.�z�D�.��y����	~;��#�?[�O.6:�$����^��o��p�V?݃r'�w)�eô�`�8�Y���~xls��/ �	a4�U�,-�j4�Nc�OP��Ei'N���wb�6>��+����B:�Tc��:��!��:S8�{����o7z�JC���8����5gf%��t�B�.��,ni��m�-��|DW5i\�+}g�GZ�R��z<���Do�#y�Dk�a�d�q {��$����(x=[���Vbz�����������'޴�9��\u�t,����4�ә�|TL�:K����t��J<H�Nm cO3��F������c>��_����&߽q�Z��Vt��SӾ�^YżUzu9�S�(q� �"�ױ9����,���{ܨ�����}�yY���{}o6g�s���z�.�i;��2|��T#�z	�������z��Y=�����׬�e���}ջ�2O�gD��n�z#���m�|{)L7z�ʍ~K �ؠ/L��J�o���D��V ��'7NkW��<�����?P�~����*�z�A�>%@���م����(B�M�U)ʗ�Z���ղ�h�>��./���s�}�ԧ=�Q=~ˡ\^L����zdEEƈo3����
,��Ee1����#z_��u��g�a?N��UD��5�c߰�o�{v*���U���vv�eCgG���x������,��T���;�ۻ޿fgd�~�R��i�Ix����\��"�"�g˪f��눒�(�	8��!A9��+�&����s����zo0L�;t���6�s��Pw��R(��"������ze�)�+x�s�Y�i�U��8�9���/	�W�9M8�g�C�z��H��f~���.3:uN�0��aE-��i�x6��R��=V�{fhd����v��k�q��}��Jg�^�;�C��Q��:n,�|���Fz��z�N�[�J6rw�wOo��HQ��	qB�Ќ�\싇����e1瞻Còn�T.ʑ�r�<k�+ƌ����"/D����`�ѽ��u'�s�Y����@�W����>>܍����=n�;"n�+�l�_)`�����n=�&lG�%,��r�0=�g�{��S�q��X��w�9R|_�H���+��f�|�O{^�k��S	%>��^�t� ox�+�rKe��]����(W���Z�q�F���������>��Y�V�z'}���ñrQ����"bK}$\A�^s���V�ւ�t���	������C�*j1u���{�>��m:��˘�3%�����1?J�u����j5��e�j�~*׋�}^!/'ldz}H�G�O|���=^��s>�Pl�$��5���T������\NfO8�k��u�}������W��"=�R���x��� �T��,�f_���ޅ�[���angI�މ]mvd�)��x�}\q>jq��k�E��el��$j�����{(*�XD�;r���;�uo@'���X‑7y�u�%߲��g(��B��&U��R�t�gC{�p�鎱�.�7f���]Vn��(,9�V�jB����vuw�z"{�E_�t�z�%>�m{n=����/��Oޠ;�]���������^����ĳp^-{����O��pzJӃk__���>7^\<��]�މ��'��1�Y��z��V��{o�{����p�x��@ɏ+����O��N����cםw��"<�ݑM<�����(�=kF����U�}=�hO{k
�O*p�Z��ઐ슏b�U��Ę�}�g�.ͻ,Ƚ{���q{G�uJ��v=�^/�hf���xW��jY;�aᯏ�C����+B�9F����J�����;�s�S T-k�#)����z�3�9���x^���Y>��x^�=�2�S�P��ɾ�j��ݻ�uϠ6G���M�ܯv�.=��J�w��hVt��ۑ���؞���I�p_�L�)�3~�.nz�8�O��I�x|�/�dz�ǹ$�U�Da�`8�%�w���ǰ�� ����>E���s㖲�7�Պ��~2<�����Ӻ���μ�gL���j���~�}��׌>�rQ�GĕFX
^�z[s�>���ǯ����T�m\��3Zw�*����:.�%~98;�p�o�c�ء���q+�y�[�:�p�q]
ox
��c"�d�9������,J�U
4�!�r��;�t��؏n��J���k;��z8Z,¸�)�M���8v	���2A���V3%�Mξ�7�v�|�F���r�rFr������}���<�=H.\��%�-3In��=+�힏�T8��z����G���w�����g�+���RM�Dm��&�̗5� ��H~X�����z=+˷����q��1���Tr~�ˏL�x�A�V�o޽�7�5d��p/'R�#���U�U���A�
�-���~�*;�W����ȟ>��>�k ���s��cW~4��d��Z�*fG�<Q٨30�)��.{Ƅ㕦���k�G��ܘm���ª\�'������y�$=p;|9@�[)Ҧ��8��� ?m͚���ϣz��j�
%�t�R��
��ܣx���������h�q�ʐj:|J�0��N�u��*��/�&��9�l��c�Ho�h����Ȇ����yF��h�/JsC=P�rU`G|�w�z��f�h�-~ �\�zl��['ND.�x�u��ȗU��οTw��G��N�n{�����Ipu��E�v��5u����}�=u�Zd�x�zϠV/;�g�=�ɷs�{#�w	)�3�D����P.w��2��ˮ�?�����C�=��'�������.�u��&I��e�5̝;�0<ŷ����Г����<�L��+�f��]l+h��,�;yw:�,E�|�.N�.��k�:A
bM����+Z@7am�=�)F�^�hw ������ݿ�J��ڎ�~Bg��+��xdA�C�p����<�/����Q��qu�/R@�w5�]�U�8��eCڙ\�l��jO���ȏI��A���V�x��$�bF.�Q��k�kc�y�w�����H{����vT�A����FU1q]T�Ӑ�*%��>���L�Dz�'��DרF�w+��x��Q��c�M��F�I@À<��`X/��i4��Q�}���f�ߺ����s�9>sپ�=�<���Tø�T��"���L��Ujr}ug���y��U��S�>��cQϫ�Q���#��s�q~#_�Dg�4���|�娛��Ϋ�>5V�����z�
��<:_��3:���H,u�l�}�޿3�O�D�ϝ<�Vz�:�w����8��#"�s' �Ǵ[�A�rs����\{�!���٦r�	OP̌_�*��gO��Q+ :��N�DҖOW�f������3���䩏R�{�5������v=y�6���c�j�Cn|O�����Ԃ�K'�����P_N��T/�
�����A1�/)��B�1wQ�k�_��@�{�z�^�KN�T�Yܜs����^o�����\M���V�
z�_w,��/�Q�)�u�R�֩�XŜ:$XgM̧tԳ�ڏuwJ뻹�v��e_Ay���ڂ��'�z����ʾ�uv��ڋVCw.��;^��Ǹ�^���y����Ҿ���}��X���T���Z��U�W��'ܷWU'!�Na��[>��y��^\,O�|rz��)Ͻ�Q=oۖ.!d�T�a�S�ۻ2��X�Z��,�
���r|3a]{��_��:�ǲ%�{LgП��_�TN�-�^��6-��'{1���|3g����3���l�wS�t_ƕ~'qu0/|�<�^�끙�Gnz�թ�_J���o�Ne6Eb+jԍ^J�Bq������|pӠ<�mxȮʎ��"��}]����ߞ�n�z���r���³���佲8�Ec���O�LN��M�Gdm�w���,�@N�B��d[�^���X�q�<;>���dn��$񯤯�{���x��^R+�b�FΙ�>�\�O��wp�w��}���o���G�ׇ���N\J��8��C�Y�f�7�|�&�3�Hݨ뮪~���S���Э�w�9R|_��H���{�'�NzI���J�f��l* �!�:[,f���������z�ў}�h����W�g)�Y�vF.��67�{�����5�:]-� ��f7Jʸܷ��68f���)*_%5�8����r�m���CI���-���+�����N�T�G����o�p'i�8F����,��ǭ��t�
�W�0۹�Ga�c=���a��9�3������g�W�;�rY�P@J����# ��9݆gB}�C�ң�C|ݵ�ۣQ[=���F�{�N;���\M�{��ǫ��,�Ȁ�}x�����7]-u���U������w�����<���p�O��Ͻ>�O� zt2n�Z��q5g�*�Cf����X[��`�}
{���Q�^���ϼ����zO��~� ;��X�rg!K'��v�7�ٌ�㱮:���q���_O�Z*�.��QH�*!�mǳ��w&�{/�Ѹ~��σ˱6CQ�+N�~����׷��ML�}�vk�9>aNu+N������y��>7�W�?Ui���Ez���5��g���Z��BW��{f��3���]2a�Z�O��N���ަ=Fu��d,�EGc�yՑ�oз�k������f�id��wL;�++�n:�t>�W�������
�����c}�F>V�:�^���Լ^G�X�9�<+=�#.�wl�<4|��{sG�;N�G�$�:��R�*6X�[�쑔�{�s�Q���sÒ��nN�\�|6��C���'�04bU�� �ݨz���=$7tn�EEnc��VYjf��r�Wge8ٍ�h�'k6�Pl������j̤uKG7�2&-���Z���83h�Iָ���f>��?,��4v�^u��G��lh��;jc�8*����(NY��+[���ۓZz�ڞ�{t�.��{��m-Z !e���A^�,a�t[}) }�$�8S�@U��!IK͜}x�=���m���(mu�\c�m\���V�;���[SN m�W��f'��R#՝����9u %<'/� Dc"�	]Hk�R�}滖q���F�(.�j�W����Z�����J��hE��lV,	�i��i����DQ��zq������ZֲX|���C�,㕮�h����t��؀��.�ԛ4�+��BD^��|���G�ݷ��_uqkD���9I�d��.69}�kEu\']�{�u�j��N���o�)ju$8�-]�&A��/.���ѩo�a�v�Z�_N�+�u�\�y�t�3{j�l� h��Y����B{�;KVAT;8��7�Z����3t��1r�U]�@��e�[�V�]����V����#Z�u���S�֡�v��`��:.�ޫ��)D�2qB�>��	K;3��eɼ♫���b�%��R�#vi��Lbܹ����}m�/����'���+�g.7��/��h2e����B����(b�c�@�	�OBsry�67o�]t��cѰ�RX��-u��o��E�=ϋ�}�>�4*	e����\����i�̜2+]7w�Z��L(Vb�4*��e�1w�ú��;b=�;�	/�nV
�q�E�:���t��Ӕx.�wr=�A���jf6�V�D��q�a;���}Ӌ���P�Rep|�u��;��+]iܲZq�²;�۝�d��f�]�x����b���
X��B��dRA90/3RLc��Ӑ]�"ԉѺ;9����
����lsFI�n��ܑ֨��?�o����ܹ�;���ř�G����:p��E[��<#ڶ=Q�#��ѐ�k�����Eۼ����p��]y�:�+���!��Ǡu�(��h^�ǯg�)8��7��\i4Խ��K�+Bv�i�ÇS���)�Xe�ܴ�j�cvg:�zwt�e�غ�n�����ެZ~en����f��؋��J�a��cEe.q�X����k.;�@�}%f��]V����9s�\x�`+-\�.��w<�N�}��v(�i]++��J-���h�f�Ѧw4X,.(��/����j��Y�v3��׋���a�Wg��D-�}���r�[
�ǹS�q�s�ٛVض	��ǖ�}u/�j��i�+d��<N;3�{$�|#:���q�~|��u�
��(�FQ�+��f�k�Aͭ��3�V�4��~˰j��'��L!.����g���C�݆Ԓ���v�����w�z��Ϟ����������"�9ę�r�&X)�����`��B��*e��9$Ns�)�H���(aD2͈Q�q"be	C#F	��@`L�0&��D"�r�H�9�"1�f0���79�
��s�a"FDf⸒i026$�8���7&I!��\q��e�9� �0A�&L�9��L�s�")s�%1�BI$�s�I��q�C�\�� �.I,Q��s#0��9�$& ���i@I��(� XB2e
Y� ��# Rh�"2o]}��}դ �Mi;P⼖I�b'%ڔ��붟/��J�����dK��#�݀�&�|�M{2ͦ��yZ���G�cg0����ߋ?��G����\2���;���6ܯv�����*�ޏe��,�Mu�b_�}�w]�rp{��$�>><=q]U阸�t%��M�z���>>Ӑ�/�W�����
�<�cر$�{{���m�>;�[����X讥s���.�Эk�����gQ�8}��G�flt�:/�;��=o���x��%GĕFX ��g��/�b};î��*��l�+�ts���
�r����V�z��g��˘}�,�ȈU�b`�\L�L���r�2���+�r�֬�G_�Tk7��+����!���#�ԇq����bi̗4��J=|����ʨ7��򴹐_M�u���j5|�GZ~�ω�>�uh/ެ�7�0Ů��P�����޻-w��dIZ|T�_�
ȥM�����!Q�j�'�>D����|O��%���������y��9�3"�|zA0��`��=�B���x�>6ר�[�;y[��]��ΘìfM.�p��d���p911{��2M"���d���O��K�/�y��L��~�s���V$�4�>к��o�Չh�V���*��w�)7k�,�#ʌB]���v�uد5��K�Z�H֣[�}���F�قa��YH�gL�X^�v-��,�=�:���v�6�a]�/aR��5��8�Z-��7̋��
6�̥�����^wt/�zg�> ��㽕 �O�U2a����[���ye߳e���o��{��k�4^�������x��Չ���M�̋ȍ�N���^.�xLxf�	tj*�1�L)��m�p�ռn�^��q~/:��3���~��9�;���ܽ�zrNN���t�^���Y�.�s�W(�w�P=��jB[�L����{>�K���G�sǲ=�p��� �
�yh>��h߲�
�tz<��ۉ��3�OO���N���� �᾿p�/z�u^�#B��y�v>�<9�q�C��jʇ�"W���'�P
|\dFDy����2�w��]�5;6��V<�WR�o3��;~�G�ï��~+#�H{��1�v�\eC�N���~/��G����G���ng$�{O��Gw%������	��d{���}�G���zM�%E�UA�p7����laNd���X�/FONq~}w�~�u�\O��NG��9��P���TF�:����+TK�"�}�[���v���� �}' ��oR�K�o��"��\UϽi�s9����4���둱��QI~�c�B]��4L6�s�uj?��ݛ�\�9��r�]�c�J3�wT���f#���V�3���vd��Q��}Iz�ź��{J�"�������>̒�.WB�3��p.�<�k�(QZ/�\�}�U/p�
����su`�=�Qs^�j�\�?��x*��?�}DL�\q~,b�gQ�ʐX��ٌ��_�o��P��Z\ͮ];��_�jzS2%��50��:��+�h\Rt�{a���ǹY����6��}9»��ѣޟzώ|};�^@�F@�t�&��z�0�b{W�/��o謖�m��UJ��ףq����}����+���>���b���~ːj!K'������Q����^�Xrg����^�^�>�s�z�z�񶽷��:�7���߯�q�@yV;�2��Ĭ�sһ|bnx�\e�{Y�z�#㒮�lc�;���
����L������{��z�~ܰ�n�)u(�>�v�NWrž33��t�䠮·qY^p���#z_��Z��}潦3��]���|�T�ϵn\��fWi���D��?�_�Ḅ���|?T@�����~'qu0*/|�<���^��f&&nv�7�p�^�}�\�����ug�\ΝE��pfT	�,\Rھ9��7LAjq궍g�q���֙��ׯ��޺~*\��z����A佥��'� �%/8�Q�;���Q4�fi��R�I�D��X�����'��)�N��imy�,{�t�S���S��G��?L+��/�TqR��,���mv���a�r}YYnc���3�Ʒc���+8�M�$�!W�8�m����J��st�U�%d�K�-���pC6ﺧ�n��}�!�^����Ly�޻Cò"n�.�����$�^@�*����nWO��>���m�MzL�`���wz��#�'�۟o�����u����pW�<b�؏���,މ���u��'}����`5Q������חS�q��X��'~��O����<z��~�N��zR������A���9��`L+�nKe��]���z�HU��hh��戫��\�\2�s�z�oO�Dw�iW��\N�e�}�J	TQ%��,��9݆gBW���"����f���hC���c#�Nu�v��R�n#=�����d�H��@�&&%z����!{7$�;����ı������k����8Z~v�}��"}�ӡ�p���/�뉨s>�V���WB��<U��Wd�������=����t�=iT?r�M_�߽�@�=> o���Pꜙ�꜠vj�^�L��sp�'�D��3�7N
�]Z*�˥��q)|m�mǱ��ɷ��M��P����fzC]�nkn��g�y��&�=0ʚ9,u�=8�JӢ�__��F�>7�W���4�X���׮��݄r�-�"7�J��w��Vh���8���9�l����4��n��	��ՠ�#��㶺�V��s%�k�;��_.˷a}��vC���F@�t�+�-�}�9A��(��S�l��aլ�i�W�Y�련��I�CKJ@�ܕǯ�I�P��w�n8����W@Ɇ�mhwS�:/�N����c��;�>I�TVlWO����Οdk����V%lؑ�ꇥ6�+�N7�����Q�Y0�V-��2^VE�f�9N��o��*/Z��U�����W���>���)d��|fu��+�-a��}�����^����pjS%`���k^�NW�'#�Q���7H,�mp�Μ����N��J�a�6�R�:\c��T�'� Ft˩/�}ʂ��w}^&�nW��}��y��\w{�m���7zy#������I'��=P&x9�L��[�.nz�<�ޯ~�>>��X��$�Y�����磭�{��7��(� �,E��U>.�Qfzy���y�=�������w�o��� �G�uṾ������x��%GĕPe� ��g��;Y��=�p}���Է�;�5��p�j��Fy�y��ޡ�\g��˘qD��ʾ3t(�q�Y]��vO���b���*R/v��ny\U����NW���C��zH���LM9���θO���fȺ;����%2%�k#��B5ߧ���m�K������ڦ�站6%V4�&R{V↵�P�[���v��AЧt��{%^��@m��q>ٖ,������n��)������P�����wK�0B���h�^Y+�f}j��F,��թx�|vH���`�å#��j5|�G_���>&��şuh6���2��oMWۇ=#١n�R�,ϣ�$�7�L��"e�����M����!Q�j�%G�>D��Z@c53�^��#��$������T�H?��:�J����å忋X�q����k�G��fwZ�t��ؠ�ѻ���'���{!������d�=�@ɇ�'�b�Z�ѕ���泙G3���״������]����wB��zf�������E��eH<|J�0�����Z����^��>a�z޿�G��r�k�xhyח��W���P�����dЯ��R2�Y:��5����=��2��zF#�*�VSF�O��8�_��Z��}��~�֧�/]A��r���^;�Uy�:����^�N��I�9�����Uix�zK�_-��DK���}F�w8?d�L�ŏo����xI�O�oz-{ռ_�z��߉�yIx[�	h�O_�t_�����>����`r��F_�w]o��w�:;Ί�t�Vz��v:�b�;*t�E�O�,^D<X���I���A�5�!A�ў�/�c?�RQ5��z�3�`�2�S���@� �o�$m4mVE���7ok�Ȕh%��h��MJ[ �Z�r0Z>��e:Pc��iv��R�aK���~yn����l�uw�:��C6�J51uL��8��ѣ�Ve�� �bR
E����	�P�D�`�������Vz�v�0��Q�,��a�ѕLI��Lt�h��ץ�d/T���*%ڷ�!��{ף��q���u�[�s�_��H�J{sGu��_�eQ:�n��V���x�Tl���P��'��~늸�;����=����I�S�v` �b�n^ٯw������j$�!z||:[/\��T;򸫟z�9��\v�iS�z�	��.���v��Z�q��zk���dT ���1�p6:_��3:���H'>��kqs�#��w379A��B��n�|}=��'냷�d�7���A�hJr�u�3���9�	����ᝪ-SQs����gޟ+>8};�^G��˘�Y;���b��z�>��2EeE��f�*���_V��7���'dx\?+�ۯ��z|{>f� ���K'� �թ3�^��4�E�j�)U����=պsn_�Vo\{��^������?P�~���U��̂����V��~x2���Y/�F�����w�l�>Gb9K�yח	?Ui_>��S��ʉ����ȏ�U�:���v��<��{��y���w'�[Ce>�W`[���#��u�i��/P{ %N�N�oj�o~�XS�
*Ju�c��5�%}�	�J;;oV�#�����Ƅq�K��-E�T�� �Ji$M�QԓE�������W��#+�n����y3�>�䰮·9>�^��}�/��\{"\״�m�>q1յ"S��WE�S^�=Ϊ'M���>fp�㓛3���·'$��4��;�.�v�"&�����1�����uM炱����D��y�05z��N�J�S��|�Kj��/@���y�@z���o7���/<0*�^22������Y���xW��S��'�vZ���W5Wy��v2����j��v�M���oz�Cφ��E��^��ǲ���R��B��=xK�ͣ��י&Ϥ����u�MzM�t�n;�qޟa_{���r7��r=n�;�F��j�^S@mx�q]n��6N�t�z�|�*�q]T��k˩����UǓ�q�'���� �V�,��K2�����՘����ߋ��F�<��'�x���l����#��B�$V�Ҝc������T���ln��ys�#��U�}q;q�a�ʀC�C���I��vjc6X�.3N�a^�Ѿb��v���;c���5G�K���޸<n#�ꉨfK( މ�c>�c�2��ߚ s$�_�`�uύ�����g<m��>��P��B�˚�b��H9�J��ji����뺭��QRuuϊM�t��ʏݜZ=�y�w� �gP��2�d�H.�O{O}��xq�ERR�h]pg�ͯ!��/�,�'�%���n����׆��N@p�O�����|�zt2n�Z���g�*�;j��<�/@��O�����a �.������P�T?1Q��j�'���|�� ;��u�d_�����>՝�t�g���3�l��_K��Wt�z�%/�^ʏ(j���~&��dG�yӐe侁W�]¼�=�b���(Ǌ����Ӂ�Zpmk���z_U�(����[N����k5%F�S�1�|�&���=q׶o����>%T@Ɇ��Z�i�)Γ��z��d��6~9R+��N��X�Do��1�7^쌍~�ޗ��V%_�X(R�T�,n٘^�9��*f�yߘܲ=>��zl�:@�.� ���{�;�R�yucx�d��\ȴY9�Q�'�̩�xXzx�J\���2�ӓ:vO�+ m0ֽr9^���]F{�"<� �mpDOިc�T/xa���7�Do����qW�S�H��nT.4���M�R��S����������z��]�ތ�G�ب���:/�RI�P�|&x;��L�S�.y���χz���C�(z4N\�ô⨣#���� �;�^��\���-.����բ�w@��=I��s7_�Q`��{f�oB�w&�͞�����9+�'A5���ٷ,�LgK�igu�j��㳳PB��;u+�,qc��!�
��t��.̼�[ѹ�iE�����/�g��{��7��(�E� �|e�0�bzV��(���D+Y���_����v�o��wZ1��cr#}Cǟ�G�A��p.J5����2����@��Dc�Zr�7��/���ym�*����%����z��FG�W�[�VzP8\����f�<�+)\{0a�����o8cŪ�o⧼}�F�p���}�x��Oԇq����bp_��D�L⽏mr9�w^k�z}� {4T�2�\��h�v��o��Tu�~��G�s��t��AmX�g�n�{{�ܯwj��h�6���R:j3pzH�~�*�SG� _��!Q�j�&n�r���^�y�'o��w����Ө��3X9�3"�g���/\X=�Ck.7�S�~�b�P7B�^�.�V�¯�_��ܘ��~�&����D3Q���2J�ѓ��>�-m�3�ރ��G��Օr��V^���i�r���j�����~���ޟ z���;�2���a��d�X�>^�렒�]Tޘ^����}s�>[�Å�^_�s>Ҿ}�4��x'��&�z�D� ��X���][b%���R�q�����+tXɮ�5yE],Gb��S.�j�M�#��t�Zye��Vr!��}��3\��\
�uN�9��)�'H���[�]r:�[˵0;�0�^�=�TB�V�����_Y�G%^��Ng�kzΜ�;��(M]��.�JA�y&V�wUnW�Ñ�w�1��XUȜމ��Ԏ0��x�6���7�뫧u�Ҭ�����i;QK�o&��\�m��4w$��Df�����.�,�&�k�^���g C�[#�ti���o7!�藓gA����Rдɥ]u裥����Pw+���̜Uw�c��V�-���ö�����WY	Yo3�,�HF�r�j��[`<�ݶ��8�d��v	2Ȅ�[�C�	6,!��#5�br�cI�����"���o[č���͇��BH��µ���(��p�Sx.�k�m�Y�wa���:`�Z,�eb���c�"�4_˫D�^���h���x�
���,����� ��Ҙ����C,o_�`q'���P�|]�:�b;�HW�;����,�;�.!�[���Q�`�F	���ﭹt��<��XΈ�<z�`B젘1��Ս������\��n[���ڳ���`��V#S@��6Q����ʇj�h��0��$hS�CTv�r���lr��#�H��L|v�Ջ.3����;�7��&:w�n)\��TSu�l\��&m-��r�RYo��T��_Y,h�U!�Tg%0k�!-G5^f�aWN�ހ^�}O������nJ�osv:l���Ш�t2��,\BݎC'�(֚�G^���˚;��d�&G5�һw�1�����R��:�U�����3:(в��uGDo��{�T]�3X2�ƶ�c#0wP�W4���agvP�l�ɾB�x��F��N�Ws	���`e�p]!"z\�,d�)
�`#�b��A^=��i>���ͣ0�N����P�S���x$0����һ��6�)+�\�nX�[���)�۾Aq���p���(�u+����%]�$��M��:�H�ձ���/	�"��F�7���v"�q��U���j����k�$�g]�TH;|�w���v���5��*|�]3AFn�igu��2*�L�.�[�ݘ*���@fc��]��u�������3s���E����6��;�#MR��MփV�����[��y{�1�rT�'7�)ɼܼ#5Ul���"�����Q,������Kn8�mK�f�M`\Pcje%g/6��_]r�8����H�j��ϲ����TL�u�BG����RÈsC(���mL�ط�/a�@��b0�b�b��-4d���2;��wp�M^)y9@�"Ƨ2���y�{�M�۹���{�84r��p�p���$��!2m��F�	وz랹��:�e"($�6=7	%	�d�L4�0)C�-	"��T&��!)A�H�)��+��4�\\���ID��MJ4̋�䑅����HL�`�`��24�$,&bF�QLP̓D��h�i1��)2�RR��!$���KF2���d�-A�$)	1��F)����)�4h�J!�$�L�b#bfeDXH�Li�F
R,lF13@�(Rh�DP�BTL�c	��L�	�Q��H�0�%��
0�Ad�i&Ē`��b�fX�%2c�E��_z���~���}�8�J��94�*�9_y�z�΢8!]W��놃TJ��Rf5����l��A�9��dۦ��dV��-]���A#pwj�W���S�'ND.��J���9�?Tw����PwK]vF����W��H��Y���󜓗���A��wYU��W�GˁK|�=�.���Q3N�򽦫���DF�'c���^�ړ�s�.����+�#�%%�l%����Ti��;>ߓ��y�#/:��{�Wv.��߬G��>�/Ǘ��\w9�c�6��>�����^�i��[���k�h-��I��;D�ni�^Qg����XY5ׁG��_������3|au̢ǉ9�U{�楰��+w���i�ܱw�z"��gӏ2�};yb/z�/p�x�G���[���9s�_�.J;޹�㮋�����Ա�O{�1�$��+����]���z��q�~Ӟr|�7��q�TF���c/ ځ����W.�pp(��S_I���6:[/5ՍEוE(�z�9��s�q�~�-����]���þ���k3�;diA��"�[���/ō�g�|���)��\��\��^����zu߼v���~����W���2Z����q�A�h(�N��Kp$�|��;�#ş�;�}��9��i:I��-urò��*�MM�l��;����Έº]�Ύ#�{Q��De��Q�2��ym���������j�).S�r�WJ�)�|��n-m�������2`3��,�{�,G%voF�VNZL�څ�����Z��[3�b�-IF��n��m_�>T|_��~K�@�a�:������Y(l�����2.�;ܢ{�r�Q�ԧ��y	S�tG���w"�u�}>|���)�.A�R���z-�껌@NG�:��`\|s**}��9�/ǫ7�k�~�:�7������d�bN��Q��O�$sn�k�r�:N���l��r�p�V���w��7ח��}�ԧ�,�-+ӊs;}
��w��z%���b�y3��t�F�gC���U/�Ӛ_���WX(��zb�;��U��֘�Ӭ�}�wߦ��3���p����χꁳ��T�iW�w�,K�k2gЀ�n���}�چ� �c�Ù^��g��bI�
��-�p�دy���3*�~.��.lk���U�]�XD쀻�6�}K�B��~=t�VS�;�=��S���,�%�"����ճ�&�>���]�,��Tz�)��7��<�w��<�Y�W�=��c�#�]��Ƨ��}���m�W��ʴ�i_�g���N���j��]tפ�t�Y���@�W�������T?t��Lg9��1�+�fs�Wj˘&)���EGq�Yn�����MH�~�8�&6�`�WL�����H͊�7�;*�q�u��U��Ҋǭ�;x1�B��Ou2j��2G`[H	���g�������co��A�vY��R��!N9��Ғ�*z/6T&��k�4�wwFd��7�7Hz�S�I�`G��Ȋ���a���߯�b��{O�u�Y���`��5}�B][ㇰ�7�<z�1���f�w��B��,�)^3p:[,f���L5�X.�R���'}����cFG�z�=�0����v��S0�\�T ؃�"bK}$b�F߹�����^�+-V����z�C"'�v�}����z�y�\7�TK�������o�pb�b�JG��k�w�1��YF�{����5���?;c�҉�����ՠ_��|T�!k"��Gm���ܦ_�C�eI���Q�R���J���y1Q֚�I���HdW����:u��8uﻮ�3�g�|ꜙ���� ����/�E_їKǨ�^��^ۏc󻓳�D��-ԇ�;t��,C�d��/:��b��>ɒ�2�~9,u�N%i��V��ޗ�Z����Y�n��C�aYֆfz3�n�k�O���τ��^���3gx��P2a�Z�T�N�|�^uԡgP��[�o-��~�o��g]����vFk����*�*�6�P�쇥6�+�	��yI��k�O��<��|"��Z�_<��P�w�G4�Zkq�ݙS���c�	�M���)�s�����p�������ʭT�r5� y�%�6�۴:��}�h��(*�=2:�6��������*臸�´�6�-�R��sR{�P\t`PW;������)����ռn�փ����:�_:�^�οR�y�V;�vO
��T�y��pG��(zE�y���P�^
�H�ZlԿ�� V&��%��I~��}9��.��fO��UV��xF��l۫�Լn]�J>@���u-���^�����x���0��.8xmǯ�%b�p���Tn�塜nN��rI�C�g�����3��K�}����Tzs��mxґj���;=`�΋>ӏ��Vz�ǻ>3|i�(�$ߌ�$"��u+�CP�9G��.��7�E�ϣ�U��I߇�G��ȍ��~w�3~0��F��%W�X�H�|��X��/wX�ɐ8�9�Ϯ�}���ާ�ё���V��iY�@��t����wv|5K.o)�����mx@]�1�oJ'>=/���F�o��*����!�s�u|�Hq9�I^OG�3�W�7Z6�Ӻ��}�}��J�� �>�&[��t�}��j/���O��Ͻ3�}㾤Y�IC��#1�ٟrմ����>��fv�-5-�=$O��HT�h����G�
�v#|_��L��>[�[��	���dy�KgP�\qh�Q�u�N�$2Tg1��4+�����G����p�n��(�f�K6CX[�p(����ug�2jy+�;3���uge�	ø�$i�:�F�u��
v�}tS���w��1���W38����[ѷ�d*Jl��v��ѻ���x�����f�
snfE"�M�^�
�TD��X�q�p�j�\ǔӊ�&�r}����=~����7��>���f�*:}�IA��2a�������2}X�mg��X�W:|oz|5�U�7���=3~���w����������7��ugPnz��O����¸�[���/���+��W^�U�9��P���<o�4��M��&ړ}\�Kf}"��N��#gv��Օ�D���Z_�ε~.���~��9Q��c�� �5g���`w�*�py�h�%9'/���C��N�u�\n*ex�p�|�=��c��;��Sו�C=Э/\�r��#v�ؼQK�3�פ���e��x,����i��^���<���pҡ����Β�b��g�>�r�|�S=�v�;�b1Y�S��'�-|�b�Y]G���1ѵ�-��r{�'�}A��9Շ��x�z|1D?S�Y����\aṃA�vy��F`�T�^�(�w���3���+��.qfTO���>޽��O�w} {_���s�o������߿�o�CB%�U8
��\R���W*�����`r��(�*�(�zN��U�d��u�Xy;ZVt���wj�Bp��k��fe�U$ܓ͜ɭ¶����W6�5�vr|Й�'��ܬ��R*�
�[�л$�Z�zR�yF�&>�)Y�F�k6:r�,i'�f	��Q��l�}w�q��\Q�a�9>sپ����9;/��t��Vj�Z�gw��Dz�G�Q/�<���$7^�Ke溱����Wq� ���٪�ݯZ���*+��#J����,ι�Y�����Q-�|e�����'-��;���f���&��{ԯ��}�޿3���M�z��Ǫ�dS�-H���"d�)����D�,��=yݞ������r�:���1����Ӿ%��F@��:��R��3ô�5�H��bL߽|sY�k9g��;��}Y<�o!*c����~Wr.!�^'�=>���`�rߝeǞC���jw�-�d�j�"_���!\�D��ӑ�+ǫ7�����)�>����p�~���.W�����魻ŕ��沤���@�|n�>�ñ���+l��R+&�n��-X�BB�>��#*�=Rs��a�F�]>���z�=���g.:|
5rXV6t;��U/�����E{����Q�1U�x�j�w�\�����^Ǖ�O_߫4�?��(x����~�:<~�Z����B{�_�7�������"�ߕ��wV��7������M�l�1�ǐ���NU���i]^��r�)5L��m��j�ww+2`GH�!����]�_BF&Mb�{97�X^�P�9�:�b�oA��J��ܠ+k��8�^v�a��*�f�ssA�ѭ�CRf�v�D߷����k#�̯_��N��~���m/�q�� �^_�]\ԕ�?Zk���Ǿ�ɭ"\��d����ׯ��޺~+>�Hw{<+���3�ກ����{7S�I/���.��Es��}~�χz�C����e{�޹c��\��Ԅx��'r�t;�#��ڇ92�IbG����F<y�B���>wp�w��r=�|}�t\�ĥ��v�dW��qWz��:�1�u�X6JE�Ol�G�C����a���߯�b��z{j�L9ؚ��,�׶_�ӌ�w��p�e�6
4���Pe���-�3<�l��Ǎ��N�o`�;>V�
��z�ў}�h�w�iW�\Nߪ����|������������h��.|�H�������O�Hp_D������_�l{Ը�����W�&���r���Uz:/�����K�j�&�tr+�#��j5�>XG������>�����V��R�Uw����%��e�v��++�>�L���d6l��1��F��-�����1Q֚�I���R�~<}	�(�̻F�}[�^I�\���x�,8�S�u��0˶�[�Oh�Z歮:�1�d���*�J�v��剼�#��s���w�#�B��e"��7��)�ܹZ�\�&ڝJ�[�]9�̡��;�X������u16p�D��.�:��^7v��@:��ȧ��:���<�:^ׁˏ���K�ײ�Ů>ي���y�J]���l�Gz}�h�{ޠ;�]����dҘeM�:<l=�Zt\V��#������Pnz'=��j�zq��?7�1���7�	���7�q��||J��_�kC���a���k��g:�֢Oj�o���Q;������w���}��#\��B{ѵ��D/eN��|�c��g��J��v{�����0���|d�t�]~ W׾w��{�;��/�uc��d�k"���nf��Z�ՙ|5.5��N��A��5ʣ�YU��Կ�� V&��%��Iq���f��^17Ys�����+����~��^���E���Iz�+]t���F}�z�����>�9+69�K���s{Գ���tWz;.������]!�Ӓt]�$�L��3��WUzf.#�З%����y�%�L����ݔ��Bo�3�u o�|}���~�q��7Ƒ�2�ےT`L@>E��wY:;�N�P�^�
}:}�R���Պ���о�G����zߝǸ��䢇�*i�Y��+C�LOe��Fw×���;G�Y�]��j�<W.�ĺ~�ۿabB^8���߷Z{�P��U�:��sm�C¦h�S��Y}��̾�ƴO�3f�JV^e]0�4A��Z�g� :�Cn��u�B����;����cS̧.
3eEp��o%QY���k|���� i֧���'���p�z��FG�W�[ޡ�_��@�N����Ȩr��Y��+����5Q�@/O��x���5}�qW���Ͻ9^G����}w�ǣ<�O���{ۋV�x����M|�J��@��"�[��t�}��3Q��C�*:�?[e������,g����Lw����A�V�p��@�M��$����Q�����B��4xr��nX�����*7���]B�y�r}��O���w��!���3#g������X+�s�4J��Ɍ�}�J�贈����M���{���#���������7�O�w���z�YD����uе^�w{W���P�����4���ǧ�oFV����c���1�����L������.;�R�=�.�r����<y�[�%�����׫t�ԥ����~/�μ��<����x�q��b���z����^z=O�z��ʑ�,��ax�Ɇ�+�٩zN����s�W�s>�3�{�{s]24`�^��(�z�x��Lr.��6kӪ���V�B�N��zZ*#���P
߁���R{�sb��j����2q�GG'rG<7����Ic$f�k��+��
��G_w�v����(I��-�ܱ�pr�=(��+v�u�ot����m �*�umt2ȃ ��p]�1��+�d���꘹��O�)���5(U�/��B��3�d�����҃g�z�<{�u��<�c�KW~GJK���t���:�q>C�&)�o#�.������R�W�߁�n�����׼VC�q��ю���A���c)�9�L��>�ޣ|�����mVɾ�Pe��Xy}^[���܇�~+=t����]�(�edO6���{|�[�+3[^d�3��p�����Y�����{ՁG�O�w#}@{����w���@����~GT������Q�ĕFc�$�T;���Q>+���i�'�wl5^d��vڜ[׫-��q�#�
�@��%�0�����]X�r�\Q����W�ە�F��4����ad���{�{}r6�4�ә� "�}DL�\������#!�wG�,]ݟF��!׭��޿3���M�z�����E9����n�u����x��yǻ��TОs��������W��z|���N�����DҖ:b"Jk����o�7��ދ�7F�N��J]7�T7ʈc�:�*T�x�:�ޏ�ն�m��Vڵ��ͫmZ��Vڵ�歵km�5m�[o�ն�m���mZ��[j���ڶխ��5m�[o���V���mZ�~ն�m��mZ�{�m�[o�ն�m�ƭ�km���խ����V���Vڵ��n��km�Vڵ����
�2���@��R��������>�����V�âB� R�
	Q@ 
�g �m�PU%@�
�TP��R��$�.8�R�R@�AJJUUER" P��F��X1�X5�jX��[l�dM5h�q��aJ�j�AU\��  �  ݍ�A�m�qn]t�jfćj��j�Zi�٫5$i���UU3h����J-�)�kL�lK� 5��UWl��6%.ZR�b�k"5����l[Pv܅�#N�]�ՕEm�3�ls�F����]&�lu��劗g85S�GU��N�5��s
UQ��YV��iV�T3f�E���)Ad�,��v�m����3M��2�QEf�Q�X!�jm��١���*D���Uk6�#&UW c�ClěP��bdk!I$͚�      T���ҩT@ 4     ��0�%T�       �&MLL`���y��R����M2d�` sLL�4a0LM0	�C`F&�J #$��D�ɚ�Q�M�6ԟO�����^q��Vs���a�W�������G� B��4� !	 ~0�$�,����/�%�HC2A��'������?��v����3$$$ ��BB��1"H)	$$��VBBm!�������@�������?��@���$��
��������*?rJ�\���?�'����&�
�����O����x�r�b�ַ��h�8��ky��&�����]ٻXؐ;�@k���24:KUї�RŰr��ݰ�PV��츎%6�2�-��nʗ�٠�5KKm-��ZU���C��"�fCv�TZ�]}��U�ՍNퟝr�U�$��)�Ť�L�L�@*˖��zi��Y���e������X2��m�I*:�]�)4i�gr�XF�j�r��|ܼg�lm�����T��pne���z�ްz�J�/4勴7B��7.�2i�t,�4Y�G.�ؽ��Z�V�Yu�-�g�^j�Us�����++,,�ܕx.G@:��N�ޫ�+��M�ڽҬ�;y���~�@0�7s�������>��=й��qj�*M��Dr3ޔ*�N�#�V:��,�i�u�څ3]ku��R�ea�6P�Ɉ�̭�mb�F
���h��
Ѭ�f�Y5+Wwx�k*��4�*X�F�)��K4SpVhT��f1�]��a���m�a,Uࠐ��w3)n���k�ޱ�U�7�����ͨ�n��U�ʻչ�LՊ�m�tŜQ�K%�`�Yf�����6�٫[�bVl:!�㥉ր��rLL3F�Պ*���� ;��"�h�P56�RӦ�G�h�r��K���a������rVP��X���� ���׌Q�֛�Jҧ��k'�sT�x���V�j��:p����j�;j�T�pm)W�����c83�i�x���a�k���j+�����̖7mJXRy{F�^]Ҭ�n�ڱ�6��]`vX�%��2��sm�`/��rd�zl�ܽ�G$�1�p�/7pY;�V�5qGi^VS��e���A$����:�l�kq|�-%�ʳwu�X��6HO�(�V��c��F��N�:9ZlK��clA��U
��;M}vr21�N�Q���j�3�I�XB��.䍥�t`�.�3Nnm�RV7��z�2��U�&��@7X��l�q*�.���M6�j�=����aX��l��[2M"+�����sv�^m;t��ˌ�.P�v
o%
%�o��i�{1�@=����,�p��B�jՓ7QgK�c��V72��/bѪ3u��b��A+-e �l�3u0ۛef��2]�C��N���,S6Y0�jm���4���os��U�K�i��ũU���Y#ܠ��{@ꖌ��e��8r��'{��]eZR��x�{�m^�0�B�Y��&H�*�'eZ3j7$fstP�x��m����m"���x��;b�N�h�xT�g4��`8;��x�-ޜ��p0�Tx]�]t�:�$����u˹H���#����bƒ^�&icr�fv
˫c�i��t�o���YcP�QRfkW��*e�W���႘��f��Kƭa���Y�)j�%S�l���"#a�K�i��.hb l�v(w[`
��Z��Γ�R��
WXjv��e1��[�y��R�����7#o~�W�j*�R�\4�^+&7��Uw�n�P
}���x��:eX�.݅B���KD��hbŊl��B�M�e�3�pkd*KtU�f��n]��m6�Җ���Edڄ�(M�cZ����I3b��d�LJ�/2Ꜥ���t^XI'c)`�+6Z�z�U�Ɂ)ڍV�st�cR��nb���J�[�)Y
�D9�aȲLu�{���;h
���0�kl哠^՚v�k!�C[o)������h^Rm�"++tJ�6�9��ov�ݕy0�R��l�+�9��iLn1"Ea�X�I��,��f$�E��f,��"�ܑ��P���M�KBM`����YA*%S_K�ˊ��b�sSI��#�ʴ5;��{i������h���ӛP8W-���gm��V,_Z
�'Z�Y�7kj�Z�嗬X�'�
ѡlӖUa�:�*T�Fᣅ^Г-m�Kr4oC�B�c5�#�HT��ū�ۺ�ӵ�Y�	}��o+SO�x�
嗛kv���8/��	Y*�V\���0�av%YM�'e]s���۱w|f�����"݊]�?�'׋Ub[`-�����gz��š�{�j�Sོ�������E�cS������m�S4�K�@;{e]�WSM��7�z�^�+�E�a�TG(+����.˲�,\`��jD�!L��+d�t����@q	��*_W�������P���3������1_c�c��7���!��w�w���A7U��~�Y�Gpl�Ͽ[�1���{ހ                                                                 �                                                                                                              ]�]	qc(݄O,_���r���=��)z[L�Y�pf[a��f���l�N���,@�X�ԵQ��Y��}�x�G��9�T�hL�����9f��P'Q�.խͺ�����] f�Q�|7
C�\.�����V��y.��#q�q�-ǚ��o!�)ݙ���Ex6�����
�	գ[ʥ։�n78�G�}�C\}h&*��%L�P�%��cj�S�{fs�V�@�}�շ�eγ஍����6�\Z��׳{tV��t�dֹ�gJeF�$ef�-�v�n�r��b�������QQ���N�yX깉�כ������Ʒ[n4���%U��-8U�J�gN���M�0�zp��;�Upnu:�l��<�8աP[RV��U�Z>�p^��ee�`ۦB�4��³���{��4��wU�(S��`[O[�:��x-Ψ69��'�&���$U��.�#��x����Z��ƛ����eãF`��M����� ���te2&Y��)��(��=Q.��Âu
�Lr�!�Ё��T  [�n�4D��Ҳ�m=��җ+x�ɹ"T��$S��'�����/����7�����t�u&���3�S�u�3c�v4�xKq6�=�q�J��#K!�3��QQ�|8:��u�5l��A�&_#�&����Oz��t�fi<qɜHO��Ч-�V]�
�h3N^'.{�%�ST��ɦ@��Qٮ�u�/vM�����!��(g���^�(�T<�s���2rf�Ρ��V̒BU����,=K�s��=B41>�+".�mhcm�|�z��<����u�����L�L�%X�8=zZ[W��s�E�9*�
<7gEYG;�$U�\iJ������3 ��2�m	e)������˜�NńU��"�Ó�
E��hئ�m4�\��}�WQ�w�z�^3�wf�h�iB�:>���L�����uL���2���[��L�jbJ=�u1�U3�˪�@�Ʃɉ�
Nc�
��␹M֭z�βΝ�j���ŏD�!��0�}Զ S�p��1��4r9mq�S����wCX��|mv�I�͋�aXR<-L7fʵܻ�"�u[]G"�N��L���sT��B;N������"]�g	��뎰��W�O�i���.)�5Y�;����������$�J�͘ơ��<ғ��V�MP�CL�l�S@e�E���'�j�!�c$�Bvb >�Y���l�2Y@\�3B���-ת�[h��ru��)4\�9R�� �\��鞻��.������7��QQ!e�9H���cF�W�qC�VmO�S��7���1��������|̓n� �c�RV�ǭ��wJ;��3��	oV�Y�+��aIp���NŬp�`��h4�v�B�(����O� 4T#��_Voޢ�"��f��B�ΧDu�h�q��;w����#m�T�6Z�4R���K��쬗4^ֳ�Ms���j�nm�n,OM�:n����Wd���/C�u����)&��>�:���K�`��Y�O��
�D��A�kd�����V]X��vP�yw��AZf�p��ƨu��3��*�_*f	�N�jV�o.e-�B�v�j
eiu������vݞ�z�M�v���SF�>�Kat��>��Έ�����������3;/7�DU���8돧��f�5j�+7
�%�c^��55��%I��c��JnK���t�ʅ1���<>����g;G0+�W�"�u�(>�U�1� �V�iI�Hܭ�/6���Aw1S�sK�n����:�i�ߵW]a�i���o3���&��&GM��� � Ĉ�_��v�&���T���0�{.c�zL���r�6��fɔ�E������˦��V�ݺk�)׷�¾�����c7]�
"(��/��9+YH�7A��$��-4!������Bͧ�佊(z,�-��f����3pQ3v�b�=��a8��E�'u�}���% ��/��d��]9D
�W�~�0#��+2ɠ�v��d#�Y!�T�Â/�7J=���#¬�
�K:K�r(�h�zz���ySjƫ��Lʒ�c��޼��*v��!MHӫ�qa�@z�7x�Y|� w��{����{�����?fg����o��k��՗� B�	x�d �$>���~�w�4QG�$�$����?�gM����)�c��ٕ�Y��{�	�r=�ۼ�h�4�Ҏ_*Z�%��k0S��w��v�+h�1\���5��7"����Ș�[�ͱW�JVnP%Q�X��'����8�d�)%N���`��[�@L�˵]}t<�����JA!2��C� ����F,Պ]�r�X$X����C����V\,rφuЅ���2���#�N/.L㏖d�/%o�uyx&�x�i�틬8�2�+e.iv�J�>kl�����c�������yZ��TsGj[���M*���we�C4ە{X��']�9���n�Ct��i��U�Y��
P�t��R� :��c6�]���}c,R<��(�V�%- �(S9tG�����/K�O��v���Xk@��* ��h��Q2[D���cn�´M������]\u ,��y}���
P=��++�!�n�/��SKLGj����a���k@����k�ץ;�4�%�փ�U�E^�M�p�vj�p���M��Yo5�e�aZ�=���)7e�jE�YD�E���%�Ѭp�5�v]�f,���`�틺��МL5�1U�'a�wA�r����S.�npB�Pμ�1t37i�k���V���U7x��7Y�x�@����M+�6�[Ё�e�W����n2�b�7R������5��)eYYIξ�7Vi��AÒ�b�wr������c�@@ٔ) _�/�:�{D���K��.�_-?^�QR��Oe3������RJc9�������}�=5u�ݲi��kwm\c�]�[�;F�5�
b��t��g!�����{������v����J�]�ۛ��ڻ�n�+��X�4���0֟�G���N�G%;Dyt��v�m�V-Pe`�7�Pb�AY���s+�;�nm�����ln�`MD޼�	�Օ��'k���j�\�Kw���y���ܭ*��{xf�U�YzRh+��M18�����|nV> �Up��������w���/j໡�D
�9X��O�J��> |r���
YZ��}p�/�bԆ�A��f�<�f���p�p�i[��LݻHٴ���ϒ����u,�zb6�wcw6�N��c��m����R,�:�7J��d�F����x��*���.l�t��ם��Wt�04T ��a;[�j*�a60������҆m�ɱtLC��]�F������x��wt]�m�w��p�b��u,ؒ��g(�[���L+\�f���Z��;��F���y'-�� �nv|JۦQs�ŝW�E;*�����a
�7 r�#h�m2eK-�I�ڋ�	��ך�mL�˄sJ����s���]
YQ�u-_^���ެ�~��P-Q�$�v^J�[�Iu�6.�4;��&o�+�^�a��3���U�76�S��
�� e�j��I����X�@*�|I!r��7Nl�-�Hµu�[+�݋7����h�/��8a�sh#B�cW�J�ij�Y|%��^;��ߊtmW���J�AK�mu�ɡW���7��{���`l%wU�a�T2����]����	����R@�(p���k,�4���`>��-]�+����p�wl/s�@\ƄV1rfQG(E,5^pI�;���5.��v_ff���'u���Ϧ޶��3(c�ذ���LC%�Fr1y�#ok~�o/ZɆ���p2�jڗ�J�1��_-&*h�����͘*3;K9�;IZ,]qV\ڻW��62<��:�P�4�ā���ιZ�Vh˫�ś�v���aA�`�$Y��3 �>�im��@	<p֐(fds�
f#ԃ�G2GZ�٠�Z���
ut�
;�HQ�XS]��+r!C;��_u�K�CKKʄ
	��!��j��LI�ݳ��̣��]�wB�.��d<,,�6���&�dq�}h�	����+V*�/:�h!�x�[%�;�:���:��I�n1�s�NX(٩�m���3x
�XE`��fu8�,;2��CB�G;:��)����@�E25�|f��Y}EV*�s�s�X��ڐ��'�ug�Z4yo�ք��Wƺ��۵���J�@+®��&̳X�+��������Y���j勫,5LX�36��*i��Tzb��(e:О!�Ub�6�!|]�=��k7P��m���ڳ�nU�xs+?a�}�h��$$$ �)"����=|�@�!����Bҥw������z            I$�Pe�1:�XQs����y�BL��]Eڼ�.[��!\�`tH�6�A����N�X�,�Zn[����"���ic�Y.[�rb�͋��uH揘Sz���F����x��:�F#4�
�Z�#����xKbd�"{��f�n����"�2��H�R6P۬�6K�Z-ʳgݡ�J���u�Č���API������ծ��wN\{��w�y��ð����Î]������%�"��Z�J��eU�Q�Ф�,��U
]T]��B��!b4�n�@�u-!I���L����n��m�R۪)j�R�5P�4%�6TPQE�)i%��Um�-��DauR�^�j��B���T[i����I��B(��Ŋ-+I�UUWb%Z��ꡒ�#T]DJAe�R,��TYUP�YWRJDVS-��M*"�,j�Q�7Al,dQ�B�}T���/߿^T���.��\��i\SWN2L }Ud���k��v���_*$w/�-O�R8�HY>]�}J,^�K��8ǹ���T�VW����j�(f�ڄ�0�T7�����mں谨O���kvjWY�i��%���V-�j]S�c��ݞG@N�6\��6(^f�o��>�{oX���i�Qq�7��d��s��٪�B�+h�z@]Y���.�Z�*:�]
�A�o8�E���R�{_����B�����g�Ǟfmz)Cu�[h�ڔ�.�o}�d��a�oǦ��d
��5��̟8t�,�M(��p�v9\o(��w7�6;���/Kfv�u�<,~���drP�)�������kw=3˜\��|ˁS�on�;C�F8V%Y����_g�k�`Y�"x&�z>g
L�I`$�	��$����^��ŕj�t��z|UlvT�iZru2I�y7S��2k##l�:���{�/��{-�ۮ)���=����O/P�����d;�^]�o����=�nb��͂�}d�WX�G.�(zo"�3�LއP�;��;N�i��W��+�^[�����7W�D�&���k,q�sו6�,6{�(���BV�6���'\�m���B�]�V�6�L���1ȋ򳵫I�,Wr~ݬ�^6��h��;���滻{66&�t��g<��f�t���?<�o��:�چ�d��<�N]��ؖz �g�����/����.b�ɡ���K�^�������
�]��:=���c�Թ����5^�E�����
���C/*�r;�իF"1��W��.��n�ۧ+�ܼ<�vLlù�����2y��/H�J�l#��n�?o�⣺�ܤ�OXI��\庾��TN�B^��[J�/�W�A��,'��y����E �Q��IX�����Yɫ�;� ��x�B�t5k�y�<����N*�0���սoc���n7������)�^��6gU�>�IJ�U��̷����Fm�Gh�����v���@�5�}.�D��1c�_'�ؽ�(Զp�V���2n�:'Oot�:ieMs����]��t�v{��~Qn�Q�
#�|(��:��V	�y��	�;˰��^ �4�@4&n.3�U�M{+'p�t�kb�/;X�e{o�1�}����W�v��]FsI���;Z��orO�=Y^�ߎ}/ܸ�����qGJ�q���/��\>31u��BI�w����>�܍[���龝�ȫO@Q�*��GY��-U@��sѢ�E�~f�4��	��Ԝ��;��l�}�2˿�X�:k+ˑm��{�m�+q��L�3��
zb�V
ΪyV�[S�?N�sr�0���G�h�9{O���/8;hyŋ��@�}r�8|Q�c5�خ2�g�K���k]ʁ%��ٙ
��M��Rh��]v�]�X�6I�q���3/ˣ��A
�g�7��5g��[���-8���iVy���zyd���Q�F��k��a�1������ߒ���S�W+���y�M&H��~���ͦ�Uy���{P�k��"�$��{��+�ag­;Sx��s��@��J�A��ʊMG|u�F/ }���r�M�W�h��'�T�3;A�֦hvĶ�]�lSs6`���.ྷ�[}��w�F�zۡ����au}yH���o8��χ�;����S�{�%]AxzԜ5Q�+"��: +s��`jq��5�9���w�Y~[��[�[���S+�ـ�w���5�M*=`�@띾զ����Pwv�#��z�BE[�ڏ-j�6�2��/%�ٻ����@R5��Q�o5�+4�BN:t��q���%�ef껆��r�"C���Iz��D�a�vjD���U��W�%\wH�E4�<�z�mo��T�&��9�c�d�WH2kqU���tf�u���	�ٺ��3�؟C����ε�J�gz�D����:��~����~�ep&�Sx<�c�������9ڻ�1�_d���S�`zGk?���nPJ�t=M�7�n��m�"˧�qtѺ���b���t�WW�����֍-r���#4ۃ�t����X�d�qUϳ컮�GlX���FA���kZY�ruwoX��{8����_=�B�v�M	�2Tkm�7XV�d��������9�.L��N�f����Nj�
U)Rղl��V͊i0�f�a�`*�&��Z���C� ��t�v�{�w1<���:�����R8���}�4�~�               	��l2,6�{l����ŧ]�[R��6P�wԴ���\����ڸ�iU��ϗNX��ܢ������I��������ZB-:X�������r�_j�l�,&����'[��$FQ�kJ�Orn��3�32������Gp.�n.m^�F�u��^C�k܌��Y���^gY�,S��*X$^�%L�QߏD����0Θ���l�i'"nB����|m劻����UU��utAeUR��?KhE�ҍ4�
IL���KA�%�ҙBAAJE�Ei�]@�ڪ��EQ�Z��VR�Ҵ�Jv�%�T�����J�IH-	IH(TE"�P�


SCd-�tSUE2�e$R�Je#��UF�*��Z��J(�RDb��t��UPU
SX5T�P��T�
`UPRR(*#U
H[-aI)P��dX�5���s�_�z��k{�g=��j�Z�\�;#n��+�e���G�� ��4p���ZI861|�j~�ί|~�H�iK�_��+?<�+���||�j��/c�],EN*�p���eg���I�?p���(�e_�?�ZvO���g�_�fHxT��[����@���_��~4vEZ�W��㏷t`K�6{��"2!��Z��7*ž��;�>g�R����@7B�W��OV��uַxZ��m��C��M9��>Ւ���w�����~��N�Y�|����THV~��wX�|ˬ�4��Ѻ�H����v�<��+h����%=��'��7����>��b��������ybD������~���M�^]y�o�hI{�)r�-�g��[����}U_���@��|�C����΅���Z�}F���[tG�;Y�Wrm��.u_�B{r�����)�́�2���������yW�k�y���~ž>����yp*k�kӔ�������!�6yX���g�u4�V	s��ٿng��(�h용Q``:,d�5^�O!��j��m���||^��-I�'�����Tb��gMS����QY�=��;�����ۘN������P�Ol����t~��;=��HY���1��3�8�!w�#��W�T�����VGŅ�m_��+�ٹW�6�,'3%e0���zg�ޝU�צ�(ue[��,=R�(V߸ׂ�{�\U��~���_�+��d��!�2��f~w^��C櫉B�RC)�C��>0�H):�M�CL�� e|��{�X��{w�aԁ������P��8�4�a��!Ԑ�B��<�;��Hu�$
I��m e���KC�d�SL	������\��0�{�Mr�e�,u��ZzJfr�%:2���J�dM��7�����_�!�|Ha	l) _*L��&R���a>0��W�߱�g�`[%�$�I6��0��HR�cT���i'o;��{��!ˣL!��B@�d�L�i$��@�$�:�4^y���	��Ha���I
�Kd��L3$���C�t|�/����`,!4�Z@��́�HVja-�(}�s���2����D��!�@�!�a���@�I���Ka�����wڿ�=�I�Cl>	'Y!��N2B�� h�Aāf*Hy�Hb�M�����%�I�Q��I�j�K�A3��h�������Z��|쐴�g��@HN!�a��e$����IwRC�~h��|ָe�2�N0�@�ʁi'Y!Ԓk��$���`O˺~���;�Wt�
����yX:�*��z�!���������Mv=łrI�wn�D덐�rK��/������2
�X|d�$�)}��g�� �N2B�e ��Z���R(!�i�/�̆�6�<�B�S��C��K� u�������$)$��d*萭Tf�|��m���B`q���7��s���$�� ZHC�a2��2�a0�$>T����p�!h[�'�L�H[	��q,Ha���4�y���?7��<�)2����!gj!Ii�`I:�L'��|�Ϙ���9
Hml�P��<��i�GXB�Zad��i!g����=��Y����a |d<�Yi�u�O m���L d����w��l`N��y$)�āԚa�'���Y�Bd�2M�VzWs�yܐ�id�I4��6��C-��@�!�&�RJ����U�d����؄n!�H1��L?�5��Ž��>�1�'T�r֌;|�س���U����?I&�B���^�2L 	���I�������J�Ih�����7�c���k_9�󶲕���f�����9g����xT����^�e�q*V�"*Qk}�V����6p���ш�F�K�n�R�r[Tc�������V����ǳڶ�r��Ne}�=��Z���_�`�]-����HǷ]u��o)ު4��j�9NuĞ�}"�9��iPV3�!���HS��?}�{޾�g�>�*�>��|��꫺��˥ �.�$ݛ�¤ժ��wg.�ߝ:��}�閫�~���jV����0�1P����̢�(��F�o���!+�4G�!�0���t2<�h7��rO�ؑ5=�ۄ`k���L���	';�y�A�>�q�8���T)��<F1]4̓%vv���H�ʐ{m+��E/f�N�琾�8�;O�%���X�o<�|�����l�v�f���%w�=z�H0�����Ŝc۩-��Zϗe�N�}���G8#�O>��zf��Y�u�0S�o�k��^'� �b9��O�	����RKl������ 0�=����I�YDD{{\v��y 7���tp�^�����M�qλ7a�P�W��;�}��C}a��A{����70}T�aa"�E�
A@a�"�dQb��UQd+E�Q���.4~OY��.|�;��dSYC�Ɋ{��~�V�~��;5~j�ja�s�*�����F�֤���;}EtVv�o/ms�k~o�d7�z����g��>Ջ�^(�yqD����N3�Fn��n��z�5�.�_�.5���9�M��ɌI�t�}��uN�}���7��sO�v�^�C��H�|�߻�]F�����&�ͻ؃���^e�OI[�,\�k% o���0�:�����������Ko���H}0Tv)�u����7Ps��n��-�fn>�G"�cm].�7YN�
LVB��s*�a*��a�Y�%�&�c��\ș�#���A���?�!�,=J7بuᗜeM/9�b;�q� ��x�AwF/z�o�H��7+ͱ�               	���Ib���`U8�}cT��hf�,��� WAń@�PS2�{�컵Dg!���N�	ӥ�u��f����d-<'+zj�.��wV�DGG���ѧlV�����X&��7�/V6��n� �U�W�=�ʫU�&]�����P�oKu��坳x����=�/���W�%�=�����:�B��(e e-n�XΜ�o{Pe\��R=�NA+��Ț�)!�^_��W߾����QL���dRB�H�*����i	I)P��R,����B"
� �B,� (,���	:�

b��UE R�JAPX()�))��'R�KT�QM$>�["��PjR�dU�#"��;j������o?�d�(��5��XƖ1��;w]�7�U�}����C�&�G��tM���?~C�I���=z�M~�3������90w���ʳ�;��@/8��0����9صHt�d��y����Q;�rSz_'��r�C�Y�7�<��ޯ(j'2�N^tm��8�ǅػf2%�\K}�^�T�o�x�o�Ҹ6[��|z�``��{�z� +L���{��!t��\������{.�u��� \�9��gw�Y/8޹|q�ƾ%�����|���j�	:A`���햱��c�6\T���_h��rnw�ګ�u�";�ӳ������ֻ�g�����vg��{;!d�����b'�X�v�M�J�`�c
�uWx�C�<��u���˭^km'߳�;�G����v�M�S�Ϻ�
 r�ul=w�-)��U���U^���"_����)�n4�G��ޱJf��Wx�OEC󜮰�u��D��Wܙs�~ݿg����[�߰^�;G�>����v��\�����8�����x'�~�/A>@n�^�1���T>����e�0����zy��y9�*�G�Z0��>Ӿ ӆ����/m1Ͻ#E��|��f"��8�K|S�?�����X�?k=�Y�{��2��N�a�����~���TA7l?7\;���Mﻅ(��= 7��,d�{b��/ֹ�����9��b_�儎�+�6$�Y)�khٽ��A=+�OgŬ`D�sv&b~j�Z�7V��o���������*ʁ�z���|U����>k��������U�=�-�t�R�FfE�Zre������us�����xS���C��oGRQ��o����'��{�E.��NR��c�e��G-/q�<60e�7K4��*�*��{�LR��y;֡��i��z�E�k�3{�
�{w���D�����Sm�ɳ�|	]�+�a��.����m+U@���;���k8���,!���eׁ�E�L��Zb���Y��r"[�dO��#��Ym���=3���6޳�/}��_Ӆچ_��k4Dd�;�Ԝ�.��2щ�O����q��Ê�� #�Xo��0F���Ug�[�M=����{��gEN�v�qg����=�i6 _zY��t��)���
4�/�=N�B��x-t����mo\"��� -��-m�80�d�rZ����2� ��e�0���ƪ�_W�}sv)�;B��+��X?])������en�h�r��r�=�,+�$����H��ʽ��mc��{��sѨ�Jԭ*��ڽ5.C���g���}�L���Z�-k�{HkHT�w���+��M|�Wy�K[=3�H��V�$S�{�W��zԊ�����9�ܲ,;������hn��̮��p���3o�쇳p�1ο�}�}��Tw��@�o�8�b���Vk��t.g�p��R�8�Y���z<I=�����(�${���֢�v�%��_e��(��7J]yM߫a inr8��y5�jq���.��2�t��wiɉ��,t�`�/}�����{AʿzsD���ج���;L\�t&I4�t�Kjɷc���>-X�,���f�gR��bJ�lm�?}_W�G�`�ߊ�A��m~�)��ʱg��
�x�W��zT=P~"��.g�Y�,~�u�{ө��ѓ9�t��p^eg���~t7}I��&�ރ��z��}�	��М�w[<� ~����t�&IJ.�-Y�sݻ~[�'����ųZ��洲��Nf[w��HWf�A��qݏj1�<�däs׀̮�z�g+rm������L�ء���ݢɞ�,"�>�#Yk,�����@�c�{߿9p��o筟��3H�V���;��+���,���)�=�{�]O�� ��ϕ��4&�=-.ɷ������h���WW�<����Gdz�}�S�M?T�~cҝG�����K�ٷi�������V꒶�u��;�d��~����e�r�
�v�&�\�m�@��uћV��7�(j�(����_^�����,��Qr�-�+V�
���ێ]H�:P�Z�T6�|+;�+�x���\���X*�F���ĘcO�]�ާ�v;��!}���v��"t����8]�t
��&mÖ;�K���*Jk`u�K���9��WN�5_�ϯ�h �              $��\�Vj�,v�S�Z��]c�3oF��Jt�j��T6�*MY�B���PX�]��V�h�3�E�3���M	���ȵ=�'����H4[=��d�N�]�-�kQ��]V���i#\b\q��e�[��7��M�� =aܜ�63Q�W:7�.gA\d�4pI�t!�[}��oyȠ�s/n�F*�1>�;���2:�IA>��ӋN�� ���}������Ū�"�V(,R*���b���UJ�M(�Ea
J����"��EDn��((��QEY��)"Ƞ��"%S`M$PR[!L����@QAdR��|����֠�El�����oVJ�$��
����վ��8��b	��GƳ��O��[��]-�"曼�U�Q��k�珨��w��{�J\Sz5r^V+����C�hMH���j³{��b4�~�Nu��쮓Y�|���'�J���K�WȈՎ�T�y4}�<��/���l*�,e�;740�،��<ɼ��D\.��N6c��p_���&��a�~��RZ?U����kV���)��K�Ck��V���c�O��Y��}y��l���1R�5����}PJ��<�On|�tf߮���}W{~v�{ 	���k�(�|��>�J���(�fxF&G���uj�C�%�V�w'��{f�2pp:��h�=����o���2�\*8u��M��>�?}_}U�쟬~���Y��'B�A)�
�W�{��K0�^�����ǥ�v�ބWV���AS7s�8bv{����1�CZ~*�<�U��p��r��r���{=�^_�^V��lW+x���`st�{ō��=�O�2+~龰'#Y����\��v���.�"&������e��ܷ�R$��m)��/�}�}H��?Q'�������;u�^Ȏ�/�n/��%i��-������z�?B4�Bz�Cg���]��Cw��'GV�S��&UnP���&����G�����^�4�sz�<����]�S�K"�&�/_5x�����<ct,[�&�Kj(&}�wQ�N.=
��;t��4Z+��H�Yz]�]JlY1tv� J7\�td�7;������)���{/�I�N����Q�v�a|����M�=��;kh��;(�Z�Ͻ
垏	���������N�����Ժ۰{����,��}.���-�v}�.eg!����]������ڰb���ZD햗��@z5��V��۸���7~�oww�����DG�.�h����{�YB�$��+��<�.�C������Ư�s�@Ю���y���/����ޚ,��8��[>p��������7�OA���@w
�8m}KGbޙC���]J���.�C����>�[`�^��(K)��
�]&�>��׶�-�5��ʷo��C�\�*~y���*�����a��������ݗѕhŅ�W}w�s@��\�-r7P��k�ч'7�N1�_����Eѡ��W��|?b�>���nH1�U�@<�N3���_S�<Z}V}hr����*Ǥ�"<�p�c��i�[�D����z:�Zr���B���lQ���r�X�����<�f1G���e��ǲ{��<�8��Ϩ�{۱|���ou��3^�OH�bJ��"�nW��u��z��ٽ�J��ױ��R_
)6�<��m�OQ0�x{B6�u��w��ػ�����owĤ���+&FWq�{
X��7��_$�s�s�|�G�3o�Tҕ���N~]�ɋk��}S�Mכީ��9ZC�U�{~�W��d�/]<z�l׊�Zv��']sY�r�3tj�Ǩ��E���s�c�d/��-6���3�;u�q�m;~ƻ��yi�L5Ta��:��x��q)9���k:8�L����h�^


�����u.���e��+��D��k��n���]-�(�0���l�ه~�(ǜk>o��B���
�묽���R�[���O"�n�ƶ�2ƍι�ü1��ds8�u�Q�	�Ϭ7�i>�	����ȌV��=~���J��0��o�v�9u��=����H��K�����]&>���`�{ix˩`��".���
�ӯIyaM>�%��r�r�f��n�kl�ʱ�5��^�y����]��J��+��".��Mr�2���k�~�>��N	�e۝�߫S\*�Tڧu��;�)]�e�gk>s�gݚm�m�nŽ�ўผM;p��y~��>��ѿ�
�y�Y���Y]tS�g}�y�%�����U�۴�����u�[Wjv}WC3|��oW�ʻ�5H®j'�L��c���V]$�M�� 8�9�v��c�)�S����֯���~���S�8�<�e=p���n��T���7<>>߅S���ϳ-r�S:>7F�oaYR�ͷt{*�G��=��l���QNFq;.��1�<Gʞ�x�Ts([�����2�v���&K��y�fa�Y�T�a�h�n�1���a�>��Х �]W]m��u��s7�����cTZX��u�z��۴�0&������e��M�ݛf�Q׬Ӷi[[�|l�.�ʙ��|��ܟ��2����x.�l�<�y�j�Ƿj�fF�+�,^i�wT��Ե��h	�S#U�gWY��w4�tyz��i�c;�[*��U�XYF}�$� !�^�QV7::�6+�3r��v�VHBt�^(�/e�f�ï��	5��YZ�~�C1^��[�%�D�]йHuZ�֪[b��~mL#���6딷����ͻ۽��:�EPq�*m��c3�G�ʏJ�̿�vns\�    wwwwp        URB�ET`RLZ�SJߜ��/iH�N�6�w`��#�+�Ct岶ա�f�6�_YpwH�Y�-Km�L\�md�<-��Y�M{���ʕ���#vo�r�z3��HXA�N�L7d�-a��)�h쐛��u�2ŀ�Ѫ�<�������N�"�ܭ� U�w�\�M�9И���*��vw�٨��X�l�Q�9� S��]7�T�NU��nv���y�s��y�wv}���@X�a�)�4��Qb�d��P�i$��"���X5P�()L��Q"��@��*�RRJE�R�R*�IJ�EU"�VR��?C�wZ߳��%x׍v���,a�r�Bib.���U}dl���k���?
DS��g���fV1p+�|ԁ!���m��7�<�;�_&O���7��ey^N��TS4P�y7u�&h�u��ܶܦ_���e�B�S�9��[u��b�_���v��^9�ۮ뀥t��ova�h�׬4�y��t��N7���t�P���8���~N��^hw�F��53fq�fM�X�i:��Qc�˯Q���|�i��;��Y�+tZa۫����}��W�V}zu���u0�W��_�ՋnJ�+L	��&E��nJ�<�Rnc��9������L�/?u��Ƭ��NU�̾|�u�ޱ���&�F7E������l*;���w��v����n�x�V��
����N����\��n��Oz��]8��݀�^u�z�СD�Z��nyP�5���^�g�fuS��H_+Hu��|��b�;z�����M��1��~����-����rŬn�;\�Y�Ql��x�.,(��ExP�%��y3��CX4��UFٛ���F��&-�oϸ��.%Z0ޤe.��f��l=.�R�+�K)	F�Ș�/�s����f�a�=�)ۭ��	�����;x�t�i6̡C*s5��cյ���V3�Zo�Q�a
m�M&=sX�/=�{����4w���S�i�°��o=���I��ѷr�+��(pw��(�]r���,{�t�fUQ�)i�/ޣ|�=�o>�3���[�	�gӚ�����k�Y���i릙�Q�)Fk���su)2��>�3�h�Q�U'��^�Q��n�t���׽�+i���W��^n�3G
0��Ʒ�C��u	�$�0OQ�J�I`��ѣ�oxg�6�"��	���W;�Rw����Ʊ�|�m�q�x��6<t�����d�RA��_�![B���*�eS�6���=&%��N�dW@.����>�R��{լ��m�f���i�x���a�L��P����+/,U�m��əB���y]�9:;�Sř}uZ�cn��W�U��w��-mޜw����>ʨ27F+�c�հ�ѷ)nyXN>t�7�9u3�w{�vr�,�ޮ�t3iN&u{���ޝL�\9t�z��Pu���"�N /k��:�S�7�++�X
H�ȭ�"�Ğ;�{�Z�R�_�G���=��ͼt����M�k�[Ǐ��j�Nz��+�n���h���~��k6y�{4pM�L�o.��M���{~���ٗڣ��Q�T��0z��m�(1�����ԝf�G��yEv��)��6�9Ϲ�z�&_������Ϸk��:�:�}�%��4����l�2�u����B�1E]d乇=1��:�1�]���@�W��m�}�]���y�v
�� e�]�������{��r��xΦu�ȸ�g���A$0�:��f����sJc�r�sv��E�>hV�ӝ�/����o��՟*�7���Y���~͗�����߷��w��޶�b��fkLo����Z6f��o1Sɗ��r�j���k�q���=�9�Ⰻ1����4�5#3��^X��V_��S�V�>�u�j�X9���v|4W����v��+w�w�WvB曗J���¦��]஥׭�,�.�X�-�ʛT��Fn�9N'}\W�
�5�6�Tg�8��i�w���S�_9�a�f�
��ܷr�Y�n��n��xtA{���f,�4�K7��5.�=�b�},d�8en٥&-Q�]g�%�{͸慎/s�_�k;+���w�_1]��3i�α��T�e��sz�q�W��yB�1�����]���µyb�vU���f�_�Ys܏���;�f�ez�J��v��=}.�{���:�mä_:ɻ:�7���^}��掉��,/U��9�"�+�<���L'1^�����yV,]l�T�7�߹
�~�S&y/T[�e-R�<��M�4��٧��M���q�8�L�ތ�z�h�i�mf'j�Ǧ4�>*��1ϳks�g�5��K{<���C�g��5��%�c��^�]�I6�}VZgu���n���t��>:���q�Ҳ�f�1�9��L<t&�KH<�;�;��+�k~�M�i�h�nmæ��y�y�ri^b�3O.��m
d|��h��L�}�W\�t�U�^�[Y,<���#��#Zڡ2�Z������q�8�}��4[�w9۶w5��W��(��9�ܥ�D{���r�3�j���g�b��<w��%w6e��.��˪7��s���r�{����-]V������Y���W����ZC�(��W�S4�ua��E� \�{kzX{�7$SyL������g{E]�r���ܻ�˚�]s�N17��;��wTЃ�Yc�=�&�:r����Yn�j���B�5+�{~�!��N%��r�|�ܴ��bj�v�_���a�s�Jkt}�W�L
xV[�}sqj"���'���S2�J�Lz������d���Ӊ�4�v�i�i1�ٛ���������wty�;G�=M�3λ��y��3�u�A�B�=��q��,��w����ǯZ�9v�5e��ڞ�j����'��I�9�q��=D.$	�s�����љq]������.�/�B�c��N9|�O����(�ɃIq��ĉS�ȩ�9"`����&����甮�������>(]���釟W_�.����u�Y���+���Q�׸��^;�~��-8;iҲ��7���d���k��7��ܳ<�6��(؛�*�y�=>
�ϰ�VZ9�W7+Em__�o��ل�3dqA�Vi��NY����U-xT��/�YTn���m��緇�w��\�}���л|������Ov���<o��=4�E�:m�@�EX�]�7j��Hg5/+3d��l�\�θ�/6�hX��X��.��!^����%��Μf��	�&�ۦ��=�
�k��T)���{&��뾂��}ouU�g1*m�4�_q �o�@����WڮV�Ʊ3;Z2[�c��5ubH�h�8�qt�ƈr�ρ�2)O���z�,W*��VhXr���|��f���QeAC�iLa�!f��e��{�b�_1��r:�9�DQ�Ӽ��               *�b����e�����Cg�[�:�1(_l��,#�J-�?�%�/�t�r��,�N�AC�L�⺖6���:������ښ�0f_p5�P�T]Et��]�р�ʜ�
,u��]f\]"Hwj������n��2g3���c(^�p����S��[(�y
���9�˝�(�n"�Ȇmjǝ�ǁe7�)��Dgr�U�%M��#s�[�7�� ��8�rE��}T.�X�������"�5JP��e�UE-�QQU���l�)�Kb�ŕT
��UC��e �Ji#��((�0X,d*�i*0�QM)t�%�L.U7vKij��Z�}�d�7���b��=��}5��O
A�p��ꯪ��rk�xM�L�����ݦ=G�v�i������ǭr�UMd�Ln��׵��w�o�y�=��q4�w�eS�篾�U�Y�|%�̧KV��#�몍*1g{�zΦ\���/��u�Q�h�7�)�r�g��|�]uԱ�TxU�1R����{S>�*�n�@��Q�+�A�药=��>�<��4�hp�ݗ���Y�ix�X�wjoԤ-�<�x����ɜ��tM�f�*�n}N��3�]\g����D�p�qh����lF=��h@��^T�cK��k�b؉gzj�F���Io�I�J���n}��4D*_�u]깉�٬>Ɖ�5��W�g��9����
�.�̥��o;��C|�&/�m�n����'g�8�=�N>N�J�+�_b��q�6������8>�^������J�w��|���=���/�2�Z��)���wk���q�r��+ݳ��E3��%�m��=.v�ڣ�e��^54<N�y�vr�<*r���X�{G;�g�M#��y,�\t�陋�1�e&�UR���Ϧu�����Z���[B����E��ec�����(:�B(���v�=ٌp�kw�5/��+�m���z�~9~3�܈�ZM���3����k�{[8cVi���m"�gĲ�~xu��<�4k�vi�7�,o���Ue����s	қ�{ӓ���?��[�]�,�\���:��|`��WO�ϧ�����V�M%8�a4�Ӕ�Z�5w�k��뇢i�n��C��U�w^�{���Zw[�w���]�\�V�f���*���Z�u�Ϛ�7�J��|[~�ٚ�E��c�3��l2�ǚ�n��o�H��q���&,�r�M�Zseꉒ:�;�����+�R͚�.[�^���Nj�?LQ�؝~3o]v�}?|f���j�~���W����xV�K8U7��чl�B��jy3�����Qx�Wy�;;�}W9Gt�-˶X��z�s�cػ�r�p�M�x�]ב�a��\�f�k����T7NT��$I$�H}����>�ut�VܾѶ���˹Sc�J�0�(�P�u32��P��+/�z��7�j�QC��+II��]�����o;3*tR^֑�K�.��r� ���Y�ڿe
��߄t4���G�6�S���"A��Q�ź�q� �표3���5�x.�kʗ�_ո>O���ts9ƽz�*��jZw۲j�a��e��mz�k=ќі�GOW�f��Ln�I�f�����gf_;f�����;�-����mg,�Y�����-۱tŊ��veD�i�篘�����U'SO�V�4z��_]�A��<Ӭ"_�����7N�ٿ���W�E�=�&�pW�%�̮3�w\f�7s)��}�{z�=M�^+��\��䓪������{����`�2��W��]������5��=�q���jY��ݫ/`le��ɲ�c�te�ʊp�V¤� ��8g��6_߽����µyj�Qܪ+�R@�\�e_��u]j��6�j�sF�9�do^ד]���&��rͦf��������(��Z1�r���z�=}�ZƱ{ٜדy��*ctV+�����p�Lv�l�5r�V^�}q�;~��i��;����}�|"̦��[�v�{j똮�rXHk��.��e�QN]�f���\�fh���=g�p{����"���Һ������U"5�]_w����z��r���n�r�|���^k���yf��>bV-�9L��L�}�<�n��~�,_0��.N��V���L��o����fb�}j�5�6�����swڷO2ݺM⦩��B����PeSQ���U}�eV۷�4��s/��W��`�y�k[����T0��i��к�����4q<���4�L���9��r����9�/c�v���W�u�����;��5e������2�Mr�7ʖ�e;�Z��tc4n�	�㾺L۪������0�J�j�
�9��xۗ���v���v����TwF���ee������Z�*��z;���:κ�6�{���蛍Vs&�lr=�e�Ƿo\è:�ě�tgξ�7S���>:N��f��tf�^���F�!�.m�۵tG�-{���V�A/�u�>������_��v��
�oj�f��g�l2��������S>���Bq�4��������m�l�kiI�nγg��qy�s��xͪN�1\�z�^X|}°
\.	u.���lں�N.�}=�]r~�+����)c�t������niU�룀��B��u�}r�H|;g��q�j��Eހ�p�E�-]&Px�]��̣>U�ʗ��5I�}�� ��~u�
��Y}yy~����w�$Ë���*����`ˢ�e��5W�o��-�TT�aX��x��U=fu[�ʆ�� ��������Ϥ��gq68r�;�`�ԣ�Gɗ�6z����t�m\����A+6Za�(��<��;�!N�w.>���P�6o�Z�Ad�k>ut��jY�B���*���p��w�[��w\m�I�6�5|�Gh�iy�Y�k��S�U&�N��I�d��{��fmi-��P�����ѡ�^iܲ1 2��^Ts5bS�!�W��(r)����e���C����˗N��_]+v�V��=��x=xô;�[��=ύ֔��6��R�u^�wi�VnxKwR��1��+�|=�T/��h�a
�WgfV@�����u�|9����j�e�NqF;Xe����t軮�/����U���G���m��ˬC�A�u��+7R���8D��q�+7]
\�"g�8C�k����Y��v�z�_+n!^�7�U��������>ȗ�<=u�P��UI�0}�.�Y����t^4�^�w2��¥	�X��]��07h�FN�y�����q"�����d"�s�q�J�S�ܮ��it����܆�ɟi(�
�)X��Ϊ�^��z΅Re)�\]���}�>��C��q4,x&�+wx �o��,2����,�gAGi��]lǆ;L�h3�!�ǋ��+J���]�U�6��E��)��`=w�
���\�	�1���6�N�ǚ�S]�J�q������v�               U3bZ�[yJ��s�˾���^�:
yv$�+�(򦭧c���*{�������˒�F��gJ�Bӓ�x�����q�������}هR�K����w���Μ7�jC�B�4Ptt���t��N��VK��[�k���CvȘȕ�X���w�8���V�so�ŉ�y�ѐ=��;�N�P]�|'i��9Vr��ȸ���*X�p�rD���I�U�B�]�_]eU��a�������]ҝj�RT����ER����+)b����QT�	m[R����(��QB�(��En��MUĤ��{��h�Y/]b�W+�� M«v�70^�\�M+�ZK�٧M�N�gG7z޳�n���e�r�]'�iQ��k�Q�k���-��l�o�8>W\�������u�K��;��,�/����xӔ��e1���#��]��`���
��2� �]+�aś9�c��u�e�T�R�h����<��e2�텯��A����y�s(�a��k��s��p�I�V�[��\o۱z���5�k�=�p\O'��GU�p��Y������:�f��3�3�Ǫq6����@�F����C�ڣg]ۤ�ԛģX2N0��4Mds4����$��.��V?K�T^�+ux����E���䊲ý��t5>��٥�A�C#���u/?`P���~:S	�z�S�C���h����MO$wR�G��#��e�/��h��z��#-uR���擿uW���=�E����ƭ�~���C����a��j�l��c�J����8���'[!y�&I�4�uYt۩2��NnX��R��z������������
(�OL�=�ý^֌�S���.��&���{Όdx)ڹm��Zu&{���?����ͬ&-楏���ك��M�Tv�㒒�&z���<�Gl�by&
#<N'�SXkݒCfUdy+��~_8�s�:�J�Z<s�7��4ݾ�N��d�VG�����v�� 944�_��։�1��Mf�`�/�f|Ʋ��=��/��&���~����_��t�^h9�=�g����/?x�z����ܙڔ�k�5^u�>�^���2���q��f�մ�e/3��A��ُ�����gP�a�2߅�
����Z�x��R�P��հ�0�>��!ɹh��N�}�5dҏ��0~9���K�Y�pm����G�ўQ4}aO>�$О�d�Q�s�9��������uBy�Fz��/&���U�^�Cy�Q����R�-��D�n�j+�����k��e\f�9�p��l
}H_uO'*��{�̢vw"�4͆��t�^�����Z	釔|&V�ۛcT�«�0��]$��ֈ!Tw�Fff��rm���5z�^�G!�H�{+x���6�q��ֈ��[�l�u���eJMgL���/;�<�tc:�y\��ޫ[��u��;K0?k��L�o�r��=��=����!�Y�i���`���_��q,�R�_	�4��I�߰_�b�n�t6z7�"Ϸ���;��tM�hߵ��z
�&^5�nn5�SA.�e��,�;�s�)����x�����������غ+H~�슑��y��0"�k#.��<A�|��!^޶J��9m� ��;������܎��e�y{՝�R�F�=�\=����f�>Q���ݿGI�1����٬(���aV<��rb̚���Uj�����wx-7mr3'����B�elڷB�c��.ʳ����Fo-P��Č.�c�JL�r
j���<�ϱN��/v�$£�+Փf��ݵ��;���N���h�XI�&h/�5Z��w��^"r�MoiQ�W�y�!֪8k��~2wX��W��А��"1���EHǂm��ք�n[n�Y��p�R�:��1���uz<�{�T��Ug��&t�]p�6+��U���T[����x��"��v�}]�3*��\�$�x�y���r���ٴ?u�-���>�W(�ۓ��E�3-K�P�)z���5.��s����bC{��&�]��@������Li�W>����I�5}W��Ԉ=Ѯ���G�(�{�������p_
͍!��^�7�IpU����¬��/�ro{�aK�||<��I�P�^j��q��Q*n��'cA
il�;�=J�(T;cn�&��N���5k�prz��#�YJ�K���W軤Z�CO˼���Z�6D�J�R.(q�n���D�5b�D((�]Ujm^ց���w��ag��k�8Mox��^��c	竝W	B<��Љ�ݗ�K�[#�����{��7��,,9y^P�[�UO�o�G���3t4G�����ۥm�E��K�n&�r!.�θ̮����)�j0rpH۽!Q�۔pp�t���\O(f۔N��<��8�h��v�L�(+v�j�:nJgT���6Ы�3V�9r�6%�n]b���ӽǍhHﳴ�:qu��'��AY����}q�M�)a8�$Uś倴��k�:�(9��V1j��Újd��)l2�.��
�}LR���d֘��<�Ρu�fl�f(�*�S���w����j�               **(�^킀��rs��s�f�̎_T�t>�]�U!kL�������E�[�:8��u3�1XP���=*L��V����I�^>�Z�GJ�E�1V�t��:K���z�\>�vc�
ۄ6�+��r��
��:�yB⦘S:m�:�����dc�o#��KԤ�)�t����s�g/v9U�#Q@���0pѲ�+��R\�f�JK��{���;��~ٽ��X�4"�av,(�*SIUB5uKt�R�T�ʢ�(�*ꪆ(�B��UU�T���T5J�E.���L�F�P�H�����N�^5�t����c��9����땉�6��r�~����y8	����v�'�&Ǜ!�rtޤ�kuPIy�34oHz'^,(���A��wႽ��LV����;Q�Fb�j��*_1N�7Kr*D���"�6���GN��ȷ緋��t֖�կ6o��^�2l[Iw{ݾ�\R՝���#��}sN�%��|6�锎y�������s^�vKG�Bm�}�8�Q[Œ_)�^���D��7k7��U(^�����D:4�{k�}��kD=c�ܻk����c@�zK�=���5��ӟ�{�f����6Q�H��Q\�)
v���y	�C�$'��K��ȱ&���@���b��b��kF�����5��P-�6�����u����~cm�����t�^9�[�:�=g=��NX�Ӡ)��X�x���A�(f܉�� �0M���{W�QMn������EY��|�M�s���uӮ�i��U�&�_]4�Hi�s���&������L���xк�9��������7s1azb#<��'P{�Z�z�������m�&,���re��o5Ώs_�n/X�jL�`ߣ�.��0����kۻ�v믲�����dI+A(ow����:��+��d^��[�X^�gm/�nOpG�5���h�V-����n���]�_�J�m�C�~t���)t���1m���*-��ʎx�O,��[�y�N���g�{_�N����T�7J1�\�\O�V,��A6`P��LX�8�k�N���s��mEa��	�I������\o��u��~^�.��f��ٳQ3G������#��]���SѨ�{[=�eq-y9Fg�-��
�l�c�{��5v|���G���6�ߛSk;��+(Л�����;�"��A#��"u����ï͵Z;O�����4���x�{��k���4sU���_��f�;m]�H�����7��]�F�--���RQ�Z�ܔ���t�˗g��"�_/45~Ǐ_����.;5F��2�Yd6�����f�m�R�bދj��a�L�+/jl����k�征SYWW�R�Q
��Z�QW��2�o{�RR����y+̚��Ϭ�!�&�]��F�(u������O;ڛ٭�Q^v{�R�!=�=x��ׁsj^#w�޹�t!�0+�s8�P�i>��)J͝�NK��k�d�DlC��,Ts���w���N����O�?�{3�^{=L�I��v�k����ɞ�YZT���5y��v�R�M-��z���mxD�B���z8�#��z%�<�<�9�|���P��٧��^¥��y�/3Z�7��:�x׳w/Yj��r����]櫫�G�� ���+��|������%�VCu^;�Z���t�����y1Q��5����r���m���Rf�3�xD�gI��+|/˴���;�s����2ϗ�"�f�/q鐎�h~��?`���r�/Xή�}3������}�Xf6+��v�O#:�ܨQ۽P�3��D���UZ>�>�4V��n텈m-�u��ޣ՝PGu�e�#& <ڕ�ʙlmwpB��	������a�W�����ừ�WD���CϏ����)sgT�*3�Wə�ٵ�h��HGj�-�RV�>��ٳ}�1��V�4)|�ڸ�*l^�{���<|�ض�����7x����E���TX�EO��۰��ʶ�ˊ�y�ߐZ�o;V`��������Bf3����!�����f���G��X�'M_n�1�C���"<����1ǯχmD|�Iq�Hzna-Rxd��߽H����.�̭��z} #�����L^~�Z��)m�օg`��{+SX��YGAd�}��Y2L�j�Z�2<��r�se�f�%��v��Si׭Sf�,<��w��&o���9��g��th��}^��H�<<���X+�>������C��^��[;#W%�,N�#�ݽ�Y��,^-)j�x>2[��T�G61ن@a6��>�޹z�(u�F(�t�.P��6��w���M�1�*VW]��K/{�5wU)����Q
��>%l{ծ]�鬆]Yd.��ܡD>�)�n�r�C�^56���5�}��\�2U��߻0!�`��If<����wRUƉZ����#����ub�� ��)�0�����	�^ͩ��m�����ds`V��`(��F�                3Q^7ך�%-�m��%�*u��7ڌ���V%_e�Mk�E/
����!��g3P��S3j���z�0���#���m�.���5Գz4Evh�ק"���\"�k9��_=�U��[����X�����kM*2��&r�;/���]�����/��l�T���e�g2*or��.m�ѡh��m���t�s4aM8�iM3���rH�I�"���\�B�Bꅁw��M-�hYKT��bŘaU

�(j�b�U+�)X�MSM(�4�Um��Q)��TR��R�)R�*C
qE-RF�j������WuM��]�Ur���i����n���L]L��MB����Cn��(PУ�w|���ߝ���\0���^��A�+.�w&�^$��_����W�^J���evoH��tkfP����MN�\� �SZC��a٥4�C\�w�k��^i�'�������4)6,(�>�u�i�ֻoKCNY�P�H�[f��H�'ө;²]Q^�T���_�΃/�N��DR ���q�o9傶&��3,T��{�3_6�}����-�PQ��xa��t������}vG��B*��)-��9V��<��qu{i�v�O�TLp�rk��X�ӹb�
�[q����iJ���֪̆߫5�iF��X��N����^�%�f]嘦�����n��;W����X��i�z�����5�����5ڷ{�w�ū�D�%zN�6FҬ���^P����wf���������{N��IQgaSd��P�{s�7T:�c���Q=�3?�;�'��Ԃ��t�i��fk�ym�C[��ķ57�{mL,8څa��ٱ-r�b�	e��.7a��wN���pu�%G2٠tZ�$����Mv��O�G��s���Nc���U�/gey�T���+J�3�̍�U*Ȥ+R�����Cڰd�hWH���Se����A��(����f�Ꮙ��&��m*�w��(��ujD�H��NL��Ee�ޱW�ả�!L����%�ֽ��б�M2��y���[�����{&������h 哞��T4BJF�n|Siӽ���sj�4���;�R�U���2J�5���/H�ws{�%��+��ʋ�B{7��@p�����Π�{\�jp�I&��>ܽ&���/�k7.��e��$�0>���o^d2�:�#%���*��fnW��N�N�iU����H��5���x*m5@����%��v&�[&�֢�x{���`�<g�}�b�ڶ�~d�co��d��~��u�l�ys����h����e��(^E7ka�Єs�|�~Y5��a���.ոvN^��M��u�X_��WM\"�}�w�e�N����Qp�d��|c}1�-!���We�8��kR��r����xq;¼Uw�ō�Z��:�{�5v�^�lTG�b�y4/��z���<��9n-���3�lKw�0�~{��x��o�:i����U�H6N��fϠ�Wl7���)[�L��J��j�(�1yX����IxF�� �f��x���)u�~�c�	%�=�Ƶ�gz��m��.j��wf�:c�u}ūV�]�r���
*rJMgʮ1��k�V�X}��Gƅ�7Vz�矡�|�x=Vy��)�g�'���î��	M�{P�ѕ��B���~��N�@/�(�����Ҫ�VD�5Vb��*<yu��u��Ts.��ص����|/�V�Cn����}�O=�T������LVux�ڴB(R��{x�c$�7�H�tF�%�
Trsn�s�J�wߪ�
�p����}�s��b�h����r�����N���/D��Ұ�qe;��0n���WZ���y��	jόo�`]�M��1R����{7~��9q��Q/my/:/��d�\eI�O���8���q
�&��e��}��hy�8���5}�>��v�\:�L�V�
J��#o[�㐗P�F����$�v����P[}�n��]������zC����o��L���}�T�wK��k���D�|H��e+�Fd��w���q�\z\X��j&�qĚ��m_)��f�A�������^�M�U�.p�E{��[ϡ~N�z��<���N�#��������������`z�筦p+��:�7e�����Z|jd~�[T����`g,�L)N� ���|n�TqJ�ۑl�:IwXro���{�<��e��9�u屔ݭ�s,Y]*=>��О6��gy���:��t��{{�&i�6�v4��R4uz�zy���;|��ѕzW�����ޏLH�^M/�R���Ng�X8�k�T����7�T�VP��"�������vB����B�Cq~��~���ԯ>�P�^صAh X傍ua�P쭒��4Ju9.�4�u	���9}�6��]��[%d����/F�8+�zz&5�;2(:����ʖEl�3A�T�DMˮ8B�A��k���+O	}�����E����6%vuj�Nb8�ww�Ϝ��Fq�������9�i3	��%A��9��%B�m[T]��le�\[Yin��d��w�t�A6Z�G�®`�k|C���s���w���               *f�1�U������JE:K��m1�/2p��H x�r1�{[�����s��֬ݟ����lu[b�$�*W[>�(�w7!���^0���,�O2��Y8U���c���w���hV�aiĒ�u޼M�aZ ��3�;����9�݌�7��NP�}�Kj3V�k:E��n�j�T
���P���+\�EėQ|���df���&���M�����| �_U�VPV.�斪�����l���Di���P�)j��Ք��b7kk��YM]��i�h���4R�R�YmR��j�	m�v��wE�E�wWwuB����*�2�R%QvTiJ���R���Zm�P�*E�J-�Y,`��T)M��U@�E��X�-UUPUP��UP�i��D�����V�CEKK����UuV�c��Oo,_��*NG����w9���#�U�^�r��B�%�I*q�G�j=�k���@��J���[s�V���H�����s�  �R^[z=�ĞUCܻ1Oj�@��Z�/}����;�cj6b��Y�������]������9͡{�YJ��k{��87�,T|;�T)U�q�����Z8<�t#�n>��]����թ.Vm��-�4u��q���I�Z
Gڗ��n(�X#v��:�se�����[xр�{*)����n��5{Ls�%߻M��Wp�nv�ysDH��dQ�<i5�*eV�r���8��}cʂ�����{OfX�eM����MX3�b����W���r'h�yw�7��+����K��W~���� h#-d�[i#-)��y��C��_SV�ċ��܉(Z��z�n?߆f�R_�*�o��5�igc��R�}�,�Cc�Ʊ8�k�뉩��n���r��[���.ϐ����C��u�Id�N�P��~9٤�/�d���y*���ǋЗikܗjƊ�����а|ɣ��A�c�����_��p���%��:x�_�0DW�[��r��+vQd��1��_��c���$����HI�D.R�2{ڰ��q����#���=^"7s�pBޢ�e/�2��F*>��_����'Y�	1��F�E�36�ʪ�Ԯ0��Z;��F7����w5yiO՝�?{I�d�7��&�3O{�A�Z`�h�?�feH�Ӿؚ}�L#�t}��zʰ���[�A�n��U:b��j�#Y���o;�k��aŽ�b* ��R�2���%C�d��sf�̘+����>��Q<�S�<ur��lz��{u>��m�����D�oa{=jhQƉkh�M��t����q>6�Gz�w���"{���N�����c�r�_���5{��`^yF��[�^B����8t�mj�ExX�O��9�=f�䞗\e���3/�n�/X;G޼B�,Z���&Ɩ�o�@�p�rCW�AF�vt8�M���,o�O�Ƃ�0�幵���ˡ��3j{�_s�#B�`��#^�7�IL7Y�yw����-Ey�7���uƝ���n���tnl.+w�Y.}m,냏��Y1�v{���x�oV���PCY�<]/6��zHS���{���LlR53�ה����<���߮z���}U9-�J�Ov	�oq�FS�:��ެb�F�Pޜ3�3!>�9֏�*�v$׆��4��MX7_��8�&��Լon��}��ks'i&Q� o:�b"�Ӽf�C6+��|���No��<��3i����!<��X�28�s\��j�%fX4�Q+a�o�9e���)�u���zj�=�]G���EۮvO�#�9.� ˹(L��d����-��Z,�q��2Iwݓf���*�hwlud�L�0��=�r�fU�si��y-�@W�5�/q���c�]������f�K�)�H�j��;F�<����ڇ��I.��[3�l��r���ⲇ-��['�{=�/�4=�����m�O��;���}{��Ԯ������a�j��C�Ӭx�e���C�q{�͡��]n��"��
|!S#+o\=��0WE1&�������wӒ�����J��@�>yHN�=�;tQ���AY�7w�Mb�s۠�;�*���8�z�̆zϊ�Hζx�	��q��T��w���`�f�Mu�B�ey����m�ݑ	v�BD�[��i�{�c�mkMx��}�f�j:k��Ŝj�ܺm�Ӭ��$b*���E̾Ӡʊ�V��whj���#���X��xp,Ѭ�*):��H_�e2o��v�s��e��wW^B�NQ�wW� �z�j��.��-S��+|����a�f%�%�F17�w�%�e���h8�v�Ԫ��sF^ד�B���e��(i+�;���U?^\�ދ�X����1�c;��po8����Z�G�?�	?��
��Ҫ�b��A�$��-���hBB��d(�HHC�1P���3P�p�p�]��{���:������&tc�xN�A��	�$��V(@�d!	@����C��a3Q2T*jC�i�����eC��J~��2J������m��"E��a:���_u�k����|,6����4L����#�P����oiC6�.W��B�&�~-l�Ġ,>z�s����C��~ߡ����I��	$$!�`�� B�!�
������?BB����?頟�C�d������Y?Y�i�L�����4~_�����d?�������2"$>fB�a��%�&O�����ܰ�������=��⌖�
��0J��^��3������`�f������Z�j]���?㒀�NfJ����ՙK�1$$$!�~��8& `�V@�IR��Уl�XXg�?�6`��?��}�B���?xBBd�	�@��4��&�1�	��O��3
���?��d�}���>��	���g�f��|28~���
?��O�[�솿�G��#*BHHC?��#<Y�?�C�h��?�I���>����G�S�}�Y<B�*�?��+�~�����!�E̟t���~p�8��/�$�&��~�|6}��� �c#���~� �����d��f?�����2�&>�$$�%������a?�'A���'�h�}��O�%���pN% O���$���$�4�A`�O�c��"�p�X�����2d�2M���~�2Cϧ���]4��@� �B{A�kR��*�vl���p_����I	zXQ�����!�H~2BBB�g� ���!�O�� ~�����I�������'����!�I�HX�?�>�>�(���P���ȓ�|�{�a����%�}��/�����RBBB��O�?i�?q/��U���C�t����I����y,��B������?���$>��Y�!����!����\����!p��T�����~�ç���C����O��.'O�g�������/���O��P��M���~Z�Â~�����ПgŇ�B���W��$1 P)3$?g�}�#	$$!����?����@'��9�?��N�����$��?0?�I�A�D�}D��*&���P�ND�w��~뼚	���A�?2'�$?O�Є��M���ܑN$���