BZh91AY&SY�Py��ߔpyg����߰����  aS��         � 
         >��@� ( P���@ �ES`�
$I(�-5�kl s� 
� �E�����X,�
P�       @˸ *�5ʫ6���2el�z^�8�j�`����z�=� ��W���D��:{bn��)���l�
�_m{��h·w*����z- S��@Ԋݎ�}��x�Ͱ�F�@θ =�EYYj�)ݺ�F�"�=�T�6K��۫m�;�Z��g��ot�Ʒ�]� &�s��;4uo{�Cůukf�붳�LL�]g=�W��[g6���W-�{����/y����l ΰ �M��dz�cw�+͡;ޢ��z���ŷ;N�\��� \;�6ɽީR����yxy�.����t\ov4�tu�ݵ���-�����ܽf�s7fuB���m�f��� 3���6�a�vH��#���A�&�pn���˗[�{�˜�3��{մ���*M��*��;����pt�۰\�t:������w�����9V�;���z�@"w�ji킀.=΀Og��v�{;ٹ��{��m�����x��î�e�I�zy��{�n�皊T����Or��^�ݪt;b��o{�S�@�鹴��9)�\���|s���"J�       2�P`  � jPPJ�`  [  @T�T�) �440FFF�h����!$����!�  &&#5?$I55U4=CA�di��h4� i ��T4��&�M��L  �$�CSF<��4b5M<�M=�m�'��zHfT�P0�12�	�`ba�7�$yF�!�$��aiUU	*�Z% ���b���8��6�
(#`���;�PT�GPz/�~p��h�@Q@�"�_��8������e���,@�1�F0�$oH��(��z�TIUET�lz�ADP=�H�b	�$0�*���O���  �l�>�������?_�5�0313������ �1�c,e���,e���e�f���2)a$�z�#,�4�LeS���	��h�3�+�c4z�#)�0��S��`�1I>eZc�դЙ�ژ�(e%M"�c4|!�c*�1�����1����Lc�C2S�(e1�`�1�1�1��8b�!��1�ɖH�3�3�$c�ь���1��F\&3,c0~��3F�1�~kM$c(x��P���L��1�2�M-��0֐�(`�p�1��L�1�v�2F1�c�?11�x��2��1�c5���h�O�1�� cǉ�e2�(�C4�Lc(gRc�f��,c$t��1�	�c�Ɍ��p�����K��&�1�f��?2	��w���8�R�21ن11��!�Iŏ�I&3H�&�fX�Bшf���S0�2�Ő1��1��c$��E��d�?1�3[�P�S�e1�C���1�G�c,c�p�2� ���1f�3��i��#�afM
D1���1��@0clcC�p��E����3cŌ��P������,�1�"c#3F2�3��Y�t@�H�`���(5���f�2�p��@�,c7�f����!�cŃP0��i�c�!���c�o���[�2G�1�c��c��1��C)��چ��d1�3Xʤ�$f�L�P��1��Lde��!�c��=��%�c���[ cc���kH�`�f���3���q:�#(cK�2�d�P�a��P?1��[�2X�1�z!�C�deb�F3ȳ�e?X�1�c��1��1�h�C$c�f�1�c)�c~icX��P�bgC���2�/1�Ǣ�?J`��c.�c(f�I#d1�e�~~�e1�`�i1��X�?31��1������5���&!�c�1�P�c�h�>C̤�2F11i�k�4c �V1�e�a�#-�c(bJ3�!��A�cˁ��Q�ge�c�2�1�����c��8c�&1�c�c�k�΅� �c;I��+�"a!��� ����B�&I<���*����6��
#I���e��@�	�c͕C c���I�t��3�3�1���2���P�ɐ1�r��b�. c�h�Q�%�b���C:�8ѐ3
�C�:Lc3!1�e|�c(� ��i�f���2�;Lcd�1�6��F2�)�c6�����H�1�PƓ �1��0⁃��3dc6�����c0f�c,c*�0c��z�"��{<PJF�4�3U��X�"�+�4��Ú�	�&`��@�(�L����Ii1�@�� �3�J�JHI�c$|��0ðcB7�A���U�.ˤ�f�-�&R��bV1��1�eP�1��Lg��ih�@ڲ�1�c&>(�Z���U��nZ�R�E��A�B��1�$�c�i#0X1��_�c43	%��H�����e�Yz1�I�I�3�+�p˥�0fj��29@�f�*�1�n�i�Sƥf�?R�c'�P��r��=Lg*%�d�4e���1���g@�cSĔ��	��ܙ �H�H�c t��3<��)�fSʅd�c��1��t��H�v���7�#2<�1�ɐ3�
�A�1�gG�drg1�	��F1��1��3�1e���1�z!�c*��2�1�!����2�?$�1�e�cE�1�e���,"�3c$�n������ַ�f-�X���2Ҳ�,��c�(ckN	�)�c�ь`��cCZ1�1��1�c��1�Ɛ�1�S#�1�c&p� �Pǉ�1����1��e�S�p�!�$��c��h�4�c�c��c�6��?1���3�1�z���	�c4f��$����c�8~�1�;L��c��(������8c8t��Yä� ��d5�1��L�1�1�f�c8��Ĕ�c�sHdb��1�f�� �251�1��L�1�ɜH���� �Y�!)�0f�dn�4�Lf���1�SՐ@�dXǩ�1���2�@�($d�S0g%�3G��1��$���,eҡ�!�� p�������&q#.�=LgՐ[8ᵰqmI4���i���@�$bc�1��#^c�<�1��Lc�3И�1��L��P�/1�ጴ��C��1���K�lҵ2a*��n,d�ܧi0�wfqri��$�hb�H�d�%�F0�R+̯Q$���3�g�l�	1�c(�Hev��9�a#�ez�c(~g�.3��4Lfx�G1~�	e�+��b��|��gp�V2̱b�ь���&�aD�E?q$`&K8��C�#�3��Sc8v�Q$	-��&*!�QGc��frc8��yc&R$e�F2F;,�cX@�I�c&i#�(c�3
�1�(c,|��Q*c��2�`��d�`�=L��qfRf1�e���洂�eVb7��4c��jH�	�c9� g$�2D�31�KH΄�$��c$�Rf��!�c@��*��2�k�g�kd�i{1�2�1�e�K��f8��#�&1�ţ�1�D1�@�l&3�����c��RLcc1��@��K��)�qEc�8���X�i���a,c0f�d1�I#fc Lьc$�ip�"��0c��1��1��9�3�`΢IC�0cT1�1��X�1�g�1�clc�)�6��h�M1���-�`���2���1�c��1�1���1�d��c�Lc�`?cC�c�2��`�A��@�2����!�!������g�c9�e�a�1�a�1�e�C0c%�3D2�e�Id�Ilc,�1�JTql�(`�̒�(E���3X��(�B�1�%�22EĖ1�q�[P�iw�d��i-�3��$g���/�i�2&		c)�D��Fk4�H��c�^��e�e#%���.�W4��~�$�ML��dYC1�~EzE�!�d��[(���
5�v�N�1��;SфiP�1�C0���d���fic���G�QD2δΤ��1�p��3tC4�%�a(�1��^1��8f�2Y��I�?qD`&1�It3�0���3��L���f��^�G�B$^`��j!�QG?2F>Le[^Cɔ�F⑃$mYe���1қ�6��LZ�<�jݡ�Qj�+�thSy��Cg�FP�	�W��g]z,gј`�U�yBI���|<���-}�"-�n��۟�/ؾ+���w�\���͋>��,��ʻ2��s;:�cn*��;7��\g�F��m�T�.�"&?�Җ*�����ٺ��kU��K�˜��Q2lwarR��y�+�r�=s�{f��ڭUU5Nb�t�T�(�ySY�Ef*��SxUQ�)Z���ƽgw�,s7k<p��%�VyE9*=����d�^]L�NL�ҭ]V-J�fl�xEwou(PTt�uf��.3g�-�eÙnr�)u�bV�'�6栙&*�L�w�ӕ3��#m���r�^�Q�3sWp�v�"r�_L�VdV�32�W3�ɋ�_RMڟ#"�V']34�s"
�_)ߔ�����\�������y����>����un��1�R\t��ӳ�W��T�哓��k�ILʗ��*L���Q/'��$�>X�Bز�ܯ_��t��仼�������鏟�iѳ�0�AQ7�*�ʨ�YkveI�U(s�T�ή����0�/���TA&f��w3I��j+�|��5�s���
��?+]XN|��9�˄�S��WUZy��wzfWn)�D�g%nt����ex�o2����
���'��*Ws������~�输�
�۹D��ɉ[DUnj�4^�ݍ�b���/�ͨ"1/��k�뭧5��T���~22�q:J�f;r}Z���٩���9��V*��2�~��W�mMl�[�)�Ғ߾>��]As[����9M�|!������<g�m�;�V��/Ԣ�)[/'Tg\�)�L�ZY�~]�����q��/L���qB������w��0�fܹ�:{t�E��Q��VL/�e]r�Q��q\�;�Y�ړ��Ye_'�t��H�*+r�)�өfL��}D�Z�Q��,��94r�Dnb�͵v�nЧ�RW�u2mu�Xe}*,��DS�H�!Ye,���2nmB�^�Y��T�1�%�y�+����I1=Qh�;c:�r�q�՗8�e��8�UV橷�K!GQu}_����D�׻��z���ߦ�T�tUl��Դ�nn�}�/�.xz�����;!����/�ާ�/{�c�3W�#���(��.��S��Qn�v�Q��;�\�������V3)��ߚ���K"��Sh܎�K�rz����o*;g�ꖨ\��ȵg��u��%Ő��'~˽TF���3=dʎ�&+ۜ�}�(�Yp�S�!D���Ó*�+�[*>߳w��t���Kw&H�s���&�V-շ:"�L���vn*�Q��P�UV�|�V�%U����޸��GEΨ�Բ쬵ʕ�B�T�e�.�ԖdA����Z�{]����Z]��.[���=�<���սJ.>n��(�(����I-7�����u����b[���ϩ�3|�m(k��3�2RM<�)8���2.L�r��e�{
�OtV��.ɴ�=�2K�W�X���)(��if�%9)Z�O9n�뵞�F�)������2;������qs��jʛ[�8�.qg_Z�j�7q��~��,�/t����*�&�k&S�*҅)S�!Rν˺_l���U�Ű��l���wO?v�v�{C|�{�N�����G%���E�F�Q�2e�Zw�#^��~~���f��|���z�O��K�=+k����U�VJ��ff�.�i5v��N��T�U�N�܉2*kv�*�d��t�E*.�*��2f�IDR�u�)ڟ�S��.��a��^%�|��֜��&�1��R�N)�����]�;0�'c잛T��ۍ�P$F����y������%�u�{ʖ��.):�ڍ�Ժ�E5;v\�a94��2��j��S�y�����Ot4<~7�������{�^u	�=�{3��q����o�3Ko�?�������y_h��U~�}��/#������uws�˞��cp����g.�qΦ��z��w�s{s�srE+S�1nvzyj��Lr�3흸M8��UVMc��'2h�ĕQ�5ieLnk�Ź=.jzgfZ�~�H䣦�E�V�b���j�'��T}[?F_^���5�?q:vvb6ʔ��&�qݳ�F+U/�Z���d�T�6g�R����8��Q�s�,��YWY(ٌ��W��Vf�V����t��;�	�UҢ�f�m=ɢ"2o6zȵx�R�T��S��ݺ])%��Z��g%�皡WT�d�d�r��/UD��ģn��,�����T�zV���D���ww>�:断��ٙ�����`{ʷgdB�ͥo>K��LS�է�mг������}��!$��}6���Si�=�gd������%�J�)k�R�j��E@�$�..�"TS�K2eN��ӊ3�1}4��o}�=�������%�ͩX�ev�	Fg]���|�nͶ�"w?�vy��^����7ճ����*m�-�p�ڕ���Q�r��&�d2�m�s��s	�3��^L���qSX�6RX��Ienb����>S�zQ�ǝ�⿏���Ov�w�_e�S]<�z��[��l��(O��#��7�f����{^�iȥ�*d���xﳷ��S��q;���'D�ߵ-���U&}S��i�Wt��̩���ێ��>;���~@�S.liџ_�~����\^��~	�/�>�h���~�f��~~*��#�qG����z���'�x��?o�]��o�}�w��R�����|~=����oz���{��R�c(�=�T@Eۇ���7�{������>?����c|�=|5/Cξ��զ�����T%�ce�[����\����7z�=}q���~h|��S>1�-�x'\�~�!竟�}<��s�M��?��*xx��e�Ov~>���ǳ�K�\{�)��O�rwk�ӯ�]�q��$�Ŏ�U)R��St������:@,���ߟzzc{�2_W���t����rxc�{��5��x'�t��y5<�ƞ�ZW���仳j����S��&ZS3�%ΩT�n��
��J4�Q�w�h�X�5Ij,��<z?�?��x{����S��f�;��n��|�����{�~Ow2��m�s���ϾMP�l��N����{W�zuK߶�5T�s���.��ݕ��ێȪY�if-�W�i����]��U�je'�=|"'������gY�_6�����6���{�}�l�m��l���~6�>�y�#�{v��w*�Ne��1L�TE(��_t�O՗ݶTk���{Z]mt��%c^#\duww������������zm��j���S����W?:#!}5+-]UN*��mm�u���{f��JU�d�D���q���t(�,�\�L��7;-b�"�u0������1h�*tf�v�3n����J���S���~}�ֈ�~��]5�ȡe��QE�9Y2�_�c��6fU��d������U
T5�Ss3��˝�:P�R�J���7�K���d�?��5���<c�j..dg��r.��Q/��뻟�����N��9�.K��O��7����[գ?�c*�)�N�?LQ:{*aBș��ٻS=�F^��~|�z�c|�_��e_��nF�|������ޝq�0�k^߄OD�|�_C�G�k�שg�|_�.�Sϗ�Oo��/s����f� :>����}.�h{꽝����S{�/���������y�ԕ���쩘�s�镫S\lbs_�گ���t�v���}}])��i��T�D�ji�2�{�ݷo�˶�u��cT��ϧ-����":�eb�r�k�ov������_��?vV{}U?�������}~g����=n��K-���ޯ��M����O��7�t�gk-e�u|W�q��__H~|ޟc�[�UG�~_;���T�Ǉ�޸�}ӕ}���Ծ +|�����=<?�T��F����}����?��{��Nũ�xE�ʪF^-��R�=Q�����/=��6�U%d�[J��k�P�S�'�rtjܖ��]�Jق�Նĵ�k�{�Cݫ��f}��R��w���m�����k��4�r���_O�Wp�S�X_R��-�ݬr�ֳf�}��������K˷����W+����2����ŕ�!��������˻�.���*T��DdrX�WYp�q)����\wW+�K)*�[9<�wtҜŊ��Jn���T���].�.�uI9�5wשg�:��3�ĔLGۦ�ܔ�ϕ��|��S��RJ2#5ui�w���z��y*#�.���Rnzn1l��IЖq_W�Ɉ[��u����G��#x���UX���ڣ
_��KPZ�J�yU�Et]e��fCs��X�����е-j����}���۳W�xA�
�D��b����h��&�yo|�<�.��s��?\��ח���lHM��^�����@��\�M���9c��M��V�,Q��b�x��,�'��L2`�Q��ɧv�{R�R�mR�*�ļ��Ba����ǒp��[������y<&�ez�umgq��m��9��^���-�����qm�$�BF�r��ض˩K654�����a�ffJI�,�԰��]��*�ݍ�3������iM�2ʹv��'%9�
�3�4��V�)���w��L�-�!4%�4���W��13�
(M����I46/��;5%�թ��
0,�Ë'qY`s���t5-)t�5�X�
V��YP�5k,���!F1)�'p���dY6
Kmnk���i�9�Rb�c2��H�e�U&b��Q�4�S��NmgH��V�+i�u5�ɥ�>n氵�Y&�!X���)���U��[6���I�S3�m;f䷌�)�Ü�3Y��t�����5��s���^Lm��P����V��X��k���m+y$���NH�BjS�muۗbۍ�&W2�[���m(99�M~3�c�5�%��b����.~�t�2�^0ܪ�ڡ*b0ֳ%j�մ��Vi!�2Fh��6�Θe���˴�%�CI��IȒ^%�]��6 �Bk*+3��<)�Q�Ē@�IkF.nMjGU�I�^KI�9`W7��
���]�e'���t���3��ylY���u��w�i�'0�׌�5*K,�@�efKk�Yo9��,�Mn��"bŐ%�2Nbb�ae��M۷loX6�`�s��4n��M�;��su���K5���6[ ���Ж��'8�������ռܩ]�����3Dnȑr$����a5j0��q�zy�'�+ڲ�plگ��vE��)�H��5�b�gnT���ph�ą�%)6�K-�	`�.�kYc	R-�"� f��
�����冚��]�`&�%�l<u[ɍ�	a�us[m������fs�ev�/^;2�f^k���-����3�Gl�l�p鹜����i-C�,��vci\$�1�6��s6�u��%�Ҍ2N�ݽ4��V�m��3ϳ4�m*y��a��b�^W��!m"im�2ڜ�o�d�k�Z6�b�xp�
6�5̎�P�����[�����A����z�\c-����R�30}����V7ɪ#s�]e�"]�]]±e��k�R�fε��5Ү�k�L�����	����;�cR�㔁�қ�b]�,�E�XT��4CgJ�c�&`�̤1W�k�<�o������	�A��Hu3yFN��  �&��M���ڧ���aD*QJ����l���8��?���pI�U"T*,�"2P*0�Ȳ����>���A��E/���������6��z��m��6�or�n�m�nm����m�cm���m���m����cn]�ܶ�x��m�nq�m��cm��lm��n���6ۦ�v�r�m�m�m�m�m�޵�	�H �� $#"�Ƞ# ���P$A���QT�!��R �	Y!RXx�#�G���y/{�xۖ�n�n�m�m�m�m����m��xۖ޷�ݶ�6ۦ�v�r�m�m��cm���m���m������7�f6ۦ�v�r�m�m�m��UN�m���m���m��6�۶������ITAD���*E
0%�,�`T��"kD�kI&��m���m���m���m��-�-��6��z��m��6�m�p��v�t�r�m�nm����m�cm�޷�ݶ�6���i��o[��m�nm�������m��6�m����wwwk�����\ֵ��kI5��5"H(DB�Cх@�%d�`�1���+:�E5j$X)��"���1��a�U@Y�,4ºd�R'�̬E,*E���(��L
h!*Q	T�E4�^|G�
"�	$�I	��z}��X�S7����t��-O_�?�ط�Z-kZ�Z�Yf1�c�1��#�,��4cC(c4�$�c�P�@�4�M4���`�2��2�H�1�fc1���a#�1�e�h�8�8��C8b�`�2D1�d���3X�3�F�,�Ϟ-KZ�|������2�1���c$�I�1���c0��e��e�1��e��Զ�kZ�Z��Z�P����2i%��1�c�0a8b�X�p�q�h�8�Y�IC�2��1�2�3i�8c(g"�,��Y��)kx�^-�kZ�ҫ����9?��{�Դ�b��uۻ��%�^f���3��]vGYlʵ�h��3B�42Z+"K�זn#��ƴ#w06+l��ݝ[�lx3�5�UŦ�[)`ƫykK������:���Sik�Q��VV�]��aq��m���e�w����]����)-��k�q�]�׳텱��0�E5��X�(�i�N��K�ð��n��Zs�͡Rvh3Xf#f����؆ܥ��\���me�˕b�"E�ЮJ��&&)������fS^1RR����Y�K-��G1ҍ�6гL[�hK��͈�[=���=�����w���ic�f(��^n&d6�.&u�֯�+km�Y��s��b�r%��+��m�gXG:�+6�&˶]%E�5&[��bn8NV��]�ڷ��#ʍ8��5��.�%�f�u�\��i.ٹ�����mE"�ɣF`�W����
Q��	ex�L6TZ�Ֆ�<lE�ʹj�ј�]MF9F]E���6�W��,UuR�hM�ԤnT����P�"�8�e�6c�V8&����G8^�q(�q����KA[Z��*,�e���B���7�;;�-6�[
X�	LhM�1t��м�m�]�c,([^4��n Ms�P4! f5�5)6�l<�����9�	߼��|ˊ�h���ڊ�s:��RRHk*Ė*U�BQŤ�Ů�(����˥���Y�і7�s#�%�����8&	�q�E+��6[�(�pך���@��a�T�|�G���v�V��y���ٌ13Z�fKKY���6���[��1tc3mV�b��8q�̽/yd`�5�j˸Cjݮr1.؆J���Hm��w���E�um"���*%�����kk(��te��6�!��:b�7.�V�r��ҥ�]�2QmZ�( a-%�Rr�@�P1�0�k�RgC;2Sk�fQ�f]IPcK�R�-�x��3b�)��9���Y1l%��`xۣ���m�L\�s6�[���5ԭn��6��pMx���c,
��m9�6`��f+I]�\@i�o*�P�*�h	-Q�Z�(F���N5W,38��3��7m��d�R�քt��gL���J��U4��i��k�m��2K��[�.�7�̫�[p�]�0��aa6���k2��]�)l��g�u�T��k]&h��-�1�.&!Y0��6Ûh�$��i�*�c6�����t���n&vi�zg�ۍ����6�7�m������{ǽ���fg32��������~�kGٙ���˻���������h��)��:�8�\i��3����h� eg����2ZY}+��cfdX�EVQM�vFW
�GB���\�LL�,Ք�][��V]j�Ynx�j۲�k1���x����74I�j����nbEm�P����$5f��	`\�Cux�S�����r:�i���4�M�iq\eV�4�3����1��f�j�M��B�1t�[l�流n�γRі%��i6��u
�R	��	v��W��sk6�͎��BWg:�%kSj�#���0�4��]6�@9�d�R���7�-�,i[*@����R��US��/#)VؤYk���+;mI���J��a���A�ɐ�-�Ű0Ho��i\�{��ֺ���ó'��s3ó�����X�� nl�SP�=JhԌ�lm
Y�(|M����ٯ���ѥ�ݶ����xFŦᇥ<DCyv[��\m�g��b��c4���{FZ[:eu+tzt��F4P=߷�E}�i��zi2�
}~�!g>8�L?`�8fgc�Ӆ٣!��8��ᇝQg�ߑ��4����b,�ꙎoP�IbQ�X���f&偭��وIg4iF�"ja�u3T���E����&�bܐ'�Io~��'���{h�¢���T��l���2��D�)�nԳQn[��Q�/�z�
(*��`�7�c�l)K*sF-�gD8�bA��0��Ù��1(���c�iƌc8�L��`�rֵ���#׍��$��ZnUS��:P`�T�6���Qr�����\��K������0�ҍ�K��&�-T��Y�C8P�4�g��M����a��76)�Xg%8f�Nm��O֮��=����9g��w��JlÆM{8��l�o+M��Q��'�τ�=!�5o�8ڹt�T��p𸩱��x�6af����Z�s�Dxl�;,�~�觇z<{<�^���Fh�q��1�����c4f��44G(ޚ�.j��7[�U
Y)��jӽ�ň���r_����x!�LN��Y;���b�+�U�6��h��m�ڶخ�#<����Y<��I��Z]M,����觓G��Úfi,#�,葵el&�9/m�2�0����+�qL����z"c�6�:t�r�nO�k�%>׈.ᣌђ}1L,};�f�OJ-�c�8��Yn���[�Z����Y	٣=@�y*�*0�&��;5ZRv%��Qj�wz���7`P&����EFs�ok�k��>E��R��ct���j.!��l�k�]er�ٶ���0�ءP�LG����e��*��T������l��1��]�.U�ǎ�%2��
L]�ZKh��	.��5��L�f�GçL548|s��hN��V��|,�������q\)��Bat'C�̃	��6�ڛ�Y��N���<�,��	�>�p��Jk����6/ΈXS@�OF��`�)����i���]���v��G{&ί���<�[q,��1#��t�;��)��o���ɡ=7���&��c1�:'�PY�(>�BN>8��i�`�8f-n�k[�|�=x��浦�I|��������I��<�l�2��'Ӆ���x�����r���0̭�z=6��<rf��E>��aщ��z�����l�d���)V`���j���MK/ݔ��3�X|V4;IE4]�kR�<)���f=ِ��g�J{��DeTD/`�d��ň�c(?3O��4��1�A�0c8f�f��Q"�[$��I$�_	���:tѿ�{�ish���{$�`���&ÿ:�NΈ!�gL9։+}Ŧ���b}��6zS��������Ĳ��;;]���n�k3Y]]%\6y>�t��)0��
(��Y�iD�tԫ���c v�8Czh/�ÂM@�:����ẹ[�i�A��"�Q��NwD��U3P����5�z�>��S���խ��i��� �1�3F3Fa �(�b\�{&�K�\L��rI F��RhtI�����.���R�L8|�}����f�J�U2�\\��T%� �`l�Hf����A�	�a��ҚLܡOL�ٞ�Xk�Ȧ(a�ن�~_��)$6X�#n�)�g��犛�:����飆I�����t�XzFX�w�⽙Ca�9�Ӑ�}m4��JL$�!,����f�<]�80�����ƚ`�1�A�0c8f�aő!4џ���?e�X����@�����gKfGf���,�,�U��m&v�/MM��u�I�l�gV�<�lh�[�֮H]pu[4�C�b;���M2�&qYY,�:�� ���z���]�%kn���c���6��R��)��i�NZqi�&è�	mԶ,��9ف��źY?�d����;���|[��qRA��Z?P��(�#ޒI8�3<�u���/r���I��c�-!�rjj�������j�ڪ%�OO����4`dd��|4tàG����^;�\���}�ᆈ�BC0cp<�杜�e��ԇ�)� �R3ie&㦤����>���M�t��R@<)M2%=PG��*��>˜̕�iE/z�� $���|q��|1����4�62&K=�z��^ �c�;0М�'G�x'}�,V�^�H���A5}�uL��fӕ�]�h;�����3�_U�vl��6��^�y:��gqo5z�qTP`��Zr��8��J{ϡk��I	a��잿W��eX�ˢE�ʖ��IWc�ֶ0�sa(2l��I8u�P`��Bg��n&^f-ɳx/C�&l=:�d���tp��Fa<6a҅��M�9;�̩���xznE�>4���*����b����"�V1]b��6���+���+coX�b�mX����z�&>cn�X�|V&1X���c�ݥ��]WW����1��+1�b�LO��X���c��~~W��W��~~S���)X�c�V#�����֫Z�'�kVֳv�&+��c��T�OX��S�)��h�c�>SlTb�bF+�S�b�b�11M��f+��LV1]Kb��7�W�V%�����+�b�c�Ǫ�X�6�=W�U���j�+V�lR&$eLU1X�z�3sSV'�RD��5����c�S��b��m��x�X��1�xʘ�Z�M�1T��S�+�Lq�۬~x�m��1X�������T�b��1�<��'��cLV'�W�V'�Sh��z����:��z�M�$LH����?7�?8��Ƒ����6IT�~�#�S������̹0KJ���Dm(7vfl�$F�q��"&d��.�Ve)��]YyX�X�Jy��j7:�Ơ^_K�W��Y��c�<���h�ÌNc�}�	L�p̋�XF���C��r±=0�H�6f!�f�0�����D�^X� p9V� ��9�W$�3;<��:Kܿ7�ٮ���ħ�P����^��w�ϣ{�x��:}�ߣ�m�n��ٓG�dg�}���}���ٝ�y��}�Z������ffy���}��}��kG����bַ]q�c�l|�8fa��$ ��,�E�DA�SG�f�SM��k[�)�Pz�'O��t�n;_N�!�2Dd��Є:l��H К?|ے3E	�@����.����I�%��Z�߆�:RD@��(��P���$�CFA���P
&�͘L�L�@���a~�˓l��y�v�ya6��#i�8���v3Z�i�_�*�=�'����?+���"�,fY#6P�BDCr��P?j)��k���� �kT#d����P�p��$��u�~_@�? �w����n9�>��0@�p��L�Y"2~Sh�MD�����$В
m'�����.���8k�l���!C�@�!H-4��vkZ��Ix���)(ךiǇ������u���ַ]mn��\c�X��z��5��Uh� �����QP`Â�`��� ᣕ=�\��l����SZy��}�h�Zn�iz#!ѐ�0
�HhI��4Y�d������n�M[m�8�;G8�p�̈�9�sm@�}�'��x����$��C/�&�3e&�M�[0(�����5),a�I���[���ھ�\����~��ఇ�2d���6��oOU�#J!�#Z����c�_s���A��=(K��� ���tCd�G�BJ&����/xn�!D��w����<�jGֵ�J��x��Z#��8����9�JMYh�a@�0(��쌓��̠��S��Z��x j2#$�	���u4�jSKu��Ě-����Q�8��:��u��b��0gÌ8���Yd��-R���U�e���[��M�����}�٪�|���l����1١�<�nwp���/u�2f��sn��Rͳn����]ooבx���Q�eAb�:�"�;^"X��,l��[�W1q�6e��Қ���S)˩uį�.�hb���Cam�"?4� ��;St�C%��ZmV�r���֘�U,�e㉮(˲M��/!�s�q7&�6����*M0>?	���;O4'(�(�A�,�"��P��� �<��R��[�qBB|y����<>
t�ACT�h��Q5�֏[P�JX
O�S�V-����A�A� �8'�S�C �dȓA�0�%z�haʻ0'����M�~J��,����E4#F��!N�#8C@H	J>�I�JD40;����~8l�~����1�Ziִf���՘�'�p�$��}h�MX>V��#M�V�s6�~H�KwN˚2����.�/m|�;���fL��3�d� x$��(�5��I�!�}|.a�����/�JQ{5+Zޣ��m��´�>�M�><�ݓf�)�2 ��̝8���~u���ŭ�>c[�Ç�ω�M�0UnQiJ:�(�2B�)�O�Hd@�05�I!�)�"�ؔBx$�y�ʩ�g�,��O"���0B�P"�<ւ	�Mm���[�F&�z!�$��mD�L�!��0�JK�Hg����ܒ$�I�>=(y;"2�b܁�!���
s�9�)nd�p:!D�d����)�D�2D`pdD��0`hHh9d( o9݈R���%���[�jΙ�Mt��y�ۭ*;�#�����$(��A��|&���ؘ$�<�
&��	"L>=2bC�{����2�5&��&�y��R 2l'�P�^��5�ֶV�5�i�m�����麨�]���GM�5�J&�Z�B�ZTqGϟ����\qű�b��1���z��R�6S�>��e<�E���y5���q4��5�cq=4o��q�]��5MS�BN	�DF�kIiZz�k��0"��֘��o���Aȹ1r`��31�R6����d���s��ل��>��Zj��w�S�<#VѪ��i�k��(�d>)�͚�>C$'>�?'럁���#f���Z`i-�f7��m{�k�2�ژ���ѩ�ʓ�8 �������_��v$��C��c�)�@,�ƞ��6�f��!~�>܍�T�]B'��"���D�M��L9`�O:-����S���H!�&D1&OJfId4���S[G�~���ּG�Oy�o�����G�ʣ<�w��&�ޢ��E��S[F���O͞i��DF�����~|ul~?:�??1�Z���1�=u��g��R�6S
"�_1�"(���˅cJ(��TEXȪ\,S�
v�E ��&����!��������������@�kn(�JRkV��Z���5i�RH�CXP��5 D6	�t#?��@�6�R��.�e�w��c�q�D�m�̱�2�M�h�?{$�����)46�,df�LCbDiU���C�q��{�_�Ӛ֍�I��)D6:�k^~�J��"���Z�� C�S�쳂L��`q�@ݪDG��6zMkh�>�qF���${a؜О��	�/���j4[M^��iȕ�eJ��!�ָ�M���G#��m4�4��PxF�PZ�"s_6m43�~��W�:�P�42
^Ӎ���jjYֶ݊��sP��kP�	hx V2H�	4Y0��Ì~~~u�b��-lx��=u�|H� ��$\Y1�"ꍳͬ�1v��$u�V�%�,��3C7";�sr����y�n�������\ǗH:Ta[0��5v�6��leq�9��.%�ni��z@��Bs�6��M�� �,ơ\�Ie2sp��W].��:�\��kM�k�d�䵵�Ð\�:�$����{,���-�k�h�Ҕu�Ӏz$�O����C犪MQDj5��4��U���Nu �p�"Q�~|1�s��М:P�D�DD&�6'ޖ�7ND�%$3��Y��BzN�'����?	�:��pe��"t�JFa|5d</���N�0!Ss�����ܐ�!���Oٕ��0����tß0K!�������ᲁ�N�{2����S�1^�i�<��	�#��"-4����M>֌�6�u92�MO���`﹝�:��j��;�bKnжi�8�y4��;��������䧰�,	���(�A$�bLT
2Q>���`�O2��\78x�h�R��z��?-����[���b���νch�)���r;����Xj���0���=��? �(r����a4 �!�����i��j����a80臾��HsE0I�<��?=<�6�ߋd�r�]�����Hx��Y��~��k<�x�rI�:��6!b7��Xv!��E� Ѕ����0C{ؿ\�����:!��D��BE5��D���� �k�i4~$�"$��M��!8��d�5" �O3��0��\��kF]L�0�8�#wN��ֈ�+ɐ58XO~_�FI�8$�C�%&	O ��I�la0I����n�\����nl�|)<D�` Pd
0/F�5� ~O0�`t��y[����8�H������Hz��+C�iN�>~~[���8�ַ�-lq�1lm�νa�R�0ٓ��V��zEd0Ԥ��40Ї�a������V����xh�F� �$�		����t0�a�3�u����!�L�F��M!��pLpNC��
�?O�&N}��m��ңt�@-l��2f�u����%�jG�Cе�iu!���y��C�O��	g!MM�؀Q�n�tM!��l����a�$К�~�sżOB�p�<=4 �����hN&�Y&FMD�t��Ȇ��2�C3ص<�&����
0�l&	F���!��_����(�jh�뿙�ߟ5I�A4P����:���d�3����C�c�:�~u�bֶ-lq�ulS��z��Jz���
�Ne3'S�Ed�zd�Cȕ40�5�.l��}d�,�e�b��H,P�5�Ω�1����5��H�E�s^ ͉��0�k�Ҿk)���SD�.e��ݰ��<K�b=���BM�˗2
��h������<���h���"��#���4Ya�aC##���O68��s�J��u��~[2j�?@��I��&����1H\j�j��澉'��0aD�
f�Bʆ�֘�1��j=C��?#�շ$��#��M�Ԥ�C�V�Ĥ%�|j:�7?~2N���ɒlIy���[�����&�(�:��&�(��	�lL�+ٻM���["fdV&ұ%�2%?���%?=o�c��-X�V'�1X��Չ�W�b��c巏��
����=o�q]c�x�LS�+1�Z�j�kn֫N�X�����V:��X�X�c�6��+���+c~1^1X�a�u���+Ӯ+i��-j�����V6�b�Lo�uXF1V��O�S�nLq��N�Ӊ�T��*���LO���LF>V&1]b��Ɍnخ6�1\c���++Ǌ��+$�c�V1T�naX�^�S�>n��b��M�&&)X��8�������)�t0����(����;�6S�LTb�-���#ת���1�&%�\Jb�)-6��7��V1\b���E�ݭV�c���nR�1X�c1�X�m^�X��b1�b�8�:�b15����KDGS�z�$G�Tb�����*ǳ�?���ʩ~?��H{����Fe�y]�{kg����@�C��������޳v�ր�x����ԥ��1�[��1����/��.TL����y�n�O��F�u��&VLb*�ڹj;��!_)ص��`�U�|{C{m�7����͇�S�Ӫ������ӷv�݄�N�ww:�%�0�CQ������!dEL��˒wrJ��P�uwT�ysjP�-�SR䐕��6B$j��S�Qa^��2
�9m��Yq�E9��d�JQr�)���
򫻔���w��;��������1u���y�=&{k+�ݫl	�~/C6�M�����x^�g]��:K�d�Y1|�r&��`"~����ͫ�B�K�xٻ��R~�y��Ͳ:4u�����_-m,,vInu�h+U��f����@���B=�e1�C��O;�δ�zbު̨U��4��Ģg�𺫙�˽� �����e^��q�h[:6�3y1��?3�b�)A�f�Y�y���|����ɮU�ҋ��U)�BՏ���E�(����l����'�K���V*�	~�����;P9�!ml�C�����b۰:jShExF�
�e6�p�@�@�Lkh��7r�\�����J:iR�]��Z�pʬ�����̗K���\�<�6�87���--��a���t�����
с2��%����	�m��K�uܡ��9Ii��9ؙ��[0�"Ɏ9�YIMpj�S��Mi���sL̪�Q��8�/���_}��}�;߾̯{3>���r�o��W�fQ���ﾯ���m��n��2��
|�c�b�u����-�1�a�3,d��$�O��c�S>��]e�ҙ�1�n���yT`:	�f��!�[]�q�Xbkj�@���Y.,2lRh�Z�d��&���.�6u�6���(V���R�v�f4t5�v&���[]�,�\���b�p�Ǜ��(���V����i�K�х��K`�D���"�Z��ɵ�Kq��9��nl�ܺ�-���!jm
,l���Ү�X�x`�%6�4YF��ҥ�:�[y���ظYCm�04��	�BN�vůF]5#�iJ�k(�	��4�5#6.4��5�c��B�Fm�dgdꛬ�lD\ݑ/���'�{	��L)�+u�0�!A��iKcg��k_{u5=�ک��l�)JsѤ�AH`�M�ge?�C����%:F"y<I6�z�[��^�X�u�1�i�i�A��՘'�m9Q��i�L
~���[q�߷��v��d:0��&�K;��������[o���Fjk���4���B���9�3�	`{,@A4oT�&��I�m���hB�{?�,�5����I���zǻ9����,[�yj���hI��#�b�%8�O�M=~M��C��k�m�R#"��?3#�4���G�V��[ך�ׯ�Ÿ��:�1k[���1�c|��m��^6�/����$jZ�=���4'}��؟���X��k�F)m��23�,���g
d0lJ'�	�Ci��l���x���"b�DU>��\�msʕuj�����z`&֓BB�㥄؇i#��[��*hwZ⇈Bքrz�xl��-sA�=<��BBBO}~�eBY�iq)e�É�2Ul u��5$�u�K��#��e�r�4rC�=d�C�Mn5H~�<&�h<�q�֔��}��?&���Qw���`��Ș4�wZA�6��(�jh��רz!������$)�8��T��s.aJ���zad��(���8�Qk\E���-���\q�k[���1�c|��m��^6��+���R �&���2YÅ0C�b;as)��&D<C�Sc't6�0"�kP�kX��h\nmO��m)��hO�6N�h���L9)O�����ld2'������i@���6��v�Yw����h֡aV]��|,��L��8Y�2'���4��""�s���-��ԓ�
	6%�i��7�'�Z9�Ґf�/R+ZxB�R�p�zbۙ���Lğ����d6" a�,:'��ŷ�z[��C��6h���nD��)f���N����u�n��������0��z�h�=z�;_7�5&�=߼�R ��(��ߙ�i��Z�8��ڶ�f��D(!��$92Fgƺ��g�k%p H��(S����3U���I�l����0�ó@�c�Җİ���;��NQ��u�=���!�0���C�.��d٨~\6u(
2���`�)������,6�$���3k��5D/P�����-��6ɮ<Q�8�S9�n�H�!JS�]4��M�23
�ć�$���񅹙r~�gd臒`�0>M�Ah���h�u:!�����Z)�:��1�n������-��>>h�4�Ae�KL]*:J�;a7f�M����ʤ����o;��R+:�=�6̩.J�ih[����\�wN^����~�����w��:��5��s�]�y��8!�5H�a"�0��5��jͱ��2U��
�x���'		�%<��n�M/)uH��v��j
[��i���e�a*�,qAP.�&�њ\5�sͯ t�Rzyf�X�"�k=[��JD�5����Z�M:�"5H�ٯQ��=��BM���OD���iz��))�xCsLBsZ��;R�:vM	�a������͈pC][3��}���C?����Zt�<^��2kS���׏f���1�Q���A�pþ�T]}���/@���B�C��5浭B/$�m�=l�����C��[`���f������̃��i�=��>����i���pC`��AZ8D���URj���_iO���=S�~c��q�-kuվZض0���h�6l���	Y" �b�aP�Y ��A�E"'������X��~�㍜!5ͮb�{#�z#4�,/�4��[�A��*?L8a����a��4\��p��#�4a��S'�<
zOW��<��=��p�v��n`�-�=�Cg�^��sSM�O��N�:�n)BBO߿ӵ���RB�V�S]e�̬��Qa�1��iu��=ﰜ)�k'���)�/��nd�k���e$u��Kӈ���eS*	!J����4�t6��:��������Z�uo��,���,�DA�Agr��$$D�P�t�/y6~����f\��լ�\<�z��St�;LJ��-��B���`u�q(,I�������?�����-�;�B�4X0�
���*ۜ5�cn|}8`&��0��h��&���Rl�7�g`��p���ɓ5q���9?z�-��f\���:�L�m�|���y#+���y����欁
!"=ݓ*'� A��ܛ?��ε)I�u��x��u��[�1�[��������[筩Jz�N��y-Uă�
)C�B���B����#��H \&\h�$�N�B!C�ʹ/�8j�+�-�.i���CXlġj]f76�*����O~�ψM>V�$�*��k������_%g��~��p�t՗���ͼ�T���^SH�lQTUUI��0�A�8|B������%V�����R �N���g)�!�Cr�(LA�򙟏G�RY�����z�5N�n��7����S�>~~Zַ�������[[�z��f͌�	��ڌ[)a�7�#����;׳']]�6hy��u��Ec�[��+\�s��v����$0X�a	`Ք���\
�+xjkj�w0����e���E�atb���Z\�	�BA��X��i�p��5e��m�Y�j���ʗ@q[F�Y�e�X���uʹ!�4����d���a�M'�����<^��ߓ�j�Ǯ����խx��5�s���Q�Z[��Р��.=]�<�6p��p��p(~�6��U��lҬ<���m�rN�0�z6�qC�Ţm���5����d��O�4��<I*�QE�W�$�~z�B-���)�}i���D�N�k�/����*e.����͙��	k\A
L�oN�a̜��~?�N��Ì`h�IO���s���a�C�Ҟ�qk~ZַXŭ�V������� �,��.)�Qg"ҙ��2�����O��d�t�d��� ����>T�x��OƧ����vl���'��^���zsK�����m�~�p����i���H������a��u�o��{������ �Bl���8_0@����)/O��UU&���L,�ɨ:��-�qb����fb(�ɣߧ���o��gDH�u�������W�knk��DE�?��><4Cx?lSB"a<�����&U:��bW�{�}���E#�����~}�O�����~|�������_��~?++�eLz�1X���X���+屿�l++�=cx���7ת���+�g$����]W]cv�m����S�q�������1X�X�11�ǌo�b�U8��ln��vKW��mo[��ݩ��c�X�<f�+V�uLG���T�8�b��Mbbuʓ�LTN&$L&'�V&&&>f�+�V'�{��Ǫ�+��Jc�oW���bc�V1X�11����1_6��[V>U1X��M�ب����+�jیo��b���#h��~DO�������,���o�$�^�2�+����lsr��U&6��c�U�_��mm��i����?6���bd���ŭ�6ڱ11�bc�|�1:�:��1��=LM�Z���OU���bb���~J��LZ��/��U�%>�Jb���n�e/D��r�>��JJ���h�9z=��N/�v�:��ձR�$@$���mg��wU��1;v�<�Y$�\�đ���Y�:.Wl�N��Ȼ7"1jQU��L���Q2s������Ǟ����ޅ��������t�f�����o����d-��7X^g��JP��翐�v�ߜ������n~�33��略�6�|۟����>��m��ܻ�����|���1�Z��Ŝp�h�τ3ad�A�Adn`��"&�t|;?���g�MU5��s3��DDC�j2&ϡ��"&�, ��˷���Tr	��"'v�2�e5:=4!����'�	���3B�٪U���Qfʻf�g�}<E�Ľq�ԭ[���q�D}��k���+s�ĺ0��<��eM%� )!goƇ���n�O���yE59՝��3f���>�;Æ�W�>�������S��w�}��Z������ַX�1n�n-խ���|��)O^���o�9�*�s��������}t	>^L��i��? ?���BJF,i��D!4�����u��j�h��(��n��Tt��Lч>�+�=95?�q=�y pw�ս����q�����ؗ�q��ϥ-km�1zxp�O��4""h3'��x#�6청����D���f��G����2g���H����={��R�ʄ���&�DD��A0ɳ�䆽4t�O��8�ŭn��b�Z��[oL�� �,�.!��	��M�����f�6�k���!����BV˒�o��:CoT���}8���N@����˅6�xi���o!�������x]�Bˎ�S1�q�Lm�jqv-�R1v�m9�1�-���B��<���ʔL��J��ݦ�4֫���c,b`�l�����l�$��*q&u����ַ�ޚZ�4��ᡟ���\)��m%�tp����B"sP��ޗܰ��""zp>�.Fl�t}ß-6"#iOs^x��S=�7[�e}����oV��S�z�5����u��k�_�����q��5��*�l�G�vSR�͔�5����SZ�%J�ؘ7�1���և.�
�2�6�n&����ӟ/M�e�F����|}奝�a]�*Q0V�w�lqN=c�ZַX�1n�ku���X�,� ��:є�J��߻H��#n?j�ǎ>�i�5����'�A���|���S�w�k��F�w�Vަ��?<�qj � JiMq�B&�~�00�������5G����ـ�~>�C%Q�ݟ`���CSE4jO ~ײO4;)lHǏH{��*�����!�r��sHZ�$%I�ե&��V��Xy�~�q����B����`�9���T�}��2�'f*1$��4�&G�$�Gc�.!�M?y��fS�<��������=~[~Z���1խn�c>���AY
�&a)����EB��p��3G�G��G��I����H�X��4Y����O\�ԥ!��l��}r�#�C����t��լc���|��O8�B����5�5�,cˆ�64n�ۙ��	[����\�v}ω��6!��L0:S���>�����l8���N�1�$e�>�0�G&��X����Q�h��g�,8C��H'8"���*�Ǩc����i�I��jk_�➘�OS�-��k[�c�X�������z��)O^�޺�2,FA�)N��t~m�����lO
}�L6_Ȱ$y������[��҃���ی���\�C��ک&�>~�z����XF�␭\y����=�uu�����ٳF�L,��5��&χ�=f�hD/��n���7�u�f��D?5̭i�&�6��`��R�g-����Á����K̲}_~�8�l���TA�t���rq�pp��<(��γ�nˮ�%1�d��L<q��~~u�[��c�-n�kb-�޽mJS׫;?��
.�c]-���w-�Z,���Im�cʈ�0�P���h��ɗ���i���fD�������3b������pM���t���n��	],�iKmmk�3Y�K���� HBO<��v%���]�P�o�Jb5�J˪T�LVX�e.	�����,p����]K�>��BO��y���%��B�^-��~eTy7<��.��Ҳg�����;2r��}<?CG�rP�W��L�\,x�5��/�M0�Ja��&����ٯ}˙��ޔC���[�?�O	�����Ik�{���➢�bh�[4!�^�Ξ�b,t�4[�?v c[���RT��@T�@gm6t�ړZSfA������7�c�"��{�3��Y��I&��8��ku�c�-n�k1oV��jR��S.i�։jܨid�u�EC�)��a�����=DC�U\�U��Z�-~��I~�� vG���W��
J)2�MծkF��A)N��OK�0���f���4���)�'R�V߳^�h�!�����O��8����|�Űe�7 6⍳SnXd[��
��4�0�R�4=���>)Æhvnph�j4�>�	�7�C��wOuz��kA�/Kz�8!��e�e�ˣ99�L4xtَ���]b��1l[�V����M�0�)�e,5�4(��?nzh�uOԗ��~e6�}M�RH�n����D�t���ç�7~�R&�I��c�wi����8��I��<�@��&�r�Қ�l���$��ݶ��Ko��ZI��,�����l�Dw����0�%t�%<(��<0����Q��\���٣�h��G���\`��2GA��e�!B��+S�0A<���z������|�c���8��ֶ1�cź���=[׍�Jz�N�ҫ>���+3V��
��s�ECcMz{mB}�*H,B	 1Ж��ƒi��a!��}g�X(�*ė2ae�mxʼ2��Rⵕ�Z�;���\[��j�"޶��zq�� <I�Ԇ�1����i�� �i዆��M�4p�������3�;�]M�C��X���s�r*R�I����A��YG|Y�X�B/�V/?޼�o����ko_6�=i_k���s�%�Ǐ5��򖧯_=~mqk[m�ŭkz�k~coX�1�z�ec0c�,��(cC��4�F!�c���i��h��1�1�c,gC�`�2F1�cC�2�H�1�2Fp�q'q�c��P�`����1�3�q�#���0c�1�1�1�2�H��1�kZ-kR�mKZ�Zֵ��ֵ-kz���Ŗ��JYe��ԥ�Z-���1�]1��1o�)k[���z��`�2F1�c0��8�8��1�Zַ��)kZ���V��ֵ��qh��Գk-h��p������Q
EET��#�7Oq�ι�<I}�&l|���u_����6�<������ڎ�����_&�`��R7k�b7MÑYd�*��y�0+W[��98����fI�j�$�* ��jE�E�S�������r�o/{�]���O���T��	��}��&���f'}.s�qV"V\_�W�n����I�Ir��|��v���a����Χ|�:m�Y�V`2ؐeѮdJ�ڰ�����wa��x\�,���j{#9���P�ЕO*���ݕ952�Qخ&9I�q.�Ɠ(J�-]t�EU��ՎnyA.p�s".u�nv��u��C��뽛M)���z	;ni�6S�ߗ��)���?o?}��ߋ唇�Y���%Q��I���~Y��t�y�2��ilYguqO�g�������,���n�z�$�w����&��&{�ٟ�_���^Mm���	e�DQ�-���C�/_ٛ�	��YZ�%1�`�c%ه	��]1�)��srY����i��6-�M�c)r�XW��wc�h�.�2������m��5\��^043����0����4�6t�h��#Im*O�����:K([P8/ٕ֑l�p8��4\��]�)(�Im�J�a�ܳ(��emh)�]p��.d֏.��4�0�l�R��?�Ϸ�}�����m��fg�o�Cm�m��e�}�}}�m�}�7ve>x��m�:�Z��1lc�F1��Ō�� �,��eI:���n�Z��`Z��iq6�ƭ�ەqM.������mE%�m9���!#v�(���]k��q����	M�j����n!��l���j���[i��X����o5�HƖ�e�$ٷt,���n�of�d;�UZ��h�lU�fB]�T��9.�K�8ë6�Q����C1f�i�&��r͜�J�v��Mh�M3cd�T��\VS���1ҡE��uҋ��e����m)��-��YG*6�_<�Bi��kr�&*Kh��&n�6����aJ]mҺ(m��ˬ1H�[Y��$�\c!�`5h�d�5L�B�2�>��#>4��I�Jɟ��̛�C�R������ǩJSCkm��x���~׭��ӏ�J��q��"c=OM�Q�ؚ8h���������!��ѴѨYDJ"%�����t/�
>�J#D3B��ϊ8��#�;;,$���'�L�<mwowM�W& �k)"RAx��U<��س��fQG�$AL���=�0�̇1[�b&z�~A���0���1�_��1lc�V���V��jR��Fe���H����!t���ފ#��L7:�Q�{��$����	���|P�a�/@�B�SqS��CDi���0���3�٣����O�_��<3K0K�?+}6zp�@IY!�Rp�z>��R��%;r�s3�p&��mj2M�L嬛 �դ�:p�JaD)�4p�aO>�iz䙙��Pk3��L!a�֌($@��?D#�MUTiH��E�4�눵8���mn��u�c�1�c�Z�ǫz�)O^��Unn�k^;��u�EIt�4v��s�3=�F��6c8"O��ӆ��@���3�w�H���^c�x���|$�Q$�h�O���>�� �	��[��7�/6�[.6��n��U����g�9�����0���
�=F���r�LJ!���xl����bl؂&�3�`�k���B$���̜f�'�!FA��!�ÝN~]�:�_�'DA���O9�Ӽ���kb�~c�κű�[�1խlcսxڔ��T֏2�$���U%a8(��}4l�3������"6�?~u<z�:�柵�cǈY?���"XSِ��v��q��b�+��W4sTO��~�O���~�41�� �0ٓ7��"��������S꒟:�k�C4���m�����f]���=�%=0�	�<�.�1�|}��(�l�Za�.1?�D<�l���%?}�����[����
!���SF�/L4�7�$�Z��]z��b�qn�ű�[�1խlcսxڔ��J/��t)��VR����Uj���fƫRk��+��1����LM5�	I�Nv���v:�uwv�Bv�b!4���1�Bt�ݖi0L�C�tINC��{����mǨWRV���y�e�ֺ��K�Fj9%5e��B�U�3u�f&��$-�5��[���1���b�d�fWW�k.�f���&����k�qJY7�6W�)��8�aq�4C�K=���D2�"Dx�W4��{k�B��՗0�Ǉ�6�͞�C$�ٹO&ϧ��Yٯ��b��mK�vzl�	􁲈i����X��4p���\s%���jQ�ɣ��:3�?k�N����M�RSӇ��BD��O�-0f�"���I�IQ�&D��HTMWFA��(�Emi�bh]�υ����;�b�H�A`�n<��m�Oæ�oέ�:��-lc�V��>6zlх)M�Ur�;�P��HD)jz�Qx��^!�V��>R�m-u�\���+t_���&��+Rj<l�~Z�!�MM|��{	(?Igh���ק�������H"�-\�Ug��<�ExBQ�iO�v���<����V��C`��%*R�[`6��X���vh������QE;�~$e�yne��߭[~2l?M�ޯ��h�ၡ�%(�͙Ѵ��N����ׯ�S���c�u�-�Z��1��kc���ԥ=z�d�Ԇ�E�AsO&��R$"ͳ�.6~����k�=:�a��&��/D%"�5��(�U�l�n;�!x�~m㌓T���U�ʄ!'��g������WU5n���.�Ի��N���~�y��f�L�aL<=¿|w�D�U��k�$Y�?i����*�m�L�}>^.�O��?
 �������W�U��X�6�y����X�^0�}a�јP�4�㏖ŭlc�V���V��jR��)�-3
�M
("~���913�]�}��&~ 0~D8t�$�͘O����8Q|��}i]i�ɉ+y6�����u�{����Jj��j�-�#q�9�y ���Դ�����S���x����{�Ç���(����s�4��6����0B����NO��w��J��I'��N*~6Q�&�їVߕ��B�0$A}��$G�\g����2�4��q�:��խ�[�-lc�,�H ��6��權H��"&b�f����v��;��ݏf�gz�4ݝ�݌^�)4 �vݬ{
cÕ�g�n�=yl��t�kV$u�Ӳ=\`�/�)�4̱�@G���6���jc7�/WK���Կ~�Bw�-�<	]떚[�m�y�ă�B9.2c!P&%�*mf�L]�+�K��rZ�:К[NT�A&M
7�=� ��QBfU�$�����˙���8a�C�ç��f�d0����Q�.�9<�h�����L?z���Ŧ���m_6pN��l6nL�W�ó-�v����6޶R#�R�M�ZޱҿYH��fg<v\����%B�]yyK.�m�?}y���(t�hNe�JY��{��ʐ�t�cn���=~qź��:���cŭ�z��R���ԯ�ySq�JH�(F#1C�'9�X=�",��L�p�D;Sw�3.\�J�=xǇ������|ֵMS2M��Τ�.�U�u�kf�_�1��_?,08M��h�z6��S��M@����xj~��;���
���N,o���5/�`� ۂ16R�V3���"�=���t��^�~�|��GjMkS�5I(��H�2�eE�W��,I�2�xx�4�2*��U}�ڵ�^�`�4Ê8i��H��1�|����6��kq�ֶ��1�1�x��mk[խkuo��,�1�ff�i��i�C�jZԵ���o�����kZ�X�1�1���њp��8�I��3�ac2�H�X�qn�kq��"�,��ֵ�1�c,c�1�c�1�q#(�1�1�c�1�P�a�<x���T�,�֎-�)kE���[�Z�Ǭ=t�#�Q�p��X��ecZ޺�]u׎���c��c0C��Y�4c8c4�D3�$��(C�@�C8�i�5<��2�7�����F�s���y:\�w��_Zb�{�^�"ȋ�5[S�[�TJJ.�s�5;�r.B0��c�p��F�+�'�:�i��ݭ�Ȳ ��t�A ���!(��8���i
���_.��V^��MB�j�L�3���망ۘ�Uױ��Sr���"�N�u�5�5ޑ�0�R���3��
j��<�ɇ�7}��4���9��}x��g�bb��ά�:��PՔ�+bLɌ��Pu�W�V�PGD,��.�X�*�z!B^?I�;�6�7��q�ff}���m��7��5�ff}���m��7��5�fQFa������Z����-�c�1�޼mJSf��sB�DD8R�����5+s����rS�D�|)�M?�!�#A0�u��������+S�Ӧ�
'�w��G�̛^�4������e�Ɣ�����Cm�� �G����dv{ya,|��M	5��#�yR�-ÈȽW��v�����D�88�W�e1�8!�=;&���>�'�"�yVf����R�G��D���ROc����O[׬z��:��q�:��ŭ�[�1lcսxڔ��^��|�m�����|�(�D��Gޢ�B��d��@�ឡ~$to��0�!�t���
j�j�������P�ls�Η:XZ�%�>q:��:hm�kґ��#�c���0L3������<��	������zvt����C�a�
W��R�`=6N��0���h��(��a��7lk�_���l��S%��|�:�6��o��^��b���1�1�b�ǫz�)O^��U$�O��n
�u"ܮ��f�ٖ
�ۼs�>35v�SN�M�\��@+&f���`��mf���j.��!��cC�t*��XA�]f�M����!ԝ:6�5����]yL:�6�ݬqUj��M0�iF�kf��&�s����,J����a�v��>z{��`	�GD���<�>ߚ.fV��ʩ�ʓ�ȍ�߭�ﬔ�>oP�	ϔws3.Q��>�y6l�'�|�M�	d��M���l��WO�38N&	MS�M��h>�qq[��yU�lŭ��"$�����f�F߿�#|�#�Բ��޳�R�g!K���֙)�Sl�]I�������?�N3�nK�@F"~S�+��w\�M˙j8T��E�_Ya�,�M4�1�|Z��X�1�c���ԥ=z�u�a�db�E����F�����n��e�~^�;�m�Pٔ6"~��;�4s�K���J�@"=�P� �4�GXX�
Q��r��3��������S�pQ�&�����������B1��mw/�J���\q�l��u�$%������]���D>)�x�bjcƴu�s��kx�7����?J����l�زaW&��M��/O�<<<8|z|[�:��[�Z��X�1�c�E)Jl���KSY%��n���)���iX"&�Xh��N��Qί8DL
a�=>��$Ќ8*�$A򎙙�ҁ��E�!0�J=5h�t��@�l����30un]�H1@ҍ��.�_�?��o_����=zڜ�l�#�(�'�ơ(��o����3�EG���~�K�h(`�w?-����pP��`T"8�f�S������Ɣ���ڋ���Y>���"�=d�a��\q�������c�-��E)Jl��ȫ=���*�{�Q`�"i.b����!D8IEUa�#�Ld�yf��й.��g�>���iƠ��k���N�[��5�h�k�N	��O��l�6$A�b0X���0Euʹ������k�G5�׾�>Db���Q�#���~��i��4��C�Q�De�Y^�E��g�\�8"R��������`��KO��[�-s����Ђ'g�IFy���(��h�8�M?������c�-�׊R����:��4�з~��ws�+�|�Sk�(x�hC���t�	���7�o9�f�7�Q����WL+ʳ���L�U
k �(|�75V��W�A�A��Ku�R�X�M�8#^S��[I5~�������}�@�����&�lh�JW��e�1y"�f��q)�Qu[-���wN㳪8�m%Z�FR��G������B$�g���2" [�����a�N�pN�G��>���Ȃ'���U-�0��"j��4~��m�6�4[K��0���Z�6�#*J{�b�N�>{qN��0O����&�xR��6�h�B�w���H��4= �<�lXh�cJe�@��j�@�#>��6O�<	a��r3���3.��)�o�-žu���b��:�1�[��^)JSׯ�Φ��D�4�'%76YM�KC�Hg�z�����G{� �{�3��&�B�ya@�I��>����N�C��ٳ٣���}�8�rҴ�Ɗ�9��}4;�4l���%
&���W����%GDm��G%�F�l�������I��#>�'y,(ԣ�rKd F(Jϣ�ER��(���X�IĈ E�����FU	L>:P�?kG�/�1�̆�kG���mǎ�?1�8ŭ�[��1�b�=x�)O^����� �D�ƙD���'�6~�O�)�߽�˚�G�<*>4rh,��kK9S���s�;8]0ϐ�ܝ�k�!/�o,���l�nuR[��4&�Gik�:����vi�=��!�|��~�_�������t���ڋ�u�jS�oCGaL�݇¨\ƚ��^��8a����$
!�����ȉ0�I~�J\�"<[:����b���-�u�c�1o��R���_^����M�SY�]Q��7ڊ,��fCG���iD�90���L�~)g�����l4d�ꕁ���]2�H�hLL�z:��
AGu�����
�<LCa�(�2ϡ,�Gsa� �����	��k^Qٳg}ږ�`�x��ѣ���d�=3k�"w�����|㙮>2?��rp�����<0�F l�SG�C�M
Yb0DҲ�(��`�?b��"��?���M���#	�����Jxyyo;u��x�t�Vꖷ�X�Q��1�ь��1�1�����:�)���|�-n�Q��3M0��i���c��H1�c#��`�1�c0c#�`��bƒ1�c��H�8��Hޭn-�Z�z�Ȳͬ���f��c(c�2F3FfY$��`�1�c�H�Ye�P��2�$��h� ��jZ�)E�Z����|�c�6���c���ǋ,�e�kz��o�]u�_:��c1�c�c ef3�i��!�a$P�!���e�'�9<G�?T�4s��f��sx��)���̵vZ�̼��]�T��ʁ�w6gsc1��!�ٳ;���.95�y��^��7-���<Տ�M���2��KV@�UUP��V\ժ�
n��>㽦�8c?;��;�v�l��կ��Z����_.�{�fxo6������|���c��l�N�Mڹ�޽�f^����oi�(l՝�޸;ӻ���Y�������嘽�s6��q�.�<�����A������K�8���stN���[d^eT�R�n.%Z�Q��cr����E/f\I��=���X��Lr�d�+��~;ޑ��1s�RP���~G"���.���+˫��b��#ֵNd�����^c�﹤��8Kn��:����r�T��KbvmIV��:�6H�.J����^�f�7e�I�˚��f�5d13.m�f&���L�;y��S�r��Б�f8���{�����gG�Z�����}��7�:m��t`��"�f)������؍�F��4i��&��)�~f�� �G�,�qI�����M�cD��њ�sK��f�V���@.��lf�3iu墷ܶ���7;t�\�p��cv�biu�bWKK
7J���җU)��ļmy�6%f�-Q��8�����&��-�1��6W�o)��)v]��l��׃��b�\m ]m���T��	u��lk�bik�Ua��d���]sJ�:�Fje��bb��ޖ?�y���m�}���.����M��z���컿����m����>˺��>>>>�9���u�cc�1�[�,�������dc�(�#v�M�Lp�q5Џ0<3@]a��n;nX�X],l�n��v���K�lJ`Q[nV\��b����M��j�YS�iTrXi���FX�]Gj�fk�t�ضద�qhX��bSk��5��Ζm8�Y�	f��[�
��n,����#J���/�.�.V9.H&.b�^*�[̖Ŕ�[��Cl�έ�f)J��k��p�B��һr��չ.l[
��k��Y���mY��\j8�vi��Q�Yt�RBw�N��l-�+�偫P�#an�j�	s�`�[.�]�-VWGFm��Ybr��q2<�mڑ͎��Y���������W���PI���A�����ہOI�����{���2P�� �aa��}/��?��*�w��lg��OU�!pO�����t����8�x	�O�G��Vl����^H��O2�G��"���Ƙ~���
f�I$�B��EL@D�ʡc�j6�.�CM.fr/��m��9��4s�R��?l8~�U���3�nbXd]�Vb��T^�(�)���_??>u���u�cc�1�[��=m�Z$Ԅ�;q$�fk5��M(�*B|�1�RE�s��,�bPX���Sg�ѹ����Nx4>6h�S�$�)}!�M�h��Fխ���0�(A3�0�H/F���%)Q.&#G�ؓG�gv�᳇�M�p���p�����զ�EK�d�X����,k8.՛�4�Rw�ko<x�x��Qx��|��ӵZŰ�z�A�B����l���	`jO#{�naN�\�����͞�׼LE:�����θ�ַαlc�c�1�|�┧��}�:��;��A���c�h�p�?L����8D�O��Mp��K����aҋ����W-ih�g~��6T�����N���2F~�g��O��wa��X�Y���Ml�A��b
S�f&��1��!�}^D���=N�CE1\'�"��Q*�׺�xs��T?��0��[usپ���MO�JQ���΍9F��ދ{���_�T�uT��k�l޹�m�1�>|����:�Z�:ű���c�-�׊R��l�"�Cl���U��@�E������}8�:�5�o��Җ��%���'JJsi���x&���&�jo3*C-�uAt�2�3��.�Ӆ7���y�m��K{U�TH��m���T��⏑��M�H�S��|���~J���J~�τtPOa�����ɳÓ��[�u���=<�O;�G�'۟�����UQ?O�><0C���)�F)�k�x������Z���V�:�1�c�[��=Y��_>�ш0��7)pv���b���e��Z8������x���6jp�f�ڗ�R�����u�#aTd4$.�פ{[�L���c�������N�6E%8���krY�Wm]GU%��Acf+��h��a,�؛��ѡ�t��+��3leN\Ԫ���S�0�F!�9���V�4~8R&��&�!�O{������5Ra���8e�����3������G�J������q�4�ƚ�>��bN�w��?z|�����x}���O�fa��-����ikU���pŵ�6�e�uUM��/A�Y���Bi��~���`p�" ��H��i�,�O�q�8�\b�-�V��1lc�-�׊QM�n](WxXT#
9�Q`���P���dD8y9��5nNk[=�JM�هO���b��i]��!���2~C}:aiD�fM�a���ѭ~{���A6K!����2-+0�P�����?~̒>��iB�^:eo-S^W!)1�3�.f�гJs���9(��Ǔ��F�ߟ<��w����k��Ȥ|�o�������ș �*#J�|��|a#>5�n���x�]Z�cű������6a��$ޕPNN|?����N["�TҨ԰��{��TQ3�KI@#=� �ǿY�~��j��e�xZ9�6ۇR(������U�ĤJ�Vؤ~t6��A��֦Ֆ���M;������>�Qz���Z�u#���X��˥�1�R:��'̐���y8!��N�BS�8�S,\)���1��5������~��_�)�5F<g���4��>8��M4�e�[�c�1����)O[z��Q$J)`Ҫ!������^gK���m�vn�����g4H��I����$'~�3�m�̉Ze�ҭ���BT�#�cTq��꘩���|IL��( �=�d�������$芿���`���Q��m
v!D������tn~�?jx3�<g�ڡ���J���0��>�~�>(������`�"f0��Bi�v������8�O[z���c�8��n����1�c�սI$Y%�5(�.�1�sVG���w�n���}��{�|���3��[�Q�gg����ij;�v>���!���X���e�i��yi�q\T̫0`�s��ӷ���E�5�����#���6�ۍ��u��x󽦝��Բ�A�ɫ#6ճi�� Hsl�tyG�[P��J[��"��M���]�5X��43-��D��6��ya��l엔ͳ��r{<��M�4~��������e���C�aDa'� ,����O-��xh?2�&I�+���2|Q�5�^����kԈ� ��8h�����њI�x(��;'?'���}��P���I̐�sغyNf��P�����؉�r�5�� �v�����k���̓s��V��	��T��,��`�����Y��N4�\b�-�V��1lc=[��Q�X��ITQ愦�� SڒH#���Z~6q���?>��m��㚥��ДO '�a�N�x]��N���f��&��PI>������a��拇������<><:}������Jxm�4Q����L?���ݵܡ�gKc�&ĤsR��ħź��/�4��h�S�⃅����oM��h��5�� �$8L�y�.dÆ�k�7����x�a�[����ֶ��֥�kqkRֵ���žZ�"�,�ֵ�[�X��b1�Z�q���q�-k-k31�1�c�Y�C�1�f�dc��q�:�Zֵ�n-jZ֥��e�1�h����`�2�@�2�`�1�1�d�c�a��I$31���c�1�e��^�YkZ���-kR-�)k1�2� �#(��1�gc���b��x�ͭh��o����뮺��X��S��c�@�2�2�q�C�8���	 `��22F1�tִ�Fҹ��,x�S�^%���� "?2ǹ����c�+��������e8&(V�Y+U�Wk{���6�Y��x���F
��|gf�v��޷��!à!�>y����>�)-�l�}�1UD+~n�&������!�9����癊����^-u��ԩm����a�:DTn�OWB#&}J�)�F�}��|��??�i�|�o_w|}�w��}�m���w��w}��1��m�w}��E��1�[�8��n����1�c��޶ڔ���k��$&�c�Y�.|�֒BBȄ����B�s�ߟe�䓎#\3��ʒ�^>{��!#�=��Gǽ�a}�a��axa�������d+���XG(KH�����릖7Pu�k-@���S~wE+���YoJ9�3n2'�����ȟC^��t���ol�T�5�M�GN�$��xw&㦍��?)O��fa�z$��T�Da�,�f��4�6��[�c�1����m�O[6l;֢��J���b;�T�O��sύ:ֳB�C�	��E23��M�O߸�r���ɣ���9���պ3sF
�D-���>�D;�^8�_���� ������SaӅ��_�>:rI�� (C�Ú����p0��ft�S�)sN�ʨ��8�� G�#�A�����kR��y���D�'D��Q6�Bٳ�Y�"+��M�#��j<|/O�*�f��A�i�៍0�_���ukqkc�1�սm�*v3���d�v����K�)͕��1��LkS����e��gac�D��J5����0F[݆�͊�i���[1�CM]*7b��lԮ�	ye��
�Z�^-�З\]��| (�<j�l��,v�ۀ��6�iX!���Z]����Mw֔ 9UkL�mDɮE-uZ�FM�Y�<�y?�������١�
��'�%��H4�~�S$I�Cnz> �
X��tw�!0F�P��«�ep$�h�:��aJ�$k�f'��g��?4M��a��S
��e��C����|P~��~��6��\����� D��ؔJLhs(ثG��[ZD�L;Y�g�J�L)B�~)�俿�^����O�i��Ƙi�#8����ű�z�o[mJz��e��L�sXWxU�CLk��|UA'��{'u!9�j�p�x|k��
'&	��4\4'���00�6nt�j~Vrj�6	ϴۆ���t�c�'V��<�
w��u�o�
d��ն�z񦶥����)�m�~��g�x~��Zb�Q!c���K++7�ι �b��������J��a�I=Ơ����<��j/�na����P����)f�D�_��XV�g�>	鋹�6l���b���b�[��n-lb���f�M�aJl�f���6��i����Ξ�zj��8~��f���醍JOX���l�p٣�e<m����)�4!��^�S�e�~��X������A|q�H[+Y����8a�feqsW�ݞ��'�M
|Y�u�5�f��p%8I�E�#ŕd�����X��Jh٪�l��z��Z�s�6�ּ?�����4^
������Y�y�#�e���s^���'�V��qn>q�嶷]Z�Z���1���0ن�q��T��T�^ѷA�U1Q����F~�|�'��_C���ѷ������X�sr�DIG��](���Y���0�T9�O�J��{J0~�=>�K�T�^�[Q�=|���d��I�_���s2�7���S؝��t�����ɣ"���~�8�E�р����`�������Ҏ+Nm��[ֶ�G[q��o�>q�-�����ֶ-�cǫz��3e�7��>M@XBɀ`�˪R���{[{n�H����"mI��v=���L(�ʺk�r�ݵ��L�u�ضVD��f��qs�:��sL�-9vv��h�L�7ջ��s� $#�6�t�U�e-R"FR�嫝���ĵٔS&�b��n	�]����f�yq4��"��5��[oܛ�Nϸ��ș��-8tg�7����j󍹳Ȝ�=�:y98<��K��Oti�5�	F6�ۆ�[}�Α��/~ּ��E�x��(7��Y�	3ɢȂ&��ʲ�uv�`���V��w�I�=��{K�˭h]5��lg��t��#nIm�X�Kv�[���0�NA��i���HTQ^^��>(�>4�M>[kuխŭn��coV��ԧ��SA�^��}֒H�DadG�|Oc)��g�PY�jӃ����Y�J"����^I�{�Su�����!a��T2!�XHO��4)y7ξ>l����m�T�[J��� h����o/��C�c
),�i�f�M�ܱ�����g�{?јo�����d�誔��AM�(a�~)驓�c>98!ã�m(�O�Y��4�M>#8�ьg�����Y$�Ad��;d��p�r6}�`���T̘y�%��å5��t���0�����Y�%�I���6�.~��������_=8ϧ�X����Տ3erJ�60��#��Z����~z�a���o
��)��
3a�G
[Y�=
8S�G�EgC���=~�pĿ�~�{=��S��ѹ��_����̹��?Z�iڒ	'����~�(����8�8��-�V�����1OV���Sf=�d�!*;�(�q	���:�|�6�����D2j||nrwzs�<��pO|��7'%&�mf8�uؘ%�蚂p"m�ܻ������S+��6[z��U��sZ�yDD���-�z^��!���Wb~(~nHc :]0=����s�A��N8�p�q?{E�
g�9M�eq�{5��������%y{��$�3J8��I���e�k|����բֵ�k-kYf1�1�H��1���fc4��kZ�c�:돟>c��-d1�c��1�c��"FP�1���1��3M�q�31�2�1��@�2�����Fh��`�p� cC0c��2F1�c0c�$�F1�e���c0��cE��$c�I1���QDc0��H��1�aF�ķ[x����k[�^0�lcŭ�ֶ��u�]qո�1Lm�bַ\Ykmkx��[�,�1�a'84�H0e�����2�8��{�A��1�����.��������e��<���o,�-v%s�-r;�n<�eH]�2}[�z��)�]��3�Ya��*7&��?}�f��p�ǹ��
7�{�R�*�D!&�Wӎ�E�E�O+��|�n+fb�>�YDE�O�x�[[rZ^�(�2��"*qVfeSQo&�6x���y�籣|��7�{�why���]���VM�]U+ۊ�uf�ad\����,)�r��Be�]��{F�l2�g�_��/^�����y4�n���vU!�;��̬�y��^�~����-�3R���۽减�yI����B�[��h�I_�2����Os�f��Zl�<��y{�1fŕǖ��)�h-��뻪ҹ�j�w�s:�e��m�B���v���w���>�in��I�e�z�a�M�c�Nf�|f�6ݽo/fٲ�)CZ�����<gn������-�7��de�k;Yy�:���3��XmVV�n5�f�s���&�K�Y��d�9X�e��g�f�0��⸣���]XLi�,���]af�ٌ�,5��Jp؅�ظ e&EBk���+qy�m+�mK��g��!��9�׌v���¦���cK֬`9D&�0�J�U(_�I�Yqμ��]�e5��h.4@Smt"hѻ�Kf`��3��u��դ6�f���$��$�&$���W�����6�}����������m�����������m�����tYg����i�|2q�-ŭn��b���m�O[z�fw��*,�-ի�Ff0��S,U旭�tn����*<0v���ݻ�-�U���]��kp�5�5n�6H�mrƖ�n)M[���(Q�1���F�1
1&��Ɔ@F���e�㔥��ʋ�p�eܴAp��G��y�i��҄kne]�kyP �U�b�bh���\��YHL�⋂���d�XTM��Ͷ��ռ1�Kf��niB�k����i�͸�N쳢��g.�Jk<�[�  �q��Y�.�F�,Ѥ4eu��n�KҮ�n�&��9!S`��I�
��B4�k��)HSm�L���&�bS��gz�����0~�RV|n���Ʀ�Y�ð�8�s�v>������mX�f�'��D4w��3��[�'�uҕ��}��o_�G�4#=,�a�4_#���ɁN~����c�6q,&%�(4�
 �MiJI��D̾�#�w�q�1��0�?��qkqk[�~c�o[mJz���� ,�/J��P��UPNY��JI�� ��Q�)�G�z�y�	�bȰ���i�z��\��ߣOfá�	��w�߬����[s?^ynf�K(|D�zy��R������JǙ���f0�
3,a���KT�w����w�k�'���z5t��6&���Nd��?p��I58xQ��0󠹯��6r(&	>4f��3L0ь��p�jַV�1OQ)�o���jI��S�UA0�
*ÆS�+}֋o�zop��`'���О�}���H��b"!o� �����q�8�����7,�����6Э*�9�����hV��O����m\��@�O6���������5Å?�<�gG_�ٕ�)��0���q���,��H��*����M|�[�+^>S��q���-�V����1�z��Mh�Ou�\��8��'�sb��~<����H�P~+�_��!PL����ݱ�x�8�Nd�6�؀͢],��E�V�Q O�Ic>�!�؉�^/M�{��o���|T}�p��g���&M���rg��t����0�PDw����>
(B1Țǚ1���S<N���g��#rh�?w�r��_��:�6`~�Ͼ�O��~(����Ƙa�� g2�Z����)�#�<m�TT�Ues�11X۬�#U���L^,9s-)H�+@���1�1�g�eV��:]�8$��8�p�l��%�Ne!���AC[f�Xp��1�j񘚔�Uٛ`M��_B=����26[�n����қ���ļJ�ɪv�#e	��R;V��tm4�ܲ�d[��\E��A����}	��9b�K6�\R������'��3]ְ���N[׿��G��T�R�~�N�Z�����l�CE
x�~���/F�0uҎ[�f	��t�;���Q�D�����ls+R�4dM��>48'�����dN}��.�V2e�X���"�-�L�����c�P�B�e��Ї�~��<��NZV�np�����1�>q�R�ukqk[�c؉��0�+��mU����+�@X�q�(B���%�2E�$6(��C44����Q��Y�#�?�pW�pRIO�БǱ�R�[�jhr��a��\��G"庺Q	K���3p	;'��4"��%�V��|����<r~�h��a[�	�Y����I�:�(c�{�%�-0�	,g�qƘa�-KuվZַV�1�dx������(����D�F�UTg����᩿R�|�v��=��e68��8m��e��~-젞ϏG&��,3��A�����O���������v^X�C)6�-��w�V���4zd��`a��U��d��DJ_?@�|O�|*0f��PK���n53�}�s�Og|]�.�g� p��4h�٬���d�%^����D�P���?g��Z��|��n��c���My8��y-��I|�Hb�AB��UA=�c�>�.k+�����g��?;�_�6��f߶��<,ke���P���b��Ɲi�i�ي�r�0��C�Սأ�{�5٫���������zG>:h���[�|��N�0i����Cgz�̌�/���r�0�����(z��[���^m�#����$�Uy��T�s]֣���OZb+|�zk禒~4៎4���q�0c����d�(��Z#	���5]Q>&iJ�s�aԊ�Kb�m,��l嗻�Խ�ٕ�f�󺆰�w6�15�ٕ�u��nL� X��P�m�:8�B�՛4SQ�YYLin��r��7r��l{�!΍K&�(1E��b�b�֦Z�tn4s�6�mxE��,.�)�T���&�g�?1S���<�	���f��/��,�¼��%$�E��'EA �(��>٪��T�F�3N���qХ<fL� �$��[��O�-������ٻu����o��Q�᠄x�f�MN�׭6��-�|�մ�>��K��R�1,%�5L�f*���3%�=݋̟g������Қ�X��g�wg�8-����V�}>��?i�3�0��!�p�-k[�c��<S���Ȩ��ٸ�)�I$#�Fl�z�^���[��n0�F�qi�K�ѧN{�<�M�y:|���--7ӡM�Z�N�������C�xoF�?*e��cG�KH����,�C����ID�'�@�O3Q�8cVb���2�J@ڦ�빫��5��m�="�l�H��DF��E!�0���ØZ�����Q�b������]�n��{{mxh6��>ץ=|��^���[խ��բ���Zֵ���kE�n-jYgd����cƖ!�c@Ʒq��q���1Lbֵ�ьc�3F21�3F2
�1�e�FQ�q�f�1�2�1�2��@�"�33�S�V|�,��E�բ�-k2�1�ec��2I$��cC#��ic,��ad�duH��Z-m��Ե��mo�@3F3
(�`�4��P�5�k[۬0�1�cŭn��1�]qվc���Z���H�X�`�4gc0���pi��0a������2�*���5VB21<�Uz��B���+n�w�%�J:n�*4Z��\����'����؇�C�]	�Mt����Ut��^�)S��b��w�ί�7�#���"��QY
�Mss�2�k_:����EР��4;͙��[�H|Z�[	�J!1x�lD�K�P�v�����j����z>>_}���x�O��m�w�\]��}��|�m��w}������}�ɶ�m�w�]���>0����\q�Z-�V�kZ�Z�Ǫ	�Fg�u�T��j"	�D�����h�h��z��r��R'x��~�o�x߰�W���
���_���a3�NƖY��D��B{���>4;� ;~IA��#����A;4a�K�L.��g����Q3�W��pa� ��*��-f��&*��;D��DD��!agƜqƚa���8fc�[�Dx񵹖��$��3��{����U�815�O�N���N�%pD���i�<��S:�#�%�f�:�ݥү�����N\�~�s���OOj�'�2�ϡ�T7<��}?I �M��.��u?*S���2(��¶h��y��y�-40�]B�����l�̐����!z��Ĺ�E�3��zg�K�h���,���i��M0�1�8�1�c��Ő��'���a5Ji����Y�q�q�����L�M٭E�{[�׮�c��fӚ�N4�)5v<�gN�jy��t���86��b�I2�y0��9Μ��Ӻn�ΗSI�q����SSSV\����i�irݥ-!�t����DdԚݬ(��a��� Ŷ���f�����P�[���R6�&�15V�jX;�2���Fb��ź1�U��4�~�4�=g�J�"!I2�h��i��g�}~��ws��6>���3��G����?�S�y4�Bo��Z�9�������TUUte�7�ޤ6���S�����d�Ӑ��K	����?�]��������ה�%RhjM1������h���'��9���?/O�.�����sxmیz�]u�1k-�V�f1�c>>,�E�I}����I5&R�DzUA�,��a���O�I�qtB">�~}��95�~��2�'���#JW����8��Y~b���~�Jt5ϣ�f��M0@��~����Ȃ�%+c\�2P������E���*`�~0��䨢�/���pG ��e>�%�<���J0����#�ex敘 �B0�=���%AU)O�eQ	g�1c$ c�8�\|Ŭ�][�kZ��=Q�����,�¼�� ����i�sȭ�5S�'|q�%��o�IIG��1�\%;[f����� �,T��v��2ff)IȉZ��\ך��[����<�i[D����beX�5$q6��Di�)�����"0p}�����{���Ie{����&k��J��bUFG�9��pY���2����h�LU(�I�	w�E�\XQfi�����|��kZ�Ǫ#׍�{�4�iDMZ+�*���9B���?~���`g���p�� $!%��1q��p�>��;�r�d�q�lBQغx�)���?
��5>֛~���������4���IӈЧƌ7��g\��`�n'�5����r~>��g{L8�	�O��
W%��2��V{�(����S���Q�x�m�<����?���ED�2;` �_���"h�XIgƌ�gi��3����||a �(�� �Ol�M!.�U4y}�����,�=�8(++0��i3b�v	;2l�i*��w���3`���nJ�Z��WV5.Y���V���<�mt��Y�ͳTn�&@��k�ݣ5���v�L�W/����k�_�[���n����S�ƪ�e���c���[s��B�%D����W]+5�yk5W�]��tƅ��iyZ�x���|���+��W�3-.(/>J�.j,��L�S�[���R�0����P��{J�=Č՟��ֵg��}��)����.f~����%9��H��O�'g�tٟ"��V��A���a%{|ȿ x�s*`^��XBX��;Z�J8�n�GM��%���=%�	�4��xy[�hM�|�h��_�N3�+Ӧ"������q��M0�0g33�OOOO��
	�F��l�+��"�Y�!s5��>?���t�!�$A􊏴��E�)-8���FB��~מ4\؞�k�iMby�?���?�|T�'�Ɉ�i�`�Z�hч��ꋎ���e5�����[+
�R�˭��ry�Q({�SML��ek�80��Cn�M��v��_N�r��ug��m���*�n��󅺶>[����-e���-n�k[(&�t�i#�Xc1%A��֦j#j�Edw�~<�g���q4�s\ms_�=׈���QJa�6~iZe�ΰ�Ǧ)>8k��B�p�д:�@����N���z��)���Ȝ�I�n�p6+(�kH�@Z�]�f�����vY���<1w͓����V�-0�@Y�2�=p�<X3:t���E0��MIP�+�׏_<��iJz�5����ǎ����>~Z�uվZ�Zַ�>T��љ��Z@���^e��P��O�>�S�ӆ���1?'��r�}����1�ǆ4cZ勘�!e�%���G&ϼ����
	O�D�+U�{�ɣg���a��M9=2^6D�s����ޟOީ�zz�)H��#5ɮYs�4��=�"5�2�U3]H�D��ȸ,����+�{��A��I8�$		�(�}o �J}��r~�XG�v{D�b�4э*�x�$�#���|k!bMtɚ$8$"$�H!D �HBkP�&�BkZ�!dAH�H��(0A#$b�&�BB	�@�$`�DD�1#"�0ADA�2D�1�`�"��"AA��"@`� �H�2 �" �$dA" �AdA" ��BD!Bh�j�� ���� �D �AA� �2 Ȃ2 � Ȃ2DZ�!5B�DֵMj�BZ�jD!BkSZ��&��B�!H �	# Ȃ"BiB��ֵA	�#P�&��&�B�֦��DA�	`�D ȂGZ���!4�!���!4�֡B!4��A� ���AA�	DH�D"0A �D��d�ADHBBi�&���!�#P��!BkP��Hȃ"	ADA"	#" �� �D&��"�֦��"HAAD�2 �$D�B�&��BZ�� Ȃ ��1I���B!Bji�B���F�5�D!���$A"� �DA� �22D� �"� � ��A�� �" �"	"2"��dD#Ȉ"0DA"20���"DA"" �aDF"� ����0aDD�$DF�� �0D� ��� �#D�H�ADA""�D���"#�"�"DdDD�DD� ���"DAA�0DFDADFDA�DH�""0D"0aD�(�D`�"�20�"DH�"��D��AFDA#AFDAXQ�""�DFDFH�A""Ȉ�$D�" �AD��AAH�� ��2#A"��D��`�"��AF�""0DdaDD�DADF�$F�F�a"�0" �A�D�"DD`�"��AFDA"DH�DD� �#AF"�2"#�1�0A��" ��"1�Db1" �DDa���D��1�DdA� �#"2"�#"$D�ȉ�"�dD�D�Ȉ#D�#AFD`�#" �#H#" #H�##�FDH�"$FDA#" ��� �AF � #"$F�$F�FA�AF��#H��20���F�#" �#�2$`���F#b2�0Db	F""#Db"$FDH�2"�#`"�0a""A�2$`�$FDH�����Da�0DDF�DA���"FH�1DF"Db#������#DDAF"#DD
�""#�FFB@1��eJR�H"E �$R(�H
E ! �����F��`��HE"��$RH�E"���R1H�-)T��i�&���ji�#F���5����)�i� �ִ����H&���i� �� ��
�j�`V`�@BA4MkH ��TkT4� �kPCZ�h�i��U���U��q�m�SH!j�&��Z�MA��"	�4�4�D �$��D�"�HĀ��"�`R T�`��D�H�L@�&A 0B"�$FI, ��H�# �2$A�K$HČH�D1"	# �F$D���$bDB"b0H�F!#�bF	�"$bB $D�H���$H�H���A"D1"F	"F$H�"R0H�"	0H�H�$̸�#��&F$A"	$A"$dH�2!$dH�H�"	$`�H�"$A#"D"F	HȄ"	"D0H�F	"D �"F	"D�H�Hȑ �$A"	 ��D"FD �FD����H�$FX	 Ń10�#�$A0H�DHĉ0H�H�"A�DH�# �0H��4��D�$H�"FD���# �D1�H�H�"	�"D ��"D�2$A#"D�A��H�F	$A#"D�!D� ��D ��"	$dB$`�"	$A"	Hȑ�D��H�DHȑ"D�"	1"	H�$H���	AH��!Mj�j4M!F�ȂAdA"�#D!5�BHM!A	��#D�#HBP�BM�!	��B�BM!�!M!h�B5�&��BkP�B�&�D�P�BM5B5	��D#P�Bh� ȂDA�$H�DA�1 ���&��!	�!��!���A��DD#$H�"� �D � ��7d� �0A�DA��	DD �$AD#P�M!� �!4�֠A! �$A�� � �A�"�1A�AD� 22DA���"�� �A� ���D��AB0@A �@֬	�B1� � �MB �A��i4�! �M&�D&��MA�� �H1Ab�b���`��!�B �MkQ�jBF�5�֡֨�AdAA� �1�"		�B��"Z�BF2B�b���2"� �A`� �&��B!4�֠��!$A ��"	HA	�!!!�&��B5	�"�M �I�j�&��&��B5	�Ad��" �DA��kZ�BiB!4�! ��A� �� @� ���M"������d��a0thZS �3�����b����1�*1��� V�������>�_�P���-������(�p�0�8�����/!f?Q��;F�g�����[����|[���M���u�	�m[�E��9/�g����ޛR�^9���PQ�@��)�մ������/��lU  �&���DP>H,h�z���]���A�!�`֤J�e�~�p؛�gk����5aڢs����(8��z�����A�,� Xz��S~>��g�w( �fZd���II�LO��(�5Ն�!��N�>a�B�7yq��ѽ����$|�?�a�dn�).r)  "�EЩe)Dn (
���\ 
��C@��"�tAh�lEYA���H44/�@j�M�����\^�tB��<M�x�EĀ�����H�B Ą��"!	!P-(CZ� ��!�&����!ڽ|A���+��a�:��H�8����f#���`U'��������=���H� *"�I�4Ĳ�_�L�b�u{8~�cxlC�8���{Y ��9>s <��.O�K��H��Hi����j�s��i���@އTA����ְ#��x��s3qsp@9w�JQ�}*�(��0E�C�
Ey��>�)��YN��z<F��ޮ��܆�C1
Q�������{z5��"FBl�)�\,�X4d� *(@bX �6�[ġ����RP��iHR�� Z�C%/C�{ �hZ%Ł�\Q�lA2c%�2�9
�(	�<4�_��xD	�z��DP;��9z�[`x'z/Cu�:C�O�?}�@� �?hol�K�ԜKPNc����fc��ZDZ�HvP�������EZڢn��A�^�Ey^�NX�8~����rW�5M�����Sh��A���%�o��)����c�&�4(��҅�6���Q� ۹�!ϳE{���Hˁݝ�Y�0L6	pؼ���Ҙ �(�ޮ�����T�t�C�:��C`�b��ür��699&�r�(tđ���F��6CC��H����EP �����	`7�������8�@m5�T �(���.7e.]a�Šx�!~p�����$a�J
A��b.������ܑN$>Tn@