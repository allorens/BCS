BZh91AY&SY�	8�/߀`q���"� ����bG�                �蒑(E
E�Ԕ٪���D�(T��*�P�Q�)UJE"�P�IR*���)I
��UTP��R��AR�����U)Q(J��H��D��$R�Am��ct;�ZaR���*��T�R�)V��T�J�B�����P%o��$�2UT���\1�klնm�Ӏ n�����:�PU8��P��+���JQAE��F�J�!("�j���Kr={Ȁ�J�5���R�7M�ϴ��2{L1���7t⫳�$��h��{���gW]ݔ�˺Ի��tkA��ӫ����;���]��c[{Z:���P�	RR�J�=$�)@�g��AP:u�gw����.���g�5��Puf���{���m�����}>��ƪ��>˽潵R��ݗ�ʭ�������{h����zy�]WaUUϧ����v��HV�B����
%-�>��)@�������[�Wu�� �B�����.��
]��}��+�*)_g6��S֝��TW��ҥ	^y��=B�(�\�����^�o>�i_l(���<uA)P{�JJUR���*�ho�JR�@���U*���v�/�y(�UWއ{�}*��H���|�>*�U秝�*^z��Ъ��
ު�/QT*��^9��*��y�v�H�t��+�UT��U٥� 0��I,_X�ԩRP����eUJ	O�w�m�Uf�y�*�UT�z�=��hj�Q��o�����<���*��U/z�y��-=Y]}����)UO}�o'�UQB��g��U�b��ЩR�jSV�f�%H)�Ҕ�(/��}����q�U]ao���x=�� 7�hd��h�l���H�(�����e;�@Ң(
����-4����3�E)J o&�P���=�;�������� �>��6�h��k�����
ۓ8�l1M j
�I�.��$*�/J
)@�|{;���m̸ 4v��@P;�p GL: �{�
 1� =�輟p ��t.�٢ڵ@��RQ!U�>���R���� �O������ .0P:�|� �6���(��h�{�������� (���
����H)*�a�	J��W�R�o�=��Р�G��G�1�7t�4ò� w�7�� h�[���v�;mP    �     j`)T�      "��Ĕ�j�      �����@h4ɠ 4  ��IR��    &� JR�&A� ɦ�#A�O���M==CL��@h�C�~_��������������}.Ƿ��=��l�ٿod�2_>�����ﾎ¿�����*��������"
��t	�_��ߥT�� ��Z�I'��QU���EO�
/����~���L4�ɏ���a�vƱ�+
��;k�L�#°�+ư�kӢ�+�l+°�6�Ʊ�cXV5�aXV5�ecXV�l+Ʊ�k�����+
Ʊ�+
ƽ:k°���k
��{k�LJư+��+
1�+±�k
±�N�±�6ư�k³���V�cX���2��k+
��+
±��+��ۦ��:cXV5�V�`V�aX�ztV�Xm�aXVaXV4cX�5�cX�5�ecX�5�X�cX�5�X���5�X�m��c�±�k
ư�
�2��k
Ƕ5�aX�5��Xi�aX��cXV��a�V5�aX��k:ecX�cX�5�a^�5��V�`V�aX�i�aXV��
ư�k��Xtư�k±�(°�k°�k�L�+
Ʊ�aX�a^�5��V5�aX��daX�5�aYX�aXt�EcXm�XV5�aXV��aXV5�aXV�c�]5�ztm�aX�aXv��L++
��k+��±�+
ư�k
Ǧ�+�l+��k
Ʋ��+
��+Ʊ��k
Ʊ�+
Ʊ�4�°�
Ƕ5�cY�+°�ư�köV:aX�5�aX��cY�+��6±�k
°��cƱ�k²1���+
°+
Ʊ�
æ�k�l+±�+
Ʋ2��+°+
ư�
��X�0+°+���:bV5�bV;e`�lA�=�l������ �����5����X�X+X-`�`X�V ����(�"� �(�"��
�(�#� V���J�J�Z������Z��Z���J�����v�kkz`-``b�`-b�b-b`��V"�(� ���F��F��F�{`%`��X#X#X�X#X�X	X�X��X�X)X#X	�k++k 6Ŭ�逕�5���5�5�5�5�`�b-b`�`b�bb�bb'L��A�A�k+k k+k+0F����X#XX��
�� ���E��T�+ kkkk;`��`�b�`�bb�b�````�L��F�l@��A���T��H�
���J����J���J��� 逵�5������������������ V � ���J�Z�J�J��Z�
�t�k+kk{`b%b�b�b`v�
�0��R�P�Q��`��X�XX�X#XX�X#X��X�k+;b``�b`c�+ 0V�F�R�R����R0�������T��T�Q��X�
V �"�� �5���
� �5�5�����5�5�����kk
�lD��E�Q�lR�R�S�*V
V�*V*V � �!	X�X#XX+XX�X�X�X�X��)X�X��kkkkk
ư0F�V��+kص��bX�V"�m�5�`%bآi�b�X*V*t�+k
�]�F�F���V�;`�b��*� �(� �����X��X#X�X(V���`1��b-b�`�b�`�db�b�b�b-bX�X���V�aX��k����`tư+��
��V&��5�X���k���aX�:k��VcX�ư�k��k�EcXV5�l
Ʊ�k���z`V�aX����Ʊ�k
��(ư�k±�
ư�N���k�+�Mt�X�l
��tư+�+���cXV5�cXV5Ӡ�+
��{cXV5�cY�
��L
ư�
Ʊ�0+
Ʊ�k��k0�+
ư;e`V5�c��k��aX�`VV1�`V`V5�ea�`V5�`V��cX�cX�cXi��cX�l
Ʊ�zecX����cX�v���
Ʊ�
Ĭk+Ʊ�
��
��
ư�tۢ��zcX�5�aXV5�XV2��
�lk
Ʊ�k��J½:
°�v��+
ư+ư�t�cXVaXV5�cX���cXV5�X�bV5�a��X���
��k��k�MaX�aX�cXt±�k�+��
��X�Lk°+6ư�z`V5�glv�A��6��k�+6Ĭ
Ǧ%`V5�Y��bt��+�+�M`V'Lk�+�+ۦ�4��JĬzk��+l���
��k��aX�cX�X�e`V5�aX�p�p#��\�^��y�UQF:�tZ�׷F-�R�+��7$��O�^,j��۔�aS��&dP܈]7t���4޷�L���b����S
=��P���(�6��iLb�m��P�V#x�(S�5SZ嫷�Hԕ����uR2�2�7ww��rd�m{M�� i���K&��4���qU�НYKbJFS�����Ĉi���i�n���r���&|�J�D2F'i,�d�nl`�n�Q핂��[d�/�r�3=1�Ŕ��Ak��W��[�L�E�h��;S]��Gw�e3��`h�NV��l�[5Q�m�u��'��i�ـ�9�J�u�9I�Z�K�3`�XáPx�����f�d��0܎�  ]v��@�86��5(�S���NE�܂����@d��K2#t�r�t��"�;4p��7)�D*�&gۛ�Tq�)�Oe8P��>�h�6�;6�
s�T���'����Y��0G�i5b��B���[{P�Iab�wuv�sUJW�Gh��eS�Cgo[�;�cd&Ƽ�1�3��hWHݶc�&�I5yVi#7 �Fu�u�"G,SH��e<�4X�H��틏F�K��%=8b�B�Ah��-�Z�0ݍ7 ��ZʙVc�������[(�V�'C
��~j�P:�+Y{i����p��t�����xR��Y�����Wh��dEQ�T�Yq��ʘ���rcmmӻ�[2�-��Xl�r&eCxN��잼�S�i��iH�M��������%<ו��)����SL-j�M�-�5���uS)���Fՙ��v+�P�nܱ��|.�{�j��e@�	(c�
��2�G�	qAD������w*��LX��T\��д�@,��x���ıդ[4ntL� ��e^�m�'&b�Rn�ە(����U���VՊKc��QDf�+�F�YV%*���X�A�����gh[��G��Gͣ�霤�˕+�E��c��;z@�]�����[2�'Ve�jZ��T��\v��ʀA�m����`�37Q�I��L�9����L;[�!ͧ�fs2��E흔r��{#Ֆ*P,��d8�۳L�p$lҬ�~�X7s�"E��b	���f���hWՐ�.�de�r��%��ٗV��u˨m;��������"A\n�+}n�U��aX�4��sc��\��%�˺���wԪkY�2-	5@�X�ٔ���*]�nKw*���s.�{�>���-&�Ųԑ�]q<٧s�@�Z3,U�#�֓�ЖL�Ms,+$f�����lyG.k�by�k#��1ZV��l�Y$T$WJ�OA��
�2�7z����$묽d�i����kD��M���YU�r��m�<x^�f+ژ��EA�k�W�ފQ<�/�Kq��@���ߚ@^� �V�03(D�0r�9�B2�e�H��)O]��f�Ē)m��m;�N-�����.�b�,E�����!߯r�k���kҡ�H5�r���Sb.|��x�p��Z*D[˒��z�VkL���J�3m�,��\z�Ж^�@3v�%��\���6n��]�a�ؒ����<�A�6RI�Մ=S,;e��7c��E܏x&{1�#�!]g4�(����X�����nL�xތ�t�ё��^�����'����#1ܸ��m"���)�*Z���&���6��ӬGw�@��[gYWq�����i��T�H�;ʅ����*M��5�wDׂ�eJz-�m!��i�)�N/��l[)�DJ�B	��qC�����Vћ�(R�n��/Zql	n`��)p��s3Y��$h�HTu�ʖ#+Dv�M����7��¦�Rm%n�B����M�<�Lڻj��h�b�h3~L(n%ek;wl7P�u� l�q� ;%'���mbXUӔ⩇r�a*� '粞+gQ.|(�Z��pAH�#L
3��Y/.��,�C�'�m�(��Q^ne�e��V��t�S�L9{)Ѧ�Ee�A@�t3p�rj���D�/&�]�R�҅l¬���IǮPs]9�'�5}��H���Z��l�,l!;"�	�|R%X�9���v=n���Kr�Tm��v�@�ém�2��le'��ɨ_��o^��õ���'y�b9�e@IJ���۳��抓e��on��	�f, /bx�����R:��-F$�n$��4�S��4�q�UAfnQ�&����C*�8y!ܺn�LJ�:siY�f7�1�*�A�ہ�d9��j�P�"+���*J��E�7Cd�Aj��\�ta���l6[��.��\�A���l82Fܛ{4m�RT%���A3�Aͥ�X
-oBo����j�Ub6�wsU�7JC%(�̣�J� k�/r �!���s3�9sQH�1a�N��<�H�q��L�����#)���L>T��8�p1W\ĺ�[p7I-[�Z͉�PS:Ƭq��*��S_U�] ����ZۧZuI%�GRݘ�a�,B���8Ȧ7Y�z��&�F#�3��k�m�BK�,�۴p�&���/Kou���C�+��G,L��J32����8��x�&��,�]ʚ�2�(�^;��o5�w�ݪEm�qͫ�]���$⑲��훎]���b�̹{,�E��@�l�����M
%1�+T�*�z�I�J��V���!�W//Lq�&��%&�4���mL��)0nP��"��N*6��F3v�L[F��I-�6eh��M�h�znmm,�Y-a�J�>��ؗf��1Gn�:��˒e+�	�oI�Xq�F�[��.��ֶ`n���U��l�Y0+��,�SU�P]��� �f�[Oem� ���������MS�pҪ�&�P�he�7�YYr�%��v��T���;���[B�C�9�hU��廙�FEsQq\�En6Q��9���Z��#s���+B
��}0��z)�n��a$��i	����+2��0��zVn��kUXV=)+"Z��?X��@@v۩F�%A5�7
6��*k��{n<�F�IQn	ؓ��e�Ug.r�GZ.Y�����[����U�;L�lk�-�:&�W$�b��i�ki�)ڑ�Ч�6�W�2̺�1I�c�1%�M�l)e�����2Gy@A6�Jj�m2ൻ[���*�Yd�kl��x�upd�YH;�;tgn���=Yo���pl4�G� ���i�w�d�L�q�u��'��ۖ���X�X�fB�*iTZӺ�C�
[(�h�X�}wp�+
l�/��)�[�U�@A���V�ٻ�7E��$�W��:�Q��o&*��^+����t�Y��4\�Q�5k�h�i�6&À�)������R#mˍ&%�pi0��W
sM;�&���h�O�ƫ��vE�i܃��V����Vݴ4�% QH�ƪg�,]���yC���jD�L�i��w6���h-�&��2�r�AgN�H*Qۄl��Wm\OCI�zim���We�
��Rz������#ʹH86U���
���a�G2�Ď1�d<�t�������ïf�c�=K+"ȣ��ݻDZ�5�]�rⳓC��Ѝ�u��{��ʓkRx�TTE��V]�汲һ�i�]M�tȃ*cF�9Se]a+��jح8�$\;Kv�6vVEl��E�ۡ��'����[
�:�
jS:���w�P;w�\��H��C��,eM!	���(����!�i#�sqǦ��ij��m�AZЕZۙz`0�T��"�`r���6���֕(����T���$_e�u�6ЫHѩ.�s4UEՅj��ڛYb�[zQ�Y��U�E�;4�Q㬆;�J8Y7h�C*?�c/2�;��� ޿��L

��%��:6���{� &��t͝����ml�m�)37v�0��tٶc���ZL@���B2�+t��ȓ
����$nlbaoX;I�*j�܍TW1$���+3��C۲ZiU�ɖrB	��q����\V��E͍�(ZT���v���� dJ�[	cq"v�MN����ۭN;��F^ܻQab�w)�7��f6��2��;Y�܆5l	j��Q<d�߬�Y�T�b�΋15��^kTmd<�e�ů���F�d�Ě�l���׮��Y��{h\*��!�,ڹJEKq�A44V�Ja���"�U�X��c"y����Yj�$���`�
����n�A�^X�3$x�*[1Q���en��Hl��vjPSۥw)���ɚճCӛ��t�ӣp���H Q�oPyZ�8���45V�\�� �az�C�Q�B���Ѕ��������K7k E��[���Oذcn�f��ưt��%2��d��F�70���#�%l"&�WXF�Ȍ^�<��.Ua13v��f+/�VfT!�	 ɫ6'%UF[�6v���ҭE�E%��a]�4���vlFC�]���j��Õ�J���n�ߛ�b�6��kT�V���YM�4[3t�x�ְR�[�]Ê�j(�Z�+�m�;p�*��PH��pxl_���cӭ��w.(#�jgn� +fF���ݡ��3Y�]�g	)��mLq<���tE5L#�	y�����nK��
Հ8'
r5���`�#Y�x��e����a�é� �)V(����l�t���2�څa��Nk!қDc2���\jԗsƍݏJ�v�\��7usF�SWq�XmB����Ot��b�W�����3&N|f X�w�1���ذ'6$�\��x۫wxpM2i9���\����Ί��@�f��m3�Rv�z�:���J*�����/"�OsRY�:��.����݌�e&�NFTɛ�hL'-@▍I��u�������[K¥#yŻr&�&�R�>��1��N=aZ�[�� )��,�;�X�:�8�Ǥ�i{1Te������0�ג���:+Y��f�������O�ʲvcE��ZL� kn��o�F[Ui�Dك�
�3=�*��ݕ����MAHA��`#<�J1�h��fj.]�҉���Zw�y`��Dv8�;[P�ʹ%�lT��Z�"؅h�`CV�ˀ^�����xԡC]f,q�n��p MedT� @׭	��٥V��.Ed�q4p�Q@�kY�H��޽5�ܸ.C���ds�ܨi콹WM�Y6%`ȳ0�/���@��:(�À�;[���:n[b��.�X��J�K�҆����v���i��E��K���(c-��0J�ٮ)�'}�g$���*�'���#��|pq�	��t�=<�����ܺ��7;���*Kou�ݷY�����n�;}.������fc�X*�K�9�EY���[�[G���]J�*Nt!̬it$�m�c[�6�ǈ�ÍnXQL�Y�JD�F7�!��M-���m�Rv��IZ�6��*�%o^��K��b�$�h��J6]]�-�M�j�w7��T�̧@��K.��Eκ^[�HG���Ƿ�E�
u���	�e����y�̌������eM6Re;Ԝ�ˢfâ��`����$z�=��-�밞�W�u���#1�2��i�1u�y�BKa*���2!���	�,,�,�:�N�J��

���/�d�5(> ���^��)���Wg@"��D*��ܸ��t֊��Z�ċ7�d���#]+��Vi��c�D�1vQѐ��B�^�8l̩�O7%`�ŀΙ��I��Ɏ�b���[S�g�>GK����{*
vϕ:�ǫ�9y-��B��(�+�;p�J,�7��H�@l��O�ٛ�)S���_03kMr��n)�Ei��`V��;�&N!���[��[���{�W��C�~H-�.��%�~x2�i��|�_�;{
�8�D;��jJ�n��Ԟ�{�^\��V�=��hh��|�U?
��%d�}��iV3�*�wF�l�m�[��(_i8[R��v�qwX$��N��y2;�FE�V������hײР��VyU�!\۫��H���(#U��}���e��킬*#\W1�Rk4��S��ܻ抩��M1/��C��lY�˘Z��k.l쫩�R�tm�`ӑo#7Z�n�]��R̺zǼf!��x�*���5���ub�C|&v2!a���MB�v�N�-_MQ��i��E�� �T3(XZ�ڵ(`Y|x�腎�[��E�*p��=�
�(��LW�ܳyc��$4�ܨ/0�)��h�$;;qYy����hV"�-�GD�]O%�!�t�w�U�b�`N3P�LE�U�"���;��7J��`��pA��Ҡ�X%i�j�Ѧ&��P>�U�"Ba+E�j;�������	ݚ3������r�\��v����j[��J�V�o66GC ��kn���^�6K�P�1� +Kn;����[�x�ѓ�Ĳ�S��cB�;t`t"�Z�2N�f]d�@��5�o{��!�U��Q�ͼ_]JR-*:�I$]]^%n�'��ε�ܰlTO8	���nD�]�f�%˃v�m��mмu���1b�I˓(-��+b�)�.�"�K\).*\dw�NV���-ɼ�[P�e:�VT���i�Z�R.��PK�ɧQ���'PCz�bK��4*5%+|���I���r��l;��a5��ع�W.�k���(�:���}��M�')�*��N8=�FP��7z[냁��0T�.��X2Z��Q^Cr�b���ԉ����#��2K^e#Mۋ�ич{���8S�o��g�֜RYRo>c#.�E^���l�6mX�i3M+�
�˥��d�=A����;i��%G��݆�_9��X��Du��븻��bޠ�uۛ�����S�ڸ�,��7�ܷq5�M���TU�{,���)���x�nҏr;ص����%��Y�G�%S3�"�ʸ晈�[�6�Jܻ�|�w�&^a�mݑr�%�������t�q�.Gؖl�B廽!�6�)�1A�S���O�����ѫ2,&+$�(
�tBu��dQ����_��ȭ��|���?�C����a�����������Jj�����]�ݵw����X����%�q8���x:�9��!�y��n��z��毻)B���}�u݆Wd�� /p�o�S*PV5b��^�܌�A��w��f���+u��9'X���-���Cg�v^�[ݩ]v����t�P��)*��u�\�]ۼ�\�}(Q�t���Z�J���%JXtƠ�)B��g��Cuq$~�]�a ,�}ک, �?Ε�9�+�d[��1�kQ�v��rʭ ���P����1��[��v{{RfS���c��L�C�`�݋�������b�3�"�]tVC�f��+ V����\��a�D����zn�J������r|���1 �i��o���}I>gn]\R�yNcn����&w.��n���c;�6]P�WM��G�g�6�Z�u0��"ⲸT��pOwݎp�3�o\��2�*
e5����J;Aͨk�q�9T�ST�#��D	+Y�%Y��k\�@�v��E�Ӎ���fi�.�6�Ǩ�=&$mu�q&^��lW�X7�X�E�d��c���g�Z��s�22���۬Ҧ��lG�������IP�7�>�[�8��S�6��>���VN��@V%�uƃ��������9ye���b��K�Ҿ!.�1j����)�R�]K]p9|�m�s�-��SJ�H�ݒ��W�w,�����^�r�di�q&��9����v@Pျ­G���]X����:n
�����W۔Y�ثW�y��l��yN��v�oM0��3���|�ҏrM��m����F��`��T��ʸ�pK�z2L�z�I�B�.͛�/�����>�h՗�3�s]��a��|EZ����N����z{��v1����*i�F3�[u�l����H+��5͇�ivn<�!��|���e^s����s*,�s5��5�����=�:��[�W[c*sn,[��}]�&g;�����4AlQwO��N�����'��4\�A�E�!v<ku�f�[��cZ�g���_L�𽕶�v����IV�5���Oɛ���\���Cz���r����T�Z���Ɵg���q�^��6d�����]X��Y�f'�!8M�Qn�8G0����,%�߲���c�.��C�N��+3���~�{YR����Z��w�z�bF���6�v�}rV�Y�(r�>*ۻ���et�y|�搞��q -��a��]��(���evģ��Ձ	�lZxg$_K�xM��m����Ƹ�l��xb,�#��1	(�NMv�t�y��ͧ���WXzRKEL�Yo.X[�I׃�A>�m�ΥB]�&t1��6�6Ϳ�K�8��7��Z��Օ�_}%�9��4���X��ܕ/�Z箶��:*�Z�
ڶ��nA-Ԯ�H`�c��&澥�w�X��Ղ`8*��#�;���ԅ�I3�����@��H�ֆ��ѫ�p�vI�[�%��{��ż�倄:o)S%��R���F�"���H�{�|���`/j�J�s,PJ�N�"ض�p�E�ϯ^'ٝ�wmW3���|�n���[_I's��rk9�S��;;l�$@��ɰ�iiG��	RY�q+[ǯt�CYt�e��J�[���!�l���u�D�k��W0X��ҚŊXz뷶a�nZ��^l7������WMR��TmҒ��OB˩k�4Y����;�k�QY>�B�%!�2���L\tq��n]�]�����u�:�p���H>��c���';{{j��o�5���XZ*�dp)f���{L������QI�K���ݗ�D�6F�6]{�A{O�%J�U����̀�[סgs�E�XSy��=y���9�.K'&u@$�ZA��0�w�h���]YAb�q1˝��b��u��!ji�'i�xf,Jr��f���Ƣ��KP�D���mS��#�]N��)]:�Y<��C��M��L��Yv�!z�t?��Bڂh����j\����x:y�3w�bFE�#�e4�r�[��NP��y��&"��佦��,�qF[�h�\�$�{9�.�ɤQcs�f�>u��T�O[�E��;�y�ŝ�o��eSx����Zֱ���ˌ#�.H�b��f��6װ��S0�"��ü����.�Ϻ�1�G�;ӵa@�;f��S�e�B�Sޕeu����^Z�����ewqJ�x�)�{���E�0�hJH��Nb��
�Vd�Y�V-�"�.���r���'�Z����{�|�X��D�b�lzS���r�T/�嗸�u�Gj����X9�u�G������I�l�k�͌�3//��lǦ��W��&�)�4�__>�7��"�F�X�R�t��l���.���p�w67(�;)Z/;S�ʋ�m����KsMs���'�w�R���˝�$H�Ø�&�Wиuc@��@�.�0JUҷ�O���T��y֝��{�uJ�ÙҗQ%�j���/S�Ts�n)x2��	e3�]��.�I�h)pR��+4��*M��&:&�漣�T�*�b�n��gj�}4� ��A��l��y��U��������U��]��J�n���:V*��ϋmeK�I&e%�u^.v���q���D.�M����.�D��"vn�%�3�˳�\��=1�5Y@/���15{���ۥ�>f���Z�����H��T�ٛ�\3���=kf���ܣOo��N��z�Ĝ��u�	
��wI��<��kid]c�u����+���և*@D�e18�Y�YD�T�=�̆����ZJYg�5Zv=ȲK�|��΂���:��xۺ�q,{��Y%%w��)cX`����h���*CI��m!�s�Q�!��)Fe�tiX[s��\2�.�P�:�a6�s���Â��]�8.��Wv�\�5�	��.V�+ZԺ��n�Wk�1Kx��{�oA�-Dmk�ؖ��)�Z���RlY9����}����x�֦8�S�'���@W\�� ��bO��v�g5H3*"���jhћ�gk�����+*R:+�g�h\��WAf�7e ��\�r���+{mr{u�"�oM�uEIˬ�{ϸp��+�o����fq�ͣܯR�������s0պ�x�3�ɽ���i������8Nv�9�v������E�P1��M��[
�D����[��Wn�{~J�ٺ�D�D�z�q���A{���2�.�����6�K�Eu�\�ʛ���V��"�fê<�}�f��d"��u12P��݌�K������\R��z�b����`�]{�LDx��7�|r�|E��\Τ&^��M��"�P�/N�;��/�N���9R)n��WB7������8ѱ�`n�oJl��W��k}W�V�:K��m��4��n�{�;u�e���F�)�N�r��R�@Qot����ڕ4;�4<El�zj�>���,M�����\�ה��:���',+�h�*�}�a���r�7�R>1Ü�8�Қ��ߣɃN�+��5��[�H�fv�H��6S�2ձƯ�ب_r*!Ur�>Y�:��k2�:���=��:�0�GO&��ƭ\䛊�ޅHV<A5������ܙ�u�e9���t(��В��Z�2g|4KI]��Vƕ�^o=�N�䓱]�r�_GQj�]$дXjucy��ՉV�kmRfY/�����4�܆k�}Rm\��i$/���{,���.;R�����,�rj���굗�7ӛ�ƊX��Y���.+��X	�77N�Hm�y�Ms2�����m*�n<�A52���s�ok�x�Ӱ��>}��ןl�<�}i�����v��K-�]>������*ܳvVR,n�]\_:�|�M��%-���GsG-]B�罞V�y�����ٴ����;+�@f2�Y:�sp>W�jXx�R�ġW��\�˗�����"��sUi�\x0�9����8��Q�,W��+FA�&��.6a?�V2��nÀu�`+p#���˨M=��Iʥd���:޷���I���H�3�wp�'n���F�:�@SG��s�O���D��oh�j�w�&�v�Zj˷�gS�jr�_n��@�v�vJؔ>"c�Zd`�4x�&���v.#��ۗ���x��J�L��e�&v\_Ip���^�j:7R��t❎�6�8QS,t�(ki�V��VN�WqMϖ`w;5k�Qm��LGg��؄�ڬQc#�eF�Ƕ�\c�i�І�u��'nMz�Qۗ	[u*/�+���q�K]j�dXTZ�l9��) �J�v,ei�Xy!۹�\�b�$L�V����.��w��m��_;�	��Ra܌.	s�]+2����ھyYR���ŕ �kEJ7����wYҁg=/�0�N9;N�
�ιu����6��Sǃ���f���3t�Vė�y{���i�������C$W�Ԑ�4^֫��Ř6�o�=R��7Ι���U���`�2�����XΩ�)p�П0-�&,z���ejQ��H����u8h��E�~�R�1_�l���y��*x�]�;(e��
f�`��`�a͛�t�Qw�,Y�<{}�{Է����f���w9K��ϱB�M���HXR3���h���D�%�h���ek���S�sP�.�ն�]���>{0���2�.�3��+S�U��;ո1��F�
{*zRY���P�8�f��鼙C��a[ĥ![Ҕ\U�Q�
�SWZ۾2q�ow6AȺ�`��o�F���+1�;H�C�@
�������`�4l![%ں�p襷׊�6k�)wvU�F&���oX�����A%�;ݵ�%�\��]�J�N�����G��o�i��ƬҾ�sh�uR����+�V롢�B\3Lٯ���e�ٕ;��!͈ged�]珥dÏ��²T�ګe�]n�'ĺ�W:ݺ��.�&�*��\�0-NM�,�����S�[��y[(�9���~r�t�7��U�7;B�\(� �z��}���z�akq;�����ց}*:YqS��*@it�fC��ܱ�V��{��9��M�%�-�9n�r��ާN*��J���7f\}�|O1K4b����'!y{���Y����]�-�
�1��n2�P��l\o�&H��ƻE�S����渤�H��u����w���9��wqٰ�/�"��)*������:S�8N��8'w��u�Z�_fr�:��J&�]��p�\KWOgg{z�LF��ޡ�A���Z��Kƹ��^U����3��Ӻ
y�&�a��%">'¼ś�d��H4lD�*C�L(��/LW�)�
B���=��QWda��.��EJ�K՞ѹ�x���T�l��+n��	�	""B�d�On��Ն���q�Hl�fH2.��觝:Y҈i0�G���#NB�S�)SIDT�(��.��K*�r�p`�0��M�$�)ڨ�,1Y���d�����U���A�`&�!����I˱V�Aq
�D@d�8��ħw(ADhk#�8�!��a�
I�v��B�$a�S�-�BI��(�[��s�2���B�Z|[�h&&޸1���(4�0�4�-�%
��U�%����U����r�@p�\�Z���̀�(D�M4X."NF*F2U�*������mF�Q��p2��8���U���9%��R�v���M�Y-�� �(1�R�B꽭��/0��<f��)S�#b3�^<�1��iV6˶�6�6�K�C~��ahS��.I�������������<k��P��4�f�Nd���aq�KLQ$��$HĠ�%��/ZUm��@����A�Y/�:��T��I�!�D�.U*��$\F�l2c)m��)J
4$XU�ܙ.��U6b��H�L���H�CeO�ˡS��P �(C%IR�m��OD�F{�'��S0�(D��M���I�����f&� �f�FM����)�R$�X���M�|ʨ�'2��ogEŀ��F	i� JԲ2*���&\a$c(�ؗ.�P�5k�A���P5�pa504��S��L�RM&E�jX�
5�#�6�m3�j�Q���<����p�h���"��i�L�U�;�.�VL�l��f$s�ܺ�Ät�q�i31�$s^��M(TJC2KIBC.FA���#���xդ�"6D�eD#q��="1W��B���T#��Kg���NM���+/��5d�[1 a�P�j;�Ou����)�i)A{�ܛ�VY�
��A�ƨ�)/���J����Sb�]R�f�&�)
���D=x�T�����d�d�#<�h�ࢨH���Mpfcɚf.��9	BH_�ߨ��P?V|��_�(���Q?���O��o�C��T?��	q���Ⲅ�@ �F,:��vU�zS幃��q�@�.�X$H��h\�`��p>���7�)h���l�6�����+&e�:v�-�.r�{@���]�R� y�q�4�%��KLg����=֝�-ۋ���1�GUn�I�Ѕ�f����p��LIԯ^5o�T��ޓ��㒺P;�G;ήLk%�!���H5�k���ٔ���\w�,i�W} ��ǜiN�ͻS�K�JCGt�ԟ>�w���|;oҔ�z���@�=�X6�-j�v��p�$;��P�`y�"n��v]1WQ���ZJ�I�Y��@���f]��uܕ�[e�ڣ�r��Z��K9�˔A�q�#�R��;�oT<�rցջ�;k�der�a�9�2`��Ԭ+��-���	����̚���/R���!����Tr�9$v���M�{-��;��b�)[��$]6���7B[�T_MK^����6�#��+��>NA��z�J�S�8��z�P��]| ��VV�+RU-��pt�ǁk��bP��E�p�4�t�x�{�n>����\q��t�8�n8��q��q�q�8�q�q���q�q���8�5�zq�1�n8�=�㎜q�q��c�8�8��1�pq�}pq�q�|q�N8�;q�q�pq�q�|q�N8�;q�q���8�����������q��q�q�8�ۗ=���ޏw���k@�-��ޏ{Gf��ƕ�-²7M�μ�_^͢�6=�@�WU����ӹ����V�B�y�[oyغ�8���ᯅН����d��$���.!�W.�w���ۭ3f.��Չ�b�,�ykN�@Mͼ�R����0�*��;�x9*�@l���P$�Q�gQ�Pn�t쉪�\��wG��]��oj�R�b�is�M�� P��՗r�vP[��T�w,L�r�J)r�
cܻ͑-�ͮ٫q;��;/���u��r��,����]K����w���MC��%�	��.8^V��{��-`�Si���C���ʰ,X�.2U�.�_2k�v��"���v�1��U��[6���w˃ٺ7*�r�a�z��e����XU�識A�᥵A�oR��f�iJg6�5�Վ����9���au��p�����q��5���B���.L�ɺ�F��9���rUa�mL���V�Z��f��2��	�ݿ:>���BjNts��!꣢|1a��"Mh�u�5b$���&r�Vhw���K�n:.�+�|3�����Bg&���'��$H���
�ñ3� ��κ'~a��o������8㏮1�pq��=8�8�ێ8�qǧq�k�1�q�q���q�q���c�=��;q�qێ8�n8�q�q��t�8�>88�8�8���zq��q��8�q�q�c�8�=��;q�8㏯��}}}}z}q�q�8�q�q��w����b��Z,U�ͻ�X�z�ϐ���F�ջ�O>�2PT���!Jm_�_AW6Cv6
�wUI9r��t�*���e�q;#������N�[��E�����v��)����]�h
nh���dA�[˩Gn���� �sjznj��=�;^R��͞ �;I�a�+�a��qXD��.��lnj��-4V�Q�&�0��XK*��je6*R��>���C�����F�cFf���L�\��Q�`L�z#G��{�y��#u�"�L�_Q�*��W�ݞ,�'\֫l��$q��݅]_j��VXQ��z؆�B��ЍM�:�0��ӝ����)� �iF2��5��ԕݥx�0au��&l����a�����=D� ���j*�U!^������.�K.�G��J���6r�Tu��N�7�x[�n��*7Y�@s��ˎr�&QŰ�T*�K�O��������W����)|�n�)k�f$}v�6����Ju�4"a�&�4:��qYz� -�#����TB����o88)�����(av���k��k����� ���t���ʫV����裷�)W������nJ~|4T�U�9��v�oP�t���uٜHG�����h`8���S]��n�J����:�Q�0��3r�0iA\�kZ:���^ڽBYͻ���I3j�����G�zPT6+���8�s�����}b�Ύ��]������^��#�3,�9\����F��ԣ��*�Hl�����<�5�ێ;q�>>��8�냎8�8㏮1�q��k�8��\q�n8�=��=8�8�\q�q�q���q�8�ӎ8�=��;q�qێ8�n8�N8�8�qӎ8�8���8�5�z\c��q�q��q�q�8�ӎ8�ӎ>�����������8��t�8�9���0^) uU|����a����q�r�E�^��.�ڳ��6����H����nem�A��6�`����m���W���l���
�� /YZ�uθ�/�U�(z����7o�n(�2�.q������ l�Bg�T��a�B�*�>�=��8I�A�M��Hi�TcCö�)]b`�s���u��%-�X>��J2���{H�u.�!�X&D�$�^�ew^��=���e!c[{@�M\dn(��W�}��J}��Ū���'/I��<��E�,��i����Q�)u����m)C���)Wq��ƍ��%�*�2U#��ib���w�5+ֳ-�rG�,
��!�` �Z��T�ĻZoP�َ��gNʱp���G{��Rr�k&>��H}K�+�0[ys����N9VP���"� �m�x��v�� �̮��M�2�(p����T˜��Y˵���l���n�Ѫu.����D�zp��7�_Lқ�k�=Yjp:yX�蕑sS5�K�+u��]��͚��Y��J�����@
��f�QJVM�=z��n���b�@�܆��[*��vpM�gm`up7�&*u��1j�Z:�͢���S���}w�E���ߺ�\{{}q�ӎ8�8��q�q�}pq�q�|q�N8�8��8���qێ8�n8�q�q����q��t�8�8�㎜q�qƸ�N8�8��8��q��q���8�8�㎇qǧq�k��:q�q��]8�8�����������8�㎜q��q�q�}��s�|�71*K����6ZJX�ɂ��R��F]�VE�����m$+��z�h a6TѹiWm`�B�Kզ�!1��՚3�ŗV��h��7ͨ�_��X�L�:S�o_t��S�� �}��G�-�뢺��t{�,�t�{il����u8oT�J�l�Z�zt+'�u&l�*�a���b��yګ��ԭ`c��J6���i�[��3
��3�m�ކ�uvؾ8�P9�q�`��YE�
�2���4K�r�\[]�<v����bS�/�;B�C�S{��^`ؖ�蘰�U��	�����̼�\�������)�������Y�8�,͂gnoSȗ��W[z��Fs�$�R	�=���V���\�yܾ�V	R*�K������ءX1�5@��2>H�]��_��\��k�z�pHN�V(��u��a�u��H7��.�l��L��2��9������=�)�%E謆�U����i�y���V;��A�Ēwd�O�i �Nڽ����A��i��h�蛥g+���+����B����n��Mo�����뼚�S�7���z|}{k����v�8�ێ8��q�|pq�q�q�q�q��t�8�n8��q��q�8��\q�q�8�ӎ88�8�8��q�q�qӎ8�8�q��q��q���q�q�q��8��q�{q�8�8�8�q�k���X������8��q�v�>�f�6"H��|���u��%�uw<��+�'"�!�V:K�e�!��t��7P�S�b��Z���O����;�F3�)�(����,�=�r������s.�թ4�Hܬ����k�C�lM��g��g�����$�P���.+��d�]�3�Nu�0�ٜܺ�ق��jOH��=���N7�|�wxۧ��͸�~���Wv� ��`w0,�ז�M���)�����,[��+/����p'f���;���
��i�C.;R�)�D��x'[�����]v�nP{���fs���
2��"4��4�tB�&Xs&�qb�:�q�:C^Md"�z>��j�T�,3s�����;P��=�ӑ�Wi�K�\�X�eG��+��T6_�T��n :�㨝�P����.T�w����7Ӳ�_c�vp�@�Q���نhţ�����Fۙ�;��5uu����˔���m��X5�e��8.Y����mI��Ǯ�Y�z�]k	u����ԝ�7��c�FT�v���Jf�(�bS{v�cJ�iz�oY55��TQ] �f�Ѻ�t�Fw��Z}7r_c�#��
�MH�5ˣz�;|��O���^�|q�{q�v�8�q��q�N8�8�ノ8�8㏮1�q�k�8��8�n8��q�N�q�q���8�8����qǷq�q�q�\c�8�8�q��t�8�>8�8�8�\qǧqӎ8�8���8㏯��������8�;q�q�q����G���>����
K����v��0jL����P��v�~�,j��r�n]�4������򺂩�gS� t���N�t���-���Kkv�if�e��v�o�ɳi՘��%��p�3GOV����W!���G��$�Xv��Ֆ��וtw}�i�;7�R٬oFM�i��T�L���ͧXs&���4kAn���Qch�o}U�c��{�&�5�}�0���J�l����s�X�J�[}
[�-ȱ<��MeR�va[��e���&���1�5��T�����W1��+��4Q\�]�f��<t��(�E��Y��G�V�G%��D�EJD5�}e��
�y�q5men'=V=Uy �ol��Gd\jZ�콐�����y%Cc�d0`��]8V���}EƄ8�T���і�$�_S|��#5ăr[��vl��m� QP��e��8��Y�����,��^KA��G3V�QwTv�冨�z�`������!wF���w�53�8��U{H/:����VC�^p�����)��q�vz�ѷ�4��`�� ]�v.讒ܫd�5�t��0�uҺ�ynb�i��άcR��x(��oG�׵�yR�j,� �4AA�[�oOsH{r�y�݇�4��]��.m�:����-��	/w���m��ɒ̸S�JSD[gn՞p<�wD����s��&��C��,U��+Ew�4Y:��nC�w�x
t��aKȍ��q9m�7	��s{7 㐼�G��'St�E:��P�dՙiowTf�� )_�t/�W)Y�2�[�R�1�D���]�b�K��T�^��ͬ�?mP�����C��.����P��u*b��4:ݮ�Hr��]oU�FR����8���xd5���WdJ�j�DlZψ��04��K�v�z�p�vtwc���$��ռ�Ś�J���l��i�����,�ҬŠ[�.���R�
#�z�v�X��eJ�*=aX4؅8s�w������ʵԌ3M���C�[�Ԝ�R�`a�lZ-w%�%��`��ӎ%+�5/J:93�o��*ˠ*�Sx�̓O"{$�o](�Y�]J�F�뺲�D���=|�B:��֤ʗV�X�
ɂ����5f��^��2�
Va���-�������6�Z�ut�=�i�LD�{]F>��T�T7�S�Z{�V�U֣f�q7�=����@vpQ�ٙr�z���m<3aD��p��;9ܵ/vG���AJpr�o˴�R7+a�<�U��
���G�͑��)�
�6����)���v�}jHҝ�8�*�Z��Y���N�Z��3����|M#6�vѷ���=�iwv�tu�/u}�Uqm[�+qK���T&-�åq��.��1"�Z�j>�X��w�o_aR���lc�2q��H��"��x�W�Q���mCo6��B�̠^,��	�ˉ>̦������r�><��!I<e��+���Xb�Y�N�G|I�r���{�H*`�y�%��Q��T���Lk��\�R�OU��ft�t�*�h� Q����ʜ�4��ŵ�E�+r��-=wkf��݆�3w��ޡ]"
�bi��E!�o���˹C�P��j����;��J�S���:,�ڴqs7�3T73���z7�r�Z�y�@PZ��%$o9ƍ֕t���9YK{�t�4�bǙP���d���_=�;�R�����O2�^&)o&d��X�{�7���5�Y�<��A(m���|�3Y�y��e�M����%e��J#k-��fe2[,Q���]�5���{9kй��)�њ	[[;9�[W��z];�w���=ko[@�y��e�)ʝػ�g�ʼ�X�N]��z�:��77K��c歧W���腙�3ή�-dHL�g�K69l4Wou��k�����|)� "<TM���1�cQԷk��31����B
-�ŇI�% �aiJ�ދܤ*����U��pF7}�R��J������ 7�vNXh��޵�V)g��2#
�BZ����!�ja9$;O�D`Ψ�3��\gH�Qً8>gp��Ms�-#��u�,!�L6�9m�z�Xc�Qh��'$�m�VJs��}QX��2�'�/(�9��ϳs^�]v�Z��wu"�\y�Y��@���˫m�]�1��x��)�^I˕0�}�\�s������w�kY�����������L2��m�+�ݜ���/,�����m��IZHEI�u9m�k<��Cb�����a�,+33Jy��K��d�]N��y�����x� ��$_��_��s�/�/�?��?d����D��ѯˮ�7����]�AERl@Ԑ Je�C���Dԓ���$"�+��K�˪�R0�AJa����L4j8���/��J��W���9ܵ��%��̮�e�Z��<�����l�K�3�>ػқuT9���*p�%�#�2j�������<d]���6�/���vC��9G��F�c��b����[�4F�6�2��e�Mކv�Ȥ�i�y���u�bY���j-ɔ�[؟!(4�+4J����]�$U	v�����لՋn�oe�9=�ko`��OhbZʵ���Y97H�r=�,��O�,���ѳeފ��)��[W���ʯ�{X�{�+��$�IwJ�eC��!Vlc�[g����S0�pm��Gc�t��N���v�1��%�t�Ӽ�o2?t���b�W�8�xo�݇�%w\�N��
�ܭ	��Fu��ͤ�w:/��SH1)�`=�t�.�V�Pem��X{�8����ⶠ"�@w;xd����_L��9�����i<�A��}� fu��,���u��ݴ���6A�`�ͬ�;}/�wK81w��qD�F��͎��ղk�;+1�j��=�*N�L���2a��깫2�r�7k�q��L��3�ou	[�6�@��6�vm�eׇ0nf4�W"�\L��eH3(8�$#�)�Ko�n�|�	Q�iF�hF�d������Y���*$$A$�!���I� �d����M�th3Q�A���1u���.A()"���Ri���ܲ�)]�fd�mۙ�Yn[�28|�S� \.��9�j*�@��(i�*[dTlS�Ƌ!�X���a���\ZU%���Z*(*�,���{,��9=��&͛6};��}̜��>�~�<�0�DQ���_��
�w�&aC#s+�l0H`����J�}4DI	�ۦ5��׷nݻp|q����	".�H+ )�"j �(�|��CBU@RX �PX(,$�V�B�P����!R�K ��1 e�J���)!X��Hb,��1�J� cX�J�&Pp��VҁmV$��N�������ٳfχ�1��a�Xp�I	9Lgۘ�X-�2�,d˙��.rЭ���B�̷=�S%�j���0jU�̂|����QP���kZ�X��O��=�v�ۃ���>�Y`�h�MJ���9i��Uf�eM��.��V�*���e̢���dfNO�ӹ���������1ӎd���D!#j��]yqT�+���v�3�h���[�UU���e�,�^=������>��t��9D�9:�.u�9J����&T�q5խ��Q
�+6Z�5Ċڑ��3,\��}�0�j�-m�*	[++*��$X�R�*8ʆ3m�Xn6G��j�U+I�h*�C�Q[E�(Q��Tr²��L�m��T*+F�2�1���JU����q�.w���쓭��9��^|j8�0ș,�o�k:6�Oo��آ��U֥oX��Cc+�i[��<��X��)��v2�7E��&9��(�E�i�l�E�)ڂ�L�*r�����&�������Z�z��&������,�u=J���)`[�v��v�z�����ް<�0#^�z��C_EW�D{:��J�o��W{X9��YOd���o<c���ψO)*�@�Q�0�~�M�F�S����۝�$���mb^���D�E�L/z��{�F���c�t65MD�4��j��KjoDӀ%-��PͶ^��i��p�o�B@�����U�j06M��4r�F� ���i� +��P&��58�CEԙ&�kjɚ#H6�I�����}8ݤ���gA��֧��;�7
��Bq�����	§��8��VK�L�x*a������mLyv��s��zx�u�=�=��O��l����<b�[������[���Λ<�g�i�I
˒��~���V�O6`�^����vQ ��B�j5n����t�rS���Y�YNݹ������VW'�Փgm=�ITC�;����E�5�o��y�X{m�]�[0A��چ�j�@��f���e�T��/~mѽ�R0���XG��u�i��A&���~ݐ�U��p�J��x��V����ȽP\��ZDW�*��l�l���bݑ��Ϡ+3��̻���&%iF�Jl�l+^F�q�g,+e)�f�}>�y�'�r�nt��*f>�ޤ�)����R�G�j�;��3�'V�t50�ڛ6�j�a�h)⊸�L���N���A�ʆ `M� �.n����\:�~ |���'je��(�}F���+���m���L�������n�z���!p�%ѐPy���%s�}2>*�qh�
��+��� ]y�6�gHE�xW��[gFkԢ�M%��CQ�yM�T�[�5,�}j}Z���T�Mb[5]ا��^}���:7[:�T�V�V�e݃�0}~�5̥�jњ�6�ؚOeN��|�6��@]����|��{��Xߖ�=�n'Cݨ;�5vX~�"��,<��lц<q���=Nq�SI�Lzx�%�l6�/����M��FgEU�ij!+�NR��ٿ��xSb�cxW�����]oP	����;�V�Z�I�9˄(�R�\Y5(2�I\�윍Ьw��s�U�U�&�L�&F�"�{)���#�Ĝ��d��n�U����|͌��/�:ʞ>�o��}���s�n�
�ыu����UĊ��3���`�}��%y���^��� }�Ҕ���٦�^�:��J����|绒�.o4-=��@��G�x�CU���<}�Ou��3�������O�@�T���V�y-�&}��?WՔ�F�QdJ龼*_O�P��f�pyug�<���I�mT$b�ΐ|�,f�Z�Nt���e`H�-�qZUD�3B��۰��eS �Ty�vP6����Q�Q�U9���C�Wx {D�q;��w�ލ_˵VC��:3	^ָ��`��>jUOi�����{=���{�Ÿk<<�&�]�
���l��_��A���1yO��'#����O����;���.�7��v)�=�RS�V]��7���MB�6�ڐ�3���uȟ[�fOgv `}���xH�!�u-��+��i��Fl��{���`Õ��r	�[��ѡi���hr���uĥ��'p��+ﾻøo�����[��{��:���M kR��R�TZ���A�][ya�{P��	�b@��z�$�q?<�ha�Y�<Nyо�:�"{�I�F�ATK�|����ơ�ɫV����J�f��S����kw+R��JU>����]\ǭ�Մ���jh��,쭳��>]������Q/^|��O=5oދ�;��~o���d�ח�����'��+_3��VrSf���|������5���B&*���-UA��ez�
>�T�eV�'$6�H�q�z��}Xq�)��Y&>8L���V�yW����y�|���ܯ��D߸U�݂���V�R�*�ְ�L���Xm��L�nP/j�bI��Ѹ�V"6��*���x�x+ؕ��r�S��+h��NοO{w"����3n�t$j�_!)F��5ٛ��p�5��\կ��$�f��b��E�D��Be%�pA3�'z��([R=j{G"u���ؚ9Y�f�[�s�mJj��n@�퉳���=��x9j�����Һ��� �h��R�P0f����.�)�q*f��K�K���D����Jj(��Z�,��&�|{�`�H�����`c9� �y��wҽe��V��\�NC��^���4�UVZ�0�	���o��R�`�\z�+nt���=v����!��ﳞ��(x�E��V��Z�:{j00-�ѕ�ּ!�w*��z�N�Y���ʠ�k�=�祿J;��yg�gxu���5*�f��5~���J���3�t8��^z��h���ԑ�)���2bg1,� ]��W�rJ�f�y�˂�ô
ܿn�,�L�9�k#���X+�6w��t��Delx�e�nS���e��_�䞕�is/xw!a�s��ή+��k��?k�x��vq��l(l~��|@��L<#���}�^s(o��3��+>g��몵�蟢�ڸ��>��*�PQ�]e�R������j��j~���8�-ҫc>��Ό�v��� .�����Ȫ�'�$�^�+p1�ӂ�tfR�`9���;_
O~����<�/.I�5�ۺ��UՃ#�Y�m0'�y��x�`�9]gb����;+^�
B��B ��Q�s]���@��V�
׊�6R�,7�L�euD:����x��.�Af(>)�JVǰV�#��L4�jAFdꭓ�m��B�L��[S���}b��[�Y��f#پ����a�N�r�����n�E̋�6�*���'픐.4�an�ɟDj�3{-+�S�}�;=C}*�h�ߣ��v������g��@���=那��2|�;on�M&�RSf��R��[>�q�#=����_,X������&�6N�Z�^N�o�4���'�Blp��ϟ�]g�y�k�����]�Z؀�f�A%�kT�J�z_��L0��]/X���78����)�7���o�FWH-����H+o�P�����>�8F�f<�h/� �B7F^ò�6`���X��1�Ѧ
��g��Q�(?i�O��U�-"�|6��Ť޽��3���%^ ��n&�]L����@b�{}[n=ZW�^�(�s/�����v <�@" qC�)�[�ɘ����-h���򨕾vBp�R�X�O\)r���t�W$��$��߫�U���8غ6I,a��Z�ݖz�ש܁ w�Ӌ7�=ˁz�Z-\�w��<�6��*�( �eǖ-ٿPG�Ӡ�5Ty���6��UH0F���e6\�-�2
	�f�0�'}T	�f"a�#wn�\:��>�t�n�hF�]� �xkv)'�&�2�+ �&��+��U�ɠt���c�%�L�^�e�w�e,���������h¼���ǯ���+7n�{1ye�)��94��e"|uW�R�p��	�h�t�llI4�2�>�(:ey-��[��X�2��އ1��P�¿Udm��SU��8V���
t�ŨPgE�t�F����;�J�{��D^y�s[m2Ѿ�2��D֩�\�ͦ���־��`��/zmC@�����]K4�T=%~�+}�;V��/h�z�{�X���"�>���[��X虉e׎��)嗪P�$�Vkn�ᗸ�V��Pϐ�vL�����˦"��G�2*��sɴ�jH�fE˳���ld.�G;_zi�v��z$5$����i9{h�JK�ns͆V�:��}BZɪ�$��^h0�U��l���y�e\��2�V�[רuax�x/t]r'�`-�:�q���ײ-d����͋f
y��0w�;��7(���)��g5��T��ق�S����`�
����C�;��r���P�0�p��-���@+��g��s7z_� YZ�7�u��ןH��GcY��h �l�y��u_��]��~��'�N�.����"@���Ru*�UVl{=����0<V���6��U�F_�Lk�x�}���J�bY|�m��g7z���^fz����%�3Qz��|W��M�RE�\o�D@���D^�7�Մ���n����+8BxR�50����dc �f���}vu�ה�O;����vO7�d�2�<NKy��O�{G�*�q��A�����}�3I��,�}��P��LJ�M;N�Z��GL<ˬ���y7i�+ȅ]���4�4>�e�� xCd`B&s5�q8��35qǘw���7�b7U$m܇Xl0n��R��&��5G���{v���h[�&#��sA4U��.��]0��D�l�}�Z�'Jn]]#S̤ر~8��,0؈�t�`�ػɻ�:o�r3�Nqj�H���r�;>b��udƇ�X���h,RW��ihwR���N�\���i��z�n5����A��c�(�hҚR�R�g�l���3{�:_1�}*i�B{!�#.GoӺ�W}�N�h�F�]��=���u\�@LTQ2�+ڸu
ejMJ�/��C"�<ؠ8��=>�,��ys6d�~�{������f�	=��F^�E�փ�B��� +���43�v���h��u�Q%Sd���E_OHFm/��H�ui���������*�Uɛ���i3�|�vqV�ܩOӺX�,:
�8r��e��Dz\��8vyI䐙]w��z�{(W����J����6��UQ�k�UT��Ͻ�|�n#�2��6���7�u`Ez�8�����p��W����S��u��]�2���%KԣƲed��x����~�[�p$ӻ#
ݛpe<7r����h�  ,S:XM
��	 �A �Gb�]������}68�O.IW|��K��;��GW7S�)h����:�}�pHM�z��U�B�ݼ[ws^�GI{��
����r���+_qM]�%��S&X#Ga��;e&k
�ݝw9g7�/�. �=���^�ΦC_eUcC��/{s�c
�PVz����˼�l��("�i�}�7�%Yw��nHܠ'`>6ߊ���T���y���^M+�jqš�"^�U�(0�	*5��Օr"�Y�ٝɃ ��$�X�jp fǞ�,�N�ť�uY8|�㶯�v����y�����{*[y���pt3�%�-8�p��	�;\�(מ�L�>X�Vj*<���͙�v��U�:��O������U/´�:��w�#�!9f�^�*=�A��%�F�22��:���m�	�0o�Z�(|�>��\���>����lz��s�����œC=�^�s���Zֵ'��t�u�*s=C�D�΍��3���.�6e�R����j;w_��r�c.h�s�K����(�N9�6���T�w�Ţ��O.:њx��9�z���Q/�{��+zg"����3��څ�����}�)��Tg&��o\k�Y���w�T�e���9V�{�n-;������7B����9��uH.q��.�R<�{�rC�FgP\��2iܲ�q\2��M|�GQ��],~S��a�<��ٳY�M*�U�M檹�y�mƏA���R�"���0\�����p��V�wQ��n�8��ɝJC���8G���S�6ȥ �z��C4rv.-;���j5�Y4�dp�r��鳋p��E���r�T!�o��:s6��q6/�mmB^�3��5�<o���:9-�g��6��,J�s
�sk�?MJf=�����ݲ�L$h�28�[6
��i�C#�#R�!E��:�0T1|����Gb�c�Ga��ۅ�M��o ��ƺ��Mou�=�t���A��DA��YCΞ{מm�-���7�(�v#w��i ��!��5�7y���	Gu�fk���pwG� ��PTJ����o��`�|+��_������s}�N��i�k��T��p� ��4�6c4ER#\�E�s��鵊��n_ɢ  �e��9鴝��3ؗmuT�+��o@�GuP�띧����%ۂ�
[1�d)���(IC@�2S�����Gt��k��&�*v���`CM9��N	�$����n�AXiv�Zl~b�c�Ҥ~�%�B��(׊�HX1�iS.duǓɏ��󒺓|wvh��L��t(�]��EO6=#�pte�.%\�!�|�Y[{�t�AK\6ګ�K>���ˁcO���Q/���uD%3��iK��޽�IZ�1;:�Ͳ0�J$��/�Y���XR�p��Ǔ�c넚Zyn�����ˈ[y�ݹɧ��.��3�^L�Y��BS͜�ǝ;�rS��
���j�׫%����Q.�ꚻ4����)d��/�����}]�X�i*��^��	,r�	�U����;�ѩ�&��n�/�Eitu�7���nYc���h��U,��[l�����_lSb��R����%iꤎX�l���ga5-��٫��iPfl��179�٬�i��kF��-nb��W�ثy�sx��X\�o٭�{l�.����U�2]3wӝ�3���A�� e[.u�,08��ug����Z�8ahξ��[4���s�V6o�`�d6l>��.nWw"IG��[��]�[�����yy�<��gv�am�����(�
"%F�D��刱j�-*֩X��6�Z��(���Mi�Mjq��ӧn<{{v�����ǌ���ﾴ*���)ޔȈ�ʩ�L��Z9L2Tm*�W˙T�:�:���N��k���۷n�>��<c;}�FsA�z�����eFu ��"ʩEVT�q�+"��c�Ur֢�['&K2Y�=��v��}x�t��$��&�騡���X,F����������*QR���H�+�u��==:x����۷o��=1��{>NKg�τF�am��LUDkR����2���DjkQ9։�Ƿ�n����۷o������fOf!}�i�,�%@P�ܶ��
��U10`��h/2��z���������۷n�^:cǦ�{�Xu���a�3.�[��G33"�Y�!�Eƍ5��km�j)QEf�T>�Ƥ�x�R��D��)�}`6�V�r��[l��ˬD=�uƌR�ZU��E�	FV���"��*bӊ�̸51�!_[��ե���ՠ��L9��B��<�*)�S���dD��Dr �D�=0Ռ�������4jih�,c�,�t೛��e���K2�*nD�������������1�ht�C�çEO7���S ��N����<�u�,᠐�;����u(�$MN.o���&�����/:��w���p��;p1���.9���������2��c�[�om���Ѕ϶t�E��v|w��A�dFC�V"�U�����~u�������~ |�8y9��L������s�\���{��>@x:����Oy}'/��3�y����3iL.	����7��9(S���c���%Qk�C�Q,�>~�����&�j!RH�R��8�A�[ď���|�����(|�/�Ҩ4�_m�6�ૌw�.�����z��,����j3�Z��0�2`00�m������@{�	�]�"��u�DQ��צs��wV$m�W���xsw\x)�<Ml�o^���X�{�o7�(��l;�8�0��l�wN(��\���'t��p��������0/=���,/
S{Xd�J���om�r\���d3�69M���{�sO	b|��=�è�I����>˜{yݴ��.���W9%ux&�!S6e���;�[��o4�@�n�m����S˹��C��/lXg���� ;H���`v9��O�zttdM3�F=��{G,o4c8�_u66.��IК��Ce+C��x�ϡ¸:�Ƿ��|��r�^(jA`�@Rc�η������v�a�y��k_k�.�� �;�v�̒ou������j�5Ü1{u���pk>��ӭ����=��ʹ�Z��>a�܎9 sr�f���\�I���K�|P:�=���I�K �n��c�5���ޣ���}���ON���\ _P�6xJH
<{Ϧ �O4����3�߾��p����y빞��vxK/��$��S��ۧ�@^k�d�[�n�E�����K��`+<C��_g&+�����N_��cWJ�$��C��~�[˟��1m�`$A��;���4��H*�5���gu��@���g�׃�5GMv+����8xf`h��|o��[�ʜ{�����Uׅp<���
`�o��5��-f�8�i� <�^Oʇ}��w��I�������V/���ܖ`1�{�F�XS9N���}F�oG����=��,`C�C��ϩ>�̀9>�a<2C�d�<s<�6j��������N��g��;e����=�ze~��"�>���<6����a���b��B,��>�~ۧ�y�",qݏ���r�;�y����Yb���5)����v�e�)���&#.t�����mNr#υ�oaa�΂�1�ϑ���L�s4^�\�x��բOvUs�ꕝ��(=	4�� �=�\�p7��l�͸��Y�F�b'�&�NJ��X�)A�u��p!��utV���vϰc$@E�7��
�q<)u8�q��+�)��٢�\�:L���K��::�؋��w���'����/<��f,��$A����9r��*�u��Ѩm�X(���{h�qu�L��eҙ�q,����fr�.s32���$bF$gԋ�p���@��]�_}6r �#�@s�n.	��sg��3˸�5��@���=�S����]9��};��v[�eFlr�z�ow�^���a��\
����d9h|�Y��Jѯ��Ƽ9�	=��<��̳��gD�����.�|��/i��Y[(u��k��u8����~�Cơ��=��b�)�?~ϼ�p&g�	��_N[�V������9�y0�;T�\=�K�Ǵ{�.Uᵕ7� ���W�=Կ>!�_`������:��̬�H��~JS $l�`4���`:���o�=U��b:C#!Q9��oȍ��]���l��;ώ}��3M�88zg�˔�z1��� ��oOx���� kΛ]�"�Y��3xm\4.'�'}��������������g�b��ocrr�[��� �2֨���A"'e�X�am2z;V(��?bc���]<�=��� }8�i�;��/b��{�-�z�����A�rs��$t��-{���$��d����v�?w����!ԥ��0>�ŶbS���{y��8|���������
$�ۮ���צ��� �s�m��I�C=����(_�������L��z煲y�L\�]?I��/������;M9!�i�Q��N�!λ#k ml[Ȳiʽz�.�����|Y��y�=G ��k&�>��&G[�:)��A9P����b�V�C����E�M	a��h��rzbs����v����7����D����Ie����RO.-b���X��0!�<7�x�j�4��HΥ�K��9z~�������5=�|�1�v���v{z;����u�@1���g�ǖ�����0����Q���~���g5p�v��<�W��}\�����N�á�txD�Ǻ��L��jwo��p;���4��<�5�e�����`��l�vGyM|������	�+c��s���u}�o/�v2<!��9;�P�h&�Os�/5Zn�sF�	�e�Í�e�	p(;�s�%f�q"k��d�����q��4��W!:�<I�պ��Μ+=ة]:�� i謜a��}��T;�@Dw���4ډQ�k�������;��Y����Ι��Ʋ�t@�$�3�{�����UK ��`;���_���_v�x>�U���^4y�T�]�Ag��8:G^ӿ��̾!��f�dxZu��ok��L�tz�[vҠ-���x �3H�c] �\��"�< >`���[S�;z��YnFK�"<��� Zf�|
�a<�y�ǣJ�.^�����[�����{��;��g�/���s�X��-|B�PC����4����(���+*��=(��=��Q:�3{h���h�K��ׇk�-,�+b,����M�ۡL;p�ǌ�6�{���={u��t�˲K�A+��<]6@������|�R!֝ʼ5|�w�:��鲹`K��nE���P����2lι���Ӥ�����A�
��5��y��� z=���vm��e��k�-��׺m�Y���^DͿ5�q�zξ@�Rت`��ͯ
i��;�E���8��d	��z믰�T��9�0#q�|2��d<��=��>}���7���P�9B[j�_����Wݷ��=�m��~l`+�N��r�>0�y�������O	��<p��4�P��ΌHhz������-ݛH����np
z��k�,�c��n�bNϳ���آ�ڶy�� ��k85׮{�}��R)9l��5�����ߕ���0�3��6p�Io��t��͠	��ʀ")h�l�}Q[�E�Z	p�e�q���0���������̱�/���b��<lh�h��|�sQ�|w-N�Y��^Z� "Z`I�2������;ə� ��>M�>>hj���{o09���TU����P��F���`cW��
�fO��Ɗ�9�дV E�*{�����n;��*T�������7��ے���%������w�DA�;���x�Ă
��gջ�6���̪�S�����������c���TʦV���;ُ���~z�C7�E�3�h<b��Wq��Ɠ�،�Qe���׉�}���u%���] ,����ҵ���j���+���1,�b�t�l�<�k��Tѽ�ug���֌Zm5�t���W7�.�>�9�ʺ�,v��a�^��-YZ��N ��R��B��M��<9k����@�g��Q��_����O���t�=��gk�}~�U/|�H��:���Ȧ�O�F��t��~`a�;������8M���Z2���or&Ȃ��5�����l��Q^Q���쉒/*��~���<W,w��@-�5%��џ}��i�]Кy�5�2�N���s�.9�ʑ�j�7X��ٌ��鱻I<�/�yC����4mY�z��voc�$xl��o\�{�\hu&�0��5ڇ8�id��="K�ܷ�i���?�[�p���_��0����p�E��զu��_3�]�׉p0�YD�'���n�Y%5K�����e�^Y7YR*���o6Y�ߏR���{y߸��F�� Un��85�ңb��3s��Z� �_[��r���cT����͚fE����wuQi�mͨ2�`�v���IC��&�9�˻7l�T���c͌�rΐ�L��9��R�\�WK���׉�O>^^����T�<C��	��Q�.��|S
��i⾬�vy��C%����U0s�����ͯ���Rэ����;/f�F��uN�(�{]�Z-�<�ww���mgv��<h�h�jED�Ѝ����)V�]X3���H.cL0�")ru&�":1�lCjV��	ZtM�1���Mޞ;�{ys�������Y��/�����w;{ T�/��Jfp���@��L��&f-�騙fkwn�?�e�4�DHČ��%�<����y�]�s�u��BE���L\�bP�(�u�Ů>5���(t���[ǟ/����WC�Nu��i��s��/H�~fh��h���"b��X�)��^h��Z�A9�����۞�ã��r���zڥ�n�^��v�~ge�H/¸�����Y �J{�����o�5X㦙 �����G�񢢳xg�ہCo��g���@�/6�p��<��2�4A��.�w}<���W-7��8*_c5��|~4C��}�Z�Y�à&g:��pu�CS&�X�,;ҹ�7����=����5dY+�o6�;��ZM�;�_;N�k~B}���0S�G�?���Ka3qy�O���m�/>�ɡA+�1�w�03��Z��]��Vy��u���P1�](x���Ι�E	=E��C�~喾�*j�Ү��z�\:��t��@E���8}��'�t���ޕ�D�,��n5��p�2A3�$"§��R����ڇt�w��L;�\цom���[����w������a4���Ӭ�fd�s>0^�~�}p:�����NW�P��ݡ�� �-��u�&b�ս���4'6u�s)������9
͓;2�s�#Ds]�D�W�:�\����d��ɻ更�V	\!��h}���[NmtFƛ��`�|�<���c�foJ�_��� �w��H1�A�\�ϙχ��޺�}y�Sl�>���{ U�a�w?��r�&�|�b] S_�����~���zx,���2�ק��Oʫ��@Ӱg�"�_;��w�߫���B�����W[�X�Tw2p�Z�>gX9��;��P搔[sP[��@����:��`�a�����6�Ƣcw{wc��:\��3v�/�9?y=��KN:��	�fM�����=�$F��v���t�����
ch_hTZ{~��I98P���t�{��S�x���iۊh�U�<�2$�w�3�0'��{_��TFE�X�$X��#1���iW�4�y�=��o@��t���k�Mh��<�}b4E������v#D�"&8{S趰_X0���D���a�8�W�(�}�����1�0�`��3��]��#b+#y<�;g��W.��&�$����=߈p�5��K>��8���ǼD�j�Y3���SWa��q�@À����i4��]�+���i.�l�>����|;�����h5;��#c���mـ�et�NW��]��~ow�%94�@����s��6a����|wrx�U0H�)�@��h�K3�%1��Kv�\W�,�@���u��Ư=�0U��//\��FD�"��˜O�`�� ��2�W]ӳg-��U�T���R����,M�]m��;nÙ�8BY�����]�u�@�!
A��b�=A��Љ"!/gy����>���M?M�,Έc�oT�u�M��wE��ȱ�v�C
 � �
������$���ﱐ�0v�;�!��.1��V�����ﾼ���~RbW�k���f@%���Z�8[k:ڟw���@@�H[�0p|l;z���PJ
z�_9k� 9~�Z���#����<����<�{��胝pr~��{i�-C�|y���6zN ��پl�-��67-Q�S/C��u*�Qa;M�<�����{���x��yU.�����m�;�ak��v3۞��)����?Ϋm^��O	�%!��`��G{e�
�ر�Fkϙ��nl��<�0S�~j��lm)�s�L6�&|����c����&�Ǩ��5�w����9CYE�X��Y͖M����-h��q�����4��G5s�d}�����Ɍwkj��9� /�; �5ٵuo Ԣo�fQ����i􏚯 �ظ`�f��,?gϤ��ೆ�܎OGa��>�N)6(q<�j����C�＾��cg렗70�o�k��]�p�O�Xm�mB�����=ŷɊ�d���f�c�ɃW�6-n�+ Y��pʻ$�3�j����Q\�0W����	�;!p)+�W?���{�T���Ԝ��J�V��0��c�g�!FIfi��fA�wۂ�d�{��<uo�X��#	i,�1X1@5g�g>|θ|>=�{#>���Z��Á&r�Ȧ�����>���]�F��.oo��gC��ɝ�}v>���H��;���7n���q�@�u@����}�D��U�5����}�����-������[��<JĜd6܄=��c�sඹz�'��群G��7�j���3ɰ����N�x�I�"\(Wy��x��,6�����覶��ƿ72��U2y]����6���YpС�1��[S��;�����|���t-�s/�+਼_�Rش��Cy����/�k���v���@��w�_i�栀���=|����&L��6�"�*\0�|a��'�6�^k�ת��2f�Ҋӎ��V��7O\NS�o_)r�3ނ�i���[�/�\��l;���\�#^Dpե�eL�.C"ـ��M�^���U�MY�(d"�m��DY?��|�i��V�FC~cr���؏EbF�A�Liz̷�a�,�8J���&���7�q��ճO/�����C��h���%���%�K�ϓ�R���o�kDf�kE0@䵾Gg�{|D�$�S�������!s���|e,�Z�7��ԕ�]�����{l�.s�׬gl�2B-(�]+4��N�U.����<e�(�Q�kiϦI;�.�U��2,�'jҭ�5��r�ĥJpΣ�ݾ��7�	U�h2����/��a�G�lQ]��.�F�O��qLUҝ�~}��Թ~z'vI=z�֍��&CU�;����|��
����0�moR��+7��(J&A�p�̓Z���4��֔�yn���[��٤��hc|�.�f��ڌwo8�$�����V�]JKT#7�\YA
�m��̻P3e�� i<�3N�m���v��˗��Kq&`o*59�;��n
/ɚM���,E��e6�b0Ta��N[�9o]I��]�#R[��^�՝3@+��u ���ƶ��Jp�_�G�6v��>�I=�C�����wn�U�K����� &F��ޛ+sb����εYҗvk�ْ9���ݽnWK�J�yR6Ȕ7b͈�0���e�`��3U���MN�rBn�����+{�Sb>��k3 ��דNK����P�s�E{�+_�r�Pn�c��}h��(ѹ��,�ָwN�&��,w�ݘh��J;�M��5%*k����֤��+�p�r�P7cU�����(`��oD�.���D�e%`�×�R�!��ׇLxTJ�����V���Ve�B��<,�Ы�]x�hu��i$��"(�E=v�B~�8���a[��J`�je;V�n������0�,>q�XҐv���D-!�㢍`F�&V,D)B�-�Ia.l: X�}�ةX�JG�X�/�m�������{��>�Lȫg�����5Ɲ5}AH�8�0��!g�w^9�_=�͘�ɸ�T�Qg�f9���:�ܢ	I�cu);��gA]1�Hz�p��,�&���5����� ���%��ӗٽǀ=Y��u�I4��ê�J�WMo�1��o�J��t�8�&s�������b�%������]b��7�l�ۧ�RK�G�+{�n*/�;
#-f��{�u��lN�9�9p<'(Or'��۠�Г�����d�J#�i����f�0�m���u��;�C�kT�em<�:�_9�N���{5��2�K��b�����uŴ;�^M��+:Z�ż�8�K��>{M�.�u���d�Tsr�G3��㰽ɢ���Y��v��RV*�,a|��{+�yc$M�R��d7k�$|�IqSj@S���o��f��MNXT<)> �+�fp����u��N����G	k;oc�7�9�<�똸y��U��Z�X޻;'Cn�py����6�K��Ć��Y��u;/67�8��;����%�2o7]�|�s��{o�:�N�}���SIc��,�|�]1��M��u�{'W,�:#��:��b��aA��5fE��	F�h6
1!W�B��q.2�S��[˾��^�sa���Kc�3�2ʦ�`2��)�D����q �4EH�-��h&g���-��"0�N��L�	�Q4����`�(�f
�mD�Pp7�-(�"(�I��N�GI(T12��Ib�J�d
�RSKWc�����U�ף�p��=g V[k5�fZE�Z��&�m���Bഢ�������ON�ޞ>����v�q�},e�OU���`9q2)���e(TS�11U���0�h�5�ON�ޚ����۷��:c���QQ��=�5�&2��
��UPc��e[R�R��N�ֻ̘x�onݼ8��>�2I�Z^�X/���S�f)��AT�DE�d�`0+F)�a�����{v��ֵ۷��:c��`A���g���m�a��ى�i*�����*����&M��:kƵ�n�G�<t�Ob���H�dY��J�s��K�+B��q��T9��.�{����;'Q�q���������k��������;��[@�5�Z.�+���izJ�=�Z����[��x�v�i"<��J&������Q�P��QQ��E�`���1Y�p�
"+l�]��kTU++SY�����q5& ��\��R�YLs*�. c�*�V�Q����Le�PUW��+DXW2�;���*(V��%)�u�;��È�	I�A>�"D�,�m*[ό�q]� ��9[�&���X�+b����!�Q��x�+�:�n�'�ލ��;��Q�KN�
�~�(�܎(�"$J�6�N&I"(�n�fo7���s�HO�`	D�	���
��}�^s�l�� �й��1&����9i$/{�w�];;���y�;�.Zk�>�}Ź,é�(�襤�C��L��C9S	�K��cI�D���/����yVwm[2�/�(���7�u�GSv�?TB�^�%����W�s�y.��޵Y�~��lDA��C�1&�ޜ���K�����p�N+XW�hJb�۬k�P/� �EU�P/>�ɳ���}�_�B�����S����w��{��XxS߸�P_�~>|!�c�+L�%�YK�Ǆ�|��0w��V֐��o��`��{#V��A`op�x�z{���ٴ4g�!N{eL䞚��	o� MT��s|>&�;���Ԑ�yol�	z��.���Bg:�;�"���P`��6�$���)�q��o9�YC������N�s�낒��3��=�i�t`�y��q_
�â���o�h^�ho���L�߀���l����}wgh� W�q}T��U�hޡ	_'���^�匜z��so�J��&9���Y����j�9���C���]?5���
y�xYi�G�,�ϐ&�R����i�|��	�����KMv.`'��J�k�[W�G�Noe[��`uצhY�$��[]��vsOk������� �Q�>�t���� �7��2��{{�k;��V��C�N}."�#�t�b��ӥ�HnT�;4,�2�Iz��]����坚���"}�CC`�MC�:=E41 wv_���Ϛ�>f��?tx����켡ʢ��|w��p��������6N�s.�v=[����$8cn�/O3�ޏ<{<b��ՒJ�u�����u�lE�}l��p�K&��Qk7$����xw�8je����xbX����6c���jtݛ�I��v8�T��FDQ���ջ���ov�^������.@�C��r|����y�>AN	�t��!-^]�A�if�m��~��"r2��"�O�v~w�喻����y���^m��V����>������i�6�g1���z��������>��~��⺉�Up�X�|z� �wm�#�|�R���3	�����|7�o�u�t;/�Of��$,e��� a�.b�CUi�Qt���1.5��P����>��eφ;��~��7�z���?A�JN/^���O�Sϕ<J����(PW�N8��_}_uR�j��ϻ�9������W�W���J�'ą�=ʮ�ϾLu����	��i�Թ�*;�Owr�g�͐�L&�s��zc4��Ү���.%�(�+�o	��4>{w�
���������~>���wj{�J	�WL��Q���J)
;W䨮V��������o�ZB��;ޑ�(�V����>���3b�`)��/�ѣQUU1,D�l�c�I�%j�<;Qm���u��=��o��jlɍ��� ��ʳ���:��S��[����]����0A�<B&�
A��`�@D ����{�+��;�T�B�=3K�J�	X g1�-�yM����0n|�iA��vL�g�͖�������v� ����z;k���aK�
-��ӄ-T��g���>$��9߷7Z1l�����vӷL@�~���^찟O���w!'=0�*�
��o��Kʘ��̞�ϯ�r�Z	���9/�ns�����㳻	�U��s�M�3.�D��L���(��7>Wu�~�j.���(�l��"�u��3D�L$�K�pq�R%���c9wխz����PB}�Umػ+�?DS�x���ֶ��F1�zg�P����GR¬�����,|�@胯�����ǻ��4cl%7.iږ�ȫ��D/{�X;!���(Ϡ^|$er�����q��>�V�|��V�_<��ZA���51���=;�ozmԯBn���M��|�2�Ǩ3w�@c��3�׵�����B���U9z�����k5X����D��^��cN�����=�q�C��|_�y�=՜5��jLH���<�N���9�'�p bۇ81�a>�}�,�
`B��������x��ǟv��o�xf��f}�Y��2��>W#���@Uv)�t�v�K�ex/�M��3*�)wgu?����PD�K��@�"<��{u����iwc[Ū�S;��l��)�����<{J';h*�)�H_7ݝ�v��ז���@�$ D:��� dMG��u;�"�*O��[|���훷��:��ڪ�;Jt�O��Txiv��t���d�/b]:�;'��p�;z7Gqu5/̹���P�qo��s�􋠎!5sb�sv������a�"c���8ϩh�-���W���R(��M�i?��=�41O��(Lfk�@��I������|�G`����q�,�A�I�?x[O1�����M��J�Ϲ�4oJ&�ˁ��B"8��u��j;�>i�02��nʽ󍬳��j��xZ}�Jԝ��֨x�LI���_����x���Pz����.��ԡl����U��H!��p�g�CJ��`�n�a^�y�R��څ6%ͩ�n�Y�L3Y�u�����g���������P�G�3E��us�t�|����)��9YE0�ރ+����p�t2���e;��CO	���n}>��m04�tF�dʗvݷ?�vЊovM�Ļk�='S�nYv�u� �Ϟ%��^��ju�jL8$%�A�ʠ��񍾡�>-�{��Q���Ƈl�=�8��z�����#�;�yz�q�!�� ,r��vY�O�2ׁ��A��3T,~dۼN2�(4�z�ò�hU�ʸ{�ɝ{Ϳr���F�6�ޒx�����L��eR�l�T��[>b��%�*�NDA�=�����M�H ̅@#!� $fwfS�˚;��L�]�s�C����)��랟L�Yjme���9ծN��&��c�����Z�z�T�E�dA�H�:RR4��^���^Z�w�@a��-%�40  �D��D�P{�y����ap�@�����4	���S��_�ާ�yh���U}��jy v��g/���Mw�q/�_N������`�b�d���!�22O9�25*ڋ�5�	q|7X���|��M���a�kc�㡬9���r]��Eqcü�������LF�qW.�3�^���� �Y!�zM�����9������i�}���vZ�B~��p�Dø�h�-]���_N�Aj�p�{��]�ԧ `n֝6[}��������?sا��/S�$S�Ia�q��ݞ�Z�g�:�<Ț���G�]�+��Ϟ>s��4H�EX�`��*þg^��~����	>����
Ip����N��w�u��z�R'v#�I���	VCl�S	�'������g�I���5!���'VIA)�V�o��@�������3>��>Ւw^�|L��5v��ώ w�L�돇����L'`}2��/g}L��F@����t�3_:�\=<�¹�ƺ���ׁlh����A��I���q��p ֠��Ǿ{Z���U$z�|'�Qf���Q���������(��O-Z�7�T��7�ۺ7�"��8����*���Z��3�>縞~���~���_�^y���(���*�������ũ!�uYn����u#\N��V� �1S�����W��&����k:�/Q�Ф��J˻��LFf�aX4\����f���[�w3��T>�
b)(�b�
b�����y��>h�Z��?[뿬!�7���_�1W<��� _PC��^�OY�M��RS����$"�aX�<</�o��6���Y�s�k��Z��F�͞Y�>���
,j��^���}>&��;�]�aY�;���k��d�Lv�e�"�}K�j�����*�5��-l���[;t^6��J3 1�h�%y���u���{�چ��0�q��͜�&�^���>�[�6��m���&kr� =l<�Ҏ����7{�j}/�v�v��ru��W9m��p�l��5y�ܚ%���e�s �*�U�Gx�Cp��������7k�Q�Uڜc>�Lv�j����~9��k�X	o��w���(4[a��r�N���2����A�wM�^�S~���lr§��7�����6���f�琟gGg��n<'��;�i��k�,Z:/7���}V�� �a�U��j��=�1+ƽ��7�vrZG{��[�>5�;���48w�����K��wO����q�TzJ�y��ɊQ�N�dm=�qD�a��=HU]Hj)j�#k8P�P���Of7��/�Tu�-�~�ϻUX����fUՊ���Bg �g�v��3Nn�����^����Yt�)�`�v^cm�l�̬��$��|4+/.��$R�g^�8�g"��-�a�8l�&`-wL�	|.u�6�Yxx����7��t0P��E �5@�Ds>s��g������3ݕ9�o��THK=8ɓ ��05��z}���e�v_�R<<Z�{�RmE7x[&-��m/�������Kx��
�B��	�d��C�ϟ��E�R��5v�x/zႉǆirÅ��Vc  `�H�$Ag�шx����Am�i�ώ]��)�j��i���W�&񺁼�N�x���^����1�ye/��4!�Z��>[^�%���۝]��N���9�l��b��t8�k��o��������;�5��b�4C��!��h�V<3�z��D���T�]��6�` ���e�9|]Ƌs�&�O��[ȇ��]v~�_�#a!���D���4��X`�	ĵC�y�q}��=M�z�+0%f�P~�h4�-w#�J�k}��`�8��H���̞��L6}/���9�Mj�U��K�&Ů��m�"W�l%v�T]��7����ɭtg8w�����4VG��>���sVX2Ǟ������>�a�����q��p��aT,A ���9����l��{�9]u�^#���;�]�����w1?R���w�I2�����pѫ�i;�k,��27tu��U!��o8Y<�Nh��D��()��+���:ܼR9���#ô�ڝ��]�����Ŝ�'�]+�F�x��+o;�d�L��ۑU������ >T1A�1�5U]DQ�>y�^s�:��kj���QG���WI���>3�/{�����y4��>�mV��a�6@��Q��������q�'�+}"B�i���MQ������c�[��W�ݫ���&a�����Oq񌀶L1��ü��p-�灺�;��Y'w�o�]��g�3�sǠ:��9Q���OpV��9x57 ��-��[��"���_�i�[�^�H3:C��|֎�qz�N�o��Ƀ�AB�Ɯ�K�[H�ޚ�ǃ�sY��������^d�Jj[$N`�g 3ni�\{�p|�q�xY�h7˕���������+R�0�[���:�gy�-��� ݸM�=��^�{�?��P$��15oOk���>T���<��|ڃdcfkO��q� ��Y�~�a�{����R�2���D_���;b�5^���r�k�j̟^/,��׼�M�FV����g�c$`��s���0�Zբ�h�5��P~}~�*	��s�7�E��lܹ�����Ã�?}�>9��I��w�=Cn/)�^0F$T=�n研
��.�h�l�9|��(	*lͨ2s��m8�[��IB�u�Ș/����{;�p��̥�����),ԋ<n!F���H��&D�j�FS���͝/qn��{�^��˅�1e�Ǳp�����ۗ�N��	�<-�����]Qke� ��EB&���[f̨
�JE@Ȁ��6Tq%KɆ�T]�@>B�Dt1  �P�ht `�A��o��Y��ɾ����������ky�������}�&�c���$�h���z�{��pjC����'j��{��6�LgBS����sk��y��^���#� ?~PU;;B�h��৾��fq�;"xŻ�q�-����IG���2q��JռX����3H��>S��Ƽ?���LE�kJt��W�zq��:d\�g3��M~�n����\�sx��g�w���s荚�����v��1G�Yؕ�A&c�B�޻뼓���C�U)0|7�r��?l��X}1���� K�%�$9�W*�=�Q����D�{9!��mz�ۀ<�7�g�S���wB����xe����t�(h���w�a�o�Vۜ��@(=
������y�|}��1 ��>3�o\���[�K�n}pu�z�XFć|e���(��o�+7KG  Խ�[�!>{��P��37�MF��z�ľx�v����L��K����ܡLN��v���Cyi|юS��$������a����X�M�7�%�S=��8��1�Wl>��ܮ���8L;��<���v�3!��0�X��F<�ߪpН�\�-l�hKu��L&w��K9v���M)建32��n]X�۲ӈ͕�z"Uz{�+-&(_�HC �r�j�A<�ry�)�{��v��v��0��RB�H�����b(�O�Jŏn#�e���)��z��n��{��0�BT,��V@t�~xORA�pv~��X��nj	�0���e3�wiO�t�{��g�vlbS`:]M����ݞ�f�����K��]�?3^#��k�?����0z���"��2n�3_^�Nѥ�w �F�36���Ne.Q���!���y���-p�0�g.g������K7�n�o�ރ�G/���=X=T;E9N%8M�}��3�^Xj��W���k��Lv$�h-�s���J��?:/�^��5=��HOp��n���#�/��yj�wx�=��q��u�w��Uqr��5��c'�#��l��PR���/������<�~��vr��b�0;� z]����7���gn&��h� �7[��]ㆨ|���CO	�w�.���&�{����T����\�H]V�e��om�
4~�HiO2���+��C�\믾����Z�L!�u��3
/���Ѿ`z��+�sz�Fr��z��FÁ-l��>��e,:����sdh�gnL;	^�8�d�Ľ��<��v9����>��M��z�js�������,��R�r�/��%�����h[����"e��E�}|������.���%ԃ�F;�*j�wt�t�L�A�s��p�=}N��{U�s�whN�T�vU��㾂��o��^%��*�_nN�SY��ST" M�v�5ل�\�l�;zq�4w	ax�GH2mȑc�0U�ö�ԍ��t�!9{����w�ܧ�q��*�1ϠnZ�yn�q��9υ��[� =��
�u�.ӕ��8��J�t,Y����y�e<�[���o"�[�d����-yi��8��Ō�2��nAt���=YVk\���ue�3!�
������IC{'��G+��c"�R;er��Z���MF�L��;a��Zw.<+�m�Nٻg楯����q����9-9��5���eн�ɸw(�$*0b�\�c�Yt���ξ#xsy9���֯��K��"$�2��D��HðM차�����|vמR�~�ɚ4�]�+�E#�#�;4C���(ǝ��f��n��}��H����=��z���w�TE�ҡl+0�wn`Y��w�}u��ko�u.���z��¢U�nhs����, %k7wV1a�xl�4Ѵ�	�]�1�J�W��f�S������A}�ͫЉ$˨�ܖ,�/�C�7�:��}ִ�!Fe8-���qOyS 4�bsn�*˩���V��F�\W~K��^�P�=��]�)��6l`�{S���Yg �@W4#�hǩय�2�mBh�o���`o^�aE���F��wP(��̺���{ˋ{\��fv�!���� �tjX�-�
����Ӯ���w1��<tv�"�L*�����&��fJ�Wf�"��I>K�͗`����a^�n���cىǉI�t�۝]F�,��*�Ӑ(�7c��s;wx���*n� �R���QÅZ�5�)�qб���iÍ��b�NʶL�ޅ�B�;H��5�ޡot�]�|H�H�[�!Zkn��Vv��X���e( 8�Q������2���,��U| ��k��T�t�*ӘW}{]P���I��� 5GA5�+<�ߟ��{t���5u��Μw���� ���0�E�&��i].3���Vl�;�=�s�wdSk�> �����V��6l�YCD�*Eq�J�v�]��Fni��J�/��V��'{k7�=IHIY�I&c���FN��Wr�)�nI�����C�5�WWv�%�!44%[ʌe�"�PJ�,e�y�����dZ�[1�E��L��i�V)Xc��-�&3:��2l�c�>5�{{pq��N�<�3A&��q�keqY
��"�h�-�T�˩5��1"�>�K2l����Ƶ�oo�:t��y$HI!-���~�CU�eʣ/V�5
��11�F5=f����d������Zֽ��<t���'�h��,F��v�X�z0�e�+P���QE�s&NN�Sgo�kZ��x��N�y"�w�Q:H�ad�(�{x����`��		u���������oֵ�������<�"��J��iJ��Ⱦ�ێl�Z�+*���ُN��;x��ֵ����:c��}���H��.fKt�%c
�h��W*�֩]�2��E��X�82�e�$k�X-�PRw)1PP1�9J�m���Ŵ7)XTPQFԻ�D)��� $	�#�1�V�����v��+������������2V4�+nq�u�4����FA��k{�˘{��믲�b+����|��� j
k_�s�t�|3��#�>�"`b�w� �����sy6�2���7��]o�ף�';��)�I����ثva��3O�s	/��6�hP����9��7���ssF�IEk�\�1���nj����9���L�V��$�k��il+�_>;�v���vlu<E����fܶ�ǧ�4� k����:����}�ߕ	����i������a�oi&N��bC
-�õ��`W����1�T/<��)z���Ѭ'��,�̎��?vm�l</����ni��L{��jqC\N��;�.myeS�s�`��y�G��c�@ն�������_��q�|!���2���}!N><9�>�`HQ�p�p���EB���;�qg.��t�~b��6|��
�q��>b�Es���O|���$_©2���Q>�@��/C����{߇җ>ߜ*�s��Q&pZ����@�9�L#z�������/�p���l����[թf��t8�;)�<��H��sO1Fr|~6i���ƹ�-�&��~fn���4���5D5���<�q��(�z�-�.��l�������b����:BѦod����X��n�#��uț������;<���hu���:\rk��~fuu�����;�2"��`����`:�����
&�H
$��<���|>G�󳮧G6�����}����l��������VJz-�Ap���51��Nސ>@+ږ�K�-�͇�H3�ZEt4��r9�J@���.��2��1^���=y�1��{�e�e��~_^w����R��Dax�m�Z��+�W��k��/�>�����)�wec
�O6�L�3�WSqq��-5��;��f��N�w�u�����l%��˸��<"��yn4ݻy";�{��t��b1Mr�{���׷��Z>i��s@��_��/����YDM�{�ZIݺSOl�`O��[�2��r�D7������"���Q�n}lT�SyD޷F�Ԇm�{P�����'���'\^����z`�}w��d*���'��x�����X�۰�y�3����%������s�[9A���L��k�Cj�3��a��ud��V�c�%�5K�,��������Ǿ|M�	m��s4b�鯬T�=��
k�%��a�z���?Y�>�Y;�S7ϧ�X���V*�v��{����r\4U��H\����'�~�6��x_���S7{�R���۴��u?f�Z���\�Y(8nJ.����T]�D�ߍx��o��l�f����� �m�P�ѿ��Z��=�\N�F��@BȪ�t�݄.|�[�|������H%����n	�u`�J�a��1�8AH�	�'$l8���.4\���f�T���������#$��Az�����H:b��R� !��
>_'����}�{0O���X�F#h"s���H�5���)���d;Շ��Ϡ�����W�
{�X����ZY.t���|�R`��%�(��>},�4����Cӟ7{ƈ垁���-W�-��$lZg�}|b���M�"�spq�a/��=U�%��򋾣Ƥ��MW-�R_��Y�����s;c�<@g������$x��Ώ�{r���cS����ir�?1�R)-�·"�\Q�nm��P��W��,b[m��" ��[e$��2��:���[a����v뿸b�ռ&�$� h{��䴅�U��GA��H�0t���Y�����,lc�R�vW(�/zO�&~�h�5D��3!ֆY��0 ���NF����*�O/���wv�n,�V�Np�7;�{k���|�	}5+���D��g�At��E��w{w��{�Yq>�s��1IA��>�*�{km�f��d�0R��ډ�z�E���V�'�L�m���(@;�+/:/�E�[��	-C\y/<��k�U�fn�Pw�x�r�F�-�q�|:�pgk~u7�b��c���)خ����巓z��:�rL�FX9���L����Y���::��<�f�#�ou�\�<���^�)r�i.�C����ХG[v�wYܣ%�h�j�E�}dHr��s�y�D�@��C�Pt0D ��A4:Т˚��Z~\�p��q�8_Y��[4�f1�`ف����S��u�a���1�&_V�קg6t�D��"SS���2��:�/t[��xJ�n�/�X�Ǜc��Z���!�5Z�J�ni���!�ܷ��l+������`���vP0��^��ǣA��/W������qy�ʋ����Ǆ�
��Y0�����o��c����v��O𔀁�0�n�F���=��#H�v�:�>���1�»RT�ѳѸ��mA7������|�j��<��=�&�Nl	������U�	���:Maz�����Ŭ��WA$���s3�@o׳�t�F�����3�r��)��˽�xǡP�Υ}����O
ɦ�\��4�!����-���Ag��"B|��#�l�M��x,.��y��,�̟��KϞ�C��|�w�a��u��>(��G��P�f��<��n��3����㴻�������"U� L[JR��|ւ�3�������_+[m�c�)��R�+���Ě)\�ߺ�lmpԺ� ����vg����.O��JY��2�W��pI�P��u�hw��`*e��s�}V��ΫRk�M��9^%>�K���}U]$�b� ���FQ`��Q���s|�~|�N�4o��ߟ���#i�ĵg:�xr�߻��Е� �����瓛�����G!�y=n���Z�[vyFW�Z�At�8��P�}k���P���C�ၭ��ݯgOO�a�,6�[�N�����C{|�G�l����P��K�t�i��q���۱|���#r��P��x�?]���kn]F����-���Z��5��屠��O�._��Wc�?42��*G�G]PĢ� �κ0�١�a���>��������K��ᴉ��VCJ�� ����`S��R<e��/b���=Au7pY�t�P�`�ϽZ�?w]����&26<C����=_��z��M0��A�=IEf�S��0{�r{b؜��{%��d�o�Lg�W8/��h�lTy��R�1$a�8�u��4W5�e8^[�1;3;�w�����֣֩އe*�vp_F��W�cy�Ц��bY\ΝW���M���0��A�R�����1��fpt��(�n���}Ճw�o�G�] ���w�-���g�0��{U��:lH�:O��j�Um�6�u�9}LpJ;�4�����:n��h*�\�/�L'e��k^�e��Kaw�:�)��G�R�Vr��.����fmut�}c|s�;��kjWutt������p��k,���X�F��g���Tվg�O��`�
�`�E`�S@1P���9�v�~U��Ǐ�*XD��^ W�2�`�l���P���PW`�|{Zd��Ӣ#��ޖ��)����]1�7@K_��c=G����a���|��B�jV����!�J�����C�-���G�c����K��Vv�k*����<g	q�0��ݰ��۱�7����xjo��+�#�����7z<loIw
ۤGI f����`�Go��zV���%�)�n�9c\Ok���M�)�hp��w�c�;~0o�����g)W�.��+OuˎW|����;��àgL�ֈv|K�y�ݘ���U7� �+«�)��Bj�����8VE=<�������VO�����μ������wN��P��
v��ז�,?-�M�͸��9�v5�$>����u�ÚY�<ER��.�D��/\
���L+�6�k�4\\C�=so{�^�v5��N7wEC�O?��b"�q��<��@��3��������:$1���(�Ν~��|�*<6{�[�j�+��X����2p΢uqt�����~�~�1X�s�/Y�T��K%�/u�c�Cs] ��fV��8,��(�i&\Y��Ud6��;��`"
���n�n²��;��!U�Zʍ�n�h���xp���K��*��PT�7|�фM��5�^�{�s�!�˅�c��A+��
IP����)JB0˥@�XQ�㶔����889�p1E�	 41SPXGCH1��DG��<4kɯy߼��̘�X�Hd�ǆ�L������>ߦ�z6�Bp.O�	���]��m�E���y�]�X1jR��1}J�g����۪!�\/����p$R�����;�K��ў�ۈ���� �����k���A����y%&���PAp*^y������%�>*�X[�Ҿ���ea�b�q��P{�V2�s��!����G@�.�t@��ʹ��y� ��s1}��8�x��r/`Y�S��Y�e��P��ܣ�bl0����p8� ��5ٶ<�-y��-��@��/�P޼�e�\<���a�J6�!�<��	��+��Y�H30�y�bPhGI9�,\����Ʌ�>��t&�^ׅ%ލs�r���"׊��>�;��P����J@��xT���&r���á!m���B~nˠ��`�l�� b�z��q�ķ�¦ v���r�0��q�]�}���	���,��%ϝc�����6���8P ���G~縩�����S����2g�L�L@dq*}��Q���^���I������G[���3_1>�(�%�J�q���T�4��^��7>>�g4a�C��W�!�U�s��5kd�w8��[I����B�^�E�5d��Ы2�E�[��]B
B�>�
�+ޝ���K{�6�jơ�KՆ8 U�ݶ�����j��&�3u���;]+�]Z�L��wI/���|".�6"���(� �bj(�g{���ϛ�_�w釈�5SJ�C�A\����p���Ŋ\�3)i�+�x��0.�ߊ���gz�޽I�5��\fE� ���<�^Z��@�!�����2����r�fQ�jV��]ٗ�)2y��l�eeou�K<�ߪ\�7�p��XBV�[`������=��sM>B�����Φb���x�ڽ�8��,��e֮��
����qz���N�����[y����c/���<Ų����&�1�9���s�9m��5L@h�k�{&��۩�6�Q��$]}��~kO}Y��e��kxCIq�B����&��߬����bk������yGvRH���E��;�@��3I��XJ�y���ڬR|�|�]�7�XKSx"e[nѦ������~L�=�:�;!��{��>���'����8)�u��[��������vs2h�������"ژrJq�Izq���.uw���	ƧIg�@�_��u��k�f]�A'��{xwH�z4�fwO`�5�ZG��{�9�^��:'��J��`�h��׋�
m\j)�lRvv����+&/�p/��=��uҔ5�}�K�]��>\
�,}��+RO�n�|�%���TF�2�e;��j8�m)|��#3F�շ/.��7w�~� �8 �����hb	��"!��� i"H({o;�1Hp�~=8�XN�v�F=���6��5����@g��N
~��dޟ4;����+�W�`��i��>�;���/�r:l�+}\s��h���[�^�~⟳��Z��K�s�8B�ԀmP��5`���W�ȅ�塵�ZQc堟}h�K-�ʴ_���߀D�d��0���ü;���y6 \T�*0��D�L��X�,��bMSn� �Ǯ��,9��S%?�(�5Y��}Y�O�V�q������q���0��\���:3����tڕ{3w��8.�1�r�9���:�e{Xu��F8�x��s����`����ށ�ׂ�e�����f'I���;���~lgw}�~N��>=W"y�Q����C׬�zaq=��2�̾�HWx,��֍`��[/� �ށ��m|1��׽6ܝ`����ʅ]Tx��n��gZ�c���<����2�D��n�? E�3��a�`_|�#9s:�	W�������5�D~���Q��qMa��xO ZR����vEk�`K�6C��y�=q��Q~O���Qϟܢb�~� Y��?'2i7o{w�� wΦ^��r�.GMm��;I��E����i�"D��Scyț��טּ�X�ٔ;e3��+�Ŝ���֝-�6"1��6�Z����Nj���\+���)?��#R0�@�!���"'|��y��|���X?r���[C�,B{��Mj�L4B��(�����^��U�biy�WY٣����qC:='�}�˲�W�1�u���=��斀�%�.��R����h:������&IlC��?r�Ԩ���僶ܬir�:�W��V,�I��x;0i	�!k����{����o�3�[�:W���gH|^�����4�*2����F�75܆`���ی
�s���;2���$a����ы�AV�"[n�j㩈��f]R�׎����O���Y����#�B����3c��>s��������Ւ|���"_g+�vJ!?��Mu@�=��X�<�Xo���d�=8))�6��g�	�k��OM�-�;�zx�[�q��9	�e�x��}K���;�÷H�^��kC6}H����iw�%���u����M�9|�iBH�}��s+`��ޞ����c.Rn�6進VW�|��WR͖�y)�Iu��]���(��_���W���/����*~��0�n�wn���I��:´�zk���H��'!w��{b�v<�Q�kU}�0)�9����P5����Ωv�1m�h��+!є�ը�o��o⣢���pLˡ�,���M�4]f���*�S���*��WyV�$0_J��@��T��ɗd�A�Z#tHgc-+ۋ�{6�䡊�1)]u�Ow[_.܉`�q=�ckL2�Z�LI6wm�I�f��TTB��m��·��'���nlji�`��	eY���ׁ;��v�at�������Wv�4lj�T�a� ��A������Q��pS�*��T֧��%�fr�RZs�|��oz��Z��;��;Kh�F�c;���Vq+����e`Zd�g;����̵��K��\��Ji�5;��E�u��%L'��MJ�Y�)ᘉu.�h;�R�n�ˁZ���3r�Z&k:�m�u&����p9-��ۦ�*�ry�ޜA\dd#�0��cx/tRr��ur�)-�ݫ*B�+P��E��Nor����tr���ʦlh����-˼�rNU��.��=���Mи*ݦHZgJ�5�VM��4����+z�s���`���e"e5ĭ�]�ð$���Jَ�fT,�`ݡ�ڔ��p
i�E��ڼ�\lm���J&4�UWݵ�/�����h32Aԗ�#�*���Z�lIj��\�2^�G��#��T�#Ćbo�v�݈��"B�
՜���}�Z�l>��k�/��t�bp�ɒ�ǲ~�eя �
N�\ =���c.�2)�M���#��3Sc֐ſaV����Q�a����tt�#KN"�`X9gwp�z��"��1^+BL��=�vĬ�U�ؚU�z���ļ��=�z�*ł{ib�ԝ�6��1�v�)�VU��ej�t�n�gq�f�uP;�RSZƝE>�:�e9�N	�d�h����[�*�n���|S�(L]]�Nf��qvbț�z���y�'�+��)S3)i7oju8���ș���Gd��*v�����,rC6�Kڌ־!ԗ�KmP�o�`p�rFq�Wwj�/i�h�K������)n�t%)��Of�v%˧�\6�"	ZP5٭�Vn�D�\�+q��(򞺶{��`&>[�M�yD3ټ_[j��Vl>��j�6���Eu�:u[wN�ܩSa��PY���z���v`X��N���{��S�ڹb�m5�:�͜���{e
�7
BD�f¯�Grqշ�"]p����iHJ�N�,s��D���]	��g+�޻��ħ�>#	9n{7��f��֍|�;�p]&&��<��"���8�ĠTYt�P��3P�I���Ʊ$��(�.9MW )��
J2��)�K���K�&�i.��b�ŗM 4q�˙���Lq�[q�v����Py2��
	 �N���,��Q8����F!��6��()ƙ�Uʠ��x��(3��NB�'�5Pb�e�.�-$)�5�R�A�����'S�Ҥ��g�_y��ZQ��QŠ�eN2���m(��y5�����ֽ�xǎ��������+V���Z1T�U�QC�=ѽ�f�@�8������ǷƵ�o����d��a	2�Y:z���#�{ )DEZ��5	DI>;zv������k��}>��X�O����
�{C8�b�Qk*�t��E��f5��m���ݻ{||{{|kZ׃ǌx�r�(�C�b,1��;����XB��^���{�&�u��ƽ=5������Z־�1�<�CGZ5�:�*��_w2��Nڋ�oZ`ui�Pr�卫��»[�UZ��N:zzv������Zָ8�,��|���)[r�-�9b�1��\Ab�Z�c�4繝U[*�*��X�.2�D+W���uZ	���)[�w�TD��ik�E�9��+�e�J�%h��hr�LL1R��TD�Q`���JR���;^�)�̅f%����L֍3[iE [A�J��Pm�,Z�U�*��۲�8��U=Ʉ��Yq����/D=�H�I��ĕ	W�K�2c��ih)�OP9#�#H@B��Zm��P��7[u���r�͢�Ts,�o�!>Dɡ��CC �`�H0�0�k��b'v�Eq�	Q�v�@���G��t}W�.��^	;������Cjsf�6�u�k'�R�,�|��D�����l+K�}��
��s����D�y�n���O�܂qYL�4���m��h��n�Z�z��{����@�樂���K�8���Ӑ.�8{Njjm��b.Y��;y�����s���.�ÿ!~��,?O0��s��_i��b�����"]��#9�R�ouY��5wW��i}'��*3�^��^u�"@��7u�|K�ȟ	�I֞N�{��eT.e�Ž�D�_G�kU�\��a�cɇ�a�eݪ�E��L�w���=3��2strz����8h��U4�3���C�7 Lx������B�Q��KhgC�;2}!ۘ1�׻��+�~�O���پ{��{6��ݘ�5�p-�_���\�C��;yR%`����0�~���	 t�>: oQ7�u},��0���Qe�������U�hh ����M����}�	�o��G7��������t��|��W�>)�VBO��r�nc{N�qd��ut!M�qݫ��b�pm�P�L���L�Tخ�m.�_��_���`��ÿ.9�:�$Yۨv��>�����ޓD�C���LQ����Vg!ڕE�]����^�г�ݝw}�#��B@���`�`$��h`0b���o޽���>|:K�O����@���c;cX�2��Y,2i�����~�^s��L������^��k��������=^�'��4�Mހ�i�t�����Pg9>{���O>������E�j;��n4y��O���>��x�z��`��/J��"5����]R�yC�S���x��|h}�B.E'���M�>���a@��u��k��vyK�Gk_om
����ż^���;��a���}���xǵ�q��<�O��a���]�)���]4c�dy.�Vp}֋�[G���+|Ł��_�{�r�=~���/���ѵ	�Xa	ԋ_��/sl
t�������G�-+*|��:���z������l0�{s:���'����w+��jB�Cd:�iq��F60��Es��r����y��L�i.�9!A�4��g�`e���%ҷw����U��<zk��k۞/v2=��ϭ���r.����FK�f�A|�?��4�5�"Ox}�|�՞�lc��3�w��'�m��qV����=-8�L;�]E��L�y��tS)6���*�K�%�쑘�i'y�}uҭH��� c�S��q���q7M,!DQd���U�l�J�Lo��B�*��\;���.KmSU��J@t�]�ə��N�I3S�3�׾��)}@>�#,�����!� sw����|�������W����x�3�_pж�y�[�7�S�_({���;+cu�4'��MA���qi�����ZA�zO�����]�eo���|��Jb�/q���A�ad�ڶ��s\6�^�a'��4"�h�. E�~T|pyB�1�}N�/�1�^$f�����J��s�Ԏ�{F=�,�Ɨ��O�b�O����۝G�'M�sb`�}�|������!���d����`"�MG|'Ͱ=^��#�M��\�P�4����(w�rx��^�Jú�g<�6)c��
w�^x͛9�o��r'�[��\��$�WP�^�1�k��(SsN�,�w��'��{nP���b0�# ��~~�_"���;)M�M- �=�>���]A��|�s����X7�r�kԹ���%^����L�͚���՜����f��7W�6����_j	��mx�t������9EY�p�H/~\��p������癳�88�����bX�v ]{��:TH�����'U�r��.�V���ۆ��v���p�o���ƾh�y�8S�'ߣUە�բ�eg!16�#�wPh��B٫�=�gs8C�v��k�\��x��MV�K�G�Ư^}[�,��}�����B�Ew�O/���b�7�9�q�H�H�H�䔌���TX;{��B��R�$��'>l`�zbۚ}�/c�a^���b��$H�r[����|n�.�����3G��D�r�n45�O��q�&5=�����>�;���(�"��z���~qAG+(U��9�2���o�:��:P�VՖ>D�A��V��`=��y�']1-�|��<����I��<��?o~�~?G�x"H�m����d*�n6,�|6W���`���k�kN��+sP�S�8u��_��x)��D�|�5�_��ߗ��3m�#������0���U���x�fˌz?6��hJ=dt�,f1�`�g^ڢ���T�Wb�z-�fz���1����5�>�|�*����˯y0h����/�x�yz����A�t�h&h���A`l35ߤ�*ɣ�UD�%��mO���(�{�ļ�6�Nڠ�C�����!]���vǇ�#�]�yv#K�gr��@��]�P,=G�G0�u�pmM�~N4����K�S<{�^h~U�K}�o����>S��U^����Exf@a廳���V�ek`�90�s���3(n�$N�2��LGL�R��e��v\]��n��q8�*�!jk
/[���U� ڳM2ض� h=�ԩp�7M? M�봑+Q�e^N}��h�5S��F�}:�we��j�q��nI� �n��p�sk�q���ܷwq�������$d ��$j ��F~T�؞���"⅒E�thp��
 x���?zo�����Ԗ,H��s��R�8�}���������p���g�юZ[��{L�y�\]�����Ķ�[�{N6��Ovn����mx���Ǯ���.�n�J�<��ǒ��ۼ�.'}
dd��k�Oߡ��O��d!
����p7��F��'=>g�'�wV����y����3�uՉ"+y�Z��&���K�Ȑ��Μ�V�x^l�!W~��+���y�k��4O�\8�0�azcāY���H.���l|C��X���ϽO{�S���3��\j|�xŰ�p)�}�i��ɶ�g䁬)��s�+�n�(_C�b��5d�o3>�델�d>o9�BHa�P|LO���C����t�wJ�ֹQDw�T.�6=K+�?��6��M������P�Ģ�����Z��Wf��xP��<��>�{,�t��]�mmA/=j ���� m-��1R3mtq A'�*(̴L�{���^���܌y��v��_��9�fڃ��݌5�̯Hlh���6����:4a��2Y��s�� ޕ�}��vn�yWg@hZ����r��b�u�b�dj˿�T>B�����
nu�$�(h<Ṫ�g7V"�����L��7�O#��u#�ַ,�z;]`��PF���x���b`�`0b�����|pf��x0�4#��,�c?.�e�>`W�ͺ�cH�SMC{de�'Y��s�m�V�B��x��1jY&���\0y����W<~�3��W��Z\���YS�)�4��o=�}(O���T�3�&(����q���5�!~�|�r���FD>|m�I*E�;��:j��H�@��=#�[�/�צ���N ��ɡ�&�\�g������sy�8=�vdf��o�mL��2�(,�;y6�Ȩxl`�kE�l؄��r�|!d�����3ӓMrSӟX UM���p��X��y�:}u��Eo5F3<?�i���|;y��D ӗ�/�&&�_�:����O��X���N�3fh�,���,Д��̦b��ã��"�b���-ńo~/�9X��2��U��|��rL򃵝0���J���M1)�[���0��ռ+TJ����	=<B�th�rel1\�^�h��'��i�{�kՀ�Ψ�qC̺*��F45[�v�y��ĭ{�j�wKJO���/-�ߵdsY�>���W>T�ᜍ�vv��X9�k"Ф�X5R�
�97����/�̍1߲��^&ض�vOB�(��(:�9Y[�vSH�&�ǻ��K�\3/w�G)v:J5�&)�Ʈ,��Y�rtu����0bP�� ��8�y� ���=�����ML>��̔+|��G����em�=S��3�����7����^���o4��p���6V� v��E�wAm���/<�2�T9�{�]U�_,(��`�����;��4S	��6��6�9�(�@��FaVc�� ot�"��u������oF�z+_��|�H�I���^9��y�]��/�͇�qB諪�Ҕ����wg!b�`� @�4��g�\��Õ�Ԃ8�
5d?��w���Á_ޡ9c.�E4s���r2����a��-���R�{��OzP�myP�z@՚=N�t�c	�T��x�u�q�s�zs��E�Gl�HΎK�72-�Խ�N�y(�L���)0g3�o� W�W]���W�t7	��u�kY�����R6���R����	��W��	>/eٶ�����N���7.��y��>�(Ag�͜�^��1q]�):A��8���{�gy�+�q�[	�Xw<��yTH�`��������ߖX\UMK�B|����u���?Vٮ5�'^Q�Ӎ_X�yˁ����Rޭ��'�y^�ֻ;^�ɗg��l2.��qp�I����Dh^5�.Ƀ�HFg��L��:��<�rG���s����VC���D�d3Nrz�0%�[��I�{cgs�9��`�����q��ZF�H�D�t1uBC�^��s��:>jNy��׾׺�ׯ�ф�S<�\U��_��.�bj�O�(v�*�����7����{۹�d.v��RS�-�cX���2���^�`��7)�B-�v`���X�q�IW���V�Z�v�6~��O���~�/�g;��A=Y��,׻�5�G��߃>s����.�E���	��݇W�ӯI��l�	i���r�TJȀف.��Fv�0kvmX��7�3�gt�5ŝ�2
�����N$�U�d�숯4��I����r]��V��0
����TC˺��X����z���!۱"{����,&ٸ57��/E�A���-���p"�q!�.5f�P�*5@��koDo6°�ᔾ!���*��xϱz�����s#�v��3'�s����{U
<�>��<���+��"G~;�06<C�wʭ�����v��X�nnp,K�vz���;�u�\����~�	G�E�C�ʳ��D�g-�d{�qGx�g���=�jD�tiq̹��c���>X�ծͻ���~��o{�����~��,�Zx��&]non�	�I��d��̼�\����[����t�C.Z����:Vg���)J�%F�Ϯ�Y��4����EiK�	��m�β+:�h�rVNŚ��T���,93.M�Ы��fo6�EoR-J�����x˅A'2��R�݊�;�qr�jeMt�m�nf:����?F�&$�����8x�<�y'6����}�)�:�h���O	�?(��R>��-�/.��.u������a
�*���H�ż�|Ѫ��f���<A�����P���!^�2Y��?�� �4���:B�Gu))A��UM�������z��`���7�b�1Ѭ<^�'�d_-��ڿ����zj!��c�uY�KO��h�q~�[���
��o���˓fj��.�8���p�vZ��&X�$,P�Þo��Ȯ|�p�>�o���=�Tx��/�#T��?�;\�h����z�^]��%�T��|��w/�.|Eyi�.�����[*"0�{�8rw4��(߫>�}�����*�\�3���5�;�>��Y�+�D$�5TD;Z�8�j�qJ������+���f����w�W��_'�V3�����//zY篥_��nଅc�w~�_t{�D��0\N�&����I����u����w�o��W_7��;�S���޺�[M�N���5�Ǝ��5��q���ea|�!�e��X�\3#��	'�A�lm<���f]x����KP329S�=��V������L�T�p��R���Y��,��{�T�n��s-�;x��H�l�a����%dM��j`G�}��Z#�Х=3-P`:���`|�]`˱@gy��{���y���L��0;<�a�a����En�r��]�Þu���:�[�������d�y?���O�93Sgv:1�m�38�R�8Sw?�E+�t�9�N�^��W=ҭ��8v�`Q��X����[t�����Q\�7�zY�����-�*�E����.Ou�-.wi���0s�>��7�j�H���{��N/����{��Ҏ���ʾ`i60Q� �Ɨʇ0�:Ωkͪ�"ೡi�5���+m��Ѻ�/<�Kߘk��_���-�u�έ]]�o�������_���D��0��Y�I��PiOY��稘�V�^�q�+ni��W����XzP>��w�|�Ķ;�];��yA�WQ ��6���!X���@�#�z�;.oO@T&��FX�����]#%�-����rs�����v�N�d�?0�a�����=U�}���k�?D;�M�}���\>�אU�0CC�繨�yiia�z&�d��/��5�����.�Z���5�������^+����?_G=�v���>��!%�9���ۮ�S��x�jӂ��L�u�]�h��C-.X�Zt��W�6��pT�2���N\��n)K�������H��K8p �!�VE�Y3�*W���K1e����(����o�����S)gt�sfPo��a.6"H%d��78%��r��󦫎E��ҭ����0�7��V��H��E�|�rws5�t�cg:}�ic�v�Dk�hO�+}�j���oN�wsv�K����A��Sc�b�b{��WdL�On˻N�1��q�ùw�p�;�S�5�,@�+mrNW��Sě��1:陶B7��^Q��q�˅l�;)�d��:�:>�Xs�;�Zn'�z�j�,�8!�r'�1ZW����}�bvMZ� }nr2�;�S͂ұ$������ѝ[M�ʇ�ĺ���7���25`��k�;*�!3�cTѕ��`��!��9�m��lM�M\׹\�ov��.�d����ѡn6��ӂ�%S6!s�E}�c��]��^�R��N{/��i��Y�V���K�4�]�U�l�s�_<L؏�$j*vȸ)a����-<�����1*�s��K����8	������U5��9GÔ�ږ�s�&'��pFU�b�t%�t1��"�.<���������-�y.�u�ML��Ү�G�#X4,5`�m��g*6�z{���A��S�%�Ʈyɖ>3�Q�(��Xx=�v�a��6��;h�H�DTL����ؖ�wm�w�5�*��5$��%Z :��2@/냪q��]�4�fekЃ��Qt�؅6�@S�@4^{�7������6�Or]��#*=&�Q��Z��*Ԉ3blp�keg:1��x�����K8�E]���c�ެ��4�Ut�y�>�����J��3p�f	�Lɞַ&Q��O��jnd8oG�x�ۍMN<9c�t�����Ϻ�;}\[)WF�\f�x��a\gi�ȳ����+qӎ�.2�OȸKꅹ���[d7����u��TZ�d]_��l��n��|YQ���n����R�)����2���7J۝Q���B�'�[*	kt5s<���6\�OgV��\E�b]|�.-��T�g$p+���Eg1�����6bw���$;!�Q�4L����y�*	�I���u{�\Rb"�A=݂��1�;�0��[��$���[�����u���w��o{ *��+
��+ᯛ�|m!��.Z/uM���u�:Y[Wb�=\ؓ�b��&q�д�G:8�5K�r���)�kv�]K���]!B�*K����%����t�tc��Ur���}ãĎ�[}W��[##�*��-�&7쇬�TJ����n�	jTW�QpeR��*Q-*�����:���ƽ=;{|}{{{|kZ�8�x<��b�[-jV�c�--(�����v��F1>��2l�};����5�x<x�<y8r�ѩM�6�\b�[TL�G2��)TE����eLA�X��ۖ����ۧoom|{{{|kZ�x�x<��=q*.F�۸񢪢娹�<tU`�ʰCUK~�K2l��Ƿ��Ƶ��ǌc��2sZ�h�{�av��.�a��%S*����r��]siԙQ�ː�5/]|{zv�������k�ǌc�pim�*_m�1v�f3�ܭ�Q&[���Bc0Rr����]=5�������k�ǌcǜ9��eQU��,X�}���[zJr�`�H�-̔\�s3�1�{�x��ʱV*�iJ�j�B�-Z�e�����5�
�4EDm�V�R�uj���\�s���UX�ZN�D�"=[D^�j\�e�y�9,��!p��[\�!ƌT*Th�8�e�O���|��;;��x��D��l�ɤ��eoѭ4���<po�����Ĉ$�ɉ��_�~��O//�#x/��"���5o��J|�N��Q���M:)��-;��<�J��9լ�݈���Қ�W�Ma>��\k�8(������M܉疫�zt�ӹ-�����<�e��B�&,+a���Z��MRǤK��\g�V@���җN����v�NX��Bu���O�uf>cs�P�U�Ї4���c�|+]�Q��f�������Kt��@���z��Y<�a�.�/C��W���Rvfg�ʪ����p0FG�˲��j��ݭSõ�����6H7�Q�_`S_'��t�(}��j�Ui�Z�޺��=��N��Z��Ϲ�F������#㳽��y�-�^���{��k0�x8�n�$�HO�=�s=�e�;�>�v-���ڜ�Y���4P���������H�-B��[wd ��Xs>�Z�lz��q���@��O��
}kM����l9�7�a@��=�)��{e��8��1�w�ΐ	��Č�Q�Y�k����o
��~�YkA�[�{�LPY�g��X�`P(�!bKTM�W�y�Ϻ<��0:OSY+*W�"�;{��R���u^�j��Os����׶�̼X��}Vj.����i�:X������v�,���s��H�FQ���g��{�����������C{�7�0�0����Q��\w;�61�^0�������`2j�vk��m�὏��Ӌ��-�@���H���c����o��s��|}8G���+�<2�Q.�Z��`:~p6��Û��a^�Q*��5_��P�+�/������o��WA]�9�h'}��� �0��Ϸ����?/�(������\2|�dW�c��C�0��v�o�î�m�{�NR�*���3��|f�2���π��U�����,	<QW����|o��L��hb��x;Q}cwu�
�{H��y߄=��v7����6y�����:hy��1�C|�*T�z 5�&���&3�v����=0�qm�@L�~��8�v���������MA���n�n-����K8 �����2~��5.��.N�WX�JC�|����^-�K)�ʂ][�3��019�B2����C�7.�t��u�$G0��QlZ}q/a'��G�M*χ��V��J��#����p=���-��SK��i�k�?6Z�./��5�)���׻K���r�*�w�vC��tcD�ˊ�\O�Mo���Ϲ��~t���/�gƝ���5o�t�����P2[��vIɪ�k�*a�pP��A5�.�X*�]��7�� �t �W{ӵ=�;�\�:1�h���bv^����ۻۜ�pB���-պqdS�&s��]���8g?��	-�"V��Ԥd1��pz�Z{׻���y�^p�P�#����Oiw�n�>��t;Cκ��ꁫ/���f����vC�寒�P�4����m��MlS�z�2*a[��Ď��i��|w�"�F;��On��5\�m���� gD?�"oa'j�լ/���+^q����Z�^�.��c�����<���Z̓;s�|��w^�:DϪ�K��\�|�5zXS>X�x|mfmU�7��S��Y�a>�x@���*�95*��X�������z�[�t��v.Aׇn���ú�:�%�V|�"5���Q�_,6��ƴ�|�"� ᆇ�������d_f{(9�X�	auE�W(P�^ f��M�э����1�j&��.�4�g
e�P1=g��#�K��i�+�Rx��;��	yޯp�7���U��ߝF��'�gp�~��r6Q@�QI�Wϝ8>�V�{�� o��FH����l�{�ջ��5�V9\0�=��Z�5P;�=�R�u�S��"�Ox �ߏ��^Q�����j7}2��������sYY�^����Xfx�V��H�ޛ�+Fu����m�gr�\��)�h���cjA]��Cz5s�[�����3��Ke+��
���ΉOm_E^�d����;��d���1a�o0�q�G� ��Y��g��[�zp�5���4�� 3A^h> s�b���&\G^p};&�޵��7�k��2ܐ���v�ƨ�Y�u��B��RN$�l��;]{u��'�>����{�I�|�s4��n��m`��##@�9D��9�Eon��oF%kT�W}�Mb��	� S��
Wca���oAB�Ox�,%g�k�����_Wgi�V���nw6x�O�M>���t����;�*�,;8Q��v���fdz�{�ɯ�!}���H����xY3yt���`ᡄEc��>cX'�w��9�mkF�^O�c2R�K��2v4���;��j>��g�{�`(�c[����r���3���ZZ9;K��&���q�^hkƭ��S�@N�[�;���Q��s�6Ȣ���&mt>&��i�`|܆��N̑�<�T��_C��͋6�m;�"� o�R��þi�
�]�=ڪ&�6�v�`����W1A��;ٱU��C.1�1U����ST�Ħ�����kS��c4���6�Eү਽��Z���(]�j��'t�Vd��&ڛ��8��Ä�8�G|lqP�E�o=���g~�wo�0�#np������]�7:}�ʓ>K)cV��O�+U���������/�o
;�Ƕ@m��5�KO�R��P�e����u��Y<~l�pݸ1F�:�[�O��vT1k]�3Tf9X�߽Na=;rw��'����{K��`��xþ��,��vG�T�y��PVe�睂)Nxܫ�����T���S�W�oϚ��z�Z�ڵ$ڸ}6�K/u�hP���J�pܮ�{i��'�� l3�e�M��}���<�1����$�=�>�d��:��P3�����7�#�,�/rp��B�6󷻓�a�YӒ���?���O��v�cf����­0��:f��__ץҌ"+}ם�=�ǳB��Y̼�c��5�5	Kx�(QmB���(��b�ۢ��y���������p��Hm{�E���O����t�Y���]�_�����[5���\�/]P�v�ա F�z��x�x1��(��p� 28�|�V�sK��kGz!��2�>Ra�Ьr���Vqe�\I��oE��;�m� �&���W�1;s���B�	R4 0�CƑ�%#p�#�y�����9���rʛ]fШx4ÿ�l���S�}�c#�`M^]FF�i�3x

(�TNsη����}~�y�~�x�Hu�����g��>W�f�B�]С�?#�Y����u�ߥ�^j�m��&$ɩ�ݻz-Vn5���XTW����s�L�d)��Se��f�t�U�`�����:��hH������3�k�&A��8���iÞ��ւ�n�Z�v�6|�·�6�vh�g��v��mp	h��6^�ʒ��`�,f�Tȴ	^W�m���_/fu
3<s�#ׂN�0���\�+01�`��q}��K�V��
�Y�������Q�Vcc�R��l�u���A�k	u:�`3ǲCQd��Y{���k�L�X\T��Y��c��}�zY�a���.�E��\�X��oCu6���ic\ٚ�� �Y���@�e�G�o(�B�e�y�u�c�+Jf^z=���C�g{�vg"��ɔ��N�eB�4T'ڪ-0X�|;���� e;h��I]����Cx�]f�TJ8�����}�N�曻\&��{Rr4��5P�M�(�Q����i�
��i�a:��*vێ��	iIei�P���Y���O��y�B�I/+�����_�{��?��v��+�C�{�D�m"C�L�7�:h򜒼ƺ|�1�Լl;��O�O�RX�UK`���yF��n	=�ކX�v�d�ʾ�ί(��Im�S���Sߋ��.P�[��$捚)�y����)a�>�J�7��لڗfr�-M�/�ݴ4�H�a���1A��r�<�H0e���Ƹ�Á���Y��0� �yv�'�5����owj����I���ϱ��~�/qu�6�1��;�@��Q�Z�陚�z�'�JrƖlʍ�1���*c��#P�~�G{�����a��y�ۙ\�Ng]}kN�L���{�$�T}�{�&B:��&Q3D���%"#VЙ�����6O7����5��3@O�a��Q�1��p�D��k���lȹ�t�`����*�t�M�x���n���l�Y�oj�m�R�ƕ�K~�q�{<6]��M0��wX�(�Y���[]��nCԭK5�*f8T+r�wsFv�������:�qkw��onH�����&	V�+����[��7z�G��a������G�D�"k�l��v�5�y��,鱽�Q۾O��U@�o{�E.�H0қ�睼7�E��g����r���N���R���T8�=�n�[nõ��a9|5��wo@��v���Q�ٟ9��f.�ϝN_.�t��F�4H�b�P(�쪏<V�o0���X��-�Y>��Y��7{q�g3��k�z܏O�S�k�e՘^�3�"�� �Vq8س2އ�i�3=O}O~!�&�{���}^���^��_���4�s2�ۛ8l��y�D�K����_e*+/��L����O���UJ��̊��ok���F� ��dq�Q��WP����_"�C=r�SK�� fNi𙺴w-p�ɭ蜑�O�sAU��Y#z�䨆��v�Kv�)��T�+̆�S�nkV�����{_���^�Qؽ�j=�ɾ׿|��ľv�;�7V���wI=�n��7V.�/��h�
���r�|�*&*�w%�0ʀ�d����ϧl-����+rU�{���*�d�\��%��J���K����o�%�D�̻����;� ���f�z�y�ٞs�<k�s�|������T3�^׸��'>ݑx;� J �9VN��z{�2 j����������D�n�i�fS,��櫷i�e���h��l�0���P��^�z�~��Q���������il�����L�6�� ���c��y��LR��|��=X�[��U���7�~�R���������'+k�SRL�>�2lY��z^ WS�]�fz�s����'�*������ׅqa���އ04Z�Ѽ2�2.S�ۼ �������lZ[o���Hq�Fz�`��ӊC6ңft���]�nÇ���oDO84z��}v���S�#|��T�.UӼK�����7i���*{="&��/ܳ`wvsE']�w����/*�4[�L6R�.֍Y�� ����i���ON��ґ(Q���/�MQ���p�WY����#�`ƒ���s�Ft�}Z�G:s3�^t�dn�Z���IRC�Olf�v�9v9t��DNA�)d�Σ��J:��m=�ӗ i�
uӷ��җ�<ԙ�d��a5�9�{��|<��*�]�ă�z�,r����|]�����4�}����	�>��+_"VݨK}i7�˺�/�P`ݷ������i��w����<tk^�<�~�iI`.��0%�p�Q����T��SyE_��^������m=T��iF��a�׻�T�����W�l]�;qϧ��;���w�W�w7^���|�����HtHU~�v�;7�nM���[�o��~���N��\�^3Lk��^��7W��uqh.�:�g�<���w����h<�OղagI�-��X�����J'h�����Ʃ�Zp��`vaq(��<���5D�W�cq	O���mC?ej����N��`y�\t�U������G^�O�Ms��R2��50�����w�4R�d�ң�9�%��lK=ޟ6Ȍ�n�0�����{�/�0��CG�
�����{5WB�yim���l&�i�Ⱥ���ϐѿX�wi5xGA[B�ډM��ŃT삩&�cF��� �,�rm���WJS,O��R�h��m�G��r�vM:�.�*:tt/��h��s7��$����S��'�PZ��z�R��X��]�o��f�,�&*Y�����]��j�44�����\�)a.��4C(�q�l�Y3�����|_mG���,V+�B�UH�=��R��.f)lpE��8�-�`[��K��2��,��A��2�����r�{�̤��*p`��t�9Z�]ٺJ�2mS�Ø�����7�p��F)Md���g��Z:���Gwٱ�R�%vs�2	����{ ukJ@�/kW8��q�+y������䱻�7!wQ:ɐ�gC"!!�Z��Gki	ά�]y��}MRz��ۂJ��zh\�2���	Zg.��գT�lG{X����+u�JlNZu��e�l��/�Vr����,փ����F�kS0��թF�bOY��+rw�A&�w9¥��+�Q[Y�]7
I��]�N��%�M��4U��O�"1t�c�-]v���'inM�e4����é���:lQ�#�4�fs4G���R5nD�2L�U~����E}�*Ԩ�LF�t�Y� E�"uט(��`�ɗY�)�[SI�� ��C�Z8C���K?o��dA`���$�[���`��R���0m[ZR[׀�j՜"�d�]�w`Xl��et�H)4���h�wl�F�����pG��-� �6���P۫�uϰ��a
�x�2�,�X�����R��{�1��1�'wN��0�W��{f��w1o���E받�3P�o�LU������C=Y��������P��c|l��ZIn�;!P�
���*eA���g4�	�Gw^�r�im;}��z�
����9fln�!�C�6.��T�p�J�Zt�]���%J��䠂b���
�sp9��і��5!��]%���%�[�*��`=NhF]Se��x�sj�b"��WW��ՊY�)8:�S����;gK�&澕��#����g�I�m�{�K�{sw=CP������K�'N��IM�[.-E���z��J���h^�u�+z*L}�<�7Z<�BT;]��g����/�:S^TP �M�"x<��|�^���r��.unT9U.�ֹ�Y�
�w%ͼ:IS|�A��ע\C�-)�i}2������[���j�cQS�.�oq��5��]���B��9��d�N���j�:K(8"�)�m�@Q�Es�d�Tnӄ��A�$��uŞ[�m�\{8�ή.����&�ր�uH%B�iN��J�Ҧ)�JV��r�ŖJ��}�"�3�q��P$�\L�	8��t5z��B7�J$���܉(0�%�p��4H<M8��k�[Ww6Q��E�n5�Ԩ����lzZ��L��j�xL� *&FLH"A
�:-U	"���k �e7�%�;X�& 댐�x��1�*�J�:�c�]��Ԩ�MfQll�Pu,\���j:�Nݽ=��������ָ8�y=�Tvβ��,���q���DA�L�ʣ,��Vk(�Zu$�yѾ5��k������Z�q�c>�}��ֱr�-�m��X%��s9*AřJ"E6�ff�h�m8�E�&M��O�''�׃ǌc���膤7֞�,ĸ��Z�T~h����!J��*ijYT*}:�2l�w6l�m{x�q�������ޣ$�m�m+��J��_R�ߒi�ѫ���y�"�}�'S��ٳf���ǌc����t����z�kD�QDkDWUETR& ���+mUեQAQ1���fL�x�nݻk�ǃǌc�0	3\�R���8ˌ+�*�C����J��*-J�(�b�(&���࡬�,������{�/��$A�#J��5Ԛ�b����2˔�(�TY`R�b�������}L��ҋ,!��(�X(��q�
��h��=CGi�Q�*^S4ي*��	PE�(���(�J��m\ۨ#4m31���:�<p5m"԰UR�j" ���T}�}�SiX�u�=�/��۹�FA�V\��V�և\�V� 6gz�we�`�BCm6ZNt���E�M��q�d�,$R��o��0�-7�����!"$ӱ��1��|2�S]��JF�la�� ��?{Fs�[��`.�b��U��Ɔ��_gs�X����@:��n�dמ��>�[��Z�^�;Ϡ�sE������Q'���	�Ä�%#-7�<�>g^2<﷊�P[�Wae��Z-0�{������y��G �7�3i�݆��`�2gJ�Ԗ���3��;�d6����czf��㻪��hЯ_��۠p�o�7}B���艁�3����g�]�0��]Ǻ�bzc�s�a+I��^���j���`����lԴ>�ElnE6Q�D�M(�&�Bu>���ug�<�~�0���G��3oY�f��Rr"�zn������F��w�$%_W��1�/�wﾹ�	�ف/��lغ�B��<P�I^��
����;3��ߓfM��6^����-�ELqnh�qAͫ/�pgD�jR�j��vsy��˺w9]'�Ws)U�ћQ_Q���+3�}����K�X�1�;�2�5�"l����Ouě�2�K�-U���;hTC4�ڃ9�.��{�5�"���c(������y�p�QYo
J%tQ�>���8zv�*Ӭ0^ˑ��2�[�ZHKRɼ���/0m'��� �|Zyr3��)M;f����[�a���C����VSS�x�| ~?w����~�헞��e�xh�f�5V�k�U�*r�I4x�J����w��>#���KC�f6́r������v��!r$f����� ��N, )/k����;���Z�Xq�1�M��My	+����F�#���v1��ܾ�������]���W�ot44��SM[�����C|��/=��<�3�/����{��c=�Mc"{Qc�
	�^/u�]0=!�3��ШY��ڃO�jL�i����,]��3��ķw��3�V�jDl�������<��ߤ�7[��KU��?N�j�o�S��6Z��^����z������:���ߦm��Fv�xD
]��p���
R�)��%ImQ��d����޾v�
`֪W�;q���ܫS���'�B��
=&�P�X���8��>���r��]��r�-=}HǼ��A8w����޳�ɇ�� �:t����Rm��K�;\�.���0톪�`U׺����Cbɜ�&H�%���5I��0��ݍ~�v���OP��z�E!x�[h���_<{�}� ��o������d�}B���5�Od�9Fu�"o��P��"�U{l�g4�gR���*2�)�F�z6:h��w�|S��!EV��,a8\Ξ���������������g���\�:Q*���n0��6�2V�}�*ڈ�w����/`3�*�����Cf�ޞ(O�w��&�'p���6Xƴ�؈]ѯ�ێ��cl��ӭ��7;l1��I9zZ�}���A�ө�e}�DUd���##i]��W��|	�.NQ�/��@��O��`�3y������s��J��^�IS�튦�,t��)l��˞1�B�SF�T���4Zsy��g��:�4�E�&�A�)�R�*b�((^�̂]�73��f��<�$�9��t��js�&)���'Uyzz6�ȳi*:�o<��vG@����t|<����0'��[��lr���ig8�)w*��&���/9߅�NsE�o룲ε�ֈ����:9�},:�7�O�e������M����g�ˉzY�l��x�H�ߍ�9�����B�������� ���) ���u����~�A{�G��0��=>q����s�u��pi Ɋ����L8�;MZM:���*Ƅ靚c!���KQ��A���,�W���}s�=��cv�h�L�Z)��1_C	l��U6��.��m��)�)�[���lk�_m��'����W[�;&�����yЖjCE�QM�욀��$8[��mJ��i�q�d3@��VR�MGǪ�1̋�%���:,Ka�ل�{OI��t����-0h��(���昈��v���{�^�B����U���˱�%?n�CoR��^Mg���۳ܮjx�<����5�ڗ��Bch
��bܶ#ukv:�f{mb�լC���8y�N^��`�����M+�
���zRW[�b]i4:�D���n1�*�Εv&U��ٲ�� �ؔu��R��Q�C�q{Ժ(�2{�S�V���1�����,��8�ŭ�i
!�zt�A$M�AE ����˙��S���swL��R<)�wX�G�ry���A�� ���3����ϧ�V�jOH9�i�@�$h��p�Y��Okp�lD�]�#�
�w��3�I����Q���8Ywn4f5�^
��e�z�/u!`���v�>�0*:�_*�|WE8	d�5LY�/x�G3�S{�'�y�46��b��H��'��F'|��/�/��u�2[�F\|1A��b��Xc�1*�($�����E��ֵSa'��h�Z7�!��z�0��,���ΨOј74���W�~��!���e:m��z9�!�Y���̪ܝ~7;��{�����U�x�[8�~�,��͢_v��7�ėNȯtq"��7��z/oRv��6�FO�O�Yܨ�����g����)���Vۻ�땊{g�U<S:2������	x������Jo^���?_^7y���~��h����2�f�C��>�E���}X���(�oX���"̎�j�.�VL�L����Y6m<�'N��D����Q�����㤸��/�����=�*4���{o��Ʀ��Ⱥ�R�gww�A^�MxT��ಣ�]�^c���a���Wo�]�4pK�7NS	�1R�������ݟ���� ��x9S�⭔�?��[vN�+/'5�s��"���r��K)���Wu�bT.'���g!�6U��&W�"�?�7��Kr�0k�� ����;�W�4^�=�3�۴9U����n��MO2��l�6��k�?|�LSsE@l�������E���{ڸ�ϷGuϩ]dp�4��n��Y��}���	;���oi�9v��<��#J�|��u������&��H1��y���~�"�=�0k�������z��l���I�hS��VwP��>�Gs�)E����o�z2�����gCt���Ȫ����Ӳ�צ���y�����nP��N��쉩�̈ӺR�|��q�9{�s`lF�.�o[����G��ET��-��n�y���m_V�mF�\=�#ݍ��"K����L�cb�C4��u
�r��Dw���r#֍�;Fv{�zp-�%��'0�����`2Z���י}ܘ��ac�o�|��O>jf�VX���X��7�B��D�W��M?

e�����&؆�ا�Y��z�^>�c�{�p3����V�s*��YwH������I�?'��B]�Zכ��g�o375\�Vh f3����V@�Ӿ���WlߠV7�8�T���X�6��N�q�T�Y��i5�PA��)M��D����/�壹�	�S���P��}O��n��K���L��8����^yV�E��^�^M4�f^��D�����i��Xy˦&� �b����ࡅ5hyK_�p�Wf0�Ss�'���G�v�3m���ÀB�f�� "�s�V����<d���q�i��-�gS2�)1�A�o �S��;�@z=7�l�G�y�u/wv&�ij���CO\��x|����w�͡Ѱ+��l1�����s0^mbliv3�C�:�[]W�¦R�^h�E���L*î�n�����b�-Q��>�B��I$w9	$(��z���6��=5���7�r�8�����̽��7c��,��v�U똴M�i��S��s��7�G�����/�gy�xW��Ъ�w:T�$�7v�v��%E�۸S[�fv���s�,8���wk���/�4�ͼ;��u`�=4���-Q��f�6�K�{��D	8��%�gY��v׈6�/h}����7~ݾ�nh�� �&M�jM2Y�� cz��NEG��w�ѽ���[��"�0�`'r�t,������D��
���9/a�8n�;��7�lY�Wg�䆥1{�/*<j�����R�c��pϡ�z1����U�S+�W�+�V����H��cx�%M6W�]�%�/HXj��7�.]������ڞ�'�ʵ��aj�ϊ�	0��H���!��}��ó�
茼���d�= tb�LףMA|g�P)%1��&V[<jmɾ�x�T�n�StS�{�90�^�>M��t���%�s\dx�у폢�]�(+�.�v���ٻj���k{��)��+��m^S���?.�㜊�/�
�4�v��f��v�,s���ۨ��5H�d�{�j��g�j��՗�R��t�m�[����7���A����$N]�4�{i�l�$m-KM�\CW�e���E��f4�r"�%-M�/+s� y�MV�L�	a������Y d7>�@�`{=\��_e����r����d*���m@�J[]:i�Nd�^�,\0�sȽF�����del��j�5���;���1�)�v���z��9���؛����I�?zn���X�A/������r�Sܮ]���g�͝�T��3[����b

��KL�]vz��U>���d�D��*�h��,�3$翼�Z���׮鑏��{M�a�8Ӏ)i!��r��9�5!��Q�ۅ4�"#�/\/c���CqWz���e�3�<oK��:r�g|���oy�ba���9EG��bSw��e��%��55��ڃf��-�f�L-��k���v����m��2�����V�$Plr�4�=�e!��x5�Fb�=�7-�9<��p����Qco־�˨�}�w���{�*Z)">��/n,����/KY^ڕ��v�;�6)�u�U�����׺���<r�wi5]k��j�M%�Y9֥i�\xw�da�c:D�חQ���5�1%��l��y�a;d塍��^�j�|����a���`�Cnִy������;ɨ�0�C���T�G�������N�FG���ӯ��0����E�ؔ�p���8 �L�.^�}�p���eJ{j�޷�}	M+�:;�}���s���/Y���>|�AP��D�zӼJ�hƦ���ލ�Tg�E��Y�n�ǟ�ų��W�v��["/�h�G�3*r�f���2��}˖GG��EM<�)�v� �7g.u׎u��.�J,����Ǚℳ�f��.���,���u�%/F\ML��v�o�{:����̼��O�E����5i�V�&C<O��xǎ�}���qِ�YF�:v�?��*�dh�|,�o\z��_�O��[��B�����۾���y��?'G}���������s�m�5'b�#;L����[}(>�������j!��{venh+;�VSc[�Ed�Sn̉�k����AЩ��ѹܙt7�c��V����P�OcW��V!�Õ��=}բ�ƕ�
l�C �.��G{p��w�������GV�0���*��deD9
����d�Ď:�q���ݒ��!�8���	/e����s�Z]�]�I�q�A�:���Zʧ��}]X7.�A�4&l�F���t�:�އ#ݢm�����m�����^u1�KK ,ꮬ�b�'�֝�B>��R�9\���=��m]�#/���ԗ)K�<��sVV��)�{����K{-ښ������+v��wk�5�f4�I�|J�b��S=���̻�_T#���Bz�	5DY�h��:B�Lo�q���t�7
CU�<n�	,�}�ղ3գ޵����L�C+9.�9΃�X��Añ[�Y��X�ԖїG�t�ā)9u)E/m��;`as<�w�B�ԙ�Jz������d�b#�bwr���A(�Q�K������0HU43gt����S	Щ����tA�3S�Mtl���S�y�ի;�z���$t+z�kDڕ�
Y�� ���.��Sd|38��+�G��MM���'!��Њ:�,�ZT�}
x�B�	5`���ס�H�4�w�yM����k`ͨh �jt��v�����������:`lT��c�[uڂ��)Y+.�XrK��E�o��mdh�#k��0��0)ݛ1t���S�۰���iU�}���1�M��l�����^�(�`�USSr�x�U�������2ŧ�Y�;-!�R�bU��b�d1Y��s�oC�{��.����.��.p`�������]K�CSN���Gq �.q��i: 1sf��wcH)��p���6��4��� J�s�iV�1�3k"I�]�&l��.4���Z7�#�����ۖ��j<��뵤��G3ܔ�o[#x������X"Y;97{Q�7��M1���f렛#Jq��M�;�\u��oh�N�	����[ȫ��J6,b%��1Y7��*vr��cʼ��C���h�K1G���H�B��A�V�R�⳶b�ϷV���癧��w2V��)8w��f=U����z�V�H7+^�܍��;�r�z�x���
�:IZ���>5�ƥ_,�S�jp��g���uu�u���uq���j$Opx�ַ�Q�/�kP�
��!i�2i��^
1V>���)�v���4ރ�}�#�O�_��A]�U�q�R6������ ��w�P�>�L�˾��:-r'Q� 3����xt�!p��b��dvv�༻�<u�QFإX�Z�V��9j�_��DU�Y����cm"��%��q(�'Q�6k�]�v�n>�<c9�NPXi�EiddT��B�X���[�ұ��X\�FW"�%�J�zǧ�o;v�۶�}<c=w53��(Բ�B���Z?f$a�6�V���D��2��ل�&�O�͛6l�}<'���y��V֊�T�1\EA���R�U-cQ2���eJ嘹.%-r�k�����ǎݻv�1���rIˈb6��+B��fTW1P�aZ�J�i�e)G����QL�B�ZV���	fN�ӹ�f�v׏1���3Zd�5�ri�$�e*�b0G[�Q���PEm+TS�\eN�f�e,Q�\��==;k�nݻv׎<c��kU�b���S\-��L��9�+���J�(�YYUR�Q`���\��ݸ�V)R��҅���-Zڸ�ʨ���j-T1�"y�0X��R��h�Kg32�oM#�P[ƤMk��mX��h����mDeZ4mU�.q�/E�6�T����jZ�R�fUc��)$I&x�q	c��Uk�z_r�:u����)(�m����r��u����1@�:L����

�\�sO���D $m Y��}���{�<�~��l�Z1�`6��b#zb9��C������籛��y#`t`K7������a�` 7j^�;�k⫎��kMc�(�yB��Q��~�a�AI��)=����\�kU�");��1{P0�ǭ9����lo*����C�?b��?<���"Pew+���о��I����d���w��_�[�@�����7�@�/�m�Ǖp]�&z�K�%�}���>CY��ý}آ5�;�Co��� O�k�@��M�w'r�=f̖��P0wzj-T��uU�ד�ژ�ӌn����������>��v�I/)߾/��Ҏ_N!D-g�����ꎑ��@���ZX������OR�EHFҥ�=���F��O�`����U�2΀ƻ�+`���=U߲��>����-����ϙ���M��_����?-y��в8���j�x��u`~U;f�_�^��QK&CDE���e�l#�W�J�4��5��@�(X z��4��I���u��Q��
Ls�őYR��OOU�]
� ���M���O)S�&�eKG���}�`�~� �#� ϯr{���EϘ{��Hp�����pK�������i�3�ǒ��CD������_�Ȉ��:{��ݎ�Uεr����|y�yG�E�k{ѯ��c	L'�2�I�>ٳef���|�P�.�^���oj��f���<��I�mEc�[�!��dRH�t
�ñ���,���SsT��C�oge�bX�� �����������HE�����j��Rrjw���"�ꅔ�6{گ=����0�M9���\l�oDއ�~��I�)5�l�	�2a��^��i�����I�b3`5�Z�[�G�Θ3S6�p�~�\��!����v�D��ЫD8�y�8mfU�#{�Ś��{�/��t�ʜI{8s�#���רk�Q��a���l�g��d	�FZ�c��.4��T0��x�gR��A�U�ٴt����ofV=[F�}@�=>�:AلK'*�`��XY|i�[)T���n?i��)����q9�I&��n֦�*�/Wj���T�d���4Z��cɦ�3�/*p���ξf�=�� 0*
�!�	�I��M���d�E�QFAF�)��5G��  q��Ʉc�h6�o�~�]îJ�##�,@I���~�Ż��o"e���ׇ�NKJ�d`�k����_YՋZc�uO�s��w��q�j�v�c�n�SM��SׯDM7z��[��FZ��m���>�bf�Ճ^�Iy*���9�5�����UU����M<ڃmG�va�;���ek��zN���ӾJ�mtsC
�%���TUw�ǏU��l�yʏq�؃��0��ּ3Z����Lֈ1%]eOp	V�z�r*|ݖ�eُwZ#f#�X=��Q]�F�R��ߓYY�W����b�k�=!>�W��<�/����Z��+��o�I�2I�Vu� d����v}ܮ|���0m�6�YVEa���B�d1��o��h�!�H�-/,KQ�|^���:v;���y�@�Y����f��?~��}[]`�%M� ǠQv�N�r���7�¬�0��t{�|]��7�m�3��ڜ3z������<:z=���ʃ��\��`�2��v�3b����x�q?9���S_�ۡy�(�|�5��5��pQms�b�faκ�Cٽ�΁�v8;���u���;]֜w���l�W�s�p�pNq'�vuÂ�f�ff��{��s�̸-���]{q]^�;���F��|��gƼ�w;�!)}Ϸ���q����� {=�
���گ�,���[�s���C7p֚`���o�%C|sׇ�	�V}��u�ŉ�T�܊�S�2�#�/�[H���8��U6����I
/�����36��ǰ�;��h@�{���7�o8�<j��ۍ+Q�
�oL=nH����n����&��̺�i���� ���c�m���6�ac���\qz�sـ�0�k}fz{�!:�+��۴�GlM��f5�h�p�8�{&�Kz�v�̎*+_�7{j!���\��t�u���#��UJߤ[���U�m����=������b{VfW�2�d�-����o.����g<��ղ�|����υMw�� :�vMJ5}-�YkW]޸��9`�wsf�"��`�M��8(A�f��Lh��da���<�N��\�9BTa�cB� S��G���3y�&)���[wj�F�]>����p��� a�a�`<��?m�e��~��O݊�#T��ZWO]d���y)��z��Wk=��ɻ�$V/.�����q[����W�B��ۻ�__��m�ܖkq� S염�����St<��0�Ώ?�^�uu��9�v��ݠ�W1s�6rOawP��wW�ؼ�k��E<��o���Ҍ���#���%'M�������e�#�t�/��#�w[=�ט�gh;���{zf9�)�vҎ��b��bg��\�|=AC�n*�"��x�,ަ�\�毦cd�6��usXU�~��m%T˽��sձ^�� ˝����
wPb��YV�ǋ���r|�*�Dq;k���h�of1��ҍ��l5\�uwW�"/G��k����ъ�B�X�wi^��łr��4�W6NnVW ���3��a�!� 5u��޴��������=`Z��T�*��u�a��5��/� &rt��]��tN'�M�-68#-j��W���0չos����~9N�h �p}8�3���N�._�hsr��a]roL�c�/4>��4�t�3�l����oMj\S��W�W�W��^f`��n�U(r뇴�v[������AL��:u��!�G�Q���I��6f�r �!�r�+k�*��e��N޻e�/SUj����V�՝�!�5;X��3c��q�"�g�����>hz�q#�s�6�+w��Cf�5R���n^�M�#�}�睸�^S�x�C,eH���vcÛ25G�jA��QA�J��-��>�����#@����EW[�0��T���%��e��-�Fv��떧f���k�v�>�˯w�4��&"�fi�Y���ltR���Z<I��ۈ�m�����z�tٔT�3M�a�7�z�g���EG�PQ�>���@w�nKA�:�/Ӱ�s�#����h��[JJ'��;�7��O>�hL�g���vł�p/Lf�RI��۾�t��3��w\z��lZIƔ�bϷ�q?���&LV7H��&�3nÒV^�Q�x�.�[HIxf$���:]�rq����t��7h,vTG(!�s+��o{g/.M�M�B�x�0�X" �d��n��;�m��L��|s�u��#k���	bP��r���C�����L��o�ڻ�,>�j��ݗa�hR�Q�"F ƜHc��p!lB\FT\.M�4�8�Ff���{�_���P�"^4�+� �G���ǻ�s���\\�{$m�M�1���e���e�jc�^����}��è�(��^�k� �28&�9�RXڛ]9�al u`m�^z_=�ݒ�r�>�j8��Ļ�*�æ��]W7�~�.��
�</���Y`�s"�}BA��Ş�\�:�)½Rr��C'��w6��H��L䌲�d2����w��v5�;��������@���]���d$^x��L���kAJn�j�{7Ȣ�S�Uʧ�qd�D{�X������
��2N*i.�˥UFb�����:�^N:P�,�s\z^��z�0iW��E��+o��Oz�ҁl%�lmU�c�O����\s�{ӷU@aǊ��bX����x�̰T\��Kp~j�X�5*����)
�K�����_���d�l�פ��`�Ŵ���x�턥��ե��;6���SRZӉ]�`��{+���*E.69���^�^J;m�͈VT�\)Q��j���[�R���ڹ��kO2���F�_T�{����&�]Z�*�Ǹ,\�����q:|��e����7{���^�z��zr��{��.o*%=���I�w�'���R[����4b^��GZ�H�ù��-�~]�ױ����ܼ��K��FFV[ּsU�ux�/���� ^�f;K�����y�ӊSw��Ξr�2ۣ�����>������s�㕵�+;L���et�[;x�d��MO �WM�N���� ��O�f��*���Q���uh��Wj;a*3������ 3������y�/^����/�([x�2�DTX��Eu���4)"���{���C��%�5�P�ɝ���*T�t���Hx�o�rvU{�7i&�j�^!W^z@ ����3���DC����^����aȝ�<�(�Ů��l-��/zgܜhC�yP;L�rj�(�;҃��JMbz��=>j���dzD��{\Ԛ���Aaq�<�F�X��ɘp��������rN�{��ˣ��Β)ǳZ�u:\E�:#r3.������3l�*#�E�(3��?u�G�.�f.�ϱ_>]۹Y}������Ŝz.u�g{��Ǯ���{g���:@ �9z�LT��]��n}6Z�_��l���S�^7"�b�zߨj*�]��D��G�Ҙ�����w&[ 5T^\Y��%eǶ�����=�]��J{�=}��T�C�xn��	�?`�Uj��/cA�f��o^obfuzމ4��R���]��MsV�d2X�Zx�ױ����/�Gm�CDCM5ݰ�0��Eh����{#Tʼ��/V.��W#J���x�v�ۜ�)���I���2��e��ZB�Y���!v켰�n�j��l���Ę��ƚ�h7����9�	�3G����v*

מ�W���t=[i�ƻ�����ܤ��K^kSj�W�5�9��)�I���K�;xwj��x,h���x��|+��t�8m<�j��=f�b5F֓:Sa�/�;�w
�@B^���HOw"ό��L��9���>�E��r�(m�o4Ǒ<ntj�ưh����˶w\Ex���>���D������8A��������&f¶Y!l�"/��m�Z�:}��=ާ-�E�R����6)�>��m;P��f��Eˠ��\�9�fy���ח��1ܧ�$�ԄnD��ƁɱO��(���������	���!�������򈤷=:WC8�o0v,, ����.�m�7t/U� �H6k�C�DM5��%���Y�n�`�F|G�ҟ`�.U`�)&��op�3biV=K�D�0nqf�i�}�}�|��Bb�D�c�'4U�l<���6�C�a��
�x-J\�`�# ��Ev�*odl��fnRf�NJ�G�=����R��{��Oea���W𿥜�RAzV�{_K�>�rr�z�c^�ɹ�oN��\�0]R�8����(�ܣ��2�w͊�Y�gf�XDgr�
�ˑ�[�t���fh�G5����FA4� �z�Z�s͕
�q��@{�A��;�JT��f#��-ӎ�֍�P�����`!mlX���H|E�CE_śOT�VKO)s��#U�d����kf�����|p�(-��{s;y`����H��j�l�đU��S���R���>��W�ܶ	)>���ع$���*YX����#kx�,c��' z�c��dtB����r%�۲���-͍�\P�}�G>�
N��] �r�vs/��vuI9moRU��%b��h�3AjNK<{`�j�H���V�c���Z�� h���x���yzT'z��X���]�ujݽʺ�)�A����ښ�L�y ��}ݶ�N��9Lg^A�����Y���ORz%&hU�z����_S��Jl�����8�G���ZrL:��{���V^iX�ь�}qP�:�C��*1j굺���D]!A�4�n��Sy��i�.K�8oE�*��3�-�q[�����Ѥ��-+� ��xu�����lSEL�]ýt��u/��㳉���@v�d����[
�N�.��4v��1�r6� 2�[h�k�6w�n\��o����	L�G�*��� �n�95��Dr��>Ա���2AV�	�uʳv��iR�Dj�#�r.�Ǣd�e�@A�d�ɉ(&�mRD[�Ӥ�̙J#I
����0ɹ���P�%����^�W��kR���m\%�0��8�]Y��s3	wCh<�0�3���F67�pE.�iO��"w��Ҥ�dr��O��Xn7�CK^�������2yv]����v5VK�^�B�b ]����(�KK�c�o6DpY��7kx]�7��P���ōԺ1;W=K��l�ɬ�}dނ��)\לV���Gr�!�A���q�k���ǐC;U4t7ҹ��]�J�n�|;75�U�����6�M� �4NY��Csc�F!kv�|���
���_5P�S��K2'.�*��
�M�;5�Z�J�.�C]�������"��� e����6�Z��u�v��Ш��0�f,��+��y�񏵵��Pw2�����;�}��v�<�a��H^�u�}Apk7ͪ�کB����,�_8��k���iȜ���L�zEwٻ�jj�ůK�$���R���;H9�n���>���TFn�����[�U/$ne�@��?>�72��u�z����n#�އ����������NlG�i�Us��9զ�..��6b�����'�t�S�[R,�^L��n�(�����������hmӒ��zbl�>@�0Qֻ���旍�>�4�:�+�+qrκ�m���2�< �uU�)(	`a��KL4a����@��4
!�8cf&Tq�8\'(QqE��*��2҉G���1$D^EN�A��1n�aD�M�R!1��L�)�� �QF#J�
(�LSTC��E���M�18�Qƛ�9�����ì��.4ʍQWM�&2 Y
Ii*e�"��b>GB	"(S��a���KQ�h�R�,mkMh�[Z����-����+�{��ZSs�%jˊ��I��&�5۷nݵ����cfrNh�{:� �յ�F6�G��$TѢ+U��Jv���\f���bu�����ǎݻv�<cNj#Z"�����Զ��2\̙er��LpX�Z��I�ZX���*#�L��4�6l��lٳfΧ��}>�g����[>���[Fwq��m�yj�c�*)���KR�G��:Mb��T�\�i4����nݻ||pq���':ѩ�h��4��V�A��]�}�E��ҙj���.Z���q�3�u��;k�nݻv���x�=���0�s3=k��kC.8�m+�)D&Z�wP�uQ����ס����]�v���ǃǌcϾ0KI˘�*UJ5`E��4x��DU:�]J��XR�\���k�ʮ�ᖢ�DT�����A�)mF�0����qM$w��Y�[��ks-k+��2�KhUV���)�Q�t��bU�+�r���,m**�^�]�
�[w0w.+A��n�J^<�����ivYͤf*�s8���l�Z�t��y�̂I���y\���z/.eq�ړ�|
��7�2�f!�Ϸ��h\kC�FѦm�q�f��w7�Γ��/��D'�DIs_��;�|�;Qb�y7�I�w{�l)pc�Lio�>"�{�5uC�].�̐';���N���n��׹|���`5ްQl��7��G�Z�-��)7�%f�wg�n���,!9;mލ�pəS=��1�FY�:y����v$���\U��b�}[��J`��-Y��j��v�y{YF�o#ڗ\6�f{MIWq���fr�����p$4<]��u��(��>a��6�1�����#��z�]��k'�Ø휹�!��5h>��0"�k��Lʶ�U{�ʚ)�B�uyp�����Y7}�P��(��HnPO�@L6�y�����z� ��ɘ�:���g_ve�SHL� �w����S�v߯�C�D���m���[탈��3��/��};�7���朩w^���m��beFIe!+f��0��;R_�iSW�T_�-��q#��NR�&�y9c��5��M�{4N5���V��@Hl��0E2���^�z�W"1�k5F�Z����]7�Kl���n�[.S�y��J�-�D�O��t!�$�r��s�vfM�%�{z�zՁ]�t��ӱ�jI����	�Ŝѽ3�Z��`����l��(��=w��>;b�yLsU�u�i|�PͪCW"���v<�[����3�Bo��}��G%o&�VZ��L�t�+�[r��A3�/v�}����.}��FfNQHl�QY��,!�4v-W�F{ۡƺl���h��9�"D��-)�F�`�ޝ�^�]�~�������W���s������� JX�w�������H:ޔ�t7�xk��{�C	[���R�;=�s7�>�6%�v5C��C�����Ƈ�������8`oܽ�nF0p�|�-t��uYX;M���bbU�Gy.�h����m�I��������Hڑ�"u>as۳e����p�wG��/*���5�6��rU� ��m�b�a��[DVBw���ł�=�s���������~[ӱ�j��{`m�������k��9|�ԇ��y���������U���i�9Y���~�ubݔU,���� T���V0��Kr�ec��$| � p�8z��,uY�J��Ns�YI������ܬ�r�R��\ƹbT��&+c�dG�|դ��#Lі��5Ԏ��٭
��5�)�_}3{ϖs�l�֛�,�"9MS��`��˽��D<�B\���-������qB�� Zg�>w����ﶎ߻��)vz�^��-H�xK�����_���/#?����X�	�Sw_����y�sne�k����r�}T/OLX�b%�l3��>���	h�Y��N�K2{�!����/�2;|�%G]�k��j��U����k���Y��2߸w8<q���|���R3��<�<�^}VҞ�I�;l���DT���uqY�"�Sx�>��	����\���]���$��9|���m�0��T�jx��\q9��v��L{}�o[:��^Ի=��5;�f3rfig�����n��D�yTt&0��R�u�6owW�udp�8�5@;�����1�M�|��v���,M��nVd�P�����2X�ˇ#��o<p���y�vܽTN���NR�,�gf���x@�W��<px�]���R����ٖ���������O�[�l����C^������%�c_#ղY�
d5�WV��(��j�س���;�{:m�߳��mw��{)���=XF�?����U��=�
�}��#p�Ҝ�b��+�P>�^�V�=,��+2{Jz���{=^�}�
��U�sƆ���>�2vg�<˾Z�����N�Ý?�{��/c7���ȹ�Y�v�lԷ{}��y�:�}�j����<Y�X���u�T{"M�(��3�s���2��2�О�]M��g���U��RW6D����n�M�3�>����#���݁ MT��gk`��!�.��
�Ў=��+c�1@z��3@=�B#2��m3i�ݭ���Ew���~=��X�YT�ޘ���
M��q@\���OV!Z�݀�b��]ӝ��,��*��`���a7ʽy'^�6���Wb�:Y> !G
	 |4�"ʮe�Jmj��U
4��@��Ӱu���S�)9�_ma�+�;':�Bܭ�1o@��g��ŝ[+&�ͷ֧����E���^su�Wq�ErZk�陬�����;�7v��๻̼�9s��"���I��nn���h���*>!~?�p�7��eR�ygz<�}@^��}�m���,3,��(P��w�-�C����ȁ��-�j�֜/_H�;�m�ު�@�����g��`6(���\ ��{����ԗ=����zj�g�'��Aew�bg`�TMBFF�v�\�n�Ǟq��#����B�w�؜��&Vu.�l��^�S� ��^wo]G;�=߷�U�ZXٳ;g$�Ƅ��`S [݅%��[=�n��l�[��Y�.�a����N�!�� �"��� ��������;���Rs�-���e3�n��Y��������j���wy{o������m\T�3}�W���7bz�ln؝�`�J�B���.}�p����{�Z3�M����y�=M����ן����叿I}~��#��2½�N;T�tz�z|۔7ԮL( �Y�L��C+�e���h<��F&�C��߂�Rm��ޛ&�������'w|K�{\�����U	�:��C�x�CH�[1P���R�{k��I��f�4,;�ƣ+��;յ>�xuw�k*���:��.����X�l>H!�'v��JY��9��~z�q��c�`�1�&e[Q����w&�����K�z%$��q������HH��}�A��1k�P��U��`> _���-e.��Y�o`�j)`�7����h�w��A+{��w���H�zzxǥy������OR�^�rU$���o��V<�ߢ��f��c<�<�u�w�ɗ~�Dlkf�ܻ��j��KFVRœ>ܶx��!�a�W����Qq���Uj�AO63�%����<E;��g;��)u���.׀/ ��@r��BP9[e�0�6��C/���<�«{z}��ұe�)��Zȡu��b���tY�6�[rBډ	��ǶF��;2�]���|;gڦ/�)�ٙ�����5��o§ˤ��]3Ҷ+{��>����ۑ�V�VPN��E]giҐ-ٱ[4n���s���h<9Au�^\�R�vp�ڎ��j�s�+WeD���j(x1�  C雽f�n��wQ_g'V6���;��ܔ���R�Bs�]����T�W���]��Y:����	&��ԃ$��5>n֦a�ۀ�gM�@��z�P]�_]��g<A��z^�gk(}4��}_H9���X�6�^�-W���UC���f	b�oя�w�}��S�=�q�$�w�g��7�ڹH��76�?`�l�w�����+��+EV�$�-�����Т�f�R���.��w׽�5�	*7M����n%��[Z���aSRL_�l^���7�"ږkW6�Z���,N{��;��~��V6�)�_��]H�ހ�
�\�M���*y��Z��Le�V���Ej�|*�����kB`�0�7�4�ln"$�u�fs�;MHs
��Uz���I��{to�-�����V��!.��;>}T����46'e��1�!u3�u]"��
⻞n&��F=�י�\�F�����{;��ؗ��H�& DM��}S�����SY�'
U�r��Q�虰��{���V�ze���5�+Y퇴�p�)j�0"�-��ᜊz�¯ X.!9^Ց,�����s����-�5�oo.��/��~���:��gYߤ믃�,:X.���X��x[�	��d����U���{���XWi�5F`�٘��l��T`&�v'�og����R��=J9uW�������L�g1a}"E^�
�[�@�'�����Ǵ���
ܜ�S�ٔ�>\3w=K?N��=u�e��ہTcxz�U�����P���X��v{m7����՝6yE���^I@(�:=��^֐��=����:>��$�E5>u}�WKw>���7��=�+	~|�a!�`'v��pODۛZ����"��Er�9�L:�N�����a^�@�|4�E��>��/�b�q��T^��L��Z�������o�`�آ���S�3��S�*��1���T��$�0/:}Ӱ�Ϙ��]�"�6_-�N )R}O�-ĕtdܙ�R��|�n0�h���"�7�Q���w�St J����;Q���?�����$wր��W�ov��o�.���M���o+7�7��	x��
h����n�@4�B�*xUbŜ�;��r\�wv�]E�w�!�+�+٣�^ǰ������Z����h��G��Ρ{DL$��D�A��mw\�0�?̡��7�^������&{kp�&T�g�~P_&_--5v��Yt�-y�Nf�d���ʘ0��۞� j����C������"fQ��#\�z�y)�K��#O!�K*�q0>��LgW�SG�i�W�f\�a���{���M�@wwKFpgG�7�ZLvY��SYڻ�f+���{/+t��꩸���5S1vaJn$����J�k�������f�%Γ���TS	�M�9���&,���Uff�P~MW���&��Kn���;	�h��wf*�\�Zæ������3sd�Nީ���k���\�R�WO]䁛דJ�O��@b.����S��5a�D���}�&$BK�� �7�҉��VN�#%��'�bT��m�4<ٻ��Jt�-���g����7}˨
X��C��E��T��g�m���L�U�E`��aZ��*���K�H[X*��(��o$�ݽ9��*�9⛧z�-���7�!}���<�c�3G�uu,�����ֲ�4wF�H��3v{:�Sd�C���[eXn�A[������'w��Y���`���A��@�N楩���pO�^_�lWD4��ݠ��P0���oWO��4���%�s�A�̸�e��k�sx��P����Xң
���E�],��L��$�Y�\١uyFqї]"!����]��f��|ńj��̓9џ9�9�>^��7b��Yٰ�Y�8��4ly>������)q��<�w؁��.mNu2l(�C�wY�Yg�I��Ä���sֶw�W���ͣξ-z�KJ�����·�t�`�v};}�����+�-����>�5��z=�w�Lo-2���@k�y��Zp�Y�5����wR*����Ɓ�V�j�{����럼Ǻv�wb�b�A��A�9~��<y�����8y�_��g����e��(��X���+�w�&��}���Z�r���ɛ�:ǅ����>�6(E�E�M����txٽ�ʞս�b�E����c7I�ʜJ�ux{	�p��X�o�'ғц7����;����rh��&d\u�;��l\�C��Ӽ��;_&;\b����n����f%
L�N��_�v�뢬qɠ�#
-ؾ�1��q�y�\EDe��;4пh��iI�k��҃���8�u(���ٸ޾u�ӏ�Q��jC��D��ʶ�yR��j��tJ�qs�xZ��1ۻ���l��/���n����C���;q�\.�ķd��h��N��Ǧ�uy�]{�n�rp�$XB�����W��=Բ�s%ɣ��/�&vZ��Й�u�3E2���R����
)��wu{�:T�1gIV&��������i����Dot�kT����t��mm`��:8\���tYv����)��тjga{�ư������fl���	�[۵ͮԅs���J��/� �4�3S��zڏ{�����/m_���SU�M�3��uդkbnd�r3+xm�3Pr�`���4���/���&-5�4f׏-�a��-iT�vV�;�[7q'jRx;��\�nn�\Ep����^-ۘ�J�rS�mټɥ��V��t�P�qT�%�J����AZ t3l4�<Iف�˺������u�y�
`��˥�U`] V+RJ��K�]�8�A� 
Z�< �[J����z༰�DuGy�]٢>�6�S��y�vJ;�05�^{9H[��@���sYNeMI�˚�5�Ugv;%���8�Ǣ��[�nY,�\Gc#O��౒�mL{�9sK��p�W��7��� OmT��]��vM��gۏ������{c}���+>mG�o��Nԓ3*0�5f6�I�d�I�Wy����7��\v�ob��p�wS}ܯt�bZ��n��&��8s���{";��s)��.�?�=��=ᇵ�lW7�i����󙙉^��r�E�i�:Oz�*}SD� ���H�n�>cθ�[;�^W��R�o:�3dwXj[�.5�u�+V�Ƒ�rI��l� �n,�+;��,.A��,,��Evg<��-���J7ƞe��3]7/�3���u�����_r��+F�� ��m��]u7w[�L�)��[�[��]��K��̽X�%ם���tJ@S��Z��Z�
�7��Yi[�
���J ��`ʶ8�Pu��|��p�ݐ��i���Md��u�!򫳁p��s��P,V����6�˛���_Q�F֢*Q�8�b	|�i�
Yy��c[+*|�1;�)����Z�nݻv���8<}0�k'P�kl�����]ƹX������̕-��U��ՋjĐǡ�ӷ��ݻv����Lx<p��?gى��R�0���FC��iE��� B �	���ŢN;=;{|v�۷n>8��� x���%�"�O���&8��PP��Q|j�hͼ��[��cӷ��ݻv����<9��R��-��V�b����EX�F(�X�QYD�DCm���e�۷�ݻv����<8d�&��m���Ԯ��*��ԩ+kEj��*6�a��d��u96lٳ���Xω��ߔ-*��Jf����T��-�˗9�eH�ʓm����:(ej�m�nV���J8Ԍ����m��
��R�R�aQ�*�S��[[m��j#[JTF���s1���J���lUYFV�Ŗ��-j�J�+��R�eqX�e+yeu7<|=��μ��J���]�[ݳf
L����s.L�.��{jԺ5��Kͪ3����%��;��3��� �=�dN����R�{�w�	��*lgg���.��^7ky;��{+�]\c\��¬��o
�6���i{*��A���vMwc�6�9�-�6���dR��ۮ�|\�<�'=���u���1ٔWGQ����A|���j�k34Y���,�����j{�sWt�n���'Y�RFب0���cW���ף�1!��|�[����ɘ��=4����,4#���A5Lђǀ�j�}ņ���3hN��0����M���C�V,}���ܽ�.{9y��c��3�v����s�C�/N���<�ѻ��g'�'4�:��0ffk-D����>J�zB�nHm-�� ����6�h%.´�a˅���ӊoӘUA0+ۀ���F��������k��`P���P�v=�"w��>����Rg�\Ssjl/L�V�XLT��E��+�a(^E~ǻz�zT�a���2P�rc�����MѡGGuEZ����x�'u+x��$����%��i�&������1gk8�{���U����W��@�8�@���³r�i��B���-���q~�pb��v/}�k�1�%�Ѻ����!���y���%�fOy����g��Q���i�>ơus!�͙ؠ�y������T���p�ڌ�\�����|�D�
[#a�Ǟ����.Y����y��P;\��ݨ0�c	 *mOo8;3JX��qp#5f�s�&�7�h�����c��*������J{�s~���˪M��vm�=1�:rC�k{+K��TjUc����Y�ynww���]���5tC�:Z�R͛���<�zR������� A�٫С[�ДFKGR2x�u��kg����`�<�z��ݏr��Ԣᤎ���.�=�k(�d���JU��f��	���n�4`�tC�K�
Q���V��K	'�ⶤ��1����'���_/��J�e��g�l5σt�$�IV��?P��g�\F�a�f�|e�=�[=Az=���{ò-w��(��-�>�#�"�qq4^��C<p������,�S�XjZRQ�$q�G�A)C����$�I�"�>���ԋ�����K9w*�B�93Zp����|�[�IJ
�b�w�o�L˺��f�e�Z�E�+r��jk�wV�扆n��3;�R��f�ޗǣ:���� 8h�X���聇L�G˧��aX72}�3�Ss��^r."�c�V�i)k��� =���Xa�0N@%Z�jlh{�[їIr����lH�j5�g=q�X�ީ���ö^���u��:QT����vA��oޡr+��v��\u��]g͕d�����.'��˷t�/"���h��&ef�K���8����6�D�7�=�@D�]�|���rKt��+8�o���!9n�Y �l�4�ٷm7|����Ðb�\[�6��*�6���W�����e�2#��W4�� �֌{c���{2���Z/6��A"��P�Q��P����c�}pMK���]�^�&R	��DE&[��s�C�^�Wx�	�$Cb�o���ê������y�)����c���l|�7O��{D�Huc�m�l�v��_k"��o�K4���u/��`�����Ng����ΓE]!�o�0zJ�Z���>�w���rKK{�'��g>�N����=�������=k+i]��h�oc����W.�}f|��m�M⭗�S�9�sg�@I�=ǆ������oU��V�v1^�ݻ���r�ͩ�Y�oOwO���[�������W�*-����_��A�uΎ�JrRP�鲛{	�/1�P�q��yG�җG�b�kٛ���F�A��\t���A����٣�s���H�t��:Ϫ�37I��%��̀`�5Ǡq0绪K��9�S[횢Z*��u��zV���(ov$��U��~���F����4��dr7p�Ys�<��sF��ߥcfa,�7n�S������x��9�!��4Ez6�v)������<�
ߐQ۱���-Y���ԇ��}�g;��r$��{9��	��ޡ����D��6�A��%���N�[�0�J���q�C`���x��\�9���^��Xeh����w*�q�#��7_��ޞ�MY)�oؖXw�u�@>�{�颔�"�H���<>C�x��zuu ����j�r�zI��R�^X�fԮ�`g|Eށom˨9�*�f��=�{���YV�h Q�ª�f�bnv���3����4zm�I��2nM"��D��o.�_�1�f3�y���o�MT�׳��R��ۆ��HMv��wM�
ַH&�� �>zM�8g]~�}�8f\wM�v���-�1��<r�)q��mֻ�=�ϼȆ���49��8�����������Ɲ����мa�Q,ĳ�s�4��R��>'��^���WuAv<Vc�a�H���b;�E�Y��㌒�M��r������˸�g��;h�*���Ur���ۆDJ�*�
�Os��&�=Q]��k��iq�J��`�bu��,�|�Nb���k}�߽a�lq[m��c�ٻ�كZҗ�!z1Ȭ�H�sm�G�)���@Ob<�Uֳ0nGՉN�>�;O2�&����|�儚}��*�6�t|&����=�������(�!�"
Y�nK�5j�ncq$m�i�Ä\��"���:IX3�]��PH� z�{w���_
b������R��ښb�>Z���hNۡ#�z���d׉񺙌m�L5�䶵Ҁڰ�ܩz%�d| �{�<�=b4�b�#�Qu5eI̫�1�@!jJ��P��~�[q��`�u|�7���*�{xt�:Q}�u���q�#�U���r���~Խ1�Vk�R�˦f��gi��[z�F�ݸ-T6��T�=�OU�tj����a�38j��ہ��`��ly�ڟ�U�.��S�_>=ԍɜ̵��"q���}�֛(6�Z]L=t2�|��m8�4�gb:N�ӑS��
D��q�L�c�E�ws��V�vp*�0��,�w�@�l�C�^3�Y����-�C�=��nj���Ӽ	�j2C�D�l��6ǒ�����z�2s���Z�րS��=y9o�f�mg�k�����L��@��ʊ��wV�������x%�wy!B )����"|����w@��t
�M5�]�z�z8代O�a��&�?U<Ȼ'[8�~����iR�g+�Y�Rz���KyU��S���0Y�\6-0�7�xD=��|��s����ZY�4?�yz�9R����㦯%Yc ��p!�>�&��#x�׽	�f�N6�f��skr���vg�ۋ�P� �:�wD.�}�έ�Ҋ�!�"TޖgI�#��8�w2/e`�߽���������q3]�v+n��
U�d�����G�m�2`F_\��LD�QY���٫Jy����g�B�����y��^�e�?�}�(��f����DX�� Qf`�X(�M�Ƨs�l��U�������l'�a+���]�4��.��i��ӹ�tU,qޯML�16����orA�M�}��"!@y����ӛg�����T�{����05���2��>�O���v��g����T!nȹƮj��FͰ~��˚f�rf�����R�������oy��/wC��; �f/�k��a�3w��읲;F�m�3�|M�z���>-E����V[�	tH������=��̟��{œ�V���MC�#�հ�w55�XL����]綂����ެ{rM�;�۠�Lg��ǖf�����J����]���({��oK+=��Mo
ڻ@fU��9�fy�<85Ltf^��������EGՑ�f�N�;fn�Z���>]w~ zyǃMV#���ܳV�U5w_��l���!�F�~���?��m��p��K�6>�OLTǼV4��~SZTI�]�� �Gw'T��3�4��w&�5 ꊷ�t�t����>��Ù��*EAVl�8ZZn#�Iv��Y��q��r�p��j��6��5:Xutks�Se*k��9�tޕ)U�.o[@�n���z�˞Ȍΰ�^��Pf��x�I�1�������"jR�g_�[�zLHJc�Ok��8r��>*��~���L\�A\M�ZE�Y�zR����i'��Uv��~�XcY�ș��)�\қJ�(__�/GDt�v���h�x��^�;�o������.��C�U^�X�=׫��p5���,#_��D�l��PO^�Bó�u�DF�b֎2�מJ�9�n��Q���~����k�3��-��t)@�z��j%��IR�韵��ent�^�a䋯��>�o��rW/����a)�̗]�7u�rw޼�9}�ȡ�'� �'��@��}߻/��:·�;_
�Gn��FdC�5\�mn˥lP3�h��RO',�i�-F��N�9���y�x�rtbW�>�r�&܏jj�o��r�pǐ�w��'����ux�l2]ܻ�r{�e/)�J�x������''q�QW�1:͙3��A�p�P���fx�:F�@NW�̇rjY�5��}�v�S�`œ��&;���;m>g��Sz�_�}��]]wOs���;���/;9Bԟ�Һ�6Rm��j�a�6	ǿ}��	��s�v3�G�0�l�f9���['�g�?1����o;X�3��=�#u�ϒ��eg�K
�E��nbliw]�)�˦]�NI��j��J��JV�z_ ��g�R�F����Be2���(������Za����+�㮙��l�5W�G�������N���nC{xr�x���H�Y�X�H�����x�[v�F��#�)�qd.��A�
f�G^�&X~<j�*��J���T3k���m��g�1���1J�k]u5�%p�J���Y�RL$ϲѵ)�]�̸;"cp5<��Ml�,i8.mHlz���k3|"��!�r[Avf+R���G��̘6uP�WQz�N��/Pyb�Y�~�8K���R�C/
�w���X6���a��a=[�{�e�>d�5��3sy�/��f�����r|�_�x��Q��Ue�SR�c�{��Y�dʏ���VN��!&�aE�|y��z���a�2Ju�����◦�����1Ӛ�	���� �������y�>�(ho�ϼݤ�OL��C<���	/)��c���*�n>�ŵJT��(ԯr9�&bX�IR�*ưf�Bm9�7��x��ѥ)L%FO�gk�2I��|��A����ϰ���c����>�m���cq�6B��:��B\u[�ѩ�N�,��f�s��y������oz�l5��P&�ݩ�nn���f������Z�x�ZR�L�o�X1�S/ D@~ƽ	m�?fV���:�]y����l�����6�d�.�����������ZG��*��� ���>����A�b������ttA�3]�;�.�Q��E`! XA��T`!X@F�օ"�B�B �,�,%��h� �"(! �W@���P��P��E��@D�Tv D����Q�UD�! `!`! `!@`!`! !7��$ �� �� ��"� *"*  �"*  �"�������*�"�(� ��"� B(�@B
 @B +(�B0�"t�Q��Du�@!��B0�"�B*0��"#�H!�F��`!DA���A�Q��z����`!EF��@`!H@F��@u�ң �B
��"�@B
���"���z�~@�g��*
""�(� BH������y���<������=����@���@�b)����:�˿��=�����@� ������O�A��("
����������ܟ�_�'����H�AU������������?G�C���`k�~���Mk�t����EAUIB@TDTVDAQ$E@�H�#!$PBE�a���A`��V� �Q�E�$�DY`F !b�Yb��abE�X���d�@YbYb@X��FDX0cb� #�a`�Vb�a`�b��E��E��FE�V�X�1 F,�0@��`!b@X� �E��$�`DXQ���`@X�`�XF$U��0,�b�bDX�b	 $Q�`�`�F@X�DXE���11 �E�U�1F��Q�U�0DX@XV@XDD�+d�F �DEX�Q�DId"HH�IET@E D������*�*h���������i�@������ ��**H
>Àk������	?����~���_@���A�h?/ϯ�>�:�~��O���?��M���PDp??�?>=}�Ȩ�*����!���}�]}�=P�(�������[C��'��A�����>�����t�ڂ �>�����AU�CĐ������'���? ��>O�������DAV���?�AU���}�	�~I���x�ՠ���������õAW�����4����^@�?����3��DA~����`�.��?�Ϯ�����?$���
�2��h�8�� ���9�>��ϗ�e(JQU(�QH���Q��QITRB��P�� U%	*TD"�
�%P�TH!J���@ET}]�H�V�Z�E;U۪&�J�e�Z�m�5Y��6�5�ksu2�n�I��kX�c(��9�';����e�ZՖ�g9H�ٶ��n]V�2�Me6��گ3���M������+�u��ն�
���ҡe��;us(kA�;��/cf׸�]*JkK2۹��vjҚֵ[%L��CP�$Jf�V��56�wnS�r���K�  �}��ݥݝ����Փ�Nڧ/f��yڧ.���*�����{�����n����'Q\�s=�oEگJ���X��V��^ݣ��r��j�n�ݹ���cl]��͆�N㺒2�X��  ��B�
.�B�{�����(P�B��z�>�ڲ/��+��mt*�ֺ�l�峯!�[^̮�m��w��4��v�U�p��m�ڻgU;m�W;��Y�כ޶�nֻ=5��m�6���f�CL���  -}+kk�V�|N���wp��y���ْʛ9=�][{�\wn�j�V�Rgk��7���hr����g�T���N��+v�����ws�]m^�k1�V�j���I'Z{�� o{�4�Q�j�jUu���{W^�U�N�[g�:���^�^�V�v�g�����cUF�/w��������r� ;�{,��/eh�kU�
Zͬ�j��  a�>+�Aھv�n��b��9�ճE�K��t�vru]۽�������w�un���W�]��]�j�pz�F�����z�]��ͽ���V����(Gf�n�  ����E̬��e��1��Ǡ�p� 1�5�����7t 7�֔ �{� zQh� ؆=z ���ڍm��u�����m�����  o�� +�%� ��J}z�� �  ��snu����x �]K� j�@ �u��P�4m�6�ƴڵmY��ť6f��|  7�  ��u�@Z [��  �Vր ��J}�� @���׭�4ڽp@2�CG])ol{wV��Y��:�ZV�[�_  ݾ� �}�ׁ�ҁ����Ҁ�2�  �w��
 j� =S�{/n  7qҀ ;u��);͜h 4{��ٚ�l؍SV�U)l�->  {�ݡҔ7˂��=5�  �X��r׷��:�ۣ� Q�7�� {�q@S@0  ���Ub� �)���*R�@ �{FRT� 4����2����6��Ѡ���R�  �lѦU)P  ��O*�@ ���~��_���7	?�࿏ⳃи�#\��0����?Z���}��������|>��۾���^� T�DDW��
����*"�" 
�y�W������������$��9���/?���FMSo�+!�B­�"�26��
�X}�*�Q���;��T]�-�	%�:F�O�	�d�y����t2�)]G�m���`F����vo��l���f���.�M,Zh7����$3�Q��:�Ǜ��
E%��7�/PØ�N�@Ne1$�5YmZc%ZrF��e�L9n,B��3ma���QH�a�V�Ϧj_)y�ƥn���5��Q;Á�bj��x������֐>SX�7.�Ō��/��J�-��{��w��C�,HQ7"0��wFi��.�N&-�*gd.ʒ�P��c��K�J=ʷ�^!��"��M2��w��[[f�Ǆ��뽛,�wJ)C %պ��ݭu+9��Hc�Й���x�R,h��)a��5r�j(��6�;��n��P����8��tM��T�p�r�ڣoj$m՚�f�k^��Su�ǵ�t��4��Sb7rD�Ĺ��6�\̗q��*F�/22ĺ{���c9���X�*n��2�]̻{z�����̨��n�\gh� �UDB�,=Ԡˤ�h�����[��Yd��7�J�w����{�b͉m��jZ�K/Ee��1^�HI��`ƝX;(ǢB��lflV��[��*Ǌ��U��yD=: XԱ)P֙XXop����K�0*�]Z8L�)56Z������4�����qX�sb�B�Q멢��l�H<���������RW���@���<5�n踑��ke	���P�����v���9+"�@J`�^�mF�09����:ʗ�e�ͷ{�&����tP)Y �(,d`B�n�F��ڽD���M�2��E1�X�J�<[u�v��Z��ˊ��{i�,y���f4��Ũ�)��°1�̦���}���LU��-:���m�t�;;Y&�����V�1����z�^��e�D,ە{�j�P�n��m��"f�Jn��̗�@�5�Z��y���z��I�՜����ЭPOJm���Xy�f�a����nt˴)ʊf�,�XSf����6�95�[G])L�ۘࠆ*�{�
"�t�J�Z�=�M���^|5P`ǈDe@n��2]޽˰�Ɲ�{W
�X�	�Z�%|k�Y[� �j�*�\Xv:7��HN\*�a���Uy5����-���,�ٷ���2�n�w�m�,d�q�bZ�
����Z����Sh�q�pj�L`��`�;3Aa��gM�Z��B;�L��7H�b�pn���ie�1l��(���	��ݸ,�(�f�4+iH�m(�7`U��i����\i�#�z"��p#0J:�'!e��ݍMd@��eu�Qu��;m��P*�j�('*&�(�Z�f&*��y�έ-d�j�R��`D7v�ffe,3%�.�f�����eJSf̫2u#j��Vc�� � �S �lj�*��A�{Vnɵ`c�N,d�	w���gh�V�Q�V4p�{v1��C�V�������
tf`�ۈ�-��g�N�ʗAAy��¬�Z��#հ�*��m:B�E��R6��5a�؋�&1J�P
��WB7�!�H,��U �л�H�
V�� �Ѥ$�aҖ��Yt�Ue�R�� �隐�$i�n��L�[��`&��a��$ĉf�iB���7$``� ��i��l����m:�F��Hϭ���� mʼ����ʒ�ͅa�:RB�ܵj-�&8�݌V GZ�Y����-kb@�V`��ًIu,1�`�)�����t�C
�ɱ�E)c�u7g6bwi�����dM;�����9C++^1��"C4����S����u G�Y�G��#=�J?��y�I5����K =Ǧ��H�l�`�*h��lF�+ �Sun+�dm���5 (�/h-c����ӛMJ:,���NP%�ֺ�MۗF��!K*� �v�а]�Б|��x]�4%��Lj�ʫS���n��dr���)ABӰ��]�[T��en3�woʵ�Y�Q�1�4��d�:�͊�9	��v"�ZJ��b�A�l땘��b4í��xr�n�s�!�P��Yo,n�+�T~�j�i[�Ѳ�Ʒt�aR
�*�魡N�mMN���Z݅z����X�5RY-�l�k����O ��k�SsS��yL��,:݌ċ����E,�����e^2nT�JX)Vi̳�&����֘+����Z��4ȅ��,x��1�ߍ�fkÒ=�S(�C�x�f�8a	�u�n����{u�M�-�(EX_n]�N�ɒ]&b{7Sc�82��'�zcd�`3Ϭ�Uh��ڵA��҆���k��v8��� v�G6�me2�Y3sZ���"7Avʳ��$�jl@��9���-43R�Sn]�()'4�b��oq�ͱ��l21�3O1��m�;m�1�Sq+�5��j�m��&�&bF�EkXN�V�ԫ�lX�Զ(P�/��PYrŝ�gDV��`1flT@���&�#Y�IFl$2%#J[�BM7����M��Y���!�eEFn��1Y����Ψ�*Rv���bJ+l�l�hKU��tY�9�r��R$�!t�Q��:���(��j��N�/^���T&2p���*![Y�h�I����u�l�!�݇Nn�	T3]7GSE}��c*X�Y��K�J���Vź�wE�F;���]�@�j�q�Ҙ�I+1C�e3��iR�Q�d����M���WCq:�N��3)m��@1uua�ٶ)3�����v5iT�����5x��Y �N���-��Lh՝���͂���G�T1ҿ�������G��]J/1�"��]���m0��;�ө7m�V�Z��JW�{�m\+4dVR��ѹ"jtJ�T('�p��_�Y���Uu4*�����y{���kg6��I�3�),���S3l\���3YS3��@��IgVEO��v%C8�p�C�!`��ZD�nUaĵ*4E�EV�ffM-�TQ�)��r��K�(�����4R^aWe�d�AS8qH�0c�4�x馰5�$��2�#�m�;L$.$��ub�U�i�F��jMgUw���˽9p[�m���p'F�M���]��pC�E>�Cu*5d	̐b��RUʌ�\�/�xU�ٙ#հ;t���G#E	����\�]�A�p-9��ӈ��Y�~n���R��VJ�����%n���!V��pI��ٱ.��r�@ͥJ��Wi\R+�1�����鵒���g	�{7\�ì���M�(�2<��wK������J�=�B�.^]k//3^`ѻ��/(�*��0i��`y���uj���k�q�sͨ�̫�o1:����J��#Xr�7*`;y�Vdڏw[��CLcY(���1�%cQ�
鯲+{f�@he����#ŇF�T ��U[$�Hg)4ڷ5J�
�Ǔ�H*́Y�	EZ���$w(Ec)P��)5�Q��3�������m\8v�b��DE�7$�>�Q���
Qz����A���iҔf������f�Ra�G��<Ȩ�4���t4�b�6���l�8�Xl6�8�C�X�u�qr���E\"ݘ֯�ţ@��2�[���ReLvXM�{N������$�뚍y�VT�î��� 9r�A@"��m�GT�2��n�PdݢO��Q��oUMͫ�u쵁2�����W��޼Ճu����F�����s"ݲ��ۘ�"��H�`LW��/0�ûsaT��A��)
�w��(E��V��  �iMǚ��4�K��u���gѶ��w�l;*�l��Ф7�G�w4��7�Ԓ� �㼛d����	�I�T�e��SU5����#w��1��9��#*d4͖��&��-�t2�xӚ�Y��C�VMM���Ctu�j�d��[k	�)�Q���jm�9O��b���S���A�ۏ&70�^fѕ�_�8�?n'��o�0�f�����HKѠ]Y�)��64Z�*�k�wW�Se�G���ۙd,æ���H���R9�f� :��4�`������&�q�����6=��"�;[�-c�`�lCDkD)l��a: `��v��0h���"��Uz$v�j�9B�Q`�&i�
���r̻�3�{,c�k�C!�+Q�7�0�
�����M4&��1��,X�@�t��q8�9K5��Q�W#;�/4j"툲�[�2�X�IL��uT��·�Ҍ��Q)C�V��y�O�V�J'E]�CO�C��\��f)�Pr��E�����"���&�:ȋ��5�<1^1L<�^#�U�����dz큨��u���Sl�`G�
海�c�l����B��	�ꤍ@y�ᅫ�Y��E�`<�j��6����[2��s͉�
7MiF�r�����6�0%e�1�7W�l�ci͚��P�2U����{�C=�C�ז-�m�-@M�u�������S3R^�ۉ�n��`],�Q$+#�Y[����g6Y��$4��� ��HX�C�����Xu{�Zx�j�r�YRgM�6�K*h��LeV��Z?؛WI��Ed��:�Ħ�:t��X�� ڥI�Y�[{��� i��U�ى�wSh��Y����C^,A�[(�	�vLj��`V��Aʲ֘�lX�J�R��̖t��ef�֫r�1n�y*Q�:��p -2[�� ��b�5Sr��)�6�ѫ��	�[.��3�(3�y@m J��^e�%|�stХx�"K�Il���j:��P�r��u����u����^t�Y(�9��$ih0<[WeZg�m3�-�A��tq���X4홬�a�f���v,���J9��w��,�FjQ7R%9Y�Jl]^*F�ͤ7%�/E�ݦ��8(N�t��cw 4�&��y{��<h$�1���G%�$+�a)M�'�ԏt5yr!�C����o(.M���[�ЌYt�,@	��4��WM�	�XoB[y�/~���WXi��)�81�V��J�u��N�`r`"�V�S�b��jƚKR��pՕ�"��[�`�mE�����xe!*v�PЦ���ƞ�N��+B�^�[I��w�ڰ�ðH��.���2�޽�����+&���U��7	 �n��vp��,�-4N�ϲ�6�F���V�)�6@�"�WW�`Z���"�#��,���w�yv�b��F�<�}�X��Kei�m:uw{�ޫ2��M6��c�ַV;t�s�u�Q�:����  ���[/]���nQ.:,���d�Ohi64�3���5�l��8v�x��V\�bl�,�{w(j�7Q��$�1|4��#�j]�BT��6�:UwrƱ6'N��Zq���v<���Ű�&���l^������R�&�p��p�wD�Ef'�n�~U��uuOf	I;�W�!>9� ��<,��[��m՘˕�%$�D��+1�h�a˰���d��M-��ݷ����%�M�ccK*g��6�Ю��'%��{��kY�w��(觩�@�TV�9��hfT��	
��[hj�ֈ�����/^��(���51r�D�ҊG���M�p� �H���w%���j����czlmul�6�j��5+�l���E�2��s/H���f���$�
���V�)Y��v� ~B,�B��h�WmTX�������ԫh�V�!K7�5�kA�6ȶNJ#)n�e�g1�p�"Ĉ]Ju�����)�֡�ѵ��"M����h�i��%G�0�ګ���qiU��y4�ma]�fa�Z�����&��f|(��4l��a�l�X�r�pme��ԬLp�cU'a��X ^}�����Y+#�b�,Ց�f\��]4-���b���r'b��`�ա(�t��4���Yz[��t�5nٲV��yg(���[�Lb ���*Sj���z]��(^G�J�ʃ��5����Si޼y�kE+�'�f+� QQM8+&4:ߤ.K-@�t&�ttFHsEd��JbcE�y3MZ��t��X\�D���3,Q�,�+����c�nT{�c��ĵɳE^h�R&A��25�Ҷ�Aj�*��y��m�;���̬�2�ʎ\u*��6K6�G4�kd�F�M�.hU!�/jʛ-e����f�U˖�&-�@YPb��F����LL٫�-�D�2,���F�Pi�I��r_��� ��h���4h[�oV��(��4]j��=�b_ģ)�2֍�eؙuwN6�-�q�Nj4�n���s%^\Z*�Eu,h���Ss�#74!.d��n�am`�]\8	���h���Vi��'Z5:˻&����5���BH� ��g�Z\�Jdů�`vN$>����z���U,&�M�WX�j�J�6����0.�d��b�!o���H�kx{b�1G0ù���*�
�NY1P��5�n�Ŋ�x�P�	��][���^�]^���p�;�m����f��*�dZm��ș�F�Vպ[�)
�6R�X�,�EgQ�;��Vi�x�֩ͧ"e'k��!����X��{3^�Y\��j+�
r�C ;15��DVf^��lF�jemF�,�5K%k�.����+�����o+hn�Ӓ�g�]�G��.�*�
MgjO�0��y�̭"Z'��n�d,�����&�0ἊR�֬�36/�N�:�FYȪ+p
q���#�RY��Z����M�ŭ�ZM�uz�i^�Wq�/h�Y��U+�+	۽{�J�ٶ�gC"f,���H�YXS�Wiѱ��J��B[ٻ���Ê�L�q�n��oo{6i)bW���ݍme5�B
�z�	7�*�(	��E�o�nP�|��8��Z��Ժ*ZV���0S�(˶x��گjV`�`����QN�s�Z�a�7��G�]H{��z��.m�r��Y�� �V7�J����ݚ�뻙;�a���A��`s,tCl5��C�囷ֻ����%mX�H� �iY$_k�� o,��i&=N���NG���l��;��E�	Cv��܌�۷N3�-�<���E��r���|�HH�XĢ4Y���ַ;��I��X9L�DNt�ܭj?#��yWv�a�=�Gy�'�br��5"�ޘ�}��hA5wR�1�9v��O#�+v�g\݊�_�e��*����9ݬ��MQ+$���%*��pZ4��N���(k$�Λ�B���n���L�.��w��Lsɑ�wxq��;�e��ԛ���uAJ�]�(� �%Ӯ�������µ3��ƕj�)��h���}�ul<^�|rt�m,�;��!X�:ep�;��5���ϲ�M�h<�e�{�:��@��܌d�f�Z��<��j��%ܣ���]̄�u�U�`�޼���V��:+��C�f`G�{ΕAht&�PZ�j�
��b�x(j�}��f��;�wv�1>�?(�n,sOl���)� TCq&c�2��
�N�f�w��������w׶�v�J ��}x]ڛ/NKo@V��YR�
��$=�sn��_Y�A��)��]w�>!2$���JR�\c�Ԧ]�l*��kN�u.���C����#��u�M�Y@���a ���X�*s^�hH��t���l�#�r��e��m��mͲ���M<�:�;ݹ�*Rq��e��%��@5��#/���V�>#�w�H�"Ҽ������3A�vfh��,^���]N��V�q��Bo�{�W���[b7�����['YC+I�)b#���a�,���K�t�,-��9]*���h'�v=�	 }z��XUY޺� ��׎�����1oM6�fϹ`�C"���G[�w�C����gq��&�b.]�ɥj���(���ol��U������b�o�!��Pڷ����0�V7�ymY�D�:��hӏ��o��+W��'���e �7t����r3د:�?):�U�Uxm����Xz����;Λ���vu����zDG��l-�q���,���ȴ�<������I�*�ŷ#ԣKJ�87՚�	.�7��'4���;�I��f�|��x��3���wyw����6��r�=`M�U�-T{����}�P8�T� ���t<��̻Ī�� Z����1:*
���b�je���%��*e�;F��}%�뻱�X�[�[`�h��̛i��ED��3O(I��X��_+7�������n�/UM
�:a\�kt�W+l\C�1�gV�i�t����i��η�K�M��Dk�ȢPh;��C2؎�W&jՆ�cyn�=1/8�|35d��<���V"D����MK,b.��wץ|���JUs�9���t�	�P���O3)�뽎�k���Fih���/-��tdZ�\������4��}�z\��>k:t�]�|�X�z�/i`�M-�^>|�����罩���ݕ+
׮u
����M�TtM�eu�(-7.u�`K�\�۰��F�r�]�IF�k����F�M�GY}�5XO��3����ywX}I+��u�o� �B	���Z�םg��W���^�[w%�1�F�ә�Q�#g��=�V�b7��G�8E։�o�4R�o�^^��
"�ћ\%#�=��Τ�q�3b��.�l�ӈi�^��$9�"fTv�<�������*����;�QV�Vfyi+����l�w�wGh��6A��Vǃ�97��3���*8�e��)���NX��L��7�`&�I)���u�>�� �����b���n�c���J�k5�dVc�c#�C�z��vf��Dt�����^��Z��I���T4*0{<�c溴pѳ��DO����9Rn��f�������}���E��̓��w��ӗ:zr[c^O����|��R��gc�x\��n�]P�Y��X�"umJUB��Ӫ��u\��5D7O��i��u�Bs֐M<g`��P��T*���L��4y���k�����1�_��v5��(�6mv�;�t�"�껷ĭ=����-��������K[uյʌ�u�j��NX{p�[����O1��f��U5��:�d�I�4�#v���"bK$wN�@�vv�v���2����KWjh�̗1��5M�����|I
,B�E{�4;�`��4[���O,��tn�	��;�Tr"�C����G��=!���T�Dv���^<�V�6������o����q�j�-0Q��l��|��(��^iv�n�]M��; L�#��y:c�@Eݜo��5t��Ăv�^�R�é�?�����
���!J,#�0+�q����Y���6�����o(ahJ��@}(�B�<|���QeL\�I2�.�����Q���u\��'1��jL��$���x�c^�b��X���c��t/jH���Ws8u7��:�X��c'i7��ݥ��Bk�}�	8Y���z��x�"sW�8��V���렚P��L3khU�������~8+T�[�}�o��Ў9��)?h|�O�/��˺wuH[�PU�Q���3|���#�jp����<��GWB�f
���E�h-wFf�ny��7��axs����v"t��u���eZc;��H'�S"��&nvވ~�Dc���qe��GI��aG�Z��-:�ɡ� 8�ǎ�B]���BG�.�	� t��h�Y',)s��0={	���\�M5�M����֒*���֪���^!p��C��{�5e��x�aJ)�̐Z���q������:B����~��[�2%�=�n��P�L�Ǵ���Z��Z�;]*e��k�?�h����b*�Z������'C�p_'b[|�c2���|�����j�4�Ҫ��R^U�+�X�Av�u�@�2;����X��l�6�;��R��)K\�|�ψy��b�"��PǱX;�-ҧm������a���h�=�6h>�ޣhZ��[�R/_Uº����a���S�!�Qc0'�4Z��t��:�<����ޘL���M�l���w�����E��u^��Q����q�#�_{��Y�D)|z�C'����6��{\D3��X����I�1�1>. 4�Hb4U��/Ͷ�u��(�>�޴�Q�u�Rkz.)�,�Nȥ��ޜ��r\�?v�<��ixf�N�޶��c�Z������@���*�	��%ct����%od�b�^����\��\��)�55��=j���v�V���u�e��f�W�kDq|��ү�>��bx�U���qJ�q��
q��Vwۧ�"�݊��'Q�95��)רM�;��)f�,�t H�K�,��t���c�;��k���H�z��y�&͋�_��t�O]=�UMY�U���8���}7�R3����"w6�7;b�V\��]���(j�Us,�XYT�aqe����|1���R;I;1�އ�3�����'b�j���t[/
ݸhʻ�1�0O}ݢL�"����^Wd�ż1��J�#ȑ�Hg&r'����]h�g��R�F��҉Ojl:u�5cd�ZM�DJm��]�m�p�t)��\9�-^qɗ��yv�x�b��-=��G<2Y�𴩉��~vn�l���`Z(�w�UvhwU��ۗ���L�S4'|��yZ��;ep�a*��b8��)Ļ�b�N��s��˱�ڱ`s��l�s̠u7���i�M��{% S��܄��t��!9/����B�=P+�So��������ڣ���>��2�s3"�rvZ.���o���]wëf� ���v���|�*�>ީc(�[`>`S�zO(P��30�3M�;L�����M�&��'.�T�1j;�:[�c��o��cm�{%��l��X#s�����s�u#�a&�
Bw"�F7�8o77m���e�Z%�S��h[9Y�Ȱ�S�˼/�0K��1�r��{�C2|C�z񭤅�]h5�t�+�^������h���mݔ��M�`Xu��iՂ��X�GS,h��K�nK�i��=����/�@��E�u�^wZm� ��N|�J���l뛦t�֋�C�=�[ ������,�Z36	�ҷUGݖ=������GǨ}Y�p�c���)��a�@���nr�S0�����N��go'�ך�W��R{�>�}o���eTP�Fyb�ԣ��Ov����{;Er�����aZd.��7b��`P�d�o��.�5�H�-3[/�5��F	+
����Ґƙ��a�;l^�!��y�i��"g�����{�ٸ[���Y	U0�whP�����ςx
�T?.U�"{A�ܸ��rW��H��woSg��6�V��eB.�=��b�|�4� �/�!����Y{����������*�Fp�vn��7���w��L��:�մ�����א�UN���/2U�D�fs�oy��'im� �<MQ{��T�Śt��{�敦ڦ�x�e�F^Oƃ���i�Xh�w ��JQq��1�h䤶5+F�QaH���"��.=9V��5�zO=�2��<-�Tt�CYh��zm�_���h�H7��Y	iN���ONʆ$�Z�6���<��\�8~�ު9-�yVm�C����۰�Z=�R̥,JEE�D�Fiɘޓu��{����݂�X̬FD*X�N��Ta4ft���gJ.0�nS�x�bp�=�����ot!��(r� �a��C����x��6�xux�,O|#Uv$�6�v�xdZ2�z��X�f��\\Z��]׍QF���� �_���C1iPrw?8�i���Z�.�w�@�X9	p����������p�X���R��j�n��S�-���/��/k&���{h`�6=}m���yK�V�o�!����hsjH��K���5��h,'���WmL�`R��,�WS>T^а;�0��W6%�|+�;@,ܵ�� �26�s�mcu8]gX��\�r�k�<{�^�;U��
��K|�Ǆ;�~w8���c}[/��0�cŉH����"�r%w;�0A`K�l��X$�J k�J�ō�;�2��r�9n#�T��������缃C�3���2Ꞷ��P��Ik�M`g��45�k���!���y�u�6�\�׎n��]=eI�;�����Ԫ�VF��;��𭹂�"�D��/t�-��ƶ.��R��E��N�"�J.�|��w��ȩ��+p�\�V(0j�y�ssZ���Op�'nٕ���}A{�)�/[ރ��G�;�O���	ܠ).�=,<��M!r/�u^���C*%�^�j5wx�3�Sr��ǌvU�o�K�����Py�����b"#p��>	�-�R�'�l1�]��x6�d�l�ׇ���ڋU�$��(u(MG��e2Y��e]���|�����U�u9��Ehb'�٠ot�h��b�(���=�R��_6�+���oM�jr��K�uZj�۰���>��AQ>�,�ժ�3q���X�-ζ)����
$�E�w�V#�G\�Ȥ����B���ˢ�Bu�s�Y.�uE��ֲ���0P��m6�� �v���\�B�+K���݊X��/4)�V�-�-�u:��1�-��P�I�$M:�r���v��p��ԝ�;f�> $f������Q[����}C��1m,;�ޮ��v��* ��x�����D��B��;1���q'��fv�S�=V��L|Y������k �z��ن��¡^k���Wj��Bv �����6	$f�Xu�VpçP[z)��.A	�.�M�,%Y�0�v;[�I`8"�-b������c�O�Yݩtj��y�|$��xٹ�Ҭ�/�T������C���Zh�4T��u�����ݖ��}�篻�[jf�{sW�UP4���0�E�-�o��-|�36���@��S)e�Ob�yæzz^�g��_�v4	1��"��G�_X	��;�n[	��++�+%�'hr��Wya��^ky���3����2�!P���B3׹fc ��(r")(�Z�݆�mh(�><�PS����0��ӦB)B�)�;�q���5/ᯢ�y:/��zFM>�K�<����)Jg�<�d1�EW>�:�ԅ�_vÞ��D,�j�8td�_j�%<�kx��J��ാ�@�K���S�&/x�U˱z)gk�z pe�6Tx�#�1�KdT�dXe�`�m�AJޝu�����������ޝ����b��}�v��&G�� ��7��є������������d;g�lE�V.i\gB'�o������w������d���8����V���:ֽKD����[x��KP�$��q�Ͱ�2l	]G{aQ�[�v���f&P;�&���hE݇�=ٝ���/��R����S"rV��[cq�wi9A��9͸�T[wr�����ʛ�;{�V�Lr0��]�qڴy�E��!��]ђ�۸�"�sW�Z�O8����W��C�ŗO-}˖J�a��A�NJ����^��j�������^�����͕����Y��vZ��K/�$3�Ri�(a���E����Ou΢�m��å����xu�N5u�[Z�滳�I��o��ߐ�2kBQ2�>r�$���COlr�=��Y so*�y�뫔=�ޘ� ϰg�[zzgi�.1�Jň�*�d���/1
X�e����	���ݻ{7S\�Jﯿ������/���������<�耨���*"���+�Ϧ/��ty���'5\�H�P�i;���W�r�m�����C'�*jk\c�s�fK�:Q|��-�t>���#��qM�����tk�פ֣��{<`1;�|�໤<���-��;2�r���\4�	�B�f]��XՃ9CT��]��{��}39�sv�<�t�y3�j݃tv�m#�;V|�8]��,��-��V����U.��0z�F���58W���6�ıJѦ!r:�`k�$��N����"�g��:2m��Ł�)ً�#���[׽�{ Q	ƺz��)Q�c%dZ1n���bǽR�ۙ��SA��o;��f�jhj7ȹ�Z��PSU¸K����Rͥ����[e�.���ID�Y�;B�E��/���ŵ�*�F�Ch���5
�����t�R*{����4.عAR�Ĕ���k�a��g��ɡ��=�x��h���U0s:s���Ø��LF��=��'�R�]%��*���+���Շ�՝�z����y�9��E�Yq�p��0��S���"R��f`"y�lfRU7ye�F�łq�K�۾{;7)��$�����H�pc�⢼�7��Q��ǃ�oh�x#�EM.��e�dZ�`Gz��"*Qh݌���%V�a�����%��Di!5f�7ez7�V>D]`��W��㷴-D��	ǀ�x��|�YS�baq�{��Ua+��>��[r���5@�����4ۼ ��6��Cg>Q�YF;z�T*�!��Q震������r�fh�#�z';�y��qX�r���F�S)����#@����5c��ӧ�d�d�l�7sd�M�7�����-��kڵx�o�]Vm�嫗H��:�#����Ϲ� ��P��V@1�Gs]�ß0��KG���4b���6�Ĉ(�lr��w`�'A���&�%cX5���se�)�<
M��,�h�S�
ܭN�>YN�0v����w��B�x�wr��(Y��f�SPMôy���Ó7fe��r|	�e��n��,y��=A�/�:��B0)(�K{2��\I,��w�AtK���~�Z`�\rKs�'\vƅY�Ց�6��z�bsI�R�[���U.�_Z�tN�[����˜����ê�̫g>�WWf�4Kل�6��e�{L��/*Q;���:6�Er⥜���%�q&��+ȼQm$�V&���X�-�R`��`���o`��z�Pz�O��7X���ͷJb�s]���`��[*�`&��ztgǋ�|�.�)��wEs������;�("!�t-Co����Mâ���''v �V�7��tEuλo`�ɶ5S$E�H��E�w3�.���\ts(3�l%IJ�;�$f��V��L���C8o]�a��L	�1��oU��/0�jnh�ʅqdn������yYA�;��3���c�缱m]hF3�PMm��M>�siV�GE-ɛ�����Y�/s�謲��h��=y�>{\���x�7e����r���*�Ǥ�|���wh��5��Ќ���v���_)���cl���j��}ƍ`���Fnѷ�ZS���횲���X7���]	� I�SrOhT֎B��S.�bSf;ǔ�{�6��X�V%k
[��0��8��\8stHsld�Of�,����s�iu$]�웎�5��+'��]U����*�<���Ws��iD-�b�N����#��g!���҆���A�M��WSw`�����{f�\v-մ��y�*.�A�Rp
T˶T�Ai���.���k֘(5X��.���ā��Q��2��tw�#71,��eI]I�F��S�i���W�˱�i���Ζ(Gqu�T36'iҡК�+<���sU���z�v���,���a���ʁ��O�)-��f
�Wϴ8��B�Ŕ��\����, �c�j�sty��AGG�փڸ�J���}1dcU�\L�c7s�7�,�d�f�y�@�f�d�g(�}��6�Q�ǖ�ݥW��i�2*��	|%��n�ɋ�("{��Dz��@�.��f����G�3؃����/:j����
V�\�V��Ǉ4������g�����<bhv��3dDm���RQ�	��n��m�kp�mi����Pm�v�U��vhT�Gq8�0M�v�X	DQ�ڟB��w3{k3n5_\��t��ApQ���%C��4�l�;���f�.�M��
fDj\$�B����yDq�|� $�P�/+h�u[�#�)w�I�*��O���,:+2��5��;��om�[�s�d�3��D�<70ږ�﫿zjm�S����"��z�2!�B�ǂoc��xG�\;���N��G�a��tJ��W��hGWq��	(�
�]l,�.�-m�,����ԺR�e����´�[�4�}�R������+) �K7{�8Cpk]�fu;5;����;��w �x���ٻ�B��Lɤ��@FU��=�c�%<���]O%�5Kr�ڷ����m�q;��J>���|���2�����ZE%�06j����ŋ��P�1�9vS�q;�m�5��H���hr{���)m�*��&J�Զ��CR��r�D{��_L��1�j�X2l(�G�g��t]CH��j,��Ys:��]$�va���'�˅h`�CÛ�����x%�}ky�eZ��_Z�x�t /�\�CP��v�
gDjz���Y5�lR���/�.��֝[$xM����<wT��J�Z�ǲii ��+M�q�y�YL!U��\y�2��`f�׈
�$�'�D����ł`)�,U�cWjhJ&��G!�Mծ!M�u:}ZL��׋����
�va��-b��;{�e���-�c�o冐��ja�Gh�3\9��f���K����X�
���*��d�7->%d��y�Ǫ���w9�U�� T�t�fj��J]Lv�]^�*�v6��:�4�V�3v���m�2�7��L3F'��{J��C�*���Ӵ&K���n�%�SYh��%��bv��\��\��S�R��)�ۧ���d� �W �Z�ջ���\{��>�qע���G���&�?v�-J��ju���%���O����7i]����]�na���A�oE�;��v�yV,5Fj\YkO���\L���샮�N	�����#;sK"�j��,����-�}m-���s��)�(%���WI+�J�w֨�i��z}x�n�� v���t�v��5A���Q � ��m7y]��X�>_m� .�Jwr���M�H��A����I�#@���� k#IJ�Vܵ(�YOXd>}�k3%��g�m�Ig%jx�����!ѣ��v�0̸z_K<�Q`ʾmM���u�Z�_{X�fs	B��\�>� ��b�J.e�݋5��]�Q9I^���I�V��;7��37���f�z{d���e�{m;��|�^޼m�֡�I���ڞm�4��qP�	Fb܈(7Ƴ���u^�n������>!���f�����[p@P'{,'�.���9�Y�ա}˸c=8�7�$^��Y;�EM�|�BC>��Mx�{�3Vu�rc쀯�h}��Wd���V�%>�ӏ��㯳���Ż��̥.Nc�Ph��0��ڠv����$A{o�/5��O	o`���vM��B�/���'ם!�]�<��<H����=)��˳��:��>�b�%�/WV�}_�_�݌b���+c�Z��1g�*D=�k�wa���W�$�]>�+X�J�������\ 5rW�����ـx���n>S)�r��6�f±���k��-��)��N�����w:�������8��'g�:�6=0��w����;!41З�^҆�B��m�o��\1Eh&��B��e��Z��T��,�g��:�T-�U�a"���w�KM�l٫�eʉj�����.>��C��A۹%�r��f�+OzO�>ۑ�YZ�[u�����g����}��[�\�Q.��R���L�']�7y\�a�n�n����M�*Z:�5�t���WX�7����u-��6Kۊ읂M��m.�`�|�$~:=s!�4�&�6��ȷv�Ik;mW$��1g9�Ϻ������yhne�1:�6��o	�ޫ	�zz9�o�⇆c؇�#�ۜ�3��]
U���mR=;m'f�����9��뻻4�����r��Nr��x� |M�{FeY�!�hޣ�b2��G4Yشm�3\#�
�������;}�m��J�6/�z�+��a�[1�������A��Y�<�@���+�.d0��|Ƿ/o�#(r���e���F�0��v��fG�L���w�")ܙ&iOP��KX���MwѠ���.����x�������j�X���;�k�	�*5��ܜ�]Mz���x���D���%����mY������U�;��l�����m�VSX`[�zb�R�ԓ0�������lL[E�<J;�[�
�i��n�{���Mhp��_��&�Ým�MA��q�ѱ-Z	��L�ﰦ�ـ�{4�Ɲ��D]w�t�h��	q�]ܯ���º���<0m�z�������Ў1λ��3�W���x��:^D�Eh��ׅ��|��=w?Gko=lB��`�hr)6_ʬ���z��각�!�Y���3*wW\�hL|���\q��,���o��@NT�10];�8/Z����#�r��\�9�dk��7m�З^��
4ms�jMȝ���3��$@�,�ŉ�_<�����_<�FV
b� f�Lѩy\�R��̀�&��J���ڏ��:l�GY(���Rku�N��	}��s1����L�`��i�̔�n��C�Ŧ��4g[/Ki��D����4�/\)9�L��KT��G�BGu�@�-���n��0��j��}:!���ms�n)`x��G�k.h�7*��������)�Ҭ!n{w�!L�C�jMQ!��e��k2Q���<���ft��W\�#�I��Z=ܻ�E�=.�V�������=O�OUv֣2Ź��z`9�ӱ��-Y���]H�O��¡�P�;���k��B���������"2��z4��M�K�c_qXZm��WC�C��kG\��ُ��!�h��+ LV$Y�=\���׹�}�՚�O}\kC�7Ԡ����q����Fud�E���<�;���!��h�yI��#:�@��
]��C or�ʂ����:"W n��%��V�5�/z3vo���8���Ǹ]D��J�C�ƶv4�홭�e�ҾC�^��
�
"��7*��!v��ݬnL��*���ٝ�-0_Cyv�J��Q��A��1Iܓ�j��N�Y��m�G�]*8�-���U����*�{.S/����yy�*­˔����GR�-�k��̭�k@C4T��<�MZ1;d �at�I[�u����\Nye�$3%k��K)�?��(���ׯX�k��p�{�w���^�EUo�=���gw�2K5�Fk�~�l��w����"s�#����M��j]K��udw�fS��N��ȩ��:pJ��c�ڽ�¥���6oV�lTw�P�k��$��#�<=�ۨ�8�N=��I���Ȱ8�H����#�Y:���]X.�X�wf��@��j�0��f�R�5���b��!]�|���`���r�#�0mz�;�]�Gۥo�*����nq��@�]#/J5/Z��]Hv+hY�}cC���Yl��v+j��1���<Ⱆhi����1F���X$��JEE�v���mV��[x��6lGژU�x�f3��E.=t�u��J��whp	��1d��w�v���Y��M�%Ճ�6㐱�:�}zr聨�}5-�7�<���|`Y��&�-m⺆�M�a�̰<(W�P�6P�/��>�����������]b^,��ǜ0�w�~��W�7�<�zp��0G)K�C��,�7C�J���x,c�;�-��d%XKs�x�& Z���in�ɝ֋�;����x�)�gw/wC�y)8��j��<��@�Hx��t�����0�支ST�³A�z��m�ʕzr��m!|ia�U��d<�B�r[�
ie�jr-"]DzI�(�w������ޥ8�Ihl�gD+&	҇�,Y�(E eʃ��f7}w	ۻr�.��7�����CR�uE��#8YOz�f26�tt03���n @f�p+n��0�_�̈�dU��`��������S7x���{��ipD.hSph4/��xĔ�rb��<c]P�h�&����-ͽ1��n�s���޼��2��P�kX�m����C[r���}��qL�#����R��߈ϸ�R�=H�7h)]֡4$;\��u�qR�I����9$lW�M��6��|��^�O��v��0�̊V��������� ":���GqA�N�����γC�6��TR���G&^+����ڞi�����N	\V�F,Q��Q{#U��`�nP�2��W���;�S�&�8d%fXڀ��;�C(�CoVe.��I���Gs�d}b���}K�gz:>N�9w�˦7��
n�(AR�h�
b���Q`@����	�b
�Z��*��6h���U��4%�=����ح�1d>s�q�n�L��E�F|�1���.>���d��U���MᛖS|/����n�re��B�FyF/W����@�\-�hǁ�g\����\���j�����PE�t��T���]٩.yx�^n%$[/�́::�;��`���e}�����gʮ���!�^g�b2�+&*�l;���H�[�E�]�|�i���D䥍TX}��2��d��
�o�	����s��`� �Z<��^��7��vp �ԻŪ{mN����U��|>�����ʔ±fmT�_���|�:�Z�yk�|ȝ�A��;笗p�(��#�F9j�;�h�v��ڜ�\�����ۣ�H����ls����wK��a�r{^����ϭBtG���˗+���]
��I��g��8�,��'w4({"kn���t��Z��v����q�Ge��=`��!�-�uts���XtliͻtOI!F�XZ(�ng�fg^wb��`���[�ބ�	 ��⇹�W=;���ml������{پ�f�����%$�����;�S��Y�J>�|��8:�]lb`|֢����>{A*Ǆ� ;�W�|�m��|m>P)L[����Ъ��NF�o�Ay{�VL{���##j%�;�������b�����������#t'7���g��d5� �޶�g$2�W;�
�P�OeGx/?��7eX�U�ٺ�j� �a#E�� �7��D�u���}oJVy�݃�;�@�]X�!-tԱ��0)ϧf!�i.;S�mh���Z��9�Vy!؋R�f�V-�̉$^ޭw���5��r��NNf��q�}w�u���ur*�ˢw��z�¥���ۺ��|ɰwx�R���4�!q�n�S���AW��}p[�!p��ws��7����Y,-������E$ӡ)hJ�O	�KHUQ�]V%���^A�(��O*M5�u�Е��N�ҥ�J��-h�rtP���t�K((JG �SCCE	H�SHR�Q�%:���1�G*]��F�m���[b��IZК��d4�!X�kJF��j4�Jh]-r�[h� �4!A@�F�\�R��&��O'����2n`�4��(h�h�@j���&���e�#��Fۑ�tE���9 ��L�+JP�AC���!h4��%]���Bi9���)��b�i��4�#���!ʴ8���b
�
V�������
8AHh)壛S�@U�F�M̦��na�A�4%ͮ���ʚR��\Ͱm���sPh9�����rB��{��
9e��@��w�K���;�:N�Z�jg����Ԕ��R�3��Y����Ǒ�G��}>�N5켮j��f��LrD��᪤۷fɮr���pt������ҕ�2c���]�������CL߼E_��2��)Z�������������0����I�0o|�u>nI�G���Q����@����*K?LE��[�~��ac6�u���A��ؖmrxW�ӫ�f�i��c��JAY��wJb� ��0D��/i��B��G{o����^���� �b��w������=�߬n\�rϕ�E��F��3>G�˖�b}�K>$v�_u+�J��q^𰬿���\��	��<�#ބm��G�"�佗eD$�1{�11���$!c�%�8��{���-�T [���{H��U�/h��7�S��tʨ�PY��_7�5 �Q��4ҥ�
򮽙u� m�_����c��8x^y,��w���R�v%o���V�>��Lh�j8f�� H�sΫ ���V�Y�}�W�e�J)>C<&�Y\�9�iυ/_ҧK�[�;�Ǩf��9_?H����_d�Mm��!�Po�q�{x։��fD.�\��'LKI!*���n]����Ft	����;���[�5���3(9�R�:����p�Pґ��  9�Y�Nb�Vw�H�"���&�Tӊ\�f��e�n,4]�f��X.��L��O�0Y5c��/���_��I/�l�:����G�O��E��{��iӻVWN����ǁ��ʚ�X�H��K^�N=�ok�ǵ<>^n��r���*Ǟ��n3پٶ~�}䶇g�B�R�dU�Z���Q�!5�Ӂ���E�+��^��N��v�� N�]�ڶ�P�>�0x���>�Ż�Zݣ�#���R!�z|�2��V���{7�����_oQ"~۩CA���,�(Q��b*�}�/�Ll:�9�o*
ֽ��}�)�d������F�%��ϓ@dƷHM6聦��>)�� ���?[��뾺�z��8�+4{tJ´�p\�9?bs�*	���N�f�	�r�_F�Q�#�t���6��I1ӓ��/��;�Qt4_x|-�d�z��:�!ƴ���� �4�ϱ�9~^5>d5/#t�9��nO�Z��^�j��倧J�x+�A��&���P�r�Ȇ���K��V�⤡�����|�Y��yȝW��e{�̟J�Ua՞��>��T���J�w�6ZÇ<]9Ae��A]� ��o�Ga��R���~?__�Wbw��=B���� ������^��-�w��-�mi�k�ۣA�:ʹ�l�gThg���<]��B�ĺ�S!�NJ���*6�5����Ӡ-�P�-�k��N�`�H���]�����݆��8�*�>}� e���m`~���Cq�?e�C��YuK�*���ׇ�"���x�r���=���7׶�K��0��Ex:�Gaʯ+��g�,o�h��9�J�K<����}��~{�h�!����c��HT@��S�[��Z �u�%Vyj���z�+a��O�{�}wu�j���
��g��]w��F{⟭���r��!9���腇���j5�X�q�MyX5S�����œ\<3��8;��B����iq��5�;/�[�I)��{8*u3�#Q�O�x����u��P߽=p	Wkx�:�\����]�/(.�[sgv�q����n)��[�!E�U��G����/Ƶ��εA�S���]ܧ�{o�Z����$��M�7�J���X�f�±Nvtaw0�Ք�$���u����*qлqZ�r�u���}����7\Cϸ�G_/�w)q����zy�Thׂ��`���*3a���l��6i]����<'�����K��yx��U��r�⼈�.��c@V����[W���l:�eG�9ޡ}NpN\a�L {K/p���ڳ�K�FI�<F�Ս��C�6Q�3H��+6���'��6:w��NmG�*�Y��A��o�82���{�j���p:c�Ȭ��e���譮�I�'�8c)ܓ{N��ɺ��\Ȱ��4��^��\-�k¼�i镋�/)B�w2�x�[�,�TgO�7�����MМ�X��j�������V����X���� �ր�^�~�&fu�u���H����d����9H�~^o2W]e�"��V(��Wx�k�T8[��'i��7�|\@� G���aV�И�߱O�������~Zc�Ŋ��,�,b� ��؂��1�伨��!�#x���^0b6)�z�ۍ#V%P�o�'�^7��z�������߇{m�5�^�pu?z�$
�K�E������ͥ�0:�����es��r�Im�s�F�D_�k�|2�!8�;�����"�5?��c�q�ִř;u.���j�o���z��X�䨳^�ؕ�ʶ����CE����'�������Ń�û��=�S����B��:�]��q��>�]}r����\K�|n�.��L(�}8���sȩLi�j��l⡨��{�sf�cB�{�ܟڮ��|�Ҫ��Q�V�Xn��Ra��*��yǺk.W�mS7�P�_7�j�]0-	��`y�{��CY���Ҥ��*����<�L�OZ�Nֺݥ�U�EdȎ6�ޔ���{�[}��ct'_�ƾ�z6�Ja,�u�Z앧A����,Ǌ�eas���]�6�c|bu�S�Y��7�u�i>߽�
a׭��C�KzMa�D��/Q-���!��p�7�k0�f�1���yxW�����.�(�0+1��l�}�0gAm=�5�^�U���?Qq�`�̊R�����j�zv�F6����xBO<.���{j'hك��Ւ1�}\Ո!����<<�dC���(���ݦ�df��5^Ð*�P��7R�a�)�V*�ۨw+$�-�J�R�z�?U�u���Z��`��C��ۋv��ߌ��}M.���wsg��<�P���_o�]<dg�יe���xl��^��Oۺ*�/s"�}��W?0)�� ;�ylg��J���'ޖ�&��w�Z�{�x��QN	)8Ӂ��D��0�fk�Y�ɖ�[��h��/i�qx]�旪d��/x������t�ҁX�R޻�L�D��z@!;�/%_�΋w�#UG�~Ƿ�SJ�Rn�}�/^=��PX��Ņe����pS�z/��������V�I^�On�
9�{&�be�bG���e]^S�q @D;e�&j+.x�H�K�YՋCNJ� �ۅ޵u��Ҹ#���B�]j.dU�:#�L�2,�p���F�u֦�����Z����2
+[������,9`1�;�Z�%j��%�u��W�F��Y��X>��pW���5�	���'^��vU�DGl]�1��R�Q�>�׫���e^����e���a�z"-է��P������>x[�6�:9y�*�w���[ԉ�v�'��t;�E�^oE���V�E�]���O�1���Ev#W�#�����Ӭ垯����01��ʝ��'����,���qk��+[�j�s��/vr�=c7��^�p�2�E��۹��Bk,�w��O��k�d�z����;�{�\����ݩv㍪�� LER�UZ�1?ENn/�{K����eKv�۷�ԉ�"���^�١w���a�%�w��ы{ 늴|;v�`�זa�:<5ϕ���}�9_S~�tM�3-��U~t���5~�ss=«[�u���CM�Y��#Q�z�v�pk�[{���r�Q��rEF�����ƍEV{�Z��LH��s�6�o��[�F��3���9N� �>�`(�u<����7��y�X�^vG��1B�{�����V�5:��������
�
��ް��4�I�Ξ���Y}����nI�1�m־��q�KB�Ì�O<�F���U`����R��L�C�"��ns��w"�Y�:�"	6l|j��m�5�2�����{Yf�q�Y𒭦I}WӺ���y�jǭ:�a�=^|�|O���͏�=�]�ȁ:d��P-��Mf'�wsA3���H�}+KPb5�c�0�[�S'��CΝWy4��W5@X�J<{��ro��0�C�yթ7���Wf�}j���,8Q��1Q�#L2^A����u;+��[�-Ŝ5�06�~���R�X��L;&���QbƳjր ���ɹ�8v��-����f�vt,5�F~֢���S˸����Z4�b�*x�㺣�u� 8:����aָ�P���kH�^�����b�{�#,�w�x4Z6#��*�VW��9�d�x��e�N�؃�i����������d��� �������t�Į�i���	��}��D��U��}u�
�_b��{W�R��u~����4�G	�N�E�s̽I�E��R�\(��>%]��Cm�̮��&;�i�'�v�ދ��;|:撚;�&N�����ޏ}����|�sU]�_�Azz����
�篏��j[���y�4���,��wlH0���Of���`ݸ�G�go�q0��xa`��o��d���֮p͈�u�����	坝�K$�ȓ^�=j��k�J$JZ.vp���w�'�ҝ]u����J�6�f_0P�f���݉�R���\��Www$�1g��^���|�=E�Iq��Է��6��y��;�%1+b|z���.�j?K��j��w������<2�2����y#]<��m���X�M84.)�S}n��VP���^��u�����˛'�K;�K٧إ;(,;��b�����Axw�{u)ņ����?l�a�hW_'N#�e{k�E2��wnk߶��f���=1#~��J��l�w�Jߤ�����fog�^h�\��q��>��KEa�D�;f�s��e�\,x}�u���G�o����ҳ�}i
�̮�w��q���c��&��.�
%��믈ȭ+��1èo�1�=�� 1y��ےu?p���61C |�����ug�+D����L�?*�V6�g6��`�� 3G���«��$|f�!�̰�4�Ш}�?��<_��گ�'�8=*ռ[���&c�m�ø$���b9ڍ��d�4��y3�]�pJ�ՈՉC�4_�?�3��tR͛�Y�"��f��Da`(٘�3%�g"�^Ǥ#���e:]y*������,t����2�^tý>�E0��AzN��~�:5.$ē:�7v�꟟<�ī7�D�W�p�<Ő�[��vӡ�KY���u�Q<�\O��օU��AM�|�)xn�Gp�{]> uu��]�Z��
������â��0�������M| __(<*q���{�]�:9wOkV���ھ����а��z�{�n�F�����wD����ʿ +�$8\�8���>�%.�V}N�Bz��=S��Y�W�����/o��yϩW_\�	�ļ7��ԸV�X@�&�k��m-v�,5~����O{��_؀\��f�O�*�B����\���W��uz�d(�~�k�aT��N2�nTf����2�kLD�LM��#N��`S�X�U�1��T��Z��=�<�������Q�`�}'3�C���ῠ{LxLSLC�M
�-Èylk�͏�~��iSn7N�b��'��o�]�He�]�Q���EK��5ߥ���.Rvqo�yo����i����G���P��2vݟ����:
K�xy��0�8|+���:��4�53��pN_�ǌ����� ��ʫ�{����(s;�9L1wAF�Q��W�m�sI�0�.wt����3 d�k��F��\5׊�|r�23��,��c�{3�c�hJ�e	��V�3 ���5ul��J��x��/�=E��[a��g�q����D�SDi��X�M+�s,�e�a��F�wWKI$D֨�1���q��{ ������N	1M��U�ff�Yz-t�{s����/�,�_�AN�e���.�	�7{z"N��6Yai#�}�ho������$ɘր�ik�"~� ��&��G��7>~�����h:H��u���~!۵��YXtaI����0��fcre�a܁02LF0^x��]y��#}Ÿ��r6�T2�}t�~�aL\����Em���eYS�j�&�0�Z� M��Q9�� ;t{��,u�C,�m
˫��E�.V���LnL��V��f`�y����~�\o-V~�� �d9�c�{���-������,��j�����;ug����;��\l����9�5�MG��J��.ؙ�˥����x:�:�pC�W���E�6^�x�{(	f4t1�i��D��z%{1��UrV,�I�>�˧�O!�ٲ�y.3u�}�U}�j^Hn����VI��T1:k^��c�r޺cE��g
�pУ��U�w���g�Z��3�wν�c��H�*"���P��WT�0�$�A�mwEM��Z�ݿ�& �mՀ�|T��q�P��3{_�9{N  ���'l!cMY���-�-ǟh�L;g2�a�a����6��A����/���p2�9m��;�L�R嚕�Q�r�.���E�A����ox�:��%��˳��,�!�Z";��_P�M��,핱�7�h�&ڭ�ؼ+�7��h�k}tT��y��ln�^��weڭIb�4oa;���̓T���F5�vv��trxW���У\���T�&AT�ן2$�av+n��n����v�Gn����:-�汉K��U����3��>�� ,�pmoJ�;8�[���s�YoL��
���ĝ����t��6����Mi�\^� =b�-<U4�hk�\u� ���`����lGݮT�s�Mu�{1`A�XQM��ݭ�'L��Q!H�N	���n5�`'oS��u}��:���R=u��<|�����խ���<��P�;��#���y�c��voS��P�`-�5�n�NF3���]ʇ�x*�Г�K.�$eD2w �F&S<�������f�T�[��7Bx��C�����|7}����;*���H�g ;[0éix3g�ogN��֫LŠ�(��@�F�n9�E�AW\�L2I��
��2B�{[}��ʹ+���t�����^=K���j�a��.�[���C(ū<Ҏ�J���≆xƣĸC��㾕z�B#:�c�QxL��T�1�۪�(�JpSʜ����t���CaE�mو�#v��b�΁NVfr�7�$�i���paM�%�N�[����u���V�v���tu���(�406��%�<�K|�:�WN�غ��S���f�v�>3)�����g�
A4���M8�v���Lv�>�m�/��M��-za�=tO}��^1��
���{Zu�Mի��-�ӝ�����˗�j�(�8K�)�r���s�I�5�|M�>�:��+�p&��:��J�m=Q��݋<X#��{�͑hw9`Sv�&�f�T�����fF4N��_&7�'��h����y�x.U�P/E�O����u:.���&��V���9w�D[���4̿³Y֯�W��7n�ݔv�5lbZ��YB�B�P$ }���m��* ��.���#z��9cz��KY�;:�o�i�h��vD�}��wK^^s;�N�4y���8��BEi��#��K���b��i��k����K]�άz��v<��uqH�=�k�v:ݳ������*N�/R9��U��N��B�l��{2[�I7`r��������&`=5�6榆�7�Ȃ�������A�m�V
�L���;���z.�A��}�W;I\���k`����P�e�<�8vՑ���K�xto5'����\>�M�^?`��e�×�,L�Z)�*��2�uAZ�&)�91Լ[��0�t;s�K���usJ>�
&�[�v;o6MA��1ƭ]��RٹK6����M�
��'mh
�SEKy֪�h�g��+O��e�M3�4[�(��-�j����U��R��V���h���kȔU�ק�q���O�&�
�dt�K˕R�-4	DZB��̦�@ii���(^G"��w,<���%%Js`y��EQKs#��
	��)t<�A�R ������:�!ZJ(��S�nA�B���4�<�� S�5h4�:ѣJi��i(1:s8�I��r@�<�s�h6�\��5HLRG1A�)
�hֹ"��Ri�i(�t�4i(J��PеˑJ���%4$ѡ"hNF�@�.��(4e�����4����((b]!��ևBr<�xKʎKO �Cl&�5�]-ht�iB�ѤM��$҅�
@�(�]:i4i�;m:Cl4 ���:�����������\!¬c}S�F4���/#5u�"�ss]E���l'Y��Y��w��Kfr�����u�]���7Y�[���~��J���8����{}���Zc�}?�p��i־=p�A�F���|����M;>p:��7�?���wS��h��|=���?��w'GrLV��UvM��Y�]"�b#�ʇ��q���������sԺ{}����	O���8�F�˕�}�
�+�O#�u|����C_c���������9��s�OP~����w@ G�>"��On�c�8��K���FA�%���:����y/|��P��G/��?���F�e�v{��@wPi;<�]&��!�4��{�A�r�C|��M/PPy�~?z��!O����p������p��rĤ�\o��Jq#�I��#���̇'�~ܟ߳�h��?G��?�i��s�0� ��N_<���˧O���އ�����\z��:=>u�����=��^�b8B�Ж��Tb�-ʯ�ػ�ܽOӥ�F�G#�\��?`��`��=6^A�:�o�{���$��{��������g��w����ǻ��C���޻����" �"2��R��w�G)͇��Aܚw8u ?F���>���?����`�~���P���v���NC��/���A�;��������eѡ��C���t � B{ۢ�j�Xh�l{݀���ν9	Z�/O߿�t;����l�A�����|>G�J����޹A�>��J�� �߹y��#�A��Pw�h#I��k��Az~��HL��A�|�@�N�����N�|����W
�)>���1��
#{�����)���<�����N���w<�'��?����!)��.~��>�p�O����?`���^I�!�	��D1}����:��Z�Y�uع�b�������:g�|�]G����t�I�9>y�}�O�t�>���R��R�9��Gp�5俣�ׯ�C�>ï��ܝ�c�%>��9�/W��B�������9�￼�����}령 >�#�>C�~�C�h>�� �F��c�Os���~y��=�Py&�����w�5�z��j���}�|���:�e����GP}�~�>{��y���~v�(ww�m
���ӕmL�u�)vk�ֱ��\/\�5�1���8���Cj�?���µ�s�fx��{*������ad�mh���ٽHc��=��]3���я&9h����0g	�0�2S���*T��ziP�9�Wӎ�g��o��2�����j�r����ԏ��Z�'����	=���=?c���n�+�{/#C��O��y	^����#�%h뗓���Q����Hs��������t��%/���G���=����4�{ }�}��o�;�ɍ�I�~O�}���������M/�:���^A�y9��k�r�?O����~�������NOg�|��O%���_���}��yKsuW��	���!@��!�g����|�O��|=�������Ͻ��~��Ə�ru=A�:N�n�� ��{'��;��:#�������t��ǳ�;�%����}���Q�~�2��ј�����A>���ݟ|�h>C�7�/^�J_ϸ(�^�#�����A�$C�y^�	_`+G=���r}����K�>|�I�&�~��PƼ���&=����%{�A��Y�=�H�,�����A����y���<��w����;��4�s�/\�r#�s�N��˨�z���.��*������o?p�>�P���.��=��:��w?O�1�L�z��{�G�,��#����p~�p���g�?��K���^I����y���@Q�?`���~u� <�=�ׯx�� 4>Gg�p�M&��!�M��G/������]W�x����=�h��zV�B7L}}���O ��]|�r}������?��;���>X�w����y��4?�h��� ��� ����'��Kߟ{��|���F�{�KOPy���j�t���/gc3�Mw�DX��D�G�]�4���8w=˯�0w>Gq�/ۓ��h|�^������a����K��:���ǒ��^^GPx{��P�u��:~BWPw�/�n���Q�y��s/�3�Dh�DA��Yu��?�䞾��N��<�'������{�A�NT��ϙ<���~��I�#A����C�����z�Hr~����?�n�ᩥ�WE!�|�/a��F�8Έ#�}�C�����	BW�;�yGp����|Mw�G%�u�;��/����u�΃����w�'�������M{=A�:��4? ����/QU�>�}����<�v0T�k�2�ul:����;9����Mj˻_\Ϩ��݀!5�Qǻ5j����@s���9f��|ndG$0�6�ou�K5b1�-�^eN�M5��+��w,�_0i%�$s��W������~��4���/���}��{���ϼC���:�κcs	�O:����?���:�����O�Q�;��?G�J|���}����9/g���DW�Un/]���;�no�g���G�߸}�����}��~�C���.�S�;�}�{��}�^���z^����縣��)�N��xw''��y/�Ӿ��
`���}�;�n��U�9O_i��c}�����~�/���H{���.�/.����wJ�@��)��4"�]�
����X��8.�c:�z�\z{}Kѣɉ���Vϭ@��~X8��T��򡇯˾��#���(Ys��&Y���]�d'á
U/ *� �'g�r�0��=(?VN�F�D�㻷���k0���7r-���N�{v �ە���!~Ucey�0�sH2g�_��.Vg���m�E���e\^��ȿ���9��F��G����̾TCw<�Ժ��9TH�4KͷRQ𻹦�xj�Λq�dC���}(&m�yÝ��#T~��ź��5b������#���آ�,gU���������9�P�a������Z/��p��܁&r�X�� j���[q�����AP�W��1�(��M�</�.y�C ��uធXk���z���ݎ�bRN����݁]����x��[X����h_-��z�2.�qŜgxNZ6�8}�� as�F�Iuc�dX=1#���yi��]Ԗ��m�ßW��&�z��̗�b�X���;u̝�բ�j�V�y@M� ���+��{kg�Gy�Y+ͱ"��6,�����<U�:%x10�`�,�� xT2�N�}��z��c��k�+n��uj��묑��5b	������*~ϭ\��qh��ie�v#��kL�����L�۸"h�1P�)V��X���]�[�xI�p���dj�l�O�gv�M��1(l?)�@�����1�����!�o����M�yLRں����(�ƹ�3�����V����P�_�P��f���t�r���� �5�U�g��J�ߗ�┛A�:V��{����z�B���)O�?}�'��4�z��o7�繀�����!�6�K<�Oq�'W���Y9R^�{�,��c�?��N� ��W��R�^^]Ⅰc�sW������bx+�݄�fR?h���J�����b²��xQx�����sn�B�T���[�w�yb�%>=����Z��F60/�dt�{��^:����ʡ��~ Q�W�����Ք��u��pg���~3kо�a��Q����-
�j��l�����r��КzfJ�;���=O��ԇע��X�m�:��f	g�3��Ya�Z���֧f`��ʧ��;{
XS��:��!^��gvv=��;w�Ṁ"�ĻWzc}��Vv�Sn�������e������1�(´�=a��5vm�F`�;~��z�vslP2���F��rƣA���������H��y�Q/�hP8���{�Y�YV7/�ˁ��o�`1���P׷�V;�/4{yk;9W��6��R�G�.�F����p�]�<�w^o��Y�(����{�O�M<%ZQ��y}�>�&�mn|��i��.Q�j�+�q*{���֕Y�=^����� ��� �[⥮�Oꅏq����Y����5�Y��������Ɛ��w/�]}Q~�,���&P��7�Ɍjy�4���9�3�����8r�G����.Z��(xPZhkMLn}↘�9c��F���wg��ȫ�Qp�d�P����{�ck���ٲC��PcIPg�B���o=N\�-n.1����;�WV���b��!U4��=�����r�����hd�t@j�;OI��~�m=7�y���鼛��B ����:ۯ�!^Z=O�@��br�z��"�6) 0m�o=�)l�u�Y�� DX��Z���Ghp������2x=CΝw���e�7�~�Ð(l� c��C6�n˰�^Pg,�����[�m��h���hh��biT5R���춷�ط�O���T�A�u�U��1\�}ع0k�c� ,��n�v�;JggYŅ�6r������8�/� �uY��^d/B�㗃��a���˺�p߳|=% �����Gܵ&��j��u����X
j�0�5JI7�Tk(�;��y�t��HeS�߄���b�7� 8j��{U��Y�n�����+�6E`��
�8����� 8L`i�γB�w�@��e�5�fsƅϯ�n���_Y��Я��k$%¸曎��EW[�y��x�9�
�+�
�����v���+v��Q�Yhﰭp���^���ڥ,rw�@��iO������1ڑ,�>����e����=UdMN�;�f�R��[�s͑3��D����=ڐ�u��>�<�}�Sٌƥ�)��`�b����Ε�)�á�N��`>��X�iWO��;N
@�[�\�J`�܍����Y�K�9����0r���\��j��k��'�\\[���`?KG.�k�v�sN\���}�e���4N�ʀ� ���_k��j���!w�GG1S��^P�&6s=O+��iE�l�H!�^�S�b~�[Z,��Cj�t� f�A� ��̎��-�R�f���l����n��kƻ�ɇ!ú�T���9�y%�m���� ���^S��������8����e��D�5�N��yR�=�F���H�4P�L�3coBT�W�1�`uq��162����\���.ﱋ�{�u�/5�M�n�zw�Sֲ�����h�5�0h�j��(�m:�G@����z7DF=�xZ����q�]�C���g���*�V�2�������$�;B:(��o�=�5m*�{��aw�KEd��������/���5�^l��l��P���Vz_+P�k���6}C��]�.��t�b��{.�^�������'X�X�<�hzo��+[�qW#p<!�j]F)�فGގ�����Ԯ�U�M�)`z�.��8����̛�n�\�� ^(�fT�Q�fC C
!��鹡M���cPc�;�^�1��ByL��JT�?a2��"V}�G�N����^�g2�|׌�(X�޷�n4�XquNj�|l�F�z��l��tx��V7���
��
^u?z�d�j�d���}/�"��:�f�V�F��UfC�G�N�"/v�AO9��!�''w���M| \X��l�GEmJw��^��o&��[������Pf��0�� �%~3������o�d�u0��ҭ����h���u�*V��`�V���.�^������\�"�O}�[�E=�wA�4�>��QV��&�9!>����7;��pH/�.F� �ք��.K���P��5�řKr�9]o��tO5%�����@6�mɷ ����w#���TA���b~<6�̾R�q��>����x�����qf��/_I���
��
u��{�k/���+�l��̊��{�'�v��ŀu�[��xɭ'�'1��yP�6Vᯄ�^���mm�c,�:#2����]v�}�|&�ۄ�	.��n��u�T�QL�J01Gt�|bCs[y�/���b�P��ه�87D��G����v�9�f�c�r��2�s�y��ϭ�}������v}���"��:Z8��(��3q�w�d;z�V��S�U�y�4��}����m�y��΂�������gr��+�"�7��q��]{�[��}w�G�P�"eR��Cܬ�7حѫګ��v@�	<�2>c��.�7����^�����<�(���2c]�
~�t���h��f�>�<�Ѯ��ES�0{yd����a���$���#nܩ;m��,��F�������O��.�M8������"��T�i�M�Ugm�����|~�J����2ø�>z�S��!:��'h���)a�R鐾� |X����΁>�cw�I��~k��i�;�ۡ�k�E��uw��ۗ����|����|��B�D�^��^���m�#-r�s��ĻĆ��%�\�9���}�jr���ZݚȒ���f������y�yo��0�~|a��X�e�f�Y�²��N� ��z���6�Zh˖a�����lT�9�ҵU9������w�WG���`�Z�k5�?���B³||(�.V�����o�x,g�5�hr\*�׽ \Ez��t~iV~�o��І�1����x���뻧WP�NZ��H`C���7�_ڟ�m{ݪ�
���;�� �"g���X�E|l=�u+�7y�Uݦ�ch�A\��.\��
3Th3t1zk�֌-�z8Q��j��u����a��k��wu�~����7��;�/^�.HO�x:���[�)x���QБ�ɠ�%�����T�Y<+nϽ`<-P�W�E���7���0k<m��ѦV�F{��r�/R����ÿ\���D����k��L���o���kH��:oօ`���p>Ҟ�wXe���H�ӧp����k禾%�wQ�R2�d�n�R9R����5���d꺋��0��V+��E��u!1�Z�ׅ5b�z�W�b�?e� i���6�Ǟ�B8��:�7/�`H^��>�mFN�A��E.��W�K�x�SO}_�]CDէ��Q�����x���)Sҙ�1u�w�Zi�n��<�~��Z'�W���J�5П[6�2e���s�ʰ�U�<�8*(y��\X�s��]�꯾�y.�����-����ۭ�Wx�����z�O�.H���36�����`�%H�����*w�F{;۾�RҤ*���N?m`Y�}�ː2��~�)�5�Z���Ӈ��}�PϹG�j�0M2���qR��{G��3�\.�U}ҏ���Xј�$�4{��\u��1� ?��kC)X�����Z�t8X�u����:��/�O��9�ϲ<Ul��ڊ�_g��d�t%���#�P���UK5�k�s�倧J�xkC�f	�_���ѡ�ԍ��q�#�����W���[S��}�טUX�?�_Gg�C{��[�z����Ǣ����q��
Ӣq(`=��x���}�P{�Ke 6���7�{姝e{��U�}d�uG������gƣ�"ٟ�3d�D���Y⾚B�yu崌�Wஓ�k�Л���bǫZ":�s
�if���0Ӭ5ẙT�]�_�;BM?W�QϝR���1�J}�2�Ѻ\=�Z�E�E��n�B|r�/i�ԅc���ڸ+��,w�M�i0VM>�D�'��C��:�te�M{�]=�p�M�Ń��^8�V�����Vz3��`�;5��ff�?DrMly���PfҠ��vW%KX�������Kp�M(�c�|0u��%L�ܝ����
�ֺ��-���Q��Rm��T^���������l��-�XB
�^R��r�].*���32�Մ��l��v�`u�;�����E�K3V>�����8��37�n���2�#g4�T|񑳵���z�nEj���ȯ9֡w����]V�c�����ِrK(u�w�v�J��i�� "﹝��m<ʵe���ܕұ�h��p�=j[�{�f��)`�����ku�.�Ih�=R!�Ν�F;U��bA�Qp�1�TޡWd����J��:z�6�#�>]�̽S�
�.3j�����
a!����g���b"��}ʶ�Z�k�{O��}
����Ȋ�PT۬�Q���s�׀[�ErL��y���G�0�O�Q�u�:��,Sq4��Q��z�n�Փo%��cT��@��ܧ�Z�C
�W'�O)�!L�{����jt�粳_[�V��Yi]%y��sz����LY5GBߞ��f8�d�W{E�;�B�Wu𣐪5p$ީx_H{1ݼ�K$�u��UoU٣H���x��)j�>��y��f��9�1;�L��` r�2\� ������*^�LK���Zݦܭ�B���׉��q��s����(�w��V�0Q4�dH2��vuZ�Ɗ&��3�yc��,�9��c����#�+��7�&_SЭ,�e��\[I�Q�wK�|�P'Fn�j�f�/����լ4�ѵlz���dW������ޢzxr��wz:{<5z�3G/�/��>/��u Ж����.�y�������oiڴL���)��N�5gm�QmK�gD��̞s���L71m�P�k}������Ҥ���G1�'�k%�7�X�ֈb��r����.���D��/$Wc4��$̦d�Y�#z��"0%�.?::b��.N+s�T�UŦ:��O�Z�pǗ�����8��n���0�O(�+`��zX��,�(+x�zh�΋|ձ�jTC��!�I���}˽˥B��@���Uwx���1]&H���L�9o6���-%G�䛳o��P��K4��r�ѬZ�[�f�6(o&:66fl_��%s�=��}���*����ٸ��e�T�c:>��-&f�]?�ʶY�X��JP9.�T���/E�Y�.Z�R��^��.�
�f��5�D�b����b���ȱ�{3	�J\SdW+�t�|9)ÿ^d�G�7��LS�A�FMj��0{�o������B�Z3�[g�S��W�o4�FN�)�� ���#F�g�9�ݗ�5nL�*�!��oZH5;~��ՅvJe���N
vs��°���3\���C����ۍ2�O�ڜ�X��=�ۙ��ˀ��uq�;�����C_h����W�}���H�����KV)M/!4%)�CN�Jѡ4�ۗ:Ё���F�\��!�Br
C�9<�e9'F�R���69�V��:Jt0�'�IX�٤�+\���A��9:��bi�l�ѧQ�4Ӥ4:�5N*k͖�M��q)G.IAB���j�M:E��d���GZ�C�RUh)КM6�iB���9��Ƞ�K��BV��A�.�M�h"]�(�N�J҆�M)�B�1�NAɠ)��9���ST.��:J*�+[gIKEC�����W�}��^s�ݰ���xZԺ�=�V��rgoQ&3����S�zJ�,5�X��i���Z����F�X�B���R�D}��[^�yz���/sW򂜫=�Ο��J�:�S�)^��}o��*Ү%�}�������ݿV�3��<إ��f���b�xh�hj��]�)�5U٫�A{с�=�/�+-�*�:k��{���Ѿ�-��mK�jc=p�`�70¬�v�����s�mw�(z)��rI݆h*�]iS�^�R��V/<�u�E{��P_�y,TsmY@f��ݝ��GG��y<z���&$=썊~^v*P��Bu��>�C�hΧ�;��Jqa�(d�u�(]�*��n�(1NfǫU*���KGe�`^��@-��WLƇ��-T�ղΫ��20L��:!�Aϳpl�4}lku4D���*^���!s�������*[�K{�ƙ�#�;G�E����N��6����b�I����z�$tp�"��u��<4�{^��~r�ads�-��`
5��2)��$�{V7y+��OI���ť���.���hwZj�m���&S�f`00���ƛ��x��{����5��ۢ�#P���ՙ��E'=�d��^����鶡�������P*�:u6��\������nMtH>�q}rzj/��rw��QV��_����8��-�T�z7�8�f�ޯyg�Y؆8A�<z���L�;:_fc��DŮ�6� �-��|�j�=9Tџ��W�D�����K_����<Z�9UtUA\"q��^��R�w���XR��xS��z;;˶���}-$j
�����弟zZ�ٕ|�yJ�~����L�=���bN��O+�{~��co7cs�v.NQ���Dz�-@E�k�"�s�CHe_ /����J��
�.�^�;�73}6I}QwQ�4'vq�m1!ބ��1B2~s0p�ݤ�l����kX�>����
��=Jh����#�?U;�Qt���;=}��(h�ʠ�vW���u��s���Dq�N��H�HyhU�����bZ"b=�D��f�����b�����~����g�j�bMԘ��f�[���]�n�ў�DPY�� ��5���T,C��V��T��l����f�o?�������-`n]zF2|W�h��=�a�=�7MTf�7�,s}s�淚�N��2]���U�jxN����:��u��ر�?#��ߎ{�)��u�ѕr����H�C�4�~��z�͠2iK1�F6���f���`��A]���UUqB��-����ؿC���;��EDWh�.im�{��O������x}���T�Vm�ӡ+F�VgK3�B��u����-Ecŭ�S@^b�����}�]��T*AI�l]�2 \��zfh��ΟpO_�2�6^(gP(9���ﾈ�����B׎=������,tB#9���v�t���m�^�[b��x�J���/�Xڎ���^�V_w�(��i���8j� �������u TAB7X���k��^�����-�\�p��ǱN��~��a=���?[e�ِeZi:�%1/)pJ˲��E׍֛����0%�n&�	�ފ�#��T{Iz5Lz�څ���^c��	�U�rw��J�֔u�n{(���N>�`�����@���?#A.�p���)p!�� XX��&/�ڳDMBY�~sp��[�"��ϼ���	E~xaÕ��A��ܿ
1��A\�nk�ٶvm#�,3{>�ٌ0�UW=3����^����/M�m�V]M^`ef�t��;�{t:S��qb�8��)i�;d�\��^�<����H��Lv|������v�-c�����8�����GV59p�`֊e���%���p�)8��ϩԸ/nB)L�pT6�����""9�3r
6���2��;�OF�H��ԃ�#�{��/vA������X}�ؽ_�8�J�w��J�X���d"�o�:k���:��x���F�r{��">Y�-��t�]P[4󺱜oٜ��}-���֜5u*M�Q��b����z�[��
�Lv�:/�A����c�;Q��a7t>+����,�3�k&�0��Gv�n��VL鼸��q��X]��,�:Kmj�';'v5�u��}V'��A[�Vv�y�����`�7�%���@l>���OMJY�^�:��Ȍ��u�����͛�Ͻt��v2�3�f�6{)0������e�/�F�̠˙��/�e�T'�O����q�^��l��~���~��ü��g�m�=/��L9�X=~|EU��qC�k�_{o�;��"�����>��;��igѹ[�6x�U�]5���)��t]P�g�AI���7i��ڷ_q�:���o����d���d� ;����9�K-�R�Kq��U����H�͡1�VN�<�j�?Cǌ��� ��[������4��m���o�M���ly���{um��8h��zTs.�S�� �YrR��8F:�y�:�������aҬ/��v�=�u���,����W�Us��\^�B�Y��~������`�NT\�唱}N�k���E�J�yI��=�����r�bc����8��[�uz/�}�<�q�Oy	y>�rƧ���������s�9�~�Ѕꇈ���f�~ᇋ~�:=�`�A����1V����Nw�S��2Ѳӷ��]����o��<�=�I��Ϣ�w��^��2��҂W��%�7�|�z÷܎9S���_���S<�H-����@\�u���̖�-��We郩��cO����4~��`��2����΍���V��cӠv�m{:V�s�g"0��;ɑ��H���R�$f�3��6Y~�Ǭ�g�Ve'��X�����O���:o����,^k�o_�vu�3Bj�Du�A5�iٓ��}��y�m�L�=�Fn�4��X�sI���*S3w��h�Z���+iڽ�1�0}�{���{^�^� �^�j]3ui�i�㷹Y��`%��{�x���Ea>�g��O�)�3KQ	<.��id�M��׏	J���l�_H�]�}�y7<�>�m8��������G3���s����*˿Sό��m��q�������;���X���ϧ@t��˸�n_\\���_j��g]���!(��%/w�݆��fV��N��<�_c�s���P��'P��6�LP����=�CWz�iW��qy;"^��~�މ���7�xʦ�۱�s������������N\ްV�A\��,=����/xK5����{=�8��ﯪ��K堥��Ծ�Յ�z�9�p=���d��QߎQ#GԷ+��!ߍ���D�ᰩ�{�L�[O;�p���z�Bf��)�<�6e"�5�7}���3���u *��U%n��-�>�����k5���M�e�ի�1����ʽ�W��^,g�:\u.��}[]�(lt�����k�G9�Y�	��L��<d�:4hIi�H��=ۧ��,{v?P���|������X�{+ml�knL��u�.֮(x�a%���u��܁�9���~��{�G�Yy���Ӵ�'�F��XEx��Ǩ$�}��<o�oU7Zo"��J�o���W�U}_�K]�Xw��`��p�9N��F񰷟-��T�͗�:�p�:r+���Z�^���g�z~���(�o�ar[�k��,{*�{K����ƻ�tq׎��r�p|ˣ�x��r>#l��zYR�^%t��,΃o\����C-Շ	���4�Q���&�TN�L�g۵��
�C��籚���:��iЋ���a�����=uO*)s��3-�]��5���Y�ק~;�6�:�f.�x��A*�׺�Î]�l �c��>�_y��0��~�J1�8���a���u���v�En��|({��@��<���L��k��ָ{�IG�:����tg��u	��F~�yd��U[WMת�)\��yB�����>vr�і.ۺr~z�cK�$�F8˖���9��5��a�-��4��%&�������U8C�fHk>�Q>9z7����E� +���ZMvL;�`�н=��o��3�wy���g:��W>�p��{e�j}oy�څPc��OM���g�Lwa+��>'�q�;YoF9.�-<�=���$G3����� �[g��綇�o��s8c��7:˛�2�*�`�Ҧ��]������ի�`�!�m1C����s�Z�f�"=�^�;(gn\���l�����g�jB���y_�����-������.��Y�v�{A����v%o�W�\�~!v��Ŏ�^̯�.�/���U�{�O�rv�fAN����OEv��]X����g�� E��f�N��}���"��ç{	�ٽ�e��A}������·�օ�%>���'� �G�v��m�!s=�M��A�)� +���P��Qg�2�X䫩�9��'����D�5E�,��Ky�;C��4�fnא�c�r4n}m����UY��x�eF��RvN(v��m�!�V2y{yQǍ�g·E�i`Ț��I���y�Bɵ}�ʝ��W6�����<XP�IFe�a��"��.�e	��{C�tp�RGov�(C�!��{.��~���ɦ�@�3E�&��%��Ğ���V�ۮ����ƨ9w�Ԅ�ݾɵ�
T��o�5�����K�#����Yﾏ�ﾈȟk��8òc������Qu���=�������`ΗV�N 'W�j����N��_S�ZB;�3�����^�P�<�����o�בֿ^�mٺ��V,�TN�����|Ë�����/���*Ǵ�+���W���=�q5/��K�fco�5L
^̕����[��g�j.h�X�G,��f����}��v��OR�)\�uc�P�{naߧmRߍ�^(hd~�|sq�b�,ξ���wۗ��D���ص�`ϓP�ڭY�.=Z��29珨Ou�s�w	T=�ld*gۈ���k�7��fVv5� �@��v��z*~�o�=?m��TAwc%sN�]C~u=[ΰ��;�����3��J|uWQ�#S#h�9{�{�?xu����üpf���w%{��N�w��IO�ɛ�>[����m���~w���i�oh�>jዷ��AC+pω8���n(���o-]�τ���gt����)���q!n�l5N�Ǩo�p��ae��x�/fd���&�Ǌ�MN*�/)�-;�����Gf�Y]�V���tB��M>�s�Еp&[[Gmw������^��}}�}E���c�N�~��;�E���}��k�i�nyy�/L.�xez��v3.����}G�F_J-���˒#���kHd����>5;��
3۾�-S�k������Y6z�����G�ߪy��w���ĳI���=Tpk͟)ݙ���C��3t��s�ً�$�cN�'[��I��)E�t��q�4���C����`F�л�޻�	��f �#o��o}�Êwcr�ƽ;�d�*#i�_=���/;8��yN=�Ə1�78���c������6��X���9�P�Y7�욤�M-S�t�n�UjR�Wf��`��j1XCQ�ํ-�ϖƤjO��ӽ3��4~>�FF?2��=~wV�A\�uy����{�/+K|�(HG���z_S7�����K���é��CܹV�4jۻV��jh���8OE�4�z��Ϊfjl�J���<U)�`,�N΁�hB��N�,ND��
I�M�r3m�Ӻ�V�5�q�
�+a�)b��<%d�ů;�v&�p����n�dN����2%��F�]�B�7Z���u�7M�A.;�w9S��PG�c��}�1��ʒ�T�*�A��)��Ԓ��l�w�A&�4�t��50��(��,Y�9�����<�|�=��e;S��'��td��&���eF{%�r��6<nl��k�˲zL�x��A�#�����Ex��ՍJ�Oɘ.>q���t��43l�gJ	�d�K�����Ww91�r� �@�&�����.nayl�Ҋrv�����E�
N���}�#Tl7ެ��
ڣu��h��_[T�`=w,GFk�W";'^�f��U�ۭ]p���9g,-����EY�vy{T�B;�G�m�PV=]pz�$�tQkB��
W<�]B��\՚��&G�+&���m�+mM�}LXEYZ}����Vɫ�G^�ܻNZ��*�VX<�A7
@�A��^�S��t��%��Ƀ�(��mW�l
�Md'�=��
�oB�s(�;H�U��ڤ�}o�m�Vu��̳X0s�%Ɍ˶����\Tfp��uz��t�v�u�y�ٸ&��Z!�b�<ˢg���=ӝ��)f�.�W7�<����-����Z�U���`i�
z�p�w<���=8'�w���É6�'Q�7k��/v��2֩|��L[�jgZ�::΅�w����w���x'�9�K�34hHT}�"��>Q^M�ٯ�������V*`�$.n������٫n��i��U��6��n���؆����%]kF� �;.>%�H���J|�4tS]Ձ��ۣtRn.�D\�U�6���
�N�Q�D|4�wF��V^wP��l`��Q�ĲT��¢�bף��g+�Nn�oV<�"8��c�����av�I8�A�.j��|Hȑy�-��f�c��:Xw�6�2{nU�� 	X����h����w:;w�N<�Q����N0�q��S�,ef_	���o���N�=�\����%��l S���KnWs|� ��2�{�R�Ct󡨮��t9<+n��&���Â���݂�eZB��O�����sk#V�����R��]\Tơ��-d4m6��z�`l����[��d��z�(p���9���&��Y�D�}g�����2133b׺�ֈpB�Jq�#u����1&D17e�.�pu���6��V��D_&f�9�#}��i��8t��s�r�AEa�k�u8ҍ��jNeS�q���P|"-�D游��1���|�F�[��J�xj烯z���O�g_s.�T)Р ����b�&��R�Pѵ��E�9qi"V�(t	�h4��Z�&�IQ�it����i)i5I�ь`���i5����E�4��-#N��(ДQ��M	�Ҵ�M)c-4����Ak46�h�Tm�Ѩ�RS@U��Ѡ(�l�à�CT�֗kA�1r�5UF�(�Ĕ���A�d9�����MD裐��
�!�M�4��9�E���Im�YJh4�!��M4�lm�Zt:u��խHi��sr�Z\TV�d�i�Ͷ��E���nr�lm1s!����Y��" �'Đ2K;����ק���^虪1]���*�+w��c�%�r���]AQ�I�݅�JXL�3%��=tՌ-�L^���#���^M��ǜ{G��q��a��[��A�GZ�#!O>����ض�#}m�� �Z�����P�X��ۜ�G�dl�E��^�������ܕ������oJ��&!T���nk�Z�'o�&Sn�<�P��*Z�N�U���6��dY�/���!Cyӛ�s���|����J�Yw�P��cݵ�,WGx�d:x73��+mvq�h��'���M����>�I�=Bb��:�"؅������#3�o��{+71=uϭE������zf�*�4�[�ug�϶�3��g�I�8_Q�焊����1�g�W��ؙ��6�y�m�].[��mj]f��ni��H�W��}�N�o�$��L������$e uusѝ��ՙ�ޜ.'�k��i�_�j�V���ܔ3�J�3������N.e[˖"�C�d��e�0Hk���-r���|Z�z���绻���v%@j#xy�����ǋʵa̰U�q����Y�uk�",��"0�p�]u1<c�%N�8�ν
�h�����gb�����;�i�9Ъ�\���n��I�WQ��8�So:�-3���b���U}�}���Y�e/u����ו��j�H��:��%K�ɖ��F���Ž2ܤ=\r��K�t���7��e�6����DĈʧ�i}^�]�s��v��\5�wh>��Fk3|���M󱔻�9)�	;��v-P=s�KVT�~�W?C��r�3�Um��R�E��X�3�<�0D�{gq�4z��+���y:��l����=�[���.�g�ƕ���1k��r+qB�z�����c�u��7V�"�y}����{�Ԭ���=��_nq�k(�m��aQ
j�&UM!1_s�T�974�uSV�=����6+?���j�e9����F�~����/d��8T��>�q�����8�q�Z:o7�S�J�xj�es8wzwMx��)@&�ͼ��b}[�5�/��rَJ��{���������[&����	�,/m%��t�A�[�Scئ�_�e/��U���4��@��
�|Pz��3�TW}��|-���i�o��F�p/m��a��u��D�Vmum袇S2۽>��f]��-��V�Q�1cｃ��쁝��+>�%��
��V
�uz�����t.��1���}���2,}(�Y��_����Y�ƈ�d���͟�� ��7�9��*�6߸ky	�t����r>?X���u���#y�MmE�ݛ�V��n%�{�7j}z��V�a�c�?cV��+Z!I�x�sMz_g�t��d���v\�7�eNk)�U	ܻ��G��1�Lc�#����!�=t���C������*ui��A�P�H���ڲ1ĳ�/��ٱ��^A(���:�OpA�V�I��R����z�͸�ͫ�Z$�'�ؠ�JI�F�\�1Ik�sq7Cj�3?F�y Àu���.X�f{�%:�4�;��U欙sC�p_�m[�52��8��l����xL.�g��z��9���\~J�잫©V1�E�^�ssk���|��M�a���G� a��5������ ܽ�2 ���ذ�@~���h��m�G,V�y�|����\y{�n�;�Q,����������X�!�H����Yr9/;��`Ѕ���<8Ռ�_���A��̗��9��5��"��?�-�K/�����j̴x�1@9�о*��%Z7=��O¿�� g�m�iz��K����#�9�U�ES�L�D��U4��}�]؄�y�qX�y|���=�Ox�SNW���+�����E;�pߝT�o]��r��]A�PoO)ɋ�]č��N�E�_N�r腲��:,={~��V���x���Og*[VX7n�����DW6��v]
g�8r�f���V�H�z\�_�������-і��n+o�O��s� �E�I�ug�l�V���Cp����x�ù��,���`�=(�o���Wn��HΖ�ׯ}J���}�m�~��g=�`��Ǳ�!�*��}�}G쏎$��b��&v���^��}���e&�Zkj�F@��7���ۡ�r~�/ך�/�K딩w0�T��2E�p>��2�� ���7]�v�i�
9`))Ľ��}X�^�Z�_�)D6Y�ק�ǜk��'�P_O^?,	� ��2"E��x$)
�cU�Ջ�fɔ�2�zk���E0��\�37�i���oU�7�vS"����=����#g pӼPu�F��#-�n�PW}��k4ů�7�q>3j�q��[��(bXo"��(�X�4³Mm2<Y���Nonŭ���"\���B�ncޮ����p�(���(�}��W��T�{���dH��������!�<�Q8�p�m�%��W�$�58�L�F�N^��N��|}{`��־�CV�k��t�yq�&5��ԘS���~���@�[�����j-�����Ʊ@+��y�=���!=ϸ�6��v0�T�=��;��dS��(P���n^�Z�Owpnkmy�����Y����lɹ�)b�3K�XFB�nq��J��p
�S�o�߅�co��fQ��G�gf�.E�#s~��>��\]`s4��Y:�(Ǿᨁ�t?*��߹�nk��v��ew`%�[����.c[���sl����ml^3���־ՙv�m�Dӭ��z�=�u����l�:�V0�9O�"�w���fX���;u#�ި��`u��$�L5׃BǠ�t�1�8cH�����U���*]KG�T�-٥�+eﱐ�X\R�]7jo��lDO`�g�x4����Ƨg`��|�t7�\.�O;]��۠�%�bVE��o7ϐd7�GY�-������eKD��Dn:���[�����������~���s�k~R�]K��|=����I�?a}C�Q罡CVt��W�s^����K�~�m���.tƶv�t7J/`;:��E��pc��N�}��/��E��d)5[��y�22g�<�`����"���7Fު�6�l#��M����y�{�և]88��n�����s7���W��V&_�?^�͋�s��;ْ�M#�g����\�ܪ�NJ�s[ʁ�pQ�gP#�ψ���EĦn*�5��}�|��i�WLD_[�[G���T����UX��Fj�o���q������YW��������Gk��Y�0�@��eD$������� '��K������^���HN[N*!p��!�o^�����m��yU���{�Aך�Π^��{|�T����9uԠ�TϷov�1��t�07�r�em��N/�ר�igg���]8x�Q9�ۃ��h�{h�*������j�ށ���Ԟ����b�Gq���� 	z��a���f�t���Y���Ƽ��X]t����E^X�a�������2�A_�-S	NWG��3)=����v�fѭ�3��E�[;*��ͳ�Z�G�G�}��N��i��Z����g�`d*���u�eT���.7Y:��yb"�*A�V�[{�&l.ޤ��������\s~!v��Ɲ4B�u�^��0���N�<�GqvRP4-�O�dkǶr��E�ݾsV��I�׊���a�q��:>_,É�[N��o�d_Ν��}�N������Q^��F2�q9�ƥ\�uڳ��o���F��Oh��Z�ǵ@+��J?d|@Ō����H�i��`5Nw-�"�C�=5�%mmn����d߮�T�{Q;��Z2/q}�9g�{�Q�P7�}��aS43r���{���4��d��08�P���~�WwQB��+F{��g_�#/�Q�WIoT�b3�����yiǵg�%�y�}�e]#ype�%ⓘ�>������pqh��̖���z����~���)����l0��/_l�oj�����J�֞^���RyJ��=�L�����a]A&�My���Vu�����EgR�f������A�W�5�����A�K�r��05�v�P������N_�1��f�-\���Q�-q�apq72���qD���x��Nd�4Wu��Ϋ��cd�����װT Ob�v�)�d�TF�-����+G �轹��oN�걬PW!��a�N�n��T�Z���7b��L���-�\�^P����v􏵍�1C��#|�_��9��Ba�qY�oUw+o����o���T��H�5�ST]�.�cZ�MySXcB}�U�9M�o�Ƚ�r�SU��m�=�^�I+��2{�	��N^�$��Fo�:?36`鯯��DB�b5Vj�"}����u��w���/�<��O��ɛ�ϓ.1!Ʒ�ٯ�D-�[p���s�:��oFYW��g���3�Ss-��}���9��sŇ�&���{}W�0$!2�k��~��=(�1�8]�H���7I�����o�W��}x稄�Q���\��^ ؏��c�h�mr���H�Ӗ��q��wâZ���v�9D�o#��m��Ͷ<5Ҕ�3�Ǯˣ^�Ð�J泬w����j���2m�gik�]���%ƶ=�h>!g����t-�ysy��1�����-��|>V����#�������o�lo�­�g�����T��l�y�To1�;�V9)/vppۼ[��hF~��7���>����ڕ�+�<��Lnz��k�o���щ��<�1��QBg+Η�zXx����'�yjz_r4F8�����c:�����U���m���V�ҩa(�p��T
��T����_c�s��.�\�{�fV�j��t�\�r+j���6�8�y?X���.�)���ﲹ���,�Y���b�ʞ��ǜ�ڜ竁���gT�����_��ȷ?"��X�)\�|Y�BN�)�)�7\z^��᝵J��i����'�n^�Wx۴;���\8���Ѓ-��oMc QB�j��r�[�~�a
oyx5�GG�����)hQ��uwws��ڂ��e75�ef� ���m߉������B&$��}��X��[�`j!Ij9�W��@�k��9H��5-���e�3�j�N�][�n�ߺ�C���"Ыǽ�~Ӿ�*���3����o4�={�	�u�� �����#u\1��Y�΂�Y1���������+>�B�5����G������NN�d�^�ݧh�l o�*�B���:#�Sm��,i��3=F,��p[����t����k��FV�2�<T�
�>��Sj���&v�a��囀.�q�l��u��,ǀ��FS譾�3�m��X�E�.;�+�vgrY] ��Ӓ	�=����җ��'�n��e������FBs���Hd�vS{�؜&������^���\
G�W�ic��]N}ę�����"��n�	�����l9),���>�Ý����|;����ئ������M�<���Eʸ���#F�,�F�Z�=���1���-}��UUW�i}��Y��ps�J���W���=�?[�ЀjuJ��c����[�T�YNw� �Y�=dn����)ў~3m��jT�׶Q�o%���UZ{��S��Y
l kyK��YY�m�<��h�PV;(ܳ�4p�5��$�gY��6(�h4�f�3�K�OeOt���{����6wyB2�C]���2��tkF��i�L}�P�b�iQ|i��e���Ƈ:m9[\^G��_5iڑB0�-./,��՗eh��Y���L�zd�|�����N����|1���3���r��;�zʹ�ǐ�6Jη�Q�m�y"�]dԆ������"��M��xdq%˥X��8^�o\���AR�z���k�]�U��d]��L9&���8[Z�Và����������gv�էK��j�u�-��[=�^���N��˃Y�
�r�������I����:�u���+S#��]���O�W`�<Aatս+��&ʜr72���Z+��E]۰4$kգoh��ۙPZ\~hl���pxfƥ�-щ�[W���-]R�$����%M|x9�^%�c*����r��9�㋶�`Vf,a��O��t.������L�������szf�D5`�L&k�<p@$�wU�=���Y��M��X��W�]`�F�#�V���[����B�����f��Kr�e��:{�
`�	��s��xfc06�{���z܃[��-��k�!`�}��F"������mK�[v;�����Bh�&:��o���}�F0	�aw'7 ��3{/螡�=��U�;�}:���j��c���6z�X�d�U��n��NG��)�r0���wB��j����GW��ũ����.� l�^[�BމD�]O޲��;����k>}z��W>�z#
�G��&-���Z��X�yս������:����D�dsǝQ���ޛeF�ʁ��H��v���$�G�G�~��@n��2km<U�bu�R�]�&���&� �w�y�!*����zo�˸�s�}n�d`d��g>!q�>wӻ�4��7��k)#̸8Ch��z����]#}�%;�tvȹ�,F[-qN�6<g�K�1�ڤ&��}�VN��g5�-��@P�����=��9^�6�A��(#zr�X[b�����0��M-,�f�dZ!*���K�	��}�UMA��_,t��9ɗ�X��2��Ģ�kx^����Z,f��.V�޾�kX��YٶR��h2�+P-��+/�����^�hΗw1����)�BY�c�9d^��4)�z�S�j��Z�M0p��n`��9�h��M�E�+yޢ�ܗ=���r�$�8��'�}�Vn���6������͍��G1^�����Hw1�����E����moe$L~%��f��@�	7~�^�s͖��Ϲy[���[�9:�Ssl+�,m��v�%��t�KuĹu��d��8u�P�	��!t��k�uhg�<:'X���7��SI�Y[!pd�wI5*!��x�[fl��G�I�~c2@��\�zV�gȐEI�$�G��Z;��hޣGä�����l.P���;ќi�
#ǣu&׶ Һñ9uiݩ��k 9�>�ǝ�L],}3]�"�������'�%V�V��l4i���1��Z�U�Em�b
Ӫ���4%%���,�U��kE�a������l�)4�囔cUɶ������lDm�;mr�ɦ�J�AM.E�mj�֓F ��ikmZ1!��1X�(��Z��cM ��r4rM툚5�"*" ��9�X�J-m�T���lh��&��t��4Q��Y���ub�AQ1�	��lkؠ��A��Ū��*h-j1�PLD�,m����� ���
#d��D:�TkN�m�lmcXب(j���5M� �v^�u�e�U�P�#�Z��]3�ÝF+sp�ܨ�)nˬ�k�4�vT����_j�\��� 㜪(�X��ﾯ���������*sc^|Kr7!�$�c=PT���W��يϴ5Р4�ʳ�*n��k�y�3���}�˟�V�4��<�J�e�5�~4Zp>�h5u�sMV��T�oHފ�LW\�ud�N�;U��l��o՞��'P�A!�]V��B�u�d�]���6��߷��pXns�ٷ��m4�exl#�:dj̓�}{B�dM(ϲ�Y�X�UM!1_s�C=�<ye��ϴowU�STh�}�oܕ���\���7�Z�ʜ�*k]�ج{w����1v+�)9�Y}/��`�ݍ~{���Y\yf����s�ؐ<ҜR.�^�<�����O��rU���w�?	��k8�6-���;�������C�T}�#�݀s�`��p���o���=Wc��h���7�����q�5&��)o�Ō��?kQ��@��Ւ��נ"�V��ײ��mK�Yh��
��\��ƹ��B
y�b�D4���Ư/��/���I�E���-�_+޼{ܭ=���$��Bp�2�+9��U��<��H���=4�������Uh�yWpĔȾ�t�Ӌ����֚���UҪ� |-�q�̨f?�T�HT��S�D��6�<�%	�_b���*�O(�
�Lǆ�紣����Ǧ��N���~���KwUz$����oלJF�3�;�V��s�=���ܠG_�(tU��/*��*1H=`�UI��&v��)�]���71�n0y�8p��Z���S7i�j�W�.�K�cG����@)d'��_��c	}�1���i�Q��:�ͺ���be쓃�k }��`\�*]��n�D�k��3�a�u{;UOf�%��j�}<Z@z�p��砥�-�ޱ���y78kbw̱5��t7d_�V=t�YW��G�K|�b�ܭ�3���c"1C���V"o�ω�d�K�0��@�k�9����q�]�+3yߎ����n"F�^��-�.�~cэe��V����!��G�~�<���,���_��R�y��Y:�Q�I�ckn�d�^�k��S�Xf;/�k&��;��0b�5�����Pb��wi��>���Q��ĩZ��1ݵ�����C�^i1��{|=�q�л�׾~��F�8-ɓ�3�V�9�eh{Uz�v��=J௝^SaY���_�?�}��E���ٗ-e,��!Sҡ�|����3�y��!N�s�n�Ub��ت�y��P����c���FWL���Si��ӟ&\r�n|�����ֻ��z"g��?VNBx�	����p���e73�[!>�5�X���jw�����e'+Ɏ<���\�&&g�=<o���҈���v� ���N�_��n���m?�b��n�SO6�g���tu[�Ͻ�������h��UӷK=�*nټ�ǃj^���Zk�!^�b�!g��fP�zzj�4��\�O]�=�yē�FǦ�7�V�@��dm��xZ�߯m�=���K�{{f�Ϋ�/0�Z���'���T�������j�ɩ�EH�y��ty-�,�z��Ń�/��"e�AЁ�����݇q�{H\䪁�"��x���� �;��΢.�U킢��XC��8 |��ˋx6pH7�~����(�{���w&����X}A�x$[P���@9�mՓL!��L�}}���z>���5A�+g���GE����fj��m=�� ��;����A�95�-hm�e5ˣ�:!�0�3�UU}SŖeO!�jU��1�^���QӼ;l��Un��y�{�z�OB��E:���;��{r���g mTZ<������-���t�(we��̱�#�l�lXO #��}����=�����Ku�K�~~������Sa^��l�b;D�������?s�g��6�o|��̐��1����w�{Вwz`餵i���X�!M�A̅STӧnk�ZXL����yF��{��݉\?{Uer�D.߈��m�P��ӛ�zf�Y}sH�h���
v�<	iNwz#��}�-Ҿ�f<�<�ϧ|�}�Oݳ����δ��D�k�m���|���uʋ��ϙ�Gg�{b+�K��&�gf���yT}��i�$�!ۖk�7������b�+7��F}�:�:=�HO�}Yv$�C���RkN�kMmE�ݨ��q�ʅ�_��k�g|k�먼gSHAG�����&Ji���TN�)�tJ�}�`���w��x.��~���מּIހ�Q�S
=�XH�M�W'|���u4,C��Fv��j�ۼ���$�OU� !Q��1����p�e+�N�]]��n�e$��]_�}� gA���$nˤ{��qo��6z,+������`�~��S<2M���~�~k]��ʺt<e���i��>Dߡ&��O?hY6��6�ǗB�)�%=�3��66�d[Ͳ�ij��{_��&:��e:���C��C��^�V�;�4;�z ���+�hw��������V��q)�qU��l�%gx������&�}��5}<ew�J��U�w�R��č1�9��z?1�{7iƽ�n2e���m�6���53�d��V1v>��>�w�ι��w�RZ�+4l��c�N�ԑf�n��X��]���5��z��YUf
ai�U�mL���6�|�t0�O�o|��@�{�"�{P���+sz_����#+a�5�SH`�z�pI�=�9ul]O��n^��}~�yc6�n�T=��Z�؝T7�o 7��=]�X����z��Sԍ��� Q�I��9E\G`(�gj�������>4�lu��0�µ)t��m�����K�\����_�3#��p��;K��,�W��������*�"1Cj���{<���qf[��A�������Ɏd���K��	Ӑ���;��
����W��:Z��}��I�y�"���SQ[|7�>Z�����)��[c��ۜt�rT�w���j�z�J���3��cO��s�lad>�M�_��p�Z����=�=��=��?{q[�K�q�#ukϧu���׵B�+�Ҫ�����'g��U�hF@�	���]Н��;;��C���J���D}��2�8y���#x{g�+�*���#l73�ۺ���4;}�F����μ����?�䙈ly}�ƻ��r���ψ�E���`�ڳ=�wb�[�v�pה~�p&�J���{��%xt�?��a�K�N?UZzߊ�M{y���ړ�N�|/c~Je���]��-��j:h��w`�+(�[��W��"�O{h\Dc�+�}�/��U_X+��-���ۂ�4���څP=�w5��!�8V�hU�t�G_�Լ]�œ�7���5���4u�O�$��%�U�
m�kJ���.���]�[�J��e�=���3s�X��0����ޮl3r���7"�� �]��^��h߳E[{���׎���|>�|��fg��]�ϯ��f?2\�)w�.�=�N^��:�y[�D8શ�R<�r��[�U� {)LB�TܬѬl?&0Rd5�+����Ot���'��y��*����[f��T5�g(�_�Ƚ~���]bE�Ѵ�tk�:�<��̫	���8c�Y�禧o�ߊ.����w�}�S���7:�u������P����Ƨ�C^��5�Y���-G$Ĥ�{����q;^�i���dzx��ތ�����`Êo�/��b�]���m뎕z�nH�a�ǁ����y�ȶG����QܫAu<��J�t��G6Y�Xd�a������0��tӼs�ǬZ�[<��w���OS�ަ�s�א�s��Nv�f��a��eyo�7����Wnя�I�F�����9m<�s��{�m�N��l�{B/o"�X�|;g��Ϫ��{���tbM��	�������V)�CS�޹N� ��:e M��<[�x\�X5h��;!�R��GYQ�r1�!2S��On��K;�F� ��-���'}]�*B�Bݓ�ky��feh�ו�`�3�YV	/��%����;r=8��^Eno
�w���{E��c��p��ss�L#�<��fr��uzsUk6��v�	3��
zX���:=pqhJ�/_��>�r"���*�(�T����˥���
޿d��j���A�ҡ:��xv*]�d�^a����@��tʱ����~(�����S/�R���n��^�|�1�ҝv{gχ�ζ�MB����w�o��z�]������O�����n�]��w��Z�k��� �?t�"v�+?S���ej{�U?c�*�j=�&l�3�rێ5Ep��ص2��",� I��)bl�( o���]t�dڭ�w0nq�2%�c���Ȟ�!ڱ�R>��7R���+�i$�[���۾X�c�G��X�~U4�+�:"��O��Y�N*��2�o@\^�yf��M���!�z��V�~��ߩ�|�et���t����s�%��p�I�b�Ϋ����j뚷��v��)��X�fu.��g��\mi��G��5�Ԋ ���b� u����5�q"���T��\u	N�t��W�C2��]텻̻�wxJ��@��s#X�� ��mC�(���W�}�w��Oe1�[��O���LS�D-�x�`��f<3�S���a���{Og��.{	�-�z�<Y��$:a��q�k����M�!'K1w�x��y*������~Nr϶�!�Qݫ1��ý�P����P���͊�`T�jQ�03W��_S��2�������n�g�F���=k��R�u�/<;�CzB�����o>傓5��M�!�kv%�=N��1�=r-s��g���ܮ�'Kix��BO�|g���<�j�Ǟ���zcĆz�B=Cީ�%�R�u��%�B!Yǵx��f��g.��ُ��=�8s�WA�/�J�N#�Ot\J`�U㱯P\�gN�]f�X�nS�r'z�Yz�;���I]=9eY��{֡������d�[}�I�R�,q0���ʈI{3�XH��ޞRf�;�z�u�;WiT���
,�{�������]w�W����-~�j�6X�]����7ة=a%M�҇/���Uo#�GF��1�_F���B�:Y�̎1�Ncs�e����Oi�yW�1	�[;�X�*ܢ�@��W���Լ7
{;��JK���oϨ}3��1z����O%��x��Jݨ�z���.�1�Ayo�ڬ�jfVc"co���}�!ړq�\��j��%G~vD��f� ��[f���َ�o�+aX�UM�@]]-�$㽵��At%�ң�F���">^탻��c}T����7�Œd�'��g3�V�	M'z:s���du��χ?w��s�9�+^�k�v��J�=��/t����m;߲'�^1ɝ����v����꫈�u��,�ў&��r��F2�)�[ʸ���v�.�v�#�8�����z��L����o�Ō��:�v���~�_*������y�jD<�ځ��w���Q��4��g�<�jQ;]�+��w��&g�OQ^���1a컢�����ٳ����Q-�P�˵F�c�l8�ʽܒ%l�$9�'o��
W�����;��!�� �GXl������g-�5w�b	�dr^�Xے��bko�pv���3
���O�׼#	�IkW`+����Yx6lf
;���G��_U[L��U�=m����4, �t�ԍ�xGi~U��z�R˵����)�p��O���u�:�(.�jFّ���K�˳��`~�C�yt�����o�'YӋi����.���;��s��6��=7�DΞ�O/)0r�Om��9�=^�4�5�����_z1��(ۛ�Kۃ(0#��:vx^>��jZ��M�x�q�K4t5�b+i�e�mV����=B��+룣װYzX!�j>�t٢�4^֨`כCya�ʵ�h�C�2�(ņ>��� ŝ7|)Z��v	��kǈ��F�g�sa+4f����画�Ѫ{9��ۺ�#c�8z{���s.���<U
�鍇��\k+4���M�7[;�jo	��|����3t�C^N1*c�c��B{�E�I�ӡ�.Nu��; ��=���j]����3:��f�#�"���X�8�B�O8�/:Vd�<B��&���q�ӹP9�2pɹr`kL���mZ�����Ҭ�΄�m'S*��|oh��vs�qk"���B�c��J꼉��V�M�˭�l�j�A�xNr��=I-�(i+x�W�{3&�j�|Z����+1��8,p�҉OE��M����uڛS�0�Kk��� �6t+L��\���eP��E�ov��5.Z���]F���U4�����Ȧ�m�B����io��Ӄ��|+XV�Z'y{��|�h��̭��o��V�n;"ni5����,�4�gY8�+F�� >�.��:-�+�:P�܏8�Kh������#e��P�{3�/b7-�o
��xs�6����C�4n�@���lob�H��JZ�Pg����®����.�N���)@�p�y}���X�aș9�������0��`0��C6!�ml��F�o��f:�Q�!�)�t��v>.�Q��`�����7c��-��U���...h�͔�Z}�d4Nn�ןhy�ӥj��VwW�p�TU$�M���c[J���+/h�݄&�#�c�`A��|���+��ƻ��f��m�i7�̴��K��*�iŊ���-[�*L�֋�n�S��ARm.d��W��t�����>U}�����|.��[}V{�ﺤ\�˘o�6.��������W_������5w��>yt�0q��f1X��Xz���'Y)u�Z�'4>]ˎE�$V��&;��p�t�:����fh��t$��5���\�R�Xٵe쥯�^Z�}�C�W�>v�^�~ʭ}�}{뢝�����S�af֎a����3|�0nG�d]�$fuѠl7b-�]����T{T����o�����TD[�j�lRK�[h��h���cQ[*"���Tch��,L�1F�h;cE��P[����ڍ�U;j���� ��MDUmFKI�Z)��j�&5�����mY��"fJ
b��UPQ�)�m�f����$�����ֳZ�i�k4TLA��f���%�5��&�*�.���)�����PZ�l�F���L��QT�1D�Nբc�ECUEb�N��Ѷ�A1Vɶ��#T`��b��h�"#cM���t�N"�j�)��MQPMT�QRMMC�����W9)5���w۲}D�:����c�t��Pa��̓���*O˽�|8#b���V۷��]+c/j�ևW�">�"�1����w�,�k��5��煈ϣ�L����Aڂ�\<=��@�����m,a���Hq�~��&5�[̖_�z��𡨑W�&�t���j�{�����ѳe��:������ {�\%�m���q�%�ܸ��3�׃rU�{꿵��Y^��*r=�glUD����\�	XL����]��
�׹Y�\�_�©1s��ɶR���HA���N*Ὕ�K}b����V%�|~>�lW/�\K�
�[���_=�2vm���c�%+�9 ϲ��
�U��JD�h-��(e_b�ؘ�B����s2����LY�^�eM�u�׽}z�X�{�/z��B�ꞟ1���8�l�}ɋ�<��fB�X}=��=���Ǯi���4���=�S6:s�s��j�Y��;t��W��C�;4]��zK�b������W!�,N���
c`����*����;�t��i��VvM�FbX�o�G��Ya���Ӌ՗�aƬ�<�1�p��'�� ˢ{�j�c;�V6��A�F���C;D�sN���4�Ǐ9���v�{�:��}�ʔ����&�ø�-���k ��f<�<�Ssm[앲�w��,n��=Db}V=��J��Y��5�H��X8ޚOF_J_c}{O�p���W!q��軷���܆LL��ݿ��j:���ND.���W����v�rpn�g蕎����8L1߈�M�+��M��\�2��<#1�˪�^ww���[�c��3�ܫ.�
����F����K�ޏ��1�y��rY���s��9���OM�F���_F-q�Mc��C�}���/cst-�*��^ѥ���g�)`���
޿d��H�T�y���x�{�V���jTlhpu`��J��N?z�=��8n*�5��U�6�4eF���^ȷE/�6�ߣK��J�p���>�Q�~��{"n~�(�Xy�OU%��!�Ɍ!��e�4q��<�|�����+|&��U�7޵Y��U�,4�]D-7�Z���W�f���!�����ً���:�#�٨��Ǘ���M�J���e�(��Y�J�[�d�h��N:x�m��#h/�����Z�/Pw&��� ��ڝ���![��j��t��:��q������������Hv�p���<�#\TB��[�@zӹ�9�S�~��eO[�{W�c|�-Ҽ�_V&��7x����;����_=�B�uu
`h�{�d�V�݂��>��U���s*��|��c'Ϊ�ǔk2p޵>v��3[��d^z/C�ף+Yʜ�*ng݌��ǳ|�&L��J.�����2���i�u�F���b`ï۽;++T�{P�(�y/�gX�k�;�rA����MHI"l֨�}��i	��Tr>#g�qNr϶�!��)�A���7Q��]���nk;��c���&�0��2>8�5#��1|au{��FT�r���ŵ��
��^@��X�zJ���z	��������zy�<�M�C!�6����ۧMyp=����vH֏7����z�O_W���5G>%ٝ��X!G*M-�
[�tZrڠ�����o��W��S�����CcS�����ik�(;�`E ��ٗwm�k��������6,v���Jm�0>�ά؎�z���Ħs,h󳪮]O�)<1�7jѳ�����m���}�b�9zD-v��O��5��@>�C��zH��!��+x�#*@���ב�Qmvs}��wW���X*k��<�:��nИ�:���o/,]��j@S�x�&6B�5�S>ޞ���UWe��=��+���ɠ��C)�z=�GMFK҉�F����Z�ѷ0�%!Ѽ�jɸ���L
�����$�utG�ߌ?R��9`*},p�ک�Y�%�Q��=Q�2=�᫚
w��ںx�e�����fIB�y�-���y���_��Ϗ��呒�
6zxWڕ�����,F�#jg;�7�|��K����=�ּ��3�Z���ٍᕇ�g�>����S��ОjVr�O�;�r2�K��^!�xk>�����԰�G?I����D\�nk
��/r�2-���y˾����=�q�=�j�i
���_vz�/��Q�O�Ķo�ޟ��D\�K� �o]"lV�������"�e��$���2xP�״¸��κɆ�1��,/��hm���]%|Y������s�EZ[Ƣ�c{����P��엧=�c�#��G��Q�0^��nDt�R\χ�x�]v�jœ?<@>�<n�>/���A�7y�̗�k�yۙ��R������R�۫AVF�N;��[z���v�H�	3���Έ�#��)�y
�{���m������[���&.ȸPu�*�5��x�V��>��2ˉ�g.�)���j=]��
����,=;�R���[��ᾨ�����߱�3���,wmk�|�Y	������Zv��~���ґꅏ���_WbGy��L�n�Ib�����r���o�M����~���.\��q�l���+�ݶf��Ugï%,�=��
��b��ֱ���~�[����ց(qr:ij,TJ�=�@a�E���6(N�عǃ��Nd\{՚%U�ӽ ���d�ꄽ:��\qk<��z�M5<���OO:;ע����:�=Y�>܂���;~�&�a�������)�_Z���\��u ']aTu����j���^�=���F�!k����qWG���=5�K����|�ޯ����3�B�  TLs��ۛ�ti��{%	��ӧ��>�ZՂo�O�����D�?mT�Q�>��>ܫ�u^���q�z�l� ���σ�nhV�1��/�,_��˿'�^c߀��1�l{-o}���1۞�v	��V@����ɟ	�}��i#�qt-�������l+*>�������8��z	ޢ����ѱ�݈ՙi��(n�	�-�l1ƚZ_n_e U��9���9Y�,��s[y]�gS���
�����DI��^��p���}=�S���Q�0O�L��o��.��������W*��ib���;.h����$<^����]r���y˶�,�]1Qϰ��H]<H����:�Ղ��{?�d_n���=��~�`�x*�簾j���a��|j�W�B��ǾVz_�.�p�٘4z�n��|�q�/ܤw��aT5�=_o:c@�3�dз�2���c��E[A5�.�����,�`�9��q�0�1�	���w��#��;����~�-�̓)���涼/羓�o�@�_5,���^k��
�Z�E���c\}(>�P�:2��f'c�<r�F�#�ǣ�鯯P�P~���u�^��T9��tƖʚ�����Ⱦ�5�T7�9f��~9����uuGMƩ�X��}����������b�K`��l�%�q�+VE�΋����
�XuS�#�#��Ċ��ʡߌ.e��;��Mz�}e*��va�:�2����A����	���Y����<�����z�1�[3i��3�.��dN�3s�3���G1w�{Ǫ)�t������p<6�ӱ�9�wh��fL�����eEB�r����wn�>���t*Yi�{���ې����8����L���EA�f竀�gj����H���u����mڕ�i��c��V��m57��x0���5��V���+�++��w��N��w��Ժ�8�S�5?K�ޠә�l���Cx�rH�5t�6�*uSh��Q�f�W�s*�w��9:D�a~�g��,ԁ?s��Ux��:���������0d���32��	�׫��S�Y��3��v�yC�'������7 )���Y�_?�~g/霯�.=���Ј������n�����Kz?}O�yh��b`<���w)���P���&}&�r�4۹���-�9�w~�]R�U�)�:/֧ƽˆ*�`-R��s�V�{�P�>����l�o�p�Wo+��3��t��=4K"���r�Y~���zv�G��_d��� 0���n���t}�IWlt�
ck���.7�Ǩ[=��ep��#�Ժtx긎�Eۜ�^��ƾ�p5�ĸz�:@��gN@aX5~Wo�S��.ty���:��h���J��O��ޙ��������U���K��vDV}g�ә�ԗۓBb�v�r}��b;��㺑��̠+M�L5Q�Z�K�xk��螹�n����jM��I��T���([k,�w�T�ƽ7%���]&S�y���U^�mDC�tc���X����l�������J՗��>k �3F�ͭt�[N�>G�'}-+�/�-L%%��f«�ӯ��ע/i���$?3[%��ZV��MY*�w�r0"���ޅRᢺk#x�~e�iwa𩓞��3u����@]��]�L���֤�m��8�綋<''پC��^^������3�j�3Q�gEFk�g}�t��]1� ��w��q��;�}Y��}Xq�	.�Ӱ;�2�����]'�U�j/+��kZ�ϲH�Nt�,�P6�=�>m�q�S�@tf�ڏ9��@c��P�d����M�^�(|v+2a���7U�6n������n��x���h/�=����Ƨ¾i4D��<X��꺐2c�����v@t}5x�����[(V�d���E%���<�9�k�ޤ'�s=$V̐��}�eH1V���WC3ϐ.�0��w.�����Y���="a�.�QPy�P�t�5 O>�@���e)�+� \S7���}�����2��5cQ�j�s��j�X�C�&!��QC� ?T�IH\n��#�R�1n��+��~�~�&�5��LW&��������	�j��N̖C<Ogt�|j�q��^E���{�7Emv�ﱉ"g;��"��_�8�5��{�c߄�7�w�=<+�J��[��x��Wz����,��gv���C��X|y�r!�Jޜ��������_���N��ފȻ�G$��Um�;��i��:�.V�F~�ݽ�� ��蚥�����_(݄��׼��L��v��\Y���ק��/ࡱ׎wѬt���U�Wr��tΫ��Yn]��)>�����&�g�y�g��U�)<���u+
{�Gs�F�?��}��B-ߜҧ֖~T�^g�~�Q��P��d���T����K�Hy��5q��Te�v���~^%�zՃ��DZ����a�΍��a�@y�G}�{E��]�A�d�1�e���s6����i��y,��f@��l�8�tK�:�Ux	�s�2*--�V��49-P�v'�Γ�Ԭ%���v(����<}�9�����W{$N���#f��'��@T]�f�&��)pu�wM}�p��9=�]�癑�����㦽LIqz<�k�`?,��#���|�Z��W��z����ZqDș����HY^�p]3�|�3���z�hI����yB�r��ld�~�.�����W63��;�3���cO�a���N�~G���] %ܴtT����@��=��<�����0|����s�>�<:s'TB��J+�q�M.��KSȁ����w�_Wf�=[�f9���
��R}ˆe���j�xN�N���o-G��}�;�K��ّ����5�6/�Mh�ӱ�����Ǯ]���1,�ՙ�&�ӷ}Y�3?<Y^V|�xz��k�5W���^ʷ=��s�.�3�t��=难�}�nw_6ŧ �(]�l��dn���*�g��J�>�'�����ӽ��n.�����A�:kzS�ϻ��j��!���w�3�P[C�p�1�ڗ_<��Kח�K&3�z|�v�ϑ�~=>LX��Ж+�7&|�@]�{�HR������l��v����@���AO�Rx�@JGYj�a�޹�J����'�!�㸩��S���~�ӧ+��Cn@Zk�χ[74+��PS�����*ݛ���.��=xj����4��ɝ��Օ;�/��َ�j|��g,�]�U����}�ީ��|���GNWx���f���'�>�]^��y^α�;�[]�@_F˨�.�P+r^r�ۘ��g�!_��#�|�A_�I���D���>)#���kǅǭe2��C���=�w\��=�E?���8b�m{#-!Xw��_�����˜�'R��ﭻ�*���@k�C��n��D:�����{ˍ_|=>�q=N��'�7ap��-Wɫw�� ��D핬�Z\7���0�Az:�x}����<��{@1__^���r�2����}:�
�U֫Z�(7���G�,�N{���΍΋}k��o�ߟ.�P���_ڮK9�rw��=���}0��3}��p�����*㮾��!$T�7{���:����;�jS���z<+/��Iʧ�!R���-���c�Ӷ��Nd9�є�k�q,*�m�8���Wl�'������אY+�c+QE�:b�h������X\�B�����릍u�&
Z�z�qu(7;���k"�
[u�ޭ=k)���֌�vi�bR�c;aX)�]�18[��ŒJ�*����mJ�S'WfX[)�=-�Wt	p-�d=7-�W����Q��%TWgM!/���v�J-!mw�ެ�"���>�`��U���>gB9�X吺]];"D�z���TNM��'�����J�/�;ÈN+��TzsƆݨ�Ҟ��
;�R���V�Wrhc�XT�	33{�-�H���r�P��B�s6��j!3k�>;��
�F�+fv�i���X�na�N�y�9)��ܯk�NX��Z	k���y��>�oo/��Z}+���&�o��r����h��١T�������j���o�һ��y`9�������N�x��i�[<��qZ�f3.�9Ʒ*E� .	�'-���=�ˬM�o�y�H���_�
���ݎ������y:�H�M>�����{�U�1�R�<ɲ۾��y������.�Չ�D���<o���Xw��"�������8^b����*Ne.L�w=B�ڑØ�ϖ���`�G�eP��[�}�T�G����F��
�PM���ʗ3���ٹN�:٠���Ѿ�'S�-}�pm�+Q6����\+I��p,���Ϥ��v9���&���ɠ�6�GaEts�Ўf������,l��ڠ)�����V�Tx��YM�뮱з��ۢ���!��m��+]u,B�{�<��f�Q�r�{��c�:�q]��3�2�:��K�;˽�tp�ި:�s�-V��3e���|�bP�W� �M�6�S���wapyp��-��U��%���W��hah��oL�6��x��}/�k��1��r���,Zom�����MЫZ�vE��m���=�����+l:1�o�/e,�ci�/`��v!��E�+u�W�UŻ�C�c���uΦ�|�'k3�m�y䷢����V��/]�(hݡ�1�Z���W��������(<\٘�κ�Eo�9��:�z���nC@����j�u�ѫ�\/O䅈�-�H��`p����hI[<w*�]��m�� U��`�h�x
��J^�Ǧή��a3��ԄZ�'՘��˽[�� ':��g1�7����BlU.E9�e�6�[oy��/\���oo��{MY
��ނ��y1mW|�>���.���0�FsndP���v�KS7v�NG����ePf)��J)�ں���'RC�����/5�6gpw�]/�п���IŢ�� �����a���� �m�WSwVޗh ����j̍���`%�(���*�2{����p��f��s�87���*���3�6��@}PH~**��TE1D�EPIE$Ah(qQ�l�(���MU4�E1�SM��$MF�9&�ֶ�3���h����-��kb�����i��Y��ERQ�V5��i��
JJ�&66���%�D�KS4�L���P4D�TDh�4�PR��J�j�+F�lD�[�f+K�"����&�(4*��b���[`�D�T�Q0MDV�IF�D4��L�%���3QF�4i�i��EkMM��T�MSDlj��i���V�N����DEV�h�5
��[kY���j��52S[�ڊ������B��b�E4ֳ;��Y����?P�P��Tݷ36E�˚R;d��b��J�N�����ZTN���v=�zI� ����=X��S=����2����ٳ�cۉ������7]%�-����ܜP�ݫ���|�\fEg���0���k'���������pdF�é���t�$Wϧ�C��l����dvi�YV�&9��P�nze�~�m=>��&:s'Ǚ����s�6s^zz���=C����ǫg��dvj��q�*�~xQ���y�B�߂R�fs��1�S��w�z�.˱Y�|.��]�p�� {�w� Tl�gx��9$u]IF�K��7�>JdX��3m\�ݻ�*�8]$ɟ������1��w<��ړ�E3���ެ~W�KnJ�g�e�׭��uk�IKF�t����#�A<^�û�n@��\�P���3�d�?�O��wq��a^�ظ$���ngY�`,���5���ǟMW�]P���g$�7�ѧ�p�ֿ.����.ʎ���<.����b���^�2}Ը	���z����ɇO�~(_�-�����}���g��f��� k�0ø��h��/�'��� k3�,���2��5�w|�,�����א\�Z��&U�4�������X�ʇ�鋡�� 1dQ��x
�R�7���o7+.��#x����N��+UCg7iژ�H�mf���ɂ�v6�a=��9�%��mr�z?������:�F��մ�h����{��,�x'G�=Bc�h����F���RW�4/�v�z?�l�y^Ky���U�R"��T/}i{�G����%��鍳�D����*��z�~��_��a�\s��Lv�:w��J��X;�6����d�����	٫~����.nw��ƞֶK���9������7�@�k��t5�4ת3PC'�ON�zk�}�#L���iv�q��y2�me����;�i�,��wD��ܤ�չ�{#؍nf�H���́�u�x�Wkx�-�߭P�k^Ί��9{�x�wWTp�����b�#{;̺��7�}��\��ٳ(X��/�E�zUZ���Մ�\s�s�ι����F��Y6�ᙺ(������z��uYA��@7���~��]��m��ߦ�P�C�B鋯!�y�*�lQ���q`;\����;�rF�<Xו����g���*���@����u��̌4<��lf�'��ن^L��E×��������@6x��;�@{��+p��d�YYH���=}��!��t���t�<�򨅫�uq�c��"F�]��ׯ�Һ��*�/��>����Fo"�H�����:�u��U���8���\Su����Q�K{2�{P�x�<���(���m��+�G=����m�br����l`�=��"ݵF����Zz���������v��b3�^5��ӪIcH�|���}{� k��M��~v�XOkm{$�p�A�$qg�Qײ��5������S��8l��q�C��z���9@S�<%���=�hWo���5����ʎ�>�u��1�8=���~ *����>�wv�=�q��H�ꘝ/�y�#y��N&ó�9�B�ӕfխ��;���6'.�F.���{�w�����M�f���j;<+G?I��B���e�i�
��8?����1��O�q���#��Cܪ0��Q�j{�'������3��X��x���.���:-/G��Tj��Q���l��Z^�d��H<��xP�{,*�:Ϊɋ���KLod�ŊV��2{�-W���_�8����~� �r�dY:�}i1�y45��OO��댿=�����bτ�m�́�="��,1���
j��j����Pv����a鼥����t慫�?-�a�]2�en�>��o��+���gnS.�y��~[%>wPZ��U�oV!��/��Am~�*Q�7�ʈv�5P.��ڑhK�o�(g-bw��|�ݫ��Qĉ�_:���I�Z7��KC�T�p�v�z�1�c�����_
μ�gW�w�В�̠�������{����a��cЯ^׿�*ds�	s+�o+��O��Ş��yqxV%s�H�������OOq�ً�k��z礻�@6k�X%��DJB�9�W�8+��cP���{x�<|��}�24��W�1���xv�~~G��T��''���(Z\���F�����X�+pw�H��ׅ�8���æ3'T%���8�Z�9��=1MO"�;�z����s�j���,��~�QW��&�����׳���Zg��o*���k�^:��8.�8����������w��|��S䛏w����^G�/ǧ=�����x�ɇ���{F{�C=�vtAّ�oU����*�Ԟ;��uU�<��<���+ޘ|ov�+�������Y�(Kњ����@{�wL�u���
���PS���/����^�x;����ݴG�H�;9��b�\l�v�|@���O��g�jz�Te�G<nB��Y<.�Ү���{:Ξw;9c�M鰬��r�<��;�_%��Fl��$��Gg�ي���7�Xר������L����w�TE�����j=�<Du�`��S�6����	e1��W�Kۮ���Ȫ)$ծfV.� C	9�_��e������
#2y*����y�ѩyO)���N��z��wJ�3�t�+;w��O��<���b��`㎹��b�(ӛ�Ĺ�>x�>�sy=I"�c���!���������t:�
��+ȶ;�k@z��>�.�~���{ U����^&��[wHU��5|��Y(1�Κz��O�Z�����v���p2'�N���Lp������3��j���ME�/��Qek5ip�7�0��~+���җ�Y�q�.����w=�]1£���/��Jgn;$	t԰+���+��DZ�h+�\���۟?�2�^Z�k)������}��o��R&�vi��h&c�H�F�H����������{Z�$��:�:�gw�T��9�+ے���|g����R�X�>	�UF6gn��΋>u�Ω��FUH����6/�Nt+<����t�a�Q�p�`q�}w�Ni3 ޡVEe����t����=�U#.���ނ�oس�/.f���82,ף�o(����B��������]�!1Nt�
�]��T�.����3YOJ�X��=�6�+��p\
�=�yܕ3�_�7��=�Z���e� s�:� i�	H�8��^������o3�pqԹ��������lW\���t��2��kg��f�1�x���<tQS8Ͻެ�u|��z�P�oپ��ۈn�F��Y�<��i~�6n������f�Ue���u��a�؝ʳ1�N�,�'aH�������8� �	�6�۰W;FI>�o��r<+��.�2�C�0\�r�`���q�>��#G�%�S��[�ƪ�;�ѷ��=�+��R����dLt�G�K�G��ڮ�\��L����->���V��<��FN��s�m<Ƅ�x��Vr�Tǥ�������˕C�>7����K�Ό=�A�r�5��v��Cq�@?�;.k?C_�y�Zk5����*�%��K Nu���=�� T)���q�����67_��F�<�6k�YP�=��5��W�< ������\��d��]���|��nw�sc�k��8)�IÇ��:�IN}P���U.�� �5ܛ��'n�l^"z=�����\<�Gsu����}�A���X4g����ju_ät��-����e�e���O9\F�ꡣ����;O�D9�����R㽈��w,4�ă��Ǧ�*yK��w7�w�?0?C��Qj��+贞��T��b�ŷ9�6�a�u��NIf1�q��+b��/پ0�K����^~˗�]��-6v��M�f���>k����Oo�h���v�d��K�̪����S��pj��9�'`w�e/��zVE�k���|�f��9FW����ϙ�e\_��
r�S'�AZ9[��^����S��\&�gL���t�G _�J}G3 �I������jM�����m�h�_>������-�#n�]����[nT5=��uɕl���=ת&��=�<���:fR�R>J�7[��9����[��S�#�kk�
���P�<Pmx�5�g�JG�'�v.	��������<(! 9��T��G<�ة���Oi����}΀����%�˒*7��b������@��ux\Ć��G�e��	�����|OY��1Խ3���ţ_9�jz���"=�$=5�*�㜱��3��U=��2.�G�[X����v�x\�{B���&1t���Ƥ	޹� /�w��B��TF̷�ò�BS:=�}=Y��<�b>��ә<=��ơ���U��w���v��Y
�_����S�	��H����*f�#�o�Ǯ{F5�����fW͙,���q��q�f�y�y�G��!F��s��+��y���\�����y�vʭ���m���v������F%~"�K�GeϤ��M���+�t��5rP��ɷ_�<Jq�ҭ��r�f~�/�}ŏL{z��g��n�>>��62��Y����5�ln�U{���}��V�ӷ��E��ZM�GG�r�(w�@Q��B�.�W��F_���:j!�x��/Y�K'�����N�;F�0��[���`�y(�7_��s�}���B�ZZ`��3�j�[~��te����+8]Ӯ���R�2&H{a�s�Dl!�7�W�>]k*Lgb��{�;2�px|��'�Y�S�E�ͫ�k[&[���e޷v�|vΎ������;�q$\�w�lȨ���E��]�A�FO
z��H�9����OX-��7伃����{@.:bz/�U2Eqk:�@�r�dY:�ZLo_�45�P���zqQ�{��)��5f��6�q�����F ��ǳ�&Yh��L\���Qv��%��c)pgҘdOwd�x���히�s��ή+��xT��e���̰5�IC��}j�$���ݽ�j��z�wF8�k�6�r�;���7�^���]<��f���r��G�xʊή�{�����W&��7�aa��7��XUiᘯzcj����N��5�=p=S�_4�:*'�'��x�ilǼ��������Q�+{d����Fy�ʠ|?=ף��,|��-q�Z�@u��B��@k�������;�mݺD�	��C�"�}V�JM���ςb��<=��N���o/9w'��!�~�����{����hћ�'o|@����%�Q���&:k'�ϋ���ŏl���ڃ��Uݪ�{}ۤ���9֩��m�H��!9G�A(u����߮yc�T߿~��꟝�7]
�dq��!��[xjn ��x{3�Ir}�nR�Y���{2�Cpo$Fծ��R�ɱb��_�V"y<_��Pg�F��e�]k�C��t������/��.Va�x��c��ws�Tn���H�%J�l�� :d#7�9���d��c�\�f�|�<g�e��nhM}�$��ґ~'Ǉ�\�v< �B��v=We��9��<��g�)O���]GW�U��#�c�g�k�ޫG�+����c y<Ⲽ���T^�;�0�f³��=��l��1���
ܪy��J<���lǰ{b�z�ݟ�=�G���>B�ċ[��֩��~˷�7/�9, �]OM�ax4ޮY�T�Mg��]N+解�\��q����;��5���٘�������rPc��E��#�羋��܌��uN�����cG��:7��Õa��1`z��&��f�.�c8�_��^�L����Ir�M1����1¢�ׅ�v�S;}��S�g�K�Ms���u,�;l����4���.o+�Qξ�[f��|w�>]���W�rYˏ9������13#�~���l�c:�����Q�qǽ6������"�������� \mI:�����c6:d�͐_UH����6,ӝ
��3�y8=�o,:�!�˯�z��N~yW��dj�*كlM���mC7�>�h`�(�b��N�c~8���P�:�`��ѹ/6�z;w^�Ű�����qK+����e��Gb9->�Ɖn�سX����*�KD��U7h��OU<����<��Vn�v�VZ��ڲ�K�΅�a�c���pLm}�	�Q�ˏUH�{�b��z}�,v�b�,T-��uK��E��������������[�(��j}�'�W�H�W�Q鈊��Vo�_z:;މX��ѕ�_{1ȹGf)f�.�� 6�]0���H��U�l���F��:��#�_�7Xݿ�%=���v�zJ��W'���}��7 ?EzIゾ*gY�]_�3	����e{ gH}�B�&<R��(w����/R������L����ߏ�F��������6=��񽟆�cy���Xxk�倩���d�G
���Tyw�S�0��>[L_�	d����=��O@��u����a�`_�5���5O5A�Md�ךኲXT���<��;UY�D�g��g~��Y�ѿ�s��Q�}6+_��e����h k���^M�_�������`����1�φ��n	�&|���r�����{{h�v��ǋ[l]�쥟ZY�*p�O	AR�'k������Ͱy@�=�$ǟ =�YU燙���։���g��eX�w#������O�s�jVޠm
�!���so+}윭8���GP���ٌ}�L��ڋ�Y������z����=K%
}zM�lc�����uxwE���z�������m䎛=M�>��Ž�77O��[ٳ�Y0ͨؤW�9B���j'XD��pP�+p(�����譟�^��8�$`C�Ac���K���7��6����+t%2�ef0�\N��UhЭ�y�fzb�DI��F�P=|]�����@���J+��:��;5��G���Z{����Vr>�D�4��IY�'G��d�ӷ�Eb����<�ں�k�zB�r=`���޵H
DL��]���//n��S���W8N��hM���1YVp�3w��}�mn��U}�L�-��fm���J˖�fl�D
��,�*X�۶P�<���;��ʑ��}�{���2f�y�� ��ێ7K�1MԮwf���s6/R~H%�9Ts��S3��2��\�ov?MWj�y�(L�Y�/!\Q�6�=��{h�yڠ$ ]����iE iz �J�NV|pm޸P7�2�{�Yma�8[jW�;3!�q�!�7�|AVV�+ׯ�4����|[g��D���te�o��+z��/g�Å�WT����Z��/�m"����ms�H�wB$>��=t�G"�2�M�l�Sa�v�+��Y�i��Kj�m��-5Q'J|7d�!�`���O�B�U9�9g�d��E�/W^6�A-:�{�7Wp�`����,�f�N�X�+n�;h���XjE�I�yOnL��S���wL-�c���7xb?nαz{x�c��&6�x��I�q�<������ې��=��n/���+�C��nb��sn�����m؀�*�:ͷ؜Y�ҳ5c�Kx�C��v/,���g��b��v2�A�k-��ר�ŭ�,�����J�v�.�a�Ts�*fვ ��=|�1C$�����~����ڶn��1{m�8�đ�P;=�C�Ch�h�+Op�;��)��9�"�B6��ݐXt�.K]����nN��� ,w$�n�n���-+_i�Z��u�5X���5"ibEq�Wyh��`���l�$p��m�f�0ʒ�� �4�mm5D@n��|C+���S+d��Ћsj\���]��� e�R�_I�TeѠ��A=5��uT{~k=�3���e囧,�д͍�]��!n�*�m��ۮ�`r}z�9v�n�Wv��N��pT�v�w
r�B}�&<�0 �}�����{�8)��z����O'��[�R���%��勷ѧ��e�2K��/�k��%'���y��R�J���!<��̃١��Om�X︰3�+s��V:��M��AYX���V��:`g�pc�.U��6�y�N�����^�5֡X��,6��z��7|Eu+��3D�T����A��W�S���0��{�W�c~^�9;}��
��7s��Ͼ� *��� *� �Ө�$��cT�M�bH�)�"���[&��b)����f�bqh�(�bJ�"���(*�����&��JJJj�v�TRm�F���"���F����"���"*�t�A���b��!�(����[`�-���	F�l���Ӭ�L�L�TE:U1P4S�:3FƝv��U��PD��[F"��"!��)"i+F
�
H�:
d��h(���M�����654�5M,HF˨��ch�l��b��i��֕&�!��4�jV�h-��DCD@ѧ�3,��9�F��iMT��1kIG�#�#Al��KAQ-:5D�%$TR:�n���s��:���PM��=�G0uJm�����=�@s8e��e�oo�q{gi�˖�Hw{i��
�DnXյW���,_�'�4��*���xPn�:�N�ֶM�r8�ϭ�e�ݲx�veZuOl>�s8�^�߳og�x�U�LWN���ZX�����T�ď}m�x�i�s[P��0�Sڀu�d�
�����4w�6�a��B�=��/���/�
��oQi�����k�ь��bn����1�9~a��o ��^��gf�\?@�ٞW.rDX�K��+-p{W9��s;"�Eh5��=�-u�������🫩��t�w(6�<��\u)���زm��{�7f�c8#��q��d��6�<yx�n���"���4Aޓ�C0q�Uԁ��yЙ7B�\�_������vn	�3��_/L鯉|Z5��}�B~�3Ȋ�ْ�}qq�1�{��W���H�o�*G���HV�ё�����"a�b���F�#�w ���k�����I�B�5	L�~���x:��b3�:j2xzuI,Lj0���[4*��d�����۰6cv�ݴL�?kG�aS1�����]�cX
�c��j���,\ 2�ɗ�/Ӕ�m&��5�rj��v��2�lu��f�J�����ۥ5�]*,ĝ�D������U�<X��������k��p���zN�`��2E�/*�f<�,���ޗs�R���*�� ㍽�|��hs�m=�]	,	�]�v&��I�y[�g���:9�G}�d{����ۦP[�/�����ٯ/��a߿�� ��*f����gǘ�nvptl��~��v\�Ou���{��k��V\w^'�;Ӯ�f�e�����=ʰ�N􀷕q���o���{.N���8pr�ﳴZ�=�~��^ٔx���V��E{P�X��c�
�^�B���]��/�s#��.���Sw5n���/��?2gOB~���D\��ّQ���K���H<���Bc^�
�γ�ہ�mj��>�j{z'k`��S�f��]�2�9W����<�_���KY���޼����63�Z�yQ{�1�2;,�}�:գ�}l���A5��0\l�z_\�赝�����8�sڎsXf�h�Ucu���6=�����j1���0r���۔˿��mTrL����#��z��NԞ�����;��K���K�=�^�z��-�1��{O��^s��A���(���l��w��/T�����#�g\�x]�xx+/ݨ݅�xj8������t�әh�L3�gu�yʿ��H��>D��j�[�N���2L������o��Z3%��.;��v�@��L��ۘ�4�D�Z��^SӔ̡��X�����^7H<�@&�O��M�����t�p�[�WM��_`ǜo���}DY�Z��e9 ����q����j���-��z�Mk���/����qՒ�z!�8�5��Y:��l�quol]�[+��}�e@��;�a�X;n}DxU��'�mp̰���\O	��>{�=�[��_e��b��荕�m}���)��=��)�����c�.�"���r��`g&�Հ1ߦg��)}��W#��ɘ�r��C��� :���I�du�s�T;��"�'�v�(���}��S�$�Q��uT�ԏ�@.=�X�f�Dv��y/�&rxe��Y����O�/�L��m�ܷXw��fJ�<����i�=���7�3�j;f����d�v50Hꭉ�8�Un9�%�6��:<�'ƾ�!�U��e�	����~��J.k V�u^�:��Tg6r	�پ8c��~3�mr}��D\�����|��%�FK /���I��R�3�[����7ОՏ\G;������-�xK��]���/q� k��A�H�9u�Ku�;+{֞�=��k����ަ4_o����-T9Vێ�� ��h���o&A���V6� �b����x-e�����-��h����%�3�gns���b�W�{[�*B��no<�S%�{T�wFu�������mvo���YÝ8LOJ�N�e�)wll��f⏩�	zi3�ݢQ��=ۋ�9Q����k9�tP���D8�-�<����m��I�Ƥ{���:�8r���9�Gn����m-G���&��>�}k�Ͻ���~��^���w+�)Cu�l�>;��v��W�U�g.#�@tsјʮ��KN=���� ���o�W��t��zx*��ڋT�l��ݗ����p϶�
����z��x��6p�Ǳ����B�d�6.9Ъ�3�y8%�pV�ê�m��ٷ�%�߸��ͽ^>�C�ˉ�Y�w0����P����U�E�ρc�������h�����ͼ���x�`.�9�ޙ����P9��o�{��G������K��nv�\���C�ٱ���z�=]OF��Q)����. nw] ���=�̖v��*�q�D�޸��M���zn=��l��}ǰ����P�Gx��\l��܁?s��UFԞ:D��&��|��m�$��ŗ>��xT�?���ڂ�{�+�WA�2�g�1H��cD�$�æꏼ���|��L�ߦr�eǧ���V?a��X
�`b����������61�WT��iU�1�)W��!x��M�8�}���p��;���e ���mp�Or�V�u�O6���W�ەF���[Ӿ��D��]�5ʪ�� �o�Q�.^p���n��m���]��5bg*�.�$�[P���o�c	Z;��6���wz�C�%d���{���q�7��QVs<�S_�U|�k�fŦ=��m̞�{c�'`�Y;Q�C|i���F���~�A��4?������?e��}qP�3,�e�X�� .�r�yS*�n{��͏I��x�
o�p���|<u_R"��u�{ѸUyž��!~�j����嶺0��Q��@z/\�)b�l�ϱ�Ǝ���(75>sz,fm���+.�M�ū}����׻뉲}�2-l��
�L�F�ֶM�O�C�ڏ[�R��3<��W>�9d�^'g�Zz�a����	���V�K����7YTņ�Q��^����a�Y>��!�{�ӕ�eR�̙��Z<�H��x	�._�v���M����f�׳�wG�4+�ϱ[^�9[�z{l�Cr��Tpö]C��PmW$�v_�U#£%�������\���z|q��f,������q]~>�0�ܜ�����u�օ�ə���!�$��J�{�a���FA7�}n�7xVmT��V�9�Ƴ<^�dq�9�������\�Q�'��Yʊ�z0���Xoj���c�"�Pu[X�l҂և�t+	�h�Y�b?%to�ƮZXJ�±\Xb۾?��Ï�6D�G�/KF��/R�bF�o�]�ڛ�}�{�m&�^��O Y(�E�Wn��r�uM�ur@���:�_m��);c��@��㜲�>:���2�o��s����j�Gc;&:�zgO�|Z;	��#����QD(ֺz����-�Z;Q�úx'J����/������r�vf6B�����Cy=��ٱB�U�=�Nxm�v6�W ��C���Jgý���=yX�f<ׇN.��$�:�L]ߟ���T(rz�w�L�Vp�.����}�g* ���e�H��{��0��\��k^Lp�ʼ�~0\���>��fn<�;>"w�����m\Ш���PS�#O��^���+8�VI&��`����彲�\�Z��Z:5+�+rX\{)\�>�د���E�r���g��.��3a~���t�8C�-Yc��|�3���_,�@���@Q���mp�;�s�=�'F���O��8��!QyךYs73�j1��w��*�/j��rj�0�>�sF��
g��Gs�F;q^�:�R���5�͎�<|{��N3k�+~��o�ё�K��E��]�A�d�:�XJ.��!B� ]���];b��z2oj=yޥ�6�D�5U��L��ܿ��_ZLo^M�v��u�����B��~t]r`W�O:�'�%�ֺ�̦is)��U����yg5x��쓪���:���N��:t���Z�A���]8ѐAZ5�	F
�u�szj��
�^�/�Z/B"���e�/iR��ؒ2�ߦ��r�Ϡ��³��ȴ�4��^(�n�*v����u���tp��]F\wH��!�`<���@���WkYK����3s;��W�|o��mܱ����p̾�Ⴚo����,��-��K@x�6��FE���mI�[����h�@�ڝ�-G=U���:���5/3~�^]N���\��~(�R���Ǭ�e��a�����mL�WOW��l�U���鍮���p;	�.���H^l���C�Ø{&3Q���U�.h��0��P�<��T�����,t��8:�KӪ+��W�z����=��C����L�����r����}DxLU�R�_[]�,.b�x��wW*1ǯ�Nyu�<%v��[!j���&�*�Nd��Jv���?����w�?l����f�KJ��������H됸K�d�>@oV���m�H
c{�
r�Ȁ���lߪ<r���9u7�ע�9��O�W֏3�J��Ƴ?mT�ٓ���q��	��E ���'�l%����˒�о��W��k�=ģ1��Q��_iV��g����W���ۯ�4[k�V'I��2�7uԻ��+>��͑V��+�V#��6k%{@>�|���M;�[-oq�g;�*��A�&��hgH3�幪����,Fڴ��'U�
�v���;,�ޭ�-8��VX�>��R��34q�a�R9gm��J��QPL����g9��?$]���-+�O��Ǯ��`�e��/�o��#���s���/{�x�f�K�^�p����E�_��#��hw{tYu_��?Zo!���������=٭)�}^3�{�6=g�.�;��T.��xû<_˗����A�?[wHTZ^�|@�<w�^�"Œ���:/8��}�4&��0�%u���-��FWfP�DPgr:j4	�~~���Y�4��s�Y�u�fj���6N�3щ0�1�	���y�1ºkk��})���]CR�x��j��ot��L�ܷV;@���}j����㱔���u�k1>/O��v�p϶f賳Gk�Bk9�/'�h�a�,�CY {n&P���pj��Ui��d?}�9�*=�/�Dz>��\���Tq��f�=t9mѼ�Ό��S���x���hLK��><�A�;f�rO��t�
�"�,���^F�v��?$;�?W��\fM���p`��QuR0r��o��w���`����?8��X�����>9��/�θQ޻�&��P*9���$�+�B�LE��͙zv�|��O�D�Hg"��w\��xC��Y��f�g#�duI��	^�f�ȨM8�4}����p2��a�J� �9q�ͨ�6#���§C�ɰG"�*�A�t��W��0i���]2��=��+q�V�U��ۻ�-ݪ�b��}�^���=��܁�e��Kpc(�>����k"� 6���@L;�
�4�w�R3�*���x�4��^��dp��(���<^�zΠa�gI�;��Q��1Ht��L���|=]'�9�^�ׇ-:hw�L�.�������c�/��!C�ԏ(}��=���ܗA�aL��{7�yp	�~��
���g-d�ʹ�x���c��X
�KFOTp����G5EU�(c?��N���t3|��^��qB�gz�C�%d��r}�&:��}���yO����,уփ�T�	Y��5;��̐eπk%����Fa�͊��3�6�>�O*��VT?Z�(�׎�f��q�7�w2x	����܀�֫�������sc�k�w��o�p�������H���h���ﳭ\�'�ƣǠo�1.�ΐkZʩs����=��uӷޔ� ���E�]�*b�l殽����&l�o�&��QD�4�
e�gU����ɪi�ڏn�b6)����
�����@y5f�POBw,5�4��_���ZX�I���A�LH����F{Խ��ɣ�h*;�pV���Դ,
u����Х�����y�^g�xҷ�CN�Y���d�p
+d�&������޳w�TC�5'�`V���k�k;�����n��Z`�|��q{�N�+��Ӻ�4	�Ͷ��إ�Ӫrc:�\c.;�z�CN@y{U�'._����*��gj�69��}�+���7ᝠ�1�6sN{P����9gj:���DrNe�mT�
�����=+�4�v�잜�����Fw���ͮ*,�Z�w�G��u:@TGw
�P�_���e���_�m�W�?=�u������j8gs��W=��f�&-��k���5C�Ȏ�!�NH�����)U��9��}7�SU��7�f���vԁ��6*i�:K�1��|����i�HO�H[�Dn��Qܿjh޲L�~�kϫ��㞈ʐ2b�ב�V�a�����q���&s2�V i�K����+chv@΍5 o�"@�R���Va�򱈼�����:�L����,�&���rU��c�r��:!�֢�v@~�c�*���`���5��y���k@~��c��j��W���������*e1���;˼z��U���^���!T���t�Gx�ɶkݝ��߼zY�Z�����Z��4��:�/, b��DjW�TnK�e+��zls���] o�����({�NA�J��+V��!��`F���g[�ke�os	M�K�,�r�Q�*acaq��Nӽ	��VA��d�p��C��:� ��R�]VB�}1==�!�� ��wH
fW�,�/�.��;�m
'Q5���a�t�G-��p){:c	$+����.�}��@�Cv�	���:����k���m�����z.�|�ų(,<�r�옭�Aog
Y	����'�Cr9��JѨ�VR��36���K s]z/p�zĚa-��{7�^�z����t�Z��)>8���Hyi�%ȗ�F�b�$���5(9g���z���p��PΨ��o���*��������NX��b�n�'�������}� A�����'=y��ϱ�fK�O��zI4�w���kE}�0������0kzqq�ip�`7HmY���'wo��{R!�f��s�����˳2�+�ͨ6��q.;����[|�4�TG�6�]p�B�q���;k%�i�m\��{kD/N̮�2z�k}�k'����X4eaip �
O>]B!�7HXu��\��	ٹC2eY�[4�n�R��خ��!G�������g�f�7�L�nk�O�}�'�{
��'��s[�2����`��/t��3v���T����Ȍ{r�h�M�6��X80�aT*�W��io��3i;[�c˫|��q쭴�Q����n_BS����2ҜܖM*뎆�8��nY�E�%��i"S����=�^`�\�@����8���.Z��K���E{����R{+�7�Nf������M��6��]8�>+�˼��S@+Lt��4�ib��F�oj������nc�:-�)v�{��ܱ��:%��[`YkQ����55�Y�����/��2�ۜ�⥷Da��)�8ͻ]�n����dRB֘R*a��+�;3w�;zjh8ŞC ����jķ��_W-��y�]O�ܴb"uw%��:i�WV ��2��9��(ţkA�lb`�thpu�F�S�oB60Gt$۬/u�n������l:fU�M��8[,�����[���q�܁�Cv���`AU�b��^�8ѡk媺j�6�f��黺GqҦ������]����k"^~���r�y�7k�g��؟'�֗n�t�]�M;��7gȼ�W��2�(��G����	�f�#�U�=k`�͎�}��0ŽDֳg�w��ش�j�y�ۣ���=�b�չb��l������0�LĔ�oM>Wv+��w������佾��k�yz�#<q�܁���Yz�08@���e��2�O�ot�J��p����`�b�{����T�v��z[f^��A���*C�#�R�q}=E۝�/���ޖe�!{�[��9��~�����-�4�1-P�LE)Z ��A:�Ğ*�Ji]U͆�����Дѣ�r�
������G6Gc!Q�%�S�(�i֊.���)��
)th��ZNl�tR�U��� �4�SAO �MU)HV��\�T�P�@kBRm�b
ih��ѡ���A�)y���cX���5J"J����ADE�r��m���U��αD�TSERE��Q[d6�P4D�J6��J)��&�Mdi��[[Jsnl�UIHֹrl`14�RLht�e
4��*合Z
�"�ذP��usih����8a�AAMPDP�@�Ϗ|>�N�W^uq�q]�ͭ([��嗜�ce���Nc�p�^�ĸ	�)8�S0>��C��]�юT[#�������Y�:��p?�k���~O�4���=V�����7�k\3��LeGge�3�wX>��;-�e���
�{м��w���Z^�懚��(w�1���$)��4���;��]��d=F��Ľ�5]�f���['�X8㪈���vdW֗��K���+'�W��9�/��\��m�Ê��ѵ����p�o��*����-t΁�r�dTZZ�ZLoa̟@�G[��^����,�}��s��/�}�S�����2��KT�0^�G�Lu��s<|�t�z�ڷ�����(�ړ��)pu�9�5�pܸ�0WM�p��u,�DS�2�֫�Dp��)c�{dِ����,�\
��g%f9��˘u�;����_���S�R�/���<��V��޺��^�7�L��wO��/�'���gB��O׽1���ϸ����.3m��w���%���p1r�zY8*vb[6`�~���&������;���LfN�X���~�-�bQ��=_�4�+���~��|��?z�S+�Ѳ����O��_�&e_��G�;�_��{c����:A7���\����w�W�*��Ӣ�R�J}�V{K@�wޣB$Uu_I f���#y�G�ݲ�W}aa�yZ�W�g
y-v)篳�T���b��f��U�D�t�^���T�In�"�5�I��k��w��}ԍlC�ƞm� �5�]��bH�vfE�������_�N���>V����.�@�ٓګ亪7���Y>DK�<⏓���\|6�|���h���	�Z2g���)�5�w��Br��	H�+�{;�L��F*��fC���.����#>=�W�>>���*#R<e��ƣ���w�R�ۥ �,��ؓK]����^���g������xm��s�^,qJ`8��Q� � LE��Ƣ;&|&t�ޡF0j�v댫x�;=���G�z����+����z��'�̋�X���]|�V����
x�T�v�k,��6�iE��ѣ_��1��~�A�-m~z`�j��A��u��z�l��Wz�
���>�
>��t.@~˭
�o�v�=�KS���\��x�j���@?�����߯�����s��:h��wM	�{e�N��z��Ll�������9V4�)�6~�+i�I����A}�l_�D�en���㄰�3X��^�<Lp-���Je� ��#z}����zvO��=[&���P;�U�TYA�W����u�k��|w��-WK�D��$7d_"<H��5f�CF�A�5��n�{f�J*����a�o3��C!�dϲ�����1�D�.�iy��ڋD��ʼ�")�e@�RB�ji�M)�f�^�C���=B9g*^���ne]i����)OuXwi|5:|��{�<�G�	��b�g�Ծܤ͙�
Y�5訡ds�Z�����L'��~ͪ���u�+�W��������uÝ����v����2&��>�7{FnN��,�M�gDZ�
�a=5|���R.�Y/����,���^N��éwu����ǜ��ݫKUȎ��q"�}<�yS���οE�'m����V���po��f��`��̀+�<3ݱ��M���D'���G���T�>f�w��1y�s�b���~�O��{�p���(<�
��w:Y�������p\&7�t�k�Tvx���u� z6d���������K�q]�oJ\�3�;$f���YF�x����!C���ɘ��������X�qݩ��={>����g����H��7�=���k
�Ŕ��:cdL9ԏ(�Џ��7%�mR�k�N�`�ӝ�{��߮S(W��_�˙��2��ϼz��~�Q��>�����[��:6�w����ǨW@�ݭ\�;��MCڡ�oy*�7�#l3�a���Z��X/���A���/�/�]S�������C��z��lzMC�M����f|�9P�T=�Ɏb��?x�j�3f��=ңǽ�g�}��ݫ6�5�Eh�b�M��LU�u���`�R�'�~˓�nѡؙ���P+u���R�4�cB36�녻2�r��$+$�Z;^;��̷&U���U�oF�e{nmx��3��W����X������vT'���Ԫ5c��?\e	��M�?+|����,�ʼ\f�.�@z5�e&�[9ݎ�\}�����~����߳ݩߕ�]�|��b��uW���?\M}iy����Z�C{�uP��=�l�����YR	[Z�Unda�qR��ڇ�@S7
ֆ��ڭk����ZX������T��(>��p̼�N�����O��A>�g{�4�}�[Q�6�3����Ӑ\mW��˗�]�⬶v�}姼R�xz){:�}����;zX��<��1{�c��������x�ڨ�^��",{%� ]��1�}�j{����W���z��0����<)r�:�o����t�wO�G���$�C�~[��|qt��"���m��o9zn=0��b�����^*1��zU�;�rG���4�[�ْ��t�hsP��_�@��Z�������Ͻ�c��i�%�h��z@ٮ�p�=�A��ж4���ZHĈ�:ey�teH5n�����\@,\쉇?F.�Q��hؙ��1 $ֽ�tnF���D��ЦRik�-�kK�S�-��]���p9�ڹ�L��]��4�˼��+�������Z��59M��1�h�pӧҳ����1��mO16�^\�Ⱥ���F�59�O�ٮ�a��ngQ=ʎ?�_ӥ��[���" tn,>�4*�0�rm���}���E�=�l^~��Ր;D�.5���+d.�IN��o� ��⹁�;��?Z'���{8K�7:+:���F�4k�T�끾�_Q2���=�.f�;��>�q��%��f�W�uz:ߖfȥ�@����z�X�ԏ�����p��
���'U���Yɭ���6!������#ˢ�}3�Q�qTFK (�WWMq͖I�=��~��<6d�l�1韨�S�͛���6z6vP�����V���{�F�����mp�;�s�&;��+��W?x�űJ*����U�ݾ�3�
Ƕ�Q1nk
�Kܣ̋k0�ެuE���:�V�1�VW#��D�ͮ���Gf��]�Kf�]��;}TE���2,�3D��1 �:����v:�T����{��ћ�Ъ#�[��lǟ\�1��&Y�*�j���LC�~2,�ev]G<K��m�w�U���Q���Gbz}n���bd�:�r	��+ n�j=f*��v���ky��ǶN��O��kp�Z\��)pu�wMF5�r��0r��i&u�"�P�\����S`��D�p�3�}��:U;�;��Y���^N��x[l��6b�V"��P:�9��o�*^���w
6�]��vmdr���44�Q��r<i˭4�=˄��i}�K�ꮄnA8�Ŝ�v��f�ԋ���(_B�����O��Pޫ�P����4|�g��l(�]}lz]�Q��7�u�=�y�P<Ѯ�� v��}�26�2]x\
gB�]ڪ"�&/Oa���N�Ψbox���Z�y��jI�}Ѯ�	�s:����\ό��=1]��b�9�zc������g6�	��������[�;�Np�ˀuΠ�}4Q� �g�����<D��Rk趸fEٯ!��5S>}�������b~�)f���o*���k���ll��T��y���桧x����x����B�Q�wMFK!11���|�ޯ�rj�q�ǲ@{���I����fzT^JCs3�n����.�����-2�QUY�?Q2X�ԏ���~�����
���`m~=�T�)?��'����_��z�RU���\z}^~W>U,qJ~gLu��[ y�<U\>ݻ�7;6�r�7O����ޫ�_����:����������`�h{�a`jss`[�<9��3��͆d�<꟦vU���~�ܶ��Ѡ���l�g�/-m~z`�i��~˷��jG*Q��������jv�I�\Q���}̴H��D\�6ͺX�to���Y>��5�ռ�v��3Kf�%QD��/��V�����k������b �y6$�v�~�\gDv8����ھ����ڣ�m���XG����;@����^�̾�Z���$���`���]��U�u���-�i��Ҋ��n����:�����c&s.{|z1�7�#%��1�XT�{Ǯ7�Lh�f�dL�P�Xg_z��#�^�1B���2��8��\ME��l�7��c}�C���z��N��;vS;�<�٬)Yz��z��m&����q<��wp*�kUPo��(m���,�9���]�yn���	��w������^��<�C9^rQ��ک��^�^�
��gj���[�;[<��/<���>����>Y�g�Z>3s���7<�|f��d�U"�'f��4�B�������\�5�4]��n�)?c����G�gb���.��.�j$w.S�����P����U���6�T*�� �y~��ܾR��Gw�&:cab��3G��ʈn�]�Bb��P+�O3Q��ŕ3����O�M���o���۩���zuE�	�^+L�s�UFO 6~��t���{;����,)���f��Cp��G�~�z�3{ǰ���>�
��&L��x��Z��}�&�T�}��)��-�E2�Fi�<�"�Jew��XU���~�%yˣ�8Z��W@@k�밯oy4xV�Z�3����"��r\�#~�����C�-�٣�vb�=F�{!C��-��6Tq��sـ�i��{'I��ړ�@)g���_��S�ǊS��NȘ{�.P��W��{;�c���Y�=�3�kv@P�T�P?{����fM���c����'�,d���5&&��
��nع�v<+�}�z`O��k�>S�7�V"����I<F��t�Gx{���X�w���U���z�+���f/b�ݢ�����Yݮ~��h���6=���6*��x�"��'����>�H:����s��+,{:=��9G�@�������Z�*�����sc�k��8�p�܍��梻/���w�)��м��ϻ��F�"�/�.}��xtgq.�@z/\�*���ٯ���/Y���}޻&��);��8���~r�0hP9�uV�???\ME�梭.ְ��uP�������)	{V�zgfdj��f���,����7�������$	f�;����&�_���ZX�^��T�O���R�j����ǃzF��ܭ���a��1����}��j��֕��x@��[�=�j��ǕW7�ۦ��o�P�5�tV5�r�� {�z��������K`v\mT�����H����"����9�)S�3;6���8�Y���������9�x �����@h�q��/bV�
ᇴ	B��ü2+��Ӵ��[�V�*������`ʒ�r��^uR��J�.����3s����Z�%󩯰�j4�G�q�ł$m��s,u��6�_rxh����zUE�k���}�a�k>Τ<7�]^ˌè�R�>�;FXqY���
�mvR���K�ظ&ٵW0��W�a�/O28��n���H�������S�]R�7^ӑ���Q]�GG��:+�����@��ux]�]�� :9��^��A�h�� 噗n����{"��!DN@~�������禢����z{>">q\.Ŝ����Z���|����C��Z�p��\��*6B�1&�{1������Ƣ�����>6-_��^�#\r�X�hl���7���v�L�sH�䉿F��z�-O�a�xt�_��G����yg��Lzt11U<+R,�~�G��d{��W4;l����^ݎ���m�M��et�������F�G�3�_x�8�0�zxTjW�V�S���h��"2o����T_���=ug��0�Lߩ*�/�x�s�J�f+��3�+5��2)��ioE��Ď�ng��Gxi�bz5���Dg�t�cڗ	�_�ҥ���O��g��҇��@�+�����8��@�Y�c�m��H�q�0�+��9�]��4�ݗ|�U�wz��p�;9}ff�����0�8�^~�������i,�W�q���9����|���B�v�������i�4������ҳ.��s����#��h���ѻ�;f��������"�����z�:�����[7���v����~�fE��s�K��q���,�oՒg}Wծ=�D϶pP臩��s�7�����쉖g��+��`�o�X��GpP�3�^U]>���k�͓�ϲh6k�j��}���ܱ��U���.c��,Ӕ�yȗ�V��o��'
��O=��Ѱ/�rE�|k�K�ӕK�ַL�|�g�����t�S)-=�k�B/�:���;��7�et4��qԤx㺁F_%�j�W�0�zwMx�<����'[�'*�d�*g��~s�����	�[8���(f�>ˎ����u�v��TZ��W�0�2r�M�/�3�I��N�퇗�̞?��W�(�}?�Z8?=�|�hy~���^,ӝ���9TǌI���"}Uuk�{gz{���j(��x����B�jy*6Bz���}��w�W���F�~]��f$z�y�F��D����h������Zf1t�ʱ����&��	r'��%3����&�~�����-��ϲ'�}�:��狜\,z6Bb~�FL����!�q�H�}R�#���c��g ��(EMF��F�[�;�e��*+����:�#V��Ɔ�s���fh� X��ɳY��֘����Rr���V8[,�F=�{^j��꫃���¨Z�E-uZ����Y�q�q%n�2¬�9�˯���y7xs�����V�!�q\�pIw6�g�>�P��⣦Y:�>s|������-����L��S���WYB{{�k��haG�06U[�H=�e^�.�U�8)�(�ި�L�xK�@�y�<�:���츩�F��sT�suz��l�:�q���>�A{���:�&���):Z:E��6ƛnGD��`΄r�K �h��������˗yZ��\���#qD����2��,�v�M�:��]+I�B�-�Y%�μX6��=s�����]	�/w��u�����[C��83�e���:Ƒ�k��B�Kd�q�|�ri�z��l̘�f%'"~{�B�}�j�8�`5�na쭮��iB4���c{��dvܱ���F"䅉����A1�{�,0�z���{үf��O�K�{M��{�z.�r��屎+ ��I�r���#�|>�5a�Df�ʧp�鶷��B�2�����]�����8�V�eEî $
��	tXn�3ŋ�j;g*�Zs|�?�3�,n���gw	�:��Nvڜ��.�e'�V�h�)_R:�eZ��8֕�$�\��H��^F�Vb.{�0jA��^�ZV�c�a���v*9o&���V�,�ώ�_�v+�g6�?+� ��F��ս��WE����I��i�W�Vj��/3�@�����7�$�Pe��8h27œ���-Uڼ�j�*�ڭw;/��&%�4� Z��,�p��� i���7���G�o	�j�X��Ky�@;�&�E�����ۣ�[:��`�FW;1�{m�]�cB�� p�/�[�9���xý:��X�G���]ӻ<�rk���E�2�ö똝Ӏ���Ktź�p��LŴ�5i�f�l��kWb��\ތ�ݨ%I�`�j�7�@oU3x?��4����,P���Ӣ
�U�K�.���>eB���3n����;��7oO-���t�]�َQ8/QVZxW&v�.��M�	7]��3Ցk��'�-� �-���8�����|��,�8��d���c�`���z=��C8���a�K�_VP�K׏b�jh����Y�j9��br�C}��s���ɇ��h^�3���oo)"�:�?L��W�o^M3�/��Z�B��
ѓ"{s��G�������=I7]>�3.���q�����x^��s|,c���7Y{�γ ۳�:w���u� �כ���a����YH�+wOK1#Z�۹�W���1���+�TM��TMR�pϷ7�/5흕�S|6z��ݧ����ee;�ժ����,=��������C���N.U�qM�m7��sd���\�("������s���0�T���wu������ (��P�s`(*�)4�k�QE	��s<�IJP�s��W,T�Z�A[.�#K˄U' �r�(��IG!�M!Z�@�).[���5F�KI@�71�(��) �؇�h�����Zщt��9�Ĕ��hA�yb�Ѡ��X�����������`�ʇ���h��`��IH�r���Ͷ�
H���rh^MR�yj��*�9�h((�V����h5�F!��QT4j��UR��Mb ��Mm�$�k@bh��(6�!BPSN-k@h�4�e��I��*i�&�Bbƣ�P��T����Q�4�%�A�ꀦ�X�B��&6X4�V��m�䜹D��A��ևI��hU"R|R�bk�C@O:��I�G�*V�/'^e-o�LT,�Ƿ�{����V�IV���oH񾼤ރ��d�SWn�ץW �wh�mw�3��c�bωK�K�*����"~���3�2k�W/��oUp��<���9�z���g��$�8��)����1j�>�OFOTuiV�~�DA�z���^J����ԑy��=����X�{�K������NWy+���yX��Cܰ0:o�-��v�7ًk��
K�jc���L?J�?G�R�;�����ǽ�l��L�U7�GE��3r�>�̽��j�
�����r�+�s�]�s�����1P�ᾀ~	��4Y{��V�el���j1���E�r/a� kߣ%=��{^�
���a�GvW.1��*=�B�9�]�3�$u����>��~���ϑ�t�w�'���,k�Н��z�+���$]��d�<��{��i�g�z�w�r��jX�:��s��V�Z����,���Q��sǼ:����+�^��}�=�T�T��t4�=r�i~�u�TE���Yl��߅�;'������ej�����3�e�xM��;��:���,x�l����K%��օbq���u4�p���u��<l޼Lk�]$����;��}b(=��	�/��h��V�z}堕��p��
%�v�U�J��O�$�w7*R��q�#9t��^���T=���c�����G�g	9�K��ԩ���o-#�w+�
���T��������{���>���ļ83ya�OȎ��w�}�a�\�|`�~���`��^�DJ��u��v��8����h��`q����t�b�,W�˙����Cu�:���!4嚁\�sF.�XM�*��*6���G���k)�%�j~��p<6�ӱi��� l�>tD��P��a_O�3�{�͹��N��ff��̔t��f,��d�:��q�d�F�x��-���ѱ4u��:;�:>f�	��΢�6������}��~����&<R�;PP���l�o�י��Nu�(܂|]��� ~�L�U�����a����c�x��?d�����ɒA;��V����}�^��pof����O��*��؊����I��!��ӆ�5T�=��}u��v~';�#��;��ܯ{��y�c-�j�@���%���6=&��ޛ���x�>˺�k������{�4����~O;�H�q�2x�� (�s|U��_j�r}��b�'b���h����gp�7�χ�+�D\ź˅V��x8���p�Ft���+�燙}��u��*�<d@U V܌��#�}z��S����ِ�H��\�C
M��_�륆���R=y�W�PeU�����k���z�.�q�ξ�8���R����TEr�c(�}\WK�I=��ϕ�O����w3s4���i��|f%�7��f�|( ���̉��:�u���5������U�%���j��Q_Z]�^��g/%�o�Y�j�fG:t����8�OG��8�ݘ�wz�}��Iܰ���V�t�V�Ki==�ރ�4���GR�Z��g�o`��9�Bo��p����k����m�f2��z�4��U�'._����]a�x23FL���S�����բO���>�=]=P���B�r]�=�[o����ͷ�{�^m��z���gV�=���0�x��Z�ϲH��]N���ʡׯ��3�inH�I��ݴщ��u)��~�M�^����5�0�6r�O��H��m�
�r�A��ݙ��\@��ܑ؆��Z���Ǫ@��ux]�]��>%٘�d�R�Ξ�6����t\9�=�b���_^�G�3���#�sd{���͌K��X��pd+��z�1T�j�^�3b�C�ѫ'Tih.Y��t�+�)��@��ea�w�����c=B�C��c��,�<W��rK�igHs�t���)'��1/��U*Gu�~�~�D����d�Tw�mVbd��*��F������:;�Ɲi����Aɜ��n�o��6�:0i�Gyʱ�/j�>����=x�I2��]�g���Wh$!��m:ko�p)>*�WX�M��]l�ͥ�
��r�j��$Vuv`m�w͜T�"��&
U�Z�;r�ά�oa0-S��>h��+�r3����pٕ�~�H�'�]'��dyz�Oݽ�R�䲟*�;a�m]n*��.��O��7>��|kǸ��`��O
ԯ���aq�˟I<�X���/����<�b���|ea�h�ג�}Yq��s�^,r��.�5�yW��OFT`�X>W�<���Yw�(�	��ӷ^|�Y�����>��{>��[�9�J���Y�3�}��߮�~o��;���8''����ye�!_GR�5}��Fvܝ:��Kd��s�����vdY>g#i�.�����>��쮜8� �=��¨u<�[�ڌ��c7��L�ZZϺ�@��v�Tl�.u�i�>Ch��s(~�,~Ľ�U��z�ɠ��dz�%��;�:������Q��%�����^ٓ����o`��3�:j=۹��%���)pu�9�5���d�����f6bĥMa�Buz���H����#ڪ;�,��P������/���w�0�7�t׋���\]�p�	����������?py7:?|]˒�� ٨>Y�Ґ�Dd���Ь�j�̘�� Og�^]a�w�L���$����*�w��@R��+�'�!�[JB��G�"��Ö��<]���ѶR5ٝ�cZ�Bi�3�N�=E�!/��t5�W6g�ՠ�/'X�ya���Ry�����+5���{Cm�����F����U��k���q�%�x�~��2��r��ה-/�@z~���f�#8f��9� ��=�c7���s%Gɨ���ָ]�\(�sā;!=5�ˉ��7=�C����59�7v��s����h̸	������4y�Q���}�%��2{WM�!���ϕ�ǾH��΅����/#c���FK��Ҩ�7��S#�ޯH����G�sT����J�G��/�S? �G�~E1�ō�J�E���%?�׿�H�$jG���iI�:-w�k�q˘�ӝ�{��
��AkG��Kˇ�>W6D]���c�S��W����x���^����C�^��G7'M}�z�;�V+�ґ�]��~�[_=���^�i�-��w���)|�z�=���_ :��	�������r�z~�Q�����d.�$Z�����te�ִ����+0���hu}���}��z�+u=���v����D�7��N��UGE����~�ЦGA��nm���մ�d�ǫ:hk���u=�������������9�q�ڐF��hƈ��˯;Bz&����B�g]ɡ���X��}��э�W��+���Qb��y���6�p��6�a�ʇ[�Wmu$R&���)`�2j��v`��2u��m��Ə^5��dY�o�W+�� ��([Z�3��t�=��*������;�{g�ը�������K�����V�Qip�7�0�1Պ��e1��ז>]�w��؝��J�P��ݜ���M��6�ux	�������k�(7��7X�l�/�ute���ΜQ��{�����j��ڮK9y��rr�ک��]x
�-^�
�6u��Y)qQ3�*�ǻ�b��v�1_y]��E�=���)4xT�Ľ6Z����m|�_���[Y�W3S'�]�V�!wѩ�꼜�.Â��T������Ċ�}<��g~��`ނ�rz�o|�b�����GE��X�6����1�0�K˙�]8��� �9�/��@3��;��kE�	U�{����De��1�O.l���}�0��8.�S��\�������#+�T����驲D:�n����P�Ӝʡ�s�NI��YFl����B�1�&K2%.�}�~�g�g���/k(�n@���[�)2��.���
���WU����t#��/C���4֣F�T�e�q��ќ�6��'�����܁=��2���|������f��v}Y���HL�[�M' ť{jfN�%p��M+<7^�����{&��C�Rk���z��o5#Dxc��^�,�r��3���7�k�yfz�x�v����W	O�^�=�hI2��Үj�j����6_='<2���3\�V��Q����w:����^��f^S�W�}��4i�z��*��G�oz�Ev�%[$���,u�����r�\�{�zcn<]�[bU���GC�3��2x��':瀯�%���c�jzlW����[p�8 �k[�L#]����NLvǽ;F��uFO =1�@�5\W��.�fÒ+��9J�nx.ݏf�G�[�||sg��W}&��E�˅V��W����</ѝ (ֵ�t���zk�2�{4�z+|�h�t�ZZuÙ��;uW�~wQ>�K�E�Z����gϫ��M߬�6$��}�d���Gw��}���b3�ܰ���V�t�Qj���q���_VK���g�l�Et�{i�
������_t��t�E��t.��왰7���#xR���S��:!��*�s;Qj�3�V���9~���]q���P�m?(5{�v����ّ}p)�e�����=*�p{_\�+잝�l��]�#�b�m!��9 C��n�zK�q>��eP���}P�^$�,��H�}�޻�6�zo���då��k�<�^#�1��G6}�'�Ĳ������<ёf���g+����'���~枑����`z4�0m����� �v�hVu7cYn,���r�ۆ�+cp���5������"~h�zXn$�;�;\[t��uaQ��b�G��v�-��iW@�Vh�w?��o����,��~�'���-g/� zk��.�����
:����і��\��j̏f��,��{{�P��"2!̐��*������^/���ÄO<���,?7��'��9�V�Q_CyV��Q��?oO"��]����~��՘y�[MG�/G�=��F-���Cգ��X��O�vOTU�ʡ5#�F�@	�(N�=�,>}K��QX0��w�y��'�k�O�c/�\��kS�c�̮�dK��=Q�t��iH���ۯT�q�q�V���pB��}�,]�k���6�~_|����d���up����3rX\r�x{�\:>�.Fff���#U;g��lT=�Zrט�W��.�=�����>��3����r+�;�r�5�|��2�iܱ�n;n|&���p�s���o�+��.m�aUi{�y�m��e-���>�so�o3X�tE����Ğ��ﷻ2�rt�w���&��TF���20�y	�þ�/:����g��n�ă���Bu찪O>V���/��Q��	3��[-GoG�%�Ia�G��Y!����l�Q���{E������"�X-���C���x���� f�����V�xU6��ϖu5�k�M.�7���b燞��k�R�;B�����A�D�*�.�#;9��t��R8� �:�n�b�����-9ǰ��.�Ȇ��g~�Lob���j���=>x�w-�*9?�w���3}SӞS\��-g��R����Lz��mQv����zn2�X�t�����0C���5��UG�vW��R�k=�M�w��-�ˏ�drZ�qJG�;����U�oUE��=�w�+��@�����}8oO}ݢpT?WW��{j@zD��T���u�v��Wֻ�^G{�����|*�e�?�ob�����5������;�HM9���0y�����LWuxX�F��/�.�;�91vߪ��{�:s'W�zuE��k�u��}4Q��/L�)��eU��{i9�`u:��� u뾿�~g4(?0�X�zx��)�Py�_l�i�� �w|��p�tdmS���l�\��{��Ո�T]ϑ��鯲X����2f 7��;�����l{=�C�;,�ݢ*�or��>��i����z*�_"'�1�R�}�.*w��Gv�Z�[���Cv׍� l�ٜi��_=��I����O�sa��j�G��Q��#y�=_�5��<v\+,i����g-Ш��Zn���ɼƖ�y ��gSB�8�'+5v
�-�Jj߰�n@�Dz��%o�����r�;\�@��)�ku�9�5�i���ʼN�u���[�y
��랲�����>�8^�[��������S����~��K�AzmX����s���GNWy\��4���3�ׁ�S�^g���G���<��1��(����m�zk��lѮ���g�/-fW�9�ז��X�������}���P�W�, ���U���.�:���i�~𗅮��}5b���S��������9�ц{�C���5�u(1�Ϋ���s�z�{)���[1޼+��ޏn�`��+��"yWJ���MG�����&���k��Ęu�hN��w.�v�Ӫ�Ʊ�;�Cz����6kk���7��[)���ux
�U֫Z�)���.a�{�v)�����N�ÏA�����pޞ�٧\/�W'N_������2��K�Qj��V�#U�wX��We��Xo�P��;�61����|f;��:o��<K�	�G� <��Э�\i�g<A}�VR�GA�:�gk���ɞӢ�yij�+P�j����C��â"�x�ԡ�'ݕ�H7�ިNڳ���V����
�	��o?�N�-���������g/�@TE� ����@TEꀨ��DW�*"�쀨���AQ�
����_�*"��@TE�Q�AQ�
���Q�TDW� *"�ꀨ����+�_�TE~�*"��1AY&SYg��J G�߀rY��=�ݐ?���`�{�w��
��"I)�P�J��T(DD��*��R��$�$��))R*i��z�z��R�JD���!PD�JUQH�����#�@ZsM�Z����	�i��3P�Re
��
�gR)n ��  v�  \�Q��e�M�4��R�� �Jvf���a�( ��ѡ��P�P�UURK�u�::  �&� : f�T d 4 	B�@�J�`�44 �lh� k@[ ���V�TUINݑ�-,�J٥[�L�m�Sl�T*��hV�T �K4"Q
�d�k�m���m��0P�p&�ڤ��ٳYI����J�J�(UUS�ENu�-5mCRZ��R��4�-�J��$*�U���lbUM�6�YT��j�����E�Q*"c!�)I ��` 42d�2!��$����  h    R&�a2#)��j4�=@ =C�S��)U5F       9�&L�0�&&��!�0# �H��QM2'�M�$d�h�f�=N��:��V��k�.��,��"u�-� ���Ó��C�?�%!6@?4$��C$?�l�HI!��}����������;�g�F0' I	$��O�R$�����5�I!������x������_�~΀�HuI��~�fN����)��d��E��/��������
��Yͧ����*�E!�S(e���n�B��D-�d�) ut�қ&9TB�n�rݙE�K�c-e�Ŋ\d=�G�dH*+�Z�^rb�2\ʧ	�rB=�pAX!���37!�E�J��*���`��m��Jr�g�C^�EP��A_e�(�el�2U�4�VSۖ����:g�����I�N-���&fS�vQ5�s^�=���ư��7dU�Ϟˑ�f4!��r�$��2�X��(�e=�A�v$bXخEoL�xJ�j�tn^��f�]��;T2��T�&��dk��Ʌ����ܔ�|6kƒ��͊P�4��=
P��V��������k���bb�2d�v��v��&t���V�
�)B[����YݷO(�8�a1�[�wB�Y?K0Ԃf�ܗ[eʴ��Whف[�oBsckk�VP��� `:o�e����EVCb��2I�'
G���c[˵�!MP"��f��ĕ{���i'����d1�Bi�����Y͚�y$�Z8�e=CC6�Լ�e�5�N�5�	�UM�6��1i���Qv,d
�h-��H��V�8[*:�_)�w�(�adY7��C2�G	��]���N*ە�`QՃj�؆�V�@�uFp�֣2X!�c�3�/�N(�L�����{�Ä�Pf埬�V�K/�.�V�lh14�d��෥Sz>I���/vQb����R]�':��Fɹ�r���z�H�!��l�ܴL4O�e�1b�61�vV6�y�cњ3+%6)�b����i��E�B3("rX���q�ܬ�mY�;�A�*n ��R���+bZE��v��YE�R�6n*WJKݺT*ۓm̺�݂n��Un<9g���#�a��f��^FM��Y�jlP���oLA�X��*�VU(�`�W�l��7M�N��,A�S6��b�߲"ɭ6ѭۡVې��4��C��L�j��e�rm�ȅQ�Y���Q_�&�5l2�	�f��f�S-S{a	�D�M��X�u/LE=5��Uz-�b&���4sJ�qcJ���e� %�p�l��yX���`�[��,ӫm˷2;ֵ�F��6�:4���IJ�W� ��ApT�Q�B�M4������*�k���ѹ`̠�Sm�&m���V�X��(7oX�d�u����յV����b�U�4P�mJ�5jP�b�l\�&{X,��6R�)�[�S`R��l�ݩ������d��Kr��7Pfh7���Did2�兗&���{�ITUn]ؽ���1��oP�u�̉v�ve�#�0݉,Egr;ӺqJ�/�[���Mj��*�GM�,�@C���f������s,m�t�:"�{,|��l\�*"��b�n�*vZ/
�o)��ߵke��Z�8Ve��%�`
����M�S6 nŖ�n����F(h�N�����:�j�쵥�
;���pkǒݍ��RW���[[�В�u 8.����l�Dh;�6��(P�]��[�����K(���<���@���G3j�|fսU����b�kYc�qmJ�L=DF�X����i�Z����9z��i�H�%�\��37aٴ�l��<[��m��r§�hwKf�D)6F��H�-2խ�����R˸E<�8m�A2�F�ݽ��f�8��VT��rnV\&�ۭ�W�j�HF'l�.��PDLf�zv���÷�K'Aѧ�0/V�e��	�f��#���-��Z��'&�uc�pX�;rG�`-۩傦]��ugo/+q��NF��L�,<�Ձ�b���ѫ1c�^h�)ht�X(iui�m��T�oU<Up��	Ӑ�Z��dVݵ�P;�v+ܫ
e'�J֛tx��m]]f�Sj��A4#h˩�զ�*l]+��Z>�E�Yu
A��K���Ђ�a�BM7��B?�f����u�����t�6E��ŸG<��ՌؐsיW��.ՠ�Q̲��Z���v!���V�4�B�Bqm]�[d�V�C�
X���Ǻܭ��{x%�/`;��ko1�ʲ��ɶA��&"� �F����EGwYB$�St�ڰ�̽�a0����HW�hBN��L�b޽�`h|s
�@[�3ot�/e,��n�2��T7
�����A�vNf5l*�PYi��=؃�u0㤱!yX�O/pI�3v񄣳�e����Y� ��`�iѧU��*L����*��Vl7�D��}e��q��y���v�u�:橸$:F��H�/�d���9B��7R���i���u�j����ȍ�1��lLI��d�Q*��A+�����uX�t��ɳQ�6��[�O`:)c�j��wSm���a�-Hnޒ��M��;Q%D)j���܌n�J�X(:��>Bd�#9��l8�s�
��ar!���D[Y0]�1Y�׷�]�l�G�+��eSͥ,5A��Eu55�5�%- fB)�m�GnX�2�yuh�	�2*�Agf�j؛��34�/��\��U*��q�-=��5�n����5i�/
�r�g�AH0\N)�:SB/a�ݢ%�aZ�t[-�)J[v4]ڽئ�ܒ����$��-�%?�����f�"e=b��maz+&巿#�H�j ���­��[.�4�Wi�)T4�1��S�ȴ=�tj��� ?�g����Nӑ"S�;T��}>�a�����f�m��Z���4*oc�ٍ1�`�r�5�0'��-U�B�mC�>�Wu�8I6J����NXT��Û����M�`�s�AX"���Պ(�H������g뢸�'H�-w]����P�L��r����
qE�S�%ZoCL:͆�'��4������]��م�ư6GX33,�a��_a���7�Z���p�.�Hn�f��G��:�^��gN;E,�_�2�G���Á����fIV�����˒��s�R��z�@Kr�L�g�}�$�R[\�<r��-�+�X�����<�e�6ʵ��ӂ�$sliy"���`b��IS9<����5�`��<y���
�����{LK��V�s���\���/1-���q.�
��8V#�%p�{�$�\�u��sq��˦2���_]��Z�.�Y+�&����T7�ǋj��Ő�E�)�y���heu��;Q.� ּ��5�P��\�ԫ:�Z�V��u����o�
�s�)a���Kx`��0t���9-����73������r�sxQ���J{��)�j)J��9�iz��,U��mi��'�I�<���fdVn������N�֛� U}f������4����t� ��_-8S�o1��������P�[ׇ4�I�����t���PbC���)�/��c��9BW�uC�W�dRck��ˎcu)��CG,4�I�+CO_;�7L�-0q�x��Un۾r���.��"��ا:r�sr����w�8ĲL�ݎEC��X��f\)�׋O]oNI��GQ0V
��:�Y��u��ĹTA�C����F�J��F�J�c�`ŶYvr�����흥�eѼ�,��.s,-��j�u���=�¹�<G`<�ի!���M��$�T&fcn�	Vɳ�����_q���#4���
��V-��M]����n���������Ιo
;(VޣN�����[�^�N9f�����v��w���	��{t��4��eV�<�e2Ĉ--��f-����aW���^�p���<_n"W�쇜����C��g�R�R{��˽��8�]/�v�`�T��u�ӳ��ݢ�W9J�6�U�Q�c;�f=��{7U�]���������v��Ue����0L��ξ�B�p��*��:/4ޝq�̆k���n�j�bF� D��>t���HI���6�vk���]�F�N�a�R��0l!{�A�B���bw��"S�Ҝ�4�R�Hyd��ǇI϶�vU���v�"-�-���x�M9�`'f�H�?�Sb�N.c�1�r��s�ݶkt������Fq(�\[:7���F{C���M��_�ۢF�v'yu��Y���C1��:(ʗ�3+k�����re39���\C�N���چ�uv�bvTh�E��,7U+[���!'[��E�{�Si�j�A�i_M\9�ܘ�<7�3�f,�-�/�y��/��J�Z+q��j�m^Q���/�{4שּׂ��Y�ꜵ0��o���U3>\V]����+�u��&��T��*����"��T��gh�!W:#y��m�����]t�M�0�M�z��`ڵ�r򝊽�%6��!��d�u4���;����N֌-Z�Ʈ���e|�a���������_a���!�T�Ƴ!vp�x���'j>�ڄ�W�ìB�Yȯ� :���ސeA�i[
―���B��I�J(�Қ���iњ���b��;��5�7Q��,���*#T+��{C���t%p�*�1��A�-WӔd�R*����K7Z�ohb�5����3u��4޺酒MD���ko8-�&��or.�ha��Ej;�v�nS��+c�X�[8�.�%Ō	[|�lWA]ה���A>��:�j}YB:�S#�dΥ�aDvj����t)a��8���F,R�1GL�C4rëKλ�U�K��pZF��Y�&���Vlw�Y
t��j���І:��p#�d}c�Hfb�|/�	}-<뜥�|/Ǵ���0�@�������tgZ�nC��vTg�����gf��C�_Fz*��<��5����V��͐�e��p'T��27>�|5e�Y��m�7�}�Vrk����=&��<x����aOjM���*��\�G*�l��t{*Pm�<���9���6&X��&s��A;w�L�����+�i�TNS�7�{1���bD#$�yi��)O���,�s%2 ���ϯ� vm�6c���;tHki���"1�X�'9�f��K������3bk�v3CC��/K��]��,�n���Œ"{��Ŏ��u۱�9p7W���"ob��G9A���.B�lϓ�N)������3R哵�LYPǷ���}{�_"L�x/`��F�����v�s��]o7�_t���`��Z���\���F�CX&t���/�l�y4uiu�Y�R��A��j�Wkܐ�z&�<�n�w����r�!��
���>}2f�f�jY�oP����I!'�(��Or�������]�|����BN��J�:@Δz��-� ��ˬz��`�u���2�:���	Y���0�:̮�W��� �v�J�k�k��3X,Uf�]�:YC���C���u�C-q|z�8,��X�V 8��{v-Ȼ�������;8 �$�.�s�&_$���m�R>O"�4S�:��ĉ��&+<�v��EOGuF�Q+ySޡ�]�'��R��-��\U>�vm9�e��NfPG�EQT��N���@ ���B�����䄐�Cy�!����t�
���3�g)R�UU��WRe��d�Xgy, ���Ko�}��P�RV�D�K��e�wmRC]��6^يmh>�,!yŜ0\���_�Ӭ�cG@�Uӄ:+FR������������+����E�N�ݚO*��6�<���B�	i���d�,}"�1�DLWʮ�c7*m}zSs�{(����xm:f����s6�ј�q�4Ӳ�VLd^��a[��PH��2�b���}k.���i�9��]hPV�O�8�s���d��[�:E<�-4����ޛ�u��GJ��jR}��r�V��j�H�3f��µt����0sa��pCjM{a�-Z�	ngVN�A�wVy��k����Ȃ\�J���]ޔyZ��0�&����.8.�3�(e�����k:P:�Z�Re<:3;�?I�;ѡ��Ĉ87$uN*ֵcT]�!�U�ָ�,��4	ѕ4M1��&B;�kJ��yy��n"+�Y��./���I{bLk��+�~�8�T�|����*m=j!��{&`�gb��]iB��ݠ�����]Zmc���i�cw-C��?�%OXz7����7�b�x�6]�X{�M��R��Σ��F�ɫ"o��
�5��7��ƺM�M�6%�E����˓
N���]�/�y9�Fod��r#B��go,�ƶ�jv�5�:e�$Qϵ��_l4F]��q�3ٵ�қ����c�]�%�t�)1ܭK*�n��w;�6Ho͋ ̐c�fȭ��L�btf�#�68Ԣp���jo��]F��jp�s��`̅�侾���̬�N����CR��㵅n�f����fޥV�=�`���[���@m�'
�uwv��uc��c�WƉb��;5e�m̹F�L�ðS�ٻӮ���Y����ߥ\��̽��iAHM�%�C��SUU�f�ʥ�;��g6��a%{>`���R�>��u�Voi���g%����wk'�;��{��=/j�������D+\R��VpM�|v�D�g9�B��?-���4%�K%j٠�;rf���"P��=�0�6�`��j��g>'4W�wCf��u0��{�V��}*��\�����Zծ���Ց����}���(ƏV_0�7�z���&�^M��D�M9+5�ФL��w��X��a�1t�2�]%n���)���Uހz�`�
T�_uۅ.��TY�M��6t]�$$VYT��hN�b��H�/@)T�}�-��9mF�t"��6�*��<��\��ӚAڶ����X��Q��ٶ+x*��.���.g4�lC0�:󶌇���g����ؼ4���7��wq>����N��������/��@{�U!�|a���l0rTT���,��;eX����u�BӚmq��FW��<�C��[�4���8������"�h��������������
��7W3�Wq�qW��5�)p�[8�-E%5��na��&b
87�^���,X�u�t�u`��BX���1{����u	��q�F��.�E��wE��h���df"8N4�=I�X��&��8��f7zE�אLz����oT�Ӛ޻��ff�[י1Ky���,:����{�2�֙��GYY U��0n>��]}ӷ�x�-�!��QӰ��j6N��DS��B�n*��]evI��Z�#9�I�:��{��I2Q��V)�]�2m��k�A�xp蔻�!�n��uM."�>�4/���xK����р�\�wRm�3+�V���&:�/U.�M���sKX�^��=���,�h�ۺ'OK���l]kY\eN���`2%���S��0�j�6)�\L�h<8��[�j��ַ��ң�Q���;
9����l��u���U��t���0��Vl}�.�oC��"0s|̜u�IiN��n*���F�����cy,�g�ն���	�㭯���X;�_���.>'��X�b�LӾb,�ӝ��"�wÙJ��.��U�ff�e��j&��Q�҅+ǂ�-��u�v�ih|R"[���Ԝmf�S!�}�U���g����橗�z���>�6K6bsl�[�M�4��1�d�LM�z�P"�V�snL��ܝJ���v�:�p������̡�"�-�.��Q,� �!�ħd<�����f�����u)g�*\Һ�,'e�O6�⫊٧�]
4iШ�L���m�����p#[D�97GT2���,k5Wvf\�]`?��#� ��fǕb�'a�!��7����]����td7����\ݜ�#�Kd�\7xS�u�n��2}܏Co��+m��z�p�V$��ݢ��e�j�yH�k�]�PW�y�A�$���_>G�{Mi��*�(�%�d�ʛ�@�����Yim�=D��vò#譭e�/�'ס�t5��]�����0����:	�8t��ޓWJ�K�y\^q6���+7[�N�6-�۸��Lɜ��Uv��gk|�G4��gR�$=�p��t�����㻆��\f���Ĝ�u����<�����R���wa�m��������?gn�ڮeC�����]#{P�`�Is�(Hŋ�Ԧ辪�+|��82�R�̱�vo.]�ur�sY�oq>�c�����z��`�)�RBgE��iތa�I�шv�ç:��Tn�<�{8����f�a
�����v>��L��3��N�s~���I	$E���D��O�؈?�����o��\=�")�o�Ղ�n��hPyj�H�����5u�5%����jI"ͼBkY��ݽ��.�'j[�.�HZ��s+�3(u͜�c�b,�[q���v�0��;-vRiu]�K���૗qk/������ݽ�l���J�VG�fd}o��ݼ�38�]o���wuƅγ�6wt�VVe�*�HcƳ�a���;��I��2�U�������Fm��d2����.
���3u_�F|�n���v�f�m	w��ֈi~��6
|��x�j�9�I�������N���:�]�l��@!��d\)��z��w6%7.�ˢ�˿��}r�����e���A��kjҝ��n.��՚����嬮\�QMxګP��+�mے��Aj����f�f��L���.1��i0L�Q55�B�F ��!0�	H��Q��@A#�A�cDw3tx�`��i�naj�C�-Kl8˖��T�H亚�-Jk��"--D�13i�Z�[k�v�`�U�l�c�`kD1�;�E�\m���cR�\�e�G+�+�i��`3˅�%�mq�U�L1@@��$��|0>7_��;�\��V������y�k�o��\������.x�q�!�d��Whr�vG��u�ٛ���ԧ��6ˏj���?.�7��;`q]KdBw��0Մ�:�1|�Ǹ9�y����c�p��{�7K�G�	��H{�ג;�Y[}�Q�ݽu���܈�sL��հkvC��h��$=Y����~[9��Ͼ{�V��m��ᰗN�⬮y8�S7�oTFf��}ݫ!��k)d���+��J�Y���$o�B�۱�����؄!'vdh�eλ�]EP�ή=��ʡ gsZ�k.5]�w0\��)��������R7�J�=:�m�����VtB��3n�j%�n�(����������⛧������ֽ�\:]N�#��XWE�a�6���Bo�hm�B�K��՛�$�:��u�\��Z��X�ߺ��[�P�}�u�Z�2i�[t���n&BIr�I�u��x���w�Zϋ�����Kz� �c�hF�66;{���w�dKbQCq��+˩lǔ=���Kx������J�bht^w�=΅Oݔ�HI�+~��r��xS"��ē���A��Y1��<���w�Udx��}�i��g��.���rѧ����.�ʩx:�T+��Wh�u����ݞB�.X�˙ǆw�\����([*�"�GR�����/�=tf!��%�k��<�5�o�pzō��
����"o�B�x���j�f�Z�T hZ&,�I���%bC�}1)���jl͡�����}~B�p-"^{���ϴ���8�s�*�h����ƅ�p���*�Ő2����A��J�@����������ɜخ��=]N�݌���:K󋷄pHl������j�7%�@�Ok>�|��ɑ^��JX��5�s08"=;\'�Է��n�U�/@�n����� ��1$4'2�#�!�Ɂ�z�lu�荃�Cx4a�0Ý�zŌe�yCv��T��ל%�3Gp�&|�b��<�E�󮽎u�_�}�1�b;�Yy$��� W7��gW<����2c}����t���5h���NS;I?3�0C"�#�6���ݏM�7�aĸ;���}����RuikC����cw��u���0����(Otb+=��Z���qUѡ̓;V�2]�C���=|�v�m�;kG͔��ίLL4��/^��t4�{s����X���c63�잴�RT�Ws��4R���#�f
���-�F��%��e��;6��Ty�pSᣅWt&Q�q��8^���_
�][�a59�]�2u\�B��7�3��b�/'K�l76����ǅ)�u,���]S�;�G!�ޕ�;%�o�?Q3�.Ů�X�s�����\Tޣse��z�eݳ^�����Lfv������L��OY�\a1��Ϳ����vx}�Jݯf�h�S�J�v�<2�X��dԭ�{�2�b�^P�x�y]�t�@�P����r�!Q�]
�s�/R��c�qwѽ��<�/}Oo+=�>L�3ݥq�����T��^U���-֭�=���_V����1�K��)M����j���Yt����`���j��BM�t5�s\�5�v�/JW0�k9��Z�z��[P&�=�l��هז:�Oa��bo-��0�<;b�N�\��wP]�V`��Dr�A�R���;�}6c�O���mu@5Ȼ�����Ut��|r4N#ܘ+^l潌muo=��;��}���7"�ϗ<s�Q�x�9����)��kt�:w�D�H���nQ٤d�\���lH��Uݞ'er��JCfX�qL����gr�m]��+y����1y/;4������rg���^UϹ��V�T47*���+-4�UwM� �b�Z��B�y��}Ձj{n�\��[	�.[{���勨̰�G&�vW30!�a�]�����8aN�Q7Q�0�^��-�=:&��R�v*m���桑vN��*����Yq3�E5Igp��֟�=�RUSB�wݼwA�W�nvf�<J�
@t�T����g:�e��UP縯oF�S
s��ph��ө���]�:�(��h���~����C�H�f�)m�XW�t����z���ǒ���&`��d��J�-�m44K[gf�:8;4����+���G�%J��֑I
�
�V�����1������_W\gJy2�{%p�Ůһ#n �N!��J��99S+�+���b7�l�YٷLwER�tT���`U�����!�v���і���<��0G��2�I����\�.���h��e9:2�:��,�l٠^eN�eܯ��]q%%wT�{X����ٺ�r�t����-`v8[<��eʉG}�w��k%%X�����|#�&�rb��ù.�͐R:�ı]�0���l��c�U��!7���*�LI��:I�I��UM!A� M�6�I*��}���4m��>XT��,����N^BdXZ�me24��e*VΘ�^��cY�EգqK�T�:�%,�q�1�V���0��ܪ���UxK�i��o R�Xr�t�i[t�U6�7IC�i,�2�[��I��)�P�A�d�ETn��˹Bn�Ti"N��(�Ÿ�2�.��С�F�Z
fɢ�f��M߼�����	�!F��b��Kw��Ve�n�-1
�7��3S2ݢ�11���nQ�d�%�c��uĦ��s������TZј���"���1��aU�V��*֗��-˸2�H��eLq�l�KkYX�3i�q��܍�VR�]B������J�d�q*.�*:ڂ�ˌ1.6��Q�֠�L��Dv�KK�Sr��1�?J$ƌP����V~��٘�	�j���nq��o�.��]w�[Cg^Wo^ޒ�n���cF���@��*��м!<v���V\�9}BiT5g��՟nz��_]%9Wﴥ�#�-c�ד�a������C3�^Y�s���8�!l�#�,<F��4^�CQӈ�[���� �c���<F��U�"���4����$�Ml>Y}{�v9�޲|��Y�u�HwTS1~'�@8����ʇhL� ��`��p`f�]rU�q�C��-Ǔ�1J��WY���C�j�>�,��B�;��=%et����,�zaXy"�d2��L}3|��`dW�!�bI�wn�5�m�\f��i�!^�̸sݟ*e�[ےP;����6��<0u��pm;�q��P�fC*����N�����Vf�^�T�b26+)��u�������5�w�~VR�qNJ�y&�����{y�9ӻV�?nU,�DM���q8���8XjsLS�#����L�7�G�~��@8a&P�@�O�P��|�>y琝�3�!�H|a�'�d������2,$�+5��I�I�}�ϟ3�7�<�Hx$� �$��zȰϔ�� �����I'�/<�y�gG��<LI�1$9a�"�r�v��� z��Hx�2h�9a8���{��:㟄��1��d�C��x�ā��!�N�|H���]��X�v��<��r�:`t�rŐ>$��a=I@��Œ��5!�!��o��@������!�!��I;I9d� �	�"��=B0��]��^{�5 t����&�>2i�$<g	�@��PIRI��Hz&��>>Yn𒜫aW�5+X�=#h�%����͑K�(��2"VH��̴8�3��+��6���#���w�,��!��@��	���RC��,%��l!��}y�G�|>y�}�C�I5'H���:CY'��C�):`�C�Xq� �N��$��T���!� �8���� g�� �!���/_<���@��� �d��r�� �$��9d;M���0� ީ ����<��>H��6Hp��d�c'l�Xb@�'���!�D!�ԓ��ӏ�<i�<�/�|��=d=/8Hc8B>�p�pya8@��	<B�9I;`y�n޸�:�;gI���zΐ�05$��O�I��>|��e�}��v�
���e��О�$�z�y�!�RJ�k';�ι��<���bj1�1=�=I'����|�C����$�x���s��yRO;��ᄛ��!
����ā�X�t�x�=`޺�߉5��8G����v&���5{η���I�z�C�3������z(��أ6�>�
�n�b�׃�y.����t�>��{����!ϖHjBk �	�	a�dB�����0ή��\w�������ԇHg6Hz�!��C�����`�9dY$�s���=��b@凉����	�@�N�"��;a>X'�CO,���M�� ����_9��z�$�휲v�o6C�'_,��|C�H=SXC����k'�7��z�x�p�<I��B2�v��RNl�hj�@;I��MHg�H_>y�u�sϞ�a��(�����r��>2CP�I3��C�!�9����}w�o���V��|I�E ��!���x��r�ϴ;H��O|����=��=`y>Y!y�����$� ���C�,���0�$=aY��{v��I;���	Ƕ@�=I���9�EET{'�s���-��u���	ϫ�9�5�F��x��Ќ+}����AI���f.�1Ն�k>姨*�)ӯޠ�:Ċ9�+��NQ���,�*�I~��w�	Uq��Gƥga���iQ��\�Y�}��Lr�ݽ��*a=v}W�5`�tv0��#k/M�ī�%��r�_����e��8݃Xν3�y��dJ�7)��ʁ�َ��Ð:��M��7v�p�v��X�d�����OY�;ݭ��9U7=�9��滱a��E��n���f2�w:a����lŌ�&h�d79ї�|J��{��{��r����o��èf��&�ŅQ �X���{�E�sjT����Xoio�E�U^lq�k��2�:�R,Ԁ��ZKZb�3DF�,��Mf�'ט��+'���y��܉�q����̉ɶO{�y#E��I�K%�e�����C�C��oh&~��SOpwv����M������|���G.��?7���]J��j��rm�� �B�f���K?=��5��_�n�S��Z����Yxs5���Lm��k2k�[��}�^-�W�E�<{�]�e�zP�uWM�י��=P���6�D|�ŏG���˂��F�E��ػ#ǧE;��{'xf�8��<qi3��U�V��K�(LE�qV�I�0���C/ސ�.��y�$O��h�U6]�V�l�X�d�w�ĸJPߧ��Ԧ�_��gQ�s4�ѽ����f��W��_D{��\S	��v�=x��{;*�н��V���|�pO˰rZ�Cr��P�|��7аZ̧�;qF�S�Fևz�s=�Xf�d�O^ڻw*�tYǝܕ3\�)���z�.׏;Σ�=+;l�����1W�d[l�3�iYe�1��ӬlL����^��2�Z��@5)��'�׵�����{�7�yK	ZFK��tܖwC_����	�X�����j��z=�h6�_�*a��@����£6�]�l��X�^�b'�W���/XFX�S�����s�2����ܶ����m��.EY�?W��;��q�j��V��e�ӎԸ��!;̅1Fj`u�u�Z����4�ѹW�9�Ƥ�滄N�vc���H�QC�F<��9�o�zo4����ȣ��h�W^����=o*�Eu�p:4Ce]P�!t��IKN���W�oA�F4�%���s�K�{fpR��O��@��5�����M�2mjN;��Upɫ�Zޤ��J�D�Wj�w��W4��q
Ǚ�a���+�VͩA���Su,�;Vp�#��FP�}Y�\��GH�K793��-��eJ��䙷�Dm�ش���ܖ�g[�ӊ�K�������>�]I�zQF�q3��Efq�C8����\�WBӴ�J�p�N,q��ق	ŉj��x�	K��g ���|,`���}qZ#3,jTҦ�f�5y{z�U� �恍�L��"�xЬ�yupH�1�%���J���j��8JJF���E�n&�0���*a(J�yHLK#��#�-IT	��L&M�Y�%`g��ࠬU�7`j�a;(iݦ)�d�FZ����CEf<*��w18�y|�C��ݷ�˘�
��<VH�1-��F���`� �-Į��C`�/�q�l��Ky�R�m���2�60�e��FB
̘dn����:A���7��* �"_��}ZV�UPQEEYk���De�UT�-F�iu�ml�Vکn5&#�pc�nB��2�-�bV�m�ʥ�[
 �a�r��m��ڻ��.�"��*��k�ն�Jm��KMːD����mը�iEU���XYn8*���l��mU�W
(�[�7U]i�R(W�f\J9J����X�[K�T@�����u�_�;����$gQ����ܒ���ȴ�nja+S������������u+��$���\�@�g���8];�X�~��bj�/h�M�^�P�q�}�,�<���;�$r8IU�Vo(�g�u�>p@�	�xkA�o)�*E�7z�n�_<��m�f�h㑄d�ݭ�&8�Fq�w��I�#�������{$-�Z��*�͜�d[�y�HeƎ��9�r9h,�^�競��������X4�6�L����z=�p�Ӄmm��ً
���~�'��)������;f^"A�"�FLj��a��M�o+����Z1�Έ��(�mNG
��}�v��3!O�=7�ʼ���7�N���Z�%�|\�ˑ��P���r�V��A�:�z���,�5�<��N�u���}u��6���-xX3=�A';�u��b
�I�;��7ܮ�<w<[}]������ܤru+�]Ϻ������}����|�ߝe�q�hz��O��Ԇ�);S8��^�N�C��ßT��Ɩ0�6Y��`Q�L�b��p2�Q�.����u�J!غv�{���>�dK@�]la~ZY�K0�;]����<۔إ���,��-۱ٕ�*vz�h{��Ub�8�ٳ�vä�C�`���Q���T��ᴴ�4|t��
,�Ȅ{P�,��/�z1p[^!�Z�����[;��F�{G�o�4l���H�`4|F�l�U����ԷV�ACe�i��/���"'Ʋ��ʁ�}zc~�ڧ�ճ&I��=����N:naʪ�09ͨ�����9d��f7��&#�p�Gbv��kL�2�Fe��8�G����nY��2�
�e_���Q�c�º��фE�H�t�f������U&vr� *۟/&_+5hPH��1����lM�umQ�CثW��qٞ�.0��ڪ�V�h��Pz���\��TX"�?q*q�w�*�b�#Svt�����%��k�O�1·ޮ�O�Qa���֚!��4a�!{�����4o0�?69|�
5K�Z���e�Uԣ�Oe�7��7C�J��W��T�p�|TQ��Y����s����;����x�qY�Cn�q!���W7�3���&���[��=� � ��`���}����t��/����YȄ��9Y.���� � �!h\K�8��K�W�G�w�V@w��h�gHG���������Z�����%��^ڼ�"�e
���5�����Q�c�G��;HTTV�w��۬"����<��A�x�6M!䅟L�Z{7�;���Ȭ��_g�rG��!$x��%Vt�(�Ҙg���RT�va�v�A(;�޺��D��Ĵ��Y�=hQ�bA�Q�N��0�w��P������)*�"j��w�f�o6j��V{�(��Z�y6�Aȍ���'ٽ��|>��{� ~2��D~���ߎ����(=�w���G�QĄhc
�ܓ�D �X��sp����û_��d�fyiF��Z��h+"��E6�{(lTj�����8~�XF��=ٱE*���:G$=<�?"�x飄y�����Iz||C,������آ/U}�v�+����4}���x��d����g�ޛ�����L������"��=9�Uvߥ��|j&5Q@DU<
�<�.��jh�]�>�J�ا@a��ˣ4��B�Ѷ�Y���ɭ�d��dny)��f��u)͊J�;;�"Q�]m,4��"�ʪ��C�T2M�Ɍu��1����{qp�V�&!��=U��#���x��G��.����.��0n׬p�`�<`#5V@�ʄHп]#N`.���׼n� ��/��f�4Y��ֆ������,j���$ih��آ0�������ZG��dAj�����m>:}<n���M^���]@�{qӑ'+f��1
4P�v�{���
z�5��KV~�![�>��j/���.`_4���%!�↭,�%��[=���1�u������6t���b���D^-�8;U̙�S'��b��x�Pk��k�y��_R�r; ��+(/g:���ӇV�r��n�r]ZO�5��阍��Iu�Dz=�q��"����Ӳ��a�����`�+�I޺&��(�!9aCp1�����uV�Y+2�����Z����5\S�Q�0�"�A������d��T�L�Ij�MGd�>!�e��{ag!�$�0�>9��%{X�\�w�o�+�z���H�
���j8uă���TBZ�+��g�,�#H��ζ-���z��C4L�/=K�x�$)�f�0��f��b�t�����n|�&f���$��b�����@m.2��9q���N�8���`��o��=b
�vIL�;�A�͇Y3$�F�gto0e~�>�d��tG�/�eS)�����ȇ�k���nO���7`�/����Ԭ���.�)A�l��,�Di�A���b��Ȳ�Y�~{Y��7eBD����(���]�M���;�cM�X�F�9�.��{u,sA���C��ZA���xBNR�4�~ٌgy<0��|<��ѳ���<Ɨ�I�&��yq��i��:�����2�?a�ӄx����[�l�T�u���x������^4F����;���.#��~ AhQ`�_!��,��r�S!�M��Jgl�����py�Νɸ������p�mA�3�R�Y����+��}� ����J~U�>٩s�UEN�W�F�L�;�p���uCN�5���,�HC�I��,���Š��W���z�U>�w~\8D�M�g�ׄ���91]�j*\����lT�&!�ur䟽m�:a����ͻܛ�������HB2*!�3gb3��/�WC�v���M�x�F��k!���ζvm�E͜�bv�7�+���s�Vm]j�F�6{��*�r�g�yש׆��l�C���\Yp��}ld�� ��	�]w?L���=�zIv&��Ʒ�m����U��B��#�D�n�hI�׀�2tΣ��S4j�Tn�w+��ճc��S1J���������μ'p�,.�ꯨYܭ5Vi�����A�]5��r6��ܲ��oo2N�0�	�6d4w�����J�N��a���L�/$��ٜ��<�ـfa����-���.s�g��e�H�X�.�ԖNn���M�P,mw�{+�%�S�f�s�s�Hn��%�:���9ҹ�Sw)��^�unϫ G��K�g"�>�}��am2S�a�ftV�M��I��|5�����5���S7�7��C!�w�&���!��7�H��-��Lb�Xj��!�*w�.YDܗT�1�¥���w4cv��I�i��Wvv��J�]H�ʩ�F�F.�Q2ڔ�G�F]�*J����9or�)�v~9CGb�AÃu���\IP�)�
�m�c�T4�`Y Q��`,QR�ҵ���_;��@�]�9�&`���I3(ٱ2�R��W����z��)�,�TU�11A�V�1���q�n�TX11��[�E��(�5���eUU`������"#���fR�DB�nd(V*�e�2���0cEY-*�[V6�R�fS2���G(Tu[`��e���Tq��i�������uo=���Ox➻W���Uszj��~��G��Mwמy�v�_[��暜&�w<u�[��Ț|��垼��?
��!dt��H�t�x=;kC�"�X�8��Mi���hSCR�lئ��b�{j}��#��֍{������0�Gg׬��*����tܮ��^��h�,�3<��_,���������Zoj�4�W�1؇7x�ҬTt��֜5�VC�a�4���i���v��]Ktwܠ��89CF�$��#UH,ש����VP7]�]��(];���G�b�DX����hڐn�^+��{w΢�q��&��*����Y�iйoA��4u�uE�:�\�Wt��K����G��k�]r>����?Z��-��X#���VƯL�cP�(� �Y��T�v?����;�;����4���*Р���8��0�Uij^M�nY�Ԑ�x�_CF���G��<<}o��1�"�D?G��ig�-��uQ�= g<��8��dQ�	dVa�y�Ϫ�#H������i8�j��D8E�Ce%����V��+q��/$��;r�z�������]��G�Q$)�#f�XI�C	�=}�/1�!�@�|Y���v��46;z�qҴ�z]b�gif���w��}۹��� �f�H���/��4Q�4�?B<�������ݞ��R��{\�DY�H�f�or��*����l���~{o�92�Y�l$��{^��߻_Q�S�bf!��%:8D>N�>���=O��������4s���4~�}&>��i�����Q��dr�0�5��H�o�=tǏ�?Bϊ?jCְ�[!f��!x�h�����H�C���0���Zy�]�y�k�|FHns�'�r�b�: ȷD\�>5=uz�Y����'�c7�Ck�ۇ�,ϊCݿ'��uzF�*��ۍr��)��a�,���k���c�]z�:�M.�#PI/��z=��~���+�^����v�^���;\5a�ƪW��/��<C�D!�@��,�#㚃�=G�_�#�NP�@��ő^(\´7Qt<�z���W	Hl@Y!:W���{^��Ґ���� �Ǝ�>"��<F'[}}ԷI^ذB4�z�}�q����0+���U��G	�0��4����d=Za�E��z�ze��#yB,����z-�dYh8�>���׬w��Dx��=�a���Ӈii~��}���x��yу͆�ƨ��;_F=7��x��xMo`���ճ�l4��`��Rt����`8K��
]Fq����q�_o��������6��C����XBl�J�amQ�;Xo��{��HB���k/k��M����A�w\��p�~�RB��aԾ�Z�ɭ�jr��c�����>�di�0�I�k�Io��y3�H��?*B�"���U�x��D.����d�G��1C��,�ψ�Ex��enY��װ2,�&����dG]�����3�o���LP"�2k:_��ۛv�$�bqٗ�m!�8�/�a���ۤg�XG��as�g6���J�8P�x+}`�Z3� W@�3M�Ұ#�ӵ[�zt�Uu�L��#!=9VT4Ƽ���gk�]�=�wp��T����*�̝�]`WG5�X2����DG�5���ʚ�8��9*}:g��yP�����n�k%�]K�`�b�vгD3��u���'�a��?u����GŜ�e�J>!b���Mw����/!�y1�x��&��^l6��w�*���6�ޖ�r���9hV���S��}�4��Tl��f|�"ZX6Bt���Y���f�7,u��i¾�>k�2�B����lq~Zg�/_Y$�(C�t~Ć#��_Q����7Ҷ{޲�܇GE�6x��a�A�L�3�~��F��l���9�q�eLPA��ͩ�}mr�n[�];&;VeOC�(6�s�mS��f���e�Ԧ\�?L|r��
�:����q�T��s���B��d�\t��H�eA�
�)�ޫ� ���׈�H�Bm�Ӥ$�=B׌�g��`ُ|�"�.?P0��'�"����>���]{`Yl"��#�~�(O��J�˄{�-���D�"bH",�D����oS0��cmq���qGMv�$�
��US}0�:&�f�_��a�#�t�u�z,���B�6G?eв1��a�d̜����ϱY�Ȋ1qQDsL�jΜ7�9k��T���uF��7���])![#��-D�%��r���]�ڂr�v%���Xrw�}��}�~���e��ެ$�
�
?y!-a`�V���uR~��gǎb#����/�?+J�z}�>�������cg=!�x�D:G4ٕ/�a���8����㘉~��6��7��w��G����(��>"��`�8��q.��G��5a�G��
�!�BZ'�#��z�_m]X��"�/�?#�E"�yq,َT�E^X�\~Ō�<����x4(�0#�yƆ��:l�h
�l�҇��G�n��K�1�G�º�v�����3��'�w��r7�;/D�hli��3�Nҵl݌����׍�Y��}9R�W�M��ԯ=f��b�:������g�0Q'��t�~U�N��1��~��@�l��Up���0!�q�qB(ه"�VG���@��%!�=��4h��C�N��	��z�K�<h�P����l"2D#晳�3�j���xv��B�%��q�e�奵G��;�K���y�(�*=�v�Fj��^�ϼ���h!R�)!s�a��h@N��,���y,b���a�����[a�'�x���HFu�$��e��Sw�g�N*;���!�~�#s�����Lw��õ�]���4�o�R����}x��j�S�"*��uz�B��2&��_G��C[��1�lV��_#å��/�d
&��W��")�0yv-$���ڂ|E�1��Sڳ�}��8�!V�mY�<�}A"r��+������$�>8l��L񜇸����_�hx��+-�����?n!]l^!�8_{��wfu,�C���R�Uw�R�t[��3���mA]r����PѲ�4�X��\��|��dTS�rl��G9Q$",��.��<q��]tQD9hi�n�cؘ�bl3�,�Q��.ՖE������v�pߺL��RR.(��v�eT*�;q�RzqV�J�v���m��lL�0v���:�wm1�$N;ٗ�;9�u�:���]��R�$6$[�N0f�1�H�}eh�%u�.�kw��Tt�q���U�c���5�EV��h�4�r��\h>�F��fh�^˼�.V���p��O��h��ق�U��!�w<���\y�AL[��u�{�uҝskT�ja̎���c[c��H��	���6N6gm.��s�ԍ4�~�2Z�l�<��"Y[M� ��!�t0�^RV��L��'%I����w�r�ơ�5ũ���Kn�_��|��nMn���"��]�;ǎ&2f�D�㴋�׭<���[S���}J���׸Ԥ0nZ��V����cWs���tG���w՟Z��I9���F�Ug7/U��1ѹG�Û*�i�:������E�t���K���q�^�āvnB��Ek�S^�EgZC��F�������Z*Qu�7����<	N]��EW@O]_^u"���>��t�oN]���"��	������C��Uz�ރW�|ﾬ��i�݇�Cx<�	$����_�L˄�&�Z*�n&%'Z^q4mE���������7+x��[�Ș㋅�FҎ���W-K�i�gp±q�hU�\[�����ᚯ	^el��(�˕ƌ�x�2/uݥ]m���Mj�LG*�3*��ʖ�!TejnC.,�kJ84[J'�������ʔz]�:���+e9}'P�ވ���5<�;�x�^������=�8a�-�6���^7���$���ۣ�$2����TH������x����7�Y������(�<Wf���
�>�(�F4$B�f�m�hӅ!n1���o��&��Mx�[#������#�0�9h��3��e1���>[�Uu[;O&�'
0�bB�
kNy;jބԲkP�b�D>/�(G��	������}:��C�|F�TY������z�瞯�\G����=����aH",�J���CV�N�{q�I�銜�N!�u�R�
*	�W�@d�g�:tv�.���U_g�v%�<���g����_�r��e���O���h�H�J�����1�5�ǖ����C�Ϳb8���G�0E#e�u���L��G._�ΑgPdO��خ�\�&Q,G�j��VI���k�HY�D4���[��P�B���x�hP�ΎG�:D~{ce
7��#�])b�zo�i�]k��ħ�g�`�,��%���a����7��'(�v�{w���ՄY��h�!�TO!��MJ�ǕU{V�<׭xـ��qu�G[%�4�<Փ[�ԩ�i�XwEޣč��K���|W7|�{2E�o��:��ȕ��2<���!��z{}���o�/���F���>0�V��Q���y�����<���Ci��M
#����}K�Cb��k�bE�>0��'�ofo��	"�9h_.��Ϙ��4]_���b����H�����?;Ǧ}hMZa�UV���E�Q���}���VF�㠷~���+�����!�L4Yq�՛��t��f�ZX��EҢc�<�m4~��秜JC�LT�=4��"lу��h�Noe��j�!�#L ң~B�X{�ψ��沂.�G,\������o4�*:3��g[aJ�MQ���)�yJƯ\��Pe�����W�N}�v��+"��|E	"�!�X����5��AG��f���G�Hx��aEE�qda�B��iR�;��q	�_j��
B�v�Wz��:5#�o��
�p��.�0�^���R��e�@h���`aӉT^0�6~��K�/����bj�,��ڴ�]��p"f����p�$:��fr��>�4�{]��nw�1x�d(�Y�RQ�;����g����s��̡�<��(�(��ٌ/+.�)ݼ��Xa�ψ�VCmk��B�1�65�~n��Nb���JȘM謖��ۻ��銇O\�N���Z���z$�������x��+���r�(h�Q?�>�|��vγ�G�.A��S����ݙ�����H������sƽ�n6}�P'r�ə��`�ϕ�U�O�3P�bFr
���>)���W���?��d\_�u���% �K��{��{��}�/y!}�v~�C-i����Ţ���V�8Q�<�c���,�q�Oɠ�U�]x�G��6q!����9<Cq����UU0PG��dW!��G�tM�Z�&;6i�����#G��������'j'��*��v�=�E4�ݏ��.��Q�/V��}���y�B{�x��6�̤::6w@�:��Dy���3鯦��u	��(�B�
kW�9SfW_��8�CAA������4{q{����T��6ՙ�ae���<h�#�a�˪��la�����H�<�DQ���.��$24�/�щx�a����gM�I$�w��	$2=��)Y��,����v}�y�g_��U�<`��b��Yt�z��@u�z����F
Z~�"�Y��%`�M�ά�]{�Ѵ�� ���,$�YpE�$�&��k.@�HicU�r1���=ΎG�.a����V��읱J���A�ܷ�ה51M�^M���81��ܙ��f��;I�������#М
Je����EX���nS�t1����ZBj�O!U�=��[z��<@D�f/8E%���kI�������͐!�X�<n��NW�����G�<@Y����n�7�ݎ#�+5�W��9MC��6���])=Ճ1iE��Fj'�D/m� ȣ��S��Y����#^�bGN������Y��/�4�;hYֳ9���_!�Hٛ������H�(�W^��O%�����\��O�[��^�����Y��6Yȋn{����$A`�d5zxd]�#�o��Ch�m^���ɬ�Ӄ0��}Wx�
������G��7��>����댘�P'�>�� �#H8�o�:���<a�^CƍFb������Ҽ�W�mR^q�ʵ	�;B��m����ObY(J#�t�CJȣG�>�2,{U���Ȏvn����Դ�5"��!�Slw�ÿh�m^g�݋�Y�F�͆x�` �E�i�tN4�ꮻ�M�C�3��!��r��}HD�m'�>��;���N<G�3P{�0�1g�]{ʉ{GA�[�<CKJ��TX6s}x��=�v�憑�@i��$ލ{i�"���<���z�g���C�K�X��Ew�\���p�s���J�ü.p�\���Y�/�=��6�a}^�s7&KH�\�6t�x�&��v���O���u�N`��)19-�I��׌H��%�d���r��f�|~�cN��_Vn(]����,/��,!�B!m A���o=i�Ha�U���!��r�PѳM�c�;	�g�a�e�2!����|��%(l�밈gƈl�/��{L��m�(p�z�y#�حU�7�g�S����7�لVwN1m��n��_ij�aD0|�#M�V��Ѥskׂ�X�gH�M��Pמi��z�'ۮї[�<wVKSS.�
�y�UDL�S����w0����z`�c�]��`��lqw�}_y�w��T�9�b'_�*�s�}}:��}P^��S��Z�)��H_�J,Fo%	T�=���p�.~3r�ף����_�+�����I�{��5ټ-�}.�@�"�,'��G�ܱ���oeo�z�M`�%��g>���y�mF�)���_�b���zZۧ��!���^q�]rL'B�n�T	�n��U�GJ�2�D�=;���\6s��*Q��W2/p�����9�U�.�%E��n�����L�S��1�u�ˡ��g6z���2Y�����Zu+���f�$3*iw7Vt^���\�8H!�2�� �TC�S$�k�ջ#k���^:e�o/��������m`�u����}���ܶ�z�`����q.����sm�^�]���T׵ǹ�&�Z��mM�ƨoH��fM��U���L�r��'$��������U�-	�0��R|�fy�%V�u�-觍W�s6��z�N���T��kd����s3�vCƜ͹�C�9�weP}>��dP�V�o�`�b��,�̗������p��B5H����侨pj6I}�v���he�`�]x�E��(�������{Lr�*���ҷ'M)K{wm��!<d9�����(����;�X�{�����2/�5��u��lM:E-B���g>X��V�dh����bކ�SG�����])�gc+�aXD�V�
���E�噥�I���Xv�}˹��4��lU]�O+������ҷ�[1d-�-P��um�A�ySv�H���w6������mV�+Wp!u褺g3n�#��K�kgTŐ�ǧ2-r�EiUL��q���֣[����`Ŷ�R��(���R���8ۙ��2�JQ�*e)��U2�U�!iq)�)��;��Vィ+E��m�-�-f3R̮F.R�eq�+V#��a����av�I��������W�������yw�n����4��1�`};�W�WN����7���;d|p�H�;R+@du�u<���� �������uM�rbG����J𜩇�`��wbݔ���5>T�Y@�<���k;e=��U�1b�Y!�WC#v��F��2;����5͵����7}��M�<U�-k��y�xvl�V�k���r��S�g��.��}�,Qw�;7�-�˖�ڝ�FL�<w��3�2�B�R�oI)r��{ɗwJ��h�83>w�=�Y������î8S�ŏ{������1-9��(s�ei�N}�W����m<�{�\�#4<�!��8>��$!ʞф�*�@�̌B����o�79�U%�ؔ���%������aWD���Gݲ
�Z�N�{l1�u�v&�eι��ϓS�V�O	�3�[jy��qHa��r��B����xv	FU�.�����M�}�������f�d9yǝpq��Z��1$��o_-����bjSW}���x�o>���Q��n��Ie�_J�S�Q��v�R�%���슌�P��ywH��4�xzRi�.��IOe׻s�$�]֭�-��z(�u:̨���;Ig26��#m� #kG��5��RBD����l7}M��Q�՜q9쳞�0i���(gf�z�]zk||���g��q�M�o��ÞY�a��iUL�' |���3����?*���~���=��卧��h�S�~k+�9�{�Efe���ol��ZvK�&(�b�-�����V�=
.�c��+4W��l����f�V�g�����]/캲���������h�o(�U�6���ѐ�|d(s�9����]qtF��.Q���#kG��"r�ԀҊW����|PW~�׽���T�n��㛥�9�ӶU���;v��&pղ�)ZI�B���[XlvZN�u�z���w�}^���&o��]��hg݂��nwy7��"�3;�'�N���7G{�NA\$��l��؎��ˊ�qhu�V��6�s����p̑�[�İ�-�e���V�����X�����Ț��=ڊ�U�ˎ����׭qYR�KХ��B�c�ok�ń��E���ck�]�d�E���s>7���U��bڊ�yI4w^�:�4n�3���?4��ژ��'�~�s���?i�2lK��7��\8q�UI�.�M�ex��Gn�LF7�Ň	��-�.�l�Ҹ+��[�<rfy���Wz7�B�i�J��j��6�__s�ˇ��Ӹ�`�6}'��6So���xne�C5_�/
kh�+�]1�޵K��!X�ٖMm�l��fE~+�ٔx:��0���uə�^*�9S��}	)�p��X�з-˧��p���6n`陳ZY[%F�
��H�R�3B��,���ctyD�^P�	!�DG9i
���S����d�x�)ݰ~ 31`�1W�T���J��{0F$l�;J��0ksգm�j�q(Vs�.6꼧���i�����Y�yWw�}F;�aӼk�WQ�8�UҔ��+p2��&kh��9�V�Zf�U��..hӘ�x��޺�vN�6p&̎�g�ֽ*j��5�7��6C���	���޼Ӵ�c��m)��G
9�H���?+ﾧ��{5(�ߋ8A���KxI���Y���$��f��:y���[�������3!U�/^�J����/ �t-�Y�W6����Cwv.za.�då�˻�P���9��;	��Cʜ���;�u���Ѣ�Okݱau㬩+��!���y����9ܿw{��hF���L�h���bk��NDuWe,��P��,^�,��A2�y���ï\]Xq�q��M�����'�9/�#�c֯� ڊ�Y��7e���Α]d��ϥ����@�x�.���6��(t_7]Y�w���ar�]��X%�P�C��=|8��{js[����)}��X�[��Y�� �^c7�VVt�~�`4/���ܰ�ƱP�_r��;;
��^�;�sx떭��BX�8���L�7쭮�2t��&���Zg�>v!��5��9@�afښ�R�P�!����d��DɌɑع}�G��O��[��Лƪ|o/?��9[x��GI��W�]��+��µ{�N$)��;'���ٝ�6��情���`�������y �k�3�E�7J����L���f�@-b)���[�x�u�v���X�<I��s�<���Z�}6ܐwy�I��b�VJ�u��=���k�<��K7İ�HX=���uB�o32"βqRZC�i�%�/r�NEn��/:����n�^>:�\t�f�����uf�yy'�e��)-E�a�]q�w��3ٷ�}pUɬ�p�KH�E�B�y�P��M�OE��%GV"��s��z�sN��(�(�rv��]'}G�D.�,��ʞJzE,癛8��\��%��m������7�(B5jh�BvZ��Oi��AkNg��sތ����5[�`5$�`n֭($wi�`����/��C��&�+:�UZq�AW}�¡��"m����ʸ.����`���������(rU�#X�͟�y6Y��H��
Wj�:]N��)��`�#�ݴ��Vi,Ӷ�b@ɦՒw*e)�V+]�-�͠��4��i����ʰ��6C�l��F�PE�U�[�Jx�2,�(^-�x��[D���7R�dݱRJ���`5/b]�Ʉ���jU2�Y���T&%@�N:�fS��A���ʎZQ�Hg«ġ�L2fg�'�(�>6mL̫4t0�r͢�̘�Jg62*��N[�N�iն��?��бTE[IX��ޒ�wJ�ʗ2��v�l�-q�Q�̭jň����J��+Y��iq2#-�b�Ɍb�(*�V9n4����bɌ�Y[EV�TX��kDAJ؉���b�
2كr�b�W-�Q�ʩ�E��r4���4T�GXQ
��Q�9�*�ƕA�A1Uߨ�mt�D��7U�3�JX�8�a-s��x�'vωܚ�L�$P����^Ȍ�IM���Dy��K?8�����:��ȱ��۔��=�����uu�z���ܣ(��9hp�"	����L������X�!9��
�۞մ��J�$�ow�!����`D�S�%¾c({���'��6��2g�RZ��x�����𙸶'h�8���
W�t}�	>�2:�4��JM�f�q�eI��Uz�;�w�]G4;3�(
��<���#ж_17}�����=�_g$t�`Z�͑-���vꖏNM)�+�nn��L���J�dY�]���Ž�=|���8��1�WfjXr_�6�d�gxY.�P��l^Af�ի;�K�ɆFk�s��H��H�s0����	�}�;��3�
���8�V��O�پ4{6]^�����(N��z׭�ܫ�mt�L7\��}m�8Ot:g{�e�~ƺbλ�����	R�泹k�z<��|2�L��r݌�?V+&�<���ڕP{��U��P�FK���άЏ`Bvbc����:F��`h���L��6��ޔVk��]ۋ51s��5�Ћ=��bO�VNI��pp���8`�GT5�`{fb�8�<�&����*��ٻ�����K�7pIH�Y�/,�)��~ļ�LR73<�>5k�kˣR��ԫ�7��oa#�_f��J��\D�����p���4Ԣ;�)��S;��v�%���e&��2n>Vv0S�E_�RF�\�U>�j������qgX&�)�sh	�VR�.�}5�eY�ᨓ'
2N	QU֞\����B���c�nT������"�\R��S���P��^P9Q�G�`HT�W�1kT�YwV��*-E����^��<軴Fc|���R]ц4Z�k�r{8x�O�0˙5'Tn�������!���弿V�ɸ�}���j�'B1�'bK�z��/�>ߪ6:�+��^��-ܾ�)h���������w�U��gg��[/�c�Q�.����$u��m��-*�a9�j�;Z.���q�ȸ4ƻ�JC�yU�'N5�r�l��5�����mo(c�G�U�˵ �8����*��饮�i�
�6���8�d�Ù�|�77\�m�|�����~���ī�\�s�(#���t"�o�.����6�yW���V28�7V�ʰ��a2�H��ֶ�X�����jب,����F���Y֮���@r����(ͪ�i��
y���1��2r�Ůr:����Ϲ&m�c��Z3�M�^��GH�'gp�s|�(��9m�0�n�OQlԭ	0��,\Y�����[�c-q���[t���:�����*)�3A��ȅ��%�W�E 71�Bl��Du;R%q�5h'�KGVo͝{}��7p����o����_����#��{@n��$�N�$eAg�/t7�����݃-c�(��љ�R��w:�hQ�����Pߏd����&?7V=1U\�X�{��B.X�#�]�&�=�L^Z������x��"�S��{vŚ����X�=#�F��y�:�d��7���E��%�Z���}U��![�w��j%
Ã�vIh�T�v�ͮ��p�sΆ�Vo�����񷐢�7�ܴ�^
iT������C��;��Ǻ�g˚F��M-��yywzp>�G��M��Y!�㝷�d\=!�Wc��3W��5���?^[P�D�	!��qyL�_=7�3�cԭ�̡t��!��œ�,\k�$3f�V��h,�m���_�K�D�=2S�*��'�R�^�ma�TEur�S�Ե�{7:��Z�^[�K��]P�U�u-�ٍ�q3�m.׆)g¢��M�ü2�k���j��g7�&��',Z��'���]ݣGKI��E��c��,��O�;\��8�̫;n������FO�3sA��7]�5uu�����7���ɚ��o=x`3tq�t��˽�-Ш�J��:6��1�-�$�먳�����:���n�Ε���]�zEw*�2�QR;��.�������#��s�u��V�.�c��͵`�x��%��_h�8�#m�w��Ͳ�3�ج\7u(�'�.>�������E;�X*����Y��z�ͫ�[Rd=�Ą����j-��|��^+��{�K�^�uk�̣��W#��J\�;�L�r�;{= ^�Z�.�V��4'�mr��Mɻ�2@�)��~�ރmGc�7���8#�o�.�0�T;o�;���&ݗ9��d��#P!}Y0CO�7ι�h�^��r�:�	�vY]��39�Z���-�����+��p�Va"v��"��o%s�t���p<��P4hs�Db6��"�nt]9���4G���b�B�'7y�!*����Ř;&֢AVn��/z^b0Z��Y�ܞ�kp��S�����pi�J����g���Q[��<D:��^^��e��+wevWe�̶�݇�����y�*l"�&���7��'}��� �;i4�|7�m�z'\��e+�4��sjXW�7E��5e�6԰�N�M3CǺ�y�v�0�I��40�eb��'/(���*`Kr�
EKe̻H8�&!�Tyl��rPP��L6���eJ�ю�U�
M�c�_Y�+�X1������x���T�L252����fT���2 �ˠA�A�[���*�o(<�E���p�q�FȠE�0"�6+�g(�Hdwh̼��,ZNL(�M!�T���f�L4H"rTɐ�b�H�l�q( �̱b�X�K*���,�'m�.ڎ���yy˶����,ĭK�e幞]��ьU�W��QX���r�.5K��\�1�G*��SF��#��6�b4���J�������k��%���\rk]�lܙ�q�jZe12ت��m��a�[-��SL�Z���aF�m�Tb�;hͫ��W�K��-1iRҢ�nX��#3.3Z�.���sR�RA��"���?X��wUe8M6��� =(�M)Wa��t����%�;]'F�{��88R�f��s'*{��b��\ws�}���3J�15��6i�=6�m�[iҮ�[]��T���m�y��k����P".&7��e�q VMD��tgsdX.��ת�w7Ǻ�`f(�2���P ���V�"������pӱ�e5��0W1 Ԓ�1f���ؑ�W�R����E)��wp��h����ww]�Sw"�ϒ�M�ٜ3:�{I>�����b�(t~Y3Iv�s��ox�G�ECE��ŧ
��N�َ��
@5�w�go�f*2zu#<�kP[���X��mzJ[��l[Up��{���aо��վA'@ތ��fu��R�;&��gT�ق)v1ҷpgY�|\\�����˷ҥT�Y�w����ն�C�6|���!ܭHde�Yڒ�J�A��4�o�WkY�w���T��&�}��6����!����-k3=˜\=R��Aޤ�~��
�8_#�ū=�&�������B�^{M�X"�+�h積^�aR��8]i�O��*�6kw�
o�������4�^���5eM��2�xa'[f�͏֢�|�fg��ۍ�O_��{Q̇�m,�y�������輗wϯ(s�� s�;����ľ�רV�Z&�m8�;8v�����u`?cC��бgw+�v<Ϋ�ÓԦM��`}�;��'ՖF�u�bA)��C��.��ǒa��7+�of*A+��҂�7G�/0d���7>^x������k�ֱ�?�Qg6���$4�8]���?�z��~p�맂�o~��8�ټ�Rk(K�����Ϗ)x`�##y2.�Ù�kH�^�f�z,8��e���'��o\����E�I=�O�_V�/4%�E���:��4�g�2�򼈌u�S��e0�N�j�
��]z��g:�s��GVc�c�Z��@�Wa �;�N��MR�U�ܻ�fi�0C�O�ޤ���>�\4�ܴ�D���Yo�ƈ2����wR����\0{6M]�-��q{�L_�)ø���ԢZ�+��e�m5��u�+
d��uν��Zee�y�)��{C��MR��5P��"p9�O���mL��+�ݘ�el�����Lm��M�Rno���`�/{Sn)�l�J]�8yN��徦����Vu���2�y�O����hz����YG� ��F,5S�6Ix-f�S�t�&��=���.�V�ӎĵ�hvs�7����+�7~Pa�P��΁����l�v��.��Q�9�qݭ�b'x�b�c2�/ݚH}�y�c8�tN:��Ҏ�ݮF�Q$N��t>�#��zy�uXzI�xY�W��F���tb� ���ΩҺ��R���C]"��$�4'[�Ӯ%�x�=���oL�a!�x��ٲ��)ΒG�B\�ݚTe��UE۹m���*���pA�����=6'zFq�cC����r�3ʡ���uꛍ��e\�2���K���*WE`�Q�<�հ5�5QR�40g,f��̐�z-�&0-,/3,=x=����=sy�½��>�z��}3����bff�ą�9qh9k�N �YW����j{d�3�uYɼэ�[6j���F@���P��]���T;��EN�S>ǐ���	����f���I%�+$�xY�1�]5ݽ����c���?!�#��^P���x���ӡ��Z����d$ ���
gf3�ή�o��4Wlż�H�����mk������a�C���
��5ȯA�Õ{��Z����k�3L�|q������9�l�ӭ#쥚]���.���R�K�7�|�5���rj�m�6���<��>��J���cP�G'ݛ���EۓX���\�w]���I��QV��Ѣ�7�2ՆC+�3��{F��\�1�����vr�Q�wx�3D��{veݥ�v��U�C�	ˎ0����U�qj��H��i�P�a׫dݡY1B�.�C���cz1��>$�b�{O}a��L7]ȃ���H�����v�Y:O\��׉i�5���є�z�����7�g0%�u�x�HT	J��K74�\��^��J�T,
����Ե�T�9(��s��o4�s��rE����_gzrL(��G�V�!���ӻK��m�$� �S8�$Eo.KG{f��5ȍYg׳MX\�ffe�
�kp�Z/l��r+��oN��f;uro�������=Z��敽�U�}����D��w�y�%�e9WS�q��Z7~+E���lҮ��2s�Q��6/�R��PC�hi�:[S��+�sr��+��wѫ�v�W�d��)r����r�b���:��4�x9��p�a�뭽�R�7�L����>�i<��`wz��Ƶ:eK�����]��x��s�s�JJ���N�J�:`���i^0p|tf���`a�
KWقhI���.�z�q(4�w�b��5�����	��w�i�O@���OU���ᙢ+4���ìl��e-�3uU���b��,�4�vp9�:2"X2�w�۶u��+��W����|SY���y��Kr�`��&��$�D��A�Tq�teH�RH�}u����ϔݼb�C�5hi[icI,�oq���Gv��oLv�gjԗ�x�p�Ʊe�T�l� "�^$h�w�.�2�ɗCY��l]�]"�$�P݃hf�en��+[8�V��5`�_a,�0�2�#�YB;U0)L"I��XM�3vn��2��*L%X���[�[EDV(e̬���2QF�SZ�t���E2�X�c��$E\�%����V�Md��LJ�]�¸�+
��6ض˷�E`�w+R�\�̳(�ss��v�-J��F���R6S%H4dA�I~- 
��jQ6����v�ffj��%���7�m1]�6�[�.�cm�;�
�\hڶ�&�(��6�3��$LF�d�.fcne+�-�ڸ�e�3.��$@f4�`!���- O�3ݓ�;Ä���������ttz��S��7��1�p��:���a	o����:���i��A��V2��ۗn7:a�t�,u��	��ܽ[���}�,���������5��7�{�iy]c/}i.Yz� u/'q.�� v���*�L	7�
����jz{r��)��5�Ȳ�槃�X�!^F}��wڕm���9Gug8��f��u�m��j�RM���b�f�jv`�H^�>����nZO�^��F`����9��ݞn:{wV�/��w3���`ys���׬��g+��H�)����N��5�7�c�*ɲb���M���p|���ܹ�qp���/x]�~<���h`-n�.�#"������Ԫ��KaΪ�N���0@}kE�"�Ӎ����Om˵���u]h�b{�xEMܜ_�����І߼.�w��x�]�i�Յq�r���OM���	�':��n���V׹�����Y2o�����H9u��ź�;�ej�7�^Of)�*���w��Vfcy� B��k՞Vyx���㣐j
�b����^a�;S��J�-�醂��ҥL��s��P^CwX��ǵ�=|�*������
�d��9�d�8�Cަ�S!��sg.��wa`6���Ԕ'Zt��j�Iߙ';o2��U��0>Ӝ�]�׸��쏹��l��C����2u�|����s�g3گ]�l�����#X���b���9��u5�Y�0���!�-�v<�t�:y���f��c��f��\r�a����-�-��Q]�]JDw%�5�Ϸ1�S]`��Xvd�[R7�]��a$�*�Z���]��_3��͜��5��|y!�����sI;N��Ϲ̩�n3+����Y��}��|�B�3J��/�\8�o>��)�=c<�#w�+5Dz��<�gc� 㦉>T�IӋ��,,���$؁���ks3U���5�"�1�}}#��P��{9���k��[ƶ�(����j��;"���ho0-��:O�O¹��y�A������ҫS�fFQ`Ӊ����sNͪy��꘴��L3�xx�{`3�yV��h�%O�yB��pM��)�D!�1x��%���X�hëV��⫝̸z��i�Y\H��aeu^�k�O|r�Qk��:�+s��oX6�eCT�$�4u&�x5�u�W�5��mJ�׵����~�7-�̌�����*����~��|](�v�Y+ի���&$�7}'<7�`ڥ9�)�X�B�q�إA;�?1T�ɇԦVM8��^�����~�ĪCj�`�Qq\d�/h�D�����%p`�O���lh�rL��껍���y9�+�U��u�sZm��ڮ�a�Q��8�����
��u'�w�qoG��P�U�>�Y�V�!��GO$�����G�6��l�33�&�ocR.f-%��eq�<��c�d�ՆPk8ffnY���xD��L�8��Ct�� ݱ�+twx����,bѳ�6]����>I+0��wʁ����?V-�^D�cs7/�ޱ�3�P�z�v7��I,2o>^�az=��0�G��pq������+e-\��]9y!�f���M]G��^���o���nfM���V�ƃi�gv����	�u�L�[<���R���V��OzS:�N;f��K�vQsC�P�ܗ�J�ê�t��<��^ߛ�2��_=�GΛ�-��ϐ��qS�~�b��$��xeb�ڑ�8�{�|�r���ūI�bD�g� 6��@�Y�B<t�߰Է�Q�'�{k����]�wv�J#=���&�`5ʺ]=�=�ێ���zw2��i�n��_���1e�B]/�,S���)�\D��Q����H���N.ףF�g�@a-���^G�����ut:ɧ�������N3����� �,=آ����d$-�p����z�'����~O�f?���Q_ʁ�l�FFu��w�w��ܦ�J�A֒Jum;�oe4h�)��3�1����;F�صڻ�Lr�;��0�޷����s�;���F��q%�;RR����y���(ּ���6���/o5�<�F4��lE�Rt<%v4nʠ�������۞|i�*ŝt�Dd��;I�6+OF���;�x���f��CS5h�$ͩ�����%����T�iD^�Z�{�J�>��Pٷ3�H���W9�ٮ�E�/f�Nj�ϛ3�n%Ƌ�	�W[�qnK6$�`�����8�{��0fޅfb���ٮ]�e�O,�B����5;x�b!9�p�j��9wL���D�l4L9��a�k�':}����gn��W|���Y��:�6�̷݂���x�WN����;��L���t�KA�>t��j��R�f�{�;���'�m��fw+wE�j��
�g��j��P��<W�b4�r�eJ��)��5^���zn����-��P%�]9f"d���[�fYg��AGv�<����rq��{�tOp���b0����㩖V9}ٳ�=�v����e��q�MV�'R�W����sBWCXE�kr!4�Z�1F�n�O*Ō,
G�;��̵]�����&�T�:m���q
*eh Y�3�e�p|�^�W��r���jt�7ܸ��s��Q��F�[q�٘��S����P_d+�6>�ǭ������~ߕz�Wέ�dyX���2κ��yu4d�k�ne�&>�����d�.H���y˨�se�I�S��p��Nl��q�E�2��Lf�����'cW6�B��ڲ5u�1�ٷG�U�]ee�����q���1s.%lF�p̩]B�fe�����.�1v�7J&e¢�����kq7�Kerʘ�f��UWR���cw
�4�VfS0cc��Z���s
R�ۖ�n���L��u1�Ҷ�̫�J��\�2��K���P���e��P�m��Dʵ���r.�طs�1&5���Pr�����Y����i��K�
�ݶ�Pv���
�iV�U��l�i���*8�բ����j$I���B�`9!�]5+�{��1����']��
��3�3:��cz�M��,Ay��9���T�
�����	�(A��z/2\O�i��\�=�@����-p�k�����ʃ�`���U�!�[Ob���XYժ�/)շLz�C��/%'S����ń.�5��Ӱl����92�g��x��oL0��q��=���..\sNZ飾c�K���A��gy�{�-N���c71��6��?�v�'��)��}�b���S2A�`}:WGC�v���ay�CB��[����-���p���Q@ET�T]J��:�[��V6���*�6����lVI*�b�-1��f���*P�yr���������g����C	K�czx�y��ɴ�'�5=u�d�������Z�4}�ܷ��q��+/��]K�zE�2^�^h0u�+.�ݺ�\j��	)��%���e�}k/����Z�h$���.���yc^�=�{�[�˻��$�3L_2����_%����YGs����R�S,,[� ��n���ѯ%�~1)�{|��:��JB�L/�x���a����Y�u�(�h�E
F��x�2���Ǝ捺a^���y�{wWR�LA,P�ѡBs�����ls�E��Tq�!6��F|��z�v����ˆd�7;RUA�v-a���9�|�%P)7���e�kG�G���#�^�+��x4.�zy2.�w��nm�)d��yMqy�t�-�o[��p���,{��U��Ėɮ��ޔn�v�&a�ǮX*�E& >h�פ���>������vIȑ��t�O'C��X���[^J.<�2w#���}��u+�S�0�6g.��'d��R�R�^��7�Ք{�͇�yA�Z:%rGk+D�{RK�����C�5�6�;�Ǚ��v����"����pew�&7ho[v>�>~.Ӭy�����Y�m�ª��dY���B�r�cW��Ò��uC�f�~��=���!p��E���uN�p��f1���Y=�R�qYU�&��;�*1�� �̡��Fی����9�s廇7|�Çz�X�擛Hwt�KaeV-@E=|�V�u��]�����F*y�4n�
�=��/|A��|�=�n�)x�~��C�uv��3��d�X�;7Цg�.*��s>�G����u�{f������H.W+�1�-z=�Si��qIK�Tp�����:��;�6o˦����^�Su^�%7]�ڪ�Ag�:�ݡj)#�,�k7/<Kɹ���8%Mkey���Mlm�^OV���F�ޮC��	�1�N�X��{�_��%�ۣQ�4�.W^���`L��r�ftdʸ3k�S!��<������Q��9��A�;��k�A�ev�F൝���`9[tŒ��f��B.�����K�w�S�#�\)�
K�W�L�
Z�lV񒶵U"���Y-bй<���*k\�ޑ�T��d,���[;�"��k�"M�f֏IY۽��cd^���6�Nb��������ļu�.ݎXïlVY��-���㐼3V�jFg��勠�qw�����I�.�	iWy*p�e<�G7"�_~��Ǟt"������:�(�ߚ�� �X�	3S�|]�vk�{��=��������F:��j��R�
/��7s�7��_
�����Ͻgy(��[c�sA��H�8h�\	��hM�#��Ws��^�N����L��4$�u-79�}�0P]!t�i-��E��Y�8]��Y�yn)��OV.����Vaw6l�'j�a�9�\{�������t�v�9{y�:+��{1��#�|�SZ>S�����D�%-�9Kyq���BWX����	��y}�)О��� 2�:�|�߄ؖ�}:��g�/���лZ��:xt6����cU�{Y�ݐ�A�u^WW)Y�Xz�Z�r����hoDq�t�n,�� ^5J�����F��øݼ�sF��N�t�FZ�.�xt��� �6�j���t��P�nzV_�B���<��o����n�KS��S|����7묫{&�~2���կ��$F�E�_!9A�*��<z- �z��������y��qZ뇃��)�����>�V���텰$����� I	$?���πI	$=�O���ű�K/W��M����Oߧ���$$�D$��#! ���$�y�qљ(%50>���с�����된��}��d�2�$$��Q"�P�����-.�*��K�Fv7��Ju�)��&nXgT�jK?�y��7����{�(Y|8�q�޾$$���y�g���o�����:'�	$$���$�I��ad������u�?�`�'�	����k�t(��$q��������O���=���d��|�g�)��� ���IxĒ�v�[�s����O�������]�Y?bss�	?���0	!$���7�_�O��DxHI!��?����꬇�	L/[�%��ǃ��N!��?�OO���C�9���9�a�gi�����XM���jT�`/��sW��U��>q����N,����� 2��Hq�e�X䟔?|>��������?ٕ�H��ʼ�7b�	6��My���x�Lր|NV����B�g.���m9���d� ǿ���r,�/�>�C�����S�a�%'Ԅ	$���$$������ۿ���l��	����vtp!��?���ܒ$��9?&*�I�ɓ���}^��$���I�В}�������<��V��3���2<��1�������C�Ɛ�H|���?�|$�a�$$�w���`H���О���^l��#a�}yi0N|�*�G &Fg�'����O�jO�L�w��
���6��h1aid����;����HY?���s��0�.���y�6&I��31���]�ŚH��Q0�k8�.x�Ө���|�����G���-�cv�̦=�4QT婸�]�,ݹ"[���;�tO��}(O̟`ϥ:�No���i%�����$��C��$��O��x��&��⊢���qM�XU�a���s8�<�'c������89��E	��?�H^��F���]��BA';��