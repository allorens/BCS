BZh91AY&SY.��{׫_�@q����� ����bJ�      x���E-�B��%h��E*٨Ze�KXVm�)DR��TUQV���3%��+f�J�)HѪ�V�}h�L����׶[���*�����@������Tk	�̒��V�j�IVm(��6�����5���b��4��٫aYYSm�m��7�-+��5���k6�e��ڌ�ͬZ��m,DfͶ�mjV�Ymij1f�ř�[VmD�ϻq���iQ��k4���Vmf�l5m�J̖Pښ��@9͍I�����  	�쾭����Ѧ֥V�9v�.��UQ�N.��j�UV�4�n�èC�%AV���V�R�(�]����K�s�P-(�ҭf���Y��p   �{��4�w�wT�a����r��:+��( �ǹ@OA�5�ҽ -��u C��{���y}����� .������� z�>��[kFI�[3fյM[-�fmp    ̙<�i�}�|��  }�>/:�҅���Я�� L�����im��ټ�z��}_ ﲀ��o�=�z�������i��������M���QP�c%j�ͶŬ��   ���꜍����}����u|��wwOo[sж�Ꚗ:}�Ҁq��U��z۽���>���w���@=ױ���)�ޞ=4�;��hh�UB��m�Zip  �w���u�]C�۠��뺠���pz�J�{���t��޺r� S���p;���n�s� P�=(: ��ޭ��@��|�����R�f�5+`6j�  ���0�盀 
�����{ʹ���:z�t�h=�����{�i��;C�^�C������@�G�� qz}޾�ie�f����hhk[g  +��*��`�������6��ov�=)T�2�񧫰�=��� (6�ndh;:�z4 A �}��&kh�*��6a� ��=j �v��}u@�F3� �0 ��@�=�c�5�@�Μ >��jĨ�Z+m��Rڦ��  gw<��}� ܸ��pP�;9���У�X wy��@ ���(��Tl����lT�Fիa��V�YRi5�  -x �0 �r�>���  6��
�x��T �]�頭�� P�F*�E>         � ʒ�C ���h�)�&)IJ�&&`i�&#��BR�       ��
���=4��1 �j�� ����h� � � BJ�mR Ѩ2&�FOQ�d�SO����������������������{��{foJ9۞}�F��E��<�w��{��{�� ��(�����
��� W�=G��_�������ǰ�%��
 ���uU_�����`�	>�>_���@" ���������������S��eO�`�A���>XG��<eOS���|dO��>XS�����0���
xʞ0���ʞ2'�	�
x3��2���
x�2��(x�0������2��)��ʞ2��
xȾ2/���(z`�|a�A�|d� <d�P�!�2����(�¾0�� x����e_G��P�W��<d�&�|`S��|`G��l)��A�|a�&T�|`��>�|aO�S�D�<dOS��|`O�`_S�S��G��<eOS�aOW�A�ʞ2����(�ʞ2�����#� ��>0/� ��>0�����|`_�<e_G�|fa����|`~���9�<a��|d_G�_�W�T�<`L�
xʞ2���"x�|��(x��0����Ⱦ2���Ϧ�|aO�_L!�*x�L�� �Ȟ2<���0����x�2�)��0���|dO��|e��}�/�L���ʾ0�� xʇ�x�ہ|a_G�@�P��E��`W�E�G�|a��9��E�|e�E�|a_�U�d_�U�|d�T<`��d<`_�OL xȧ��fOA��� }��za}2��/�(��*�(�� �� �*�(��*#�*)��x� ��*x�*zd@|` |d|d|e@|aD|aDED~�|dD|a`P _Q_�|aG��|dl�� fP<e_�Q�|a_W�U��`G� 9�|`�<a��|a�aG� <dL#�{}��SO�׿�1�2�~�-����bl�L��E�Ĉ�m��/AB��-g-]��t.V͎*���mf	{%`ߙr�X�=�W����Ż7K*�I�+rLh��К֍��2�&9h(Ʊ����d5y�ݵ��P�.���l�̩�f���P�ym7MЀM;v�p�Y��i-Ril1�����*���dۻb��j����,r��[&�Z6k(�wp�i�����
�6�ާ�p+l�c'H��W^"<EfZ��^l�]��XA�P��3���b�Ŏ�8tQ�L��j�pK��sA�v�o��E�Y*�d/C��{FI���2��V�FzG&��H��7�5�1�-:{3"3j�0K�J��.'�hY<5�ݧ�ݭ.�_<��C5 ��ң4n��e����I��5�:��#4�[v�.�I�m��^%6˕����¶*�<n<4��r9��]bu�B����~ \��֠J^	,��wk�{1�	��P�"���M��%Wij0�U�R:.�w���zpT���/K�3j��^��T�XE�X����r���^cM7�퓸��%�FoC��m�����3r�Ov������hԘ,�j�T�����J��t��F��H35�M�VR�Y�E�,��rJ�c�FTŁXv&��aKViˡ��,)�u��}lvݦ��[�b�}�D�K�d�Ưk7�U�o7������)$�uu��hv�`,��A�-�Z�S	$�@�+��cYY��ӵU�ﶩl�S6��I�JB��u�V�:���*�4E��c�&(�h#�H�4u��qI�i0�ԮB��U�of�I,Q�@b�ޝLcA�X1E�(B�R�(�:>���u�3>4��d�#��0�#��v�u�=�WP�q2�N�j�B��G��.�d�V�u�ْ��-��hd
��{w)#���L��G2Ø�;�b�4j�f�˖E�Dӳ�	zf�@�,Y[�E�آúr,fDk4�[����Q5c�u�.�s
ɵg��)c�����D��`Z�m�A��n鹐CvF�J"��fhwu�{,����ZuÊEtT�Y ��f��M^k4�Xo^U��L�E;���-{���ҶV����|d� g-�x}+$e'l�&0Sv��wa��Q݄8)	54�s-Ix�Ճ3Y.L���	���*`⢰�Td;[��&L���h�Q`UP=	f�Ǵ�r��M��:�*�D��7oV��&�o������pb�#k,kLe�*��l�5�KX��usF�Q(�e�m×/�jȩ���rPf��̰ʹ���z%�T�j՗�!3��Q��C6c�.۬�[�N�ySX��ͥ݅�nkmkf�a�-�`4��cKJ�^X&l`=Q��RUĜ7y�Ҙn�EJ�`�f˵-I���)akk)࡚r��U$��ü�g���k@á�E�s/l�;�8�=ܼ,����Ru	�E��Z*n�U銒q՝�L8rX�n��ZLm^n�H.�zt�ե<�R.��T�(<[-�5��6n�l��Ӷ�%JV^h�1嵓3|��4�J�*���h�J5�U���P�XMY���v�ZB�g7�ń`�72�ۆ�.��ƨb��!7l�Y��3e3���2yVҋM�{d�Q=�x�NH��nRO)�|{��#�aZ�9}�S˷\�t�X��MEJQ��y\�r(�[��D���Ni7�6��������`�w��$�BP:73��ӯP'{��.	�1ԭ;��7Dt<��(�/H�t.��mRbi�9���&�h��m��&�N
�@�v���%��� X�Ɂ4p��J�*L,�B6K/P;�6�ə��Ų����ʹ��Y��H�ӣ
��œk/H}�Va��XdtE[���ls���״l�\��.��Yt������9�En�SV��Fe\*,&V��TW�i�J�՟��Lp��s�5��4�X�!�5��cct�U]��+5u(aķY�q��9��mLR�i�#iPq/d�ɲE1�ݚCĶ�XQ�RS���r�H��e
�[0j����`�@<*i�l�,�VSŦm�B�4�����![YE� zv7*�@�n���q#�n�9�6��g��Ei�r�T:
�^�pR��������[���2U��4��4njzr�nF�45�i[Tك�0����+J���5�k���f�%��S
6ʚ0��هv���]v���j����F��i;�sJT�z�Cf�̺�����aEp����6f)Y-:�ʷ��"��wgL�%����Z|h��5P�|^���yX�љ��X�1�������5����G��	ݸ.��E���k^��=!�%�黙��䳶B`���M���ك15�`Z��0�*0��%�Ӫ��	 J�*���-U��ט ��ثT��-�*;���2�Hs*����,��V�b�2ô�;���ܠU��9t6]�V�ڽ3Q�ujLR�oiu�Jl���hhũ	"�y�iv������BÖ��Ѹo&�k &����L�vI)�+A��Rֆ�طi�ǲJ62�ۢY���������W��v�)v����ud]ł��W:�r"��/^fV((^�:����e��s!	�ܺ	�H��f��o5�Y6%.I���֖�:��U�f�i�SGvf��#��!,[��V�Znf]����f�hC�zwf�3�wo>AdPU�l25l(\��w��B��b�f�ut��>��I6��7rJ���;�o!�dJY�5b�#,	q��uG��5��՘ʼJ1Y�7J.m���t�"Ԁ�᱗�v=�n�*�B
���h�'��ɴ����6�A��W��r����B+=ה�M������"���tm-MY�V�o%�2�����Ѝ�D�xo-�? �;|�L,h�-��(�b�6�ns�����%t���*�U�T�Iq�.�3v��Qڗ �Z��0�3 �S啉1���Jʺ��WmV��� i�j]�����{��Ho��4s��e+܆d�B����{��6��&F��N�୹)1l��!Dm]=6p�6%;`�B�Q����x�-"+2��@�%+F�i<.��=۴17o-u�_%R�l�������$Nb�����
5Q�� ÅՐ�[)M�O6A[i^�5S&#��-2ӼS�J$^�#�순&�fj��3(�R6v�/wtX�Nơ@���Dӈ�K(C,�
"��©j�La�8.�mM�âZCUU^�1S��Դ�Y�]��w��s5U�X"���\ӕ�pkt�^9��#F��+)�F���SE㘝�7���u�͌U2�[v���օyt�݊�V���yf٤�FB������2�:�=U�A;Xu��wJ����tMa��^�N�
�@$��HF�Ii:0����kyneQ���Sr�.L�u l]G@�{eՆ���^^j���d��ҫ*�宬ݬ��!�Y�5�x뎌ἃ�#���S��I�����fڡ��j5WBb�H�r:a�+U��\��D�vI����sTnskr�a�ՃF�y� �oqǃ	����K8#,�����������aެ����hn����UrvU\�pF�����0���6d�{)ㆄ��CV���������G/0�;z5:�RA�m�����J����wE:Zn� �s*,a� j�Lүe�iܺ���8Zj<���(Ҳ���n�t/<�ANcq��@[�x���TŸ�
�Y��@��Y@��F�7�7c�aU�\�V��44����#)Vd����c-^��	�E�ֆ"D�����fV�[.���^A�H�e\5yRT�����#���V��A�i�X��H`^��^9��� |\҂���A��	�J�\�P;����Iuy3c)km�j�E�"1�E��wK!+X�(o��f;�tK�-U\�Z���7hl�֬��f��a0�de]�u77lb�-0�Vkp՝ǹ��2}y���u������&���6�#pd^��j���46��Q۔���r��� e˫���h���);���ޭ�f�[��,���J��`��u]w%%e���</xk3W%oX����7��J�z��e��id��t�����F�u�3v��(^Q�X�+��z�un�w@W(,;�sw����|Y��M��t(�%�^��m�Z����Y���m5D�/]@�Û�r�]�cB�T+\��{�MK��ݪ���X�%'�%�a�d��BEX������[{1��1K�ǤS��y�v�,,vN��tZ������&��%"NR�w��	�Wz�4�/B�����,l[G4&�l�?�����J�G��N��+bu��Z�9�������.�y�1�ݷ{��i��
��9�`�n�^>艹���:CwXË��;�pYu���ihX�뭴����r�Y֍������Z�m�����E��5u6�,�fQ9WtȠld��,�����cu�,�c
������ִX�Tf�C=�]������p!u[1Kqi$=��#�^��4�!���8�*���Ԛ�� U�滁������M�i��Rŀ<�Z޻�x�^w/�jxE un�.�D7&f\#Rj�8Veu�z�@���lj�f+�XmG��)���S�B�Yj����Gc�eX��c��m��em��*��,0p�I�-�n�0r���D񱕄��i��T�a4�yU�"��r�8�7X)�/"r,?Z,�8�n����5���i5ݼP�U}�Ze��-WˁR�6�1sm�X�0���;�'�&=����t"�u5��j&�ea@�������a�kJ�UsF�X\X�*�ʡo-�'t�m �ss7E��
3c �f�ݬԲ)� E�'�EI�!VpY�4r^Lɂ�(�`�j@��$øQfCR�����֞��(��fj�Q;�a)4.��z�a�ssT)�d��1Xy�-��T��̶�7֭���'�ږ�kçl1M$#�-Y�֔*�K%9����Y�F ^�T��Iz.��1�䴅���/�JM�qѴ��94`S.M������ȷf�)&�h�j�ʹ�5g2�(���E�ɲH�gj�P��Q̽-ԩwk%Fs77F���[CFE�e� l��V�� �
t�區����uk"Src��&�sA�&�vm�%t�X83ma��gv��&(�X:��CA2�[/\o3A�T癿]�D#�ٔ�n��;L����
��	7����^��
 �q(ՌuG��ӺYjY
j����dͰ��`��`�/c�a��,�Ϋ{MGR���҂Pu0���W�B'��"p��oҷ)ӎ�h�B�d%v��[D人�VQgH�9[z����#y��7�i��˹J3fp�"�
���ൖ0�n:;�٤�f�t[�kP��t�N�Ѯҵ(�ę�vt'un�W�����:��ҫl-�Ah��z�n��i�4�Y�G�/w"���;9�4�#�;�Ei�G%j��Xe�Ȕ^j�g,����a;4R���rp�@���M�%�Q��v5�Z�R����I�-�v0��9��@�nm�ɶ��-�e��y2����H����%��!j�	�%�D�3M���Z��TYW��2��Hd��U�mb�,7���Y�C ��Rf�� O�8fS�W���V���7,�F#�{�A�0�V��*'�
F�ېiw�ݼ{`���N]jL;���D�dp���_S��E�:'�5��΅�6�IKr��+5)���U�*�6�ԃJ#B�BHʸ�;!�r��4��Z��.��P����2��a�2��ܹWE�W�Q�Ũ��!��ܥ;{%�����e-�D�����	���Ħ��D���<��p�ri�p,���9�z�Ve����Zf;�S��b��ތ��3m4�ǘا�Аl�R�)%��xc�n��[V/��fĬ�0�P�N��^؁��>ɠ,)�k4��+ͺ������h橂�7jP�����̢�W*��5%���nin��)�9PY;���KX��op3P"�v-S
Vѣ�a�����c��jyc+Io���M/lk��&�%Gt�m�MD�����1�FG+6+��j(*�I�e,���w*�6�"�-[�NE����u3�> �^��Ȩ)�BXd�T��(��uF��5�v��H��`��Ӈu��(�xތ���u��J�l�Aw����ٳ{n����h*.��`:E@S��F7Wy(��7��M'&��@��*�n�Q�/,�L���ۻ9F������cЮ /n��X���JE4�41\j�&`���F<��8#�Ȩ0���-��FD;WB{�(b�2e��Ϋ����];��6eh�4�y�����N��M�:��	ȍ�zVjeS�U�[2��4��Q.�.fp揦^\7"kdd
PU��x	��1p+���yW�vY�g6����4�L�����7��ӫ�o��p�ލ��q�0�'�$�2��h.ǁ�"�B��(( ��e�eQV5�� ,y�\0zK�0��'���&��p5Iڨ�U��	�)Ȃ���&��Dg��yig�=��&��P�6� �#�׈�ز 1 �	N��1�#|=�U�Yb�����Ć��|� ����\�3K�� ��aڛ%��LS4>߫ft��Ѭ, �-���AПZ.�a� �@�އs�w��]�b����VZ8�'iZ�'�,�0(�a�	���5>ѨטQx_�J�
���r��7QM���pM��Y��&(�	.̀�0�*�0�Da:]E��&&�*J
˰
p� �1�8���
Md�����a8XC�%Y�<���U0��&�GV�1SR#��@z�Z3��66�(�-˲�o�{��5���?����� �����>�±��_�Q�#���ڕ<�9=����U�n�]R9���5T�KGQ7��"3M[�M�аsw�I�W�o�˱S����9���9f�����n�S7�H�/_b�5�<sr�{�{]vi�9�֛�	�o���$���RS�;;���Q�uv�mSPvA�e�.^��B�R:N��8G\����]}ov!��T��9ٓ� ��Bt,`�U\�ύ��*s�L7aU��7	W�d�Lvh`i8&ı��G[�����zd�2��k���R�KgB��ol��/��(�m!c����32�.뽷m�Jdه�	;/�8n[5��gvr�;��#D���lʼ�xʹ
Ĥe���<� 4���wi��>��]����끔�.;Idٺ��s��"`���r�Ž�/mL��ɫ�e���4ktH��(����"�怒�h�g91�0�f
��駽�f�Q;�U�$B�o_1��S���U�⒲ɂ�'&�����[��q`��\/R[V�_*ھ��)q�-P_#su�������5-�Em�^��*�'�	�z�%���Y;� ��v�+6�[#riA�
�$䯡����Mf���R�:�,���5xpv���1���.��D�f�i�;M�N�E:{5luy��XQ ��f�K���e\�o���l�@"�-u7|r5KP��*�����r*0M��خ��Y�sS��[�Om`�8�×X�Q�w�L���t©w�H�bJ���
v������n��U@��=+UX�y�`�Eɭg]-�*ga��,�K�v8.q��0�{�8��$:���G�8�r�ld$48�h��X�z�q�fQ=f�2��2&6�/��uM���\��bjxX��e3ڙY[�]!�YBQrWWq���N�q)�{���o1�����3�ӨU`&�ν�^k�E��\��Tu��rƭ��^S�d��d�l�"���={��]�vU���I���]R����\�p�ۨ���u=q|��8o�.]N�Ռ!�侤��
�u{�59�O����J��p�isw��-JĠ��NL���ş�0[�]��]UQ�]k7��%��W��8����+�Ew���B�vn��bT�\Q(�x��(J��@gb+�����r.i�#�f��{c�"����ɮ��*T�*^���<�O�X4�S�2IR�4h^[�I�c�KV/�J���"��4sRif4Hf�"q��j;f����}p��t^m�u
�;�w.���;(!ð6�b�73W*4���qAe��\4�ILæ��"�r����<�yv>����'=M�%�f�P��ҺQ
�.bV��,�ط�Y�Y�qc�[����N��J�ώ�w.��,*e�t�B:F�2]k���z�Bmq�,˺ �j��c���BIb��攃���㵱�tf�>k/��0�N���y�mSe�N�2P���4�Zi�h�e��}���J֕��l�7S��( D� 庵��ɤq��l\�Dr�����r���t����M��K�wR���a�5K�*^nP��=\Y�N@.2��76M����Vv.Un���6�(,���
��݅���`�"���L합#!u��!��3c������]���;�m
A�Wj��"��Ӧ��j�w�F�t�Ti�*B��pr��4f�Vuͱ���ad|G ��[�n�qi2�ׂ�[�,��k�`%���%�n�;�;B���7� 
W�Y\\�eXX�x�x-u9�r��t(�:�1�����\uc.vޑ���$��u�_&��,���{��Hz�*kv��ۙ�quIu!���h�5���p�����A��
���Sc��E��(=e���D�{+�5bu^_v8a]6tU�;" �Ӊ���sO`�!�|�YXs�'jm3��w��t�8�o�wu�#G��P%����Rf>�w���w��.�j`�6������Ӳ��$C7�Ԑ��i�/�]K�|��.T�0��k^�v��I�-v�tŧ�"k*���,B��)��	8^�VCo�E2��'��gR��Y��N�WH���[���ʱypX�t󡎅>P� 6\���o8�]DHGxay�T0v#)���$g�4�l͋i� )F�_P,����o�zed�\t�K��7or����4Y���P��� UuڳY��1�9i��Va������e�A��w J96�-��Nk,�D�͛6[�r��S��	;�#d�W��E��`G��eI�%��kR�>����D��v�o��lNHe�'O3�8ދ��oB��j۫�l�	�ydd˵�����la:*��&����.Am��l��\Zϣ#&VR�������nm�K/�vl���	o�JK��`�;�s/fKϑ���='Le��D��Ա�95���˒e��	�%��[JƃvrJ�i˦�y�6�pY�W��Kk�)SѺ��c{�Y�6bܖ���T���]H�5�:�FL�w� ��*r˯l��b��-�U<"�;�I�-�o;E��/���j�F�R�|\�n�+�}�5�8�:��­@� ��Z�u�ˮd��K�[W��V�S�^�57qsvM����-�ís�[�2�Ds���{�<��J�!!��(�Fj|�p�O?�0{C�)0X��v�z��R�E��j���ڙ �n[[�1�vö.t�X���}:t X7[���ٿwn���ԏ'q�����/UƲ�n\�ܗ�g"Gf+�kL5��oP�C{M�c�m� �1m�iݛy�x�ge�+�oa�q�$�hE{��(j�G+���u��)�NC۔"���.	q��'rE:I��[��-e
ߵV��U�[�d�l��D�����U,�g��j2���t�wv��zݻ�m(C*��ط��hm���xN��-���W�/�\�����pǛ�m	-��8���U��tܓ*sV��t�)V�>vqW<c7%�Y���s5J$tB>h`���o:�նu����W���]���Q_4z��%�vպ��e,3������3(�� �uV�<f+�[�(T��)NբN�;k��tH�}6���۹6�,��:>�*K.��EL /r����S�j5���/#���e*\jpP_��a]�ՙ���I��>�5]��2Ig$:*�9���0$�ˇi�sN���$�k�)i�����Y[z]gp΢�9��WeL�Uq�jұ���V9v��#a̽A��qm��Wbӑ��G���}oT��Y66oK��h;4��E,��fW^�A���ԋ��øl["n]�4����:}7�m.֕����W�.<���6��Cy��M�d�`�(�][<wTZu�{Y��i�Q6��v�iFEt�P+Y�kp)�8K)�T�%��eA]������h� �̗���� B-D�ɦ�u�Z	�>6�M�=��uf��L숍��GN�^n"E�N�gww���Q� �=�C�&�Vb��w8��"�Y}��!���k�541s	����3�U�c��ed0�1�L�S/V哉�6,�u���/_C�H����]sV(�Q�T��u��7���}[��"��-��K����M�],���ݛk`[��ub��v�E1�E#���mb���$�R��m�%�t��K�y�B�R�0����.[�I�̗A �P���m� �ҵ���
Xq��X1K�6�v�Oj�1�����r�gR��IjmY��������r�jq�o�4��9��������
�l���'zЧ(��,�,m�<�RX���E���-��.�cv�TA�����O˅l�u"�-5E�Y���ٵ �u��N�Vbm�Y%ˑ�/��7���\0�h�H��ջ����\��x�0ҧx��}y� P���o��Wtf!6���W+��Ҧd7vxh+��k�h!��V���t��$1\�e�d��Zv�p�cޢb˦v���v�u"�d�\��'��݊6gok��[E�5' �l�F�:<���\��
,�zX`k7��c#��͝�2� �!��.v-�<�%E����0f:���O���C4i�7z-^�k�X�2��:�3O2%1�u����Go�N�Yա}���q
]uS/�,c4^�S��xڇcYz0�I!�l���,���ծq̙e���|u���HN��nj�{V��BT������ܴ��]�p��W���2͔R��`��02���^k�v�KLt�S	���uѾ��p�1�=X��IJ�r���).V���BU���KF݅�oz>�����<K72�;��U����4���l�j��]��j1��f��=��R&�b���3�=WJ���2G�J�`��^:U�
�����8Ty�M���̙�ؙ�.;��{W�H��Fج��Mqi�7J��*�2��!$�snSTX��(�ʹ�3���)�j`�TC��J�H�w҂ar=����=�s��[�Mɧ7��S���z����_j�����j���Ε�����
�� -�l"��I��"�L�]��as��G>r�ۺr�m���nu��+��#����j�Cd�����dI 3�\ne-���+8V���Ջ8� \�����τ�u1�qZ�mf�+D�2سuQo��t�4Y�'ERټҶz�ܑ���:�L��;�|9!.`�-���n�w\J�:�2�A��\l���}`��O1���^E�R�>5Յ����×��3�k5+�(��[��;�+r�� }W	7I�j��5$�D�����,�D/�Q�ӹl͠�1<j�%�{"���D;^к�A+5K��o�y�o3��'}jr��^ء��JV��6� �J�u�B>��ׅn���"�2���,��V(Hl
M�h���K :���ƝٍG�]��,��}PP�f_Y�g\����k./���*gFo$���Φڜ_,|�Y[jZCPoGG�����w4d�w�l[��C��]6���*N+�3�ջ�q��oOc��f#E_&R�of���a�(t�R��,����u��#ȅ���c �_S
,i��z1�{0ԏ���܉2d�c6I�x���ZT2��L]��ROuӺ!��MH]�Vm�G�ؔ����Op���Uģ����#�7���U�ɞc9e�yn*�1ɍ:�-�]@آ��J�g;:�T����Ïc19�͌�u�E��j
��ڠq�c�M�r���FJ�p9	�`y^�m�Հ��5���Z3����J,�K���v]wE��\Yh]`�%����Y��'l��� �e6�X�v�L9X�yWۜj��Z7r�s��I�^g|�
,�5������5m'N��@�ĊX��]n����3p��S���3K�M�˒���u��� -9w-lחL��&D������͂ؼ��F��
���XU��I�OXͬi�������BnP[.S<y���q�]���0���س���5���3�c4˱������3B�5�bL��z�sG�+�6e��W%�2���\���ز�6��\{:W,�;4�M
�Ҭ�uts��ц⬔�#�(*^n4~�4S�^:�u7�N�}G�|O3�/gX�-����,���E(���R�N�Mb}����wH�:4(v����Z��`ٺ�*=��8���-�P����Y:6�N`��Wvc���Ν3.ȼi��pna��0�(�T��侬,�/6���U��o,nw@6���	�`V�a�T��!�<���5AϐWtƒ�E�:��j��1V��Pb<�g���"��+i��k����Z��R�#��I(���mK�⻝0j���e��F@���n��ܾvv���Ჱ���+�i�w��n�^�EBB�����l����h���+';��:�>^U1��v�,y�|֢3c�ṖM��jZe�ZW:K6���y<���]G����K�a�9z�)��K8�p̎����Ց�M�.��	ǉ8KR�T��é_`;S3a�҈�Yͭ�����t�[��hm�`��@�f�|8�n,��8p4eX�2�8g-g*�\T�>v�\Qt��"��{�blh���S�8K�[3m����� �LTzm��	�e�@�>YGN�Z�fV��&U=���2ӵ*5�ns��n�t����؝Q���^��۹�9�:��X��&�#�1q�1C�]\Z��2ch�ȱ��ʂx�ww\G<��Xu44�n�\���[�	��T=���Ӧ�Y�*qXX� W�;��͕{ѝne�t����cf�c�H0�?IX��C��pc�]6_fܘ�$�xr3�p�|v�A��8�o��P�GZ�r�+5�Aa�X��7/zi쭛v�*�[BӾ��[��}R�R����������:�T�sr"�$�I$�RI$�RZ�LA|�O�N��#�y(GnK��9$q9$�D�I$�I$�I4�@���:�����-��Z��֎�`18��E�=$�L����������E�>�zϽ����>=d<�4?����O/~��^���P��z��G�}@�_U���J�ԉ�z�z����������'��<��P�A��(���~{|�]��= ���>6��OR;́�=�!�S�}�������?���@AD��ȿ?���	��?��/��U�/������??�������ְ[-�3��f�Q��P��]�S��H�bdLt�,���ë���>�m��U\�2�4�i.����A�&,ڻ9;j
�7;Ě�f�>���f�.�#�QR�}Ht�f��!�p$65S���C�����1i�u[0d��ٷ���Y+� {U�A+l����� Wܹ�ȇ/�[ڽ@+�q����B�iɤR�����&��C�nV��Wl�^e��غ��e������!�֨�����A�2ȚJ�	eI}B���0v�쫮F��5�<lڣǈ.1ۢ1�c,�bn���#��ۓZ�d<\�o��+�L&ɁUaYµ�hi&��ǣo�b�g�<�V�p�o��)E��M9:�Z[�~�5z3@�/�H�]�=�6W+9
TC��RrR�H���5f��x�^��K�v��Wc9��'�_A���KcO8\KC�k�#��Ss��W��8'}R�(cw�o��j12�=���(�l�Iu�7�nA����{m����o#)u��G;-����7{�����0v3t�u8$��̷��a�f�E�-���g��w�U�Vu����?e�Zcg���;p�-�^	�hg�)��A.�oZ|y|�&r9�}W������2�ud�P�;̏j�e�^WR<�8J:���˝���t �Yy��WN�R��ha�ö�Z�m�Z4`c�lWJ=Gd�nתnjj����oN�⦲�-��`�Li��Z��c�ssn��MG�hҧ"�=Ǟ��r�}Z�7�L�D�S'������,9qQ�1�W�\:!�μ�\��$����X�LW[XA4�APZ�G��Z�qt���[�Wr|��A�F>�{�>���=e뗬��%�����67��OxWX�kg�K.��O\t3�v�Ob��N���Br�h��Â��b�GX�2�b�"��v-�W�5u"Ɣ�X�����n�������*oG}�5��;6B0.�*6�TD�q(+���{�^ՇI�P��-�������#2ݣ�se��ٵ�;��+�czZ\P�0�#2����n֧���
nu�Es�j��Y˨a�U�ul҇�7>��b��v���j:,�[ƯHى/�:i�na����f/WN7��5�2���Nn�]��8J� ��F&GJ�]�����C�߹�ڶC�Qt�4$&��x�7w}����Hkڞ΁Nsm��������[pv_NL��Nu���INw��9�|����B�K�W�����y_�w$e�K��ţ�`rl�Q�{�bANe�Hkf*�w�m����:4;���E���xSJ���u�:t
�;�fu��ϕL��U��xNv2�E�z3��K�}���H���:�A�ɨ��w�a��3�%��w����pы4ogCL��m|ZF��6��j�-8��i�]��C9=���h'Ve�ٙ�рf;�WMM sz7U��	Hͼ�|�A��n.�����!Ճ�E��Vy�K,5Wu�Ě;G:�n�W"��(EB2Q��8Qp��֌j�J��SH����9T=w��*�b�H�u�'!�f�}:�ǘ9�[� ����S8���;˶hʤ���"I�[P�������Fu�2�/p��e��to.�VJ�żēk,t;��E��2:p��(IK7�K��-���1�Z�["e�9Y�[G��պ�O�SV�č�$�de�˙Os�G�k7x�;�b�J�T��")���V:f��5��@z�U0�Dil���e ����_%��R��R�v,w=�`�:�u�crW7Rb+��p��-;���{���#�����v�� AQ�=ki}�ō����	�.�N�;զ�D�C���hdCT�l,��O�s��!w�V\�6ix!��.���]=g���\�e�*��F��h�ĭv�_m�u�f�aj}}�ݯhZ�Mu����V����A���9��3^�E
���*X��B�����(U�tp!��Z�i�.,a.d��wӡ|�	E]ޞ��f;����1)�V�������Ǜ�e*=�2!�G�VEm�ϳ��h�"�1�9W��as���D�c�6��h���?roY�2�*�o.�6��sI��o6��Z���1K��6^� ���L6��n��tI�
v�\�}o\{�K�6݀XY�V��LΪ�qZ2Y9�.�Y�@_,�v�!Q�d=��]Z��[{v��`�R&4Øp`K+�Z��8o�P��+�s^�e)�s얨��=l����̏�����H9�.�82Ns��v<K��6�k������2r�W��)aF�p�V�Ӂ	��3T��­����3��k�5�VaWX��Z��P�\��b�WD��"	&���r��������,Cy���R�Tٮ��?M&��Eª��(.ú�&��,6X~�o9���R�ۙ��K)�i6�G�ï"�G������l6��n�ԏP�ȯQ�������4 ��<4v�m������s//8N��ڱt��`�ōT5���1QB��b����L1�c�3C�-�k��*�-Iq��"�s@J	+Q���Y��7�:����Z�FA=�V��oK��f�\��򻵎P��{��m5���7�Y�+(D�UB�zY�ܱ�sJ�%��,]�� 
��_�>�Ȓ���j߳DK��f1�E�]�VL\J�s8��]��<&�y�el�k廐ۑSu�����;�k9��{0��w������X�}I�k��-���R���)f ��}���}���(��ɉnkr�C.�zܥ��t�b��f��ׯ�`��d�I�K���a�r�B,�s�/��}���U�/$[C��|��E�i���{����%n<;�ǧ*N���lPd5��-�p�Lx�Z5V�#l��;�S��)uL7y�NJ��	75:7���f�8N�M\��um��~,��(��l۫�ڱ����pIt�Y4�>N�����q�x�C2SӅr��ê�
��A
�o^ɥ*�Z6��B�u�<N��Tx��!���6�ӻ�_d�Ms�*o�ב ;�e�v��$�Ug.�j���'}���Áf�{"��һr:D� Hb�K'sb�nD��wA��d�.Jr&h˽�S����c��p�7�q�M]q�2�j�2���BA�	,�U��+QJ
��Z�� 4�a����kf�k,�du��������&�Tݍtҋ��Чa�0=��+
���dlI0��ou6�>jb�;mؤ�b0�Y8��ctzV��V�կ,u*@"/��ePb��ew+���-������Z�D2��O0�=4�whΈ��֡�A�8��.�
�ـ�I�Uuv��Tz6nʼ��p�[N�=�KM!�tj�Xw�0����nF9�%�<U���}��
�==U�����Nmv�0�ٳK�d�w�);/�1dmao�1�ӭ]�Q��7Y��E�/8���:�E�i7�6HP��7k�K����n@Ŧ�R,w�^[N����o���]��[��k�n[o���jqr�@�W�Y?]���8��'�J���h�S+h⺴e�K��F�jJ�h�����j�}��P>*���VP�� ��v�s�P#�e=f�O��}P���a�����EH������:�T6o(7���K�xa�zv
��;\i��[5m�U%�C��*ծ���b(R��i4�;Y,AƎ�eN�KZڸLIM�b�'wg/I���;� ����W7l��q�jVC�2:ww5��V��N����n��ȷ"��HWj�M9[w/f2��������E�6�7wi�[rVʓ�9�ɜ�t�*t�3[Y$��ɡ�
��5r�r�Φ5G�<���za/*���V�T�)t�\a�_��T&�U�64.����[11�B���7��n�ރ�&(n���'�h�9.*�fY��͖��a��
)�n��suZ�pHP[��yU*��D��>���B)����UĘ�؃�1�������hP�ms�:ۧK�A&�a77{Y� ��e��P�������¶�}Q�3��W�x)ꂊ��1�t�uN�@�1��3S�u�wq}.��.�3P��I��񒮕��]��w�ۧUq�k���>	/�<��nP]���۫�sn%�˕����L���-г �n��fܥ�Û�2�nU�B,\-�a
���o�	�1��p���f����l����A�j��`'�'H���P��B�@�b�cVsb���سm��cj�(-HEf�ܺ��6�ƣ6U�[�'#`h}��8;�V��pa�[�,�q�<挦vJV�����xJ��U��;�y�AI��x�{���W6��:�Ύ(g],��zX��\r��2��m!W�7��3}Ȇ����)hGY6�	�h\+1a!�1�����Ûz뭾C�˚n�v�mչ�|�d���/��o5��ː�Eغ�
ӆ�,i���faZ�Q����A����Gwq����>LA����`�����B8�c�W.:�P�1�\-��@��ggX�	b"�vu4�dS2wX�2)�&%�P9\l_:���[%Κ���q�(�)
�\��F�f��y(=0W`t��U�m���P\��-��{\�}[�b0d=���&j_Q	슬N�B[ް�Ә�wzY�5�6��se!c#�ݪ��8j|��ԓ���t��BĚ��+4�V.�^v��Z�i��Sn��y��v�����ř]x*�9M��f�R:�^����
���P�����kNU�!6���Φ�
WLoڢ��"���R���b���{IB��M[6k]��Z�@�^]1S2���ϕX;��fk��B�)ʧpCH��d�/����#H��E��o����LS��!�&s���I*<��&�I*x>4��üEbA�c5��cnZz��Ԕn���^-*�=ۛӳ��o�����m��T��ZzM��8Ь�S�!��Pz2��/{;��Z]iry����
#^JT�Ma�W_A%���c�V�X2�YZ{����(i��GB�u�L&������wU�[CKG.��$��eծ'UfB��\.4t!����F������2�H	^�:_�\"+�E)���>C�0X�is�w�-N8h&�<^5�~.�nC�<GR��͈K
E��r=:�A4w��w�
�dPi�!�2l��ӱ��)Hɭ�ΰp��J��xN
�����v�Fh�#��F0-fhľ�����k��ƏE��fP��
�Wnݛ�2��'_]���WZ|�u۔H0٫
�ms,<-����a�T�H�Hxe�2��I��k��@5"uw$�#*K���Z���-o�{+���}�a��AaU�Ց��W{�z�C#˻�%�L�6M"��v���kv�e.9��3y�ǉXL���d"�3,�1R:�F�񇨠�o4���obo3��wG5�:�G�P�)C-��|�gU��q�e>�-��o,P�H��xbG,D�uZ˩�����ZNa�u��
���(!RaxD���5�_k+R71�r��q�A:m֦�U�gl������W�v�0����t8ٍF��ݶ��kp�'o���R�n��R�\U͇�lE�;����Wv3M��\F��ң4�ƻ��bf��#� ��znLW��wK9��cF��/��uL�78��uW�jf��|ɧY��]{|:i��I+p"�i�9Z�-o��<qY�|D{h:�qʔC9�g$t��� ޺�= �f�ϑn�CE�������Nu�p�7/���ڄJq�)]�EU��c9��U���kT7�a��;GN�Q��V#�!7��i��Cn���r�k�DY�˼`��)�8��mV[��k�N���V���c7��yq�XЗ`O�KjVێad�t��Tx�`�������,j����݆��5N�;9�$cU�Vv��t�Q���Q郱Fz�)��1��4�LV���Ü��:ή��e�4�i3��k
݃�rڔD�0�9Y�E�����H��_#m�1����M��%Y�
�S.�qe��1t�8�[T���4˿�"�G;r��f���Z���պ]�#ʾ�w%�h��u4��G�p#M��EH��ͻ�2k�d=��I��L�lp�0Y��i�{���#�kv1-mv#`iC�V2"��wJ��J
E��t�l��[yHq���oRFM�G$��ujGS�����GO�>g���!jF`6��G�*�Od�&=Ȩ��7~a�|n�.;u4�-uCo�D��9���ha7���ζ�V'mf5�!��:X�z��73��c6����bul�[v�)K�]��t*��C�c�i�1fV�U��s���/a��q������Y��X�VIFҘk�2���29�9^J�iK ����2�O!Ĺ��Ͱ���˂�=�ooYC°���Ǟpsju
)���#O2u�US%Ǧ���������۲ 0��Wv����1e�De�K���_f1n�m��d���q��j�<�3V������ZTf�U�����u�96��۩2k�$��X�]�>�ng'B�=nV��|�2KL�5q��˥E]Ǘ�i�!)P����X�9�Y�r�uaw�|DJb�(\a�mv���h�u�\���Ar�tc	�{�wy���QiYN���N�ߪƯ��,-6/3o�ا��]́Z��Ѳ�EX�}��r<OHʺ\|Rv�:mA&S7��y����
�NJ˚�T�J��c�d�Γ,,7[���S��^�̢l�4$ѕz������� ����$�����������`���������������}������}��o���}��o�����}>�o�r~=�<���r�4�F64�.T�%�"��OѤ�?@R��������,Ƙ($��e��'�0H��jDbR(a�F���J�d��y" )QC /���R2Z&D�E9��1Qa�Ir3T�BF!��P$��	�D�
��yf�Y��qRճ)��-��/^�4l�kN�jeV�^>Zg�#}G�)7�Id�4����]ZH�Y{��֊�VMUl��W�C	���f���\¨{EY3�v�'wNa�
6�:[�5�Ń�掖��5�����7,���۵֮�~CtN��t����V�����Y�G�&�D�Z5�rJ�y2�K�q�:wY��E��j���u{@�Q���k��f�m͒V��j��V�W0$,͘

��a"�b�c�Bm���e[���0A�;]18V�����T����e��oD�x�=�-�����7�hd���+ڲاclR�JwEWL̹�d�n�ޭ@6�;����ٯcآ�k��wmk�t^�-L/&���I���)��jmZ��ER�{G*�����:�i�,yϹ�Q�q���r˭�0E�6�Q��=�*W/��P��elH<��rAяb��D��=�Y���T�c�lbU�u��koj�+"�/l3�rĭY�Ms����oP�I�V^f�t�J�r!���7v�� W\�g#v�X6�$7�J�GB7(��\!�Zl��2,����u�oH��F���p�[����aV[T�)�+�M��b�ˢˬ���s���5@)2���d�(��;c�qW+�q��E+�(j�#<�9$�R�I��WR���akc��ZFG#h�R06�"b Y�b<�T�� �C�	R�!�A��z7!��mB )#�"i�K)�܋���P�aM"$�3��\m��.hƛd2�L��T`� �rNU`�P�a>��Xa��Q6�1"B(�I�2c$H��(a0�ZL�柘m�bQ�
1��m$|�H�PN8�
B�i�b@��ZQD$�d����j�h�M#D�YMH�)�a^5A2��I�W��	� ��xB\�>svqth֧cWmZ6�]����ΜL�؂��_YԐE�z�[E�(-f����Zb#ջ+���gmMcj����EUQ�7'[Ztw=q-dմC�l��E��?|v��X�Tj,QEXΪ����T�E�n��X��f����Fk`�*�h����6ֻ��ŭEEQv5�E�+���
pl�5�d���vM���Z,`�Dkc]nh�n�:��D]�DU�S�(*-cZج�llVlꠊѽX���&�*h$���ӋlD]�Gj*�b(�c�V�9{/T�U56�TUm�AcMm�E��c&�"�����\d�B�����=�li�тi��A�Mcma�(&M?EӦ��Q7mEthbJ��m&�Z�o�'�=q��S�j����DQ՚5�F6����LEEUEl�l`�'UTv��i��$B½���0+� �j�'"@Q��1 �o�2Ai�G^��/�Z��ǝ���ޜ+&D�C'ΔYo`c�nL
��l�EV�����}��u��;�Z�s�ή�L(ϩ	���D��$�l��H�L �!�A��1�E�bb2|g�AD!�H����D�8ES��v���R�p�7D��7������qk�͏z�A���>O�nB��Ў��a�F����ֳ鲔�fz��ޭb���I�O���>��dʉ�)ה���u�A�ɜ�s�}�G1�s�o���#�<�h��=�8���R�a�Py�'��Θ��m�Hl�)��.Dp1��#o�v	6�޽z�iM^~`F[g���)��Yc�`5����;,�Ul�2h�Ë�L���7��ؓ�n�{�cr*��U�EǟA�v�0��ɮ�.oz��5mf�'��0��i�gbz��x���L3�^}�{8Jq�3$��{˶���/�w����@|���o��K��O=����:�~D-�9�5��G>��y���y��#�?{�|^�&������o�_)�=ٷ�5}	�z��y�Xa�W['\� ��P��G�%�hc�֚h�=]veh��Ңl*����4j��`�z�����H�����[MmË啓���2�p��]��*�Q>��l+������w@ѕt0��p7�X�c&I�_]v�N1tx��R6�\ۏ�L`>�rN�N�2_E��=Y1�M͈ȳ8�X��c�π�>_X�r�]����Z��iܮÓ��{ދ\��RB�;�&у�j�����1WM����G.��y�Ɨ�7��ڼ�~��ޒP��9.JR����pU��þ�����8�NCD�4��[��>�>��v���ONj3�ZoD|0�!= ��jr��+̝�39qR3�|A�<|O[^Q�!�VFg5��Ӓ����(|�P<��^��j3}3���wh��l�sELB���\�##W�sj����1E��#��E7p�0����Aį����h^c�d���{i͙$�s��m{ep����\�pe�%ƽ��Z�^瓦�'�K�l1�h�$����r�����%S��6����6�ɗ=#��c7ϻN��<F��s���<�ٶG��ݏ��Ds¶�
�����B�TVQ̽Z�R��wAޛ��&o��^G��b�������~s-��Y��y��]U��l�a�8Y�G�ΐmٳ��e^�FBʚ�O3��n���O�Ƶ;e��x�e������	�a�ñ��S)q����׎^E���m�Fe��X��v��w:$����OO������M��I�y��~����u�ma�uW�A�א��y�>����Ả'~9��=��+$X>�ga��u��wãfvF��V�<�;^�Ǽ�K��G&��1�=L�����%�Ҝ��^��
��]4���3�u����6�L�_����9�Tf��*ޯ��;�^��]x"1b	繧�seV?u��~��^�IQ	5�����v��{�C;�l[�a�S>s��U=�j||���{L ����#����~������-K�H�_�f|i��{���#}�V�<}C��n.}<W��zQy��ל��}�t�v�&��J��G�'� �*�{�>=�����#��觻o �%7L�+�c��Y�Y����%{҄���_�O��l��!/.�AW�U�ݎl�U�Zp�ew5:����΄R��&y"]�6y�{�F]pK�m�yMK�n
�Gp�W㓢Sm���iB��d��r�N�v�p�n��_u:IB5�s��x�^�,�2���x朻���
�m����f�0�y�7��t�����l�x��>�ѓ�5~��5��0�[�E��朞��������t�@Y�43���ƙ���{I�T5��l�C�[�#Xc0H�m������H/'I�_���m�F{Z��^��ܧ[�����b����:Sh�����Ǎ�$�A�����6����(|b�
�[9��*Qz��zC{�WFO�9�nx��<]�ꖔ�i�43C������U�{tr�W���)�����8AE�d�j	���
����7j�>�@i�OE����%�u0�{O��UȜ����6ˉ���;�{�^���߁��l%n�}r�<�Nz��=r9V�wk�"����nO{�||~�3���>־��b��?K�Xc�{�4p�]�_��3�	����s>kއ�>��	Z�H�ȹ��Y�X�M���ʱ�YFc�X&���=!V��)��FN'�YeԫaW�*�> �W{Cl��Aܕ� �LWX��x�	�f7c�1K�w-��`�m��֘�TM�P��.��S���|���H����t�9���c�@�ni�S^�����ιA��f"�'DY�k�8�W�/_�É���e��ϵ���ˉl�e��^\�s��?$ܗ�)Ń�5aρ�W[Y,z:��}���ȳuڇ:Kvo	��E1�+�W�#ǹ�v
3�~�����"��Ɉ���&�s�80]^�<׍��]�++��:xG�(�ا3��:h37�F�g?U��(|�X�z��f�{H�^�G�����z+L�ԅ���������	��:�E��B26@m�n�����R����UFރۻ^�������۪r;Y�uA�nH�m���vCi����<>����Ԙ�C�ށ�-�w�q�5�j���� C���m�}�I��1�Ŷ
��w��qvVmfM��X�Ē6vک��2�8D9;"8l�� �E�����9܃�>��E�D����L$6ɟ��6C	 �mc��m�.��كkj�sT	45�4��V'�t�+��[ ��#1��5�:�����;�j�j���Z�v��6�^��$��5f��_�(\�]�me���<�b:����j=���Ƽ�5�T�,̶�Ei�I�d��S���6���o��Wy��ް>���;@�� �}A�}>��4�����:���R�^^���X�!����Q'��q��	%_�������g +I9G�[]ك����ΐ",ϲz�������5����b�k�z�W2����ș����#Y�o@q������O}��{�8=}��<N�P���q� �?l�*>�!��R�Ե^��WL�%�����$������كӳW�U�����
��<���x��	�������Փ�:Nj�iȆl}Ũ̶��z�IR����Q���4�����
q����v=���mNR�z�eE��x����w�r	��S���(�SӞ��ٻ�2�I'B��6�)n���w����]�3�|A�F������{᢮z��3�333[�4ǖ�Jb����u|}=�n�zwz�{�}41ۢ�w�H�]����=+^�Wm���Z.e��-�Z���Ū;٧oŹ�cz�m���n�Z�z��r��ڄ�\^X���,U�C�{���br��W*`��-��IkY�T^Je�.�u�gr2��=
P;��Y�;���<�">�Ϻ�\�m> �z�T��9������o���U3�n�������_>���u|	5�=W�n�m7@�g:��s�'f_1��s��WDkp��!�	6���2	&���|�Ng@�<s����:m�^�����ܑ&1�l`m��ݞ&�p��[����=���[��/Z���ꕣ��N&��N�e�^���_E�ڝ碤>~���~Ǖ�g}��8���AZۣ>߫�2S�����5�b���^����Ӥ���[�>�l�<���t+%��O��W�����=|{�m�q��q���=N8A��pF���/��BS�K������{:����WkIc���[ܟ�d^��jF��њ�*ޯ�;ڕ���J��3��׋N�E�W�k�~�z�5�='�E&5Q�A^<�����}�7�{N(��BI�(��Ix_:;H�s�D��X�2�hc��v�Ie�oh��ٓy������a��$�9e��y���ص�Zz,����]Z��O���+v�;�c�r�GG:�⯲�9}O!��3������jtI2y×t�҇nw����G�u7C~����C(S�ܗ����#��(���r3'���*��nl���T#o+����7%�������}0���ǻ���`�<�Mt�bW��A�M��Qk��;k��WL�L�
ݑ�LO������@��?�.Q��P��w�u�+޶���۴T[��o[;:�n=�p�;^� �x�{�-v�
)׫�S���<�_z���v�9����^��xVtbܯq�{�龕[���9�Tz�Z�����>[$���sV[�����L�p�+iu��ъm$�n�h��4䚯>�rXaژʙ;��sn%�p�7xC�1�ϡ���n�$q�Cl����o�6���:N���oTa�ɪ� �u�/��:��t�Kλ<:1�tﲱl���a�,{2.�[����f���n��tr�^W)������e�S��PU�+.Fa=��<aXg�t7Hv�ai��(^;�H�����b��8��/�|pc�-�F���,WX��N����u�8�Q8k������3M�G�ִ�a�n��e4���eƫ��q8�&��c��[a�$�\�9[%�L6k.���Ǔx��Zp	�Yj�޴C�7�{݇�{b@�f�=�c�`)u���-��ڬ�(�;¼=ӜS���q��42��Ǎ�����}�~�l���&�,f-o�zn����u���s�V��A&NR�?3�HMx8�.A���/������۾#��	�A[S�����k��2V�&�N��7��F1qW��O�����*�l�r>�^"�m{�J�h}�ɲ���*Ƿ'�AVs�p���R{R�Q��������*�Y�僽'fM�e��u~o�c��r7{��Iy��F@ا��:#�Q��w{���L���b�����DG ���mWt���Rxz��J(�S�/>T��OW�{�3�]��:2%է�*��ʋ��0���jI=m���^?PA�!7�ǠqA~�NmS�[��k�{��ZŹ^�R{���<wӍ��*Xd�B�}$7P��/YG�Ď���#0�Y�=�mDo-��۬�6�ԑ�����pb�&��^�I�˦@�E{=���w�dh��	Km��q��{k�4�hf}|��(������:��θ��ĉ���Y	�H[��u�|'aavQ�����}��7��\v=���v|�A��M��^=�=k~��\�4?U�ت�ٖ�z��!߿���6�6���8C�󄫬�3�C{���©I��}ޗ�dL���Z�́������>։t��`BfC��=�e��G������Ķѓ�����c�j ����9�v�9�ѫ���[���&���Ah�u����׽ ��1^�ƭ �s���^@�{*�]�)�[���E2zh�7�|[��1|�O�x���w6�[���o�{9�OF�Gd��N׉�F��2�ܸ�ka��'�qs��L3f=�ѭ��4e@���k��<��Y�O����9gzMb�ꂡ����x�}�
�x��Sη��|���t��40�	㻇^�`��P~��c�{�GϿ�>I�~�����|}�����Ϗ���������>�o���<���=W�I�˕L-�Ӈ8���4�C��'��Dȶ�V�n"�t�6�u�<�52�Ļ��Hk�#��N�]�hu�y�&E�󩊬��f�X�r���	���}"gỬ�sPx#���ƹ<'!���fv��P�*-yI���%ӗ����L��*
ï]&�W�LX�fE��e:��=�g��{�M%����9|T�t��X#x�jv�&�'I�/�9�s�p�c6����a�&�Yn�(V���cEU�Yq��9w�+��.ˆ��vGɎ&�}�R8�W���ے�]�8�[�)�*����ck�'WED�.A���쩔Y�z,��;�$�����^�Z��՛vՐ�fT��9�VsͲ�^k5�F���:�Mw�`D>�)҅���7@�ۡ���l-r��	����h�W��x�1�Q�ܱ���_;�9f��	��NZ��Y���\�w�-�q�'l]N �n�K��V�(��6��.�T���]�n��_q���\_��A0�i�-�>�T�I.Sdo����Cw0�yz�����r���'�v��-u
=��U��wiM؄��w@�_S�͎��
��E�Ii������'!�i��4Ł��/j� �o,\��$�]�=7rA�S�B�������E}�t���\
VE��+b�rܜ_oW9���;�/5�ukb��3qmo�&�yx�mQ�f��Z.�|�{�m��I � ���!�8�ޥ�
�����\�ȟ]�����\�cm3���j�������[�c��fQ�+@Yd�1�gf
\�(���\���W���]�sI�*}�"����r̾ͻ��;�w�:Tz�(;%��0[�/_���ͧ.��I:Ե~B��(U�$@y�ܛB�)�в����;�����j����T{a[R��V>�J���k6���V�i���X�V]$ɗ�b�q.7y�͓2�Lؘ.�\�L=���ms�����D[xG+]Z��+�p�\2��+h��6�.�om�_��Ү59\jo*�4��૚�&VG[e�Y��^n�W]>��[��l�`��a���^l��),�;7�nd��F����tNP��;e�$�I9[����²�J�M�,^��&�#��ML�v��&�!1z��p�g�ڌ�~�yR3b��]©�#��[��U�0j�9E���p����E�N�XꇯJ�zבͰVgau|��l������kt�WIEc����r���;�[��R�]��)e�̗9q�V��J��\�4s l6�d׵���U�AvM摲l������ i3	<���!����vA�."����O�l�L�ݒʝ�K��s���6�J�yn�S��5tA	��lK��Y+]�\�I�1��Ï>{|5kR��_l�eWh����E[���v���|,s�!��j�v1���̒zM����[Arq�.NI<�e�U���~��2Ȋ��E6�h�b�ITD�jw�j��QQZ�5�ڴm�Z���0ZT���5TF�b"����LQU� :0N���5D�;�Q�d�)�Tb;<A�QAh���-�Ӛ*�`�EUucTWlQ���tuD�%KZ�q�4|�ص����"�m�mkTT�DA1U4V�ڨ��W�����Qٰb����U;h��U)�oS�����%1�h��"������(*�"�*�M(�X��tt�1Ht�D�TUSk�`���V���Q%�[�+n�*h���v���t�F�q�v���֌U�-ۮ`�(1lLرEضw=�[C��:&*^v*����G�gU�Ψ�F��n*5�EV�_]�DLTPĆ�Zt�TQ���c1Ewq�#`К۸7`��k�n;�n��ͪM9�!���ۊ�z��h(�\Z��jb(�e�|�	���l K>{��^��m~@ʴ��LE"�k���{�����!����m,wh�f�V摤ֱտD���jR� �)�g�K���|~�\��y���s����2����g۵���	��5�_w�ů�>ZK#��b�Ճ%F5s��Ow*��A�C�F���s�T^=�#w3E_I`h���r����Ԝђ&�g�?��|R�7�:�xv�$1h�v�\�h{{��3�)	�."�RR͜A�z�j-�g�y{��d�(%\X��<t�Wm����,����l	w@`qm�����J�`��ء��!5��� ���+�ɫ�����M�G#�����>��,�u�9����80_��U�@�� }�dޑ��DOY�ƹ5*�diۊ�W�w/�7�@L�Oi�W��Jy�6�kKJc���(!xW��f���әT$e]:��;z�����BI���>9�N�t�e^IR`-�;'������{�Q����-W�7{�&le	K7W�c�����;��O�b��V �"�-�Ú�Lap*pQ%�nM���쭆��f���9��~h� �}1��}�<�Q{T�t�/�ŧ匤�d�k�E��B�������u�ٽNP׽�a���l�&�v#�\<2נ6�i��j�k�a��y��G����ʴp������9�,�=��m�����^>��r����l�FDTjΆf����%@�Aipּ�ذEK^��eƍÑ`��E��s�N]V,E�+��:��1�[s:60CJ�ӳ�t���bto����Z���d����4��o�a��k�-r�أ��|w&%ݘ�c�t!w(��w�	��PSw�oT�ܙf�Z�H�Z���m��o?ܺ)��p{�2r¢1� �H|�6�`3��οn/��r��7����L>�-m�$Ë>��'cӤ�sG�6����5�5��|O��[��+q���:��]W��qa����k?GTkݴS�i��
�"�&+����1�~��o�����[����X΁L�i�����7�#Y+����ėme��8�w�ȋؖ�n~�K����e\��%�G�Y
�!;>S�{��B���>��Uw����YϐvJ��~�|�4?j���<��������/A��.�g)i�C`���H>a[�ߔ��=���Ї�u�e���~}���3��p8^��%r�W�3��3gV@�t�H��\0��.2��y��zor��#��f���蛄;`��r�,0�z�YW���z1���쨸sV�`�!��&��W��w�+e^�u.�K�BbS�@F�g�-�n�e�~&):��Х~�I�5x+�i�p釧�ۡ�]K��)��h�Dy�7�+����4��\��DP���߫*��P9;8��y�R]G�,"����pbwa��e��y�n׽�D���dS�̌������Dr,t��0�]����N�	�y��pjf�FT��&N���`ԧ^����y��:�U=�}R{)BN3��I��:�ܭ�*�?�������mw#�r#òso��2Ob	e~���j2IqM袸lN۶�v[�%}1ݙ�kX +��ǖg���4����x5�96�<���ԩ2�0�w@�Њ!_���T{L������G�>�~�བྷh��wȳ��݆o �sL?�S �y��,�v������;�V�Z�v�ǥ�6ĺ��4�x���J4σXѓT��vy6ּ4s�z�W�����V�V��0�:��K%s�P9�M��iIcH�C	�xwf��|yp��>`鹽�K�h$��ձ&����u�yN�F���:�`�E���~�]i�Zhr��9����9ؐvn�m�ڠ�� ��@P[��[$n�`9�;��+^҂^�K��N���!�C黱}��f홚ա�U@`�#��&,᰹Ɇe������,�o��k^Ɇi��n ����+_nwK�v7��UgiI�:>�(��C��Cߦw�ay�Ӫ�ͧrSxwH�p孓Y��\�do"]�a�1�3 ;O�����uLx� 9x��'߈NG�v*1�q��y��*s��O�<"��u�P��1߭������%�N��EBs]�9������aW���N���	9���^��]?]B�k�rC9'b�T���ӟ>��u����u��Y.+)�r.�:�Wh��1/n��T[�v�K���+9ڔ��ɡk�B@��W��-;xc��l������# ��P@A�r2�'D[*�	��46#���2��㿃���ǻ��)3�7�z�:;��k�U�k��Ƒ�C�P���W!
�k�o�����go#��R�*Z�3���������;|��t(z��"iZ'*Z�I���a����WB������׷�ç}F:`��aV֭c'��U���xZ��C��ig+v������6_���P�hRp"x�K3�2�n�_#o.k�y^�a6MФ��=��Ip2$�e��Gb�j������F�S��N�U�K,�N�-/��e0M/�Ҫ�!+�p�����
���E�8!<�ހC{c�O:�gh{(�c���خ��j=-��P��I��U�&�\᪢���H0͎�� �(�aeR��;N�;3��6�j��r�D�,�=�E�Ԣ�tS*[~7-�̽�0l}���w��,�f`���<13C/G-�逛��P�xi;����^�9��ҀO�o.�R����]���9QM�
q�Q\rOn����}pǝ�4�Mb4Al��o&�m�,P<v��%Q��Gs��t;��o?�@��=2�*�q�?0��-ZY�����Q�C�^CƲ��p����9+½���`K<��zHݼ�g׏5�
�X��>���-�	]�͆&���]>�u�y2��\n�8��:�d�4�Z�)�Jr���9����:�8A�gV���S}������O��J*A=����y���]SبmQke~35�,��p$p=Y	���M�۹<x�ӭ�֒ܳo=0]��(p����N����Y|�󂁫�`�^�B���Wع�{^>�S�עfy�ǲY�5��ɀ�぀�4B/5��U��p�y���*��u�z�T��������Hf�Y%?Yx���H��	��^x���-}����]�-��:���Yf�z�-������@DԜp,*���L�1;���wA!� #��i ��H؊���Q�>��NGf�G:�c: ��Z}�AgknO�Qx�pwP֝�4�}%��U�B��K�����pc��vޓ/^t���k�e��iʈ��0�)��>>K���s��Shԕ3m�3:oD�01�!�S�����w6�s��
��ڣ8n�TŃU�*Y�P��1q��X��^ �m�
��b��3��w`�1@�5zњOŰ��Ƕ�>�w�|w��,-��	����-�;�qm�錄s�Y9��&%�{	�W)Rk�Dv>5{`=7f_�B�)]}��G\����)�$��[�������Ddڸ:r��}
8�YK
ǒ" @m�7�1�S��7;`��x��Gf�c�x������Pn�d!Wn>��=rkh�p�n��3F����u��6�y^��u��q����_�W��_}W�>�(���vݛ>�L�cHB{$���Jt�ħV�E2�RJ�c\vN����M�E�p��e��-[���.��;��T�3�.�O�$Î�2�����Jඋ`,j��K�BVp�N�^U�g`��G� >�������z���h�����uL4���/@���rb�����V�K����m
�Vu�',��x0vo��>p��r��l�v?|t�z6����ǈ9��V��x́����%q`�ÃN=���,u���n7��:�Le_�6��u��{Zmb�6z��I���&ޭ\�T��i�d;7_C{�n/�U,ͣUrz�^��<��=�o:2��2��n��[����Xu�e�`��W����sH/����;츌D��is/���]����t�ki�=K�>H�Tk��po��ƭ�� �i��_�9`22Ȃ"C�j{�[��5��y�C;:���FyJj�T�����H���s��4"�3Eی;���a���UA=������˯����M��'�"��YI�e����������m~����f١����Y�(z��f���ʛM�Ϲm��x��S11	����=ϹEۙ<}��O�~�Za��kҒ��ש𕪹r���e���y���"���
�G:X���Ιs]��;������}�4ղ�a=F��;zU���b�����:�P�^s��V	Y��4Pf{����� �7�4�˾���"~�c��g�C�Ir, &�=���*����g}�˴��_�\�o��H�x�`L�#C�["�=Us���E;s]��MI�[�a��\�q,�X��bz-�f�2�dgO<�����'*.B&1��ݮޜQ��ʐz��U�PB}ka��P%� ��1��c���*.��f�+�U$�8�r�7�����[��(2��.:�1=#��fg-<ɳѰs�~�c�&):�dJ"U&�d� {OBzή"� ��~�͋a��9�$Ao@Pe��a'�=�v��	���$�^�Hд��7��H!�e�l��߮!�y��'c������c_|�~�6�<�������ƹ����F�)+�'#c������8�\�	&������nok4>6����}Y7�u5��$fv:ј�,�w�#��C�׫�{<���)�I��9�a��/��H��g\��C��tJ���\�S�4ǡ�On~{�n��?��*^Am&G%s�W�\��a),k��Cx&��f�w�`����I�,���J��;�Dc�R��Q�*�$<q[�UΞeV�����}`+��?��f��1k������9;q$I4]D^�f���r�{L�dJ�][��!��`�Z\Ű���W�P-1n-;-%��s�$|��u��EN�U�_:-,8��f4�����Dȁ���,o3��+YrXey�t�9�^����������~i��)J���>|�y�,�ۄ0nM_0tɤ
9�z`kd�n�2u�Y~��iA/l���5!���
M[V���E�_L�2��}�:�g7�9����C���XsP:�a?Mk�U���bv���̞,���j[X�.X
�"]���4Ba <F����d�n�6��o�X4.�h�x�l�cgWb��'��r�c�LC�l[�¦<F�'�_���o��V�nD�;KXnglv��D]���w���o^P�Hr��n]ݡ�y�xe@lg	oR�#u�u]�8�����s̽c�f�cNd����
�W#^eP����\'���>|���Z�o���N���χ��#���ܮR,3��h�!k�� ʅ��+	Q�ޘ�V��Wc����%x���L<ï��g�|p�k�~��*ea��q�:���d*����oe����V��n�5�4�r�K}�.�VMФ�ח��
<[˄���=�y�Ep����B[o�^�]Ach׎}II�gIH�Ȼ}��xU��v�!Ŵ'H>T�!?�^>��ʝצ���k9�-XI�F�d�����ߘ,�7�8b��2���P�;�&:D�S��p
t����䦅�c,�}KA�;V�ޱ(�}+��Dx����Z��=U�]��B���N�m�b��m.]{7:8��� �� f�[�t�]l5�b�e�fRu��3L���I)L8?E�w0��5��f���|�Ȳ���Bb3�����լ*��)d��J���(�aa�]`�L�i�n���p��^sf];?H����ݕ�;!��Y��A���z;�<�_�N�)�~9���PX���f�j��n��ճ����G;����<|ɵ���v�Iu^�Qo�)yժ�\�2���uO�J"�xͫĢ|v�9�ݕ���+�_:P�^�~�􎀎~~A}�i���~6~��x���wO߆ѽ�)�g���a����>��:��w,�^��h���1��Q����������󭁤VzXm6l���X�v�� d�1��:�l����&g��{%�׌a��j��p56��"�`�����e�v��w�;�37p�H�O�^=%�h_����xt�/ϊ�nq�7f�R�ye^�+7��J���j~?�^����~Y�h1��@cn�$>�D'��b�)ǵCT�J��g�3��e�W�%�4F�����D=�	=��{9�CZF�f��X*� �����ө�"nz�2�vg\g}��x��@<����Xy���ʿ\���Cj룅�
�<޵)�AX���^!!�Ш�Ɓ�75ɝ���t�qY�j�7����y8��(��Qmn��]m�#�؝�r��RK�]����TXė�;�#�?����������(��@�	�y����-���6�n+�c���#�Y��0���i�=�������M+;�Y��&���ʮ�w^y��ț��ٟ+�X�ψ��~�Hb̓���W�V0E��Þ =��#�5��m8�q��	-��d�h�'�(�0��ǡoV�^����P3�or���j�%�u��ZޝB�u�FB�/���!8�&i�>$���R������L���	�aH���Y0s:�7��3w�Q��N��0��iOb�"��14�;�讑L�-��� � �L��&�uZ����5(���ڄ.�m�Lpc=���I��F�|b�����I�E���r�hY8s�mvo+a���w�����4l#���b7C�ݷ���S �&�p-�Bǩ�Jjzv�gv>�/��n�K�]�QB+���|@~�0�`e��i�p��n�R�ؖ������Ğ�v���fz�3��?Ј$�o�r���)�}����[x|{a���[	��Bq��?�fY3�v�w$�#�y��r��S*I�j��t��b��6�~W>��^��ھ�}���執�����>���~_o�۟o�����||~����Ǟy���>�7j�-��o�Lٔ���FS��2L%(���w�J�-�lV�D�5 G*Mr]" �����[JKA3r�u�W9ɪ�캵�rf,ԥ%q��.1��6k��,i�'nP�|	�DL��D�L�wF�{%���Y3/J.�]_6���x��A0�C7�DC�M��2�5�ڥݳa<�U��i�3�%�pc��-�&)���+3��uҌt�z�*�9��-�۹�s����O)���,�b�]��X�߱h	ݘe5��.巚l��8�0R�C�f���K�D�����mU+Ĝ��+h ,���K��{����X$i�W1��G�7.\\��&�f�0�s/�g[���sMbƱ���u��k� �ɺ�5ס ��&|�n�
��VN���;���'u��c���a�k5�or>�,_K}A�!i�.���ms�K$��j�uS�*]�ר�V[��D��],t�0��+wO<���QW���Jd����"-��T~�R��|W%L����6�[]��-v�f_vV���(�vh�H�Yщ�;�8���Ȭ�+�KwY�*pc���&\ut8敖�{� ]_e�G'����F�s�E��k��j,�{L��Aw������T��F����$u�4��ck��2-��Ѳ&`k㵎v[=+$��)��(�=8r/��E�GGq�+F)1_bP�1欷lo\\�*�G�9��G9<��]ˊ[z��p���D�5o<�;�o��ڿ��7��l�ٵ�Ma���
��>�˻�
�q�}3��w`��n�7�tw��X��>�K�\�Nӭ3CQ�[p̦�d�>�<�O||,�8��^�'L��Ҹ��5����|��۬é3�"�W���(q�2DJ������kɒ����\:9�r)��÷�o*���&���N�!u��׻��X_8.Md Y��(fR�ݧV��UZq��Z�摽�qS#øE��]��t���hd&�i��9��vu쿂���9㬡-����9�p�S,C��N��.�4��4,�%a��:�N�3P[�U�'i5R��V��Fl��(��p�H�;ML�wK�[�1we�,k,8tL��!m*y�6#�Ma�p���h�
�l������P�aAJ�<r�i��X(.��N���������-n���v�k=�XrE��<x��h�������R�Ê��ai�r}:]�R����jD^����l �+3�YO���g;#-rMXN��L4�A��Khl&�6"���I]2v�y�_�0���ҕ6y�W����;N�pSI�N|*h��˄_7r���^��e�/~R����;A��;�-=���cknuZ�7��BM��h�yw�/rS��<1{�nf�lE��S!vv�f�Ɛ�.4���"��Q�Q���Y[fs\b�o0JM��9.nI7�I$�������}�vld���`�]�f*x�������q+���]F�EtrOv-��7rV��8�;kF��ZM%d�ifִ�m�q��tM�k�J��46��[w�tE���q�f�upa��4a���-�����;h�
֢x�'���Uv��{��/[��\U��\]rGHtv�7c5k�7h����0Wkb�m��GF1�F���m]b��g�UEyk�i*�Mz�n��,]�*�;�F�\�Ǣ��E��͢9�љň��TU7���WGCE��G3�;d�F+1�pn�F�s�f�t7lG]���\OOlS�����Z�޽c�"7�Ѻq�혩&�p�m�m�zM;Z���;n�����.8㪩�g��TQ�X�#�v��7kb��E��7�z.��]�c:`���T�3D�+��3�Z"��Kn�4[����+��vϨ�Q� �v�b���B�"�3�kE���*�EL�hV���5%��\ELm�щ�������CAz�UTz�%f��^�]c�:t���޽q贱o[��)6�z�J�}q�{��j����T���������(
z�=�'ѷo�����|Y���h4����<|��=�� �YFဖ�&�D!��Er�[Y���&�g{ˠF#�v֞�*���x�FC8G��&v`Z���uk����aqR�������g�D��#"�(�!��m�!	X�$#L��l)!*F��ݮ�n��׭�����
AH�@�E��A� ��>웅j�;G�U��ٽ�Gqֵ��˖JI�vп~4�<�j��:��΂���Ë>�|OO��ƫ�K���Hwnoje����h�"��Ni����43�P�&v���.��|7���s4���:��=pL��2�̽*�z�X��V���yឃ��w��X���k%}��N�L�vo2�J`<#ruE�Wco^��\4����؞�N�C��4���,h��8��}c�a�_���y�d^�_c,R,xK��e��c���{Y0&@��A)�A�r2�6�֞�<���� ���9��l|Ē��(�k{=M�S������Sx���*Ɯ0�qB� Ũr�W�3���l�dgO<������W,ϯ^y�C��Fe~s*�UnI��v�nż�n�!>��ըʒ5��1���2���{�RQU�,6k$�oN��/e� Έ�q�1:� i�d���\�������1IՌF�+�I�)�g���򚣥wMfgMeuj���#[РȺ�I�r�`���
~��=�1)�z�����j͘���t+�Zj��+ް�ѭ
��7�HQ�>�(�<�(K�e���v�����f���_�0G��d\2�K�xZ�E�r�ڃ�mû���v�;ʰy�����%���� ��Pw���B4���Mh7�6̢���Ί�e<��i���@��>��V"��-^�ܧ�ۼ�;��2Rz�y׈��v%�TK�K���\�J�Vv��E?��@�J- � RR*R�0�Т��ϟܔW=�z,�h�����"���"lg�w-��r DcH�!?C�9�����M&n��;s��>�܀��!f��'�)��� \sr��6�zk����Z@�g\��$��[e���eY�9�s��zu/)�F���vS	����T$��Ib��0О�nC〹.f��*&��Z�3gv���W�����^ļ�5�,ى:��RX+���K+��~`4�1X^jcn+�Z��@s�R�Xnc@0t�y�B�c^�ٸdR�9���Ng��t���ϻl͡J��*���WvZ�t#[Z���4?�����#�ѩ��2����֡ڕ�C�TD����y5:b{��/9Ŗ,.f���KkW�@����Ɂ��<C��P���s�:o7'��ׅ��������i��l��Iz��^��f]��c�)��y��."tC{�ok��~Tc�_Gr���x\ܦ]�.ÆdYx����TG�v����U�:���-	��:�u�oP�-p���ߚ�2��/���cNd�� Az�W~���5�1�����������vi�ҙ7��[{H��\�>|E�nM5�	0c�t�dР���3S�z�2�J�՝q>1.<�V��pt�[�8J�M�O��oj�4�%�,
ݛ}�����,����u(fl<�0X�1� A	��^�͉<�L�fp7�N��~��끠F��!@�V�F�H���	bA)��U�
�>?�����?�� �W�4O��od�5՞����%���Q�]s�-mZ���xaV�D������B ݞһ'�mf8t/gM�T>��>��0G��5�3����W��y����6xy�De��X�P�n���gT�m��߇�7����v��v�0���m%���zc��۟W�8;�^��~]�=��U��9� �$��e0L��|��Vc��`��L�w"��ڶ5[��M+�8�3�u�9����b�O�L��c�:�:Z��X��ɴ�L��ml�D+�T<J�������gp��j#�.xd��=�F	�.�Z5(���T��7W�r�mB�0:%97jv�v�g{PnvmeAC1i�!�uzc��Oa�F�N�⮗��O�a(,[�+ɳl������V��S��B�u�<e�yC-�"8F�P���T����ZJ�.B%'�wܨ�K{3b{���|�Z�ŗ��9��8}Ǧ�-���k��Kb�-,��T[#g�o=B�uFuv+`���y�r^�ʸ�n��t[Ӡ ����:��:� o����^W�^�R��i ~�se%�u����E� ����(Kd��N�G��pTrU�,�"7�*f.ւ��T�#�������y�P�,�SA���� �4fB.:V�V���&��<�۳F����ʻt��-PN�Sf;���ꯓ��R`h (i(U��R���JD)(A(EH��Fq��ϟ~�=�������if��e��Ri1L�.i3��%���3b�;��޸���~q]L�\��nW��G�Rs���P7�B�t�yo�~�^=%�Ĉhb�'D[��Ž�R�-s7*�Zj����X�za��\LI�/`mFozЕx2��X��A�D=x� ��N�6��8���3�LN��@C���Ǒ������sld�7hkO�p�4U����9���Q��Q�ή߅����\^��,���,�����G1�M����H3���~���؞m^�uvZf+I�hZ�`��G(=�|�b�@?���5��j���V��{^�4wS�S��^���Rõm)�W��)��A�Fi=�Q����ݹ��Țy��^���-ꨰ��ꩶ׃X�#h�hZ�P�	��Ak��� �Q1,O~H�2�J�]�v>753�,o����j��9���_.w��5tIvl�� �iH����>9�N��~��))ML�M�Y�rT,���,����_O��B��0T�uL C)�`� Ì�i'�1I�_����a�l"d ��e�`ʜJ^�+�S���O/��g<����wsרʹ��eZØ'�D�.�����S���I ����E�f7j2��+j��Cz^(����#S��.K)��������Y|�,RW�nM�%�o{H���8:B�����������i h iU"F�PfAI�ZEB��G�o7����ʳ3����%v�b�k�h�ȅˡA�i�4s	U�V����ꦠ4�l>�E�� �G��M�1��r9���S�V�-YhƝ��)�꘮����m���\�S)�.O#��z<��[���G?���+S>�E&�!�7K�gcM����jAl��^Y#YK�Qܫ�$:~q"Ƽ(����]��p�A�pנ��̉�Ύ-�{�B�RuAT��>�=X��?0�M�_���4��B��ٶv0�l<���IU��	��8n�����ݘ��B]��>�2-���@�k-{�=>�3 sh2��Ǒ��#�>���F����D�;�vLR-�b����]����A��m#�`�i�x� ����Xk0���û>���Ͽ���Zo����8>.р�i0�́�#Y+����<woUj�ǡ\הv-܍�K�=.�Ҍ����*����"O��/�-���u}��G��y�x�[�a�.˷��S]c��5q�������� �#.�kM����Z�l���I������=f�h�d���Q��[5ת�}]kkF((8��1b�d��g�f�2�|�K�%�7��uj���^i��G��f��E��_����"v�ћl��}&�
9���("{�G!�)%ׇ+2\�f�l>Ϡ,q�����P�׬��hMTڱv�V���&v_��n��Z��=V$�T/F�P�u�F�]���E�$���û�f���&��}���{��<<O�J)H��Ā�ʉ�*(�*���������y��qC����L(LϮ���LE6�!>2a��C-A�z1���l6.��N��tn�d���7PP�Y����I���.��<ɨFBosS� ��1I�#"S���5���뽼F6{&wa�׹Ӓ��Ql:9�Ϲ�
��)�V\&�/Й'a�8��/2fE��]Y��69i@AҤZ��T���GN0�vE�*���$Ƒ�q0��|6����)3�&�U��z���z�P��sz� �&(d	.�&��p�6S����שr��~��~U�"|�D�^m6�^9�8�(�Pݓ=#˜��4���{^4�ƌ��'�{�bHi�*++����\���u��<�М�Q�F��aG!s�w�\�Qp��4��0����zIOot�7��q���4���m�tX/^��F��$닰J�t�*�u���pQ�=��6�Uv���s��ʩ鐷�� �ʃ֯sԃ	�1�͝�E&0qƒ�+\��\S�����lKw'��[Q�$��֮{�=��~%~��s���	��{���x����;����q�n�ã�Ԩ����L4r݌�L��)t�c7[{��΃��C!W."��f-��e��)������Rec�a�+�x��5�0>G��q��.v�w�9�2���FF�r�.Y6�z�$�W�8����z���������^��PP � L*� �BP�# H4�� �(���~/�W+�Y�ὮEctN?�C4�j[��@��^�9�"]�Z!7�y�6ߛ�q��'��cҭ�+7k4s����[���	y/޳���P&��A��\S9|�K��7�b��iٳz[5Of��μа��<�
*1���;2-<w@$?�w�z)K�{��o<[����&�'Ex�Pz���ή^ȍ�3����F�ڨ�{k݌īCϥ��  �r8P���,��(<98O_�=����7v�;p�����|�,b1��2=���w⦠j7�ʖ��`,~�2ot��˴�mm&ٟme�໧�k�kp��l0f�ܸr(�9�Sm�~hq>���>���Cr.����ʘ9Z�/3Efꎮ���&BeBѡI�J9B�Ǥנ1��E=�� ��d��8H?�����p��1�S��ODj��h�f(Bc�c�%�:&E/��z��	��
`%cm��LGvj���,2���` �@X��3��t�N�1�d�L����%)�ؾp�Q	�����i��[�*i[}�w�T2.�}�9=K������%vI��vEM�hԢ���-3���{<Gvk�+=T�t��շ�\YV{"<]���֬F�NS�%�r���سٮ��o32Z�EJ�43�=+j�#gR�;F�w��:U�27�O�8"Uo��^�b	�]�C\��*��Zt/{h�ܕ&dJ�"\;K�V��ԋ�Ǯ��0-t�/���-�W�����|�O� $�)@�@%���ZJ)�R�H`J&��������޸ËMJY��5�w��LBvlg�巽0t�p�	�O���Xd����XM�5�<�я�M��юsO��#)&O��#��G����K�ʒ��;B�ٗ<	�D�g��U��w�#.��4�Gs��@�-.{q�������sL���7�ތ��.)���h���v:s<��t1A/t��9���6���������t��Қ]�b�G0�&/l�ٗ<�o��_I��3��i3��%���z��1a����3�*š�%X��]�n��g#������/�P6�p��\%�^#�\����:"ذ]oɢ5�fc����˽�;*%�y���S�1�k���t���dn�0�C��C�poU�[v��"������.���-��m%o7ι����(4|�7q+d�Y�2v�����~O����No>q,
��t4P�w�y�i�m�a?ԟZ���L�Ѣ[��Yz�-g���SN.d1q�loarҊ`X��y]cռ*������E��7���g|�"�0�/Bti���8�rڮ��G�H�K\��md���bb��0ko����qM��d����h���u��Ɖ�K	݆���#�:䧨���U�)��\N��4����X�N�wrQ5��V(R�ѿ;����������z�w��HP�H!$�,J%	0@H�3"�
"�w���}�>|�?>}�}�~>�}�H�b���8���=R����I��~&Pd��4��(�0�z3/��4�_ ��{�S�n�T2�v^B��י���(��S����dQ����N(��I���(JS]���ͻN�9݋-���VsmS<:��� ��Q<��BW�0y� 皽�F޼��'�9�N���*<��\䎈3Yii}���R��F��Ac������~b��;Q�?v4G�!��T���왡�ƥ�=��0��p��jc"��,9�p,�}�ǧ�<0����?������?$%����TF�v۾^�<��ts)t���,��ǇpFi���4�>���gl�W�O���?}D~eF�-��޳���`ٰt�4z��/'�$s)p(��zO���v��v���C��m���;;��t;k���O�:�S]{���úJpZ�&ެ+��cb�ٵ㵹X�3{5��[�V��n^E�uh�!��c�(7�ZbKoP1�^�'���j����z6&^��ؕ�ʨ?���61���?7�o���I�����7#��<��^>~��]�M�D�|�
�g:ř4�Zq\�iL���=wf{ ��J�*&�N�8]B�3�֫2�:�oZ}m��Շ��o��C{�������X�����$��)|�gU�{����4ͬ����
�li�J�����8k��s�y���_׽�^�� �D$A�F���$�D���ϯ��������}}�N
���δ׿.�����O�c�LL,s~ڑ���Pnv�ܜ�B�A�!����٨B�d�;W�K�i��O�����?�ӂ\��6)5�����-�P^�7B�S���Bq�֮o>��}�����t�v*}4�6�F]�[�Zr�O7}B��h1�;�.�}ݘV���Q�ൂ~�c�~��ez�ukN(�U���ŮU�A#8�Y�����O���8E[��WA98`�r�t�F�<�!��W�nB1�4���$'�5G��Q�,��c8�`��?\NU-�7ol��\:�[�����S�2㜌��ƞ?�W�B��p%:���Au��в�%��b��D �BUc
jӓ�e�eߧ&��s�>U0��Bˁ�Bێmm��۱zd���+ut_l�A�$�X	/+�'�ӌ'ò ��]8ށ �4�#�B^C*�&�HO����Sp��tN�7֌�|g�L��\&�n�I�"h�8^���H܁#����Ӑ�1��T��n)��y��S+UCIʕ�V��"�<�4�Z���4]���}����>�O���|����}��}��o����}����|~_����ʭ��*_6����5)R�R�m\ޭog���GhO�k�rX�we;����u79���ˇ!� �9�w�h�ú�[��m|£Պ��@��nSW#o�[����Ҿڗf٣q����㲘۳�yn�]2��Զ>�ؽt{+�9��*���U�{��y���FSF��"��6�.#l@�����sXP�va����m��&Rs������4�"�u�Qjq�9�z(�y�V�m�C�]�#FZQ�Xz�uu��D�u�&=��D�t�} w��/�t�,OR��Z�٧)��@�]�]_���huc'&0\�8m�1�J�PJl�
ճ+G-q��/Y�XR�x���)�ˬ�\8ň�r��o�q��|fTWXr��[�*G\��'�Ɛ��{L�i�=��\�aE2�d����u�9e�ԫịq_mӁfHva��3�i���lZY����t�_R�	�B�r*5��b5�"����txieR�}27��\��r�&ObØY�◠L^+�a�z���)KOe0�&Mǥ�w��**]t�ɻ�ZO�}d�)N�����$��4۴M˶zme'�7d��t\F�AQ�|����cs��Ko��{t��O�M��K��GnL�+�t�(�Τ����PY���>[B��4U4 ��R��\��;�7����%wWmk7ӞS�<,bWZ��#.+!�iۃl[2�p5�4㏲�4�V&R�����,&������"���۠���uSGQe�'��N�Ƀ�vKçA;V2]�q3�n�Js���*!�P]�6�e��d��t�kr�6.M��r�;�D,l�.9ۓ�o�ÂV�/2�Z�m���>��w�i'�`_�q�,�_A�S����L*�;lÍDK��9χ��7rP�-,'l���������	=��% �5}CB;�;J��Y��9��u҄��mY�ZhX�.���=	���cF���c��ܣ�H1�$�*[Ϫ�+�F�	�d���CWPء%�0����wcf:o���S��y�Å��&.�_k���V�G5��ve_��c��A��͎�Ǩ�ތ���T���H2��&tR�.n���K�z��V��A�K�ʻA�&�GA�XT&���n!�R��1����@�.��F�+zK;�#\��Qn��|1�kU�GQZ�<Kzn��es�l)4}r�<P�*d;5)�Fl0$&�'���]9�u��5�oռc����l�z��C\�t�çy8���2�,L�wX:��Y3n��4�;EjP�jp�U�ؒ���A�Jm��r��ڕ��W}v���t��ʂ�4=�(/D���g��B��5���y"���Q�恜o�+],�i�L�S5e��k�f��Ǔ�m���rI���H>����g����t������3���i���|mTLU�T�tj�KI�;X�kZtb���G����[�rU��m���z�i��mޱ�8���:C�4z�S�PW���Mz�R���T����ֆd��kՉ:�%4��AA=EAELQLEU�q)[f�v�&*���B����^���A�]G����M�X�Aj����U�Ě+Eu��Z
H�E����m�X�ĥ�	zv��艠��&��Ѷ
K^��7km���:I��:2]&���b4j	��фꖂ*)���41��:��t:�:]	k	[�⊤�z��vh�I�A[���T̑ؚ���t��Bj�b���i������B&���m�����Bkh�h�cZ��T��)��#X����
��"h)��[�4�TT64�j%����m@$!�||�}�ɶ��%���Wڪ4����j�u!����s�A|Ah��\䳿~����FY�Ӽ�ƽylCjn����7ڲh?ׇ���� @>��a	A�" I B�I������a�*��|`���8�wb��A~�2'���h��,r�'�	I`#���"gB<��ח]�H�ff���,�#[�76���;%As}�`Q���.�J�¼���U�Ӎᝪ��܍�ܮ���J�DRX|�7�ku��>��1�05�w�+hێ���8d�3ݧc:Q�oG��Q�'�4�+	t��\��~���N|�P������jup��y��]��8�q=@�	�k^ǉ�i�&���Ǡa>�/��̃"]���	�uuf��u=kc�}S�?Pݖm���1a^&$�v���D��ޟ���<Ft��<����gt�i�hZ=A��o��	�3�78�w��vdYx�wH$=�S�P��ʬ`pB��K�W��ۘ��1^��%ğ�ϙ�>�H���'s���A~*���nY��%��C�U���fN� �E:�k����V��F�.Ǵ�d��O.e�O�/>�kjQ�	k�F�R�ˌ��O�9Tw�k�&�ojD�:��zq��skb��t��0La�s�(�'�{|�ܳ;��nR�=c�7Q�o��ۡo{��J���g^YŤ��3h)�Z�Z��N��$[�;'i�:�ӏ�6�%U��<�[U�����jX����xCv�|ѡ�4R�p�;�y�����Y��\..�(���u娓���:&mo�x��O߿��ѿ0?"T�B�X`< f��0  �k:Q�����m��	-����ʀ�hR{�r���u���v�����yҶ��Q%�-獇�Y�6�zx�!b� ���D�6ħV��5BJ��l�8�}�����ӒUM�����-���n`�^��NPu^�9���k��2��� �%�u�n�e^IRaO�|��ɊB:��h��򞵝�*%׋�D��>�L=z\���cH��%��vEL/�Ԣ� n�eyu���!�_�&b��ܝ�����d�	��Y�s�c?M��M����aF�������].�Òu��+�6��^g���1����|��i_ka���My�zz����/wbZa�}�͎i��cBtvf����Ϡ���:k�V�?u�֟����k���uΒ~�D���}�9��6�j-&m��
Mk
��{(%�¸�A��m��l��0n��U�J��;������%��Yـeoyfn���t�Lm<u>�3�ע`i ��ƌXgbo2o*vꛓ\�9���oyd�Gy�F��%�^�ؾ���r~,��r	��<|�-mD~3N�o��j��B�k�ez2��Z��	�YC'٧����)�?���;����%tS�k.�y�iOA]��m^�n�v�%5Z�����B��J�l��k�4�7�p]CL�	R�®F�
≆WkGЃmJ�95�n��{�:�ؚ��{��� �����ޠ�|jm�}�T�}�Ӳ�bM�>������y�ށ�L$��ĩ�{�ڌ�K4��cn�$<�_�}v�U����<�
ݗd�4[��"��lK<x�-->C ��{d����l�k�l��l�%÷�q8�z�z���Y�)��Ro����"dW��C�aR5��q͏q���{ۘ��+�����C["��^��f4 �6�2F�>��'ƚx]_:�����{���V�^G+�=�1��2�����T'+w\�W���Jl�L��&�h����#8��z��x/���}��kq��v{��E�/3pxaw聼ul��7:	�&%�{	�V�I����Ǌ׼R��g9���W�mL4�:����46D��1vl�"�	�v��$��?7�S��ħ]�͉�`�Vll�Ի9��R��1	f�lBYŽ��\���Ř��������c���y��	�}[ULd�oh�D�׃c|G��&�R��0��Lav���4[!�"mLp�A_ၛ�*��l��f��bd[�d ��%�?"H%�.O#���?`h�|�F�������*����Z�cڶQdGw
K�o�����)M�5t�o2��kK�i��ޟ�Fk�{2�{fKr���y��|^�(_ (��qvt�R ��*U>Jn�e���-a��SK�����(�]�a�F��\�*l8^S�����'5W��������>�f y� <��0����s��S�E��xd���]�u����E�H�R�}Ӛ�n}�gǶ9����G��&�+����|�̜����"���}͍vr�2rִɷ�W>�j�`��q���՝�5Z����5*�����ϡ�]�v����-X1%�}e����u��!���U����2�2뵽%�>��ԡ��
����<g��~7��+����x����kZ��~9w[w��{}h�����֮5Y敚����A>'�0'-"7�+\��̻��kF���͚�Q��s�4�Ά��H�P���2�Zx�w�tE����l�w���h.9�	_�s��X�Ǧ�.��<������wO���wI.�(��A�r�v�}n��Y���|��dT��!���Psb���dp�aqlSߪ�|�vm�0�qi�b�W(5��=f�2�y`\�NV����k�nG,cN���պ�V���.�ap�y��j��0�z�Y?vclD�C�z�s�co*���O�[M�Ӊe	�
���>j�G���<X��ta��1o�J:e�{|��1<��d�EӮ3ݢ��k%i@]�Y�R�yd��R �z�#���8Ab�\;�3Y���tE~3���/�ͱ}]�wvV[�����SsWcF�����j��N�U%�E��v�dO���&P�t�:Z�i�;r|�:��Š�-5�U_�	@0�P	I@
1 }eu�ű�9����O�S�=I�5�8�/G��^j��H�ޅEÀ���v�H�0�n�9.�ۉ��l������D�V��j��GH�Gd[B��oF�3��q�UgVn�����{3kU�0�C/,3 wQ��	�����&�����|��.7s�IX�$�n#ۧ�l�?���v+�M�:�COeIOV	�d]`�Ći���G�����X*Ę���Y��9�2�]Z08���t��`z$�XF��F��L)d.yn ��=��愥1���kkv��=��emn�;.R8|�|�"۾mm���ޮ�f��B̀bM���,2@�w�^U��أ�]����a)��j�nX&L/"�a���/?�u����f�*�˝١���5��|]km�/c��{	A/l��hF7{��P�f��0�V�й<���-��n����n��P�b�`Z��@�����4�j[����-^/a�ɑ.���`l_s�UV|W�3B�	�3��L3-~݆m�۔��_Gv:��;`:"�bޠ9ų��~h�Cf��Xo��v�tN�����7<���xp�zJ��ȣ'd��\k4NG��\k>���G�{ɢ}�s�z��N���(]_���q�>]x >��ЮٳAv�OԬjc}�0E4g�o� �H����M�}(�|��֙�������߀ �{����<=�`<<���W��Rqvr��T	�b��y/�6*1��oS��ۮ'͂da�a��6�$�|.�u�vi�;yA/7���[�e�ll�$!\LfJOa�0K��-Va��u8��4�}��~�LLx��s����{M��[�>�t�צ�KQ���P��R2'���]��~�y�;&��h�����#�2�WB�����i{���㦿V�)������9ﮎ�1���Sp�=s�6��T��MA�����L��hRp,J9B���&�h��g����k:�G^�=`�ms[�
�cP�}����CH�3�^~BS���N��Q�:JEll�>���y�j"�i��rqw;����z��Z7Џ���_l>T��^{�k��锝cY'Xܽ6�I*L��*ͻ^�i�o�����d����иf��.�`�m�������]0�#�E�^�m�~ܣc�y<V�;��qSjv��yA�-A�6�;�B
��8Bn�&n�2$ٔ�&�:ឫ�ދ�J���V���e9�%�ҡ���]�\>ߘG� �lhI�>6�<x��>���GoiMO��|����mF�aѮ[{+�Gsc;�.�����j����Q��%{!��a����*<�{��pnId���;��jd�yѻl�=�\�r�C-Z2�F$�_m�̲,��R�*/�C��Z�]A0M��4�o�?��ЩH�D���������z���+�zg9�r/7v���w�C�v��/^Y��ʭ]砲4��� �ì0���x�K�W��N��Ύ���d��ke`5�	�Z���{8�W��~�mM묓j��U[[�>mgJ�&�l�t>��vd�C�]���6��J��3��7����׉�i=r�K]�!ޯ�Y�6�3�����@x!��9_������5��q�6�?��)�� �3e�u�Y@�{ي|�[���읞��q���F6��!�ɉwA����%M����t���sv���~�fy�ii14�����$�B&]���N�Muc�0>D���>���ʇS�VM�0�/v�LSL����ӈs!��3E�,x��(r��h͋O�m�����sK �4�
�W[F��P	�3"��o:;�>����zl-���q�(1���\��M�_�#������J��q�KcC-���kNln�=0d%�k�B.=9^�XÕ�v�7��"Sm�5�����z3/кj%�G^Zm7]�n�����`�as	�`��U�C�Ђq@��I��M����"8=s6@�G����6�2V� ����\P|���7	;ok_�����_s �Ѯ�_�'n�LD�9�i:0+�3BR��߂L�v,Al�:�ct���u��P��ԏ-����#N���d�(3#F�-��q7'Q�b��;_�b���w�| ���G�gc�r���|���s� ������]�!�����aC�N= k��(����F�],�Nzs���^����w�<�cA%I��Gd�S�p��G���l�C6��S�vK�B�3�#x�{R�mu��;��<�E�!f��|���:�h��%쾾G�e��BG��D �}9'!4v���'jz���6�HnAl�R{�%.�7K�F-? ��.O#��a��?KE�/��{��z�&ͣ}�Xt���>����k��SM�;H�vvQy��5�R�PK�O�؁��݁n�����sWW�7'���;E��2�v/ŽS"5�u8�M�:z���~b�ɷ�
�y��N�4g]w9��u���Q���5�Ct� �^�;k��%�_7�ZIa�Ʋ�i�qх�2*l���2{��L?ˬ/t	�����.)���t�x�	vO�7�䨧��$]�Y|w�R����
��K�6��rŨ;��}��9m���z��;��Tٕ�Of��!,b�A���"�LQv�2�[��C��1*���V�c��,o�����}o��h�g�XŽ���f��*�R
�TQ0���aY�ҝm�4r3[�Gߊ�����^� w��tۖ%k���u��9��o"��r�f�˝����7�]Z��\�Ƴ��t�ܥ#��V�a,�.샶�|N�o�l�OL���y��ۦ�e�X�*(�ک��s��}��Gt�TS�܎�ͺ��~�
�w������"_��e�=\����|��
L_[�:�5�ö��ؠ���]-E\���q�C�3^�W��+si[r����<��`��������{��LlQo4�;���׆O.[�Ajy������R�Ռ����2^��7.�­P�FtcsO�o�GUWk�SD2��!��'��Xl.�LRsc�JĪL)��8�uW� ��������%��2���ʩݥ��]�V��js	�{bS���DJ����o�c�������¿�kxP�O�Tn�մ !�d��m��n�I�1����)= �4��az�[�7�k����Cf���;n��2�#�T�#�}�YWa�i�)�~&-�u��)��V����fpk%�������mN�fU�����4L+�߂j�k�=�R򟫨У~;I��J/LEe�OQo#���,ٺ���m�mB��0�xw�e������\����:v}*�K��_�a{|����7�"����T �wۼ�k˯.��+�,����F��O�x�N���{M����&��9�媗��*��|f(�������izռ��:�Q�4ҏ��o�wb�w:C{�[�q+��p�1�v���JY��{[բ(7�xx<wa2{N�oWņ��7W�WZ�Kݾ�{��<k��>�y����Ƨ=#[F�䶿[/�ә���9�Y����}���~��a(%�Ts	�M49XK��\E�k�Jv9n�7jh�4���������L3#+)0֮ҨO�Z�	�i�f�닏 ��s>0�;�`6Ŧ��ǜ����R�G}��[x�n�a����3n���w�E�L;z&e�N�� �,b������e�W��x5�>>P=��I��oO��z��Ⱦ���5��C�p����������][]��]��l�tM�������@�B,��̔�e��7cs ��Π�����P��j����{���od��ךE�ۦ�t�îyg�XXd������b�u�G�J�����Ǎ�	ۋŧ�2�d-|N�#�WB�Rq���,8Y�M�μ�ߐ����`�T.{o�e6��fZ�]ӏ���c��	��NԷ5?)�ɐ�U�B�ؔr��=;��4��)흚��i�Qb"�w^f�����������P��~�<���� �'IG0,�%B�6sxG�������}�^�w����{����}�߇���������>�O�����׿={r����������
�t:�x�3���:!�5�ᒏP�7[s�{3��Vs�+J�b���.��
�96�\Πv��
�gAYT�Ŷ�=0"���y{c�KŲ�q^�K7�����Wء��3�0�A�m��`5�t���n�C��Kh�o%�I���wg]�W}�oB�]��p��7]y����B�����K�К�>�XR���ʰ�j=��f	��]��+sz����,�j��(��
��7��*r[k���E`Y�����Wkif�6����`���Bo��a�c�������WSM�������|f�rL�]+�
`x�Χ��"��1E���eaL��d�o�G�-��w��β��q+Wt�8�w��.Xr×�Q/f�U�Q��X�`�� ���7��D���ٷ�M\7��� �G!x~�.\���sp���*��=�����.g������p�⭑��V�h��a������,i�|s�\j�U�iʔe�"6s�r5oi	�h������F�+�]p���hN�x�'����V��gT<6F�v2��7ָdV�pm����*����ߚ����˯`�Ei�8�*�U""v �	&�%%����i5��[���'Q��4γ���D�
���S[�f��X#*�Ig0�s�ôUf�]K1[��SY�D1�՗�rwů������a�{�ݿ��3J�TŸ�\��0Wnm�7u�����!l��Е�ܤ=.��=7�P
ժ�|p�����X7��{��|�;�C\�٢�tS}^C�e=���� P�6w�w+����I�C`J�Le�h�,��V�oT}w��un00� �L)r��b�(:'�ڹW��]�u�{��f�5�n�ʕw
j�\�r��J	y*��P
���
��b����?$�<�af��Y��M�N!6��%o1nT����Z������6��M:�mM��NZ��m�!԰e�M,��Y�c�"����0�l���9L�k7�[��6��c]M�T����V� F²uU��v���%�&�{G)�tTY��ʾ�n��1\�Y�	��#C	VӤeJ���6p䶢��_C��$멅hl��'KYW/k]�� ��wy�e3���P!�au��v���wP-;�\r�AV�6��H4����o)���Q���&�{��h�gP���[QG��Uժ�G�F8@�_eY�IqӈK����z�Tә�ܷ���f$`����>;X"��P$k;r��]�j�d&�lZ��.Z������:�yn����tt[&�a��4ne<G���c�I�Cj��[o�bfT�ł�l�n�1Y[���wKy���p=�g�T����ykoM§ZZ�m����,ǋ���-^��3��5y�s	E�b��ЂN�=x�-�
;���yn�9�Ⱦ|\̗�7#���!)$��_U�Uw������[��;��
�����
��AElg�C:4�5c:�b�ή�TIV��ޭ5t��
KF�j&"`6��a���$�"��M���6��61�&��h�֨�(

�"j-���Q���b
1�m�6mJ��:�.��5AZ�ES�f��-F��?Y;����X����Q��(�֖��h��MDU6�itU!QE�i�$�1%h����m�bb�MSW�]j�

X���"J�A���ڪ��t�Q��'�CI�QAE�:
SZ
~#GF*&���h�*��F�� ��&�Ɗ����1���LAAT2�PV�h��i*�� (���tĔU%QPiİ@hk��y���w���s��o{�$`~l��UF��%��%(��c�?4�+��¿bnmn�����<n�Vml#�W���pO�����/�Z�s�J��������oN|͇bv��ʺP� FPR_�����L���m�t\	Z��)�TaP Tl�[2OOO�{��_P��>��Lٻ����e!��+�Z�&��w_��0K�"����&	뱠��פ2����I�7E2�i��aC��{7���{��mV h
o��ե�2r��*����`�W�ekPv:��!I�=�O���ϳ���c�tz�b�-�L�w4�;��f����li���`&����p"��fVg���=ҋ��}�e�dZ~k	Ab�w����w�v�}���0un�V;��~�8U��/�B�s�{�!uI�8f��m%I�!dw:�WC��8������>�$!ö�*��!J٬��W���N�^^p�_hLK.��-llɭaD��t���uO��ܶ�ڇE�~3~<�<�X�ge�n���`�,BO"��O�ٶ�/��h�T��x�}�gӮK�lD��|�k3R�������u�2�
�uⓑ����~s���L�q�7�|�=���󺬮�:s�+�1�LP�7`f��PŰ]�vS��~�XD���}����f�D�cݎɺ7�ѷ�����\���݃��rhH�i��F4c�����-�����8�������P�`̤�Ԃ���.�ɵ�δ�2�ɴq�'}٫������ot��P�����l�f��A��aep@\���<�������+�kN흲��}��v㾽��t̸�s�h�*i�5L��J��k��f�jW�f�J8؈v�������<��s�3_�������;�i�(_I`J�h�%�<�ͧ��;6�<�ղ�Ŷ���߻�H���/FQ��Q�*�ӯ[�m:��l�2��6�5y#��gױ����*�;��0�h��|�|�K�)�hs����6�.�[�:��d��щOҌ�Trz�c�͏;�ޙ����9Q4?��xC�f��	f`��[ ��U�OЂpK�$���p�4��zf��f�-h	Y<�E5��1�I@���sǆks�r�+�LѮ�]����pd
��gq�|�O�%���{�-��g�z5�I��:���s���Y_|���?m�^_["��U��.���pa�B���2�k����

���Kn��#Ϣ���[�v2���XKL]n7UoN�6Ԧe"Ԗ���*]��!7K����e ���H�bX`=�6V���.$T�*V�]�H�����~�<�4�j�6��Vzi�j�㲋��5��%Λ�Z`��z}��t��^g.we1�;�`)��xv/ƦD��^�M�:z����'-~Zd���yyx��N̷�F|P�v��y�6�};�����J�%�:R�/�N�Ǝ�]���ʘ4�O�O��٠��-L;+�]ɹ�)���ē����}Gj>��;��;e1�Z&N�����I�-Y��]��/qdr�1s���э{�V� x=�s�����q����;H���2
���D���d꼳"�1%�v )|T�؝]�����{���I�G�����A��qO�i�;ka|�d�-�W2���5�K��G��3؄n�86��H�v�1\���-@��q]4�^�����8�V2s���}��~�GW��&F��A���hE4]�2�Z}����,�{�m��wZYe��v�SoUG,ޚ����жC�F��&0�_��m�{�_� fY���<�EM�\��H�ִ�k�ک��nK����ٶ�<bL��u�d!�<�lKت��v�z��ڡ Ⅸ�Ũ�Pc���my�M�7w{{�+�n�3�;?��1er��I1c�0?�]��"�䃷9mZ����)L6uŭݝ��������D��z1���/P�3`A@��`��v�ɨ�t�5l�eY��qZ��:�q�%�X�hR�J����8����A˸u��!7�{�ȼ���-T���WW�����vC�!!d��nr�?1)�FE#*�i8���oE������z֯�1zV��V�W��B�H�>�5�Ǝ+�XMA����\#0��i�u��`s������ڔ/]z�r9�.^�B�Iuה�C��6\������%��p�Q�ի���y��V_V]cp�zo�Zs7�Bj�=Oj=�u��]����z����g��c��7���C�b~ۗn���&S�qK�� �7�3����+�	U�!x}�g��j�x`���0!��� �y�d	e^�5ݎ&J{�f�s�o�9���Q���^�r���#ks�mvoS��Ց:J1�&��vd박�M�L�l�w�i0�%s�In���f�&��'u�gN�����{�}��p���,�?э���t����З�u]J�,�z����g���;��k���S�C7����<ʕN���]�����=@����!-\Xc�L_+״+v!��<i΍��ٛz�7+YBͺ��:���{�PK�X
��I�a����%�Ø!İ��p����n�[�}�ٕ����|�L3,�7(�֮Ҩ?Mlz/��5mR��z-A����5p4���W�Ϝ�$j�E�x&�6�ba��U��f��nQa@]���h~�B㩺����6O��g��_Lo�u7�R���u˝D,O~!9[)ٹ�Gz]�xfE���HzR�:V��ftrz��؟p�b^-����@��eϚ�vU����{kv1��7������2��VA�yY�!�f�x������摢�j���\��~�����U��>��J��n���.�_G��Ü$r{!%+�̬�y��eJڏK�ǥeL���p:���dՍ]�W�y���[qnVX\�܇�[d��+M_��U_k~V�x"�U~^j	�z9��rE[=]�������( � ��B��H��t�P�:)�0Aaa��@{���=t͝
�=�;��w]�M��n�*���T��c ��H��Q�Co�H�.:?���J����*���^�fI+��{ٳ]��	e!<�LcwX��nj~"Se�!2�F�'�(���׬z���W�
z4#"���ۘ����̙&oO��ʘD��� v)��%1�1)��),:Jg�K�I�\f��P�i޺�|�%�w?nO���T��x{�GT�p/>�#o��7s�D����\�M����>�s�v����V؅��¼�JET?���k3��]㠔۶Ο�n|�ta.��lڞ�M�w������f�s�ؖ4s�Q�NZ��mxw�� ��Dp��B`&��]��]D�f���{�^5Н@�s��X����Z~k	Ab�?7x'���!�{�ɵ��<������r=Z�3�Ѡ�1p����O�1����k<ل��zYΪº�Ado�6A{�!�p���߁�Xp0A)"?�b��
w���p럨LKgl�je�ΰ�J�װR��)�C67����K��_[>|�r��}�ۖ�7(Г��)�����d6\S�\�{d˱z�wM�ycej]j�\�6:�mgTD���Ag�_d9�8�&���Ŷn�z�����:�3���Q��y�VH�lg�<�2����rʸ'N�.	��u�Z�}�xz��'��55�X<�C\?��I���L;6�ϲ�m���Ll'�8������0���^Z��e`�wD[����c΅d�67����O@f��<�D"��a~>7Vd&l���w��S�gZ����s��.��t:��^}�D[�u�v<��A,#C�q D�������J��Z�ѝ�4�h0�:��`��8�'��i/��ӱ3����҆Al��$k]�3��:�Y�܋^���Z{��1�,�4/��5⮂�����OÞmᵡ����1x"n�f���A�@���O�1�O�r-�JT͘a$Z��j�G(={6q<�>�A3�����rh��ْ�n�&9t)�*g�v��=�+��rkX%s�^<�&�@���.�%B�~�+�.��f{$m��
� ����6�Ϊ��|?!��s͏߂���"�sS� �(�-��s(�w��V��.c΀⦙\�I��;��<�z2h!D�f�t��cH!kݜ��Ϛ�쫭z�;q<��uΓ�u�.�,�%I����<��ȸu���<�i�Y��>�������O]�^NɵzX���iA�θTX��;]�֛ދ6���8#�Q�lmln^!��gT������+f<\t��$ɖz.-�`ŷ� �q�bܚM�W]ج�ϝ�0A�]/d�Υ�|�̼X�m��M�֥t�4�+��ꡞ���{�׷��R���'��$��9��o�ȥC۴XsQ1��ϸ-���\�jPzĎ�Ⱦ�680^O�m	��a4��*]���/A�����^�|UF%�ͼ�����1#9�W�՝�����s?�傂��s���<���Mݪu���/+ kt�s�菶�ǈ���l�n����Q�����
"���=��?.�@H&����p�*���g�g�B'߰��8�'w+��zC�}UH�طvm�l0n�n.��蹗m|��hZ�+x<�y�2o�[X�����-a4ϭ���t���8�b�a��Y��z7,�1gmk.n�vB�1�ԉ������e�h��s4�����@�r����s�<h�ge=��	�&���|��3F"�D��媑����9��>,"��.��#Y�T1j`��DYz�oy$��bء8om��'s�8�w���
5�&:�uN6ۜ�@̳B+�Iv�T� ��˷v�����`4���'�7=ĭ��s�����U$�����j�p�
ޜ�l�U\��mV4₃��1`;���5�}��s����=��fD�f�E��)��i"�`�8b9{i��-.�C�ks��O"�X�Ae�����̡Vt��:���qO���g�)n�#.>��&^���ͱ}�|kH:y���jDAh˹(os�\�Q{���Vm}��DG���&c�5�ށ^L+�(�{Ù�uzH�	;�c�?��� �ǚm�]{k�me<GHh��Q��� �K�]Z�,�˽6����k�\��s��?�w7�o#7ג��lR�'��z6��0TŐ���������'W�ХbU&���8|��C��!��%@��S����;���nRK��v!{�KsW��2��1)դhZ�)8���a��ЊW�#�<���ûZwW7�##ZD9!Ĉ~v�ۃf�L4�w�Zi�b�t�Z{#��m]�\n^q���h��Υ��߭ᄍ�B�3cH�!?W��#�{ K.�0�eIOV	�d]E҂�'Ҟ�K�3_���ή��kWc�)���~e�0���aZ�Cw=z^S�ul�[��&�0ʵ����;����Y���ե%�+��칀YaE��ϛ�i�so��0U]w�"n�l���ZǷ���P؞�aE�,��U~WZ�|^�����>�`�6�g�>�7R�,�{&���Q�U����HY�-Xs'\qn���A =���z��^�%�s_�����>������ꊌ�i01���ǧ�c B`�Vm��m�5�W��7�w5Fu��Ӳ�cP�φI�chr@��U��]����;��2�/�U!wA]5^��`�%�Na��PwP�H��xxj�.�Sy9C��k�㊺��6x�rPZ;:<�諭�h�+�5�Mzw�l�rﶣ͏_dS���RV)�(01b������P���0�ٹ)��bR9�5�`�f��R���\�԰�Uĕ��m�s6�15ژ��P�+t?��'�w�5�n�\7^]�=۔X�_}����#R��b&����=���g�rӲ�E�P�#<O�@:���*��O�C�Ų���n��S���^C�5{]tr)wg?��$:�CHD˴��-����5����j��iq1�(��E��E��ږ��ᨛ���i�̵G��\��
�W#^i�m�P鋇U�g�`���$�i��%����{�'����fpD_Y���XZ���:�WB�KԵÞ3�^j���T:)�9Z�J�yȷ7��[���SS/0Za�[�|n]�;R����%6}!3�F�'�G(]���׺f��0�*�κ�v�����`1m!8��@L����=�y���Ǽ�%:���	��=S�c��3�V�W�hC���ǡϸ���=��qm��0O v4;��!'o�p���ǯ/{'c�1���)�$�K�����i���M��*�D��,����`�/?}����؛A�Z�?�/�p����������G�"�XR��s�|n4H�K;qfZ���l�U��ܥ3I{jxyC�d���+j$�vݧ�nu��(�1����J*=����$���ʴi��ic����q�dCb�����j�zOGD���1\�S�A�*��A�n��� �A-ˆkj}O͸ܛĳ��X�����v�n^��)^*N�U����j�7��9�i�@>�7�O�a��Vp~�����Q�^w��]o����CULW���vJ�/Adw:�
�w= � s����|ygx��²{�X������οP���[TZ�XMk
'�s���NU�3T�:&���W���}}2����5�ÐY�}�"u|m�v���l��Rc~OO���rakr����s�Ӯ�tkO�\�1a���3_�:/_9_���˷L�	�Eշ���sM���f�s1c��3���Ǥ��j/>â-�P��g�]�bµ3��"�l��Zd���G�S�,�3�m?n�s&�;}���q` <M;I}����2%�<��/xY��fjYx;�U�E���:�E����C[u�36)f�����\��A����>�Ұvr۪�K˩��«Uu�~��֟FFS���s��[O��LنcJ)�e�Pw����������o������}��O�����~o�۟o�|������?��wz���X��d�F�uE�O�l�����.
mu�9w-4�J_-[�G�]�T�𻓪u�>��5��o6�Z^�A\)0G,���4QotS�\�r۵�qT�&��yF�>$��c0�W[�3!��
y�;,��8��:.�ľ�9b������}�}���ӡo����ճo9���z�ָ�]�ugJg_�k9���%��j�*	�&�K�B��ȄL�r�����5��-Ėr�Ռk3s�sN�f�]���l��!��hIc�0nWr�����b�ld<�R<"�6X=��A�%��vA���a��y��� Wr����X�}�ga7y�gw�[յ�\�%i;��Ŭ+�� qWwX�U8]H��'0.�s0i��,�u��Zn�2�gU+K�od(���Ul��)"��k6t�1A�~�ǉӌ��V�iw�����nd�3RkD�^��}iu��M��צi�2o3g��|G56-��ȣ�8��2��Y�l���+q�.�S���:�l�oa��X�+q|��J���j�gJך��s��%wxk-�t��nE�+��R�!#�Z�v�}W'�ԑ��/^�Vd�1BB�m^:x:��Ss��Ȓ��𹩰 ��LI�����}M�G<T}(�\l�-�uso�4Fm ��np���]�.�﷖m��k�z�a��/��#�|��]�Z�ҟ�t��gh��+(^�� �;����m�x�E����h����~��3�߻�r����̉:Y=�,1Kp�XAQ5T9��7��ֹ��]���"��籔ɒ�7R��'N�Jj�)��o�-h�ػ��I:�h���]�,Q�]_9e�lL�P��*�;=t;S���H�n�����M��摜��#�Of�����be�����J�UǱ8�:�lj���V�ѽ2���w/�s���r�$��!�to椯U���S�i1f.�3�y#8ekJ�9�t�m����[k'��У�z�ا �q�T��� �h���3��h%X�e�*��>��\���x-��.� ���M|�܂���xL#Ѐ��[�.zk�Yc�fP�z9�ֱ�rQɨ8P��/�ꎙb���|�/��gFi����"Gsu��_��f��k��o�*��dc�\�LY���N��Af�j]�'B�.��mEʸÓ`F�՝�����H;�g��zr�Q���v�mB�����WL,��X��oQ��:��^9���Z�^�[.��+���n��q�uڦ*�N��S�����+���V"�_�&\�\x��nt��ǔ�xL�J��b�5�js��"��Y��Rnd�[N���4��Wn�V�ӂ.�Y�WnX&����)t),E^=Ç)��t��� ��\�����$��4��޽�w���b��������m�� ��KEKQ!M%�@���i:u1I$PDz؈
"��-tU`�ݭU��x�'MD�uESD4EUz�֐����b��訊:��z�ڒjj"��

��)��"������2Dt�X�բ�[�3ф����[Z�$�����UQIitDP�'F��Q���ZZh�U-أcU�i�P�[>cvT|C�����.��Y�T����F�A��Y�t.���5���ޣ�ש:61E��!��4[Z΃b�Z4Q��*���:�'A�h:����F�%i4[k^w��۸��׫׬QS7Y)��j��(
�ֺ��>'�����Ӝ�{���>�;���eL~z/cO["�b,�'$�����2�#��]nq+�Mht��p�-R�u���m	�D8]������8L��aJ��OV��"���h�����J�`���z}�D�����j�w����B�Zy���k�N�+�`��f=���\-�=1�	�D]6?~
�`"�s��D45��&h=ںk��p��X��H�2�%*Mv!zN����|y��xA��Ivl�0�!Sy3�G���W�D�Dk Etqt���<�%:]YrJ�[X��Y�����9ͱ�����u�ܒ�JaR�]���&H�I>9�NP��O0��cϟ#Ϣ3)�g,��-����т=r#YT���jOc
�i��&t��O�)�+��[~)IZ̺2U���s�v��G׭������<����G�]&%�:�����Ad�����;i��	���K����Z���5uzj�c�@#l27HN7�t�u��>�gcf���K�M�[�����.��͏�6�ﺣ�L:�נf�X��5���l;���\�tv���z�Q1y9}�\�{�x�2<����o0��U�!�����	��v����ŀ�?��h��K=�U���h}��vtz�A�9�H�1в�^*!�v�x۫���i�������M>>��dJ�66y��uhUǎ��FJǕ�MLuȫ	)���gV�1�v��Q�v�6��a֖n�+y��	��M�x�)��r�m�i�x���{�;꣭=�v;�ׯ�d�D��e�'���S��bXo��Iy��\�~b������!J�W�EgLa��z���-gd�Ƒ^ԍnV;�7<��hE M���_v-'`��^-��6o��9-SK�w�/ V^
�ȗxCB	��)��N6ۜ�G�,����d�j*m�e�x����ܬ��t��nݧeO�i�ݞ�Ǔb�S�
ϐ�a{�d^�Us����8� ��3\�J�ʪ�ǹ�Z���t3gW����zw�X02@�	<�|Ǧ&nA9�.�����]�M7��j��^(A=��BF���v>5eEÚ��fpP.|�"K�T�xM*݆V�s3����콆S&|}��ĠώI�Rx#�JĪ0��.�ƯuEê��q������X��uXT��1^mB�s�l;h����2N��:K�QR�'b:q�T�\���C�&uWt9�2U�R��>b��}�F_��xu�x�љ��T�`c1Vt�OV��݁���}�=}����ޢn�#-�?������YW�COeIN{|�5q{B�pڧ�ߺ�m���!PWX��������9`����=�@��SN��w��Ν9|٠e#���'e ��OP�n1x�n�	FBe݌h��}�`���/�:d�{x�z2�m�rt��{�.��gg0���Y�q�4v��G�=�7�s�ܦŦ](�!� 0u�t��� sO����zk��z�Ϝ+.�b���U�Ǡ��[���i�^�ۆ26��w��鞎E������\����+��	��G�!��0�6�Fy�?:�j�Z��㘉=�{��ӕ���XⴕE�,�uj�Xa{mnip������fC%3}SyU�[xuhX�y��m�����,`�	�[ތJ|kʎa'�N����߄6�n���ݬ��>��j	�TZ�!ٺ�e�0-C�*7D��3�a����9j4���;�����S�QI��LܸE�O̘.�q���d3d�����bK����p[o>�o^���;M�{�{S�z~�T����ϡ�=����dpoS��ќ:���1�ss�q�u�����CO.�C�X׊xn�dg@��B,�{t����ߣn,�}�"�-��Z�[1���K�*�!^�k�7n���:��#��&r<�kBO]�&�o��p��k^�WzEu�Զ7.��� ��H�~�~Ş.�{0�.:k���y{z���c/���f��*���k�M�eN�x�%۾4͑�ٛ�o�v)"�c�]7BzϲOd�w�{j���n���I���\��j>�|��)�f��1v�ϳ�t�m��
u�sV��]']0o��G٩�ʳ�gG��P��=:s����@-kL8�|/��d�F��ɀ�η�xش��մ'T�@�~�
A������ٛ3w{=TKD��S�;�m~N%�b"}�{��A�F��P~B@MDħG���`�����;6��Vo�u�������K	���l�!�O#�y�!GUx��D[Lo74A�Ҹ�=�+����E�tS$���|��y���^��7���W��~��mEQ&h{)޲�j=q�t;&6b���J.�7E2����9�gp���-�	�`��Q�v<�t�vs�i����L�fxХ�M'p�������֔+�C�rq-��6��;B[��l���kneAi�����j�����J�/A[�twB�7�ֵ̗��Q�F�>���_V�_.p�n���(�yÛ~��lT6�S*�OV0�P��~�w��-L	��O���N�Z
n��u������� ���!�]4ód\8�^5�:U���h�2�.�I���e�{zO�W=�K��L�@�Ok������9�2~X||��Vx��!��K�p���ι��٭N�NS�J%җnp��5KF��KHsJ�`o��2�FZ3�,fD0����Y"Ow�C5#-8���M7Ћ�&����{���(�쎻�������k`vrQ��kk1t��'v����&�жI  V�W���ɾ'�T돃���O:��ǥ��@��H�m���Y����0:.�=�Onr��ͫ1ݜ�]eBdlwA�A��n��1o�סo�#B񊏰!ͫxcOX*)��.*B���٬�A
e���2��uE���wW�2�4��UHѦ9�!{��x��yvF�͵�ᗩ�<Ɩ���Ysb�}<�7"�F����fbTSئo�y��չ���ՙ]��ɪ��b��e1���R5,�����=2)�	X����x�MY/���M�V&{n�u�G"O��+��S�)tf=[է�h�>1pXp�������}N�cX���ѫn+�['Q����Y'HĲ2�
�(�|j�t���bA�	��;\Z�E����V���ޭVÖ&���,��^~��;�뼔�e^IRkk�����i��-��2ޞs���/���D!��a�t��nOC��I>y���a�E.��N-0-iF�gj���qS��*���C΁�j�H��y�~n���������M�d��1i�c)�������2�
��s[��v4Th.7)�#�O|=�$N��U$s�GY�w�<�}�z.mK�2���ա9�%�V�QZ\^���1��t�l�pA��hb��ԣ�n�Kzc��b��d����=��a��gp�^�� A��Ȗ�Z��[��έ�+|Zo��D)������D�~y���xG�����Y5y����P9(��fkƛ�6���&�n�Yu�r�]Q��㸂���ql��a��y�MƦD뮘�g2rI�)�0�OT��m�ٳ��,���a\�Ժ�����d��1��#4��x�~����h˩��=�I����Z�S�a�➟�_��=_�Ӝ������+B��7������Yߑ^}u�X�ێ��fO��hm�)���4����b��L���M����F4�f
I�o'o�3���pp��~a���Xʃ���Poj��9��G����*������N��w;�����y�Ӷ��+�#����������ʣX��S��Ƿv>��B{Kv	v�l�~���7�o]�ήB�!5�H��+7�yLO�(`�$����a[���W>��l���3wwI��k�XoL�r�tŨ%r�W�FC^�2΁l�G�H=/:uH�!ʢYz�C�:6�����pv�y�H�O���n`&U���g�v8�\�C���P-�}�0���y��0���yGbꄢ�7�QuTRԝB:�u(孓]ܶQE��8�H���#���`k���f=R^�s�r�us�{���A�F�F�b�O�#�ֺq��0�>��D�q�,�vھO.����\��_iŏ/WV�����L�Ș?��kſK�ҵ�5�ɼ�a���tr��],��ٕ�P��Ҷu��2=?A��tʗH��Qjv����m�0�3N�^-{�n���"΁[��ؘ�v��"�öKSh~��<a��t}��U
Rqu�Q�qa��]y����0"�[A���H{hNPq0�2�m˷�Α wJ���L���
j2;)�6�3<��g�6���C���F4���L9�ݐ%��P�F�[��cѱ.�}�mͰ`���#m������O��Ґ&��K?!u���ݣ�6�_����~��&y�=�E�N�5�|�al�<��):NX�*���4�#q�D�_Ƹ���g0���J�Q�s_z�S�{�4 vN��T��gO2��>����ON1�1Yg'�;���ݽ�ACs�l#�st8�~�n�̝q^'�k�J	{e/�^�G.���L�8_�w�~I��.�j	�`��<���� >�̯.y�m�J������`N�ڍ{Vf�!�4�f�Q�]ًX������b���fq��x�	���ss�<�o��kӊ�x?�ь-Vt�a���P���Sg�]X��3�O�E6��8�j�נ�uF+�ȻR��pp�7En�K=v��T��{.��{���Bt�T-vk��#Ve;�ZI���F��೻�K�W�����;_GI�*Fk#Jtr����iƯM]�_�V$}�ދ\�=�S.��M��苯9�tg/<���ȇ��Դ��Q;��<$�wu�YY�|�7���cY�t���9@!�?�'��u�-�)�dg�`L�\5i�Ɔ5�yM#[�}���-�B�-=�׶�fG��/��\���.�1��t��>זq�GMFƜ���]�w4�E�A�8���ǿUV��Si0:�2�R�'=��&E���9U�N���H�(�x��aAi�9�c%0ø�Mh�	�F�'�nI�;YOם�3Ll�mՠ�c1�z����v���i ���pH�U��G6��%4�i,����f[�9U{{�;���8c����S��)P���ǭ�;1�)(!2��;ȹ�]�-�u�Sc/i�6'��rom�V�w/Q���2�d��]ʼ�����g��T��K��a������d3>2|:(�J��㷛Z�7Yhx�y�tQt��]yb��F9j��;�4\����s��v�Y����3���y��F��wt����҂�t(~n	İ���`Ȧ�ÖD���.���92�m5e��G\�۔1����M���~���~�E͜t@�)�Y8�(a�T�vΦ�����p��a��V6�U��q��qҘ3�n69�58�6��o:��J��:ḱ�qqn=��5}Nj�N��1T�z_a͇"v���yF���y�Y?���73����ηj�\Û�l��Q�X��y*�r��e=�E��i~���"YJ�[�*�}�^� ���#�>�6�S*���r��y=�{��(	��qlӻ�ˋ�:p U,�Cb�>�Ü�]ٱ�(vl���P�z6X����̷��9��҆<�}��ӯC�sI�i���;�Ǝ���^}��Ɋ�.Q*b�\Qέ�{����R�B�)��^=- w/4ߘ�%�>��ź��Xׇx!��nkI�Ʈ���ך�����J����t��;X��Gt�8;�Ӵ���H؊��щ�B�}��:.�j�i_u��t!�XQ��[�GS�=��/�9i�+�KE]9Aw
��O+�ٕk��k�e��i�E���#Yۗ��=q��9�r.|�5%L��0�	r*(K�$3�I��_�ѿ���a�L)��u�AG3����E��q�
m�1�>�VcFK�"CGwwGWX8�x�A�P��#��ݿoV�^��3��]��q �p/���r]��m
�|	ӯn�����i��h�g�晔�'}-pR�������L����B�H�c�f�<�Q
�Y����٠�0v��p�t��;w�OI>r�D�P��;��'c�������uh�Xe�[�BsF�(���GWt��،�����g�2!�0@�!MNapK�$�3L�JW����s�:zkw�H��S�Ts�­�5�5m�6Ö�@#n;]�L�ۘ��iH�T����\)������.q�O�yz�W��w�{��-ƲL�O�c��i�*�'��$��:���kdu0؁39=Z�t��Y�t���G�Ȅ�Sd^Ȓ�/��>�,��1i�Uc�; ��ZB�q�W�z�]��hk/Qǐ�D����|�-�kL9���i���}
=d��4���sT�w��=�9�^#5ֶA�ϺsX+���oL2�b�dv�����3�C�W�14KsЦ#�V���i�9���V5�2�����W<����v�,b �H��{y�}���Y59OU��uW^���]K�G:E-1%�}e����g=Z��a�����w�5�_>��d�`DUff�]�C��"Z�=4�t�=xK�>N⡴;e'���
$@:I�Qn��c�q9D^�*}�]��~���@���i�u��8�m��	���A���B��.��]���K��>?/����Ϸ����}������}��~�?w����z{��Nv��cA���n���gWs��A�t���e�����B�����0;�}K�,rl�ĨJ�u��~)�T�K��/i�Pc��C�1��xf�����ָ�V0���2p�Zp]�Y����QX�$�	�CBi��mʛ�NK�7�ʓ��C(V��N�iv�]ȟ[��+Pi��j�=5@hg^OZp�J�� 4�Y��*L�ql�W-9.�Z[ws��.e�4�����g(���R�o5�k2dyz�K�\Rz���u5���3n�Y0��cvÂ��:�{�Sא�&�[ɷacڜ��XzI\��F��nV갖4UVh�����EBvwA�2B��6v曬x�gI]�Dv
�˻�����e�+�;8��Q_#aɐ�c6s��p�z�\����e[<J����zE��grczZf�N�,K�HA���e[�/b�wz���YZ� r�٦I$l�/���8�{��ޮñ6r_;6���cs�A���m���er:�HTUlf`!�;ӕoWY�jK�.�f��,g3��26�V��%=�*ΛN�:j+�LN���y�	X��:�]���u�Nw]dZ9�v����;�9�?$U����%̘�1n ���R$�v��]Ț�f�a���w�z�F��#����o�;2�1܊��{�sٵ��ڽٴ�<c28H��W"�@���*U�2� �$^:-��V�K�$�\��~I9õ=2��9A�#e;�������oެeE�I�/�(�}�)ڢ����8���9�B��$iu��Jg�e�M�]�W@����K�1��ؚ괒� 
�vx-�+�Vi����j&�`ɰ;{[�^sp<����cf$j>]A�,!]`u�B��cN��n����y��׷n�V���Q��4���S�8���AYCY�����(�ϟv�ލOK�C���~^5\�����erm1˟(�7��E��WNղq�ٻ�u�l�E}W���7(�ݴ�Rz���f��.`7�
>V.�CUѾ���EYBV�d^�rj��n��]EΎ�X��v\W�Q.�W�9T
��{��h�����c�OЍL e��5|N<��٤,���T�*�Ȥ�<Ź�N;l�9��	��g�X��k���N���� W3��m���o����ڻξ8��ᑳwtFS��Y<�ubYz<�*݊�6�y,m
�7U�Y��ܮ��ٕ����#}Y���\�gLN�En�w2���vꗃ������V�F�'v�EQLfĩI�?<ŵbs�L@�Q�M���|a=|f\ݼ�8�>�%>t� �:�Z�/�k��P�vt��<*ҋ��%As�T���YT1W�ٳ�t.134�4�u��4���n�w_"���Y����6����1���r�eWd��>&�ko6���y�j���-���%A.�u -H�|�qi9 <�U����մ����U�Z�ꈫA�m��=N�JH�6��G-5A�h֣m͉��S-���kܼE���4R��fh6��n�z��K��1���jZ�k���F�*��������b� �(>6�(4�*�(
J+l_[1���1�$�RЕDAI]:�c�t�kUU5��z��$��g����;h�����o���#�i`�(՗N���T�
(���4��h����m6���Ɲkz� ��U^��7X��5Az���U=�C3��KִoVi�4j�
��q�i���/^�Ԏ�^�-WGh6��l��t[we���%1�����~%4���4�k�:���
[6GZ�����Q%}�����HS��b0���Lq'M8�,�.�BF��q��kF�ٷz0�e����D!��ͭ�:`��+5�=+���|�ٛ�ә 3�ዯ��iݮ�|���XF�p;M�Il/[F�0]$|C�#FJS�y	<L$�B�aR�
yRp���UJ_�V�������'Z�P�W�X,݌�*�%��sC��;�^�e}�4��C@�q�10��=W����2�5:֧�[95�s�9�}�v^/�i�m���π��B-�y�Ų/`U\���6OnQ@w7ok��M8��(�U�!�QW(5y#!�׳l��[:y�������p�y����H�
5��ʐz�"����PS�Xa�L	eI�r�n3�1P憴j���Ż3A��=ܫsy�J�DIp���-��FB��!�=��L��J����x���M��P<�_S�
����Xrޠ�H�	;n@��	��]2�^s�XH�]T�q��[
���&v:�Uˎ|�a���WN7�5�d���!���v��7:D��T�R��L�%8�ۘ�������n�:�M
��_=;ݼ0��"1�'� �y�d	e�Ypѐ֓��Sl^����ܩ��O'��S"��&���l��J'I@�B%�rX6��7Zn{{����7s�����;"J[I�Q��!��]Gq]���oC��p���,��o?���cm%U����y/x��^R�j�a��d�DYgm'6�^��+��Uk��Geeoq�M��l���g#�Lpꗱ���Mчl�"P��y'�t`ʽ}Ӆ�j9K�M]�?�+�g{%�v��,�ikvn�-����3���� ��:��;��f�]�a��Z�7c����]J��vN��R�&ΞeJ�Xo�m�>���Ӄ���TM����=����Ԙ:a 81����pȥ������I��c��֪9�od4�Sw`yZ���~����~�id�2��x�>$W��am��2���kݩH'��k^��e��ǧ�4�Oq�f#���O,5-�CǠa�E�� �%p��`h�o-u���嘽�U����e�_�~���6�1�0�uɈ�qL�χ<���"w���qL�W� ��������D]��Ƈ��,ȶyݑ��(7�tE��x�������;}����z�Ǭ�������:��/�u�2
W�K�y�`�U�}��t�����U4��*Fz�K: ��닋����ۓM�J��� ��HZ��)sgr���j�ؖ�����g��UE��]�@��O��s�|d�&w����d�L���Cz���)���k�i���:�n���}Ol��L!��	᪼COb�`��Թ"!��m�Xn��6��F4�ou�ܥ��i��17�_Q�SK+M�k��v�<��+tʴ�����������+����f��{�%���_�^�ݬ�%u�R�Tƫ��zx����zk[e
�+N�`d�}�e��c�KD���<"�~y�3I=5�?c~�%��S�\�wB�|��X��xB���"�C��@)�C��+� ��0��]#Y^G�2��1,��ye�IR�8��PYq��܂c�6|��p~���wb��S�XU<1PX�d~��F�X��i��r��k��@�. �;��}��{E�0�"5�8�ݾ�*�S�^8�z�|LZ~k	AcK�C�4�ފ�IMU��g�fh�*���<���cH������smŒ(��F^���S�!uK�˱�����\��r�&���9e�����ں�p���~��Ⱥ<�='�N:|V��oN���N���{
�x�~u	�>TC�` �~����4u�y��]�q؂/[zB�Z�㯦�v3ݭnFMA<j}&=侷mC1���z*��q�}G����S� �M)�B{<�;p�dw0gh��-��]�̅���
~�������x��H:"ۚ�X�hׇx�ǡ.L닊��5iPZÃU�^�Si�mF�+���cn�$>��@2N���h{|���m�~�l`4v�f�Qks\��s�Ac>�6���F��Z� m�Ä�H������)�J�t��eL�*�2}�^�aw� ρ{0�~[K
�tw|����:��zV �P�d�Rؑ��EsQBsբ��j�c�3!�{8�nъZ��	�%<����a��g���P�M>�9i�Q}q��s����w3E��KD���/с4�r��R���e��WP7}6�ĭ�(��!�,Bib��-9�U>�z܋i��mӷ���ϕ5�/3���wk�"��0�C��\�o"��e1ж��>E�(M�X�_"��0��i��:Л� �Gc���SNj��.[-)A�W�_���	�7�쟕C���˝U!�TV6ǰ�3�Q�w��՞l!���sS�����7q]މn��<m����]����S�s�7z���ٵL&;�#�d.}Й'�9�N�)�%)��;$>�dCn��=x͏SEA�͜a*���
��2�>���n��nOC���"�xr�,�Xn�J)D\���֢��ѵټ�����=�y_��'���4/W���:���A~�b�i�dR��͓i?.�>fG��V�i������sO�����X`��,"�@(֘r9��z%��S� 5c~��V���|-��I���s�
]p��	���I\X'���oL2�[��Giso��������x�bt�ח��ٳ3.�����$/Y"�MT����-���ͱ'q�Y'}��5�e�Ġ�c%Ѕʾ���)ņ�u���m�zI�"��+�]_,�'����nk�Ռ�[��:;}��e�&�vn�=�«�n���ZZ�_\��'p3��_�gR���M������fμ���f�P��v�;��Ȼ����}X�~=%8Y��諟��N��{f�=0�2�H}؊��� �곚{4,�P�u�KǓ�nK�0��W���}| ���w=�>��N�˙}�$�~����gv�`�ង&M"���'���;���픜O�L(� �b����d�n�=�3��Rku�>��~a�ם9���T��_u瓸h�]�8lz�z�V�v���P&�������t�:Ac�)��V6W���~���E�a��ƫ05,�O�وF�w;OC�65֊x�̰>B-�[�"�����R��u&�����WV8����t�*�b��Pj�FC^�2�⚽����Vચ .�ݷ�:�5�?s�
���'"��j��[���Z�,�#X�@�c���s6�����ӧ;�A�à��&5�p�2n��_��02�%�"-g��P��m:�[R��y�Y�k3:h�T�C�Ol�>��(R.��y(jrG	���s�Eؼ'-�����>�)���<��&�Rmފ��t�Y�F�^R�֋�I���$�3*� 0�Yیt�?a#X^�^v<�����N�tg	{5L�l;`�E���{=x���1"!�Rw=����.��k�V�N�| ƺ��{nm�.�|	���veM��7a��'�,�f��>g�}�a��m��!�����C-�v��}OQ�ظn~|8��k赍�\�6��/$M
��_=;ݼ0��|k덟����5k�s���L_��v�΍��r�Ҹ�jR������p��+}>@����y3r[ֻ�_lMi��n�h��t�ɮ�U@��n�K��:]J�}��P%=]z����C
��rptǈ��ڡڹR��4���G+2!�P���uᾬ���0�=�0�8aǤGb��@���x��'�Rۘ�T�j[:��M���V�a�P0�1�H��<@އ�*���@��{w:s������w\0ή���^��XH�H��`F<���	�7J�m��g��4�㝸���$�LG`��Ns��c0,,�U-��<�0�����W�ݝi�K���7O�1�۝Ñ#G����/�/�?��������r��K8|EPҲ�8�(��w�$�m��+B�V�'\��1���V��uVC�es~�q�N
��V4�h����v<��k��,a��ڒ��VsVۉ�xz���E���;R��d.��t����|�N�_s;(=G:<�=ƴ�޺�/M�aՂ���wb=7_m^��C��TD��M��?*Ӹ�vз΋��'�P��^P�0fG�F}1wF!�i��]��>�J2/fS�m������2�v�����ľ��!S��~��X���
r%0�E�q3�LWuޞ���cڳ���.A۹-�c"��6�+��V|u����E�]ծ��v��m�<�E�&�ԫВ�ګi�M3�;�n��V-Zv:���.&�;fi���>��G��^�j(c	R�2	%S�{:�-��ݣ͑I�)�r2��l��u�h�\Q����nk+颞�{�z{��4����6g!���h�y۽����܃s�Ad7$F��t-��<mlH�u$O(֣�-�qOU��8���z��B���U����=�]�h�aE�|��Y���k�`��6���p��0އz}�bz=>=���ֈ���F�z��\̂8YՃuv��el��ͮ��$�#���`ƥF"��Xq��=v�l�۱��q�V�i����Qí��j���P3��}�� �d3ic�݇w�wmT�n����m��$-�34J��m�}���V2e�f�2��7yT��������������e'��c�8�/���c9e.��Ο�b��"�I�X�q��7S���f���z�*}��\�惖�����μ��՘���K���7-6nr���l������]a�ڪ��ǅn��ގ���Ǆ�Y�����]9�H�Oìހ�}�<Xƞin�V�&�٪�wOTN�P��QQ�;g��BꟊU�yF�n��D^����#�����Uy��Bwns],��`g,��R1�b�.�����-� ��̝��,k��GtzœI$m�m��V6Y�C+��Bgu�y�M�A�����P�xA�!Q()��=j���4� ��v�z���aVQ쎣ѣ�HBZe�춠Ux�J�2�B3>;`^�ud�LCC���4���;��ˇ8}[�:;�8�CjF�t@�J�I7�<�^\�,O����~}�/�0��D�T�ۆR9�<��ǰ��.�_-�97w&P�;��+2��ض��vCw�@{R__r��Y(JX�Xd��ܗ��g3���6�;��B���1/���eΌ�}�m�ۂ�cN&0N������vM}�;�)�:;ZQ����	ǀ���3-ˍ?w� �H@~
Sj����RVܸ��i���sV{�Q����+�$l�f<��.�e���[W���)j��nf�D�"/x��DM^��y(�%�s�l,�n��-�9�"�<�B��MU�9]��o[�M���rU~��һ��kC7X.�96�����& ������o��}�R/�=�/+�3F�����=3��v,���g(�����p�y��,Ү�/�_V��4ch�v��'�ۄY����3[��Ϩg�����@�9ؗ�d��>훩FMn杕�ݙ�Z���e��sN���G�q�6�w\�܎��j�^wnF�p=��B%������1�:U�V�B/���M3-"n2j�M8�ż�"@(�O4[j� �:*��(�ޏ?�&��d�S9'0w�0=#��c��m�����k��s�)�zW�[��T��/��[Z%$�j�
��6޽��34�儣Ζo��V:��ג�]�Qv��lXW_g]��gD]�f���"��|e�T���CV�:Ռé:H��T�<�G��1�s�ݘc���L��AeŮ#���T��.��U����n]tk����G�7M �'�w+=3��#"��{|A�QR�7>s�[d�����	-��|)��q(`Wa�8r���h��B�	Fk�x��Hۼ�x����"�~��H0^i�]�Pna!|6��c ͥ%v���V��!�\�輍�ӜKg-nS���-�H\��m�uWN�l��{�Fu�э&ؤ���T�"g͵��s!�!2-Րe�nf�d�4=����y��6�AK�\�G�q�˔���<��6ԏ`f,Z�wٽ��<��~dB���Q����*K�A��|��^��(�	ӝ�NOv���K
pdw� ��&A�ʮ�ʖu{�Z��7�~Y=�Ջ]m������(5����Gb��J���ڲG��������g�����{���w�����o��o�����}>�O��������������/�/sX��s���X�:���uĈ��;6�9.� k���ِ]��:�J
�1�Ln��=g����R+���N����+X�I)��R���
;Gr��d�yCǴE�M���[�ce�f� ��Y�j �����ڃ(�l��#��>��X�ĥm[�缽ĨQ.�:7�S}g���DtIڢ)�q�Իh�c[2��p!1����?2|)�� ���Г+Ҵ�d���g`ؠ��-D���n�k{Y��YG1��D��5u�B:c-˘I�V�.Ǽ5�`�w]�Ѯ=�|lk��]JK���F���U.�c+�n�qp.�p�&o,����wb킌`M����5;Ek�Y���v�C��4�BRj�tt��o�Jqn�������h���,������!Y$�,h\���.ڥ�"�������h�N'�Bm�����w0�Q.7\%��.���K���h��L�[�IA`�6-ݾ�����wIG+�?[|椢+�֣6u��;�ٛ����Ǚ۽�"�!�t9.^=&���V/�
Th�Y���I*x�Z�X �&���\�}��Sܙf��\�m����]՘�ɋ�[}�
�Mf*ANt)�b8�6��J¦�)�b<2�J�`9}P�V�	B,$]�bvx;lv�o���U̴{a<�3��db"�����j�}Z��a���ʹf`�µɼ�]:�ȋ��8N�
������֕Y{�H˺�H]��Q~ӦرJz��~�Q9ɱynM�ǐsomݛmٻ�$�9��؀Ly&�ʛ"�z�F�WcM2�U������N4�p�6��w֒���u{h�bpݴ�ǣ�uۙpzP�O�Z[�9��CU�F�Z� �a̙�ޞ7-bU��!D�gWe�L4tX��jt]r���ө[�V%찤"�3g*�Դ�����Jc+��n�DcW��A�!�P�n�d��88��k����ֲ�.�u���'ji�ݮ�]⴩v�F�y�t���mb�bܷEy���od�,X��V�
*;)A�e��س��Qf�t#Ե�I�r��V,#e��!�%�e7��r�JI;N���l��L@�5rz�$���ossEԍ��`��u8�w��;ݚ�qĞ��+,�+΍q����6f�؄)Uӫ��<��q�d���u�E�Z�^7�����O��K@G#��mvmW0/��ӱ�^5��.�@z�hz΀��ۜ�/c��K�C�YJ�5�x@��h�=(�卫H&��،j�M�.Y0�[/3���q��۫Â���9��u�9Y��Q��	ke*���R�n�Q�1�=m�	��p5wv�t�G �#Zpa�9Z�}"�ó��2ƿR�S֯�*j=ݗ��#	�$�����!û���a|mA�&��Y�.�^+cT����&�H�n�uj���A��
��Q�:�����TI�l�PE�X�Z4P�N�`:)n�'C�j�)(��a���݋�z��F��PPQ�g���GIv5��Av˶���[�{kv�K�%�1�t����4���Rc��4]��Z��յ�1I�i��h��JJ1�kAV���۷&�։��z��m�;���ꍳI��l�j-��E��h�vƍ;V�+I��l�l�mSl:"t��%4m��4�j���5Uu��m���QlUu�[v�b�"�N-j
�9�}u����fۤ7���nL���m:��ܫ��e.f�̫�Nw7�S{�8J�;\F^:r�v�3���8����t�����a^޵��]�l��t{|�G3�7��(E�r�[��q�S�+ݼu}�+�(�����g�W��@Дx<e�}hta����W�Y�b&(���$�l������ [��bj�D�۴��i�����+��EY�Ҧ��ܝ��xW��{��x2�Yf�|ԃ������gSs荈���U���nތ�C�q�Q�# �ɻj�.R�m��u���s��Z@���i��* {�53���nE�ԑ�5w9�2��z�ܰ����l��oyj��9�j"�"���bĨȘf�옇}Z�T��\7�����r[BѕP��۹4�}]�xBnM�.Hp�EJŝ�y(���&z#x$󣠞J�%T�w#i�	�xi5q.Y�)�7"�gF�0I�"��Ot���$��A$���t�<ޏ?�	v������^R2�i%�?�O��k�I��)�]�o1	��.븽Н�k �O�<J��u���ֹV�V��*�%�s��dҭ����L������J`��̳�ʻ������|&��sMҊ�n��D��g_"ɏ���;�fc=:�w��
�<����OC�lH��ܪ��>�evgѻ<�	Q*�_������,�cG����Q���N[��y��Aہ��j���4,��kc�N��[j"nk�{x�ەͶ�z���)���Wycp��d/;Y8��L\�e�Nټ�Qӷ{��F�lI;��mt�`���o@a���b�����YZ@�95qݽ��}��Z�R���C�fT�ɑr2�쁾b9�GX7m�Nh�����sp�N�k�u��ŕܻ���="�Cl�ë�kxw�vu��/M�����L��ȭ��K�߱�{Ʀ@$��I�Tu��nm'Sbz�p�d�hb!څ�!&sf���n���FYyĉ��'v�5cBaMQӝ���n��إ#b��#<��Ⱥ��{���tC�+���Ί�/f�~��=�ϝȬ7�|-��#b�ϲY�uze�k�b69�ޏ?�qsϗuʧ�(_�z�TN̷ڣ�<����z�U)��,��c�Ra{ێ��]�]V[��E9�����a�A3�(���ꔐIu���m������+���0��w#=�ެ�[�2\o��H���:F�<V�ekT��&iA�!:+?�t�i�Y�;}���x�,���.���Ȁ�{{�*�t�5�4�ڛ�Q햠n�0�����*�I|�y�'��N:��T\d�!e J
���=j�fM�9�T0��u]����fi�1��/A�V�kgͨD�T2��;w�p��cS-��їǜ�͵O�<n@A+r߇b���M�K:I
�Ƹ3�KQ=M��O��G������@7�n
��T�����IS'g��(]�=U]\{#c��?�gd�.&΀ُ�p�B�)��?~ڗ��vgX��?�fz9����xŦRT�[-�,��;nS�7@an��&s�7�(
#OO��bi�����̬��K'd׎���#�%4�]��`�mq�3^�EeL{f6��}W�w���9�DA��u]]�ʮ�^�I�foF��M2�Z�r�nx�a+p��gӷf�tG������wQ�|��?��>1l6�-^K/��7�l�h��X�~�j�M����*��6�-ּ�#��F��w�ۇjT�2�z��.�2഍V��U�"���Un��Q��"���>�l�&41�s��'�o��kg(%_��4�vMt�Ck"�Yk���ܭ:L]u����T`o�y�@�v#�2�l���.�죝���d���'��)�4%�z�} ���|3X�q�g���\�J��9����3Ku��q���v����ܤ��D��;��1�<$�<�5U�o��0���f�Nd�i�)��~�F��"�h�)�-΋��ay��]�(���w8Zm�ȉ���h����	R���N;ה��>��Jo��ϩ�����dP_�.��?O.�F�aJ�_dEJ��8:��a�Eo+��ν��G��E�t:��߄V����W@�d;Kئ��k8�]^f�I���vd���'�o ��A�H3)���m�I@�阍^�_��7�ܟ喙	\O���W�o'ۖ�2E�	!r ��r�x٘��\.�]��(��D�w�!е"d6��U9̴�_�����7Ryj�߳��ȡ��=re,����j���%�2�\h�s[pc��a��	ʷ�j�loa�԰��`,�3��b��
� PY6����nK��9g܌�^��m�;��<��q�&懊�����x�R�������'5W�Rp�~��5�2��A���.��:��q�ڒ��v7�bw����w��t�=��[��­NG'=}fz���v�z�<E�U令�Ҩu�Ih��狅wXifgW���g��/�|�yY�L���ܙgw��t��g��5��k�	q���G����f�a�K��e�E��e�C<k�^m��:v+y�����%!���z���St�h��1@p��D�6rr��t��Ƌ���O���$wF��8hx�c ��"�\/[S�]O_lvu��1�p2��d�$O���Ѿ��6��އ���3R��J7�vk7�>�Wx4�+4�p��k�w	�KU2hK�l��w7�1��_O/Rg��-�S>٫}�$��y��w��Հ��;�C�{2�v�2���}v�@��=ܘ��qS���������L�~v��o]��mu8��0cwK���ac��Y����T'x�I���f�q�QY�+���z�q�O�Br�t'Ϭ/ϫ8x�;������>��8fP�-m=s�(�W��-��
��K�876Qj���i����A� ��2֚���<Ks��w����d//鹧2�:���������7�#�:c������t	IP�eT#rv�EM9�V΁��tݼ�3MQ'-f����!xb����GI�IU۽�V&�n�wR.Ki��������o��.@�#lDm��)+c	P[&|	%��G_ozx|�N�Ij�ӝ�����G7�LWnO���Yxvy+�y�eVE@���w�7ѽط�k�{�zE�w�֖M�����FO�j��&���kc-�`׋ܫ�9��	l��z��r����v�k
�C��b�;�mb)d��n�S��4|/7�M�'t��4ù��8�a�<�il�]whc�F�^���ͽ��$�R�⺒&�M��GcT�*i���f���&ډĸ\�:<�����vy�gr�����?W?�����N��,u�D��Oٴ�4�MTrh����9]k����Yg���G�� ��G(�ک�+��`�5/	�j�ZN�Zt�ٻw�y?��j��"��e�V��W?�Ef�0��4;��FnB�
뭛���>��+)�N�^c�8�`P�͝�)_�}u������K���7,P��5ѹ#�h��%���Ê���_@�p2�d��z���p���4M���d�w1J�J���;2��C�V�:���%[�n�n���ǲ�Y��6[����A,rH�;�}��C���U��7�ڽ��W�`�\g��:�09w����ȶVRח7��x:  ��T�5k:���*�<n��Mߗ:�>�E!V�q�RGF���2�GK=��n<񪬝��o�����
:�^�3ڈXJ�(2OZ?z$8?�|U�?��]~��)^t�W"3F�X��CjW���$e:14�j�����?(��|vx��mn�S������õl\i�	鮾s��Xu����_VNk�o]�)������#�aW����Qߠ��e
K�}���V�G���v�m�O.�p�����r�#���y��eB�m����4�T�5����c+����0��Щ�?����i�>�;�ي�����E�nT�Uۍ�"�ݝp�b3���ކM��9�}�F2P�K��R�>(�2�j��w�kY� �+��H�9�����vξ��ܨdA�tmo�{m�����5���>�o䦼�wS�s_����-���F�`R���Xv��f��	N�:g�J���Z�����K�B�x.����D�(��ĝdQUY���E�̧��|�{dt쮎ʮ�^�4��.ău�I�]C����fr�X�P�!(pQ�yfVtq���Y��T�03����5n�Wv^�7AN�e���n��؍@X���K�3��3�#�:g�$���䷆�c�����	�K��Yƅ�<mu\�HXCO�����a�	�oM�D����<[Š裾�c����+E�L�ד��0^���� K�`rT��*��9'^��E�qx�ʧ��VL�i��xZk��S��Ď��%R���W�oT3�\_��ۻ����bՒ�]1��muFE�+�#�T���<��i�}��[�n���^�����e��w���q,[p�#�M��͌��k��I�+]+fD+��VմA"��}�R����F�Yj�{�\�,��fh�5(���eF����_A��:��ّ`)&����j4����2p����ޝ�<�E"�J���9������ޭ�ܡV��b��*P1�Ż�rԅ�j}�ۧ#Ų/'�?^�
��y_��k���$#n=��Ԙ��u��\���E�⭔%@$T�$�0|�Z��uِ)"��5"�S;TT�[ٛ[#M�"�C�q#�I7J��2�[!���F�-v�ε+�F����wf`��-�p�#���/�J=��R��>==�+d:���e���Xs�i�y	C� ��g��*���A�J���ڒ1�������;}l;�Ҹg[ 0O�����r�t�';*�r�:��a����{$Wo\�7�ҽ�����!��]�l��k�2�C�`�v��u�w��	�����s~[�y�sr���9e��T��S�~�6�>�FѠ��I�r���ѳ�p�6�!���z��h��CZ0�Ƹ
�*j2c&�q)�Y�5��@o��i���mgEO�k�� �L����FPG��2��x�싼��.֟��!rEhJ6^�ŀvE�{	H�#w�r�v>�5���s��E�k/�8M�YЛ�W+h@?�y���������P�ؼ�GA2I����`���qᲲi㘴���}=�����/� ���Gڑ�$���É��Ko���aHo'Ȭ��1���őOOr13��E�c[�S�M뮰7o0��\k�T�i��q6X��/xrf3A�����4潼5&׹�%/�*!́���՞�=�x��Mu��+Ġ�JKi��ԋ�s l��T��:y��h����랉��0b�׻�V�.�nN݁ Tә�g��g�z(өf��3��
��s܀yA,�������/��'��F�M�V6�e��>Hk	���֜��������&=��m���I[J�Z�J�K�l�׸憛K������-��:���-�࣭�u������+]�%�s�[SW�W��]�8k�����D�An&5l����e6�c���������{||��w����{�����Ϸ����}>�O����g��<�ח�w�ً�i���7Y��s/�5�9Jه��v��תi�YP�j�/�N��ǌ�73�q�� ��(N�7v�(s��1���aԜ���a�,w+#޲M3x�e�K9Z��C(�L�hX�����ui��h�\Wmæ�$ͬ�ZRJK���x����]J\s+V�����sq���.	�]*D�f8�	5HoKZ9�5���p���-TT;��qXF�S��`=ǜ̺����*#u�#*h[���k.��bq�#�<9R��o�c�S$�F�Ʊ�*�7�nC9��3 �.�I�Uɕ�v���v��1�����/w,�H!���|oH�SH���Pr|����ܲa{�E�I^)�R,�K�Y�8T��ז�&���Ͱ�s\�S����(���v7�J��pj�=F�P��1�n �Χ��C�۫H�S��-�9أ3 0�7u,�T�e��ޙ����BƝ�u�qf=7%�Ծ��'W����gy� c���31��(�H�{g3�]����H�2f�7W�r0��Ѝ!X�")���쮅|��ۘ7onW�*�G�*|����(�D�ĹZ͂aa�q0�aF��l:��cs� �W�!C�!f
��>((�o�n�R\��0�d&m�YGi`+F��E�*'(�2��5�R�j�j�*ْ�wcc�e )���p�,�M��s
��>:��ǩ���gY�����Ok^F[l�ޞ�f��C	�D_kм�UG@	�f��������]�A�D���]v�h�}�֜���+>ُe�R��-VG�k
�;��l���B��c�ܳ%��4v�\�#tY�f�s��͢�$��W�����6��\N�wa���6�	����3]ƒ��0fP9��VEc����e��d`��;�.2�3��̭�Q���:]=���Ƥ���Z����X�,_E]�"z�U�y>��$�r�*��I�-u�óو�z�8�ٹ;xRxzq�`އ�>���f�ԩ���u�-@��sk�4�^C0k-�'3�=q�?�0d̡~y���3콰�(��9 �#q��+F��R��\���頜{%�^��H�e�l�8��3,��x�a�֊
��/m�����ٰ�t�i�;�B'a���c6��(�	�;��7a��t���b
"W0�fȭS-��齙�o�3�Iʵ��h�XV�g%�tP������[a��=�����Ճp��{�m��%Z[.�:�T}���Y�(�	�Һ�{��2�¹ �j��a]w�bZ�C�H�v�j�����w�/q��4����7NA{��,_n.*�ʓ[���B�ؾu�����.�\q��[�d�S8*M9̗���lݢ��93P�d�JRA�)$��NHw��ߟדOW�W�:���-��wd莍�E���[Z�Y�_6������v�]c���gE��[,^�WmCQi����GZ�]�wm�i4��X5�mm�b���QV��jgժ:-`��Ѥű���qqE}wL�ն�Mj�뻵��n�bJ�m[J�n��m�h���N�z5���Y��cQV�V�u:�A�n�qY6���m�ƺ㻸�-n���:ѵ��݈�h�1�� ���=���qݍtlg���{�j5E��Q�]�X��m��f���j�Qk�tQOX�Z�ŵ�u�1U5m;6�F4F�f�q����[%�Y��Tlu�cc�`|�V[@�������gAzĉ�Hp��`d���B�Q�Zm��}��ը���n�8&M���or:F��R��gє��Vrť��ҫ�7 �!�+\z���w%��WuVU�'W�U��������Dz���7�ئ|�-6Ԉ�2$	��n �P3� [�Q��x�Gm��d�?~{�RC�fy����������2��(�km����d?�r�C�[��=�;��ر��j��T�1*�����j}Ƙp�gC�o5��G>m�O�5V��qG�>�&GL�}����H��T�2.r}J6��7�fJUP�cW�}�{}a�L�8%O�eǆYoR�жy�e{�N�'�H�"�6Ŧ�뼌���3W���)��3��c϶f��w��zdT�w�y�E�?y�!"X���^H����w@�L<+;�`ͺ9��u`�6�E�����+�Gkk�^�G�cɰ����]�ӱW>#��\ئ�u�m��F��4��hy�w��V�'܋Ee)���K?�tj	�>8�����X'�:;�vgGke�*z�\{QB@�C��$���fڑt��K�M<3<��E4)ڽ����AB#x=ܺ�Z"�'�HY@���䍁'n�����p�g�g�Y,r_�O��y��h��9��*d��ۮĲk.=7�B���:�f�,��[C7������,�����*��_�Eu]�A�hդ/��K�a���U��|����w����b�`�-��Ʊ��ᡑ�wlVv�	�aN㞻5�Gú��6�7�T���jhG�>��=�T���P*���#++��'�6�Y{�;=���՗s��p�U�����EH�n��6��,a�"e�[���c6��8m��G�˒UA��î�N��m��ಛT�Du�mHȉ�ac��3�b��ٞ�lO�p�X=�N���ۅ�.��s���qu�خ�iμ��NA�o��*h#K���Yϝ��w7z��\7`��nr�����r�D-�����L����IM%ܻ�
zC-؎�|�����<�ܓ�y���	P̆�2��a+�DvH�4y��;��Z̓4i2�1����A�A�&��w����̚��b1@Cy�F�n=�iWG���i����R�I�wr{!���C6Cm���p8)����Y�g�_q��͆Dp��Y}�6�	$
��+�?��V:�s8��Ww����]a�p\�ò޺7���;�հ�ິZ�����k�o=f����r�u|(�K45�	��Xv�^%�D��W����S�;%�Żǟ L"&�6�p�f�g}Y����t�N�Q7-j|�:0�c���d����.�Z�|�:����q�v�����9ӻ;�7js���P1�d�7��Ɓ6�tQ��02�-��;����`n�eX[�ך��b�{u�2��q"|Vx���?4r�T:-̕��(��y�Y<M�OWW���Dz�(��∛��e�GU�ATD�.�/]*z)�2X���_��'X]�+r����
����3g�2*u%�/�=B��j]���vw�ޞ���;�`�F���Q.hag�
�� ��#֭�\��ΛJ����3!����3���J�AG��}բ~'�!��p��P[���b�H"��Om=�x�I�%A"�9&�)mӮ�ȑuݏi\㬾��ݬS�A(A+b/�}�Q�ܒV�*BDϛke�����ꈍ�2�U�w��2<��c��ڕC��\��Ԏ[jR��7o&M�ˁo�8UI9�א|��0��pKd9�oG\x�U�U@��K*z<�lif����\MȚ�C/.N��M�zV2�XS�p���ht\�*�b�P��LY�ZkE�tNu�B\o
�a��ᆲ����e;�S�js�CHG��q�� ә�2�q�Wz^���^:Z�e��e�N�w;��§e�ޚ��>���'w:	ܮ۬�Wc�=��A��侭��AS�~&����U���>�$����ޮHq�f�U� ��0������0+�;\��&X���g�37��1�o �w��Ou+WA� Csi�n��z���u{�_z��v���\�\�ҍ'�0����o��Č�#��и�i�u[�f�z�2�
Z�d/2Y�3o�&	#�������ܽ��mtO�+9^�g��Y���V#�������O��ȴ�?ɩ�G����n����"�_m5���CS�V��n��:=��3C��n�K�P�v�i�|��ٰ|{�H����=��C�J�ML�y��k���_u��4ә�%��JV��}yjni���
qA��h)���i�Y�gzq_!e#B2#ݤ+�䕣���}�4�b�����>��K)��g� ��5ǆ"�R�-�ݾ�qM�Ո#]Ka����A.~,R�W��e�+����{�E����&�hɫV����g>Ce�#����(��Nl�ת�[^�9э3��gB(o�v��3����ћ���v۹����c��BB�:�m.���[���_e�ʻ���37Ӳ�'jZ!6��hؿ�`���T��q��܂<��<�BP��n❟T��z9k��1�ٷ,�ݭ] ��*:؈|g�Ғ�Y�,�Y�Ӛ�]��ϱսP������O���ĭ�zx.�V:����E�2���2n��#����d6��9��\y�l5:;pY1�2��|�E��0�x��^�k����]_U���:�$L�t�GR3 w7G�WC�S۞���r��Y��l3�([��N�KV�(�xbIݓh�i���p��4=���K>��]Yxs�ZAƝ��}�=;}@wԑ5*_�9�\���[�8t�?>���۞#�=`8:�\e�.���1~R~��?��ݟ�#&�8KAU��҂0�fDye�7��d
��բL�B�;'�齅$h����9с�³@l�U�ѧ���G[ӆ�,Ԃ����?[��8����$�g��}��֕Wذ�y�l������P�rJ[Ǭ�2���΢���`�
�pV!�M�;��'�:�2qV���m�X/f�6�����E��e-��u��:U�,T�J�W�Qy���/����Ở<�gLpi�@�gb���p��]A�|�3�.5�}+����ڜ�� i{���ȕHr�"���b��K=��/��5<����Q�����>�S�7.=��"��)o�GFm�L����\v����J�ӝ,x,�O�љOV���j!^���J�֨qA�N�âά��ͪ�SNd
ڧf���>��^�Km{�D¾q-*Sv�ps�\�`��f�Q�� �܍V�j���9�5ԭ,i���b��kd5�G���������%]�I*�뎺u��l���ye�����.�����'��5�C�&Ԯ)N%�bx�������轄�����q�zj{��V��$A �o��*i\������?
������۳��ۧ��{�V�"�5;���OP�3#�lOZJi.�����|sh�4���#d9���MDxf}�ٯm�l������tkty>�ݫ)+����A��A�Q�;2�Mx�^��+s�g���n�-����l�6Զ�Q��c���Y�nN�-M*˧Vs�\x�[O����R�h���r�� �$U�<�f����g�����ۜ~�o�
�ݮx�F};&��;*�rJ�L�V>��v�_���͉q��Ë;9O�`Fl�7q�is��ӭ'p8���B�T0~�M�'���^�F�O�w��Y�p�
��O\љ�7���/V�oW�����a�=!�����s8:i�kY�"��v��I�~�a��|2R�c�t�d�p��� X�c��8��v^�	�G4VV��3Y���i�Z��ϷLfYy��E Q8���ъ�yy�>��s[j�v�\{����`��E({�jf��2�Z$u��HuԆ��0�$䇜7���_n�&���o�8��=�\PJ�ODY��R5%��}�1��4��wf��8ᗊ4�[/�ih�20���,A�;��V���i|1�"tc���RLwmEn�c��y)�Db2�B)�T�3�^��:�Pn�|��̲"�i$=N@��W�������g�Md�<ֆ/3�G��F�|2�M�K��2�]��$�v�ߗ�ڽ�"������9���Ô���FԼ�h�`��G�YѼ*iW������cvl��lVx,X�j�F�}+�I�	z���'t�w�}�_��z��p6�Q�1���.I���r�H��'-ԪL�-�p���\(��)�:6ۄ���;�AR��$�&���lY�b�ɽ���ώ�a#��2�#c�fQ:�뒏B�17�4�g�K�;���ٽOd
��1�	pB9/��<.��=@_%Tqts	�xG��/�Tul���"��A��B��l��6��H$����T]���;���ƿ)?�vA��!���c�#jk��\�x���eN�Z9�s���-�N�.�d��3������ߘ>�`���ؘ��v����ٜ.��2�*.�uv�i?NP`�7>Wtl�ӄ�cǚS��i�	o=�Z��]���
�<m�@�b�e�I���rA0��cM�h�QV���uEu�
�J�'a�W�0�xVv+��:3-��w�@��{<�`n�.lԻԼZ����������-ψW}����RE�Ma�ý�v'���y��=�����,5F��:	§��=1���iٕ�;{B%#01z���~-�u�@��]z�D�D��'%(��)Z�-o&��ϵ��Vg��8�o-��3���f�D�C��EG����2ТC�S�W]{���YV:ד��t�v`|��4F�M׶��x�O�a���[�8�(<K[d�����L�����<R�(" �JR�k�YsNv�g�i��G7��3b�g�q�RNwTd@�!]rF@��hT��Ww54�#[5[J��j�%�ս�� �$�Aߞ�.-�V=�� �:��EIT"d�|���������� �T�L�Ǘ�%lD{m��Ғ�1��EU�# �U��#flٮ�T�}-t�u�L����P[#�O��
_�d�2{6���b>��	�O˺�V�*Vv�W`b�~��;p[1�v�M���P6-zZ쟖�����2�Nһ�{�/�Ŏ��WW�^2+q�ڞ���5[��)��cQ{a�+�dO��&=�@����_�����JC5��7<�]Ub���w�Ҭz�����dj���y��� :;��y�Y����r]>	����ɝ�O�dZ�]Z��<�Q�������İ�}{)��G��;��䬒gݽH���8�U|�yz�e[�(v���;��vw�'3�X�ʺ?�]�"3� ���w%��548�wuw���}���7;��jkq<�+�c���8�g�2��W:�kW��$b���.ɻ��+�3O��d8�4&r�>٘
��f�;�YS':fv��(o�@i�7�$�}#�3�vr;�#a�Y��Iޭ���n0�T3�M4�ӝ��I8�oG��G`�>ȧ��gB��e&�x���NsTɫ�ͬ1܍�EĶ�ވy�MhO"�YJv)�CUf������S{�m�;�F��]fצcɖ�jH*�;���i��F<$$�wy=���N6�1����w3hע�'Q(��J<s)�%�Ec�����������w~9v�i�}A��P��xG�j���Cja֖G����e\��N������&���v�U:�*�� נ("�B+���W��o������|}������}��o���Ϸ�����|>���};����m_�S=zz���s�tB>�7�98��ܴ���8�]2*�9�#�X�����l�u	�(Z�t�5���{ZΪ]f-1աPB�e�
�}���(c��ݰV�8ӣ0 �h��<ݿ�x���W`w���X��nj2~��6�0���-�W��2�½��I�����u�K�%p��*pI_e'd��{�;�GEG��.���#��LXz����n����Wz�p��	�w��
��oi�j�$J{t��\^�}n�!���&R�Y�W-q�
x�K��oF2[bĥ�M�@�٠I2�䘀A�rJ�{�7A��i
4��9�@�GFu�#��ʸO&[��d`���.�R+�����l����P\9;!���Ӵ���9Z�1oJgD(�0#�û�(dPN4h�ٓ&X$���[��>���$9���M���G {l�KԔJLމ��#�6
�QX�n�ݣAt닝Jڳ�����u2����m:5��.���+� [��ˮ#�Ն���'��q<l>��^c�RY�N�����3�_T�k��{��C'iJ³��c3T�Ұt�`b�xo�:-�a��|+�g�[�P��u]s�G8��9S����E�$i�.O���Y0��z���9�m�V��IV��G��R�ܱ��kG�$�#�K
���e�jn��!pW��b���<=�xކm�ǫl<s{j�j�̣��]�Ej�F��zr�˰�\�ek�y��H�> J�\��s�ODb^)9l}�	a��6p�{���`����Iz]fgY�ƕ�9T��#���2w���,����/fD������ܠ�WC��kA�7�M�ࡺ�Лh���[Pu<n����y�����Y��x�2�t7�uowe��S"��q����	��x-]�-ɤ��q��Wt���R\qZ̄r�;h�C1�3���ټL�Rd���5�Tu�]�-�k�캙Z�X�鷫���3hl�uƶ�h$��G�,R�բ��|,7׫����6ЊG+%�� (���^�)�s�!���n���)�Mh�|�[MU�wt�_!�:�u�<��V��y5��aKOSN���x��Fp��K���f��3���Y,��v$���]eА��l�άKp�@��[�ҙT���7� |��5���s�Ğ�wG��͍Uw��+�>�Pf�]vXyj������e	�c=���<�����Ze�ф�ٸ�օ��(F�)��8q�n�]D�x�&�:MڮJ�x7(i�	Ү�R�����Q+�#w��;�r�f��ZYH��C]���ח*O%����e�������§:��,uA�۞����s��C�]��V$d�\�jk�	Ĝy�!kJRA˓�HRRI�_���AZ���Z����m[��zޞ�i6��A�4kmiѦ#L�[X���ݎ;��cm�j�h���(��mE�Q���[&�i��cEj��Ez�Ӫ]E��v�k�UMWZ���]����i�ъ���mLQVڢ;`�޸��A5����kh��d���v&=N&{(��5�v�UQU��P^�jz��lѬ�ڶ��+���fgX��j��U�lݴS��tb�4Vٵ��n���fm�6�6o��z��j�4j�h��jձZ��j4��qݳk;&�v�ފ"�*�h����P[kZv�AX������s^��Gm�d��Q7�Q׮zɚ�Ѻ*����\��D�Ov�#On��X�.�PtcF6Ŷ�ֵ��bkb�3>���}z�ww���Sya��͵��z�2:c[�av�`G��5˧;N�k&��6m��k��A�4>������~�'�Ǣz!�6��Ɖ�1����I$����u��l���ťQ��U���6��2&����Ƽd�<�l�f<��s[ѧ�m	$��faင�~]����/ m��\�e�s��Rl��N�;�h�R���Vvv�ia�@�9� ��g���<�}ֶ'�%4�pdٙS��k������d��N��ų+a�ˍ�b�c�����{_��C��1=$��y]�S���^׶�8�p�#{�����2�p7S�X�*�i�M6� �uO�Ƶ�P3d6��������FN�sD5۬ͥ�{���F�,+�l-$�v�u1��4s=�p �+6���m���f�g��)q���r���p���>$�du1�VV�ju��l���v?0�#�����ӱV���̲�;��Y{=�����}W'��E��f���u�`
���n�<���U���O�*˖���W3/o�(5m��]�0k0����6�N̶��-@��S,������� P���Rp�c���6�������VImg7W�E���Ï��HN����w�\[��Cc���h����̸�~$u���)�3̺MS99�ٽ7�]�v�������KX4i��7�&5�PR��7/v�4o���}�È��PH�I�TK�Y�
�X�;�u*�����Eؼl��=+'��YR���Fh��yUْK
��� ��e���uL\^���U���	�f��gͱ��!qR�T�쵻n�":�Gc��qP7v�:w��Dk�$\�8����	nH�5��It��
`<�������+ �ө��@r�}l{lʮ����]@��xƎk��m���}۸��m�B�:��{�A�����vE�t�4,����	��Ǌ�<wN�oV�ޮ��=���ɫJ�c����v��+yܩ�z�a��L3n��GN4��n\�����MS�ӛ����#��~;<�}�6�n
���a�pp�t�b��y���N��{�GL�ufOe�L�F1�����f�_w�nm���u�����ytw�e`l�f��[(��r��Ch;,�ӻ�;�-.ڶ���6=�A���frFZ �+)�vW[��J�XTOHO�D�lݷ����kf�5���rN,M��Y^'���WA�=M�4z[�h�}���j�M��u�E�8J���\k�"��������4��퓎65[�;���=��Cx��-�A�����p2�4L�A�STu�����l�n�ע��+�65ۗ�h��Q�d�#}ã2ڔ�U'��$樼'�:q�C�;3npw�		&Z&���}|��@B�= ���W\U+I�uW��5���a?R󕋤�U<}A�~��;S�x�r	b&:��	B�GEQ=y���xD�l�qXy,�7����[��/-O�i��e�P����mW.5��A��u#r���׻���hʡ܃�o/�x�)���5'[�٠�������ɹrDXD��t���Љ<�_L�]ZKw�ؚ:�V.�L߶���
�1��%}�D]������6��?J��F�VJ㾩�g)F
��uY����c'J�n��\p�`�vo�gh�4��KŹ��@Y�%��{��PBV���n/W���{+^�F1Q]f�ҝ��L�A��^l���[I�p�ݜ�H��B��,��若�Flv����$����\��������#���P�jC��cK1��o���{���Ҭ$}iE��*Vvϻ��1m( ��d�;B̶o67�7:�o[�y]ޥ~ZަV�3���	�?o�����py@���n��kv��t�9��d��;N��HW~�$�v�������q4�q���f�2Xpw�#�lʟ��ܗ_�&���9�ח�`�YD���__L� �'��7��8�q�Ϡeǲ��{�l��Ǎ�{"��L�n���;���)�0���c�3��B1��3^Yl�; �Ȋu�%¾��|{2�l����!�#�2{E��z�?�����՝{�������晜��+������D�cy��ا�q�؃����y�Q�ۦ�E����;�wH8�ĕHo��VRח `
�C\fMK�ʞ��`�BDy�[�L��G=2����$"A�|�+��gg9�w&TR%�;o	�	�U�7d��Ya�A�w]P�W[Х��-r��;�Ϲ"��W�Md�8Um��R>�]V6�,>�P���ӎ�c�\��]�΄��ftx�(��m���~�d�n�lMv����!�8�T8̫�)���73���L���i�c,��9@{�ud�\d� �m�A)����/|�vοN^���GmR�ve�uB�U��< j�L�˪{b��NQ�l�N�鮡i{�OPHʨFg�n�S��g
b)�Ȩ�ܭ��bz���N������ɹĚ�MU*I)���N�ix�3f��"vQXk��ܐ�8�ddns�AK[��KzI�����zjn�����3D����;npXP�R#�ֺ���J���b�=��m!u��>����&�~IN_�oC .� � r:�D-���݊7�kbzҕY	�gsf�ȩ݋��G6�[n!���Z���q-p��q��`�s��}l�.��B��L��;�u�]���M(��VN��1�a����{��������q�@*�#�cks����EF�{���T0Ƶ�7p*��9��*���b �6�K�P��*����� �(N�[�R%�$��t�.#�wj�*�D���阓JY�B�l6�o?9���ɣ�B�kLo9{4=�8�:/:o'��]���|i>�'�x��2m�|}�#��j|��W�G��s�3�v�%ೢ*�`�+�l"Ggs�eqU~ڛ}�G?<õ����
_���7V����tw���op��xP�n2Ih.��������&?�7Ft~�q.N�3XN��x�#b�����/�H�Q�S�����hD��f6��C���齞�(�(�{�jf��2�zm(�d����s:h�i�{�ok���gڭԎ�q����:�͞�x�(��K�a\�p�M摇�W��dQR�$�8�TQ�����p��H�YS�սS�7�o��+�ħ�����%zMA�T{2zi�M5��vf�ч��sVso7zĤat�\ m����CiHߘ�T*\�T-6���Q;k!Q͸��;T�gS���[#�E�m���ѻnI+�t��|N ��e*ӓ��Oܤd�]BP���x�o�%���s)lC.�b�nftd��=�>����̬��5��X�YH� �Q+5uP��AWftp:C�P�_�-}=j�l����"\�P��k�(��~T�Zt�㧱if��D�$t�A�Ox��z�����?�/��}Z~����g����M��⠣#��r��>�?f{��HZ_d���%�+��U�������� �磅��A��1*���.��n6{e�7������:,d�j�՝{��1� ei��&�����*s��������R�Z�ŢȪ�����{�b�""���'��$�.l�����ҿ*�=Cdu7cϚ6"&�U��g�<x&PI���ß��=�r�}^:��?���\��y�A�ԫ���w	�3�F x����]���Mx�*���ph�l�G:8Eȏn
�������,Ǟ7�߇ty�)�|�!ެ6-�O�����/fv� �"x��tTk���^�!f�R�j-M-\{���6�%�ޓɢ9�{���F��O&��S�Oa��p��
��1l��.t���=-��fT�t+%*���K�S��;����!+�f	���W3zb��`���)&����w|9�9x�nv^��Fzw\"T�m8:��޳Ժ��UcY�i-�2�&-Y\���7���X�>G�[�Gx�l��d�6�1���X�F��i҂[c

iR�%����R�9�gFM!�\�-���Nӝ,xs��:������!Vw$�Z2����a��h�>�9��fd�;�5Q��S��d�,XD��t� ��|nk/��;9|vo��5�(8j�n�j<�b�]FH����oϧ��vZ�o(��<ڻ��gM<�V��� �������N�j�E�tWF���q��&`�u��/����}]�z	Q�EXl����-�� J�a�:T�njz��|�p�.�^Y���x�6�'����!r~�g���Lb@�Uh}Vvwc�-L/�#�ߺr{��䒺_B�;~���SK�lH��j5N����T��������-�oW��RK0gE;�nL썍��ܗRDԳ�m�[��e��e��vN�N�ي����@�2�q�k��3"���ͳK���{����pFbgCָJ/hn����K�����ovP�޼�.P|z9�s�vem�9��l�,z�5�_�9q�
��ѯ�+�X�>�Hs��Ļ��T]���r��`kIV��:+�|��}jSժ���=���+�#��h�!�s�
�<���MZ�ײ=
H�i���wV=I�׽7Ј�Hm�m�?�!�K�{ws���Mw9r�_q��N���G��~�9�?c��7�Wg��8�g�wF[�*�_��D	e�������μ>�'�tlvZyĉX��ͱQ���ȗ۟������1/�~M��)�&�����;���rw� �*��[e-{fs�h��ܼ���ql�%�{�p�D��OV��Ԑ��:x�X.�g������矒1���z���/v	j��VM���B�h�ó��2���v]�6��'�v��.},��A���#�`��j�fŵ�s>.�[���.+����JFQ�P��;w��`�g��NEc���	�l�_i����}aKT�ta�m(�s{=$٥J��T�S���F���lV���
ڎ���}㛧�YrD9�˶��wIHr�28�˨�7���轖��{��*�ɓ��WP�D��2�i���*����]kk*��$��]~��4^�z��h	�֤[�h��Qΐ�,���*H�"�N�y�-c*�q�w{��vP�TŪ�_>��J�nӃ���z�*�L{�wa؝�ы2z�;wҢ1Z���[m8D�A\���F��q��7O?mvoS٬� qn����[Et�-�l��b��[�%r��y��l�2r�'@fW�"����vmtl�\n#��]���6����4��b_��>���]�T�����d���o�F���E���!�2���̥������P1˨��������}O����~w����5\���2)"�ٜ.gZ�l�a]��Q �����ބ�{"���o~H�7`��~�U,}c���\��R>� ��}��d�f���6�O������P�"��<2�Q�9Z�H�2���$(�L����ӽ�잇��0׋����3{?:=F#�U��f#Bf��n^�Ɗ<�T���Cv����3F�h�:Mɐ0ۗ��y���C��������ײ?�
 ���*���{��Q����SOG��|���Рd%�fE�eY�f�dY�d!Y�f� �Ve�fE�F`Xi�fE�`Y�f�e�f��fQ� �eY�fE�VdY�a��f�dY�fU�d`Y�a��FeY�fE�a�f��e�f�FdY�f�FdXa�Fe�fE�V`Y�f�`Xf`�f�dY�f�dY�a�`Y�f�`Y�f@&�dX~~8>@@�03 (�2,��̫02�Ȱ��0,ȳ*�2��3
��>�.`Y�fQ�`Y�fE�`XeI�fE�FdY�fU�dY�fQ�Q�dY�f� �F`Y�f�FF`Y�fE� �`Y�f�dXee�fE�V`Y�f�`Y�a�I�fE�FeY�fE�F`Y�fQ�P& &UVBV�D��@�Q@��@�O�E��s(��a� =a�}p�Ua�U�  �V@@ XeUa�U��ª�*�� ��2��ʪ�*� �Cª�  C*�*�2���!���*�"�� �(�"�"�(����a�a�a�a�a�a�a�a�a�a��Y�f�eY��P�2���
������|߷� ��Ҩ�0 o�o�~��������������|�����`�����!����T������G�����@
 ��������D~>� ��@� ~���%�?�?��~�C�@P_��'����H��������?���>��_��`�C�X����G�PX�P( �@B�P&@�T@�XU@�$ BQ�P%HQ�P!EP%�P%U@�a�%%�!� aaD	! � >R���X_�?�{AhPD�@(
D�q� ��o��������=��>���Q@p>�����~����'�?��� �����=���P_�=�����{�'���
�� U���h���������Ҡ�+���	 U���&�����}�^�A���~τ���$�:y�<�= �
��?�����~�� �
������d����������?��?C����?��$���C���w�@(����?Q�����@p_A����h|�&__��N?���V�?��������	>��
 ��53?_G�C�@~�8?��>������b� ��I�8?7��D��������?!����e5�l���Y�]� ?�s2}p$a�$$�Q!R�@O��4i$m�R�$UP��H/M]��Z4�"EM2$
��%m�
kER�Z�R�$��}�.�FͭJj�ɭdZԚ�Im����k	A-4Z���km�i�LѱM)J�KMfjі��l�*�6�6�H�Zdm���j��1�Hw�fk$$�Y�YkUJ�M�ض�ֵMZ����ԥ)U�ڱ�[-��ͪU��U���2[J�4���%kjC)����6����M�ڌ�b�mZ�Ӂ�22
��  j��|�^w=wl�N��ݺ���w�랝:6�W^�����z��v��n���ޭ��^+���CM5��lwww.�5�k�s^���wvu��vꕷ@˵�κ�N����P�M���V�V����  �\=
(t4���z ��=
B�뾾�z(P�
(<��(P�H�WO�u��^����t붧��˝.��:��tޛ�Ǯ��^�Gm�z�M6�{�ދ����ex��kdm��-�����   ��ϯ����m����S����]=�{��޷S[�n�@VOW�zxSv�N�k�g{Yѩ��uo=o{z��Y= ��M�u�l���
t�G���ݩ]��9� {F+&�Tє-i�  w�U5����wս{��C{z��0MR���{o*�l���{�{޽���:oK�����kpB�:�Z h�-� 5�u��F����l�-[l,%���6�   ��*�uΰ�il�N�(�W8i@*�,�D��� �-�U�@7.�4�H;K��@���  ��픭)�e,�������  ��Q�� wawQ�P��W���kB��͸���D�������e��
�R����(��pV�v�im��U�b�kB�m���V�  ���@i���kB���ű�	���Glm9�t�>� ;���]���� �:{xP� Ł���sҖY��F�l�f��,a��  N� P�w�  �xۇJ �ظ �Yӝ� �{��tPۯO F�={�\z 7a��g���y����y�ֲ�d��cL�,�ִ-�   7W=(} +�X�z ��c�`J\<�@�^�h4נ�7= tn��׻� )փx1҂�iGzS ��MǠ ��̑��XV�kYYY3�  ���(PQޯW @޶�B�h�á@��p
 �/p�=�Fy�z ��հ�4�p�n��w�   "��1JT�� ѐE=��))P  "�������`4�S�����   �� �#M 4 $�DM�R�  ��;����o�ߜ�ߧ��'ɹ�gJTּƛCɷ��I���|�[�'�s�g�Zy�I<������ !$�H�BC�HI?�����`I�I$$?�������a��O�ݹFXv(/�� �n��6�AV��[�ټ���1�;N70YJ�{r��'5���b�1�~7�Ls/E֪h�0\�P��w����5hy{z��]];����"�7*ŭ��F4=��Z��tGWF��T�\�T���%���*�f��;���`�b7��<خ0���ˀ���ˑ&+>ӟ]��6�=�m���欂J��t����TF������\3�l�V(�k��2͝b�[��T��:[���4��fG*��t���y�5�r-=8[�ݵa��S�"�&�6F�Y��'\כn�F��z(����4�X�Ku�S�V~�n)�I��90/�`4��Na1D&%>/�I�B���ˬ�,�\�� {%�J3�n�u2��������\�@}�KHO�+"6��?kIH�Ȣ�{N�%1�6N�<ʶ��f�%��²���e!��m���Ez���f��n��w�]\��t]��H*v%���4.d����)���[
�V�U�J�T�#��OT6wkI����N��Yk �4ǩC3�2�0SktT�#�n΋7�$XNG��yDۥs-kR�W����dJM��h�r#$�Wm��v6�{�(�,33li���uxA��k7V�o1����i]	�͇g��/����kE]L�̍��ۂVZʖQ�ݧ.��X�8BՈ�R$J��Ã5D���l5�4B�;Ske�݈�:�rJ
9c353u���YYYM��jZ�&�,a
E��+V��BS"[��sjT��"�W�"�=3-a۩3�H����@Cb���D��t]�5 ���޷Ah��	GV7t��ug��B��W57�3+r7,^�[VTV���h�z�Rx��nL�u���򡆯!f�v��1¥\0^��t^�3f��DW�- �ip$ڧ%���JP�]��g(�8�ڻR���^6�D�z�̷�U�Y�������Տ5T[��	��MlkrVpn
���nV�� 	��r]���� ��V^'��A�G*U&�
�%�[�W�!d�`�l�]����ӽ�c[���b[�es�����t�.�sE����V��`��@p��.�m�F����Ɉ��G�'��-/�Amd�t0 *��R�å�j��# 	�.e¦,Q$NI�60����q �����]'�&�|�	r�rO���5�[�F^�0��͎�)�G(�u�h2�k�]v��S3N\2�+���۩۸S�D���i%i��KS�W�q4��$�:$�f��e�婻r�V`m囑��d5 {�*)yt͂��%� bΨ��DRd��,"B�mI ٪��6����kn�@ժC���^�����D��B��̩R��v�޹.R�MV`B\�%��R��r�ߞ�3&�R�X���6km�͕�9��Hbw���^f �f`�W0m<���a+�%ڱ�r]o,�,��Y�K���~jr�)�,�k�.����<�&�Q�Bĭ*,F�J��9�D9��r=�@��>۠�Ǽ��T���X�J�f��Zn���NA��6ela�.9{�#Ů������sX�f���K4J0XÎBjd¬�G"S xef��i�k�.� S#0^Rv��Mh�|k2ִ�<.�\�
k��6���Ӭ�n�U|�;�k��ai�c��ir)*��GDbହY��r2��0 kR9�����F�u��Z��২����\�vU��Gb#Vͽ�^�$��֛]����[.T�!�k%)��Ud	�,e1�,p�+/ ��g#4��5�ZVe���1LfGr��E ,�2ћeѩ*^š�RM�ɘv�6n�z۳D��%u2��^�j�2j+&�z6Kd����2R(-{�1\[XM��x���;n�x��귷Qۈ�E.�,�/#�=����{�H[d;���:ؖ�
yW�$�[M�����M��V��X�38S���
3�QԎ��H���4��� �Y�Z����3d���n�e�,l���G1�a�MS��U�55�Mw�M.ŷ-�nl'V�2�z*�L�ҝm^����C�ї����R�8��n��L�EޠAݡwov-�-�6��ʊ����<�f��eXu{��(EA �\�����0J��L�064��,� �.��,D�3�ܶoj:�D��|��	j���,{���c�4֪"VQ�3+#�`[tc�o^�d���kr�E�*���Ɖ���(m��@�p��fà�&�c=���c���l��6S��옭f����m�(mܒ�9��͸\T�\�ƱX:�U��&�6�tE��+D�x�1�K�l
���h��R�Ʊs��b��3\d���[c��bddgfQ��L	���׏k��5���7�����i'�s.鶭�VIR�SoVݨ̆k/YK����Pj�^^5�@���!�L�6�i�]0�r����r�S`�L��G~ut��\��nh��鵱�Vq���ἳX�׃%f!B`a��&�Lj�mCO���+A�JC���#���]lQ�dz����dQ曖��QqE�Թ�6�q�A�����oq���w���Ѡ&e^(�\��b�a����-�eDI����FӼTӴ�G�h��Z������^�m��Xu��Jd`�`��fH@���i�˴������scЅ��@3&C�8ժۭz�^T,K�X�AG���X��i�(��۷��2��eԩ��>�������/�U����-́���n�6��ۧ��Ze+�n��X�j�խ|MEmh�v�5��b�g5�#wF�M�S.�j�$�� �meӓ��
��7b��T7*`Ѻ�\@r���N�W�.=��M��]<���%bd+�p��B/7��t�43�흧B�n�wRL�/D���rde<Y��N)�t�mEF�M�[����e�w/Q�c,�*Q�pJ���Vekr�I���3gV7)�,f�ܳl�
:�d�)cAnC�F��R�d�v�m��V�� `��kuX��19D3�ij��9�Z���m����,�� n��˺��uk(����C��oc��k�TUs	�[�^n��4��M�0[Q!��J����*b��1���:8��A��~�"c)Mƶ��bh�բ���"Y�t0Q���n��L{M��b��r[�-õ�F�{`)�67N�/1a����m�;���f��Hc���BY��iԱoHF�$��ܡ�q`!�3Dw�J�f�,�%H�/l���JQ��ToY
˼Z) wXp=!Qԩ+h�f��n��D�N��V�3��^�jЬ
��X�EEW��\dJ��Dܡ��<�F�o�d�ШnJY��4�J��z��c�40�M&�8�Z�K-�.�nкoj̽��%[�q�BB�GOh�n�G�E��+�v��E�0�oh]��֔t����5h�������V7(�O�bW{{C%#2B5�IQ�F�^lu�!�,��V�*Ğ��Bq�G�^+^�2��]�AR��)��6<f��\�6A�Ķ��5��I�!2�*#e�����qk��)#�ַ��V�����X�Q�1v�5��l�2d�ֹeh�e��r)),��(;H�Y��76c n�&:U��EԶ��U�u��Z�X�2憫Q5.�ڗ��!Y���{��Z�kr%��f]ڨQН�%������v놾�v��^'����Y�lmb��g��%�S�h^��4eɢef�kZ��Բ6QN:�H��w�q'�����TFj{eU�&d�aIv��8�q��m�r�j�MܣE��b�nU��u03fD�+�Z�u>ko5�.�%�3��!���E�lVpܓ	��.,l�Dޜʟ,���1U����K,I��ًc��.���4[n�9W�ڣ�.���t�)�ӜKkv���C��5i���	�IS��Ғ�X-ƶ�7[g �t���'�(!y����^3��ݴ���X�Ĵ���)�͍���Z#�Y*ˉj���ڃNB��fE��]3*�Hzr�ր�o��$���R�1�,�����r�Y,����#	�g{����W܂�����nKI�m얨ۡ2�\�ؤ�NR�Vj�h�	{F��x�&�kW�$�V��7n���Q�<��Ncݱ%�-�bIS]ؼJ��/n��3���e�j�q]�$}y��H>�!��Z�ǌ�0!w9���ǁ@��ۥn�lr޺��R8�����9���2,Gn�A��]m��t)��P.R��I.��Xm�*��S�/Y�d2����L���K�#kH8�{00���{��^�Z�J4�f˭����g*�>5����Q���+YB�V�2h�^J�ؤz��2ҩ/M�]En�JQ��;��b�굀�5-ò
.;W�*&�D��f��P�%��
G�ejڐ���M�Y.޼V����҅����76�D^V�L�˺7Yu�����0��ÿnf���p��QՇ�[��͇Pa�8�弘�4u,t(�ȵ(�\���B��
�%V�چ�j���٬7Tô�Q`����7�n��W�5�E�r��S@u�t�M���<��3%irл&��N-R-�-V�.�loi�*Q�����V�+ð�j�lM��2F4�D�E�J�s2�b�opm�O6�)6��[I�V�s�D��-�w�*=wC�G�S�ȶGqŷ�*�e�im�J�D�j�q���Ϝ�5�q�j�*�>�+�+��d:� <�v��f)���ͽ�c��k ��Z$nc��f�l�e&S���:!Q��*9X�K�.�*ml������.c{�#�t���,����]Z�&��3U�i�f!p��¯�^ �	���'��S� �i=�wv�a���lޥiU��6�0�
�vNV����بl�y�C�nwX�ͥ�)����m^��3r�R�kv5�I7�Y{+pY��5�2�'���)˂`�lTm���3
��N����;�0;6rRUf��E�-Z8+CY�Z�<BU��V�L���2��� +�Oj���*TuV��%��i�Po���2���*n�3y��u��1�+��C�{t��r��AЭܗ��+uF�
S:���@5���4��t)���Ŕ��Z!q���Fi���Vͻ�NTF��eT���V�ݜj�T���Ы+	b���4n�S`�m��i5�ج��?@�ҧ!��L���ݟ��pe�J�0aW	�5�A�!d�J��njHD�O�u �����.Xq���hV��o �A�s&���aY��*1�e0��a�T"9`:̷zhI�^������Zp!�r��n<x�ł�(@��IR�]R�&��P��'`p�;-*�Ŭ% �C�,�oX�1ۢ&��#dXӼ�0��J�
=:rބ�2���T�#G
�yV�7�7Y�$�e�j�@2��Ե�X�[����j�"��#MH�Uei����&�)�����zي��\�����Y����W[$oYm*"��Y��p(t���P��qf�
P�����I��^��՘�2��2D����
ڬӄ���M�s	�SQ��^��ڀ}�	�GL���$�x�:�9.��ZE��!P�Ys\�Q�4���&��ۚFL� owB̨�P0ŝ�kcGtڀ�Ӱ��`��z���r���0Ѩ5b��ܒ��lݙz�k��Ƽ�va�ti� )�dͰ�WY�80�4)�d�E��ѡ��[MPZ;lV�ԍ�a�h��<Tݭ9@R\�c��)G0]k�h � �5�n!|�̴����Ў��RT��S�[�}�VU��nJ5r,0�C����լe�y�7�%�7���[��f��B�7*Z��X�Pޕ0LW�@��tL����b�DH��e�L�/0Um'rf&����Yk]Iw)K��h�3�X��>�V���=R8��1�m�/\�)2%�E֌�5��T�J�z��'�-'�[r��ATNm��M'�Z#V ����E�lm=��Sr���'خ���Ōn�Ne��o#F8m]at\	�)`�se<n(�;{�0f,�aIV�vL���QU�L��
K��{q6��B���9���W)��[n/�X9s5�i��pLt-:��]�a�;b���:"z�-�R�����᡹,��5�l��5n�4���]f�i��Z���#�%�3T3,՚b��2�Q}�f���StsM[�����A1�6QYŌ=/
7[�l9{.&� �RK˼{�ɔZX���35P��1��l�\u>ۊ�!�R����@&7V��ͽن��q!�z3iʁan�[ Ɇ�S�Xv��� h����o� ��.`��D���L��T���h|��XF��R�Q�{,L�v��i�C����v���Xn��2n��r���ʼ��#ah+p��H3.jGrۃEK�t�$�bM�Ee
R��f�eh�e��W-l���q�׭�������{���[G�wLE��̽�����L���n�]Y�06�A�kZ�uf'Zȧ� $g	2���o0ی[z ͣ6�f�F����L80�Q@�UL^&�̏E�aȉ�l���h	h��q�t��[�vd%�A&edYna�ۂ^U�d�`6rܬ�+m��q2��L���0���`'��*��V,Fhڸb�j�Ȭ�82�,�28�v+�O�n�j���F��ON8�a�62fe�
��.�@cLU��It�-����02tm�9k�[t�m�XX���x�I�"�il'k;A��:���-e8/��q"�y^��[
r�0^�i�)��Tu��CE�,+˒�N�gT{j��F�2W5m����&_l謈�c�A�������\Dᷧ��X㷿0|�KSy�
�v�����J �C٣`��嶟t�w/$K�Wu8^@����u��|�I8���l��ۑ=�k(F)��6ΗZr����-Zg�e-��d��tV��Qy�[7�k�K1�}t)�6��23�e2��yfV;Jv�t�� c�&Gu8v�������S�M`�y����)�Wrċ*�E�݀�t`�ћ�]jz�+Q �}vi��$�5�;E+W�4��)�PW;�].H�K��衮��ֹ������۫r��2����T0��oY�O��	b'"y�6���+���t�(�>��n�*Ս�k��;.d=s#����܆����De��ثg�9�wn�xYiK[ѓ�P�� ��.n����#���{(��h�%ܫ[RҐJ�1��q���}����H)k 9�|𼃱u���v�+�7&�󻙰uz9�!��:ɶ��n��Z����sb�0�eI�Ӥ�$��b���^�]ȕ���n�\.�C��U�8n[�+��̍�nZX�s彆�m�GW�+V�"tcO������l�<3P�EO��)�KR���ķ�ՂQ	'Yv��C|��7�P-�39%o �h���P���R�۵�"��:h�LӇ#��,IDr>��u��7��w�K69��F?���(N֖C�!Y�����:Mt1�\�m|��}�gy�
y�e���.C`i1��w����8�i9(�TXS%�̂�B�Hs{E>��ӓvX����k�.�q'`˅G����
eEXYb_*t���W@v5W�E�43�Z�O*M��������>W&K���7�����6�n"m�����i���b>v�|a/:Qxٴ����nF�m-jʸ8_t`�U��9���`��3�����ޖþ�%�����;јj��&˥j6��Z�V
��9�ʛ�6!][�% s7�i댷�ki�yc�B#n�0�7�-Z�>ײWa��O�6�Z2�cr'��V�X���;>��u{��08�6�XJӛN�N��L���gNC��6�p��vm�[�,EW8���	�._�ТA*h��sxR��L.�)f[�"�_f>	q�))��</[U��Q��@Q�Q�Dl�"����twdΛw7 �n�=����8�6��Ы�e>�]�gRDWWs�l��hǑt�S�yz`� _wr���w[d'�������I�^����Qt"�B�K�|;`�w3/+���Y�iv>o�
�;4v����yR�K��T����K�g7YIfr�]J��k��V촂�4�l��Vsʘ%�)��J�����RR��O����¤y���a�S�Փ[��*&�mf7܅ �C�}P,�]&�u���);�Y�q��0�_k�{u�7���U���9��*v������uw)���v�+��3���j똬so:�X��,�X�oBࡻ<�=nWƺ�S��!95Yuaf����z���&s�7��g"廎�P��اM���4��|��u����3�Ylpz�����澭;8+�LLi�[rt��|;K�VR?e����0�b<�J)GU����-G=�u�q�`b���R+"����q�场�bs]�mu���$�b����-ֽ�n٣��*���Pۧ٫$�w,B1�T�L�P?L n��v+��e�Aˏ��3�&Gٹ���l`�]a��gwylT<Ѩ={.�]+mߓ�z�{ϸۊ����Wcv�=��:����6+i_T����sD�J8��.�e��uvq�'�)�i8�A��k���)E�K�SpԬ��X�*��]���aKj��z*�܁����U[|74����9M��ʅαQ�T7TI�2VV\�����w�5�T�G�,X6ɮ���`��!m���j�|�9�!wy��.�sݟp[�z���┼{�Vm<��]�$7��p�N�g*��c')�`5:�:a��k�)�!��{�8���Vk�N]���N! ����f��|� ��5�.�
#�3 *����i��@&\�-c����#�l(�%.t֊,�y��E��g��i�����$�H�why��];(wp՘�Feß3aA���jn����k&�u�]���H��(iⰙҳ2�ЂĶ�s�L�]*d�wv3��J%���`yg��f�)jǯ�*oVu�����y�.�Q�2�3v°T�ߟJ���G[s&TҮX��X[E���{��{\�CV���˻KvK�U2�7���Qf�%wu�}��u6���B��9�]���5����EԳ&P�Mʚ:�Ǥ�s%D֊Z����؞I�|��f����t](���tt�DX����Zh��Q�8�v�c�;1ӳ��{�F��5$�EڽE��iP���`=�M��e����Q�} ���V�߷u%p��Z�nv� 	�`4��F<����S�c)�˵�/kj��\�ʼ�T�_���>��w�����G��^����ˏ sh��F
��eS��4�ڇ&����WI>i��y�H�N`|�О�Um��Z>{���s%���.ٗ��T�X���(�E>�-�<{��o��j���-�;=���U^�0� ɐU��c�q��<�:I{�"��ٖ�L�on���vGW�b�M�#�5�q���[Y�6;��b�j�n�ƱZ�N�a���*MQ�5_,�+�9Xx�W��׶Fwr���#�T�`$�:�fh�.Ad�j�ȷ�l8� ["�t�՗C�tV	�Y�¡�Z��Պ�̚�>�u�%K�Xؼ�Ȧ��[!*��.��؈geK�r{9f��w�m>�ӋI�R�i�wR�ڔV-%�ox��vCcKm�����˦�O{-�P$�*�k�r5��^eN���*Z�!/f]r3��|���G�5��Z��4��gS�-6,_c<��҇+��^Ɖ�@Z9�Z����3�����x5����e�`��V)+�L�����rT���r�h� ��n�͋\��1�]�D U�'���X]��`nJ�����a����n�	��pɎFOP8���&�A��X�c��sw�+q5��}w6�h��{��\0��fot���8V����[4��Q4e-uv�Jl�m��(WS�G|ypt�'on�+riS$ݡ�#f�6`��t�E:���P*�(���0�;]mk{ef���=KD�6da;��mm��l��s�NK�y�ҷ/y�Bc�X�Oe��l���{�w��Fu�ĺ�73v�쁁36cձ�Ւd���V0�Շ#D__;�F�vkqf��W	ܬ����N�q�%]X
gQ2p�p�.)`���2]T�!]��G
�0��$ �8t�Yj��(V
v#��p�&U���I4�� ����� �g,Y���Z�9�D�1J�\�����/AWө8Ok)��	�L��W7G%�K�o&�t�}Y�A�q��T������<���6a�f�s�"Qe=}�0cʤ1��ү)�_l��.���y�p�1��T������6�gHSzt�|�	ge+E��Y�/���۽մ�t�>�e�f�n�y9�}�H�<Ɩ�|�ԫ [w�UdйQz�
�OT��u^�`�?�27+��w�lA'~�P���8%�7z�	�z��6�n����*���jQ�I��/�hC+ݱ�����zk��=�ħ�+�c�]36�L�碬�f�*���4����)ܷ���F�jyx,�#s���Ea��ٝ���Z��:tu�+��Vx���A^T�2+�#�v��N�޻Q-��B��}�6��b�����	g]���HHj͉��cN���`t�d��VI��K_^�齜�:Q����o�[�غ��e�u�g���ű@SVA�`��~��b/^�v��d�'H&d7g��Ժq�U�F��Br�����F�=�
�+��d��ue���&�v@�E��!�t8�X�-se3R܊���^ur���w�f\������;�H��o�Y��Ѯy���ݳ��t�5�*k����H.�w\���;�@�y�I�J[ڎ�p�E+��ɓ$���RG`/A]��٬����ƣ�k�B��ec,�D8���G���fQ+�iv2������Ybw/n3��S�|~�sSl�S]�yy�q�����N]��C>�E�d��:e$[�=�+^GۍGQ��J���4����v��,Y��p����R��]��z8�]t��5�k@�����c#z�|�q��\�n��9Ǽ腳+�6qމ��v� ���a�qS��B�����QN���l� ܶ�VpE��V>�y"g2(���GXbd��:��ͦ5�n����5b�Y�֭_O�,[�(��n�J���i�WV�O+}� b�5����Bl�vie� !�F�ۆ(M,Ri�4�����谽=����X�֣2��Nj����������\ʷ�����+B.�T��Bg�ݵ�t��w^F��ql��/5ʉ�[�����t0V�M��.�%�u�c,����O��Oyի�	�w!Ce�F�b���M1�=ue�vYJ���šw,Σ�6��(��ϻV�-�da;F�����H��/�X�Rv���k +�
��[�b'���y��5�z$��Z �ԅJvA[&T��)�1�u�u|����k�O�N:trm1y!=���N�m뛉�l��5:�+�`����r=	��5U���v���
ʂ��.{��^���I¨���N
4�=9���\��k�lxm����ۜ�V����la=j�[��v��YN���cDMME�"1\ɛ1%a�0]�❮[$r�K��їh�wi�Q1�{Z�N��e�l��ʔB&%E�.���˔��Җ�8�<l�2��]{:K=8���6}o)��>�;�=���.�Abq*�FL�
+����ڋ�*c-`��_n�]����S���;�ۢ�Y��#�l��l2�W��+\6���u)Y���S����l�\�S����5��b�����l�<!ާ�؝r$�a_k��u7]��1,��k���;��W�Y�3�)Z.�CXLM�,C�r�������3�PM��PT��JT�-���o�J��]]*�U����Μ��	��hŚ�Հ�ȡ��*+6�Kn��ɋ.�-�*=�9ۡӤ�L���Uq|v���Yz5@��[~��e�Ʀ�_/F�i���Ӡ�\�-hlE �I��\�ʹcL�|���/u\��A�t�"!8p����)�oP��n�2s�߲W]u3yr�t���j�Ŋ�K��PJ��]-p���*Wb�}V-��ϋ7K9��1DN�K��vS�*��Z��	Z����[�0��ys�j���z����^��R��=��2�x�lGpM]_Y��q��p��i:Wsc�E((�.�T�)����ky�͸���pM����V�S�����Y�6��(�Q���`/�\jd��@X*]�8�[���|��}�Glر ��J�7e�\�:͝(�j�t�X�q�Ʀ��{��Kdq�4����Z����pp�2w�14�j^AS�0��l���i�!y��@fF�A�M:�e�7{wA�V��ʜ�Ɖf.���H�+3����b�B
����WS����F
<�r��R����np���B��Er��Vg9ս �v��]h�o!�I�kæ!6�r�2�e�M�r��]
�u|�pCb��H�i����]]$W+��st;|���[��nV�]�N%҉�n��zu��f����9��ׄ�a��lڎ���{��/\���6V���Ec��g��SI��s8\��\����M�K6;y�#�ՠ���牮�.ļډp���4f�T���+kg6��5~�7��ᾟ+�Z����\Ӳ	�W9��v#͡Ƿ����r'��;|���U`���\�n�����{�{�@��3��n�*�>J��|1��L�]i�Nǫ�SN���f݋McXp� �Y�+f,�W�by�k,D�8�|�&l���%�Ts{���{F�B.*k�{&�rB�X�:���8�)1�'*��w��IkzWN4UC�����+.���y?)<咱���g,��kq]Ǧ�{Yy��&-P�sv�Gq�Y�t:��r��*��鯴�2Z�31M�LVs���1��T;��}��*�K��o�Q�-,��W;pVhX�X�>m�;���w��V�i>t6��e	�<��c�E�����o��$�³s�ݨ�@��U���|����+)�!��͹͕�� wSZS�ur1�d��e��r|�*̱�`y؄خ!j�W9 v�p��rl	�,�ܦ3/�%u�w��N�>b����])���>F�V��79��e�sf�� ��:V�'^\M��;�ޞ�Dϯ,]X$#�ѧ��	r�b����ך-fKl��6��ӅiWmrځ����"�%�Ʊ��Kw6ڍMvp��UxvD��r���[��Kz5�G˭�kF*]̥u#ʆ�[��WE-ԭj^Ù�{$�Υ���4�å�Ś�������=�8X�T�[	Y����/�mN�uE҈�vD8�9%�I��޹W�T�2����6�p��a��q�;�Y�/���&_oIRJ{\�hu�p�K���o��SzA��"D��B��+k%�Ϲ89f��ǅ�,��٨i�WC�p�g<����b*r��Ny�I}�Ef�ޝ6;<�I#W�h\�ERqeHb���&I��l;f
;&ȦTrd�tbU�;dr�s��v)?�U��BC�@�oZ�}��tk��u�����k�cV��ٽK�u�?m���Ɍʝ��]g4�Y���2E�s9s�r�-�F� �$�I���-�)YՌ�s���΃ʊ��8�^*}����tF[ʒ�������v�\�[j3���E��)ӎSJ��1�m�kp�Ǹ)���*��7�U����1��1�y�R�&��s����m� n�c�z����H�r<�g�.ŭ躅h��u�,o��o�[��VIq��v��w(���JP���˙�5��f�bq�g^�I�d��wB�i��.C�����ݬVH�1	���b����m|���P��ʟEuَW[7:H����W)��n��I䭩��|��ǭe޷igӛ�L�����m����� ��Lvӵ���VWRmvI �ʅ��t�x-���4�Ʃ(;��̐�b������<Zӹ|3�d�樜��L��[[Y��^��ے�n�����%P�y퇴Vi��H�[�k��:�Q�i������,���͑��	ӆ��ђ��v�5o��CO6sH+��Y%�qϕ��|��ܦ��� �7�#=O�䎬�vn��;Ʀy0qt�7�(�|+P�ÃX(n��nF�����Ez0�PV��/9�ޠ�\������]Y�Ҏ5�
��Sr��KR���a�W�f��.Ld5����N3�LRm�b �N��!��ٓ�Y�L���.	
�W�����6V��&#*�F�P}���}yv�J��̜��Fs�sn7/Y�q�)��ݘVn��t�����:;�Ct���A��n(�|�ee�ڊ.�P��M'���$Ƹ҈^>�k��8D%�<'`F�X|��jlT���8�G ��*=�Y.�4٫�vC��XǊ9��&�?s<�TKTR�㹤v�� q71��Xc��ۨ�r��z�,�;]`�r�V:/��G�'��;���%tz�e&9�y-^�K��ϋ�r�hMz�sj}2���]y�ip���:�=ů~t�%�q����(pv�ŧ��q����.����:��l�<+�� ��Jǔ/�gH)Ӽ]�g(�r�A��0�o������Z��ܘ;�AӂƁJ�V��E��K�s�:)@���	Hgw�i*}�����z�n�X�w�͕:De����y�k���y�d+�}:���J�C���텝{�J/r�����nKż2��s�L����5���.���⾗�Xs*>x
Ӏ��%�H�N��4��u�Q�dh��Vc���B�J��MS��ST���3�,t/Fb��z9�ڻ�J�C�+%E)7h��#��`x%�gl�=+N��2���K��X�C���Y<Y���}d Ĳ���.\�5�;WAHh�2�:ya����[��u�j�1º�u��tӍ|6��%���dJ[�LA��Ѫ9z�ۥ؂.���en��;�޴�D�Z�a�����1��S��Vj�R�E���%��\N���ǹB:�y�݆D�wtn�e)յ��ծ�Bnv�\�1�E���1���M�w����ڵ���Vn��Z��3;y� �!Ô��rP[s]u�ͬ�л��R!=w�U̙c���z����Tq�-d��s�Y�Is��kvbe����oc� �=�DYE��;�ewD�8�]S��0*ٝ��η(1k����N��{����Q���<��0���մ��&٥��xR[g8�xT��Y8J1���#���"�M����ږ����:@jJH�A����tc�w
������I�u���В��&VmL��K�Rt�^�OK�*[o�\��څa<�:˵�qH�j�V!H�OS��eq��QZ�R�2�z��Һ��΅dʈR�n�n����!�b����>�05�S��齑Cti���;���Ü��*�h�Az���PD��R�o�X/PA4%��3G����*�ȡ׳�əz4����컺ZE��J�7Zr�X�JT���!�Լ��,���c:���mc穂w�;��V�&�E�gf
�Zn�(��2�ThU�[������xc�j�/n�O*T5h6��N�h	l�A�����,���#i:biL�T�%e��t���V�,�5ˮ6򯪻]����wM{�X+�6(.Y�f©G�/�Gw�^^M�J�IR�n�yk玓X/���<�q���iU^��qŚ��[�a���v
�N[���1��VWd�m�Z�웬�R^���i�&E:�#��̮a7�Hb�`�:펊�;:��K�:�3,�v@u�7�/��23�6���c��i�Yv����:�\+�6r�fw��*#R���z:'#�[e�T����[:B�5$3��|���]���d�n�N��:j�ѐV�����0���jgf�� �� �:m�N$no)�h�X6(SXR4�;�t)RTu��
㑆v;�(��oh�7 �n�XЛ����k"�1+E��aK��>tR6�Ϛ�C���ɮ`h�}��w�YP%�Q�- ���$�k��{�P]3���;R��r�A-%��|��nL-ǋ)th
,���>�n��i8���n&(��Ƿ]`$7�:��Ɛ�or���1�����Ǔ��W%�!�4�-��qn[\�ܝ��U��[y���k��g8�+�.�����D��KhA20��!)��[�6��V>��Ƕ��s��cZnhK��ˣ�.᳅]�9I�7vQ놑@���j�.�+(M�+�2�2.��9i�qΉ΅��v��{sv��}���c$��w��+�j�{H��L�]ӣl�z�J��ŕ�	o���|��dHCJ��p��:親����:񅦜���Bv�5��%��I��b!YJ6ov�,�4`���wb�J�}�%e�n-���!J��כY��6V�|(7juł��0��E����x��+˙���n*ɍܼc8����s�P1weY�W0Nn�����m֍���c7hp2"d7�zh�)
<ˡy7)�ĺ�>�x��Ҷ���XT�fG�xZ;�Q�ޘ�[ܝ��f@�ֽՍ�,�m2z�.�h:2��}��`���Ar�@<t?�9Pʏ�STW)1Wo,�.l�����b��<ǲӮ��m�̭f�ؐU��<������*��SW��Uf�/�AB\��s;�c��Ţy�d��0���#yn�t��]��/�eD��R��g`�&���3I1��kl�y���@���$Z�f:�.W]�^�Ɏh��z��y�59f̏q�{��֜Y���`nr.m@%������A@�"d�p�I�qѝ�C���i���/�&V[&���n f.Ǔf��H��F�êc��7)b���I�t7jM����d�J�}��]8A�n�5���WhUԀ��ӫVt9��볍J|�����=�U�W�0�þ�:���!�ɫ��Ѝe�&�'�����r��룤>T�鄣���7+���%:�v%O�+U��[Y�&��Cx�CG�"�WK�=�v}��b���3�:�#�ը�"9�]��1���t�a�b�TS%����e�d��t�dR�/��N+3�*�M8'6e\��b*2���Qf]�|Ձ@Zo6��C�Q��x�SK'GgR�/�!0��e
�/��k�w�jE:���<��ʾN��z�C&�ϷuuN��Ǹ�Nk�jś�3�:��"1�n�^��t[��1���*��kuYMw����:R�@;Cxe`��ǵ����*�Y`����h���(V�X�vd�؅}�����9���n�gL���A̺��ע;@c�Jm�o�g�*j�)e����ok��R�V��ô�6��/j
�8�5���'��vYY+ }��v�*ȉ��ifkӢvլ���c�>�EѪ�	���;M��"qC�!�k�&�V�N���g9B�Sf���'j�y�يj�B9HT�4��{{�m�յ�-��-G�=���8�Gp��	JԠe������.۲xp�zT&�6Ӥl]Pn5S}���ѹ��N�DC{4�<�q�����^�v���7]���q����"w3�}EeCΧ������-�ލ:�~wf��Z������ƺ#DQ����.��f���75�.� �z#
V
�kTc�v�&�r�#�������:%�}�7v���f��ۢ\
�A�U��s��'$n����Y��]R����1R}�s��o5�"��pJ�I�K{�c_+��p�pLv;xl+3u5��Է�XBvsg���![z����+v;|��΋�^�$��s��:i;����x���M�WV���p���y������+�iʼ���ku�S!;'O�oe���'Pc/7+�H�v���+�T3YQ��h^���7�3�%f<i�qR���=�r��Z�k�n1ݕlf}��Y�o\�C�E�mJͶ򐺽�4�By,c3�����
-K
<���b�|@�!�A�h^[1��+J�P�]C���Բ���5�9՜\��P��w�3��ݮ�`l�$M��$kˬе�[W���wzֳ��.�f�ۃ���F�]�r�Z�RI�J����ٮ��t&.Vq��c�W�5u)H^na��q`���oU�Ia��J����Y�V���������y��P�Uzn������U7�fN�l�M�mcAPp���DӖ)!2�ꜥ�)_V��C�+c���q,�PX�e���%��+,4���:�SD}"B�hs:�T����J�'jx��.�p��b��im1�=�3����D޵S�SF���˔[�i�Er	����GZ��+��*n�ٶ2_<���!r��+d�yD�jL����*ͮ9��nM	p�lN�P�
X��Xh��vq7G,)��+�ͽgrA���U��</[v��)�q�������N�ɫ��S��"�sp<�gnŊ`0WvE��*��}&��	x���B�59���M� m���`ݧ@��r�Ub8�~��JT>"}�=teu�|T�s8e#���.��v�u,��YHi�1���g��f�VX�Y�Yt�	+�1k��	{�0�|vmF��e�B^��]5��^_s��`WI`K��4�,e뀪�*9Q��u���ٗ}5)n�ۯ�L��&�����H�`� OtޘJ@ԙ�s�n� ��"���z:`�����9�}p	����lӸ�$��}�4�!�@d6:���ME).a�����..�(m�\n�|&�ޘHv^k��*�v� R�Ƅ�k�f*ժA]�^A���Q�F�J�$V�]z(��*�t���.)3����^FM��,�J�m�P	^�h�C2�u��[��YJ¬�Ph���ɻ�SN@���K�b�Gh��2ڱ�N1D�iɆ�vy�����\�{�ؔ���$�)��#��B�v��K�5�q��E�	J 7i�!�3ol��7�r��I.����p��y)C7�R�2�eB���N�p�3���3����Ȋ�{787u��U@^#ݱN�v,k'(�;����v��L�+j���Q�;�Gk��*��hUj��Mb�N:�ۢ�D��o&ӭ���2���ƃ���m`�X��`3a��Ŏ�&[{�]Ѭ:��e����[9ͻ�je�S��Q�W�Oa�RoԾ���,�޺�W!3v'�~!�ti��4th�0�y/��7F���F�����r��r�׺�n����,�}O�ҏw�İT�U�ng*��zr��<M5�J2�mo[𬓒����.��j��V�sr�|���΢�`�k�)�a�w˲Uн�wR�7��҂��0�S;j�t���+ȑ�7V�qQ�K4������2Ģ��M��t|eji#�I��=�c��I�Wk��[�Va���!�ݔ%g��o���8 Ǳ��0��t��kt�o)�M����[��d^�\d"�>��hAd�Ԙ��1]�����r���j�"��f��e��ɬo+��*�&���ǩۥI�J"鰆���޸%�]�2�ӌ,Z���J�!<���|+sssE��9�nU�����f�g=�q.�7EI�jZ����{��\�� ���056ɢK��v9A���C���wk�<<�%]����xn�W�.k�SM�hr*�T(�Fx:��p��+^9��˱�гL�릕��OEk��u}`��u,C/���H���ԡУ{��c��	ݫ7��H]��4�<���^���w���x7��Q���.��;R��j��6 �4R�uL�҆L��=]�C���s_L*xA�ۣ.�3�g�jq��S�E��o[��r�P��Vǵŭ+��4���Ґ
�i�j̭Cc�; �G.��,YR�WY�IV�R[X+�͊V��)�mbul���N��3mb���ݔ����«�08�r�p��6#*�Cεf�ۛJ��4��N�(����6)���{5)S%�Rõ:�$�U���2b�`w)YM':�ԫ�Bh�)�5��G<5f�yg�� �	L��C]��U�oj�ʙS2V!�a��d�k\A"�>��,�i���Գl�6Otu!�R2���8��E=�I�L�7�x�Y< )G3,�����:s$ol��.}W|B#
�s����Iр��������zI�t���G.�90_w*�b6ܥBS�s�P��qp�Np�J��Ls�}h��:��g�Ǝ�8��75T�ӲH�e�^T�:ih\��ҙ�i3�U�K!<��..��o"t��7�,�*��Z�W@1!!v^R湗̨��\�䷀"�r�r5�m�ze.n�0C�4��.
���r�Q��RmV���v���ٸ�� 2�ua�تQ]g�\[�[����[zqmݎ&^�6z���6�3j
}K%��������U��/������bYw�c[y�^�uܜ5/�I�C'��B}�a������6�z���5���� !$ܗ�����y�o�ϖ�G��F�/�#�R��-fth�
-�vu��巜���WR$y��*�j)��ٝ�J����:�ʥC�t�+{�vuK׉oR�9p�7)�Ϋz����SYC%��lE'K�4͝C�_&Ӡf�FV%I�z�h��U���Ʒ��ㇷ���צP��'٩X�3���ts�/ነ���/(�|;�pr��=o�,e�e����5u��Y��ɘ�x̺��V�8)�9YϮ��2�eW��J��R���ˠ��)��yy��At����s�˧\h�V!*�t�fS�:U�ᳲ;1�|�e�]�	x����p�I����E�/��eH��Gʲ���1�[]�3��%�&��p���;�p�k�I٣(�J^�/S�zQ��������Y;6qZ�]�b�Ul���,S�2������u�Y�-�N;��Qկ^��.ar,��n�=�t'�o�Ԓ��yc2p=B��#��]�m�	,���a�f�*�����^Iz�M�jdl��]S��S�@c�h�!�+�wd��1�	ǁAV��ܥ�#�����_#���ؽh]؜9��;���-�޾���zL*��/m�� ��Rh�QΨsf`�� ��9
�A��*KZo(�p:2�EF�l�5�,,��' �tu+��C����4�W�'����Y6�j�+-�Ѻ���5c7��h�訾q�n=��� ���`�m��-��KiR�m+KJ��b+F%*TX��eUp�����Rմm)h�-��.Ze���Kh*�[ml�Vڅh*�Ym�"�bZ�F���ҥ���B� �(��ܶ�F�Jؕj�-n%qIR�b�nZ�+�A&�c[j���R���`֍jԩKA���ji��[eT��բ65��*�[KZ�kmR�*E��Ki*4��B�֠�-h)�����`��c�V�X�2�fR�e�,�m-.�-[K���QQ2�iGV�-F���Pkm��J��)V�%�%M[��J�UX�q�V��1eBʕ��EmY�DTa��(�����"�
)U(�R�"Q�Ak*#mb
���Ԫ[�k�b�QR�[j)[P�b�E�Z�*�U���5�M�%kQQAcm�B���1�Ɗ�3V��ʣZł�-cJ ���O�o5�34�<��q�+^�J2��7��=CK�(]�n��ܚ�ӭ�@]���_}+Ңؚp�1,s�u���c�z�s6���T.���������0���N�.�����W:2Y�S؛[�;Ld��T����΂��<?A�B��{,���c��7�}���F]5�^#)Lݘ!��F�Ox��=��ȸlp�}�l:�>�GTk´"׆��i߄k��t�ff�W[�=)��^�*�8��s�U�$�x����	��0Y��<MK�\<��Pp���H$�[<���K�(|���������wo!�lS�`�W;�泐��ݺ��&zuD��j-�5�����=B�N��t_0<+�ߦu�A���|��3)��4�{���S���4�5�y�#��Q���o���hu0z��e�[&�\�D�t&�u��;s5N;�g���g�v%2�7�S�Z�ϑ����`Y� [�v�q�oa�_::�i\䭩�C�0�$cZ�錛��Y��^��3����:M/��$뤸=u�F
�� ��hu����L�ϳ�pi�q�Pa���zޜ�8굇`�� h��{y�+��m#U���!���4[�q陸�o�Do��E�uAf�jG�1]�q��wy)�����'yU��G��7ݧpb��}����#8��v(��O�Αʶ�X�-�bu�����in,.�D1�ª���������k���.N�	(|�J�I���=9.���TǨ�����1�{ȫaO%��S<�糆=�54��͋3�W
}�pIt����{~n��i��a�E�����Lv�{�����%�Ğ��`EE%f�X���E�Y�9=6�X�aӴc��)93�n�0�^n��Bא��6C9�{�[q�L���O�����-s+�;����INK]i$)^O��22���[��8�l�+� ��"Su|�=��,Of�]	N�;7专�C�Ѯ/�Ewϟț�7�0(g�����lUd��E\bg
c�ǛSG�TÑ7�
9�Kh�\�o-�G&�+�+˅�<�#c�|�zMo'����t*�*�֊���5�kl !���{d�����=�&�����+x:޿l�YޱƺUg���b��-C U��h�^/D��b���0����]�rk��O]x:�pU��N���g�����\�'��;iMǻfa<فUS�/�Z��]�e���G}�{�e�g���Ρ5�֕�r�R�R���l�v��O�gfIS)T[�����G�CK�Pn(��	�)r+-��Up4h:ּcL�F�f�
R!��7�&���������%��^wS�:�Od������Ò�H�va��&:;y�k;�N,��d\�g)�^�
�v�2F��:.|�aj����ώTCC>N%%�#����e�3}o�-n4��6}\B=��+#U�Ck�b�[�M�?G�+}Aؚ��1ͳ�"1�֗Z�v���܌�Q,=�t�[����Q�)3����~PB5�^oS<����_������t�Aʋ����9��jw~u�_ͬ�uU�g�s
M@���Ȧ�#���{��BNx� ��Htb�CT�����ȅt�g�hF��>uF��3�K#�Ű�p��e-Ҕ'9C����T(����� XZ��2~\�E㷐g��
��˱k>���9]�嚕�$F{���rG��@i����}'Ȋ�=�Q*~ے,�a>����.WL&7�]{#!7�gd�@ ��HH�+�pW�G��;�N�t_����f���$��t1��0�!�k�����M4���3�|Q򱦖*5������nzԸ�g�A!�0��/<v��ށ�ɚ�_a��ֺD��$C�w���.��c%Fs���]��."b�MZ���\�'d��b���N�-\r���� �0�՛�qlY.F��n��S�Q��*�ǣ�B�gtk����Y0�)&!L������i���ݘE^�^5q�T�>���s}�B
���kb�H �z��2et�m�|/`t���򜂞eNJbUSa�'}�R�*���#s�E'��}�,'��n��?���p�l��၉mx2���F�r��E�ڄ�V���dsa��q�5��z��q�bx��]>x�B6c$�L.�8�f��õW^ujOx�� f �3�����ݦq�@�'�H��">T�1QI>�l�V��y��p��#ǀ�|t��]Ya��b9�u^�?���4�٨.�|�0�PK�⮁	1��=��V��PR.��߇R�Q�c��Ñ��0�.���׽{ƯM���+¤6��u�:�CV�����'���Y��ih�Q�S"'U�3geZ���0iіW�S�Ay(��{Ц2]�]`�/I���D���υs�THɻag�dn�S3P�q��}���T^�Ř%�2��_;�/��!��6��f�fLC.1�m}Ǘ��	�ZeXCz����zU��لڱ/�k6'����H����5t��
�1��c���x�u^|P�ۯ4��V��������cg��?]�6�ꂄ�`�Z�� ���x�WE��z��qb�#詩���*��n���2�I=��]��kc�ά=C�R��U�	���
x�PLa�E��*�	�> g<�#�F�gE8�\

���	�o^T�[��q ��m�o�>����4)��z����/QB��hB"�2u[�Ǟmv��5;G��\��8O��l!�S�Jή�;�����JD_����R��"��Tg9S��o�'X��h�^���O&>�|�V��ɨ�ζ��[�&���25�Y�6G�2BJ�X�2X�27	�c4����]�#�Z��tE(t���g���[��;G��0��r���cQ�����^v���-�� !���<�c��j�e�┾KGE�pn����\5E徱����y�"�n�5��8n��68V>�6�D��5�Z>>}��v�U��*hT�y�cJ���@`p�60�,�DrN,��̀��w���d�(���ۡ�sfX��+{'�7��iI˜�hD8q���sYS�ycb�sS��;�Y�Fv��:Д�w���]O(��s3�]��>�|%[W����t0p9�F����].s�������%�:�O���|+���*�˯>�)��h���*�W�0c�S]o�A�å�;U)�#�(N���p~�O}t4�ū���e�z���a�U�dXvzJg;�3���&�U��Xu;y�ƭR^oZD���5���"�x��N�5����m�wIs�~�>��ǉ�W�:+���B���ݔ#c�2u�k��Ff�+F u�s���"y_�0T�7<��t��ݭ$�t���g���r*�Lʃ��z�y.�N��փ�L��!1�s��W�eD�k>㠓�.G]t��^?w���4�������ePOh���K��OL9�zr�1�rP�L��L�Lu���]�\ų�h�B���wi��n����Ĺ�C���N��tS��Sj��-�Eʖ�]��C��?
۷�T˯�A L�f���S��3��ϱ��絻$��Ȣ/�)���SQz�V���?{M*���ZM*�<�7�3Z�	g��L��թP��Ҝ�(��wv;�A�\t�w�9^E_�r�} ���F,��Y��޸��Q���H���[�b0�R��D\k \�����U;ŝ_Ձ���Xl��6��K�KH�G�'������I�C!�s%ê��F �o�
t<,{�4]u���}\��;qiꝆ]Jݠ�]^T%�<��sE�.�xfpK�Ȉ�9�|��9b�(P��< `�0r\��z��D.��ی�%�OMoNs����Kr�C���-�ѣYڲ���%V1��;�QPع�*l�T�]�T���"��G�����^z�+�)���݂������q�YY�y�2z+F$�d���m����c��J��
�p���U�ׄӘ�y�c����2���5;���G�������{�e�nv�x{� �������t �dn�S2{]ÜB���W�BY��ߋ�y<8�WsM�����ݠ�j�9����{�ғU�R���� *:�	x�Fh�ʥR��\,be���(�$AYڧE��^�p_�#O�|Liv��"��r��T!�M֒�MeD󈑲@���ͻ��A���)�0�k�DD~ʫ%\�^N/HG�Lͥ�q*%P�u����Y<���Q,=�&�y�B0�@�.����n	���i��Ǡ@�K_m/�����x��f]��u�\6�B����#�Ȫںl��g:��?{K�Z��	��s.)�ZZf�!]9�Ȇ���C44΁Պ�g�9k�̅!	�]{(Z<]�b���
�s�@�=s����r/��7��]�QXf�,;:s3�0x`���_?�g`&v �ue����kK��K���l-h3�5�E0���%�ʲ���t7y�m�%���F콿lK�ov�R��!St�]�Ɍ�+{+Sw1TM���G�W1���M+����;Y�'vL��\�x�sz�A�;H��!v��y����#���!������@�����˘x�o�a�ʚz���D�A�	�d&�X���U@)���Ch
�<ҝ}=7Uvq8�N����%]Z<d"��Du���C�3r!Ү��-�T�<6�b��g%{�mm�7Q��f�6^(��tj6jrT��A4�d"�K����x(bu�"U���.���1f�٭)��n#Wi�3��|����YF<����g��
�3>����NDJbUSá����xyM#�y��ݘNCj��zM�,����I^l��ݕx�01-��)�xT��&��Y;kv��ކW�.�0��X!7A��Q�u������`����f<.�\��u����Klـ�V�]Eq���}Ԙy���43��S꤬Q���f��㒧u������ǕR�����WVX`tX�`�k>8��1�#fˡ�r�N���U�0*��3֣u�<~��^g���z,����5ׅ:�S����L*c7���#8d��52;��',���X�p�)��<��˦��q���;�]��XzDw]Y�sR�}h���=&�â�5���y�N��Bz��37X\�X��t�� �s�N�l����]Fh��
�PM�*7�3��*Y�^�q��vXt�vf�� ��k��Ÿ�����R럁�n�\`D�VV�1ǳᩉY��6�`�S	��+ve�8����T$wAs̳�<�{��7f��_���]4�6>�b̘[<�t�3P�C�t�6��Z�Ȥ{7y>�Y#�p���L�;U�y�_Q�������/�}��&=�d�X#�����0!�A��%蕞�����ҁd�� ؚ<��*�*@�9R]t�ݔ��w��ܑpw =��!���8n���z�r-�!Y\�"��ó�I좷��s;Soس��h����!p��D.4g�+x؍���`FLwͻ��v�J !F�]��'Y�G�p�,j	ˡ5Us�j����gʌ�֑�*u�X���_���×�,Q��u�J�\WHT����飢."�K�y���&����.q�c��)��nn"�,�Ԃ��xg]���u�sƅ��1 YU`�Ch{���ǉZk�Ցݐ�{nce'"᧲
�o
���b>� ���`��g�W��M=C����$5i�z�p�	�)��nj�o��af�/�K�%Ay�Ӳ����p���S�����L��r)2W2���=����8�Y0
n��0�ٜ݁�xH�s��4r�	����D�zc�2˭Ty�9�6�P�[S�3��OHr�Gx��Y<�aA��V����;[�$]4oteԎf!�=�~#~�c�c�ca�Z}��^��5����ԡ���}���b^П8��k�q0��M�֯⪡��IŖwp��F�$�Y����q�r-W�8>��&0l㋭���0�܍6�o���N��*u��N�x��g!�tl���ً-����{E�� �5��ã��� <*�*g\Z���k��:�V��o`���h��Kk���n��,��_`_����B���݂6<*����"��KN�0pY�.�,�һk^;S!ݙrkb�ѹ0��XB3�Ǉn�mk�P�^�밡��)��ZS������^��LB����}�V��"�� �a��d���'�n�;�q{�Orr�TP�������0�؞�s���)`c��\(&h�5`�*�qΛ|T�s��\�������w�93��%�P�km�S�S
+^�
�Z�n�Xp�<n�W�]}"3%��"�Ůvdλk>�cx9�n�~���P�/����/�	��`��mn�.��'h5*���at�wW<����N�x]�.���g>sv��0͈s�X`�r�Ҥ�ѹy���t[V�*j�/�7vȬ�s30SJ�.�;�,�8HF�u1/OVݵ6�Ū���J�n5��$Qג˙&lP���ʵ����:����p�'sZ.4͎wt�Mձ٩�ɏ|*�lcZ�\;R��*8n��7E�ڶf#(����ʄf�f��S�H����h�P��5*�IbF�����|[޻�I��Z�2��7�.?v�L�R�L���+rH���`���|D���ޣA� ���j�X����9̲��M��ii�o@A�0nE�%�m�8�]�v���^�+h��ڗ�ԣӊ3)���:+C��I�n�ubŎؓ��[N�rΘY�i!�2�gj�5��q;"��h}���J��zG�r�R��y���Xt���㻀"au&��htܛ"B]�V��\t��J���^Rٹ.J�Nҩ��w�؛�j��M�]��'i�)UǶ�5��n�̍�0�{m�ؼv�8r8�^��v�a!gl��dwa�_�w(��󺐫�cRѝ�M���wmc�9���0I`Rܤ%l�vC����qe�����7�Vv��%�i�U*���z��@��:��KWu��+c��`��v�@��{� ���f��9ѓr
��6y�o05��v��
��s*p�iO��X�ti��\��c1;z��:�4�m^;v_df��޵��|_Sʇ�e�.`�&w �@�8]�%K7sY$װ��V�2��n��]]M��w���ކ�0�m�����Pۂ?^��
�w�6 +l:G��W�ff�rwrW!����X.V��W�Fd���}2:�2�i8`�$�`�ym�wi�aC���7�c����R�Peqv�+��0��;�(,��g�9��0��#�׆��Jt������� �n5R�l��w��2�=ҫ����j���b��4A����wh3��n���2:=�|/�Sz
�	7��t�&�酣EQ�`1+�W4+��Y햚��:J���Ӵ:�I�ëC�Y�;��e�r�+lp���t�&SPi-��H0>p�.��ɴ�s�����G{@���i����G�%r��kxho{{�s�we�+��X���H��_7�wS/fl����>G��6�2J��]E��(���B�\�1$�Ln�3~���;o��.S}�z�Jb�� �em�\��vU�$��ڌn�F����7ʺ:�cNV��)_eq�V�z�)^t-��l|jf8��}��qO�{�v�	]���$�5�Ee�e�˵�D+5�ʕ�V��8m�Yu�B��ې�Rf�4.�:g�t�%�_"a*���<໥]&ID�6���9>y��Ch�ܛ�+THT��b�7$��@r��d
�:Y陼N��Q�.حR|Qi�3�l��(�
�q�sv��Z*	mTT�QQl�TUh�h��`c�Z�QkQcQ����JEX�����VT�(�X�,Q+Z�r��XԢ/��db�c(�#$���Z��m�m��1�j�j�M\ʈ����mc�cYQ-�Z#cZ�R�$E��+�(�
�1b�1
�SU�(�¥1���m-Ke������k#m�Z�J�SMm��\�*ŭ���l��j[lEJʆ�b��5
�*"�J����b�[�*Ti+Ej�[%�D[cF�`�(��Q`*��P�+b�jF�VZ�-[,`��ETR��V��R����ӂ��X���V�iV��,QU
Z.�X�*�m�A�s-�c��2 ��Z����
�DZ���b�-���ikF��Qb���*��UQ�j(��*+mPb���"5
*ź��R�[QQ[J**��d�J�#EV
[IR��/$P�L����7O2��7�0���N��C7mDEaB�j�7Eу���I��uuYPe�8�VY�W] ��	�vŤQS8�5n���{��u�,��?����1 �k��:�$�l�+:�ai��&&$Z�ݲo�M��y�LT��{I��i��'���,���T��wRq�g�b'֠O��Dμ���;��w�s��&&*N�fE'�W������d6�̖��<z�H,�~�`�'\bϘl��`)9��e?2k)
�k�~a��M�$��g����<����鏄���s=�RݿE/w%�=�	�Ɉ?P�w����Ld�oSL���I��m'P����_f ��
��9Cn�HVb�Y�8����*N'S���V�F^'����"!��ё"s+�,�eﬣ�J��	�&3�L{>�@�:���xs�����Xy��A���`o�f�I�11�&>w�'Sl+
�=}��m&Ш~g�Y��ɉ�1��]$\d�4��}d���0"~���A����=���R�eg��&�3=�z�V�w�q��q�=��%gR~q��s�OSĂ�0���l6��$���Ԋ(u1g}�gl�+4���������c���L�_`�B���E�S�Aߟ�����UPE��AO�ă�~a�i�g���D�'�3�J�n�P��&&*��i'�Y<?kz/��gY/�֤��<H,���5i>q�>gwj�R_�~�\�귯�Z�EO�~�p��O�#�:~6�I�b$��cOP��Ă�������1 ���/S�&!�3�Y�%�=C߬�N!YY/�wZ`):�N�5�:��B��O?j��ۯ���{����5�~@�یt9�4ͲT����g~�>a�`,߶x�&��K�'��3�c1�~�Ă�!�1��u�CiY�T�$�
�s5��RuL~I�u���*s�ߺ5�?Զ~�&;ޭ�ϼ>���
�*�⯬?Y8����J�^�|����&�>J'��C�6ϙ+o�k�&��ɤ�:�q'�_.01�I��2�g��Ag���:�a��c���o��޻���n�Q��k=~s3��13�b*}�s k�E��>K��+�LLd��d�>�;I�7۴���K�9���H>��<��+8�Y7��4�2i�~d�y����d��J�R|�z����=�������d�G�aƂ�v�'j�GD2�;���q���cq1��c�!�`i�wKn��t;6uݼ�:1�v_[�sS�̹�']�n�e��A�{6�E�-�8=rPE��9\�eq�Y+��|��9�Iz�9�t��ޭq�6�ﳙ�z���s��ӂ��y�wMj���4�^�dդӌY���I����G�tgY.XwX��Xbu'��{`c8�a��s}èx�P��sY�!����*E��&#	7�s�|��޻������gI�
�Y�p2��"�g��o)��0��{ԓ�6��i�����5'�~�T�O�x�9H(q����a�$�������ƞyw��^����=g�1 �KChT�!P�v�?Rb��̳HJ°��>~dĘ�M�:�O>La�y�!����O7�h��2T%��I�Vz�Y�Y�퓌Ğ�\�{����ww�:�����.�$�iğ���ԅf$��}���x�Y��C��z�$ݠ�(��>eq �Ȳ�̼x�o�LLC̤�}�&r��ә�i��/�o�_p�����[�)~xgƭ�)��������Vx�Xt�Y=M�̜q��~��I�+�&&w�Ę�}OӶM��8�e�&�=>�2�[I����%H(fS���~d�I������d������z�z�����������g~H,�~a���~�T6�P���i�!����M~�R/S���u�?&��%�y��Y<I��<;a�)
�\��L��)
��m�Hx���>�>#�ge~���Mörk�3�~Ǉ��8°:j�N'��z��}�ِ4Ρ�b��
��Y��s�O�i`y��|�I�*w(�'P�ǩ�3!��XT��4�<d�_!T|j�W�!��Rd�h.V���?_����{ϯg�x�~�C��&��%@ٮᡓ�Vi���2B�d��g��M$�?8��s��7��gRy3�km�LH.�9�u<a���<��H
,A���Ϋ��'��L�ro��ˎȬ�"9���gxͿ$�L����ܲgl7-�$~CrٟRx�$�>dڳ�J�ua��u����?d*N!_̛���
N!_��I�y�B��������nb�>���=N�|��H-]�#�z�m&8�9��=d���wCL�%����8���%���8�0����Ă�5N���P�n�9B�^�����:���^G��xϮc�L@��F���ј�h<�~��o�2����ûV��]B&[�����\
��@���\S�Sp������\�M���co����v�k<&V\ǥCH<+�@�:9�Y:����4���ܫ��m�w��J���5mg�w2�����wmg�fdt+��λ��{�@�fwo9��iY:�gp��%@����0Y�J���m4�L*�������=a����3ɔ����Ag3�i�g�K�1Xx�I����Q�����I�7�^�=B�d�'y���'�J�ۭj�2bLNr�C�*���g�D��_���z�3�%I���42c+<a�1'P�d��@Ĝg�!�)�5�!Y�~��ْo.���������K�|��s�LT����=a�1�?!�P1YP�}�4|���Nk2i�=I�Y13��Ag��3�xw�CĂ��xw����@���2b��K����c'�Oݛ��Ѻ�~x�q�t�({���1Lò�I�`)<f�]?�6��![�q�V�����LgY-��}�E�d��Ӝ�$��1�d�Ow�l�u�'�޲|� ����w�<O�qH?�/my����{� ��S��MO��S�����H�N&̰��Y�.Y��u
�n�d�m`,��8���q�R}/�3l�����m��ed���!S��aU�s�M$�u1��ߛ�)�z�^�(�G3�u���f!L{뼨z��Ă���Y�i�Cxya�¡R~u�)��C4f~d���t�'�̘�˼��RU�����O������x�̕��5����Z�s^k�{�{��>���T�d�+6�~��������j�Rq���syP�ԅge���g6r�g�11�<f�.�
�(��O�ă���3�c�'�{�5�%C\w��z֖P6����f"䂩��~ԛ���1'�sYN�b����h�:�������&�b�����X
N�41�&&r��˦VKl���I��d���ӎ����L�|=�/ѧfgfC�
��׋�P��O�C�N�����O�b{�wD�x�Y��܆'�|� |sXiYԕ���3��D5�*E�7;�u'�J�Y��p7�dĚO9M3L�-`/��0'���Z�rcG���mg����e|t�ed�;�|���eI�q'S��aU��0'S��6s��&��+>C�o��!�:��Kg�~f��qNwX���V;��H:���v�M�d�%���i���4�}�����%]O��"QZ";2�.��sf]m7M�7m�\�����X�o>��5�֣��c3�n��rӜ�X˶�sX��S�H4�cJ���f���۬�A��NB��wjFF��e����RᚲB
`��$,Mdm/���^��֞�0�1�&3��CHbJ���bLB�xj���O�L�%|��q42u���ZLI�/,�s_jU`)?3s��^$���ON�:���1�La�s!g�?EK��zy]nޢ�Oy�iu�g�Y{��P�A՛�f���L!�l�i ���S>��H/��̗��C�<�5�|Ɋ�3�}��8�:��߹���'P��ϵ&ة��"f#�y+�ϯ1N[CW��%���7���&&{d�ٓL�%�O���̩��[Mr�]�f2UCG���C���5HVq?0�3��6�Y���4���a���CJΤ��O?���%��1�ϰ�f���	�rϢ�k߽���'�R��9�I�,�&$���^ځ��4��T�����^d3l��v��ʆ���I����ݸ�'��1*z�7HV|�͈���f �T����<(j��>�r��s���q��=C9�!���+=�͡���'ﻁ�������/r����{�����=�[�sk��i��Yj4��xғ_S���܈�@#�l8=�>�U�bN,�� ��"+�x)��b,�3��;��b��zd�ɥ�4�_��u�"��jf����N��*u���'����lݫ�NCkop���n�uƀ������<.ڸB��U8�̉�V}#[���70���;����pJ3<���n�ݮ�f5��=�����.Aj�QRn��hי�8*17GR�ʰU	>�*�c�0�ݙru^���0��U�d#8sW�n�z�
��9M�:����S�ݑn�~�V�#�d�w�!J����̧�.���&��0�Sy���VJ���G�y�� jo�b䭢�6��6�5�](�h�rfw4�ե�|�qNGlk��$�2�_f�r��'
����Ę�4vk��ٙ��d���|���_W�&�G���H��XC�vd�*��za��}����jܝW�GJ�\0rR\ ���Y�=T���G�ǥOe�qT�t�,�\JB�����26'���9
q�kbFHAO;�rd����#�ň��,36FD�����1���/�NL쥮�
��`�>ۍK�Ϊ;;�%�Kt���n����y�@u
�$Y3�fUB�S��8 ϝ��9�v�CwPQPL�\�[1(��WA����4�6��/`��������e�����w>�@`���E����[���;Z5t��
c% �m�L�בS�ey�n�š�ێ�Z��)���*�m�k���y�2~�qzn; ���~pg�/�/�5�.o�qq?/��Ο��K�e.����Og9]�Q�/=C,���4��I�}���8�`P?6�d���U2N���W��*��ou����T�sr������7=+F�˂�y�F�:��p��Mv|�v
��3��i�I��㾵Ź׈���h����Z�z2w��Ϸ�K�Sr�}��;�!t7v�_r�E<ܓZ�ˣ�$���&{Ptm#X����p�Օ>���M���z]�m���*1k	�k�m^���+R��q��%>�����NJ!����e�W[�i��b���K^L@Ö�lRg-$qخ:����;49ՔhN*��qU���ƀ1�شg��>�ݦI@6���ү&��d�&L+� d5��{�< 1�|���.Ӌ�ܚ���T{�i{����+�7�=ϻ0�ͦ`	h58eL�(��'�}�R<ȹ]I����С3/��	T�|�3Xڳ0�ѓ������:#���A�Zh�q��.\�v��P���쨎#>�ԢVD�,�*,3�cϜ�dFoAy
t���z gL��-S΋i��'�c}A+m-����hE�.w���nFC���n�
�����0���ն��Ka�*c�'t0{c+�T��(࿶�n��a9�_��˵:�K9�ug��.f�$��-�T�}�����:I��|�͇P�ÙqO--3S���˅���W�YQ���D6�h8���x�̣�g�^!6��v,$3���=�ϙ���۪��&)-'tfſ���9�Gt{τ&��������$y8@i��Vk�Yɫ�Mx���D�]/QP���o�I�C~u]0�ߡ�^�M�L���H�5�B�����t]?)J�al��qO�Ж�y��:��4X7��T;!u�k*YkĘe����L��X��0װ��c��NjW���k^��X�m+��a�du[��&GP��oe���&�c���2�a���04H��51 �,�n��ŭ�~���L��4
6\�L�w��\Pdl���DO�	t1��.rV��*�f�U�Dw
>��e�P�<1�4a��W��5;�`rxFA4�d"�Kσ"�E�Iࡐ�Ds�8�������ڭ�r�(�&:���>�N�GX.����88e�7����B{�y*�E�ol�no�[� O��羶�u���Њ�]�~��!z�
�ϳ_���4�9���V%�(\�wjc>���W��`�sʘ��a����twnm4���v�R�ۮ4�ďeB��	QC>��8�~���J��!5�rއ]j��Z�tOY7�Y���u�Z7�)���Ț	 �Qu�����������H?Lfٜ)^�Yض���!��Q*�,���K�״2\�[:�ʎ�s	aHqn�n���Zvm�ZB�ZGz������l�b�T���OixS��q���C9��9���M����MO��3�~}rz�*��������<,3-VآC�]d³L[�-m�����ә����3pp�p������KF��v�:����� dr���3T�m]��oe����c��<[O(��C�7)�W*h� ���	�#U4�=�4c7�SK-o1LWR��J��r�p��;�Me���N7��� zcDή�^�>�>��Z����}	MCz���廧�d�Tc�<�H� �ay��D+��9;c�f�[��6�Iv��!��T�t|�#���|25���o�:�l��� 3Q�I.
Of<��ڌO��*�^���)�.0���t\f�I����r�:�SԴtN�[Rq1Ia͋\����]Ǟ^�,@�,	���nA`�d�\l��V�7����6o���q�X��d���}b��r����P�M�W4Es�����L]>U�܂)��F~넎9S��E���A�g��{�׼_i��9g�e�>`��eT��0ӪGG��z[#����#�9{�j6f���|inՌw* '��KڦE`��:"�<N�P�#֫G�sl׭<.v�J2d�jV�2W{$q��owc��M^P�f\�t�x8B��]����u�����
�Z�F%s�7C<ΞZe$�U7�p�w|rv�u��������D��^����l���Ҳ�b��n-�)�W����d�4�=j�*��IŖD7G��0�[խ��ĽDa�o�#�-Zӥ�5Ӱj�cN��U�ذgf��𧕽a;���sOL����Tqň�f�d���)�wu�+_���yϞZ;w�(ҁo���ʸym�M�<}��\���nvE�J	1ꦷ2�;���ڠZ�w�����U^3ˬ-���u����O�TkÕ��b?@�074ڙ��ka��N�C��u�}�1��޴�9�L�-��P�۷\2�$�*�}�<'�m\,�X�ν�����g)~�st���������*����[���R�='��^�E��f���n���չ��x�pG6H�9����T&�]E�6���˓��>�q����$�"x�\��
g4+����{�J8Y�bK��bza��}������'a_a��0S� �ƙ� 9�dꓭ�n ��!� p�o�����"��d��Þ����9�XsFv�M:y]9jQ��uQB���*@X2�o����?�����ڑ{d
�Є%c�{������n�J�v���z�\�WXh��6����@�^�B�S��|��+��!��rW�h���Bk�m1��m�W���-���	uǵ������a�����W��G��7�?SV�����ǥ����9-�*\4�9ߝ;@C��`6�f_�]�th���qH=�̽���n���d��v������&ʺ��������(�]���A�efӉn&�n��n��ː�v{l�]�'�?3�����~��w�05���//�Qu�n�U��;��Qԩ�al_���=�;z������N�8�8�'(��|��5s�W�"">�Ә�=̫6�߾O>3h����fC�b�̙S3�
�H�� >����Ӗ"��QD�/v��yכC.@�kf1�I�mOL�[`Pϡ�s%�K���5 ��;Q'v��qx�����j���?SB�=r��t��.����|�zMi�
f��I�ޭ���g���ᇢ�c2j��U�aTtk����	�B��o[;��S9�\[{rs�kj;����؂�u�6���a�����ɟ��2�V��. S�7M��0tt��a=qz�҆��Ƨ�X��'6;96p����I�qp^\̣��#�A��l�V��n��{;P�B��:�	4�|�3M����`ꩪ#W���4�X���+X|�u�<j1ۻ�,����q*%��%E�{|�g���^B��Me�|U�&h���"]�y�@.���&�f��㹡.w�Ȟv�g΢Xz2���o>+�ڰU%�o���t'u�r>��.�z�:ʀ*¸4��[^|�Wb����}~�φz�뻵Dp~���
���9�P\��vY����Ɓ���Mver�������9���u�����h��̐11�f�4�!���bBfwq���[X�qCu�����[���3)�wĽJ��!�٢(��ã2��m[��N�!�c�yC3���5S�����LY���Z�ᶤd�Y.��[�gR�����v�i�;_V\����fi�i�{X�c�j����<�I��K��{��K��4�M��p͝�=d��R7{D�cɧU�|���I��E�ym��*�SO�\��$^/��YV�,�{sWl���癪�rFLU�&�9��ʶ+h�"�E�(�]��eռc]iM�kn���ԩrB
�p���]��X�p>�d�ߣ�VfϮ�/c۔t��9��9O�� >��-D�E��Vӌ��3�"�Z�M�R�O���!F���7tIڝ)�[X��Xƀޏ]oR����r�E�{�68�!��Z���JL��ڕ&�um�%�RwV
�矵���B�Z�K��*΄y�N]�.=�mvY����.P�[�ev��4Y����PWy����!��M-���o�nY��V��E��~]�.�Z���"{G��d�&/_��6'=�d��5�R���p�Ǣ�Wv�B�]�P�TfƖ�ِqԎМ�{YK&8*d�X6o$v)�e��n �Ya��ھP'�m�7�hdi���rJ��ؔ�y��(������[����#�"����Υ���$�b*��v����.]��a�g9�C�E�aJ�;v]M��rL��j^%��f򂄑�X)T�ܷ�-�AǠ��Oq����$\n�0��*M.Օ/A��f����{�S�!`Ji2.Lɝ�2E�0.�]�X��N��Tbh8����(]�Ge�G�$m̙���%#�p��(Q��㝠V"Io,�bw�-O]e�[�l�F�`N�9��%gt�yB��A���������_WG�o/M�40��4�w+k�̳]���s#@-�WJ���r���j[u���t�6L����wôY5���$�gm.�Nf���7�v^�薻|�*.=��g�g��'����\5��S:��ļ�kP$��5��3r��V�:j�ͨ���N��v���F��Ֆ��k�}������4ss9����2�OX�P:U��7��-T\�g��e�2��33���V)�ʖ���9-�Z�b�*�F��1����䱙�YۜݾR�ssA%3�C��Ev�#8�Ӛդ1v��Y�-�u��P���x�(���3Df`�.t��P�A��uz��jN���>u�)S6rp���%]�;�9T��5�W�ԗ���m���%�	a�Z�oR��ckw�ޅi��T(W.&m^��َcĥ�􋔨ʍ�Rk��
�ZI�:g41`��'%[�m�r�����Q[B���߽���:-w6��U��!T4+\�i��&K7�AKWh]��2�O�� �  �E���KJ�P�*
�U%e�m�����j9j�(1�ت���kRҡm�b��EƊ�"�j�
���+1*1--j1QTdFҁZ��h�iZ�cDE���EV[b���6����b�*EF#mQEDZ���X6ҷ*��JĴ��,�Q�-�LJ+��"�lQV�EH� �X"�"+V�+EUU�ZQ����(�X�QEY��m+�\�(1�R�JFՅ�UZ�cVe���1QQ�Kn����c�b���PDZ�V�Z�"�b��AQEF*��[B��F
�MX\lEH�R�����-A����UD���R��H��X��DQ��DA��A*�B��71EPKj�E`�l�TTTUATݪ��
#UKm"V�*"� ��dƢ5�E\nYEDKj�2�MZ"+c1�U`�U+**(Ͷ(��*��Tƕ,TEDEҨ�TF#Ң)�]��,՗)F#eh)�W�Seئ)� M�o �!�$�����} ��R�.{p��L�7f�C%#�� �NV�w۶1��X��}��DD��%ܪ܈�7������̝��K�yfs0M�O�ft�$�f�V�5>>K����2���]��Q�ɱ�#�z[��(��x�M��W�d X[}�'tW�����e�ؾ2�Y����U���nԐ1�@��v��rG��C���M8���t{��xf�xv8�0��\f����6!�t�f}�u����UW$O�O�]�K�|��,o��31��߸Rc"xȎ�H㡍��9�Xe_L���!�O]l.�$��-YV��e@b�T7�od1jv09<#	��!b^EЄ��B�"oc��d�&B�w�[�]Bl82�z����O5dQc�g]�B�hUɐH��Y�n�����HG�}��	~�羶�z�L����xv���]y��.�za�`�N0�k��7/E���J��gڝ�,!�.�:��B��&Pc�D���\���b�-{�NMb`�P�]u֐H.�8�b$K�-+s������i�z����,Ҽ�y(��`Y��bT���1�R;�W銚��-��4�ҍu!u��Z�q4oy?={tS�&�g�𝳕^jb�*4Z�p۾�o�^��Ͻ�]�Xݱu,�C��4:j�9z:�	��]��X.�7Y�6
X�}o��5��c���JKHw4��ή8�&�d�,��9�_}��_S�⧹���o!|�tn�C5��6����k�'�g�5|CT��̽����A� �Ѽ#i,�%�XK�'����j�qpX��rTXr6ݦI�)��N��E��5��Rj���׮��e�UX(K z�c�\���KJ"y��8�wIe�5�J&vr�a���[�-o�S�B9T�H��h��Y�Ж`������z9Js� ��G�%0�JO:v��;����u��Q���!��6</1��!<����d�z��;iyNu�3�s"�ț}_Z�~��F��X��Y�:[���@�{�b*���G�K�WM9��pPU�E1Y�9��C�>�]+��0H�UO���z�r���҉�PX�ԫP���H�p�O��j���	�0fq�'a[��lHަ�6�);��Vi2��J�H�{h�}3<�W����H��-���ϳ�P}��_�Q(�W� �k�y�lzSe��ևO�[��Z��I���CWH��6��4�n�J��G׫�$�ix�n��9��}G6W^u�7cy��n:�j���x���:x�.�n��t�pc�]��[�ԹIv��.���+�NF���x3��岋f]ԣմ!��׫���7)�>v��+$*_�Ry���g3�1yFT�Sj�=�?ʯ����l�E�/D�����\AJ�a�s%��d�����2��(v�>�G���g�39޻���q��o��efd)�ed9�^۔�]̹����u3ꇹc��b��g=�k7���kL���)�D�I���]����aՖ*?�uغ��F�V?�6�iW��DP�\�h\����ƬT�˭W���z�^�u&g���~�My
I�sAy��4��k����FRڷ�;��$��i�W��>���a�9��S9�d9T��9���~�X΁e��R����3m>��\���^�w��Up��x+)��<� �w�t��,\^�sq�phrŎJo�!p?g��C����kKg��:+� �\��ളxB(�bW��{�o��v_ &z�]��Nt&�Qn�}���uF\�{�\#�S�\ �q@��vs�\�v�h����_8���(-WpTIv�o��^�>�LFE5nN����ߤ`���Z�^����g9��	�<&��M/��/蔅�\B+�:rvaN���3gHU���3xeb���P���& D��2���҈���]���%�

�z�[��v��V:qv ��N�7$j�:�댧�\���|MM�Ҷ�`������]��^^4m�d�H1l�1wI�'�!EN���W��e��d�k�O�2c��=t5~�>�#�7ջ�)�Y�8�z�?��
�`��}]�)��ӓ;)k�FV��{%8j�t�Ts�ze�׈X�m�;�0�n� �5�Hz+څp��(4�w\�^�G�vVh����)�N�z�Ct�ˍ0
�Ai4�O8ͳZ�N\f�[3�Q�ѻ���&v\�)�N��F��}3�^EX���G�BqN��K�|��,��*Ë�^#�9�EM�P�mWHJiL�I�ɖ�ԋ��*���w��n6�'�m>hl��k�	^��@�Lu�&����Wo&��̗�K��I	�4��@��p������}\��ɜPSX󦦏�mv9����f�-����o���)���I�µI�o��ˠ����e3�i�5Pj�]Pu�k��z��u1)y�s����r�6��EҴ���`fpڹB�s���C���Żu�#��E�NU�n��5��C�4��b�ގ}<�q��3,�pg"�:CT��"��Mّ�I�Y�p]ϘM�C��z�z{w*�6'�u-�	��u�$�{���[���ky�	�7�Ζ �y�8��8vX4hr��A6I.����׶�y��"7�j-K�$LŝTk%�e����wm�m&��;��B��d\]��*�KQ�Gpsc�	1�&��N�-*�I�����b��>ɼZ	EϾY�v�MA�������n�%�k�-�3�]fr#Mm���3���ren����x�l�+.7"���ʈh`�q+$9`$���K�2#{ ��/�c��t�{b�P�,�s�G^0 �Ҡ��uL�U4!k���v�1��a�L,;\؅�}�o,�x��H���W�d.�`�ⴐw
�>����~�S��
������B}bvB��w�g�bJL���(k�5�������鹄�K!������rm�}�0˵�)��Q��u)T��y5.ѝ����E<��=�=-��!�׎6���s$��dO�M�tKꥋv�z�P�p��gS7��t��m�;��$��|��'�N��g�����s��S��&�Pg�=[!ĆB��(L2.!q���v�`l�a|�dbo�0.y���&�lot��9M*���U�D�4�E�gw�&2'���H㡍��,`53T�n�!�g��;�[:���H�j��Mw��_.U���>M\���t�#Ώ��5�4��q�7q��:� e_n���J����Y\���ʍl�7�3%3�:�
MaWe��~v$/NQ֞QE��)@�c�Dt������	�Mc��]����zp�����h��^��n!l�X��sb�JH�e��&٭����
#m�E�K�霡���Ϣ#ﾈ�k���f�0�J�9���ֺ���5�g:F��O-Q��3��j��^\�΢�c��E�_���)�x}J;�;�7j��_L',���v����_��tK�g
Q��^��Gqd�c��ON�Xs�]����X��>r�WyS��B�'(X�N'gltYXL�e2oRk��Z�# ]F�l�A�lg��q�ĉ|�V�]Eq�L�&��T�߳��oե	�!�d��>�TE��hi^-3,��n�����s�u.�ݸ��42҅
��{���/:OD��f����_=C3��K���#a�y�Z�i��t�5������J-��pJ+],����u�}5AJ�Ɲ�W�H��Zx"|+>��q�҇��3Q|��=ެZvΗ'�`��\>�ja0��n̴����"f:�|��r^�؈n	��H�X��ۮH�	tZ�̘;<�t�35w>}b_cy��+���yF��0�y�-��d�c��N&е�O`��S�ڷ2)����B�oC@᫩�N���g�,��v	oW7O��wt�.�����{7�wH+.G���y��lN��<=Avmֳ��^&�~�ڞ��@�k�P*�锠jc��[G��cm��˄��/i�:��}��8��h�O��q���v�\�ԖK�GJۺ�l}�;�{�VF�S�t1%~�菣�+��*k{�3'+�A�Ԛ�1q0�7���Dm��+0H�UO���z�LwE;���������(SI)z��� 9|;�x�[t.�c�v�lF�Hަ������6��Za�꘶�n��erͱ'�4�����D���^B�:�i��i^(�wf���*=Z���@��y��R�|�:�r;t��
a�4y��] � >A�m|�^��v��.Z#�RJ�a�s%�X�ٔ��|B�$T��,8��;�V�h�n9�#�ڸ>ʃ=]�`���s�����̹���/gSꇹ:O>uH��9qOs����汼�� >8Y/"����CC�4�)qۨ�j{.�F�˗K~��t�����.��1Z�鬞𮺖he99��|�S�ߎZ �i0z��UT>���	�p�Ƨ&�!�����83Ie^��}K�q����M1\=�(9�jY�03tڙ���C�wڋ�>����ɇJ������ְ�۷\3�F����{OʆQ��<+}s�u/x^fd&�7��}%�݊����O�Q�ǻ�Jj�g����Б=a�1ҍ���>�kI�-�����ν;����^�/��)Y7I�$h�@Ý�aUs!ݳ�V�]L馆��~�U����:�1�;k�G��G�P�wg�kI5"g��t�Ȥ���^]Ʈ^�/z�}yP��87d^��:aN����:�Og�v1�v��]5�ʅ<F^���7r�2'[�7��G�߅uכ��g���}-��V�����t�gr(+�硒P��!W�cHq�Hb�,�[%��0��}����9⯰�Y׹�a&�l�c0�f���A��:�3RM�Ⱥ�!�|r�!q)�E[�b�ϡ�+�u��h�;��|�S�T�wK�����Y������"xB(����x�����xA�jڜR�VV���㻨8n��X�n)�)��7A(���@yP5�Hd�E�P��uuzZ�cAkTR{�twJ��ϲ!��絻$��@c�Jf%-��"���b�TLv=	��.*�ֿ��E���I�S���1��`\6�s�"� P�c����������zR�U�{c,2:ɿ��3Q�jvd74�)���|��y��EVt���9裣��I{�~����ۊx�bx�'1"2}�&���I�Cw2Y3je�叭P2�Z��+8�ɩf�	S]9!R<P;�K��;�=��Ɏ_�o�y<J:�i�!SL�Y���a�SY�e��B�O��ls�5��i�T�݂�Y�`\ݶ�
�SW!��\�w"����$��R��B=
^��Kp\}�='�0-g��X�M{�����UW�Wӌ�E9�^���Q�
�Tj�Jb�\介��덵����囐�wdE[��ds��R�Nr�)���qƔMvC��^�B�i�5���A��C�۳�\��b��W9vyə��G��YX���ʕ��k�g���p0뤵��+{�w
�W�*4�IKc����4{*T��ff\v��8�1��ΡAus�ơ��s.�0��>E���Xtp�����)�)�8�Pf@d�5fN�bM:���1���6��d5�g#I�+�o1���N�L����� ��p��Wh:�J�r��J�����+ 2#z3��kKr7)]hJ;�iu��="�x]^�M"|<�	h릗���_\Ћ�s��s� ��a����3w�͵̝�r(�.�ώ|�4��@�./����U�\Q�u�oϖWb��_u�*�Vu�x5��U�\�ѕnw]3�p��-�M�Q|z|���K!������W&�_׼����ɥ��(��uMN|����5�Ѝf������ݻ�g(1q�q�
&Y���H%�����6.x�/����^G��q�C��&�}&6<��:*O�[s�%��+�:�Ҩ9:G\�2�Kd�#��;|-%v�;;<^�i�oG�2�qX{��:yg�G=+�^������mj��%f�Gbq܊nI��"��]�\SZ����{��:fͼ�oK����d�/�:����A�U�����R@ϼ�Y��g!"�m���+R^��O q�P����pi�ϑо��v�؇U��uײ17�d�*�d]?lb�K{��(�$M����&��`�dE�gzBaO�t7Pf�łc;cq�R�kpa�]�;@/�/�o��#���
U=uB<r�Y�j@��b[���Fjک���K�@J�;dF��]�CSG�u1�2��}���ک�/��o��f@=����H�ji�ng�s��eL&%�n��������~zM�>uvx��ܼ���my���Դ�����j��f�	�xT��*��1�U�yS�]�+��L���'��:)S�1���^�C>Q�9��LwY�*D�ҷ0�ֲ�?ݦa��P����n�RJ��y�c�40t��>�TE��!g���6Wd7g�g	ڸ��VE��ԩ8�j���d��g1�[�������	}^g��z,���:�W�*��~74�����v�]C�fg0�+)B�w&�[z�T�]�GM��*�s�V�-�r>��^
Y�坠R��42��U��P�볋�4��^7Z�w�d�f�o��|TCU�-Ȩ��Pj�tL+=�e��
���|��c�9�[�s�WgKl��ܨ���KX�t��^]��IV���3��"�9۹z>��ĝ��'��G�ѧ<뫺��|g-љ���h����qgeΝ��e��|!ɡ]O��^z*�����݄29���G먒�R���;z��Ǆ�R2s�^���2��r���n��z��X%	N�G[Rm�ʋbn�^J�q�!N�\·��Y$����e�-�s8Q���F,��M7:�Ϗ!���j]�9������;��\�PU�Id�\�+)��P����i�H�wa+R�����ל�����ި�U��}��6��;��>���
�b�o(�T݋~(U��S����̶�|�:�s�ͮ�sYw�j��s� ����涕�[F�&ڏ(s۶����@f���/��w7�ء��̜�e��O�.��9e���'�H�Ǡ���k"F�����Gf3�m��#Fb͈*#���#��hx���X;���m�M�Xk�%������RK��{5���M��<�N����U�4�h�[n��<���u�:�^S����[ț�����e*鴞����m�n�=f��ŜN�Wڲ�|U�x.�1x� {,t�#�Jx�dý/�F���l>�g��ʨ��XW�A͆r٘���s���KT�9U�~o�7�2�����q�Vr�RK(m��g���ѥ*�U�[��tNRc�M���ŕ7��6:���.�{ư\���n�̗pn^o@L6:I�EY���-�u�qGx/*|;�v3t����T�1���� d��JR�Aܔ�e��uY�+]**}��`�i��ᑷ�f(R�oD:R�2ٸ/��j�Y��T��\�c��$�s#t�)�$��e����Б��\�i+��B���$9m�3Y+�5��@b�)N�)��
�э�,ci��'�c����$�wCZ��2�P�lg��=zV�6�Q�A�7���)�U��n�5����=�%.��wy�
���Mr)��<Vr���b :iD��u\Y��l��>�	��(ulw����g1t�!���=\��NE��8����o"�[%�2��Y�v6P��hVHa�ɭ\����	�W�����EL�۔���ĭ�R�䬮s:�Y(�`��2�|��#{�pɍq���o5m�tV~1�Sʔw����|y��o��_�Qtw�ŭ�r_���i��:j�2�vL�n���y6K��I�uæ����q��)� ޽.����%������ˠ�E�ڂ��o�.fk�� lq�Z=�P��[zdd�����w�jC�u�w��߁b3�V(��D�lUAil`�"-�E�mR����ZV4���5�0�J�*��U|̈�(���Z�L�\��R�TE�A��
�hUEb"�]5�1QUq(�UDUDm���"�3�Ee����,���%�DQT�TUKb+XXm��Pb""(�,Q��`b�b1�(�P"V�iQ�6�(m�D2�X��2�[H���ecT[J(��X�&%30�EY���Q��X�$UQUQ���R"0UH�1���j�(��ƥ�b�"�+mU�5��*"�F �UR�PPdZج�U�%�XŭR�X*�H(�0b�ؠ�iWz���Q*���QD`���-��%V,A���AJ���(�]	AX�&4REV1�(��,���Ҭ�mA�Z(��1EF*�QUkQX*�,����fm�{��ϊ�7�0/.���<S�ԝ�p49u��[��ÔL�����/K�ɯm+ϯ#��F��(;��?�U�}��8���^��\6G�Zal]��󐎛�����x�ʰP��XO������Yl���o����C�"�w��Ϯ�\2���`ӣ,���H�r������b�S�����Fu�El�����U^`�Ë2aG7{/�B�q�K�o>|2�W�A-�%���j�x�>�n��z�@�քk����Ȧ2&�W֩[Ѱ�#�X��Y�:~o3�*o�������=��;D%z� 7S�F �r�
uB���;y(���Eg$d*�rxl7B`�64��D���w�E��m��f�vb�#L$��|/�{�
��������qI�>�rdn-lR�|g�k88�U)�{Ζߛ�A��/�"��D*Fz'{�ׯ��\��$ra,-�c��_����.v!�X؉��_�J��Y�[d�����W���íz ��v��V��Os+0ZO��ϙX%�C��ۻ\.wί@�N�zvXh\8�l�$���9�l]EcpѶ����]�lA��ݐ�{nJj�F�3.m�s<Ī�[C�>�a����^��]V���j���L˲G+��َ���x���t�-����ѺV:���VC�V<���y��V���k�^Tx��z�mM�'aU�b~p�*��
���M6��J��V� ��H��RxZKV�G8��+n�2�:-�SC�=�v`E�����{���P�q\�#����v┿O�q!�Lc�*pҼ\v�mI��;�=�~#>�r�9c�1'���>SL�_f�AmTtk´*-p�����:�}���=���,�D)Um�����;��n��c��j������Ζ	��0Y�<MK5��b���3��(|Nd\z�<����:���fU���tl�9��Z��n�x�{��m,9ƀ���{O�����+�n�jٍl�ֺg��J�3Pua� �����}�'�g#���	d
�'�R̡:5��UJx&�u�<f1�5���kd�˟��WQn�}���y(<6W<���-��� �o e9�cb�6	�dW+�G�݄5���{�v�l�×��!1�s�B��|�{�fxpR��G�nZ����+ ,%�Գp�ꐇ9*)��Ec#Z�ǘ��wKT]�L��9�B�G������<w�� @�'�T"��}ܾ�n���,�6����Zc��"1>!�W�nT��h�����;�0��CL	�7�R!ppf��}�l#g)u �=�*c�[�a�8R�v���Z��b�X�nQ�m�K��g��ORx�IϷ���j�cEc��gvts!����*�u�oY|�D�3�5���gGOGhFqg�0Kvr�j�Y�tf�Z�(KJ̮$y�ɽr>������V�߫ꯪ���8'���g)�G3jL�j�s����$|�(�}��JDĥq5�Efu&�Qg.M��)�|�w��#��MBE������;��#>b6X۾�x�+� ���˹��O<5�Pߒ :Tի(���s�7�*n; ��n����������w�����-��iY��V:���BH�V�M�r��M"2}�gɫ�8�`P���;���F�q���p��CJ����y��^Ud�QW�N�.ǅ�6���6�c�ި\/�nBq�a:z�[�Q�眖�ؼ�*��=�]��v#Ш^�Pj�]Pp�Bĭ}xMc*�Ή��=�6[�D]͸������J�ڟgz����g��c�KP�<N`?z�f�U}uPor�����^T�N�܈ӆfo��p�"�:F|ղ�4���3۷����!2{:��Η��ų�����b�=�5<	wW�7;�c����n�%�k�l�L8����V-�~�Z^ya��ȯ}��/��W�z��[�CTCC>N%d�,J��cϜ�����D<�7�#P���8pg��;�`�1�i<�#��w�y�o'hLZ�Wu8J��C颇J��t������`&a�\0CK���N���)�óo�f�f�@�&e�wS�������R������1��0qj �/;U2ren�+v��b�s��_U}�yN����[�V�ߦӼ���!^���(���u��G�#[�o��c|���,Cְh[���y�N�Ej�F`�(���r�������\�|+�����ve�TyASF��u2��������3M�~�eڝ�Q,u���W�}a���&:+��! URοA����Fs=3e��{�v�e�ِ!t�1ι�b��}+$ɕ�_r^xϕ)�#\Yѭ�=%�nf� �	j���E:wJ��Gt7jH��O\C�R�M�<f��ԕ�m�5w�c'���+��H\�P�D_ț��I�A����-��SX,e�F\���p���� ��j�gq��v�m��V-�خR=����ډ�زf����1Ƙ�=�N'Ҽo �|H��6R��pa��f����m6bޕh!�'���)^Z�H���G��R���Ք��XC�������i�.��T�w��=�d��Vfj�o�O\#��)�T�Ҙ�Umә��g�wU#c��cD"��a��xH������*��@�Wr^\�]e27�)���ژ[��Š���m�����M�:ӯ]��d�Y|9A+�t�5�L�(\����6[/\�s1u+�法����K�U��NyK���^��s.X���d��������v�!\�C�0z;)L#����Fg��s~gy�g��Z����j`��}�
�\V7��9��bT���d^�B�6c'bRc";�� =*s��\QN&:��w��ʂ[_��x��CC����*-�Y�i`�qY�{��0����'ڌ�F���8^TkI��FuU�讷�7xN��Qu�3ӪM�R�7j��0\�}��SL�#���|�4��rL������Yv�F�3��"��o9TN}:�����2�B�6�w�=)�b����>5č�T�';��vid,V��oq����_[i�B�**U6*�K�{�B����i�u��_L��8=�$��,;�Z�I�R֨}/���U��T���c^���J.nMC���QrO_����ȷ^���d��&�1��b�V;��w����濛cn��hJ���D��D�s �mq%0��1^+�"zv��.���yhð�/y�ܬ���gs���	T�s��k0�N�h�/�zp��Xyӣ�k��l�0��ty�N�M��3�c�n�ۙ�,2�t���w�U�7���[����g-%��S���n���;x `ݪ+��直���ς�Vh���)N䤆�����R�t�,���x��	���%3�ٲѾ�=:�-g�3/�+>caR!� ��'���i��H�y�UMN�q��� ��R��͋����0�D!�_'�EO-���܊�4I:ƅ�	���v��;ˑx�4'[n9��{٪�]�o���%]�UD�u�;����gx���ē�?jp��`M0孫� _d�2
Ww�\'�i�ˎrj���	:�?K����gz��{��l�y�!,��k�}��p�pт�:�{��Y��p��y|$�MK�-��S������~m�i�'lV�J�r�&Ųg-�>��S�ݔ&��9����|i�~����*�[�:b��7 ���SMdS:���zUg��w��n��-ʭ\�ɡ]V�����d�5ܘ\[툶�����5գ�����󡃴GXoR���n��P|#
	�Uܤ�u�ז`�eNj�ob2��{Uiz� l�y,S��)�};���k�ʜ��\��Zԣ��h݋�l��R kr�
��G�41����kYz����K�E:{s����e��;Y���W�}�{�E�t^�2��z*��Pf�@K�#<��>��&]��^䌵P�����Ar��E7Z^M�]3�@��P���#��->Ȟ�!�:�vcRSӖ[R���]�����K�2�䙨���9i�J�Q�4��*��z085�Jֹ|�鷬m�N�ɹU���bR�Uʄ��u�@�z�i���Ui��s'4��������sl!*���S��3j�%�e��^�P-GK�]2�"j�q���X�2����x���@�.UU�{�zc�`z��ء�����9k~�l��sJ��Zy��T�H�4��o�\H.���Wi�gĮ�E��Շ��eֻۡw��d����H��DK��bv �5���x��؍�γ�q=)�gP��"Wb�k7��C�x��Nz�o'�|�e��Lb;���{�I3��i���o�ՙlh�1�y^Hr��w�c����GYe[�G�g^Fp(�rŕ����d�@�6��Jr[);��YY���Wq�`ͮ�@W��G93�xk���1����sd.��������<���eHV�^����+��}�Yśй��w)M�J�����]OZݻ�9�.4����#�	2��xnr4���d����r�3gt�?n2�S�ƙk`���۱sw,���MI�z��gx�׋j���5(����Q�5.�3��"pn�7��Ln�θmu��+�'l<����u�j9�3����o��ƁPpc�(� �i�.�od5���뾙�/>��K;j\^�Zp�'_#oZ�ʰT��V�ɦr�e=�W}3�@��U�@��ԩdLwm���q[W�^l��>9�G���2��>�����*��&�T.�5F�c7�-U�@�I�oJ��K}��>�K�	�|�4Y��H���n*^RA�4�	�IE$<��瞪�Um��3}�ަC�������� ��14�X��AJ8rJ�>"r���}1?$�nW<�!�q���Yo6:�v��z����m�RR՝Q�av�u|���#�i��X��"x����,�n�O�?z�2iۮQ��_��:�E��"�d�Z �N������SvR��K�k47�z�:s:Χ�&��Z�%��m+��^�V���s�ųMZ���#��#I�h�c����Kc��.nJW�	�r�]�����H���.O:���M-ڱ��)K�5��Cb��/ Uo�UoH��*�<ѩ�r�Y\���bQ�.3�����͋�I9��jr6#�	���'\�����sF&Y��d�w�䕮#l��嫫Bʄ͸�����v&�\�8��e�WJݽ9!�@�'9\Rݸ6�����:�����hvB}mB��W���Wt�^�p�v1���u��-����m��������E��	B�O�_q���X���xe������O�\VV�����
+㬹)���ǈ������-�R�s���t��6f�75�9������"�� �)<��M����4�9H�c|���Y����V�ҭ��_i1��f������G��������K{��d7���z&}X��沈���.�}�v�yI�g4];�剝�4TN�@U�%��gC�u{)�f���/8�
@�����,�G��36�d�]{�G�n�Ee�,`��-�ݰ�yp%�Ϟ��ͦ2�r����՘����k����n>(2�A�����8�s��u]���9uR��Q_O7��[�����b�)����w,�8�m��V^���g��$�)9a�+]H'��R�c�}�wč�7wE8��f�Bd�)M;�r�!}�T\��=Η/��"��$��u�Y�jIЯ3D�9��x�'Λz��;BЕG�3���n%3�B<k��'-wM�n�N���O6�[�)	U�(�ρf�W9.���n&Y��sA��w�"�C�s�Qcb��PB]lL:5�
�]A.)q�M�ӽ����%7�Q]A�I��s�9]�I��Pą����j9��c�9_۹��]Y˭�5Bӄn9�:bcqH&���ƭ��z�9��S����'q\Sݽ�����x�vT��R/8jR���ܢ=T�@��e?h��&���WX���ލ��|6%CDЎ�a�b	�:7��+zZ�v��۰��2�ӽy���J!py[eU�^�3s�����Js���^����x���E��r��W%�����R�Jop)�e�|4[,�3�U,���Դ�a��ؗS�>��k���n��ǒp�)M9˨��M�$��U80�Q�i�/ �`d���Vm0�w�հ�<��y ��zd�u���J����������+	V[�,lJ)���\�G������%u3xa��5Sw+jQY�!�o�1�&�n����6��0��k�2FjA�W*�{�0��U�3~��*#�u;��K�����kt�pqyDSQ���2�V��^Y�2E[I��ǯ@�w��޺�Nn=qR�wz?��1;����ۺ��:�0�`�vd��E*�Y�Ԭ�CY[�2;<�����'n
����YnY_`鏙A�++i2E�s^�gR��us$� {�3��!�|�rr�tY�k/�⺈u��L��M�͒���z5}���Wt]�1G[]��-M�˰�v;��H�]�lK#4Ԥ�����,�,�3��I+v�g�æ��I#D�]p^�{�_���~AK�u6�(rkT�17t^i]!�֬K%K����T뷱��g������n���ؾ9hR��[����M�P���N�7G'��Α���`] ��+�c�/���Kq��K�2��Źs���{��Pc}W.��J�Amf�4�a��x�L��Y.s��[�a֚L�EԤ�uy��k6��B��n�MZ��+���Yɧ�A�iu�̹&���BD��P���X�@B�;���5�!Ư�u
��M���豃�NѲ��\�n��'j�b�lH����wO�vw�P����	`���V���V�<��]t�
����k�v��ΕKopG���������1�z�;5���T�1�fl�v8g	�L8���|��� �+t�}���fJ)
�8@-�-[ט��}1��b���o$WrN��ǚ�]p|�N�7yE��`y��,���N����]��3�«�o+�!����#������zf��[2���Y�t���F�cƤj`�g��o1ܥ��)\S'+%�C��rZ����g&�7g� ��*P�yw@1��vUl!X�ve"�eԮɢ�e�V#�TΦI��l�s �5�aѹ�x堻��z:`<�Ï'�1^��g^�28\.�4=�¤����<��E���551��O���v���T=�s;���MF \��t*��q1Ǯn��l���8��=�vJ�(3eѣMP(ܩ�8m5��uM�FSJ�j#`h�k��v�z&V�xZ�xv5��q��U�l����de��v�d�i��݋4�r�.�z:D�WW�H&Z��s@8�Y�;��f����!r����7����9��uk���R�os�w&j���y�luv��hL����S���1��j�@�jնĊ[(��Z%V����V(���c�D`8���F*��J����ELJƫ�U�5�b�\,�(�QUAm�%�-�уXX��DPKleJ�J�ҹj"��s%1�Q��U�[Zڢ�f9�UQ+DF#"ʅ\ˑDb��`��b�9h1E5B���kE�V�D��X�s1R�DADPQX��h�"�"0QX�h[b"����\�DQEcm"�#R����(�e��E1�+PU[h����i�*"2 �
�#��#�E�""�Vcb-J1A��UUDX�c����TAQX"*T��"�*��+H�ZR-����(�(��M:p��eUT�b0TUT���",V":e�*��)��1.��EV*,��eȨ�QQX2幉1�X�&[ (�9��L.�v���J7���<�q��Yx
C�>]
Ձc����U�ZN�.k s�g+Fzy�&]u
���꯫����~Sa���&�"WaN[����Y�9Nf��ulVV����Y��w��g�������/��>g�^�:r�a��v��fy�+s>Y����������Uy�󊃨͂�s��A����q���uڻ��4�rp����V'���zȞ��"u����b�k�UQ���#���Y��d$���'����H*�7j\�F��K{][�(�ʊ��;V���8�Jȉ�U�zT\����ǅ+#���zGo��a�_�O����zWc�o"&�R�������f)a�8��a���V���E%��qD��9�%�ft�c:��(���gz�̎2H��#q֙n��7T��ݙ"��.�Ns���+��2���!0N�N�tz�N��_�|gS�����ʓ�c��5Ͷ�6T�˶J�n6��X�'���η�u˨�Jn�k����8@#3��o+�R0o��H:�ｆ6u���7-�/1y�X�C�1���c9]�_as@¤�(�R���9�O-֡b3�� �]�1:��c�a�!�$.��������:���\ڵC�1P�w�/��[��3�y��.p���@��Fk��vVG9�4�l��NP]�yi�a+���rj�oy��걁�ԋM�8C7�8L�}���Δ�uX�|�qJ��C�9�WYE5O��א[����\��2��nR��{wB/��J脵��/�����oz{7���yS9��溞��cr��� ��἟m:�A�����p�)Q�_՝�4�w>��q��*�Ӎ2��W�!�9�H5��T���ܲ�8߽c���	9�X��%��S:�^~����,V�Iy��J����H+�H����텑<C��CQ���nv�gCR:y3ܫ^m�YEq�[����g{��*��?�aL�<�d�;��g�m��4�v�]��<���[�&��i�0���W�=_�eMlM�xur�`�����f�v�5:GG9s�4Q�|�֍���Za�k���V�xԞ��m�B�n`��#�oIg(/�6����<�&�=�8%,"�+�[���ՑT�s��� Coq�J�J�v�af�QGo�f-�VS��S�(F���K\��������W��9|�'O,d��&�!�k_K��}��[Ϧ�W˦Lß��WK�k�76u[⁇�㚞�9,+�K��Oq�h�3���4c6U�ɳ�;U9Ҏ+���h/��Ȓ�D���p铐�����]9�&�����<�7���5P\4�����Eu�U1D�i9�p��Ѥ��7���nsC�n}S+JW= &j�)v�}�;v���&�j5�
��]�Si�2�1�^!�P�MC�Aw'(.u����5i�Wc���5�j���r�3b�$�\&�|��s�5OT��ϠBk��_fҎ��n�[F;�#X�❋�Nm��AG;&��ݑ�xg��W����)����qKv���v8���eκz�3��@��`5:RY����8�݋q�������[;�����U5r�u3�Jby i�#ͫ�yX�@�J��X�n�Jʰ��
�\r�\�^��+���P�܏�4�V��E�2K~�7ם� zY�:L�gf
�j�g��z�e�]z7|ap�%��J��nո`ȽN�Wu����I���Y8Fo7?}�}�\�n)��{�;>�
�m�޸x�Nd��������>��hP�'b�D���.J��Nw�|�kx���s�9�eH�t�s!v杽}״c3B�q�vj=j7�Ҕ���-���1�߽�3�������?u��5yгMS!7����Cz�Y���F'[�]-�Ci���gi�G�8~�S�(��t�W�'�۵��69�D�$�j9�?C�oq���1;��Rn��5;�
[<���Us����"$��_�����B�Or��=��t�a�G;V��jԉᵷ�y7*�_q���{���e��I���p:3�z�ui���z-�һa9�p���v�\���Ƅ1�Mľ�uH���ef��)u��YG4��2�l�luæ+�%K~����rCѪ�}o�����1.��;ӶKk"f^C����+�V��l|��e���A���Z�2�=&�sޏ8ߡ8�¥�,����%t��i�QZ�V.n���rˣ����9]�\|���Zϲ�b�=�ǳڡV����c��̤��8\ꈞ�2^A>5(Ս������.�F�� �G���F���<�
���}�UH�h�w40�D���jͣՐJl�⹋�$��0�B32/��\�ӧ���Va����Y'*��/k.�E��MX��ؚ��ۃ*�c�H7��!�w��˭���4xM�������.gyn��k��u�L�3Y���[�c-���1�ޏ�۾x2��&�':�0��M����!�A�c����:�՛�ms`��,�cr����v�l�Y�0F�_��Vf�ͦ�q�z���zITU8�����1Q��.Pt�5��3�|�n���<���+�'#�%rCy�;�qY[3��Fne�ئͶw��w��S�л;�[�|��fTu\�!���0�D�W��s$[�i��@�i��ܑ��Օ�������坎�~��QԄ�I[+�F��ӗi��E4�B�7
�T.�ꀠO�4bĎ�F���]���m�ģ�=遼..��XՔyk�u��UF����ee,�wwͫ�fҦ��T:� �u٭�[�6;�dy)�7eY�L��{�nF��*v���ξ�j-*N����<�ر2�oq�n���6�˦i�PE�0��/�}��|��I��ޣ�{�J�e�����l�c17*�GQrL�j@yvƩ�w�%j(o+q���pA<乣�C3���TCv�}7*���xC��9�z=���s����M��ψF�s6�%N7�!��qX���ŃB�.F����UܗN!��R�|�\�F�q��I��syk�|5BӚnz�qN%�]y�=���<nvd�Avn���e�9]$m\�Vk#+'Y�1�_+SQ�눐�N����[�5J�ڮ��t[\��ឱ���k1+yМ*z�\���fS\����%apI���-]q:���bp�n�'�|�W95�M��T���{;PVғT�w�N����m�©�NS�|ԭl��~Yn��X��|�?+��#t���ҫq��{=2��5eK�?b����p\��!g�����a��FL��KOH׺g]6��/&�������ʌ���C�H�Ҵl��D@�텼���^f�ӧa=��$�\�屍�r[n��NՈ�Xk�i�[�"��gc�	��3�t�H(�]��Y���M���}C�!�A�����vm����Cܨ�l)�2R�����nV��&$��ڌ��I�㝎;\�ִ�{^���~��Bi��Q�<ey�U��f��ɋyI�}�ƕX.\>���i��K�׼�sг)#A��M���4��=����Ì���*�����������V�;w�`�`�ASj�ܓ;�˱Oi�eOb��٥��]�oq����_6�����k���{�]����vs�c��_L����K�¤�k�K8�吴9�u��8�N)��[��_ba@�T��Y���dL��CY�-
��]ѽݝ�W^f���HTB�������[�!�v'��c'�8���opq�� �)��q���0�Q��� u�)�Y���f�q4K\d�wN���N�+!��K �H.�{�*�J_�z�3�����]p����X}B��Z�gKԂ��6X�E����}۵4Q֌�����r���ީ��V�f�p�1͒�{ ����a�l>\'s|�.����J0ک��g�7����d��+�ә�#�.��B'���/}�D}uz�S�m�sʲ���E�)��r��e��N<�����3��8{@\��N[�E��ڃ�V�^'6�Z.��n��O9�s떽<ޑ��uC9Q�ێ������ų��16Rpř7 �,�+������\�}�z���C=�ξ�j{>]�������	�uI��� �G��6���p����'ڮ��Y���7�)L:｝�6�v�y4N|��s�O��Oz�g:�����3b��&�&�}�Y�/9Q��W-��F�z�jK�1�#�_{�����zҧ��t�&V�c��҉B�ȹ;��a����u��\��i���g!V���Ժh�d�m��$?�̚�j��%�aZ�k"y���޾z���ʱ�(�p\�r�M֗/~]2"WώP%��ՠ�y���]q�|��)wLn0��ָPG�]�@���)et�kk8�ւ����8���	Mt�Őd`(֦E ��53�Ey��<�9��k#+a��n��Oy��:�ujB��ٛ���)S�����)	b}q���+�X�l�$�طm]�XV���}��s77�ӌeONZFV�ۆ񼉹T��*/�0'�u�uW+��nqG^vԻ�.M�F�`pk��Z�ks����_��W��5��iĥ,F��k��%j(!� �Ǒ⩥�o<o�o���LTB�%85OU�ġ=y5��2{i�2� �Pw�l��C�Ȇ+��[V�*יJb,̩n��9��s��+���EMA\Ť���sù?9���Q�z��0&�¸�ȑ���|n�_"���m�vg>�T��:p���v���P�Ǿ��!̯5�Ov��<��&�9�{��Y�36��o���D���ዌnz�On��/�rk�Ω�7M����Z���m�&���R�i%}��|��eG;�p�jػ�S�%�B��YJR���#xғO෠#9�TV�/��ϒ��G��`�{�%[~���ateFG�2�^�(vv����ݷV�,��vwU�K̤�~F*����c�����M�ܬ��tlt�{�19�ܤ��R�I��m'm��h�WӅ���.���Uv8�VfU��f�+*S�K[�*f��n��5��Z��wj~�ꪜ}�C�����׆dj{�em�&ruE|u���i�6w�!p�8��ڜ*���]-��Z��gljMDK�����u�Y��y��nR-�A����� ��G�9��Y���7��鞨��D �h�=��S���V��	z��U��g���L���9
����R鞠�e	2tq��P�:^�A-{[m"��_^�\rO��e�{/o���1��IG���Ȋ\�j�{xwSDZҧr\�ܮ�|�j�܄���C3����ݥ*)�*�E���w6���+U:����"I3r�̂�����5��l��cyD	y"AY�:��f\p�_�I�/��B7�����c��6�zm�CU�enFc0G=����V������7;#�[��]���ˌ��S���t0n�x�ݫ����}�-[�����x���޵��I?j��3邋��I�I����m���P8	[��q��빵v�f�F䃅A�h��1�����
�rn�]�5c��{�K�v�*�n}7u��MgH*汔��/':b�\���2nm�}����k�%�LT�mܩλ��W	�|9��F�m�aB�Z	D�(��W�r��a.�fC��p�,���A˙M����Z���j�2Ļ%5JkmM�ppC��ܱ��>]�-�������\�� ��6.�w��$�O�f�4�K����
WMX+p���e���jT��'h�X��u�w)�sGm�ghLΪ��`�&=��[�k��&u4�8�BX���� 8�(\�_%u��@+���Ќ�q�khT� T`pT��6�P�rf�-��-�	�خ���F"�D�f�]҇U�8�&��8H�ͼ"X�q��VҼ��#c�f�M�|~G9���	����.]�e&�̇�,Kp �:�$��0h`�N�c���^!������w�{oE����n��xQ����8��5w+安sm���yٚ�l�d�ܤ
�)T5]�r�T4*L����o���s�*砫_M�e�&G[��z;�]��e����C�^�o���\U��I�Ө��߻�.�Z��P�F ʕo˙I�X�{���op0��Ҡ�9�S՛�0�Fn����%]s��坁GslC�E�Z�"�/���E[U#xL��@�'6��j�xMۈ��!�Z@Ǎo=X���ܭN��nViLP�|�e�1n�}P�Ә�bՙ fS*��ƫ�E�{8w�9 fL��=���I�`�4Q�a$�.*͒�V�n�k�0m�[���}"�u��r�������b�#3���7�O9_�F1)��/[�:�X�(P������DC�f����̖��JN�5��	 �R��o0��2ʚ�^1A��Ff��=��Zj�{E��Ƹ�-G�/J�K�wt�g�}\2��B�Ju tv���X>m3VFT�K�Vg
z�N΄|9��9#���vq��9ve;�N��J�45��SUf}�0wc���l���˩�����)=���¡���*�O��٣�V�OM,�b	XΎ�V�9��XWYk^͡ϓw�bN���f���ԧ>�D��b%2}����]���&�s���;9sˢ����P^uM�*��㦮�E�ؾKG9����1��꺰�Rk�u5�9����"7A��҆Qv�+�W��.�'Qm���G�q��Tz5�k�`zlNb���9O���b�Ε,����H����o94��cl�+�ê>;���\�#�f��WcmR5fm�mݣO���U�n�fr�{�ĭWNbr�ۥ3�a�5��b�p�xI���C�
��	�.�sq����nXX���Νv�Z��.�1��P%��!���� �p˶1i;(��b��:�I��efҳv���Xq�Kޓ3�ۜ@�4_R���|BE��/+� T5�J���b ��#mKh�1�eh�Z���X��J�<LEF*bQA�PV�&V���Tb1��5��Y�F�W)`��Z�A",r�2��*���VEb(��cE��*��[LF !Z��+ELk�UR�*1F�Y�-�IQ#Q��]5b����UQQ�D�b�����Pb)*YR��*!Z�AZ�FE5n��9h�+�Y�b��UV,U���R)��T�1��N"���U�&4b�ѕ�&4E�FDF�\���Z����1��e��@��V
��FT�LF1�(���T�ETU�Qb4ʬq(�UV)�V�ёs3+E����TKj�Q�b��[(�i��c�V#�DAU�eDB�V�U�Q�DP�+-���2)R�#l*�1�AW��$�*��m����"�uo@�����Z�B��j�h�'%�1v�"ȜU]��*÷��*�{Cs;M�P�U$���ܲ�cx�iq��ѽ��6-$�[n9䭨�bk⧪quļ�&�d�:���3����+^�&�;�r�]�N�8@�	��V�s��MK����v��� Ns�[����N�oG�S9�üu;��6�`����|{�1�������1�}4vwK�|�e����ny�~�)n9@�he�+���\��Y_KU�ùV_�W:{�Vr����\�9hrA��5ŭ9S��M�n"�Tm(d�]i�������%4�9�E*�V���L�Ի{�zpuGt���-
��
�V��T..:�:��Ƨ��[��s��,gVSZb�T�]]��˚:�9]�K��W�]�x�]���K{�����b�G$��5S�
�����l�3NL�@P$�"n��K��Os����G\o� l}����mMF�ܾ�j�p��ڞ������094�;l���-����趇[�*^�6�:o׼��u�/z��%���8�U-[݈AQ�9X�r�}�V,�5�����d��a�f�:�0�/�P�q;6bL�'�o+���F����	��R��^�����~%LLF�S"��'m��œ����s�����n&ޛ��uä*�P~?2vv$��Q�۞�ΕPêh�+t$x�o5�vͶ��
e5)GN@|5K4�����Ԇ��ϊ�U�W��y$�S�5��cb�Z��hu�.��K������]Ea��Gs��j�,��(���q	�	'&q�NF�x$]��z:�5�֬^�ųd��vX��X�M��͍���;����;��ێz�2�v5�k��g���6$�����Л��/4�v���Xh�sAI�{�n���{���UgB��fs�d-�ߏ'��Qx��\�e����Kpq�K��Z�f����!�pc2���C�Z�
���b�lj7��R�%Qy
��;���7��;v4��!f'S;^���',�b�s�*�Ri�����G$�R��Y�X��yՇ\�Soᕅ=�X�')7�`θ	�uzZ�E/S/��)|�kOe�'�71�̐�@�-�>����5�Aru��;U�a���U{q��c!�|��3��&�9ٓ�������%��C�w�\W�Q����E��w��q�Ħ��:��+���9��x-6'��&��%���D�sk�}�m5�C�Ș��k���ĵ����w�=_�$%��P��k'�܈}-��'"��"��z�����h���Q����(��zT_�ʸ��7Ar�u��{�����*�q#ΰ��d���������o&�/��_0Od�}��C�Y}=�|�[�!�C�L�Z�>��X���v�D��O��
��[� ^V`�S���i��anۄ�̜t�Ȇ7�l6zm�|�Z>�ij�t�
�.�̜.�n��s$��<��F�I�e�1�n} S����d�8�]&�Pÿ�7s��AvV�qw���(��3�4��Ym ���bӴ��:�L�i�ꐝ�e�YE�t���^�7v�����D_����Ъp�3z��>�v&܁J��ke	N�
���%9��ߜ}F�ϠK����W�LY����j4Z��ːYD:��2��VmǴ�B�7����$=������q���r'w�ܐ��4�;�eУՎ!�]0C l���|M�F���Z0zjE���y�J��x&�*MN.������{k�>�y:�f�tr�1�6�j"���<�ݜ�N���z�۾x2�ۭ������F�6���嶀�Jj+K:V�����J�oL�ڜ����59��p�Ug���4@:'�z1���i���;�i��q�(=����W���UǷes�[����?v��^��rJ��ۚNNDꊃ�̖[��=g���H��B�Y{S|a��5�(��q�\_���Y_H�<R�T�ܨL��z��h�unc�Z�g{>/U�����Ƭ)�y��B���n�a�v�.�K�%M���!��}M2���v�	B������k��>�d�I���/�v:�6��
o�!�k_K��|�6f�.�++��q�����I�Կ���D�����y�5�g8��6�~�G�f�Ҿ%�ے���˭lS�NT������������.u�c
��5;�l�U'֒.�uؙ�,��;
�M�m^֖�9���V�,4i�ɝ6c���Qs�Ln'-�CvO��}�)������W�zⰎN���6��u{/a�X_K����t��Y�!��t�S��l􌎘H�]i�#������ЦV��2�OJ�B6��ZM%�%�f,�=5F����3�-7�p�2��I\􀙠�3x�ێ	������t;]�v�H�	�/�/!�V������$�ue�u̒�2��Vw���WN
}l�i�	'"�M�<��Q����OT���Z�,j��(����6���{��K�S�c�q;�5��ľ���2���6Nu���N�L���[��>�z�o|U3�����z9�Q\$����HK��Z�p\�D�w;�ⱘg0��\�*��z"�'�s̭,�r1uv\AV���vm�xH:�N�ԣ��u=�ȑ�b�I�D�\GUrs�O�mo���8�c=k�v:^X~L<�_*�
�w��ˡ�L��r���v�hJ����&ݝ�&�;1��k�z���ͅ����Xڄ�:r뤶��B��u֋�H<�.�t5�a�գ�zay��9{��Q�<���*NX�t�6�/��t�$��fݲ���w��',�DFa���f�֣{Ҕ�u9�H�9M3���C|�N��rM����2��,��+�rӂ��1צբ�R��쥸�g"�g>U��
)�*��QOz^�tT�Y3� j���%��K!b��}-�|�_6��������ݯJmzoB�yh�Ew�%�DH��dB	�U�~����#����vK�h��5�fv۶�j��"Rsq)��O�����pA�U����s�Bby�6U1�.�V���;!`�䈨ںq���;��J˾IB�.�ǜ*id1�ӝ�m�n�S+ ԥr�I��/�[�y�狍��|b]/Ȯ3֑k"f^1�S���hT�_M��[�T[G��憔�VKf���?����Bf�I�r�Q��&7�l�(�vD�N]D��o .�ȍ���;�\"��ɫ��Sλ����,�4!<O$܊��C�Z�|sk	JŅ�3]j�#�AC�t�*М
��ػ/{�/�;�@Ъ�n�H���^�v3ëdΈ��6/���F���C��4Q3&ۖq;�]�=JS�k�du�����*��EF��F=��w��Z�+�WyK�N��)U�w������1y:N,��fʯe���n��z�q}�c�#^;C���[�����:�fsW�uh۞��-�n#v�tg=:��t�Y8��bNL����/~.we�b'u}Y�Y�Eto'��$�*��l�}�b�����r!;���n�f^��W��:���d��,ަ���}}��t�U�^uޥ���RX�'F>[�&��B�L��Gc�Y������)��P���j5�[�k��kv���쇯E��zf[F�qh�Ϫ=�����2��FP��dڴ��wWE��A�i��G�cZ3ӗm��E4�Q��P�g�(K*�$�兙�1-�wN6g;��6��i�%r2֧�����ɹK�;�P"I�Ֆ���0Y�mm6�
�	[9�Rd0�r\��ft��6��Y�ܪ?q}(c�n�2愁�It܄���x9[B�^f�_EW�S�ζ��Ae�Ω��u[���C�/�	���{6��K򼮛yз04�қN�
C������禤W����omV�4ob��8[���[{»�v�˅��d�ŝA�ﾃ�1��_5���OM����F�2Xi9�Z�l�z�[�1��:�v⋎��o�����K�K�)s�)-��	4�f^1�D��gGb�;R���ךa�,b�!��uU��r�\q'�����~s�ࡽ؝w�G0�-��ded����2Y��F��U�".9���;T�D?95�_;t��lYmr����Ĝ�m�8��g�xj�ǟ�l�vq˯xj�Nur<�r�����[��x�
���N��L��.��2����jx��EMU° ���xғT�v��Og���m�ϊ�u8�W��M���0��W�ݏ�t�/sǻ�a�|\BM/�(.�?��G����.�s�W��$�/Lm��䄤��ٻ�9����U�V�NON�:��|��4%�M��9��P���p�}#Ok�<烯�rv�ʑ�0z�3����]�%gE�1z��l-�,[X�4����j��7�c��׊s�7��m��*�OvM�+ާ�-���5�b�Z�����z�ڲ�,d_�Pc�w����td�+��<G`"�R��s��`�K��Ό�#�rj���U�|�
�k{%/��uU�ikq�V���}���|��dC�L�zV+�j��������{�^v�k��:��P9��r'��{-�Ci����ZQ��fvTU���evU�&�=*{��n³f��o��kr!��m{��O^\���Q��y�4��wu)gRn��8��5<�7A�R\.'��\��gK�2r�`t)���͙\��(���i�ʠ()t�Ig���7L�CY����4��[.�h���I+�7e�� �T?��^P�^U��ڦ#ȝ�F:;qF���mާ��&�n��4��vͶ�-�J��%s�)�ȥۣ&6�+ec�|I��ק��
,6̵����lW��(��yЗ�W��@7���	�}�W]�O�%�.Z}A�����s�[���AS�Ge��\t�Vs��<�9̨	n��}Yܻ�b❋��m���R޼���Y�۽M|��4��� �۶0r2��D��M���(���u:\����zL [U��;����f�j�frK(�0V#�L��=��s��
�0�w/�,� ��FBż:�(��V��9����ʢ6/W��<{d�^�	7'���;�=�6��/w*��ƧMn��ܗ)j�w�Z`��u�'�g0e靨�.7WV3sKgr#Jw�m���@ª�K�˭*e.ⷰ�4KZՃp�y]���;��և�������2=�ǹ����z<8�qU�b�2��-q�����oP�~��q��'�7�`-�+=�9Q������si�"�d#���Ӄ_��K���v;a����+=�.:G6��0�p=8���Kq4�E2�B�=ӷ�f2*���5�\��$[�3&��Aw@��IZ��8��޾�����׆�3���Z)��KϦ��B�Q|��	���\-R{��T��#0�OQ�2�g-8J_^3;pݷ+a}ƾ
JNr�G��#�|��+�Oզ�ɪQs��Ƹ��g���M�cm����M�w`�U-�]k˂��@\��o4*��:ꖯ3P�z��	Jr�`�LI�s��F,0�C���)m�<��0Ɓ�\�Y�א��ڠ*,�o
U���o d��"anƣ�h��������CKdG.���ۛ�3h':��,LYgՋ8��x�)>Z��!=�Ѩ���� <)M��(Þ�}v�F�����I�/'<����:{����q�(�n�5F����e&ˬ��\��n��y���ӆ�^�sN���z�Fm
suu鷷q�[X����7sJ�"p��.r|���R���y�[�b��\���ɰ��\@T2s�V7y�]����f��-�M���j 䅅x�kT�˝��c�;�h���N"�Yv���/r���V���(l�qN����kU�9��Lإ��c��rVn���Λ��bj�O^:�4"�}��`J�46���bފ��	}Cm�C�[������I�jrM��-Y�I�fj!��B�Uo<�b��PW]����}�����U�D��
I�t.B�*#w4�����p�պg<}�����c#K�i*N�׻\0�&Ҵ�W]���z���2��w0�[w%1��O1y�͢��wT�%���;����k2�Ic]vN�Rz�q���2��29�6���9η��T��0�O�K���1����7XX�{
Gr�ۥ�:�Ӹ��e[5״5u��9��H�ӝh�dn��>�7'�Ù�e��Y����������+�Y��T��.x_c�IL��zkK��a�-33 *���ۺEc�mD.6 ��t��(<�eJi��VĨ�F�A�L��f���V���b��>��jy��i\�0�|�[7��@�HO�ǩ ̼>�>���wC�;x;|���V��kf��vâ�b��.p}���d�"=ѵ&ê�Bu�髞��)�c&	��ѣ{)cr�u`p�����Ɩ��"�� 	�n&ua�z1B�y�D�p���!Kh\L��ACp�X���sn�C{��ugc�}$o�ޅ'-�𑎴e���VmjE���ժ��m^v���s�R�pQ��A�Jdww�]5P�S�=Q�	� ~q��LY��<�N�.�r}Y@'$�[��oZ}��B�J�(ச�gk	���a��Yu��Q4��T��,�>G��k�r(���)<5�K@��$�I��}Ӥ�vGI�Cs���{�ܧ`��mU�tn��=��mCkBbp,f|'�8�() ڽ=���{�L�is�6�!�m�k�&w8�w,H�We*إs��8�9X*�oj2R!�s�����V����ܩ�H�_\����+���t���Em��
�t�i�!�'+6�h��/��B��9��s&w#9Z��U���l��7���Q+
���'f݇��"w��si\a�,�,�����%�^>6��g�LZJ�Ƿ75��&�y�f����Y�7l��|��^�;ݔG�EU��(�����2ʪ��UMʖڢ(�����#[�0Uf4�(�U�FJ�Q��QAejT*[QVؤ*+��1��+Qb1
�"���r�ŢȊf\��3LV$�mR�DUZ��h�A�
[Z�1C-�,�ʈ�r�2��Ab�A����Ĭ�-e���PPWV�D-��@�b2bULq�P4�+1�S0�6�bcU�" *����W��
�V�a�`�.e%lX��d(娢��PY�Tb�9V��L`�X�ˊ�`TZ�HT�U��V ���b,�F�@q�4�D"2�YifR�r�2P�Ld�1ҰT�U��V�b�5c����lF�f���+"����h�����
�"�� �RE$�T^<xl�{P;�R�$9�;�ԝ7V��D�;gw�l�`a�X�4����U�@��2������!"Q�״��9�}�q~\�d��o��7�8���9��l�luæ)	DJ]7s�V����m��pڸ�V�����_��f^D1�V1+�������\��d�}.�x�;�=r���W��Q)�T�����F�B��$a��t��;w��,_���z�ۻE��\��a5b�Tã��x�P���x7H��z��y,���>�=q;�=��\���t^���<03��snƫ!�K�W8�l�p���؟]�x3����n'uy,�kE�ݍF�#�Jm�Iv�eU>�I�i�a�޷�e�s�a���ء����ɼIOU�5�#;��U�/Qnw���'{��۱�b�\��-�{�������gi��}=�Og�ey��ҋ��ڒَ1��aK�]8�����p���n`T��w�E:7֡,��j5�0����90nM���%/T�u��Z���g�=�0@����}=�j�_������Z�nW;P>#nT��[H�C���!,=J�b��͎V]�da�'���//P��u9r[���/�ک�������s9=�BY���&V$��ܹ-�O&��b���}�a��=X�>�d�u��Gϱ]��~6�ԲP�QL��'�V��{8�5GFk֤����z�>�p�9�yp��"P�9�I�׸�c�>�9�f�I.����c2�d>�׌���z�r��ؾ=B¦0�¨c��=�yك��L6A�L�|�4u����1�˙Z�`S��X�^�X�p|�a9$��g2 �W3��K�}�����wYq����f�"f��f��'�l��}As��	\.3�	4��.���Muw%ƟF=p�;��-��o�7�Wqx鋎RO�Q�I�o����{�?I�iq��V08%�y8�!�J��S���}kn.=[���MDj��ɲe��J(��q���V/�I�mƳ����j��[U�}ֲ�朘��*/���C�c�$�F���x��gS�-��'�}�]熖�����V[@�7�(L�`_(���!iᏥKj���}Xe�ǻ.D(�f%]�J\����[�"�Q�^1Ĭ����:�tyvu����t]b��pl�=|7�/��N����v�y�����8����Q�R�\ͧ9=�AA��|C�eـ�@��WKt�����m�©�N9����M��nOa�	��+oR75�Q[�1��ۀ�n��������Ң�{	���F}�f]�\��/h�J�6}4��}ݝu.�|$�<����jX]�N���3��xګ�����V��[��������α�ܝ�y#��:=Jw�S�q�1����$M������(�����C��j��g=1]�A��S��}�R��U������K�{�+Y���oͦr)�qV�l.��g�*��dH����ֵ��q�a���Ֆ�g��[�>����
���kI7wI�8EޠmaZf�˦z��$�KH����K�¤��k��Ν�s���Υ��T(Mvb	�|�/�ʅ)t�Ig0�n!s5n�<x	����O/:�WOY��v�6zn���
�%Q�(sp�\� �u�8D��if�n��&��[!����)���m���]�����*.{Ќޥb��Z����_ۃTR�-�4P�6l��sa乓ԣ:�̦+U�n��b7��F:y�<�E���=!Rĵk��4�e���Rkd�Ε��iш`|�(B7���u���=�D�4��cy�;����v���Kbz@L�f��m��㼱܊�TL�k���E�m�y���������}a�K��8E]8���TU�	�;��yiud���\�L�I9q�%lTs�;���6*���+|q�-{�YsMP��{'�ԢP�s�bp���zafa��Ѻm�����	`�������t�M.}��Gm�(>;���̓�M�U&�wg9ˊ	���˿���h��޿��t����#�����o�Vq��d/+w�RN���"b���ka��oZ�|�v�,����+a�]ط��|�8���=����J(�- [�����;Տ�9�i��ŝ�ʍ�T���\�C9����$[��i��o7�����&�{5�Wݼ{���;j��zf�Wu�Q���-�M2}12�؝�2��#�N��������Yiv�7�`�t��M����������l>�a�=(�R0-���v'٪E�*R��tK%�δ���i+���I5��r�D�+2�:FR2<ȥ��UMzqv�]5�E䚪����`V�����h��1s�"+k+V5�t�es�ܚ��zV+�G���Q�|b��%/{}�驅�+�s܍(rX�ާ#[��m��Q]��	B��#ώXa.�g�x�}y؛�֯
�_��}�>�׌��Cv�Mʥ��(���vW�f{֑VZG���s��[��T�S�����p���HR��MD���i�d�w�D�T�C5L�p�7��NB��C�k���
��T;P� ���,�����%W��ծ3���Ϙ�+ج��ǳ[��QW���J�0�$7q=�󫌴z���R�3b�I9l�+u���L���#��6+��M=�>���s~�/�>�\�נE۷,W(����°��Bq�"Us�9�z0���scms4�Mc�̀ъ���=iv�*���Ɲ��S�.1���}��rz'��Ԡ�1"��4���#8l��|�:M����GE�&K�h&�!#Z��&A{���G�<o�)��̙��9��om{N]�W�˺�ݺQ���D8/H�6�P�� ec�w��O���\�IΜu��	�v)T�K�̊hO�z�z�9Z�$�����-���ߙ�_��h_9�uU]{�VA���o]fv�$�4������nw><������!���5���E�'u�ʲ#ب;��fu�����8.��o�<�t�T+,��-��2�ڑ&�x�m�L!Lh�v�hyP���Q��x���p����9m�>#��nz����[ߤ�ϥ����	;�#���.>ݷ�ޤ
&w϶���O��{1O�:�Ra����D E��p)\<�^CS��)�2���wA,�ܸZԻ�/JV�k4<=����~�;���}�\M��ѐ��3U^K}�3�7s3�_ȧ?�����=ˢ3���ɼ��~#cʇ�#�Q�Y�z�|=�#$18%f�uW�뙑�
ѽk���}��7�������Z�ϣ��S��z�#ʇ��dWW�؇U�ss�!T�2<��\|�ށ2���u�3Br ^U���3�Rg��jX޷=���r,�=�Kq�|bI}y��C�;��\xP�&'��T�f�Xd{��6����ߞ9�Z���?~?��[�"d �ǓJ�%��"3�q������iR����1���T�C}e�2r����D��Ly�&m��
S�YZٷ,b���l\��{!8u�#�k)�<]���j6]>X�c��3m��V��g��;�e��wb�t��WL���f<Zvr"f���~�*�|��39��E\:�U,�-� N�3~��a�אNB���M��������K�O�z<�*ޥ#ޚs3��_L��#U0��`��M���L�%]��u���ҳ=�e����*�Y�25W�{�3�Q.�{{j�®NH��)^�0#`����E��l箉9���7���f�b���~�����;A�Z<(�����vNK��uؐ��މuY��������Y� �6���6}:��lo?\�S$,�w��~��]#�jZڿc���UB�t�.���y���>�T}����;c�9�����N��a�"!�G�H�]���R���>��U�/O���]���u�T�7TZ�1p�����ܝY�ז}�}\l�P�\w�o�����R�V�9���}T�H5
�T���LzC��].<�*7������z�+"y߀��xx߮�q�Yv�\���4  )�~��=��|�{��֣q:ԿE�Q�<W5��}y.������?�_�G�ë�1�����r�����{v;�&��^S���o�*T(
7A�(��Gz?�md�	f�Z��`��-��l��vЈ���A:M���@�]F�#���J|f�r�v�VR�*�&�QqM�T���Y�!tn:wf�w��v�bL�ٳ��7�9�0Cp�������\n�+ɼ����;S�s�6<D{�#��3���v��\�<�o��9A� X�LԄ���z�T��+�"��58��:v<������~������I���3,���ޏz��z�q�<|�ĕp*M쁀/�\41�,�n��s푮����V�5ef���EN���w�����t:��Й��|�SvdD�=�=��o�צ�ٳ9��e�~�F�5�O���G���H�{�fsվ�Ϋ��BB�RUUI�����)�G���ߢ����B��ʛ��6��2=���~�Wxl1}3p�p���q̥N$�6�j�Ho�85���y���Z"��F5����fP��߰P~��C�ߴ���t�6�������]��<ǀ��N�#�KD\S]�;�c�zM�%��?'�ʜ��U�~�ւ�����{7�7 �w�������pi��v������}�>YL�"����f�_/�������_u�������u?[��lki1q9B�&��EG�I�,߭��� ��o�yƙ�>�S��}���.��qݵ[η-ݹ��_[�I��,�r�"u��3`PPȖ)BU�����k�v��;x��V���-�tC�t���cf�P�9���.���c�u+�z��������{��˂j�֮�T��!K3���!k�#�[>42]^vvvA=l�q��C��6<�Ҽ��◎�����ƽ#�eS�p=],��t���=����쳶t��^v<.��"x(������^�;��y������Ut���8u-���@�?e��*h�<1?PJ�[Q�_���镟O<�nׇ�m�߂߭��;����^��83~��k!_z�+I�p� % �zE�<�A�r��5r���nD��NuC��h�t���B�ǉ�2��u'~��v�\C��&��<�%�dB��x��w���G�ES��\�f�����n|�bFz}�3�V'�!����}j^�Pb� "N+��)��]�xjl�Q�*���˺}OQ��|��ᰝ:;�����V'��O��0�̕]�Kw��D����n���5�h��"�7��#�����=�ʞϽV�0$1��J#KW���Sc!�oY��k��Q�Mt�D� �T� �V�l;�6#}\s�tG���z����΃��cI�;���|����g��_E�\�[���W���O�Y�s�z��xo���62c)�ޗ��Ӹ��jf�$_mď���.�*��k%�F�jX:��"����fE��y Bgh�EN�_;��>��3a�7��[{��L���]�b�r���UwB\����o:.�;���VZUy��e��f@=]֯nV*<H���p�|��p�&��&���f�c7)�W�	[�g�O�q�fT�E.=^r���'_!Y��h�B���ǆGL���H�T�7*Y�qt����:�����eי���NC���ز���/�>��yC5��}Y����#�|<�u?[@��(`�F�,��OV�xm�A�k�n{�	�ǳr���69��}C>�e����rT�*��zBk҂�>�c�����4oR}st�g}��d7�{�b��ú��~�^��"�{��#<5��W�����z�"A::;3�;���W�(2�,Z�p3}~';W�����=:�׷�:/�|����tҷB��D��?��ϯ�<�۷^��Cۉ��9�þ�g�bz�ͮx�NE"���^�f�5{U2��ţ�t��k���[�<F��mNrۢ20x�T=C���q��{&�}/��p��q#�����GZ�ʰS�������f)��w���O�Ұ#�߈���/��v�'�}���^f�[م���D�p}%߸o�vǎC�;��wإ��:2 7�^��o�ߒ�ʾ5�"kz ��.%�
����(R��\F��k���ݍ��n���e���;�y]c��'{��oc�1`�E^I�[�+2f
c��i E�8�oD�s�q#8������� ���5�g���e�����q��&�L��գK�j�|��ut&>R��V[�Y��ܹ����h-��Ja1�-�r��E/�9��Լ��ͬޕ��[���fJ�<���>��5�f��*���l̀ZM3I㦪���(2.�<�̏ '6HL�yڜ�R� {o��d}.�K���rW����X�Q����l�B�@���Y]Zb�Ǣ �da��EY�����.[g3xd�"{qi���#=���X��⥯�H>�Zvԇ+p�o$�n�A��1hY�V������z�
=�F\����gM�]�sq+�#k"��Z37>��
S��۶�.K�?d�L�P��E�x��4�!61��9m����J���]��KB@엙x��k���Q����F�[]V��b�"��}��oq�*����<��[
���Jn�������)�{�t?>���|_j0�+h3��d�U�.��]Q��:+��a҆��QU�����z����0ⵦw�x\����g� e��D��}F ��b�4��y��K��Į�d����n����pܭ`�K�T�6v���f��������v� N7puY����)���Ź ��6��ƟEXX�Y��V� �q�w��ۼMmWC'b�\�K33��4áY(
Fwb��/V��-������kN�@;��Y�0@�j�Yh�\�]��-�!�)����Y�Kx�����N�3�v*brh3/�H� >Z���5kN|nT.-���������i�RJ��Aq·xl|o��hW��lx�u���?��da纶Z6��WIZ�La�Xz�N-�pv�Ut]���m:���)Z��ֹ�.��!foC�,��ܶ��V���3*�L1M���T��T�9�D`�8�=I�R�XY�����X,\��w_<�Y�p.W)��ݧork�&v�����G�+Ub�/t�f���G�f�9�E�����;�uڦ)���i�S�U��Y��	��11I���V3 n�Or�d5ʗ�R���qY,R.���0��W.�H86:�rs52J��4#���u�����խ��Ux����k��$��G|%�$/�}��%.[A_\ɑ�׌��K�2�o���,��7���v�r&vf�s�Z��Ɯ��W]1�	SiÿI׺������U`���/#ps��h;�jg'�ۣ��F��Ay�7��u��4n�Y��i��ח�X���r�o+���m/�(n��<��PN�[&�0rړ9�;{t��9@ૢ�֨�s��2��qTƗ���Ã-P*�Nu� _dٯ��ykj	�&LyDZ�4�ܣ���X�,P1���V�L��,PX�)E�fab��2W-̳�X1.P�1+U�5*Ĭ���Lh�
1FaG)�R�T��dL����r��Jъ���-U1�d̠�D���ZU2��.R��[AE�qqZܲ�֍jŅh��m���QU�L"�+ዊ�U��+3.+%k�(1�j+KAQ�Q���]0�AEFE�T�V��1
�E��l+��bTs%CRQ�bJ��*��b��0[�6���[`6�V+J)\aX入[�22��`¤�s�jC0̨�Ķ�CV�R
*�+SJ����#[2�nQE�ƨ�U�1+���Re�m��Ԯ[�l����pS2S�YPY�`(�ʺf��ʺ�Y̡�
�H�RT(���1��L�0E%E&&	��(����������	�g{Nd�WJ癮:��f2RGj�r:+J��z��Nd_Di��/���c�05�p�X�B��j#�=�����3�r��!㼛ƞx� <�C���d3�Y��#$1���p�s��Q;�淸�G�Vzzf��H�~K�~��z��zw�ϱ��T8,�{"�w�y\��I3�����-n�1Ӕ8_�L�"e�HlМ��n�NS>�&Tz�����㞓UR+x���5�'��g��{�FC�\U�A��&%��h��R��a���.e`��Y���\O�������݆�mh�t�S��<+��d{޳3���E\:�U(�-�������E�G[�s�nڱPsݣ��gܑ�ϡp�#75~���Z���L���}3p��\�L����ŀI����4�����|�Oy��7-ll%^!�mǗ���(k�PQ�z�O��N����T0��^�zt��5���{!r@z����|:s������^nCߓ�b������G��i:�@哾Ge�����Eh���v�,���C�6z; 4�� �fϥ:��_s���=��<�]��C�\W�O�μ�ӻ� 	X��}5�!�����]#{�9�����Kɏ=���W�4s����a��u��S/R�Q�3�(�˧K�'���(��]�����7E2q4G�u�m�+A�,5&kN����U�ڙ�y|\R�XjG���.�'O�,�G �Ve��Y��p�6�pK/�����U�8]�����s�����y��G�s�F��Gn�N�*`wHn������,���������*Sq-��hx���z�g�q�9M���t_�;ʶ=�fV�y�S��h�� ��ꧢ�Q�]���^	o��=T��*�c�x�|8��=���/�d?�ő�W�\�ܫh�4 +��F๫���D���MVJ˪�PmTӧޫ����##�c��=��y\3�W�4����u�e��0��++<���	
C��HzO�Jԛ��;��o���;S�s�6<	Q��t�+bF�,݌ݎ���N�������`��s5! &�z�U�r⽖ޙ��o��G��J��^��%�1�>�����JkG�~�~��LIV*L�D������Y̙��}��qx���Z�ފOx��_��Z�]u���� g��Rs�]��uAҙ�n���_Svdu{<%0�<�e^������}�bᡌ��8߱��z����G��H����g=[�W�����Z�@FS�̚ճ�l��'���o".��Oi�2Spq����{�������z��=Y�]~i����c��*%-�{����~��Zŧt!o�\n���+�OE��{+�e?����4��N���h�]�N�ԥ{�y���w���;�lZ4�^az�[Xi�m]ղ��']���4�S7���0q�[BS��gZ���J��b�IF�e0�����6g���j:����/�x[����z���]І׬PL8�wv������~��.C;W�1�t�P� �N�#�^��gN�;��nIw{.L'�ʗ��Ý޼�͞���9g87�Z_��^ ���遇[�Z�~'��P�D�p�����,�G�|VzL��P�&c1ۣv��x�X�d�;�m��
ȉ��8{�V5�������eםU��(c�+7Q��֪��q��4{=l	��b�Nû�6!���:�+��9������T�%V����z7�op��g��iOz�=n�M ���p��#�A�`S`�=�V��C8n�u�Z���k�zI_�\�
��ī���s�
�Ow>U<�Q<��2���~�੫����Ҡf��������G�-�b們���E�.��a�r��5r���nD�B�v�+S]~����*�̝�r<�/[�)lz�������@�C�J��	w^�k\��T:�{�rߪ��G<9��U����M?���9��K��\0@
�&�W*���~�>����Xm�$��p[3S7���k����N�v��uv�9�Sɝۡ=Y�x�����]��%��[ѽg.|w ;n�>f`����)��bq�y%��x6�P�7a匲a�g�ĤFd��h���v}
��Q�z&��#�d�&Y�����;B�5��m�Iv����y�
�{����6'�f�X����=>��u3%U�A̓��r�dv������.C��G�x����Zo�"�^��u]�����p^�]N��V�\:�3���?<l��<X�K誙y+R2$/;�SCV�l;�6#~�q�1ު<{�ȣ�w{�G�.\�gM�q\��+>�T4\;�)��;�\�[��څz^C+���\�3a���r�,3����W� ��q�7��qJC�`^��!S7��ѫ�J���؟L�&D,��Ǣ�y7���X�T���=�xW�O��雇�ʑp��n$T�2����������̏U��l�2�A�︓����yC>���d{��g�ɇ?[@��8::�w��ߊ�/W�#�	�>z=�I�L���nC�Oوo��s>���4u��N|���pפ!w�E)��E�^���eb��@{�ƃ+�^ڞϖ_�o~��Y�u~"5�E��G�dR����7� q�� �?`�9bٸCw�~��� ��_��EK˭��4��n�s+;�cӮ��}"�]�h�u��x�T��fL�*cV�hM
�@G��d��I`a���-��Vt<�a
�Y�z'�X��r_����E�̘/<�\Ӑd��\&�y�o&Ћ�&�h7"���%j�F�3u������t=dQt��J�t����%V=!�b��έW-���q���m�*Hg�s��1۷\2��*�ב�uq^�X�|2��������ԣ1?W��h�3�}�)Q`�/֧�߽�js���<R!��F��E�����[��u�O���m�+©=���<��{��r��Q�����j}%D;�S�mԜ� .(/�J��Ϳ5*:�z���G�J����4FB/2W�/�hx{�<r�l_��Vþ�/~��;�F@V�F�|�}}�Ӟ�xIC�g���9u\iJ˪�v���O<G����s|���^�x����O{ݑiJ��/��X�2M�S0���! g�߆߽jk=~�=:��4;�*
�-8d����GAk�7�Kގ����4�w{�a;���wbX7�UP�9Y���_�9Aޥ�ϔ޴xW���l�{ֈ��E��\U�A�Bb[�@�������v�p�A�@�M��i�����]��\��6����@y�WO����fg#�슿�W��}"��$	�f�b�y�u�v${�U�ػ���yi��M_�/��Z���̟o�_L��r/�L6R���b�þ~۶�Xs�T�0��#��C��+�&��9�(!u��Qf]��Y���)u�^����K]�U��z4M�VG��ww��8�v5�W7�h��"��r��E�j;��n��msp�� �8vBs�5��R��ٓ&e7�PZ#��*�|�����}E_M�n[`��J�׻#����O�P��S=�����5��|_E���1���Un��^���r]l�.����������^nC����o?E��D{��4a�T�����ɻ�)E3�~<���ǀW�Y�����:qc�߸۟a��?	]��҃y;ɝ������d��K��䅑�9/2�KvD/9��>���-�H�X�g´���"9����m-�}��v��ߓ��ߋ��#~h��KBq�2aU�n���w�ϳ?4���������_��}.���.k�/Z��W�7Ɣ{�̭��8���ǀ3�ꧡ�[)W�b�=k�b��	��eOFӪ��R�� ע^Oz�ax{��	���,�;ݮs�U��h҇v����}�^x }U�뚧+>��*���i�>���"O��=�<=��	�M\3ba��Y&2Ǉ�ᖯ��y�����BA��b|��t�I��AZ��>����������S�kok���#zy�����yG��s��9�|��V��/���B�~{�x�+�@�Щ��������y��\j��F����~|���m�5��)[��vk�������l�}�*Z��@��αgCu!�X���m���mu>��U�X�Uw�	��"�a04�B�V5:�͏.��¸L��p���Fr�=�,*�_��捿��c���Z���g�=�9C�ؘ��T8�� �0G����{kM�%��hz �<��~Z�]u���� d{�u'#�nj��WL�uP���/a�+��/����%�n���D�A�b�ʚ�?7�llG���xw��H����g#վn�=M{�o�f�X�S��l�5�P�6=�P������]2:{H��ʛ��6��=������1}2������=�q��������gª=�U���>9��D^�l�k�'���̡�o�(?orkE�	�M�9�lG��{���kh�/�A|�jȚ���k��{���m�.�e�[����Svd�x�9�鱞��J��Y��zd�=���>۩k�(�������/����΄�N�z�"�sx$����d�.�����;�w~Cb9��²7ג8g��l=�Џ�\N]x��^�O�w�[��<�]fx��\K��c��x�c"b�N�����n�+κ<��x��ϡ�m�^�á1;<�޾5���Z[�(�=�zQ�Ƚ����^��]����ź�����A[�
����R;�P�~��t�R��(.e2������Ӂn"��'
�v�L����4��&u�9흗IZ
�HQ�&D��%��M-v,
i���Q�v�XN Nu:���EDlF�����a16��e��.�f��ަ�W�\A�v���p���q~L�~�p��3���u�8-��V�:���瞑������o�z�`�c�3q��\��Ϛ9�ѧ��B3��s�"����(�4�m���u3����G8��d 2�SR{�u#=8�s�v�����1Z���錌d�
��b��ȋ�Ha̿M�.)�������M�G�50�)<�fG�5�x؟��ψu����[ ��P�hy\5�ɕ�ʤ�����{�N����{�FE�r+!��p�:t|hO�(�+��fz}�# lL�Ut�#'��3;�j����-L�Q�#>��,]y-���z����w�#����S��A���dn�[6}]h���1�@��T�������B��RW�;�6#b=\s�w���}���K���4���V����Ql���"�$_�cY	��;P�wldgt~b��{k/&˸�ٰQ�V.3��<������x�*�B� B��3~���M�J��wv5�g�^z/���R�r]��nY뺟Bn����L�k3oە"�S �8���T43.Ȼ�|���{鸫gZ}'Z�tT�Ik��9�j�.o�6n%��}��o��_�vD��:�KI�e{��-�Zv���y%��:�#Z�pq��:���Kti]>#�L���T�+vdZs�e�t��':�x�f�q�n_3�!���Rf��c�ef(�"�=�e���<F5㞗�WAk��������$z��E���(���=.�3����Q�%IO�zQ\;B1��d��{�~�C~����7�nh�v\����n�h������E(�Y�.�U���WI�,�{~��Y~ �i�dő�B��~�^��,ȥ���@NQN��Pkk����V�?���S�G�C(l�W��V�n3��=;��}#Y髒���^����o��Ϣ���;��Y�4�T+%��.�n�fu����K�����}~��7/o��,PP�܉�Y��L-�v��߽�js��s�?
�����~�@n����E{u�j�b+�zg�*�2}���	d/z��JZ���V��_�ݍ	v�&�=��o�A�ι�~�^�O��"����b�)D���j"O��7Ƈ��~���U�^���b��0呼�\���{�ԫ;��t���3_I냟E�?W�e�0a㼛�i��*��7�!�	�ளt�5��y,֘^�!�	���ϥR�rr�߆߽jk#��SӰ��4���63}<g#�pGN���Mx��ڪl]�c��,��n��JZ��uƓs�Y���ˎ;����oR�)���*�^�G]�|T��&/��`�i�#-m���OBym>���:�ˬp>� Ĵ��r�=�2�]�k�m����<˕���p��Y�y�0%�s��Ӌ7���}���췘�=���+�L�%�Bv �[�S����Z�f��J�971,��.<"�F=�*�O?Z {�q\z�qN@c~Bb[�@��F��,2=�n'�r&W�]���Fϑ�C�Gyh�9�~x�c�������-��F;������Kg�'�$4':�J�"�G��n�~�0�MN����ï���Nj8���3�����̟k�.��A����9�=U�U-f��Ho��ѓ���7-��22�d{_�e�]?C#��̟o����s�=ֳ.ϽL�R.���zG���m)9*�}�K�NGc9��l���܇��1��P��z&�p;��{��_�&�;��C�+FAs�dO_KϮ�ç; �n}�{3g���)Ě�wʻ|{��3{�\�S$,�Μ�{�Z280;�B��^��n��=c;�-�҃����:/ٲ�-|d��d�3�߰������'��hڜ��n�qS� T=<���ec��z�喷�Ay�����Z���sX')z׽B�Q�4��fV��qO!�	����˪��+�?Τ��ɅY����y�8tc��V˃3���kx�I����l=�[xi@�6��}�D��dZ��ڈ�sEeM�ݝIwr�O��eޡ�F���t֨���cwQ�u�)@���ѳ��r�]��L�����on4�wR�A��kJ�RZ$t��Q�&��Uԧ�����
- t2�Zr����܃&�+��m�Zm�kX[�|oMk"�h3��m1ƢBf�V�b$b|)�V$�]��nK�ż�h���d��A�%syO~�ަ��H�$�6 ��U���NJ�F�*�9���S3�L��)�3�t<Mr�u>�B-Fl�ZƎ��	U��Nb���8�*�gb��s���B��-�S#�����;�u�Zt]Ih��MU���b?�k�M�aK;L��$�(W�*F�N�s4��{�������f��ӼY,q��q��d�}m��lp�]D"5��̸˘N�K����L�m�B�����u�s2��:�ږ��{��3�>(�g
���E[i.<7$��sV�k��$��[V�B��Y�{]2	6�{��;�_>i���풹f��ʽ��K����Y;��1���gh�lt���YRՔCο��yf<B��ͬ�OB�h`�6%Z x�{)����daeY�hY�>�_>��@3�Hڊ��ɮ&+���������7��4���0U��;k�%���R�-b2�4����2:�;�a(���gM�$�Zi��X��M�Go	o8�[�eK�U�b5�$�)��x�;��	 e\P�W��'5q�����VsW��jZݏ��)Q�q{ж�f���W/Gv�tJSw&�r��YA(�ͤ��a9uij�ڹcu<U�	�6�q�ƺ�g'!Z�,E(L�ܼWgw�(��3�������cm��H�av�Wh䱒���x،e �ov�e�mD�-�d�(# q�Gv�Gvہ�m�pʚ�*2%���hZ�m����ظ�
�Ӆ�����!:D7�{�!R�waul92^�nV۹��{�[¯���pv�O�;t+HJ�it�e�.`k	�)mZG�6WH�*% �n��e���(ɕ.M8~ؕ����P�9�Bj�6o%W�M�4��nRU�K�R��WwCX���ݽ�[�L?����fƮ�������K�[-;�*��^D�f
4���Z�R��2��1 ���4pr�F�R3����wp���b�����頻%�j���}����mv���=ѣ�c�m���ۈR�
wh��	��c���w\�{������(����WSbt�c���n��VӴ�E��q�ֺ'PVCv��2�;������H�	P�SӖ����I�����M�s�M���Æ�؈���z3�e�p$ھ�@qh�0nq���I⼵ːcz>c$��1�PtS �J�2���8�#���{n���z��EW ѧ����Z}-�J��^\�.�_��.f��;>��K� ���_^*���VTPĩ��SY[J�+\q�b)�#K\IY���bfX��4��±C[J�+"R�"��b��-�X��e�	P��a�Ԫ��Ym̹h�"*��Uh���[Z�K*6�%q+3(�s)�YYF�)�C�f#qffB�L(�B��2��SDˍq�n[�q��E�e1Z9��8"�ĩ+X��J���TU*,�KM2頦��U�VD�K��[W�2�nV㊸Ȳ�W-��-��3)�df4*(T�11�&f9W31�R��r�"VJ�"���c�h�cm��Ri��´�"ms3��QmaU��R��(��ZG2fYE�W0�cCLh�eKZ�kT�,��X]k5��,D3Z�V�h[B��-���(�s1�F�31�Y\B��FbT�X��T�c�B���kR�4�1&"--V6��Ukt�kQ+PZ�Q����kC�cU�ˋ�V�1�b��i.�r���U&������/��rM�a�3�J��p1�;㻝�|MZ����֋%�Κ�αR�ܰ��A�S��3v�t�eb*��a2�J�p~�?�n7>�7d
'�(��'�~>��xx�g���b��ݮB�
K.�z�S��~�p~�"O:J:	A����]K��!�^Kߤ��#=�<=�cާ�J����}JT�^�lb0T�rӄ���3�h�Ȉ1�W�_����τm.;]|�;�߯�g�z���@:�n�����kJzs�8�95p��:���lNPb� W��HH	����[r�oM⍸�����&��ޏlԚ�{>Lߘ]�c��u�������3�>#�;>ly��Θ�S׵�U��lt׶��x�E&/�\y|�-z��Nî� {޵$w������ :�&e�^��uqG�Nw��CI�;�}ՙ#�=SQ�*n~���W�������g�Rꜻ��&��}R��{9D��Ͼ�]y�:U�jn�#gL���eM��mg�d{����z�����c*}�A�kԋ3-���2��'�C�4kT?gүf�����Z"ҧ�C^�>��B�zU����P��S��脩ğo��hl_H�=�C�n�g_P���soq��-A6����pqzDk�ޮ������V�qʼ�,�Cs�W"�Kxx�o�?{*t�siu��	Mm����on�+�@y:��OJ�N�(6sӕ)�`�q[A�kBGq^�0ٸ�����Z�]�O��u.����ņ^v9`�E	�	�]B��2�я��K�p�OO�Y�:�R���G5�7>>۩k�(��������94U_�
��z���߹�c�Z����s�������?������߲�u�Z��r�;�=���w��,�Ĕ��_���A�9��Ş�ww��~��]yqK<{L�=���tt>�^-G�ԡ���C�#E��UZ���TE���IK����o��կ^�W��
��묮���tr�5׾x�U)�t8vUzv�ʡ�=�ϕoé̬�瞐�/H��2��å�]=�k���[9w��*�8<Y��Ȣ��y8�X{j�Ҧr�\���v��kRyV\��C2��l?[�U�S��i�ۦ3 ��R�4@��Dʧ���
�,�ڿؗ���ͯ�N���/���#������{���9R����8�0�	��=6ؾ��B��#�kJ���b�A�{���ȧN�����6'�f�X�Ͻ��O�F ё�	zb~̧x=�Ԫ����YB\ϢR�#"G�.���ſ,������GD{�8,�w���� Ǯ}~���\t9o�]s/�!]�f�6m���b�s8��6d2si�s	M^�]��r� #�`/�����m�|���i
v�1����xS��e�;B��K������ �}�Yۍ7��<�.��8V[�u-M���˔��:�2���N���3`�I_��~UR4_�O�f�vdD�8a
h2�IP��؍���<���\��gZ��[PG=���=���8��'�nH�P?u��L�ߵC�3ⱴ_:��#mac��|�дZ���5t�Ϡ��ڻ����������㧡�{E��g���k��4j�� ܂��Lz����奮3�;��pO�!�fT�ͻ��
������6��R-S �H�dO����e�M8�ܬf��G*����	~����׎zu��P�~��V}�zd�lK��>˩x����s���We^/d��T�����-�p��Dy���f�=Oوls����F�-��˚�N��{��x1��3��Z��o��t�'G�t�t�/o��-�߸���=�#��C���-x0�ҢEK̝�g��4���Wz��2!��*�S>K��XŃ�Գ�Ѿ��93�����[��*�1@fT����P^���>~��'�ǖr�۷\�6eQU�t�>�,߬��ck�z����`�yi&�S>G�Ȑϭ�_[��طjx��xڜ�Dd`�	`�z$������A�ԃ8��k^<�B�'�W,X�)�w� �7\���@���$�w8����h<��ܾ��P�zr3@��2���4�o����+��Rة��6�N������!�Mzp�}�(X��4#�G�V�����
��7��\
����;&�G*~pRחeA��-O{�%���瞷>~�S�*�)Ϛ۩9D C�����]��qy��"PvG�z�dX���^��{'���C�ݱ���b��ҝm�x�R�E�fL����X���� uNf���]Su�չt�C�y7�<��C����:(�=��s�Уț��Oޫ�=�#$x_��V)��J�"�B@�|}��6��SY��)��s<'cn��~s���׬{ޡ�{�p�=L��L�!��|��ə��C�o�n��	'.�c���;�+�yn���޴����=�Q�=��E����\1A�3�^�ax˭�R���9����xŕ5���L��n\z�hlxWO�Ͻ�Y����"��U�%���VA������ٔ���>��}c,y��r�CNn&��3�����L����7��r62~>����cdi�ׇ�
}��0*ٸ�o��7-0l$׻#���(k�P^��d��d)�γ�3^=W��t��\C�AU��rr}[>��l�M�6���r����b�S�ZdJ���E������C3RR������~���uy�n�COl�N �m�Tgj��G=�1*ɘ��#:�Ɠ�V%�JڜP�c�_*d����]�� U�n���Y��7A���cF��V���(��3�rd��om<�A�7����gr�}�r��C�U8�9��v#�+F|G�W�g�����p�Ŏ�x۟O�ǒ�$��$���,.�-�뜟Gz������|}y!dx�NK̪��p`wd@�^��������f|�;0J�{ө^4{+�Fz�37�kY��w�27�;,-��c4�v�Y%�8���2/L~�}J�E��x�Ԕ��m:�=���=~���X��kޡ���yٕ�g�*��8�2�N৙��{ʼ��Uv��N�Ԫ��S���5藑=���/��C�u�q��,�,����K����w,G�����%�~a(=m/ܪ? ��3��{'���у�����앋t�w�ڿH�}�B[�C>ah�20Аo��|%Z����\_��ص�����iʜΛ��� qV\��R����c���t��\���g�q��.wNn�Ǉ��C|J�쾍����Cvג[��K�N��T�{>}^@�<�pYG�������؜��11%X�q>�]�p�"�¨�����0= x��\41�,�ϣ��u�_�=�Z�G��Rr=v��S���+�ɞ�K)hg_����&<��j&<��PgA��2�E�Y�Gp�� Բ@�s"����K�ܺwF��o{s�o���ܤ��Av�'���W�6$�1�uC8q�z���p��w{	�n�U��D�}�i�4����_Y��N|�����s���-��1�z8�C�2�xz��7jF}!�P�hd2���~�ǀ�=��F�F?{��t�^�Ѵ�f�u}�l�jAOx��wѯt���!x&T���z��<���g�˞Ɂ��z�ex�	�lϡ�0&�����@���{7N���ߩp����	���c+���p)7������V(z��'�����5��q;P�`��k��c�߈�+��qʸ^�FOYE.��n�\���q:�U���� �G������H�5���C0;�+��_��X�U��og{�O���e$�ɜ�ٹ�N��k�+�T�l.��[�KB?�q9�t�i�~��b���O1�����@��p6!~�_�C��5���:��ˊY��d��� ny���A�e�x��G�H�s価���h��$7��J\�t���'�����!+bѢ{�\-+�!�֦^��G4g��9��T���~E��N�:��3N�Ɛ�s*9ߤU�f�E�����yEq���=�x-��,�;�##���<X)�܊!��:;�3���ٴ�G�	���1Oר���������V��к͝(�R� �į�)�7i,�W�t�k�������<���^<�N�LX��o���Ď�3{ןJ���J�m)��e�ok]�ɏ�9�g�i�;-��9A�}�L0���A���ժ��1cWe���I�����r'!�����?�֧ɅZ6v�.&L!�����_c^TK��so��J�*w�|�/�����L8>�쯼f���4'ܣ��>#~w֥��-� Lq�/uǪ1@}���t�⇡D����X�!,��`�[g"��o=�|�y���3|�Og�����o��E�vufǯd�xWy~u3$Е3פ��Y�%����+=~Ćê�G��LiO�-��9����̢�3}R���uRQ2�g��ّ�H~
wa
h2�IN�����Ǔ�]������{��G����
�菄�ܑƠ~�|�ב�j���Y�{W��`z�̽x��U�W�u��C�o�w���}U��x\tK�QJC�҂U߮��h�/̻u�r����t�����Y�ǕeS��'�}9��̩ϛw����|�Sq-n����9��#�'�O�n��Q^ĥ�j;}�v�vS`ޓ��ƼsӰ��(g��s>����L��usg�u"8�2]9��;��4&��՛H{@�Hs�2Vϲ���G��*��r�~�Cb9��}C#}��x�☕���I���\���k0P��y5�e��0���^B^p2�[�K�.y �(ݳ���Jw�'\j��fNS3қ�i�M��<��3RAc�,�ze��p9�=����^QR��]����;7�ɉ<��l[X�[�_��������nC�HBt9]�OWKϢ��=��� �!�?�b�����B�}��!�|����=9�麏f�O2Ͼ�M�-�\*'O�W)|��{V�-
���j���+s.�;k��}}�"�;4��JC�t��{�~���'��g!�P��8.�M���9��J,:o�d�Ofi{��F�sY�^���nf�<R')�FŻL*t�xxڞYTA�,�P�U�"w�_����q��n��n�����_��Ǌ�|�$�ϥ�O{�'>�i{�{=n|�v��]e�mmԞ�=�V�%ы7�Ȼ͏�>�/�W�ϴ�9�q���9>�p����L�5NOJm{a��I���߰n����~bPd���%�5>W"ꛯN�ܺc"ۼ�ƞx������Sd)�l������#V�xE��wKvW�Q_W��s�na�6��ΩH���3��o�o޵5�c�ߦl`5~�X���ye^�d�G��=�C��z�Vy����ma�6N�&s��򭷇Hkd���ه/2��L���+�w�9S�;��>o��=�D�w�(�W�+�b�LKw4@���^�m�O�E�JJK1GXU9K^���0���'aͽ�mӷӸfV���#Cgm<��(l4��v#��<��
9EG��56�������&��7�8
Y�U�;z�OgT�n	"�%M�q���������Ż���q��=c#�۹�T�v�R2Y;�P������<�]L\7�2�I���σ����]>#�����o�*��z�3h_$`�Q>&�w=���|=Bj����v����&���ɬ���jG���3'�kfVd�MO|���=��՟\�:�� ��l�k����^�A�Q{�=�CW~��;�\�G\��Ǘ|��M�zg�����|��T.G���NNO�g�t�t�c9��l��.oL)��ʠ^3Y佼������6��C�=\a�;A�Z2�
4CQ���׸t��d��]'N��k��9��v�=s~G3d��w山��+�Ϫ��^zKP�>��~ʠ�����\��f&}�5�zz��+��|/o�v�S3q�g�]߰��;,-.�x�hڜ�۩܅L�������}�ĞHz8��Ƚ��.���_�f�sX'>��^����yV��+b<�)�Dx�=�8�k�����'���@pƖ�uTuO�dgݔ�\��J��lJ�N�0NF�C��f��_�KG0z5z:���L\D��.����K�*�����~���`���z��~co�t��,~ܫ�2�t�">�2���ծ�nj���V�z�.]͞~���tR������}���z�Qgc��|8�f!@ƍ��죕��v/.��ЉMN�dC�Վl��q-���r<����\-�{2Euu�9tCO�2�}�ⶃ�:�ѿ���:^b/�#�a��V
`��3���jp�]!~K����~�w�]+Z���Dڞ�CS�s�6<{�#�~u��S<�����ל���f����G�=�>�V������ܸ��i隗Oײ|�����c��u���{#���bbJ��t���J��TѤ�K����0!n���C�ȼ��j�6��{�g�zꧽ�4wĲ�>�	�cj���Aף�fxՏP��)�22C#ۿ!p��T���66=U�{�ëd"IJ�}۝sz|bO�ٛ�L��xUǪ�sB���@4&���Syt���!x(eM�m_�d�1���9)5��7נp���</�o�X�����ԁ�J������.M>1��s�����>����ew	�G�̡��
�^�>ߥ�t\�
K ��C95��ٺ�y4�i���}��s,���eR����t��Oٕ:�Rꗽ^�"<��'��E�� �'j.�z��Tg�ڨ�ZB�J<�E�/��a�d5�g������N��lG?\�V}����!{�'"�2���~/y~b ?��J_��W}���wv��Wq	m��I��I��O9�M����.K�sg]=B�w�1���t��a�Dgt��F��|���>u�	y����k�.����zի��>Svc��DݹCݱՄ%Ř� ��|qB禎ݤ�W(�ލ쁚:�݃u5n>�ئ��j�w�]��Ė�C#��	V ��\Z�cH͋�ޗ�?^�N����;�VTP��B�;�wr�_sb���`�y�8Wv��iZ��rhY�F��3gXW\��řx�ϩ�n6l�N:6Ny],��E�8;`�l��h��R�����s4��2��s��B�)F
׸NR�s��x
dG�LHA�ohI�:��F���ow����̨�N�X�M��f�K���
:E!���AQ̣guTA�J��ա[2����7\�!���ƬId�ڛ���g78��b��S�����D�����`�Z'��%q�o+ xS���f�\��qR'$'t��\����v9b���e�0mF�����
�W�Q'�em=��ol���j��2f�g�[�jp�/��E��|�V�rTǨc�i���ok��W��1L����r��k{�Jׯ�S3[���s��&ҽk���g=r�6Ly+Z���:n'���v+$ޙ�����"�9�LŶ��p��C�R�Q�j�9P-�]���G�r{%-(��4-���t�(p��ћ�9�؅���B哥&�V���c�I������P�HZk3�$��h
z��M{����ր�Ij���93��Ǣ��Ъ��׃�뫣]o��* ־`�f����,���2-���܋��C�ͣ���]s���T8�깲�]�Dh�X)�l\*��l��3�>�d��k�����S����<�*�^�n�u�ӻ����E�B;�!������fn��Q�q������>�.Ǩݕ���]�`�H��
M�6Q�������*�� �#h1C���Y�X�r\�r���I)���t�cUa)�Z˷���n�Ȳ���5�Z}��<� nw�w�l��ţG2��6�(�|#�r�Υ5r<%jɹZ��68r��3T7���'707����W/O7y�n���c[r""Bh��l嬰9Ti�dq��S�k�Y�Ɣ"j�L�be%O�:�"j���v�!�gg@�Қ�-���1�4]��ۮ����z�������eN}SB�v�sԎh&��qss��aYq�ŻM�LNI;��k`�yI�'��-��R��T�3Ff�aU��
둹"G�B}gH��N��Ș�˄��d̵c�[�Mփ��_;�1;˄.�nC���f�e�2V����z[]�t�P���7ƛ�a���I5����j���L���EF�B�m%�C:��z8�`$2��Jf+̕7L�]�őnR��4PrM0��]��DH����ǅa���+F��)QT�խhUQ�2��q��7,mZ#R��[��P�,��X���������&"*n`f�����-d+�33*\�+,Xی��*V�-Ƴ-kZfS��:�X�r��R�)mY33*b���a��l��,+�*�[�#��j*��FF*���[Tm��E�.Z���4�a�RV[e�-IQ���R�V��QeuJi4e�
�%(�*��Z��LfZ���6�+FVQ%T��u��D�mF�A�JZZ�j�Lբ9�,�Ъ(�m�Dj"��[j%V���*U�*��B���#lKV��Uk]d1�T�i�0�m(�ԭ,̨fR��m��kZ4����h��lKJ��Q�XfZ�Ym*
1�j�)h1���R�*&Yq���Ŷ�V�j�����U��Ƞ"�6�mmmam�kA-�R�mF���DE��cb5-����J�����L�q�������v�K�D�.6�����Zh�&�jSY�^�+S�7g7����6hDc��DeZ�Y��{ ��#��d뇗��0]{�ᰍ?֯Ң����zO�?<�����cGo"'��y�A-��d�C=��.|m	���LTF�-�4�-s>ߕǓ������*�J�U�E�G;=�k�c��k ���
7j�r�p�� e�����S�S�̛[$st{2]w��.4������#��~m��>���l,%��7\��y�����/�T�m߸μY�פ��urruߤJ�t�W���߭O��C9TÈ�@�C��f��昿a��]ܩ�7S��>��$+�Sl�׹0�$��ӱ�5���>9�c���q�����!:�ӨJOo�)�ϣ��!���9)�%�q^�\R�~��:tw�����|�O(�͉�_\ъ�������Ϗ%�|�z"F �#�3'�qC�5��FHl%�r�Qo�"�=~Ć�:��D/T�4�'�o)�E�熎�����(nI�#ͬ>�I�o���s�5�P��C*Ԡ��>δ������/z=�#�*�ã�G�ȏ{�s�~, �º�D�%yU�0|721Z���m�Ø4倚Bã�m��[����+yN����y�� ����	�,֋��CY������$Ybj�����_&�KNYr+��z2�=.-�9�=ܪ�9��t	�v�*��~�(6�p�Ld].iT:̈����}33�۹�2��4n;)�܉�۽J7�3�Z��$�I�Mg��ǫ���� �x\tM��qJC�{骅쉣�46��w11w���%K����;�M^�~�g��>���Rۯ���73���R`�[��|��^ �n��rA���v�\Sw�7�����rx����Q�s>�������us��g�$h[�/�r�w}ꐆ �#d���e�����L� P|;o.Oوo��s>�6b�{�-�H1ϕo�K&Aj���]��.}�Yƽ!���Y���kӪ��~{G�^՚s;�졞�y�݀=��5�G�dRϽ�8�f���ū�K��5��m
������ޥ{�\�oy�,Τyq���� ϡݿo�u�ς����Y�F}۷\1v
��<���o��9����|�X��T/,�}s<w螵3p�ؤNR/��i��[�<FǼmNG-�##�K��m��sw�0���=��r���L���w>����	�i{�{=n|�ي}+b�)-!�ř�1\&m]8��S�ZO�w�e K�ǲ�y9N&��^d=������߼r�Lz�������Wj�2�
R�~���J�3�:�%k�:�N̘��w^�� &�����݈vT�^�Aa���O��yix��<i�0�=��P0��Mw5lo�AGfiúI��k�AIt*w׽[��7 ����}Q�ûR�[ä\�J���w"��I��[kU�&	��Z��l�����9c������l7O�.���mL.us\��;�Ώ:yb�ɡ}�{�ۍIOxh�=t<�\>��~�!����*�S���R�D�������_��
g�zM�F�{f��➝�L��j,����V��Ṡ8�k���;����	l�ي17���о��c=�I�E'u�����gإNǯ�龜zO}�Z d{��Ddz�qWPb�	�o�0���feM[���5�*Y|�ǞD2�I��o��G�ր�ǅt���fg>��"��1�N
��*ys��&�ʪ�H���К�f�c,2:��9�8��P�{֤{|/�2|�k�
(h]]�8�����xܡ02�~"��z�[��3�ʙ׻#���(py�Q��۵�!����V�CГ���]�a�mP��C
� m99����g��M�d<���v;�.ksW_9������/�}�K1��Pq�D�~���{Eh�<�چ����y^��j�Μ��u���v��l�7n^A�͟Ju㐾���g�r��n[ݺќ�*��&J�]��q>���[��50=u�~CiV5��qԂ���m��E��r���M�,��\�%Ƅ�DW��ې�V+�)Y.�Qq�t�,tkf��n�X&A�J4���~Ǵ"�c�)��}�Ub�dN]m��9��|��];i�J�Dv>�"�lM��/��Xa�?|3ج.�M���o�zu�������'�ߚ6�;v�tF&����u�����ǰ�
��w�۾.���O[���X��kޡ^��Q�+�����0:.��(Iu�y>x�2�5�R���!�}Di�s?�o�^�y=���t�<e�EOd������r�5H�+�E���~�3�s�U�� �T��Te��U�Pm�ӧޫ�q��/�M5�6�)<��G������q~�o��E�<m��N!̆;�s�9��Z��e[��1��w��ݳ�q:c�:�l�~���>�=�C×��<u���z,;�_ϖ
u��5��H_����&X}��{��oԟ���t�G��0�����5�޿\yD�
�3[��f7����Ǧ%g�G�jV�����\43�|�/=~Z���!��zԐ2=޺��t<�p��-Y��*��q2�W�t$7FDK#ؐ�hd2���l?Uq��z*F�"�*����#����Bn�gγ®Pm]60T�jn�#gx�^ʛ�Q���l��S�\���*1X�=8��ǵ���R�p�B8���t�(2y��?IW��G&Jg|[�-e��H�j`���mN��a�eh�(b%'�Sv���ԕnM�ǜ�8m:��з�L���\�J���7��#�n�|��l;��c z��gq�������|��W��w�S��,N�o�b���s��\-�&��q�9���q�z��C�̡��
��z$�~�q�G�P� ��C0=���&�{e�ln�[��7��G���rp�Η:��*s_�]V{��r<��'>>۩� �O�!�^�����r��������d,�G�D��8{7=)�x��?\�Vo�$p�W<���C����V��	{���yX\3��q>.�T����Sn.��gb�K��p��Ҽ�U�l�k�qP�ݥ2k��x#M�Eq{�}����k�8v@z(z�^}{vF@�^���Wy\xI��F����|v���<�h�0SW}���,��8q�%�,%����p3~��Sޓ��d�w������Mz�Lvّ��xzF߭�-�k#���X�����`�	d
s�(�<��|cUL��*�;�T&P�A�rBߤ��ȝ���.�ny���w�S宯��kn�� NTL���v^{xUs��9Ĕ=G�W�NE�3�no�^���>�t�G�׼;Ƅ����9��,�?L�uR��g����`��I8
y+�`��oy�)f��d�91ٔ=�0�z�O��;$�a�M�U��*��e��l�t����I�=��Y�~�uj`��9�FP ��x��v��58�Էz�b�g&��N��c��e����9����� 6*L�Q�M��s"�3��[�~�|�y�؏��8���B4��6z:
=x���&��C��*����n�#>��K��O����$8��䢪�l`}�
��><5�{�8,�{*z�V�t:�_РI
�g�ё��B���\_�S�͡w�Ɯ�ZV��K�z�?^�^O�|A��C+���G�x�!����lMP^Ur��KW������3ϊ��|�zV2�IϛY�s��c��������x�*Ч@�MT/`~fi���E^)�6�x����c#r��ZT�����N}�2��^�½2}�dtͿnT���<�NӟR£
;tl��$K������e&�9����sӱ��k�������o��a{_���3�~�F�z!W�7��6Y:�VE���L�!�S# ㎽>�������<���l-ff��8[��ݶ����ˋ�<_���=]/"/o����-�߸���L�Ё���39��'��X��^��Dj~�^�� ,���=8�`�<:�*�?�z�^}u�4'ދ����ch��L�mi�HjU�5*QT�l�$	q���-��-0�Uʂ�ՏF��D�q��4�q���~Ī%x[�p5lO[���b��+�GF�Y�.��.�
D9����/7M�HKge^�+{R{&�.�ǰ>	�{Zq°���5��=�3�ۙ�k#ҝ���G_��-~��;Y�GfUp��*��M�y��'��:��6}�0Y��-�����jD��^9n�
�)��6�#��<�\ut��K�����1O;��08��Pt\
w�wh�L���ϥ�O{�'��Q�����f)������=�@>��Q+����[u/"1`C#� [��/��l���nΙn�����C�����U����9��nG�Y�[v�o��K��td n����\<��n�;�.�ȶ�&��O�o�>'��8��5A���(�,�w�{��.qþlx\��k��n��R&3�߅ĉ�^]'n�En�6=��nk���͟cC��pY�dWe�1�q`1��W�}�\c�
�9�u�>4� ��	�&�a�r��}�T�z��������h��{��DdG��p�3Ǣ���&r�fg�a����h���C�B����L�~x�c��@{|+��{ޮ��5���\��*U�*�U{$T��hMW���}a�ן��3����z�D{޵#��ϙ��&�V	�^��v��0Ā3��!A�P�K b�.gh�=��uzvޞ�Q�-�!u<GH�ؽn��]Y�-��QC���U"��N"$�"SJŠTy�����1(n�T�/N��\�e�]M2F��Ĕ`h�Fm�8�oe��%K���2W���f�[�p�<0�|O�T��]�o�1�n��Z�d{{����j�y哋�K�����W��N��rO\���$G�Sq�
\����V�����S�98��R�M�=��u���܏o���B7���C=��9��v>�X8� �'jȞ���Exx�]���U{����sɎ�Dvu���ܼ��fϧS�-����}גG�`a��-B����;޸�p]��~���e!��xB��&�]#z9g�g���*߰�؏;,"��x3�ez�Y��]Ј����x�;�;�� ;�G�XJ�����]? �z���˚�8�ֽ�~�>U��c���Y�������=�r9V�9��<� �*�TB���|��^�qޯ l��Vϲ�_�|g|�n��y�/��~����HǙ�BZ�C3���<�:;�u�K�h�^�(�m�]��TJG�X�����-�����W�cE1�hH7��D� ���s۰�.)m�Wx��{�}�.�V����zL�O�θ�#�y:���=� /����oS'�A6�)�⢺Xn��+K}^+���`�+{4��x�r�F�`;۷�;��Kj5cIY�@�o�HjL�/_d]9��r���+��G��Q�� Ĥzs-�R���odR�hh��n]c�٨��F��ި'd��O%KGw��x��8�t�_<|P���7�M�\U,��t�tԸv��;�o�.��g�������/ޙ
�K����Gq�a�ē�&�y�ex,SP�l�d^G��T뮿 {޵$
��-w���E�LO����J����V�̷S�'"��#$2=���T������Egtɪ��fk����;��H�|��}��� �6��$�:e�F�#���"��~��D��Mo�z��]�}�y�T2!������Wxk�6�q)ѬP��J�����؉���^������-XY��/�����dyz���e�m����I�˸�^�@ZN�3Ӟ��S���qF����m(gDz�9ӱ��{ߤ���t�O�u+_�]VG�^�<��' �n�w�r�u���gU�({@�B��p�dE��
�#���'�/�b����>���=�9G=��͑�-L��q',Ȏ/��{�֟[���%�7LT}���,���v�����kf�9��v]v�"L�#�7�z�-��rh~�#�����a��yD��!o��1k��ޫ��a&�">�EE���\�����~{\���RrgܫVq��r[g�p f�騐D�4mR��&��RK������*f拋��kKI�buX�dWBB�WՑ�/�����|:���κ�:�.�W�V�7r'�GK�,d,���R�wM��*',�(`>���3��Q�[��s��A�%^��Bh�_eY.��V}�g���W�i���c[��zק�x:s+"y�7K��_��-�����##��s�?@�:�e�-��x{�� N��Ʈ*|Ps��2+��j�gӮ܉ȅ���k����S宯�����>���"��U4Q��#;��p �Tw��+����9���ܘ{}����xv�؟��ψ1���y��>�^�>��E� �T8���p�"�9&��x�3�x��lG�:!3�>���ҹm�xMp�{���G����Č۩�*����n�#"Cad.���ſ,�{�^����.�#���e\��yUi�^��d{��=���)�!��HWU3��ȉ~
q�vOO&e��K	U���K�̏w��N�m�q��c�v�}�dQϽw�R�j��D��VG�꽕�%�Ysʋ&������+��V'�7�R�6����=�����;�R������U�U��8Y+{kI����ݛ�I��e`�)�	����y�˜_��G���� !	'� �$��@BI`I?� !	'� BI�0 �$�� ���� �$�� BI�� �$�� !	'!! I?�!		&@�z@�$ �$�Ԁ��� !$�� �$���H BO`I?��d�Mf���@
�f�A@��̟\�#o�5�P�Ql(	Ukl�4�J��Q*��
��RA��P�.�5f��*��iE���(�������ى%Kl�Pͭ�,H_s\k	��V[,�R�C�e-�-i�(�n���U�֔�h�kd���ٵiZ�{���liIY�%�[3T�4�[[JK+l�)���m�[%�idM��Zұd�[m��[B�m�6�R�j�2�ҵD�E]n�¥4�mjm��R֋*�U�t{�%���b�j�1+�i��W�   ��}e|�����(y]���sAҽ�Z��V�I[���@]�ˮ t��A��@u��S��43�۔j�l�NR&�3Tћb��VV��u�  ��঴Qj�� �\�E+�x��h���<0 (��(���x��(��(��-�� EE��� E ��x 
 ( �����  罴+5��m���Z�e�����  �� =b�j+��Y�v�bc��Z �Su�C��EX�8 U��t(�+04�WL�	�S�%6m��5Cc����  �@ѽ�X WU��� .���u6�'9��s�[�ǆ��@ջ�V�zzP��qT�=;���h ��K��iZ�w�-a��U	�Q[e��3�  ��/���z�hz�� m{�敶���N�g�B�{�ZmU�r� ޒ�VM G��T(=-��� �3�t��躽e�[J[=�9���k�lwg�  ���j�����憵B�A�( nq�{�J�:�:��҇�Y^۴�[5ZN,�=.��5���j�-i��
tW�y��{b�m���t�ckb�[M�e�����w� ��º�t%]�ڸ Уm;��4�OMi�=��C�,��� Cz��usݻR��׭�g#;�޽5����ζ�{� v���
L{�@3�Yj�D�2����  �x4�Un�[P}45�f��䝴���wp�S^`a�)-)l�`t-X4�]��d���]
�w]��5�-��΀ �c����T6�kk+-�������  y��u�hn�Ҵ�:7{G �Y[�ծ(� ��Jz
k^��8������]�����k�,P+��]@�����^��CQze��m��������   ��Y &��t4[69���t)���٫�l��:]��]��J9K=u��Aб�޻[�A��Jj�����]`bM:��| j����IJ� )�IIR�	� ��������ԙ 2)� �Jz�  �{ҘU4�# �H�2�j(�C�?�����^�xG4�߱61��٦��R���fk���u����~�����$���BH@�a$ ؄��$��$�	'�!$ IH@$$>���?��g������wF��p���f��\i^ ��&ڀ,i�Y������m��BI��o>U�ϝ�t���i��C�;�xw1����8���p>� c̐'���2�l�T�VmܻY���|&�;ceޱ��5Y��݇u ��:�e��ed5u�� f�"ӻ��'fkX�`h˄2FVh�+@��)|��*CcLS��N��jzv�^3�4�eܚ �)ů綫TtZ�����L1y�v�f�`��6
˕<�����I�VjzF���x	e�/ �]�J�v�DL��KnƬsjX�V|~W7v�*miu�3RE� j:"�L��Fˍ^A��	�̀�QV�@7m����JD-t�;ݱod�w��м�bf���C(��yNOi��#Y�k�: �����n�Y��"��I Թ�[��Y�r��.��p�2��m���fn�Dї�ػR��]9�5�̉͡��I{�[ҚS�+[S^4h��QQ�(=i�.P.c��Jאb$�jGfLf5�2��S��4R��H��h<&�wuM��A裘�F�D�V�
*�iS��eZGcl���U�[JԔ���k:�	577T1lq���widT�n��Y���w)]$h��gj@&dxڻ6짘N
Ԕ�ĐM��G	�)�!�,��>N�4���GwH�`齤u+�ַV���x�+9�!��9wJL�2�h�/h}(:�FZ0�d;���1R*�D�{1��j�&�Z�`�[L��h<^:�\LƦRB��]H�c��!�H���;҉�ї�N�W��+b�k���w��r��H��v,����ʵ��45xꛧS�,�*eڬۉҶ"�6��GJB\�n�lS+CPf̩��(��4�L�C��*�f�Q��ܸ�aݬޝB����6%k�Ay*5�3jU�(�)ͻa� )�1�qhfU��w`D�����S��2�!-P��չ0��qP���w�J�϶�6᭭Uu��SD�����j�d��V^U�4Ul&eKz�n;dz��c��KU4�P��2�o49�byA�mԙ1�z7A{Vn���#�*X��Ϟl���|�[0�H֭fB�)�p��L�ބ$A����~��R%)V���B��j�+2�(nB���B�j������n��N�M�F.Q�%��m�0�߆ZX���J�1����3L[w}>�Sp����B�f ]�V�9A�1Oq}A4lEwS(+
�X��U�,��YbR��3�j��U{�Z~�ɖI��x�Ӵ�f	W3I�:�؟+L&�)�*W>�3SY�5���f�C�N�[�v�'[e���e���2Qz d���*J�[{������ۼn��jV�R&�
㺺 ]4hTd���C,�xH�SҨ�$�2�v���Yʻ���x�g|�~x35芋�_o�+lx�fe���i����J���'Q�9���a��˱i�C�![��[{,=/m�#m����u=�e;���Pո�2�H*H\�Ƚ��׬��̗Am�3 �d ݒ6$��sfɥP/R:ƛxd�	��3�R҈en(�YWh7D��ݽŸ���$�Ok,�jv��g3���4��:&c�V�X��݈p����f]A��-�.G�e6fؙ2�9z�m)�y�HTi]���={3*� �A���rB��e�i�����^nY��CE�P���K�r[�d�vأk-S��S�0����kW5 ��T��GY�q��g	Ӏ��ס㗠|1�#�����y燷91�v�n��*-Z孕��^ƦdcQ��6���`P�M�Rm�05Y��z]�N�������L��5Q�3�7��#6��w�d�����
12Q����t6�I��d%
�KI��Is\���Vwi�(X%B�-C vE�����%̡��
��5"e]-N�,�Q�e=�y�VT%�Jr��V�F�$��V/0S�k߈V��2�%	M�%�hD����V�2!�,��b۔66rc�E+�PѰ˵��^�YBT�^T9CU,�-�I�kkZ�+cH
8�i�!t�Ż:��vV�Q�Bc�[���rv]�32�ָ��`�E���QR2X��@-nO��l�ǐu��r�%&c����L�A�1d��
hj��c	k�*��6U��JY�7W�.l;YZ�(��e���U�Q�w�2q]�)]!y6l
ܬF�˲�9T6Q���w�S�ع[�0f"�.9��K�Q�#4o�uwkg^��x��+le̕v��z�X����>����+S5f�;s��2��ok�l��@�cq����k�k/�$^�,cT�Zn���@]�/��(P�-j�R�&��O���q�CY°�����}���	�ϕ� ��V�H�V.Ρe㡻��TP�&f�?�5�[pM�X3"i|Fy�v<���㡙Je+� ZĶ��G[��C�]6�1��t���-x�Y�4JȀ����t�@�����v��WIÒPMS�(ԛ5�T7C�J��8�)�xS��b�ȴ������J쓠��v�cĎ��R���܁���l�hIe��9�5�&�bO	'1̌՛���+v��(I��Z%zf���6 �i�t�Cuj����g���2Z�B�*<; �B�P!�����p�ml;u���Q�0�"X���7A���y.�X��ņ2�nڛ�ܼë	x܅^�#��Q.�j��nG����18��m^@$��v"���Sj�)`�U��q�I�QZ �ܺx�'>x�
�
��h:���Rڻ�o�0��xg�5n�2��PhRϳ�D�SE��j�1,��T@�R���R���5z��Ij�ӆ4
Ә)	*�N�mى7r�r@p�@��Af��[Sl�!RѶ����ƷJ^Ah#��%i���q�t�N�b�X�弛X��TXl`3�mV�IM�fR
��+ ��^�P?�d8�3N���kn���$B�1��*�{bB)����E[��0�[P��-(�(�+c���>p,] ��ݣ�,�m��NS+!6�*V��x�:��i6(�Ԏ՜#jeD�H�&Q�c$�i:#5m�k#�u%[�{x`��m�b�A ��K_���������"ԫ	��=���/ ��)Zm�7Ğ�L�.<X�(���e�łˤ
��'��~U65�ٗ>7�L � P��2d���ވ��+�t�ǯUې���m�m-ݰ��SN*1 w��75�Q�l���*D����a�m0m���lӢ��oM�F(�^c�ǤȕK��� Zl�Q#ۏ�u�m��n7*�n��K.ҫyl�V��X�ک��a;w��U�D��ݬ.¦,���;sq��VJt�쥚Y���$'`b��f�ɕp��k8�� �AQ��"�,�H7�tn6]j���+tG��Rw��P˱6�՘KE<��V*��\Hk���h�6�vvTu/F����۷����l�SCj����Gt�m7j�XWeh�w$$��3#��l���W�fh�ws{Ա*����)�� �zq�/�IL'�6��L����cn���ɪ���/���H��E�
a�V���&��+У,���u�L���Š]�A��#�$��$����%D!���@��fا����Y�l��;�8J��Ud�f�����*�V�Ya-��٭ɹ%�t`�m�׫VC0�����/�^�KU5�kL�*Jү]�[et�)�
������࠮�xn�	�Z�e�f��oxl�N-�{����8ZY�c��R��*�]�ZR!-Z�̨�M	��:f�ޜ���nvHǃ���L�*f�L�m5��Aţ�&mυ#�Ց�vKvf�`1�N}�;��4�z��-'V�k��C@��8Q�nk(���ɸ����9�����2�d4Y2Ar�1�.`�jU`,�ݚ���ALd� ��`�!M�V8�����2���@3z���	j��cB�iJKxv�ٚv�A�V7>ݕDe��¦j�\�5ʑ�����-���d٧�ƀ��Y2�(��Z.eh�w$ʶw)fRD���N'fnZg���[@Sbkykg%�45j{�;�vL#n�h]����c�@X�r��ԑ@���Y���QnMF�P��)Z�af�cR�=�O�Nb-�!�/���-�����cN��)E%�Gen�@�g]ݸ�%]�%�� -��;�h�n��[mm�6�Ր%�Rw)Rt�N� :��,�Z�M�*җ�h�}�i-�B�H�F��h�n!����͹����+,;�k[nb��7f3�z�Ԧ��(�Z�����zhɺ��*L�mPeHe�F�%	�s2��i�@Ӗ��ZP����x�Y/i�P�oGs)�!��B���!��l�i��6zFC�����:�
�o3ƓAǫAT̘�4h��ыk+x)�)��W����W�	A��.IB��]n%l�FV����+X7-� -�ګ�`�[��N�aE���ᶥ����!I��tB)vr��nX*ʫÕ�b˦����XuM�����T��SѨ`ڛIS���4--Ne�w("tQ3u]�ZR9A$���⼂��wt��-���'���ġ�ݹ{/��q9�Mb�r�KEkd���|�>�8ia��V��d�yl@��()t��O��*�����B��v���:u�Q�F㴫Dyi���@�%��]˥l/�n<D8ra�b�Rb��P�BP�L틧�%"/%(1e��U�D�n���#�S�������@���P�loɲj��.$��X��L9��6v�!��u$� �KE����ڨU���0S�p �⠰9��T�U�^=��T�)WDlӑ1>
�Kl��^Q���F��	�L�*��)Ab��yz!�*�x����0��T-�FP	�[_l�7�T(B��6�#hmYA[�/+h̭���2�-Q��OF늆��V���]�Vh@�Y�[�7!s%�r���%7��T�iW��d�ɴ��a�g鬙3'�5��c�X����L�vl:�C+#$]��5h��:.��ݠ2���a��=�${��2*-^V�'�7/�h:�^f��x����R��^ �U��ܫ%bN�ML�J�>�.���d���H*�U���c�G4���*�i��M�hV�u{2ee���5D�/k;��d�ɧ��jM��ˉ"2�jo�krX،Dlb�Gs6=3C4X����:۽�m�f��f�}jڷP���Y���B�4o���B�bnF�V[��K�A3��zH�7�� Öl^kk+4�3m����.�.Γx�R�	(��0�wh+��)�AJ���:�2�d��o6�2fl݇,1�3�Ɨb�ݒ�W[L�ޕD���cz�{�� �m��[8U�v�*���n��6����2��. ��LX�;v�6V�CY�$�%�Y�|�Z��7���q:Wq�v���ı�W�����a  �!��7oMP��U����4K�Sb��Ԃ�C\��Fn)�+��Z(�+V���;t�F�H?f�@l.�X�h�{����!�����m�u��j��D!�r��dQ��Z`�a����չs��t�)��4���M����[7H�Y_���F�6��ӺoE�7��7����r�*���@#��i(آ�y��ŭт�@Ƽ�;2$�d�P<>J���4�N`���7Q��PVH�͌leǳFN§m���+�EM�.�`�&��`d�(�(ͦjņn��yu+q�Yu�@OeZ��8�0SS4���a�eࡲU�������l/�T�TPVІ�hK�<��vrZ�u���U�υq��������j��qf�t�oZ6�{�*-2͔��J�h,'5\!�.Ƈq�J=�4�/盶���k��¥��Q1j1�W��m=Z��%��Ekm0�+pĖ�[��m�ӓI���r�.Pn��R�YI\�����#32�C4��t�EM�)oc��<x�<;���Cp��c[O-�
�V��ӯc�>S`ע����l�*�v�L��iŪ��n7���!٦���Ь��Bh�:��7�Ks�1J+C.�R&�ͧ�EA�5�aa��v�hR����v�n�lՍ�#�T��2+,k�4K�{��.�������ncڽ-��Ԭ����f�AY�I%�)X۴G��agr�5�խi�+�\�/BY>���д���P�	ͳ�=�k����aOȪhF��K"�' ����OCՆ��#�`�- Q�LmYN�p"��9[0�@�cr��8[�����,��x�fJR��i�Tsm�è-J�Cr�I0Ue �����z�X���ͅ`B�����z)�e(^�Yx���/i�媰Tm�������!v>ƈ1��˳�`�����e+�v�43
`75�f[��&��pS.�X��P�fe+b�[x��\*M?�kO*f���Fn*d]��l0-�R`�T��s������$֘<f��g�+@<�YY���ǵ*xF^�zը�bL�X�kj�i��μi�f�ILY��0+D[�2�ŌTu�
P&4]<���FJո@y�nd�-Q��=�.Tb��6���M�ka��{d̒��M�?�9Ĝ.>�a&����=j��X�x���o&��oYV�����Q6k��*�#Y.w�4J�ԿYi�fgV��]K{�̂,Ӹ�V-������p��Ӿ�]|���]�uk8�0r�{4���"�����퍏g�<�����E�`ۚ=�������do\�+�T��n�u��S���m��JF��;Fbܓ��FL�\�*<f����(10n�v�p�e�#�C.��9wгB��WK ��� �щ_isu7k�c�����s���r�q�^+F
Z��N܆���=[��F4B@I�v>�b��3��a� ʠ��h�2�.�ճ'�.ԗI�ъ�����],�P�(�w�fy���V�Ggu�hMjĻ�B�|��
�}�[b��,Pڰ�V��a���<�I��������Y���52���.}����X���c �6w�����:�T��^��P�4!v���W����cz���=��	s?�0������ᵭ�����z�XŮZ��IΊ�n�6r�:.ٺ밉Lm��%j��`8�g�����>F�pH�.���'q^�7K/��3hxV�ʐ~���~�h��wœ�to�l̹�^�7|q��b��Guk��u�r�c��������]�ҕ,�˶A�m�Q�*���
��KG_�H��M3�h�+D�_�e?���J"��q�{7�fA3�2��M�uX"JK{L�#lhWVή�B�;+
����U�m���8���\%ō�/�mj~�%�MW��]���(�R�.}ٗэeY�&zߠ��O���N<]w<���(�ټ-�Q�]헔��Xwx�$7:x�ZR��f�%�6�D\C���8�-;�Azԩ
ܙJtnu>wt<|�Kk!����Mk�Gn�R�i��\������2�gOK���V��S}�FM����Lz{�-����ڒ�I]a*�osھ찚D�S�7��Ѐ��'�qf3�wG��Hvn{��뻫<6��t�={Gq�dc!�8�+�'�C
������_��r]��ג�Ѵ%�v�3�s<1v	 �y�&Y(uӲ%l?=V�u(^�}ա��O �N��'6����X�X�F����
^�sj�8-��/EF�S��%z8r�{N��d�ۄ{ø<���1nYr���C ��V�����E��zr�o�d%�uȞ;ͧ�]�<�2+7ك�	�����A�_��� �}�<c�������E���כr�ۊ#�K��z����V5��TB�9��2���y����3�����h���̍i״3��6�A�9q9w�Z �򷱚�A2M���7|�ޔY�R<j������s4r]�7$bE����r�+��r�k�����<#)�Ł�(�8��;�د,Aq���6��G�tr���o0V��]���������-��#R�l���\���cCIe�xU��#�)d�,w4�9��9�g����Z�*j!�lr�+�#�;��7�q�����`.ӤYh�hp�_^\����|H$�=\�)n!�;�c�9�v�\��ͥx�AÖ{uNoXY�U�W�2.�Au/�1t����6���E������8�*>Ic��w#��η�ZE�������h&�*�Z/�oϜ;�l�z��6]�x����\��u�M����n�6�����.�!�(�P΁�	2�j&�/��o��me;���Swp�G-�&LΟq�(ܹ]Zu͙�6-�c��GuY��v�D�m�%!���%S��ެ�����^�t�dV���s���N�[ԺZ�"��K�h�;%:Z�؊M�3YV��wVŜpX�x�,�,�1w �
�[m��[k�Wc�mރy�^�V�OlJ�M�7�3�N����hJ��+|4�CC�k�}����t��΋���7b�����v�z���S�����aH*m;yXe�.z�����/�ۣqҾ���<�����}�h��]��R�E���EC�g��i;ƌ�5�j��-.#�(�Z�]@�a۠�Nwa�k/��SZR����H����3>Ͱ��������~��L�wV�y��Sd�>�U�XiS'��Xkw�Ԉԫ/h���	6�� CF�*��Q�.���@:��0�+vug^1xTxsj0�hwU�6���7K��u^6($m�2�s('���,��O["�To,ש��g�\"+�]ixUى�a;���]n�Ώ�f�\X�>ă���J<�>G����O')��z-6�����}{�S������D"ZbP>�V\��G(��*���Ys�����s�Ulw{�A��� ",�w�w[���E)r����C7�SX� �*VT��Npo:<탣�4]�b�s�AHc�j]7�	�t�LE=���3w!����Џn-^���#���aֳ�ת�ns��yz ]�1�v��68^,C�w}av�q�M�4�9��[��o}��R����UsY�/�/k7���n�
���F���7��4�Z�	�-1uV���kN�:��I/�����b�i�&�G2��.�r���3��}r���]��-�g=���c�r�L�h=��u���Ud�����{ـ��P I���{��NĚ���G{CY�o����<��y��u���u�B����Ik�x��6XW*��rxi�ǷT����@N���R�nz�C]Nn�u�ws_�P�"j,���ԡ�`���$9�y��j��7Y�� �8�Be�M����BՕc+C�m<��S�d�i���K�ί8콦G�N�[���˨��M�NS��-�c�`�����4�{����vP�ۻ�HqOVlJC���,B�@Q[ٚM-h-+r�]�1.�|�m�f��X��a��ƶM��n�����,��Y\���ڔ�d���AGF�uB�njξ.�񳉺aS�h���2���v$��f��i�e7�c�"����cs�2�%mE֭����{[|NPcy�u���~�*5]�H>��ߖ���'�(�Q\��;���k_�,y(�j�*��A��r5�:�%�t!�?{����!�hw��Ǡ5J�L[rKۈǷL\uh� �/3U����
�A����\]�h�W��Ւv����e���+X�7��ӭ�ZSv�$s��S�r0pEZt\�_]����/\�����N������,_O�F�ZK�;O������h ��P��wݶ���@*�2�.�vq�d*�r���|{@Y���`Ko;qOT�=��n1P��5�oF�Y�4-U�bZE��\�5 ���[����qum���R͎L:�u˹`��ղ�a秄r�w8;�P��\m�.��`ѧh�+����!��:�C^�f�On�Fڸ3�˛]}�u�Cz��8�w�6����ڐ�b�7O�i�wk�:@Y�/G%��ŀ]����ܥ^���ai��[�k�T]ojO�OWN�K�<t�;�xq�i��Gv]3$�N��B���y�f^u���!pb;��ik��-���݆'��t�Z,9e�F)�O;����L8K骊�g9����K���=���9�Խ��D@ަfoE0�n=N<��Dɱ��1f�2�"L��ڇp���K\������Q����qv��4OF+%����Q���=�{�n���_a��oHU%3Q�M�wbOՃ���._-3}�u.���S��Y���	yD �<q�5�ykO
�d1pV^Ta\���*��ͧ��0&�8�wigtw�Ou�1�{�H�Ep8Nv����N� ��/��?@��ֽ@���	[�j���ou��T6u��cFu7�bA+���*���v�`�1�`���}���ևj��i�ɴ�eY�g�2���,}�yC
o������y�0W�e�6����+�cw�55��2���SPؚ�3o��d6�޺傱��8|���s���$uЖ&K�U��cKSpM�B�n�]�e�;���R�_C۠��>�{X�~[��ry�e�͋��Gȥj>�z���文,Gj���zQ[�V�,�.���Gu��4јP���Ŝ�J!��޲�����5nr("!�\$�[OX�-褦�5�}� �v��bQ@yn'�j=K6�h�ܨ��^lޣ�O��{g<�LT�Y,��1Gg�U݌VιJ�.r���n�<2<�-�ݐC��c��l=_^3�o��� ͓�;WF6vL2{RBp�y�Qx��쓼�A��v�K�Y�Q|���H��N���G\����]Z����u)צ�M�kM�>����l%��	=�#D�ǳ���7�-���:��.����(y�s1�wLˎy��;��+��樇_N�Fg�h�d���v��W_L��zٳ�u�R*���2��v\��W_,�ê�"�i"��Hޅ�~��j�Ҭ�Z�K�����D���gv����d�qw��ʕ��M��!��#z�F����H�i��p۾&*�W;���v� ƈFg�Δe�����K���pm�l���cs�����l��X�p�x�է�۴��=	BVq�!Ds�\|]����r��k�e�|�Ƿ�W�T�{��/^X�5�wK��WgR;�ݹ@'ch�b+s�A:�ݶ�ծ�Չ6���u�|�p4ʾ����&���q��$��pY�1�S\5����D�]�<��x�g���ٗ�V:v�<�����Q$�	���i���Y�(D�[��Xl㩄�J�h{5e#�z�*Ǫ��Π�������޳����g�S�[��òV��V�)N���}��8�t^ȧ�r+ݡ/�s�z,
��XV�6�U����h��Ll`���^�k7�Y�q+K̩j9����g�]��� Ȑ_f�����6&p0��\b��wJ��^D9v�!�q�6#��W0�{�y�P։��̺&{<K�n��H��Lo��stʋ��G�fzz3���ø���N��܇F��n<<]գt���D#�A�MР���.d�{{PI���vMo*����$ ��� ul�p�!$����吢Ț�z�����||C-c�ۣ��z���7���4o�΄!��<�)���D�*P��O.#d+�V�����ψZ�	c�����ق��}V���� ��v\<&ft�x���|�o6I���l^��U��aL`�B�ɏx;��rԑ�c�Lu�:����x$<�;��n}|�Y0#������R�лlvR5�W9� Z�_
�����\��5���koW5�����]Dnyj"&����#���]�Q���8*͘8$]J���Դ�&n�.��{����wY��ݥ���&%�}or׍8��.І�z�"z]:�]V4��=;�QX��j�Dm}��'7l=dfR�TX��mɌ�}�{�ǝem��츬<�r��;Ӟe/:�훝b�-"��(l�a�i]f�2ѹ|0�[�<j����`�O�ZI;��ì+ƭ�av���l@���%�tV订)�#�������f��
��0��z�3n̅�+��ƿdJ�f]�&�qX�pp��,�e��uA��c@�cc�'>@s�{l�b�ݢ��.ú:i`-ӻ���q^RV��*øg]K�M観V�����̩�� �j$�Um�h���&��B�ޏwk8E��Я��u��G\����� ��o����ɾ��4�H�Ə$��屽`�U�f���cp�8��{vҜl&o�}����{Jb�]N����t:�Cӥ�����|TSj[�4.�!�]�s��C�����UN飮��㑋Ch�:�j�d��A�.#u�n]��2�Rφg%wM����R�p���Һ`Z�Q&M�f�7\���(����yV����������h��y�-��H/\���nL�[�oLW�1�5� a��M�AYh�˩�>��w��4(���ӄ^�|��ʳxkfK0�,�Y;0���Y�0䝢s�im<5�0Y#hƟ�h=���k���yj�$��yh[pX �р�יh�`�5ß}6��}�ޢ�n���"�z����Z��C�\a��c�:7py���ݒ��NA��t�u��v��I�����̚LL��Q���r�S����v�*PХ�*7�S���Zh"���QMV^ed
�ښ0�I�s�+هN�y�8s$8�x��_e[���:|���8�@��z�٪м�'n�]�7)V2:|�X(�4Q�DP����1j�j;�0�Q��yQ���M�������z�-9�+��6@����Y�e���U�gs�
g~oFЙ�����DP�Ŋ7��՘Lm@yi9���50Yᒊn7��eP��T5��I�h���3W��]��w��'p=<�㙺2�W�SC�d��{�1��� �+ �fP��zKE�����C
�J�])̇d�}O ;��vfs>��r	�<�o�j$����O���{�[s֬�Y��x�����R'.2�=B#ue��szY9���M����h� �m�52�YdѺ��C'!�N������j�:\��-�� 2�h��ν;����؛�%�EZ���m�n���t��-�n�8�1����Y��q�6��C}7��w�[œ\`���N,��;����KAduc6a[&�w1�]��=C��@ۜKDs˶�ݏ�ͼ�|��
Wwk��n�x{�4J���#7:�+�;��u���u�`;�[����+a:ﯓ�j.��FeջB
�O���ǧ���k�ѽo�R�뛸�5Oo��f�Ԅ>�tg�lZ��%�1�y���U�r�ܿ�x۶U�q�ew��+��n��,�yY�����w�s�w�7�o��_o�2���Y�}���$�BC�BH@}�ߦ��z��L&��so����x*��!��҉Ҧ���Z�X���]^a- ��[�î��QA�����&Z�̛t�
a�RꍮGZ��E��]��U�VV�n+h�7��Zm����ngV׹})b�ۋv��ϝ�<�2��@�A��K̓�'u6��F)����Zs��ݦ��-�{�O;�H��v��f�\�T�%WOKx*u��A)S�bP���<��r�A���Yj�}��h�5��x40��{��A��q�w���dM�N�t��WdQ�����-.��7�G��+k�|h�(5ܰ#���ֻ�i�zn��/,��Lo�����6��/�MVv���w�f��}���_j�I�ʮ��5�мV#ԥu����kN'S���c��ͥwO0ؒ&�z�`���p���Ti��NɄ����	Y���lY�g1�b7�h�9r3T��>#R�u�� ݜ��L�����9m�4�%Yg�8cy�0t�]짴����e��Od�_t[��4�)ڐoE�1%�{+NaX�1�F��u҄���	7;��L�Q��A}�������-��]=l�����P�8���t�3\��f	YF���_#m�q�vq�,�)	����O�p[[��c토���tL�ы����\��7B�L8�k*��^�K �4G�w�K�^��Dt5@ۢ4Oas�7ٛy��y��`����0��_jaU�@��+�������T'kxS{L��̨�<A���#.�|p�Zn���{�O�2ኼ�]���0���mׇ��]�bu���wӬlxOdu��u�v�Mi��ђC�6C��V�4Ŋ��ھ���@��9Y[g)�R��T���`��	�T��w�۵��a��ۜ���X5zF%K���U��r�e���D\�M�qT���J���6�/O=J��8k��{�`��c;+�� ���Z���t��f���8��2����Ch��F;3ј��z3`⟚=����6���\����<�x<���G;N�s=n@�xǧ�{y]v���jة���7jGM��2_h��׍��p�H�\���.G6�I.���V��V�ӧX��bi�w��Fc{���t	{���tV��C4
wCj�qZ�`�i�\��o��՟f���`��>�v�G�3�8L��y���0�)�)W\���[F�T������4���5�ѱ�%`�r�5Tc9��:�eo3���2޺��ըws�����r.��D�P�w��� �ޠ�ڂV�\6nvʛ�]��1�T��Z,�O�5j���K���u�5?'���4�^��g��T����:f�Vjc���ފ�d��d�]N�y�X�d�p繁S����A���ݢ[�/l�:%�wZ4;�
�+uǛ�N�)M��%��\�������<a[�V�˝��v�b=������;Q;�!YG1Vᐖ��oݱ,����b���u�X��z��܌jY5�HI�D�;!j;���U�WB��ݹ,]���aP�jTZ�'N�
M-�'eR���;eĠ����2�q���p��d��Nv��^i���.�r�ފ��!`�6����]�C�߻̴՜V�Wtv�ճ�)k"�"����K�l��[����f{`�g�=#M��/1X��s��h�G���s�I�K��8c��t=��o{��B�F5!.b���ke�A���m��V�K�HH�6pފ�N7e�Dt���pWK|�Wg�9Lx�XxXi��Q�5���)�U����Y�.�s[�(lE\̎��cm�Ε�0-|���=}�6;5	1]X�zGK��S�̑E���JX�eu�뻡�9�b�Y�Ď>���Y{٢���g'`R�a�"�d?66nrs:�Oe�Z����FRl/��n҄��Ev��0�8�plkYͮ�J�HL�Ԙ��Eʁ�������a7q'�]� ���w�M�*
���s#�,}���3vL���m�85���|����PCI��N;7�6;RQ&lh�Z
^n�����Q�4۳�� f�1h' H��z�MZ�nA���1��]l,�י}��f�V�P/����a�9 WJ�<p�G>�l`����66�
i�Yܓ<k0��KZ�uEcB6y�\m�;�@���ɝX Em+��teV��-y�h�jdM豢!���& ��2,y������g\�1�&6?���������|4[[KT��m���U�XC�;0μ��_X˸�zsh�&}� �{tx��v����˫
:m;�<C���zƟ��z��'��#�V�x$��5�(�*�H%�/�Q:����B�ޢ���j�iU�����oj�����"j �oZ�����9#̛W�jj�#��}���S.�
�0]^u[��nƬfH�P����"ŀ	��s�odz[�CjT��LB�JX�w� �	fv�U��=���;+�����2-�Q�32l��L�",g7-cOU�]���6�s؁��_+9��f��[y8re$��}���k�6�Y�=�4�ޞ.���_N��u`���V��R�����u��rڏ1�&�RvVv�L9��c>����7��Lj���ی�z��r�LR�Bm\6t���] ���z�k-�2Ve.�i��h������E�:�'0~��۵���=�!�ѢQ{[x�g*�?��^t�8�4�`��K�yZTN��h�b/n�s���U� ��[�r��}�UӋ�gL���4"bb���rm�)hЌv��V5�ʆsobؕ���yq��<,�C��ETc���q��G�1ץJP��{�t0�r����\�"M;�8�7��pO�Qy�bJwA�U(Cj�򭯚���I���1����0�f�g��9���8w�������ViǢ�I;�M���m7��C
8u&��t(���"(WSk-a��;��3N'���~n�.Ž��U����Z�Bޘ4�ë��}1l��c�E�tj*6�ɝ�~�*ξ���ޓ���'�u���d��.Y\�l�V���7��[z�˾
���Ȏ2;;�te���j���u��T+�SB�f�N�FpD*���+s;0ܠ�>�\���β�x�LG�X��/�t6!�/�-�1�y��� ��+2å�Y��Fu�\N3����rL�z���'�c�Bۻ���s�g�{z��ZX�ih�0�̐�С��F4�U�r�H����ݷ0�m-�:�X��w�3��G�A����fÅ�b����. *4�P0Ȓ�W!/$s����Il�3;&+�'�m�^z�\��vV�O�|�7D�*T����$c.��Y�H�j�s��gƢX8�;�ʸ���xѼ�Y7���<��÷N����n���m[���czr�s�YK�cq3����8凒�R=�	���(����`D.j�/N��MC>�:�q�5��6��c���w�fގb����*���:�7��a]���݄�d͓�Mz��Tɹ3��|�^#d�����.�	^��reg*7]�l�c[.��}������7Q2���BΙ��m��;��[��w5�C���Y�5b�ʮ�#O�eK�g���d돬�iW_v:+v8��MV:[ΐd5f���Ep�F��n��{�K�,��֜B����S,�@g-�Ӏ\��;� ���86à:���Q�:çzm�����*\�uwe�A�=C����P�CHΣw�MjȲ\%�n6Ȃ��M�qh�A��E��x1��R����H+���@����y#]Q=W�VB�.�m���^��D�2�k��&F�Ǭ1(�����w�OU&#b�ޗ*��ֵ870���]�ԙ�*� ҉�AafP�Q�����%t��K}ʱ�m�L��Y�7�/��fw���}VcQ�|_Q��2W^�n�t�+�H{�ǂ�H�h��WnHsڗ븉Xϫ�vI�$�@��1bid����L3�M���γՑ�6l�(��[a�{f}���0���/xL.\рհUa�98ib�Ly��+�vԻ�q5��q���\��H��-U�ʹA
��6�7�&v��nཨ�z��+�0�=欹��b�feø����UW^�@�s�^�c[��]�V�����5I� 9e�E�]L!�Be攂]���Xw�&9�pl_5�7���(;eK�J�\+{����W���b��̪̈́�2�g/v���|Kt%;ٮgjdQ����
7�̱|2��LJ���,�dy��&��SMI��y,�=G���NH\'�SFt�'��߹�[}�&)!�M�QMt��V˗���Fy�q�.�T���.����n�W�z~�u����P�b��er�u�F�=�f���,�*�}�R�
i�(W�x���gM{�y�콚��5ĺ�d���sF�{�<��c�p����}�n�q���y�o�η�3,q�@��[s^�0�٦)@��8�ɘ�Wf�������]z��"����S$[�^��P`3yRK�m�޿��U��h�H�ٔ3�By)�NLct>�ҍ=�)<��^���;D�Cr�V�oHȂ�yxZ��=�m[L�<p���޻�$�:��e� '#�X�'7�&�@� ���:�����q;{�.{��ۛ��iQ��Ks�F��0�q���L��&�&i��	��-��vm<���Fp�i�pl��Y����*i�]�G�I��:.�s�TO\�̀�$kJf�kp,W���"�[�5f��&�jQ�h6��6AO
j��|ƒY!���7P5N�F�g �
�d���>0��Çf�z�'���2+��A��B;��`��.f��1+;���]٦U��D&-p놹ˆ���K�����}�y�;��c6e��}*�l�dj����D�X\}},����r��ρ��*���w��������4�ﺥDGd7�������B�BS���q�j-IQ��6�vॉ'��M1lA+%d�v��ע������_��f&tƶG�j԰q9�C�t�6^��4n.�(f�5�mH[5�i�:�{���+�	�p̫Qu,�O����c��I(Ċݲܕѽ⎬v+b+�.�VsouA�ש��.��]t�ǸB)�d�9��Zb3�pн+y
�:�;����{|�v\Gba�$󙸐ܥ��HƬ����A�,����y�6�N�t |v���#��#rQ=�Wq�Όyb:��/|��}�>'�}�o[���KJ�g�]�U�5���<	>Cj��w��GD*��3/�Ho.���Y�
���;�d��gM��x�<�+�%cRܭ˾ˬ��Lmg!�c6Ib_ih	���t%�H^$�[p�2�%�K��)U��/j�.yp������X|m%����)ѻ�k���*��p5%�|��X��N��r�"�v�N��7F�y3y�1�{l���'�ݷ�\�5�wq�'�ym�P���>etF.\��������.�p�{��()�k��Z��I�Yd��A�J3)$�>��*Ҁ��auc���u���+$�%����s�̜R4o#�.�i�ݺ{W�n���9Waj[A�Z��.ˮ���-�X5,ق�G&;c7��F-�j��I��[�w���Tz�%7|�qp�ֽ)�ⱈq�̼���W�^��DOp1�}�7h}t���o#��d"��3�q�X*7V�&��C]�XPP��s1��h0�U̰҉�z�d��Vkr8=��Ī�A��I���}����<�*`��hO�"�wH��R9 gM*��_n;�h�\wO�� J�rL�j�"�j4W��$�!�V
f��-�	HS�b䜂'�a���
���o��2��?m�=z�wV���l����vW�8d��t�l%��"����Z�r�2�c|q
�m�M<��[�|n���	]1Ÿ�u�H0v���n���|%incEn��.� DV52�u1P�]����P:=���������=��pU���NR�T*�h��P��<@��{i�z�{u���D�m� �G�tiX��NL���)��&&�p��7��!�����Q��׃�����ו��\�֜��gJ����cB��D:n@,�ňpH�%XޡE_G�+�C8��Jz��ga��BW+:.4:�/v��	dn�L�$.�0K�C�-�L}�-���Gy_L���̷#u���U�i�w��h�ۈUӂ�1������gF^9�s_��9ڸ(N��3D�:vAQ�֚�8f�|�E<_�&@x��FR�ύ�ƾV�&���@`9�-3�M�ԟn=�^��������J��|Bhm��j�4[�G�.{��nߣ���L�'\���Ws�P:������Q-n�S����C�v�����
�z���2�F�؝�vi�Gr�/�_).b�e3�F�j���&\�d�	Ekj ���ŝ��7B����n�Utx��[k�0��zw�5��N�����=+r��ר�w.�|�`Rʦ6;�P�A�)�g/!��sGr��Ȩx(Z�EWm�v��1��	:��YyՔ�<�t3���x��;_a�����Z3�� eZ��A�8�ƈ}�լxpb�x�H��҃��ؗ	�F��.Sb����k���g���r��e�Ro:ߡ[z�.��W��e��2J�c���U�����u-:FZxu�&��e)����/�$T��oq��M>;ԝs�X�����0�IV:Kw�����eǊl�[�]�����nY�J��=2��^����}���>�����S�Ӑ99��85����w}��"?�X��vxX�������1���*ї^�Q��{x�+;:cgX���::;4G��x4��t�3w:�Α���%�Ĝ��9�p�J��̜��9�}c#7S��xT��h{�w^�f�¯�x���tDR�l��(�|��n�tb���f�.����x�;�9�T�Q*����,;t���rv�g�#[j����k�o��;��@�S��z�:��G�.�+N�mpQK��0���ld�o���/�<&/Z���W}��Xb�8��EEW5���	@n�C:�!�e�+S����z��8�ͼ�����^F츪<������@�r�yS��s�1r�.�n0+����%}K��vقgMݵbԃ˽�$�e\�[���ڷ0u:)})�ô^pJh�/-�@Ԯ�=݆����R�X�*XCB�h�XE�b�py�����:��X9a�齛���%��.d[�f�/�鹱%�*���gu��ʙ�l,}o���H�Z62�їt����B�3٣O�&���0-A�whr�0�tA�,��o�*K�oR�Є�[���_V��>9R�\��Wm�[�˨����z�����q�y���mf�]2{���E!����g.����9��]˰���4�+�ڧ�����붑��:�����Rی�2�J��imacj֧�bX��+*-Jj�E��k[([)XTjQF�*�ܴ��,�m�jT�֥����`�6�V%�T�Ҭ4Uj,1�
1`�(����-cV�,�-T�iVѫEZ���kiU+EW3t�p�jR�h֌�EUQUQD[F���e�Q�0�V�GR�6�-EkA�U1����c����m-(��F�[X���`�m�X���ְ�KX�Y��
�Db�Kh���Q��)�Z"�*�����al��LmZ+F�(�Dj+h�IYkJ%����TA�FjႋAV��������MG#mEX1Q�Tm�*5�*0A�[�+U-J0����ŊVQa�
&5AF�Q�j��f*&Z��Ti��IWV-��5�h1U�Q"[Qij����Z�E���Z����1T�UF(�eV��X���j�Q��Vb�U�r�cmUM��c��b�jV&��*�#Z�����ؑ���-l�(*�����<��cx�+�)q�k�:^�S�k��2����Ӯۡ��KOQ���k(�Ó�6����޴�ʰi�6�;W���qN��b���Pcw��s�CHGɇ\�V������3�*��ēҭy�h����-�e7��	��Rma淒wP�+�w҄���P�A��I
�Y�I�IƆms8M�Ħ�|����v˿Vjp{�vV{]ј�ό�h����b�$D+�p�[ή��t��a��"�����3p�U2=��ƽ����7�
V�$Vpi�~�]��u�����%�o�{5� F�iֿ�Z#�Y�i�I�~9��!�(j\�,Uv�*�7aG�9";�/�al��}�B0<�� ���C~�X::�L�_�E��U��:3���W5ӥ�u�+i��<�<�ýgnŴ�?^U&������ƒ�ʚh,����,���z�����]��fd�dn�C>\��Eܣ����U�&\/}�WK���%�re�P��mo�����H�n[3>w3�t��	���9�pU���F��P�1�;Ԫ^��kqJRе(rA�3�e�s��-`�����P�:�<pN���?gV.��zw\:�d,�{�f����~����~��'F|X������T[�Rҫ�v�%s�y��S'�޹<�Ѡ��A
*����{;8���gY��5Z�X�P[�˔�т�j�,C�6�{n=��ZX�z��;�Õ�fTv)��D�Ek�gb#bw`�K�e�P��a��f����S �C��b�X�f%oiE��mNP��Sk9g�>���]vf��ػ���d�UllRsc�3eq�`��3.����m��4=�u�UV';�x>��mG�6��)&�����,q���wk��H�ǋ�E̼we�0M?��W3�O�D���|�S�ր��oz�ݺ���kb$M�]�Q��cwQmec��N@��9�ðJ�����^S�Υ�sXx�$��~-�m۹vWECn�ZWY���<
�.E��PR�O
g�eD�����C>�,k�S3ǽ�u1i�^>~~�k����8�>s�<B� �q:�w�\n�K���=�0��oJ�rVD�]�P����������}�\�|<1�ѱ�:�"�V��j|�^Qզ�t��K�5�x5��{���g��z�����&�`���s.���^>�j�T8l7�����c��l_����w{.��XK�������q�%�
d���[^J4����/�7��j�kx/�|S��Ev�4�
�6���m�T
7��o��N{����]�qg1�������2˄P���u��t�b��˹d<�
#˷���Wm�r��/|`�ۊ�wT�r~���!��+��%�G��ｙ��1�jԻɽ����Y�o��k�z<�j�2?_yC����u2������$X�����$fW�SZ������.'�s}��.i�R�5�!��^�0{���u�9���v����\{rN�>މ¶�;���}�Qr��̩cU�Ev��@�ܶfw1i�P�B%��O2��h&��k7��~���2	��0�z���0&:U%��%ᄹ�T�`A�`gQj,�C��ޚ��WjBs'-v���Z��)�Lý�=��Vo�E����$�z?0l���7ޚJ�}k����[�l*F�W4yO��BN���
hĸ��mFఽk��d�*��Ԟ���
�Q���돃>9%ۉ�	��(�x�xV(w�b�,����Qi&���ߚ�.����`�i�J�w ����r�	[p�{�֌ɷ�Yy9����{=h�vg��
��?����G�"��^��P��+�3���^
mî*#������z\�̮��;{�Lm�zG����l�t,��h�f]���T^�� �@�im��jr�w2���~t���,�7�`Wg$�x��`��+H�٫�w��1g}�5F�LY�r�᫱2z����U���Zb�76r��v�S�]r�z�F�d����X�`�r�g9�����)���~5�6�\�|����6���l�w�\�},n����xw��U���pЎ�S��<9`�$F��]��V��_Ocm�c��0��g��$�^u�@:�g�R�ê����v�Y<�v��I���hs���S!��B�n�׵$#�z)m�,@���[�'սB����;﷢4�Hć��Ϩ;�j�ױ����?r�D��L�//��g�?�\��q��*ӌ��iz}O�w�'%A��6�.{c�g���l+tq����^z���[Y4t�t)�|*�qhG{K��N^Xc������^�_��yE��o�!{�q?z�x���� �+p��9_g��T�u��^�j���q���_��m�����r�\�dȟoC��O��gۖ�����d�v�����Nת>���G��꓂��WJnK�-�����Q��^l��|���֨mf`���:���u&�m�YN"�B֧L#M�ޢ{�{5B��ڏB�n�&O��4hXK���j7���Gn���\Ǹ�!�/�H�}4ap�y1�(��AczOs;�,�nƗ-�^�R�3[�3���zZ*�b:�������\ൻ9�vm�d/%��1�;6�=��Ksg�>��=�GFS[�<�b�z���6��!чd��;�]u6l�sv���+�s��m��닏��\�z���&��=n�]��}�B�el�ٞ�x.�BEז��iM�2
u�6���<�#ʧծ˧D-�|���ү��7ƶh��S=�7	��q�W]��w��_�Jڗ%�ï������u�V]C�v��VXʋ�5{�Nж|�oM�N�vl��eI�ħd��\��{gY�.��<g˛���~s>��֥�21�G�C���C��WS��ʯW��f�j=�_����ܟy������i�m�ݓ}G�`�|�<���4L.�:�̘��Q��8��S���fT��������Ğzs����<;;3��[��[�8�g���emy��O(�ǂ�4}��-&�:����N�S��V�����	!�i%�f�n��3.�<�37�����GhvB��1Ĩ&]��`��»��;Ӊ�-3���tU�;����݇\��iZ��!ٛ"D^�=[���ϯ�bv�O.��,�n�o��w:�<�7��v��v��z����]���R��[둕���\�?	��3ׯ��ɭ��c6'�����[��R���z�E�"?u-�$��i�~�4�{\>��Կgϣܛ#�s�Nѱ�+q�2�{dM�[k�,)��ͳ ��l���ΌǞ�Vħ�,{ۭޮ��L��G����;Ke�c�����Cy��^'�F�1.|�wtҵόm����1�Vz�Ӣ��ik���Wp�foWB��^���!��g��Rw>;U�{ٟy��ׇ���,裮Z��(nF����o�.��l�뒛��8N�����u�;�fDF��C�����mv|��{�̮�{�����$��K��s��v��s0k�h~�XJ�=8�$G5�������u}�g9����W�'��?ic��su��^.!�M�@�}˦�9���6N���s(������˸��z;�����y	��<�y�6۝֦��4.\c�j/�l�њ�����(|�H���ǒey
.w���2hy���v�C����L=bu�aqm�sV)�ݻ�43���2f_�`�d-��<��25	�`�G~��iJ��1��Ws�xX�m�.��%k=��IҺ~L�,��CZWIu�uOf��soRF}J�-��3����~�2�}��R,YKw_���������>�y�</>���1%���ԧY��3�J��~>.�9�;���I��{Y�x���c5��Oӌ��v=������*;�v�O7N�wK/^�2�fԞ�������׾��%��%\w�'��gv����zlZ�i�[.4�@vb��l�6ܷR�r�s!��m���q�>��}��3�{Ɲ�T��h[�c�8f����j�/n�;ns���x����	��h�iL�m-�)���uu\YM�V-u+}9�o�}4�o��tϚ��=zKl��:u�]NITY�{���z�y��β[�HWQe.�O�n.�P��uǗ
�p��mK��8vӥ���<��rP=��ǩ���\6ʡ��a���y�� �(V.��OQO�H�YEo�0k�5�<u+Vy��N�ی�z�t՚C��Þ�Q7͞�]�^��ש�6;�u�+jjl�zd�}�%sU��ك�M���=n�Q�:���wy���ꋏ��JK���3�d�`�szV\��Ϥv8竏�n�=��{�F��!4��B9֦����/����I�.����#�0ě�����ݮ���_��u�U[/��F��8���İz>�U�ݔy_i3y��S�;�}$����K��V����𧵐�]fٿ?@�u��S���S��V���+��𿤛(O|앬������]T�,�o�Y�=ǯ���G�LH{�}N�����wm�8�[��o57�~��{�f�G��}�1r�ʷo*���6lI2��>#� �p{('yKu���s�5�/`S���<��ƅ��W�'p��t��F���k�c����x'���t/=q�nu��~��س=�j�PxZۺ��ĉ�J����*��9O�8�^��=����8v��js�2c]\��x��k%�ަ����U6��ڔ��)�����U��rx��:�uf�H��y�px��R��=�o=�n��^*:o��Y��`���oi���1�y�S_��+o���ݐ����2������uJn5냧�J���.�~�e��39�was7�:���,����IE�w�։<z�p��-9s)�*�����z�A���s�n�`U���f�Nv�^�fa���l��庝�;�A��&86�}D��W0^����蛆��j{�]A���zd̂Anl����ݝG%
t2����{a��z{�ہ�:���E��\�u���{�{�s��;�׹�|��
�{)���*�����l������-u}N�����+��n{�m�m)�Eb^��o8p��q���]�eӢ����4�O&;��^�ufb�s�q�'=c�L����他;!k<qyJ��cȡ��%N�m�A]��3/����7�'q�U��%�^��=��Ǿ�QYm���`�gf
i�e���#����>��a��U�@>�,~Yr�[
z�v s�٦/���!�5��3�hզ��J���m����%��;'78�����b���"�]govrrR�qY�^>�t�AR����tW`�1uA�����<�:$τ��|�:S}���ǫ���ȁ>2��x$i����ܝY�޷pmԺ�w�*�X�h9��.p���Ǧ�u��.�8=��5b��gΓ��q��&P	�_�n�2c�ڛ�)܌b/��׾����0s��p�瞘Ϸ�_���':ڗ�G����
t�#؇���Z���vý��&z��{-�~q����v��ήYΆ[�1$�dK�JS�<u�{|Wl��nm���~�ܽ��3<���a���zz�i����!��Y;��v�u˼jܮ�L_{\;Ns�~���}6G��g+�},��m�j<k�XO�cl�<;ų~nZs��z��R��3;�\�	}"}���s*ݾ߂λ~R}��`���~�W�� ������m����{`�^�o�w폂Z�]>������:˧ꭼ��6{<5���w�
�-�ٹ�+�h���̀4�,�V�,�ʝ1:�]�7�:+�^�.��R�B��rg�0P[Q�pkG�1
�E5��<>Sl�t,�X��pS�y�u�]��\Q�{�ǐ�{؏m<\Eڄ�L�Oz�Y7�*]߱��j�Ot��H].�x���6�6�#�"ek[��A!a��"ު�g�B�d�8ރ[�d;�ij:j�W@V��ci�/5���'90y��,�q����7fgEqT�K�w�;�Y�{Z*��\��z�gm�;ePɳ�/ҳ|^,&R:�+�;C�^`��{�9 �]�J��"�D}�	1Kq���%�=����Si��C�|�oaO�Z����>ޮu%9�]b
���0�@�,?N�3@9�����(^�kTu{V�ɩ�J���8�����7)*�֐oyJ�'� �R�!n��vr�>��v�FJ���T��R�֪�P��К�H���v�8>)[)M�.}pZ����u�_
^��_K-K
�/R�Bf�@[��Ő1*���鲂����n�8ȋU���ӣ�3X�t����+�#:;v�.��2�,;�*�
�8���<a̬���D���.�V˽v�vpX�ڈf��.�CS��>��TYt��b��'u�k�N�Z��>f�	�. 5r�0w��3��W@�rZ�Tq�fɑ%�VZWepXLa�Z�.�9X���h�5�WQ�|i���M׻�x}¹�=��Ǳ����ܯ8�:e���8��rG�^��t���.ٛ����Ԩ��{3fI׵	T��Y�H��`n^�*(]JM�6_}�r�<�mI����Q˖]��Aƞ ǝ�Y�A�����M��{ѧ���:�ynəi޳�x3X2�՘C�yݹV �2r؄���П9�uҁK�֗��6閬^�����U�t>ܻ��öɹ��y����-eI�6ޕ�7N K2�e�����4z���7$��ܢ�^��$����)���:�tW����ܭ�d��W�ۂ��&���at5s�k����e[յ:�
L5�;�[��f�+Im��u�v>=/D��p*h^��r�s�:����I8��wc���3"a\gq{�0��=Y�����fS�t���0����9!��j�5.�hQ�U��}�˜�Z��K�d�W���:�l�w{��,:ۺK���u�Y���̶��7(�/3�r��Y�Z��䭊�a�ݶ�+2�Mp�,t:��e�������v�������"U�Wj}�Ci������fA�Qȋ�9����=���^y�f��+�&�\�
�3*��^� &*gѱ��H��0"�{[	}�#ǐl�� V��j]鸮v��ѐ���7nKיe@�pҙ�*��	���c;�gmR��띅�{5��rDA A��4�Z�ҩ��q�-K-d��eҖ�b�[5̢"�3��K��U"9F���*������h�̶��Q�[*�1DE�_SnDE��hT�j�b�J�ѭ*�Kj,TW��-�`�X(6��2�U����]�*KR�h�K+mEZ����X�e�7j*�EĨV�Ic�xTƨfa��jQ�Z$Q���mb� �-��Z�(**%�c�m�Q�˦�%eF���4!Vٙ)TRe��*
�aE1�l��idTQX�1Eb֙j��j�TAE�J�5��E1��T
�A-���m��Q������U�YmE4R.ڨ�CY

���e+A+(�b�h(�&2���*�b
�jV��DR*���V
�eQQE-գ�UAM%q���Z�Ub5�Ab��[e�L�&(�Dh�Z�1�m%DfS�",�h]f.1�SME�V1-���m��Z1���#7-`��h����
�����������]��k��^f{�ǘ�z{ZM�c��؟���:j�WcYFS�5*�n��X��{�K��u���yE���kp�߾�ok�8��q��'��|�ʹگ��g�c��ׇ������?Vm��=�����E?4�����ړ������q�t��fJ"�a���q�!�>�J��tZ{��	+����Λ��?sS�o^����������r�[������8x':�{_\.��-��9���._��6]\5yN.�����n�z�� �=a�u�v>}r�1g2�*f�����z���UcR�W�3�#����!�I���	�6:���y���Z׳8�u��R�yӏĭoQ�I%_�[���ӱ�q��2���T�����|^��0u��y�{o��}�ѯ8}bĘ��p�Vמ�9z�E�~�F쁯*%���9�O:��y���yL={/��*��q�<���wr���μn�8�*�͸;=v�yn��ۓ�s����z���*��*�������{��5l������n�,�n�8�lNl�Ec�9��o.��<��7���;Y��bo���=h�@�g?,��6��<��=SX.��E)�j��d}���>��}���g����+E��Eɭ;zw{��R[ޠ�F�far�|�쮅oﾪ������z0�?�{�Ld�a�o���eCyձ?z��τ�U��a�b���?w��7��['
�kW��w���ӳ`Or��uzgy�̮{ު^�Q�D-1��Is9N�}#�ޙ馍�i�az�����ߤGq_L��8���u����pؓ��5��A��1�Vz�ӯ�t�JJf9,K��F���)�'�8��y��:�7���{0�mG���ZV��B��wk2����ﻧ��c�����?c^s�b������SӦ�����R�8�2s�ˮ�u�:��9��;���/����m&���a��t��-N��wV[��r�[�����>!�_}��
�5�%zvwU�~��;.��r��I/k �.İ��:��t�{EDߵm�L��vx׳������w��3�.<2���D�nX���g�I`��l��+ܥ�z�%���B?T{Qgv!1?�"B��t�N�C��k��2�bu+<]6�t4	S��Ƕ��ق�wˌi��j�n,��=�2�ud#��;�-���B"ϯ�!j���{�{����%~^��P��%�3�  �Ec:�^}K��_�g��߶#\�b&6C����nD*��a^���N�.tI��˷=����[�۳0oDh=�s�l���rV\����7���y�{�ߡ�5��]yr�fzc�ʜ5�7���������+!Ӂ����R�����z�/��;=e��[���۝l;syI��2�Q(קKX�����#^�����E��^	���.���q�ގuZ���oC�4'���F�g9��I���wp��W��{\}��eK��"�d����^���Ō��ۖ����{$s��L�(�;�ae�r�Nhd��΢�y��~�m���l��jt����}�4m�/)Qg�U�����N��>Ve�]R�Ke���v6m���%see�.�E��g���5T��3߾ׇ�=vs'y��׫�:��A�尜͇֬��f���w\�\�S=�&�&w�dm�Y3p f�����w'[2�b��}���P5B��d9��
̗�Ye>���HDN��K�҆�s�*�u�ndV��ز=n0�6�i8�4�ūa��7î���t븯�����U�x_c]:f���z�o\���g`tB�tP:���1K$�@��'��cb��}���u{�Y���}o��v]D-�.|/�GV�v�N_w_YC ����f�4�n7�\�����I��K�*Pl;#�V$�M{BM꒰�wU�m�����sͩq��WzIZ�:�=}�6������El@{�xp�}���XN z�����'Y8���a
�ɴ7�8�bu���?$�I���d��%_��z���|�o�d��@���@'�ǽ��C�M�o2N��?d�+	�_YO�X�I�OY<t��	�!����M�|��}�=gY?!����$Ĭ3�����W���S�o�+�����G�?���~�l� �79܅C��%a��T�2h9�4�8�~�+��s�"���L��I��o��q��7��ԟ�q&���8����۪7���4�?}���|¡��a�I��y�Y>A`l�p<IĞ���R'����$�d�vJ�s��I�񓩳,:�~|e�n�������^>xw�߾��4��	�s�<f�:é<=��<M�u����:���������0�'�;�I�OP�l<d��y�I��~�x�'��L8��m��`m�U�_����������~�'L��	�|��i'P�n�3L�b��VO�'P^��$�������$������N%Bw���y�'7`x����1���>'��B���n2��^��-��yW�e��[K��{��F�۶������jUOrh�;O�~$�1���]�W�Y
9y�v�o��k�Npݗ����>�y�
b��G�EO�a��Gy�]}�o�yP�8�ц���fB�+�A�}M�ru&-�	�w����=��g9ϯ+�c	������'R�3�M'�gY'�Y���N!4}�*d�&��2OP�'R�����I�7�d�m�x�}N�q������������ٯ~����z|��'��;��'Y'��%d�R|ԚI�l2��4���Y��5�Ad���N��y��J��8ʛ��:��k��;�o��_w��s�8y�=�N0�s�:��~�|�Ğ�2w�N��?f�J��CAhz���!��&�8�+$��!���}���J��zk���v�;���y�~��%I�?2�g;�'Xj}�:��u��̝a��O�<=�O�7�jN0�Oټ��� ��+'�R~��u���HQ�︁��4�9iuvФ�~���=�v'��oC���'R�7�� u����d�d�M��XLI���=~I��������{��+$�=�J�䆒��� ��Vj��;��I��j������8��w$����&2O�>�8��~��񓌝�~�<I>7�����&�?��u�O�4��p���M�����}��:���.L{�:�^��~?���	�Y����z��l|������q���̝}d?�2q'��xsY:��	�ߞ2m��3�����?>��u8�~��쵟��޷��k����N���=CS��*
�䕓�Y?e�I�6aa8��h݇Z�q���!�}d��s�OX@_��~�����
=X�Y����7��Ld�M�w��u�d��3�'P���w��N!�o$�XL��aY>J�Rq��j�j�q�����ư�!������#�?�f�~���j�z���_6����c4ý��u�w�<�L�I���T4��6w�!�=d���Iԛ�쒥I2{x²|�@ٖN2z��Q���@���~ZM��}����UW��V�X��3�X,t���4��SKҚtށ�z���юKw��c��nA9�d<��� �2�=a��V�%3�z3��ц��{Ŏ��5ҌX �3&:W�x/���^6�볥���t� �K����:���ޞY��~�i�i����}���q����/�{��x�������{��M����I�X{>�a�I��&�q!���T8��;�B������i$�O�d��N>�,� {��ڞ����^ᱳ����G�Y��z��!�ٷ�M��OǟdY�N!�=�:�1+y�:��+�YԜAHzw�?$�'�X~�0�I�Mo&�N���,����O(m�^��R��F��?��,?=d�6e�'�����l�d5��'Y?$�d�N1�	=C�79�Ad�����|���{�����O�{�^!ÿ�����2w�W�? i��{�N2t��I_�'SXOω6��0�������q���=M2u'Ry�'�i��<��D�!�>�M�}�
�P\9^�K��Z����
?}�VC�;��Y=}I����>d���P�06yI�Y4�Ĭ'�Ri�e�d�%M��0�~rI���I�~�� �p��ep�Q'���_g��o]���O�i�Xxͤ�!���u���O���u��ԞN���z���d���Rx�M0��!�4���Y�I�Tы������kWM;�,~�ݩ��ټ�{P���
~�AI�'�s�`N$�3�u�a:��هY>|a?w�������w��������Y6���R��#�~G���!�]=���K��5p���~���iY�x��w��C�O��6}���'�s�0���4}ܝ��:Ö�d������6�I�o$������������F�$���R������&Oz��!�d�6LI=C��8��>|>�C��J��=�Vd���;�'P�,�=�w ����'�/�}��KG7�����k߽�����Sj���m;�d��Y=aRz����=C��M�1��'p�����k!�Nyd9h~d�'_�}�rAd���Y���﬏�bSg��ҩ=�Zm]h��Khm�:[>&�xI���tN���<5�tZ��'���}Lsqm�v��nϴ{%o���GY�~�����3�Y�U��}����	;�d��N�O��!����2aQ��4}��,V{u`�X*E���4��Z��Y��}_W�>~׼����<��8�ɶO��N�l��y
�>Ne���>��!Rz��d�':�Y'�8�7C�i��7��>d�t���?~���u���U>�8���Ϸ�y�=錚I9���M�i'{�$�u��M���!>f�6syI�9�%ABl�����Y4@��>J0�@�i���8�z��1�~�9����g�_߹�~ǡ�M?$;{��I����m��	��d��ý�:�d�&���p'P�'uAI8��7�T�&C�ĕ�䬚2���|�g���Ʈ���}���}{��^�m���퇶�|�~��H~�βN�C��6������O�x��w���x��ý��C�M�x	Ԛ9�%ea?�ǧ�~�]se�>��}y�%d�Vr��N2|�1�����2q��}��B�2m���$�ʇ�s'Xu�p�1��)N�!P�'�,��p�I�#���;�}�|ן�oZ����O'�:}�	YXO�;�,� k)8��ό�j�Y8�h��2m��~���Y?0�{�u$�T4�'X�L"Ô?��G×+�ׄ]�_�.�c�����T<d�T;��a�&�o0�@���IY'=�,�;@���&�ɾ��'ߩ�:ɶI��ɦN��J�~2 \���	+���fw���x�==�AI1;9�>d�*���N2x���y�+5���I�O�d���g�M��4��a�I��o���	���<M�u�\y������\���=�>�od���q�T������	�;�2u'Y��'�2{퓽�z��'��笓���~�x�'��O�P��6��g'��C��fX%\3�zn~>��;������}���'PY?My�z�u���'�:ÙN��'�x}̝I�VCg|ì�d��'����Xz�vJ���n���~���B��(~J�Q�xk.�K�in��mE�c�G���odT>�{��.��9Z�fh�
�#���.������ĴW=ȸJ����� �V^S��\��,�H6��oU�:xV7Ӷ½����v��^��ݨ��H5ٮH�c&��|��6���x}�c��y�8$*q���C(~I=eMM�|Œg�p8��M���=C��J��w��a��M��a����~���d�'ϩ<�쓬���>�y�/)���뷟r�%d���̬�a��!�i����	�4È)'��p8�ԩ�y��8�ĩ���:��k�2N���ì���w~y��Gn����7�������k�RO�S���:�8���*O���d��P��bN3̸�=C������?~��N2�=�
���������<ַ�����g�{s>��9_���=1��q�{�q'2|��{�I��&���B�O���d�����Y=Aa�-!�I�nq��'u1�|���I�V����v��45n������=��~O�Y���	���P�o�̝d�'����'䟎���&�����3�d�XO��q
����2u70�O�q��x�睳�p��˭���� �g���߿]|!����ف�'Y>|C�}�>a4M�_�~d�'�|�q�d��I��2��'5IXN!�5�T&��
�Ԭ�]~����5�~s�cswݺ���Ӡ~I�OS���~a�57C�d�O�X|��,���u�~~a�9��?0�}N�I�� }7ܓ��O�i?M�$:�i7��,��|y����wY�����;��<���;�ԕ'RjeĞ�}�c	�OY���Z�8���!�L}d���d�I����m�Y'?�4��?w�'Sl� ��|���U��>�����p���y@���X��J�$���J��VJ����u��'=M~�o��d�ǟa
�ɴ7�8�bu�;M��I�������緙w�=����=1�lR9܅C�OY��uY6wxi�u��?d�+	�A��d������'��:vj�������&�>a����'�7�<?~�֍�9|.���t�	�q�똅<]d�t�.��`��%�7�סX���G�^����t'��<�c�C���q�^�7�D����j:+k��C�Ŏ2��}�&�-��)�w�2ҝ�\}�p��1�N�_7�X4�U�5��n����������~y�q�_�~��!���Pd}��>��{��8�����*d�+���<d����$�Ͽd���9�rE���C��o����8�y���s�~sy�z�<����;��c�OR~I�X��>C��gXO�T7ϰ�$���u����q'��w��I�'���RN�o��%2Nnd�Oό�L��}�~w����u����}߯a��O���6Ì&�߰�d��y���m��/�y����7ϰ�	�<�d�T&��O�>I�*�܁�'�����u5�������n���{���}�����{q��M�r�~xɴ�>a<O���I�'ߩ�4��(�7�z�Y:���I���Y��$��u��P�;�q���I���돺����οu�_Kn�|?}g�����?��O�L�M�d<gY6��:�<J͡ԜBx}�*d�&ϼ�=C��J���q'P��u6�<c�r����_k�����w�|�9��2m��w���N2s�O��:�<vf�Jɶ����4������'SfY��4n�Y&���'PY7��J��8ʗ�w�ٿu��u�{w�����k�~��O�i�L��d�a�s0�'O�w�8���O��ԝI=L�IX|�j�����Cyd<M2q7��I�M�XO�Y�s���os-���b�վm��?}�#��u�N$�*o�2Ad�s�$�a��'X|��OzY'��O�{�Rq��~3y%I�AC�VOX�X��N%�}����;�w̻�n瞿{�ӌ�Hx�5a�i�u�(q��X��:��hw�!Y:�]���&$����䟙?p�O��&�y�P����5�T�$5�x=ֻ��W���5��߳���������=M�Y'Ru5��L����N?��?2q���s�ē__Y6ɦN��׉?$���N&�;���s�/�o�}�Ӕ}#�w�.�xھ�҅u'��z[�9��
;Jw8v����]l/e��P,S~�ĺo#�4�y�a�<��"�,��Ĝ{2�P��=]5�b�h-i��MI��U9q��*�;p!��nqZ΃F�)���p�J�c\3Gx�d�ұ>��_�}��UU�{��s�<�/aXOG��T&��+'�,4ZRu'�م$�'S[���'����:��~���<~C�gY<a;���&�z��>������5߾�u��~���9�/I��2m����q6ɰ��I�4sxJ���oVN�d�P>Iğ2�'=O&�:ԓ���0��N����u�z��>����������y��vc&�Nv=Ì�I���u�d��?��2l��I�4�IR��=�VO��h�N u��SH~�����ҏ��@��W��]{<S��c폛��߾7�Ğ�����	����~a�I��p�'x���T1��=��HuY6wxi�u&�?d�*I����h���OY;�w|??k�\u��=s�[��}���!;9f�6����HW�6�~{�d�����a�I��&�q!���8��;�B����o&�N$�����N:��7����w�+�{�u��O�@�Y8�ğ�Sq�������&�q'�>��l�C߯Y&%a���$�N�'Rq!��'�d�+Ӽ�'�?w>{���.s���ޱ�ks��{=a6����I_�'�|d�{2ì���o���8�~�O��I���3l�b����OP�����LNyN�|����h�7y���2���}��s�/C�2~Jç{�z��&�wdߟ�J�a:�>���m����u7?Xm�M~���'Ru'��|��:����I�aw��y�kc������zi4�=C�S�O���|��=}I���2|ɿ��<`o�OɦN&��z�&ٹ�q�x�5���	���q�|sϻ����/}�s�|k�q2|����	ԜCa�a�m$��s�s�	�;�d�'ϩ<;� z��O^��Y? y�'�d�!Y��O_C��i�����L��Iz�_��(Ungc�t*����b�W׵w�"��W�̌ײ���C߱\���*�?0��hV�е�ǏB��li��7$��.�N�N��6��g������j���\Ř����C�L�𡕳��*J�Pv�
5��vжi�Xse�j]�����g;~c�����x������.�C�TɈV�G�䣕�Z��Ft���#�}|�Ly]H{��n�}sGX�;�߮q���3G�l�`����6��E֪V�΢�{lx{� c{՞ۣ9�9�5ݶ� �|&�pm�M�[�9�RA(��j=��5���	.eJ�_v��[�@U�����`����<���F1�$��Nsv�V����q�`�l��pj��r�÷Q�>���pB�C:��yM�/�,��|��������Q4:�Oeq��[Ư�ݝY��&M����/��ď_��B���{
�l5������"L�W�(h�̢7Z͚<��E�b��!%1�W>��Jp]��z�R��^+Q�}MU�mm�0'��9��r�W�ƃ&�;��$�uh�,=�����y��|g.|l��N�T/fr2��hT�ReFg-�4��d����t6�9��N��fOy(8\#>����FTE���/�c8m۳K�v��y'u�9+B�؍>)N뼳��J]�.��G��J\"ą˫o,��6�ѐK07g?r���R��T��uۏ����U���>D��[�q���� �_��D'(d�W��mn�.i����Iu:���;֎�_e�	z���9���2�M^�E�Z���\�ˇq��/
����(��;���fx�^�e�3;��ޅgC�i���>�23�D�T�;\�VX׊�oed�"�Z����tL��wq&�-��{:�����ٽ4���M7�`Gq�,ĉJ�ղ��6��v��e.��~ҧ6����29{W}C�B��3� &�ɍ���r�fIo��J��u���h�v�:f`�5����R�ck���UK�/�6��n�@�f�J��>��S^�V�7�\�<<��ýZ�ډaphE�tN��iK��<�3��ܽ�{imypD�Oj��v����,�� <n�RV�;�}E�{5���(�%I@x��X��
�<=-���o��f�H�Y��t�w�Ѭ�{I�r�(��D�eJ%��E\]��ݛY������m�����83-<F[��
ȷ&���[��]��n%�*���ށ�-�P��>�p�Ӌ��#c�=ӕ��GGh��|g.m�s�v�߹�ޢXj��dB�[��N�%�aˣ�x#�L���Q"�z��D���L�f��F�˺�CZrN'=�t+�w���s�\v\��3�#��4����-�<�f�7Up͕�^~W�`*[��5�Y���\~�z�O¦��@��҆h���2� ��y�ޱ�w+��j��]L�m��d�$�����D"�m��f #*��mCm�PX"#!mQ�cP*e�b�&!���@�am���r��Rz�qT�d(�b8�d-�5�QTUF �����J��b�ڌ���֤weH�b(�QED�*������R��l��b��XQq���Ej�mV"�J�UMR�S31k�KJZ����Sm`�-c�"(��i*��QY�֨����1�1�[J��
E+V"�l�k
�A���ӊ�TDb!TDGvb�1c"�B���Ɩ��R��`��b,f%AET�و�+Ո�����
��*�Ȩ¥DB��E`�U�IYQC0�cFfY�*.8�1��J�Z�ʂ��]5�fdZ��-(*��������kVK����%�UmD�2��*UT��ƣm��jEP,_��,��-�pd�=-Ps�d|<����KqMDB���;�g+
��1}L�����<��Z�Ӄ�ŕ�Jq�7��!	�~q�u�3����!�
I���*$�
�l�d�V~�	�N�ٜì�	����|��~;��Xz�����5'Y'���+'����VM$��ڗ�����ȻƹR����?C��N��I�=f!����ʇY8����0��8���������;��u���ì�|a?y�$��nw��'N?yM�V��l�~�w}�������a��H4��䟙ܤ8��:��LI=C�����'��a�N%`zs�%a�N�!�l���>7̝��c&��{����ڽװ�w�}�}�oy_����x3��,%��uu����3�@�k�~~b���Q��t���ʂ�vV�����������t�3{��D_�=G���������V	�e��tvB�x�K�Z.�e���:�YS3�#��7�睉�n��$���.İ��+Y�ugu+`w{A���U��{�j9�Fy�`{[���]�!�M�,K�yR���ٌ��fȝgӌ�O�]N����k���#�e1r�}�Ye���F��D�f�:��ͼX#۶���̣�{��V�j_�����^~��5��oo�F�
�k:�aAV���l�h�®���Dz}�#�'(W`7�wa�
��N;G��z��w�P��:L�HF|��nw�JyY�)����u���j�����=~o�x?uz�<G,ݥ�PҼу�,���\����tw5"W��"��  ��|���<j��|lF|�CP��t�	�}���T��/sN�W-��s���ӟ�s��q�'�����~��q����s�m�R��ӭ}+�a���:�ͿK��~q��۾w_�{5����E��8A��N��|�i��`��Ԭ��7������k��f�C���M�Dc��l'�k,�,�p��n_�˜ggH�n�}��8I{�,�u������_cl�|;ų��	Δ�Ǉ�{��^�K(ՙ�2O=���/'�c���t�<��Ke�Pu���������|F�}o��UK-�c��בN}�����<���N�a.w�J�0�iR���@�7Yf	<��k���Ys{0H��=n�\����3Վ<�kA��5��'Vޛy!\E���ٴ��~��@�]77:��Bw����㕤j���3�� ��Eh�Lb���8Պ���7���
�"H�(J�C�e��5Q�
���z�C�ꖓ˅�꾼�ޔz�o�r��x�乮��/����f����Q7s9��=4.�"�v������{S��O����lg�Bl���,��|]}��p����X�6���%�櫵��g�V7w:�ב���2Ța��U�Or�/yl��O�[��w��3���w��n�Gr��T�сQ���]�;��������]�u���ӽ��c�W����Ҕ�&z�kb=���b�D�{2�f }w˻�E�F�	�Ӕ��_��}A�;���+��.����ą��+�w5�������i��T�8_�y������_݇��+�3r�4�u��}Ϣy�2�}��o)�ײ�Ϡ��3s��rMѐ�z�f�����DUA�c[1g��S���u���^�Wo���y��8�����ZB��6�͈��x���kR�����Z�}�P�uD���{��Y�r��gsN]�K��\��@�=�6G��=j����P�>�[fO��Ә�'�{ue����{�$s4��	�6Ol��줖/a��P�R,���3K*[��gu�)�&�G�Oim���eXJ��:h��s2������Ջl�̢{�w��ZW�Ʈ�vgGȬ�|�Z]k��Ў�x�,�܅��?:3����C�}���v��r��"��GaI�>NF��8�W���V�����Bm�zVUx?C�of�������c ��tsװ{�f7�Y�N������ꝛv��*�&�O�~�)�ꌽ�=�$��j�{ـy��ׇ�n����$�ux�.��â�a�}]c�?g�y��۩�lK��6����;{�/|��\釯����ψ��|]}��C�2Wg�>յ�����Y�7�z��`%�S�t��Y���փڸ]}�`�]m��mS۷/�����x\�I+þ�=bXu�V�Ƃs��=�����D����)����8�����O�!�	'�]K	Z�d�n���Yb������1ƽ�R��W�������%ILo���g��y�{+��_vtW^�E%�('������[��ۙ���*��<��B[��d��j��lڡ�(�ݫ�w��(�Kvu�xd�P59.Jk��qqz��h�p�8n���VL��kvy��dy�Gl}�_f\���*������y-q�X��6ߜ'�̚�L�P��Z6�"�=}��z ��Kս��K�G�}�}_}�w��������3]�V�����ɕ�f�����m"8IX���>�+1�n�z�1���v����*ُ�ǫ��+�F�a:=���{1��|�����>{��\ڞ�~��%c���o���r�}�p�{��ܫ��v�:o�}&���r�u-��g�?z5^-�^6�+��<8�Ex�.�+�z_E�`�z�c�g	��a9s9N�	ޗ���W���8�W����ӯ��'b��\;�����C��5�z�o7��o���ܥW��,��Ի"�+�a�.�a-w�J�M�zd�|=�nj��!	G}�o�_,�d���pv޼=:=C����y.v+V�^���_��?�$��K�r�9÷m�XRI�X.oed��l��>tG3��-t/��.V��2
��x�lV_C=<ڞ�畂d�u:�ݐ��4>���c���]j[�ʍ��l�s������p4���ǘh�_A)��q���P�������{0=ۧ0e��ݞ(r{�m���vm�Ï�;������0�I�>v��H�V�X9:�+�5���G�i��A3����jo�q�9��k����>�����>~_�~B��	�j����v�7w��I{X.K�a�vL��z:��w`Kct�Ř�u.�fW�W}�n`R��+��C^Oz���u^���w|و��m��=��]��S�~�>����ѯ����b����U����9이n��}Ԟv�K���9��ռ~���s��ur\�4)�͛�f���� p��PwR�;=�^X��3�=�x%�<�З�i����q񿾝���Ğzr3��K�j�8��$����F����N}�o��s�o�����3s�۾w_�{,{<�X�/�[<���d�]l�r?A������;6�߫� ����K�8��zy�\[o��y��2��N�����������)�W�l�3���ۅʚ9N^Zm,��Q�w�s���H��x�W@�R�|h[e��[/�70���tٹk��9����#��̦�4y�?_����gd�8���=��S{A�#�։��G�Gz)rg�,Y�:���0�W���q�.2v	�Yسm>7�ζ�����^V��{ma���m��ݮK��[٥z1��=ʞu�Ԉ"��j�U�o��W����×	3��ƿ�t�A�����Y�:u�]N��`T]��j���o��W�����Wp8%�c3����{0����ӿl|�<��72]'۹��i��u�s�N����P��+.od����=a�Ί|�)�~���������:��5���u��yX-��vY����]^�M;�He'�Ǎ��t�/�vt���'y�%���}[}�jB����k��ck����>]:��{��^�ك��eGɺq���G��~�NL�4����`�=K�:��)�{Y~����漢�yE�^��o�v���~X��L�!�	'�K�`<&P��^���w�mb�*ݍ��uI��4��I�3z#Oc�[�c>�t�vw�`��PP��&�Y��+�k����Y��6i��*��ps�g����6�i���W{i�����2���J�C{�l��>G_Qf���V�i����p.��YH����∦�`�:�0,�`��O�5v��J���Qm�p%5����TN�o3��0G��[�f;����y;Y���^Y�����-M�5�/~ |>�}�0��{�J'��c'Zy�.Wٞ����c ײ�A�q����e۪�\z)��a7�23�:/v,�M��E�z�'�e���c={ �ɭ�סmy�n�&zϥ���Kq��{~w����Nץ����C�����kRjn�������ǪJ�����d{.g*7�� ��C��oR>.T�Ǎ�.�9c��x�g����:3w�=�	����W�N����sB�n���N܂t]^��V�e��s�09���e��Xآ4�$���������.LO�_�֚�M���I�\�V9�fy�ڛꞻ�۫�w��o)���FP:w�o�u�&�L�#��J��o8q����S��YTn�=oy�{u:K�fl�3�s�:u�u�gMu�u�c/1�)̙���T�3�J��.u۰��k0�\��{UOð��[�G�gd�.����]�f6y��w�A�}�<��tV��;YeC�)�=I�x�0:���em1�bm�<�nݮ�Va{�m����྄�O�j� n�Fκ���D�.Ւ�dTF���J��\|kޅ�z��|��� }�����Go���e_h._�I/B�%òV�ƾNuh����ʽ^�t|%�}�^Ϟ��������2<S�}!��m�%Կ����^uH}��A���sw+Q�ڟ
k묹�L�kGG9*Ja��͏�_Z�V�`����{G����5׫�O��*J���w�{b/�.����Д�p`��Oyg��ϽJg݇��=.������ʙ[�_?m�*5V�����Fd�ͅ�7�zr=ݭ��8��~ڣ�������Un�ެ�b�q&�LI~�%{^�lOy���u���4�l��?�>�˞=Y��'5�~)���Ӝ�_��{��v�L�ܘ}��j��ǈ��dzeѨ#��}>Y��f�lgy�\��n9���g��1s�]oqLVV[Q�(�=��az�:�)������ٱ�J���G���uvQ��YuP\�6��3啾P^��N���[�+/_�l�e��x2��óV���7J�6�&񐻪m�7��L�u3�lM��l�G��uG�tx�ذVY8)��I�lt�}��ŋ�Z�C/�Fo�>w�ԯCl)��V�1g�� }ۼV���/P������t쿗S��u:�6����p����cqK}s����]�J�}��{�a����x#��%�b�u���x��{+!�^�;����lb�^��oJ˛ٟH���=a���E�o:V*�yV �Ƿ1��鿳�?})�`=����畓$��s�÷A�xì�-&�^���ø��o`Cʙ�/vn���w��߳�%�T��^u�!Ao:���3�	����	'���6�+�%�[��+��J��~�{�O�u��|�۹�%K%o�fʺ{C/�������G2�U��Nb������V#�|,G��%��D�O}aGWyo7v`x�*my@N�^�{������$c|�7��;�|�l�xK�]y)��Βz�ǫ��wl;{�I�z��T�:ÞzpFv��Ӭ���>�=�����9ӎ�l�Q���h�����c��W
�3i�c�;5����.�]��տ����k����-�koaŊ�k�F]3�Ze���0��x(�׮�g1��"'rͮ ����r�X1���ӷ6���7f�Z�sh��q�l:�a7Q�Kks�T���b�J��˵��˫�vS�A�: oO]L���a���Z�fs��[�m���uu/BX��e�y��C|���X�u�q��T-rt�.Ae4�a�Z%Gi%Ц�����ƺ}�veǀ/D.�!IC��|���@�)c�;N���n\уk�RӼ���V���r�(ʊ�2��[�ȵ���_8ܥ]iΖD)��}�����M4�wʅ� U�s����[��8�n8��v�wUֺ��y��X�2��qU�ށU�����.�/Ue��յ��Y���u6:���lv`��g3�X��&mQ�����>a
'�n�٣7��K�0���P�K��a�7�^[��4��5M�3�BhAN�=Ӫ=;6�2R�of]�:��@hh�7����8p<Ug%8X�p]nfsku7Sɢ8״�7ͫ�j՜ܽ4DqӈQ0�8m��nΘ^�����x���N�w�%\-3Eݛ]yʠemX):`̡j��F���<�=�ԿS1����$���0��]�����&l��n��Ya�nqǩ�/U��Ʃ�@�X4�׭��T�w�:�i�H<:\6˺ �;k���#$������a�:���}�d����V1.&�l�=B^=.��9�%	ܞ���μ̩x-���L̆�8��j�$Zڨfin�!� d�g]�K�u�ޭv�Hmw��t�8:�˔��]��Y�5XA�9�+�����H�4>re����#���k�-�C���U�,�ܧ��0��(<�����@c#�Tӗ�R�7C�pp�Fp�:Ry�ᰫ����3[޼i�f�5�~�I�r��Af,Y��˥��5*7�q?��4���Dި�1F*]�3q�.�v�o�[��T���0*!� ���S7Oy����:XvGj�_�������S/y�l��Y'��*���WR��bX�n�7[�!������-�]$l�+������{�-Ҳ֙�^��F;jr'���ͧ6��f&Sk{��g2b�6���GA>1MpYe��<5��m��F>�G:��(j�KWo :j3�1"^K�s�{v��JybWZdͬ.-ч���9�3�㬞��;�˻�O�&�|��[���u�J�O����WR5�lB�7	�Wv��ms�$���iM���]R�����٪驡ق]���}*��*����F�
<�aI��F����
�t��\��&5N�N�E�:9�M�}��\��1���;��sV+�0ZK#rf��d��]��E<���x�]���N�=/��t�ǘ>
�����1
�*�T&!\aEb �h�R�E�"ʂ��0Z��W3&"�T�Ԕ�b8�F0X��[P��n�9J1�1���DQEW,Z��EE�`�1�i�
T��V",���V��Db��(R�UR��
ʊ���R�X�֮*Ȣ �,-�,Y�D���#�F8Յh��.!T�VE�

��3-b���fU&%�J��r�Wz��Z�KiDAelTDX�[DCVQdQ\l���V"���*�E�Ej�]4FR�[e�*1�1���q�P�*�1�֪1�(�X��Հ�b�"
�Y+r�\�UPF
�[L���D@UD\h��Delj]ڨ�����[�GT�"�����dU�Dk
���GhQ��U#wVPb��"
"c%��� ����҄m�3Gl{M��Q������4.����%O��/��lc4{�W`�024vMڍ^�yn'{��S����\F1j��]�J�ʙέ���S�Mw�瑏�I��{�D�����yS�E-�}Qfоuٶ�^��\��9�l	�7Sw����L�.����g(fgҽ�~5m�����p�\4��8��lc����W��}�'�5c�t����B�m�=�-���!��Z���o[���y�Q��z��1Y����i2}3�Lh��3�ɪ޹�ia�4}����0M-�������g��fu�=@��@��j�څ� ��N�#��5�4�%}s��7�$vY�tewfҕY��o+i]_wJ��=���}U��ك��{��\��پ�l�����&}�Lstհ�NA�B�W�δ:W���gM�]�}�f��/�˥Y����{�S��v��ON�{p��^�s���u�p�ޥ��ǧր1��R*m�ͻ�xd���B9�F��-k��v{�K��R/n�]�A��B�ڴ-lW�� b��f�G��/�V���Tpk��L�ﵮ
B�
\�h�׉��y�Z8o
/��#I%C�w_��|��-e��<�?�>�	%�Rf�a�}�N�U���Ft��P�r�j�٪8��t�#��bC��m�u/焠4m��Jv��:nGc��;Ϛp:����ｭ�)���X���wN��8�o���w��k�ts�:�����y���뙽�.����3�����=��50Oqv��h��������Xwx���筍~���(c�^zyx�o/8��\�*�{;y��2M�{/��;e`O�����sղߣ�~��-% i�������fzfl�{�֥y�=�C����6�qڌ�w���t�Q�n�K���/���&���3�'�3k��v�a�6/���Oj��@�z�ῼܴ�S����%�'Ń��ΥՌ?s�{��]l]�y��~�)��0�ی���ټbP�:�z�߽����+�xޘHԤ�*�B�ǉZU���A�ع��i����BR�1uݴ��[�2Y�0=��ҝd���r�nн���h��k�����fx�'��Du��yg��8��'�5��ɑ)Υ�䋐�����V�籋��qҜ�yo�諭����/]M��'?|l��il�R���/g��{ս�6�8QXx��p��K/	�y
�GÏ�;%�u}]}Q�>k�{�e��>�-�ԕ*:�|z����pن�Dozҹ����B���?=�^������8�����6���I:��]�a�"�B���t��[~�٦��2�\|���t��6���/�$��Rz�N�CY�e)V�^�4ܨ�'�}]�����=�.K�E٢C^$�*eE��Z=F�L޿E멝ǝ`�fXO]+�m��L��{Z5�KS�ov�t������q��5�;��Jϔ��
��Ճ7�g���%͑�Q�i�NB���׫���{�r�s���ʿRG���7^X��b���
1��^�-g��(r��^��gܳ�X�,��ݞ�	�OG�)zSY�=�����]%|A�V44-�v��1��p5�y[�]�z�;yŉ��F��"4�ݿZ3�A��7��p�̹�羖��}�gY]35�6��9�B���Z�{�SSt��ᡧr�p,�wZ�P���Us��k}��������> ��ty���I�p���oQz������y(߼��	�����E��Qk�FК"�X�t^fMu�Lw�@���Ԭ����4���q��޷n�X�j�=��vڞ4.�c3�7��������`�����������x�R���g�q���}�\-d��R%wP1-Ӊ��s���Z�,�?<�}=E{����j���Tqk'8�ogp���o���D�|.����Ou�I���1=�l����x#���Qt�0��`Ӟ�\'N	ܓ���k���U7����������\x��Zʮ��D��'���~^�i�a~}������2��]��Ӳ�	�����J�\kO���j���z7���w;���(��N6�O�y�/^�e˜Z"����� �꿅=��}^9/�kpʏ�U��t�����e���t�m���j�ם�%�':��h~���">�VA���[ǪR�޶[�F;fi�踕������I��Ρ��iA�^�\�-8�=y3���6�����R���\�����[+��C��KyM��*����?�����u:�sf���6O[�(;%����R{�G����2�g�nW��oB�����Ug@ep�x\�����D�O}`(��-��UY����Q�l��Sl{)�#F��C�b�������������וJi#4C��b�}9'[�w�f���O����:���7��#	+}�W�A};Ū޵NO1\[+�j�L�{s!��F�D౾r�Nmy�"yx�s�K��.�w/||A�z�r5�G�m:F:�|�_���׻�
��v��Q&Q�֢ჽ�׹�Hq��YG��P{�L�^��B���t5s����K�`���=�M�x���vf�l��Ү̒��$�;�b�ή��l*�#l�:��VЬc���w��bΒ�5־���$�"��X�_�.r�Υ�ҟ��I�z��d�\f�Q�J�����%��f߽g�G�Q��� �;�Y0�ST8�_4<6
��l��xi�������U)K�/�S�n �8ܕ���/9����^��3iz�x��qN�ϙ��{��ˊ�����x7�*���=u��»���^h��@G�Ǟ�᷁~�5�|ݗn�����h��띥�����|���$_um��5}��>�v��7}&��/��UQ{v��#�]��W�ܥ���̐Xd^�68�\[��;�4�1Ԩ����w:'��<�����$:�*��g�:�/>�p����p,+ղ'~����3{��j�C��5�%���x(S2�R߭����rr�g��jo�nVs��n��{�hw��f�4���B�Q$z.�T�b�C���!��C2[1M�J�e��o��Xy S00�kǀ2+�r�ù2�h�����w�{�p�u	�玷��볪�5I)E��`�nVD�L�W0캣��i�0k��5��c7��<�KOu��������f���IXr�`9���%&�>���.�Nʣ���j3�r�Oj��&�%0����f�ޙ����Q1�)��9y.C6��c��S�wv{�}�x:�/�9�hN�{ �"�*D�w��_ݾ�@
׽qkv�yb3�{�m�o5Uw<�=�uK"�#�x�;�=��W��4��_�>�R��2�.x�ME#��뻆HB��}u=�L��v!��R�D�oK>g�
Rh��n,ɺҺеNy=�3�D���d������t8e��6�r̵\hl�&$+�f���{8�ӣ��(#�ឺv��u���v5� �eskݹ�� )��[����q����A����g�) g��<a�x7MYx*��,yX�C��[��������3���}�`��n[3�ŧ����e�7�,{��^6;MYx*��ch���u��[嘮�>��+�&|�P�8�&��L�r���-�xEŌ�G^z�u��U�6n*�Y+_���4�lP�,�����C��&�z�l�4b�\�r���ǹ
;�^W����2o0�f
AF��p\y�:X�5ʢ�T��<S҉��9���~n�1n__K[y��y�/��:
�c^�Di��%���lS*��)�g�sW�m�=�n��>5jB�O����x*I1���oKχ2��[!�rF�/����s�A��ŔA������A\K�-��{��6�٢U�"���}r\j�S7ތ�
���7�����1�^��W��"�?=k��A�`�e^ ���IS��ç�PؘiⱧ��d��&M>�Qf��_rT��f����:�6�lI��c�$�k�>�Ǵ�f�Ϧ'A�]e�4
�Nh�����,���%ý�GZA�k� ��ye}1U�<�`tE���1(1�)F�dW��r�}�uö���[s�����,;�Qv�۳y�8�v��whF����c��F�;B�Vܓ���#��3��/x.Y������^��o��#|}�I*R/� �\E_�CiQȞ{mE�>�wIXjd�`�COKTun??�ӼH� �R�2�N�E���R�^]7\2�*�2ϼfo�Rz�{���;z����&��;�7��6#�#��ץV�6k����T��\�<j�_,���G��bf��XJy�q�ݴ�K���a�x�E��,����^�}�6�j�2%��ztz�N�6�������Iۘ�]j7,lX\Zo��Y��|7s�:ѡ֜��5g���}w�]KE�5��8*�u+�%Ca���=�"۱�`w3�'7=.ա���`����e���Z�"h�������YR��,��5"9�bly�3)��<Զ�W�����q��q~�^4�iE4��O}U�b`���E��ԉzWџg���ߚ�[�-�QI�J�E[���&��2!�J��=
ٞcW��p�4�]1w�2�o�^��b�Q̎a2�KE������V�Ξ�^K�Y eN
�D��1�RP�&�YS�٦���DS�/@�|�lٍ����!���f_��s�T`\�9�b��aS�Q��8+G�oRM�e�F�Bw;��ٜ���4���a�������9�4�"�
7�E�Ϛǲ���C�(� �V�n�q�; ��2o,�3��_}_|��n�\�ɲ��_�.c#qC3�a0��9�Qoet��gOb,�(�9K�y���8��5sYe^�Oح^��<�!g,'HKnc�i��BÜ�֦()�~����c�X9�0����o��- �I�c�<�
�+M��ӳk ]L������ܙ�,��!FwcQ�s�̹Ҷ�'9���@�P�yh�H��P�`]��=@��V��^<�ł�\-U�������W��NcSÓ�B���l�B[�Ieq�N���w_ެ�:�R�!�`M�ڿr)W�ɕ��s@�(f|][D䆞��Wޠ�f�a4�<���U"�c|�߻ymI�����.kH�7�
V�4o��`ؐ�ԣ�}�Y�+Q�:Ǩ�S���-����u�*�# �4k�}�Z}�V�k��3\��>��sٌ��x��x���sn���`̨v�{����|ѵ7>TϚ��o���f��ـ���/�7<�4�M�5Į�ji���]>��>�u�F��%VZ�k��i]#����L/��ޙ��,9vG�]$|����s٥�po��{q�ޛ�N^��ޭނ�Ƿy	p���p����^��f�t� �|���x[�-ͼy2?�t]��fi���(�k+�¨Ń��݅�-3%��}/���z�[��f��.������0s���ka�������{�ދ7�}&�?yd��K(��|_̸^��C}��>�Q*����ck�\�W67��z��u���C��uLP��*�6U���k�j��p"�W6�,�}���އM׌�q�-g�a��NP�Υ��ҟ��{�<6�FGGB��I!�5[�3[l�<��sL��\�5�lhZ�g\����f:��l=�6{Î ��=�p/��n�z��JI��]5z��+ǹ`����#on��ϹE5lF'�ܥ�D7�`�XdW�<ҟݝ���[pΤtd��!{QL�9͇�V�SU��ִ8ս��)}���س�0d���_�v?.�t����@ޮJ�up�p��Z�V0��wR�K-��:�&oOu�e�՟n�M۪0@�k�����gK�����[-��>��mZ���wcG'��"xD���d�`RF�Q�Z;��lp��c;d�W�/3Az�[ot��a7��G���? e�2χ(a�eه�UY�}A��N�z薵�IʈP�l=Ғ�6xǝ�Op�$�0쿍 � /�J�����K]$�@K���5G���p�%��T��r�ø��#>��x�:��*3,e��*֚�mj�|w9��d�0�d��<��}fe�ol�s���
�O+[l`���)
]..�6���hC��y�k.���_y����C��͓f��b�I���é�iF�5�gigдP�<��#n��m�wݝq��X��_RP��9�|��-09��S�*R�e�{��N|�wjcB
�V�E9�;�I����*,/��#F�Ƈ����j�d��Јv2��p�[��q܏K�.3��C�lr4~��]��J�G��j����Pt�o	w�Gq�:��1Z�=i���b�9S;`B���tι�WQl�M9H��83��&/��/c��sʽ�*���I�8�f�ݥyZ��'��X+Z�%ִ8��v��S�N�n�"����i��2,x��[��/�bU�|͆����%�C$�Q ����\�دr�T�]2f�����H�5��iY�Y��f�ӣ:�@`��X����]N�ș�Ji��C{�	Z��\�l���̽A`��RY�9Mo ��z���7����]խ��AvDʋ��ī�ð�yp���o!���i�x �`��%9�:�Wv��«S|.�'�Ԧ��̖�5r�'��u�M`�5�#Hnn���v��c�D\�/�JR�`Fd�®Vsp����42��[�M�������Wuj��/�۩^վA�d�E�Cw]T��E�b:��^P��BZ�4���*SU�s��jh��B2�T1�#8+���Lo�B�5��S��aWK��q3�� /�0V�n5��R��L�3�R�#U;�w���kR`�*�!����,:J���.5��X��p�%��N��ܴT�Z��1rX�kk��^՘�I��ԻΖɵz �坡��E�`�J�!��VPтn0��H�t5β��A
���x���ð��ll\�J����2k�1B������옸ک��Eoh>E�T_d���;���u��Ϸ��bi��6Sx^֤o]�Q/U�q��otT����wtH��N�����C�o�+�8#~>��vr5X�=�-py6Kuˎ�@b��j��fYc�H,l�yË���6�2�1�'��#��>s|B��\�I���v��e_&�f1��3F�9���A�/s J]7}H��c^�c��*d"F箖�2�m�l�j����u{���֩'��:���:���kk#� ���������&�񪒻_��<;\���]�[��������h�zY���F;�f���1ǉT���y��x��s͌��j�m�����)�h�[�\aN��T{�9ۯ!����'O��,�&�������t�?{��}肇�X�Y#<���"M����⑖�j**�r��B��F�U(�TX��Qb)t����(��*�H����A�L�1EAUA*(��N&5��Tը�.2����m�L�
����]�I����UF6cX�bȬTQ`�(* ��[UAH��(�,X* ���F0��"1b����l1Ĭ�kP*4�6�&DE@U�cPU��,V�]0�,DQE�TUb�Q"�W)1X*QQ�����b���2�DAUE�h��Ab�D"������
�FX,U�*)URDA`���L�k-� �Y��5h""����i��ŌV",AVe������"�DQAq(�QJ�`�*��v���|�>�Pl�]�ýoBNU��������~��mp�g�/����&�̮��j(yR%q؞�s7�� ���ר��.Wܗ��۬����ᓪ���S"���	)5�%��<qt�B�gh���������K˲Q#����g=���j�zY6�nX�f>#��ɢoY�>yӟ��<������/�tFJ��TyT�I�-�ș��[E�2M���ci���yq�7d�+�"�s/��	+�gݝbg�}h�YK<�Ko��m�V�O�;�T�c�뤳��ݗ�xO�^��)�/c�\��Ε�s睃Nn����n�X�Q���6��ob��׆&���kSn����-> ����.��b����+�c��sϚ�7�u~fQ����L���CI{SN��A���PS��o��Eŝ�O`�j������*�����J'D�QjZj$���d�ݕ	7�z�l�4b�\�r��S��myo�����|��E�HD�^:څ�\^\�/܉u	�҉�bM��W�����J�zV�P(_,8=i������rZ�����N�Y��o�>��ߪp�Z��د,�	��Y �>�[��š�b���.<흜/�M�ᇝ6����8�|0F��2컿��t=EÞU�@z�w��{��TF����NR�Qr��i��ڬ��Uv,�>���4*]��޴�t,�eL�l{��j�feV����F~X�6�+/'<��{=h��lP�d*P���i���U7��U�G�f-�5��f'[��ۇ^ʱ�X���=r\j�S7�L�a���D�"I�-$|7;�&�e�o��A̮:^s�5�)y��2��d�1o�ˇNL�{�z�b�WW��M"�.JU�J��Ր���W�8��>]�Qf�#��<E�b�B�����[������],���%��Oɵlq<l�[j,9����1�^8jDE�0c��c�Vh��`������>�E��'K�E�\2�/�x�;�����=�^[��U�Q��j��2&I�#��	��� �-3�X�g�"7�W�Kx,?_��M�ݰ�`�)�^����,��=�ȼ^��;���!�9A�W��C�Éf�{�}�uON���+�3��nWbcn��K�M.v���c����pQ�*�����:�\֥�J�E�qԷ�u�]�p=�"n�D�]�hN&o��p��M(��^w�xh��1��ƶg wL�IyWE۶�;<F�P��Zf<�Q�#T��~C��:Է�E�Zsw�J��M�ۺ����t�s��v�ޡ��|�+K&�աr|�e�h�!Lջ��y��0�w����vc]t�Zy��(���诤��}�}�"ٙ�;�=��l���y�Y�Ӣ`��`.�0l�"}|��4��N^	���zhy��;����y�V�w4r���#�=�G�'��+�O�Ze��aN$t=5"Ks׹��zϘ:�����z��	7pO�=��6
��-3��j�> ��ȡ���x�;fL��J�{��]�'e�ׄ��cH��N��~�+ygOZ/%�,�t	ik�
���+�/A[!�i��U�A϶�C�|���d��Nx(�[ޯ}%3���=��(�A�g�^-����Y���7WޝMv.F��X[Hu���Qk�2�M��;�]=P���:��y~��{��]�΅�x`�R��8<��i?4|��q}O1�V��Z�:�!9X�Fxf�n�\�l�0�.TŁ��<�y�ZI�]�wX��l�i\wle;��TR�����WIB��"�l�B;��φ�\m:�.����A��뼙���qv��7��m6�p)/%[D�S�:%}��pu�\��^���8�[Ѡ�}v�"�FU�u�!s.��/4!݆]h��-��S�6;�{��
�p�x��~Y2d!��x#�}#���ݵ�aB��}iv��/8�k��e_�߇L�!=eh�~n#���wA>��E���q\t�}��S���=�w>?���)�>��q�Y�^���ZE�o<�����=Kv��(��mZ.x����`PS���o�p���ǔ͏z^E�z��X���X��ه&#�t�[G�m��s|
^��=�2c�P��\C3��+��_]��0E�'8,o����r�Bds�[���ɷ�ta_���;�V��k
�i��sσ�L/����������^�xV̀��'=0�#�9m�2l�ܶz�L�Dl�6K�
o㢬�����	�������ԫ�ꗦ��f�)2�x%�ý(? �˝�1C�*�6٫�/��5�7"�k"mvߦi>��Y�+G������6�1:����X�����G�Ϯ�}n����
�OQSn�q�T��)5��E�PPv:��_�iE}��a��u/��L�<i��bz}�;�)u��exM��ϊ��eUq������Q�#떜5�e��
��k��&f�4ҭ��� ��ď���PL��c�-��k�[�Z>�q����7�fk+B�M��e,U�;u=�z��z�ͧJUGvb��>���0��xU�XgN�Tn����4���˖�g�{�;s`3_qf"�YW-Yd�����ɜP׻�F�����R�	�Kִ���ڴ0W�u �kl+���E�9u�5b�qM�|�6�����q�����^�胵b"D���O%�]L�3r�R���4�4f\�������=�����g�	�ޟd��o�%�X�C�!}��Ik��T�m�X�:I�<�kc��=���C>�,k��fx����O����p�L�Y�d��u+�oǂ�Ɂ�6�nr�i�b5�*5�Η,��`�+"�]�^����Taπ��>6����'h�@i���/I%7��e���k s��;e_p=�gIAnz����.��Ǥ1�.��ѳҵP!�����K���U��L�4K�\)�;�]�_�^�Fk�G�B��J������Ͻ�+i�t��"�^�֦������u��zx_����Y�W5ӡ5>��My�$��/�{�w,�vu��l��&|��/�Y�WL�}���ڬ����x����蛗.*>/Ӭ_y��©�C;4����'��|�T�L7:�OVJ���K��7l���38;��O���ɲ��2�����E֡ln�
~���*m����m�Y���˩���vn5�8�
�p�?J�]��7�8<U�(0u���-1���h��A��Xzu��|{2\�Е�����C'YgX�+�L��\�>��ݫ-1/���SSѼ��Ϣ{q�29�Jo���@���*�Ӣ����𪖻*�Ԭ���A��I���d8��̇�uKz�0�y�ɂ�����`Ǜ@���k?&�ȳ��^8�����V�� {h��yъ���EOLg32�aW��z�>���|��:=��Qg��,/�x�A��v^;�9��By����s"�_��6�δ��k�P�,8��˦��8���Iا}J��N�)��j��ܘ�2�����V�#��`d����xm���)uHő��\���l_���"j=hp�A/�q�<��6�עU�"���a�Is��2[9.��D�D�n�ŉ}�4��J���kD�F�!�xg�W�=�9�_�R��?|e�K^����|�槵b��Wճ/7�Dv�4�GJ%uP�����l;�:�>���TɁ�v<Dy��n_U=�pz�6>�JՉ�����yt�3�6JO�B~M�g�Eq�Y�	�J�|��;������:ٚ�o�������d�H�dK�˰�����������3>n�*e�\*���3�`w�1�cZ�x)�&<�Z�6��OI?�N���=�,p�-Z��u�`Ӽ��DktVi̮�M!̎~�KP���Z˸{��壔�FL]P_en=C9�W��TV�p4C|C�0s7C0��2��3j�t������� ���g���������S��5��tT�dևB4L�2N�#�j�쥈=أ,{hOy�T���X�f]��]�$�c�ܯb�	��X}p7������Y�+���x���0jit��Y�rʺ��?A|ӂ�vz�!c������L1�cb�\M����7m��X����#`礫�h+v{x����֟Z^՘*�Ԭd�_���^����I���Cd���>����c�sS͉�=U�6\@�+ϐCs�+��Y��_���5"8<�$�ۦc �/g�<K:�DIo|���cUhr.���j�������h���#l�|��z��	Ĉ�wm�_�]����˼��jP9p�u;�U���`�j�f&f|+-rJ��>�CgvU\�`����}Ƅ����^��#ܚS��P���&^Ka�S��ނ��t���]�ͅƸ�q���uO�y����dtH��n�vu�i`|���Ʌ���Q�.V���AL�t�"ɗ�¬$ޏU_�U���x��\���f�q�R��=^���{P�r�S��ٺ��
��H��5Ss���ȡc8J�g�d�>�}� �����|/4[�'zF@���"Դ��V.n��h�휀�����3w�y�Z�~���d]K�0��M���.;`.V�ۙ�.����ٗ}J�5�Z{�����3o�k��o+u��ޚ�J����������/3\����&�`u��Q/U3Ϩ&E_���НC�7���/\^�f�6�7�ܝ��Q��J��jZق���Z�:E�b�B�>o�_֨T��9�Z���}k���l���ѿ,Nӫ�\�5v�zP����B%'�yi!Z�rW�:�/.��^fW��/}�Vf�N��Z��RyX=���S/%[D�S�:%v$D.�Bp�[e˵�z�p�D<FX���u��B{6�uq�oL��H��2��z�}���E��kkj)��</�a���rn�hd��#�xvS>�KȻ�v!���%��)�E�Τٮ�u��B_k�y��4f�\8p�.��/B��Yi���2���P}Ҹ�}�3�w��wk�Z����A�=]�P@��{T��Y��x+�����_���]�����".}��}c����R~��9�ߍ����=��6L�Z'��K�-���K2�l*��qڭV��K�/�{"}�����"��-�fpw3����d�s��z��v��W}Km-��TJw|���N���D��U�G�)X���L�ualp��,B�����;C/xO7}x��v�]!W��4��p����O��7��iAIZ�e>��᲎�\v��o8�v��'��|�ͯ�=�=�nv����+֨�!|��dYO�|>_��S�>��-P�G��p>��k>�˧s�>u,x�[��=p����e��[I>��"UN�ԫ=Ǡ���}J��C�3=�^�L<S�8�_4=�P�����A���珱�}J��>GQ�WUW�TGuSe22)��Pd}�՞
/�n�7V�w�u�A�:�0��T����qq Y�1ݗ�݇��s�</�I���c2�1o=�d�����^��v�l�D�.�5�&��au2�P�f&��>d]�Q�����y��+#��O\��9�pE�a��fq���g��!ӠA�f�WK��,����7��+��hf�J��s��3�rƿ3<{�S��9r��tK:l�3==v���"������WH�I�)sN�]��~�N/4�_s��ȃ�2�����;~��s�'.w~pD^�`~4�C�b�;.��9^�-�(��,RQʄU�3;]��n8s�z��Ų�a2No `׫����x���,S�"�gmc�p���nx�C�A+7�V��IG@�X}�6En��-�n�J���0R �Y���;(g!����ɎX���X�z��T�cn���ß݁��'-6����o~ui�z�K�1�u'�P�`ͳ'�/e>�:��ua��z�T�Io���$))߼��ޛ��Zw�R��G)�  �e߶��z���E�y(�����L>�@^tyT��ष�<7w�Y>�o*�moim�޶��4��ɭw	"ęoJ����_P��X�'KڳK}^y�{ڡ����W?�����~Z�{}ׇ��ݗ�g��gK��7ln��ǳ��i�*�,N&�7)m�ݬg4רr�b]���Cb�7-�ꥯ��d�p���/N�/1mw��ȷ�+x� ج��3Cb���O&`��ME��q]9��T��ַ�-F�^@�^�7�kյ�k���oM�F�>�%��-^@^�� u���_+�z���N2Y@�	�����U��3/圼�IK��p(��0q��c��\�/܉������f�����魊(]��,��(ü���b�,��a�GZ^Rآ+��]���w���t��[�\�Λ\*{��9��Ü���{=h�v�Y�uk�
=�痧 u��7�6ƶ
=�2ݨq۹��mï~�i���>�.y]�<�O4������4�cY�b��T":�qr��Rٴ��9u�$s}��[;�%B��'���GA�Q)���y�W-���}�m��]�}�T7���{�^�u�(k{\�v8�[|7��J5ݣ]i	�޹ha���5�]Б�2�6q*\�V� тc�m������zg>���"�R��Osb��;�K!�-s��U�єT�#f\�^���D1���w1X��Wi���ӓ���SZ���^9�'�pFVG��]�*㺰���W��b��\
�7
9�
�¨��.6�=�;��ޤ��ֻ�+ԥ�v.yx�hhҼ��mֶDy���1�nr�n���ݍ����=y�h=Z�X���eC� ��t���t0ŋW�Z�{�
U�ϸ�h)��b�fM�UlQvn���z�}9��x,���?a�]0a+�-�Wj��;���N�i���O w��S�C���P;�����8qb|�rv� m*޺lw��,ù�5�wj�W���c5�`�7�z�D�3���N��+�fis�ta�e�z�7ӌz�C!#��!赝:�8r���_d��ts]�J�c�ݞ��ͯ_���_�:n=�����qjU�
*�i.�[;K�v��!d�E4UE+8�Z1nZ����R���=���~�5��<>P)�n��`^���`X;�OY%�/3�e���0^������Cݞ���<�ܕ���Y~i��%v��<;�αz�j\���� ���W��^�MN�ӓ+�� �I�EӘx=b�,g���`m<e�U˼ｦgIx�d�8t)�l=
��&�R�hou���7�p��2ճ;�ŏ2m&CJ�@t�g07�m���ѝb�����気x�k
Ɵ��e�.���Iv�2�%+4J��N� i��r��]��ilQ� 9�;���6x���˛�D*x������K�8�P���FX�9Ջ�2���e��c�)��0r��1K�o�y��0������{NZnc��>]d͵�Nh�-����tp�sk�8pڗE�N:,`�U}���%�
zL�[���2����c��ǈ��gR���N~������s���<�= ��ϖ�]JKp�Uw��8U*Vb�ԙ{e���/N��^p`���vn��fU�9����݂B�wL�;���u����h��n(��6���i�g�U�1��G�7/&�Oz-3�
\�<�$��[����i�«�ɱLw𧳙�i��|nP��P���)yo�\�V4�ٻ�<�@�JN����"������u��#O1������[5N����p���������R��H:4��+�ˡ�>u0�+80�}��nin�{���ݎ�{n��ۂvMZ��m�ǵ��:�9b���"#x�=�j�P����]r��B�"X��N�{$d=�(X�"� K]�M��&�iA��¶���3&`�9n�~~㎎��iݬ~�n�@�A$�RE"��m�E"+��j���"#
��֮[+UEMZ��.	�E��A\d����[lQƺ�0U*ł1�R6�Օ���+-��V��U-h�XԬ#$�I��Tm�X�eV�
,b��4b�.
�UF*(�QV�X*�k�*�,X��2"���U�ܴTbc(�X�-��"����i�EDWLuf
.Z��Qed�J+V(,U�����X+KAc�*��Tb ��r��)�b�*(����b�T���Z!Y�nZ��
�a��YP+5h"G(\�ڪA���r�-ueAUq���ł�Vд���b����Pƣ2�)dL���5TU̱A�1e��(�+T�T
ȥ�e������5��R��I���5l���H���<���́t� �G�ߗ*?xS�:�բ���=��Vn�P���_bU��,�X��9�3���?��;�^��D���R$��x�XB������N�0k��^y~X�1c�3n-�e.�|̿w������KC��D/���Z\+Qu����yla�k�x�/OJ���X���jS�<���U�1�V�0Gbr�&
���IW�)�T�"�g���)��\��vĮ�"�8{1�ʅ���=���_�ޫ��4������<��i&x��+��n�^�v�]�<�폟	1�w�Z����ϦV�6��&�t���X����{~��u�u��1j�^��9��Ƽ7+؟����\���ȼ^�"7����z��*�#]I�N��r�?W+��_J�<j^;�ەؘ�卋�-7��m,���u�X��:�W�)�#ݾ�X�i���[X}i^>K�	O/�o�5��^��e��;��}v��������K�v�X��{�\�ה�qt�Z��hu��Ɨd��5"9�|a&�筗Ӫ͏��:l�|o�ʛx�j[����xOl�ި͗���F��^z�����g)e���ɛ���jma5襾���&�/)ʱ��K{�����v��j����sC�W33��v��Xg���/Ԙr�~��b�.\�lwp+LGz�7Z��bj>n]�ȱh�\�v�Z�u���W^}&r�Q�>�L?���N\�{�����ƜK��,|�v	��G�6�\���: �����^]Z�0S�;�	���M�hW�ރ�i�a�f�f/�4ß:���@������]��=vM�:3�Eu��QY��'�$>P\�����3}�	��s�G.V���
g�ӭ� �˘�}��az���j:E,�8��c�c���O��GB�N+G>^J��}fw��=i+��V��e�@�J$�3���ƃ���<?�Z�����^W-
���oܦ��"�f��1
8.Tœ`<�s�ZI�]��=~�K�.ˬG3vP��'#��J�@c[K˅����J��\�E�,P�ZHP�k��u�\�K`��ɧʯWe���V��*[��Y�TYv��e[D����rP�nU�&��+o� �ޡ��4]8�P]JRmm�6��f�Eܴ������>2��4�,�;GZ��Ů��}�7}��y�Q���!�%꿩C�]i���3�h�]�f���c�,U����~�t6<�+m����ґ�)���Y{�wi3i/�B���qU4a�X:K��.��I�D�=j̛�E�2�i]�;܌�f���:�#(�/z�t��JD�TnW]�En�����\�m�׊=\�	��"vA��4�#r�g�k��o�U%�_��ѵd~�x�w�������C~�aϮ.�$���l��}��#N1��.@��;{�͊$xҚg'G��ǋ��k����t�X���j��ܤb�f��Os�6.��F	����dn=��6L�[=]�&u֬�'�)�|xU�u�`�[=�hb皧�#�Ri�0�K�`ܶc�v}�t��	���9�s�G�j�,�*\_Q6�7�z(�:ޱ�Ёz�W�[f[;M2�m�e�w9C�RǎN���OnC��h��S.�΅��8M���Um���q�1C������X=0�l59BԮhhOJ̠"�[~�2��ly�Xܟ9�Bυa�l.����q�eUq�uDu��ecC�M^�e�r%�[u��	��i��m��oz�� ���,26Y����"�<=�\\Hf�we���|z�nYy6ϳ�z�+a35�b�׾��_[���Q�����H�%��&��k���)�Ꞽ�zv=�^�[���rY>��qw�yrr��5�O��38߾�o|l������+�ӵ\��p��8��7�1��F��Nz�������O�H�t�pQz�v�vѦ�4�&�Kq��7�N��<4ib��qO{��i��Bړ�$��;G�3uu��bu��Я��ܣ�i�.-/�y�G�o�ۆ�Ek&q���Y����w=�2S�I���P�;���n���X������b��dW��p�L�Y���MsJ�r)D�$�L�fa�mv����k0�Y�)Ǿ�s��W��aW�y��]��	ڑu����yM�#c�W�"�[G�<Ԧx*���֢�z`���*Hң�t���4�vx@���`1�\�d����w�^S�"�g�g}r��f��u�ȁ�U��y�u裏>)�RN�%��δ����/��l���EX��jjS��k¯�=}��{Rt�݇z����x��P�,>�M_��H�����r��ֺU׊3�eY/$7E�ƭ�o#L�vdU��[V5�����0{���8�ݚ��"��oi����p�C;iU�����-��R9��W+�j���T���lPf�1��Z|\OV	�����n�EX���ƖzEy�� ~5��MYy�VڙU�c �]���Ԛ�2WNfB��^Q[��Rcx����1�6�r�+"a��g�X��������R-��Z�o�y�c\�(�BzU�4o �9[lݜyh�Gt���S��y�������]ڥ�r ���q�u�!�����C��ve�I��
�z�{�w��B^8��s$_�'-l�-�1��E���l��L������cZ6K�&����ԥ܏�8��A��Kz�z�7�TD�9��:R+GO��x/0(5ϵmB�j��� _K0]�����ϔ;�}�*r����(�>	4�v)�I9���u�$�j{��]u�s�sW�m�=�L���������v�}l��͚���^w�b��.�\���ϒƻ
X��L�u<��Ci$��a�<��3~Xuw,�:ʈs������4�
�����DPq_�ƃ��;�z�����/<��/�{pf��9��1A�ɹ�V�\�&C�XP�))4�U2:��C;��~�:�>����Z	~ْ��3���6��.�x���Y�)�{�����)>Z)4�k����'=�ы��]��'}jH�mR�$wI\P��+�9D�������a��ZI�৒��m;��;6{p���ɭ�3����wSş�tU��	��h���$؎����;ּ���p��F�;�fs�!O�Oom(ii�=�mv�{.-+�}p6ǈ�^-�kݢ�~�(r׽{Z߃�{�YT�"�U�|�^0ڌZ�]c��]�j��bͬ�i�]m	��j���P�9#�JƼ�]�B��ԛ\���|�P!�)|#飳���7(]�]�2��ڍ������Լ7;�������K�M�Jp`o�v?�T��=>�v��"��}��ȗ��[�4����L1�cb�r�T{ւg����}�׽q�^�mK����En1嘚����K"������ ϝ�������1 ��矊�4�\���r޽z6�a}f�\M�3�������E:�3_voI��B��r��9�%��j[��aqv�Ol�ެ����G)M�|U��*��u!>�V=�־�h3��N${Jq,�ȁ�����h{`�j�f&f�|����9��wog���xJ����NwȪ��P��N:K�p./�����a�����,��9�%�0bۮ��(�8M���I�˰���,��3}��&��+{�t�fz��OjL��i��gFFW0�T�.D0�8��u �u�z�^i�0��}pD� oFs���jq���7.`�Y��Lۺ@�:Q+�f4�d{���%�<��/7{�D����������ޗ� ���4��^*bp\��&
�Z��H���B���Ue,b�_J�&ޠ���6;k��dKgƏ���Ѽ�W�R��9n�;yCs���y�ճ�3ۍ�7�MՉ%6oݙ���tg��)wjw0�}BVk7;�m�>�faG��5�{�UUJ���V��{�h��Kb�nh=ss\���g�ɇ��}��vn;�=��s����\Zԫ�_}�=�	k�˕�b��>;�x v/U׃Zz��wn;p]���P�r����wFb��xe[D��z�BD��/}�����y�oVS�{�](��$<��O��]ȅ���ȼ;����x)_�rEg 2����ԩ�K��pJ�N���vC��i��)oZg3%�Ps��3zX��+�,�Y�9�Q ]Z;��%��/:g���c�)���ߊ�3닃��}~u�=V��כ�jg5��׹�^"}υ��9�,k�rByx�ۛp̵��C���.V=*��G_��h��Z�-ڦ�zJ��u��i׎�3����dn�C�3�o��ܰ	�u�N�Qu."���u"y�1l��Uu����E���W�5e��yi�,r٘�f�KPϦ˝ՠOT;�v�z���\�Y�{/��C�93�/$sXT)Wf\i�Z���jfRǎN�����X�����+9�����+-m3\^}U��
T8��S:���[�QE��	�ڜ�a;�H/B�z�]������m�����kSBg_Zq���ڞ����e�_�HY��L��At��/S�7�S!����=����(*�y�3��ֻ�w�[s;޻E�!Ov|f�9�t��h��a^wm.[]���]�,����ه�*��r�<���k�<��郞��yo��߃���ެ�'��|8_����t����1%��搩�w���K��v"�as�Yfj���Q�ߺ��k3��"�0��wk�h���Gx�TxzrC��۹S�3mJVOd���	��\{Zj��x߱�k֡��H�.�<ZZ�S/s_2�"."�S���p�6�0�޺vG-�.�s8��Y�.���%�X�C��WC\[�E��MP�v|�/��np��	�ѕ��7u�`�,k2�p�ŧ��8>�p��m����+m�Hb6M��HQ��}K��˰�_�{MH�}�K�g9���YbU?&�z�U+׼�ړݮv��C�yvaϟ� �
�H�k)�
��_k>2f�R'�'�)�޺+�V���

[���t؟Ih鿦]Á����H��Y�^�r��I2���@��Q�x�4{����`�8�AaXr��r�֥�.[ix_Z6}�	���b�*��'���Vi��>��0N���;��ȏ!�8>�My�$�e�+�:�XgX�7ּ�.��l�d������o{x��Φ��n�n;���g#�*��/|�Evs�U�q�wW�+�*X:�m�j�о��y�rn���1fa�t9ݞ;f/e�>���\���f�e���mu���{1�Ʃ��o��(�*��~�U~��ﵜ�}uq�@�����61\W�m��U�e阜Vt���v����\x�i�-+����?kMc�Ƭ̪�K��Ȯ�v��6(�T�㠸��u��њ�=��M;z������*���]�y^;�n�o�t�P�.
���}L��ȝu�	��\�y�U�ϥu�^3���+²&qz|��$�zS�V�P�����v���w��*F���Z�d�Rޮނ����P<��-�uYx)WwmA+��@��ԅ��2vŹ� �n$p>4'�J&_��xQ�yY��N]0�}�8��4�4����_v�V�;�U��5�xr�<�V�#ө�MΊ��w��P�V6z��{&�^�J�j���Q�����^��B�K��L�sW�Sn{*Ƒ{z�����U���!O�S�����>wD��(�ia_���ƃ�����=�W���д�Ч8��9�b�3i�ُ^�.�4�zﭛ2`�na�ht�Һ�GR�gk!�����Y��"��__�p@h�y!��]S� �;�Vv����C�]��<���dna���fͼj�\��Q��:�������֮�$�Ԃ��t���;��Q�v�s�����Jm��o�x��W�>��8����rV�x����*�(fO_��X|^��!:��o�ੳ�� k}��F��iu��.�x��R��X�%t����dm�琟�����)�m��ǐ{~�+�B��ߩ�n�_Ev��(����R�a��w�$͎
yf�D��ཥ,�����.��~��;����tS�d�Br%�!�I��D[�z��Z�fj�Y�>�xR�Vyk}����·�����G�����\����9�^/R��v*f�����W.a�:�"u��p��:��0U3鞼�^{s;k�0�ܱ�g�@����Uv��-�hK{����u�4h��Jω�^��	uS���ײz���]gE/�o���k�zpu�/s_��7���>Se�@�+V�g o�1r�]N`d�:g (��w��yg�a��y��d�ۦfS��x5-���^OƢ��6�]g��{sO"��W徃��;)��M�q���G:�գ�_'VJ��c�3k�?�; v��m���ɋ��U���%�4iƚOJ�{��&_�,i����1�V�?|:�u���e3�6s_��P����[������6��R̴檜�3[8:l�����=R���3Gv�9��\��Ѧ�
�@��}u��y��(�	�/J �������î���1~�"<���V���y�Wr�e��׺�7Ye���z��|�_:��sEb�}r$����+�&l�iOI�tM�'�RnH3�&Nd���/XA�5�	,b��6��rߑ�ɘ�e�lP*�ؑ���n�n�9��J�[/"��� s�*[r��K��G0�f.�O�x��}s�.�|��&E���n'gp\�Dn�؆��.�OG�Ձ| :Pϕ:�����	���ZF����n�Yx�+WKV�9lٵ�PvW0���aY��y���uQ��O��xv��/�?<�CM�Z��c��`[�XZHq1�Ovy�b�F���Й$����h\�(WHe��.[2�B�`�8��*Q���Wd�E*KǍw��_u�b���Ej[�[ȌXv��du�z��n�X�O0ڹ/��y	;m��Gq��z�W��w�,Wv�O�JH�;i��#���ՖJKn;C>�l��2�y��qTw]���形n1d�g��~��"�[��չ�>E��|;7(����zɱq��h,�8{r>�?7�7�:ێ�2�5�l+����;���ݭ#��fl�����w�T7�Tk�U!���@��2F0�ԫ3v�9@�59��sR�;q�qbr�Vߧ� �:�W)�}���7�]�b$�Z��sx)A^]��.�����6�}�9
��u��2f.�D�B]n�j,���.��sVu�u@k	Y��h�]�aYf즶v���O�c�¦9�]��V��7�:�J��	� �7ҝ_Y���%|�X�w��x ST⊭\��v�69u�5&�:����CԊ��Ͱ#� �lP=V�8Z�H�YԖ5y�!�-���>�L�FL�B�\ޮ�v\�+`l
�%,��n��D[�u�v�3�n����d��lJ�#RQ�/�]I���vN�i�Ɂ۠"vJ���j�T�m�Ŋ�p����/i�����#:�8A��f�m��+,d�x�Ɏ0�Ԧ6r]�Pq}mWn"\��s.'��Ǒ2���7�@���ۧi�xi
�;�]v�!}P0����J�6_�D�>�z�N��b�u���p�8lҭ�C�&�.
vw��ov
#1�1P�Z���JI,�J��F]V>k�-�Q
sYS����
��Y2���a���J��G�LT��.�i)g �>G�R���_�_[nY+�k^=�]��u���j��� ��C��8��˅?� W]Z�E)A��Bޡ�EܛS����+i��ΧD֙נ�]3���>�Ga߁z�ф7÷X) ����礏k;��C��xEޠ�֞��sy�xI 	Q�RB��,�%and�eKL,*.R�f2�
& e����In\�I+#h�fep�
���j�T�VQ�&���q�ՊŪʍ*�VH
�D�++�P�c�(�OYTa�Y���)RQQk1��Ă�kb ��H�TJ�
���*EEƪ�1��eJ�8�-f ��*���%(UH�*9m-DUJ�TdR�YF�I���*,Qb+�eEQ�E�DDB��%�m���j
��-�����E�TL�S,��!��e�J�eK"�
�*���e�(5#���2��[`��1���JʬPVڂ��V���(�HԵ�J��
�>"� ��7/^�XN��o]x��e	|��/Oo(��ؚ�7���s^�o��d'��2�=���g"��9�^���_�}�Β��p���9��0چ�	q�#���]��v���&f�l�a���
9]5�N�?d�����sU=ʃ`�{Ob,��h�r�"|C��ԃ���SK�?/N��[���M�Ü�����+B�,���W0v,xi���(����eȡ|j�C�F��u^�w��@5���E�����"�^�S��*bɂ�����Α��z�7ΐ�k2�Wޣ\�����J��t��|�Z�u�"�g�%	k�������A�/`�Lc�8	�ݼ��u���j딦p�wFb��x�m�COQ�B����O��^�.�0��g݄�낟�/���w"���@�#7��\��i�y<-�4�3[���%���*��Ev����~��P�:��/�����4綠h_>�'JzT��������Qǌ�/ug��:osn���^#=i��u�L�_������_�=O�aeziqὴ�洈'Acs�cJW�_&�{��C���H�����@�Yg^�]}��^u��]�(�Eo�IM��tN��;�ӫ���ۅlk��F^8_���R�s
{�.��]4_�/2]�[W���u�V��<����:��UP]���g3�1��u�h�q����ѕg]1�m<�{o�����+�}���QX�����[����+��^��e���˲7>n2�}6L�Z'��K�-�+�����LI[7Q��]���Dq�<��|���5e��Z\K>ܶfs0�J�9��uh����&��l=V�u��"�_,��1^ !m�p�4�X6�2��s�-JQ�\T��۱���?߿~�/S����ې��-O�h��S)P�w���[�QE��L5�oK�i��:��[���L������v��Yb��7��\��WK��uDu�:�uJ��<04��u�wR�FC�Gۍڂ!�f�A��0���;���t�+���8a�V,��{ ���yw�e���]��0.�ɵ��o{<o��5�^j�Q"\�@�&����b�ҫ�_#�%��o���*V1��O��Ӂ?[�����8"���I����Kx�S��=�T�ӌ�"8i�b��v}B��Q(lcw\��X���W+��+�~��-l���gyr-=�^�g<�=с���f�����iWi����K�s�(��VD�D��I�*_��S:��q�å�r�]����ce��z���Y��vU��*��l컅\M���[<���¹�����C������9dޗ`��f��s��Z�"�~כk^��S����_�Ù3g'su��Z�����7t1�9"��ז�Mc��d�M���3�Ω�zO����,��.�8�#@�;��<�/����]����#']�������=�7�`��n�%�d�։)�w �K�`�$a��=��r��G�e�����aIk�{)��4���
ܰ���5�{��r��.�x�)Ȝ�T��4׵���,M�U��Ԙ����Y�m�E֪��]��+��g��}�߹n�z��5OZ��]n«&z򧻪Q��y#�\�q�Q{��R/�^<e��G�^ǈ��y}�g���m�6�+���>�?l�X&`Lt�])CU�dw݆탃�ؠ��fc������6O�ɛ�ϖ�x���7�e��+�Ǖ�?F�����	�*Ɇ�D�E��t��(6��7q͹ωJ}Ss�u-��Lý�=��VojT��U��-^@a���6)�cI{o�b՞m�}���qPyшI�#2��u�����+ాm6Lz�b�%{R�]]]u�Ή���}}vf�r$s�Ƅ��D��xV(w��9g�<l<TF�c}ޤ�s������v���0;��p(-��8���L�ϲ�38�Rޙ+p<X�v�MV�8�-�yL����������cff��gQ=���R=��L����C�qv�|rc�w;y�� e��w�썏m�lůL�o{=�M��7��N�Kj܎�<���Ʒ>�P�N�:˚�%m�=�֌ɷ�Y���a�E���^��^&��j<NN�@� ��S>�C����˧S˾Sn{��E�'?{Þ�Y�O�>w��o����v�ɒ���e��4Ms�I�G��Y��\wT��n�'��h��^�Vyo�;�=������"��}�!Â`�o醑�K�U3S�u�������ۗ����}V���.��TɁ�˱�R��I��OJ}�`4��D�y	�ڛk�:$v|��O=ֹaϷ��V�S@r��K��]���i&y[@�t��}M����PS�}�A����*ڦ-�TW�	��Ѝrd��"-��b1Q�i�����ٲ6���=�=y��m�k�r������h����5����7��:����6����]e-[^�����k3�x���[�L��L�#�S;Oó��D�jc��`�O#��Y���#��ܦwzX�֜�,>�J�ȗ%�/ײz�C��9N�P�VO.і�{��rWV�j�j�ӷp�Wa�Јҝ6�9�=O.
�,��o�S�YjO�Hy�1���)��f�i%u��e�}���)�0��Rt%�Ol��˺��g$������n����t��wʼ�;O۟��{�K�:�b�#��.�k%����8�V'��ܴ?u��,#���.�Jǡ��`7[Lzܞ�e���G^j��I~+�3�u񄝤��N^	���\[������/|�)�qЮr�T���X;��ѝ�Ŧ�V�*�S��5"G�R%�z\"�N�<����
��-32A��.�Q�=-�w�����,4<l�K�Cf]�x�ƚOJ�{��&^Ka�S���E���zx̷���!������E��p6���Ջ�c�����fn�&{٤���Oz��(�L�9���F����
g�e��	f�q.D0�A.��A�K~X��������ݘ$�tc�����Nw��(E�;j<4͇t���:Q+�f4�dz�a�</��ޕ3�|�,�S�cج)'��ø�*y����I=)��1D��F�����m�DR̘�{����\�e�emu/4ˋZϥ���"�g�(K\E�%���ü�i�����r�3u�E$��j%5����~A���K���k�3��xe[D����]��)��fu��ô2wF������F�m1��g fjw3�Wӣ;ڝ�A �s="�ܤ�l��)�n��A���}hbO!�	T������KN��*lh*#E.���p:xQ׭�k��'���q�'�w7s�HY�wUzɞ`���'w�����ۥrv����D3>	��w��Jr۪��ٷ�xwW���.{�++P�{���5�8`�����Ұg��J:GƊ,�6��>�ԏ	fV���y��[l~E蝋������?>|UJs�b��`Ç���8Fx�)�c��B�+��ˋ���0����bT�HnE��[��~��G���K����ew� |�p�/��;�^��NضQ�לba�����"z4���ћ>�l�9��8/צD|;/�c�dn|���(���A�ט�U��qg�f;�0v�R��-D�>G:*����{a1�����[t��s0�Xz�	��utUu���u�ǭ7]� ��p�M[H�!��2�<i�Z���\�����g�YB�{U�a�sz���GoWh�܇��,�ˍq��Vژ)P�.�����J��QD�f��"n�&d���y�����yq�I|���C݃g��J���t�=㔒��������A�yg����aPD<�խ�v۵"�f�a������+N��`�������5̧�}��V(�C�ٸ�
�Y�}��;�z�qB�cޱo�k|��l���̣�n�h�>c	���u�B�ظ���D��f�|A�ÓGf^S��A��F|�07gB�ȱ�/m5�V˷ti�4�ˢ�C��f��Tv��K����A�8y�����٘:�O!�'�sk~�i��f�-���^	j��$KK�	��򡺯���̸�j\^�y�ҍ��p,�ž�!�"��.����#W�����T�6�T��n��# �4��..A3�*%7U�p�,k�,m�^��6���\W^�l�^���g�.���f��HC].)^���U��b�f?f����e��Tۚ����w����:wڼ$5gF|��o�C�l/�xg���Q�8�_GӋ�& ��X	��ܯ��k�%B*��`䔚џIh�2�~�����*8l7�}E�7�vx�%��B��n��/֦��Go�/��>��� ��[A��8M��Z\lDq�c�
�>Gst�,mS����_��<k3�<���[E�2�L&�y�$��L���$M;z�ޡė��5�KB�V�9�R���PS����~��:�Ɠ�Μc�a�o���b�y7}ϵo�bmi���4�۵f%�Z�5vXdWa�`�!�A�L�����r����r�4W�Z�|�N\�_1�Q�͡ދ7�\�C�2��*f�@,�q�o;"}x��j�ۛ���^"�����Eٖ��J�秶ѿz�K���-m��I�ʰ�����=�비rR�^�ױ��� ,uvGw-r�cs)��%m�}�W��nDξ�E@��#�n䨐|�Ǫ֘i�ɲ��^��0����~:S}�M<�kTns�j�o��r�6�\��X��̇�RިY��\�
�I��E��`|e$�z��&������z���g5�L�jlo�
�:1	:�楽]�����,�@Q�|��%�d��wGD+�m �r�I����T^�w"FqBb�J&X�"�?[�٥՞��<�k��xRv�|�K�����Q#���iw)�����3���^�����h̛}�2s�O��}�e���m��=j}�֎�wh�����e��p;w5{�6�עU� �5��ZW޳%�A�Y�2z[��d�s�&e�s�I��� ���h;\wT��z�H�=2�_7�W�~����W�8e��%L[~28�P�����%�µ+�Z��u51��G�٧�=s������8���LJ��D��xd�',Cbe$�$^+!T�6�����m{YS=+>k��k�ޗI[P��`蒑�)y[˰���0/z�-��vc ���:<���(Շ�[�nyOh��]�
_ w:�@0ؕ?a;�ιz_��m7�=@o>��9�x6̖�2�ߛ+5I��όjd$P�6�}�B�up9����w��A�h�����r�!�
��+x��m���y�]�;�Y&mYi�o��f�_���-v��)��kC�&Ć�'5���Ok�W}ר�ڪ�W-W��g��->�$���ꜜ\U����U��Z�G�r>�_��{�U� ���j�2%��V�
�)�]i��ueL�N����/&��Fڅ�Z|�4�o����7�嵇֕ᒩ.K�yx}����ă�pȧ�[�]^pwR��jx�WIƇ���tf����D¨QG���-X�b�䫾^�O��2�Q3p�h��I{t�NU��5-��0��W��`��&
�]n�y��x.xvR�lz�)k��*��8���ԉg��-�����h{`�j�kp��9��Yӓ�K���Q
����/�J�ʨ8�Jޚ�n�&1�Ƙ}w|'l���q�^V7�5S��Go,���]�����Iׅ˱�N�Cؙ�����S�O_H����3z�0	'`��\��W��S=�-xK4M|�.F�\a��]��^��#�e��9W�ґ������m,�A������������W�*	V�6�X�P��ʽ��ʽ�]+O��D4��3�f���v{6\ǎ��y*e�����Dh�eO��vL%>��Ѽ��f�)��@��^��Ky�~�|����q�nw�:��᭱YW�J���:���=k���Ϯ`�Xe�@��J%b����t=�w�g����c�7����{A�r�}�$�}Q?a�M������>�D�A��-5��gBK����7^�ZP
�2�.�� K����qkY/.g�%	k��r�Z����#:Ln-��l�G�A�i!R�3�f��z�Y�3�K����wFj�ʶ��5�[}v��=��dݏ���F:�!��D5،��7�}S����o�Ȟ�tvLO�n��LOG����t�ew��Gh�4Y���Q�^��ygò���zg�����+)<i����ק��{hO�v9)�P�{1�|��#��c�P���C~�x^+��$8�b���md誰��s!�;׸�>+����-����\�������9��V�2��:�߮]\}�7S�ǰ{.��#�^2#�^1��=�e	�^�c�$	�#=I�x�[�ߠ����Ŕ��0�/���Y`�Z\K7-���aޔ�߀��U`o��C:�H��%#-tF���v��7�pa��k�@P@����_a�u�+SO�b%ub�CB�Y� >�ưR��1cn�c�/x\z�|��mH,�q.j�SD�Va�MmC�L�E�p�u���KXv���وC��T�a�t�:��Q׻Bf�T!_�;گX<aʹ��O��=����ej[�;|D�i�c8����h�◊�:�U�;��{sޟa�*2{�I+��,Ně�T�w�iAWaS�WY�K�KXwP�!V����7�%��<۲�D�q��@���wsh͜��vU;�Z&5��Wϴ��];{mR��*VR	�#��w=O!�p&wL����a�g��[OA}�ʡ��U������oN@.#�ү5��"~l&���lN: ���_m�`��F��{w�<H�!��1�s�wat�˛�C}��iwj�<V��<%��k8{��vv�&<x5�Ǵ��^�߆*���\l���t�ÁL���,�ز���.͟��Ar,|Iz�^�7��ha����KAg^�]���V�Y���.��/��]-��ގ-��8-�󵩊�(X5�*�E8�}�,�����N���-3.��s�vܙ:��ƒ������t�UI��m ������F_Qﺜ$;�iNA@h&��;k�G���.51�<�V��=�t3�K�ܳ����rv#���B�0��B����J�z�.�F�!��zbk3�����#��WلQ�|��.:u�TY�s|����;Aʰ���\;m��T�ggH�z��:k�=�o\5�I�5o��Zy:{�|/��D�ˮ���s�/_P���g��/0�m[̄e�Ȅ=t͏���w4ݘ��n+w�M��t�c1���Bi����l�pIf%\'.)DbC9>=B���#]��i�8������P�x�ac��G:�*�{�ҕg͛�\��o���<�����`�G8��㨳޹�r����WB;��^o+����;��j�<ի<qb��ʬ�[o6��г� �����"�j��&,�s5?N�����3q&�Rsy��XT�,�F��@S����}�X�<��,p��	H�Nr�S�� i�(�=���S�`y �j�L}�vh"W+�R��*V�4�buwt8Q���H�u�U�cCh��ƺ�2�\B(hoL�b�m�NM��qI8`޻�]kvh��#;2�@{5ZcH\�jU�g1�@�ٖ�U�Pf�' Ų����s���ݛ�e�-tz�-����6�u�^�}Y�ޒ�əV�����z���!E+-���/����Z��4��Z�H4��٘]�g*|��J�z���H6�u�s��xidQ�J�K�Х��RB����>�
�I:�}×qyq�o;�]a2
�����%�X,�ޒ��}�)�����j����̽=�%.̭�����v޽�}u޽���oW}B�W[Gڞ�ł"��*T�`�	���V�-�KU�B��s*���K�Z����ZT�*V��-����[ekZŬ���b��Z���jۤ��2��a��ilTd��-J�
�[A�m��±T��Q�#1��ƃJ#�TplE"���KV�-�r��R��҆f2�֔`��V�mh�laXeH5���SqҢԪk��-��-hTZU\�\�HҪ��\�cjѴFV"*�*)F*�Z�R�-+eZR�+U.6.5�K����j�E*TZ�SVS-�ۉ����\j9K2�m�D��l�YjR�b"�Z�2��%kaR啭b�cG+kS-eT�����4U���#�#Zc.[�2�ش�b�,��TF�,��
�UcJ�[j-�,�r�.9#ZV�ʋQ`�qL���q�b�kn8V�kQUm��mDQ��70��*���EA��@�vKR�;�,t��c���� �)�#����g7bzh8�9	7���t
�^�c7��)$�ޗ�|�똳�T��9���m��垶sm-�Qm-�,'C��f\>�4�[A��˖�>g+��H�H�nk���]C�oWo�ې�E��q�U��R��&�}��Kų��~�[r��y��,Q�&g(y9|��ٞ����@�::������KG�GSٗ�`�f�h<����;]v�pK�
�C�M^�F+��%��5��Xd^�6;�\�'H����-���_���W��eꂂ��uE�wa�?[�[�oz�ݺ��ӈ;V6Q"Fm�܏k��k���tu>kR`����314��dx����.N^�"���O/\�}B���R��Ks�l�z��F�o�X��v}B��Q(ln��(y��g�<�[�2��u�9��{���Ջ2+�p[�v]��l��K�E�ע�>W��ԋ<�r���E�ճIeř/%������#��O�ޯHj΃>ߦ]�q��4Y�v]m������pC�C�d폕�V��h�M>�)+r�9���)5�JG�f]Ï���e�����ݓ�q�k�qJ�HP
՜���c(�}]�w����4��ws���.���{S���$VZ[�g�߫��Y�0��z�=�پ�ZT��xJ�4&ә6D]sۤI�}{�0*gvFx9��{K���s���һ��\�=Z�^�Ks�����z]%k��r�~W�ԕ{�A���ؽ'm��d+��U�#㷚�x�}��yT��c��-��������[�םBH�&[ҫR����4��۵�!�����}[5ײ#E�R��ϪX�c�|�ڑ{��^:����t}i:�)��w�;Բ����W���� �5e�]`,j�������lP^�{v��x(c�+}�e���7��ZC��O:dzL�;e.�wp8�Mߎ��O���z�Ms��{S��f�<p`3�Me2WNfC�S���{�{#r���i��`|C>�1�u{Ζ�}ջ�[꧌
����H�Wyъ���Fe?-��"Ȅ�*��dC����L=�K��IR�%�Kʎ�J�����x��H��hO,�L��w�g��<�N^���FL�`��S�Vq���<8],-G��ܥ\^];L�w.j���G�:љ6�+6�v>�'8��oI�\�9�{������Z<�#ő��\��B�;}i�N�����r�Ac_S�9q:��o���玡�ܰ��ߖ�m!e��[��oG45�e�n�̘+CY(�(�D��%�U5�U�N����F�����V�����;h�X�ۜ�����
P�Vk:.�7i�Yn�[��8\�$R-N�����G3���8#�{�fJ������e��0�5Α&�#���
+�4���I]�4��<3�GGr�*<<��~ ��IS߆L�L�0�5�JM+�du-���&�5��eR���wD,����7�ufmdYS&�.ǌ�R�%	���$ۡ��t�6�5�g�-\):��k�����:X��h���á�lR#�ܔ���eG�r���߹���t~��6 S��WmPgm_���;��ʬ�4��>U� O^�q��ڦ��پ�!X��"-�N�+m�5Ҷ�!��Qn��
ߒ{G�g��v
�[݃p�n��Y����h��`�ǰ�^�E/�ۯ	�-�J�xd�.����3ۘ���\�!6�q�z[xq�b|&Xְ�~r�Y7��v�x�Ӄ�ݥ�ڕ��a)�K�4D�r��&N�=��̀���� ڡ�:�axw��y{}r�)��n��nt%�u5����դw+Z���Gθ�K�n��N^̧��0��W��Ҵ��!��K�}��4���Et���<X��^�C��(��F�A]*t��sz���(�Pa�;�/����j��N9�Y"���[گ[{�zǂ(
ok�l��k�r�%|vS�&P3y�����W����M4�dh|�#ᰒ���/��=6����/GF^W�/Z���L�vq#�=5"^��S�O�=��x�M��p_aW{c�C�v��Yk����6GRv)P�U�i_�MC7�0�z�Q��Y�NQ��,ϥs��z
�Y�OZ.U"΅Ƹx��#��T;�u�iUPs:�d={��z�f�lW�da0�Nx(�[�] �{�Z,��DӔ�x���X!ͭ����"o&���3����z�:�bz�N��s�Z���˩c�o�3;�s��ý��p���������{�k:ܣ_EaI���p�&�%LB�r�)a�1��Vg�}�d׷7b�q�ZW[\]�C�������x���WP��히JZ��Gv�ݽg�yz���՛^���2%%Ii!�W>y��2�9�lVy�U{�'Iѵ�z�3��r�W�鏟�V"c��Q�C���m�4%��WI���w"���ɒ�צ��;w�V����L�=��UJ��g��6����;GMY��C\����	gY��4�d�ŁT�g����we�Y\�b���Փ� {g��U�ia=X"{�*�l�������Փh�3��S�7��`�8����\�R�b��haD��t�&�줥��h�� 
��:���l�o���{���w,�3l�#w�o[]�J�oZ��ge����5�ﵝ^��Wb�,rX�=��ȼY���sn8F���S�[��y��\K�\iٽPL�}�f0;׸�>+���X���ɵ�/5i�75��o}�Cms�w���$i��Ӛ:l��e�3U4te�v^��K�7�e��w.���M���e̹�7k�����J��)qj�B�E`w�Y`��q&�0s0��R�׶�F��y�6�n��A������v����
[h�$#@�2�8;M2�Ug!{Ȥgz�7��&���q�K�L�:�����z�xm���΅��,gґC��LP�⏫C�Gf�>|��F³�O��i��y�0�jr�r��킇�3�|8]R�pGH���*+������bil��wg1����F3��������SW��1X��%�� �,3[O�����D���;�	:Jyb��қ���
�|�0���uA�����!�����c�׭xD�aEO=��ԗVΌ_9��r/��^�n���Ө^
��Қ�l�8���vә��sXt�q�;�b�״Ӭ�E�z�V�e���g6�VXw�v�ms����W�����g�m��][)[p���r�
����}c;ΰ�
�2;>3����7Wu���ȿ�Ķ8%0��Ul'�*�L�g���1.��j|x�g���\{�2uNT_[�8���O[��{ۮ�(߃�Ak5�\�`)����61��C9cY��d`�oQחؓ؎�~v��ʘ���8.\;�e�̓d���\U�N.���>W�5"��u��o��xv���xqR�}b�j��z�!�:1Cؙva��H�+a#�<ѽ�f=F�r)-��G�6]z���M\�$�V�������ђZ:ne�/�*���t�Ձb��툺�t��E/Ӧw���ޡ����.����r�֥��r��h|x���=>6O���>#:���]�+��E��D��n'����N����_/ )mK�zީ��0��g{xM�W��Pͯ�!<�5綥��[V9�"��u�ò���¨�^�v��������AiQ���8&���Ҹ����t�--�ةcU�2�"�a�`�'�5�T�ٵ#.e��	w1i'���.��zwW��67Bc��c>�xa>���e�,�c�1.+2:��x@�͢�X)��s2}�-ꅘ}�O`�n
�xo�iZ{�V:}�t/�O��[=��ޔ���Lyt�xKX���i��i����v���;b9
���g��GH��ܖM��rL�f�X������bΩvQC�ޚ���'^��@���{i
٪�]ǘWG�k��u�Ău,��,�Q��:���$^��>�nɮ�P��H�Wyъ̝B3)�o�X�YD'�:���a�y�_�r!���2��&
U�`�v^;�98ОX=(�c�
���XU{�݆̅��+277�������_$��l%�L��qyt�3�ܹ�Ҷ���FF�VP�-m]G�����27�6at�l����@���I�k`e��p;w5zq�b/{�b�+���m��P���?{�����%��2Ɇ��h��~���FxrqM�mn�d�/Ӕ�����/�����K� ��/��1mܸl�
e#JM+�G����{�nW9��J8�����W�m\X*d��"�2%K�D�',C]�|���'׵u���]v=<��J}:��X)�V*��
Ϣ�=ֹa��t�����2탒R#�����Tk+���X�"�;���G���V�$�u�}e���yt�pL���m�3y�>�MT������'�{���D�5��R>��U��K{·�`�c�긪KT��Ep����Ae�
�Vݡq�u��:��C�����}��U�6(�_"�:��+NR��Vpcv�ξR��9:�r��@���h�ӫz��%��Er�,�Kf�i��,�p�\�5╴7.��^�T;3GJf�W�[ICb����؈f9&�{^������4f�h�^/R��_z�b��:��0U3�ב
)£OWMK��>bJ���B:���?�����o k�o\��v�}�^�+q�/�10ye�gV`/��ܓ���9��}&�/k��j�E�����M+���Y�^��/�^Ė�����^���RupUB�`�ZU�2Y5�jD|�$��ĻV] ���^�G�v.�{�i�|�%�"n����ו�Ȧ���E+�ܦaN$wΤKҡM���=��Us.!ۮϠ����MK+�ެL��gՖ�Mo�:��T6`����K~zj��]I]	�e�7��ԉ�%�,��;.�{S����l.5��K�v#��r�r����6v�f\�'��+���_.4��ڢ��8&͊�����;4M4u+K$���yk��L��xm�Tg*j���hV�C=��-t�B2�\�ذ<4ˤ��z7AO_v����z5�.JU��@�<��u�X�}��S���9H�U��i��z�qr�^�[�$g� ��� E���5�7�n�B�)�|2ݦ� ���e���"��>H��]cd�ٔ/v{	��y�t�V��yS�nG}�:S�r���h��֡=����-8�=��ڍ����P�C�q�^���͈o��Xҹ�����!�w)׏�۷n��h�.fZjF%�N�w�p�����������ֳ�yp�Ev�Q����S7:�۱!���״=����B.��KI
�Y�J�:�/�=~��8J�Gb�y�vPz�gF'���vGT��2��9􆞣��%Q�$W�Ҳ!���{��
t���ɮ�-�m�2T��#XGI
W�ܑYό���!��`���
�o����L�{��]�F��e�f�sW�[μju؆oK��Ab���8Y��#���ۇ�0�*�qf��]�����}3�X=��ۙ�޽��åqAcM.��<����_�w�at�5��Z�~A�z�r5�~���yX������k����0IvF�ی�1�<a����m�uٕUG}���7EE�fB��G�}w"��Ƭ�p-.%���*�}���5��s��]��KP�6\����v�l�Ŕ��-^�m�Pcؕq��u�K՜��<��R�(xRǎN���z��+-O�%�S�Z*�x����n��V;j®b���u�>���w5�]E��Hs[ԨU��IL��w���/j!�m��-۾F�(8�U��Q��Y�M�R�SG;Y�[��#�E&�m�V�7ۖ�#-m^]�`/�	����̽3�P�tS!eo�9�~.���8��kZ,_�3��QE�za0�S�8��l=ٳ�eڬ7�{T&/<�K��z�SȚs�S:i�nM�l�I&v�!���Ƈ�����1^G�-B9�`l,��y^�3���J��R��#�<��L��v^v����ͭ6���;�z����v�n����wYy���C�O�Q#�R9D�]L�)�c)�-��q?[��R���ת1�:;7i��Io��$��~�o l������>�L����61��B̫�*�32Iu9��~����<�fx�Ե��ȯQ�r��tK:l���qH���]���{e��/��� �̎�t���RJQg9b�|�dA�˷�������X~4�|Y�2���Q��U`B�	�����]Ak�e���u&��邒��B*��`���Z0Ih�U���ǯ����z+��4����Q#g�{���~��<^���t���r�Ŝ��Z��'�k{�}0��S�sz��R������Z��4��q1�Io�xem�Ȩ~���w���8;��~z�0�q�7V5�d-l���Z�̷s��̉x���~�&{1f�G����pk��D�lrv��0{�	{����OE���!��u�.���c�_"���p�������tlk]^����EĢ���洊d�h�}K�0ɷ����ƺ΄�yIM����D���I��|U@5Q�8L�b�\��u��(n�4%��.���5م4���B���^��ln���ފA�w}�7�-�1l�;��)X�;���-�ml��
��m2<IÐ#m��M�3+mP��2���@ɥ0=õ.��YgԼ$�w2m�ԔV�d��wj"CE��k̕sdֳ���G�L�:�3ø�V�t&�P�'Ћ��A�K���c�C�mS��E�}�����7�8Nƣ�-�.�ɼ���-۟m�,g.��a����U�_�����ĮpB��'�<9<�n��0:���)O/��q���L�A[�rk����u
vl�8�{��w���>�U�L3&ܝO����ң��ۃ�V��
9�Eչ3΄'��vܗG��m]�xj�͞����)kKIr.����R���¸��"����J��-6�n��y��V��`����?P����M������΋=fϹ��6ѿk�0�v���3�q���OxnV�m������0�o�<\5�[��8G;f��t�R�� ���i�Wu��5�R�)Ԣ-��W�;y��O�
��>�S�K>�wV�n�#��&��7���-!i�U8v��<3	�\R��k,,F���[�WO���R�˾��C*��|�N_1϶�]��.䠔e.�ŏ�muY�ۡ�O�����'o�p�����L���+��zm���o��zmx�հ��h�ۡ��y��s�&�n�x] ���Ƴ�5�[9B[{��W6���d�	��f2�&+.�qԇk���	�5�����xH"CקYs���B\1I�Z�� �d�����JͦqB#�	O</���>��U�7Vͻ���Ա$ Q� �r�N0#ڸw;)�Hs<�[�	�O��v�{���6s�t��C )��{����#7LTKN	��t{Y�;R�OpY��ɛ���bɂ�p�"�؊���B�rv�l8%	;�5�v�wr叾��5��V���s�GV/��/.�"iл[5����Wj�q6�^��{W;��B�Pi��p�8��ᮂ��$~�r���ɓ�jk[Jă6�������av��E�S�Y�P�'��e�c1e�*)w��xc�G%'����4�OI4z��(�x��V�J�T�3��|ނ��YW�V^�]v-�� lL � (81}��[�]7�� ^�o���#�˧���epB��*��S��c��>��e�K�]1�~~m��8EQ%�$��7)aUR���K��S&-���A��Z��ESMA�`�
��ډ**�ڊ1"5�ҵ�CfV*��`��-+h��\̥��AKB�T�(�m�QF�cj"ҥ�鹧1+�Y�*�\Y�SV�J��b��bZR�Qb�F�C,JT���R.���J5�-��Y2�1(�T��K[m�2�LK�� �0��)muk�[��M1J�5b�L���b�Z�+Lj�5-�Z�P�T-hU�k��+*�(����P̱WLq�ʨ�#KDYmKeAUJR*�b�c��H�F�*��k*6#��T�t��ٍ�-�TYF�
%�TaV��-�Z�F)
��E�q��kK��\J��1��j6ȍJ7M�"�������TUm13̢�YUD.9R�����e��T*V�{8�%�-Pz��[%g��N��ct�Հ�
��9 w���ǹ�3^>P�
'�#�.�|ic0+ԧ�v�xO'��D�x�@�.�w��c������g�VI�dz�
��r��Lrʯ���G��ܸ�'?�q>Vt��c�f���a}=��v݌��og��߲�"{�D��V�*����t�h0D7��l�ws��~LM��u��)�x��5e���'���Ϊ��z�vԚ_E~-(#+p�`���b�2]NfC�S�D�;�,B=¬�J˂���F�U~��yDp��zbKG����/ m�-��ΌBN�85-���,o.�zo�!��a�݇c0Sͨ��?<~������n�D�҄ō���
�����|n�z�:�d�_+0���s��Qh$��Iئ�U��Ӵ�r�	[p�>�X�ޖe��-�ͮ�i�}�ͽ��qB�X��G�ݠEF�A-��V�Y��9��<�L���g(��;4J��\���>OK�Y�Kg3�L6&'�D�����8f�{��0ז�D�S馆�g|�S�5�W�>2��H��_d�p��*e#�[�����nԻ%ɉ˽�e����H��� �.+n��<�s4�v92�B���A���i�Y��cv�q���u��V�xrw�0�ZsΞ�3լ�|��rpw�T�ň�����~n�w}s ��\�3��f����}�6���1<��l��q�N��!�~��uԾ�͉c}gVj������aߤ�kF	,NN�������+�]��-�z�"J���f.Z)4�k,_��׬�Û��&a��2���q���=\Zy�w��<��z%��v&w�$���yh����	�qp��}��@�e�L�z�s�j��[�L�hn�`p�$ƅ����8�����ei�I��1e�7��s�a.�����p(�bu�h��c�p�^�"4z�b�kk�T����v�>�y�o���z�w-�O<��f�|�v(6�z.���9M.}l�h�8�i�ǳ�Z�M���~CަTw�o��4��ԯ%Ca�� 5������K��N&��K��<�ӴI2���u���#����x��+J��Y5�jDs���Nm�3 �/fS�����o,�����]�EI�u_J�Iϊ=!=<�^:_{!b`���N$p=5"Y�p��x��,�W�{pګ�Ҟ�+l9�U�hl<��f&f}Yk����I�Ԩl�w�1�z�L	� ��l��p</�owCݤ��W\���cʶR�ہ���u2�*��=��xg��b�R���<ΰI��yj�<V�gV�V�iu����_����y�(^��y~�+_<��뽭d	^��v_p7`,��W'�T��Yv��C��z�MoY�y���Z=�G20�d���[��A[�OZ/%�,��p6�����O}��TJw����_e��]�.	sY��(f�a��b�+{� L���E��h�r�#���:�F��/kFΘ�_s�=e���'HN�oɥ�ɞ���瞵qB.�\�؝�ϨT��/1�n�[�'E�d�M$��[�ȯ���t���C�'��4��a���i*C�_�F�,k=��<P<:�Z��H���N�w�p������[�*����%�W��ݓ��� �%���\�B]td�Y�i-r��>o�]���J�Gbs�/zV���wUM�cy�m�X��O3�h����b�D�"d�8.��@�3�Dx�Y3A�E�c�oZ��poL��H��I��CORτv��,!���?�Z��Ϯ9��P����g�$�4���[f�V�v��&�`�^,��#�oj���(N3u�s����� +D�܄>�W�./�'���Z��Z��u�Ք�� �狄���:h�%�o~5�ԲqS�g�RL���X�gw0��sI��쬜K�}A�OJ������POo-�!�0�&ڵ�T���[�SO���f����R����Y��h�%='�!]#��S��Jk�/��k�G��%�,��o���J+$:����2�U�	�Z�k��-��ǣ\6����Wx����~>��Ӵ�O���.ޞ�70���r���R���ujW
\E�dy]H��xՖ}�Ĭ�M3+}�W�w_��z��u��凨d�s��z�ܫ�p�l�Ŕ�п��������NlmK�Y��"�;A���c�k���X����z�~�܇�Yh�x�1/R�}̝���/X�x���!x ��e�oiEL&NP�+�`��͞�,]R�p5:�*{�{Z'����� ��I-=I�u�e22)��S#얼"�l�/�V����+/w��GFGv��R=��"�	�c�n�2)�[�x�)�o8U�����~�=s[���-q�(�,K���y2�
fbiM���q?[������.R��ڹ	�o��ّH���I���2[ņ���AY���\�`�L����;�)�%
���vsj���<♞=�O��^��.ɖK6�t�	`_xM�Ĥ1y>/;���{/��M��kiY��v <�T�ݡ�Y��]w\6V�Ca΅A�T�R���6(%�w=4����>Kjlӹ��v��MƵu���x��̚��ds��p�A<�uX۠l��0"����m��z�ޣ���%���w��S�:\�9���+"�]�^�՝���]�q��9�٦���k�lE��n���)2��>~�3������I8��f0dI�R>=/ZyU�����H�<E���F�ϼ�����{۞/z�ڇ>ޗIX��,0U�u�q��_����x����A9.�7�:ѳ� L5�yT�T��%�bg��x���g�_��$���jR�7�����jI|I�[ҽw,��?]x�8�U�sY���X+��e�ǒ�X�w�)&ߓ��< /K�"������7W�J��g`Ӄt՗���̩cS�8��ʬwqk��<���w��kP`ܶf ��->.'�&˄o�/N�W��U����,��nv��qe'+s/�`TXr�M<�i�c:�Q&C�9v���x��{�O`�m����Ǚ6ާ,ʽ��:'Y�VZ,��,�$�zS�V�� u��l�tb�d�Rޮ��>Y8�o�"^�U�{�$�����4�������U��˲��ȑ�P��zQ3�G^l6�6�pkI�1J��a���A��g "��a��4b��|��{�}76�T(�H�V�����v���}��v-�G��
�\�i~����|��`��Qxv�n��y�	�֐կ�=��z'y]��8���Q�Ї8f�"�vI�����m�z������QIih$�Q���\z�?-۬w������wlb��#$����������.�l����Wő���sR*U����eS����6C�۝郖�y@��:�U�"�����d���-�ϦY0��a�k�"KK�L����0��zE��!C�^3Bb�O��0k2�|e��*b��ɐ��0T=��yn�+h�L�m����ɻ���.�iL6���Y�A�}S&�ǎ	)Z��\~#0i��pl����u�x��ne��d'��g��:��z3���5.u!��$�x_T}c��ǹ���X<�#���wT�֒g���\s��u�2�.Cp����Cz�'���z_��篣|��]�d�t#D܆�&�����:��a�ͥ�})����I�9N��/�9�s$}n�z�q����u@h�{#�/�GH�������u{V3=�;�[���#��ٯ@�S&����B:�;O�߽A��g<����nݫ�歉%�uh������=��\�c�x�qd����`{��c8�V�d3,�V�їN ��=�� �8ʚӊK0�Q&��<1�9�>�3�zn2ܸ�݅Elt�J�~���dxY#Rv9uԋz�^8�ǽ��'V�]3� yi�J�dKF%�C��� >��A�n�D�]�o��Ұ'��܍m]ޒ�����f㬺�����Q��*�e�D�z�`3��)ϼ�$��30S��_�FLZT�ly���������~5aІ�Ժ���(�qV�,vq#�MH��_lf"�n蛓��>5�I[�'������Ud�I�����l}�����|� G��{r�������כ�+V��q�^��xL��ƘZ�oS�����)��l.5��K�uEC؋.��񙈭���[Tۙώ�37e��'<r�oz���h�(�t��{C�|V��WW&ʋ�r ��>Aa����x:�i�ߏGB�Ny�W"�`�\�Ot���Y6�-xg��4�Q+����}A2/��C��|�C�I�a�"�%-9"{�e�l�{�	
���<Gm
�Z��-$�.�]��������x��՘��ԫ���,M��k<XKO���@p\�E�,P�ZHk+���댼����Vj���
�+פD��F2��I�J�G��<X*�b�ku�@��X�3��uc����{��~|W�g�9y���C�6�����"w`�ő�Ϭx��(�s�����w��Gx�������:�T�U�J��pݵ���O���,�>������y��-Yʶ��QqLP��V�2��	B�"B�tW���/�{N0mw�.�:l*��/{��4 :�wW�7�
V��i�!O�GH��G��q=z�n�;�eV��L���.9��g3%�O�v!�zX���X�{1��x��>��rԿ���G�:�nw�|A�xAP[�^#:�G[��>�8��������������Vvc��>�c��a��c�+-b5���[G��eU���j��e���8�J��P0^����1Q��l��\���ܰL�X5jW<Ex&G���;Ƭ�imt ��C:�ȑ��w����\7�~�g�Xz�	��uh��uU#gf�,�����ힴ��Ú�1�?
�}^�h"|�]�s��LŴ�N�(|�X���~[3���Yh�aq�2�F-Z�v��G��(��z�&�J�"�
���_�iE��59C�����ol��f���7K�4:����������ѼeUW�TG_]�V|��SW��J+��%��f��Lt��}�)���u/v
��hK���-��`�0C{ك���J����ǌXKC���c#�r�f{��x8�m�M��)��>����;���Ӱq��Y�����=3(̧�Or\�r��Z=L��o��8���*p����O9�
ʗO��z�\�JG�<\[A3/�we�wa��;�'�;}Z��\�[��;��'����d�׭z �^�$K�\�Z����̱�Җ����l�4����u��<>����/���a��3����`6C��B�j%R�
g�[��gq���y~˓����Ϫ��rƳ.���b��dW��p�	�K6�B�K�s��W���>%��|�Zwؑ{J�cKU�s��ȃ��]�^����2���c.mz�U{�(����I�wX-3C/ׅ��֢�ޘ)+ʄT�l��b%��l���y����1�.�F�i���ܧ�����X��Xτ��D��:.��`9�xd�G;��xа`W�j^���ܻ��a�}��L�s��%�Yᕸ��U����cz)0�c��^zt7x�*�wn�c�lHf��Є�C~��~��%^xs�Շ��-�bI)T�H�z^:��p	�gN=����ޕǺ�Ռ�	��%�2�w�ř�(��+�A��nw�d5�Si̴)ظʛ���@u})�r����mumEqV�b\��.���7����suwۼ$��ގ�F�N �m�]���yY]�N��D
ز>J���s�y��e�ff�v��-S���մ���G*�����
���`j	a�[�탟r�T����`�.�/N���ƴ�Id�c��Vb�>�u���Yq\��)��J�AB�a���E��#�\���뼠��w����}�@��غ頬q����p?r,��,�$�zS�}�/ l}ޤ[+>��d�8\�T��"?�.�y�y� �Oմ�?~¼s*�`>)<~��<�|�n��ݐ�Q��lx|��a����Lw{�y�Y~��]Y��6Dq�M-�ئ
U��N�7ٜl�=	�8���PJۄ{ϭy7:+>��<o�j�z���ݠ~dh8�5=�ՏD���1嫻b=��}k�T���mî*#���a����-�ɖL6&'T��d����ۄ�fsZ�&��s^�8�w��uD�3*�iC�yzw������W��ɋ}��Ga��H�t�V*�K�w��c5�2b����u��V�^O���j���ٳj��t����L��}ґ~3�墓K������,no4H���9m����m��]�3 �M.�r�x��Dad]�4�ew ����n�^v��`3���K�A�]\C��n�(��Im^j�6`�F�ޮ\۳�.r$_r;B#�;V��Ek��_1Q��c=eзh�uz�N�VC47�T�-eݹ��Zi>�����9.��F�PRo<Ƙ熞#,����3�k��6�&=�:�Aؙ��&����FT]/�,B}1���,�Jy�۸���I��4��׋Mu�6���OX�+hp4!5FzS�w8Nuu�P�d�p�ͺ�Q�Ts�hW\��ʍ��k�
�����Nٴ{,qF�ՑIl�], �t��w0�_gm�Z}#
ʘ~�����ِ���#Au	ڂZ�lwI1J�1��r�u�4ە+�k�䦁Y�--�@�=�Um*�q��σ9Q+fa��`J��f��:�75��z
�#�����v'�׉�s��n��Uto���>pz�%��N�]��Η.�K�՗b�-�tNu���e2$���rf����Z��(�1_a*�����I���]J�yۤ�(ʬhL��c���!)����+�ϳxMl^fZK	z���jo"U���_��(9�g}��)�!=Z�L���W�T/�\��$�لP=�+C�.�i��X2Q)m�EG�d5o6�xi=[P�S� f1v!����eBŅ�t�:A��.�[]Co��3[\t�8
ևt�H=E.<V�ڍ>���2�Xa�ΰG���9ޫ�HN�6�V2%J����9<]s��q�M��F��������Y��jQq��4r|:��������l�i>��80�����V���v��W��'Cc��'/��J�FjjtՐ��vt���4"z�y�A�js�X�����i�s(B�=-jo��E�>~TgΦ=�F+�˘�a�{*>Z�4U����ʹ��}K/��p�����������;;{y�v�j��M�T�)�x$�8'�p`_fGq�ĥ�0��3����S����ε��j�f�<�i[��/z���b������(�˛�o|�d��8�lJ6i���K �B\A�/�k�����KZ��,��F(o�6'2�HK�н2�˝{�jħ�\]�R��V���nZ縚�qD`�x_>�7�ׅ����7�]��}�8����DG��oN+m�5:%��wv[���1�N�-���W ��g�����������j�
$Y�����f"�̇k�A��b��a��`[�p�.��\���f�F�]�k��kC3p3���ɭN۶J}wָZ�r�P�_�T}�)�h@��u5]B�&���3�ZNE���p���8���D�iii��O	��߁�#�+s�2�Ś�X;|�î���z�39��K�iX�7hnGlG��{�8�=��	����/��49���LF�(��⧗fn}��C#N�S�zz�O8=�{n�>��ͽ�HI��4�o�(�F
־Z�-�V+*�m*\(c�+jhcZ��R�mQAJ�F�Ab������*��m)jP��jT���1�VѥJ�%H����������*5M`c�s,���TR�V�Yl�e3XT�5h�c�P���*�X�m�V�\�R�j���q�eAT��
E���"�*��Z,Dr�)P�[L����e[[b�3-�fbe�Z�k�6&��*"5
��89ff\ȩ��p�
%L���Pr�G�꘺4fcAˉ��J�[��[5j����a���6�i���Db�-0m�c�k���+���K(��-Qű�m�c,Zeĭ�YU2������3)T��K[Ŷ���9\��ƹr�r��i�0��c�kAS-Z��6�l��b�J�N8�QD�E�-���iD��V[EEUF���iR�U�Zŭ�LnPJQ-�kYuL�V ��m*�b���KMe(QZ����QVҶ�[Lf����1EiKj ֢�1V�У~>���=����Tf���%W0Nɽ
� ��ǈ73�;����^Y��A��*�
j��V��eζ�.�yH�o�r��z����]�8$�G��$������M�I�����^Z/-���w�98��*��c�'�:��⦧��tUΘM[�&���$��>��L�^A��[�*P��Ǣ���et��gtWm	&�ƶ�Z���}P/ӭ����Q�#}~����dnʃ15��k��K=��{Ǽ���<i��+�5֘cr�ņ@����ɾ�{�	c�늯��+2o��!ꓚ���/j̪�Rȡy�p/k��ݎ� w	�}��uT�*�N��'L�Â�sS͉�=^Se��7J�Cs�1_�5��ŌvMv�:�	/n��Kt9�����Z:���|���7]�VF�M#�S���N$w�$�]��n�mf��9Z�r����#*?Pc`�jό����\��4���N�P�O��=�p䥛��ӵ��هZ�_i�f�l�e��4Î�c�t��e"�]���UZ��h��v�Pz��n����$��-ݎ�v����0�o��Q����AL��؋;�2�-�^x�Q��g{�R�ۙy���/{�%x�f���%�9yǮ���j�ԭv�:� k.�tBxw��qb�˷ݶmm1ܳݒ�����X��8��uy�..��"5=��~��;�*�r{�˂��>���>s�xA�������/��g���U�r��&��2͠�au �u�z�S��;�VV�h�u�ظ�!E��}y��5�j	���$t��T�k(.���[�R�/�t�;v��[#��6�{o���S�1
9n�,�(;yh�H���B�.���	v�/E�qx;���zU�_��~X��/.�Wl��	k��r�,P�ZHV�\�k���[����/�2�ᄯd���)_�)<�k�1��(^|e[D䆞���;J�!����]�r�x,���Ś5�4��f���C/ך�5�����J���i�bCORϣ�v³E�wc˭;�]{ދ����)C�X;)���3�o:�C ޖ9'�P�f0p�YԷ7����� �sf�#Fnu�.�o�L���=i��u��2}~u�=W�iAcd'REj�Z{�.���8hw�A __�v���WO�|V���X���?����q��������K�⣶�*>ڜ�o����ǷBk����w)}^;�R��R�,�<�wǐ�V3E���ϼ^r���{���G�i'OS�Ϛ�P��|�
��-�����a��@9Hv��m�=I�<M�k�"<bû�[k��r��Lޚ}We3r��3r����pmN]D�%��7�(��������j�j��N�0�m:�_gB��/��r�ګ����f�K���a�6\�w]����$}Hi�~��תv�;j+��t΋�-O�p#�z�v�e�a�t�r���:�~��s���(����^wc��"��mJ��z}U-<��"�
}Lĭ�(�Ͻ0�Y�����hx�����p�D]en���q�Ǒ1�a�GJ.,��3���m���覯}:�Y]�Tfeݫ�//_��u�A�b�"l�c��v����W
	�x��ϻv�
�9�Y]�7��,���Ib���
2H���Sk-B:��D�b]�x�����̰2�Q���q�Ƽ��4��Z�XG��y7R����<}�fq���`6t_k5�K��a&Ko��i�����,��y�zxQ6�^�K�s��;�rƿ3<x5-x�^���ù��%�6I����^�IM���_|��o�Y�����y,�L�n
2+�1*��2��O�0�b߯n��ͨ}woXh�,��i �+��ˬ����x[�Q[�%*W&c���<i��������.��.��|u<9`,gp�֮�k�:m��Ns�r�Z5��z�gD���q84ᚥ�h𡡟r�^]p�q󧳎퍻\
�Gp�_>�Ge8�2����Tk���K���\F�+mc�U�] �C�
[�Q��6�[Ĥ�%wty�]-7�˸p?R��H�@�ؽ�\�l�*��2��Y�=��c�+Ԧ�+�t1��tǣc�0.t4�r�֥^]��~�l�j��<�\��R[��>������ٺz<>�h�(is��X�Ce�+��r�α0o�yC��j̩c�N{��=9�o�bM�/��*�P5KG�/��o�(uߏg�m�?v��YIO->ٲ�J����Lׁv�5�r;O�5�sN
��,B+���prt�uR׌��d�p���Ӻ��鞽I]-��93��x�xz��c'�c>�%��AC����΢�I���9��T��X����.+�C�Ž�]����+"a��q}���Ih��~`-�x �m��;�o�r�R#��i��;s�kv1�|��%.'E�ڌ��.T^�U��v^;�8��WC���w����ڎQ2��;°(w�b�,��a�G�Z���2�qgf�l�lj�⇩v������������dd�h��&�Eg�9��(]��H��v�Y�]=��<�ҭ<�ӏv��[��	��b�U���.i%���L�6cHi�O�v��(/� �;�/v�[>JL�L�֫~
��K�П���H�,����������>{_��v��٣ҕ�K����H2Ŝ��řsk�r,��%�_k�͎������jg��v�ϝ���ۇ\T<G	9��|'��,�L�L�a��ƕ*���+s=к'��ԉ?x�y
+�4)mT'm(�iB���@����P�O��ϱE�K�vs�{Җ��@�T9�i_�L�����l<�Z�v�.,2`z}D]��mD���1�Şi2�}���J�O��,���2��ؗ��<f6��û�x�+�ws�.0�.탟IH�bJ^V��>�I2�!�g�Zj�k���ն
��O����_lֻ�L3Sś���V�F���I��_�*���� �-�~��J�9�'O��%k�i���{G�g�xqV��4^�h��x�Kv�����s�f�DծN���S�z����fU3�ב�n`gەؘۡ�� Zo�9m)�Lfu���~�ii�;~���XCĬ��+�"^L��ν��/�Ez�6:,���nZ��>�T��s���_yｶ���j��}^�z41PA
]���C,����D����8Z�c+�W ����Gu���[��R��&������[�֭����ڍŸ�p��ۛ��={B.um�D�Ү>��E�� ��,ԕY�M�7t�1�!F�дÍ�O;�;�w���f�@���Gr��
k.�7'&�c����{/}�y鮤��m���x�)uw���>�F���ӝ�Ɯ걦�W��{=�-G27:�� 23N%�P��`�T{C�{P�����G��j<�*��M'1r��GtM
���a�q���5�l�fJa�S���:
�Y�OZ/%�,�߲�|��TԽo�TV}�b^#l$D���v;��H{3�fNv(�[ީgYS�f󧴗��e+�t3�b8v�&}:�#Œ����w�\ǫΫZz�joaZ�uN�6H`�H�� ���M���vf���Q$��:	�B��|�OQj���W������'��Y�%f��1
8.Tœ�9Αi_��ywX��	yݛ٢�^X��$3Tq�jW��ŀT˅�+�v!)h5"}-5�Kg�&�a�y=y��	�zyMCz4z�o�����g��eg�]�b��m�Hi�9(C�"!�	�33�vǚ��8�G��۠��=���Y~��b�/��R�"���L
~J�o��ǥASu���q�<\e�b���1�OD�� �^�;/gze����n�.�F���XŊs3�E9ɑq��M���́.�8�n>�F��/*���{����{!��-�|����]W�ۜN�ڲYp p���O޻�<}���eRoh���!�u�:�G�Y�Ww��[λޔ5.}���c}�[����J�3ə3��.�ބ`ǋ�(AF�~��B񡞴��s�Rd����G�ԕ�)��}�9T2�n"�d�b��� �U_�w�2��~k
�>+ppC�������#u��+Pdx�D���f�&^��$�#p=���3�L[��u�өT\)i&G���2���K�ܜ��Ri�0>��Y��K��,=C&˝բz������m������޵I�t�˵F>�<�j
�ٖ���L��a�t�r��:�<p{_a��ד�Eƹ���J7�;��YWO�Vڈ��&��f%oiE}��a��	��h]r ם[��|n�o��r79�3�}Xi��r6
�!-��a)g��:��g[RM��7�+zWsҷ�ȃ��,q��6;��ZG��\\X(&e�/�~C%��{��'�W�HL�zݟu祝�]�7;�z�!�ᲉĻ@����O&^Цd��6=W����	���}��j����
��$9��2�)�rm�u�?z��ٞ�<,����B?�Ooq8R;�s��O>N6�ܗ��<^z����&{��ې,�b�e�Y9�u'$��݁�u��\�`x�L�7xI��Go/m�|���X�	wN&�Kdi�޹�Υ�b.kd��o�-�ύ�@�5�5~V�;r�����zM����q4����9c_���=��b��dW��p�	�K3���)�<�'��<���G�h�iW���o�GVo;{�+"�]�^��P�jhe�\�mwz�Ou�n˳�:+ah�g���U�:�Y�7ґ/�B)i��մ
߱x��y�ǫ�r���^�#�o�WZ6}>�@�p�n|��c����:�ڄ������GÛYӝ裏>)�PI�¹,0o�+�j^�܎U��	]h���P��wt��PY������u��v�;՜�`��Ə���>�M=�I$��+�:�X;:����=}e��O���ѶUeN7s�N�"��ji���x`�e�CgN��_��H9�C;+}��hsٚ���sNAU�>����XdP�7l#b���f`ws�a~SΙ���>JW�jxQ��}��8}]a`uY�1�,�2�J��(v7ȵ�:()��nt���ͅ箊B�DFl��|; ��T:>���k^�0�גJw��s9��J�P�OR����Ն��;t���&���z|��)�x-���o�{v�^
�y}J��k�W����Vƻ�xի88�t��K��q��7�ׅ^�a��g�X������[h��Um���ѓ2=����7h<�[�킇�Cm��+�p��>Z������ŊU�,�Ӫ�V3+�cao�#f��ϼ�bw���t^�S�':��eCA�`�	lS¾#�yq���oД���:��[I�:��^����Fd�謿�s��P�V6z��T�gnt�}��qqK�BL��·n�6�עU�"Ĝ��3%LX�[9��1Vja�~���ţ���a�f�I������b���m�Bv҈v�*+�B��<p�7�=Κ�|��22YH���Z\+Qb�b�x:�S�&*��+V�˾�%�tMyװ8�2%K�&�&
��RK�E��\E_�L��g�G��\�]�ͬ�a'�'��ڥ�	�W�P��˶|$�G��,^.�������O+��q����3O.Gu�^Ϛ�����x�y�o�V�F��!�I��[ʱ3�k�? 5�~|jt��.�A�a:[�N�K�D����vX+= 2�EW�˨��[���a���e[|E�K���-L��9(�j���Zc��wior��[�m%).������m�>О[|�}�c�t�S������l\��D{ʊ6��u��Z��#R�z�����S�ɔY��¶�'��m��;���T���E���,� �s�k��o#��\,�������҇&m�B�ۘ�]i�]E�m��o�Ų���3|�s;K�������ǀ,hh}���P�U��� ��c�gT/<iW�9�<�~~*��i�bz\=�_�����<k�/+���z�`.�0���<E͸�ۛ}~Y#���a��f�.�=>%���~L\]���ƪ�k�!4�R�;�-�a�A��U�
�O���Х�T>��K4Ӊd�ESp?T���yq��U��x�kc.�U��T8bc�p:����*j�,�9I�P�w�f/%�0�vz��=X�3�E����@��"����̣H�a��"GER�koX�37�l�a����[ާ�qu�;�̬��C8漴tϝ�&����+�6C��ԃ���W�uZ��;P��vd@iMo�g�bq���e�:�]lC�YGo�����g�=��=���	!I��B���B��$�	%!$ I?�	!I�HIO�!$ I?�	!I��B���$�	'��IO�H@�p���$�$�	'����$�$�	'��$ I?�	!I�HIO���IO�BH@�zBH@���d�Me�����f�A@��̟\�4�z�  ��$PU@  ((PUP
	 
$D( (� )@�!B�J� 
�U
�F��J%m�
R�J�����T��Z�Um�Z����)]���V$E)*)
�� !SL���bPB6ʨ��H*��R(R��iUR��THʶ��f��+B�"��k)
��%���j��J�M��T�Zh	T�-��I5�
����7��J��clQ�   Z� ����=:� ����d*�vhp�C5�\m�@*eA
��m���g@��SwZ�5.�T�#k��k+LdNڛa*�(PQH�   {{����6ŵ\�n�Zh�Aw5ƅBkbТ�7[��bN��@�6�������1M�)�V�L�E���N�L���^   	��v<(�B�
p�(P�B� �u(P�E��gl�(PQB�
��(�((P8��
(�P�wE�P�B�
(C��;zoN�j����E]��r��\�ڦݭ���*)DJ���T)^   ���V�
�����Uv\�á��we�F��r���T���L� ��p�jPV��:�Tm:��X�ԩ80P�J�Z*� ����  7{m��f�F٠5�\6��N�KT���J�颻jm��M �ls��M���htk@�5-lV�U��պi�Gw-iI	%U�   ^4H�w)Q�f��P+s�u*���v�fu�٨�Uӎښ��gn�[d뎠���q�δ� l+
5EY2T)!mI���c�  � o1ݍ!�v�hi-�ڱ�����T յ��R�`Q�1��l5YlV[j�5n��С�]�6�Q��Z�Ă�H�����%%;hѶx   ��١����N��� �̀R�[-P��`U(� T�UJVwS��Wn D%H��FE���(�-�   !�
'�`C������F�0
(6+ J{� Ҳ�[�W ��m ���"IR�U6�QJID�   ����  ��j��� T{���9��Pb�� �:� u�
E�[ o���b��@h �Њx`�)P  ������ )� ����@M E=�h5*�� &�$̪�� �
�R��0k"�i�H���{�����"�#��>|q�=�w�ߵ���}��IO����$ I7!�����$��H@�2B�	�����_坯俊������Gq���*i�E�T7 -��㈞�%�J�J�Tk�Mq����M=�5���N�SJ��{�D���q�ۦ«w v�$�˳���{N�{A�mj��K�r��P��n�׵ma������ v����ܽ������䬓-A�阍]���G.�kE.�fƦn����V-A�V+����A1-���R�Ĺ.m�9��zF�ԇ,�J�;���L��f�֌�V� �0�W�%B�2oCQJ�#D�:�iZ�1]9s ����"a)�C7	:�=*Jmj�oh�Oڥ)�+X��B\)�`Y���j��cNn�r��i�,;ن݁���w�R��v1R�r�[�u��i�X��Xk]r��Kn��77����e�X/��(X�U�b��͔��	��E�fH��,�I�+bzޝ���T�ɵ��*��'Hv�)mp;�K�����O;����2�e���4�م�P��m9g���(���z�X�!��7�F��B��A�ܱ��M���i{�ׅ��׍�ڵ�����h�H/h��)[�(Jor�u܍^Ò��T�
�(Ո��Y�	sM�o$"D58N�4�WZ��Ù(]���-��
7�`x��J����Y����{f�*NJ��S��Fn/Y::]^�����%n" ������^�j¶�/]-&�4f�mn&��kp'{��/6�`L��4XL��Ƶּ��+0'��ā;�s3"��n!-�r�ݬ������fbD��Ŷ.l��[X�s�C:��*�����	��_}�G�F�lu�H�zq������v�9xqcr��r��Se����7jQ�{�,���d����1��h��Mo�� �ie��J�#�]�mEl�ɠa�P��v��0�m��Y&l�0^����0�x�yyB yJ��w,]8�!ݚo6�w%n�I�)�-�tEa�`U��Km�u��i��P��`�b.�DS
�n^s��G�ֻҤ�ۥ�D���֛	f�}�B�t���X͕/6t��>̂���Q�@]�l�Vi�Y{ �G���X��ɗQ��sZyCUԫ!c8t��j���j��Z�:rT�J�ۗ�>��p6�̂ܽ�6إH�+]Ç	1�gf�I<6J�������]](�QDc��:5����*�tV�2^!zt�ZX-2_hI]J���s�.�Ʀv���s�,悷]O�+)�
�϶�)3`8�j��b�Cm�{!��0�P���í�2��؜Mޜn�#A�H-�&�ڎتn�GuDN��Z��u�f�.�Uq���b����-i�d��V�q�f�w���R���y��i������U��7uu�0�L����ӈ)AZ��
�j�
�oiۃ6��n�n��T�[�F�t"��� m�'�d��p�\���	v̚���j�	�;���ιR�;F�b�*�ע��*�u,A�J�5y�ҧ|hV2v�J|x��:)E��yO��c��t�6�a���v;�iVXY��)�F)F�"���\�f@�řz�D����<��l9`٘�����Ҳ�Z�sj���t �q<ُ6�9��ş#W��n�
j�,Xd*eVV[B��2��O.�G/S[zqj�5��̽���h����LLŪ�5�,�W�V �(n���qZ�KqkRb���7*AC$�{�
�n;�r��m/�%���43�&��;�+o���!2*aЩ��-SD��,ɿZ�q�HnW+|k8e2/oS�@�ƕkz+E]�Y���z-�<�ݻ�30��'��fnr���n���a���$�D���o`�G�����³.mLF ��a����&&ڇUn�/,�w�Ah�f�B��Ѡ�oK*�dT/v�ദ:s4"/~��t�rZE���%��)q@P�XòJ����r�#�e�7f�ޤn��ѫ�g4�)#9`@�H�	C� ���dw�^jO�IGkrh�8��*َ�n
y����f'���	Ŗk1+ �v�m��u��ڳR�ə�@�k;ل����F]l`uv��hٖ ���X� �2��%%P�ŷ%�պ��l��2ZQ̢�kU�]+��� �bmފ4��%�:pY�[yX�9t�Q��P}ycE�e!WJ��(͂�Y(�����X�ʼ&A��eS��~VH�nU�#��Թkem+�٨����KaN�4l�=���e$޽���m�"fĵ�z�g��)�Ey6�Ǯʔaû����V5���M�x��
D^r�M�[z��@6��>Kv�d�P�����)��ea!:���	�(!�E���"��3.A�k$����]�&�x憷Be�1�=�v�q��VΪtB�ch6��b#t'l)Zb��߰�ȴ�2$��p��VY/n"���Bf
wEʔ�$��Om[,d���:�Xz���TMo���Fm���+$+0���zA�v��2�Vb���Z՚��ұY�6u���tz�`�4���Ք-�n�g)YA7I�ȷq�v��F6��lY�y�`�ϵ��ݤ�VIWj��wUR������#�s.��F���ཎ�7�昅=��V�p�(���nef���R�kw�Uh��Z[�eaֶ����NU�M��Š���3��c?&�f�]"�f:L!�	��B�Y2�ǎޭsF�N��ަ��Ubܫ��R;J�����`��*W21���:�S�n��T�2��j�5&v�E���ň�r��Ui���LՋO%�)K�I�tH�̤r���>/ �Y\:ʼ���!Z���6����&2�fK9��p�5Q�r����i.�{V2����s���|΅3pid�ӎ]�(fX�l-p0��ՔM;SSx��:��;�5�)��`�8��tfĄ����ay�T�o ںOv�j�-��nU�"Z$U7(�4҇�v�4��/
�++ef8bs76j88]�s(�N�hm<�gm9$�]](Rչ��V���K��"��eQ�]��c6�z��5aa����M�Zj>Y�ԟ:q��:ҙ�[v�Ls26�oc"$ܰ��`g7q&�8��^]-˄�t�d��nm<�X�N)X�o/�@b4���A]֌�`��pI򻢪i�P��AW��F�����>e�q�x�x"M�!r�3��t���2�v��� �sK�^�J��e���[�%%��b�Џwp��bXʈ峥-4]+�T�&a�n%�<�@�}���� ]֒,�o	��L�K<"�U|�^j���D
(<�o6��b�
�"	E�:�V̐���s&n�sZ�Z�ƶ��%K��5����*��ZY���*�W��e���I	�1S�o0��E�f��(4�x��e�lt��L�ٺ�e��H�2K�J�r��!c��T�d��V��e:A��L���������E_o�h�φ� <�3��V2@K��ۤ���Q�ʊ��`V���b�P4Bc5^�ML9���b��6�f�h�w�k	�KpJ,a�(���cN�:��w�����9��dQ۩�+]ef�?^a���c�T���۳-�[���ܺi0lG�l�БysV�����f�m�7`��D����*Ge}�(��U�f�Yy25"z�!��uyr�d7�EZ�j�V;���2�̙��cr��k�(
F^*�V�1+f�1�t�Z0��x���ìZ&���6�h]�J�-��!�.�fpV�M 5���8�&�����̻�R�2�Gb�F�N�@U�D�M'iL��[��(��GB*� ��۹dj!����܏CUp�ڱJ����&���5��k{(�+_kЕu��ٷ}��<�X��q��m�ћY����7�Mջ+�ܺ�F� ��'t��
/��+I�����^�#���a�*�����,%�n��/A�ʈ�4S�f�gUw�k55�Y�I�QØ5Z7]����F�4R��|�3U�Ν�D���1h��/��\��%��M`_\�z0Ϭ����MͶ����b�kkU�HȦ�f�GZ���iv�̡z���[Wr�렉XFĊ���nc� 餲�u��Gk�Nފ�_j�h��D��W� $L��j����74�� ��kS~XP�*��0m�7��r�`�0bY	��qhU g ���jl�7t(Y�VK����ʔ4�佼���.�[���1�E�-⠯�SF��."�)4�L���Wz�#��SpmT����t�1Y�+m&	�b,G��)Qͦ��Ճ�l)G) ���79�9{YO�T5f[�J�{Z�ض�0��X.'����?dX&�=��O>ˣd�xւ�Ʈi�tJt ���eLڙN�Y����P�e�`�T��p�ը֍��˫u��*�&��'t�&�^;ݻ�As��M��i�jZ�{x�9��fE獄un;��;�2�r��v��CY4ȼq=�u�`����aK-r
�`e�R�]Xo�X��^���t����\�o):X��ܩhŅ_5��r,���!��o+Lk7l�RSO�ME*gL�J^�� ���6���1mŻ�h�R?	���b��ɮ�t�N&.o�؃�з4�Ia�渪.PT9��-O2Z���Ej�H�����Tڨ�N�ϱ��6.1&�IFQ�E��I)�yAە*+_mԩ@�%���k�)���]僶�h�[�
��K�����c��yO1Ze\�k%�L��w�K���u��2��`��P�WOV�s!Ե�kG2�����^b,ի%�Y�K����4}�&#ivtK�8�+r��U���xN풲�`/c��USi�d�V��ѿm1��d�x�uv�כm�(Z�7Z�w�w�â��I�̫А�km�KZ5���ħڱ���}�i����FV�-T���ۂ���ݵ�و,�8����v�-yA6�l�f��#�0����ZV��X�fd��6��8�o\�{��n�ŭ�@��2�u�;��.d%���$�"X�V4B;[7=Q,�J&�6镈;�Dl����h�M�ZĶY�Q�*���匚�TA��@DVH���BHp#(V�̆�8A�a2�&4��2��Ss7�`�B�hld��F�Ur��L1U��Zm�f� ��Ù�mՊf�Rk�w��2��g�Q% 񍣌g��+�*��մL�6a��-V��ߤn�;�f�P�A%�̲&"&f<#uݚU��-��5n����F�$�<��D;�#�0��������x3�o!$�qf���ٰT76-���oAՙOA�2��Ԫ��l�yY�:ɝ��$���#����g�.}J��j��Y��qE2P@L��Z�� �Y�r�E.����kK�!qP��U`�Nh`���U��L�	^�����j���ֈp����Wtv�I)�~� �����W5��e:vG`�+8���Ũj����^��U��WE�#q.! It�Ɉ�N�z�Vۼ.��j���V=�z�a4)�
9�P�sdU*J膩-f�����?)*Ȗ�)��2����٧2��4jX�m��@��)�`h�/��[��A9��M���f歼IĞ�0��>��4ɔV+��a��ji�U�*j����R�B���8���pM�JN��/2�mZ�Ș�m#E��T[���ĳ��X?_]�A#C�U�ɢ�n���"�惢�T�g#gmV�4�9���c�ٻ��l��B�wQ4�VC	�ہh���p޼��d�&S�	��KJ�h�;A���y��F�ghA�g�,ۦi^�v��ƹ�cBk���y���[5-�J�,���y �ۅmǉ�;�w*Z�Ze�s7���Ů��e_Wb	��-G�]��m.&��컶[��SW�`��"�`�7EX��tU%k�es�+XcUwiI����a����Ce`��DiZ�,�Lx�JnS�C\�*���+��y������Aз�q�U��B�mWc4Ζ043,�Z�һ ,x�BUEYOk1��;�ʺ�m���U��U��R��i����o�;�d�b�]R�� !0i��T�PC&����HS����ZS0��E�5�eKV��V�8j'P{j݅ti@m� ��9�Msc�i�7�L�p����v�ߦYr�����2I5�)��� H4�G`=�[�S�m����r��{ ��AE<��k�̘���p;�N��F�S�U�U��Jt'�L_]Aq#x��Ԑ,�@Y�k0��]�efb��Dj2f�Z�y�vuE=9BnR�6P�qtҺ;��)��o$D[�y�m�<\G�� x�E۴������yvX�n�*m��˾�O<�����D�Ms+��#HE�-�I��v�Kk0-�<�D<�`em�Ǽ4��5���t�
���ś�d��%��æZ��Xc͈a�ƾ����]v�Uc]�Tƻj�kx�jK+*b4i�O"�q�qC���-Ԧ�Hh��
A0��˘�Გq�)��ۻ�ͫ*Y�)<�J���������Sø�uH̘A�NH-=7�2��J��(:We�{���&w
I�Zh9t���b
�����D�+3D![CAr��V茥�%6�E�	ܩ��hJ̎�V�L6��ӏ���m��om��I40�3>��c�4i�fɘ^�GNټ��pGE�ר�:��e�X�������4S�wk5��t�7Lշ���	�)Q�RH7>�ġ�&f�"�c�)%6����ܮ1�:���RU�X��'_K��90���M��D�3VCSR��xg_7���ͱG9_1��ni
�\����Y4h6����.��TS�^�\�Zh��Q ܝ{��2'���d�K�;d�Z�fvv��\�{P��k<���1,�T����`Vd���+�ma�����,��"�1P��!����X�a9i���ҧ$6u���Z�Pyhh�
��(W�Nf
�1��
�|Wu^`�cީ�g*��K@�esY��@�S�B=!Qg8����� �����e�-��M�1�͠�.�,{ ��#�y-}�����/��RR�#�4F1����e:���u.Sw��&��cm������\�k�P�#�+&���o�������kz��\V�b��_��7rt��2��O���s�*IW��>�8�q�r�n�t�zzk�ˈ�Q�ԛ'���=������ 0���\�����:֠z]b�dN�[6�����8r��7	9$��)�*t�#�f	Elc$�6�]L,�����Ǥh��1c�j����ð����������0�{s��*ʽt�Hu�U]e⒧��6�.��=�	69�\8�ж�3�8@; �B�S��b5�	E�M��,9SE�õլ����
��&���c��(ks-�<gq��ܱ±˃��KV\���w˰e�E����e���b�.�\��ruI�y�m�{׻͜��t�"��D���U�Hl�^7��a���ޛjam�u�9�ޅ`]���i�Cq��A�*9ٺ��%�AOU�w�e��|`p�0mѻ����Moq�yGj�}�����Gb�e9]c��6��	�ng�(놵�}���K���N8Ԇ��ȭH��l� $���0�j��7��������+���މ9��ఫ�-��7[&��^��n�uĳ,��շ��r���J}���Df��4���N��t�+��Qg(����f���+���ls� �<�M�:H�H��ggc�6ݤ:��wZ8r�&kt�P��g��%vFiS�Ұ~#��qWUvdMKCsuW7��,���
x��M�ͮ�����f�Ǵ6�v��not��A�&`�W �f&�ً5v�]8����B�;p���C�zs�캶m�Z���z�̡\�a�QJގ'P��˝��<���{K�88#1�h	�����έX�����t���N�)�z�e7R\�V�L�}bT Z���6�,v3�[:�D��N0t��W�P��9�s���n��� �%[Ig��(�y�p=ʴD�������]���:�h���+ѕ�إq�8�f<�m6�im�ݜ�_&�9��e����ݡ�&8}�E��.�I!�齴�p�z�37)R��ڧ�k<d���p�t�� 	YsH�tޅ�N2M��x�	,5�6��c�x^U�iaȲ,v)�5A��5{C�kP��#w��u�)��H,Փ���0LJ�)3D�¡��j��/\���E�xs��������7����&Er�́�ܺ���n7dZ�ܼ�>��#Zi��X6-�]��Wn��>jf����[�D}���	�a�����0fʽ<�\ĺ
��8ez!�v���:��G*5��ۻ�TɄ�Y˺ �����
ӫ�^�Î9��d�����%OuP* 3B����+N���I��0 �/5�<M�:��m�����p|�Y�-)�=s�J7}��e2u V0�޷�QBʲ�T5n�bc����n�0S={��kqy�b���ƭ�d(�3�>��[k_�1Nypsu�YfB��jͩ�.�O%�L����4���F7������Z�e;��̝�b������G3H��3J���|�K���<�K��[k��8ʆՆi�P��Z�:|M�[���u�Y"�V�=����ox�r�8-���2����5V�K��L-����6N҃�cw�("���U��=~���6B1y�ʷ����5qS[�>�h�L�eES{L���d���6�c����.rL��Gz����+�]�;��nɽA�*(>o�,�b�/%h�;�,+N��|��Fq:��_G�]dqt�,.W0	���xYV����5IВ�G'�ӽ�N���G�le���` �'��Nn�rOT��4�e�<��"�k$���_s�ƥ�̈�S\�^GdX��c~m�nwou�됻��S��(�Q��:�bUd�w���6��Symg���C6s]4W[|Mr�����J��l�l�Z_p�u��/&��۠�k+m��wñ��?k���[�����(�KW�E]��Q�"n����u2;6�ܫ����7$��T����KZ��#yb��fp�$���ab���%���녅������'ea˃JI��	s�ާX��Ӧ�ݞ�4��z��P����.��Y�=ˉ��tZ�Y-�2�]V\vyh�w��q+ЫA�ٴ��뤙�Zx)&��S#���V���TS펽�؀��`���C����jb�X��=�/��LRs�S�)ЦY����n�E��I�X�]Ֆ�Kx��9�h��<$җ��U:�h�E��V�);�݄^�����*�;c7x���ȉ�����9�եz6f�y���I����U�)�u:�ټ�Hh�/3r7��l��n��fI�
c�����8t_L6d��rp�Ǣt{�6�myiq��Q0�ݱG��VU��/S�@����Y��U��YF�;��9��
"袻�2sl���Y|��ah����٪�s,�i����*Ymdy�e� ����ֺ���_X]��k7f?�B	6�b��5�М��֐׋��nef�h@Ėw�.�����`�bҁSf���sd�PZ�*������J�Q�_Zq�|;�WH ��\�����b�|�n撪�wS����Lǎ���6
����Tn�̢�¬:0W�v�pl��v�]�\"]��Db�'�n�h�ז	�]�t�2
Lp�Of����E�T��(�;�V>�J"��Je�XI��Y�N��GJʄ�xjw�F�o㹭e���&�T��k�F�Z��k1�����tS����2������45:.8Q}@�!݀�a�xt1s���v��`�7C�2�rKxS�V8��}9l�q��ױR�ҵ:sk�+�s^N�Q����&;��i,SF6�O������r������4��B|�'�STB�˘s�f��*��.�t]��cq��L�/FI4�� �@;}F�f�mA�ջgn�m����f���V��Ej���b���C�6��};A�bhμC�3:�ۙ�rx���u�ԍ��`�֌�b���Y����]��L�]�s'#۬Ӯ�Ӹ!W���Ǝ�cPc�diw��������k@���7]t��� ���.�S��V;�6e��γɵ��(v�yM7fRV���
[RMYY�r%|9��h|zhyYZK�P�BB֦��]w��{ip7�a�Oj*����`�Y�*�`w�F�&e�Z6i�������8�-Ui�du���Z��W	����ͯj��);x[~��$�9U�=AM�n,�M�Z!�HMϴ��C6���Ĺ>ͣ���G����B���mU��kKPP`|M5C5k�6Wn�d�t�M���c�Sn�g�l�\�-�%���]{-����G*�W���=1E%Mv"���]�9��8G�R����F��ZD�G�,��옜̩Wo-:V	1�jp���p�o�J����̢f.��kh;��`%��kh�o!�;�U֞�d�!����pl�%J(�\j���B��Kmc4Ee�=K2��5�L"�8�|�k�d��ȕu-˺TI{t�Բ[ef�����R�<�j���G�SZh�+J��8ŵu*k��nvӵ��6���.�C8��y�\���W��Ͷ�tlw" o:\��}:�i(0�NY�n���m��]�w���<<fIiJ�6qY<�5�����Ҽ�n�mZ�:{�������"�� 4�Y*�Xv]
荎�:����j�K�O;�u3�Y7��6�.|M�6�����#�ٸT����5r��D�:�/aw�8���'��G�:���v�@ �1�X:����{�ݸ�5y't���y[}Ye�a�M3 �:�o
=<�<V�l��0�Y�%���d�Ԯ�Bڧ�Z�zGm%�&�񗐬P��5�t{e��]J�n��O]c�C��3��&���n+�AW�gR�|�fPU5AtT�Cc*�A�DV����7�r�)�9h��,��x���62F'e��.`��āݬ�n�1��l+#�XBf���K6
��]��l���)�EY ��C�t�k`���^��sBa.�k)s�k� /�gu
���a���\N��,���VuY��fr�r����ө.����2��5��)aLX���7&s����9ᱬEd���)L�h�fi%�0]������Y��O�v��;��9���S<)ʘ��U�[
�*�=�m[�7wn�e�@SUؤ2Id�K7�6��(���9��Vp���/o]> �f���s2��'�l��0�kAZ���`��C+,qOB��j�`u�*��c�xi-wO9��'��Et�E�>�V)�L�FfY��l��u�����*�s]�Y��E�S�\��t_Zzp��5��6�o�W�E�`%d��(���K칆N�C�[nb�Y@o7�.��D۴E���/Y���E4F�f�/(��ދ8�i�T�{^�.������#���͌��G�]j�̙�Xv�{w���b�
��M�ޗ�A�J4yWp^�	{���;���T,7-F�r�|A�<1W}�LLi�@cvI#�oIwJ�d�WU�W�a��F�q�-�SE>5��wTZP�w��&�s��P�j2�����7�:T���KE��f��-�����=�D>�v��cŰ�@�Vړk'mZbSa�l��(�H-U�vKo�ڮ����#�1CY�v��']�	���\�s�*�$��ԝ�&y_60n� u����j��#����Bs֜�o�fU�lz�H�w�t����IS|���ډ����۝��z)�n`�ܐV���rl�vi��ǳeص�Ҍ_7l\�b�Z�&�m�1����Eh�˹NSYNG��&a-�}\�+!����L�/Uk,*�m�Y�d��V����\�Ҏ�3
��b����[�����#��.OB��T�ݳ�]��Ӽ�P57,WaG�����-���
�#׋i�1"ZBV�L���jE�w�ݚ�I�J}I�B��9Gy����$�F�VuP�F���ɯ�%$8ߌ�f�[j����K��^1�����L������[�aGZ����*�V�G�ni1��_q��jT4��'���h�.�%��s�[�א�Ƀw{�q�%���u\�ܠ��W�)��
N�A4G�<pZ���w\��|�r�E�v�c�4�3�%/&]ix�C	�G���e��.�q���X�� TԨ�׌�Tl�e�w�{���n%�Zr�x[��kݣ�蓜��(�K5�:ff�:xY/�t����a���kΰ�Qy;A�c������;/�0�n��]��ym/_���='`�mG��*�B�wf�T����)Q��Z��Ɩ`c G�Q�"ԭ�#��6���e �w�HfҡԥЧ�pϢ���պ�f����ɻ��%=���ʺ���Pu���H����^c�ku��yN�w�l��bWs=J���ɺ����겍��	��l�b����}�Z��h=m�{�8���_�1�.�s3 �wGm3��J�BL��{Xp�8FyX���,�1A�N�V��Ԣp�$r�`��+�U�i2/n:���_���ْ,��[��D�����sVN����遫3�d����R�U�Aqf�+���n��ydč�c��]��]���칶L�&��i��ǜ��ݺ�S�"���k��@HF�U���S=�PH<�ʦ�"��x�<�N�R�����5��N�k�,kY;�a˧û������k�� ��գj�iUig^���_Fr�U2���m�DoqM�\�<F��At�G�F�NfP�����]��/9m���D+�uy�����*�m�C��n����f�*�\��}�4�D��������O�ӕ�qa��ۮ���^LO#��"�S���Rb�2��.�����N��IIi�台�:�5�/�M�5�.�%��8:�����7���	U�Mb��1TeF"�znNȆ�BP�p]f�|f9&�a�iڮ�D���hb���]H6t��A,f�(t!]��V�#]t^ް���
^_':�u��م�Z��V>#]�guv`m,ߝ>����֬ӥ3[����=����aVs�f�̀0��YH���N����1��yz�C���B�f�gF���x��L���1�+bQ�k�M����u�'1]i.^7J����4͘�>����)P�(�R}���� �㺢�6����{���.S�P"E��7V����N��j�+����xf���r_�s9� ˆvƷQ�I^��0�wh�9�=%���s�4]�Da=RF�������EC5XVH��0;��Cq`�U�S�]]�����su��j��Wo��L�[�u�n&L�S��C�D�V�2�%��`I��^٭o�.��G�-�p�zc�"W�Ȫl�;˷���=�խ�#�+rEv��c�ȝ|9��y"g�e�1��+Zu2�h1����H�m�\k_����[|��I|�oq�6�-���ܩ��J��Sޫdֹ�I"ٸ���K$8�IV�E�gNeV M�Z��f�&-ѩ�-�=���3�XO.�q�f���߿�		����$�^?ky�����k�*�YB��uv�c�\�X�jz�u��22q��:Z�nn���oc���Q�)V����y8�\3vD��G��&�T��2;�����)���.��컳S懏�$�*�ߒ�4��G\=�[���wSM�mV`'"�K���z���.��l�������B̖Vvԡ8�:��n1n��q�Iu�e��xMǩف�w�a�sU1i��u�0�^<}��M�HiV��,�g����Vރ���Z��Mvz��6�c�7o_|�X{�;���5�ԫ0b/+y�2��p�@��XK�$#t��v�����p�8Q�7w�8d밸t1c.���93���҉�Y5ؚ��C�[j�=��eޥx�h�KCf���Y��#J �m��^���G%�|ɬͼ��}�'Aԋ�L�P'RVEr�#�.����E�ݐ6]�������N��vp@i�`�wЮ^��K���R$�B7��1`����D�M-��դ�Tu�w��y}�0��Rmԓ�j�kz+�1%��X.���rW�����I���]��g�;��:�5"��w�;�^RAy�%ڒ����B�sk�򸜏[`��O���
 `�Ŭu����t���DY��-!J�� X�N�j�z��G�b��M�='�Z�S���-)j=��De�	mWV��&>�(h/� [[u7���3��8���awW	*ظ:Ú7oi]eyVh��.�b���L#�6N�M��6���x�+���6�(�H,��ʳf�fwj:-��!�v�_K�b�ƆФ�B���� �y��Qj�n1p��wL�����|���f�Y[t������W�7�u��Գ��q%VӷWQ��w@&ec�Sd��);f�DZ|)�p�n�'���|J�<��s�Sc:�tx���`r����`����.y�f�SYb��*4���T��v��<�E��!�܅�� ��4�v��h�#�>)d��ZЫ�e����r>tn����q���z����?A*kSn]��3���b_�KW�NIJ�f��bY������.�u��}lje���gh�>�R3GF���̫�lXS\�me���p����<k$�Ӱ^0�ݟ+����l�H�����Po��R�C��0v�5f�n��+��̽��*�
�ZVJ%���=�1s��&���B�;fnI� `�>wA��9���t\*ڹ_7/�:��Hn�y�ձM����ֹ���v�T�ά��Pi\^��lN�PZI���/H��]����p٭�|�J�'��Oz	hWSsr��\T�X��u趔v�0���<��}w�ݬ����J�j�V�Ҋ����虭w���)'����8[�1p�������򯕻�6�񗕴�9��V��`�t�wۡ5n
@�va|Ƨɜ;�k����6�$�-ފ�4Y=)AID٫|�zkkv������R>ͣ3����*��Ŕ�2˦��fJb�|��(B�Yu�l�:h
�npc*F�w���^�a�m��lY�Q�=���dg�է�P<Ғ���iRuÑ�+]*��U�*�Ee��tDR�r��wu�W�e���ێ]���/�.e�S�^	��T�un��]&l}���-� B�h"�íb�Suj�k[��m-��zP5Zv���
��o��eI��m?��ۺ(ݠT��_T�(v�@��ՏG�w�R�I}�]�o]�.�b;H��b�&QG�a�gR��!���MЭ���\g��o(��pګZ�������f�t���z��e�pZU$|	hCt��5x�� )N8�^�����Ukq����B��ui>�������Eb�E����kDI���3G�j+7S7�7��'c�4�7�9���w2�.���uMRCsht
�u5��-Z�ԭ�����d��!��oQ�vV��`3S���o6]A�uiJ\�l�Ш��ꛙ.�;�/C�+�ad0ń��Q���]�%�
'�����]YG>Dۧ���,�(�û���g7�W'7VHRj�zZ�C"�NJx��ո��2��IFL�����m��7V����)�f#�<�}��=úӦ�,RTz�}8�D����ݪnf�,��4t�E�]m֧op�y���e��1CB��仑Mz�`�p3�GW�i��aR���G�[h�4rR�;?%l�v��S��WB�N
��{b�A}��ܡ؛b�<��NM����W�גݘL�=�_Az�k��L+(X��`0��I�=]/1�v$(3N��:�;��ʄ�>��G�N�e��UՒI�#�Wc�&�p�QR|�aGfc�m_J5���*B^��dNYr��V���ך�����!���#���i�����EcBw��r6����_6�t��tf�I�mM��R�{��q=���a�[t�����[�Lh��>�A;ל{yC�Bl�w�O�֮�[镱�ԛ���D��b�k+L���[M��6��զ1%�g�&\���}:8̑��%f��t����+X��lwn��/}OU�!�% �d��gtdv,p���2l�Wܻ7&4���Vj*u�k.�+Z���L�T���\��q*`"���TjŜ�RA�&k�'(Ŕy1{zy�p�Ϝ�?e�[d^õ����ǝ�I��M�h�K,�8oqF�w{h7t(�-o�������1�ƪ���X�ӕ�=��_r�hbz�RB��w��V��WC��t0�.�r�S]���)�|UfX�S"v��zL�(r���f��n^͠�ޭ1�:�c^Ǻ����<�s��JN�q�K/��D�v�Jl�Xu�[������&5�M��$ⶰ���m��ȸ H3S[G��FpTU��W���r�\Ks��A��N����ά9�)25�m��.���˻i%� �,�*.�K�����sh��M�0jT2��x�����n݆p�G5I��v�|2�1g1���1�R_>[Ŏj�u%���JY��cA[W
5�g�@����D@3����o��R�Y����v�gD��|Ν����m#B���y�"z����Y|/m�,���S�v+��R�w�Y�]EM�tifb|�Y�����ݘ%�7B�t2��B��\�2��ӕb��ۙ�0�$�ۡ��KH�v,�7�HZE�=�@oD��!��,��S��hǵmi.�P�aRI�c���w�÷M����QQ�i�gcS)�������g:�6�:�VB�������.KEf};�1��/�\ν��'N�s�r�ș��{�kf�⭮�Yؾ����64L�e��$�i��C\���<3�N�M.�u�Z����z�Z���V� ����K6u:�+<6\�x�}�\�E��X{j�8��AGN���ؠO������g�ˇ�v��X �Ad��ߺjìj��AJ���&X:9a0/nlB��q�{vŒ8�7���eA�Ő���	R�ɭͺ�xsM�5���e�ŕH�ü쎨�֓��έl_�zU�̕��6l��qݧV��k�

ɽ�a���SY۷*6U\��"��W^l@C�s�:IF�+,W�/��-�`u%*�JUÝ�����}���Ʈ�܂TS����7ٯ�a2\m=PkM��y�lf�e��ofWX`���0Kz����Vb�&�d��{pE�W9rꪜ�9v@�#	Foi������@><�,ͶN&����V�&[�sV��py|�<�xb6z� ��N���@����X(�<	���;lO�,�K�9�kLđ*U�K/��qv���t�Q�����.i�05] ��C���cƝ]j��[
�V.[Z�=�6�HTs�Y;B�#v��t��Bdsc��y)����X-�n]Ct��C�3�L5,4�r5�h3n)���$�w\�/ɮ[n���Է�vh�v�}5��v9��� b�Y$��W(�������]��9���x��p�]\��Q���:ƪ��I�L���
'/8k�y�W3fI�0�-��-$�5���,u�A׶�Y`d뾾"�K|Kv����fc0��W[�JY�p�cO���٪���wpҖA��j�kT�V}��t�:$���0�R�����g3�6��f>��A���P��'�X�y�Ҕ2w���q!���:�q�]�w+bIV�D�oj�5���]Cji�d5d�p �k5ݸ��W���p�
d�`@v1Kv(�n#;��*Q���7�}Dr���)�� ��[WK� �P=#Y4hg&��Ry���ƺfWX�oO\��=��I)�;�����{i�F���m�]�hl,�R�FO���m��2&9,*^i��V�f�a�vnY���ut�m8T��%f�O��#/��Ij�?�|]M��k)U�������9�luʫf����h9[:��(�us�V��W+Ä�t�㖣�ge]�GN���k��,���Ñ�s%s)��w�
��ήUd�^&�J��EL�p��;�3:�=�L�ж�G�YW���e�7.o(_gi���3{�u���#�(b��q����z�gB�"
=�	0�5���J��0�^`����UgV�dׂ�QÎ�y+��F���B����p�I�2��k�[+���7wUx�έ!��C�K/n*7�D��F�{�S���"�!q:^5��5d�ltM�{wY�Tw-r��ÙV�&)K��FO�:ﬃy�;$��yG��U.��I�GqթE游e������F����[iVf卫�\-�u`����4��f�d꾲�b΅�t�Kmҫ��G9=�Qnjb�;AV�Gv�)X�u�S������,�c�s���r��"�� ���`ѧo-�K:+kR��,։���=`�!޳�YM_h�X篹�p8 ���ݳW�������IVw*u$��gw]1ɑ1�D��y�8� ��/��*o�)f�Y�X
�JM �M���uNVag�(Zk�	�%`.�컚�ύh�PD��2�/{Հ��rK�hI�v��k�ÝҸf��w�	���[ө�j��9΃�;�e���YFd����.ϭ�to�))1��yA.ؔ�<6��p�GL�FJ� �,5��+O]&��B�++HP��I[�e�q[��o`��K�Օ9�L��r��Ú�҆�x5t9�(UZ�P��	yEf�mf���52T}���m��8�΍T���n���:l\ ���wP���I�����m:�%��Zp������R���G��v}+);7��o]�l`�ޣ/�>(�����$���\��I�heu�Yb5�:�Z/��u��z��nwp�h��3�7����TE�ܜD9��ܮH`��R�U�:�l.eCHXrGצ��u8\t�jw[W{��K�H7M����s#[�Bm�ۻN��BU����˓���,�'H�b,�X�6/X�A����nL"��u�W`�K��z���(�]�D��k{U_(�(��"���2�6k�=l���T��,F��m<>nYۿ���&*w8]&�.i0�C������6y�,�qw([�I���M��Zc�ȱKN��f�щZr0Q��Z����%��0nZ�)��״�osC؇&�`.��v�p{³V_OF.>��%̑-�.��d����+:������,���(��C���*hȪ!�5S{Z�������S+\dT������pp��9�ņgu��+s��Rq[jQbZTf�M+��A�\���%�[�kuV��B��`o�Ifu�L�g�����f늝Kkd�De���
�#ЗY�8m�7!���[M�ֺr�|� ��ӷy/Q�)K�SH�%�L���F��b��Ks�Yڴ�u�ڗ���T�]]����\Jfb�hU�P��bf<6nK�u���������{�pm��ж���}�e���]V�u�$��ZQ�i7J�qT�:u��*��*��j��I(H��[WM8_`SZ��R�d�t�9�=s��)�Ԅ���穛�\�?d�i�j�:���*��e!1V�Fn�;-�4f�,�ާ�e��L�t5�����*��ڻ�m|��0Y4�(@�v6���ʚPÁ�a�٨�c۽�/	���[ioW��dv��x��ky�s�w ���l�ҳqQ�q�R���z��kV�3YK�S�xԮ:IS#yr�Lã5�xx'�v4�^��5��f����.���ǆsK��a�SrT��0%7�������s9��Z+�Z;Y�T�o���v����m�[�uw42Ҭx��
�*T�'_:��]H���}�0iU�ǧ�xD8\A�Ǧ��OJ�q�e�;Wt��B����$�]n�F�B�YAjҹ��CGS�hF�jغ]t:�TЯ
���;��<�[�����f�X�'yv�M]���ca��,X�$�o5�z�c$u �s*V��@<�����Q��k2V������hېÒnP�M����6a�b���z�d�s�ZS����Qf�׸�޳����s��V���G�q���N�nCo�&�6,7}C��k�, �sF�=��zi8w.����ph[��3op;�í:(��b�'N�F}�M�7j㉊��R��jtv*��d,���g��X�鲧s7�Қ'u9�"�6��N�G2��׻:�aq�(Lv�G ��ܔv�6��.(�ʗB���˷8�X*t��4%�m���זp޽���.b�E�J82gW+�КƧ��L�6�m�I���+~�Y�DD�������.='o	����G��Ժ���|���+�݁���Vi�,uԐwV��gq���ft񉺔�!�
�24���<�|*�
��+��6�yZ��U���[�����ʷz��9�Q�jܳ�D��XO� /������Ɂ��Y�64�mڝ&�w^]�{W�T�泆������GG �.�^��5���KK���n�����6���V����/;*�r>!�ƅ" ����(�}b�-3���݌pG2l��ݼ��Hv�h]i�Ȕ4�*�ͷ7S��t��}�3J0�Y[�:�4���}�s�s��F圵Ks
C-8K���J��G�!J�����P|c�8g%����,�u�Z1AP�ͻ��OWH�����b�P�W�z��"`��K.K�C�h¶���^k8h�:2�kܧ�E�IǼ`]J�@�Ȣ��ݶ���*����U;�Ip�͝�ͧyY{\�6����V��}�WlYfK��͵t�8&=��o=�x
6�6ls��}���_5�y�j�+�VY	Ót�f�+�JT.����!2f��XzLr)3+	�6��ԕ�frT���}��2ҧ�7NHy:j���nc
]Oa��:��{�S� ���h�|��7t� �kfڰx�-�J\���R�!��8��ef�(�^��Я�n�u���t{ݭZa��1v����Зf,@IMŚ�q�z���'�j�ׁ�턴�W)��킛�L�s��{]i�Q�7z�##J�%���h�-�S^�
�%��,օ.%�UiK*�mk[(*�T�0Dm�5EKh,kJV�m�0��T(�J#,��J��BҌ�T��Z�VT�TDKj��bѢ�-�*�ڕ��bԪ�j*ъ6ب��JĲ�E-�h��iFU���*VV#YmjXZե
��j�R��jUAR�R�Ĩ���
-�B��-�lU�[kZ�"$UYZ�U-�UKKX+k"#[Z����VQ�*DZ�����[(Ɩ��
�E������h)UEiU�"�@b-J���R�UQ�"l�KB�m�A�T��-�l�ZR��5m��*�l��aKV*�J��R��-�KZ�mZʪ��j4*Ū4�)l-,�,Dj"#e�m�R�e��jU��Fԭ���V��6�Pb"��ڢ�[F�*�-���֌[V�X6ђ�Pb�jҌE�����"�mD��U�JԶ�j-�6"��D[hň�ڡUJE6�YZ�Q�R���ت�AJ�����~�������[�2]�mt��pn�q)��Ah�A�D�8`�^�#]�|e�[��!y���1ˣ�&T$��P�Q��X�B��	�e+���w��ϡ�1� �ؕpbݧ;��_�$Zif�?@���*�Һ���#�Y�q�����|ː�Q��LZ���l��շ�eVM�Akګ�9�:E�̭QϪ����j�%B1�������z���މ��Nyj�ظPr/TۚݺxqV۝[/(�I�
��:�Wr�ǂ��h�x7SGTm� �9:��'��ä�'��t���x8�x\S��n��C^z3�{s~�SwlZ���֐�)�2$��e�5���h�7����|�n{�xmXu�2�'7���1�fi<�R��C^��/=Y�3��v}�h</�����V�KYp�^�ĩ)�̶���q>��Cz���Z�1���Βé��y$�[�ό�56��}
?y��6�x
����p����/R7�͍� eq#�H���m�� ���e�
,%�jL���
���5���x�8��v����nm�;X����o���1��c��u�j��Fnm�mk��&B��t���Č,	.p��T��L�qܨ�Er6��с�c�w�vec�aէ1m�6�����յ�����|��{<}��(�Q�ݜ�̭)K�i��Nt��*{X��y�i5mi۝%#�>*��}xbw,�����s⧧v�||u�t��<�9������s�M/:Z��N�LL���Uܥ��/s����hH@��&ъ�jN�vy�XX�cY���؜�S	=d�"��I�{$t��A���U�s`�#yk�z�!c	X.�~�����c;����s��5,%3��v#�Ld�,���{��8�QYlZ)Vd�O�`�{61�Bp�k���6��p�\���m����u�[��#��d�dKJ�eܽÍމ����HCW:��-Z#��I'NYe/.��dݏGsy��r�gWbZ���SաJ8zUG���8�E�.��Bh��@Ⱦs^�س�;y�)N'��T��!��4B�,��c�÷�@=<�x��p�\t,Y�s��%up�X�.��VX�c�����I�b�V��,!��3]�=M�+�P�mz���^w� ֠ja�'w;����,Ki�7(7ݫ�����8��۽�ܝ7J����Pz�P�d���3���ң764�h`�m���踅ϊ����YI]��:6�ٿu<��Ӻ�z�hf-�f�wg/����ڼ���VKP
#�o��&���oW�Vn4)���-�u*/k��/m:今B�������k<�6ͭ����F����L9�s7��i��1%8nI��j��m��Xg �ÿ=V����|��g:j�b�6��Ȩ��X�l���4�&0Q�=L�i_��(%����ݼv��Ӽj幨���7��^�M#�s�8�h�Q��	e^K#���-/bܷĈ�'���m%���+�o����p;jC`ؤ-�|��;i�
F^V��z�[.GU�E�0l6��N�G��c:K�c��nh��R)�����]3�!����g�ڙ����n��I�^�@�B�uh����o�;��*s�ow���|��{���Վ�`*t}�rWY�����m����u͠`r�[�;t��,�!����`���#�NS�LΤ���ݹ�nt���
�Y!06Fe̥��p��u�U�5*<�X�@�����`p��6g��^i��h��J9&U����u�*0k7�:�TH�)A��d�oo���QXZG l�t' +^0a�g���Q�jƦ�%7[�\˛�y�ͩ�j�Ӄ��c���I�1�gfˣZ@�m��x������#���(�*�=u��
-J4�#/4T)7��ʫ*�+��C�$Ӓ%ǈ�+f*�ǟ%��$�����E���n�`�3U��nB]�,���τ�u=�P|�.���s���e#,�yR/N[�����
<sl%�Y�SiWF)p�T1m������"� X�^�%�`"�X��nhm	nS9�ϳ/l�-�{sM��vbsY��.
�ھ��֫VC��C��VӷZϰ�7FX��������Q���x:7�߻����[K�1f��짹L2s�9^�;gu��۽�\|�bE%����n�b�c��8�8\�;��c�|�{/�� �����QN-s��>
�j�_mr�uG��|�xO[T�U��7])���{�<��n��}}qU�ck2��
���Z�L�S��T��& GW=�ڇ�[�Y���bFb9\��(����wN���Fm^���^r7�a d��Bt�a:ˁ�Ά�v��%�Τ^� �A��{o�؁�*����\��uJ��i�ܺ2�O�E,��z�s�q��!��4��̛�Ej[�F��5j<����ƚ.Vs7Ĳb-M��ŵE��	ڷ�eF�F���Tbj���U|o©��"I{==�t�ċ�֤2[N�T�r�t
rX�,b����ݨ�:�ġ=D�l>�{g�ma��h�{�%���/��؞R���XrJ�rڠ���9��)����9��3�ќ���k��Cڀ��԰�ຸWꠣ�/���߱�hϯL��?�79�=J���6T��t��4�EiT&
:��PCƕw�E <{��x<�1gV��h5'}.,�s�i�^dک4ֵ�1�{p&���H�J����0e�Ԉ�T/@�ve��S��!�֚�i,��۠�Ӆt�ln�*υWP�2���i9��S�e�Ė%r�Ư�)�Kְ�Ҫ`_Nr�q�By�\��u�d����GL9q�P�X���J�ҚDJތb����V#y���8.f��wU,'LG@�qY5Խ���\p�4�O��Y�ac�/"���Q�T����9���45nw	�<j><��9����p���tsi#5�ИΒ�aae�h�C�c|�r���,�-Ct�3]���ɵ���T�iW��x9 	Mmb�S�,q��eS��\&2��rJ�z�`�Eu��juv�r�}u.�y㑞.����E���3��I����q�Z�<�i��ʨ2+P������b��6���u�Ӯ�-Oe��v��0W���d�~�0����|��u�~�t����|�ǂ���u9�npP���W�ݭ�>������IևU�U�r����N׍e�&)~!FT��,۪�`�:���l���U
[�Bg�з/]8�<[с3c��26NmZ�]�A�T�:�A��K{;�ȋ�d1R�^�bC��U[��߱�	�#δ���R��u�*WkgoZ�|J(�I�(m(�UhN
T�a��c�c��b���,c��ǖ �F����K��Z��a��ͤv���,uz��AI�h����v&,���{�땲�"���o�CGSwDM��,���c�g6!� t�0dԡ
.�/K��L�Z��hb�$X����a\�l�$�l��i�V����0o���VyxDj
�5����T�=-y|��?#�.���j;�᫷3�40����h��Zz�����FI&uūI�̓����jm-_s���NF�`3# R5�h�֣�m�w���bl���6�N����f�zW#m�p|U]�+�++�p�(�wH�������$���"���2qC��)1jK��$�#�ѝS�Eöl½�<��V��;(9��:�B�/�<;ݩ߮�wl+�h��L��N�`�V�b5Y�ҁ�N�3N�g���S���HBTJI��5SV��ruW3N�p�It@�q�2�c��\_���`��ʥ�)�W&�܇0�LJ���,���Iq�3��,�UՏCMU�J�U�O�r>�?)�D>3���^�+�AU�urV��ǳ��Tc<<��o:h���W��/ƺU%�=������<}=09�Yt�ξh�"/��ˮ��U튰���gؼ.�kʛ����7g�(AW';����%��L�}ŠjU�a��a΂͆0yӉ��]���LՀk&hh��}�U���[����0��su<�r`nu�S&1����O�r-m\#՗�O~����α��/-U���1�M1_�lMv+᳾j�ʿ[5�؇��E�0Ǜ�{�|�gH�J�C���w'�m? kL����쵟*�9�4��]tZ���
4��5nRt�ܰ�ʄ�>��"����7��n�Їz/Q�ְy%b�P�v떵̍��csot�����,���9��\*����(�L�-��>��+w�k�&4�)����ŝ���F#�f���R�n�Cj��T���%�a׹:�7Ya����8jҍ�z���'L�-�t
v06��EBN�W^�|;��W��أ��;�<#�7{���J7���J�`:kT�Q2�J㤪��R���WP����"en��sބhDLy�������W��@Q��y޳�<ݭ��0ciVxL�M ExԄ!���#y�0�s��yro_s�I��[.c�L�/�s���� �=R�n�1<�FJi�]vwj3]�$�$R��q6s¤lv:P2�*�c�b��tʍf�����)�U8�p����e!Ud�R��	p��u	p���fjZ���2BS���8)�@:-T��b�jH��,��fQ�\���|]"3˥4k�V{W��z�76_���;�,C$���p����䯆ƺ;�@͈��Ĉ^:HW@���%��$�.��f{<��7���KJW.�(�a���'Bv�&P����	��TtK�cb��(^6b���ء�6�4�Oc��E�)���x8ڍs�
�/ͬ�������:�׈����[���˗1��KI���]��Vo-t���WL^�01z�Ƶ�=����c1�$s.e-�O�<2X�Næ�eʶ��ppm�3;�	XwT�SaV�z��ą���l�����4E[aI4u��-��C6���l�ws���Ԣ0FI�"0�RD�$g?Uvg����
H{,�p1�[9�Z�5X!��y���˫�sW��GRB�1���mnJۭ�~�X:3{x�HCg��;fF�5�:ERؐ��g:j�-���̚�u
_`����t�X}�病���uO�%`;;n1��b��}����w]�����P�0��%myU��╯	�o�9�K�E���4�I�b��83w�n4�Q�f����x���LҜӁD��9ٌ��(�|��c�3�a�9�Mv�����qFJ��bڭ �{ҧdvI�ꓡQ��hv�C��:x��|g�n��l�ܡp��uY��Ʊˀ`S���X���ڍs���X"�$j�ڍ��L�:s���'�1cʮ��#U�g�3nt�oy_��
�J��9��3����L*t|r�7����P_�V�WEZT��|^8��~��ϯL�Xn\�d�ds=�+���
���4���}�K}
B���H�{�t�>C�G	ګ�t�~�$_u���S.�R�޹޺5��Pa[��1J�,U�N���W7X3.�U+1^
h����0��3G:�A�{�r�TyVT�U.�72�V>�V�V�VmI.V�љ��[�lʖ�k;���[S�>�a�`�v��� �N��^�ϊ���]�)uNrv5ȗ&��鿆+p�3���/8�B�������E1�:���t7U��}�/
(�Ht4b�3%�Qe
p��͂�,�����NIN+%��i�������QK��=Ň0�9�u�RQN0�~��p�K��D͂��O�	����!<����%Ҹ����C{f���*�b7����8e�ܾ��]M�:b0T
��y�+Y��s��n��[J~��ܼ�g!��d����hs���u����Gf=�#8���J7ϭK*�ն}��L+O��c4�Ү
�������Nv%����c�G��kt��(��<�߼`�_]W�\�SA�`ן�¾��+(�j���Z6)��V<$����L��G
���n��7�d��Ó�W�v[4�h���^{k&Hr;������=+]bNf��fo�>56J��ʅ�z8���g�6:hf��g���Y��:
��wY���I51h:unD���[��!�npuU�[�����NE�Ӄ�|R���+a�ȁ�Xm��[����#se ;���c//�F�gm�kyLʈ7"��]�E��d4��T0-��
��(�m;��{s�J�A}0 
;}����J%�ƵA����h�{��w]��
����$�j��_
t�}�Z�ܔ�\�Cz��G-�+����̼\�X�n�J���EAN���N�(�{��6��V��.M�D��m���:V:�!�t�C�lj��qw{X[�B���aL�.F����[���X��u�d�r
g�(��ti g�ʱ`oP͜F�ֺ���p�Ծ����5�ˡPdtCZ��.�63�g7�������Z�z���U�A�%n�eD�.1�y<MwW:"�kj!��i��̨>�ya+w�P�ڴAW��C��Z��^5�AдU�s.���mn�
����|r]]��v2���Ǒ�WU�nSo�n�
��jȒv��7�Qk�+����15 �	��c���O0���w�m��&]�h�õ)\��5��E�4�n�M��$��Wv�+�KwiM�Nm��xc����]���'�*��p	��?���0L¥]���di�gv4U�e
ɩ�DPj��6��'���f��^Jq���W�z�1=Q��=���
��N�v��F�]s�L@�k�k �p'(��5GwS��;�[�pb�7�>1촏l�������3hNǔ�V��	��d��%���չ��z��P��#ۄc�L`p�_��a��B]��A��V���I6~";@n5��d��h�q>�0>�Y�&`k�}"��P�.e�i����Y�X֋����܎݊#'JIS�ܭ��,09
J�0��@��B�T���J�8
|kj���/i���E�,�Ŭ�%��N�����i�*�\�_	��龍�®K�0�Y�y�S!�t((xA��䷗7[r&:ޣ�ث���4��&Z!����;��ř+Y���|��؞���q-�Y����'���8*���a��}E�3
�Ӫ\=���LKE��"�8R��n�f��Q�aRN\��n�EN�Pս��iUd�
�:O7��kⵜ���lvhkߚ閎a���M]m�W�}��1�V���I[*fkV�
�ñ��E��¸eq�i�� ��m��6S�ȳi���˰dg��U���h��T싎2wN}�YDN	�W]Ŏ՚����L�z��̩�Y��Yok,0�i"^�[Z:��8�Ål��,i-ډ�����5���u.P��l�9w�K�0��玫��F��^�[��5r�k��7��ԹN0˙��c��,�&c�%�D-�ɐ^�%�C���7{(^�r���6��,�|^���ð3tw(X��F��c��,r�Wj�+�P���r�d�D9ۼ�E�Whz��ޕ�X�z��WH���^^.�{&7��Nu����s�C���Oe�}u
���((0EDF5���Q���1���1���YjU*�El�D�Yb֋m`��1b�4E+b�h�Tm��J�m
���me-�Ukm*�[Tj)U�()Z����Kj,��Tm�m�����QU2�����rU�U�h�*�#YT+TX�m���+d[E��֊+KU33"�j*����(֊��10��Vҭ��6�m��i����(�+��X���L�QE-���q�!��S-��iQUX�U�e�b
[
�j"
��-�Z���ԥ�J�Zeı�T@YmQEZ�E�j�UQ�"+2�Q���V*���e(V,`�,[h�2�����T`����Uih������DV�pLf2�"���Em�5�EkT���U�DU\��ʋUQJ�$Z�Ec+ET��1�5����`#�)T`<aX�>���r�mT�O9��f����%�puU�\Xy�4c�i����7�0�>�ԏb\�z?xmC����')ҁxh(���8q.R�,c��8��[׊J}O��L�gb���p���^�:����WR�����LY�	��޹W�W5[�N<���<��1��[F,&����H階���}8�$�����
���+_Spd�����kZ�(d[�~&k�
L��]�I�q�#�=ꘄ�]�2�R��@��7c�i�>��f˝F�ȸ�lمv���;�+&��%yBp!*+�B�̚��8����=o�B!I��M�60J�fK��S���K�,�>���F�P*N:�,���x�;�i�������˻�3@fҌ�܂9A���e����,���!�x�v�35��,�[j)q�,��7D���jFB������=���C�K���֧|��k�[P�SO1�6�v	��轅��Z"o�غ�	�P�Z��M�������b|ch�X�d{�����Y:��g[�DM����	׶*��٬�qu6C�v���-�x\�����o�%�e��3;����͢xcU�췻q�����E�h�;LU�&RY�3\kL����ҽ:
�|�����̷�c�E�통
��R��t�����"7Nj�i������7qoA��@n�7���]MEڵ�$�e��v�U_�M��$#{#�nq���A�}A����=���{fk�d�h�`h��<)��k�PtV��[j2�y⺕[��t��-Y�W*�R��ٽ;L�*}q����h�x�=��jI�91R���xk|.z.�[���8;�؇��E�y�=m��2�����˵�I�}�$x]Ȧ��ҨS겸�V����>��8mZ_p���}�^������#D79��I�^��c|�#4�W��u�`��6H�B]	}E��>�]x��{�����H�Vpe)���<��-�p���N��f�b�3%��}v�S�z}[�4�;�$v�]6M&����1^W����ݭ�Y#E�P�V��Q���D0o4���)��zi���&��0M��3�C1J:S �]��6�*Vĸ�W��V�M�]���2^�_&R��T�L�Q7��H�Gc�-�2�݃:�sq��,��ȝ���k�s��ED�����q"���P���q�q�w�lY�6�Q�|�ǅ���@et/��p�g<ժ��G��8/�vי�-%���s�]����Tyds';����a����8�ˀ�>j�,��r������\�8,۠���r�;寙�U�ƿ�S����+]cx����#A���WE|���N�_/���U�K�l��ʁ'��1�^	��o�Dg�"Jv�|�g�xJ�a;lD�1�f��<+����OS ��#�x!���Ĉ���5�+�W�k�UP�(d��fǞC�D��;��ʑ��&K��'�&-I�'n3=T�d<�:"�uu6A�VR�/�_�
���A�C:�dSۨ���2L����c�Q�T8XmeE��� L\s��.)�{Ѕ;��������S��w���\�����߶�V��ۘE�`����};���U
���̓�x�a@lN@Q&4V������V63m߸�hC�z�����H�g�q�8��彳ܻ�H������P�_xXUt}�ѫ�v�~ ӈc��+�"./�D�W�NV�t�jS�!a��<� ����6d�"����V�'����Q/
���c$/gu��Ť�s��^C����㵎3θ�A��Lҝ��б>� �
*Է8K��.����d�)iQ�B�N�@��-�P���`c�n0:�vTo�꒤đ`��R���d7�&Lv]�m������@�	�tR�R|�m��b�k��Ve-��9���!wk�T�K<�/���Ŭc{e��)���*ɗ�Cq���O���,^�Y�(�8(�7/r������k�=Ԩ�]3�W3s��
'{-r���;
�U���.2��v,ϼ�Y<���|FA�_�D@��:�S�k��"ܬ�,b�x,�F���Ī����uV��x��`������ãUE��Y�m�{��\�
�J����{U��I]A�zN�)ZB������W�|jI�()9뫇b�(���ƅ�o��/��.�%�w�Ez�{�������a��N��]��[D��e�>C�G��H�횫cQo��]$,�~�M��C�&{C2+$v*q"��<�b��R#��p�T{�Bt��'���u�p͇�(�3��
1m8Qv)��:��	��l���^B�v�.T��of�=�C�C�G5|S̞��$R���xM�����|��wy0��!��wڎ�%�����+̌04����0��t��>������}����N���i�ј����9�ue��|�=
�X��-Eň&�{묍ݥ3^��^9��nOoe\��]��ݴ��1P�7��3=�aSW̬cƛ��\*ŏ{�©9ؕV_���;V[���<h��!�ܶn+�94�5|��{W�^>FW\�$�tP˯j`g����ݭݏ�ևx/e���GH���d�!7&(h�]��~����]��y�1ϟY�M�Jz3n�v���e�A�y�b3�8�9��4�p93��V�L�W.ӽDn�u_����N7��ŨQy�0�۾��f	{\ҟ*d�Q��U����lSYCa��yF��}���+�� ߊ�@�3^A͝��I��} �����^��4C��8U��>�x�I���8��H�R:�뛊&��{j��ʅ�z����:�J�k�.�����Z�j��lZ�K�<�P�ʋ4.��H�Raa�p��Cs����Н�;	Ȱ�N�{sErtZ��
�i�������Ȣ�w�l5^\�����¦��FvOOg�b���,c�0k��o$�c�)�Vǋ�S�*�{�c��!'n�1Y����L��ح{8���g2�����E�髞r�"���X8�́��Ȯ`Ւ���$m�k�S�toֆY�1xn��笎ŵ�����w�gt�d�3��ڬӌ�#��c�P�s�*�F���E>�9����f�3=>w�˝F�ȸ�lمz1獄�d�;5�]	���*�A/�wo_^&���L�OA�u}7\�`.��h�3�.�����S���7w�:p���powjȫ�o��]묎�yֵ�8�{�&(V�t�8b��%��|��ẕL�9)�x�NFh�M������sw�^���5f��4�<
Uuro�X+x=E8!���C��3��X0p��(�	�
ˤ�{�5��M�͗��}���^��/m>D�(ĩ�
2=�k�1�B�`���Wr� �vL�Ai�0�i%�^qsh�ۣ\��~I�!�Em[��Uc�����<�N�?+�|,g��ִ=���l���g/�9�W>��dH���P��c�;Y�n|l�>ji.�;�A�Qd�)MP��%�U	ϲ��ɬ��qu6t.��t
��Cs���̅27�N"��*��oz�0F��#=�W	�}A���ö�S��?���tx?1qJwi�\fv�VX����H�X�#�S<*Lo�F�h�{o�}��g�4���n�VqK�.��]�V��ĴW���~5L]mu�=c-��!��V�<�R-�0ǲxDo�F-}�cY��b�9:C�5,�qX+�CO�蠨��]5�����ľ�fo�[�%��NCѾKЙ�ŵ�uS�{0U����v/�QU�a�����v)ـ�M,P��iX�	���&��L](��5��s�5ni�RB�&j1�(P��;<.�H��#e☜�/|�ʉ �ט}��3֗s�%㋚��$8D����;´����ߎ�p����$Qd�cG�oL��tG�neCo�↔��\�m�$3 �j�I����jw3V�W^f�Oh��܌�����#L����_.�Ǝ�,���U:fۦ��@Q��+�Y�O����L���Y3�4��ƭ�J��{�0o�$��6.��y��߲�8v���Z�&%BC���~��F6�\�n7*lt���UZӭ.؝��N��2d����jF�c�=n�`O��u�*%��|9�9<����M"�������B\j�&$C��«�B\
���c@'^5=쐔�F+�KF��<]�쌍�	���1��	D|z��h���@��p�����$�1�<:^)���&Գ�N6�C�]쐢�S9�n�D�N$G �M+�P��՗b�b����+n��|�HFDť]�(�U0��	یʤ#!��@DP3S< ��jE��u���d�~�\���"\�	�ʅ|0��7�mƹ�p*��TXN��b���u�lV�1���/^�;���- ����6/�jښ������a@�����4p1k�nc.n,�(P&��8���$�+*�8����1�(`�2�7���)X����W��7+����"��s��[�N�3x]]�X�+O��ؑNb����gr��^���C��`WE���O�t�����r�� -u���({���g}n=��p���f�t��E��BpӒq��g�=aqŊPy�NN�3�p�����tA�2c��~� ���-#�!�U�+�v,=u
���,+��HՇ3�����i�1��N\�]��#�%�vS�*�5�l_N$l� �<�=3���H���eϩMVӌ[�T}v��G&�Qp�f���RaL������4�`�'�:7zf��&f�z�"B�s��i�Uڱ㖹Z���t�,���#��x:l[T����҆P;#F���17�z�'$ڡ�[Ǻo�E
��UFϪg���}4jH�X���!¾b�$�(K��F���#/\��W�R���sIm�0}�,}԰`t��p��UE�����xasO��mS�vJt�bր|��D��ɑ�'c�
��S��Q�ba'���v*��W����?�⌗�"[?a��ӕ�N��`۬���,����{bb�4ri��#��&C��]��j2%��۹7�Ʈ8��GR�]�!�����w@н�x�@� �N���r�b��U
�x���<�"bA��X��q��I���A�b\wL�����	��p!",�A�X	�'��fr��t���K�ꥎlUK(��x�W2�J�%��I�=DX{�7k�wp�I^.x��v��S�,*�Z{9��ǹ�H��Db�s��ӽkq�ّ����ܬK�r\���1I�֕��Ƴ��۩�C��vjvkQCrUPg���<4��-�<Z�}U{�U24�?Jy��7YȊxfp^o�>l�t>�]�x�h�CÛ��ˮ���Ռ/|~��ii|V8=t��S�t��>��u�%��H��Y�[i�-G3X��<�A��0oU%����p�k�_ԋ�<�!/ӥL��j�����W]]$�)`�_EE�����7Y�J��8��7����bǼ��.�P^eb&�8~��b���rSٝ}��no@	*��lf�xf���5��}��9׳&���<��/�,�0��߬g]�'�k�9���-	�0̅�ϫ76�Sљ����^��n���DG"��2��ʁ�~�˛(����"j��0�����6hlt3C�z����7��f(�O�[�/�(�
���uZ��!U�[��0�%9�V�jw�n�r7�{����R��Q���`�a7f)h��MTFEpt�zi	�t�X�A@�[���S��ނ�Y/���IfTh������91�T�
7�N�|�����]WS��&�Q���A���	^�ɯt�|�w�h�;��
�6Օl�����P }�>�q:*弉X:��t	�a�kjQV'��G�S�|�F���>�me�=�e#�g ��k��3�����M����|�nۇ9��u��s��k|;�4�~�����Ը�r_#6O�V)Z%�E��b�-������Y3*�������yY���z��/H�rV�����Q�|-_���BBZ��z��Sr��A�>���3���$\eF�6MWbI��ط7J�W�ʝֹlم{�<m;�X%�9��	8m`+��y 9jDa��J�U�Q>��==u{7IX�]��΂�@��[�)�l��Y�@��)E5�K�{b>��u9\��"0�t;�K��g�A����8��!ֽ�������#�*����ې������+ʡȚ�j.���� 9�����v���k1V�F.�.U���n�,��Ԛ��/��P�VQ�$/�JBZn�Z������"�d��n�/4�R�ʀ�_���_X��e^/�����
% �w�oP�8�mOD��g6������ӎF�nK�'N&)�_@�j��&*f�e��F�@�!��e>��Ɠ���r���9�
#E�<*9�{�i�!�W�TvXr,�\{�| +�ʧ�9K^S�%����nN��yk���٧����i��9<ՠ��E�F���*A'���MG�E��@��M�@i�He]��Z՘��4鱹L=�{�J�*�oJ�H��P���8�HFV�(���4:�F��j���:j��"��Rv����GqP�SO0q}�+U���@�#X��owM��ՙ`��F=�c�{�-�VB̷�@�e�u�`�n�8��]ʈ(�%�1NS �|�5)�Y�{��L��Z]u��<��Z5xe�J��2�o {5�Rw3�r��ڶ�.05N�Z���4^���V�:��#�������&���]+����HhR��\V��H�YaA�E�['�%��,�����j]�L�v:�x���y�-�|��˻kb3�n:;��
�3#Z��A��ê�5o�S��@�9{\n�$5r�.R(�+�_Js�Ti%������ʭ�����g2}��ꕔ��ƙ8�2�;p���Ym�N4�l�P�����}]���W�8b�HIm�ۋkd.���\h\��͌�\��S��H����i �����wkDr��3{uK��r� LTV(v�
��OnUу[�N�a��%6��hA���ج�ir��dw,uC�,|��6��u;ovEʑ��w���.�:q�H�X�d/0^��]'�E����]I�{dpC��Y�  -	.�*)� �j��;�N��a�:Z��xm��AGD�,��e=2��� TG]^�����F�R�K)i��eq7A	h�1����;�/{<�*{�{dk��>"� �g�CY��S��1���`�o*7B�3/��vY����]�2n�8u�[}��۔�Zs �����I�.��I����a׸������=��O�@�+2��u����2+����]�]9{�"���P���[]��'�Ŗy+P�}��䃵����$�{��JrWv]�)5q�9�5pl$�d|h�W{��vSƟM����b=�
�b�'�Cx�N�_��c�
3"�������`[��}f�ӎ;Jк�j�DM(4� q�|�L#jN��n�h�+�JR�{yq���@ƶR�#L�W�_�����]'ٚiu�wj��3��/�l �꒴�X�+���f�^q�|3M�}|�ό�eF�#}!�9+jX�8��C)�DĹ���ƹ<�����c��:�M!R۸���<�
��rȞi�c����Pv�4�,E{�ʍ��6�e|�/*L�9Ժ"t�͕ě���ҍٶU%,H�۠FT�!j��#��s���#�����>(�Ҙ��Nd8n������`��u���|r�p�܊��4{�z�YN�%1�>��a*�kX�"��Z�FkU�]�"�44�����(	�y������&i�P�9Uع>����5s�ȭ㗹K�߮t1cᅫ&���Wn]����C5.lޔ����2K�`��,�i�'�w�U��J)�Qq�c"�bQV�-�R��cZ����UQU�%��U�0�K"������YQ��Kmh��*G#�QƊ�E##�m+-�RV �$�TAQ��!�X�fY�1c�b#iQD�
���V#b
+*��"*�ƋV �х��
��cc2�+-F(�6�DjUb*��Q�AU���.`��L��KJ�%m���[j
5��"Cƈ��jV[n[��J��ʗ-�r�����±QA\�b��E�TG-�m��Z6��[+[E�[q16�(��Qb��E1(��h�jQ��"��r��Qs3�J�R�ŹC2т�-�`U��*+�a�F
*#�,QC2�T`�q�Q+Q���j�R��e*,b�Q�#mb1RⲆ[�(��m1�q�*X2(�X9hc�\eV6��[��Z�"�UQ��*֭jA�k*��*(�-����V�U�kU�-mp��n�=<�!���Ekד�.o�w*&��9�l˧o�(n&9� \^��Y֫�9a��=�<׭��H���~
�R����Z����~�=��<79z��:�[;�v���pz���ly��xo�K4��X+�C��@��>ߚ��}cG�Y�����Ȍ��}h��!�t���ڌr)::ӝ|��8+����&��	�����0<!�M}�k��\'P��ȤGS��dx(��W�A���q��2iE�'��|�'�w)�;��7�B����C�R~N& ~9�4ϒ|�M%G��`V���_�T��&����w��'�=��s�o��Ӵ_r������|�޸
ACF�}�m����O?}�^Y�N�è{9���9i�jɈ
)�}?w�Ă��ýɴ�'�v��f9�X���ȸ���ި�zb�ؾ�w_ﶗ}�����A@�h�ڲ��K۽�a�Y�&�1���t�aQ`}��0��Cܰ3���S��ņ�8�3�{�o1v���Llx	���QF������{O�{�C�d�}������4r���+:ɽk URq
�["��h��}HV����0�8��_��<a��B��7ܓL����ׁ�������ȯ�@͝(�~�8�+o�����?%zs���?jɈx~��a�1�q'��.Z,����1"��%E�La�
/���p�&�����'��R����;�}����M���������m=��?ti'�z���$�}�>!R�<;���a�P�~�O1Xo�Md��ÔRc���1%�z��Xq=ݚ@�R���q�L "@�$}�Py���t�h�?yƒÞ�CI�'\����a�a^�~�5�,�%v���C�(���p4��eC��a���*��,:�H,ǈ����E'�Cz�`t �� g��e}J�8�ٽ4g#)-�qc�&@�~߀_*����u��q�u7���J��:�m�(Y�n6�`�J茊����&k��{�:E�ӽZ�
ީ��ǧ|�U�a��$D���8Yi¦!9�jzF�;78k�݊6Dt^��_~�� xv�McE�Q����a�O㹓�����D��q�?s1E$����蘅gY9�a��p��
��ֲqI��a�{��T���!�4�q�h�ϤxLxTU�4�3_G�'yp�;���ė
z��i1�T�m���8�E�V2~eC~ӈi ���Ϸ����@��f�u
�ݲb=����:ώ���4�d����(�z���p������G�&�m��d2�½�"O���\C�)�&'��l�R�4��Rz�&3L��$��N��a�RA�;��^!R�����{a�S���6�Y�g�J����RE�w��u�Xo~W����� zc"C�w זzɭXyy��JɯlrβT5�aY?8�Y���4�2u�Xi�0�z������Ag�����N�Ag���i'����������x����-Q��#�c�DG��U��>LH/��6ϐ�?0���}�i��*bw��A��Ѫ��0�����Rc��&0�TP���I�4��+:ɿ;��a�
��:g�W^�2j.��M�% o��l1����*�:�~��
M3�>�0�ԅC����x��|���~��񇩈i
�<��Y+*g�S�i �Cs,X�I�ɭ_ɤ�B��Y=���说�����o)�"G�G����7'�$�
��Xg(�q��﹆�<J�����u:ɴ��Xq6�R{�����'��P=;�6����I���큌�&8���LE ����{�[�\�o{}����~�����b��!X��I�9�'�z�|�H,��ﵢm�%E����u%zè{u�Y�Nj��N���<��ݝd���O�<q ��4O��zɧ>�_�������3|�������a�
��4�Y�����s(�S,I�eCW�K�!Xq����>a���3l�ΰ��~�a�8��{�H>Xq9�6�8 q3��{�7����ft߾w;*�J�|�錀�ި���x\�:�!��$�
�a�9��=a_ƨ��:���ՓT�o�H)+4g��|�ꐯ��m�&�u�&!�)1�0�be$����.�|����3�J�A�:3�oM{�tJ�MT8�A]�y����h���1^�aY�5���;�3[��J��]DVV��]�����%�`�V7r�Go�F:Ĩ/q=�ɡ�	f��EA|����h*� *�kvJϥ]���{����W�� x����o��}���l��� ��1 �O9̆س��a��u6������$�}�+'�$�
͚�g(�q�xo!��zɰְY�J�]oߵ'SĂ����kϏ߻��oi5�s�Ͻ����k�2<:<H�M���� ��:����z�H(jy܇��.!Y;�3��0�(}n���bAN*���
�̰�:��a�r}�<#'�=�����I*�>��u���ݞ���K�c	�����>Bp�܇>d6r��OY>t�|�O�8���Y'���L�27�@a��I�I��VO#�ǀ����]��o�+o�_՛�ծI����c>d�ְ�Ì*o�>CIv���6�8 x{�!�J�>d���膐�J��grJ��+:��y�V3������M!_�fd�� +������Y���<�K�i ��7�t���aY��3�����É�h��&�&��&��uH}�5u%bͧ�1<��J�I�+<���܇��ٹ�§<q=�6n�Ū���v�w��D�<;$D{��;=��@�WL7�Qg���cY>LH.������/�4�V�OO;�Si�I�>ͤ�
�S��N�`�B��{��P6�Þ�{��<�5J+A=�|m�[����x|�OU%}`Vx_�J��+�k��6�wf�l���8 m+�`~�q��*u��<5Cm
�2yۮR���`����#�xD{`�Z}�ߘ?�?�s�|������O�;;ܚH)>T�n��K�B��;��Cl���xw�3�z�3Hy��H,+u�C�bAݛ>��H��+Kg�~I^��>��j
����_&q�`���<������M�Y��I���6�{���#��g�����%`*��u�;��g��x��d��ɶ3��f�:H,�LOǴRbAa��Y�}���{ʶ�˃�
�/��1R�>�?Y+|��`��*O����ϵ&�����Y:�O���`��d�������<J�?�Ch��J�g~���OɌ'}�$��d�.��0��H�~?���|��9`�����Dd̢v�K8�V����+yp X��&�2x�nT�ub��b3�z�S�83!����F����T�)̽�V,�mϥp��@��y/VƎ�sc܅��p�C*s���iȳ�.X9��y2leR=8r$���-]Z�V��x3x�R��K��@���?�".�E!�3 u��*oT��.���IRz����Xi�*J�����ֈ(u%z��N�R��;�ya��@���F��>d����\�~��k7�����}���&�M�c�w����T�4�u�B����릲o��AL}d�L��(bJ�Rq�7�6�R_�[*�a����3l���O�@����=׀�;�����;�w��}���ă�뛇�<E����,8�Cԕ�|�{Ch
(T4��I���N�B��_Xi�a�r�;C�J���1I�*ANh�}G�� q�%|���wVr�S�IXq�&0�?r���Ͱ�:��QH)��C�T<N!�<��C^�+bz�>��>J�����ɤTXT�'\I��xH<�ɡ��<xL *�V5��P5N�c���߿~���~�qc%C���E����O!�ri'�w,�O�w-�+��S���T�Ag��{��ğ�����dX5���0�����״Xi*OSlՆ3�I^�]g�o�>����Ҋ]������>�@�>�׃�2��o�y�9��L*O{���C�f�xo���'�>�@�N!S��w!�2��>M��M�2~�4��w��u��3�R"@ xDxg8�l"6����Gﺫ6��/,�՚a�P���ɽ��g�o\�i��F��P�|����~��E�a]v��i�W��wRx���ɳ������<���(��������1�|�l.Ԋ�x��m���"�g̕����=B�0��Vq�0�S�t0�?&0޹�����x_��hq
�CßkR|ʇS�1����k�JŞ&�&��6 
���w�B����U��nL�����a��N!��CQCG,]0�
���.��Qg*jZE�N�!�T����Y57�M}HV0o\'S��>��*O���#÷O��=�[y�j��`��c�~k����m �@�39����I��^�1�*J�w�m��C��a�1 ��O5a�CI�-�g�A@QN�d߹�����5�߂�k.qoAz���X�]e��f���XEv��fn��]���	��i�M�{���t�[Ʉ�`��>��j�KUq��*ϷO�a���1M�.ٲm�v�V�`��ّ���,�5�N{�M�����*�]N3���50E��PL��aK�#oI��W��}�ӝf�,�������xL����'��ri��]�s)�;�R
k���hx�����CL?*��g��i�f�͜Ȱ�R2Oh����ě�����E�C��z{�~�[�e���{�U|�P& p=1��h�� (��ߟh�|`T�|?{�l���܁̫
³u�{C�4�2V�riU'�+'{f$�6�0�{��a�i1���:�H,�;��=��/�ߦ��^���>{��{��T8�E�S=eC��t���V,��� x�'����l���{�i��T�'\O�����O;��Z�VMw�x�}d��i<��mE����߃���^���B��{y�g�@�*������!Xi:}c�N��̞��Ğ%E��c�a�y�B�(��4xý�ĩ>L}�� VqRW������P�s�4��1�������m��o:{��IO8��ǽ�>Ͻ�.e�OO�4������H)<C̥d�s$*~՟�i�'���~���z�]�l�}�b�R~�'�����}�� 	�8������pc�>���W�}�]��bAg��;�0�0��|�m?!�������E�w� ~J�0����L@QOȤ�0*<C�N�rO�f�z³l9Gm�} Lyǽ0-,���A�SA�s{�����~�����6�a��!��g\a�?s�o��a�:���C��i �gu�P�<C�*);����OS�)���sTS�4��*=��3|�bMꘋ0��N��w��Ͽ_?�����u�t��iQ�d`xF����yǌ8¡�ϰ6�z�QgP��d���N'���Rx�r�s�3}�+���I�8��̦3䞸�IQ���k2��
�|�o��<}�s;O'�]��"G� Lx�
�0=��9>T���&�H(h7��&�0�������2wVC��Ҥ9i���ɤ�7?w�Ă����&ӌ���C��>a_̚�4�^��~���~\��띿k�s��}�8�̕�;펨�-�VT>I}�݁�*�}a�i ���wAY�����0��Cy�5�ì1�ņ�8�3�٧������g>߮^}������+��T&��tB7����Y3�JT#���t8/���1��P ���o+E_C͞�I1�Y�w�	*p�*���M'9�s0Z[�F�|���짛��Pf36��U���&Z��$���#\�++�˅��6vn�i���Z?{�������j������������u��Mg2
�����*��>B���ְU'��l�Lg\a������1����<a�q1 ���xé�8�E��=e@p/��7��[�G┓8��gީ��f��c@�W���|���VLC�(b,4¦0��]$���˖�'�0��LH�z�Qg�Ն�_Y53�T��Hj��{��_�
�|�}�}{n!F�������Q�܏t�PN�3g�:�O�o�4�Xk����� �C�w�'�?j�����m ��ܺk%E ����8�!�Re��N�É�4�R�-,�ދ6����
)����L "@���I��g�eCI�'�����m�W���M{��8�]���>�AI��ěVT1���!Xb�]���1��(i�������qz2�~�����QD02<xL l{�wi�q�&�3'�*%C[��oS������(q%v���oD�+:������aY�y�d�6��+:��� *�*_aI�c�����V�;�~�~�����<�+v�cY�bMS�LC�*/��1��*7�:�����}�E�'b�~ͤ���d��^�*,4§Y��㴚B�zs�5�,��ì>�ݼ�{|ۺ�m��/�G��c#ޘJ}���t�i ��h����2����P�n����~7d�~I�6~���H,o��l�T���~�$�<a��bT��=M�uY���'�m��O�}�}��rW�%E��ۈx��0�������Mj��܅@�VM��d�
}iY?8�Y��<CI�'\��va��zɳ��h� ��J�~��I�(�{���S�_���鄻�k,�?{��YP�;�`o�B��Y��sl��
�M3�4�TP��M0��LCN��i�CF��8 ~J����ǩ�La�Y���%v�p՚Ol1���>��"����q{�!~�gy�5#�'��=9��*�:���H)6�8���7�!P�n�����1'��
�z�����H,��<�QN�����,X��8���]���W����b�٭�`؉f��^E�ײF��]�&���Q�/�/f��� ���3gG]N[9hc@u�ל0�1j�V2r��l�R��x��x�Nzs��ͳ�.�m��N�rˠ����k��-��P<8�2��0y&��;��ˏ{@�T�:�[Y�x{� kL���=D~�� ��3&�@Qa�*ϵ'�$�
�����N8��~>�@�+�J����u�h
/S���8�$�9�tyd����{��~a�Ri8�����|�A��Z~l;��F�-/�@�� {�.0_P�B��I�>��YI�i ������6����u%zè{u�Y�Nj��a�����ݝd�u�
|��ă�{�5�Z��[��[�&�߇�p2=�3���:¸�St~��=a�SMd�QH.�X��ʆ�p��B��繁�|�I�}�4��1�aQO�f ��<&�a�� ����}���Ǐ���:K[2����q�0 P>�2�0=/��&3�5��(~I\Cg,4��+1���B���j�#�N�Y�Y1UI�`i ������0���!_P�>M��<LCZ�g��~g��y{3�)��x7����� (��� D,�OܺC��1 �Og{��x�a�<�u6������ (��>�VO\I���yE��0�V���Y95�q��(����<��9WQ���ϙ�{����}����.�<<��~aܤ�m�n�:��=�3!�TR
v��L�����k��IRq1 ��UI�̕�C�+�|����o�O9��n�[�}K�&~����>Q�|)e�(� l
��$�vu�����4�u�� =�I�>d㛼�l=a^��w�i� �����l����\H)*������R<& �u�:3���w}�u�e��qT<g�<Ld�՘���|¦�fXz¦��`q�,<��P�,�
��p�$�S�L�w@i8��%풤�
γ�]����B����4Ͱ��Ri
�G��s����߾�ÿ�׿~��zm��*�t�1 ��9�t���sWL+?&0��LO�1��S��E �jo�u6�S�bC���ԕ�6������J�I�	�j���^ ���É���l��r�f��߄����*�?W�</�C&8��i�@�WL6eY�J��{�5���іC��<e����i�aܤ��i �I7ϳi<J�AO��$��*�7����ן�n������}�m�'-�Ȯ^�5:\t4RĔt�n-�X�$�*ՇVi�/'�Y,,���3��I��ܦ�����g9�J�0����n^�W8�2+�v�{��3"짵gPj�:�g[e<�Kw�����0Q����z�/� <!󖠮l��� l
��?w'���LHl�u��I_Y*,��$�x������m ��0���q�@�Wv��l�%f��1�'�b&���'�w7�B��
��?}�]��N�]��Z���Y���H����C�2w(�}�1 ��{t��.�
�9ܟ*g��y�������Z�É������@4x�(��Cso�~��w�d��U�,����X{}����4���؟����`ןF��{������g=Cc�1W�a�NO^àwo!h	�1l�[8��f���sq
����cw�HҙФcB�L�/�9sb)����"T<t�[vsa^�RKia���H��l���,�[,�=��X���֕��	q-��K��*����3N���I`��?*�,����t-���Heyx5����S���SqEggs	΋�v�H���9�3�g1c'�<�ũ�U�'�11^���ܚ���ݘW�D���}�����u��Y]Bc�BR�α��."-��1`�m����0ԑ�[S�����s���nQ�d��g��Uf��ޙ��\l�W������(X%��7�vv�<�8ʐ�b4 �aQ>w�z7}�-��q`�a��������b�{��e$�F[� q{[���*��y=����57��G\�q�&�٢D��ᆣ{�RP���jodجJj�=��	���z܄�<D�I�/���ޫyΛ�z���{��>/��z����_
�#�P�::��eN�Z�\S4aZ�<��f�Щ����\\��+�*��W�%q�D�Ó���5c2�4a��JVܶ�M��:f�Κm���R���IDr�xѥԸ� +��g��F��'�� �����Xq�Tz�>=���[)08���;��eֈ�n���[V�?�5c��� ��rWv�ͼŏI�0�4�B�X9�ũ��z�h^C�u�&˱u6�'Tߌ�Q�u��cYH���[�VB��}���ȼ޴Ϯ�P�_���_Xu�'
��6�n�a6�_Px�q�i�o�+`Dd#:.rf;�����u\7:6r�a�����Ȑ���;=���JH��nY+��n���Z9�
��*g�G�'�F�0�;;~y'=���܄Z�
��Ȝ���y�<)\Lu�B���t�/��J��4�+��w��L���������y@&�c���g�1��fˁy"�V���<~�3�}m`}�n�x���w
Sks|T��4�A�.X� R1(xu�'6�aZ���`�,�@��	��m�kX��p�τ]�Le�Ro��{����������c;��TG+>$HT|'�S��y.`C���2���D�i��k�]���v�RO��a�[�������+�Bo5��ը1��W�X�V�jv��N��7��ٮU�����A賩���e�2<�z4E���6�,�Ko�ݸGMy��Nx�[^��:��;J��hm��<��SZ!Q$�W�"�@�B��<`�����Z����:|��s�}�Ⅾ�t�6���B�..���1�F-_k�Vb�Ѕ{jB����P��
�ڵ''��ʟ?Vˊf��jJ�i�����qsN�0΅N���14�F� �ߤS��ٲ�c�ϗ{eӻ'00M��MI�J���Ҽo��}~�hϯ�0zP��WXt:T|+�_b����V=rqzT��{qduڃ��j{$%9n�9�Պ鞒���J4�w���Fys��4�z��8J/D����e��[��(�Z��z�B��L�7z"lb�U��G��.��k{/��o��
 3�݈鬗�M�
|��,�y'|���亄�ʨ���P5��tS�:?$M+�`!;��:*mO@�*cfۡ[��)��q�v
������&�ܞ�"����h��M;r;v��U\�'`U��v�މ�G `�=g���P#o��Z����nV��7ܧw>���M4�d��V�YR�����A��k$��ӹ<��maj��[��
us6+,j���Q�,]3���)]a��u��we3��yV>G;�j9A݃��Sp�����mn-qE]�G��x:\qn0J��ʇ@���һ"�.���L�	�&֓{��E�a9��&ab��`�Eμn�L��m���('�,�3�p�u-���n
�Re���Qۮy��V�uA�,�V�&��y�s�� �Z�?��R$��K�.�b8p+�om�3S��}��AU���pǳ��){:���Y�SJ�Z�n�B�V��Bl�J����T(�ݻKp���ʠ�9��)4�4��v�L+oҏ��ۋ/���]x�_�p��s�]k�f�շ��st���/��7owV����u3������G5!��R��)Ȝ3�L�����&�T�+[pX��S֐��<�,wnۆ)�<$�;1�p۹�Ae�z�He]��ؘ���'Xw,;��}�[������p��ep!7�;,��3i�Ch���^ް�x��M��Zal67>�vҭ��r	\��.���L��XFӃ�m�[T`Ud��,/l����{L�"R�V���nvm�n�n�������LĄ�t�|Fl��.���#��&�r�#���Gt,/GX��>�y{WI"�c2S8>�N��7-ʂ��$@�4j����V8XV�@�A�od��j�����\FcNA��
�[9_/\�;���=,�L:�fg;�CZ�
�o�k�K�L`�Y��&ǔYe�#�%��y#�.���2�gu�����;�Z;�*�ʓ.�lF�mb��V�T�b�&��Y�5�b�J��wj����LQ1���t��xn����t��Նɏ�W_H8p>�k]I҅m�eb�X@�����kl�.��ITk�rU�T�J�Q�p����j�H"[�uFe�WXH��h���-�l����k�#OHG�-�vͻ%� �]��#���Hvl�)�Y�E�[Yw '��77�K;n�`R�;0�{��� �F���C���S�n�JΌۭ��"��w�fC#�+0��f��Q��������X�2��t����������թ�4G"�H]i! /.>�W;;]A��*�P���mH�G�5x-kPp���X����p������T�gm�c�h:5Ȏ���8(�K梊=C���hKS��q�7U��|һ�=�g;$��=�t/�U���# ��6e� Ĕ�.�MS�5%8%՝�a�;[%�܅��k�:[��#6���9Ga7�[z�����F��ը�S����t���ޅ��Xnu��(\u�˰�I齒��[ۭ��S�o�ow�a�,�աB��� J4@AL��-*.Z�#W-b	��SDAX��-H�R.Z�R��J�V5������R��Le�
"�؃**$bŬ�Lr嫍UD����"(���F��j�5�b*��mmX�YQZ�%�\1����b�5W"��L�m-*ւ8ؕ�h���(b-%��Lq�QF��(�.R��ĬQKk�C��%1����-b��DVcQs,B�Qb(�h�
�D\kjfe�WJ�-ZՊe��j�mpiE�TLL����V�&!D�����"�D��(� ��1*�řK�1*�3\j����mC)U2ֲ�PX�J���pk+J�R6�r؈�e"��b��F�Q�j��*�C�,QFQ�Ʋ�j��Z6�ԪZ-�T����cDs
���`��cLi[-�Z�[YjҲ�X��[Q��Ke!inS
�QF1��m�ʱQEc�TA-�J�TV�e��V_�u�+q�M� �g$0h(��m�j�s1�z9�u�K(�.�{s�z�B�gGӅ��]��z��<�ݲ�Q�yҿ�<����E��b���1��Ίr��%z�Äf�2�*���p�����̰٪�j�<sN{��#���R��s��Ϊ�.��<-Z�#e�J��N���twq�'���R���V�,�w��7l��f�*W�<)�O� ˣ��X|�U�X}}g�Y�V�-�QуN1�Tg]�ǽ�G{��i��aB
D����b������h|��~�=[7�	��ꊹLI�ڤ�*�μ�v��+�s�+���
T�'<��W����'��>��P6���tl,j���!�6-��&�`c�n3z�x�[3��W�,��&i)<:�!�ݚ���16�UC�T�!+��S����NWaQ#S6˗�;�J�^�(Ҍ��+���%Vr�U1WR���Q���؞r���7�Md!��֍Z;�����65����ӽ�z"�G	1`T�������z����7��v����r޺�k��c��U��7,=7���n]�10�%�0;v��FV4;���|e�
�oC˙$ڄ�Ǣ�#w׎���V�v���R�3����n�g82���T3��j�[�f��3�1#�_?2#&�n)]'�E%r;�k.U���l�7����W�GD)�z�65e�0�YsX������/%v`Js? <<5ަ��ki"|.ū��FzMQ�#A���
��c�g�=�{"�R�<�W���z����smœ���Q,r�(��V5s�AG(��AFVS�����`m۾�ۮ�i�oc���X&���!.&��X�I>���/���c�������g�5�<�DoH�F#��gw,��`���Q�tK�L&~�F��j����US]��G6<�G.U5QĶ��Sиd6�nIО]M�LG@�0D��b�ȵ}}tn^�W�A�,�V\T�=r�v*�z3Aw�FS[v�����8u�5��MuÑv���NĸN�f�
��$C~r)]r��Ww��q�o�ő�x��	ـ-�u��њ�ᚼ]C0M����곢��O%(��%/��`�s`T�YC`�b�h�vؓ�טrH޸������9�t��{0�^A�RG{����R�A��V�)��-�䜣>�n��{j���1:p-ŷ{�h��v��'�.ݫ�F�A�dl�\�IW�VԧPi^#(�j"�/O`K�l�C�Nmm7yn4}��Y�\%�]�b�l��=<}��G3�b��)��Z�^+��SzoI���N
�sF�h���/CL*�%�>�J����m��:9y�H���ʠ�:��1���ff7�:]�QX\t��a�8
t/��]�t��Aw��vDVgm���� �(ͼM@�W9�;��v��M���f)uz&a�A�N,WU�9�t�3ft���=w{S)�l1.�]3�`�,c��8��c2WLmt�J6��z��=��{RI]�E�(���n&,g�n^��r�\D[��b��6�``A�=:f��|��H��*s��<Y(Z�.�D8��DYT'}�^�`]�^W�e12���ZP��AI݄�R;9�(�8��]Hzz��!,b�ߩW��|p��k\���l½Ǟ0��0���+��/�V�(��;3��njyBP� t�T9P�k�[�dAV�b5�Y���TZ�UQ���^�jF���{���ϳ�n�T;ƍ*�\
�p_�ǛCJ�J0]��&����%Χ'(�P���j�i�R*�gr��a��0�Nx��WCaW�z���=i-�PMXC��g����y�ϻʸ3��C�6�u(G����֯�ȋ��8y�OJ�K������VFŁ��g^)�4�Y�(Km]Bs��C�ɦ<1�b����̛��ղ���l�ܒ��&�9-=a�]����Pk�m$��1��)� ��=�^KV�~�:��b�;۪��(�Q��j����X���6gJw+��0�d��w4{]4�4$�tX��s$�Jd�Uc]��F���}� <<,�5�N���������*�t͊Rs�(_��S���bt�a�8�'��r�U���?/�������%�(�P�W��Č���XP0��70g�BT��{Q6���\�d���Ӏȳ�q����X5��oj��WWb���-�ǂ<�O��t;�ZׂM��W�$�Wc���@�����dd�_B���jY�FA\5�s-�z�Z���P?�h��v�ٟH���iŹ`E�B�i΁��Κ3��lb3[#��7�"﷊��]H�G=s}iv�:��MMy��5·��`��Z�L���m��l�;|�r�aL�k+t�|����UB��9v�����V�tͧL����y^��R��3�P�� �rs/�z�.Y׷j�ӭ��!��"�+c)gjԜ��*�4pC��O�e��G?O-v(>s�et�x�e�t���j�!�"+�S� O�����dcަ�-�k�.��M�u�zW��a<%�]�/�0zP�Àâ�Q�i}���;i��rh���m��9~��*.���5.��.�Cz�@+-Y�7�Grg3�5R	�����)�>4�D:��GA�)��"��c �>Q�1���\cmg>ӛ4jOnLG� �5��������Ό�b��]rݫ)����3u�I��I	���aG�kƧ�������<�l�癵1�ؐB��O��T�G��͉��]���]J� ?Tc�#���K��v���
.Y��w�&�[�sN�5�W����i�/t�S��⾱�5u{�D3�+o]��;>���&P���,��{:����a��$M�&������[Ţ�ਈ����:�c�q��}C�zwɊ�L�J��YXz�B
y��[K�{J������zov�5x�(ӵ[�=G��mP-�n�8R�U��m�`��{<#.Z�ih�b�e
UZE��j�}mX��	&.��q�z�+��K䐃�!���;�x��07l��f�>���c&��6+D�0�k�l+=8o;s�	k�����W��1Ѧط�`��b�~iϚ��;��*TY#؟�ʲ����q䐪	��9��Q����Ę��H):
��;��k:12������;k�9�ϸ��fd��
\��Ej[��Ѱ��8���6-�Л�� ���Է�>ڞ|0L�7sjz�H�4.ʍ3�[=�0��w�#Ϥ�t�>���dg���a@V�*�p�e)w\t,cNOy���;��P8��@Oz�q��K�/C k;��hFFR�&5��n\;��&l#u�-��R}��	�1J�T�
p�&����/��<<"ά��KwuGΨv�F�%f�t��c]a#��mu<4tҹ�S�®��W�3�i��<���*G�X�,c��<��k��lO*1=b�:$!.]6����=��ՋcctvY=������Ç'Au�Z�(㾙���qӽ�{�D�Q�LL ���'(h���j�֏Q��@ǫׄ�A���e�Ϥ������=65��<�z"�Ϯ��1���t���@bg�b�Qq��Fg����K�M�;0p&{C�B�D�M-�U�]���el���U ��azx��T*Et�j���G;
9D�}+��Q��S�N�=���n���ʭ˸���(O��U.�����c�$0��|��/���nw�L�N��&�t�NF�O�%�$���k���r�M����T�9�I��V����S|�dn����x�����6Ty���q�f�rwU-:b:C�49غ�-EǶh�ec�eF�����{����WLي���Z�aUnB.���EBhVܷ7�Hתz�Ƞю���]�}�LNÖ`��EP_yGL��n$hq�{x��UlRb�K�3"S�V�o(�Lgh��^<����5�:=ۈ����J�T�HìN�(����\vI���q��`GGd���^�4��PE��-���[ܞ�[htd���{���{����MO�V����\t����0��l���w^!/S� 6꣼�;:3Z�3V;�G����i�\IF�`��P"������Ì�^�7m�<k�9�wo!hN��[YhV�I��^�E�b4Fw���;Ffҩ��Rb����)e�^�eZ]C�Vr�!�/����ݽ����޽*v�k�ݮ�h������+h�e��>T�bnFT�,���sx�*!�yz�qIE�n�ܝN�o<�'!Λ�袇_�i!�a��^�X�QN�����R�>���ZTmt��s����3�`�,c��8��:gT0$�11��W���6�.�C�j�o���N1t�0ى�*����bm�R�"���X-���;!=P��;u�.]��:�%&eq}�>���]A>�E��Z�-ֆ��̔�(Y-L�UGw(���_F�d��H�};u̗ە�x��o�e\����k����گƘ���sǼ%|�t�V޶����﹭\@笩��P�J��:�9P����n����P-0��o���'z��(�e��!�@ԃ��#z��-F�
�_S�Yz]�{��W`蹰R[B�cQ�:VX(��H�Z���_}#�Xq����$< =��h�rf�pc�d]u�J�x"`�cۣ���������3������L&S�v�V�=��:P2�نi�l�w{BBr$w��J��=�U�A����⭕[�r���L�!lc&	��\S�Ab݅���܇0� 9^��R�<h�ڷ��^5�yB �ԳѸ�(�C�ߤ6l�E�<q�LB��y��������o�4Ng�Gݸ[R��c&3�I�?X�ɿTِ��#`'>��7�O%�B"������{a�����J����Ǩio�G�ɥ**���B�!]"r[�������`k�R7f��/ś�' �e�M���Ln�?Wk�	{�u�|�ig��s>��+�,˿x�y�v�2:�R��R�`��F��*[<�;W��l�j����Z>>HXLol1u����/)��a�b-��N�����k7�����c+bh�9��73�x��D��s���_ADV(Q�>QǕ㗡�q�v-:t����,�k~W\;���@�g�j[���e
���l͊�PN\ـ�ʵ�n��5泞(�:+q�D�S�B��2ó��LЕ���X�H��6:�HR�S�7ۚ�{W���K�����h{x��)��sU%���+�׋1�vnm�w�v�\}�-t��Z�]**��8�����1��]�Wdw�Vgq'�*0$Ҍt�}}�Ѭ�(���� x_:z�4��d����:СML��B+y�U=��:}�5�`�+�w	�TKI����s��r���Z&`�Ҭ�� ���B�B+�62�(f����)�G%m5�J��y!�B�<�L��F1K�[R��{�Z9�U�Y��.=u�CֵO{�ܹ�H�b*P0[��W��Qe���r�1�R?�.1�J���ٛ����N��w_[|��&]��fo�׍O���`�C��u�y�S�O��U�p8Vc쾹�P��7����f"�����{*=��Ҍ�(��jv��!E�3�8�1Ǯ$�dྺ�p��of��h��o��S��G�V�Y0�N���U.��v/a<V���;��g���P��2��]"���",���Δ�O����~"����ҝ\�X6�f���U!��	�Vy|Um.�+~y�uL����}v'/Lk�j^.��Y����nc@,�c ���6��꬇��KH��ҵ~>ݿ�e	�2��l� v���b��Ҡ2�@P�Z����;�Z
����}��d�t�y)ѱa�y��G,|��Si���ӽ��MY�+zr+�wc��$\;��U�Z['n�U ���<�s��	\n����=�J�΍��O�ᱰ�����}_U}]-kOp�S0~zptg���=�hC�}7O�f��}5xldϔlN-�[��i̸�/n�EЕ�0W?]�u�ڎ���C.�V;Y�3FX��Κ�O&c2����4���x)��fvL[�.�QB�&3�T���*�μ�v��Ψ�;*"%��Y�f���v/yL+O��)��*�U�P�G�2����i�q�!�:l[Uo�$b�2��R�{z֭j�m�ݛ0�A����ԭ�-:�X�?#k�1ᣜ���[~ߎW��Ϋ)w��R�������c�Q�t:��<��Н���
���仚uzx�D�/�K���w<�.��R��8݌s�:w�LO�|j8I���r4긽��Nwu����MB�Tz�|�T/��F/c��U���
z<o�Y�1a�y4�&Ş��tm�����:�Qr3Р9� �b�ĻQ��MQ�F�Sy.7n���N�vj��]Z�n�^�&�+�U!�J$E�.)zyM�ÞXZ�u �:�+8-�u�U�!_Vw����R���Gm/c5�<��U�jƪ��aU2�=<�7K��z��Ֆ��"����}\��3��!4Qn�ja���y�P�f+����N�4�?=a5(�et�n��R'c�|�{VQQ#���`�9���c�ʳ�nv������β4�dYL:��{�f�J�-��CV��Oޑ�̶�|��a�1��'Y[Vɛ�ggv�I�>�ƀ�h^���n�':����<�bƘH�t
3fݎ��	 ��������;T�ݕ)���E��I	[E*�6j�mJ1Q�Y����ێ�Y�P�Ř.m,J���lƬn�QՇ�R�7H�i����}j����Y̠������bK*�B	E�Ǘ �qjQg���jK�c�)�����n��7�_Q�`Ieg��m&������	5�f�j�����zUf��V�{���N�Ӿ"����synP�D?&�};D-(��%�6���Ѵ�p]$�\�>�����Kc������[�۷e��_->�����&7
ܻ=#U����Z/x�����Y]��v�؝�u��
P��43�0�u�E�2�Lu��*�t����"+T��*���+�@���pD�]�67{7�Wu�*6,���w���ws42a�:��:������wX�i��a�q��P�M���R�*�Քx�nY�ޒN71�mwlA7&�F�V��+�/�6nmn������)�*]�U��cbz.<-ʽ�����][�z�1H� �������!Rs��Ð$e*9����#�^���l����S���(�/l��D����Ԃ������,����m^�i��fV6�@{���b�,v-9�I����
��3��E��f6p����������kr�4�`��;ӷ��,����R�e ����];(�U��q�ce"q`���E���N�+�rdg������݂�5���PM}f�vYlu���;��V�²�WQ�k�Gٷ��KR�1�{�m��K%۽z�m�n����&�������e>����_�h'l��<*-�z�ý�3���`�nڢ�u
;��sd����N>���V�
�/�\
��.��H��U��g8i�X�YX6?�/���W��~b���1�K�|��C[�fa��tu-�.�d��rL.�R�� �ͷn�Xt��u|-F�]q�����ָ���w<!U��%i�:�BMhF;.�Z�cQW�Cܸ��'R2#��
��؞JJ1nԘ�]5\�b���Qw�I,
���µXv�S^�Ay��"�s��d]p���l���ɣX��O,!T�+��.H�_48�h�� �2�L�������A�>�j<�����Щ���9���\��(��Zt�v�:_��/O�T���j�y�)�G'��x���+^����
�;���3��P ª��Ӗf��V���je+�DF�F��TQ��L��(����hR���*�V��
2ұU˖��Q��,r�QKV��r�1,b��e̠���k[kKimK%m�墪����ֹn	b�����%�aQ�e̫a�W*!Q�p�*"!r���0P��"�V3�F��%F\��E���LQ�S3�m�Kl�\�E�mE-(堦	U+Q���DT��LƆ-KR�R�JU̙�V�X� �[�)X��ejZf+�ES-h�Ъ̲�S2�L�U�6�30�JZ��Z�*�ƣZ��)[KF� ۉq�fS0�8�mki`�,*b���.8\�UU�\��-��.#�i��fe�F�2��0[\�Qm���J.6�1ʊcL�-��a�eJ�s*-l[�(�ƎZ*Q�\q̩�d�*6��2ڋ��L���TY�s2�b�R�,Q(ʎ�-(�m[KVU�--@X�0¥�L-(�ܫan(����-�i�$�;hc���i�i��l���犿���J��9��j�qm[}u���&ȝʧ�6`�@���W�<��^ޕm�}�
;�G�������S��_8����lB%�z�lf?x�6�+�z��.�[S}��7ܱL�m�(�����.�L�5�~si>���%��-L5mc[��$#hS��c��0�8�3R��'�Sa:b:0D�U�Z��6f�m,jˋ��K���֒�$.�~Y
���E�4�хU����ݨ��&��� �gMa�T��ܨ9xj���ƭ-+���$A�T��I�bY�>Vc�G��f ���=����,���-+�"�&U�[�5�'Ղ[����P�qC1_�a�lI��l��B���#v��o�3SRFMu��Fw���;�fm*��U�=3�B�;r%��<6�q2�ӻ#GYgPD��fqP	#�t8��F{��X4{MY+j+V��ǈ>T�b~57�>��/^���ae# RGGZ��`�.puU�Iש�a9i�ѭ�1K}�蚨s�`��z9��0�}�p�Λn^��(���Nj�/? %�|Ōx��:gT�0$�Vb`LK�}��G�D�]�ޒbv�6��@c�\���{�\�Qx,��Zoѓ��zr���Q"IU�9�A�9Kѝ����2[�el��:�y+\�`�A[LS9����z�S�6�	x�um�3���=r�c�d�$�Њ�����xX�-�ɒ�o�zD���@��f&/�]��;A9zf���."-͍f,��Y11>ܧ��$pm�,��4<�T9��!Ŋ��P��NqyPB�b�Z�38��P�
[/'q=k�XV�L�0���%..���fP���9^�^��8T�5�E��df�)�A�䗆ND�L��[���ܳ �ᰡ;�Tr��T*�i#Ǉ]4�݌[�1MM�1!>so�=eՊ�X���*����w�>���А���K͛wR������焵�����yz'[�Q�`����#�!o��Y9L�C��DM�~�AT9yceNrFuI�go��}�!�p�]$�}n*,a�5LB�Y�u1jS���B��h��z�ځO�ZF;1$I�U/�O�P�S~��!窲6,Cs�ΫS}���R"%�-���-$�p�Zv�+�Ҿ�TpSW5�BG�^T��
�%C� �����Ưf��;*���%�0먺s�kV�h�u�K�[0�<���Q��t���
ϑ�.�`m�r�)�t������+{:P�����'9�X���䓶�>:3�`�0�MI�q�Y, m�N�ۚ�m��suі�W|��@�Tp�S�m�LfΆ�ih���`}�g���O+=k�}�-J��o���݅�p�q]v,�0��.�a +}�{[�T��ъ+&:B�!�;~a����ex��LOe�!=_���Z>��U^�a�as�X�{G�u�Vc�����u�
4�7:�[ǘc�ݬޞf�N+V���+xm:���2u���P��ӧ��u�k=�X�F�W��x��6��Zt-֜���:h��7L�FJ��ˍΔ�^��8�&�ة	�l�X4��j��>e�x�\�x��K��u��uE�"1gu�rR��V���f�`S�5�m
���v�����S�i�N���
#1WT�	a�Sj��EQ�{Xh��ˈ���Jg�H�nHBM�j=.`㳨���S�b�y�N�jmNd��T��P�s�2,k��˭�hD���aX�A�"��X3���s'Wrל�5��.F�c�-�a�}�\�a<'��v���S�����Dl���wu��Ғ���*�.㝘Q�kƧ��	NF[��q:�R�r��YBo�]X�N�"X1�%w�&o�0�,Q�T�҅�(�[���z�B��L��L�e�L�Y�n�
��J�u�j	�,v͢OL?Xr��~�`U��T5nW�uk0����f%��G��/(˳u7���Q�=m�ٽI\�Y�.�؋��l[�/���7��A��X�40�,b��(R.�Z����3�6� R���i;�,��Y}˴|=���k&�R�D��������G��D�7�P�x�c������$�,WS�$�̨�ԍ���y+�A����;C����H�8(�f߼�:��qkg��J�����y�K]*8�;!@��i�T_��:^��Q�O<�+ipo�c�O�<n��0_�t�#��ʵo��H��o����bsY��K����s��Ϊ�C��C������On���ڒ)\#���s���ѽn�dwZ�}7O�f��}5x��)B��N%E���(j:��A���o¤l[��<7m�F8�8\�����R��	�y�j�4]'����wn�)���V�ˊV�N��T\6$�{j�Rt��p1�8�(��A6����\��Ӑ�K.^��;�3b=�Ej[��Av��t1�>��{�d'U�m������f�-^�t��u@��h)Y�[�V���s���X�V�w�d���-`�+u�H��R��)P4ȧ+9�Ӱ�:���T6'��+��B�"�vH��疸��tm��%pr+�:i,_�k�/�o	�� �؏01ep�o3r����F�ԋ{S�c4�8�; f�)���)N�h��\�媙@���|{$���lŪ�ݹ�*Myh!��AiU������J�7U���i�����|Y-��}�4Ң~�LTY�x�K�ŕ\Ƽ3 �n�9����=�"�f����y<D�ot�J��&&,t�.���.�8��Fn;ߥ^��78�����n���j����J4��Q*�i1
E�0"���_C�$х�lNOO1]�t��Z0��j��kc��[yHc���Q"/�J�zyM��r��Et�j����aFxr�0�ǀ�5����h��Q�7��ٵ�k ړx�Tl�IbhYf!)+'պUn�	9�I��md��t�l�bR�j�����aN�P�ؗ]h�*j*<�w�aʎ����u[U�D���ږm�k}Y�6=��
Ì�nQ�˩��#�`�U�tӭ���̼�x�)+�_i'�y~��(���Y��^�Qcr���SXn�TXM�n���v�lG{}��'Ux-
`ƒ�qm�������/=w��*ȼ����U�-'f �ۺ��gt�pO;i�t��a�ª�jڱ	�){ţb�JUc�}'?����;��W�����ow�`�3y���-K��m���%�m�7)�w-W���?=�#�J��G3�� ��� ����2ю ��]�1�ܸ�rz+u�Y�������H�cZ��B\9JGD&����K� �n��t��Y�}�ȿtz��:�VI��{�
Y�`��R���?#`ţAl�׽5�5	U��X�)1J���\'��,/y<�9�uy�4Zx��o�8�d#!*T
O��6hlt�����ؚS����M�Y�ʀP�О�[�-i-��*1E���DB���V�o��[��'!ΛVb���D�UC��J��F�����||saӫBpR�����=o>��r�������L��0$��:֩��Z�Ή���BD�$��B�Y��]�����f���qnu��b2a�����"����A:g@#��J���EZV&�q���|+�}�ܻ��CO.�~Z���(�±���`n�eHѰMR�n������l�8xz���ag�*m�8�U"��6�]��N�d��c��9���� �B��U5�njsZЛ�(��oM�)���@�k�=�t�eS����ϛ��М��Am�K9ɬH�����,mn�/�O9*�J��/(���P\���).AV�(e/m��+�]{����Lvmy #��]d�\��{X̵dz��wT^���yG�^֖���GvuB�]�DG*u��X�**ic���,���]��Ƣ�����ܚ����a�C�yT����Pu'Z��a�8��nm��[\�L�Ҟ�/�末Fآ�#;�xx{����-#"�]]��@3}j*0��b��u1jq:
.Z��U�f�س�����֒&�D�6.�ȟD�B���`�&=�Vő��{>�Q3^�uz�xw�Mc���}�m�[U9��=��*V/��kʛ����*x�_�N6>��+�^�!/׍gY�������6l!��LW�������K���v�x�s)������U�4QT�\�`[o1�1�!�ߘN��}�Om1슈Y����\-ա��N��;���!�RXv
H����s�w쳞���b-�6�<�R-�y�=m�����geoP�y�K������"��5'pg�J+Ŭ]�5������K����Lیs�-:t��G��X�ް�.2t�I9�\��;E)�T���(�]�4�FɻpD���x�\��ٙTVk�|�7���/בixf�y�Bb�ں�T)�9t��:󱆭T��X�=] ���tRU��^3����P�+�q�]g�j�p����uG�eN��＼-�T0�d��>��n�K@��$ms?^�(��C��l��ge:Tg=����;�/ѕ:�����3F��&-1YGlCP�
����m���u�	��	-�פs{rQ޶U�����"J�r,�٪�ˎ��3�qT��z#6�9���xLk8����*�''}ε��X�=��Fx�L�W��쓤,"��E�_�������-��N'��[,Q�y�����@�7ҭ;u�*5�ʒ5P����J;�d]�+-�:k���OZ,�i������xГ
.㍘P�;fXɮ���Vx��]�n#K2�+�7�au�ˎh��Dyz5N
��J� Vʀ5�(C�Qr�'n��Y�6�[(Yu=�}ī*�+��w�'8��	�+�LΘ�(�9&����g�V�q]�����ȵ{KX7f3������B2r �#�8���H�8*R"��� ^v��sD��<�qD	M�]�([u��!��	����zh�QvEl(�V��=v{g^���<�����W��|nӔ6�.
{\#nZ�ڮ���\q�;��:XoqG{�Q�5VQRt]lu����{�e���Y^��Mזi��j�f�IkR����R�z�"��ة��e8�:qc���y���N7]�|qi�۩'�ŵ�T��:���(z�`w��y��^��T,��̔�|�Ȍ$���J�R9�B=݀�n�v"�wii@t�̎PL��"�F�;�a��L�@4��Z��xoz�s�:u�z���l|��@F��g@�ͼ�q�/��}��	-*<S�*{w�d(����S?x�mϗg�����}�:%Z]\wy1��>-o;���Ȟ��|Գ���q�H�w�^��;�3B��(�
*Է9�4�����WfC�:k��kYĲb�*(R�a7{ҧdvN�)Y�ZQ���X��>�;HD��TL��a-�kR-���NX���dS��P�|��y.�k�U����.�y�j�M�\��;��9��R^�z2����xʊ���X�t��/B�,ߵ���w�yq/{��!Y�7�������C��4XRp]\+AG������ǎ��V���;7�lׅ����l~�6���٭�8���2�%�b�ĻQ��MQ�#A����Sy�(�MMɮ�&5�c8��]"�C�D�����tTÕ�]3����alq]*��.e\���R��a�2�S���{���Cl�U.����V9��>�S#��������fܪ�2���1Y3��L�3��uޟ1�Ώ�+�]o&?p��T3V�3�r���v�N"�V�jJ���k8Y�"��f�(�k�f���]q�/�S��̑ҭ��/ ���*�;�i��(rL�n6\����e�ۮ���iJ�{8Bٰg�>kpG��@��&�����Y�c]����b9�)����OQ��H�[џ�sX���G6=��Ì�Sr��'��#``�"k��]�ۙ
{��,��)!;��u!l��#oU����uh�*����a��QQ~M뚋G^<Mrm��I8���3}�߷6u��m*�Bŏz7��9AY�>}��Q��=��q�F��Q�I#�6��`�sJ|��yG�(��ѱO��
N?�ݶ$�mg<�̓Փ�l�qf��۹��Qң�P�W��f�+�#2
��� �;s���nS��N.)�J���:Cr�S/�6hlt�%C`�m/x��PW��9|x��6x�ȋ�d?
��c.���L���U[��߭�v�a֜ڳ�ï�YSZ�W'�L��ߜw�����7�`�JᠡF	�x��1NW1B�Oz��R�"bQ����8������砄����U�Nzu7Έ{h'/L�9Z%�E���K��uv-��+w"�?&s`g��vB:g|GQ��!���1-+c8���.�.@*pD��"�El����5�:N�9��\T���Rz���$m�����+2��y3���7� �+Sf�.@�;���pmM����qr�{\�Voy�1Z+SUW��,U���X㛽��iݓ� ѫ[up�Q/�&���	m	]V_]Lū�:�*1��MEB_4��G�v�>y�A�c�$E�h�Sd�*�љ+��%YG\�i:��v�1]�.5Ѐ���ZL�T�uvE��(s�����KtwE�vw-�.ї�Jj���
���\��ո�P:þ���f�$�P��3d�x�y:���$o�-W���My�z+tҧŌLq(=�j݄��cr��s�f��G��3=���St6G��Йw�k�j�nmJ-��,0dξ�j��+�c�tޓ215d,dǫQ�ľH-%���'�AsD�����r�K��;;�\$|�(Wf ����i#4�x 8�#�F�Q����r���'�*�!y�hf;�!���!��o#�u���	X�ɡ�G�H��튒Ӯp/��Rq;ٚ%���K�cz40=X�W&u�3'k�aS9gJ��a(	�>"�7�G��c��ۖ��r�U�t�i��sy>��S,mK7l]�� F�i�J���;�[',�u���8u��+lSUX�OE���(�oz�4-w+T��g5;3�2�`�b벒���{ʱYbu<c����"z������c%l��X��B�e�k:��Գ����
z>klR�Y���S�vd�[x��x( �&�
5A�[�]�! k.P�]JG1D�0n�F���ɡm�"o*�i��;;{��,����*�Ɣ��zڳJ��B��޻��0/S+3����RB1u��p0�о�ܐ�R7�wqҩt�wv+^Y+���
��As5���kz�Ђ'1����~ڊWN ���/9�~�#��'D

`ޔ6��t0���ñ� ��6�r�E\y=�b6^�y{i�N�`�.�K�l���)�s�κָc�}	�dݶ]��wK�Oj�Q��]�1���>������`�rMT����YZK��V�)��W-��pT�Z��2�j���N�d��kzN��3� JӾAf��j�c�_\7wEH���x�w�M��jksD�L���������Ί<%��n�>ceՓ����>=�_n�u�R��YR��]I�\�[Y�,	�NFjð�|oD�zjҸ6���6��g��͘�V*�u�P�wQ�÷z:�\H�l㣽PSӹGp޼gpg�Q�svX�e3�!���t��㶬\�v�ֺǉ��ɞ�a�5��b�Y���ͼǻqF��p�P���Z7%s�#��w��}��G}�h�@��
Ž܆��Rl] ��O2K��.���Ӂ���-�Q�>�;+�S���.��3��l����g5��TV�e�[��MJ�FR���ڤ&S���j�����Ʋ�s&2���PFKV�)DDm����ʊ`Ԫ�nW*0r�Lƍ��L����X�ET-��F��h�Q�1���J��%���Т�e�9j-�[����mr���2��"�Us.V�0��m�*��S��L��kQ-*��cZʊR����km(�X����-*�+UV�KTqK��j!R���ʨ�̸�-�2�(,���J�j.\Z�̸�kEQhŶS-Ɖq̴m�01��3,��
��6֖ҴEU���ڶ�T�0��QRڪ.UˍEc)mr�lJ�V!�qDcram˘�E�s1EZՃl*Ʒ-�,l�KV��k��J9)V,m̨�̷,�KlEUq��m�5��++m�j�b�J�.7*ڥTYm�*��-T\˂�Ѫ�L����6�F���E��e.f[*��JcV�84���QU�1ȍ�D�9��2E332�����5�a����.YL�`���b[F"�+mT=���������x�����Y�MR�ua�P�Ex1G*��K��R4�9�ͽ�ﴧ�`�[�u'w9VJϊ���]�)uN�g>L�&�_O�P�%��65�ڬn�eH�}=ꐄ�]�sb�z��h�F��Q���y�h��T��ٳ
�c����ᰡ;�Tz��U`Ԑ���!n��N��\Uh�G��Zh���v0r� �k�=�����0��d���� �B�L�X{B6'*��P�ItE1T�穡�Y����p�J��5�ʹ�^۞�P!�s�cw2�X�iq�@aTd�ChƊ�$>��yۄ�![��b��N���"sP�T%3WoH��f�ˎbh��b�o�O�����^!����x���U�do/a�n@[��B�e��^�>S�
5wʰ��=�����L����myS}K a����+1^�<���~5.�eJ��]�jU�~j��ś9q1��_@�j��6�G(x+�Y��G0�Y��,u8��/���8��2Þ��3s	��go�'Kg��gj��1Vk�#E(��b�rx�O{�73|�q��X�b�guO��!��M�5H�|a�_�����^�+8JTrͯOn�SUd��[���Y ��|�|��=�M���5���6��4n�͎�4�#� 0����ټ�d�ʺ��`��L�2r�]"튱Z��T�;�Ӱ�Cm�!=�МU���W!��;PK��<r���(��4Ș$�29%���y����-Z�z��\SÅ�_pٜ珴3n1Ȥ�Mis\�=��h�=א��飢��&���"mM��P��0 ���Y����+Ͻ:Jz7S �aC�No.^�ut�$άcҦ9�l�]
nN��c�=�V�U�����>t����M�b���5�`�+�Y�	y��Y#E�R��v��*�ut�P^�;�W2Lk^.-�%v���0�թ9:9V���(\�L���b�t�X��=�#[�#��⫹��ƒ��&geD��Ϻ�(
�gJ�	�P\�ʃ~�hʫ�L����"䮄���v������?d�R�D8j��.]��fhK^5=����s��u���+�Ì]�{�Lsh��+�a�bE����N����K=u$^ҏ_����K����z�#^@o1�!#q�㫺U�i+ᱬ
;�x�7��H�����*da����P�!S�~���n��zf�)\����+��a;q�T�d<�@DP*�
:%lW�Lٌ�p~ף)��v��<=ǒ�����
�"'p7�{dȂ��";�4�pߕ�ۏwC\Aՙ�%�ꋃ�OO���[�%����+
�*��}�.lَ�)H�C��8�q���m�Jsf95�
ض`��6x�ݾ�j,���Ut�orV��6�hi���HHt�R��IV�T/f���)p�T>��*-:C��H�]T��f��|���+N�"����jMq��w:���zj��p/8�7:Y��8p;�k�m�S{Uއ*u@��n!(�Z���]z�Y�}Zt�!�����Foc�^�B}cv̌����u�u�C�����aI#Jޛ]����Hص�{�m�F{N!��`��b��iAO`�6)��s{��7�-�܆Üg��t�X�3D:~�R�����TU�bL`T�����j�1�V���Qpf��;YЙW�SW�iOA�"���� mKs�h,��՚��锤���4�����M�j�&�`:T����Ѿ)Y�[��bh�]T9����L���BܧG�#�_r�\!��
��S�#X��0%�\Ōx�	�(�$:��=�+13Ї�qv��iqD�W��0��	�F&眨�;j�I�u�^�@Y��r7c�7�W����RԾ��%z8�w^�U�5\�Q�#��e4ǉ�O�o�_�	u<����ν��v!�t4k>*4�J�b,{Eu] .T�����Ww���nP󫙚�?+ڍ�];��TcJ����!����*��ՙ��˹�)JW͛�sPv�q�� �.��h(��כLu��(ʹ�����@�Ճ�r1WS���v����	|k��ks#��}�b�U�M1./I��%T+�K�d�h56��
��&��ַSR:*7��҄�=��4/d^*Q"�����L9Q0'�=Z�g���c�mma�:�
(�Ht?s��.B��80�����8MFÀ8!*%	�[U-ʸ�9M���h�(��FA���q��7YȊxeg�6�>o��ҏ�>WD�sz��>��u��#<	�y&������u�4���9�,}3G�xJ��,��z���,T��(Y�1uC�bz*�;�c3
D�DVEC�����e��n���TX�:�aUnB.���EGL��=t��վ���j�H�,+�u}E}�|B]
�!bǽ)��/��bU�C���>U�#ȟ.
�H%��U�qv�WЄ�^�4�+�BVQ�*���ѱO�*��W�{n3�pP��]׽K8�j�<ï0��U�N�B�[6��f���L�C�f�
�ʗl ���(t2�1'1#.+�t`ڤ!Fr��<�y�z3͛4ht�^V�׈��0�-�|+=��2�BBǲ��b�b[��uj�j����]�I"�� ��nD�\�GcYCO��=������MY���R�5�N�N9l�6��f:�LR��A�PH(����_vs�!F���1�LY���l}[�ό�ڗ8;��1�fo:�{���jR69�~d���puU�Z�[�a9�Zptkj�R����uq7��7Ft�'�1��
�z��	�N��
`���	��+9��&=1�2!�N�֏/lrsk:g���堌u��h��v5]J�=9�tC�U�>�_�EV����U�f��o�p�!l�ыo69d!�H�0jP��z�}΋���C3A�|[�gU��5IԺ��j���LR��KS0u�ʮ�t�*F}=ꐄ�]�r����Y���0�zh�Km����0Y��Q�f����s~n��ҏ����*3�TP��g9�����/���i�&��6(�
� ��,͹P.��B~�}����9	ȑ��j5xpO9�lb�{���怬��i�M+�k���o�L�
�;�Z��Y=��sk9��;�#���hD�z��j�#iƊ�
 v��A�����?)�D>>���Ť�˽���6Ү��輄���]���*?�����])(,1��I�qU./r��׊��u֕�(z��X]�Z�\��\pǔ����n�O�bG�x����κ��e�,���fg�V�Qo	#S�S��.>�ֻxR�PK�R�wo�6i��.&ͭ�,�����ď�%[,���^�u��m�2����w����WQ~N���^M`�qu7��!]�3Y-΋���t�Bp(�X�4x�#{!�s�Gt�&%͆0:q1A�_@��W�%�E�YG���Y�sa��wg����6�"u�1�{pL��� {��}n�C�v���;]8�Yڸ�m��^�7�ۙ�L�ߓ2J*߾;k=}�P{����[�n�!��lC�R)�<���f􎵷F���n�Op��HJ�AT#��>3�k�����U�<8^%���㗡�q�H��뜺ʎ�9��s��;���v݊�[�aP�b�@�(�$Q�L���ųE�o�u�}���:�^v���r�k�Ʃ��[��N��:Q3P1OLЁ�6D�'E�B+���:A�t��G�5��sy"Gf���J�)��_���b�0�R�hL���Y3�5�+�R�܎�u.�S��g�I�(��ɱ7�`�;4��U�F)B�s�25ɋRC�}R��B�_I��H���^si/M�b��Q�iD�nB��@�u�*�'�E�]tʌ��{R��e�0�������-:�A��j��rWiT�Yx��Y���.jH^�h!��P���&Z���XmF�A���-�����y�c�-f���c��;Ǯ�).�� ��X���!צ�<�z��� ��Vouٴ7�v�")Oi��a*Ȩ��QDȨ���aL�(K��U{�\(���(Ж�j{$%9�t9����j�m��έ����f�紻-P��h���MF��1���Vp[���@���O���w6ݟ)6��O��~�s��7��H�:A
�3�<J'�X䗯|�hoSw;^�ʍ󃅔A�J\(
/�rɇ�t'n2e�|!�MT�"TMp��b����]
��=j��ހ�,[�x��ຄ�Oe�+��T>�7YP���ȉ�:�׈�"w�J4�}��K���a��W�L������zo��q�ntl1�\8��F��U�U4b&9f�98�5�sIB�<Y0�6' PS.,V֩{뭎�V63m߯v���]�1�7l�73��Ĝ������9"���O
r��)}�aU��#b���{���C$�eT	&́��2=��8a��=�:X���;(l4�U��V����V�']7�
�&$ᮨ�WVwTx����$�s���p:�A�ΌL�0�5zf����]��U��'�/���m{E	ui�~b��,�\�:b7yk:ڎ���h`���O�Վu�|9����oQ�7¬�X�ӻ9Ð �Ȟ�SL��B9���b*p��Iu�X��
U�u�4k�2�+7��B�\�@l�y�V�2�0$z��&�fn�=�kt�;�Q�"�uf<��mtض�Svn��w�{v��e��r���.�&0��\`|9"ھ�K��3�%�t.�V�s��9p	r�1cv$��k�uCby}�:�ú}*��iVı���(!Jz�	��؞r���y'�ֹ{�@Y���A2j�nM;h�=|�J��q��^v�_�e�;)�<Ү*y��o���t�ǜ��M��Y\ۮ3���Ǖ�GŷO&�������b۱}~�j23�h�o7�r��u��%j�!dە��c�3�<�ꅄ+t�q.rư���(���c��*���$�׹��u�p͇�0�y�1u*:�6���Q�. ����.�k $g2S'{f�EP�����i�A���yȊxg��xM��O���t����;�0D�E��	����_���`\�OE�Voa����W�G6=��;3��nQN���#c�p�D9���3KRH�P�~�b�1Q��eg��6���T_�N����#���]Fe<;9�T�6o�Y�����e���Y3VAz����z��
]�a�|�8@Թb9`G��B�؍��ct�czU���:�K8z�����\����B�t&�뉩o����._˖U�z®&��4�c���'����!��ڳV��b���]��rF�B�짌����W��4��J�!bἻ��{1^�{e丽�`���d^'L��DIa�0�7uo�c��4,2'��q^�Ʉ�'�q�r�Z�߶�⻊B����x�N�\.	�!�Uu��R�+T'+Ƴ(�B����U�p��%"Gr�a����Mͪbg*C�N��ýf�A�f�LՁ��i~�/]�����%^����ڷ����YSNzf��U[��߭�	�!֜�N�U8{��;���rȢ���Uv,t�zi	�N�2(>���DK�����F"-f�J�Oc�In��0��S������LU��W�KbN]+���.�������`{�!2��7��T:j��Ez�X-��9d,�3@�b�J��CBұ<;6Iqe	�g��k}���ض���/��3�&)B�	jf�]��n\]H���l
�!(y͝8�G�)"���̈́e�5�Ӆ�3�E¶l½�������K��;�TgQ���Z��v�^:wuY���X"���H�F���2���*V-�3���{-��;J�U��j�	��g�������P�n�]7*�b���ƥ���'+�	"e��y�{�<�NPC��s]1�������9��ҝ��Ѩ�N��%�$**�� l'꨹0����c3�U��k�<1ҁ���×]��n�hOz��}P����[e��$4(��UW��e]���Q�"\#(7�9Ir=�����'��S�+\�ۙ�F�lK�6��*�"h�� ����@r/�EE��41
��B�7��H�7�gWF�%ǒ��1}/����އZ"lo�4]u���|H^5֔x�×����;-t5�Y1V��TrQ�(JE!���ǥ'
�b�h����������Kr{uƱ�ͧ�QYg�����`i�2���1:Y�×�/�^��3`�ʛ�./L��-�p���(v��*��>�oLC�u
�.N�џC�k�;����"��� �lLV�s=�f��Ǆgs%��`W`�91b��m�E�o=�zЇI�!��oa�T��cp�U���R�m�¤Z�"a9�Aek���q�U�\_�ס������xp���[R�=��u׾|:��L��Wt*�(��&\Y4/ʴ�@��飵�A��x��6*ECu`.��X�׽WpqK�Wl���I���\�M֦�����1 �N;J�w��F��c��z�n\c2u>Yw.S�v�v`kk~q��`�/8�R�)v�V�ss�R��f�jq۝Ev4���H�f1)��)`ٽ�$|}���=�\0V�7(ԭ��[�ء����:�J�&�]�����גP��ʝ���v��4�Z������2�b���|	[K�}���@h��\8��2L��=�6�]����I�OUj�&��l���fI�N�Z� 4�'Wf�A��8�j�u[6�Crm��2���o�o Վ����Z�jC��y��	�B�v7���҈U�}��C��n��)�Ә�Yɣ��[)i����Gz����D�Ҍ�R�+��7�}�
�j����|+0����ѥ	��i�孙�RZ��UN��Y�Ӑ�P�հ�Rb��&�Suq�n'twٷ�^<W]��U�0py��wqgfF�3�:��oN������@�8Os�E�����lގ=��G.�ރL��sј��\�^��=�9�[�n��Ƅ��X瓬ؑwNW,hvp�4�>�S=�:(�7BݥMC�Y��]�i��U̾S3Q�[o)��yf���vt�n;,bSv��"*�h��)N��}+F4g�Jµ[�N���O%EÚG�.Ә���s]YN��1�<�Xh��;s�U�����w�=N,Ǧ�:��)��gN�+@�K0����Z�>(Ʀbz<fS��_i�0T�wb��:�kI�V co@ 0	"�*
�_%�a�qp7b��!�����x���S���*Pgl�F��F�̖�y;2}����{�M�\)���D"1�p[F�Bfnf#Z��y]�r���έ��o�e��F}�lA5ܖlvX��a
"Z��#|w���Ij�l���52@O�*�X�9Q_C��i��v-|�Z��]Q��Pt�L쌞�`�� ��fU�C�����s�I&�=v�nk=2ػtWlŖ"�]����6��lgs�[]�ǫ>:XL���T�wRTà�э�p�mM˄$�����`�_^�[�'i�����yr��5D�\��W:u��h�������YT��v��6UݨYھ���+�N���E��e.5���EN���z�/ ��^�����*�&�A@no*�H1���4yu f�Wݴ{��;�*�N�u����e�r�(��1�N���,#���l���4g=�cع,?=�]ae�z]l#���WH�LWGfB&8�BB)r��R�9Q�kp���tySE�ظ�
V.���Y�7or�5��� �R6�RȎ�m�-�	��`��s���b�ȭkx��f��*��5уD8�n1��۩ã)r��'E\匬�T;���q�ڻY����9U��u=����)�Ż��m��B�[-!\6�r�2J��՞�:�\m�ׁ����|��M��㟋jX�
�cX�RĎc�iQ��\�[�kF�\̘�q˂��eE�&b�mJZ�-��+XY��1�d���1J9�,Fՠ�J����L2̂�e�P�̔����-1fP�Z\V�&�TkF�)�d�*���"��-s)V �.#�Fe�iV��$�L2ܳ-mKkJ���LhʢPUF�j[ieq�ZUp̸R����[n#B�+TUT�mm4(Ĩ���Z�Z&[�V�3kF(�W2��T̵E+R6ְ��s2��*�Ķ���5U��s&6�TY�ff"ȵ�j�Vթkr�X��DeW0��[�L��(�T�ڭj�l���E�k�q����ѹ\��V\�ɖъ[T�ʕ[ec��ƶ��Dq�JQ�2��Ȫ�KcL��#Q-U�AR���U""��Ԣ�6Yna�fU\3婡F�B��}1��啪s��cg��ų;AEѮTq������L�Û7�N�����2ãL^���\$(5ē�Xx.g�̉9ɸ��˧��ך�x�\��n2'Mj�
�����h@�T)�8.�ǲ:�q8m4q#�>��Z�����j&�(�'ōg'T�Z��J�g�h^�T�2A��Ʀ��ܚ^��t�P�v&�8�jNN�r0�J:S ���b��}R�G��onz���UoZ�bX�R�u@(7"�ХJ&��q���t�S��VBx_���Q:�����3�����H�+n��*`��Xt5G¹�_b>�C�o=~f��'��ꑅ��&]{�gy��:�s���ƻ����A����cΖ��7���#��
�emJI,�15`�)Ŵ�tZ���]w�B��oǃw�&�[�aBP���f:u`�����O#b$��q�V//�ӛ��˨J΄z�/ԗP��yU ����h�\)�K��勻0�-"T�S
j˱W�61���n5��C�P�u��:X�1p4s�Nn7x�5k��N�|���U�ܒ���Z�^o�L]�gQ5�x�(�s��f�����6���/6�˚솧�7�pȘ�eB��V�j��'7[	�t!�HF�e	�)>g�:�&� �wIc���,�p�%k ǯ$T�RLkSjiA��N�jm��E�w5�������s|]�*4𹯸����,�p��RL�$���\�|Ѿ|-P��G�����[+ӻ9�?i����k��)X�(x}�l�.��hV*���le�cĤ�������ve<�u	���t}��F�8;�������C�/���b�rϥ�nR�J�5�oc:RTa���&4�U��V><M��T��9�V���k���/��a�� d�w��c�~y�k:3ɕ�U�4e�fj��+�UK�~<��d��>�=`��(��e�5jz1��mV�&�`g��p�A����Ԯ��źl���<��]�H�Z9��6}^�DE�,3J���r�i�NV�XƝ�	��5�)�ѶMn>i#�.'��������R���	��16'�����mΗZ��,�]E�n���^=�l��929�c�;ا�^���&&Rjj�PQ���İ�y�ڿ{@?�Q��a�ADVO[�78�x��pL[t�i�p�����P���|�@���չ�U�)AF�rK���Pa���Sx%�����)���4/dX�J$E�	P��EL9Q]��"wb���z�ڸ/�$��ڄ��RR�B�&�<���};V�'��z�Ӌ5�b4�1Vy坉���El��B��@�O#9�S��͇���`U2�7��f�t��n�\��yi(�V$�d��848䧰�
WZ����`f5[Ũ�]��Нp�G�.tO&$%3���#�����r]*pa�=͂�^��;. �%D¨�����ڡ���:��Nj ��:�v#�۝�L���)���}.	q��D���t	�W��v�&�☟d	�3
L_���:�seФ#����Φ��af�;T)�8m��|��X������]X4�0�U�W��,K��?%��Sj���V��v^Ax�Zs�8��j��{~s��3�S
��7�x�u�ҮX��Jo�&���$�X�,S���zd	�Sٝ�W�JН��wQa�vtcU}5j���J��M͊��k�����o�Q�Z�<�to��:�!<A�0��ݼ��;=����xPr�BVW�a�z��	�@� E?mu��3(��=�z滳���G*C�J�xw��Cc�������۾��/L��xk�T�絋6`ڝ�yun�f��=�V�o��[t�
�e�j{"�kk8�EI����vb���Hx�{Mx:X�Q�˅:���q�p�f)��ₘ<G	�ʼ�k!%h�uϹ�`�]x�2E,��:�;�u @y{�cͮ�l�o
N�2�%|\��c
�=�-h]5�0�p!k�4B��[	gQm���c�]�c����҄�B]NԵ��\�c 9��0k�������uw���F;q���<�)Q�B���:gT�UF�Vbb�N�|�z�ƫ�Nz��D	�����Ad;䱄Q�Er3ad�%ˈ�s`k1`�m��pHG�$t�x�b�J�r�W�@��:;���F��X�cm�P�-_��ĨHKS0l{]�����VP��^|��l��_��De7����DMP�,R�E�N�k\��f�+X���w�*��į(J�l��ǌ]`��z�Je!u�T90���e����@�k�=�����S���>}�;��#��륝�)qG(K��$P"�J���r����fҌ�r�y*.B�2"K�ss�[*��ƕu��t{qFʭ6�@�P�M6�X����H}}j*0�:�J�.5ƭE(\��e0�LY�	�QbZ�Ü%Ъ�Q��Wą�]%�<���^����zv�K�B2|��Μ�6�Z�,Io���ʡ��S�Gkƕ�԰S˻X</��P	E�D�l�s݆�@�^HĢ͆1Ӊ�r��^ٞ�VR�3�S8�T_O�ڬ(�6�6��,���/Zް�����eom4KR�7������LW�N1tlV�zh^�|E�8�,gT���'u�P�(���f�9^�;H�5��vը5ك8PܕΑ&'���ڭl.LY:�ڛR��R�fIEY�^̴��h8g!@���nLCgo�XN�N9v�7�I�s���m#�bb��x��ݡ��X�rCϪy�om���b	�"��1�q,�m�uǒ[���7�KÕƦO�������-Z�>��>���x��7{��kdlC�-��Փ�'j1Ȥ�Zs�hn�����
U�bmţH{ї���ciߴ�cR}�":��~�v`-�5��F�ל�'�ޫ�|��B�q�U
�V�R�������2�ʼp�3�%-R��zoϪ�U��Mct�Md�W��Y�|��K�&`�Ҭg�N�8���M��͒��X��;DFBte8P,�Z����k�X�	v�F�1jp��+sլC�;׳�ܙGg.��D�M/Q�2��)�R�y�����@�-�t���(֯)�3gx��p�9��<��
3k� ���J`t����t�Qv#��P�;fZ���N��/g:��jG
��v�78�l��6�S� �Q^�S��9��u�� �j�=޾Kر�ѧ���^�(F�g8XT<cU%].�zM�t��}�u$估ÕmY�����f��e�j7�ܽr�݊�d�8o�y�\*�[;�\�����m����h�8���K�3|2a����Ɏ�z��Rm�"�7�V0�U�ъNV�;p��d�t�x�n�D��n$E�	�+�DGN�������s2R�9���D���
��W1����?	>����*��h��<�G6-nP�8&�5�&ycM�]'����*cf��V0��7����;�p*cu�����$Td�%W<�8إ
����&�,!YD�(�|��:x��ׅ���^9��}A�p�M���JrePCf��/�Ƿ�'A��]�Z��½ZE�Z�#IάK~>�1�`��N��s�Ӟ0�]��=K>:�]{�{
z����C�7HՇѻwo�hجޘ�9�ѥ���r9��goc�w����ph�PCL���V�ˊ�w�&�+Ѓ������Q�����v� ��<;��k:0&VMVtє:L�xX�c��O��lc�g�{Z^#c�ed�f��5nA�!��mV��``v��:�vz4�f�S����2[�+k�o�����v*�O�v����5j�<�c�A�NVb�<O� u�=>�`+��r�ݸ~�̬XT�lbJ�3`';7h٦���7�������-5�6�O�l��>��¡u�Qkؤ�;1ܬ�n�����-�(�cn�q,�i�\�ҐM���_Q�ݩS9>GX+\���a�(�y�|sn��8�a�Z^��W�4���j�a��j~�^��,�R���	���������rͻ����s�U����1�-`5�d&�[�;ا�5�e��.iW�o�6�g�նթǬ����E��&���3'��ʎ�}ba7O&�������b۱|��x�Afg{�}[%��RBr��ˣ��ڗ
��v`�	���xн��6^U�Ҳ^ϱLF�Ѫ��%�<\��6�~���#c*
	�},�D|4{iz卿y̢��>X�֤�K�|'g���}N��i;��u1|�̶��
�<��aОz�K��\?y���yG�Q���(4�V;+/�uZ�}��Dqʚ�T�S��s���gw�\6.힨��S���J�U�a��� ߕ-�^]P��Y릠�~~:�uh̯C�;3�x�D�P:�Hm��+�� ��O��T��+�cƛ�U�������![UÌ�:&��ZE�HF���丼׈K�������эU�Ր����ܰ��;B��+'ti'	�U�&�Z�E�3HDU�@QK�/q-�cRkR�W�&��"T#gN�f�-�-����i��̴�Ż�Q�{�Jh�۷-�͔��yD��YP�R4 �0ܗ	�����I�½�p-7�3�l��*�RȐ���Y �Т��o׆�'��0����<~Qҽ�~՚T��:�5��=�A��Wi
A1��L�ў�ۛ�N�F��T�!)0)0��F6lt(o�c�s�/�$�X��j�M)G_TZ�=4�h;
�2���B���%����l-�=�D;��l
�+�b�ԓ��+��i��������\8^~׷��t�j�O��4�t,���,b��8��:gT�
������X��lI�/jV�';˱�|���HW>>I��YUe�3X�l���:�P$6�``A�"GL��c@�Bu8#��d
gf�W�Om�c�DЛ�r���`�ү3)�0a����`n�eH�����'/G'�\��pwWL�o׼�s4k\���l½Ǟ6����.MD�݃��%+<���W�$A���aʅ���o�݌R�Q�2��:P2��yEN��K��Sl���h�ܬ��N�hN}=�p93w��|:'��������+1.݇��X�4�߭e
�aާh3[n�
�6��G���;F�ݤyj�le��/����dJ��@�{*�1��u���c�D�{�Vl6�W�v�9ZV��x����fҗX�#x<�g�j}Z�M�OP��僓��+F�r��#2�*�3W{��.K����`޽��huˤwl��a��

�Ț#mE���X$ _Z��"v;G�Y��О�D\�DA�O��b��t\������;�I�?�|eR/ƸbZwWt�K��L�~��,��ޓ�id��DSm����{a���k=���l�]t;��z{�3�!��t �rU��t͊_T��A|g�J�L{�n���.&]l-_�f"����C}��n{7۳��-�z}H�*#<\<*����go�'KdIZ����8Vi���)ᙕp�^ؘ�5葢�m�C��֫�s�w������LC�v#-�Y�	��^��;)�@��Rtfx��J���\Z��}m`}.)�q_OM��y����I�q�5x�3N-���N��Zs�77�\}^�[E)��o��b��վ�u-*6�0�,Q�n��5���F�v���N��7U�n�*q�W°U�W>�9��6���Kw�'��6�Y��iT�k��k (��W��8�o��]/f`�Ҩ'c������˕e�k�i�r��ڗ��y�?�՛t�E�3R�6�0b�oO�{�'}�@��>�j��Z��EO\��oN�޳#�&NnfE�9R��9 ��c�
���ⓢs�E��u�G�r����u^�s3+-i�ν+���&�MNc!��\$\�蟸W�!A�B-*r��gjԜ���e?VK���(��ȡq^�Qq�,T�ԷN��h�14�F���Nj��]L����˅J~S1`��P� _��S�r�CQ�q��ojsU�Y�."��j��q?`�ಆk��l^�ZQG7����7��No0S�>���+��WL�����O�����.��@�]ӝ.%P��_=�L�"�<�N9ė%'n��]�9ほ���H�AК
�t�Ն��w>ٴQDX�����%<���¸<�ЏC�]��"]BO��P�#%��i�t\�\���) �%�vo�6��LF��ӱXhZ��8ۍr	���ʋ	�.�a�S��Tb�;�G�$x(�g�����qun����M�צ���s�,�bN�qn�ki�\lƴF��5��R���J�H���W��j�:��Y7��&��u����jDA~n�n�H1�k``}W�W��ɟ(����5a���{�3׫�
^��ۗu��wm^_V��^��Z�Й~�8��c5�$XF�윷�/p���,�HНW�FJ{��v����Q5���	�������y��V	���BXM�����:p|��5���o�=�d�!�]�)`V�R�m�Y��;_/���T���Ჺӧ#Ϭv[��2��Y�����F��KG������B5o^0�(+l_���X�rgq'泰�D;z�������6���J���O��"u:��Ҍ��۰uV7�����j;vc���5d?�t�����)��ÚNN���޸y�����r�a���.�1�!�g	���!� �X!��˳2�r���Z���G�^U�lqV��cV)n-��a���[�tz]�7NN��ZL��	5;mό���.�/BDMX�V�a&i��\h� 4���t-�\�ǥm�5��(�O����q����)��-ە�p%���L�]��컣t3erW�M$yP��gU���{y�lVD���-� 6��퇑XAN�[0@��vwԵ�h��j]Z�����v�$@�ѬO�����=x���̡���5�W��X�/�sj�^RU���ү�ݦ�:��v�a�Z�޻���p�z��jƠl+��+;*��eL�y�'���	ɚU_d��ī76�[,�q�ӆY�mE9hh�Xg`�t�\���H��k�*[v����F��o�L���6���3���QKT���$
'��5V��<uat6�J��\�:�<�x�����Vmk���DcG��D��\�ĵt;G����o���;�� :K�޲-��B�(^�J���΅`��ncB��jJi���������n��2�j]�����!��rխ.�)���gLu��ZH�a�����j^^���DY���굟.�Qbܼ��Y#��GW6h�P��G���7w�-l.�ouY��N�����m��o�@�5s��H.��z�W�1|��h��7��ް�p�/gW7N��mu: \���|iv�fv�ZL�nb��.�bj�v霹��)�b����ذ��ȇvY��9�qQ	T�w�Vn�X�z��p���lԓ]	Ҧ��Itd��jM7�1�#��G[���r�J�|�������Wv�j�M�+���y;��� ��Y3�6��0��ښ�:�5u��Z̵:^�M�N<]t��E�����{�\��Gn�"�AǱqT�N�X�51{,ec�$��%�S{��8���D�D�8���+\s�H|�Vm<�]qXn��Ӕ�B�C�F�ss��J���~���a�E�:&b����n*;yv)dY���wWz����B0�;�& �	��{y܊��^��.���cT�A1K;�'��t�f���8�jj	Ӄyuι��:袊����$��&l���P�3�Ç�ߵ��\R㘋*���aE�5-J�TDF�a�[m�U���Z�Dp�����KZ�mmmQ��."2�q��ڸ�%Xڵikckj�(�أ��q��2���������s2ەJ�a�֥��f��UkL��W��,̨�[��Q��cme��C-e3&S0�J�P�\-ƴD���*f%�f9as.��fS�VU�b�\prٖ\��5��TF�\F�1��B��jԶV��U�&-1s�pR��)q�,jT�L0�-�kL˕q��ʍ��s0��ږゖ�r�*�q���Kq2e1Z�H�hZQU¬�ʭ(���m���\s+++ik"��Z�����ZR�1��fZ�	K����"��\��B�K[E�i*U��Kr�8�Z6��ʫ[-(��*�Sp(R����n5Ti��LL�6�֕U�[Q�R�*�RQ�U*�Dej���,R������s���}2p��x�J���xS��L���qA��z����K!�<�98,Ѽ����ۉAW��I8K��W&\��ERKx� ������pJ�gk"��MZ��X���Κ�"�h�m��)�,u1]����D\�<�wꊹ$I��ڦ����A�<�t`L�0�5zf���Πn��W�+����<���
*T�8,�V��=��(STSw�1ڷ����k��3��KW$�ޫ���׬`UC�T�!�paX�V�q�.�.RŌv���sǧ�����$��r*[����Tݣx��Uu檋堺9���:z];8ō1�����-%��y%��-^�3 �n�9�N�)��i��&.�'.���R�3�0
UރWCp���:BM�7�X�7���ҭ�a�jz<lk8&�sL���������/+*�γ��S\L�F:�.�a�h57���Sy�v`�w@н�~�J$E�%G^�Fs����y���o��=D�Ң��cQ��(����r]*pa���-�蚌��TFn�ƈ�Ď[m�' bjVK	Ӽj%�{_%���XLV�}a���.�ۋޠo��ʔ�;�${��e�mN8::N�t=���:ax��m�t�:�|5Ħ�p�3�Pf�S���[foU�I������3�ؗ%��y��A�y�$'>�����$n�2[I+=�p��g����#�f�����hn5ǵ�Wc������>k%T>�Ր��)�ޘ4���cC�T�:O��,}3G�x`�W唅��Y/cWVS�u��	��6JVy�N��>���F�g�SP[������	�%}Ői^�m^9]L1~n�TX	�}r���p5��\9`U/lٿ{O��}���x�����ߌ,��cd䘼׈KН��n�/��ɂ_��4�ʙ7�~Aw����9#p��z��,�j������{��;��2lmm�gMb�jan�6oX��R*��jp۝���b���z��vx������,v[]EI;��Κ��[�V;M�T2���J	tKE��)�$����km��+&����ѕ�oD���S�;HX�U�%7̱&EGF��]Qģ|R&-ani��-�M7q���F(v���7Hpy��Q��T��/Q�E�a>rv�h���Ż�`�k'edtO�G0��}	�����oxI#�ĆVEj�Os��Zc9�	|el)դ f��w���3�g�,w�r���-��-�]��:�dA[�AEC���[f�vHB^��7�چ�uί.�Wu����#���o5�{�7� yR�%$�����Y\�{�)��D}���	��sPu��mܼ�;�&�aǅYw���֖=�t%��^zJ��Q]�^d��d�}����T;,�۝R��i�T�&�E����Ƅ���U��dq)/����U�6��Z�*��E�{��'q�j�F'�����H�P3z��kM�˯:.��.Գ�m��Ŷ�ߥ�x!���N �|F��մ��gV3�`��JM�E!,cd�P���"�0з�C��Φ�Q#���GD�㽛�ƭ�0�^��Ȼբ�<�qx���1m������&����x��h#���&��g�Hu��`Mb3{��{c5����6�{}��GvFE3V�Ζ�*�*�5^#\n���C1m��gIA��B���E�Y�t��/�wZU�>Κ����G�gv��������D"d�u;={�xX�H)�m��ಸ8_�T�":-ҋ�
�R4.�LVpW$��+|�	/�E�5�%�p��_a6�-X�Y� �X��_`�bi9��=0��j���^�Wt�#M1��w�C����dq8�9v$3�#%���7�T�퀯�9�Y��=���	�o+iY�w��Z�Ђ���k5$��-��;o;x�;t�ho:N��hK��C�u��W�e��ȋG��R�4�GSo@馳��<v��:uj��qti�K�Q��{�Ţ�s�.�6K�*xi�ޙ��s���Y�K\v�w+2�oS�I�s�H�#q��!"Ҋ����o=��XR��J�	���qk�<�L��W�q�A�t�ų��)ȵ3�Ԥ�¹�9�Ʀ���+�M�W+�ϧ���^��V�zqh�mǰ�����GR,k��4���v�j�w���� ��g��j.&����o��L�+��^PY-++��ߥ�8ވ�i��ˢξc���0O�[�����j��¡_r�\SWr�ǀC�
����M�1^d�	/Ե�̴6��p1�򰾬Ӈ��+5��꺱j%���1��.�}D�ˤ��5[���Cި�=�i�H@v=/�(8��Y+0����p]�����϶ɝ��M����l %�8�[K-4�����9\�� �#{���B�H+5���nhY�W�����>��Lbp���P�K�;�1��x�g��.��_mr[Wȯ_�)jN)�Ns5���,n��;��K�:���mpet��V�������FY>��v��^'�|ع�]��g���4��i�`�[K����������5��������u����J��㷝h#�ó�kh�K7�Κ�e�u)��QRg��[����\���WI����9[x��t��|��9�{u	����"k.ڊԙK!�(!F�����4�xAa��i3i�L�Bk7,����Ռ�EI��i�+�P��!��B�VeJ��bZ �2��G�중���X-x���#C�� ͊P�M��2]V8d�l�+�7���z����ĳŋ65�6X�<�68h�%֗��#ڬw��LVI���U��(��y�.�&n�p[i�LhNb��xa��7&yW�5�͒�خ��[��w<1����(�V�ё<��
�7[�f��z)=��Ѧ�kE�1�<�	I'SV��:����a��C$��nD������g|�N��I�����rl6�Xz����gj�ʸ�y��) A�T�Iwq̬�8��J��6�j���q(�a��#j����9:�I�rWꮩ�w��VAgK*�d/p渉��,�Ow����bZ=�%T$sv(��;�ॾC�/��=�"^�(�3�pn	%n�w�A�
��B���h��Aͯf�Bw,�0�n)���ޒ⚮!��Q8�ж��3�N�+�OTފ��S22����\�9�ir(FK-��<�p�y�)���j�o��h���i�����-��glrK��u�*1�i�{��`�b�ni���U�\n8V'�� gZ=�(�}%!�'���K��A,3�K�Fٵ�j��B��Y�ǂ{�$z�i���4R�8�`��M��3���z��c4�;"\Df]��2bgb����;Z�Zt��Mg�1�Q�e�譺t_N�)�ێ�ͳc�fy�`�"�C��9�t޽%^x�	�r뒀M;�,٩a��e��z������NHHh�5ڙ���&��j�,gC�`�V*�fP�Pk
�㥶�)FN��E$D����?FVl��S��V�T��8���Y��n*¨��/p���,��i۝;�h��oD�hN��!bYV�TI[���ש���\��+zi��1n�i�ӈ�='���BC`�x��:	��{N�]�40ʊ�&N�m6�b޳��<N����z�c�]޽����8�DO���|\��l�X� �J��7���Ҝ57=zct�e��1�{�J	]S�$���V.Ʈ�*��o�rL�R7y��4��qGV�E��&�r/�%�0G�]^ݎ%p�i;��)��g�u%#kz�郗ͻ��(CV#��@�꺳��D��q���4���X�DIt�ȼZ-��K8�x"�pq�j�5ڮ�c�N��L�ܠ��V T+y�)MP�����+�I
${GH���
2�]J�eH�g5�[8�r��l�=>@���J"�!J��ʌX�Vl؎�qf�c�aA��7ji]��;�I�!��!}�����n^>�`b�]��@6RCOd=2���(u�C2�I5�}xY�l��J�E��p	�R,i�.�z�K��
f���x8�xqL_�R�Û���U3��:zu����$԰����5�M�ŷ��_u6/�m�h�;�_��6����2�.�o�\�s�k�;��ތŶ3o�e�^&�t�Z\<��~P�Z���\�3¼���׆�5�Xi��x�ڎ�׊�Ӫ�Y���i o�U�v{��
�4?:�5�a�zi0�c1|u��*��=�(#����|�燺{��Q���(�ͯ�H-���d⏮�]������%�3��i��u6�t�Y�k��t��'���H���coj\��x���r�}[++��Z�·!j��)]���{�]��8���MJ�8#�|Gl ��-(�jNR�C�9v�o���0�k�[]@y5o������x#�|}Ƅ���:����x�l�iI�}��g�o��|,�R�X ln[�t|�
u�P2x�czya�2�V7�W-p-�摼#"�d��-5���9N8����8�}���d��#p�y�z��Wi��9-����E��dݘ�c݈͜^��,�Åݒ[J�H�����oET��O��k961+����5!�~�M_Yb꣫���)!3�w'�q���ʧ��4`^�z�T��O�1���u1>�i;8==vy%���V�`�Eg(,���f���z"���-��Kf�y���b��^�E���7��W���	��hc�� �7u��!�����nT���>�TIմ6ۜ�د8�eĽ��Ư�
�ث[��U�/�tj��ls��9/���^�JR�I�9��IW�q��{��֠q-�����2�5{7��U�5F�}Y��a�W�v�\�m�m�{�~/X��[�;x��j�čkƽ�aB\�(xߤ�Ќ�~�x>a�X}�E�Ѱͭ�of�\ve�:��Gv=��+���&0S�<�୪I����T��I�\�-��E^�}���!�s�[��U����ob(]��@\a����}�S�2A�lm��t8��8��en&n��c�-Zt�%urͻ�=[T�`�үcZ�at,jYۉZ�5T�Q���-aw
�xQ�ŷ�9c�����s��:L�:�$�$���Q��v�`iR����wa��וTW��Bv��(��k=���k<�ǉ7^>d���9(����+��$ef�H��BCt'P�l��Jmu�����S3�ӗ��ۼ�%�免b����K^9;=��ےf�HZ0�;�*Vv0��w'�v�cU�y�,Q:��x���GD��ДC;z*�5���:��\�/I� ��];��M+���޳�m�����n�v�Mi�e��I�N2�>�8�ThIW~�q+Ư�Ue�l'ڳÝ��NU\O-�w���ݩ��`0�^ӒWU�'Uߣ�Y�AgPh���<�Qvt#�}&�F�4Vz��(�!��sv>�Wq�����ΞQQ��ق����(�G�>�S�iU4B��4ue"�θ�e��躩�\��6�QԵD�i��41�b7�Mx�U��M=R<\�s�|�p>��/��f�U,�Mk�.\��ŗ%�ru��z����c0s[J��φ�k��Ug�f�GuU�J����j�e�G/�<��hC3��ZtR�(L\]=M���z�8�Ri���ZUz,m���S�7��\:=�QS�.<R��';}F��(�%�C�ڙ�}\\��]��P��`ԭf�C���^���z�U˥֞�iS�@�g����y�ޠ2���)��Xu��v��mD)-�e��a#����Y[�m�.��hZV�����6`�F��-A��ـv�[�(�sv:J��ﻞ�(^0�d��F[���)����@�Q�5�8��nl�Յ�e���+6�%>�@���$i�����Wf���|��$iKN��D�;�;8#YWV��¢sfK���3q;�[���7�E�B[�����l���g%B�w9�;umKwyfZ�k_Cޡ�Yϥb �C�O�]4j9=�ozf�6 !�S�*�m�L��2�	���;���Q��H�V��+@��z�,qV�㇑O��CYF�,Z���*[�a퍫��u	҆N�*1{�R�sjp��Tެ��{yO��oU���1�&~GWB�������]p�#�(�Lp��j�y�R�0I�Fbմ�$�#�4,�:�>�\"�i�2�ݺ�f*tu%#[$���I���Yث��Hq�
��&���뱗ni5��e�U���{ܑ��(t�k�4�kt���2k�ά{�/k%7vK��l�ד�	��n�izX���ٴw7j�����A^E"��8P\4���Cp�L�w����:$w���--�v�\��K�' �̝���i1����fb��d��U�t�f�3Mm��b�=b�M��,�hy|p|@:k[��!�VR��esǔ�h(/������p��"���pp���:��5�b���`2��t�d��*�8�a �?j��S���a��G+FF������}�V�	W�/����E�[HZ������F�W������:/Eiğs4��K�8��bѠw�#x��"����P����V���E7�cV�t��\��鮇�V�X���d�u����<�p6�v�Ð��۬'���ێ�i��H�@���H����g��#���Ӊv\Tֳ�Q��J:Coi��sBW|�hm+��ŻJ��02��o0K(J�w��>��X�h����d/[u��x�ܾ9���n>m'}��>j����5���^pvwzKOY�4���4o���<�>�䟤�cWm��ݙO]N�t��dI�$��]vͣg� �Ň�x�����\��>�f^�yQЖ-��nA�\x�^��+�7�Ƥ��M��\���%O�5�5��`�fv�g�TV�1��;��%�}Oo�D��9Q�]&]�\�|�Q��h��s�@x�/7XӔ钖��%T���4�H���r)�[}��������bQ(�S-D1(0L��*��1Dij-Q*��X��j4[B�4�*-�Kl�)j#YhT�m��)VҖ�U��s+�U�E��kh+JQ�*
�r���ƫ���Qb(��H�$X�JT�%r��Jڶ��֢��k2���ʈ�*kFҌ�b�K��i��q��E�j̹R���KJe�q�*��k�D��Ņ���(&�n+j%��KcZ��l*!E.Zf&(�YV�j�VմVљk���S�����*�KUU�bʊێ
cKcq.Tbʨ"J��nYDR�l�h�+mem�k��r)�"6��c�(�s2eA�D*�Z�K
�DZ�2�V�Q4)h��L������5���2�jcr��JPh�J��X�Z�[bVTUes0�fPQE1V���+Qj�Y)lD�Qr�E��PdYe�QQ�\A�EX��c��1k�1�����Y�b�0�e��U�T��ST�������`��Ra\wnj�@�A��M��]�C���v��g�x��R��b�݈��^+:"<̜���1��o������6�p�mM&Fյ{7Χ��ڕ3َ�I�aO�S=��� ��:K�{|Ŷ��m皾�j��Gn�cpf�i�><YPȺ�C5;��ծ�߰�`�,3�K�h���3Ϫ��l�/]=���y�Vn$h[^�J1��[U��F��S��"=�^O�w�����|՞�%ˋ7�G6$����N�yZ�e�vR���8M��7ݧ�H/��gv�&C�;��2���=�E:��3���Eçĳ�iQ�m:Gu6����)��n4�>RzNy�C�f���J�}�gx�}�-��|T�;i�m�Ż;������K6� ڞ�j,]2r2(�����7HM������F�Z�q0��Pf�SfL	�����S�ҪJU$k>�%��u�*/�Ev5t�Tf3#(�y���v�-BjU�&*Z�Pʲ����R	��0���`��'#��e�\��V���C�1t�+iq4��q}[�M]��Y<7���Lr�X��Ķ��h��[wv
�9�t;�u�<4mw��l`���7�s)�oq_�}�&�J�3��vS=ޖ��q+,�d]��zy̚�t��Ų��˹{���`bp( �Y#���廙z��Ὥ��_R��sܠ�g"�h������a��>����f��c�^�2�"\�]��g�*5�)MT4-���+��L��ɱqg+eN�ZB��&����19��W�^<�qL[jh&�����1�3�p��H�$�+�U4��#]Mcx+71f�׊���{:�w<��M�����o����T�S�jm�b��o�k��b��M�e�G�%�����7�^Q�M{ư���:v��[�����u���{�!��xAߞ�x�n�k�٫����&1�H�8����{���E�ӓ�e�9��<�����i۝;�Γ�oC�qS|�ڄ�ڝ�m5�қ]]g^sc_N��5��7L�. [nr�-��#(徠B���ݫ;CXM<�����.��3E#��I�X�n"v,�6�*-��wXet�k�����&ErEd��T�V���M�ӹ�h�=4T�,��Ԅ��4��$�~�Z��+q��Idu6��4�5m;NÝ:�ȡ�me>�Kkw�$���P���BE��ʞM������6�n�:r��2Ԅ���F	���)�7+���Β�zbg��V4�Z�����Gyx�����f��X��� ��J̼�,����"���";?kį-�*�&��Ь1��
��>Oj�� ٭�(��Kwԟ#(�u1KF��-����;O�s���
-g��b.�����(�H�%%�"ɺ"�X�Q�p�-���9��F��r��b.HP�4�A�h�7�2$!��v���5}��*�P��Wb�B�ڨɡ2GLR�-��j��pV#T��'��4ue�[sV{'��D�Ƕ_��X���o��)�E!�9��u5�W�����1Nt�r�,�޺��	����@7W�s�$#��:��#m<���m�(��լ���2���^+�����k�
&IiG�p�3��>F���6������}�,���^��XU��㡛������4����٪�g.E{F�	R��"z���2v�D�t�wG�{���m��6�����s@pu@�T�wT���o3jꊙz�J{����zv�m�y܃�^�~iu��v�>���n4-���D]4�jێ��X�Vsս@f-���g|K�R��f�os��/�ꢗ��/g,��Ii(c��Q�:m�΋���l��*my��n�!�2;y�	��i*Onc	�Iގ����^�������,7�-V���&;�To�]�Z���;&;�.���Mڐ�	�-��iM���.z��
��^��Z&-f�4�b��4�:Z��]�mzBؤ6ٗ�8�h�Xm�ޢQa��l�x9�Y�ś�`�mc���Ѥpz:a>[t��)�V��-_��G���q\��~Ʈ��h�����u��mܹ�����g��mާ�*y��KX��Z�ĬG��J��6�jll�]G:7q�*x��)�ʣ78,�A�}z[�M�Ha�.|R�ţ٬�h��Ƭep�����M&ILj��X9�|&��aY�X��R(��ǰ�x����`��-K$��@7���D�M��v�ѻ���!r�o���/7/fM<�b�ī/G�8ĮI���?K�^>3~�ʺ��:��s+��������h�>�Ѿ�c�w�D߱8Q(j���2/U�w7�È�P���z5�fV�}m�7
�y5w-`x<^T׈Q<�4u`��
�{bq��x����7Ť�\�o;(V���N941���+�M��B�D�udM��98�-�)�D����^�sW����h�mM&Fյ�9{q����Ծ�`��P�%.�
&�k�6��{c5��A���m��캩��kj�w5���*�w�Uקv�
�Y�o��ÿ�Q#gU��R��ԑ�ޓ��Q����x魕8�emU�gj���U8���y��"ߊ�8�o��g:j�͉!��Ӵ�
՜5������Lw,�H�$���M�A�v��mt���hLs�&�:^�Bzӣk@���zT��9o����5����4I�oyK��0����v��^UݙA��ǨT޿K��װ��<6-tOtų�`����gv���(��1�*����a��+�u�XlWr��u�8���ؔbˮ�ݚʕ;7U��9�"+�}�QDZ���a�����z:i���i�nt�Ф��bĻ�LU�R��A�ڵ_6J�/��Ɋ�M���SK�Ż�����<�a�oN�]��H�\����9Ж�LH���|\�;���<��H�I]�$5�#�Q�Ź���N���>㒂S.
��%`]�^)����D���Sُ[R:���n�}
Ƴ�x�Ȱ���ƽ!�b��	n�>12j�U���b=Oy�:ֱ�;m,��]��9��d^'�P��9��C��1M�����+M1J�Po��x��"Y���4�PA�{گ!�;��{�C��5�e��6y�T+y�)�dS~��9(�UXTOvJ8a�6�5-���h��Y�1���W��e�1m��Xlֹ�M�]�w�}B�ì��*�:#V��o=Y������^w[ck��݁<f�+S�~��wuG&T����SN9��wTy�CWV{����^�O]���WVo��GF��;���U��yf���AU��F�C����_4o�;oy9���j��ת�)q�IW%�bt��v�7��S^'�,�|�͇����.�6<_��3�뷂��+ �MueM�=�iK�)J�;�Zk��������O�-���wm:l����ɋ��I׼Ua����;z����{�G�,��x�HC���/D�����$ķ{���.��6PG �m�|�L��N���$��Z)o,�-��(���Ĭ��'���i!��]4�sX��{S2κn�a���RR��i�/���}C��!�(S,�4�ƛM�hʵ�L��C#^S�ȳJ0-a�S���;+#�@#��(3(e��S�j��K`��Ru#V��X�x���Pu�D9{/=�aH�wf��v.Z�Bj/�]mZ���X�V�Z�ͥRT!{�n�������1Y������%����Vyh��[�i���{6187�G:Jn��lb;&�*&Vu,9�]�m�w�56���rX5p����=F*w\�Į�a�oh�̎e�Z�,�n��5]$)ad�F�V�:}�S9�1!}Fܘ�S�u��j�& z�մH��U�/[}�4��況Bb�d�J�}C�����[JE�9���sť�m��K8HER�U���r�w�\hGf@�����h�����)˜���rBs��c��$�bN�@؍T���hꑺ-��=���]g��|n[񰧽$[-D$�G�QԦ�>�Y<�t�TF��z�Vk4�z����Jz���ȡ,x���ܭ</����{�j�����s^����lk�vRxv
K��u�,���m�y܃���.����y��ՃqR����9�fB�5�P�u$8����۝7o/�̖ܥ�&���[�I�ȗ�pd�Q7ԦaA-�=w4�Ġv��Q����l�r��:yµ]r���yN����,�:�t���M�J�;Mࢫ�i��M�ηڬ.n���s���Jp1s�{��Ν�#+7�hvԆ�ueH�^ұ��Ϯ�*��`��4��V,:c�T'�0T���UF����5�\q\��?�Lͥ����-��~�9gI����F��^��<v�:��3��!��{�p�d	��˖�,�p����[�b�]�#����n�a��ήa�Ta>�e���<}��O7�W1n�i���N�b14;jB����H"��[�v�}�46\U�3`���'���56�ǎ^��GEu�꧹K�]�]��{���pb��Q����ڲ-�ƓIx��oY�ؾ�/����E�E�>��&jKd/s��Uu	j�G�#�^[%V[$��ݮ�ɩ����r�GV�U��f��@����ꮍU�9������3��Ev��	��GJ�e[ͻ�8��
$!�7 ��􌗁R�ð��=�A����}��;8�����SD(��IĻp@o;�cʭ��:��y@-�M6��S#�S8�	�� ��(s����m>+�H��qZ@�!�9
R�d�5=���*['R�+~��U��c���L:��K�������Guћ���H���{��^OP~m͓$a{���o'��B��(�W]�t[�z+
d�F��hwo'l�E�I�B�+,�R��N�Kܝ[晡U�
"f�Z6nȋ�1<mt^�4z&�,�ƍbX�1B�얝�����}���֙!���;��o �����6IL���Ƞ�ɋ3-�������	ݵ��׳�l�,9�ǭ�X�����iz�)���&ѵ�����q#C��J���@]6an�T��q3�۞ݵ����!z�L+U�����YΚ�3bH{Z)P��f�"�=�K�xQҡS�����kv��Ӱ�N��ѕ��4ˡr\Pb��˭v������H\�W���GSozi��-�M;t�Ф�����y�T�v�n4�.���P�b��@�ރ6��[�f;[#1hG�����)Y4�R�H�#L ��bm(߹?g2#��y��麪�t�Z�Q�V5��r�:O�Ԡ���%E�T	�O�y�F�wj5�u�D�N�6}
���J�r
|�ƽ!�u]t-*�Wi&�]z�B7����p�����[.��n�E�p( �P� >0�ToE����[x2|I���ґ�a���_ct�rᒋ�-�\3&�Aom�Q�Du���,rp}�:�y��r
��� �ذ%�ZT���wjC�T�c&9``�r��Ot�����a���Uh�So�y}��i����0",��4-���v�#nںF�}7���V�1�b�q�]G6�jY|o����_v�n��=� �3i�j�[g�����9�X��vd�v�+��r@�̦yP�����o[k��Fc��u��v=r�u��~���jMC}s�©�����ihu���Iܮ��-�5)�*�}��P��-�4�S!M����0��;��������Ve
-^�+M9�nvi��ZB�ZA=G�$����۠4[̺�Eۂ嫧���
֑���k�U�Z�uأ�q�-�{p��4s�kE-�\#6�/��vq �9�e%b�-�7\��ۉ�Dx[���l���Zml�o����h�
�htwP	�H��N|&u:��v�,�J9(i���[|�z�:8�n���8r;3N"�=Z��'6�8ԽB�j�c]v��]�k���$K���x�,#4�TH�脆q]��ܻ,n]j0P���fk�(��:nZ���F��aפ�@^�P���7"��,�aO���T=�sf� �u�Zj	:Y[ej1�Yy����8С�ϖ�l�����u�DS��F��p�v��<�n�6+gi�wt��Q�*�U,�ut��[�9����'`P�;Sݬ�ȊSK%Kc �\;7���MR�l���l�ǣ�a䳭fS�|(#��F�}�@qkl����|Sᖱ\Z��&��p'TM�e���,�B�*B�@&��e��(�|�ȱQ�wZ���*=��e��4�m��=q�i��MS9K��$���9-eu��9M�:Ɲ�e�ܠvgmY�r�%����
ԅc���Z<��襞�Ռ܋A5dQW�u�p����LS\^��<�Q�wr
F��V��^���-�g�6�hcu�)��
FV���i�ƒ!�̺G1�1'E�Y8����8�&7��AWXݼ�R�U۱�d���t��0)+�goTl�/2�-�-�]H�$��5��;��d���g�L5�$�ÎleKخ:}t*�.�O]K���ђ�6�[��.+}��|��u�U�$�2	o4�qNu���m��]�DY�ޣ�Ku��Wױ�o^�"���Equ��*�c)*[}Pv��Ⱥ�=I�f��وu�N���vv�i�m��{č]@XT��H��|��')�̪1�e��y;�v��qؕf^���R����Q�þ�+:��p�W��:ھ��4\)�;P���i:5Sءs�
*���b���\4� ��/���!���g%��������_����e�ʘ˩s�y�Gq�orͥёNjkC�}����x�_PW$��Z��d[�Ge����-GGS�+sU�sy}�am�̙� ��U
$֢�ӌF,0ZTq�9V��KmnR�����H��VīѥR�l�3*c\�KkU�ی���D�[V2Ҫc�e*�Um((�m-�(�hƢ�,JZ�%am�R�J,������Z��+TDm��Dm��mcrܪ���cR�5mlV�Ɖi��XU����U�,K-���U�T�,aU��[KZ��QE��U���m-Z��S-[lUR��-�iJ�
�˘�31���������K+j�kkQ��F�R����R�UT`��FT[Tj�b��Q��Tb������D�`ڡ*Um+me�-�Q(�֢-�k+im�֣mh��Eh�D���X���V[km�Uj�6�-kU�mmZ��ԤQUm��,�E�e��T��V%��UE�-�mJ[J"ƔU���6���Q��jʲ��(�m��kj�4 hD��77w��&����ڷ�z"'Z�*V;��Z�ͮ���E�Sw,��65R��!؆Z�+t�xsD�& &�!��r}�[S*�+��^Po�e[W`K8�i��Ì߭�x��:e7$��WR[�lה�)�Y���[�qH�M�>ɨ�y�m��+���IB3�_�1>5W����C���W�^<.)��v�$���K����_�A���S^:�5T�77�b����VT*r���h��(	o��=��Ư��]�8�BwmM�RN��DmT�Xŉ�D�I6U%̔�C�k�>����k����:k��W�5^���*�i�&�$N�e�]Ud��a�%�uS!���f��Κ��Y��,[m4x�UǒB�)���VҼ�g���m��o��Nn�):	Wt��RG��Zq P[DR���
��Tu6�t�X9�s�R%��2�J3MvKL���A�������lɤ-��)�4�m��j剘��Q�y���^�gN�}x�e��F8�ǹ�!s�!��g��W�E�wUr=H��@*����Cr_oB��I�JVd�tc���ۖ�[Е��5j���2���U�:ɴ��� K\t�ŗ@S����x�����W�u�|J]R�����%H��cP�cQI���J:$�ڐ�6)	��ݞV	Έ�|/oWs|Gj��ɼ�^��q8y,���0�1�t�v.��]r�K�<alwC�%�cW��r��^/�^���T�/^d�\���ZY�mqzZGڜ�*�Q�IWqĬ�GE���[�a>՞�{3���]��y�p�=����q� e{T+E��w��Vr��iYBڻu;�'f�3׽ǫj��)Օ[��'z&���A��n#�oT�sd�_r3���}��ti�)`ؾ�=OҐǞ��(S@�����hl�[sspv=
�T�1ˉDJ�l���72�؇Y7�u4U@�U4�Ļ��8r�b�x�[g�Aozj��4��|ņ��{�i���s�����+��k%����~ڙ����A�&��v}�h</���X}go<��k�=�S�+����!�9��lBV�ژ����B�:Cd+hf�d�Nu$���q=�*��x[A������i�/��B�T��@���ρy���,�k��y*|en�Z�
�-^싊2Q[uc����6��/�m<8i�����4c�$Ld�"�n9~�\y�;k+^c�mIa��X�*��k�ws��7���<�h�����������l�A�m�d�n�P��j�ֶ}8��g���P�.8�y[^�U	�nJ�a��H��tO\���r�%�QQ'�ki�ӛ�#+7�E����3s���%N�qT.N3��Z��l'Jl����\�2�k-x���bhv�Ȩ���Z�i嵷gx���m��|T��N�sƋO��6����D���eDl�=W��%�Ƅ	a�R�)E_7��5t��D�?t_	�E�t�=oM�ZUK	�����WU�%��J�q��-��ŜΙ��]{�B��#�Ǿq8��r�Ҥ�AY^��unԼ�/;A��, ������eWRK�,�e�`�]��8���AB��s{@�#��](�w�ʻ��V�
��ە�)f�𒊳u�9���-�am����!n�쫗�sS�!6�[SqՉ�U��θ+���S1�Wm7��Z����G&��;� �������Y�d�m�|اrr\ilk}�XyH�	��$R��yA�>��������(�h�x4)�n�A�����)�D.�A͗4,�<a�����4-���s*�p�J�a�\��)!����$��Y�19�yدl��mM&���a�w(�Gq\�%\�2�5@�7[�ͬŹ�ݑ�h<�+p�
�����-$o'�f[F�j��Ц��wmg�k�ŷ��C��b��em�����E�0��	#l��}{5��H����Q�����1��D�0dA}+M��X�Hl��4	�l;z�����q�3�5y�>!�{E,�5o���s,��9Ҟ�-b���.��l���i7My�n4�zJёNr�.i�u�"��`�BMbIW�4�z:�{�Mg1n�NÝ&j]s�����M��]�%=#+�5~��RP�b��Gm6b�C��������V�:���	� ����*cMYaGy�c���E��jc�����O�!���΋c���h v�xEv[��T������i��wa}O/�J�^���r���Aܒ�>"�E �!�OV�-jǼe�tD �Zq��=���-�x�jkD�r8H�類r���^:F�n��-(�|\�;��dNI�:Gg]j�m`پ��c��roͻ���>>�BPJe���X��Q:�	Q�{;�2;`kį-��-�~O�X�rlbW"����5� �h,��##�a=������/�U�i/���K+ �]��8�����R
�a]��_+��d������r,��ת��̼��g"�o��v��!���Ǵ���v�\n�jk�����oA[��)5u:�`���V�B�%�B���ʦ�
8j�&���э�^v+���h�UT�i�Ow4V���#4RÛ��SF=U�F:*��bN�%yiܽ�]c;7G�Y��j��s�o���.�x=�Gۄ��֛�bi���f���	Ͳ�{ۛD�%~;�Zk�>���}�5`�N���z0�]�"Է^�xu�A]f�V�V$z����Y�����;�*@x;��=q���5
֚�{\���ȩ/wG��7�3�MA�vv���n�T�)V����丮`0J�Y{v�ܹ�B�un�w�W5{�)9���`��mK�+l7�ͨ}�qZw�j�,; 귎�7K7�Κ힊����Q�=\T~��Ơڕ�p���;��A��|�������tk��L�R{sy�poD�k�R��n`��I��ĳ�Q�R��z�%��L�֩F����:�I�8D����BE��a�����Yu�����Y�о~R�@��/�ūYK-y���� ��fPǧH˭�j�ke�%w�l���,h������9{/=��=l�ќY0ZU7�k������m��@O8�_&�.Ư=o9Vy4���z�N%R����G�g3��=i
~�'RWU�%���V#����|��L����=QYJ��ŰRD�*���(�{UH殇H�Wq̬��-,L�S�fr[�=i�}���<^��N �X$v���]�O3�B��K��A���wh�GK;�����ޢY|�P�l�5���ʻ�Y���X,K��q\�*�Y������=�OՍC~Y�p<��ˬ�Ձ�i���3�*N<uջid�<h�����ѻy�_M���B]$jL֌�q��/Y:���*E#��p���vp&�Ĵ1���*��Q��GVP�ܝY*,�pg.�M�M"������qX��<����d߹�׈UDj�}��y'�fzD�"Ϻg���4��|�n^h�f�P�sǝl�i2�N�/�R�P�l�EZ������l���o�>���X�̫��v]�]��G��0�%�����wmg�k�Ƿ��gA,3�I�_l*�Op}Iv���7�De�sE(�KEmU�`����\6ul��Vg ��6���_���|�t���(J�;M�ܺzp�2���5Z��q��#i��M[A�v�N������4;k�ӷ����vj�/�E��R�0қ��bZ�)?&��K^'g��������v��=����0~�'�LU�Rv����,޳�X��M�l����&;j�6��o1�S��FZ�OP��^F�N��,����<x��¯n,&���pE�I�Ӯ��:�E|��g;��9ɁPV�ֶ ��ܩ�����U��}��L��q8'�%tyk{+r�b��P�"F�]��a*)E6�H�ԑ���R�3/���������?=OI?^�ii$��@�!��8@�i�M����C�/q�K	]WP���XƮ�%8���Þ����ґսT�+o��X+m��k���a���̿��lE�S��=GQDu-c�L�iee��^���D߱8����G7
�,�G�i�g�� ���ƒ�r�}�qM]�Z����E�k�(;TR�QFnaل�^�J�%��sXVz�M�{t����Bhc�x#'��f��L<�7q�xZ$Կ!�Dj�MyY��nk3�V���\Sڔ���y+1;��nRU�*�VK�x9�F����VmŶ3^;��AĊ�V�S������/Z�D0
饷�x��Ճq:P��N�u��!�֐��f��wIR�+8�+�a��I�}G-���Vn4=���8�qB�M�����F��M�m�7oL��:�339wq�+D="ۣK����իpef3~E�ѧ@[/9��C��b=�8���ѓ(C�t09B�gG6t�Ϫ��p㕤(I�&G�mٮ�j�va�Ki�Dx�\�x�tzĜkN�H�[�Q�;��j�a��[�;+�P�.9���u��6w}��wA⒞��˧�[K*Y�A:i�M��i۝;��2�8�����Q�X��|���U1J6P�,��Ku6�t�X9�w�Ӯ��b=��2US���R���O�_IF:�mzC`��/��m6b��c5=}�"�;gv����`Z�Am�x����� �5(3`S�J*������J1V�;D��Q���:�QYlZ�q0��Plk96w/=}Ƈ����+�n�HI�S����v�)
�e��v5y�d��l�O�^���T�^����g�7M�;#�S$�7��-����?3]���p���dX��S��-�>��v3Z)!#��E_��X�Y��9�@���{�Vb�cV2�l��k)q��#	�ՀPw�r�7�o9�#�w��vߔ}1zOU�y���E�Lޭ���7z��,�PJ�	.7�/�0A���[�����a��e�'H�N��	�w����RD�7�����'2�-���i��'�}0ɗD��խ���X/nq�]���X��@�ܱn��]%�����Bރ8'9+IWf�Iш�.��Q>᪽4�`�t{ټ�Fe-���6����qL�;���SI��!�O9�!�5W����{ l*�;N���-rHF��W����͹{]����.�GU�5�����%kP���F}�h�=�2ܯ:���w����S�bő�8���Ǖk���u$8�`����ڡm����V�N�j�q��*Vh+���]�0�HAmh�Bu���V2�(#����Ӡ�ӛj$%���%�-�F;sXK:NoE�E(�oEIW��-�Ɓ��pJ87���P9^�g;MƜJ;g�č�$6e���t�8�r�`�w��#�K��%��X1jƲ�K^ ���tI�!t
C{t���sٸ��L�f�W8���G©@��+�|���O>�l~��O��H@��	!I�	!I��$�	%�$ I?�	!I�IO��$ I?�	!I��$�	'�@�$��BH@�BB��$�	%�$ I<IO�BH@�RB����$�Є��$��$�	'�!$ I?�$�����)��;/����,�8(���1&m|����j�(EIU�Q(���T� "! R
T(�����R��%RU(�TT��*B�E$
Z5�QUHRH�(*����H �`ԊJJ%$*�U�Jm�%%"��U%I@�U�T�7���H�SZ�=5TK�S��&��*�E�)D*��dUTM`���Ԩ$�)UHIUU%Rc"B����TT�T
��D���S�   `�{�
�lKm:݊��r�+eٷp��ˣk�-��lZu�v�v�:;���u�̜�i�ۮ���J��L�;v�:�V���B��I	)�   X�������htҫP����]:�F�7T�ٺv��UV�*����A�)�i��Uu���ݩ�5�Ź�����Ӱ3N�Sl-ª.��%R� �V�   1��ַ���[u��9]�ݴ +�+We��M� t�m�6�+�fST���[�4�2�q(P��СB��7
(P�B�
��B�(P�B��JEQE@UJ ��2   GaB�
(P�C

 �B�
p�(P�B�
(7�P�(�
;���J՜8֜�ˡ����[:��+T4�wuS�m��[nq�����hn�R�I�EAU(�K�  0: ed� b�EP�[0
�A�jR�6k` ���V��2cE
���F ѡT%QHhd��P��J�  c�(m�(6�f�A%�� �֡@(�a���؀h�M�
5VUPv��@
�ʕ(+���BU��7� �"����
h, UX� ,` 
Z�*��0�0�!� � ��5����*�T�  7/)C@�@5��(��V��ݘ�-�kC�F;e�Mt��t�(t6�R�#l��'q.��v��"����]�7f�m(n�(��U�]��������  �����t��gU����R�wZ�WYІ����J҉� �ݲ��a�\��Á5������t�U#N�ʪi�sM���C��
T)TQJ
)"��A�  Ǵ��Qv8:�u����YV�J��4�4)v��Ý�Jj����]��wu��qѧR�k�lm+E 1����(YÎ��wwv׀O@2��   ��a%)(#�S�#$j  ���R�   S��`��� a i"&ʥM#0��SR�
�I�g��%���H��1!DG�Ѻl�$ڎ��}�:&"�����<��O���$�	'���HH�	!I��B����$��		�yϓ���?�O�'�J�K/2jv`$
�Վ�PUl�H�cz^���+F�{�0�7,��[k��'koY����ܷ�Lp�](T�f9W/3���jc̉L�b�Y�ּT�c�l2��4�[Щ���XXؖ�-�B��1���Yb�*.��
��{��	F��J�e�ڵs �쓤i,�w��v��e�7-쒓�{mh��ÄeԼ��*+Hƞ�@F�J�ɑ��he�r�<Ǜ4���qѳ��0��c$�v�8�35�B�����Ae��6.�u_�	�^�r)��^6�p�艧g.K��!舂+n$�h(�/4]�["���5�n1�jGV�l8ۆ]�M��4l-��8�Ǽ46ʄ��t�f���(\��3a��m����e���k(T0���V� �������+�v�S��Kt�5�(����=�
��+�M6�Q"s_fD6L���W�%��LX��/[�P�׫,�@�F�R��G4i��5�&Z��
T�a��;;v"Ũ�gtú�t�ԫ@��cw��sFF,h���S��S5����P��,a)kQR;����Q�d9G�ۄnGV�q�Լ�&p���{x�K7Fֆj��EǻY�d�M�Y�\�;I�3�WQH�J�se�c&;.��%�"�U8��t2��H�>��<T[��r�ų+4�A�^��
V�S�F%�F������cb܊t�f���e�2:X-��-�$����]�Έu1Y�7�!���BХ3��K�l4��㬺����3Z-��v�Q}z.�5��!�qK�z�h��D\�9���t]]��c�}�`�	;
��I&Y�̘�0B�D`���U)� h�YzK`�V�I���v��6Y����t�u$�Ah�wp�ײ��ђ���Ki�
���L�A�u`M���1�YX����� IG$ON����P�$��p^�MyAc�]꤬�c��*�ɦVX��R�볱�grL�wuh�����|��u�0}7rME�[[�ӷ0ʎ����u��)%mf��e�pZG]���mR�-c@|�=u�a��!nX�;q�gV�3ցu9h���jڣN��-a����,ʙ�p�z6�T�F��������ʬ(�o	��n+�A��mbI�qn�oǦ^9MVe�bU�^\�%�G4e:alK�7wU�c!���լ��M��w�S�1M��֮�+�h�^lh]�٨4���v^0.��hz�����>�\d��6�cq��ujK��Ђ��n')�X��ڳ�d�{�c��Xq���g[e�'(I�n��J�G`��i������x������hOmJ�����,�Bb�NU�GZ�*Rɸ�-{$���sQlR��u%X�8�����cq��*UjRܻ���T0Ѕ���FV�{a<
��S`b�Ѭ&�5Լ7�)��jM0hj�XCml^hB}wc+Nd��z�0nJX��
�Ӷpf$� eE�=.S�&�$��g27כY*��T�%�dU�*=�i�&b�0k
� X%�@�,
����ǆ�(���YF��1�OL����ǁS6on^��V=m
� ����,	W��-ufj[{P�^'��F/"�xY�V��Zv�i^ںҧ�iˢwv�S���D��M����bw���cX�ͨpLݬ�V�
������,:��Y�iL^�+��x�B�Ks�+(bz&�p6S�u.ک5-�he�f=yzR�jY*���*^�Z+t�4�b��n����) �S~E��;���)%�QX�Tw�ܩB�e�!��ˊ�a�OyN�Q�rh:1e�GE[p �4����B�ۥm�SA��T,ĕ�,㤕#��S$n�y T*Ȳ���xH�2�,6"E�.����˸Rh��X�v������X�9.�"wRb��a]Dj�j����\�-�ۑbDۤ6SI��		��k�σ��J)��V�����C�ϝ#[�#p"�l�D�����*ZL�A�HJ�[L��M�Zre��.�����Xq2�U`�E�
��l�Eܦ����r�B;�N�0���5�J�hň}	c ݼ�t�:a����N���U�8V��V�`F�,�Bf���OM�����݅aɘi�m[3���E���J��N	)�U�ц;�seZ�#�mXT��˱-��/"���)����܎*Eb�Ǖ	��Z�x��b�5�V�-AY����e�(�m�,�ȴv�m��[˳�+��t>�l��3(Y���"˙/U0!hr╖Kr�������3�[{[��1k��B�,�YE��@���)���i�A��U��[
۳���	b&2�2��5 &�BUʷN��Y�b�VY\ �����6�;�	�J������&ݍ
��U�R9"�m�G0����[v�FЛ,;�6�+u� 'Oh\�o@�D9�����;�]��ZT!�'�����GwW[QL҄��� � ��x�aZ��Y������QJՌn�6��6P�m�֧v�P�����N�kV&l$X������
�&F6��j�(mލeKf��@�w6L��) ��I]�Vsw1�ˊ�fcr]PƤCu�27Y����̹��V�}��1,d�;S	��m��{�d `n�D��) ,Ӹ�.����wF�;�v �j�.� U������ۚ�JT��c��T����K��A�qm=��0^��KP��}���J�܊�(�`�xNZs-%iŐ[�V����e��2�,�b[vȎ��l�,��&LT�yv��S6I�r;���/�U�bT�HIcn� �QP*>����U�T)S�q�ڤ*�e�3bԀ�cl���4)�*�#a��0O���i�;��]&�oF���U�M뱙���hhPdm�/Cv7�b��B��N���E������[�fa���j�b������(��T7����R[kM��'��dQ\1�����MV-����+W(�% �FV��Ҧ���f쬛�/hU�A��K17*)���
h���`�X~���-
&�!A����5r��Ih��G+v�hGN�����ڎ��]�r��t����C�̤����!m���ѻ z��b�T�S�vV|�mA���{t[A�Eî����f����ʹز��M�Aŀ�w�h�鷘�R[���7	X�6֓�����-�"��ԩe�w"�\l�d��8Yǐm��aЦ0�2��L����_v�����-�
6�1��[Ǻ�͋������SA�xb�MZ���v��-^oή$*f=�IՔ��.�ԩ�R�[֜N��j[s
L�n�"�\#.dۤɬrŝ�`w���&Q2g�Ì�ֲX�8�k%<��/�uB����Jе��LL�4.���%�ҳLE�vUmh�Le��")�O�U����X��
�������/f})-Yc���SÀ��?�^Y[��d�f�Ak]ȶ4r�ʩ%�6�E�X;7C��աY��s2v�7�h�&袱:j�J˲VJd7E�]	Z�q3��;,U�4�nbG���[���F�;H�,���бyE[�JU�#-!/� ����af�]4�ڹZ֘�fo c.8wif�i"�����M1���c;�2%x.����3p]�7M����,d�fS6�	�dam ��۔.�4F�w�QI�U�,_Ck�i�惓v$���f�*/뱘�=�w�2KR�M�,k��ʲ[���ecX�hh�a���]�kr���Wi����`ԕ5����[d���@ռ�l4�nۼU+��h1X���FSˋ],���[����R����m��
�{+��3�2�Y��F��y*��:Ӈ7lf�۷��MTK7`9-P7P�����Y36 ��Lf�4ic���1+��XUn���o~L9*�m5^�b%��ى}�
2Ľ����g��S��6-�J%Ll�Q$��I�JR˭o��*�ڊ2^Z�NE���5w����M�D��RF�Jv�=H����t�{�ȱ��"�{F9M[ii�Ԥ�xͭm�[u>H�qZI��B��D0��T�c�x,�ǵ�k�XZ���c pBZd^V2Q9Øedp\��ܑ�f-z]KLIj�M[VM��Yu�VHPBά�r�Y���G����0k�a���[��U�Q2�9�%��9ב(K炵^Vw[�t�=v�L��(�ui�7f	ڰ�P�\�4U��[���5:��F�;2��qa���pͩY����2���F��Z �ֶ��Ԥ`�IƨI(�AV-b�5j[ZnTNZN��D�n�<ު;���i�5��a�I\ګ�)��yaL��$AY�RFݲ3ڈ
�Q
ʶH*a�� �5�����YWR�*��{Qӫیh/o%�l�t�C��R�Uy��������bA����&7�Ș�A6ACQ���:B��eb �<�V�+M˴El2�LƀŅ�P��R��ҭa���'#`3r�N�(^��3�e`)7
v�~!�{�
��wGN�܁�#e��m�e�Jj�7
M�F�Ɍ�)��d33*M�cy��CiY&<��˼�ݽF�Ӳ��6<�H��mǬ˨ό0�ʲ&��*Kh�&�\QkVr��[���N��;m� u��F�"�5�9j���J���ڀP���4�T�[W+h��� �n���)�,�S)B(f��Y��*�u���
a0��"�T�M��jZӢK ]
*U�ܢa/������9��ݵ���4��	��LhXZ@eح0��u[n$3.���E��{i�K��U��
�֖�eSHkaR��A��Z ��Ɖ#JS��7�U��Q[���������u����2�2�'sYi�L�bA���[B�!O�����O��z(�B��,]��ؼ�4G1�`��H�f�к�NŦ���k(%���bBab��=Y��[����t��7�[Z�oH��ɺ���sZ�yZ�����;��˗q��9�U�:�=�g!�T2B��*hD��1��r��e�62^���EJwj�B��(�UP&5;�,����ʏ�dn�.idm��,��ζ�fȵ�Չ��S��]n�ۦD�{iY��>��;�D�?L/1C4YG-,<�+d��ETX��J'\5j-�qQ��k�m�U��b؍�����%v�b�P-M�봉��)�5���AR���m�TI�e��S��۫chY�X��yA�Fɶ�{*ٻm
k.����r�0s-�B���F��&�U��J�M���� 5�*R��($��O2����D
�I��(��V�
ɓZ5��$�+[��f��H���ڻ�0ژ��m��ڨ� ����f�-�t�Ҩ�nӲ 7�X���ӭ�JvԚ����Z�u�y��I`� �bsIFa�/I:ksm�S9�<۵�$+M&�r�ѳ�'B*�m �c��Z�[�`;��˽6	Zs�V8H�rk��Y�=-k��V�d�Lh�^ثj���]A��ɥ�9u����,4�U��Ł��zK9Y���ڂ�������Sr��IPͦ��Jf�5��&`[JV�²c(��Q�ZN���r>��XJ�4f�֍�%���Uj�{a7nJ��q%�VT7�Ј`J��T�f�a�d��r����d���u�cN�iL�v]T���F�j�H	iC&!MeM�12 x��n5Q�;Q��G-�lZ-������P�P��n[bɦ��[��ܵF+���R�l�&��.�m�?Xzr�J��,t�ހ��<qf@�*�W�U�H����D����C#��it)=R[^U��g]��&ܫ���z�ԃ��x��Ah���-fV,[^�:��xqֳMJp5�b�Z�+i2�*�j3�+B�i�[$�洤Y�� �71B���sfF�7	����n�Җ���ti+���mH��T6Z�f]]Vj���ի���eh1a�j=ӛn6+ܳ)��O��x��SU;yH01�]��p^:G ?-��L؄��nb�9�K�N=��C�(Е!t�6U��ژ�U�G<����6��!�@
�oh*��{W{u�h�BN�+�5wHE6݂{iG&о�ՅX!P��e!vu�Y��*(�	�̿���ݏF˧�e6�����`Trc�i=h�pj��l&���e,�30�B�eͬӴ �A�S:/,���!�������0�"�iP�0�D>��W� iN7b��W�úv�f�nYL]Rn�7U*)�K�����K�u"4l,�P܆^]�ۊ]LC���t���z-��ia��$�)�XYs.�l�l]���č[tl��Wz֥tE;D�mk31bĨ[(J��=B�Q٢vh�e����W����u�7�Xy�CM��
{&ڢР��A	 ��z��$�s5�M���)�pX��+�M4���0�ǚ��H�	�[@92����=49����!W���
�lS�d�6�Vj��r�,ج��i&[&����x)���H^�K*���;X�T�y)}.��q3���Jb��`�2&u\�!Yh���E��(m�f�Vh�t�PnM�@����M�Gk�$�_b�PYu��Ř�X%H�>t�E������m�-+��D7�2H/Y���Z+ot�m��`�vy�����f�$i]=�7��,��Lz���̛��2�����9GHI9�"�8��4p+�A���s/7���i����d�+�ݶS�����y���x�Qw����Z�wN}{3�</�ӧ�'3�<D�^<-��jQެj�Iow�������G��s���'�5h76f�up��.в�B|����.�&��['E,x"�If�o/�|A��M̮2���"ګ��9�z��u�\Ĳ-Z�Ven��k7r�WR��b����X�F�O�C}�u��]C2��؟q]ۢеYJ�ݭ5p -�aA�{X4��T�N�.BZ��wfe ��+e*�n�Dc��u��=���˳J���rfv/h�T.�w1-��c�w��!l8�kz&�#$��@�kx;��3���㉻au��F�r޵-��ZHԳw@e�K��)wX��{/7�/t��|���<�'-�yL�g�c��
��	:;��\[�e���Ӕ�m �:��#�3Q�D�[�η���:'O��"�krb�:k��<f��!F;[�K�� ���ט��ԫWP8��^Y+���N��-
�/_=��I��NtA|�V>ܩCFk�(+돻�N����ܾ�О�o@i�Č��_J�7-#�1>sV��'Z���j���X��_VĄ�+�If�����1��M��b��(,ޙK�f�+�Or��g`H�80�;��n>��M�Ϲ���mG�[HM7i�,f�w��F �&��-��Oo��]�m�ؐ�X*���k�Sks�}Ε��]�故8�/wl*ۅ"\�!WN��;�X��p<�T�t�Eq)Ϲ�/9R���a��u���+��3U,�@I�qԠ5Zj����4Cyk��)d�wj�Z+�[i�l���ߴ���2��Ft6v#�)�m���dMVԳ �x�{�ff�-���fP��b���M]�\�Z���Y����8�R_��Z�;|���y�];����d����`��P�)a,�zz:�1�y�9R��oQ;����Gr�t�.�������,��-�6�^�Mvc�U��ٸ�o� ��AҠ���2^!���eh��J�1w�5��n���ؙ��\�hV�]��%��.��wT�1�� =y˖1\�}�Eg�j9��]�͖�a�ݝU��޸[}6�����'o�յ@���U�wCm�5}��̋2>��X��jm:U��ȡ#9X���R9α+�ew=x,ԏ�;��3��˳MBt����<�Hus��v��V\r!:��n�|DdΠ�]o��Du��=X��<G�i��h��s'8{���SYg�{�oXU�ƌ��w^�X���e��%:��*b����J1Zѵ�5����{�-Ǌ2�ګ̻��}]M������T�7���l$��e�B�ܑ5w{�;6���í.K;~��Z�a��8-�mL=YC�X�f�.s6��S���9��d��ϑMڣx�l�79�u��p�'���ʘ$зSJ�*��rB��ۗA��Nu�lξ2gki��%��݉@$V��qn��\4ހk8�d
4Rv��1�F��8�G��q��Ṵ��cW�Cb�X�q���1
hF��Z\�� Ӹ�]ol��۫�7v �5OT����ZL>�k��[܇�.����{����)�uf���C�J̠����ܧ�,5���*P�C��g��NQ��G�-�uH�����2�Nm��)B�[GE�ʽTՊ�������!ea����ġA��gV	Ԇh�,���ǲM��^T�>.���p_tWA�xv���gfb�e�-��%��3WrsZ�B��p�"��/��6�\=x�m�w��N��:��c�Ec����.3l0�X-]%O��}]����#��z��j��b�u.�2���5��d�ޘL��e��|++S�����7f�v(m�����ݙ�8;uk#Z�CF_"3&�n����R�'ZK��X�L�H�śl�XӳR�&5va2�b�;.*������$ y{�F2�U㲙hk�g8�D#�ֱ$�Eu�E	��;~Z�[y� �N��nޓ!}ģ���qj]g	���v��t�C�_j���B���E쬚;��\OW�m��d�KT�Z���=���w� �/uu:T��|���p���ޮ�}w��grkFj�ЋE�u�7ub�6�A�1�q�o����z+�4���}�ѻ���F&���3T��+Z���]v�ᣉ�t+�{j��{��9e�1��l)���m�}�l�aK�QyW�\�GS|+9�2w
�2+�6�v��Y���;�EO�������'Yb�+vx�Di981���9�R�eм�tҹY�Gw�F���T�lZ�ˆ��eKdv3}��.Z��m5��>��Q�r���v)�dIա̾���oq�ۮ.�<�i��bmT�%/T�Z�
c9lIt�Ù�]�[���2����C)��o08X���#�[o[AYMC����sx�4�xQ�/��G�w�:�q���ӫ�o�P�Z/��������w&�]v�'�$'��t���-V=�}ҦVy�D��u�"୨`����*k�:�!y5V��3�Af��k#����[�aC� �_j�_e�n�H��%�މE]�Bf��2l�R�tF�u�+9N�-���EP0��
�v�Xp(�.F�,L�e���[53s,�h_m!�
l��]�Ṷ̌�Et�D�W�	a�湍��z��v֗}JY[�]b�Q]$q����nj��W��,A��`;��\�����G�!O!���⮼�F��{�gSh�>7��̔)�ͷ�^n��=������w,��Q�&;�8,o��x\��K������ւ��Ѥ��K����
5��\��s3c���:@�]짓�Nu��nwˊE�ӵ���F:�mB�K.�X$��m�5=��p���v�8��\Ģ; Cq�N��7�F�r����V�P�ˋ�N�� +��b5���}r����{9���aA�J�ֱ�ޜ�y7,��.���D�k��m��{f,�(�����:2�5��0��I.�������v��k�����+2;>����;��Au�;�hS�%�N��]<NH%�Վec62�l�ˤ��$	HuP՘�:)�'��ee�,�L.s�*ݖ3Q��,.yE��W��[ə�e)�|�BM�R_`��k9Uft��q�1�V�����CJ���l�oWv��t-Nz�� �SY]|&]�"e�������|�Mi��v���(�c�C�w%���V�:l�����^�~�]��S����r��o��rP�R�w@[/���)گ�aHܕ��n��f>��dl�����D������e���]�l��u��x�O���|�|��m�e�ۦ�g=y|dkZ�{�B�gZ�,��WW�B.��T�#p�.IkW9��	͝������V�MN��Fۥ���G�:��Z�{Y��ټvv�d��q� ���̸��$CN�W;�$>S��\���-5P�23"l��L��=��|�gV]:P������b�b��y�i����p�T(K�G�i&���֛3%J��|��q`v�Дl}a�U��Wdۦ1|��q�\{Z��KV�-��Z��;��}��P"�q��n�MN�q�㩣d�R�w��u�ns�6�t�����m�tm9X����i���v���`�̾���s-5Ҋ�ٵټS�ެrolTk��}���:�b8/a��(#!���J�$f�N��J�^V��Xl^E�m��)��5��]p�Ɩv�i�N�H�f�N]���ا��e��W���WM����_-��l]�nh�8��}��m��Û�KY��)��k("Aj��}���	qC��U�Q4;�-�*e�٢v��˴f���K��r��+�f+[�ŕ��դ1��v#G��{��У{(X�I�Ǘ�b�0!��Y58� �)�X)�F�:;b�\�%�V�G�W�)�8[�����X�ﶁɻ2��k��-�5'[ړX�Jc6��
��Z:����8�KɊ�/xkN�����)e�9�U�V �V�1wfpB"�e �<�3*�V]3^l��efX�<9d��-m�U�(������3��9�;�'H�Cd�{Dy����Hւn�:kj*R��,�3����V��c#7݋ep�D̘F�7{n��@ۗW��u\�����z���
ҷ:��LZx&p:�-���e�����2,�����,�I㹉[DaS�lt�D�h������[��~�Erh#��u.�л�ivn��h�=R��t7]*a���XG7�Q��8:kxα��5�6��XƧX�u�:�f(���ڛ�ΚQ��}r�Vt�Ǎ�d��iw��md�#$����宬�Y�>�+��Ձ��#Vk��c*�h�2��JnfgR��£M嵧�
Y]Wkot9�uup�.�(�ؒ�&���M��W3$跚鐎�m�;�x޶V��JJ���u�c��Y7��#B�`Q��t+��VR�w%��a�x��+3:(�ʔ䌒��E��h��Β���u-$�jN���ݨkS��X5��]�S��q�Ъg���Wl��yic[k�9Va՛q��'�ۓ�0�;o,��(UR#�*��v�jR�x�N�׽�WRX�֌���ga�a�&�=3��sr�\�mt�$���WM����}�}�pwZU{�ĉ�U���u��]���+-w]�Б��o2��&�>-��-4�9@PO!}&5��B�\����(HX�&x��ÌmQI$�Yp��C�.�
�g������r�|슘��ջ@�Hg#:"ji�z)�Nm(%�[���4�8è�6q���)�X#��ǠG���',/cڿh�M���_��@�
�������&�"U��B��i��o@|U�,ܗI6��-ử�8-ȳT!V����@L�9����Y���gb-�N�w���J#�aSa��������ݱy�(hwt���9�jr�P>;GEl��_
RK���(��,������X��Z]�w	�fM�ZT�=�yy����m��e@��ř���/��׶��N�ٵ�6Og��1�u!xnY���[��2��պ�l�.�1���p["�j�N��eG���y}fHD��`����j<������ө��߻�ǟ!�c���a݌ۚ�huܴ�.�T�c�рW�l:5�]n���2�h�U���Z��.��! ��k��X��P�O��tj!�#=w_�kMLO��4P�N�/���ܭ��/�&:����՝�.Zʼ�`�� �r;��WD�� b��L��K�2��ޥ��:Z���3r����j#L�^RVlQ��!U�`����Xug^'�����܂E6���y��-ۭ9�h��;7���r|���ڐc�i��:���v�,��l7�Tq�ģVm���V�fe�hDfe=F����R�ky8�QR���q�Zám'�x�nhn�y��}M��^	e���9�'$j�aV(���w^�r:5ty�]
��t��jvV��e�wGqeovɾr��O�j*���̭��w�m��5w�"��|����.�n�yW��[�)s�Vsӵm�&%�(��V՜��s��
��D�h�N��;HYK�UqX�Av���u��N&�Ŕ�  �V�Ds|�C��b�����z��
����
�p5��\G�MmoY��b����6Q�����y�LFӦ�m�^c���\�2�e3'1Ǳw=���"u��|�&+*��1(ì�>�ў��J����idຘMp�O�;(�Hv'|�[�{rR�o(l+���WigY��+��K�N�n.V�u�8�G�9C,�w�j�(\�],cn�ڈ!(�E]���{�\�Fu9)�<:'q
�����)܌RV��q����ӛ�!o2�m��Jk/7놋��v�o^��l�7M�lZ��M���X�� h%��t�o�sx�վ�ٺ�e�󏷘n�"e=Yo@��;�;�v��y�*(�����-A	����u�48#N�usB܆�m�x=�w�N�7�\4��^��K:��@����*o.I�p�V����<��L4����ܹ۰���4�7rݞ�i�LG��n�_%�]l��̏3�wv;����;�uu�@o4"����VeLۮ�k��N�L
�:
�3|:������d�!H]'E!����1���bzk,_kP��ԝ�R��J�r��t���71as<-2�A�a=л�D1�g�7%s��h!��$�=sh��9]�c�v1R��AꥺE[��H���0�7��{�����2�^]���7���]�N�9kx뚹�3��֖�}W�}���n�T���J�*�S:n��w9o���c�|����.����Z�N��+w�
ٗj�[޾��T��Ά���0�j*>͝E�̂�鰍/���E��t��eNgeiH��}r�C��;=l�{��<qV՜w�[7��+��V3��͈ڊ�e���Ԯk1��y[���/�[�7{|�Zĝ��w���"��W�����8�DQ�)��LK�|������]���聧��CTy���)����_gU�
���l�ٷ]��M�Cv��8B�]
x��*j�]&,�qIJ��I٤c��K�.ƨ�s���K7��e�E��wǋkT��s�SE6͠��M�w<<�nmlr�k�mU��Ù�靽���M�Ů�a�bu��T��;��>��w�WX"
T�bb�ds�,fIQu7�q�GQ�&�7���ʀ[ۜbr.�KA�]�V�wMȟ=gd哸��j��yt�y$u�&�n��|8�gH���oj�¥�W+�(a/[��Y��ΉS���쎲`�������I��V*�]��燖qEZ�]˷�L�K�5y����� =�C�HIK���}�}��l���^�n�B�W6�R���(��3��_L�峑m�%��2ڶ��F����a��?��BӦX��p�Rfw��(gQe���wZ��IWΟh/�/���]���۩R��zs��a��7E�Rr��{H��G1�Q�>ev�F*'�j��Ar�f�,
�B˔y�Г�C/N�&���_R��L-�T��>�^=�������)&ۇ,Zz8,��8(V:���������9'hT�}�`��9�f(�dV��yoג��A"=*0~�"�ޛ4�6号��7@(u���e�c83�D6�Y8���wT�E� �J�F!�	��V�@�q�rT�v�z�f�����󺽥%�4����u�9\�p�e[�0�%�I̖�f���vβ4�?3�'2V5פ��N�}W�z��Kc1+��c����U4x�*��[�(�U<�r@R��|�3��A���7\Ü�\���%7�ꗥ1ؕ4�v���o)V��y%R���l�:�:ێ�@y����H��f��/������J{w�i�K屋n���ړ�Y���z\7u���q�a�(�"�٣3Π�[���>��L���;r�@�q�o/��{X����1e���ƃ�w�q�q@h[�K����ǧcG�Yj�P���6�MX��aЗјܱ3B� �>dLN�٦��-2q?	�ء�.n��[E�f�H=�9��8Rm���%���9Ɯp`��ŭ���f!Y���7�=�O����WB�FkN���ᙴ6�P��gp��׎X������02��塔%oQ�`�+#�V��nZս
�%��bc���p@�拰�]��m��շH���Û�W�.Z��i/�/7b��tgdg*���hV2��q5tS:�z��0��74QÚ&�:(SOEC�SK�y2�К��z{���_]3[��-Ϥ�9��{E��fU�����Ջ*���ވ71w}\�;��0tP���C	�	^�������
9}��VD�G-�n��k�s����[4�B]WUe*YZ��P��5t�ڍ���z��`>�)�Jۨ6�68��8��`�c�:;λ�c�����Ng"�\��٣՝���ΆM
���7��K�0)���&7:2�:����#�٩��l��L�b{P��a�'->j�=��R��Y�ܻv�'V��G��بiF71�%O�b�"�*۲%�4�| �|�e[d�,�\��A"ԝ�U+��'n*���;��T����Ѹ����4���4t�Rg�{�um]q꒕E�h����
�K���*�ˆ^Re�[��/�Ω]f���*^cv��1fj����2m�]"��v>��^Nu^o��mάʝ͕��f��%��>��f˩�Q�W��sd�Q��V�=��v���1���V�ueFs��N�w
� =��>�V�,�Ӻ�s�[9<���̣)�r�;I��;X���Go2]q?;�'=���ᧃ`�/��L Ή;�0�}{,)@̡���VBZA����YIM�
��l�K'j 
7j�v���fr6�w+a
`��Wc,-w��y�N����U�5��B��=��|�5�m��r��ck��(K�]X2�{!�3���y��>'@��>O�w�Yl��%���euc��Y|���u_6v=���T7L��F�j�P���Q�����2�Vڻm��ա�V�tb�z*�Y��q�5��3m�n�}�Г[��������v�d��wv;���TcO74�u��e�K4����&�|L'��2����h$6�{��<��a��#�LѮ���N"Nޔ]�ݸ�����ޙ�3	��"���*�X:��so�[�/R��].6��0�l\�n��'��2�S ����u�4����vA�3���v*bʖ�=*��w�9�4�y	;�/�l6U
�R:'z��vf��⎐D�B�ha�L"�n��]���Rt�BS;:�|P��s��hm� v' ��z־^���|)�JL<�k3#���(�Ų�]N܋�f2�j�⼀���n��,e�P1tZ�,��AR��$%����V��!�L��"�Pua�b������\gi�´ݰ��Pk��0�'�VS\�@�e����z�8�=۪gL�Shd8��VnP�>�2qw����;+b�Ӈ!wѰI�WZ#`c!��o� -�8���K�x�Ԋ&���^V��>݉5Y��k
{y7�l#vM�s,��a[u#�|�PKޜ��]�6^�Xk䴎�R��53��=[8�;kY�^�3��'����z��tɵ{w�ҋ�I�b��5 �Z8�-_J���V+p��U�8�wwJ�G��7j��(���Fb�K�tL�����9��3{ݠ�sc�Dt��U&f��K�-�%>��P�#�2�65��q�kb�1RI}��.ʁ*AVy7,��� w>7�3m��,����5A�.qMv^1�[�_M��gY�� �qV�tn�JA˩����g\Y�,vIEk�x8�6X��qvC�%Ҝ7VImP�~�p6�=1n�n�M�|�'�eŤ���e2�n�x��̭걹S{&�0���]*�����7���4XȆ�5l��(�ql'����%�jpI�ۛY�ö�1���F���3���WK��Z���	*��L�p�h9��FQN��]y8�����ѕ)�21�3>�*�,��-�L�b��<YJ<��݋���v��%�sv�řd�)vt1vlA�G��#Ȼ����s�����!�4�4 �s�]�T�V��C xF��v���i��}e^�w��Xq�2N���	��f��jj�����j�.޸D�b6ޫ�Xĭn�n���6NR�!p�bf����n�'\3�
��(J������$�M�4����ev�jJ63x]ռe�H�mΫ,�����`�HoX�.%Nި.cɡ�������lٔ�Ffgm:F�Mjެ�B�mX��	pޖM�j�R�']�e]J֢���KZ�#0��i� mp3�f �de#}j���ؑ������`�Q����IGqu]�����1�ͱvs�X[6�х����Qw�Fj!�������{Yp���-,�nN�N�
R�Nt�Z���A��4>�c0-�f��2�7˧4J}�lѵݣ�&+:�9N�z������P����Gi�T�ʒB9ꩻ)h�W"���=
�X�U&����]Φwsy��Mu_:�� ��OM�zͮ4F�S��Y�kBڱ��U¶��n*�q����zq��ǣ��z�ӄҾj��=i�&�˚h�ws�Zwi�4:��Z����mS�0)�`��p\��%�;x�M��M���]'|�ݍ�%#���U��w_K��[���Ym�����P���P���KX�	�pz�1�v^�R��Rtv8�̦]2�^�B���6j`ޣI�W8�rv:3h�t�8*�֌�q�JF�hO��F�v��:CO(G�WP���	b�Ǔ���q��#ƚڵb�κ�L_s����!�Ӝ�޳���5!���d����\��{8u�s�ͅP��(SR���<�q+�l�#n�xػ��7�n�U7v
�(]^��sGq8�uq{\��ƭ�ַ.�ă��Մ�5&�5��Y��F��| ����4'˖�]�f�Qq(�]LT.���l�yظc���4��[�V
�
�ˊ��sIr�{wya��l���5������=��dF�#�fj�ct�t��/tʲ)�wj�]�+
wYWk��/4�W$P��)�,�Z]^H8ƭW8�m\J���1�d�����9��W��Ϥ{,���7#y �v����O�w&�^L��!���YU�Q(�.�θ5�}��ޥA�g*�.�����0��2�%b�Թ5w�B�Gu(��f+Bͬ�U�Ҥ���㕚�YKu��C8Hdo��l��4���W78�����L8EC�|��t�ӻ1��^���¥�w�GWa0v�=rbs��L4&t��Y�l��E��k��[�CI��u�Ҷ:R��lVVg�ia}�t�)h髧k��n��ׇ8L��Æ-���3�.�ʗ+m�Ի4̙[5��V�'q�Ѕ1A�$f]m%����Q����z�u�i;/���Y��Lf���k'9�3d,��:��v��ug��t8"%Q��wE,�px������3'J���3(71t��Yr¬	m1I�{m�Ε;�r�C�ֈ��4@9A���Щ�sPl�Hm���/� �;�����:�q]V�c۫��Q�rS'�qc��A�h.{;2���wc�F�����=�I��;ћ6b�_a�܅�kD41�(�vRłę����Ws��huǴ����=��U�<�6� ˪�ؔ��vط�u�OR�;w>�E�{r�soQ
�z�T���3:���/�(ަ8�ԕ��w;��ӫW_"]��zeɇHR
�W��A����Ȥ:�WX,��{6�j�B1��Vr�o!HL�ڥuf�'������LB�N�;Mu��₉9�?��?�f�⺻�<y�ސٽX��'l"폚���t	�bc�X�n��#i�b�Ar�G�r)�kKp�sh�G+N��%r��v��m���U��L1��fk`�T�>Rq1.c���!g���|TMu˳Cci;��.��K���P���rykvW99�uP�kz��m4�Vӻ鹪dt���RZ+zY�i�ܽ!k�${ѵ6��Y���
��eH5�sGV�L��h-\3�3����`ӡ�\��5���%g�a�$d�NgR���s]��=�,��z�}�;��\\�wj��}ź�Q�r�ʱ��8M�Y�U-��}&���l�Т��B5�kwk�5kTl3κ��n�i���ق�=��t��#�y�-Qv�M�!�f٨��2�<�I� �hD�Cv��wݼ,�q	�T[g(�fV�:/�aӟ%��!H�sGb��[�����U�:5�y%jxj�>�7�o�Tp�Ǯc5�'�b�{��tή�v��FmvX��J�c�;s����m8ܨ�sd��]��F�pٶ��ߋ��a7D�)5�>�bʹŝ��^oRTq�}vث�i��-����bä�e>ƴ���|��ܞBnQ��3%L|Ƈ��F������mƛ���b�G{L/+�os7��
�N;��W3�p{��uE�&4�z1�ZF��",�<���"��sR��O�-q�u��Vm���4�Ѽ��2ar�
¶�ޛ�\��D�œ�ɵ�ޚe��1��^��6c��¶�AF+i�H��/���b��s:�u��*�tֳ��r{k��;ɂ�T���F�a!8��xcdu¯��� 7\��k���	���z���J�(�4����PV�+�#�6��>�q�PR"
��0��4����F�6C5������S%X|�T��Z]�b5��M� +����L	Q��+Oj��Y 3���s*�s�w�D,��{�v�����<S*��r�U>S�&dxu�)��ʲtR霻���r���Z�ݎ�����jeN\��m���t�
<3��[��p��ϩ��^;�]g�[&P�dN�r�1W<��&�m���U����g��6Mw3p��κ]}d��t]���nw[s�RK]��f�'�,ý8%��{Q���|;_#8�o5�V5���jh��{r��3���@�{s�٬lHUx���|�yǺ���H�-�!��JCQ���5����=,d�G���n9��Z�\WX9�B5;[ʔ-��s���غ7t����+���m7Q����!W�S�Ok�weӭ���ʵ,�σ�,]�x�kT}Ώ�2�p�lUҰ_d;חx�5кu�+ܢ�^��t)ԝ�����pn&�ܷ�^��!GqD\����[(V7Qd��yӬ�N���7��H�:�Ih��_=9[X�!�XZ��*.�g_]čæ�k+�U�$�cN�N�U�1���vc<9���.�uV4Y���Vԓwr7nn1�QU��b����j�jő�r�;�"�uT�L�`�X+P�cwD��p���B��4*�Уh�X�F���,�Bw:�������9H�	$V�U�gRs�[!�\m,�V�n�i\u�N$Kx(�}c.�r��<��kou�e��|��IC�5�n�˼Y\��`��U�L��c���nY�_:��֮�G[�Fmr��rݺ\��\�.����lt	ἴ��]�4L�..���V
��ӊ�2Mܩ0��p=���]�P}�.m�6.�������o0��U9��-���f�oWoww��R��S9[k�]C���a���{��@*VL�Lq�h�̺ãk��jKA4�oUb�Ε�1
���۝�ut��O�'GϬ'@�� �JW)Ry���m/��ye��hqі���Z��i��X���o.ؾ�����P�Pe�X�u�,ǹՓ�gxQ��{���|��}Q����.
�j�N��͞�k`K��n�X�0sʷZ��Bh�0t;��^��/�]�V�r�yy�#f�[T�M�f��tm�]g%�+r%צkv`�s۬|��cb�W]�')�r������azin���4�U�ǚ��3��y��F�fpr�Բ��I��,o~h�;yR���\��s3h�]���[�f�۬[۠_0�aC�� ���U�p�ή�VՈ�*�a�_T�o+�s��X��IUa��c��xuPgtm�Ӷ�}��F�v�z�h�OB� ����i�y��.2u��]���?���kpލf|����o�(��U�R��� w�r��-��Q�W9O�w�aqVYC�0���dM����-��7�p���٪��n���w>�_䄐�$��>͖����@<��Y��x塬�
�����#�#��9Qo+H�Ķ��gZxr�䨗g�'�lط�\ܖ/Y}5����ݮ���>��X���j7�lR�F����x��F%7s�K"�DH��BAk\DK�C"�p��7M�ۘd.�ĳs2M�m��9���:v�0��(X꼲��p7���͵-�r��*��P���S�q��v��}(;}-�]��6�]ɡ,�W��ё��qq�yORi���f��GB��C��/I��an�Y!1d}���~[�R�;5�\D�ٓok��b�n��N��FgW
��ke��w�
J̷����,��O:�]
��2���򴾘�w�5G��[�'0��}ƲN�*^��.���s�8�F,)�O��2�jF-���4��g����i��rgu�<i�^�s"�D6�RlEU&�;��J��|8��Wn�g�Á��nȲ�{��MeFn���n�k�ǝ0�4{\{k��V�z��j��m�E��
��7��wɠ���{j����yג��1t�{���F�+5�'?���tw�yjs�Yܲ���!Y(�`՗��q$f�ycn>�'97#�Z]���ME�d4�s��絽F��� �7����Qi
[ -�;w�X�U&ݷ:�Uŝg�_ Nl��̥nW6$��v��{.N�I��>\��*�'�#zk5��fH����Ԣ)mH�Z�+U�Ŋ�Y�.,��/�W,�dX��i*LQ�3ut�V(��P��n8
+\���ѣj)YR6�iEH��,PQQ�PPL�k)�T�(��-�E�9VU���UKJ#U�#�1YX�b�R�T(�Y��K�E�J��ʭ��TDc5�����TV
(Ķ���CT����X��˂�(�؊�1b�
""��j��R�kU�j�j��т��("�A"V�rʱTc[�Ep�EJ�s)]f:�Q5Mj��)�c�h(�2رU]\�e�R��ѷ3ZiQ�* �-����)�1��q��T�*)YH(�TMYX��"�5���m5j��*���mӚ�[U1��r��Ub1`�&5T�C-J*��5l%QW-b�"�XTT�F�S-.]h��VZ�X
�k���Q���mX���L���[�kSI�j�TQq*�"
����Vi
���͓����}{�w,�
�M�2�\w�!uÛ8�z-���z���6�WNg^T�/�s�3�q)�F�xruڕ�rd�ձwW�(�����YdL��j�����hz%�P�S~��*��U���*6�����d̫"(DqZ�n�4���ۍ��]��L� �� -���Aީ���#5�Rp:rX8d�bv�b���;�[Z�{w˩�*r�����a��ݳ��B��{˝����t�ɢ��9�b�|��K=^*�8Ü�q��E�x\q�)���zn`��.'v�V�=�t�ݒ��HbA����l�P�_:�.��aYcq:Vճ%��mf	�(��m��Ta	��E�6}
 �A����HS�@-�\�s��Si��F���Y3_?���U�Y�WN�ѷH���>)MD��3U=��d���2���W���`�]�Lo�R�բ����x��,��f����p��O�>��<\�k��g�-�X'a�j�뻆D��-�ܪH���I��S�6��P���k�au�2t�
�����f�}.��g4�iӳVlχG�,�����qF�ϔE',��������������{�&���F+����oI=��l�����Tk���3M���*��<!;��V3G�		YWb��1��g:�2�G�<9E���ˑ�/�����lԴ��x���|*,ꊀ�!<ǖ�9��%N p�F�ms�wv��Ǧg���j.�O\#�c�P�p+٭�\�/'�wɬ�ԍ��T�1��܄�X��/`w�+����\��Юd�o����D����ޏ��n+bҼ��aJUY�3�c(�X����=x��k,+�����\�#��}as�����Ӻ;�^p|����Xȓ�g�t�>�8^�d��)�J*�����2�qZ��ڳ��-�E�7u`�� �J��*�!�xT=����2~�R�Ռa�>|��]�u�ﻸ�#XX�<@V�?y�y��!8Fm:n/Ν",���N`�D��*�I-��Vn=QkM�@V��k�fw��J�]X��>��Z��!	����x8f:{��H��3{����<�``'�C����<�բ+U�8s���1�*�Y�˦��������oa�tj�n��q�V#�)�	����Q$3��_�A�S�J֬��ΐ�x�3o%:9{�P�qnt��\�m��%cݔ�&_�0�Yqo0��"����.mJ��uX�OV�3)���y|w���.h�Qf����Sϙ�㬵qt������Л�a��M�r��b��뿄L�+��޶����sU�@T�J�b�g��8%�9R����E�ܺTŋ����ԎP!f!Iv���j�12��Q2{��p�l�2�Bx	}vE�I�����" #���!S�1T^>�]����^i]�i�q�
�t�@#�f�ͨ��7n9�BM)�)2��1��sƚn^6����'ٷ9�t3���@�y)q�	�л�sZA"ո��-����i��P���>�
�CMn?�>���m��Jj��
-Dד�L�G��k6�-,�MK����=1��ڬ�����^#�vP�^ʵ]��*�Y��Ts�;�&%�L%97wVJ�6��HmY/�EL*����EE9���p)kξTg���\��~�"�Vs���!{�*�t���L���!��^�q�Q�`ׂ��t�K���s�{���'�U
4��Ω�E�T���"�*�;��kEqFP_�ԵtsΧ8c��2d��Fv$�{,��C���|�`UT�����N��t����60�FOM9��O9��f� f\b�����%v}�EA)@M�N�aӾ(�t�oc}�#���/�Y�^�Q��cL��a@F�^���u+f�콁�ߔB:h���hy�+
���d��zҝs�B!�$�-v�s�ڕҷc��1Y/��1��5v�+r\�S�oH�w65{}b�L�Q��| ������DN�.������^\˿�zhx�`�+�$�#�:���9�.�U��t�P��u1[wb���7�=��O��cJ`�d�sq�R���虰�_����B��5o$B�O���
��zgr�T.��d��$ґ��Kt����w&n��%*&/��W|�x�U�l�y�%}�S�(���;�G	�D�Uf�Tdcl�=}ᰧNz�g!~���������r"�#���i�rȊ���"��Q�nM��&庥�c�����\�b�z!h!mui�ʚ�K�p�y����7��5B���ݵv��0�֫�q*!��3��lVs�&M�MzW����Ƞ��0�p��:d�4���Sj|�`?9]�+��[�����Z`�/��x[��;�:����w��b.zj�xqsG�d�=�s�����`�|���_�����X������j���ne�����������:��e��/Ŕ���_t�����3!m��8�<�ֺ�8�Q�{_)Q�f:�ȡ��lɆhu3���UK*g"n�B�*!{�f!�r�um`�Y���1�����6�x�v�WD�o��)�"��
�mM�aG��7��:ؾ'H�PxjB��К��}�#s�9�RwY�FGi�3y��1��9;mf����.��6��/r����!�Z�3oft��p��y�z��^�6����}귣���K_Eza�q%M��Ae��UCM����_D���^�.�ndb��md��凞/R�T�j�¸W�&ݙL�΀�k���|���/�u����]��,�h�9fs=����:�e�-��[^r�>c��j�X�и���P�%�]��o�؉��W���r�������cu�� �H��P�� ���!��L'��i
sg^ގ�#�l��}è�!�i�n�O�tm^�s��FJ0cH��s�b�8>����|�j뤉?z`n���%P���%�8p�,&��I�*s��{�0��b�sE��z�lsw�K�p+���.�}��%��UBq�9���5�qg���dBKc6=c��g#v�N�еM�k,���A�~�$��Iq�0Tk\�7Эv{<VC���t6�C�j'�y��(語�2X
�oG��i�1: ̔募N�[s�_�\�%��!���w���)`��w[�<Dzv�½I�޾��T-���b%xZ]���dͱ⛶:Ξ�v�1*h��e��[�.$��������.�jy�ʰ1���%�gq���'I*��+Z�7������vH ݠ���U.���8��ke�o�)�s�����"�8i�v�A�$$��)�n���)���p��R�ި���U�����M�Vf(&3hqnD5��j��u���)�.��%^;^*5�T��S]t��'�ܽWј�A�p��4.�yBq�r��ڊb��y͗%๪��Xeo��:����U#��7�=r�dX̑���J��qF�ϔE',�J���� t�\ݨY��J�i�L���� �J.��C�f�8��W�[�+��%����mnb�v�i#��Ro����8��,��~eP�5u�ӵ<5��,����}H�����~Ē�C�.՝Oˮ���v���c:	������<+t�����W9,����jLJ����ډ,��r:�8<'�f%R�M�dY�(y`�|��U�a�5{�X<�w܃:eR��]w�Y��w�1T�ڄ�u����\U���"6��=���Z�^U�i����k�h����뤑Ց>T/��ht����7\�8�3��rȒ���a�lUÌ��k��D�V�r��t_R73>��p����)i����p�c��=�]���sU�m��qK�z�+X<ѯt��kju���ӽ�"|-y��j���%X�**�A�}�F{��k���C��g7��-뢙�l��
�:����1��7�sQ'��=B�4��P�W�WDV)-ϭ閣1�FST���J����F5��\��'�F
�`�(Q�j�먑Ʀe�yj� gU2�r^Ϫ��nAmwjbfr���4�ݗ�}�����n�ȅi���N��="��g�+1V[qI'�w���)�Ƚ�Ɲ��V�5�iE��f�I@�6J�\oPo{��ŗ��:�o,���Od1���\'IFs�3i�dZv�M�}vE�I�����#v��w;��f%�'=mq�`��ʃ���t7������.)F�;����8,H�3�q�w�3d1�/;%qP�W�_4Cܜ!�;�M��$�R�p�д�Ȃ,�@��3Ie�TBY���v[�f[�cn-�dBqv"�Y^ͶB6Uu�5
��&�1-!�7�ϫ{Q�m�?����Y)�������&̋�D:�
�U�R�B�;Ř�]�.fo��\��9^p+��i�ҫ��u�fŭ������*�_TB�ؖe�A�誘\,�"L~�p�e=o����m+��'6j@[�[���kCGȕ�9�iFW����n��f꧛�>��گT�tj�>�����E�_�;:����}@e�����7�S��v><p^�^w{9���JT5� .l��óu�c��$�͝��D<��)`�l�L���-͘*���&�@g��1�J7����S��>��])Q���Dm��]=��bQ�Ψ�戥���g2=�."��kmv����<|Z;rt]?dmzf�l]Cq�6Q8�q�/��򪦣<Z�=a7|x�uE3:;�m����c�9�5��b�AB��4OI/��{�EA)@M�Aܲ�d�7�y�b�f���#6,�a7�G�#>+���s��3�v�k�lxK����o7m�\3yj5Y0p��J:��S��u���5�8Ɣ>�l�#�#��N�r���,ҘꞲ0�7gtf�.<�
+�>�<�V�~zgu�B�Z�|;�n���&IR�7�����t���L�ŊN�؈��s*�FrH�}Bڥ�؂$�p�X�rE��9��W�r7bA����6|�Ⱦw��%H�����i�nYj�ݝَ-�k��MW|2T=�a�r��Hk穭��m�v���:�*��������b��RE5�66��I�/���Cuvs=�d=�Y{���@�T"�}- �z�c�5�����v�ڭ-RV#5��Ԫ�B�ؠ��0��ݵ[��S�ԅ�;W�N���ݜ�oy��,��\lz��И�˥Ɣd'����g.��+�����ja��3��lVs�!튨[�ɸ饟\uk0[��(i\�ݭ���
��?y��\��Z:E���|�x[ˠ������Al$�j:Ê��<9��Q�i9d�(�Θ�89ל�Ͻq��a�d,y���|��^�B�/rF����`�@G�ɪ&�uNE���'`-ΐ��uɮ��g�}:�+9���aZ����K��J�/�>�ak�ؕ�@2t,6[}�B��eq�U�4
��}�^�=t�=6c2B�e��*�y@z��E�8��!L=toz_7��U��;�2rԀ-|-W+¹&ݙ�;�C��M^�Xu�p��Aَd�Us�y�1�wq^�c�瑿>{zs���ꋈZiI�;!�30�{y8�O^��.ӎ�`̫"	5W9��HF��dn�g�cu�PFƮ(%��#^Ӂ<u'���r��3+)���5��9�a󰝆�é�δ�o|�K��ACUd�|�Q��'sz.ˬ�$ Q���;�]KB�cv��Y��>h �Lwa�N��Z���|�A_t�w��:nr̜�����`��E���.�����*�8�E�:��o</+`L�V���G�h���]�h�}ۙ�gRC�ն#��p���x�������ݼu7mK�`�Nt��X������t���ATo�����ݞ�^���7�p�n/a�Z����w�[�7�u��ǰk�‸���aƬr�Æ�r���(���u[�6�e��LXۃ�8����
�g��ƅR�P��u�[M]EX:5��lɹ��F���W��
��wP4]$-��`%�Z&-�
�F�3K���EU�*�q��ٳ�;v.e����!W���$���31�d+͗�R�:�ɜ�H��6(m����C�]P����c�
g�(�s���Μdo��w��i�qk)�S�ӆ�\�Τ�wP���=��������j�{�c��E�<仆��ͣ-��i��%��������ȱ�#(f�Ұ��Q�Q�4�wMl��1�vT&�����J������&KRm���SP�������D��H��[����B'l��%���	�ݵ�q�N��L���I����g�e�Z�^��\�E�U(鰤;�=���=t8k��z�#M6�l0��Zc7���*��0��S�3#0ov�]{(�D��:�.����v�O���z<�غ��Iu�{H������U�iܱ�ʙ�1�]Z�y�����T+E�P���z_�f�t�S�ea�&��D��!�wB9e�Ǝ�Q��L\�.gn]�L�÷���Q��%��pd ��(M�7������y�-�gQFtA�uk��nu�z��5kU]�\�r��Ja�˧&��i�IJWBY��>����&�q�=�Q�i�Y�,H;����l��=h�Ћ���vX�˴k�:[5ڗMH�
C�n��"EЦ �ܙ����䭘3/�ڀ_7��cB���:��������M&������]I{��V��Y't�@�j�ONB��;���l����ܭ7�&FM*���@�r��T7N�%��׽�%C
��PkS�w����q�Y�ot�[�9@-�g(��w;�n�;H��Obn���<𰳮r���#�3�]>��ƈy{���.� ��aW;"�OF�]X��&\���2N�=7\�;5��q�.p5�֢�p��j�ꛜ�m�S�S�T��vVPx������ң�)�ښ����|���vۊ<��m�wKiw�vw��}} X����Y((���+�ۃ�'��o0�9���Q�-�����L�N���]f,x����$��[*�3�/���NNەϖa��7bn���̫�qo`�D��N�jP�'#}ri�ǋ'$v�ՙ��gAmk�3�]b�V�h� �{x��ju��R����⛏�\�]1���/q4	�`Jgm4l����O��>�z4��%YSx�}'V�q������¶v����\L��,\��ZG]Z�1ʖ��7P�6�q�}Y��_s&8c�X��d0%/����;5T�+x���c��E�^�<��.^sҴ]9@�g�06�7�Vh�g�v���Ӱ(���v���w+ޕ"�eE���K�����X�V�r�Q��(�2[d8[`���Qћ�[���\�wMU��.e+�Dh)d���I�`�x�2���^>��èvΧ���	O�[��N�B;|0kb �V���n#FwV��++�ONwi�&+�OkU���^��*�Tv���� za���;M�^�������d�h�^��Vʱu�V'	.���+-J�WX�E�S��W��)��Є��@i����5b#�4�w5���s0m!����x�!*8��;��Q�R�Ʀ����p�GZ��[�g]?�V:q�͜$l[:��6N�1N�I���5��o���;ΧW��E�Ɯ�tL�6�+bvH�U�]��<L��UJ�S����<�X���gpr���Z������;�� 7��\�s��B��������~�M���Jҕ��H��c1\JZUTDQ�)eU��J2��V*�U�c��(-IH�+R������R[T5s%b �%IDm�h-�:�[�IT�T�2ҭ�F"�Ԩ
Q�"�V1[l�X��4KZ�Aj�Z�؊�H�EDAW,�j��cUX)+*T��
�媈�Z��"��DQX-e-*�,*V#YZ�m��*�EX!Z���e���E�Q+U��(�*��[Ab�kFJ���D�qEq��eb��*�ibɦq�(�EQWM�*[*�DQK*�.ePZ���Z�T�Z�5�Q"�R�YUQ-���Z����J�X�+X-j
��P++��WL�`�3�PTJ�P�n2��TcidTDX+Q��X$Q5� ��b[F,�֢�(¥�Q�J�EQZ�Y,DU1-*E)YDTbꁉ�k"1T*�PqiUQH�ڠ�F�KE*���`����@@�؛˽.u��r�u�ۡ�ʅp�1eL*p�u��BHs�}֟Sw�Q�Ԏ��0�=5}��p������-���/� n�b͏����>��<��7������W��jR�B�*�j);�/`���^����X��a`�4��K8���e��,Īi�l�j�X7ya4�h/%�v��UWu=�H�Y<�����8i��r�+#=q�Y�%ӑ�wa�݈+Znp#l�WB;NIY�W�X5��e9nt�etgE���ǧWey�^ꂽ��1��m�̐�	�}*KUI1In}a閣1�G�OW+�sp�V_j�EѪ�G6����5�^���t��Y�$,`s���}�T�:v��:���%�9����FT��$��8���8؅~��$h3 �s�*$�l��$�n����OY���m����q��`�U�BiE��f��$� @*�C7���zO��gI;�����F�{{��zp�l'9�a;v&ľ�"$
	K�X�ń�"
z�uO6�1u�Hds�1�\`:v���핅���!ͨ��7n�3�C���[Kk��=��V�滼�3��0��w>2c��/_N�u$-c��L�ݴ��ڸ�<U*���0�;�;�״18�|@{��.�[6�����	@�Os8���F�(AO7�+�G�i�I�ݩ�͍���;��v>m���PreO�$^�lqfO���@E�w\���O%.!���1��&��k����LNHՙ5��ι���[B�3��d���'��꒡��E9�劳y����tK����A�틠pt�F׌Q�gza���k]B�;y7�|�9���uڜ\f����-k�][�#��h>�1*x|�
ڰw�����w[�Ku7��+f�q_Cؠ3.��0�9C�:f��-͘*�C���S���ú�z�1�W3�X�}
�Yq~�.��YE�.uF'4B�6�3�>�'�zo���g��X��6��j8��͚غ���L�T8��|�r���j,��Ns�-���we9b�����V~b��y����O͊t��{:��h%!7"d�O3�\�m�v�b��h�N���g�kj��C<B��U��1��S��wb^���S`̫"8e�u��7nU���<{���p%��P���L�g���������c�@ΈPSʫ=u���y�3ww��`��j�El�0�,�¦UZ-��ԏ,�7��}yOj���.Fv[�c/�9��g��������=�\5�LꚛH㜛;+yv�v�T��yj�Y3��Ȝ�$��]9�e��Ձ�5|Ee��e��r\�!F���,i��|�q斀���:��]=��+w�%��:�C��q=�d��F��3�k�D����2x.�փ#��s{�ړ���[�v �����l|�N�#�|�M�T�9n��t4з,����uUQ[n�k�;�+חMi�E
�@���� �Y���էʹSP�y�ɡ�T�0�̻g��8ة4:$3<�&�g>�T�b���&�[�v�f�4x���m5d1Nj�z�W�C�W
�_5ﴠt�8�kq�9MW�N��Y�gi���&.'/l"�Pvu�E��8�I�$ךQB�i��C�y�]����b��X�/�?i���~qǭn��j8��#tY{�ٵ��U(��v��n o�\�PF
��Z�޸y�b�V�]x�YpT[���.���{�@��S/bTWC�u
�x:��з���*;yM-f���vyǼLG5���2򃜷|Q���i�9H|�����.k��A�����S�=�F�(:2�u���杩.�^�.(�_U�&�V����hU�#�[�*֍��z�nϝ�
��ܻM��]F�k�|�e��h��=�[І�um�ir��-�Ϡ�5���0C���\m�8�E��b\�,�L�ʽ���b�'>����4�aQ߇k�8C̙7�)䃒�����fh����}��z�ݩ��4x4!r��`f��P��ߗ�{�_s��y}s��A��k�B��H��Z(e�>.g�k�G�~p��P���Rq��"�K#46�=`cu�PF�F�(%��U��|j1�����!�G�����<#g��a��:�:��0����X�� �Ȉ�����YP�\�و#�ҕ⌕��7�]���Ұ�#*���Q��	���j����`Q�>n>f`�:7H��RY�T'pn��{]6�2��)�����X�b��#1HD0��A�( �,I�s�$�sծ�!Z��u!�OP*i�0���}��K�T�{g�<��_���m=����)�b�ҵB�;'6���.�â���dB@s��J2�C8YÆ��b����a��ù �,
���8��۝�7ܣ��Im�Hz9Pf���t1E����c�L�u`�"�l��YO�4�vV[�V�h�?>�w.����f%I�;I��S�f�P�G[&t4ú;�.���֎�q��]���9n�]gW)3f�pǪ��8{��Ļ������XS�E����d���9����mV)x�5%�C���,�����-�{�1��~�GK�<p�˔���Iu	5�S�-��QC/��j���U��u�iwK�T?ld4g��>�.^E�H��k�))uP��"��<S&�����O\K�X��q��jA= ��@S�������c�!Y�����X�s�	I���t�	o�����"D�O��6�M,�3}.!W�aV��½r��jxn�t/}��M(�|�"z�P��&{c���{���t}4�=u�=xe�A_A~�a�v�*.j�Y��g�õWW����Î���Iv�w�9�=7�5��Q�XCB�6���k�:�߷%�{���A��3Ѫ�iY`���"���U4B6'�ɻo�b����������w6�#�b�����X��2���������i<���:Df��&<�mcP��B���t�Qd<�y��!�r�Dv�{��見�)-ϯ�L��V�m���j[����\yN�ON=��ͽt��X�i�H�h5�}AX���	�e*U$u@ٍ��:�:㫶,��V�Y�*ŀ�R�G�҃��l����ݾ�u�u�D���/��wu6�*��Z�����kr�R7��	p�7F����B�)M�g	�V�z8����s2t�``���U��dI[�0'�^S���E^�9����:/s�&ɕW
p��zK��IE�qG�������#�����Ȏ�E�.�ge���V1Z~ͮ�e)5
��7�_�[��)����ثj�q��������D�y�*kione+�Y��UA+�c�!���9��/,�/�Ҕ��W <fIp��IxX.�:V=7a��$�"�dT�:�����+|9;E�eC�Qi۱����oz�gc��bkyl����f
V��E�4Bܚ�@E��뒭H�kɺ臶fV��;ټ��5�:�4.ۉ�_-��Iﴆ�S/�nT9�x�F
�~�7o��V�0{yk���;���y��nY:���c,�N)��b��Y�Bc�d_�-U�6�����-7�'1P���HV;�,-tK��θ {���j����(;L����n���)'���u�3zv`QX�N(f^XY0��2��3N8��nl�WO+�`TAN��w����u���_��b�-δ/*��5ʦ�����<.�����<fs�Q�@�����9���v���Յ,���v�y�(��Suv�ҭc�5IDu�+st�x�"[Mz���×����1��̬Ԙ>qma�{�9�3��t�*��uXO�h�}kWA�%�ڗdD�d��6�h�j}t��iS}a��Zg��*�k��<Mv�ɳvs�q�ddFP$<�(�^��[�R�:�Q21P�(t��*䗳�T�_�޶��;��<첬�ܽx0{<�,3�PV՚�(%��?6)���Y|�c�ą���۸Xhc^��kX�MVH��Q�7N��j4�c�coꊀ�4Wiec��2��3�+��a"�{Q ����1����J�w����ӠݹW�mOe��(Gf�\�>3�	/�!��T�9ǊM���r���Ψb��;������S��a�Q^M+<�V�~zgu���X��v��8��>N��46蘿D��#{dUL�s��i��P�`�A����I>�m�ۊ�W+2��s�3V]w0j�B�!���t������;7����Z(�1ƌ��	jN���E�׫�[Y}m]��
�����:
PM�D"�!��������x$����<�a��s��b�Y����>�sn��R��JPT���j.��4�w��`�.zY�����3vbf�ä0ۮ0Û}� ����2��	�c7#~FG���3X!�ґF�j�S'R�8�j����=�{����G2�����mAute�,�SF�^�s�.�.��Ƚ[C�I�t�"ʾ�(�6q�γxt��ɢ:�%�����;�X�Zf.}�k�t6E'�X�����ǹx�ǽC�����޴'iY\�bs�8Be3�O�����n�X��F�t8�N$%�UP�)��u����Ld��z�y���|��y�&.��I`��v�[���crFΜ!X�wu�`���iI9��S�y���e,���١�@����!1��+#z��Δv��w�Xސ���S���j(�͈U�-������g�{Ҽ�<����vRqTh�G(������ͺ��������w�\��w��v$�oVq�dɽ������W��7��U�<Y,�{q���i}�LJ�������ذ�y�+>�=�S�@Ƒf�4��g��
�q�}�5�r��A��� �2;�'UT)djko�cu��*��	�i�&����w����~�1j8��遛F��+&iE���!�v��Xu<C���:0'/������W�/�;zs �5cҨ%Ჩ�+C�L��FJ��;g5�p�?F��iPb����S�zj2gn��Q�)���� �ᝆ�LF��u��}?=�x�K9t��ϹaN�C-��GV��c� �)Iv��_'Z��k*VR3-��铩^&	ͬĹft�I���:����J�{ۈ�կ<�	>�f���&��;o9��{"�QU[��L�bgnu�;�V��k�Z�NWd�(^Nh��G�@B�/�=�xJ�.LL�X�=�t�o�2-�ʎ�
)P�X�1kn���LB�_G5���@d���P=��Y�H�'�U�#w����{�1��-���xi��	��a?&.{�3��^խa��3�(vfP�5�v����g�v�M��p��!R���3]�=�Ӕ����l�}	�0�V�{,���6Wi�tvS�U���+b�����M�&��������b���.�#Х(�/�M��)��ن�nd�r�cx8�trr���N鎍��sZ��QMdK��.���C4tٙ��>�J�����o;���Ӹ�x��"�đ��d𗋳S;foA{�"�}s�� �n|�e�
��ΔomS��t�:3��v�X���x�2n��D��򼦓X	�J2��C�]��JeP�6Q��G��P_l�<~Q~������Brݺ�_����'��ϡ��7�5�y���� �;���5�.hTOkI����X�s�]=��	頍��K8��amae�fL��`���w��5x�:I"�}�<��W��4{��߆v�ί��6{G��7���T��.ՠQ��j�͝7wgD�@�f�ޮ�+�]g	u����m�Z{r�q�Nl
';�f��@�f���۬)񕣺��n�e(���'�S�@&н_?���}UT���H��rzͅ���o¤х��H��w�0*�!P��v4�lh׊+��Ø�P��R2b��b���P+!]K��t���c��V���k�nMD/M�OZ3J����ތ��j,��`����Dv�{��金��>�u�jm��[C7�!3U�'"����R-8Ql�)B���h4!�&93,���7P�;J滩�46g����uǎr^����>�(�F_��2�_�1���2P�Z����k%u�s�uwS<�Le�n�T�Y��u��'d�v��Ź���,;��Zl�Od��W-�]�V3΁�K�rK�-u�_��J2�cs��v�#�lV�����vkr����L >�7�)�iw\/(5��n��=���+r8�nڃQ�{f���]�x�;pj�oG9�p09�BM3!��&�rk�@gu�V�s�9VyT;���H4�f��dF3��>4.ۚ�#c��k��E�6�C���+��[_%��x�N�Z=j
�Ai
	/�z�;�xN���Em�tA]��|# I�oZ�{{��붖� ���p�vU5�nKC���X�;⣽݂W:�n�� EpA^ER��zU�\N��2�L�c�d�;�ᒕ�ֵ�`�J�1]�C]t�[����9:��ֺ���h�C��2>;�l����6��4t��҅7����=��F>Vxg�F�*�M���%��7i�8S��١(+zu@W]���7�_<ݽ�{�v;:Gh<��`U26gZ�-��[�y�1ۆ��$� �g�*��C�VڼΩ$�ti3 ���^*�B���vD��u�N9vP<�S�.Ό�A���e�Mݎ�*����U���v]�����u�\ԟ66��6!v�b=�*6:"��d��l=��5�����qh@J��nVG!��;(�9j��J��9/�;%�n޺b�AV 2\Eq}N�=Q��Bh�e=��[;RٹƓ&�\ ��j|Qa�]؈&Lo�v�*k��C�A��N�����sM,���@��NuF�z8d�͏�`|7�L5]m�y��R��U���+L9g �0��]�δ5d�q^ݹ3�=��v�F��9ˤ���@k+�f��}Sl%�hܹ�v�Jm��cl�˃��
8�-����crڍM�Ӕ�/�/�<�;�o�(��j��z�����W�0��NN�b�hRR�9���.j �p�=Ў5�2�[��;N�]�A�؜�'�D۴�-�{��z�xoN��[�x��`|�8�u10+�]]�(u4�+�s��KP��Y�����$4��]���&�U����3��s\���
�.3\�t��!�4��1����c��n=��S����׆�������RO!SQm��ܶ�`��d��zr]�YJr�
���u	]2�8����ʚk�q��y|��)�Ǎ�H��jK5z��\�T�0VNX7�Cy`�ߢ#�7�5B)n7Xw�k5v�����־�s����[�dhf��([�&�ks���vs���t�/�ӥ���H�������JkB��'���]��v�S��Vi�k�� �{�^����z�)��R-`0���+���"���D(jF��Ε���Zu��	��x���u�C5��L� ��\Mk����סVr�1�����ԟb��|g�x��*}�D[���-����m ��7vk�[.��c϶���x��r��]�x��WZ���%���(�n�k�5���zw ��n�D+e�J�E2�'e��՜�5���]@���@�y��FE����I�u5M�gW��D{(��
��ӬP�P�o`Su`�sqbhVg[��o�)�V���c�uH�ݪTdj�Ů
�l9�uR�QB�f��C6�=P�YN�C�wq���E� �i�_����<}���^�<2�����k��1��[)��=�R�"��>1h
,S�"ʒ��J�E�

��m5�mPTm�J[b�!X(�3-U��4��#"�m�h�(���P�B�Yiee�!Y�DQ2�(Ԫ�*�1�J�Cb�-�e1����Y,AU�(+R�Ab�(��DPV���%AQ"%kT�dX(*%aTe�F�\���".R�Q[J�Q*E�*"������"&��%e�
�b"Ŋ �lQP�DL�"����`�Q�""��Q`��EUR�*�R��ȶ�H�m��b�V(�X"F+��CV�YZTUF+KP`-IX��QA\����eƄS+j1��EdD*������"[*����MZ,��aEb�c4ц+
""*�UR��!ie�)V��F(*����"F��ZQZ�b�4b�9k*U
�j�1WL*��Z���`��V�6+JҭJ�m�kF�U��(Ŋk2b�h�am+R��9KZ�Z�iZ�?�|M Ʈ�r��f�#5�SΝ�i�N �e�z��ە�-^�Ѯ�����ey{\֫��:�Y�s'�#
;9�N������ݾ�Sg,�7�5Q�yG4�2Z���c,	��-���>�êGE����GD�J1[K_c�s�}[tE�Y#��Q��.��D��&��}".dV�1��6WF�����ΫZ�,73�b���*E��8љyadt�谶X!�{T�8�KqF�8�ɸ�۪�-0��dT���΅���u���Tj?d��i�����8�M��u�l,�ԗr�bX���9;wb��()P���>��#N�[��XԬ���\*�AhN'a��S�U��̸��?x�х}δ��s�v/�Y���Xke?6)��������]�Mwn�3�����f��,���P�@:wǰCQ�����\�}�.�'h+�9�UZd��Ձ�S�x�ڣ�rO-�<]��7aʿ3~S�|qB;0�\� �4ޥO�eU�-ԣ�f�(Y�H�!��xP����W��YohB�ҠӅZE�������4j2����$la<��R�[�*5=�rҭ7J��:�Fk�E>���� ��uJo�e��E�����R%�-�a%��~&2�Ox���\z�2���h0LJ�~G:���P���+v��Ș�"#���S��`����v[��������f�����*��hg<R��Y*):@(VÙ֢pJ]qv�{����{ԝbksTU�_�܆�em�f��3��?�߱֒�W*#iި��L����;��F�/%��n�O�K��`��%עe�V�&S����Uom�6�Ȫ�ɨ��r���{����qN�yLi夆�~ÞA2m�1�wK����Qu��Y�ҮEk�N}u;���Se1����Ȱ�m��	O�;'/k���w�z�Z���V�w`����wQ`��A��i���0E����dA:.���u��tӱ����fzM0�5;էs�<�M�H�C:p���;�e��,��TM����b�Y���M�.���#�Q�!m��H�.�q���Y�U׽M^�X��)�!֭�<��}6�u��n�/̙�y�p��y�[�V���⨘6�k�FǙW����w�Z�Ԯ|�-�iO$��U����l��/�K��zp��fN_H'$�k�<����bO8����A�4g�ʌ�Ú9�f�c2��0�S�U{&���緧<�����1�Y'H� NP5�@g�}���26ܮ��!v�}XtS�n�c�t��x�^���ǹ�$;�)�"g_dNM�\.�pꫀ]�^C��t�m��'�n-�K�"�d4���[a���_JёIhrMX�CA2��,�8���(u	Pf�(���V��:j�s�1��M\R����x�+�f�Muw�>�F�{A� �I��Z�=�T�)T��M�z�ڍ�s�:*���UƠ�񡕚�q���-C�W�`�FDK��pTz0�y�A�N��v���RS�/&Zfd/t��������CV���$�`t�v�*�\�J�%B9��5��P6\�����L1U\��y
��
1����&u��1��#��+��UBq��v���}ۊ�+7]y3��bf�Fq[�T1qǈ���"�ӕ���D���@C���L�ML���W72�T�(���yD?Fެ���59':ڶd�لu9�8�R����A�L�a���.{�uzעF�-��+��!�t3��8h�ܛ��l�6I
T��<���3��Y�ټ��Y���:i���w�H�>�ؠ�Hj�/�狑�/��4�V(a=����r�6�ұ0n�h��f��;^=�T��67%8ԦH໨I�R�C��ښ�ۥJL��T\��M�Y�@��Κ}'�D&F�0V��D�y3%�u��7N⎛��Z�Jx_��]{�X����8/Z +
A\��i�r��z���w+dG���?<���.�p��d��k.r�]m��s�@F��x&t��Z�T�*���ӬԨ_
�ú�`N�{����)�L�i%; ���ukznb�8N��{�{�j�_ ���]yD|3eA�"�띀mH'�셶dYS��:9Y�:ױ�N{M�ڝGҼ4%u�^w]��ΉA�yM&�A�tj�G�)��U
~���z�μ�J����ձ�V/�9���+ۗA�����Q+�a�~����`�8+-��s,=��q�O�7��帔�����q7ޡt���頊0Y��P�[XY��wfB����p�_]������1Pv0�=(�[;)��ivz�ڨ����u�1\'��k�^!�qnE�%��)_��cXb�xG@�=�:%>@V�?z�mt�$��.��q�wV4�Q�ۼ��Y=8ד�+oG5C�mZ�{����"�H�G�����I�fU�3s�7L��CqAҤ^
���N�t�!�+N~Gd���R��*�:���Rp��w�Dc�e�佑x�BGl9�q�Vx%1#A���eЖ�5vq���z����o]J�����Iƍ<iZ����G��`���-Ξ[�,:ݷ-vܼ^��^�����������蠀kM�[��v
;�n����}�V�> �K}��Mѕ���&��l^&���Y<r�ʝ2�M�,1��;t�ҷ"��U�{W.{��(4sG]\�>1[`�RZ��v�w]��;µ�묝�� �:o\���������f�oܒH��/d�N{�+���\AnR�9��y9݋�;v&�v#��NMs�ta	��E�$�����$��d\�:��]F�*�'h� �C,:ӚzL.R�Φ*��l1�n�乬p09�BC��#�P@<<��+�\<�v!݅�B\��.�S�]�����Q%��R�x\�>�ƅ�nk\�Yn��I�)�e��S�J��3�c��u;��E�������]E���%9d�"�}��Y�b��j��C�nN�'	w/'��=��U�7�rwa�����]�`����Q�%ՇAa5D��s"�6���(K��U���V����~�(ץ�ӹR,�8yƁ�yadt�赲��{T�8�I��*�RyԻrb"k��琰�ms�u�+�Ħ5�]�Wޞ�-��}��|l�ӆ9�Jw����Y��7b�p7`a��HY`d*�P<3������+�Z>u<ޡ-R{�k�W��؉��W��Ws��¯ϝ��\靋�G��Dl�S�"�*M�jיK&z�'�9�5nn�D������������Ue
�w\��j����,��&�����Z^ow
�f"3.=��˩�h؞�x��1�=\���A9��]���;��w��R�-�gR�zo=��e��ɓ�_����Z9�*v�a?�G`�HM���Yw�N��CQ��7�G�#�+�'h&`�Ӷ�;��9�V�='���F=��驙}o���&��-9���6���90���(�^إ���+U�
is�
�H����	F\	3��e8��K����(��V8U�	>�:��=[r�q�~�F	�Ih�J�{�S����;�	D�<�t�y����j�W\u'g�ʸݳ�l��͕��{�R���\��g�-�0�}ϧO�����+V�*Ô�m�*|������P�^�,��:۵�)�=�Mt1��n��������๦(S=/+RffP�>�/kT#����`a�	ݳ�6�XSb�E����%i��m-�+�4���.y{~�S��@z =�w�ڞ,�M�x�.������¥rS�Jҁ�L_������1�3�=���\���,Jt�]HG2�20f���w]�S�<ܲM�V$#���ˍ���L�~�eۘqw�H�觨?�y�P5��b>�e���U�V;��E��
��Y`���n�ǎ9.xvG�l�t��s�gle!�d�]1�ٔm-��ۄ��w���=c|���\��K�Ե�g�{�:����v}���f���9�ӄ�[��s�C��ê'W[���[$�Z:��F:�r�e]#3�K(������<:g{�%2X��'/�n	�:N@���+�Cȳ��8�t��7.���`-��yÔ'S3�.v�&���0�i�{�8]���<��P���D���9�I`���jA�@���`�mXY#JC�/�K���{�'/�������&�����4��ĽD�����;Uq}p�,Z���zURq����o<��y�k�I\U��{��to1=4�.��;X����j�`�p̨�Th/�m���3��b����,���g�������W��P&Kw��5��Y�ʠ��.� {c�LӋ�P4#g��;ŇS�;g$�̌�Xiͻ��S�P���*̲_%&���G<A�nb�?@�T�FJ�3x�G.��B�� 橔�usM[��{�~�]cʯL�G	�+�B�p@�O��1���>��Q�w� �<vx�Fm�V��Qn�d[�J�_�5=�+��[�0��=�!b����<{���%�@�����~���R�ehs�\E·��y��;Bڶd�لt'>����z$��n��sd��(�Y�bڛ<!��\�zǻق�;���AR�蜿mL�1Pe��Nٸ�%�K#]�2�C��t�FL����SFih��e:�R���=�Wr�{�,��v������D���eڡ�H�:�lţ��d��j���EI���������}=J�F���H[C�Ɛ�Jv�d9Άp��y;w&�/���b����S\Q����M�x������e��Ͻ���2���a�M�q�}̛bΰ�c%����c1�C��z ����^�F$P<J��#�͝����9��[���QMo�C<}� ��^��%{�<i1
��y�n[ɴ�ML�_��f3l<7M q>�'�W���$�:�~�Cn�9��:`�IXr�>a���&�}��T����k>}��� �>��~抆��K�Ɉ>RT
�ϻ�I�+;�&'�Ri4�^�M�����
��S?�=t������u����&�8������u<~`T�l
s���\򶦩����I�3�q�Y<Lv��O߲i"2q��6�L�#l��3I���m&����'(AJ�O��g��Ag�,�Rm*A�gRc�P�y�&<g�|�����q�FG�������w� m+<a�u��<d���}�:���g��'P�VJ��w�AH�i��5�Aed��y�I���a]���&�u113v�}`T|�P�I�΁�]J�u__ڐ�����i�>a�1��0��g�Ol�Axèg�p�i"�Ĭ���a�O��&0����M�RW��'�ϰ�&Ш)[�ړ��"���S|�i��Y����&c��7�_T��t8_=�g��gt���6�ٖCO�A޲:`��VM�Y���Sc=|5T��J����~CĂ�M}���RTf�VN���Y3��4�H/��������y �g�b�o�~�D���o����M:AC��=J����)�&�:����ɧ�I�7���M�? i�������{@�q��5~����Aq&��|I�hbC�oZ�� �Hd#R[Y�n�僚WXj3Γ�Ăϓ�~��)?%@���i�?$�l?!���1����v�E�Y�7hf��Ɉ�xi�d�_��vCIY*�3p�0�AH�P���	g�'�G�~���>�����yp���FJ|���[q��-����h�6��P�� Q���yw��`l�|[�r�j�wJ�fjzv�:{p�q�[53Ŧ4��
��f�n���Y�/�b�9������{6s�Z��k���R,l���8��y��ۤt�fN�{}7W���xx��<bf�>&Ͻ����+����i>N�!�w	��
�ϯ>��=C�ć��:�b�0���@��1f'�����'��I��%٬��i:�Ɍ�nÉ�*=��Y9/�M}�b6~���#�l��=B�����d��AH�;�$���8�g���@�w,�x��:�C��m'�+�Oe��a�X,�+���q�&0�_���K��D#��Gvґ���}�n��殾3�<��:�I�O�Y���6����=��d�����I��d��=�@�S��ߵ����q+�u����=`T=;�?�11�O2ĀH��e�w�g%+b���{42��$i���>v�H.!�C�}C<��0*
q�a�N��?g<��"�Ԭ>�>��1���r}�<H-g�����E�}�ڒ��zH��y���Ц���H�b��}3/;?]$�T��_�3 ()��hu㴂ʆ��d�����˦�*N'ɉ�~é6���/�;�Y�8�=�ܚg�V,�ɞ��(����7i��ڿ��l�UN�� 4��u��ĩg�+
¦<dǌ�T*J�~��IP�)���v��4���Ŀ��f'��Y1��P�����I���0��N �π���l���S���f*�|>�<J�3��xÉ�<�O���wZ6���1 ��kԋ6��J�0��Leg9g���J���1�VN�M!]�`/̞�C~�@dA#k�o��C����	�"f���8�2T>e_Y?&:`T�{��6�ɉ�X��R#'�����H,�ý��'穉��o$��'wCq�q�PS��Zb~I�bA��N'�D�Q}���������-�E��I��G��s�
�_��=�=eH�q+��a�M�f�1Z%gY3.�}���N�R�l�7��AH����D��Ăʟ0��Nj�a�,��'�w�ߡ}�nz��%˧~�?Dz���β��Sxn��+u��|�i�P���g�i �O���<O�Rxs�M��*u�O�%B��h�y�$�T;�a!��)��>,U�?�<Ur=�ԭ�r�����L%�͹0��9#iUs�d���G�u��m�,����R�< ͧ.F�7w��R�Zg-���q��R��Y�brõ���W����=lł�ua�tF���yQ!����0���^���T�gn����[&Vg����\k���$�I�ּ�������%@�\�i?��g̕�ܧ�a��0+��g���$�1���g�}��g�:��}���m �C�}�I�u>C<��4�"ʃ�J�;�$�m���߹|��?���Y
��W}�A AG��"�e��8�Az�'���,ĊR�ɻa�z�Y1�c�'S�>7t��W�LL>��R#�o��Ă�!���Y8�LH?����\��Z������9�;.�� 4G�@}���z��AM�{��ԝL@��S��O��`c�1&>�OPĂ�'�����;5t�.��ɉ�n���u�2��'�M$�+������޹��{�n}��+�AI��kG�?<t�SӛͲm�'ܦ�~/{�c���w��?$���?wA�~eCH~Lg��E�!X��h��4�^0�<M3L��$�&�Ci��)�ߣw������}�io*v��| �A3�ف��P�7�3m큉*79�4�y�'SH>���i�{dl���~O�����+�O=�Y��M�_��� ��`�%�
�Y����g�4~ܕ}�-���~}$q�vn�H~O�Ğn�?$YP{Cg��hJ��W�y��&�*T79�	��}i;���6�^�d��AH�u*s>�<vϙ+��8��ɤǉ�����^94uݭ̴��~dz�q��Y�AH��hz�1 ��l݆j����7Lv��s�1��2�Y��٤�8���=?wL���O_'f���Lvs��8���'��b�^�;��SMo�̳�#�'g�eM3�K�|�÷hJ�d̼w��|�J�Z��
��Kb�Iǎ���L�~d���=�q���
��36�LC�+�'���m�e@��9}v�}]mv�ݯ�������*�;<����� �a�{���xΡ�g~�8����"�E1�aS��?%B�ey�V~�R/ݲ|�OE"�Ŀ�4y�g���A��!_4�+�\Ҭ+R5WO��l�2��/G0���I?!_��;�m������T��a�����3����~Ԋm'P�<;I�H�����1�d��-�s�L@�R�W�Y;h2뙆{����}׺�o�~�Ն*�F�ykB�j���rqN�RJ.�bNEN�1l�طMh��FuL�L;q�\�ͭ��'d�^X��"+3R�n��'�������ҟS`�[��ĳ�9�8�m�����V;�bFr�u�I��(��Y=����=����\��b��+C�F�����)�+�j�Ctf����b�z��e�x�%@%�;khXzc��b����S7���,c��Ƿ�C͹�X���aQ֮2�D�0�7�a�;�o"��S.TMm�vu�v�='ݒ�ݻ�S��<��t�4=W�k�.hʘ���x�4+����r��7d�sh��9�-r��k[R��v�P��H`;y����Eqօs�T���7�A�ۇgi��t!-�G9�_g���f�ZA���Y�6�AԹ��Y�]@2�
\AV����guECs�`VRj�[���:7VS:�WL��8̊Jx\AnX��&��_fgG��� �����"����e�v�撬 �v�,�c���|�z����n�*+kv��$K��}��+�L\-�'S�x�Sܓ��`�j̩�ͅH�|Qĺ����g5Xt^���5��j�u�Z�c��&�͔)����6�K�AY����g}���on�к%��'4��oS?\Z��Ԫ\:�)l�=x��
=Pj�2�vorZNSt���N2n��X�],42��J�cr(��@��o��<�J����˽`���j�D��,k��P�L��f�a5��Qθuu�¥^͠,����v�^�T�;��>��������5�]�Wt�q]3;�X�%<�H�����u+B|1ds�³?�حNl@[�rĈ"�t[�撶>�ʘ��e%�B�`)'��]�]�ťs�7��}M�V�F�-]W԰˳_
g�7]�g�+	*���^�u��;��=���@v���$�������fX1>�w�;ZB+�)���uxy�ś.��e#�����smF�WB�qF��ً�N��c���/� �-�\v��9�{��;/r�[�:�v`���0�Xxv��� 71�p�/cȃ�-C5_b�L[9�T��ˋ�Aa�L �[
-92f�W ��Iԝ�oV\��;�}�3u3��+��$u����V79S�*�,e:�wl9����uj�Ĭ��7`%�d�4���
���u3��<�D���b=�B1N��n�7��wU��.��uvM��gbGs�]�����gB�^aJMB�,��H��ѮN�[j��rs��{�h����yM�H@wood���THf�mb��q��ɬy�%�7è�j��ȹ���'����� �?w(�K/�O�))�zW�;�_�.�R�����-��3Q���ٗMJEe��ԔW��|��Oz#�äն�P4ĩ�z�;�E��BE1.�tt�y:��[���u]!�N�Ղ;���X�Y�FUӆDZ5P��"Z��*�TX[�bbT�(֑*Q����؈1e�USYp��+*�T��F�X�EU�J�DX1D�S-��A�c2����TF*)R�AT-��	j�jDUQSV��Y��V�b)�S#XU��kTU)b���U��4����(�����Z���j�V*(*��"�-�`*���eb�b5�*���+i*(Ċ,�ѥq**����,�*(�R�U1�b��Ub�+���ՅTU�uJTDDm��DPV!iEV(���eUj�"�amF"
��
"V.\r�+B�QE@F*�ƵF1��b�J���[*
2�̳DV#RURَ���2ʢ(�b�Z�X�Z�V�J�
�[H��n�V���j�(�-*���(*�҉�DPF,X��Y�����L;X�+��� <@��J�X�5ǧa�%��n��=;�G]t9˃}"�l��Kf���枔���d���������9<39�HG�(���n�������7���q�d���z�~d�c�?2
OP����|���AH�ܓoS9��Y4�1'P�h�Nr��H-`V��]m1�����ʌ���E� �G�� }�c>O�bM�E1 ��������HbAz��a�J��"��w��|�rΡ�ɴR���gwu�
��*w��4�X�sY'�:����z���}[_[[�W�T��}�2}�*#���l
���'hq%v�ɺAg̨z��|�i�B�}�N���AxϹ�!�<f�Ğ^`W�:�&%a�w���aXT�y�c&�=J���2r����}��k�ABk�q�$�C���M��^����.��R�f���<d�75g��?2��=�4���?!_?{�4��ֳg�a�z� �����x��m1��?f��)P�YN�����M���D���A�<O����>�6�R�o��Sl׶L@��T��+'֚���Ax�g����R,��bu���%�����L'��M$����{�����PP����ք���wis�������a�$�~ސ���'�3ÿ�M> qě�gy�Ă�w���
������gSb
%H/Y�=��>��`nj��z���SɪN&��%�=M��~�?��l�ϣ8wã3� 
"�������8�l�W���\H�Rz��w솙�J��~�͞���0+��C�~M!���<�Y4��ʇ�����Ag��Vu����Ͻ�.�C_|��*��H|���$�p=��>C�g�bR��<�Xu��:�>�0�M�큌=;��AH����;���P8����ܟ��?2VzN���>�ɦW�������$���ߟL�J��/�.~��@'���g�z�e�Xi��l�zȥC��<�v�^$YS^�)*J�����m�vɌ���m6�^%d�湽��T���9��O�PR,7�,�ꮾ%�f�����~���d�;<��=J�'7���q
��[&��7�2u�1E�dm�����{���hq߰yCi�/�*
u
�$��;�$u:�.��wxW�jb����fm:�π5��V����#/���O������l����r�	�zh�t(`�Y��8ѣnj�������;et|"�0��+��1A����p��Da#:v����zi�}9���ٝCA;�N[��%�jq���u�9��}U��U4�uf��3�O�A|g�?g�&�X|�2{9ܚzϒc�T�o0%f2\��~d�R������Rq<7M&�*�0+�Y��N<t�/2J�2W�75�?@������s�%����f����u���J�LCԕ���P*8ʇ{�&�:�ך�Y��?f�a�f3�18�^0�11+�,1�VT��& q/�xI���}���(�H�+���)	8O��5�}�����M��P;/�ў�>f3�J��rE;�'̯����&�VuĞ_�+������m�ΥH/�aXz�a��19I�dR���Y��"��)*J������_��ۢ���5�ϒ۫����8���}�q4�H/�P��2wt�B����O�R,��!�bu������Ch+��~w�<z��4�|5��&�0+<w4�1�bM��2�6�ǎu�禾����w~�㇚�jAj8�,>���r�b
z�N�������'�����T���\é<xÈcL�CO��&=eC��*�Y�%�����O4��k�jO<�`T���Ǉ;��Pۼu��u���5w�$A���Ͻ���AH�I��N���VJ�f���a�
퇛���O��?]5�PY�*h<��bm ���s&س�8���ɧ�>C�������$�����m���W�U�&���$x�>Jç���6��d�y�tm
��݁�4��AH��7l?&�R)4e8��d�1�a��'�d����܁��g\C��Èm����}��l�D;�E��dF�˖�Ò����O���1�3������2)P�;��Ԟgu��>�T
�wY'���옟��4�H/R������TǏ�O] �|��8�N�z�<=�$���£�2�����2��p��2�C<��8Ο��x��c�|=�M$FN8���w	�u��M����Aqs��^$���Z���R�S�j[?&�8���l��R�I��@������gӷQ�1oug�0����g�1����a�J�X{�uf�1䯧��'�_����CiY*�a���m"�I�|�5�Aed��y�I���a]���M$�bbb��� �F�XpV��f}�|,���Pl�1��u�hr��� ���X�ʜJ�T.`3��}�B5�bP��u���ߦV[��vih9}����p��_%��ή���L�o;k�b�*����h�Qv��؆�ui�4\pZGQ�Mt��~������a�ɺ��@�Ă���1g�<La���!��z��6�_�u���&�(Jϓbu��}�:�B���Y9��I�*
E�N�������Y���?&�_z���O�M�|>�Mh��/� i�M������q�e��4�`T�d<t�g䬘�Ϙq1�3��UH/��o��<H/��3h<���h��eg��g���m J"���Ë�9/��vb�bX���OP�;�����M:AC�P<J���O1�_�ZM?0*NxoO��L~@���
Dd��bo�3�������ɤ��M��:���В<49�a�}'�ﳗ֨�]�}G�A ��T����bAg��{�C��P<��<g���3��!��Ę���(J����Y��9�4βo/�
��!���_��{�M �Q�7>�
:�����k#��3*���4G�ʓ�k�Oܦ�u�v���u:��u�&���%�ژ��|����u��+i����t~a�c1�1 �a�{i��T��5��
#⏽'����韟w�rcm�",�I]{a���m
����ol�M �_!��%Mv��c=}��@�w,�;�jm���=9���~B�`T����=k�%a��3�11�%�E�Ox�9��D\4����W�j}�'�4�^'�t1�A�%a�Vi4�����Xo������y�l���B����&�������@�S�����g̕�^��'���
�ӿ`�>��%���Wѵnd�b�������AH��|k��dm;2���m ���h|�'{C<7f:`T�s_h�'SĂ�3�h�=J�߹����I��>O�wY�&;�׬� � �������zd�ʧz�u�ֽ���dĝ��4�̙��q%B�d���d"��C�$TW�'ݦ�|��]5�Rq>LM�?aԛ~`T��f��Ld��a��>D�(����Y�˫�ֳ֕e��?!�￼��$L<�~�x�%H�y9�h�+
��2)P�+�Y�ZM$�TP_�d��Aa�@�_�N��ڲb졳�����I��K�����5������}-��G����uL�G0@����LW�]��@xz,�un�!vۼ"�˒�hܶ0�ðQKE�a����0m_��}�9�,�32v�u`�Wڰ���r�Yݣy�Q��eo	}�eoI���r�sqd؛�Qַ|�L5�㣋�G��k�{�����i��5��x�a ���Yĩ���4�q1����S��A2{��F��:�$N�^�Y�4��a�&�1����R�~J�+'m&��Ű��O]!�-��{ퟯG���c�@�#HwO��i��|��b����L
��p:�ߙ11�=�&�ɩ�~�M�x��{��O�S����=|I���r�0*N"�?$�bA���Ϸ��w5�V/��\<����$Y�DDA������&>��<����P߿����q+��0�&��l��-�����I>�rm'P�Y6w������ߴL}|H,��|d橦%����sߟ�G��[}��޹�Y&�h��&Е̛Cl�� �'Ώ7��0����x�>M��d�M������E���l9`|�>�Jj�� 1�]E	~s��v�_unf�������>�i4����@��,�E�x�P8�e?a��0+��g]���$�1���Y�_)
Ϙu1�{�3�� �Cٟd�bO��~�OR,�u%w������}������<9w��s����ɤ�'���}�ے�T�5��i�+&ZN3��I댞�w� u*|�-����%dǉ���L~@Ӊ8�|d��ד�Ia�nGǈ�<	� F���tt)�c��U]�kVM��$ۤΒ~��3��$ӶI���A��'S=;�,���b�^0+�1&>3�Zz���z�Zz��w5t�.��ɉ��8�g�ޙ�}]Zp������~WБaM��ؓ�*V��6�X!��Z�ğ=t�S��d��Oܦ�p/{�c���xw����W��~��͡�?&3�l�<B�g�S�Ă�����(��G�(d��w��6a]���WU��C����T=M0�*~~g���:�
�g�f��T*l9�4�y�'SH{�0�@�^�;���>d����ԟ�^0*y=�Y��M�_��#����m�k�TG�2��z��7>t��a�gs!�q6�_�L*b'ğ�C�YP��@�VN����l�@�P���&�J�����i��O;�kĂ�ԩ��}�=|p��>����,���~���.{������x�B/�'�m��:;AYI�c�ܕGDP�R��yTg8䕌�s;(����}ҷX����0�J��<�/���]����,<d�/ ����R�N�8�7D�m����lP4:g&u*F9\���_��{����{�$�����a�o�%��2��UD�E�����dz�YN3\�~{B:��^��[U���39���a�m{��3<�u����1cQ�]�
3������O�\
�m6{�}���*L�7��y6�{3�<����]�X5<��em��F=Ϧ�|��zv����I��ϜL�Y�E�{h��Ü����"(:۵�R��C��������Uˋlr�Q���e�ծ:X�v��>U�T�#�W8z`a����C�p-M��ࢢ��d�9��#Lt�I.�A2Qɉ7���:���
,�M�x]av!�A�M�E�)�q�u�a�@�w�׫
|�P5��5�]�\)�W�(+�]�u�q��I\�]9�z��L�%
�����&2{�y�X5�z�vl:���e��8&Z��X�����W�'OEP���]�)ɻ��UC:P"[TMvd����8E��UR6:�q����׭��y�����39�ky�;�ym򞓬�'>;D���^f���>~k���h��
j��·6�~�[�
��ے���P@J[DںAmd�y�c���&|V�w�R�[��E7��e��^��+҅��6�%���SX+�mvQ�v�w7U=V���q�r��5y���Z�Ҟl�C�6��Ղn{k�����w$�!s�߼=�x ��O#j��w��g�*��ޕT4�)\�}4][՜t�/vd��rNHG�����W_K�����OS�ze3�k!�}/������b���"��+�zHr�tw���,zT���$��qId<�gb�C�����&���`
��6�dw�3ѓ�	%�y����r�̿��f���L�L�t���%�O0��*�l��y׵a驫�D��ՉR�5�hR�մ��Ό	�蠇�^>	h����H׻��s	W�N:�l�H�dFY���*��[Z�{w˩�*�l(0׀=H-��t�#t}#��du�;��>���QU��q���.*�A���zN%p���*9���f(K*W��7��\)��24Нt��V�=������9�ճ&��ڄl����	̜���#o�yC���5��$�Πh�!!m�zB�NҌ�9��f͝	۴&*y�{$%�;1�X=I�8=@�k��w'� b��z����U�
Ц�u�ʽ�x�Ú(u�����X��B.��˔Xw���c�b봩3(��$��y/���\_u��[�n��jB:D��t�aҀ����jK����ޒ�-�x*J�2﫬��_,���\��ݣ-Q�]u��!�m-��oV�J��D�)5���R�p���_x{���z����23c��7U�1NQ.��%@c�|yg�G��̵�3��hR~U�&��nV&���ɚ]��`��F�X>F��v<̭J�+�_O�/Y���%�;7U˛���q9�q���x�;�7�|�+���J(E5�; ���8�7_e�T)�Y������:��깍�u#���r��*��w|qs�D����k4Q�F���I�T�q�hv���ljK��/�;������F�e�_'D�}R}<�=NhL*�L�M��@f�0D �a߸��o�r�h��?d����	��}�h�͞/����_�����[XY�}��2<��P���}�
� K����<܄n��cX�@������8����^���{��WF�6W�Mk�|ȳ}1�q��'\U�7Ԥ'W�b���Ѷ9	9f��7��"��΋NY�u� *
�@]uɋ�ؗ@������!�D���]X��>�=2�c��/:T�V�6��v�r��0��"�����������9o�7jfx����^�����ݻ����{OD���ݗ7���|� 5�;��C������:xR$�k�����J�ܞ]a����Z�����OM5��{�,q[�}V6�7�|��f_2]f��#����QW���� =�z��Q�m�h�~��:�D�1�[j�:�pk��E�Q}Q��ϯ=��f+�ЇΘ]:���/�葠ϣ��	F�Q$3S��_�Z�j�v?	�ƭ�V�oM ����~�L�WX�g��?&gb��B�`�@э�=�$��]q�J$m[Sݦ�����D�u�s��#��p��l/o��}��/�,�
)%*2H�9���:��95���*>��e�U�z�]o�m��#�f�mE�n�É���$�H��A p��A�:l�sJ�9]:69d������%�R9Ě	�臀����k�e��Q$-�Eq㔫u��{��f]M�~�u&Qf�w���E%5Q�G)�'Z����`��䱺z��@g����,�}`�x�G	�9�~�d:tE�Ւ��vE���u~t&sO(Ȕ��'P(7�����:��u�i�q`t��-�ܣt�P��F�	��;�`����|��;9M���y`�;�(�sęnl�V��*)�ѱ\eLk��\$��5
�3����Qm��TE�����\�F��5�5h��s8FW��H��^��]�5���ᴒu��6�{[�9�����v��Ԡַ�ħ�o;1l%D�I�N�TE��ՙع�]C[�-��&c�+��`��Q�㹑�  ��k���g]A�U_W��F���s*�V�ɉ��*��}4E{kf���O�iAR��9���9��\�
�cE����J"�0���C�_9���t�U�����g#�F��
ׯ�_@s��J.v����N����_^E"hgQPJPr�n��{�����v��9~o�4�S�i�HfH�"]�Q+��!W�Uq$�ك��t��_����r(-�v��\�C��V�Y���5�1�>�l�"@kF�wDV^Q�������^���w �s.u�jn����t1z��eN�u��g����F6�ƥ�݅��j�v��'a����W������H�<��A�����bo��ی}1�0IKbt� �PA�>�3���`���ݥ��sY9~��o���E1�t��i�-�")�ݨ	�p��r`��s,��˜e�_���x�5�~���^�MB8!�s���Ô�g�m�=��85W���g����m�\쒀���6%ƽ�T�d���n������q����\�5�����GZ�]nJ�[t	hXk(3��G��&�{Lu�l6�{�Y<�^��1��a��x߯ ���S9�{/�dYU0�6����s�jVhK'Wmİ��+�7��H�]�tA�o���u=�.��j�{@�'���Ĭ
�t�ҽ��x ޫ޶�Ry�b��iO5+�r�T���5��.�"�k�	wUTw�)������8�ej�����5�IcqEa�8���������(.׃/���Ua�z���W��W�Wd��ä:��?X!�$�uNA�G��1���d)x����9f�q������xT�^l�k8]bŷ�zN�t�Gh�}�l�3OYĪW��ٿY�#�{2�z�c��C�f2�R.��w�UP�c���q��ua��:s��̜��	��+bs6�)�gFu�s�W�b��Ы��f�}&p9����UI�:��$���Օ�M-�E�I�ns}y�'Օ����"�Di^�gbJ�H@����T5UA3%#���oWQ��s�r���oˊ��ήZ)�^��WP�/�I���[��x(fÊ������V!3U�I�`f���;
:��<���6*�K=~3<T���iJ�nK�n�U=:���'�l�6�����gǖ��R{
���y-4m��m�}�92�D�9�(��B�o�9��9��Y���\oN��Ѹ�7�u䥕6.��&�Z��c��,�k\hp�@�f�a���Κ	�JT��wCza�G�b���J���5�\�zk8j\���u��e%SZ��{t�5r_&�T�w���Pwb4��bʡ��{�P�lly| M��>͙q>̚���{,'�7�g�Ӎ��@�c��i�ͫ4��Lܮ����wu�˂+�7|�Y��|��b	�f�aEf�"T�{��:z~�[uل�"��T"��M�aj��b�ʉkl�e�A�8�\�c���g7yݖ�1�=´@*d�;���tq�E���Ҽ6D�[Ӱ�Gv�%��;Z�Ӱ�y;{��FԲ]%�]��㻛I#w�3y��mq��7{�S�����yi��V6 `M�2F���Ȏ�ogHy�.����/G���9�`ν��0a�O���m�AWEay@���X���;�j즳q�|u�����xSڋV�\Iw.�H���{d���{�G}x=D/����
��	6��ܝ7�����j�;vR�tC㽹H���	�p_<�rmOh��u=��W��[�}d4�N��%DOkͽ�z����-2�����X!�.OFp��Wf9eg_>����5��p�ў�.�{JE����=Mz�ѕm�Z�O*]�5ekT�.�6Z���a���X����G��&^S�}m7CX}aC�v��fgV�M^��,�l��^a��ι��"��Fr7J��:L${�U���<���Ui�Vq��8mj�rٳ���s=��ɝ-��W>��wkm�R7���V�馶sKj�՚s�mV�`4��ً7RB�`�ȩk��c�oCɢv�(x�VT��k����"#i���Vy���
���;��-/��Ѭ��}��r�2�D�k���Ұ5���a.��%E�t;iS�he���=��kW����܂���B�!Y��R�x�1�f�p�;g,m�u͖���i`�[le뭦׷Jw�2�Er��ml�9���zkZ�d��ϤZ-��a��.�ښۤ�S᫩�o�'Iv�H�}c�����X;+y�i��T��������K@�j�f5��c����Qg
�=}Yo�C�;�E��.oT���\�}��EvJ`WEQ�!��-tpFP��U�S�]wun0&�>A^C�Yǰw�Nb�G��V:��p;Cq�<ˣF{;�86�^Fnp�⦩夙J�p��#��ї�����EY'u-f��Ü��L��Z=Ys2��9���:�>s�ۮ�c3&"GBvr�C^rj���v;���f���	U��QdEW4Od��NN��XUfSC^9GBe�vʷ�s�n��r����QbK��8�2��ɴڍm���tt�qûι����3%�Q�o��ٝ�#|�<�uقS0��S����pHFj5br;3�Jc'�JKB��4`�X���-k�#Z������X�1R*�UT��QV�`�+V�bE(�e��,�kdX�X�+dQԳ�

��ijT���*�"1J�,���
��QV#YQTX��b�DE�.��b�ʢ.�+Y�A��UX,VEE�H�b�U����*��U��b�5TE�����,U�"�L�A�b�*"����A�uu��PA\�i�VX���T���5`��*��Ub+�QLeH���"�DDX������+��QUQALJ�̵�b�*Q"�(�B�UA]5f%AE���j�4؊#���U�h�u�Ȩ�
-J�*,���T�(���"�rءR��X�G����`���[��L��Ps�C�9�!iu���:��F���	Bu`U͎AZ)n�Ә��1�ytmܮ������+g^�O��]E��L��S�Ry��ݼaH���S��=@/$v%�)��+�v�42n��yu0���aJ����c$S�!�,�әf�;9��[`�V��3�d ���<�����H7���]>��5٘����C�|�>QbyIJ�F�}7+^��	r�m��:�RZ��I8[��Uڳl��]���Ú�)��� %vVZ}��к�)cӑ�Yl(��3Y�-$˰b}ύ�c9�/��n}s.��uL�Kj�1��yJr,�1��X����L(�ؖ����g����M�Vn�N �Ĕ�����V�U�M.κְ���&����lκY���d���MwFF�`��x�9Y�r�U����?�}c���}z�5���H���(z�d^m��w�e�M���OZ�]C�|hL���L�7�Φt5&V0g(�e17tv���gC^�9ue_3x�p�v)��LW�'�Ơ����(�x�	T�Q-CyۼEH�"�;�S�;9|zf�"��I�u������s:�J�bp�� �M�x��k�^�sg���*�ـ�v/��� �iw)�:��+;����=ݍ�,81U��P���A�bs��"ի�/���"�U�L�`)O�7�x���Y�<��j�%�U���T'�8$��Cy\����`lNP��ƛ�vۇϊ��	���'.��t\�n53mw>F6�&s��7��{�V �</����I��,��u�;���E���Kw�e�8��0�za�t�@��o5���.��S��4r�3��Ҫa����~KDh��gťBa:��K�9k�T��0ev�9���[�����]�qNv��3���S`���B��]��H��b�f앛JSld�]Dк��{�n���(�
��RF�<�jV�$�ӬwB�
�i��ɜ������&�o�E�N]�ҋk�PR�	�8_m�/�^]$����5�Į��^���u���7Š[ύ�nq��B�4�g�Cf+@�&��i}aq��`�:��kp1��rhݝz��
���r���чkk^�6���h(�7Me���ۧ6s��я⻳����)Nt� �fwL��[�
�{Y�;��}�vCzA/.��1�\���И--]��=�K��ޗx��M_GvM	�2�f�]�M ���M���c�̞aF�P�9R��k!.�:������U��Z��ub��]kXs�T�]��#�|��-HD��e�o��s��O���!z�R�-��\s�ˠZ~@���y�F]]�������s^y���Y�����2a[�ToD$fK��6'M���Z
+,1�����9S���,X���e��'�:1��=������]�z�����,���|så�2�bo��v�1���*��7���k<x����"�@���\����|�䛜۠���5�}�y�0恞���RHL]�M:�`���t&B	n)x���m��1�:���zԚtjy[�Y�VJB�#�Q|��Z^����ʙ�q�Z���RjJ7y��i4z�=8z�%O�}�h��	�盨��.���Q4�?|���ٮ�m����Y��g"~>����^��ۜ�y<J<^e��飥7����햵� ��B���"%E�54t����I���1+������ 9��z�k�WQ��ǩ��,�k���G�<��@��a>�(��#�����_gu7��j�9X�9���c'������NO�H�R832��*����[uws�df;OhK�c���mx[��+OD:��h�Go�'��u�2�@��u�l��*�4��޷�/2��<�C�{����&��$�Gf�]���y� �.��X��Is�M�v]���^>����LMi�8ͩ�<JC'}	��T�-��;zM˹��'���^�Ͱک���2�P�ڋ��+�9�/���5����P�5��SҸhJ�63���0��b%�$>�Z�Iգ3!<ĻƁ2:��|���/M��c�e�<ޕֵ�5甦�B|��+�p[�^���j�p{�������U���=UK�[��.�X���ʞ���r�e�Ov1#�YQ]�΋M��F_�e��u7;�Z��p����^,	�T=[BZ$����Cl�����\;��D��;ͻ�,�;N	W����D^���{�pq)p[̬E�Ɏ18�q*�O�g�o�~���+u�v�J<�nP9����*�����-�$)����f�.P�gKs��+��]��s�۷}KB������Ч-���}�L�d��P�fȿ6�dZ�8�;BP}^�/��\VW��,b�M����wv!�����X�i����������Y��FKs��CM2��]����n4v� ��w�D��zo�'n	!c�:��y��U�;,"$㭝�A�zZ���4���9i��%{ �@hGUuX��Ouٍ�����-�����;��sc{���j�;�ە<��y��a��ۆ ��SɅ���T���wc$S�rͫ�5�]���[����^~J@��!^)� ���O��W�k�n�`=0���o�ߗ+�������/B���JU�F�<�jV���Ya�u*��[��T�TU3���]�N������
U�#е�J��D�����9!�9z��w��rL�-��>7A���׺V=˺y�|2V.�g^)���;�
k�%�M�wr��:���r���`�ӫm��_<�G�{�.��������h�@ĠVօ��p���pv���p�i�un^����H'h1S���ǹ�D>��n��<�R��BLI����նb�f_o~��ǭ:ʺ���Z��_e��ITզRl4��}������K'�5;�Q����L�M?s�k2�=ku^���~�u��9���M����"��=���;��5��,Ҥo����ʳ���e֫�~�O��PyYGƼ�.�sf+,�䱙ۍ�E�3�>�*3D�9X�]=SOcA��f��ڳUsv�gq盞�,X��NjÒ+�Tf���HY��-|5�ػ�Ov��J�	��ƶv�Y���tjPN$� ��'�grJ.��e�ѽY�k���mӗ����M���)�CB�1��fޛ�V�^���	a*�*�1��j�[�);
tI�(��1E4������(�L�J�^�J�0ұJd_W7��ݱ�+-͛2$�巹�+�Uʟ�+���༔��w9O�G�fv���a���v�O�j@�}t�#�U��4�)�o\�d������ȶ�%g[��.èѼBP��;�1���#�+>�xv�Λ��Z�<�$���k�*����9��L�;���*�f�Fw+��f�;}.�T��Y}�w];oC��a����+�5�\�DM��/��d���iZgK����!'y��cy]wc!tl_tknbeY���˽Z�gz�8�iڋ���{h�f̞��М���|���7W�Xѻ>���riYo���'.�����E�4��QRu[
.���^�.�F�����i�t.��&���禚�D�T�n����VN���/�O�f缶��f�I)�9���廋p������p
�2����"=2����Ǣ��J�Yk(��}λ�z��N�b�a)ɻ�
o����3CY�k��H��.Q���ƽh� !`��4���Ĭ#�6{��k��y�[��z�I��d¿@pv�=T���~�{{܃�&\f�w��t���*|�C���[���Xr|q\uVV!2U�|�Z�۫��b\�K���z�q�|�)��7|�f1�l��V�E�xK�W����k�6P�Uj�3�+��XB̖���Z�n�5]8�u�H��auI�םu��s�z����ұ���&��i.�\gr�>R�$�*�>"�/�����c,�B���_m�7��<��&P�8B�� �%��v~�����縘��dn���p��	a�{!	��B@�I����Ȭ�n�(�Fzh����OABk�o{''I���a�J	V)u�U��}=B��^U��^�.������s��;:֭�t��h��T�uze�b��-�����j��$��S|���zW�vv;�Ӈ�$J��=�KJM.걘v(����L�1{SU������2�tho��Ӆ�%�4B2c1SV�j�Z3���9>���a����(v���*�v(Ǻ��t��i'�ݥm����ō�Ǧ��L�މ�X��٥W�5���~�%���rd�C͘Ϧ����ldX����^#`�M+r�'"�aR\�|\fMn��֝LV��b��nq��s]*jak����k3\(�@��aM�䔙�ț�x����4�����
��Y���]��S�2���Ll6�@T'�*�j>��3����j9��6^S��{���L�!,���y�^p����ݶ�3hDoor� z�-���\���%u�;����;7�:o�dS:��Vm�g9W��vr��fL;��6/gs֡m��p�t��}�=���L\Nf�|�c�Φ�
;ɱBC�5��d����4�3u���ʹ�b]��uj������4R�M	ifL��rR������_[���hv1�;t�S�C�y�NF]j�GJ�R����˩������*��g����j�z��K�o����ܞ���E��b�Q�N��Bs�*n{1��ѼFz>l���g����l9�g��gW��_7�X�ٞ8�T0r����{5Y5o&y�r�XM�c{;ug���ƪ�P�p��ܓ-t���S�r߷F���M��;z�{.�9����Ο]Σ��O�O�4���ǻ`WJ��7v�����M'aGgZӇ�"Sfy̸��.�c��vw��jal�i,
S�a�<aM>��S*%Eʞ�E�à�u�g,��3�gѢ
^id����u�w`+�&1d�m�n����k}�S��:v՜	�4�L�uo��g:^ '`=%�%z������r]�U��-3�7���Z���<���r�;O'j��V8�ޭY;�,��6dۤt����O\�8t��L�ۍ����
�qJ�����/��Pq��[�{÷+�[��U��{��u��@��HH:�_�-���SJO9\�FAz��S{o�����̡���zӰ��%-h��]����C&�¨�Hv�2��s��V[��i9�n-���R��>��u���;h�Uں37|��+��X������P]�5�2�9��`����$ĸ��TMt��oa�ʋ~�}���[��]��j�
cG��_{p�m�bA_n�_&VK8��$�[4��0�e˷��2�o:�XsO)Os�ΎX�}�ВΉ\\�Qs<�i��3+y
��;�Ľߧ�Z>��2� �M�����v���y��y��OZʵ�b��ڞg+Qې�yΫ��WO����6�"U��b2uXS/�b�c�텇$V-s�6��uQu�K#n��S���|�Cm9w֛�ƲT�r�nW��B�ͫV�4�_�ݘ��F͖�	gњړN�U�a�(\��hh�9s"�����<��껰7�4�OJs3����=��a�:q&n�"e	�|���6�W��c�D*���z��A���9-�E�̢ޘ^Gz�^�?&���m:X��U �= ������pե6��)�l��k�Ʒ^��7+v���.���
)NN)H[�,A��;�)ͮy�o}%b	�w>�:7���ېDݬJ���4/��x��or�0�U�c���c'wk)�iLg4qfUk!¹wK�o��(î���*����hb��-��ۼ*���ێ���60���諲�X��bG2�ћ�k��}�\VN�1�����]]�{��F�v��}�� ��DC�4�Ju,d̾sx2-M!·=��-p
�ٝ��|��X�\���jV�൥���s��v�o�LEt�K:�D�=����_��%>�І�>u��.w%Z���%�t��:�v�wJ���*ssru�lW68V\��bE?���+�Kq�m;`ضܬY����-�1��X!��&v*�V�i�P����	ً8��@M�V�����GhU��e`�6D`J�1m:�"R*�vޑ�úU����;�2���c!�)�����j03yv�ѧo�W)��A��m5��v��FKCi����ae��|�!}L��w�&ݥ�tWGZ3.F6��ּ�5�>�������ړ�s۽a�)�����ٓ.�C�W����:�s������S{z�V������n���z':v��Y���+,�J�vt5�E�H�׭Ei&0<�j}ѻ��zr�H]gfL��x[�& k�=B�NWs�U�
t��y��o�;�{��n�W�Z�xЎS�s+5ݛ�Е"'3����X��Ip��٭��S�=Fٽw��k�#b��'J��r��MM5�U7�d���,]��R
ã*
U���^1�%� 3-�f���4!��1h�����%�oC�5�f�*/VC$�ê��ݛ(X��h�w���-���r�N�}��S�B7J��2�C��x�333����;s�m��hP�ܰr/+�k�7,�ȥ��w�t��y<8l���p��6�������͆J楣��j��,|�޾����h7���X��x��8�ٮT*�ѣ�@�2�d�=�=����u��r�CB�V��vLo%˔A�MR�q�u]���H�1�td6o�F�YnZ�wms�5J�U��G9�Y��֩	�V]���ݸ��{�[r�]��Xzՙ]��tǓ��L�Rg��=iYҌ� ,e�����o
�'�c�8�.��+$�ʶ�K�i�]A����3B����w7WNE�.�j���Cqr��T: ]J@��A�\�39�j�+�cJ�Z��h[����gw9
ݟ+����"���̨*�5��b���Ţ1�����DFҌ�2�[Q@̢�5��"��V����VQ��$@�b�5h�X��ư�Z�$D��X*)�L�jն�
�UdձE�*�DF$X(���TX�� �D�3,��I���������ګE�QV2#�Ub�*3
�"��VU�(*����"�fVѐE���1a�����Ub�A�"��8�UY�U"
b��(�AUQ�!�Q�ci�1
(�U�5��"1UD+TPDQUA��EDb��X1ED&6j�eH�XJŊ�SMb���IF�*��B��r�E��E������QDA`��騢Ȃ��&5PD��"+YDr�E�%J�h�c)�**"�8�D����X�������#�J�FE"��
 |�F�y-�up�]��[�^�HؗRZ�;.w]���Ӿ���ժ<��C�̵�ɔ���ǡ$���Wcb�'���T���Oxz�b�K������*���ě�v�y��`�ΰ����9�h�.�_[C���g{Ba�J	P�P����A�t��/�y�ret�d�ܙ~���KW5"`� �U0�	������sx5���M D�,�Mr���������oN���ƈ���Mz����R����J��~
{�d�;�8�EOԳ}<7��ZgK��@�/o>���q���N�R��ș��^ou�M+ޭ��j�8�iڋ�y)#Td8��.g���ᭈ��jX��`]"�a��Ұ[��j�t��9�`(���NL{��7���w���IMK��Os��s�7�ߋbG>7�A��28Uc�V���bk�ni�j�Ԉ[�R�VZ��U��M,�gAˮt���c������{���^�doc�F��w>�ٖ�u����U��2�7J��md�.*��ț݄�nw�wJ"WA��ו-�:�w)��;Gl�X�g2�r��,p�Oד�����uA�>�6$0��Z��}V�\g��X,���R�Z{��h��zp%u<B�NɄ�{0�D��Ѐ�DK"j�ܠ�����C�������t��Bhc�k<-v� By��Vs��f����a�t$^M��V�����k��e�<�!��V��㏆ab�Ϛ`yz�w��\il��-ߨ���'�+�>x�Zz��fE�,9Nh4����٧�8T,两v�԰[Ss�)��1��K�aL�Xo�{�gl�yV���u?85}B�:5�-=^ܳ�6��䛜v��;�
�'���f�Tfs9�-V1����`\��}R�U�]{a��0�ӽ1W/,h�e��݌L�a���J;�Gg-Y)R&�<_*c��2Ҳ�cUIB��c�B��\y��9Ln��`�凥Ji4z�=8z�H�0�\����)�.���p�w{��yP*��篻��)�E7����ߒ���e꺞_,���7���˝�{7�hK��{��.5��Щj��#��r����aL�@㹱C:Iy9GF$��w"8-�ߎ�ɗ�:� �:EOE*ؒ($��iYkz&[�'3z��ޮ���ys^*Ǔ9p�����;�Q+�S��'Ј�7ٜW ���Z~������a��(:�Z���+��R�6b�V��U�i0j�+���#`�$�t���UriYw��y��0�V�]�D�g���g�<><߻/���)�Е�^���턗8�j�\X�"D[�Z�W3wjͰv� ����6ۚ�)���/�)[9��=�|��T]���ɖ�fi�%�A��
��Y���]��蝭F�^�Iu��9z߲�V:α��hZaE&�4��[O�2���Eb�y^-��St��߰�ͱ�,J����ipޗֵ�/%N�4$�d���e=�+^b୰n���׎d�o�U����]j�+oÕ=xK����"zr�k��[�%
��cwv1Y���|&�c���!��
y�g���|�ų�57<w�H�=U'�zy)��g��k-q߬8<��K��1�RK#2�_0fU����IB{�7�񽝰*�I�tj����fjޙ%�b�o$�c+��7�֧��]9ϱ--#c��v���[v2�k����Ӹ�9��K&'2;[~����x�5�a��6�sO�.�5mj�n���M<�}���;�SSj�P�Ad�\a:��L	9
:���h�dB$��x����vp�Ncf�f|6'-7��Si�A��~Q�ɼ�<Hצ��oXShq	��.�����̝㽝�.�x���YoJ��vvu��V��9qWS*���c���b���	��b��Ry���aS�j�(v�o:��r��5���W��� ����L,�oJ�݅c��u6��Ⲱ���u14��QP����C����BB����-�ٺ��e�\��VL{��Zn2�G{��}��C�vX�JJTFǏ>�Z�8�����&]6{�ɜ���lm\Ղ�-N���aE�<JC'����tK���/*/�k��]��t3��S�2�-�|ks+�9���jk�J��*ީV����.�;�.y������	*�L(�ؖ���k��̥�P�pf�w{
���r�Оe�U��{�V���ykH0��{�vY�q��F)��[��6�[	!��� �ӗ��p���Ntѧt�Gz-���+w]/WK�ÜX�%�sn�h��Į���9�gaS}I=�����Z���#�tr���dl�c��;5�W:�%��Ɩݝ�ưǫҌ��%Z� *��昉�19?�����2Ϧե�P��s��S���>*/�{qs[-�sW��߇�P�l�/;/[݌�����ᘷ�s��9�Ic�|��N��M�\
+,<�j�!O;
e�����o�ǻ;aa�8��_&�Pl�v��ыؔ�u��"h4����{Bzx�Ko�|�̷�94t�̫@�m�qެ\õ���al(P�odK�|�ؓs�v�/�]}�m�d(*"!�4��hL]�MO�]�s����b�X�wa�k-�q5�T�yZ.s�*�i�C�U���η�RD�=�@/���+�7��䖫U���(��q�1U7b91��}ɞ���Լ��G���L�j�SdXǕ<���q�����}kW%<�"�~�4��y�ҴΗO�H��!�(��Ůn6��]���(nϭ=e��w�q=���C�v��%��\-��,�z�:��"�ܺ�!��ڇ��]k�x�7u��X�O�!�]��vwP�l��:�T�����<��令����WM9;.|�M�5]�g�^.�&Ϋ��e@�w3�{�Y� 7�h�US_ړ2\�UQ�{"&&����z�0�V�~�����
�&��[��I˽ۜ0�.��v��h��sd�2�����-:�
������Њ�Q��O�s����x�ӊ)��Ue�𜧓�=�cG�Ӕ��P�z�%SR'5:7+���qW|yw$������̱��jy��
�W�-�]��y�V��]FfOi��zqZË��9�;��-a�y�!4tTγ�g��i_y_f]���S�lF7]�U#���cغ�yٿW)Y]�&����addy����Z�g�*�h��b]��ct�_L��ʟ<}-Xz�,=݌%�Lv�z��k�i�ք�#n�<�	��S=X����|�L�Xo�a\��������Mwc�j���Y���toW��P�P�Bo�ܓsQݢ�u�oEns�B���S�{�kU�����7%2�`��gN��ۇ�W\���_�t��uk,T�Ջ� "D`�SMR�B��Y|<�o�C��*��ĝ{�yD�xK�)1/1��9;kl��Y�Fҫy��\�]a�d|�v��7Lv���&c�y' b�T9j��F�.���}��0N]y��c}��F�l$�3*ȁ��)�m��'aGgXZ�U�D��E��VJT�[s���11�8�d�b����/�J��N�v;�Ӈ�"T�4DWJqm�Mt��WլLjv=IeI�{����2�to�}N�Ӆ�Lk�y=�*�i�v���m�oD��}!ms��ۼm�r�v���K0/�Z�ʵO��Y����y��#`����dvi\�A�%!��!�c���MjVj�יO/��ݨ�	AKA_zf�5����1�^�G��="\s�leMNEC��]�n�:7A��l6�K|v���}��jh��t{[a�.'/V1����T�L�ؐҋ}c<s�_�����К����77�8��V���n�:�߻�M�&�6���5�q�]F�yj�ͥl��L�M�̱*��Փ�V�oK�ZÚ��SA4,��I��Ǘ�XV�/�;��Kq�]����A̘���d�ɏ���b]ԉa҃�H�u=���%�Uv���bEty����,_>o����i�q�ʲ��=���	�-� ����
_��#-Q�>��Km�b���i�M�`��f�j�����U�d$�D�����$U�M�KC�m.�G_9����ˇGJ\�R��Z��Y乣�6�+Y���o���	�z��|���\�.�ck"&�������+�����m��$�w�	s�%�6n�1һ+/9�Ņ;v`�>is�2��)���_����VzA�`���؃i��Ȩui$�]]����ޡ�.�|�ء�M��sG��&�]�H���oc�iTѭ�Ϲű�8��&7�e�t�V ݽ-ZzT��v��j���gx��훓�W�ܴe��t(�:	P��,�U'��a���+�8OZjF����jʓU��~zp��ѢHO�J�P�n�U.뚪���#JOSɎj�jU7{\��2�8�{J�x!��R l��>�P[[f�8��oL͈�N�9��&P��q����Z�^e'N�hЄ�RR�4s���	����I�L�yS4���-�����g{k���a��n�|n�ŷ|����j������M��==���X��"ʵR�//���#X�����k��K�ٙ�jֱ^Dnbnr����+v�W�1�v�y���Ԋ���F�v��[�'�͍��)��DUC�O�U}Z�ѷ�����߽����t9sW��-N�����AJn)��@��S��S|�ȳ�e��VZy�	n̡�2�$s�t��
0�2�s]}}�z��匄��ۙb[��Z�珂J���&��~�S'j���y�,Ul���n&�{�m�g3O�#����1�j0ގŇ:����g.�)y��7�(��wY��J����kT��1{���Fj�(���C�;f*��v��w��~����?6���Z�ڴ����~ў�{I�Χ��W|y��E��z9�
e����x,����x�r�����N�:9����3�2)�\���cˎ����o��	��k'9�Li�=rn��H�Z2����㣰J�a�ObM˦ל�cB��l����{V҇=
��~�];u�������C�� ݽ-][����18G�]�ϠF��5�Ξ\s"˛��{�p���1焞)H('v)��&`S3W,
�u2)��jE�Bn_Zzr���+��S�-�t�0wcSe��ԬW����wT�8�$�����qJ�N��,�]m�5)�S�,�ꎱ�_����\��T��u����u�8y"p�>X&���Ғ�+��u}ӻ̙Up�74,ǌ)��=mᳩy)�q�ZBn*c*u��R�������ߵŷ��/7��K7�� �iXL�t�� n��̰�wbq!��̼.���a���vȾZ�m+.�n'�V��z�F�)�����i�|�V-7~�d87�5+U���
�&����.�r�V,�XVY��s�%�mQ�&�[Ȱ��Z��zV�R{�Ш.�)�/:Hj�V��SƎ��\ۓ;f4?U���QNWAj��[��S̥x3^���jQݘ���j�d]M_q��a��Ō�Q�V狹�2�*��1ţ��9C(�yZ�t��R�%�oW�Ol5͇4!��*g���k��&�u�<W"��x����_d6�y�����y�s��\�8Hn��g,{5��Њ��)cVM����^�ڹ� !}I��vq�;��WA	�9>�ve�Va%�3�x����ïU���⒊��)g_y�X8�?��Ӛc����gwOJF+a,ȧ��.�@�{�aЫMq��;3r�R���!�J)s����W��:`�P�/����K�7�/\�]�lu)�Qa������8fo)�e�����"v~K�c
ݼ��oLvRTL;���W9��OW����;��]� �oJ�2��S8f����>FSt��iK�[�,E��S�u&:]+���[AHqngS�JA�.�K���ʹ�(*m������;_�F����J�c��T���q� 0�N��8\���^fkimt�\��ꋆ��n�E$����'MN�AWW��bx��S5��G�����fQ�W�fs�3#48�yR��z�����V)uJ��:yw��.�k�5uV��J[��}1����6Lm�嗻��u�Ns�҅��q�w͒����mXb�]�]t˰�I�ы0ե����C�E��|�ۥx�)�i�Wmm�yfk���;r���&}�{z��&'�)[��G*�<��H�KlU�K��;����r+:ie\|����)q���v��gm��x����)�'{;��jn�]��g�ӣ۔_Eke��³�@u������ݎfrԄ5�i�U��V���DRw��Э͜n>�i�gr���=v��jT�Y���E�M7�)é#͠�-e$�G/Nc�Y�bM�dt�g�ZC��>�Jz̚Yg(`IX��;Bu��w.�9�q<�&��&��곮��$,�L��5�:��'���w�!����kZ,�p(�gm�c{��Dd;2�Y�e�/�Nv�&��:��雠�	��k�w�8;r��W�D���hn�_eћ%�������֚`�J���~}.�Z;��S]��z�����\r�o.��TB_k��;zG���e��[�Ү�)��#�pS=�S�/�1M�x�u�jr��۶����izfB嶭RQd�"�hJk��JZ�66�#g�_h�d��-�Ժj�ܹ������G�j��v#���"�pd��.��W��|Z�.��U���u-���a;zN|�{���I�:�G�R�|حڎ�r�0&۝����Y��,��S��n!�'���R��}{\����pMK��m\;˰��SN��m7:�j"��]7f�O#�Ī�ƶ[�{JO�\�W%��h�� R޺�rX2i1f�3z�d��7�T7�/A�3��̬��a�cߥ��]Y'7[b9�kp���_U��+u��=+���'j{B����V[U.;<=��|o�s�=!B��t5v��릟3�)�j'�9pAv�����ܶ��o��*s����:3��#�,����+�1gowN6���a��0�AZFOiĹL�u�$��	'fD�I�ŀ������*0R�+1AVEĬD�)�Zh�QZ�TTb�m�T���l*��"�h镈�aY*��T��UE�X��5f&
�(�uj�1%��j���limEQDը�¢,F"ō�hV+CHT��.��+*� ��UDV)[�Q4U��+Pc�Et�f��2����#H�2ڢ�R�X+4��U�T��AU%j��e�[i�SVE[Z���YP������H��TKVR������:��`���3��e*#�UƉm��4���"Z�Hc�˘b��J�0F	u�c
�KE�Eb��Ɋ�J�m4�i���>�Z��UX�L��KGNZ�F+���b�v�f��{y33�V`Q�W�nt�v":�h��	Y;��Z� ������y�y��ɩ���w�bU��B �z��2��ʟ<}-[׸��.3z�i���{��v���羛��L�B�qΗ�D<WxN�{�������rx{P#����K��= �1�R�P}C!	�	��nS�
-`y�鉪ɻ�`m�/���j�oVJz��9�������Uޗ��uU�n:�x�kB:v�[����}�ۯ9I߂�ε�e_�"`�%�oz^�"v�t���k��]B��ݱ]*�[y��凥&����ˉ�x�;z�R�v+I�$6��tF����Ie�<�u{Xɧ��S�(uM�kmq�m�Wg��,~�Zw�X��E��R�����Y��]$m����U�t���v��*V�u���6
BJ�A�٥W&��ʈ19On*�#w�w���̦��sn�))PhO�ĭ�	���v\nKUa��YV/�̜������E�n�vw;,%�;%g-+;TV,�;��V[#�h�#��sk����h�6<p/N��a+��l��1)s��P��A��ٕ��d�p��u_<�-�y,ϐݎWn����(5�N�"��%Փ�����:���f3x;Ry��|]��u�.��f�ۚ�)QڟB�<s󩖱ݥ���E�u[o�AwT�$��lO�Qt�cx����Bom� .o�=Ih>�ވ�m#�L<���6�Qɱ�tX]7z��d�C˶vy�wFY��fK2<ѫ$eի�����9���l[˛M�=�\!��]w2�L�����̟B�Шݧ�u��%4�iꖞ�aꚉ�Q���.h��c:��8��x�nv9��b�`�I%���MI�Vb��N�L�I����ߞ��b���:5�,�\{C[8?L4HR��o"���[�h1#��2����M�ogn���Ux��Y4���i7�3�q
�`Z�D��v(jx&�+��GgZoe�n.�N#�\�%5�o�GU�,�:0��)+�V ݽ-Z�Ҥ&�<ny�ڑ9�͌��{�T���|�*�
��^�۵QXN�ue�K��o����cmPrZ�E�V��ܬB� ��	١q\������J�N���4�F/��s�e�4�N��s0gw-F[�<���olڽ���?�¼z�lJǆ�^�]����[��㇩"Tƈ/�	��Lw9J�I�0�+I�V�|ؙʱC��ئ���8z����%��aexN����*R��Jk�M	���7l�v� �ɧ�*ҿ'����x�}�B��73(��;�ܲ&r�c�f�\&���Z�S�i�Qb))W�؎����;;���2�*�i�����j\��wh��u˚����Nb���j,9��θ�����甖���.���E%0��e�Y�
�uMrL���ύ�nЇbs�h�*��U��B���}^l���O+-e{9��sh����A��I}=�::�7���[��im��eʷ��}�V���V�A�YkyA����y�מR�M	iE��<)� s$B���*�t����=��gWJ�u	�����M��?r�{ퟦ�v������I��s��Sʘ~)�,��t������Mܺ��n�J4�͂:ϯ�h�$������xߕwc"u-'Zϯf�dI�|�f�O&��RB��W|���Rt��R�`�٢V���\8V�{�f�6,���P﷾�
Y�-ǝ;���W����������g�?N�vv����^��z�G.S/q����gl,9�Vd�A��9�E���T�Z����zX}�g��ϟ2����_�{���Nf-�ɋ��}�H�u4�{���s^Z�un�+�/�;ns��Jb����n#s���Fgr��ο&�v뉏]@�*�}%j�vs"��]���䵉��3��y�Rv��~Zp� �0o�,�J�0�B�X�vBoST��cv��=�=���}�Î�oN����F������;���%��WWU<�����P*�fr�݃X���9�V����(!D��٘6.���l����6!���.{A��=w�eޭ��j�8�{N���W�w+"Z.��5w��rF�-��׾��E�¯riX-�v����nh����k�ڃU[|���vXsJ
TF�sn�5��K���QF��7:�\�8d�i%��<��Y�K��ppK��Hw�w�9�ʦ��_^�$L���wKHy.N�5���;\)pjjx{e+ń�j;�gk5ӭʽ��k�-���Z���]�z�ME�yqA9������X�&wVWM�hI\�ݫ6�u��ql����Ahl؅�4%<�WSW�S����:;7a��٬�wTזs2�t�cx�X�W�܈}�Ï��;J��v�o��"�[�y^�Y��w���5�D����E�׵��`�,Q��u5˘׆�m������r2�Ս�|��k�e�<��T'�k/!>����b�@�ٖw�1��ī9C�t�_�em��KA�7m��ʵ�\%
��`n��+7��/�	����b|��/�Aӌ�k1).Y��f\V��]�+���kglU���`�g��B��F�q5�JP�0fU���8�r�m��޾���cǗ� �}��:�f'1������m����caa\�6�);B)ϖwV�ظ��;Vn>��V�i>N:j��:�<�ҕC����^zRi>��v;N9�ƗW�Τ�R�1j�^���O�o�準�]���*�3�Z��ʾ{pw=����(:��@+�J�5����)��>t��p*�Ms�IX��Z��>2K���]7\,�)��O7>�#��V�4*�{;C�c��[{i3��[;�򫫹ꖝ�<�&^ft�!�pM�A�2y�=�i,��<�z��Xɧ���L«�:曧�a����N��������|���ޑW����U������ͭM���Vk��i_�����F�HH+�sȝ�{��8���:��:3h�]w�U�sm�))Q)�Е�N&�cn��-1�9a[������kɾ.�v����������AJ�иr�lZ�ke��ơ�\�Et�}���C5¥�S\�2�QtL`�����I��f
��l{���o���Ed��ym)�w9��QI����z�j���U�jkc���R���"̹V�Ƭ��V�z_XZÑ��g�X��������Nى�y�%��3�����2D+}r��N}�Z��D�d7��6�$��U\�1�]�<�\�x�/���_�T��1=q}Bo��&�{��'�حL%���Vl���j��)��w,q��W��Ң��5����Q��0�@����V���~�����}�%Jf��<� ��ݴ��5G���}���h���Ϲ�R�D+�3�:�{n�(e,$ΥG����R���V��V�u�I��VX�\�
u�L�xo��v��ƫ7��1�p��w4Mp!��m�UU�u9��C����>v�R�)�o�7��*�*���已��R�r6���.�	�P�v��u|��M��9\�(��O6���q�5gw������X)u�LwT�J�J��zZ�zWYQ�yo<Ή��r�=��=�"Tƈ/�	��Lw;�W�T�u_,�/�gE�Q)$ff�G&pt��[�v�=^^JKC�P�v~�k�E������܌��3s}�
ź�B�B��V���2�=��.'��d���z�[�ws�]����p�Aִ�̤��{N�))_��H��|�]`�y��k�����U�\���ŇKBu�[�}:%fu�Qx�N�0n�E��:��{\�����gt*]�49&XlL��v�Vu"8�aY	골�d̬���ݽ؎��A����wAik����e���ȧ�Wׯ�B���wz�ZlW���z
厦�X.�5����1��$̮��|蝽VO)˰%����vvIR.Kq�	�G�d̾9\2�A~�Tm(:�|۰�Y�o��]�@5�y{6M�psH�yj<�O?�J»%e0C�ا�Ku^�������5���
n:�ih�)����|�$ʗ-c��W{�xhJ�?)6~h<�5��iEL�����0��{���(���}�����8L��甎����=��?�?f�F�W��Fz�/M�qJ���[����쫙�~�=R���]=V#���2�g���,X���Z�-}��+J^&'-g��N����a�!��q<��S-�r��]n��{NP�&���q՞���ƪ�J�a��B}ؓr/�5w��o���_$���k''�y��֛���p���U0����w6���+}>��MJ�`̫"+^�O/t��(���.%�>X&�ע约���)��!1�8�&Զ�X{�1�O�J���vnN��(:�e��($˱�uo��e�ΖVd�ϩ<�4�h���ב�f0��9��^�`��{V�Mk֒`n+�3��m��<$ۈdǪ�p�:�r��V(Z�+ޠo�	�]�r����͸�[��\T�9��:��"f�v���4d�c���������j˦gj��
��1��RY@�]�9k��c&�8�{J���Ч�V,�qְ��m�q�z$O�-�x�6���V�{���4�ǣ�c�i�Ta��Wf�o{�����f��u�t�}��ܚV[��l�f�.�Q�Vn�SbsX���mڋQ)o�>ծjV���;�(nt3t�Ê�mS�LeMeEK�e�#����6����-W���Bܚ��#=�3b5\�H.b�r�c��vU4�����҃/�0W��`��m+�������t�/�U��U��ޟ���糫��\��(<BCi�<�Բ�3�3�k8������+O�Z�k2����s�V����k��r�Z}L��|�ǹ�DMgG<�>��0��*7��]=V:em�ζ�����f�'ꏚ>m�yZϭq�Nxq�gz���t��W���::�6�4~^��5��<��f�x�:��'.�Ѹ8r�\0X�*�{Z���GƘ����o�_fö��$�TT]:�9����gi�!�:�,VX�����s�]�5Ը�YǞY/f�}�TzYs;���]a�B�m�	[Sz-f��Sz]I���'4��ߗ����͟���:ng�+�cz�������8׏em�й�S�l1�0K䛗M�9}�,O�N��.T�Yue;|�c}x�J.��eΌ��Z1'�
�i�@9I�Q�ֵl��D�*�Cͥ��cs�w�1�^�iX�+7x��Xy�������r]��M����q���<q�;"4@=�KJ�;�����T�g=}���;�=$э��*#r�c[ؙ��uӰ��t�:+�! �>�(-��U.���q*X�ϵWSJ�M^�'˶ܸ�!�$�C����/,h,�v-��P��v�be�����w��w�:x\S�!R���
}4EQ���϶U����WP�ޭzϭ�:���`n�U^nq�Snk�+����љ.��x�;���L5x2�P�p�tΎI�m�(�}1� �!g���y�t�U������eM0�V�GIowi�}�A�38�su,�Tz�4e\�tp��Տ�r�bC��'���\WG�<K����s�e[i%�D�9������Y��N\j�)j4���ae�fJ��b�� �$"y�[*�v�)y��st�eAY��;�uӝf�����-0k@���7i��]C�vr�� �l�ٻ�n�=:�@%H�T uw����p�yb��̋�]v������N�tZ;�tR;��WX�ܸ��qWe�#��)�r���/l��h`Fi�b5 ��_:�Y�x*j$.㛐t��k;��nǘ��J���A�,����,�u���JBH��h��aZ�w(��FG��6�.T�%[t�#ۃ�	���b�j�D��̝���|�On�z��#525۵�(+Bز�W]����Qڒ��`}b�U����T�� �fWbh*��|+�h��w`�I���JT�
�)�نD�ù�g�.��E.�p��g���p�˧m;�O�uy��s1ҝJ��@Y����F�A=n�9[*'��r�ڨ�S�a���݅�e�-H.N��9���W(r�D�\:�+�ڗ�W����Q�5��^f�JYMN�&�ޒ��4n��:{zA�#-m5�R.� �{�yX�]m���[k{k����u�+�� ����uU�m�;�r���Zv���H��Aݎ�(9�݄�@rn���Dz�z5���Z�.���.�)p���85�b�ˡ����i�r�g動��lC����J1��G�x����/_r[�e�5��G�\��Z�y����nց�k�2X���ކ7�\�Z��o͋8�'[�O��จ�}��A���/k�K���w��{���ٙ��!&'GW���J���SY:�؀��[�����Q�)K�wu�%����&��6�l�9�)��yq�@�K���bH��#-��Cq�b	:�kQ�fS�YmvwV#�}gT��Ae�wQ�Hv�9ǰ��>��f�9����2fv�#Vy�ł]������*X��O�ùȬ�8�R&n�����l�8���`p�L�4�k�����mВ��L[���л+�����P���ֳ��F�n�vL6;ۅ��:ǔ��f\OwmF���k��P1͐����z��wV]	L*6Yu�ؗ�_S��^��0Woˠq2�jZ�v�Sua�K�+�wJ-b�
��n��ݥ��qЕ�B��ܾ�[Isa�ҧ��T�n���龙y��d��L���zVq� ��:�vL̡х�Je��78mWo�e�4�:A�ve)��߲8K*fcs��*��1�s��C�bt������y3V-���ak���2��$�p��HP �<��ۘ�f>�K��R�2��yC��R���\�r-WQ����
���
N��r�=�x�"'C�D�ST�A���/��浻�P�v氺�p�̧���O�	�C�6|��@ZԱQU)iV�b��0\A+ZYm>rEba[W,�B�X�Ub��0KV�����R��V**Zڃm�b����*�����c��c.F(�6���ڭƦ2�3���LL���*Q�b��!�r�̊���G)b����3*�u�¶�Z֨��X�[V��6ѭ�ZP[[Z�-�U�����b����q���kG*�m1��-�+Z�V�X�i�j�Ӭ�+�3-m���Q�8��#h���F+���2:�W.�qĮZ6�mlX*֊(�eU��YR��ej"*Kcj�f,0Q����,4�q�am*[J�KEj�������mE����iuq�s5��)W.ED[J�U�(6ֲ�iR��ldZ֔��e\JTmYVؠ�kjQb˘1��Yf�����o����m��}�um9��a=B�J�����L+39.�B����G%�<���x�)Y�n�+�V�
Fဵ����.l�u�?���ճr"�=崏-�MJ���k֘QA6"B΅ћ�T.w�=ġU�娱���[^9�!<˕olj�tx����5������$�6$��UnӚm	ifLߵ�����U��*�P��U��Q����b'��[����T��s=���4{̈́b�������Xq��V�'˥7�����]���Z|ʎ|�^$���)c��f�Ⰽa�0
�kn��=�9WS�.Uzt>�b/����S)XR�X	�X�N>��Of�ˀ�as��{��^��0}���k�u�^si	��56�u�+���L�S�܁T���e�t�(Mwk�[*Q#���LwT�J�)X�u�=-dn����ꬴ���SS�g���q�ִ��Z#|�X�Js�Ic�X�V����)��2��Nk�w\)�E���8yy#�JB|ZQ���3kz�^�n��/����aѵ���Z�������\�ڒe�;vjM�m���.�c���AW`צ�Jb��;x=�+��MB1��ӹ�FMs�tr#�]�J�i�o#�}{�MGܺ:�ܭ�ť���
KyoK��%�����H��ܭ>�rHw���ެ}�x�t��f��'7�����{�"�8/e'b�)��#NR�B&�c��"z��I]�ٺ�КW��Z�^e �8�iڋ���1;�����zn���3��R��}��
�sA�-�PN����\7P�v�e.wX�z��Տ"ÚpR����kһ2��3�.�I���wNL�ܵ���٭���s(s�5���ۘ[����/�d,��l�J�/�!*ͬ�-a��y�A�����`�AQ4�M�A���r���A��PX,�p�<+��	��w6�����KNd��~*�u���!k�] �QFkɫ&��24�"����މ9�u���zd�RV�oչD�8S����>�N>|W�U�s����c�,��G��,Z�hY���i��mIe��Ӷ*r�lT�qcd����3.uF戠�V8��v�á۳l�p&Azj!2���pV�(��<v}��WδP���I{�=`����#��i,BnteH�,6gW9ݳ�b|sڝ@�Åz�x�r#��@w
�t��d5�5��8at河�.L{�5����m�J�"�LΩۂ3.̚��L�=��q����Y�eZ܇��6x^:]f� F��	���x9 �A�f���Κ4^y`Xe
��U���J~lS���e��z�<����ỽ�L�e���狰;���<m7����M��n�+a���&���ar3���}�튤�	��v��T�Az`�s�ӕ~f��7��(�I� M_��s�����̅)=8��{bT%D���N3\�l=�
-�PH3f���qL͆ޚ�I��N�[�#}K366���`Q��*e�9iV���`�3��IO���	{v�Lݚ5�CiԾ9|�5v�D��	{B$��A��>����z^z[�Y�{�'CO-�|өnej�h�UN���¥�JcOh�[1��g'����av�lyP�MB5*���5v����tb��dF(���|\S��Sb�E��������A?I�)��z�J60�TԿL\ݎԄLݘ����v8��n�����:��$@���¥rS�M(r�Tt�{��t<�����H����n�ר�F'�G8�A9d�(�,鋃��yʳ^g�G�w̮��3�� W9;(Rd�ں�d�%�w9���r���Qް@���ьKmP6�`�s\'|��dr��,��y���Ou�ys��M��>�۶`�dvɖ��\�C_>��`n��U��.S3�pw��@h9{��%�[٣z�n#&��s�������_nr��R���'������,(��p>꜊��q.�z�����[y�w�2X�����O�J�W�	�<��h�t~s+�Q����3|[���"�>G�vu��SzhzGP3����N*����4�z�����8��W6�f�i��0�ؤ��S�[f��yW-W� �����NH9!!�^�L��&�:z۽��vȳ6��n�����+k�9��$�����Ӟֺ�m�d��'k>M��u�z�{$�yS�{��:(h8C$�s��ּ��.���]����cj8�F�GJ)���ǮN�,W��{��*Hb`f�4�M8�A�4#G���7�Q�MP*�ڸ�ށh.�Ks�3�v��Ƀa�vY��8�	)�Kر�;�s���iϓJÑO*��뜃��=Y[0r���uds���� �9J,TϹ��z��N0�>v��A�u�]��13ub��=�t�o�2��q�pAJ�Gx�I����$#"�֐��5ԸM����w���s:��2 �2%:��9\'�4�_ܸ��9�]�2��Ð��g/P�u��t��}F�jE7M+bv��M��z0녹�OL�;�"F�.��%�22��������p����k.F�uGOX��f�*j�s�b|-2����O�q��7<�q��v̛cj����[�	�ݔ功pE�}�r��}�3j&r�ǻ`��9;J3��:�YÆ��zr]e��.	
����N�W_���Q�����f���䁗�u�1�G*a8}ÑjU� �V8�UX]FAK""vn��n���b��ߋ�	�O>������̕~͍���wK�qC2�@.�n�N�'��U��@@;Ps=L�P������n��aX�;�61ϔGv��A<`���U��B'l��2��X4ڹ���vB�20���H��z�Si
�zR֤Z�zx�,y_�n��2n�@R�ս���v��K���e5�ʡ.����i�޴E"�=�f��VUj�*����wخ��j��h<[�����f���t���H�o�;\��g��WQ��ȍs�_>��D�x(��(�&��Μ8id��a��;�[�8�j��U�"����m��v�z��� >��@6;����(NXM�F���Ӭ�.ak��Q9g�*�}um겱{���Q�B{j����b�V��uqIf���̒7V>�&j�YPދ�:�M���OK����O������l�<:�F�=�16��N���^������i����N�t�T�򹗽f��-��^�EI�����7w�1ip�'�5�P����\q�R�Ga�<�
��
�\�����+%f-}�iљ��0齎P��}L�%P�^�A!\�-�>mxw>hVR[�d��;ц
�]���bf�NE��THmR/�ZQ�t�k�D*#A�C�
�D�hL�~���#{E�y9�5�����e�<༐��*��9K�=�}���>[�V����{/GX-ݣ��4�]]��(�Yr��U*z��	�;mP�@�J-=�0��$��4Ў�*t�4$2��vl���+�oO�Bt�`�8CQ��2/�=)E�T��&��MԈK�3�B}�m�uL;�C]�zv�`�����چY[����{z߼oV�|k��Hz�";�Y�&�]�YY�rU�Q&d<Iv�2�s�����f��dF0z@��л~Ma�7�<̪�k!�ت;�o� �L��JEUu�e��c,���u]@N
��'L��A�신{��Y�+��tXh�]�Z����h{�s�V��\],}g��)k��}4PU�\J
+���D�i�u�7.N�A��qTe��Y�܋q�M�eXܝ+�x{����=�9\.�;�gb��J��6�/da�v�a�Ggr��UI�y�Su�u��ZLޝ��Gg���M@�0]�A�P7W#���셮It��QFkɫ&�ܨĩ����
i�,T�;~�l����Wr�����AV�w��̕��?�����U�s�r/�Θ92��ȉQ���b��n�dT�����/ENTm�S�Dm�� ]=���S\�a�s�0'4CԡW�z���P��n̈{�vا|!2�����v%�!��\��ZA�|�o'���zm�mv5j�������.,����:gb�GI�
���^HU�@n�-�v]/�0eٮ(yǷ	reY�0M��!�ܲ�Ӿ/qǏ�ݞ��&�$��R#%o��;��j�V�0�u�1�<�#l�#mQ�ct�1��G1�m9W�Tu�PNDu)F"A� &��=�ȗݽ�G�U�v�TM����p$Ⱦ�-�k��k�����ac�ZE��1�kmO���R�wD���D�"|G7"b99�ZU��t�U�l�y�_Cj'���s��t�̈Qӱ~���r���:��6�m���^1�} #�/��y�n�gE�#�^�r�QFQ�]��r8�K�]fr�<��F��fF���b#��Ș���/����h7Iِ�5�������jzuniwOu=�v��%I�׻u����k�@��5������z�^3L�\����kd�V5���M�����:y�rP��˻�ލ�G+��
-{$�2��q�cw	38�=&�t�ܵg�{��ׂ��{�X����n�Ynݦ`�I�,�N�\9��-D�%fA1ѥ�I[ �};ԥ9&�ldMn����OBnx�E�$��4p7T���P>�>:����yp���_wq��������E���S�[���#0X�w���Ő�p!��\��mx)��[7[�{żzfs�i�6hKU�s�=���H�Yӄ+�s���K�X8Q���H�n}p.�����%����~�r���gó�+U��Ŀ#�n��@��W8��r^J�E��˒9f*h�E`�%�+���Y��5�K�D���Y�l%�vw���Rz�8G�Ԣ�����s~�+)���_C\�R�i,CE ��b�k����xTW+C'��Q�^�p�0���/2��J�����<��#a��ӃZ��뜈@�n#H��$F��m\s�|�WWpzbM����k 2L��IçtN]q�.������ ��g�^3Z�.��n�Ul,QR���u�k�l-�����y�T�tzm)��
���T�q�{vtb���{²�u��|��rq��\�n��ݍKXKW	ձ�#}v2<��u�|��/��|:ڛ�ִ���S�=[̾).h�Yp�f��x����հ����kM�Z8��DT��`��\n���#�:	Cu(��M�"_yf��5$�w�Zbcn�EP�
4����T�j`4�#hŏ��wi��ș�ؙ�F)�'�U�/v�Ou�A����	�����S>�)X
a8���b*$�t�ik���K}��Rc���1�ãE?{]xT�u'�{�B�Zۄ���)yB��Ha��a%J*��^�&��z���oVy�/#8'\z�;�d�لt���z��0�T.w�̠�-�KRܛ�Ў��7k�lrv�`�9��p��ޜ�Yl�\)�JE.����Z�o��$��&X<�]N�n�!���6WA�v.��9��{�k��n���;����㗾�#X#>}�P��Ӟ.a�a�+b��"��&��S����Y���=���aA�������GlE^`���_].^�.��n�v�2��宭��l�w���(���'׋�&ڰk�+��o���D>N.�	��ͧ6�9{Yq��0N9m� kE('a���h2u�1z�BP�/��F!�O���飆u���t\VXY�I{�o'��7�n�o%9,�k�T�����D�gue$�r�U�����e#�NCO]��9��=ݬ�JWm�;��1ʈS/��;F%Ս�%7ҸTf9^mu��ΉO+�i5��in乥��r�Md��R�avC��F���7��� ���ט֎׬���㾹��;g�#��=x�;��Y{*�'gq��1�W3vC�#��;g�������6�K8�{a`�Æ�Y/fF�˺/v.�k:�wH�C�t��3(��1��T��+��@6;��
��F�'��I���.�r�.xB��k��v��N�^���ix�]��dO�z�+�(r�Y4.�f+k�S��z���k��}��q�&��]���Kt�ׇuΌ}�uͫinj�seY�7>{�S���j�x�V�iۦ���@�D+N�[�$-~���Z�9�����\$k_�o��wL��r^ȱ�IE�q����8���+��i�DMf����Wv^v\�>*s�L�5�
�pB�q��;b��h�J-=�0��%L���V�Qְ��$� &oh1���$��z���%p��!�dZv�N{�Ҧc ��Ө��KZ8��4�m��co5SC�%�H�;M�P�C_3{u8��᎞oq/�3��j�;p��1�(l{�k\���W��r�+�9��+��5nV�]>c�gZ<.+��U�׳.Έ�-Y�s�|���Wm�[��`�ȭ�nRI.�<gs��B��K�G���'z����ꚱPIJ�H���&���f7�������n�Yu/aH���c6�p���V��5o���ڴl�0u�v�% mc�tt�[��iu��W[Kb����p�S�{L����O5��j��ˣ�&�I4�����0�:�es��*e�k�}o#{/�NBb�7W{M��D8�@�����s6Q�:΋<3�丯��)c籢�huQc���<Βe_*t�#PX��ה�R��v-n�S�X	R�t+f�lK�f���W^�5h��_,	P��V��vZ�Np��e��j�=h��S'�[Pj�
����`a[[�[;�(�8o��e^m�gh�,�s�x�'f�rRż1�����s�M�8�'����5��<�e��_8r��Oa�2^�1��lv�!.�P��ů��ӏ����ȄЕ˫��4a������t�8�tR�X��Q���kLR8�	B����ެ��.�'}�v퍂_\�����,���6Y�6f>�����Mb�mc�V���=��jfs������":�a����L#��A�F�f���
��G�p������m�$�F�X�wJ�Z&T�J�7��q��k9jN&���V��{z+��Q,״�%��%������h���c�<<gwǃx�ozo%���6&ewa
R]��晹K7i.ߞ|�)��Ť$�O^.
�b�mL�4 �1Ɣ�δ����,�d��8��F��{�؊�c9/�l�C��w=��V2Ë��OA}:���ʻ;`�ɘ�Ɏ%m̏�quш��f2��o���%ī�Ӳ�q��A��9����]��V�	�v��&pqh�&.��!f0���fֵ2��K�<�`����4,�y��(ȩ%���7w�Ǵ\���$ih��`���ԇ �xc�HJ�l���y9�yKg�xө1vS�5�H yu��e��T���8��Lǻ}w�}>6��9'*|�U÷%Z^\��9l3GPh��S�}���*Q�� ,vj�ؚ̣}b}ϫ#[ռ
+\~�wFo��súi_R�%#}Co��f4,Us�'V�d�o*�U{t�+��8�q1�-lP�RR����/�@/l
U��r��!z�[R�x�OxEQ�����w9������S����v]>������ٹt�#�yi��w�^fV2�S*�Kٷ�QcB�P��޴�gR���XT��ЋqP;\v�RɝW��%�ؾ=X�¦�8w{-�y�����M�=��p���u������W<�v�YFu[j������9�^\=�&7���qBW|�%�VޔG�nki�T(j(@�?�4��³T���-�ee���F"յ�KQ��ň�Eb�j�F�[e
R�&eF�h�\��Z1Ubbc-Lk�
ʋ"ŵJ�j�mh���`̸j���B���UE��Z�ETB�b%�WM��Q�cG)��m�"ŶZ�Ŋ�.e�Z%��ҵ��FQm����e����T��[�զe�F����U+j�S--[j����,��Q���ʵe.\2���hֵZ�J[q��4��Km)[j��[T*��X��+lQkmkA���iKb�	q��,U�fZ�J�hi��k*�33M]YVJ+)i.�&[+Z��J��dqR���"��X�2�e�-�jUJ�[DL)D�t�\��������*�Ua�
5��m.�LS-t��R��0�Yr���Ū�h��*�MS0�Zѵ��f���Z��Q���+�J	���Q�1][�����$ @!��!?���&&A�=vG����o);Md�U:��s�ǽ��B���5Y ���e��ޏe���ѼC:����X�:�8��.}���(�;Ǽ��N�
�f ���D}"��}�0U]l���=~9�o¯���qK��=�5Vjc�6F���ָ��	5�0R�;qS�&��hd]�)�%��:�16')ڤ�j�{�<���C�+�Ma����q-!���~�ەO�(7����*F�dgn��b�r�ǻ|C6ҫ��ਚ:d�T �C팰lt��1ep�6`Inub=�+��bw5�v��4�2��{h<�7W!�:�8-tK�"J3��&��s+X���P)��XQM+ǝ�iC�����H�0ײ9�em�>����s�#�c��Հ��7YC���[������#a�1z��V=)�g ���6��t���uMr��̹�
��+;�����n�%���1�C��F���-(*S�[H�%���>3��XU|�Ee�[�����a)��Z�If�~2��Zn���5Ιز,��zB�g`)s$`�$�dڲ&��5�o!
v���;��Od&�c�e߃�|X<l�MmQ��r	�t��l#W�Gn�+�Y���4���
�q��і��`F���e�b�b��[�:񕇋����Q.p�/3�_�%)�&�)�Ѵ�Zֳ�\�aOe��+w��-��Z���ڪ��~Á5/��'#�]vg'�p���Gh��LC�]9(���ڇQ��Ι(�]�}0Q��7~r�̨�<�����b��K����^g��4���p����^8�O��.��
:�u�ʜ>��-E8�"5�}��W��+�[zd�cpōC]�D�rs�ҭ7J8�r��tf�$v�<���!O���37a��b�xw�@X� ���%�{�M�#�/��y-߇���/�9���.��y��d:;5,[�DT��pX�Q�A)	�y�2���]���T�������{��Y��1{Z���D<0,����sn�R���qD�J
�:py0�z[��:��5�m]E�(.C����őI��tɡ���C#B��S~�O;��g��u�i�3.;�����Pˠȡ����$��q��IiD���Ld�D>����)w[�`�.�ٳ@J�Ӹ*^C7�#�8B�u[a��8P t`Y�ȣ��K@�U���欷)}���|-�8���Y,��~ߚ%]s+�V�b�;����Ӕ�v݃lN�/U)a��ᖽF3�*{���!�J���m�v��AM�< ݼ�nvj:h�V�NL�Cޱ@��Fh�1u�J�y�,E��E��gvnk�I������ �Wt� ���B�=��m�Z�T��e�+�L\�"M7��|4�PU�{�F�J�:k�S��`�9�Ig��[��򅧻<�r%t`��m��^�.}4Z���8�̜� ��rB4}����m�D�j����A�_�VmK���0�ڱ7�F�緧Zڣ���0S�δ%�Sѻ���X�)�c!��A}�B�D��T�:���4��.��t_���iӑ9�=1��_cg��LD?ENfe�.�!�V)��:�O��i�n�!�n�"s���~k�u'�p����X�3�����s�LAr`4��FJ�bǌ���ƶV�L��﷛mۂ�zg�W]x��:���-4m�L�?�����ҟu��E�� ���.�p�<U����[Ύ��<E �PdX�ӕ,���LI���7V^Hu��YqU��3�R��Oeѡ��|��+�Nt�wlɰ&6�N})��AؕP����үN��ԯAf�$-���@rv�`�9��p��zpK��p��! ��dV��9��D�j�e�orK={��oהo�7=p$pst㭁��n��2���u�OfW(op<�]bqp���{�X*����mv�[u��u���$gj)=rHG@tn��T1����zA�]��W�յOu�&��Na]���ac�:K��o�I����|>�y�
�W�)c����x]q`��e*����u{rCTM��TG���n�N���51�[�EgD5�p��lo��w��2���go�Y��.�Q�5`o�gi��r=������</3d��\�%��]�k���{��i����-*@i\�~���p��$w�ٟ3�|ח�=�7;g�R���/�;�s�D�y^R��K]�tit�\��k%�B��a&��}�z�oydT�L���TE���P�A�ŎWL�j��Px�<�NL^�ӱ5.jq�J��}7��9_�2r:-�Q�V�A�}����Ćh{�J-Fy7�S�9w��䤾�;;�.+ԫ�l,��r�Xz�R�:�@}���P�;��h�o�V'ݖ��5�mn�.�D�@�Ρ����/�d��GT
��旎�O��c��V�����J�ZO���QS��ms��H�x�Bp���
"$����ׄ��D�2�x"���b6�%pm��V#�M����J���t�\ C9+�2��Ҽ���-^/hx�����N��~~Ig�2��S�&f
��c19��gTJ����ȼ�}HNԶ�`��`]F�+�a_�3;��R+�e�;����vƧ��m)��%%3�4�'�l���'z|��Qk�AQ!5H��ZQ�8GTD-�	}!%�r��.�\�j�F"4�j���WL���K��IU�����/�dB>ۅL����x�sWBAb9P4zR�0F�����S�7S�r)�,��P����ѹ�!�C-�����cd�F���N{�IXJ��ƽ�;�}��Mv����ب���˾}j��j����K�= �� U0R�$�Ϥ\�:�}p�K�[)�)���Y��b9�cI�7F�A��~��us�O<k�R�2�";��6�>��5��ʣ��ɑE^��ي��7'X�Q&�T�p��B�75; �=�FW+X95�����!K�E���zm�ʋ�Q�E��X������,�D�tɠ�>}�tt��,�6�w�]���9�=�ԖfZ�}h�}������(���yݑ~Z�W��QFh&��jhĪ�%��7H�jM��ޡ `�PZ1ň��@Oe3�����2��?D}�ח��~Ŀ<��&�?nb\eF�V_i��li΂'��_ܽ���|���Ԃ�ܾ~��s�d�Tq��R��_r�9�NyF��S9g��&�d�,vlg9��%W�;���JÃ��8]a���{��z��d�k'JރM��44]%e]�3��(�����&�5L��*�c�}���~�%:�{銓����r}���G������C�V�����$��}P�Fⁱ�^��j�U~��X%q�m�U�G»)(����8�z�A���/�:�&%Y�D�Α�2����ɺӧ��t�ődt������
��TFu�f��{�SCZɝ��'u�������	��.ç|X<l���]�r	x��f��Ì�ys�������T��D�@�CQF�O#<�`��1�nÕ~f��_I����`�bc(е�Ѯ���C�Ԙ��J���Gq䤎7J��}�_Cp6�Ѕ-�XZ���g��Oe��Z�8���J�Bg��D�RK{��s�>%��w���t�q}�X�ט[Y��EU��C�؛��n19��!�J[Nό%�c��l#���z]��$�Ft���U��1�<Lã/�U��G4s<+[�4�Ѧ���9��]B,�Dm�$S��u5��I��;"�=�r����D<�^N�X��Sb�E�(����Oo����u,DtЮ��=c/i�Řְ���hLI�Y��Kwxx0����4�v-7�@�eL�&��#]����S���^~�u)k�(>�*��fQ1\��!
�٩��}lk�f┧1ʢU|var��>�2����f>q��p�1����ȅ76���z��~9��ߺx�(&�0��� ٠�PdZ��R3}��=�c����i�^12p�ԿC�5=զ�T�s*B#3^�X�zO'O8�ͻ��G�u{%)�"���N\&�Y>R�5�z�͚�էf�=�#tY{��F �X.�;"�jN��<[��Nٓ��2���7�9Q�eފ�G>���+_ob�/Қ%]q�0/
DTT��k�uWr/ <��0>�d��;]Ҽ�-�+t�d���sWc;.9Nḑ\�`���-�Y�U7�C�8�h����:F�L�Ф�HF��'�L����D����y�;>���Rf�G7�=���:w���gسɼ�/�V���G��"C�{��Xɹ��}�z4j_�R�q��9>�Y)�"Or�p���k�]q�.�E�ǖ{l���N��A>7`�z5�F��3�A����%���k'���6�6�{�豨�Y���:�����΂_���Byܤ�1�X�@�v<���}~����m�2Q>��*T��W^:=��A���ު�h_N���|s_@L����E�(�3
ݺ�V����@xS�I\xSY)�Y�s,*��+� 
�i�툒�\j:*	�t�ښ��������͚�NW9h�̌��r��&��'m� �pN��{pZo��fV�k�rS�-�qݻ����:��f<�Am�f`9:7O)��9W�OR�����}��j'��y��ч9�U��vJ��ݒ����8��OvHX��1�K<�RdFk�w6y��.kn����x{��=˂�0����ݳ&���#iϡ�8 ��@��"˵����U�b�����$-���C���=s��͛;��ޘst�.,�0Ff,�74�&����B`d���UƮ�tm�d���lP\�9��r��y�x�~��4W��朞ś8�����U�#VQf����\Vz��i�7%l^�"��'*�6��oc�R��%$;	g׋�{�*�F�[�c���&W�mټ��gÇ�t�u�����b��a>
f2�-)�U+�7�|���J�iT����vB�20�8̂d�4Rqo���{�����;���+H���z��\�(<�)MX'Z[�F�Fp+���[[�9a�ޮ���i�Ŕ�4C��������F�酱~�t�=�WG�^x�=i�l� "�(����V��#s��C�+���/��D%���q�
*�q���(J+[����V��ٵ]y׮\�� �׏�- �ț��J��vN�ǩe�ĝi8!�s�c��A�u�r����`-[�Ͱ��Z7�s������7�5fN�Fp�5�Fŵ*=
ܨ3C<��L^��.��$3�
-Gy7�sY]rE�m=w.��=�cً1*��ͯ�,��ܧ >�<=���lʼ�v�_^�{T���KZ���ww��㨚3�'\���^:%>@V�����l_j����9���ș�dD��FB�jۦ�çH�t_G�..�>=!��2B53=л'�y�ڽ�7[̮]�´;���;�-ϭ閣09D�5H��ZQ�t�q�O:*��eҊp}�~��MkX�}Q#�zft���k`R͝�9/d^9%Q��{�߆��	�"��i�:e�܅O߄�$0g�{@��N.�H����q*-�g����A}sKV�.}Q{w��g(�/N������m����OUF59�%tRޮ"�:J2�D�ՙ�gU����]EX6���;j���d�F�
��L��|;
���w)���ƾ��U:�C*k*6ͳ�؆�ޅ��y<�+�H=H��Ad.������j?{��g�V��e�4�c��CE
2az�1�Ւd��\z-�If�߮�"7\\X>������*.��ә��Zä߰o��zr[襈�����FN��:xё��k��˭U
/��)�w�s��\�#Êg5�7��5�i�\�!3z��p��dN^�q���nLI�rT�p���Oy5����O3>�k!��=.�͗�buw��������`��~�#�����Jj��N
�NY-H���c,8�{
3�z'��X�����<e�5�s"O�}�Eur�;��%�t(�4��n����9ۍ��ۇ����*��w�A�2����]o�-���;;��2����c�	����t�W��M�>\�"�Ȋs�Tc�;�c����D�犊|�F�'%b����
f���yo5cvbj�f�gg\g��"�*���S����B�Rq�l��6F��{yJww�c�ǙAM�Y/2� �.r8*�mΙqg�ɻ��5Ιز,�U�fvc/�z)���9>�|�WWqC��w�dUc:��V�M�N�aӾ/qW,���G*��I���
�zZnp�p�n�ب��T0B�2Q���Ls�ל��6������9�WhZө11�J���b$(�.���Q��(� ���n3\�o�hB���6)nGsE{|-���=S3v��`Wp�+�V�/�KT
��̥��s��yE.�Y�o��t��ީ۷�D
J&x3��:�C�U�{��S�54�
3;U���� ��Rn��{CH#���֛CX���|��N�R�9�q�=� v��ե�����lԺ�z����Uo)�p�t��O5˥���X�(V �9	w�R 1(2��7GNU�R����o��E;����u]jt�l�@��E�\@�T�H�
pC;�0e�DK�ݩ��'9|4WtV;�"v�Ԡ*V�.N�������7�>}ʷ�Z;v�}�T��WJV���;X\�v��6NeBŞV��8�c9u���2� ��N�ƻ\�z����δ�l;f��ǆ��e�[������p��:�["�P�^��c*weLȔ�m�|�9WD*��k�3��Z��.�iשf�R�h��
X��̾����Y�`���n�eHv���9�y���P���zc����SI���ȳ.N�[��m���!Zz,� wk*��tKy�S�S��Le7�_Z �����ՄKkS*�b`.����0 ��r��[\��.���y�]�Ku����9#��R�u^^X[Vґ� T����;Gzk�;�r8�kP�'P��ãh��{++���(��_NL��W���ʹ]
GO^ѡokd'c�3)\�\�sB=| 0��h.C��M��m�N��!���;h�!KKn�B�"ޭ�FX�(g`�#$�n�h��R��ޥۆ��IZh�L^>�|OW^���������R�<]_b�Y�۝F���S�R�g�<)�*\ͦՉ�����:��i7l�}ܧ\���O�:˽���n��f��\��U釹)��V����-x���oJ�zībm���_^[�1c�!�׌�tBY�.Z�t�-b]��m��N�՗'3�q���K��m�}9c�|9ǃ$�T覲bս�Ev;\9})�Ph&fV�WF0�����Ft�4�����@&:r�S{:�툆�.��7��ye�QY;�;kkki�l���\���U��8��n \���Z�H�yu��ŏ*�Iս�J�n�L�!{�	���x�(�W@��Y��uM�3���s_<����tf�5-���(xn:&����e�k�0���v�2��?Y��S�u$���V�{��M�*����VP���Z���h������VpA��bl\& E��ePꀮ��e
��ś�׼7�(��5��;�
pw5F���ռ����p'G��Ֆ[�|΋��Y�c�O٫v�I�P@�<K{��؊����v$|��e`��|����N��X[X�+@����j6�W\Ev����Ǫ�3�n�-��ȇ�����օw�p��8�p�-m��P&��@��9��h/�қ�+�9�Gw9Xs�*�f(�����w�8u���ԎJ���wu*�SX�Z�B��)3]R���Kn��Z,��&L��ڒ�[Zٖ�+�D�B��(��TiJѩ�fU��Wf��f4��rբ[R�T�Z�*��P�t�\R�Z%*fTp�M2�R�
R���[��j%�T���ijʥE�K`�Zښ�e�i[t�2���+
��l�̘��i�ijTl��k+.f#T���fKZ�J�[--b�Kk`�&)�S-Z��Db�0�+Zܦ8�D���8i�R�J�ZT�0���%A1���0ȩ������DT2��Vښʢ�kM\��iS1�̦���X�*�YTQp�t��[d�ljQ�[D����q�":J�:ȵm-�i*�#kQ��e+DQ*�5�+Y�Q"��E*\�b��"*86�c-m3*,U1���A��\%���\e���#��Z6��E�����H>�������A>�[��\��#�SwS�4΢�;����j���\;4�ݓ�E��py�V/����U{W2�bq�M��:G���\*���ҧXb�o�*$�QM�D��݅��~ݛ~H'Lt�4�ձ��TD����I"E>v&���j0�6 �	)h�'d�Phxǹ���:ޜ�_1<�z�_��%�Nc�Kvxx]0��ޕo�sA�3�ձJcOh�[	��2x=���3���gܵC<�#�OKg���*j-ʈlʯ'vϮہaM�u�BO)^�Ï�[�]�d���6�	�ξ�
�OE�q���&���A�A��Ȓ0���-E^˾ӳޡ#����y,Z�x�!�ʐ��׶J��x��k��$�����)�䳀�o
#�x!��]�=^;6hK�ӹꕐ��9�8B����*������k'+��a)ɻ��U@�DןuNEUϙ�1rX9^�B��aq��b��'������m��n}W0^�o���q:��8��io�p��3"
�dm<��&�tm̛�Z�F�]��դ�[�,�U7�R9}_'�8��2o|��HD�:Qyz�ۻ�$�>/6Z��M�Z���0�X���o�.�z���]����e^xL/�^=�Z� :������Kg2"�3�KC�},c�|)vD;V�+.�N�3��;o�s��������\Tl�AoU�:��q(3sP�a�>�&�RF.}�ӕ�Q�V�v��ڤ=fo�tA�r�9���%~�ea~ֺ��GS�dp�p�r��o�JIĺ)�Q,�Q��,��AC "Or���ya�x�ۣ���u�n��(˙�r��b�2���r���z��1�Ov(b�qz��k�>G�n,%�
Wx��E�O���Ҽuޛ�]���<2N�@�� �9�Ґ�4�
)���N�합�2���<�*.8����w˫HU�Xx0Ŧ�۶��GF�_h�8c"�A�Fc.;ӎ�p0�Y箸��:;.8��G=9P�����D�,Mq�q^��DORI~�7��,H�7δ���k��a{����v̛P�q�p,���ї��O�z���w��� ���#
����;l'IB�:�p᠝��4�ޝ�7j�����@�~_�����]�$�o�$.R��臻��l�d�R|�ru1X&Fl3��s6�4*�.�}��?��wM{N���پhW�{���ʄ]�G���83�ˡ����Ar{G��`s{M��@���-��q%Ǳ��mWee�c�_*"���YOU��osD}b�i�y�N;�v����z��-Jw�� �:�z��N'����vn��b����Z
�/D���A���z�we��0�_���4zX-��z#�C�au�7!�:l�>5��@Q�ۺù��5�&�)��19�q���x�;�7�|�+��i�`���hgڨCv@��s䭛�p�A{�y��8���>�g�tL>�S���;�s�D���M`&�[�F����;�E#|��:�z�'b���i�*]��e��V��F�L-�U,�M]�k˚�Fa���֎Q�vC�N�5VA�PW$�}G�:-��B�)�JQ���B��̀�K:���gy��'V�aS�5۳��Q�!�u�y�����~ܪ��W�r�U�a�Ir.h��UC��U������e��jj�_���7P�;B�8
�ѥ�S�h�=�w4#c�ք)�9�{�l�P��鸰��"��΄�.B��=!�+��_�j�̿{��9k*cN������>���Q�P�O�*����k�i��]U�G';�_E��w&�Z��cn�H.��4�̳��[ ��l��%�pJ�}d�}v�_�,�^�БS��q�q��(5�3%m�(Z�/�[�Q�^(m��~+�/n���%�6��,�U�z�{,{��Q��f�[Gjz�]��lB�W�kU�fJ�����+�e͎��_F�2�ΨƦ���ɒ�g��u���f�ObF�E�w g,�Da��q#A�BT)D�#N�b�+V8��n�@�t:쮉��j�s������Dz�_�U'�f��$�@Д��1��T�;�z�����=�'��Q5՝\����:��!��=)E�T� ��h�� Uod,Pk�<��c26g���nB�����&eY��2��.G�ÛQa;�`75�9�BM{�`�fv��,����(��c]��<｜���[֠�8���J�#�$�%N!�r��B���S��GQ�eT�P�m�̺���6&���PζC6Uu8*'�tɯ5B�>����U��Z�^]�L�����GH�1� ���Yn�B�o;�/�]�Ȓ���j�S["uu�N�P��&�T�c����(=�X�~mTa�g|]��\�~��
�{�z�;I`\��=OQ(�8��T�8��0r�C����x�㸴3[��?<�����ohL�5��Ar��h̘���:��!b�q��0�	\l��5��/
��h���Z$��"���+Gi�H;f�vy��{��-��c�]����#UdP�j*�h�%�6˿�e��q����ދ/�ƯE����W|��\U3���Z����s�}��b�����I'S�{��^dB�*,9���[!�W���̓��-�8��"-���:�,a6�iGK�#U6�L��֛�<s��L�_��8tL�j����V��O�xŎ�h���b�R��}V[*�X��r0;�]�:wŃ�����7lFL��Y�ݦz�!�#TK��ath�b�(� ��g�Ls��r�̛wNm�u�1�)JI%R�5ݚX����5�1�����d�7Iht��Ÿ�k��h�n��n�s��*y�n��j|#����k��k��fb[-�6b0�08��)S<��Zz�lr؇��\.�"z�Ş`oPG�0k�E>t'e･}��R��7F����=�yy�����dL���;;=�S�Y���Gq:k�����ЧJ�H!k�f�_PЫ=���u��}�l��h`����ǝ{�5�7J!�e'T϶ۀ������6㩵ݝ��,z$�N߾
�5^<9ϰӫ����j5��Ő��0�.�4!�A���E՘����繓�N��T%�^�@�����^
���Pˠ������$��,<�$*�v,K���U0�� �2�T��WU�Kgf/}J@�ѹ��{�C������E.±���\�O��:�C�,�[�tl���\,��!ɭu���0�}�qr�sv���3��ei���v��M�'sGO;Ԓ��[\T:^��:�}[�ڮ9ۼB���G�p!����Ƽ�P;6k����
����9�8B'��Y9���r�7W�a��@���7ɪ&��Ȫ�O��n�+�
^F���gs���p�Ǫ�u^6כ&��΅�/m��"x��}Х�U����^$.zW��-.�A�ߺ�M;���1;6c2Y;��*fFP�a��|�<��_[o2�쫴o�1�<OYi{��2 i�P�q�8�L��� �k�0ny�q����o<�畄�t)	5�c�����bz+'X8*N
��z2���( k "L�*Nhya��*��Fu�$�S���s�]����Tn\���|�F50.�~kS�%V��z�*�te�^��<�6������WYh�*��1��q�;���%��1aM�ϣϩ�+A��[~`�={&y�h m����t\q܍!M+
��/�d0 ������$Ւ��k�5�ӍU��P�L���I�P�a�|���'�<j{�W5��IǗ=ؠ�:��*ﮂ�4�jn��.�֨���br������)=�Ɗ�]sN[�ܻM��k�e�@�r�I���J{g��$NYSW�kK�7��ȇ��|8WN�u�7�6����զ��R�`�s�MqU������3��;M�d��nEײmv�Z�J�x �;+�Ѐ���֑p�v{Ycp'\z���7鍨E�M�_F>���m�����(yb�-� �/����l'KM:+t�:tЋ�1q��wZ9��VٺD�G0��)�"	�:�W�R�6��!��ؠ�T����s��s�59��5�1u|�#��˨i��qU�3w1��Tyg�G�lfZ�:Sՠ�(]�̶T]��!�ݡ&���Qm��/@��O9��8TP:l̎�>��M6h��q	�؁���Գ�5��X�;�61ϔE',iP-uI}2��1\�f�H��2�|w��>�pQ���|�r��Z�YZGYs|e���O+�h&�M-ܣY.`��82���b�v��D��1�N�T�!vMo��('�t�4WL�j��EzUa��}��=[�/�X��Xw��h���82c�L�v�q�.l�{,��8ut�s۾�I"�����*�v�b{bU>�`�f������ƪ��i��;y���?CPC���-��ёj7h�b�Q�P��ƈ[����Q&�Һ��!^�;�G)ѓ�v���o>���#�}��6Ṇu�6��.*�α�+�s��nXK������'nW�Y��;�D},�������]z�V5��h9�v3��_���FSD"�p55C���V�\d`��Xz4�tv�־�x���Y���Ngf�	��>�A�;���4��	Ӥ|�/��rȗ*DI���[��߻���ݱZ=I-�)�����tER[�=0�Zr
�Ԣ��B�*���]K����}G<fz�3 �+��r���C53<yҥ�8B�g{���/��_G)Z���۽=����&�y�gb��JDH�f�k��Qb�M+���#���v/扳%I�{��kn�*��z*Ԉ,��P�I�}�$�k��@���p�%tP[��gZ,����ȼƕjld�]FU���s��9�~N݉�/�ȿ(�L(�S+IG>�p�跴�K9Zѩ������k�[(8C*ڄ�$^�5�y�
ht����P��v�}��MN"��N�TgUQ�%�B��@��;�J��uD���<.@�ύ��`�����>�"D���]�1�S���`��gS!�IU�X)�Q4�KSB�SQs.�/��$�b�������Jc[�	���J�o9.���˝��!��y�fU�{Ć�(T����VQlp�.������!�c�--_KA�5eHiYܥ;��]�ԎHoX�g���ş�V�V�{ף*��&U�^�w-9 C�=��Tt�K��y�M���n���'g�֯��,>fS<+�*��Y�{����D�5"��θ�����n�!d
���W{ ���]a�:�(=�Y{Y�}omѳs�$Y��{�:��+���j�*�����@�l}�_�9��c�,��D�\�~u�
��c�;n"%[�a'OM���c����\GE�[�-N��qO�ح�J
�P�,d,���j�ឥʹUU���['�l2tb��W���e�,qg�7|x��;�:����0F��s�����"�]~�����My�*�cүXPM�rC-:w������N�[5����9֞�j��2���	�|������_E� B����x�����
9x�7��{ʚ���˼�SP��r��������XRq�(O�[2F��$q�W���ŸǅX@�ԙ/4(�hr�Bjn���";}� �V�a�1֨��W�x�R0T�':�a�)%�	�>Z��k��OY���Ed#�΃=Ѯ	=����{J[�X5<��d���4��
*���i�,O%��w�ס��ns�pK]���FYTx����j�m'v�΋v�etPP��*�����88k=ZD�<TҊݏf�Nt���@�����=+����_e��p�t���r{X*&��@%��ޛ�[�7�%�Ww>������K�Kv�9{�'CMrȊ��n8*T"A6�]37|)8�Y2�{o_!�rL�˓�K|搷����5�;�C��/A;�}p���8�U�Y]zs��֣�rT@^�'	�}�5�����޾���#�n���L�yX7���M�پ^��E<$h��mׅO�)��P>�(��.ׁ�^�����J�Ը�ĖwQ*-]�~�Ԑd$K8 ��C�1�k�yʳ^g��٩}Zw*VC67$a�X.Z�1���� �0��gu�Fyt�]E��'ɪ%�L�UG���.B�+��R�0�+r*�K�����
������Uӂ����[<W�o��+���+����j��5�k��N)&���g�6�V���o�EO���[�2��G����)��}4Z���8[y��2[{�Ex��s�/z����̫V�7�*��Y�M}����8�U^ŞM��x-���}��G!fm��;* 5c�B�b��aS;O�<����?+��k��:BH@�Ą��$�`���$��	!Id$�	'�!$ I?�	!I��B����$��BH@��BH@�����$��$�	'$$�	%��$�$�	'�!$ I?�	!I�HIO�BH@�rB���$���$��b��L��D�mx �ſ � ����{ϻ ����&�|�@�4�V�B��L�- 4 (  hf�*(�H��`�! ���zC̶��ڛT�U�Y�ZԅA��mQ�nL�T4��&-��n��M�m+m�L
ֶ��4�ٵ�Um��Zm�R%5d�-�U��2	m���V�Y2Ͷ��"��-�cͦ%��k[w�J�v�mG� =݅��4��J�w:8�[��b���+]�� �0Ӣ�݀���Di��ݶBՁ� �Ov�f�j���Y[�0�e; Ν��tSS�.@]�N�έf��ػk�͛m�� ��hz��� \��ۭ�е2lsq���ӹ�4L��8�5҅uU�m6��Ͷ�mi� oB�X ���v�
U6�w�
 ���  R��{� �)Gk�t  �);�t ޮ��N���6�F���x ��u��ݰnݺVᵵ�;��:�]�En���m��TTV5k���jݪڡ˶]s����۹��Z�ٻ�T;�v
]b̩JX�l�  l���Z�sv��v�j�ݮˮ���mmvsWs�6�U�[]�����]wiѝ�w,�����wGvkmU-�7;wZݥ���d��r��,��  '\�Yݪ�jh���Z���9������r�]Yݝ6�u�f�][2m�]�w6�wmvƧl�m�wt�k[9��g6wF���̥�m�b36� �y��6���۸jn�n��ۚݎ����s�wk��j�]�Z�٪t˳K,�rC\���mgUu��cv뻎�lV�j�՛�� 69������k�\��nv�v����������ڭ�ۗsk�k�vN�f����`��h6�`�3��Y��ZV�j��� ��:@v���˸����(��:��Z��uL(.��v��O}@   &)D�4 0�i�bi� ���IT�� 40@�i��)��%SC  �L��  �~�T���h4� ��M�EBd	�)�2jj{T��z�P	�z1A&�A��A=#  y	� b1��8�H���0³�o�0�akM9�y�o8�j
	����� �u���Dx
���S��!�UJ���h�h������	�$���{��H�C���+!P�]��?��Վysۀ
�	{`M-,����(���8&�p�K$�Dt������b�w���K?i�>׷r��R��a�Z"��q�L��G����jd����N�����eR�K͹�)�{��B%�V5���̧�i��Jϱ#�5b��z]�Z�+⁫�v����+KT�V��ѭƮM�J�0<����J��N�޵
{-U�g ��)ުt\{x�Z5$Q�j�	L];���
�2���t�I�4��M;�����ɧ�1�ȍM�2�2:j�j��
�D+9j�8�T��(��K.*!�[�m];�
[��&,���dF�Q�/��2��Ռ�S(�4]	yY�(U�^-�^��3�O(�)���#u)Є��w�kSn�ҾSf!��&�Ch����F��F�n�U��=�ᡩj�B�f�iU�7Y����B���9���M�m!V���R#�
5�����o+F���1+�Rn��T�$�L��9mYt�݇�A�1,G�����w6��#�
5>хL;�G]���k%c�u�Qj"���"�f�4�����2�+u��q8z�\s�*�WJ�)e��!�����R��0����J������*���n��E�0��ae74fd��f-k��'�nS�l!�vO�k�l�a��J��2P�^MN��˷�S��\yz����-�sd�wDi��YY���凮7�&ִh�SS݅�6�Ԧ��@֐��ѧ��[�{YC[��dkIa��d�~���߆i�Z�n��1��Z�[�t�V�о׏�cx�	���P�iS���,ُ&HV���u�0���[ԝ�t5�ޏ�m]3�4�ڹX�̔���ҝ'��o!Z�j����%�y��!d2n�ַ�(E`����n�5h
�Q|:�򤻗4�6w�,ͭ���N�e�U��j�&���(+�PI����:���h�[�m�^��٠r��/+=�z4Rx%u�ZCd�ު٢�[���M;չ��:��e����Tl�\��e��F�����3N���Jͳ�!H���-��6�j�x�`k/j�Eaxt�p��%g��:��n�E�Q X΢¬ch>v��v3��f�!�n7l�j<�S5��͛{�m�ݗmT*��Ŕw�����m�"wk�*e^��D�n+�m][gK���h]+ڡ�ˆ�U��=���v7��7���ŧCq�s(�$u�7�%qۡW���R���7��:��q�컬T�n�}Y�j|V�Ir<���������6ᢦaD���-Ո�n�(�R��7(!$�E���#�r�l�k)�o�\�MR�j�X�R|�4��CT��+wJ��%@���a��z�mmZ��=�XɑVۢ�1N���S튞S�;r��w>jdy��]�dIF/j@r�#Ǌ*ܒ�m�3�#抷,S�1[Yu4^[�~�h
� e�]K���)|aK[��1ZM�aoJ`e��'Y�[̬u�F��oK\�v�֫CM�v�F�	��HP챽��a+�.��76�R̔A&�����vESBܴ�7)̥��]۶Em*�4RE�zNv�٬��xS����m)�t]Y! �s���Z;�h��4Z|��VZ�oZ[�&�v]��2�qz�Ua��-��bP��:Ɓ�5{Pᕚ����Yj�a-Q�l�kq�XVR�>8 gV��^Zo��u�j��������l6nk�XtQY��o)�1rm��:T�*��
��9�[�N�:��և J[��	�*I��A�R���j-;�/-���s]fT�.�)��ܕe�e�tՑn�l×�^�� v���	r�!`�$�X�,�YY6�b�/"�j�L�ѴOn�&˅%�H��tB3(�wf�RǧVU�.� ֢�̇6�1ǈ�2Z�(�"�3z�������&��њ��%O����]�pQ��������x�>ҭ<���w"̄3��d&�Ln�����{�e]���49Ыl֬�K�=y����4��W1��nm[�0��rS��PmA�K�yYn��[Z�u)p4��z��V	�1�.a�xiڼ�髛b�U9�W���Ҩ��f�E,��}�=FR*�J��-t�4����������	�d�Ȏ��*ę�x�Gj���S@|���M�Pp㽎��/L�T�9�ӡ�+oZ�Q���ME��(�S�å�/-a���j��֮��1��Y�.V(���	3Om�ݼn-�4q�XLA6,�p��.��-��-$���
�c/6��E��s���Jȿ��Р�-M�!,�w��� �a�tiĞbׂ�ئ�(V(�]2쯥l�-�Op��Ss�w��ܺI���ֵ��j��yrP�:R�z>�X�jڎ�;�&��֭�Ie^m�b/+�%�����5��ŽدT��Bh�ͽ�
tńKK0V�D�Q����Z��/^֩/��fa{�;�(�g(m�J���9��-�1Ҩf`��Y�y�bH���
4E��f
:�F���k3h�m���t^�R��;���ګ���wv�9)w$��f�Hj�76�;�\�RXw�f��opQ����Z[5�%me����T�u����SZ�O2+����ⴎڢ�(�fVdwR�����	���-U��%4�z�2�i�V-����
R��UU�(�6Y�M+�$�|���Ymޙwj�U�����bRԥ�Y��,R ^b{�m��J�C.��ð3}Ĳ��m:��랶�����.�d�3~Zۘ5J��6�e��1�[���i4�qe�s"�7Z�fDi`ƀ�S.K��ҶÛ�$Jܢ�����V��jee��YCl�kB�e�K����D��Ö��ԆZ+I�.H��F���ّ^�5��:�	��4-ު^���M��y�C�n�m�P�X=J�"P��捭��I�C`d/����K�1I�Ҡr--J�K��S�����`�fj�Zz�0�����Z�a]�On�\����Y1�`-�k���8��!tB�C)]�x�jHn��{r�ƪz*�٘���uΗ��J��
Ѝ���|����Y�Z�'{y�T����j����<��;ޣiō��3v���r噡�I1f���B��.�xP��7�^]
$wlm����-��YZn�#��t���F/��-|+���E:����tv�����,R��i������h�7��r�<��t ,�- b�N�Wy���6�1�G-Jij��̲��{����J�p���l�p�����dt�7�L���J�E�K�nR�f���anh�n����MA1E�\�GNպu&.���B`�w)]f�{s+,�z��+�U�X̠Ԙ":4��gf�[2���[�b7�u��އ�$�`Au�vT�H�W��$uL���u����p�\�W���k|U��݌�(�����PTW+K��.U��ݚon�b��y[P�"��_�SO9Y��л����66��Db*��ș�����Y���5�]�Ձ�Q�r�N"�9k4��+"M U�9��3���U��ț�/�]�ܔZ��"h����3vA��2r�=��0
Z�z)�h+l3�u�\--�ƞWf�%Vv��cI��U+�H&�AH�s�D�P������Ŕ�������n�ջw30Rۣ�)>�o�b��ȩS��{��Z�ܼ�V�F�b�h�pnm�y��N��jn;�����:�+�K6�ű\d�T��cl*3�GRU�kT�#��u�F,�[ i����V�=«��Z���Ȇ2vQ�`B-3FV�ߒ÷YF�hVde�t"/��y�S*��4Y1�j��][�X1e:��ԝ��L滦�7�W��	�y(^;��'�I0ś�O�9�K�ᰨ-�[{��H�֎u6
O	��V��2���ӬS
܂���
T�*)�f:y��񱂭-p4W��6�7�Ȱ�;��sK��(�Z�{w�f�P�G�
��֫i�7���{t[�z�qS1Y�RQ�[&ٹ��xҗ��)�h��]y��Ӈ
y�u�am��V�A�f�`��7H=���]n��ߖ���Z)�Ɲ.�,�ɨ���s	W�j�VZ��rw�],c�6���-� 8f'z�L��欳�F����䡪�ZM���fZ�J�VlD� 3#����0�Z@�ܣ�y÷.��4#�ٴ�b�,/��tz�eL˭�6�xցX�S-���h�PJ�tūc��{��q���KN.�L�.$!� p
9xJ���mLBD�d4�@ٖ�D#p�N�a��P��4�	�v�ذ��a�f�f��#/t��-��)���p�t[U��[Hh��f����B��]N���R�YH���k
V�BTp�M;�(�0c�3�,Z���CCܫxq5h�k��k��Yކ��[�:�4�����&n����W��pdܵ�vغĚui��A���S�f扭��/U�U�ٮ��%c̬8
J�x��|JݬXLZU0Fd�n`8.�n�%.�MS�*���z����,��m�Se�s납���NAj`�{tj�̛���3v�uq8���m�Gp��7Y���+zWU�Z��"v��V45_nd�+e`�7�s�l)a�&Xm�rX���5�8��fԄ��y`l��y�h:{�h��ʺ���f��!h�5ی&]3��XGw 5}�������q8�e��"�ރkŮ�
�g��-�����hM(&�Y	�=�������Mq��,@���0�b�&��SB��+��g��'+����)iK��Jۊ�c@����mv5W�^���P*P�����Nwq�*=��(PM9��2R
�N�M������%F�>k6Қ�!��8��%l\�k.fqAa�rZ�e��O(fR�&d�����O������>�=FRh]���cD*�X�!���Hs�c^�� ��P<KU��n��e)�5r��n�Vܭ��A�V�k塥Ov�i��V󆬖�j�U�1h��c㩤t��4b*�4��{G�f�Oj�x^_k�Ɋ-�{�\�iw�LQ䴊�і�&p�z�[;��U�-��n�W�q���W�w!�l��_9o���ee�pw�o�Z�9dQ��db�%zP�����B�.ojO��orfc�,�/��U���u��h�v�AtDNY��(k�W��X��/E>).Y9*b�_S���FtUb�Lg�g�b�f|�W�oZ)�Q[�@�\�z"�v��8��o2��ېs��3U'x��/F�JE��`Th��Ց��Ӈ^�W��86t�X��c#l%"٩�X�UJ�)�@���αdj_\�La�[b���P�s��G��� �5��@�|3��:��7�rbZ߭8�e���#}2\�1���r���NB�k�{���P�;W0n��6���3N��$Z2�[��QW{kS<���.X�n���Y��`��Z��}E��O%��R�僚 :<����̋�vÉa��3��5wۧ����`o /���wmBZ�����$F��Z�״ `�<��85�3pٓV˛�f���%_�9O'E_x�S�|�p:Lz��\�{i8K��ֽ/�
���ıI��i=s�}+@U����d���J静���*VA.�&)Q� ��ą��\�9�1+��.���r�Ӳ���0�kT;,a�vK�c/@�GL��� ��'��S���S�Ԫ�娮��u�:�"u'm%�%�a� !�[9d�j�"涉2��͗�0-BS<�uS߮�Υ,j�Oz,+�x�����%k�Z��en��@��`�]أ��M�y��8�er�T�Ǭ(]_�n��n��v�t��eh�ygFO��Э�iE(�S�2�Y���t���v��]EZ����k��tu �A
���u�-֍�s���Q�c,��$�K [��D�SG�բ��V�$9e���2��c�`�2�d9t����1e�������)�+3B�WqԾ8�cf�E�Wm����7��Jh`�`����]��R�3�);��Mi��T���s�����;+�l�>]����|�}z�-kT��`p�"�70
�kO�{ls�L���v�|�F�Ӧ�0��L]��كgZ��d:���=H���W[d�kZ�ڼ�����W��<�ZT��^��Y��b�]����u��L3봄ki�:T���T2�$�+m�wv���0kt��I�S���8,�*Nc�n�&�ֳ�,�V��H���1��X�R����"us���gf���1T2��ei��'Jn���<4�J�+z����0
W�d��,�I�]�,)�tc]�
�n��d��,�f��
����Ht�"4�!�WDk�Z)��
p\��ܬ�z���F�� me�� �eL���@�S�v�F�v��C7c�z�v��Pti���-.�Y�]�˭[������R֧t�^8���FɳJԍ.W.X�ɽ�^�WB4�+M�nZ*d4�-fV�X�"��M�!����ɲ��+�i���]ԥ��v����(Po�闊rJ��]�zf�)|.Ch�����c�JK9��Zr����̨3J]$ϭԔ2lq�8�ik��.�'�Ŧ���V�*bδ:]`�kh^��B��19���(ueF�{��{�nN���ǃ���=�m���n\�Fv��a���c.1G�#-V�qؙcmZٴ�i[B��m�M���,�,Ć�Q�5,����S�&UΠf�Թ�f鉌Xě��b�)��|Ɯ�ǋgk���UxW�P:/;�&0�����E©J�w]��S
ҭ�q�e�n��mL��ŇV�+2�+�g9=s�ދ`E����ɩ��(|�[����:�"��g�_Qs�J7��f1pdS�?�ƪ��_\�q0��b�����+��K�pl�f�,D�+F��ŅK��u9�w�m@r4���0�"�[W�M��\�2��T�v�Em>��<sU=��e�۽G$���Fњ��,���C8�׺�^+�frx��Y�����r#Y]�6	`A�@��5�,�7d����X��QJ�����k�Z�ob؁���dA���mvSqw�+�a������q��LKu�\�5b<1��v����WGK�������;�¸γ%k&7��o�Jb�@�/{�p��[g8iK'd,>�"[C�T}.یJY�����G��iׇ�T@k�Ӽ8�p����� \�o/v�S\��)��Ҩt�	�����|�%]f�
�<�Na�n'�;*W:&�;�v����#'�F���"�4���!lPTD[�/�"�JN^IY�NʱWEF$��(��wuH�m��f�U�i��Yyy0GXl�(bۡ]��"�j%�Z��tD����w*a�1b�3�R�JϷY�V�W[W*
�6��C������JO�v�i luz���J��;�.��c�x��2��,���t��e��.��yw�Â�M[U-T��}՗@���)}���En���P#"�6z?��뉝̭��$hY��m^Y�Ԑ�2Rm���}��F����^��w���^}�{��3�����~[����O�'��2R89s�\�r��a=��T���D�۬�ӕ�|�"Ѱ�"��:�:y��	i౼���`���v�=)���Ǻ�KE8��}qJř`w]*�X��m%J4��-��5���$e3/U*K\ۑ+X��8.�پڽ�/D�EW^=��Bf��ƶ�.�E��dS1�6�� ��mU�CV.�}��������܊���snˉ�p������gm������M�Xno>����k���{���9��܋}�-4�X�5C�R�xۑYu�yS����VRt���*�j�.pE���&�D��6�E\���!{�,��wd�m�(��s7��N3��wiߖ�uΞܵ��Z�I.jT;������c�ӮA,��� ��*����]d��byiX�,-��o�.��]���;�f1���ό�n�6m)b�G��2���ݭ���i�c�ܚ���Ou�㳭�x�$]��;���hfm�@E�	y*�F����,p��F�V�����3��?>]uwz]��E�4�X"��=;�y�̈��M=D�����I�7rnc]s&�_j�NJ���yİs���xukJG���>W��w�\���UwG|�H��f�`�
^�R@�M�.V����=��� ��vg%�_d��ŗ�pS�/`Il(���)k���N�9^a� �	�y�5MV'Y!X/p�ҏ��+�9m-�;��B�ۿ��h4�XO|�"�lL��eo	8��2�*�W�Z3p*K1�ǲt,�&+-�k9��LZŤ��R�Y/^�vq��7K���$���v+J�������=��ni�N�l�`"@��L�j��n���c{8\�C��V+�pkU+Z0 ��`,4S��m���[¦G���e���]|CDi=�T�mp��w�c����P<��E�J��1�oO�̧��O-�×vTٟGO�]³
��͵\��z�j��*.93���6�IEf����B-�٢�U�#15�E`�d�%sLg\�I5��7M�Od׵���eg^mH��3�jg�J�5FD��6���ms���i�����5r�8�ȓ�΄X,[�*�i�L�Wƭ�K��V�U���vPv8;B��+�C:6h+��gU��]M3x[7s3^]
P��4��`��A��v�Wu��v����6�O,N�h�a�W�hch��h� 7�"���5Q��`Ey���ռ�I�(]�;�!*E�u�EE�]��ǏsSM�p�˵NGV���(����;��4k�l�9�Y)�:*�s���|LBH.�@���j�Y���n��]��tN�Z}}n�EX�e41@Sݐf�f.� ��5�u�/*��2�����Mo&�T(�ۡcyʾ�6�/�E�]�+�/6��H��֖,�ݗJ�w��λ��]U�D�Y��Q�v�D]ɐ��'EC����^c��zn]�ur�+�KO"J\nF��`�X��;���q���n'm9��{w����y7m�;\SN�Λa��PO:�άKs�Ekf`t9䭱�r���6r:X�7��J�T��.�7�b<�>jU�a.V�CSE��j�bkU_%��KbjE�G�� �k�S�;��o��\,\�I��lr�u����G�% R��ʓ�!��SnX�M������^:�;�	��y+K��'8�Ԥ�I$�I$��L�ʕ�%ٍ`Jħz�R��ЭB*6¾�Bj�u�7nBt��KpZt*N-䷹^E��q�wC,�ղ7�5�a��t��l���<�Yaĸ���5[IoW�O��Ó4�jwQ�c|�##�;���AB�u�k�,��J�z��H)1�"���y^9�Xp�|C{�d�}�k(�1Čr�E�	�S3ۻ��CMfS��X��ETA6d�R���DEA3�"�\�v��eD�2/�pٕ,ck��o�S��� f}x�vֵ�����vr�(2�*�qiP��;ױ��j^��Z�[��a&.]i5`eL��j7�\�2��nƨF���'htI���A�f
V�n.��S���IS��ڄ�*ZѪ���������k"�54�mbqJ�γVW�K�-S�-Z�G*�8��ۡ,�,��㌹r�;1�sf����{���,��o���*r�����R+-�9M�u5Vq�C���_v]D~Lf�HPh*�G��݇c$����_P��"�VuD�G6��1��K�y���w�m�ʐ�)Y��������L�޹�Ρi��he5�mpmKi�Z�:��IfޛAUᭇ 
�]�����Y�ٝ��;��ܤ::s���5"�t�n)�V����N�YY��T��$��:�����&�{ي)[��I��:�޹����̨�2T�L ˑ�%geԁKUE�d�����^�x)A$j�e�Pg�^ñ��Q�)��:��f���Uס���K�.s|��{.ɫ���l�\vU��a���oi[&5t|~����r\8+�F���PY:<+9UNǆ�,K̶�[� D}zsj��
�U����wiuM7
��5k&.tr�F��щ�k9[&wEޤY�I�c�(<m�J-�縬ݷ���� N����h,�b����&�l��n�c��moe����:9�׎�h��	�s�]���Rkp�MS�i��3X7�z�5�s���)zZ��Oް��E�F�R�)fRV�:mB�uy	��8|�^�Ŵ8��n�r�<j�m�簶�3�u[�~ �]� ��iq ��Sp}���PsN)VF�À����l���Yc�q,m��$[���`ʼ%��� ��0¤luY9
8L��
�X��eb<X*ZKe�Cz�dg_V6��LWaw�u6�X�l%9ou#�Ax�E�u�k	R �Cw����hmZ���H��W`8���dj�yq�ɡed㋝��iy��!���f����.٨�{�Tр���d�\RP����M(�e�i�;9o�HF��ב��XL7r���7[��]om��k������M���m�iT���с�t\AЫA����B�����[��c���UȬ�&STdz1��J���s�z��-����1n�S�������غ�nS�p��$6[J�ʝ�.INt*�c�Y��s�A����7��9K{�*0�oK�"�_у���;�J��b���&u��oRCv�F�ׇI�N�b$$���joV�qpYۯ0Sz�Y}���u=�$�Z�T�Kl�\�v��+5k^*U�m=�9����ud�S{/��3[7��;y�쟂�,w���������;�⑊?���7�nA��j���PP��E�un������:���fS�#��y�U���K�=��O�f	$㢬K�p�n��Zw�d�"�+\T4O-Æ�.�Z;�WXz�����2:y7[ɨ^mfWV&r�V�����R�ȭ֘��UQVG�1p���+C�y̦\�oi�N
 �E�2�Mx]ܣm��X�����ͺ�Q뺝�]�t����R��t����We�j[��ʻk��U�:�=`NQ�l������Ûrdw���Tt���/�vv�pVT�m_r�z�qJ��败[��Q��kl f����`���9j�3e�2���=V��q���u�Z�&�Ԩ�c=���g0�y�$g�k"�k�u�0NS��u�=p�j�h,D���f�GPnݙ��C8�R�hq-I���G����u�4�P���s)�:�7>o!qꡌY{�����n�R(�^�z7����b�j����mko ��2#\�ʙ,obf�УVG�sy#yj�s��y\���i;ʆ���R�������P_+ ��jZ��Yw���|�upV���=,��a|��`c�l��}���r����;;�m�? ��<W ���v�s]���e �k&Jڵ��A����Kp���G��v,�h�`���u��v�V���|�R�]��S�pv�������xRhԜ�˳����HҼ�Υ޺E�x�v"��q�c�M�~L,�X�&�6�
¾�N�I"�DN[b�w}B��\K�Ƕ�>�:e�81D�`��74S(n/�uݸ���M�$sVaF>����� ���+8�P;ܰc��ky�i5�3݋��T��˺�X��Q��;ʥu]f����qn��u�e/5��0u��"a�J#c,(�eZ�)�W#/�I�m�۳��h��lK��d�Je���]��J�w:�V:n<,ɵ�8�V�ٶ1S3RC>ޛ�j[�[J�Ko�b9o�^����|��F1٩���E�IN���-l4�6�VS٪'�gGB�0q7���"�3�@�,��bؘ6��@j3�[Md���z��z���従q�w�7��b[#dN��(u豽�jq	Mw$��fU�p��Y�eS�4k��Ф���.�=�X���E��y�]d�kv��8����;RDm�T�g(�a����36�a�{3 ��uwsP�Rż��:��-8{����/
��D�#[��ۂ�!��r����z�Z!�Rq�y�6�9(�*۫�m����CKD���v7�\�
`��re��*0r�jł५d�1��]�� h����4h�i[�qa�>W�[t�����+n�r57P��6l⡢��}����M\�=
�vT��{q�� �5��Zt)M�٣Q^O��Tw�4�*�z9������t'��ɓ�V�ќ2���!-u�1���o-D��Z�w^��j�!nR�g1K#��x��y��r��qZ�l0��kr��S��wR�eNc�\�DV���X��Ma�a�:�B㥜��6X˜�֫�Z0�zc��їݙ\p��F��-�#KU](L��.jE-WP�2evJ�a9wQ���vt��j��4�n�1M�0s8�]�.�)�O:�m,��I�-+�/U�'f�h��S4�iԕC�����a��`u1$���*��W�(����\��֋31�P�F��������J�u��b�ݽ;�e�h��qm�B��S�9m�	��]^,��)+HT�UՃٷ7x��.����ӊġ*	Y}�֢p��G�����*���q���k�W����v�F�G����+�����+5��r�xwY1�[�i�08B+������6�J�d.^%��.���'�ҁB��yX��(�"˦L��cde�o�wL±5$L:��7�Z�A��ؤ���������Ư�M���.����R�>[R�T�TXۂ�QɡVνF��b�:pi��c"jx^�M`�!�cp�Uie������)�bǴ��^e��c+�/���EZ�#�����2�����幵��C ��4��s���4�w3��b��9}b���(�s��0�Uj���\�V�yRn�얒�����)�!_b���4ԏ@��Z%�{�N�I�tK;Q�𦬮Sz�7aR�<]��edVq^w��M��Fr�K=2m]S�6{l�H�5��N��f�Z�,�{�uqX����]&�f���ӂ��)�T͊���Y�����d���u�\�`g,�ؐ��շ�it�6M�����I݉�˞�Q�	��&���G3�39N���ةk�{CU��\L�ѽ-�抸R�Ȑ�cpҝ��n�ͭjhP'tӷt�ԕz��31%���Y��e��|� ���s��rI��I�h��u:��륃9�e�2�@�2���a��U_Z1fP;�
�
=>�M<�����4AՑ��m��b@9�Pǯ%���M����uG��X9.c��e['@��λAWo@��+d��� 9p`y[��<�:����:�ǹ����ܧs.��)�D��r�s�Ǫ�7t����XBF�RF�I�(mC�E	gyf�W5��ɵk��{�8a�*�\�2�Z�l���b
����M4x�uk�tQ��ɻԩ���s��ro{�Ʃ*���e�D�X��
T�k\���Pw��+O���Z����L���^;���mI68��n�I��Y�%|�`O�+����`WV��6'��l�G�,��W���i�@�9aoj�%]�P��N㙗rgte���2�늦7��>V��KڗK��f�.-�&D��V�V�5�̛�n�n^��V	ۚ����NNct����+u�y1�����_gH����{t���@h����d�kkZ��B�g;R��Ց��G5SY[ty'a�����讓���ce��Tဨ���Y��+2��l�Yg�D��Bt�JZ�y]5������S5P]u�uc���������K��w���ʐ��F�F�<F�^u�¹��7�4�نVYu���ȣ�m�\�9�kL����MiYd�w3�B0���e�If:�K36�~ ���CH�S�V�������ΠS{J�eEi	��	��ek�F^Kw�8 D �+	z���-�����op�&ܭ�ԱA<��q���1�̝�ռ˜4�F��Em���	ݨd�O�)��T���p���[u�F���ΰyp��(6�n�M������dٶ5D	�R���O��Ћe<޼�U��ꨗ
Xt�y�9�/��	��tTA " b#���|iA�IB"b^c��h�;|3�i�ܔ)��=V�ӵ��ri�^��vT+;�w��A����Qp�0ܙ�V}���ib���H]�/�.g�ﮜj�7���L��\�<j!W�����X�#N���WW�I���Z��֞ġ�pF�]�
0l}�Зj\p�����q���u�䎤�k/.�ZՔ(�8���$�DC���2��6��F�AX6�圛�����"�J Ĳ�ݐT,[�{�}��^]or����B\�^w"�!jy1v����\�����H�C��,^
����Qt�l�"Kl�R;��"��u�Z�kV��N�-Q|�b}��ރ����j��YC;�k��/�Τ��V�(��|&Q��af@����ڣ;σ�BT�#��h�Ǡ�?�����"�J�dќ�����n�qKK2�̧�df\
�5'9��	!�%�v�6ftY.��o�uc���6F81\����<��TUH��"����EU�@�A:�pDVe(�ʕX�"&5�E��Eƈ����;�QAT�j����j� ��aKX���H(t��.5&%J����֢F6�DH֖�-��1TB�1gM�]!SV���.dę�����(Ĉ��(�"T��F%j�X�+Fu�W(�n�m�!`Ԫ�h��TQEi��"*�Q��E��e���4�EV"��eCF"*�EB�UJ�Q`�e�G�{�Ϝ�ֽ׾�����H��
Qx����p��J�����^H�=~�C�	'�lpν��I���}&3~�5R�k���a��&Va��jjt9u�ߪ��!���Ia�[��y�q,a8��r�*5 ��"qr�GT���y�s�G8v��ʎ�t.�^p��3��صչG�)�z������(�hjЌ*L��V�[�$Osս� �~��>I7x3r�V�|u�a�J0g�8"�P��j����a��\��������e��)��>\`����������I�^r�&5��)ʽ������E̻���Sg�;T���R-36|dH7M���ܞ_|:Mno�����1�wu���o��ӽ��F�m�{�_����MK	J�":+.�C6����+6�Kjٺ�i1;�aP��B7��v�LL;r�]�:��!)�$�K�-}�`c�K�\ȷ=ue�k�u�x6�ڵo8��p]�*�T�ѹt:��Rܩ������k�#� ��.�C��s�,h�`'N���N�MvW��[EA�P��va��}�����.Q̊ڝ`e]�j��T;P��Tb�E=4E2&�)ͅ��������u���������Ū�ؽ}W���Fd<c{�R&���Gv����bI�܃�y�"�j��{���	hNf�����iX��S�7�	�;V�ξf��<I{�[��*��R���/S�R�vΈ�x��a�젡�r�T���lZC:�Z�嫾bT��Zq��:[��z���Z�l�}�2�"5ک�ҩ!0r�E�e��/B(A0�]���<��%J���B��0bai����D�R�4�Sw�/^wK�EHa��x���A[�v�]�M��33�ԡ�����
f@r-=�E�1d@VRe�:��F�l�5���G�DĂ��J��ogv���y��#�9�l��Q��_A\�*��Zbl��S(8�5qbv�R���' T�A:+DN��<�ߤ o�s��:�߄u��ګh�H�q���J�z�{�w��pJ��f��n�� :ě�r��s�;�j��͓^�#��ѾG�}�*x����'�,�l�;�~��.�U8*��������{Ҵ����(y��S�2��+�O�n��k�e	Q!F�ĺ��I:���&�ۧ�6�ح���xK}nN�|�S7�$�3w\�NG�����L��V�JG�����IͯU&������=�v*��o����-j��uz,d󊬾�q�߅e�X,Z�ǯ�h��Tl9]c��b��SS��%Y\s��%��>�;qX���j�pc�+"z�#!n~��l3�[�m{���z痴NTV��ajl�!}�f^�i1��b=�s	&���ʩQ<���1��4����+/�^�k������s�5�
���%�7g��i��U�S\&n��*�i�Ri�ā�r3�dJ��<��� �6����[Kzaq%ߨ:���ҵ���vA�&�u�L��l��\�[8���e!�*�f��1��-$	`�C�L��'�Y���
��6��y��).��d���'��V���*�n�j.	�1=��{oMfh�dl�@��fjl�L�H�!�8Ӟ��u�=��uu�L4_d[������ �G^��Gif��;���'d6
Ws.��8��Tω]P<ckuK˽��q�Si?Q�?Z�R���+t5��`
'���8m�e'*'x�
�YǍ�-:�����\S�9�a���۵�	�Y�7�@�50@l$��6q��U��r�u��8�Y�B7Yq{|�/3�C[u�������T.�\g
tf�d��4��\iW��ѐ��6#=pj�h�+�-�Eu\V�q���oڞ��	'�Hr���˫ݧ��cަy�/Cdfw���P��FF�rr���8�O5��4�M��XA�R*,��!bUK�,�]5���0��Z���wۜ�.	�		%�.w�F@Edi�\�w��s�k;3�F�>L����r�	���Y�!��;�4��QAe>�ڡWS�.8(����$gec�UsY��޺x��c&�VEo�T�g��ⓥc�<�s�o��R�P�ѹ'}D ��F��S������u�\w���It�
�����+�=�i�0e���j�3|�!�����6��X||��`�-EIN�.+\�{x�1@;I5��]� ��K�ΝFD1s�uye�|�e�5���H�������iP���*Ҏ�T����)��-V�+q@�a��hV�*���'�|T]|��g���ZX2ݭ<M�ɻ�*��2*;.^���]1ѐ�݁a�b��J}�Zx{^YUǆ�Ђ%,67A(�1L�M�c_W`�荵uF�C��$�Q�S{��06/bQ9�!�-�~F�U�s���X�q���ۂ�F�i8�q&k�3�f���My�7�'��������gK��7L��FM5kC�.���ē+"A��l,��1�{�I���hܯ3�bc��Dn1!���7TL�\Bc&ÿj�7<��zc��I�͊]�X�7�H^�t�{��ѩ��1t���P���4�F�,���7��=L7��(���'g�8V��s^���6�zq���Wjv����8��+����*$�=c��(WL@���q&z����pm����o���^5<�VE���Z]����͒��5�+�P��}�r��mu��c��̤�C�]*���Iw�ω]J�W,A����]�í['%wp�Y����\e�ΞR.WF�W�m�p�);8}�JNŽ��?}�WA��ĩ�uy�Б�{�i_]��mZ�
�U~&v�FmĚ���R�(Ovd�X�!mp�D�Зv���ül���֓�.,t��:�57�� �\��.���6�I�ZC���y�j����$�,�\1�i;��/Gl꼻��̇`��L2��;b�>˲���hR1ӛPE(��;J����4��	��x��ᑥs	&�&:�����nV1-��̯m��p���,�y6�{72h��el���a�X���7ފP����)�
ո��<�n�u>�!&�J��X
ofꛛF���}�gsn�gh�	q�k����Z��d�_=VE��\���ս��z�}�_�|	ؖ&w���N�X�X�X[Jr_����+�%�eK`� ��L�<�R��n�<�i�Qb���U�.��:�Ԁ�̇K�(�?)�s�ۖ�o_�ꏏ��\'�Yc�E�����ad�R�Q&84���b���qC�%�y�N�c�q<ikO='���cһ t9J���9�_@��H��8�z�0G�����D�M���i�aq9�=�:�
�o|�1��Ta��V`?{C�B��]u�"��S y}�(PA���
�;��oی��ž�Y=z�:i)�~�w6�BJz�ۭ�F��-Y�LAm�Gh9�֜��S+!O[Cwo&�o�z��,�Gc\r)*�s�qk���OoWV1�'o.�P����2��E�[�g{	������]r8�^`�b�q	�q�Y��CZ1f��#=f�%�|4'!i���C�^�!>E��|�o}"d
[�����SZ@Ư��I�֓���%�)]bp��f;����x=ίx��oi
}��z.^n:���6&EtX{�3��K]�s6z���<$2jJt�d����A��X�Ǔ�N�lr	�[x�R�����F�0Ǝ�VZ��K��� 4��b{C��]a-H�/���&�5l��7�t}������3���lX�J��Ɋn��f	}��̸�%�Kdq����׮���n���x�$"�J��eK\�L����s,-	z��mm9f�H������(c�Sa�[��
u�ᄆf�5��V�+�p	�����nȣd�9e;p��( :������,9M��+#:1WoQ�$�1���ܫ�WU4Sb��cA�n��?�J�|��S�/����wZ�;|�(Tّ";ᢹ<H�\���Hc2���gN�/�&i��K�:�*u`�4&Neڳ**L_c/��˪�%F�r��Ӕ)��تf.����#�u#F���9����;}y���o*̺cT.��ݫ�a�InncY=Y�z��:a�C/Z��l)]]���L�{��tp7���=�n���J&k4X4��u�}ݹ�\��҈�r*J���{�HU�G����[��k0����Jk�̶w�g�&5��;��؝���\�؝2�x�I��+�qݡ.�Q<f��y�������	��wK��2{p*��yG�S�}P���}�#pH��]E��o��wG���T�/�x��k/�
�H��(T�f�X2��Tf昁��|*cQ�>d�w�v��e��3M+���S��-#�Etp���r\H��C=W�α�u[���/V�o��1�K=�Ε�[��b��Ԩrs� ��:�wAi�_��K�j�u�˩�m\�Jc�f)�Eƻ0�
��n�1�P��fڈ�B��c�#u�-Tt�&�[�B��[����oi�j�\˼�Oq+�%ik�Ŏ�L��38�vT	�"���Vz��Y�J1<����,�ʶ� /њ�lv��)b��m�>XuT��C�z'�.�־�i^|"�	�p��e�6G��\:�W{A���#!�o��}���hNަZ���G�[V5j*�#�u�+r����V�b�.�]���%��Z3 ���I����Vd�yA��ΆK'9G8gl�f���y]F��v�_��'��~� ����X";J��TQb"�9�UG�(����LTX#�b��+"��i1�����kaX���0Q"��E��((��0h�cU0�6�K�M�M(����(�����+D��J��"�V0�)Z"ZPYR�,��"d��
�̈�9r"�7W-�[��m��b��,�J�L���d�j6�ˤ0X�mT5lR",G�������n@����UF5(�km-��q1QEASW���emm�c+4!�"�KE�iZV�aY��+�����������G�?.���.��e�n��K2��3 K��w2޽�����S;����T�;�^��X�����@�.�u<�c��MEs�,u� �e�l�����վ�P>[���&��������'�(˄D�r#�qEtw�F��+��죜h��{Fmn�;�4��Nl,fr��ޢ4�g<h����{��R�͋��������%�<'y؝���
��-��a*|7y�^��ތ��ڸ���뮘Y�'��|��0�BL�ry�;��x$���ܺ%�R���~�V�<X�OB�����-��NK��1��C�>�����})�Ѱ�4	-��{���G�����B*$!��{1��`��+�l�rc�n�uM����Q�8Þ��p�Fw^V����V=�'V4Z��U�+�������5����&���-Pr͔1}��p��;�b�`=�j)0�!%��E�����G���xWu����=2�ޮO�����|�0�<��������mvë�܌�|V��؀.�E]%aSf�od�8�30�F�ȾNw
�Qw�-9P�׋�{���;^pu���NO^�R�íU�Fs�ǅ����-:xk��3�VQ�Y,󶟜PΦ���~��&�|J�Qԩ��b�؏2���_l�<�V�	fv<���X��7�6�f�x�|s�{�st/q�v�-�,������mvgN��G�HRF?�"e��N����dQOF;Ք��(�X�����\���Zc���zD�Ō���.&L�_wa�r�z�����;����l�o��2B5��)lYYrl��N�D��ubU �z]�M���$�Ԛ�Sm�S���m�t{�k>�33�����Ԯ��W�~�l�{)V+j���܏2�h8��8��2%���Ȑ%d���5�=�%"w3K/��4�z%$��uK�C����x�&a��n{�{��߰+�|1z���e�ú��ʗ1��H쐲93�u	��QwLLK�g�r����R��#�
#9�K�ȣ�h.L�;,����z"�i��sP��(:������hz]�tw����ӌ�����[Jb+ɖ���r��x ���.a��~��m@W ��::��_�Y���	n��tA̽�����>jr�1{o�V��RD�-�%�^NWN�yq�,��9��˯�9�Z~FMel�J�Ѭ��bQv��g�XDƟP���)Ҧ�5�%sO�q ��~g�5<u�U��Vx);�����/fT�u��]�qʹ�ƈ4L��_C�p�jL���rV��N��*���6`�Gj꼕�o,��w�w�'�l�#K�w��	�:ó]�r�e�%��R�p����1rv�.�P|�]����Y�u6��\��@�M��cj/.�ED*�/�E���G�Vc�ו̒=�ny��A�3�h���Q�%�2��
ܚu�=�##BO�Ajz5�I��ͭ:�{m�R�\���[Z@�j���̬�|w���"��b�%��!����ISC)ٔo/!�'���*�.��X�B�l#�n���(�*���0�]�U��Bx�_���E~������;�Te��\N+6����77ệ���e``d��>��NJ���آZ��U����s"�<23�:�9-$4֝~���"T�q� �t�1�:����V�wW�k��.��w@�� ��1P9躽����46Qqz^Y��{��iԉ���	����7s��JW�fͬ��֖�*n�*5{��ޒ��c�m��ˢ�K��ג�V�1ft��ӈ6���n��
w�r�N�X���Ժ�V���,�WA�����6HB���&d)�防�;ګ�TR�����Z���țbΞm!���Y�s@�Yz�`����~����4?�ƭ3��o�V_x��HEh��R�&�S�+*�c�5�M�Ŭ��T�����<��oO��ܫ
M�q,L\�ke*�6'�̘��.L��dǝ��An��2s�/��\r[�#�I��uFe��	��dO\=��E+�Q|.W6�qt�ur�K��,��N9�*J:w��v�D��Y�e�-y�����Zd���b5;�I;1�$_�i�VvY<Ma���*z�U���=~��Z�OA5jF`���[��%l�O5Kf��g`x���7=�0�I�wmөg:U�+h��H@`�e�\�O����/�]�ۍ.��E)�[ܝ�g"�5�ͧ�]=O �&��+�|<��|����:�ڷ�����ױW��1ೆ�Fj��r��&��ΗIb�f��l�,�gs6�K&i�Fn�Z�b���(�rخ�m�8�c��K�7WrBm�V���C�W�3�9-@���$6/2�� ��@���]���a��RK���7�ir��(�V�.��]u�Y�����k�[�^}J���d���ͣf��Jh������w�q[c#���o7�T'<�_��Cm���~
ϫ�k���K�����X	mw]��s�	�7-�VEi�x�y)f�?vW���س���/34��N���1�yq͑A����`���Kw ����(F�l��%XQ44���Y;�k�X<4�|RM��X��=�u�f��[�� �m����
��A�F�"��;��i�θ�0����D���e���N���w����Kލ���Xg0[�z�����,�Fj�x�D*���ԩ����Y��CA��ۢ�w��� �J̍�)�ќ!�O����֐���Y����%l�����s���^1mM.&$�G3�C���eCc����M:���T� ����wJ��S��y��%��򓨩D��Cb^&�"�����3��P�:��MU�;R�	/��:�-���i�~��Vy�ϣ��S�o�#�ݷ�l(�����v_�]�J��qiٍ�{$�I�ͫR�^챹J5=qctJ'1�ӛ~�u�g>G4{|1e~^۪�z�	�ڲ�F�8��̦p�{q���1�;�q�fu��Ty��l7�.���%����G�፫˹W39]�[{^4T���2^![��m�N�؎������Dumm�o8��AE�0�����ϰ���N�Yݍ�ѻ�����%��(fX{]���Y}�XZ�sT�m�Iū���,�O�g �x�h�àW�:��e�8��*;��f�p�"��OC��I���wX��D�f�A�i�l��GWs>M���:��̂�\J1��DK�C��7uw�� &2n�[�5�dװ\�q���!��,=� Y��<ZU�n+���!lE(	���= ��ۛ8�-����b�^Ĉꓸ��;,�N���`f,��M�@�{�ޘ^�Ӆ�5� *A�X��(���S둒�OF:�`CZ]��sq�/������YwApU�5�8������O��ݜ{����Ҩ$9�w>������,C��P�q�yQ]d��=n����g�vk2�WQ�}!�İ��owMӌ��<�!`G�ǳ)R�V���ܣ9�QF����yi������
��!N<%�ډ�0m�B�Z2�sM,�T0�V�5NnJ�k{EJ��l5ı�P{�{��� Eb�q����x�f	��B[zn��+��{��e��'�j�\1���Q�ZDs�u�i����jX��l��,��L嫔�_���b�����TBj�E���M�w���B�r/r��z��t�t�� �:����n��ʷ���]�5RG��A;P�,��=7x�)`zB���.k��77�z���W�0IK���s��������p���?�+}��j(_R�5�Ȣ���G�Ek^-��S\o �%Cw��(���y�GF9��|򳫮\���7A\�ض��z���"�V�{Z�/��b�hi��;���&�r�#�2>Rʇ;�͔��U�eh&�5v&;x��<�dQ�"���"�5�z�+Q��՚z�Ah��jKs�8�m�ͩ��T!�r_W��]����A�T� R���4V����Y��h�U�U�{ҹ:�(
[[���MxZ:��QZ��Ů��㝑��XH]�p��8�ʕ�E�1����=F��A8��J�!+b��RE�Ji--MT�i8�^od���T�*�nƅ:Sκ��j�rS��_c����5N����A<�k�4�m��D�\�u��B�YIȡkr����̘�0���ǅcn�ghF؁�ݣ���c_vl�(�.�!f�A[�1�bf�9P��S��l2���P�:�̙�i��G��&6o��H�������%׻up9D�]/bоZ��m]!��&Yj>lL�R{��&��X	ܧ�p��BO�`H�h�̻���5�
�+����$��V&��;�7����5�1ޤL���i�R�^�:p3+�B���� V�`�v����4�Y���t�&����K��eH�W�q@��+�C�wx\�Ry}$�ːkDEƥ]%`��h���Ƴ�AAtY}�A�@�
��(��=�ݎ'�%�^�2�3x[�nRL\�&���5�����m��e]-���횼w�1{��;��-�O%�f�Ab"��EK���n��S��F��0�˦cS���e-I]�*�eyM�gc�P���9��M*���q�����s���05�um����t���B˒�}כ/�4�W���Ad8qQ�XvP�k\�e��jY�uՑ��8���Z�8����'fAv�Tsz���� ��.�q�xm��)�Ҟ�H�X�*!��Ǫ~{�C�XB�b������̕[������+��-(�P��p�--u���mh���FVѡKlMZer�\2].eʱ�m�U��EY�R僪�����[D5n&����.V�faL�a�����̸e��0����TեM&3I(����Z-*9"�նĬ)m�-+[QE�'Ne*VTkD���V¢��T�1�(��]%n�[u��CN�i���`i�bE13)F���ЬEH�P�Y����M�YQ��i�qUdb
Xbef�k#R�J�H��f��j�ԫ��
#�I��:j�*�PTՕ��T�&3-���V�՚�`Ub���$��LT1�cR���9���z\Ǭ�~�o�5���h�WgF*H�[\9b��
gZ��u;]���<��=��9���1�i_-O9W���q7)������
�t����]����Uw�����g�-U\�(ʘ&�^���z^HQq�z�$\Kˈ�������h�W�=��5��;p���'$)�R2H�O���J�L���/{3�Ռ�Ψ�g�t@��'���W*�l�@ovjx>��v���%Q�gq�vAk��ɹ�'7����m��,�:+'��]y�I���o�U�:r'u��^����@;8i�]5���M����V�7��^8�K����<ך	G����;�|;Lu^]�C����Ba���{���PIr�^��SV��m�}Fv��V�eٹ�m9X�m�'ʐ��e�oZ5��oIUy2a��;xp�A�R����6�v^�ybt��S��w.e-մ�kN��]ft�R�_�舥��I�s��W��Ws�4�yC��Hdkyr[�Rs���Wȼ��xg�K�	&���3��h�@��N'�$�J|Jxy��;��sw�6��m��?*�TD��MA�vx,�r(��m��,`!=/1!H�"�bJo�ýG@��zVu�]���.��w.d$T�C}%]W����P�Oz��j�^:���]*%@R!p�x���F�1�0���Bg��=q��5V�T$�B�$���ǲF��;���f�w on�*~�,��׹w��������Tn#��[�5����*W�wl��2��)�@V��{�����mNo��>P]nv��ݺ9�������V�*rm�]9�����r��P"B������=u&�������;:�N��$��{�7x i��I"sDgA�N�:Ț6����J@���mn�z��<�ќ������}����4
���sf�ph��vv-u���Y��H��^�ܽЋBsw=�Uj/�3��e��X��7�j��m��9���h�]�z��yc-)S�.y_�+�|ƄޔQ�OB]YQy���v���<ɉu�1S�-��HƳf/omk�e���#���x^���ar!��gϖ�bR���:�E����Y`���5�������%���e��}oӸs��R�(�	\��|l7Z�C������	��WH�wm����"8�c��ź�ч�V419uE�ۍ�{--�)��I����lٚp\��?KB�P�L��ծ�;��si��$��_D{�e"Z}��E`�����hژ�s��N�I�̲g=k�����B6�p"-�_�;�Q�Ta+�S7�3y�����yPYJ�[�5�W�������s}���(����/,������0�k�gtkE-���QN2B�H�G'vu��`˩���@��2��FK�uJ�lj�6�o�ZaZS���@���X#�PEd-7����}-�앇x�4N����gVh�E���%3��2�'�R���.�D0�O5�rylp�m�Bx��V������\:	�;[AzY�o�D����H�<�u{N��y$����*ca�sh�:�@'���ņ��+E.-fE�U�eŝ6�jo��o� p��n�o!w/$5���(L��P�[Kf��򾯾�Z<�lu���z֍�j5�=<�ēt�f����|I$2�������g��P���7���c2��O0+��>�%Om>>^龿�5�a�ǻ���G�g.FL��t����.�=;'^=�m���|����*��>O��em@�}���5i���(�D�9|��-��}v'y��|�M�ŧ��;)dSk���p�R�)�y�l�*>�\x��9N>1ೆ�f�D��k�6ߢo���0ǞtU?]�Pw4@X2��zܞ�a�;,�����w.���*�=C����ԭ����vu���r���bo5��h-|����p��sw�Ʊz����)�'�r��`�)��]ov�c�e��_>��ְyI�(&f;��r4�������� QNL��?I�]���uTXŏxF@�M[LǓo�7���W'�ӾwD�z�Q���⠫C�4�p^�����۪^f���j��Ӝ�	�|��[�޷�{��\mc��x�5�{�:�.�4�| �{JD���:�)��z#��x�A�tμ֙to�W�g���:Ј�->��4�c��o������0��1�Ӣ;'���d��r7�
����ܮ��Z*��<Dw�BR��!�gy��R2Q�:�K�����M� ��o^�y����X��is-.-�U.�Im˧8���^'�ۣ�ոjp��.!XՉ�B��M�R�囏�{w���Qg|Cx
�V*x�Gyt�"3T.]GJf�x9ܙ3WJ��H2�λ#8C���f�ib�K)�_p�*���G�RuW=�>�;�U�R�U�%F�"����D=�`�oez�X�چ���iSv��V�2��m��x����$;���F)�9(�T �Un��$S/g�9g����%�A����(�5��r�:��̮#�NC&w Ft�J5��8���&&���V����TjZY6[�u���[Gn�f�|i���y��3U����GM�������$��8�UM�˒7=�oA�Z�����/��\O�Šқ�ݝq\�8d�d+s�hE�QU���
�����9$�Rc��Ѓ|�7LF�����ut]Lɱ�h�f��=��Vݲ38-yE���2�([K2�O\�\E.$��[����&�El�Ec�7r��߹.Q;�kZ�y���w��q����G��p�����o�m��A��Q&*xE��F�+.�^kޣW�$X˻QN5�oK�q(ߧ���|���/p�*��ڣ�5Viv�����8�p
�)9�UjzZ�ZٛU��Vvz���Cإ��ϙ�ֺs6�I���
V;[�1]gu�qD�p�.wq$�҇�h�Za~������"c�W,Ճ<����2 l8�ܑ�+.)f��XfZ��Ƴ�w ��א�T/��n8�̊�G[��@���h��Qp��j+���j��a�"g5�[x�ޞC�=v�7���)�u-�U������8l���xyw-�̈1��u���6�%�ʓ�����:Ͷ5n(�l6�
�y�oT�C\��-��z�t>֠�v5�<��J��W���3-�����'O�{�N�K{9�}���;��c�Gl�f�"p�E$�]?w����s!c��b��`��@iA��u층�7t��Cơ��:\p���]Н�x�_��>)n濷�8��7�	��;w"�ںQW�g{G9y�6��<AsCڞ��iW�9�܏������7�#3*��b�_�>V"�þ��#��"3�g&�M���Eo�/x�4����r��9��';;��ƒ�#�'psU�=a �Q���+S=��NSᇮbBTo�G'�i�e��	�9{g�Hd��N��z�E��]�t����}�{�6g"Ç��L�s,�WJ��G1��7�+N=��Ʈ�Ui�c_Rw`b1�\	јR��z;$�T�
Q�{��ՅX"j�]�lqO��{ވ�to"��Q;�����c��I/.+�@`)�{����%5s�2j:}n�s��A�u�������+ᵋ9��:��bd\�a�\�R���SKKe������t����wz�z(���`���'���x��g^?K)NQ���o�E]��pۃ5�,/۪�>�|o����;�]�}��S�(Ôq ��{��L'�+�v��\f���Q��dV�\�i��%�[���bO���'f�v�����}�a��x�h&i���J���gK��FD"%��ތ�5�W���<�w�Cq�#�����"��I+����9�O^��Q�Z��U�W�#�8�Sr)L#���o��n?�����j�u��.�1 �˒�i=���:=0�z����sU���ԕ�S��ed���z�6�^���O9bǢ0�+���d����ŵ����>TP��+V�W2�iާ|��J�Sr���Ss.�T����K��M'���N���@&����K�5�w#+���"�C���*ԓ��vދu�n���`.��[g�f/y�;�Nt��X�4�ֺ���v2��݇���<e��a�[%�,ݙ�lSӀfjL�j#H�Ɯ�%��i�HB�P{��Z't�\�s\��u��7ya�fT9�ʢ� �u���S�����B�N�N��(�U�3yO�@��3��v�u���%tV]�X�onlw�z�6���5����R�J��h�iN�ԥi�U�g�]^b0b��w��2���̛/ 2
��`�'�[�4(��Ry��.9��u�²�S�غ���t�����j�*���\�
��wtȷ���{ƥ�5t��ʬM.Ç"�4��8�\\�������i� "��9�4��r���al�4���GN]�}��m�n�	��X%4���x�NFܸ��}J��i�m��3��.�^�o6r�r��t�������dͅ�}�Y�_b�[e�r?�Wʶ��j\��������t�z�%ÊV�MP��L2�yoඵs*n�vl�"���#9RV5�mD���W^\}VێMv��d���LQp&��^%X��o-�nc��$˶F-kz�V�x��{9�t�S�`Vb��{���;f`;�;��@�b��X�6�#����!�c�X�a�G�G�x�U�o8Ҍ�-QS966�����g�y[W]1޻s�K^�y6��a�v�Ok�#�f�̗#��;@t�t×[���U6�������yZWVlR�.�.�'��ʙ�� ^D��9��I��7W;�m9�&6�MD_�~�7A���k�5�\��I��(��\����*.&�X�GMf%@u�)�V%al4ɧCJ¡�,��\��e���4���QIQeeT���0�4nR�����X#RcXc��f3U�m̨�Me�Ke`�sԬ��bi�ueejJ����H@�P�nZckE�.J�RfU��11ե@P�M&�B���LT��L�M%f��&	4���P
�L���0�T��-b�m
����L1�3ιկ:�u��]��mw���/.*�7���q+���	�AU�U�q��х.!/��舌C�E;�]��aW���.'�2�F�+��>�w["�K��[I��c��1�Ǔ[�!�&�%B��S�AE���M��/�
hs
;����.a��^��&�e\�#��B%�����Ĕ)�Mom�Ry����N/iu&3/zY�Җ�������{���-��\T�j��$ ��m���=��O�w�ٌS5%�	�6̬פ���#��rvE��m��(�:�=9�^�K��P��2I����#r�k"V�d����z�$X�;�=Zg*�:2�p;,	{S��n�eV�W=�Ԧ�oX���g�ȪJ똺y Z���9��}EMu}�(G�O��so����wT��;!�$��b�(^9�����V=����\����G�舐�D�'��=����,:nۍ}W�UgD��j{Vŭ�/�p��\�A��.`��L�λ��`)i��X�.c_+����u�8teqD�+s�֊u�s2dm�m+�u��)�0�E5~��v��'x;�tL����M,̻3&�H`Ĩ>�4.�E��u�x����e�Ğ�h�r�~��f����+CzYb��;F8�^�㞶WN�5.o��^+������5{��#�\QV9�qJ(%d��2Dᲁ)ϵ(ޞ\`�O�����b����[���N�X����G"/�ȷ=������9u�p�kT�ge�5�A*U ]�ܖf[N�g]����7�	B�q"b��.��E�b(=�2>3�q9�;莖ѕ�;;��Z�eF��İt�;60����9?UU�}�V�O"��f��
;�r�t;�Y�q���oC%�7�� �kMJn8T�\O��#2�'F�d��e���\�M�v8�z6�j8�FHS����vn�P�\4�Kv\��U�(��jP�MnݳwQE�N��9Ot���L�������W83�.��@A�fd<|�ޜ���Ζ���{�X����Vt�x��Jy����Z�x>��ǵ K=[`����o&z��Ȧ��(�W���r�,��<�-GN�Mnƃ1��j昙q=�|�.��diW��8vk;���}�~O-\Ri�j��/��V`B,v��G�2n��AgKm,�	�$S�{YWՅ��:�l@[��������%��2�	��q�-�q�:��+D�W��Dzf��{B�>*%1���{�-�A�[���f4�WJtIq=�i�"rg�Ps��.�<KѲ�!;=<;�*#9�}ԗ�'��x���.��F��>LQ}H���U�$�d�>���5j�cq!KTҐb��đr�64���s9���]c��k|t�R8����A}�=yP�t6��$�j�N�����ÊgFI(�*f�g� ˣC-y��,w�	Q��<����ƣ�;P�3B ��)>4E2'D^����m�ꨱ�<����ǥ2�J���-��k5|�%���/e����:�J�v�9��f���J�[�c���]���]�b{[Ho���g3�罀��ó/�kg*=�Qޤ���w����Z�p�����ut�|.k��
�����DG�q!�����^�Ͻ�!�'�OhzɶN=���C�N0���I�&���Oa:I;O<�����줆g�v�u��ι���Ǔ�:d;a�t��fI<a�u��m'2!�&�>C�) |�Sz��i'����'��N�3�>��:��y���>�1��v�}�|�������B'Xz��6�0�O����t���Hm��ӌ&�>Ͻ��<�w�}�y��8�	���0�<d�CY�i�R
Mr��O�6��M�zϐ��x�)�	3�F�yLD}1�?O������_����@�[d<fZ�zɫC�@}��|a�OY6��O��N2m��z�q3�}ֹ�\�Ϸ��t��|w@8�a�N�ߺ�!������PRu-�$�N{��d�O� ,�d�����=�7�����|���&�:gӪ��|�Z�6�g��I�V7a9׹8�V�8�I;���ORjء�d���7��~s���vq.��^����4��H
I�M;O��6�x��N$����4�k.��>��$�ot��t8¤3t��}�1�;�ev���'�����7>��2��J����8���Y!�)�	ĝ���ܒm�a��� ��0C�����[��g����o�XVN�l�d���$��g�OM����$��N�O��ChN��,ā��"��!d���
�.���^|{��r��ލ�{l�<|�ER�:�T9O�@뷀w:�U�탅�)S�(m�����x�7a2�8�.Q�at�u-�l��٫�j�ˊ�`uPė���D{љˉ)���I��^����� ���&��=d�R�	6�yd�t����|��d�*u�$:jd6��x�n���w���$P��N��H}�d��N�i�J�oi:��N��$������4}Bt�`k�8�f��o��{���3�o����O�t��i��
w�I�3vm�V�6�^�OX
M=�P6��N�s�hv�0�f�o��=��|���_i����$�g^P>I=a���&0��l=ݐ퓈hݜ|I1���J�g��'Oi:���������<����ԅCl�I�C�6��uO����Ld�h�!�����8��vC�M���>I;I���'�I3�ws2����}o߷�~ ���a�$�5ֲHe��>d>a����I�M���1 ��q�׉�zɴ�=��R�/k�6��~���Ϲ�x��q'ܰ�I'I��[0=̐�	�,��:�x��MI<I����M�@��>��n)���3O������I q�����!�d�V�[�ɖ�&�~�BVM�O5@�}}�1���y��
0(��`�_2��:�x�zϻ��O�wg�$����Hs����I�+	��6ȡ�@�� ,&Zx���O~����y�y�w�>���'I4��0��q>�>I8�����hOyN !��2L>��t���
�z�-	�6ɫ`5��~��B����v�8Ai$ù�#�q�.�6�M�mޜj��5K���x�9�ݲM�s%�܊�1�/z$]��ޮ�)RQ���ԍZ�t�*<B+&�e	�&J�_���z+J\}3��a?�v���E�m�i>{O���$�Ր�7x�<J��@�$�׸i��O,6�a9�}�l�y��{���y!�ȱI:I���=d��Y'��{@�-�z��ĨM�|�{C��X��N��(a퓌��������_<��;�^���~8�T�l���C��}/��&��'�$�z:�����,8��'o��Y!|��0�a��c!��>yϰ���y�u�%Cl>�� ��'���0��~�?\d�d�י'�&ӣT�2_,wa����!�G}�y��������
i b��>�M��� z̾��d5倲v��Y`z��M^gI!�������O��O�77��l�����ո��{�*|j��	�����5���XE��|¤���ͲV�)�J���J�x�Ofw���wם�{��)�]sλ�Ϸ��O^��d:O:�� �M�I3��q��G�C�6�,8îSha�i�J��8�Y<d��;��{�k�\�k������N����ô��:=��L�!�|��I���Ԛa��=���ms�z��7������$�.��>�}�+'[�ul�@0��	�CYa�i �!�04���!��Ԑ��ya�3苃^�9���𿩂�����i	���M���8�k�z��O^2M�xZO�'i��`M��I���5>�;C���Oz�Y*I�������|����V���vC��\{Ի�A�H��Nm�X� ����u���& �2r�u�	�����:�a�=kx�."k3ݰ��5}�Fs�X��9�����2�߻����L��C�N2x�㔁�3�x��v���|��N�N��OI��ْBje�3�C�;I6Ȁy}��dl����io}�xO���GTB���x��N=$<����d��`q��7�<}Bd�V�l'LĞ� z��Y!:����sZ�Z�������I���Ձ���fB&���$�zO,6��!�8��'^�|�����&�NҤ�P�Cԝxv�����\���߻��T���!��I�d���'�{��d�:C�ā�$��鞲N0�w@�$�7���@ֺvf��}����@Y��hN���`aﴂ�yo�>d���)8ɶO����������I�1�x��{��|í��7�٭o~��߀��f���`x��VC�|Z�&Z,���d����I�O���d�'���	�ɣt<}H���;��s�����1���v�q�XC���q���i���!�XC��|�$���<d����È2w�^�������O�k��O�>�1�}���YI8��Y8�q7�q�6�$�P�.2OY7�0�8�3ϼ��<����IM?{&=R'�mz��s�O)�<b�	ĝr�c!�^�M��5�!�2���!��6��x�a
}�>���af�/�|P���{���n=�RO���z��`jwH
q�;�8���1��&�q���@�0��o��ßz�=�Ҝ!.&:sy�#�8����׫C��w;�Ex�B���8��:����n=l�|���T�̵�7�\*`'�}"�=����xk�E.G�F��{�cr	����_'�8��		�o���y��c%d���Xd�&��I��Ohz�':��������Y��Cl�!6�S�`�С��O��:�����3o�c�?0�r�d��dY>@�&�XI��d�	�5��4��V�OI<�H���s[ᷮy����>'�:`)�����l��ݛI^�M�
N��5-�l���N$4e�i�&��OY&��:�O��3��/[��{��|Hv���$ěd����z�\�]ٴ�8�j{x�Rv퓫B�XM�;�&2`��_y���;�{��믈vΒu{dSS�&2N�t8���=d�'��C�N0��6�v��|��O:������������ε���^o_y���xH}l�����m��Y�Om<d��q'2����d��R@�����i'��n�P���;y�3<�{��?i<dY�>�ܐ���� �P=I���|�>����)��^�1�O�+�qj�UW��w�c�J�]9��O�A��-��xm{�z��`��>M��1��ʁ˱��y75�cc3�<�c.�Y�=l5�b�W!Zb�'��2����̤Y��+�?X݀/��bK��]yߒ��~]����o��[���a+�$�~�O%զ㲬k�a�[��J����vP)Nۺ5m�u����+���=_}���, ������o�ȶ�IB0)����ͽ��[ٛ���tS�sVߨ�KIVT�Kj��`\ 
�I�!H����k��O���@��`�|њˊ�r�.��Z����l<9�	F[��I�n�����܎����(ʽ]�L�pW�.�cd ���a�Y�T9JȀ��Pˊ�t���qz�6Y�If�W�;u��l��W���˷=[,;��%��̚6�$dG ��q�h)ͧy�:U�i����]m�=M����,:m�Gwi���׍����nF�dN�����&�Dj}ǅZUuf�.��C�
X����������c����-jߵ�cq���(a"�u���CsjF8�(�Nf�k�C�v��0��Vh�md�:��R�.0�pI�h�7O^7v�_ҟ�(�r쬃z=������9�s� N>��Z�� �����.��퉷PR�P�<�P� �����H�F��8Y9�M��5�u��V���-��t��}�cJ��*�R��vqK�6���ih��@i��J2����v�7���{�����gޛX��,:��<������<f��)/]u�6��eE��Q[׵8�V��n��dL֧SR�th�֤���3o;����Ք�'c0ķ��j����m^u��G6h!�|K�N�-B��o�A����z��F�{�"�$K�ڴC���F��c��:�r��M�@�K.(��iⲒ��H��<��,��%<��
�q�7�[S:����8s�ű:6�F��WN8��S��k��8<'KNBk��	*xkt�PJ�Nk��-�H�x�ޝM���^ʕx�Uۥk��۾�Yy�{)����Ԟ�gs��L|q]�HF��lKڹ4�L���[�2�t�s�M5w֖d����Ә��4A�)'V^m*W�u�e)�.^�f�YA�C�dt�X�͵�S���{�����r�5A
�佺�4/����cF_w)iL�Ju��F���4��K,rz�bayݾ8co��nX�V�o���0�&��|r���Ǎi5.$�[�<IMyiH�rs_�vf��p]�{�����:�f���w=aۋFJ��u�Sٖ���e�I��Ʀ��ټ<��+���3���5�V$�)3=�hښ.� +���i�vI�,"9�{Wy�\�@��I��v�Q�S��Vh���5-���B�a�5�̫Y��P�M+�V6�9�q��-��u�	�K �]�yT;��gLl��	��N�+5t�/V$^�^=�v����e������+;I�Hcb�ʬc��cRc%EYz�H��4Ƞ��ci1
�J��I���0d4��U�%`��T���L1��8�)Y�Zc�P�Z�j�
9CN���CI�Qt�!����f$�,��\`(ա���&��E�a�)�X��.P��
VT+2�H��fe1ҲV���(��$�1GYa\IR%[
�]Y1�K��e�8�3T�-*T����3�bQ1�Lf�a\ն�h�k (��E2٫[LI�W5��LLM$�ji1��ҋ)�L���AUb�&51�72\��L�4ӂ�N*���WZ��XQ3V�(T��Y+Ҁ ��*�?R�`��us�&��w�of�w��2�+]X�-��(�t[r2{+!m�7V�=���}�W��X�����^�\�cp���%����(1�v%lQ�,]Y��{��m�C�z�K|����p8PG�GKσG�
���K䯚��ۜ�=E�93���s
K�^WH���.���)������~o�a�q��"6܍�*Avl����x>���`�>C�B��e����mu����<��tO�>��T�p�ʴ�PQ���1"�[�k	a79�>R�˛�'!�[�X�*9Py�����.�֩,��z{��	 3n�h�|}f5b@�/M����(}y��u]C���j9`:f C����ǡ�%���izM�.��@�ܶ&|i	��,=e��۔E^�� <���x�Q�}؅�gΌ�ćH�i)e�KU��.�!��*���q,����Z���C��ǖ}�)�#�v�9EZ�G^��j>�qǯ�6�'\�=M��1����ǳ�(,�N�s�f03'4��
ґW���n"������׶�"�t4P�Z����BwSy�j/)d;�OJ�GxE��\��m�W��
?d@/�?�WeŨs������O8�������<+3�V�S,U�Є^�vx�=g� Ż����4ظ}S����o�@�*�m��U��w��#�I�O�kr4>�[�;�G���^�Om�5<�V�#�G���0mY^0-�B
:�&����e���.>Ҽ�	�����]�`�#[f�S֎մ�kj{���}`^m�Hk��\׃�^2��*xpH�U�׍b/�w�AO�DØ�vn.�ɕ.J1��k
��.�*�X�S�PQ�|��^�r.g  t T+G� J������ԍ<ᐆ[7�]�䝶�kr,�mC�y� �J��.��B��=�.0{ؙF_���[ʵ#����ܢ9[�	g5�`�ȍaR������B���o�sk2�q�bn��[Em5��0�1q�w�Y�f�c,�}Y��Je,�|7�B���{��N��)�����I�:\��z�22� ����4g*"?�������)�l��Z8xt0!)���G��\t�r�����Oތ�װ�F�=�k�dY��b"�UwL]0	E�ثSW�^���!ؿ|5g�V�U�_W�4"�>�)�K�؁V����%���۶DH߆�����j���I�YJ�@��V�<f}5I���컫�xW��"m��X�4|9�a�U���S�/{�;��~ ?�@kӝ'#8]
���뫩�*���h�^�)2�]�ܯt$iq�v\�B��?��w[	G�ǯ�R�β��Vd�=Ӳ�h��W=�a3���pG-��끌~ӕ�����E�Üs5ꞛcC��>Y��\�ۖ)CP?���ʥ��7���ks�oV>K�_��-�F���l�v�Ŗ���շZ��cZ��ǧøGƯ ��\�	83wh[͋#.*\���ҩ�� �ý�v��zvԕ��ty>��򾪯��qI� �,_�5 �S�%�H5�w
q�����E{F9�~��=���NE
�V�Y<N=T���q"���	F�h����{6����:�y�wm�����O\�́P�e+�53"���ڗ�RF��;�MdT��r�/lU�x�>
���\>&D�(Vz &�ͫ�b=	��vL\��}'z̹�FX|.z�8��πP���DV�K�������u*�/-�������2e�����f�=9G���=�*�Ҝ]6t����t��VW�XP�G�ާP���������x|�0��p_:ϋ��fuw\�_��=��]$�,�U+�.��0 �
���j��v�9�U5ŽG,���֘ww���
�G���x����6��X���rd�F!��ђb�la�;����9u�|��xT*a���y�q��'�4���K���{���rfU��;�o^�4�wN܊Z�v���Ե�w��}�:Tmk�C�z#�A'���q������R�WXK���]���S*N���(���v�~���>T�A?�W�?�S��,v��Ȉ��g5�>��{�V߉�]=���y�Jn���72)���L���ʻ�c|ۡj\n�4��==����\�����&����)��٦��N�8���V�;Z@�MU�:�`Ѷ�N`��1U��-���m�����6��'�3`CL��" 0����w7�z;����)�f*��V�_:�)�>�Qh��2骿[՘l��Ƥ�{ A��dm)R]p��S�m�F�|��X�!2t4�q5U��Ӱ�}T�>�����;�%T
�3�fzw%�l4��G2G�w��Ǖ,�m�k;����!�	�ʽ��w|k���[uJ�溔��֧���3�= � <���Jw^��jZ���{g��P�a�V���e�[2����o{M������/�z#�̧ۛ��g�w"���53"��A�������A#��-���b�wqܹ�ڨ�w�y�t���^T�N`8x�C�U���#�p��4��J_n��s��^�P^ }�Z��[[�1�DT��fj�q��-��06���5OʉU��aB	C�T r�BV�&���Gl�df,�AҡY�[y5�Wd)ȵ���
�[r�^0�Xa`�{jDX��a�(�u8�TJ����y���F�8 �O���Eo�!$_����{Py��H�$;иR�.ba��W�BƐ��;������ ��.+�qu�GX+	���YiA��<px<�e��J�L����n�q[5�^���luxk�~Lޗ񊗒ಞ�Cx��9ޞ�,y���ѹN�FU{�*oc���[�����5�6���y����J��仅��A�X����w�gF�} ��Pي�,ɩ�8k�����j��`��p���9��]�>n\˾�Զ<�ıɓ�N�{ވ���Mm���`�ȋ3yC��m�6kÆ��r�?dT����W�S��|�nWT�&.`J��qtL�rQ��]�UmCY��U�W��:�*{=9e��w�X�@W�>(�H�U�����T�x���m �E�ʇ��l��טF#�U
Ch�B��=�.U�=����-h3�VC�j�"��VR��!� �Z"�c�D7O�)�)�N�B<<0_��O?����
TOJ&��*neH�ݱLE�arll�����t�*�W:5 L�;L�T �����E4�ZCs7[N��@�����9V�MX��VP"���'o���N�x��vT�玱��vxT4~�ς�D�gb���� 	�Ϫҥ�@�yP< �����"(R{x�~u��=�X콋b[��guړڅ7�h)+�B�W*R�(ɉ�#�xo*�q�Ϲ̣���lYԹ낤,��fڽ����xm�*�{i��V���I?*���5�gz^��M�8> }�d�I��*��:�.b0�$��n�zy��=NՏi����}�����y��l��`�TV'��̤2H�W;9�W:���{��/v��[��p0���\i���V�nxD�l|h���0���X���Py<�\�a��u�柯�A�f°k�����vҮ�U���b����t5��r{�b�Z�;T*�ŅF(�H�3Z:n�k]o�7�c-{H��r������"*�DL3[J����пt�zʜ�����E�5�����ybVA�ƪ.�\�9�%�	UD
��bu�=�i�� ��P�`��p�p5=q���C����͢�+߻{�(��ѭӨ�ϯ_i����*��E(�*��ß�])�����u<�Q�����.Rkeh����@;v18�6���Y6���˔$|���Pլ���0��sV5�S�H�nC�Cc�*���9��՝99'����@U��5�x�l�Ń���?u��5:�j�x���É����L}ޠ`C� �V���W7���۬����-nE�<�u���L�ȑ� S
���W���W���..E�>w��ܔ �P�����D+�R	�)K�GקC�l�^����!�!�V�^�x*ypVW��2���].u�qos�[s!�o�H\�3�4�<�)T�����V:҇G�W��K�o���^�Wx�����S����0i�]�P���Vr����;��Ǿ�Z���R����_k��y�hUD˿r�,�!���>��
�~53]� ��j��uR�kWVt@�pP��b�{��,!�����T\�|���c!AU/>�O;ʦ0��5�댍p]���Cw!Dá����-��6v�r��o�������hU͚O=�E\�p5�Z�wIփ�n,�Ĺ�&�7��F��Jyc�9����� �	>������+�v�-�RgU=!�)N����TX�h��2��ڸ�'�A��(5`j0T����~��W���_�bb�Нu��� C��X��#�-�d�>̭uJ�A��S�"��n���Ns�4�z�0�]dX� �n�/�f	�R�_�o��4E)Ū':ٲt��t�H` �H0��n�o�Č�/��3�0��o3�ma���f�̄�Z�����TM�0p�hR>j`�4�����.�+�P#!�RA<���,�^��'!o��_v�'�yh�DU��-�'� �C��	u�զI�)�Í{��vY��qׁ�}h�,p�kTk��r�"��x���ޝ��{�eT�G`>"��/�]�Yh҇>Q���U~��~�[���Fr�XmoWm�#8�.zp<�뿤,Dƞpq��3�w���ӟ/�A��L���}���XrWSB}��YEpa|Av����#6�~��T�_jѬR�ޔ��XT����+@�tb�o3]ͬ�����l�]�uD��-ɍ�ק��[{��0��2���`�h�"i�*%B��&Z˥tCw�lѨ@�f,�&���s���"�g�3Q�n����c�P�Ӝ�+\�ht��A5��y�+'.��ґ�i��s�B m7Ǝ��b>�)Y���}�"��/�����Ƈ j����eR�0��hьA2h�k�R��M��{.Ů����zԲ�¦�ov]rK@'�PT������]�.��ӻDM���m:5eb��躟fj��+H���ĻK�CNளs�T�=->�4�i���m,��[��K�	(�.��@�
%#W��]i�\�j� �2�1�XS�W�X�o_��^s}3J������N��$keԎ���Bq�����WtҌ�[ꊬ�9w���nR�:�磆f](V�v���!��&n���K{f��ƪ�2��L�FM�:�]ͤ��X�DcYՓL�-���g�K� /��:�B7�7�V�fbW����|(���S��[���W-�E�W���|,r{{���\D��Z��yYw�J�
F�.�/��Q�)[/#�W��7���)q��Y���m����n��>���e]v��X�6*�p�6���[B$%'t���&q�2\��Gk:���Ԕq� ���u�����L$���ɵ�R��p�,����/U��_��k����V��1N7���5U���l✗
D��4k�Uh�o���VwK9%�A�I�Naur@�`=f��
�=+(t�2!��;Qq�6:6�J���6jS�}����EU4\�i����4������7VB*�ɩ�ە���y ��9mqԾ�͙��?��yl6�**7(��X�b�Um+*Ur�8�U�D-(�f&,��2&ZB��V�TT��ffaq�(�`��T
�F�l��b�����ї��Ze��,j�3&%J�J�**�n[J�FcZ�kP˘X�R��`fZ�*DZ�hUdU[k�%f2����2�m4Ԛt�R��J�$�X�����J�
�m�j[�U\DMa�"�eEա�ٍmR�cm��C-1�mV��k�fb[�2�"ۖYZ�H�U1hТ��Պ��Pj(��\əɘ[`e�4q\�EZ��\f �Z�lR6�M��j�WH�1��d�-��p�PR�-�V[1(5( �UX��.#���m�[�H�TE��(�~���,�~y�T�&"6w;&����;R�,jޡ�=�󚩶��� ���c�E'������yr�0�!"G��#z�߮ͅL�X4`���M�ʹ<[�{����^<;��q���
D���6���'�5v3��ɾ�a�U��H_�/�m�5/��vѯ#���p�������V��Ic�e���b�۴+���we{�*u����xi/a_�)#������X�e��
gI�w���q�9����Y2.�]ަRwr���"8xU��K�#���|'b��_���G
��څw�]��%wN6�`5��Q +���
@ �E}��_U#M��Mv�����%��1�-
�u֪�טF#	T)A��xjo��^�I!�8o���y<�e����X���!� A�F�+ߗ���{����΍xj�Gl`�0PM��
p5 �}<���[~����ĵ��b!�i��!�Љ5;-k]פܶ������w��[�����֧D^��/��]�|��i	�]�%���<Xa�af��%h���=�Dh:x&�MO�u��V�[Lв��*�5 Lv}�J˸2r��b������}K�_�YT�W5���˨ω�(z[�J�/�z�S���N7�<�u�4hS�F�nꁮ���o��NCM[OMܒO^{��m`���yP⼕*�¸=�Dt,���	:���9g��y� 7���,�^���� `��W����^��O2��އS5���Bo������+�{
����
�X���y��l��6k�ݔ�im��XΜ���S��W*�<n��_�$`��!<`ѽ��V�y�S~	^�=�0�(%x�kfV�)U�9Y�*'�F����`!�W*^��0xՇB��PV���*��<닉d�o�	|K���T��U���Γ���H*1@x��� ���<��Mg�%n�XzٮY]);�]��"_?>@ᆆu��0�r�K%�Z�dX߰W]�v��6kZ�E�qJ�:�^5�Y�R:�a-����k'\(/���,E[Z.s�C`��R�*��{< +��"��w�sqW{ڑ,R�	zlJ�$�F�7Y�«�wW��5��J@���3��ˮ���� b���Bo\�����OZ���|cKզ�]�2=H��(ѣR(�y���~xʁV�E|�����jڝY#���G�������pt���ΜOi�'��W���lu*�������>ͪ���|~ɜ�>4�K��o��Z%�^:�8x�ʳ���<ߦ�.��ByR�R���
�H ϯ�\���������ށR�u�Uj�V�����ג�3�㣉�H����	�;��\���è�{|.�_�{�uђd.鼽���6z�qx��Wƅ_�8��u��J�rF������2�U�[�������
+��m
���!Ժ��Z���x/9Z�:�:)�Vj��96�]Nʒ�X,��70gU���'
����TU�M�sͪcF�pچĬ�sr~����q��'����G��v�n]pw�ӡW�8�?$*�VF�a���4��rM�)��hp�޶1��+ƺ�u,�����;�y^����w4=�"�7�8�N}����*j��uW��p���j�������J,�m����=��'C*2��7�"�@v4���m	���Aj���B��M
�jz+�i���g�]@��XxTJ�����]	0���90#q����wY�aę�rUNu�K���W�L���r�Ӿ m˺��|�M�^�GʬQ~l���V�@���*�j{�5/o�뇮�.�>g�?5����g�Uˠ.���	 c�4p��~���m���p��z%��;^F�W�s�լ��.U' 2�$�D���1��zʳe��]�����2��K7Ij+��J�\���E=�P�M쨯h��N��м�)��ʎ��ebG��X�U��b��staj�C*�V���=�PE[ ��x����R6 鴭�M*N��Aa�C\:_�D���v}�K+*�b,*��&�@�Q��z�sR���m�=�{q5�O4Ec�A�!q��^�� ^0i��VpJ{��=�H�!t�p�î�8��S*,e
�X���	W�4���kÞ#+ʠ��EȈ_o"/,.�˃X����MU��x�Ęl����q��g R����/ގ�a�'|j<��bY�N����o[L�'�r��������u�^s[\k��]eѯi�S7���~񗑜!��ޘyv&��r#��Ƕ�Lt��ʪ�\T�M|*8+,j��}�}� ��\O����S\�L�6Mw�xh���>��������c�c(�"�b�`������κ���,�U\�87ޑP���0���p��"F#L#�zgPI�q�\��n5�u�V�/zD��)�}��.���늋*�&��G8��hSOk+0��G�#"t�8�H���39s/3#2���ps���f@��X0:�B b;��[��y����hX|�[Qo�WLTP?��+����:��
�
�։=�Q�)�{��4�/���A��.�3Ɲ/.%��[2d h�
���M=ʺ��Dz�:�j�7���X�D+3�,S��[x�neT��� �6k+W���<<�o�5Uir7zzJ���ȊѶ"�wu���&��2�UB�q��S��=�X.��=�$x�U��Z��f*g�vTP:����x�#%^�L;#��ڝ�.�%���pʇ����ZxW[Ȉ����A�|"�N5��&cCG�N��|9\lpb�9�r3��VD4<7ƽp��q�b)-��..�Rڊ�t��C��\ U]�!UP��c4�;��Y۸��$/P^ �G6�;0A����X8�
��=�!�.S�4��<�y��tj�=-a'�K�-��H���[fm9����&���T�u)��+zL�weȧt�?+�ǲx,�S��fǆB�r���H����pG-�K�}ҮE���h��n�H� @��p��U��zХ��]�;�l�oGz�p��� bj�t@�j4x*gaZP����痛��=k >X�h�hvf�\�6�D�+��6�Օl���4Q�[m3�N6�V60��:��P&O���f�)\�͌�/`qZSZ�q}a�dP{p���>�U�3���S�)��<(S��=a6���:G�V�d�Lav����k��>��<P=N�wSڰ�~��n{�s�.�4~r��ET�=��<7�� �I"�I��ܝײ�������yE�_�*���t�Ӊ��� }=�=��tq���z�'��c���>4ܰ��B6�� �Pv|z��f<TPH�5whPS���Ks�����o��,��Z�p�.wW>²���tۢ+i%ud����.����t�1V��tNX�u��:����IîK�������=.P�nݖ�NW��{���{�ڦ=���g��1�oޱ�D�@r������o�F��:�H�y/��㕧��e�&1�M�ݝ�����@���8�t4�_<�++��]`K�(��e��8���a�X�6���Zi�y�R��Q���]z����G׽�z���dD/�#x���Y�PJ��P��"�ܣ�aH���bV�+}�� �z��~�����Sӛ����e�A:���ri#��6Mzz�;����Ɵ,���u�B5���!�D6�f�����۱.L�}����0z_g�q(wYs_�ߞ�=�_�� B mb��V�#�ꧢ�C�R�C�6���p*B����*F )��jv�8:�[Ơ�$�.ό�9�b	�Ʋ�
!���q���ȳ�fVub/2�:���p�s4�j�G�\kd������\���h���7|��,qU��SD��]��rK0���-�I�Oυ�\�w�?g<��4�禣�����vL�^���Ҽpj����n�'�$=OUq5­�d:�"��Bڞ�d���{��'k~rl�;�3�&3�.��.��g Z��P���z��ZwD���u�<�܎w޺��@��%WZ��n`T�$e��P�/:&���b#Õ�U�Z�h!��Z����+	��[*F���{7�~5�9�n�#N���p4�W�XP��<B���ADT�y�����&�%�\�㎠<�֋�c�Z��V��{��6�<�0Ue�G�<�vt�HO�`����޺l핦��;��vy��Yp��=ʸ(x�DB��E����Jkj�3Z\�h �e�Ì����.�08\<�{�+�q+Ɛ֋����H���]K�oN��c�J��ֱJp)�1��cc�X�v>r���k����oz�kW��Cm��˹ݡ1��w�!���	0�Y|�ٔ�2���5H�_�;O�ߋ�A�C�����w;��@�%m�V���+�����Wk�]��f��2X����bWz)��^�*5���3�\���3�zD����@�EY V���ga�is�rg�91ǻa����&X�OY�
�L0|h'`ux�9���q��:��=6�u`��K�e;�����q +��
@ �E���lx���Ie���	�p�WLTPj��i̠�%/��,�@�7ّ��/s}�Rz{�
�<i������7��4��l���\�!� mV	~�=Xލ,���gƍJ臟e��(xxj�p!�a��
TO�Ajyg���I�W
�h@/
�n�j�4�\5�5�!<�]0^��k�=Љ�b�ŀ(J(�;(yg�z��j�M!C�d�Q�����k���+��(P���{*\�|��;O�KV�1�鲸�2'-�=���v�L�[�{�x�9�v��Zt����Qב��0j�7�M.F{r��k[J�nH*9XK�t9�{B܅r�]#ǌ����u�'�;�k�ܴ���,�B��޷���-=���u�^.z��͹e���qr�Ab�)�$���Wc�IFq��j1�f���8v=������=|�v�,**����<��Y�P�[���5���"��⮆�}��dwEp�'MַFά��O;���-���;�s~���T�)>'i<�ܵ�7nv����ɴ�����S�s%��^3q��
�N���r���],�B�I�wZ�}N�Q�p����-��5c2㶨F��#+-�[Fw���+�ۢ�q�W��,�)��:r��Mu;�=R�kx�,j�Ֆ�GXD�mG)�W�if��\�{j�n�'��f�}]qh$��_c�0梋����r���'�Tow#Y��,p������C��h��#rs��]Z�>3p��yS7n	r��W�rp���U�Å�nE��+0c��ՠ�6��5��"Ή'`�W3���&���Q����˄n^�t��q_J-g��4^�8�PN�0nE՛HnB�钅$��M�ج8GH�=�;B�8�w��N�:�ͅwV��{Kj9���o1�o��)�*�WC��u��(m[����ҭ�B��(�ڵ5�-�S-wNhH�3EЬ�iҶyOe"�vV3S�W��n��F,�X�V1҆��b�fl�ժ��V� �j�N.bT2��:����r�Gtg�N����x��0�D�i��<æ�Aw��+���=�|��oE����[�#�v:Öi�g{�%Z����o�ʠ��Xv���q�ouG+FE����WJ.*~8�'m�s��ѭP�!w6����|Dr*���xUaQ��o9�q9�z��zts�OhZJ�ٯ[|Ot���UF��"���6�.�\�J���d̪-B�*��V��+1.�+AIV1u����X�3
�h�*��q1&[Q�++*�D�1���9�el�R�Xb�F%�a�f�q,TKmB��R�Lq���@���I�T��4�q�Ŷ\ZUU��-k-FĴ��.d
� ��PK�*�-Z�.�Ɏ2�j�1m�1P�P�D��\Q1��%�T+5��6����L�r�bV"�Z�C"ZeS�������֊#-��-(
��Z̴�m+&8�ܦ�*(�iLe�L*���j�,ĕuh�b��S3F�LQ�n(|�?Z�Ad=���3h]�fĶ�^���/1�RvL�j�WZD��oU��R�D%���ZBo��g�*]v;����djTo�����.&�a^$��=�/;}��'�hӿd0�ω�SK!�01�}�*�~$P��{��:�e�=f�*ӡV5��
�'(�'+�"b3h� Ō�ϖ�(q��r뙗������U�`�]�������~ڷX񤔃�]׫��?V�� �6�ΗQ�3j��A#љ�8MN�׺;��c)�<���0"kH���i�$�pk3:��nN�R�x� m�B��C�갦A�5_/��]�/x����'���-a����h������fN�!ƃ�d~�x/
 ԫ&\T	�[.@�cc" oz���F���H
��0|<��v�-A>��u�3to�r�/����)�u�x��྾�tq5-<��YA?K]|���nV�����BV������𚷜�ґ�� v�P.+�����7����7r�JV��}�7'���;��$�B0G���#E�FoyH������_'�>�~��|�Nx^���D�f�Ko ��s
dЖ:Լ�G
S�Nm;Ov?e�Yz�^�T�Y��5��X�56�g��'��6�� ��6,��,�O�.��t0S������>��a���,U�Ͳ���,Հ��o�\;���a�Cur�ۘP��tenAh��J��!=A��Q�(74c+�&$��Q��E�0!�󺂀��<+����S�G�he������Sʅ"5]M*�ۿ�����]	��@�^"���ORD�$|��������l��Aj�Ve����ML�渵T��m�觛�������h��V��[5���R���V0��*A��;�+$�hU�q���x��ŞuĪ�qTm��=��u�o�(�t�`�����7�g���b�5�����T���QR"i.���ge��w]yD�s��S�j�y����G_۷X�f���v�H%Ȧ��{� �T,΍W;Y��u�3�_4�$�e.�ս[v��])�I�_TE��Ovvr}T}�:�tU1]�u񪙮��*j��uW��=qp7-?gt�.��ǩ �w�/�
�}���b)x���~Uf@Ge������'��L���,y���I��o��G2�)�r�Iމ�9u&�P��i����l->*~�ϧ�>�jo{͊��b߻� �hA�w��*��U2�=�
)4�Pש��M�Kʃ��=t�Y�s$p�� !�����ͣ6�ڣx� K�3�!ԥ��.-�V��A5������ɵ�#.���#�|o��:�+Q�'\�I����%a[w��!�&ƌ1�e�]{>ۂ�hظ@�Z�&]��z��o�~��4�Y��e�"��>�P�3�>
���xn��~�[�W��E��v�GV�����[��q�I�]�FU�9Sn��&�6diV\�-�֛հ��+��}{)��;��J�ae���'��k:�AN��RA/����/���ɺ�D�Q�Y���u澺E���^�cV�̺6�:	]�w�eL�w3L��;	��w�/�\����{�,�d鯻<��u�(�XB�9�l��#6��,{o�V.�tq��,U�/];����T/���HR%�֋��L���%=���Z�ұ�E�$�����s]\k��]g�:��թ͞������*��\`��B��+�	�k���f��(�����ٛ����U���&�}�|)���viW7p��ܛ,]#��{vrpҝN)��8]D*�
��L�`?	�-M�8�)%�/)�j8V��:��K1H r�
�Hw7����G�#&���6��#N��ܿ#Y�4�seֻ���ǭ#=\pi��pO�k�1�u�ts���_sM;�՛S��9�ɘ�nW'�L��Cy�R4��_<���p��*|D�Î��8<�6\+����,�WˊE}�G��R-7�g�ʎ��{��Z�D�Y~4|x�f��C5ؘ
���� �!�4��&�����</n���y�4xP��坅ct�����)��z	�wc;��CN3^F�?qX��޾���/�z>�lw�`��U��0V�:@�0z��s����5zhyV�h{|Q�c�RM|_�u� �.����F�C
�2�j�!�o����e����I�H����F�>&���t����z�>�]�Bs�����:#�a�f�*�Ƽ����'*R#g
�}�"	�92_����!v`�8��Dc�Ǽj�@�!�x<q:A[}�K�Z�Z5�׽�L}w��P�׎x��\��b�Cnf�sT��'��`�ł{�=�ӪE��f�Ĺ�����Ewg2ɷ0���)dJ:鄄����lE����~�=��� ���z�x�[xu�p�3u�V�=b�DBѺx�<0؝]���)��!uմ�l���ꭘ���|Ыf�N(Oʗ�N�@�dٚ�6�܉r�ld���G����S�*)~���VLb����J���η�O��?�������� �p�9����k���q��֣FI���@PM�5��x�og���D}GU#���&Ծ�Rn�P���.����:���d^O%�zY�)L��/�F�;~' ��]p{(�#a�0{�����6�T�/��$`�E
��F��_����`2-#o�{P#��O�yPU�0S������-��fz�7'y�4��B`� }��c�8L5�>*D�S�SծCo�����,P�<s��/�y�p@��60+4w�ڸ���P�_^�]�Ll$k�n�yN�� ω��Y�~�U�FQ�U���gײ��7�A�N�e�Cv�4Y�E�ox;u��	��9��e1�{�|7��(��MGhGw[x�5��p醴�̨�K�vZ���?*��񽓧��Y��Ɍ�������E񡚠_c\)��+����3�Rt\�-�;u�F��&�F�4+]S��q�a�*��L�>��ku@=�e��pk�\�a�!�K)��?ep8j��k ����OKyM�)���}��s���y`y娻��-�5�X�cm�9�׶dO��q���!3��=�����,�	��u���KC�y@�Ύ�-��)ض�js� ������CC��}<%2�:�i�h���&���B�z�Rc0��GOpN�]>�*`Kb��԰*�v��SU��| ���k-"�s�:�-��Q����n��:�z0"]]T�>�"��]ν��Gn!E��u�
�*��AG筐�"�@���,L1�9��3�a��y\'d�^^�g����$�����`�}5X�������u�;J4���1:J9d��|8�6�%�����9��%v�ST�z_9'�����rO2���Mr��Sʦ�����a�5p�����[mn�i�v����;��A"��dS�^��R���p�iSs �%W�m�n�\��$��0_��B�!�i}.��Jລr�g�|,�R�;c@MY�s�&c���,�tE+0`��_y�UXP�#4/=�]YL�O:�y�1V$<ƨMo��X��:��_]"�k� ������97,W�xx@�
0�E�0��Ȉ���1}�<�r0�/z^I����U��pxWBF�t�]7d])doh�>�~vV{���tr�g�^N� i��U�{ݕ��&�E"����/��7Z��[~<�`�xtF���Ҡ��pTRb�2o��˪
P��è��w�\`��B��+��|�i���y��xp$]<0�\��v��RR�p�B�q����Й˴j���%��iF�@[}ԓ��rR2>;JkD�ou�'Ե#�(��q�]��v��$��7:QH%���7�O��xr�7>��tj�D֪��
<@�eY�p����p%��R%�<�N�(8����B�<*����؀J�m�nqi"6s�v@U�\Q²4�,�S	,� ЃhRN�o6���@ Vqa�����qmM��5����k�$a:�����=�����F��X¸vQa	�J��e�
����b��	!	�yl�6��"<�DP�r臙|<3�s���J�h�ȀuBl4����8�s��󂧁8�Tb�t��t�7{"��[���Ԝ@/,NR��s��˪�r�T��@��������v|M1P,���{�[M��Dی�1~����R)`�7^H@��@*� cF��za���7:��qlL�1s��)�U\*����v&�(�f�wHAPw�YuZ�46j+�L��-݊(x?{2�i�̡���������G�]��vWLSR�	
Y׹�Fj�0��i��\�+!Dj8w�)y�m!:���5�ɓ�G?+���D����\p���Z~��k\�������݇-�g:zz�6{�f�B4��^&�e���_�h�Yq��f���޼n9���3WZQ4�,Տ�ߞ���.*�$?9|���5�Ӧ,��,�C����: ���V'aӚ-�'�#z�b-6��n8ܹ�<��i�ӕx)��\ b��:p��Et3o����z��.ү"���q߼~Օ1�F]k(��ubǒ��˝蟻X�_]Y< �I��A���R��a�W�O\��s����y&\����K:�U@*:�������u���N>�k~�ޞ3B|�{�a0?��|M;�`O�@8��5�4���)DCx痧Z��w�u��Wz����4h�I|**���(������:io�����(V��<׈E��B�;j���uy��9��WVRϧNጥ�4�����ҕ�v#C��9%��j�8�\�����ټ �GN�o�8���|�g3.���b�c�]*x:���~��X4+W�j�]�=�	v��-��6>6��Y;���!�gp�e-�\8fB�娮����*�Ȫ3}�Gd�eY!�p��Z2�)��ƛ�)�X4=�εZ)@~cϷ��O#+t�D���0tU˅X��K�+$��	Jg�u�u���>�y��4��V4ǵ��:I�a+����v�E�ŗ
[�i�>{I�D�A�9~�&��(��u��y�F��.��<��86Ҥu!y�Ѧc����1oG�:e�UR���V��r�7���Z����EP�+R��w�5d��.2	�VB�Iqi�w�).���v����:������\�Y�@�s��gL�Vl*�KgMD�{��H�����U��\�
�^�&3��*>P^miT��ͻ]u;2�m�{/+;�t4>��J
GM*S2>gsS��M76��.n��8�,Y%�Yb��!*fon�);�n�P1�u�Q�[�/3`gwJ�7.8#�B󹆆+��j#%$b��Vֱ�Ʒ3�Wc���s �OZ��E��kjv�pe>�X�
���6�nf_b̑��f�<IP���0oV<k���Ү7�'��u3���,�))qu;N��[sC����i�0�T���s��层Ryǋo��al*3�l�7��b��T��jX��6�*vp��u>�%�V�}��O.˂m�<��d�/2����Y�s�ю�ڈG3N��בIl��`L������k9��p7^�"�����N5��k�Hq�d��sr�	Vm闓o���qk�n�zGZ�ʇj�E���R�ڽ�yQ�݄[,s	�\f�֥�G���Vn�m\y��Uj�\P��2����E�[ٲ��/�-n�p2��Q3�������)Z(��]��w��u{�<��^
�5Lj��2ʱS,��J�-�J�(��kc�TJ�rٔ�mAQ\�e۬Й���cm2ԭ�2��.c*�b�̕���DEj�+X��UEX��R�9h���K�q�\�"��4F,L�Z)�T�2U�� ��e�*
�D��rƕDA�V��b(�b�(�T�ł$P�r؈�1T1U`�"�)TL�C,� �m)1V1���TX��QDUUb���MZ	���#e*"��P�fR��"1QQQE�(��F(�5�,��E1����AX,b(�Ո�Pk*�F#�*�("ux�H�_���1���mI\)c�鶳�T�<k^����EDŊ�B�R?�:���3�e9�F��O+R�p�P��1��P?�w��rr�}�3}�ǧ�|7��ʋ���¾QV�@Su
�kC�_��/7���,O}�
�+������"��PX�kz��Ņ�D��bs�0+����÷�Ʈ��N�7^���d����TZ������Kg�D�q�ug첆�8T��K�{|.�\u���<�)�F�e���u�j�#H#�+�*�t:҃�jA�-xg������+�P��_*�Qv$$N%ڄ����J�s�cx�y=�n���O�+�y�AQ���{�[��W�*!��v�bw�yn�ہW��C���һ����S3�T?{���d_b[��(������㪖���\��4�x!Iu�׾5�>�Ӑ�X^z�ML����l2OG[MX�ܽ��# m5Kٛdۨ����7���5g�V��a]�X��!2�|���狱�y��ʊWE|e�8��>�?nI'�b~T,�^6,�W=�e� �W�څ��Qڃ.F�A�3�.e�U����R�[�#�]���
xW��M,,�;�q��L��k�D�ۂ�G�+��XXmŀP��>��"q�K��k�W��S< ��PV���u�U� c�K&�� -��^�MMw^��%�R4�H�@���=���S&|�LUu���F�J��Q^�Z�4g�V[Ľ�8����<���D���`�T����*���(/�˾��*���+�{��D�U����p"f�G��F��B�49W����%���cFP�
L���&�����i*��|B�uw���~��HP�_C�cj Vx�MK8T$*<���7�,f�C<O�U�v����j�'�,PESԜ�@�v©��]���o��ʸĶ�e��Et��#�v2���7��[x�31�,��%3�xc�,�����A���}��Y��(h�Y/�=U�_�"4 �ћ��*ޙ��$�4+՛ll&~���R�  �	�G+�e-F�/��`V���6�7f�x����4P��Xj-H;1A	6���-�㞎^S�L��\��#ƶ�]��/ǂ��]�gF�SS��o�K_|����_p��lT)vs�{L�L�Mb�y�MyS64�>Y�s��.��ֈ�ς�3����QvC�L	v�a��v.in>lԳf^�O�n��U{�+)��u��������3��j����h��@����
�w]��ת�5ٕ��(.�2�[^�N��@P�)C�	{B�C�J�@��1p��S�fnp���Uq�3N���M6hќ�������V.�|Hh��u�V��G�:��}{�Ԡ*�`p���O҈#��H{�pe��j�k�ʌ�v�M�O\%,���;2�m`��-���a�[��9�_H��0��?��dyc���P�*�f�PÌז�w��M��H����Kbe���iK(�藹��S�݃�����XMnUCʡ��t�c�QW$ ��`���؍(_��g�lF<���ف3&�;~�6�@�s�t�4wK��]��W��®g��఑������x� }�#��߽'{$��Q��G�J!j�Ռg��ѤXݘ�><�yȕ�>��a�kC&���H}�}�jjcj��7X�t��W:�`��O5Au���c�|o�r���6>%,w"��(�v��8�R�ܗ� ��W����T�^�X�Ƭ:*���P��JL����(�у��quiW���4�}���_��VS(�~���PIY6J�Q�yC}a�Kq^�y���9�NCWԩ�p��Kg=W]�"���b.��i
sz)�	�H)m�T��e�L�j��g=&F�s:޶��x��(֓ ��ե{�)��F3^D�è=����D� {�k�eTlQ���~�r����#)��l��/~�F��������i�K�bɮf�f\FĽ�\>�8�7�km��Jp��h.����23�f���[���Vnn�l Aj��n"���iLFCt���ÆT<* �/��$��ї�=���^�:�S:<�'R��f���3vx|�Ps���Q�D�=G[�ޭ����ׂ��e%JǜU��k����6w�� U�����c5�yQ�?E�@p/�o�'���Dƛ'��a:�X��՘*���'�̞٤�ZZc;�c%L�w2��=�
���`��Լt-6:`ȗ��*�]�\�Y��Pj�tE�.����cS*���W�_4�����}H�Μ��G]�r�z5�l){n+:���=�2�Y.r�M�N�]qJ���6����ۮ�nAW=`K?6j3��H�],�`R^�����hԓ��(Ou�����o���+�3��]U�b/|�ZՂ]%z�>��֕�=V�/��];�2�܍���v�	����r�	f��ﵤ����Q���%��Wᢘ��4�J���:�*3��0u��O.�'��������k����G�	��sn÷�H��ǶVIsE��̌��o��!���\��ia�/�/���b�}0���5ь�@��s�m�\*�[jn�y�������Xy�-���z#sG��=������>
�5-H�Ȍߧ����GF�k�}�eM�\s�+�`�k�������%x�ˠ.��e2A���U��~^�`R�
���ٛ[|&+��U#G��?�k4D��@�C�pZ������i�s��ǝqJ�'��$w����x�DCZ���3^��\!�z�n�5����)��w(��Vl��y-Y�M�D��s�Y�擗:��eA�@a�8p��xR�em��6��?���zG2꥜MJ�`W�Tx �ˮ�Y��,P���A���cjI��C��8g�yy!����FZ"�����owb��޹ޜ��}B
W��A�B�d
�b���t�C�Ά��(P\�m��yи9׹YQ��L�s��_��\<R"�'[�
w;ӸX�
�*�\�Ƒ�Ǽj�4@Ƴ�ùufV�Ȓs֯+�j~wL2j�Ϝ<lxX�5 ݮ�^]��to;��=���/a�"�f�ɛ�Ϊ^W@t,ux�{v�I�>|�j��X���lY�0���;�&6b�cy�3�ךN=�mp �	m8۸x����hgRؠ A��/�?�U�ڍ]^�?S���I�ryPko��"��˪[R͍ңk�N7��@�E
����ظ�2�WU�TT^��2���^��ЎV��f�\�{�D�QK A�*ۦ�T���k�ϵ�L�����Ā�����g��ӈ_��� �����_R4�.�ҿq�f����9k.L�8���E�0B��	�qFD��-�b��Z�ڜ�Hm�#���}�����Z�DP����+�㢠�/�;��5;��j�9�����
u8 �\�Z��6hY
OQ�r�z���5~?0!C*E������1K(�0<�����dY�)��KI������kH�?�T\���� bʡ��3��B�C�*Tq���΅L�I�ã�,P��֧V�,Y���`�d���3j<$�ë?�3{������X��qj�vV�*��GU.�M�˭T���V:�ʷ�%�@�6,$�{@{�o��1.K	��O�<���$"	�ݻsA枧������l��s��-*�y�[j�C/�M�������p���[���V(�R<�97W =Y��;���j��ka8i��{4e�~*v��rm���r�q��en��.���1Y�&>ՁX.t��}�������օ*�U�׵A��^��_Ё�����x��6{�_�U�P�Й�.�*�~������v��ZyW��*�-5����J�;�E\n��`_Ƹy@��2��/�4ĕJ��EK�׾ۃ(�4W���H����Ǉ���ܫfb�hVw0�g7wnP��є�d�PD�y� xT��Dyx�SRlO�EX���aB�5����#k�ӟ4k��T�w���g6�������~�Ŋ�]	f�z���+� ���b�iR[ӽ=Lz֜��"=D�z�pp#~&K5�<j�粼��T"����y��) t�S�ip�ܬ�}��l��3ٷ±n��n�����<l����`�)�K��s_Y3*����#��Ŷm��{#�ú�����5��Ck:�v|U��껫dC�9��ߵT�K�?_��c�0��y;3-W����)�V׋����6	�S9.#*z��������*���P�v|*���K�w%��DsÆ��zE,{2��x��;(�wd.�ql�9/��ԼtM#�+N�Q��szǩ�|�_�*�@.k����}aAԈ�S��VMq������o�vh�.n���?*�?<��¹���+�����Ă�Jh���R�..��ֈ>�R��e�����k )S��=��wܳgW�����*UQ(�f��X�E=�r;N�?7��׽;���#�Σ���	��AQ5���G �j�+�atˊ�>|�C(tڠ���KE�f���5u�"�>��v�Nng��mQ7���a����*�Ym\xA���
�Vd�fV�L�U�҇�"�m:<���v;fE�3n5��>1cٗ?47����z/g[[��E'��tK�U��m��\���9���
64����բ�i')'� X�E���iyK�#���*69ZQ�<�7�&�E꠵p�V���{v4��=�� ����/{P�X@�h�M�+�{"ꝑE�0��H�$E��ӱ�xIVk9&h�َ�r^�}N����v�O��M��yPk]� A��t�7�������W.Avd����Yt ֹ���)B
��U�e�4�v]�����B�쐌R}�[*C���o*f���-紖ݮ.oj�e�LN��<�]΋E ��Y���w�Q�����W�jq�i�5|�XJ��	��a6���j�[�0i�>���P7�ӦL3�W�4�w�t�GpBo-�\�;��/{N�U$p�G�[�P���ⶺ^�i�1�-m�2moU�K��9F��l`{���9o*�k�`�\s�q�`���wLy4mr�{Z>����ƪ�f�MI����Ul�S��Ws���:�\��>��1�1P���Բ+�a����#j��fd�Jh���;�zG]D3i�D�ַ����Զ��عV��Z�M�҂�F�ᮧ��Y5�ie+��&FVI06Ĕ�1����ӳ`6�_N��]�&�v*J�;��voC9͸������u�q�u�eЇ��d�ܜm
��e����4�+�ia���nEME��wT�u�CNm%�+n�ХeHnnl�I�w��bP6=�]���҅�ʅ���V�o�s%���1+n&nڋ�<{[���1Cx�YI�;�ȴ��Nt��Hc����b��rvS�z�X@-�Mˡ�]̯��eަěXy������PT��F����m5�F��0n�L�1H(s����O1V��r��n�4���oq4�Kǳ2>یN"�S�gsXeJ͑ȯWuh:�D�����R<5G�� ���Eb
,�TTV�TEdDEX��m�0Q�E"0EPQUE��EDF%J�VVTX�Ub�fYA�T� �EV��QV
��TUQEQUhĶS.&e��YR�X�PE�Qb��TEQX����UFV�R��+Քbi,c*Q5jȢ��-���	(���("������R��fR̴*�(2�J�A���SDb�F[X�V�VE�Z�
�X�-DE�Y0`��A`�(�ADQQ-��=�|��Ǿs3ח=��71?���dSiR^��(�X�_o;��	&E*��R��rt��i���
_�ؙJ��oJ*#��
T*���4�ǒW��������@W�.��{���V��2�*���CȈy�^��}rN�>3qV�]ج����:��D��t��=�7I�{�a#�@�ZXB�2����`���h��u�V�ҭ�F�Yۄ��=���ӷp��2�K( C8x]Y�:u��V���j?v{d��%\�O��t�ml@Vб�L�Kr2�3hN�9[φM�� ���Ǚ1(@�I��+��R�^��uӛ����e��#}S{N\���R�;� QF�`�7��{Ȉ��I�
>��v$z���E��j#�z����b�K���#Ps0�b����[~�� >ap��x5����4!��X4 ��s��,�_���u�w���|N��Jk�W$Ȓ�ޫu�t]�r���
�,�M\��hk	j�g��l�E�����X����lZD�O9TS"���;"�%͑��J��Ds���)��։Dէ��E���
�����4&��'C��6�B�r6a�z�"��_�����gOOrx�yY�{L�5��f��R�b�M�5��Ơ�Sǽ==�:C,�ү?��<1�L�t��d1��sB�?O{�� �|Z���ۦ��L�"�����rN�	2S=�7��83�� '��Xc���JbʙT����lKa2���K�u�/.��P�5n��P�4T�,!�J��O(�]���N{�X��	�4�_�� �E�(S��k/��P�r �Hݽ~��bǅ�Y�&�y8pE�L���@�%z���q*�S���	��u4�2s�#��Os�;�*V�
���m�j��dI3Tm���.d�*�Ļ�����5{��r�|�����m��<1s��|f�v��k�O$֗8�m��ĕ�$�I ��w�#�MBiU����t�c�QW�2n&H]" �6����.2dVeNQ������x`$�Ze��(")���������׾��xHH���Z�Aνh`C�8e� ̣m���=�F��)�Ǝ�,�
�eU�5dߌ�T�qX�ͦ뱽~RG���� �R='�ɭ�e�%��A�z�%5��xe��l�E���kt���Ǵ���c����?#��P�X�H�m�3|�� }�-f����i�Ց[���=�����5E�מ[�0:!H{�����w^�j㋫]{F,3Ʋ[ǧ4�WdW��Og��X0���\":��[Xi�7Mdnvm����ED&޹� �5�]T��:���xz�A��k�^[1����kO��Cwŭ6KJ$�;:�`x�<�b�Ψ}mW��}{i�U�e��e9����4�
��ﰮx��z��w7�]�{\�eG��
�h�"J� �	ܜ{d+�t���]z=��|K 0wy� xT���ر����7�y�<<Ӗ������
�"�(Q�oG>�����1]�d���W���!Y��A��Ã�
�d��5ko��-��s���Cp�a�a�~9^\0U��i�L��7�zn'$�4|�P�Vd�xKk�V
��<RT�xy=�>9�鳰T[���)� ����Y�[p���M:���ƙ��<$$�3���\�o��!"��v� ƌ�xR�/�M���E��M��-]�Mі��Õ!�$WFSy]k! y��m���f܏=���X`�S4�ゖ��5��]�qC>��r7���?{Ӻˣf�z��LU�T�Wq��@`�]ܬA�R��j��dד��b5�Ͱ/^d0�7�Ɲ��Z{�)��>Ѯ�{�ں+݉v��t�Lk}݇7g4-T����Sa�3�|7�ˤ��T����:��Ґ���p)�|���Xᕹt���#t��YCÙ�f矏��ZN���S�+�ƀ�dx��P5��٨�,ttVКԾM�u�N�t�;��0A�T�o�2t0B��W�d *z���G̥n����wO�v�+���߅z
�4��p�՟_�ѪQ=��(�f���z�
�k�]�
_o���T�ۂGx+�WPa{��{����������ԭ˟�=>Q{�f�OT5��AOR#c��u�/>[$�����̩ \!��^�T��
Y��֮ �}��:�ɲ{�Vz��HP�V(>��j��t�-K�u1�����f�<wW��l���Z��]s0�@�����W��>W��"�=�lAU.�A�*�Cc�m M#�VR4�豲�{T�r�]��U;�P���U��D]���rU݁�0��,��`�zt<B���pkH�p:�c�z܎%����̓����;4<�\�Lc�-R�#���6�[��!�C���<��}r�$#��u���D9j�:cgb���{.��	��\��S0��ÖR�5�9e�,%��x��CQm�9H����]_�B4�	��Q�q�$�8��D/����,�c�4X�^�c@ �1�pÀ\Է��.{NÉ���\M���Mm�<3�W%�K����׏��!<�nx��{.
���K(י��s�^&��q�1��8��E�I���]�YH���������=u
B��)<������{@�+�*g��J��*���E���T�"2�Y���s���j{�&6zn�ķs;���"�c#CӕK��;���d���K91� �|��T�G�q�b{nU#N�eF|�)�<O�)}�����؉aYV�{8V5���0]̔�0g׌�wV�U�-Թ�uv��Kwcr0��A�]���s6Mm�tRp����*��j�I�w���l�z�}wH2yP4��,\?�U�ʶ��x��3�ح�2w����#�^���׮s#>�
4�G4���y�I����5��:a"��>�x�1�������D
s��0�^�A��>@q�lL�lB~���YG�uީ��z�/��Y���M*�C��)P"�Z4׮��]+}~�>��`��*�ʿ&�ǃ�&��W3��*�\�e�����=���4�}
��%
���n��~Vug�@g�fն}����s�����fˡT�4�~3MQXo�z�L{���Ct��i���˯L�82v��;f��:�qm���;�Y�y%�Ky�j��N��p��c��o)����L�G��P����s��M��1v
���p�WfZ�
�|���_Qˈ���8|�S�3� �S��h���ԋ/��=�l�o�&NԊ�0�R��u�W��V����׆��d	��\�|J�k�w3�g����@^���Y�<E�n�e��u��o��H�u"*!�|���E4�f]���I����b�*\�i�}T�n��)���_��	�$E�R.EN�:l��r�����4X��ѫ�E't��=g����9 \�=I�ؚ�q|7%ge�u��&@�5�P_$;p���Rq<.��������5}\������0��U�i�@�f�s�]i�lS(��r0�<�O:��Q��;eԫø�̸�J�"���)��K�����00��K�w*f�r0�>/�.�Pv��o��7�wH̙�t8�>��4�*A�ɍ�;]a���v��t`˨Z0t�Z�B�qp)8������23=]���qK��[]��y&�I]�]0���*m�έ�֥7³�"�)n˖Q���W�h-U�)-�]��p�q��ښ�'9ee��x�ޣNI�wn�-�{���Sp߷j+*�_F��@��6^�|�D7�˟�6U�"u�WZoç`�i�si�z��
܆C,V�'D�HmI��L����q2�,�,�\jz$�t�r%�-��-��[ �Q��f�xh-�.^���8��f�۞�J>S�<���S�O�\�v�hO׺��Ӝ�X�]��$T�7V���͞o��1���2q��K�@WO:�gL�Fzc�{ U��<b\��i�#�^ed�p^�N[��Se���1��PՎ. �=��Uҗ�iw� i<R;K���<�*�b��Rmh�=�îd%G=��#��=*�3kFU^ �B�<wt�������g/����+��p�wKm�%+Wi��e��d�Ѱ:Ƚ�y�f��]��]������D�9�b��hc����:���s��8�V�$F��*w�O_Q�q�B7�[Q,u�FagyS�
�J�}�y�o��ȑ�v7[w�ŭ��pz4� �[����j�����[7T-��U��z�Gn���z�c,�������|Vݯ����z�ΖWKjt�{��ɣ�4g�����);�L��*��f���kpOΉ�^���V��g�J��x	g�ֳ��O�;�c*���E���Jw�冯�a��F�Yp`�S�d���Ƭ�:q`r�V�Q}�o2 ����N(r�N�&>0t����J�ɷ|�p,y{�m�1,�&�|�u\e)d��a|%ՓD�&��3�<��.��3���2DV��6w�$��7��G[k���͐$}���j��-T��v�x�wP
��0ԭn��j��Q&��y�Mڊ���cfVw�����SVa��74�uj�qC;u��㺿\I�C���<zz�'�|�{�0t�S��ԏ4��P�u$���n�N��Yt�$A*�=ҩo���[!�Y�K}qmֵo�wu�u�о7J����֚]���t�f���2�ᙣI��Bn��9K�Y�y�3A]��0��X9��C*�8�`�S�Ǵk')��"ip�V�R�o��p��w�s�oE����M��u��
�}�f�5���ò-���*�w'� �]��V2n����F�xx��Q��x�+^��ߥ?�4Cb�N��W~��~;ݐ~�j�-�ΰ���җ�uw�8ʼ�ݐ�r�LK�|F`ٗK���=]DYy���w^/l�еQ{K�X6*ܤ퓮�ٕ��re��]�7\����vt���%8U[Gݪ��Y{�Q��m^T��%m���^eɆJ��JSܷ��ǻ�҈ZǢY�VkeDrr\�\�1;A�u�;SzLT�ᔆt��GYb��f�6��+"W++:Vy:|����VS)+�f�]�@k�䘢�Ow��X���U�Y�G�h�DB+�BMïn.�v�,=j��9���-T�֖�s��c�[t�0��
��\b�qmk=�[2&3uԚk�&f�m��:ˎh��ȍ�I
M�[����Ck�]R;'r�����*V)$ff�V7�u�x_{o�{����7�N�UTA�b�(��A�SE��L�A`�(Zʪ��W-b��ZX��`���WMAj�%U�Q�)R�����X,U�eQ��D�iF.�UUR*��X��iխ�D`�"���PQ`�(9J�D`�E���U��2�Pb��"*,Q����H�� �����)Յ$`����Z"1Ac*��TUb��E1)P�",cQEX��",cAPEP� |(�����H�N�RB�֮c"i�K��\�d�C���`&�+�iK�c�t�)��}&�Ŋ�>΋�3\8ƌ� ��m=�w�u�|o)&Η���
4�>��Nv����s�Dp�L`������E�H�CV�X�{��"�c)��'��j'E�,����=U����{m*���Hzbc�KN8��b[ �"28u�O�tk%���� �ھy��(�[ \��%YSz1�̥.���X*���=��@� �Hҗ8VL[Z�����.{'���W��ЂA�v�:�@N���Fߎ�*<�� �f�N�~	���'��8�hY1��[��Y՝؏'�1��������ː��mӧk[[�	nQ�&8:�����YfWV���:�ԛ��ɵڲ��6�=�ݳ�왒s^Uv��xD5"�>�^i|�:,U������,���R����w�2�N30���94�-��,��p�1m-~����,Č��c��`^'��c7�Y~�Q�,���ǵ���}L�m܈���[Ҫ3��U{RX�x��h�N4
W��yw<��(�Bʥ�=d,<�/�'�t)��u@�G.C4#k#f6��:�	���߱{$ߵ�.yPy��1Y��$��q��1�/�}�����^��|�
6t�`W�Ń��=O��F
����ö2��1n���Ok�eu�U��(��4��j�|ժڊQ��=������������V�\Ǝ(YX�w���*�9�ԯx��T�]��F��g���W\v�+]L��\nGv%�Ic�ࡺ�>�|&1����}'9y\1��Z'A������ۍ+^�Lt5Ғ�6�I�]:(@S��]��D[��z\\�n{5�^\]B���/�r�t,�xw8M���s4�$����CP�<�+�������{�%.���C=w���H���Ί�~h�ܥ\L��������5��r���ET]�j�C�*���oAk4��K��Ó1��+"�	�����׹Â{��,�B���]K��o�'x�E���i����yl�ܷ)�7�t�8�ÛtiF$��<�=��IWT�l��gs�uD��~*��Y��~z�,x�Q�q�)���q���V�/���]�!�K}+����=������N�n>��u7�q	-�ߴ���Ϡ��05�����O���یu�Y�^��C�����=��t�'�*'�H��E�:{ �z�7�4:�rj����(�}p�{��x�Z�����s*���;�SP4��ץ��V*��/	����{Ԃ��s �9��9=ys���cBM�t���&������.�_x2y9�8���'>����F�u}�S����
���Qce:��d*P���:�3⫘YX�ػگ�����M����9GC2zVmI~�0�R>H�Y��-K�Z�h܀�.v���՘c�"R����R��o(u��\���aGa�\N:[��i��Q9�'g���f��0�4�;�qh����e�6.��Ĭ�sr]�\���7��W�g2"���켲έ�ȣ��Zi��{���Au��G^�_Q�}t��l+�D+��"��L�X�[@#L����+�b�^�%n�8�&�Y	n�&/#���u�ز�'�=�V�[�/����>,����S�ZO-M��q=\ҫ��cCZ��"qf�X�.�?P`�[���&ޯy?'�ٙE�^Sxe5ܯ��䋙b*'�2��}Q<���c.߰����\�z'�&6��ԗUʈ�6�F�ڣ�����t�
ٰsx-���߸����+ozY�vh�F����L���{��%CcV`G]n��X�g�\Ewvdu��P��u�.��J�Ӎ���;�A$�ջ4e�2�.�jx�)�t��5��5��H��=��[t|_��G�zN�렬[��&\^�<�I��=��0%K޾�E��]M���k�D�ԣzL.rr{GE�{t�Ђa�(�VZl������u�����vה���G��)m �`�Ġ�uP9J��ߤ]�������A���z�wr>�\yyUG)l�r ����VN{r�r�1�hOvdѴ�*���>�:���@��&/r��/�:⪆���w$����$�&�)s<�J�ZO`���1<��ԓ��-e����ܧ�\�U�i����T�`{�K�fXY��'ۤ��d���@1�`c�RZ�\=��}����Q�08��œ�c�%��7�A��SK%�4v݈�fu���a�`B��v�^�&�R���G�j�d�Y��΋2߫}�*4&>|M���N ���kw:�Zڷ�1хk֒o�bc��U<go_�,q�dF��������(	�'vn�M�7=;_���L0�1�z�]:f��v�}�l9:��� ,��[����kܻ��{�ֆ"X*��-x.�麮�ҵ�WC[����e�wg����qy�_0�A���tr/�9���KGf��,�Zj%m$ �ˑ�%¬"W,։���=M��qff�pK�PҦ|J�/�Y���{)s�~��\�;n�Q����_�L�
Lk�[���N��`);����|-m.�2-�\��Td�5�@�ǚV���1����3q:L
LV__W
�Ĳ�Y���^*��b�Z�]g!u&�r�Qf�S��&4���z���Nc[��^.o2wgQ�WM�<�\@J�m�������,M�Y+.֫���oJ�V��҃Hi�n�[\�Iی��.��(�N�p��K=����`�|5֛۠�С�n�,}�Ks.����'~��5�6/�3��FD��Х�C
e����h�)��OC���Y�ڔ�'{�khS��I�n,��Hǡ�a*�W9(�Gx�l��LB�2t�ȕ��{�^�]�T�s�zB[E���=�S�=i�H����K\K�2jJt�� ����Q�z��rv����U�S���b�Ya�m����qo\�q���#�*7�c(�,��e�Qã2�c��`��tW#��kZ������* �����8m�r9�I7!�y�'�q�)�e'i�]�%�7M]��s-��&rvr�hؔO�@1��`��QL�f������f�L�֖�jg�od�0w�zss��ߨ�^�<���r�kzUҾ�"-t�K������G'v%���,���йԱ����v�iQ3�/.$�v��p��S����l��=�N+�a�ŵ�(��ga̮�������X�O��\0��BT��ٽ�W)=�޸����"
��֒O�I����@���.A%1�iʨ]:���ͳ���KD]���,eް�q�\�	�ٙ�$�=��r�1e��w�X�!�n\w�����f�	%\aE���ݙ��m:T��	I�����5�̻����pP�v�q:�������.��\���b�;��@�Ģ�:޲�ff8�Q��"���\�yDu������[I�;�U���vLjRpH˓�y�)b����{,-��hVn+l)e�OQL��lMec�p��'�>䴁*�2:�%���S3�oO
�9�.�G+�Q��y�5��,���T��r�E)}�Q�fú3V�ri�Z��Nw�ecTw+�rx�T ���H�=���D���S�Q
�Ô�
L
��t��2`K�ڀG3q�hЎ �&�#�]c���~C��߭�[S�R�UU��I�L�? D��e�Q̓�Q{�~S=Գ0���S:w�h�]�=j)�L� *�%a$0��P@�u�uC�r-B���!����w�%"4�!2���O�_]��i��y?Y��ko�8,5�����<Z�8������z�8[�d���|GW��-8�}�^H��'� rETA?$�F!%hs3�"���!���}#F�U/��p��<3}q�TA1��?J?�(b s����l�X�2[�lԍ�1����5�3����>���`�t�J6mЁ�]��� ��c(
�I�Sƍ��E�D:�R�
1h��r��Bm��4�e[�yT�P|�j;@ULۥ�I�ߢmz����{�j5I�C�Q�����An�|�k'���H�m|BATA9��$f;���A��5�b��v�q[���ә�����rC��y�=�/a~�^�[�����l�a�{��C��3���Ƅy���B��Q���Q�^��7Ž���,��r}d�P�r1,)�����P�sm""cPѡ~F#�0 AA!����Wy��,5���"֘�%��.!`�h������)�R��BC�TEQȠz:���+�:�UJ�����lzl^�O���~{��do�7�;9�s���8�6���|ޙǊx�w�R�����.��p;
��#�)�杠*�'��-Ɍ
��>�[3=�)��5�L÷�B�6(@z�U(AD�o�����t����eo�w���q�+��:ڀ� �p쫏����xԺcf��'j�RA��N�ł��x��5�����}�Gʞ���tx�Z���*�	�wSYp�wxp��kvW�R^s[&��B�*�L�?���)��`*�