BZh91AY&SY���1_�@q���"� ����bD��     7�}             >�   4   4�     QJ@5� ����z�¥EU��v���ت����I �[5Zȥ*;gmEV���`Kmcm�RX�U�I&���l,�5�6���J"�����Oi��
�F�SE�3U�I�mK6�3f�j��iX�Vle�j�Z��RV�����l#Z�a���(�
T��M�6�͚�w����`�Z0z<   ^{GԂ�sD*��Wmu@k:�Wu
�T�tР����:5ݨ:��h�*�Ke�gm��X�`k,Ĳ�m� �   ��( �s���l4��T(f�Р���2�J7#�ҚV�vu�����J 
�U�����(�h �]���*�-f�E� �[�  �;�JR���` �M��x� U��q�� ����:
�ooz P����ޔ���{��M�ory��(R��W��@	 v���5Q�m�m�[kkx  �<҄�C��9�
H��yy��M ��<�2u@#x�� �)\�j��ޯxzWM(�[� �	��E Uw]��h���B���[%l��hm��   �}| �s�ݐ)l��

��s�)N��� u@;v\tc%-Ҹ��)WO6u
��+A�hY h}���5��Z�� �6��1c�  �w� R���҇A�:��*���-��T�I�� � ���֍�nX���+�  �n��JYu��{g)z̖I�j�M���e� ���
,� � р�1˹@ *��P��ٺ�%����4��Wl �n 
m0 +�n�E��F�-hU�fm��x �  7�� �M�S����@X S�  ��\ n�����B��Ҁ��Y�m�)Zmb�Ԗ�[+<  s�� r�� �V ѝ����u���4`�����@�us����@gDY�6jUS[fD�  ��� :����Yv�B��j�:�� , �s�@ni�F�;�     �   50T�H10d��0�i���)IJ���  M10 OɄ��T�L 	�` i����$�T      7��U�cRb  ��%$P��2�@�@z���G���oqں9�j�޳�N�6�)���Տ{����������������* *��AVS�  *����G�?���������3�����
�?������ U�~��J��" "�����>���~l�����'L	���W��l)����e���;`O��� ��=�l�� �ʝ�l��>��U�x�=��l���;`��ȝ����{d�G���=��l�N�G�A�{a�G�Q�}��l���/l#���=�/l� ���`{`�� ��=��l��*v���;dN�S�D�<�'l� �����2���l��*vȝ��l)�;dN�C�C�'l	�
v��l��"vȞ���̇l��(v�'l�� v��'��;a�0��'l	�(v����l)�"{`N�S� ̽��l�哶D�;e��*v�� �{eN��T�{d��E;`�>0�"�;d^��E�:a;a� ;`C�;dG�v��C�)�"v� fG0(=��=�*��*����TN����N�T� ^�UN�O�(�l(l��C�� S�U�Q�S�QS��DS�")���"� 'T{e {e{aP{eP{e {e@{aU}�>�l�yaT|��>XD����D�T� �U<�"�ʀ�Ƞ��
�ȡ�;aN���;`<2=��l��
v�����D�;`N�C��;e�S��;`N�C�v�=�g�@�;e���;a��v���n�C�@�;e�@>o{��`?���ӜG������u�D�~+��61M}���c즫�	,R�λk}3u�63�g��� @{V���ܗ(!)t�޹��Ε ������j�-7��:�����9���|;��N�B\�J\��^ g(��o�"*d��Z;�v��8�Q:�����a]6�����2ՠf��wL���EQ���!{t�b�y�o!U4�r�`�nY���x�T1v��]�9�n��
<"=m�Y*}���M��dH�Iڴf蹥k�m�;tD�kt��9��8�"
Ff����8�l'`�<��uq�	��]��$Y/��n�׾L��2Y1���L��W9�B� ������_d�@��0�	�k���v	�WY�'q�d�o7��-j�!,ί#
�Ӡ;�Ql����]k���(����F�.rs��']�1�����_h9{:�QDW FNCzqmS��v����{����Qn�3�����t�׼-�8u�m�b
F��X�k�m�fc�����䨗Ftx���<�Te���-��Ӛ�@}�$:T~��l�(B�n",���@2�1�:��֜�0�x��_f�c[wz����e�&��b" A��z�U��WB�aB�in!M��cp�k�W��˹��Ze�+�Y��@U�[è,] �PZ��{HQ�}ʘ�o<�pr�t�t[�:'v� ���7k�8�m{q��l�\���e�Qǈ}�"=3��ڹ��@	�w���쇉�"E���N�������|��qnp0-x՜�v���j�7{.MD�иM3l<ub<�0��ڎ2���iw�0t��Y~\� ��z�Kⷡ�_1p�o��NBܻ�RqMj����u��x��ӳ�[qb�l����t��1�#���ͺ�6��l94nV+���9vn��}FB�5r�' ���y����ɚ��ೡN3�Lc�;XE�6i{:���ܨaܛw��ɗ�8���N�1�yr�{5i�m$�إ=��]�X��Z�����λ������j�;�Ꮷf�[�Or�������SK�,����~g*���Ϩ=���䷒ۥ�lƻ�f�CAΫ��cwr����otÝn\l���b�fY�U�q#��	ɸ󱄎��;1�'T�����4=^۶��(�>}�7\�#^.H��Nw!�:�'�B�c���=kwE�[;�	�'%#<O�R�{)�K�98�ܲ��<�u��&�y>o;k3�B�>�p�'�� f��qig S�X�q]lwa�*8��d���#f���.ꎍ�Le�;FC݄�=��y�3t���Սُ����97����x�n�\��gt��:�C����8��b���v�/qth�l���L�TW����rn.��ݣ�I��ǖ,E|~G;��''�77Bۭ 2-��{�>6Q�\'wh'Tȭ��{)9�P��ι*����7��n��5\o�<$�\+�_�mUK&��=�1E�<u�tJ�|�:gi6e=5��L�[��n��!��g-ҹ}e�~.�������n,���]���IwR�����0!1���+l������i��B�-l�n�ۦ"Eǲ��H^Q�uicy�g=�>'��&vedj�L���o;��d&��҇��:1`%�.W����	[��X���9�Z�܇�̧��y�4���=%M�p��wH8w������������۝�������$�9C1*$�@��pֳ�S+4^քvn��r�	 @Jƭ�0^i��3��X��Y��;�X-����	��{���{�.�	ٚg+c'#p�a:9��&�Xs�H�L����wc�2�I�¸����z��uq�e���4��v�.\����\��ʘVOmj-���s�.WO�/q���B�h����ɚz�:��Fպ>]���{e.�+����δ�׽���AÛ��ye��.���x��c�uSN#�4nRY��O%��.Y�n�ͯ��A��g&��L��$�*�Qt70�K�ɐ&��Μ�Dp6����(�E�ޠc9���ö�bl\̤������M��m=ۯ�6�y3�d�J`&�{�
e7��4��W���Q�/b�%RA�vE��=�̞��[���못�+�{�n�T���N���u�C9>iq�cT.W��mv,�,�h8:]˒]�M"����5t\��+iŀ�t˛-vUz
E1t>G���q�n�wFޣ��������U�@r�������r���٣Y�U�\K�-k�ՙe���O�K� ܝ�7�P�[!�����@qTUg�Λ6����9�^�U��{�Lu�Ý�q�ӸaM�%ζTGU����r�:�}�e�N3�OTOz���(0y�����LzW]���������Z�- ��o-ワ\��AW'-QsZ�4�c;�d�,Y{93m���͏Cخ��æ6:���n֨0k�`�mǻ�^��Ft,[�'�i���U�~�Ƌ�)��gA8nL:9G�Cݚ�=��^�l/���ys�RGة�a����.��~��ō"��\�b�!���ŴyGhZ<�iŵt����wbP;�f5�gb�j�2��%)��Z�u�o�;�/�V�`X2��g9�m�}��g7��!un]�uNQ��ړ�e�z��6N�W��=���n��ыX�Cr%	v��V�K��sX�-ж.�&wa���:�ڶ�k�v����=�wPT-�����w�ۗYd����˚C�l��v�E�V�l���Hl���� ���٧'�j'��^�����1�Au�Ɣp� E7j#���y�gN-����m�\mH։:.澯 ��NS���:_C���uT�-�,)�X{6-���zq�I�+�{[�o:8jāZ�I�uld��[��O��\�-hn���.׃&��3�e��1�m�I�Rfk*_�:�7�AH�ʱ��,�yb<I�����v�V7r&U��sS��'�a�9�P9�9��WS�P�9�ٯs��v<�ZyKߝ&eíU;�dJ��Zꙺv,x�%����A��CB�&�^NĎn�W5�߶��Iߗm��C�1��r��t�p�%��7�ݫ��%aN�;f����x�Cp��n��w���p�Z�
v��=N�-U���4k��w�|��}X�>}�yeҚ;�����u;S�*�y�Ë�by1sY0K��ć��^��n��G����P-�J`�7F���"CΈ+�zO���ux���t׀ݢ��M�%#��ͭ�vJ�a��ӽ͙�;���\n�����yu��������7'wn*��ݕp��3>[z�8|�8)�\�eѯ�w�5�.cSn�]�5my0	4(����x֝�i�r}S �Efwk����8����5;Zp�B7Fp�wf'�A=��؛��N�qԶZB=6� %�w.i�<J�ѓ���%��cÀ#[N��*@�m�!����;,�\�s'���)���j쵱ٴ��~�KS����3���9t�bOwn��ѻ#}����eٜ����]�f�����E�6�-��rq����Ný.��m�I�t�FqrY�nH�����$����:ta��7
 �΃Nehmy�@`�K���#�kmax&kI��|�$��>�&u�)�1맮���:�jv> L�e�l�.]-�R���cH��=6��m�w���G:
<�o^m�\彃��e�ёt\��Ԁ�I <�5�YA[��b��[���3h{��q����́�v+�Q��Swb a�Z���n�Gj'TӚ6Z�ja�c��gZ�+Om���!p�;P�E�.m�\�������9}*�{����Tto��d�����'���P��q���v�'`�(��+�"�DF��B�}����+7+��Z�zSץ�ۉ�1��f<I��7�&Bn^络4��w_��o/_�dS�a��f๪��<�3/xu�;�Kg/i��7�X�m�&X{.�K�.n �C�k�6����baG�v��	��;6^]�dlbN���w�ro,����p�:����K�i�e	�pF�i)�����C��`��҇�����ʖ��Cq��+�Y��T�Zk��1`:��
w90i�JK���e�x5mc�I.�
�O1"R\��BZ�D浭��,��7�<��T7�>>4��3�^)	d�2��Wn>޵W��7����5�ź��|����O��]�_rX�܃��7��֍��q�L�6���bB-ָD�Fu�E*�.#��2<��ƍ�/.�h��3����F˨���>�K� �o(�N�n�T�ؖj����gd����a!�:U�hxyڛǜ�Dx��ހW��6u}�k붼���� w�E��<�ڱ��/�"d��HX�x��Y�Y�6u��:1b���w:rg�}ͅ��nlO5���aC�coL?L�{����������7z�u��Gd�"x%9��=|��Q`nG%v̢ٖ��R��o�K��3&)sn�O"T���"zi�k�m���	X&սǆ��`[f�Y�K:�ţ�	4�"�٨hI6Z�p�A�S6���]�BvZjt��O�/��w+3�y7������bC�f>��W���Qո�l=[�ŀ�����{����U�cڛ�:t��[��[�; ��q\i�K�A�+"����Dsj�sj�Apt���f�.�����wp�"�ΐ�S��W�M��-�lR�,���3��у5��n�K�j����[�a:�K�6�w,�C�ESw�lؑ��P�l�� ,|���c�8ZӤ���rS�9�;gor�ɢ�%5�nI\���eQ���wb<����:�f�8�M�ԭ�m#�(�6,#U�{��o7n��3������E��n��v��A��sw�|,�ӱ
�/�TȕCF	�ݓ��L�[�&�5WB|��C�LI=@�~Na�{Z��]"j}�7�o����h-�|lnh�˅n^Ì�t��䈫�K�;I�Vw xek�p뛫�}���MXX��i�v��4��d�K߯qy8��k��zw6�	��'�ky��8�!�lkO�I���!VmΑ��;(s��@�'k�0ku�1��X��r��fqO���{��0M9��E��g{�^������q�<3)�a.�]��ψ嬋��V�XN�P��1�,���n�A������dA��shhJ�Jt;z���ڒZ�,��X�z�η��8���'k9s���s;hx7�m�l��lmGAmM���rո�8m���q��G�ck[OblH��N�q���a��r��BK��������\�"X�4"B�hѥ���&9®��!9�R�˵'�mR����p���xdl�� D[�����ܩk:�kw�m����.�:���ͤ�c@sqT��^�dA>�C}rΎ����
	T(��hހX����rSǃL�Z�WY�jF{Aie���˝�9�8yLsuք\nv�ݕ��,�+Ǥ���܉������'�6�EL�c�g8®�9��K�ww�W��2��e���D�m��(�:��2��0��}�$�[;b�c$��;�����.�Q�Fܩ9��!��4Y&sc���s�J7;}3R;Ć��n�O6��g�ғ�N>��7paC��K����Qiu�&��l��8��v�+�j��7����&Xxs�����.o��Q{c�NL/�+͡7DRn�אl��[he�)�rh����
�#j�⚠���qQp݂�:������5��b�"��Φt��k���.��N���7_�X͌��X��Ϟ��'C�������Sr��N�}�G����D�Cj`eӦ�����{���"����rM�H�a�Z�fn%[q���ܓ�۹>��0�SR4`�/�i�!��q8v�;�qKNEm�����B���B�ܖ�+2Z!�E��/6�im2q��x�K5���p�1O�ɜ��Iݚ�6���T-�3p������[Aѳ&1�̰c��բ�f�s����v���;nm�7|6��C.C��"sQ0��VW7���=
���V=)�z�\�x������v�+���Y�t
>�z:h'uW���l͕���f�zȅ�uПAT6�p���aؤq%�;��������E6b!a�/z/3z�5vL���/p|&�u�i�,՚����^l��4��p�<�TA��b�{U^��Ʉ�CsV�n� X�`����Ck"ӍI�.�L�)�l'Nm�d1�q�ұ����Η�P��3�#L'LOy�<k�H3�DݪN�Oj�d�m@�3QH��v+��n±���R�NI����/bM� �_x<�0к�e�a;ƌ?���xĻ�g�q>r�x�z02�g��r�%'EI��4�
�QX]f�`��+���9-������9�,�\�a.�rF�����20v��2�I������i��$��^ �g��Z$f�V�%y��I��=�ϸn�b�`h�O��"����&t��(�w� �4����'�S�6�@�6^�eQ��%A���Lg0PM�0���(Ҳ��6Hg���#�7�rW$3Oq�Y'N������F�}Ua���o=!��>���V=ѪhI�Z��l�/��z 1m&��@����צ�b�U���&�C8��lx&��^ ��,vr�jH�pT�E.2j�j���8�?Ͽ��{���~z!{�	������k�xѿ�o��8�\4���-���n#7��w;l�|�]t�sTR��Z;�)�E���TSkU:�D��e9��x�C:Ql����&�s4��Fh����6QC&R��=ׅ��+#՜�~{��^}�N�1O	�y��w�$�4z-SfӶ��{�N��!�=i8~5�sq�_=���&1��f��z�Լ�tO����>�&N�De�W��)��:��Sհ;̿�Gk��[JõF�h���珫	>���ܾ���վ�����֩pɏө@ge�󦩔/)�Շ�����Z�<�R�>ŃÞ�O�����ː��?_q���s��ن���� ���&��z�.Ώ��E�%x�O��R��mk��P��7�v�;�I�mM�F;���=@J�+��x/k�c�����mA�\r´{�f��X���œ^>I<��'��V<��j��Y�'V۳��l������w��O�dD�UC}Y��s�Y�KǦ�����sn��g&6�ߨp��۝�L;Q^a>����W,�o��ѷG��}5�K�×�Gj�+�uA&A�GB*ݤ3W'�ۮ��͖���˪�L+�SӾ�=��:|���3C�𾕮��Pf��V�<��ѳC�f)A*��*�J���-��|V�FxEu"^��xDs�s�H�1i�fX���(˃4mi��z`�,5�
��x��j�\���q�qV���+z�
7��N(�N�{�+�=|��H���j�h{
�}컮�4^Ц��N�^�wd�vv��ʆ��>K���+U�`�v�S��hr�ˍʴ]Wj�{��NL�<���5�V7�e��BJ����Ҕ��D�a���m�kӶ�O��Pi��mŢ��FlQ�뜍Q���������E�Ս��fp�b<��2d~�J�B#~���gˊ��2�D�}ñ�GH��Sa����X�R�wV�n��śyy�e"��R���7jH/�a�4�oRK����G ��s}����{�RD��}k����������U�l�|ٴ\�X��1H{�7M�Tچ��b-��J_M���2��FD�F�ڽ�^������G7f�&bq��=�c3�J�J��:���'��5 P���Pǹ-R煝�c���<Γv��Z�NI�\���)��"6w17B��pf��ߺ��`y/i�M���%���.��Sz��d����M�N�.����a�ٸ��l�ڔ��9Y]���=��u�y�tR��RP��������l�X���ǡ���lD�M��y9�]�����x����7��M��Lpv������ዴb�h�	$~�����B��n�b���w�3U��]�����%��v��^����A*�nt���kF�lU��}S�+�i�γ���>'���lk��n����D�E��N��ϝihm`�7iL��m9�
����4{�a�c�4էq?*�]!�q�`�����ܣ��:{B�i,�tv�|��:���{�3��r�|����|�{F�{�s�ruNwO��y��zIԂ���|NtR��/Z,���T]��v�q��R��W��rE�K�w�M>�۝�Ň~+F��'g{ޥ��&��'vwD3{.@26'V����j0�^�jc�m.E�|���O-����jù����]u���:l�Mg$�7X�����|Ď�ww'Q�����z,Q@G"�5;�7Ԇ�5d��d��,�yAǸ��l,^Z1�P����].�y���W+�[�)E�rՃ��<R�|o�~�q��:/=�fp�}��֟�ޕ������Ա �a�ZB�O,����S�����F��0��3�\�R�^l]��7^��cj2�UX}Ǣ�*���$������ҋ�-,�����o�vC��[N�m��W��`~,��|��
�6��=t�Y�@f����?J��|���I���G�A�	�F,�v���Y���(�w������Z{eS�f�wb���q�����}��եcA�N�����[h�(�z<=�m)��)ts�H~?l^�vc/*��}�{=��?�ЏF�M�,�i2M����u8��Ϗu�Ȧ$r�E��Tg#q̘�g�q3��{m�z<V�M��ɝ��lj޶�]�ۻ��
cO�y]Vs���X=�T{f^1�D�����5�G����d�.l{���]˪���*�K�]s�]+&B'��ntG+H���Xǫ�����E�$�<93эz�v��Ku������ê���]M;-)>H<�D�fw�0�}��^�'��1f���=��ޟ	�ݲI�cN.�n�MЇ�e:bT-��T�g�Z�1�7�qntP��i�����mv����葮�_M��!��w�0F^1��X���_=��ݖN<I\�����9��8nN�v�����s/�.�="u蛵��z���Oqg�����q[�CvV-<:.o����B؆���j��9kE(x��n�Cv��~����R%�x���a��xFr¹��@���'7�rz�8q0����n��0�i@�9;
S�⇼���O9���;��s��{��L���.���Cٜ��l����}������b�Rbȓ�bZk{AU�J��j<q/�n�l^߹��gR[�,[�b�I>ݨ��-i��5)�DK���d���4�pE�%��ɻ�lgvG&��j�I]�.��k�Í�2��|�KN۬�u�}=�5�r�k�Z��׫��xz�^2�\�e����8�d��W�y�N�'�����-2#}jZY
�ӯGk���2����k�����2k!M���+P�A��B���2fֆ������v�.?��2������qz�Q#hk�̓�;�r8v�z�,�>c��_Nc�.�O�^�}��E�;�h��U�Y�$Q�$TM6��:�/QsK=q��WK�Q7ղ�^�F�<�z��wCӍ�qĨ��חd��RQ�N��G�I��G������c8I�����5P�;��v�ESj7BN��{ӂ����nG�`�w��K�7M��ޒ��YOJpn'N�L����sb���)C��ھ�zK�3�͘薠Y�z���Gx���}đ!�f���.o���W�dn��=�'�Q�3� VGUQk�Bm�ᚉ�.�3�w:gN͐��h�n=d�������(JFe��ԸL4gC[�4��2�����1�a�h^)�ݛx�m���9���>-9����U�a<иq<��-ɷm�bvy���g�b+�P��.��7�Z[wkT�]Wm�P�Ks��@I���%����v�Tn�|�����;���^[�ᢩ�E�R	/.�؊��^��W��G(�j�����Rsf�;.��8�sNыtF�`�N�G�y݉Ш+��|���`�h0��t#��*��G����Ի�g���e�X|���f_i��Ի�v�ꐒ�D�;�u'
ӗD�ש�7�;�ү�)ojuY�7�����ХMW/�N:��-Yŏ1�-��������fΞ�q]��R#�x����M�:���.M�qаz�����Ń:k�'���|}�f����}#T�� �/\?g���9#���ǚ��]q�CǮ1yv�د@��K��/8pZ��CD�<�G3ti�&J��w3::�3n5U�c��,�pK}m��N{{K?
��෻h���<gQ3Ȏ��OE��1���V�c.=�u_i+�]�.��ڗ�I�R̂��iV^����� j����"]T��VP�}��#9}�ξT\i�����p��^�7�����K��hQ˚5O:V$Ż��B����i**��I����7��HzĽo�g���Y&r-l~�v�����ҝ�l"�=p#
>��¬a<3��z���r��\7@�6y [d�`�m�s�S"�~��$�[+��^�͌Z�üs��ٳ��#l���E�[A�S�q�\7��k�!�v��%�a_Cp��]�Dj��۬o���o�t���WK�^vjB,A�]@��{-@���][���]\�>���Sީ���b�EY��5���s���*I�G���'WoY���Oh�N�'p�͞+��\XW�N�׆�+��÷��D�
�t5g��Mn�{�k��Dc�x0(���X�R��>�F޲��ے��{��Ox�=�/7��9��>��m���۽��N.�l�8��O)����n�fFC��g��)| ھ7��,u���~�����g��V��ܓˢ<T�pfU���ӵ�v^�x�4�eP�m���h(8&��FɮC=�mi�4j�T�W��C��^cvM��9zyUκ
�V'a�u�v?��JCQ���V XP{K�X�ϐ��S���*�쉪���S]����4�����6����rF�ޘV�Ķ���x+׼�f���j��5������,��c�L�s(M�Q	m�T�}�J{P�[����@^���G\��w��w�����l�'��Lcy��J6��s�z�u{:#;1e4�3�j����7<|���Xx����Ή D�,��������A�u��S�-�ĸ)����8���@o�otoϗ��M��ɾ*���w־��ђ~�f�-����?1oi����,V���d�7bY�"�5�P.h�n���<v�-�XgmgnN�x'�a�h��z!�;�<��Ίx�;z��;磧vI��@{F)�3�؉�0U�b1W;ꓑ9V��˫���Rx孭i�yvD9�o��d��	.�����0����i���u�}�:��=5Uf�.An%MY;ֺ���e`�J�X�Ѥ��#�{.9$�<H���%+�kK&�&3R^�[�m��z~3�wD�!�Gf�N�Tw��S��m�+2=�p]�L�&70��ʹ̈́欔HF�r�t���6%Vc7:��]�U�i�6���WwΓ�����ң,캺1[����9�*/��-�,횷FdZg� .��֞������sD{m0��}�,�?S�T
���/�3}���Y�-��e�oTGE֛��ӹ,�f�r�[]��"�j�iq���G�����%ݜ%:$�EdZ�J2�v2�c�eC��_��%q���v�G��D���{�^r��#�j����y�}9�]��xT�Iѽ��է�Q����Cc��J�/��y���R>��xkQ(򡋹��{v��$Z[�ܝә�������]�3S�>���>��G����@4i�:��./����0��ٽ�:ꁺz�ȗ8"�J�������[��k��r��}W�xx�W�OS�R�<�`�mU�+��PY�Kwy|��z�B�����w0�ͩל۩�D3K]jK��	���N;'���])t\�]@^���1EK�A����n��1M�Վy��kj!�A�U�}�<w�޾��ԅ�ʂ�2�v��zȩգ:I����b�Jm����/f�gc ̷թ�z��)�:��ipz��ԝn?'�{*l3���|�K�夈�*�Zi%��ّ1�G3m��wXn�7�j_l�~�geCX.�[�*��N�mˇ7dBF�y6����©61�Ot��v�{N��NU��L���6N5S�j��.6����c:�P`;�k�U��gkQS�|ky�2�0�Ϩ�q�,�ʇ��ݖ1�-�%5�wP�J	j�n�c6v	Ԯ;��f�tB�T�6K��[���?`�M� 3��s3��nn<��r�=و��͋�J����S����K���ˇ;���ZdU�q�2L����N^�h�6�3��*�7��R��a6��XE�1�KP�jk�ʴj�C^ݶ[Α�ڃ�[�:��ڼP��}8�޶���W��-����u�n��;+iȮ��ߺF��F\J���!�����z�:w4}>{���L�y&��[�Z���^���򢖑Ӏd�b�c�����;��n�����o[oo�%e$Mv�}���f<j�͎��G'��=T���9]��d�.x-�4:��h�D����D��������ԫ\�;�I��>�;T+�,�z/.��LY�N�=]ۙع���R�ڹ��^ʊ7��t�P��{�m{9i��{L���C.��}��Lm�|�w:�eq���b��}��:фA���Z�V��͡�.�0ʊ����xc���w�f��J�v� ԍ��Q�Vȑ֬\��s�\u$�k.���! 7�AB�>�=�
=�^�Cw��;@ju�6�������mn��a��ޔhjOxo�ىڶ3(S��J�
5gu��L��8�5QKΪ<�웛B�f4��%�Z�0p[)��=���O�n�ӈ�+��萷M7}��{��K�s����^>v���e�i�=��B׎�����mZ���W����e��`��0T� �4ܗ�\}Z��=吮>�=�����E�o��x��%J���E���r7���5i��:r@Γ��u��T%���sjS˼>���& L����ӝ��s�oA�U����U�f�W-���s]-��c�]�2uɻ�^n]E��Azc��p�^��L��\S$���2��˃-\�5&��')�OD�w]�g�mUtȣ��q�$ov)7.�y�MͅK�U����dwe���R���W�m|:��. *�� �	�׮>�>G��)�{��h�a|����J��d��P#ߌ��C��-�@�Ru�z�/�C��'�u�/�{���!�_1ߎz���=w�|�����z��"������� ����w��	���("����������{x:tc��$n��i��&�kD<��)��s�{��h]�!|e�΀��07��[;V'+��W �h+o���ڧ��.ڦ���'F/m�V�v���{�V��=&m��g��Y��3F.+�*{��.4����A�f�ʹ������:<ϯE�_6�7D�*m�{�t$��R�{��`81���EY'mi����Cd�T�}���k����6�]=����xH�b���mo���ף���@��7z*����1w"�Z�S�)�p$�f�E`��T���{W�E��DҘ�yk�sQf��@���]��h�{)�L��gH��M�|1��|IuS��6U�ӎ����w���|5�N���I�8b�n�97�N1��.Wbg�zh�꓅����g]}�M���.�V�,���4�ۜ�\��Ƹd����$Ns�R��y{2\������&;����g���i��)&�=5�.�]��o��
��{9�f��Ҳ��R�M�!�9=a1���s0�6��c�d�
L���ǡ�]�T!Fެ�����-~(I��nc}�_�*�8�X�*�c[g˹{wN�yq�mM�sW��t��p�S��qQq���ݒ;0��#ֶ�w�J��B��d٧���uJ}[��ڂc;�2��Os��B,������[���ЗԴ���r�%r�R��P��Jf��;�F��UMJ O�v{��Щ<2�tp���Svt���\�OX��q�fQ�a�qj����Ҫ���9d�h=�rz�:�!�wZ![�g!�Mѕ�L�e����nJ�T��c���0Kg1��U��ދ"�+;ۣx�}�!)ZZ��þ��Yn����{n��'�+e�r6Rמ�(��}�C�����;�u�a���4�\M@�]pfR��+�x:N]��Av�.�]9��m�C����~���M�(�	��21�?g��.Pʣkb�W�����V�T ��t�$n2tv�Ov�� �e���,���P-���^���={f��7r�b������ ��=X�u����!]����p�Z*ҳ��5sY������*���9�Y헽ְf�� O�17X��5�=����؂^�P�����w���ֻ2[좝X�rt�
��{yK���Zk��;V�o2��YݐA�]���޶�l��}�����[�D]�26L�8˸�䖥��ns�oC5��Q���/])nma�� �;9ME];z�>���r��Uc���H��OY�W�Lc[��WF�	����0�e�Qe�R��A�qus�%nG,��򇈠����4�f������Y���;��%ʤ�\���QF���S5��HZ�W��[a�:�4���`�Y�E��Z_)�q�i�Q1�2M|�e�����a�����r�&Od�Ϡ�|"�|�����1{���]���rL�E��aL��G�_\���65,�WN�oyW�4em���k^e�����0�ƭh�n��g7\���Ö��:��i�?K�B�>*m�@=�v=�u*�Q:д��4�Om�J�.)3�����0�Z�Ғؚ��б>��k��YDf�����B��@n�p���Ua3����W��@�aL�E��״��w��З�//r
�Y[c�a����mtE�ڥ��I:��fV=�L|��,ܽ�M3㪶����|ZW�3�7��ҍ�ok7r�#�l�m8f*�ͻ7!�+m�2�7ݥe�v�a����ީO9)�9�.؉J8BLٲ����>���4�aH����ʠS�4�I�N�69􎪙7G^#��C�,w|�1ނ*�j�(I�v�룹��B�W\��s������goroW�\�t��uͭ�)�@_h��{WF�%�����o[V�!՞�W���4^ݷ�J�����#g
�v/8��Wڵ��%���&9N�b�]7ky����K,�5�>i��M�k�w(�=�ѧF�e��UeV��n��;(k�i�5<1�)�g8W�b/���QsnX����«q�6���;E��S�N����ٲu�ֆ���Ǌ.렾_U&4��!.��b�����A�_4D-��4�����X	��P�uwY'l��ܼ|ȶ�c�d��87B���m e�˝�Mb��9�U��a�H쉌=�}�s���Z���G��&X���p=��0��|��߻\nu�i�	z�������dJ��48��1��s���ut��u-,�h�t�96vvr�ip��^��{����4s�w�B�b��$�퇞�E��p�{x�[��e �'/�;b��t���.|����}3�D�u>��(�P�gv6<sy��!ce������9L]�=j��N��j��D�a��������c����#R
��L�.�`.�$�k����Bv�<�}	_�F6v�ߜ�����Յ4�w������b����.�5G��+���jj7z�c�|��۾�m��AԚ��;�yn5��Q��}6❸�jjc��E��A�/�L�/�\[�٭�.S��};�f���;]h��[w�/ E����!��.M��G��B�ZUjGΏ��Ten�3��j��v9��t|��T*g��և�%{���U��!&������됾�e�7Sk#=.���TN�!��9:+�����WٙqN��5���)ޡ�L;c�PvW֩s����1���F]��z�����ܲңs�˷�>��|����9H[y�\Lc��*�ޞE���u�cVF��9qR󊏶�7w}N�P�U;��i�H��áʳQ���`z�{Ӷkع�iB5��rMB��}���m�i�b��ԛ�B�+��v�[n�ah��+Bޭ��Us��M0��e�wI\�5|����w�=Z
�5�ZG(1_K�/�a�n�Vҹ���@�����G9[|o@��q�.u>�P�_\�����-ú��)w	d��V�=͌�\��8�e��p��t�.�N�Kä�m@i����Y�7wV���G4ըsy85�K�;$�a/x|}�F���[��:kK��4M�NEǛ*d ��Ϊ��^K���f�<��[ְ��&r��-��7`$�^ض�4�b��Gg]]|Yy��{q0'_;W�!���G5�}ȔѿIO��E�+r:�uj�jf���u��R���ki���@އ/\zNPo�0�ɠ��4�J�.�7�=���	�/FksN�.�n:���a�*����UKFf�O!ܰ��Yo$����k�)�@��:SµȐ����*�����'Υp�_�wb���;	�ᱎP��[F,�����ⅺn.��=�6�+!ͶB�q.����r�����l��<������pF[o�N�<(��S돵%y��>o~iԱ�=I��z���2�ZH�~&��,��S[k6��<0���\M�{銺�{��s~0i��x���{f/D2��Ӧu�}�m��[� p{�7��Y4����!G�U�z�i��}��s*�ci�kN
�b����	-�u�NW�2Ʊ�'{r�6�����(\y��G>�S�|�~�!{��p=��وVV1l�;XޒHM�_1n���l,(��T�c�eo�Z�����*̹�;�t٦��i-[�4�2f��*�ێ�>���;Z���3�;���GJ,�Dj�K� =V@"��(f�|5���^���GV�^� 7uf#�qM�)�t�y{[��6��k��5x��x{ᩌ�ʥ��U;Wch��䡽k!��7[&�"�8::-g-s��On�
�EK�w[]�WnӂBo3sStuR�c��m��Q\�eƞ�9�?�KK�Ys}ui�@��������|��%��gs⩼��e�hN(��:s��Ю�տ3!׏w{�����m̛P�X�f�ҳOP��V>0`1({(�U3g/+P�N�����iX"�6Cd��j��i�b�s2�pY6��{�׳��ya��*�etE�����QԽ�LQ�\^9j�D���o�jL6�ś8Դ��2u]�ݿ�����9��N���o�ќ0�4�什��q%YE����p��&�t��R
��VT�|L
��;���l��>����f�Zy��J�}c3���K����x){���l��
�+�d���L�gz�7]u$3�G�ڻ`+��6}w��Sʝ�|�O[l.�������JV���}�ڶaX$�7N0����6��+��'D�5�%X?��z�K�tf�=^�ۦW�Mx�-ƴޣ���qu��5��y����)�"b����;��vmtU���	����=n�6��������S9B�퍹�IӴ0�EV��OF�2+)�כ[�p�"<�g�1'j��$��^邾�׳��[�� )��b�	�8c�v�����[�=(|�u���f�~��VYb��*��D���ano���[f�q����	A%,W]��0�]�Y�O3���^�~��1vXG�r�U�}�w�	�er�=z8����\6.����dF����_.�#���6w��F�O��:� �F.�h��d&�mV�!`V ��U-��1��b�L8�/Uر��?-A�\������_^A�v��=d���q�򑔷wH�͠�����J>�N�P_e�/�|y�3�Q�N�{�.*�Ӕ�I�-�^�P�O �X�L�PK�'�f�(wlś�1��Y�)��e_a&����׶��]�Aqy V/��^�B$T��Wg�پ}��<���G�.LC���oH5a{8̶��|g^� ���Tn�ܣ���#��㇩آ�e٪˻�r��\>�.��8�MA��F�0�3�p�]��z�}�e��a��j�Iڀ'`E�L*��/�����C3����ˆ���U�3��e�+�ؐ� BmU�M�j�CЖw������=3u{D��6���PTΰ�ljl;L1#(\0D�旚-��,�A���ϰ�V�;P�F��.�N�{�#\h����"���V����`�,ɓMjS��bT�0H�W�9����}.�����O�L�UF^�មZ��W�)R����&����'�gh�=�YS�\��:���GI��w�C���Epu"{���٠6wr;��7�鋴S�kq�q�7	�KSL:Q_%T:PD�/rw���^w���:���dS�~�y�Y��sz������m���$;�vhz�[��n-�&�9c��5`�_N��'3��H�1�eb��Y��R��fė`w���P�E��Z�*��WT1o�^�f��������$;�?<���+��� �O�N�c�YBf�H���C }��_���0��*��<�7
�.��&Q�����sY�Y�+IH�6N��:ql�Y�Z�aOZ@Vb���é�놫���qb�q�����&b�Cg]<�`��ɶVaϹ��7޼�y�G)��d��M5�A���,��S ��e�0�aN�L5���wIIR4���U�v!v:�a�c�t�(�;.����C1}�;�s/#�Z��F�����:�2��l�İ6V<�ɻ�{�{�<��tW�����=����G7�빽5��}c�D�v��,��v������wd�B��x�Aɲ��{|mޏ�R�b���n**���>��}�[ꐩ:���66s��æm��pJ�v�il�Һ�egYxѵ]�1f�
��ݖˮvfb�.���UtZ��B�b6�Sw[RdJ1S����sh�ܻ�-�|�R����8�{(�8�UO^f�5�-��%����ۧ�`�s��HSwF���.�օl��MVv�Ԟ�8ho�O�7�_i}.!¯�4�H�н�]ۚn��t��B��ך�Zk7��Ra����L����L،�2�&�la^�z�+{
����`Th�~��׳>��Ȁjp�S3��kj�Ѵ0��t�3b�����5R�訓yR�#C���58�hU��<������S�f�5����	Z�օ�{���.̚��n�+����7��H�;]�L��h�� ?wH�Y*َ���7T�9U�ܫ�g�P�E�WǤ4��Qj���֍�C�*�ζ��b�u^ې�ݭ�Gi<ҕ�X�JM��@} �{�t������ �֜���=�Rq�A�6�SQ�s{��m�wo_e�m�لh�G�}��Wmaq�ƛ��2
{z������6�F�?yV=�ú]�.����ܞZz���/o$k�G!ܓ��ڂ�o���/j}�v�v9���$&+�K�T�9��+@ir�,��{�[�[��{��-p\xE��v�������.��vv�'�޺�Z%�,���t�	ߵf��SIU���9�����{q���YD�cޙ�A�'Z,�o;�pm׼ȘX\į��Mx^ófv���>���3_�r;;\�`����`j��YrOuR��Qb"�~��<a�'u�7\��
*��g�Z�6��3�����Ȧ�玢Ԧs�}[�=ܓ���lmU�3���1��Z�e���6���]<��j�>X-�nY�w��&j�G��q㫸6���jt�d�YRR�4�&�tY���z��d��ȳR�ӶV^�q���r�eg#X���8�_.��ّ�����\w��e����| (��s�%�ʎ�<d��q��on�3��#�$���{|g���R�%�����_of��\�z!x1�r�lg���0�QY�곯���6A�l��
�Alkࣈ)�$�����F�������"bv�z�n�|�~0����٦�,_s���t,�MC8>�>*^ٻ��v���7 ��1j�`�jt�����v��~&�s��
��G�W�������W��K�?{��?��3�?����~?�������|>>����Pk�_1��b��d&�P��m��&�H��-�:�"(����pH_�T�9qT�A�#?�@�a$����K�e��d�a&�i��e�j8"����TM�nX~��GFA�j��y���[6V3����/v�YO���}���ZM��	�if��ؙ֦��d�T��d�f�T�]���6�^��5h��V;̬m��B�"��ν�#�����ù-�[T�i���A����Y�x��qY_�?$�c�V�-|z�u�`�v���F�N��z�N��G�2�5��_�����x�����l�
�����.�fue���3D�����uC=�!S�9mMެb��-:dL��s{�b�U�|��<}�`�#p�ʗ�����EPfm@�vU�u���-���>5B���i�E��O��'mP�����c �u���Oԏ���Ƿ�����+]���_cO7����d���I���e�����-��ی�/�����Ӯq���J����a�I6���6�I���ۓ{��w7�z��0������0w[6ڥ%L��Nڹ�Vs��5N<�:��v��N��D�2�e@��5�t�u�xlof�b�pWGJ);v�AJ|���Е��0^�䅝����T�o\oY7���,ͭ��o�q�-��*�d�]B����c���5������E�¸�o|d-����uR�VnՉE�9�\�H�!P�G1��i
'����d�dOs�cB��Kgۨs��F��z..W�$�v�^��u\���,D�$��p��1���J�b`�@�����,~`��M��j"	Dт!!���C!�L��(��p�i��X��["�a"#'�< O 8������&��IB �I�2�,7��b	�q��H�'�O����e����f �b4Z$�����M�)1�HGW\�\��땣�{
K�4�UR�!My�W6i��.Y�ē�E�h(��kED�t�.���[��馂b-h**�����h��\�L�\ت��*����Y*j��KI��+�X�E)m���b
b'X�f(؍�����`�ĔE�8���Uu:���cQ,T�V�1T�U;:�h��U$�F�MV�Qb
"uA[`�*�j�JՍIE��E���c4[h��QMPl�+��u��;S�ry-��(�����MQ�Rim��h
h���UIA����HSRQEE���m66�
�SQ�-q,T�P�QM�UE�Mmm�63iuQDDQDb,j���9��LA��DSELCM5Tm��ScmbF���H��R�Z2UE@kj�8�(���$B4 ���iI[k��($��p}��Ee'�5o��7�]d����\(�Ԓ�1�nL���ެ��1u4����2Ŕ�����*|n�S盙�',�ɑ����e6��\�p��"�8E����_`��η8����5L��,���I���&�y�EI�}��b?a���5�����nϰ�N����G�� 
�;B26u�7�L��0z���٦�u�u�N�jt��|{a�0xF����x�D�c�f7Z+�]��fȣ��o:����մ
�E�p}P_ϣg����r�EiۖNZ�ޯW������6W���6���g%bߏ����g�-0K�2�|nQ˾��(����g+�s��O�2�"��X�>{g:�����ts�yRe�lߧy��Q�'�A�}�a����`��l�3����n�Zݓw�c4���͙[�I�{��s���v&P!u]a�4W&�KU������K0�dFNu�F�����˃��Mз���*�V����i����|ޱ��	�m�]���'�0~�_{g�?��sXO7q���@���8|���i�%�ǣݶ���S��![DL=f�t&k��훇��]��ˮ�Г�4^�9H�6���4>�$&<%NcȽ�M�*��{��b?{�>����/C�M�ɑ��nв�c�[[���ll��g�f�[L\������4U����Ģ8{����y�U�'ޏ�U�)ӽ����Ŭ^���]��˱ُEKwG�:_���E�^��K��>�^]5���K��ʔE�u�����W�Ǘ���8#��$d���D�VY�"�ټ'Ӳ{�{ڸ6����0Ow�?J�վϝ鿕Էe*�O��$y�^�g�Ƌ���s���xIC��"��'��r�g�R�ҥ��G��p�g|QCh���"�O3���� u�":N�-���-^��?qʿm�4�&!?g�|/l���}����^1l~�S�<�9�%���{o�۠���ͣ���0w /ް��9p7���׽�d��s}Z ���d� �j��z.\��}��>Ч�[Ƒ�Cu�E�A�}�a�����
y��$�:�P��}*#=C����~�{M�Sw~�.��٦v�Ju��qOc�u�Y\OD��U����ovf�7�^��rA��Ͼ�>gb���)�b�3���}����Ź
��׹���U7β�<�~t�&��ْ�&uo�x3�?Ok�yO|�x�҇Zu,!����[����{g <���F�Ǝ�{��w�LPnb���9����e���(r��	,j��^v6����dy���q�s�������������@���7�<�v����%����K�k�������8�Y���fŴ��x3�_�/LxƦ��f��~�kE�����Պ#=K�{��Ţe����������z�++{ٞ���|�<|u1k�S}#���:B���c��Y���o�n�j�I�ga���}(�w����s�����z�=+����]��H!��?]����V�N��з���^��?���) τ�xc��x��_N�T�����l��3]����\aV5�ME���W�*mf<���H�r���p�$G���:.���#�M���<�(u�c�7n�N��۰/��J���U楇O^�.��s#�-ԛt궕�}v�%sm��s6��^A���g�o~��d�e��%�7��s�N�(��0���ȓϧX�k4��Ww���2��s^g����c�k��D�vj���̮D.��w:e�1J��1�3n����o�H)*m���&���`'����U��=�z�*��D��D50��}ݓ��7gsO��7�	�&M_�g�}�i�oQ&�[���ҧc|'c�Y��w�콖�O3���Qx<w~/�>��2�����h��O|C��	kh���������ޒ�>�з�%6S��)i]�xu�|<��`>g�¾}�=�o��:nyo�f��Lo���~����t��$>z3<�<����Ur�^tu�j1w�/�I���$���b����;>ߜя7�m��t��ʳ�]��p&m��iw��O��m��\� {@����	��M��&;zc�lܹ�q'ތ�;�D�����1��^l��b���b���9n��V��yx��0��^JǒG�{�k�2��/��;o����q�ŴdV5TU������a"�2�oQ|�引�h��aH�;�ϣH�����r�J�a�wr�r\�C��ep�(���x*Z�V-�۹X�z�l�°�2wikJ��L���pe��UKU�pDuh�a���x{�c��VU������"�:�v�N��w�
f!��Vh�}b{�]3 r���ٚ���sP�x�/s��G��Ƽiں0K�:X7���{ӛ�`+�)�c�ּ�5�2��|�Ò���g����c��j�ާ*��@�{b����^���O�1=��!�|�s�<!=�0u��Qy��7�{[��H�{������9�x{�����g���1]s�W'7�.�����_��c���j6}����f��^��Tnc���s������d�S	�TP���_�g���p�:��{��x�Ɍ����zx|���-������ Wv��z����<��[ n��=�_Vo�Ɏ�u8~M	l�&[kd6z�n��u�=���l�s����y��m[N�9s��}�$�&Om��w�<�L�(#C���c����.��ч���� R2��nim30�y�@������^�0v%�ށx�u��9�ɒ��_��[z�DJJ��o�ˍ��W�Z�z�v�JX�Ј��r��|u����%�{�2Ԛ�ۉ�6XU�m�.�ve27�͑�,�sd���U^>��8f�F��=�S&��;�湽Gk��O���]�{q�k;kټʻ�W�Z�OG��i��e߽/$�-߄���|߯}����A���/n������cU�B�y<��(�`c�������mﵓ*y�L���=���qԸ��=���p�r7�8�s콠t��;�;��}��sp�G<��썬�_���ɢ�� bU��Et�y���Mv|�aq�mR�1O���#h`|+�<'���R�wO��'�:_���W!s��S����/;��s������_��`�Ab�!�:
��ճ�ˎA��i*�¥fpu>s���k{g���x�9����=�9ϻ>w�g�N�Ϸ+�<�#��� h��pl��qs���;4h�=u.f��hb�Ƥ���0�,������,qj~(���������t�ٷ����7�U.r�1^���D͎�7u5����9�{�4�>k��k���2��fP~ԨT�n�r��z���cՙ�4-v�[`�c���'gH�
b�rm��U[:	�`�a=/scȅet�b5�Ѥu^�W�p=/����f��u�Mu۳�}nA۹4�"��n�����{��y#�B]�{}�ÎzC.+Ft�Ǥ�5^|���3MBG���~��x����1�rsӏԝ!�E1�	#���=,A$�y��C]9�q³+̽���'�Ñ��������o'������I� ���-��ri�m���t�J}����\<��^7;���w�uzLp�񹦽Ϳ&�B{����mu��y|'σ����{��wK���/�Ym�����~��p>����V�}>:<�BK'0g��'@9��W:=fW���ҫ�U������{L�����;�/��<Sv�5p�qk<P^����.	Ӽ�̯����
w���Dxl86Wy��y� D��f߻#�q�-�a3��=2�N�%���6P�]U�V�=W��<gQ]>]ӏ��E�g6P;����r�h�(b`�c�}��Q����6^��5�S��&�o���zt��hb$].��њt�^���ؾ&5�p�-��4.��қ7H`�[��*��@����:!i��2d4j�u�����;��>��X7�J������\�'�Tq�D6��lW���ٍ1�YӾYo�u�hl�롕�h��g6bDu�) ��.yu�r���ޮ�F�ؤ!	;�ᜲ�	w��w��[IZ�������m{o��-di��(���������y~�]%尡C�ǽj�@���2�L��Ṙ��B�	��v�'����M��_f��+�n�;��rɃU\MTޜ2_5��ff�}����i�k�L��<���`ޭ���]�'\����G[c�g�l`�-�F��m$�9:}7�~��/��������B�3ފK��.I�4\�!ψhL}�s��,�n=��Ɣ��m\����>Qx��k_x�v�\G���f	Ӎ����{7�֫o����:�m��c>JZ|��>�<�^<x)Ӻ~yT�ߞ�#����D<"PZ/vu�cX�gvd�"��e��-Ք3 ͮ�nEG�)�hy�/�n�.���׆β��4�O�<<7���ȉi�NwZ=C\��l��؂g�C�ho��=/,uY���u[�8Nt� �Mm�K։"u�}�߲	�7�1MA�c�����{�E����Ѭݾ�a$��4���{�=��{�_�h5KEaUP�+b����g`Ϯ���#���>�ט�%�n��o�f�8gٗ��[��م���g���]e��ɑZC�ޑsp���m:w�t�u���2��m�6$YsLj�"��{:%�~#�c�C�L�$�nv�Ҽ�9Gd(�������o����\�%���+��t|%!좵�`����b��-_��F�̷8���av���릆>k���U}0߭+����]J1t#G��m漣���I��g�y�C`��L��{�o&1�wd��W��y��Z�����L�{����7z}��p����Vn�p:�.>�$��\��;az�/���7�Wahܚ�����<A�Ɩ�z��'y���^a���E�&�#g_���Ϩ�.z����z�o��N�w���}T`u�a������!�9��oX/:��F��[�0P\��)�ʢ��z�I��s�޾�S�?!�Kr�D�����G>hܙ�&�bXTo��7ч_c:�.�����Iͮ��%ww|�XȅIZ�ԇ7.P�����/�4�����s��*	�G_n6�{��;�&����HÞ���8��S�����%�g��E�3�`�>�-�fu�ozXʣ׽����1;�.��`��2	&[ke��φc�8[^���l�8�.u^G�b�5���:�='��;g�{��0�a$b/��^zsz�.b[�[��޵��h��0	�w�oN���A���Z��Ȗ��{:��������ݞ���v��D&tĢ�z�7��6����>�Ï�W�+t!� M0�y^`]��|�;$�i�:��\��f��i:�2G<�������|â r��:��\��/ޙ7}�ifmc�412V{���T]3�;���y	�h��!�`���-^׼Z����ԧ�y����������K�d確�8C�`�����w���������>>>>�w����x����~�H�t�1߉׼��w�����䣋��]�o�@�x"Gc���!��uu�V>�чʣ���`t��L;K,I���&� ��gy���oQ�^�7м�����\�ǒ'�t�n��n��L�V�u;.N�&V76g�S,�V`29�%	[c��{�����{c�h..L�uO1;m��7�0y��'�B��v8�Zy�	�o~ڶ0��.�ic[:7����]a��d�%�(�i���F�v�S��g{H;ɱ�ѻnE�!�#]G��A�u8s�2H�i�F��dΉ7x�K�{�K����qZM�Cd��@�aY���z�sy�a{|T�b@�]���g�ݷp�uҤ��G��i�x_�f�i���H��%S�0���C�ig���5�_�=�?G�Y��Zr�ݮv��A�a=���l�Թ�i9̎�D�ƪ��ڮ����G!��=I�#��3��ͽ�ޡ��ָdV��GT��}�[�sT�5vٸh�z�ͳc)C����7D��{vv�DV��N��|[���s�p�!�v����,%n���i�0����{��[�U�so{xjV��JfK�`��s��7�z2�'�7w�ͱ��(���>�2���K�6�<��#63C\ꄍNCj] ��i�Q��7�s܄�-j{�t]�f�N�ǡ=�D�f8�*�4��SY���j���;KY��}�o�b�'~G���]�c�Ζ���ݸ����>���y����f�����Η��X=8�mF��w��?����R^�����T0M�r��o!Έ�yjһ�Wb�>o�,l���}0n\�x���gRū��c%��8w�N�;\գ7~�{�#Xf.�A�p/p�u�?�`x���������j7�&m���\����v�N�}�^���U�z��8��&��5�2`���H9�?Jv{����h}k[2���a�􂞘 槩��ט:V�rks"�U�5�����M�zfT�bm�gl� ��ٷ4��#L��z͚�b�m�J�=Ϯ�=��K�0���r������Z���蘼�O4V쫺·i[���'�+y�VA[,W�5�]�Zq��0%��H]�]�}]��̓��r�@�_���=f�q�QP�;���ǦS�����CC�ջç>��/n��2g.dُ�*�)��̕�����rLyӛx.�C"��B��)�4Pb�Y�EL��ܺ�6i�_=�S[r�v��`������z�E��kA��Ǫ�L�f��^��c�Ђ\9���/W�~���3н�V;qLݪw|�����uLDq�oE�;.���k�w#�3QRWL��mr]L÷�o+++:j�1Kf8[T�E��e=�eݕ%�y|��Mڷ҂�*��l,�h@�;ã.�#yw�6�ʫ��s�_M˜ة��f�@�3z�k������n}�dTA7�ũ���5NMf5�����EM-I5D��{�sb�*6��r�ME\ڪ��PL5�TL�"֢���4a�����Z)�-�F�L��U1�� �kE55U1�%N���*�y��i�l�`�+5kPcf/1�4D����`��4F��ƎŪ�Q�#mFڣFy(�������
li���*�f���*#X���Z*&4b*������0r5QR\Ɋ*6�1Tb*՝��c�U&6�m��熢�yRL]c�
:�O98�ֵfqGFM<���(�bs\�s��Y�w[�g���1�U��u֢���\樃���s�Z��T.s�ؠ�#p�华X#�1��y��"�<3ns��8.
�l\h�Nyu�Aθb+����č�'\5b��b���n���]i"8�8�����G9\�#\�')ֶ�lD�ñ�ۜ�mrn\.���\�n,����W�V�䎮p�m��9X�:��-@s*8\4sn[�b�k��UG#I�qE[��M�9�z�"*��b���V�h�c��ն�����¥��_��s�{�~�(��y~�eM���r[�V��kó$2T�Xկ8��s�ۼ��hЩ�/��n�\0����e��O���e1=�3�s�a����L�1̛`�t�!� ���� ��N�Muc��u,��y�
��]��	ϯ�¦�x���=��OE����ӻ����$�4VPB�)-�l�FlZp7�2�
A?f7/<>�U�m&ae`\Y�x|�H�흷���O=ɐ1�ڒ�m��X�[����3������㯶�o��PJz޵��xȧ|�mV{G�U@c�N�zGq����M�S��ڻ�*b�"�+f�ؔgQ�1���o��� �f�q~�Hz��o:+�'9�4+�.fN�댍s��>B	�O��Fi�W�F�]�n>5�l�AJ�py��9�N����TD-��ٝJsS��7YĎ�*�����>>ħW��)���J�[X��Z�"���=�oM�+	>*�#n�s�v�х����f�tWC0]��0�}�F�|s����-Z���c�Z"�sF�Qn�黤�Ǣ2�����QC�"��Ӡ��:[�L`m�nO4҈T�"�&�~/I��A.u��%��=��׌˫�s
Kf�Hr������Nτ!ٺ�μ��U�0����?��J�Ý�7nͷ;�҇�嗢�gݜ�z;t��h�ңЇ{"�r�V:^��w�ѕ�h<����כ1��� ���s�����8K������m�2�)Y�L4�_[�OEN���(���l�:�����"�{�q52)ZQ*��{{b@c��ĩ�w?e�����#�@�;��`	wn|gaA��n���y]�6��SX�o^���5Wr��T`�Z�L�K�Y��y�s��NF^2
��i��$K@x��ԉ:���ɩjّѵ;zz.'54>�om6bS�1������/<����G��d�q��o�ͻ�[jX�o�d��熶�t�����i��@�$�ߙ��r���_�9j����g�t����/b�TB�؝�#�� �cZbac�R5����/�Ag}f�˱n.;�D�U��N�d�m	���;g�%��2�������������󣋳Won�7-S�3����
�[�ۃ!�tF~�ߕR����)'��I�|!���ߓ����v�}�o7�=CP��<��I΄�+�R3��3g`)�>zw��k�!S�0��Mඁz̞t�*��S��@���2{%�[҆�b��t�p�'��hH�3��{k�������|>b��ߕ��T�_�1V�^o5tu��ƻ-��MQ�A箈A�=��Ru`bT)\�,)���mm#z-�������F~v�����b�l�w�$�:p���I�����!ʽ<�r�Xu/e�V͖L?�TQ�t"k��|��a��6���4�-�|y�N�v*j�^PtdΊ5��ow�>���Mʱ���6�Jh�����7U:
D�VeY4�^�f�<��{�`t>����<���Чt^��$���� ��xk�1��ry��vi����	�{)�F|)TS�o#A5��)T"�[VQΞ��Σ,l[A�t�zB��q��[p����!��T��0?�fw��B���`����[R�u�^如s_C�[�	��*��G4�r��xr��c�C�����+3<����+{;���U��Rޛd]cҴ���=ҹR\W(���ܠk��ʿE>~oNy/q��s=0���n��3]�f��E�Y�����O6��5�v������2\>6Ϙ:nob��y�־Z�v��kU�N�c�����.�TXZ��S��֑ �MV�z��|��}>�|l���\�r����=#���Bը��:�eҹ�r^��Q�Ѝ`!����L%�,ۇ��CH��s./h�3?	�68Գ-�v�a�GR�m�Mk߸ð����k�]9��o"&��;A�\�� z��gRg<�=�ȉ�	�;���2��'V;����rxM���A���Z���ذ�.R���8̻Ohv}���+ˋK���<�j|��6nq�o��Y��s��78�5�;"��ET٢\�+u>
]<1k�	��027mqL���_[�.."�8k�t���{�,ڂ�+	yyt6���s�m���V0mVS���1�:�P��iW'�ڥ��K)4�C���mT��j�L���k����>�,��(< ��TG#.���U�:��Y�x����E��Lt��Ǖ�(�꿳�ߥ;�f�^������� �x���F��q�髦/���E靼ۖ��i�eW����gkw�pl.]�kߦ��2a��jR��A���)XJ������xt^d�6T�6���OѬ���?�qD.G3��mCǑ��d&UiW�'�	i{��[k:v���!�ǧu��=�� b�Bq$>T�HOex����k~BS ��;pcL�� f�l���w).P���EP����5�׭��Cj	���By�c@!���2{�La�ɤ�W�/�μ���'[�Q-i�7E2��&��(=��z�֏	�DB`��W�zݳ�&,�������'���<�EL-�]`�L�uv4�r��kÇ�v�����bM�0�C(`nm�0)�4(��'��]/g���W��]&���F@�y���}s��c�q�[��l�ܴ|�W��2i���;4]�`X�x�>�C�?sߕ�/��zVl7�bn]���Vu���.�)�1���kv����^�-zi<�(���Q��x�4�p�4Ɲ79w]ܯ�v��U$��&C��y<�,�s%j��c1ѩ��MJ�u��Sz�h�Pʪ88"F�w�II�B�u���j�l���$:�`�ӽ|��^���I����3�8��Ha�����f�U�QkejUk
�=+�	���	���E�+��ܛ���K�tn��'s���t8s	��P4u|fFN�Ζ~?�c(\���$���N�]�:kA�6�l#ӎLG6��f4�O0J���4?����[��6�e`�[�<+54����fT����!� � LW��b���GD��ż!��eL
���O�L5v��0N\(��׍{��M;�������� ����>/��ӱ��a�s�Ϛ��n�"3S��r��9���zǣ���4��h���,x���R]����a�\�\+��.��OJ����O��,= C��|U���%Oӕ��4&��+f�;(2o�Z��KV��[�k-����ٞXe �t��q�,�a}��-Ucnv({.m�b7[��m���g�֣fٲH��뀋wl��њObQ�aC���Ve'��Q����08E�Ǽ���&���V��;�q� !�=E��	Ǝ1,���\�I��7��<�ۼH01��ol�ǐ��6�dv!5X�jN��(�eś���+���=�B�w��o�z�F�65zM��"7Zt�e�O��R���8�80���/����.)��:�G�����K��᥈��k<n']��/U��{\|�և�U���=���{�.͈Lk;�!	��O�)�|��+]"�W�T�Omq>�k���bX`����涰Z���W��lg��&c>��`� Ì�u'�9�NV �"��׈��6|�LUJ��ft�VF�\p�gy�<��G��-�&86�ܞj/~:�k.����'���`Ӭ�9m6f^ �h���B�׊א�%������G�J>��p�ˢ�f��i����N�"�͑�]�f��n�-��Lw:�H�6MA-Q��؟T����O�h�tޙ���ɔ�F�3P���c]��L���b2[�Ҫ<fa���ݛ4l0�<����t����o�ns���~�f�%�ܡ�hZ��S�1�����������`HB�GCoM�JŒ�qb՜��I���x���?0:��橗d��d>��NF%��h�	�-C�9`)d���S2�z��)vD�(	@E|0;(������mA��wPny �\@�.�8˱`1�h�F^�w�N{���'��:���q��~[F��g�I�ON6ۜ���i�3���{{u�L��?�����yʆ�r�Uwt���Q�w@�/��x�O��k�������d{��!�<����V�-�Q�3�����h�'���1Iud��F�SJ�QKNԫ������ci�p@�c(�"þ�)ႋ�������|���zq��{���.��tM�3x���bT�ŝ\�g�ƵXLT��_�r�*�-?P�)��y�>9�}�-Y>�4�L�.˼Z#��Ku��e� PY2j	d����=��U��_ʿr����2�������m?�e^����I�W����N��s�XզO�xa��C-�H�3ю�Ơ2��͸f�,��G�;4���R�ggн�+C�qp�P���̙��fPe{^��JD�%Qo
e��R!��4�lF�vިl�QK�ƳǤBoA�,����.�#�Ħ���L�.�w�4-?�6�!��^��ֽZۃS���s�[�d�J�ӭ萄c;"��C)ۗn9��Uԩ2o2�[�[�p�t���ls9n��E�L���C�[�xN�!��'���#���2oWv�P��vm�Cgl���u��JOV��"�<�<9�cw�+��A�+�*,|�R>��ny�"�6ED���w;�n��5�F�m&Ves�P�r�̈́���v�����K���)�?��4����Ϸ~���Ķk�<�(�гf$닲Uo5]<�o��XH�����=�p3����K�����Ӛ����|M��ɗ�)�5Uէ����{��\vX�V�*��-L,$�Z<�h��}�f��5�����wm� �I�����\z5�x���;J�KV����^3���CWr��F}督��l���KM����k�����x�$�F(O�C���<ŵ�@P���m�2)r�Z�2�\�YPK�Z���ud�����AOS3��ba����k >�?5�l,Nkj@f[]�XsQԨ�k_ފ��SA��0��Y�ї	�CvgN�kUK���^V
���I��	��omu��Y'W�,��2���a
�3*:��o5�`�lN�q�cn1��D[��^}�)?���C�(��a�2����B�Pt���T���
�J�@3ǲ3�A!��9v�tE��{�m�n�C���c�wt�;�hʬ�]�
*����^=���֑����%謐�F��q�逯t�æ�G�Q5�/xZ5N>���L���)Ĉ��Obj1��NT�6�c����֮/�KBUz�����p��`i��+��uj՚�}���Mm�&;�j�}Z�(�'j[����`!2ot��2�̘5���go��{vH�x;r(�f:�=[�H��v�֜I�0/��4�%�,t��Z��L���o]���	nC�%?%�:�,wkZ~��X�Y���W�F<>@W����G7=f�F�CK��Ȥh��vcY�~/p�5������AYׄq���Yz���N�V�u�]3y)���w7 7�e�GK�uO+�Y���~�����$��xLf��@ҭ�9aOU2<�8��_ eC(��f?"�E�О�h����Z��2�ʆ��:mn�٪�������oP[��i�&�������ӆeXĲo&X��RJ��q�{���mml3czN&J8K�r���_J��	.����q�B��F{"���JoX�ʱv�9jw��-�%����;�hN��:����ʐ���ׅ;JU qWK�zO��(,it�~`6jKt�"�eXg$Y�/³P��5�|��̛Y�}n��.�56¼^ˑ�y�]F���u/�J��e{�� ��ʌ����I	X��`��j��C�0e��=4ڬuo��2QS� ��53r�rb�;3f��vk�[gY4����XE��=w	��Ӡ ��c����tדێ��o���r�)�e��X�t����(�{��}�7�k �K1/M�gb\3o�h�\F�cvz�y��i�U�%�T6�ݟHv�RK���ID��;D�zN������eP�<^�����#+����b�ŰdX$�J��{omy�$�k��X��K�I�D��S����q�t��˥�Zộ�:o8wK�a�r���!4����l��=c���C�w�F�vIoU�Ayǔ��b���.�A�~��_$�酝nB��;N�`�Aziv;)����q�ߊr�7��Ǩi���~j�?.�o�X����.$�I��c��U��<�UFa��=}��;�]�j.�M4h�|��H�P��#pW�,Ү(�t�s�����B�c���>a�<�=���ۤsg�����Ă�u��R�0j�;�	�%�11��te�[bJY���f�{e��{ؠ�ev�D1@��j�r���>U��?��+���,/���fp`*���I�g�I}�V�����z!����'lyt�ɀ�-���[�v��<��rP2F��# j�d[�އ�<�O|�&���-{ei������d��3L�Q����kl����=��4��Zy�۶�;�htO;6SKLv4�$� ����>1)��ˤS*	*Mm~�<�ee6�٬|+��tڞC��y�f�;B>�_BG��d�q�&Rv/)�����������3Q��'�ףU���[e�q}������!��1�a�0��\��i�	�\�w�8��iV�f*�Y���^\�����<z<��[_����r9�6s�VM77�L�F�m��Z�
��\����xo!J�YK����8�;�{��@B=�:�?s�2p8���W�d�6�ŝ�7�e>��"�׌�ƳГ��ɷ���/�c�RͻP��d���!��{�^�O���������{��>>>>�w�������>�73�nE.C|>�}���քG귎_q�c��'�����}>ߞ4�)�f�r��w`c+�z�S�c�'r!�`�A���XC��s��i\+)����O�A(20�]�9�*���~a�Ǵ���mR�ݥd���JqkI�@��#�p��l�/��gq6��mNŭ,*܁m��;5�Ƈ� Β��c;��E}9��J����ү�Հć#�z�o����xw�I9j�w]X��ʣ8��!��᧜�5�S����u�$���u��y#c��|0�ο��΂�����j<O(����r���m��.��Àk�S�����=�}��͵�#&���}�)�D̔�Ku����,Id�Αj��}eiws���Ǧ��Av�efy�`���o�W���D~k:���>>^�ϭ��D��0f���吃���KK8��U���+��譞8���O���nq�WW�8��<���=��bc��:|^իh|�h=�A���2�7PJ�%F�$����2ow���w2��m����4m�[�v2t���&�v��3VZ`�\y���)f�b��{�2ރ 
\ƆjԠ�!�w|h�=��ՏQ��=�k��s޻�X��k1��Х{(G$9��'���e�j�f*b��nW�}�d3F����Ϊ��`�`YxS��{�)�I)@��(f[�B'7LT��FI_d��� ���㾬t��?t�41����<I�����v�&Xyh"�C�~[s!�O�L�*�R.� ��NK[���op�P�&��Im��;���Y�r,y�Vnx�ŹlwZ���'�S�3oD�}[�sml�&�˛ׅ3��5]r��u�6��Z�t��6�a��_
G��w}�v��թ�aK�=����E��k�ޞ�4�����l^|�@�N�3N�C�m��tW�FTp�-�W�;���Z0ؽNwM����l���Q�Y�UrF�<�P̓]+�訸y���@�`��
�U�6!{�tq�ц�c�`����@��5J�h���ص�	�!E@�b�I�&�$�lV1qY"�en��0��\�v�*l�U58I��eٳw݊f�V ���ܩ�'+K	X�- �b�n��t��M�;��j۫���FjWG���D7�����Ӈu�:�C2C��[ً�ǥl��8ˍ�>��v���$�/�J��'��W�=�������bUS������"��r�˽pw?�6m�t��ON�_?t�o�Aޭ�#l�:���N���O �ӳ[�6!T� ��o�-�]�� x�{[O�Ҟ��{���7��=�W��8nk �z����H�-M��{���D�������.EΥ���\���o+�N�jt�y��x���7vV���pH�vVa���v���s���xE�}�W2���zz��8�W|#l�Ľj�B���N]�J�ݺ��`��(�Q�H$�mV�֯:�ֱ�Zk;T�Z4�QTPU�q�V�v6�y�nFlm4A�ƹrӊ��:�nlD��U�㪮E���������6�� ��*���Ƣ.�*-f���4p�զ`������-8��-%DM�+��]q�QkX��p�#ZQN���Qh���E�(lS3X؈"" ��PZuQ�U%�QMb1͊�*Y�
f(����X�x�!*���"*&N�0D�Q��"J����`�&��AQT�5LU1MU��2DQQ31SLŬPUAQEEr�O ԔEQQUu�54ESQ-$PQE5SEM�IL�SQ!R��&&����j�*:�\�b����L\ښ*�b*��ĵ0T�514�S5DDA܍USUx�B���������a�+����Am�	R�"e�ƫ������6��d8�+��� �7w=��%t^��n���#��[Cn�/Tu���u���.b�rT&��EHS��A/ȇ��	��-ˢ�kn��:�΍�s�}�� �W�}�k�3ͫ�]ʴ݊�{��v���Cs��Bը��@1�e�~'�նj+��~������D�6��~�x�v��v&�~g�[�d؟�2}��A�����,�p��`��(��,��'�y��;yX����v���Agh������scjF�V;�7<��hEx���އ�{5�����ך2�~D9���Wܥ��l'�A���3ä���kz��t�]�;5;x/FmS�j|���	
��n9�(�A�e�@��qϕ�)��l��1'��+v~��
ݙ�ۘ3��v��sFu�n!�+[�q�A�%p�hH�0Y���V6�T���a���
��W���r�z��𨛐�1��S���t�('�� d�ͳ��>5eEÖ�+O��U���Ͷ_ז{3�������ps�e�]���Q���!s�D ���'V1*�	TXS ����43Q��6vR�¡[T�p�^�ޟH��(2�t�Nې���8��LZ��r{1�7�ӵ�sMr�I鷞��!;q��)GN0�zg���x<(��B��?O�qn?�Y�0󞐈]���9��<˳32�����������U�A���wf�:�u�]Qݙ��7��8�e_�]��q�����H/t�WWj��!IL��r�u�.�jyո��A�6��sUq�Z��a�������*;8 xtܚ����5������ӏ#g�i�����|�7����7���6yC�;�$��p[��>jw��@��/��o7��F3�	�=0�{�mѣW3���.ν#o��6�&���*Rz�6Ⱥ�1�͈���\�����=�y^���&��`?���ßypi�B^q�{iT�� �&^� .xk5	<�ܑچ�٣r���Y6�b��kf�>�Ƀ�cza�d����ɚ�D�qD�E�Z��Sa]k	�{���'�Qp�=��jm�_s�:�8���!��-0&5=#�[ݦ$��n�7�~.�����������j)&�{Q`��ƭ{�G��fr69�6'9�fM��Ø�2;Fj��79���um�hӠL;NW��<�˖��z/�0����xG�#���K2N���3w����|�śa�a@���D�1ǯzDg�hv}C�����$�bO�yT�~�����y���+p������{|�W���@̋!�!��4�F@v�t;?P�-3���%��n��{�W�a�{�/\>d.}Qx�׻�w�D<6�@��,��gͷn�}��A����h����]~��H���,XP%��l��6=�K�:��bPC+U����j�	:�9�VN�<T�	��0hɵ����n]ogZB�XǺ�D��Le;��J�Y�����%��zݽv�w��bWz�=����1�� #@�� �oS���+r��������������5�ѓ�{R��κ���)4m��F�1�.�2�o\��Y.�-���k�]�����׍�#�<?}�mCƀ�"[��#|��t�#yO��^��ǲ	���g<�dQ������f~���L����r0���^��u�/�α�t!2��%͂e0MP��w���}m���jkwd8��� ���fXz`eUqε�5�%�ƀ�zA钝c�IӁ/�L�%I��qO>��/z��]|�����].V6��шkw�n�.�)�%P�=�E�F�C�Yp�;u4�6	�5��٨E��W}�1��A��l`�΃��`&��4(��P�⮗�f-?5����#-�M�R�ݫ�u����[LXC��p���L6����ީآ��M�-GNо*L=��8o^(�Y�v�6�2zw\\�WC��Y�S�	�0��t<�~1���:��;�~1���Ʃ��W7Ŷz[+�T��+������>��]�v�s�@8+����.���&�0�Uv��Aa�z��k��"3r�~�8CY�;ow{[��`���޹C)��v�Z���ϒ� ������`�%�d2��io/TϖO��������O-�ÇG+���j76��
��ϸ�g&fڬ�ě
��I�3��+���(�`pQѢ�k{.�� ������ (�⒋��Lѯ���m��)����}��z����5�,Ľv8g����u�B.]��M?#���"���~3Cx*�}"�`�IHpsA1^�tE�noPgb����>�L�)1���b�{��q11�kObv3],�c>ݬ`�#L�����m�R����FFb���"vz�Xk��n���
`|`~05g�	����um�2�;$�;I���$�dD������ձ�� ^�H:�a�W�WN���b9��N�=NlMO�����4�W:+�~�Ƣ�=����:n���=r���1��t�S�`qm����]:#�X?m��Gw[ʘn/I���BSe�(2jњOr��
�=�Bޠ\H����(;��^��h���J���(��svA�y�?B	�q�d��3L�Q箘�{j����R��<B���틫��7�.�5�/tJvl���χcO�d�v��?y�Juat�eA%I����Z;YJ�d�u�T)e�k��\� �̛1��'Z�~�}	v?7;��O�b��~��u��jr;1�ۚN��g���}s�2���R�@��^9w^A����=���#9�B�^��� 8�����tO����y�3 �B$�U�J��yKa˗��&�g-c���Ư��������]�@��5.l�Ch�A}oV�Y�Ƅ�9um���� ��R��H�7��x3 =�z'g��F+U?D1��w!Y��,P&0�>}�l#�#�1�nc�w#�K��0�w=�Y�J��f��ctŧ匤����uf�p��C�!��4�^Ys��~t�`QGZ6w�k�`9n�s]���E�e��]y>;��b]�=ь� !���?s�cfؕ�QOc.����k<�^�NЬu~]�� ͵g�JNZ�6�~W>5?�e�v�;�]�_�?��g3���s�<Ãu:�]'��n}�R)r�L8�X�	��m�Q\�_�?�[u���ݽ�r��p���`��&M>����6�����Tׂ�)����0�8���L�kU&�[7%p�{us"�1�P/a!��qF�?���1��;�Px�T�)�ۍ�-[]�����掟�y�!�;��\���I�����|"a'W=8�nb�Ƣ�|l�.՚ݙ���LД�T[ˑ�i�ִ��O��`��yC���ב��%�˽ˡ����u5s�7Ǧ��� �۠ŉ�!�H�3�͜eY����s�{Y��
��(��w��S�	c&.#'4wl>ɔ��m�[��?˿dy)8`�U��H����)�K��kC�V������~r�X<\�r9_���������{�*�M�N�=�X��U�����1u� 5�������Տ�.�t|5��7�>�*"�����H�(�)B��P�D"� o^�o=����{��}_�#��f<�y�����ơ�O�u�Nm@�T�V?���;�A��X��a�g��}��h����9�e�#�4�k��\��+}b���
G���;*^ڠ���W=s}��v@�N6��:�\c<H�ހf��I�r�gd���	�}���aV�����u�B8���<�j�rU��:q���-�tczm��H8�rHۗn�ŵ�l /2q>����P�v�&A8LRn�I��@؃8^����@܁#}B~�/=-r��*�
޾�� [�8��ت}�RSՓ6Ⱥ�7b-#kǦ��;�?;�U7��Qwc�۴^W�|+]����5����|���$��L*��+��f�'�	IcA�`��ٸ N�	�'m�{**�2�1�i�Ӈ���,f#�7�=άWB͘��.�TXU��e6�����r([L)�����ﱅ����Lb��i��2 LhOH���4-XQ+\u��J粌ZuB:["2:Vf���;��,�B`��k!d"���w+,��Cܪ��=�>�G��|/���B¦|0�����1ƕڹ����,�q���x��ZO>�]�P`��t�a�Q9�u{}�d��<��̂o�^f:`Gy��{���wS�>{������kxdT������0Zvz���dS��.P��8Z�u�߿�{���u��=���"IE)V�Y�B�R�ZT
T!G�;Y���Qu��}B�mSZ�
�i�&��s�C�����.AV��7��H'COH�w�*�/53N�Άb��Qa���߉�v��-�tg/�~����wv���y�3�$V}Η�#��E���78���a�h<Wt�C֕!�f]�l����Tb�pքZ�����H4?j�O��S�Vln�3�`������B�ך����M��Vm�s�FyT9n��r�E3�~aV'sE�MF5td�[`Ԥ-{;ޔ(�������vm�k�ݴ;�G\=oN0�ʛ�6/H�2!64�)�T��q�4g.ǹR���X����o�~�~a�NWK�#��
O܊�=Q��4��)흡�q$>TòBnߙ��YH<ꭍޛ�������(Jee�S�),o��ߴw|-�GYh��ԉX������3�k;'�"wQ������hv�wL��=�f�'X��W�T�S�_8���N���y.��t���sB1Y�jvC��6LG0E�K��>�%Wey�.�Z5(���U�ӷg�x�G&g��&,C�Ƈ�/h�)b���پ��S��͈@[�xv���Ȝ���9�=�Fl�b�a�ׄ�u�k����	P4,J$���a-���N�+�++����E�F��#wPa<>�y�޳��cn���X��ͪ�ɼ(Eu�c��~��Ā	���
��3 ���<�� =�ף	�(Vj�yo��cÇ��DC64�[�`&��4(��'��]/e�?5vp��d�%��KEI�V܁S��8��g�#� 0t�����^��.��`X���aD��
׻m7��\��m�n�F��ͅt;����<���|�߸�~/�\�ê�r�y�>,xT�ȷr-LP�N�xZ���S��.����ܳmt�m�u{�0n��r]g;NGP�]}�c�-�f���f�Y�I������>�z�0�k�b^�;3箱�7R�n��_q�� �?[�y/�����`3o\.}>��C��LW����e-�r����gM��81�<i���X�B
P�/?gx�͌�K=�s���ci`��v�s��:�����S�i�{�����P�X�Lx?�?^�Z��ʧ;�~��C�׶���3�����"1��Y�ϗ�~�P�C�<�R�_ˋ�ΖV�?�͂22��S���r�ұu)�e�3Q��m��
�m���*���	�$r��ŧ�z��^����-�â����5?I���߬���`�V^����o�]�������b�z��o�@�)��^���Mop�8��[��P�Y
��r����}CQ�tY�h�������)�����b���OI��Ģ�>�w���ٮN˾N{`���0s�yD�k�'��{�﮽o<G���
�
ҊP��� ��J�:��j���ϩϦ�u�pI��d��z��ƪ�wF���Mh#(2j�f�ؔqW�G��tq�7�R%�l�V<Tm�Sx�n�hR�K�"A�[ ��U�OЅy@�1,��L�+�i5�Gc�t6���T��~g;�T_yjLA� ħfʘ,c@#��?D�I��K�B��E2t��䦉lN]أ��wisq��M4��L���&>d�_s'p����#�L8�)>F;�J�PM�������p���9+��++�h��U���vC��׃����rq�=�T/�1�
*�E����k�e��L����y��^���İ<���8��80�G4à\1��پ�Ÿ���*i�@e\�wj�jY�W�H�P�?s�|Hw�H���%�?|9������:�+���K�HW����v�'VH�5�&����I�X[�M��W>�j��+b�ٶi�=�]���R��k���D!Aμòt^�T7>׻MV�S�1��잜��@<�.,�<��%�e�J�y:ܹd��wjY�y_�1j��������v��v�I��Fi����&��:c�_��Wq<.l���+U��[�H��lo������hN2~�$�ҝ����w"��b�1���o*��>�Ҵ����Sz�d�X��,R���7_\��L#���7�ݮ;D��~8q��"�'����g˵wo��<����������@&
F��T@��ff��.�Gq|�[��/<߃ˆ/�|�OC�>~�����mH�J����vM����J�:f�tL�-��!�5��L���9�I�_�)���"L|e���/���77�B���<_v�����\�����4��Iv�8�5r2�m�I�m��ȧx	��	s�^�1�kM��0�!�^&�ӹ��CP92jJ}��XHγ�E��dw���ڎ�]\Nsr��3U;�B�s��
y�}�l,Ed��r+�t�Z�;'�Z�,�.�g�zCW�����(����e��p��*.W�3��]���0LO;H�:ɫѐ��e�d�'Y���DD<�=�ޘMs�r��_��"��J�"�}�0��v�ְ�?���M�����w3�g��Ϗ�)�.z�6\s����B�'�n)c�����2)T��~�a�vE�*�����H8�rSe)��+����_��-i�o����9�{�}I�0a�E��XH�b�z�[�	��!�&�-�w;o9z��7���"\���<��˰�6�ʒ���5���x1��#iz'�C�3��|�^�/G����������w�����z<|}~�_��\���Eޘ�Ma�"wD;�is�Y�v9J�oYK,��"H������r����}��q9,3�v�5�J�q�z1w8u���U"��(���nzֻK��d�K�]g�j�4���ï'
�5��M%�h�=��ҫ��]F�t��#]3};m�Kx��6�Ÿ&���_:�v�q��}����\��h1�݋y��O=�3��ޞ~A�ڷj~�0�Q3�c�KᓳO��2:yZ�23�8��5b�Y��Y�3��=W�o�ܭt��E�a�i5U\ ����>��öE�n⽾؛p�ә�dCy��q�+cR�slZ����U��ra�g�V�A����se����H��^*b�;��SC���N�b��|�+}׆��1s�(��9��{ƝQ�Y�('��۫�����Ԡ�`����8��u�W�&��J��F�,�˕�-�]��CL�2��i�?{�{?Q���di�R��8��k���'�޵]x�<:�Q=��=[���q͏���{�"kME�J�V#�=ۛed.��d�;9�Pv����ΆMGW��:馴�(s���:��d�n��8^��0��۱��a�u�fhi�?
��I&:Kz��[�Ss�9{���2 wk�oY��E�*�:fJ*j���Ј>R_`��U].ėk���xm5#�W8x��y�1n�IZS�G�����˾ynm�fa�7��u
��K�=+���:	M��X�܋
�L9�f�f
!q��l�w�mѧ�X3��ڝuC�;?X9�i��y�Ɩ�ɕ��2֕��:<7̻���Q	�9)�\ڭ�Kڭ���2���op�f����V��<���zjx@k�F�آu�$,�y��s4�6�6��#���v��5b.eT��q[/a���\�x�f���w�wԬ��_oK�ƬdDnΗ{͉G�;�%��JH&`�漜7�`���^Ž�DY���VT����r+:�����mЧ��;׳��LD4`�VgE2�kYFm�[W�Қ7�\�(`�2LӼ:��x�����u�cr+�(2�ybP��l��9�E��"�hf���R��ڵ
����� ]'f�p���6+cH=%?ܸڦ/s6��Z�wɪŝgk�����ۃ킣�;��'��L�f�|0�$���=��{\X��җ�ɤ` OU�-&k�ڄѷ��w�Ŵ�#��|^�ǀ�6�S�YT2&f[솱����r�k[4���B2fyڷl9U쏇�Xu6�a3���.�˿���sC�0t5���o��ZL�i�^��{2?1��(�fp����T�����rHC���躶�����V���������9yE�y�3V��\���ٛr�uք�Q�-˵�޲��^cǮU�A�2�;���O�^�|xe��o��w��j��{����z W�ۛ��mW3O�M���@$�_� �E�BEESQMQAT�G\3ITUJA2E5�E�UEErs4E4ED:�{T����Q�"bh�
H�*��Y�61D�%1M4��1���h�B#N$����Be��"&j���i�)����j"j��"��	AQ<Ϊ(���$�������*����&�*J���b���`�M:i�f�*�I�����F"""����)�����h��b��(���!"��� �(�����&���"CN(���$�����b�j�����i���"�����I��IM�F�j��� �*�*��:�&���	�"��)����*H$��*"�:�*&$��"��c��SUo� B?���>�䲇��+jtML엣rbD�͇*�rkK�n�kxۢ�c8���v����Q�sK��o��e����~��@��� ,��2B� L""���}��f����<Ð�^�{�F���L*��\��,ܤ�iIcH�CV�W�v��1n����f��%ĩ|�,7;��_'�����г`ĝqvJ���e3��*�c�'�2�u5wj\�[l,:i��
�-=Z{�ʠ����������J��7g8�F�JN�x6ݶ�?k�ze�Q�Ѝl���0��g��j����T�-)��~[7!�jnn��;�8%�2�PAtN>�i�e�;�c<���z~�&8y�Ƈ�Pl�Dx�P�Vm�C�O���2s˷Y:�w(���]��f8��f]���8:���yw��gnUz��2�]cTS��"���S��)��EF6��a��C�wH$=� ��˱���,>m�1V�R��i���e���!'�z������آ� ���B�U�V�=�W{UW3s��q%��y����~�f�;kܣ=��Xd�=TI|��j뜩ljԤ-z��W�g#�"'Uv��f��v���P��q�Y�~��a"�*׶)�M����~v�1N2@8�=$���������xvv������X�͖ �Xp�x�R@@7�7����\��>ι�l	�e����]���Y���|�']��T>���f$�r��SU��[�`�⺫zZ"0f>�.��Ԩⶒ|&<�"2DuA��yZ�9��v߻6���?RE�"F���$A���Z@b@�f��7��Y���n�[��-���BSe��&T-*���r�ߏN��H��Ol���f|��Y�?w*oū�������8����{�H�3�O�Je~/�%�b"�]���z_q�=�;Ȩ|.�Z
�|Q��.��4a�����E��0�ƀD��ק�e'X�%�u��L��*L(?E�T�u��MVɪu���g;��'Ɓ �6;�����D��#�(�ahԢ���F�s��]�;�֪�)#~��-4̆"��$}	F~|ǨL��dI��*��].�_`g@�@Q�)�oouY��{�5��*�a��~��}�-�?��_0>OPey}~�dx��s<����|2��=zu� �[ʔ=��u6��s�qͥ��ǆ��k�Ř��u�LN�)ƣt�0dMVf��F�ƭ@mV����+�t�{������U2s�;!w0A��9�3H7�[	1�ݍ��b�u���̱�p��r�o��O�y�ύ�a3�׭3<��1a��X݋z�6�m�C�;fDt��{&*_��2~���=���g���D������p�*1�1��ض���{f��K�Պ�)��ŪՅp��W����ǻ=Vצ��p�:�A8���)�{�E��<b�S��غn���b�]]fO{S[�������i>t�5�����>��@�\��ωs��aٖ��D����ΰG�� � 
�(ReF�	` ���"D�h�B �P�#��s>8<W��~����[���<n�F����O�!�Y� s�~M�g��0T�z��k>~�x��N*��70{�ո��˳�ཫi�y�[�]�XȖt�52;[$�'����H��F^��;R��`�d6w>�qf��,5 �P�P戮
��ˋ���;�3����X�1�5Έf��̭�����8񜽸�����6w�l�ʭN0MI���8�i�/�&�#�if�wV=X�^OނDB:�Eǧ�eV0]bv+��BkЌ�ɪњOŰ��Ƕ�x/�+P�T�8�rͮ���k������d^�U�OЂq��~	�W�F�^�0Bq�3���~�]�רw���4W/�+m�<�O��f�=Wi�Xm ����z~�N��bS����<�Jֶ׃ot�ul���BV������j|��5��٭�Д�l?X��>�,Z�.���+ɩE��淮Q�O�I�S�c�bc�p��G�e�[w����Bc�E-��DC*��гoy�o�3L6�q3 �&�z���R	u��w ���[
���e�Џ� _�?7�sx�I�<$�F��d��\	V`��d�E��Si�U��Ex�r���;�
4zj�Md����.����ְ�O#���8�ߐ��TޜjS7��#���YK0S��nեZo"Pe��Òu�Z�v˽�7|����Ü��V�����?��J �J �
U"AJB%�Q�B�d�
>z��_�Y˅8�xk/��ɦ=�u���/5jF��)�����IDô��g`�I�E9�эy�ٹσH������Ҏ�<��	bA�X�g�'-kL�z�s�S�i��4�q���6�M^��ٹT0l�$pt�a�]�OC���Bը�Á}d���|� �O��wVٻ[�g���K��C?L���
B����R���g�O�:��v�.Qw0!�!�dU*8��۲�0�2��j�~���#������}>)���6����#ύ�s�,tJ3o�8��]�hA1%�I�b��9!?{C�*�-?k+� ΋\{��gL�u>�~�_e����*zq�߳����R͵�@%ڀ*q�j�#.�o�i�����zۗ�8:�|Ze�B"5�=Ų繫�un��U�H8X�2n�Y(5��>l[.���:Ff�(�}��8���n��N���`��>�ǆ"nB79�^�'ְ�	�8�Q��7R�Ɂ�1��4�T�vږu�c��*.��6��?`r�Ɵ#�<?ܩs���~���Xߚ.��K�?��$]��A�9-��IÀ�w�I̼��#Q�TfY�s![}�S,����[�ç s`��,���1��Tэ�`~bw����w���-C��=6-_GR����6���s�;LNg�nr���V�괿_>|��{�:�}E��(�
,J)(1*��_=x����g{���;���z�(R�K-�������9oR�,���nK�r��V\�GGcP���~�0�͎X�N�S�	�U$�ߢ�g�"�F7���i!^�Vfm#l���^�9���S#��&X�b���)=$Mpg�>���p�p�O�ͳu8�y׻M�3�`6���9��A<�@��&��vT��~&m�t�n�H� ��:%C:/2Yu�|���ڣ1c9u���8@%�C���	�I�'�S	^�+�����o�),r>���Uw��ޔY��F�(`Y�٫]��5�0t��q|���FjE ĝqw�UR(=0�bʾ�|���E��n����ف�,A1�~b��B�����:;^��傫f��w5���e7,Gu�qCtT������\��z#���69��r�(U#UR���31��a�Wes�;R�m�Mk�wh�#��1�U�`�Oއ�1��*�1��\�Ϡ��͜Y��\�<Ec�L3$�v���1%ڀ&Z��ܘ�c���l�w�?G�}��ԟVlS,�+25��<���$���Q}��룜j�u{үpH�M\oٗњ�qjfVR����4��T���$S�C���I�M�U\��n�����kG���6�ua,5,����D�-fmY"�]�S��KǼo=o{�^�^�ux޼�e ���J�$H#2�J�CKJ^��~��b
�����^a�>0�6nq���L�3"�x����TG.�c�E��M���L�1��;AC�oh!�4>B18|���騼{m���fA!�vA͌�iih��)�++�[Ԇ�;>eq��t�Ú� ��Xt�����%<5�2���U����`�M�w:L ƭe
VTu��E���^������8p5�mȭ����}�`���'M��m�&��WB�	��ZT)=�9B���cռ4��; ^�f�ătX���Υ¶2���{^A�sk��_�ħV�X&��~��ǯk�<'m%�7h��ʤ�f�gz�L<��C�8#�ƃ�a#�פwL���I���z	*L�kN��s��oO����9M�Ӈ�>d�o�>�ρ��H��&}�]0�jQu��v+/q�vM���Oѻ�Tڼ�i�W�r��Z�AQ`|>d��������� �(qYҵ��>�8c�s�7Ԍ�;���,J�0�ԜK����uy���~���٢���q�ݕ8)F��WR�8�z�u���~~�y)��u��O
Ul��q@�y��ͯG��U���-c���I.�(�5ޏ���d��=_��'So`����a�j��N��/~[q�b�M���7�zn7�T=w"~g�5���>��c睳;'Y���C�>(J@(Fd�7}|�׭M��Ns���v��P��W3��|�3��<y��Ԩ�ը�u6��s���<^�<n@qFϜu~�0��.�]�f�L�o]��YN޸ɖ��<��)U�9t-r���]q�}w	������kݹ�`��7�Uu�=�A�?S�6�e�ۏ@n�&�'̣����>�rb9��K1��ś��);{x>�0Q���W��c�����v?Pݐͳ�(�A�$@;t$f�\��6��Xwѿ�4ӯ�p�]=~�����a�����f�X�hnְvN[#҈��������վ��1��R3�E�ڔk�2�|�02H��I�z/����=�Oe���g�=qn��!l�aT�#X�Aܤ�����U�ZgK*����>?�����u�ԩ�Y�'if?)���9m��a]��z3aUjp	�$c(Flb|ǫxU�)�޲}fa��R���c������\����Uc�w=7��!6p�(2j��4��a���t�	�pBY{2�ۋ���C�>����@���1 ��dQ����N+�bY'HĲ8����c�������w��%���N�qc���ᬞ������-^��{o�q�EW�j����������:�M�᧬�[陠p�ٴ�<�Sy��2�3U,uh�Г��j�wl���F�;�yx�2E1x�,4{�J������
�U�>�?RA(@)P\�����λ����_6ַ}�3��X�t�On��!@��D�fʘL����"�l�v��=(�5I��Lw\\�� m�7����)ĥ)��Gd�6=C�p#5�fֿBR�ja3�fYy�����u޵l�{��/Ϝ����!�J�v�� �%�X��Ú�1��ϑ��=����r!6�64(9Kt��j�دd��S �&�zb���R	z���Fi�������Վ��c���ًx�<X���m@�yd�GVM6�j�k�vQy�R5�= Tw:lw�1.��Μ�	ߺj�[�v,g`����b�!��;'�S�+�ɯ31�&����I�XZd�ի�o�Fd����6¦���8�?�~�i�Y�1�]����OC���B�xL;��5��hP�e�"����ި˕��/u����_�8��us��2
�ĉ�F ֜���hv��6����G�u�t�;���9Ŧ�4�%怳�QE�9���#���#��0(-#��&V9�p�D��2 ��5³P�µPd��4"��ba���t=�W�R�{I��A��G�[7{��}D���ɥc�^�����t4�#��i>�!c��,x�ޜ�L0p�ՉmL��v*�ȱj��U����R�:�^7�g�=ajYFi�u �k&�x!���&\�~<!�6�{k�1��b����l_m=����J}�jyv��� � }B��P	���Iv������1\�6-���ǻ2�3Ei�]���:Q�e�}kס�6�fy�t�h�vhǶԲV�D��-��R*��i���=�\����kW�AA�x� ɫ�d�ԑ�g�Ν���-�9��ݽ����}�ŕ�RO��c0/|�5���\�nr+�A	���a������G%1
����;�sv�`����r�3 �]^3	��o����S̙��:\26&Y�Uz�|�w\4�R�j�{�|��)�D�L-��8�:���\c<zD�(2�t&v�zz���aVт�/�3��3S��u�Ps	�{��#"��I8�ӌ;�Ӎ�Dc4@L�W�+e�[��h8@C�c;r큧s�{�Re�c1C�J}H�����[��͹���ܬZ�SB�V5�\8C�@���Иs��,���7d�OD�2�:;@�^ԚGB挷]r�(��UU�^͜&m�"�++����pC�P5�=ʄ����4�j6�L(�"��jy7W���,���L�ݾ��}�ȞM"X�k�co��h�	��=ά�гf$닿�~��TM:y(����c���S>��΍<�-�U.c�Բ"�^�V�߱rwM����;p���\�}q����LQe��;�R����,��8�L�W�Zû�=�2��ƪ���-D��rdB_)A����76ֿ��i�}�҇ܭ�&�0��'�q3�C��x{��ޮ����m[_R,><e1�WZ�+���g�(5
�B�(y|}rĥ�q��.,=��d�Ɏ�z���0��wqR�:�[.��NK�Q�$,��x�K�s. Q�����y�����pn�/fߣ�2�r���Q�L9�J��˦��;NW��nj=֖��Щ��g�2�UO�m����!�A��~��?r�u���8��F��z&o�GDc�����rf�y�%����2�}J$�cpy�5>XE~�s���f�C����X{bZaŝ�hZ�on��!Ou�e��"��؛xn����	�"ˉ�)<K�=6��h�d�c��;Pur��������.�l(���[�_��s�
����8�sE�MF5v��v���Ζ�7a���-l���kaU�k(R��뇭�@.:kծ���?`���E�bZ�/Kr��B%�xfη��nj�3�d�`�	�iP���ȭ=;��z���e�_�}�N:>7�+F��{�GHz�L��W�i�O3r��/�%�c�q��� C�������{|��>�w����{}�>�w�������O�����i���-P������!���2�Mt&͝��>�7G��b�n�n��,�ެLv,���W��2��0�A���t�c�)��%# �yH�ٗf�.�j��`u�.Tz�ea�e�����ݽ��������!��w�� �4��=ѩ{�@��ZG����[�p�t��7)|�_��+�N�,D��<�b|��m�>^0^xs���8�ʝ"s��QMj��zX�W�{\w��+�br�0pY�o���5U�X�ܽ�TAU�����������j
.��Գ�#�N��q�d;��h�R���\��@Etz]����mOm#����F{OڠSE����؆0RĜ֞�df9��p"U��Ϳ���yu5�j��w�F��I�^�Y��C��z��#Q;4-M�w��b0��P���uon{����:'�!�X2_|����U�i}S�,�yyy�Ӿ���ȶ47`a���ZL��hޭ�5���1� �z���*�9.����:���gzL��uٽYΎ�[����Z�3��-���Tp��t��J}�f6�S�9�G���^Ů��| ��M`y�ٵX�	��[��!5^�`�{.�D?����q[k��I�Y�+�Z�z��s���+��|I�>�2vv���5P���c������pWC�����|^���
2!*�srr2͇h`u"gi���q�����$���X�<E���Rz2���0~$�����Jv�y]��6��,��%�T�3��p����N���΄�H!��l�'��}����.�Ʀ��U}ui�۷���__|8�ו��o�^���Dꮭ�n���n�獌�*lj�e��\{ɬ䱄c�?X/h�{a��M�G;}+��z����"���Ȗ�3<�
7��jX��9w[
"a(U��`��y��>�.>��}K�q�8c޾ń�'6��,>�F<���2�I��g�Ģ�Tyv�1o��Ѩ&�Mv�֯r-֠F���*^���2�����ِ�vYN�Q�ao��r�e���L��؈V���^�s�����{��ŋ���u�b���͙Ωl���L#V7�vu�ʦ%bȄ�"������L��*(.�˥+�Y��쳼OpM��M����k��t���m��ԗlm"t�ٺ[��b��{�Y��m��ō��8�sބ��z�|˂᜖ht��}����������''��	u�#L[u���p�lf��gC~<۲�evʹM��v�Kb�`��6��&�^J]�5}sf�	�<�l=0���٨��w)ݎ3�M`ѯ�ܥ2XQscf�Qt��k[��E\հ^H��R����Vp�Aw��e&����U-��;�u�N�����QS&s�HB¥��b>"�����kꏫ_@�U��ٺ��=u��μW<QC}lG��**��H���gEQQ-IS_-TE4đ1�SE4�5�5TLQ,T�b$�J��*"��(�j
������*"*���
jB�""j��"i�� ��(���(*������QE5T0�P�E5APG �UCM4�AASETQQAUEIIAACPE4rqQIQ$UAE�O6f����h�(�*�(h���������j�J)��&*��	��T��<sEI6�ST���RD�-UMUQAILBA5ACT55EQET0T�UEQ11�b�����"�*")�lSEPAI1T�L4QD�ͦ�j �"��(!��4U4PT@TMD�������"��
j�J�(�)��A�"
��(�J������i"f���z���yގ���w:�Z����"���mЛ��SM��������D�+zۺ���7�;!�0� �5��7q�J<eU�1��uɒA?�P����N3#���� ������CC(�q���br��)Ϳi��r�攭�ӕV)|�t��>^J$8��r��	�B~�pF{�׻�t�"�7E2�w���Z�ު�Bֹ|�:�jw)s�ȼp�Q	�k�@3d���vz.���,H�]�a�(�`�MKP��7��u�0�m���E7b2��`Ӗ�p���B
��GM�&n�2$�|̪���&�l�Y|��j�s��ٓ.�E�洠�]�0�r;`>��y�kP��ʧd�Wt:&s��ѻ��p��WT�պ���F�Gs��t;��@����n@qF��)ټ�22���Z[��2)y8{���LV:�5���V��r��.|�Pq�^��;<�.�:-���Q��[��1�؃@����u�vN�FL3n=nt�+�I�����������>΢����z��ag����6����#W�0���򁩫<��־][��;%�/���-[*� TM]��rn�b����(K0^DN2k6!�I�w�pr�4>J�/`N�k���j�C�J�#"�d�v��R��z���	��`��k��鮬p��~0�1x�j�'>a�*�S�v�K�fd�α��3e��i�癛t_�S��.���ï9ּ�&H�hMȶ��f3A�'��7����v�> a8�Z�$"�w���	g�C���eg�;r��ڗYSdr�bM��N!�����-�u�t;����������|�2��C������}? Um�2���%�����|�R�_ʹKL����l.,��<����*��V�L���¢���S��[�a߽�'BP�8�5�R�E���z�=[�&03�g��Uqb�jk��\3P����4?�����	F<�����h��҉O�J3�.��a��q1u��aΥ�cռ'���>��l�DK�:{�@���1}	Ǝ1,��6�wA�׳�i���g�{��W���VpVW�
V���bx.͐��;A;$�'�Bl�I�s��;%GF�s���S�]"�PIRkk}��,v��9�_����a����#�;������K�:^��,�;���dx�w���A�$���PT�H�Kh��Laz����B=�M�Y<�*�����-7=��KrO�$�'�uL1�M���-?,e ^�����a>=�o��fv
��z�WŴ'a�צB�q#f%�?Mķh�����/�k(~�[��z	��r�.{6V1��:���VK��w�������;��;�|�O��W?�7�Sh��Dt��i�oU�"�'���+�ɠ���q���Vw�-�N��"����1(NWb�u͎�;��`L&s�x�L��2�ꋳ��85�j�0��.��cp�9�K�I��jH��vY�Z��~��Þ��[�e���W���n��A��H˦kc#��ҫ~��� ������{~���5|2-ݛg�����6�/�OC��i��2O	��`���>Z�W��V1�@�V٪���:�G�kB⟃��ƴ��~}'�DdT+�yzVˇs^�{��D�N;���i�D�	��-�ܶ���s�<h�gh��� e�M�@��#��d�wJ�r�T�dlwPns�dF�3Eځ2�Zw�$=�W�~�-?V��V��A�}����������Zb`�랜m�Y���e�f�0y��!��;+|kO��32\��n�����8��-���E;�e��[�&�}]~ݭi� ��Ŋ�!�ԹթZ�Tg���~��Rϻ�d+�r������`_|�Y����\��u�Z�����A����Ƀ���w�\����*��?ʱ�k�l�1pBby�Tk&��NGDG=�s���n���m�u�kި���*�Ja��0��������@� �/�?H��.�jdz�Ez�K��힍���eۄ��SsP�Y'�9�N���ҩ'~����C�����զ<`6���7Ua_��݃���Z��f���XTؖs~4�6r�}�G]M5�_^B�MpÄR�gC����Z%vY���::��@Y9�<R��{��>}tCv�ܜ����T�wv6c�k�K��A�L�\�sݏ��/���b=����m�n�u�����A�P�A�v�؆�nt�wJ�˘�LP��BD�7�3�R�����w�oՃ��I�;�����B��F3�	�϶��5-C����=6Ⱥ�09���9D�l��T�J5"�l���\�T\W%�0�������7s�XCB��uN�a=㒹��qّ���ƶ3(���y@��5�v�|�D�ƱD�~=a���*��J�]0��hg�gO�8ue ���-š��7���e$+�a>/w1��sۇ��7��ߎ�8ǟ����'	>:~������*7H�՝�,�1+\u�˥s�PK�)~a���+��=�~��?�5��{=��f���ܪM
H]�_�~�u���-��,9��T]��ݢ��X��0��͗���O*aE�Sxv ��:����V��2�ǝ�u}���rK�9�k��	�*������*���QE�z�;*z������χ<��
�|/�S�
�8��u3�e�LC�fZ3}�1���jT���}��CV˴������L�CX%bO��,�k�y>�8��=�� �8����L&-M��b���"��`�]:��[ׯ��0I˦[ƴM�B���0�V��h�Ӷ����"�c�J^mmZ�*�=��j�Y��o��1�y�F�=��_���S�f������̶jJ��24���a�T��i�7[k����Р�F�p�y��1���[�n8��B9�H��t�P�=�L�����������Ty��%��7�!��6{uQ�ml*�8�1oQ�RTu�׆��	��SؖxBmf��:�to�^_.n���8�v���]bv����Jl&dm*��$V�Ӻ�=[�k�Q�f=z�
�/�]��X���na	�=0��;�P�Jce�S�JK�"�Z `J�1<��)���m)���xb)��
g.H{����ێ���ݙ%�/X��F�1��{�\�On�mCV�aO�|ᮢ�ե��NF�#�U�����ey��qW&z�ԝm��7nX!�R�xc��ԏ�^��$����2p�σ��B�n��f�nx�h�{6gE���r;��0��B����-9d\�+���W��w���XG�:mb�sI���f�jJ1�B��'f�Վ���;BB�w:���p;��@�^�<�9T]��v����m�OasL:=Ô�f�z����ҝa<�V��^��\sHWrͱ�APiQ��LQ�O����t�=�_��X�ऌ{=��؈�Ob�W?�����We�m�1b�Nͫ�w��:��m�K��)vܿ���e.�e�����T�A�ȬбF����w���;M�v�� Ʃżv��:�)W�ͧ|{�]��������q��F�����T���x�	;�k���f�z�6�Ĳ����>�u9YŮ��]�	lW,�;�Qeݒ�K�ge���&4?��z��?	�|�u�w@�yw2��x��2�q�#79��;�r;k�W��D[�u�v2:%�,46��ƽ�A�5ܣN%��\c9���,��$?x�pG�b_E���P�C"Y��A�=5y	��*r*�S���9�E�^����#w3EvI`k�e9Aw
��ˇ)i��T+�>�q<(r��~����~0#��s铎vn}��k1V�J��� ʔ[���{Ȳ�ٵ�͚Y�����/oʥ��H�x���,:瘸��U��;��Jl���ɨFW�h�~+����RP����nUt�B>�<�_�U�ʅ�I�<�A��.Ǽղ�F*��A8Ӷ݃�6L��R-��Ơ^{{��.���ebQ��b#��ܬ��J�c>OȜ��#�a��w�xU�a4,��=�-����1�}�N��u�Z�ʒT������=�'%��~Ly�f�Bu~C���\Z�T�P}+5�Y:�K�f��T:1�\�Z���!1��W\9�����gOX4�x_)[Bc�ƺ�Q2����Ǐb��T�P�R]\�g/u-�a�{�q�
[�A�n _����{G�/��2F���b�	/��8d�����:�����,û!C��i'�9�NV7H�Am�Laz|�>�h��[tLm���ۯ����baS�%���Sq�t�/I���ҤuJ5l0���˪ӎ��'\�e��a�d00Y�q{1,���Y4�}���"�E���Q��.�[3C��$UL�ͨ�j�q�D�/��(��}]�4~]_�:�r����2k�BO�oZ��g�=�J��|���qȗ��s��l��n��#a�:�n �_Q���4�Υ|z���� Ij�`�|a��!2׿���3͠���������
и����|QӞW���y��o����;�޳KK�nH~Gi'�����^�~娽�q�C�h�Xh~ò�Z�{�K�����Y�����̕�PnypЊf��0�[x�:hw�_�KO���.'�0߷���P�tq:1�&s�N{�}�i��7�Iv��q�j�e�;$��j�1���C�ً�snzo�_�I���-(4T	!���^&����kbt��o�<w��;��1�Q�.2�XDY`s����sQ7T)\�WL���7d!�9i��X�>�xgt�e��:��6�E򺇬��K�ˀ�~��n�*��هFvv0/C==8xǄ��ͼ$�"�0%���ܤYa�&�D�4�ޑ�|�X�E6�.�7�#Poo���){]��ه�1�+�r���1�`|��N\��u�ߥ��������{�Ԥ��r9踆$�� ��|jʋ�5l���.a�!�s�#���m���NFo)&�u¦�S&x��B��yN�%B�)L%�.���z�Y�g�[�t�P�o�%j�Й�5�.�^����	�{bS���"���ӌ$vE��S7vG?=ș�61Mg��pׅ� ���v�<����|~�	����-����:F�`ܬA\�F�=�mY֦]}���8 ��:	���#�}�YWa�i�)蘦E������4���;57�[��'u��i	tO-	q\�
���O�x�QO�t2$���y�m��¤�WFgk%X���� \�y����#�'��ݚ ܇ǘ��L7L@M��z+�w�\��'���o�"y{�w\]����]<�o��XO��֚��j�����m}�?ON�]�ط�e���ءڼ�dZ�Z�?J�)�ze/����A߳�0�8���4�����#�)Tj�;�]�U(6���t���y�����-�X����x�������v]�H�"���]��nR��_��V�k���D��Z�a�g����7D9�&�pʡ���3���ɋL�*���$��gF�-����ר��Qza�?g��ʆ��Nny~�&�p-����,r��-�5�,�k��jR�m�Mk�wh�fX��0�F�b�^5i�;�|�@]
I���hP�7���>�}c�����@�f8���jc�&�ij���i�v����aud�x�A�^%�>0}��G�u3ǲ�{�tik4�����i���q2� �e]ok`3>�A��cvR{��Ƕz�𴸞c�i
��Q���|��Ȥ�A���:3�ۍ�M���tS<��!�{��.�r���>ڿ���L�T�6��:U��J���z-�C�;��ٖ�Ca>ݙ�;*w�#t,le�a4�Bv�S�Tl�soA�,�	�J�'�G(]�Ӻ�*���SM&k__t6q�xeϬ��E���!�C�|Cwb�j�Jce�S��RX&�ѯ�,ku�=�i�N�����?�-�tqD��w��'T(L��hv�{�e'Q��hQ�Sa��9�[�R�Ϩ2�c@�I�s�8i�4B}���c�`��t���dQ%G�{)9���,ڼ����A�v�Wt�it�|5��WT�YWanĘ�^�)�B�J�����׫�y�mh��~��U���NT�|�A\w:��=a7{���ݙ[�+��}�v
����W�n��kY�����i�����۳��ڕc���;��nE-�&�l���ʆ#N�@��-A�6��A;66�	����j�ɝ�޽��!��B���(➗�1i�������2��8�s���9wJ���Yr�kJ�x�f`̱����seN�'W�SlP:v�߸�0���Ԫ���� s�qn��vw�f'݃����-������f�M��-l�J�a\�W9NKԺ��T�Ӽ�!�]��L���6.�`�>��G@t��;k���f�z�6��e�&6�:�p���k\����d-��^�3�KrY�����$������=�MY�sZ�un�N＾��{��<�E���2D�nk�
y�x���"�&+��}�q��u�v<��^A���^�I���9\s:'����~r�������$=D'�S�m����~ǆ{�BKv���0.V���{Iem��^���ui��L�@vI`J�1?g�9�~:!�7R�~5<��L���V��j�tD&����i����5>�zܙơ�*fӰ�#jq�j	�� �w��ޟ�{}�G����|��������o������*�\Gz�t�rʔ$�v�M�z�
�1���`��]RִKߴ2�]��f�6��W+e��k�^N1�Ύ���S�9#=��=Ɖ˜�]�s�hD�Z�a����n
����"��ZX�_��v�ΰ��N�p�ı$n����P���GL�DK6b�#՗�MQ2�^n�p����_2���{R���?NW 8g�Ky X��7|�|�,
oT����2T�К늟����ɱ���[�)r�f\@ظ&{)�1ҪL������ԗ6��N�:�.�;ܲ�X۳���G�G9���Tsl�T�L׾~s<�6��`��WU��=7bT�؛Ǻ�ɱg6�˨ND�}h�dC�4��X�V�odm����OK]�i9��y��cGw�<n	Y�N�E[iG���x�=��\��"K3G�c�����8��)���p_uӗy��~���L�q>���m�|��lJ���<FUq�`�	4�gKݕP7i�H�w�50`�/��nh^�����ݾ�gi_-�;��K��{0�UWM�u�S�����Ym䅎����K���U�n;9k��y�s"���R@]��3��@g��!�ï�T�Lˉ̚�H�}���d��R=�+�]݃��+�9��û�F��o�������͵��&���q��}�a3kf��ݽ45�����G<7 �9)���t��7��o��s]d��9��; ��w�*7e�a>��Y�ǑQꏁ��L�E8���|�o?+(RS*�yθ!Cg� �'�G��r�Q��W����eq�e�z�����]w�X�#g=r����}�.��.<U ����!�t�&���VL��x���ŕc��䇌 M��[rA��D3�O�O[B9�|�X@���r)]>�>�(�ڂ�|]�rӪ]``�OV�r�n�5k���_�R�P�W4�LW[��]$l�;���5F�:ߛ�v� [�RV�b�6v�<x K���=�7�{�w{xK+�ꀒL$|�]Hq��7�+)�Q��Y�Mc��F��Epda�Z*a�_+�;�}�o��qI3���ޟn`�{rY�݄)0����w! ͭJ}��'�{P���Jy,�ui�S�}��|Q�x�y�#V-��š��tرt07�{�X۱W�^r���p�Y_�SР���0Qz��ev��a��p1�y��:�__;�v�g,��Z7�:����i��Zz�\�gZ���"2h�ֲ��z��k�fc��rנ�H�;ܲo)åG�F�9{��(������1�x�1��n�ɹ[�==�.8;[��&����z���c���fѢ�XդřU�6<g�Nۏ�����7�I�j�n�����{
;�ut�ڥo�l�J�5W,���cN���\7c�eL*�rf����mِ��b��Q�)���\k5M��yrN��ngf)�t�F�QM7��j/13M4T^1��((������
�h�d""R!����(���bh*!��馢j)�&)ѤbJ(&��)� �i�h��14��QQC0ELZ4S'6��P�DKCK�b ����Z�j�(��*&�64�LkTQN�]Z�"&���	(�j�fI��m�6�J���f&��"	�`��(���"��!��������j�c5O1���(m��CQPRD��ZDES�F΂���"Jh��h")�
v5I4U)Cu�E3UD��kZB���j���
"mU&�J���+l�E�uTU�%P�PV�
�"S�:t%$HR	������?_JL)�H,��M������Vt�|��#��,��wn)KKv��Dy��	��g�	`����W�;�?��[��Х�韮�w���0i008���S�q��3��;��"Se�#(2g��b����gXM����k�ݓ��	]8�sݾz����� �d�,.b!�V�"�b�g0C�a#��b�D�:��H./��3L�J4�����9�<�{w�H02|�J�>��^X,i9d��A�VUVμ�l�C�:^�ħI��Ju`.�L�#I����j�p����0�m5M0�dOZ���wԙ�����0�9*wI����'+t�T��j���}.x�v�9����f�[�^����~�צ�>�ٞj.u7���jr^��,���<��՚�,���OdWe�p��R�
��E��'ֿC��'�1,��&���W5��(�P�#YC�˻N0�\�Ĝ�7Rs���c�y�|%�5}-Q��2'}@�s�5��o�&���ƤS�Xׇ�˽�n�r���Xuﭩ�-/��a�oW��U,�[���{���3�,�?�w%�^��ǥ�k�c#;���c��I^Q%��Q���}=3�}��Y���jpwB���(����y��ӊg���JL)��7R�+g�YáJ>�e�[Z��Ÿ�W�XЖi(U@�-���j���I�u9ro7�F6Tݨrn˰�hC�>��k<Ѿ�/U6k�፧��W{�/+�9Or���$��vۢz>Y!ֆK32-
!g+8�Q�YT�1�ｽ���_M�ﵤ�˵�n���df�W�P&+����-@��q�������8՜�(����M"&>�ǆ�";�79�2#�O;	�b���9�O��]V_ik���,�wKj|�^9x\�w�pqE�k���GE�Ӟ���2�4�.�E�9-:kb-$᧦���;�Ӻ�GN���{�킒x>bO���l���z{rq�$6A���Pי}v���#����x5q3�����U�-�ˌJ��1���Y����\���[�j�fI��Wa�A;Э�� ����J��C$�m��m�T\9����(>�\bˆ����y�?C�_WJ{�`����͍B2={��:w��u`bT)\����窡��?�h<��	|7Lsm)!��;����5C���p������L�ۘ���F���'b:q�t�WST�ٸšgf.��u��zG>5ÔL9��r���:!��ҥ1L`&*�t�OS,6�E0����{U[��b^��p	�L��?�����uF<9N�!��COeIOS��j؉�h}t��&�p\H���
�炷x��6��h�S�)��t ���+���gy�v����]����G�f���5�����D��$�]6TX���;��Վ��3U�.��7WX�'l�ՓO��T�m���qJޒKwo?��vcܔ�_~�~]�ϣF-H��e72���}����6�M#iz'������� �k��`��xhO��hQ���H��u�e��u���CCrRykU	<�JK�;P�Ri��+,;�ѱ��&��O���j���W]�)�{j�Y/V�Uk��M�u�]>�{p�3�[�q�_j��Λ���׹�H=g���|}BzBm�ڨZ��V��Oҹ�����`v�kg=�~�J[�E�լ�[k6%��Y8?���֘��R̶�h��:��C.�׾0�8L�s8ԫ[ʌ���ږ(�GR���g��H�{@�x�	�y�:��ʖd�_t�t��,(q�.Ȃ�y.��Uv��Gu3u>�e���C�[:yTI�<Ě?4�,"��������gג*��M)g]Ϝ��-��ג���]��8=�����ϰk���H� ���)<s'jR�S��7Q����͚@�r�}d8ƶc�Gd^�Y!F|������_W:)�~">�������6��N�#�U�'��ƭ�9@KcV�!kߎ��ֲ�$����`}�q�l�W�8�����Bv�o�z7�>�O��mc��$��S�WuIeA�Ί��{� ���v̄Vg���N�{Iȋ�]C�S6��!�[a�t�䍽Ch��'`}�lݧ۵�r�1���^���y�(y�0��RU�x�,lY��2@��T�5�nP�e6:Dg��W����`h>Fg��X�6��a	��-5���h��R{�P�ɦyg5O�Zl��A���9�]���k�j�3)Yv��Ųa�=0;+�4��O5?!)���N�+�Չtū��k�����Q:tw[Ď�ѿQ8(uh���dx~*cCy���^q�[���/KqE?I�sѹJ��n�d]ctS*�IR`���3�w0��ipy����*/�W�iUX<fʘӏ��\h��Ȥ��~�3(�����R=��t$�����y���v�ް�ˍ;��!01��+N҇Gt�������t~n	Ļ�l��_�U%f<���W}�-(��������I͚�`Z���w�Q���Τ�t;��@�ۍ'u�;�]w�y�Z�'4ÇBj��~�a�O���OM0��]�M��
�Z×B�)����ڹ�j&R�S���ݿz�,TɼTB�
�$t$A��v�M90͸�7:m��eRbr�4�N�D��'23���-mذ�/�N=w��_��	�y�(�y�{�G�>
ycSVy=K���4E�{-��A��k�L�5s-w�5��đ��ۻ�z�d�,tt�~��C�"&�>R6���4i���_��W���2A��1���G$�Ւ ]_j��M>��s#4P�i�����w�j�%ڭ� ��٨_�	:��Y�g��U'��ʸ��<��VǤ� �b�t=1l��dtK�{��h|.:�kY��f%3���j��^��/h1��X��F�$=x� �����>/����0�c"Y�H*ft�h7��n�1�簩��k�;Su=�k;�sN�f����+(!\������ڨ�{w	�oa�LdAY�M=r�xd<�ƈ--$(-1������^ܙ�Ԕ�g vPej-�g�w����j�C�][�q��[�.�^_b�O��J�!e�^���=J�%���!5���2t��ټl�S��9Ő-�/bQ�aG�1�煸�  �d�,.D@$<�[ ���n*�k=��@w�1T�����u����:F%�.�����s�:�E|w�@��
%;6r���X��iݥ��J�i$�\����>y�Juk�S*	*Mmc��<͏P�=��'yk�{˦�x����������͊aS},�H�a��Q���'(t	K'�kc��Rm�z��Nt�[����SF���`D�]M��7gd������n�S�&-?,�~��D?!�z��¹�r�5(��|T��K��1����rd�;�Ձ���}�p�P����)��*�߽*����������0cM����h�&TNU�+��M��o��;��u��jB:����� �4�V���pʦ,����j�N+8k6*CQ���.��s={��
�ܺ��{�2E�RãZa�a̹�ud�wk�N�q�E�f��҄��!�)�!Q�/�Gun�<������tX��/�GBr����T���F2�察�d��Fcv�M�p7�e��DAք	��-ai�oVύL3e�[�6�d<~0~Aw�h���x��o�-K��Mv�G��7S����K�a��5����>��{vV���h����.���t�R�������M5���b��B�u�j>����I����0� %�A~���0pxD��T)A�������^xS^��a�n�uA�`8͆��2�V��n���K�}���]:t�@����Z~Ar�>2��o�Ô�'�m��'ٖe�3L��T6���Z��YK5[pe���m�4S��6E;y��R�c��["�&�	�v��mj�'��rN�w��\�ws�)!�������[:3�Z��3��^���@�!'�|Ǧ.g8�;2�Тq�0�/u�$�cQ�A>������-�gII���zD,��fq�@����6Ǫ�3��z/�ﺊ�ۦ��e2F�������.��.`�W�PBO���R5O�z	:����2�s��ܾ$)���(����Z�F��|@DB
9�N���͕�nJ#��Z"���s��G�;v�p��DZg|u���'�׷����C��}��է(�+������ݝ=+f��Q�sI��+7�_�/f�3�}��c�&):�bT)\�L)�\[gT\:�4˴a�����V���{�sz=Х���;f�p��)���Й'�1)�FE#*�qc4���j����;W���
Qm�q���cH�H8�C)ۗn����I�.i�$�,�q]�m�R��[�F�如�p�;�0��B1��O���~�,�v�Q�x���brb�N�3U��)d=!�6Ⱥ��4��^�\�%��>TXX�!�(փ��П���߅e�"vZA��Lv�Cy{:�
�����$��IcH�C	O�ێ��>6σM�\��k�Mҷw��v2�Y�r�n�'b�Տu]E���J���e6���k����n�aY+�����$y���t����T��k(�1��ę��"���XOҹ�r^�K��'[��p�O���Qb#s�0e"�\��'� >5�,�hv�a�@�T��u^�v������|�*"gV�Gu�nd@��<^�:0!޸�	�y�6߯*Y�u}���ܢ������j2,��`��gB�g�S�K@dv�ǌ�0@�?�>aW�p�:j�U\��`�׆�8^NI��׼s�В���s3)� ����¦�l��n���{ӯ��5��)�3ܣ��������"�^�w ��CY��jkh�}�����=���E�{ɻ�_�ƿ���Q��5�b���X⼦��1&��Q��h�����}�g[��ݝ̞��f�Cj
x��C�Pi��I�ʇD����f|�e&��j/�&���Xۭ/ØU��@MFc�_lkH̎A�vA謐�r5�q��t�îyg�z��2���9��7rְ��>�]�cǬ5F5u�ʖ��ۥ!k������-�J�Q���A|EX-��հ�Q�n��ShtS>�M�~�1����b�d�ӵ-�C��M�	�PL�WB�ڱ�j[JZ�e�Nb�ܚS�p� N��M<5��;@@Ŵ��K�8Hg�+�4��<��Bc1CT&��+6rN&y9��R\�`YB*�؍�Ǡ5�з�x���t��xL�c@#�諞�7��wy�����n̤�o��'Z�)��J�
�|��� ���H0͒"�ڙ�)�>���{���/4�j^��5
��P�N��wL-�]g�tS*�#N�@��-A�6���]�����@�Ï}��v4bf���@L�{
6v�8� ⮗�1i��(,k�t�~jN%ע���l]��m`�<�׈9���j�.��/�vT>�;�m���k�3u+Dv�����x�Nx�=P�䆓G�i�[�<!S�^+�r^֥�@C�k�`�%��ͯrs����4�&ua�I[��1�ЬR�|G����MY��:���1����0c��]tgj�����0^8g��zz���56��Ӓ+@��ը�u6��s�pՕT%�O'l=Q�E�'�ˀ���
�tz:��ؖսTZ�XR�XW.�ϛk�u4X��gd<�|Y��e��D��^7��;����@AC�0�y_掯�;��:Y��_�/uc��i�+�&���5c9��1��@��jw)��1a����xy4?��SVy$y]�.?X>��Bsz�����=Q�uHf3㒋�g��qhh�D[��!���xA����I�F5ܶچ�G�w�
&�u�v3]&�����`��H�D��v����;��/O�ӑ[�߯�u�GW<3S��D&��5�{d^������ͻ�Y�� ���R]����$ߪ���x��:t��������Ň��P���Pw�s�/���Ȫf�;(1ƅ��!�do'U��$]���Xs h�_�t�T1U���)&0!e�_y@���J�%��ƕO��f��7뮽!X�-��zPb�h�'�Fq�ј�oV�UX���	�ix +�����C��W�Qp�vj�.#������Tfh�$����vv�v�V[��Ҥ�˓�j|�T���Zv��`��	V5{�j>`ܤ圽����y���+?iu3��
W��f�Y�M���N,�F�`m�˛5]�����i�7q�(h~���9��bY'HĲ"Q��b#��s�:y}4*o9���6�ї��'h�vl@Lk#q�!#�O=y�%:N��:!t�e^IT�����W5��î�dp�ku�^��&+7�����li�r�cЃ�f>�$wQ��<�)9X�R���k�z�\Xꈛs��EgZ�t�}��a�� ��gnO5�uL5�mO�ŧ�b��]�_k�\+�u�� W<�'	M0����C�>��=05��M��t�v}4Р�l�_v�㍌Rq�����!7C�J;��$:yĀ/�G�P��B�Q���>�<�5��8��h��i3��A�5�2��S�K�e'-x��y�+��f��Ͳ63���<~.�׻���ի��-�4���{�е~Q)�Pc�^�ǧնYj�������61���QSI��428�at�scO�?6k�'��4��N	�#4Q1\�_�9e��Q-����'ܞ�����$>�)��/G>08���j?}������s�v�n��;����=����{~������{�����g�����-}-\��Eȴ\�����!�ʹ��5^~���tv! �n�n�F�wv���t�=2��ʃZ�7��L���[R^	���\�jj����,��Y���g/ý�u���ϟ-I�hd���ꤩ��q��-��!����m뙡mM[�U*�n���梞L����t�Yx���]�VwA�7_([�ނq1׷&q��ᜨ��N���&���1�*.��*]�+�Cvr�b}��ƍ�,�&��Db�}H�]@�Z�Lw��\�DkB6���I<[��8��o*���h8�i�5`��]�xlM�Om�u��$�9�+���zg'"�-f�wq��r�M�SV쩸%�'h^��۬�����Rv��|"̣���N��y�7<���<�Ei�}�XW�z�*SMd!�B�W@��6�>��^�o.��/'䪑�s�Ӧ)L��r`�Lc��r�-�½�}����"�Ǖt�M�]f����ǉ`��k�L{]�յ{���e؇K��p�V�_;���LZew)�刻1U����8����=�ߩ���Mi�=ˍ�N�1<�Z򖙁�CmՋ�RY>�hK<C��ķ��+5���9��w>[�w^�`�s���B97X����wS(�&�k}���U�)訝��l�dJ�iP�,%����k�)<k_,���qHv�hvV��5�S���ky�z������{7�(5n���\��4$EK]�֍�z)���_{r�:o�w��g�^��Q���jA�E1��<3��F��t�7���]��.վZ݅?G~ʊx���c1�������[�PS��Q�\�R����Եcs�gtu']��y�.���Y�]/r�}�~��4�lX���Q<��}�i����z��N�6��]d���ZI��%f	]�pi���e�|
ArjD����a�˻�T��)�P�2��z:�5t���c��۔��&�r�Zk�,�+�F�L�Α?Kn���sG,��y/7;3~�)Ǎ>�젌��fi���#bf��+N��հ�d��Ǵ>����B�8K�3�|��5�"�g�ܯ��b��S�Hs��VK��;�-Y�]�mB:���I��2�K�vJ׽�o<��Ɓ���/j���gu�v���B艾�x~�i�rW`�L�=RP��e.�K�Ml��|�<V�.YC�i����t{��nVCb<=&T�\�V�{yH�I��s�"���|��c��&�e�Q)4r�K���������+�{y��-[��'ĠwҮ��&U�J���.nH��+:_l�*�Z~�Ӵ���5z���FS�����%0<Z��s�n�
�9���s�켗�yaRX{�jJrK�����q�/MX`��L�R�yv��wo�E5�;�}iw��ud��\�Qv9�����@�&H���\���>��o�"(�����2RSCCB�DDRU7�Z� �9�'$�M�Px��I@U<�]d��U
D\�j!��CD�kTLP4��S��Jh"����*�[P�C�rR*H�l��CmF��l��RPU�5EEաy	�Cl��5��!��ADIAED:�%��=X��Z�.�ALBPUIV�x㖊i*�	��UF���yk�\�AE5G'��CQ5l�'%��g���CZi�B i3����
3}��F�^��f�|�ƨó��񨵳_/t���B{ѝ����4��Y���p{��ΰG/�^�~�y���V�`��(�M�S4m���G0��EH��)0�.�R�m�e�|�'r��s��^�>������ܗ�_�l'��<-q��/�N�v׳�~y�i�&ݸ�f��b���]�{Q�gj�F��5Y2�"���<����)�0(F0�=Ų/Q���9�	�A�Ku�@u�A��!�pd��3��3gW�����N�,��y����fg��c��=Zo(��M�EcW��	���ըʒ����;�T\9�p�ő
b�4�;�y9�vp��.)�P���5�o�!s��c�1I��T)\�L)�\[E��6�5v�V�l�0}.���8����MЏ�"<'d���gL��xNI�N��j�s���mq9�pn{Ns�^��a��г��!F4ä;��ܻpmΈlԩ2ݐ砢�"����n��5�A�<�܉�lA�.͔��m� ���B~�L9�C!����3uB���R�R��QL���4���|�K�J�Iq\�6~}����n�ɬg]��Z˽U/�="y��U��-B��O6��4��0L����><,:?����x��ɯR����ǜ��	�Eu.ed˫�*om���ͦ���.d��U�MV2q�����u��|�|��� ���U~�,�����b�iT�������M��L�v�V���H�w�G���;��}�xX,�z�^uCe�47�b�?��'����u_�>����i��f�I�`�E�xZ��R8�a����W=�}��RM��s1�A~�2����[Z`(LhOH�����
%k��� .{�PK�XU�V�tƞ�4������z)�1��c.{�>^�!�#��#c��bs��;��j:�l�k^�d��E,�z�[�r�S��UK�z�^�9�"]぀�4Ba	���?|������;�b���ws_A�f��,��3.�
�	�VWˋ_~~!7��(�Մ(�O�>{AF�^?R�j�J��L� ̋/�A!�4��v��-����:��U1�s��&�����is0da�̄��'���{kv k�� ���d^��P�y��m�W�b��,��m���Q���3U3�!0��a8�̚Obj5��	ʖ�Ԡ,~;2�Z��%G\=ip�8c3O�_i�����>Ɋ�T6)�[pL a�s��d�v���?)�ɐ�i^K�];Y��5�n�΄��~];�C�ᩭ��/M�8��s�mF����h�6�����L��3/՚���į%g�*^]lk+��-!^Wn�=�|�=��u��9gvYv��E���" ��F�����=-8��R�m��2o:Ƣ�2��1���\�G�!
�<R�1��E=&!]I�n\��t�_EOi�v��i�?��Hq��}j2$~?��M�_���5B*�ߡ��cξ��{lw�!Ŵy=y!YL$�y�M=�
��Aͮ�O:[5�а�x���pc�:��T��¼��)����� �6KT�*�<"�Od��XIu/����"U�0�;"��5�2���n�eC�n�`Ӗ��]���;pq���F��t3[Lp�Ƅ�M�;
6҇@⮗�1i��%��0��%�C?���
ͳ++X!0���^`���΃����~�SlPNо*L='�s'���&��K/>**8i��چ���^�����;Xtz�Z�ڴuQkd�N0��v��*;(�'��N��z�n�F�i���_��Ϯ�;C������a1���3k���f�|��LI�e�,e��Pݶǻ��@)5̬'����>�z�3<��1a�v2g�`>�E�"���7,��=�s��Ƶ躞��U�!�g�I~,���8��	����ź���^��$�.ڻ�b�XE�9N'�*o^�c5�!���ci���H�D��v-��{|�~7�����/ȏ
˧B滕�r�6v����g�
O7�jbCR;wj{_�C�'b|a������T�k��"�eDg{�>��ޒ��-Ytu�umWJ�bwia���sE�6从hav�HW��D����Jk	���{�σ�z͘�
q���;��?�ש2���C!4�l�ק����H���4��%��
�TH�}-t�G����X�"k>W�Zf��= C�����^�S��[�8�5%L�t�	B���6�y�W����;\_�P�:��J�>��'ƚxX:E;�a>�u�+EA{Q�5��Y�ܚtt����5�]���ޅ��kBSe��A�Z1)�Q�aG�1�z���-��<���0D��@�"��<\��Ξ|�C�f��y��!8��%�t�K#(�k�����l����{Zr࿍��y���c�xvB�D�eL&����O=?D�I� �'X��nI)��n5�����c ����P�����x���a��ʆmɎgݒ��I��e'b��E"�`�f,_ZZ��zUY��[#�������"=>"Sm�c�\����uL4��&�z�F��S=�R�}�Q��_�R	z\�G#�<O��4�1��|����X����WՒ�eW����
6�sUP�]�hF�hdk�[Z����C��_��*,Ht��
#�u�C�<�C����7���a2Y��֙wء�U��^�>Ma�	{[�%,����=�nV���Y鷕�^h�XƱf�����ʛ��{���2�0����@��a\nX��T�Qi-a�u�%��K�-Aq�*{����vmz��&�S|��Wn�K��:%������9���]��پ�����1F�E�8��T�eJUc]�wJN*�O'�W>�j��(k��c'��:B����a�J��ϏudL�|����OBm��BՅ�uQ���q��Q�֒�a�#hC��o%$)�}؜�s;$���������t��|�>˲}�v�^;)86˦��b��5���YE��A��S����/a�k?y�,�8��V�`eHL���� ��$�x;k�<٭��ˢ��<��ԅ�U��VW�`�1�A����0�Ѝ�lNs���ր�o�E[�L�.���c�4/gJ�j	w� �Q�d�կ��m�׶C3��B-�y�-�t�(���bYB퍢H�u�ދef;�,U��H�i��eC�|�П�]�Y�71�u9�G���#��4��D܅��6��PS�y�;'��Y��u�*�z�8�nb�Գwd.��L�s
۷'�f�̸t
��$���8��FB��2ǲa2�-*�Ҩ��O���^K&��M���:�[!u>��ƉE7�(2�p�;g�;�vBnm~�Ƚ�1)�{|�.��6K�(ӧ0?8T�A*��^��gcF��Fn�SU�����f�Wih�n�B��:pS�aX�"£�l��,�P&�U�7Kt+}(����[���t͝%!�Q踵v�Nf�j����'"7��x����6�v�L:!-��o�����ٜs���g֡U�毪�-W�����!?5�~�qnt�T�?vx�s�+���ݩE�k��F���$M�\��L��a��x<05�˚��`�N�{�w�P��\mC��1Ʉ�A1L��n��q���y��6�8zd,|G"�&2"�,�ǃ*158���
W��L*�J疡f�'����ơ���vm�|s}NŌȌ9v	l�jX�p��0CP`��1�W�X��Nl���;'\]����t������<��y��qDR�Ju�������@��,;�?zƕ����
%k���=+�ʂ^ٶXl;F;Xb_���z�6oLƞ�#9��"�{����+KӘ!~��ᫍ0��FOٹ<�7�P0k��Rg����w4u�e�N���f�A�^�^�9��;Y���w�s�˝#UґQ�3��+a�$�h�rf��kXW�1%ڼL�z&dO���5�-��4;�����x�q�o/�oC�z�Y�0���D���3���C���tG��&z�0J������9�
�[���:�^⻮�ɯ/,ڐg�'U?x~�](j�#�6�lYb/���9��UOGYX�z_9m�;j��Z*N�Ƌd��0cu\�����i�K*M��w�c���ڔ{ۺ�}e^���[����{X�	�J�n��*�X���WZ/�T�x��E���s�?�VK�z�=�l�D<6�A/@����ך�i�wd����������n��îyg��:.'�w4^��	�ܠ%��ڔ��`�P��on�oD�)z5sz���_j�p���-��j�g�lyx�A�3�}0��ن�	��10�,�CJ��Ц;xk X�d�.������V�o4���Qm%ĵ�����{�����U��
5������>��'��B*�j�i�	���H��gc�.}�K0ٝ� f6���wL�1��-�$����Z������[�.p�j�Z{?:L4�]��zHN�k�F�G���ϯr��w��_`Zz"�jb�q��dH��ΕGǍ���;�EA=\�*gl���1�p�;w���t@�p2(�1���R��~|��f���mP����N�M����o�[l��<��g��	=� `P|�oX���eG�^��vJ���4=�;yc�bJ��kI�����ѽV$������-嬣2uX.�'�<�8L)3��sd����ƞ���[,�ZF4���en�Bsۤ�ө��w��P>,�{o+�C��}%,J[�&%Uta��2�T���:�� "�T������z�PH��
�̋�O��#��D������f���f��=����\��ϧk���c������4sa��a����R����YH�ಮ��_������Z�ʋ>��cb�h�ٸd�YN��{Q�c1��.������l�����^��H�Ly��֜��6�O���D��mK�)�v���B� ~)P���c������e�-���mB��y��+(�փ�:�*����u l��y!�����D�����P��=7�	���٩���l�6���ٴ�Yh�gńa��v��ebdA"�k���͜��]�@"��H�X����d�Ӛ)�q�ħ����;��t�歁����e���
�q��#*�Ŝ����\�4�(kGMd���8l6C\�5Й]>�n;O�jDs�J��J���n��k���o��gu�Zʛ��)�k�����Lz`��J�н7�/
U/\T�y[�d��~m��V�+Ο���3�6_Q�ɓ���7GH���V���{��[̍��hd�h�����{�S�����\�5{�S�\F�lX������1Zo;��-��F��UV3=MU�
���9���:B�YM�o��t�Hr㑓�ly��ٹb_d���P�u��8�k�k���Ac 2��v���O�J^�LHȱ}5=��f��Y���+�=��>����tÐ�ƽ�5��`g�qNe�c�U��[�5�H�鞳� W$���]�����3u��f<��szշL�Yv���Წ�N*�9T%Kt� iA�>�A�\	�$� ��ﮱ��8s�ƤA�pR�����r�,X��u@3�$e�֥$ħX�9��9z�p�g͞m��v��9����H6��s�e�n�ySk��Y#o�>�4W���Ģ���o�MY�+� �kR����-Z:b[�����/��9I�c�M��02�@��	K�Z(s����j���0�yn���|�x�'}�Di־[j�-Ί��Q���P�fN�Ɗ���+�i�j�רy�����oX$��w�T'jޭ�4��ϕ�,��0h�Y�_U���w���@��^q�T� =�<F����]5j��%F�;.��k���������/���8�o4���:q/0�ci������N���?��u����Wz�k�ِ/y���!��BR����R:Yŉ��{��kX����Q7���cڒ��ah�T�cH=p�"��6e���m��cf�2ň�w�բ��y�WD�"��G+Ѽ�ᣮ�L�TW����\���4�&��s	�� m�p���Q����|�k���ߪ11o6;��rM6R��u>�E�H[��m����vW\nv��^�s��o��)%a�T�"e��G;�/�ݟB[r��L�yه~,�"���=��⏅�؟z�и�ڔ�-�zzXc��F>�4X�p��4����l'��0��=C�*8�:�%Iw�[�᭐���{ԈYOW!���p5S¾�{ ?���%W�џ��98�ܢ�nˋ��|��RO�mgܧ]�t!_�!�0F�s�j��J�,�j��7�����o����{���o���<}~�W��Y�S@����B笣:�.�#����l,2r޾�a����]ڤ�V(��zq�lf�fp�C��*��ݲC�+�����;:+��ҷA@�ƥX��/����u�l���U6����ݽ�a���Zm��$&�̣��'�;�:��K/t��P�KU�0rܛ;��
~^�����Ov���b����Ϫ�zdd7/�x.���j����O\���q�u��;��E�}v��񇂿c�{���V�^����D�=��;9��(K�8���x����'��Yc��۹}+nqs�
����*�n���-�H�d=*ER��QV/c�����|��z�2.�Jvy���ҫ��4��\d̀�Ū��tc��B�d�����jWg�4�t�ia��`�Y��`�q�}���Y�l?�̪��&�L�o	�t�r%�[�a�(�Q�Z��n��G��1��Ox�!�������Ȟ�}��է�Vb�^�UJ6^	И,+=�ߗ(�֎1�����V����)���[+Z9��܅���(��X"	�<��S��^>��{$O�]��B��{A6M+j���~YF���~���`;��9Џm	L�n�X�Ob8�v��v/�EY�t�A�!�k�-�.��C��n�����wZ_K��Om�%P�-F	V�T}<�9�{��	Օwo����ל�ǘ',K��}Fד�LӍ�/�������=��'�`3q��l�ĳ�7suѢ�������"M�#VL�}3������vp��J}�z�p�k,�U7shuD�)�o��|+_2W���KK��W���<#i|#Kf�yP����ǵ6lF��l$o��Sx;]۪'S�z�P+/��;��Y$VJ;�wgM�������"K\�T"�[�亹��7��+�º�N6U�Y-�	a:��&�;�
�<����^X4��k�x͑/z��,�5�i���؅�3Eq{�r`X�mt��*����{�I�s��޻��Uo;\��
��֔�-ʙ��WU^>���O8��L��w^��s��n��{�Vʒ�.�i�t)�Nլo�W7x���K:vԪ�a	�E��	��\��}��&헛�Q��7�=�l7U��Y��|�Y�t��SX�3���Ҫw��PQ>�nv;�3"�}�!0�{��v����C�FRVj<v��1��tX��ٱ��@�8/���9��{�ʘ84>�;�L����2�x�C��-֐�SA�UkfK��iϻ��]ɫ7xM�N�v�6���/�A.D�Ž�m�>��ا���e�u���R��ͱR����[Lu1d|����v���v|� Ŵ�Gyo��{���J�I�c�VM���h`@�w@�w�	�o G�ڶ:�X~y�//�/n?z*����h���ѣ�����y�y��ξ��u
P��PRPA�"
<C�F��Ҙ��j�i�������R��	�B�%4�tP�IM6��U1TP3-@r4�Ts��)4��
Jj幌�%#�a��yP�JS@�5�D�I
t=sSUEQUG0������u��4����Q.�CATą5IE� ��CF��T�]i5B�41HP�m�)(�"J@bCc�M�MA�+���Ph��,N�A�� 9�*�K�6�KO'Erُ�hnם����quG�s2�ވFК
�;��u��,�;78F��v����GL}}1U�(�dܕ�=���������od��g�g��ܿ��#l�t��ހ�\s�܁���]9��ؚ�ֹ�}�}G�ņ��0D��|Ǽ��/@�b{��h��+4F��g��2D�����h��6�}�����,ϱo{�6�ڡ��x���Q�x�p�l��Iǚ���ק�
�q���`����Ӽ3S"F����ں��јHy�Y�TF�L��F��C���箺z_�觌�z�k�7 e�ϱ"�������;^�72�5�n�;�/-\K�쳑O��~��.�&�5��Y�h]2Y��������Gh	m����r*i̊�t	�Jڟez!j;��M	|]���Q��_o&(g�0��T"��n�i�zi��vT�g�WB"7:�#[p���Ғ�0��:	%P~���u�o�b7]���~��7{{X^���J֡���Dmh1�ġ�Yo�YK&[���z�=�d�����
���x�u�	�4@s�?��s��>�ΰl�a>o�ǳ�����{�5Ϝ~Fxq�E��vj~":to���yp���ơ�
�[�8K��)z���0�~3��^�pV:���$��#��t���մ�:�*�������Y�Z+���}��hO���Q�Rk��i.ǹ�<����(��n���a]C��|��'��d�B�3��\���͑��7es�n�y��k�a^�n3�'��7�-���\]D���ӛ�9L�	汽0z2���@/(&�Ud���O��`G9KD��@�_WQi��[��/�.�g�H�^�سy��� ���Hm��ۊ�A2-��Gnn���*UBg�	�>疩��Sq~��Kr�I-�6�����j�)����;�쎀��]��W��{�~�Ĩn���e�i$I �M���{��9�S�����m�tRǗ��;�+��X.r�tg���6��޾/ܑ�YZ�:G$?��W,�#�h����CW3y��?��Ez�Ѣ��}s0$�bb�9���eӭR����r�!=�<��Ef�_!�<���^z�1_��M��1�s4w�Q��w<�yBg�1�d4���՘��i�}x�T��N�'����"����)����k�{�l�RK�;hD�l�8�ɼv�Y�wd�V)U�TM3���0�Z�o��-�s6A&�Ԏ4�fڹd}�L��݄m�E"����weG
��ؙ��U���OkIAw�A�OZ�{2ni��8���5�F+�᝼;E���W>��j�/kd�
�2����� �߱�	�����դnY�l��(�<�7$��l���#\�Mx�J�u�nM�KM0��.wy�����]�~�5�O�Z#��@�mS���	-jzeRf9��i�mv1������H�˨p�f>���Z�7i�D��z��9#go_]^������T����l��st��F�caL��e�����ju����3��:�i)⻥v<y�ٷ����m��<2�>����Rp�r�8�ǥQ.np�H��b�i���%si���6�EUnN/�7�8��	�v���i�Ju2մ8�Ux���涶����KY�f�}�8��Z��j�=���M���s*}��)ǹ5�˭Ŭ�x�把�_Y�ںF�*\b`�T�����͐��ms%����u�pܞ�e�>gp<�U0���o�z��ݲ6��������#~*J>�=��`stF�K�Q��e\�fu��嵹�q����<��.n�v42�ù��1�J��)�j«����˂�tm,1�7o�u\� h�|}�.��6��5��hFX�ҧ�tL��΍"�0O��"y�	;,H�P�y���} S��Y��iV�^'�-tI"s�s�2�y�Di�唵������#���ݕw�R3j��{R5��no3#֊]�����h���<��L4��u�V�Tl]��~C6X�G��q6���+�#�).��
����{YJ';_o,��3�� l[܍L�]z�(w��z�|]��+�Q�S�]w�v��Z����uE.�y�OL��[�,m�v.�N=Ⴌg�}5��9���W���y"��5A���r�Of@�nH\��56؂���QM�˛���ބM�|���*BD���\g����4C��/�����M1����E�t�dU�_йW�m>�d��F:�wT�þU���)�m	_�"V�0���]u��O3�=�H�:J\��؞\O�Z�<w�3���s���8>c������� ��PV%�d�(~�&�R�>u��m�q��Ǘ(�M���0:Ԫ�\�^=+���>�[d���5��7*�#g,�~��41�к�������WbK�kXzy��i$��I�	�e�1U>*<�Vk�>�j�0����oP����;*��+]�"uq-]�E�ގ��dv�^�ކ���͏0�
����M*򅋔dl6�f�Tɫ������{xҵ]hl���7�4s8#zb�p�D���Ɋ�7wWSK�����w�˧+L\�F�a�F�$p,�1�X�#<���j����n������ŝ��\d��H��&��nds}�k��V�/5��0��xj���)��Ŝ�|��øve��;�OGc�^�����˱/vW�����<�:9)3u�ߊ���L��cj�ss	�{}�Ȉo������nÆx�9��L��N�<l5ԂP�M��ˋ����� �1d���{��XfJ�%_��#�^^p�e���{��k�ֽN��s�r�;'7gp�0��QKGpO���xj��i���8*�䡑k�,���Q�����{{�<{´�uS>0�M`s�,��21��Mُ���M��v���v^��R�R�	������e����%�!T��႖$N����f�f�c�t[�߁�����IIP�eP�nN��W��ȫg@���N�gS=��ƍ�5�ţ�="��3�x�}4�v��B��'�u�W�n�m2�����=u�ܨP��5��xvH�0�u�|pwJHK�ɐI*�����<�3eee�����wx%��~Kjx�@eϤwQWh�*ۻԛ5������e���MkN�5W�F�ټ��Y!���|�\y��d�ճ��hON8]9Ѷ*zɪ9�]�Y��ku�y�L���Q���~�0�/#��a�
���ţ����;�^���>��7��/���i��i���!�<�z��J�m���rG(�N�����\F��$4��&����ȹ�O~��N[�6�升Bv�u�FDzC��>ɯ2��4kal�a��S�Lt��!��^}�N��Y��C��(u�a�S������~�̐ռ���gnUԜ�DZl.LP]�ݜ�ƅ��Z"��b� ��)��z�7�c������9,nܓm��I����s���e�G(l'5�1d��4SC�v)wi��5yI�v*m/M,l�6�����l�(�]�3��ٵoH���Ϗ���k���� �-���m�������S�m\IU
㣷��>!�����xVkg�n���ǆ��ʻviG��˳�>m8u�ׂ�����q����T#�(�l]���
x�3�N�����ϯJ�	dy�/"�����g%�X耂5R>�#1�GGMsl"Zݣ0���x��n-1���	� i$m�6��+�j�K�ŵ�߶�M,���e�Mŭظ�D+�PSJ	=KA��4�A��2n��������#u�ǆ�h�r �ի֍@��J����z�n�W>�έ����9F��*U?!V� NEH�T�7�7�|ڔ�k���p���gNٷ�ѬjV��>��s:{��uB�Q�ڤns�T��J؅g�j{N��`��>m�$��l�f<��A�9f8i��G�b�j���|B��r�W�UZ��_�ia�ltS���ͩ�ﲷ6���y��н�7vs�gl��7��eN�k��8�x�Y�������`��{�m-ڐ�g���/'�Q��_�E�X�t�&&��{݌뢤��+�>y�s���jI���s�܇����h�~�Lr 9���T�7@-��oM0譞��z��{D��8��f��a��Pˎ���hܷ���kS8`d�>��5R�ŉ�X3i6�?"6w�t�4��w�n��j��.�a��d)[=w�*bl��#5��z���/ݛfQ
�cqݣX���2�7���]��tOv���[A�"�����;��B�0���<�y�e���t<��0�۲�'F���=Gp�Pc GzZ4s>�V׮y$�ב�'���:�m�`���<õ��@����ctr�	惢��1�j�� ����L��W�����j���/^f�>�~����ꧠ���=�;�00��Ev�
x��V����e�L��T=�ډ�����b�;���h%�nT]Y�����<_g��6���!���5Tu��]B2.F�|��u4�S�=;iI隼VFP�0opה;Z����D���l�f��gD�;]O�q�쮠�8��+��/��+�4�G��Ut����w�q�dP��׹��rF}��Y����%��Ep�������-�ֽ�Lh�j��[$F�g&��L������攎U�[�"0e�)Ϛݝ]nQ�_g n�A�~-Z4#H�!]��w�t/_�S�eƤ��!��~��]�M<�P@�\�B6����Og;Hۮ2�}1)<%I!���jF庑ّ"�$��L���O�C.z�:�-�����#lǷc���@H��=cp�u����M����ʜ
S�@`�����v�,��u�TJ�5.�Y��ie�����{�p�F�i|��=>���:��v%TqtMJ�K�٣9Ww���ޖn�Q����W͐�?��cj�}���2vU��z����3�oK/N>d��wA��&��a��ހÝ��@<����M"�#"r�+��d��-�K_8�#$��P;Cg��}#G3��16��z�X�]�3���ԧ��ԡf/��a�hg�<{�~���>��⌃ϼ���Ϊ�m}��x�̕����fQ}�߳}uC���y����l�*��� ��S��Z=��hܼ�>->8�F��Mj����XF����pu�LCB����u[{.���շu�q9�ޏ�ｪQ����;<~,�`���p5!�̬��`ͥ�z8ω��`�N�>��I��Eh����Us�	ʯ!����k���A,F�`d�D�y��WY}a���fz��ٯFz�������#!�*Y���)uu׻^h���;����e�fzI�[�<��M��E<�z�BP�rk�1���g3=34�7��/!�Gjn�G���V�.��^Z�sNdl��
z�?y]@�鍮yZ��[N��GB��,�N�V���ω�fUͽ�[<�`F.f��Pf�X���0j�����?p���v���0�y*����܍�M+#\FUd�SY�5����H�z�<D=q��]�p4BK`�$���
��6X�&k�I�7�Q6S�ӂ*<�-�<p]E�n�%h�(����72)D����b��1��|O_O�6�
 �>��6���8q>�u���_�y{�����w�����}�>>o_�������Kr~�;���D����������!�q�/3fp����+�咩�V�'���=�s��מ�N��p��Lo�1��}r��V�l������ػ:�V�uZ0��#v��6]��[i;��Ε��7�ɣ#�ش�;�#���w:j�Ѫ堻�Ǒ�e�U(�Ռ$U�/�;3ԣ��̕���Z��(I2�w;�����,{�F�!�Go0T����K�s_v7�\4x@&kփ>�&�qb�:�v���h�.MP��	^�%i�DbɃ��骙o����̺�)WV��ˡ&*�M.KL�%w������(e���m�S�`�[�:�7n`5R��kOg�WKXF�W�-'�vX���o+��R�T�].��O,w��t[9�G;�o$P��x�ʛ�v�ӓ.b������.�wO���78�]d�(�=�%`�;�MQ+oV��u�閯-9��ƕ�tӺ:��#X� ��ɀg��7�eh��s9_gr��VH�K'G�7E�Q�3�J�T넽��ǽ)��us���%�#��p�1�7%�<����#����}s�e��h� �b/N\�qM�;���)ۖ8���7.Zl%��>w�L�0�;dY/zS#��
�8�i�ʴ*VD�]
{�O+N��k�����/�U0��5�ɟ5t�aW�>�peЦ*��Y]p� ~�q5b�����Z��_F�=�E��W���Zy~Чl�8�S1Jb����B�_W[���"��=��,���W�*wК;yƖ�����'�t�	Ɋw[�t�@@��qH\c��}��8���:u����/����}R�dH�����������̗[��|!�)�5�Я��i"�ʯu�� ��M����sU��=3��n�����	�1
&���� w���Q@�H|��
��s��hg��>�f�rU�84ӹa�eG�`,�P��r]����n\Q���Sκx��t�9miYZ\�����S����u��ZTjC�/uv��1�wn�Җ�ȵ����QM�����[Z5Ż��{���rr�UJ��V��qnWJ�m;ǁ <�r�9N;(ԁ<*��i��,�;����nm��.�~[�(��F�/�w�S�Y���m4:���u�o�]l�}���M3��j8�M[\V�V{��8�X��1ᾭ���j�IpX�mخe䪫*��.�Ufut�l'�5]VONTu�lJ��!+�Fv�'��t�s(ɻ�4/<�
.;9��|�,�}�r���v�~�u�e�ը��-V�q;��cN��sV����3!��&�4G��P�I.�j*�ݏP)�D�f�m�n�`Y����9��,�P����v��uȜ}�gH�_oj�q��z�V�]ؠ�I�����nQ0�Zh>�ϔ�9ם�
\6Fn�.��wFd�6uu���t�C��X׈��s��$��fw�sŵ�r䋭�/��<�۳�]s��)��<�n�AHRW{.���HRPV��
!���rնi-�M1:F��#�5[gA���I�4�n@�Ll��i֓V�7d��!+[X�����n�:�C��1E/#I�4����@[S�jZtg[A��l��4�ѱj�m���Z��8����F�"(���bt4GF��N��:ClRӤ�1hm�E-.-D5�fִ�bڶ#V��4Y5�M:��T���0r��1m��Pi���-$M�\�\�4Ѥ��+@b4D���CC�����Z�m�EV�f����Mъ����(����4Q4d֊4�8ѩtճEU:4���
J��h��g�()�1!�`��h�g�w�[���tWF��E��S��@cbU>N�V�J9�p�ٸВ�Q��?��)O����lZs�g8���]��Np�3��$�l��k׌s�8���ߖ��G !1�I�p�"�2
�2�H�$fT.F�A�D��W��j�z��2����@i�w���+H����=��W@`��m�+�WC�,�L�TZ=�U��3]r���W^E,/ ��7�Oޢ�_�F�ON1���1�?o�]��ɣ6hl���Xo�6���
�����o�7đ�2b������B����>:��4����pѣGG��o)�/�v��we��[[�����#�0p��S8ь���>ّ�$n��G�t`�n�ǥf��C��ma9]۩�}����Gt��7��W�Fǻ,��xq�[F�g4��־�J}�鸉����\�w��ċ���',������9<��H�VJח:0	g��  ��<�D����vtEB�*�O�T�#'x�=hAbm*�֭�W:�:����<>m<�u�1����G�p�ِb��\d�Do��Au($�-=�^>���؆�8��T�k�F�D���w~��Fk����H��ۮ5�k�3Ͷ��V�.�`D��m�;�x��t�î!v��ҫ(]"�"��p+G�rfj�F�!k�o.�+�DK���4��J$��F�p'r��l��A�򫈃2Ex��:�E:M'.��{�~��?u��d����T���P*��+�Jqc�~ӥ�9�R�.�Yk�Y;'f���E��/�`l��SN��n���jE��H�g��� 4������vp���@¨�EH��ޖ��N ����Q�Ԅ2���i��ڼR���w�X�#`���N��X��-���c�!������qH
���/�EMir�[Yϝ����޴��rѽZ�z�#;H�p�M�v(�X��֒�(���
G�M���2b�s���a��V&�C�q��W�hу�@�S�[�+Ɣ��N��Pӝ���Ɗ�tu���<Æ(oC���;�w*0WPe�OK;NMs�v�FK�f^��;���`�lm�����>ԯ�V��;3u��{�&"�N��~�}��eR]�;BLt��zC��`�~+��������ؖȍ|��11��:�t�sL�wx�s;d���9��&k�{1���*��2�:�*��Q���^^Ow;�d�j���#��fg�\�?Z4�g�t�'��ݕމ�V��Ma\^M/ͲmF��т���ew(!��Qg�����Ue���Sv��
��!@�gLp�w?��<�tQ���C \v�"�����&Oj�����[7g�n�̴��W�b9m��\����b��^��z��3A`�a��x�VV�h��wa���AۯA����R:�ms��>��;�_A����G��OTM��#RYC��9��ˍ��n�7���];�v��[�OhagAd���~-Z/��[��wM΍n��	k�����@�ʏ]�K�g��("��6F2f�t��t�V�0n3l]�!�$l�%IƸ��S�n�v`$^�aЋ.�����[�(�c-���n�@nI+ҧ�6vک���E+��~�����S��C�ҏ�_����fek:���\�^=+���)�h(։��M��F̎�Ξ�q��a/�,�:�$ړ^�*��D�4�z=!�6����\�o��u�9���5�bxL�5�d�e6�^�g[P-H�ևY�`ھfȚ�Irz��M?,y������2W+�;4�Mg+aj���k���*+�Z���˺wG�݊f����p�!��wf���֎I�n�}�x���޿���ϽtT�Py`/��z6J��';)<�9�^�WD�ٽ �c_W$b�n�7��l3c�5�>]S�kq��L>��S��{y���W b�x����J®��7���ͣ��C��D�k�4*:�O.���d
�|�x�F�˧(i����l���Q8Y��K�Vk���1~���9C�����sF��C��$�rLv	�E�n8c�]�H��ʚƋ�pΰ��2�<���ѻm��@�H�]�/&f�U��[��j:s��!�*��M�!>�a�\�X��͟�?c��|��p��Z���~�ot9�x��މ��&��S�O��;� �����/r���|��!�ՠ��Q�_%���ԭ%��yjni���
��fً�3ϵˮ(Ω��w�FDxv����UhʨF����7V���H��"����/z�^�\�d�x�[�÷{=��GJ����9U|572��i�dadm�V���ގ@��B�� ����I�겺"����	�cE�iWu�4Y��$���t�sܻ�����ϑ��p��R�<���'96��l���Jd�k*C��{c7�����SNՆH�:i:�/	 �������b;#˨��0�y*���}�/]WN�#vj���f�&��8��_$3 ��"����*ձ��-�8vm�'խf��]=n8zn7���ev��H�rV��Q\u�^=�<�[b��+�x��q�gFj�or�}�冏Wg���
 ����s۝'�Ȧ��g�5�A��_�kc�c��]�\_���v�ǘWCK0Y>~&�ңWw:�DU��7w#v�٤k�mP����8��6����7�v*:�/\U��ޘȑI�f�F�TL���'��H��=+=��[n6=Z��gG?g�	{�	W�7'۝J�������	~�����mh�|ӗ�w5��w���g�L�l!�6#d���=���2��	�v��\v�e�f���	��+�u�h����~����īX~����&�z����en)w|�#�����Q��onP�sr�fQF}�/�%-�V7�Q�r�2Sl{x�]]����yu�F7R��.,v��xzĪwO��G9l�Z�f-y���81
�L���8��o�N�k&�Cݯu��V��DO���%)��[oh,���2{y�:���$���Z;�؏Tu{!�p��ԑ043�t]jֺ�ؼ��':�9q]�����+�E�VR��s��X�My�Z,eke%q���6}�4Nu�;����P�ց�iPH�O�mH�e	� ���pr�=Wԑp'���@1�l1����M�Qq��W�E4��ԞSq�}}t��q~��Χ��~4����p��Z��l���q����3(��Wi�8鮖�;��D� �܍V�}V� �r)�Y��#�r��oS�""�d��:c������A*������N��t�?�nj��ɽb6+�!�������0���V��	�����xn����I~���Y�o6���p�1�ǲ�϶��m$��C-����c�Ӄ����-�}79���ᡎ��}Hٕ��s�;Ȯ�-����K�v;���ֶ�����(�=yF����&H7�c�Z�l}IQ��/��ixdO�Z�u�\��X�)��:�&kk��*XC:љ����eĺvNcl���d��^��f�����lQ����Ź<:�r^�[{�������Q{�v��n���a�}Gls}��7��4h�ʯJE-�� ���LHrn�H�K2��7�Á�o!��7�d�vN�@�\[UG0�'�ER~�9�^�m���UFt䌽����0��!m*��uκ��Y�A�~���Ӧ�����[�4W����G�+��U���Gj���S�ʹ��0l���GU���,�v$�{ޕ�3�M�Z�Ы�~�'aʼl#��k͕�n��!���+Ј�i�崻o9�Q��z��(6�e�ZoKfQ5uY�i!�dq �@Ч���Ŭ�Ә�=�ݣ#��j�	5Tu��ꌋ��,���n��޾��Ͷ�?t������aĕ=����ǲ=q.gu�v��-Z+-�H;=U-�_ece������6��N�L�����y�O4�= ("���C[F�2�p�z6/�%�5�]��K�`�����/��^��k��6p"@��r��������Co�{����"�O���d���zt�C���!f��ױm�U���w0B���_KM!��L;s�&�ҳ�u8m5yW���R�׋6h��+m�r�4Y�o�j+�/	REK�5^|�Z��u=��q�����j������uvt)�{m�����	���&J��)"tC�ot9J��ܪ���}��x8�W޿�2.�nم�_��и�ڗu�s�D3�&���:{�o-��/�C	r��.u��g��8� ���wӓOo3y��2�v�w�H;Τ(`�q��>`��o`��QW�6���U(�YzM���P�]�+ʷd�פ���f��>�v0(��Z�5,���mb�&��\*姫�/j��u+
��=M�7�4su;�Q�Z;�/�4������4.4.>�Z��rtoa�h1�b��S�du�ݣ�H�1�jA�Z��T������"I�z����/��h��n�NɘB0�WK���,ꍁy�� ��$���=�����3�_a�{�j����ҝ��'�_�8��eOx�H�e��o��z�PU�>��X�$�K���-�:�˸u-$��u�|Э���W=�q�®!�"�'�@�8�U��Dtۣ�r��ܴ(��[t��G���C^R���M���o�s�l�7.G�*��4�)6������pA�Y����ں���s�(E���X�\���ȼ:HF�|ok�Qh�U�����)CA�E�v�`���d��)i��j|�[O��4�@�gg�/#�9���y��C�<㰺����ё�t9.�pI��@[w"���*���-&�7��4F���#Fި��#�V���(V�Gx�U�}�ܖ�Y��eg�p�쮽�"��=4�\$FH��u���\wJJ���R��̓US��Fm���9S��s������W�^9��T��ʸW=9=��S�u�oR*�n�!gl����A�t0�B÷��wA�#���<��*�rEkW��}��M��I3��l+�����I�Mo���87gh��9���&w�=O�wM��`�w��S���vn~�r>�۝y<[�\�3�
����H��n�{f���=0�w-whqf��`�fV��}U�#s��ͳس���{vd�%}a���r�j޿J�te]��0��5��do����k���x6W��گ]�ewQ��!����:�Z���*�����m�<7S� w��F��tɞ��G�≘��<j�<5��܆n����%���NW�|��C�	C�G`n`�H��nÔ7����6�7�Q�w��lF�n�L㭘���Y�d������l�-����u�3D�;�����Қ�-�6)��U�	/0�8���e�6��F����f�{)<�H��N7v
26)�r�wB�aܣ�b�{��Y@#�+{t]�9�Mx�C�l����s d���:�*���u�w��L�j��
;7#5$:��M�A#� fڊ�l"2%��`��.%��ڈ�g�<,-���M�Qq������kp��m>����33ܝ��ʮ����ٓ�~�AQ��"'Ǆ�ַjU�b�UWӒ�=�ו���s�M=2v�}��M[<�9>�T�7�?������^�w����{���o������/���5=��Y��s�:��dC��T����x	�ͅn���Hy���'��j���Ao%�eX��x�H+���cY1��u��=�=_wH���+��(��"��Q��5���
�{��˻��g�u2������r3�����p���Y�V�2��"i����و��i\��>��ǎC5�$~[seB��;�M�G�n�����=Z��^� �;%@U��+���f�{7�f��p�H��`�]��ݳ	��������A�h�{Jg2a�W;�e��kc�,���U���ƺ���=��5u.�����ʞMJﳻ�<����N3�4l�5�&��,��@�l���E%��z0b�ޱ
ꤩ��Ÿ��k]t��LM�'�Os��κ0�X��+E�x)���k��7^�^���E� A`I4��rbw)��iz��<~�4{��{�p9�ow�Rt��8%&R�����NỊ��0�O7)��9��������ѵ���s��c�m�^n�r
Y���ڇ-%����*1��_up�SDTrc���h��N���&�8��cSû�+�i�s7:�ŵt�Y�}�&�kYm����;tإZ�)Ѭ���卷��3�[ú�I�Yz��PX��쓳@�Rק7U�F�@���U��KW��컖V�{�=�{���v=ycS'��:�2n�չC��}RL}��=�	W��i��o��'��/�+7�l�"��Iܲ��\uKc�t]�,��X[j�{Q߃�*�ᬺ0-Rza��CE�[�2�h��x��GY*�`��klr���:��8mJ5o^�):B�.W�{\���M֪"WN�K.�k���UJk��T^�	i�<���@�Y/]�t������43�0uk�;#�I���4��8]���]�S��>���~��!7��y�(�=d4{$���\�d�y��,���)�[�����cÆ�����osZ�H�6����#�*#�.�$]��,�$Z��lN.���ox��Z{&-��gz?���|.+�˥bf�"��slǧZTkj�(�E�u�"��$o��Ǯw�b{W���yX=;�
rw �	�K�ٹ�څ����F?ֲc��nq�w��:LKZ:�ۖa<\0������#6�1��ҝ>98�r�Zo[n����Ӻ��r��\F:([3�F�R��ts����aATO=��{&�{�\O����Ϸ=�ƯԔ�c�pym8ڰ�ڔ��p�NEL1�~�n�-A\����e�u�I�u�d{�{�$v3&r��
���.S�+�8�D�Y���_L���M��y�V�.v��g�����H�W琗R�\$ͳ�}z&^=�U[�(U@���XVR�6Ƽw��Ӹ#}���fn{[��6L]1�y�5=�:��g���>��Y}vF�� s�_�6��=ʫ���g�fԗt�{���|����x�E�[Yѣ��NEk;X4Q�
W��涢�%kCI�U�"MAE�K���&���\M��a��F-L����b�ؼs�scEj��F�k%;��)�9��:�:���M�F(��J
�j�X�tZŶ"�A�9m�l��CAKM1-IU\��0E�M$T�r�(��`�� ���+AԴ�Q�M��Ж���cG6*��5Qu�IA����USW0��� ��Ѩ���Ѫ�)*���vƊ���ք�")��V ��*���ت���&9�sb�ӶEa�& ��ö�Д�T������4cl�r1��7�0�v�����?��}|��������Z�P���N�	FƆU��X�ra}�,TUGUX�M+p��$�v˛T��Ṅ���m�͝C�&���ْ;�����*H���}r�Ɨ�E'�\����{��f��3t����ܸ�m�,	>(�Z�6c��S����f�fg�m��w�0�8�s�A@ۃ>�Od��ir�[9�|;eXu�o;�崕\0��f[q-�w@r5N̮�t��v)�\��%4�u���/3 ]�f����{����8f�a��ȍ�T:M��<y-i��ȵV��sN��I���=JP�L��C6ޏ8(��"ƽ����/�/Yj<����L?�
�ږ�+���vP���Z<�o��@~�sbF(�aha2�O=�f�Û�#���;*� � ���Pc�t3��9�jn�f�������et�s�����'�à�>�'�q�y�~�g���>��5[��F�1��;!�)��Y6���'�Q��{}�j��������_���j��L�ZqRn�mm]�瓶�������@�|ޮȻ�-�Q���F޿��Ϡ�=7�D{�����P[��L�9Hz7����^��k��F�m�#���X�u�}��*���ȁǳ�%��}���q)���)��g�����b�'Å�x�B��F�"j�2�GP� نb&��]����{�²�v��Dz��_ʠ�5��A�Lơg�FE�ܢ5����Ea��Q�s�颥%��z����ǬA�;�/�6+7|7bo�w��vq(<dt����~�(�d���k<�p��Rr�S�����#c�Q�іF�f��$l��$S3�ϖ�n[�⡄55;;�TVɬ(k���0��d�0�p��݄��7$��Z�-�}q�s�7lQ���ݣX9�C��u�c��H�[l����~���y�K���y@�n7]���|�V�)�?Ha���@���t��fz�ؕ:w�z���;N6�d_WA�8�I�x
��0�l�Cv!�oTl�
�����5���;��	���-�ޯ�˹E[�oc���#6��o��ekh��z��k�U�x�5�7V��J�����J��2
�E��ň�8�)WE��s�3m_`�z<]>��n���0U�7�p� ���f�ps�;`{�5�ZV\F����!�u])�Yu���?8��j��s��	b38W���;;C��Ǹ��u�܎�q�%����#�#�Wj��u+
�<v���o���du��v��[�󰽄/p���\�4�i�NV����6a��y^������~G�6��$!=���93�vd��0d�Ƹ�ǘ�R�[�VXE�sM��3�𑎛%�� ���/��:�`F^#`w��l�ZL��5}�u�_����P����=*ǘ�g��@��f��׫����ҕ��׭��GU��e}gk�y��q�'�y4��S�xC��	��^�X)��D�m]�1��n&�7���AM+��.��yjni̍��ځК�ufQ�����QF��]�ե>9:���+FB7>;w=s��	�������1R������0>�=�r�#V=�� �L#ǒ�sOpC���;Nٍ7&��H|����&��"2a(�b �3�),��ǕU�M�f����}�`�D����L��,H`˘��a�W*G9��d���m�/k������C_�C�q�{��(Ǵ�3�W��Z�96��^E� Č�����9Ž��+����N�t��n�~T��j����}��[����_
�ٽ�L�$�}pp�l����ȭ���_��.�-�b3o��Z��5�9��;��K����;dw_O���
A	�e�"��{^�C���q������$�}�;�uXH�\_�����+�k"����]j]:�B�����&��K�ݫj���K��&�I�4�wm�n���#Ed�-덝=�tu�,%�Q4}*����7yc)�S(�qy)��b9��q�����Ԩ��nÝ������NOmvML�ի�~��b`�nQc��Fl�HY;���MLǮ�7��m��u1�}�e�8�gs�{t_OPg��8C�6��X!��ŵ^���۱_+ލ(jo2�����$HXƝh�gb��-��6�<<��0�����������3����̤|3����Ee-Qx���X>cT�lG6��;I���/����M�ܸ���9����ރ/��"k�E��6{�Vm^�D˽�N�>��xQ���m*w��mj��_uR}AF{�r�oO�Y���~
�Gr<�e�&aХif.F0�q�UqSC_p�.]i[���7\�_:O���4�&�~����RB}ց�@��#�������e�KKf�/�my�`���{�	����	����YA;�1����ASB&���l�]w�wo��]�q.o�QB:��a=�����lrE��$�dK���x�x�÷s��"��@/��������ݐ�f�3�ۂ��Q|ְE�{Xq'y��%R��UO����]����׻�����V~�ر��1z�׽ ��t�FF�<wJHr�28�	��	�3�.�����=�A>U��F���ǆ�z�6�SH��a����j��f�הg�2�ofl�7m��Y���׳+���mrמ�R��7���O�Xox�nH���nuu�	��G�q�FΪ�4h9C{ �2Ds�ֺo1��R�q߇���n��h���/����'O��V�]��U<��?��-���^����s�Mc$:yo>��o��\\��űpؽ���+�$�l�*eh�"z�p�4^��_^n�A:t+u^����c���;~j��K�
2�� ����-+�Y��ޕ���Է�}b�7�h�ɸx�Y:�7�����;�L�mq�o� 퍛���7��8.1�|��t�@���Sny/u.����8�W��X�����A��6��O~�o?��ԯtu%��*T�f���.V;���c����A<�tQ֘�el�*I�~���RDK��6���AҊ5튴l��l�=�H���Of�:c�]U�&��#����!�o�40���ѯD��̴H���k�{�51}���7��\i���gڭ�����PJ�z�n;�b1c;Q�l�*�^��7y�����o( Ϩ�T�i ����20����]z�I~��-a�Iun"&_�r��xw����r3�,��RR�йUٓ�^������{bx�y��G`����$ m����[JF�xJ�E1�8�jWs��v��fHŷ�9���P
P��o�R;��ѻ�$��*��V��*("Af��;��Q7��U&"��1^2\SH���m�*��U&��M��c	CZ�}j�̨z�(s�	��zE��Y��"�����,Ԁ�Ul������|�6C��2�e�֥�}]N�;/%Zf��_fnum	��cPF;h�����5q��Y���Յ�����"Hw��N�n8��.r7v̪�/rT�(H�ܜ����]�ӏٝ�����m�zx{=z�:�v���1�|��Y��ծ�{q(�T�]��
?�!���,�ռ_5=X�N��
����]��N\N�;M0�<�Z�QAV��t�q���Fk�ıtL=6!�r���L�7�
�|Ioj�J/ɗj�{�Z��I�=M�	�%�(��1���	��u�Up�e��VԶ�eӔ4��to4kGs�h0�.����Q�A���0��2BS�+�>�\N��T�lWv6��e�ӗGtl��3��.gUǡ?C8@���ά���߻�D�o7Y͛O���Y��!�}bGr"}ǘ���|��!f zJrY��,���4nW�Z��qoe������VD�<�}{jGF�k4H�X~���[Y_�;�����'v���U1y��Ȉ���h\6��R�T�͢Z�/d�j=;U��`C��q���O"n�T��V֜=D���{�!ɫ�=s��M}s���ݳ[��E���<'M��j�h�|���֜�u�������\\�%�PDR�)u��*�4Ӝ[���:�ُ�f�`��z<�8bĸFDv�����*�eT.��R�B��Py��)��nܬ�~aQH	�u5lへY7>tDXD���܂��z8����^�>�d"�x��ޭ��b�MS�܍�3MP:���J�[o��%����[���]�=�� <�$��?_�W�o8"�Em	���*11����y�z�F��=��zIV4���*V?�\w_O�����0fM�avf�ĭ��R�;<Ä酪{6UONw��3z�"d./����鬎;�}A{�-�o���P!u��յ^�ȥ��q�kI��n�8�N�*��ޖBs]��j�p��FΪ2��f�亊&�����}{; 9Fu4��� ]'���9h8չR7'۝J�aj�zw-�y�Y�muV�@�1"v�cY֝͵w���T~���U��_���o��Tߝ{���{����c )������*-]�<Ӡ�x��(؇r�g�8)��r��f��v�T�p�2++& �ٍ>�wJ@��-�,��h4����ns��8v�-�B�9���ͣQ����Oǧ�`�a�c��[h��B�1ú��.��7����o�:�P/�>�n�ѳ�/�u}v|:�Ӂ H�m��َ-m�M�S&�nw"�H��3Ge���D��u�݂��S��Ү�
�79�� ��:�Ւ�v���3���X��-Y+s1t\���-osq��7��] *Y���
��D���ٹ:�:�2	��nS閨~.��eZ�����p��7-ײ�Ղ`=�ʛ&�\f��P����Y�]6cc�s�ws����^=�"ת�P��¨#�D�Y�GT9�/c���q����k������YB�4��ݻ��+�WlE���o��S�nӶ�_H��jW��Z�\[����h�J�*���N�i�5k���CȬ���v_41�S#>���ޤ�ۗ�m� �]@�+��o�M����ﳗ�(X�5���9�W�vK��V�_lGjv̑�w��v{�0m�w�����$6��uOpZ��W�e��܇�S�
�{����no�&�9��f�o|������M���٣7��{.{#����VÇ�pn�7����M~��\�?�o�FXtHGG��He�m���&� �y�D՝ڗ�3p��vɌ�y'%O�����a�ޘ����f�k���^Zk{f�����#�9�~s>�G�H\�^C6.���Ϊ��B�9��N �'Q!��=Q�8M�iG�P�L<�� ����[��dZ�b$D���늍��{��A\��h��T������������X^��x�c-��y� f��k�=�]@����=^c��q�9��1s�du3�L����њ[P�n^;���Y�[����rJ]ø�d�f�L�sZN�&�*�wr�_gg��>���l��
paǌZ�h���!縐�e���s7��������V��X4X/Q��F�]Vfw�9�]%3�_m��߻�v�ބE�$Ϭ�C�I��~w�����;���S�W�������G"�
��@D_������	Aߟ��<3���L��2�ȳ*�0,��*̋2��+0�0,ȳ̣2,ȳ(̫0,ȳ �2�³*�+00,4ȳ(̋0,���#0�ȳ�L0,��"�0,³
�2��2,��̋2��3�0,��2�ȳ(̋2,��
̋!"�+0,ȳ̫0,��"�L�L�0,�� ̣2,�°���"�2���
�+2�ʳ"��㇁��"̣0,���̫2,³ ��� CR�Eze�P0�� Ƞ�� �2"0�2��2�0"0�2�00�7�@�\z��Ua�� *�0�2����� ʪ�*�R� d eUa�U�  � �UV@UXeUa�0�UXe eUa� !�U�  �QfU�`XteY�	�f�FdY�	�fU�OfU�`Y�f &�V`Y�aӁfE�V`Y�f &�V`Y���?��Ǜ��|*�(��L 2_�ݿ���z����{og��oA?�߫��������iloc��N0s��t^�y�~�PW��?����� ������_��#���?��8���	�%�i���?z�
 *��������q%�@����?k�A��=���h~A�X��>�"��)" !B("� �D�!�(! ��  HJ�����,���
�(ª° "H � "J���������� 2� ~I ������_���~	��DQ�h
Z��p�?���������~�_�� *���?����O��sП��#����_�'��~�����(~��~�{:��܀�*�@_������������>���>��*�?���t��>�0�o�����$�r{z<@x�( �}O����C���}����������?G�?w�~!������$�O��C�@_>��D� U�׀��|��)?R��&? ,�������?����a'��� U�j�=>�ԙ��@}ޠ������k�AU������
��l�����/�2�?�b��L��[]o��� � ���fO� ĉ7|���@$IB��	
��TTU��IU"���E  AJ��I*TID(��R�	D�J���D��Uh2)f��mmj��"D��JIJRR6�m��UJ"Zb�Ȋ"DQT����6�TJB�J֑J�J��� f}�;)Sf�m�a)6҅��1Q�6d *+fQ%�Z� fЦ�)"J���kH�!IA��0Q	M�Uh¡B�R��  ��g�ۺ���t�5�ݺ���vt��v��5.n�ګ]�V�w;�ֹ�(u*wm�
�n���[Wh�c\�A����+�6��\ڹ���.�R��X�$$��`h�W�  X�{
(Q&�&��+�/m��7�������X֝R��m�1"��y��և��l��V�jN�4;i[]чb�v]v�v�ն�εr��+V�seګT�m���:ۻ���R��%P�EA*�  q�H�˹�]�jݮa�8�w[�6��\�lwn���9]NΕZV-�wZ*�iWs�m5��m�H��ځ���wm,.����ln�n�Eh�ݨU6m�J[4R��*$�  =�r�K�n�e
:����]�wV�b����m�ۺ٨4&�g\���ZUۊ�v�J:��ͳ&۸�t�-��;�Z�qu�J�*�J6j�J+l��  ݭ�� ��ͥ+�.WV�l�gu���U����Vwn��SW*-�9v�M��Qָ�.�[�VB�Q�Z���*�ac�D��i������  ����wd�ζ��v*��t6�Ꙏ�s�裴j;[:�V*�u�3���v���l�ͮ�(�4��]kZ�2�*�� �4��JD��   a���]7Z΅��jSn�h�uk����i�q�һw:�Pv�ki�:��@m�p: ܇  50  ��P��@��KF���  �x@�S  �L �b` D�  �����  P�ݸ( ݲ��h����N�@5��
@B��   .�  ۣp  3J�  �X�  6�8  �� ���� 
��  �4h
kN�
 hY'cV�*H�J�P�h�   X���s�� �@0 ���@ܮ t�4� r���A` Y��  ���&d�TC 4hE=�	)*P���2�d  O��)F  �~Bl�)P   ��)
cUJ � Ğ��H��l�$nTP��Pa@ъn@�x6���vE�~pجEc[���������������*�j��򵵶���նխ����j���z�j�ٶ�����������$k�1Jg���j�<T�@В�]ڕ���e҉I�f��(Z?����f�"ĺ5y�������A�B
Ӡ+�2�5�H�C0�嚱�c��@ƌw1BN�v�b��(�X0KͶ­�t͔o,��1&�l�J������3wi�ɩMxKŠ�ۙ7)�tK�{��*���8��jf�$*Vŀ���uf}�Jۛ&d�j\�i�"�z,��Z�ݛ����M-�z\�2ywP����U�S��Dk���kh��{����]ւʰȱ�Ĵ��84؅�#��u�If�#Gl^d��d5w2<;�ȥV�<h귱U������\�[N��r�R�)�Z`Rx(a�A����Kv`sAS+"�JhlA�6VN!�S0�K�f��v*&�M�Iݬlnm�ЕXY�2@���p:�8S�5f���J�&�MVf ���.�NU����z*5�*F��;Yc6�D1_����eຘ��4Ih:U15�^Q߃��&?��1mkG	AMQE�w�n$�;Su4�jU=H�z���fU�3hn`�m�EL�$iqL���I�Рw(�{x�m��d%�B�ʌ�y�'�@�o"v����G(Z�eV�w�.�nS Q*1�+*ںz���R���o&a�o!N�Y�>wW���q��m��6�+�۱3"x$&r���K�Pxd��`�� u��1�.΢�'"ou�5�+Y���n�N\(c���ZV�2�իݲ��cY/CD<�{�V�U���7x��;�Mh�L�j�r�YP�05@�����e�&Vm�E0*L�Fo%&�jHУ�$4
���n�#CE�b��ʫ��
!�X���#n��{f(,D�T�l#��iP�X3z��4ӽ	�HP�wz�J�K1����E�h�J:�w���Jn�Й	pk��(�k�)�G^d���*v��ZI�a�W����:�����l:GI�6��A��k-�X4�T�k�iܱsD����V�m�'�L�L�+�Q ̗�}�K��F�(�e�AK�A���,)
R�l%�ݪ��`���&�1m��Ȕݠ�)�K噣650� ���PwVw7eu$���ԑ8
Xe�Ype^�]��e㰘�t��`��#G��V|��]أ����(=Rn�j�����<�q6.���mw{�"eP��YH�I����J�v�a[��$�f�jc��%;6"���Lٰ*���,La�,,�t�h��lS.��^˭)ب6I�H����J��WZ3%2��ƌׂ�b@^�p���tr
ڶk(PgZm�Hȫ�sL;f�%���F�7�&����%zf��YJ�w�Bm��-a�P�e㛺5�2b�$}�-T��Tx��%�D�n��x�ڻ
��E���i7�KԬ���X��yn��`������DX��@٨D3h�Fѕ���A�X�j	ڨf�,�-6H�V�":T]Xsr����]#hM���Ͳ�F�M�
b���N*9�X�S�b�٬-YzV�S�V�m��k�ku��Z�mKi�cU�Z޷��,�D2b{5�-٫%�[jUڗ(�V@�+K �YCFAI�U�8��nO������b���e�G\a�5y��XIa����x�/���׷3[��\���n�GN�[%f�U)2ʤ]K�ZV��U�&\��
&h�ݙ�X�oI���fn}h)4EI��˭��Ӧ��ҕd�wi��bX"#j�b�x�Zb�Tk5���A��V��Q��K(�0�mfPJ:ԳK�.�0��uj��cv0�8dL)��(�UƉ�k0f��T���',�,i� k4:*m^j��i�V�j����ƫa-`x�6h�{u���INn��p�N�.�Ri��W�����l��[�)0����&A���sm�:�5�q�hJ�$�,@�/PӺ��kJ��Yl�6��XJ�(�l�b�J����MS�Z����@���2��6�Hnc!/rF��u���2��Vc��,��$��k�І����bTB���6�+nAD�gUd�xޛ�'Z�)P����5k&�����z`	Նu��Ҹܷr�L�W,c=�
�y�.WP��M[����ґlX��i�Y�U�j�|(iHfT��Q�e��LҊ���n*�QmJ�MU�(-�P��F�le�i/o :`e^Mxb��A�*նbrۙ2�4�.�\�-�e��ҵEy�낷5���X�(��ĉ����n�,cKr�|j�t\/��t��K���c7#zS�C4��X��@�8�B):��TO6��[��t�,�EP��5)��YF�� A��Sw2��©�M����.�c�Ƽ[�ƕ��Fr=zj����й(��%
�3v�R�򴕆��VέT����ێ�j���F���0,ϓ�Ϩ�flS�J�Ջ{>�^8�vWr�&6�m�0+v�#z�n̕i�ъn��Vc�(t���	@+��ّ��Ry/e�	L��T��;L��c,L�����M3�sr%�+4�ǘC;*^c�Ni���p]J���$y`O���o/wv�w�.���+����'t�	f�K,�ֆ7c�	jw���R�lh�MlR�245�ц����$�hbȎ�M���j������I��k��:ޢ��-��b�@�A�ځӰnRMFV7un�kR���6\ј�7L�򝌼�����amۛ�,�M���LA��U�@ԇN�d��Ur\��������E��:��Bj�YM�y����r�ܘ*P̀�&&��L�jf�k"�|$WQ��[�Q�(JtVӕm��[�J\�[�D2`��:���iL�-�S��,r�V:4��/+��.}�mL�ʷ,����b%���هb����lZwJnKG{���$"3)�Ϡ���ώꗅ奥����Sl�Dm�lQ]��W3	Z�@\����I���vʦMsHFc�f(s'd�raFa��2��1���#�涣��e<,���{�nV����IFK�p����LNe��E��x0�ʚ�=�ȋ]Vn�w%�H��]75��[5�����!j�V�KG~Ci]-����囄�j1��ɭ؁A���G��e�V��aw�V�v��.윬ܧ�NI`Sٛ�ɅS�*�1DN1虮���t�f[yf���[)����uiPm�Mh�����Ymk���B|���� e�ZtGY��wbƊL���Z̗��,�)c[V�0^�m��sp:����e7�##A�qDilͨ.\ϵ'�	���iM��5b�@��1lY(:��x��6�Ŷ��ۑn)4L@C�ķ�iI
�o*Q���E �
����A�5�/�1���n�fY&�V���S�4sfS�wq�6h���B\�rѩ�0҃Vi��T��/�)��~�9-W*�B-cDӕ�nf��1D$��m"si�"+l^}f��EvT
��:Ķ'�jݻP�YJ�i9�����ą`e�ę�ł��՚(���]+ۘH\at#b�q�wq�yA(�:��X�I����evA��5Xiҗ,�`	V��8���3*E�<7�Z;l*��h��Bp%I@r=ǲ`��V��[sV�eKJ�V�S�w�B̭*ՉhL�i�� ;�Vi�%+�2�p]Ve�jm)]Ԭ��gR�B(���m2��2dy�
�X&]��
\���;hV-^��n��1���X�5R�(j�rA�R��P9��~l�c�����Qf�m!��U�S�nAZV��b��nl��F6Lz���):�$vc,̫F�}v�"*՗%F�a���+̐nҘ"�[�Iu�(�!w�#&7-��N�]KlHh���c	�J�+-
��4���{á�@�x������s%ӈ�Q�d�s��6f�--��-S���6�3&[�mie7EX�H�569�0��2�嵩�hU�dSt9):��kM!O~��2P�PiU�V!m<�7N氈��љP��ԭȣ��ԩf��q�5ylAB(�ԉ7[��@�u�hvJ�6��q9ۂ�$�m�d�%��[y
a���5�7.��j�ZZ���Lm�?ku�!,����8���.�Ԑ���=95�f��Wd�[{��7�Q�t��4L 32ً#�J�N]��F����*�)��߯&�z�É��	{m�*���6��]YD݆�n�"\֡��0;�e��n��q����� �P�y5�c85y�ٻ��6ؚ�0����JE;������zb�B��]�[��h�ڋ(<?h���(�j�L�j��
ܪ��*Rl��f�h�t�15��˙XX�·���76&Z*�՟X� �DLգj쑢�5��~*��+k,K�0��	U�ںTE+!ʗnc.�I�{yӕ�,KkQ���q<�N�)fR蚴T΃���D�¯6R��m�d�j�V=�����@�f�D�|Uj�i�ӈ��z�<���2V,����GD�U$
�V����ӹa<�"��e��b;��n�f]&͓�z���x�^�Jc�7Y�X_f�Xؠ�&bx��A�t	�1��(oc����d+J�����Z��$�O��������uwiSTt��
@X��"���Ex�w�a�C6onn���Z��f�[�����w�5P2Y��S���q�:[�pC*P*���3<��*�X6	n!���]ۀ�#4�H�M4��b���.�!� E�LT2Q�Pљ�Sv��ee�u��X/��g�(�/5��J��J6�(c�Z�X
aX˫���M�M�h����G���N�oC66�Øv��4�+�Ϊ�+&���%�Fi���f��yik0�Ss�yZ7j�)�ndA��-f��G�˹[l*����hd��d4��6�X%�2C��(���$��̣hif��"�!ną7O&͹I��ֺ���*�s4-�ZPY�jG'nP���wa�[������Y��#�+�4�#��5qR�5��Tub�:WH,����!��AJ���4%��W�V�q�H�ׇ��M2/�IZ��=ڽŕ��gbS{J���8j�L)yak�J��U�ONpP��{��7�mǍ)m��*��j����j̚��p��:V���xj�I��t�MDi��2!�F�y%%07$X5�㒣*�J0���&��ʇ`�̎�M�KZX���:��pYJ�Tz�,5��+R-u�]#�t�V�M��6�e�RKo7E�aXnY��z�����5���m�i͊��6e1`�M�W��z����f]9��Zv6fFMaN�4��Uy�4թ�����kA�M���UkF�ګ��t�3nV�6&���׬G�LB]�4Cb�[X�P��5Z��S*��GQ�ɕb3L��9�c F�M�Vp�z�hl�XI�2K0$UF�l<���0E�)5of�eJ��]e�,
�o\�
{��ە�'bʘw/(Q�b�*֚�5*H��W��<��0�z�.�l���M�2��,b*@K`=����+�
�i��,qhVh���4�}R��u��m=K
�\Ϳ��B�1[8���9z�:j`�F�EQ�YqT&2����FL��ե���X��J�Z�[�ދ�o*�L����\����j�٬�@�Ѱ�.V ��0�I۽�����9*S���V
1���֗�dJn$�ժ�tmm�fe� �!V�K�bR�F���)�I�j\��Y&6��G�V �7k;��"+3/2,�7y�B��T�|����֕W������#jأ���ل�=�.b6�c�z��IK�ۡWC^*��D'ƕ��:T�Vb�Kn�-�[PV���H�u-�ǩ�Y4��պ�m���q��X��9ieD�L�f��8����G)&��Af2���jI0|\Q�ZͩL�F[NcW��R��)JZ�8,�a�N��m�M��f�߲�@���մ5Q�M��^ڍ�l��^T:B��ob���ϑ'^XWt,E��Y��I�bv�#�2���¦�[�Zf��+�o�o4GGK�Ǹ]�����iP��z�W**�������46�RՕ�jG��yj�	���kd�������j���\�+�^���̔�4�8�yE
54%a�WSR���KsNMK�`�R�Ԛ�&T?0㢄����f�sf�+�*�bYn<�6�L�!cE]Vn�b̀ᒢ2=y�X��RA6��fiʓ#�x\�Z3*m�6`@'�5�E���GrK�%��j�m/��%%VcF*�D���f޸�h�d�5�j˶)�zN���HeP2L�WIь��	��6��,w����{7�4.� ��7�0d�2@:��_J)$�ܨ?m�6��ťD�B��J"Rŗ,�̚�^*�'XwUf
0��� ��7s\�.]j*�>�#�Z-勏��2Ҋ�ud��L}h
Ae-�(Sku�e������1��&�k�i�Z�$�gf���R",�C���N��q��-���{b�VnlB|�m��:`�6�5��g�
s�VO��Q��|żzh����(��R�hӕ J�͍u #�I��R<�L:�I Ԡ)��o.bc�]� ۷aT32�v�d�Yx�Lz�A�]n�7�����*$�h���41�C0*H�ئ�S"y��:����̭$�>,��.=�X�R�Z&��V�K�ON�p��mmMIVf�u��[����6�ӊ'r���ޅ�M�M9�4��7x���˶n��ں��V�x1:���4�*f�4���E!T��#���t�Y���'7�v�'w��v5�����^�k*�b�r�i�{aŮ�/�����;���z�����n ��-reݮ���X@wM�޻�O9]��~\G,]+{���� ��ȶ�;9�Z�]�۠����?���'3D��v���1݌ED�v��];0����i��z�W
F8�+z�7�K?`�dҟ\׈�f{$��+���Q}׎>�h����t�f�[#aI�*�;-q*ܽ��<���W�sJ9ǀB���ݑ^��rΞ� ��_j}O�:X�M.�<�(H)�LF$�y�R�uy�K��,E��1�+�6@�[�fAeuG|�X%�RN�qd^-����2���	�J>n����̞��^��Oȇ>N;�8il��������!�Y��xPz�Q�-�`����wv���w��pd�D&�f�t��Y�&���s�5��y4��R��s��IԐ��\ý}�I��:[��
��ނ�t�לLѬ�Y�^+�3I�i��y!M��/T�HF�����Hik+Qna�,f��
���]{�]�q�as�s���۷���ܜ�k��j.#�í�iO�R�q�T�h<�Z�����!r�s�ǏN�Pȏڊ�u���	�VaϜd?��k*TT�As��x2�ZC��Υ�Ra�\�ݎ��ۆ�p`e��x9d��a؆Ṫj{�y�eA1����U��G�P��\�K�����ż\>�`׳��r���]nP`
@Wk��5��E]=����/�KS�]Tw�9����d��s}\��]�of�XOSG�j��Bvt�ܲ��qu�r���x�
΀��4��f�3gl0k��?������M;z�+D�g&Q�y�����2�=��l�t��E:t�a*��)��x�H�"��:�*p�ٳqnYO��:�4�sF<���ǽ�谔�P�k�f�ُ3��Rھ��E/F��Y�s(cO�tu��>��=w`��wz"ν�}����8.��F�f�����0�梏�!d^x敽��Y�2^%���N��zzmG��+��Q�[+��ͮ�X~�[$�~j�#U�%yR��ڗ�7UG���
��@8,=���c7����M��&���[n'���F��E��ͺOdW��WҠ>;-6ֹ(�k�𠃡p�Z��Cr���W+�ɸP�#H�v��f1ۅ^�\0f�����W����_P��G�woO�{���f��Vn�.�EP��ﯫ���u�粤�L[��eXN��f^)���*�<e�m��˓e���r��Juf��ɽ�3�R��܌e�^�J����}���u�Hc�4�qѣ#�NQ�v;/m�PS�v�+���J�f=��}M�l^aB�p�R`+]����V�m�"�z�I��6�%W�.���1j��.�{(Tw��3K--�W�{8�62�[�uwH!��ͤ��H�`�-��Vg},���bn�z�f-��u"�9i�oq����j>��Д�Ph��4��U.��.D8#̒�b�!���-\���r�\��n8ż�4���.���u8&��}%u>�scb�<Y�#&�l�WK���1��>�U��dZE���YYH�0�x>U��G��M���F�x��J�}���v���;TH����S�6z� �g3�t���w�QoeG��B�V:�*�QryZz��,��Ϻ�]]*c5z�w���Y,e��Z�#�D�*�r��{M]��j��tx����-�#YG!(�خ[Z�Lu��8�Ϟt��A�j�.�Db���kU(F:<iquk��5^V3����]�wlpߤI��Kj�3]-���G,ցF�a�}�A���C�]ѷ%���.c��(<��9���N�byN��59<+@���0�̨��!)ܗ�O�WI�_<廤�ܹ��%��/.���g^�g�.R����8�ގ�ӟ�K���!-�/R��\���}k�-���'Bp��]��5�a����q�{��ֵ�w��Nc8e�_�{���,���ܡY��
�3���\/�`ܾ+i�J��/c���^�N��\y�%�j���
�1���@�{g��Y���D-5J�^e����z��^���8�Vs��R&����EeCnb�e6fVs�-���+��P�RJհ�7�$F�K`�i����| �x_�ٻB����=�X��:�χ!IP����1�yZ$9�'�|)<u����YvaU;d٣��[dҗQ�+wȔr�����Ŕa�hqGɴkb�-�r닥ugj���V�2�+{�"�rɒ�u�Y�yV�	N��;��T2��A��>ߴV־��A�[;��l�t��bU�|�O�=�P���b�Z��������J��-s�[��.�/%%J�3�V�wR�j�0kuݯ���'�].�y�)�j�$��&�k��f�sq�$��Pږ`�Qt@�ˋQ�;��"w{�btP��zs�4��p��6�����6�#zV��4�%j�Nm+MC��k�Uv�L����i�1K8E��|b�Ǫ�L��v_.��&]p�5��ln�HOv۬͸E& IU�ƻ� c/��p���R^i���V87�F�/]�̢X=�X׎[�a��W�a����]E L���!|�h�7SEr�o��I*������;9Ab����.� Õ�9��������Xlǘ�߬��״�Wщ0�&فYl���j��e���5����h}�3k����ʹ���9�J�TKw8H �k�����;��Mi_ep�{I=���^Iz���0�"�h��m�`����,�b{���ף��)r�~qp��yx��WWdԫ�����%4��պwY�Q�-�u��� ��[U�C�p�e2�n�:��sfm�2F]���)D*6����2�CA�
�<l����/	sү#� ��JQ�a]Ѯ�>����;���@)A��7��܊UN4^�1k�}1γ��Bnb�X�M���Yd���{z�ˇ���L�Le�s�S���/uC��JC�s��8�N�5��n!i���I�u��/9�K%%W�v��ᬭĲh���p�5VV��K�v��3؃ݾ|�35�n�♆�z��2詜`�l�n��*��>��V�W4��K,���FV�s�e��y*S��NVv���Iٸ�`W�:^vD�Z"m7�����B�68k�.����WA� ��ȭj��e�*�fq�Fм,�9�Y��SI�t+���L��]]h��� R�Q`�oMC]x�Y�O���ɔ���ùl��GL��]�`9��C�&�j�,�S��P����P��O�<l2�fe��R��A���S졦t��n���O��ѝ��Lj[˷kz
i��ູ ��ݩZhJ�tڶ��f��%�3n�*.��ry�Kh��9Jǚ���mV�1��W�Cť�p�@�1����h( 4-��)�G:Q��F]��u+z��eh�x�p	�0��O#���7��U��u�KvH�$~c6#��s��ӎo�]�ȵ��C�㺅*�������ѡK����o6�mf#A.W-Q�����nԻb���➤ءL��e�4�]��Y	��qh�F��S��!���̎Y��>���a�._Zb.�Zy��.�Eԭï�Moe�l_[��j�jÁ�*�k�3��͇e��ZÁ`���×,e^�{&�ij�v�z�8��/��얋w��`Mٮ�^����l��^��f�#�_6���Em8v[���%����!9D���!�i��eS�	6]c��fz��Zl�J���������TQ��,�{*�AeC�5ԛ��8$�;�����{�ܐ����}�u���[ɕ/`�kj�)��J��̍o���/a_@���V��'��ܺ��s��z����˾��C ��h�*����G��Y�Q�6�����S��wc��g��wX#��I��8#��w�A��)��:���ud��
>�ɫy[�c�\�#}�u5�3����앓]���I��mR�"�58��ӝ��_u��>�؁,�i�sWY{��N-Z�s�mY�W���q�qVjVc�����ƚ�R��*�i�l7��ƴX�m-�U��7��ϩYWYY`�I14>�"��<��d��@+ �Y�zq�@�Q�ڳ��̪ڜAӇ�s�Ӭ襜�*ݽ��7V��f��Ȣ�֧���^G�U��ӵ�SBwQ򖻔ݣ�=���15�f�c�0�{x�γYZ\O�0������R7�B����Ԧ��F�2�;�]7��LK�	Jt�?;�Ks9��[���p���)[ϊ#e��H�"�Ǹ�=�ɮ��#(�r�U��C.Ho�u"��7&���ʟo,�򮖸m�k1�;���V�Y���Xj���Owv���ֱW�s�0�����'%!CE	�xoI������4n!�*ܬM�i���p�]�:�ř(N���osQ�[�5D��۫Cw`��[�[�]��c�eI�$JƵ�$���7�[����x,z�b$�X��RP�Z2��J:Ko��'fkW�b�Xnc9a3��{���=X-uS�	j�P�Y�-ҙl��*�t�7KtrMW�:�3�kQ�5N��U���D���>AH�Q�n�O�j�M�Tl�3Y�ޒ�n���m.��cw�Ct4�1�W��B�bϒ�j�&���>e�0���]�"�f�oR��X�p���)�m�*b�n[t.d����Gu�ƶ�6�A��u���;�r�����T���	\�P[�����䠷V�<�&��u��%2�v�ow6�k�?c}�0sw��V�*/�7)�Ĩ<|�w�+��HXB�s,N|R��C�++Aq���b�88�Ѹ2��֛U������������"�O:̶��v��O�
%<��u+�+y7ĵz�P�pge�ԩ�R�X�t�����8*=��8S�����$2�ʴ�K��t�je_g�&<�z��o�D,���X,<'{����A����eG٢�����ns���b��aa�h�Sirkn�[�cI U���cZ�X+�ՙ˳R�?t��j�F<qǐ�eV�҅���G���hMc��y�+�d��N��o*e�/j`��t���W��,SF����f�nVɪ]�M��ϥ��6y�u#�T�e�����b�"�u�t��H���a�R�`�G�X��nB�̠��m��}]��"��b؋��͕\.��8Wn���[!u�Z�S�>[P��>b�Ύ��̬C�=�FU�q_ 2cF��8o3��7w��I4�Tn΂ˆWc�}Wf-Q�m;2�a�������9udZ���`�s9'����D.���}��eÆaǝ�җc��
��v�	�
4�*����A3����r'$|��r2Qit��2��me���a�)qE�z�*aDG|��&7�y{\�����hTt�]ѽ-�	�88E�H����:@<5�@Hy�W���t*KR�I�P�Ef�-V\G�M�J�MÍX9V�H(�u[�k��SU��A��S���;v+4
:���Mc�6���<���x���J�0�Ԣ�<o�V�%L�n�KgbY�o/pR�jF���a(WO�>�������
��9��,�Eie%/kQ������	�l��Υ�@;a���=(*e�kOe�BC�=W�9 �M�ٶ�}#�K�g"�����0���#쏞�[s3�f}��2�DHQ9��Ν�h�+�� �`�c��n�K��g,��('q��R�k�4s�
�W��(0.�r�|�MaU�c�$[F�Pj._����Wڵ]3�CR3~��%ed��vF���`������9p9l�=�����f��.� ]��B��,�o8�7y<����Z����Xz�9m@���}'R�$�#o�aoW[�ۨq,�a3 e�sv�sޒ�CQ�'n���v=eJX�ӵm� ӛ�$�.�Y�!#�+�١#��A��3�7��	Ao��Ǹ�)�R��>����5`^Wnu�J��u�QL��Y���Wc��wWӧu�K�8/E/�ĳ�b�c%��Vʜ��ee2������jOL��0��>�I6^4F?@�YO�PXiJ躎�0�sq�\�(��p��1�Xk�58�հ�۫����%�ov�v..Xºٮu��B�U�t^TG'+�n:�%sM"e4�L=!�ڡWQ������*Nγ}���C'K� ����n���8�]S�ݫ����»dy+6��^j3E���m�]�h!	˹e����;��K����7�u�@\�Dv�&��A��7�tR	)���T��cEm(#
�<W.aY�ݍa2L��\ry|qYo��Ӫ�1��'��n�gj�,K�&eHL�z҇��"�'X˔2�8��h ��n�{����K�l����:,�ҥl�޶u��!*$ę�X���=|�
������vN�R��T��0)Ӹotqa�s��⛙�����n_�6�QW﹋N���'U�(�&Bx� �����˺�U1���g�^��{�.��ሱ�Pߥ,�:������^[�_sn�5R�\�Mr�؟kF�L}�׬#G�ueX`��R��[`����� ;��ٛծ+�����u���Վ�L�p��{yc�΂�C|)�q'����;�]�q��M�s��̤�fRhY�����~�c[��y\��4���^�ܣ�أb�l��Ww�b��<�G�Bt]�d������.��-���e����؍M�<��v�^�)���^���y�!]��m%��g�t�4��x�yf+7�;���s���C]A�2�V+#=ظ�NL�G�i��ݼ1s��\k�����l��K5�Ƈ8�Ž�>�ע������{����6��3��E�Y���n���{س3���R͡նW_
����C�!a�'�K`��מK2�+�Kp�41��O�C�U�����*4�ɲ���?��|>�����}��G�}\���uyS9u���G�	�%5�xc\Ff�_>]��L�BĻ�ðe_L\�o�*v�q]F�s���׸�@lp�nq�u��-"�t�k��,hj��%.�ݷk��b���b�X�ڔ!zla���n�|�S�܃J��nާ|�^$������F�_ʅ��拡�Bڸc��/o�V�\t��b7�v�z}i
-պ�g*[Y�k[��c]�=ŷ:�)G�t�kZ�3�Hy)ȣXⶍ�s�G, <(�Q���c�|��J��[����=��`ֿl��;��A~Ĕ'{�ٷ4���F���hn=����S��3�0��t;.�]�[�����`�a�Ly���TEL��᭝�he�lt�kvj`��ӵW&�u	�eY{��ã���iΦ�%���N(S��W[��U��:U��� ��tU�k����t� �����fN��T9!���;�gV�v�fծ�*�mYȶ�����lӢ������7M_]1��Ө�3m�hZHv�p-V�x�S��n͢��=E>Գ/Q̣����cGC�啯��ah��S5mn���׻p*���2�ջ\�|+6�a�b}g�Ty|��q�F����W�֋t*�+G��]ku	#|�-[Xp��Gt��,�[&��;�a�PK1�Ƚ���K��v�7�X7���Rp�C[�s޲�Lqr3�N���2o��c��9hb��6���V�Tj5�Ӱ#ᴰ�����Vv�Zr��������P}z4��#�Y�Q3���ie�F�D��\��{��3
�ۭ%F:}1�9n�i�.��d���نۗR����j�W}SfDOJ��V'I1�śK��1.Z���<{Ϲː	֔7{C{bU#����n����Z�&�ʷekK�Ql�q.�;7t3��GI�Y���U�GG,�_�\�6Q��o{&�@C�I�j ��gƅ���p�V����*�4��oS�{-,� �����T�s��[w���R���rZ��nˉ_n&�h���N�t[*\��a���D������������'�X���ڇdۢ��*󔵐Y����c�k�uX������b��L�F@я{Z�!�jR�U�k:u�+����7��2DF'*_ ST8��ı��`(�`Am�*��
�����Ʊ���t;��#�ĻKC���[)���9j�<K�������}K�{)�����,��K��w�y���W&H��F�OI{� ��Țgs>D*ks*��m��g.1���5�@��r���QVGj/�3��正m�����6�J�t̪;pBJP �R��s'���iU�4j����0�Қ��j�Xź��>��t��.��"�v���z���n��=�׸�oyU��Cj�Y�tG�����1��N����!��c#U�沅X��8�o���k��/qo2�R�xCEٮ�؍`�ң���(vˁqb�9J��~f��(�&�Ӫ�e�,D���W(���X�ɽGy��iѳ��9G��V�^� /�dw�{�
D���N��7�]�.J/���9���]/dޘuYSzS/.�l����۔e���iLd�eʫ�C��u���_S�]��E�v�<�˹BW��BW,ptv��V�Ş�*�:��P����$gofl�r#]��>��=r��8xZx�����ƀcC��J	�WYi�m.���M�IPzNu<�2t&��$-�]�n,���h�hV�u����b�P)��m|ύ���V�xi�ڻK��G2h�o�Vչ �. �wi)�Bl�wo2@
��ӥ��'n�{O��G�����Ac����,u������������̨j�ن�㮞e���C�XU-�p�ᷛ�.�W�V����ݳ�b�*��K���q�e���YG�Ev5�!)C��*������];wO�l%�
��3�ӻ�.X�Q���f�
�l����.;Ԥ8�O	v��I���X���$�"8.�����
{`�]O��q��Էn�x��2pL���9e3�d���� �Eom �4-ꌄic,	�n#��u�r��Gv�7]����������5�+��=�~܊%K��,x,���34�9��,�պA�(汉�m��)n,N���ST"鑪�����*�Y�t���1FF��{�%n;8�Q�������sV8�lf�k����#�ޓ2��ދl�ꨐ@�33���{(e
[�[U���tC#ͷ�<���i�سX#��kE�3o�/�R���Pc�E�fj���j"��������@�YQ�N]��.��Q��Me��gL8�bu��<nâ+H[ɩ�o� ���ˬ��|�ͧ�-�5�xs~VkB"���ǚUZK4WQ��,t���̮H��>��nfK��wY�%^���@ǭ�1�jS��.�u�v��v,-\8(�������t﹭�5K�E,��I�چ��n���!j���[����x��q+�i����E)�5�:�����@�Kx�ziB�qt�S���V6�P )M[�WX�h%�Y���ݻ<H��c+����"�����m
�Y";��>�j
p�������˞�}XZ�#ۢ��J@�4pޭ���u �;��x�ҳ�;��$��a6hz��憼��!]8�:e3����/�yXoup�!�r&"�"r���������%����MRŁed��]�*k��\�1��P=��REK��j�Χ]�ف��պ�5�SFf�\`B��5,�Km�݋y�`@��_sJ$|�%X�x���%�=����j�b��`ж�Ex�kvc�U��sjmo,s���تsP�:�ڽz2���ۣu�9�.�|����b�홹r�R�0˴7�B����"���*3�L���'u�{+k8+�� [jiu.��Zii�wZ1�z��Pƻ�����!�Ԥn�"�$���e�̮��]��QIZXR"�;�C��'=�)L-��y�&��8��Ʌs,
�t� <�m��[���^u,��y�������D�&�]G�u��̖�^J�v$��=����-�v�)�mQ��OX0�-����V���U�Ӣ���S2^��a�ɸ]8j�*�V��r�����i�W\�:7�m[\�@*�䋁)�%"�XQ�ȱ���wu#��nq�ANb�6��g+�{R����d���霅��+)�M��9t�S�]eJ'Z"]�����%��gf]C525�{z��`�c�9���yU��2ts��*��C#��om�;�]�mֺ��
��$�)X���)��-	�8]�n�:�b�̺nG����qq��C���q��ʎ���bȂ�X��#7>�����TF�by��ٺ9Fz�I%���Q<#�h嗷E�x��N��
��_:�SC8�Ź��pemL��R5;�k��h�+l�L*Bs5�4.�=��R���ݎ�շݬ�@����yo�ȓ1ղP�#+��/��"3��.Y�����:�B�iһ���K;:�q�R�`�%eo�"�v�3�n�X��\���U�[<6�N�W�/U .�nm�k�K�&����`�X�Cҁ@S���^��j�nd¨�p���@��h��+L$��Dr���c"(����8�̧b�U-��t@�]�}1��g�WX��8��˔�UI��}"�&�3��hU�f�����)K�h�_3m��ֽ��7s��nT����Gp�K�D沧�.b�F�� ���b�MFV�븰�������m�Iѻt��l!R[X�
ɤ3��dH/��)ժ�S��	*��d�k��r-Zn���-��s+����S��'�`:yb����v�G���] ���	ԩ����y�%ekm���q����l��7lҺ�$Yw�Q��m8n'�e����2e�rww_V�F��n�P���Ncm���TRLN��=#պ�9ʁ�t��V`Z��������1�us^,�i�[�}!�&zc�q��Z�"�A�������d���ȪQO�����k��U��*rg� �����VU�+Ry��V�`�Xz�[a�=�4b��.Vu7ʖV�e\g�(�Z%�v�fZ�<Z��	��"'���!us^�m-F���c���m����)T#2���ٵ���v&���Ô�}÷���9%g�OI�*TWN���V���7�ę�A蔝fb{yۉX�G���Jn\|�X��|�ҰOg�e����~ݧc���b�w)�(>���1�a���(��Mƴ|���턩�͓�+�a�����*�:67�
Sww�+��I��'+��K]�j�}�^u�Y�>�l�Λ��+�-��-ڍ�WT��vU֨iST�If"�j����,��(���K�������6�kh�ޜK�1�h��.�p�v[�q%����CQ�-o��ɾk���:;=���V��4o9_U��gV��a���u��T%�m҃����^�sc�Ve�!}u��N[>�7��|M��O��3��qk��*��:����q7��IU_�v�F���|�����|��)���<���L������T��P�J�5�*]6��R��6�4��6)�9�a>��c73e�bL����IV�r�Scv�,�2�� ��r�1:��@�C1��l�kYw��lE�ܻ&�h�/D�b�6�M�:����.��kh�='Hq�c���a��Nh��dG��kw�N(5Y���6ja��h���@>u��3�wKql���X,��Y�j�� #�7f�J��F��W-d9���FM+��;7"\VU��H�.9�	"%ǟ_7hЩ�+7e���r�	��.��B��)ؒ��g1�.�^Z���mo0=���+��;�0�	�G�r�n8�Y
 ���2�TT3oҦ<u`8���$�B�������E��ں�󄓨⬧F��V���6�ٓ`�D8ak0ե��gV��e]� |����"�2+~Q��)b�w:�a�})v��ZM�)��Jc��^W\��/h�i�UاQ\/�pbN�k��e�� 
�/:cZ��fn�MV�թ�vA�6�x�ˊ�ձ���9}&*-gg>��̜��W������M"V�g���![b����!�qN+}��OW&M,kAT2v�V�+"Ƥ�2��tWS�p��V���CqVV$_��F��U���'�b�Y��p���ݓB����X���X��`����E�&�Z��[v�&���g-cΚ�}0�kYe���e�(y谯ub.b)��*�9�sB����T`�@�K��c3�U��:�[aB�6bPnB��Y�>5���W*�5�EN�����|�!-����az��ǡwۡ�A	M�gv���x�yv����R8�Lh���:�T�z�,o^�#�t|vnTǣ:XŴ���L���V%��S�+��*�,������� ws:�;=�i'MѶ�Gm�r: �ݵ��(� ��U�0�{�M_[²���u�9��m`Cv����j�- H��'����I*,ݹYǆ�ǺIfM|�WR=�Eؒ��O���㿻��F�0v�mm����5�BV,'w�Q�O4K`Ս�yz�
�0�.��룒l.�4S�E!B`ʄ5�:���V9P��u���,{u-<�����q�n�.([wu��j�m:k"���X����,�뵱�]��p�KU��oD<Y��:���r�]ǲ)I�!9�ܩ�m��7.
xw��l
���HvZ�Ɲ�Ħwŵ��r����0��v.j>���nR�f�2��m�ѭl�%�Lܾۤ-���X'I�X-+�Jd4{\)W�����k6��z�J�."u���?�IL�g� W���~Xپ�ݷ����H��ƫh�n��&��\�X�k�C.�6�|̓����W�&�{2�7� (heh@�RG�����X�Ny�tޣn�M6�g*�Kc������M=�X�Q��e�H��\{Uػz�k�oV8G�9Q�gw�+Ic2�,D'akHj7%eaӎ���.dE���u�~#K�+y�gA�-�:��v�N9O��VPy\�+E�����^#����֍���ło�i/�e��J�5Xi�Ǽ.à*�5ژz/�T�)���Dk�B���/FJ�\���eMf�yfTy�r�%v��u����Жmd��<�4Q	"�QO�8�ǧ\�h<�2W�B���k�1�x2cV& �E�+Tc2�;���3�^3�G�]&�[���D��G;/+�|�G�\��C�;uYU��v�֝�-m���%�]nvu��"B(р�0bm,ث�wu���i��x�>qQ�P6�oRǎ�//8o`S]��������h$K�:�켁X�o��Eu�]��u s5n+C&Zw��BeՆ%9��n�fF�ze�ϸK֭����Q-�HY����ʾu��f��q�wYS:.v;�*ð���Y���\T릚.8q�V��isX��e;Ɗb���j�p�A�DC;~������<���̍�]��\{t=h�-�6mf���XN- :��rfŗ�*7@$r�t��� �reȤVk1��m�������˝f&,���]E��+k+ ݮaҜ�M�n��Ts��0���|��ł녹��9�����Д��t�aL��B5UѾ��$*�-7�k�i�^�i�/86r��Յ{���4��̛$��z��3h��=R�{Za܆�U.���F����Z�g.T���ثl�����*Gv�i��!��,�.�V����*ƈe��(}��q۳�n�U�#���� 5Y̫ت�S��4��.�99�f�L\�n���x��4�����諭���}���W�^�}�<�U��TޮT�����yZ���L�7��m2�ްl����\�6����v#f��e�n�}�k;�|2w5�n��P�N�\OR�oPA�-z��Tp�R�[`9��m�-g��,Wi��Չ�^}��V��o>k	ַ����eAr���Qh�=�W+����Dt�$� �9;��Z�>ǒhh�I0�`]n^��ޣ��Nt�XhF��ՙZ�i5K�1��x��!R��Tq�η&�k��q��\0D����A=�:X�0��}��yO-D�X�b����L=�}Bݱ�U����V-��;0Z2j�;w�-�O_�*�o��+�h)w"��3>�fR?Nov���K��87:�WS!�:e1�ni�m�7z�1�n�|��W��4,e���AǂVC�,�״͓���kCh������j�YK�[cM�G&�Wb_k�����ڱJ{n�Nr|��F٫��$��i\� ����hb�3��ȳ�i��s ,�$�F�S6�iҺ�䓶��1]��lWN.}7=@���:��5�D����:�Yt2��x�,���RN����IP=�H�D��V����L�]�ٗ��Q�[]V��|�䭃��o�L�5�3hf�v�R�b,�a���P:0�;�i�;Cmۡ)���]q������P�ܨ;J�VvC2�*p6�h�=u��".�w����Ci��(]3����GG9��	.:�ؗs��\��t��C�G]ۜ.ݎ�ѹ3r���̺h�q]�wnQp������n��ܻ�s��];wE�s�swus��wv#��n���$�BF�t���5̘�s��q�����q.�\tgwt�
e�.�0n��Dr��N�`E��݁�ݻ�ct�� 9�t��r�\3���w.\�K�D��N�sE��
��wwqr�9����M��r�gu�㸝�+�컷a���$a��۴��(�Np�.t�;4�ݛ.q��������P���Nc��ɛ���B�\�]�\���r�7uuΤF��7���c���ʉ*RC1AE����:\.��s�9ە$D�79X].�!\���w]��Y+���7�����מ�W.�Cٜ��sim���;Sb�!��ێ�_���y)�>,-ڡ!�o77N;wَ,��b����ox��+�����m�qR=�����Z͢�K�s��]�r�𻖩���H5��{�>���í���-\N�s��_o��~�y�{��J�7N�ڊ����s����yps�������o�A0��p�
Ќ\6_sQ�\ٽ �Q�-Z�����{Ԇ1	�����C>p�\}b�cڬD0�ZbC<�=G��~=@z�Jٯqd���^����'יLĮs;P�8�8�U�i�O̭�
�I{�|��=�:��} ��!g��L��_�)DÆ��2<�;�\K��z�}�6�V��X��a��r���_Z�;��Cq|Bޅ}'s�ി�s��Kc��C�H����靖ٵ�87]Wu�n��g��aA��_z�#B��NG|_�s��^�`連C�'�k����Ǎ*�θ�+v��s��3Ԗ}Fg&	��|^--���Im�*�4;>���h���W�R�Ӷ���Gͷ�}��.hi����+�g�aM0I���![⇃��Gkz�V'�[BL������$�l{H��Йa��[�2Q�	��`h�]�i�e�͗��9�7ٍ�q��[R�g�N�L����p��X��6mo9��t��f�9�n��R:[*w3w�Oj�M����s���
X��O�	�H�s\���ワ/<��U����p�3���q��|�(~���`�(�$��v�	]�˫[��e�_q~�xb䍭�}[
�zu��mW���3���7n�鿄��[��զ��}U¼A��Q]�ԅT��`�A��hd{0#�Ý2�Q!91�BN�ƫ��=�u�&�hj�k�A�����F�m���D�K���Xܒ�R6[Stm���s(�n�S�[ h�� ��E=\O��,��|{��o���[������6\c�_�3����ɪ��:ɢ��1��}b�3��f֊t< ����%4fW��l+ݢE\����}��Ý��ڬl�`�u�B}�_rW�P�;75�U��%�9B?)Z#��0*O�X}Ԝ<�(C\���թ�n�ϖ�������γ���ޖ ��Ofj
�E������OTƀ+��eXHT?nW�ڱ�#��k� Y�2��0�\��Y�'�(TYy�yW�4$�����w�*���/�e���?�_c�t�������j*��a�c�3����{�]����ո���:c6�h�a��+�{+��-�	�onW��W���e	k@[7ƭ���c/26T`s�˩��wh��!�o�K�D��}��m�(]�+C�\c#5e�������I̛{Ǹ�`���v�o*u8�}�gWu!��s^��z*o��^�F��:%��]������*����U�I0w������[����Z4	�A����z
NW�h_LQ�&��t�Қ^��0��y[Pxs�.��Rz�}���+�yO,����ݟ<C5SZBj��H�tWo����ײV��6*ǒ��no��t�(�����ä=��gU�_Cd3�t�{Q��"�<�G�J��#n �?��0�Ӑ��tߴH�r³^��J��І��XCV:y��ew�z�kj�ᾪ��9I���7��Iz�!��2�fǧ<�݁��\׆8��
����G��0X�e���}�|jĪR�4I�Q���IzV��n�#�].�~����߫Ϥ+��W�!��b!�啅l��N�!T�J5�]H�$	_ɑb�F��ᵞf���̾~��|<���&����Z���8��%���W'ćƆTR�����)_��=��J~"�o+4{�_-�3�v�g]��R���r�̱����Q.��;�pCQ����_�����Y�/�`/*W"V�f�s[e�Y�E<�JlF���� P��-�59r�^QL��V�J��6���M�9r9A3�]�T�js���N��I��3m�kAʁ�sѨo�lݹ{���|EX�ݢ��8Q@�ܝ,��~^�����½/�g������:�ˋ��5ܰ	����S8o ��4�ymÌ�rǾ��m�������U�:��8}x.��s,FǓ���,XTN;�1��ݻ7ɕ�T���k�
vt�tݡ�_EI��Χ,�w&q#��4O��rT-�;b�v�ãH}�H�t���hފ��W��O��Q��r���w�:s�ክR��K��^��(��^~x;î�r��gb}���^��^!���ٸ�t�]uִ=i�Zy}�������ؙ�t�^ڮ&`�c����.+��ܟ����b����Cw���G�3
uko3����T
ӂ4�EN*�aua{�������gN���M\Ǚ�YY�����S��f ���j�T��m`�g�t�aܻ�O�~���|�_5ojD�=~w�_��,ϝ�K�q�\��JXU�G��T�<���5��}�CݾB��K���ϗ�N�EŚ�{��>�k#'7�0Y:��D�t�'��X:dSҬ��&nW�(t5��E��f�@�FS��;��rW�df%nU0����d��wx�+z��o�,�k�;]�!?}c׾���ף/=�=:�ۖ�'�D�xI��}S�U����[|�e��w9k���>K{9P�S�5��+Տ`�M�T�e��͍�Ֆ�'[���mw+5>Q.g��p�a��#j-�#�i�R�#N�^d%�� Ο_!u7{������J�MZGrjǣ�_�vw(�7�#��xBn`�̳!)��*��M�V���Q�-�H�곂�X�a,4^���^�y�VY�1�J�?B*bY[}>˭��~��ѿPJ�g�m�t��J��F��woK��|y�}rK���`k)f��oƑ�(|f����\e������U\p�`��GEV�^a���1ϓ5�Z������iКKߟs�1�^�1/�X�:y��uw�z��Ǳ|i�$���kՅ������]�CN�M������z���7X#�Wzq��p=G�o�A��Sp������Q�[�~/���4��aH{R��M���9l߷;>�T;�g�p��h3LcڡU��-�W_�kY�CF�09Y��!d��d9�N��)qi{>nc7��|R�b=.q���Ռ�}����T��ά��S܌52?w��f�}��� E��n'f|�0<,W�7�x�};��)y��/��Z+�oǤoe�<x[Ѝ�#�F�J΂�=ˁ��gB{�����n�^T%\ׯ�w�<}���� �Z����Z*>Í��_lʾ��E�b����/���&�atʰv�>��.ޗj�b��*2�0�T��X�$��CB����¢�(+�Ei�����@�W����f%!_Yii�M{��d��Q�qH����������%E<V:�Y"��1\��[�}ܵ�\��t�+
��R՝0���m]�b��-����R�Tƻ�}�{��r�_���V$(�Im�U	�yؘ�D8��O}�t�ҿ@iq�V&�;zu����!�{p���l,x�(OFga�}G����ǧڭ2Õ����>���P[:<.�i�#
�Kz��� T�r��J����n��0�{��Ph=H��m>��ei���j�P䡞��t��wI��(ǣ�����������A�܈1�Ƶ!@S��e����zl�����]�;���bF��͎[qт��(�\#��pvLa�;+���5So�e����xug���q���t8������t.��Wx��%�&�ܥV�$��?	�`���T�z&uάg=SJI'5�Ǧ�픳���D����M܁��6д� �E�|�<p�\��'z�]�.�V���EԢ��G��&�ɢDOt2�OZmK"\�q�zsG�o�M���S�S�,o���w&�u�_<��66��َ�[)e�J;�Ԗ.嶗S�h��X��n�F�1s�-�;R���ᮧtT�\Ue�����\��g"���&�0}�}��x-3V��~��"��%gT3�,�Py@�WpN��,��ä��+̷�4!�pByxط/R7j���㏯���u����'cݞ8A�ƪn���l��g{Np���Ϧ}a!]u0��(�\nZ Vy�1#,�3�n��y�r\�g��^��J3)�~]��[�	5x��TUu��s���ä�x��Bq�h���.�{s�,p,u1�W,ט��(G�jt�!��l��R-rZ.|�YtV:�T���U{���v-f�)Mˊ��t�����c�|Y5�r�{�;>��.h{pu�sU����)$)&z�5Z`���vg��q�]7���v\�:��&+�k������^6ܶT�_f����!5w)�i���QxW�l�݂N�z�a�o8��g�����O�Ô-9��T6�����m�΃��}��&�4�$Y�Q$�V�E6���7M�u�S~�"��,x_�z�1�r<t��Ry[o�6�%{����
>׎�>(�є :��K���2�f�ޜ�V�J��q0��,�_,h*�������P�m�΢ggܴ5ޏc�+29^����枬���s�#'�=�1XZ)f���s�z�!AzG��^�݊�s���!���P�����y�+�o)���5�A0�50L�g#�w�Z]�w.+�6��8�+��e�7x>�w�d@����T�Xh������g���x.�	����ߩ�Y�W.�`�Q��yM�G�τ6|���o���Ђ�Jja]H�$	Frdz�^C�+g^�]��;�mM^."�4��w֟��O,乙~&��$n u��9��'A��}7޾�V�yu�4+�T��uQ�:��BÓ�Z��{�0X]
$.a�z�	ō�����M��_s�rk�Ճ~^�7�U�t�p�ޑ�3�� �V�ϯ,׬4��Y����>��cdiǉ�UU��?:^Wj��v��8����㏮���;�l���z���|�64����ySdhS������|e�]*��q�ҫb���\�2��˼B�Ȟh�B�}c���3���2�c���sF��Q��6i�B���c������w�+ͯ�1���dO�l�(��i����e��Go������4�٫�F�ĸ\PzQ�S]�z�����Y[�uS��|.��:ԡ2j��+\�X>�M��T�e�x�_�|.�t�F�����^V�&��]���&ՙ/eKO�v?�0����km�x,����|�p�*�iڭ$$vgJg"�`��ez]
���[��+k,�7ӳ�����y��cHe 5��خN���Z4��Ի������8gYmI-A�9�6%,(��]Ǖ�F�o����D�U��c�^8:�����T#�H�]i�����w�Cy��Q�bJ�{}mi�X���QZ�Jin�j�����~�ݚ|�����eXjmw�U��`��6��}}5e]ixRj�k�R¡�4&^�Ȧ��0.Y����W��[4ҎI޽(�����x�J�0&��;GpK����'n�<�NC��R*�D�j��Wos�=/U^�
�����$8�	�Hv3�����UC��]h�u='����w�z5�g&?����y���~�grީ�3I���e�
d�$1�py�ז�<߽3R���)"d�١qZ��#,;��?e}�m�=󖬲Z%o���E�Yթ߫�|֙|�|����m���
~B�i�V/*4/woK��v�}�I|�-s�y�˶Oe�rˣ��8���&��aA�Kl�3Vޱb����{C��{pB/���gk��9�=�]���J�.���偅�/U��ד<߬}�m���}��c���><�Ѿ����1��[0�����т�]n�e"ാJ4��#��3��Ur�h�M)�S(PoD�60�� �9rk�{���A��J��so�×θnJ��r�Ӹ�Pj��w;�|ڹN��Y�v5�哟f��\	+��d��h�ZXNQ�W��5]�&�˿#�l�n�� �a�J�p�F.+�k��&��[uM�:�f�}r�I�u9y�_�U�$�o���0Tͱ�V"�`�c�����{|�ۋ��(ѽ�Pd����R88��������y���J���"��ۊx��+-��f������%�Mv�*�*�x:q;2���� &/U�dz!Zw�M��W���f�Nj�P��=���e1q��:o�<��}��ZD���U��������)82�}U��9a��7ӗ]$ӹ^�_
ؼ�xm�+-�йp�G|A�����0uŴխ����+D�ח�`�M��kGi���^yPم-Snp6X���Im�U	��;��,=�G}�����J��!�����/����9��ys^:D;c9��W�k��O6�/�m�t���Ľ�s���M�ʫ�����|[:</��G#\�*�\~��Ds�0��Mc;���x�:�w�"gZ�SBjF���[�V���ϋ���a�J��>��v����תK�9qf���7�F�N8v��o�,�[���rJ��R�f\kC*K�*9�9�m�3�}o\�#�ԏ�����X"e:�S�����g\��k��q�����j��7:e�P��i�0�ϯa�O��������O:�V'Vo&C�h�^�ǀu��ޢ�]ut�c�z�7�5<�3��.�մC8�0��Iw^f�/	\��X�J|Vp�}a6L���}87-���3��Ĥ���n�ygF�u �ŔTÝnb�P9�ݶ��w��X��^JY/%6�����i��n镛l�R�V��2Z�
A_,;�dCo!����PV�vܱ���odm���-R���P"���K
1d��ǽ��̽�i�	o�]V0���"��Nأ�y
��"Jȵ��N���͖����
T8L���5��=���L�q�|�t��g@�`��hVu�д+X�@�3,�1�s���_[q��Ģ�Gڨ��A���{3~q9���m��]��e�h��vR8�����g&�ut)����ܜ�܃oS� ��M5�̬�Ȇt'�_�Y���{Ҡ��ݙ�����Ԅ�+W�k�/`K� �l�l�|�&�Vn9�W�7�́nM����t�	i��z!�V�xt��-��D�U�Hq����r�7W_rD.��k-o��k��oe�n�Z�J����g:��̀L��F\�Z�v�t0�-g���o)�(�6�Pu��&��.xw��#rq�����,0�)V[Gz�P
�|��"u�4�,r�d�3n�$FV7ҳw�ޙ�{͘�r�נ�vcP�l7��� �^�]�Wɲb�2q�Wz�!lZ��e�"����[ʶ-C:�-m����mg9����5���w�C'�(+5q��k���le���U��Yev�Ok��|1	��Ʃ���;�����(8Z���:��/̨���Q�������)R�.�Ν+3O,��'8I`�|�mr��P��,uA��,�K� h�J=����a��C���K7C�vy��}S�L��Z m}�	��V���b:&`�q��z�'�MbZ���Z��j;�8`҂�+���C,�<�@�� N0$��E�N?fV�ɪ���Wʗ�
�����GY����[z�\����E��:�R�uM��x�̩�.���z�gO�6�Md��2*��������c�=�1xr*f��A&��0����v���9�ѳ�������g�4 `�:�*���6�5��l<����e��r�I�:���$�An�F/xT--��'����E;U���*v���t�3\Zw��:�!q�jr�J���of�2�}bٳ�
�:����:'�f�v�k��E��B�J��"����knV���Ģq
�^�*��V���}P^��N��հ��z�&�����qV��u�5�׽�_뮙wq e�sr��9�MJ�uts��d��!�wq���J@!$�.vA��MwnXI��2MD�@17.č��2���H�\I�Nr\IG7" 3;��M4�)"��ЄEs�9CDbJ
 �c
H�;�� �77%w]�RIdRu�f�E,��##(wp��%
gu�$w\bg72d*$��K�r@�3��b]ܙ��&C�FC ؒ��w@�$�-;�Jr� �2ʆ]�K����;�� �n�r�%��H"��f3���]ۆsu4���P'�?
 M�Wgב
9�����o}h���K�u�u�̺SMC𛱌��OgJO̕75Ss�9��uWW#�e>:�������_�x׵��;^���h/_{^"�~�Ž_�^wlno��{�u�����|	�'����@ђ��I�����G*�C��{�޲~��Ȁ�߫�����"#��+;6ϺrD������h����o��b����/>���צ�6���������oKߝ��o�߭{��ux����:�7��~5�}[��o_�^7��k�������փ}�;S��Rf��k:�B��U�D��kO}_w��~�}^�x����>�m�ۼ��g����ssn��~���r�˛�^���ޕ�zW�x���ƍ&�ܷ���o��_�z�z��������{1IC��� ���]�o��>��@P��x�j��}���^��_��|���ߊ���}��꽭�\���������m�|������k������oJ�߭Ǯ����7��zZw�����ͽ(� ��'�p^�S�}c*;}C�#�oM��-��{����7�S߯��~7�����~y�7�ߏ�~|����ѿ��}�|k��^-�Ͼ�lE}^+��}�y�����ޟ�������m�x����݇歷}�"D_'�������;��̫׿�x.m�:��^��i���]ס�͹W�����o���6��^�|��{~6�x+������������ε���t.���F� �5�}��1#�>c�F"�DN���z�����J���=>��~u�~/k�^���/��[���k���ϗ�W����z��?������B����3��@�TG�?|�}�G[���������}���r�y���^i��DH��*�l�޶�fbJ�v*�j>w���|<hߟ�xޛr��y���~��j7��ok���Kwη�ޯM�^7��W��痥�+��=�:���������z[��[߯^W���x�~���RD1}}D��rTfzprڟx{S�k��}���DAsP��">��_��G����_q�� BI����[s_?���_����m��׋}o-���w��j����7�:�ߋ�ѿ[�c�X�,1#�>;�^.���y��������lEz_����5z������}[���/{������{o>��[�|��Š���޾o>�_��i���}��7�nm��~/K�oO�۾|������z�O�H���#�A�>��By��:�U�b��b�֎�uS� �KP���/�QOy�,�iw� 0|6n[{,�aza{�v'X�:T�2����H�B�q�/��1>xx��e��:��j\m�k��I�}�6����C�g��.�)6����o��w<}����vǶ�	���:!�G�~�!v����zZ=}�����x������okE��o��꽷���j����7/�x���//�|�龯�x�������-��/;d
?b*hG����~}���ݙ�O��o�}�b�����}}�h�'��ż���W�so���Ϳ׿Ϟ��a`�@?�#��� ���#�G�>P�} D1��"���>��"4G\��]�#�:��/�g��}c���LE���W+־����x����y�ү��s^������żW/w��U����x������i�}m�����߭�W��"+�����}������"���H��0a�4$��4�@�_�|��h����(&��7��=������ѿ�7u|^������EDW��޼�KO��ܽy��彿x�W�<�����y���?�y���|o\|�G�}�P�_�eP� &�g���(�}� }�������+��hC�k�߾^��W?[x������nW?���׵���szo�^�v�?��^�޼nm���x�}m�Er����ߍ�η��1>b�$G�C�1~8R�w�>��}��ţx��������W����}�oo濕�o���7��W,}_[y����_��ͻξW��>���깹|���|�\��rE���\�ЁGԆ�� �Ə��G��}�����حy�������z<E�?~��*��HdQ��i�*��+�x����^-���������[ڼj���W-�\��U�η�x�}_���kگ��7�����x��y_R}��C�W{��+~s=�YV�|ER�����~�m�mʽ޿|�M�[��n8���
������J��#�?3D}�߬~��7վ_}~�潷�����������^=��|���ޕ_�����7����� �W�5�I�s��Q~�c�#�>������xߞv�}�{��+�ѿn��{W�O��������6�����^�����~�z�E����ߟ�����W?7�����������?|��vo��wdKƧ�{}��PS�T�E���L}"Dp�V~��ȏ�9����?Y��H���Ƽ_�{��/KF�_�<��_��h�/]}[����^5����_�\��~�����/���o���?��o��-�\߾�*��k;<	�ԇ�_��ikZ���}yh�����H;��y�:!k�v�O(kt*LB�nPH�W}�_^���.Ի��[n�#�}��8�m�Zݜ�8��<�y����W9��Цu�U�z����ݵN,�.�A4rc�pZ�����(&#\[�|o~�䀿������`a���>�o�O�?|��4s�P�7�ܯ�|_��5�^��W�/��5�ϝk��_[���_��ѿ���o�{o���|����k��[��1&���(�H��z�f���=��}�����o���k�޽z׋��x��C�y}�"�Kx��|�G����/��ۖ�^דo��_�ſ��v���y��o��y��z�u�o���5�t��}��:[ID��}�����G�_}���~5��k��_��^U�lDEB�P�G�}��g�꾱�#�>�DN�~Z����y��������A~����5����|�:����ͻ���_W����>�U��xt^GA�
��3`�;�K~+����z^��ߍ��z~����u�z��޻��~�J��=yoM��w[��n��|@k��|��H���1�}1������o��^o��F�/��}�|_�8�D|�lL�FY��Ƿ����?Q�5�W���gήX���k�_���_7u�ߍ�[���^�z���o{ӯ���#��k��@u������" ��곣F����>����������-�}�8D��>���g��y�ٺ�vb���_��#� x�Ԭ��E�$`���zo�x�ϝ��\�㘴��}W�/<�?[{U���{��^�����M�#� #��ITxG�G�Ξ���h��>��e6lb"<��$�7�/So����o��+��+�{o����>E���������_�k���_��W��߽�o�^5����w��؄PH~"(�����t,���<G�x��~�������O�������I�/��,�j����#� /����}�">�}1z󯭼񯿝zU��������_��-��o��k��[��ux�����j��ޛ�wv�_���z�o���E���p�� ��ZDq�Q=�y���W�{LD��}�������F��Du������oK����r�W�U������V��_�������뺹c�|��ͽ��s|o���o��-�u�6�;��W�h"$A|��4{����oU��o�(W��-������ѣr���o����8�'� >�� v���D>���ﾷ�}W��ӝ���o��W���*�5�W5�}�꽭<�~/�z���>�
�b��&�?Z�&��(�0��4w�Ԯ7h�:_������}r���w(o�x�_��U�y?�.�'�ʈ=d����w:�mw*�,4����1mi��k��;L\��=����V�wω�,�0r�[N+{�2���Q[�TYIΘ:�~���k��o�ޕ����}����oʽ^�����~�M�>k��/so�����D}� ���ʾ�� G�>�ʼ-�]�ֹ�����ύx�W�������D�
��λ}�U����"o���؟<�K�^֞�{���7���?�woK�Ѿ�v�]ׯ޷�^-�Z>��5�H}>������@����W�_˗��?>�z�ޛr�Uϝ����נ}D���p$۳��ޯUfr�\�`�������m����~���__���-�ۻ�[������+����o�:�o���\���?�y}[���������k�_�������n~5��:�������c����܏�U��f�������޽���ž����nm��ʽ�}���U˛~<��뿼��^��nW˺��<hѹ_���W�ƿU����/����_�|�\߫��ޕ��#��cѻ�V^J�x��~
������o���?�}��V�~+�����|W���[����U�|~��W�������5���o7�׵x�?ݽ߿|�����r�\����g�#�R$� ~��)x}�����B�p�}u�2�t�������j-��������w��|�������Ƽo���~~�W�����_?߿=}WŠ��:��"8dǡ��\_*��Q�P4�]^>9�;�{��=M��S��-X�������x������uׅ����.^�w^v;r���gf�Q��E3^�mi�$����������k�<�&��2r�.u�{[����L����u:�ъ��ߓ��Y�ǹ�#�I�*�-��l�c�]���voݦ_jۦ��RU봏N�%=:���W[>j�ʷ#B�EĜ$o����+�b��.���\�̫��\��(�f���EX�����~~�l.��_`w�|=��z�k�������T3ޤ-��5*��Pr���p�Q^
eם:��<��F2J-J�茎?X%��׶hwgq�w�t���(�W��IwWNJ�*�5�6�Q�95��_SV�u��@2_���/F�O�V�P���KT��+x6	����ip�a4�k��9\=�:'�v=�T�Ӗ�W�Y�&s^}G�5��x!Į)��5�X7Bݱ[���O���O�|�$j�S聓��q�U�}M�ƾ-�c��k��g���/e/���qV�mcnUx��t�_N��%D&�mm>���"���gJ�_��N�����M}L(.�ޥ�v����4A���HP���d/�p�\_�%w�t�w�����Z��i ���&����`��M��`��W��F���ֲ�H�o��>��dN9o
��5���oMF70��n� �,	�T��l�~�Bdi�-�8>��]���R��3}t;V�Ϧ��z�_�ک�:ɣ&�~�V����Vֆ��<�w�����Ç�����^��8t�'�=�x	;2!�>���u^3�,�f�1ώ)��6�Ei���{eV<�z͆��S2Pw��>^�{��؝a	ڿ�{3��@-���|K����!_v>�����R��b��`,�^�+���<� Z�/%e+�H\�1[w� V��88�2�r*h��SSi]v��nN�C�v�Eg�F�T�!sZ��<��X�Cos0TE�#��1k�-J�8��Q+�.-�չ���GM����� ���W��ˡڬ��W��$��X㏗$<���e)FeK�{����{|��J�&/�{_έƄ����EWY�����I��-#�~��,�o'u�0����BD�#7����L�:�B�x	h!Pǵ.F�j�x��'�}]�-�k�P��\��.I�g��������ٵ��s%$���{�w2�����rK����,�R��Ӿ��^L�eY�n[*[��L^W[6���G��y��k��V|B���Eu��Adq�T���?Z��W������p��1z^���\˂�i���Ǫ]bp<+���4�I;U	��H�[A���X]��������VMR?k�̽|mA���8wQ�g�+˖&|r�VÙBU�ûX�
����.m�CL�\ZO|����»pq��|�����u -��	�G�� �J��Əs�n1�S-���)לk_R#�_�W���\��>��9�xMށp��I+O�5);����Y�z��m���& �hx�r�K|����3��ų� ��[ռ�{�ٍ-x�w�VîK&c�~6���G�����w3-�W	�uk\��4#��n��{)�2���'K��oGm�*X'�6��A���gS?z�B�1��	m4 ��7��=q6�A8��O�[^"��Q�;�Wrϵ4�ֽ�Fۘ��f�/B�_)�Hڀ���S���&����(�C�)U�b���g9=C>n��g]Ϻ��BÓ�3���:�]a�+���]Y��Պ�D�i;�-}���i��V%+��2��\3e��蓳,�����s�pw�,D�Sf�'�{��γѠ]b�:�Z����~t���z�W��g��᧖�?97�Ay�IIr&�f�n���t��:�'4����o�`�G1�O��q^�ڊokqd3[��NY�<7-�e*�>5K����k#��'�K��P�U��1�39�d��͕�<q��,K��h�}�1���L�rgo����k��tH�f����o����R���{�o׆b6sԕ���K��)�g�jP��C���9q^����t���I�ӚJE漏h��_��W+!��*T�qHEnV����-ØFh�nw y��[���+O�g}}l{���5���x~�V���e2������뎭ו�(��2�퉍]p��K�AbŞ5�-�cVZX��7���'Q��_u}�U*COՃ��K5{!μy�r�9X;�\y��x�m��gYa��=��<t7K�T���z�O�ن��%(R�{w�=�m:�Zי�>���L!�yD��;>�X*�K�^D�����4%�ڹ���թm*�^�u%~�+]kZ�ήů���v�3Vs�w��XZN�y�0�ܠ�>dm��������m�dq��L��xu��0V}Uŵ������N@���Ϝ�3_)�GҼ��H����^��Pg���q�+x��<��;e��grީT<nwX[\̙�uX޹�Oپb��I��5��;H�'Y�nX㾊���}���}��$M�;�3�w@�S�Q��6)��C_Ծ宓�J�r���|٦�"�Q�x>n���(���M�������~����D�C2���_x	N���҉� �3V.����v�mv>v��)���j�4Co}z=��6<�T',>��[�C���v����6��mX�fMhx�ez������1��n����U�-�����o��0<����� ��)�B� ��A?����E�"�ˋ�_rʇ<��&���,y��Hv!�I��)��S�cچWb垑���a�)�ݥv�X®�LN"X����~j��+N���Q�6�V!�%U��F��|�:�>�C�nҜ�S�5�2��LO�;8UQeuy3-�-��͊X7]Jz��e�J(�3�#�-4�`��Mi������ws�/��}}�;�n]l7u�@���c��.��x�/R��Rg���	�郏U;C�8�˜��mTK�l���Y�
�VU��!���ՀD	����B�*��J����i�
z���)՘��[��5�s�¥Ʒ��������{t�\�t���|qW?��--�0;�Vq�[��53����W���D�gS�����/=R���й�\I���TW?�k��E������}V�؍q���X}�'�]}�ھ�=�c�+��k+KebB��%��2��(x��fI���D����g�U�q�n��`���9� ��.k�"���8�E&�~��d��n奁���e��@BI�'���Xv�_zUg&�_���L��齒,��!���7�-�&O�s�3×4"W}��:��j�a݀��"R6��J��~�l��wL�]Y5H:[����𾢱U3�:�K���k��"*h�#�,&�|��Y�Uh�_W�pGn�'�|�r�׏��55PE	�=�n�1�rbV'u�9�g`��; ��V�yY�}��9�<����N\U���n���}\��j,4v�}{��F���zE��]+'^q�2��,�5P��H]D�Q�ڱ��W���7/x�O�[���P����� ���Hk���k��*�3rHR|ͅ��Rd��1��� ��trc6Wt��T�G�菢>�ue4ޗu��r�����5iX�W�������� a�5.�*j%��Frf��`Jϻn��eg�v�o��km`n��;����]���Z��d��=vY��v,�2�~��Z���̦mx��L`�]S[g��<%�pv�,M��"��K�0k��-*�;x��1uN�gث ��P�>4<e��+�����M�_�z����話�'��}7�T��V%�G�����omq[�Q-Ҿ�s��y��d���Em���y����*kZ�	��}V}��ok��n4$�W�(��.����Ec{וz���|�.��m��+Ҽ��A�rt�]!S����%�z�cζ���3�LG�čm����
�=T�|�W�[��FQ�h��2�+��Y5�2�"���<��h��ٵ��\���
�g��Vo���}vn��^��c]�li{UG��1��������Cr�R�}��Մ[����U5=�:�PA�]1�axd$D9T�����Qe�U�����7�>�����Б�srR8՛�^��4ȶ(ͻ,��E�.��v�$
Y�v�TWvF�NB|�vB�l��XT�>�w��#s9ݏ5��G��]�O�VmyJ��E�_fݬBg���o o3���U�S��e�]�/��c�(�=��L�uݨ�XF�Wf����e�5ƺ���|5-
,�r����Y�a�"M�M=Jǘ�y�.)��v�)�����R�"j�?H�d\�C1��k�N�TZ�4�ۺZLSGJDm�O!���;�k�Y7"B��a>v�}<֌�sC�Q�^&�	��7�д�En)٨(��&h��Q���.b�Xv��EV���-^�!1e#Z�.��ʃ\�j,yYʠ�PR��^T7Mt2�2���u9���r��%���ɶ{�p�:W9���+{�]��+Q��]9}z�yvv�#O�k3`j��̤^���:q��4>$�g!�Wbk��{7��wA��{uqշ�r;�cDt3L�6B
�)jt�N2:����ff�C��;���nj.� ����V�w[7Iֳn0�9yY.	��b�{�
�����pJ˻��go��/&�h��4]v>�V�=�\uq9�@F��F���ף^���6�+���)k	oػ8i����u�!<M ��`�G9���6]�d,�+�T�%o�Ŕ��XUܚ�z�U+/��K��>�V.��	��B�j�S�i��Ҏ4;�fh�ԅ�;N�oa����-W\�����Cs��	�����K-�R�����p��.�P�=��f�-���eg*��7�0ЮmӅ� �(�n��E��zi��;
��ip��MwB�d:q\�<������A�
����4qm�����ty�GnvLr��x��6;���',��1�v����<���	�nofK��w���΁�+je���g�7O����a�u��C��
�F����YJ�L2j!�]��[�ɏ�~�Ls�h�Իc�5zeiQ���d�$���'�e^L�=]:�bQ�RnwU�H�����L�9�ݐ윛��MZ�~�=����6u!W<�&z��iv3�&��5�{٨�[��N���୰+R�\��3iW���=�ID�v�*,�����n�
i^֌�h�{�K8�]��q+�Y��a�1�yġ�ٺ���S�)�����{n�;�ЗKb�t���ϳ5Y �Dgr����B��/�x��gH;a��V9�ILKT$�/�nM���N-[۷ׯ k{6�V�`�4Y��',T	2o)G�K��A�F����̣Wt�4ԝVg7�� �+w}��
���������jؓOg&Rʾ��\G	WB��O4N7�A��Ǣ��RF]м���>-�)WuNݎ��L�x�}]zbȯ6�m�x��ؠY��A�,\�g%����$*�����n�i�(������wA]�]`�@�pc�bmݽ�E�Bo�S7X<�\�q�0*$�H��d�.�hF$���u�d�'.&j;��b!31�PF�d�Lɻ�Ji��g:b��;��˦J.���4&�rD�19q���RDd�FQK�t�wGP
;�h��@�bK�أ�C&��Ś%�0�B��IK˗nt�v�.'M�Jg:�ۄ�B%��fI���DfL�L]5�n��$�A2Ҙ�@Swp�	c"��c&� ��`�uى]�H�Q��)s���	(�2HW;wA	��"���9t́�#���cb$�"��
V8l|l
�k]���tp_,"�r�������R	]���N��-�Y��,��u����O3��|�Un��
�����
�쐾'�Y����?^�����rI�
�4M�l-��χL���y�.�^��T�!���;�i�FL�����4csK�D*�&|r�V~�P���KԳ��<��ِ�O��%J��E_��x�0VT���ktN�ZY�A_]�V%R�mb���
��i��4�Uxs���P��?p��V=��9�"<���W��d��O+!zU%h���.��ߦ>�굳W�(��t�Ӻ�����|�`���.�r]�/�׮���c0>�v[�p�l���C�|R��1�k�q�`�OP��j͝t{�5H8�եJk�d�[�ꎷw��0+`[�]�%zK��u�-}���4�]��E|��^*���>����!\�~ǽ�XV�����5'�^ ��V>u���x�t-Wl�����{]y�U;��kvDH�x������7j��
�X����#��fqC���}�L=��O�<M���|g�1�J���o75��ҽϏ��Z��p��X*���T{-[?����ۨ���z"�\W��D�=�����+N��k���b�ܯ2߃�����yj�6����/����Y���n���5z�D���H��r��ڥXh��J,��d��XgU--/�'��n��ɋ�}-������M}#�}�]w�����X�M̓uBj:�@��?��꯾���'�P�E�?	��[�̜
>�왈���\?|�i2�υgm�m�zЂ\f�*��Oe�6�����y����I`�'픗3b5�{V�wau�O\�X2峙��mG��4�w�B�w�b�G���^+U�8�ʆ��T9��q�⠊��]XX��C#�-ZI��y�ڗIh��s�"~��z��?]E*�Q��QZ�F�錱���6�^y~�qjAׄm'�w�캎�j�S�eC������y:����&����|�+�>�Ée�}.���f{���?�|}w���~�-S����3<��=�2�Wʠ'kd �[Œ2X�t�3"����w�Y<�x��5ޗ�Z�:`��������Ө��;�g�We���>�".3��g�Y�Q4"�X��WJ��S�"}�V=����C�K5H�U��WF
yi���4s	0��� q�|�Ty%���Q|�υ�c���e�e��*5��ȑ�����h;j�p��+m��!�K���"�+U)n��'�{�Zz��ʍϛ�{��^{���bU0�=9���F��!�rE�Q����kx�Q�\>��wϏ9D��Ǭ���d�\�*ɒ��7j>R��3�>	�+����ZBݑq�)0��J]�V�R�'��n��x��mhR�Z,^]��j&N�����,�3�R�������7�;-+�E���u�Bj�/��_�W�~N�����r�[��]��Kz�}r)��ԵV�q�'�cͪ�7̀�e����V,<_��$쯦�>P[�٦5&7�͸4#}X� kVTb'6�����{�M����}sa�Yؐ5j[��
�g�^ب�U�"0�W^,y}��?���&������;>ϥP�!�I��)�t�1�Ml%[�<e�}ڷL�+���G�������Պ��-X�ճ�GG����	��^K]p����˕������cz�����pf�q��%��#*�*�<�ٔ�0<%Y��Pθq_5�~]��v�B�=��<�������Ӷ���n�ϱrR��KH��iF+m�\ڦ�r!M�����L�����{����>Z<3~V�_nF�ȸ���R|���V�HrkY�=G����wԇ��F��X���{��_j������܆
�|Z���+����i<��o�;ӶKWW4��L���ﮪ!�-�1Y�Y�&s^}G��>!�Om�{Άss��c��}���.72�:A�vt�"@��깩B�9�z{RC�a8;K�;�ʝ8n�5�ښ5��Vh�ͬ�'�=��IK��eNsN(c6���[W�����R]�\Fߧ��K�ؚ=IM�d��m��܈�`�Y�o5��v�ia�2��c+�F>�UU}_}�xѕ3ӵ�`�P���`���fld�~�*�3�����|[:<-�v��y���6�7��A�X�-_ ��`u"X7J+aݪ%}�MH�O�xE�'�[:G*�U�_������5�{����N��Ͻ݁5������ �`�&�-��e=U��&��녁��;Uۃ��_0#����B{�$'!�%s������Q�~+���E�V�� �-���������qf�\.V���L���4j2�*�&��Z�4�.URE=\Oۓ�.�*��*
��=��U�+-���x�!9z�n�Y��wKo��|����K��E���HsW}&����E$��L��2������Mβ���|Q�_wx��~ϼ�ݏ�G&�T�Pn�4T	�o,�"�g��K�a0�Ņ�n^�0ڇ�-�c÷K�t�y�W������EF�gs+�zo�m/f�q[�c�l�Ͻ�BR���Ҙ��֪��W=ϻ���nn��没��e�f}ֳ����>�����ГW�
�����ܯ����� mn��u�5	�����E�4Ʃ!Q�S�n�����b�U��v�ct;#�{��:s	�}h�(v64�z�{��?����=Q�܍��vpԇd(�t����;��RwndR��&���[e �فVW{z�_9\�����>�۹=:��u~a��y/~48�X��s�t$K>P�=�Kd>�2�S
���%�!�z�jU�{�̼��w�T��n�@H�j��.\���{N�c�=��4{��[�����<j3*�-x��^�Z{:�B�I�`�i�2�b�Ub������`2�[-�W��7���L��V�B+�(���8�|�puIk��l�0^wg���^�/��j�=���*�l>�%�Ζ;Z�r�g䓵P�)�����q�-z۸ӳ�{�{Ӕ>�ss<h�uC�w��ޣ���ŕ�b\���?t�@k�%�]p���ח�o�4�d\.b��u3�~]�k��.}C�}����j掻��JS$��W���Y	��ｧη޸�����`�o$�"<ՏF��s�E���;���~*w^�ǔ@�ݚ�����e�9��d��}�+�k�"d_��5�YS�ji��:�r�1u{��`��᚟^=�����C�C
��^���U�����M[:���f��^'��ګޑY˻t=��`Ƙgr�ǭ'%��9�a����pMe$bORܼOn��r@���Sި�����5�n�~"���ca�烹�i�w��Gm�������jJyw���o3���j��T�&�ח�vd��wgg&4�wu+��|>���%����Y�kb���<�S��Q/O��k�`�t�]X7��f�*�x˦8B�<��k<�n��m���L�r�&������H5�KR���c��$��cVWy�O7����E{U!�Ǫ勈�T�_�N�+|��g+����4)��m���w����=�Kx}2�g.R�q���������Z�= ��i��i��Q9q��\+�"�@�"�"�+6����{��vqX���xe4��x�bUK�t�]sT�dď3�ڿ�e�������76G>��u��*C\�F͓�K���O�l[\���ѓ(xj��r�`�}�̧#�wc���Wu���q�&{��f��!�UX*�C�U�X��b��W^���l2�\����6��g�_ ӅZ"ӗ��_[=
Ƅܪ��6�ӕNᤛCF�('#���`�6��U�~��������z���ӿ���b�5`5P��zW��^=����yV�Δ�ӹj�2�R��!�B�*�������18H��j�ܥ�	��)�/��ڧƧ�*��K."�+nf㔥$�NJ��N����멏&@���>V��7x`Y�B
o�3,R������KM��=_#/2#�/k늳Rf���T9�<^� ��х����U��\�Br,mm�Ϫ�����f��z�hq~G@T"Η�gޗ�Z��:`����Ϻ�ql.�]��>��*��z�p>��$��w�]�uEC�-u���
��7�ڜ��y���~��܇��R&���U:�%�����a�X+ݾtry�(>H򔾞��hR|��r��UǱs_on5�2���˞7�x���T��x*(�%W��J�*�T��P}����X<��i��ȏ��o�=�X�|׽Vk���ڹ\�?RJ�/��\O��u�E5�Q��.��[<[n�Y��К�������K��ƌ��e�X�����<�T',/�z�\g�?l�w3����=Q�ӳ�����g�uA��<����-r���V���kgQ=K������&�#�y�1�p�}M��=B�N&_�>���Y|}�[��k�7S�y�g�%P�!Ӆo'�i�Hk��k=^����EIک�E0Y�&��k��V:]z��&y/`{p��<8�ǻ�I�u�w�"��Y~�Q{V��ï��8��Kq�.�U�
����ƹ��ގ/<��S�����FI6�\U��/�M���
���i�%+Y]ٹΦ��O�>�G@�1��e��g"�j�*�wv����=������WXJ�ec��'N���">�Y��ڢf^T�.�!�
�:ji<�P��p\6{7���� �/ۯ2p9V,�ˬFGC���r鳒���ϡ<���:d>'��
��](z�^�����ͱ�vّp�vN����dH�)�O~ξ��G���i�l��{+=��E-�wi�32�]]!�V�
�Ǥ��u��_q��܄�_�^�/»��8�h�n��!W�!��華����_���ȬՍ�9�>�˚D>�{|�<�[~�������K�+
�a�L$�CO�iڑ}�U�����X]�-]���V������z�=��8�����B%�n�VD�j�\�ԍ������wS�����<��{������¹�}��mC������	��}10�K ֤*�[��_^eJ��'�w�0���n�oV<�ft�t�|�CJ��';;y⾑1����J����gv�������F4j2Ҩrju��3L��s|�>bY�fV�c�}�9#'������6�o��[ku�������:ɣi�Zɿ�ǳ.Ca���:�\�b�tS����M
:n����P�ts�;P�Opqe;����uΑ�B�?7|����5h|)����qљE�>�Hegi�P�ݢ�i�@��`f�Or��¯������IjX�ػs�D4��Z�Ҹ�������U}UG�Mw��������U�6�S��6���_d�pv�=�zN̈t�5e��vfv��)}�k^�û7 �yW��.�P�Gya���C7j��w4�;u�/��ut��=���f!<9�����P��n������5Ѫ���Oq�v��9nB�u^&��*���b���~���[��ῳ��un4$�\Cg�\�ǻ���!��ˇ{ qgx�ܭ���t�U\�~4!&�91wBD�B<���%�0>�g �5Z[%�St	�/is{/��dVM��Ye����e�����L�
��Y:�e�:����r��fQ\�5[��FQ��=���Q&�>�X:SKکo Me_:�`r��,W���d�ȭt��4<i{�e7o!��5�&��+J��\D6)-{�M�x�4��w��|��;�չ��x̙�叜Bp�{�0�m\=��_X�f�\�eBs�H�h6�lU_oU!���N�����u7���}����>OW�˖ ��s(@1ɯoq�i��,�j�}��]GW��m�kNo���9_�r��\�W��������9J�M!K��o���taIe��\��S�5��kZ3ǻ�؉�n���vZ{:�y�e=d��|����}����.��(e��PA���׉l�gw�����G�΃�����9�E���[��K���F�=���^o�rG�n�˫Gŋto�۝�ry	,���`��/i�*i��}�x.�ܼ:�~+>��ɱ��/j��n�9К�TBi$���5�Q�L��Q�;�5S�M!���k;�282�0Wk��5r���׏��m.���w�vċ�C&��c��\��'�S���g��hxrV�Z������h4�{1Z�@{��bmv*Jډ;>�����]��JW��f�F]����I���ͤ/�W-�]��'UCQ`)�NX_�X�<��͡j�g�f��L��n����V�"�|�xV��l�qxM�~*��x������i���{�|����.=��3^������B�v��iU��/Wxϯ'Oz�u�v���Q9q�{G�f���*�
�i]��F'���r�l�̣�ǥ;oio��{T�;���.HQ�-�n�F+���jRP�v�3�������x
�λ�~ؗ���=���:}�ׅ�N��C5�e��Aӻ=����QR�)�xR��*9�z����lNn�Ş�]-֝�r�u��:`=����IK�i�܋q��	ݐD�2�Y�J<�_5���k�$��Z���3sSg�-�+5,�W5.��C(	�`W���u˫�W�:'��W��~B���6����e�!m�Q�:��pa���c��r�m��S�%3�<Yi�v��Ssn�2f�a�2I5��^��LX�:2��c#�%o�FJ��t�>�f$��6,��&��of�ܳ�c)j7,���(�ޑV�AuK�`���������7�uk<�U5@��W�Ù_E�R��kI9� �l����u�͍�2�֔�H`�2vú�f�JĤ���q"�����B�u��I�2�����S�^�����}�a�xU�(I�2n��u�Oon�@�V$Y����Q��<�:F�"�j`'�lzC� �z���$*�v��K[��j���vL(wH���*���y�h�tW-�ѥ��5�&�2�7o>*�:s抽:$��v���(\=g�̭ ��ى��F�Љ�ˡr�S!%s���S���^�`�=v.�"�ڴ,_|��gUL˂���Q*��`��V�$�e7Z�fL���]I�#�����/���U%�:�S�C\v4����R܄�����'�E%j�p� �y��%t�oI��]5�c�J�+Ս��M�ymH$3.L��Θ�f��cwC�ҫ�*V����ݙ��G4��QQ�De�s������:���ú��L��B;2�qX��+eoO��;��p���,&�(Uѻ�]ܱ}�ө�d3 ��̺�ie1�0�Ð��[6�����ƻ;�s̕��ůx�2�vw6�+�X�hu}�SŻ���2��]��v⚭i<�&��W�W���d�t�L5ͫ�XcV�-깫��B9#��q�eH���uW���9��VҖޛ���4���R���m��Y��˭S�N��W}���1����4���l��7��%,�v�p����9����
G2�ݠ�O�vL���*����Sl��8�v���TDᴲ�	�U��r�9�ce&���>V��6MݴxK}:R�+����]֔;�ؖȈ=��Ĩ�at��b\o�I����[�iA����N�$���ƥN�e�_S��qj��Rjjʶ��X�k�)\I꼂��1�7�CR�]�ؽ���	.���R�D�.�ŝ�(=���z�qf��RY��}is�+h��O�5�>uy-�]l+$k��v��0��Vx�H�}؇v
����vq�|�X�|v��Y��^;�#z)t���*�N��Q��*�|�e���j=#��Ӻދu3�;*�u,Oo�λn[�7|b��0�Z��,.f��ש�!��S��Gk�Mi��k�Z8#�v�N��ζzJ�_��?��?߬�F2Z2cڹ�(�#"H$��]�Λs�`�"fB�%�ۓDl��e�4!k��@Ȋ�2dI&M�Ka�8�)�,ؚ������1���b�D��b"�4D.���)D2���Ɉ26"� � #�:������C2�1��d�c&$�HHa`h�I��2����DL��%wr҉΀��1��f�F�,�0R20RK�`Ɍ3$aDK3%,�(e*� j+-b����;�gYǻ���8��
u��Xw�2F-�۵*�\�Q�U���l����7�f9Ò�0�[T��߾�����o�_�SN��6������t���ӳb��j����P傫T9u\E�[,�tM*|�<�5�W�� �;_V��pܶw��C@ޘ�[ꨳ$m|���ua`=z�&��{y�e��҂C|ج�z`��*�r�����z}�3�M`�":tq'�1��V+;5��!�WË�=MW5���rυ���j]�d3^�7���F\*�����0)�^x�3��Y1"_���:G@@��X:dS=/��0V
�-�T8�^�N�C����o`�t�r��*�Gi�H�/�`���C�_��_���܇�"����)�6d�.�xE6�_Ω�
d�P�~T2H#^�V��3�#,6�n�����z�xɪ?S��a�|�,��Z_�)B�R����?!`R�ԩ��J��\-om{^O8`��[�.J�v��X{S�$���,q?X	:�"t�r�e�K��B6+;�WJ�G	�VI��U�2�=�EF'�c�6����<�Rs�0��[�C�v��Wq�q{ə�}������eA���I�3��!ꬠ�0g4�ه
��1).\��Z������n�xu�v+zt��e�	ږL@�V��u��Wl��j�N�\jq�vr� LZo5����ٕ��19sF��r;7EM����O�������G���JL����6�ի,�>�棔4��]���OR�}k�{��ȷ���J�|k�2�3�o���q�Qxl�k�j?������uw��������������ޝu����Bz/p��0m�j�±_ڢC���������g���	��q���w;�d�:�v��^�x���`�.^���ï��8�8��EW+�x:q;5g۹i��K�̶��+�ɲ!�m�qQ铳��ܷ�/�j��l�׷M`��HW�CtN� �����^EI���x��������?a�#qlu�:������^��3�kހC�x�(E=y�������{4T��֝<
�Ǥ������_q��;pw!��_���,u{,>�K�mU���
��KlU2h�L���h�$hM}�[Ӭ�^���x�\����H����	dSXSV�'�$����͌���U^g��|uѷ,S��^�{v�j2f����v��G��c�p�B%���-�M�R6��J�C<x�{׬ת�����/����So6馤X�뗱(ɋ9�1�w7X�|�剫;�G"̼]t�*�9��R�V��q+��6際D��̧/Kd��/�L�~X�^3*B�����;��:.�a���LYR嵓렪L�B��GY3�	9�?�����ܝ�n���.���sn*t��=�P�u��w`Ma�_W� �K�֤2bB�C�+n��q�L�k����V=3��aΙ�uĆCJ�u�9�g`�.A������ϻ�',rw��z��˂t�
nݬ�]�}&}±�Q�L9:ۭ�,�B]i��u맶�G6�]*�K�(�V���/+®�5���VO��mTH���M�9�sمG/sӬ�8+p����$�U��mh������Ω_d�G`}�k�S��2��=�ܻ�8��}��5�vn,���,�K��P�}������
CyJ{7'��s����R٫�q��a�yq�bt��{_����q(o�(����5֔�*X�0�fE��IF������m�[ VyT1
��T�u�A�[��w��^]��$��ؽW�e�»+�{�P�Gh�����(��Io��U�����Wq3�®<?wvˣ<�\W�^)��߆.�_f�Bn�F��'��K,�+j中5^�Օ\��.J�T��s��/���B6�n�G2�.�Ct��$S���Me�z�ٽ�Tyl]v=�;�Y��[�Yx��#�9cB�s*Hf�}�v���f� �*�5Ï
�LI�5#�K�H&u�͈�|���5῜��9��.�\� 8�-�[�5L�3�9�K���M����W꯾���L(���uY��v�b�ؕ5h�pv4���=�	����-齺�>�z��6e�ZM)�����g̋�ψM?�R+mT$#��M�ţ�"/�Y{r�LU���^����s�ټ:�� b��`��ܾ�d3MrI�	ϊm"G�jxP!-"��ٽ�'v7ז��h�(�Ɔl�v�:V+v�<9H�?	��m�=��l<��Hg�*>���xR�?2ǧ<���3�������K>��y���1<]�W�fp�
Y8�Z@E��%iY�ڍv�j�w���"�s��|���a@�1Z_坽$�F�s�F͈,�wO�O"a3�����w�bO~���=�gn��<S���+E�|���p��b��d(���;~7R�#"~C[��V���ceɽ'd��v���n���;�����e�O�^����C��CG�Ta�o=�Q�"~�5ddֽO����x��q2�r�ih�^?X�ˢ��I�!��A<gL�/��&^fH�c$��ҶU�ڇ�ϫ�PI+�j{I\.�4�-,��Ytc���9�	rDI�VK��6�auN��`^���<C�n�w`�
P��` ��T���1C�Y�j�N*G}��J:���3��(��g���{9e���}��W�7�h�o8}�&$2	u�>�f֜�o������[u�P.�ʘ{#B�Ǒi[����lԜ�r�s.+}$��c4��C�}��h�t�T��4��֯0y������k�L�5�/�Y}=������*":��4螄~6;������P�`�J�.H�qOs��T|���!{g���C�5���$R����4�a/���lJk���ĸ�a��u�y)v�<�̕n���t˸�8*_�vlC>��}�7���*�C�]W�!T���L�0ߗ�����7rw�������P�;��?�g��U�yU�@�������;s���}gC��^x��U�`�g�Mݐ�軳O�����Fn};>�X]ib�jS�~>���d�ޖ���I{���"��O��<��Q�|�wo�^���_!��a*h^�o}�W7�^�xi;�$�U�J_C�����Kíx\邒�����p��/������c��l�|�����V�(�a��Z4*K���jr�K���M�(���c���p4�z��R�Ι���������cRug&�D>�Fe/k.���o��KĻ���}�բ��R�����G� ՜�l�
���1�݈g�p���oi��wr�/{��!h����uԃo]"WF��$A�4&w�q�c��������������}:_���X���꼕X��{ΎO�ߊ�#��_s�H�1)�:��2w*8��!:�bŽVj�e��)���9j�>�G�*ï�c�:O�+�������5�U3���%����K�׵ϛ�{7�Q�����w�W����&�XDPj%�j�*�j7��zhӬ^��m	1���zާ��lb~�=�j���<�W���sB�F�_u������8fѥ��iN�����,7��1���uN�v�ۨ�x�z��I���Kp2�s��=nm��T����6=��+��j���t������3����B]�qӮ��|����.�͍o�;x�]�}im�Z\K��T��_�wv�Tlwşu^MsK����Z�>���ߔ�����-��/ӀǲN�Q���pJj���n���+��K}�+��s�f��j�=�}rU۽{N�U��s�5ٞ�w��V�&���R�#�k��y�T�N���G�	H}��U�|9���������$���΢`ӝdJ7�I�&	�YH�����ˏ���q5�ф�x}�MS�;Y����j���l��Y�Xw��9g���E�wf���!�\��Z���3Sx�G���+��m:S��ou)Ώ�>�>��OJ~)�>�>��?���鵏��Wv�c�F��܏��5_�]��-����q�X��~���'Ly˥'S�6��{'n���S=�M{��*�I�N/o�曓A��?��S����˰�蛼T���/.�`���g	���7��wީ,ٔ�l��4�}窳W��ȹm���&6Ө_�]��P�J�;Şo0[c�Y�D)ߒP���bF�B�̝Y�e�~��7�u�͇#�kl:L=���!�ݢ���ו)�8�������
�3��V	���֭��MF4q-s���q��>
�T*�ɽ�e@�b6�U�gA���M�]��9��/���帄�-v�J���F�>ѽ��z��������'��G�)�ʘn�[g*��yF�M��Ի�?/z�<��u�Z��W��3�=6���<�UUC��b��dܻ��웬�m�WcwdNփ�=0;��X1Y�mi^��ƭ�>1���.������R�:Y��%My���oj��>f/T�w{�v`0S���ʮc*�5������q��
Q6�TZpUǋ\˂c����f���m��������|���d��t�����z��W����v�H7�A��2���$��f���9I��_��o޶�xϛ֯�u�����E}�h���.��y�O����{Ի���+��l�L~�&���P�����%��>���5U|'yu�/ֺ�ڗ:qC[\*�ű�7��Ec�)��uOQ�^�г�j���yح��Ӯf}U����r\��nU��N�'w5ӵ��Oq;	�P y��N�X.�+�c7P�ҽ��0L���F�>yx�<���m��P�`o�����YPf��0zN���<d��%����U��w�t�G�3X���I`َ�τ"��bݣ�w��z�����j�Un{���o�Ӱ[ݰ��y<�O��[2�5�c0i�?\���6�˚;_w�Q�)4�;��޻�8���^y�:����rh��Z�x���W�pP�;i������n<�"�q(����h�ۭEԂ�}�1G Q]�4ִH���2:+���,Y����+��ֆ�/H���9��Z��3��zEe�a>TRt�sO�ҀT��a}��x0��]�T�]�������W=�]Dzͪ����E��_Dc
O[�;�7'F���$rY{�yu�Rw��/	�Կ<A�~a¨�&5������U���iJ���k^+��o�Գ|�sN�s����W��{�(oZ4��'c��š��-�q<�(��fq�׋��|������N�s�%\�o؍���i�r����N��G�����U3ެ�'��s�Z��=���^��!�yk�+��ʌ��C
oOj[�_SY�;��e�6��>�Y��ҝ��x���iw-d���=e�(ݚq���,ףx{�Վ��D��
3��N* �����%�ا�:�\�߻�'�C�1��ް��uz��3
;��٦�)�|�֔���G�TCi�q-����˄�_��ؾ-�S+�`c����^u]�/#Gթ��<.���*�5�m���z�<���u�ґ�k(\����٭A[V���C��ޜ2+��m�wqV�2���)���(6c�.��ކ�j�h4N�����!�׸V����Q ��.�ʈ�1��R��f���i�Q��-݆���
wZ�9��O%��P"�mV��[B<Cv�z�?�  �j9��`n��_@/�}��4���"߼����t�5�Ɖ�T�O���됫';x�AhE�t�x�=`T����:��:���-��M�t{W��ru4/j�:�|���}'d������0������c>��^�(��2��q���9F~����n��
M6vt����з.�.����z��環nj����p�L�c/��De:�Δ�:�X3�h��8���5������K�5���� ���>AX~�R��G k�{�F� ,:sb[V5}sn�I����n�-���I0�q��/BrD˿,x �e5P�Co�fӑ7"���\��������ز���M/8S_&��iϫזbl���+�AG�`�=_DE���̳�jћY���.���;�)u����z� T���>�����g�}6�.߰�md�m�󯤩~Ȳ��S�l'�f��#���Țܘi����ln_h3e&�Fr�
ݭ�
�ٺ�K=pA��D�	Y#�s�X{cJ�oS�Y�@�|�d=מ�A{/Һo�^���ņ�3�-Q��Z帺�؆l����UI� �L��q�U�}#�훣i��ѵ��Uk8��+��N�o��$�1���;�3h��iE�P�ҩ3 "r�\s�{bsZ�r�Xy�\�"�Ń*:T�d�@�8���P6�U�-�mcJ�CH�C��=*�;�Qtk���p�r�7wYYӪ��Zk��ٙB��{{�i�ż�6���e�S�ZTv{�v\#iE���&��ŘWx���V��^d�*�L�@�=���rhC�jZA�1>wm�k9�-P�]Mo�ى��w.R�f�)FY�:��q��^�}�;J��N���{�!B�яy>���>�Ns�(v�-a�N3�����&�fC�D�_֧\�v��T8պK1���b�m�R����LkC�,�F7�V����|ER�Պ5k�;eZ�>jm�#�qq��u�[]���,�7[uP����}N�N�S�0����u+��8���^����t%�:O���#\L�2�6�Ѽ�1���4kT�t�|�#��
���Iv�ͨ徨��#} h����<�վ	�XY�vt_r���7�2�wfv��ۧOK쥽Zӎ�lT,g��u�悫�Z�K�t�����d1�۽��;l���웸�ź�NF�M�]���&^Ѹjh�q+�İGm1�vxr%g��s����1#.�h��%:f����ŗo���~�C��3�t0��v\�āuy�5m��A3 Π����Y,�O���Ez^��mǓ���n���/�T���-9�(��Xz�ǉ���2вP�kn�3�F��Wjǹ_^��2�K�ߍ
�!��Q�}�>'��XR��cx�}k�+h��e�`�b��]K��Q4*Υ�\��;��8���렇Z����t�<��u��:�Sv��t�����r��s�.Y��rr�Pm�T�7�yr�r�B#ɐ�ݠ�	�E�)���VY�J��s�uq�o=��2�ǯno5'%s���y�:ǀ�T-$~
�AO����	n���Q�!�+�Va�]�#qK���x�(�º���ː=��y(��m���^Q�m�x���A��n,{����A»�TJc�抱��r�20��wY�{6���yp]�2�6 p�u}-����t�k�L3���ҕ��oc#�[���e���ee���up:ZV�؃�`]��s3�-.Z:�ʤ�76Z��;(�b��X�\���z��27d'��b�	�#9���s�i�x�]6��5V͍��^*�>m�u�E��/��wA�ˆ*��x�bB�VM�J�l8�����*]�Gko��E�n�S�����͹OF e�پżY���6��|�K����A�.�Nq�;-����e����w�$͒MI%4a�b(b�36IzpȲ2�)��"�cbDL�L�\���7@�L�f�E%I"`�J$�I���I���
b(B�L�ns"�fD�ȔLA$��` &"b�&&��F6�4�)02�2JfD����a���[�Ң-�(���4@��ed�%IbLDL@��3.�"2DA�%�dRL0F�XÜhd�P��Q1s���PA1H�d0d�QBg7':�l�J2
D�2$B"���I��L�a3D�� �AE�AS]n������(�w9I�I_,���C	o3BZ�d�k#��eb(v�t���.L��-�f.u;��}�����|���>��^��3�����^�&��{]�}im�|.���#N0.箼ޫ�:i� ��~�A_{:v	T���vǟw_� ����aT��'#޺o-�3��ۜ�;:FC��(���=�?g��s�f��o� �$��Y+�LWE���OPG*��������-_�-��M��K׾*�z�՜�ݫY���͖�i>1�9b�;����\�]�χ�t�mِ��/����ӥ�F['��ʹ����.��t�`�)I���%�/f�:[��};��M����\���=�;�n,��6[�����+d�T��X[���i�i_�ﾩ�XS��gM�xy���}�M̧�dw��+��zq�~θuc�x�=�~�{����Y���=�Y������&�3�A�����<8�<�K�m�:L��3�n��y���s�������]�1N�b�i��|kih鱀�K��*���Oz� ov�vշ8�qV���/W�J���h뷺NJ3�Tѵg��*�v̈́��t��i�Ut󷠚���꘱�2��l���c�thh��mv��N@���UW�f��Bm0+&d�>.�[_ �sQ:�/>nu��ؑ�_w3�}o+�zPT�[T�5�=F�-���T���A��/)F��N{��/:���{k�H��Һ�\�j[�Bj>m�8F��ȝCb�z�_N����v�u��.�_�yɆz��8}���w{b�W�yu�8����q�g�%�Ô\,ۋ�ճ集�q�*}{=�������^��{<�.�Or����vhֺ�!�>G�/���8aGO���������Q�i�xϛֵ��1���ܭ�0<��=syz�)��U���5'�aŵT��AX�-s�2�c��>����������	�/�?-���e��Eu;���\'�q(���k^�z�QZ�{�Iz&~�Y~޻yT'��>���_�Y��vڭZJ�zXY�'�?^�W�gws�]9�����p���rC6׽�K��)畴w"���4�|�A�T��E̶vu�ES����O�K޷�lK�auϑتowGv���{�u<4][X>iTI��n�6:<2%{�%�ޙ'J-�t�����+�n�#T1N�6�f����1�p=�6s75�/K�Уv�367?G�aVic�5^��DR��:��oێ��+���Md
?kf�k��#l����圹������T}-�;Ƽ��{jޏR��4orR{��x8S�w���w��>�>���M�u����v=9����s�Nzo���p\�ڽ���P)Ŭ�U�^U�E��J,�Xů�G�^Zr�4�����SW~�.QX�gr��������Dc��IgJ�3k'F��w���F�{�҉/l�����]�sҺw3�{�	cҡ��-�S�������tz��ɧ�zz�KJ�i���-��ē�q�¸�tDƠ��<MyK^�������U�"���m����ub{���-�ﷱ���B=]�J�r�����(D���w��Kry�/���kO��zޯ|�z�9�yK��网�ÙuU��w�fIY��)����vmNJ���F�1�gKYh}���sɧ�v��f��½���gy�`��	�����tknc��'��i]'d�1nz��"~�+d1=�&�#٥��*��	�A*�V�q��+n�N��%-�1�W1��.�:rfM�.�r�+2)�;�&���ްg;�5ju�q�foo����������>����������}J��~��<S�i�Lja�뭶�RCα�m����S�JrÃ�V-EI�����i^��TW�'\3��űQ�6.[yr��'���[\[Ц3d�g���޾s���+�Ek�����]+�Ÿj����y�o22"=�Gp�g�x./>�X5]�Pݘ"�r�W
�,���~�xTBk�]���^��q�=:�گo;\��P y��yn�X�5XRw����D}fz΍���8e�+���ʒ͗A�ξP d��zV5;Q�Y��얳]z�q[�ФM�b���q�ǩ�P�����aI��;:{,WV�Nw�՝j�ָ�vk7ی����^��xWɱ��DeFKH�j�qj.������N�3�n���F�j�z�>A\���_k���{V&��2Ȓw9!6��"�q�Y�s"䐘����3��.��7.��y���j�� qZ�u�)ԣ�mb˻���$�7�5.̔`S��R��jga�;��;m?)/!�u{e)�[�	AnӞ��N��]W�;�r�����<A9���/���٩��W��F4]7�4�a�.1�î����)a�/[��^ ���cʬy�ß4�)�����/��s����x�ɜ0P^yx���/i�c^��!UwJ<գ7<�\�����f��x������9��>������=����̫>�V�n!9���m@��`-BϪ$����:W%v�gm������s�:�֕���7����Ս�k�;{Փ4�I�^c����:�_KŶ�{.1��z���y0/��xvf��8�w,cډ���J�p�''-��������ӵԜ�������������m1��P9��jqBWe��lW�i��6�ǬY���V�z9~��VZ�����B�vО��)k�gP�ܹ��]�«UfÛr�WTw���%��w�$y�t�5�/��|���2s������3��~�Ҧ�'zt�]�b���d �A����ݧ��#Hb9��V	�AX��b�I��4����S�W��[a�67�e{F����h���1I>�`��G���Vp�hN�������a�����S�[��+ݓ�����g諭q"���,�bE��?W��;��)̃���������u{��m�Z%g=y׃���;T5Yރ~�F����)�޵�&�l���i��L~��W8�
�{<(c��@^��{����Y����Y����+�`ϝZ�5"�$]	�;�o���2mel}�z_�[nt�s.ٴ	�zj�U*5���$��M����O�~����b�{x��z-�RZ�x��^��}��Z�+l��o`=�_J�S�h���yJo�c�^��ٶI�����){q�*���Tj���M�8F��"�\������D��[<at�lRf��"���]���/$�Z��9_���;�ob�x�#ǚ"��1g\z�Kl/I�˕'.�ӯ\f7W��k����=��D�彚7	{B}�{ >�y��bʴ�V��>{���}Qw�ݙ���g����߃�e�+�$�n8G�ϩ^k�������qI�γ!8� �-v�Bi�;�~<��ն�������B8=3U
�	2��m*�	%;�W���k	� ���i�J���C�Rm��Z�2LJ�ݸ���&r��<]43.��}�ά��8k	?�Ꭻ�.�؇��R��#�WՓz�>�c���'ܕ{=L8<�d�8���c��l_�/ +Z����j�6�u�3p�'흀bݹ�E��{�z����ۧ�b��TsGڏ���}������
*�p)�yJ�b��5�m��i�3nC����	Yi���-Wi�
"�A���~�K�r��RZ�6wnoC^�xT6�Y���CY����l���?�{%ګ�s�Џ��>���\��+�Hi�V�c�m}oG��ĳ|���>���}U�}��� �FM7����c�ڻ���Y�SA�i��^*Ư{yoF�֞��ur��FPI@�2id�M�t�lc��<��aS��^,�K^�sN��ʢ1٩,�Js���@?���j^f9�N<j��zr��sO������f
�T4�-��|���D��e��d����O��}��\�n����ܜ�HUu1S/�V���=x����aT�1�2�SK��6m��O�![�Z[m�y�-���VtkWS��8\�{z�9�S|�x�6���)�Q���ڌ]o,���r����������~���]-ec�=�>ݜ���u$�w�3�"����p�A1��w�K:v�r����zj�篪��N��y����O��e��*���nt��Vb�dBv1w�u���f���֟O3ޮ�����u��ɽɔ[/����w�Л΅�:S�GX�w����݃*�:[@��/d��y��&n��ĵ&���������x{�]���++ȿŻb���t�c������\���wg[|�[[�{w�]�kaV@
�Fͥ�+!�����_OVM��q�☨֛����o���_{|r�����n)շD�6�Wj+j�����å��طz�m����l�PwLљ�~�{}����%�|ORn�O�o¶�L�d������;����*�}�׃R�̹tr;5���P��]|�@���ݞ�Rj����P��;�DS~����[��)&�;�GdE�7���qY����ez�+� �1#ߠ��^\7�<2i����ǐEB����P�J���V2Ը�ub�[��c��q�����5��(Ƿv�^���N�ّ�NҦ��ЌT��+�nt}���;H_�W����m
r*D��&7*-��)d
?o�d�@����=+���ق�G_*���w����p_��m�y8���>�(�"����&�	���/���sS�R������b���ক�x�c>M�e�B&Ptd��>��=�IŇ���!~��7�S�Vy���ӕ�Z�����>AX~�R���n�z�!R�3�m�6$��_���S_M�ʿ�S�h�oji$øe�y�UÙ-�y�R��w��s��"�΋��o,G�|r�4�)禓篼�}��s!�p\�0�?U{)PM��q�#��w_����=�ћ�Kqs�Ns�Wk]ي�)��ym"j�͵[��������x���r���K��iM�� RU�Nߞo�c��p�3js�]��������}�4�>������_a������b۩|:v)s>��gN�oC»c��~��6=x��}�;mn\���T��Em ����<=�Z2��͠����6���>�k�sw�2�Ɠ ��S/�f��w��9��Tn��Pv��h#�4z�Tb�G����H����9û����P��W'�s�l�se�J�ʓqۛ�9��/�QY�r��`�O�r�?mUez�(9�>���� ���WwnT~۰��^.�I�Ǜ%�����]b�l���"\�Dℰ�6y��ލ̃���0���9��k����k6��ǋ6�qz���N#�հ~������S�H>�N|��	3�'z�7��������v�P y����w�}U�ehu��3�%������e�)�V
K��f4��E n�8�����\G��^wޚ-�c�m[c��PO|��^�z�ĳ�۵ޫ'�B����=j���y=˂�P��������u�aY������y�7�Iph��}('6��އ�ѭ�:L����X-�_f�0K6�OG�:�����p)�W�8����^�Z�ݎdqE��/��^���<A�̸�p�T�gP�:��0V,yo��*�E/g��W
���$XD���9�Ivc7�9����/D�<��<U�HЍd����U_b�]��w1�v���`we(�_�g�����ӕc�����uP���;��܉��v�]�t���	�4#�C�]�6��dE;�VJDw,��5 յ������.����Q�`W���ӱ�N�]���c+��od�"_`6^�鹪P�lX�Lȕ�H]I}��jj
�dX�r��{��G-gӕ��1�i�]�a�s�[���t͠�����麬���ufI+�L�3��zGW0r�t�7��P�Aƹ�H�Tv�Ka';��VS�\�5Z�2�αp����.LRӔ�]���P��/7�ֽ��FçP�pУ{��J�����7�x����o��+���"��_>�B�v%�G��.sө��4�1�&����Ӯoe��w�6n�_C��C��l߅Z�_[�J��X;�;7/�p�FE�V 34G�?\�-F��[ʨ�������#,��>'�k�m*�wu8���%v�aǼ���2�<�\)�f��Xy�'-�5+��Uo��р4��۽��f��^��0��}k��}c������;{�\c�&��k�Z]�����b�᡽u��S		������'u8 y����=����轟!ְ�ͤs�b��y� V(�5�gUɘ��
ރ�9s���]k9*k�S���{��2�o7BVm���m`���W �:1�ŧw��0\��;� �R;s�Դ�cGS�+�;�Տt|���m-a�L�&�{Lb)�ٴ���q��l�K�$nP{�ivv��ݮ�L�m�.U�s�*=����su<<]�]!`E�B�wz����o	�'h�;Lhj���E�^��z���t�Vi�R�H�1�;�n�����;�V:ĂcNڮ哸��Ȯ
ڲ���Jy�&]J��K�m|9�r\P������)ѕ����3W��+�=�v�wB�l�A��7���9��\YO��f�hf吺����ژ
H�#������h�R��Z�`�uI�>�ҫjw����4|��۲oe-:"i�V���q	�����J%�A�����b:�[�Wos���z(��%wa����������� 88rC;�uv��	1��cs�h,!Y�V�lov�ZI%l
�j�8	�`V�֞���)�c�
�ڵX�;���5G��k��k8����)�K��h�M|M�6��"T���v��u�+KW� [j����sAR�ςS2^�)�g!a3=�/�d�L�(Y$:'�{9kW_p�z�Ю����F�^f�p9NҮ�:���0�8-�v������f�a����F� ������f�{#��s^ŵ2�A۹1ا��wyu���R�\��r�(oIu��ܘ��a��O\E���W�.�D����=OgtTyV����DM��.+�m��J�!t-���i�+�P#+�_%��/��%���y}ʁ�P$�	(�r��h� d��@�!�d,�L�Bۻ�)�A(HĂfIDL2wp�s��bLDL��4��A&�%�.\I�00�� ���*f4�$�w@�1$� ��0�@�&�h�`��I��E.k� ��"H�f��cb�%!H�����i�2'u�1)��J&"�3@�5�0d�)��D�A�]�4DH$���b$Lr�ġJ���!�$cnt�1�$�bIwu�I*"LD�	���T!@2�#(Ќ ̌SA��9$�%$�BD3J%f� �H �QI}��mڸo��SS�7<w�C�P���"��k��1�v�>5J�b�n�J��eą�$5�#D�71P��|o���!f�Srk�������C{��^�%7p�(�vDơ�𹣯�5T��o��y�'Qw����]�g��ɒu�����;bw���Ŗ�p�w��ZN�18���~���N©����md�l�}�kW��z]���o��J �aa��3ؽ��S;�:+'�$�K��;l
S���gNr�����};���쨱c/d�e��Ͼ��V�g��T8��.��t��AC�owmQy����EVm�>Y,׭�=/[ϧF�y�<�����@��ح���棵�w�����]�3����}}��W?nw��^�����]Y<v����l��]������t�0�-�W�������7��3����#Fe�����;���'�(,�J�bo/5뇁e6�\i��^���Q�}�㯙TM��	t��̓�$���[�E��k�o�1ǵ7�/\��c� l��3E����NwA�NWEsIw�M�δSt�E���,��|���k%z��M�R����7ۯ;��I���6ΐ�xfM�ۺƦ-p;.1+9G�7lC �Yub�.��U�]M�r*�5ͤ�޷$Yz
W����Mi�~�x�F�V3Mw����fPGJ�l��� g��4�sc�����*�^b�\�X���ϫ�(�#�F��6>��^u>�p�z�������ӈO���3�
M�TC�fF;5%�+�9�h�VV��֝W���1Ed�����}�5띆އa��q?)Bb6��]�;�q��5��M��A�\������f���˨ojjL��c��&1��6�x����+)r-���(-�ϧ��\{Wت����^p�5A"3ڟ���p��Z��P���3�"/=�g�%y!9��s�i�>3��߁	��#���6Mi{�ߪ��n�C˭Q�Uip>��+F��a����oy�Z�ٻ��Dz�����\&��5Gk��x�όu���>�~�t��k�~[Pa%��{2�)������J�N�L�cγ�t�c��ً�z����\�+ ���
��K&���d���n��=���BivS1v 4��0���U�f6�sq:��s-���XRi�l�h����6�����ZUl�]�t퍗~)qU��n��m���Tͼ�@2�U�R��k�S��܅͎�S5���飣��@��q�Ӹ��ܬ����B�u3L�l<��.>���V��#����>��Ƿ����yz�m����k��"_�����*2M⣝�N��J)���[|�}2\�]��=ûڇ�s��L�`�h`4����Y;Ou���l�ĳ�y����=b���eE�5^X����[�ɟMcl5��-����ʒ͗O�t�N8�	\5^�?O����MP5�+�YOv�{��}�Y�QP����q�Z������ӓ��oދ��y�&ٲ{�^��ʇ,�!SY�'}X���~kޙ������٩ǯ<�~z}���z��3>=ᾓ#2�d������Rfʁ��rV9��mnV�~zSojjL0�;B��=:����Y�x]1o��P�h�����c��~89�~�<���i���A�k�v�����	�ݥ���2�WJ܉��+"˭WO/7����{���x�;@�HJ�&� j-S�[q��z���]
���Θ����ӻ7l����S��W]-�*�}�Ir��>��k��v8�#{|�i�]Ò=�/�%�<�9��GR�^,���뻇����h�>,d�|}��w�����S�W�Q����3�{�Z�N���	:����5�Oӟk�x�෵=��n��x��|f��:���Sq������כs�Uw�p�ps��w�ļY{-%3B�&���W��O��^�Xqo�>{Ν�U>���;�ۃ{^�X����H�f���0}��8Ԝ��ڬ^��Q���bH��ˉ7} ���P�_fy��.�o�O�*�G���P�ᖯ�ǀ6�P�8LݬnUI9���H�>�~a�/X�N���N].w[����>�<+n��Ӵ׫-���`���;{�WNy��vl��<���ݙ���~��fv�[�����|ˮ��O��Mχi��$���_?��z��t��7m%�S��1�׏�;�����[�q���)"�1���"�������ΥI��Pݠ�:�j�˭c���@%�+�|Ћ�S^��<zY����D��!��2&�r��s��f�e�kɃ�k�z���h�0�pD�;3���;7GG�}�t��d����`l�Q�9��Ãue�`���[p�n^��^'߷��m��H���yߧn\Ҹ�g��C�B��UR�|t��K(�}��r-��i��j�l}�z_�[aΑ�m��;�=���l��o��X��Qr`��)�W�8��όƼ�VE��T��9x�6���-<sI���� �
� �����w()��fLyh��sۗ��4��^��;����'KSύ9�7�W�h��c&�����t�)�nNU��+�9�imV&�MR|�����������c�S��ά�v�C���s�z��5�=V�܉nNv���������z��zh�n���-��=��J��3��A�����ʴ�p���9Z5Μ��]�D��{�	WW�A���v�j��դ���qʿN%X;�0�Z���>�"ө[o.F�p����:�<���~x�E�~��W�k\��T=��.#�O*��5�xJ{,㪸v��{[��֩6V��KrqC�6�G�����s��ٹ��W�!��B= 6��T�Lcjs1l�FX��w4���Y�F��R9ݏ��An���,�z��u��5
ʌV7(U��Γ��3��E�#���}\n��u��B�ƴߥ��"^�-�f�ϥ]�'�)0ġN�f��r���'���u��_х�Qn�������7��e��G�ޱI��ɒ�Q�=����O�q�������;�Zo��8k�ʆ��>��o�����r���8o��Ewi=JvO�KԨ:����i�ᦱi��(g���y0�8,J�ޟ_T���v�Ʉd�Ӟ�M�w�^����/���iM߶���{����\ UpS����W�Z}��T8��GOq�>>�-�4�q/wt�f��^�'v�r�AԃM3��B�5����	Ժ�zY0z�ڨ;�����>��xv2ıң��ׯk�����s�/\8$��ak5��O�=����$���c�Q�+�����i�y����G�Ǘ�;֪���R��9�媯>ɒuՉ����m���_�gE'mj�՟6���e�T�{wv��A����]�M�J��Ԙ#s���9���*Q_|�?q�o��]tX���=���W˰0�W1�I>A�aC+sU�V)Jg�������lP�wb�f9��Ĉ�Gu%<��{s8Xޭ�_t;��"���(����c��s�Yb�0�	���0��YW�l5ýkϲ�ٺ����d�Π���m��9Ӝ�٪�%�vm�we�'�S�;_w{*#u�l]��;��o�m\�f�K)*n'&�uğ`���M���z߽��٨���ZLo�;W_x@�^1{�xx�%������[~.&�1Z�b巗J�e�	ᩓ�:n�s>�9oBvR@����Xlm_��o}8�+�;VR���6���ѻ|E���4M�|]���b��K@�G|��sH���<9��Ϧzڈ���6���gs=�KL�#���½b��	U}��5�O�m�z�_{Ԇ#�/39XYtxl�{ �zn�f�<�.K6]�:�w��*�\���[{�p�˚JNa~��j�]ϥ����{�oT�,��y��%���-Y:�،n�{z��/�����uϨ;,x�ڵx1B�s��E
�-,���j���v�ӛ�\!��V���Y��a<�^g��$�/�@]v�a|{��ʈP˥�XG�VG�/	�R�u�0_��x�,���'XBVʟ-�O�ɧ��o6�j�Z���o���S�#��j�_�����?g�[�y��9lJ���]ٞ�Wo�����_N-y�T���M���A�xV���_����m��D��j��-�����b�{y�s�z*�Mꝃ��d�{3"����[�r����F��%sE�|���;,=�y}u�RK�v�ެ�-͋TU��������M�;��c!}�f��Mt�v�^�o��B�UU.hc2r�w�ίo�N���3m'r�ټcp^� Nt{$�˕.w�:�{>�n�)�k��cגqǟ�M�Q�{l=�ں5�lY^�9�ZXi����]=n�b�ŷײ��*i�h��|��՚~�
��	؇�]ez�w<�W��-l�Ƅ��i��[�^��c�����A���_nXSk=�9]<y������n��{���U&��q�>= ���3.�g���.��<C�E������e]G$ƀ��@k5ǵ��G:�[�+�|�2S�ǟ�{�_��cӹ�����d]ɮ%�e+ѣ�+Z�6��yZ��ś]G��NS)���=�J�ǫ��g��ޗ��y;�}_R$�O�K�x���Y^c=���6Ͻ�yJ�un��킺sśN˯�'h(�w��]f�F1�����[�#v�1���e��� �/�{�;��$�e���'����ؼ�o)D�v�͢}AЫ^����=����Ӽ��5��q����$��kڤcz�L�'Yk�]�¯��չ�J�;���7����!,�U�<����Q�ٯo���E4]o�х'�-�����@ߍ��n;�ث3;�����l�wܲ��,u�":x��>�q��9�(�1��{��ʐy_�;������ws=��og�xE8v�]@Yr\��#a<�5��E�W7��^e_е�bn��jÏ�_Ӹo`37��[�}`b-=oA���FS;wQ6���b��V�N��d��@v���;�G_�(_[�BB�|�����6:u��v����I(q�5�0ru���Q����0��Xt|C�z���O���k3�ۅ^1�J��z�[�˶��9<�g�)��I��H�[˭�{�wKk/7/m��SD��gL�3�k�!嘆ǽ�wJ�o/��Ƚiv�%�����Mj��B�����E9�N<=[�	��ݩ��KU8�d����Z?G����{aI{��S?[�o��+�Q�=Yٻ*���׏\X���S(��u�)>;,��o�~����z�M�B���X�����t/8�w�L����-5�:�l��<�(˝qQ^C�5��w�=܄E{�/B[^tZ����܂[ni�=���
z��lG��~-��pכo^pk�k�~�t��ղB��{��=KQo�Rmm��=��4�^�~�}y��&�@��-By��eˬOo�Πh�d�&ǝ ��OR��%�5��a:e?SZ)ȹ�����g�%H(���A?��}0zy߻d}��qO5�77������}�������*#(?���A7�>��_�;�p��<��_������F�DI^�E��54D��B��8|��l�#YZp�]]�"F������9T,Jʷ��tdDz���6�w[�u'Ѿ\�˩g
T4�ļ��o:d!�H�B�hEd-����
gR:n���љ�8OLe�o	�Q����Wm+m�[Ξ�T�$��e�=��\���X�:�y�X'6�>�*��fJ\��{C�B�M�]ۯmb�[*��B��3Y�z�z[M�wl�����A9��� ݫ�h]Mc����)>�W�2u�3*��8;἟|mu&��R��T��t�fK.u��E���q��z҇�w���Y���/7��V�U���Y� ]�K���)F��u@8+��+�S��`�`ùwn���jcqd��#�Ug]��z�&&��Պ^g�OY��KR��I���σ+T�/��"���{t�[)�:��Z�9u���1�&�\��!��/d�9t��](ns�	Fj	#'oN3�.��j2�����̊� ��E/۱u� &r�e�;u��F$�r�rquлA��靃�ް�.�1�zm�g`ǐ��۬��J�Z��ĪM��w�*V��[�&�^bsأ����f�cx�w��d��>=�3��0�Hr�W(g׊��r$��V�q�\el�n�)`�fXv�{����D^e��4��(& |r��}��2PN��|�<c�e�,a睍p8j:���Wf��Ʋn��!��J�v9H:��v͏g.�|�K�V�1"�d�Q����|�U��鸎)Es�R�q���:iO�-MV_T�|9���Hq�ٜ���Z�o����c�G �6ge݂CW�6o��7a��<���C׋ʇݗ�W���M�ړ�������
�z��W)��Wo]hW\n%A��捿/�'�����YEB����.�I\$�%\����B[Y��XF+]91�s�;�e���W��`.Y�(�Ŏ Zp���2h�6�7���*18@k�a	zw5�ӅS��S�%�@�'Dul>�;:��*��ݏ�l����m�Z���2��N� U�B�@�� Nއ�2���n[��@�����09�#����!v	M��2>��VF����}�y]���Q���Ͱx�5�]�@����a	��7��aε0YJ�g[��5�;���2pl�uע*�.;ޠ�����u�Z�����#n�F�J$=HNܣ[@hY{�Uɢ�>���`]0���a�����OZ�e��Iu��f-��QɈs`��o��*�Ys(�.�=�:��&b|'9h��k��w�>R����T�{Q��IK����Cg�6� Wc��h���B�+|ݹ3��`�,��omX)��[p�r�7n�-���o����.Q�64���^{�Ž�ǛqyP�\���Ȳ�e.��s��{ڤ�Ҕj��:Ȓ����	m��:������@'�K"BēH�߽�R3>w
�h	�bIHD�/;���Ț!��J"SL�$�nffd������K��Ap@�	�$��+2)��H�L�;�I��$c!Ewb���QA����i!�b�P���M�cMݮa��))D�A��dɤfě��h������C2d$E2�f���^D^wP��Ҕ�J�JBM%4I��yκ�a��#d0c�WBE%.��l9�7utE��q�t� 	I�v�B�ݺ1�4�H�:�D	��H�)�L.까��02��f
4��C$�Yy�"���=x�k�h���W��{�޷~�fm������e5XT��Oyh2��tC�jF�(�^eodҰ�ewI��8�9�IE�}Yع��ম�w����K��¾M�C�P
�e#1�U0��s�
c�X�O\Y~�22���yz<�m�v�W�J���L�li�AdA~����(��oȏg'Je�U��x�m��BI��y����^2�<^��;��A�t_��W_nP��<����I9���VX�>��dc���i�6ck��7��z�a�trm�|�ve�ټ��`��˘d����v�*.D�c��o��]�=���F*y��jx�*�k�/S52��{۲ȯԓ��N�����ּ������t�����]���e��w�s<���
t�3o�W��;�}��{����z'������X�t�O��<�)�����5��X+�)A���q��6o����a]�zjfHGٍ�Rl̰�_קv�e��s�[�����Cy:+�d���5RL�����X��ʙ���u���W�����tf�e��k�(H�+�dS|�b���b��/�	�]o�P�']��K�뫔eF<�k���z�6����R��%�Wthڤì�'���ڟw#ͪ��;j�;N#3�u���Gz�Q���X�P��}�g�:���?J�-\�.>�EJ�W�8I��bt��ٲ��D����M��Rҹ��S)�$�J���`�M��h5����T*J�6w�z��z׀������^��M�~�tf�v�Jzj{M[�N/5��2��-��G_�f��Ͷ����ެ'�}B�����	����КJ�V߼cֽW�z_��c�gla��{UK�G��1��NmX���"��W؛W�EM��-��۶�Q�PZ�{��*SLž>��oV}N=���׽2VԳ�l�{�~�p�	�Կ���z�+����;=�o�z�mBؠ�y���b�^<��烺]\�J��p��eP޴h1�o}g��b�6%����N����L>��
|���a��|�2��������cb�RŻ��!�p���^5�a�xҵ����{�Rb}����|7��ZZf��ٴw�R�j��C��T���.���jSKy�6g73���=J�;���זt�:�ȳ���v)u��;>rY�Z�f���T�_\��K��&�w&����%/TN�q����\�_�8֜����֮Սʸ'�p�^{}]�gf���v�Ȫ���[�	�G����{��_r��Z��'���ݚ�Jyi׺G��ٯ��G��T/�T��x�iCn�/%���)�~�kk�5�y��D�[�e��WV�լt��My�U�ݛ��ǧ�Wͦ���ۗ�_;ɍ�>�{���*9ٰ�.�����r��|�Z�i8��2���`n�=��m��-=�7�#L�CG�I����īT���'+�~�>G$/N������T����e�gs�y�D`�WQyw�{��]w*Zl��nJ滵X�{�t�p͢�,��z��t���T�8�N��u�7@p�����J�M�ޛW�Hm<�KRN�c�3��<�V�ʇ#@�Ϸa�:އ��}�I�=���E���,KW���3Q8�9ע�M�m��^�Ӥ�skD���|p}�t���R����jj�pع���=	��k�0i��&�Y����1�M��yR4Rƶ�q$�_,0�Էi�4s��ң9���k�u;���(���ã}\��)ߡ�e��}����D�)�IK�=�W{��k��wt��~��5�oC�^;�0�	�Pɀ^�M�?&I=Y;�^NF����><�2=2y��u�9ڷ��p��fP޴v�^�v����������>��1�S��/;��wwS8E����Uf��v�fߣ���1�"=����ZSj��nE�S�5��:��!Zr��o�>K.�@�>�A�}��>��L�W���*s�Oab^�y��N�D@��]'(�Gp�
;�N+�y�4�^�Ojiju��8׺�l8��+���C[��v߫��D�����j��ly�-����~�8��|U� kkO=}�5]oyUh|�W���'��}���LTF���o/蕞�^ټ��RbJ�|O'Ǖ�Jz��aA~��}\��ҩ�[��Cm��׸�q���#p�c�z��9�^�^�4�ޗ	�VM������ģ�����I� �Zy�B�5��CZ&�n�zC׎-lh�p[-Dȭ�ܟm�ʄ'�W��g�=�'X�j�ە�d�7[�MnWV���#Zu�i��O��дZ�b��pu�T�V������:�r��x���-���NX����v)�x9w{=å�=O{cFL����������cWωf��ڒT��Wv���4.I����{J�wY�75���\y��z/�Pl��t8��'�n^]o��6�u8���Ҋ�m_WkV��r�{�8y���|�>D)߷CS��������f|:g&3��~��y�ލ�
t�{6OrJ���{^����PS�~9�����T�0�+6j'^��B-����z�z����ێ��=��Z�}�bH����)���oU�����^�]}���{�Nn��
K{=6ˣ�[���:ѩ�y�X�^��K�S�M'�����)~�q�y�Ґܥ�޸L�U�s�Վ��ۊ�����g�-���[X��{��~xg�72f��G����RXN������ޯ�f��^t1���Rt���o�r��=3ݏW�e���ڣ
7��M�E�R���G�%:��sx6�Dw���{�xP�W�׸=�ܦ.߫	�j�W)�Q�֓բ��+M�jC�U�h��2����k�m�r�R�� -�ض��[m���׳�Kh�ZKP�jc����˳Ҹ�#���l��uL�f{#v�Ԝ����UٞG��T�({Gj;����.�ɞ��B�������uK��d���#�.V�R�߻ҫ��x�{���{�9������m�L����o��0Eim9Urp!*���P��;��K��wv��oݘ�-n�I3����X~[b��j`;2���$cU;;��^G�,]����]I;�^t�����׶���}��,R�b�(d�Ԝ��f�4�����x�잁�/W�z���z�<�^�6]8Nҁrk��W�۽%y�����/wԨeN�Ļ-�k.���ݷ�2�ޕ	|QW!�.����{�\Á�Ơk�qU�rޚ�{歬Q�=��ϩ�^��Rs��7��n��<��ԁ�zi�u���������wI��f����ʽ3NCK
���c��� 9y�P�]|��4�O��V���/�F�Ý!���C��v'k��6�+��C/k�E��>��-����A7>�Rߕ[:��՛I��ŸW_:�5�imcВg��ʊ[��V����S���i�մ��ȒSt�1�-Vr�n�#��r��U���K׸囵�
싸��>p̭�!�0��V�YǷ�e_��u�\�2:��_���nt�P6�W-,͋�j����oCaG��*bT;_:�/()��zI����c���&��>�m��K>Kjk|ؚ�7���g��,M��{��_Oz#o�E[��z�Þ�Ɩ�o��|���5]��Wz������~��f����\�d�K�iqW�O�\�;���n�a�t�i;�i�����������c���*�*�G�?y��L�]O\��,a�h���j�l�q�s,�s��a�W����.���`
�s�u]{�g����t�����4{�ޙ��<�;q����n��WYg��;oixm����w�R�v%ש֞iI5�\GGT���Lyd��ۭлm�S�v���e�ѝ�W�uR/61*l����\fh��E�w�Z=�:���mt�=�}q�W���o��Э7�2I��eb�}ݓ����?E��n{F�L㘖���}V��p7����wOqSΣ�A�i�w�8o~�k�W���"�^�_��+Gz0E��y�w_nD(0�2���l�:��IOޯk?tq��!�	���Q<�{m�1�y^w��
dD�	�J�
Zk�r�����C�s2j' ��=Y��G�6�v��L�+����W.��*iԑ�ڜ�RҫR���ۛ���e ��.*z�E�Qf[��u�����c=�G��w;�ر^l�<�_��Д��L�8�OV��\�k��z�2��"E��������������y\���F�O��躜�����3]	V����C�%�D@�Fa���u���\^C��*�ߺR��x�.�e�?���3{G0�����SGs�գI����F�uS�.}" nG.%��ll�{�ѻ�2����S�]5}g��Q���|z}���NVo���:o��9�Z"Kdi ��:�w�}6}����7�WE*�:5���j6�+�7�t�'��g8��XC�d�E��E�j*.�R��[F}C��^�Q�>�XoR����H�|������4{�@·1q.�8U�W�����FI�g	��za�f=�/���i��c1�XA��t/Ϩ9���;|)��=��������-��A��Y�`�[՘n)K��Up����V<�>��&��=�w���@;s����e{��'M�vU��_�G��}���g2�ϧ�ߢ���*������K����+`il�!=���vn.���z�[T�>}�*e.��F�·<�ⅼ�˽գ2&���>�~�3zU1M�2�	��U����vo�hQ����Cλw5�_M��f���pJ�|��@t�ܱ��Dvq�{�s��vME��$�Y�:�j�x������ ^���b�x�~~jY��,��_�/ƢNUϢf�z�SQ95m#�3�N���Zj�������G\�+�w;��
�Mx��p\.��2�����1��ݛ4��O|&X˩Tp_�.�S�ɞ\aw���ǁ���Jڏb�i��%�����:�x���|Ou��= ��詞F��e��=V�/tu1�����K�'9�{tu�^�ᎇ��f���;Fa�K�����AR�Ѕú�<w4�ܴ+�-��rMC�}Н�����}�Ь\�jd�8yT;�٦�ϭ���ы�%%!u��mA���ė�~<�O9�}�@=7�De��
%yH��I`O���r>��I�E��u�#&��s�N�b>����Ou$Ttϸ�8�Fq��#/���s �P��U�n�YOr��wtie_h�c}<GNm`7e"�g��#q� �/�����l���9���;q�\dM5�����H�Fgc��>t��S��D�榅�'K������r5r�q{E�ϑ)$k�j����I{H�{ػ�ѷW�q&��(f�|9������ީ�<'b��l����vk�n��R�� ��97�U�u��	]�̌�yR�]�.M]m�_t�QU�9�%��md#e�	f˖9�pҺʹPk+R�˘0l�VuLd���O�������R�&�&}��&�fT��c�@�񊈗��o�K[7䩎��r8_r���Xt|̓+*��H��Y;ç@�������K'j����T��3���*�{Қ}5�x���aȚ�v�ή��u ��}|��sC7�RB�%P>M��u՘n��@$؜�5��1&�Ն��C��7�~�^O���c���e�NZ����/�>��GO����(�@Nfǔ���\�+��`˥]���l���n���7�;�8�w�������z�����C�:�Zx�3�'ӝ3�F�>���z���-�^s�p���{�����cvr�ڷ�2`����}�?.�Rz�c�|��O����	���2\��p����!;}|��-�����L��gc�Y�؍�:њ}���ŕ:hq)lA�~4gj��H�V��F��
�]:"�n��)�oSRL����қ������]hpF�F|��#.�t�����tg���s��2�d{6�3���Gv���i��>Α��n;��:�pF�B�D��	;Q,�ȻUQQ@+t�w�N�.Q���]e���ɽx (R��̱���2̓t����"\��
в�iƜ|�G�{xM�-1�1�>��W�YY-���&E�u���&BF�e���1���%��S�9/�3 x1|�"������Z��>n��u�掅*�M�d��eYyDb&�X7S,�%��Խ��cȻ˱Of�2Z�g���D��q�9����\5�8Ayd܊:ڐil٦`���օ��T�v���7�to]E��W�2qy�í�JM�k�ŮU�}�P��m���vV+�9H�I�]�Wt:r�Pc��5g+r�Y�ՔU��8�� l��-�K�����P�g�Ÿȅ����tŲ��Q�xn��Sr�YP�B&t��&�l�9��;qX�TDT�]���u���M�}���X60�,���_+���"�j��60�.�n��K�woZ}�u�h�4��v�iih�6�#;VTK)*�gWu��*�]b��l]CLB��U��N�,�O]ɂ����b���%ῗ
!��\�Gٙg�^`7�q����S_R�׼B��%]���؛�aԻ4�N9�l����=3�r�w��P���e��wO�xڑ돑�j����׹��{i��C��q؛)�l]�-NDUdS9��T�&�����=�4F��>�=c���5��c�.K��+��]
5t����&!��L��pJZ�R,usf�
�:<mu�@�0��̨o�
�����t���6�K�\�t��Zj�L�̳�.ز�ra��s9&���il��` N�ބ�i�a[�7�Rފ`o����!BJ���S�NV�t���^;&�'rz�Y�����ٓ-���oɧ��اP�7�ڴW;n�� ĳ�� +�Fc#4�����U�itx�CD��;���}ݵ2��t�n�t����w��b�%8��*�L�'v����HU���a������Z�ʊd20�g&�V�ܜ��G������:�����Կ���M.���{2�ЅS�����<��+ ��r��P*ڈ��w#@�iw��4Ύ��qb8"t-������W.:nTt��RZ�sC���L��f:�aouZ��at����slk�BYI��gv.}�ʖ�����D����߱�;79ks��^�y|�n�v�G����������6򹺶	h��8v�ybĬ�#j�rP�)�`��od����{x�,��u�-�n��s�Y���k�+fP{}�(����S=@nT�+a�#�W]JYh�H�:�y�&r�TV^��G7G\�w���[��,KMp=�D1�|�J�+���k5nd]��T�]M^��z�b�7���eC�Ƭ��B����aƷ�B�m��vl��ǳ�U�e���!�}B���n�V=�V�Yu![�z��e9�a����}?~~~�����P�+�
Lc��%�\��H���%(k&�;r�P�%�HX�b�! 4$�CC`ѡ5�wy�K�r�@hԦ�F�κw]"4�	/�]ۉ�b-@�5	�d�Ir�d�O9ܨ�(�DSd&�B^wR4�"F�E�`�J0��	"�G��h���&Lb	'��D�	)�ΔdSD��8�ɢLf<� �����K`��1���F��;�dɏ:�I��i��b�a�1�u#&`�a$61�RO�(2F1<������.�Ćњcb
$@/�!w]�w$��p0DQ�^.(�l@�PI�F�%�j6��t)&�q�"�;���ݝV>�ӑm�$��{¶P�G	�.�m=Z\�V�:v�/5�5��e��d}ۀ�5.;jJM\��7���ngL��<t~���:�v�)<^�Gl�wܪ(3l��F�9^}�'��{
P&���q��6^������:�qQ]Ԅ���h`�<�h��*�;:�r�<�[����2W�6��\�a��rt�Ax)��H����0|�ւ��lx�������U�F�����C�	Z�*bz��|���D	�`�����h��3Q���ˁ�j��uz5���^�>��8��'�g���� ޾��s=2��d6F�=��A���]��|j��%�C��!���_����}F���=�� 7��N�ɚR��Qe�Íw��DoE�ۢ.ed,��U��+��]�l���7�.;�w;�7%q4m�P��FF����3��{�z_�����k�n�{�:�����mp��OMƻ�����]���]'�\���{��14��f���tfO2�i�z��9\�u=��u����=�x8zWo�����w�}�G��_=�ZB��_�ܘ ��vw�ݚ�;����>[l��\2.3cMGgD�������yS��,�gN,uO��I���� �o��5�@�/�Y��"u��I���=YB�Uε4AC!����mܻ����[}�*��B���S�����Ui��΍��o"4��9+6�r�l�#]s"�grEt[|2L<PNd[�A���w�?w��*�����PY~��,��a���P�U�I|J�Kz&�����������G,VEé���)�b��6�B��/䝻�%���Fv�}{
G !���:�e8�[͙G`f�ٞ��0�q+��������wq~g�@p;g� �x\��w����]N.�{��qS9�Z�7���������8�>��\�9{�>��}�g|�͌=�k+23RY����$��� �A�G��+���,�sBr������z;h��g}��gc�JХ��6��0�\�5�,��`X)(䤧�L���#��^9�@w����׳E������W�P>;�C���f��DU�p& �ZM�vW�F"!3}�5T)U�]�VMMO�I~v�w/N780��u��LMC�.isG�����A�.�{��N<Fy߬o<q[9�Noq��n1�Q��[gǧ�{�t�`7�����C�%�����;��v_e�Ў��)V
��SGF�{��F�mr��wO"x�:g8��>�$'{�5��𮬨3���::�卽kq_w9n >YR��:�e�8e㮹���H�W�L��=v��칕1u�]���k�,��m-�����K������v�u��+`�4{:�� w-�wsR�6�/��ŮoJ�dn9B;w����)-�1\��h��G�	�g|6�
:�	����%OM�����w&}F�����~�F��NnTm���td����������K�k/���i�}�m1����������J�Hs��:����F҃rxl�7:���oz���U@��ہ9��Va�R���W�E{��{Ր��_=��O�{ù�4}�C��v߄��ʱp��#�,����\l�T9��(�Y+4��	륌����
�O��ϧ��F���{�� �����;Y��8���L��ϴg8��9o��y�r琾��R7S<�Dap-r��3�Y.�3�ʣw�^���gOb�]Q�v�6.���0�3�z&|=��EK�����>ɖ������>�������ͧ��L�'�\�$)=>1л�<nΒ����t�qS<�ֺ�i�������c7��{���L�z�'���G����נ��[�n�t||eSJG>�����K�!Sц����MU�^FL�i�N
G��C�����>�N�p.J5�J�3�U�i��<�ʦ�פ�8�O�ϑQ�ـPX�(`��$�x�oʒ��tܸ�J��D$hkf��%9q�X�Z��tKN�f�ê�#�k+*�o9��sgL���K	<�_ݓo�;�H��ub��j����j�R[/�R��N@�]*Ի�{,�̓���㧏�I�'��ډ���s��w:@xW�Qp�p(�� RC}c٣�l��r�G�B�[|��Z+���#�|�&��<M�XTC�WgT�lt�3_9�Y\�n�vr���S�Zso�׹jE�p���U?J��ll�,cȯ��Az_[f=����}�_uA���D��=�F0x���y�	��#���_uLr��DĔ�кN�`�眮F�.W��GO+<n�A�i]�:��Hq.u"W@U�P�TMB2�����{]F�����䩎�����9�U�ǘ�[��k�v��'��x�Dq�S���v�����TT���8W���&d��ie���H_�����ܲ���ή�������=�oz�SĪ��l-���U�x<����mU�+=���sT�7����}���q�,�����J�ڼr��	:���$���~|W����OIӚ_�UΦ�z!��\^r��W��晑���U\��ß��Q�MY�3�'/�a��nO�}*����i�W��=�w�����BP1J.���W�ú�r����M�C8���`u�%b�N�#iS�k��|�.b�
,)8�Ѥ�&r�B�Q�}+O]b�9droMK1�|�細n�\��3��`f(&�z�Mt��%gF38<E㡂3����,N�R�'��"��[�]�;��+�c.�p�<Ne�f��,O��ȩt/F`W���G����3l��s��[5�'�\��M�u!�}���YS�������Fv��uR7Z�����y��g+ss���BC9�EǺSs��õ�Z�բ�o�F]�$�!q�P��kͳK����m�sF�y��NT��u�?}����3�qy���S�熚���R,t�!o?x`�y˳�}@F��tT�l��Z�<e��9��i�r����l�wܪ/��-���O���l����NA���΁!Jfn�e�F;����&�{��y���ޑ�\��}2��No��3�5�U�:��F�� e��.��8��J#Zz{�����l�O^^>���ص ٖ��9��{������d�_" 7_	�beum���L�cY`d35=Tj*s^>�2j�E�����[�'�uh���镑 �l�${�{]ET{�#�@����7t�˯rӗ�����f�[U�{��/��5��X:�&Qd��3/������?k��^��v�;�}ni=��ՠV�#3ƣ�[�+w�7��#M�B�VCH������5��CC0��_��U��\�(i��-滢*r1=bF��̗Q�ܴ}�A�[�h˙�U�\��H�l�K�
��}/�]xF��~�M%
!��蝸ru�2;[H�t�p'?+���/Mj��U]��Sݗ��wF�J�h�Ϻ���T*4�̝y�W�g�������Q7�G���4�RW�����_�V�����1�}�n=�����J�Ǔ]�z%�ѳ=Ztz��a�����V2�;���8%9�scv����w���]]��?b���%�e���(|�)�7V%\g^�fϣ'2���9�}^��qR��-� �+��ek��*��9�+�g!�./к�f��\;%�.W/�
�Yg�:��'���^���T��Pq>��+�R W�|�U:ܟS�Ųۜ�m���N�\�(e�2�u�hGn���fJ��>���S7NTgѳ=�a��nK�ۑ}q�W��q�W�z�LX��Q~}�m��|����izM{�+�����3�\T�)���t��}V��p>�_�ql�P�r73�C*k�쇋3#˜�Q�Ӈ��F��$�2�����R�q�rY�愿�������vY��rtwݹ�X�tC�5������v.J4�U|e�"E��IO������#��<*c�T�������O�Y��/&��,�O��e;��Up��\��W깋��9�b�%_��ӹ���.:�+�pc*��C;��2	Lkzv�WK��Pp���빙[�>�^!z��5���#L�����j���^������q�75�;��ef�+�(t�Q,���`�ZHҸ�^z��a��/*U{S���W�4yv����|���Guh�o��F��T��9��sPzH�f��3N7x�l���Q���xt�+2��o5q	��|z}����9X�~����$����h���J�Y����xz�
�B�O#����q��F�.W�n#�y��zs��s`G�O`[�m���SH��G3����%6=.w�	��*zo_T���+�1i��F���m*�t���g��V����
r�k���W�z̓H�;Q�o�=�-e��Վ�M�3i��Ua��F
�j����|�$����)����o��X޹�s���UL=��aONx�E)zyB�y9αF��.�g���=sw�<;���{�������^�	��顟B�T�ad�"�\Fdø�X{&�k����1�T��� l?I��˾�U]���֧���N�<���\�O�e��
�{�8v5��l^��=����V'Q(�����w�L�O��2������k��y�~�	ވ��*��" ��赅Wt��]�i�G_s�eXӋh頞i2�Fۤ?8
���>4��ji;-���B��8��!4�u+���p_>��N��'���H�y�*\�#C�n��u!8��f ��M�=U��L��e\�/~䕏�v#�%%��5�p#�?rڬR�W]�6���]]�g�G�0���������
ׅ�,S�1�{}S���-\A�=@Ζ/��g\�Z�=V�W�\v�zj8���w�QU$�Kcܝ6W��9zޘ���F�A��DTĦ�q�c�ʞ�*���K��_o�Q�B#�x=�<�{��!��[���Т�GЋ$�3�yT9����������fۙ;W�޷w��q7<��9��;ﳨ��ʈˇTÁD�@�
�紼Gz�k�^���)�P�X��h�sCȪ���'��<M�XT>��_�����i���3}��GU)��	� ���!��"g�h1��c��g�Ʃ�}m���m�s�p��ȿ��~���߱��a5?�ӈʭ2$i1�FQu����B,:�ۑ��[&�ح��^��\�c�*.r����uG�S�Q4��;��;����K[6���'�3�fɠ;�Y�)P5NF��wB�:�{��3�q�T>��k�,��d=#�c���z��a��߱R�ڤ�)���z��b �Z���
ܷ�ԥ[����j��%�{+@�]f\���\��G\����k)�{��z!��q�)j�U�:@���|��ހ��jƾj�_D]7ov�Md����i3k5XbA�\%]&fي,���x�W�`���M����WF�y�����i�w427�R)�T�19ܾ�<lW�a�s�ǉ��A��g�5F���v�����u��t4;�����OU�Q#n*w�qY����2pm�z�e�*zN�f��{m�s�=��R��9]�w2��Q�kf^�x�?WS���P��0b3��J���b��ճ�S\����� �󟣇��.�ձ����<�a�B���3�m�߸�i���_��-�ȱu�2\��~�L��O���n��樚�s��m��]]�}N��/�P������{�^���^��|c[���^]�j��.��]j�;��#̦���×����ž�w,����;�y�yP�P���##�m�tgQ�fQP�����vFt�/=��}θ/D��+�]瞮�3ħ���55���@O�Ρ\T����]e��:�v�'����,�T<��L�`��i�3�Շx� oW�X�3p6[,{�q�wRs�h`�sζ��^X�l篫��No�|u�cL��w�2	3�9�c3�/uú�����:f;ck�
3��gf>�`�����y[Av�h��[���k�lf��SWUͦ�b�2�s��.� �;���9������iL���Vز�]��$Ί�M8�I��w��0�^�ߓbb���jw�3���,��	Q�qod��s�0|5�c�A�]�v���7~���bnk�w�W����t�wT;]Q4̖i��:LӴ}[-ڎd����������O�(����H��:a��D��σ&�}ՠ\u��ә�`�l�$uW}�,�*r����|5H�o��S�v����q��F�6���wR�k�ހ� �uNLҖN��eMz�9��(Vn��*1���GU��^>�o���{L�~��ѷ���/�@�A����Ϻ���W���/�ƦJ1��A����;����c��~ͧ�]]Co���c讓�K��и�r7'��*P5<�{^������d��za����*{�N����1�����yYjG\X���ۺ˽�ɛ����n�r�M	�ׂ�ÿT��d$�W~߯�Y��a�`�j�!�� ��xܷo�������u./�.����He\ȿB�Ne�f��0��p�>��\��T�l)�^�T�i;�W +ɻ"�N�'�S�ų��h^��h_ا$��\�(e}�(�#�2ǫn�"9z�n_�Um˹�-+P�()�&qG��9�rN������N�a%��>t�V4��%b5w&��^�cz��>��7E�YK�9M{C�����d#�슕��j\�ٜ0f�=���f�D��q��� ��5;is��٪o7���}\U��F�,YLk�Ԃ��7w��+���r��m�^�g&$o"��Q���l�j�\xg&�������J�5S/�}�)��}�-ԁ�wZ&����xk�X�49몂G5̤��ݺ�%X�P�f�h�����Y�ҍi�A����/�큕� \z��`��K `}��Xwm굪�@��,�7¤�y[��(�H�Ȫ�{œ��)r����jb�"�K���
�[o�,�b��-]���sB0��ziӡp*��%���PXZmGq�<u�D���_To��KDĉۭ�LP���o�����[��Gi�g]�$��N�n:'(/���a;�o����ݶ�^��}�W��V{��H����A3k;�u��&�u���^n�@u���ZJ�9���b�V��Ł[}J �;�!C�V�S�h�߃��#( a��bb����]��p��Lj�/#w}���E���΅�~�����lA�؛�ճ��J���ޝKu��މ�un{/�W�5���mC�t�q�QQћN�o}V��(�hu�'66��[T�,9����B�l�w8�e].,�4p�c��1bB�o^��F���Y`YQm�ƶ	̋�2w)��[�e�H�\V`���sm��/���ܻ�Ȭ��k�����&>��E]P[p�j�X �ԍ��c::�nŹv�K�
E���4�[��sS��V�X��u���7�dN�h	c�ʝR3V��e�����/-��T�H钆ܔg��7`�^)s�3]�씠���j��U�`��ͺ=J���[}��λ�N�X��_Msy"l�^�9[@9�ܱ�=T�Iu��r��5i.h�8��	J_lб����v��L]�D݋�7�;�jR��	�W��u����t�l�LT�@�R,'F�qu�B���s�q�'�ޕ{;����h'X����B����1*d�Tn��8��D�=U�c�-���r�4=<�����Nh8p��rĬ���=���㢸��L����"���Z��V;/��F6n8xLղ�h ��s��>�x^ޠi�G x��ک��x0S��wb�/�u�`�g4��0�M�0�SzމY���u���f+|��S����4�gY���H������6 �?K	�Vzt�	QRS�5ceT�3!���`|�C�ʽ��h�(k�}y�@r61.��n^��m���z��k�m=�r��މs!���xz�7]�2��0�4;��1�����p��ȱ�Gi��r��'9VC�sUg���y'��r!���J�-ӺƯ���3����{S��|',w�
o��8v��Ԫ���<~��'��PO�u��P�7H4L���țBw]H����R�4�ηF���s���La˪���qݣ��^5���� EC^<��]�BJ�uwq�w�u�nF�8�R���c�\wE�Cy�c�pt�]�5.�u�m����u�j �ˣ;�N�Q��g]�I��Jb;�;��8�.�C�"(n�E2���.�x�#O��Weuu��J.�0Q�n�)K�u��u��.u	���yܡ�x�r��S����#(�"(��]��*�]΄�-˞9U�;\��Es�ú�w9��(qwts)���j��u9X��+��wx仲s���wm�N�ܰS���r�r��W�͍�y�xƩ�w	'�D����/�UP�-<my%xs��֘�y���F�C�F�c�+++E�!��w7>{/�e�0���֝|�Tk+��ɕ�Ո�T���e�������8T��ٞ��0�q7��������7��h%۞��o�;��u�נ��2pt_I'�e��T�)����.n1�X~�OW������lVG���M[�s�W�ht�l��}�i�;�<i��`LȱT�\}�E�����C]|4Nsq�]�[x�tS�j%���:(����o�ϸñrQ�G�*��D��䤧���@�~��b���ڼ�A��x$tOc�}�̬ޡ�\{���:�b�P��ʌÁ%��iߊ���{[��b������9�F#q�\M�r��y]գI��u��LM9��r�N��~c�lR���yA!��#��X����&<��h�m�}m��i�<}>bu�k����ᗺE��շ�'�I�=�QH�D�HU�R���Ȅe��F�n!r��}�Ȟ>=9��^r��h��_*\i7�l�$0��A��wk¾�;ƅם-7�鿵�H���Lg�=�vN���e�{68�y<h�����=fIA��fA�0�%���u�oٯ�N�}d[B�c�Z��S���չHK]���4e{�p��nƦ(	��z,�ܮ�B����N�f���r��r�0N���B�����w.�f�kje���mQ/��^Q�n���}K���!���f+r�����͝��N�V�+�&R�n�_k<�o����H����o�����������A�Ĭ��{bs+����y>���ܳ��y
7�7���h�ܿ_B�GH�:�o�t�vU�W���%�� �.;zr�+����yYs8�9r�+�V#u3�N-��{��Wi>n�Z�5u��z6Ϥ�ϕETv�H���׏�y�8w�ex��>�ÐOq(�A��\�;Φ�'>�ew:��o��Ql�Q�z���ߦP�Rp����	�
���8$��re��0��WK�����S�Uҋ�>S��,���r���α������fX�:X���o��A�����z�,h���l��Г>��Bp�G����]!��oLR�T�qe�v�3�T���G{]v��9~w9����\	���﫳�#�u�΃���HY����&���䢃$��0�qQ�i��M���<�3�js]��+-���uݷq<����s�Π��ܨ���S��TL�A±�{h{ݙ�-�| ̞�(	�%Z����F_mD��ZG��+�<w��wYN��0:�Ӵ]\�����]͖cX���Bf^d
��2��岂7(k�S2�"�aʍn>Ea$7Œ+:��u�!��$����m�y�_gs�{�V�#e:�a�I�K���oz�=�zS�n��I���(S4g\��8���kY0����f�hbW����Q!�h�ѩd�6����%]E���?�L�����x�"�[��/���#�J���ُA�m�mځ�Etץ߭=�U
.��k���22�eI��m?I\���t���?������rm���(^�vÊ�<zq����@�N�j�'lL���1Q/k��zZٸ���ϸ�v���Mx�$v�8�׻G�;��B�]ж�q=��<�:����A�,�������T.}��W4{�7S~��TmY���)�v��q�o_e��s��o:�u>�OC�����j�+�������x.��ɺ�C�F���Y�������zw*���h�P&��'z�e%�}WD��T�{�Z�2x����}҂����W��]*zN�Fl�7�w�S]���.+[�5N���(]�M��{��7�|n㓗<?T�O�����>ܖ���๊�}���]�j��n��u��S�Ey�X��+�b��z�
�{��E��Ma��@rx|6�gG�x�[��Z�^�5�5����[��}�WWq�r����/T�<J@ò���~��h]�`��dǋblۙ�tr9��σNՕ�Z��Ӈl�8OF�e�1��&�F�;V3����5�2��_j�m����Fu7o�Q����3f�1Vk����%��^p!Z�:�I�S���m^���ʉ(-�����LY��c��އ�&v��|�I��l���P�j�+�nȸ���}}\9OR4��P��#/�I���/Mu��5Y��������Tmќ�q��n1��~�OWa�#����S��\�աEΦū�h3�7瑙�\I�}
xz�t		Tu�L�<=j�t�X�n�
���/O�d��/k S5){����Y]�oY�5�|f��l4���,��q���aF;����&�����e��Փ�ۮ��*Eɖ��wH¯��'.:��v.K* 	a��[� i\�ə���zWE�^m�{�=U����������������cs��I�uAñ��L�f��:LL���^�<><��Տr�������W�zF�����Q<�σ&���Z�����g�U���c�n������4˞#�*�7�)h�Q�\o3Q�ھ�wu z:x���Pꜙ�އ�N�$+p�t�M���e�gg¥�`��Wq�>�)zo_e�z;����&���y��I��YwW���6�l�C�˙5���������T�8'�Q��޻���}v�Q�i;k�Z�&�<x��]{(1�򷢬��b[�a+\-����G�r�S2탁�C[�<t��Y�Z����Sv 4�Y�J�9���g+���"E!V5תw��7h��:�b�[���ٌU�4ѣ�k�Sm�s�h41�mS�{Dd�{#R_��^R�ʵ�ky��$:R�'Souz�i���ĭ�za���������I�ݦ;8bN�r��Q�2����t�������ܪīμ-ߪ|p2}�atx�q^��+�l�n�ɝ=����
�~5� tg��:���9�K��B걚}���Ű�)d�\A�~"p���N�V��93��m�t_R�F�y�2�ɺ!IƤ��Q�gͺн��/�S�u׸S~�\�۝G1���`���I��3�tꑺ�p9�F������������q^��\f�N�
��{{���8�=�˧�x]�$�DL�ugC���SZ�7��������P��ר��
�8��{�:�~{��E5pע�MB;�(��}$�`�,_�*�W%��)��>�ت�U����^|�>���({�h�ێ�q����;�\�P�J�,	"EA�IN�O�z��˖T�t�tM{zJ��#�%�^s��VF�*��u p�C�P��f��DTf����v��Ձ}\��
-l<�Ȟ=<�́���>Wq=����qwV�&��u��LM9�玽S߿��J�͚H�.�]R���"�
[�';��;�K��s�򽣦o�X7��;���\t��9ϩɸ��nT�G^��E�������c��Ү����,m�:�ˎ��(�����������fu��R��ݭ7;��}4N�]]16���iʇ
($��3�u| {=�/kA�<�y3Q��4j6��l����=Ǐ����+XIs�>�ޥ��B�L	��=�%�S���&{�
��SGF�_��m�W�{�"x�$�B�:��OJ��PR�D�ٰ�$t"��A���k���hM�Xov^��t�}��Qӗ���P�=S�&�G����==fI��d�x���1R�^Ec��v��*6��6�{׷k&����w;��U�:��;��;|������A��x�Q�lNa���h]>&�X�t�j��7������"#U��{���=��G�c�e{���7ݕaŰ�d�q!~Y���9꘳�C^n�3^�c�x����4n�^��e�1�ֽ����ڞ��nV5�]�Y)7����9~�(�8ɭ���×/Ơ����8J�Q��p+˝�92��/�u�T���w�%mf�AP���/s��pU����p����3�I�82"���>ɖ�끞��.[���)'�iP��e��N�;�W�u��{}S��'�,\��S<��k������o��W��ڄLT�r���X1�h�|��Wm��v�=~U����rԈ��1�U�,�s&[٦��t��S��_���naiɖ33Hj	�=~b�P�1�ث��>�g�t{zō�Pm>�"�3xt��ir�F�ӫqU�D��j�s5h>��At3���tt���uw�C����[�h2N��a�*�S�M�e
�5�=ۊ��cH�;�9u����u����<�{��z���*&�B�rQ��IZ��_�[�>�b��3	lz�*A]Q���=N�o*'���Ds��w:@xW�Q�XeV�g��X׾ħթB��o� ���9���~�uc�E>Wq=֑��3�+NC�T�j(� �]�i]���-�M�]5�j#�AF�A��DLD�Z��Ō�fq�Ʃ���c�0=����vUm�(� ٞ�z:g0���;}U�C$��U0�l��+�и��q�Y�:7q.`��z�\xɪ��S2��=�/ê=�t�&�F\��3��;�/k������3�}������~�7��ï��r8_���nx�|g�އQ�2]�5
Y;P_������CS�5S�Wȃ�1��Hr��'�c���ѿ�u ��py�q��}�����m��W��/R-��}$���3pr|����{O#��/r�p�	��8�@�/��'(���jz]<�F����O��쏕��d��i�ޯ5�F�d�#�/���Yip�g�-i`��Ԥc��ÖxF��̧�܌��ՠ֮��C�em��f�`�)����3|M�4'���b:����u$��J�'��3�:��7[J��V�Fz>�k�jK����-+���x�>�
�d�w^�q��:sK���n���95��*�����yt7w�~�i�6������˙���8���	*�[L�T���G��#�Y���:������+�wU��r�F.3ީ'��E��Ma�����h�n)D��
]k@����v��}]]�}N��>��H\bʝ7g�J��?[��S���-����j�s��UL�5@s�2!o�-�e78難/Eu��z"}Z)o�FG���)/���x�Y�K�k�����hїP�(�#:zgc�����Wѝ#��Gm�r�W:����ѓ/�;��4&踜�����ҁ'j"e0�w�L�<=��7�7V&���>�'�ӑ�[�U���}Ð
.�k�-�{�6˰liA�`O�J�66[,{�q���HM3j\�Ό������
Dܻwvu�r7�aW�q9}T�8�YP I|dŽ�.��9�
 ]y�]�#GX�r�ě��}	���<{�ln}�[��{��鿺��i�,�" 7Bt���X�3�<QYC7u��cKU��:R�
���5�4���-�c0��\��G�(�C=�Gl�y��E+N#�����O��mE2T̫��(���[Q�z����m�7{���LO��������&;o.���55�ұi*Q�ܲ��qڅ�5Q�����f�ݙo���Ȋ�T�kߝG4�~���wפh�O���=ԉ�G�d�����j�L��&�"�{��H�f,U'��<<T�1�*7Jxe^���q��F�j���wR�������3f�d�����wO%�o���ĽRg������¢{k]z���J^���q�j���<����P���L��y7�A���/X�_C=s&�Lq٨>�p��_�s
�k�?��7��(׸�s�gwO��8ߕ��?	���J%I�T����ƞ�J�0�@��ฤ�I��F*:+��v��ڏTպ�]w�����������UbU��x,[�T��х��3�O��C(����v�R�f9J2���OENփ���`
�7|=��x�DwR����f��_�G�d���z�.�q���S�R?�~��#���~ʟ�n�je2W�W +�&싅S���S�ų�mօ��hw���2UmGL��喆�,~H�@�=I`_U��zg�P��G��MƹL碝Cgg)K�;,x�<Xҍ�9t���U��ϖ��Jb����L��gC����1u��sx��?F��z�GI{t,��pt3E��0�/�_�����`�|iت��|��E�Wu-P��v���]r�,xE A9�2��½�� �%���1u4'��I�������u+��g���>o��&Z�T�56C�ؘʳ�ř�p�qAG�l;ڂ�6.�� _���ܶW�+��/���w�Q�rAڃ,	�y.�R�J�pE{�U?<��s�>��BV�1�9C�$�����g�a���IXe�?�#�qگf���3�{3mT�V��=	�AW��$\�����s+7�aW�@�t�Q,� rێ���h~]\�ML���ڿ�M`Y��^g��b7�\M��/!�ޮGs��Ѥ��H͈�'��7�Ldَ�+ش*�N� l��vH��[�4�{���o5i��|z}���t�`9���AI=$@���_��nP�h�}�$�o�S����/�
��M���q��F��}D�8��Ɉ���P�u5yo\QQs�d��zsI��Ni�+�Y���|6�;ƆW�-7��<Ɣ6+�5} ��x��U�3�+�1q�����z��ut�W�Q/�>']U�~�O��ɂ�ΐ�����\��ˁ��Oe�������=��y�M��<��9����H:x���n�zjůi���sI���3�R��qJV�Y��hܫ��{OF>��������+��pJ�mϾ��WW�&�k�.�S�t;q��y�vz���J�l���HHVˮ����E�}���|�W�c�ވj{���u*�e>��AVnj�:��2�T%:T(T��y�|����<ݥt���msG��x���fj�Ε�{�ƙ�;�K�}�zP��^���z1E�0&k��kj�X
{��fU���M[u��T�V�=��Y��л@X�g9�!��7zcK�V=e	i$�=�G:��6���@�o�É�ӷ�u��f�̾��R�&�;5����Z�3��
���u�����H5�2�V_�
�ˢ�����;���r������>�V���]ރ>R�����-fӭ��\��0�\��;�"�8�p[:��䍱/:��̂��J�Fiu����<��UtR��F*�v�z��V���A�郹(��D�$)��ݾ�f��bZ��-Ò��m-s�6rGy�r�#�JÊQ|+}�h��R�Y�:�w���Z{�e�Ց�ݕս�c�<n�[�*��4l�Ԁ��y���ڍ�=����\�:�$�(�
��r��E.},�Q�-����8L�v[CH����1	Ġ2a�����[�%dO0:Gkf��pLK����ׄ)I���[�6Ѱf��`7[Ρ��H*�Q�.q;yBd;�P�z݌b	Ң([7�������
5[I���J$@iAՋ�̷�-�5����!�=�K{%2G-�9|�zѺ���UV��7XZ���.xz�=�t��!OR��"{o�-4��������t�V�I�9�s"�]��sX1�M��L�G�+�]W�b2��.��c����Tz�>��ӫylXW�`0V����t���ȸ�f��܊��i���6�Z�3*3�Վ�X���-����E���@0^o6�Gk�g�=7_�[�Z2��-ۂ$ψ��x�&&�ͻآ+'�,[�]��ϖ�2��vz�`fd�b�A�ʕ���}oz*
r�{xy#��f�<��r�;iV��`���uQI��66��n�f�
J�������;���	ӕ��e�x5�y����Z.��q_"[3��wF�����m��7e's�آ�B�3�4�W-5����lB좆����:2��W�; +t��C4�v��Z�k�UwW�gZV�>��.����K�ݲ�9��e�-̎G�9e�%.�9��}n��N��L]�O��$5��f�]L��ۏ(�t�-�9B���jѮ�]v��9)�B�w���g ��
�޸�k�3o,`��Xo-:�w�Fg6�<T;�r�(g*V���yଦ/� �E2j䭏Fm�gfLO�9Ǯm5��Y�p���[Ȩ<V�o-sCh��]�Tv��]C�䒰��CeӁo��.��t�5��h�R�%E��V�e�'������܍�+�֙�v;�|,��/�@:�I��mV=Sn{� 0Q �R	 �$�{�����rr��r���$���s��d]�W,�n��sN�3�Ýe�ط<�<e;�C��;��n���Ww.w1�ԗw�s�\��ێ'j���G9�x仃��1���rEλ�wWJ��*滸wA�Bt���s�F-r��r6s��.]�sr��;����Jw]��s�����ۛ�.��K��WI5�wq:tK�.�t�Ÿ�"�ݢ����s��k�uws���8�����je��'u�w]']s�$�G7:�K�ȇv�[��ͣ�.�;�7v�w9ww;5���WH���;��1��m�u(Dp8�$�v�s�]�wq��n�]�.��N�N��;��WwW\����뻣wdq�"�p���s]�DI��t�k��q�\�:\�ۗs�K��:�� � ��gȪ�ڃ2��$�� 䭙���S�وi͠�rz�t����;��$����+�i�V�P��n̅��$U���gV��U�1��Q�^�F�{	´�/r���Ϊ�@����b�q��j���?Pi%����e��W>����p��8�~��V���ģ�K�Q�����'�=������xo�5����+��Wy��W	z^���X3����%�n�Z:S_��)�1�}�,�S�"n��}�}ԕ>�`�>���]]�}M\f��#�Tῢ�'��c� Ζ.�ykN�3��̼��F^8qU��ew�O�:��wWq^��C��ޘ���F�$������gi�(7�B҅�.�����3��+�=)]LwW�gD�9��!�;O�ntq�88J��S6���7�GZ{�~ѹ]�O����:�:eqj-���Wv�M�;�>�'�ﳨ��ܨ�������I���q�����*�@�Q%����~�V1}O����ZG�3�+J����^�9ٞ�ކEEpF�䝑�5�k�25
ETOQ-փp6_3!��n1�AJ����	?O�<��Mz�����>��1�|�q���o��pv�����s%��U0���"bJ�4.���k���^���#b�f�l��>��|����v���3&]э�C;Ƿ�S�K˞%z�w���q�:����{'��<-��)�*��t����423�`+/Ei1�6��/ۥ��(]n�TJ��^�<����Nٮ�����ﻕ�ێ�|�O+<}���K���
t�&��'o�3�N��{<��<<rSC:N8�|��R�ݛ�T�o:��Dw+���{�`c��0�R��v�\��:�'}����h��^<w�;��}�d�;~�ۇ���_}����Π[��4�;����n
W[��g�:=�'�R����A�?o��~מ��;=����'�h�1��z�@��K�w��t�E�ԧe�?}�֕ϵx,���1`������:}�/���GP�M�"�z̘��mhw&n��c��Sڨ��~��|m��G�N��@����pIS��{���UWgg��ז�	���۾����r����uX����1q��7�'2���|'�a�o+���}����5����gF�<�>2��_���;�t�i��.1eN�JN�����b�l艝�X6:�}g�2�2����V��"�x�d\y�nw>���]hp^��hV#�� tzF�����N��=#:.x�ƾ����ʨ����p7��?F����Α�磶�OM���躨u D3>������_��F�Y�I��"������~�N®+bJp!n]��u�_��PP���.����YU��:o/|2g�C�-�!�AV�KC����t�%����Y���ֈ��\�S�{�������2�^�X��6�YQmr�ؚ�-
�M��_O�GX6OT)`��2��ʡ�T�s�֮�7�7V&���;�R'Lzt�a��J�E),�l�Ϥ���W}m�@6
4��ʌ�& )\f��e�c��:�v�} ƞ��7�������==��>ζ�oH»:�}��LñrYP K>2�H-��+��2�}�zJ���V��ּ����rw����1����{�����cr;�t��w\7�WTK�����Hg��&]��������h�[1"���xפh�O���=ԉ�}�|6��@�� 
��Vc��m>f�}�#4��&^ӣ(�r�+���7���m_Q��{����͟��:����̩R�$ې;�Rf��'@%��¢^�
�J�u)zo_e�{�����/�\�m�F���&�.�{�:�Ti�4��(n}���X|2���f����#�^,�y�"j��:;��1��讓~�p���7��g��O����VqS�pM_GVoL��o�y7��N7,+ʯ;�]]��}#zS��U�Y��C>w��x����m��O³.���.5��QXtX4����iz�(u��ZU��]-�X! ��TAp�uu���H��ݫU�5���5�^�J��~��W�l��_D�<�M�C۽V����+S�U�7R�q����b�]�-�0�����3�tP��Ч�:�t��bۑ�d�����Ɋ�a~���w���|=���3�;�oMaǓ��s"�Q crh��������7�No��_ڎ��V���%{���ݑp�u�>��F-�6�B�
��B�l����3�>��.Q(e���څu�H�l�Ϣ6g�;�����|{|�k�ޱYu�6�'c�Y���7�On3}������/���2�A:�*g���V������n�3��/��+*oٙ=�[�L�z��Pea���+�\�9xϴ��[�����b�U.(�O�N��^���,=�X�&|��觕bS��}�Lgl�8��w��3�0��pp���=vM�=3�~F��
�n=����GAr�g��A��6'�^Ds��VF�*��H6��;�rY�Ӻm��Mxv;�x<��3:�'�vW��<��+����y|{���t��W�����Y2�E�W��VvǶg�^	�S'g�����[���G���#�c'���ǧ�{��*�u�����z=w9�~��
2�k�@�L�9�Z7��4��}HU�ԩ��s�e��F�m���Q��θ�/��<�|�7Ù�7��w�&�2f�j[~����gt-��O�_��$Zyl.�Z�37�l�!�aﵝ�3_MS�s����Y�m��􆶦ұo��Ɨ(� Ԓj�
� �.�O;/��(p/+֧���/	����8�g�Nq=lsL��;9fau���;Ƅ���w�7N�����4�G����{27����M��7��7��\f�Y�k�Y;0�>�1�j������\�F՛���R�Zo�f�q����C}wB��Pu=ǀ9�������A���%n�3(�U��,[u3��r�7U���J�S��t���ϵ_����zUr>�}C��v߄��ʱ⇔�b���У=*���t���|6s*�z�%�>8�_��w��:��'��kRX�q�O.
�z�8�%�}���OEhܭ_�Ã����z|�2�]��Fc˝�<�uC�&�����]Bn�|Y*�i��F�}�Q�W3�I×2ǫ�3�\T��K��O�N�����z��-(5�s9|��O�==����o�u��{}S��y��:X�ʒyO^��>���}MPҽz�?F�\{����wWq^����i��2��,��X'W�^ى�N��F��Ni�ۨ*R���{���y��v�m���}7,��?zBH�0�[ѹ�گP�0���N���+� �*,�Ý�=L���є�����I�5�p��{iC��z��*�{A%|-�C:�n� �e�
v.�N��tw�l!p�r�p�4�4�g�R�n�]X��&*x6�]>�W�N��X��^��^ģ3V�C��}��U��?���6^}n����w�}�9<�}�@==�5T��Z�s?_�:�n.2���UHu�6OR�SRX���e�X�}�\M���i�7�g�_Z��)H�sE��_��2�i��s �P��UOQ��|6_1��R���B(g�;��y��'`��r/)���m�s�s	��u���2+�2Y�S��\���@�J�Ռ{����2�{8��]�w��<�+���_=<����d�@�@�N�k�e�ۈ0�hL��xE�F��3��s�_�s�e;^�R�*��ΤpQܮ�[n����7��O��{���aK+|�QIR�6�@!#�}QQ/k0��{�߾�ۇ��_e��sTT<�����4��VOޛʿw�_A^Pt���� ��V��6WVa�/Ohpy�Te���O��;3�B+�����d�
JU1>������ޙ��Q��a_�'����.�='O�6_��1�]/m5땝�G�����;�'x��+��q��曎6�����쉞��R�;Y�=�h��?iB��-Q�ә6�H�ې�����ln+��,���[��h���j��I*�Jh����}u�R�23`�<�q)�HJڬ�$ɩ��9{L^b)56l����
�:[�\E�^�����I]��?���VU��,]f�=�:x,���۲70��������8(uK���uo�4=��z�^_�p�"�̸�0���w�n���y�imw�z`ZV�q��0+�'o��|���>����˔=��N���M��R������g������\�o�[C����X��{�WdL]؍��)�ܾ���q%#��`��cw�.6Oxt.�H닔I�G2
�{Fy��e�,�7w�F�����^I����{��2�0-��Qq��j�^��hV����$�,�ʡ�L�<=j�SubH�n��ut�v3&}=zy�/O��K;~�p��f�v���,2��W�-�W��S�y�C�J��c�2�tIN�xw<�h�oH¯��'/���p.K5�U�:�3�U�m�a����=<��}�p,}HhS�����պO���ꉯ�������M���y�'뙮�LL���q[<�n3Q��5>vǢu"{���}Ӏy0�4&�u�zo'\������D�e�!#qd��^�Q��-�D%p��o3Q���*;���Օ��t�l���z��6�ҭச���uJ�D� �K2�gg�w�[}K�J����D��/fH\�1� �R$���X��̼�w�{��ƨ;;m'�q�F�gc˩]zk�reύ+z�-_ͳ*�aN��oI�u�Z�fB'��y���䥉\1�[�>���5���	ߨs���S�����*_�������\v�E��ިw]*w��y�;�Oj��6��z��r�d���9T*4�̚�0���Cs����a�qO�����}����9��xg�+4��?G;�����F=���M�� ��i���ĭ�za�X�st$�m�/=;1(ڟw��Զ���۴�{j�8lB���c�Ҝr��:�X�w��,�ˤ8�W3�ت�U���kЦ�}����R�qR��-� �s�g���Ů�bT�7�����Zլ#UZ3��ob�[=!��}�3�_�:}3�I|N�����vE©���)�b����=�k$�r����g�����[|/䝣��=�2�k�;P�+�R7�l�϶g�;������6�1�#�����]rNr��p�^��Vm���ޫG��I�Ip��%�Қ�S�V��O{xw]��,<��rx��Z2X=�{�qx}�=�z+�� oNB;�(�[����y��J����rh��<S&���+���uX�k���oGS��<v��v��>���F�G�+ZDZ��+ߓ�������; _Y��lh���z5��us�ʃ�⅗�)�N�����r�a�B��[�B���$z���/����S9�;��{l��H0�p�1�J��QfӘn��u�[�y����^;��*-����{����G�w��OĊ*{z|�����#by���<�edoP®=ԁ�n�C3�j}(u��׻!/���"�c`s��+��)�iq�����/!�z��O:fqLt�G���^3�jM�]�Z&��J��@�I��}��h�g��b8ј̈́��6��ݳuۑ�ח�QJA�4u�}>����3_9�Z6j[7��"e�!R���6�Ɵ��w������ԇ����|�o��>�D����{�׀�4�3���]�
�\��rgE�B�����W�U�{<o���H���]ф�Q�����=��d��Y;0�7;|>�eY�mxwV�(G���-m��b����Lm�����7�t-�Pu=ǀ9�����oz��C��7�Z}�R���>�0�	�0��f����Y��h�����˪�Dc�evՉ������3�7E��*�=[�F��ѵs"�:x�����̨s��v�^�ъ_��w�Ϊ�Ḭ���Zױ�~�@�Լs�r����jY�8�#_l�8r�/�~=8�z�M���Q�L���E�ɍ�=)�]�
#Fo��%n�:���+#����y1뽵Sf���fk��$�oh^�loI�=�ﯱ!��}�ڳ���i��>�'gr�ː_ѥ7$��T0�ȥǄ���\�]>�]��WU�5ta]���8�z	H��!Y靚���Ez�G���	���u�ﻝ�^�]z��L�]'\���΅q=G�a>��o|��qv�s�b��R�����t�<�����)���ՌǷ�8W�x���J)OWnxO������+u�G}3����/ѧ����_���c=��W��^�7�)o�Q��`t��Tq�c*��a'A���]1$�9[u\E%��{��3�y��/�[��f�%2�=W�a��.g�o@�(�$�A�p$�w�l�ԝ��uݷy�x�9<�U�� �|�&�pP��:;�$y̠�%R�)�����u���l�F:����Q6�M�	�:�������=Zzϙ�9�#
��u��e��24��UOQ�h7e�c�jo�����y�Qf�͞Oi����cǽ�����nu���2%�|�a��#�.������������^5q���hu<���3<:�9\����1Ǖ.N2_�uG�W���M#,m}���g�0o�0߯?c)z����[�Y�;��o�%P���uR)%L�ګ�����o�6��[����m����խ���խ�km�[o��m�[o�km�[o�u�խ��u�խ����j����m�km���ڵ����ڵ����V�ݭ��m�Z�j���z�j�����j���z�j�����j�����j����m�km���V�������)���-�0,�0(���1$�ޯ� 4
QCfI� P! �JT��	�T �U@P P

 ��(�P�J�@�H����R�*AD���T��D��(�QHD��T�PU��U$���U@AR(�EUUJ���E@=�TT��T��R��@�J�U)$.�J�*JJQ$P��J�Ѩ�HTJ�H��(��U�@��ED�!���  ��S�[������j�sI�v�ZPA.�ȴ�*�������BU��JP�PmJʚ��J��	TT�%$�#�  �=26�aH%U]�Z�@���:(�Պ:   (���F��&  :�49뫊(�ѣ@h���h��F�(��4wUD��R� B$PI�  �zF�5)BJؘ�P�I���6�j������f�����ud��R���*�$����A�����*T�)
%G�  9@I��i��-$ձT3I�� 6iTS{k�a[CN�TmȹV�A�vv���\�hU4�(�UTRE)ͤ��ZJ�   ��kv�T�[������v�M�Ѭ͈j�wk�ĺ�6��mӍ�u���j����IZw-���Lj�ځݔ2�ƍi���QJ�(���2%*���  ww�t�e2mj:`�hmwm��������3��S@�jkq��i�u����m�7Mw;ws�::5K%mm�v]�*��[cTT�*!*�(R �  ��{{-���ѶF���;�V��6�umvզ�-�:u %����ܬm���� �`ծ�4��GUݮ��A�p� j����U�J(�[0Q%A�  W��N��G5+[j���t�:�i�[4���ik�]�vP���ӭ5���ZFP���[MS�n�KP��P�v7E�ܮ:Ԣ���EB�AO   	�y�U1�zj�C[�����
u��-�u�ݝ��wm��[m��v뺭M�̛��AX3)v:: �1U�5vݰ٫ct�tN����(�I <   ��Uz݇v'A��Wl�q\4(nΩ��q�u�Nۚ���L��m�F tЪ��ʷ\
�*�Q������Wpu��WV�4m���S�i3*���F#COhaJQP�4 M6�  S�A)R��dh �?j
�� ɑ�M%LaU5! h�┼����.b���ʆ,��X'0T���f��y����������BH@�s���$�I���!$ I?���$��$�	#	����_�:^�y��߽��oު�,��d<A٤���k�����K �9�<{A�&o�W��,��!���Ң�����K�����xq�����IP���J���7j!d�)�D�)�V?J�Y�L��X�]SS ݡ%X�n�v����j���{�UI+@{�Q �J�3Yݍ,��h^�n��A֮�kF��KN�--��G+;�.�H��4���y���3N��[j��R;�q�*�ɛ���������*)YB�p0��ܡB^�#F���l�� �:�S(��d �8�br���٩,�)�0�T�B-���Q5	���H�5S۫�>�m+ҵ��5g���	���b+1&c��Xu�oQ�βmeZ#V˨�
O^��ZbD~��e��6��6cR�
�n�lG�jY�b�mӶ�S	뺗��ݭB;ǩ呅ᬋ�CWcs�&L1*��Ǚ��Z5z�B��(r�������N���s��f�,^\�t�5LX�S����p�u!��Dt�d�z�K($����Q��+ja��ݘ��]�ʮSe]��KʝG6���D�knL�$e�N��eV�˺�ؘ�j�)���#�N���!ʎ`-틉���Y��[���<��Gh�F7I��v5)��J&�c��g)�����ڂ�h[n�yY�Li���MǤe&'�c�Vs���$~O��b$7��d:�H�(Խjn!��R�S�ln	k�T�bա��*�ýu�t'yI�K`��j��J��ڛVKAk�B���me�n������Y���
���m<��������h�bͭ˘�=H�u��\ۚ���+4��
�Y� �ݹB +S���ƃv�-|���7fWZ٠$�����^?���R�bx��F|�
v��k(��W��v3Wck@�����=��]�7M����A<�����I�崴�L8�� -7�r���fn6\A�N�nV�j='T˼	�\�y�Z�Gcpݦ������٘ZǙ�H��nR3B��]����2��Q��9+jih��m������a�e]-X� b���W�����O��ilˉ��׊�EI�&��LӒ����ۚ0Ec�aa���Q�z�i�GE�5f�ޢ�r�ix	z�/H�����n0�b�vՐ�2�n�pe,��D1,@��YIIR�N��Msua�*k�g)�9e���Zl�ծ��ʱn���FƊ�E�-�X��i�:1�l�A�e�&���k4Q#�T)����%m1�N+�Q+D�өu���J]����kui������sF�)]�F���`��k��8�V�9Ȥz�����T#Cj)5j�V�J�cL��vֹ�\�LT�Ʊ̺6^�ڶ.��u{K�/��m��m-ySm�[O �������n���z3�/�?��`��n�f�0)Ҹ7��T�xԺ�-։��5�"7i�v^X(&Z�$\(���;����6ö��lC	�y��˛���e�W�	�Q�W#��B�\�u�O��[����Щ����T��u
b�&i#2[#�l�u-�R��ȕa�Flړ���ibd����KUP��X�M���v����U:&�@�CZ�f�8���Wv��Y���7�E��{�	P��1� �:j��2͚�m��`
V�����7���V2��a�ۧE-lX�/K{HK��XKn�YD���: @�Hڽw�y������ba8��81ʻ���5i�e'wOk[�p�J��r�۵O!��f��Z�u��T�2��g
Ъ���gfao�ǳ5]�]7\y�:mw%���A�u�3�������o�vV�`]fq$�v����lPՒJ�(!��/l��)�b�՗A0�SkL�k�l�]L����	[F�f�n⦒�A��wL��.ZW̵oU�&��dD��#������sn�Jb�/b�F�k@�;�\��iM�#wn,G�OK���^L�U�:Sl!�rܣg!"l�E�ŤY�,۹��b8v���	 )�%�{��Sr�i�H3n���ĝպákT�B���4n�Z��	42�m�E�p��h�t�c�_�+VQ�Gs.�� ��yCK��� s2�Ӓ�\���"X���[�sl�yo2&�Ƀ~,�h^Be`׷Z�۰�
�驁5��Ҵ��͒j�sk�N �=X&��2l�R7v'X&ø諈�P�{�]���2
G1��R�P̬;l�z2$����9v�&�)ㅔ�ǫ-<��E��i3h��M1���j�YN��ƝՅk �����'k
WP�<��9+?I��#CkS!\���-:���\���k0u<W��vJU��Ր��o��ZY\m�Gh�T7��`��i�;��p����@]7���"���R��U֜�B�x)X�X5��e�Q[���<�ٴ�h��Kc*�n��Y8s*���SI��_�^2�+E�5�*���ՇR���ǌA��6wvmk2�|��-���G����AE��K����X�2,l�����
�e-�iY�݇��n	�%�5X��ݲZ��j=�!�fЕ�U�����݋O��J�mnpl�u��8�pܔ�F�!h�Kou�"��eI-*�m0��kEj�q钅K�W�Sh�b���[i�
B�h�wE7�Yo,�uպD�o�V��J��n�m˚4[�R���`J�.��Ӎ+ç�0@1+�)����rVIA�p$j��d��ٌn������oJ���˶&sv+I�9Z�⬤V^Q뛁6�pƥ�Ӹ��K�֎j�YZ�ch��M�W��g���^���5`ʳv�a{�u7�sT�P���w��3٣T�側&ȁt�Q�2��L������{��ˢ1�D�԰�nQ�����[oM���Y���f�P�Cm�Ҵ��*ͣX쥯M0������v�bJ�������^1����4��i��O^�i����-�ˠ~�7$G�_K��0*�Xd�T*�iV�e��l���p��ۚ���яj2���],kz���X)u�[Zi���'�$-:�� N��)�F����D��mZJdv")�m�ge���
��:���4Y��J�zE�~��3�=�k�/��J��޼�"�5c�/�C1M��*���8�md�S4d�J�3@Db���l�xE7�q$:dr�X�Z]ؚ�V.�q[�Y/"��Nm����[�jmn[Wgl�(��W��B[k]��4cWxq3)�/2Շ���1f8�X�q
T��Z%���w&p�K9 n�,�{����_#��
I���F�k��C,f�Ef�4�9:<�ϲ��1٫M��-��v�O*�A�bw�]���ӹ�L8�VM�n�۫pUKR��V.�j�e�9*Y�**'*�h�I�y����׹٨�r�i��t��1=��%��t�N������-<�-L�I%���v	�V���/	m��jE����+ ��*"���΢C�dX�Q�Gr��d�f��.�i	��uy��!fR*f�Z7eT�{���]�H`[��ChF�(]n8��8IWֶjǵh;�v��WW�e1������D��wc32%��ڑa�f��	�k(ɰh�Ղ�hvѤ����H�f� �%:T�z�V�L![*���r�TyY�d���[�,��#][�������)�
����-Q״�u3��&p��}��ɾF��xj���*e�bh����̄����[�S+U��0R�nG�e��`k�Qn72ᗕ��Kīm^C�35���0RSj�ܫ�(`�X�5Ň �SN������E�JF�Sd�`;���sn�ĆaŎ���Fй�Z�=̉+x��
GV��^�i1Yݤ�|]����RF��(k���I-�|K�t�/�����S
�]�5�'i�uc�l��CC
��\Ҵ�wۂ�"�S�f�awC]cOL:�^a�5��\�Qݦ�`\���p)wӤiض�k��PpB��xM��_m-]#}g�i�P���,�[B��aͫPݶ��6A���T�#�	w��깠V���(ݑ7C5�4f��gu^ơJL1��{>(��,�i�6�U�owZRˤ.K%�B��N�6��Ykٺufa n��T���K�5���Ykwj�HJL�IX޶Z5���1c-�akV�SN�� oBsF�f��(�v�xj�Ab�ƦLZ�c�E`V�MvnJ*�S8�Όk)E-I�����-�uJ��ZA���r;q�PU�׀X����G�N�Jԭ{ˠ�fa�ll��a|����36�X�Ok'��e�n���v	Y�Z�Y����=���n+�hiͻ/�"��Y�j�e�4bUm���Rw2I761�{j�����@!��C2�!v� .��Z�*��,���ӌpK�e�+�]�+Gf���%�uh��P�R�
'	����n�Y�Tnl{�ծ�S:Ӵ�3;�̙Z����m��Z�:�V=�X��;LS�n=b�#�w��l� �[�1����Q�R���n�C)���v&P�sE���$논��t��gQ�]=��:Ŝ����.Z��1+"���X���w���������m�:��ZE���4�uj�`��U�f�6���o6�6�(�#@����iT�KR�Y�Mr����X��	[%��nm��8�ۘ�ŅbsQzr��V[	�4��3�MƷF�gC+�7s�Iv�Y�^���GYu�6:��1�DSL�(�F��ܙ�&�')�Y}I�J˴��9*�+��]��deL�5�n����j���J��ip��h���U�u��ٵ���D�c\�$^���Ќ��4��ڹ�K@����qYy4LGd�E�Eb6�E-���hx��X���(����Q��X@qYD�v��ZU�1�TA���`e�к�&��Y:�������f1�֤K��D���@30�%�7Gu�D]����P�[*n%cv�\)�P� p�m��Tr�HU\3�aF��V���YSL�l\5�r�CD1[H�U�5`�'%]'����T�!���-]�E(��ֲ
�7�Yei���р� �4�b�e`P̔�X�t��4�t��"��j�0It"��`v��î���B�Յ�-n�$K�m�۱I���;�X(ʵ�F������YX��l|������l�����j�5���X.E�\���۰�J�aDu��i�w����R���:�2��9R\N��`�#���]�� t���$TMc[�$G���֫)�����z5;^�^�)k���X#��ݺ�e�q\�4Fk�KUݩWN��Ѹ��Z���|�������e�2M�X�f��ڳ�A6��	���Ne,���V 4^*˂:ǆY�����e̠�����,��h�ab��q #�h�穽U��Z��U���ա&?�IE�E�� YfI��oov!c5��[A���T�*�(!cEf4P��ѽ�`�PY	��Jr�]�WB����>����9���k�D�F�l��6�)���o�z0�ܣt�`�����.b��<���Ǭ��
�:6n�P�d3ym�N��j�Q#x���Մ��J4�Q3j��^]�{����Į[F��S2�*+@�����f酹)Ʈ��R7Oq�{�%�b�P�̽ԫ`
�u�����ƥm�N�Z���[r#��]��K�jV�-����[<���
+��]��h4ͥǓq�W��#.P�膞5�1[ҡ����,V��na�-��46䖾�n�M�v]��ىX[7�w,�HY�XjMh'��͉ʕ�2|�މx [ �YJ�X�l�"`7�b�k
��%n�e]���at�V��'����e],^+��@�D��(���f=���Vt�%�����c2\�:���+h<�^C����)��jT��5҈|ފYGX̖LR�6�5j�3	��B�ٕo>ʡ����0bن^�ʕ�"��f�]4�$)�mYh׻�e��j!��g(`�+1%�P-��N�%8�Ѯ���oji��&��[�#bUQ	0,�l9x3s%���t=i��&���+*1vŲ�,�<��Ӵ-"�&�+�&m�h�/�~Хy
���Ņ���P�\Ә�[#�{5��o�f��FV刚��m��v6ء�/X��­�skt5�%y�^����[��h�˥lkt�l!���"���D���o^��"��^� ��;�Q�+
�Y�m!��f:��� kܼ��v�ь�*�Ԋ��oCh�+�kK���Ra�@�;t�{�(��fA�b+F�f�{z7�`�m��e�wA��1��ۭ��C�.��J'�V�8x*�*���7+���][�fm`���QCH�dY�6��۳D�qc{0��
���(��1Pa��l�ŗ��ݲz֓j�P<Y�-�+�gl�@j
�Y����OwY�U�U�� lʹVM�݌���M.R�gD�~Z]��;��_��M	�n8 �X�lg6�hQ�ئ#i���]]E�qZ��Gu���h�����U�N�Uf�PUyn���#n^ek�4���I\�]%5�^�Q1%�n2�d�AFZ$[RYf�����a[QkM�z��}�`��(��w�xj�rā���	�+2�r3VR��&���kq{�;J��-H���q� ӫ7��
�uz�d�!sBSd�Nc:�ԩV�
$��>+1�?^���P�X+����-�h����(݁��-mZ�/(�6"��ǅ�r$�r��X,��̛R�"V)V�j�5oRʻ����p�7]���ASn�ƴ��]<I��ʳ-Mr^�o�4q1�jVm^�&��c�êľ%od��ӻ��V:M7}��-1o��U';A�ç*^e�[�-��J��+s.��)���y���>[q(�vT�o�U��W:�n9�r�^4a�rٲ�hI�����z�6D���܀@�ކ���B���o�m'��!�NG�yN�:� ���Ƭ��7JP`�����JK��.]_%Rhݭ�J��N������~���%pL�h�U�Z���q�}"k$4HR���`VJ�����ɼ1)��6�֚Ô����eZ�]�e�]\�ݦ��r�_\��+/�QhvپU��P5�`�Vop9{�햂<ōk�9�ll�����kb�VT{Sy���VRiwY���S�P�|*MX����EՉ�*�]�����ͨë�v�_G9
���܋S=�u�Ӑ2hw��S���	T��;ܵ��v��7׬WV\ı��թg0H�bVV��/��V�Pȉm.��O4Yz�unU�Fc3e��(��_if1t��Jug����(�q6wZ��/RKS�X�y.�k�P��!v�7U;�h1�&-�aӿ��O��*D	�c���oz��'I7�+t|�ԩ���N4޺��;�t(E��wlo����&i�x��j{�O�R��[�Jť��������J���i[�ѷ_P4n�s��Y�^�:�,Q�k�]�]�E8�Ip�:�O^.rb�&�=�(�!�u�gۅ����\P#W��PQ�_ژ�(�ܗˮ�B�=�4n��M(�:�;x.۽�_
�b#"> Sd�d��[�5���m�g��V����(�0Wq��:ثR�U���v؆�Kܙ�Sw��
��I����7*����UbfJݺ��G@���-��K���Xn-��5�7�Ԧ��Z��۵fq5+(�ל2�ߴp$���@|�!�� P����kr��N���G9?�⒯��1Z@�j�*��9������zk	���9�
	���B���Sw�Im����&���Y�B�[I�LZ��5����ջ������[�����w܊��ӥOV'��T}m��]Yb�b�`�] �c7�N�@Ba���2D��~Z��>��֏�VQ���*e����ƫ�p굘u�B抋��v���T���a"���m����^�$�4�]\x���S�C���n_ov��7ɻ�\$>�C�ū3Ga�faݫ��ѻXU��x������R��]�i�|,���oy^� �)��+�I�E�`�U�m��%�F֥
!t���,��A�ս���"<y��{���2�)���6,8���_qሌ��̣%E&�)�|gi{j���c+��A*�gm�N;�T�#���9��]K�P���B�q"�@+?%v��֜�������{��T�����RqS;|�yX5�;�m�Zfz,�Ǔa>�R�|��V�nq�MQÁ�'w��\��$��b��Q`l���������T�.�v�B���єt(0QUc"�l}w׉U����DV�XpcX�ӺLɂ�m��+)�����4ed]θֺ��U�ɯ\�X�*�z2�p��;��Te�N��أ���=���яr���C��F���9"nA�G{W�o�v�˽�˰�������+�D׵{q�jET��J�%'����U}3�d��ݷ�h��] H'Epg��O+>��}ԝ�;��:�cT�w]-6ص�q�i�_G*W"��[�3iW�67��B���(��l��-�O_V1
����fھ*��3y٭�dyv@���G�YX������;�,��r�?�
ۤ8+ƭ3���WH�4#
��/wy��N`ض���U� ��:�vFub��1���/wy�\�zW�n-���5s��h8� ����صԜV��Bx%�� �T�9���uݷ�����F����;V[���{�>��:�OD|
���j���3]�gm�7WJu��Tji� ������PRT� �F�p^�K�}Z���]n�W�.i�F�uM�:>.�a˫FWKX-&�9�j�M����,{AN0QK�ޘM���R�67ݽ!��A�=���'d�aN��0:3�v#��M�{4hK��d<�������v�+Ĕ@��/l��˼)g�h&A\Y�0�B�U�f��ʤ��P_wow�z|&]Ӧ+���d{�AT�3#��}���2����r�_nuaxWPs5�Q�o����S�D��])i���*K���
�e��ئT)%�p	��o*��n��Zǽ2���f膰�=([�/l2�'_������'���ȋ.�"�㗴�b��/uc���V)e=Sl�{^t5NGA�t��k��v���`Q��Tu��<��S�կq��PY��=�npx-��[#��XhYZ�p��Ʃ�.|mъݝ��齯%�8��3���e���%�RݠYb<M6CUZnuE���|�$�rV��Ѝt/*��5)븮�P)�/J�'�V:�̫�g;tii!�a���En��;[���'~,:WH�H��[H-/j�b���3�;��&kGt������^�mr��%����:�*Zn>89�_�64h���Q�p�K�G���yk� v��R�omf[L�X�Ѧ
1��wݔ�����Dc*�ѿ��C���NY,a�[4����:1J�n�釟;�b�zmYL���ef_Cn�`'FRYSm|�?���\uZ!�)��owt�1^�5;X0�oE;sSXڭ���6wS;����e१�4MshX�JF.m ����]tY�	��k�40��R�ٗ	�8IT�>�cO0����t=��.�rl�Ҧ�b;��uΥ���ek�U5da��˽x�[/u�!�v�"�Z�L����Kػ�j��#���;o+�g7�n&��ߔ�q*9{}���W1Y|M�+�#��4�� �;a
����ڲ�ň�*���b�J�؆T�gVԷwr)l[���Dj��U�~��8Y���i�H�e�d^��؛4�]���g;��]���:Iމrr����mu�z�̨�U��NyPP��naG,��ː�w��
Zxk�u��ǫ^l�w�������u\�J�S�e^@��mu2n�t#z�o֨��^�[K.�����x�<iGh��ۘ���q��Ю�tݹ�sV�����.Q@�'��dhJ�4\}�u{@^ԥe��r��.d)X�7RW+Ht:�xnn\B��h��I�*�Y�;j���8�x�p�z����5�L�v�rx­2g�n��n��,G �qt���q\;Y��x�k���.���vm�L�穔����Vz�urF%k��{(%Q����s���Obπ�;��r*b�N��{z�|�*f�.6�N�N*���}yO��x�MU*���YGS	]k�	R�,0V写�Y!gjiK:��ҞM݃R�r�!3!b���BK�c���wwa�UtQ:��Y +X���K�dJ��swOH�<ȗ|&5�{�%�w���1*K��̥�M�>�
�+�7+�l�ˀ�>of��6�CxV�%}uzܙ2�7�9յ��I����W�0���Y)f3���t2�p���Z"����k<��MqD�)����ؖ��/���-�0\���l�6�m��]�jm��$�op��Uqt�0�'��w�/���<�Y���S����B�d��Q7�w+"�mLx��`}tp�G
�' '���78gUͧD����s5���
{�
�.���E%���Z�r���ںo�(�e�ssx����(\�ި��n����k���8�*+Ts.l��Cr鞥�_�%ܤ�Ns�d\/�f��q����aXN�<��)}�a�:n�v6����'�_"�Z���-r�_^ե���o�!�ֵ�Uq�p�_m�q"�_3�!e���e��"�j)�X�.�����5�X�-��t�D��?�^]�4���d��8R��+8Y��̝&u&bE�Y�4�>�� �s,7f��^�6��5�a��z�Kx�W/MJ�N��.]�Т�\`-h�b!D.�r�̅0Ulu�� P��]4�u��h�`\����U)Z�J�̓\�bgm��+y'��'��>,��pU����ZR	�u6�th�ƧPʾ��N��C�C������F6������R�c��k�{,P�Ң�檎�M�tҖ��V`�D�����ƒ�stt�6n��O-=��*���]e�	G�Z=�H٭'���b����.�z��Y����{>o�r1c�e2o�s9�9�*^֛&)����ʃHV����,]W]�RYa�Tu	[*fԽ��){������r��%ۼ�#��6*ac2���K���	⧭�����d�8����j)}n���`�[�I�6���b���'!t�O�w�]��<P��씳b�����ﰼ\M�3ku9�Z�:��}�-�H70^4F)-��,R�/pK�����t͘�Tk~��.�ڷ[3�ٖ7�(� ���[x#1�DS#��2z�]j�QF=,fʌ���Fj'̔hIO�9ێ���V�&�Q�D����^��*�o	�t��7�d�Q��`CeC�SA���j3pm����Tj�Vu[�yT1�\J(��M���N��{�L���9u.g&����0���ҥ�W�ݵ����N���}4�o�����f��n��}t+���k'&�@��uw�VV���/{������C���˸FT��?�����r��f̫cq�ǻW�m�+���U7�TV�+m�'���I�ك:S���!�I��S�!�z�о�@κʴli�e	s�9�U��Z5�A���GQ��;/8����/KX�M\�����Q��X�QW\���<�\�t��(��Ǵ�9��_7Ժɮo����-�[����p`���{7���Z�/�l+�Tj�g�̒�|��J�sqش8�71��T&d)��p���U��о�5��5���mN�C)��vVH����zV���/p�7��u,���o[���́�#��(R���WN���2�ښ9,`r�V��+���!��W5�V�F�f}��>�m��Y�3�Jp�C�h��bʰ-kf^/�al�s��&�pۭ��O��o�J�P�W)���"y���'j��i pv6�7H�WQ��"؋��0N�:�ю���X"��Z��T܆�թv�\-���L�,]Ewy9��a�J1\Co:����!�n��V�p=�dT�]re]�!��+�R%c���u��o`*�qΡX31ʶi�iD(��|��-S�����wu���;��� ��ŚVp]u��0����5�Fih�LQˮox����^�Lw�U��1\7: U�L=���:���3�.�p�η��o�.f�*��X�3&wv=*�9��L�r�>��c3puX���U�V}�FT�엷���{���Bq��u�)䫕��v���P����C��Kz�L�G�]�.u�|f ��(1h�Q�:إE�<5�y��rۭP��Q�8��u�ۻ9g�<�L���4�����z܋UIiT�}���ҋ�#�hx���W�!�cOm���#��ݪ���"{�Meg-��\���Gu�kS�L"t[���08��I{Z�e�7���^EuF���Q�Wv�!;H�m6S��Pl�n$A�cg
]���zT	+�k�wF��K'1���󩃴���'f��bS��@<!�}oZ�K��(D�J	�O�t?,�CՃ*_;��:欸S�u�ӒB�9��aܣ�Mg���TW:5P4k�C3+���V.�`!�h�yy+v:͇)�\+���2)�G�y��s]�6�k	*�e ��a^5U^�8�Zs��$@�HC���.��fٮ첰��R�2(��%߀$Wd�<
=+r�H`oj��y�s��1]3F�b�Zv�Y\m}�ju��e�̌jYAڧt�n����m�f� ���C0F��ֻ�hݬ�lE�ɶ)��
_B:��@H(e���c.�N5��r8t�%-;�,��:���yG�Ғ���v�n�C*�F�7�\4e�]Օ�vJt�w�����Ȕ�z��ɏ�C�l3Z�-�AO��fp��G�<[D�e2c��Zܧ+Qc+up�5���WG{F@��f�����8�ʾ�%pU��U�AuG*˂ngeٝBX�.�p��^��A�Ѹ� �K\ɜ q<&�CBÂ�j95�n�b�+N߷k����/YF�"�lsm���ʋl5�:����WJ��6��U�t��=m�+� ����ݖ�;�r�E��΂���q��M_s���]��lͅ�b#Pe��wp�7W��)�-��NʆC��G�8��{�G�E�����c6�\�ee��y�{	o�%;:�:�0�|�S�ۛ�q[��A���������V���M�m����赠��A�k���o/sF��ҵ��ݽ�v.�4�w�E���M2�L�t�께1��#��p\�V�,�Z�۾��t�3(��/�&�um��Y��8�Á�Lt}}��;�=�>�rqZ��-o;7K^�-&�`r;��Ŵ�O��	�hP�u�����p_o"����gVoar:ɖ��c�����q�F�R'p8B�Hj�}-��4�dٛ���C6F���5��)��w#�n�mB���s6��cv!�[��Ž�S� �b��+m ���4u�j�J�u�5�ҙ|�G��9�u�ż��@�
Χ�\��b����R�^�u��%K{CN��cV%Ƹ`��DH�Z���|����  ;�SD膽���[,�HA0S�����J�7��)X�W4k����~���Ϸ���		�	���W�}o��ϛ�(����E9Ҵv$4�nʄ+��^Q���:CmT�j�����.f�U��TN��6΢m�T���-�����;{��S�4��Ԫ��z�%�yWf������s��R���a�ʱ)evҼ��I��i[���eg6��ZwE�	��������M����為<S�9�6mm���ۖ�>L�tԸ� m��V&�	V�Y緮E�@x��3��册W>݄nixDt]\�	˳i���*�\G/�t�h�&��t�du}FV�\�Q�Y���hz�<�[Z	=/�#F�K�h�%���5�>1o=�X'c��Dʫ�fRۧ@�L�ͽ}˭��A)u3jHv(��1vï�������CC7���� y���+���nѬ@̲�?4N��^.3`�}YR&��� Y',Y�pg:�f;���H����Dt�&�K^^���=H;��u�{�\������[�ZT��y�4;^��Ed`�4S�2-�6�8�r�;u��D�Gu�B\����cpT�z��bk9(p�Ю�4iR�Z+n��Y��Ou�4iU���5�)ֽ�JZ������WhE^�h�:���΁
��Á)
9[F �::v��7uuGw{4����[\�t�M�w)�b߂i��u71{���Hma���^��b��˕��ۆ��0(Tu"w"�Y��A��p�ήw�k<Ud�!���E����M�N�nS8��m>�����f�oU�Dn��ki��PY҆�d-#6Ȅu2��gr��Bz��4&�Y\�M�u�yr}�v}�,���QO]OP'W>������x�7���7FN��*+�����ҫ�m������ �Ƕ�KJ��ń��hrl��2(�)��q�����M�|�����o+��@evVry�N�,�Ȧ]J�p��p#�g4 �a�9LC��v�ų�٦[�B,�;���+�#�4YY�q�=vU�3�#p���3l�����y�z��3��&�X�2Mu��2�ewoZl�*�b�;'� ġ����(�PWyq0�짺��$,1 �5yJ�B�P��b�*懙E`cq�(L+��8r�w=�g�\xi�(��v�Dڹv�6�(�5���WC��+�IZ�چ�c	�o�ŻG��� Ʀhkdh��+e�����&ç��۷�=}B� �jk���
�ʊG²��	�-۩ի�m*��q
U����� ��\	��ul���u�;6�RA�a��4*���A`pp�Le�A�n)��ɡ[t�RcS�e���<��}æ�5��ڢ��Q���4[�kw�_ZP�V�M���)T�S>����wl���ܗ�7�
�x_u���پ1,V�+2u6/�@ �0�eJSŕ�kT�7���E1,�ϭ�*LVk+>5�i.��w��^��ᶚ"j�U<L�|����(�ιF��
ʜ�X�޺AلN��R�Iw���(���8���n�jk@@ʾd#A�;'g#W��\*���ڨn�fµt��[���R�M�qīm�*"��w�]%�f��]e�seNl���vR±7{!"���K�Q`
J���/ol;�@�Ѽ�Wsª��k�ZfR��Й+��!�4�!u]�
�����m/��YR��v�v�SC�@����ԕ�	D��-k/��M(�45�]����d���u��Ja�YJRz)���橝N��f@���|� ;lUc{a�g2���lV�o�*�G�o�)�պ����7p��"ˮtj$���W�M$	ae�1=�����q��ɚ>�'YC�}��b����ߐT�=�	t��D�i����1�uv�J��;V" �b�f�Cb]f��ԂN��CD$���kJ�zⳕ��R�wm��=73��IG�(��
y$��zَ���}z�8�tho�� �Cn�h�]��>0�Pp�]v��CH����tel	ږ���
3[��8�,�T�KTW1��6؂`�k����w���J�;�\h�xi>|�:Q�&��e�5�(�o����NNm傖$yn��WѼ��ZM�@*�k+[y3o0�`]tٓ���`��(��f��-OHWz]:�j��p���=�u�}g8T�TP��Zų���bԂ��R��n��SZ�[�ro��p*��z��zkKc4ep�*ǩ
7h�/%_���-S6�I������I��na#�Ö)tq�}�5��(��"�Ḽ��n��3pՂ�8qͶ�T����2������E�;Yf�S��eɝ,u��w<1D�si2�5�J�]b�s*k�J�@���v2�51�K{��;u�fJ���Yn�ޡ����A�`c����G�,�8	��9*�kh�麨t�B!Dv�z�!�Z;ʲ�9a_E��^[r�wya��X�(c/{�Ä�bj�Z�>U�Kg�ҽ����h���fI��6� ��86���ٍV=���JH*ၓ��»ioM��́�c��P�F[*���.ܲ�tj����ʔ��v�9qq]�u�6:�i�����JL��N�3(nP�"�r����Yc��+o,���s���ZUZ��t���4��Ư�j�Y.�XCTQ�w�J[U�	\y����9�T�`�(r��R�� �̡Y��6��=�pD��ꔕ΋�o��Tv��:��v� ��ʼ�'����:ڱ"n��+�R���1Y�Ffo �_wu����ۨ�W!��B�����:����!J�a7�5�5L^��}��ΝA��j9����y���&;�'akIb�iΫ���	%�]Εu1�|�DX�W�V�퐳ڧ6��B�ι�+�^��@JlAm���:�6S�i�.��'3)Y� Va�����\���/
�#1�k�X �4���Ofm,"£Oi٥����a.e�Bf�u.�V�k�h�q<{6e�9$k�6J<�;���,�Z�y�
k�H���T
�ݖ0���I���[݃N����A�g4�lj�wZ�|�ia��R�U�]�}6�%�)!�����>�YZ2��Ϫ=��lk�K�C���wB�+i��.Vd4��tF���r���͙��Y�VD6��]�`���l���s��S�u�>Bl�&a�,���3s�B_J� u��aK�]�HY�yG"�Ȏl���ӂ����S�M6}�h���{WI��/H�}�n�t�9g9W�>z�nTܮ�P��t����5�*TY
�B�u۰��kG�$�Z���=����O5�T�����Q�W*4-����戝[Α�d�qwd�.`����7v�l�����H����+~o�Û��\���3��T�y[��+4� aӖյ���N�k/KIiƮ>��`��1L�V�1�w+#.�ec��ҩZ�tT��9�Ґ4yXͣ;���aAn�Ȗ. �Xi����dW��3>��F��KV\<@�(��	%���y�^�e���:+a�ݒ�764����v�����v��7*3]�f�7�S��}���.gg*X�H���1�ŀ�9S�1��2Wn�DΆf^J`4l�Õ�V�Mm<��U	&��Z%��4�E��x/����mX���N����"�x��b<�G]fܺ/�=n�V��aFv|pA�I�n�	�@ܢ٨�R��p1�Z��5bO[ͫ�`�H��ބ�:����/`���qewr��!��3���@k��۝�o4���#&�!v�4� �
�:j��$d�h���A�3�n�
��
�[!�ۃ�v�d��)����x�S��gn��]�:}�z�͗�CW�xi��ú�r��;dm���I�J����i=��bZ{}�)����&�M��Լk��kQ(��2�&�(a1�Dl�;���� �[�R��z��Bf���0P[�e���y٪�q��.�`R`�hn�Q uj��iu�f��Hb��]�t̸m,�gEd�r��NX��T�u�1��b͗��ؖ��ؕu0��b�Y�)�m��{q��F��T�G텭�T\1�yt�ȭ��;��V�I;:����\���ډ���3�U��U����L1#˷/#��H�T�]��,ƭY�s ���Z�jpÃ\-���K�)�v���jj�t�ݕ�G#�q�7�V��q���7�Y!Ie�����;�>[l��kV+�C�����mjü7�j�mL8J�s[Жؤ��F��k�Ak�;R�W��Q(EΒ�Ux�\V9]/�Y������<xT{�z�jf�s"���t���9+# <�rxp��r[�G\�nP}H&w�dI��j�-[b$·��{�2���	p
�Pv\�Y��)���:ܼ!,�A$8ن��U�S ��vه-\J��֣.��Hk3Z��l����qMێ-)�}Z�
t0˾C�k���z��`�ua���v���)+��|zu�y�YM�Bշ�^ͬݽf����	,b\�d5e�����ƻp�L��e���#yF�,!9�#n}ͦ��sqf�΃S��9�����C�1�Rl�SPP�ѵ�om���n��@|/`V�p��JN���o:d���.�I�u�F��Dӈ(�u�'�k@�Nw7Y���}��3i�1�(��I��4��#��RX��V�	��1��� �r3�B�6�nX�e?�k6p��wW�!�*r,R��a��3����� �YYu�%͙
�U֍�/1h����rH�]
����;�t5Qu�Vj�)s�E˻�D'E
z�2�EI׷�c�
�Ĕ:��7B�ݡ��R>W�v1F�Z��XNs�)�vxrʼ�N�jr��WW%�v�+�H��T������t��mȢ��q�u���j�e1Ka�71u`���U�v.���`3�9�#$��sU�r�D�-1����I-[�v*�
w;���d�W��>u(��@�[.�B�wS"
��Ij��u+�m�)�J�,�[S/��e0Q�$�������4'��W���#]��ԛ�cޫ���Ա��f��'m�����
o:��շ*�Ǣ)��gl	Qoz���Fa
��M�x:-]3�'�r��ٛhm"A@�''u����������B��͹�r�W;i�u:��ZY:�\M���n����NN�iC�؀��\��u(�V���E�Ж3Z���#��y��T�}h$!�՝��2���]Ӂvr��d���������i��<̀��P�-���;����+���=,���E�Įge���z��=9ܔªTEW��v�T�;$��uo�����o7���-*4M�ܔr>��_�l�c���&�&TV��������h��z��gQʆƭi'l��ڪ"�i|��4�ەy�qmM�R��8"��A�v.�[���*k:���'��:�n�F�
�Nm��#H��v3�n튷��4����b�Dz���rb��B2�7B�aNn��/�AR�	�\���eh�o���Ƶe��o.��v��$�R��>�ڸ/���*r��t�5�tbD�2F'lu��Z�e����u�� �`7��TөD��s^q��F���LT�8k�4P����V�t����q���n݈*K�}�YZs��9զ�XGe�ۻ�dM]�^�n2������S�a,E�꾷�sJ쫈"�.�hG���c�����w���uz�TΦ��cr�z�����p�H�A:�.w�3{r�s���N�d�
�N�����}#h|�Ӿ2�{�#`�s5a�jPЍ�U�v�h��7�PG7WK:���<\���
��Y�uHn�֗{#�(˥��@Սr��kz��%Y��'˹K1�����������e]Y5�]kxw$��J(�:ܽyA��۳ �����5&։0<qݣY�,k�[c�A�D۝@�=�zS���v)v�լJ�[���t�2���b݁�j�Z �AS	�h�@�@��{YZo�
���t��t�AT�F�#,�&�Q�C �5�[�k
%]����u3J���.�X�)��Ȧ���2�V�NpoK�G`<��ˡʭ�w­�	ֱ [�fr�)��8�:;�p�[;.DG}R*��K9wM���+z9�q4M��-&vFb,�9`�Bg�vԼe�Rek#�]<���å)5�R�o1f�qG���cM$ mZ�0s{mWC+��Ko��Od'YH��8V��j�a9`LQ������u�c-�o���
ܤ	��@�r���ľڸ0�\��Қ
�k9>��e�ρ�0;h�^@t`���I��+��vƙPe�I��r08�۫�e:�>6������3�[���a�ЁBlw:E^VT3R��qQ�O7�l��t�t�|;z�/W�Z�Pe@�%Z�1ahr{��%�x�����U�?A:�n^��'4�Y�\�V�#-�h Ŝ��Tf��\�!�oR���:�S�ڻ8��3��h¯'Y:��k�ͭ�{f.5[�����U���Co�?�x�*5iY�5��,]t���>�.�"I�O#� �jN�2�UЃ_f��P�m;��v��'�>�n��c����ӽ�X�N�l�VpZnJ�p�ȄE�k%R�
J4]s[ש�zw�+���gEF�T˛,C�c��r5�Q���)�\�M��<�pm�=��6�%D��a<E:�0N:9KKE)��\��叜�����#���#�8A,�rcԇeBY�;n�;["���c��75�)hv��.�����p�(��=f�����j%y��T�����{����zD�J���s���V�I���՗���f�;#\�vn��"��+���ӌ��}��T��o)/��]�i�h'�ԭ&�Q�W�^a-��e�����>�.�nc
�Qx�$��k[�m�����
?�������ڪ�ZW-��v��<%j!��f����k �x��f`KM_a����������Dq���7۪���jV�7mm�,���U�<���oNӃ6
��Jܺ��.�x��.:dA�,-�u/���F��U�.v�cS�xCCkT��Xy^�+�r�sM7X���c��Y&�aV�t��N��q�3���W+�l�y����ġm6T��i_q�+vͅo7:�p���+�gL7�KA��&������]f8V[�1)��7�l��6�i�bܑ���J�f:R�:���:M��I�)���R֥�2�q@��@�+�ڶ-��X�ΧR�?����Ҡ�컱�	�ѥW�-��ғUj"Β�6v�~��	֑�s���$����6sMY�T��\���VqD�ɹZ���Ygy�B��V�:T����-���__>{�ReN�P3���?��=�JdP���rS���hL�"��;m\�Y}�ݙ@�yq�[�{Rq˛�K�\��ѝ�ǽ�6<�o:bd��d�]���z�i��-�l��.�.3�Z�o+�N{t�m���D"y|��+&sXU�MJ�R��AǫZY����<W�O���� �l�.�]0�K1�i3�喀��un3���6΃xB{1Z�ӏs�����Uq�>�k/\�,l�٦̬�f7@�#م����"�v�N�J˞��?��?bV5�L+Qűm��̋���˖fPp�b��X-�J[nfLiQb��EV�E-Z�k%+�dq����(���mb1X�e*aZ���V�-���[*֪���(�m��\j�"�e�Q�֢����ĩR�YkV[(նZ�[,�Z[iVڢUk-�h�&"��1j��Ҵc-��Q��,+\l�-+[QTQ��EV��[F�J���+Ib"!VѪ��[B֨��DVZPLh
�h��Q�m-h��("[P�klm�UR�Ҋ6�R��e`��h*�Z��J
V1�j%�T��V
�����E)e�ЫYUF�2Q[B���&8�c`��իT���b�m�Ƶ��m�lm��Z�kKR��Q���Y(�,������h�er[��,P֍�>y��yS�v઺sE���l��I�x"��28Qݟq�ݞ���wm����R�*���Ǳs��¿Ζ�A��rp�%tL?�R�{��5���Z\2�y�,��3�Š�]�}2���5��&;�`����*��u�E)a��
��c���}��ی+;�M^�Lz�Xy{�ȏ�x u��V��v*��=�o�ӻ�B�7yGα�'����J�"��/��+2��Q+�$60D]�[�W4=����s�S�~��t(X�^#="e�Ҏ~��]�����ȷ�ΕaJ�����]s��t��Kj�[T%q��NW<���%*z��B�/�����$𛜷���{��g5����I1����.K3�V_V�����sq��z���w�����#ް��mfF����<��F����E��r�HW��z����Y��/	��&,�,'�PcR���{�{j�k���d���(�U���~�P�i���𑩘=������)�{U����6}F�-Log�3"�j�.B=X��>��B������EV����}^OM�����^5>�/:�h#l��[�ӏ3G��w]�s��������!�º�#M�����i�Y�}��L�j�m�c�lLTR�VQ�����K�9g��?�4�Y���{�[g�5�QS��t�o�֝����GX�<BK��j2ܩ����׼�Wf�h�(Ȱꎅ��3��*��P��dk���u����j��Nx��}�{���׽ء�~�3�\}�I�DP-���t{�$�z4�kײX�(�y�q(��,Ғ��74p��ͮ�ϞiT��k����̖<���ß]"ƐdJ��3u{|�[�q�)�^xu���n�y�7��\�����*_�#B��2�=l=��V+���D//S.V�T���]S�����v�����3�<�B�Ӻ+�N0����}�sk���[и����e���]�Ƀ*lE�ϣ���^f��S70�5���/���^]��fP%��~,�f�	A (�u�
���wO�{E�^��H�Q
�K�i��|n�ymvP�x��絙ñ�C�W]h��Ą�,����U�6+�,mf��b��Q':z�+��׻��OZB�����|݆v��@hS���̮�+�aU�@�Į7'��)=��}���x�(�L�94�\�E8��N_��z���)�Ϗ�j��<�^cO|����@Τ1�C�(�f���',oM�n��d�V��n����\N�^�J�/K�=H���W��e@
o�%d�-��ï���rc2v���*�ΧN��C�������k8ʂ7}��[�3Ρ���n�!���fa[nܜNM�����{�~�{�~<z�!�|�`�{�����X~L��r:~�_q'�^R�cN����E��L�}qS�+��Z��՛������	Oc�==u�^���,Z=�����E�_b�9}~��K�J#�U%*�U+Z��3���_�jbcJa��3�zA�b��}�m��x�����z�°��	���3�_]����uv�A}޲�9M|�I�k8ݾ�y����o=��|��	�p�&���Y�I`|g�-������ ���Z�7m��H�wY�~Ӱ]KN��/�ʼ)':-쯃��������kB��_�ԝ=�W�����$gυ��ɶDX�y��3�s2�]NO�5nS���nk7��D����v��}f�L�q1���}/T��G'嬡�~�<3�.�*e��䚯�|�	���x?H�}�hT+h]�̫����r,e4���z�ײ�p�T�?yOE<pI��$��Q�=�3�n�O��/��� X��Ʈ�*�}�Sg�c�ek�KY�����шڡ�s�"��҃���V�Q�¶)zb�	�����ۭW�����']Cs���ww/��+�b�ބ��Hwa//$�X�m�}�_E�ݨrV�wr�J%�h�Bmc+q;)��e�����]�c�M.� U�oҳfZ�n[1�dw��ub~���{���S�pD	],�U��U
co}p~|�9�<',ҙ�pTX�I�<�X��erɕޠҭ�}X��e6�e�q��;=��72_$�9X�9G����=�8�;�$����:NX�	�)�T�Ȓ�P�r��*��9.ɢK��͇Ғ�Y�����tL9�tD�`�����[ *�`y|��H�j���� ��.RNDP�K�+펯%��N����<W��^�~�C��<^����I�9�����ٛ�z�ۯ	�X��m+�%%��-�tJ�gV>�����U�P7^^�������n�F[i"g�51ݶƎ
��W�gL'����4���T�ْ���
��e{��;8���خc�-]�MP~�{}m�]�d�f�̇��~��d�cj�m�{8���<*y8|���+�0�W��w-S�)��ԅ麗βR���Z)q"��޲��Eޜ-�-)ܡs�H�z.Bsꚠ�E�ʞf��b0}�"�ϯ�R����VU�&�ZG�����5�7T�OM����. 
g~���9R�I%�� \E�:�]���O'�ڟ1���]�2�`�D\F�n���1F���Ԍ+L��Zh�;Q������ܼ�IVQ�e�V�����r�����RSܛ�2��q�ۣ~��`��ʞ̕n�^2�z�;��*�;��}O���ޒx]�/���)����e�4J���y���[T��o�	joK�Ǐ���&'��:N;<��x=��b�V�ut5͡Ng��k�C���w�[��r���Vɝ��9S��ڑ(���)���s�~\�L�;E��;�a��3��b���w�dZ���)��
5�p�ӯ�*��uiW����=Z���3q�q���j\�̩t�݄��z�nў�#��<�q[�P���K)^���n���_I����S��J���7�Tͬ�� ����E��z�]�U�ʡ��Lg�O}ݳ3�u�!_S��Yܴ�}c�����X���rn{__yW�,�{!��t5M��43�0�g�S��\�>I��	SvR���et����vk��Dfy}X���w�Q�e�i�}I��;�*�ņ;�	d��GZ�an�
�\��'��!hZ�jec>��-���֐����޺lw�k��zɝ��xc��B+�!����u���1��\�����(�i7øՎ�8�^N����Z�Z������˷ZR'F&k�!�Jz��E�{]���Z�{~<B���BTB��!Җ~������#�Q�ev�WU�E�/eS���$�����O��-�c�<@��z��Ҽ�{�t�z�y�Ulx�\���U��Y�??I;|���{!U~�tk�;�_T����p\x.*�늏p�R�ڄ���§�:s2{b��=w� �x�\�>ͽ~���T<#G��;[���z$��3ͺOҝ�:������3��}*p����(m�C���CcD�Ur�}������,�&�����0�N�y'<ʜ*��۱�C���S�)��n�|�W�X�}x��k�xfa���'ӣ_d痟T�x�Ɣ�3�t�T�¹x�NW�W�>2.���F�_���{��7:��oTȵE׿<���͹���֭}�$y��+P�(슍=���~c�G5���f-�r.�����^�8e=�Z��+��gR1�N�U�b*Y�[����e=���Řo�h�bL];sQƀ�"Z�chO��BF�R�z�Gn.�cT}��R��M�x)k�+2��d�m`�����ݜ���6M��&%������[����L���K�r���I�R���̝j����Dx��>bH�_�()���K��OV�!N��N�~�s�^��λ�����ϙ�Ѻ�r&m#K^��ލHISn��K�̔���k_���_MU�τ���
H�4�08��sžI�k�N-�߮��^S��=�ڧ�Y^W9�����l�n<��9�7�~Z��F��3�%�\��}���oхNy��~+ir�ߜZ�q�G���]��Ǻ9��J��X��٪OR�R��r.q{�����.��Þ��>�݇S��p/U<�����ȑ�����W{d��qS��*9Jz��m<�s�NX�ڷ:t�KAl��/�:�B:_w����[&��\�ڞN�>����]z��x�~ؼ�,L�����;���Im��T�[97}����;���.9ш�z�j���ClxH���z`���h��s����J(G�έsB�7O�ʔ��K����'��q�ʌ�,)�����T��T���$��{VYO�m��j�U#uv���%)l;h��6��yV�ɚ�r4��٭�'���r�U�^m�,)�R�M�l���W=��2;�χs�W��.U\�U-��I��D��s�eN��۱�UΟ���v�7�K��t�3���<�=U�>v�!S:d�N;��Mbԡ�"��%>�����*���F��.�����ǝ�N�*s�^L�{'���av�������E�}S��S�]4(����>F�����S�힩s�{�G�\=v�}��֛�ykr�uL�}�2�m�R���Y>�+J�ҩ�x^�G;=�n��λ'��<���-�9W�rz*�`:�;�������X����<�̤�t�tҭ��r:����?R�r�켮�*4�I�~����uޟ�2�K��d�wl��y��q�r��J�}�p�����v���^��0f���5s<�;��L~[�2��о�(]?F5�1����s��}�ߙ��b}Ҷ��ʻlÞH�����Է���d9�&�4��C���v�����B�����N�����z������i��w6����Ǽ�����u�R�@r4i��^'T�sx�z�ؑ�Y�J�,��ٺ��]��ᚵ6iIz�\�Y�f`����R"�J�<�LY2���'�M�&�z���2T�oW�k�T��C{����D2̱hU�����D��{�q�������rq2����}/�6NX�yl�I�=���K��_S��Uz�w��9�������ƚ��{=Q̉>w�(�I��:]��T��s�3'��N�ok�ٹ��^��f�>/ݣ���'Z�]}���={*h�͝L�oLj6}���(�n�=:��X�N�����g��<���3��߂�{-{�QnȒOe�mO��D5�[����s�.���!�b�d��������3��{�5�NyyU2LQu�v+xA��#]*����)n�L��ɽ�|�t�y���K�yRח73�S"Փ"����GX�t��zp�G����w1�r�]?A�^��ӳ�v����9Թ��eM`��k�c�ז����1�M����K?;���Ó4,�k��٘w�.f��k��96��i��QOb;��y��K|W��}�z�-�����Me`�w˵5뻕3f��G���h�(Z��:�ktr��B� $�Ӊ:Y�L�)�2��ᑛ�|������E�����iV�T�	n�9Oգ���@�4��a�����mʙ~[�K��������yt-�w|߮��xq�_�Y¦�P\�:�\޼��l�૝zڶ��cU�2�M��w���>�����!���~�W�0�9_��W��V���+��Xt�__s�~t}-�|�61m+q��w����͉�]���Ԯ�^���n{����Tx�/}n�b�z�z��2�n�SR�j����Y{���ױ��I7|��<��]��据��L��2��+tCz�}y+j���:�2׹��zI�u"�Xkz쮑u̔���(+� �����p�N��%w�c�눹�>���t��y�6'췯sү:��5G���U���z$���<�[��ܔf�)d�۸���^?��B��3�u���}W,v}�k�A��֪��uG�@����-���t�=�Eu9im��L�d������8zI�(�l4[2�P"��߹�U�9�}��ßj�W�T��G�v�������O��Zty�C�E��E���	�}�*@B��>�6�F���̚c��6s^َ<��L7R����#{\�
�TLκ(�ij�Ҷdg��%��du�i}Ub�N%�|�����W���t��.&����a�4��ڥ�={|��Eu)j���l0e��q{>��1u��F;Z9ӱkh��]Hy�n�CVVwe�c*����h�v_c�0�Ѣ�J�:݈�s�uw��b$�\6eYC��uJ���0�fԎp-'����H�w���ޕ�b�Yz��빐-�*9�N�LVv�h���4�s�SToR���aS�n���I�̂��l�3P��%��[v�j��cK6�'�n0��I	uѫ3`����]u���T���kd��
]���;���6h^�x��P��f���gϞ�Ct&Z��!�ɁϖJ�ˢJ2���B���@�h	p����۱/��䍦�5�����W�nl45K����c��L�V�&�#�S�ľ4�����s����(���Ɋ[����A|���o��F*ɂ�f4j�����+Ʌ1G��BL�m,�wV�R´-�YI�om�jW.�eэs�2XU�]�4�/L��1������{�
���w&��#�N�GIf�Q�X���7�ѥ�*�+
��Y�B�d� @ϝ�]VФVfnum�]v��u��;��v*��2�b8M%������8� l���kV=��Ad=j�dK��W�ܾ������@��� j�sN5,볳Q]:�:��H����5g+��p�n�M�{G;�x�2�+)p��:��:-�+05dr3V+
W-�������uj�ɉUՆ���Y*�d�R�m5d���0&DΜ��WDĐ���pJ�J��환I�\\��^�m�oe�Y��]�iǍX�
,�!и��"m�]��Ğ���(�]��a��ʽ��e=����6:��(jD��ӊ@�b���S�.���d���癒a��Wƥ	W���8�Q�8vk�Ff��O��oKa����F�l��{y�H��>��ډ��m��u;Zn�����m����2���z�lW����כ
���K�4��e�vk�a�4���'��w�p�1�9�+v'�)Ru���^e)k%O�C;;%��OMMq\�߳:�/x������9��Aí]]=֭�/����̒����6WP�Q=�)Ү����%XǍ���zg$��2Ԣ�n3�g&QZ�6i}ʹws����t2�B��ao@b����ƶڼ�Ў��d��sS�P��F��s�`BXm�֍��p��ݏ,�{�����γdfd���XA��74���pt4�64 ۘ_І�4���ihڍ��Z�R�,�b���*�q��)h�-J�pD1D(���(��ŨVѦ%ƊUE�ĕ25���2�U���V�,��3+�a[K�PĊkADbZ��Z��Z�Yl3("cU���*�Z��-D�,Qm--��RڭlTb%DYXV���V5��mU��Ҭ��5[�G�E�iKj�)Z�P�5����Em)F,���kj-eE��(�EĪ�X��m���
0�U�*�%�ʋ+U�Jմ�ڢ[*)iE"ZUZ���-eah�r�WnZTp[F"�کc�%�Ҭ���eE��­
R��[l�c\V����QY�\j��ڕ�Akl��*����)m���q(ն.`3���K�e5RjU�hV4;�VB
��M��A�vL:p�BW�*�7ݸ����{��eaS�)�3y�NH$}ǘw�h�~��^���s����m��j�ϔ��<��S�0��p���QnWS��������U��'�64��_L劽���xs�;j�Vg��2��r]���Jb��|��˞ym9������^,ތ�v�5�uپ��
�e����܁�~c�Ts^T���bվ:��{�T̹6���^7}Q��������Z�{u��S��1+qj��B_d��Z�.�P뛍������t ���g��Ʋ;��c)�r����-���=��:앯��nB���|�?WJ�SV�`ƫje��7�����d�\�y��5�v|_>F5��o�yFz�)�Jߧ�V�E|w=����oE@F =�5�n��Qy)��N�����(m?F�z3�۪['fab��=5����3����琛�^�'�yJ�܋�^��������KQmH��¬�t�<�/V�&��A֊ڳ@*�N����z�2�T[�3WqKYȿD�w��}Wy9r�S������{Hpɋ��Yۂ�]�S�J��4aۋ}ø�<lж���y�)YQ���kU=�I5�xգs�ݓlZ}�J��d蓋f���e~���7�߂��	�j;��n�w�J:�}G��6��hS`k[�d���H٭���W�~�ټt�m�@5���
.�*K\��r7���'sj��8G�NI��^~_%�h��>���v	��y����z7�}��*-��:T�%���~�T��M6�	�����g�L�mgy�z誮\���#�S��9����!�F^λ�͓�g��&G�Vk�}���/=@g�󱐩�|�z�WKo�9g}{���������+xJ��#\����S��������Nէ�{��Y��^�/����Wg<X�yN�j���{�Ne.w6��z���o]��ן��gw��nq�s�"�2%U2����=:���:��{��
��ߗ��-/5Q�E�g��u�ӕ~���S*]S@�;/rm:~ζ�Q��Z�i����Ch�����ˤ6X�ٰ���aڂF��ltB_X/���K+��U��^o[�O�8�<�G��$�d�+Z7�D���%��T�y�Z�=W{�WiL��C�q;1w:jܡ���wN�|:1/�#�.�n��Yl�mƎ{�c��S�Jkv���Z�?R����շG����i�}9/9и��Tw�'��?eww���fgt��/�qҧ)�L�B���H���z˞��k˷���'fzc��)�>��BB/u<�����V�t��]�V'�=4eW:ۯ/E�1��%E�U�3��'��s�Ý�*�jN��S+ɺ-z^��3����/k�3�!��I���3�ݑ�|�zsI�*�VI%���Y��1�O{�?n������uC�Ov_�N� ~lΣBuw�@��qU;��G�NH�������vǐ�^��=��ގ�>���.�:5Z��}���?8��2���4g�)��/%��;U;|�'/%=��B�]����\���l'�OM���^Φ#5�GA�uf+?����G��~V�}�=M�clx:��y�{���T��mȖ²U��H#qoج�%7~R���Ū�w��y!�
8�֙��B��w\�Ke{ez��f�C}w���J �u�B�M��C�Y�&�:L
d�I@2#��=ݬ�ב�ӝ����ӓ����b��Ʊ�S���f|�ʀ�9�iA-��r��K[ILS��ތ�gNO�z��Z3.�&��}��c�7sҌ�sGE��ǺWwy��Y9���$�^�݊?o,�����Q�v�[x�μe&�)�7*���y}�&w��E�*dK�^�v�Y�'l�r���+wmL��w��l|�r�u��R)��ͬRw�{<����l��1�z�U��-��u��u����Ku����3��=Z&s�0���_]��j:R�o�bʃ���[����Y8�o�:I�'jox��O
�����D}_���oz�����g>���Ox�bs�~d��9�P�'�Xy��'̟�y��I�oܒ��Nxk$Y;���d�>��݇��d=��`�+�����d��ѿv�|�|M�|��v�|¡�s��J��}�Y8�����'i�f���d���$�'�~���sv��N�aԟu��?f����޴|��(}T/�7�}�����x��I�V����.��$���7�PXO��sXu��P���Rm'̨k��2i��׹���}�C�����<]���_�1�;�I���n_��6�i8Ξ��&П���L�P=��I�:����XI�C��'S�I�9�u��P�=�u���'�X�`��y��*hi����<���Z[��1���h�zl뽶�=C�6n4����[��}�q&�	!飧k����xP{��㹳B��Ƹ]E|.��9�����b	$9�p^oL�9�]��{&�4� ��[7��=��s�G�bR�2�v��.�n����r������,���O̳���������̜Ad�d�C��J�C��'u9�'S�I�=5�:��O���&5���}|o6��	Oԯ����Oܲm�z�<�+'�Ʃ6ԟ�q�	�c'S�,�	�?yC�,�&�p:��O&��T�I�T�N$���`��)z3������{�|�����u�N�0���a>t���rM��|�2J�L��C�VN��L�'�N'�Ld�C���C�,&��o�2u+/��#�{�~��~����{���OYSZ��L7�q�I��̝a���d�wnI>t��|�8�m<�2J�Iš�+'�XC��O��2M!ļ寿~����߹�k_}Ͽ{��
�2O^�߰8�Ĭ9��8��P���B�u��;��$�'��� m�OY=�܄�6���
�4��~�*M$?͡Y8��޽���0��t{߼�����Z�`x��>N�d�$�~<��~d�w�8���CG3�N2w��@�I��s4��O̞�� �Ğ����p���'�}�V�?~��y���w��}߯��{����IPP���hVM ��hIԝeM��~a�d�f���:�����	�7�u��F��x���>���<d���������ۙ�~s���wo���d�o��qӞa*
&�VN�d�2���I�y���&�^�u�'��d8»d�{�:�4�埙=a7�:��?s����?����uw��z��O�;��8�6Ş��u2xw��q~�T�'��VM�d���@�&�S����Oƾ�i�:��=9��]��Ý����eA�#��nn�ԇ��`���`�������8�H�̟ �Ý���N�Ld�I��rJ�$�^0��}@�e���d��y��q	������~3~/%���Ig�ݴ���}�wzi�mxK]6�p���i�3���Yӡxwn�S=��)̜��+�,�ia�*�FR��as6�e���I}�͎����.�}\n��6ҕi�>���"�h��K�Z��t��f�����:�.˵�2v�p���=i�&�6��ֹ�Ğ0�ZβJ����a�a1<��Oq!��(q��o���Ԝ��'䓉7��d�~4k�>����OH����������>������,:ɶC�������I�����'P�oy�IR��}�:��+��2u'RNw'�8ɤ�=�)4�n_�}_~}kR��L�����~�����\I>{9dXz铩�d��'��2q���|�d�'}<�@��2q��7��!�k�u�T�s�:�Ĭ�;C�d�+������x�s��o�o�����@�'g=�����}�I_Ri�iXO�~g�C�&����q��7�O:��?jɴ?2u��~$���-~�����:�&��P��_+���$�\��+!�]���4�'���4ɶO~��'�>�����8�e��Ԟ3ɖq�|�?ya�a?��~I��~��W��߅Pa�O�=^��t�����Bi&��a�x�z����Y9�	���u���t�����O���VOP?Oi6�O�8���C�~d�Vq�|�?0�
I��z|o��|��}���y���I���d*M�m+<���N����u�0�a�N�q�����P:�N�>�}�q�|��J���t4���N3̲3�'<����8���s3�^�ӛ���I����:��g|ʇ6��῰��Y8��s�!P:�����'Xzs0�'�m���ܒ|�'��$�	�_���N�����C�u����_��'�t/�O�R!��J�$�gP�~d�|7�!�N%`y9�%a�N�!��d�d��9��������i�'���4䓮�g�߭������}�{��7�~�+$�w��J��C���T�Aa���d�y2��m'��6��&�7�!�N}d=9�2q���}��Bg�gΙ8��W���[�G�Ryv󛙟���fw�C�p����m�9F��H���h@w�fޢ6JM���i�k-H.�D���)��Atd;=]뛻vnCu�Ub�i�
!�r�R�ŝG���X�!O6G�0��W�;q]����IXC���8ԙzWj�Y������sz��>���??�6����Bu�2xs܅d�O�?d�	���'R~d�N2u<��6����g����6���-P8��l<�r���w}����k�5��z�ē��i�'���s�'S��$��}�M��O{�d�C��2J���Vm
�Ԭ���m�6�L,':��{�ݲN38w�9�|�.�{�Ͻ��<��u��M�I��8�=v�{�>a6�fd�=��I��i<}��:���w�$��y�T�&�$��J����&��9�2��>��_��}�w����I?2b~Ն����� �d�7��d�z�����'Y'�8������ �Ý��CL���u'�<�VV\���o���~�}׿k}�JɽX�OY6���x~��`k���:��5���'�5�䒲��s'Xu�s��̜AHy��8��y��}@W�>�i	�k4E�POǷ��IOVgOY'�;�p�����Y"����)8���3��:��C���2z��>7����'�=��u$��}�:ŒT�|ì�AHn�׺��}��k�7�כ�?2m*�Xz�Ӟa����߹%��9ᬑd��'S��d��'�~d�!����:��$��d��N���ΰ��QX���Q�{��yW������'��x��T��a�N�By�d�'4�����d����$�'��$��N3hO�?'�Xq�z�=C�N0����x����A_%4����|���ovN��|�}��m'�.j�x��t�0�	�<��N��+!���>I�Mj����d�'���2N�|��i����6���y�q�|��u�������ϖo����OBQ��+0���É�'Y=���6��/���6��<��:�2OY����8��x{�:��M:I���>@�>��$��0?R|�O̜MSo����s.�޳�m-�c�=&��\[�X4�4c�iu�y-��.�~=��̎
&`���ʛ(^�O'7r�����<����G����mH6�c����JY�n��N,G!�'���3��a[���wi��穾@.y��.k�ԃx	�����-���T��_�R���_W�}����?w����ɶOS�2�RM���,8Œf�p6��O��i2u*{�Y	�a̧S�	����N}a9�u���~IÖ}���W��-ʝ
��s��,b��������q
�z���Vm��;�PRL׎:�!�7�B��'���!8ì/)�l��7'3���}_~l������l6�w��N����I6����$�$���0�&����+'���C��l?$�+Y&�����Aa6�߹$�+�k!Ru��P�}B����X�,r�y��G<�F9fl����I�;�^�i'ujI��M��!Y&����J�I��|���,?ZCHu'�ˌ&�q<��:��&������R�u]��D��z�w�c~O�UFN2|��n�T��;�v��O̞�� ӶORzs�XN&�<��	RM3�?d��	��Ь�Aa��C��O�}/����������a����0ɿD֯�Щ�	�t��C����{������~C��Y6�y�i�O?2w��:βz�����&��O{��'�s�IPP�Ƙ�#�
#����q��n�����UT�d�;0�OXu���Z�8�N}��'ud=��8�=v��~��O�O5�:�'�6���'S�M0�;���4w��qw��k��w��[��{�����PP�����>eI���u����'4�{C�d�NCd�铨y���I׌=��<a�I�^����@���:�3�uW`U���Y�������v�b$"���C�:s���&�Y*T�OT�ed�8��'_���M}g��:��9� �d�Z���Xxw�z��'u�������oY玻������'�R�r
d����d����u���$�XN��vE�~����&�>>�:��C�����OY8��� �?_���{�R�r�^��u���knT�Ǒ�L���+i�-��X{�:�d��[w��QTtѭ�u����p�:O���gA+p��bWn��5�[X�"gӽW�����$i�ۼ�:�����u1c0�̷P��|5^�s,n�"ʹ��d����UW�U4ï�Ϲ�}����IR����$�	���0�,';�P�'�Xo����O���'o�%|d��Y"��l
�'��^g����}�z�|�BS���7zU1�M��N��@�x��7����u�T�ϰ�'Xs�$�M2���&�?y��'Y<��$����o!=~d�y���=8p��^k�׺{�~�{�6�|�Μ�����O���l:�������/9�$���7�PXO���N%Bl��>I��eC��=d��Z�4+�
�����"�~Mݢ���埜�������6����l�'�a���=C�N�>߸i�2q����Hu��.j�x�P�,�~d����ì�J���?]U~��HWߨ!��d����Mn�ϵ�@�M2t﹤���ϩ>jO̚J�i�d��L�����P�N�?oܨ~d�'��$�d�Vz��8��y��:�2OX������{>���ޝ��y�������d�&�I��rN�O��$��0?MRm�?$�<�>O̝J�0�aS�(q�kƇY:�ɿ���
����ҿ�]�n�?ޘ����=I���5�$�Nfd��	���	�L�ɴ���<�+2��Y:ÈVC��N'�Ld�C�������b�O����䗿~i���w�|�Vg��T�I�T��B�u��s�I:��fN���N2}ݹ$��'�|�8�m<3̒��C��>ed�����:���~���>_<߽�}u�y�>��m�z������I�����'�<�>@�'uC��
���;��$�'���oz��v�'�O;�B�M'�9�$�|���R�Uc1��w�h�Ϝ�VM ��<C�N��$�N��,6��&�7���~d=f̜d��>��@�I��f��z����{�u�ORx�{��>��qt?P���1}����X;��HU�8���h�f��B)ٛ�+�M��m��&������5[å��օj��' \B�氮Y�;�J�q�[V��:=7h?��{QCRf��D(�Ԩ�4[���n]=k��Cg-�@dM6�Io�����U}e�>p޽���a?0���	PP��B�u����I�|aI6����$�>7��:���`|�z�f�d�&�M��A��>�U
�C�!z�׌��:|��M3�&�x��I����{��N��s�%ABd��J�Ԭ��P6��6�	�M&���RN3Aϲa]�u�����}�]T���<�9�翙o��I���N0��M2~I�y�'Y�&س��0'P�'|��N!��2J���S�+&ҲT�@�&�S���q�I�_d4�_~}R�o��1�	�n����w�?o������0�	Y����$��c'|���r
�>Ag;d:�̚;��'Ry9�IR��x²m� �X>��������+������a=�O3��=Bt��<v��'P����OxkY�IR��9�:ì&'�;�ĜAHy��8��<�p��䟹�O�'yP��>��[�I��c�~�:1��=�!)�Y6����'�'�S��u�����ܞ�2zÉ>����'P��Y%J�s��J��2u'R�O�q�M��O�_U�|�����_�Ix_A��1�y����'{�I_RM>�,=~d�y�d��'��x��C�i�u�Ĝa���~d���|�Xy�a�IS�ϲ�_�z�_�P����y��O�������a�'����|�ٯu�I�O��+�M2u=�XO_�x�2�M3���8�}�p�x�ԝI�VM����<������_�6�N�s��~o�xO��y�7�{��|�>C���8������4�'y`|ɦM��~����ԟ5��'�e��Ԟ3ɖq�|�?ya�a?�
�
�*�o�~c6gn��[���9'�m������8����Y�I����Y9�	��ì�dۤ�y܁�	��}�+'���Y1�����N���x}��(���ݾ��|嫣H�^,�kj&�v����å�u׷0�$�&���0�\I�.*s�T��iY�.��F���cz�̫"���q���5j�7{�I�:��q����^�g|�h����:��AJ"�X�]֫���l\ԹR�DJvmūAj��{u����Ҙ]Z��wd���u	��j)�()6A��}A��X���X�_�F�'P|����X��.���)�1�q�ȱM��f@���v�xW�M[&>�gfKCF�x�b�*ײ^�LӺ�k+'W|�4L���H��q�Я-p��9pރ�KڗszE|��V�hT�p�nm�|�m��,�Y��+(�8+Ai/.ՠ��v�6c\�WT\��k��X��FBV,�؊�O3N�.��a��1!v��v����K����w��eZ�"3�m��R�c�om,���it�/�W����I[eI��.wd��>���=�gY틦c�K�����W�$v��(��Z��x�ȁL�%'c��=0���t)�uh��)�� "�+�:���	�&3|wTY0�JG�(���a�8������Q��+:n�r��:P�y��F�ي�<��͆����؛��;Z&�V��S̩�D(��l�ݣZ�K��{i�G1��8�
��[p�u�[j���ƱjHǩc�6�z0��Ns:v��Lg������ |󦕖��.;,���=1v	i'Cze/�VU�;�M��j���fҡ��l�N��4��ƅ��ކ�YnL2����ܩ[;��7A;-.�!�]�:T�C��tX�2�뭚���Ru����ڂ�C"��^|K�lm^%w�2ք8�	gj|͸�U�R��Ҹo�5˹��j5+������c���ս&*������7�+Gv�f�(�R�V' �Zwe�䚱j����нR���T����i]Ѩ�o���@9A.
�=��l�ʮ�[i��M���,T6�#�ך(}dcOd�h��Q���!�Q��\	�p��j}Z��V�,^�GOIyv�e�4.�3v��:��3�%۵���ɸr�w=���vV�[�.�ۼM�bͣb��t8�4�"�K7�Nw\b��f9X��}����J݁�Gq�vlKo6B�h:����7�8Л�nhXxiew[V-�u��z�������x�Wm\�rnܣw�E	����ᅖ��|t��X	�+.�XB�|^�������<9��l	;R�AJ�¯M�<pT<y�F��ݎ��(����r�/�8��V3m^):�������z��Xk����[��D��Jj��a7O���[��-�)����Y���j�"�G��N�!�[N��m[Z�E����}6�|jT��^vL|D:�o8�zJs[�	��'\=ٗ4�d�uq��uuJ��w��v�5GQY)����g*�c�&7�`Um<�����������m64�홃J�he�R�Z
���VV�R��m��5PR-am�A����mkP*TX�m���[D��V�������l�-���akE �lRVZ�R�D��V�VT
�V��V���j4+"���D+UP��Q�R��m��D�jVQ�eB��%*����F�J�ՠ�h�R�mQ�[kQ-���V�jTVՊ����(��KJ2Ѣ�T*%RƖTPZ�ZũQ�+m�YV
-j4j�ch6�YY)YciZ�e[`҅Tm�Q+kDcj��F�ұ�T�%��KmJ�j%��0�m������#l+D[J��kTV�Y*�ڃj ���)T�+F�QZ���%-���-��Q���R��ҕR
+
�Z"ȡcQT*�iJ�Ҫ����KYb�B���ֈ�id�m�D���-eF�j��*(_�|����n:�@�:`XrkV����W9�;�(�!�f�����9���f���E���D9�`�л�ٷ���B7���k|��y����
��~ըm&�P7�I�N%g��'u9����=�xu���'��Πu��2}>�8�>|�$��`m%dĜfo_�Û��~����{��sI���ԇ�}��~�.2O��1�����*d�V��	Xq��Y�>��~�'wd�a��ì�~I�O��$�:I�<�8�q�}���������kw���߻��Vd:���i'Yᔆ���ԩRM!�}?P�~d�w�d�V>��:���9����C�s'ua1��}�4��Ma,����8myz~肗��w.�����2M�㟲J�L��i�'PX~����'Ș0�I��~��~I6�7�!�N}d=�`|��N�!�w�	���_��fw��l�4�o�>���S߿yd��_��Z��ʫs�Ч5�i���}�^�v-v��ӽ�ͽ�R�/�痕2LYS9'�݊U� �υ8��oLE��/n�!�w{�y�Z�c1n|�\��)�݀��82�e�{�9����7.U�~��W�}�O���Kz��'�L������R�w%�j�wz7o���5`r^�;��{�4�vSr<�Kt��~�5M�1,��oHC^����`j!��R�)%ο�s�n����X0ZC�\��{;p���ܓ�+Q�op.8/�k���U�:�m�K�V���m�ԩ��C�)�[{�e^��j4�b�k�k*�`�3�<�׽g+mL�������ǰ���R�!e�ö'T���b9�s�0I�25]W�1���6��k�kk<V�T:$��������#�$.��������:��q}�1���B׽�;��=G}�>�O�{�h-�I�!;���z0��=+���� ����E�X�U5�B�n�L��ٯ{��}�R��w��t>w;�%<S|��k����־)U�<�g�΁�`��_�5ul�����qfs�*�&���S�󒲷�`-���H���&[�n�o5�ے�:�:�;��P���NH�i���6D��y�w�����B{�~>���t����l*~q|\�qU�V�WL�ތx������]���=l���]}��T���:���a�D����dr��פ�]�{-�Z�7>^�7=���nU���tOd�pF���<=ٻ���/�7���7����G����k��2X�u3�E8�}(�+��ǿ{=T2~��VNyy2LYS9/�n�:�m�#S�G��9��/O��Z�{���Aਨ��Q\wkx�E�ou:��'^3	=�ѸUz�d���x��e�g ���6v�v�V��,u�YB�W�� e�=o��C1����Yɋ7]e:�Ĕ�Vb�VL��m�:���3�]Z�������{���z���lTk��������yoI�꩑jʙ`��8[� X�Dx�y�x�ٹW~�Y�֪��o����<��@ϫ秛��g��o�o��6x�SӔ��=�ڼ���G�j�w+��z���{sŲ������n�7O+~rj�e��	}]�^���w�q����Oi��^��x�)��rUO'I�~+=M[���S,���#��ȫk7�>�6�P��Q|�Fs�xߩOU�C�[<b�����緰��V(�tc*C��T���'{k�gq�C����3������/��ڞ(ׇ6�x�
I���K9Ҩ�l��[��ԿuJY9�\��U=�M�J���x����qw��R���9�M�{�Ϸ�}bQeH2������X/ɥ�w��ɼ��T}7�M�Ry�/�}p>��P���נ4��CR%��*�=���t���s�H�{S��$[I��>�TxA{d���y�;���h"�$���^R�rk�r#7���~�{�;d���{�F.�1e�=\��lK5Ю����D��:����]z�3[��n����Re�]����ꪬ�^���-���sk��LfOd����1cp��r]�]0G���t��n��w�����J}��_=S�_�ΙT����N��hm��r�� i/+����	�����q}��O}&���.Ni���D7P�w��S�n�͏O�����|}�V�z���x�7�=�;ӷ2,Bv��˨x�����{��2e�N�J���[��rپ���O�{z) �O�'���[~])�Z��rUO)�B�l�]��T��6���P��p}�@VE�����d������/j\����)n�O<�ȳ�j��>~�ɟDY_��ur_S�"�L����_�|��U2⧀k��zTnܦ����k�����{7eK{���
q:NS�/�W��%x����AS�u$���	�*����Qˬ��>�\w@<�}�:Ny�Z��{?�p=y]��% j��AYo��Q�Y%��Y-�)�-:�e�۴��Vb������[��x`�*�|�w&�b�϶8��ߨ�7Ql�^��|��-�0��|��}�/"�.�ܤWJ"��<�H��s�Rg`Vu��cR��Yo�1��ꪯ������Br��?Q��m*�����v�����.�Nw��@����n�ѹ�Q�vڱ+g��xN�?�_)zr����g������>�2�2�V)�k���96_��zy�K�t'Х��7�B��6w�V��)��{�s��Nï|d���S�{4�9���h���w�}�� 筀+W�s�帺����a��D����]� T��N���9&�/?*(BT�w��=�����M��ގ����\Un�j]��_?	G:g�zk�ʵ�N�z{�����F�~�m�h����\���ڧ�OeM9���4��V��+�Ĵ�u���N��M���m�8:��"y���]q��!=�;L�'zn����J}���<}�)Ɣ��N�����w��揳ܼizT�}�3ˏt�����w9�j��bʩ��t�_sk4x/��o?j�f]Ak�x��k�!a'nˮ|�R8.�.��ݣ=�=�%y��Z-�*Z����?���=��-9�AGv�T!Ss�|�x�܎Ǹ1�N�t��`�����2�V��ٳ\�fJ��i@$З��N�+]�ls'�8����W�}UU������~c�R78{��y��f8o7��G"�2(���g&�C���$Mr�8�߾�7ϑw���s��Q�����'&�FOM{W@����Ξ��l���"]������Jkv�܏(KuK�9y�ʴX����_W�dj�0=ez*=���/��:�w=&�݁�G{�ş8�a{W	�廊m���M�=����Ol�>���ުg$�&O�13�"�=V�������K(����_��E�S�S�Sxd){�%�O�[�VU^�Tܯ*{ɏ�s��6*���:�n'���I\�q{��̘��<�)N���+*��%eU�Fe�s�*�&���G�	�y��(^��W�.|�[G�*=�jV�vy�������t~�����;�,����:�������U7y6�z��=�tkPp*��~rP����@Wa�%S�W�7�uXvX��_Kʂ�+n^Tԫ:�6 �8���@��+���>���X���
c�7����ò�\3_N������H庙,6��e%�5�d�FA }���O��*�:u� KfÒ����ﾪ��k�l��5�w�vy�Y����<#!�����Idh�p��6�j^����tl���7��'���v6ǃ���������@p�/s\�ڽ�3'�����T�-M�qo.p>Q���;�ׯ�Yy�W�iU�{�`o�Bfx�5���ݒ���z�F�����d���rO;f>��������a8��v
�>,�t���9�P��v�������"��z��xd��?f=������ʜ�����}j�����V��ǟKQ��{ʏ\ʱ��Dm�4g�[8qo�zWF�����eKhZ���Z����67��+�#7�7� D�̏��{�Ϫ�d��ꆜ�ٗ<_�]�^��\y�	~�s;�&�����5���]y�U8�')�.��j���յ3(V 6V���Օ�z-�]/w�o�[y�2wz���hZ�~�Wzu��}X�߲���hf�(��}Fgr��j�u��m_�F��w���SX��Z���I[~�Cr��J��q���W�`�w���\m^qޛ������H�=D����]>��mq2\�W�ȽR�=yE��o�pTS���8����V:�}�Q�Y� ��}��_}��r�=�8���r��ǳ۽�����Tg���^�����uow����3�X~0s�zq��;p�r:��ev�W}���yx+T	�R�[�[,�mX�5��?js����C���*�S�o;�M1z�+��}=�dQ���ż���{�����j����Zu+2��*�,���r#!��K���e�{QOo�y����y3�y�|Pۡ��}��>7Y+�{�~u}e�^�Ll=�����Lfss�cR�ڥ��z����{��J+�|d��lD���*��§��g�N�y^��y�b^je!n��Ï�{�eFU�;�lh�;��ʺ��3�=��t��_�*n�A�����s������R��*�>�Ը;����3��'s;�n��t-)�Oy����j��4�?SB���y�܁�%8+9�x�^Q���6^�|����m���Y톳f᳒���h��}��d
�ޚ���bQ�o<��U�B�M��׮����f�O#x%��7 �v
:�D[wk�їul�ai�+M::��]�\'�!T�+(��v�<��ηP~�������_}�}_y����o��������vS1k����I���)n�O<�Q��[���y� K�=��}2mrT����#�_����*rj�����Ƶ�g3�>g�\e8��~���^��u�v ܇\N���K�z<�z���ع��OVfzL���_Ŭ]%��ǡmo����꼧=)v��$w�Gh�����(���=���~U���v�fWq�L]��F}0��t{�4�'��ؚ�>�`M��Ξ������y"�*�T���6{x��t�{7���V������w�H�'���&�o�{n�4��z�!(�k�/mB����<��Y�??I;nfD�\wufrH�����o&������һ�����e�~}*{�P�r�Wo�ƒey�ގ(5�\��<`������~꣝2���ɳr���[��c�d�6�ɛ�n�%I]Z�S��ȹA�P/lP����.Z�S|y@ۘN��>��n�5�a�k�K�>������Q���*��*Y�ŵa�i<�\M���ŗX�1�sU�Y9�Q�������bΧ�nn���*����(���������[�s�.5��w~���(m�����־�|��D��4D�Λ����nX�����g�7�eG&M�Q�clput6E�<�����`q1�]�Ͻ9�N�~m�%T`��k����c�)�Y�����
�c�u���_ٝ��'j�����ߠǝ��9�_T�1eL�S��S�[�&��������]!�?aNZ�=2��l���׹�~r^��ȕL�N�8�:z/��n�5����px��on��@�w�R��!��K{�U�������N�6����^��S��� ����j����=ҚU� ��g|�2�>�fu#5������g�j� �je�^��������k�{�Vrv���t�I��ISn�M*�OҶ���~�0y��T����q소���zK>�����Q�k:��=V�;��ߨ���m>��O����W��"q�m���o}}�&3F����.k!��8���
�T�b�5�
�pp�ia
"GP���bJ�w`} ��V��Ŏ���G�)�L��n�&�S(�%_a���T�
g?���*��}�%k��"e-*�^G��ᅤ��+ZP���,�}A��+���ҷk�wF��j�*=Q�-=)ӽ,vb�X@�Z]׼�M��}���T�n�|�'ƥu^	-t�@-�2j=[\�p���9`ZX����n��If]��M���쬄H&�ٸ�$�� ���/l�&�K�1�{{F�d��-���=�k����g�G'�&� `�90��Sݾ�p��������~I��.ڶv��Lи*��7�x�L��$^u�i��M3��%+m(漾�S�]��@Q·w�{� ưtKS��v3�-��l�@����]{ 9�s}�V�:}O

���Ѳ&2�sƫ;��7����'����ʔ�m�K�]�k����Ve+:�M��M���c��<9\+�3,J���$�i���֭fV����9y�R�ȋA7&6���}3�`Cl3�� ^�?>+I���&lÖ���ۜ�7YyQ�V*j��>��}7�J6�vR���m�46��'�Y�'}��Oio(2�wO�ǘm�2�T�1;���焆���N:�iͽ��.�����Z5�`�n�G:��'����WwSz�}>66u;d4C�Թ\�nHn�-��W�@*�;2��:���(�=��(ѻ�ؐ�E
��������b��Zĥ!�g1�ZG��1=R�VY�w�762S�:0�@M-��jN��W.����)�:FWA��}��W n�.r�Fڨ���0Z�^]tV�D��u�lҢ�&4�5y�C�{$X�f�;�61H�����w�9��s�I!�YLb�si]Lbc=8Pb(�l��ɝyg@�/��<�!�-ЃH�C�IR�wp�:NG�`�i���X�F�gf�ٱ����l�.�����j�&��t��VW6�|g���b�ۿC�؎.���%�:^�TA��$��55��X��o���A3ٝ��R�Q!.���r�W��:S��u2�#,��h�8��gs���Fmh��� }.�����-DT�yV��o�@��@�l�Ϯ��V�}��c��uۑV���
h�ʲ])n��B�J�L�O�E��=2ƸV]��<9x�:T�f#;��xI�ӌ���4����A	|��`��aLݹ�+X�i�ҚɭX�E�;:�bI/�r���a:�m8��z�%��s���x_��	/���U�"��}��mՓ������K�A���1tQ�Y��g@$+h��L�P�N��Q�f�Ǵ��u��g(�r�Lt��u���I\�.v�y� U2:ϲ+��g�S�:��wk�w!E�A"�<���^I��m 7�m��u��Ś)e�9��(ˢh[��)>��8��<����vY�7ln���,��a0���NzX���(��*�F��5���*�kDA(����*֢��(�(����ʒ�h�X%�b��*F��U(��Z����m�e�Z2�*� ���U��KJ#e�DE����PE�jѭj*6��*EQ1Z�)R���Z*0�j���JJ"�j"5"�ҫKU���l�2��UV��Qkl�Z!U*6�*##m@b��P�m�(V����Q��PR�*Um)[j�X�P�F��mmb�mF�()b
��� ڥ��jVZKP*UeH�j­,�c�+V�Q"��VE��-���-��(��+Z��YVҰ�*�����VBڕ��HT��Qb�JT��[J5��(UbժҖTJ����eV
�`�jV�	R�X��Щm"������%�ʅTDT+-�kAQ#l��dV[j� �_@P���:����;�ۋ6l�Z��KQR��WD�	j��h�jS5����VSӖzml�:��л%���^�����W�ܵ���}������Y�v7�_�K��<�yo)Y{��Y�=�*���&�{e�d�D���i~��΋-�=Fx.��n���%e^�N��q�Y$ݿ3d�]���jRd����UO]{��|}3�ꓭB:���pe늝�����&L��]�ֵnt���/?"���mU\FpN�������f-���a�s�׽���yL�쩣<�sTP��xF�=l��\;ۜ��ɫ��[����g�w%S�.��1���z&��mӱ�<]����L���v'ޗ����}r��q��级	t�����َʪ!��W������V��}{��(/EF�Z�j���S>}�S��NyqH�T�Y�]D;�'6���3��ۢ�F�D���s���.��s�v����O<`�ۚq�5�9����j_We;��k2�N����@�+Ѿq�^pW�Ӯ��p���P�b빖����y�\�]��6^���h���g{�b��V2�b�vq�A��z��'���Գ���Z<v�#�d���y�b�8��7"��u�v�f�u�n] 6�\�Mv�]0N�yl�l�2y�ﾪ�����ߺtŽ�w�sr��k"��Tv�8Y{-[��fǳZ���j�%��~n���y��d�_I��.���uNMS.*��K���ם�E�Lի��).�q���]9�����߮��xOd�=P�����j�����ң'w\l�n��IL�M������k}�7�k\��k�z3�nޏS��&o"�4.��{�<�}����_3�n>R[�]<�+�>ڏ�v/K���Du��@!�1����tݖ�|�=<B�U;p�v�|�V_�J:���뙸�B��������ޏ׵]�y#[
��lD��[�e>��zj�#�9*�Ź����a�	|ڧqfV��=$��)<,^�/j����9�o)�6E^��ls_g��*.�?�|���NfOd���^s6�#�G�ׅp����;�"O��J'�ʞ��p'�@����L����p�����T*w�KK�����~^��tK���/W0K�e��J�us��ۺ4Y�+�m��,�۴��|.��$$�g9ÁY6��tZ���t�Y���ɳ+f��G�K4JǂQ��&�c��V?�^>��Ci�V�8j�G�J.R�����5/��A7?}j�e�{h�5��T��o�	)�/$�r?�S������!�����\���clp�t5�k����O=@g���l�OQ���6�u�] ��~˕��1c�D'��5�%_ßm
~��s)��*����^"�>���B߽)�j�q�E/˪g&���kX��2���³� W�=�cҐb�w��s\7���[��]R綦S��X�nP+z�K���v�ݞjK����_K����u��%I�����9Z��2�>}�V�&���W%��oS~���>.KUp���?k��ջ �nB�q:T�?}u���`R�=ܔ�xwB��9�.��2赝&�f{���L�_���J)O9�;wa��$��lck�/����s�`�����n������O-�6��P��X����\��$�IU���S�+�\���S���#���5��R�;t����Ec��+�r�|�й��]]%ioS����-]��Є]�s��Y��8>�{�ѥ��3hSJ�,G;۹�C�qP�5`Y6�˃S��MY��x������AF��=f ԇvn����%�rм���眍a���j�zt�ߪ����輽'�ӒOq�ղl����s�z/K߻�$j�����ݵTv$��=����gow�����D��K�/���S����9ǹ�'m�Ȃw��H���s���6x���������e����_}O䳦__$�G�{��m���ŎUz3k�86�ӗ���ڦnc�w&WH|�Mͣ��l`s����z4�(m�	�j��j���u&Z�'������y�鏘�Z��=��D�Uۧcn�pl�s�x�*�/�x����~��֛W�sV���X�Q�F����n59U�v�6�M9D6w����L�ߧ���w��*g%��wTС�fZ�u��%�}����	���[.�s�O϶z�\��kݔ�Z�]S"(d�\��q831>����ܫ�hbQ�֪����թv�-N�.���a��5X��x���6�%��i^�w�;x"�V�ƞ=���ka�ι�vo��5W݋�{��AӍ���� �K>
������A*��Z�Z�Lד>�cj�C�_Z�b��T�2k��yl�C�V@92�7���(�8Mɷ�9��oy����}��w�d3����t�j�� ��v*/e���_���Mn����X�g�v���=�M��P딩�~�NW����E�^�������z��:g���5=��13��^r�8����zڸ�5�슭�$O5���s��{���׊QY�rs��9�Ы\��ߜ��ҽ�^����S�(����첔��T���w��Wq�G��'YW����{ɏ��7������a��x9ѵ{����U����5:>�(�dws�T�YW`"��g��;s6�b����n�=��f`3O�����#��{\���4*��I	��O��.�g&�����I���|pe�p����8'Y�8j�;�[^���.��w6���1�=�4g�ܹ��<#Tz�'e;��j1w��+���{f��W>��૴9�uRsfU3��D�}Q�co����HhDT�[C�sk-�{�.���� F-ɬL`�͍=��rS#4�;�:�a{�Mt��;�@��KC�B�=�>�/c�v�i<cg�ٻkH�:�^h�����d2���u:�
�I�v6Ёʝ]�Q���C����^Ru��]�&1��WA2�����}UUW=3]�fws]��O���W[a=�8GJoK�y8;dCn�~���Y#�=��{��']Ef�g޺p�ɯ=}Pɨ��d痕��1\�8�$��n�}/�gg݁۱GxAuG�/�t������'>��y��l7�+���B���Z�?�ˣƵ5/fS��kX�tzu�����\f��s������(�#:����mNσ��NE��MS*;k,���އ�C|Ίs4\�r&�������{���Ku��ɔ�����=]R�S�X�>|:�tz7G�!N
.�M������vτͼ�������$��pQNf:NXgNS��U1(/���w�پ����f��
��!'���?����b1ܜ�3��ټ��+S�+O��Xe:�ބ<�cLy������:>U,���<xg�q�"����0=s�[���p������e +�/�s�/k܎��_!�=��~�k���'�����C ��*�ޞ����Ԏ��nͶ/��RuO��4Z*�oW}�q�w"�)�[�8'���{wWU���L {�ʅ�egV��@Tcz���,�6��K�� >�}ekL�yb��C�l\�
�A	f�_6ﳜ����C6<9Ra[-��9w��諭���G��ro�����kӅ�{k0��c'^�0O�c�%�2|����t)_F����knO%�d䋰�_�B�,�R�be4�?^�A[�Pxe(�4&:RXϖz��u�v^�nq�߈�et����P���0��|�_[��3.x״�y��p���Z���on�˝9�f�/7���>���ؙ���@��D��M�
�g�L�̽��*�ʽ���o�A>`ʍ&)��*�`�A�U���]��)	S�T���D�ݐ's�]�ٶ�;^����Įb�
�p�Q[oSn�����^�G���o��NT'_�fq��%�={��&xg��M2Ȋ�F��*Pʢy�ʫ���|K}�T����j^���u� �L[E��m+�sЗk�o1��LfT�U0X],�/�\N�ґ��V���rOg��J����}�0$qV�R�i��n��Gj+�C�,I���Л��3�ko��p�2�K(V��������T��O�B%Z2���-�]b��������<��栍���M��*�j�(�C�)mf!���5�K��`;v"�f�m�Ǣ���+��7�H������p�Â���3�m2�N`#El}5T'�q���r�D��s�C���>x콴�4�y�m�s����W��Cr:���E��U���J��G��^Z)4�,,\=u�ǌ��=A�����;/57���w����u��:���c�Sī�e�0mu���\�^�K��+N��A��wd�����"]�7y�'�X�.�7����\N�+�l�J�W��y���H���Z���{J�c<�I��(ڕN���jP!�h���9]�[����gU�Y���o�����ќ_�I����Ʀ��\/O#)�U�X�pm=� �徶�KV�~aY�@�9{�0=�N�sL����I�����pq*�[	�%(c��R���Nq*�.�+�(�&����f�3G����W�*Ħp��w�<t�"�ר� zX��YS�SM�4��}�.�@�<<�\��9�V��s_��g��B�R��F���,���!�2�������q
ṇ�^�ל�6�����}��.	�U�0R�n9k ��W�3�c��M���c�n��b����K<ދ~���aWM]�����dt�#��,\�
���\ϲثo�W`b�B�+�����[������j�C8f�c�},I�+!/ttOT��;X�|7��[�N���}�8,��n��>�	)f4���޽��`�
�Z�Ia���h[��\�)��|�֫��:�[���u��PoJ��\L�ytAi�6�{���U����{ͮ)�*?�l聫K�5^|.��'՗�:�z��&2e��b2a���Y�ym�k3��2�W�B����)��_=>wzγFmӛ��O\�%\��U����[��;��Y��O�'Cf]*�s���>���Y�E�C�
Ӕ��4�8�j�Z�Yv��#e���m��4��I�Hd����%/�U �y�s�E�	�U,��N�v�O��s*��#����ls](]� +W�3�>������V��k������n�D�zɾ����{Z���u3l��U�#(���ئ`Mm\�V_o��О����q>�G�7���1�s~����
���_9V����E*�0�ՖNz�x���g��J_��9���u���,���{���U��k����!9P�1�:`5m��i�N���q�nzN���C�K���g}���Arxe|��)7)W��9^����+.u�*�=�Yԁ����~��}}H +�������*�&�)�~��&$I
}4�q�*��^&Ghڵ����	2�D5>����3�75x���9�k��u��/+̗�vI�e���[d�wte�9��:�%d�z!�T&[��<n��r��Vb;��[�����\|^Ɍ�1ս	�*�r5����m�}��RN��:@UU}�Wx�}+��m�@ֽkt��{ǽ5*��*�-���k�)�Nӎz�'�7��͵��Β��}χO�v`t�<5�E^�NPw��"<͋P�U�F��\Uӫ��9����O{���.�`z���>N��=N�	���]��ϯ�pL����K�2U���N�~cϵվ|kF�>��%S�0��Ӱ��f�2�����躛�L�4&����]�[���̩2������~�̺k�l+�=��0��.�`�9�N��p�x�͑�~zeFU�/}7E^�J_�Bh16��&4���S�'�{�00�'<�I�^8v��ai��y�X��_�L��>�V����"v�8=�F���əST�*[X;�˜N����O{��J�x8y�fpɗ�B�wB�k��=,I�]���W�{�q�/w5�E~��C�M諟�^d�	j��eLPn}<��P@
:��*�������'/,J>�qcj���ݝdB�wL�Iy:�n�S�pmeK�5TĄO�ȝUG��Q( �XW�7�lY"�ݞB�v�p�
O7�M
5�hҖ!3pD�+���,���1ٌ����p�/(;�y�����ᦪ�^�g�SZ-�f�u�K��*'V��G6%5�"<�]�z�i
��u�ɮe�|xe(�G����L�s�%�*��Ы.�'y����m{s,��k�����*�>8�I���i�vG��!�����I(�<Z��f�һB��g� ��Z��&9�|�E}x�Z���sJ��	�`�T������#b���il���L[�rt]�@�sU���t��FgB�#��('���j�ԭZ�G0`]O,�h��ζ�c���i��(]6�B�$wt�X���/����߮bv�sU��*Y�y�=h�����7�il�]e&1�O�{km	��>P�'}�)��'BgV>L�]jv�g��Z���<e:�;rr�Yu'6�]#X30�B�n�]fJ�V�ȔT�m40����	�M`1��jf���G[��G��`�I�cn�o)���8���|c5���0�Mc'v]>�(k���&ѿ�E�((�J�jP�6��Yn�)����ʾ�-1c!jt\Rh���^�y4�pt�� `D�&%}�� 0p����Wn��䉵}dk��N�5�v�K\h�e]�guUΗH�)�O��I�t5�Q��7t)��:��]��>�l쫗|�Mps��ц���w]ԥ먖wvUX������{w�;D�v�P��b�q�ʺ��%���sa�[��tp����L�)_h�훰�Lzo�e� ��Iu��g/w]Kw����;�}>
�a��nAlP�Ί�h�����ӥҦ$:����ǘ�N:�8^M�̹(l��҆�MF���,��G��6'v�+"˄&�K̂AJ��p��ߝ��8+�JK��I����0XS�Ujb�Ȭ��YUv�$�k�a�ռI�a|���8�5Aa�~�W�*�ѽ���lf2քeEPf���t�X��"�M��M,�dեd��#}���o18��̃���_Rͮ��&Xƌ��D�<ݱ��x�\��z�d/�.U:L�[s2��LɁ��������#�b�\���(\���i*ۘ��Q�Ӫ>�S+j�L`�N�,�4��JTDW!ճrJv�J�&���t�pj�=��T3�����(쁏����k����9�����D��u�/V�vg�Sc��\�ܳ�0(x�A�m�s�WYّ;k6a�}�y��i��=��Pζ^.F,�MK9 �j֯�'<���I>��(��|�r�f��cL����H�����+t�%v�'moV(�U��톸d�\l����
Wt5dr�gS8�Z�s��}�KV{zX8�Z��@�BJ�Z������\0���p�n���+�lε�)g�"��;� ��m��}�K�Մ�&�c^5���Gt�Ҷi������_ԤTE*%�
�e�QKB�Z�iR���[l�����A)H��Z�#mJZ%e[bմ�R,F�UY*%������iK�$�h����@�6����E�+
�" �E[(�T�b+Z�EKeH5(�,EH��6�(��խ�V��J�Z��cR��-�TP�`T�0�T[@�m%b���R,�m��EQ�*��ƥ[UB�j"�V*��YR����ŴhQ��ʴkj����EZ���mibѶ�KT������
"����*��l�X��
T�,PkA�#l��l��F2��j��mFЪ1J��T"����V֒TV�Zƴ��R���F�X��l�DkX1iQ��Z�DX��U+Q��R�"��d[R��*�il��V%eZ-�VQ-�R�h���*�H�kA��+X��Q���c-)l(5
��m�T��Ub5�jQAVQ+*

Q�l�0�Uk+jQe��cYm!Z%H"*�EXV",��EJ	��`}��Tn�2��,���̈㒲�3��pQ�4�.��*Y��� ��l�V
K,���̢z]�	�pj��ʯ���).��S�2���K���Н���neUl�(�s1�p�|y�E`�n�[����#t��7�h�� SC���p�����ew'<΋�P�땩��q\f����<��L��V�2�~��1�{Miz�LpR[�<2��@���W��C�����V�.�� R���������]J�7p:�mGJ�*��~�\�����^�յ�b�蟙(�S�^٦�T�<ƈ���);�ܧ��7A�����m!k&���ػg�	F�u�����kxß-�&SJa��q���H���p`��}�-z���<q��&l^u��$��	c��uu}��P��=M|�.r���4�o��UR�o:��`9��z)�͇~���}��|���� '�D���l�jc3\q���:ϟ����Y��b��e7D��A|v�yVo����H���'Y*�*���m�u�[���<��m�o���]�:�qnR�p�R!�8Aa�*�v�w��vX֢�z�ǂ!���X����j ���f�ڬ��S�0-g{�<�^�庚B��m��^|���H[��cB�֍�n�%��"��hur��X\.��r,�(��ʽ߯�M�Cݡ ɫ�����*wʳ�_�>�j z���[}��Ҥ�8���}U���c��;���1Y�5V����������d�[&��mjp�RJWA:A�4J�[}$���!��i��K�^�S�Z)W8���ȧ�O&3*y�,�  �+˒r����_���y��������>g��*�׍t��i�.a�}1A�*z�1c�����sC�s����>�WN���\1�Øx1�2e?�h�r�>�qu$��V���M����2z�'�I�Hx}���V����c!~����d��8`�C/�t�b8��U��o�N�z��cǚU�[l���]/*���eH�ګ�bB��8pd��k�y�{����w`W]F@p�B7��vY�Oz�D_\UǾ;�B�����O��������EI�]�)u�z��xE��(�Ǆe	�����*ݺ�m�x:�+�9���ޜ<��ɲc�c�c �T+��g�X�z�j��9L���['�51ݵW�
������LfT`��������g�%�R���WՎ�O�JOo�J��]|�̯x�XU=��j�I�1��� �b��M
�P�IеU��Mj����rz�s�j7�wP�bW���C8�U��m��Y}�h��X1�Qp�V8N�O1�ۨO5z�osk~��M�pZ�S��������][���V=�gF�l��k���ыZ$�7R�-ʐ#/�}_}_Rq��nd��˯~���^U��qڹz
ƀ��!n���ܵO�B�\=���-;�nԭkrfS5б��e^#Ħ���T���ZU�e8����O]�t����������E:����1���92�EY�H�]0�m�Vn�eR�[����>~�O>��;
����O*�K��f�U2��#��G�y@+���M���V�)�tp{�M*܊c7ŉ�N�)=�V6�\�_��T�#����^ŕrP~b�]�w�{��>b��v}s��{b/Mk:ⶾ�oKf�k£�zJ�U-L��Oiݞ��������Jyf����U]�Ϯ�ƫ�B��]=qĠ�e���`ZT=���k��:'�����\P�7�������J]���ܰ=W�3�=kf�������Y�����A�5F����Z���.�E�@�-L5�)��\��"�[��^r���˟k�9� }���
��z@����S	��T�U�#pF@H@v�{` ր�t��5qul��1򡃢�-\w�.�>uqu�@K�٦�{xN���+XElj�#j��#<{#9S��/�4��{wϿ������T>�Y0WS��+�Xy��NY�%R_IY�)T�CΦ�{�q���նp�p���2��着�עfE�z0��t/���W[�Q>j7��t9V����EzB5��u��~O�Q絻��Vǡ��\
��S��5�>����\�E|�dP�1�:`,�i!:��l�6��;��AP`Bu��~2����$��UMlJ���M�U짳5=p�߽��ǧd�������O��5�G���dL!�S#)yh��R�S����R�n^L֧&�½#]���;��d��_w�����/�-�x׈�wt㞧�}~P���}����������HmWK��Y�N�����_����|�"���j���xTk��s�����*.1�E��/CU�8�̺��M����qh���A����.����ͱ����
Ur����	zL3�j"ϐ��⼯.��ԯ"S��~)ɑ�2��qQ�TD5w��X/C4�u�r;�xA�s=�쬠d̅�����x��K%¼�}y�)���TxzrB�*�j}���W��7h�8נ�$��Ȭ�2�����ݱ��j���ͬe�+�Hk���,X9��!o|�S7�Z�|�Kq����z�(ŉ��O9v��%z����l�b��Sk~��;nmp	[e�ݕ0"�u��`�c�."LU�p%�M`�a����UW�U��R1�~X��H�r,MݚL��򮭉޶L囹t�^b��.�ҰL�Gѝ�������觏��m�TC�)�����c8)@~�%�T���f��o�����+��U9����+���T0-"+���[�� *��1�2�����:�=;�����JJ�7���:�9�:e!P��&2���k%��$ �U_SԷڴ|��y�^��YT/��A�� ��1��.��҉/�|����4݃6�O���Ny�۵�a����VZ6}5P!H<��ww�c����UѠ5o��ъ�8=sz����'��=ņh����j
:��^�J6{-
K.B�gj�C�iA�9�&���w���Iڳ�M���Y뻭�:X3ؘ|�v_�y�(+�R��n�`5
/Пk��ϻ9��ޥgD��ê�؝N�C��h��R{����)/q�MK�<R��l?6Y�MTT��P�5�̥���)���3Ӟ�A[�U� U���mq&|NR��������Nvs��띫�{-�Ek!e�>",��<���FV{e�Z��t�D����vN)�ܭU��${�-tݻڗ����O#�u�u7��v�!f���Mp�T1Chelk3R6l"�����r���p�N[����}���_H\^�Re����.�쬥�*U�G0�5�[����N5��6X���B�����]����Ԙt�b>=),��]�J .�. z�l��U38��(t�u�������~�����x:�8�Wt4�>%�GnA��D�Ɣ����S��87��̙���6y���r����4�K�ž�+��5�݆'UD�3*�_e�X�����l^��Dx���Ů���a�ه��|k�SI��	�N���/���Lʨ�_��bE�i�s�e������{�f�f����TR朙|��S�g_�Ǭֱ�����6G�� �\6#W^�}��w����^nZ�4�P�-.��T��[����O�J�nV�*`�.���U��M������� �e@�ɔ�B%Z���i0��^#��h#���:�3���%o�f|��Rt�X#!~�hC�>}�(�9�R_6���O<O�(=�t#vz��,x�x�>�#�mB�yT���*��T�n^g����4�9~�s���w9���}Z���/-[�5�OYjmg`t�1�o�r�����nvVִqc������M��z"�d�͋�}�)冄2ə���Fj���L��9��*�#��&o,z��C�,�̢�����X��pF�^N����������nrE��}_}_I�<������?��AU�`;���-�o��'^،5�FǏ�8Vf�9��5�Xr(��xE<�Cڰ����jP!�h��O��t_]yyT]��V��)p�l�#�ڔ�X>̗���q��{s)��Ⱥ�]d<����MLwm\8ZZO��5s��k���&Y�yW{eU�J�p*~JPzxT�z�����&���I�B]�q"���3�̹a�Oc��`������qr�_Ӑ�.B�@|�ؔyz^Y��s��z����M粶U	�i�CR3�W��W´U�Ug�̫�e�]��$4��c/��=oc����_a2�����6������ �t������7[9�̙O���\��=�W���%e��'���DU<�E*������s�G*��Q�(t����{ygَ/K}��xX��D�gܞ1�|X���"��'՗�S����;�E��o`%N �F��Y9�o�h��)�B�:�\�Tɧ�;�e�P��NsX��%c�;y�4�[{��F��5닺������W�/�܁�r�鹧Boe�?�ڹ���Г0�GkȐ.�f*y�2o�c��?df��Xj*�C�/��C�p)��ÇGR�P�&��C�a��r�Ǆ��p;���u�$º���r�}HJ���Թ��������Su�{��Sk,�>�F�ځ8Y�pLF�Ҕ#�M�Y����q�bѴsp�=�lhޫ̬�Į�_`�3��4�|�������#�!�Y���6v�p��k�����P���-�F�u���z��o����-���A9pR�WQ|�j��/�.�E��z�5c�nod�k�w�o#X'��<���*wd�r��F
�$S�R��ֵv���Q��8��\ɉ����w�u�/��ƫ3�|���r��t�oIϺ 5,S��3=�yk�o��!7��{'��:�d�'����q�}i:�]{2�|Ҕ��5JV�~�muG�s�D��P`�X.����p�qpuw�x{*kc�'��b��J��[�4&�K�kF[k2�^���͌%�	�&���m��u<�:�0��i�~�x��^y�Sn��z([w]+ڐ��֣�$[����|W�>%��pSttU�߆����-뎄>k7]��w�f�+BPl�M�Ą��OƲ��w^���0yѸU�#���B�Y��ͿL�D��;)�OI(���4��m��u*���i�ӋA,�V�`�W��Tssz��:��O���v+��M�cu�����kt�޼��<s+��_�w�X�ytk%�b�0��ҺW:hK��,3l���m�E�]�`�]^`n/�ꯖ{c���c���R��5�+�\�^�"�jq��u������pnW&�V&����Ѵ_�O����b֩G(Wf>ۃ���#���`d�~����AV��6+�ͻ�-˺V�m8�x?/�����\WV�p9\k��>�u�UVF���]j�9o�f��|6vy����aT�Z�i{�C�pp�]"�i]w]�����m�m>qaܲc{��h1*=��^��1��9� S���zx��a�Uձ��ɒ��ҼA�魥���b�J�6s��(o���z�&�营B�uP�F��x���9������^1���&rd�ʛc�/�5Q�^evr�`ZFW���
���+o��уW����#-�C����{{v���x�˃�EDw�^CO�"Lc�pmg������[P�eI��[�%=^ÃD��Y>��Yc�^|����o���IU%�E|�c�i�.k��:h�Ǳ�g�D�ix]u�g�P�7Y���w~�;�g�w����.;����U���������,�ꛠV�p:���׎��.cWG���s_�#�F���ؘ�g�].��y�+#�Pu]H:��އ8�lp�mf���g-�e�)m��tw���7�3cȳP;N*��X�b_"n��"�h�[�����w?�ܤ��l������>�;�*T�j�A}��'�,q_n\�yg�Y�����}hQK��U�^!�lQ��)=�qH��bM�	f��>�{pI�.�}N^���r��o�Y�2�A
�H�e���q{�=���2��M2��p�^\�#0X��c�%�U��/+�b%f�R�G������M�6����L�U���R�W�fR��wqL���ޑA[r�
���u��>�x�;[/c�w{���ЙWz�%�<�]]n�Ao�������W\Oħ������Ad������[������åU���O���ϒZ=)�u�p ��C`��0�������6�pt׽js���[-��;�(uU�ɡ�	�0*;p<���x�A�JBE�����oMyB�vzI�����ewY��{���f��Ź�p�Hk�>Aa���2��<��X�1YWP�Ν;�7z�xȀ��}絛�6�T>��]d��l@������7����vv�ĴR琧Az�����}r�����U{���s�*L�q�O&3>�@A+�:mJ�	O��r'���[ko%՚�c�|�C�SF����DU׍Fz�j�
S\����hȯ[�WT;կb��E���9�Tj��VVa��(��wt8�v���j	g��.ˢ+&�Z�%7��@���*�xu 	U��Sf�NG�KPԽW�U��@5���K3�VtWUܷ[�pb�B>*oT�c?�}� ��iv4�p�״��u�
ށ�C3oVg45�7b�Dji�3�������l�z�uV`��6cE$Ȓ�{L5��`�ưMt뻻53����Tfe-���S{:�Y��R3��ʻ��mQ��^n�J�����E��dn�J�`��I�Vu�2�T�� g8��5��΀�Pڨ���%jNu�Ŭ3*�-��u��u���wZ���V�[�j�{oV9,{V)�]Ζ���+�:��!�����ܮd����z��j� "G��s��_wS��E6��-;�\5�~�RNŚ�׌�-sT�1G��ǩ�V,ڗ�[m��n�ŝ�N�!�%'ou��㙎#7U�����2Vr�P��w(g[93��k��&�!]ͅ���V�|��X���w;�%W[���9����͝�ιnE������v�N�u!�;�%oYgd�����R��.����8���E��w�.ҵz�5��Y�!q�v���fP�(q|/���r����fDm0���h���I��8�%+-CÆ��+��s_u�[[2^����j�h8p�mBOr�`�MX�A�Y����a��/w`���֕8�v�w�I�Y�S���v�����p�U�r��=!㦆L�W:�9��C�Z�2���{����\�7M�-�J?9շF��e��i�H�\�AiB�]��3;��"�$����W5�v3!N�-�u�ݜ�a�m��d!רIC�^�ח�`�Z�W^�*6�ݨMC��[�S�7d�h�|�"�����먣�*l^���\�'t����%����>W]:�!��bg2,S���M�L�&���4��ޥ�hE%,[o(n��iͨ��'IB���w���R��X�܁�c��}xi��]�g
]Fde��Y6�����]r���â��q{��6%@ٔiQ��%�3��i$�V3��C�Y��v�o#١n��:�{}YYʉZ#7b�/*ͽ�^T���:k�.Ji��1��(J]c�յ�[ڙrX[0��g��.�p��rɦn��K�lB�C.�F�+�ޮ{Z�pۦ�� �ᗶ��N�\�	��D��}R]"�Xi-ܝ��f3��En��=����D��ݑˢ2)��-��3�7`'R52�v�%��B������ɺڇb��^,�2��ưT]��+Vt��$�͊j���2��;+��_Q]0�:�[0�Ӈ���m�í��Q�N�չ�ڔk���.ɺ�[���ۢ�����m��D;�n���3'8�]�;�����0�j�M8%�T�q��6C:C�9˷ia>�Ƴ�6�ǧn)�cm$��l`4�6��J��"��clF�JU	mmŶ�Hȵ"ʬ*ŅIR�E*����j,i[TU�X�c���-
�֒�,���Z���b�E�Ab��QkR��UT�5�ҰF�-b�X�T�X�Q��EQ-+Q���%aD�0�*
#++"Ѭ�4���aQjX�F����Y)i(�!U�H�UcF��lX�F)RVV1
ʨ�*�Z����)D�)U�m�E�*�V*���-��R���+�Pm��T�d��b¥d��Z�X`��j�R��R*,*F1A�EYE��J��IkJ�Qaj�J���UB�,m*VJ�ŭA@P��QB�Y(ńR6��E"�լ
!R6�X�#�g�G�U[t�C��֝��ֳ�B%l�b�xnJ�cf�۟'�M�r`уk��"f���?(�Hkj�)Ȼyty=YF;�}I���_}H�z�N5���� �/�]s+��
�Q�<$qW�6�k���-8��=��_�W?7ȼ�'B��ޚ�����i��gA�XRk�{�d��s(�b&L�W\k�ԥ�}+�y����2�'K�����*z�_T���|��2���M*?YBx��s0n�I3u�C�|h�-��Ǿ����7L�N�9`W�',x���Sʮ�!��5���򥋿uM�����|�/�W��l�tDZ� U;��	�`],'��vY�Oz�D�$�"�g@��n��֚��j���-�a��u�kR�cF��?o�t�z�oy��մ17�W6�Wwf4w�+�"Z9�OƝm����|%b�����^���i���Ah��v���M�Fq�JDl��,��%VK�|����o�J��]SS2��#�Eg�]㜚)�9b[hؚ�1�S�SaK~&x�\�9��`^��P㝉�d�&]��}����{�çܹe:r狆�,bƫ�Y�´U�#�|s�k�U���0Ê�2�Z�c��N�J�a��n�R������^${s4B�S��\�;y</u=���4ؿV��ɗue�I�V@F�#ū]{@������]�`��$��:+lP��\A�����gH먖b��Y�Q�s�*��5�۟<���uE��������9�'��{��G��&m���ʞ�n{�pY�}�h�Tl*��b;.�T�ޙu�lw���ί��W�����%=�N�$�֊ߺj�>|.q���U#��.aӱ�ٛ�7[��t��$�6���&VR���Iߍ}�.��O{*�S˝����ә�c��e����t^���dh�а/�fB��F�r;f�V��K'̰�N�s��L�I��f�k��:?F:r�tW)O2�~���� k�-(GǦܬ���q���;���S�/���)�v)�/�-9�w0�2��i�dus�%�Ԡ�ڨO�I�������������x�cx�V�Ac�`��**5<D��b�"�Yr���=�-����cx�����l����� J�R�"Q�\��`
�}5M��A���~y7z!�"����`�=ՙ�
�N���gtTOW�@BAS�oIϺ 6�}�>��D���klr�T���Q�9~9:�=e�Z������
��^'�\�E=��"!�`�嗛��sp����/zٱ�"�X��\��A�����s���'[���@Z�/��X��-�71��|d�Çw�$���o:�k`��:� z�Η^�Ƌ�,V��N�˵YC{#��Md���;��j��|�;z�_wi;�V��sm�K��o�ޏ�d�=&������Lz ��XX��W�xe]�ʚД2�_�d5��-#��b;3������������v�}��,���w���{e�_!�__dd;��z��7������T��T�B�9���I�u�xWz��<RP[S(ƼzA2����M��I�n?x��-�C��')jbcS0gK��NK����*�ȏ��<�r9j�E�d���m�Ƨ�]i4�V�냫�[�^�"��=T�*�6�S:��z����}��K��-h�|[�}J"V�G(W7�%-�8ꩨ�3LN�x���e��){��l�q=�`��y��}O�UGl�<$9�DCW?\�c)`��Y�d)2c��Ȼ��-�ܳL6T��)D.��6B�5�㔨�����V�C��$�+��Fg���d1�xK��sz���Lb8 �X��F��&����fF3��|�~ORA�=I�W�I����7�Ph���M���)P���P���^&>����~��5[~W*�urn5���P;zeu�_Y���Xq�괵([M�w�8����k�ずj�VE7Rܩ�w,��n�,�M��%w5]
�A���<���v*i�+^�8^rԱ�z��ZH������X�u��]���3��!������,�*9���^evr�`ZF}S��
;/W����s��� *V�>}e�|�>+����S�3���:���~�&2���~��SS�a���t�t��W�b��l"*��#���������PgtTI��F�*{��%2�\q��Vf��P���:��LJ��>3����Y���y���ь�e�r�o�Eۛ�x����YC��ԫߧ�������)mAGW�!�X�
�CY�"����Go7dr?c��f��dz����ۀ
UNyv���U3|��H^+[�O�0�_m�HV�L3�o�5bU2�UL֣�){T��xF|�+����Wf{���{��t��VÖo��͛x݃�ʻЕ�^9t�{p%�2��k3*��&}�Ja��3ӟzEl�]���FF��'���U�LO��}q&҈�����i_�Ê���*��PeT5�.E�3m��i�<��'7�X���o���}w�3�w�e(���ˀ]�!�E��wc��+)��(�t;	M����9�f���˒1�p	��;�N�c�$��^|�[���)v���cSjM�B<��kp�y�իո�}J�,'3�:�JFL���9�k��/A�ӹ	Vs��N�6 kI��������neM�|v�[%Ȧh�%�Q�"�0��Z-�Ѯ�v9^�����9������R�{<���[�0{�����f{;/�]�x��"c��'R����랗
����w�O�Tz���H9�|�߹׻��s	r�}/T��]I�k(z��������E���
��ca�Y�qo�2�i�wN��=�VWL�<w<d�Pkکj�R�9���N92�P�Pwu��k3{����	S�~ ���j�_o�T���#�Z�R�i����(�6�ϳΡZ[�G׍�\���	�`ژ,���}���MЮ��P>��3�G�e�V�M�ߏ�i�>���G�*Ṣ~�/A�� ��9�T�h�QэD�/1���¢��o��{��8�O��IT09v�m9`W�',x�x�>�!����*���׭lT�����(�<�ѿ��Q���ﻢ ��0��dN[ *�`y<�Q�
�
<Ւ�m��秊%[���6��7+k�:����oڦ��^�^�>����_ɩ�D�M}�hȥ�v�`o9̌����h���=i=]M^�IX�m{��w��7A�ڻ�l���9����Y��_�H�k���Զh}�mv�^"EJ}��P��Ne�<s��\��k8�yYK+�2��K�e�m!�xbj@N�z��B��pM���EZ=��[���W�JK�΢~5��S���-U�s�`�_=��:����/T������k��cG�E^e�J"���#]�q�h���ƹTl����¶�L�]w�f�_H�&�δ=,O�EiOף{��^��Q8$9n��}�� G"s�kj3<��}�|�pw[�)ӗ<]CR�c���x�,V�\Z6Ϣ��wx
�JXY����=ǻ;}��	�-�F=�95AH��S��ɶ��b��}2���\iLe|�?]��,�G��6��z=�u�p�N}�*���j�Y����;	���-]��,�p��O���&G/��PTN���\ʥ���2po�}�����9՗��L��:N�'��I�:��y�jG�a��l4������[��J���?<��9N��'����8[~�G��̮Ô�-�d���f���1Q�Y4*��]�\��ڃUm�ݭ��݉��������3F���g��s��[Ȏ%�^�~n�#t���e��q�ߣ�lEYe{n=���f��@���t�a�2d7�mU��<𖉾+�O'Y�W%5��-������7)�o�ފ�ʵ:ӬO:uK`����0J�rv��Qu��jP�����4�:DAg)Z�	��.~�k�7��<h>�4q��ˋ�$�%�P��R�U�T�j굌`i����\ސ����³��w����1�y��"B�L�#�oH�0A��˯Ze��s!�g��t.#w�|�
ˇV|����}��v���]�(�^y!��P��	ʷ��FS	��yfj������|XBê�!�b���L9qK�O��*�
�o�H�=[BE�ީ�۷R��lR���CF<es�4jۂ��;uA~�W��w�x{*k�}@�=�p�R,�����g��'Һ�ͺ�=T׺ |��^��˖���q`����md�~��-��U��˞�;�sI�zDM0�\�&S�
�S�5��gqu�xW{&,�,'�PcS��}�øg��w��?6+��T�:�i���bsS0{�tT�פ��o'(;�_�V3y�&��'l���2e�G�-�]2��
:�R�Wh����UmN03�Pm{5��W��3��r��B���S�o.��}#�x�|���!cS�f�-m���]���a�P��w�V�+P�u���>�#�s��"q$.]^��+3W)1Z��Xv
��k*��44Jοx�]��촺&&�5=A��U�=���E��]�t;�}I�f)�ݻF���:;&O>�S2�{��>�;{Ɯ��g)�B2a�k�v9��=��:�ռ^N����(�G��1��#R���"7Yh��X��۔�)߇��M޽����sȍA̧�੊_D.�|�:Q�!����bn5�&��J\[Z�q/\��b��[Y��d�.�����@р
��$h^�&PG����f?+�9;�䋴���:���'���+FK����O8e�E�^�I�_��2��\��B�x��T*j<_�osdz��\I��<6Wy2`�,�O��~��������`ZFT����[rz�;����=�� @
5Y�`*��ybT����>��̎e�����I�K��v�W���/�c��T��$ �~E�+at��R�.��Pv�/�w҉5��*�ҹ�����؞��72P�n�;X�DWpy�όΰ+���tR��+��Fה��t]8��^��Q����$�tv�T�'/��>�c��q)}P�#���Z&W~�i����������?Yڲ���*}0_=PI�'���^���쳇a�k�ހ��u����U�gY&nܺ%*�JN�J4��;P�)�o/��bX�"Y��E�bViuc.+ɩ�w �%b�����'��9�:[�ΎF
ᚦ���q��ЀT��<P0� e�33`5�`��V�uk�l요�`"e;�cX����=��yr�N�C�*�Ǆg���1�5�`���ړվ$� ��W�%R�9t�z�N�q��U�:��0�1"x����v�O�׃0��^��i��+�И�3藆=F�`U�ݖaw�OL��u�,�t�W<��J��i�P����S�h(v�E��z9Ww�eR�� P�=���f�8�Ȏ���<S3�Lf'���
�
s��N�q_FD��c�A��Ԯ.��iyiN������Gy^#�m���y�s(9���L\����S�/E{�f��<��s����7�g��0e5��
Ωȋ����=O��CN�D�=��ȍ��w#�=��{�M�q�R�
�OC2���ȱ�54�ꗪ{-W
s�b%�8h�w��t���^�c�?  �2�� }����]8V����|�i��ek�׍3���,�ae���[N�#������=���Q�~�,��e��خ�������Xe�O%[�\���g�C���컬��I]��ZS��%d�)XE�х��w�&�$���~��ެJ�� �w��CY���&���{ݠ�P���/��[�{[�SPҿ��o�����4<
-���G6<ݬ;>&�w�\��L#,Q�2T�˵��.-J^Y��������h�,#�r�i��L�M���\���̗��r�k�Rs�7ɻ�;Ԧ�82��$���P�:�^���*�%O;Ȓ®�<Av�2��9!��LlG{����%Z/���z���}�V��� 9E�7���T��E��b�w�_��Ʀ��;�y[�4R�ұ��ٴVW�CJ��U����3���V�(�Ǆ`�/Ixn��.4�}��zJ�v�|��V�f8	}�w�+I]�,����|�W�bP�A|&�vg� �z�F[i"g�51�X����D
��:a=�m]����~��B��Y&V���<�z�t��(�嫺����o�����ث
��k�%c�����;�K�f�]�*[]�o����{��+�0�{lLj,���}Pԅ��g��*�>�\*�V|�g=��v�p���`q���@�r���m�3�z.Bf��E�ʞ���m��pY�W���J3��#�yݩ�rMO��8��mѿ],*x��w]}�&�v�ʴA��Wq��s��U�OG����#B�n����$���5�b�m�bu����ޝ�K�x��W���
Xm*v�۹��O�R	hOJ�[�gLݔ!7Q���S=�4�Ea���6�&��j��t�����.�т;�{:+Ρ+l�H�P0����2�y�}w]A�Z�"�s�X�ϙ��\�3J7)�vQ�%��=�ۧP���K�"�r����lF��4Ӿ��w=��$U�9EY�o�r�-6ģ�c���s��R/���Y�6���Fڷ�C��
�ui�RT7�9�+�z��Y������\9شp:�$<��ŧk�|x����-�Eln4/����{w1�v�S�ܛ���K]�Bp�ɁfQ�IT�,#j	7�LȆ�j]�5��F��*ȸ�M�8qNNݑ�nf`8�N�锴N//��]+�[J��Tpɻʂֹn��L'}��Md��uz�LT�����n�C6�[�kp��`[7����9�2�$���d�'���+#����iAg+������.�R�7�W��ϵ:㣄�Wo"���fשU�Y�b	�i�v��J.�}�����b{�(�]��Z�9`�/�I��]q��V�:fguu�QϷ@w��Ž2���=c;㶲vH�I������&���H@�i;&t��X�8���R��d�y�۔�m0o�b�&[�U�A ��
���͖��i{qd���V�xC���9������K1�mI�t_k�踹����]�B��Y�	�ʵ�/�1B��eL���˦�h����)non���CD&��q���#a1���4�����P�Ӝy� ���Qu�9M͸�RT젫Fu�R�j`	��Cb�Ǡɝ�R��Ӌv�9�C�.ˎ�}8Y����̴�ɋG�oEX��|�8D��n��Y�	O�N���7;�W�������$I��Mu(�xml�N�]��+���h��	�^,�K�r5:���������Bv��Κ}��M%���m*˭���`q+mc�#�WL����)��%@���Νl��ΘڮT9n� �Dɗ,5��#��X�@�­/�U=WҊ�t>ꜘ�Z�K	|�0y��MuBm�/6���:�Q��J
1sk�)�����qc��,�ݒ�<�s��9ۧ�B=&��G�Ɠ���c��iq��d�v��V#x0�l�}��JjT�����jV��7�w>�g�ݛ\_U�x��8�p��r��h��J�B�%�Y��t3F��W3# i��y%�,��\,�=���F�<�}�>���M�X;r�$��ûf˺���6n�cU{��͛�d���;Lwu�v�u�\�yF%�1�����[�w�e��ʦ�����]z6C$j�����S�^v�[�/N>X����@�R�{5��k��ka�/����8O3*��N�j_�	��*,4j[(�PD��QV�J�PX�l�cl�N"�q�b,�,V5�X�V��UV�AZ�b���-���(ɌYYRQ*E�k"�� ���T�TYP�b�EUB��Ƥ�VE�V
E�,QR�D�������ed�P%eV�.5ELJ2�a���`Q"�aX�"ŕ��aF,R�jQDe�Z���²��DBVH�J�E���E��T+$PX��UaF)r㖩R�*�CYH�Y0��U�PX"��E"[`�U`�KYeȲ��AX�����YTP*��r�,U����`���q+�kU���c-����I�Kh�Z�Q(���h
�2�6�1�(�UbֱC{n���s�ޖ&uJ�V^ZA�E�w'ӗ	�8�󽛍�S�I�qcŭ���d렃��,��K�e�*c��{s��"��,އy��u4�\��D����N�bo�v��*��"<.�{��ޓ���x�\��.�D,�f��
����57���f("�/s���g�x�N��#�~�+J����j��f���U�b�s���WK��2<m�y���~��A��,Zp�=���4�L��'�駈��Hd�`jyMT��\�{�������kn����Ô����� �}B#5F���$�w��E�O<�ȭ>�)�i����ǫw�.��4ǩ�����3�x yBZd�ʷ�e �{��z���[::z��+D��]j�j���JCK���;M�
̮�J���Cc(D]��0�۞��O����: 5,@��0��&b[��{%�'�|$EO����������쓒~�WF}Sw%���9�����LSz��J+��ʸ�:��=~��+�=1�r2y��W��u�z��%�աK����*��+�\iU��\�xs��A�=�+w2�V]�i��&�e[T_+���#n�
�묰&η��54+�Xg��pm�׎5��=�v�zg���$���U5�J��9/x�ݣy��賃{X9��MHv ����Ĺ�=kd���H]l�ǹD�o,��sV����'f�b2"u9��E�)���GB=K���q!^Ǫ0k+�L�;U���Or�9�IPݭ�ӆ.���y3|�d�q�I�]�hJ=��qjbe53�]?zE;�rr�ΐ2!푡�ӫ�����^���"�d,%B�Ю_O'K-ƽz�2o�����6)f��6�?'$�y��^7�;|4�F���~��}����u*��[�T��0��"|ǽ�K��q�4�a�>��CS���}3ᗂ�*;e���!ʻ�>Wb�rM�|�V���o]�M޾�]6}�}�VG��9�4]p�`ףH�G�����߮����Z�tzF)Z��l��\+�L;=������<��ys>��ET T�f��<L�Ǳ��0����g��q{y������G�Κ����,�O8`q�4_��h��z�C�]cYf�M�轏�gH`�'(�������'���[��(LSb,�TqV�R��f#�UC�����{��z=��0�,% ���9fC�)*|{x\�iT��Q
K�i�廥�+�:=].��1 ����s�R���5�'G��ո������i�Q�hP�z��
|m��(9�'�g	Fn��Ѻ�9��QK�w�ܷ���)f��xWGyZ,�>�R����e�|�Y�o�
�C1<��T���jY�h�2S��=�ؽ���ҭ�wPlWbS�,1]��6,Z�]Y�{~�)kn��L��RSJ�3�ۂ��y��9a��q�LJ��@�:�0�/�(#��u������_f�r����>r��qS����,=�	WS<�o���7V.	�^��e�	[����j��q�չ-����Ր�|xxG�z�@9��C�/�ʦ����Մ�iMɸ�{�Q�H�*}Wʸ*¡�[fCټ�J���w}4\�>[It�a[��;��\��3޽�`��1�ߋ��Xb�{}BW�ee-LLiL>^�X�;���Bٟt�o�E��O�U��'l��Ds��\�G�N��8�"fޗU(Ͱ|K�Ί'�#��s���7�=i�1^6.���/.�&I<&҈��t�wOh>��-sv���ұ���S�����­�3M]����Ǜr������~���g����(��HH���x�$N�s�����pLfY�N1�x�^�4Co;�1�-��x���7r ���c������䙠�"S�X#����̼�S�n���K��y��ՙ���W/9�[��C�E��l>��G`�P��8a��l���M<S=e:�Җ��I��Wi�:��r5�:�5��}���y�$�Ni�U�XϚ�i�ž�&��^l:��0�q��Mk+	���]�������摡�
�2�p̫��j�r,eSMM0���KU9��@6x�m�'IJo�9kԸ��c�0X�����5t��p�}�����L�}}�������>)��5�f��7KN|��=���0eOU���phz#Z�%5��_��=�{W|�Y3�>��r���B��E�)��J�Rއ'�}�+��G;�!g@��}�V���74������F{�y~���4���UI��r��PNX��۵9� K}�%�ƣ�}�!{����f��R�E�ۯR)v�3NC��A��0��F@T�[ t dA쥷+z��p9#�:��tO��"&{+�;�����X���g;�AZԠB��x@��L�Xf Ȓ��٣`
e�vvR�V;�^>��_�?�ۮ�l=W�5�|�a�~�Ѣ�ǎ��<�I�u_\g ��mg�[�a_���Ƈuf1���p'�̔:n�:�+4.�+���m�QM���}Y��&�ϻ�PePʵ���caՅ��rMR�����z�[Kw3�|P��Mv.p��V3�@�y�q;��z��,�����Z�o,�S�9��[]P;:湵��uWD����.�q8�i"gh�T�T��S2���d���� �.�͖�%cО8�iw7k�i.��[�g�����0&1q��W ϯm��5S�qM>�jB��w^*�=�l�-�)��{y��$�W��oG���Yn��p��	sT���S�3rm��F/x��.я���>ײZ�=�݆�.L������+؎O'ZhW�E�7�N�$�ֈ��]e����Vu�n�.�Ӭ^�,�wdp�Q�r�'�4H�eR�WeW'�����Ȉf����̭�[o�V9��8-��1ϡ����Mc�$dr:w�ZZ�z���x���)#�$�ڮ���>�פ��WX\��y����%׷�ޗ�V^�������ۦ�ߪ%��ha´���4�T˘rz����к���ɞF�2t����OE�����MT]�Ì����"Lw�0Dv�UL�)}2�����u��~���\�dp�� +˯��Pr�^�Ly����n�D�x uAv�z�!j��,ڭ�*i�v���Pz��Ǳ�]y����噙�*LT$ǱL5�h«�,��['B�r�H�/V�b�gI�E}¸��U���C*�P�����j�]�<b�K]�f������eS(TA�Vfc�sMD��K�.x�,��m�Ku��$x���7{�hk�r�د��S��U��U܆����;�w³;�Q+�<�����Ff���	i�~L�P����ԽK�������!�u�z�F�^��/I>�ત�»�y�����8����=�:��̔ �ǎ��4:ɏ�P���Z���0�U��Yb�T�^W�%�O�ē�׫����?zb�SՕ����>������:s��X*uP���W�����2���'.I!��Of��b��!\�&8��e=Q�Y^�gq��{�'�^���j!k�2yy�=���D�2�ΊH�^6�2����{K����Ʀ`�������H�u��'��������GX}*'�^�:,�L���	P�5r�9?,������s��W=\�����E.��o>����}��];z<Z#E��Ғ�}>EV�=B���K���۞�9���3<Y�(��)�e�e�4�p���L�8gׂ�#�Y�xHr��LWb����Y���v�M߼��5�ǐ��@���}��9���S�!u���t�=d:T
��g�c���)���c�m�v�}�Z�KuhwF�]V@�ܤ�e[P'�����z
�oT�qm�z�&lEud��t�EU���";�y90��l趒嶟y"�5��z���t�ku��f��iZ��c��ٸ/����E�D�zM�}�ڄW}/�ͽ��9`��x���F *K�W��@����̯	�9� _��*��E]�əST�(����|�������|k�g�y4��y�t���͞YW��v�i��p8�P�^Nzx0g�b,�TqV�T����a�R���z�*�;���'nG�%��ڭN˹z�k�����唕>+��������9�D�"����j�����^��0��)��IV��UK�5LHA��Ȱ�ve������(7o��p���F����o5��y�ϥsyD�w�3r�;NX]�߬����
�u�aUF��Ϩoo�^��Z�T_>�j�����(�9����Ahe�o@���:�.�ż�@.5��lA����7;V2=G��}�T R�<����{�����e��C�;9��i$��H��3�>әWpU�3¶̅{m	N�/	��C�Ǆ]�e�4�	��E��Wz��e�}��n�hX��ǢW�%/:�1^�	:\ka��-LH[��t�~�}��){R�6�!���8Ǌ�'��k-ȼ+ƍ!�N��vƤo"�i����X����z����cz��S���)Y{
{+{nN4Sۓz-廯��B+�6[\��uə�5��ahۥ�;�T����0w8�S�U&�6t�êtų ��(�aƠ�dE~�bi�H�����*x_��n��w�����ו*�Xt��t��b�oѽE���9|�UnfA﫮'��3�b�i0�7	G�,�Ih�u#�Wv���������}�-�?YǶaP�5��7��k�xW�΋A;�w
��0f@�{^����y����z%˱܄�����Hs�0�.��U8_qϦ^S9AVS���(�w��$�~�
�h�C2������SQM>���
��"-?-eU?G��s���qPf�=|^3w����w�j�O����8Bͺ���4���z�ײ�p�m�(�n�xwv��hG槎zy1���S�u��nǹ(P��W�r��=�Y���FQ��A��l3%#�y��3Pej�#������ H��e���خ���=��z��97������pu�c�qd�~�D�F|�}X��e6�݀�����oz]��{y~��S����h�'Dei�tA��%I��r��PNX�O�w�Z��G�nt�}-��w(������ʛger<ZW�3�e��AdJX�e5R�<5���W���� ��}7�_��t�^�3ztɚ;/s�H��
@���2�{�P��nQ4qt��Z���"��fՅ��0U�z7t:�H�NZN4�x�8@ ߝ@���}�\��F�K}E,Α�{�٢���U���c��˖3*N�?s@o#t��A�u���[����m���C��֥�r���� ��S�.�W�<=g�L��/�ۯ	[b��J�ȗY�Q��WuK5�	]��פ���6�{�{N���}�'=51�`���q����W}�2�'!�ik*9�k�e�1ǝ���h_�*�WC���Wg�x�S�~�'cѢ
���k�V=��r5����Rsfy���Vqs�F|�p���b;���qM0T��'���������c�w���i���#�g�̫����`�	�\��MPR�.vT`����1{ǣ��黰uM~\�Ξ��6}x��#����Y�ٔ���Ue��'�vO*��u�x���]��N��?.L��,��dp���k[k4������Ф�ƾ��4G�Lt�aj-����H,߫�>�����޿S��yU1�X s&CD�h�GQ��1���*S�**d��bz�b��ݼ]ze���X8�d�#A"�٫�<���Z	͐+��$�����˽��УY�����N�A��B�4��Z%fWU�AU����p��S��z���]:T��!�#S�,ۗ@VW.��g1]��%�e�-*n��e6��g�wN�Yzw���,����0RQ*�]?a�42�ل��g����v�*V����w��������_�~aWg߮��r�3-_��\9��O\�HeT˘fQ����-"��-M�͍�礎&[�b\9v�*� 6��#9(�I��#�2e�Sќ����7��t�7++eLD���	UP𞻃����4ǟXyy��%���	i�=��k�/i�u� �l���:��J0h�H� ����Ue�՟%!���vzΊO��M��n6�9	�{�؟��6 �eMս&Uo��pu�C\�Z�xL9Wd����t�!7|���~-f�+�EZN�WG�̔ �ǏD���P�X&�γ��(J-Y�����P�o6��w_��f�\9m�BUGz)}�R�=��(����m|�o��ł��wGr�����=���ؼ�h���T¼F;x$#�.^)ą{)���n�Y/x�t���Z�����زNP��p��F�^,W����}���^��.�jbcS0x���B�Up������
*=y�	�2���j��%8��\7��6#�"U�Ҝܖ nv't���v�=�<̓mPU�Ѽp@/������9��һ�5��p�|�������4���^�4��jy6���u	�IZ\{��]8eg!��Qx��� m�b�/5�0���i�|3�!^W��ò�5՛�j�g�t��CI���z��#�u��!�F�b�����+�Z�y3w���jcvbX�]��vn�7d�0s%�k�	t��Rrn4���7.�.*�ޱ֛͡��V)��Oz1]���u��"є%����թ���EuƑ:\щ����1w�,�Z��q||)�~�
Y�����V�x��\!�d�*W=��#�_4��[�k;XS�m����&+�tb�܏&��$xv�)�c�3��P�M�P�-��u�����b�����U+j�N���>�ώ�'4�S���v�5�'c�|1@̑b��>\����N�)�0rdh������:��m�a���𭏌]Y��([V�%�v���n��� 5����@t��Z!"q��W&-ي�%��@v'-1�v�tNee��,��a�[�E�c:��U�" �o=�w^�K{��R2�G�#˪!V�B�>n�h1ɳ:ؕe�P�*|����+���.�	ҹ��^��T�(�ԓ�6:�z����d���V//d2�@%jeL��q1�0f��Z��[4kw�J�կ4p݋�yRb�b��U�C�K�
��A�>��wd^�x� ���2�#�K*��Uz�̡�E������b̢�N�N������F����Q<U&���&!V ��9�1;0�.�1�*P�`V��t+���z����*Ò��h%}�#�R��ӳ���Re<���vN����Jʌw|Qg������P����Rf�,s&
�c���j�VI��pTu͆�3m� |U*뵷���[�X=��Q�q�r �����]���t��E��9K( ���r�\��e�}hs�c�Z0�Ѧa�ES/WT�j蜾r��<E�+oC��:�-��Bf&���+�uu�0���Z�*��Yg`<�cV$�FLn��,Қ�m�S�N�Ln�Ye]pk��{�0���ٷl�z�+;�x�<���S*b*�R�+�ƣ5�f��$�do<�{r��(C��������lÕq�W���٧1�Ԩ�-�
-}\�����	��E��Rwt6���Bql��m�g&�9���N��a���CӠ��4a�;F�[Υs����[���-΅�NY�fѠÛ��zWQ�,;[�-��D��n��D6�wc8�^���]��0ֈ`T���5�,�{��s��c�=��j7��������)}�ު�mL\��r]�&6U`�;��aEDEw�U.�Yb�>�e�rh4����,fJͲz���#ufH5�2)�]�#�WryH��Φ��e�4����}�|a�UUP�PXT�-��YQTUk}i��$��Fҫ*e��U�.fb
ci[lR
��QT�ZQ���c1��1U�1*#�����D��*��UZ��*���A����c ��P�eG��8��bc�Q`�Tb�����E
�m�)�J�������`6�1�V�h�*�&%��Xb�Z8�m�1�E-`�#(bLk+����qZ���K�,��TI�U��X�P��G-U��XTY��E��nfZ�����QXT-�����Y���P�ņe\���(��q�̊[a�30�(Q���\ĵ(�d�fZfZ�`��rٌiLeV`����,q�(�ZҍE
�301R�J-l���.91�-Z�Z��fB��#��"�j��C�Z�3)�.*4(
� �콢��9������rnҧ1uvq%Q�k%Jjf�xt�%a8��MD�̄T��w��VcM�U��\�M��o'�{	B���]羶p���m��;�=�jj��r~�-ƽ;���#}G�.<�C	\ܨ��x;��Z����cZ;Tdh����}U���,Bl�Fqٖ3#������>3����`f^�S�׶$��oph���J"1�]c���40!�ŋ�s�ڽ�0VO$�,V3<zu�VG��9�ʜ1J!u��GJ��C�����7��ؼL���=��k��&4���;�soa��Y9����}��+�@�f\e'%��o����"}����֔(�����]s�[�^�ܞp�;��dKF)�ר)>��O6���o}s����	��Y�IA�e+�c�WyB`ɱk#����y�;�EŴf�<9ev�ž~â2���=�O T����*��ybT����
C��pr~v��A�����m���xS�v��FǪK�5}1!�H�Pb�
����m�u��>WUfw>�k��ܯ�{�qS�eUIpQq'A�8��8����o�u�g�P�����ڙ�H��y��O����\}����R��Z����n���[4ON  �ʺ{N��fgN�:������}����t�mB�i�{��
�6�L�zc�{�ei�8�h����:�Y�š��k��+�h�K(�8'�j�a��f�R�Ĝv����w�D����;Z=|�"J�r��AS��t�WKUn% ���o�!;/F���̦�0`P]��T��g�}7�,��]��Zz���y=�x%	�<��8�����C��(wV{i�^@i�Zd+zД�\�&S��;3�ׁ�L��=�׉��{$�B�9D�9��S/����h2}
ۊ���LU���[�=l�kr��e���|�����l���="������</�}^�h<��a0i
��YZ<�u�*���>/�ϑ.�:�y����¾�3 ��q=>�7����4���%&��xՈ�R0QB�Rƶ�[�ׁE0[ *�Y���{�q���OOoх[�f����=� :ɘ�$S�����e�}X2_���A�4�$d�u<rm�c����\��/��n�ٟZ��׳����h��E!	�eD�/,���,g�E4��ꂉ�=��6���6>�3��})ǫb/r�]&�;�ّ?��N�f�J'6�^�}Sf�^ž�2���Y3%�Mu頇�@�t�/�+�K��cu��w�ٲ�t��vj)o�oT�4�j�Q�քtm���I����;�]�VsG�%���6M�t����˭�[rFq��r����[��Vw.5hĠ޴3v1�����)@�
6�������X�b���R#�N�u��L��S�O��c&XD\�,W��WO�Qw� 1��	~���,��߷;�`=>��ek�KY����i˘{==�`ʞQ�WS��t�d\AZ��ٲ�N>�����s�.�'�r�|x1���d�u.��\���)�S�}=W��d�W�ޭ�ފ-.2�P\c�a�uj�֔=�a�tD�0:�n���^����~U�JW�]gy0����Wc�egDI��:/-�M�R)v���a��� �wQ���w�5K�Oq~bM=�� N���U��y����m�{´����a��3֬Vs�'�xj��{ͤ��(#�S��N}�`R�n�%m�x:꒼2|����J���R���'����p�1�y���X5�{E��=Vob���KI���n��/zΙ�w�p�4��f`/�o.rސ�a��[�u~�V;�PYO���u'�{��[aWE�٪��QnI���h�no��<�ٱ�K:�h��n�=\ *�ؘ�YO�A�4���ұ�y�3N�C��g���mt�pt��>Ү��x��өց�w�M��}}�IjS��6�-��W|�D�K��7{�N=R��J�uwS�Z�*K���g8���5�҈��:��U�Vۮ2� �-�p�e_\���[J����dXe:�;�C)�VZ#���s�) ���G&�����Q��m�J\�Qz��x��������*��ɶ�2�bߡ|�x:N}m��a�g�-�ʼG�#�����n�bR�Cd�z.	����KT�<���Ǣo+]���2e�ʢDpGE�
��M|H�eR�Ws��
��^���g�,9�%%�a�A��*��*�G{/�p[*b#����|��< _5��%zz\�7������-I�
��;: kي��镽�8���
�zJ�g�apu�
���=�~(��e-�、�̾s
rd{(���T��t���D��}Qbь�s��z�C*e�9S�t�!6�
ng<�����f��di*���(9Wj���a�X��W�c�ϨX��Ճ�yi�ûo��uٷ��r�*��+���o����4��9[�h�
5�}��i[A{G[��tS�V'�*ޑ��5}R�T
�uU���/��JCOs�C�Nc��x�>�̣�gw��BJ�����lg�.��_��`xX#����Mm�qunK(��n�xHz�@�l�o���v���"��p3HR�ѷnOb�v�
��Ho�*�����M������-��[J��E�9Y�Wk1S�6�:͜M�����Z�oM���T� ����r�7:���&��tW`
�fk�Y,v��Xe��D\{׊7e&�Z�1�����Sմ6/d���1�:`nj�(`�Uu���2T�tk�a��	3q����,fy-g-�(z;�Z�]f����K�x�}��[��'iW�sʗ)9=:��{,�-�>8�(ҙK�D�{���9v+5��{ڐ�	�E�}�ya��>㺧�ś��.�LYVXN5/���fyĽ��=��om��L��ޭvf?�V?;��K|�٩]9N�ڬ���_�	�(.E?	������t��k��p����*�����r=�v)�x`����<�*�ʩ��7Լ�2��:.	�z� �
�}n��,&P��9�ҝ�vlQ�g���ey����/��pe;���T�u��Z��n�G�������*u�o{���d��Ev+UD��C4��u�Ud}�P����pT�(�֪i%/s�J_W}4��t�7�χ�ڀ��r����wt�ӧ~Nm�00�s�싙�>4E���j\�]�<�>��WF��&PUG���ulE]�ə5AZ2��`�W'�08�	rX�VJK���g�˕�i�;4��W�E��u<��]3`�Y�(�_+��|+�v��)x62�jD�����`u?mz�	��,4p�K5l�ՔUe���W��3p��AY��_��Z�U3�VI�T.yu)FP�.���,/�������q��o:;�����GtY������5жM^����2���Vzx0d؋5�U���8^��۽��q���l:Ө������ܞ@0� Qׁ����}�Q�i���u�g���G��9n���c�Ms(�%�4���>>�*��ʗPj�bB��d]+����av�
�Lz$v����ۓ�(+^&;�*wL�J�K��s1�Ϝ��Ӗ�Wr�C��js�����]Ը��7_�R;���"���W����xj0eWtD��R��ӡ�_��}��ܭy���.�gM9��O"�	�=Z��4ϕK���y�Sō�Ռ�S�Zz���J=4w�d�3ٽ��`��^�]����o�/:���֚�}�T�pz��7�/�Z��I�n�M���Q��3�Uf�r���`��>���E�X]M�u���e^T;�P��E���g���^�ꔹ0�S�����H���(�,J�XV�LtK���0��ǽr{��E&Ϛ��j�׺^S�ߡ�ǇTߧ�ۙ�q��X�����LW�ւ���.�/�B���^;l�f�<"�Q{�%�J���)����1å
32������vS否�U��.�'R+��EN`p���f����wr�9��E�F��Uw �w�l]�0��F姼�J��ur���`�+�ڮ��vp'�v�ɼ�oF6��%����� ���!�q�UC8�b[�ި­�V�3���X���s�i�F���a:NÕ{hL�7���$U4�$eNS�>�dE�w�^�\�]a��N��ۙ�F헮��,��099���,m5��z��z�r"I����L��H���im�������K����djit8S�3=WW\�.E����C�N�:�z������8�Fz6^�j�R�9��z���9�Ld����nw}WN���<����&ʋ��/n�!SǼzE2��kƜ�ǡh�O��S�p)�Ⱦ�Y.Q��ɾ���dk���VY��K�����s:�&S��hp�9Z��'��@�J;�X9��}1H\|�@����
�Wlh��f�A��%Pp��D�r��P5=Y��Q�&�	�}{OKje]�����]̭uD����:&��0D�[�ǆ!wؑ�w�7OQk��&ʶ U���yj�e��D{�}�WQ��V�@ua��U^h��Ѝ���q� �ͺ����K"�R����΃��.:�NG�l��WK�7��U�4X���l֚��f�bKK#��<N싇�n���{G�+������R�6����E��	:�31�ms�X1�50'U��pL�����S
�=J��6[JIӋ�6=Ij�!|�<#*��zNWD]yyT]�����2%��*���{Ћ�6��o��<���_W����u�Z���2��{'����}ph���'L��Nj��ƹ�g{Ԣ�l��*)�A.r�u~�X�JʽU��53+�.J��A�S���&�ߏ�<q�B�t�3t��L��V�e\�V4�`�ʧ�� ,Nj�vP�0T��DLU�\-4�n���ޅ�`��hÔ�k���J������̄��
r����׽:�X�m�s��������4��a
�-Y��w(pь�^��"&yb��軧��y�2>T��Wi�>8�T�#�@�����ƶA��T���%T�7nn�\��<z�*�i�\�����oV�Z6}ё��0�ZGC��a������&z/1"�Ӕ�^]�zD����/��:;�Y9��O\�>�V�:����K�|���<�3:n������˶:A��ۜLwNm�D��e��a´�-A��+�uw`����|��tM`˺w��vtz��/fItd�[���DB��V ��19�x̌BցWeNV����H!,*�k�A�A�F��Jt�L��Ur�Z5]��=�vMՌ��s-8؝r.(m�X炂K��)�o�]q�t�V���|�R�.����x^��wY�Pr��@>����S,Fr,P:�lh:o/>�{�R��p��c�E�?JBΐ^����lc�3�'/K,Ǘ;:��/�Y��E��1�}���h!��j��GQ����� �����}e�Ք���=�g��3�<K,��$^�w�p�or�g�y!��".��ʷ��D��\FklO^�����>c/�I����m�����Ņ靆��*�s\�E=�(d>iΘ�[���)�27��Z�i�<���潭���=W��/{s �Y�p���Ek�u�Of2}��{�|4w1.�y���{�����m��{�^V=.>M)�~��/�جת0k��78��wt��8�o���H{����^����A�L�׉��)��<~�x"�:���H�ne�w�����_��j���H�u�d��0z��P�F�u�ӡ[b\�LK=�����<��kq��e�dn�y�������h�Zu��Q����Ғ�}*�U��/Z�N��s.�����x��/����c���X�+4�ަw2�V�죦x�f��n���F`� #�6�
��[�~���w��ʭiu���{jOۘZ�-M��B�h)];i���;����q�0�T�Z-�룾��6�iq0��mv��:m�
��*-)���%�6,xuyp�Zu����kӅ׷>��p(;e��]���v��C�z�!��{���t9J�T\�`�5�f�N�
���#�s9���)}��f�s���p��n�y�����@��]"�A�4���9nz������u<���7�"V./��;��kL�e��mllȜY���25�,���r��ѿ{��������7c�J�M�Im�����|a�ê���g�	�����T(י���u��,#nw��0�9^�Y{����f:%��Pw0��0-#&(6e�Ƅ �Z��$8yjT��)�M�y�}�����=�5�g29�B��~�'���ZY�^��lxN��C�l#��)�e�c�%�y��r��
��owX�:�D����c��NXgk>q�TĠ�p�GE�ȷ���Q��)	A�1UF�_{���{G��}�%V�J���N��r�Β��mS82f�[��9��>�߄��l�j���v��%�C�f�@��<�]US�Yd��^��ق�yى�ݝ�Pc��
4�e�eZ���e��feR;�V���Y4���5ν�ã1X�r���1r�26�k��'z����Jȇ8���q�]��\�N��O�6U�-���#��z���YH?���\�
�T�i/_P0\��V<��\M�YL¥5��]�kS]؇.]q�r#S��jsڗ��Ru)ws���:���#�9R�a�7Vٵ�ٽ�)z��$h^�-
ܬ��7�l���|ݕ��\-�i���
d�o�Ǚ��Ȭ� ����hJŌ�L5 �3�ʅ� �!�ի0.Y�^|x�VZ��1Z�x�_v��Xw���C{ ��s-LJ��	VHvd�w�����mu7Ŝ�u�Rt�YK���ǽ��t�u
�s*���[�ּ���P9Mc�H��<���n�$r�`��jm����n��ub��ٌ�;�Y�~�w��gQ7;���̔���΄�R����h�Y&f�BΤ�2����t>���*�pJ�-J\l<�&�mҦcۀ$�"���\_,��-��M��w*mz���Iw�Y�P5�D3�Ү��jn�v��4n�*�И�G�����;�;~$�0��Cl*d&u29%j��0s��[;�v������Y�on��eSr; WLmm!�V8�������yml?6�t1��6u }î��ZLM÷@f'm�?aK�N\)�Ĩ���q�]D�9���|iKN�9�H!GaWy|(�:�v#��0}� l�,�t
}D��Q�}N�^��ye��F�v��`N��V:���D�v�d�����ԫn���'f�eر�3K_ls�F�n���D[�FÍq�W��{�.��y���]cv��2�VQ���]��ɹ΍�J��Ä�{�D�Ek�f���ީ���(S�u�})SM���-c��
l��ޮ��3�4���u�%4�_b���:�F`Ůd�a�Q�n؊�d�ڢ��MVaV�М�.�+��ǖ�
�{0_�����{t�6���Ж�c��G	;���9��Ԟ��� D2h]�:�}�{����a	Í���M�,[C���*Wv3�A>�><;z&�{�mѓC�"��ǈ���ffӴ�)��zsi�$y�A�fn�۝���mv��}��v��n�*�쌅��fL�v�.�ԭ���AS�`��$8 ���:�P���o��^�u�ўnJQj4�L��A��';eG��ԙɛ{Eo>P�����*���k��{��}=u�=}L����q	<W&Ͱ%&.unjZ��P����:Fh�qn����'6^rD�6�RV冀y������E��-�ָ�*��L+r[��k�B!*Ɏ�X��;��R��ƹ�$�4]ðw\wܶ�]Λ̈́�#1��ق���[rư!�[6� �`����wf�
�_+��b�i�(�zK�N� ->٪�t� _7���i�s���\�Vb6�P�-a���K���Ь�K��&-��Y���#b�8�d��."%\ʘ�hT���F5
�c2�[k�"�9�6����R�و�k*Ua�7,1�[��Uˎ2��qQrٌQq�D�R�ٖ�(�R�X7�J8Zfa�ʢ�&+**�0qX��
E���Z�m1�
-�fe
���J�\ɕ�����Ƹ��2�l�U
\�iS2�1kX��K����1Z�L�堉TkE���(ʨ[f%�9KҕkF\��b�����\��,Z�D+�D�q�)��Ķ�QA�J�UPh��R�T�(Ҷ6�m)Z"�6��r��2�e*�m1�V%�q2��R�d�̨��()X�3-*�(��D��҅H�ijc
��(�֥m�Y�fR��q�r�S#b"�q,Uĸ*��XV6Ѩ\�*�R�f	��U-���Q�e��iX�.9���ư��1�ܶ�ʣPEq+Q��0ŋU��� �-��@f��{��b�E�	1m;�9�{ow�;�X�3L�fP�y'ϸ��,d�$.��s1��0Y�1l�ʏ����~��X?>Y�m�dF��o�/:�����X��'�~��{�}�}��E�9ɾ6�T��پ����}G�i!���/�եc.<�C�qV����i��z�6ojOzf��yۼ�	Zi��>Z��M)������K���b���a��Lt����l.��k���e���t���UҮ���*�Y�k�
�3 �-���7����+AA����gUZ��z=~^oQ��Wz9wlLQ� z��C`�&�Ʀ3��U�F_,I�RR8��׺ϥ>��\M@�-�}h<�|R��)	�NS�*m�c��p*-�z�nzzzuc��We�U�[��*6+E�ĺ l3l��J�,g�E4�낳�(,������SG�kܽ�D/�^F�c�M2��vhV|8S�3��^�~�#9�YB{{��$��Z�7Z+��~��觎zy1�,6`�.�`����q��o�惞\�G��r�v�Hv||�i��)���-f�~�n��r�Ɋ:���_LGw�z��#��^s���c��XՏ�P�9i�^����lb�q��eG�&̣6��{y\�{J�[��C�Է����^K��5sv�u�U}o�Lذb�WS��p�uJķ$ʲfn	~�����-�j�j͙���{���WlT���o}�8?>A��]TY2��D�FS��c��"΢�͠t<k�w��z�[�� {A�Q��D�k�b�{����4�Ի�����G4=��K��,
t?}��x�w_�U�D��G�O����p����i��g۾dܷhI�%��xb��v'�Xf�������'^�lٮ���ϗ�L��ԗ��g66��uKRI�h�
a0���&�����_��耫�/*�+�<�3�P�%����/%h�P��=�D�>>5+[̮���e^�d,J'�bd禦;���Æ�3	��\��6ώ�[ԛ�m���X�fKa?vd�zxT�W��jfW��p�Ud���p�zd�t���Cb�޽k �42���z�`+"��FU=\  �bsQe?��ZVp�=�۩/�1��	J:�.U���j4����:q�Q��3x6=�=徺M����! �oԧ9ܩ����/x�`���4�����՛��IJ+d���i+sVl�Ϧ��"�zvn��\h�ˣ��'IG��Uq�����^�&���~^�8�7|Ld{�1�Q��(�W-�W���xf��ń�70u,WJ�u�uA,��2��if��)��pt �	^.�N&Y��.�G{����"�e;��_4�H�vF��j|�c[ �h� ΜX\u�#��{9�o���g_.&P�&��a,��eH�m]w���h��yׇ<�Io7�2fx�;�_�
7��5�聙��ӿ��d�Fa��꩙]��,Y��
�͙[Z��ţ�%y���~���*>�,U�pT�ӛo�Q(5�E�F2��>�z�A����7���������z��F���п�Y�V����]��k���q�#9�X�x.�Mxr�s��3����#(c˂�L��ՒkX<O}n�E�AʻW���jѪ���R4ϣ�p��ο[�2�_IV�0A��ب�.���!�տRRt��/�>�a$O������^��ڛ����C['�yF�RΖ��\FklO^���.�eȳ�Q��Lv�z��O��H��߶���hlS%01�0��P~�<k�N���S6N�����3�|=�=���Ag-�({��E*�)W���d�ޗ��,Z�\l^���&��ϻ��Y��~�lݩ��0�\��ұ#�γW��g(�GPfR/+��#Jj7]��WP�%� ���]1ynI��W�j�@;BR��p�q.Q�vA�a[��-�oo�{nR�԰Ғ�y��I�	�`���N;��qa�;J�+�q�ba|B���!b�ާ��~T/f��g:�e�}��Y�՘_��xR�dŕe��JjdּM�}U�����\$+�^�+��2�ל�kٱ��v�O_u�2�>>���]羽���,>����G�G�iR��X����xv���H|��V]�ln窭��e����o/��Dp_ʻ�g�<�k�WC�����|��
�\����N��0Óp�:��w3^�^y�7�І�|ؿt/m�H���y�y��@|6Ki]��\�`�5�f�N�
��"52�N
��J���ޞ��u�J}�
�4��=dJ@�M�i���r��ϡ����x"-�z����� ����<�DUS T��F�����ǭ�h�7��dɷxt�,�߲��Լ�]��{���;r)���u�w�h��5��M�8�b������=!��|_��܌�k��Iy�;��<=H����O A (���������R̞�6��b~y�E�^,��E�s��~C�Q�k�-�� rW�[�+EX��j$>�n�\�����G�����]Jh�����/����16��3��g�m��Q�����:�]�S�U�޷���f�m��/D�1�&_b�)��o8�Y]����qO��%T��өv��hmd��b�{�~A�X��ն|fNx��o>�eU��ہf�	ﻐ�2��Q%T�_9��8C>�q�I�9����s���Sՙ���8vWX��b��^��<�G��t�OV�J��:�뽯l��i{S�'���h��u3����ub���^��Ik��yi�GE�ңZ��פ'~ۛ�[|��"�&����^�ϫ��u+��3�Փqұ�TN���;������{Fbi�ђ��;U�٦�T�^��=Љ��fq����0&:%~3*�6fi�W��Q��ԓ[�����Z*V0�P����2�m���8#0=9�����O�U^�h8�����v"�Z�M�|r}w�����.��,��|�V�d����ު�LW�X��ʻ��}����vr�`���Y�K�$�{���p ��C`�=��N�=�M.��a|}|y��r�,�c�A�%C
�l�x�Z��H�)��Ӓ������ɶD��'�p�,y�2��oZo�x�nv����1>�q��U�p���1�������v�+?�^ѥ"�N��GV���E�.�+)S\^��۸eA�K����S���~H����ەL#���i�-�2�Z��]��ѧ��&*Gs
=�_	�&�6&D��'t7��K��_���}��c�H059A|uA����5��o��Y+U+���c=�.��舵<��=O��{�t�_L�5SHЫ)к'��uu�ߩmZ�|�S[�ڷy&���K���Z����!�觎zy1�S�L� �z���c잻���o:r��S�
�||�i���ek�׍8_��.a���A�'��y�ᄮ�ŵ$YMjnxO9�3p_������^EЮ��&����8�GG�>�&S��V�r�>��҉j��g�ǆݛ{kt��Qnv�Y�=�J:1��v���C=�pwK$�p���kv��C��)�ը.����;v�|΀x:�>�ז�ī�eȸmi��sv�n�T̆yz)Е8�	-����.�K7�tN��k�ie�/*��[�5�<�Z��>~��GE'�L�C�/T�Z��Z�T�<"��w�
������aC���@T�w�pOyc��Lv{�d4��̨<���۬����Obd禦;���tA��G(c�w�j,�q�B^Ld����|F��o0U��Gt���Z��M�Vk�ڂ��x(�MtF��p�������n
��kr;�&��#���oe�z 7INщT�A��\���#�/y��'��y��'�3�we����p'�̔/O
���U��SS2���d��A�Ub\w�=ts���v:{�{Fxث
͖�|��C��0���'ݏG�勇�s����UƑ���/IO��k�<+Y�Y�r�~�E�2�ۋ�Yn��`�	A����'�iη��䙋|�d�z�S�3�Y-v��)uG<�&
Qn��7�B���V��6��=��O/d�����/��}�E�V���|.qʙdr�����j��I����t������^�>M*܊c'��7�;�VNyV3�{޷c��G�0�=�+|��#.;���U��{�J�l
��=>�wz�ӣ��Y9瑘`������wa�Up;��fL�~�ȥ=�B5f��^�0�v�g>�,U�pT٧=n]��2,Z2�p�A`�y�١��Ǽ�!���5Ҟ#B���Un�k��n���۵��K�e�Ve�Vg����������FPʩ�/�U�T�j��IuK��4�77�;��)ょ��1�R:b�J��]a�W�v����Ȳ�08�՚�I2h�͓�2�>�V.��ү#�����R]�Vn� �Գw f��S�ۀ���E_3B�Kƥ�xz�=i^��J8��[d�R����ݏ�� �೽۬����޾}mg���5�Cʗ��Zd�ʷ�eQ�R�T�]N��}�0��5�h+�zu%�*sqx�F����C�G|+2��Q*��CcE�UNU�'>���B���Mܮ&Kz�P�S�wӊ�-�>��gÏg�h�8�/��B��^o(G-��O�=~/:����=W��gq�Z�ű���1�>+qC�j���9����M�[�P�w��ʺ����M�����q�96-/!x�0�}��Y1�e�F�>v���X�����iL��^Z$#�K��uw图�ܽ윟&�½*5����;���z{���Ӥ�r���|��w���g�{��mK{��K��5����\����~�zk="�׵Y9A޿"<�j�ΣH��$�%t�D������
����C�z�ڜ`�;��&���U/.*��|t\kw<�꾎f���'��}*�֊_\��ňK�0�&�S�pw���kӅ׷&c=C����L�8�~bWǬ�
��!ϮEw��>f���f��E�9������J�K'c��h�]�T�;o�xQ,�6��W�_rс"�r�޴��Kԩ��a*�V�gTU�����6��q��M����ѧ|��R�0� �o����EEJ�]�Út�iL���g�Q�غ�,Y�lk@J�z7��-�\�757�Ku�^{yI���H��Ս ��<5���ۂ7އ˰�_Vm9�����5!�>4T T�f��<L��=l<��b.�d���}t��]N�Ok�7�g���T{�Pq���y�3�O'�
lСJ������+%����z��=�#1�H<�X�y�Y��ל)xo��!�q\����(�#��*7]�k3�.���;�>R�*�UM��>����9�D�CO�'��NU���K�5LHA�g�U���Cx{=��S~�4��B��UYbEx��-��r�}�2�2(��P9a�������^g*ԩ�����}1-��@�:�0�/�(���8z���3\T}����=}�b[�bXi�@��=�l-���pe
�2�� ��g��c{m2;�%$��-j��>|��fRo��~kj��}`Ҙ�|�}~��:A^$�V��yP���Q/h״�sT��{iY����:���2���o��Ӆ���i!��L��V����̿��{�[n�Nz���m�O�e����Y0���=2 }�>��J�T�e3���2_f��(q<���yk����V�{+w��a"(ܵ,�y���o"���lL�MoQ��Q���+Ve����5]Q���2��ʗ(wN�Y��FS[@Z��_=�1�Y�烹��ë2��*`���[�Z��Ҙ|<�NzEo�E��Cxn�?G+:�7���S�I��Ͼ�Z!,i;�:���t�/��e�q��*���f�{b�=ex��q��ʳ,J�ٹZ*���Qg��`|bKG��l �d6=�
�q��&ץZ+;���5��?bL����4�U�6O��������yJ$SJBFT�u<nbU�4�;��Z��D����Ѩ}zG�4�K��aK���D5n`jr����;�&	}���Ni�ZK��4��1��]�1輭�TfN7��eI:Aߖ̉��jt�4�#�l\S;&�_l��tk�>i��\���t�Z���~��觎z�y1�S��`Ki�ެ��]�s͍�6x�%
���Uo�*����qL�~��M?Ct��S�0�z{ ���[b;�c�ҽ���G�����Z��\1e�Mv��O��:j*|"U���*V�e�Э���6{�N����0l�$�K!����VK�C=�pgtD��Q{謽N� ���(��7L����M���)���hi�n޻W΍��'oC�����z�#l�B�\nR��YÄ�wM����L�aԜ\²���3/����]_S�i��*���2S�ps�-Cm����J�c�o�܄m,�d#��DE�s{����}nl��x���.ps+5�*�B*����h�q���d6����5����
�s�z���H0IF!�{���wMj�Ҭ'���4�k�gm�0Ѓ�������#lw,��]m�\�ʜhK�ݷ������>v7��MRt�3w���1��m�]��I���z�VE�2�/9�	�mZ���{T��fK��:aDĤJﳔ�S)�uՕ�q8[��u���/���)�ce�]*uђ���^҅e*�ϮV[��>v��dު��^�V�K�� �6:.���e��	��2��:v+�e�YT�1��������b_Sp\�`�����I⣊e��Gf��T�2���uX������� �-�4��I�u1`��f�g.����Ϝ���eawȹC~�(�˲:���G�p���}��<n����5�q�F�LE�'uA��7lY)q��B�-����{.�U�[w�v�i��,R��1bӫ"��͜��f�;}������a页O��>��I[�x@ް�u�WR����up���>��l�[�c����b���@W8r���U8f��GT�N��W�s|k�k�'���=�Ǩ�����$W3{�m��/�hs\D@55�\��x��^�A���f�Zi�J�7�0�>��-�2�Ed�O�-͹g��ԩaGǺ���sҎN��c#`0�,��F\ݷ�Ӭ
�6�(+�nїr���͜R*�k�����\�nW��l��^HK���Mr��Oh�M�9V�js�p� TH�[�[��Q�{OV���.9�u��Yk:Y�$���Y�Wo��6L��I ��9�'cp7�4T�ͮ�����<QA3����*.��[cT������>u����y����ĥ�,�	�\�!vBٔ����� �FwW@��j�U�J�{���X��Ю�"���r;8X�����M�Canvi��SEõ���;��W���.�]���c�S�uȾV
ǫzds�BM�+��t�˺6�Y�ڴ됕�ˍ`���]�bn�H�j9�8�n�����ֻ0mG���:��>��X�u�;��晥�J-ڱ�vJ���,��Yq0��e�'���w(���2�d�hZ�hhN��"�͗;���&BXGխ5o�U��Dӽ��e��^�z�e�Q��J�C`ŭ���8��e͖V����@	:�]�
�'e��pդo%���;n$��ˡ�;���ˉg�w�+��ɼ����E���ڻ�8�«�]z�%� e[�ocH������X�(7�1wn�"�?���߷���b,�UҰQT[ZK�ơs.
��ZfQ�-Q��DT�,k`�ê�ږ,�ֱ�p�\�C1�a�2U)KJU�\���&YVR�ҫl�-R����Lfe���*-*Ң!Ym1���5��m��[�.Q�Z�c�V�F�8�\VcQVcL�F\����-
�n&T-�E+R�J[m��ԥkKP�K`�̸�Ze*��FŨ���+��i�Dq�cC-�Ekj-UƸfdQAq-�˕+��kLs��r�T�Q�)�������f4ʪ�mj�T��2Ե���2U���Z-��i���Z(4s��-ƴ��cL�cAĕ�pl�Ɗ���Z"�\B�T�[X�(2��iD�j6��l%������,+����1m(R�\V�4��d����-�iY\���9)Ls.e�im1.-X�R����TE�m�E���emr�"e����[3.E+L����'Q�n3���!㖑���-��I�����s�6��Q��g
�șc�=ެ�>栙2��}�rd:(���E�4m���}W ���_w���u�'�mY/-��p_H������e{;��2L�Wy�s�V��sh��� �uS�l �X_<�S��}G�cQW���;�Vx��e<�\�F�Rsk�:����a����"��/�
��/*�;��C�����\ziR`��2Y��b�+���W�]^�d=A�>	�L����q��F�D^��J�!iu˳;2b�>]�,��'j�'!��(:[|*Qۮ�����|g����ˮw�o��LIk>��iOcѷ�V,YK�IX�1r�]N`*��r���� 2�ؘ�g|=G՝4�w����{+e	�i��=���5ZU�}B�U��ϑ�qp+-к��!r�Hۣ�L�N����_a2�����S������Y�uG<�&	��&��)x{�����wi�~�*-)�ۢ�&}OE�6r":ȫD�Wi��s�D�ؑ�r��xF���J	�w/;���z+Х����'(o�}S��29���vI��s��-��5݁?��
�$�7��:TL�y�ʔ�2����
�N��5.tn9܁k�'�)76�:}ݡ�o˹�R��:��x�ɏ��/�u^�B��:���9��V�e-�]�+�˞��&�����> v�?��ZEʻX-�W�j�ʻ����R�
��I�N�w����̷�D,{(��t�i�5<�?Ws�#0�Ifo^\��ff��h���=�U��l*j��f�،��b�s�����~�%��h����^u��J����ϟ��1��i�4/���,����ڨ���4�eԿtak�����l��;�r�{��c�`���pR�WQ�$�kīw�,���'�8^!-��?z&}d2�W_�˝��DL�x x%�@�*ޑ�`�T���]E]W�>���aeJ�~Ovc����n�
�"���Lw]����;�ةe��*ޓ���C��Lz����[ǚ2N�!7��{'�q�C��K��,����Y�i:�]{2Pʇ��&�~|��U���Ҩ[�8.��q~�APy֨/��xg�w�x{&��(z;�K�r�{I�X��
�����7�R�(�6�j�Z�q`�i�u���u�d��x]-ʸє˨�g���;��t�y!^���^�gqڬ�xR�dŔ���*je׈S=��6R���w47J^l�>�M;w��v�Y��o~��M��'�ҡ������&N���w���j^�y$2���ebÑ�V�O%v,��-�7����bgq�@�Ȧ����&�;�`�]����^���N����2w]��c�>oϳw���e�r��#��������%��y9A޿"<�j�ΣS��g����?eYnx��m�6�Ϯ�
1��v������_[S�wxg�=6��w;;E��'����|�1�����Ѽ6Uޣ2��]�u�	_S�0ßM� �:��qs5�.��v��T�V�1�a�:�)��p�>���Y�/��!˻�3�v+��X��x��a��DyS��r��Ryڏ�����u��V�i*�=d:T	���ƐyTҧ�L��
%xn�q�ɾ�fN�փ���3�>�@�UP�R]�O(*=l<��&L��R@�g�\��<���bb���D�������4K�[�gΓ[�i��p_�f���hW�o+fi�:��g&O�f������y�;�����C�2�(7*y �^�?Z���������#-�C����{z�v���H}:�9TGIy?P�>.Q�i�+֍�+��×pf�~�E��Z�S�.�1S
��yT�د-��r�}�2�*K���:�hԥ�����%
����'SÊ�U�Prk��o>���i8ϐk��\�g1v8��y�c�@iH�Vm�R�؏���*�Z��F}�L�r,M�}K@;c诵6J�F�/�lY���-���:�6�����]���2���Rz��Ӥ��[���]foy��6�}}��=R� 4/�%�>�FϦ�*C����:���;(��`�M�^��g�;Ѝxܝ����o�j|�c�X{:���=�������R�c��߬�ԅ�Y3�+Qė�er1&����sj��]��[뻭�x�V�ؘ�{^�t��
�g��Ş"�=Ƿ�]���mO��<�0����M�ټ�~�.^���S�����I@m6_e��6�^�m�t͢]�cT����coo��\T�]p�W`JP��[�����SJa�b���T�����#{��E;��Dv�~j�!>~�ȋ��]��%��jr��i�-���y(6��zM�V�ka�d�2w���Cw�֊����%�K�Z=�
�`� ]�!�q�]Z����]0/�\��v�9�)������W�T�ʴ0�!��A�x=Q �!#�M���2.�G�Y��'���V#>�9c����4�Iv8�+���!�p�����w;ח�Ȃb���̯F�� ��'���A^�ND]'嬡����=R�~��|١Hh��q%w<������j�I<o��R�͔�){��֜5a�7Z�D���*r���Ԍ�'�P(���sMāM����r��m>{p��|l�l��4lt���U�jr���6jŅ�B*w^�gx�Q\�j`0�^��Y�E�����,nqҚ/!N���YG�����|��-�׵-W
T�?y	���|��sh�ͣ~�l��;���� ��IB��_���H��gyt�+�.���q��uOg�>r��ٍ�Wz6<Ȋ	pG����z��?1��}p~|�9�x1��QS���^a��<9l��N������evH�k� ���{�K�V�ؿ���g�� �
���Wt�x�{�=�kZI�7LN��ߩ��A}=�F�;v�� KT�x���eK$!�kgU���^��|�/��
�o�,'i�F@r� oK�媙�GƟQ�2XG�̚��G�����u��q��j���o�g�w���@��<#�zG?m�eQӵ�T 3/Mٞ�9�"@��J�Ȗ��OƲ��J��=\�ס�Q�_=������T��mLOw0{0/�)�Ϸ����4A�Bl��9�]����p*~��C�o�J��]��q�N���Zlvl�O/�&� �����F�*!K�+�R债��[���z�@ ����C�H9�����8k�)�Ve��G��[�G��z��6��|߷�����l�%� źs�l��YDku�B�"�r�'M6�w3�S�7�n]�fK�e�=��J�����aV�z/��������5��f�{r��7��3_k��>�\��9s��H^�Vy�ܼFB�U����qp+-С�Ia�`Ҹ�t��=&s�����H��[d�MPR.vT�7&�Q��9S.��x���a
�.i�b���!G��Gt�V��W���
�2�z�;�.�A��Wi�>8�H�ú��r�Ƿ���fK��퓼��%Q>Ċ���Ү�O5�X��v���d�����è�X��\�sk/�j��J}�4O��샇,��P��d���'�l�������Ny�S^��5�����} �}��W)�̩�)�\
��B�ل���#9t%�R�{S�eO,��n��RԠM�a��I�����a�iZ{F��2��i���̐��[�Ġ��j����A�����{cj����i�x�X�~�D��U";C*e�Je]F��Y�_�ۿh�;k���J�)�w���M,W���<��dG/>� 9E���	��ͻ��{g�E��G�\e9A���X����}��[:)>�O����W�Ց ��dx^d*�� �̥d����f���Zav�,Z���^����]S,��Z��]�
�[��Ւ�u��r��w�k�2a��3��������]2�Xm`:4�f �s�!q[��us�_ZYǮ��¹H�*J<S�?<v^��N2�ZW;ǦT(>�Ը䗮@ŏx�k!�Y�2������{��O�*�r�\�E�R�OLҀ+��?o#�]�g�AgLB��\0`�u�~�x^����w�x{&���/ܰQ���&�&xn<n+z�z�#y	�>�I�L~-b5�����R�c���SAx9M�^��)y����\B���6����v1o���U�xR]옲���Ձ�n�t@��S��W���Į��eW����МZ�����EOMezE;�rr��~Dx*z-B:)w�t}��-om8�$�K�J2�J�t(�j��Xd�p�ڜ`�;��&�����{e�yқ|�8�N����G	GE�Wz��7\)}r��W[���0��"Aθ�� "�Ɠ��� ��&{b�,Ss��x/���a�xHr��K$W{�l�k��3��z]���z�t�4G�o3|�0�RpT�(�ֻ��Ǭ�J���ˢ�X�T�k<�^��h��݇��2�{��/~�9�����5~�����]2'Y��ɑ�Dk�x=<�7޵�3��ޒV�ǽ}�樇���1���wƁx���>7���ݨ�6[�71��:Xh��,���H���nY�Ѵ)�I�P�#��R����ۡ=�h�1Y9�\ w���[|����O�]*;��&K]�����SD����r���$�<�˥}^ðe���(w�A����M�o��P�\�P�Z��F�}��k�X�w���y��'�uz#��`��Y���~�^f�������������ܞ@0�G��k[^�go;����j��UYpŔ�>=�.B�u�s*9�B��~'��6=Z ɼ��AR�x�A�z�&$<;#�C�l.��jS�������<d���J��
��=���F_��ufk]����v��������|fu�X.�b�U�{s���!��q���Z�BT� �F�hm9�*��� �e���߄��l�V�/?�*�>Lp�u�`�FǷ�O$߼�)=\¿WE����"}0_=PI�'��{:�uV����P�V��WW�&/b�M�O	��JeB��G��o,��xF`��i�|/��m$zb�̾�W�N�\}�g�ft�,�N�׍�<���s>��J�Uv�C�ka�{lN�����`zs�(+v�=��z�ʾ��U��Oy�%O�^b%�\j#���\�FS���z8����P*��i��+�u�v��3�(��4U=q�)�wq����n���k�x�)��a;�ˊ�4�n&�Wmgx��2_f�����qr��> �j]'Dr9Y�Q�X:VrtN�o�}dW���68�M���\*��#�kZ��,L�K9l���ΐ�g"�i�<����l�LW���U�e�z2�Z=)�����m�ٜ���6���a0���{bz^�c��
����d��R��JEh�O͎>�i����M�<$}ǟc���2:��~ڭ�����<ҝ}��0���,��j� ����p^��7VQ�r�K^��9^�{�
+h�ʊ)��R�A^�ӑI�k(<�`�.�+�F��B�2vo42�4�=�s��[@�r������54����-W
s�b=��O&3�W�g�w���mk�ך����=�
�Q X����
�pT��3�QL�~���B��V�.P}����Ś����N�m���Є����S�t��UWlWYT)��@�7�8�x1И\��o\��u��{u����:p4�F7aS�SL�(�+� ��{��J��n����z�;s�A7�0�������ʗn��`W�',x��%O+��,.�<W��vQ��W�g�M�`�#<�.���q[�Ī�CÝ�UV��j2�W��@[��צ�6k���z���E]�؁g��!b]�1�Bi'������������v9C`&Gmf�Di
�ռ�;r�%��������:G^=�{-����z�' �y&9`��3�X�Vu���a]���`��F	�^�9�9��r��np���'%[ ��f��Q��VV��߰�|�]�k�����9�Dz��%1Nbߤf�3�6��]p���G]%x]�=+�Wy%pXu������(9G�Sؙ4e{��;���a��s�cG\t0��:f]��%�%C��̔<��T��U���ڳ׺��S���=���q������_WE����Q��+�|�`.�0���kތG^*���m���^ �}l<j,�N\�p��l���d�ǓX�i*I�8͵b��<���wۨ�Z�Dz-�r\7)���{loы�9P�ʭ#Ƈ����/0�ä��~u�}>�u锔��%S�pM�N�"���A�S�]�υ�1:Aڽ��3lgn�/�#���C𾠨�"���U���'(o�}S��2sUc�^��AO#�/μ��3#;�m����SB��L#��[�{����+~�G���F�J�|�˸��tFs��{KF��w�kF����|��T�*ת��o����$���$ I?�IO�@�$����$�$$�	'�!$ I?܄��$�$$�	'��IO�!$ I?�BH@��B��$�	%!$ I=IO�BH@��B����$�����$�$$�	'�!$ I>!$ I?�b��L�����*� � ����{ϻ �����Ϧ|�(�T��
� �PP P R�� @ R�)&�%HC��!@U�TR�*D�UPB���*DDU6�!��*��JR�QU)"�R�UBJ�(*JRD�!T�R�IP��*R�B��V�*A� � �������D )��R�L`T�ʔUf�A������*"*�� �huB�#$�͡�X�(ڱ(�6��ֲ �M�l�k maY֪FA*�JT v�n�  ���(�  �@P   ���� �R�$�jP��CkhƭY���RP�U�(kAW  ��hc�UL��(�a�j��`e#f���b2h����PS!Q�U$�d�6�  �t�ҀBR�����m�VaYP,f��X�"�� ��eH�U
� �+�*�Qk�P5c�0�b��P�X�Z�!F�UI$)$�  r�&� �`d��-X5)l��[0��E��l�
CX[R$B���  ;�E(�ą"H����EY�J����J�0�@�U@�p  �R]0�m�`�ƅ���i�khY3l*�*"1D � ��P�XҠAV�рmF�Rֲd���(ضl�}�� ����*RSQ��@h b  ���*PѦ�L��i��&�# �D�M0�i1=%6jjl��L�=O'��S�A*�=F��M4� CF	�i���4MJyOj����3P  �� $�IU*i�&10 Ѝ}m�^�j�-�۱�S�H�%�a��D�#~�AB���R�ܪ�(u��"���U
�� (HH���� � ��?�ϩ"����AB���
�h�*�Y� �
����t�mf��xz7�6�� ���:K���A1�i��ܟ�*�1	p��2�-i�):�,�ULތ��i�׉�*fk���NV,�u�,��|�)LC��K�nDt��nS��
p�B����5��'*��݇ɪCdT,�ff��a$1ɶ��zN���%�a�0GƵ ReU�c	57���@Qm��v���N�ͤ�f�dt6+�n�s@��CGS�"���e�y���gn(8u�51C��U�+�v�V�z�v��
2M?��V�7��٦i��V�c�.�-yX)PQ<�*����0,z���u0$	����X^�p�wX�} �b�]����7ZHg%�ѥ���	���S��	�]CIP�h�Zt5:5�S���s���3���yZ��1��*����� 2�Ө�D#fe����j<��vȬUI�1������KCq<�V�������+E��P�4I"���喯u7�t�Ъ"d�3Qw��@O��8�9�ƶ�\�Y5e��f$ �Ykw��	h�1����2���Di�J��'�H�#L6�Z$)b�
�i{��p5���;�(n�!�zg�܊2)�+LԹ��hY��F����o���v�.iV�ʗ���a̽�njӵ��Y��,�V�H�x�q���aw)M�ˇb��Xh�ݼu2�hS]�n��:�Jճ\�v�h���ޠJM];'s4G훬w.�\���P�,��ǷX�sLr�)��)ŕ�n�`��+wK������D,�l�5���Bx�6�V<���m� x+EbZt���N��_+u�'�ȧy@���n����+��gf��j6�7C� �[���O2�OZV���/��ܗ*����r<��N�tw�qk���ˮAQY��DqK�Q��0m�Y�q�v�^YB��yE����V!�=�Ph\U% �LVh�q����R�f�
�.=m�k]wÃ�^L��ǲ�iF��wO,:n��tp�w3ct�ʵt2�U�m�W!_�
� ��Vr��	FL{L;�MM��=ݭ4��^�!%�������*�wL�p[����1{�q�л�i�x�۰�f���͡�3�ѯ&Hj��@�+E�)�®\��*�u �	F霢5n\8ΉkA��7mm(�2���ɦr�K �Y�S[J��&�7u�T�ܭݨ�CV`�{���H���&l����,����W��4��Pr<�	�l�/&e�b֙ˣ�Vd�S�Y�J0�V�˲�Z�R�Z����x��
�Ҏ�|�ҍ�}co2�����96]�`j�H����%�����O�w���i��a���z�*Aڬ���m��z.CJ�V��"�ce���KtYY��+�}oj�m*�j9f���˫d����Te�h��予MM@���G+&=�.��t��;��	K#��[LI��6F���z�vΖL2^*�K0l��wnѽ�4b�$�[n��M]nf@k^ە!�MP��jcz�+u� �xD��k&�w�ޅvwT y�b����E.j�,D���7�>�4bP*��+����Y���-@�� oY�X��[x��gq|>��2+j��9���%6����h���f��⢅�f�,����� 6��Ǫ���s,���D�-��h�t��k̸\D���.^b�]̩ywl��J��wM±f�.���Nd���]��`�H��u����!5�-z������K4͐���J@C[uR�
=#Qb�D��d�bQAح<�ъ��5\��,�s$S
����U�f#��
�t��,Hm�q�![���zYg���l_>��PU�L),c��3[������hF-7Se���nQ]-�X潔�GM��]f��k�B��yZ��vs�s��eұ��\*�驣%[�2	���!KF��u�T^�=W]n��O<�Yk�I��5эm�=���}yL�zr���EE���f��+$�)b)�C0օ�w���1ѿ��vJ�WM�M��P��ւ�+w��89-
g�(��w�n��٣n^�5�>)��ƻ�towQ��,I��5!��ڴ�1!G]Cjm���D/�n�A+S�d�Uۊ�pUEtB��rD�V��W2\�tDq��Y$�5v�ZӏK"�d��R�LQ�h��;�&�ON;QF�1Eʶ�����v�t��1�6��7ib�ܺ�2���P^��(�O]�gW܊�l%o����̤�a�	�LQ�U�5z��D����1f�Q�A�e^Deչ[N���u�K�')kģ�tk	�@#�:�x�`w�!/ b��[kf�Wj�hC0�h�+k
y�f,j�l��%�#qJ7(�0ф	!#�e�f�e�8���^�54mMn�5��z0�� �8Xe�5����*���-ٵx�$�^�,��23���y��g2:(4p]�^�5U��Be^f!y�<ȖԨ��6,��I9��q��L�lQ���8n[��� Cu�C&H�+`���J��z)U�b�6�ɹ�Yʿ�j:s$���P�>u��+Ce������ܗ�� �f����ḿ=�e�IH�|��r�f�׬���qk(0�#�+ot�^K;�&-4N8�J�^�V%����m;t�Rʲ[�[��u��g`n�ڕ�X�ʺp��2R��V` V�n�ᬰ���S<�W��Pe␥n�8���N���5�6�#X ���	�e+0g)h9]�$�Hy��7`T�b����C�!#�J���zL�B���]���1edj��%�p���tV��X��J�$�kh�#���),�r�
m�ĩ�
��l�0��wrc��T��G�.��dv�Q<ne9��[[�PDmR�2�����[���H�&$:U2զ��ݔ�I('`�*�8#�:�7����K`V�d�
�l�-�9�Ѵ�I�.������b�1��n��)4|�/�I"hKe0kjR��eaJ�K��pO������x���U&�5N�n��R��]wjzC�|����:�Kz�DG�lh<Oq�t��P��8I�N�u��fe�����Z�HϞ؅��ZzDZ&�ݦՄv��Y� ^�ذL�*�-COdh�0N%�5:Ճkl�X�j�l�J��&$*u���1�@�����wG�ٱզ�Z��w+qUO ���舷�CP�Y��F�wؖ�֑�[v�ǧlw"�t���;��	�jq�,�yTt�6��t��ʐ�#�Rl�(��R2��d|S��)Yus]�w��Q�x��R��V	,'��F���;�������r�n]��a�2�3�n�3VFRU�P���l��Z&����I�F�"��[��y��Vƚ(�md�V͕���U����%�1m�l�oor��4�6�--b��˔h-�xYx�1i!n��m]����ucCدh4ZZ(=���6�9Ja*��Қv���{I�ZƵ�U+.������;[z�#iU��e�-K��\J�%ۀ=Ⱦr�[�lT��Ɋ]KT�ʘ�$sn�\�&�c`�z2�	��ݽ	���Ƶ��YZ^ͺh$^-���.	I��n� ��]"o$xt��vikRZV���[R /f-YN��g!�5�h�l���ͫaˆ���Uy{.j]
����+��^M�<�zvc�	�o��j�a\�>YdSs(��f�̰�N����Kn�(�Y���&^�tM���ðSز�y8���Z�譣��W͝�v�Ϧ;#+c��͙f��w74�Xuz-<sseh���R[�7V6�ee��@�n�U�r��˃[�23��5r`M3[N��*kJ���i���4�ܥP���,�F�Z�� 9d��2���-�r/�#+q5�'T�i�ݬ����!ӹG�G2���4N�2���7�R��0̺�[�-E�D���hl�V�:��,�И%�h����D�	�ٺ� ޑ$�HZh"�8MZ�]Y��^SԳ�v�T����iZ#
�7�g�ߎe:��E��:Ά/N ��1�m�J3sZ�-6��,��l����0qu�������S�fe�հ�b��͚�U�ɠ-Y�]�'Mb����A�%a[�՚���h��$�=єޱ���oq�:���4A!��˥@ZN�5ʙ)����"�	�3ue���e��֛�[O>w��sAzo	�-L�H�A����һy��C2����oU�׬��E��I�p��8�a�Aa&��v�Xz���a�9m��'�ܹ�Mf;64M�,� ѹ!��Y7@�F�ʐ��7`���ͽת��BAQ���m��^�Ra���� ,���j;�F�t�m�8#�]�tj4md�/M5Ov��?B2�l�X�F��D��6%���Z��^����j���+����V�
���J�&�W��\�d��w�Q����t�:�o�9����6潙��*�.�ۊ�\���9���ioJ<�m�yqpzc����	�+��LoD�Ծu�d�ڝy�(m����jP�e���IsBN�`&��<����ot\8a�(��W�y��ڛϰj<u;��;y X��(��֋�M��cG0GN����;Ú�k�2:��%6���(��X�ma9;8ڮZ���-� v��0�k����;;x�"+��2
�g�IW4T�ð�(>w@�$^lR��)��p�޵�ɩ�ٹd�W���n�x�VL�e���H,M�O5Ө5"��ڠ.�6<���Z�Gc�w���;0E��/����&0uu������5�]4�ˢ�n=Mq�ݒ�ԙ�v8×[|F�3tN<[-���M?[Ϋ�'9���ĊJ1�F�ٟZ*@�y=[�Jλ�l,�T%���[/l�I�!ŹAh�1`��om����)lP�Vꂓ���O�L�/�#���/�i�0��b v�<z�'n��uH�����ӌ���"z��|��̽9�.�Ħۡ�o+ U��u���MV�}���
��U�B�j@���uf�]=]�Z6�|uwj��7��6%��k���:�{�\�B�5Dn�Z�ĥF�;M�&R���I��4�C3���*´��W��Ţ�v��b������4��Z:���c8��v����z��F0�B�ԭ�Y5T+�js;��u��3�w���׊)ٰ��N#�f��bD�l�Mwt�o4u�d�m�F�f8����u�)�C�,s3Tzܻ��y	7/S����ҹ�#�̅�I�v}p�eū�����;{hK�,M�ıQ٣���b�M񲾗��xY5�t�N���#&d����]<L����̺�}�Dƺ�Ҏ1�:"N��x�(���,�۸�P��;1fҔ!�}�6ԭ"Ȼ{�%4��y�kI��e�s����\(����n�ɡY�����R\4�sf������rc��PUҮV�kTt4�l�vr��¬�N2����\]��7X�\�Emt�YQ�ϋ���������s����'3B���p���'׷KLg.^��j=:3��Z{& �y���{*�z�6�ݾ�C�]�o],�H_R|���kX�����	9�]\��A8���Q���7�*�K��J�v�Ќ�&������u͞�&K���V�c�-<�j�����^��UΆ�\ѫ���/Ws�SH�p+�꒷c赹p;��+�H��_p��uܫ�6�NE�!���u��_m$�V���T(spL"�4�+N��#��`a�6[��cHΕ�G	ZM�te08������d�6��)�J_F^I�7�/5(d��Skgc�|��.����r�&��V>�l=o��)�I�	�l�S��.1��DƎ���V�c�t�9J��w���6��waYy�M+]�A��qK�γn�>���b4E���]��[.)I�����E-%�us�D�j�$[��)�����%d%�A�P��֫�ou> �5���]��AK��m��'u�s/	8'R����©�W���*�N��^虂���w����;W:NOwD��z��L3�*J����V̭v��֧Ug!�]��T
>���2��v�i�6	q��#a���3B�[s�v��}|��+��s/:���Pw6N-�H��K��$|g�+�̰y�xK��7[�CM$�Y��p�'
v{��A8x>�����􁒊���p!���&񕱭�����\�Y)��Pm�m����N$�5�ve�q5lbŻu��շ0>��G�[V�T�v0�ܖCv]��Y�H(�b8���g@Rjh���R�ȱ������I�n�M1�[�����"�e�4��M�;�:�ii�t<�i�;�:�\.�&e�t����Q&E���6b�@kQ�@}o#��!6Q�9h�tǚ�;��J��fߌ�录���W.�{t��IƷq�p�D��gU_Ӯ�ݖ�	79A[��_��Çϒ6�P�6#d���5s��F \���hw��{I�<��:��9��ӻ��9��@�G�&`=�zLqf��քtH�Q�Zp�k凄s��1:��*F`��#�盝�o�j�q7B����Ͷ�8+z���Ő�A�,̝�5B+4ٳ&��]6�I�W0����=��t�!=؆%�Թ�s��E<}��id�j�����`���(1����5g7�!=)�i��(�d㷸޵P�n(Bղf��I ���y����$��A�<n�:�kKt(U�oM�)�WN�Y|늫)d])/37�W�ʖ����)�qQ*\$ J�MG��C��ʷ�H�	�O.��+�S������n7�e�1!`] h)�R��B�X�>���k��v�Lݳ���2��Ob�LU+1#/݀�tp�GK8����������.�-�
�d��vd�%Nˆ��¶u�jsYN$�UJ2�1�j�n���ʤ�q6���79��@�k˂g�<�t]���QCR�r�-gu�-�x��3���r
긒��]��X�j�]�u�m6Ї6�@=hݴ�7�NW�u��3�J�oONqh�K���x>��M��c�[%h��Շpv��e��un���.ISo��I*��T3[��Y����q����2�]����p��\��,^�eڗ���i�}����岫M�T��(.�'�
��"FC7~gw��5�����%�]4�׷m��s��י2��2<��"�T�2x��G��v$0��6�#�d㵖p9��Z�pp︻@6�J����A��I]�1�-�[J��n��9�t2�u�����J�{�v	�ԏBy��{P��h]��
�[5�.`�����%�n۝t�I�2���<O;
P�G�fD�@��߲Q��.#u`�6o>0Ӽ9ô�`��J�}�PS���������>��)ѷǷz����Fzu&�Ѡϡd�]�����o[�!�EG|Lź`
��Ʒ���ܮC;�ЮP�Nc�T�ƥ;��cL!��"��:��sė���s��,c�a�tjf;9�լ*:}@��*�H����ͮ�;r卾B�@8���u��J�p�7�V;�"Y|������j�s6���MѼ���Ƭ���q_I�NbG0�0sΎ��j�4�M�@\���}7Io8�6иr�ꙍ���ǥ*���J[I��r���T�v�RT~�:�fˍ�N�d��'L���>[�+��F�>7�QO)�b:T����{-�
C��dM����ɻ	�x��RsL��Ϯs9���F�Uo19�Ylߌo���WX����ot�9���*��\��F�of�2'F�U83���r���!����bzϐ�CC��Bt�$C:[+*X���鎱q�\�A�)��l�#��%m_X�j�Z�w Yk�-�O���{޺�wD�.f��=�[�e�Y�ܐ�8Ea�����3oiM��$�uy(.��O��@r�q���:�;�N�(�+A�/���� �h��Q���E��!S+�*��s"n�|t^q�e��6��[OBm[�}��IK��e:�J���[Wj�iIV��m���G۳�[ڝ�����B���tZ���g݂��-���-!c5��:x[�r��2>8�ͧ�k�v��ڛ�!��	3hd}JS��geY\��3U��j՝"�K̭E�l������AN�.�J-������EVǦ�-��
�v��ܑt������)�	w]ކb���h���0�F��e�:�J:�Gf�f��;M	І����m��6P�Vz���i5d 7C��Q@^&[�|���"V�oPh̶/l�L��dY����y�u$Ĺ�5�7�+kQ5�؏v�#%eMvh(NH�nݮ���U�U�Ծ	(V�%������"�x�v�MN��]6z�*r�וn��e�����jt��3H�"�n\ˣ�G�ф�:rB�K��%N73#�����#�5��%�Ơru��K6�H�mIu��Z�Sh��ß�5��JQ8yɝ���ʈ��*��;4���M�-�)�$�7$��x�ؔ\tf_`�d���n�b��r[���ݾ�o:t��M�Z&��5t�f�����\��t8��gi�(�gl�CRU��"S8������(�c��}��;�mVY���X�U���B7l@*r��yg�1���E�����gq�x�e��.��G Tp�_[F��Xj���|ގ��jvb<�\��!�쬮��:�ە�Ef��z.t��*�u�����+��0�MouP��>4;T���?����`�G����F{TTAC^I
�\,��(g~5���D?Cv�q�e)�L6K�P��0It͇%շ�~?*q�U8����u�����"¹���;���R9z�>+.����M��`�k ��\�۬��{X�Ʃ�ї:�m�uCƉ����k壩��+U&R��7�u`�Bna"�Vj��-�J�Õ��V�f��d�{�U�H��f�;�cD5��K��R�˝�*���]��6��x[�Qӕ;;:���"@��� �z����4�&��=-�TZ5�w��;�$GY���xy�ҝ��7��fb2�Y�ѽ�֯�N��Nƒ���W�r�ܻ�f�r3�a��&�*���5YѴ��ȷK�مv)�K�����ٛ��rF���;1d��LH�����0Q8#����x�m�N����@1@nջ����ޥl2k2�d���\�}vnZ �&�k2+!���o7��6T��̷Đ�9�h�$��Y��$�!���,�J��v���W
�AWA��0轢�J����0��pJ��1������ H��[�+�钬[�X�Tt�]���ѭ�5���-����y�7�D��o�x%�5�(;�ǒ��Abr��"fB�+8�J�[B������J��2䡖������Ý{c���v�Ґ�(� ����V�p&T��mw*���uGGP�`+z�\�؁G�����ks����f��H,У���s���N�@�sY��`�kl�U�[���������:8��L(��r�P[�G-���=@OK��n�P���"��tstP2���![�C��!0c�Ul7F�ͨDΤʮ�*�	�$�8�h㎻�`��*������a�/�\�ֵO�v��j�8vL�n�^K���i<��A�Ӕ4��G��W�C��t�y\�\��h�̾�^k
�%���G����Y	�l`K�6�vK�s>u.����yg��0CkTp�8�e��`gH_.U�u{��g+,L��6@]Z��S|ҧ,�`t��7&CƮu���$�ʇ��TX���r̥e`�]�vs]�4S����$����w�>�#M�N���
kyfS��R��k,Ձ)��L���8z�j���޼T���u����
�u<]y�'�f���2C:�f��g��ي� o\;l\6Q��m�ঁ}Y	1����`���(_r���}�#�Ɣ�Fz��%�c��[���O.#Ö����O;PB��-�Mj�$ц������ ��7C�lU�M��Y���GLGG/
ɒ]��4��A�&�l�}��A�����[>�����k"Q�ݳφvJ���1�Czv���l����H��5�|@4�5tUe���t�_tN��1�3�*Vӫ��|����ۜ��r3����2S
b49B��4ԭ��4�'6����oY�O,A�9Z�5E�R/6�) ��!�P���wyws�s��Dn8͐�bP:ᅌ�)]�'��J���+8h����y�
��
�WX�}�j%|7>�o-J/��p}���;�����{��:�ȴ^o@��u��ՆQ,�W�z3�eՈ�vD�t�;@��3��\�M&c�9gKtA׷�V4SNN��x�0	�ٲ퇖��\3S�2å[٭6���L��԰]�r�{57�	��U�@���:��Z�`:�Qi��h���̣�.T�+�7���0a{���P�%!�m�D��sM�Pr���U��	4Jr���Eiu�7T9�z̨�R�:.���-˶�3��s��Yw�j%�<nd��'T�S�t*ZgL�[�������St��0c0ݵ�,t�ZXr����l���z#���Ƴ�7l�i�k���i�fQ��bޔN�h,٪�=��@����f��V9ޠ�̎h|c���_(7�P;N���v��t{{V�w�����B+Knp)��n_cͼo�N���ن��X���E[�5���f�U�6�T �:��)�%��;��v�@��=�ֻs@�݊��u���<Oi�Wj3M����7lѧiCY��,dR�L�:��!CD��#3i�-�w�7O�pv�a�Q���7�}��6^�޽�pGqd�����U.Z��e�ͷ*�3i�R��&m���V�# 45K�Z��ͦ���5Z�1��c�Q9y��gMk��I�w+F�,��|m���d����w)V=-���CX�^
(a�ٓ�U���w�,u��v*v^��ŀ�5[Zz�J(�i[m��zr�Z{��5%�P�6���3.�Z�95�m�k�H��ɲQ
���U�'՛�.*{u{|��ٗnY��hª��s�oGՕ�R��ܢ��D�6�]
w  �oo�w^έ�4ѷj�9�����M�hr�A��-<�PZ�U��l��v���Cm�e�^�z@l��BT�W|�M�Ao-Y�*�y�0�eֻ���\w����u��[��@ʺ��nb�	O�Ï��bR��}4�-��XY�[��B3���,��d-X�T{�]�e����lV�]%�E�c��)�tx9�ajY��Y��Z�|
�,;H�U�+�<��}��<B��7�Ǫ[���::��FU����k%�y}Wv�d��+!�eb�,4%=<k����\�ޙ[��hrX��QݱDi�^;�*�5��e6TԈ_�����(��	�ԙr���Ih�5P<{�v��+u��[ӧ�=Ӕ��٤��f�g��V���"Y��B�h/hi�q^�\��$��ݱn��w�fcS�D���| '1o+��L�j��Ë��}�b�jX [uՂ!��.�<��Zٕk��/����^[���\}W��{����]J����u�^�6Y�|.��\��Lk�%���"�w5X�4:��X����9|�k��37B�����T
�O�hm�.9�N�D��5�b�}(n	��ρU�\B�KHv����Z\ø��#��'�5��ݙBM��԰�.��Z�l�V��P�oH�-:�3�q�rq�x���B�t���K��3�0FL�dݻRH�A�q+���j4��^�g�z`�+&"������Q�v큂f:�xJ:�u���31[Cp`�RsCE��E��U��Ɍrz1+��6�ޔ6��?7S��y�a[ڋ!���pݻ
��I�����eѱ]����j�b�������n�4.��*u��FȗoTŵ'䅂][�z���m�칝��!��U�r����x��Ic�?���K[��=mv��pv�N�6�˺����@��}F��{�����V�Vۼ�1�[��`N�Ӡ��3/��C2WB�"����RQ�uXtN)��D��e�"3Y�V�8ہ����,��w�i�h,�BT��lx�ᆝ���Յf��Эeַ�Y�dV������un�=�u�g^*	��LR�?Dwd�[`Lͩ =iV����00��*�_�k����`H��ʝ����dN}�V����<j���H^�u�>�LE4�s��b�]μ���2����È�u�R��à�˦�������1�Er+�짷�9Y5�����j��r6��fRO�l]�V��ŮgZyh�}�n���-�%c'V䭬��Ƥ�m���R��f�6A���8�yc��Gɺx8m�ѽY���Q�V1�t��]���5�ș���b��L��"�n]
�V3��V�M��bj��$GD!��թ������w���5���#r�6 �n7B�ގ�H��WV���J�z�����;�6Ձ�mي9�n�r�]�<Ըf�t{V(8�S'	
���I?&��������x��r��ּ�d��v���z�m�Ks ���h�tzN�A�W6�+&u�k��4�ֆ����V79����<ej��m�Kt>fE�2#{�9��"8�u�C��wCU��a4����U�\�n�vÆ�q��#���d�݉��:+����o-�|W+�p�}z�CeZ[��y�ᜫ���F��)j'�UdW�X���8��U�z�{�Q���]Z�X��|igN7}1��Y�n�P���^�B^.����#ԍ4��i�r"�gu���kGU0��E��#��P��F��r���$�u�L�Sph4Tn܊ɡ�VaWoq��]/k�F6M,��+���B�s����LK�H��w8�,��&)X(�&�f���[J)��S���A�&��뱛w�����[�,� �V����,+%����n��\.���	Y�c!]
Z9q��t�����+����O*��ф<x�Je[Y$1X���7�FlV��1Ҩ�(@�,�Hf�SkQ�!�}u�?�����q�&�mթj�ΐ���)��GR������[أ,�+k���j�ja9�N���^+�^��b�g���r��]���9�s`X��h&�̩���H��g;R����sd�؀�%���+{`�uc�$�cO���C�q�����g/#Uҽ|�qQ�zh��J�����q�W4���X��#�C�NU�Y��E]'E�4�OM.���e)Nb��ζ['wW�oa�h�~Vƹ��$�)wȹ���&���
�o�i�P��8BZA f��̖��Q��|��E��1$�h�}[6K��O������O�-��5q�7+!��bP��l�3�$k���<Ձ�L咭��΋��W9���8���֥�mg1D"6k���%�#��,ik� �."�Q�S�0G"��N�����[}���WX����>�{G�B�>7�^9-�Eu�ՔA���Vڈ)v��5k����W/���%~7X�Z�e����5�Z��v�<L�9R�ɷ5AX�v���ꢢ��nY�e/1��k(�9�b��vbe���uJ�uAM��Z����ǧ`��ܤ��UU��u�(��ҺR��+m�3�R�-sR�T�[s*j�y��Ҷ]���>r�����-G7[7Y�&6\�d�+Rѕ+Um��Ko.�kUFڨ�ļ�k]K���[+�\4F���n���|'���|��w��3Y	��K,��e�gI��m��ܼ���2���(vN��o������g5ȥ�N�/�t۷1�+`���-�ڥ]ψ���0���/c>��#��#3i�|�u��}��b�t-�O�+s��g7�������L�z,n��Z�®�o5b�>�S��������ٲM�F$k�M����oL�m��c���*
�%��Z�O��LV6n��ּ1J�7T;7&Z�h�l66�A�ve56�d�6���]T,��Q�n�"��_�T��h��'wݵ.��:X�!%+���m��S&����q�zyw����T{I��k�2�ܪ�4D�{r
T�Y|�X��ֶTj��t�7n܀A+���2,�}D�V���ju���-�n�ہ�WOd�B�mΆ�&�%���s������G�I�殣D���_'<��K3�_�E]{���c�
��#^j/8*��V��h~=�g�D�_3�#������ܠ4I���K�Ͻ{ZVv�B*U�>F3]쬍��t��{"�f��:7�VsIL1Z�U>֐ј9��'8��cU8{-j�bh��d�SSSo_�<�2e�kk;Y��s*�D���Oik}��67r��fz�^�ND8��C<+��̀��n|�#z���Wݺۀ���A�4�pXm��s�D"j(�5n.�̜�1x�P�b��[�劌���A�|�H]
�z��Q����ԟt{{k]΅�­#�!���{6챋��v�����d���fkM�n���������Km`j֜w2�o9�c�f}��ӈ��MS*z|cr�qG���ίJ���Ư��wy�f�+���y�I?i>�x͢�Wg��pm5`嚊m������:�<�ek�UóT����O�Mz�M�3��qű&3M���h5��wC�O=�zD�����Z�,q�\�SZd܆��c��x��3�d췩*ʭYk�EN��	�%�{r�1�KJ�%Fl�}ou���>�C���_,'��-7���(�ҧڶ�Mry㱪ީ�\�h<w�א�[>~�Ʊƞ\j�/#��L�q ����/ao��yݏ�+���x�5	1By�=e���Q�3vi������n73Mn����>������E�� �όg�ML8���S�{����ޓy@�-�]�Gk$6؛��kk14��m����}2!:j���DR�Q�����1t
�c$<�J��Jx\�(�b����4�b�;�+#,G�<F����+7�&��orV�Ǝ��27���8��z5&k͞Ճ5��S�`�!�Ԟ,�xˋwr��"_15�wu�[����g��Lqչ��1('�떮���f��#:p�+��2�7��.�#�Ϩ>��np��*�ie0PSK���Z����M93R�4�C�6-�sv-8{= =���⫨#=6���]��0j��V=:vu�i֧�D� \F�O��ϝȳ�2��reK���&L�}�䧋����h���5\.jn����7P��e��iؑ�(8���dxc��xx��-��^v�̪������n®<4h�
��bǩШ����>\�HD��Ϝ���a�jϕ�s!a�Q:�r#�L�b|��ш4GX!���d~qFY^����9��k>ogt�<��*����t8�G:3�&�ؖB��R=��{�ky)��%2*�ǢF���dQ"��5�S�3,��3w^r9qp�G�qӍ�.�,@�P�J�_��dZ����y5K�0p��׌ �B/H6F�ȈD��O5��LQa�s���>�0�w�6�u���M��l�O٘+���v��)kO]�dR�{(���]7�E����<[�1|z��Vʛ�����'K!���8-���d�t�Y�yM�(�-ރ�op�>�*ǉ��kЄ�T�י4�=" ��^��;��ٓ���/��\�I|�CR�y�rׂ��P�"�|r��6��rD��<��$��@\|�eO�ˇw{�s���Vj��D!U#h)���tO�t�40��\����^�صw�׈�3(TbY��q!�TN��P"���ي>w�@�ۚ��&�&x��H�� GQq�͟erc�g�������;{�]Xl8���Z��F�p
�=�F��w5���
L:0��=E9�Jv(2<C�U
��ȩ����o��&��ˁ<F��� (�GS���n��\���}˝/L1�(P�tz6"�� d�B'Ďf���Z�P,��3Sڻ��p9�+o���R	=-�`w�����������,��]x��rb��}3z�wGM��Z��Y�-T�d�/�\2��.��^�@y�T��G_�;���*�A/il�u��]Bq�LǇVRm�<L�d�#`]u���f��2�GN��ڂe���D(b<���>ӱC��h�P*ʀ�c9�n�"�)kT�[7���:>�>�Ĩ�����M9Q���ٮ>s�zk���҈�b,F��^���̣�&B��3sQL�U��[:�s��0�f �@>Ңl�t�DΉ�G@�0)5Bc){n��m���ؙ5�xX����.��p7t��� �B{x���Y�ӓ���������Y##���q��A���]��3y�`��d�3�9���
�-��g*�U�"���Σ[.���qB�r<��u����U���΅^0n��y�##�"k,`εr)�w��:�} G��W��"t(:�j	B���p6{]��(K�����V������@���U7�oT��(i��Mэ�%��1gbc�B#9�'ʏ��Fn+ȸ����>z�!����[D1���i ��n�q#[A����ŗ�}ڽnV�V@�}�l����P���x��
�Imj�D=9�=�o+���8�f�d<=9�Ѓ�:�m]��'���s@�>F�+֫�\��qZ%��Nr|g��Œ�l�&����x����Ϝz0��.A���D(�>��fBn�6�/l���ghL��G�PS+2T;1/q��iVTK��O�Q�A����/�q����}کS���72�:��ogt����1��>*B���1JTj��?����Ɣ���hz�f��b��=#p�B��>7�6:�f{��[�*��m:��N��:�c����^ً8^e\Lx^���ܣb�nk6��-��Z,*-�)r�fQ�Z5�u��ݭ𨥩��wK	�mB�[�[¬��'[���A����O�R���6oHB|@�*�)�!��ޗs^g���^�+���j:���mϮu��0���j��Ȟ�f��(J"IX*%qU2)Qql����ƃ�3�w�� B# D<#d�q0�T�NEƈ�;[mGwgV��@���Ȱ9H�2���pG�A�\Z7�B�{��f�{���7����טd|l���L�r���ҫ_b~��x��w���*��i�P��V/�D�ȅ�U%v�M�m@*:o�  ���g��5g�n}��->�sy��7�݊�|� =<#*d)s���O�#�景�ZD��o4����O�1~y���?u�'�||}�q$�t�
��l��s7��._�Y4+%+������TF)��Z�*[s��xC��=Z%HwK���Ѷ$Ɲ�ͭ{�7��#���5>��xV�i��c؜�� ��?<�Ւ�A��>�x�"A"��9�#���3����ÃE��������^^p��R�ňY���B@���Ɣ>brFD@�9eE+�2C�x�� �#`���ٝ�}�����#��=2n�z��\C-�P�b<
cK�ݹ�;�Ҕ0����P�(�nTLS��-�CHs�z��E�����=�ϦF	ؑ���>�VD�*+�\�:o�m�>s 1d. ��zv'#ـ��b������]��3�ݣ-�+�#��>!���F�8F��.B�RW�g�U�b�nc4��"E M��p�{5��a�P�tg��"�Nﻋ�EY�d X�������������x��>�H��A��4�b�M�1�m����-#3`Q�j�9p�,X�����������k��F	|�v4����S�"��kX4S�6+�C��
�YŐ��y����feI6��1h��Joum�k���qk��v�<b���GhQΚA�~7�ۀ���#)�Q��$7ۄf5�m��5x�U.�<�Է��)�#{�w�{Z��籘1��˽���V��cλ;`���UM*�%=��k�8�c8���G sM$�ߥ ��>#܍
�w0c���Y��c���Q-��n�>r��d��oTrv��؞��i��,�j�&v�f��}��1�չ�ծ(�3�O\��
����C
4�8R콶��N��b3#n\��o�ҫ7,�V��n�3���H֎��p��`�Zv��0ݭ3���6��Z�ҍZ·�7�G|�Bv*H	��uŌY�;�������/�ܮ���Xޫ��)��8)ʂܩ�M,=~���قE�����Ń7yK�5�m��C�fr�kdYڙ�h/���;Y�*�`l/���{��툁f�&���V�+�x꼦)u]Ҹ�i֪��h�00�꾤⥄w}8|�^԰�����S���-�Ҿ�j��K�7
���C@u�vVԜ�{.�虹��b�z��

; �ڝ�͚�v�2���|8�����������xi����d �b�^4/wn�˾��E�ݫ܁�A�
ڬR�)�k�w2���u�yE�[����� 2V����O@��oIB k2� ����\��Ł�]��K��P��۝����-�vy4�u.�Fl��{�q�</ӻ"�
��/|rT���CX�(�{Q[ΰ�d�B���x�>�Z��a�p��3���I2�N�BK��.�a�	�����w&Lq����NTeeb윧mKY��5�<�W���eݫ@z���^U��&e����jZ�KJ�i�jsS�63�嵨��Q�kB�KU�ڰ�`KI]���5��z�m��6�m����U̵ɛo��2шsQ�]��:�m
�C ���h�l5��uh�hփ����2W1*ڶ�"(�ō�kujV�ڵ)Z(9��(֖��D�D\,J�ck�[�iv"Wb���ʕ5���QcuAu+�k`�f��ԮjZخ��gk���rf��em��橛Yv��ѥ�KV�Դ�|�g���ؒ��Y�B�!�D{Wa����"�4��" ǎ�{י�����-��ɮ�O���~M�z8�0�**2�D���Y�h��_n�^���w�n>h��->�߉�=���S��=}o2n{��[�[�qrn��@�p;�2Oxp�(@�G�����6��l\�Xn��/T�Ď"�����ٯF�G´���H�_t�>����=�5�4�AӢ�����X�B���BӢ�U/�xv;M�}�p��{�$3�
=rU�X��y/+5cFQ{2��7�t�D�t(�ϰh�P*ʁ>dc5-׌.���֤��CG�C�A��ȑ��$\��:Q|�CCg=2d�m�\�sx�y�y��C�:# 2oO��B��\+�Ŕ7X��w�z&��V����������v�}�@�04q��g�
�b<cVn�{ɴ�G��3�^�!��:�sw��-s��?'�1ۗ���Q �4T��:ZY��Wh��ZZ�(��ޠ{����ɇr�U��Ӆ�5�X�6t?h�@?C���J���/�z�f�Jh� �~k��EVP���*?�X>�/����P7��a�نv��b�iϻ�T������9�۵oW(7�x�aʏ\�Ke]5bx�X΅^0n�9�:�w{��'��>�G+�+���F��~�ʁ�q��=� ���S�$d4ri4��c�G�N	h�"c�m�+�;v�u�XTo
����u�Y�v�
���'�@p3��<ӻ�nqtE�ez�`]E�
�@�Ș��T���)=ܝ���[ܠh�����#OC���>�%C�ѐ���4�['�]ME��|�d[R@������G�䍊t��*6�Q�5Nd�۫���/���_N�r2y��BT�򛿑p��1<N��i��O
�[Գ�-��ȶ�.9��s��4�O7C���P޶Z�{��r]��x����:!'�:=�B�C4ʍ�U7ȟ/H潽ї-��;����B��_6CJ�U�΃�b����6xx}T�w��B�>U��� A`�#����UnM��%������"�l���|:�쥔�j���>	e��g>i¢��2jγ� ����B�#JGlm���!�n��\�ǲ*f f�v*nd����^�����}\9�)��kQ$����H�,�5iV�\ �5y����י���tC�P��Dn�p��.6$��b��ȋ��vUS;ۏ��G,��^ϕ�BR*�M".8����\Z9ز\+\���i͉~�>p�`s;��v6@��i�X��U�EW����f���j ,$a2u,5�͋4C�G��S|-a�����/��u0�evz�ɺ�k6��m��`���zB�&�NB,�l���R8%�����V�FVi��84�ջǆ�a:(h%��j4CK���,��L8u��G�tT=���ѷ֛m���\lJ��A1 �b2�C���NG��v\�4��uj�ߗ�P�,#�DgP>���e�@�fv�#brs*�=��0&y�h�-졶}�X+���x�*�0�55��[�s �EOGGC�FEP���r�H�  �l:�^���&(��dtD��\Rs�������ªӷ�o��`6b$:0��7=L�E�e�@�K���b1Ov$���is��@q�*ܨ��R'}��4�b�E�O_%�lD1|$K)}l���+��K��*}���U¼�v2�0��e�N���ŞY/%�hj���>����2�`�.U�N�\�����|/��ɶ�u1��Y	=l�Q���ݢ���
�"l唢�٬�<sjw�W��t��~��t �>5��}����%LR9}ۚ�\稛�de�;PxW	�E��b�}t�+ʌ�Pѫo7�t��D�,_�&v�(k��Yα��~a}��&hw�Z�7��'�xU��(�==��R2�G��n���+���w���u�7��s�>��8�)Z���LU?yU��>yݰn���=�V �8��hDH��Q4#p2��8�(���G(W���UL8����p;��#��taO�2;��?%鳮�y��џ�v�����к�������	^Y��`Mf5��(1�al �h����:��A-[�n#�HZ�[��rJ<�P8�ӒDȎ�He@�G�.����>d����#er�����_��@���j�yt�W(z�(�ɷ�˿vvc�n�Fһ����8��my+��c�Û�Mm�b�:���3n����X��N;!Ӄ��r�z��S"�s��!@MÎ��4\��*�F3�7vb�ٽ���F�cNQ譟A�9�����:Q����dÞ�U,|�"&Kϋ�B
8B&t��!AG�
2yS~5ɽK��Co�� u���Xt(tj/�4���4Vm0�&v�l�<��t���5��cAx��`0!Y*��c�y��4:<�@�'���B�6@�VF�#1����� `�U�ƹ��=��0�4v�����zh�g�d{V�	[��3�����:�ea\hK^/�;ǣV�H�EW>�s}���EQ�O��S��41�t/ݙ��f	\�s[^S"c���d(ظ�ѧ��b�(��+h+9�3O=lL��F�J�[��,(�c9nɞ�s��f��"L`H�T,���U����aʏ;�{�bg��\z�%S1��S�!���kV!��3��QG�ULf�rYk������۞�?8����V�Qh��Q�;��k���z�M4!�FӟLl�,�!nO@��EEB��9��:u��p�#�ρ�����z��X��C#�!q�]oM���bvϢ1�i�8�=>8F×#$��i�t�wIVϳ�[; O�GgI�d(_Wr�U�l�ѵ잇f��*�^P�c�бC>�_�aQ44�L3�-,��ｪo��q뉢9��z$!P��E��g �!���'��k����&���B�Ģ������h�љ��2�bD��I�J !aNH`��[���9 �:l�4���d�̜�Z��9�x�����*�m�<��Xs��v|б�+W44z������[�zȯ�����x/V���&lN̰͊�B��F'A��O%p��-��UJ1��(��ϭ̓jfA>#�:�I=��4�@ؾ��ߞ��̽i���(���$Ϥ`�R��V�|�X��Y��V�G몘(�A��ʫb�v(�W���)]W���bW���`b����>\E�"��#=g���A�3�b&ck��U������`B������=2΂2S�n���p�Y�!��N*�0k�x�ņ(�Po�ϕ�]��u����qCb�����n�� �P2%�P�2�Y�O������}O$k5
'j'ц K<#*d&z=~�"wH���a1S���𥉉4�f��>��u\O���E�@�fvF��n�f5Z2.C��p��od�@Q|z7�+�27(�ځ����s�((tD�*,i�QXFEQ�>�J5�a@�����@��5�;;���C�sX_`��*�R�]��4r����+r�wan�fnmh-�k�]ñʻ4��S�y����SvS��Z��S��sq*_�{�e�n���s�������1q�Q+]z`8��L^��<���/�(���6�c��D�(�g�,�-���N��.�l��c�G'�X�
$�V�D�wBp�GvÇ�/��׭QH�kD�[44��}8�����C�_7��>m�9QLd��5 N�F�Oi��I20�	f�>������)��m϶���x8k�"5�X�\0`�e�f��5�W]ɽ��߅h��w��#j��ϨT�b������,$A�qxΧ�ň�n1�"΢�,���Ƣ�ض}Q.!8�'뵭9�q��\�$�	�**6�	�k�n�e���.w9vg5(\���O����db�< ����'��y|Uj(0S}zͼ1��7!Z���9��kˢ^�������3�T��v,�j�ː������"X���N�S�Ć��YЦvP�}�at]�喾���zMRm��Q��yA�cR����Y;�"|O�]0���b�����Bb�\yeϘ_q�8`���,`�t>�q�/+݋3Z������r:�bc�l�L	�n�[	���.;����{1,�>�ˁQ�L����f���b�{w_ p`�^�ˆ 0A��&㡱��YQ(
fp��D���Ց2N����k��V��<�O˄��i���]ɨ�xXGڈ낄N���

;�W�,޹�{��ޤ�3�� *�`�F��%YK����w���L���B�(�EY�QXG	و#A�������]E�Ă9��q�}SN�"�p��*�#1��������ԂJ�aR���{���a����,	�wY5Q��+176��5{���ų�>ܙ�(����Dw�e�5рn�:�c����sK�:a��MW�v�vA��#c8m��yf�	L��]E�՛��7�mҽ�m�.�#���u
�XV��_bSL�R��svt�PM���il�W��>3�����cCG��9{I
Y�ޢi�8�Kˆ*���0�=��9�����é�X���i{���3�����T�|��a������oxj�\�<ާ֊����Y/!�q�J����^sr^���.�U(��7�4+��-t�A��T� V���9�ȦbY�R���C�o
�EU�7m��C�i��1Ef֪wz�ـ��2��Ub�K�{	�uk��.�[��bTt̵��#�0Q;qA\��4BY��hs�wo��*��EJ�/#Kpw/j����ie���9�ЬS}���ꙋbF$�V�ko+!�cw����`�wl/�Ʃ����]��M�G�	�}Ֆ��=����ss�^�Ǐ9�����ٓ������e��]�7��`�V(����d7�J˓��[��lar��d0\�Wurj�Et)Շ).�s6��fk�����r!�������/Fs����ӵ��BDv�<�&�zq�/j����H�E`76��j�X`C�����t�B���N�kT��4�wҧ���8�J�r�]��[�PY9��	Өl��l����Vlia�b#3��2�^
bgIG+(^����tT-�R��V�I��8R��;�SK��e�f��z�����&�j��5����+��Cu�g�+%�f�mf�A�{b6�+��w"�q��3�En����%7q����2c�S��N���x��&�h���������݊]��Poaͪ"���������kR��ZV��֥im*�S:9mV�ҍ-VԵl�Z�[KJ���+sD��%�(�F��e�LT��+mm(湶Ѷm�cn��TZZZZ��6���ь�^2�V�[hV�.�E�-j�[F�TJִ-�R�T�ڵ��-`���Q�h��&�U�Y�nQ�rmZZ������Zֹɚ�ZZ�6gs��y�sm��6�PVյJ��YZڢ-��V���������>��ף���D�f^ta�)`��\4�<6Ф�[���ބ˖ȸ.n���W�|�����}�AcOEM˳rrz�~�U��ed�y?+���kSĒ��%V1R��`俔�������)�X��Y�ݹ��**7��^�* �8��g�I~�ϗ=�X޷��y��/�����Z��ötV�>�wK�C�X��k��~�������Փ"�P���Ă����;d�?!�� �O�L������Y;�̟<w�B�<a_8���V}d�C�y��9�}��_c����Z,����',0��Vs�$zμ��ήa��H/L�;a����É����T��6�\x�_&+�~߹Z���f|d�w��[������Ag�N�UH,Y�a��!Xv�ϟ��AH/��'H
,�L��*OP��%O���������;�߷�3'� ����3����OXs�8�X�u��X}aS�
����>�È
/�������R�{N�{� ���=�*|������>��߼�>��N�����c$���`��;C��}��?!R<V�E �?QI�
�Ml��0��NYĂ��ݧl�E9��ϼM�]����|����T��w@��N0�|d���X�g�J�����)'�VOYP?%2�_��$W�(d�!X}aX��|�R��M���;�;�]�s�;&m��M3JWOFN�@�v�������Wc٫i�v<	�N=!G��Yzy=�c2rýӥ,�	��; �Z�G>�����:뿟>y�w�R��N3��P��L��+'�j�W�u�Ag��o1��v°�=Ԃ�|-2��w�C0+Y���+���ߝ�{����x�)�A@��38ô�
/Z�̟YP���d�Ş'�3�$�
μ�dR(��*zϿ�8�Y4�f�a��i�Yλ��������~���v�O�
.Cӻ$Q���!^���}R+%g|rO���"�X{s��u�Փ�釾�d>~���+9�PX����ww|�}����>� �}��u/� �o�fv�P�iP*AgS�'L�;��Xq�����q ��%~��I�TR:>�3'��<}���3E�v����$G��
��dL
A}��3�2��0�²}eH:�!��� ���E&g�JÓ�2(|I^�u�8�Y�':��:!X}aY���޵�����ߞz�&�Y�=>�����T�����!P��Y�t�Ru-��i��R%eO� ��X�g����,�<��}�n�9���)� ��|�q ����a�:L�_X�>�d��ɒ
N�hy�A���a�5 �,��g!��S"�R|�����_}����>�����k���הS0���'Ψ �������'�d=IR:؃��2z��2Aa���g�J������02=���Z�������L��
��� ���N5����Z������~��oӭ����.gl����+�+�,2A�i��a��Hy�~�������u����z�2J�̕�0���%x�l2Aea��<��VXW�X�Y�Y2���*A`>ڐ~R���8�P�}���2$&�~����>s{���Ar�C�v��C�.���au�ch�O)ʯ�E�xaf�|k6���{�%�j&a�#��%ҝwe�Vwv�[R�Ԁr&�v�n����Hm������|H,�?��� ���3x��fF'�Vs��g
��@��2^�V~�C����ӌ풤�l�X����{�Ͽ���Nr�z��a�u������~s��P�AC�\�`�|e�@�3��� ��~������!�J��fH=��&!7=��y�_:����q {�C�&��� q����I�O����:a�'��i��?$�UXC��������:����+2!m ��
��T��=��q��*^S!�J�/G�C!�%zN��H,�P�b��}��H{i姌���z�s���ן>�������R{틒���0��� �@��<L��*Ad��t�AHs�t��<N�d��$�
μ����3�D@� �P����V��w�r�<" gi��\ ��J���f�*A{`}ԃ��I�V�O�T�ʓ�ϛ���R
z��,:II }c�ԫ&5}OR�/��@��6�*J�Y�l��VT�홇G�t��
�^K`,��Y�O*J�H)�N��+0��l�'8��9�g�_=��u�=~2q3'L���v�i
����C��?Xfz�̝O�d�°߹�)�}E�a��`�P�%gl2d��W����w��n���Ag�|�}��B����Hwl�g+W�����÷�Y?30ퟓ0>�� ��2d��H,>�ʐY<�<�����矽��/VJŝ����������$5�N�*ߔ��
�C�2A{O�퓌��Rz�|`V��HwiS��a��}󾞼�������4��]��I��-ub���d�ś��u!�vXt�+�'k� Z�g^ֻWp�z9n2k�ͥk�9ɪCm�r�_�:kR����.z���I>_�>}�<}&H,��x�Ԩ�8m�}k������=���T��RT>ZACĕ�Y*A�g���C�T�$t�_U��̙���S��C��@� �G� �C�.�;C����>��Y8��IR'�s�8�~�aڡR
|:�f~g�fّH,?3��w�_<����s��AH>�|�;a��+>�2$��ξP���q�
�\|���;�*��$<��!Y���/�R
AO{������Wլ�O�S\�|=�q3'L��������AM>�v�$X_,��;O���H)*��?l�@QgE�O*J�H?��x�XT�����w�{���{�y���P��C"�`VN,�퀯�B��;��}�d��Ӟ����Ĩ�twf`x�� ��d�����$���J��r�������7�?{��� ��J�RVs哌>��:B�}I������*AO�Xx�ԅa�wl��'����̕���E �z�?����u������ݾ�>$�O�v�T�������faQH,=9�C���ܰ�a��~u`d<IY�G�N (��9���
�U�2y��+w]|�o��}����~a�C�ﴙ��VNKUT����� �N�@���3�a�8Å�@QHp�i=eH,�VMݒ�g���8�Rx���~��^�����v�ݓ (���q��
��*A�P���~aX�sX��*)^��&H|�Nyf:a�� ���>9'�Qa����ۿ�{�y�����g�S$h���a�Ag����J����*S$�o�Y8��
�)2Ag�sPPS�O�R
|ޮ"���&�｢�fV��Ĩ��/2��۔�6z�T��+ �%S��@������6�y��|�hN�Z]�k-�[��PɲP�҅�\C�	�}UUs��������:z���}V���̟��fed���jwi ������A�él3
��*Ag��o���Ϩ��'�]a�ô:�W=�s����? (1�#��� !7>�q�Y:�fg�Ow��׌+
��Ӵ
��X~eUH,��fmHp���
öq3?2T�̛yz�o��~{�ȧP=ꙓ�T��X�JŜ��=a�AH�B�yd���s0��~�*A�~I�V���3��$����Aȧz���,�<	>y	�<x\�ǔ������O�I�TY�L��9:�
A�ï1�}���l��J���"�P�>��O�|��|�κ����W߶H,�
)Xt̐R:ج���B�G,�Ïl�0�9a�����u�θ)!ζ��T��Ώ�N0�P�8~�G~�﮾y߻�R32q8���^���$>��ö�O�8�P�1��T��L�P�3;d�y��3�*C�v ��%O;���{��<��U �����%�HV��a �~��C��E'Gt3'���RvJ�ߨ�l8�P��(fs�&I�)�a�=d��9�O|�;��{Β
AꜴ��
���g�g�:�g_Y�8v�~�4Ȟ+@��9��Y[ij��(�$`�}(���>�{>�"ٴv�P���m��R��[�pP>~��:D��uןɜ���5�ஆ�u�y�A����Uڢ���#���=�+�d����;a8 �(���fӦ��|������[t}`&U�GU䝋�3�ySq�e�ww#�*�������K4e�׽��}@x
5|�nQ���W�r'A=>@pG��u1����xz������{��b"��>��#"\(Q��0}$lGK5����R1<�eD�Q�O�S�͈�U�Z�D�)���of�ss�B
"p�=
���eϭE���2Ǳj��7��� 
��R~Z��h�z!��x]��\�g�}Iw50XbAΟQ.6P�ƑqH؏zE(F�R���OS4:l��A
')Тj�g��}N�64��egR3z��5)��9
T��V_E��T��?�Oɻ9��ё�2����?-8,Q-V
2��P7IV؛zЩ��G���u�Q��dml�t��P�^�p���ő1n4)Tz�b�^ny�ڳ��!�KpVUe�gE��'�:�IMؑ	�v��)�[Оa�P��;[ow���]�{[�-���_f�7�+58ud��8N8�?������{������A;T���Z{��AjEq�EG��[o[xځ�B<�n���@~p�L�q~�KXkG˅+c4��qsQ�E7;hH�ل}$�� dtѐ��FƋ"y\�*dع��'Q��=��Xo�b�\�UG�4G�X}�;�(�����-����E�>Ss�������L@Q�2��r�{5SY�dF�z��$<"�Ν���>�@�;�D����E�V9Su}�)�z���H��#���Gh�l������f��b�j=aDq26�;ʅ"p�b��\zO�n��ꦵ7& h� *ٌ"I�.<Q� .5eE'>.nN*]���ws��.$Ga�6����&8��Qx}+�_y�740n��X�/l2��^�v�R���{��WS* xxc���XO�_���}]��ҭ���ꥧJg;�cⴕm��l/kT�*l`�������L�'ɺ��9�P!���#�+`�FEM�Q12:����^�:%��"��="##a#��ѳ��v,��&�V�bJk��D�:��Z�U�����j���u��*���1�H�<��q��U3����Ao�΢^��7R;E�tt��Y]�mr�$�F�zGG�%�Ȩ��(�0�U�q�@��&�,ݫy�(����"��,J��$��ȃ���#�GQ�Ǝ�֚۬���u\_g�s1�=�v� {�9�x�wL���dJ�U>�*���b�1U��D�T����j�Rv����F��ؖrc�P(qP'��ta�:#��ucM�D�P�4�b�n\����rTls.�F�D5��J}*5���q�8�y�.C�2k�vE��Z�o��_fҤ�e�K�w�bW7��&3	��UgJ�l�]5kJm�;L�q�;�1��$�ޞ���I����5ټۏ|�>s�'čf��p��L�����Px6���ٝ�40����p8�ÒD�}A���.��Rf�U��P/޹�>�\g ��H��"<��ntMd��Vߍw%�����8��r,D��i�H�9$۝�
v�&�kn{�jn�r"=�F� �0�L���Gi�ˋ�u��R�N�*�\>j&Wx���� `�Xt.����aEzZ�(}-]]���!Ģ(Y�qXG	1OTS�d]oyD{�����	
3@0�cӢ�6E��ϔ27c:v�Ļ�ਝ3" ����#N�D�|��<��u��&X�u�������4��"����PTN��Չ���3��I�d��9)�d�����9�ח�}���Fv��J�r��=6�B��]��j�*�p�b�*�Ϙ*Sc��6w\s/T]�W�Ig���<=S\�7YC��dGcb��z>�^�P@ѣ�H�g�ԉ��y�����R��%��T�uk���6|iV��� g���/�ۼ(j��#DMR$3�팟��iͣ�T��]̪ǉ�E�T�� (�Kh/����g*ei~�]#��Ғg�js7�訨�tFF�χ@PC={>ʕ^�������I��<#"C)�B��>�� ���'��;'4�bz��l-��R{
���c�ܴ\ h���7�����˜�1q�!��|<�=Լ���0�4a��b�pך���q$�úD�Q�뉚��V�C!\{�6����DC�,ZgO���� ̅�ÉGc��d!��%V���|M(�BO�
�%,.I[T�72��k�,ܹ/�J������4Y����X�ܬ1 iU�ɠnlkE��}+��ٸt�"l�J�阄�B��,U�u�}�mN�Λ�%��!m�颖K�4[[�����N�Ge.�\͵�:m�)"0�3%����AV+jj��i�\o�&"3��o{jݽe��g\�[�$�^00�֙2�36��_W��1�)d+���a[Qh��&cLܵ�h�P�O����v�7�%�親����-
���IC�+[��I��U,��
��U�ܒ�¨$��{]{\�F���΁�|�	;�uoW�uU��2 55�Zl>��������`ϕ���]J�s�ھ�8�m]17��K��C���݈\2��X	9���:-[t�t\�>ۭ}Q$v-�^S���c�ю��5@�t�⺃��\\�:]h��}�0$<L�j ��|�+��6�;Khy�ƣ��B�=�W�⼌�Mv��t�&�t J�
N�^�ݻ�4k�D���S�M�r��8�f�i�Ca��EK�(楝bk,��7[3�a��*�iA��#��X�4���P^�F�f
7�k:u�]NH1��3��5�j�S���짛7h :R��l���3"^+�z�ݣ&���V=��f�!j:���w)&z*=�T3�t��]W�P8�$A��;!F��B�yFW���Nn@�;��{���B���g�[��� �nP�XM��jP�¹�Gbټ- ��M0^vf�a:ڸ.�K���Tj�1P"@k����D�F(3s^\��CX�s�:�fk��:��qX6N���I�d�I��-��SY
�g~����j '&ε[ZW^7/8r#R�����gJG6�o;�:��\ΡBA��^�#�O���43��f��Q�x(( E���Sb֪VնT�f�3[�G\f�V
Z���C0��MlZ��֨��5���.�:��QrZs2��\�rW-QMv��(�֥
�
�Ŷ��v�k-x��\�iQ���"<��:���kv�gQES��R�Z��V�]*��g9�ܢ��ʶV���E\6�r83�u�w.�CZ���hѢS����ּ�.�\�7'Z�)dF��R�����j�s�nq8�ev�ys��P�j�lh�Qv�J���Q�pf��x2�1mh�r�(Q�֊�ͷ��}�$���ˣ�/�K�֩��/*d�ll�m^T�I���.���~U_}�}R'{����B�����UЬ޺C<��i�i�f:#L���f���H!���>��
=��7L@6i��T�,�2s��.��lϐ��l�!C'�G3�pX�]*�FQ��jx�VKXg7/���WY�F�`t\L%��x��w�E,���i��"�2?�G��On�1H��"��8z|���WDF��­�N�>q8N��`���-�GM��É���>�;Q����fj�d�3��3BFN�3�%ǲ:��}B��SWX���gk��N���ʎ���9� 蜌��ܙ ��!�D�{1���Z�+Ce�}�|�HZhB��}�
<#(�yֲ���5=q�w#�X.k�L���ϭ�1�>�G���6�o]�ݍ���,�:,M��Er�;S�:%Ǚ]�uc��	g�V��f�(Kę9f&I�"�Ú�,;|��e�ڶ�V�-<�LŌ���N�}��U_d7|�s�"���
����8��#��*vP�-�R�ʹ3���(���C��(�q:D�v-�
+Ȩ򱊔n�i}�1��Ҍ� YX#'f0��2ϥZb�BʊIF����o�O�#���kX��a#NV
/
�1�DujyϪ��g6��l!�AB22�����D(�H�������i^&�r�a���M��6��"1()��8�J�`���(V���^��ƀd���>���ᵅ���9���[��Hȕ3�o�u8�0����b|�Ϯ�TT5�j���k��Yv,]��������.��=Iq�f��Ȩ��(���F�x�w�Y�����x&h��e{f(�z\��8@�Ѯ�p�n����Y~x��el�
�UԨj6�N�w.���]b�R��s�T��hS�Q]�,u�P��|���o�y��h��eؽ�w#�]צ���}���U����>��/����0��~ *W��\両g`Xgz{[U`#���"]m����ג"6FO��w��^�֜��Ը[.+�Q6v=�Q��l��b]c@fW��y�Z�z(c�H�	� \V�N�G�EϺ%�p�c�tn�t�K��]��C� f�9)xd
�D�������qs+�h�]==8��Ǣc�<ˁ���$#�������Yk[�0&�F#H��2⸈�K�j���(��ޗH����Og����U�Q�nFy"}�ѧ�`�XG�u�F9�物�όۧ���ٮ>�GB.'F�Y�{5x�p{�V�&�W��L?���K���b`���6�E��f��k|�Q0h��ֆ��L�Q+��4p��Ì뿞bS,�iWe��O�:�լ�[
����Ez���9{�ԓq�'rM�f�/�������f�.O�D�b|p�	�	�j��0Y�qC�1K��Hٵ��f�ц\}�؜X��ĕ���E�����/������sG�qA������������b66yx�!yY �כ0��ޜ��������ENq�����ܙ����\��
��G��^�Q�=���;��#j�׼��đ1t&}�n6�>��R��
ϐd;�K��˾�e%�	,Na0�����3���Ϛ�V묢=�לn ^��ߠPg���p2fxC��=N�4v�Fx˪kzR��yy�QRgEh�P���bVQ����p㣳׵��E���s���Q�2�U��n��6"28ޙ�+t:^��".�Î�Sջ�h*6)��״rAz��R�b+oL�Ýւ�X��'gQI��TZ�Υ�/��j�	:Sm��l�j��)u�e��f���n_u%����u��4���fC�
�����`8���)  z@��[�5�m�S3}�90M�技
F�XT:3K�(q��Db�������ν�П(q@��"�ʀ.��L�C#���b��u��|6"*�+L����i$>6ˊD��GNI[���P�PGF#�cd����T(�����C���U�j�7u���8I�:Z4!G�:i���|nu�(�r��m��/�g:W�)�cCz��Uo��
�"�V
�0z"��Y��͚4�Sr���{ �tdL5�6�$iG;�K��rP��&H�j_�ʗ��	h���uQ�*{��c���w��U�%������Z7Dt���E�Dj/O�<�C.���0+��\}�αHČ���ݴ�LzŉWE��Y����u�]}4TI�q���M�l��7UwtLv�o%���n����l�6�]]��1� �
��s�� �����n�"�l��6\�#$l�>�K�du�2$3��r�+�l���Yx�;A�9�;8h�P,�@�R�a��X�d �^8�nbu�6���xг��d,!A��O�@�#�3�Sn��Z�'cήD�t���f�!i�s�dG�G|�ȹY׋��W�t2F��tFĲO�ԏS��(vȭ�X�]��+3����.)�!�e�2*��̆��m��И�P$B�:��,�@[�ju��V��J��)��2�2G@#�9��C@�!ve��U��<cH��S�m���:X�L[c�
�� ��Z�&�MJ��ʑ6u��>"##4�v=|C62驼�'�z7��]J��(�ţaCS�dџgTW�
�c����J��� Р���"��B�eՑ.��"���[��*���s�u���RK����{ޮ���d�l"}1�ۑ5ΔV n��A��y;c:Od֮m	/O���0�>QT��K�F���Y7j�̬�H0��=4N@V0K���	�Cde&�P��2��^�Z����\~aa�	��-�f���j#KƬ3s�=&�f�4)������0��~ *W�����9�1{m�)������*�����y"#dd��껬�y�jDa�	$9�JvgbD�G v��W�E��+zw3[qb������C���u�q����e+�d�o��O���LG�@�,D�9�8E�(�X���6t���ջ����s�09�4�O��e���&�!O�$W)5�k.D�-9��5����K��d�j8��7��8Nr�N串�hu�Z	��f�f��-�k�&�l���1�b��i�kbb���7����{ރIcl������PZm�2\w �gb|4�l ��La�N�8�GӲ�ܶ����tU��J#�n�y"x�Ϡ؜�Kb.o��{������=́G�|}5ձ|����q��:�# "n��]�]ޮp|�ʳ�x/�������@x- ��/]��՗ى3}��I�șD��p"	�󂈨0�F�8�j�ܝo���c��� �:��G���S�x1�>~�ml����B�#��t���,�&�F#!��&.:���'$��6�;����]C�厨�U,+Jv�Y���G���չ��&t�5�a�Xj���_x��g����?�p��SP]n�w����0gM	"cjg�Pn/̨�>L֍�b�oܤ�A�E��ﴭ�2q��n���pFdD� ,>B��F+3F����na�Ou��cgML�D��Wu5�� {r��Ħ�z��:��}��x{�ދ�]ɸW��|�G�N	�H���q��9*�T���(a�NL-J�rr�����rpi�:�������zh���1{�oq����!P�pdL�\h�F��B��z9N��U�k�O;��g�5o�0`���4�'�
#W�A�2'ȸ�i�I<���1�E�s���
3O�[�͈���k0�2b���� ��#�&}��@��GU�B�1��J�8p1������s��"�C팈�_��EG�&jBE[���L3|�>J �p|DO��S3��OD�}2e�"�:ȡ=�[[�׌Rh�g���vA�F�OH�MYL����!�j��>CdU/����8\	R5�Q�4���Vj7^���S#W֬��]��6T@Y0���"Xz���[z��ӝ����Y�4����f��ZvK�qL����f����K�dlè��C�着���onn��2/\�p���B�|Dr>�;�I#`,�t5^�r��ˇd(�#dR��F�� ��k��9�8s�"�1rj�a�}�ȓ�Jg�%�kB����g�^P�M�ikF?K�]ft�e#A��|`W���>�.$Q�U�9e"LuK{���\8
���]����U�`֭����[����T4�۱��E����&@73��v�w9!���x�ff��ȹ�K��Ѕ��(d�܍�q7YV�{y3DBdav="���#���~!i�s�>��v"M����Fy����D@�YX)���^>c<tvEW��t���h�@�p����0Ȉ�S�L���X_}�p?1]uz5�2���ɢ�䄤+)n�9
[��B��ޫ��ū�&q)�ZE�޶ma���s�*��Z�Z�������ݎ��vt��R<��	j�2p�/``�{Œ�Z�.�G;����t�U�|�T��w<*�2���e+��Rt^�c)\��j(������e���t�޶���f�� s�_F�)[c5��x�Y�jc�8_M��kW��4��w-)vu��`�W-˖����
�}�WMR�:��T�İ�T�}ƛ&_[�	�����1��nl�By�-���s�+�i�swm��P<�b=W�īu-Hz��	�Kq���T�+$-�oFܚV7{�X�V*�:mC}*^�9wV���9���×7�:�Y9�`޻w�����Ȟ#��!��~�	+���D-\���:[�4󩌩[AZs@�5@�5��h�O[���o��cy�f�V������:[u�)����FM;�*wJ��b�a�t!��R5�V� ޳T7Lvwz�=� �lz��nR�q�8����������T\�^�uu|EN1=�����Y��E�N��faM��8��Jݿ�v2��ć"�Ō":��469�R���Av����]�15�+�Vݶ9�b�����5�V��gr�ϛ��}��S�+��s��4%�G�2�j�p��ː��֍�p��_om�L�]�lepr�Q6~�����T���m�
�Ʒ	�ou[�B��m�>���H:xN�n��.�g��ۍլ��º�Xyy��¡�*�e�5�N�e7z���<��T��pS��f�IT��� ���"Η�h����I�.įp�����B�%��"��R�^gX��E�Eet9Hmt	짃�򡻴3�ŵ:۸��u]	�G]�r�Ͳ����]���h�b�i�Ek�)e�j�iehmtY[Z�&�j�e�;*-���ث�Z�4\�%Im����E��6m��i���V�n�Q���U�vΥB�*U���j'.�U^g��Ub��[AJ�[^6��	.�@ܲ�e��m�[R�Pmj'6�E��Ӛ���&i�ڦD�R�9fT���TE5*��6�4w4��k�W5��o:ڨ��k���j���lXZ�Җ�X��D��XW�sQQ[��m��kU[B��n<�Sq�g&�nЪf�Qm��-\�S*Q�]͢ikl����}�2�hR	Bo[2�-�y�zuҙwT9B�r�
��\�E�W��=��"����z''#?�!@�6�1�I1�G�!5{�5n;�s騁4P��k�#^t�x���X(���dHi~'Hՙ|v�>sB�G���E�����#�E��Fr�Ƕˎ�ƹ��L��)]	�-�������{O�N�'Ӑ�����0ĸ�
f}Q!\��7J+���7H;����Ǎ8�ǠXg�
*v	�>�\TRGZ�.ӄ���NaC�K.�$��7P,��i�Ț< A1�*g�u@���:�G�<5�3B�#Vmo��Te�:�����ȌƇl���+��q|��Z9L�Wy�Q���
�d^�;��{��`m��@[�"/ߝ�ݏ�Y�ץ�6�@����U'P�%��)�},�r»׼��s�08q0��X��=,���3�9��uv�]Eh�p��9�.qlȯC"h�d�%ܨ��Y_��� ���i�w�Ga00~
��H�c!GVOD��vy.�}�|79%���#�q-����������E���Uk��N��}��3W�p2�F�r�H��I�VȿQ�va5ٖs�;5���`d�Y�|�Q�z8h����¸��E��fy�r{5��`�I���)6��̶l" q�1#�8Mԙ1�;jQ��'7�1�.6}��@�l��1�܌�,GG�Vϡ]f�N���p5B�l���U���b4\��(Fip��*��Ou�	��6$t=s!D�zl�J��q�B.�ws�m��n:9; �>�<DD���
���Y�l��^u��7yʣ^����t��8��t<�V$>��.�g��|��I�j/��'�����Z{q�o���M<pA.jr'�Qbp�s^^��Jfk源�o�*Sn<꾑���㶸���kj���r����m��k?�=�uz����? | �ϐ��V7�	��j����BY�S9��n�T���jg#]�{*���,F�#hڡC��5� ��52V17W]����e����Յ<�
�>����Ӄ�._h<w�N�\��E��tԑ0�ϻ�Ȭ.6�O����E{��k�-�,�Z�\���xT�
Ѣ[4$�"��0C�g;$�L�/Ud��|���eB��`�Gc �>�
�8"�u�'��$R�v^���K��>>�ʹ��K���Gd^�5����2�s��7q�2�5=^0Y�GD�+��eDv�8i���|�4�v��(��`��.B�.A�e�Q	�}�峰���f���mF��+�"ͺK�>c�B�ָd1�y|�����4�Ĺ!�SD��8��_�s�u��::&�.tYt/:gi��fQv��r�/Vc����*���,ç�i��j �7��M��(q�˟�꯼"���n#c�*�dA�>،1��k`�o�}�0G� j��Z{�5y?{wa�����1Xv���&8�$>6垊��ރ��U��d�����+��X�,�Z1r�<�>~ڗn��S��W@���zC�(@�)/�n�]ۻ�:ɑpx�C�B�ՙQu�2-���Q�B}`G#��4�'if[�.�����
B��0/��U�ׯ�Q�I
��2ݛ��y����������^��"Ip6��#2\R���W�����N��!L�ĵ�ʫ��ԋfY��xO��l�n�W��<#a9z��fK��;��}5|����@�طQ`.�K#���Ь$���w���e��>�b���x4U�1P4`�e��zv��~[��N̾ŏ'7	��8'x+7��Y�څp��^n�)n�ԭ�vS��.�����J��Y��Ěr�m�u��'���3��;�� �L�曞�*@Qz�����T���\jN�G�՝��'���m|��C#�X�$m���Ӟ���)
�M3C���>>{�W���K�qW���7����"�h�u����Kz>�~�B�����F0s��G�b*'��C"�#�ԑ2,}i�e޾�g#D1�ﹾ5p�>���Q�X�� 5��wl��ѕ����Q�eEr�!�$"�N�h� `}��q� �]���,|���q����\C-�P�b<�����kq^�cƞ�������&E��Pc$��)�CLC�"+�:R=Tp��ik�g�r|x��ș�CDK�Q\\-5 N��"dUvu�x�����= �c���\|�*�z�̶la#�khvݘ�iFʻ�k�"��.��n�kspc�+J�ч�Gqk�}��熓۔r�ù���7p0A�o1�}i���;��w�����ƨ���\�S�+����T���tO�7
�~S���3dn�DR>��Cd^�o�sk�(�*�n�cG�z�ւ��bю�hY�Ot�<��^��\�����q����,M<1��)5�oP�7}�ƅ���)���f�O�������D:���Y��>�a�!�9�����d;�؁�2ӝ�"<3ۄ�����t%�"!�H�4�b��m�tL���s���K8�S�hFC�*A�Fʔ"I	���[@�U�[<��r$ɨ�p���4�����������ZMbC��j]_w)@�>��x����9�ͣ�KgQOD��z{��W�[�DY3�
=�L��1���PE�������U��+���	�rEz�+x���kW�5Zݙ/���Z{7��YF��t�JL����s؏ʺe����B׼�p����b�fe��+�)��������<=�g�u��}�NC�8��u\��&�!"�d"�r3����wus��	Q�C�,��d8�!G���J혇		�'39�Jv"�����'�:�
#	���8(�
��٥����QcH�.b��*�}�_"��R�g|H8v��2�{���ss��U{J��n�g�m|5�B���xV�����x�\\�}>�*a���-�(6�P�(Κc�^�{�{�T-g�5aNU����Y�� 2��o)��-�Q��
��R4Ad�0�Ϻ��\8�O�����|"�����G V��,��'��D�hIEG��ȟ3����f��7Ҥ��6�����u9����
.N��:����t��~ύ4�v7-,�Q�=Yg�`9��.��1-��_oZݰ�K��� aT�Z�!u��Ƀ�v�-�鼦��e����Ù'T���qe?��O\?��=*��n�}��*�����g�"��N���F��c0�o&�tت����	2�y��p�����GvĊ�j�Wv�[���
�}�B��:-Ӡaaq0(q�ȷM�"��:��g�q�B�r�	cOP��T(�mW�mTک~�:�va1zZ�K��]u,�TEӏrL�]�]j�1.ƣ^�@>�
�������i�WO�.G
�'��t�z�ɦ��xwB�F����l���|6g-M��Nk���5`��Qѕ�L2�'�Wu�'b׺�=�g*��jk�Cky\�F���v�&�C�!��r�Q�WV�Fh���X�
�[����G�Y�[�Pۛ��9�퇩�8������;��=�:yæ�f�ĸה� D�dg4'Q39S)�Gh�#�g:��*�9{�Qʐk"�j�x .斤�I����c��U73M�
�Z����x��)S,]��z\҃�t���G�rG�evr��M�nd�۾��"�.�i�;�m\�OOcܹ��^�&|���:yU�=����ķ{W3	�`����R,��ʡ|�r���j䦟bn�A�E��4���?<���hL��[����*� sG9:D�˕�7�.g�^���t��n��zB��H$�Ӳ�:xm�kh�!Z��-���(w`�4��_79���o#dN	�bԷ���ފތ��*[v`�&���L�Y���d�
�l����rT�쮶�S�s�,ue��x�%`�6����[�%oN.�u�*s;X#��u\�Nf�P&�)+���U�>nc��"����89���c�B�m��7��[校�9����M����o6�W�x�1��2�B8ԙ�v��4�'�@ˬ�j*q�Ԇ+��Y|sv�ģT��wf��[}tI�61��Ʈ�>��v�C��x���=e=Y7���QS)o� �V���<;^XL�I��Cн�]�e<]]*�rɮ��� �I���l��K��k~�zQ���Y��Q��llArG9<�"VK����bý�|�sU��>uK`�pІG�������z����o��p3.c��cHL�yu����p�Xф�	Q_no��d���c��>���d�����|J�ȗvw[5̀�K7#�Y��9�P��I��@HvͮF�b���M�A�
� �f�$�\-������������8����p4XS��kd�p(�^Pc�5*(i��$)m���N���նە���X5u"w��6��͚x��2�J�Gk"��ㆺ�X�rO��G]N�[\.�W�Y�2��T�8#�����N���c��3��%�K��Z=�F�0�wc?SfVl�/nv)KM��!�,��Y����Ɋ��/6|���(T��~�w��W89-�e��% 9M�/fv�ʛ�+�t�.�pv\��=���Aoa1���F^�5�����:��	pRl��Q3m݇6Y���V^��Cl�|,e<p)�D�3j���K'|U����Qyp�=�~[Y�fM�����J-C���Z�,Yn
��ڝ���27:v�]�[�#�V1���"΋z�:�56�-��}�S�)
l˴V��H�٣�6[E3�e&Y����͙N��53z�镎S�����ؓ�j�iS$��Ӫ+�*Y���`V��\u���!R��{pܮ4r�ã���K�tj���{8
��ܹ(O={s��B:Vphn%O;nbd,NGVx�Y�F�J6go`��)������ �(۱cS��qqY�2C0��o/^��1��v��#t.�rX�����mӧ����ϧM�ĚpTI�en��R�݁Y�8�9���u�aZuv���55e�7��R��Ax�nl��8P�E�ѭ�v���_�����S��ޫ��Q�ڃ\���-L���g=A���T�#��*�K-�T,�Ee��i�ZW\�4T���k2��,)7��ʔ�6&���$-*����7I�kQ����vr��������r��R�Y�)NR��v����5(�k0��֥��/���)��]��1D�yF˅�A-cLҸ�j�1SZ�*Vr��Z�
�o)D�Vrجjm�x�u�e���.��%j��ZsR5��ʜ�H�'-E9R��ZЪ�֙�m���ƍx�S�amm�/�U9��G5�Wb�&lW�]v�֜M�R����K[l^P��L/5�X�[k3�cZ9�EÎw:֏[E����E8�+�X���U֯/֪�ٵ�����矟�����79�i\)�-z�\�8�diGr��.�wN���EX��;�=�5J�&�O�f���&�.��hԅBq�V�SS����'��G�W<��D�o�=�G5n�+���I��; �]t���r���GV������6��wH\%�NP�r[����heN��ZiQ����6cFmO����=ʸ���c�|�E���pC+��5Au�ܪ��
v*w1jN�MCG�sc��OAqb�{^��{34W=@��F�8�8״]��
c�ˮU���t�0+cr�Vr=�y0kj5N��i��I�´��ղ�s����-�QY&s����u�}q\�b���L�����y�*�ά�Pa��&���ͭ�O$�c.yt�����ھ�H.�>�ow��K���b�J��$�+=yws[����xE�f�����q�X�������I�8����Ӱ��Z�EV�+�yM�/x.������x�yA�z�3ӝ4K�`kI�îW{�"�P��L�6�.q�rPv�*zҔ�WV<��Z�^���Q��0c��ȰQ޽|����dS"N�L���R+#w/�[enZm���̓�A�'z|�¶����Y���-S)c��6�6�������-��75|/�k�*���#�,iф��� ��>�
O+F��-h_�\�]�@̓���L9Y��˻��s����J��Nk[YMM�G9g~��e�g�e�(@�����<�^�U��ŖT2�H-�8V��6�ƚ��V�Mi̾�K>ީ��i�5}��Ck�k"�6�����7����z��e��4�Ͷ�P< b�������j&��Rԫ���㲆g#tnh�ȼ����s�0����}T��ތ<0��-[M$���a�dl�m��T�f�M�p�wsʹ�.�x���}N�f�ɕ[,�|����!L�ˢOC��t_�V�,Ïc۷�Ғ�E�YQ/6T��XϫB�Z�\��1bgJ�*t��{�pGTX{�V����l��/5�GD殥��.o'�CcH�	�K���M���SLH�_Gvͨ3;9�M*�������س�l�G�L�=�@|u"���-��靍qO6�^?T�y���ة-jt��q��s�1}�
	��٢(���j��sk_�s?��?��@F�'��Zڬ+=���ط7�~S�����8-5\�G�>�{$�C"jz/���嫱����.�b�7Im��9��'&c0WvZ�Of���Pއ�.��Y6Vr��a��7��n�9�a�C���^E�M{T)X^j�up�L*R�^(�7F[j����L��bV��D����::�%&iږT���)�3����� .�{�/fFWo��T�����}^���W�*�A�9^�g;�@PY��x���꼑L\�c5�����F_n�rV�B�D�ѕt��u�H孂˺ϴ�5nP60�w��B/^z]�<�u���}H�D�Zu-�zB�(��Y���$��U}Y�YͦD}�,NR�by'��tl��s�r��y����Ќ�Y�͚9<�o�@g�n��vg&ْ�1m�2����3�^>}�8-�-ZW'���n������-��B@�!��z�w\�ֳ̫7չ�p��1�<�
����E{Vm��/zzf�o�3!�\�S���	�'kr�js�y$�ig�t��Z�z��2����kicv3��|)��p�MoEe�]{�Ƈ�X���	�jG�����/���k�F��^uôvp����*����}^S�C�C�Y��ԽQD��o�(�d߶&%�-<+��f��e�3y��馄d�wrm��oaʹk�Y�"�^8�KD ���&�$e�n��M9�~�����)����JVK*��� i�^j��o܅��G�?d�oc��Mz��-HL���E�4���Y��=no.�_>����nhc�_Q�^w��|��_>���9��)�m#!3�ku��m�U�Pʱ7O,f�����p��Yk��N�/��7��^��
��s��m{pMo*%��19b�*��P/<������r���3�Hڤo�Y���ɎI<�0���]>�Ys��>��+h#���ȟqo�]o����IfO2z<��-	�|�٧��Z��Y�ʈ���.�jE٭��Qw{�ʛ�7�uxz���\���nq��Y{��̥�nщ�T��m	]��p<��_U_l.{�G�|��c��Ӽ��U�)��u�MK�i�����ᾁ�l[�w���N��KU3%k��O�
�Ƒ���.��aź������Y�L yX*�Q�e)7H��xZ~�S�VU����n���P�Gz_0�+���{̉���58٥&�7�gBu"��u�������<��;���ױ�d���N��Wz��%�ݞ0E�8���T�ż��.�zE\��7:j{��:b�l.�T����»3�4�o�,�u6�{��\UҌ�����V�*}�Ge��3�"L�MM�GV�wy���ϖ���N\�����Kf��{����Θ�$ǫ"�O�0�����n�6�Bm,�f��r.���އ�����V�=Z��B�X��:�c+[�!�U�D�y�W<7��=�s˛DLDQ�:Z��tNu�>n1z��/e�q�[*����:�e��KyLf�������oz�~%E�8�q��Y��~s��ckHn�k���g7�p�ku��J[��;ynD��?�W�| K�	c��ˡ<߲�+�����@��]b��{f��o��@��ȆG
�V��>-�LoC]�����^6��cz�>)h��E��kQ�dHnz.M���a��QK�2�U����KjS���u��Akݮ������Z�rh��"�Tꃆ�;�%Jz���p����,�[�,s'�f���J�+�U����*�7�>n]F�AJ��ku��N��|��N�Ƭ�v��5���N���{�p�p!���:�pS�}r�AE^�|����Y���>���M�Yb��5�d�"ln?��ֺB����h��;<f�V��Gc�[j�q��wU�Kg8�!���T�u�(m%s=�����*�����fכپ�t�%O]�[ʼ��*�e�c���B����>~tU��B�Q�����m�|�-����<�YN�;7.��+z�|���x�U��HIW�8D���z���z氉;�sW��-J��ף�L;m�x�|�HV�]t�͔��*O��C����3�t�|���,m���~�a�n�n��^�R�8v���_8��'b�Sl͝j�mE�5�&��d�N��=��z;o�V{$����Dm-e����=D�b֧���+����G
j�:��QOw\���F��
�E�y��9*�S����S�ԭ&���wH��60O�]Ej�"+�����K'��F��V}K-�l+4�;�K�&(��n&��չ���-�-G�N(9�a=�w����A��bo���7�QCr3���kdU��ev�K���FKu�7Fj~�OZ���zV>�yV[����ė�8g�xbvB+f���s��=��/%n/]�j^��7Z��L�5�tp�h3�;���{�l{h��kO�n�Z���2�1�[�{��8=.��{��5���1�G��f�-�zz#�b`x��J�R�Z�f��S��%k���I�VC8fM}���Mҽo�h����ۣ���׭���T�瓡�`шۂN�C�ү~����۽v�fn�xɵ�/���se�E��L�
���^�`�Y�\�c�b�MN�bh2���`S����oK��hEȪ��oL�L�u��+9�2s]�i�C*C.S{S6�QH^Z�$v\;tWP:�7p��y�s�Y�ڭ��F�� :�1a�L���I�}����� ���j�]fZ����&��6�r����{P�^�5fXΩ�̦�c�U35b$&���p*;yԴ;�e���ھ����T,����f�o���j�j��ݸw���G�j.�'1,��႔�W�LWJ�S�p�yw����9&F�S��i�7��cndM�m�8%F��������Tr+H����n۳>��(t����9Wwx�Enw}y(8f[ޒ�vom�qKy�wO��H�+:�OY�`9����lL�=����c���{�-��̱8���)�����YY}�3���CS����U��\�N=Զ����mm�W56y�Ѐ�C��;�Ҡ�(kȱU���X���`��}�u��S9Pt-���Eu�k�+��#�F���V��`ͦH`9�*9ڥ8�����%��
W��M�c�s엷�1�&u�R�p=�ۜ~��a�X^��1^W���@��r��zÅ��5o7�n�vH:�Vۣj�Jp�7"���+!���S1p����.+�$�@���������v�ǌ��D�.�Ʈ��WeV"Nq7Q�J����r�/�ݎ�J����u�ㄥ�%K� �0�Ǔ+�>�:C�(֋V��J+��u��|J
�ǚ�9lc��Ί�0�WsW��\�mqUU�UQ3fJ��G�
Q�ECYb��m�X%J�B�XԢ^lq��)fyo8ڣl�$TQV�n���Ӎfi�Qc
�fj�Z�TDU���;6�g�&jnm5F�Ъ�Palڶ��m�љ*��%L�yj0�50QE�elQjڛZ��U��cm��0຺�J6�	�r�\keŕb'����U��]y�3m�V�><sD�����* �:Ɲ5��2��63�m�r��QKj<�lJ�sTQ���5�]9I�2�n�y�&E�q0��Tk)klG�涖T�����/[�iZ"^Q�<g9c�#Z��P颂/-��V�T�g�x�X�UF���ѡC,	��� �{=u;6�Y����kM��{%�c�WZ�K�׹�g���m�3ߗK�=�O���r�"ϴ7%]&f������:'�н�)q�RgY��Z/3���o���{�K٥�e֬��<�Q��V��$ۋlq|6��'t�o�E�\i����y�~ê�@��9<gy�
�Y�5�S�yY}��K�7͡}�o��غ�aw����O���rkX-�|�w�X�ў��.ɸ�5k5��+��Rއ�{60!�+L������M�4�2�o���G��藛'������D����ӣ6��0p�#"��ڨ�3.��{$�w���6�f
���Zvu鋩��7bwj�|:��㊗;�c
HfgWN�9�q039��7oz�W-v.���*�.M�w���������w"�SCf�km.s'Km:�b#B.�ĳ�v��ŭƋ�;������۶,�P���(L���v=5fmo��%G���L��j>�X;�}�:#\Q�OL!���F�OR_m2sU���x���J5��Z����uj������+r�h�nh%��\�q[IF\��:�[a�q��W�1�����T��t���=2y�M>�Ķ��	+���7}\��u:Ҩ�d��}���[y���9�O%�Q�{��)��.9�G$t��^`�T��f�q����;��i>�/���{�B�nF�G�� �&ƟvE����9q�S�L������ ʎ�f����:C�0���zAx��(�wL�i�����3zm�t����(�0�YwkV��͆D�5�����J��d�)���}�f�mц�v���I������#4�v�f�,P|��;Ӕ�8�nM6�\b��]��C��[�H�h�K�ӵ".�7��f�ē��me<�9���1+��=��N�B�Ws=ܳ���/�b�n����@����PT�I����������h>�<w���=p3R�mZ��V'+˪��Z�i�I,����G�i�k��[��>ҳA�G�l{�7�v�z{ݳ�r�7�.���i�����KH���]��	b�B��)�aRZ
¤5��la��=m=���F���m���t�^�H��d�+�5}�xY�Z�sG�n��p�F]��r��⃢g�˼ޜ�V핯^>��V�dp�ܛQ���v��g�~ɘ��ɝ���~�c{e���!ٝI�)��\�y"����j�J���]`�陻��k~E��툢��g����,�����Wf4����?��:4��9��N����,�I��-(�ԝ�U�aDS�s��E�Y�.q���V׊ت=�C��{�q�L�L�uV,���9����1�o���F�b(�i�p�+6x�w-��P�Ve�!��e:��{�����GW�&%{U�����Q��j�T�,�$(�c�gN��U�8F:�p�Ζ�����ʵӁ����l��F�I�V��"�u�M�_W/���}��q5��{&���鷣��^r/�B�f��jV���CS��	]͛sIe[��y�}����b�He�1u��
�Sf�f���6]��W=uO>wҪ�UtX��Ax;=�Wy��7=��L�9��ކ&���,Y��H�47�Qo��\����+A�Z�rǴ�+�3����'o��8����v���^���1�'㊳�jM�>�xsc�%4���ݯL����#��i�
�_z����U��{�����g�}.bt[�Lo۹��V{�WO4/�ط�Km�^���1t���d�˺|7��a�VT�@G��U�v���&]yIt��)o	��0t������V0� ���8p'j*%+Bo�y=\��x{�U>mWg۝>�ʡ7Ж��@C���y5S6��o��T��ӆq|,�e}�L }{���1S�1S�����f�4�7+7����Ux:��VSi&�l���GeO�j}mrn�u���S�]���yo��*|y�ݝ�=3�8��_1����W�H'��U�~��r
ݝ��	����)��ϧ�1Y�B+,�P���{�7z��٫�)�g3]u�5ҧԠ�]���6 ]��떶D1�.UFU�Z�����z�39H3�?7�7�[�Jϰ�B�I�_t�R7��\g:˖F�[���zPFY��*��JQ�瞩K���}�.�<�A��;'Q�eXL�������d�Mǽ�����V��J�źȬ �E������Q��f7�[��� ��/$hK��Jl�c�\��]�n��ڕ��ȋ��2��|�=�w$��k�U�S����;�q�(�d���w%�0�m�{�9����Lps?Hr��#�:~ڙS4�K��Ԉ�U�'�Ԧ��WJ�m-��(#;n�LX�����|���ȇ��g�J��d�ާ]�SM,ۮz��V��4�wP���Lͩ'^x��t^U_[���N�0+c7Ҕ����n�lnK�3���u�C���u�Č�'G�H3[��Z�r�9SGe��aWRvXE�Y�k�
.���I	K�i��B���1_�iˮjX�6���@c�����:ׯ1V*�X���'#�;Ź�O^)��v7¢����Ͷ[�6�8�t�֠p�ғ��W��ِ�~��;?��6w�{F.V�x��k-F��'��o*����B�j���Z�jm�Wj��^�5�bHm���=�
�����;�bO,k��Lս�Ҳ��P���B������&��:���]N��G�W�X^��B�5"߰�W�:���C��ܬ�ބ2���&f�&灗7ջEh}�{��b��6�_g6�Z��n�;�Jڕ�����Rs�uS9ɵ���kH�ܬ��Lf��{�}�S�ua��n]��{�l*��t���xSP�Ś�����3�3���VփN`:�Q֨Pg�I�= ��l������; �3vTRnФ8��ի�:����h�D�A٩�r{U�,����;����5I��L��_H<��0m�+6%���Y��O;�sz.h%ڴ�����3c�WHکr����xı�=I�yWJ.�6�$���1Kխ2u�X�
R��[�C��5.�R���/�{���/�]�x&��JnУ�̣Y�S�4҉%��=1[^����_JW��s�7�-�Jl�V�kmI,V����V<�2��S�[4�pG+e�*�@R������4�nZ5OSl�˞�̹8�e�[�;H�R9b��c쮭&��wa\���W/kՊm�[�UrƉ��&q�j���c�^�۽{V���c�������'�`i�!v1��V;���G�{[�I�l'�ވ�#V,wڼ]�u%�]X+:�t�mE7�r1%5�c5ܐ9e����T����5]��qQ���,����t�SZ�z1�t�F�4��nG
ckU�7ve(�:���U��9���^=�{'����KyFb�����7�3�N��1m�C�}��Wu��	ު{�)�'_[��oK[�P8X�z����jD8�z^��nS܇�!خ�ۨ�b��n6!�p���+�뵎�����䣶��B��15mri���� �l���Hb�X�Q��2�|grwf�L/�q���p�	-��L�'�v�U�uS��^���W�7S��dE�ͬ��m�En6����%>p��������ۄ_X7�~��LiAۄ�t(�&�:���:��f�'뮥VGesP:W�mꜱ;��W]��)�ޑY���h��v9QLTF�<�����/���}b"�J��:��dw�7`ۗ��o;k9����HG�+G�h����V3�c��&*��t�,]��s�S@�s5`��%e���qy���n�p]�y��_g�غǨ���c������2�1�5�ޗ��<Ɍ9X �X�,����x��u �K"�chb�jC�ݙr�����H���n*�u����w�������õ\pr�T@	\�ȓR�,+�2��:�ؒ�"l5��j���2kB���Y4�cm��w��(6�'`�'����8eg��^�is2 ���$/��WGhIݏy�h��w��ew�b#��т�U-�#=�b#}2[�}�:)P���5���a&��O��I=����	�&mn%�2��4X����+�<V��ǫ��
.<�r^үq*{6�pX�+�4w4��)pN����K:j�Z�����6m�x3.�=�í��̽7v�r�iZ�]oRL"��~��� :�V��t')�w+�qW�ʒ���r;�KW5L�VXsJx6M] �ܤo���T�mǢ��&�XlD�5��Y��S{h�u����Ϗk��GR7`6�.3Em�s�����^��eD��/�16r8�!�U���*3�5r����L·k7/2� �Sl���u���.��X��}�P|�N��eArn`:�w�t���E]�:�:��9�W	�Kj�BH���//���]FK��Y�rned���� �z6�%ܻ��D�h�}&>9���ސή���˕�}.>��Z�Ic�r��W\v�S$v�\�������{�|$I0 D"��R�E��UP�X���,c���ea��R�*!hQ嫛i**�L­�t\�i�Z��X�mm-V����sku9���J5��"*"�i֣iӞsdQ9̡����n^p�R�X�ګ85ұh�8�喵W��y�����R��*�z�b���ʋX#�ޛ�Ӗ���U9��T5*�#ĤxԩDFjs�u�W�[o6uJ	�U`��+QPm��ԋ��V��V۶��t̡���c9M�6Ӎ��J�Ţ�����QS�3�����[F%B��!�U����[,T�Ҷқdj�Af�5�뮵���S�%Zδ���Ӧ��n�eMS��Ԫ�K
-��*��6�V+�c*�(�֋�L�a�n� U
�+�⏝m{ko�*���it�Ɵ#��&+������Kf�GvTle_u%��=�WُSu���y���k�9��b���T����i�NI�o��u�;�Z�5��-�٢f1�^��qa���UF_�R�gt�����nwq��SwE�U��KOo��w"�].7�r�'Y[�.m�2䬍�/IG�ݝ�I�3�d�Y�oDp���c�E�
��=]Y���"�H_e�󿧽�!C}���bE�Y)���I���1c{��	\zH�x�h��k�i�C��؉��+Y=����>�q��"g�/��0�@�e��-��\�S��2�-��I�LX��,_)���SAE޻�A_��Q�񎣲�[[.�c��.��j�qV0��1���n=����ݞ�q6+5�dnP�l�?�}�8�=� ;_����^MP�X��2�}mf����χ(Z���iJToj�)j�r&�s#ԬbFx���%�魨S\�s]4�Տ7�C��V��M�B�O%�Yz����V(�gvw{�>ɇE7w�y�
2�ʾ|�FZ���6��B�_��j���2�3;ZN#l�b�ZsbE�F���\�
���u���ҝ���Us��D�8E��fȣ���I�غg��eN�G}���Պ=u�n�e�'kL��ܧ������"�]j/ss�lPF��SH8��ۘ)ȸ)^�z�eݢD�vt�W�ժ:��s�vD���C*&zK���ε�ܬ�0�a�%�� �uk8����<�TŐ�:�N[�[ˑ���L���/_e�`yS��(��󪖷yŶ9��'�������4r�=5�
�Zy)�k�ƾ>��B,�(��<�<6��I��$Ǽ�}��������`����v��SU�X��cz���6w ��}{��~��.dP�އ�!-FlV�Pncg[���6�nz�r�<#َ"��f��nMbM(�D9�&���NT�oF�G���W�Z�L�-MDsY��u]�&��X��b\��fa��8�qo9u<Z�0kloUM��J�[ǍVTK|H=��b��$������Yw{�Π:P��N�6�aY��qJ�{O�ڛ��S��j��|�|d]8�Qt��n�"LR9e(����ߖ�v�;���%�⌍����P��n�t|��{Kέ�rH��&*y5�R���ȼ�x��g��ZUr9�y6NE9����A)3����y�]/W�+T:yż�ܱ�#�WWݖ�i�/���SJ��8`h�{]�Ej��S�\�rSt�u:GE�!��M)��UC*ٽ֓�/1H��ܭ�� o�=�y�s9�m�R���N��-���-����eLn��Vf�rH���o[��(�[A�9@�㖍��E��A1��K�����fT��y�6a��cՂ�8j�J����� qtr�>ǣ�=6KҲǓ��eg�a�6�U��V�7:R�i���%���=o�O��1:��<��A0�N����n>nI�۹_�X)�V6?3A��;]�J���4�#�>Q�X4���3=��=��'�� J������A�⍌w�&jC�hIw1�U�-�)k3'x�Z��)5�_#^�󞖮���9�ٽ��ޡGf��,�6��q�ŝ5O9""�.d��.�*���ӧ�C���t�"F��(��^������S��h���SM�'k.v� uG��iY���ږ����w�OYg�94]��1�e�#.��VK΅�p����Ɍ/r�.�F��G({����!/��;��FL�\4x��!�yxU��"wԳ���؆���>�/>�Pʜ���K�B�ys���[�3����N�J}����1���H��tǷV�����*/��mW�T�HhŦ�fr�+50;�dJ:^���N���EP�}�-J5y]��$��வҶQn�W�0�^����q�[��[���ŝ	Q�pZ^�:��W�Q�u
`(4Ӟ���2��k�
*�ͥ����5.=�)\;���+�2�g�OMx*��oP��>Ӄc'�.�2m6��b�ӳ=�к�I���P�׋��7=y��ViS3)&3��R23�Je�U-�v�X��$㣌77���9K�;�����٣^y]X)jVG`��}w5�Rg�t���hY�|F�JeR��lgr�N䚷�Wv�5l���l0d�VEv1b�8��kx�e�d���̒c�.��I��6}O3C��l�v�T9�=�ɚ�v��������r|ϟ���3�20�؟2�Պ�F�+��T�q���T�>kk��wӢRc7>�ٖ����A�F3�[[tz^�����y��w5X����͌��魘ZV>��rv�v�f-����N��<�A͟/NuU]L�����i�L�.��z�w����6��˓t��smU��Ϸ���HY�t_v�oRNGs�@�s4���C�"�$VaհGyoY��|׹u����B�ٮt�&����~�`)���]/��ǈt�nY��̗u��
�N�"����%�PC�;Z|��n]3Q�e�դނ�T�j�%��sD�I6V�#q[(�i��g9�fl�s9=14��NL�oP�E�(��+5?�n}�ot��fwv��h���d�{���dF�V�⻨���ξخ��Y*�����Z?�)3�VP��<%`G�oK���i��g�]sFzUt`�/F9�u7X�"Jx{�[5�^l���糱n���u��o��e%p��(t�l��"�kWͣ9���˒�AФ���	�|����''����E�+��K��|}���X��ơ����J��q�����*�Z)�V��X޹��^�(���^e�.��k4?�R�%��isd�Mg1��jٗ�yڗ�P�n���N����}�扮�ϭ��o��c�YLɤ��4eq�i�y'״���7�4��%��m�l(��Z-ec��P*w.H4r�V��>c<��V��T��1Me����hކ�ٲC>� ��nf�of˸"�=���R�ps}n�6���6ѧ'�k+vu�o;�ؽ(Fp?/L2՚Zڡ�ʍ{*��e]���L��X�X�މ�܈�{��Y؇dq�}��g'�V~o�k�ʵ��3��b��:��[�!��rLR�I�p��sV������I��Z���"�@��"C������io�%��-i%��Iv�[ ��N��"�;`�F��A�,\V^La���̻�@�5q�:�:,��nV��׽Q�}�e�_
��otb�	]OV�ʌ춲iA�atZ�͚$'�������.�uR��%���yP��BR���g{Ȩ��J�<�V2��:�.�jS��ŗ^�\���joo�wYT���T�J�,V�Wʵ�y��@���ݎ�'-+��6�%.:�OJw�NS�Oib��R{"'е�ֺ�(k�i��8�����۱���]!P�K�;������D��4��F����6H�ڞ-����oFL�Iu������.+�����4s�F����c��}�:����i�,U��@WgV&�ת�M�z���$���T�]b$�`�̵{��۝�7Hxk`���%�|�������|!��=Z�է�W��s]s�jSs"67��|eYo��`v�],^3�1LVg,'���]��wH��F��r�ۛՈO�Q�Y��J��c��Ϟ���U�n&h��a�^`���@���490��B/~����w:<.Fyr�v�3�HทY�\�kU�.��/)�r��oI�����譩�$�1ӳm�B���-��&�JݾT�'�76�0������8J,��a��*ɕNM�M���ZM���Nw�(�EmUԷ:�P�Z�^gb��;H�d�=]��nS�X�ܙX3��5Y���K��M�m�^�a�Gn(�Y;ky�S�A\Y��/kob��4�f�Y4J�ӈ]�l-��;�hu��m_���k*�Qqd՛�q��S�q:�.�Y�&>6F�,��g%��X�;s┲m�;�3�R��릚�M�� ;�fAxGL���
�r��|��b�JoF��8"��;�q���(�:���>��o6��0�ǄD%utHE�G>�����Je�ܣB\�*�ZS��Γ�/�{��4�����(�%;P%&ܵL�r@�U�Xw�47
	~X�R�~e0vδj�LY�7 6ս�4�ve3�#l��+�sc�.��-�6i�.z[+hlr�Rn��/�I�Y[a%H�ɼ��9`uwg]�-�h%[̚=4�@��4s�Ē��)H�R�Z�Q$�VU.eL��Օ���tv�����ջ��sVE׬`1n-B���f�׷���u�>��ҙ�/74	C]f�;F�kK�"�R\9s�.k�3ox��v�R��8w	�3�;��FN%�ūD,Z�
�Ib��C��]r�7*aY��e�i���fE�L��jX��il�îY�"(T����؉mE����Kig-�Rq���W�e7-U"��ı+o.3b�-E�0ylb,u�#ͅ���u���*<�.EE�[K�W�.��r<���Md.��LW%x�UF9)�VҚ�\��Yuk�s�mT��p��nl]��#�Eٓ
���9��ԭ��eMK���Em*ƣg5u(q�[b����Z�kUq���(]e4b<��Db1u��lT]���k����X/�Ƃ�4ԧ-S��lNR��A��nj�m�Q�I��YTVs�0���D�Do,��S
F1�-)��Rң���險��AEbb����]Y��k%V�H%�K`�*�#+9�N5�Q��9B��������?�Mxo���"/W3�y>@��Wa=:R�C�(9�HهQ�"�5�trc���9�{Ƽ�Q��Ww�l���Ov��"]q�27H��l���6LT�0�R}Ȇ6��˶�UT�o}�,��`�sz�3R1��Q6^�y�o���7ۯ��ϼ�2�����Q� 5�.����-�oFQ��V{ӓѰ:]W)���#����雫�ML�����"vu&ZthV��s�&���\��Ź�[ːk��&�[�"�{�ECA��,�^��z����YWQY4�71���Y0�}�+fؔ�O	ST�.Fi;�s����sv�K��n:�ӁB�V��-��}�ٵ�K��ɍ�<|h:vr�Ф�ms2���q;`�:��8�T��;��47E�]�"k�rS���"Խ����I��F���1�V��u�Kk-6��Db�v�ίs����֪�US�Ks���P�3*�gݪ缦<[R���[�<�_�}r���qٜx=踩b䫀�*���{�x���Z镌`��6y�iu�a`�6���m��iKB�[��b���b�F���q��wI����|���탩+�u��V倞�a�v����==�j*i���p�

8=�:34�A�;�^ӷV{�6�1���I�5��h�-=>z%��9�0RQ�6�����c�ޢ��@�3Φ{�V�.�� �b��F��A�Mߔsh����Mਯ�ϥ��ß9���/�N�|\�n.���ιܳ�r]WD��ɶz�<QH-`�՟+��7���l���#9*s�-��ܳ�]e��Um%9[�=�Ѣ�
�AP���$������)y�����:.�.E��b(ԛ�ֶ�*ɺ�����ў�m�)��z���`��O_�.i�gz�j�q�#��e�i/�Zn<�]'6m���QW�m���7������T`5a`q�P�K�ԧ�"ʩ�ڑ5}ؓ�~�-�3`�y�Gh�i�7;j��T��������j+7���i�qjW�rժ��ѻR�"^Vͫq��t�3�"���ؖ�D�ȴ>jV���&�eh�;D����6����E�n�Z׻km�[��&�B�J�渇��ܥ�v2��ϨR���@��o��[�7�|�N:�W�v)4n�&��ۇ7Z~q�@���n���*ӏ+�y��#(������lk�zdR)�����['y�9�s+IDk���k�|���/$_Z�.äv%*.Nݾnt�����k%v�3ʝ�������{�jm��sg_e�e�6�������&�C�7���hx��ی
C�X����̥����6|�����n~���_}=�*�
a��{/%-m����g=�+�]�IV�f��{�{dU�"��Ab�wU�d��:�^q{Ӟ� &��{���{05#�軰��%v+�9oA���ޫz1[Vc�΋��|��X��7йY���]⇣�'���E�6k�u���R�I�:�Իٚ,n�Qet�!W�S��f��|���-��t7~L��60���3�E�eg&���cF͎oGk��A�"���9�S��\��d5n�kF���}Ű�z#Un��-_%4�M�����j/f�;9�j#�$^��f���u��Y�(쎅��p�y�=[�I|r��5x����IM;��9V}���n�?K�5�t��\��e9;:��������SKΩ�R�{&�k��LX�s�WlAPɡG�Z	�7���(<�*�q����q6���S������Uk	[]먚���.V��+�Ʒ,q�Q�_L�.N9g6����\���3�a9#p��ӽ=����vy~��'b|˧[�lƷ�4�_.P5��m�D>[B���knv���j�6�V�t!����/�yj�������D�rgg���Zh����gV\^��`�U�u6�4n�s��ɴ�k�<�~�f�|�j~sY�qa��+�6���8=4�w��'����d[]�m�ǅ���`�L�gwRP��"yO�\�KC��9����uy�PiAb��<tG�.l���6�d�9�zu��L��y�;7TMH	�dئ�,L��un�匱���:��Ԙ��7�+f�����֓�H��jo/,�D3�O�j����o+���8ٷ/v1�k������Sf���HV�'dVu��@f8���[��(�:.��M)w����d����K�<b�{��?Y%e�F�4�7�޺���u�j���0w�I	t��: f���iu��O��˜�MҶ')�U���W��UA3G�=��!�� V����ʷZ�<������Bͧ4��fK�yIA�gRY�QO�н�I�q֝���%����p�4-�w,d&����9S	�]6���#�^	�C����>�����1���Tg�?t�U쭘r�cOy����Ԏ�����􎑾m#��7Ox�p.<���.�4Ww�h;�t�cw�x�4o��z�.([���ع	0IFs;�S�^a����gN���9���˘���I�$���ޢo��偵k'%�i7��5��3Fy>+�R��#������:�qz��j�o���nZ���|�l~��eT��t�<�஖
��S����V4�h��3}��8F u)��86(k��|�1Pe���r���#w�F���A���ٵ����ê��,�;�D^�잛��t<�[�K�$�c�7�7���i�g]wN*[�Ƃ���ެ ����~ٹ�t,-�E%����|%Ut�w���%ky<��V��ί<�ҥTx̄q�Ưh���������b靻 ]����؝F,��������rR�.mB��}�7���GL4�喥+}���Ø�=rnq�p;t��7��g97��7���A��eQz��-��S<W�~�J3�u��'e^���D���yP�f�����9G
�oJ���.T�}g�گ���3k�S�|�{�ʎ��nW5�G�EWA��;�6a�oW��P�G���B�m��9�su36�k�����C�*��<��T�l厞i��U���H-�/z4X��Y��L锳;����4O�_*����p��΄����s7r8��@�̤�b�':���o��;1�8���eM=�g���bo>V_,k.�PO8�(NtΣeڮ�����bj�E���0�<J��׳2�WW<:��+�O9v��0�3
6SL��pX=,���Sg/_t�������͹.��,u|�;��%UMRn��(�5�v��{��.�H2+G/r���y�9�3
�V����u��� ��Z�4�}��:�L�T;V�)�5��ʾ��*k��P���m�m��˒"M:��yz�]��s����[-˯J��'>�#���|�ꆲ#^�Wo�����g�+t��p:�+<�uV��+o�r�Zse��J�}�pb�P�u����zj��bh�m���nU���O<�ہ���"����s�Ѷ�i�e���w��,��Y���;�L�@�"�ok�LY�$�Zpwn����ç&�e�n�����7`5�*u��x�'��pq�zp[��v���"�%:j*�8�[ǵ�^G��Uw]mv��
�f]��o
O��Q oW�O7a���`rF���V�z��%l2w�ۂa�u�e;���(�E\z����ͽ�oe,�yc9z���(#�#����p��a�j�	�lJs�`���`)��,����e�H��I�r�(��
�,��QV�U�(ތۈV��ζ�x�O3��"�FF�v��ܗ}���K���+;vi��M�6���5�$�+�_TIμ*'[nŽ��f${� |�LB�n�w׎I�͓,�z��t*H�uŞ�+�!�I.n��v�-�u�@Ey��Z�3��0Q�8cmn)��9��-��7��e��ë(�u���ïE��������F�u7|6������<[/e�e�K���p�zt5��ަ��;vL89YMRKud-e�2N��u�Kb��:��}������Z�E83��u!�Eo "Ɨm����5�u*��/Vh�:����R�D��8;��D�E/Hͽ�ӄ��(/p�Y��N�Q7����b�o`�v0b� M]رԶ_W4e$Mv΂�n7#�p�\$θ�VA	�2����bj8xf�"�9[ur�6�qsJ]�G+�Kՠ/�Rԕ,�zed��U�{�k�:%� ��ibXun8pCQ��5m [
K7 j�k�#\rv��K�Bw�ʷ8�U��J癄
����=FQ|�ϴ�lTEv��H-��w���-\�uZt�KP�z��(�a�������W/��x3#�ͷJ�EW,�wa7���u���׷hM��cw��.ʗ����F�{Нt�=X�,�5�lCr��:��N^G�6Jj��9��=���Wie��=C��QDX�KR�-P�͢��m�˵���--y�`�TRҖ�EUE"����]K�U���26�墜j��iU����W%yj:�ҏ,ڱ���<�r��D-�*(��[Em��Qɒ�v�TȼC<x�U*�W5^5J�GR�xi�׎E"�h���F� �:�*4]ӞN)�V�xʘ�0Ug�<K��q�jZ�ګj���ۖN"r�u3���ݒ�ǉ�q�A�� ݩ�����"��D�)yx񜊍F�msE�yn��t�kmNn�x�R�kiJ��b��lx�@ ��!��?��t�"���w�M���Sx��m�^H��y��6�L����1���TRe_~�l�o�b��ۆ��;�'#�{���+2�v��61����|.i%��Ƶ�M���R�E��x����nV"���fVe�NgBb6����#%I�d�=����k�����5��x軧�4��==!�l�c���4���;E��b�'N(V )���#GX78���f��#$��t-t���t��'�wU����f?r�ߦv��CD�r�^����5pXDh&)�sƎM�Z�����K9'Y5���pEf��9�D�{.Gu���r���Gay
�7�b�A�X.qK�sv�k�{�[,�j�Cx�X����oQe,BR�2�)+�]�}��N�I�GU��.�8G���4�,f=�ɣա�{�iC�Uң�!ς�Ǯ��-�>%��+7����tRѾj�:/Uzo�l2�Տ�N%ۓ��{1��F49ޜ矯펉�xW{&���ζ�a2n7�`q�9�7,<~��zM�L-�լ���37+]�%��ڀ��|����U���b���m�{@�lw!w�s`�ٲGhb1;]
I�X��Orf�K�X�E�#4��VV�ˠ����jy�3>��|�>�Ԭb���hCS�x�"X�Pj�皚vxp�Y�7:����V�Oێ)Z��%�

�bYl�_ix[�и���֊�Z�8Z�N�z5�AY�C��YWq�Z{��T+x�c�e.3rۂn��`d�^viZ�E)~[�9�񬛳{�9Q��#	���pG�Ƒ~u�B�n@�6��wuO;orKG��;*���L_$n^R�L�p}�o5����.s{$V��I���!RW���{G�{Zw��UУ�o{=;��ͤ`HkL��NoH��Y����)c+��{n����J.8':K>]/o����Sr�כ�����qr��B�߰!���+���������u����#���� q^W��p�y1���V���~���m#J�r��q��������Zo���}:m�xK�q9��:`Y��l�b���	{/[;���ˡ��5��Q}���-;��M����h�=6�N�9�����&j�{!�[ܤ��a�<�jd,pݦ��E�ޥup�^wr���5�\Ȱۡ���Q*nr6/k[|�!�t9�f�Sj��F!���"sn����{o
���D�mM9SV�Xsq�9�ҟs�!��/��}8R����x�4�����[�멘r]&�W�&E�]1]��9I�&��˫�����Ey�`�W5�Ր�y~�!y�Ti�/Q�S�W�^�M�X<���Z$��x�k��Gޠm.�y}��r�O>D�"3f�Mn��ⶓ`����8U������N�ޥd���U]�y�gU��f����ޥځ�ƫ���F��؜�D�H�c@���Fw]�+�]�K�6�[�+��V>� �����C��jm�j93���/kV]*���y���f�����ٞ*gy�;5|pa]�/� ۀ��rT��VL]�OH�*��N���"��.s�c�Ԍ���t��m��6�g9>�ط�3]5i��8m1*z�wu�MQ���;����J�\ϩ$��,���u(�q@��y�=��i�7*�2�ms�����l���g'����ƪ�i��6J�kP��+Q�{D]>�pt6mg=����w�غ��*��倲���hyz��<y���TR9�c����_<8�Lйh_S0奎��i®`����Ķc�4}iԻU�xB���s�C�	�)',��䂷ժn�2N�q*�b�
�x�.�qԼ����5���Z'Es�Yז���4i^�q�vEt�$ErW<E�dV�)4͕�Uu�/q�/��t����p%�g��;%EA�),{ӕ�ٳӖy��*5ڨx�Uڍi�Yn)� Ξ����Ⱦv�Fl^�Lw_[i	�!��;�R�e.�S#u���F�n����rt�l�.A��}zv�Jw�"���n#i�k}^��M���-�լ���ܲ�r��P�v�Y��G�iц.�+�a�xkΟ�PYB�X�j�_9�^�7%��=�(�C׳L6�-yޯ0:����HIQ^>�Ԏ����M)�mr��q�1d#��NX���tY2�g*s����%"���;C�9�/c6,u���P��K)f��f�7ݬt�DZ����X/k�����Np���eI�mk���KN&w�j-����9m���=��F�'h��%�������_���n�<kv]��d��OY��I�*��n��at�3�JE7\*�cvDUus�P�����,{[]M*�G���ü^��o�ӪW��V�/�Zכ-�T����NF�ҧ���[h	�Խs�`/��KD׳��1n�8���`ܩX�V�{��\o�(q7N���5��As��
�,��7�N�~��7-�K_a�C�s�ٞ�˹M���s�4���qK�.�'�Y"�*�[�C#-M��N�=g����'%�n�w�ѹ�<U�:�_�'�^��x��?gT��B�ч��tt�8[#E;�o39�8�6]�k7����̆r��LN�2k1!���l[^��-�UI0������Ù��F�����|i�ރ��t&P��O[��]k��t89�a�C��B���9�R������r�]��e\5#�n�Q�R,i87:�̄�2����!�����r0G���Wo�J>���੺|�+����3L;�9��{�0��{Ջ���×v0�')p�5�M��v0&
L�	�@X�ޔs.ǜ��r΃�'y�Oz���a����o�|���g�I�o�M��`dlè�t�ݽ�W���w�J��5lu?��7��]�����&DV��e��A�[�d�pAݎ{{�,��G���j��v-Θ��'�s.D j��.Z��3W�Ђ+Vx�u��oF7Kܻ�қ�x���:����ց\;r뱩�%�.�ԲWf���� �	�*o;UZi�٫7���}��M�7��˩�M����֦-��x�>R�t����m��3ܞ4�8���doHnZ�i�ǀ�&�8G,�o$�w�0�XøD��ݵ}�>��=���$�q�h38{�e���,�-����4�/�E��ڷ��٭�ɺ#�I}�P@t<��=T�eA�Ѻ�5�]�.IC��Q��K�a��os^�2�)bT�펱���&�hV�yܮ�v5g�c���HQ�Cb*�;�����nh���:3�R|�e*;�h����Zp_O'�|��wƢ�V/x��,
��^i����[�%�n�a���d�Λ�۷*3*�q�8�<{C������T���M���K~�c��L�f����ٵ<�J'y�4y��Ǻ�fhU׹{�4f;[&��;�s�L�]��ę�J�H�ﺊ�BY/�,��	C�|q�%�[*V���z�N�S�<&Ӑ9w��F�4҄�I%RQQP�����(x�e��@�=��/���~ࡱe�������8c��⟛���3��	����Xy�ߥ��$�p,���:� ��t�I�a)�ycm6��ܹ�Ю9��*^���Sz.��W�#��i�*_�r^R��3�Y��a�
 ��WG���OO�%�7��
 ��* ���T�ȔZ��?�\v�U�?�_Jԇ����ga`ߘu�P�ި�(c�Jy�>��I ��\:
���`^U�o��@�Y��"�� ���]oX��>~�0n;*Jv.e	��(�cZj��V���T8@AA��H0
�%bHe:]��8�%ôIt��3�QP��7�)���v;Met��j��a#���끳525+��v��z:|}%gxZx�h�(u�ƌ�v=M����<�U��j����
�����rw�S�r���z�٥y����z�aب�(kN1�1��2��ϐ�X1�<����|5(�
���������ê[�ޘ8���;��P� �D�q��EAAB��md���Z�ϑ�� *
�j-��oov&FC��K�w���ɤ���a����Ӆ�Ɖ�P� �

�=�o���ި�(]�j}6<������O~{t��27'�7-D{z���Fo���Ò��<�)�	�lJ�wi1O��^��(o9�k֣'A~��TD8/�p[�L
���~�Z�=�#�t��aۂ����!��q@��n�p�9va���(����#
��i��eDACy��wٷjJ��D��Z5`5�r�H�C���̐�D0�A QH
�(}�/�� T�؀n�^���Q��:ȗ���8PoX�����]a�BA{�ؠZ�Yc�.�p� ���^