BZh91AY&SYe���֭_�`qc���"� ����bC��   w���o���UA���b�P�HQJh�$L��%J�"m��
�IQ�i5���jZ�@+BmJ�FL���lP�����*]���c1��Rfm��6��f��Y��KI�m�V��مl�jZ�)U5C4P�R��֖kmhVU�1+`-��Q�m�>틮���j���i�-a�@mki�k-j�l�lɔ�Vj�m��eU�lX֢Y5M���D�f�mm�6�m�Y���3e�hY�g޻��l�ګUFx   q��4 T�۵]e��H�5��Р���*�U�T	��Wgs��(�m6�u�t�։u�tS'RT:4�K[&�42mo   =��ɬ���F�[jZz���K{�$�)�y/L�*[Ǜ��h��oS�z�y{eZd%�B�����K����)=Y��;��ޒ�/kj���[�t�J�v�^f�Y��­eZ-Em�Z�m�  >ﴥB";������v���;�4��!�9��[k������V�OXy���T��{��ޮ����{��B$�m�����R�P�z���f�]��W�[b����5m�֔�  �Ϯ�,����r�������=���V�i��ʻ���l��{��^��2��o7��m��٪�o��>�U��]��B�q9Ǧ�X���==*
�T�����46[�E6���  }}����*oW�W�]�zj���دY��v�ts��RT۽�w�������y�z��IV��J罶ӳJA����Fֈ�x���*[�{��zi
U���z��)��l$�#l���  ۾��IJ�L���$
��c�㪒�d[ޫ�����01���k{j�ޞ�y�z�;c��ޒ��m+k�ͽ�;4��S�z���p���^�I)B�4��#cF�����jl�&��  �um��U]Y�췞��ƛW{O=AN��k�.���ON�g���R�T\�ܩJ��͹����M*i{�\�on�Oy^p=�9�w� =���m�j��j6�4i5|   ������F�k|�KǠ n�^��Ǹz�z;`z�s�G�m��W����xn�CM���Et��v��i�Sy�4�lZb����[d([�   }��hh������֪�m�]�A���h��W�UF��{�4[x�4�d�����
P�Z���'����b֩(��,�>   ��] ��@�M�C���(�������t㧠:c�8
u껇������dw��T��Ǫr���     L�)J��mLLLѣ&�4ɈE? �)JQ04ѣ	� �d��JT� @    S�IT�       �? �US��@    IJ��bi�Q��RyMG�f���䟛���?��D�~2)Ҭ��lf�T�H�ͮ���ϯ��|�����������*��}y��@~T��P_� U�C�?����/�O�� 
��*���� *��>�T�l�������?w�?�����`�/�����������d}`~�YX\Ǭ�(zȞ�+�ʋ��+�� |2"x�(��
��� ����� ��*��
��s��������(�*�ʠzʋ�e =eeW�U�P�Q_Y}aU���E_X}dE����G�_X}d =aP=a =eU���E�	�"/�(���*/���"�� ������L����������� ��",� zȠ�� �ʂz��z�"z�+�ʯ������������+��2>��>����"�����"�������L>�"�� ��
>2(>���
��+̪�������">����*��(>���'ݕ�)�
z����!0?������#�#�#�)�`��3�#���#��#��#��d��̏�/��#�#�#��!������+��+��#��!���� z����2��>�>�>�����z���z��>`<|�z����?���մ_�t�q\���8����R<�Yx(�]���jЍ wf�J��POfbU�qͼ͛�����ᙔ��Ӫ[*�h�by&�	�ܤ���(�b��H��Q���{
�M�
`���'7qZn�vXQn՛p��Ƶ��\0�5�P�E���wA�:>E,��/�u�\)�:�Qc\)��ޅ�P2��Wr��6�;�^(�+sR{!�  ���F��X����B��8���
��;%�9J UD�y.�l+��.�N�f��4�ڕ��C�3r5G(4N�o@�-�1V�+k1H�q(YD�,g�))(a[�$<�`)9G�YJ��u�y3�y�8+��a����l��XIn�wId�`#m|/�{p����r=�U�*�y���L�nv�l%���M��K��V�Vf撋TU���cZ�!!if BP�Mn�!��$�u2P�_	7q�zG. �V��M$��O8s��֬�r
�h9W���
Vf8e�%CyI"%�C"P9�M	�%�4�-V��$h/�w�]�$
I�>>F��,2��u&�e��0J���zLԊR��6@i����R��l��	t�<�'g�q͵�Lb��H����_�ͅ�\���Fι��֦ҏ&I��im�c�3hP8�v;xsh&B��3�`���Zh�#(azV
фH���t�]%\��z�YXH��F���I��2���TU�!FmAd�ͅb�������o�nu�Z�֬@�����h�95��*��X5�0���1mڕ-�M���O-�u+��;�w(i�w[2QD�$��=�
N�����@�VA�Eaj ��� ��bP���m]bA6��#�{�0j�P�n���^*�����֘E<h@0�(��(N�Vv�D��n},
� GyA�:�� p��A�C��v��M���l~5��H�T3�ԠU�Y�F�U���8l2���	gVj�B��dj*��[��f����5Y��x�i���V�ƳZͲ�)n+,��&�e7�~P���ېMT!��N�1�!��T5�))��N��+aT�תCv�M���J��(��@��$c�����X�T���X���������U_Z�7O�%Z��Yg�օ��$�
�h�G2���u�QD[�
f���٬�ģYL�B�6�`����F\heY����)fk�W�{h��nL�S�-�^a
���Tz��wL���!����^�,I��D�!X�ժ�,� ��a���ŝ�<`m2�M���
�����A�K�9������tD, H�zƩ?K�0�[u2�E8�OM͕�9�cni�[w+ YPU<����		Z������e-�O�1�ȴ�J(�[��^������wD��F޽��f�CR`	C76�
U��q�'/o^ВPђ�!���f�Zww0X��v���H5Kd
�6�_\W[Q�,$�l��c�N@	��%�X݇E�2m��$bI�(�l9YcvȳZ��Ӊ�8iCe7$��XPBk������m)z��kE�:4�;�,m�)I�	Ll�e�l��d7�"tIװ�Tb梞��,D��oD
8ࣛ�LL���fѤ�9� A���j%tM�j$wv�
�B�c��y��J�6��[.n��v�%٘�۴��(̵(깫-	��G"�d�0���v�j�)�EI�k�vK{X��4L��:0+`���ܩy!��mR�1����7�((�d`�(�!Ш�dX!�n@��p���.�Xkr^�M�Q��e)(��Y���Q�sB��7v�Z;
ʽ3j'��fR[Q ��j�0%d\�0c�u@3��įD+fk����,R�N!w&��pZ9wX`@�$k���{���nn�n��2��35���ckIR<��PX����B%��b��V�����)lT¼22��Y@MZ��C&�
xM�(T¶a��m!�={0*܏t;X�ʘF�)�ݢ5c�C�`2�"�n��Z��ʶMBu�mY�e˙"�%��J�1��ڽ� ��	��P�pn3���i��O�o4�9�Y� �B���su���"��r�1a�u+W�XZ��A�X)�#�O�-R�sh<�E�1��rb{�R��-t�\n��Y%
W\݋�b**��s3hL��]����q���n�v�P�v�����˱(RX��#S[RmB��©�W-�_E���z數r�K6f����M{�7n΀өXpk�)-6��I�{�BE��i fd$�n�ZX�:1�%�����eø��R�I���Vѵ)�YdJ7n'u36���&����p�����]����u"����Jk��a[*�n䕛�yP�q�&�- ) �	��ii�rd&Ҩ�m:�s�V�]�W����v]!'r�Q���M�Z��kf���By� �ɼxrm��B "�r����LT�n�\5{r_�pm�ΖVB�LR�[x,��^�
��条���1��#�H�af�7��2�+���-p�����&��9�vųpdt�5��5�ǵ/l:�u*(��r�H�ri�B𼼊VIAѵ�lz����˼ �jkOI�f9`�7��J����.fh�
Yo2���0�-Lom���B���	K��s�xV̘���hJ� ����h��H�4ix�\�CCX'08c0����Osj�&�9�RV@FţY�d5w$z0JYX�3t6�Kͭ:Ó	&佌	�)T��hA��B�n�L��X�&�Ց�r�I��,���1��S\1�h�e4b%Bn�MLצm
J�ޥ���hn�Ҭ뭺.{���3�R��̦47��4��*B�tu����f�j楟sU5p�Ӱ���v�-7���`�N�ҒGt�ݡAV�A�u�h��U���3�D�;6H[q� �����[��-X5�UdkUL�/_n�q|a��i|
���T��chM؋�Zi��}wYN�ŁK�W�f��PœU��.^ t�˳Z-�qi����0'Y�����&��$�T�\����)��[A��KN����n�ʐ�x��`�3BM��Ժ8��{X�K�$��7`���"=9K!U�CB;j�p��z���Y�RaCA��Y��恗�R�։���@�,w"��O�G��!o[��DԎ�Ǔi�V�24X�τ�yoh�c7&�IT��ͷ6��ѣla��K�ʥq,�R0\Qse윾O�����vp^���V�T�3h)7�FYt�ZYr�#��ˍ�Зn�Z]����F�ȥ��b����&��g� r�n,�[��)��ۺ��`�-��#����"��na�|-6u
u��=��X�L�F�XI�JD8�ǡ��Y��Ź@����x^ۧ0�bZ������\]��!a�h�uD�&f�z�4�XA�E�Wz�vP�g�t���5��H0nĠ�XA�	$=f�#�`�
��lm�v��엣�OSX��2݈el�JmַQő���F����kc��U�������$���m�
�`y�2���f�lJ
Cm�lb�*Olס�ujcIJ��i�K$KP�1A�l���r�"�f�y� �;۶���19B�d�A�����d$�H�p�6qS&a���e6�ѥ[������"׊˻Tf��c�k]1�,i:!ЪQM7�(҄K��u�F���+���^��0^ko��fh�,�²'�id��fb�A��ZN�%6��P�96�/oR�aLvC0P��B����n��XIAb2�85 �2���z���c%����4�a��r0�bO�-���v�x�f������W�p��M*H�W�ݛ�s��	ȵ"�Yu��( �s�`���5o�#Sq=�I��[��"Ʊmm���	��]悶�C �d�^QȊ�&�����% j1{!$�ـ亖-m̔Q�kr�F�[P�X,f�����&l����̐��o*ຊáMm�2Zd�Wr<�y�PB1��rc%h��;��X(��	V��p��� \�;E@�ۘ����ïv��6�((�B��݁&��u٘ΝJ��bh�A�^��)����Gv�jF������CA��+-cUp�l���2�9���	3Q���(Q�\���Swe���Bt���-$��b�����m��&�j�K$ ˭z���t�N�kժ�/&ź[�jnQ-�J���Cq\e������1 ^�6fKh��!4Ek���bkxr�%Yr��D:#r���P:�E��@*ۺ�[�-:BVY��7Z�Ll�Hi�MmH΂1^
�B�T���[i-�tEu�E#�
�f ���f�k6��P	�a/*@�<���u��D�AH�#�O��;] C�jV����ꕘ�ͣ�0Pe�@[���d���U��Z�@��b�yV6A6��+���P0�������ԭ��sH���n�koB�wh��!+ɯ�6na̫
��n�]�Cj��{����˽�e�.c��*
E��D FاT���)�V@b�m�H+���_1�Y�ڃ%�Ea�+R�M_�n�o(����}�5LV��,YQP�1kb�l:_�-�gm�$�.�`u�֟'��l� �6IK&��ݬ���PF�]f�^'���Scu�/� �J��s)�t������96�[A�H+S�ٽ�,,=�E��zЀU�kk��5�d����}�)���V�
��B�\�������D�[���컊n�O k]�;���[O�S��|��)��f�k�U�vi�٠E4S���Eͣz�7%=jƪ�f����seCRB0T����^	n	���:��ǹ?�7��W��������L��bك !�N�ځ)��C�Å�ܥW,d�Q�+h��QaJ9�dō;��5���݆i�Nf���c/	�$^�kL&�K��sL�ɸ/UF^`�r��ۄ=������ówfϳC��c��CEZ�eD��;��+-�ڠ�	��Y�L�kK���e\�dKM'G%��Q�z՛ղf�i�.��U�ӱB�ɂ�\�Z4$A� �f(�����V=A�A��QW�b�ǥ����p w�e"_$�^��Z�iS	�y#6�ڲ�Z�V7�2�)KU`{���D^m$�m�o��+{F�HGv��)X�Z�/Ca52f^�������˥��(�Ac�u�(s4�;v�|�݊�;�k}�1��W.��f���h\�Hh}d
�_�YYx�3A�ihm�4p��u�,�i %Mɲ��^'�Yؘ���8���u�SA�,P'+"����c�T.bE[�@3�v�hƪG��1�V�y����࡮��9%&�ݺ;mf�:����K�b�XɇtFU�L�nK�j�]ا�Ԭ�(�Zkb�eܥ��oZ[� E��[�%>i!s�o���������]G$�T-��s2B�m�uB�*3PY)��=�#�r���XWB���ŧ���ʠ�1����[�1�#)��]�w�e�5�S�aP��z��j1,�V�y[�����MM�c�Se=n�=9�L��X��Y���E2m`I�Ÿp&�l-��hK]�h P��+ei2��vR�j��m��[>��m�/�u9�#�vH0(N,�-�0�6���*��/�kڷ������Y�}ذk�8w.�H4�tX�����{s7U×��p�̥k\V⿷�IOe��͠�[�O�7��ϐ��s�ʭ�%G�`�Q��92-��2%c�J�h�N��t�J8hF6e% ���ȯ1�X	�����Ƥ�Y����n`)z�1IY�p��`���k5 `
�r�!g`�9L�қ��lV�G�l�&����v^ō��&��:�G\y�h���x0�9a	��:�m�
��^sMՎ�A��R l	�;�\S�n��]n��C&���lz�"�*j�q��MXF�j�b�-7�����&��;5���4�#�J���N���cT�M���ǌU����#"r+��m��Q"��'\��[N���e�	*L�S[v�nڽ���g�V�Xׄ�@CZ*���:�ocԘm����%a�T^K#�#�4Ay/DPڭ�,��{��JhQ�gfݷ�Lɂ��FK!b�B^�j֑�4�xҧ�Vh�$�;CY�F��J�-�&�r�fYVq����6��+Y1k-R��)S�ZN��e̡��!ц� La6\����b�+��U�en�d�C�m�dЪ[˼�A�i��KI����2��{��Ӻ�(�f+?]dGe�� ����%Ռ�3k)��b@[ʗ�R4��g
���$k,�xP�&�/4T�i�J��cu�;H;���i���ż]���gܺu�M\��2Ӊh8�*;Q��[W���:ˤ�Y�6�0%�%��[�_<5-��M�KUh�Yٛ)Q�f}����7�(�l�������K��y�	N�Gj��2,ݽt����jL�諟
Ct�����*�S�oh*eC��ֆ����Kc%���X�1�V�����YED���׆�\�1kjf��GL�
\���4��I��%\�c��_��	��C6�ZwCC+ۃ [RU˻Z�ݠ��Y"DҬ��z��W�Q�e�A�5���Mn���%eT`a�Sp'$�,Sor�d�aת�$��
�����W-�C���eӐm^2�qܰ�mp.�s�>��,�:�Bm�»�Yj��I�I͂�61k�;0R�:޽������-�hU�C����T%���f��ugf�ҲF66壴�.��|MeL (&'e��Enm��EB������5�/^�J��wwG��Ws�Tȑ��y���P2��^���րd[Z�7s��[Эrtr��G]3����hީ�qv�f�RS1r\��F����E�eWo	)]���X% ���@�>��/ͽ���~���^��@�3�����7�����n>c�Q�Tӵ�˵Q����eJm9�H�c�4|Kᖳ3q(�GE���Z�V�bh�$�j���\�}u��=�k��u�Gej��:�����2�k�[���h��&��[5k̺U�U��[�VJ�ue˔Ẽ�	ś"�J
��Y@)3�*��P����q��]&
U�� }7���{� ���=}��^e�x�>��ʮ�W2�TD�����k��)Vj�} ��y%dᢅ�-��<�;˄Z��3(�98�YC��(���Z�q�}�h�����}si�l9�;(���W_pe*��'�va���.�jT:�j�&��B<�nR<Z��ؙ�}Of_*Z��stؓ�U�2��vĵw,Z��B<[��f�T�?v�A>�X�j:�A�;2�u7�%���M�1���K�*�����j�4����81q�u�Gn�U���S[�&s�p�!T6�W�L.A��B�Ì31������w�k�����@�a�&��3kU(l�8��AǺ0��2��R���Aߺ�h���8�Y��RT���x�ح����i3@QB�����nm�&Wj��#�T�XjN�;�9x�q[��Ζԅ+��*��͔Jc�C�౰V���ۛi�o9ys'�e�ɀ�91}iS
J��;�K�uN��]=yq��˖�c��U���6�1���MR󘳷��l(��ʷ>���U�U��4s��l�u��E����⑱��Xת������yzzlr���>̛Ɨ��κv���i*�y��{ό��b���#j��q	�+7���[��d�� �g0�F�7���������Uw���Bv��B�������
ng}� f:��B�T;����v'v�]�0����o
�a�qrk�f�ge���Y�
�9ʳxM�[�:�:�囪�5�/�D2a�[u°�v�T�"т�6�}���p���M4�h��k��h`eo/I���x�Q�#v���s��.pIO"�Np�����y`S䁮��un����-Yͦ��C+�)�L���墮�'93�],��.̦��p�M��Xr�7au�wZ[�s��ѫيC] C+1v�R�V�t�֊v{��;w��+����8m
\��v,�dR�t=u�3Q�[�[%�O-_-��㮸����iuˁ�o;}��z�<R��#َ�Ox���6�gU��[Z�Y[����V+ؐ�f�c��+"e�;��J��yxV���%=Oud5��,8�m�c3d���c0��A�5�(Υ���-�`��r����Uk����l �ЕH����f��ER���,q��"cw>`��n���_+w���ͦrGw�'-}�*qR�Đ��I��FҺ������Ɨm���d�U{N[Bp�ʫi�g�;�uۦ��aާ��nL=7XԈpҫ�r�����.%D �H�9�t���ά�H� 7�L�kW]p|�5�c>"�8]����*��W���v)e*u��9r�6ޚ��ǐLe��6�%��kX�[|� F1��ה������mځV�'��7��������.�2��aUכGq�i�D����k���j�U�(c��Iv���`�n�E&�(�	���.�}�ا:�#�̬;$1��pA`5X&\v���;����-<��0�}z�kc��f0��I�nԄ��
��(%��+� ԏ����n���B�Ԓ�r�K�Iۻ��	jQ���)Հ�,'�_n���:���6+��:�>Ҳ��`G�5e���Y��+���W,�O]�gi���r���vi��H�k��Y����-����̔�$K����p�ޅp���k7�N��Ε��]�y��d~���,� ���-��m(8��6�Y�t_����nkJrR��ng7���4�ٻ+Q�]h��C�"��B�	0����/`L3�fw-��eF�j:�!��B2��l!�v� �W�ƫ��73�_W'|�.�8Ưv�������m1�ծq�K�,�#�sU����d��t�0r̢Y�z�;̧��6.�<����|:���+H�/r��wǝ��6u�4��7�b?�eJ����	�x�7ޮ:���u�b�׆g)�ub�4���:w_F7n�^Q�(�<���N�15tl�۔�Qwn��/w@�&�x��́��|��%i.�����1ݓōY9�Y��j��q;�gK+LT�"]����+�T.���gO+�e�+rS:�`<������L��)Jv2!W-s��SF�,f�s���9蹲�Wi�nGs+��[k]+��K�|7(Mݫ��%լ���N�9���u���A�-��}g�����;)� i�4]���Zۘ��KLu�nޛ�^4���}P�[hS��ʲl^?3�p�6�[��V\�E�d4�vqW��gT�&G`�0����ӨC�Z�O��&Z�LVl`W
��YY����v������T�:�����x�'�\�����5g����&J:�VMa1����\�E�a��GS����w� �(����0�9	��*��A*Ǳ��p���J��wE��*��NT���h�k��kg=#I��W��3�-�V�=Ρv?t��B�r�B�Ra�gR�+ut�����`�3}����ʀT�Y����P�j��Զl<���p�x���B�B+�>T��Df�&n���(�ı�E��o��`J�+,�%�Ֆ���^W�Q��=���=yQ҃�G}�ͳ��,����fZ_c���k���U�4>�������-�m��|��ɚ�1,Ĕª�ko��9��wR"��p�XT���9�vv�7�Mxsngu�V���@-7��豆�wrBۼ��f��G2>���G&ژQd���N㛬�B\��h��FgD� %��qK�&k2pwi�_.L)pv�j��Z������=��Pc�ū�3"��DC�4��OFDAͭ��;%��\#��T6c eů^��m�HJ�T2t�K��T��a��M�F�e���3Ii�RV�
�-4�Q_s]�/��*�[�n���P���4֋Pm���b�h-�Vc]��|��wWˌ��'VJ�cO�k�1�rI�g2z��>�c`׋�D+�&��0k}��I��;�S�r^Y����F�';:G�wW!�#��v�h79��/L�S��p��6��Ik � �D�u�;ٻ���$�ͷ�y����,��9����Q��4�S^�ұm�J��ؑVӻ�5[9��e�w*�BsY7��H��E/�Un#�fL���w��n�l�J]l$^��.9F�%�q��.���6:��%��ne�R��۵vԖd����ȝv����̈́vm��ܬ%�ؚ_"��lMs���t�.���W�2���#�p��J��!ַ1>���5֦�bn���T��� mm�*N��Y���]�޵[�k����;x"�A��G���tY���WBv��E�Z��f�t���S�HR
Ks ��P�Į�`���I�:Ǌm�}��@�{1Z<&;@�K8��{D�I��0J��
�%s�}i%�E��+1����n����֜V@=�����T�4��U�U�[�����$��wp*�-A�)ljGN��l�W����͛K_hnC��L�A�t�����`�IJ\�7�0�����;�_Z��V��ܳ�%s�M�2D�
Jwf������o5��lX��1;
G���Ii�+�toMHű>ޭ�Zڋ:��Z2��B#�n�J|��,����sCv���XfrB�:yLu``�r�v�{�_ �MP̲�kJ�h�<M�:�	$�z��z���F+��d喷��&�x��O�$�c�h���΢�=�3����^} =��nE��A��d�1̛����}j	/�ɼ�~�� -A����f۵��U2�[:r���e;��o�{W^h���:��⁇���d�A�s��6���R������u����)�l4���a�]Fn��t��vZ�W���٧e����7�k��em�]n���չ��.m����R<�zʼҦ��*�T�T�cz]wueJ�v,ECt_�ɧ^Յ-ʻ�[ u��owhT�.�p����<K���ѣ�8�a��F��i���EC��5L7+D�	v�i$�tUgj���7\�p|؞�ֳ�����s�<�;��pBh��̠�\x�A�2�ż1�|��,
����N����P�rlp��ҳ�U	�[����Krӂh�>�7{3��f�NF���ʻcw�6�gChPI*���.��`�zG�J:�.���h�HNÀթ^}&N�˦�6�ZwA�;�1j4!�=ˑQ��qu��ki�:n���Aښ�i�t��kr��θQ�́l��o\�J�x��/���;�)Rח�Y���/uN��\k�� Tp�J��H�w�2*Д�ھv1��>f��F�ɻ
��i/w�\�:���D�KGvӱ��Lbo �[8��2�*ݠ\T��p�#���fu��9[��̵-U��_uSǩ�v���(���9ټ ��0k6ָT���8�`�����eg��L'Z6$����ysqWR]Qp����1#�A5�d��v�@Ey9bͩ"R;�\�-��7a��L؂b���!����v��a�d;v68����jB��IA� |C��N��`�v��[6�8lz^�rv��Z�L�Vm�"�$��o�qkv. �\�{xU���I=9c�'�Gt����Z�(�=��nVX��T���&��HT�pB�cb�-,��\��ǝ/0h��VJ&�P�J�mG/��/O�n��ʘ/Tn�muf������®6&��bG6�����t��zByts�;w�,���m�����#T��I�W'��6?�uS�[u�b�ھ�BTǝd�V�q[qG���7>}f>�.kW��[����7�VX�V�>��!�;�謤M����D�Gy�OjDֺY�ԭ�u:�cTE5���0[�l�Vu.�LJ}�6�,6�1�n�xj:�y�����.���:�G8�)dN�j�A�����r���5�nRZ8�ҝ��	�6��o4b��%�����'���U���,��U�\ԯ�s�wg��m�����؝�+ե͜�Z@�T����v��/T�
���z�^y�%��qnja�<���Fz���]�$�ð�E	+���Z�h]�A]"B�8�XY	��s�L��A�6��T���^�R=� Ԯ�7ˋ�<Ö%.F��i���o�)ǔ9v��GzA�7 ���@Rw�g+F���]&a}B�}Vĥ��6mt�iq�]℄H7/�W3z���E,;V9�tc�EV=�D��)8�T_Vv1�&�-m����]n��z�q$*B+��m��9�x�C�T��5�ǰ�;2�Ḟ.�2�z4e������<�����
 �+{�f�������	\��!Bѩ�!�ږ z�C���@��e5j����͙������pB>���j�m���������Q"��}z�<Z!�h{d�{�u �%�8�rM�a+FwK݄��F�\�7t�YV1k[ƅ$I�JQ�K�c���L�����F݄������K�ً]���T�������gKr�W6)�l�,�Xows	ta��d����5G&������[)Xڏ�����.�٦+�4/�#N�, �ǙK�ȯr$7��A�nb��mÍdJ�b��N�qN������a�D]p���EՎ����1KV.j�-=�ζ�*,���O��t^x�_]_�iА���Z��<{�p%�j�N�ؽ�re���vU&A�����m3�n�E�RE�Z�����ū�d�T�mʗD_�%�63_Esjm`�
���U���K�U�8�C��XT���>|j���^�ȵJ�ʘ���56#e6�P��=W���w36�.��֪̭.G]�6���S�e�TQ��)�
�Z]d���W	)1b�Z�ݭ��qC8�%����ny	�u��m��O9[eS�J�Zk��o6m�0R[Ը�w���)�d��Q�r�'P�67�L��GuXƔ�́�]7���r��ގS��MG/0�B���kY��(X�pK�K�Y����)���Y�_N۳cil��Ħ<kS@���2�8s&&h;p��X\��7��@R�\2�3m�}4���/�`u]����Y����g>:i��Y#E��]u�V�d �.50}�Բ%�����;��s�P�/�<Y�U����C��P3��,ZܫDg{W�J.��v2W}�q�shm\�p&c�����D��M��D�t�K��8a�}(�����[T/K�x����3ĢD�fi�IZ�
���4���q��R8k�;�f���AK�(�g��zh9@�BO�6b��[�4qZ9�f��q�IxUY�����;
��1�KD��A��P��r�C	�
����&V8��od��Ҷ�f�HHg-����E��<s�z�aN2z��A1t�����Z8�9!�Z��52�ѽ��N�98"�2��]ޘr>cGf�������P��E_��5��Ǜu�zo��9S��]^7mS��R�G����5b���
�3vUJ�8�R�ibwo1���Z�ǎ�L��W��"ǴHa��U�Y���λc�ڌ[)@|�������(�����6�n;�Y�O)�K�ՙ#�I���z��ƀ�#�M �eB$5@�F'Q�*!D %6h
RӦ�h��B��2�`�i*,�@�ɰ{2�)��A�}�?|�u��k��$0T�����Ւ"
�> �G�LI��4U%H���:���
��wnu�y�αh�y�������//?ڢ�����?��<U@������~E?������DE�������ߟ��~^w��o��|?��y
 f;�1T�E^N��Q���^�CN�/�Z��j��[xlV��o
w:+U;i��\�#��T�)ƃx9�ivNB;'w�1L�S}[��U&��k܉J�l�1�h���=J�66����MzF����ض��WT}v~��'�	�mI�{�r�����Z�}js���B���aJ1���c�vQ�Q�`��4�o���]|dJ�O�dv�0��T%��5�x�o*�r%+MU�U�5�Qkd��Wr��\<�Lvc�u+��<wqmգ`��kkb(�(�ݣ� ���t��/N����p9�ɏ:qxp�$q���v]]��M:n�4[����]�rtl��\�������:��j�9��ӳ4Ξ���ԃ{lv'���� �5z$L�Q^�7yE�G;x�˥os�Y���dD���������[�0�U�OT����i�i�S�qP�}�*�Jl�	n��iퟤߔ��4�{��c�Msm��Uh�*�I�&�s|�+7Zjmg*Sn��
����1��J�Lro=4�=U#�d��%�ХN�*�a�ʞjј�i���q�����a#]��1]d�Q�HI�g[�C�$" ��N4��W����P�ã�v�ø�nf4�o*Bb��8��.��8ze��J�S��]����� 9�#ˈ�u.�f��\�ɗ�(']T�\�Q7�SW71�؟q.��2����;z+�h���\�����V�u�;�4�La�nq�V��1��P���s�k�]t�����T�ނM����N�m1pk�w&����-jҌ�jX��죦��TS 7oI�)<��w��6�붰�4�TDZ�q���$bܤ ���� ٶ���+iu�./S�[���3e��:a���^��5zw�uv������Yh��͜��o�5r���,�5�M]L��p�v���F>`f>S	ٜ�Y�v:���S��^[V�^hRs��Q�ĳ9��G��]�'J��1�� ]6у..�E��ю��'��q���r���}��,>�)@���*I�+WVq���;%�Gs�̿��hv���+�/08ԤU��
���XiV� /��� �W��9)t�e�ǐ1�]�s�
�U=Ԅ��ӫΥVۥ��mv�3@|+Tۈ4[����MEj�s��\�]J�vu���	�@ب�	h�Xޭ�i�T n!(� l�g-���1�Bl�{��A9=Q�M�#j��8�m��֍��E+�:�9���Q�*D��?h��]�U�H��9��(��&�;e3Sm��W5}��ՅG�S�ń!�_R��i�j���M'sea���km�q�ͷ��ԏ*�Wl/�y0w�1կ��o�u�p�[�hS�8Aʱ�%����E��"����Gw�Bu���	8W��x�̬�@��7�r�l���5�:B;���{�*��M!˲UNKr�VAE�_eħ�]�Wgf��"����Zq�Q���,�J�����F�/gA2�jP��0�L�$�x8��{&��R��:�(n���flM���W��˫}S��S��H1���WU&!��y-u8��#N֣
���	��Ғg	�y�Y�{��D۽�>b�A�9͆pCxf�� ��u����h�k���w\�Ч�A�"�s�X�+=��ɏ�p�N��N�*�>��*��';g^�X����c�:FpT4QP1���<Wj;fM�/hL�r����h�ЉK�t����αq�R�����K�7ww[Z�s�W״�̺h�#B��6 9��B��s�3�dڍ#{*ġ���ܭg��k6�S	���6����;�r�hk%�lT��#�Zgަt\��s�'\q�҈:����dw��M�ne�Ah�1�8�R��Pj1yq���	��4��g@�,�)���8��u�8ɬ�K�lj2��ڨ��E�w��Qo6�Л���^Z�G����l=�K����ő;�b�ܧ�"�k6ޤgt�������ӝCJ�C��Ap[ǚ�v�D�Q��������-��U'v��v*e^A�Z.�_W>
^��a�b��3:<|e���A��p�ٲY��=}�*�]!4�]���<*��q�6VkX�H��\�vCw�B}F���dk���;�3L�z�;v�Wv���䓋�Bu�����'C%A&u,o��gYG��1K{2�X���9Ws�9�1Fw.X���l��Їu�ey�!��qIN�������4v^�9�Q ���R�g<V�[�ki.��4�DL�ڠc=,�B�4�oPlj�ݽ�>u�3���&�{n�ӭ=y N|̼/:�͗�P�&Ibex�+;��VrQ�T�Ӱ��\�TmQ;pp="�t+(�C|����Į�[��2�t]+O�T�"�ֱ��8�'av ��,7wç.�:EB����W<���%3�Y��Q���z�;�+�cXd���J�*����mn�t%�Ύq���H�{�u+Չ���K�r�P������q\B��so�"��fp��s�oMX�����`���&�5s��٠�#.E������{��\�u�����I�Fr���;v�Kv�b�]zX�X����3T��hA�V�( 4��\��1��7S`"qLb�Щ.wz*5s^��^Po0�����X�S'w�A� �c�zx(��o�E�����un7�AƸ�cG�W6�;&_.�u ��������$0;x�&�>�>.�"ֲ�s}�������֎�L��P�s9M��.�S�:V��Q������\��g�5g�;*fg��C%`���t�����j�I�f�z�#s6��w��۩��0��`_ky(S��E�6�,u���������z�2���Be{�����B[��s��Z����͐�3��u��*Yj�2)�_s���3hI.�2�'��tV�Gk_�N�A�10;k#~wՋq`����l�L��3�,|�}�:t��ƺ;�܏���[�jXQ]p���ur�w&��n�R�yI�����*�%i�)�)�V:�Px.`vZ��]��1�ח��&ր)q�Fj��kaON�X K0:Z�d�ٮ#�ޫ��0��v�����]u����@'8*�N���Z��q�
k0�����'*\���H�m.S*=�Z#����Y��@ƾ�]5���ýXd��Vvڗ���a�l�Y���Nu�	R7�p���I6�DUp��ʓ"$n�%Ŭ`ܺ�J��j�C�D^�}�P(n����uÁ���@�⾂.�})����\;�7�(W@�8w4�i��XM�]S������:�,��LYeҰ����/�=���ӎoYɬ� �D�l²:�݊��Y6:��׍���� 3���:�vW.��JT���ԙ�^���()NR'w���yy�%�tˮ@ugշbX�Z
��5��ͩ����n����.'?�rֻ' �CN'���ͧ]��-ҌC%�t�K����A
��P(�:�����fQ��8�(5A;�C���),
�Ev�,�5[f�Й΅lQmpv�#���j��J�K��uhS���V,r}��ޮ�x���X*�=R� ���)h.�8��<G���6+aj�r#$��XU��̿�#t�A��+tk�� �*<��)����}��X��.�Yx�!�T�m%�Sb����f�D�&�7�n�M���� �I�޹BC�st"�V|�MWbd���)�q�ksF���V��6��՚h��v1�ع2�V�,V�R<Wt(s,ZG-ڌ���fG,Mt��\�M���l��#s���4'rWs*,���l�ƻ�g|'KۖfP˧Σ	��Wb��ƍa�^���B�3R�������/Q���f�qf���tȕ@oe��\���to(�'ؖ��]�w��HY�A��s륙����qKȱ��v�V^Ο>\E͆����`�,���;�p蔍wq��{��N�4�
DiP��;w#tx��{��WU�0�G.�ѫrgY{�Z�0v�.�^�Ҕ��Hhԧ�����d��cw�Z������G�D�'��bޖ�>�0)��$%�E�T%s�_>Ê�Y9E��6Iym��J=]7����
H�U�6�j1Y�X!ѣ]P��R�$�5ee<��g��Pf�� ��lN��{j	�Z�Dުݝ���E�r�2�a�y�^Wq�qο��P|��%��y�KQ�<�I.�6m�w����е��r��R).!<Y*�l_m��1,��pc 9m<�Q����rh���Q��(�Uc`����+����ٗN��a�T�%smTXcΎ����Y��/QҊ�}�{��,S'ບր1ݝ\v�L����,%����<g�ݝ�Wɝ4ٔ��Xr�J�����ʜxd�b�D3llD>4���;�!�qk5L�wn#�т���L�^qG������r�\��tەWFD�E�I}w�t�ʣ���8��k���v��K�<]q��P���Bɦ:��=R�:��� I��u��4��Ҍ��F���G���5K��#�<OE�{`:H7;)�~���	��W}q7ҌP�+��� ��G�0��7MC���@��� �V˩bG#��c�s����u��ia`Z�n$ٚ�C����t-�:��A����ԫ�f�o�ܵ�	�檹��c�+�_:aR��$˽�ʡ�َ[K~32��1�n��_NC�TJך��������P���h�A��B������}C) ���U�,f
X�w �H�1�]=�]��耵�
�����Y-��ā���;r�Pt�t�	of=��nS\�	1�Ճ.[Oȵ����Gu/e堬nV�O��y�U�K�t�rŮn)Ҟ�n.�V��v�+�X��n�9��7��Gp(7��Sv$J.�ֳ8#�A�t]�P쇴H����D��N������\F����Rg��bmJ���|jvd-̦��1��Q�v��7ò�����W���Y��h<ё��R�)85;�m5� mJ�b������4H�Iv���_���/��ڜ�����5}&0�%�pܝD�����p���Ed����@�r��%�Jc��6Ƞ�pS��	�� ��OL*�掹:���T���@������&��9���ޚO@� #�4���d�P`D�	���/��"�Y��z\}�0�WWi��s�u2�=�S�1e�4c�es
��@Q,���\���V�d�#��Y]u#::��F�6q��\��"A�:�Cǥ�D`����ݰiӭǭ>�H��9g��l�ƭ�N���3�� �;t��b���/��;_M��pr�Ink�wj��.?A�)C�����9v���������w-�/�#4+��r��rŦ�oUJ�t�S��!li��2�z����7���T��u
K���X#�km��9�wE/	��ul�)�|Y�ͨ��J�cz�'C7&k�U6#Y��;b����< p�����)�Ǵs��!�xa�;���c��Z��2=�����B��x���:��%���������Q�Bu�*� �\�]�����[5�GJ��q��Ec��+�SkivqVn�ñ�l���੔ӗ���DXr�f�\��`ƊG$�vX�U]*�;N�]0oM�J�+�Yv��O�8�7���L�b2��i����S��q(�]����/�Kdk�	dLC�h۝1,��k�I_��@M�bąȆ�������n_D.	�5bu�%6�0�p!����)����|*�udb�;(�O1��B�n�վ�4�U��K��K{S��C�aK���ZSJ����4[x"=�ʡi�rR���+$�u�q�+�Ш��X#kT)5��]�5��~�@��l۔,"d�[Ϩ��'��ku:U�+�k���J��m�{�=�\�=Og%�I�:�Òvb��!���}�CFs_�8SX-�`ު\��de�cg]e��EsL�B�)��6 h�ۡ	#[�VK��Y:&�l���ia���om�f��DtT7o5���]�è�p+r����oST�GTr��\�DӴ�U��Ⳡ�f�=��y�8�^��+[��4����Q����F�ἧe�w�2��2F��pY�;�Ѯ��ȨN'��xM�םB��B���j9���,����ʶ�@i�I���-=�p�>�vᡬ�n�s�J�oנ�Y�Va��$i*�<�ac�|ƻr�^��V9�޺ʹ��'��'�R�wh�N��3^�h."�ЧlXK��Ն�����}f J�,Δ�g��W�ۗ��Rf��ŀej+
��$̐��7>@ٜ�Jgu�o@�A�,���q��M�<�u݀�6b�b��a�)�]���9��۠���k()�s����ou�)_I�o��)�9*��p��\��q�n9�hih�{�H�T.�k���J_L�k&�����(��W �VR@s��X�Ҿ�읜�X���1og1�t]I��a������yM���&顱7yi���S�ܮn���zoѐ��Ee�\��/�2(U���"�m%�P���C+�u3�Y�]���yJ �mh�3����	;�H��u-���k"]]�!Û���pF�S�[�'-n�;;�:��Q��?S�o��P�ݺ��>��#�33��E�]u�q��s������v�6�P}�M]�Ű��Lc��k�E�|�1.���etdͮ�
�yp�Hͬ�5�`���V�9k��y5�a�Ӯ[EX���"n���.;�>������� J���������������?�����~��_����������Yhق|D���_*d* գ@B�/�PJP�R�o����P��]��l�pJ��o�G;"h���0�:�E�ԛG�s �ݢR#)`F�b#Ya^���4�G^յ�JU�������E�^���)��e7�MI�`�V�X�Y��*���I�r�{u��ΊLEfҁ��8�g0����IZ��B�fk����u,GS#��Zd��5�Q!$wu���V�}�m�\T�@�x�fk���^�+#]M�JHj��;�>]�r�U0^T,����ݧj�[9�6��KQ��U&ؔ�^���i�l<�ܒy|z,t����=!w5m���UhD�m�qw\�ށ���˭���J�8�|��N�qt�u�{�j�,�W���}dnvk��ch@����9L=��0n�#C����,�Cr�o^6�m3l�͒8�b�4Ӕ[���J�r�]Z�G�f�k��q;b�v�(w�T�&	�?(�ztf��7]�&��*'�ʳD�]��еV��{��2h5�+�h;�/S�-}�\}�.��X�Qv�Ħnѝn=�]b��2�ʿ�䐲6����fˊ�Y��V�UlM5���3��Mi���ض��ԦY�&04��6Qy	�'������ H�nD�T����e�#���C�l�ӋO��}T2�P��lo�ѷB�i�7��5%EU (��g$�I���4X�M��1F��h i�qӠ(2��y�'��y������G\]X��TN��Q�E��Y5ۭɎ��*�tk��G]ٱ�j�:
���� �㻍�֞�b�����c���S�mcg��q%�G=�]Q��-Z���b
���틜:�uF�mSPv6'�ۭD��P۳O��l���4lU�����u����;Y�b����u��ɮ����kl�5�Z5R��N���nj�7n��k�ۻuѮ�ݹ�ݎ�����w&�DZ)�AA�q=�vŌ��tP��mv�]v�t�VڢۭX�v��I��WƲWn8h�\GE��V����Z�;�E=m�tkw�a{n�K�b5ݭ��JAh��V����i6��AwqT�'�ƢͲS��ET��i��x����A�TWN �4D:;�� �PV�Ţ��'"(��(h��5�jg�zkHSmM��M�����JCX��]u]|E�����ņ 4��T��Cl���Oj9�o�\����VVu�~�˻�T��xzG��.�&�]�XMڇ&sWE��&q�S`4h�TJ�g)!*���Y�U>��إ^Ǥ9���f��k��O��\��Gzo?�"����+���`������>�n���e�Ö�˵�����)�I�o��_��i���W/�O���nN}��8j��ͭ[������y�U�����z����j����K�]=���~ųm{#u=(vw�{}�zE��T����G��:��{mW�}��lvc~"���I�>[��ޯx��ӳ]Q�
捆G?�j���C���an��l�o���:�5y�~��x�����OoЋ/�|��Z��`��m=1����������K2y�I��Q�7�{��� �\2�ݎ��`�o�Gy�-�|�e�.�-_r��{�|�T�~\}/�ZBs6g_u]\�^�S�����(o�)	^%"����Y�	��s�:�t�t	�"��5V��E3��%��'*���V1������=��܏�/˱>��sC��Q��s����(<$�6�nC*v�a�*R�["t��W5[u��E�ԁb�EYT{9�Wcs6�[� ��IP��mFm{Q���k�p�o^��ފ�q����Q����論�*�W�)�,^���3/_Ouͧ�����<�2��o|fЙU�)f�zeQ]2��}bɗ܌{��ܪ"���Ɍ�1͒:����)?+�Vp\��*��zq^�q32ĭ�wW�o�e�׽|���yB8귪R��޿	\����b�nDI+phwIojޙ�|��=E�:�9��e�w�[�_��g�Kl�F�`�T��N�Wd��g꾪D=�V��'
��=��}���6pzJ6�hS0s�ן'�݌���ҪK�;��.��D��4�]OW�ޛ�F��A�/���n�2移��w�'qߋb�D�^߼j����y�����f�
��座?}�}�y{]NY�mJ��|��U�6}�|w�����yնwZ:hn�ջ�a��׉����M�8�R�Ư�b�"ɵ|ͫ}{��xW4���m�]F�ϣ�=���L5�jV�+4G��b7���u'J��%#�}�.�Plv��ƥ�� V8{�+ *�j<5�>���ɛ]`4�1C�kܚ�����j=Z\/��8h�JJ�ᅰ�J��d鶰;���<��ǎמj�[ M��D����K�����y[_��op=���=~�^C=�q���cϪ�;�������s�==���Q��e]ׯ}��V��;V�$Er��qF�S�*1�;-w������S���璘�r
�k��2{���Uu���
�?��̻~�Y�7'Z���	����u�ǜȣ�S��u;;��5|�֋�>��gS>��݃��%��>��>�^��<�����^���E]Ay�`h¤qG<׳��ؿM��U�������}���l{��/*XP����Y��մTt�A_��'L�=7�7z�u���uЀ8ѩ���#ķ/e��z��ڮ���?P/|�;�Rs7������f<��熇�R�k�<���n�����\[�����3�O��ٞ"���J�C.�tVtt�oL=%ڻr��dEBn
p{U�m��]{}�6����cB��<�-6�uo��l����\�<�������O�Qؒ����ՠz�9�8L�I�1���Dzym�u(i _�P�ʘd�q�C�9k�<�{�qm��mR�6�Ǐ�R����^����{�y��+v7�e���k[�B��9o�=�{ͯk�̽�^Loa79G�g�i�=��d3z�v�=����īO{��B=�2�$0�R����Uۍ�~R{�}qz�yv�dJ��5N^�oݽPe��s&oL�.pգ���U��.��2c0�{�W��mW{Gݕ��[N��h���]_�yg�1�܂m�]�s�s����#٤��<g�F��t��1���w���ϻ�R�k:�[�+��>=[�������;�
�5h5<//Ə�,��>S���н������Ȇ,��y���2�ݠ�K�q_st�6ӱ#���'��~سZS@WU��yVS�"��q�s��n��i���%�����gk���;w^�}'Z�d��`�9@�rc�h��M��׀������&L��=݇j8��y�o��`{x���r]]Yo�����u;r�����3��f�^���A\h>2��&��+�Z��Z�G��y�~z� �۾��J�����5)�U�h��"����a7VV7r����	��9�v2������񲸱Sb��<p��t�sG�yD��VԵ��,�B�F����L(�D����H��4�tik�ܓ*ߞB�]�EbD^/w_Q#ق���F9!{�T�};�κx�6EIykf]y]m�yK�/�8%��ᡷ3U�r9-m����.Ǫ��Rm��5���Yus�>|�J��
��7޷���C��&	+���j�{_������5W8��������}\��ǘe��f���0�v/{Ջ}E���Y�0v 9�U�0F�v��MT�����VXq�dǄ���3�78�l�NVm�e�wgk�����2ǫ�^�i�}8��P�p�[]�4��}wz��y{\��1��u;|�<�s���=���ː����N��l��8�.�T��V.^^�Zfb�)���^>����Iy��B����Q��WJ?k�Ht	�)��M˸[����}�U�G�O��zvk<�Tz��~������ˡ����ƽ��fMB:���-#�<;"v�i�}�3-*�ոl>�Z��n��=��j9� ���թi}ſ�e�|vm�&Cr����Օ�L틅�lB7.F�̥��(�޻��s.gj7�O[p�7��1��и*Yb���PO�S�T��~뗤߄�OW�����}�����t*��g�v�]˻@�k�NL�����`V��m���:t1�=a��R����V+�y^i�w1�yޏsd�h-ge�����Wa1G������<W�sv������W�ި3�:~��9�]�eU��h��Xߟ�/A�ev��+�;ǌ�Y뎽����Nd�Əd�������Ӫ������ӯf��(_hn�[~M���E��|'3��eɔ&?��Ө����xť�o(ϵ��x�=t���=A���	�d����eŻ{|�VC��ipw3E����mJ��X����~A蓳�p�����/�6|�T�X�me�3n�z�C�ȕ��齖�WRN�z��Q�zD�����Ԗ�.��et�8�!������[Tf��Ri��{���Y4,��vNx&�>�L��;E�	�P,[{u�{ւ�+���dc����.��$q��\^#���}W]����-��'D"�T�l�͵N�kɜ_��V��w\�� ٪4�ENō�{�򳷱9L��W[�#�0�Ǯ��	�2L=�5��û��}�����V�����5�������!U�4��-'ޓ���	�{��^ѐw�?W#68�sœW<0�D8�tSw�^�O�{"�-h�ẚ}������ע?V���g�/q�X��7ޘT�󥜮D����r��Ԋ�\���F��NzT>����I��ho�I�s�t��"�3���{!k�n$�g�����V&�����s�q��Be����[��[�̞���ѐ�g��\��NcӚ�O�v����=�9*�'���=f-X��^8?�B(C}w�p�w��!4��n�O����ǩ�T�g��oM��!�Q�#t3l`f;s�>z�΂:�9�c��ޞ�=��g���o�=;*�ȼ؆��?c��Z/��c�b��~~g��\��*��q���ΐ����N[�>��M3���[�zof[TA�q��#��|N<u���/=�g*���9m�ҽi�G�axT�b���р&ž�T����:ѝ׆W�N�:9C�b�}ѻܛ��{�Қ;��M1����k�u��3�ҽ�hXa	��p֚�Q��P
1�j}u�(}�keM��hD�x���ycʓ:\\�Uz��̯r��u��	���Z2�|&w4��6���0���7����.�/^]z{:�_4>�o�=�pe[��`c�S��zk���L�������ە�}�����"��뿽g}/�m��8�uo�}N�sw����?[��y���:w�'��:r������-S�I�bOp�LT���M;��_1o�zѪ|��2b��0�0�(��W�N�>���~]��z,~�J���_�\��c�	7�Q�(�]I�ՑP��Gb�p��vW�q;Vd�z��P�9���ߒ�6n{wSJ�nZ^^L'[�Y ��Ւ�b��(����������oT3<M���.)�b��S���aS-�2Ëe�zF��4���q�����'e�f%ս��<��\��u»TT�>�ʸCw�_��p�����<eE���l�h�nRPy���녖-p<$Ӝ%go�«UsQ�t�(�q���v�ЂZ�^{�3ME��F��4/��>U��W^��%Lb��n�Ɓ\g%����OYfjua��b6���nr�OC����/���J�y�F��n1jh�wg��s�w}�W^���,�}d��j��{ʻoc�tZ��r�������o��{�Op�w��]F�u���A��
���u3U&,�]�-�~���I�Z��7����O1���9�������?W��G^�m�$_b�g���G'��E���|�e<�޽/!�'zZ�\��f��O\s��0�v<�UZ�s�*ߞ}մ���G�^��SԵjDe�^��>({()W�X�]2��k^j��G��e��1��+#����O�W^��*�5C��)�GB}ӯ:z;f��κ�����W�U����'�N68�("��.dl6|���3�?��N����_�s�0�����o�K_��y�����P_�G~�[i�	��b��8������|P:缱�e�W����!�G%{p+�h����i4��~7,d��29%r�R.;�t<u�[t���fe�ch_�5���-��%6rgF����fm[��H���w��Ӄ��f;�2��jr����gpu'��ѱ�����ݬt��{e>Gg,.T3b�U�|j�^�qj��: .�ܷ�����Fʴ��u���O�x�7n�{��r�</:�sw힧ҷ�<����y�^�4n3-�?@^�^O��_�r�U\��J�޹:�4�� ��7�`XcbGDi$c�t�q�q��D�վkv���b˃9�_{UN���cϮ���#��t�cK����/���^�)�����y�M��୳O,�=�dSe*xrE���u�F�t�n�û��NmF�|Ɯ[C���D��۴�E~�VRJ������t�g��7�#O������U��+l�~�mI�7�G2=�z~��u�d���z�7~����!.y.���Щ�����{e�pU������@;_L�_ۂ�{~�������g���<���w�x���[��g<{�u߶��U������O�fk����g��z�6!-/H�d�{*�\�Bg��ѐ�G8�}��g�ߞ�w��������7�����	3�$�Æ��.GE�}xw�F��!,sE�(���#��=���e=+itI�S*�~�RV9Y�Ǘd
A���B@��׷]䙢�V_^1KL/���̩�ɴ�8�n�'1
Ń&+���HN
'�_��s���W��¨e�sUc��V���X�#B;��:V�\0�ʔ�pɓ&�"�W�(Q.NغP����4EYJ�n��#��C�\t�q�Sr71��]9�6�9�U�8S��d6p��v�(�MM	S*%�� �޼[���ik`W"��S�Z�1��E�d�Tw�wpҴb��D�֝-��ctv��Z���jkY��o�@�Pf�
:oj��ϐ��]iMJ�'>*�F╝�sV��F�z#�����cbV���"��HnEYD;:�ɣ/�0����[3XF7B+o��z�w�tH=��{��%q��l�Q��Z�1�mѷrģ�
H�+�Ž
I^m���b�3�9�N�^�Y��jSN,�ʤu�����Ί��v9�*�tb f����a�:�X��q�k<��r�ua�*�q*��	S�MtE�K���-��;D��4��"�|S,g4G�7S�'V��5[U�-��Qih�t����u��ع��K�%4%{&�Zńu���T��zb�!	Z�h��O^Ժb�Z*�;�ёRۤmޢ&mZkk���:�K2t+v��p��0��TĢ�唻�%�>�Ս\d��up�/�k�g@Ύ%�nnܾ���7G1a��XF�m���n��j�R�v���C��=�;���u;u^�Ëe4X?���w[ՆID�:ō���֢��a|C�8��uj�/�C�a��hA��98�-��b�É�������{V�WHc�m�"�����H��/���V���"�2F���V�7�4)�\S!�Z�&ή��b*�쓲��=�r�kB�g���C�m�=�@��QY8l�#0Vu��2Vw�V���FB4�1�YN��"򝩼�1g����=��b�-�(oi�\�Sjb++R66Q��0��4�6�A�0���>�:�!��g;6�*Rl�y���ܛ�G���t5�3#���u%�	ou�*�q�K.��2������Wj���3ei�ȑ�XZ�zw�֣�NP�F2�wzfd��7���s&F�y��F�\ܻ�IH��
Q���Q���i������cyj�il(��z���6Cr�����qq�)�i�*��ʝԻ��:�|Ag�1,��:�ʼ�P&(l�1'[�+�ޓ�S� gR�aZ�=: e����ՙNV;�j�C�h�-�w`=�#j`�ge����e�4�h��T,��8�y�4�W�JgK�x�b;����:��wP�q��qv���Z�����~�@t�hi%�v�n�� ��w(�b7ҟ`�A�u7o���	k�R�l��Zy��'�b_u���YC�c�M��;U�o��$��߾���y(��lk�u�lk��w3��[��w�z����v����lZ����8�6��g��n�t��q�-.+����ָ�n
���pn�n���n�u��౎��F1�����N*8����qh�n:���=�5ڱ��0y%��I�����y��:��UGOV��c]n��w������tu��SAv�EU�bj���;��G$[:��I�wk͢�j)#Z�tUkOc[f힚�kkWm\�S%[4�:��w�S�Dy�v5Unv�(�4bM8��4�Mi�v�v����Nmb*�;��q�v�7X�ݻ� ��c�<�Qm�4Eڌ����:�lM����"�)������3�Ŏ����ڜED���Uh�Ή�<�v6�V����%Q�����"��u��N*�h���j �ۻ�ړZ��lSv�Z6;���-D]�3Y�UQV�+s�g��������v�P�I��Z��̏�i'I˺��[����Is�o��lݮM_M�*�İ&���ݏ�oհ�;̵�`3��&�`k"�:�.�5ႄ+���(3�#bί�������j�S��u�]�E� �6O�P��	8���}�g���l`�"Jm>���]By�}���Cc�?OҦ��f�OY0|JǓ'Y'�9���6�3*��x˴c����`��
 ���y��pq���~��_yR[�
�b2E��j��{�]���Jhz��'���ݾ��&�^2٭z�K7: �N=90�}�-��~0��ag�:���_e�^�t[ۺ�c=�M2Ƨ�t��*Q�Zc�#Cq�{��Po+����Z�HJ����� u$l��lV͆�ʯq�R��^tP��m�yNu�TI���;�j�9�Zk6u@�s9mD�U��fzQ�׏&o;K)[.ƆG�_���(���Ur����uP������s��$i�=ʛչW[�����|Ta	����2x�Λ(����죞Aӊq��|�rmݞR�"��$%%d˰������ۄX��3 �1��P�A�<h�����[��Lo�/ɿ�����ס�S��.no�4�k�ӷ,-�c�+Ӯ���b
�Qr���5x$N
G�e)�8���=޷J����B���(j�]�f�u=�BR�M.�/���%�Ӵ���7.rͮ���&��� ps]�$�+;��)[r�IV��<Z���W��2��Ɉ;.$�7�Y̽n����q���=)��9e5%`�#�{�*;�J���*D�9ж>�oQ�1�\L���hr����s�ޘ(w�8�<��+�%+��	�����Ѥte*����eX�5��í$0c��щP�I��l-�h/B�Ϯ+�lK�8��D3��%�#쟥i��t��2�ӽOia�7ކ3b��9���d��7 u5*����XwME� @�;#���x���˝d�+5"t�l��B�������C�L��;��<�+�f��r͎Ɩ�e,�Ⰹ:���d�qɎR���P���
�H྿�߹�,����h��_�6�n�Y���Л�
漎��u������E$U �N���%Α D�Z��t�'b��z�+�t&�ַ�'��g(����o���c�L�uO9�N�G�\"��U�����T����߽^z��q�LS��*��e�l�`0vl2$K]7�9M��H�T>9w�ߘ�
EO�[�2ᯉW��Z�p1
���T�
�2��Z��1E��YB����]1
~݋�������9�#znr(r��J]�-��gu�p��Et\jL�jÛ�'��V��y%��2fJ{P��(�,���e�l���H��C��:�;Ȋ�gx)�%��h�ls�o�Y�:�쐸���3�if7���FƩ��4.�v�n��T���
~?�����̏G],�<7ߎ�'���(�p܊�*�\]���m���M���df��� #�@ş�}fp�l��Z�.F�8�b���We�<B�£�Rt	�j�8�z���V���Y��b�n�|��}� @*e�e� ��d�f����\��L{�V�
c׆a��}k|T�j�7BA�~�S龘�\r�K
,�]�r����IE	�����]=�.�C�*��ƥ1O�QR��ʹ��*q��lT�����Bg�w�������&��3�KF>���8dˎ9j����>-�^�#4V��	&p�z{�W����lF��7��T�k��3 $��G��J�
�l�]N^���q�
�.+˚���I�/�Uj��������':���4@>�A<��l�kҤ���s�����R^���T.Ś��1�ɘ���b�C[�Z���@�&^>����Rv -7�sE�P�u���Z��W�u�jr��\�����V[�I���L��Ɨ�J=^�N�"uPK��"~���(��M��F���Zx�?8��x���5��;AV�v>���ｏl��^w��jj��Q�ն�"������䦣�F�%��Ι��;6��z �S65j� ��Ln-�V"hK�`��3n�&!YP�4��ͺΙ�>�+����|�,S�R���@c��#��[.���M��F-d: g6\��g�\S4x%T���R��<3�f��ȈQ�Ƅ�p��A鋮<+��}8�}p��dz�G�\��4s,Hnl�<�5_t����1����f�|:1c`kf5�X!}�+�j-dX���4;����vF���������d ���{h�X�C�sy�`������@����z�f�G��pt�iݝ9��;���o(V"�i��&���w]uC�o��xKܨ�#�%��6l/9��q��t�>���jҫ�R����i�,�h�s�o�=˔U�B���,��kT!f)�*/Jm��<z�P8p-�ř��@O�1�f����3:ݹƩ�s�S�m�>V0-^L������r�/�'W����C����R�lZ�˸�FM��%9aiT��Ji���N�X�7�EŴ�DY���q��>$_;�͓��y�KG�����y��jX4���QI��>�=��\AKn{1�91��޶+Ӕ�p+�c$��(1�uu���g�bDP%W'�:�]�w;y���c�f|����
�nWr�ii{�`���x}3��u��������#$� �����:iL���d_f.�����u���l��R����.�*�>u�)o���j��{RY9;l�����a�Dp׳��e�zR���q��.��4�j�4����y�EL7sN��xti'�`h���C�*8��;�&�����~8pjRZ���,T��mP�*B�}��[q��{��r�0~�z�ݖ� �4�5�!H.;ʀ�<��M��@Y��{1���NM.���\_Pbe3�3F{�V5-r��0nb�5���q��z�؝dz�lσ�iE��	S���-l���B)H�ѽK_K�e��@�"LW��g���LA;ǈ�;5K�z.��7�_x�d��G�����j��L�e�nc�$h`0���v�ɘh�;����W�͔|)���>�R�g(ш��P��{���}NP�	�h ���f�H��[υ{&���\G��P��<4�PS��c�d��3/.巌;aQ�V���h�"��9x
�������3ô2�TŌ���=�4��Щu�1)�nyL#���Q3b�Zܾ_#Hy�'U|<�U����$c����IYz��>�"�ђ)�]H)�T��jKGQ��b�c�'u^txh[�,֑�Gm��7k��%I���O��b�k��ϝw��O�}t[��i��ՃrIo-��t3m3����'*IZ�oFI�sca��
o^7L�����W��hj��k<�^�z�n�F�ww�+�<���ߦB���'3�T,Y��Z]�����s�1_b�n�`�Չk�6Fh�\��P &���*4�;��`&���`GD�r^Zz��)�_��Q�s����;+5)O]x�MSÏM��R�?�b��By�m�!��O0nP���Tuz4(�NNj�{>ɂ�u�%�>����W��ҙ�M��I�~ǲ�{e�F0��`o�~�-t�k&]��%<��ADR}��b�b5TE��O��b·��7P��q]�#��W��6�� V�dns�hܬ�S�R}���ʴ��e�7�d!0��`rJZF�	�Q�ʀ�ޕ>;^Y��}��8��P{��k���c;��V3�P	�k���{���b),Չ#���N8�㼟�TY��4uF��z�;e����}�^��OB	�T	T�m���	�ֶ|�C��5a�������z�ͭ4�c۔"���Tg�^���^4%��������[C9�P��{��.��7
jh-����_H0�������d,��sH�ޞ4$8�G�ϳ�`%�7$u1��z&K}W�1gH���ƶ����mn�@�	�U�)k���c�ؾT�ϝd��坯���u��?G<���3�aO_;�+��j��/۬;��������˫גv֟�<����L��#u�-Q�3kv������I��޻WĬ[)��g��i���`�m��Y֧2RP�sk;��%���'j�gFC��_U]����2��=3��ީ�2���u��0w����g#O9��Z�=�;��e�U�����^&Y���4�*�ERs�LLY�,����1f򑝞���,�{{����/J,�[�G!��*y��|�:�aN�~�W9>jw����]5�뮋:�\Z}��۽U
�d0\�n��9ȓo��.qP���xDz�>�<r"_[��*˞n�lQ��{ˁj��ث&,���j�M|S�MI��kyB���i��Ǔ���	�!Z�D�k�����|�c1g$���z%*�G��YS��:%�1.�k�b�OخEc{n��xv1d��Q���B�vT7����c}fpЕ�P�r���ص��%�9�E�4���B���\���}�d��D�Ӟ�Xx"pS9�'�T�=K�˫$��1�Ν�7����M�N����p�:s3��y<S~�n��~�b}7�ˎZ��0Ȅ��_J�=�7��D����¯X����:�1���:�C��޴���b���=L��=v�r�
.D��w鴩Da����wu#9�f��]L��)�"��лdÉ ݪ���,���� Z��pN�?��8��a&%���k�����-��e��Ga��\��U�/
u��e�!����O�,�=8��!��s��*��6��۫[h;���҇f�w0KqlV�)��o73/5դt�����V�M\q٥-Z��&��pv�\��j��u��aYX�.�����z� =7�|{y����5Bl�r��&`�WQ�]��J�V����Gr9�!�ۇ/�؍���.�N��<�'����P4A^ �N7�}3׮������&ԋEO>F�ֲ+2z�f��?#���9��Q�b�5^�@�lJ��@Pv7�ae�\Ӭ��۟0t������r��9t��$�Z޼UsF=	5%�9� ;�@f��ͯN���N��$|tW�m�yġ>X�yRz���W��-F b��s=٤%t����wT+���������G\�>O�,x���!�sg<��C@���*�4���`�s,Hnl��&Ե0�5��#։����S�Y��`��c�9J	��q~ņ��jJ27!�J��x�bD�>��l��<��x&v��C}�n8!��<��N^&�C�.����]W��o�&��AmU9��+�3�j��.`}}��?3���۳U���8q�����5�g��@*}Y5��Цٱ�HȨ3P�bA�o&����:�V7��
 bʈ{8��,�*�����"�x�� =Mgo�o@�7��@i���#���aN�},��&TE(�w��[�u�5i;Eh"��A�-EoL�+w' ��ZV�p[%Ϋ7��BC��I���Vn0%mv0A�Tޟʉ��@l$�:]�ms;S���_}��U���s[�Y��@�'XW��p%Tȹ��>�ɲ'�/��N�~K��8�>��������(��т	�)��6A���:MJ茎�N�`�޺,N���W>ŷ���g%P�k��
VN���i���3^�Sۯ_�ǶQ�R�x����"0��]��sJ����'�b~n������q�{Ǣ_�$Ono���)��]EGڒ��:�gٜ��<v�P%W'��	~H�@J˶W��2Z2�ד��d�x\��ey6�# �����}O���ウ[�^����T�kS�xv�)�n�WW^a1̖�P[��vG�� (	���+�yP�<��x���O�Ck���f	�%)�������ʒs�[,���j�ƫZ��˱����U���_x���
ˢ٬�Y���mnu�J�>T���v�f���OۅP��f�$Գ�j���!�TЬs���+��[�j��<!¾菈5���n{;��~cY��8��dXܔⱫ�z,A��#��˃^pνu��̀�hj����.0��fù�b��w0mq,0�v�X���i�17A܉����a@!��w�i�@%+O�a�--�5��gy�Z��m����c�X\픹Po0��ʸ�u"�ٺ�O	��>��'H8�W^*)������@��.�7��pa{JE�+�l8��f<?Ͼ���㙯&>����;M��E�W�'C�P��������&v�'��k1#kw{�Z�q��n�_�V����t�>c�I�zԅ=�j�ܩ-t�:�!&�p��LQV�����l�>V�Rs�������ۉ�/.Q�+�^׾�_ݱ
y��	�^��yʑu�Ɇ�X�bV����;�/Za��ʠ[�6��t4҉bȫ�9�7���\�(3h�!+��wǼdl�X�'1��i�V1/�I������i�ېLSy2O��Si�l	l�T�{�UV6�ӛҔ ׾m��c�[�W6rh��w����w#�_a��8�B�\5_�TZrsU�V�}V{l�fM�h��G�rU{c�*0��g��-m�' �θ(�(�����}k3�}<��W�'�9n�h�sZ�5?Z��2.��u��X�5���,C�*(>�PY�[���B��˴��?]�K~�5wӾ��G��?g�+7��=r?#�l!��Uy����w��9Xܣ��bSe�o�©�<�SvGI�\t�N���u�c�lE%��%$vF�@�|�ߧ���~�w������|||}B�N�L�Tvh̤��ZUb� � ���t�f%�˅���6�U8v���V��ޱ�Y]�ƵҪˡ���s�˛���M��P�i��ܸ�C.�n�v�}����J�-^��3�3�ˬ�z�����A�l<[5���k�S۠+����c3"�3[�x��\T�S�iH��S�=�U�3Q���'���t�G2E�#q��pҙ��E�v��C|��ż>[L�-ݣv����b̍�r�&L;d�'�Nk���B��u�Ҍ��^qM0���zC��s��F�5��P(\��}�:�vki�o[;بwUصt�;�����;��Fm�'c9\��m�nl,���R�hqˈ�A���ɎS � ����[�Sz�2���#�'{q�*`W�i����1�b�LNnK��S�j�W#2���Dte B�����vbY''�(����jR6��鋨����$l����9jZs�Ζ~�r���ގ���9rfe�7yk[v��#�H�."b�EE�-�UW#J=�jj�b;ٲ���QA3��u
gC�3Fu4vy�t�;����:r�����2�Q�����C�$�kኸ��̫��2i)L-���P#k�C�6�q���F����%��I8^ w��ז�(�����U�<9��ѸB���ś]�����چE��W�WJ�o8:�F*��t5�������Z⫙鳹�j��r�Z���'^f��mv��L;�,N�jk�a5�s����A3>a3���������I�F�e�N�gK�qm�"FnNj%�ҹ�����~ĥ׿u�ͥ���QK���}�vz���Z���h������3����u��m���*��0ӈ[�޺4�9#/gL6�^;�B4Ȳr����VqlT��Й9c�"Ӟ�6n�S`�@���`�0�^U�ǓfD�ss+L
�x�������'}�*�F�ǻM�죍��0�ѩ��ʯf�*C�c���#�� ;�{�-GzI8���S�#��5t���oT�ҝ���q^Ѓ�G˅╢�ɛ��ah��S���=��P��h��.���������M�
��"�O��ׇ�5��Q����3m;����I[��{�֦ywm̂V�C+^��*�5�x��(-UmR3������k���i�n��c��֕͡�l��͍\�N��4���|�9���o&��o+��/A���P䃫��C���oKS9�W\������ԇ����)���
Q]��1�ubWTv��)��S�F��v>�&FA�WgSI�;s�q�R�ٛ-9���MΑ�������U٣OC�m���$o/A���0�����/�#{pC��W]�&�Ѩ�OkJﮌ�9nS4�����o(�[r�Z��ع�sOniV\��n=�����W{C����	][b��vHD��F��w:�fj��=S%tC�����̏�].s���!�J��WsԗB6�h���]�r��m��`�+/�6�=��OmB���!"��4��4d?��q���mX�:�����KmT����kQ["-�j�;j�f+Q��l`�*�kmQLlDd�5��b�����l��v9��剈 'cEU��:�bu�#`�h�Z
��]js�&�k�N�;mU5��<��UE4EACh��[j;`�4m�����TEZ��E�v��5�kk�mQ�MS�$�ٶ4�6�A��E�SUcj#Zu�4P[V�$���q�A�sA4t�ը5�6�mLwm�+�5ET1���jF*6MP[i-�j-�%X�Dl�6q�Dljd�Qj��k��s�* �Wv*	��1m�J��"6m��X�b�lI����h�Q&��3%1k4�U5�b"&��lb*J�"j�h��~w�~&�)nx��+r�M64!��`
](�p�5���0Y�<0\h�ⶓ\�:͹,\r<�֛�j��Q3Y��M�%����~��`=ZV!�L�@}�P\n��C�;���X�0�[<�^���=׹MsVk+���lj�z��9����:���Y�K�P�W��<�ƇX.g((	��.z�%UsȦ�1j)��q�4N��o��Lyt�J����`0Ze�9���23��b涇w��ۼœ���T^\��6Ôt�q^��*Z�R�2��i�Fl_*��d�����5�^��E�#�ׁ�m���7)~��T�(�3�r�z"�5��hP'T��}"�,EŞk�V����@~�r���3�G�O�S��[��B��N���&[���s���}�����U��@�֩FNPjV�joFC#x�����ڼ/rB��f���e.Q�K�j!t�;ϹM��w�9'1�^fg�(�ٍ2'�{�0%������*�I1�^���p��W��r~3��XE��î�;��#��B}P�oG�0�;k��%8��)��Y>�L���籊(&ѢOOdva�!���&'��W*�q{�0­ݎ��-�M��P�	�űf�S�Y��{�I����=�b�;܁��2'�om��1[S�)����x�ʺ�[ʲ`�D�pd�mn�<'G����l���b�3�sq#�Wb�V���X��:�Pα�:
egi������TL��'P�A�P�]hT�X��7Z;H�ْ��mq�3{v*2���H���Cb����}���}��y��Yܯ�>|L�c�ס噕M��+e��(��2D�_y���x5ջ#�ǉ�l� �랴�+덊�^�:�K���6T�r�؟�߲��蛘��.9j�FY|�<��_��ewlmP���݃6���}��̦�Ԧ)��*S#����h���!�+��.�я���6ټX؄�sez`&%�=yɨ]ᓮR�a����+�"q����U�S�'��.��5^��r�|��F�9s���(�i��e�d�R�7g��N���%����=g�N�9�q+9�1l��j�.���*�q�q��LƵ뭛.�t�� �%`��)�2k��Y��*M΃����ގ*���Q�]�@x�{��@]�
A�dH���\Im7Zi�$���\,����}/&�1����F�
�[��L���:D{9P�@�(��Ij�,7�:���)��Y�MO��锋:o��=�u��{�/�n��^�):��O����)��WQ�hs=_oZ���e	��B'!��P�	̏b���K��C�X�H�?76A��h�Z #��a{>�Zr}Kf�-z%��[t�m\C�X���!��pt�mڥ��54�S�,Է5 M��mk:�f����r��-`C����g`�uU�T�*O�����iwS+�l`N��Cp�H�8�g9T΁3�+0�����6���b6���T�t8�߀ xs��-I��(��xl��a0v��3*��mF7Pݙkm͂Ɯ�a7 �����o��P'���W�說#G�4?W���(��?lf�#֠�3a�U�^�:lg�3� ���N�BT���ru� ����S�ѥ����EစB����s�hQx�C=�TM9M9���x�/a��z�[���&�׊̱w�*!�X��A,�M��W��*�<�8T�âu� �:�ݑ��%�wM�|USs��۩fV0��nr�E��mk�;!�2&\��v�~#�kG�x*#�.���1)�����(���u����2�[l�~N�n!���ͽ��qlI�E�˶�In��_���W8>sJ�|���t\�G�]q�' ��������b�$/�Z�<����$�@�t����b�P���e��1���;У&jjI"K]���@9��� �3��~wx �
|��Lq�G�����;7��l�w�~����&;7|&�>/�/Ck�<�C��.Q��w�(����w�����~���iy_\lu���C����u�>�{x%�7"�K.�G��*�e�g�{L�-�9ƕt�q}h�	�؊Ƽs ŗzh�<�qĪ�1V�a��.b���ɛ�\CZl(w;��˚�|6��C���a�;�q��>��<<>o{õo.&�\��E#V����Ag��W��]��N�Gx�<M`�Ǽ��o�i�^dgb���	��^\�[�LJ<�T�V��Uɔ~g~�3|R��@�z]�\��������m���F3�Wf�,\/d��Ҩ�t����\$�g�yg�v�J��,L�d^A�8]ϖȱ>�4�)��<���U�-i�߽@���ȏM���3G�	C<�a��pw{)��@-�ˏ]ɜ��E5���<������Xc�7�-��僔��BPrJ�Pf\y�������ݶ���W]��yq����{ݾ[��o���8$Q�֤�P9�CUʒ�P�V@�1q�PQ�_Y�&�L(y�����aS	��5~@�
�O�7�5?A�'��pD�qq�R�,���ir�]wf�W��w��f�=z�5��}�®��WB�k΄5{֢Y6�-�=���qp��yƩz�L+�����n��;6�{#hDO"o�x��B&�u���<�:�TRs~�"�J���q�ID�k>fc��'�[?W؈ہ~5�P�5-�;@dp.~�O+��!k��cq?xUQ%d� ����'+<�eN��owM驔�s��YP�j�n��D�X,��T��gQ��-�y�e3Q3nbSynw� :G����T���z�J��D2Tc�7éR�$������a�if�d7{>9t�G�v+ˀ�-w;|�ٻ�ϵ�����Sr�x�<���/P3�U�9�s�_�8��`��/"��d�2t܅�n�ϥݪ=�AK���͆�H�]I��u�X��_��P=��F!�)��^��Y�8s�׺�Eu'�v����>]�Z ;�&�ܢ�G�~}l���7�����L��=w*��,�ۺ�]XѺ֞[�!R%>a���Py���i/a#%����~B����C˷A<O�0Dg��l��沉�/&�S#c�ץ�:Ob���Gq�v8�L6��4�[>{�S\Ն���ݍt��#S��A�γ!4�(�f�=2�ɪ\v��<��4:���;Q�Lh,�Pǃ}� G�:۲rv��A��{)��X+U��<`$N@�";��@k�6��Nu�Ŀ�\rLr�8�z�kjó�T�ǈ�].��ΰʎ5��|]v���T����D*Z�����ی�M���gs�yG9}��"cC�//	��>�ĩ�Q�|���0�R���	�+="!Ɛ�w{.�����ݛ9��Rrf��}ח�Tpj�!�d���
,�;�+�Tw����N�I}�g��n|�F^@R6�e�	 ��/��7(^���ʛ�nD�^Z����2!��IL�
�zb@��Mda�;.�V�~���\z���T���[���\�Y?�`Ӡ�=�Z_�E�����Bܫň����4�� {�����f"�s��ӎ)�׹#�����e/���lr�-k���=�n�-~$WTK��ۼ�"��2xy^�k��b#ǆߪ6���{��yЃ({O)�+�9w�z?�Dت�*���_�ۘ� v��s@\�P*_q���5�VT�����{���2�ƹ�׷�mGt��),�zL�8�VT0��v�O~�Y�0[p��`V����'��N�#oe���yݎ8�b7�8Ǐr�ׯ���c�Vʯ�jB����K�S;St�p�J��d��2�q��9H8duHf�7�I{fP,`Oǟ�%>�~��}79q�T�0�ӸIa�e�UA��`�Y�O�^�_b����B��&�jS�T�G��my)Z�(�	W�y�s8�w�Z��1�n=N��Q�1�� �yM��|�	��ڈ�[����`��Ƞ�y�-	�2"X�;���՞>*��"�!��Z}bE}3��s0����ƅQ*���].�s&)N���sY��m&��i����x�����x��EV�(�������}qB�:|~�c|]���q^Z�}������5�ɨfd�@#��!I��:����GQo�j�"0���h���7�,�j.���(��r�U��$��?V	u�hq�Yܼ�[��a��4}�ڋ��cA諏[�g9n��bz.(�&ﺎ}���| �������
��vw����e>EZ�g�j�Mw��yW�D���G�P;��|��W����]Y����<��te��;�yp�{ӆ3??7�?Jdz~�@o��GT'��/A�=SV�Ú���RbQ�Ȱl�}{����i]��3��z�-�3_/T��tIZ���ͭ�|}{}Q��i����w�D��hD�sYIb����=�>iybL�bG	����'�4��Y��s��.8��Z�n�a��Lk���ʥ8�د���g���P�k��V1���^��_9��f�M�	��uH��_(��W��B2=j���k擾~���{z�I�/)Bfz��80$��ˮ�P�V�T����D)�Ia���fW9�P�QV����_���g7��4�UݵO��ɲ��%���h��6~����cʈS��I�'1`J�����nc9	�7T��#z�ӽ�4]g�9C"G�2ϵ���v8���VA�o*������T�\���Oع�n�&/�L�_{�*.���Gy*��ؕ[r�8���2`�-熾s����ӫ!cQ�)U��k�N�]��6�.w��K/r�Ml���x>�ٷ��3
1���F��R��D�-Z���i!�ސ��,@��9��=�]v��U�t�zxr.m|j�ӽ칖����pFhY�H�Tʎ�k�x � ���;C34�*ak\��8�����;�4�C=C 3_x�|@��mC���������16�ŗ�a����Tډ��Z��r|��3�؈���=��2%��R�oW���Hw7����'Pf&�[#E(g��W΃�IN�C�p�V��ނ��7��A\G�X����^�[�0.�T�Uړ�(Χ�K�si����8���q�8��;�	�ׁ����!�qyP���b�/pA7\�h�]omY
�޼l�A�U��G���F������>�=ҁG���'����w����W��S�|��+y.��`�����>�g��"2���H�R��;���S\v��y�Q���Ǥ3J�A���0v;�4HQ��1��r�����	��wH���[�fl���u�6���{���
"}�0a�ɒ��̗�����a<�=�H:���;����NC�gnT��"b܎�	�. 3U	��Zq(5��A���f��a����y�eI0S'�U_g�����"�y�#�>k��,��ԅ��MO*K�
p/����N>��8&Y3�ܲw�ѫvpqD�_��ڔ�)u唯�=kxj�8�ڊhy��W���U�.��t��c�}�orX�ӹFb�t��J��k��׻�{���Z����Xͽ�\�vq��&�)��i��TR%V�z��:p����t�p<�ɘwϨD}�<�>o�<+�&��QD+���whu��Sl��P�2�⒔ͯId�e��PD�qq?t�
��B�[�`�ě=T�[��K�7e��"�e��K�MHt;�^���f��Y��y��u����k��t�o�	�<\5O�h���u�d4��fFR�$�XЃwO�z���:�	�N��TRs�Ȧ�E�q:EP�u����R_ݙ;+5,N��|�+6��;_n�7�x�
��@�9x��r㰣Y����j�6u�b�}�g������cOu�f{W鐕�����|G�r�{̂wu^��^ ���|sc���w�XQ�i���U���$�eA��w���(>I�y�Zڥ�ﶳ�M�b��SSU��d/L�W��Iu��{�E��� 7��,{*�`�#L��=�˷�[�cNuΎwn�1*y=�S�J�����d˜�M%�$d��1�)�+��;{�Z��<c�5i_�wL�Mh$�4�Aad2$GC����ؾU�C����v�8�{?+����U�G��:F�y˪��_1�M,&��qR
mxЗ�+�������3���F�1a�T�q�.ف�)�Ή�t\u�2���W���Ũ�'9��
��TKh�'>�!�ߛW�«�P���)�޹�r��e�9lO_Y~�g<�����:H�ʛQ�>�}@α\lY�٬��t����޷�l)����k�go��p�s���^�g�z��3�p���x{� &�����rHE��š���j�a�=`��'�H�������_g����Q;������A�7�5��1�;��y�W���Ԫ�׏N�J��~?*!-[��\�˳�Z+���{׳ߺY2u��}=�tO+䷽(�2�f�F�R��z�ק�"6��J�av���y�=��vC��8�W�c�#2&�C�A�N'�G�L|��:qj'ɩ&n�-����9�)�K�U�Q�o$7�0��A������"Z�t�;����0L�2�|���ul<2ڇ�T"�>`L	��7.���@��1J��̃(sJ)9ZH�ƨ��S�&f���v�w��z�8���(�똅Ҫ���_P����q	>��.5����IA$�HK�j�C�ͧ;P'5*���M԰яL��E��i��hb��[�i�vNI\ɴW=�v�ި�|�_2o��S���,p%>D��b�S��c�VʬZ��+2Dǜ�U�|=.gkpC-[u�����2�ΏPf��(��B�V^)��ħ�*�X���ڋ��{}����z�^�_�����=�o������{sa�R�ٍ�$�mb�`�3v�mN�� ��۠8q��S�n��;�ħ]/�b���rEWSt��J6)�_v&�![�f��iɬoe�t�K��aM��ݻ�{n���CI�&k�O��ٵJ���C^��t�np����59�g+���vI����\���ъV,�dT���۠l1�J��7q�>'�R˭���u^v�W+M҃�U���ۡ��gv�-e�E�� 1�Ji�5�ܷ4��X��
��"�PW�)P�f�Vg�����
���q3��]�� ^�͟Bzq�%A�r����P��×ۤM���R�h
)mrː<y_3��Sʅ/)���"�W��Y���Y\*�bL$�溍i5n�v�J�,�%�%GD���k��ӊ�����W#�B-i_@i�[X��G�5e&�C�ؾ<���F��O\�{���u��u��������c+MlYȩ�{�j}t��b��%�������ǘ*;��vxՊ�C�r�#:��|HGv�N�R?k����n�L�-(3hnn��dV6֮�ZŦŲ�{tvR�xU��~�%�R
�fH�V�j<;z�X�,�/]s�9��y�i�-F��Z�mKb��0>�c���i���RKx�W���zI�9^�����keZ6E��I���ق�T�}����Ŝc��2R�ؕ�VH� \�/�ut*7��NP�"q9rc��VrjԲ�l�U��	�wS���;u����D�t�G��}҇�w�����)29���k&�'-�|����N�z{��Y�[	�EW;Y����i��0�k1�\h�ܺF�*ە;7��T17[���� �[��U�u��"���*�ஶ��2�^ٺ��/5�,��CsR��Z�/���"���ۺ2�_4H��kZ��u�Q��1���.J,�ʷFvH��x4��H��Б9�cib�uK��L��#Wa�E��u�b*K���W�ɻ�/u	&E2�:����2h�^�e�:��J��z&��I�c�J����4/rQ���R�sk�+,RⲶk�:s�WnN8���%�+�̒P� wX���9� }-oj�dq�xl:�(@vQ����+CM�sJjΖ��WV{�m�*ʠVn���u��ʛ��=�zvAV�K����s���X�O6h̥�(ݑ��h��a�:~ѕ�K~{�=an�B^w
})@M,�T`�yMl�+��%
�����V��N�/8�V���҅E����Ϣd�`�Ե�c�k�< d��+�|M�S��uzQm���nܬ�']l����3m	+��n���ʃwn��j�Z���x�6��l5���r�4�HI�w?�]�!ѻ������X�Z���+�e'C�ssj�QҮ��+�Z��*?����/�W���j�Q��10UTi�"������mT��lf���1m�������kPKSF��%AT�LM]���kZ��l֍5'mՍEkEQ��5ml�"�m�TF�kq�g�MM���6؍�DTZ�C�6�b-�b0ES�b����61Eh��6)�TP�M1���j`�Ί*��5�F+Q��Vٱ�F٢)��lh�j�*66�D;b*�k�kTV-0Uk;:���l���[EE3���k�FƫX�����[b���mCQbuSQZi�ӆ*j:ڧb6���gc�J����b��ULCU6���V�ڱDM$4AkUDX�Z"
���l�b3�DF؂Jh��V�D�m��5:�&*
1�
��@���l\����5�)�^�Ի��A��{�\��{y��D?p�f=6 kK�/k&�Ǯ�ӝ��9R�H�^����1�e�q�2��_�����0� y�n��d'��o�C�jz��7'�b����B��S#���>i��^�]�W@�Z��~PL\v2����]�X���ON�W�#_���_}�u'b��B�Nx�o��?EV�N���.�.��D<�)���AF I\#OHKW1���G� ��b�U)q���'�
rw+����jV��!o��琠��5�A�J�� ���ɘֽu QqG}���Q���;a�I�f�����*���|7��f�H4O��V���(w�jt	]^TW��?�w�R]��4�qߺ^�� H��S^lK(IU�@3z���5��\O��J>���|u���C��Ż��**Єk"�x�d���[,��V��ҺϠgCށd�R�/T��Gɑ��G&�G��^۲�s��F(z3�L�O����32\*���0v��H�����1�se�f�UȰn�aY��:}cX��N��|�8�د�Ԭ�n_�������&�Фg ݕ?uNS<�Uw��N��b4_z�ȑ��)�_X��-�ƽn����������� -��;M��\����P��Mk)LѴ�ucR�j����:.�Mj�\�t�5e��Z������Bb����.�{��R�Q�ޛF֎�B�\�V6��1ζ��i��U��2"}g�v�U��踓\�b���1�O�wm����o =��=��k�<S�"�߇�Ji���n��&ނ�y^ŕ���<8e�8SϷf�[?>z��=�舣ց�B�ߵ�v�X��*X�b�/-͟���X�Ǖ��O���b+�^z'���Y�wg�Ԩ>�����<���1��&!7b	U2.uE6�̬a^*/&��ﻞA0�5E��U�ۭgC	a�4ܻeL˞����=!������S�<�<{y����4�5����135��=Vp�S�lK��a�-�
�mj��� &�-��ƑqniQOrz;Y��tD�b�f�uwe�|e��Su�Z��*@,�\�W�4��D��i鉏?ٝ����
9=U:1!k�=M���B��{��O���]�0�^<�:�)��Q�$��ի��bT	=��tt;6��E���U-iƹ��Q�أ�-8�˶סw�|��-�V��>��L�L{ъ��\�[�k(�4���J�nttܯ,�;T�֯qh����a�s3vUF��]h?g�ÇN���䉂v=ʥ%�#��ܙLd����'���`���[Rf�����2��sTB��v��݂.xH�`S� �T�7;��9S�B.�k&�K�Z�Im޾ȨGƁ�����bVeһ:,����G�[�	WV��!���S�:�NjA��v�����K'��m�ݺYI�m��@ױuLG_�]��Q�^!����^^��I��#��N�����a�Z�ͫe������(%*4 �@��w*rxw�y��.�7�?0OQ̻�,$C�!F�ls}��q������(��2&�YV����@�W�B>R��"3Р1P��A�c🙬��dDg���X2+��m�T85�؎a���G4y�����H��SA`�U����t �J��������s5W�BVC������@*d
j�@d͇�rH�֧���X9RZ���tqT!��/��9M�r���Tҩצ��uy5��w��^��9Af�Բj>�}�n㜘���yB��[%5��);rNC�#\İ7�!�2jA��\���&�)D���92ۀ��k�wy�%)��<�f;��y��f��	�;��Q
���Z��V�P4#���^S�|O)�w�\u��k2
h���P-�9�\���{pi��������ׇ�Ⱦs�R�/�=�hW$�/^)86�E��jY�U��ŧ �*��8�X�뗗��e�|apSO�2}�q��X���|�{��u>���h��s��az��3i��H:������1���2]�ǰ��_���y��&�ň�N+c6�����kJ�5�u�����KL�-f�9N����f Y�j%<�N(e'Y��*���N._qn���.����2�WZ!��5]�Л�U2p����5�rc5{l�Z8��a�+�������0 {�
��(<���+ 7��2i�Ɨn¦[I�E�2�r1qѭ�Gl���w�3�n��ʃ�/�F���1}Y(b���М��� _)��d��˔�^�2Yk�������1��(�>�Y@���w^�I0"0.a�x�~t^Zu�;M�0ő�s�kg�~��\=�ie[�٬�'�gA�����,+`���6��C�|�MT3�>�i��)��Iډ�����/��'�>)uZ���u��"r>+y# d>0^/Z������6�Y�{2w�Gr����!��¬�p���{9���.,tP��C�R�PP�	�F#b���{�.�+0�Sz��+,��b��"ϫv~���wyg�~��?����_œ��P�y��^4���vk�5��e��ܖ[@X����wx��q8��E�!��*y��x�!\"��g��y��:�d(~U������N��*���Bp�e)w�VH��΅6���s
I���`2f��u�ٸxiP����	@�n]G[��S	��{Ѓ({���ퟰd��S�;V�a[�p��z�k |B�On�њ�2D�D%���҃<�-�v��p�1�5��S������o�W!�=_��Z'^��j=���3h:J���BCs� ��f���Gl!�]��Ɋ�b�㧶�5����` ީ�O���mB�F\�Gl_g��	kU}P���3�>����	+��<��v��j�K��𹊄ZY{:5�>��ز��[�]��*�H�߁�?F���^e|;OeĨ3}��ܚ'��1@.�mj��E��.|�T�`b�z��2��}��$��2E�M.]k^��[[1-Jr�wdpm����T�0���,y��S�Vn�������pm'�أ{/��m�j�aDa���T���w+���2���L(R���)������&�>�I�����=/��-�uM � |��7��<�/95�2u��\�A��<2@B4��m�5�:�5Sw'2�O��l�5�QPHkOBZ�虏5�_v�����;�Uʥ�fջQ�g��̤e� I�OV���XJp��͒���r�CE|WL�yT�k^����钬���9欅%��x��J�U�渏44gyX^2�E��U(��)�*��"kY���:_��.;]'���9
�6�7\cK�񯗨J>퀊���T碳\k���%�o:�:�P��_-L�U|���8,<��Z��F�J�zMi��.�QQV޹�}�FY����F��m_�s��8S��MS땮��l���q�qxrS|��z�qY@	'u(����ǝ	�Z������2;gf��������=�o <��y�������{�/+3CTn'�=䈑9?�v/�'���:ү�O[4�������JWI�VŽ�8;�ȑ�
�Y�cq3���g���Ǜ��\D��Q�#2��旕'���K�,�����ㇶ�(�X��� ���Ax������j���H߾UW�WU��wj��+��nl'���QA��/x��]�����;�[��As��:7��	xN7�v���@jl�=m*���ܒ��2��ߦN;|%�y�5��0��U;��G�v+EP�!W�
�T�����]M�8�	��&J�=dO��J�k�⥓��O��q��̱v1dH��w�4/̌+�? ��L�ؾ���|mס.��VH!��m�%��2Ϸ�/����y��,{r�{�sa]!}�-)��������}�hs���^e��܆�cŃ磕"��%9a`����κ��4�Q���;z�j�'\�����<���ey�;�-���x�]ޗ�
�!;�����pE�E�C����rz"���\s���\n\AR�m Tx�wO�|��q,X{M��lj(���d4>���/m�˖dx'ċ�񮺝�jI�V�r�"�;��Pe�=}��uAB��/��Mg�sق��͗`Y�ECs{3s��n�Qx3�z[�y`��f��/AF�V�~.^SWN�g��fl��|��p�g7E�\��&�o�:(�_)��;� ������
%*� ��=��w�>���F�3�jv��V�ۮj��8���T:�ڲ�H�Ԕ��@)��Q�o}�Z�;����웼�"�vj��^�L�����T���8���cǌ�b���j��ߩ$��a��i�_�n���a3ѾU*Zfm���{�?��V�[�����6xv#�vy�]����L�ػ�:�,�'�Ozߏ�Ҡ�W�⦧'��]���/�,:�r�D{=;�𝡇����6g� MKC�;�mu"!�c�`�v�0*B�/�c�9��P`c.{\�B#z��S�Ʊt��I���Q|s�O�!�8�pw�����P�8�3a�`1��I;�k��>�A��8�vy��"������Rj��-2 JIW�˂��iCK�u����oc*r�SB��F}�3*��۽�F(7,�rH���s����%������y�c�)�P���x�ʀ����@Gg�����E��T��9�亭��v��s�DNf5ai=X")��ԝޥЇ�yzEЌ�L��H)�dԃCz%k߳�M@Z�b�Ǔ���C��y���r��&�o�p�[A�J��S⌺ïk7w#�9�:�6��4_$+0v�:E���h�������Wv
��z��/i��Fl�������".�Q�X Z}A}�x̸��U�~_W�<��7�B�d�p6�9cWǧ!ᭁ}����F%ґ�0.����=����]��ܶ���C�̖����e�*E6�3����v_5�]hp4�;�W�)f�#�E�a��9b�������r�9�b3���2ik�Qi�����,�a�ME����XgƏ5�)��d��iDd�ғ�i���
��N�׽Ʃ���I�q&��KP�u7@�����`�&KǓl�-��9З�ɦ���K��0��.u�n}��zX�$r�\���,g�azDT�Ud=���]u��S�R� �g���0�sT-�����M%�ș,����m�u3J�iWg*����.ҧ��"�#A���x���<�Z)W+��B���#-ƕ�&��9j{��0������������|y����33��������.6�cJ|;����i�΂��%��:EfB��W����#A��Us�J,3����'#ⷒ2�ύ		��n{��H�Uq�<^��YM��bf��x���1�>��L�B�qC���z튇��!���Mɸk:���^Ⱥ�B��>Ϳb�*��vx����� @R�6t��)@����S�8oI��8J>;[H������}���=��mC���{��*�bԕԘFr��Î�K��4.[S04@���<��[��MΜ�\�yA�1�;}�z��!�k�W� =��xyF�GzKK�!��d3cn�����3��a�g;�&Y�2U	����l�V9JW�#rv�k��}��z؋L,�LY�+��zo"���w��<O}ИTNS�ܒ��b��<7Ӂ����=o�M����'U�.��Uo��+1/.�n��U�ʯ8`����s��K�k7���Y׾�����!A����Dz�T.�1\�Pm���)��)z��Z��:̐�8��΍$���������NhF�<��C纡�my�/[>�� �~*X��t1p��.�T�zN�5��&\�1E'�Ķ�v;�Ucʂ&�~�~�Y�=?P=ه�5�:�a���A�l2f�t������K�w�|�͡Z�;����rV��R�I�i<ᅵ׽�/�zB��ס.�.���G���i��^�̢�<��ؗ:��Q������e�1P�<#�{����t�ۑo�0�z�^���ͼ�qjC�$��M���*Q~�V�i����1�E�K��G_z}�.K�'T�Т0�	xM�0qz�y��ɤU�F\~�<RpA���Ә�1C��Ld��0z��vơ���i�Aͺ.{��<��y0�<.��#n�*�\�dT��3FP��Ѡ�n>I���P=pi-,�g)�]&Bj�\X��oO���]ڤ��D�w�^�ɫ?쏮�\0���bF?mMpǮ�уp~x|����{��{������7��-e���ae�*aݱ��	lW�� �4���ؖK0)�)͊��+6̢�ݸ��.��b6�Α�{��qٻ�O~����8\R��~z� ��( � �	��u*I{�k�n.o1��/��5��}��+d�oW�:�n��EQ��e���b��.����m{�����ɫ���9�a0r8�7��1cS����q��s[�&���Ԗ���,TD�b_J���n����5��8�?H���U(��O����w&�D�]`�x�y
'r`h��X.�����;��/����IK(O��1���lr"D��!��m��3�����Ҵ��ord5Q�=qkGRp�{�H"I� ��Mj�酩Ј��r<B8�������W3U��~zJ����{����; Lir��<�"�>���'�G=I1�|lE���	������,��ߟ��3I���=��g0��;����
�u�iu&}�"�' ,=ۡc����P����;�Q�-�E]tt�Y�3c���9-;���أ��߬^9��Lz3��������_������A�^؍/ڞq�W#/�vv��{n=�p]�b;�Z�lu���x��}����6��X�ن����6é8$��77l� ����R�l����=\�<*J�ۦ�-����{s�Il��*�tv�RSA��)�vVR�l���ym�岊ӋJԇ2�N����w̵��1�;`�Q�u3E�ߥ��@�[S@�W��:�n!��L8�6hG�^�Y�w�"I���3��釦'�/fX!�5f��7�ú�xu��}R��1O�����\imE��X5��9w��)�����Eۻ�������z%�k-�+�O�7�k��Ɓ�0�,f����s���]m}�'�hlJ�
�Y�LnK��n��u�H���x���5QQ���y��&P�+��;�P�qn^�ڑ8���V�;#��I!O:�݋�vK���*��N.�s�r��ʀ.���I?��T����r:X�d�5<�>��1��	��V���Ƿ�$gx���;	�N�,��<r���2nqrS�wfVk�v��5���]��In�tk	�i�(�>�r����6e�e<:��%�pL�R�Wg	|������yQ��y��ݥ ��O-�(�ΰ�����Jj�oZ����g=��Zי���z�:����Ȩ�������F~W��:Mx��ݩ�8\b�ԗE*7ڔ�z��wXW'i|iǱ�\����<Ł�ē�<�%z�� U�ә�s��|��7ʛ����^�&%ծ�ѵƅ+Wi�_ѫhո>*[��p�bpu��j��	��n��]�K�t]��j©�_WTѼ��ְ�JZ�}>ֶ�.Ƥ�m�AS�p���y�(��f�V��IZѱ�/���ܳ�p��ȵ�Ӹq|p�6O�9�����ʹ1U��˺��F�4��p�nG�2j��ټ�ؗ�S�1���,��^]��RmVPrZL��-]Y474�*��=t��RjO��1	(�5}*�J�ݐ�f����up+�*\z����a6��b�K[�*y..�����*�޴��K��T!�]��g��M� �{|����ھ
f�kU��Z��{(]ηkN1�Gu�!�mK����MK�}�+��m�Xr_g)s,��1yk%9����vٚ]�efu�.��.�Ϥ��XVPk�[��1�{6E�}h�����Ke���`��rЍ�#+$�wƆsl���ƥW���(��]���|���ٖ�r[M��WR9Ф����ۏc��ԇ������Y(�3�o
��O����,�G^,��vG���y�SWUq;d�<ƻ��`)�i��=���u���êl�q2��T�۔��y���R��8�ӏPb}kb�����)��m�p�[�o@:��ħp�P�{\�pG�V<���R�綜4n��ɥ�I�ݚ �*�&�<��=q�/�-�NK�$��v���fS�u�:�4
̷��\��vF�����u.��S���L1��cx��o����㏎��%4�|cUhű����DIvEZs�mj��Lԅ3ETS���ZR��jتtSU5E�4kF��TmmU�&$��d��-gA��""ccIZ4DA�1M�:���(��э�����[%SSh��
�TU�i���Um���(4��*��J�`��uJu��)�ld�Ec����h�*�))*��h���Bh&#��Mm�TPVت٬D�EX�j)
`���"" (����3AMG)�l�
(�f&�
ihm�QT�M����"$����&���kjb"��)�����U��;�STQ�
�)*�&��*j��gHv�me�ET�T�S�j�4������������E�S����󏄯���eA�U�/��'ky�g	P�lvr��(�R�}��L����$TxpДz�b���E���evlV)����"" >��� "s�{��YB$s��y���lOʕר]v��`�9a���ĥ2˟����d��3��v����wz=�q�t^LĝF�����&/�^�{�+1���9a���Qsy,Mm㿤��</Y3ԩ��&����:�q<oi݃K�Kg��Gx&{r0/�d(�u��<��^�D�����(�zQt�����6�O�<-���ƞ�+��K�U>COO:5ǰ���(��択�MKݦ��=��lE�9�]��ʵ�ʽВ1�!����xvW��wn�e�[G,R�DF������%��J��8�0S�i�0���G|�;čз�Jr��Z��0��Z�!H>�ʥKLЕ'L���c�εڠ�٥��k�3�{�G'����wS*�t��,��vI��j ��ِ�AhO�G=�>��}�5��6�0q�v3���v��zjZ`��o�C�ByI��ٓ	��pGW��vq�$B��
��<�c�9�g*��#wr�U5�k�����܆<w��|���0W��ڠ�
"Gt�;% NYb<`�y3(_�}��P['��K�G>M�c���:�������9�n����H���`9r�f ���R���������;(@�SN���ei��uC[�jh�srwI�x�����`
��31�<��>o_<��L��+	l{Fb�i)�K0f<}��s�����=�3{���Qj�AK|)3V��� �f�\�D�	E'�e��P��T:��4E��SȤ�	��W��5�,d�4xfeT5�i�+R�X�"���ԅ<�Ik/W�.J���t`7��:=	�򪸛a�kS��zKQ@y���'�_ϲ��f	;����D�~�^�C�U%�T,�!ɑt#$S,�*AL�3nA�xX�/��[�,�ٮ�;ʱ1�4�9�u��zy׷ܕ���uJ�
�q@H�U�r���르��ǎ�k�Q8�9��m�9���U��u�)9�b�M���{eO���y��1�qIY������,q�V#�/�0Z�����J��U����ek����U�YX�X����v=�^g�׾��ǹ���)�ts⺇V��������N��;����EE��O�������P)�`�;�7=7�v�d���y�[�T{	L��7{Ƒ���Z��E�O�]:5��Gl4	F���C���1I |F�R��Wҥ�7R'=ќ�Kh;����)��cFs���D���hL�x�O��3��X#� �gޚ;����S�2��gy��'Lni9Y�T�s7����h���֚��6^�Ýz&ʝ���s4�2��]��llU�F3��WHF28����h�1f�<4�'�l�.�N��}.��PR�����9N�{��� <>`=��u����Ͻ�������4���¥/.�?x�MW�~��*N�;dr9�0I��=�e��ɭ����[�׸����k���{g�m~���_��3�塇a���z����ܓ�u5��r�S��J2-��F��	U\��5^D0' �䌅�|qߛ04�67w�M�/�Rw���6�_���ˮ��)�O��>���Fq�7�^_w
-�՗{t�;�BC�]C*���ퟠwzq-��t�%cц���Y�DQ��_1��y�8�y�-z�5��sTU/-�_e������Yu�e�nl�XN��琎f�Ķ�#�0�X��s�s�������*�Z	�Q��5q
7r�n��7���R�$�D���OW����]����|Э���!��.bW���dd[�ɁyPS��S��������f)3�ee#n�?z��k5��Z�8D��b}�"�+7�A�ߟ�����'�,�]6��K���wB��md��ll.���y/�0��9�B�k��"�b˚�g�v�9|����������z��ӳK�gvq��q�%���m�d]�w��S#�2��tv^�JdFd�/������5סq����+��q�t�v�z���AWl�Lc��%��(C�]h����+�ұLɲ��wd,j'] ��j�UZ��3/����x ����ʫ���Qi�7������4V��Mq�h��3(��J|��������<�JΝ�+/ɖy(�����$k2D�9X�Su}�<���P��fQu�<S~�%!��3JyQ����[3�i�7/��+Ȇ2c�B� ,1�D�R|r�R�߼d)�S"��LS�C/R�qS4�{:���ren!�q��lm���舖z��f���,�fEq�~�=p$���	��zPY�i0���K<�y�↳�k����!��h�QGW��)7��sy�t�ݘ_�z��*�ߧ����N"����W��a��<�}�d�U�A�J������(I�Zd��גb=��x��sN^X�z�z�'U�A{����d�65	��Y����%����B;N����ZCs��d)�x��o��i�zxϣ�X��3͏fy�dԖS<�9k�fe�춫5�}��܁;�t1�5�岋ZE�X{F9�==�m���+՞xV�]?\�nR+�H�=�Ɨ�	��,��\{a�ȈQ��Md�����3!C��]�d��e}1��d�/���1Ӻ�y�e�PM������a�t�������pZ�W[Y�� �����|�1=W��L��+�ie�����ϝYb�r�q���i��Q_p�=x��.�P�,T��Lَ������0�����g��C��p������;_y�%���sF��SJ��XL>���B�&�#i�k!S��DoI���Wm�YC��1\�����\�`�0��bNH+�Y��P_y-�wsC�zL����������}2p�	�,��A�/_ ����!����cV�s��Q���4��4t��fD��0�ͫ�k
q��d���4�lU��%�b��S���f��m�*�Q����� +��]�H��|�ZX�\U;n��T��AU0y�U6h��s����z�����_��G�`a[����ux�t�"睺SpzV�rz�46�D�B��j6���[�%��&i��>�����T�V/|��R�t�A��V��ս�z��u=%�{��A��u� �)�6G�9z��C�V��h+�$�Ӌ<c�l����d�aڭ\�I�e#3�ݽ������r]s(����a�I��׮1�^�|9�������Hl�?�!��;��׍���K#\���v9n�*@v�b����/�h%]7�C��!�j�>�v2ä�V=�(������r���n2�2��ԫ�+$p �mÈsǇ����b�����oV!�_�oB��aDN���MSڶr9{�����4V�/�AB�Jxv���.#,���CND�EL}���7��� fyoyFcC2�qa�}�Cȇ�I{��t�/-�>�ޫkܕ�<岈Y^�z�]q*�L����h���,�K\�ux��35���y��	G�yV*ivt�s�-��e){�^�y3tUem9�^�g^=�#(I����KC���L�Q����!nz��q�!�򛡵�jBY�v��(����F2Oo��K��,o��U��("F�#�Q8�A|�[�]�o`|))�xBw_�;_q�����C���P��sx@�����^�t���#Y�m�	���(��j=��7\��F�����knd{�FfUCP��R1M�k�rH�#�ب*�Mc���|o���:�1M��M%2�	�!z.8�	��]�S��}��<Y��)�^��M6gS�6�t'2���oc*�`�3V��=�q=qp��kl���(��R
|��o�aV�s�ɤB�p�c)���d��s'��i��!A�hq0�ܟ[�����k�����U���۰I��YFd�O��u׽�)9�b�M�T�=��;*�l"�L}I*8<�#��_0��};�@��C�ܐ�yp���U>��<md��сB����̫i�W�ZR�-���gΟ��h9�;���PS�<j�FJ�V�����C>�J�F+o:�ޓ�rTx������ֶ6���mB�3˹��oh���wE��DM��1��%p���yE'���������a�3 7�����;�	R�������K�0���%�����&�kh&���?���V�޿�4���))����Ӯ�O�q�Zt;%^��FGsu�|��!DR}�J�砱m�r-�e��a'v�넮;.�������Klf��Q�<`R��oG ��Rhz��0�ܺ
�<�!��Y�*�K���ɷ\�u�SLI�q��dz�Gr�w��ʱ��=~�J��e�2��AמΑsJZ��ٍ^?Tk�T}���N��ӶIm���sO����΋�=s�q�]����G2�E�֕|*�akL���kg�t9�q��������}N|�'��4�8��:j��ƕڷm�v�mײl�V����b4:(J�研XgNX��' ��-N�2�z;��1�ʦYB9:���⡬��ͱ��w�<�*�qF(L�s˾�s�Qe������8���#=����Y�����|���V%��Y䧽$�2��<������4O^Nzq�^���JW�u�H�.t�1g���}�/2jM}���N����n`�WW"o^U[��^����.��jKl]7�+д��[K�E�ya�)�ޕkG���+�0-"
NW�2�~�I��i kv]	����+�d��%�*	H�5IlpP��%3q^.VJ3
��j����UW���Brm��3��f�e�� <>=��}��Kwp+fީ��f���<ڢ}:�ّu��)�SX���Wr�[So����;Y�τ��|���LxA�NBS�nP�y/���U~��C��uپ�|h�v���i.\_�tEo�1^�И���yB�߫H���G:">��,C�:���炵c<��������*`tcR+6�X��z|�S]cP���u�yPD��G]jDy�ڨM��}��'��[���g�����س]j�b�&�_�̢��J|�����?eۭ��{y�n\E�63�\�z�>쉊R��%�e�2A��c;��ʱ����]�;ӉL#Ft��kOE-��/jt����Ȓ��OO��Ys��3�<�S��pXr��>r3<����i����H�s�b���!�x�n���U�B�����g�{�~�<�<]�ȺS�DU,��\����9�B�s�h~������N86�GOE-�(����x����c���5��f?*�(��'_��)q��]<э��Yq�P�~z=̍����Nd��b�{.֞��8�J���$߹]}�1�s��7~̮(��lzG�y[Wya�(;�/3����类˹5r�B��I�n�jm�Ӥ�L�u��{��0Ŝrn��A��B�w;��@�V7;2�k�#�:N��T�H��3��B` ���������=
s�I�) ��7��0�C��/��<&z�z�	:�n���j9��MSkW�����A�Cw��V���ut��P(^r'L.�_W�i�ʹ�;X���5���fW�]z� �$N}6��Lw�Kz�����B)��)G��L�g��_�=�v)��pq�L[�FEN���KޓZ�K:=٤�E�5,��ϫ�}�sӆe�����W�꣋�o��o8ٌ�q�H�]�Z�^Ø!��	$su��)���'C�h��0G��s���G|��R���u�>��n,=��-�rz�P�m{��9K�!���h���S��OJ2}�d��W_fx���#mT�Ƨ�S4�^��Tv~W��,��4�7�+��"�TBV=uڮ@��s�ݮ֒�ңf~]�6h��yY5�ǡM�_P�4�oc{p4�p���c䭲.r{+_@��"��쨇�o���	��c>���]z���ע��+ܗ̲�qf���q�Q�.��R-\��St��u�+�8���KH��T#}��U�"�����J���	� a2���0�vk,Yo�:x��I ��C���r�G;����;�F�˫_,�J�7��{m��uїֻ_�*��(m��d�9�Ļ��M7�О➞��¸� uhŵ1�w�j�:t1Pйtq?6��?d���5���V��?{���{�� > � $ O��  �g3��>�#���_�}��1:�j�6����lfW�X���?��24GԾ��F����԰Ni�5(;!}��=wI.)�*���S�-}l>*V�4'CV��吖{�.z���[�T����¡�'���{;	�^i��]�� �G<�Gs֭��sYr��HP�'��=��w}1$w���9Q�$DC;�YTv��>4k����7Vy� �c39쪎��T�����Y����c�4�<��kސ�j��>\hJ��Dn�Y�;��]���g�v'C�mAW��qɍ����5E�xܢ��<s� i������BQ�U�����n7#ҭb3�䛱���wb��V^W��,�<,��&kӦ���W�;k� ꀜx�����/#'�+�0��1��Ɗ�%��h�����^��I�YG�x��4�)�jDgJ(_���m��z��e�����a�𬟥�����͇mU�A����n��l�8�'�6�U�Mq���hR�_�C�Cȭ�y��z����S����W���w�;E����,��B�y��{=>�W����������������18v7���u���ow��ճ6B�u$&5zT|�AwYj�T�Q��#�9��)r��ֵ�jd'Y$[2����+�3�V\*�%�� _L�g���8R
�k��a�Ix�%�3�����E���'XR0g)/��/�N��S"ڄ1�����qM�3:�a�2kTiNm��t'T�����o�j[�986��*����7BE�$��3/�m�ҩAt��X���R��P�{��	�+{��&Vc��>�L�e��;-�il�(q=��4��B�=-�ܔ7YAs�c�ܭ[%��,��#܉+���9�V�� VԷ\zm�o��Q��uO��o�m*��Sϖ����CJ��ķph�۟�ex���Y:�P�>��ރ:.����^(�R#3`k�6����.�M���� L��ωV�'o:�@�:0v��2��%�p���n=O�c3K���%O;���=�����z䬺m畱ӧC���33�*�o�� �2��EX�����>=]c��.S�:6wE{AR�e���T��"�s�G%%BN_WR=����t�d�]Jʕ��X �o�l&��S-T�ol첯kV�u�{��?�������* �7�ۀ�Vp�Q�1V+�1P�6�ˮ�2b�Sw�^����e](����2�u2+mS�����V���P�X�Yo���Wy`Y�I��WU���v^u7�4��MŔ�L��_Q$[z3486�� ��H� �Ļ#��%��u;S�� S�V)�_�L��^�
����X��D��oϸ��)I�ޡ[u���]-��2�o	*K*þ�����QA�\�Hk���C��r��C"��5��� D���y�����9:�,ܻ�*j�C��4TEܢ��64�������@;�ipk3�<خ��c�j��S�w,Ε�P�"жP�3>��5�;3�L-Wf�"�wYU�Y������t�&M��&T0����XL2��R�AK�6���׌!�&ͬ]�iAiԗ�	��>"aŋm���ح:;%M�oS �� EMD�b��:�e>Z6�Ucx*�B*�(j����0��rKк���5�c��Og�A2���l%t3S���b��[βlzT8b����5(]e\\�FcZL�!|\��g�$H�
Ӧ�u�y5�|�����i'W�m�i��D3��9uD���s��+����zb�{��AR�Z] p�a�0�¥?Ht��MF!���Q�k��9���b��#�]��Y�4wf��r�m"�5�sZ#�*-�����vbè�ܨҗ�n	x�t*I�b<���\�f��usw6�>%�T��x�ƕ!.��̧QfU���ێ��of���b5��
Cid��P�.����`w�hw1�|����i���s0�F��9ѝ�� �H?A��h�����d4�&�(M:���F�b*���Q���+�b ����������b��*���j�b�"Jt�&hִ����1%���"��kc�D�A6�E.�L�[�KDUEUPSӬX�Ѩ�QPDh�6�*$��T�1PAUKE44TN�(���S��EN�h�&�F�	�T���44�QP�,E%=)����ڬDQTLQTR�b��R�*�X��M$CM#]�
:�MhƵ4h0UE�@Z��jآ���$����+b�Mi�E4D�
ClUU4hЄ�b��f� ��l4ĔUUQc��$�t�44i4j�cX���b4j�k~�C����=n,���۳e�6�M�s��U/��O3�*�h�D�_~�X���������A?d(P(R�D�Ȝ*g#���%���N� SO����&��m^��8�U��oC'��1�;�S�	�b��<k�����7�P)�+Ipd��)�=�qS��`�:���f���C�Y#n�Yxg��`����y^7�f�I߈��?%f�\�������1�8�+��Ư)߭Oe�z7^��'I�TRs~�"�k�y��0v�B.����RVdY�[�*�ƈ+
���DF�t�f4q�o�<�ۢ��B.xRK�J-?,��Բ���$��S�ty�& f�����7j�^{�G����8-u�NޤQ��:�$.*X'��m*�yb�M���>@�
%�y�*in{͐�Lޡ�����5��*�	^��j5�a��wGҟ��Q��M��2[��-&f+���OvZ��{�a��Ť#C�`x�bT�޺�:���v2��naqJR�*��i���^�G�ʔ���$�Ȉ�`'DÎ� )����.�_�j��vE�j�0[i�.c��NV�����[<�^�kg���s\h{aY_p'Wg�2���G����ڽ-�a~٧�����dig<(�Mz��J��=I�2�{0z���{Qeܘ�C��)7��Ծ�H4�fъ�-�}D�j�qӉ왓8u ��`�fN�}�du�>x���է�Hn�<��J}*K\}c&�V�gr�=����k xe��6?�W�U~���Qi5q���Dwu,bӌ�j�H[B}5���W�yx�@�<{{�N�A��^�6�_^���y�]\�X�^����9����cmށ3�2�͗�b��yܖ�0�{�s��;s�X9����+�2>y���'���=D��FrU��$�/m���|�aAw=Z��O^=/�cU)KYB5p#D��$���_���&����7��Ų����޻��ʱ�>O�L���#���']q"�7���X���3d�CHm�NU��-���=K�Y���EBW���PdT,^���"�DY���ӆ��$?kd:ْ����F���6��|��Cе�l%�+_����b���a�j����	 ��h���A�K�c�}�:��KcX�e�x����YB��*��gT9�N�wFvo�PǛ�{�{��?G��3�^�)�M�kQ�[#��1鄟l%>D�+�� M�'*�ܮ,\�������bRdtd��e0{�$xg�~�2��"��eL<gkw�Dj�y������nLxw����SZ��r�`��x�t�Kנb�cL����
%���+�ķ�s�g:�Ń�^[]�D	�^qB�CS0,P�V��l,�^#�R�U�cL�γ�
y�[ߠ&�]�L�{�Q�Y�ݮ��?a��8�w�Vq�$�wo0/i]d����eg�Ħd��>��0��{k?WO>��}.�a߮�?Ъ��G?�<6�F)�E��Z�eک��{=�?��N���R��.�;A�z�}8�R�j��0�J�z�=�7��5�������9�S�ӡ�ZEP��2�Z�a`$d�Y�3�H��Zx�Lx_%��7�����Lh�%��jsb�}�3�
�O;t�`ޕ���q܆XnY1��E_y�6�:A��O2��{�����BBg��asЙ�.lTS)��-��V7 /ԱP�U��꣧��:>��C�WIDn��4A�(T��)��2$M�ĖN�w����+_������fv��f�ccg�cTt�����u��B:�>T�=y��U��v��9+k�?��(�su��\�^���$�2ς�wI�\�G���\`Y%9Kl?4̇���a����
-µ��ݒ�������	� �Üц���1�j"N�9 십���ɬ���\Jn���9��ȼ���sj���ჵ�4
ۮ��<������Դ���"�S�T��fej�+�F��> ��ܡnK�����m䪳�\�9kE�'���������2R��Y�^�
�����$/�b9�i�7�"��ǭG%�xw>\�A�SB�؆JR�mL�y��ͧx]�͔yn�w)����\}���L6<��O5K��53LJ� ��M�zD&Ր9�AYB��.בSW��N5����D&*KL�f���������{� ��Y^-}Ҫاn|>�4�J�9�:{d],3Bb�-}���r~���2T�Q�6�nA�A�S�l���TC@v�m��Q%�@��T�:��v]��ֵ�HՈTȹ�J���N0���`U�'pN�r�/�b�*<�vy��#^c�Kn6����S	�:�V�׈�UJn�	U��:�9ɋl��.5�}-�gv�Z]b&*��߮nō�25#4{�!�5�L��Ң�<�)?5���k�^�0��y�׫D�$%��i�m�.NQ|�L;��B32_�*:��e"�ӷ�	�J�.�����=�0��fmצxLS���)��'T,Ch���oP�>���T��o)�6�k���_���m'���H����ŧ}1,p^�T���	ސ��@S��w�J�L���ĉ��Ã�ε�7�g�ֲ����9��kQg�g����۵��]����HL.�>�2��3�P����nk"�AL�v�5	d���$U�wm9M[tk�XkCܹ�6���3��cE@&��ҳJ�s!�Wc�Tm��g�z��~��=B��?.��O$�-�T��%����۳��E�t*j٘{�l���}�Ur��U]I�MǛO�`�`c�����_��>���/������?1�~��r$�zG���v�2C6�(,'���蓨pms��ٷ¨O׏�t?��{T��\��ְ���ʯ{�eJ^��?y)A
�H�^�7|
��_y]Ǣ��&�x��n;6)�bx�w0eq,H	M���>�Mg�jСvM#���0s<��VIF�^j��j����O�`�۸67ޒbCr�|��Eis�z�h�q���My��X��=C��3����KBj���J���&�����}�-Ff�ٔ��'Nv	��k�3s��5�zva��<a%p`OF`CߕGTq;�Ew�Lq��ǌGj�C�L�ry=�b�u�Ν�PY���>������r��'�p�e-��8�T��*]���/��%�p�)�fHœ�&��qI�>���qH��qv� 󜅧5"�/�u�/h�"�<�5�Q8v���ע-��r���<}�8�WΜ�c�/Sj��{]�	��kq��n�9�֞��Go.MV���!6c��Z�M�J(��n�l#zO�iP%� �ςh4dp724C�N���?�eZ��
���5sٱ�'��r�E[C5_G+$,tH��I�w~~]��٢�Fg����)��/�P�\�a>7��[ �,���f:�<��7n�k:����,�8����p�8��r��n-�dG�g�ScTq�U"�jR����������b1_m�A�"�.,���j�u����]W.���+Sg#D��Ou�p�����mv�������L��=_J���o�"yH�Ey*J�W��ʙ�م{�g
 �7S���s�-y�<^����jđ��#A��t�_%�VC?q�*��7t-�QiP��'���lsaz�������`�������K CWt��]E����Y��wI�|ha���\	�vr�ŧ�#C����BUV��P��p��ĿD��]8�Jc.�	sጫČ���ܣ�b?/8�P'e:�p�s��s,�Gg�}�8˽��R����<j�۾�~�?��+5����ex�%�������(��E}%A;;��/��X�p�Rc�}�
=["���	���11g���/�>�5'���s���-+o��}�%�#�Y��܄[4����@�6�ҫ��"�/ʮ����S3X��b&@�~�}��!-s,C�uP��r��`����>���s��{.b�\|SfE��ԍ�r!j��H��2k���M����ӕ�`��VBʗ]�H������j��])kԥ�^����ݐ��m�X䜄U�Q�!G��#1������S�Q=�7&�t�SH�-�/���zM̒��D�$��]�z��$���蝕��c�!~��������7��J�m��)���V��B�P���yB�߫H�_w1�-N��î�?A���ѷY]�=^GA�/��C��Fy�:�~��M�`�2籊)?Xŕ�{iV��°޲���:jwkP�n\#�Z��\La��B/�U�Z�t�-nfW>�S�I��9�j��͍����cɏ<�����VHA4�aR��%�e� ��|d3o(E�v�|��z��'H���F���s�>�W��m�����,��,�����jZ*��D:j��3D�O�j:zO�����RϚja��q��杠��	S������Wü�����Ou�����8�E'�g\��بˊ��U�-+4Y-x�ђ���Ȩ	'ê)�p<2��.̸��4o_�P.Z�3	:�Eό�	�J�.0��r�j;�e�%��B���{7�����p8#Z�����p�E�q�Ƀ4�����cK�ye����[�J�R�U�p��������|���v�__��cދ1��� ��(Q�@Tv���>����yyޚ�l��A��~!��܋�tq6��?��x�.��p-'w��(VcC�K9��%Ԟ�L�<����j%J�Y���r�
�H��Fe+\�޽�uֵ!��N���q��EB�t�;�2y9�FWVf{�<����*`�nɎ�e�w�����F� �/�����[�}R������o��ɚ����5��_��hǯI�,ޑ�> ��D��"'���(%�"��dav`OǘV�l6���ݨ����.A�]��R;�8����O�
O>蒵y/�g�F�.s�u3U{,�y�k�}&�}6�"���F�ݎir��{���A�|�_��:~��c_���!ˮs1g��ެ�X!��+�Qk"�>7ln�46r�|T ː��˫!��+� �0��wb9C2��=q~F[D������ޥ�5O�f��j�mn�!4��m%�+�ǽ���u�B�ڜ�n���򤰓f��;ut:͚��z��8-k�i�ܜ�9)���^3����.1����������C�e���*!�Zĵ��b��ّ�F�9.�����;�����T��n��%����c�
�d\橶��̬`S����ad[��{�˶7��c���Hv��*���ж^�(��P���Oe�9aET��Ji��I��;G���J�w� ��h��;�y#�_dKG��u�<b����/�K�j����ig�0<���Kr�׿[�v�3ަ�_���ռ�s�M�q�i]���N!�k/k��Dce��z�V�G��J���a�50�h�wz�W:���9���ړ�n ]��4w�����5r��ۖ�쩊$l�u�$�U�Ǣ���JN/���O7�]V=k�_��k��,��T7��W�P�	ej{���u#��J�q����Y��[�ϸv���rHj(��=BTq�M�b�[d^Ҳ��a*�v�q�a�
M�:�s<��]���t1��R�׶B+�l�r
K��N�hJ��Dn�Y���b����2���u�V���-`�g�W^v�j����v4a�sZ��t]_x�dq�$�عc�g=��WV����~f�NG��x��?u�=������ތ#�?v�3�^E+�^P�7��/q��Er7{�&`)	=c�>�R;|����s�c�C��㾻�+*]��p�F)�}��͵�Tc:��v<`Ÿg��� �?G��#���G�@�xH�<�d����Z�8u���v�I��R�?_JFhd��k�H��/2>㹙Uw��ܰv[ޭ�Xc��D�C�?H9���o���t����|4�Q����~�u
�\�ߓ�=>'������g:7y�Pߥ����d�����8��#��~X!f"فX���08����֗4"%E��.��ƽU�m�S�9ǋ �룇�K�:n�]��v��9�Z�|V22��n��X4Q(	�58���X�M��x�)����X=��J� �E�q�xT �EM6�P3NX����-&�y��]ص�SC�8@�s{�t�k&G��+�������̐{3{:d��Q~�㭽�=�g��(2-��r}r0�n��GGw:^B�"7�U;���M"�d��X�S�s��6�k�k�J�K0������t��頍(�.���ۘ�_�6--5/�N��� ���A#8�-�Ү��2�-�gٷj���!��z#p���7�%�Y˯3�0q���k)q={�pQ�n|h/@|�Ǖ7�k|	���9���y5'/P�u��rn����}^h�pj^=z\��m�H��(�s�2�OT��T��{!��]3O��"b�[($v�����XkS��hK�sЗ��AXݔ(�Dc�\E�*��"�����C��:�T�����pt��kE;��wv�<��K
���žk��<�"�8}&���N�5"c���lb�g/V�Gy�!D�wv>ﺅ��N]�Atäx�?Oسb�b�s�}�-R�b��='���lbӌK�[pzC�zMV���'���Ĵ��e�ɆA�I4�+<����4$'�Ց�=��s�3�C��e;�2Xf�!��>�O�����z|�|�>>>�VH��m��fS�Xt gB�57�	�L��*ʷ��<�̓��NW毆�uL�34˘�iX�-3]K�1���\t�;��rh�x��՞1�k�n�������㮎i�m�����Ʈ[*=��ōm�	�-!p�/���i�7�� �YW�Tvƶ�+���Z�	h�����c����.bp��5;I.34nK��|XJ�uĭN��������#z�����@�=�̙�y�[ܵ�*�tRja0�E���m)��F�[�����ѽ��ځ�qܠO&�[�
�"}��SM�W� |�ޭU�tԔ̉���0]�������n��F��a�Sx�]��0C��,L~fpO�={8�[��wF(���@ݜ�N��LCnS'����&v�u�u��V��nl:I\85һ�0`j|�xdv�-g
7���̢�N����|1�|�]^���yGV��oX�"��/ճ{2����܌m���F�}ٝY�n�2C+nl<7R���*ٳkf7p�f"[��2�YXrk�m��r<�:v�f�����\�tOr�d�xC��=�(��J�T����U�A����T�>�­�n�2+�;4��s@�m.2�ϝ�;*k�Ҽ��lrVk�������{�����L\R�N�-fPݑ�u�He�,�@*mHr9]�|E�V��1��hT��R�[���q�Y�\�'.��3���jĭKx���&M��D́���XT�}�c�V��"���3w�㼦�.�ح��h�lV�T�\h��Z�n�;ծF��F*�� e��J�*9j�SL:k�c�Z��o�!x#�vtw3&]�G��S���U(��K%N�,�wP^\�A�s�+]��^�ɛ�ef�wI��I��(�::D��T8!vsw`9d��Z�:7( 3���s;I}:����f�}��%���O�X�Ճ�u0�T�~wz;:�l<�e�إ�Ao��R��*�}˒�-�f=çt�scB���mol)H�5nK�w'�5e��d��x644NOhc��z%,�ec��_V t�@tYP��^�u�ݪ ���46ƪ�����ywe�(=�Ju�h1�U�S���\��i�tLi�V��v�l��� x)]b�%}b�2�)�
�5V��Nt�X8�TghrXj^(��ڻ/Q�yӗ���&T�*�ؕ�άnf��E�������bJ8֡n���m�F�V��=�Hx�W镏¬�Ya�&1�#�Yݎ���
�;4=4�CYH.Ƭ�]���'>������)nm^�ԉM�.���h�[�"���,Zu��eє�=d8�=�����4�;� �Y��u�8��ks1 M��l�O(Q��6�?7�*u�/���4̝Q��b>�>�M�f��
|�C�[��:����鷱%������Xz�v�jwdӁsiQ=( �v2Sܽf�${4�s圦�0R3U�s�  h��J�#�A~*�b P��x�}�E%R�l��TQIH[(t��h	��(֐�F65I��4:q	[m&������E1%DRS����5������*�����U��Չih("*h�[�cX����UL�֊6ͱ��V�5�h4mdvآ�����Z��%j,L�m��*

&��qIO�Iv֪"��h��Q��X���b�*d�Kb�f���,X*���>��jkaѢ"؊�(�����P�Ult�ъh6�%%U:�U4�6�M%;8��O��8�b�RQ�bJ:�Uv�c���Nؤ#i�����*�+��[U[��ICt�"���kDlj�&��@QTUI��D�SED!��Z1Q��S6�Z����4֍���D�ַ�7U�j
�*�����:(#F���yulh�&�!�����D|H��>���F@�%L���	�ڦE��xz���z�d��Ԥ�|d��a��[F�� �} �N-(\\�9�� �l���$P�L����R��W�x�'(����9��ŉ�U�R�P:�A��w�>u�Hc�M��?c&~�<Y��M+��;�c�R�w]��CI7%��"��<�駁:�垟�H�:D�Şk�:Țs�9��v���Y��C҅{��us
����<��>_p�b�~�t����v�#h���+ɬ��1����,���t��۹V5xB����r$�Ӑ���a�20y�O������9D������uY�5+ʁn��Kʛ#Zv��.p��
�NR5�)�+��:Oe	u{әS��p�������0b�H)��S�J���F�ͺ���Z���=�OخEgJa����
#=�=��b�s1y��4[z4�N5K��-�5�ڽb���4Y�Ǐ����lŵ���Ǆ�vK�2�6/^�fe�5����}��n0�|{��������@2��Eց����Y��
|[evw�~,�ݏ�Ǳ+9clI�̸ �+�7h�~��a�	
���_��f�=��qP�]B{Y��vg[#Й�^qR�<����g���s�|���@1�_��ߒw�S{]�
��Gt���޽6���L>��۫�����ٜ�(8,�Z:�';�A��>]Mi��2$��ڡ<���f��ss@YNG��JRз�l���ɚ�
R�F��c0�fm?� ��nj�պ�%Sdݹư�a���{�˿�+�63[�Y�V�|��j���n�Le�X�>��EWa�.(�\��H�d��F��M?j��Q^�ċ]�!�����Ȧ˳�n��5̃ds]	�/�L�Ne����6.�J�.6�.�/i��_y),5�w6��V�����c���y�ؐ��`��>�ȇ��E2�Ӵ[��%��ƕ� �$��i����Vll,h�&�����f��A�J�u@�!I�d t�g�4Y�}<�MUo���`��zV��x������?G��2=+�P^a�^<�:#�O�+�ױܜ�OF��o�+�B���<�,PxŖ}��i�WI��jY�W�%�\�G���'k�\��ʻ������e���εz�#��$i6	w�>�!��
�`�9?��S�3ϑ4o��.r��9���O�b�N�Ｊ8�֯���a���[�r��\��p��K�&rI�6=����pC鈅� (��e�XV�K�Ɣ�WVz�nd�/�%�y���G4��2�������ǁ?geD;�	��y@Esgʽ��S��+�Uc{�+m�70׺a��\#�6F`��B��^�%�.��ȂW��[�F���ԅ%�v4Dtm�T7�]�������K:�m5/�ߦ�j�kh
2d���)3�l̬X��之�v��)����t�yfG*_�׵R<�#i��U��c۷��+.��P��o�y�V��E���\���6�j��>Dݭ�*6fx����L֏R�1gjy�g��@�lN0�~cd̷�5͞ysdy���א��%�7�(�P��gZ�������:Zg��Mt�s���u~2�×)�����"��gI�7�0���\N����w;��B����z<�EwS�k� �P��38��{��ጩ��E'�.�m*?1�9���y��G�N΢"a���!6�Q��О��ꑓLhW*v�a1"4��ߝA/�)���-3l���i	�<��Ļs�6��t�ף+�?�/�����ϟ���������1�yؚ�7��za{�qoa���T��= ��
��B�\w�J�L����/��\a�l`��nz�
vz��k.*t�`�%�(,�;T�5Z�Z�oނO�L ������/2��S��U^�MOy��=�س#��"��qϼ������o�=�,�H( ����b�5�y'k��ݳs�^�+�񐒇��>�?eO_ԃ\�	�L���f�ʮJPB���V��4<��2,��n�XS�턝�����{{Rԫ�@q���#r�뵆J�*P�R�ѝC��(�2+��\�t�?���uҳė�3�����7������^a;(U�:����%Wlע�KHTO�Qm�׆�fT��7�:*ڂb���Z������L�X����O߯��v[�;��1��l����6L5�*��[�77�������z�j���(9%_��)�j1�XU�l����ov��}1�U	�9]/X��.�<��a�Idw�'C�#���?�a� �����~���l�{]��B�Y1���Vw�}�Z���uW�M}�h��!��P��s�]"�FH��WW�����J�QD��̸���4u�]M4�X�XG*�l�����7M_�?��>M{����}˞�|ĵ�
!S��@��T���+�'^�LRsϚ����T-��e�QS���@��^lD��ψW9���"����I�g��m��3����Jξ����B�GR��me[B�oޞ%�2;s���>�!Y�d����kf����g���R[��M�uJ̙�<�T��9\��-As�Ŵ:��t!�������e}�S>���C��e��h#�v�ڙ�C�,'�n�)d3nx����F.:5�/ep���V����=�.�#�w����*-��U�ѧ���_�����Zx�`��t����+�4�����t���~Y6��	hBu.s�R�|1Y�{�M�qg�s�pXʽxƆ6
�Z#v�s��ڛ6S���q�	X.�jyW�3$K]�fN�*p�{����޻O�ԗ�4� ��U4=|䒰l�>�Z���cr:��.1���S=�~�쿚�,o'؞G����8����u�m,n��58=��V�Ưb`R�y�w�Ja�ا��խ�=�Q<�²�������m��4�������܇5+��\k<�xr��8cm�<�i�|s���'��41�8{�I��j�}\[����z}��
��"�$�W�#!g��H�/Kk����R9�����۽^�F�T�$�LZ�|{Ռ53z��	��a-e�Bp��g�~�'�gmz8�tT�c;܃�R.����{���e��@�DQ��r���	�?,�B�G��aޛ��w�J�ǂ֧xx(�BC�X��WG��A��|���q��m�T#��'_t|u�1�ߠU��	r��`�=��T�.�t%�\M�����f��܎ʠ�0w�5��!)���(3��gE�]�wӘ�4�?Mכ��Y�g`^P�H̩�+�<F�.�5~�Ȟ?V�D��aoq��w�ϲ���P����;��b�~N%*�>Jr�OP��M�d�c�~���{6�E&M��_2�z����=t�?�/i�����Ϻ�2tX���������3�1A���%z43�v"���}��gi'ݏU;�� �r�A� fT�a�Z��لw���uj�w�ծZxYo)s;��:0�Be{�k�2N��a=��EX7f0;պ���PE�Gݿ��{M��T�L���6Z�b�&����"{�z�l	x�Z��{]��*���Fw<��X�!F~W>�9X��5ې<�ĕ��)N��6(���v��v1�)Er�n~�w챶'�y1Ǎ��F$Be��/p)y��C����6�yO7��A���jSr|1R����m7/P�8�R�6Ջ�yV��5�̨[��x�ەr�>�O)�ĊC�їr�sH�d��g�N(kg֢_]�Gy��$:�k�(�CI��Ŝ��qɓ)������b�yZ��zt�z�w,2�R�Ft훬��g(�F��^O�"qCE�/F�Z״TQr�u��`{��d�tRӥJ}�8���h9D��&9��	5M�C�[Az��p�d@�PzB�v����ӟQ�K�e�W�=[�ՙ�X��W�0��O�����>����@o�DiG�:M�����,�y�ʼ{�Za�v��y/VL������v����y�,�LfJ��^�):�1ھ8 C��k���˩��	�����dS��ڏ�3�)�ÑS�z�����i�y>���œJ�Zލ�����k/���{ϖ}okMi}�� ./�]B�_�
��d�ٗ��]�z��hVwk��Gf�&�*�y�)�ծ�w���/p�I������L4��#��C^���a(�8��s���m�ԑB=�R���vիDI�!���J�\f,=?n�@�����g�_P��S��X�����%lRF#��m�O�����$nT��Ȑo� ��GD��.���F���� �u��,��l�X�W_�z��u��Mw�@���B�T�	Y�!s�4>�'�Ӂ�1?�,�9W�2d5ब�F�/3��.y�{��X�4_^:���y�/�B߭bO���R)dw��
�ʹ��N�Z��v":�!@� �����3)�pT_����XE}��!:�K	 V����m���y|:��m)h�!g�xc�h����'�ߢK�30� ܶпN�F��٪������^_[5[�%����O����M�M|Z��H�c*Js�I��?6<Hg��\��GN�<x|�W�k�M����I|tJ|���٦8�����b����Zk'j&��i��5oܼ�<�1m�E˻�m����8��D���Hn�������=+�����/������P~M�CޡK8�۵Jy�{
ui�\�Fa�Re��q�<J-7P�����70����/jd9�Z�*g($��ʗ�*@/Z|�X�$U�O��\�*a)�Gt�N�8z�=�8R�ʟ7�k�Pio$W=�9���w��D�V�G��P���EnG)d;�Q^H�b�6�Z�5ӶY���>x��=Q����Κ��'�P��W���=�zl��n���������r�P�b5�qk�b]�sZ<��3��!['�)�:�-�£I��jbH���:�Uɔ�˙ߊU=�D�yL����ϽGè>u����;V�h6�	��^��`�q!sp(H��*ͅ��#�i��;w��#���Pf��4�O�ҳ��"ظ��a���#�b̥�2������.0��fù�b}�v�����s�9o�-,y�F�UB��Vd��>�lR��xJ�f�Y���w����Iuu�!�TN9���o!\��nS����mR���E�D�]����ܲ*�n�m�K��5�U��Hd�som=��ҟ�NzB�syK��>�NϙZ��gM�S�+&��'�Z�W�K����2����'�y��ӬB1d���z�ll�x�S����^~�g��2z����+�����+��Zӯ��'�{�"J�DgYjn��s�9#oa/(���#Zբv 1���V�r���F~�'Tk�.��٨��}'bAv�I
@mc��J�D�<�:K��X��Id��/�+��.|)}P�?�M�F�=�=�C̅Fډ��i��Q��7�omJgmu�O��}T�"
m��_i��L.�Q�0XEU٨,���7m��=����mum�N�U3�9Ms-�|Uw4�]cpȊxy�ѕ����f[O[G]�<�.iw`=��F�SC���̈u� ������G��ޯu��S1�xޣ�eˏ�-�߳�G�����{�ԧ��"ʒ����чftNU^F3�U�ͻ�i�0,�+��ă)̄wV_��zЦ��͸3|Ê���|��/���D��B7�!S=�����1�Y�t5OH:���7{���3(D!p*7�N�b÷��|�Z n%�a�s��_�a<��㕥�f���l5�uy��}����H/>�+G?@��͜3ڸ	 ���3Чj������q�Ȅ���z�_���W�x
����A�x��p��,O��J��,\�>Ȣ�.���3ы7���֑�P��ߔ����#�?	�eJ��+��g@���oZ��������j����` �`��?e'�6�����5����&�cy��LN�s��*��T���M[�2��2,���iB,�v0z;5�t�n�fl�Y}M=7�F�L�أ�-�[5�|�Gc4V��E���&'ۼ[�$��-*F>�I�:���ڵ���rٻк���>��ڻ���/#/���>�ҧ(<�c�%�0�S�9ob�s0,�U��7��%At�/*�MX��Q�5��3�j@w'+ĝ�f��{̣$^I�C������,T���ʸ	~���NT��:|�
�ݥ.�2�D�t�	�S�2��h�;���Qg��{,���H{��m�	�d8�ZA.�u'϶�jՊ�b�J߽�����z~I`��U[�9^D��5-n0����^a����6öA�;���������g�c|���[�	[!Y͡���5�\(fe�*�e�DV;ǟC�f"�Us�%\ɛo��M"�������D�u�ש����wy	{P��'Z�^ePm·=>�x��h�K�^9��\椻�n�7�q��&�6�4�֎��3�����!�D$k�z��JQ�k[���}~�_�������yx���|};k�*tX/�t�-9�����8�ڄnQ��((��C`?����b"=Z�U���,�g׻�����g![.�f��tp�XN�J��(�&d[�+����w���"��p�i@aƯ�s���$e�e:��kP�i������약[Rw*G��-_A[� W�����fT�R�FW�;ʒ���Ry�^�pK\S:ͷv�ΗBd���C���2Ό��NiD��0B6�l��5�5�,��)�Z)�71i��;�(����հwZ���<9hc��@�[6���iF;x�Ck�ɨ�Ph���b�R�q��<Us�wef�r�|@ٖ7U�L�j5�{c�萨F\��1[���[�鄇3|�oUpJ=�8b<nf�gm�.��>�y��4��p��I�یL��[��v��6�`���/����Mn'*]u�;��ԣ�����3���@�	V�cT$������E�و�%�TU�M��z�9��#Wٗ���F�ֶ�b��u�a��a	�S�e	Q��#���.n{��Z��2��Uԯ,�`�o;2��!>*ic�-����KfV�O��9IN�J��qb�): *� �U\m���fb����ǰ��)�e�Eչ׈�ۜ���gq�O7��}y\,.�Ǖg�\#�֮��o���Q�z�,�EP8�V�ދ���!UՊ�����M�u3rOs!z=��k Яn�a�kc�z�1�_u�b�SR�R�u<��������̬�Y�ê��Z!"��d<�Q�l�c�ʲC��*U�\l�8vgf��ݖ�����t\n%6��}�E��8�����TN����a$��}������(	-���F��FE�]� R�D���Mn�r�*mS�c�^�ݬ�C����j�4��dK�*Zs%M�Xa�Y���.�[�me�m��)�eP{��4:M�D���ڟ�o����$7(�w���T/���YY��
}e��o�Rv]b�Pc�� ;�����C]u�(�+$�0[d�H�u�3鲱n5NK��46���Nu��&TS�R.�@�ǅ��Ig�n��/�;�2�����ѱ�1��;{ˠ�i�<(dK��i��7r��y[�H}]7�v@�hP(nr7ҁ`��Py���m�Qg��L�n�����F���Q�1����tb{��������t|�yWY}(μ�C���Cr�QY�Qn�b�]F�	x�j4�0pv�N��5���ɾv�5�sgZ��]�;�b(��9���q�k�>���
*f}Ƕ۽��ac���e�oC���6�u�uN�ɴjIG���%n���Dnk��Np\�]�*�b�qn�+�5�u�Z��"�c=����[X�3.��wާ����T�V!�I��r��(���n�[��p�0�ΒP`��©�gT�ȡ��
m��m�G[%A7���w
ں�:���E��qs�j��k�c�&U�O;Y����	���:�����_o����q�M1Zp34�-Dlb�#ͪ���h֗�y:o6"��f��(�b��(���PSQAQTT���A,GZ������j�;����Z
hѡ�,b����"�DDA��j���FƠ��'lDv����QRD��.�]�Sm�^��k�5CDQmѪu��U�Dy��1\g[jj��ѧ0E��|��j�u����I��N��փ���zլASvq]&��3O5�َƂ{:kF�����]�b����l�Z��csvn��(f�k�6��Ǒ�kͺ4����3th�1ME�5E��
-��kl�%D5�]a�h���DEh4�l����&�+ll]f����������ZՆ�P15���1Tm����m�����Ѩ)��n�4��mF�Vۮ���D����a��{o�{l�ǂ� ��ջ.|b��P��R���c�I�i�f�3���SE2E�*�9����SA��wa�n����߽/V������6��~�*aM��&U���W�����mAI5��:������=9��	���ZCbR m�O5-i�J"s�\e4r��1]�9�-q�bv��n��:@m2k��p�\�S�.����m,&rC1�g;y���w�G����d2����]�fۆ֣������1�&�wĞ+����n�������P�i6��m���v-dl�Z�v���K�@k*c
�f�]�y�2�4��G��eg��a���1{"���ҹy�#v]t5����AUo�LwT�sf�E��ւ��9!��n𕻏�ǲ2~}jm��ț2�c��{�k��������F6um�;z��C_r�\PK,�Vu+���ҫ/pv�귴9b܃="�J3l�;��z�Z����η�*�"k�J�x�dwh�����:��\e�������4�w�jW��{�(�r�ć�$�����l֌�JU��yD-�s��H+o�Qqy�H��V��e��dƫ���>w����\|4��-N�9Z�j����+�K�ݐ�|R�e�l�f\L���r��u��Ѵ����c��{u7��R��_Sf�	Bш=q�>�]a��*VJ�}K�V}��Ѝ�昺��[qΥ���:�y����wg�X0�׋�Ÿz3[��J%vV�5��/�ǧ��yD�~qf e�7���rc=��e�q���Xp~��k��%o�K~��r���M��fv�a�}���[�&4C��:xM <;g^�d�3��G��D�Z�Wr�
:І�M���9�'�4�ڊѪ����z
��V]�2�\r�`�Ŷw���������jc'���l�wD�Oʷf�oskl˛��gL^ȹ��9��_�j9ϓ�+�ԕ�Q��5P��vss^1X��>�.-�h*H�uf������=ls�I�7s"zd�dB5�	n���>�O�6)�v徉VxV5�d~A�W� ��^`ut⓱[/]z����r�x�-!̲��ؙ���Of�fy�<�I6>¹U�|{$�6�n�k#	�6�q�0���[��Q3d�
�I˦b�.���$�WK���h���]!��J ,���#�Fǽ��Y�F^e��\�r��<�>,Uγ�J�I�S3%�
������tI��P)n�cT�pH�*����뎘��<�{�k{��i�y�K��;��y
���~�y�F�^�e#��K�CZ����_.C���eeqj}���hӣl�_H=5�'�$�%QV�u#��$��>{����N*�#���}f���4綔y�wX�K֤�%s��ݽ�����f6��U���q'F�Mt|א�Y��kM�-i����6�1Ɗ����zF��A�}�dH����yxƥ��T�0Sl��Zh?$Atnӈd��l�v���������KI���e;�)�D�["�^�;l�#����}�9-7;��c��V�X/+v��Vo\ʎ��υ�m�h�N!�,�ї���h����{�=�x�uܭ�rR9��[�y�x.��cqz��֊���o״���U#W����a���g�ʵIw���օ6N�6�*!�GLD�P�e渞g�����5t�D$jg��Mf�Le�nT�^�����vv[5g�ԫ��pM�Xc5��P	3h�Q��
$�q��k6~/�wC�ƶ���gX+@A%Ps}KMmW�r���W]Y�\�9[2��	�|����Á׌�[ntĒ��0_,���ҫ�O<nI�O+N��xgj�Ƿ,u�|�c`&sD�t�tY���8X�-�{������=a���'V-nذYwt����������wh1���0o4��d
͜:3�.��>A�|9V[\;��:ћ�;r����A�%�?O�6q�'�#o��#sk�U �u���m�=8ӄQQ�q̈́��<��r�nL�@5��Q.1qB��E�7���HD�T2[����X�X��2|4�J�n�S��Q�ݻ�.�M�v7oD�r�Avgѧ�&�W�ɝ���_s�xd�Stc��`g6vo*�Mʉ��6��ȋ�������S�WS��S�����W'2�E��d䞜�
z%����]�����5�X�����2�z�]	��`{$Q4������]��� �]VV��̙�n�U�M�L�6Gb��WYw����w6gj���3h�=���jqy]�W�^D��c�3]��~�.�O%0��X��"��u���S0T���w^f���"ezV>H`ƽ�np�m�6�*v�n��F�'Y��P)�p��О�ޛ�q�`�bUۡ��tDG�PEQ��3|����W-���
��ϝ^7.t��pva�ө�O�ĄdT�����u��Q�7j���[�4�IF��*�^{v�[ +9�əUڥ�j�]!��N��xzM�Ӳ�!�>�1\Y�o��	�U����wQ6�p��E�i���m׺����Ӥ�Ϸu6��M�A7KU�ILg�4�ʁ���n$�9�ܹK�RF�l�v���LAD=��j�J3��;0K\u�5�f���)� ��8����~�~�+�'e|����J��^�IOa�����w���om�(�ז��t܌�q��Í7�6%Pը�J��ZyګqU��>ܢj�>��tĒ�>�&|�!�t��q��K�9k�)|}���"*��\�fO�S�cql������'�jW��Fy�׭-:��U�[Dm�E��"���Dp�K�����J��:��i#��xv�w���M�@=�":洖�X�{U>��=�Q�%<Q���wr��L@���Rh�D;��|�6��o�,����D�ږ{�+���F���r�7��QL��;j\�|4�Jd���.@	_�>pl�g��W�u��N���:�	�ҴQ$�Đ�1��(�^�n���R�KcX��V: �ޛ�jz��Sy{�~U��3��a���.z,U͒�zfJ���9Rzy�^�/@rY%\���{BX;P�j�v��:6�mx�!S�y��I����M�?Wq�A��kR��T�����+d�]M��b�c�n���W@c�Wj���M��,�3%J���v���(�JF[2�����ֽ!�gKS��s�r�mK�� <�K�)��Mo��4�s�x~��+�L��~��۽��p�X�|�Z�}y�O7��{�+A�}Q�9z{&��7����%iJ�a2��{3�c�Ƕ�A�V�)e�8�� �ͻ����drU�g�'&�?1/{�^� wC�#��!�A��x�;F_v�\�=5$nt����ZZJ'=||��v�ֽ���^˸�쯻�5!�w�;�[���E�n�+7��֢)��;<Z�=����� �kP�̸���"'t,���L�;e9,fQT�t�x+,�hH	��ҹ���Ȅ�v�m����1`�r,ݴ�x��*ĕ1��7h�J-x^\nG���ܢ�(f�]�� ۷����6��Lh����һJ������9��Xx��#�qe�S��5�o���������O U�Y�j��r�k�UI�����g���g��Q��#NH�^�����{�ᅻv��τ�n���~y�=�zw]����'禶�?+÷�㪬��)	�B]� �<�������2��h�Wx�#Y���ܞm-��	~Aܻ �K���~Q���-�X2��P�E����b"8�u<����?�"/HTQ�h��P�fQ��2ᶝ�����C���n�g�ޓ���a3�/�NR�EH[n���ǺZ�T��Ď���i�ع;�_O���«����iY^�@���;^J�(%���9oW��;�E\�΍�ݥ�g6����o+7�.�T��B̝��ڱ���^���^sGH̭1<����2��z�:}����\�
h�'r���'|��%[���Hk$�ͮ�#x�U��7kyU�̖��̀'k��=�bö���1;sZ�,Z&�Ht��@DZI�ܱ�΃t{\�[�M�b�X���*�@�[��!�Ԉ���60Z�&8�¹�eKp�dd�G���-Y��57Pn�6�l]c�u��c`3/y�t��NWuE��v�>��n�gC ��ڃ�r�m"�r�D�ȚΨٮ��Y׈7$RhY��G�j�6�k��{!�/w�E.���c����;*oi�o��J�~/S��=d��a�gf�ڎm�*�KA6�q4a�����kJ��ě�h%]��t��%�g���cku{�얐�� J��~<V�Q�<���7c�YV��h��u�L�*�:ZqMB�/2�,���g/��6����F�J��3��k�=����2$�ę��Sk�.m�t�n��� �6�-~�����m�.���o%�h����FtQ��v`E��u�@��hA� ��2=�8�d�e����"紴4�uPֲ�Ҧ��RG��n �l
�e�z�ݨg::�>z�쌸���zv�\>W�ԥ���h`�y�5���Ah�'�$%b�Lr1"�T.n��G2�E����j,y��O�U�jrɉD���M���vꇈ��O�7Z6+&|�wEbl������Q��i�Ux�e�Hv5Z�&a���n�_��mm/є٠�5F�ʹ�:���5����xܩ�5���8����ثohK=<N�����ۈZ�n@�М������M�E�r/+��'o,X��v�O&�#�5���~�?~ܣƤ�*��%{�!;�QR�v�k���<� ^os����������wP��S^E]Gc��P`D[`�O;��s�z��[+�Z̟%wU�6�>�e��p6�H��CZ�J���h���R�M��z$�����֎(�x�U�_�S�ձ�f���½}�������3���Hk�i1������$d1�ul��X�ʂo'v�5e��"���n3ޠr�?�'���+&/�W��Lz9�2V�_+n���vc!`#CƼ�sǢ�c㳲
p�O�5�b�
�k~�&;�V�	���kfӴ2�|��ҳ;bwK�R0���pfp3X-4!��]^������&K�������~��V�i\üĜ�h��6�#6線YoH��,��y�T�x�m��>��WjE点xތ�o+�@�04p,}i����]:k0�:M��{��4�	׾WS�f�b)��� :k��q#$�M�M�ֵ��V�G~�6�35�ȕ��\������ehBl�%YU&-I}0e%;�@N�������a�]\6����+�D����Y�̭�u��ͳ[Q��`X5Y��:4Vh��.������ã���M�;m$��A������S��ou^�4�L8�ZO��j���3 ڑbɞ���=�s�}ǬO%������M�i���Vp<3X8u�:���A��*E���{���Lw�e���O<���9�ε�����>oLϥ�`����6n�󋻗S.®lV�Y8Md�>j5xb��[NѦ�H�l2��L
�Gu{n1+�G�T�t%�ba홑]���Q���ّj���������.�oƽM���mM�6.0�P&g �-I��9,W{M�C�Z�[�36r�zF����3�:�nMĬ4�q�(�+�EǸ�,��h�=T����#j��+[�[�m5�"�;��}#�p��z����y����/L�މ1X+70�w[�����?�+U�3X�H�O����z}�^�w�����������ċfz�z���&�{[s���(�o0୸���]��wD���� g%
֘
��c�o�Q���ss�Υ*���U�;����ְ�0{��Ȳ'.�y�\�9<�PJ y=�6iT'4�剮����+$�yt�^Ğ��o�\���</�
�iLF%�_.��ұt�\c%�vep��&��(��?D��$�������Mn��m+�T��0mb�Ȯ䮇S������,�a��ٲm#.N����M]�"�*T]����xD7���#V�kJ������8�)�hcM]3��O	Xs��Ţ�n4!Ҍ=f�k��J�@�-d�J��9��.y��HP#ܝ�:�u1��57�UpQm����d2]wU��7'n���x�ڔ�̲���{�{��k�P�����w,����p���9�5ΰ�ɷ9�Z8��Y����ծ��O1/��xº�B�چe���7�,��m�M#�wqzm=ډ�h��q��O`hA��t�X��Mwf<�ǻR�E�{�EKC|���:&'9X[YI��nīۆ��ť �4����;��]K!Ւ�ֳE�=g�0^qb<���ǜB�F��T&M���Xĵ}6��3L��*JF�m R|�w+�0^w�%a�A곒�u�w��J���6ƴ�dr����e�@�Lf��:q�����q�s�ԡ\��ԫ�Ue<*�k���0�z0��"Ϋ:]�'��/�3K<�,5��w1�Bɸgf�'	��a�4���j�&�R�I��$����:��w��4Vݖ�Q�zWj���\YR���Q�2�V��J���J��u[
opa{�E���Y$<~��9�rp��ʚ�r�0�+��RR�N�;��D�k~)Zם�� V�c�߭�� �el��w
	_Q�S�L����</�{�՗�Bes�Ѵzn'�+��������u��=l�����x���7q�2�Φ^c\U�m�Z�n\u*�x��Ȧ��w30��c�rtAU�8�}�[|�����9�>�h���6���e�w�˩V����M�u{�����:�єe�B�E@���J�����y���t�2�{�*�|v�etɦ9�q
��Pڻ��l��T���Y�i��vP���-�eS�.�yne��f���* ��%����75�u�3:Em�8(���Z���eV�=�۵�j_��A��ӡ�fgM���N*z���ul���YV�m 
���\2�0�*];�Us�z���@����u����Kj���yI���v�(/��:q�R�^>��l���$o.�}���m̩�t�o���t��	X�<�o_�]�֖�P�ʱL���wH��[HûP�
yz�(��^b�&�Wc7�T-<kH�Z��ՎCw4#�iVT�|��)��v�jTA�&[�P�[�;�J��F��WVUGz�N��_��H"����8K�݂��)���5h�C�@tn�Qu��I�q�֪�,`:�:::�X�EgZ�<Twv�Zwu��xIC4]SF�1����X��
��EU�@P�l��F�"��*��lQlj"��4Ɩ�uG]ۭ[6�ДtݺӢ*(5Ѯ�����]t�Q�ln��q��WN�PݻT�g��E���wS���DATmn�m��cPn�6%�I�n�#D����u�k`����혣m�+Eti�mb��n1����������v�Z���4b"&�1�j`�i��Ѡ�$��Ѯ��Nѓ����n�I��kU���Eѧ��v;f�ja)�N.��wcv��yƨ�<�q�Wv;mQ&��5�IIѣ�CC�v���CIIӫ���u�GE:&����EDn�:v�th�űvM�]nݱvwm;�bzzttqA�DN�F�n��Pc�ܘ�� ���ӻ&��&�[tu���s۬tAւ���AuG�Q=����D��n����U�Фo7��im����tv��m ��K�f��s�-\�'��Y/��DC����2Vf���ۥNPD��7d�J穇z�v|Y��gN��K:�2�[,��G�G�K���M���y:�~KLò��B|&���W�Y���a���̦��q����y��y��LJ�P������d(���6l��20[����6�\�k�>ha��3��޻�A�^��Oc��~�g�C[��cV��u��F�g̩�̒��2.T�;���x�u��1k"笎�`̹��X�3{x��6w�;��b2 ,3y�ql}㼘�K&-M_ׁ15���;t�B��n�3ճ�!ԍ�ΗC�����X2
�7�v�B�5f����@��e�~n������r����D7�mb9�p�r|x�|��{$��ha;��uW�m���,�=�+��h�*u<1@X�bq�!�;nK��cRsV��"&ꑳ��t��r�54��u<��|v+�F4��T�p�z�M�:�(�Ҹ#��\�]1�|�n����(�ە�a�]+��k��#��#
�G0��LX�.8Wo]��w$��5j٤C݇k� �8Ze�ʾ����[(u�o!R�=��T�4z�VXv�Z��I[�X���om����ho1�Εq5�\�jX0rC%pVLĵ5ْC�{f�������ݔ����� =e󛷽�!矼�fO;3���i�==����f]��"F�:�ͦZ�BBpyŝO����Y��E�PS�ļ�l�}�$�4j�j����r��������sϾ�H���\�\���m�u�EW��ꮼ�θU�o-$��r�<��3�NA�g}+�:�4�g�aq���s��#p��J��z��o]�^�b��|����Z���n�*�vn�K�y�^s�-ƶ�������gۤ�h��4c�]�3:��q��y���s���"X�46�rs0!�~+���z�#��6g���T��+�WZ���r~z��˞ŭo
�j40��ؾ�7������6ɦ�����:8�e�w��Ƕ&�ǯE�[k��ps��[�!�I��mz{s�ݤ���D������f�o�t*�c���;sp�;�N�TtFB����%��P^U��<�F�\�D �l�Lw��־ R�E�r]��Z��0徜��.1ǖuCB���8�\�շ��sk��EA'<�C��Q�|�;��Z��%�Vi�iwi�lϋ�~�Xd�ک�*�X��BNMS"����
���wn�s���`�R��)m3�߷(~nh�����^����W��eLM�P��e�n�n����
�jY��1y��Tĝ��OտRn�k0���]t.��z"�Y D�����3m��Ӹ�;M��k�f ��Gu?;Z�9UK٩�bvE��o�G=��7�z!TPQxiUX��?d�\�n:�v��vT����;�e|�;RR�vV��n�z�ڬ������*�fJWwv۩��.�5�m,�TΑLn�fLܽ�����;���)л,��«x]�)ؚh0kO11��s�s)[ӹm�=�!���M@rF|��R�l�U�ٸn�og-ķ�B��:j2��������E��qf��J�M"�QK��������3<�hv�S����u�}�$x[�뵋��Ngͤ��u�a=ٮ�5����w�2�Z�I��u���;L9��k�<Zޘ9[{uԭ@8p ՘�h4�\����:���:�7yQ��A-^���{�^�"�`��	�O�[�槞��ӗ�Q����p�S�ؽ���ɾ�|�'�8���P0A{ɵ����=�0YTn�K��dFG:�M[���Q�Z�|S{ue�c�����`h8+󏆪�[��|�_�d�L���W�PK����L{zrw�����y�����B�֩��S�����>7�@��f������M�Ưj�2vm�K�f�苾�ۺ`Jg�c��逬�5��`|�=���N�r���+F; leG��:no���|9���y�C�.�����5���w���<��\v3\�G`� v���i��N���\������8jߧ���[cT�p�e��yf���������?���\\4�S��/H\A�.�v]�"�c��5ҍ�5�gUZ
�qGh%s����E��s"��ǹ��L:}B���o$�3:"�
��=�|u�h&�kt���b�t���\�e�:����C[�Cw%�6�q�����7i˩�Rl��#\.�ŕ\���tX��ڨ>�������*�u�י�R��P�����A0q��;�γ
Чwf�t%��G�(ѻ���[��i�N�#�D���(��Ps����X�b�x��Q+zKa����[��.��SM����X@�'�x
J(��u��.�.���5B�r��<���~����?^!�,����`W# 6������]k�]46C�RRA�3g��a�ڛ�ub�z�{6I���V�p�4?�+T^�4�*!Q�]{gg{S���-��E��K��Y�T"�[�Y�ϖ��h"d�ǭ�59m�KT�;��{8�ω\�m��r	y��wc��ȩ�BF��ѻ��6-L��5���G,�1�[Ӷ�6��4
�X�
b��sZ��=���6�aՉ�{�����F �c���S3���T;��m��^�l�w�8zˡ'�����V�N�����I�E��\�Ç���/�_�m�$KYظ�^v`��vLd�t���M��6y�<˪cP`,3v`^�>�=,o�D�?��g�[�a7��Tv��uS��m���8.��`�K�E�yES�E��a���U��`�7}�=y>�GQ�y����n4�uŔeù���Ei�����V���@��sT�SG���w��0sbJ
X5P�ïK�u��wװs��1�u���V�[O��6+�nxh�ޑ�ܳ��y�P��t�Is�qʌə�������k�q�g[��yG���(��y���Fi
��n�r�F���.y��3Bc3u��2�����s"�Y6�m�	��*:@[o����Ѭ`>�8e��#�v�}�o�Gsf}.S�%jUZ|�s�jN����5���2}X6�'=o��QxFvL�{N�#S�ِ��h�'�"���B����<D��w���蝼�4QIP)~������$��P�/d/��nc��p嵯�����m9�;T����1�r�G��f�A�[\��;�-�S]�M�(�f����4�[�/x���"����	d*��Ԣ{�*Mr��'Ṑ�k�;s�\�#��(�ͷ˽�n���tF�������s�O���s+UY�hYV}&)%A���T�2ȋ�c6L����fj��1��^XE�Q�VuK<��]ǘe�4�=���gL۫}g�V��gx�K�1�K9�W�L��Q�y8S�ᷮ���o$ڀ.�+E`i���:�\�PeАY��nw%���S���Q��n.�3z+v�sdC�O�q��ԧ�;4��GR��oM�mb����:�Ζ�Y����2�3�!�6`�H�(�X��7|��%rR�w�_3��ӿl����ߧ�y�\f�?N�h1F`�5���pD���Q�bng���5l���ά�8�ʳ����d�m���0o4�+陨[rD�?Z�9����x�C��k4Էv�����Nם����u	���e�\����*��EnȀ�b�+�:���.3�č~��Γ��}�Na���}:j���Cڸ��^��*���t��!��PvTcVUt-=ZY��յp5�W�r�� {M���~�~-�I������<(v(��:{���7·�\i�Su�8�i��͹�T�{�": 	���;���������漾�����8ME_���ߡ����"�CTy�P9Dĳgn��R���6�[{�>7hh��A�Bm?e�����5�I�8;�R�[&lą�쥧��R&i[���Df�s2��7*�6�n�Á
f��L�/h�:E��h���^��aNA]r��Q�|pt�t��m�I�˜��%Z�s��UN�N�o��=al��-fHJ�ӭ�e��9�4��ݨ4�aSF�u�ԑH�����wB�JD�*�uW�Up�N`w~&�\K��ǻ��gXF��V����d�:m���-#JF�F��{t�Z�k��q$�e�U���wL螩��K�N��]�mY���4�x�T�wi�j��3ǚ.����M,���6�3s2̍[��Ɇ[�l��]U�|��.��JVq��>�G7��s����¨F��ڋ욫�/��T��	]>���8�ڰ��B�g�g@|��O��v�k�h":MeɈ�1ʇrն�{�m0���+�^>�/��������§3�hs�&��������\ZV#_�{�����_�^{|v�u����v�J�����/��Lz\k�& }� @Vd[����l�~��C�US��\|�y]�E~�/��V��\�&S�/��bU��:�[���+��P����iyi�m)���Y.M�\LƵ+���8�`)�W�w�g]X_�Ͱ���8�æ:=u|)&���RL֧342��u¬s�u;��lV.��V�dQ.�S����VѼ9����̢�8J���t��edt�1X��Xn,��}�ݎ1�=���Kv�L��V�♺	�����L� I��:��ؗa>��^�E<e�pCZ�2$�.��H��,���٨��R>�.�v�.����!���˄�
���~�7�N�Ua6��]i	�+^Uv����R�r��c���)��]�#�ͽ������H�*��s��՞()�(9ƖhJ��j��+�{�fMڼwi����<ʮ@tZ�%Xg#g���좤���Ѫ�.�Fżt�/'t~����q\��K�4����ҔEu����'j���F�o5v�t��܂��7}ݙ&b��P�4?��Հ��~�������-�*%PqM���D�HNuA.g�ղ=�lÝ�%���a|�cT��k���e�T?�9��G8�nؒ���j���i��6,t����ہ���N���,@��z/��Y��\�߻ubS�/4��\z�(�]��9by�e^ؼ�0�ӽ]K��wNn� �vq�mɪ�������ө=U��_\�Y�ܶ����|�Z}Fݛҝĸ+	��r��e�WdC�w]�1�Z�v��׸�%n���B"����ZR�{��W�zw���AÑ�Fߟw���,�u�J�T⹔��i�=#/��̇�q�������>~[Gʏ>���k �gn�U�M"�%l��d�2�9Ϯcl�{�~-�˺}���>ib����}�o�gl_9���\�٦~��wԺ���s� �N������ՆSDڹ�8%�@�8�8�ox؆��������9�uԲ*��ǫ�Ss� ���:V[Q^���*~���d�0:O�X�(jT���~��a�꽯�N����}9}�OP�!9H^ �Tӭۺ��#w7������&�B�~����\�n����i���iZYB���z���ٯv�##euuq �\��-PSj��pƠ3�����>��|�~�/W������������	��ϔ�fߕ�9ptijnm����G۷s�������U����4�[�By���54�����B�)�e;Ks+{5��jRr���Gy�����fM��2d�d9]���0X4xt�zVC2G-��4��5�e�ݖ�	Y2�]���i¸:J.�q�g<��q��4+�Q�ʹ���j��5�@���n�`��$>K`�د��,�v�b<u[����"�l��X{�ST8�͂��E^W0�5��ʱ@��
IT�+�V_>b��0V��+f���s�t�*ܶ��Z_Dzo_������ȧO��g���e���I�>�grV�U+ jX]�M���p���k��#[}�LfsF�T�c��B�b�V��>v#���'3{V�ck��TR��Ǆ�V8-��{s*�躶�n������,>;r�S�[��)r螒��t74��{*���f�s�Z���u����݃b: sB�9�D��X�ny1�a]ڽY�gw^�M+�L�i��P�o�����ߎ�h�&�\m��}CB���%eL#{�Y���<fQ媢l��o/*��[y����3�c������C�p�S�T��V���r�&\�ۙ2������G��7��� ���v1¶�ӏ>���@��!�m�p:uܳ:�3��$�Ȟ����w"Y Ɔ+y`��\��glreo)�]v��;(uZ.H�ԛ{�n�Ƥ{]%|�����]��G/5��mmK�a��ݫ{l���DK7��7�X��5j���ӏ�N�̑YY���i�YBØx�����b�����8Ws��XA�+��
u��'ӑˤh
�¸��7
�m���C����7�bN���>��=�j�&r�
�XhTJY<l�k��k�e�>Vꢤ4���3�GP_t�k�,e�v8�0���O�;-��ԩ^.�q����@�%�����K��� ӫKDޙV����TG5̼Nr-R�;���ܛ���2@��
�t3���?c�$0��Y�Bl��n'Ξ�W���|o��Au�pK7��Z���ܛ�i)��,����pM��K@�7+��)��h���jen�c�ڰDEڔv�g7辅l���m:�3>1]'ʍ�s�7����i����NX!�W�1�#]z�b�YUs����<�U�N¥�*���@��e����U�o1(��uY7���\}�윥cf!�S.���i�	9|���z�!Y�qB�tg�vsa���H�q���V��t,K�]4�99+tꓲ�I��ٓF3۽�4�˙�t	6u'T5&�G^V@S�؂������9yXYnr�nd��G�]38q�'4ʶ5��l��*!RL�PQ+�0Ô���uvvv�8KRZ�o(,굙8ef��@�x�ǘf*/-c�p�02�s��)�+���jS#���n��![W,��]������u�V��&�]�kI�6�ӻV�]f�٨�h��F�8�u�ۺ�m��lE��[sh������+��"v7@hu]��u�����v��n;���h;g����c�tU�qغ��l����n���cU7Z�飢���gZ���]���k���Uݛn���Ǝ�j��؛]=��c�q٭�d��u݊�
��ŵ����'Z֞��Mi5ѻb1Z���s�ݝqt�zz��
5���n�5��u��c]�ݴ��u���|�qݚ5Zb�Z=6�n�5�1�1����j+`���ݭ6.��ۋ���&�Qm�ETZ��clcZ�lc���N��"�S�: ��j�&����o.:��#�Gcuݶ��I͉ѭ4wnۣ�j��pv;����v-��:�Vv�GOq��Gn�zݎڻ�t���u�;�ݺ.�]�Ѷ�4u��֧��v�wn{��i��nƋ��&��m�7X�E��������;�67v�gln�i�X�s��Ѯ�,�GqA�Ѧ����;����b!��i�)[#�/W�4Ŗ8�/��=��$Sȷ�a"]d�d�fN���jPؗO�������WwN�8�T#-�f.~I���_�};!+5@�x�e��M5�LS4��NO3N\;Z'�!ہO����e��u��7o}��¶�d�����m�_FXp��M2|��ⴈ�uy�"�A�ԱW<�<����~��N���H�A5�;����@R/%M�6�r�и�I&ܽ\�Yݨ��9���~����\�l���R!�O�q���Jpvn�wedP�3ḦW��U�痖�?\�t�hq��@��-�r�O8��6�E�aӕ�;Z{3��ߕ ;y��ݺo�jm�oc�v��Q����g���;U���L�Z�'���0{{�Z���]�"l�i�}��q��͏6Pk{�WW�к�K�&EZ��N�d�v�̗��G7�0���ͦƜ���[F�5�zF�%�zpwn�޴���^wf��;Z�>���1s�m)�QJ�ٛݜ�{��)�Wv�+s�$6ELJ�e(����44|�Lt�k���p�
Ԓ�!l\�����b���L&:26gu��f��D{��ԮSC�= Y2d��8�\Gl&b�RL�㶍0�j�G�����Q�!�6/tƢ����_\5��
���sWfto�	 ����5���ޔ�l��y�`P͐Fd���gL�@5���EN�M���
}va+���~��Kt�/d���h.�]Nת�5��*�=��2����yܜޒ�{*��{���s՞F���*������T9u��v=yS*3!�5�cz�Z��1uu���I*$�Y̒���¯n۫N��]uX�rܚ��B�1��_�j�O}&�:�%-D{l���6���&K�	y��F�]�F\m�Hxy���D�ὉߥW�"��G���A1��8�r<���z�{����p�h��#��V(�hn~����`#����zm�Y������N)���Y�6OK?C���{�(���*�2�)1�ƫ�#x꤉Fþ�����IX�7����긍h/>��@��X/fD�k�t���"V�T�\9�5�A�c+�������Jgi(�+���|�u��{�ӂ��X�V&���P'}7�-�V�-�2C&��,�1K�S��ݰq��Wqի5a쭓u��MQ�0έ�J٣%�g;tn�#]��c&�V��p��g<�@ً���|��>i�z�U@��f�7P��Q�%���c����35��wv����W^&V���������o�S���fczsy�y��w��K�]{��<�d���|p�A����&��mTtw��u���.~�|e����/�\3��� f�OɇXk0�fD��k�0�r���}=���c��V�r���uf��!����E��C�@d]�-�ع��OQ�j[M
�-������]t �@4�r�R:c��j�!��N
��v��i�QQG�[���f"b�Hl�B�˶�u�-�|�P�79`�|y!=ݳ���^a|ۘ]R*+�-S޾!?���r�b��i��u�[B<��w��FK�)y��c�/r��*��t���(���Ɩ0�2�R���e��;w'�������Ur���
�V}�4L�������ǵ��e��׮�=-�s���v�EܰB+�:�Ԃ��lo��J�d�C'AFn�qy���C��Z��w�+��g{ݤ��1Y�,^��gi�2�'X�ena�ue5YW�+̕��2�yg
.������B�Qf�����w(M�[������c2ӏ�����&�˟��4���3���Ys7�]�>����9��D7@�ɥ�iVR�ϻ��{�RU�3K�� �.V�J�[["��pf:�:������n\h���kK�AK:�#�l3�uy�H���b�)C4�Θ�`U��u)��2�
�)��s�Vu���y�]SU<�D�\��:ݹ\Bއۭ3;k�@�)�ܲ�w��@v��9�Չ����2�~�ԚCnޝ���
Ovvi����MI��m����j�&I��������HȎ�p��N����)ٶ�S��vw��f{3\֣ͱp�������@XNE]aN�+C�oWF�GN�����|�I��3�!��6q{�nM{P���}����:f��[`��X�q�!���#��H�r����W���)0/�[� V�O�u\�鄈�]�����/\U�^e������VV\��1V��T��-S�d�]��<JWH�چc�c]�K/bO
�K�!�����)_;����Ϭ��y"ͥ�U���aAhZ|��i�˝?�fWH���	�U�o^���{�"���7��l��B���̗�-�p�!QT���K&ܑB��f,��7|�F��|��O|^*MWpŊ�W�$2o&�t�2��m��Ρ�7�֜��J]$��ΡWU����D�Գ���>��29�v�����33�R�v�������&FC]�T?s~�} �7ŀ��7�87�[��ռNг'h*�+��
���e�K5��C�I���n�Z����LG9|���q�#�
=�f�M��Ups%A\a��-Vّ����9���l�Bdz�p+x@�+������s5,�]y=-{�Kk�u�\���پɺ�j�.��!��Os6u�wJ�~.�.Gs�'�P��E�*-�Z�ey�?\,L��g־�=��
��LA���d�h꜈ ���:I���B�gõ��ò͐���H�w�/�'��_*ж�j'XKN}���F�i'�^�n1t;9��,C��S3�E��F��%1b�����Q�P�2<�5�ƛY[5�.��c���[�h9ٖ&
ֺ�c_U�vU����0K|"_�A��>P�w����f�'�������L�[����^cCϧ�Y_:��{���`��ʽ���cuV0LY6��{���1�ݫ,�YB�6���	���i�;6<�baLbÞt�p]����O�-[���N�.�����L��Ӕ �-�䪖�i�.�����^i��ݶ�={0�P���z��ǹ�hlDoU�@�i�����]y��ʟ(mM��֞=
��&�`̫��Ź�]ɢL-?ǝ��v���E[W�p�Ә���Ϣ�=��]54z.8�T���˳gxg1��1CH�T�]��9S���}������s����L٭���=LA�t�j
9Y��77GqUV�'c�U3m26H��[p}���`?�rjq����k�N^���IUk+�^K2�Ӧ�mY��~����lu��^iZ͸�F�e6�+V�~�^�;�v�:�7��=s����uzH�g/�^V8q�#9�pU��fc����,����������b�<UC:��׃����{����{��;�!:�f\��z�*��Fj��pT-u:������8���E7nYWttV�wV<����-�\�!�����m�v��� PM�mCK\̭黊�I�P����i��b�y�@��Ȱ+s�P�.�IMϵe9��{���ui��j?}��Wޞ�g����T����wqq�r6u"�(����<����w��MKw'��P��;[@�?!�۪��1:���6����	�5*&H��;yz��i:�%�U��V�<4#� �bv���ї�Wn��p�9,��D���&�O
�H��Ֆ��B�d`�~�x�H~Ƶ�D��yuLxg���>��wU����6��
�m�ޏT���|%�P���v�r�Ϯ�Ħ�H�M���i7Lc��>ܐ��S��%�b��8遙 �F�I��|��}�>��Ȱ���z�fd�*#��2�3fN��%�#���4��X�����k�~�d^=�E�WP`8����w�6��K�<xw:����#��i�Ԏ��l:�t=^K9dA�ϰ k9n-��q����&vh�֐�r�1��{Z]��HxZc�v��l���}�7
 V<��gV�ۖ���9��1o��x��T�\��t�M�^�'0�f��1�W�)vz����S2�I�Go��y���B��d�oqD��â��Jo�>��wv�b���E���-l�V�u#e�����k��|����K�������720�;adG�HO$��\����Ɣ3��2�o�/�kWF��e��QoZ�\��"��9<z�\.�.{z��dCGCVw6��|�^Uf�QC�T z�B���)�*V�}��^�c$^T�['�=�۽��ުH޼y�eBr5O�-��Yhj�'8d6��h˼=Fkw�����]�W����lS[�ː]ʯKS�����Ut�68�#
����Q��Ƽ_h���%{Py��|���gB����<2-9�~�t�u�1�K�8�N�(y�%r��4���p	W��S�\t+�A^��X>�9y0�Ȉ��	���9o�b��PJ&�]��utk^���O[�����8K�'�נ�n��3�J�ζ�M�7��Sݴ�꘨Y+�H�f�w�=��pmض�6q����-�G&�ɮkx����t����>�1u�$:q��jw[c�f����*	|jeL�[}�Hf9�5A��|���</�:��](Q�6i���e͊�e�l�uΧDI¦s��7O�2%3��r$�,��9A�p>����yo�J���i���~�U��r����c6������� 1������~� �ω��}��1�.���z�L��&v���?H��&�^/r1�'g����Xs�|	7>}��s�^��s��n�Bk&U��ܩ{(�)ܟBIVW��m��qޯqk
���bg:#�Wx�����3;���aF��ځ��x�T,�{3%�t�)��!]�u6J�g�cJ��m�z h·�����3,�.�j�'�|EyDݑ�/�ht��މ~芻�t(�>��3�ϕ��G��-a��&�	��L�#��ڗs�[�xLNOI�v��AĪ-�2��X7p�r1pK1U����8�x(��tW�����I���4g��9�fUx�x�e��-�S��h���P�������NWb�:&X�&�\I���T���^���SA6�~a�[��'���3v�N��icJ��^\��ޣ�Ф�z^֋z�|{
�w
����L��~���sޓuEܴ�+rI�klr��t���?gD�.p���*�l����n"s�5޺�wfGD���qM���&�B��,�q5���׋$�rw��w]A߫�V�"��|�8�>c��/'v�Ɂ��:U4�s�u����%B���!��#Np����o������]M?F��d7rz�{�DK�M܀r�A'%𿝚�]g;-u�mj���WKn3:5�UY����?VN���=a�@�)�q����k��(����|���Sг�z���v��/�a\�Vei��u��Gk��6��,)o`R��oZ�x7vM��n5yG)�]��o؋l��M�;�e5=i,Sp�N�_P�*tax�:�ul��J���\��l���nq]MF�1���x{̝�E(/A��3�Qy�b���6��3�����L�w�ڍ��\[%��z�[?W�L��e��7ʆz�0}�o�FR�́��9����$	#;��Ё����4:� _ww�_������w����q@W�
������TQ��
���8���������d%�	�	�fU�VeY�fE�C!(��3 �#2� C" C C  C( C C" C  C  C���|� � ���E� l?�X@��  a�A �=Ȁv åȀȀ� � ʀȠ� � � 2�2 2 2 2�2�20 0 0���**
��(� CJ a aUa�U�  �D �QU�!�eXeXaXe|eLȳ
̫! *� L�2�ʳ *�!*� L L�2��ʳ *�(���������H�����2��0?�@s���u����7��W�O�������P/�7�{��G����;����o?����  ���������b������ U����?a b����P�� U��������|�އ��z}��?�O��o������o��  ��$�J�  P R  J @�( P�2 �0   C�B  P ª��H\��@�@ J��J���  �����  HJ�� ���J��*�H * ���C����'�
���(�B�~#����/�(>��������O��@W�����ÿ��~C�D���C?���c��rx~��D ~����I�={�O�D U�� _�����~( �����|�" *�������x���_\0�7��O�x��_�� [�C�?/��Q _�>����?�?��?0������	?������@W����h�������'�_�1�`�O���g����>�z�o�I��|" 
�	�S3��~���<��A��o������@DW�0~ǂ��������|?���C����(+$�k7��T�Oۋ�B �������/+�=�J���R֕Z�EHT��EJ��J��TE*Q�ٚ4ٔ�����RP����YTk�MU�ڦڵY��m�cm���+j�m�Ka��l��mKj����Lm��[[3sX�Zm�֊Jk[U`2ŕ[��Ԙ�d�f)Y[i�Kk-%Mm�j���hY�j��7Bu_  ��S[m��9ʥ�c��*�7*��e�Uhk�.��)u&U*��nR�-kCwi�`�Gf]۱�5V����&Y� o�袀�}݋�ϼ{���Ѭ�5�k*����Vw]��un3�GC�,�u��:5Z�.�XV���[m�g| ��t�gժtn��ۮ�Kb�[Z�w ص��wv�90�e�ݭZ֘5�,f�5Zڳ6ۼ �{[��2�M�k�Aul]Y��9�nEj����퍥�:����]Hd�mvٶɍmlkU
��  @�{���Jĭ�l�2k���E�b�N�r7wRٴ�M�*�9�5�n7:;��6���� .��mX�nt9)��%�9�Z�g&楺\ꪥ�jSku�6�`Ӷ[Sf�H�m�6ڪ� �^����*�*gU�k�n��\eT6�Vѫ�h�Csh:$.w W(]*��&��6��=� q�R�-��Pw\� �[@�� :gp t�� ���u݀ [���%�m��[� =�: mX� ���@n� wg R�� �� ���.��Bm� ��4ֆ�"��x  �D� <�@�pt � j�#�� fb�PX�T�0 w�=�    S�)J���0 ���0�*)#& �d`�F��0����JUPz�      ��%*� �     "�&� �ѣ$4'�bh1���e*�� ��@   n��Ï)�g�f���r����X�b��E�=YD���ʓH/������QP���k%�b���#�� 
/@���E?bA
��?ɏ��~u��0�a@EB	��?���*�4H��	XTDT/��~3��U�߿����H��&��v�\D�vxO;�Te�H"w�{14�f��۔�^i9D�F6ma߮hM?[#Z�6���-J�-wBK��V�ڲ�S�@Jŧo��.�׮��9L����!y��5Q�$k,]-	��\+��]q7�h�/����ۤ�+TuaX`+��(*H[��ݴ���w����(R)ѽͫ�`1x��"��'�ͼ�M��w�����͓��Y4�Q%�E���eSI1{�-f��c���;tkp�,?i��B̭ �vU��5M�wHJq��ݨ���b�ZR���^bb�3p�i`�[����Pj5tN��6�#"��rk��$�Xٍfحf�̭�	��0P?

��PRҫQ�R`�CbB�[
m�G]Bq���y��^L+sC�x�sj-�Ѱn�DQ���;Y��wH2��WU��3����#`ڶ���C�e�lX� �SSX��.I[�e�*��u71 �1n�D�;e�(��5వ}f�ͦY�N� �f�n�9�P�RdT�i�7h����9�R��s)�h��n\(��H��]\�u�j݀FEɐcU*8�ݤZ�1*�ţ�/2����l^�b	�p�1RGn�j�*�D�{sV ��e����5[Y��n^N/�nM��FoQ��n�K1� ;AM���l�k���U+Ӧ�`��p�1�Z6Tťږ�ހ7j��zu�3N�)	���ov�,��@�z0���K��}���Tq]�
�(�z�FJ�x���B�j,ڹ�(�L�u��U�r,u�2= ZV��.hLַ��b�00��H���[L�8BI��-;O���x@y*�X�[up:��lj��Ǵ��W�1ڨ����o�������r�eQ'���ݝ
�n��+{7�f�[ H�*̩4ni�O7M��`1 ΅�d��ie��7�'���ȷE
��4ͯ���Z4�ni[6���������BQ�t5�x��ܥ�A%�;�2�I�N��h�2cb:&��vf���u$4�Z�!pUb��hc!��K@�hM�
�,ܖ^QE&�U��z�\��d���1�b׷�n���
�b��M'4V��YR�[D�+$]�s��譫���L#�n�a��E��y+Y�:���m�R��b�j�ۉ�1�*�X.��tb9n�in�B%P*�\#6��:1Ғ��H1`f��gwp[*�`5���ea��XIA�5��M��B鼂BY�U�B�_'���+U����i��iif=��Ս*r� e���Rf���31-�t� .���ސ��U�$S.eP�v�ڗ)���i��R���VdV��
�Q�3S9�a��v�hNi�e����u�6����U��R@e�6��O]�jۺ
���x��)�6�ܠܚL�1:T.^n�Y���3Lҕ�H�WUZ�We'
*��*MYI����a%e���Q�j�Y��`�ti��Tn2*��,��(�֖�b�����Mן60nP��nM�L̠��n 5҈���.h���((Օ^��K�nG���a�V�/
Y�h��mQH������Dl�e<�i�9A"]ɨ2eD�P���gck�1^��-�e��qA�+�I���#�9s�ڍ\�"���$�u� [ͺGZX#�Hs�QYM2�d۵D,4V�hy���kF�P�b��vZ6�ثu�ÚuQ�1\�$añ;�
�d�t����
9���V�ff� qֈ�sZw�k1-N��>�!��e���V<��C��݈�;��wBTIɺ�坶2򃶈C�U���Э��n��xۘ�Q:+�i�[H�+N(w[ߥ�{�AYE�=�l6���
L��ݬ������6��Z5�ޅ���ɐ4�.��ׇ]�V]ݼ�Y�)�Ȋ�f �URHȣ+2�X�,��F�uZ�B�+���cGy� ��<�9 F¦��Q��/�ԕ�e�b�mP�s�9�-7��o�:f�Ze���S(���9J�TU/p7L���.^�մQ�`�!F�*r&���fT�iôf��R�VՌ���]v�&�K4� ރ���񥌆���O0�����0��٘���
v���x�:��UJ��Wx7U���^�m'�+Պn�j�żY�Ζʕ�,vUu�mT��T�Y�W��M�HO�dn����Z,�SH]��ˠ�u�i܏p�٨��w�,]��w�����N��F�8��pQ�ɣ)a����*xUf�w�3;U(e��H���LjRe^������.��U��!����e�ԭ�U��@�R����:r:⾑V��{طJŶ-7zY�dSG��2L��SYӹ�S�H6�\��훡Q�f��2٢�'F���*�u�Cr������dovk�X&���t̛�Z��� eaddB�Vp�ɬ�wpn��2"5T�n
M�kݳ8�
vq�4��Ҩ��ܭ�1��ۺ��e �Q���M4�mX4�,�-�o�����l�������3o7㌶��{���ܔ���j6��l���x超m�@������En;*e�/Z���4�!�&hY��4u�B�զ�Vܠe7Vn�ť{F�Ce�Z���QY��ݶ��iX�Y&��4��++\`�N��n'��*�l�[�`$Чi��3@vZ�yF���!YbB�MP�ց�o5��7m-sڥTc˙�/Ff�*��Rя2\e�W��J��֯e�f��z��fY��PJ�F�edu�o*ͬz�-��V�<����Y\w `��o/͒]��[��c�&��ѕa@�Ky4SiU�k6���۽�'r��kÂ;M�dєAϴܷ�7w5�c��"��j,PB��F�A���	D�ѧ�m<�#v5�(��Š:�ݦ�U�a͆�*'[aUz��xF�b4b����WI踩���m�w,<�H��3X���	�f���x�������$F��nh��m]i�V�n/�	[��z���S5]���y&V�u�HT�A��ڙO(�؎H��y��l�t�����z� ���%��jlk7,^�GE�Γn���TL��\���:M����(��\!Ꚅ�I5f��{�_cY�ϗo�!���P}��(ҙ��O	h�7A�{�*�#Bl�
����n��%:C`�c�i�� ��4b[6���$T/tZ.�ԧ10�VS�Z�K.�M�hA�֣]���)[��6h���N����"�oI�B��r�n�ݭ�f��fdL��4�E"Ŋ[)�$GsA��y�9wX'lůf��m����D],-:�8j��l.+X�K�']V�2�i+?A�Uֱ��v"[�6՛����E����]6�$��UȪ�V��������2�ЙUj�(�/�+���/F���B�J�{��v�ݕ��[��ʶ��xm�e2����%$�om٥. �M��b�X�'ǹ�������YF����vF�zy[�ZT��D@ۥ1nl���gVn��`ӗet�'BƘt`�["�n'�؋n�� �!Ѥ��EKr]=���3(�
5E�G�D�q��0&B{%��$K֠�,��)V���F8�ƚ��b��Lc*����ac��q��itJ��L�DJk�҃z�E
4͖��V�V��`ղ���A��x2���I_n�}y�RE��SǺ�&-�ˇ�q�GxC-�X �j���V��H�J�^Z�Li� U���!�]Q�[Z�h!�&գ���a<�,!	���AVUǢ�u��Ӕ^�ZH$��d�4��)e�sy��Ե����@ml�S~�x��7b���t�4�*�hWPؓ�ib���V*e9sjk�a�Fhs1'Wv�hH�&�"�%(*�G�B�_��4��YW[
�L技e\��,�mM�E�yvȹ.�^�a�3�#>j:�Ҥ�F��2���**ͥ��%j6A9��Fԓ20&�	r���v�^����S �Med&��fX!�eAnn�Es8�\ŖV�֍�-�k-�8����D\vH�-[O1^��!w����V���0f��T����IB"yZy�~yp�0?�X�5��ߵ�l蘋+�Q/Y�oe�F5�!̺R1vê;��J�p�dW&�m^edf���Ge�;�Phܫ�,Fe�V�V�{�Љ)����u�e�f�;M��X��U��Zs�fݵ�\=n���ɂKWp�r�<�j��+�z�C5c^��
Q��8���̨B8�-n��6ZۥMӽ��8�/p���2V��0�(��B+��n�z"��
�^lfc����OsvJ3c5�Hb��Py�'!��)]�30\'�6.ۨl����Fc�+�D�mo�3�9� i<��i���+j�)�SOPy��^�衈.@�&Ȍ򈁊̛�(AcaI�m���o"��d���B7\%L�j��a(L�	7�6Vʀ �w1��T������=b�`%�L�A<���h�4kn����F�7��ϡ�Զم�h�,������v�k0V�:�Dٽ/QFƱ�c�I�G��:��Y"��xu�
7Es5�<�iBr���6cz�;��:�5}I�S��b�~��#����j�#�Z%�WL�x��
�Q�ci�e��h�D�*5�^qI�Ň�r��'��F�p
V;d�ܚR�!+6��m�fFZ�y�*)�5^�*�-vք2�Y5�w#|V�<jgmf�l�X�r�;@�˙�me�V+O2T�%����?4^1���y#w���,��7Մm�+ڼt�9��!���Oe��R*�N��"yeS&JW�����7���@��ٖ��=����cW9A^r2�"��3�+.�5/R�e��3dk��H�C��}�b'�5�g��.�b����x��ҚS�r�]N^a0�k��m4؇���t5���z8	ί�K�{l��*(��
�]��D`�W��P<Y�wR��f�p��܆�^�0a��3w%'�:<�h�v6�ի�טr�v�'_#(�� jԶ���%7>��L�I�q⛡�gt^�]�"!��L�Y�n�q`�xWRЙoh�]�"�S�"�[�fV�H��5Mgi�U�/ZϮ�;�*�uv_	խG(���J(򶲭�fl�0$5���%�7[X��N�6�,HQl�P�õ��Я:�a'���4Wۼ:���;Q�ӕ��*�J|����.��lN�ǁ�%�1�bz�3CO���*)�-���V���Z���NEY���ۧn��6���)mb�-���G8N�1��x�FSJtw�/�d�P���[f��M�C��b|8�wS��|W_��Ʈ�pT��@�E!���6��f�@�;vE�gi�$���:κ�m�*(̶4kӁ}ilYCo�M��R�]A3�s״
�2�l���d1�b����>�J�ᘃ�#
��Mǔ�ٲT�{��Y���ֱ������;c1�^:{|9!�У�W%���ԡ���+T��eCZ�d��g5Q��� [�����,�I��)v�P�<���7g-�hLj�o��2�x�)��,U��]F���5�I�u<T�i\;^QD(��(ش!K%�[{.tvet�_\���ur8�L]*-�T�N��v�{z�2{Ė;u���1[t�ʜ��t_Z���NGs���æ!���55U�@���Q����{�-�ibP.t�П]��ح������4x|�1]"�K�.�ULͥZ�(*�S�E���2��]]�7QF���2=�=]ʺ?wo�mi@7k�޻�	�u;��JX%��Ԟ)ݑ��W#t�.X�AyY���e������������['���Z>�W��������$Z���L*�m3b��5�e�Ԋڧe%6�ګ).M�]l�����$;.�S�ݒR�V+D�K�۽d������4���f�NW>��̊��"��Hl�W��S����-����,�H��G��hPvet�\�c6�� `k7�k��
GV*^Eק�-ྭ�e�PTs,�׺�pF	o���V���m��M�O.ξ)�¯��P.mZ���p����&�`-��]I�H\�.�2�%�z�g��n�4�V�}ӏ�Kl��u�����a8F	E��J-�8�23��
�Z�С�p�xE�g%����l���Y�1�c{����k��En�WX���.v�S��d��fXq�@7ϯ%�[q��ovȽNZ�MQ�
�����b�.�VvI��ʣ�}O6Ȭ�Q
a���LK2Io�M��W-�s����LNҢ���(K�GnX��``My��"�[r��(�3F�����pS� ���&ϱ�3:[�`݌�����j�H��N"�\hT���"��]CW]Nv��$�vvNT��-��D�!u�c�:�yk�J�yxLw�^C@h6�U����D��0�7m�;���	Eȉq��T�C�uv꺒�,�Ι���B�J����Kwd��:�t��d�;���V	.T��l��AܗD�X�+����@��Cݼ�8X��z�m&��RXv�g��MB�u-�\�V��6���]�nV�Vu.[}��h�+6�GtD�xH$����vtj(vb��@YX��Ū��}��5�̔� \���-��*�j�w EKY����z��j��h֗Ø���ه�x�&u#�!�S��eM��d��B��\�jl�B6�ƺZ�u�%wl�ͧ\�-�Ip�QWZ��պ�g���EQ�c���$;iL���^<Gk��	��m2�s��Y��c:�#����ώlTk��K{u�fn��ղ�o<+>� v�.C�(m�q�ͷ=�P��^`p�|r�8�aV���B�{
s�Nh ��,M���v%aYp9m���FД']�+�j����Ԗ=Էzl5�Y����
 X�y��YGZ�H�N�v+8T�zö����[��k0�����JzJ��nKp��tb�{�gϝ\��TpDmp�X���΋ec3N�3��>F�g\�c�E��ܑ���WL�U����xp`�c"=� U(�����C���Ӓ���R}x�&��_�(J��)�Uo�y�+�T-P�H2@����m���@m31�ds�IP�e����2���垊e����pA��Gޱ��*� W���n�N�����J,k�P�������@)��
�G%/��y�hv_Y�-C8�3��7�*�r��Js�t:��6Pw����,��r���I{FY���{Ν�Yu�@w:�q�l�����]EG��N�hJx�+��֍�>8@�i�{u���
�"�*bK�+�RR��*���-�H[s�̜���]-��N焭���Ir�M�Ɗ�A���Y;^" �=�o�%�ºڔI0����O/j0��ܻ[KF�+摺�gy��c�m��v��Q��c�X,r�ؕ�k*�7��#d��,
��e�@��9���m�"�r�x����a�}D��{G���
�������m>���P���F�2� j��|zk6��<��ԣd��~ۆ�Ar�\��w�@0����ou⛸���ز�W��4*�8*]��U�E���4��>�Yh�
�X�<HV�ZM4�Q�XR�W|��h�\�O1֩�'��!$oF퇔�jT�ΏMu&�oP��%��5�%�%�0�Y�FN�t;2��^��u���ƕpH'�vcܭ�}-U���d��}�u3��Vf��R��c'��-.�+\W��W�-�q��DЕ�
�B��90WbfN�b�*�v�:c9�y�b�[�F9K�'{}&�Lbz���I:^������}ʶ��
�K'V�ɵ�E���>�Y2�0�R�ڕ���mT�w^�#꽀bN��9ZtVq,�p��묫�k.�Q{Wa���s�.��Wc�ac���к����Ut��oo�9��#������mv^gi��	X���y�(�x���`�a�8��Y(��U�� �v�������TT������kI5[�aṷ��N���_��<)m��B��Pc�lt�o��u��M)��E�涌��Ԝ��IWZ�Ҹ.6��ь�Zu�ܾ�k����%�XN`����S-��RiS�X뇸5W&N�\�� ��Ғ��vlf�2���#H]Z ՘�ͼA���{]��t�Xyy09X1V�	X�7��t%z�⋧t���R��ݭ"v�ssY]��[���R��,˲��Ew���
�gٸ6�����c���ҕB3&6
�Op����.�ʑ]�X3:k��%c���:�.���5��f�'�oz�9]#|��Աݮ��<-����}+�PM.CU��j�cEm�ʻˮ|���ˎR�`�^|�����MJ ��*��f��A�v�w��:\&\�1�ԭ�3��-+�z%2�/�s���M)�����o(d��̫��T��_g+M�h��]�sծrPX��҈rˊ�C�aX���S�]�;�������o6��`
��S��V7-2�5�ӓ�ܝ��`�'te��6�k��Μ2s�zXt�
!.s^flE�Sx�}�%�(�,Q�Ja}�6 D����c(�d
��P����ut�wl����i�y%ʎ[�M��)sY��v��8(�Z�/:����]j�@�Hn�'2���cF�5J����:'�}7[�w\*����b�flF�ʬ9\�&�At�)�#�w[4*�5f'X�+ u��c9;`�k���:�6iL���ɓ��]��\z�ʬ�V\�{��O�YNf1+'Q���~=��H>�j(�h%��K��	�4��YMď[Ý�T�+8�d�����7$�������A�q�nzқ�ɷ�A��Z�XPEP�|�)��b� ��I�C�wF�i�?*_�V���;��m�9â�bk�Y�^���κU�)���sEuL�d�ݡ�W�pw���=̱Fd
�n�A,��]��Zlq�3J��WQ�&8Z�4�)^%���
iy�4p����PT�Ø�L�8�h�H��a���1$��>h�-�+��ôX�Nv�ǹ���p��2�t�j���et��!j��l�x-��a��@k�-�AR@k�F�M�B�4}���{D7y�s�Q��I&������\̽W}|��v���P.�����^��;z�Hqq��'
9zt��"�ɺd&l�<t�A�v{ma�K�q������і�n�n��H(��Z�t����{�gkR�n2�FnRf�/5Q
�Ի�Ao�t�_$����g��;{|>�wJ��tGF�d)��"�C�Q;Ө������}�Bo�^⩉��N�sR��o���^m�+�-G-m��4���*_',V�z�4�+�:�z��or�S�����i%��P -��e�e�<:�KV[
)wv1+%��![\ <ݑV^�V�� �x���Z���\��5m�H0���c�Yz�Ns,R7cNHU���鯺�َ(�u��xXnM�T����Wŝn<$�6GQ2��&�����P��7�;�N�ںv��3�wV�*����B�Q;�ؓ��Kt��5a)r�n�����覑�F����ʅ�`�PR.����M#.#�>V՛=��M��׹��P�����tM���{65wAkOB�5R�����lp�l'����Z��uS��8�z�Z�뽹���{��6Aq:E���Pv%� "jf=6��܎N��A|�!*�	����cpΎ!v��żYڲ{~�DT끔�O��q܁�ݧr�g�gt���Oq�0���&��'&c�����M%{:A�՘o	�k�������Y��N|�kE?<zb� i�9uv�G��Wp��֮Y��^��T����r5W��Z���m�F�H--5���U�5yRS�T�1�:���T���4�ES@7�WQ��qN	���nj6k7��ohܣq�-s_#Y���gb�5����/iF���c�]���ӊ��T��9P����s�׹���Y��"�ج��ޗ�x(�d��"	(�7�s�zR�$mr�m�ʸ�R碑�;�WIQE������r��t�C3�v�����@eKJ����YU,Ǫnpt;��O�9lg(�N�$�2�
ͨ�7�%�k���M�qr�u6�Qʖ/JS>ct�2��=�%���!�s�[Aj?Z
�ۗVT��|mK�:;��(.���;�+��4��,�u|Hv�h+$*�|h�'I�Q�k,Cl����J� XZ��cz���Ԫ�|;4�;�Ym]s|�5u���Ɠ���R��±���ynŬ|��tl^b�]_<�$dui�ʦC��%�Mj�N��VVnp���'ܨ,�ҤB�I���B��NH�;ր���N��1�V߂�v�-�6]�EY�%�0$D�:�w2�M�e��
q���2n��-yWv/��{4��Qhh��pA���4�v����L7ͽ��X,a�u�5ʦfc21|�L�q�&���v����x���Nlnl(��y�o:�$,���\���Ef�ab��7qC\%���
�����d'X�V.g:f�B�K:�(ٚ�#EIh�.���.�7�����
��E���I��}�[@��b�j�#)���"�<�r��m�}�R�)m`�(��t��D����Dp�*4ualg<z�Y��v���p��	�AKCB�-�Uӽ�RW �*9rk���;j�m]�I]�17z2���:XT���Mw��Ո*�X�n�n쾺Ҭ#Ԏꔟ]@ ��[2�VuZ[�R�R���Xew*�@Kgf�G��I��m;J�8�o^ܡ%k�p��Ag.�X:�aj���0�6c���h<`�5b�Z��vѝ�&�>e¤�qY<��+�D�o�RqS�e�P�@��ob�V�L�܂kA V�5b��-k�n�޽=@0O�Qʋ5vܗx�rw\��H!�.�n���A�N�jE��c781#�]�<�7���^Չ�t��4�Ϡ�n�{�ގ�Iˋ1�۽�9s::��Cm�nb��җmIk($�r���m�L�+��T#���Bi2�ݤ�@ӷ٭dKPA��Tʼ�`�aWC���U����~M�t��9�ZX�t|c�{ �(���e�]�[k�Ch�B�c۪;8��>�/B1@,�!dӌM=⇠"��kKmdz��6���h��lC�
�կ��'5[�"f�FU= ʭ�TřC�e+
b�l��Ę�]��]Q�EWS7�n�d�6i WP�]��c6Խ�>gm�E؄�����:�Sh*��mf.�%���r�<���[��n���%`F�Y�h��fC6�^�͗���ӯC��ɬfˤ(�gf%�T�z�5�Ylwk�:t���h�O!W�n�V�u�o>�x��c�#�;A�)wDˬ��7��ЖXwWZ/a��O5�լ�����6i�����l\���Z9%;b�����m+�o�g�0�h+��Ձ�L����r�+;c4�}ë�7�������gU�<W���k3^Xe �_%�0�$s{{��8wX�ڔ��i�CNf�o��)��)�{Q�M̢������%Yǥ��*�5�{j��u���5s�N���ja@^�G��/��4�nr��m=�*ݛ*�%�wvVWU��cHs��x�]����V�%H��`d�n�PJ�B�a�tiɘb�uw3S����m��e�ݫڵ�䳙�7��ħY�x�}�k�j�R��ൽ�*hݳ�8U�yq����^�L��s���$��)��Zm����w�`��+��h'�R��sij��#���M�5�#/f\�v_�2L�pD�%,Ʀ>�업-�G�����Y���E\{�3]U�2�L��9h�LX���B�p�ْ�9�ƫ�4�&U}�Y��:��O��$��z\es'q�%uh13��}2]s�]ž�3������ϹݔKżݻ9Y���7+ep8�$J���B����(kLs����F��7��f�};�f|�t]c��ܠ��=��w-͵{ӓ�rC�K�l�2ET���0�*�u�X�q��U4��3.�m	��`4�T"����q�f����%u������-&�@��ƴ����9�ʝe���)K�de�:�H�.�J�6��5��6�Ƈ:.��}uה�Y����k4dAMb��.<���+�PHne^��J�g9�Z����%3e5i�a��]*��{͈n�RF�nԻ�N���pb��p����
�.��n\.��0[ܼ�MC��&����l���q2 ��8u�����cv�	%�N�G�-6k�y�R
۲�qS���\n��++���u*��j<R�7�.�7Wܛ�NDAv�r��Ǖ�1�&�l���pֳ�֎J��}ʮ'O�I�3��+e��g�ʭ�TE�u*�l���{�������	6�u���J��8�Ы�2�"2���.�iT@���..y#w�I�n�@uLb��WM���A)Y�wo�r�]C��$ۚ�7�����YMj�����Q�'hd����%̙Ww�wY��
����3�UgXuҝ��[�SشL���c�iK=C���fe]�A����5@�4j��N�9�j^���J�����j��7RқS(��%�3d��5E��Wmރ@��H��1wS����b|��x詂���h��z�S��E��>���� ����z�0��;��ѩ��]��P�kD�u�;��H�Ki�������DҒO��#��1X:N�+6+�΍��%a;u�y?����ʱ�[WK�tGLbƠS�.��c�=F��
��ӓYV��w֪�$gϫu/:�M�n�,��.\l��A�sl�lJS�S�v�'�R���@�45\�Zu������s�/��M�N����,;/Z�6�R���ym�*z)[Є3!-`��$t�J�`��a���h���Qy�N]�cG�.j���q�U┮�]��,FP�:�W1���m���ٕ¹f��Ya�4��[f]k��vy��l�����{��D�%=�%��|�vR_.��v�ݳ��eLC5c�~�(1�]4j�"�<07���܎�)(W/�쏀�C�"���� �j��'�V��
�.�c9gSu(R�hZ�w�"���A�5t�\�T:tvI
����	���EAaVe'y�&�M#�Pg��$f�N�̡����g��B�z�^�����l;�b�>�e�\��1n�,M�h���ie�G/�v���Nt��g��{S8�"g<��w��܈�@A�B�E#+�L�CR��ٖZ�0Z:@B���u�ON�)
u:LT7���h&CL^spd!L�������e�N�3�!O��b��q3M��p����S޶��}eip�X�73@�%��O�/R|��A��S�q�����G�T�}� ԕi�Ā6���i���wZF�(�-�]Y;j'�����wmB��`�ē;9�*����N]�����}�]���U���&����쭴j����O���FWT���%q���5�fJY�;�,۸LD���\���z"h��l�?
��1y�{D���wg,i +�cV����v����{������:�V�"�X�A��ݱS�@�<K&��X6��Jq�f9�X��-��Q��	�(��qF7�j��Uudr��QtǺ�=�<_c�by�g�����}��  >B�(�4P�]�9{���N��NQ�'N�
Ќwn]̒�2uf�wU'3�R3s��N��'\�i�8`P��!Ŧ�D�y�,�;���w���/��8sԜ����M��J<�1�;�z{�˫p�"����8���[�$ܝ��'����A�D��Y�����,�����l�a����y"{�:N�w+�\���t]Ԝ\��r\<����h�\uw	�YyrnL�nYj��)���dh���3��Iu �G(�S�rM�	�EУUB�Q:r��,i!�2�������eF��Ebd��j�PA' �hU`�Qʍ.�P�5L�z���V������?��&��q��"���D���:��ݨv̮OĶrB�GXz<8_#��J�*^I�>�������Y pT(�OƼ
��bh�&8GGq�Xx%���Ԗ���t����?h�Z�+���O0������S��3�C�j@H�I�� :J�:*�����j�UY+�)��?�T�p���Oӊ`q�Fk�(ţ@pZf� �Hj:��λ)����>�yx��^��xerUK�����Y[��+����\���ʗ�"��^�hW{u@!^5{k�{s?0jj����r���ͷ��IpO��
�Ȏ S���.�½��ón?k ē�Y�.v~��!�Up��ey�����<))ڟ����]V�fT`|b�o�0P�C�a�۵9{jp��E�%:���y�}8Y�Ǫ�rzj���E���t��D�S������4�(;q�7 {�<��yKi4�u�G8��,!�r��F�[�J�E�0ж��E���3%�a�D�X5���+^�sӕ�9�3�2�bC�a�{ӂ���y}��Z �]C�^��VZ�*�=�k�,�'�`Vaъ 1��Y�!����P���1�s�����Ns�k|�Ə��"����v�k�P-��c:8�C���7}|�4�o���P �";�Ҁ� �l��Z��/�S��o�����!���8E#� r:Ќb q���#�/j�c ,��ؿ�A���_w 5�Θ�ML;D�Z ���l	��x�C�F0b��ß�]���Q�(Kr��LW�	��)��'o1��#�d�#�QE����18¨���"Q�B0FA�9Z޻oR[[�Y?\������)�d��ۖ��@S����"M6�9r޿�)#�(�g��bjb�2�8x�x�
�, �󙚮��?�Z0���W�a̺��Y\>T����>"�47\�jz,ԩ�nV�B9�����-OPP��u9˚�vɺ��x'�39�zwd����BϫW��X� f��1ֺ�uƪ�^
`���߼q��z����p�4_�]*�ņ"���ᠱ�L�WRX{k`H��J�]��)���ac(S���n��Pk*�0��RFc��'0���fD��|>xts����MluIѨ=����\�{^�l|��dS�ň�$����4`���8�F��D��k���0��\A5W/�
��~���Ը����tS@�]�����\�9�٢x }07L	R�Y�ӱg�ܘ�&�֦&�8e����1�r�A\F�A"E�,Dp�ݪ�\�ʾkl-L:�눱^�q�F ��i�5�P����|�n�I��Wݭ�����"D ���M遦U��?�pi��,m_��D�z�Kk�EB-\&%�		Mj3bY[�AϬ�a���p2�}�v*Ny��2M/�PTz+�.�D�-�6���٘P2�������NY�{�t)w�=���T�8F<���Vt�盭�$d(c-��~��B(p��l!���?!����3���Հ� �Yю�cG���V�V(��|�P��������(D0qURqW�?u�Z5/K�ĳۗ���k3zb��A�&!����< �!�w�Xx���tZ����e�]�ӯ��։���7Ł0� ƙFl���>�  Ɗq	F�=7΀�U4�ӾT�"���< �(G	9byNN�;uG\v�����Q�b��S��BM����̺�yF����5ck(If�Lq���g�`�!�>Y_R�U0��Y�u��G��|Q3{���j/JT<�x~���'��f9�<�3N!��Cb�b�;�X�F��֜��$�� ��������#�l�>4!�yY�w�0�&\�� Uɽ�%�[O*�Bk�1.f�J#�fgeocpNͶ�'�i�-�o�Ε��Çxh�T;�
Ў�7����,^F�Rq��O�PD8Á�A��yX��U�i�U�µ�lAf�����O�j�����{�m�*�6�����Q�Y�-*��v����mǼ����WN�2PB��5x;rDdp�w,N{Q]���˞H�]�U� .8�ʊF�8D�(N\�������r����#@Ҩ�R@��@�E� �#!F0D��5�����5c��v/��T ?#�͝L	|~۩�o�d+v���I�cZ��t�f,"c��&4�N���'^�9�\�Nu��X�T��N��Y�� *���6�Ya�qw��%ͯk�����9P1"A�������۔GL)S���~��]&�m,�L�ޜi�\���Ӿ�:����kc�[���U���b�t�U�7,-���JS��p �2���9_.�����<��tyݓ	��^u�g5��'4S��_��_�4�k��G~l:~�U�@�./;X�.a��7Z"x膏�X��ɋ�F�����r��.�I�ו�Z柽=LW�T�P�-�f���pT}d��A슨S��\d���⻮ֶ��G�8 �i���c���q�2j@�$X�N�1����$y��>�*�\��V�A\�s���Y�W!�p㞦��X��"��avtR��Y��gG�,/r�[���ٻ������%�$��C	E�v���8)�I���K+�2H��M�]'����A�@��.��*�����if�o�΃��5E"��9!�91 ���H��	LgKb���'(�?���ɞ$N n׼�S5�*�SHR����^*K��fB7]�E�X�#�ĉg�St��
6�,�E�b����Ș�����g)n�lhdH&���.�h�K�m�H�J�eM����y���CjTw��w:�}�z�]
W��V(�p�x�#�o����҆�m�, p F��z�CrɌ����C���]4Lb
c!��XS \j�R����i�uɊ�V�5�X(���|88�f�Q�[�9ص���~q����j���4����  �j�A|朾ƚBc�F� =0� "Ƌ�N,��='��f,�YqM�f��C�>r�P���5Tֈa՛	~O�N���ٽy��Kja�#�}03%"��|�+!�LKn({o6x�OZ��q�á�"����и���T�,N��.�JbcC��'����Y�S1�Lh�;�xGʵ/�G��[�#�b.aȓ$�[?h:@�h�����;yS�N�]
���1�P�ᵴ�V��`��it�9h��$�F�2)�T�V��L���`��-QuS*>���⮹$Ѳ��f< �\��uWe[�9j�q����؝.�!�i:û(={�u��X^5�g�� ����,v\���S0)�so7Z�X#G��B�*��0��G`�$Y,C�ѽ�z�U%��`#�����ډuE�C#�#rP�3���1�@�j:$�U/���jdC��������DE鋃�\M��-T+(B-����MwFq�>~� (��S���i�U�N��(���Fs}͵��>�*9��)Wf��^Dp�WfF/�|+��ʧ��=\���
 E�`�AQ�ȵQ�,A��ڛn�)��OZ��,��W�&�����"����a�g����w�`�^��S�0�����Mg���8��w�=��{��b���o+��\��4�
��t|p����D_�r��D�=�N2�bgPdc�R�U�/V�׹�鸦��]qy�NZ����[z�����0�i�=3h�˒��.�jؔ�ݓ�"�
�/'f�ƴnz@�{Q���	�"�����!
�OO{��{8*U�LV��x��	�~8>H�]n��k�|���u�w�n�Y�	�Ǫ��� �X��APcJ������i���iPl�Y<�0a\�����g�� MUsJ/75M�����y+5��+<t<* V8��[t��޲��~�́>�\)��k��V)��f�U�\*q"�Fio�m�u㣂�Ei8����e��P}�)`��u��
��r�/�c{#��f-�<�}_HA'��Y��>ڷr��q��½�t�}R��2"t�  ��3�QL�@�a	��ۼ7X�F�A(B��0�1uʈ�~�x@0���q��w:��W�Y���
�̖�z+�8���Ɲ����e.���Ñ��2gj*�Ļn�m�Q_m�o4*	����)l��C���وEiT��V�؄��U���^@2� %����\����-�dg�O� �:L��D_��˞��ε6����L��1�ܱJf:���0�����59�w�"t'�(}h�3�Pܺ�1L�L"�dLj�#޿U3R�/ݝ�Ճ+�k�-V�� �f�eu��OM3E��zDb��λ�8%,f���G~lT ?eV:���%��)%	Dy�t��8}�Uǅ*��HO^������3W�a�N&i��n �ܪ��7�#c���d��A�[��Zۦ���#�O@��|�>Y�f�����i��Lp�4W�3�E��,�{jӞA$b���K�zϬ��ե\|�Ѣ	ZxXbqZ~5v�
���/-z�;��5@�J�H׀k9gDK(D�l�5�����G�8�Tq?~F[�����v���P����d�T_�v��Y}A�7�����:��f�>ej��XT�O8PY	�ws��֊��:�֫tY�����r#D0��-D�h0�k���,�#�]Wu��;�Gl���$n�j��1�.��ܻi.B�R�[ڂ�ke=��U�����@����	_�o���4	�ڝ8�����7֓տp�0b�7�NH�����sv��g]vj�^�M�1@�C�_	�R�;�Z{�r�W؂��k=K����9Z��*k��.%�9]�ي�#��b���m�|nT�ler�7W�:�t��+�X�dy0������9_P�<L���]t&wkF]�M��9�p��,Q�"0'W�^�B�����Em%zb�u=���0��CL�ǻ�b�Iَ]7��c�ݹ����� �d۲y�es�,�Z�5��h'�rZ���K��e���7Em22ލ�0Lx��#�'+l�����i;��Z��vI��~Tn��Ɇl&��2+��2��u��|�i�\i4�f�+��AT������W@�r��3�|[Uuv5'��T�ٽ|�H��n��\�	ܔ���%��
��bOF�����!^!�t�7	U,-��3�O!�튧�F�6�5m�ss%)�Z�7pn����C:qx-��t�2�nЖr������e�
����B۔/.�jQ1i�Qq�"���6�Ĩk��{�[�{ap���ښ(��hgr��)3��=�]��3�hpR81��
;S�v�t��
� �nP\FG�Qk�`-^ƪ������@���x��j𽣻"�%����
Y +�3l�Z�M�m�r<Kn@��Ʀ�\����E��[���6NP�+l�E�e�F�Y�e�n�A;�W�ա�:��c8����.�I�۝
IiX�=�]sfmCSRM�,�:�:���L4f�����.��N�����}���`�>`��(��vƪR,E]�W����	*�,�����BBK��r�)U�-�DK!�-D�3$�0Т�MB�8U����D����ĕ�A&RUJbDK�uJL(%-Z������1(�R*B�:�(�q%��'T�ցdRI%X�1&J�4���h�d'TE1*�B4��F�':u
�$B�-@�A;J����r�Tb\�Z *QAfq��I�	�%EF�8�%43��BB�4�bP�#��E�0��E@  �0"�$Wޡt�iV6.���[���3-<k����K��:7��i��Ɔ�$C�&PSi�����"|]ɽt�pI�S��< xI0�~;�
���P��M�����0�����W��$��Sxw봐�I�]�B�������#� �����A;�����Ʌ�O߽�o��aw���rNҠu
����s��<�����S���y�9ߨ~��}\�@ G�|F���2�|����#�`������{O	�!'?Sz=�S�;J�~ ro�N?.�O��v�ې>$�p^N�ra�o�ʸ�>�%��A}���	��U{m�A����L���������m�0�� ���{Bpx�����s�q>��';N���~q�&oN��I�q��_i��� H�Eߟ}��������?~�qΝ�e�r������OEmɅ�vS�aw���ݷ�ra|�;�"o����?7�Z`	�a
�+���$A{▔�i����o���>�"�#��<�߶�P>����i��'�C�iP�697����w���}}�񾸟�����NҦ��>pxWDޏ)�*|�{���@}E�������w�>;�}�90�o�������z��
aC�iɽ!'>���aq��������TE_���_��H}Cȝ�~���w�r��������&��1�\���tb~8������d�raw��}�$®�<A�<&�����9�!��i;N��?�����G|���z����}�����]��M>�m�0��ݻ�F$)'~� �۴���c�@�۽G&�Bz�r$E`���Ah!�6��s��4�3���{�FK���h
�@D�H���$}pH|O�r�����s����¨|q'���<&���Ǆ����NC�N��y�HyM*~n���DA!#�Vtz�'4_�g�ccR�Y�_T�-�חJ�0o(*e!����<5/�z�p4)�������t��|"\]�FqxnЉi=in�5Ph� �t��ݼ"��u��V�.��Y����O�U���RU����UPx1_PS�$�+�;I�7�1�<&@��x@����5�w�?]�x�x���I�!8=R�q �C}u�Dw{t���W��"#|F�qc��Z8H
�L��m
�@`�@�+Kɜ"SIK�eg�+�Wi'[~ש�*�yu K�
hm�)�u^�т8[<��3�S�iʡ�'DH�b�m$�ƾ�V���f�=ƥF@t/���(]��,pќe��;���wY@P�HU��[��Xu�=r�!�ǇզE�U
�J
 	ZH�
.2+��L�XC*.xLE\�Ԫ�f�9��<�!�rUu�7��ԧ��EE��0}�o�Vzhi��?cS
n��L����n�@ͳD��Ъ�C������(����ef9�(���<�av���q���z^��y�ig�ֻT�yR-zunh�/�hE�0��&Q���ޅN�5T�F�tNG�e������N��f�*�0��ȵ$�4߃�Xi�G/��|�ٽ��0�b�$�����x��,�l���5��I�<d��NMk����3�R�@�n�V#�&�5ɩSܞo���>R�9H䮖��F���ny=��K>��x��>1�r��ڃ����_a6k�_t�䖛�:1ʏH�כ�i�t���Wo��=R��O�<�i���u���1����2U��p��=,�~��52�>��ڠO���Rny�R{��O�:��5��px��K�:��ӷ��ߏ�v�!�Q��gb�s��1��7^U�_�^� �WQM̮B��+�����Ý1Nʜ��SlT��ˈ��;Vg�"�	��mf%��<I&k��v�du �����5�5�S����L���-�}�vP�[���Z�2&����7�7l8/Ro[�k\;�c�<��ٮR�+�ó�������eV�f�I�u�J�.�huC�I��z�!t�cTi���!p�*��̎�8|�n9l��x�=I�
/F�䉸d�W�WO��YTm
^�����H�1��6�iOgc�X�_^Ӏ��MTŤ�0�
2"���WK�)%��v)���t�ћRm'A�l�VV�r���O����n?r�����r��F��%�OVת�&q쑾YyؐO+�6�Ԩ�.5E`y�[�7�lSy�+㈽�S�iBmv��S�U�����.[�:�e+f��s agfn2'6�����)��ȡ�]�k��2A0�Z��2�V����%%�y����>�Nv��ս�޴��jxc�W�Y�+c��+�����cv*je�m�lN#P�]oe-�ry�Y��],��q�o��������\��G6�+U�0N䱤i\�'V����F����
>��9���0��)���ɡ8�d��j\��G�H}��!����L����M+.&q�����ʶ 51�X�)S�a;�c/�r�1��ge�p��X�CS����gu�T��ݔ�P���`��xohO��#o��ˍF%�QZ��Akp��!V_��rz�[_�X�`lD��qw�4��	% ���g=���D�t��8MjJ ��#���v�\i��JT��6�:C(�t��<��;�5�4�C&�rDO��ת^������y{=�ks����m��|��>�sh.ہ\���5M0c��9a�K�{��1�E��{�윯osVv&y��r��J�m
��#����)[��Ă���ϟ'$��QǇ�5NWg��(S鹫���%���qt:q5�O[C�N>�8���	���f��x
�r[&�M��4�S�j4˰��Y�L�{M�i�%�����O_��y���u����w;;8�'A���¹w5/p��bJhպyT ���-�}s�Lo^Jn�HU��W0�&���㓮�ˑu�x񛏏�j,ϖ݅gjj2�J��[.Hb�Y��-�ޣ@���-��y�I,r�N�0��6���� i\�El��I� ف�J<�[�۫9�T����N+�v��ܥ7.8��|��������}WG���D^�V#V��E�On�eʿ7�uǰ��Nc`A얝A��:��X��x�޵^2V9t>\,.Աܚk��5�ƴ��mw8��]�
!A��{�z�tҮZ�U�lY/�ΘR�4�*�;��p��\��)�M�<��C/��5A�FK�V�N�rO(S.�"��7��T�TWڵ�}6������'�$��ٟ�nb�:Ό{Yщ8�'�]����I�Kl�|�Ƿ�<V���/	V�3*m�B`)^�z5^��z���/��䧱A�[�}]��WEI���u���v�{�@���Iyn`%�O���w)'Gc��U|�rN�S�Zg��+��Nxj
ٷ�P�>|���Y�}���Y�$_�nS���P��t��Y��D����&�^+���L�\{�K��ʗ�Y,�)�6�R���Zř�[��灜�ڼ''��o�i��p���W�5�]��t��t������b��կ��wA�SG\Ȧ%�̪��z�o=攦pǻ)LQQ+��Q�v��ݕ*�PUmw&r\nw;A�
7!��F��;u�dSM�.Nt8�S{S����kҡD��{�'I���Ф��+E�Эv�HS��zD>}��s|�E7����]r�9�PkV[�>s�B8������t>	��d�/����.�;�AڛRV��.���ָ����,#)�W]mwm���#�t��'7؜�}&f��`�Z6�
5B]���uN�{���횳	z0�=��e	�kH�:���h���+ն{��]m+�t5/\O�J~B��[
�	�O����G���n��Y�9��fyY�'�Ε�mg�����f��ij��̓�%��9��/�Ϥ��T�&��+�+��G~ɫ�:W� u�}�Vߧ+�9�y�5L�g�1׽�	�G�#qN6�ᬹ�(-�����ʑʴ��ϲy�+��T��u'���Y�N�°�8��Ko�5i@�Z/ٞ#��#QVj�]�M�7HG8���[a`����\�J��dui�^	����)�K�$�u���o�f��F*�����9�U܏��ꪫ�ۻ͌>�n�<J®FR�yTr�()����^*K�bٷ2���U�y�t}���0��v5���/n.���'ꃱ���8u�ZB;�U��֓އ�L<0
�͖�j�-��qW��>g��أ�r�ܟ�$z��u�)�꼀���z��p���0��;yH���|3=H���6O-J�d��چ�]92�]-yg)�ܧ����M]�=�=�L�
Y1AJX��)R��S�J���n���c�9U}+è�g�`�y��;�ly���4[����o��{>�
���k`x3u�x(>�t�k�1 "-b�+V��!&�2�ػ��u�b����d�*����}+�[�Y�@.�0m�r���sl�Ś��J�X��<]ӵu�5Y|B�qp�GEV4�Q���nk�!��,ʴʼ�**�.�5Lt�8�����%�A�K�.�GzBU�e=�SE`r�v�6��(s9��v��oh�B��	�<(�u�Ϋ��ꊶ!��I����0��^n_U�N
MGt��>�XP���i��-�y#4bټ�i Yj��Ǖ�wq��2P����qC�!F��S��"T냶�S������?7z�¼����+!�����TU.=Rt�L�fJa���8s��L�Ո�%�58���d9\K�+N�R�{�=��4w���Z"B�,���a��a%���;�aG",c�f�(��]�Iy�%$��r.�:�aȗ}����W9Э7��{�؅��(�!�Ԝ`�Z�*mEIgRl��i��u"<k?z�Xqz���5�ĕ�����"���X#**�����%6C|q1_*���}Or�����]z1.}"��S!�A�8N�=��.;2�Q�ԣ<Ȅ�w<z�su s��.��B��$�`#\0Q9��qb��O�󚸵R�iX��nu��к2�%X+�/��L�#c�����at̑��{�.����qI"W#�B���I
/d�
��E�Er��J����]*􃜾B�_=��d�gxjڜkB��s�S:�~ϑ��v�m]B�Ⱥ�w{ ���d]W�'�i�2��9��{ʤ��! �b˺[�m.��ݬת��vaN��}b�kw*�T��4�8q��6�>�hwo�
�-]:F���ڗJ�k����ؤx㗧V�կ�)ZpjҼ�^���M2��V�3m��K�)K<��*�H��
�nmz=��dx}�� � �ufĩ3�2�3PZl��U;+)aDQ�*a��ԫhD���iZD�ԖrL�(�P��,NҫE0�p�9�N��.�EZڬڡ�Q�VIҨ�"��XA&]U���KY���Y�f�L*�SK�A�f�J+C*���"1%3(�D%TZ�+&d�I�&��ZjI�"��KMA(⵲(�s�\�R���.�S�����Z��ZfH�mP���$9��Ve'T���%I	�� ?O�{��Q�j,�_f)�.�'��L��˕ιZ�lQV�n��U8̽n�_��U�}۱��xo���xv?��"���{#=�O<�k�=����s���X�k�80����u=c�]�CO|�g٫�����G2��ԇ�����<���2k����W�;~z\��J�n����3����ք�/8I�˓/��V�^�[���޿����:����/xO4�Uv&��o8�b:�s�9��ލ�M����N�j4�1	��D��v���/��#w���m)�u9�PT(1Yr'zw�ݫA����j��]<3W��w~�0����Q��M{5+���W���?��A�"����t"U�9��2�7���@"Y%�?1�p����؇$ðe����Ԧ����X&(3�.���VQQ�Q���>����]���Tߴ[�-�ޅ?F�74��M^�/c��0*oN�j�l.geD�7�ݖ	=�����(&��LÛ����-�\f�����z�$�K�ٕ�j�:,��TB�ә�R~�9��OzU�=➷��L�v�a�h����S�{���~>;-�ݙZ�G�	yC�B3\s��u���uhy�.]Z�<���2pq���1���SND�;��37��Z�˂��t�l�g��I#����3�-[QٴJ���0�W�jкS�N�>���:��3띏�l(]�<����ގbi
9�EV+����H5}R�-���ʐ[�go,�.�rҝ@��jޥC;jgr�R���ؒ��}�@�Z�6+Ë�=��d5�&��^U��a �y�?z��-�.z�͘��"w����tc��7º�[
p�uo%f�s#z����M.��i���1X�e"�hv�����I�u�ﻖ󸷙c\�3G���H�9j�������ż�ı�̫GoҳFmI����3�=򈦧�O.R�J���,
��4�&��k)�\�_�&���[T(�8�ae�v����u8�R=3��55mu�ީՆ�tó7�ӓ��ױ��|˘����L�W�vN�Ko(Q����`쨓�W]
r�h۰�Z�6ХF���,�!�e֬�Z�˰��{W[��D��A��;�ꉱ�V��q��#ѫ�yʖ�k��m���UU}�^�Z��^�*`ڒ�q�f�V^Lf�U\.�v��B�'�x���WP�×A�?v��}[r�ڇً��]�g���^b��4	��WU��r�}�0�e}cئ�1���M�TW��	)����֫�Ӯ8rL��q���K���s5�ޠS��l�ޗt��r
6�ͮqؗ^n�V&UE���o�ؓb�e�t���/{�V�}aqG�h�S\���x��׼��u+(�r3��s���o��kh��GLup�l)s*��ص����L&��׽���7�M�Qd᫽o&��A��1fb��\��f�u��tiEy�a:�j7RV�%V`�JMK9��&��ָz(=[Jd�&�!
����F�~�����魻�i�;���迶8�@��5��-�NRqz�������w��ʘ�u�¡�E�Ɣp�Ux��c·��}�z�'G=�n�&�o^_9�3ҶE:��[6zj��Z��9�}�z+��_e)�#�C�㢫��m�FnV��c�0��Yw��Q�H�{�<��J�Y�W8��{`�yg�
�	���nC����廤�k�����3+ދ+Q���՞|�k/���{5�_=��i5f1օ~]�o&�e)W��^�V�ؓ%'���B�{��zuK�+�=@+�xa�ja���C��*�?n�ջA��lq��&����/��(��e*z�\�
�n�Yӛ���EL���:�R�Q�����l"t���+FgFu���~�����Ym7�C��4�F�l:�v�)�r+���	W|������r;�6�����kN��(����ֆ��R��N[�aXPc"����闑����Ԏs��H�50��	x�?�*���!������ϝMMC�&ه-֨=��a{v��Oz�Z��S7�\�V󣣞䯖��RK.�|�?_iU�+�VQZs�����O^ߣ����u{���>O��m��a������s��kyw4�۱�(�zKi警Q�E~�a�*/y�#Ag#^唓͹k(iE3 t|�>��+�ΜB�g}g��70K�ز.���`�57�	-_�CY�nL�3ݒ�ۺ$*{QÝ��K�w�^I���	�����\���g��э{�U}��U[���g�5���{�Dv{�>Z��y�)n6V�^u�\̪m�C��"�L6g-�*�QV�f�쥥ɞ��G�n������?N!px��-3���Eޭש�雥��n1e�S�5���ӌqY�=���%����deҾ�J��);s?��\�|��Q��B6���@iW��c�Hj��,U�|��32��~߄�Ծ�V�i
-�6�D����qm��ɑ�!=O���L8���u5Qz��L�Wo�n5tn����#��;���}ly�4���1����������g���/&A"yl�����4���!)��U�8�z��;��7���k�=�K',g���<5᭫W�v�P&W��5wVȐ�vr��#�ꕾ�~�1���:Q1��?nt�{� ��'qZM�.-E���2T�sW�A��Lo���83���������kW�>N
~���9tNe{��Ɵ=��.++�W��@��m*�\D�y������!���mc���~^e�yNu[�n7����ڦ�*�4�LI�r��|O��V��K}`�5�P|uy�͘�7T�6q�������K�<�+�w6�QC��g5�Ĺ�oTm��h��6�uv���|��F���9�v�X�9F��d5fv�������O2�����Z��^�7� `��W�J��,M�;R�T�
�u�l4n�"�M�4��鶀��3ӎ��$(oP����>����N�\�ﻠ��B{��T����T@��B�n^Y����%m)/)*��Ew7uM�7��R�^��+�n*���P4�#��Ly���}xj����7��^(\7�+�N�;=��efp�������s\�9Z<~r�mCR�d�*��K��I�1*��Ş�x
GfԴ�~�J�6xF�`~�&~u��:·�}���u�)'�{kk��w�i����oכ���{£Cϝ������Nb�}1�0{ ب�s[e��{N�y˓Q�OdlΣڞ�($U����tǖ磫�q���ڪ��.��/!N>�Lܖ�n��V��;Fk� ��_�'�1�߹���@O	��6M+��p���^&�wG���+�n���'8���{Y�?��>������y�����4�����d*�*G�����,㛽���3��'��q���o=^<��#�󮍕$g7�ߪ���e�A��o�G��gt������V����WJO�P����[�H��K����a<�J�of�c ���Kl���<|�.2������\�N�o-
;p�'n�Z��M�N�?ZM�=*LdVYg�r�GF��kB�M�ӵ�k��SqR��������.ƞ���s�f���kŽQЯ���{k޶��9��*f/K��K}�9�}�C���N�۴��&�yv�� ����/�������P�}�j�\mX�L;�>Y5�՗�s9�\Xk�,]�/���9h_(�*G�b<4�A��d��f�详�u��b姣k4��������)�Le�ꔴ����a.��vC&����d��N<���+7�4xmi��i�sڿ��<WY���k�h�xd5N�r�͛V�y��ku�]�^P�o!&�oܕ�\x�Ї�6�p9�3E*DM�r�P]rh�7��ҩ:�[�0I�����Sx���}9�P֊��sO6�����e͕
��4_T��a�/�9s��)�[�9&���u\l����KB(�YU�!�X�5K�n�%u�ic�l�{�Բ����ܵ�v�{$�V��f�$^۵��z�R����'1k��C�M)W�c�[QV_�e�LF��]�Q�il��j�X���6弝��j쾬#S�[���MT}�_NR>	"���oa�7��.N���.���X��٣Q�|��=��9}�4!-lU�����_g^��Ф�q��9��q&m^C��Ƭ�P[�it�2p���d�����ŗ.�r*nǳ��5��fNB�k��A��v��@ykau^Ԥ֨`�e욟N�1��σ�QLA�ΧV��Ϡϕ�Ԗ����)�jB[�p�yBɦB,L<���nR����1�h3r�+���w&w`��Suf�/b�F�%�>����y�1r�!ت<�!)$�Z�5���-�}aԸt��H��)��hMP��mI������?�N�rzy�%nf�o`i&q3���Chܢ\��"����2i������^r��B7'=����t����OV�2��a���A�xW�T�Y�eE^�]p؎M��w�E+�=l��K��Q����V��ZV^��Ww��� 
e�Mg*�PB(���X������u��R�3L�B�A�	2C,٤�Aj�bs���e'*��0��+:"J'
���.�ʠ�"Ҩ�C�Q�ʂ4:����1R�N�Qe�VI!�RE�"����3�eʈ���ه4�YE��R�,�\�):ATD�iP]R�I�Y�E[Z��
*�Ҕ(��L5�j�"�$$�d��Ȣ������H\9��G�~��~��t�앢�<�����*-�}D�	Ӈ���t�J�ۢ�|�R�B���}�}UI�$�j�漤�h��޳�w}��\뽊J�/�yIA�^�k��z��9�˞��,	79���Ԙ�T�/UI�8��G�w	ݩ1��w���x��!�7[��RL-}�{���e��VPt�����n-0Q��C�Z��%Ꙏ2��:�wbc���ъ�\lU&����{|�I���i�F{�ݷ��*l����u _֮]��+z�������|'�]=��-50�;��)(	vX�ѽ�hS{�⫐���L��9s�)�Q���2J���7��z�1���G!Y�E�Bج��1��'����5�t^^}����f�@/�K;}ZB~~m�;gkS���ƔT��UI��E6�u�u��K��ӯDk��UU}UU��O�Vb��+^��N��\�s�Y�_:Y/p����_Eh=pn�t�6�g\9?b3A���ޭ�<rS*���0Q�Rf��;f)��T�86���8�N#O����W����6=xp�W1J�r*hG���ש�	����7H�kr9V0�HѶ6{з����M�/R�Oi�Y���֛��=CT� �}�����fyC�"��V�ϝi����I5��C�r�V.��+:�_Of��6]���Ŧ����Ό�RɚV߻�&Y�������|��˵M�@U�>����]�I�����k܂�A�����RVw)��}8�, t�6؊�rt$����f�W]xi�~��GK��%�Wթ�=�R��&��W(�W3��t��S#꽖͕"�F��]�����ݵ��su���u�B�D�T�*��a�.���jOz�a���N��'�!���d�����<��d�I��Z��d�Va�{�5}�����/��=}A̍N�tr���9����V9pqdj���)��'�ь�������Z�#z�TYN!no7"xU�!VԔ�mO^�aSn���^H.P�L}��ٍ�'�^�M~�}�_^�_B<���C����Qo��^��s��6���H{Iuo]Ym���^���]&����9Pi}R�Sԫ�~�϶F�Z��m�p&on4����D�\z�N��)d.g��:�7G��z���ث��J�\dn]Ց
(��Yoȡ��C6�3��Л�eD������u|�zG�ˑ3T`^3r��C��ج�f�O���1��ݫMob�/M��6��l�5s6[|��i�x˾U����S��m
���)�Ǒ�[����3�ۆ<7�uoR�,��thѫZk�"�{��{�B�E�O^w�<����g����j.(�M���T5X�%��c�Ժzp�c��l��"��������[f����w�;�+�V�5����U��P&g*_V���b�N`^���%�$3n{���qx��Hq�[�T<�=F��Ӆ/�(m�I�p$
ݭeܣ�T�v�Դ�Y��Ċ @���r��輼�Ykd� 5���n-��K�!������zS���{&4�݋�2n%��� �St�q��w�U��4�'ʜ���G�\�f.Lz&A�Sn��1iL7�Q���J���k���*��3�\����c54��n�K{�U��y>��z�-��Q�'�;Z���!GԦ���NnY��L=�۳���w���{���OV�����c����]��!7�~�����~X}:�>ŶG�p'[3�Y}5{����F�P!���CRd�L��\�jI�A�hΧ}"��e.�{1�Ӷ+{]
�coe�s[��&�.sn�kkv�U΋udMVZ�ʍ�n�ظ���'��6ߌ��v�Ҙp�&[���Y:�p��t35�X�Ey[�"G��RX`�Iù�Il��}���%���I����o?�������ɒOV�L��I�k��l�Z>����aƽa��'����}��ǟ4�.��-`F����s���b��O�K!�9siś&�L��/ݚRo�S+���K�Y�F��p�$_3"�㙵����p|-v
��-:33ާ�%��<�mmL7`�d�z~�B���JP����܇�$߭��1�G-<�h�r�)�0�\=��K1g �-KLvt#�ԧ엮����Z�A-��/v>�4ڕ"�\¬�4�r��3}�5{u=��Ҷ7EP8�>�n5���xL�0�Y�)rB�6`�㞡b�GF�9s;4J9�&h%�*W=u�F�P�����ՌM�;C6�tN�.�ӎ-�m��V�H��+��r�{����NL9�~���꧉)��b�<?}���)�ޑ�wb��y��ym.)�ល��m_�nmc�ߕiy�t}Hv.��I�9ɪ�޹��;?c`��͠Η̚Ӑ��u�|���.�i��B�?A�s$ι��~�=]�=ⶫ՞��t�*)��UxTo�#�=W��^�+Q����P�)�)��R3��V���jҍ˦Ul�Յ��%����s���{��QL�I�u�Z"���׽�B��Yo�ʹ�#hfŰ��ۍ]mr��!Nr�ݓ�޶؋x�{u�j�7 m^��3μ���q�e��b���>�i�{B�]�:O�)*gWC^@r5$��.��ya���NhX-r��a� \)��rۜ�G�}}sKV�`z.�V�n$~
G^���@J�.���s��V�q�5�;P�q;�îບ��f�ۥ�����L��4��A���9�v8�tܝ/P����i�]B�b��K-Sy��kWv��:�.bw���M� �7W�75��:Mֽ1�ޮ��#5)M��;�5ҏ��W�c!�{��w�^���Ž��Rì�����:-y͜�PV�X��+�T}�Qm[�g)ؑ{���M'7.l��FN����b��*��Ν�u}�wi{�=��������v��ݧ�������Η)�X��{���)�x���W�凪�9��5��svZ;�l���*�pճGZ���!�Cy��sGg{��躔�&�2�ysﻣ�D7���F�h�J�[��p�vs%tB:�i��j2�5S�4k,���zBc%Ʋ+&1��ҥ���!ۮy|��w-�|���&7��Z�p��"~�B(�Y=�1�5}�g,kW��dZR�s���Cg��h��W׏=�Z�k�^[6�Ӊ`qP\��\�Uہg����[5��O�X�~��P�ֹ�y��!�>�S��F�q�};���� �%�/+��^g��R�|2���o3؂�"���R?[�g��D�Z���眡O�ߩ
���R���3��F�qm(&����޲(^c��[}�m6��A\�'�غ�������a�;+24����p�y���V��ewu���N3�O��UW�Z��������f�c>���fZ�3�R^s�Kڥ��^_z�ڑ{**d�]����o�hպ�؞9�\�[?^��]f<U�jp��٧��Y�Fm`J��a��S;b��׻ݚf��\��f�(��Xʕ�.�b����i�Z���&�l��+|�\`�k�4ǻ�S�r��h��,崖QR��u��:�>��˧+�p���9��Z?F\�%�09�_��|��r؟�
�2a9���`�d�fj���u�iW�����=0f�^M���=���\�5�%4��ʃ]tĥ��ạ�G�����L��S;A7�,6�d�{Nn�JD'}�s�{q�uk��,8�PkE�z�+�m��[�Q9)A@��dM��h��� �y-�^���#�r�]�n��-7�1W<��=O�9WMa��aծ�T_*�z�P�Y�e���;�"�fb�W�����=�sO,	��fԡ�wh��)���k԰B�cI.�wOn���X�a�pK��l#��`�4 �@U���[�^.���ɍ��d��  $�λ�ڒ��d�Z�J�z�l���5w,.�v�0�KX�X��Rhq6�
��o��-�f���B�en5�ғ�b%q�yo��+s��b�I�n3���q���Wy�1R� b���rV�u�"+/Oq+
�ԃy�i�G0���D/�%E��H�8C���܍�~��8^�j�V�=Wgu����U�UǨ�r�kNEu{��T�� ��E�����w]Ꚓ�f�޺.f"���dV��W��.����̎QU�.�9��&�M�Yr���K�TEJy����IPr:f%f�]w�DQ�"����I]���[]fp����*�F(gNt��4C;���a�9W�mQ� ���Ԯ���&a�]n'K_h��0�g�*"�41wc5u��f�X�y������+)R|�]�2Ļ�X!��e@��{�>��>���1J��>���|o*L��[��>>�k[b��V���@&,��ӛ6Q���;e {�l�jMvvI�^jeS�X�D�U��v�4䗛Ⱦ��|Y,v&/,�5wHi�Y�γJ�b�;�vd��<��̲�WQ�a���s��e��K�� k��s3��}�ˬAX���)a����++{k�s<9�v4|�nZc��۷N�s��T��_PB�U��*��Ի��/tq��(2�����^k�ͼ�|%�u�Wmu�\����D�-���0�>�%Ԭ:�=>L�ŖUPUghT�D��ir$�8�TQ����B9�5)P0�`�*� ��)"�]P�\#T��Z��R.U(�*�a2�(�%�a�rQkR"�B�-��R�9�#�)a�#L�$-��UZ�$]B��L@�QsKi�fBU�Ad�r�J�:vr͗9*�g-Xs��	$�Dr
Q
��&WNY	��P�ʋ�t��fE�E�9Ȉ�Qt�,���"Ԡ�QÅQQ�uH���r�R.R����~چL��FK���L��`Y�J��.�c��L�%�-��=O���\�9��}����Q�z��[�y��\4���i�њf����|{1����ǌ�Φ=�*KR�#X���1��f"ԛ��\��=�]'Αzk3�3ؤz)�m�_�8չ���scO��j�]a+i'���%^v�yr4����W��z�A�t�C�����,�K]蘺D=��|���If��w(�,3��O��u�B��>ҏ]��c�SN�xM'��?nS3O�__Q��=��:������m%3*�js1��|�r��w[~>'� ���~�Mj�T�/�?��� �Vj��K#j	��5�����=��L���r���N.�횾H{���]�KsVmY8՞z��Q����V�Zċu�L�H\�KŜ/���UU}�ť���t�U���GH�c��ʞ3�CYF������)S��8ƹO~t�ǯ�)����pd.�D[Ik��BS���OA�܍W�r��G��xg@:�NER�kPn������S{k���'E�z���烵X���AKp�!A���{��nR�E9Z���M�gP;L���!���<W�
*���|��fb�3�M1����t?[=��~�����iR�����s=�+}�'{h��3�q��m���{�(9�5D^�w]�:0����N��jzr����{�f�СG����-}:�Y�{vt�l�؎����*F�Eg^vf�[�s4�`n��WpY�����Nj�&���h�E���Ί^�+h�Yu�}U�}C�%Oz��3��~��~�p�W<��J`�{=�^>Y��o����>Ϛ�//5Ζx�Ӟ���k�P���E�EO\��D���5��91;c!���V�*��#���Q��t���&N�n�˓*
�z8W9=fy�.��^OP��}�b�J<�rk��.��:��o����J�q�C{1�J/{g����l��]�1v��U	=���-ZT7K���L����ƚK�X5U����)n9�����Z�SY��=�n�D�;t����L�b�iU��~�6�	�����ɩÄ|���zJ�;F�UĻ{lY=am�k���^��ٗ[K�7�"�KT��`#�C����n%ϥa�m��=��b��c�N�{�" Z���5�����4r�3>�6���s���|�N��`��M2�j�oc%�|�h��챾2��g�
[Zh]�s{ci�O���"ewL���OqT�W�[-=�;s�{�0gt�|T�y�DvY�-a��I���rX_$��*s�wΫE�?7[x��GѠ��w�v�A`<�d�+o��u�K�}�R�p�>m[bF:���
���6��Ӏ��xg���U�yh|C�εz��N�~�q�㳎?W�'�4vl������D0&Z�b�d��3��Z2].]�̽ʇ])Qk�A}�rj�<�0���9l�5����	���-��RT���2oj1;���=5n�%�U~���>���\�įE��B���;��E� �lJ_��MU	���ع���~��g�w�ê����Rlh�oný�"�d�u��휀P+��r~�:�����^{Ҝ�ү�W#��������}](�os=<�c��d����aS�4�i1�z�q3O;�s�lZyw0�Oڔ�h�����S��=��c<]�8�4��~�t� �iJ?}��2��C]3>�u��uEP8�6/e{gm���G�w2Ό�re۫]�Uj�b��U-��q�b��#b�K]蘺JC�\�z�ܫm��@�����_N�P�~�'�M#�-?����[D��]��Ps	W����=~q��J�F��2���\#�;ik��r�+/s{����n�N����o�z��������O�h,0*�Œ�Ԡ�no5$�.^Vw)�J4]o]��##��QĂ{���L+�Y�\f��UMm�I��,<�i��`�]2HM6kQ��O���[,�"��R��O_4�qӤ�]?ɮ0�B��+[��z����.5쟲6�y��P:�8%�[ٺz���vR9fF=Q�r�{��%q� �Uat��8ͣ�q�*����6��G-uZ�Q�ԣ)
ͿUP1�\��ϕ)��҅�l��RX�^�a��3����[SC�*3��У�/Ԉ��d��5�F��+4�W�ˢ�prWsV݁�&r��#Z��h��c�VO�7��([�HWŴ�q9�umR���BB%nBj`�7Kblv����D	��w�=+"��"���c:4��Ή�!8��v�T#�2XhֳX�t��3��t��ʥ{6�4^en��Y��g���ݗ	D�IwY�;�T��ߓ��+-/��O=wSp��~��[~Nc�'��rp��)��{�Z{���9���|��F�����#�]�72���R���fvl�(�O6��F��'�^~������� ��}��Xz�>���ܛ�Z�ߓ���t�7�0/¼�aE��n6�=��rז�7nJ��Kط�Z�ٴ͛��0��l�ZەQp;��WD|c�����xn�z{ޛ,�&n�SQr��'LM�긶����
�)��L��\�s�X�R�?�����o��U�̧=fl�὘U���'��������ʆ��F��w�1��Anf�=u9�o{VhC�d�����靖����d�TR�z����Muz�Z���_�˅nbV�qÞƗ��ۇ��b����B��Z*�w+���OUU���f&,��}��q����Њ���gm������ĥ|���y���8JϔR��h�w���3�T4�?G��Õ�g:駇�U'��z!}OQKٽ8��Kc^�V�콰\���~��v�4�>�zq�CP��E2��b�|�o�M^�5�n��P�
*)x벉�%�V[���7ؤ�RB��Q0�r�ڿ�1��r��R6����^�.� �xO��]�]
}"R�\�;ܝi�zBO��ꪫL\�j��|�\�A�v�v�ͺ-m-�Os�x>�1�mp�����G��DY��/�.�CӬ������ˌ��4y��v@ޫS��7S�q��p�w�w]���i��I�Ĥ-����,\K�۞��J7'Z��F �i�-��S��=�"B�)ODY�X�~o��	��k�$^���\gS�#meNV�?b@OA��6)�|�AJ3Em�	��
�hJ�����h ��VT�s���#�۹c{ls3��U���M�}��-pjWe9l&�(�+��������8��k�����nG��^���N�ʵ艚���I\�ҭ�}Y����1K�B>VR,���Qo+��c�3�Kr�=˝�5���w�>��謶���/k���M6�:4����v��U.WS��M�L9���gb�-�����\��Gv6ӝ��	�3Z1Z�*�}j;��wns���?l�O/���z�DE� ��	�2�Ʊ6:t.[x��UwU����^�ׇCCW�~��hl��W�s3)p��U�X.����O^V�e�P%i��

b��V'�3�>~g=�}�Vi���zeyGC��SV��M_F69��'F�����U0/�-}�������R�ZzЗ�FT')Z<�9wθ��9>���+��������9�;�Iv���ί�6l��Լ�J�N�Յ�.֕�Ƿ��I]>��ea�Yvr��N)8��aN��X� ��ۈfV#��{p1é��Ȓx5@U#�%����N\����P��:��#n�n}�����R�ŷ/$�yXN�9�����
�s,�sq�5Zǵ�;_j)I���O|�b,�LϜ{�gǙx�6���^U�J��~�����R��ֵ�j�K,cm� ���tI,����FԵ�@}��]i]t',:���n�k�3u����7��J��ojވ���T����֘��x�!��]N�һML�%A�\��1h�������5�:3,�"��Z4s�%H]�#fZ]�ڹ�R��a�U]��5i\��Z��*�R�(���*���E��`���s��w�&x�[[]����e �f�]s���Y���Y�C���IȌ=��B�::�YVY��k���}��|���e䍻�Lv��A�_B۬�:�3���C����W�睹@[�bt�a�e6�bZ�P�'u���"R6�a��a�N���*(�[\�SmS���t��U�8[��Q���S�cvD,�L^5��i�{���#6��� b������(.FMM�D`�Q=/ ���M��t���k-�jR�#�b�ܧCt�<\ģY��+T������4fHoPr�i_�nH}�6R�Qܭ2�ٱR莓� ��V�V��=gA;���Қ���s�ث��g��i���,mc�%;����.֤S���".�Q*��Yl��d�%��k;{�I�I��%k(R�qg[r�m��s��[b픫v��W��Ŧݸ������c�u�A�&T]�ӹh�<2�����;�	�&�dP��_�A"�դ��4HȉL�+��f���) Ī��s����͑sRAH�����E+E*�SN�
��P4�P�!Y�L��(*C99ZPDXQ�DE$�j˅uP�Ge�uB"�AR��M%iU�DFJ���9Qr�$hZ%®%F�Vj!UUжX��a��Er"9E$*��Z����L�*�j���P�	r�*(,!	��B*".r$�QI�)"��AT*2.&�\*$���S/��~~��+��Y^�<�=�Ɠ���{P�ƚ��K�wEk���v��R�W9?�꯾��������M�hs�r���Ɂ�`�|!��cJv���#��t�r�9C�M<�L~�p�V;EV�����>�F��q�ڕ�����9	�T�u�4�Cj~��WV���S��f���t�aN��V���t��sc]��;��t7�5�@��*�x�V�ThB�q(�����W�=J�l�ͬA&Ƚ^WŇ6�N�-����*S���/,�7�������z�=�w��\~�)�g+�t����VJ�PlgzN9���F���J�?L�����,��o�5j�]$�`�u�^ZC�C��_SU�'����&�i�F�8@��dډZ��"!�>�	��ha�(�.;\n��,���qT� 宊���
ۼa�^pb����`�8��[9;�#V��Ӵ��w�n^�n���'�[�wh��9:oj�Ǯ�tb�BH?]\�p���|Ş�ꆷ����J�j��c��6��H��p�%)V~�xof4���<�H&��ݭj}9LQ� ��ruBL>;���Z��k��$K�\�s�B%�
�0�+Ꞑ~��*L����=w���Ŭ����i�Fw_=^H��ޝFm��=j�J�8�����tT� �~0T���:�)I��-e����8�<�r�)�M$�>���^V������dl!��7��ۗ�Xɓ�ܮz�ˈ��KR�����/��>�ؔ��DLK����@o3H�c�rm��csQRnn��i������п�f�k;5��t�r�mŪ�/67�޵sH��K^&���7=�<�禍������~1�>��+�g����v��)^�3����Ǘ�^*JXuz��e.� m��S�~�bst����f��֛aK��>�7ً���*"������3���M�ʽ�c�����L�'Ut�h0؞�p���ɺVs��E�6��N�EH�&��Y|�������u� ���[η�O�_�]�ۺ�y][��׸!��;m���7�Sf�L�5�n��P�;浄���W�h-������R�w�m���(m�q�O�]H2&n=u]�%d��T�	e�m��R�ʼe7�o2���=K'�IH����\�`'S-�=h���1�9�%f����i�|��=������X(��^�{>���L��aB��n�&��/���ރNܵ�YH-K��;vk@:�����f���4�K��蟷�iM\�53-����D�e�a;�g"/��IU�r�j�WM�T���HN˦ȱ�U� ��])��Og��F���8���먽��Ʊ���0���C���b�g�ݨ�����+F��vwyJ�>�9��ǚ��gn��h�k�׍=�Ĩe�V�5�5M?S�^�}V6�	��|f���t��ھQ�'^m��=�����&~n�%�]��n0�Vkd�#��1�g��q�S2q�5�kT��Y�p�ki�=�{&s��Y@
�2y�j9��N�}�1ϸ����ۺ�����B��$z!��aڏ:M�+��Z�,ߺZ�)C"ʺ���ҵ�NE����F���r��l�A�4�.�{�[��5=tה=�>�$�r8Z��;���=��>��2ڞ����n�J�[���ړKz\Y�y���LSΰn�j��7�4��6�j־f)�dr'{~��T�т�IJ]�b��CK�Sin�-V+�e�^s���Y#��q�/1Θ��7J�7mY}ϲ�[�␧��q:P��N �6�G˚��u�;ڤ�Lͻ���3���
�\��Wu�C:��")Iv;ez:<�����������~����J�����/4�߃�z>��;8�'x��z��'��Dz�Kέo�g:�ð\s��E�yk�G9���9)�m�ۼ0�^���ȝ�U�fo����߉!�D��7+#K^uu�d�FF�I̎Z#,�&���m�sz��^Ň�$�杷�����w���>���o�r��F�ܙ�tz�;�[��n']�)�a��vFؘ�{[�U���=�;�M�?mG�OW��.�����mB�o�������jߊ�F�F-��i_V�|��4��<m��f5��[.�;�r��&�R�l�������uрS�r��r��6��](']N�d�*�{�7��O�",.6������ϴR��!{؇�H�d��@���"o.`N���v�-������t���c�/�T�aS�F��Kr��;�b>}o���HR})�쨩F��d��V0ϖ1��$�s���3�N��eD�1��]eӜ*l���&��9Ћ���u��=�W;�2��xm�;�~^M6&qàT�yQ�n����������'��)����uV�+��=�4c��h�s�]o�������޹���te���2�8r�>����O�#�=ٴ+f.f���*�&�S���"��}s/�N�&tV���\��h��f��3�b�$ak)WL�p��D��sHX�jEؕ�}˧U=��l��������HA��m�S1ik~^��k�˙i&��kb���y�����ޝ�IN̯ރI�vj����R~��Kյ�T���'+��;���gռ��t�"��{|��8�O��k�Z9����={��M��C]��'Aog�:�525Bf�m�Žr����J2�m�@<6���mŊ����^I��xͧ�Q������SJӎ1�OZk�����_W���Q��uQ���Jyb紩�W?:14o�3M��8�
���w����io[�A��L�֞tiw=7`y��zϩU��@�(���b�|��	������rng9�kX�-�+!�X�zy)[�:�b��� M���`X>�ib����h�2���.�)(el��J�g�	�����6�*!zlďq��3u�9��V� �Zޝm^w0+<��fNZ���f��6��j?m��W�Mᾷ�Ɇ׋����bd�ņ����>��H�*圞jf*�/�#3��^`33����f@��:��n��>/���qM�|i��.�ŉ%�i`���yZ���<cI�;�t*g����w�<���:��י�S�c�Wo���Q�U'�6��+�����9v�LS��y#�A0�`'?p��F�8�`�^�*��_-�}�͌W<'co�Z�
��dy���<&�kڲX (��K��׆�(vX��;L�`���}�����NyՒYA���2�b�[[`#a�`�5��7a�a�pEn�Z�(3A�;MnF�J�c�Sgsԫg�
�:1Z�������$s�������QmnO�Y�Y��m;Ԯ�.���ir89Í(�U��ȝ��4˖�����-;�~�HIʽA�m�F�M2�aŹ؅C�ގ[��>���S�K���Z�b*{;9��Z���{�.�Q�tc_W�=��7
�z���b��w�-{����+�����e[h�������YC��h�U`o���t�Rٳg��Jny����@Ҫ���I��\z ܅Oz��
�5�}�+�=T�Z�`	S�����J?&���Uଫ:Z�����ƑBQU�el�~Y[E�*,�G4G2ة�f�w�p��$����FMn����"-.�l]�\���0tFu�:h���Adv�@�J^�4-Q��O,7D��!�����Qj�!�1� �w�k�0ϱ�ǖV9`D\2_i�J�l;3F�v�-K8�:�vX�����n���3
�DZj� ��t�`䦃7/N�;���#]S&ٖ٣w�3F'�v���MA]b�u����/��(b�ݯ,J���`M��F��,�qꡋk#":7׮�N ���X��$�1�)"�p��+��cx*r�,�0.��l�9	��y-�<��~��O�k3��N+�ӆ�7ֲ�p�Qb֪V��2_�÷n��,��#�QX�����0nj�2�����e��l�}�e�"�(�73���]�9�T����X�:��q�O.�Hjk��w4����ȩ�SB���"�Lr�or+<e.p�G�GB�+�l��MϞN�H�_8���ƙ��Nކu+�Bv�[ӵ�ق��Gm0yHx�2��q�+&�{�ٌ���١+�~q�[L�i�p�ڋ���[-�����ҭ�9����Ү��/�f���')�y&�۴�H���Ǥ��n�v��g]:� �_�]DǙFEy�+#�ܥz_wn��M�Cp����HsV�CǕ�+"����t-"[f��9�E�PsA�j�.��yԛ��8ۼ�kp��e-<i꠵{��zpˡ��˶P�d���ޏ�����tm�2(�'y�CP�H��͉9��p���2������Xw����Ұ�1�Q�i���,����i�7��^�G��P����!xԥOw��_J�i�p�7ɍ4�D���Ί��4+�a�XD�!A�����B��_t:5�#H�lE�R3�,펷 ��e����Z�jt�*��ռR0�F	V.�PW<�
P)�y��9�gj���`��(���ɗeNP��|�j�y?\�?�fˤ�VB�s�h�%"�D.d�(�˴8��JQQ�ir�V�U��jƄ�B
�0�
�E�J�]RT���Xp*�"�-ah�Q�H��(�D�A�$��ò�˕Ar��H(�*V�q*"
���41l��"�\�B*

����RHG*
aE��*e�M2���UfQ¨�aɑ2"��v�V��A�p��(*�(((U2
�&Vgׯw�9��k�ya�\�̉V���r�䔗s����nyL�չ��������淖Sa���[%�K�*��.RHc�sKM8���R��{�V�w���#�#�ּ�B��}^{!��v�)����������6��pz
G�ܸ�v��W+�l�ݬ��ǹ4�J�/}?\�D���X�l���7g=����<����r�i�Fз�Ga�����y»���+m�z�L��	YN�R.Ԝ.�y�R��g3���-��ދ�eA�Z���Z�u�x�� 6z��,���,�G�M
{[���r���Bo���R�����u�fAZ��pB�5�6�W�+�Xқz�]L��b/v�ZyLK7Ȣ���3��vW�&�VKӯ�����.��鲤9y�v�gO�9���W�A&4�,�t��b��'!�ZO����K���=V��{��n��K>��N���%O]k��-��^i��ox*��V+![��^��m�ر����������ُ$��t����-��Z�&v�kpyĕ���w���z����^�������uxk�W%L�2O��Ľ>?b�/�r�yܨ�sK�����FT'�IO�T�l�{nڑ���qN��Kx�.7^�h���
Q9��Q�t��NaK��z��V�^�?h�����ph���n���[q��r�J����3)�O��˥A�-2^TyQ(���ct@	Ӆ��X����ݮ��<�{ ���|Z��0�n^�q�z�Ɵg����t8�T�V�j��;=��?��8
{74r�������s�^�r��$�A���N�f���t^�)�����ː�V�\�OC��h8��nLa;�S?)K�%BU:�Ξ����xB���4XY�9��%�u^g�II=�z�W�����:�z�:��	H��7]���n�t_���v<���P˫��2b+�{*q����ݢ�]f�5S�\�h�N�����n�81q����ՊZ?f��`�og���3��K(��IQ��>�稉����e��^�էP�S�Uiݝ!�L�VKk�����_�k�09�X8�`b4���m��I�|{�Gj��rdq�/�MZ������br���h�ٲY׾��xy8��b�w^~����-W4���Y���f��9���˴C���A�O�QU���)�������S�W�T�Q;���ܝo�ڔ(߻ʍ����~kP_KT,���Z5Cb���!/*�r%���j��h-�g�p]���<���{�נy}c+cA������\QxⓍNܕT�q;��t�[�e�n�+w��~�B�d�յҜ��-f�*U�*�[�<u"=U�\_R�J�
[�\wX�o�݈D3�'x��Ͻ�����d�F}���e��BF?�;�M�$r��ܾ�]յ��"fO��(��4�/�tZ�t�=�k��W��;v�m�Vm�fhhV�\4#�Y�&i���{�'N^fǡ�9��Qȥ���o�hxE���d'U��mZ��*����f;�K��չ�>iV�Gh
��6�m~Qn�h�y�����4��ƹ�W���c6`d92,?�`c.�{�'���bs�n���x����H=&n����Ԛ��v<�f�b
/-+�]R�p;=;Z�*�q��n�5C'U�;!�lٷ�i�����꽉�R����n�*�P�c"��ci�X�ˋ��Y����W+��Ff����4��} �}�9�F��ʸ�Z�7��"���,hx��=�ޫ�^�>��欫�I�����@�W��h�r�2�ҷ��2�����.�N�B'�=�S�1�9�{�o\�T��Û
j���zW �#�dq��]�pp��Uw����MU���u�GBZ��v-�� �y7(ޗX4�2>�N�?!*�T-M��&s�􉦠�ˌ5nb��u�:UH��=��%?SßH�r�W���]uz)'�V�Y�{��s/���;6�)^Pc��<����f��1�/wV��9e$�������;��
!ҭ�e"��]�s���R܅k�\��<]Z���&&z?*�Y��Bu<q�z⮳Ky4]���ǖ���M�xS�6���_5y�N�V�2Q���H��hu���3�E�j�M��I�TM>�9 r�sG9�.��ִ�mGB	&M�ڙ`�ͻS-a��d���i&h��5�@�Cqt'�<���6�i�[�P|}�Of���-��x��'���$˅W^J���e�8zU�O����r����Q1�[kP��߆�t�
�$%��S�gO\_wFh:�.3k{y>��2�2�����&�G� 4������7��,����ы��0��1�6c�7���1���b��Ko(�nn�H+�A;�#gW3s��6�󋭉��F�TdM�X%�}w��Q��߮�o����<�2�T��3T���;�z����\�:׫�����tZ�y���s��o�Ō�����>f����GJG��M'��r֬����^��Q��Ո�X˲v��x�x�ͣo1p�1j�B�n���*Z{�4q�g3ɸ&�z��j���mty�)���J��3���u�.N*͐��֧-��q�w�o[Jf�JU���4r;�MGUB�S��[��ѽߌ��,oƊʳK> Y��ٞ� +z����M���sfs��K��cw?�Fd�c�:�󕜒-
�����Y��u	gQbc��Jf)�ϖD���o��T8tc�����T�)���%�.{�t}�2izi����_�b����Ȁ�����^MD90�O-�Y���{�O}�{r�	~�Q\tc����tC(paH1�>~�UI�s8�{�Na ��9<6�B]L*�u�a2�S�@~ ���}Y%��9��4o�%�n|h��':�=�0vG3ʚ��4d�	dT��ž�b�<q���R�*��F���ʻ�Eb��DHJ-r�5v�!萙Cޙ(���L�9�`�w�ܟS�f<�]=䗿KS��>&��	�w� 8P��PZ@��:+�)��yOޥ6�z�%g�F|��ӡ��r�e��,Ls�3��{�m�'a��6 �ٛ1H�j�=�*�PC!M�����'95>�/}G�{�`���7\_�ig�u��?��K9Q>�@��@Y+׻KG��LzpX��&��$!��5����𚙌��@��}o��W����Z�B8�̘�(^t�2f~V�S���_��C��Z��I;�,T��Q��J�����"|`C@{r/Aq>�}j*� �p�s�j/*��w��>�1i�{E��N��s����c�g��e*��ЬǕM���"|m��P|���ף.7|g�[>���^��0�U�n-�y|5]q�_B"ݚ���s5�\gj�,���vE[�n���X�]�i䕗�Nڂ��w^*�d�ʾ����mr���r3�ڷ�+�<�_W�S�,�G��N�=�@����?s���z����t�h���{&3�3vP��O{�/���x=ޚf��� ��>r@����/혔HW�.�R�ً�{�ǾӖk�f���w��!B h��8�=���y�#�ە�[���σ�UC��L�L0�)��F?�����M��V�����i��3C�*<���dǧ����w�3/�Q���tǽ�>���=��j�VџW��ߋ��@J�����-����~~��d�"Z���"b��4Lm91���R~���VL��~��.�������l;��Fr��m/ܲ����?�,�����V��=�1UTN�e�o�Np+ r�Ph.���}�O�5��Sݬ���Y��5��Uѝ��Ո'd�z[z�]7L�k����t�����gp���Ǭou�J�EN��D^��o�����c
��
&^�=7�mV�BvPξ���C��a̜!��-4�nm�9��(�E��-
6 �aޗpt�]��X�n�TO����iU��W3j3�T7z� @ͧ|�`ˁ����ʐq�H��+��^���B;�>����!oF�Ch%G�Y�7��9e��ܪw�l��nj�c���D�Gw
�h*t�םj�Ժu�x�B����\=�{P�wMt�HLl��32� Kj�e�׭]��HF�89ahu�-���9}�ju�
���K
��!��[�)�@N�M����#J�*����;�����n!@.�k1�yr���v^��_�h6-Mn]+j�zwh[S���Ź��#mdM���Еto�V�Df_dե���jik�kU.*�J �����A�˺�\��/�,\�6]�U��]Z��7qP�ͫ���Al�}�z�`�w��+G��D��;j�w��f O^�ү*���[�l�Pѝ8�;0ݩ3:�ov�i&���c5�<�i�sn�]4%��.3��iy�s��&,���Ҧ������̗º���3{)�*�[C�.����o��c`�qs�@�r@R���h�Wab��Ѵ�3�%o<���k�X�V�u�%&yK�d�S��"�wQ�1�0���Ҝ���8&��E`�o��[�/k\�i��C*h�
��V��}ƕ�(��nc�e�J��w��o�4q���:k�A&2�,�j�)��qR%��t �F�[h՞o1ƹІ�b��x�`�u��ۛ�r��z�6�!��k1��lvH�t±[:�	y������8`�H[{���uȬJ��GL�����V�R�5�/���Q����j�T�8�N]�Sr,V��Ab� '�P�@PDQi	�\�.I����j�4*eaW4��Z��qV��T�:�Nrw\��'8Q���yq*J<ʧD�"9�\�:G���Њ�B��\�y�EK1
��Q\�<��' .RT�$�
��U���e˅Er��M�\*BH��Z�eC���F�NȮwZv�B�T�D�m(�w]�ZT-VT��[	ne�U��>Y��]��8iN��*����D^�Yv�#<⬞1蹝F���(W�������S�r� +����f��xz��U`S�4tp�a���tE##E�_x�+���u�5�}���Xb�00��3��@��Ϩ�����E������e=�x��ў�ˏ)�\ �j	����0w�+��Ll��	9麙5;�ߗxO�z<Pڋ�u1˕B�G�@�"�}(Q=�UݟwxŽ^��FY�o�&�o�UuE�`Yc�������>(H͛���+�{� �#�ܪF���N@���&�dq�m�}~T.w8m׵��l�!�*5��7�P��1���"-���9���Rm�;���¢�l��B�M�a�T{�<yX���/���}�Ѿ?O��:V��c�}�W11�,��c��cs9�s_3���+���L���|��,P����-ڇTծ}J���3o��_L��23]*W��J���;���ɩ��,Ҁ�]lf�W[��c4�ݩ�ĕ'��n����dx�	�1;���S��驚;,{ѥ�L�L?b�>A��߮,T!E\�@�0hgؠ���i{�:��yR���π�7c|@��L֘�k�a#�$P�C�������N��E�޹a|ϳ�d#�Vy��^,\+�ƶr���ͻ�򷽫;���"p�zf:�3��c�gB�F��U�e�����|?W�����������(;Ʋ��.ү��&�ԇd{��S��y�1^�S
���Σs�I@�g�����{��a܌٫��k�g�&+e���b���
�4+��:'@��(�������o�������Fd�x�dЋg��8g�v$�6:V�#ugo5���C� �xU�
�q����%��XP�S1�W����C3�}�+����g+��λ�4���u`M5G�t��zT/h٭�E�p
zu������P������ͽ��@�P����c6�t�Ir��T5�ݙw�c8�)���:�Iݧ��)��ʊ� ?��5�:q���3�;C���;ټ���� xs C�urb|���+�1�t������䐀�u $��f;.6��RC2�*��*�?/8���_���H�� +�� �»u~��UCHM߻}�}�L���rG�x���i�T�9��B6��)�'����r��*rͣ��Q�?uzⴠ�Fal��R��#ew�!Q��^7#7Fn?sYC�<vb�=86τ���zt07�@�,�9�9��U*����ދ�4+���:=Jk[;㈁�9(1���vj<�{}M{3)��d�f�m:��A[�,���$Bu�ĸ��]��m��x�i�P�$����5��(KYW|F�D��?ju�d������p,��+V���j�aov��׀�T�L岲���xLiP�ǩ+ҹ�q�<4�
�$Ji�q�ʋ�rP"�6ɝIH�m��QV��\�?W�K���ׅ2��ܘ�(^t�0"��#��y�Q��׎����鎯��'�<�_Aמ
�����6��Ô\������1,�4���:"�)���Ş�^�Q������z�R<`�@���T��X��)Ю2a��68�"���"�X+����q�dg��8S��G��1Ε|~��b��8<�ӂ=�'k�ى�}<D9�jum˨Ҹ�1�=�TW�f�U����N�>�}=��tR3Ơ�ve�'�zbZt@� ��0=��������VY����x�0�9t�bΌC�9�n����xW�١���,)9ezf)��*f:�����3�2�*�W���IC�q�$�=]6&�����5�c�z�Ë�
C:��EM%(����"�vD�������-�J�1�T8a�"�]�t��;��^��+'GRn��\Cev�ˡ���� �L4/J�E��P���Z�X1�QuBV�i��&�E�$;���ו��cGdUdƉ�MYa����| ���R���T�ʧ��c������0�kY~x����b _�Wiڿ6����=�����څ>��ι"t�yM�EYU	1��<�xmZ��1��>�1�93W�ì�0���p�	�������^�*����4}��\z�&|b��w_��8j;fɋ��DD�oؒ,
�蒆��"��h��dǳ�KrxFB2;��{V�O�;/u��{3f<r@�L��� !�teG���8<�s]���s��1S�8ZuP��%5�1�H�;��^/o�ED��q��k�q�ѱ�3��x!�S�T+i�@��`�>�c��+ܚ�l�q���1휨�np��rù��_��P�_���~<a�I�V��V?
��$l?	��Xr4��sq`$c�Xq�]6��(��t�V&W%�y�PM܎}ڡ����{k5�&z���X&"������-L૜��iѻ�&�t��H�-�f��T���"�������-���No�]~��uz6Ϡ��L�Z�0adl�1^��>��0�{��o0,"a��$�c��,�F���&.5�P��Uc�V���p���|&4��#����1T]Cz��.�{�����̔| �$G2�"BjxI����SWUg���vJm.��I8PΕF���D�(V�*rxh����}Fa�=�sS���ɑ������9 ����u<���J4Cr&V��>�{5��w��Q��V}�cY�i�x�l��G�Q��8��
S�����l��^��1식eɝ�<�/T{g�ε�a�מU���~����V�s��P�G���S[�N��c}� ���wו�W�����k|�z��h�荥���
T7�������{d�$tO]&�\};�f;�b.Z7��\�]ĳnw0^L�aI][%���)J��o�xm�t-���ި��H���ɨB��#|Yy��o�j%xz&��ݵj`�)�S=����L�!)����� Wq������KW1�j,�j����c��2�ˀd���%�mt�gyS��� �P�댟	����z�xK:�f���fk�붰ǣ�xу�b��:�'EP<G� ��,���@����%���θu�π=�^� �ڊ��j��{[Ǻ�o�QS�9�)�*)�	�����I��7Ǳ^�[\�b�H1�zJ+��3Ir�Ld���s
D������oo�s�E�x��S��|$I~?>9��Ts�h�vF��5�H�A�gѷ�||�X>��GK HL�3 �6";�Ĩ�>��6*����jk�uj�Nr�)���Nٜ�a�/��d�w�U�`��x�����wR3B��r�1W>=Cj(`�cH�i�%��	��N>I�)q�;��r��,�ϵ�Os#-�_��K�;+w'Y�6s�遼q;�FY��,��j�z�6�u��=w?yК6�A:*��Xb�Ӿ7���Td����Mf���]��CBp��D9Ba9��X����L&nJM��1�x���U\��<DN��{6�,0�U��6��$ �����`�38�T���3�(��}1��L1������X��P1��f�g��kz6��%���u��@���مy��lp;sH�cvs�N��<�s��XF�7fc����G�t\�:�W�΢�����d�;[����q��T�0`TMI��'|i׹@��X�O���^G�w�j����/�.��u
��7ԫ�+����A�.��1o]S���=��@��C�ul\���q�@�{*<�l93iduVɧ#ף�v���B��f�k$yK��0���-j��Xjj��V@�N��}�[ڦ�T���7հ�ή��F����/6�[�"�RRs�ó�ᛓH��� �za}I��l8_��F_�Qy�|���UI�1Q��k�&����nL9@���랶Kz^���[�c�jb��aW�s�g�-���^���>����d����`l�u^Z�����\x�@�?b�FŊΟ5�W�<s�E	����=�>}�B�()�
��pڮ��P*v���#����\�����w:0��>.,t	V�#�߫*9�*�~��=�oo ��'��5@p�xP�!|���/LW�����k;��D�7�aLW��Li�R1h��Y��'����$z*�'��q�%��q��g���8j;f.bp\f��M��������d	d��*�����u��ꌞV<���3��G�4�~�j�gi�*W�>[J����y�o`�;��Y��xo�n�)fB��*naz;��YIpĴt[����QrY���h�1���Ӈ�c�ɟ��F��5L��� S=�Vxm{)��ntQ���5٫ν��9t�d���_���!)GD��x��D�lìs��W��o&���pz�x1r�N�8" 	�#u����V^��ޡ�q���6id©��W��.��cYbIL���|���9�U@&�w�jS��'����#~'���2��"�9�=���]�+{�i߲��Lg�7�X#|���u�\ ɏw�H�1��;�����Ly��$�nG�԰BaM��(��|wo���=�!P��	��h��_:��c5N z�j��ٗ���H�Sn�?>���Ht�	70��	]_��y�������������`�B逌� ��= 5�(4���ݗ�W��W�Ȯnr'��?�R#g�R��V�Fz*'d�{�Vx��,bG+�$�M*�u�+-���ڹP����]��0f�f����\�=�F��(1�h�Nj���-OD��uk�j��n�ާtr��K�ʕٺ݅Sh%����pUl�������N���˹��F��1꣹�}2\�+���CU�\Q�����V�����t��)٘��s�(..QW
U�v��^P����l���B��e�@����aDtSGy��i�]r�7�vZ/{v���1-(n���X�s㔪s��&�l��]��K�eŴ� kV��Ks�FٝV+V�أ�y�a?lL�֞b�[�>���s�<S��¾�i�A��8�{3���nC������Cz�C\�Q�5:Eu�A�	�wjKXν����
��K�]�|,�:e�׉F���7R�|�x[B�=�}���R�5�)hp'-e�ĈO�=w"��3g*V7a��\8�d{²J�*�=�@�$^�}oe�-U�(l�@�'`Lw�-���&�sѵ����oR�xf|��lJN�WfZm}
�&٢��vd�Ԝ஻6�A��������R�s;/p��u�ds7�Ƥ��6/V�D��e[1\f�P�2�8�Ҫ�-�Q���x<�9e�o����%Z����]�.l��ˮ��bJѫ���"��?R�����I7ټn�;"������9묶�o�X��و�x��;�[;V"�|��\G��r�oV�����M�*�i-dU��o�D�7W!:V9�3(i����q,]���d]륪I�]'f�7n�m�*��O@�We] �:M�s%\4��D��N���fm�U�U�Ǭ�	��^�GZ��|��E�{�u�Jy�ц����B��B�3��\.���HKg"&�Ҝ�
�s�p�(��E�t���vU�t+�F�"%�e� ��UE;���2���*+twZy+��e��G����J�w' �+Nz�9���vV�^`g�n�P]��9ʂ=͇�w%Q�sʎTWe8�DE^p�".EⓄ�����t�S
a@Q�u&�t�("T�EC�^�&U2����"�T�r��Q�"�	�;�N������
���'Ov��(�\��"�fr�)����   |"@&L$}!��I�aY�u<�-M�쭚�R��GYd�2K�:��x����qq�zs�i̟�;��V\�х�����&8�5�1���TM�o�0�o����"�
�NkM����r�2.�T	�a
�7�V�a�>o���i
�d�x�>���:�N��
�d`a���ݙ�э�ã�w��.���N��GBI�o�o�N��.ҭ�P֝�W�ߟ��F�FzX�GY�2�TbR$��o���}�[F5y�S�4"��{�
�TZ,V)����e��@��io�������|n�G����l�O��2����s	�Ee59d�����>�l�	��peC�À��gê�:��x<%�E3�p_yM{��s�b��"/d*�.t0��x:���m���F!!`��#��<��:��z� w�W&��1����V�1\�͸��ˈ��{R����k��n�9.����wZD�#T�lJ̊��i�������&�t���Z$���N�NY�OMV�h�S Faד�ò��ef\I���\��U�Aq�>'���K}�b`q��f;.#kDna�5L�Zj���84Pr{�~����j��eXۗ�ZdX�+�)Bv��L��&}%�I�̩�ꀦ1�s��R�u�{yez(</ޜF�&�ŏP[޸� 0�fa�|��l7��{1/r�����{� ��VN��
�~/}<�@�,����⛚�� �V>j���B³�誅5�-��� o��3_�!W�s5��P��rǯ�c��Zs��a2�'<_U��V|�uow�ǡW�H����'�x;S�3��5Ia"��{�>>��x�3�*�
&3O�Lo���b*�1�,o
���+��{��qV��G ��@���xՙ?�U2*bqc�Y��<���CW,�O�!}���ZS�:'�s��Z�0���m����s��8:���6��ݰ3�-!�����y˗]��R��%we���ð���5��ɋQ�Xe�st:�YW3x�#?�������)���(�{����B��5<���b.����|���Ȑ�+�݊�I=����xcd����Jr���y��A�&�y�\8�u?�F����Iz�q�~�g: .g���z+ѳ�w(���}AT>s�P&6R �q�b�O@���^e/G��c�P��ܚF�c��� ���&): WLoTo��/u��r���������0�]P�z@>=2����O-����'�|<(��W�ë����g}U}0�|9��ޟK�4��cL~Ŏ��X�4.(ر_gO���y��q�yyݲ�Y��gw�w�24��ШG�5<na^�p�3G~�c|+]
Z;(�枮A�GMx�G�xQW._��J,*��@���j���~��,�-�f$����B�wX+R�	o����V#�����H7|4�լ5(���\��Tӽ���;�)��i�zJ�oqWv�!��vQ)�럲�S�?^��b����xR��`u,*�[1|r~��%�|����}uP��qM�V���c��:�F-�)�	�"ё�ϋ��r�Sj����wP��P�2e����GnP��1�y�>�l֬aF�ꌘ�t�c�U�Q���
�����Y����\j�o����A{���1ӹU��"N�몉��{Ƭ�����&�����^�y6<�pϵUGX#�h�Q3"$��^��+;�����K��0�_E�1�8<,>���]:��N�� ��`��%���x2y�ƣ�0�r���/aT1�n����͝�o�WS�7���z@1=8��@�}2��!2[�Phz�=�}E�+��_�@#K`�t�&
��ño妈�تzn�G�[�z9=�|�E�}3��|�;��/2&Qu��i��l.�5t2s��w����T��d7BZ+���j-L�!�8%�+����4�m^�E,�F�v�_�I�kl��?�K�1zV����m��5,��w<P�:����W��L+aTp��d:�9�&&4���c���/*	�]�Oӝ�lߤ��10�S
d��2��ȉ�rƲC�<$��d,p�y	����^��]U�G�5(}^���0QP(n� �����k��x�O��g�s��g�C�	��3Qbٮs=#j����淜{*H��C2&ty�A�:#\�kL��UrXC��p�W���w�{�#��Q�bc:l��Ss����a�fF��½!�s��7�c�L\=��b�u�c�K���% T�|b����*8m��=^��ʣ��s����u���Z����3��P;�ٹZ�+}�䎰($}a2�ao*��,]��,{ǆj�f�D%<�7x��n�7Wk?1���l�5XzO��ݟb�+q��ʇU]�k/�볢�D�..��%���1�Ίͅ��^lR��,��W�g?���E{��p���M.��[��]��C?:^��R ����[Tr ωa���߁CB���U�qs�f��@ۣ�֯+{���D�1��#��A�:D�<zp{���q�.��1�f<zQ/���0�K pH���[Q^s�w���?4��p�a�>%��@1P*:tc����T�Ǧ[���=�,r64P�P��rY�z@^�0��r��O���^�E\�Թa�e�mZ�ఙ˨^5�)L����c��q��NJ�;o�������	�ܡ�lH�9⇉��1��Ǹ���+�:��2R�8��E"ɉޞnb�'����秣�a:�G�~��IqJC�`z:pKst�{BhU���fl�Z��R�c�+i[�닏`�{tEt��]�U�mF�Z��6�/P�|�W�y�
o�J|���V�O���`�!]��ǔ�[5/I��I�W�܈S����ep�(��W��`�Epwp[R�=@	[�8��s�/���	�|4;>��&pFGX��Ҭ�3	����*,8�^�;_.�)j����mH��1��x$ao��Nt\3�c�:<���7�@V���cb�c|oLnzP��z��vL,,_Z�#�{��X��fϨ�&�P(�xz\Ʈ�1G��h��q��M���8X�� k�UD��f<E����b<�N_&�)ƍ��7����	T*�?�1Q�<�S$z�/��M� �/K�4X��]L!ǕB�����?\�S�EÎ�U���l�qC���nP�*|��P��Cr�t�5��Y
�Vߖ�D�Lp�k�ò𱱆Q�;,X���&S�����j]N+�ȱ~ HA�Ì*ʐak��H����:}�ƁyG���ֲ֬\0~��i��D+��ք@z
~P2�MJyA�q�չ/)���5��E�bw+���+dS�����Wnr[��'�:4	1���s�g�,��<G��W�Q���ѕC�U{ܒx=��Ҙ1��?�%�R�FŊΟ5������pǶU@�,<|+��R���U�z�e2߫��ۤ�7w�����@z1գ<oT:,X�(t	�c��kOU�:�7�wz7ۭ��@�ۯ�؀�q�lk�/
_w,�+���Ns�ޯEY#��=U���8<�b��/�'YB-�1]�q��o�zŀ7�P�*��ި{�L�s:�{�-�	�͉���?��� �H�E*�ڪ���Gu� fx��`�d����;*�j}<���ǰP�4�G��F�S1���쁾����@�����Se�����XlG��E��e�d��y�r=&: ������B��R�T1.�/�ѩ��b�B_;��v�ţ��LIƆkz,↮��/�r4']�&l�U�:n-owrh����m�`²C�F���F>�d�_ 'r��U��k���=�T�͏�<��wӨw�#�*����3u���͂=Ӣ��(G3�s
�*<���P�[�����u��=ا�'s<���ǌR���|(Q<�xÝʤa2CU���\c2`[�x|/�ꉊ:Ȩ�ƉCx�F3�X�=9����м�y]]jэ�O��K�<Q1�iύLvۨSR��5�ak�=�!U����=4LKc��#ł0��Bt���X�$_.r'_C�]��E2���Cg�$��	#QCѮHt��g����i{ㆎ^�n��L���*��|C��q����w�7���nz��x
���:�p�v!�5P�ސ&4�<"�M�9z߽��}��"�E�N��4=��Z�3Zd]b���(6lP�mNX�BzTU��³;��A�N��"&�Lh��I�#�<aWt w>��� +61���
c��2\KE r�.aNh$̺}q$����Rm��6{o@ۭ��bG��z|)�O<͓K"�bU�Uk|x^%��9B�x��M?gg����Ǵ����i���;���{It���jm����pM�/si�L�E��z��G	��b�B����DN�����4�����R�;�1����f7��0�����1C�</=4���T��6����MϾ'@�A_�9�U1�j�v���+LU��΋��}��o8�8����Xh�pO����e�����z�#v�w�߿~�K!���
e3��A������&�s���֯ �z	~08�x(�u��`	⸁��Jٍu����9�܇9%Ԑ��7��u \&&��&f;=�\��}��R�U$y��Q|,W�LLc�ϼ@^�0�d
������E�+��X�]w��v�?�nR.4(m,Z��vb�61 �3m}��E��ja��(�v����Q*�;��B(��B�L�t��*N$�EK���o��s,�L�$��T��]}��o���b��&U���j�-���� 1ƅ �\5Ee����ÀR]t-�+�2n���L��4T��9n_��u��X��W�RCu*g_n�����fK��Kc��i*p�G8wQ���m�#td۾��92=��4�>5�!�!<�˲�/�j���sjw�<��E��)g��\��=�SJ�\R�^J�Xx"J���ge^nBjh�%��qS�rB�o i�.� XĒ�ͳ�u
�;Ȁ��6����~s�6��|a����'�h}�[���l*GF��{��.�b1DU�U�l_k��-ti�m��\Ô*L�������� BS�7�)3�ݘpZpP=X������u�5���}v�TY�
{p��.����Tni)�G���}��ަ!,�̣[M��U�#[3��}q����Aٜc*������R����;��g�SśK{0�=��N�N�v��q)q��ZvZXdk72�;��c����p�JS�Y �P���3�#����zlnu2����/������7Ѯ�={m�5r�<��#��ሤ�Q�3i�ϴ�;ehv��Ю��9�#I�yr�����1�r a[a�KGR��:�C���f����.ʦ��,ù��ZlZK��%W��8� �c��RT������/B���/�Ձ]��`�1�V��*�Q��"8f��;�Xt��v��/k������%�~�ݔ�cv�SF�d���M�wI$i���X��1ٝ�d���*;g�[L�&�>qӍ�V9���%K�i]�0��7�G��C�cr��4�Z\��(N��s���y�������I�;��:*� Y!�Nj"�v���)˧�z���w]�q�]]�8�K����)PN���R��铭��74C��p�/uH%2��A4$�;����'�{��=�tE��x��'L#��R�K��g���p��$��/t���֛q�t�B����,���;��'wL�.��r(r�p�
��̎D)��C2���Wpww'r���{��j�������V�'p�u���R�8c��-3(
��JR1)�D{2u��n����t�4L��-4���L�0��k(�U�����=W7DrQZw]=���)�G�XE�,�uB"�p���s���B�'<wp�qvI��3\M���U��&��I�Bz�2�kB�VQ|n�P�ť_:���ĉ�QU�l؄����!�kD���n)ӝX�j䶼���hX���;��G��E�/�K�T��L檨��E�k��}Ͻ��.�1�0nX���5ơ�5P��Ǹ�#���{��1g�`.���	�� f�b�������J��5�C޹���G8gLR�����]_NК:����Xb��;�c�w���7�׶�%� &8������Js�:��Ҭ�3	�z���ٙ��3ޑ��7�5l��c�t%
ayN�`�՛�9�����<şA��+�G���3Έ݌t�����d���/Hk��՜�(��x�y�U���*�2���L����c��#�rg���U؟�	1����*P1��.xm}r���ٞ5���Z�M�S���νQ֝PB��H�	d*�?�1�x<�=�-���Ĉ��V�0(�B�q'����y.�k����v�q��W�P��\�t���q��&f���+)�4�����*��<��Mo)]�SHc�=[��W:0۹꟫҃%q���U�B��L(8���u}W$
�WT�b��<�K� �h ѱ7(QR�ja�[�b�]@����o �9�y�8z.K�Ƅ�t@0�׋�Qωc�,��Ǿ����{ϹY�@��z3H�♊�*�B�0�]P�z@^>?
ۉ�5���/��	��	��FA���M��0r:bɛ<G��h�o��{;�/J����Ʌ�11���E��SbhرQ�>^��={���.A��p��Ф30̍E�Bc��������U~�c����=���1�X���t��$^�����U�~�>���u�
��T*1H�6����fѱc|X��N
#k4k�=^C�E��-<��Dߥaa&*��Q�YZ�1�R�x]{��<6�=:�y��W^pE��A̙��#�3I��L���i<��G�~<�ߦ�{�0��b,����yތ���fB�u���{\wz�41��Mv�QW����1岅�Fχ몇1}뇄�s:�2=��;�y;#������Y�e#�1�&7.@�$`�3�uOx�Y��\�zs|`-����� ��,1l��;�ꡨ�q�5�) �:���MѤd yب��J8�7��u��Ӂ�'�68�����>w-L��v���վ��^?u�3_<������T]B����b��bi�<��Uͯa� G�2&� �9c�jL#�ϙ�Zj���_�Z�@�M���Ƙ1�� ĩ���X�D�5��9�r�UU�y��g	Fs��>�H�)j<�&(�G\@C4��'9����r�j�?7��#ў����@�o��{��,��^��ST�9�2���/y�懈>�'�4LN��x�j�c`����1�{]�<=�w�� ��kxq(�g;B�"���z�{/�P!�8nI���J�]IZ72��}����I)��-��w9QGJ��g>Ę|Ok�<�:������'q��љ��J^�Ys����Cz��2|X���\�ߪ}����'�r�|���X|#����ǋ�5��>��H�逊 qn���;�No,'y���ᢾ91K&:����,��c�q�O������V3�hȫQ!Y�Z<��騲���3Zd]�wmr��r��C�_�{%
����U��Ɓ�J�|P������ĕ]���<	�dK(0���|�����{q2�	'��x�퇷�zv�������ƥ1�s�
�.��uӢ'qTe�-w>����tFb����;ƾ�ϙ���-+ŉ�zxU��k|�����7� �I�;���蹎�Vc�U`��:TlˍF���z.naq�W��>s"~'��(hW����tN%����e~տ�!ׇ��'U��)KgsF�Gt@�WP}rMFL��;������w��S�E��훺��-E�>�NZ��2C�)se�kF�7*6%g.�ٻ���=�N��]K�� ���n�˝Y:*]�aC^�ܛ���Mm{���$�����:��,�q�@���)�[�J�G�υ�����D�{�,	�� i����84A�^�b�1^���W�4���^P�T&'��>7��0ŗ qr�k���q�;�,z�Tz�=~�ଙ躄Ϥ��d��0�a�.I��{9��������#΢��j�`������Ŀ��
/��J��ŭ� �F@�1��Q|M*�P:6��X5���������?�e��^��椇�s��`W�(w����V��f��6����b����9���Ny��Q�k�7�Q�����;=����x&4*%{�Q�����������q��H���Q0�x+�L)�ӂ�':&~�_�V	�W_���J�u5չh����9)Ŷ��K�P�m7�u��+�	�u��rru��,iވ�l��96U�w7����/s2T<��s_)"{�F���ܼ!�fUp:�Ą����ޘ����b5W:�b�$����Ǣ��a�z@��1��(	�U��G���vt�_j����ǩ�Ұ׏�,�;��9�UA�(c���ƾ�b8{k���=�ٱ��qc���-�̆*Ɖ��$�0NnHw4�)�x_�>0�Sc�&|0xb;g���AUB����.�(p̜���T��V�x �hx{��3r�,pC�0ė03�;\.ߚ���ωǠEOeEB/��V|�ɤ@c�|e�9v�]O ���pм�D�1�C��I	��*�*
�]P�r^�׶���&:8�Z|N��Sc��=6�<7�a2�iױKѾ��*b���*��'��>�F�cԦ��lXS^G�{�r�kq��ӆ����ggʬ*{�9��2�VL㺙��%ѭ��5R�4�Z�w�˙.)I�:"
�hٚl�f��f:�,������ǚ�od�~��οS�NC2̎e��Bc��(­�7�Z�z�ϣEњ>g�U�ԀF|b���,кX����o���?+�aѯ<u�Y�ì���]k�l`*����,G���A�y�k�����"�b���uP����b�1�N�ex@�V7���.�������s޸w�,�\Σ��$��9����q�����'��W;]c����?% ʦ��c�;EH��tμ^���͌���M�Ǽ`���o�e�H#��7\�c�y�~G��	YcQ��ޜŋܘ���f: �Q͏��r�X~��z���}�T�����T�����	k�w�o����g��(_��������ʏ3���3�w������%�/�LF�V�+n/sQ�������d���k��..;��Yc+t:&=������P���\�:c��{Y�N��s%rV��2���az�!W3�(x!�1� �N`�B��j/�*�ޛ^wV}9ݾS�gǥ2G���Mȧ0��(o�CE������V� �{��OޗF9��z$�?{��RɎ������sӐ�W�kW����,:&6=�z��x�d`�����Q뫖�R9�*�m}yQ:����	���b���`���zw��c��.�������xBں�7��M}������ꂈ�y͟�|�o=���ד��'��N����Pa�~����)<9+8�"�e,]�gN��
z{��Δh�Y��9�5e�/\�r��p]j���"y�Z���}L��3d�B��WmZ����n{9��Q��xz�fFϣ�<�c��'?^�L�RV���y�>��n?�3�:��W��·e���I.�r���	���;��{u<���L-�;�^�+w��} *�s�4��p�h��ÆF�����������ڭ��^�=s�1a3D�/LhY҇��p>��6�Ƨ貓���w��>}��5&� Mf�,����[�'�R��)��#o�a��}�WPS��V����MA:$;�9�U1�j�tƪ�v/#�����>��Cz�E@q�ỷ'��(hXX��z<��2q���8�K�����)���b��fh�������F�y_�۶�@,6pd~1PzY<��p�}�q���; /^o��V���W]E-�.��D1�D�\I`{� [LT����>{�t1U�_ziQØP����%����3lW����S~M�xa<tn@4<*=s
�1�V5u	�Ia|z��5޺�o��,��J��,�G�U�Y�����5��2F�@l}̱�]���`��k�%(�����=h����(1��}w��<L���\:�f�K�7 ܎�	�[��z'��d i�������r�:�RN�-�(��_���r��d�Ʃ�,�ᱻr�aw�� z�:��ǌ��O��j�q�,L򢫣�P(X�p�<\+���37���]�㌁��Q�P����������X����X��Җ���P��T�Y8���"�������>t�?;�{���z#HG��9c�V��Y�F3�Di���HW��L��z=�w5��.���K����=P���@�K�Շ�׷�f��j�zHر�x1�e��@�5���\J�1��/��c�W����8'�pE_z��Q��:�x�
F�&���޿8��ٞ��ϭ�l���Ll����W���w����!��P�_f�V-����Ի���,��tOCb�Ŋ�`Tb�z�|���������P���O�Dʪ���V��9���X�9�����%�PPլ��D]�&Xf�����%o{�yԵ���8�P?\���X��B  ��TM���[�]���h��̬�!���@EC���ٔ�q�8b�~w�䚇�u���\-nU"�%���L����W�pоz�`2��b������\�T?��s�ezz��@ 2�EC��"*�rF!%hv���4�!�?��ۃ���$�vS���s,�m{�"N�@EC0<��G���l4�[��w����fo�,��{ɵ Y�kP��І����<xsb1k�G���w�?g�r����gh���w��R� &Q ��eEQAsb�
gq���l�4����AĲm�>U5<���$�/�86�q+�� j�Wt�J�ߢQ+�����B�O3�<���#/���:�TT-�ˤ�E�i��i�����r�| �~GE�%�d���/����N`>��݀�m��9��vx�nF�PP���9x�C���,��g"�$���C�#�P�{�{��"��N�&%xPk�4�y82,	�a�?
""*��C�4hF�����P�č����.��SM/I��Rdd!gD���!&S<�X�(qPEC6����<3�rT"�G`&��v�9Bzv��u4�l�hq�x%;�8����
��^�{�bڞ�Y�)���+��Ċ*7���#�G�L����$z�	_K�X�C��OC>�K���7&ǀ46���D��"�D���J�AE�u�~�x������d>���G�����������m�Σ�`ϰ2��"�g����n����7��.��
�!�Kۨo�!DP�X�`ރ�<�W��˗V�EC�x�i� .�p�鑻k1vW!l�Ώ})b鴂 ���H���G^O�rE8P�u]�