BZh91AY&SY^7�^�߀py����߰����aR~x��             2@�   fԀ
R�     z    �    a�B�     P w�� |   ��=�{w��.���z�v� w��{n{��ޞ�twg����'{�:�= �b�/�������	�������
�����}��>��u�s��[uA���}|�>��ͭ��W}��Hz{�{�t1�t���   � v >��^��v��{�{�B�F�u�Z�\�>���N�]��O}�>������R�fy�د�o|��1��ׯZ��p�����o��U7�ut�˺��]ۅ�wsA]���-�  � 6��k���l�v;>�y/.�[�t���wKN���<��a�:��]���k� I�P���a[���tƻ�s���nMW;����	s��m;kv7vN�wx��  
 �͖m�nV��ȷV���ps�;�5��ݬ�ȧa�V�\�Ñ���E��6曐���Y�s�����緑��	p%�mn��u�6���\    ��z�˹3���5l���vY�X����g- wi.����\F׽ݓ۠�`ǹ�)��js�su@˵�wsg%ˮr�@                 
� �@ �             J��Cz�R����#@ �C!�����BITHCd�ɀL	��QҩA���L��04h��@T�$���U4��d    ��H���A��"12��ȞBh���i�m=@U5	��J��z2  M �?�%~��ċ�/��8��W�?�?i��?vƿC�E /x�/�  �eP@ߐن�m���m��_}������Z�\y����q��*J�{l6������prr\����`�4hd�����n��'#�����������s�����?���̽��z��L����r�L�/��B�d���9ñ:��������E�>I\��I��x|j{MMN�ZW>ӟ'�=����ϱ8��ݞ���E�"sǬ�y=d��s�H$h�q����>�9Ra&x�	����j>0�C�p�s�,�"NFO���rz�{��>y ���ȍ�?#%xOx�����g�zWL0��J�RY�G��$���<�t�������*��[��F�'��Y4Nw��89���ȉE>���^�M�_?y�!���'Y"#�L �"=��Y],��NܮGbQ|�&�I����w���r�j">�_?z�`��N�)rWK������Og�<�l�F(�����%>ߚ��nJMۑ7>�"ܯ쯟�JD�\�	�e"b�N�l���%"[�H��W�5�i��J��ep���"q�H��,o���ԤKrR'_�"ܭ87�_?>��~�\�DŔ�2�_W�J��1��N�+Ś�4�e�����2��w�I8S$G"Q�e'�q�C����)͕�9�<�S�d���*������	~j�������"50��vt��㌳�9���%C��	"�mW����N�RmM�WK���Zfϯ�Rl��u �#��݈��pjq'^�M+��U�G���#�GH����'��D��#�<�Q�3�r"�$��]-�(� �4G~����4��~�̃�$;��w�vC�5����c�+}$=~��w��τ�f	PK�z	�~��+ҥvT���%��r�Ԯ�euei�eo�+���%S�YE�*��p��X�vV?M0�\��ʼ1�y+J}:�WVWm�F�+��93�ܞ�v;9��2�R��R��;)gNy�ܐ��$9�{.�):�Wvuj��=֫�'n���$.&A�g%|���2�U�ʣ4�*[UYR��9�}/�BӅQ;9tK�XR%�N��Q+��&��$�ړ�yI��d���'�'�'o��4�Rh�M�QXeD��-3�5I��OIx^��8�3N�#ҍ��~9���J�����7��Bo�4�I��I��8&f��s!/�$h���C�D�T��̻��$>rN������Y&�ݒp��'�'�d����d�;l���d�y�zm�w��~�w⾲��<$=I"F�I�md�]�����u�<���C�¬�$-%��I�54�;�&��&��Dߺ$�5!�&���=�j'�J���<�~RtKvG�I���"��IM��N|�=�50��'G�,�	l%��A<xM-<> ���'-�|��7'���%	�I�Mp�tf��H�ޤD��Qϛ'�I�'��,vM&�Ӈ'�ѨDI~'�"y4I<L�"%"#�
ԔrY,N�DE:P��8���(��DD�(OD�c���4�H�9Ԛt��<W���"w�&��u�t��	�{�ݓ��i+�"&��(��:�#�
�b���ji^�(~IGN����G��"sR|�p��M$���DD�0���"'lD�$�8C�Qo	������'zL�D�x���G��L9�+�$H�$�(~���8e	��։P�	���'ɚ'q'r����K�I�9�4���jx�ː~4얕gG� �'v'D�+��;:S�螡�vv�F�D��gY�2��r#��O�4��M9s�rpĞ(j%7R�������Q����r����JlMd�7�}�3��M����8�L.��5¦}�0ϸ�E��N��=�+,����<J���0�o�Cđ�*#�+tGI�xN�ͣ�$+%�#�TF�z6�6���s�jp�~?w*~��;<w�Ƨ2':��|�;֧��C��?i�85¸&���z�K􅞓�����ӽN��N�Wj�p��:`�";0�,�:]�Ng�l�,YӅ��<� ��D錇gj",������TDs�A9=RF�#�TDdN��<A��n�|�+"#ݨ�LN��J0G""�x�L�2�gȍ��&-J����"xY
ʞͨ�+�O���SRt�$DzH���p���n�"��i�R��Z� ��:[u(Fr���mDL�T��"7u0_T���Ƨ=�"2�i��TLrH>�DG{S�B������"/�&��4�=��ϓ��R�g*"7�2ڔA������'ީB3j"w�!���ɲY,���W�$��=Q�����^%'��Μ����|�o��!�9(�{>Gҍ�
g�=���H��/��Ў�6�ߒ�7�}w�%���;��+�qډ��t{ҨG�>�����&Ʀ�������d؅3�X�OC(�t�fs��FO��m�j��WEv�'�� �|�Gg�w'�Ϡ������K���4NH���+���%j1)��:^D�Υ`�L��v��;.h�RY$�;Q���G9;�D5�h�j�SUSiۏs�=�{����O��(�>�ʨ��r�>���S�*s{S�$̖˨�T{�����j&��rM2Gd9%^�=ʏyQ�j/jSʕ�{�9p��#���>ʏ����=MN�S�/��Q�TY�{��S�*r�D�L�W<w�5�	��Y��.��Lə2�p'��}����M��t�x�'�uw�4jg�Yz���T�޺�������"aݕ'$��{G{Q0MʩꞍNT����S=+�Rf��مz�Wg2_d���t{ʏ�����������.r5!�;�م�����G��)���;��o	=��N�T~��� �w�����;'cR����:\Z;�^ ��G�G��_q�U����۩%��;�8wg���<r�<Tە�D��jY��e&�쯟����"'�'�vI��G��+��~�ܝrWȳ��DѨ����G�K��D{l���R��#��:�E�],�������W�<�l�F(�����%�g����H��N�DE�Zpo��~})�r�&=���):e������o�"wY^,�5�ic|�����e�DN7)\����>ߚ��nJD��D[���+��ґ/�+�c�I�M�N�l���%"[�H��W�5�i��O���eY>�ܒp�H�H'���*��.J]�ݜ؞g���Y�̕E��gy��'�����jW��"50��vx�{�VO�$�O�?s����_s�eQDߦ�9�>��4GY]/&���۟f��Ԟ��rAȏgQ�lG���S�u�$�*�h�X��Ӄ��I<q���w$�9"5:rDvxK�*��Q㼃 ܂/�G�T�z�?i�A�;��첾Gd�o������&��Ȟ�~9�ό�L����v	�'��[*W�J�W))�y+J�[�ǒ������I3$rU9*��t��X�}�eq$��z�WnU7*�Jǲ�N��Օ�eo�$�297������S�9#s�.Nɜ�����]�e�."f$�b��W��� s�/�E��(��)�nT?����~0g�����=��H`?"�2�4��������`�lB�$b��/7�����A|�{�Tg�ü禵�9�x�S�+g3;�m���(�ȡ�����4Xs���	~�vK�����d�]9��������qޙ�o��sju�=��l�1�uG37{�s9��ߑ_	�'F��b���V��q�u�ֵo�o��j{��'�$/�]�)���n�Q����S�γ��^��/R�yԟ�ç��u����I��GP]�uh����s]<�d�����������)�N�R�q������9�yN�߿>�pB���#[���{y�iw�~����ی�;���N]����}{�u]�}�7v��=��Sܷ�8�Nwx��v�5r�{í�;�גuU�>�P�������wz��rў�ګ��1��[�)��3������?%��e�4��/�������-��}�ww��6s�p�����ݎv�Z)6��{��t�s��#wû�;��9վt�Yvv{x��o�Jz�ԫw�O�������7����{g��Ky')�5>�j�nQ�ų�t݆Õ�o����VW�ZO�<���;���SMZ7��/����w��/���>o���W"��!^}R�������F��(��>�칙_}�w��5o�q�<TsuY������Ow��輪�͛�}�]]�g������N/�>qTq�*m�E�
D����������_7�ϻ�H�(���O��$��!�=l��]�N}��ݜ��v��%��99='�Ü6��9�\�ܺl\�h�����r�/y����,�}|N���|��oM���nz�]=�}蝰t��O?L�*�����wuU��C��[��F�W�z,zFߙ�H����u��'),�_.ɮ�{�^R4�K|���������DM�ﾛ�}���Y�*֫�;7�ÝI�;t{�P����\��n��}um���Y��&{`��޳����_�]٣g�{ʿL�!�!�Ƕ������w���ّ�cu|2�9H��w��#��9�g�œ�z-�������άsdI�A����t�q=8�=Ɵ2.���4޻�.-�=����^^Q�ޫ��8��>��mԏp��ԠǬ�<ۇV���ֹ�"d��4oI�K�Kq�������/h��ԙ�_�=[C��̂7ȟ�����Ns{�47dn�����?�<�$&��:T7M�{�-���G�����1�i��#ģ�.����	�{��cD�7Yx�R��>���F4��z��7nz.g�x��&=JQR�E�4/�N,��+�j}��Sn��#��r��'����n��h�H�^��F�P�P��Nk5T�/x���awM텆�� �ш�˓�)�<�d�q���s�?#��a��>g�aϗ�W$�߷>F�D�ݧm�x|����=���*ĵ����[$��h�5Mo�xկ��D�}��65y��s��@��64�R�S\)�{�ޏ�z6^��|6�S'��7~���W�dQ���������Z��mEn�����[�rxC�����1�p���k5ij��N7���wg{�8V�_N�ƴv2�μ����K�q�G�}�/(����<������E�#������f�M9���?p|]c:�&ÛD��%�m'��*%ҫv,�J�N|�9��f�^)��w�J��ӂ=b��������>���b�Gi�T�#fl*��D53�5'�<��s�*�nu��$Ʀ��v��f��|��pw����R������:iF^��������#��V�B�.<�K��>3��)��Æ�5��^C^�=�[�ԞC�E�I<s�#��\\���:#�/87JQwK�4����q��7��=7��_1�i�-=�]L�wM�&O,\5�[X���踝���R9͚F���t�^�?x���s�Ӛ����:��*J4s�w;;j��W��{Izs����6e���9�ZPs���zs����<����d\/a�mul�y��8�)ӭm-C�Rb�!\��t�~���m�x�o��s����4p��i;m/E�w�߽���"�'܈GkĎm��&_�9����̉d��H�w}�Kt]~���ҩ���*�Es�oH"�cn�������:��uB�^��v����݄�5u޹��k٪\K�G���b������c��G}��6�I�M��0��Rn��w�Nj�7��h��R��9�j�U"��-Bu�"������ߵ��Dڢ�ߩ�|��K��M���;.���C�>eNc�R���/t�.�����]�-�?o!s���_�Ù���-Ih�r�8�0����������T#~�Nw����S����u6�Z�Z��i�`��~��|%��Y}�Bx�dּ�R���S��+X�8 g,�eLV4I��I�uV��5�Z�"���+�zn����I���)��pM��[���9-ER�W�n�6�*�7j�|/��Σs�o̩j5���㡼�->ӻ�=��rps�)����~���ozsKx�'ͤ��~.u(>����~����߷��6՟/nT�o����:���0��;�|�jm�l��^Q�Pߙ��)uj&u���W7���2��s-��9���'-�}�����S��Wa��Wxy٩�ݳ~��G��Ա1�b�H�ߝEzv�����U�g�&�M��6'z���ד~o��2i�3�s���Q��_���aɛ�~��Ct4]g���y�$;�{y��>�g;�M�Ӛ����G�����8�;)��E���5X��m'aRF����#��i\5�t��nF7stn�h>�����������Ӥh�����|��7���;�<	��3���t�xOkR���Z�ue�tDe�>�������M�ѭ9�_�s����Gnm��OH�\Ԯ�(�.��ӟ2��KI߽f����M�8-��Q}�/xr��W�P���s`��pC%��:��r�l�(A4���d&$7��jW1��k�vN�y�𝹷;⻛�����M���iv�N1�����lԌ��iI�2.k�dp�"]�Q�I^{��sr�r�5�+��:��ݥ�'�H0汞�\O���:��-�4���I��������v��je�����I���+�du%,{�j��Q�Þ�'x3K�f�o���+ϑ/N�-�Ώi�e���5�j�R��s�Gz�ӷF�c�ϩ��Z�ʇ�V�^T5����
,ל�hy�mM��������q�V>s>D�n�Զ�'�����u��T>��C7=J�v����3^�A�HN�������fq]��!�p�|/�{f�I�T�K>�}g�5��#Ck&Qz/C�M!�E��mY~�v�D�w��6���ؕZ����PkI�7�To���o�$��{�*Q	!z�q#�F�7��x��l�q�Պ��7Y|�N�|7>��M�������?Lޢ87�����y�q��X�~^D�s�l|E��3X�=8?S�^Y�9ܨ�^&[M�V��;��>��Ʋp|��<T~�i�Ry�VqjK�/J������9����]NH��+ϙ|ǫ��ю�):��I���|!��o5���\�g9��"��l�������Μ��!<���뜱��?��?�_����/ה��tJ'�������:�?i���˳��z��)��������+{�7]�֡!��y^��ui�����q����&�z��w��>��|~Q�?-��z��7c-��ci�u9H���}5����QۧWx�.ol���}'�f7vk~�����c}�O0��;{�ޑy�͕��͛�M��{+��������̌�&����m�8�N-Q�zߎ�%��|�E�h�5��6�$,hi&҉/ojk�o݉-�R��E�K��>;� �9��%��/��B���x��'q$y;��q�p����>'��A���<��w��������۴��P��]����u����`�Kޓ����������^�������'d�����zO^�=��}�w���>qw��,]WӾ��5/?{�u��Ts�u�O:w��r����^�/u�?V۷��}���~_Wo��+�_��{ͬ�6��ڟF5}�����c��׻{��^jN������[o�sN�<���s�o}(ߖ�޵'�������|���άw��[�:��+|�}�,B�9z��MU)%T������̹�m�W9z�ݽ;�d��=/}�^�˚�p|�۾}#��\���j����mK%[٦�^�l�oQ�9w�����!P��نzwC��N����l����R�FHLR45D�I�m�b�$T�i��$��m���dx܈r,�D�-��Gh�qa*1�c�e�hḏ�\�1uI%�I�4�T�JA%*[���4���Q7$����Q$�T�i���Kbj4��+u�Tr�d��J���,����ԋj(�F[�&*���+�c�?�]}xZ�$����[1Im&��LWBD���捩j�z��Tm��k���Y�
Ec#r�W,c���4����M����Z�����
��'�n�V7D�*r7��8նrZ���ĭ�-J^��m��2�ltbjZ�[cber����krj���#B�D�T�zf�=[+J�/F���V�i��*ӏULqF���n�"�m�!;"m+�����T��i%M-$�̒YP�����J�)_[ѼX�O���WĖ֤*�lrģ�n%[�&����*Q�[Y*n��?WIj�$r�ƙ�V��V�#u�;*�Fؤei�V��P�i!�B\VDEi2ƪm���i�Jډ ��mtTOW��pI&M-(ʭ��#A)p�5�tq(i����UkIU[�k+�hӷ5�H��줴v(�"���j�q�ؚ�6"���8$����n��%��Ih��UUji����JH��D���;KcI��5\m۔eTC��!_�Tkc�""w+�Ԓ*pu֛LybVԛ����%���%j���"�^؍�Hj�D�Q#���T�P�J�r��7JH��F4Z��3�J=rGJ�QW,���knK��sf��m��8�7bR�J���cRA��vCK����#r	QU��wm��X��W!%�bĥLEE�(X���eM��K�qĔ�+ph��*�ڧ�.��TZ�+���Ĝ�mmKA�J��rd��d�7��z�8�p��"NT�hn�*��)�p١]��kna"�m�V�"b ����Z��"��RK�X�I�]n%&*�u�\�7u):-�����\v�E��TO]��dB�tpJ��n�8����r;d����Ա֑^ɭ�rUdؘ�U)��ө�ԝ�ᥩcmW-�uĄl�kk��$[��\�Ɔ���]C�-�EUR8�ʙ�v�\E��I�B�ƷA_}��y��nn��-n4G�>���V�Q6�X��D���hw�j�#~��[��k�8q���쒹����Sr4��K�c|[o��F�DD���1i��v%a-l�S�V�č��������z��=i%+�VD��S�Iۑ:�X�[�#^eK���%��\ɲ$�X���ާj��l�	F+]��Ʋ9jvy�Si&Q�j����&�v��-5�&$���f�ֽ�{�y�
�+�W�t�f��;��vO��9�A�@��d6J�Z?����￵��-���S����y1�9����S�����ǽ���U�U꫊�mUz��U�W^Z��U�*��*��*���UWX���U|���U�[U^�U�*�U_-*���U�W����EUz�����Ux��Ҫ�E_ff/U\Ux���Uz�����U��	���>��@�m��Vڔl�e��1d܍�%Y�4L�&�&l�ZSj̭����[Sj�� ��Ow8l������|��mUx����[UU�Ҫ��UU�ҭ��V*��m*�V�U�*��*��*��*���U�+J��U]b��V�X�U�U�,UUX���U_-*���b�w�[UUu��������{����k��{�B�"�� ,X�ȋl���i63+b�d����72�X�l�	3S[3��fa	�V	�{ޝ������gUUTUUTUUTUUTUUu���\U�U��W\Ux�j�_<[U^�J��b�������\Ux�*��UUTUUu���[U�⯸*��*���Uz��K�v�UUZUW�Ҫ�EUUEW��g��jM�+6��&��y�il�� ���V��6�556��7P�}�����������*������*�꭪�U�U|���ZUW�ڪ��UW�ڪ�WU궪�U�mx��,UU�UW�ڪ�WmUz�UWQUU�*�qZUWʶ�V����ZUs31V*�꫊�\Ux�*��iZ>��T�T>*}��[V�8�[jնQ���C��7,������ؑL֊6�-oV[5m�Q���7�˜��ra�6��,��1�[�d��[�fQ����Eo,ܛ�g-^X��đ* HB��q���G�ڠ* @���������*ƿ��S�~D?$����������4�\a�G��"jNA(DN�4D�<pNP�|� �!BX�X��X�'O	�<i�4M<"h�	�xM4��8A(D���D�J,DN	M�N��0L4�	�$8'D�:P�"P�� �"��N	��['�"Y
��	�d�C����D�H'�DJ,�Oi������D���DM�� �A �8C�Q�5u�0h4�;ž┲�*%���m�G���!�d��� � �蚂s?��vd��7n4���㎒�k-Q�`"��G�	F�h�ċ�����jg	PXR%$+E�wvP��:�mTW"��4I�n܊	`��<BC,�lY׌�4���� O��*\"B��H��t�g5�|"�C�ǒ�Z�RWh�L�#�Hr$A�x�n�AYa�4ݵJ!dD�$B�Z,W.2CY��PQ8��2��y"t�MX��[��]5��w$E�I�C�S�9V��G"�ULCu�X�F!�R�L;�-��4-�V�"�5�,l�'ԉFR$Ə	�K��1�b�A̅v���l��&�L�ƋJT�U#����-�z��R���)F:�:L"�Qr���4D�M��Ph���G�v� �� �2�&J$!4�k�b��x��E ��B�R��`���Yq�4gC��>r-$���֍�7v7	���-V(��9��;kN���Ș�Y�rc�F��F�v������P�rlrɶ[+$���D���ԥ�W$��R��"x���ǫU�z��u�!�Y1��*�vFV����S�lhvA�j�eB���.T��� �n�iμ��^:T�N��-�kXF&7t��Kd��TKq$m�:���b�kdq��B-���8�,��Gg�j�=�(��ck�5N=u�h�T�ېpjԡ	 �Պb���8��+SI����5=���?j*��*����>�>��b���b��������> �b���b��������>>>V�W��*��*�������R�Z-l�������<��:��<xGN�_��ݭD;�\�ԋW�DI��r+`\Tv�A��
"�]&2�lPi�h��s�,�(ڶQ��nT)J�b���1��<c��S��+,�cq��bV��2'[�7%G�����"R2"J���8���r��O0c�����LP��N6�$R)"c*������FǬ�4Yð��O~�a��Wk|H���G�n�����f�2���
46��g�4���Q��+��ڗ6wHHh۽�ɮF��gG���a�TԆ��x�$s'F��g�.~���2؅r���[���L���dH�e��#y�|�;�L�6yq���T�D�&1�+�ߺeh�̺��`��:"&���i�<t�K�aA(�ƣ��bXĄ��"�I(P�2ۀ�G��LPٓ��Id(�v�I	!,΍|�R�P�B�ݼ,b6���檡
�%h�0ѸHBA�Bad�86�=��&'��p��T�b[�irZ�)5&����dm(���0Y�_�dx�$Pa�f����C�}�K��6�>�vQ>�n�ʙ��.�v�<F�̼ˍ8����:�8t�g���e䖤�T�V��XD�I�����I����G0��(i���?h��T���g�g��e4�kO�B�2�M2���~�:!ב:&񕖫�6����B9�&��fz�3�go�.�!!�;(a�SO-^lU�28���r��졦�aĕkȑ&��puD8���%I򼮬��hp�%��4�:"&������8C���HI��B,U��I$`󯙯�D�V�I�7�i��vt$5̫��۳Y�Q�!
n���m�B�q�lx�WXʲ$�-V]JDq�� Ŭ+UÕ�Q���<��#�H��/�6I44d�P��с�=I�p�V����U�V�W$K|��ǟV�fv9K�7\�ڍ��ܰ�<BHD�n^�yI��c�P2� ���(�UK��X��8�u���1_0���u���4M��&�C�K!���Wܒ�#�$�Ѷs��G��p���gOoh4T�XҤE!FA�E��!��l�(�(�ɚ�!eO!�ƉȲ�[T,K.��y��N$���*�n�%�E�O*(�֝�(*�(6�(�I�8�3e���WĒI#S5�ae G��IJ�H��*-,�8V�W�)��<}�I
7�h�v��VpӦ�&"�����IR�'���8ņ�{;��n^��^z�4�S�dj�U�O���셕�&땺;�6%��tDÑ�ٱ�f�<��ᳮ��dh����y��<����E�E�iJb�MtS�mlm�Đ�uX�����x�48u	�|��a,�f�xD舚&���><xGN�=��QA�H�����=�$�8��$�`u^a*��ʭ�fΚ)�K�\��M�I,rP�鹸�۠���`h��:	�fؕ�<�/Di������	^�D��?�d�V2::BR�j�;-��,B$w���%��~CtVa�¯�zW�_��1����$^�pÁeY�����R�a"�R�W�m�|�/�m����y扢t�i�<t�]�p��Ve�M�$�8g��w=����1�&1��&��E�>"�j@��%��S!HxR�I�M��J�9��~��4�a�{��Q<M)�$�cE�1.��F��#�V��f�i+FL�aUQ�Bqr�CCC��m�:V2�!��W��V@�j�lj�!��fWvV��$����-�[D�|~x<�i�gq� �4�x��'DD�4Oi,�w�Jϸ}VA���z�D��rE��$��<]�LLHM$���)�C�x�+�d�B8�F��$K��S*�c�JX��?!�*�
,=�ƸpЕ�5*��$�K�z#m�<Bţ<<�Sr��)����ؠ��ǐG��qWk�V����k)8i_+�[de�w���l��|�/2�O-m��μ��8�:�8�,�}�����+�H��k �Ij�ei�Qd��j��1�%F<(UV$�")+�C����K�4�P)
��Bc�!i:�h�Y��!�Q�#��,ĳ��C�RF(��{ ���ת��Z�r�-ʒ�dE���D4<H�ۨDQȩH����Hډf��UQ*qs�;B�ԓa�h �zr0l˷47�ԇjȲ��Y5 �sl����=�����5F�[�Bb2
2X8��%�1,��;τ���>}��D���ݪ��u7[�5�j��J��I*D�s�xV���I,�[�d�]@��D�l��,�A�]�����[HѕT��r��=Y�"�L��ҎJ34����q������<�μ�#��ӄ%_g�N���5
bŐQ$���
M���"�Yä$4[�J(8{Q0�*��Ea��@jERx��]���\>I2;
��=;��mc���{�Tl�:�<�&�ǩ���Mn!�Y��4�Q�V�-�MN���-N�{5S��m��0⼬+�i�EJ�$A��3��"��v<N�4�0� �ٶj���q>��C��/G��yI�b�a��eG���W��|��O��4�"�Ķ-�Y������ٴ����bKb-�Ke�^%���i��KO%��an�M����̖�/�S��ꓤ�k[�Դ�aM%[L?��?0����i����&�&+�u?%ul<�G�o?2��+ߓ�a�-?<�S�y-[�[N���%���R�Ŷť����b�cZ-�>FVŦ��irm�KL��ť[L|�NIl4��i�̝cIXK$[�̘�ش���ZZ��la,���2�--�-�g��vu��H�N��xm�;#	��o�Y-�'KdI��,Iҫ�$ꓪOu'j�q�u-*��E�V�KL�[FSϘ�y:�'f��屶1-��-��KckbӫĖ�KKy���[�켮�;�N��*^�_e�~d�H�D2C�%)Y׷\���Ʊ���Wɒ����ُ{�0����w�ْ�H����Vw��U��_O/%F�RO;;���:���J��?�=�ӰUt���j>�N*4j\�B��}�7�xF���k2U4S��α�/�����kf�3{���z���׋��N#������z��Iԟ	�/qQ^G9����(��Z��M|���C�i����{m�1�y������y��_k��������=_����w�5����;��!�v����=���~��򮢭���C�ݭ�����߿U�����������T�q������7www�U��|}�{���uZ~��������o9ϭAӮ����.�����<�4O	��D��x��atU�*������8>��Ksg�+I�ɒ��gF��dodzc�\k��YŝN��s6h�?,!��Y�0�+��c���ε�'�Q�,�'1��H�\dpyH����p�m���e"�m���2��I��,]Jmd�Q�/�qR��-
qX)�0��a�!� <��C��e"쁀�``[p����M5y�!H���!m� ȆH0��n2��	�� � �4��d~h��㲌J8%BT>eu�������u�\u�^-��\E��IRn4�0�0TT{P>;[.�wi�_��s,����$(M��8`�Խ�v�{�ItWHw�U�"�)� �ٍ5�H�M�Ef��I�\�CH���e�����U��B�#�On3e�s3��,HG�����:�rIa� i�ܤ����J7P�
�~�%a(	4��(�0��pS:B }B z�CA	cC�70L�%��*IUc�����`-���W�C�cƚ2ݖcRi�20�EC���ʎ�+k�10�VD�ȧ��6��.����y�yל=<���g	T�b�ST�I��ik��]5��ZZQ��(�ֵ�F= ���
'r�>��9�<E�C��q��#�ʊp�\�����e:�ǏK"d��`�Zē�tQ;Z�˒%$��Ш���|���`�x��[bD��H�HF�*N��"x�le�Lٗzԑ̠j }(���
z4�"�"x�D��p0��2q!P��W�\8����B%:��>�K�Қ�!�H'�^�J�I�8��D ;>h�D
B��_��c|XB>@�M6^��'G� H�!�&b9JUĨ>s���L֕JW�)@�ˈ4�h�Q�ԨZ��h�����f�M13�t!��x���Z;-m5m�u���CDh���Ze;��gq�6� ��õTSu%V��I	@i�`0˚Wc�H�&ݦWdG�Ӧ[G�2���~~[o4M�hi��(���Wo�E�}B�TTT�(=*Ut��*�����D´�?.T�ڮ�Dަ�MF���`� �Qq��FB����N"g��+�YD��^0@X|P��ЃgHɖ��md�8�� �&�����i�ꦌd�~2��`z���	�V!�+�3�b���EV�}� ��f�5o����<�7t�4�D�Yn�FD�|3t��'�� ��S�1tPxJ�`�e�f��$0����z~���$����0�hz}���4��!J�}�;D8�и��xA7A���J�-���z�vTs�$���G_2�.��oͼ�4DO	����4�gM�ߡ�>���VŖ��$f��O|EEEA"��M�E�L!�FQn0-�7^�a ��Xب�e���G��L*�QO%5Pb�Am�b�1�d|��0�~�yDUm�GR7���
#��Eo5��0�Com��Fꒇ�8b3��A�A�A���3�+��K$E"�H�aS)6��ң��e�GE[h�"4"(Y�
#���?Vb�PZ��C�_!�EV_Q�jA��>�Y
٘HT���F���� #21ZVO�M�U3QM!��*���8$�?�EU��n�n#�ɚb?h<ϓq��g�%d=o���B�`�a�CA�Cd ��	���6����1�%_�El��y�\eo����yמyǝ:��u�59*��1�a�eo�phb��BBI!����QQPHPeB�Xl���+u�p`x7B�H)P�֌�O�u��M e�K�\�f�1�ZH(9�.�%���10mi�#K,�MIe���!�Hm,��%Q�X;�@<0<D�R� p��ƒL+2��r?w���,���.孑���T!�$Cz�1�Z0J�z��"D�H�H�1/MÄ�u���(��Q�������4"l�Qe J;h60�|���<��C�|4GP�j�X��5T8B��r=>`b;I��	�͞#�[>o�e8�&t�8��i�F����Y�}gM�3_��8Jt.�I6��hu\�0�gK<���4DO	���~<t����=�`�r*1�V��V��DQeI�wtK6�)c�:�aE�,)
PS-x��["�PK2�#�X�x�h@��
B3M������m��,�T\'*�&푑��K)�*���8���ƄX�jI-X�!�5 �^c�8����@�o#���5�!)h�U����.F:+FL�28�QIP�Z�v%�_1��d�=BRe�lC�>���*$���>���G��� �ż�j��0�2�G]�̮�����WWd,ޛN����Bp$B_0����敊6I���a��ȉJڢ��%!C���Ӣ�Պ t ����5Jl�o�F�)S���8�Yӎ7�g�M���v�fT�tK��]L3����-�R���D�����-T��1���I	$��"q��1���fJC����D�r:�$(�����w�>�4����WM���ˬ�����yמyǝ:�-�)�"l����lB�~R3:��h����*�(����y*%�C�����: �I&��rA��n"+ʔѥaP��YC�Z�b���U^p����o��	�BH�� kf���#Ѡ�d݅�Zӑ�m����P�֓ש���q�Zc2�!.TA�u��H�i�S#dP��WR�����ЛSl`�Tp�P����|O���[� ah��TT�J��29||Bly��⃤�=���5$$?�MP6g8$$"�tA/����\�.�9s��D����<ˊ�*ʬ�h㬭����Έ��"xM4��ǎ������fedf�x����B�ʅB��1%�A�mp�S��3?jJ���Cx ���Ś)�#�L�A���c� ҅�����8cF��խ��l!�{���� NID�ň��A�RB2�$hMBY�b���_�〸bŁ��g����v���=��Q��K���<�D�C�0���X�2�����Y�懦CL
 L0�� Ha��P����8J�"T��kg���ڰҙ��v�ӿS�D.�eN��z7�|X�{Ƈ!�D:l���8d��GN��"xM4��ǈ�ٟ��g�Qr�7����Z]^F;=�c�08������.N9zn�8@!����j44��>�$eex@������o��2#*] �-*ے�1:�y$�0������L���!��[��V�WN����2A���:��T�˞	�Q��JP� Y�`:��w����Up�BBI����C�냾�X���< +)�aڇ��Z���YC`Q+T`�A �V��c�݁dfCP��y�J�T%ۀ��C���)���<�! 7 ����*��S�6Cd~F�b��+��ɤ�#I��U�ii�-�|��b�b���|�Yb�-�KL�ش��Z[ؒ��io1W����=���uN���q�-�-"ZDZU�	h�i2����Z>KF��ҷi�"өh�د#��ul-��o0��[�-<����>&I������'K:f�m�iiii��:�-L�+b��ؘ�Z-�-�[&�&#�|O����kD��&�a���~Ki��iiiձk[6����kb�)iim�kb�ȷ�\���D���8lk��='K�t�N�y�:���k�]Uuĺ��]RqIڝ\I�[��U�7W����8�*�)�؞c��:�]b���e��X��b��^e��mlZ[ؒ��io0��mlm+I���d]J�uI��]R���'��>�!���?���@��D�g?�����
2)�-�pj�]v�	ݲ��.���L�6*����Ө������1v��ظ��ws{ԗ^���c!�4z�o)H�����+,nDUq�H$��5�\�v��ܥ�t�E>U��a�v�n�YM�d⌆��h��v�A|�Fs����4�I۔X���|ܬT��X�I��dn���wn�5�# �&�Ѫ�Ś�	�P����V�'	2��uR�"��'Ɲ��;Ä�LH�:k4\���c3�d�+Lr,U�P�u#��5=&��!���#o�qߙũ�G����Xw�<O��o���h��_-�7���o���P�_x�5H1Ѹ��qs��1�(�yP⦜-��&���b6kDArHD��Ա�!�Cr5�¾�!�IE��ֈf�����>p�G�7�C��O=Ӊu�}��G>��{$v>��qi�g$���lHLn�_p��|�����5���cL�y�gvO�A�D�>7�����^#�V�C6�2�ro)��ۦ�|�ţ[�ɒQ�9���;/�����w�����ԝ�]�����=��꒽;���J�dr�^�Ϻ����i��d-}���>Z�iEh�-�G���J�k���mX�Y6;	%B7h���j#NEE�K��n�jRR�,VEP�F�)W�8�HY9YR��WJ��bz���6��TЊ��dqRBRD�I�X$�jҸ��CEUҋ�I�Y2����$!	�8FՕ�1����6E��eM��X�eר�٪9[��H�Վ���ĕq5(V�S��$'�*�!F���HR�bu4��v�V�7m�I�se� ��U����#9�o]�~�uZW��߿o���߮�����{���uZU_߷�����w������������~�߿e���ۻ�����mUz����2��)UӮ����.��km�u�p��x�����5�?��䲧�&�#�S�
Y�Q'R�EQ%kUlCR��0��+�c��r����@�Aѕ�BP�bb��*�)�@��wFȐ؆!�!�Q��86�c;�����bU6!���T7aej�뀑-n:�JA�di*��9V�ܱH��jF�ɬqGh���WM4�M.!k��BctcN	R�F�P��K](��Hh�g��F��ǃ�������rnL�����_�C�����f�3#C\�8�� ��V�y��T�UCB`|A�	ǅ�Н<�S!D{�ew�L:Ӳ�F���h�tw�#�LP�D�H<�1�(m���cd�,v��������!��d2f����o�D|��j6�8�yF1c�*���d�Gl�д5��q���~?ùs�3��a��t4x�ԪÝ�#�Z��<�<�-��~t�"h��CM!������a̦��[����1��Q���%<r<�FB��I!!A�2I>���|I8|���P|@<F��Eۂ��ɬp�H�.�Gᠲ)|29]<~��K�F��L��EUzC'J�� �r?7Ad�hkRBIm+g��+Fʺ�����c�jH7
��[`����Ui���k�C�<�˞� hˢVd=�8 P�����\n�d�CuT��*�N�<e�d́������h|�M�8@!P����I�!!uxS<|U�������D؝6Y��OM>mo<��<�Νu[�*ҷX���@�jd�#p�4J��d�f�7s��c�H����� }�*�3�p���61�9c������:A�԰�+c� 92<l�BX�R�Q.�Y^�&B(1�C{h@4@(�A�n�b�b?�1�/�Dh�lF��v7�����B���N{ב�n��,�����G�}���`;t�~��_�Vl�ձ��*���:}$��Ay���q�S�:=��WJ���T�V�>��ć�=����ͫ�������$���C�Va�ʺ�h�DuX���Z��U(�N ��X�l1:J��J|�ϛe��i���>[�g�DD�i��=�T
��L�gc�1����Jwј`Y�|Y��b��tD:J#��$4Dp�ξsFXa�VjՊ�ܑ��;��e�dlB:����K�V֩Vh!��Q��"JEm�٘A����l�A��2`L�x0H��d�@�h��)�I�l*�[FH�-8W�� @��c�=�(�	0��FG�p���*B�nՅ�O�*�r���8(tE:<��������й m������@b2�� P�6P����-�6���69`�|64@�Q��><`�����嶷�u�q�N��-�gw�����$5���*[�Ir�{*ějLd�!<�E�EYx�B�V��W=�gn��U���Ê,�bwY)Wy��d�ah\tDF��ѦZ�
�E�!�.vdFq�ð\]Wr���#+O"�
��*cl��,�����K$nR9T��(wn�ID���ui��U4�M4�1��G����NH�H; ���ƛ#��]D��B[qa�{�1�Ə�9%.��RP�9�Z��9�D�h�10�
 *'��plb}�<���7гOv��}Z��a�HY��|p�'�7$����'F���L�5TV���LD�T�=�s�3P!�6@�R�c��4<�CC�� ��Z]&��@ֶIYp<���<4�HB�K���:8t���%�% a�=�`{c	%$jY�u�"B��+khZ%	,�Y7��N��
�W��e�)(!�.Hn&`�P��WŔ�>�����~	(�Uh��%W������~y���k[μ��<��QŸ��1�7;֌��q�c�HP}
���\��}Pj6RŇ��!��%s�ݔ"�m��I��(Heu��%�έ�����?2�DzǊ���4l�vQ%QQl^Ok�X�}�Ģ p��Q�$�U@�A �5G�m�� �-�oz�m�d��A>I�1_a!R��ʀ@�ΰ�F���[O�	�ڢ�T�	��'`�2�,��1CKDJ51�=�������4�LMb����1���No�:�x��ی�4���;�1�	6�!_IG?@q*Uxź�c9�<ä#�}�U_qim-����~mkyׄO	���������%ѹ�F	�g��1����8|YF��	?bm62�1A1f�"�"��`�Z�i�I��j��օ����@�ݦ�17�d������I0'��5�����0b�ː�aT�5"ЯF���$xQ��P�a����`,0@���^�i�v��!�9��J)�Lg�����j�iu���'F��:h��k���{��!ǖmH�^�&]B���r���J6���h*U62%���yc��� չ�M#C���Ɵ�u�_�-����^y�t<xGJMADg#eq+-�n2P�a��MF1�c ��P�W�:Ob1��^�.�g��U��	mӆ��Y���Ic��a�b�2>�[��R�( ���^��N=�57w��I��\�Wi�=I��#:J8?'Z�2c
b<i����PU�)>� dXUJ�����>|P���#��wVY(���V�y�Rq8!����)VRcKa�����ҪW�.�9 x�#7ӻ�=�֟e�ow��&G�P��P���Hh|(���'�J�0���`:;�>v��(b�2�im?4������~DD�iӝ�!u�W%2�Q]j�[�zL�-!�1���h���kʞ��4h��f�k���
!c�8�[ېTݨV&Iq��^�PD[��Nc��*��
4��-d����7n�+iU���X�U�D'j�h��V��W]r4�+Hđ*ltJ��Q\T-!%�f}���1�`$oi	��4&"�4�H6�%MG5�cn't-ҍcR��όfp��a@gG� {a�c	8:�è�A���;$�!�5r�	��(�Bؒ%*4�h�=!|Rϫ!q��2�Xj����e������	�&�)�<�pX�`����t'H����Ѣu����j���g����%X�H}(��U��1�*�p, <$���2�U�K�u��!��$�Q�o�1Q��u��-����$$J˒���b���Q�d��� �2�	�lr�鐢�PQ��c��X<��i�UM!���9i���$q��y�����ͭo:��8�]������$�H)"C��L�c�@��_I�Vʀ\�P�1�����Eɢ��;`@��X�t`��tm��ף B97a���h(�$���E)h(>c�d(u��^pѪ\1�s<��L�c�pt�2�8#��<> Q�_�|dhvG/����:�Ϛ?��ۅ$��eQ�+Z�؄�Q(i�`,H��em�ᡧ��QV�C�C�45�@�A��Ns儈���Tdo����Johz[8��7>��T�$=�$7�5�ˢ���eفӣ�S4|o����Ç�#F!�(�8&h�M	�O�`���I��ӷ:'NDzN�ķ��-"ص�el�ZmlD���/y--���ka�i2�RK"�ڤꞜt�T����N+GH���-��|��Zah��U��R���6�%[�-���J����y--�[[[̺�M-����2�--�--������'����Q�~i���>KKE�R��[�ml6�NI��[�6�����X����I�-����KKKyl�<�#�0��lZZelZ[kg��='Hh�:>N��::'�IѬ'K�'Id�,�C�|i�~�!�WӉ})>���Rv�����iV�%��iĶ�e-�*�	�؞{3�u:�KK{�3���b׉��id�ش��/<����a�\�OI���ӥڥ���:�-"\�%�G��E��{�4�������BG�T��m��w�5��f�ߨ������LY˴=��$���N��K�cS��جޝ��W#��S���.R���:D���!�f�V�����l������fw����I�g>�f�y�)������}�9�|W�֩�w�]�ˆ���A>����/���⭪�V+������������[U^�W�33�7wwy���*ڪ�b�����������\Ux�.~�g��4�a�Ӯ�Z�Z�u�q�N��;�16X��vvM�1�c `NU�n�)���I��m��!��$����-�i��LT��Ғ%&�*����S5�+ȤR����$@���|��/�!`p"Fd�����q�������<Q���R�����!,��%�D�O�*RPY�kl�<@��l�D�6�(Ns✓Cr�E}drv,I�H.�'��2:ǣ�?t0t�H�*d-�D)�G@l%� e �]�[o���C?%Q!BL-W��L)���d>C�%>�u�G͢�y��Z�?-���^y�t��bcuLq�kTĠ�wY�"B���TTV���d6t��d�]]�M�U,����:�y)���w'�ګ��a��e�����&�.�zD5
�Qi+����/p��QSF�p`6Bȩ�zP0K2���m!�������)V�0B��S��F�CrL�l�������I[(�&�J` �0-�?�As!)��u;O�J�qpÍ:���+��D� � q��2�8Caѣ��!*���`��%����2���*�VNE0���j��V�ؤ��TS��G�Ϛq���ߛZ�u�q�N��T�~��&;��K�H��Hrm�\"z1i[T��٦��SY5�i&:Ī�Svz��4xʝ�9tT�$M@d��##�\�l"4׌b2�b�f;��QE�3uk�8��lS��8���X��sa%jFp�c����9]R��ĭ��#��(���M�հ;f�[HԷ%�?y�TTV�����Cf`�b��V�(ȬN��x�K$MZƬnIm�BK
�kAb���lɲ�n�B`���b���$�K����I MĢB}0;�M\08qM�9�CAd>��|�ႆ:,��:��A�q*d�1���=�ӽ<+H(8�i*J�2�s�(}:b�3+�L?1�Ƃ�&���	�t��Ho��Ue�N6��煹���!��utY	���FhcC�Z�`R�%�fz]O]�KH1��j�%�䌒��6Id��U4�Mx���I��?H�׌���두��
ov:h��6���;h�,��K!�%��o?6���ַV��<��Q��Ϥ��!�]ݨ�vj[��|���x49R��ĒI����Y+kdQW*��2��;~�,�BpqiY���"$d���6�j�et�0Cq�oYF��6biH&%�������p�`Y �)��e#��!��I-4`���!�3�d<��2��KBH�L9TP�zF�JlB��8P�"�h��èM�h�F��]�����$���?P9C>z�B6뾛��ve2��G�v%�R��a�q���]m�ߟ�Z���O	�����;w7JϦz���tϯ�(���n�5���А�J��I����c�x��,�p�Ģ�Oq�G���L��I<�Ώ,�m.f�$-��b�G�f���� ��:~3�^��&s�(�Y�]l�<7ʪ�t���yY
"D���R�x��RY*��J7ULʁM�K��x>z�ۮj���(!�8���Tܖt�!GX����n~w*�ݑ��I	�UJ4����H5�F�$
&둳9�V]�p;dfݍ�b@��8��i>�n�I�/���4'H`�C�qL�$�rg��FC?A��P�(�8C�?��6������q�N��;N#0H�%C���(���	�g�3�i��87	,���� AشY�m�(���б�%������,����Ȋ��q�
(.]�r��n�W�N.gKV�`����3f����a�a�,�����e��>�v1��Cc������6t6<�%M���a��zT���h���>)٢n29Q����HC���8���4�AYA���dс�d2FUQ�����,!�p��Nc���U`t�,Ï4�/ͼ���Z�[�8�]��.�6�I�n�\18"\Jkѡ�!�+YaZX� �]d5�����""��Ԛ���%�Y*��ws�)�i�'.UbD�R�a,�u����;
��dmTݵ�֥���EhHL�ku��+���32�HK���xC*�j2˖�U�LFiK�ZgC�����1);*v2pu�~;�uUF%Y�ۡ���VȫEy��u��c�����a 12:� c�% 遒xZ91	��2|���J���:Ct=�8�)�ӵ2SZ(,�N��M���e�N�B��Z!��6[��O}�33V<��?E�;���	q��d��`�! �n:X�YaD���	e�n%�%�G��v<�х�2ąa�����R���~8�0�`0Ye4`�.?8���-kykyǝ:�8�p5*B�yr��[#!�B��F�Qr���"���8���Б<l�� �� �CΜ�������,ɍM��q�W��B6r���-&J�Y_�h��x�%dpsca����Cc��yd!�v:p,��t��ET�L=6Np�xPB�v|Sc}O@��t		�D	����ڌѤ/NF�����%r�Vp�+ʥ�O�A�F�2ra�����UX~5AD�C�cc���a�!f�����/V��g
�H�Tw�w�ni��%񔠃JA�<S�:�~[�Z�Z�q�N��#)�#>ٙùh���	(J�����幔B�J6dr0(�&w�*Q"B2I�}_�m:q��wr%�Ì���Cn�p�cC��::,���z��dq	^��V��$�k���\�����	A	����qA�
� ��E�6�pJ���]h�zy!��>�$��y���IM����{d�VK)�]Yu�O�C�t���B��6��C���[�󲾩%J��a����
);	[��d1��cC�C����0y�:
.I�GCN���KSZi�c��2>[,8���[��o��Z�Z�p�t��|����,��8̭J��!c)YH@������А\THSap�!$��J�>��`�?
CL�:hr�4C�^+b��i �}��M��%	$\�_�:�~�`�;H�J���HI,u�1�Qc
$(7�ܹ{�-9t�����@'��'YS�Tv=�u#!���fvpM	D,��O�Í�u���/�M?�yÓ�g���� �B��_�s��pu��	"P�H�o	�b�j�Ta�|�J|�C���L:&��	�a�%cZE�il�f-�KKu�Z�:Ɩ�KKay�žb���^d��Z-x�b�a}��lm+��Y.J�"ҩ�'K�u%�'S�ڼOy4����L-%�[l-�KJ��y<�F��V����ŧ�i��Z<�[,��[�e�:�"�o1i�Ly-�--l-:���Ka��Œ�H���--��G�Ǒ���Z9%��ka���ii��Z[3i��h�ص�屴��4)��#gG�>>���������yl[�y���Lm[o�ehƒ�Il�̒�Č-�KD��K�N�:���[���uO���q-4�Ku���,[w��f���X����[--��[��KKqy���akċu�I�1�-����t�I�wT��:��t�!|X�����!}�f�Z�L�78���*��U]��?-�ǧ;N-[q���%�W7��d�u��!DjM�d��RM �]�J��ޗ���\��nQcj�#ǳ����WX���'��k�.�,���TX�8T�.�x�ƚ|���7vD�KTO��Y�lBP���M�q�ה�VHj*{i#��ߟ&}�L���1��HF�k��*�CB����3�G����	�����(����E�r�8�ZS�n�Kz6_�����Mi�DM۳F�㗃�܇G�ZW������!T�@;�<wK���4�Un!/�8��������A�Y�p�K��:����6�}�-y�X2�SK�4�!����Cqs�1f�D��B���+gh���j�}����s��J���OZ��Ã�}�3���g��"���SXͧ:��a��!GT��O6i�,�4��[n������^k.�s�5�yV�zFb�#=�7���o;��!���^<ya�'���
8pY��/��˝�3��N'.��f��܆�,7r獷�-8�!�un�n�ABr�CitMb7u%
���t�C�-9�(�|�b��\�g.jW}=��֕�_=y��jy��{��ߍ�[ﮛ;m��JK�z0�++&��!�(��y�i�:���'�}qn�]���ݻ��U=e�ڽ#�>L�������:�Ć���
2�$v�$H*[tdn�R)�6�c�NRѫK2�A����61�F�W��uM�Q�%*W�h�EI!��۩H�E�"F��h���Y'�����%������ɵ�zT�U��R�4�q\�n�:;���dN1���Q����(�n$�L�I1�(����uk�"J7$���`�H���S�%N�BlI}�kI��НL�V�ɺs���'�͇vp�����(�͕$��Z�ؠʝ)\��2�VI?���x�?����UqUⴹ����www���b���������������\Ux�.g��׻����߭U�W���~�~��4��i��i���ǎ�:zt�Ӈ�l����)ȷw&7�WS�֥�c������ej
�����I*`ڰe&1B��"� АUcLPph��<�8��THլ�����i�m̮DR��`��%���e-$��ƫ�J�]���co"n�r
r	�lErQ
B�\\�	e1����xp���D<��<�&LI��}	��2:�ۡ��>r;����	¨���Q(1��cp�.]��$�04C/G*���;KV���c��(��z�W/lW�h0���		P��:��
tCE`�C��!�'M65�B����$��h���#	����3?�SQ��֌Q	4$�%$�D���Iá!��:9w�w'�B<fa�&Q��֎����&ҕEj���`�Q�KiƖ��ߖ�ַ������g�ݲ�0��vֳ3��`Z�h�&���TTV����C�����`��l}���J���N즾$$���H$ �ʱ�átT��m"8�G���t�U�L�S��Q��4<}�%������urJ,�ӣ��a�@;e�K���WC�0��<��I�p���Z4UcnEh���L�i��i����$���HIi�{�?8z:���
`��gy'���)��J��$����Yb�e*Ir�o����I4փ!E�����O�Ϟq�ŭo-kqÎ#e���Y��g-��O[.���m������s�#C��2Oh�B���:G�0����p�H��b�2�p8L�0C�66d~0��v`B��F��1��ut�]�h᳙r�5�d�m�Б6iJ��R�87�3�B��g��� ��}��"�j���R����96��Y�d���u��0FL�p��8!cE12���}�	,�C�}���p���n��Ԟ��IUӈ�+R��u���>2q�~i����ϟ�~qk[�Z�88Cg�\�ȐlT2�goQQZ%B���$��,�]�X$$z��M�{u���g盯�-�i�h4D�{>L�rcLf"
D(�(�죒	��GI+�LfI�ڼ�q�i���E�3�������Tp��!?�ܾ�0m6l�/n��Lc>6ڛj��:C������z0��H�!��P��;x�:�G�А�kG���ScV�ԧ�l��<!����Cnƶs0���(Xp0d�4�M��ϟ�[�Z�Z��#��K����*�&��[�ySxNR��C,IЬB(&!�L��\f��N!�bq#T�� qb�%Ck4�h��5��6�Hq�6�v���r9��F���T��QѡNw�[�4�)q�5ƥ
�$�b%���BP�U����Ғemm"QT��i�˲HKL,��go�TTV���6=������$�1d�!Q�)!&�BIh��f��.t�b½t��Ⱥ�+�D�/n�XL;�L�x���Ē?�4 �`3.4�@�!W����w*��&� ���P�Q��>8L�`p�yU�p�S��f�!&*=�(]pt`~���]��l�����0��G�`��0��B%h�V�^W��b:<#�~�_��2cT�r��Rbte�+� ����g���.xό(������Ƅ��T<f�ĜJ����N��6Ӎ8�帷�����8��Į�!L��s;�/Qi�Ѯ�"���$4XWN=tx����G��O��t�Ad8zxpy�h��0��8X�!U����S��P��#������AZ'VǗ�V��0���Z>2���k;�!�"[&
�(�L�WV��"VZ���\ySi��!�L�4���t�h��eV�#�OWXy�ȏ�kZ�/�O��C���AD9����*|�էD�6h�(��i�u��?8���n8q�m���RRc!�=��QQZ,�xa�CU��&%s��j�R�YP��z>Lq�����Y����CF���^��ٰ�>5͆��B�*���:���߇X�W����˲+��B)KB&[UHK"�ث)W���vP����|Cf_�}x`�wFN�����Q%���zB������;4m�D8��$�T����Y��=6`~y	������U��ڔݐ�5�$Q?���ES������CF�F�y�����Ÿ��������jQj�J�®IRJ�[�J�����А��_h�o�I'�+lDE�RFXW���8cǕ����N�㲊�pCN舕X޵��T*J�Dۼ2�pt��O���<pY�TF�d�9B0� tp���2BS"N�ms�*|K,�r����!𝉓��j�4���B��1wx�.��y�����P]%GA�����c�B�!���#�V̘u��M��q�������F���8đ�r1/�uS5�qC6�x�U��e"BhS[�!�Ou��(��t�1j.("�\!�J��Q"�VX���+�Jֽ�ԑS2�"8C��$�8�ձ8RDĢ��x�ɒ��w�� �ɉ���m�2�o*P�X1R�ɐ��E�һ,(�N�yRĐ�!!S?�a!����t�A��BXoFO�=�(��Px/$Â
"���S�f�y�HI	�@��:�\�O��b�H�弫u���2򺮼�U���*��(�2XY;�0`���Lb� �e1�;��㑞fi��M��fƜS��,�Ť#�� �&�6��̹Urيb!21%1��N������2B�3�bJ��=|����:Q��_-�~qn8����q`�u3����d���ѩ���b0�lr�Z6���TTV��8sF�$$W���xV��Hj����-�Q,u�L6odeHV�V[Y�E�ҸW��� ���e�����l���>������,�6@�!�/+��GZ���脝:2B��'Hw3ں.Y��$���W�b��DĘ�!HU6������L�U�
��r�8��櫑'�͡��-*��?U���L3ݶ�u��Tv���귇�|��2�2�Ki�i��x""X���ŉ"A0DN��""xN�� � � �"Q\�0KN��xD�&��h�&��h�"h�x��'K8"u"'�H%�P�B"xDY4��ӂp����,�$4D��!�� ��pDO	�D�:ɧD�f%�P��,J#'�'�Ǐ+�l����ml������\[��n��֋[�<�4DD��N	�
AA��3'%{�������R��W����V��#�����^�߹׻����ڼ��|�=�}U��nt�>S�z�M���^? ���>�q��{�!�5s��M���꾼�3�n���ʜ��Ʊ���7f/)ǔW=�޷ nm�k�]y�j�Ώk��>�e�Ws�m�?x?oM��s߯����E���w�����������~����9��g����v�goﳹ�u���W���ng�g�������֪�U�[s3�~�������j��\U�3?g�������֪�U�[s3�~��HiF�e�:��[�-kyky�Gl�n��**+BB���a|�Ĳ�<u�H?��;�BP���8#����p���ג8�hj�~uL#Z��9U����oT0���4�>��H�Ib�X�c�I6%,�
�BH	����Lş�*�U/
]��aal�<=CIf�C���'�ԩ����e�Q����c�=a�n��]�]h��^�p��ݎW<���d2S��o����rd"��:gNg���d�Kx�߉C��D<Q�%�[N�<��-kyky�Gl���1�����ѯ}��!���.��	Y�a�e,ˀ����Hr�·P6CZ���Y1�L,��A����$"6��؛bCc�n��8`��)B9��A#�F����NLG�6X��,��:B����QUD��GS�<|�~3�xcM�Hm�CL�oC�����!FtC[���Y�μ0i�`�`!>����U1硷e��VX�I�y�|�$��d���m��4��?8�ַ���q�q�͊����ETdCX��d���Y���6��؈�% sl�E��a^�KCq�OD���I�v�J8� X@��y{9�b����G�, ��[e�ݘM�C���J8��je�1��I��D�J6��8�(�4��"!K]ɗk5;�"���$8kXGc�Wyd�;!ID<���EG(�U[+*P��j�*&+c��f��#����G�m�n�z�%c�Pl�7�%~���IU��t�.�
�i�q����ZRl�8b�U�)+ߺ$�h�m�ϤDLa�����y�u�+j��}*D0GE�$����ϸ40�d5(��Y��8h8~��|��,w�SwKKK4�'��NnV�֢��`�$d��._|d�xm��5��d�H?x*�)7�BI'%E.�e^m�L#�~e��N���8����qa�ܭ����y�1�1EU%vpz�C�B�͔ɠ���X`�{$�!��zI܍衁e����WW��������r�"4��2�2��#e�l�|��D��?q6K<�Ҿ+�*�q�V"�L9�F߫�b�`�u�]1g��s��;\�)a:���u$Z�h���1�hNA�
.�����Ĝh(�`�ߜ�D��Y�������$0����a�q*G��>ض���2|�>a�u�^[��8����qb��=�L;�0� ���5��*��p��iLi$*h�􊊊К�)5XT����eh6!3�6<z0v���ÎK��E��񇕗�t��+M�}��nA����Pe���)P<���lDR)�I"Cm��ʢ0�c�ʚ���x�TǕ߫�8¶�N6�䪐���Ҳe	X��&0l|�oB5! Ѩw�Ezffն0q����&������M�`��(��8�RFHtpp4>��4�a��/��q�n-����ON8C�l�ů ��8A��X���"���4<��T��68F�lj�sA��L�� Q�~A�Pa�C����s�U�\�tb�&BIɎ8J�r�<q�bA�Ɲ���J�
0���7�����$K$y�ߕ邏�G��U0������2;>16�s&��;�n��i�UΨ�J��qW�6�E>!���x���t�x�
4h�.�����Z�Z�q��kyP�a��e�5T�7H�T�ͻ�q$���ʆ�8RbHJ9#��A�TM&48K(���=#yX�X�F2ۺSuL׊$wDh��Bf��b�hB!H!��*�7r,H�ڛ���ƈ�Q؉Y[�"QZ1AR*�[j"G�������*�U�bV�-J��d&C-S���7��ۘIm�lpl��C����H�-m�4KZ�q4!���$�HHe�$z��#��|�}�	
�{��`Z#��9 `ǟKZ��	:p������Hlx��IDh�`Y��у]$��$^P�M���\q��
lmR�>2j�!!�p`�h�>>i_���oI�����$��'����8Ԅ"�Id�(�W%�\���ϳ���ـ�ǣ���ٓO��UP��讜mao2�m?<���n-kyky�Gm�Wah�Ja�a�BP��"���'��J��++U9	+F��z��52�x��`zV�)gT��w��VQea�U��WvIل�`p��>e���֌���bܙk,�`YF]��t:�S�,v�2/�Z���P���"(1�VQ�`�	U�W�A�G���V�%1e�
�Uӈ��F\Z����a�90PUQM��E��,����i���K~�!��L�\��+�n��G�Gi�^m�^[�mŭo-o8�8&�4*�c#/G<ݢ��T�T~:>4�.>��c|�Y
.����oW�ⸯ�Q�~z��0�bQ+'}�,�$ �rM�t�<.�c􇄡���uuD����&�X� ��	x4�BL�Cm�~�D F0������I��8v2i��7�Y���rKv_-�=\��a
�H�x}���6n�h�����r}\;��<0��y�^m���Ŷ�ַ���q�:3�/ߑ�xj�kX��bE���V�����p��B9]*�Ԭ�lh���5<�xkݻ�{�oc�E��Lf�,��7DU�7+#�"��s����{��1������QAnG��H`������>BީT��]�9_u*F�>m1=�𯂐����	RSАM�@2����	RA��1+�2�����w���2��{����˾NF��4�x������Q�L:X����dDD�4O �D�:"iB"'����,��AA:"%X�%��'N��<'�4�4M�xM4�8Q��"p���<X�$��0H"'�N�%���t� ���&��<X���DL�tD4DN��D�F	��bQBX�FO�At��G�`��<���[.�u�mku�x�ȵ�o�����O�"xzO�'(AA>����RϖH$��T��ֹr�\���n��������=3z���D����wr$%���a���s�L�J�:V�e���$T�{g.��X�+s�&�Q\n�{���$�K�_��izD��\�?�{N�r��y�n=O�%m]��=[�"\\6�C^ʜɩ1T�Y22�-H�AƆ��m���4��p��AT�"N���b$�5]�2}j#��	<Ly-I
�[7g]9��H�1si�]�b�pobz��T$�*RA�6�3B��u��e��WD,������i�ѯQ���n�ӺU��q��D�N���;}'r㌩�<�3�2}��ݰ�����X2p�Dm}���L��POJѪ`�;H$q#\$��Zi�ܢ��\t���չt�YsjOMs�4M�h�����;Xަ Y8��9���ΐl�Bp�2[bBߩtxh�cA�(&2�����E�Ac���%U!&��a7���!�-9����(���S�]O���|�����Wۖ������q�jK��s����^l��lxz���Ηʩt������7&m	8�O�'�z�p�D�Ԭ(�IKr�+H��܈��bNYH�j(�q�ԇQR��!+H�VJ&(2F�*"MVʪ��!J�D�ݙD�p��^j�v�'�F�vF�����T���!���G�4[e�qI�)Lm�47%�JV�n��1R�k�BV�$�|�n�2	��$5lm���
4YcN��I)a��M��ĤlhU�G*��+�hsPX]�r'����XC]��j�|eϰ�e�N]���ξw��֪�U�[s3�~�����~�J��[Us3?s�n������UW�ګ����M����~�J��[Us33��i(�K4鎺�ۋZ�Z�q��}rV�3Hx��+,���G%%uZ�`�;+ʨ�CyEc%B���M嬉��N��c	�⍢�+$�U ��!U�������X:&�P����%�T҉(�'+��5`&�6��m�\T���:�I$U)Y*�ĪuE*V��DՒ�l�P.��6��.�|v�QT!�H�!V�!\U�m;FI$(�cIKF�T�f#RI*Q2�2l�����x���l��><�~hc�$�gć?'��ei\ˮѳ櫱���cy�H"����n{><]��c<�!x�:��!;�M��F�F<m��Tl���U��~7���~Ʌ���$��ә�T]\�;��i l�>5͉���#+e��~�f%����-q�	�WnT�VY%�4�	���0��|Vݥ��6�lT�YTyϟ��Թ�½+�N��>q��[y帵�N-o-o8�����#"ͣ?<5(�Hu�(�����EEEhD�kV�%q˞��*�s���af�hxxķ��qq<Ԯ1�I��٠�j���I���D~�[-�����c����� >�_Y:yѶ�(���j������arIm[�˗�X���0$O���x��ټ�����UVT�ņ�t�z0�N��g��ߒK���2�ɣ⇡�	dY0�٧N'>�UXW�f�GXq�\e���qkuŭ��qa���H�D�EJ;��{﨨��	+�=��(���X�x��L<l��A��F�y�gJd%xs��=	F�������v�n>�2L.�A��[�B���W�jJç�G�{U�u��������"E�X\��Ϫ�� Qг��Á�H_L��lˣl��Z�}]̩qP���+j�vW*�PK�ŏ9��
h�2�2�-���?-�����u�q��[L�a���R=V��1�6��Q���D'��O,���0w��AE|IB�B(�)]Hp�24!B>�\�������(17��$�8q�4�:�6x1r��m�T�'䮜e����T*����l�9,,������4�g?�H��$qc�H�-��i8|v3a(w�Э���`h��7�zL4���!��l�A�h�ԄVxx��W]>0���h���|�ϙy���q�n������ќϷ�U���'�6%D=��H:���WԱ7�I�ՌTrҡQd�B\�ŕ���4L%�B�A	�c:���&�(�q���!3QQ�C�"�?�N�Z��$�c���=t�d�$�J��y*�qR��$�Sr$�"ALv�X��ثo��h���	�ܒn��je�`9p��(�Ȫ�B�b�ys�n�N$�Y����k!%e}[A����2��a'��������!a�V���!�a���>�כ�cY��fߑx3�����$d�Lx��|l8azD�$Hמ�*��
*2�����񌏆ߐ��L�gRB�����b�(���UbPj(Ab���Me�P0��Y
�{��"�E�l8$q��el���qkun-��xC�luW'FBJ���%{�EE����|���_tp6sϙ�Ѳ�V���L�#Gp;5�M�/W�!n�qI$�:$��C��Zd�m&WZI�UW>��_֤�}I>�`|�t���=���B�_LIl�UUm��"Q��Q�T�M�Q���
Uj�ŖH4�n�����Y�6�p����4��̏Hd��xi�pۆp�LL�����Q8�4mS�㗋n�m�i���l���q�n�ż��㮣�6��b{/�0���Υ��QQZ��O��J�y	 yIc���t0=��N��}1����jV�+�3��g���L����C�y����8�e�1�ʒJ��H"*HKmt��Fܪ����Y{�BI$�5F��X>c��-.�ۄ%��uɧa���ѡ�<Q*��MPl���N�		`v:4�IC��A�R�8C�C�H�eNM|e���̘r�4Q���[e��^q�n�ż��㮣�n���4#!$�H�c-|�Ѫ*��������$_�ehu���5EIR����Cg\�J7:�)�)�J�IV6+v2dd������-���6Xb�	�<5��|�tb@�a���$IcͦH�?�E��8y���̖>65�F��%2V�[w���?xJgr��m�� ��"%VI��.[4xr6�9*���	�I͆K�CgM&܅!e2Y��-�����[�[�:�8�l9%�s�ulDJ!�$*?֚�\��zcSwn]z���&X�(�Q�&:��TUR����l��c+��5\Z�Y\�E)rl|E-�9�%�3�kXDm�4�W�Y7������c\X��Q&�*N�U���pVW���J���i4�R�uԖ�{���B%��R�r೻��3z6�.̓%�E-�ZG"Q�(�qȱRd���LI$��A_N�)���3Vx~W�W�&�c��m�ؿ;~���o�K*��B��cHIfi[w*��"Gۭ�>GO<�^�:1��牔�����o��aҶ;>%�U�}x&|��-r�����z�c�]~��?�JO��MؑFRLW%PIZ'(�d��"���~���xឨ��U�Gi�\e��_�Z�Z�yky�]GXn�>�(��Τ����*jQL����**+B'���zW����!�+0��D�B@�9gI�F�I���&�UJ0nNd�Ae>s�a���4ߠ"D��f��l#	�/GoCop�Pg�w��Im"+�%�r���Ik��VG)AI�u	�&rǉ�G�Gk����h~g�}�B�Rߜ<ns�,�c����gd�a�ϛ{��6C%ş�4��p�0�h�DLD�B�DL�&���<tN���8%�AA<h�Ye�%�b'N�Ԟ�i�4O	�h�""i�<p�&�D������N�"i�"h��0L:`�D�L�<P�$�'�:"h�ɇD��X��P�%�P��� ��|�%<�4�<�ֶ^mu�\qku�x����4��6�έkZ�mo���ae�<x��ǖ���JyoN#���!� �����o�;����{fe��<��>�W}�y��/(��%��9���_c95����w�^%�K�,s�˨�S��ee��,�tמ��竚��~�6�gD�+ڎ��|�`���Y������;�=M�m�_6�����Lԙ6�2��p��;^�I9}]�w����;��
L%�?g;~�����5�=Jo{����u�{��j��w�8���Ͼ�t��V�'yG��ۯ`��ӗ��̼x3���}w���������V�\����������UW�ګ����M������*��iU���ߦ������U|���fc��M!�i4�L4�OǏ��K[�-o8��L��"RIٜ1�
�ўخ���*�r��᱒{�k8�
��\�*��0��U���с�����m���������}	T��18I	h��*��,���X�E2$���}��Y��{�8|N$���^����n��:|�AӐ��y
h8i=��l-�a���5[9(�s��$F���R��(�����OJ�&�X�,هO~qkukq��uci�q�REj@����RA[�D"ԙ(���^�EEEh�������{*�8S�GaLl�'
���cz=U�W��9&�74W�E�2o7u��6��k�#��٩�Su�X��������Ĩ\/$�d<p�v�A�C�f�!��<���i�i7����K�5�$��N�$2�`ېؘr}	�hw]�~M��OU�m>������]O�U}�	��n�?<$����Z��dˇ|41�Gn��|����/�8�8������|t��O�II�6丢JZ��i��X(,��)\�(ȱ����1(�
�R�ƣ!cu�J�����l�cYE"�]�k7r�NB��9U�NI[�V7q��$��(�%H�V[cĐ�x�)+�Y�����6�D�cJs �,JD��I�86��RX�Z�j�H���x5�rwa!�a�d��Jv�vlc��}��K�YQ�� o>Ӆ�|e��N�%LLU�Yq��]��ð����!���Ҋ�c���!��BCE41FH�馸H�?E���߃.��Z�<b��2�T��F��c,&!"�X�P��.���2ߑ��{��z2`��DV�Ea�,#,|�e֖���[�[�-o8��M�/�|��,�2`,�g�QQQZ2�GJY�+��*���I.Cl�����|d��l���;td6��(~xt�e�UK�v�<P�B�t8�2Y	|D�t�k98��Y<&���J�,R�d!(��1D�+H�v��M�	YO�t�>B^�H����k;o����|��>i͇Ct�߉+V�,���T�b|It�a�m>�d�+��gL<u��庵���󎺎����1���yt5�����+����&ʄ�+��/C.�.�M(\E3����/������Ȳ���6�2tv0��<��ǼYuw1o�������7�i�����A�U����67��"Yl#��x�a��ɉ���i���%��e�t�4?#��c��9	$!!49.#a���!!��zG��'F���|>o���m��+�Ӷ�y1����yռ���Z�yky�]GX�^�������]����O��2�kҹS$J�n޺�8�68�Y�3�?4���mtu�B&�R�n!RFZ�Kcp�����Drf�Y��,x~|��86h��\;L�2�d,���׃��5C�pd��9��B����é��r28m>J쓟��_�^�䑡-�Wﾁ ��7-���f�߈F�9K�Z����'�[K[��?-՝6zt������̛���d؊�$*KH��]��<zZ�����Ҭ�%�7��HX��	*��i�K#Ɔ7���B(��Q�K�d���8�8��[	�h��<В�"�b�m�UC��G �3rq1T8�9��V�2D�Q�T�+[�۷b��f2��Q�R�k��d��"�~��TTV�.hՏ+��!�24,��%�dm:aP�6]T.Q23n���d�����ࢡE%=�v�Hdc�?<�afH��s�a��c�6a�����O��J$�S��Ge����za�ې��|�7������ã��Ҍ��K��V��R�p���K�G,���f�.l!�j�t���$�sd�T�-�"X݊A�٢!,�qOG��R��p����p��:^��pzO=1�^y�庵���󎺎���y �R�B@�v(���g�b����U�U��
�Z��t�+<Mp00y����U
$h���LO������|�Ҫ���q$$���z:q��@��BM��Y�+Q�`zǂaHu�}�Q�j�U�!������E]���xU�������}q��OTa
���F���mQ���m�q���m�Ly?2��ߖ��ukm��ucd�6#"IA��$RT&T%T��=��TTV���U����Z<�	%�*T)������:pm��̄fM���9h�l9�XO���o'�O��JVZ�)(�mX���J!Y���}ri�K�]:+ɢL�c�kd.�kc�O&�W��Bb�2�fA$"_I �m@�#�z�!R�^'�>C�H���W��$�<i�[N2���~m�խ�ַ�u�u��ĩ�Ƥ��Z**+F�|_�I�J��a���,��>a&5ND6l=�4��%&L��g]�݂yr	2:�YQ���,D��k��]N�l�u���)��9N�����ǟ�8��5D�dlKǌ�}�P��'�!���3�HHp���g.`o������p]2~�I�+Ƽ�����zG��hlrdr�T��cE0v62��d�F�d��6^ɓ>&�:`�C���4N� �D��h��ӂpN	�� � �	�(K,D�K8"tN��D��4N	�xM4�8P��"`��DD�<P�$dK;�%�pDO	�0L�Ή�H`��DDM�"A4��'DMD�0��
Ģ�d>A� �D�H&G�y�|�u��ukum��� ��""xM:~:~:~:[��,�ǏY�Y���߹�s�ݴ6���t�Y؍������{�g�nso"�'8�C���_�Nݒ%u��<X����֞�,�{��yw�V���(ĵ�����Ż*RB���MZ����5#b��آD�̮FR{���3�qy����]�i���S��4B�jON��]�g���۩���%n�+��R ��ݱ�Aj~w��;��.&�2$���@ۢc0�Qb�)���G���Ɯ�k0_>�'�/�BQ�
�e,P8����y*Ж��˨{���mE"��������Ѣ��\)�,�����Dp��b8�j- �	�X�4����>{KA��̜�q:J�V�3k�a�Q��y�VmhQ�IN��ή�o8rz�7�+���z�2M�Ll5;Tu<��I�rŶHW�v�󆿸v��]c�I���7�r�9ɣ���q��s-f�� N�SI
�	"�]ё��M�V��)�2��Jd�$DY��ǐ�!.C5d?���y��\e$j1�"xC[É+$���8����D�X�[DQ�M��;95/���x�����ow��9��Iw�_�\d�sy˰��wi�~���,��{���g�y�K�o6q/�|�E�L$pU2-BU6��&�K���(�v�V�`�CQ9Z��!jE�T-m�im�KMm�ګf�]�l�*b-e�ZE�H�Œ°x��#V�ەUH�Es�ؑ��4�\@��q\zܬU�Sj\J\Q�)�2��T;1&�j���j�(�b�42������'���NV[Ci�&e�b%�����FUF��V�(����D^�ʚcHյ��:��aZR}y�ƴt�w"�"U#��I"'v�.��*�]���s��\�˯���ӟ�W���"����\��}������*��iU���񻻻���*��iU����ۻ����"���Us31�}���K4�L4ն�����k[�:�:�/�)���q��N��RD���D4P��U1�pc4�"�RCeU� ʱ��!v�EH�ܢ$u�7�+TiZێ�!EF�B).1dh���b�A",,�X�L��XWI�[R�Z&+���PD��v�Є�UHMEh�����\�n�.U���]�rS�**6�F�<d�QU#.LT�/o"-�eF�r픨$���M�(,_�Çn���*�|~��Q$��[l���3?׺��M�Zd4Bd���xk��(jm��,�N��������Nl8>�Hoz�Y$���7���ԕ��$��y?����
1KD���2�i�E�h��xs�p�R�]��D�?zT���^F^e���y�������k[�<#�$��P��#[���b"pC5�pօ|��Q8RV�I�!s��D>eU˼Qλ�������ꔴBI
��>�zHw	&l>�+g��WOEb�#U�+�¹G
�Y[��0p������&(7��F+!�d,�-+.ac��jr�k��!��1*��������2�^���#���gOԿ�s�l�`ɇ��&�D�ϛDH�Q6�ai�����6�����k[�:�:�+�k$�y			(�{[<-��`���ܕ'�s4<	���z}$��f��j:?I���΍���e�~���R<��������H����T��j�i�'RU*4�~��q�����d����c��$��;VDǏ��|pi7�p�JҮ��DI$Q��~������7,,��e˽��$�GOG Rp6ai�̼ӏ�ͭkuky����l{�J(���K;�$$$�9
=a���ס̕E˺�G�
!����UIcm40�BC!����eg��ٌ���T�IF( �<꼃QpjE#�hIrQEGC�\�*�1��b�6��_kH����8�C�}���I��y>~�`��❏�y3�j�<��c
Ѧ�$��O�e2�32Z˴W_��H�j��Zf�u�|�\e��~~mk[�[�8~>:x�� �}�T��UD�[m��Zw���b�$�D��.�:$)B":��A�y����5A��� �"�\�R�+*��# ��X���
-�&���+�bI	%�D��l�T���F�u[9l[�Z��SN(���h��px��!�j%�]�А��w5�f�
�
8"V(�m��ePy�y_*�H�������<Ĉ��u���u~�H��u�|a��'+�m�u�H���2v���=1���7^W�e��R빞�2⼩���=(�wI}4�lv�^���?�8En87D$)!J�!�Ŗ�%��F��J�PC&G��mT���/���r�t6�hr<d�Jj�c��>�lˈ��.��N���������[�:�:�,wsQ��h�q�d\�j�P���48%4�g���ʩ��|���Lˢ�l���a�u�=�o����n�x�G��C��~z�y �vw�j�Ԓ�����@�Ǟ$��d��t7�����r\PY&� K(�L� �c��8*%b�I+��&!!)�e$�e�eT�M�j���xQ��������$R
>�Z5D��9�h6����f�`rsړب �����k�Y�t��+-���[Ϳ-n�o-��㮣��>�J��MCX���А��				��2U*��[u$����f߰�a�C�!G�4=8��`<<C:/�8����ʩ�^,�
�[�����dWkhP���*BGJ�Hۓ��'�<<<(6s#�{�B�J!ww)����	4:(���	A��EbS
�Ur���l���VBN�Cm�����ʿ��ҋ�����:��O����~e�[i�^m�kukym��uq�y�I"D������*�7			�Z�}mK�]O8p�I<:97T�2HO����ףA�.�Ip�QH!�1� � \I$�BY�=
z�_a��PU���$��>�,tgE�����?K��[�����Q�U��9\�lu|gj]]���܏D����X�'T�R�:��HE��I ���6r<w���V�K��7�tb2�?2�/�<�Ϳ-n�o-��㧏�����ҍ���Z�ӵ�'J�6
jD��-�)q���lUȆ\�db-.Ab��]�D͈��q�����G�R�6��jr�UU������y�QE�ۼn��E��vZ⪦(���*V��["!��OL��d�"4���ݓbO�$$$%�9�J$��Kq"�h��E�b.G��:�cn�B����RbC�*p����>�;��]G�Be�L	��Ÿ��sª|��"ɷӦh��ˈ�h<M�^�!*Q(���{�5�Ca��Zp��h���x}�����a����I����E�(�b-��F+dthJ̪R���lm������<�_�xf�>d)>��t��-�[i�^mk[�[�mo8�녚Nh�_��T��$$$L��:+Þ�a��!��dUJGez�p-����	U(�$�l`Xe�4l����>V�J����͆Mq������~�ګ�~ƔCx��$-���SK��>�=oϟ��5�7	.M���q�R�&��èAfu,��}�$ftq6��B�=�@�o���0�l?4���Ϝ|�H�O#�<��D�B�B"pD���&��pN	�� �A%�e�&	8"xN�xO	�h�pM��4M4�8P��"`����x�	�,DN"iD��0�K�!B"pDD�:P�#R"<�vD�<'��&�����(���O�A<$,�D�DJ,��t�O��?(A(DN�4D��>y�ϖ�+0��,��q%�b��s��w�7�������|�sݬ�bJU��N����ݬj|�x�^;"^w_Y�j�$X�S��m��m/�ݫ�(�������>��x���,=U�ݝ�v{�\r����$}�6��K�%N|K��{�g���x���Է���>�����'�?uu�Tj���W���������w��e�8���w��^r��������u�D{z�ծ������l��o[�g��c�����j�|��9���ԤDY������~"���Us31������"���Us31�n���������U����������𪪨��fc���u�Yu�][kyn�o-��q�Q�;P����c2 ̥~�ca�
�g�Į�GF#+f�I=:�Q��E�Z��k���}_�?>�P�c��y\���X+%�D(�ױF�H�����O>�H�g䒽Xj�Wյ-ؐbhːɨ.�G�2m��<
�~\4:�2$�
Kj��ւ�
�c�Ea�0�?2�^i�^m�庵���y�]G\e���k���LV�c�I$�������I$�B>��68;Co����������ʰ���b$B8�Ɣi~���9! �CΓ�$���8��k��CN�J���SǛm��Ӷ���rIk�:d^��1�4=v��I%Va�|�t8`h]�8\Y�G�n�7����v��C�̺��u��������-�ut��7��%:�h��:'�6�o"5~Nl	Hs75�B'J,�uő�NpE����ɨJ�H�Jgu��� �Qq�Xǖ�k��*�j��-�jt����|�k3W�GS��W[BEJ8�*��n�Q֖����V�T�I�m�V�dZ�K�$�H+\K`$���*Dw�y�����ᢑdZԅp�	��#�T���������c�&�VOv�!�$!$�Ξ�a�&����q���ӠeΣ9㡞�It�RITCq���������l��t?p�����9f����`�c�h�������Jd�$�P�<�9�F�8�����3L�MIC�����[�ZAh1Xn�h��Q8�V["���"n���+��ӡp�V��&�H쯺}'Ȋ25��w�ʲ�#���.��6���Z�[�㮣�2�»
ē2CphBʃ"���q��dX����P#�-:㐳��`xc�J�D*���HS��@�X��[	6l�b!D�%ʴ�|�|d>�	J���||>�I#�$��z�Ѿ��d68G��'=w5�.J���k,�.Q��T�(�E.��/Nrl����Q��r�C��d��d����2�ǉ�N_�\<=�b"71rT�T;V�e�v�O#m2��Zuն��ykyg��N�<#�HS��ɍ�	<M!�M`$gz�I"�G�x4����Ɯ@�7��Kß�tB}�M��'���h�w�&���0���K���Yly�)-tE�]��K�K���{ěiM�ǏM���-�l�BX��#n1�9���rf�2v�#	$`�
��!��گ��_5*UQ0g�^�h�g��q��F�e�_�u���-o-o>q�Q�g/cr�1��/$������J�|�ԁ��^/�g��g��ի$iDDG��Ti�g���h$�LX�
A"�n�7O�w���(�®��v=M0:��5��C$d�ѡ�l��0u[�3)�$����UXq�?�Qgr�����t��4Y�$�n�i��T�A%H�zV�S���b1��Bf�8"�8e��u���ykynܟ:�8�.�O���L�[J�0J#�ġ�7Sz�r���Er�]��K �Eh#-��u�ېZ�V�B�`�c&Ҝ�$��o81!^!��f���n��,*7V�U$��*I%j#��o�����HX��F�eLHL��+�.E#����I$�iv9��cn���HDQ�JiR�8��dQ�݅��V�R<�-��M�p�����V��|3k���7H-�S��Z�]W{M��HI�B��v麺�/Kz8�x�фԓcҜ��M�Hd����-��jWB�|��������6�� ��[3�}�DK%��-!V:ƪ��lA�l�ԢMA'P�#\�I:��2s7�xϿg���h�B`���|�kŁ�t���\i�[����<����u�q�k�eCHH:�x�6��H�=v�;�rˉ'�������U�lg�w��N�������T�g�*<�=�10�ޗ[:ƕ��S�?���x|?{<;��A���H,Pm�A�TKR�)ZJ'Hg���\�N����I#�� L��U�Z��2B�2D��|29WYI5��}3&X�0�6�+e֟�~mo8��yn��\Ge�.����ap�B�
�P���I͝�ҥJ*�!�ɷе��8P�~5���ʞq��͘�J�[�n~��s9���>q������v�v���Ts\�HF��?~�h|fO|P>��/G��b?�4w�w��z�a$���$��?Oc>;����יi�`�$,�3<#��u>�U-[VՕn�.4�y�Yy��y���d��[�i�Q��La����#i
6���I!@�����ee]^��=;�w���>�@�F���&�H�)��HB4�up��Á�t������i�|�G1�G�|����06t�/�;��*��s�Y��Q!êbW�n�]�W��<�6�KW<������� c��m�x����i�$�	�~�%)UF�`\O�������s�G�ꠓ�?���$c�(� *�d3?��-)�6[xDT!���m���֚#-5-&�K&--E���MZb!iiiZZ֘��4E�ֈ�ML[Mi�KKH�i�ai�--Mih��5��Mh"-��LD֚#-54MD|sn4DLDD�-M�"&�"I��q�ƋI�iiih&��I&��m4ZR�h�h"H�Zi���ZD��)i4ZI4ZIiikI����$��I���đi����I��i$�KA$��4՛�ni���LZkBh$��$�%��I��-,�M<�ZI$�k%�Id����&�I%�I���H&H��I	$�$�i,�I	$�"�6��HI$��H�I%�I����L�6q��M$��I6�M,�I	$� ��iii4�I,�BI4�I�ВBI	$$�H�M$��4�HI&�I	i$��BI��%��I��M$�I!$��ii�I�I��BI	!ɳ�I	%�I	$�M��Ii%��KI���I��I-,�M,�I-&�M4��h� ���d�H���%�ĲM,�E�֑$ZZD��ZD�ih�$��Y&�id�I48�9�4��id�$���4�ZYI-6�MZZ-1D�EKM�ZH�RAi%��I-,�M��M,�K"idK"i$�R�&�,�MM����-��g�L#L�1�LF�4kh��hѐ���FF�h�dkf�m���5��lF�y�<4hѭ�k25�5�l�f�f�s�<�M��I,�M��4kl�6�1l�1m�M��!�g�fF��6F���dkl�fѭ�5�F�4o��g6ѡ�FF��M���[di�m�m�[b5�F�#LF��5��6Ѵdki�̍6�����4l��0��dka͑���F�٣M����F�؍F�hѴi��h�dh�4b5�[m�l�lѬh�dkf�m���5�F��b͡6г!6І��	�,hX!���cB�h[4,��1m�2�y��(�hi��d!��4!��������&d�6i��42kcMm�i�M6i��Y�ka6C&�M5�Ma������Mf&��d�4L�M�L&��L&�&���dm5��M�FMm5�L�bhi��l��l�bkf�l�ͦ�&�k2i��h�M�Y�[L��MfMh&ɲi���5��i���ɣM3Ma6LMlMfM6��q��i���FMa6L�[d�4ѓF��k&�̍ƓM8<�$�i��q��i�4&�l��i4�D�MM4�M�M&�h�i��M4�i6Y4�I�4�M4�i6Zi�M4�Mi�4�I�M4�M	��hM&�i6I��Mbh�i�4&�d�D�M&��i4�I��i�4�D�M&�M4�M�MM4M4�4�I�4��I�4�M4�i4&��&��k&��i���4�&�M&�i4��"h�ɢ"h��"&���#&�!!D"D#$B$B$B$M-"�h��M	�4H�$Z,��Ț$e�Ț4дmhZ"-�C�<��Ț$Z-D�dM""h�h�DHZ2�"�h[D��-	�"�dM	�&�"h�4Y	��#&�"h�H�YD�FY	�E�Ț"$Z6�j����H�HkB��h��K�L։E�4YB�ɢ4,��dM"�h�$Z-��hZ"��DY	�4,��-!4HMCZ-	�B#$Z���h�4D�4kF��h�y��H��h(ţMh�h�F�6�	�Mhi�"h�F�h��4К2К4Ѧ���4kBh�hMDѴЈMh����7�h�F�CMѦ��5�Z5��Ѧ��-5��&-5�%�-��"kKDAi�kMm�ih��F�a�{?c����~]=hSM	�����~�EP#66b���Ʃ3�i�o��{s�ƿ����/��_�9���?�������ÿ����w� 
�����g��8����G���'����D��������l��GU�s�l��������5�x����a���۳� ?���+���_��t��?���N��� TC�)BP?��	���c�~��,2��Q[@��5��0~O���?�!�����j����T�8���� T2���������m���+���HD��zs���D����s��i�k�ֹ�N�r�_��?,~�)��\� �����1?�7���E X�� ��� R"(�@Ъ ��j ��UT*(H� �b�;m�H$t���� ʻ�S��6�+	�@P�?���q����`���$�l���%�m�hZ6��H٘�!����>��w���������^g^���̏�w� ���[����?��i\�����'�Y}�m�����?I����������ʅ�����u�@m���O��.��w�3�?���}��?�?����d�O������O���P?����G�}���?����(
��H1���d������C�S�?����8�� a���T@�~���_�?����ƚ�?����?�+��J����lF�	����AGNV�d����~ e�_٠�⥿� D)���~ѱL��(cͥ����C�4����v)�P�y�?����o��r�8�>��?�=A )r�?���?o~_ܠ* ��fT�f#?�6�J~ۤ����?�_��<X�����@A��G캟�?���������|3���?����7�G�C�?!>

���~0ߪ"c�}����~�jVV��5555)Y���SV�Ԭ�E
�ejj��Օ�[SVիSV�Z�jV�Z�j(��jՔV���[V�իQZ�jmB�j(��[+R�j(��2����2��aY�)��mYE���V)�5b�AX�VVj̦յl�V+���VՊ�b�LVՊ�eb�X�V+��b�X�V)���b�X�V+��b�X�Q���R�(յ��+e���)YJe+)L�e�P�
P�
�++(��(��YE���e��Q�+j��+(����ښ�j)�+)Z�ڲ����VVԡJ��JjQ�mYYYYYMJ���ڲ���VVVVR�������������YB���ee�(R�[j�ڲ�eeej�Օ�+V)���ej�Օ�(�����B�Y�V�B�
)Z�յj�VP�P��B�[)Z�2��Z���Z�b�
�����++++V����YYYZ�eeej���Օ���VVVV��YZ��e5mYEj�j+(���
V��Vի+��VVVՔյejڵmZ��Z��X�Ejڲ��j�V��VSQL���R��JV���e5emZ��X�V(SV+��b�X�VV+��X���M�Պ1Z�2�F�V)��X�V)�+�+��[�[)�jVmX�Vj+�m[V�mMAX�+e������5V���V�SV��jՊ�+j�(�AX��+)FQ�+(�MAZ�P���+)�
�52��V+jڊթ��VV�EV�ի(�YJ+��V�EjթM���R�j(ղ�+)��P���M[VQ�(��ژ�SPVPVQEe5���X����
�b�(++5+��m[+��m[V+��b�X�Q���mEb�X�V+jڱE
�b�[+��b�X�V+��Y�R��5mF��څb�+R��jՕ��SVP�[V�R�)��+SVթ�P���5f��YX����R�څ+(��Z�ՔV�YEjjV�R�MB��EejjՔ���Jڅ(��)�+jjڶ��������[VVVVՕ����������VV���MYYYYB���ee
���YY[+++(�������Sj���L�P��A�)�V��(Q�
ڲ�B�2�L�L�P�SVS)���jՕ���Օ���ڲ�
5jڛV+�l�V(+�eb�X�PVSV+��b��b�X�V+��b�X�V(Պ�b�X�V+��b�X�VՕ��b�X��+R�[S(���Օ��)YJe+)[R��L�
P�jڔjVVVQ[VԬ���eb��(Ԭ�mEe�VQJڕ�)��B�)B�����R���emJ�J�)YF��eeeeeej���ڲ������YYYYB�������+(�����YY[el���ڲ�5b���)��ߗ����/��l��
�� *����I��������_����E�H���(��Fa��f ����Y���?��<�6���?�����s�S����s �k�~��PI���_�Fe%!������?�Rڸ�������?��?�S����BF���2A�~?��px�������"�G��#����Y�8A�?�#��|lԟ�%w�?�.��֦�O���������^?����R�F=���rE8P�^7�^