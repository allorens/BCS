BZh91AY&SY�Y���R߀`qc���"� ����bE_               �ֶ[[6�4	[l���1��$��D�Ym3kj���k2�cM����Z�M��mL��T�Օ��+6J�*"�"QR��E�t�h����Ҍ�)Z-�5��m*bkZ 
�fڡ�Md��jQ���l-�m &�V´ه�S����m�)�� �f��c�.� �A.�[f�
6��Gt�%Ck\ݶ��m�.5�Q#Y��[23-�5�T�m�5�2�M�ۼ  �<����cp    ="	� @uy͵}ؖ�m4:��`�ݺ����mC޻�zڠ�[w[-]q(*����s���k5S6��흾��5m�*J�l�+6�Ե�zR�* ����E)@2��y������Y�ϯ�@ ����>�E�d�eUs������^����_MQ���GU��/������;�� z�R���Kcl[f��+>}JT� {��|������ GU��G�
���o���(��t�ڟ} 4��n��� (�_y㮒�44���J)ѣ>��ux_C�י��@
�	���Ji��mMkZkB��򔔔�{������y��ڇ��y��z>�tP�;@J������A@>����vi@<��� �(__>�����{��@
���{�+Fg�l6��6�e�U*���JU$ nX��Ҁ���wm��������4Q7�� �����PzB�� ^��^v��Dt�ޞ�4 �{�_  ��>� 	�S[Y���T��Sk�*T���| >���Ƕ��j��3��(g}�=:�un� ���x��s��r��z �z��� -�[a6ՍfV�ZJ�_>��J� ܰ[�z �\�@��
���u9� q�p ��: ���v�}��x (��:ݴ-�jى��CK,����ʕ)E {��}�&V(���� z<׸U��vp ������O�E�����wu�� �����`h��V:R�fl}�)@�� � �\  �]r�:u�混����8�ӡ��e���� �v� �\�T�L,�,�!J��{�T�(��>�9э �ou�;��
�8h [���:s׀ {��c@����AΫ n�   �     ���R�#L !�&#  "��Ĕ�H      �~��R������    ��
IR� h   � ��R*j��z&�# �����T~�$�ڧ���S�oISC52I����������.]�����χ]���߀�����>u�3��}��0����^w��U���@������*AW�?����
���?��w���������U<`��*���� �����_�ʨ�/���������g�1����lc�<c�|c�1�c�q��3�c8�3�c�7M���l��1�����18��1�g�1�c�:g�1�g�1�ǆ3�c�1���1��c<c�1�c�1�c��1�v��1���63��1���1�c�M�c�l��3��x�0q��1�c�plg1�c�q�c���g�q�cxLc8�1�c618��q�c�1�g鱌c�c�q�c��q�g�1�g���q�c�c�zxc�3��3�c1�`�3�c8�3���=<c�{g1�8�1�gdOS�D�|eLe`aLa<a1�xȘʘ�8��¸��8�3�)�)��� � �(�"ccc(�(c
c*cv������ � �*c(�
c �(�"c*q�SGCG���Q�E�E��WI�q�q�q�q�q�q�1�1�q���A�T��q�q�1�1�q�<e�@��*c"c�*c
c �*cq�S��Q�T�D�T�T��f�A��T�D�D����A�A��E�Req�1�1�q�1�q�q�q�1�1�1��@�T�*c
c
c � � �
c�"c0�20�0�l	�#���)����!��8Ș�8�����8Ș�8��c"c*t�8ʘ�8ʘ�8Ș����C��Q�P���P��aq�1�q�1�1�q�1�1�1�1�1����
c(c"c � �"c
c
c*c��L``dN�S`N0&2�20�0&2&2�0&1�D�D�T�D�P�1�1�1�1�1�q�a	�q�q�q�q�q�1�q�q�q�q�;`1�q�zd`eLaLd`\aLb`eLe`e`\deed�q�q�q�;deL`LeeLaL`d&CGSCSSL`N00�2&022�0�0.0d1�q�q�1�|eL`eLadd�1�x�8�8ʸ�9D)������0c �*cc �*c�*c �cl������"� �(�(� � � �!2&0�0.2.0�2�028� �E�E�@1�a�@�T1�e\e\d�D�P�U�U� q�Ldq�f1�q�q�q�q�q�q�� �1�d\e`\`�`d �D1�8�c
c"� �2.22.0t�8��ʽ�!��� cȸ�� c(a\aa\e\d\a\laY�` ��T1�e��WW�@1�Le<aaC�
c�ʦ0����c
�(0�2c8�=�1�`�g�q�c��1��������1�c8��c�8�3��3��Lc3��8�3��ǎ3�c3�8���63��l�&3�c�0cL�1���1�q��q�`�q��g�q�g����cό�8�1�c1�v�0c3�o��1�g�q�`�N��q�g��g;g1��2c3�&160c3�����3�8Ì8�3�`�d�L`�:e���`�cx��8�3�c8�4�1��1�c8�3��c�1��3�c8�1��q�c�|c��c8�1�81���1�c8�3�cv�3�t�1��1�c4��1��8�3�c8�1�c8�l�8�3�v��1�1�c8�3�c��Oc�{g�1�`�1�c�c8�1�x�1�c�3�cM�c61���1�c�1�63�c�1�c��c�61�c�1�c�1�c��q�c�q�c�1���:c���3���3�c�n<q���q�c�1�g<1�g�<g�q�c�Ǐ�1�c�q�c�zq�c=����1��8���q�g�1�`�1�c��c�1��q�g�1��q�c�:����.��~o�������wμ�f{m��P�wfӟ<��Ƭ�
6���2���8%䪙��[�m#7�B�jF��������j�L$�kV5��l�����$Z{a@r��uj�p�L��;�n1l��9u�R��6&����ٮ�K�I:�t��4!ٵ�BY�Q�r��3km޲�1�^�+V���q��/	�,}���ݵb��j��@��'��:��_Y܀�P�۫0�m�׀�wn1�Kr���q���lf[�d:��ԕ��Զ��y5�n��+T,��q�yv���"�A>ř/��6[��[�y��v�����0������y픅Ap��B�B���7f�;�#��K��^]G�Ii
�!SY���d�gZ9oG�ע�T�ҔK�*l�S��h����(lFr��WO,��swe��0� ��b��������eLJ����@�dA�R��v��4�[4����Pm��p�n���tBpC��W��h�@�[��B�LHE�`�Zk+\�1n޳n���W.}��m�]0��)�RGwe�[n��6��5Nر LVEp�F�V����<�u��d�Ĭ��Z�sM���3n��6̘��9x�z5=Si-����U�ѵxx�=̫�b\@��&fc͚k��[)�Om�uB*@-q<�Д�h�Z�5��&rm�Ob�X��Ͷ�F�GSB;��;{(����=׎�X!F��}A�/t��^��d�/��9��У��e��Nf'W ʤH�A)ݼ��:���V6B�7sD���.�,͠��b�M7��Hͺ_ɠX��Q���X��lA�|`��{F�m�s2�	Sl���k7]���"#d�ِ:��P�����f�M�5TVF`�ï��
��K"S��ol�D4���9��uE.��1^�wQ�ɹM�V�� ��h�c"��&�����ܼ�H�xѣ� m�1me��
��hZ.�*GUlz��r*�58Uw�+�,�Q�I�Ä�e^�x�i(E*J��fh�m�!�Fj\ût1mE��.�P[qV��w=���;�R)��mĮ�b7iP�u�P9���t��C�]���4*��Ŵ�P)(��@Z�F�[J�[W)
�T{�T�km���L!+2��梅��e�e v�*�m^�����e^�tV&���Z�&�/w�,W���Å���S݁����[r��T��K����T��a-Z��y&��Bo[�t
���XdA<�w$�cktP�x�<�:4�[wyGQ�o�*��u>��K�[ZkrdW+Q�;piPͨա����7H
�[�m����i?c�	�����B�ũnҕ'�V���3Un���[�ь�Vm�㲸��A54��Χҍ����b�[��6�I�6+�!�V�ߵe��@E�56*��n�Q�\�_�M��1a�3��^���imE�,��a`x�ջX��d/H��,	"۫��0ѭ��e+��P)��U��X�5ld��ܺv�e�4�ǁ�ø�.�ٴ2!-��&��˹��[w�6Ӂ@�I=��І����-�df,zD����5�՘�Q���^��Oob�4De�cu�D�Սls��\OLb�KY���j���6u҉U[�u�eL�u^Z��q�3�;Ό��=���v8v��Z���jm�$�x�T9	P;��dy{
���V��f�8�3z�9H���㤔�$�#�B����t�
�pSj�O
4%���5���)�[��	��j��Q[�d�uz,8�檵W����������0�/��� �� ��:ZѦ"�� �Kf���u��A�e�����[�L`)ik/2]m�����r�GdCD.���x�ŀ���Em;��1��󈨢{EjQ�lo�f�^�wQVYkW[Qަ�b�u��m���Ef[�yLV��/2��I&n��݌ֳt��q��c(L���ƕAz�+uK����U��*+(;�E^�D%\����Ьhȶü��		P�w�h���^֍x���dj�VT�Ġ�p��I0���a//)f�yx�1a��bE�zCv��������>2�#��.��ot=n@��A���3X�c:w�Ŏ2�c�o�U#g#YE'jثj��7t%+^Q��(�-�Z��^�{�6�"�[u���F���P��ݑ1e,T^�W�,���崱��C<	��m�T~&i�����h�Cؕ$��b�mI�i�d-����0��;��&�j�X�5�U�I��W�¥����y��)��M팗b�P9�:d�%ı�i�eMYua��e���V]bx����!/j��!kJi��������2ɬ��G^[UZ�����Y�������Xr��;1�ǡ�\�Āu�LA[�d�l�;������NM�����zP���Rh�J+[Ѭ �.��Xۋ3j�;r��w�3[�FR�EU��{�L�y�1kH�T�*ho4]�Mi�Y,���6��7��F��4e`�Cy��K2�`n�7hK��Y���q�a�z�c�-���9q�eV�/׎h�)]�չ~��ۚ�bj�\iX�[%*�)��aP�֝�eI�z�<e�ꁢ$��ܦd�����;;��!F+`UJZ�G]y�Q5������Y�v�*�fz�ۼA�c���U+U�z�����d7�c8+)ӴvKA�-��3&�ʔ��vZU��T�7lh�H.�JY��03j�*F��j�S��K���Mr�+�&R�=7ui��+nrYȭ���!h��U�A�TQ;xDj�4�L���b���oӸc��D��*C1�Ou�UR�Rim4�u�L'rVJ�%cYn����Ղ�kז�[X��	}�3L9��a��-{��Ҩ}0��:���-0,�<t�@R��'r��U�H��ěGB�oaŋ-��I��R�GQ67V�V���QV������B�Ո�,�bq��ɗ��V��S��Ci*��؛Y�iB�3c7k���U�-��Y�z�Rt�i�UuL/Q�r�[\�\e^iF�u�:x�ë
�Y6�ϬV����\�1���f�����7=�d��)�Z�1�zv*�ה��N�3�[d\A�IehucwiK5�l!��:�����֖�HH�u�y�J=[l<0�*�%G��u�cK�R^����ëd1m�sA�t�Ư/e��:E�wR�P=&^����- f7wr�@
C7�M�r��v�m<g\Y�H�5�L��If%��X̳�N������Hbp�kdT���®����j�^�g*R�oP̐��/J��wQ��٘
��)I�������i�U5Ru!Ce1��iW���&Kpht�346چ��Rb��/m�[,����E�
U�Hw4��M��zӬ�A�%3�鹴�%�"���93��-k�c6�m+�7%'����D����.�A�
)�*\x�dm!cm��p0�������sai�+��SY�J��%� ���6��B�*�6틢�������ˀ:�M^��x�fЖ��?]��A��7, v�F��]�Lc��hI��sF�qL�H+��<���݅���CR���/,�i���U��ӉM�Ht��\x�o����ɀ����+��B�J ��c�*+�y.�����T6�`�M�A�r��� �n���C���"�ƴ�.�R#*�G�kn	��M	47��:q��Y��X��Q�y��˭�"n�e���7�Y5 �b��1ڱ�L���FI[�W+m�իL�>	*w����S0��b��E2R2�ie��n9C+[�AH���~�+C#D��Ь���]��xGMlE|M�M
�¨]o�Dy�,)�2��!	Ð���m ZR�]��iJ���W���u�2�dU)觺V�B*�_Agp�F�\�Sq^%�V��[�4�nd���-R�л�=�b�4��k2���T^ ��ۦ�ЀBkN�`[q��^hk��M,��5o�o�L�����i6nӭ�'KLQ����f�yY!z1]�nP&i�(1�`��A�ݦ%T`��B�Ս*AH{���+"��a:w��:�ZO �q'���a�n�Yv�`# ��Q�KN�2��S�[W2f����sc/4Q�(�*�ֶ&c8ʷt�<R�̲*'d;��^[4ۋ&Qc5Mf\V��h�>�{�_KǆF%6�b���;&�ĥ�Q<�i�ښ��U�C+lۂ�i���5�Q�%�x,|ݖ�k��K%Kw�'���y�PLf-���+ꕛ���pĭd��P*���/2mK�mV�m,��[inb-e���6ۦ�ͅLq\Z�5���Xm�٨��޸7���N��M�u�iT�%��ȩ��K'h����FZn�p��@J۰�V�x�J����V:�Hm;Z7�Q�*`�9�+�d��q�G2!t\�GbP*�ݤA(��+�V���Vț�s1)����*?S�K%�t0���e�}�jca5�����>5�n��9m�dE�.ho�2���u��܆�˼���:^�-�B��X��GSG�>�����u>�2�۹@]�,0�n�V镺c?�	�Shkc9��Kѣl^a���q�á��	�rݕl8�,j�G�bי����V��S'�kCwUڕ�4Ua-�ZӶ����\u�$��%ݛ�40TM���L�����ٛ1�iV��H�)b�t�����=������$ʷtpZ?i���e��_ԆS���#��KO%���2�QKmec̴���^=��bj��T�*���ʶ�%�V ��8��G4�+]RU��Ɋܫ�w���^�w��m%J-��j�Mՙ�*���h�w>�Mn��Z!YomX���H���4�,���0 u���u׎iR=��vRvh��MVs�;u�T�}Pl[i��*"h�,����f�x�r�%��:��k8�ܽmI����9�����EA��<"Z4̡Ta&H�ʔ�8Mm[K����B��/$O5hƕ�KAɏi�J�@�p���f`�.ejt��j�HnͧR��ʵl1%��#76�"3]�v.�@ظ��\v���7�KCv�A
]҇R����-��[CP�����غ��1�Y��{6P̶�C��_�cA�n��Cq卽�0�$��Y���P͠�2ֲ�w��0Hj�8�9�����k8c{�)���m��<z���\�@�k4�sD�ګQQ&ޢnz���B�L���
�ˆR>K�kU�����~�HK-��a��fS��V�z�Bf�$h��Mr���Ŭf=�!�	�pY��R�D՝u�*�u�m\�%�+!�\��� ����	 ������.RYÂ4V隞n�)U�X�HK5m#1����Gh+�d�v�g��NV��5^�ˀ;6�ЅK�Ќ{���9�hn\z�|A��B9ݻ��'I�f���n�ڈRf�I\�Q�j?��Z�GU|�����(��"sQHō.DU۩�0�9���c%���]���^�J%->Y�)KJ.I��%�Y���$���'���t���T�"�8�l`�v����3��ׯ�q(�U�d�2�[�v�h�*�싊�G{���&�N�%�t%�GYd���k+�ҡ�D't��/��%��zL'
%�n��B��Vad���l�:O{I�[���8L:�q����J�+����EeiH�9�2(&^������b0�PL�p��\D<��D�)I.	�G#�X���Ԯ��4�'�#�W@iO��n�5��w��9sF.k"�-��$�7���bI8�)�Ib��I(��2JN�����ꨎ��iE1FL�c�Y
��513pL�fYD��2Y<S�Vt�faXٷ�X�����K��f�wYF�M�t/�<f�8��	%��%u�j8��Jj�$��r��]�J��r=o��gplč�:M�:�$��Vw�f��x�CG3fi�I��w+)b��5�SI��Ԩ�ͫv�6yn%ǋ�>|��\�H�ھOۏuu,�?]ꕫ5K���/M�n�7n��
�u�)͓�!$�;
�	:K'a�B2�g,��[J�k]]6��ڊh̎�����2��G�d�V�Dz�=ڬVĦ �{x��9u逩Y���Ȕ]�	p����y���GrR�o�:���5*�����q��!S*!u�����|��T�K�mu�h��LE����%�È�+E����Fu��oL�J��N¬�=��#p�^�&P�8�ӺY�1\��fWtoG��" �ŀ���sW���V�qNYè�'o/2Ũ��[!ȃ��O5�WI�iF�庫vUNP�$uv�I��-Kv��R8�<�֕�9�
<M�t��ip�o�eB�Z=fa�b<���;
'�:�ӵ�OB��J#��D;�3(i8����9�o3�^�8�3�p�����c.�l�7˹L��2�Υ)8��j�J�Bɚm� �R=♐�:�&3	�e��:@i��FB��2L�|a]�7J[ߜ�]'jj����hҶ����Y���\G�Z:�H"�q+gp��̛9�2�6Y�]�͈��u��C'Zط��b@�]�vNF�ä�p�#��8�Død#\[d��G��)��չ�3,��K%#�n��,�8̲l�	���C����ڴ2�3"{����V�fs%LDPV�skJ}��9\D���&͢�S�,�,�ͦ��I4�$	m8���1k.�%ٽ3K'0�S%��A;�3��ҡH��2x�2Na��$2(Fv��ueB�l�wI���3-0U��"�@v>ڤ�KV�Km�đ�	
�!�R�2Ѻ�sz�.��I�"�%C.�͆ݞΡzy�E3��E�Y�9�hZ;�q�*���)�����R���|�U� �LmtԬ�v�u͌�f�H�^q��d^�>� ?��#�_|�'���[?���4~Vޱx������6�N�ͫ��Gj'�M�R&��mj�]@�f��f�x*!���{Q9���%�J`}��R1i�X{��.�}۸2��em+p3��Y�%�,w9�I묮�������N3\�:�Qݰyu�C
y�&Vq�.������~�yD��ӌ
��.a��vqh�3�!���M����Z�v���=�U�X��o~T�m1����e��c�#i\USw//2�50�
�(���6��L*��(�&c�SF��{m>��u�iΫ�޷Z:�Eh6u��D�0y|�1�u/L�����+�	ȣykjsGA�s#�ս׷��V{oc��C�M����6;d�9.��$gN>�4h|T�<U{z��1�R�-�dޕ�r��kT�wk���Nq��!$[m�J�X֌�9�QM�{ٹ-�YB�c�[�rQ�]�oZ�w\o��ٍ�h-Κ�aHӷ��M)�eKX��k���/\�3�b�U����j2��oc�]]4m>O:>TEڏ*\�gl{�q��4���yB�z��N�y� #i�(`��u���@�R]A툛�aѾ�P{�i�*�*[T_D�<Cˏ
ܹqքs9��WAy.�1�˕�L��1��K�Q;�NsWרot��G�tyE	�yN���eEy�󴳰Pו����,�ԅKHR�M�ɳ��]���Fi��[8X��n���/�&w7f��i���q��as���� ��:�I�V�&��j������T�e�Z�f�#n�lI��܆��긛=�/�L��s���FX��m�]�J��&��g.�G-ga�ho�Wa��sA���BQ�^�-����{��6�>v�����j�U�V���`�Dl�Z��S��J*�k�n��������[�|�p��7H��g�g&�;��)vG��Lر�JqET/:�VS����ݧo܏uE�]����#��]rC:[gk!A��R�xBm��B˽�ib|V��
s�֙�'w1_Čn��:1c�e���h{�w�z��4�v�EN�{�y����nA�]�k�� _q7�R�I�QZ)M�o��y�]����	�Hu����զ���}F�`,0 vQPWc�7]j]o�"��2L��H���'Q<
��|��r��ѻtoJ=>e��k������lm��Uu=ϏnE��wO\�j�9$)�Β�V��%7'0U��NX���Y}g���Y�i)7sorf�OxWfDJ�Ϲpr��*�^�f�-�&E3F��Q��6UՄ�/��ŋ1�&zщ6rߞ�e��A$ĲoY�zj�q?�(@�#�������v���OB<�������(���zU��En�!s2�Ur����d��ɂR	����;����6���.�e6V3+��Hbݖr�M�6��+���{�!Zv�J�8eu�x�ZL7�x��o�Ofl�d�wUSI�כ �ѝ_�(�C����H���{u�yy�v�[uY�R޸� α�H;\��|9:n�s]������Wf�Q�{ ���[�`�c��r���oY��An,-�ƭ+uYXd^�ۨ&�v �Jbj�R�C�u}�k��}�O��P,�N�
�+B}���֖���)��#��ټ�����'7�JY��/�����j�.U�Mr�JH�9���w�Z��Kgz�WwՎ���1�E����}��_c�;�7�����B�6!�l���5���a���+ s(��rjӫT���
=�x������8I̲z�f����{�\�]��ĮA�J�o��r�J1ǫ2��y}��QX��Q{ˢ������n�=�g�|d6��ǯ��9�{��O5Վ4W PD_3Hq|:�Tr�*A�MvMD����������M�z{Q��}�x#��6�(�jqi|_>{��ӑ(�ӳz�V�7�T���PL�ۡ�!�Z����c,̜g����U6;דA��u���Д���T�x��K)�=]���6w=���r�}��-��4N�KNv�4:A�]�I�Z����amY��9�n��Xk/uը��d����-�r�Ξ�͖�p�H��=���PЛS�3�v�ac����_����疥�G-8�Z�ĩ�+l�%n�.vu3���ק��;C��'����%!F�yc�f�R<���������*>�BR�o)��޻;{sq��0UN��kE��A&S���}�ŵ�Z����v�zmFd}��=Г6Ӿ�ƨ���{C�D�"ؕ�uE�/�B��n�+�5ť�������Y�yyL�	�{^F��ݮ��hu��*�v=r(bW�	�g��/�啕���`9�ؒ�.�(Q/d�u���0ZsK-WmM6nVG��٫!�A�0�p�a�˵�|v���(�-6o�u�L��c;�:�]��S�&m�I�J�Y���9���������R�L͗���ԏ]�=�X�?����2
fwT��u�Yf��WcY�����{iIB0���7�3���p�sF��gx̺�h���R����5�����b:�&����ɉ���hh5���R�N�r��%�	�{r�A��H����/=�X��Ä�嗔�h�{i)�.ݳ���M#G>���vΙ0�}�Vd3�o�P�#&�����]���3�݇p'��L���ǫ6M�Z���kkEy�E��ow<��T��{�ܚ�����{z3+W^���Ы�����t������Y��ֆPGe�Q�.��}:�a��.9�襵ۀ��蹘3]�I�z`i�����ծ��rϬ���pc�C��WM�6f��]�m������v7X����v	��4�
�&Wp�Fi;Z�.u�vR�OdGI޹����2�`6�� �Qm���W�[�Γ2�m�eQ�.$�[�sֆ�#jWpǳ7#��O����|`Y�2�5�t�&dN;��Us���i���qs
lْ���. �ͳlq�:՚%���;x
=������2�G��%qCb��Ii�ҭI�)�ut0ݛ�b��1��wy�/��4��yK:�y͆f^;D�بj�gh]�>\{�M�=��+�s���9�T�qgTi�k�^�ZƑs�4���V�__;�J�n�Olz��n�9�y���2�n�Tp�z�M`��E�a����o�s� �oroF���V_7�:��ʝy|EA�N�2KAkߏT��Rs��$��.빅����ʲ�����A.�;���m5�=����M�z�]�f%���J�(��ҝ�.��e]�^N��kD�GɎn�EX`:�+y�����jS`�ɽ@�.�ΨUw�P)�Q����
����U۽��#	G'>>*��s�z�[�9��+6�L���X��g�m2%��ˏF��@�Q�o�nņ�pPid4�r���2��y��c8�z_��:�s�X�N� +�f���@�&�	F-��K��*қ��;0nh�ₘ�u���]��c���R�&u��T�+<����Śŕ9f<��-��]�8j��|�RAsv��
��Y�F�9t�Gt+qT��5I�a�E�׊�hQ� ��*�U
�o_v����r[o`t[~E�^,k�Z��л6fc�a8vB�7S�����f]geq�4�Ӓj�x�`!;b|	�)º��K�ӂ��v�AeU`z�ƭ�wp���а`:�i���3�M�(�κ�}\Y�3;S���m�=Ò��ɡg�JV7q]n]�ȑ�\{��K��QB/+��-��w.��2xM��c��e��܆��o6�^��R�vt�{2�oN�ɽگ����ɩ��<w�.Ĩ*6⹸T����b>�m<�Y{},B�VM��&�·��K���g��=��E�<:ޞ}����3��ŗ�w/����c�j7{�=�\Q��ue�ڛN������`Pv�u.�"���W��.���`�4}"���7K���ﬨ(ǫ�w�`g.v5x�5��U�j�t�i;k0F���to5��3p����}�o}�����x0+��5R;�Am���,���Y�}���k*�Y���z���`̻n��7HCB�2��H��bу&`�d�78K���L���Vɒ]+�ۏ��S\�OF��N�puaw��+%.�`��I�t��9.n��љ)�sˎ�5������:OD^��;��*�1v���p�$sm�U<�갵�g��z�9���	�P�j��'ưf�ȷIK�Bd�zcȺn�ͽq�!� � �+nc�u��o4�5��5�kѴ��i�F=�k�5I%�^6�>�K�t�V4osR�t�IǛ�ҳb�\��΢�%��0�a�d�si>�2�#6��2�{0)����b/#z�j1�v��&ɗ�t�u2�����1:YÙp��n��D�{�Wy=Cن.<�+:�uN�\v��[�'b�M#Jk[Ș��h��e�/�Qe�L*�en�8P������7�w:)�ۖ%�'[&G3�G��˺���X�Q�>۪"h�i�^�-R�j�+�^�������z�ÉC���{w��K:f<kR�5���Ы���&����O�=��M
qL��TwPD�LѰM�R�:\�cj��$-�%l4 崋l�vQ=�&H�tjVn�I�!j8�b*����ĶvS��0�LU檝.�a�u��,���o�F��!�K;M`�dQ��G�Z�;0N�bQ]���������:n5��\T{�ok {ݕ{$��gwu�7��Em	i�l��5�Qלּ�Cz+ED��L�פ5���d��g	3�����a*3cmG�1]����n󓪝�M���A'��{�\}��)�.S{��(Wu5v�E����%"(����K�O�n٦)WA�V���nۨ`]B
��V1b�}݋._,��WF����tK���t=:��w�₣�7���3��N3�Q��C˃�a��h;�2�X$�ޡ;�7�#���`ø['�f#BYZ��1���l+�c�_K�ZB�0����A"e�z��{^��|����1f�%���nrƖQR�䷶Z���jU�Q@��ˏG	ۮ���}���,c�i�h�Y�Ƙ�l%�]�����q��s�"��j��O�F�d�n��ʭh÷���yV��;��:j]y)u��zZ�oS� x�G�^��88ݮ[΃ێ�I����.�M��Y]���\�:R\�lإ�_R�U�b�$��-<�{�����vި��8lT�e��7���T��Y*5z������8��\Տ���t'�4��}T8;���uN��m�h�^�PH��[(�*��P��敹�[��e�x�lq�1ۻ9��:�܆���(!�2�.gul!��+��Cym����=��SgB��]�������i^+��=Y6¸g1	Q�έs}��z�:sێ��l��}�]�̠t��U��"���z�P�r�b..��7Y��1�0u��:Z6������b�8bQ�;��}O�q̣ۗ��<��N�o�v�͎	Wm�%j)[�.�X�z�u�X�ӊJl���JN9��C.v�wI�v��������������������{�z��>�:@����A���9�z�y��>|����|��{ =���Ͳ3W����sj_����XuQ�P��;���}��
uY'�ހ=��F��rVm�{��N�1��8���>1�鯛�^�s�g<�;�'w�G�;d��Q���>�#o��s�pG'�����ӻ��� ��p~� ��� ��`]�����x���x=�l�r��l�9//a��$�w��v�ɣc��v_����!69��a��	�p~sz�:G��#�|�ط�~�����|>�{���;�O�!��g:�������u��D��Y�/�I9v��诶��)���@�5́�B~�0i�wK� ~8A]{F!�#M�Vl[~�5��%��G��rs�z�\3�=�2�yw�N��� b��W����;�W�F�yQ�� �p�* �����}�
�'������0S���i�
�=����������~��T���x���٣��-2�S��F!�/���	��W��سr���RL���l;�NH��S�"��}�m;�le��o-P�="������7�.hv�f>��ǆ��	W8�C�F�J��d�6����Z&+����m�t3������,�9��Ǳ�]�\
��ls` �H��6Q'��2�-<c����fL�l �GI�9���K��-6��M,[Dw��wl'*�sl��OLQ(o7>�u���L��89�r��F���e����)Q�8^XH�N.b}�Zޮ�=�F��`؜�q^�6"���g�qйw��[��9�p��6�Y��ԡ�U,]H��]1�C���d��>���A�lؾ
�sŚ�r\Œ�c�O;x�+Y���<SF�itY-��R�W��N]u����m\��w�*�S���գ���MJr���7�ϵ�w�-k�W��]��<!UEXy\E�r�������\�tYd�K�)�5��
w��o�Y���H�M��=��ԥ�SI1.�IE�o
��d��,vnާ�p�j�,�zs�>79uǚ�t��G����h���7��-���U��z��N=�zq��u׎�:뮽�뮺�뮺�㮺��]u����q�]q�]zu�]u�\u�^�u�]u�uק]u�]|u�]{u�]u��]u׷]g]u�]u�]g]u�^�u�]|u�u�]u�]u�u�]z{g���]u�uק]u�]u�]u��]u�]q�]zu�]u׮���ו��9��r^�k�z�|��,]4{.��yx����kZ&���{�S���[��jaVeɜ"�P:րU��H�Fb)�ݬ�uؔ�"^e��[�F�9SA���8�!��O����]��E���k;��#�b�u��r�wO=��/!̩�:�m^���q��=�Y�|���z�����Ғ$><rq��q̝�<��ȓ�7�y8i6o���h� �8b��>���ԩ�]t^��a�CJ)|٠������Q��r3w��]��=n6��1,\���S�,oHi`�M(2kJ�#�V���g��Q�8�4��]N�r=FYƬ쮂Y�
�aG�#�H[�y��%�ZݙN49�ӹf�#�z�w���Y)u����Et����³�@��E&�A��a|�f�I��>����Ü�Ʉv��k����9lʎ��ϡ"S�3�����6W6Ť��9��e'g4W���\p޽�[{թY����*@֍73��o���GW^�U|�wv�:����M�K�W�0>̧��B���Р�NA_�7y���:v
>�Z��.�q�GI[H��O-k��²]9\�n��<��њr뿝���z�g�r���,�j�f8������]u�]~:��]u�]|u�]{u�G^�u�_���8㮺���u�]u�]u��:뮺뮺�u�u�]u�_����]u�]q�]zu�]zu�]u�u�]u�uק]uק]u�]q��]u�����u�]u��:뮺뮿u㮺뮺���^:뮺�V���P4�P����cv4��{��-�\��m��������m�t�F��d�������5敤��6غ�}O��Qf��IT��v�\#���1VX�ٖ�9+Nr뭬6hZ�|��Ix�1�����`>Ʈ���xZjK�ƓΦ�U����\�ևr*��|�ݐ�y�<TU���׌��'3"^2I�B ��.��}]z^Z�}2c��"Ia.���v����\naei�U�Kf59]X���$��R�3��{е5�UQ�u��6�Z�� Fe�Z^�!��9�y�B����y�1m�xy��ek�4C"�k�9q�}�MP��Æ�؆rF⇒:��MH>��*6G�2�F;w}�^�O9Li���}:{[��5��R{�5귨,�DSYi>��^����<4�}�41�����H����',ӭ� �!�CI"��J��њ��l$� "����ɷW[ܕ�c�
��w[V�=�.dV\��V;X�F�OX�������<�!6m�Dir���	O;�D�E� ��Y��ݼ�j޲��8�靭(â���Q�sӣa&��Iq�J���5�P���^gOB�B8F�Rp=)ne�	k�'rr��c��:���P��:�ՠ�Z��ʮ����B�W>���b�g>:���D�U;Q�iGD��o����	�_pV�<�(عb
��ϥ��]ǵK���i�&��#� �	�O�g˅]<��f+��������q����]u�]~�κ뮺��]x뮺믎��~����u�]tu�]u�]u�G]u�]u�]tu�]u�]u�G]u�]u�_�����n�뮾::뮺뮿u㮺�n�뮾::뮽��oon�뮺룮�뮺뮺:뮺뮺룮��,�����g]��n-�nQչ�^�A;��qX��2c�`����,�ݾ����1�ɭ�XV�',�r���c:�;	c<,Y�H��:��/�zq���h�\�޿7t��/f�e�r�^���nK���b��#�g�;�Q�8�yk=����dM]���zkpX.�$�
Ȏ��A���#�*�}��%`j^	6ﭜκ5���4KN�=��6#�ő_T�{)s���q���Q�������S6�Wzщ������X��,C����P־�*W�U���j���jS2�,�Y���5,UV�d<3����ݙ�sXV+F�����R�pe�[f�d�析V�Y�C�u�^�&"͡��6E��XZ]�GT����N��Y�����E����N��|��������!�x�9YvEL®t�jr�I�.����5ykgwS���9\\ L���H�yIR�e��v�D�:�"�0t-�ۻ�q���0*:F�8�sx�z��<�J7;�tVk`���+��\��Ȋ���)�c�M�A��8X��Hּ�dg�^j��H���z�7ʮ$�m���!������o#���}X��UU��R:�~=�8?]u�]u�]tu�]u�]u��:뮺�8��:뮺�u�u�]u�]~��:뮺뮿]u�u�]u�_���뮺뮺�뮺믎��n�κ뮺뮺κ뮺�뮺��뮽=���ۮ�뮿]u�]u�]u�Y�]u�]u��뮺��^g�;ۛ�<�y����n(��j�ͥW�Y�%a�i�.v�el;Q�Մ��j\�&g6'i�R5XLV�,��gTU�#����mb۱���1�]ɗ�`�]Ma��!ϨvJk����x�Az�����[�X��&tl	�-,��|>��n"�锈޺��[|]�&��h��Ao\��(N�R��wh�J����\+l�=�jv�uc@էO�c�(�!c���L�mي����U�Rw^=��2<�{��nw��L٣u���u���kIj�ʗ��RB.1�G����S��آ�J��Z��XF�VY"��J�!nnV���/P�)��H��a����38��Q�wA�h��XMaP�W
��a�*F�3@��\n�er-�h4@|�_T���9[1�M��R�W#$�c����6��G��'M�5���&A4LIs�鵎zJt�Нʎ�\��e���`_]��֦st^R���V�W>ǡ��������=P)�yCS��m��v�����}X��e����hɘ���P&=������v̌�j���d��K4�
������[����Y��n��dAu�dԫ�6������	rWfwm�g����Ǐ�]u�]~:�:뮺뮿]u�]u�q�zq�]u�u׎�뮺���]u��]u�\u�^:뮺��]u㮺뮺�tu�]u�\u�^�u׎�뮺����]u�]q�]zu�u׷����^�q�]zu�]u㮺뮺�u�]zu�]u�u׎���`��W& �B!>�]�k/C�ʍF�6���&O���\�i�Z{;RҗVVV��EPP䶮[t3�7w��ek\�!{���Z��i���oɡ�0v0
�����c���XE�hV0vmq���Ip�Y[�m�j*�r�pMJ��y�N�`��OmN�E[������gN2�^��]]�ף:��Z����5�W$�P���c5P��|I�׍IT�5���a2�]�;���GrehEAO:���Ӵ;�B�J�} �n�dswk6��>�������� �⌬cu�`U>]�����V�M<�g�T''	�g�p	aF���s�3E��S�虐���9u�b��:��N��%��p���.��������ۻ*���v-Uq��FnU�^w'�j�;F�g�Ϻ]�̚F��dR���=aX��o#�D�;�^۷y�j�1�������
TW�����8����v�5�{ʴ�7��{���d�)p(�hlyE��������O�s%�% ����h��q�h�P��!&�V�2[97�z�J�fk�b��@H8%V������̲���Z�s�j� v;͏h�s,ɋ�V|A�Anaq}���2�q]�i�G�fp�}!��«7�1L��z%.��F���|:���;������~��뮺�㮺�Ӯ�뮸�뮺��q�u��]u��]u�_u�^�u�]u��]u��]u׷]u�_u�^�u�]u�]g]u�]u��u�^�u�]u�G]u�]u�㮼u�^:������^�u�]|u�]u��]u��]u�]|u��]|u�]u�ו�����z<��UAj���
�ibR��7W��pe����v�9�"]4Bn��Y�#��R�f֑��_-�� ®Sz���h=;����:yZR�.���[�7�F��I܉Y�;S�/�B�`ˊ��R$��L�k4���g1wI���Iܤ
�ZU}D}_p����(,�_o};m�u��F���A�c̴��T���%E��;���Y�ܡM�x����nb'M�-�ͺ=��WMDټ;�zX!Vsv��&�Ŋ\�kq�]&����C0���Od��x�Ǵ@8&��oa�e��q0ݻ�\���c2�_hՙ��!- D�.y8�g
�R�,�+F�{�vk9���,�ln�jtpM�pd�N}3e�O4��.����Wvť�9�(b����#ԝJ�U���+��Wk'1�=���C_V4�G}GK��I2X-p��#|;��=�\e��9�믾�>rX�tp��0�(ꦆQ�a����r5,b��E<���O�<���OFv�yI�**�k�m7}��.i�0p��Fn�r'��6f��n�Ww��lI�AowM�������̧�e�ӭ�n#ж﷕V,���p��z�L�V����pib6]:	��N'WU��f�����2�d�a��R�7�N�J��Wh�<�G��o�B�b�[Y��I}��Xm���$�=�W�1�e˝YKNu���������Rԋ�R�,���I��0&1kD�C�Y;;����T85�o@�L8�#�^C�Sn.W�Ɍ𵸪�r���4�"��X�&�|
ݥ�����Lz��J���I�@�c���r̸7��5�z���:�G�Y�U��Ier�:�{\���!Ź�z��+
�{��tb���܋��i�9��]zʵ̖�[�{��M��Qqˡ&3��ݚPݗv�,�������LWX�yԥJ�cn��9f�Ӛ�*�����ld�����p�θ��Tcf�G&a�k�Z���J�Kk��R�vd�I�{tA�]� �����u[�N0��Ղ���� ]ݑ��@�ls�4^��1=�}%���b��� 1��N�����p1�\tm�s��W+~��?���(�z��)pj6�$;��]y����od8Fѥ0NK쥶/#���G�I�Sc���fø��M�Ԏ��~�5�X�9$�0���8�LŽG
�Ƴz�X�n��T ʊʻ���\�|��G_��oNN!����5���7Z��XL�X��x�P��*��o��fI��ș�F��l���*��	U�u�1��8J��Q�쭒�A\hY�c�o{x�Ӡ�DqV
��w*�¤�1��zXRl����Ц�=�:.���A*fc�d3n=i�ָ�>y��V�1ٍ�49��D},of"��o敭}���6FL�d��OL�v���><���te].��H�{V)�%
�9�b�*��v
�d�G�@���8�3���,�"�5fj���Z՝�g$�T�軈ECS��cRcy�6?%qg�崳w�]�yF>��=5
����j�e���m������,�n=�r��^�/wWˍڛ�u;��ɍq:�׮00T��W�;_��B6�EYՏV.��[�婇na�:t�ox����r���-�¬�;eKF�.�,*��B���%sQ������{&�ޓ;��ra��b�5*�k�]�C��X&ܩ&�ҼF���x-��]jf���d���j�6(����n_)M^eLX�QM5ύ,����@�� �af��q���׻��;O���)J����5�S,���ݘ�wcǚ�j�Q8��+uV���(��P�}-�Kue�Y+Re���u�$�
�UUʆi����6�,_2i��g��+4Z���h�Yy�^|ts5��űΧ�����A�D�KX�N��AA�t>��2�pؕpYvG-��z(��PϮ�s�]��Q.����^88��CI�;ᤳ%�\��w�P�ĺ�OP��	\Z��_b,Ҩ|���B�[��M��,CC8� ��H<.X[��n��b��ش6bH��q���#�s{L�cHV�*�2��ک�ʾ��.�nvfp��Q���/9�1�6X���t�Nc�����Vp�q��ipMb�|X%��Ǵ��dSjhvZ[�q�Y�)��U*�B�F�ʶwt��}��ƞ}y�:an��9�8�6��NW_L�3v��\��f":n�hK��7U���3c�e����,0���2DW�x�Vu+�2���5����W]��9�Kl(���ۯj$Uw4��3f�/��fwZ=�:h�I)W������AW�)�__������M�Z�O���o�w���s��{%�ٝ �*N����n��rƞZit%���r:�v�]Sf�YK���-JM�ii&e���W���i6��-���hlA�#n��Z�it�؃c�ݣ5����p�՗fL\bK'	�u�in+��ͦ�]�u�d���v�el����x�	����^�f���u�,%e�6�r%e����s�y�KV������1�^�H�CYM5�YkY�lK�$a&L�X�h�4�����#s�Gd�B�\h嫶�XE�s�2̣έ�Ia)1c�J�Ά���Vťm��JY0��v���|'��,���tc��!ek"3:�:�\h�0�]�������m2�.%�$�jE��_Ӻ8j��NN�xY�cr;��voaΟ?�����KU���eIvu�Y�M#o|�v$3JG�4��G�d�.F&!�wlʹ\�܄z�(�&i�����l�=���=�zmJ6W*MN޶&�ˮ��C���]��6�YXMͽU��N�+v�΢��x���M���G�Ӄ�1�t݉�g4-�[���J�&����=���8n�#�-�'�XO���/찋w��Ī�3!�r�L�Y9L�μe��޸���P�&�y*SCV��k�H;���Cq3}�yy9b}�"=Ž�[m#z��	��XEt�}4�� ���BqLa�#�w�T�Xt�M��6WEF��s�Q�7۾h�c24�`ސ�nu������<���:��.��5�D�1g�	7�7d���-��_h[���6.oq,[��W=�e�zƩh�q�`�R���%_{��]a�V
}�4ȹCvh��
���с^}ww@T�}��&z�q��˭Ɣ|�+V5}�v��ki.����qB�a
)W]DM��mJT�<���f���z�&f5DY�Rb�ҥLA6�A�&6��)md�hi��af���<�Ye#�Y5c���fY̫�V:"4�͋*�9���cY��$�lGӬ#"�\�3++Knљ�b�k3)16��Mb�+vؑ4v�cv�lVenЅ��4kV�-��ӭmR�릶�Xj�;cm%&l�l����]��a��b�nT�l1��f��kE�
�խ�e��ci%�7-3�tĹFEan}3�,a┲WI3v�6�0�f%�\�mn�d�]&�p�t�v���i5�m�3�ɩ�m�cf���e̵�Y�����bǧMKca#��:��ۤ&�����iZ�Wj�١U�b�&�gk*k.l�ԙ�lոu�l%�m��goO���)#dd��t�f�f�.�� �s��Z�Y��4������i��͇�<K�Z�[��M������@�X�6LKj�%�l̫K%t�v�陙Y��$��e�ŚIu��L�:Ԇj�eSQ�j���ce�ͳ�j�k.'f�6�#[3��y�̰ոv��JF������{fդ��\��M6+2�hB�깙J��LM���6�fԕ��n��#"�\�3l�R[�fe���$�k�fcl�i��ҋ\�DF�ٱe\�)��l�9�R"B�٫,�r�&��Fda���et��IV���%���u��
]4�t���b[v���������Ω�VB�F+��R�%i=��"�wn��_���]C]u����t�O'���p�M��ǫ��֥�!�'9Y�b���5��wM����U�;�w�٥^8��㏏������5�_C�pD�!T��KʁNH�#M4D�r����8#���"�G��܏-���p/D �)��@G'����8���eJI�1�EQT�Zœ��ͭ�������uJ'L�E����qs�����y�]�}}{~>>>>?���k���QATt^�FHN��E�s:I�3\��f-9�xQ�'�Y�k9׉z˗�y|�\�߻�n��y�w������r������.�rB�t�"ƵE�!�~��K�ӑμ2�z�z�|���n��___Gџ__^�\���޻��O,�$?H"�O�z�x�ދ*H�γ�/C�w��gG ���__��������u+:�"B�b�ȑ�E#��Ku8�cY$$"�*���}���Vέ���Z�Od�QQ�	�U�d	䕄~�yZ��V��w�	Q�ExQ�DH�Č�V$Ey��ʨ�('<��}���%��Ɗ�L*��$T�0�#���(�����y�q���OoU��UY)j��	�6g3�&G+Icum������ya��5UWz�یm(ͰT[�%�1�a
Y�k�|����k�>���q�,Dվ6�.𝮉�^�I:�pZs�eJ��'>��0헦�f�s�F��"��b�k��e�gbiF�78k�;:l��m�BZ���6b����k �V�`F�f�k�^jΞ(�p��K�Xm4t���J��cZK�m��f�[i�ѥ��f�[��Yq�j[�G|8?��_� �Q~I���\X�KER�am*Ȑ���2�������⽚n��g����O,f��Yjr����o#s���g��2��_/Pʹ��m@�Z|�V��AS�=�]3�Q��E[�����GU�o}�@6��z5	��t�ޝr�����geox���X�����H���P����)z�-�{���9�V�r�s���<����y�0���.�ք�O� ��m�`"_xZǛZ�����}ȕ�Uޭ���m�� �]����>��޷7��N^�Z�}�7��~�>�f϶Gf�P'���՛����2�S�Y�N�v�b}�,/}���S����9�gz/nI�/_ݦ�7+�:h�q�,��u�P�E!���ט>e�M[��_���:���6�{>�I揳�eן�&xu�����{��vx^}k=���5�N%~�s<���߫z��^�=�bv�շʲ����q��O�TƄ�ָY�[�*;���y3y���/�H3��.6�� W��30��eNބ'7/y��|���f�]x9��t�bSɓB��Wj�%�����+�L����y���\d�OU>�8 �{*��~kg����/��+�'���`���(i�^�"*+�+�חh�}�1,{~I�^��w�]�mN�U]_q�B
[B�@>��ϧ�x{����w�u>��ޮ뤍�W<y�~���Z�F��!]�Q��`�����w�����)��/�dD/�V���+7���w�C_�m�Uݽ�+�iK;�`\j|7�fvy6�/��5}C ߫�$���.���+{�=����b�SQ��P(`%�0z�V���D�n5��p?/�]7���s��Ş]���(���k�����y�T�C�$���p��]��Q��ޒ<���nW���c�/m���ׯ�߳,zˆ�h�q��s��朖��zﳮ��w�XL��w�Y��oެ�\?y��wذa�x<��҂T�sUp��wE�ڑ��άF���yd�4�[�dY�ژ*�J��Mª>�̬�,I�������Nv�Z��\g�Q/�H�N�nN*��Kҷ���])�n���<������)����_^��˙���,|��c{��a��>���b�����v��̛�s��g��p��Hkv����ᶻL�����/g���=�Ϗ7뿇�l}=�ջ�'޸	�5ET)�y�N{&73s�^.�n�c�*:�������G�^C4�F��y�{��=�])�<-�5�+�{+�����sI2�h�A��D�����>����oY�՞́bAa�'~�����G�K���J__�I�����]�^2׫���]���´� ʃ�~�=~����o��>���{5�U�~{�~�m��|H'�
п/Z�)]Ofs�C8'lO1f�ށ�DV�@5�����/=��(���{��y�_��
e��@o��}o���V�_���Psk�,a�{���}A�����WK��M�Ѿ5�n�U��r91N Oo4��.�����wIR�:֭�2�5���7sr�'7mڎi�G.���kaRn�ؾհ��g����}B��^>=�DOo����40.��=��v5���g�]�ś0�0�R�N��}O܃������h1^L�#����tvg������oӬt�P��h�g��:0���),Ee�S�{o�ʯ9�nQt=�L�>|�v���6W�|oV7ϰnt��Rw�}ݤ$W�@�|�z����g�K��m��C�c�����쀄����:����O{�z����9��wK� 3ޓ�Y�'����4G��V;�c���oz�ci����U筊�SE�4OzfV��7�6�u�F��QLs�W�w：�w�i�b�>6���K�$�L=�E{������=����YT�I�����f��P�o�J�5\�W��Ϣ��>��T+����u���G�eM�~��~��񚽍r����4�x�����k�4�L�8u�v�y�꽈�v����z�xwk��73,=�v�$LǼ�>�o����z~�[!�ͷ�尾[�U���}��}�p����'yN�]J>¡:pOQ�<B/���\��`�~�y�[�#ն���Es�mL����9c�y�k�"��g�gTy�ܝ�5dsfdS����q���*�`kgf�2��jyk� E]S����^�;ǁy��f�4Ԛ�������߮;�rDP�"/ѠPƩ�64�M�cu�.���M������@����B�M���b��߶g#���9��^q���ޮq�(��Di��֗���H��z�l��o�*����Nv���q�pm.��2=���%��ʕ��9�w�N�&�x>k�����u�1m.��2�5Ww��-\��~Ƿ~jq��~�R�^���K�M�M���,x������g{{z�H����O�lI�fW�uS�sg���W'�����E~��et��/�p^8)/��w
�M!���HO/���]�鸲�w^C\�����5zz�\���@/���&y�홪V���.=�`��]���W�-PB�"��\�����)½����x:�߄��ޥ����ѷ�>��)'3��וܕϷ�気~`��
:}�{r6��]ם���HnN>��oM���S$�`��>g�VǬYSr�g�Qy3Ǌ�I�v���=�J�3�_�gX��O�c�3��L��o2��L�35�������6]Vf%�X���Η�ʤ:��Y��<��$3�
�������=��:|���S{�}���z�|#�o�ů����~2��O>����9Sϳ�S�i��S:�*����x�����,��C^��f�γ��N�g������hp����&�w��6gB�]ꎈG�t쫺�%�*��������SB}s�gw{�h/z��;M_�Ɔ|FPHg��6�s����_ �ԝ�z{�þ�{cʺ����]�p���*m��ۡ���eyt�3����NL�ykt��-|�b0à�`���YH��φ}~�U+��>y��k�;(]S#fUDxW��Ｔ�-�9�'W_|��;α}��̡�X����t������^[�����^�:�FF�JoK[�ow���=��Ҍ����g�� {�o;�-�3���	n�I2�W�4�K�٢T�u]�z��y���=��5���f����r���R��r$���!���7�͒�����w�sq=� ����n�:���v�Igھ��	p�R.�;��74�}}��-�E�ҭq�!b-@h��{�y�QL��$�g�_���Fz���Ĝk9�9�!�\ƲO�-^�ު\'����Z����1ù� �oރ۶��:���{}�M��e׳��{vO��P�}����ސM�>o���Kۚ+޲��������k���/|��s����Z��p���ܿ��ʲ�Q"[A���!o���0�]u��:=�<�����~��}���r�����[����(t��̠���.�ua�H���}������]�o�w	zi�~�%�y��|����f��,gK�r����K�'���^�Oy�g��b� *�5���s;۹{��cT;4�p��c��|�y����WY�>fPe}�w�x��R�YM���y{_���d���k��Ue�:vk���%�h�'{:�>^K�����s@)�<:H�(��k��zj�SV�r��n�V�큿eK�'Z7�c�ľ���#�1��!�2�b�p�#��7�_i�]Jq\R��4��5ȁ�[u��'e6�;�y]
��d�2���\�WtNq�������&�ޛ,�gU���ns�ˎTL��f���Ocys����Q�|�7���_2�y�$;�L���L�0׼������9��mP�h�U��
�����`��/Ij�}xk��MS�L�r�����s�=����`��=������8*���q8�o>���k{�_N���h�= p޶����7h��j;�?���L=�/=��n�z�X}Tk� ӒL������J��������=�g7:��i��;̢�F{Yk����������|�`<���]y��Տ�UF��^6�_t�ԫ\�Bv����i��;��4׷#=$�;=�3ϒ��2�i�->w[>?c���>ϙ�q]��_L�Jn�yR����}. �Z�ӗN��![J�9 �<��h�碠(<�V�^l��@�&�3��C�<���Rb��sl��3CYԃc���y��W޵���<E�X7��٦��,��5oc�}�;x^:a�cqq�Nc�ӡa=�Y�-=��b���w�v���;y��Y+l+� �4x��[*([~�I@��Ù;{��֊�i�E"�K\��K�q3K4��k�P�\>J!�@�7�������������x�uOhC��ty?*W��ˀ���6���ïD�M�ͼ�����p	��PSՕl~8o�$Gf���ٽ�d�gr�g��b_y��O� ����^p�Ԓ�!o��k}����!�Yp��*Z�yG�+��u� ��hw�vW�T�s��������{���ٷ��TY��������\�ۯOgw���x4�h�2��h�!Bǽ�@�zЂj��9�n�9������=�5ޯ=�]�����t5}�	��,C��?��>�	�{ZXq*<Ή��{���4�[����������=!���`�?��۰QS��]�t>��MP�
&�ڳש%n�����b���h&�v/�3��{�ӟ�k]|�zگ�w��_@oj͏�h��+∆�F^[�n���!����͒1T�U�w�{&�zx>�(
�C*S��+t!�}��t���z��W(�2W�c��!�뺹�wa�x&��������a�n�:Qź`=�6��_nn�^V��s�쳂g���x ��ʣc6s�+��ʿ-�+'���&+.o��*�2�]K��	�8-7��g{����w�9g�5�n�d 9�=��T~��
�z7�F>�+G_��<)���; �U7z��o^�Ϲȏk��wF��&��lj���n�^��U��t�s;�[��7AO[ڲ�oR�x�g �W����^�B߭������ڙ࠻�V�$���G�kg���=t��t\��s����7��A[������*s������[��H�6ŏZ�mБ������+<o�O��w�����U�Y<���q	���x?���Z�4�|ϚV�����������c���w.���?e�q�d�cx_��l{��"�K��9م�������[W�e���������0��w�����q@��E�����n�]�$�.�10��P%|��9�#���㝽�&����j�K�-}Rn�l+��.ZwB�b��ow)��KU^��L��]Wr���,9	|��39����,��]���f�ː^�7����xu*��ef���}b�5���Ӌ9���"ݫ$#]�u�qq�μy%�� �ibT�ư��F�+n��m�x1�s�蓶�����ԅeaפ���%����x0�`�V&F���`�1�[�9J��vB�u�n�ݛTJKX0�z���chR�.�_���/�3u��t�7+�����q�np������j*����	�7���� ���D�Sg~5r���+Y��1T�.��/)YI��n��.!o�gq���@�a��gn藹��>�1��%�)>ӄ%����Nvbrm�e)`�)���vd�{�ӏ;땝l;�71�V��/��w&6�&U��Awg.�V�x��az�Ղ\˝c�R`�0--\�s�-�,�{s0���87$��P��[�R��}p��s������\]n���rs���.|�6o�@J	��ӉZ��ʵĲ�/T���q�8/l�˻��^"h4�=w!^r� �,��������B��|�ٴ��:NڱƊY�!Av��*/r�Z��w���@�m�C���/.-�y�J���w7�Ӿ��^�����m���U�t0ss�|���4���6���+��1k��N���bt4���܈�Aΰ��xʘ���Sv-�&�q�/jt�軹@,��I�wu�kW���ɡY�E�±��9A��\�V�F��X��v�!�n)���n�N�C;�x��ZT�p�BnGx�An���x�K�]Pa�(�;4(���]����E��%������_o���k��̜THA��]jw�^I��u3��w:2�i`�Grt� o���P�=՛�"��M�f�>V0I��:,A�fL�������
팚���N�g\9f�A��p,B�조m��Cy�l��0s%�K��_�$Dnq���a���=��W-"��!�8�+�勐E�(փ���Y8B�\���,��4�uލ���ѧ��Qi�u�xZ�|�I��գ;����̾7�vN��ˤ[X���u[D��v��hm�zEx��7�bɳ>j��p����]h�8�l��F3�Y��r�$[��CE�GE�ͥA�Ӑۜ����t���jT�v[q�*����q$�
�[�S�E>�sdE��Y�f�k%Y-�������������___G�}}}}�q��h�V�U��R��*Y�['Ki��āTQ^l�:��}��8㏏�����>�����p���UK̈́�X+�#�!dUX�U��E��hЂ��������q�������_R}��s����h"ק=Rp��jDj
V�I�Am��;�y�w��ޜq������}}og��y�GW���I��:^U�^QE��91E�8Wە4=���?\q�~>������zs�#޸�]G#y�+ѐ�0�=^TAT$9ǄE-�>>���q�q����;�=��p���:�l��*����$#�i:�N^A��֫b��)����Q�����HA{0�ΰ���DQB�Ϊ"��g[=�[Uհ{�Tِ�TEW�A�g@{����D��"���"+Ȥ��PPc9���<��	�NQ�ty�
���ZE��&�'���T]�r�0RI:G+�aH�Gw�yu��1__U��Wb
Χ:R̙�X����K9�Ƞ���x���3�3�59ߞ�}���Ov|�����t����4���4�sf��vt@}�ny��]�,��1ŀ&ϥEs��'��s���ƛ<�(;z�>��o��y_g�gϝ�_=���ǉ���t�~z~�h��K'w@���c�Qly����0�@Q$v�Z�g���I�כS��{N���s�q�������Xw�(�]�囼�d��Ǭ�U� �>��L�V�(�]�������>;k y�\X�u�^� ��O�2��h(x� �����7�'�P�s�cC
����>xk�|ƹ��������l|*��D��_x��6�l���k�����P8@�ǂ�C� �����m=�.Pp�f,½k䀳��}s�y-�°�l�*�u~�eof�
^�|y��_à[8b���m)��o{���:|�]�@%��X��ic��??��i�Po��� m�|֛Y!�5��y��CykxY�@s$B��7��g�@�d@G�TxN���=}��z�vk���9�q:�3�P��=h�|V��� ��p0��	��$�%@�ko.�)�9$צဈJ<0�롱z⡀�l�g.C�3�Ǉ!
������^σ�>!�A
,@F7O��3ժ<=���}�gWN*��Ý��3e���lYR��m��1�<�Ozi�#[gşo���]���o98Q#@��?}�:�6�٠�=�a�NZ{�/8�j�=�����P;=ٱ=�M	E���;������[�λ�o¾��0�=��C~��?:���~��w�u� @�}���r@6�� @��������5�)�k{<m0�{ޠ��9���l��c�]���{ ost<r�3�)0������ϼ�5�����/p���3�!�G8w�g��0��� ~.xV���{o��>�>t���n�~����Ǐٱ�.�ރ�sN ;�<.��mYĐ�t��>����
��*̝���(�8q ��Ob ��k�J�'��B�{���j.22�s�C�A �@�s �[� ;x����>Io�|0�������Ѻ�a}��G:���ϳ8�oo6.t�����9����kb}�1C���Ģ���ɢ�q� `�{ d���5�����c;<�7$����^�{ @�y.��:b@L��P	�l���a c��~@X��@�U�Y�𶨁��,x�׍�����T�x%od@�`4��>u���g�����J�����U8��ȅFsi��~���j��z�_	�@B�P@E�_�۳��~���%��#�>�]��>�	^�t��V��sӭɫ٭�3���8Cl�%8D�'=���#�p�L��1�Q�Ch��vh޳N� ��>�y1���"ܬm[��UHze0��X�.���	�+!���`��|��G��}�'U��Y�.)6n��p���e��yr}�O��Ꮴo�WG�e�kD��y/8]6t��y?��^k�<x<8�y����8�y|�Ǘ�>��J��U!i�ܓ�u<Ө��_}b~�����@R�+sΑM�R�U����-�Sy��I�.�����^D��	'�3��ԃd ��s��}���l���5{K�W[r6G(����vߥA��F]��^='��"������/F�a<��j�] e�،U�T�����)U�"�&|�Np��%�KWM@L���탘� G'�H����p�МpK����b�5�d��ܭ�ƫ�
n.oZ�v=�
ꑒ#���	�R���26X�=��|vGvۘ�KΪ]fn�s�į��#!���EH��N�J0�>>�1�-!�����`���d0���^�-q[S�!&i�&��W�+�y����G������4Zz8dsc3�ad�g3��w��FL��ָ�]��/[=0fe��'��j"Zߚ�����m�ƭ�sJO���(�#�F�M�����O��e�-�H��(��f�8����\�Q�֒�Y����)dxS���.g�R�G37E5��`�,��_�Ε�����d�p�q���Ӂ��(�>lzL ����!�� �1M��-��Y����Θg=x���8%�|�q������P�0D
Eg*0�
�1e��l~����G�g�^�$��>�s�3�<�=��j)���A{hf��11-1^��۞1x	��ٱ���?cS�X�,X8&v�n����3d��v]��%��%��r}�Z�C]��;�-�q�����<'�D���V���|���<�cN0�_�<`�C!u��`K�D�v[���r��v����-=���_=��f`ȶI��7 9�� �O$O�/g�W�5������گ�k� �/�}�uƼP�u�|dD�u�[T������c��L��H$^ž/=״�ʅ�R�D���6-�հ�g�<��יٖ��3�w���0mj�㝛r'���-��R�wi���{�M~�9㤡�hǘ�F]���z��i;�����+�u������i�.��=��r&i]6��!�ߕ�J���^�~Y^�ߎV���I� ۅk4��&��w���"��@:��Y��sp�y*R��%'�wl�	|�0ogLxT��l��Ì(4^u+��:����1�[�����V��O�o���L[����h=�M�Co����.V��н����i_��/h�wB���Xy�sB`0��N��
�MB|�r�]�f1�v�����!�O�w:S�h�L����=b�t��Q�>&~�>ʌ�6<����5�ǎ�݉�)�
��]�%��&^p�s��2bM���;j���if7wh4a�T��7˿�[^D^�{�9�i}�}:��]��ȇz�t���ɻi�^�ðҫ�;���y�Q!w-]�ԫ�Q�Yg{\���!���hM�}�������<맡�ǃ���ğ~|7��}���~�����!�!�~q��I���یl��4�����p��2���dw'�ݜe�N�߷�B�C�����a�g ���k	�'�ϾL�_�E����9��J4��Y�h�*{����q�RF��
�y�ԥ Q�Z�5�x�1K�/�ٰ�_���s���:w�mA3h=�ǌ�����0�[ʳX�,M�9����d��M�H�`��ߏOˇ�u_o^�����! B#(5F���짇�{:g�>�(�+�ɵc�IL�Fb'�r!��4?S�	�:�e�l7��F�1c�L�C��I���_��AðP�yK����p��4�=�e�9���bex��n�e�<�ie��h�3��?�j�~���X�������:8*����.�S�=��ku�lDϨ��ဃ��W��_�K�S"ʦ����/'��?��߰;i[��z��t'�[���v'�V��o�L���ð<�L��L��{V���Nommrw����hld��h�(ߵ��ӽ�_�d�H3��H����6i���P<|�E��
+�w>5�&�W�}��C�Z���]Ӯժb��f�x	;��R�L�����vev��M�E0�/" P>,�yt��%�Fiݒ"K����%&�w{��}N���{q�s�ܝ{޹ּ�+���)���c��������C� ��G��/=����`�s�������g��[O4kt��y'�c�J(��V��Xo��׾�SZ۪O�z|6X����j!랽��:;;��"���V`|L�?�ٲ�x����q���QӖ*`�w%�l*�X$���R�~˟�#��ä��X�q/����Ac	(�>����4���|�[4X&Q۩�|i�d�A���e's��?W
�/���$hN�PƵ8j%R��b��V޳�Ԁ^��|����ئ����f �ߎJ`�`��>��F�2*�������fBL3��t8�>�ăQ�v��H7G�����1��bd����Է���J�l������sP��X�E{i>���&�ב����ڙ�De�f`Y��OP��j��YM8�:2��^x�Ki�`�<�O4΁�ܘVo{d�ّ]>��Θ���x�˕3S�ؖ-���f��|\�N���`@z�Ih�l�[��-H���FL֨l�����l�[
Ӛ>����<��H���Rbm@��8mp��ޱ�2d���إ��Fs��}�Rr�ӛ����]���0qÇ3y�u�=�-�f��7��7ٵc�\��S.1V�M*r����׽@4�9L��Ʒ�Jn�Wo_O��i-|���'���'U�qM�s�哯�{�Q���`�A�a��e�2C�x=}?9�%��$�M��4��v
_���nj�h�#)�-�I#zkf�Ĕ{\��Ƭ���I'M��)D@g���*�	��� �o���m7N�]4�hf�,���W�Bx"*$������ �F�[�>36�3d�W���N(�&� �Lxj��S7N���zu��'a�=���r���;Ս�7-F�j%�����;���.P݀a��U�,��)�k�[u��]�Y^t���n�E@�j�q�,~��)Qw΍���˫��B��#� �Ywg]+7Նf�L��Ň��d�5�V�M�e=�^�~�q�=m-���)Y!)n��ؖ�]����3���{�K��Ȉ�/=����f:/Sx�놣f�7���6�E+�d�����u|����vj���x��,��N�E�(����<Z���7C����r�nV҄.[e��q�����Q����۟K�mK���_�x�:4�z�l;,�vQ����g�pe�jj'��� �3�a~�~"lk���}.�\�};)B��.a�>�x�yxƖo˹���8˥����������N4s@z]"y��Fʋ"FN�_��<܋9�=���yS�B~��rk_TN��ܾ�����Zj[�l�[؈�T/�L�o:;�g����+d�k�7��7��q�kH������z{���[�/�}��2�.Pr�x;3UѸ�(p��	����ݏ�re쫷��>}��տz�|�����BHa���x��Ϸ�������~��뽳<��f�m������5��a3Oɵ6�
ДqY잌S/��m��([�Z&< Io"�#9�L ��˔��L�a�����[��4�d�{��S ��4�jV��=�%�arl�,gyؗS8ssȒ\(��H0��|��S.k^6�����}`�����ɟ��yÍ�o�9���n/���Z}q>n�V�-�vc��ʄ���X0g�C�[0d(�(}�t�h �į���}.�U��mv�(k��A�8����{[+�Xu����U��>,������u~9�8>L'՚�_�.��.����[[f���/k��,�$������s��Mg������yV���U��/��X�,/�{T�R��|��*�v6�zr݈�f9�5Ā[��V��a�D��b�ɘ<	��l����sH�vտ����v�����ݳ׷)W��%
��~�7���1?o���i(�����v�8��>ݽ��d#��(�SG.�uz�[ɵ^/`�6�PZ ���S��6F������V�?E�'���I4����S�y�j�=Xx�����3���wO�\j��}w]� z0�}��B�R^Լ�>�Fz�4{��X$�x���}*^ʰ��;rí
;�;*N:�"`h�i�^Y����s�"��A%�°�u' !��V�9�@�r��Z��}N;�{�z�r�(����;r,��)�"OZ�&��Sϙ��0�ld��x�x�X���"L�:4��p4�7��l"/	�/���ʢ����Y��#�E7mO=�}�j�g6�t�(���&݇�a�<�I�m���[M&�ǹG[a�ˬᵵT�<r�l��5�1S�'���C����m�<I��z��Cj����l)f3�^�u�	񗿷���uEIA���ÿs_��_���<�k>j�XGO��\�� �%�n�#L�×�:�]��A�������Z�qc�h8��	�pN>8�\6{ �	?S9}dm<L��l͞��'��k�lH!YO���K��yWG��~�h��Ơi ��V8�s\4�u��^CQ͘r��]�t�4��e�&��-�C�9���}����~���!<hh~kE#[����pu�U���Ե����p{ֱMeE� �6dC�ސ<#��6 t��O4�!T�;�uz�ej���rmͻ�.�᩠���-���w>{���,8�`�j��i�a�3~/����(e��Ժ~}m�h��Vu7�s{d��Μ˭кYwiN*�k�h�W��Y�mǦg@�]���dzw���']�]�*�x��T{uܹ	���H�����t��0'.���0�0�u+�����ߞ���z���{͌�}u�?O��X ��:P'�����U�?&�}���b�55i�Yis �NH�m�,�N�Pz���@�o�ʼ%?DK�;��EfD䖚��̼�pw�c
��!$aFL�y��߹���D��{���p�ߪ"+�v��RY��w��ɭ�ācF�=`�������垂:��[�A�OF�>��G��2[�?ߗ��+s��nkN���^+�}	Ɣ�g�{��/3aNv���d�
������=(i�w�ze�<~�>�����jg�+&�^�қ,n:/������Gx��j��l7��ۖH*��k������f0��>R��&�swPn����Hs�J���T(ݐ��m#��.V?�7�=t�q�Le����A3�)�ٛ�pDU:�n|e`��Y�S����C^��\�a��#(d�׃��p�^rD��E�v�B:Q�9���m��zi�%���S��c�@c�ؘ{�;cY�����f�l�C�,�}mQm1�n=���k���G�P�����w�׋�u�����Ӝ�QZ�c��z{Ϣ�������9�(���"� 0�W6�a�=Jx�aʬ˽���u^WV���K,��[U���[��㨧b�\��Ho6��{L����1Ҭ��<r��^*�.���3�G���5.Y9z15n�Uv�f>Nΰ�Ǘ9G�VP�q��%o�;Daeh�G��>)MLc���E޴�vR���}?l��H9��c\����$%���5��ɭ;��Ͼ	�������G�1�=y0�Sxe�Z�ѧ��OI�mAg��k/!s�7J��N���
�\T�P��vu��
Y���=����h���P����:�Ď��5N�@N(�[�֫sq�;��lJ^D�2\�mO��������9��M��P]�w�	"���onfE��fͤ��U��ޞ]aZ�S"{o^jc>]Q���L�#6Ѝ$��I�#2
�]}�ǃ�����w�����,��cc0�����cea���.�g�"흉�vD�F7o0�s����sf�/&�u#;;�,��wڅWrW�l�0�*�C5<�:���)�H�E�C�D�
��Yܻ9*	�����D�YE��c;��\�M!:�JQ�D��]�G ����8KϢp��.�X��[��ڽԩXD�f<�"M)����i�eMM��R8��kW;>fe�Y�l���z������1k�=�Ŗ�{);����*�b�f]���
v�.5q��ŬG�e+7e��:�\S����ϖj�6�C����w�u��u��|��`�{+�
�s {]���#�5�4"�N�Z�t�w�/Wk� |Z���3^���d�75�tS�SG!��`Y�\�yPy6�)K|{�l�ӧ�p��t:U*���Q^���d�m�dۑyZ�7z��4��X���2V߈c�/��6�F΄F��D쵿RGj���\�RἎ�Ǐ��Vi��� �B��wt�BZ��t�h�I�_)�+o��d�;��'�"%λ(�u�
z�â�r���2٣��Z�L��u�;-�8�r{4((ԍ]c���ɳ��yO�riw��k�w}a'5�P���b�7_m�]ɳ�j}�b�t�+�K^�ԑ��֬=�7����{9��C.p�8�V_Z�C�6K���eL�mLM�j�RD��18wp��ۨ�m�*6Am�.�lD���H�ͷcz�Y��Mθ�Ǉ�zb�Z�f�
��,sv3��[�>KX��j�&E+溭�.syn5���l�5����僳��	���%���ȱ��y��o#މ����pв��af�8�F��peM�M@�������-Q�N\Wk"^�{ב��S����l�����糷Q@�ǅ�f�U���v�J��9��j���A*�T��a�`_��j��@^Zt�ʃ�H��a��� �F~g(�H}�_�=�1�����q�_]}g����J� ��D^�#�	� �����ގPVp8�_�����8�~������T�+�&���9DTD$$��Rs�!�Q�:<�]�{�y�E��)�����~8�>�__]a���=�Eu<��8Q��"�H���TU�<�s��}}q����8�����a���W� "��Ң�XNE$�6�F�%^[:���۹�y`EΞ�_��?\q������__��}N�����_ A�3��U�6@QF����������+%�9Ƿ����8㎺���a��<��W�E^��1l�"*����׎�=�T��'�����ȣ�z������$���Ⱦ1EZ�DyL��y��~�+�,��^^^UU��TQ^���M�H���I`�G�Y"+ʢ"��(���Y#�SN"��@M"	����ړXa��5[�.�Ҳ�uk�8J�6��k4o;J6��ϾL�x�YI��5��6��9t*0cn�.�[��Pg�)\NL2AXi����g%�L��W���֝_L���r��Ylm�e����m4�a��an�VȕWbc1��Y.�,��]7Lyv���+z[�kuG:�f��J�0t��%������mВm�T����Z�V�Z�I��˫�3�t� �撂��Y�<���<��Jj��$[� ��rr��:�x2!��NC�F�ł0�"����'V��{�I�zԹe�����.��(�-��5|%�a!%���h�M����������Ogk�� ��)��Lu�L ���8�r��h�ė���l�x�&��gs崦�΁���_���]ő]�/=1�>���Yn��i+)��sSF�\�_�.��9�<�\X�s�έ�=N��{�@���������t����x����q��w��{�:�N�1~�����_�,�ȹz��D��{6z)G���>�h۫쩝[ҽ�2�{K52�q��'���i�<��D�y�|kc���T1��r��I��o�n�Gw��H����K,,#Ks3?�����L`}��09����A��̂���8}hU9��R���J�f|��m�@�H���,]S����c��gE34w7��"����g�께�ngD��f&�P�q�j�p������ ;�u�E	��Aц��4h�z�~��Z:^�Fn��z1��%m�ߞ/ޣM��d���_9�$������`愷����s���v�6�4x��9k�^��F�T]z�]�&{J"�[_pV}^�vg��>�
��O,�����?=��NuX�*dt���S��z������������5J�+ǹl���= ���R>���)�Ə����m#ܙ�3a'����"oHZ��]��(J?9���$.�q.�K���Xj����Ǭ�A�{�� ��Pa�XdR�@a�  �z� '����ʩ�����ool�P��+j�H�q���|����kp�5�Yp���_�q�i	�U����)�2���(r{Ɯ�$�M|���(�*ꡏ�5��0�M�w��tt�s�Ջjs��.^�@�QtX��Av��>�g�Ѳ���S�~��L :}/|�ݧ_�_�׆���Z�w7�x+|����١�2�K�J�\��6|#7�cK�=[�m=0�7\�kTb܈]��rhw�]��w�N;���Ga�x�� b�7��@^:�����i�P�7��f�Z�u�BM��Q��!fQ���2�=�Y<�>����R�>���E��e�\<n��R���C��~	ߐɢL	i#�����i��\��j<x�A�\Yp��:"6٨���꺦���vf(]��z�/��x�6��;��-��|�Z�[�c��}�K�4�����5��[��>�P��K�)���Rɠ�M�/ ̛�'�nx��-�d�(w��H|��-��7K����w�o$ꋗ���pG{��J/�_��F�$�/튔�Z$*��-w�,|u���~����V���M>��mv�l�1X_JH1�x���Ai�엻Y}�y�&��U��k�O��5-Q1V�|�����J/|}$�A?U{} ��Z^��Շ�Ӕ���X�!��;��r��뭽[:�2�h�ܹ��o/�[�����l ��r � ?��dA�Pa�g�u"=��^~|����o��~�ı����o)s�/]oQl�i���X�� ��f�s��r����K�OjnA�2YO.C{�؁{,G���Am2Z�SX��f=**�?����%P�ͪڶ���&8uԉƯ`aOْSH�'Aa�a��(ߝ�g�m	a�zȎ�J#�Iͬ�{�n��e�c��,y@Ν$��Ʉz��ڸwlX�e�K�;��Ha�;��g�l��U�� ��y�{�o��-k��)!�ߌ?K	��r+ͯ���A��d+y=:��"�\��v���h��(FP�;A];q��.C�F��B�?���[�$D� �1�2��TX���M��j%�c��rB}�Ui���^ Io�
�,��6B\2f�Ȃ�-a;ϼ�&�)�i5�Oǲ���X���ڪ+�F'�F���j��d��E,+ڎ&?$�οN>���S������iK͝�Y�i���q� _��5��xx�˒y�a~��O�}tsb� ��Z�kMN��ݻh�I8�Z.�R������&c����쬇Ӄ�VfEθ'���O�|a�n��s#�	B6��%��6���Kh��4����cN�f��WR�zf��_�CJʗ'P�×�}�����UG��^z�_L�GB(~
�݋2>��ʞ,��9���l�Cp>;v믶n��2�[
���G>u�,��>����(�a@�P`�tY�
$0���홡]:HALG��O�{m��;���Ϸ�����{��]r�Ϛ<�e�X�-ݰ�%����KK��@���OX�>���?Q��@'*�ސ� H��E�PD,/�9�D%Ѩx	[8.@,/�)�6:v��zr���״�l�� 6q&ɶ{�;��~2 ?]��C�8̼y�Ũ�`>S��7@p���Ti�'����̗!���P�7%�)cbn�x��=��8^��O���]���,r?�r�i� �U�`?>.��{#=���v&1Y�ԙ��i��4ӄ��~�=G�ǃwL2h��6�3�����N8����O�D����i�QS�;��<0�Vtz�����S�p��*"3��I_ʟy�}�oU�-z��S6�T?�sMK�9��4W�ç�o+�L�#q�3i��̐u=S��17Pw�z��.�� Yt
��瞍 �_%u��^��9<0-!�{���}"�z�)�i>��~m-�3}�x���^;�6kɣ.�@�>��k�"D!~[� ���ޢ@�_��\��۳Zg��[�ro��!Pʃgyw�[{zX�Y�m.�z����D�l2)d�� �*]�]=��Ec��8+5�|��>R,�x����V��x3�Z�ԏga}���Uk[�����G�[]�������7:��.����x��� �A�x2�C��(���8?z�?I��J�df��~���8�ix�B!mB�V˴:������?���_ZR���k�"��զ��cx�����hg~~��m,���l$?~~�v�oC�n��+Y�޲�Re�l��e��#M*�m��G���<?A����
�t�t��vk���=9�6T!v�R��~��_���Tk���"ðlwcd��Xӯb�^5LY����_!��*Ydx(�Y�\A�H��T�{�cK#�>+/&�����X2���;��Z��0BN���К7�̸��Y�&F&�f�6E=�Q�:�ow/J�#�����T�r&�Z�w��E���H�<SG����#��=��0�܇2Zw s�UZ"Th���Vs?
��C�*:j ��%tH~{��@*�M�D{���V�8�u�m
i�FOq�mu��g���Z����L��H|��ч%���|b�1kj�pQ[NM&�{n�U�n%�fU�1�����$�g��-�`�0,ރ�^N�fi����󼘄�]��3�.װ!E���n���oy�R�FP�chM�11�7�ͼ� x?�ɼ����fR7#���'��
絴=s�lI7Wb�U�[p�Z�=�&csc�f����1��̳G�*����No�$�ȁ>�Q/�}������_l�T�9�����g��:=�ͺֶ�h�*� mf�8���k+AW��� C"�0
C'��E���"u*!J u �+��6�ɾ%����SxI�j��?�"��>5F���5��{'=�D�k���a�ZO��in^w���6n�H�V��^��j0D�y1M��q��ۛP#P���	=��x�̈́��k"���H��Qe�'�oqs3oɠS̠\� ��"�f�;Ֆ�^��uuhB�Iu��)fKV�qc=?���jlӷKxW�q2�o��fU��l�S���je����;�5�:�]�R%6R>��$j��j6� ط��Mq���~�:X���k-�lR��X&�[�4�>��f�X�;��
��eGE=���ơ�3G��7����LF�I�t����34a҃�t��c��O�5Dt�&!���"�ؠ;)B����7X~��fȻRL�/W�����d�80\ioM+\ps�d3��z�a��y����<�7F��.ۨآauga��[��Wצ?0e��52(!<L5?rIo☗ǥ�&}�7��L}n��*(np���ي-xD3�	�}!,5g��5��09oip>sH����$6(ȃ���a�ϧ ��p��^����}M����5�u�lێ��B�O&X��뭗�u�K(��4B��gNt*�U%!�e�m5Xk����Y/T��}ٜy���S6�9ښ���d��L �%�ZMQ�T����7���D�ոJ�U�c���`A�`Q��a`��`�@�{�}��I+�T�~O�}���;�a��$Ӯ,�o@oN苀���l��{�6���<����t�a�F�Ck����ם/P������'",W@�6��b^N*��6����{��j�B#���=b������g�y络q=O�Ǟ`�E�����J|�:i�*�U��2��<F���w��`��.k&�Z&�|�ߒ����;���	Z�z����{O�`���)i KD�P(�;m��k�4�S�[F�.W'*+�+�*]>/����T~!p>�]O��L�*�=Dx����8R%��)����D0;cG\��?��uY�,���X�fZA(�d^|��s��x�r���h`�8����)���m����+0%f��΍��~C�J�`�-m��-fdN�/>�;��`F9M��UO��ϺyUЫW�$V6�U43I��٩���mش�"��Ê�q�1��+���:�@�y(�F���H_�i!,��O[��9���~�us��W/i	�@��4P1,+y�%�������/�.����QW���M<%;���gfaΙ�ZdJq	9lJ��<)�Vo_V,#)��R����E^4������ַ:Z#����R�ٻOU����ͷ�N�����m�}݊�.����w�B0[޾UuӮ�_&V�|����>������?��A!�!�PS������y����9ᐯ�B̅Ys?OE�?xP�������-��AE�r~L�kaو�c���U0���n��� \5V�[q�G8b��'$���,�̹�6�9�yS�H:���?r�l��d'���X�:oY`g����=�	��;:hw�$�ed����g���X����jwj��8`�<�9�{��d���(	a��^��mc��1����l&�38kGAJ߃����(���z�,ݱ�]�i���X�d"obh�djS���1��ֳ�ƠEk�C�����..��g�\�����[l7��r�_�����3q� ��=C6 �֛����<�|Gs{g���bL2i~"��q0�����k=�l��+��=���Խ�����=m8y!a�r�^A�	S@un�`p���L`�<�ٚ<��s>^��/�sB�_F]n���D��p(a�����Qx�e�W�����+y2�s���cv�:ڽ}�'6�%{go�a%mT��֘���m 6���/����I�:���	/�mMQ�=ī�Ȍ�j��D��i���&�OW�c��E2���k]f׽~ϡ�9��7�m�p��%e�s�
����ʍ��ND^�D�>�L�wV�	������_���Ŧ�\7i��3:����@ƾOFt��������}��3{�:?J��U!�B�S�"�0�C�(r���='�y�u���XZ$�?_߿��^҃��D�10��r(fJR��f�CS���d1(a �D���kV�	���3�Jc��ցx�zFuK/0���;��5�Q`�ۥ�<ȭ���P�T�z�&�b�L0�e�n�@��p#���%Q�VDS��Vn�����TI�8��� �O��F����ha0���1����z0-������V�QU�]���
Q6�L�On�6���ݷb�]��W��0�n�2a��G�`B��1R�{=	��'&o<Vf^'b��8S9�[v�XM�!\\0{Wњ�{����˕	�3��	ֵweL�O۪���ד�fk�0͘��:X=R,TmHs�qZ ����}0�@�gŇ0�s�U�5��!��Y���.1�j�%�j���Z�%�xP!�u?"��e ���W�|�������+�+��R��H�i��f�5�xwli��noe �nq�.���{�c���{�rds)���I��	����%�m�S5���{M"#����6���8�H������ǧ;�O:�gQ��Ψ��=������^�ħ�K��:��C\�l�l������n@�;���h��A����&s�/ fL��+�a���/}꾵�jo:&�ZS�)2���F�[�����Ѽ���h���Td��JhK�������X$$�0�D��AAQ~�����>z���,ʽ���>��Sw-q��B��[�bRgD��/c�q�|%l��D�߹��|�g[��?`���^�:U�@HaP�Q�x2#�ox{�r=�����W^ z#�4�s:cuＨ�@D�q�_ �?HK~��ow]���b�D��H��[�L����ze��Y��-XB�� ��v����bq@g�0���0n6�5����|�����W���u�� �۬8H��7;It�^]�kEzEk�)uV#|k�bjb���zOMÃ�Ǔ^��oL�:��$���u囷�H6s���e�&�F��-Ë�q��˄��4�i��N;mɯ[qb�5���s�0u��W���VR�Y�������H~��,����AT���*.�F_�ɁM����I��ZX���CwKp	n���`�(0��G`��~���Y�Pu4vf�~^������e[������±�,��'�$x��9	����xղ�2��
9Es
�Y��v�~>�®K����sMĨ���~���eN�~�q��c|Q���3bl��սs�)�MA��Wr��kf�0�[��0���{9�Tΰ��jh�s��N8�z��ivS@�^�km���U�#3ѝ7�����z<=�x \e�v�<�&�Nj���zgF��+����*��QÙP���+��+����#��Hc�#[�B��W�]�u[\�W���r��Y�.�+n\T�u� ��R�aګ�0�p���uh�A+LV��Ǚ%����r֐TY]rXp��qũɨ�ڒ^v0 "�A,Rڸ%u6�aY5bt����F�ƛ�Y*�u�
�����]Q�ݜI3o�a53��Z��f�a��
d͍�N����p�"[�#��s�Q�Ɨr���ē8���wG]���ʚY���n�ؔ���{�İ7���٘�M|1JtvY[�7a]o�\�8���u�o�8�&n۾�^� ߶��኎v��x���Q�=�w]%K�0Dܢz�/o����X��N�N�v6�3�Y%��
ۈ�!ZV�M�W�/tЋJ�:��͖s�9V��J��^���CC�.#Ҧ�|j�J�܇;�n�a�n�A�iz$�m�P�(-�|w�23Xb��ҥ��p�q_aqʋxXG�_ͥ[D��Ƴ)4Vn�4���3obu��t�1%ː��M	6�|����8��U�����;o5��]`�$J��|�CL��d��w��l�R��*��;�a2q���'�Ug�;����u($uˉ�u����Rڡ9>n� �,;����KAi֛���#��VL̒m�F�52�i�j�%�'~K�&4��(Ŏ� ���U0��*:BE"�HH"���#��J�KF�F�����\��[���`���v�R�n��q{�c׮k�
�ݝ�����m�pr���7T�Z�2p�v��d����=W�%�����2.�؍�ݜ!#mu��]w�B;z�\�<x��bرT�2��r��5ܨ�I����i��f�q�zD�YZ�����ʽ���k��V0�q�`��f�i�יԀ�����(K�1vE�t&�Nt^c�Z��ՌD��W��I�v�(�Ԧb��YN �����ݽ}ɭ;������
�s+��
�"4��p�z7�64v���n<%Jޠ���Y�E�����j�V���@���k)���r��o_mm���Z{3�3�|��zo�a��f:[b��q�)�
y��J�d���5vԦuí2��aG+�oe���[�p����U�-�#��2�����8�C��u7IFۻ��������:hj�H�	f�H�!��.4�ݕ������|sfm+�k3k���B�S���,�'e�M;զ$�]@u�e�Gsh]���>U�rȗ�"�Z7p�'�&�4���29f-��p�+oX;l�$��[�>"?}B��aA�""�+����z**"�+�yPL]G"�	:z~?^�q�}u��������JH�\.��us��Ԁ�¯��ш���r$M���MG(�
r}q�����8��}}~�����W9ˇ	��XȨ�(�!��QVN�D�W%�.�LDt������q�}}}}~����MTM1E*������T�X���2N��*�Ղ>�Qyߜq�����>����}}	b(�D_�E_ӧ"��^�tAM �b�"���8���p-�W�ȣ�>�=�>?\q��������Np�1%7�8���@�,z�f1 ��:DX�����<
"|�����o���q��������G˕E����V�S�6yE��UE�AG����Vɘ�ŷ������*(�ϒ'���Bʢ'��}�Y<���r"(�O!UG��
��
��r�*���y^UyQEz�$���2E':�{x�u�DyQ�_l��#�^�>B<�����<���t*�����Fk{8ʊ��0����<�����8n��li�1�/��7ՏZpi�	���x��x��J�ʽ(�*0#�PNՕG�=��{� |�c�̿T�}� q�n.&�GWJ"]�\�_Y�Y��V@,����/e�ǰ��=(b�Z�桬�\��p&ؐ�ų7�zЙ�
]"&�7�P��F��#
QTե�d5���y-êX	"{<�(NY��Ls��WT6�wwT�^��e�Gx�'թ�0`�)hZ��VZ\h�Sv6�
Atq��9���<}��9�D>&��b��Z\[���*i�Є��f�wf,�-m���%IH�Ym![��7��$;=}������}�7�a��W7V�:�1c���:a���[�0�cq�����;=��:y�9��ۥ�+r�&@��\�1{�	��%մ��EEJz `fj֌�N������]��S[�m�gL7U��*8Z���T{Ͱ �I~5�b�~:�f�+�%qcI�*뫔Vdk��d3��Y�}����]P����g <<���~a�[n�޺*�ܖ�K�X�y�hI]�N2�-p���P(\8Տ,���,D{!���<D�&�(�>�b=/$����F�������_Z�[d����/^��R���a-����LM���-�H����0�<A ���v���\��=�0'e��+��%ɀ�o_a�N�t�^c����(�YZJ�*Z����dFT�U!�XdF? ;��<����~o��?��G:�?�=YP#�m-$z�~�A�Ml�c��f̵�F]���#ёK9딑O��iX�7�ǘ�z�oM�w)��W킘���M�6_)λTRь� �H�(>�����ݾy~�.�g�_3���:�G[�R��j�v���j������J�؞���ʠ]��Î��\M8u�v���Do�f8�_�����u6L���ʎ]��ʔY�i��1��_к=��ĸ����B���͍�B/��Y[�{��T�,�ۿ��>��%�@mW�B�h�+�K���q���=g������8�����B2_f�%��=n�uel�i�U����~xx�˂L=cA�:�fZH%V'���W|�>9����}T�{5�jb��p�	��cDw'�������.Y�'\�1؁����TV��-�}��axx>4�t4&��Κ{lq�e=�S�>c�����a�F~B�����_��Ȃf�0M���M��[Jlvo S[�`*���z�ĸm�>9��0:9�Y[����-��.r����%u�'<4K&8齖�S�%2U^kv?7ᜇ��I�{�oq�c�WOyE�)���>F��L��W	�,f����$p�[[�����E;9�z�>�����`RA�!�%
C
�  �$�ð��Q8�(�
�ulw_��릒��t��n.�rlf⶛���Y46Ӕr�G�t�'���D� ��"5{���5�`��n�Q�=�,����i�����b�-�:_�*��@ly�1��)g&�6/	+&�C�r��rw��m�h���}_Wi��u����^Kp�WC�p�����P��Z��3��լ�'�τ=E�/�y���C�y4�9���d�#�zz�
�G^�$�RhV�:�z�|2{�2s������)u4����!Mdy����~'/^9�Ηb/���^���gM��D��ԟM��Y\��>쩷3E��Шa��M���ç�gTA�J�K���r�����S�y�*��Z����`{�föﱶ�N�b��}�diW�֝�[Bh����,��;�5M-7���j^]�G]Q������sI�ܝ�
m夊��`�ik�����΄�$m; Z��p �e��-��o�u=�u�xZ��2pΫ���5�Z�� ^���v�A1t�L��:l��N�H��X�Y��E�%��L�xr�G4�̠��1�]r2�v� ݉5��2'�d2����-]��y`@���֒����jaK�tM���3�^����܃�}�UIYT�$���Gl�������>ȍ�`Tv��Y��4���q!/��eD�g_���s���8�k�q��HV�gP��Ͻ}:?@��`�@2T����/Pa��>�zw�^�����5�5��)(��hk�r}v�'�y�ګ5	�,R�O�v���x}������P#Z�4'_5�U��׃���Ph5"{�K���؎ũقv��_��B����5�aqW�~5X�H�ͽ����-��ٹ�{��,�Qi����ҜֳKv�9�|-d�`\�n.Fk]7 _׮.�y�Q��b N��W��z�s�7m���V���y�#	5 �s1�r�C��٧�$��Y�r��=�t���R�d���a>��ߛx�S��J$��pm�78b�Ս�:��m�i�Tqt�()(�����H�c;�������z7-�ϺぎO�;�t�2|��j�8�u���~YϹ�����<��gz��\���[���E��'�^'�=O���H}'TĂ���nql�6y�:��r�.��</ܝyRB�]���~���\�l��q�1m���w�K��ė��-!�Kg��}%S�Z)Qy4t8фr��b����1zVس�鳒���#4��V�ɓp�������2�zz�c@��F%�y�0E^{�����:"�/"�@���4~�*��J���	5�_{3Gb���Iٳuhۮ����z;����z�̧�9�W�{���T�9��Ha�W�Q�h�@�������~~�(�u���������\�+7���[\D�83ɪXv���uGHȹ��Q�y,�1�[�D9��B�r���w�۴��_�$}@�>ciف����ps4Fv�[o]�ܤ�<�t�o� �y�7�f���iUφ�w��kf�f��]�U�ۡ_9�x�|��ei�dv)�$i����!�4�h*}���P�UxeB��{�T���f��ɞ���d[77=Cb' ,ѳ�5�ៗƻ�V�y����5�s��(�Oǟr븽	���Z��˘~y�$k���eXH/<ֹ��
��	���3dZ����ps:�WZ�թx�"���lfb,���'|o��m��7��P�2�a�ǈi�ij����bWk�\���at�!a��|ā��08-�%6sTC�mh�����m��Bԩ.��G���B��A�B&=�4��yY�� ��ĂƟ
Q���p�f�V�&�ݢ�m�{�d'@��8i���ն���c61��i�w�C� Mz�pb�V�I!3�h���-�9W��wn����N�e���6]��2�3�_T[��l~U5�>s�|w��ͳ9�����Zݬ�T8�E\���i��'H��Ovfu��ج�s�ee�SY���ò��F��{�x�,2r��/a�=�1���1�|F�������/���&턀�y�3Z�i1����9��|�e�^[\=��[��Y�[c7����� �~S؎#�um�=��g����V�?y����73�d��H�88~R��-�7�0�-����i���b^�ޅ�ת�.j�lн��N��*�?��@����g�����CbD�|���xse��6zq�:���8a�f���oO1�����qڼ��Y�c�?*i���!�hZ��~S�k�ڞ쌈H1u�7��;5�h��f�x��G�4�:`m����5"n�K�G�����hF�d�Tv4.\iۙ��c��I�.*�lc?�V��� ��n��b�bL2��l��[��(��5w���]¼�C�zlp�4��8�zm�6��q�5��
�d�i�!����]�=��(Z�5�ӎ��Aj F'��®\qỳ�=-p��N�%��t�]%���^��$ӌ������r�m����q9>/�免t�O��(��f���aPB�����&z�wP�&�f'�[�f31�Ⱥ�F��mJD��}6f�.�0T�α�/TH���	M�����4�k�a/N��+a�V�� 7��3�mG��]yߗY���|��.� ~��x0�B��0�2�0&������I������u�I��y�~�~>�g�.nɐ�&��"�6�G�e�sm��
I	�rm"f/�B�������ǚxu�&P7Y����Y���/�6g�[��
-WD�wٻ�վ�Toa�⬏0%di������0�׷���r5�8��1���'���G
��`�6=�I�N�͔-�ʑ�>c0{�0�p�����74����,,�a��%K�Y2��{!��I������G�Y^��I����n8;L��$i<����d!�}Ny5$As� 3�:"�9Ĉ�ds�s�ሁzqŐ$�zk�}�ќ�U�i�{2GK��A�d;��96�8b�4���O����u,�b��[=1D/.ˁ�Ux�w�C��N�uʽ�%�%�����8lO:'������o�������L�Y��s���yܠ*�2���b8�ޣ�v���k Nt �#2���������[�R�GM�$A'���i�><�xoD5�Xe�g1-��>$�U��ѝR�@�zgt�blK��uM�*��F��]�@��f�8��*_��{�F�^�T�Og3Jǌ��+�F�_2[[�Z�����{�������=�	n�P��}y��#V���:���c�m��\��#���_|;�U[����	X������n��1_N�ĕ��)�_L��N���v�ti����]��C(�C(C
CМ 8x������kRH}W�N�g�׆j5��r	�o	��oG0���n�+w�.m�m�k���v)�1=�rH�޽�

��[�6�u���I�$�N�Q/D;M�:��[{aq�'�ct�AGF�V�;�q� R�-M���=F���Dh�����99�/��R�S�Lv;e����P	N���7���y��}�JF�
��ez:�ȁ��K�U�M�}osݎ��-+�S80���#�@yW,g��1�[e�G�'c�0r۫5�ᙚ#MY���$sy	!}dN�����Ͱ�F��L�f�L�(����uǢ���]�_���E�}��Ш[V�Q�A)�J�7��f�H~kCE+!�����O���R�^�:|*�)�5M���1v�ᝏ���X�顗�k�J+C�y�9:�V�P;��>������� +T{���ܮ�����4!mFR�m�R~a(,�E�׬/y�=�ǉ�I�}��� ���Ň���5s�U�zv��(%m@��*���z}��G��������d�9~?�dm�QQ�����K\�^������ �u���I4ǧ���<��ݲjfĻt����aO]��˂^�^q]z��ha�>9M��ENl+r��r����>�%��n=��<4�d��ÂMp�?H��a��Jx2�2$0������ݜW��cY�����LM��<��D���u���s�Ev��֤�e�]�SN�
SV@wN����������]�������K��cV�5�Z��s�cH�"�3b�?���-Q+!��Ԓi7~ܿɚ�(�O1k����d�����6�7oVp�t+�Ԇ(�f�j�)�s�[+���dz�w3�m��i�0I��D�]>��WɊ��>9��.�b����:@]���:�Wo�dC��F�����f��^�h2��
/��3�n|�U]��@���,�
m*�SF���e�[��L&U����U�����n��vhi�[5{�N���	�/�Ci�N.]B7V�ں�Bl�["}����Z٤�Vq�_�4�'�}�sÿ́�/ꬎ3��:;6げ8ͧ�i�}Mz�V�q#�M�Q92.��B�A�t�"���X�U0�|&j.!���6�9�����>��x�K��{Ұ���4�ge汗�2���a/��$dlZ�!�&0F�>3ٮ��>Sغ
��o��kG�D�,��r'"���S$U����k?�{8�|��"�%̞@�|������x�᡺K�:��9n�,���x��f�����{�gTT[9%?,v����q�-��m�yC��u��îs�G�>���O�`eda��R]P�J�����޺�H��g���o,؋nQ������!J$�i��\ü��)��m�q�h���I�"�^jg�B��a5n�H���.�Q�B�Q�}�L{c`g���'y�{_���˥KTލ�Z�3�`X��YCA�k�#��d^�u>�����F�G�|NߵřW9m�|�kp�����F��#]"�OO����i}L$gyɛ�Mz��|y�;4~�CM�D��~��"��I�~�z	?<���ia?P�����@�P�Su�&��	������Y+A�&4x/L��c9��'�`�ܛm�6�ވ�s�ͅK�]�ohV	�ֽC��+ԃ��]�E�H�v��g7�O�Iņ�����{!�b��@W6��e�/z̽j��*ڋ��]Yq�?KH(;��� g`N�+�Fy��ɪD�M�S8����]�PF�����V��0x���	�c�����*}R���Cٳ3�շ�E�f�'��RsaĚC�^¹���3��:�+�"�`��ܫ�U=��vC¼=�x T4�HcǦ�ڡ�MDZ��l]b�՘T]���c��҂)٥׌ԋ��g�V�j<
i�☤��9(A����켭Cʹ�<�u}����+�Fl���&��k��ĥ�|��3�m��^*]�X���*S&D�r�F:�ۦ�����z�kH�����Y���!�lq�4]= :�2:�j�zU��QG�I��k8-H�q�j��=�G.LH\I��l$�t�囈^坤�ͧ:���E-�ʾ�B�H��@������r���G��,���7e�5:*�f	�B5m��S���WL{ۛ��1�ٮ��[Vx�G ö��m���;M���3�2N����L.-�v��Є�,b�U��, ؊y>��]�%�s����.'e����7�A6��/K��Ӧ���9���j��C u�j9�)��
�H-�Yl�j��;���qc�ǀGr���90$�wi���dɅ�&_Z�eYwn��vZr�����O��bJ�!z,���ʪ�Ɯ�{a�ZrY�*_<��7��yz�k5��A�,�т�����ƂJ��n���C��*���ث:��e�n�'>;P�z���
}s�2��k��94�u㾀��ﲒ�x{�\�[}me���dI���y��ݢ�Zeב�!p�v���8� �~6;1�����a�1ΩX��`�Oa�e�lvxq��PFí�ur@�H�q�Tb�I�C5��6ӫm0n
���3a�9�d��{,�kV�����F*m��u����ע��g6m��+b�m�9qͺ��+S�����1͘�
Z�NC{�9l��f��(��6��R��fj�G�9y����s{�]�^X5�]�9+8�����1�M����]J�ë��e�qW*59tCJZ�;�l���uG�Eś�AJ�37,T�p�9n��5k��a���oN����Ox�w��hT�]-A�i�D�)Z�,�"f�(�=��e�fVn��y�^�0łu`/���_.�/vp�m�BC����`nA<�����f�q�w]�N߹�c�`� �MY��t���^-k���o7��yt�u�Ǆ9S1؜z���-��k���[�DD�/M��FA��Ѷ�֥5�U��AX����]+����;{���ml�*�ǋ9�����ペ�n�^����g��&��2���e�Χ|�)vz�7L�hN��k�Hg������u�W'A6��Z�^��`�����:ײ�۠u�M�/z>t� ��ղ�Ef�!2��	ݛ�����^}��bt���]����&��	jD�W�=�∪"-Iz|�P^��.I]8�^s�󓏏������}u������EQ��8O�xd#ܨ�$	R/
����y�Z^t�~{"�<ν��y�w��q��������DS�9��ܫ�#u��AxQQA�H����%o+���~���x��q�____�>��U6�%���kU�FȨ��"��2t��Í���;��߻w����}}}}q�Y�.r���N����(�ʼ�()��Y'*s�&�9rx��������q������=����O�EN^�B"�1"��%�G�Ǘ|�o(���p��:��x��������?]}}q�Y�އ�Q{p+�9+$y�G�+�G�U�U,��T^Uy��H�G�r��$U�><DV�&�DX����'d0�*Ċ
/}z�~�j�B*r�<zH��U�Qy�_HEx�'*��B
r�/t�<c^���6w(6(D�@lEU^yA,�'�=��CN�h1�j�38��.�ҷA\Q����B/�.J7�GhAv�Kv�e���HLp4!I�"`�/�v��;�N���Ӎ)�OM♕],ᝎ<љ�n�M{�;"�z�2-A:rV�V�/icq�h�R"�`��"�
B�IЗ�[R�����Jk��gMƓs],�K)l]%v�m��Ձ�����ɢ��̻b�s͑�]�n�l,�Ĉƚk*ˣa�%՛#����k�+4��RL��T�ӎ���t:Fa��$hS3�}s�PF�l(H�)P�	?@����OF7Y�X���G:E�u��c���ql���[��q���}|��f�h�hǝ�����[��j��أ�Sh�y(U�̐C�֭�Z�.}j��Y�ʭ��*?o�>H~ a��iP� O6�`/�Έ2���}�	�Z��9QM�w�$��G'��KPvR�/�b�x��)���c],�L�^�C�ߩ����q��w�jP���R|��8��Xh�f2Z��q�R��ⵊ����w�Mr��Z��C�nhn{+���y=�3���$��|#��D�Q\��oF���h{+�bW8s@J��Dw'�O�V=�f[z� >v�3S�{�7!�l��7�x0&�w��X�"�W�<�RDx��;W���ǧ뮹�����r����E�-�.����9�pd����E4���`5�����L�~-������+�r���Z�*V�H�f����W��'M��$���f~>�p�<(HO\�mg�8�˲l���v�q��!Ǌ��7������!�ޏd���_�6�h.d+y.Gru^������j�Y��5|������mC�?q���gVo(7y�Uk��j�yj��DEs�d�mxiBޙC���/�Ӕ��o�3}��:Uy�a�wy{CA���4D%��Z�) ������������ҿ��d!�x�x���u�;_��	D�wG�����č����s��ZZXq&rz��*]��h�3�¹�S���k*��=�����[7�5����4�Y�o[R��lNv��3�l�A�\Ike�b%Ǣ=/$v�����K@��'[ ,z�a��2v����,���sz�Գ���گ5e�-�*��
^V���.��:3־�����C�E��pz�����ZZ�Tk8��B��Q�:A�{f�hn��;&��^m�G��Ov����-��f���v�\��*�T�%9�fջg�������i4k���6����D���̨�+���ˏ>�� �fn	9k�=�'!,p+XNF�ƥ�~=�&�R�Jh�3�W=����N<����Zx��}��yǌ�e'�n�4�#��y�4�2Ƥ}b̊遝/�&��{��sTSWS�v��#��{�a�!��݆1Z��c%�6�����6r��ٹ��1��Lv��fd�Y����ҙ�ǝ�ޕ9�0sBu�ZEK��ݱ��Z7s�<C����J ���j�:��c��xz�3�Q�޿w'��e�k�ws��as�7&
�2�;���i���-N��d}W�����v��;�w2�b�q=|&Ӽ}R�koz;��XZ8uT��A+|j#ٌU��6p�����C$1�<L��=@~xml7Fo~��_y@h)1��?���ϛ5�>e�B[K�ֳ�F�TYQ��Gm�@�NS_k�P]zۼ���N���\��7w��a�>�`&�&�i���J<��f�/�VJ�ε��9�k ?H��$�c;�ey5 ����rڪ��`���q8���ߊ#玲���C��9Ϝ޷�V@��l����lֲ;����x�ƹ�����h������J�:��C�@Z\���{�pp�K�'p'�_<��i�m�y7�&�	�t"��69f;��Q������@��+E�҅����).$��}'e�/ [GA���R�ѝ����R��k�灵1Z�������}6��v��~vY�	���������f�"]@����ozm٧��L�l�;q��<�T���3�$Cl<KI	�+{��I������e��`c �@ͩ�7��!��iSttv��#}��JQE7���j�i�6����Y�������g@@���1���m܍��L%�ܱ3ʉ|��f�a�-�ڃ��Y�L_�7(LM����7�)�m;�,T\&v����lt*c�l;�å�oOb����k���t�Ul>���G�Mvi�\�vD�:���'Bs�O5�q�Z6S�BWh�v���7Y-�s�˶ﯧ��2���0���x2�/'����,@wjq(�W����2�5��������ԛرwe�M]���yTt3��vWg �����T�8�`��Yc�%���[�K�O������ӭke{���\EXn���[�L3�13՜9Cֻ���j�x�fNe����s`2�D^C��j����.ZR���k�[<z�(�e���\�5�c�׍�����kJhM� қ�q����6���X%;F�}<��Zh8o���$�w��X�/�z$��b����ázWr�21iɅ^:��o�cZ�M��,5�j�'��hp{���Q-�ˎ��w��v�D=k9s��@>��R.��[׹���f7�Al�A�T�[�Pk	�-����B��p��tDm WH���L5�O���a"����_s?0�.8��}�]�I�t�B8^f�ip�8nP�ύ`��|p��
�_�u�g��y��,�w��܍B)�	%�E�l�,ь婓7����r~���L~U��<̈��S+
H)�ؘƘ�|2D^F��U��?`�������V�Du��}������<�֗���v ���e�X�m����wm�j�����6�+A���ܭ[��TY�6+�i\�]-{��T~0C$2Cz��t<��{���([l����B$#�>�m�h�ȋ	�S㮡l�<��I8~������lQ~i�ö439��H�n��}�}��'K�.|�Y{�u�Z��P���
ww����g��,��\i\���*!Vl�l�vC9aK����A����"��wXo��ym�ۃ�J�R-c+���9���k\����Qn��i0�/�<���h�s�>ޛ�7��\�C¨g
��lE_[Se'N�$�<�2ĉ2#�l ?��=��潑�r�;��TQMz��"]%y��,3]U~�!Omn%Y^Xўܥ�u�0�vn���޵V�l�=L5I员�s��/��J�͉*��։��j0� �y���.�N8�=M�s	���̌ݷz��(��So7]�>����j���k���_y���e�~����f��:dC:�A�e�3Ϛ�WF�]�@|��-�ܭ�c$�t繵��A����^��ew\�j	���jtqW� �'ac������Ƿ���}��ǿ��1�7G��:���I�X(qojݦ�s�;�ѷ׬m�Lv�jV��*m�y�ٓ�|u���`���Ԫ����T�Qt]
/�KW׎��.�b�uK�J�w��i���t�iu���O����G��Cp��2n9߷l�{���0ޒ3k�5��h8Z��ե���uuǡڪ��*��#�:ݺ���
�5;�	.�`�`c�'5�|y�g:o�-�4=d0-�5F��X k�cWan�5o���=������d�5���pm���ϖ���V�R��d��O/;}��l��L	�d�ͼ�q�gD_���}��k��@b�Wm��{_^��.�ƻ�x'%t	��*avw�8�/�q�0�2�ECA�h,�]�P�*{%wF(���f��\yN����#ɸ3��b8���Hm�nl\�����V��r̶L��$�h�_ʍr�5�7!]wV8��E��_gQ5����y��oE� �|�w[���9��� !<I���c.І���M���Ҫ��ɣ���c_rޕ=WY��v�4+S2wz�E'�g8|�釢�z�C3�	�'��q�{k3=T�+���S�8n��`��/�A��ػ��J,���b�c�?36'E#����gi�<��kfcr����%��g�n�!5��(�k��P9S��\�k�qfe+s�����ʽ'�#O��@E��u��V�S����v��r�j�ֶ4jݫM�o��q��ƻt���Au��2_<�w�������Fo˧�~������!�`8�4�����?>��[��/�MUĂ��n���јԛ���ȥJ$�'��峵�f�N_��_-Y�q�'�Ҿދ2��[��%���r�21��p$sJlĠiS��u@��bҭ�Ld�I[����$Tҁ�C�Q�;�Ʊ8��X�Z�B�����U�Z�TM���Q���v��m#�Ű�ã*3�u��Zq��4��G��Z~|�;7!4�vm0�r�4�Ǥ ����4�����p�s�P��-���������ΑM�}R���u3����jx\D��}���鼏T�F��ioV'���dx�0�ϸ�/W+]8�cl�; �(����[�$�m�#��g{y��b�Mo�C��1؁˯9�^�9��7���Pl����"���L[d~�K��Aץ=�~>��&$�`��,�qIE��|�plb���C�� 7NM&��z���;�y�m��iO&qӱe�[Nն�W,/�����
CJ��	����MY�Հ��EE	[��\O}Z�	1�����%�$�tƧd���Z/Ef��F!�J؃M\[7H-�Tc�]�3���Q
�%�^��E�,�q��5*���}�ޓ���� T��E.��Y�u�ם���Bd0��])�ݬ���,��+!��y�|ߟ~g;�o>��~��<�\� �#�<X���*�ԙ!�aA?U ����ܼw��>�J\T���L~U��n�es�jBm�2}pqD��z�H4����ٚ;"���5�_�Ǯ}o~��d<�Au�;�e?7��˦��!�1%��t���{1m����C6�N�K#i 3썩�;Vnx����N�zl6E�Yr��q���s���S���	n;m8���g��C�(�o
��%����8�3�M�ղ�{/�}��{.z�-dL�5�|�����'����,Ԛi]�x���_��q{dܽ8�|u��U_��d�Q~Ơ!��S��ϙ&�k�}M:�V6lźМ$�m���^�������m���v�3Qq���A���zWG���Έ�wbE��N]*\�ei�d%TaU��u'�`�;�6b�Z��`K8�����ѭ�f��/��ʢ�f�ER����:j,��nƞW�ޞ"q=�����a1��n���f��9�}=�9�#oz���3{>�}�)�4j^��bz8���Q�E󓱎�f�)��j�k���Sf7[��Ҳ�(���G؛���;�$6a�^%��z�V�`��w�D���ݟ|��Jv߸}\�_A�'V�{\6��E5�\:�njƊ���`�����nA:��n��n�Z�����οK�a��80�CD��?�m3ݹD����G���ٗ��%P�F�q�D2E�^�a+�f�9�b���f�%y��/	�����}'��4�v)^�η�W83�FO�y��!�E�:��t��m�e�D�qE�-���Јpp�{�x���&	�����3c;8��6َ�kN�׫��,P l�J,��3i����9)��N�z7�wm�Ӻg�A�ݭ�D���L-�0�4c9c�=>w���f(J������le����'GEH�S�7�%M"W5�Q���4j��cInn�vƁ��\�=A����N)�_Nvi�|��/:<����1|@�E���r�q��,����]?y�({���s�RhP�罫Z�Ir�ӫg!{ZlSѨR���`׮8����kγ;*�V$$�{f*��D�6P�Ɗ>s��Tz�Y�	�Lv�SH��w���h��$���*�����]�U
	����V����<���JM8�Srm���p�^��X��T&�{j�m'26W���Cz������O�
��B���H�EyX�	ǋ&Oa��ݕ�]Ҟ�ߎ�Xn{a�VaAv�p� 6X2�}��{�Uݓk�j(wi$��e����"�fufÑr)=�_:�5o�+���7~go*\�5���ݜV����t>Q��x��{����M�؋lgJ�+����33Q����][D�|����(���� 0,<|<Gn��J���� ��Q\�D�ra�蒣Ң��݋7��LP-F98�� 8ȹOC�w�Sw�2� ���ca�·�y�&�ɀÚ����N�k��.=�ᅧ��r1���S��Vp�����}�7��L���-�!����}�R{:x�o�u�\�̒�Q�;ev��jB�i�!��'��.�X�pS���Տn��,�e��>�ѻm����1�+X`2(���t74�h�Fa��k׃Bӣg�l����	�ț��Z�м��c�H � ��e�`4ΓO���o���I�����W?U�^m�TQ`R�k��u�eP�O��&��s��/��#��~y�q��6�љWf-h�P���\�DY%sy���8��<��ZEC��ru̸bWO`���y��Zy�&�z�G�=�3ŇѾp��z4�����3aj�,�ו����5ILp�sъ;R�r���o��%�\�����G�.���{��z~����0���X*:Q�O��,,'�����!�u��\D�٩���`�X�u���XN�V�kNi�� �m�Ox��6�SH��m�wUb�$mL��Һ����R���n�c���j�sb�Y<�oR*/��4_[�7�iat��͢^+�d��3�'�n�k�鶳�}�W��%���Eu����r�4;F:�S�lg�r��y���;�����ԞD{S����l��pvq�����.3����o4��}f�ȕ�ME�Bu�W`�S�w**�4��E
�ò>��l���_�:��bM�J�!uU�Y[w�a�o̊��.nI�YRd�肓�ݤ{'lS�[��ɖ���ț����)�(�|������Z�o
e��<m;�{��~U9�,���IR>�o47KUʷ)ڱ]ڕ���iY��m��ԣK�Mʬ3SΆ��+<�S�&pW����)���`y�jL,��U�Z��1ۼv�����dԖeP⫵%���]�@J��]q��H��)�)�*�}��ɮ��\�I�Y�3*4��g�l�{�Ob\)Cס��,�T&�TC���6�gV����]����n�Rk�h�����Ole#��zp��ȫay���k˿|��B�N���Ob�`�F,4���15e�G�@&�� �tlK,bc��h�.�ͺ.ƈL�CD��?dR�y�٢̅Ir�\R�As�dm
T�>��С�+�\z�4L��_3n�Z��
�V���>�\�t���7M�Knq��>�j�6+$gtH�j �0�E�g��a�Z��KS1���Oq��
���8M��չ�!R)�k��km"��7}�9\��.}�s�87+pLS���GL2��ӊ�U;�샭D��3���λ��#��5�^-I,�p�/׺Nl�kk�Y�-��:�[]�i�۰�p%�p�ͳe w4�n]�n҃k�㩬wт=zE�DR��&��GNc��3���{;9�[��{ Xа]ꤶƾ�������o����#�����c�Ҋc@QS���ðv��*��g1oS�a���2[���N����m�/7%�d��	kw��e�`:�n�=��
3�ZM��i��|��_��1�[��f˾�����j��8Ӻ煙0mM�Y1s�V��mT�a�#�������0]Ԝ-�X����1��4d�;��}�][&���C�/�'9T��m�چ���������<��x��O�ћ�Γ��w+.*+ʜ�
i%16�}2A�6^�d�-e��!y����C*�l���>S�U>0E�C�d�(�!��_@^�V���	Ԕ�QO~?�ӎ:����ϯO*yyu1-��������P^�AU�S��Uǧ������\q�����Ͻ8U�C��()a9E^�jy`����s©���߻�n�|~�������ϯۏW*Z0V{�$��XJ�T�wK8�'����.����hz}|}{||||u�믯�����9ɪZ��u�¢)�!�Y:�I���$ER0y$�+$�����v�]�y�?}}}{}}}x���������r�J5J�
�"FEQEH�?H*��<�������������q��׷��ׁ�t^N�tG�0�$�i�t�bG��D��b*�X6NC�	u���
,�C�i�I+l��N�O�3ǈNy�zj��<��E��B���)Qz!Z�Q<��*�
*/[
�Aj��2tyEe�S�Ƚ��:���"w��T|��$UJǅ�����o��o;X�V�G��F��N�Pd�k��<�u�\��{x��� �x�!�d�p`M���u���_y�?o��TVύk��z*���tE�~�y�{`���4�v��6l�,ŵ&���P��C�a�Cu��ZY�34ܣ�Z�A��9�]@��kw$Pl�-r����������g�]ͤ�DȾEYf�ה�lU� 3Q��@�����T�"��b�Ɣ�6U�ݡ����V4�ѭ��<�Eđ�H�������5���&��l�_ͼ�J�Y�5�N��u��\�pe�����.X�Z�������MK8t�Bn9�p%g�M�sVNCP|4�6���P[TER��m�B*��96}ȗ��N�Q�������_=&��#Ǐu�W�]��KD���ڭ˲�jsZ��m�П; |siFw]��j��cnk�.wu�=�p��]�aՙW��[�����"�k
�����U�"�+��6=\o61{M�6�"�F�]r��V�+֔iJۣ�H<��{f�`�f�lֱ˚�-��d�
����gkEJ(.�>1DFMC�c�����L���N=d0�����7�f�1#u�����+k�d�Sǯlw�e;�^N��E+}K����F���S�-�k�V=/,�`��]�5%�Q�ً��(WC�8��a<��qj�~]���\�ef�.˱�ɍ5�Y��t��l0G�x��Ha!��y����矛���T�
D=cK�G��g0��A��z���ԩ�<�O�XcQ�eߩ�o���*�TS,��8A������j��ιz�k�/��G��F�W����|��[e�;�h�wbř��a���ɃJe�X�|��|A�!8e_�>@d�2�S�xY�:Z�yn��=����B�jr��K�HM֤3�/濠o���t{�ѡ���Y�)�_�7!aY�O�F��D�p�LyeH1�i~���ߟ59E�A<���QU�
5v�ݲ������uJ��v�%kIm���~�����f�gEW��C47Xw��N|b]�ū8�׻���N�U��6y]0
H_<��/��{���B{r(�8/��5�j`��p�٫e���Y��A>��3��}����3�1-�Lc?7N���J*�O�1����:�q�;��Wt�%R/��헢�q��$�Z!��4�}���A?�G��Jmn4ܟ���g.���?�wK�h���m��M~9^���������*c[����^5��Hm�BU�:ۏ��n�V[��[��{J[�Ņ=�qU0ͩ�(���d���Ӆ��^.�����U�@�{�ه虓�XW�1A�h�Ӌ��u�9_F:���₦�ao��I�W�b��z�c;��rn��� z�b<�M/�x?
(�AA2�P��5�?����h2��d�o�E��d�٭���%���ɪ����#ي�dD��ķ�|���u��I魩#���{�',k��'A����n����FrRO	ok�n�C��m9ͰȬ�(Ӳ���P�,"�+�+�5a!󉍀6�8p��b���+���U'��|O�Vf?����vTaͅ,/dpI���q���}�c?z3����˗�M�h/u�$�j���t>�٬0R~M<�u��Q�Y��:���!r����<��>"��,
�X�"5�CA�{�>�iG�e�����z���F�Ƹne�Զ�5�:��_��A�]�t�`��f=�m��0��]���^��v���K'p#ِ ��9�p�/��"����&O�dSU�[�O��;4��a�/{S�x6�<��V�}�5Gw�C���3���w��)�y�Ц���ri،x�oh��?fs�1���(P�Ȕ��"����9o�d�����	�Ow(_�ZV��m�m�7��f)��^�'�N�y����{a�5� Q��3�⫑ ��\��%0�W��\#�I�?L�b�v���1z�����]�ҍ�}{Y�9���Z�Զs�]�z-�Lյ�O~9��:y�)%�{�����C}�!�]y�|�<�l�-�|x6�k�]��/�ݵ{I���6���]C���\�Uff�������"��{��,脜���>�1�dC|�L����}�u$��<�s}��r�DKx`g��cy\&vT��d�$���A�����3��!������+#uH|Ż�Z弴�P�r&r�)ݧU���iX4|	ߕP������[ʽ�x,I�M�-���n��A�m�y+|�,��OL�&��9"s�3E	l�VktCĂ�uj�<G��	ƈ�I��N��h�J(��ٷh~3����$;;�ԽS�^�%r���ӂ��c	�p4�)����#�u6�p��\ei�ˣ�eӋ�u_o���(���$����3a���F���%F����Pi�[k�ʛ�f4��ȴ.�Ža���fv�f^~�L�B��A8��[ tA�h��4��4hCM��p��c����M]�7�o��9��"���\��
3Z�4"��3|�j��.S���H4�㶼6 �x��F�|Q ���0�k���`����T�Mv����MI�����4#��]�%O�cȨ]�k<��~�����^�Ib�y��G9��2�J�壗��s�@�o�>G~���ف��q���X%��x+i�ir/�p�:���-�H��� ��}믜�_>�^oQ����a�=*��I�!K�0��`;�1��c1؝}G�y��G���Q"q������T�֝�\�CMo��k����2(�k��qD<��oj߼ߋ�_��/وM�K�>a�mg��ꏷ$��9j���0X�I��]��7����������4��^�����@}g<���2t{�iX?���O������L��p��v�F�ʇ���xLC�N�
�"��{).�M����ܘ����k���쬹dT律��W��tM�Cd�SWˉuD�%o��U_�~�Ā��W����~�w璈D_��\r�{Z 7�FOl�b=zʊ�l?��=v�N���/}��ư4���N(3l0��;[
�������	�-<C{P�$�Gi�4st���$�-)=3�[�[ ��C	$�>6�ᬬN��a'@��� F6��v!���D[�u��V�q�R)_�ϵS�5ll�����vW���6*ן�Y5lC6���hN@'�|8F��骐�}���M����6�oj]!f�ݹ��I��ސ��.��V;�aǍ%��O��R~����^��S��s7������O㊧g��ugF8��sD����b.=����)i�&V�8�M�tT�({��<������1|[���?]g+��0���~k�p�"�cu@�e���
u!a�����6l�K/,};=��t�f�;Y`3p��l�^_����x�N��s�	���כ�����`k�"d6S�Q;�m�z��ٙ�ug�M߳	�`�:O�c�KB�S֠H�w�����f�E�(Z�{{2��_�foFP��W������^m|�Wg�����S��5�/;ܢ��G�;�f��V���2�L�l�""!S]s]K�#x��t��+f�����/_�+a��5�B���*K^�`�Y�	^>�d0��k�`�z|'fV�����l���r!��vjq����^�ϝ��{����S�U���F� �*Rd�^`]h�����Z�u���`�;^��ɞ�s�29�YV�rw��޼�3Ֆ�HaT��	��%�9�+J�p ���򦩢�I�lo~^�Wmݍ�՗;���{A�1\�:��80���C�O_ɗ�A^�Z(q%�������~_1Aβ;���)�ԙ�u�L���VZ����p��c{M�Ɍ������/��h
���#�G�� yÇ�f�H��R�(�����ߒ�#��!��8�Yi$�.`Ҕ�Y	bY��R�������>��Sο��m�T���ț��9�Z�{��MZ����u��֯���`bN�p'��{�}�;�{�MI��ow8�ncw?`|��v n�$��bnY��nzeԖ��u|��۹[�����
m��=��P5�/�D O�r�Su�`h����k�V[������k���VU��*nuS��9wΥ��R�#jj��.�*��z��޵����]˻WJddm�פ6��5���y�07[��g����\�y]я�V�g����r��/�{�c����%�C�[���P�&	�΄�Ȯw��ؕ�}���.���ñ�1�> =��P�����_��d�?{3��o������W�iM����w0���'t�55����"9�9U[����9��-�������]�w�/�x۝\?]9�힏Uq��f@�L8�϶$ԐD9�a�O3\��|�����[R�K�v�f-sf���p��n�-�k+�y�3����HjQ��Dt��WKxn���EBc�/'#����ij�1����y �#�߿��KKS��' ���{:FǪ���r��غ}"�U.����N�}��QY�z�ռUH'�`[J����a�zAq�i{|����oL�qx�^i�16�`��������r���h�ٰݣ'��~�����;̽A�]�nT^.^}�g��\�3�p�δ8���%�d�M�h�H��e��5sP^ԃF87V6?z���V�ׯ�\ıvjĘ�Y��$�.l�i�����O��b]'0��]�����]� m�ȉ$�����@z.8u�R�E)f���- �؟$�U��$�hY5�z�
A_�ַv��ؕ�/�s�t������]�m��rÁ>��\��ܜ遮#��w7m��ݭ�Q*w�#Uמ��І&!�ĥεL�+�<�w��˧6k��f�`TwSC�I~	ƹHA��}�d�ܒg�<�6I�]5'#Ԇk���f䭨կ��U	+�th������:l�c;�C_��A�E�ϝԡ��c�F�����s`!A�'х�uu�Ή�[�����s>�y�{����>�>uZ\�_�v#Řy�a��e�*�G|���-�d�ff��Xj��1����3ea�vX������o�V�EO�.g���ez]W�&��ET`�r����d��Ay����Լ�u�L���0���;�� �<7z�H�`��[�ݮ���Y�Գ��jcw3��i�|F�ōu���Ѥ������5v8wp�D"�H.�yOۻ�շT{gѢv�^��ICuWU�yT��ʻ,�u�0z������@�O����s���*0Wn�!��;�������&w@��P��*�(o��ٽ�09Fx�z�l�뭳}���f�C�V�����3ʹ{*�Z�.�ɵ��;M��F����aJ�A�$�ztb-�S��P�3Ga,[K&A�s�ɥ3v&���B��t��_\�@�_�S&���<�x��g����2��Z���'=u'����D��P���.v��4Z|�9�w(��|+w�o�o~v}��>�-Z�C��$�:�ؠt9kH�j]�.6M�Iv��fq����Wk��3���V�'@���a\E��oF>�e�(W��!��z�0�'knVr�O�x�	��v����OW�^z���\����	O���q�ig᫧$[>z=+o�ﲻ�S�_��R�(��,�ӤRy��Z����wS�$%���:��޿`������l��8��sVdC'OY�R�-֞��w�U��O���x��q8FI\z�Vם5K"v����T\��\��uud��YG�� o�v�����3�j�e�뱺z��;;�Q��Or���������*0Mn�y[��nX�r+bی\�|8U=���� doG��/U���b��8���-����O��aZ�1�y�yѾ׬��œZ�ofT�wg�=�k p�V��t�~�kY�M�{W�K-�~1lI`[*;��;��~�7ݜ;']I��0� wt_tsߗ���-#���Q�J쮾l�7��^�� *��ӑ��>2�z�Y��E��Z���>�ӑ��gWL�i��M�5��@Tp,�r��+���3׍��UM�����Kʌwn	�����Wg��E뮩�}\�
�;e+���+d�A!sS�{j:S���m<�kpL�B�PX���ۈ����|hM�o��������[e�+]�2��\`�pھOr�\N[�����B�u�΢��/����w�nXXH4�ov�[c��'=�X��	�ui69a%�@-T�d��o<�#�-KZu�ނ�)G�����^�D�xo.$�6Ɠ���@Wz�F��uź=�#��w<t��d�$��w"7ʂ�fόΩpR�����✻j�ٜ֠�-�{����ӝ���ұ�c�xLr�ږ�p��4Q�����a@�!���ǉ��g*L��(�J�Y>����6��JA�#6ҽ�:�ܰ�Gv�h�&np�ݥ�F�v.E��s�P�}`rui��+5��}�b�9mv	���ƚG�Fu�y���˧K��w]Ԛ�t+�Օ�,a�Uݳ�c+%�u��'�q�m_�Vh��8��� �#} �Z��w&�-��������޵�'ǹ\�ѯp�Rō�wDiݺ1�IA��NT����v���/�Z���%a�g�+�|���гm������eY���تf
V�٘Q@���"�rS��+6®�Æ@�%N�䢥!f���,d��\�ɚ���ݲ{�o/�@eLBv����j��M����+������YX�ĴT|��qWv��x=��>̾4a�������ۄ�&<�ڢ͙���_!�I���)�������ڸ�R�vj׫i�ƛ84��_a�ї܈�15��u���Ubg��7Kzt�{E@]��[eҢ�+U�fmN�9��pC�obG���"�V.�x��*��7:�j��/XY�9��)gpGX����_j�S˰E��Wv9�sc"{%_>�W�-N�]]{+N*zfތӄ�'Ą��i�L�{d�8s-[l6Y�����-e��:D��ٸ9K|^��`��j[����=�2�N�#��8��ι���}.��{���b��t����-�����p�~m*H�׀ﯘ�[�f.ss���jP��UW��p��u�7�cח�+�/r%-�T����e�]ݍ�Xg�u���>9�U�S���Qۣ�c�{yjYb�<44�gS�T0����)w��y��l�z��݋48U�M�:$MԮ�Q�Z��{^��ur|�Y���+7�x�����2���H$�	↡�I�DN�)��/T<����+�-�� �R#׼��w�����8�}}{}}}c���8yΤ�9�H��bS�x|��X',�R]]<q�q�����믯o���?�gՋgD�?'G�i��@xDP�R���p�I�'��x���Ռ�I�����]㯎>>>>��}}{}}}f�B�^�� �����/��o׫�'G�N����(��9�r��\��������������������s�.�_x�%}1�r�� �
q9���E�2q�G��z�q�������}}}{}}}b���p��� �����(Oӹ�j�����y�OO�����oo����ק���(9sۯ����K�.G��.�`�I�~�[�q#|�U*/|I�ǉk焬@P�	Z�*�*��*<��D����<�^dG�^X=[-���x�s�PPCYS��x��L�W�2|;&B<)̈́N��Z�^S�V<�TDX�)ų�
T�^A{�[ϫs�c�W�~_{ˮ��vzM���H�e� ����ӱ��5�����M�1�NRc6XR$u�-��l�]-$,�Gk�`��,�pjUJ�5[�v�5}$A����Nݛ+
�x�2�[���A�-c�r��6��[�32��_(վ�]�؁?8��*OLe�M36nô�ˤ�.>[疒O]G��4�4'����I�$�Edn�VR�d���4e�Y\J�7��:��]%M��GU��,d��ݙ��)O.�\���2��͕[R	1�)���d�7b� �Дz�|��������u۩1��El�9��v��z���%�R���B[�M!
XG�KZ5Y�;fBd��k4*C1�Ѱ�Fh�"PrKEөm�@{��?��{k�7�-�+�<y�$8��B����kl�����v�'vkthqO�;���)x�5��E�,Y��p�Z�������*v��}k�d�Pȅ:�5H{�n�8_������"���63Tc���:԰�J2��ڽ�w`���փ��$W����������[�՟x.�n/i�2mOV�;5�u��Ĭ��7={i���xZ�V��Ay��5��7��9���fc��ޕs<7l��f^��h��R�,y�v�)\GCi���nhϯ�۹��_��-��٨;�O!����T�Y��`��(���k�����[4Y`n3l��L�g%T�꧀5�%�2��	���;i��C�ٵŷ��J��=���J�g.�,��2݄_6�vq�"�{2��mJ����bU�/�l���n�=���β�kvn���n��֍>���.lݨ-�9[|t>���A57ܬ�=��"��4T:����x�=��<��Φ#]�m��\�ƴ��ya���*�cl�X�(���y�c�ϋ7������g@����]!_yr�8���yF?ay�&EU��)}�S v_1�$�f~��n=s��f��v�%�b9�v�A�"�i>޷t�o/��Y�{�#@a�9�bp�4�Z@M��jg�g��Z͢�wq<C����@To��P�>��wEG;*-e呁���&*&�Wc���i\�����z�Q�g�w���1�E�wa��u�7i��F����<wu9SPW=���s���m�5��w��[1���;�(�&��D� ����)=SW+�Oo��.q�-юk�ve۰�l:f��u�N#y^O���U�)��1���֐�����I<�k\64���=���AJE۳���Hz�.��q�嵤�[�&�[8�Tm~gp���S�./��ώk�uDy�#��vU�O藫w�����L�w���m'�
�[�8�:q]�n���I6b�5�%�㠫�jO��_f���Ú�Q�H-�@V���J�T*j-�KA=�'s�{gR:*Q��^@�z��iW:[%k�˕KI��7��lf�v@S�=������m|뷑g�?sOE�|�ܕ̋�.0,s2�e�tǒl4Ǽ^.����Þ@V�!O�j9tJ�����-�lC`
o$7���rv5�F�nneOJ�A��ؕ�;h3Õܥ��
:�)�ٿc�<��֮Ј�Qy�Q}�Ex�8'���Ϻ�z���]9�6r�&Щ���)�}������%���}��ߎ'1��2xY����z5.L�xy��Mcx^�O\4c����-����	��;�W����;e�Vg۹�V����8�
�T{��`i,����I��<�S�����=Z�}���o���\��W>8�Or�mWq��7s�V�/M��[\{k�\�����}��_O����M�V�b�xI�׾��z%��[ُUoG�=���^��<[�w�q���2CB���W*�^m��v3�trS�+�äQ��4���M���������L�g��e��ݱ8�,Lj3��"_L+�����G��0Ews�nb�w�P�<p�WH;M9�����q��7;X,�'`=�@���+qB��L "�w��o�l:$���'aO� ������2��:����Ӭi�z=x1��x��bA�Y��8���34?�;�w�4�0�HL���V�tW�n�<� ����I�����B�tĵ���Y{ٷ÷qCG�vg�/���f�j���e�ԟ��{9F�nż�l0��^� ���}Ɍ�WI��~ҙm�?Xc�*饴3o?)G�%��+��g���X瞅\�R�a):�B��j���Ż�b��ؗmž+��~�.��6��X[6e�KNE�^�
�Gg1ĆuS��{l3�:��"�y��`��_!���KTVq�kC`�Ɏ���ڹ��7���F:�n�@O�-Xk{;b�x�'`�?��/dRJ1fG.��/�����9
��˞��um V���"��<;�����*�^�zs��߇��V�7Xb�y�wx��,/�|�_7_���(y\'L��T��Ǽ�til:L����e�:�'`��{�]�A��{�'TW[x�5�|�9>�Phot�����G�(���
a�#'̈́[~��}��زev�Ձ5�6�jf�l�Iz�k�I�^aGX�h���q>z�@~Mgc�^K2'�1W@�m�c�7�N$����n�~�~f�ًi͈آi��w�z�C���M�e����ߑt�:�l�����L8�^�Գa�Z��)r�]{Y���G0�\p��;k_��n�m��~�,�;���
vw�Ԫ}r_T����Sg&���3�^p~}R��f8��H����e8��Ǹ��u�0��n��~UX�����n`���	x��5����:�]�i��Li��0�d�v��X.҄ڨa���,gϢ���#v��@kl���v��&bq>]e���<y��/O�[ɽ��k`ǛvNs{3IdM��������,K �j���:���x�t�{�����ӂ�I�Y���r�
g��q�)���pD md3�����/��|�y���~�ƿ;TaN�>u:��٩�E��ވ+FX&���ܬ�^������b�l���:B����8I:0{� z����j�x��T�U�q�u�*"#Y�]��w2��e>}KvT�i�]�9fIu(��\qZ��M��ӥ� `�������I,2oz�������Ϯ�����1�4w*�h���d�>���S�Y���;U�B���1J�SO��1��z�<ʞpK��ӕr36c
��焽ʮە�Ws��T_t�ߴmK��A��|�6��b���7r��w��0!�a��w(�͍��r̅�I�y�.`���7��ٔ���u�h�]
��r�|ģ$ן�c�Hg�c�_j�;eN��5q����)=�l.Y�r�{P��au�+�&���;�ow�]yH��W�9�KS6�2���ҙo�2x*��zЮ�v������+sUΊ�eG��4�H���[>���C��a>�N>����I<bǬ��nz5���@��mȡ�y�k;8�r�bŻ(z�ۭ�k�UV���89�y`n�Y�1�����5�3m-��F�����v����5ǧ+�����D��������k�������|��tv7�9C�۾�4��Ϛ���}�q�3����7t�g;:��S:��r̗96_E�{�Ѵ�	ףG�~��CC ��Ͽ:�������%�晨ݴ+雭�����`���ކ�(��<+�[����mٞ�jpg:�Jw�/�,M��}��f�2��P`�">��y�z�\�"H���/���$��o��ѱ�x�/�!\�J��A{W,}���[��,�2�!g<�f)[/tӰ��Tv	�pcpΰx�]˯j��ط���OJY�+�bKƓ���oX_��f����=.���6��v��R�.&����U��vZ9��W9k[m�
���,;��[�uN�k�OM�L�R��ۍ�e��Q��c� ��޸��%�/V�-`兩<��d��s����7��G���B��^���H�M�-خ;��K(����L�~ꍧ莶���=�U�͖����$Y���� |yOd&�
f$�j�dĶ�j
�_��J���Td��Q��"�&��I�XГNz��t��ֺۭ9���B���k86��X� ��l�\��z�[�DS&��2c7݀�Z�W� �b\��!f��T�s�_j�����y�4%����<�{��!ު-�y*v��Y�ٙ��w�Q����a�0K6�'���ʈ{�iʯg�7���.��k6Ҙ�v>�Q�g�;Ӕ�����7]�a�߉f�QK����Cm�:�!��K:��m�����vWc�����M���0[]�'0�nK�_y���)+��Y�n����ݎ}�����xx3cdٽ}c�h�"��m��9JD�-����"��p�tחX�DXz��iŰ�1���z�~~N���QR�E�'��[�u�Ot���[z���'��E�r ��i�A�6���(G!83��:��'Q�~��^�p��~̃��Q��5���pyK14�r���6�e�6��(mx`VsB/�߆��;��k~�]R���(Z�dj��1�S�KЊ�-q�әl��ܨ	��N�@J�^�g՟6J��xֶ�CbÓ"*��t�ZM��|L.��R�Շ/Ѕ����q�"|=MCW��{v���ߨ��N��T���e�Y���B�˒���hy��5�ۘ��f,1;���o�s({��܈��>a�N�G]ͼ�
�V]|�n����ď<���?���*���3���Xi�����ɯ�����(��f �M��4�J^ɴ�WRu�Flg�.�Lr�BHNLd�n3���x~��ھ�Hw�)޻p��$��ϕR�&��}���qºT-��۸�i��2	*���X��w�V�[�LIme_V�30���������m�Q��\uS�я�|©g��T���g��\�`Z��+W|9u_������ɯmw;E�Òׄ�®l�g��s�w�@D��t�v�6�QuY��9��{����+��|ݼ�HUI*��ӽ�e�kV�����fl���t����.�W���OtH6I%���3�i���s�:����`�:d��X� ��6vs�k��2�מ{,-����qJ��&�fU���|=�3�3�(<O<�)�
l�ܐWJZܹ8��\�m�XPn�r�)<�����7��G[�yuJ:���3}�g�5�氆�@Wq�y��L��®��6��'�L�[���-^�M`��فZ��X�N��:n�8I!濒�ܶ��[F�9��CS.�*��F�R̔�2��Dy>�b�����ᙹ|��c�"��1�{1I�*�W����x�}�C�����L�]T�z�hp;�
��u�A�y�|�a�OV��^n6�WR���Y���fx�Z�[�{$��\�jGTQaeDL�h����7�|�	��w�G��U�����f��Ϣw��os>�c�],ϰP���!�-��L񽽶�t8l���A���u��W/^Y|1;o�}R"��ݵ	4��U��%��S�����z�ẙ��)��{����d�?�W����`�E+��dj����˹f,�bA���=�}��]��7�J���i��pf�L8���ל6lJaccF�y�Q�y��H4�@�oRd^Z���*K?X�Z���D_s��7�#S�����
ԍ��:��[��<��z�fV(�y�ѸX0
�d���y�-}����lzU�����[�8��)T[�L�"3m&�劕�.���;��*�NĉJR�C��H�˷G�����of�%3Mtj�V��vQ�I;Nv	�x�N�EG6rQS����+me�Ia�r�7d�*/0�z�`�,_�ۅP�����s����9�E��CZ�.�P�j�=ٓ��d��૷!v�oڭK]$���9�̾::�uFh���8Ő�z��t������}������� ��}�Ħm���qQ�f�,�+���D��&^XxJi޺+R�M��o_mɼh_���5V�9�4�e:'-�FG=������3����r�>+�V0��g/�s6i�	�wfh]�b��z��]�:g9�Ƭ�ge��j5DF.�d�QޜcQ�SiX�'�o>�]NM���+)i��ןl���Jm恹bc��\�;͐�u�&�p˒pK(�=��k;!�hͭ}7If18�۰.>�Z�i:�h���.�r'pTtNᾧ�6-��t���1�at��Dj)�M
�w��{p�>�ɪ��o9�s>�U�v� &��ğ������J�A���:�̑!u�A�g;W�M;�OZ��d�jcs+�V}{�On�4P�)= �v��|Q����*���I���4$j�׬�,��i{�`���yF�%x���:�6��s��2��-�vO-r��5LS��#W�I6�eU���P8�*����omwE�|J��Z%@-G���$t����K�~]��U}�n�v�sEFn�ٖ���<�!�S��eA
�"h�mNKF�*��=��ǔ��x짯~d�Σ�<��b4=���h��3+
�׳��-V����i}݂�/(���S8a��N4�w9�q�}׳v�qU/U_�)�;�J��Ӷ��x6�ǂ�Ճ�VaAӳ���Ӊ������G�W�fi/^��tOX��/Y���n���W�U��6�1VD'��Yn��=�;B��Ե�ݮ�\}��?R�܏x�DԶ[�7R��L�� G��A%�������F�ħ�zݥ
u��ԓ��T��,�t�0���Q���*F��#w8�(��*N㯵���6�eo��}&�	r��8�ܩr0͈2�G����^�1K�I���ŕlp���x�47B�ro\�4	jn��T՘bcnҢ������\�87z���b�Ks�Vs��Z�+淴[�o�j��S{.´�@��at��d�블��y��MPnPU!�16�Mrօ��E���x�a_��7�����,�T��f�.jbE]d�O�=��yj���6]2�Ac�ݬ*��qԬ�ђ���\��c18OG�(������XS��
Af�PIy�(�f�y���c쾒��9��p�9PtO$�Ƽ)�{{&�Ӑ�
���X���Ax����y�v{u�믯O�������qJ:��8+ EyI'2(F!#�@��~�N��������Ǐn>>>=���_���O�����z$�"�æ�)2�G!�`����*r9u'WDr
����������������߻� (��b,b)��VW4c++��!��Ay`������������������� �8Sʄz<��"7�)��B�dYm8�T}�<~��;��Z�$���,:}x����������ק���>�W:%	�G��"T�Q�`ȌT���P^�
5�9�&k�r���Q���Kʮེw��x�����}}}z}}}e���\�^�i��[�I'H�bD�|v�٫ ~��^N^�F=�p���AREQABHD���B����r�����c�f��YecR�uW	�[')�DZ�&n�=^�H�<�D�ZǤR�P^�*��G�VK���<��f�A߰�X,x���N��b���.��w��_\�fZ��Cy��\rNu�:�ͮ	��o;Lܒ���c9j�E���g6���bG�����<�1��q͒�y?��Vb�]]�����`��|Vӆ�ױ}1�Oς.��e.5���ޝ�ݷ�j��ʀso�9u��=6ºr�)��뉉J��*q��sW�	�ax����^q�g���X
茫� NvD敹q�"��U�F�ǽ���9'*q�g郴~n�gb?}��gv�����e6�=d�'��By���ܩ^�)w����K���v4�h2��^�󝥯��8Ɓ�5����]��
mLX� EQh�}����e/�.c7�/�_I5�U`��g�*�:�T�ǻU)ܓ��"`֞=�ct��r��cΡԞ�'��5X�Y���o^ˉ0��f_U�D��o%ࡄ`N9����UJ��,���>����ĭ�U���>�D�{g��6����Q��@��K ������{�#=x���:,���/�;��1s�o����a�]}{u6�tW:�w��Ø��xXx�a!��Q�B! ����*�s��*7ǔ��(�M*�<�,Sj�:u�ʙ:���Z�,��l��sD�L�Ts�C��=�=��$x�6�g����7�Ġ��7.Cv��x.�ޅ
*U(�����u���q�)@�i�xS����RY�saRq���{�*!����~E�릻e	I�$����73�Ζ�g:���c9��K���MO+v���E�i�ދ�5��v����.�j��x�W��aG���I����l!J�~��4�ۙ+��݄S�I�=����+�:���!)v��zǼѯ��[	��gpZ��t�	�������2��ayu�n$s�w��Y!s\� ��-��������A�����1�	���oK�i8ў�k7�ױ�<�w'/�y`'b{������;���Xc^���n�#Yy6H�B��ǷK0,��o֠P�O0��E�a�9�A�$m���D��@^��_��˘ﯳ̽����7�z�٘�Ok��w����_�͙*O
j������H��
���&%��qv��>�4S7���g|!w.F����.��^�Lޓ<ID]�EƐѐ��ϷgM���[�j�O�ne��r��+)��I�t9��c]n�J��z��ԝP�C��D�c��e4���߰��"��G�>�6LP�2�KfZXŬ�mo�y<���Hik��b����7h���nW���6ƺ���.L�9�����W>F:��/]>;B��=�'#��_\�CU(׈��b��W6�k�pkS�!�ܡ�:1�u�f6}��d]"���U�5w5�����M��L�.�oS=z�Zn����i��g�i���hڅ��dě�9��f��:���To3��d*fJcI�ƫ�r�󣫻׵��S��p&��z�<�	` 8��ыn�lTdp���W}�G�X�-�G�i<\��� �̓V�aV^�m���r8viq��-���8����r�6p[ͻ`��u�����}�o��?6�7F�����!~�=�w����9�Ԁ�������"I�饮�kbC)8f����xe;��5��濹� N�Y���}��<�!������%�<[�b&�H��9�/^t��������u�iL3�˗���W����D(��ߔԶ��p����׊�w.|���/�����>���+a.ͻ�VwK�Ќz;:��Øx~�G�$x�v�}��c\�A*�Pc�Q��QN����S����p8W�&n��n�� �Off�z���P�0����ޥw��;�D�'+�o;�^��}�]� n.���{�c�0x���L�PKu���Gg�S�D7>�F���p�=��d�v�ߺ�}N��c�X?ry�^� ;
�wsm2A�Ч���>31,(˱��V�xЪ<�3��{9ʹA�˪3��C��Wk<��]�S�g�ewU��S�?�J�K�k��� -5�H�-��	L�̀�ԁ�!�$5k���jI���D$�#n$�-�t� ����il����Q���Lc��뤽��@9��w���0���mmU��k^�{�B�Գ���}��L���3.2i�gT%Iq}����}�ۓQ��f�:k�����j�s�z���$���`,��yy�c.�swy���9{w�B씅�&Es.%u2�w_j��^42��bc� ��
5���7���֦`���Nm	�J�ɓ$R��'aU��og6z���}K�\�Ӝ��V����c̐��,��� ���5~3\+/���{�y�ZW��9��m{�Ҭ���5���;�o.dQ�̺Y�l�p��.H�\8�9�����J=�1wJB�f��}m=�N+�L{��2�yX"[�z���.q8�B��\�K�s����٩��Y�)�=$�T!��c�fy�.���E�mMI&�J�ҳ�'Y����֮���:�v'����j�;�1*^YԹZ�y�xM�@-ʀr�Om�{ި�Aa�2�<|����;`�mT�\�:Ǻ�ю�U���/0�ֽq�3M������tƫ��쾽���ɀ��U'�nnjͼ���zX��Z+(���g裓�����ίf��
ک��w�����Ϗ>9������KW1�-O�;���Ϊߧ�|�?-�Tl���5b��yG���2K�t���<����q�Z����z���f�� ���2�VF�M)O��|�������*���Yo��ז���/�A�J��p���(f�dT��t:ON:��Ԧ��@s�ZE��#��>继�>���}�=����%fx於�Ri+}w#�y��fi�*]}���k� �;�A��-�g��-㪽2�5v����P3o_m����9�]�����>2�ͮ��D
T͎Ē�(��'f񨧇׺ى޽~����]�����j6s�$���ٿ�{_�c5�[*u��D"ߧH1�ׄ�\	�`qܪ�޽���2��V��}[գy�j�fݿ6�4ל�E�`��E��Ȩ|���Fsz�۲�_b]Ւ��n�CS:����г]o0��fco]�S�j÷u�;zo�\o+�4�BrBl=x�i:b�����m�E^/H�J �1*0Tb�3����yZz�9I{�����ُS��^�����."q@�y��x���oq�Fu'�߆=�V�K�R�&6�v��eѼ|��s����.�S��D�����u|�GO�a���">��Bo���AM"��Ɏ�-Wǉ�G�`s�F�3�aӃr�����6u�kV��,dN\F�4���_��Ӕ�C�c}��B�il�~(��:�������F�h�TM�VM5�0��	d���[1����k�z�F��-�+�����"}�t�EF\��WyR�v6-[�uP�.X��Yğ_���R[��!VИ��Kϊ��k9u{64a.�b_w4Xw�^���ב D�)��.NG�9G�ՠ<�xR��0��Q��TD�R���D��ƴ�F����+�W��VRzk��yu1�6���������ʡ��r� �5��y	� ��+�mt�>�Ps��FU����w�
g\�qh���O���7���/�/{�2�:7u,����1�z����z`۩����IE�ڶ��1���ɧ�c��J��hY����1 �4Gj��l�#r�?r�����U���/���q��~~}��^��nh���p������&��kFٷμ藹o&}���~��vn@KԩL�}۹8H�C�G ^0�xZ���J˅%h%��o���x��5e�ESs!��]��kR��>�.cאb��]4�.[�֕Y9���t��sW<m�o3s��՚y����W���J��ۭh��.�nYj�3��K����%���=Dx׹V�/��������UW�Ȩ����
u��T'\>�	�Mw�\$�]���t��W��,�g,�K����ۨ��e:�&*,��o,���P�V���u.�5���˺s)s7����-�K6�b�a֠e���T�pͫdFJ��S,Q5�7�*wq����b7I1_F�����a����������2�)���N����/r<�Ʃ�w��y�P�4m�hN�r����f/���!ls���`^s|�Uw���^��GO0��S�{�� ����㦿N��űz?}۫��UDf�� Hy_Wյ�ab������_�w=ݍ��p���(P2XNu@�k���9�^�v�ٻ�y������w>��(�9�$�b��r&���r��	��CMn�+?fR���ٚ�m�[K 
�'����L����t��I��� (W�Q�m��������R�C��l.�� ��VY��������b�Я��A���su����\�fH>�k{ � ��'4�[oz�gH��\ѻ�8��|>#ц��/��I(�/�k
�+�'�w�G&~�߂I��{7�F]ʘ������7����J�f}�L���L� {�C�y}6�T�U<�e������<��ڮ����7��g���f��Ds�u�*~ja��yO�o��tG���">k�-���^������$��<�ߦ�"��m��萫�1�J�)|9-�2���*�n��tR��^�N!MGw]�Ց�f��Y裙��<@u��(T��;t�Zfp̖<M��9f&��46�������xğ����gkpҮs�-^���ek��J솶{���kf����o%;�)��33^��v��@M���Ϲ)�릈y�!?[�"�z�"wxgj�r̛�T^��-���� %���(M�;�Ll
�V4nϭ�j�����螃�t3��V���ᣏ~d۴���j��WV��Ō�:{E�<���A����`S�C�bw&�v&�gWmX���)F�d�"������σں�m��Co����۷.��2�/�[��t����̸��6^p'*�N��h�;b�'�@����{���3��������Dy�坏>��.f�X1Ud����1n�8���]���#�껧�ln*<s\f^l��s#'J���ά]�B�b��:D��f"}��+#�#��gX�U��k:�[=љ,|�ˌD�Pq¹����C���3���Y�d�������d�kUT�d�pg��.�է��rNཿ3��4�=�����y\�*�4�ͼ��2�]p	_
����:g��6��X�##T�6{�&bmӪ��ͻ�
��M0̀P���"{�uO���Ԃ�B+���4;����oWOtΑ�V�>��(��l����)ΟS�;�9�F\t�\eZ؈�s�ed���ʑ,2���l/����ў]�^%��(��)�k�OQ�ӽ��Z�LW':*,�8%���4�x��a��΅	a[U��*��ǹ�{��j�u����"Co���K���kIGct�S�^G��L@���۝J���2>[��:�>�]t��đ�p��UJ3���5@ڝ%�$z�9Dn�|�
@�Gm���pd�f��x�[\�!O���7�Z�ќ�=�V]Z���q�/�|mVS;z�-�]��qd�	]7��:M�Y.�b�Ч�V��̾�%jw6��į8�wnP}�{@�Ǉuȟй}�����!�Ӟ��-qFq�y�b0�-Q�q��]Eg���s�\s
��� �-Mi]cij���v�<��#4�s���]d��`*&K�v�������-|�-:~:���yZs��X����==Ƕu�Yg�H���ɱ���PĳXM�csD�oFd�?%w���{��8�ޱ�&1j�\]���T�� ��sjt���mi���̾&��k�������a�j���It������`�Lˎ�+�ә!��٧FiR���������r�e͋0,��I\�rx�F�%���54]u�M�N"��ȧ.\��:��-���!�GrX��V1�uY�a�ݹ5,�h�r3;�7lvƨe&y����%g�q��$W{V�����A"�ks{����(MU�.���f�NR�{m6Íy�VQj�	�E�B��/J�L�-6p�z��[
�A�n�{4�X�X�O��/Q��P�R�"m�ش�6����%���(b9�$[]Ju�\Y!�괉~��eL��K�:
�]�n�J�v1���(���ΨE2f`�x��SeVʒfm�F��.���}��dMz;�v��ڜ��c��թ�ީ��#U-`[xi��8ŋ��A�3G��x9�&����ӹ(�T.��k9�^-�v�ǜ�ʭ���Dn頫��۬��mi{��-��Rka���V ��ZhTw6=vY~�_-}O��t��o��EY��6Ѻʌ�떨��rԼ�vb��dd��^�f��X	��*�yd��R���Q�n
\Mv�nڹƓ�A:CT�b��[�6���}E]l;�4���ԭ��R��|kV�dL^����t�QY����{%�Mv�Ze���r���ڔ�wi��8�f%w2���l+�UΡ�5����C����d�%�s��<�;}�;/{�*˱;��ƶs,�pf��v��+o��Q/~��Q���${kn&��c;*u�}��&�V�G0)AXT�y,�m�L]qD�o*�{.�><#��U^ڗ���K�7tR�lC�Gk�G�L
��-����t��MKV�ڑ�2��fv:�؂̐[Y��Ж֝z-����-�V���d�]c��vi���/6�"u���]|ߙ~�}:�����<�\�O�è�~I������g�J�VBN�/0y۽��;��{g���=>���\���r�����#Ԓ#[E�%��!%�S�x[XQ�t!	r�������������������O.�=��b�џ�tz���
~�b2�	!<�Cb�$����s���ߏ�]}x������\�T���5��0��_m��ш����$�$yY9$��t���d��Ƿ��Ƿ��]}x����?H�yJ=�u,����TP$��dT�)^�UNT�:n�����������������/�RQy��'��k�t��aZ�N��/}N�Ƒ�;�nݏ���>�__^>���ױE]s�s��Mz��$dʶ>C����r����Ɩ�}M{��75��ǧ�x��u�%�XhAV�KQ����r�m��$�-��_RQE��t�pՑ�$���H�$��,#e�� Yh/��-�Q#�^���$a���:</
zHIF$W�C�Hύ��e�Ԩ���B��A��͸�;�:d���=f	-;H�1���ٵ���l�#�R������]��敍���2EAN#þ��`�G6�^�k���ßm�=���L�j0�'�bY�ˬZ��W�]}T��%�hv�R����=���.<�E���Mv�dƊ��M�d��� ��YM�v�vV��	߬O<���.I
�l��GWY�$eA��\0e�IY%�M�V+v.��biqfh��$³���Xl�=mi6n�j�Uf'Jk���4�IIuH���4�oѦd����;pp��$n�l��XLGa�M&���%�"���('!H�E�S3k�f̽��k�il���,���X32�Ȍ�v`�Ւ����^�gW-��7!����v�C�%ݥ�u��oj��^��(��}�͖���ƚ_H�!�Wc*ى�k�n��^�d�{3�2`��@�Z�3_2���d{�;w�v��f+���}�὏5�鴫��{��v�`�:e;D�t��f�Yd����>"9Պo.����Ўi��,�qz�%�2�*m�����yb����[���/i��V��;�����;:��z'*���f-���Yͫ�9�F7�u��r�3���*�6WEGUC����3;�N�p���֍[CZ#�������3�W�����x�����37��X%�!�H���HM�Ly�O��b�u8Z�fǵSx������|ݏ��o���N�&��y��I]⧐ ��9�{T�����q�&���*,�RoO��'�m<�}�˭������J>�����QFE	�Ϯ����m�� !���������������A�vг�nCq�����G�7ME��&�=Ի��\E���G�?�������55���iS^���A�}]Uu=/����3S�͜�0�r~�nK7���B}v
N����Kr+�Y꣠K���_3w��3߲㷒�US#�Q��eq��wW�W�8tЎ���n;�v�]fƷ�͹Q���{k��T�j�x۹�k�@@ed��OL�0V=�ԫ}����<7G�ː�?�X	/��iN���ө���z��V��g�b�5�K
�l	��a��U����^S�v{�%nӍ����g�Vj���\�pK�q�x1~~��^�L����]8��N�������䛷;W7"�^GYΚ܈�g�W����4���̹�/����cb=5�[:��k4�f�T�(�Ĭ�Ǵc{,1�q�<��1S#{)%1t�Se����-ͱ����t�~������ǋ��2�mjfb]kSEO&�j&��f��pH7��=L��9 �w|�d��8aj��p����VV2sj����^�#����}hG6���)�<��c�;�N��;���3G>*]�,Ln�������>[�L�؁I��> ��;�.������Q�ش�//zC���<F�����<�5�l�6�l���D�N'��9�hŻ���w���5��s���(ѣɛ��(z͊H#}� X>���9�} f����2X�gJ�|ئ��Gk����P�W뺼a\f��+����Ff>�c��D��x>�`K:3��2iKʊ.��]�m�P�:�>�>JU��\Z�Qz��h@��5��ēͲ�WS6�����>Jn�J/xXs�WNgl*{��w�>]cz�)�뢲��7ꦚwçC��)�;bֳu�@$�/t�f���s�,���*[iSH�:�4am����<���I�$�I �}�Y'W�Լ���V�dom���L��k,�fnHe^�R}�0z��f���2&������<c�)�(�:�ѝ���$M8�N<�ԵIU0#�0���;�{�W1����}��IK*�']��+�X��m#
�"!�_�����<�!����+K�����֜��6.H����ܥۜ�1Q�Mr_3z�w\���=�Is=����|��������K�k�G��W72���T�n�������n�u��y)��݊�s���72��o*�G���׭���G�C�_F��N����ֺ	G�Y���㏖�%���Ƶ�-���������l����z�V^���w���`I�#�k��6�����Z�[��V@s��2�b�OVz��?�@̧�]���dl���i*+*�9����o�H�`�vS� 㫠TV�W~vh��y[a2��C[����q�����B�;��g0�g�;�/t�7�M�40v��4!�����{U����������3�Uo����,�SE�f�hYvyL��*<������mCCv�^�N�x�~�*�m���w�g����K %{��z�v��9�^~B�sO��;�xi�z����i=&���u��ےJ�a�-h8&��Uu��ZВ�*��@���E�6��8�/��~�<�x3_gE��$����k�����q��r�rY8<Q}{�uK�;)U�O(^��܁��OeAE������R$�e�Ȫa�&uܞ��P�Fm�i��յ��ZX��j4�[-k(@م4�-�i����}�~�V��1<4����5ZU�ޢ��,ќnZ���-��zwq`x�q{ ��vjSEe�;1&A.6w�*:`uo��_�͍8t��^���:]�^��<�0��5��ޝP�-yz�˥��A=5����_k;>=wd�zr�W9�o����Ͳ��8%�5��q:��6�;c�H	c�]Y>~����l�\x\�d5�J�uy��O:�V�g^�Ժ��*���.z��B�̪hݕ��:�k]��<�!^@�Jvg*�R�M�C"�jw.5]��LG�=t5@�5� ZU��S�z`}��_����}�35�}#a� }����K��(06� |]N��S{T�DD�����ߛ�e�m�h��Пے�}lD��!��b��J�N������2i������x�=�YUm��	O5B�=�:��r��V���{��glJݞ�ՠ����>� �kJZ��=���62�u������5�d��m��BЈR�׼�ݣ1¤��N!�(����#��	�h�z��3h-��Ζ��y���G{	?��g!�=�����;%]bu�DGw0��A���*_w�{�u:�}5���Ѽ*�G8Pw�ר�v���TM[L�ĴX���#ڨ8��Z�5��7}�*�[y­x��蚘�O_]���ᱸ�]��}�w|}5�NА�k�k���A���[�ـ�Rت!�Q:2�h��.�U?A�w/\����ɛ�^���;�Y� ̿�'���NH��B�>e}28������{�	�JjȈh-��y��پ��fU��J�M����jp�GN-b�yc^�?�	���dz�UHX�=�*���@S�ۺ�H-z���%qk�9sي���^ct<���kTuw>�N�[l'��S�x��.V8����p��
<��{{�DU�r[�'�˪m��P�Ӓh=�ȁu��l�Oe�U���1s�{��hU�RѺa]N�m&���W
���i<�V�-�yYW�VVQ���w�C=1�s�e�Zlod���{!��}�YCa<9:�Λ	��9���ӍR�곝Ϣm��$iŋ�T���+9���y=OA�6z��:q)7�����_f.w�i�aFji���������}������_׿e��������Zd2�=�2�j�g.{�U+����m�,���{�>uͶ|�T$!7��\v�J�k�ᷗ��1�P2�wf�n��{����Xb�<<n��/����W����E� IE�K�ǋ\w�nG���W8�����?0�q��纜�+p�4Hݞ��yN��==�`��7{�/��z�vn8򾤄׻���a����xx^�<չ�B�l�h��oFo��`7m;QQ۷����-[b	;S��ɦk�G�/�o���h/�Z��>�ث|����� ���_�������c��ԴQ+��/]�F��K�u�͍��>�^-}��ٌ���Ϯy�9��
��5a$$�"��_�.���&zu�
�a�?=^���\J)+�p�sr:�-��³�������]E�E��1e������q�W�c�]�=׺�ظ:WV�L�i �1\9_]�����6�y�F���Ӄ��ʺ�O3�������cl�Nv�D���gxK�f��~��~�SQ�,��=T[�]��f�c45-،ˎnqy�qh��������j�uiM@�T�6
g�^�=�Estv�O���!H��I�~���p}�Ǭ�Z�+v���ʡ�jph��,!U=�^�x0�Q �1�G�t�V�;4�qx�*��5Uk�FT�n��^�fⲣkjv��	����4�[N�7x�v���w6�����v<�j;�5ج��|�-r�>U���y�~��=�w_ή�bW(�)PI�*�4\����Μ�b&�����y���[k�i5�|�z�1o��iTe��]��z��̠݇O����&���"qy�s�N����Ƶt���;O��x�v�X�ӯ�x��l:��kD[x��>t@qU�{�����ݾ&����-T�J���&M��96������o;�Prt�oΑ,p��6�b�W�v]�[�&gtT1I>�+2W�G_�6�x�(�ں�������FI�l�|��=]�-�яmd�u���f�Xd��b�,���
�����������'�,4�	�	 ��0�z�����|�L�Sm�B�Fu�TVn�����ζR!&��@$��oW
`�3?-��?�l?_�M����])��n�i������/�g�g'�݌n�O�9�@~NϞ�NᔌW�ϕmx�7nW�*��l��݇���_Vt��Ϧ�/��?cSw'wW-�~����l^�on{���ջE�t�1�O�9Ԧ���vG�!�Lz�MH�=xk�w@���D���M�/*�֜�gf�Mx㉞*BQ*��<�?���[�>pd�h&(Md����}uݵk����7������1��i��2e�n�dL3���L�����{��={���)�\�5fD�݁��4ME�xT[E&k���p���N���o-}|��ȥ���mcl5��>�=/��af�=��<RJ�ÛLU����V8��`z�Y�g�Ie�:&ϭw ��lk�dۜ���vKP�ok.�����i�݇��5���A��-�ɉ�-4��u�#�����b�Υ��s����Z6G	ܩ�z"���n����D�k(���9Bs��af���-�^��;J��h)��Gď$+v�2�s��@{@v� l
�s6@�]�z������2 ڪ����Q@�3"X�u�җF0�����,~��n�j���PXr��������m�hלv�G�b�u>��gt��U����j��nnk3�J��t^tmj>�"��z��b�0WwKQ����N�=5��8�o-ξ�/�;u5ϙ�`�#�C��*z�7e��Asη�M@;����{�{�<s�)�9�#%�*�CVj*�[�_Mf�bA&�A��$f�y�y�MuRa2w�[���~�ѽCvu��]��Ė�Yջf:,N�=Q*ic��Ǧm�^{9�Ԥk�?s��]]
z�<�'ܼ��{���kL�+� iه�q��Bi�;U��w���.�JO�=�}e{�;>~��g��=D�3� Ƹ-�L�V{}��z��iT1q 乧"ޭ�:���
F�p���ƱǮ�a,��P�޾�7�.������[�t_bR��7�G6^X8w{�]n�\q�PU��AƓ����ZLSO��u�V��r��6wuD5iW�Lܼ�][V�Z9<"V��<&"���0�-�]EK%�r�t.�滋w����L��t(��C�h]���b͌	OyP̲����ޝ�Q�{C���-A�a�kU�c�N�J�5��*�����g����'b{@����Y'K�D��A���pwV����}ӹW}�:�X��hN���m��PQ[ۮ8+�����U�\��㮙�n���1�f�C0n�un��WJr�n2��4����ys!�y�5[}A��������{�#��\�o��K9J�z�Pn�Sb�a
�$6��Y�
K���W�ʼ�y����jmJ۾�3�,�#!IΣ��L:��o{�]��
aG_$79eݽ����wYBv�����BQ�uYW�-��.��U�[�/�$R&�FbJ���dG���욖>ڭ�$����������p��W+�s�G:��攷U��>R�I�n���Q��c!Z��dtw��lƶ��d=#�`<��j����:LUj�n�δr��#!���v.�+��6�>ix�	��F+q��C��iV� ��yTn�Vc��Z�5��a�I���D���~t!b�fsN<H��ڢ/���˓T�^)�ʣ��=��I��G��y�z��̱�b�[���'+8Kԫn�	L`2�=�)3�����V^9��f*Bs����[l6��v���������Kz�&�M�ۼ����!í��7l)�B�[��]�,�o9�mijۿ�Ƕu��b�Ң[+@��7�����'ԦM�!�m����z+�6f�l��<5��\X�Nw�#��N*����8��ϋ:��Mkwj�ns��V48�є�\ɀǂ�m̩ۡ�R���)��H���	��b��S&͢�����-�*����x�n���#�C)�����fh�V3,����Q��Y��*�S�Ko#�1�%��a3䷪���S���)d|�:�ĸCǆvYgS����ۂ��	h-�n-��pd t4���X��
����V�2��\�l��)F���r�e����|�>J��ig4���1�VQ՝,�1���Rf�`��;U��r
	0�w���RULЕ�&�ʕ��%��_b��]`�O'ܸ��h���1���	H�,|ĸ��m�
|�u�+(-o^=t�\�� �._nѱ��B>`��$�Hx�.�}OM{��´���,�DlX�=>:��������������ב�?�Y	g|j��R �lP�ux����P��������������������������u�]�^{ueH�݇d�%Az�N�9p
��(�����������������~�
��l �A?Y��5=�$�鐏<�leh��g}s�Z��耺�QǷ�����������׏����
w�I屝��<��C���o���2�=!!G+��ק��������������$>�?��i=��d��� ��X�t���w��(�z#� �����S�v����������u��__By�*���驽�"TG�FO�}B�=)wUU� r�L�F�#dU��\��N+�v'BG�E� ��P�{J�\��c#!��2-��i���+�##I���y��DA2�:�o)��b�D �ǈN���i8Q��&뷯��;s��c�u���s��e�Քlk���,�/Û���0��em�k,��o����Uу�<=�|��'�o;s��|���E�R*�ҝ!*/5�e��(`�K
��7���YN�J���m�;�=n?���B�v�uy�z�U�V�J��۸�k�f�V�g$R۳{��fR�^M���\X|%��]O��?��\�N��S=�m@w�5�����e꽴��Q�^jZ��m�Աfp��ܩ����ܬZ��ӑV�t�(����n��=�8���>W���\nn�!'�k~}Ro1�O���}�����ʔY��{�3������f2W:�����$�]�t3�;Β���̩�o[y�4>f`o�+m��l� ����"��9��n�;~��㓱1ԙ��oN������zZ�gʨĻ{N�fO0��AΫH�����t^^�v�ow�t�.)8�j���b;D�i;et�}���wE6^0 �G��WS�u��;�~ZH'�z�����٬���}�þ��vo-����!�e�h��[�j��L"HOu��']��#r]i3ٶv.-6�E+�\�8o���g��r���r�ڜ���?��{����"��7<��;������y����<xCq�-Z�P��,&����q�.Y몞�M�-�8��w-��8�`�3��=c��H�>��F	�����o�6���NG� �e	=>�P��/��ݒ���9�T>�5_]�-�2q_O3��Hs��|Z{i�&6o���=l�탎*�֒!n�۫��w�yal�6�3v��^�K�Z!mn�vuE�S޺-tV��ftIf��x�[���6=�K0,n�vs^�,�KVˮ	M^�,���/k����6�a���0y�Cu�������N�j��ـ�k�����
'�+2���4�,#���L^]�)�VSq�n {-����e\^=^���u #�Wy�b(�jv�q����ut
�����������o?��T/��P��vV]Y�A>���m��L����LI9ݓ���L����)2.{���}����ػ�+�;/BꈅM��nf��k^�ZXu�_�*δ�k��!ve:���4B��n��6����Q��t��m��P;�z��yz:�����<�d׃0k8}��Μy?���ˋ#a�d����ٳ�X	4�!���ɐI�C���U��ēi�ZVنY���)�<��ԡ�f����۪���a|�4c]�$���9,��E�ʫ�žt2ϟ���o��᯲/�G��,/b!���P����U�O���R��s�y��������k�s��4�dc��{�|kօ6Y按�q� &���.7y�lDf,��c�����U�V��b�Խ��7G]N�$���ի�xs��z-�D��mE� �,����U�j��;bё��n��ݜ�g��}`n�w�POl �p����%���
�3K5�x�-)?���a�zI�^e�7�ϓ�mg����lvR���n=L�b;�|��7彷���������+n~���$*u������9$�7��'؎l�i�����i�(q<5��Δ�ZQ<&U82e;޽�&1/i���b�����%��0�AD	�����K��������Ⱥ������ь�nSz���m���C��y��j]�%?�k�D�2���ff�Wi�d����}�w���B��~m`�]�uךˤ��oW��4��v�� ��e�ǊR�}����<hr�i�|so&c��ofa�����;uV��Y�&�NtBI�-�h�#:Ǚ��pS�46<���E��k�__�#�>⑪�fN�z�SYY��q#�_+�S-s2$���dݣT�G�́{�ޕ�!,q˩{j7]��n�ÑƋl�?�Wk_f*כ�5�D����+�ժm�������Rf�q����7V�S�m��=�8�{�3�J�vG>q��w3�j�E�XcC�5�w�{�7�ҨX��T�Fj'�>���jT���4�EY����xߌN��z�w|���nڕ?\m'��2�k�^-ƪ���e1�n��|���[x���ű� 1r���T+F�cgi��X�U�������ѝ��:E�E�ɶ��7�Xۇe8��'}~�X6��\ͽ�Z5�M�3s�BvӴ{����5Я�$���%���};g���`>ҷ����L���3�,܈6�e ����nt�績�M����_�i�3�^��;���s���}v�
�a �;��;5�8���>�z�݇��ob5���E��r�'9h����A�v]S�c:�}�m���/^����j]13n��=�J�SK(�K�K_C��<)�cr{�޲k�Ů�Rgb��7���TW����
̱Y3�]������P��GZ�g�<�e��pu��&��;��.�1�Ύf�;���qy^2�z�UR���)�v��c��=o]7��ZV��4/ �a
k�z�z��U���a ��p̕*��ᢟc�<D�M�/�S�����j��L2��#jW���Wsܔ����&r=����;9�P}^[zN�$�>�9��њ\�<m�� �I�V:a�f�5]w��c}���.�	����n�y?<��w51 �\�� 3a�N��<���]�������e�jf��^[bsҳ��ls7S�皘���L����*��!/�����2$z�.oSj�7;)l���m�e o+B��G�T�֥C�A�MY3����_3��m���e��N�}yr�Gi�=0<�2�]X�����Lk���_,lO�a#��K��F�����ٕ>�l�YC(eϋ��c˄�3�A�mf���Sk����w)���F=�ݏ�=¼v�\���ԃQ�t�Ugp�K��C `��e+��ܐ��ç�Jǭ�7�y����ͼ�{��C�%�c����l���	`e;*�q��N����\Ӏss�+��'W6+�sAۢ��|�\��l���{�Em{�^a2Z{+��z��ٝ뫓1������q}-�#��'H�/L�L�QU��2ܚ��ۯ2P��n_���-I�4n�|s{��х]�}�=�1¦��U�t�*�އ�^��W�#ו8�c��;i� ę�i��4�ù[{���lGȼ8�Ǟ�?V�057}�)��z�����뢺b�x=�¤���"C��x!�8�j�ݭc�{lzm�%�T"�2���vAs0��S����.�8Ы�QA�w�i'G4&p�m�kK	��{+�f��d�g�����" a,>�A(N���1-.���7J]�G^����!��;)���{���8�U�3u�ݯ�T7�n���>'���:!(|�Vю3�L�C5�����q:��m��gI[z��Z�ԫK��") �I���B�`�������uG���'ֶ}R��Hlmžt	%PŻ�sDev6�wk��Fw�WD�Ϯ{��Z6��Z�F���ٱ�V=��y��ٚ��Q�2.����X�v�`u<��(�mn�k��܀��l�X7�+<ؔ���6H���4ҥ.ӻQ�ۊ�"�pf��l��؅��,��j�R��&,Kڴ4c^�Q�znn�x��>w*ٳY���][Y�;1D���&��}��+���|��7/c�E�@ ���}f ��(Ȯ��a�-#��ĕ-��݇�3�8=��q���o�dϻ��t8T���uz�m�bu4�sXΛ�d0�����Ab����8���eÜ�3G,#l�k�ܮ�5�Ϛ^��֜�9w/�pU��8�:����=cb:��H쾫��`׬���{�v_M���Y��s1��$V�1��i���5Ĵd��2�j��j��#�����a�`��=g��f[f˹:��]SG*S�:�k�#t�*��L���*�s����^�&q��.�8K6	�p��^ �=������7E\�L���^��n�>��S4`�j��0������_���_mN�!W�U�}/�S�:{��HW���#�����4���1/���yJ{3n<�[5
m��l�������Z�ʢ�Y���˃�|�~ΩJ�������mEj�yZ��Nݡ/[��������� �i�Q���75��Q�zw���vN�����#V>]��Ҳ��اy�j���5�=<�kz����y��-y��Oە�����X��-�������\��-$㪟a�f�2�{�Jz����1��ܱz��y^��M�R���ix�zjֻ+�j��br���Ƈ���R��
�'R�wf$��(�P����0�h���I(����>���D5�*���y��;�J��`��yN�j��T�j�-N��) ��q�a��FȽ�L��Xn�\�^+��[������]ʫ◇4R�#n��V���i����&�a`�͞B��s�i�;�^�\��%���Z�g{��K���D�7���淀�������ז�x��|]�U�o:ᮥ�4g$,�`K�2���>�����-Ȗ=�صfoN^t\�|�F���+k������@�ԙqp��+��X_ש����O{�Ļ�K`P�VҾ������������3P������{݂,-4Zh�XI4Zs��������#w���VX�3��]X�Z���i��su��;�Ri{�vy��;V���U"��u���4k��=*DtHx��\K@^>�U��$-����t�R(�$"�o��}L�����,կ��QʻCw0k���w	6�wi��=����+���LE����>�mn^�9����ܬ�I�'Asgq*~��ܦb��Y�@Ny������a��P~7w��	�F���f�,�c{E-[7	z=*�w��l�_�3<Y׃���ۺZ[�ݜp�޻� `��Vx���K�����	�ѕ]�J�[�]ɯ:y?�c^$P��B0����!�5����zi:x<�U3+��j/,d�Iܢ�.�k]�Ö��p]our�;y$.G�_l�������� 49��m���.2�Ӂ�·J�^��:�\���G��ܽ��-,���>�W1���h��Kbv��+S��G�#2��z9M����m��-����F�T~fp*��|��>n����c�+tޓ쎱O��/�w��o�v�ަ�j2��f�m�I����"#lBױ�4��f�N�ک}�~��{)�v�9�����0��deM��~ɞu9�gēޮ�4�⼑�z����h�w0���7�U-��7Md���u���.k��N�*�
�޾���N�`x۽hVˢ�w7��?n�w�k'��������u�k���P�oN��c9���~���<%��<�{���񀯿1b�����t�>?�n�	_��[�U��	��D�	ʝ��מ}������?������4PAW�����?�~��/�����D D���:: @���A������"��+L ���+B�! !
��(�XBa	�!V�XB%2$B %�P B�	PB$� BP���@ @H�N�E��@��!
���" @(0!* �����@��!@�� �J�!(@�����H�B��< �P BA@�	%D� BD@�E$T$D�P B@�	A$D�R%F%F F$G�������������������*u����	��
Ȍ!(���� u�B�B�!����B,!*0�*��H�!����XBaE�$VV�E�$V�XBEa	U��8��>A�/����  *(L(�$��w�������聟�����LG�����H��?��� ���ˮ��������~_�����?��A������@��`�P��@���e�����C�A_�?��ȿ���!��o�����O��A6;�WG���p��u�H(����H
Ҡ�H+H�@!HB�H�J�@�R@�J	@�@��,�)2B�"ĨЋ-(Ќ�@��- ��,@�(�
��"ģ$�H�
��0-�J0B-̋@ʉ) ���#"ҭ��,@��J1
�+�-
��,��
��- ��@��Ȓ0�	ċH��2�������"��J0H� ���,0,��"Ҍ,�"�*�*�"�,�,0,�4�(,J2��,"�(�	"ģ�īH�	ċ$�0,ȲģH
ʰ,,Ȳ@�ʰ,@�*ċ,��,H�(� R� @,B-(Ҭ��+@���2,J4���,��	"$@�*2H �"�@�!*2 �H�(�
�D�U9*�*-
�:��p��_�����"�( ( �����C����_�����ð�$�~��7�\����A���:����|;�'�?��#�@���������U��?�O^�t� "
��U�H&��C�p�P^�A��_B@D~����8���A|�8���<O���}{�`x������?��� PAW�R�������o���ϡ���$���@�@�<E~~��_���
�����P������.�p>���?����A���ߡ'���&�
��"��O�@��;�>A������?�{���A�����T��s�������?�q�O��(+$�k+������B �������E���/TRUIJ��TUT�E)UTAAU�!
�*�Q����B�*��%%*RJ*�%(�R	�������$Q�(�I���$��*"I UT�B�B =2�*$T�DT�A*PB%B�J�T��T<�IBT��EAH�H�(�E*�B� 	AT�D@�H�(EEB�	UU �TE$�J$�����r�H��  w5+aQkUZ���5��ILڋj����-�j�TҩhkLa�̔l��0�[K6�m�3f�Uj�BBf�i��&�QYb��J��a�J*��[�  ��(P�B�
h�E
 �B�:îΚ���R�&��EB��e[��P-b�kc4d��-i�ٍ�i*54�5+5�HU�fQQUPD�  �iZ�SRm�f�j15j��*�֒���6�D��IT*44��a�SHSEkZ�ت���*��*����  ���C�4i�-�m��FH���m�EV����
�$4dj4��B�T)i���А�U
U)"�*T	D.   Mv��dY�Ph+Y��1S-6��2M2�T5���j�Zhfkac[j�F����R����&�T��R��	()R��   #���@S+Mȟ�i��Sj�I��Z�TCUF �iXP A� b` f!�@1��UP�DE	IT'   g  ئ C`��k  �L
 h3S� � 
Y( b�  �` E$��J"R$EBJ�  �� .�@ �� M�i@ j�V hb�  S4`h �f���l4 kk  �
���B�*�  :@ �`�1� �f� ��� �`� b�Z� ư
��0 �)� 46��%%J��T���� j�E J� 4�1�  4l�� ��� P+h ���  f� )@Z �ia� ��P   S�	�T�E`4`	���a%%T@ h     �$�L@�FDd�M2&�Q��O&����~%**��&#&�0	�	��`5T�OJ�d<P  h i��J���P       j�m���U���9���[,�J9ML��HC �d4w�ye���>�ꪯ��\&���R�1UAy��ȍ��*�t���S�B*��Abu����c�?̟���}a� �5DT`��J���#D�.HF K�PE���n��R�?�]|��x���|�8КD�:C"a�떡ie�H"/��Ns��G����]ޥ��o	�&G���Kk4��:�Ad5[t�8^�
�9��dh6��X� �֙���d�4n�����cCj��EڶT�s,:0��qѽ@e^���ԔR��4�̫̬gwv_�E}�ql�Y-c3
�Wj%͖��E
v�5k�u)R�\aa�́hTv������V+�Aj��%<���34Qm�aSĲ:�m�2��J̀��	��ۮ%�KySX�]�i����SjG2D��f��Trl����V�bmՉ�nZ�в]�X�u�h[Dƕ�շ#*-�jR�tԱ�j�+���	=���+V�i��I�=ϐ��lK�2�(A��X��J�&�.�1B���ƈ�F� �N�g*� !�吶+"�-�wv���4�к�r܅5�+*CBOv�r�EtO�o��Z�՗��o2,�����WX�oo�V�r�Q�4h�e�s��9;�K�`�i�Vbj�dJ�ޓE�.��É�i҅�t�T�@�P(����7G췰�晸+Uk7-+pZ��	��ۥ���ʶ��41M5���Y��L-@�H�Lj:-�t�f���\��Bə@A+Ubܰ��bì̠��QըR�� �/,��ԡ����c3�,݁���ǔ��ѵ�[a�B����ě����f����r�L�vq��if��)Z�A���ګ��Ѵ�ZQ����B��3C���aS�T��l�xu^��q"�PލmV;� ���(�O-ϙK�E�H��6��%�M�8e��fm��Ͷ7,[��v��M�������FcUm�Z�CR��N�,,��&�:Tm��
ǌ�nJ���}�E��r��(hX�cW�ѵi#.�V(�Ԍkm���`���iJ���W���ܬi$�آ��:��A*
hQ��l-�BFT5�2�0�.ߘ��-�a������c"!��J-#iiY�o*�q��t.�i���8+����[cw>����YY��da
�XCwyׁ���)V�F��<�jx�f榅nˬd�U�i$����N$kn��jֶM;ܖ�̣�t�	fBP}fҔ��.:�ތ-�b��31�:��:�wN�k��j򔶩۽�Z�U�)5L�؝"��*�v��F3�I�I;���Vl�^]tD*�Cv���hb�Q�+˹�=H)��0��mi�DhdR�Uƴ�ԫ"�E/��3U!{`�X�z֋����C�k&�1@�(����h���Ōd��EF�����'3e�v2�CRIMږ���oh��
�f`#	d`Q=�6+�@"U�`���!)zn�LxYf%дj�cq��ufc� 5�{. uM�D�)�N��j��5yQQ�6��ۣzKV��;�n�+S*T�@5́X0�E.���M��FҒ����H�e���*���Q� H\�^�d��/6R��]c��Di�b՚�O"�-�oD��@���`�iˋZ�$�93�[�cr�i�E�����n�G�/a*��K�j�Q���&Y1�ǰ�bU㫕\�Yq��4F(35�r����r�9x�+I�Dڙ#�#"�a�Xݺ�B�*�� ��*ꞭȠ�ks(�K�F�ؘ�Z8�d��� ɹ�R71ctGa�n��IԗJ���"K�.�$�E�!��bP<�6�������,W*T�{��r�=Wor��b�[B�v��+�m�)KԀ��ֻ.\z.�.���d��f��襹��ժ�����kZde��Ð["��m$�47/m}li2*4�51 I��uu���)M�jA�Ck�6�E��U�fU)�ч2b"�l��ë e����Q�{j8kb8̲�fء�n�Z�+NHs�oqhw���ʹ��I� �����5c�@Xhٚm��ӗ&�S��&I[�kJ��Wx�Tb�<VLGs^,C��D��f1�E운<�u���)�����z�(��X]L\�w`:B�����ܧY� �����0������hT����2� <�ފ;X Юi@f���m�٢L��^��D�ˍ��qh�"�Y���h9Rf8c�ra4�ed"�6�b���@kui��ZL�N��(9X��杛M:��f�i�H"Hl���8��2^�:�j$���Z�f�(�Q%j�I� �k"��мFl�V���T-м[[PF\���0^(�e;�]^:e4�Kv����m��3y �D��� 831C��]*5���H���n���k,�ұʹ�m�:XՋ���I��.�I�����VPp1��4!Cc&t7A�[.�]��1f��a��פç_$2�\I���4��,�%9�1�#�%)QAr�U�������SB�͡��5n�+	�Э�u�C0��W����A�u�w=mS�z&����!Km�������]��E:�ɠ ;��mnn�M��X��[*�v)CW�m��v��w�Ԥ���ŗ��pێ�P<�Ů��t��fL	Ǚ�SkwuV�]��HQJ��2�[�7��n���wz�Â�b�kI m��]9z.*7O-]³���	���K@��ZIfeҌn�
@��8d6-��_��34�i�e��u��<�QƲ� f���:���ztl�iә�SgTݥ���,;-�Tma/eGW^�[�����T��ŗR[ZL,�YMm� ��]D��	�X���A�M�B�*Ûp��F�j�`�V�܄<p|٢����{R�J+	T�@a��a:��u���:[�
��zF��R[��3r�y1$ckD�m����b�^�����V�R=�0�*���H���VA�콈b�^eԊ�+% ��ѩ#xX��@VYd�tԫ]쎥n�`1J�B���i�16n;&b�I����T.HM��jb8��5�a�%�n���N��ސ������+f��7��������n�7tK�`9�7`��B���N�*�*�^��B�x���bQ2X�F�|�G��2d��SoA����i:uc�6����H�f�b �呱^E���F7Z�imh�]���f��Lm���{(cّ�[�L�u:y�;?LںLh9i:��(�;:�b�*�:.ޤ��H\�^ɸ"�Q�L
i��isZʖ�#0 ����K]�Z�Vݩ�im(���1�������e�\GKĶ�!ͬ
��Sq����;r� J�lKW%�1��#�V��b�n�];���Ʈ�P��K�n�Z����y,��@2i�-�{��+�QV�� �ԭR�i���oiT-k�Q���w`�u��)�-C�T�R��!b��J��Q5����ɧ���R�+3�[��*H��,ҩl�$���N��7sL2d�a��#-Il�a#%�����%�Kv���W"�`����$�յ�#��I�/in5iX�MU���%���.��zCǂ���CpLWA�"�|>Kԭ�o[�&�jt�/E1�.kbn�ZK�0�ݔ���[ �VC)���̭7{�L����l��tS�B�u0�����(51-e�f�t�5�zM�m���L[L�(l�C�#�*�=Ĵ�u{3Y�Y��I��\�q��v����h�b��jQ�RQ	7j�SH	�(Եdՙsp��HR�(t�Ըm�W4L�1��Yx�u2�2�M�wvi+�r�nQ�sh
��j����.���	RTY����ث��3�,��d[tʨ�¯lY�nK�ޑ!�g;L:z��[A���Y�I�k1S��E[N�J��^��AJM� �f�ê$�;7�t��+N�b�]�!����ҋ򠼕JNQ�<:���ϴT��ʌi:,�r�gl��бJ�:˼�j�>�E���,��\B�a����kd
�QTR��kib"�)7����2��t1^�b�#Ai�1#`h���Շ,ۻm��jڶ�B�L0GPWF�E�%^'5n��Pڴ�0�Ou��ڬEf��a���dh�Z6=\٠-�#��*\�ըf��:�ڔ�h�؏]� E���2P:T��1��54����x�k5�x�*�n2� ��W{�ubRu��nf��t����(e�`�K�1���ZK��!��t��@ �d�fҀ�g�̀R��Qe��CD�5dٻ!6a)1yӯu�l�YR�Ε���KD�hc�%kDӄ-�n�TiL����77>�m ��E�.\�oE�ڷ6��I�5YGl���V�����0��a�m㥨��V��q�;�/N޲w
�e��ܫb�ù��A&5�(@ޙZ�3��U��e���"�7��QQOi=XP�+)Q��e��ˈ,ȳZ�~���~&�j��^b?Dt���XwD
̓ER�]�K�#6��3�+>ܺ�a{�-t�#5��P��Ą����ҽ�sn�ˉ��.U�浌eYO��G-2u�Mԅ�B3��5l,�oR�h�U������[��S)Y2��ne-��܌;��P7�h�[[A�Qi1T�6�Pk&-�۬�#���Ӥ�T
�>E�ѤM�M쭗5�a�?�ᬲ7R*t�*���h�(kx��[�Y%E ;�B�G �������I�=�,�#��)l�l
��@)�mӱ���.%r�b(EG+H�0�b�]e=50��X�p�j�����DU��f��U�
n(��&VK�f�۠��HPL���I�lf�o]u��fS)S@�����y�k�r��fm��jl��'�h��.8v�&䢈�sPt%c7��A@ì�c��H��0����V�,�a�4]e��U�}�j #7-�!7Pf<9ͺ�uP|�r�Qe����d�6k76=CSU�xе�k
ޜ��h���fPR���IU�^k��W��!����n��aaD,�w�p���!Y(ҽ�j�xv��ud$�q����W1H��X��lᅁ����!6��R�@��7�V�/v��$�(�TϷ]�b]c!u���V$�ٷ^0�4�3-Z���D//�\ cGp�ǿi���P���Z�(��{i��;��3p��j�,j��6��<H5�����%�D��]�8�FU�1S�)�Kt��.���@�]FRa\ �u���V�3D	�����D���Vѱ�C��K�Nh̋Rby�Z^�xà��G���Aj�h��ֳk6Y�Z��ŷ�������H���(ڱ��S;�.�]��flA+q�	� Z�o5滣@�QXw[���L��^4�2��%��)��6n��ݼ@�TS�m8���V�n�i`ɟ.ć�t2��jW�2)��V�2��(�e�Ц]n�L��f���-�Ek{K~�Dh������n+!�l�en#��佭V5�o�4�܊CREIܻE�P��J�!�r]�� ]��-�%��O�Si������Hg*%���V�FL�j"�Lҥ`�䬴*dr,���j�(�Rd��Q@�*�R3v��C!}��i檺0��Nn��4U�,P� �[6흔�R����VÊA=gj]Y��%��ei��L�t)����0��꠫5Q���`�!A�V֩��iH ���͓sshM}���M:���Ql���欀P��h��z�U�"��<��N1�Sn�-`V�M�:���KO�l�S���[M�7RbbA&^���ڱ6��
��� �fS�>g6b��v9�Q���7@ sMv��b�[y2�� АFT�\��{W�/Y�4N���J�r�%ͬ�J^Yj��ZcTU�'Y��n3�F�M�o,�ˠ�[���keI�؃t�H����6JpX�Sţa�l(f���R��El��D��vMk���cbW��f�g �Ԟ�xi��e%D���J�X�h`ņ	T�*�^��A�Y��L�Ib�e�ui!z��ݭ�W{i���Q�%MӅ
���E��l���$�V��t2M�q��oQq�õb��(-��1�4���6X�溳�]�u����n��_"nd1i��
RY�oV �A;M%�����2���L�r�oM�����ލ���K���lW5� ��wyű�'�N���i�Ie �G���z�k5�:@�&��jM������j��&���%�C/��&`��3�U��h�H�Ƈ��A2޻�e6@ @��z�E�u��o���Oev W���ϭ�<T�n���r]�ote��{�Z)������B��J��]�S��Ju$sM[۶E�e��T�j��:͗�[�%knm�mee!�Ga�B�V�ɔD�P����b!l)�i����F#��6Ց�����7j��m
��c䶯뗇1"���#�r-�$�r�T�y��(�lh1*�wt��>�e
с��e=�U�vwDX1V��Q��3S���ڑ:фm@7oK��V�v�9V�E��R�m�iRB�zR�hR9��1�v� �*����IN�Xߍ���F0q�4�V-�[�2���B�[� `�*zkme����2A���f&�+7a"�����Ǵ:r��O" ���1�".�. ��݋��0�2ҁL��^$�s�*�L�mN�֬29/4�Uεpf��-0՜=�h��U�Յh?Ct�W��(��m�Bƪb��Ѹx��V̜�n���8���8$�
%A�s�M��c���hm��/0�5���yy+����X�ӈM*{>M���k7��v�(�ɔM��V�]���$��w��A�gK5sK���gU�L�}˵��"V�~�2�u�:J��,�/��:�o>4�}���E^�85��`�99͓�u�{S��ҋ]H=sR���Kxy�D���`�AԽ]�W��j �4��-ֹ-u��j�r��5�u5w-���;]���v�ĺ��z�t[��\J� ��'֛_#��{΅�n�n�h�����ө%9�p]����Pr락����ɏ���Y��:�k���P��s���̓i㘗f\��8���:,��=�u��H��e�tDN��+��8(�v�r�o�*vi����K'#3�u�ur�Z�>@����Z+����x�4�s�0m{\�qޮ�fP]��왩5�:��A�<x�m�;Q͹@v,zlt� _bs/vuǶ�c7WRUf ݡ�c���z��Y��'�6ݍe,=qs�`F���v���ܾ�j3�ô��:��%Rr�aˮ5�����n��;l��@SƮ�1p���9�V.䢝�Z�>;*��X:]u�!���z����`̡o�
��2��x���紶�v�@��bnܦ��B�kj�ۮ�ł�YV���f��T�d��ڵpS��n�&i�wè�����V���9�M��́�u{+�e'���7l3���g��$$�;[1gҒ⍚�%��%[��yX��	�0��=���\��B=�7���YI�gvv�6�� �=EP��_T�&�'n�m�y�F;x�	��wQ���f�n�L$�Wː֮ěݺ��-l��=���DoCF�*zp1e<E)]������m�)�'H�73P���',�w;yR��	f��̴���F8�P���p�OJ�z��y�[W�	9�v�;L��R�.)[[}N�$�sj6!����VC5o$P.��T:ID��asf�Э��1�Q���vR�Ւy�z�m��4��'F�i9|bo�"��7��k�M��5�^�S�..�F�nr���;Z�J�['�])�X�W%��.�`�� _#�����p&�u�*�y�>�F��z�y��8̶��wY�Q$EFI�����3/�g���V�:�T�lwW��������������E^��Ë�CNu�y(�����=� s2��k��Mս�q��6l|^,4n��V�i�Z��r�R�*��ķ�ְ�8۠��3�����fU��=j�c!t<�|�&nvv�+n��sY�+��K6���N�_]���#��΃�Ah��2�
��7ʳ���4�sk���g[2k�+�Nݹ%���&Z����(�*��N���ޤ$���X�uh5��ٻ3h
k�7Y�o�hz���u�_,�:f�:\�;�n�T��Ŭ���e,�³��Y�s��`���[ۙ���7�J4�
ӹf��)0�/�C!�5������cZ��+l�#�F�R��ɻu�wf��e�+F�|Rش�\� ������;st����Fٰ(j��tM��:��1�q�'M�\u*^]�󜁈�&wn`ct���R�۩s�6�2Vu	{�Ӵ��NMmD�\egv���*�Bh����v��i/�M�'�u�o�k�}G�ܦ2�+��Ω;i�1�[�N0�-���6�R?e�����'05؉���j��n�����8���-=e�Q\3���|���u���$LF {{��<��5u��9��>�\�KB,��@�qIͥft��.�u�Z�U���0���z(F�%V���j�/�A�]Wn�:��B�qZ�P,.�w=�j�wɕy��������:z�����.8����V�=.�i�gX�<�+:W�	�������L�9��Gu�lA��(���N�/-on
k�
��k�e�Ѥ+w��K�IZ9:�����hac!L֊
��	㕴��F(���nP�Վ�Q3x�q+{ίQQJ��7YΗIm�ͽ�El�%J;�����֞��d���
�����^P�:���	�هo��t�t�:r��L�j��-*L�k���]1��n�p�lv.nwAK��y;���bW�9����s*��or��	��w}:���4��M��9�Z* .9�_eou�v���j��ŋ�����A�]���m@���Q�%�O�,2V[�T�Z�A4i ��4c�\7��Gs���|;�j�R�:�k�BX�c��"�B������6�-�\E�u3���ܨW:%iq�VM3⸾��FY��+��r�e�W@\l�&�PT�%�)$#�M�egKme��L���CrX2:�Hj����~m����ky_i�ҩ����M|s���׵��#���1@�Uo8���RkC�
����óy7v���\�-h<־?j4�u�qU��/���/�]7;�`��fRk�igO;�o����	��;�z���c���ЧXK8��:�"�Z���UokC2������Ɏҽ���KfR���W�U�6*��+V��VJ�Xz`Q�tgE�{k'a����Y���j�
ó��Ja�}���YGr(u�5cv]�t��#����W\룙n�2����]'r�̢qaaM�֭�M��}�X�o��>3n�3Ɵp|�JAT�gFF���v�Y������Ǔ;2�m�6:`-%=@��t{b�}�T��iܧ�����K�䚦Kw5K�Q�x�u��1�X����OL�N[֋[�\�����Q�9p�;h�lp�M8�2�=Pm��w�6�v�\�[wg�7�̛}j�ԹWZ�J�D��tSpF�-L�������b�WG����)f�|ᓻ����o��ZWU�55�2o>��X���
�y[�ŷ��������X3�T�n@�i��,N��ܱ�Q�
YA)�k`�ȷj�1XA�*��C�k:*)�#�k)" =]3�R�ur��d�V躀�n��փ�����J�µS�6���I�@e�Y�Q��CQS "�Su��%�c�����@��
F%+5.�Lc��SEbUr��])���C��/n���L�gY9���0�o��+9Ļ76���@��㡔F�-��l�B�Δ��8��ΰ�w�J�F20��Xe���,ȆZ���2im�m�5�{t�F�䬚U@ܭg{����S�rI��0E4%ޑ\T�G�$&el�ww�W-;[�y�F%����-;q����b5P~��U�(��dn��E�,���S5�F��IQn���:��ԕ�����m.��;l؞�ɖ�먖w�V���Mn�:\�ԙ����ԅT�)��7�j��yA�շ\�;�+�к7MZ�h�׋�@_�
9OFQ���\��:!iճ(X����hl�{_Cm-f7,�To^�*N�ʽkiΐ�Ɛغ�82sum`����U�u��d9��t��a���;��,]����3�)��9C��V�{LGa�
��V���N�	6=#~	�u���ol��u`Z�!C�੼���q�vmI��8_',�jcK�T�7���������V� ���Ϝ�}7�����=�[�l<z�3��C�&�K�LS4�u�.sJfI'�(��j����죸{�����y+�kU�1���V��wg�,.���X�6�<b�6�D�]��q*3j,2Ħ;X�έA6�ص�w܇	���q��bհ�]�BX�uͧz;8����G��M>�gS�Y[`�Z����Z�sv,]Ju���]a�]H��z���}����!J�}4�=��)v�*����՛��85ʱ֝�E�����sy�{,bhxoE��z�@gB��<�e�C���zحMn,�i��5��ƣ�u-zXD����q'Æ��f���u��܋��kju��ѽ��ν�*�$,�3N���ys\��|;Ugo6��c5��nl��[����Go�񭢉���$졮��Y�­��h�hh�r��Ce,�v�]��2��oP�����L9\H������;�DΫ��_a',���4�Q�����t�Ai�������,�mn�$m�9�D��(i�X�	U��Q���rTml�qj� ԝ����b�˯kx����3��c�Y���Tm�Ηl�E%�T��פ՛��Ki�qw,�-b��[1b��mRnՒ�fk�Z�VXe)�[O����!^�v�]��;�_<�eZ��D�;ݕn0-��pGKd�>��.�YNoU��#q��šc���#��ƅG�v39Ԉ׹�m��з�L��(�t������z4#}��b�����3�7�M$3Hb��w������!iGds� �0u��q3�ʥ�#"�x�\�a�e���n�CֈbËue�1b��c���&E4�Ф{�>�"�
���A��\�uy�=����)��_8u4�_���˴�����n؝ơ�"q[�����Xi�1a��+ �"+���Yݚ��2�E����e��납1�����k��k^+�d�
��l��q�O $����@�#�L��F_f��I���r;�hgGu�՜��쮩K�{:e��jF�P�0,����)r�C�zE@ʂ8r��ʴ-����g��{�h�n�V�Gb�:1Dv���o�=��]'t2��ɰS{��f]����d�m��`�]3Jvo#	}�K���1M`�&��\�����n�\�V�����m'�ГH��Y2�h�t�\�j�NԺ��t�o�m��
�jU���Uy��Dڊ��0>X��|q�v��ײ�lP¯J�Oxq����Qe��<�_q�Q*H�b�ᱶz<�y�[m�{H"��]��D��Iͽ�e:E��̎��%��{#���i���ܥKT���\8�xs�s9��o��t��
[�3͝RK�b�<���br��6'7�;]��静}ΤO���w\�:a��Qw�Y;�b�1t���WdI]"�.�'5-u�B�7;pA�[͊J�a�]�����K]�u��G~�<Ec��W����]Y��YWWi�ؐ����b�C�]
u}����f*H��jc;FG�sys�t��یV�������J`��l��ۚtV6�q{�x�-k���s�.�b]mf�D�8��Y�Q�#��&D���ѓ����i	�+�o�N^<MW_J���x�0�ޫ���ce.�U��7p�����em�nR����Y��VsS,�܁���$3����"¡[*�]cW���)+�s��qbT�xj�V��U`QV�pR�W����b��6s����6��}�\љb���O�lr��:u�5ڞj��,'Vf�)2��q�O)�ZU�����@� r���^6�����f({,!�'��UɌ:�FqN��rI���n��\dm�ػ����v��N�X�^j�ì�[kWp�J�ء�酸�]m+���iF�ȝ<��8�A�Gb�,�t;
�ރ�ݶE@��,
�|�d9�_p.��j��I�k��ʅg<@ڙ/�0T]��uG�b�ɄNX�q���5����e�unifh��Z��/2p2i�j��)5��!�wF2�ix�U��,�w��I�	8�LN'v����(�ύ�|wsh�@H+"��,�S��KpLU׶ĩ�mYn��x��@Q�����ޞ�S����w>���t�D��١\��Ms��e���rV��4�c�&�]N�v�f,�Q<��W�]�C죩�,GW[��:�U�X����ݠ����T�537�R}b�1���RL�
B��Qa1���UVl��'�:u���k�V��`"�B�k���5��u�-��VQN�v��e&�$.5��sI���[�R��-W��J��䏾��ջ@���O�� 2̫C�q����~�Z:"̷Z����aBh�\,�o�n�=������ӥj���z2˩�%5�X�-,��Cf�fb�g�]�ۊ� ����t����7U-�ΎwgHgn��ٌk{\�6����uj�8��F.�mNK�<1�fۆ��H
f>��'�E����G�a�r�0�X\�0�Em�v*W��];E[̩E�uoI��t��r��5U��r]C�_u>�jn�ʱNy&�uauw�`�r���|���N�����v����x�l.�j�Z{��o��4�[���p��*T,l᤻�;��{���G���%Q�CT����v()a����#�xiE���w �ıu3����+���L���R�/6N��.���ƄS	vs��eM���F��ĳ#/۬�o����y!���*K�����KM�'m�ldނ����/��AF��ʵdIܳhR��=�lvi��e6��㸠쳢j&}�����Pt�eĬT�y�og2���OA����O��W�������{���7K�rT�Ĝ����@;��c�;�W6�l�N�2�$�wS�J|gJ]u�wU�ٕ�7�"jT/��j�;�}Y�_��-��q�Ӧ�|:�S���Nz���:P��"*�.��V�UE�բ u%�i� U^�����^��i2_�����^D���w!���Ľ�И��;2mꮨ���8�&ul�|�Y]u�_#o1�@:�	�����S���`Hqt�q�������v��Z���]���].�����Lʃm�V_r�p�w��}ض�i
а���`����uԫ����]��$�����4Wk�~�р�$���μ�_W5�L�P�B�b���%��ߠ�\��͎�2��7Cw�am�-Z�w�87l���.� ۣ)�|��r�)�[ 7)qcS�j�u��dA�n�L�.�Ǘ�$�,w="�� ��L�6�>�Ph��v*���4n�uE���Dq۳:u��7э�[���)�;�v�<����5:�VԢ�vIk$*�A����#}3v.\cf\��pc�]&�b}%u�����+Y�}\7��1�u
ߩWu:2�X>w���ڃ���{b��d���2^]N�ٙ)^΄ �*E�3w���Ȏ;�������z��!�a�pO�iEE6��s�KV�_v����暛n�t��]m�K;^�)�ݚ�¾5�&�yX�e�$HM��Ԯ���aCr�*M�!���J�7O��X�&U��j����z���|��u�cv�1�+3�rS�E��}�I����ˆ�[��>i49�3h�3h�[��,�"s��&��;E�2��+�~<�n�f����&�>[[�?��ہ���+��,�V]�u���9�NlP��;fp�͉�$�Uؠ��)e�9W{ԭ��>h!뀼��O�����y,l+��p������X�tm����ˏWU��VS�X��p�f���@��:qk�<�]�
R�WM4�+5eO��H�i�[Pq���q=ɉ:�/�e�l��S����L6�b���P�P�o`P��rӹ�ܔx3�^��zU^��6����#<����}����fx�����XMޙ��m>���H���6��nm�lȦKf�i|Miyg�À[�
�#t��30��n�v�q%�`���[-�h�YR˝�1I�����],����ːԐż��2A��!j�h�#~=���F�a�s�F�$B����}��:��H�m���U�w������C��Ҽ+&S���e��ݵ�ѽ��2PY�������5��k^mk�{N$�"���d\�s��uWA��ILM�VC�5�C�yڭ�.i�GC�ׁ1i��5�o&�&��ܫ�ꐢ-���{�-c�����a�9�b�x�o1:�Lǃp���@��v�#��P� �K����|&�D�����,�����B�['�T����J��G6M�5�s�^*�b�����Mq5:���7���O��L����o��\Th���W$��R�M}��@Q\�"$�VKo�^�ɍ"�������{�Z�U*H5�{�*c(���dS�yT�2�.�VT�`1Z]����u3�6]�p�96�a�z��lo_T���v�#���׮�fJ;$�k��'.$٨v@�n�U�ۮ�mq�ڒ���b|�,���əz�$4�]طB��]�a���o��o5%�����9�"%��V�c��.eJ����p�W��Ɔ�vj�;eo[ߟmQ�;]_B�ιR#dҤ|Y�$ ���	(��� �lի�rY�o�I�n�D=� c���-J��+vT2�V�&�LǕz�U�]
�Z�jb���iʽ(�®�/%���:���ϵr��"�r<�}\f벛Oyt���u)ꥹ|��o7o>�mɿi�t��[Q��(K8���������kG8�)�	�n>�Vͦ-v+C���/24���.J]g��%_X�-o�~HFЊs����e[��)V�����dE[{#�[yq��6$]��peW^��1_Z��|�dm�ٛhs��T��;�v|���|X%aU{NQk��G�v㐕/F�A���u�ruZ;�1A���1n
���glt��z�9���u�_D�5�]�꾺��Z�wo�;Tq��@�J��5�V�mM�<��>K\x�ʹ�\�/kq�L{u�c��L
\�R���j��mKJ��5/�>��+~9��Ł,yX&�l|OL�־=֞=��QLc�=Vz�Mfq&���D	f��i�5�q�7�3(�X5�h�]X����>8����W@^=OjX�F�:()uط,on��n�R���q6�T'$%�+v��Ƨ,�,eQ�ay�/���ɡhck��Z⣬��/n�Ok��ا�f�%ݢ���1ޡ=XjŻ���H�楪󒧨a�u�#�a�2�Ans���#vT�9����n�c&+��b>��o���]\�z;Xa��b�N�t�	��.e� ��w ��]@.r������/��) \��7+8LiGm���]��VN쵲�u�f1��[ai�+Ӡ�Z��j��7Թ.�MW�>��ڙ7nΝ�Im��b�v�G@��u}�J�B�$���P�ԓ�CNF���uh��e4P\������)�S8V2v^<�0l���V�t�K��f��p1�s�0;�u���u�p�y&U�|�]��m�#��v�Zw�B�wq-ja�P˟G�8၌.�88��&ͩ�Na���4D�Qt�rj�vԗtc�\��]��nV%/��K�E-&vo��r[	et=���w{8�B�RN�g�>�/;�ը�]�6�h�䰵�1J�cl�R�!A%=�xִ�M;Xu�x�������bC�ա/;���'v��W��wMu���hkOr䠎�Ƶ���)ڋ�X��r��>��1�����6��H\`�T;�+w�)�X��;˾j�%�0�k����7Aw8�4p"X�+-�v�dmI�����-64��1d�Q���R�v��1��`$v�[�͏�-�iE�b�6�ovofV�`�Ro�d[��{j�V�n�pȏ�݈ي�����*ᨙ��\n����[r�z&X�6f�R|d�}�#�K����^=nI�l	��h�{�iD=�4�\Zf��]�����9�:h�j��;�!�p\ˊ�K���X�1��9�xowe�m
N���uo��"*��=���[:����U��tS�����q�;5����T嗢���K��Lh�!k�7W�^F�uu*t���0ݰ��E�9'�ݢ�ݝ�ÛæM��rbu��z���Q�Ì�
�6�o�_cX0c ��6]c�z�U�N�&�Ю��&E�IΘ1v�oVW]�,��}V�H��h�F��N����.h;��ʟi���Ө��O�|�QX�5Ks.�����W.��)�1M�{"��z��ɸ���%&�7DfV��:���U�7��r�/�l��XɆ�H��Sm�)���u[An��,�#9���(ϵ-U�f�C��H;��Yb�׼-b�4]����>�&��{��8�Ͷ��oս���u�6�|�Սx(���m���Ã����Ǿ5tx���3*��"�|k�Q�V:�m�\�H��˦vs����u(֚X��YB�v�yi�ݴ��/�U4�x5)���t���c��$s���N���r��i�����sf��Ys쾔�3�n�����k������1����mCa��|�:���^7٧!�{{Wkh*UA�|�b(�"��N��������l
��P�f�e
,��K��2�xC�1e�2���${̗��}m�ӊ�����8[��K!Zt��\�:�]Hs�s�q�j:�U�(�b���ۓ%�ծb8,�ā��o0����⑮U�=y4/����β��K�����[��b�n�}�9�sՅ�T��e���@=��+��<��Tc��V�ݫ���6&�a�C��Pc�qvG;;����9�$t<;�Z;@s���s0��#S�®�me�V�I��c�Q���{Cs{���#�%nr��jN���w�V��'GBuP)9�ՋMnY����\'T�:5\���A[S2�(��L�i����K۳K���9�%�>�ܨ�tk�Ӯ��z��b�ACz��4 �}ұ�.^먮�gkK]ƍ��u��ޥ��<����/:�o.�$;{3N�ԅ3k�
Dك �:�*|Ŵ /��WWWZX�(�D�2|��N���)��=�l2N6#zՑθ:����؎�e�d
龩�J��sogR�ĠJZΑ�"�K��ݜTz+DИ/Wc�`���4� ��kͮ��Oz��I��:�� uqb�u�(,��/	8��8�c�űbh9����c؞(�t'|�5�Lڮ�j^�Ǆ�LfZ������#��wS��M�E]��L&�g�Mvh���]N�b]j�����>�ٗ��Â>{cdmw�� �P']�t,�����R[QJ�1�ެ�r�3��l��+|�]���f�`�f��N��^�v�u���tż̬"��B��F���t������`�w�]}",�:����E��n[� g*gQ�ȽR����-"��e�&M ,m�n�$<�ty�ַ_�YU׼8G�rK����6��7�MZ���9�3[�'zG2����٢*j�޸����e覊j�LHs���ƥ�.D����B�S&(�I�N'}��xyt؟6;1ŻWZ24=�;����އ����H^,��YI�ކ�t�k%+�MN���ǩL����aP��&v]\Ҿ����R%�k�BҧT�����)�5��}�g�Ѝ��M�0U�U���	��Sv!V�r�.�[��$mĔ�X���mS�/z;�}K��p�Q�����>�K��s���rM�蘩�m����\1�/�>�pC\JJ�2���N����7�W}��=E�"�vv;WI��(]�F?���Y�>q*=#�"�T*�����5���rl<J���s��+WJ\ӎ]��r�$��׷Q�E��aV�:|�Ӈ�
b0�-	5,�X����<���w}��{ZFuVh�d�ޛ0���q����)�����RG;WV��P���� ��ˤ�h:y\Yف-c&�Wrz�rv0پ�h�VU�����M�L����{�9;ӻu2���Bɒ����{qhᾭ�g��E��K��`�d0Ƅ3FQy�R��sz�d�R�ڻ���P�@�(�$����0}��+ �vHv����g �hMT��[��u>j7�5A3 "	���+�U#`�S�7���u��l�Gη�Zâ��K�S��淬
�fn�jl]�|h�s���MrZ�R�����3cP[��VYESΫ�:m�����-�o����ۻ�� S��J���6��c�E[��]0uP�l��&�a�������t���P�D�d�+�Nw�ۗ\l�k�3 Y�f��e)@8^�Kї��PA�-��b���U75ٕ��ǯ1N�2k�x�6��w���7N�5j�󭜛�V)N� ��Q
�Q	u�q�@�qsΊ�㜳w;��m�' �Rc�w�Z�t��0��T끬p�Z�\��8��RWE��\	L�׶{��u��EiS�lHﱫ���9�g ��̎��J
�l5eو+s�;&pm>.�`�",5�o�53���ӉmYi�U;�wA�z��epC�Jѝ��-[��n�5cW�?�-<�K�q>�IT�e�b�"kZ������Wb�ާv��\zX��5j��yW�$�ꔍd��$h���c�Wb��d�C{S)�����O�e�d[����B��\c���\p]"xj�ʴfAPiN�cC�>_jtk���AV]�z���bBJ즩�Mv� Ӊ�ˡ�R��W���#�,�6!���k�����]�}һ��b��Z���SI6=�]�2�,��,m��;���Di꽠�ۮ��JX\���؝<�����/mI6��`��ә�ә�1�	����n��b��R�oT"�^-����z�{��J�@��5��ԖZLR�OI�^�###��7��{-}�`��%���]xr�"�of�j�T�}PP�ֻ���9e:�wJ�S��5^�W�w��LԘ\�}���C���r��[�A�h��sef	�Hx�m\_s��e�˘2�̔�I�f>���N9t�BTM�a�Fղ!�Wکl.�����*���i�hu�OuI�u��[����M��λ��}0uEx�����goJ���.5��mw]k�"��G��])W�I,Z�L��oo��Ij�=�bxY�����f^r���r�Ad��V�@�e���`��%��]e�Of*��8�b3�G�ynř cn�U�ݸ�t��Ǣ�q�Q���t-a:ؾ�g�ʔq�;oKz�c�b�݀���н����e�Q�.5P���r�P]���r�#]C�bQ���+��.B��:����=�OK��$b���{���Ԙ�8�5L��J���t�����լՍ=ns�ud�۬>���wg���j}+9eu��hG�R��� �����2�i�[v1����h�s:I�64%��n�sY����B�g^�ʷ��M�:٨�1�tz�&֮���:�X"#؆jP>����>��k���flO�I�7{�dU�k�B�3���h*|�g�����vv ]�+s�5�K�~H0�:��,��c,��a�q�K[Rf*�[�:�\� 5���',V����(���c�b]��1�M:���B�f�Xy�ʙ�*��ej�VP�M	���ZR\\��.���a�ٝ�M,e��v��o)9٠�������R�y�i1>������:�V�ׂge��gI|����K!:gY�z*]'����%*r�{Mc��۠�Hh҃��^�}��Hj��Ŕ�����i<��Vs1�׏����`*�,VN�x����:���dTSs{�&J:��]�,E,ɼ�]����o�#6�mN�i���xp6A�71c�(�ge���A�`���y;I�Q���tpg/��Uʢo����:S�������T��P�8Q+\�^%�U��x�3j�%��(�\��=a;ݼU1%���*J�܍N��{���8��i`�Ô�h�Ι������S��츖��m$9M"jj��4�6���1w.]�n�v�gF>�OF��N5}0,d�FXN���Nr�%I�nۼ������kѻ�t$ެx�͙}(�埢��.H��]�����}��x���˻ʾ�j�I�h�z�.z�3L*�8D%{��a��:H��+ҍ*��/G;�S�A�T^��q�/E�q�DG�D�D�G*�����K �S�NFq�r7B�C��E��3�Q�xcWػ�tw3n�x�B=@�[�����"�d�+�9*ww*�#�r�T5*tkr4�E'u-Ԃ#�V�9)�;��U��	0�+������,X������]�B���N�r��ӹ�����Ls
�wq�]\�\��.NAy�=Nr'[RO"��Un�K��V�Y�R<�R�Z�^d�J"w<4p�,�e
��%$���]�'q%#u�hE\�:k��rѹ�s���w=w\Y��r���<�R��f���.`U��!8���<�IF���������t�
"�H��2y�EC������C�����]Rܾ6���wZ*QS�ؽ�H��_}G�%�pb��f���oG�L˾�*�[�؟Q5�$��EM����tp�3)~�v3K�g���f�%���=��tP���}�9uOr;E�i�>�1z@���z�qY�7Sϴ[������N\�h��ԴUFT�~uA׻'ޖ�
v�aHi��}c�@4�'n}��2u�a��`�_{�銸~�
kD"cK�\�����gr��	/���������W��AN� �����F�Z�ԇ5�v"���Bc�%����ƚ�]�*]�{ۺ����a���
˾^p�����	[΀������L;�4���c�c��ݚ2��:H`�c���`��oa�P���y�[�x�>��b�衵�|�o�c~���//�!�mO-5ۮؘ�෵V�|��vz��C������H�(C�G0�[j�R-v{k,{�~Lw�[��7��}j�VlC�e���5Ɩci����<��ա_pY�g��V��o<=9!�׆}Z^�]·�����|(�R��#����d�Tg�����6�,ȨR����3h�M��7�q�Q�9N�ut�S��br��[F˫��J�
��>]�R������{6ʡ��q!Ԋ,�8p��7��gh�S%������{������sÝ`��F*��ש�=M>��o�ݙ]p�Ͻ���{�a����W�f��^e�[�i>��1.��:��}�Of��J, ��qR׸Ӆ���ʽ]�/�����1����s��ͺ8b��[�4~�!��w͡�z��ʴQV��:����O���>x-_-Ƹ�;����:��N�
Āo�*zRf>�������T|Nn�_Z�����i0����\~��P2|?��e�l�͢0Et�,j:��r<:����eeRϷ��69��!<j�h+*g�^�*�Pě[�Q�M����D�T@��@v�����@#�A����2ӨKx�=�d���<Azĵ��0�#�QD���Jp|�e4@;<2	B6�U��P��ӯq�拃�����k��ؠ�]�N��[����:q�17�?7���(KtƽL�,w?zwX#���zE6������G�40�(��4�[ic�TQo������|����x/=;D�z���o��ɊgY�N� ��������@��^�u�zC��,���ϓ�3���Av�̅n�p3Vd6bl��k(�E�Ϟ���;=�49��M��� �����_]�)Q�e��x��ls㐾˂�b�js�]����v�*�`�;ϲ��a
̍j�\�[z�JcV(��g0�7��7��"�ʠ�p�}��1v2.y���ǯK�X�Q���N��텍~�=c=�b�<7�
џz��CV7�#,�.�c���#��*��/�j��#X�u�ju��0������@_b�i
��Kw?O��W�}�,F2]*=�E�RD����W����[u׷�t>�Kt��!X��~:��Ŭ�W;��><�+��Ng�BSpZ�t�
Vp5��,��-*�q.�pw��U-n�[�����I֯���z��v�x9V���>R�yUvMJ
�F��u.Uk;P̧dL�jk���wR�+��"D�(�ϑg`@�^-04��Z�3��Moy)V�������;�*�+��s%ƣKKgDc6�����kE�V莂�ƅ�y�ئyAN�V�Ў��������l1�I��^�}�}u��#џ���	����thׂ0,�[�v��7���s�n>�y>����5uÕv<'����T���S�(���&����X5���^;(S:=��ZݞÝ�Y�;�}�me�Hנ0M��+I]�U>�Y�c��������*�f"r��K�s�)�
ձb�9�oy���v,ds����vm+����Ӱ�Ƥ׋U�L��>�M������R��ޅ��Q�
�U����� �Q���7h���ș�o�U�;C�2�Qj��Ɂ�E��xW������
A}�@o�5�lfR�H��9O[*�A��Y6 Q��"5�x%��D�ro}�X�t���^%��&���}��Y� V�o���pw�Yx:%�)�j�ʾ���*�Տ֥[��u,t����`�UU=�x@�������O�n	�D��׈-��O�n�ll�Z��b�V��级Ex���Q���fbx�jb�4^TÖ�H�� ]9DFj�.�%�z�ɒ����X~�s����T���}+��� pW�����ٮ��({��Au�����m�T�p�������#$�1I[3����$8\�8os��n>�`��Y>�Y,�9�{����_��c*�'Q4�yϩUM���s藆��<+~�L`�"�{֜����g�HT;����i��䈬��0O�>�[5 T��*g��
��li���⎜��/��;u����+JoPa����˄��j�]vscFb ��ո9|��������(Zީ�ۜjW��8`n�6(���_ �L���-s�F7c0	x�6:�`W�ٔ���M�:\-�Ҍ}�;�[�������쁩0B�hػ���%�2m1R��u�Wd���p���E!�g�۔����H���;	�o�Y��+�9㲍1��f�����XM�!�a�h�t��}�dH��t�M~>cqf�H}�%v`��΋ߥ������XuJ』EΪ�ɍ���vS����a�g}��e��Ud�`��������OdC���c�(f�(\�,�F���^;�Ke�=��
�]�{���=���J�ι&�$�p�����zf�269*0l=�g�9>\yE���b�� �=c�ຫ^���XA�zG�#�d��8޸�[�~�F��韶\��� (�R�U�T�~ ���疯�:>��%�O�{�@�[l��⎏b�04Ƹ%���2ð� L������c���v�|�5�����1�g��1k��������B�M4���i]����s��>��Q�U��,zB\,ڌ��^,X���[LA��/�|�X����9K�L�v^��v��urŘ�N�
+�����r�O�����ڗF�YoM(4	���NoS���+�ө��J�+�:�p��gR�/�i��B�mtC�����0�p�k!aڙ3��H���NJ���/vR�}��򝘟K�>W�ag��dc�,w\i-�P���K G��Qy�l�Qśv�a�(Ӡ��nj�k��p�P"b�/�7�pe�x0꺮��uo'������`!���p-zkq
��6~Q�����j���oE���b�b*�*�C�Ζc��5wP|ٞ樳��˞�K8��{y!:*��/MX��<}bqk��+[�r���<}I���woQ��bc��K2��w,������O�O�뮙�^��� ʭ����|��q��8��=0z��K]ƠCE�G�j���u���^�gJ9�{�ً�7h�w_Yw��t�{�:��n��u���~=�,Q���X��u��~�&k�~���v��_s���x�#�T����붆#��oZ��L\^��'{��Z��ݪ�#��Ǥݣ��b�{K�����;p�b*�!��"�e��s:�T\�9@��g�h�N�O<ѹ*�c��J.6�~����?��ke�M��ʀhþQ�]c@<�`G��K->n��v�q�7,�`WU��0_|�p�k�ï33-?�Xm#j�Tu]j�Մ>��\�]��Yt�AHJ���vJ͊S�ݹ�n��C'umN�B��9v79�o@r>��t�3��3������˞}�����`�M���@�?8mg���p\䉍��Nu@c>�eK���@��q4@�Z��T���vJo+}��q�qyQ���T<��,1��_ؤ����F��ؔ0�i@��wG����;���B����o�(�k��U�/9`)Ү��8����9�&��a����i{�(3w?L=vi���z�
ߝ#��j�������Ze��"�ktָ�5(�6��n�� 4�8|6E��@��4꼑f.��W���Sǯ�U/2��D�8���{��)/�f�ր�H|�+C���f�v�E�ߵ�<-��0��Šǳ��T��y�՘���L�+X���ꀣ�HP�z���ź��Q�,F3P�̓��vV2`ݝ+q��"�yD�I^�'��UjB����}������xil�r���g�^���yfҬ�Z�����qm�	iWᾺ�q����#����P�}b�*�!~�=-3�c�0�5]y��A>�<�����V�F�j�9|�ub�GyY�o`!v��K��t��+�jP���Ȅ%��������sއ���V1��o�˾� +�q��^�2��)r�8�W���C�<� .ئ�����SM�w�V����;R�h�&�ۤ�*��]g9�)ƅn�ubd��VN�IJ�-��3�\�wyI��<;՚�h��K������hw&|�5>־��45�䥪����]X��un e�6���^�#4�p�S��3�`��$n����|�!uP��v����{�9ڙޱ\C��݉�-�qǾ�ׅ1Z:���\!�9�G���U��Geu�pǺ�w����� ��M0���5B�~���(��,꿡���3��K�wO�����8�d��OV���<���}m�I�t�x�]��4�}�m=0�1�� �ðf�F9r���ۍ�����.cډJ�ו^p�j"�0膼�P����3<�g$T*�zY�Av��g��M�f {�� �T�;7/��M�lƲ`��b/��9��)^8���Τد�L� 4^����M
�������~6�G��tߊů8���(���4���>�#/R"U�Te�Z@�d��~�b*#]�P (߮��_g��qtf���m�NQݳ��x�0V{����+O ���U��ʄ�]�R����c�?r,�땾���#�+�}!�rs<⻁�]�n!�L��u��4�<���[@�qꏭ��hv��[�ĝ��V�SWq���f9Y����*xC�O��đO:�o0s=�ݚ���ۚ�*J����l�{�`*�s��f*a���cC�5�}ؠ�=g^���^[���wi�:�i����l(רLлM�PV���,k<!7�<@��Hp��y��{���+Ѹx�Q�uk�k��y�=���m�{i�$Sw<�Ԧ�]	�i&1�'D[�9��;�1a��F�np0scyDC� �|V�5\I�N:��>�[��r�c�a`��i��>��c$\�g{z@��^fw.�y�<�[vUv�)�}�ŭ	ʷ)�;Чf�-z�W���Hu�Y�0��7_i�,e4�:�����ѝ���^��Oq���!�VH�6����"\d̏�dk�Keg��W�DQ«_��충�*k/ށ=���p�a�?2X���N�*��μ��xS��`?5��7N��-�����7wޥ�z|��WP���}�P��� ��\+>�qT&��`k�C2�-�.�p� 7>�\οD(Wu�����:�V	|ǘ��3�Ka��"��k��nK(�z焘��8`a�Vv�g���	��0/:L��a��μ��·���"�T_�1n�R�8��F�uN?��6F._ŗ%5�e�<��y�ٻY�KBT��'��3�fE˺�NÚ���F8L�C̣H�Zѳ�X�^���eK}n`��s �[������C Eg�F�u��h��^��d{�I��8Ov?���N�.�㻹G]cJr�mx2���?,0�pK7ٖ;@F#�=O׾��sa�xJ�M�{sU�L�V]�#��^L\����F�i���ǵb/�Z��߁ꏻ7��m
�X'��	iL<.�
˫��Gz�g��	ʀ�ʹf��z��Y�)>���▫?>W���!g!X~���X+�-g> �b��������z�k�i:+��p��Z2�xt�y~ӟ*�ha��u��=�Q�6���M��Lܠ�s�,��wa��o� ���}�]Wrт}�e蝘��(�`��K����q��2�	��;&=[���O݅��p����䄮��ixj��·��c��2����>�ŝ��v�=kl�Qw���Z=��ǂ3�f�=����ԺqL�}BN^���{'U�c�|���`:��Sվ*Z�5/��z~�Ÿ} ^�>q��Z*?�� "�c��~Y��ʺs��Q����Pv&�$o*4���.�T���5�B]8��`��0�v���ٷ:�m��+���ʸ:�#:��[��r����6����F�;�������C�ե�875��92�ڦ����]3�^u�{�]Zh��v�!�����\�����tCo5�r�2�l���!.=���Ǚ���4�����%��L�����$C���T��e���㩳��*����2�k]K(�ט5p��֨.�ljM��B���'V!};D��/���u�͚�!.���i�[YC����{_��7�*m�nF9�\�%��5���8��sPۼ���j�E8� ݾ�;�Rj�u���u�ٔ��J�T���\��,���'N���m��P͢���%������ ����t=�LtEL0 ��a.��O�(�1v�KB�ә���)�͞�w�Edt���+�u�,���;!%q�pQ��r��p�2m��u�]�t�+y�/�WQ�|1�2�r��_I[�Ա�bf��픆� �%�wu�$����]�]��>���vj�1ӝ��-	����{�V���aR'z`���Gi9�R�*ZO)N���k������t�������^>���K�d�-�O�w�wL�bR
�G됱WV�����N�*w(�Y�GoT�o�}�]�i�#|��BT�ﶎ�8��-�f�&@�Y�4rsz?���{30U:�C��_�R�ws�F�#+����FoeBSo&��	�*�4.�o*�v܈貚��=D�����nq�oWn���c;��-�gv�IQo$�m]u�=������- ��yI�G��Ez��sp�elb���LH�!���o��ܬ�9��=�{����̻�#O{1�F�c'�b�a0/�Ļk%�X�l㖖.3���5b��n�Pv����}*3Q�����'|'Z����M�L�7���$�#��%���bX9���eWgWK3�gXV��!V]�;��3*.R}SZ��4i�$������+V)����+hnn	�`7v�.�Y�B�(��������:�!�P��>����1W�>f:Y-Fv��� b�tVk�#�l9�'-s^s��3ǰX;h$��-#��ll�+O*�w�>�"A�����V 7Lm�uٔ{�qZz'\��b��Ltu��[q^띌a��EF ��\�_'uBa����R�6�kV�3b��p%f���0���a�eܴ��(в��ӵ�r����(D����F�Jh��b�Ѵ�Gvtdک6 n�`��7��8�W.�]gj����!��^��XN)�̶5Υ���1!��/N�1S}:����W�U��m)V��P��=�a�;V����K{�5r�Ju4J)��[�����l,�&�:�=��}q3溘I��*u��Un����XU��g�!��
҂��UB�_:�˖N�qpĻ������a�D���z��G����B�wr�t���O9��r���wJ�)�T�"�#+�N\#��A<�Qp��U���B�ZI�r��y�P�Rd�^���AUeIw��Ot"�Q�����H�DTQ��K�*�-uĜ��H��(��Brp��<8�xG����Wt�+.�拺;��洮N껞����*[�㹲�''t��I#���z��w�{P;��*2�1&W<ʽJ�腓5�4�\���e��#���rT�UA9���n��y�Tr��5q�˚.#��qʒ�D��z9ݑUz�!&�ル�F��UE�($\�h�U�^��$�>��E������.�9,��+a�t�'�����nwܑ�Z��F�#�{%*������_�V8�@x}!���~'�©��ݲ&��w&�w�����������)8=3��>��P$��G�<*I��?�<&�=��^UޓHO>?q�7��|vB#��orN�Y�7��kZ�"#�!�*o׾�oHN��y�����xv����ό~y�L.���}�	ɾ������}OI��~��.	��ǈ����@�I4���P�����aT߇��Vn�7J����L�F���H�"<�0~<G�{&�o'_S�oHIϴ��Ͻ���;󴯟�����7!8�}����`�'y����9�����ǌ�xAC�^����l��w��y������E��/'��7>�N���n�F��G��'����w�ޞw���}I<�q�OIɾ!8/w}�����Î}�����N��?w��y@����+�4�w��9BM?S�'��;���o��� ��f㋗�Y�.&�^&�3;�葧i��Wԓ˷����|ohx~���>�v������[�S���|����S�aj���?����۟�!���$��}���ߝ�@"��C0/�a ��w��i��E "(}��<!&�����o�w����=x��M>�÷'���$=&�ROv97�'ӷ�����C�kϿ�7���L.�?[rI��������\�Ǒ!�E�z��Z�{�`��!@DB��봄�<����7V���xM��yO)�S|O��!�������A�߽�r�����s�r��'�_~w>P$ߐ����x{탄A}��.w��-=�4�p7����N߽��˼�H(~K��z�cʸy߾x܇������P�M�?���<Ʌߓ{y�{������0���P'�ސ�zB~���!������#���މ�In3�,�C1����#�@�I�����SI���ݼ����O�����4��=''����|��Ӵ�뿓�������x�������s����i�O��?�G����{�ǻo/�>�㠆�Բ�ًQEmr�G�s��w+�||;�ǻ>�Cד�P�$��Q���ߐ�	�����%C�<��?��_y������v���zO(ri��ݻ�x��<!�5�����nBw�F2~����Ǉ�z���￻���%;����g��۱��HlA�΍e�r�GB���0�x���
V��Z�/Gί���2:��GhR���n�V>�w0�b��K��۱�����:�L;9P��g������y�X��n�C��W7�XO!�8�7�F~���~��>��Ü��?#ǈ���a�����$��Wy�mɅ��׸��S |y��h~O~������>���pzO)��׻r������ǅ��Aw��!>���ў���ǯ���g��gG�"!&���ű;{C���	��<��}�z?�L}C۾!���s���z��v=��{C�c��ű���o}�N��7��~|��a���Y���v�}!� |��#|BA�|�}Nw����ݿ�=$�;����I��I�z�����q������P���ǯq���o��;����˴���I�>;{y7��?w�?�����]�����#�x}�{��f>�")4�?w�y��?�S��������a|~��Ħ����}OHy@�C��������;z�'��P#����P��@=�˿>���9b�<]��}���SN?��<!�4�On=�����$>&�x��Ǆߐ�������{��>���ӏ����9�]��}y_g�=��a��t}O����&�D����$DD���bV�������ϿϿ_�&�yCۼ'�ѿ��aC��o������;oV��ߟɻ����
xM�	<�߿�}v�@������{R@�}O7�<8��탙�ih}N}'�~��˴����׿�||�G���ׯ?z�����bp~�����1><��`����C�=���]���=�S~O������M�	<���xy��s���{9'o�|v�﯄܁�/����DC�ȶ�/�!��.�QJ�W��?��ߴ���P�i�<x�������(�.��3�������.�o�O���<���gӷ��0��~8�����?S��ѹE7��ｼ����n�L��p�s݌ϳ�G�D	$���y�]�q���ό���8���[�i	0���P��ʸy�c�xC�i���֬x@������~B}o���Ǜポ;N����𛫱(��-�_%Yٌ��#��"�����
aL/��;���agz;��N�C���S�}q�����&��ǗxC�<!�<�,s�Ă�v����$�P�|��;x@����|>ѻ�n�&��$���o��Zk/.�hI˹�5ğ>��� ,p�r��5�?a�zVArD^�ݷ��̺C?=����j����V�h̘E��9on)�˒K��G��ј�����-L�����Z�>�|������W��Ǩ9��~z���|�$�?'?ۿ��N����1+�^>pxt��w���>\�������{O��ﯣݏo�ߓ�s���� ��">B#]U)���������a|��'ߖ��÷�|{���_�>�����E���V��n�xLW%��vs]M�<G�9���l�Ҕ����a��V�'Z,�Cz�hS�I�2�R5i'��f��ӛs7�����z���ޣa�Y�@[3���v������Ú�f��3ђ�+��2�u���~�E[���G,��4�U��1ױ�����b'�.�L�8[>�����e:~͕�$hٯP���e.Ucg7F�ɞ7����$<.U�iǅd~�fo��E�w/6�޷�'k�ê�Xx'b�#Pq�������#�'�8������y��Oep�r���{�ੂ_[�\��a}��`>��wjB�UR�� �"n�^����V��/��v�kaLPǼsI�N��h�޴D @e٭��; G���p�t�Wn �
u^��E�]��j��6s��5$h�u�G���(0yn�3β�׌�����C��Iv���Xΐ?���[u�;ۻ�)æ�C%x-�]]�B��%���e|f!꜑]�u�S���,���U�+z��ӥuw:p�v�v�%��o�*������oQ'�З��ΡY�;�����W�zC�=W�;G��0+%y�$���9��0�̩o�~U�:*�Rv��6]b�cY.hxm�X~�yo	^��
��6��F;��85�x�6X��6�^�����)�Ӝ8�+}*��D:�q�u�Gܥ����Uo�r	D�	(֊ӈ�kz�p�Pp��A:4A�L���unPH�6���V�H�+�5s���{��'+��h��=@Q��
�>ݽ�@c5�ː"C��M��3����
/tg-�����۟^}WJ��Qm)�cdO�aFӉb�6e����t`���AH����h.�w���!�QKE�(8rUZ�³���yc��	�(����(2O�j˥s�9�m�M��Э�].�^�(8J(]N^p���Q�o���c^�g�x��xڝ��{�gڏz(2��B�^T0��c���].���V~�|<�Ϟx�^�;;�B���5�XC�N��u�l�����Nb��ǿ/���)A6����^ɹK��g�qq�='�]�}������z�����~������������:ur���e�F���[6�Pg��c<�a �\�L�U��+��rX�vR���x��;�y[5�e\4��{��7�s���y'�*���޾�>�r�B�b=��U��_M=Ơ����!րVlC�jLõ�>�?%~~����ަ;)�����n�`#��X{5!+b�K�W;��h��,R�؇�=5�Ȼ���m�G���[eú|,�����s�����Ӗf���t��g�����ߧ�N��z��[��=܎��*j� ��Y�4�7�z�N{Sdp���#�_�`]�.�դ�~��ګ?wG˨\�b	��`9����G��9�ӯO<�.R�uw3��i���H���-�f�ly1?f�S�"̤*	�bQ�6�(ʬ�;����O�cD`�j��Fm�LS� LJƋ:)�eu�K*�U�C	�)���]��EQ�%�-��?X$�d��5�Pߨ���t@z��9�D�`0���{sx�5�րC���X5g��{��/��\n���-\����;��f�D,�Z(Vɾ�y�Ţ���bu��?��ܷ�6/N��� V���Cz���#�Q3�R3*�F�u.&��⩱WW�r�׊�H�@�B�ru���k�)��ر�[oz �[}f�ܼ�[�VX�5�i��R��x3�3��D�e-K�5@�y��`�!�iw�U_}�kG��ͷ�O�?�]@��d�@���A�,�KU྾V
5���2)�ך^(�Q���\�}S�����9����u�=){e{M���}.+�=�YV[x��������Ρ���(l?�*�4�,���E	�����P��.��U�V���ns����ӎ����W�P��@*�<DK�x:ގ�6>?o=+@ڽ>�%�;���_rc��<�'�x���a�z_�҂�]�C�^3;�|����iz�3Mz���za�+�����"�}j��q+�*ϴ��HU�����\=�YI�c�I��Յf:ל�ެ�����pY�dֆO�{��qzi�>:ޯNx�GkM��:���k���&����Y� �j�U٫�B�����l��Ԟ��z�m���a��q�u��"�z��o��6�`i�G�a�0g��Xɜ^>��y�����=�e/vs���(K���X���N�y[�:|-�g���hk�*�}���+6
�ABK��/o1��L�Z45�h�=��������Ұ�t��'9�W7�q��Pcwpn_7I��!�2�9��ל�E��4�v)Aϫ���ݥ�,m��v���/�`W�L���!�Zظ]��g�}�UU���}�
R#�B"�t/E+
n�=I��z��6���(���G@�%��#x0I!V�=���t���N�n�??�tqz�W�1���x��u3�����̼��:���e����\����>��쬂�[`R��:�^wAp�k¼�zs��ߝ@M�wj�/qc ��/���T-o��	���^�|�Q��y�./o���1����D8��ش�,B��ڌS��� '��"ab��������7���<3�~�!F�)��BǷ#<q��0Q�2ø�r����Y�*�U�1�׉�JY
N��������o�x��/��'0�#
��|r�P�]�pJ��M�0�W�
����pD�oMcv+ҭ@��=�Ta�l�B�t�
��/�0�k�ڍs~���.f���W�b+����"<!�>�r��Tý@_�:�:��xV���J��7��s�x����7�p!^`�K�X�U�х�C��iO�m�<&8�}):O����@���1A���
?����F'R�}�J���]�r�;�����r`Be����t�49�kN�3WV�o��O�=�(*b�e��=��**}�qK��0�b������a�ZS8b��&�E�ȟ#ה��vo'|9��C���
'����ꯇ�5�9}� �����m/�����k���v!ܢ5�/O�jU�D�o�ghK�\�Q/0S��匲�Z#�P�}�cep��L�@Vz�x��WT�@3$�<|_c�|<�r�ަ2��\Y�
#x�j�ef���eWr�N���O�'�/�rDH���CPv���Yp5����4��s��Z<)�=�E!g���Y�*���עq:'���(�RO{�@��`7�ǹ�Y<�%�i�7��ţ�M�;���*�:]�αm����}�U�>&�j�����X7<�3�`a�.�c��c�xf+��e�സ@y����P���]Dd�و�wLQXbyr�i�mQ�snA	�2�N�0�2Mfd��!õbc-N�-1yW��r���@W��x�d*��Ly�%�d�H�^���xw��UTFA���:�l���| B� k�h������HRFA�����5{����̟zZ�)ի��<<�*�CƗz��r^��}^�Nr�.�ǻ�`j�hR��N>q�<L�z���9Q���ܼ��*t��+w���KF��p�6rȝ@��󖯧a��UV҈�{,,:���Ϧ�������`�+zWG^`A��n�ܽ�V�2楗G2�oLk��P8ΖWS��_}��Wಮ�����0A�/a�VT��"��*�=��;�,ڈ_n&�
�\ck�޼!��{����v\����-<+E���*�(8R�9xQb�j~?=>�u����Wˏ9&w��c�T-��"�n��R�1y9(�?A��]"B� ����p�n�e� F�� ���ٿ��K��'��}����J�j������o�o��r����}Ok�����#��@]f��/�U�|}�c>�F���gM�j��;�uЕ�#��_���Q�$�4|�4�|��:��_h��8D��\:�a���ޔc^ ����~ɓw������1�9FC�ѿZU�����E��uow�}��s�Ws��?�yW�gz�w��X�*`�����1a����{iͽ�y��˯fK��N�i����p������E�l���0J[l	��}�n�-�p�S��k�u8���4���C�"�5�/޿]c�O�c��R�)F��c�2��UyF]�������1��>8V�x��7gAWȜ��RW�u��5_%abV��D�)��͘�]ǹ �(�#���ҭ��3�jr�W[�+J�2��oL]���awu]�'!�vEV¹��|�ھvU��LpdG�+��������W��}ZV�׭v6��]���D��m%(mX>�͢�r���h�Ή�s5�YRkb�� nL3{���)�M��X�5�3�'�g ������M( ^{A�e	7��4�,��?M�G�<�3��@bh�>��X0/��W=^|���*��PC%�E��7���>�h����Y Jh�	����9�"ё�����RL(�~~�!���9��VSa�N��z��|���@?t�[�}�QM�!�,�Y��*�X*bhcޝ�b�&�|�&�܇�A�#�oV��!L��䔂�����ǘ�S���W㢷�5xN~���}�kȗK����@��g��N�[g�K��o��y�-�a�i�����=�5=ׅ�O�����X꼝�y~�da�Fܦ']�({RE�ț�Qꖮ<���uڨ�߾{�Ι���~�/�a���-�t��=�B�^�]�|��g��w������8*
��=<�C�L헇p�~L}��B�}uv5�p���ƶ��W�m�fm�yBﯩc��[/��S���LI3ϑwyVy��_�6"֏�M�ҵj�w�(��F{bw6���7:=�!]Ƅ�8�+�!��z��֬p�Q�m���}�qә�����;'u5y���}�����j���y8=U��-ӄd=J֕Z�wW�cM�	˭�y�4q\^��Ԗ] ���m���gkv�ʛ�73�/��ѱC�ڃ�	��B��b�_b!֎�ceW3J.8�������>��V�H�%
	�)l4M��R�#!�U�b��>�ռ��֎��9q�RŬ.��R�+��С|,�]83}�q�r�Ӗ��JV��Η�\G_[\A$W�%�_|a�I/�ch>"X����r���+;��HV��(�� ���K2�l-���깏���x)�ap/��oj��vrʀo]����l��@L�y6�9��زG�8v��)�F�"�J�+�8i���po���)�`4���6��C6u �j�vV���RnU�ws���$��@k�j4��q��X�Z�U��E��$Zj�Y;%���e֣
���X���*?���,f	u�wŐ�7�8���ks4��$b�&�fU�W���7��r����*5�Ogd��O���k:�<쑷�����j������+��R6:�{]t�F��Z��g��Wn��']�&1-���uˬ�E+�`�#�
�c����o�/wB&o|�I�ݰ��WC�Ԥb�z����3v�p��1�u|c�V���m]����ķ�u
Ut9H=`�d��1tps���E����gH�Ha9���%���Φ��z>arM�(򷭾��|LT*R�W�Y�q�I�hZa��iUf}t��N�r^�Q�{z��+��dz�Y��2n�+��s�a�6�X�˃Tf��������4��AL\�r�rn�^��K�̈%�v��rK�YV�k�x�wjwDt:�\m�U����G�B�h
cn^��sF�=�*$n��ʳ@����YZ��k6�qȤ<�d��l�/YJ��� 3��8)�R���T$�C5ݷ6� �zU�;�����kg)�\5l��-[#�\��|�v�[i ��$�oZ�p:�4��Vq���@��ծ�>�9v�Z M�[E�6IHh��C:�&��pQ{B�Z��gj��[�sjM&�
o+2
��c=�J�)5�"l��v9*V@�h�]s�t=++��\y�बW˛�΂�sut慦�Hj����L��;\(r܈nu�ժG,��e#�����(�	w<�����-�ئ$����dpK�I��%���֫�OKC��1�=v �ON�m��tx!�Rӻ��ږ�k�R`Ip��>��/O��������g���.EfUEZF}$��$B��U�Ȥ ����Nz�V�]Y��L�!�(����x{�we0���|u�RK��Ȋ�ؕ3E�.�t*�Sg� ���(���ׄ9�'Ux��Xhrs��!*s�$�����"�:BJ���q2���D9Q�**��p�ʏ�1�*��u˞�wGX�r���AAd*3@�Q�ؕQUȊeEq	�D�Q5L���ɗ�p��Tj�]�G*�L59�'��A"ةN�<��R�"�fā8�jI��¹TT̙d'a24()8AAd4��2�Dʎ˔�UQPQArPT�,����șEU"�]�QD+J�X�SL����4D@�� ҏ���+��{"�g�����wi��;�m�+�hB��KC2$U����V虄]�7�w=X<x�z��������ž��[z�����R������p���7 �m�\7�J�Q<7�F�C��L���M�}��5��5l��r`�C��Y� �m.U]���(&���|���f���=���kT"���ڣש�]��h�_9��d�����N���Ƶ�;�Ȧ"izW����}
~���o�*za�s짞�ªgEp~�v%y���ܡh���Tޮ�,q��W����S"�B��Bu���d\�L��ZZ>.z2[��\D���[���W��ah�%���?�tud5(V�U=�/ک���˞}����$V..]v}��OA w��3ʗ�d�lu�N^�t8L5�^�ǀ��(ೣ�x��A�Σ�������z}J�?BU-c�n���*mD^��+��7�͙�F���+�����U��y�B (�[�,����r`%"�<�Tk���;���2����~~ك=����5���Y��ָ:ԋ3�`aFl���b_�Q���O�����Ei0Wu�ds7�������h<�I��f�;J[�m��0�kn�^q��(��%\��(��9��5Z���ٰ��H��Q�.ﶲ�Ӽ2�iln�u�&��GW�k�\6�̂+3̾�N(f�_om�#�ޙ^�qq}��_UW�Oj�=��nR�,K7��a���Tk�zUi\ i`��b/���S�L1Z(j�lٝיݻ��B�%�������C��i�\�*�OS�{�o��ȶ��Q��w�y�:��>���V�:�+�W"�K����!���I�9�͟?_-X=퉟x�j���m��]s �s�5(:�c���q[��\�;
��1�;6wkR�+�ʻ���:�39Yz��\}(�g{�X���C�_l���=�io��Npu|gw4Q37�°ƬCޝ�����ҝ_���u�:��z�oe���r|�,w�r���{��B\���꼾^�~��g�}��xos㩤�/���ڋrw��oo޹5��Ы)i�p)��=�_�z*{�_�q;�g�;�a������Ҽ�7^�~NΖ�;�c"����*��tg�>�go�%�W�U�k��Arp�n�q�D���(le�j�Jp� wh��c�<7�뺝~����{��âr3���4+iQݓZ���^V9c5���4���:h6�\��t�;�{�5�����W��bg�K7MNzj�-���������r��rP������:���E�ʳ~Yrnߨ�ޙ�yl�hEM�K�5k'���ڜd���N�18���38���co��Y~^��4w��u5
����_b��uga���â�/'/7y�x����Πkw�U��k�8i&3�x*��-�y���z���^��Ǳ�<,�\�O#�K�V�������34��7�ö|��6.�/u~>�"�?/N���@�\W���Xx��� ܡ1�ښ����m��q�������L�k����7�e}�����Ʃ,�R�#S3�Xh����F'qk�̓�.u�LF���!mtV��*vY-M�߆v<���x���.��e���5e���/`eDf�t�˓ݍ��Ʃ(�e�t���|a���ȅ�=8�1���e>pL��kX������7<���N����k��j �梽��lulP�NT�@����Ue^Q�VN��>�Ti�w;+��g2"v͵
IE<����>s+�a�T~�7(�����}ֻZ���TF>��N��Aumi��\�]���A_λ9�J�ݰ�=�.Q+q��Wﾯ�着����{ޞН���Y7�d����}9���Y�?v�Ĕ]�EVw��Ԩ���,��<j���PUo�#�3[2�o���M���$
��]]s�H���Y��\c;՝ݒ�ֽ��J�t�]���bM�vR��3-Ɩ�-"��ne�oz߽Q�n`;0�-���_
ܧ*�������ʮ���o����6��tJ:G���Ԥ��������b�:��0���;>ua籟z{�8�y��V�F�[lg*�g�������q�t=n�iK&ϽS-@��|���Ez������v���lj�Y0c����/'|���LlfN����A^۴ډTW�ژ���@p�w���F��P�Oo���2�xc��+��w���3��%���+	��N}�r�W�xגnf���Yo�6����<�����5�֢�o��\�e`�Ɋ�*��6=ϯ�a���(�9[V�b��@71��7z�r���ҝF��j��r
R�Z��1�cN6��m?��Y�m�{��٬�э5��($阜�%��ϫ��K�T�rr�����j�Y=}�o����W�Tx������߅d~��>5��;�����r�������s7���`�٫˻��=M>�]�����͏4�m說E�~#nh�i{��c��{��.��O�A�\~�G���˨�c�_P���ϧ�z7"�kg{n3���{������;ok��Q{6�^����'��;7��;�|��rOi�G��������8q��fֽ��߈��^��v��2�p`K�;w}���ySh���&���3�Vv��]f�����^��5�w� ^�!���|{�{��پ���+�ڿusH��Y ~���r�9y�6�S��q�z��f?�s��u�0�3���)zۉ�b�&/e�u<�s��~֭����2�c;��ޱ��zIbg�z|��kחZJ�hـ���s�\d���^n����X:��¯SۺK<>��RC�|7��*>{R������ �|�*ڍӬZv��q#S��3ֻ93Xx^S~��t�Z=����jܢ��ȫi%Nw�sE8��w�^fc�ݑ�/�7h}8��a\��6��{�u�;?W�U�}UnU�l:����9�bt��1�?3�j�������zV�;~H��9K�|�/Ҧ=�}�cu���[+�w	�&��jL6UJ�����_t��r/�yJ!��#���#r6�C�d�Hy5c5 �j��`�|�쇊,6=K�Dg�fj7���܍���'��@�^�S�����}4�ܺ��\�K��l�|����-a�֙�y�&�^��juv� [�� 2�\:<���ҩ[K�����:����^ߊ��y�gZ�g���w���?w�}���9
�;�u7�v�~R����+y��ƽ
��p��(�=�[��z��ע��r�m��\drWsE�On�V���څ?{���vqs\��d�"�쯇Ip�7�֔_��^���wVΥ}��V��\����ON���1�~}��gN����H�׀�
�9Rm��ќ�qgQ��HjA�3�W>O�m�E��3o<=�=����gV3W@ڷń�����3��"�x����Q��������h"S�[�o1W-Un2��}�u���p����ع5s��\RN����l�0���ﾪ����|{سH;_�[6�d��j�\���<��1I� ���ݿy�Ѻ�YuPo�b��_Nc3��GE&��_s�y|��~Ђn^^{�;�����7%zW/`�8���5(�j-��A��g�V�I�O�6I�{����洯�r�}�H����;韃��.̗�Ԃ@{��uv0���~
uy[�����=�RbZ�MMfN5����{��A��^>��M{{��M������f�����Cڥ:N]�[ۘX�����5��%Fk~���Q����'C������e�j+iַ
�ȸ�@>������WL�ֱQ�5�X��>�D��<Un�"�\�_<tI�y�^mL��|�|����O=趈^x�@:�s����S��S�}W������Tj9��@6���1�GVi�}�*]vT�;��6P\���t��&)`yɛ֭�F�B�����kn���Y�!�v�`M��T�w �ڻ��l�-Jt�Ŕ��Q��&�l'�c�n	r���Pt^�բ*��G��po�%��\4'n�M~��ﾯ���L�m�膩Fz����L�F������\f�2|��[���q�;ω�mxI՝��΋�R�|�	����s#(�z+l�aS�R��.�����@��z�Y�<�)�.��<uu'�=��.�h
Q�B�¼�+|�m�{ڥ�bH7���~!v�G�;潙O�6v�^���|8g�z��}α�������&�!pvm*{?oA��}�9�>��E���'oݝ�\.O{8�5s5�VeU�Q��)�����
�����j�x�/����^���_{Ͻ+L�+�G����1��s��3"�x^3z�V���;�g�ߟ��s��t�ōܳ��(�^��Y�{-�)��3�=UVrb��v3a�r2;�=wA]�a^��Nz�Y�R�5s��ȹ��y���k#X�����A��v�J�n:��Mfu�"�bW@+��8�3�����Vx^��Z���j�͡�/*JvuI�d^;�@ Tڿv���)t���"���M3++�[�cX�s0�Mf�`���Xvk�Y�[]��lq���(��������u����^�~����x?5����������ٞFV����ޏ��<+���Ôʘ�d-�nY��{ ��&�J��=���m�8z`�e��ɉ��}Bj�5}��ě��
�������]��ښ4�TPۯ[w��ߦr'}�a�[M�*����[C��O���})��y�V��!<M׷�&�p;�>M�x���0�Sak���z�5�
��㨫��f����񭩊���.���*u�}G����{3Y`�8�������pײ�W�����/�)�m�>״u{iu.�c��N�����[W��[Q�{�\��6�ݶp��E�y��Z�mVl
~�����m����ϛ:�19U:�������b�!Ά�x��+K>�h��O>�QF�3�-7�]���\���f�N�}O�2g��W<�C�pO�%4'<�}T�yԱi��9t�z��/�ޕ����z�?��Y�s��'K�g#M$�e�t&gPs0X�Aޔ̛�]FΒ����u+��Ws3W������!Ւ~MM�k���)��O�}�G�}i���b��E�s��ө��D��yzP�ʺx���+��<�r�.�m��~C<��5�=y�3�S���mW!K��v��aE`�w�/!��}��I�%��Bs>�[C��΃h�%��}�q�g�;��~�v�B�F3o��{�l*�nYہP4sv�T�ʠg��7��ۄ�4sf����M����}���Y�xt�
�f����ox� ���R��� �[�⛱k-l��s��KwD��8�H7�_Ba�Xya�F*�J��//5,����M�Dy���9���څe��8��u�Ҁ"hɚ���y��W"�����^��pQZ�9��nc��3�)�M>�z���rs41�F��|�~����sv�ֹ )�oP�Yfqe��f�=E#�T��Ϳ��(��^^����[�$q���$J)}g):��`?ͽ�GbE>םz�vZOJRɼ�-Jg�q���H�h�W\�+4��K�As���pbkw��rOe�&񴍱��.:�8��3l�nJ
��=�>����1��2e	ݦk����>�d��FL�)<�૬��|�w�z9ࠏˢ]��
�E۹�����0k�8:t�k����3&u���#n+R
�6�twŎ�ߦU񡽼r��VS�t�^����-�\k�;�+F��Ky0��ʖf�b�����GP�$z,ǻ�ktM�l6V�3*f�@d�\����qi�ϛ
gd��V���w�I�ud�İ7��F�B��;gs�l���p��I[yH&!ɵ��6�U�f�#�2pV�Hm̹���LL��J��k+5��y�ƀ��a��+;��M���f��ђ鞩ù�׏ԋ!�z�^c�ɶ�Ϭ�9kRI��2�+0f�^XS�pF"�J�&�r
-�S�\�o2�o-�;���^],�R5�qƍb��ʚ1��+�D�,��J8���D�Re̋��"^�Q�������2溾	��62���+��B�9�����wr�izV�5��]K4�W�9�%w,�;�W^DHY���sז)��;J��˴�V��09��S� �W�AT;���&p8��>2�#έE= nb�fv-l�L}� u� ^�֭��|>D�9�QQ�pܸf_\WG+Ov��T@8�?up���^$�W�َ3�B�z���f@@�γC��D5�sgȪ���5�VX���*ngf�+
��ݾue��P
�_������;�e �@�� �����$������:��<XE��w��r�X�0[�bj��Vx�j<�N�4�=͍C�^��Âf�����V�s2�u�LW��1�HY������S�{N��h|�_(����R"k�e^M\�w�Ҧ�4�Wl��AX�.�#F�4�m1]���;K�،1��/�vnɴD�	��1�[�uF�pckvn7˺����FMT�/Kq&�oiKi#W\�p���}�W$F�Y��+O#�x9om^�)�PB�K��**�'+�Bt�-���i`!J-�l��b��kTB���P�CL#fΧ��9Cp��K�w|���z�Il�q[�x�F�5����.�I����&�,e�픦�����J#N�f���{�wƮ�q��В�O�Xeb�S���'^rF�h�F�mJ��X/����,-��ij�����\�%��
f:;^Ny}�mq����E�.6���=��l�ۖ�ywZ�꡻)���v�eϳ�&��j���̝X����Zw��P||��5E���*��ʠ�Yr�"�P���Z]�i�W(.Q�L�<��������YQB��䜈*�a�AQjF�e��8�U�8�
N�QTEL��T�p����RUv]��d�8'"
�ə�3mZ%����W8�A^eSi�p)�Q�C.\��2�PD������,����ʸ�p�(�V�hI�T�("��P�E{�E��A8P��-H8Iӑ��r*��Ue˧I����,�I�4iT�
�D�E�"�g �d�G.PEAT9
�7t'1����Y�ʣ���r��hEjr�AT\��M�8P�z���s���HNh9�D�@�(��� ����'�xGHH��eD'�5"��W`�m��� [�]�{��cxiQ�p
�������s�Q�n_�@�&N���g�����g��<���G���3�l�_�n�G�ժ�u�^�i�YZ%o�.%cR��
���w���3�{���W�A�w���s�[k~�\f�%p�m����m������uܠ�Aխy׻X��~��3~�1�78Ԝ8����v�η��r�I��,�)��Z9��	5�r���'��i��_�3���ʃ4i�$������Z�Q��:���U��o��d���Ѯ�kse+�E��<R^y��ᨻ��6f��W�)N�(��;��Gc.��o{F�=�xǢ1��[�աw&���ޗ���f����gۄs�{L�O�s��g����!�Ҟ�|�L�5�w�;a��s�a���E���
���ţ��T�0�%�����M{�ϵ!z�����iz����W��3Cl���UtDq���{���M_��m}��F�:\g�ډ�f2�����_��Ɋ׭�Z���@᜚�%�<�]��m�Cu�W�m��ŋuNY�]'�έ�Ӷ�Vci3p�d�KlJ}��f��"w�{�+՗QԿ���noc�κ�n�\��]�[�3��a̢{t��5ǹ�ګ1�*�ubME�磌�	�fw�~6�R�~I�Y��W=#r��bc�Nf�i�}�+�����n�tB�z�N����|jY�ׄma��k	����Wڧ�ml�ؙ����� O_��;�L���|�;y�ݛ��Ȩ7Y�7�5�2�\��n���Y)�y��v�.86^Qni�g�+�S6�ܘ�����c�����>>�G}�υ���`����,ō뱜�˽ׅ���yu�
��p񎻈*Ү��vQ������%�ۛ��כֿU��𧻓�}_Q��὾\~�y��w��vn����8�/="���%p�{N|a�!q�N��e/c��)Y{|��pg�識����c^�p�pp=�ӊaeԼ٣��=;�z�.�%��,��M�������f�0�~��*J�}��}�k>�OQ���8qk���
5繸�s7E�um�M�u^_���w/H]�����%��]Lx7Bι8˹��L���y?J٪3�AxK�q6�A*�s�[���P̲�݅c���W;0�T鯻DT���B��L�FU��X���"���^�Ro���s:H���6g�;�Z��������菾���'���J�Yٞ��<�}{i�mT��ڤ=~�J)�<s�U�X�:i�����U�۽3�c�ۏ;�g���j\�L��8i�,�YD�&�vL��d��o�)D~3�M�ۇ�ᕴ�i��۩r'�e���F{�$Е�{ಧ��T��m���g���� �v�]�*�~>�s�NVݽ*�]m�:��#s�3�ָ֢�w�'��z��u{Rbڳ<-<��Q�}����oV׶���W����BnM���P��ة,↽�`��^��<������b1&���0�s�*�a�ɸ�ʚ����^�[+P�VKw�W��Q�8CZ�Z�t6�a�s���y��(�-��{�'v�|�~E]�������^�;k�lk��vR��M��ݗ��zKWx�O.-��"�OQ���S�z�/���Y�n�byp���9��S�QM�y�:�]}efX�1�k_ӹ�ݩ�1u�I���J%����k*�.y�	�x���8S��(�1Z[y�Nݤ��FW;��U_W�b��/w����������}�EU<�����_:�>�y�#��;��kO[]|^,�<=���N���{pn�d�"�����Oot�S���wry}���Ə{�"�O}Ӄ�����8�����y:O&��O���|yz�tB�U�{K�S������[���Y6���9��tɇl�5����-��זP��h�Ny�>G����������ׅ���=�m��V�n3�U:�|=�u������^���;k�_�<��I���o�m?��t:�h{q�`�W:(V���w�G����9z�߭�N�OV����XͿ|�����3�V��^�^T�a�k�k�>�L��gz�W��\E���P��8����ctH�l��z�a4w��!����3�=�W;,�����X.���	��ō����^�v&���~����ǽ���N���ט]LU�՗Q�$}j]�BgR��O-��۬	uE��Fέ�;%z�/nE����t#~�6,�;]����	j�Hn�*��4�2�黧L-�OEF��2�Q�n�
Ke��@��&惪�G�܄(֫�'v諭���m9W��t�{��6���/���>��<{<9��x��SS��<�:��}V0�3Ip���R�A� ָFjo!�baׇ�#(N۶w�������y	yݚ����}�~�nc�T�ά�ze��a������GjD3�ÑĄ�R8�y{_TI�^��[u��{o����W3յӼ���;+�m�=s�t�}�ߧ|�@�	�|�?
p߼{�Ԟ�JuN�	�S��嶶�s���f��W���@�r�!����9N(��)�X��>�8oi��3nW*�c[;�=��8�C}Ke/�s����HI�ە��y�Im�������*��>�������Vv�>�(CO���#��$ߔ���kd�}�}��v���~����cno�:�W^R؟:T�|]N�96�&���ߏu�6���������[Lu���/��Vn.+�Y�fXo�<�i����vm'Rk�O�K�%�(M
��%�h�c2mf�t���l��@j�gW[׮^vX\aZ'{����]
�R���b(��������j����4N�<��FnKM�a���d<�����:��+����s������N{�6�m���tc�1��/.�ʴ��}��O�:v5:	 ����g�����[s���f��vN�1�=��	���� ^�������v��U\9]�H�.����7����W���=Y��p�~A���\B�0��cw9��4��y�"�\2A� �ZO?p�Y�5�N����M��q5<��,e#ᔻ���<�E������[�����O�����}��Wz�*���M<R������OTͯ8S�iR��|08�W>#зCM�?=���p�~F��n�9��m���}o�|����v�l�}��x��]L46��;�v0�� 0���Z�}�����ُ�i,��>�]K)ʞ����oh(��)��6�f��d�x�NKL������^w�][�oi>�y�q��4Nt�q��;�|���{��S��[�k��әs�Ҕަ�����k+��RɄ7��:��_'C�����U�1oN��yP&Ʃ�����%6���O�/R���+���w��g+�ꪪ��ɿu�6�����m�����um�5�^��g6^��D�q�F�ހ*.�A��g���E�nz�����p��B���N4�/��i�2��-z'��U�~�k^�i���@~��ٹ�Ў�WՒ�*���˝s���/=�޶�n�Ϸy>s:�1��������)��kέ�KG?f�3�Y��rk��mN���e{���7�i
�uy�n5�nxj��w�k5�=�~<��nOyU�sj��L�g2r.3^|$MzO�́�RY\��q��5)k����N�w��^j��3����K%o4k�"��똵��L����o��mf��^�P\��bUk��#}��M\�fc���o�*�.q:��dOl��z�i�r�瘔)��kdz5�F'	���Y�9 m\&Ԫ0H�ZM-w)���������-_����)�xt���x���S>{����
��U���h�*�5��*��F��J
@^�|�=�%�u�u���(��\��1+�[[Z�UW�}�Ս��z�`�0�k�:5�9�n��(��	�a��ı��982/�{��iǯ�E6����akYn6���KQ�)S��&�{�pw�'FV�H��^���=�`�N0����jT�r[�iW��/ ���&��)�K����R����oi��1��HBܖ�+};D~\fj��e�C�S5�d������]�1�w^H��;�kz��zȯyu��MC^���q+�Wďju���j�u�ג_��Û׷/}�����:p߫�������&�s��X&�!=�� ��~���s��b�OY�nN����n}h�3����y���;��ϰm/Ed�2��i3n��TVg�y�V>ϻ�v��߻7ޣo#�	�!�.gv����Y�t=��+Z��ҕ=�{����j>-���4=@Y��x,P�ݣ��j3⡀�0Z6������G������zV��-_j��衕�5�*\�����ӹy��W���;SW�(>�]�
�Zl� IS*�]�u��iǺ��3J��9Y�;�'�jRi�[���U��_^�j���{�K�x>=Pv���.��loirӃ73ֽ�1������&���_�kC��h?r��x{����Ev�6��4��c�zm�7&�>��x�L�C����W:����{��}7�[H⣜6\�ݼT�B��e�f�G�Ҧ�9�S����3}�N�X�N'�S�V�)o<�Dϱ{��f���nc�XF�y���9�����|����>�����x�B��
n�U���U킯Z������R�����n�&gٺ���~��_G�S;ݷ�	{����.���^��&�E�<$����q�PW�������ޗ�<���ґſ//u�z�\�^bi�FT�y^��"�{���\w;���J߇V��:��]��v�C������Y�}^���叨N��)�W-�!���,�)�^\�����(#n]H�����n�egL��=����m5�5ۆ��oq��ouuJ��ߝ>�v�<q祽�_R�Vҕ��`{�79�v�[/�eͦ���û�Ճg)�h�r�r�u1w�AB��mś����Q�����ꪯ��w����OV�̧#O�>��:����eeu�����CLz�N_/�hUl^�;4y�$�����'���n�:O.G�u���zT�γ��Ng솳f�o�m�Ւj��ʎM�1$U��Q7j���6���S��U�q��Y�vbw|_v�����U�E�QOs����y������0��3&��S�Cd9�f�8H{Τ&�zŖ�,��/����z]����79go�a���|��7��H�4��vԙpr�~�~�mE���߼Ǭc��9��ˍ�XG95�ӈ�����G��[�*���׹�Cme����L�u�G��lk�e9��;s�s
K���M�ݯ��V
RW��P��7̄}E�`G��xǠ��Ɂ����y�mTc�:���]2�����Y�A���Ok���ot�}�����X�qR�����}yw�����̮��Z��Nbml�� x>'Wc��V��ڢ.
o��ۖ�䙺�Xkv�u[�"ݺWp�N�#,�B@5eouY��,�#����X3���GLu!��,�V�I��QS�U�
C�@p����8$�����P{J��؍)���u���^�5�n�K����/q�n�X9����9�ǯz���3lܻ��4]�J*[*����$�h�͆�ww�n�ts�ԯ8{�[�_�.r�k��Wr���a��`�W���ʘ�R�d�
�frv�Sde�&V��wR���!�5{c�t���U�R��nY�R���]��Ϻ�q�ڸ�a��6š����� �iu']�Rܣ&*��Q��i�1�'��k�\��j7� n��=���#BZ�u,��A�_KtCpg�6���{N�_]FT��ee]�I�ᭁt����Vk-�t�
bPDn�7"���i����l{�)��,��#��]p��2�*�#1e��ۥ��:s�>�=]��7�VU�
�qaٕ֩�*
��d��V~О�]���N�����;a�w
��s{��������M{{�h7G;B c���Ked�a����<
�N��T� ����*mn_4J3w ��Q���-�E٧BU���;h��lӈMYbQ��Iy��Ҹ@�:��X��E��R��wN��˾��{>�m�9'ʭ��q[�k�i�����}�lU�b���)9�yj�x�a�NP�Z'K�f�n���`���a9��"嗱͹K�*"�;�Nƛ�c��Y�%aN)ZK7;�V:��̨��k�	p$��]]�n�hT�Tp���j�Q|[�j,����ʉ�1�`.����g���4ݚ��������J���flY��5(q1�#.��Y3qbht�w����]��+4��)h��7��h"@E����c�b�T���V,��Q-N�K�S7H�e6d/���V��ՙr��UĬ��FP�v�YV��Z}2��Ӝf��6wu�ܩnr��IG�!94�{}�]8*���p8�*�*��u�m+u��ʱ����@��(�{zJ���,T��U�X8�n�h}׊s�y��\a)U]il�o�[g�K�>��i�H����޴�;��X:/б�,�{']�.ռ}���E$e�2������[7�� ��J�50�I��z����Y�R��y���3F�����nMރ�*�{u
��.�\7���fۺ�������n+�`�.�3E�P�@��Ҕ���t����o���hf��\�ۊ�p�1[S�Wv�ɭ9��{ƭ�'`�O]Ge��yCj���^�8j0`g)��y���%C�]|;O5��w5O�5���,*Ŋ]�r�j[�1C�#�K,]�˔8NkJ:��.fO�W3K2��'}z��`Uf��F����*�χ>!Gx��4���F\����z.t�B"�����)�A�w<vS(�B�z�$��2�BvQ^�ʧ2(�<�
�]�.W *����*�vQL�p�R�ȪL���ҦRH�U���㛘EL�
U��T\��Gg9���샊��r*��s��Qr�5ȯJ9t��t�j(���t�!0�r�xX�r���ap��+��A�NȪ��9vY$ki˕Y,�.\�Zq� �JG!T�P\��.^y�8�EN�Er��7@vTʠ*�l��;re�($9����s�r⋙\�EQS�ug�LI2�D�(��벀���bv�!��E�(*�2X�vG��A
�Ԋ.��s�,�� kJeQȵ.9:����<�\�.��#�r*�\�]�Av\��z�H�R	>C�"������S���y����V1���I���QtOs��Ʈ�*��(-qWN�"����O��fs��\�h��d�~����RL���ՈO欌]22a��>�Od��<��>95�v�+���C��X@{ރ���c�o�_VWz����U��J��.a�;�}j�T߽t-��N�����n=�(T�������|x�{�e��P�Ja�{�Y� �E�ƒ�=G��.�ܥ���U�sy���`s�Yר`��}��*����?���]�|z���ڥ�*�����ٵ���|<Wyv��ϟ�Z^J�J����i��N?1��'K��̤3��U��]��󙩞�o~�Y6�2�5����v��� 2�]u���vr�z��Ͼ��k�1l������fW=��2㨎3W����ۋӻ#�TS�{��UO#nw.�5�^���CHT��Y�:lQ���V=��4��6})=����u�㞻uY�n�ũs��,F�Cހп#�]@y$+7�	R�1�Sy��ɐ��j����P���ҭ��ۼX����̎�	��;c{#��f[��+�������|T\y�[��}K;�g]�v��wE���Ms�Y�,9R.]c؂Ժ�W������R�������
�Ϸ��ϭ�6��P��½<�V�bt�c�F-=����2�}P���w��ٮ�s�2.fG��?��S�۫{֭b�/=��nL���g�A�*���d�^��R0���y�+9:h߫�{+���j��ȅ��{��6�W���C�n��ƖIo^)�Z�{CQ�1�F$��P�@X��C1�p�ׇ����'_��L�[��j/lZצw w����������(1Wz�����S �͸�?Q��}t�~�b�*<���kbq�ƻ[�4���ք8R~�*�ZIr���[Z9������-�Խ���Ө;^�+*Ҽݩ�����vrg�>I����ҠJ}����{GW�u.����{|r�i5lo��+����:��5<f�q[\ͽ��W+�m��"��g�b�����3ZMj
&��t��;���(�0�'U�VWu��>�jr^{Ǫ��5�s:�}��eN0|��#���/��Z�M�s��M��ǜ�-dfM��	��]W�Ǆ�.3d|�>��f��n�}WC9k����Rɫ�#�����.�����}��K�t�k[��Os���U:p����ڽˁ�[l!�z��)�����?I�½����=<_v>أ/�gmv=gA�]JG�K��v��5��fJ����Kٮ�J��gN��촖����oΖH��k)i�n�n�������f�=y[#�;1�N��V��O�H{'j��n���>����������Q���.�����.ö_$��W{~35�{GJ��O�/r����g{���K�Pv�;�ǚ�������B{k�3>���>W��t�}�O>�w�h��K���9�ū�꽊��I�����mk�<s�{%�Ө1|�Z�oU#7��i��y�}KЬ��W�þ�egM�z��c�M�S�<=6lcq�&`m�O��6���O:K�+��t��8���ϕTe�X,)��R�J0lG�~���
�d��'<��Ө\�l5e.��{����r���.\�'yԢ���e�b��]o�����U:����	9I�3��L;|[�)�vl>��)�β�k�,��V�L>���U}�A���x����/e���3��o�/u�E�������U�1�n�ִClJ���N�ɧ��&2wYf��K�%C��%ۻ:�R8�0L��b��\��]1�b�6q;��؟m8��Z�r�ƻ���]sC�tyrK����=�.�ԗj�>^3����<3�ޜjh�;f3qV�Ȟ���J�1h�y�<��;l�����x}o=��n��u]�r2����6��{��y����������Dvߟ4$��3ӹ/iթ�Ƚ,�������uW����Bw16�ͬ�N�#���@E�2o��/�SOu��7�����T��G|9��씶/�:Owǝ-�f������d�9��ߛ�o��ֵ1�1ｗ��n����9��9�ݕ	�y{�W��������:fL�@�����˽m�~j��u��+�)x`9d�����:��O4�f��n�c�I�e��u��yY�T>�F�uR�Bf<3�g�Z�/0Z��X���Yi��i�܆�6�dI�N���4$��K��3�K�����}cK�����Wmc�5޼�ƿMŴڞ��$��ڹ�p��]��r��{mv�����M�۲c��:�����L��ɾm}��~����U�k|썋�>�OXU��w�L���g�Ѵ����|`����S7Q0�5+"�u��+w�*\]d<�� ƷH�d<@��uo.�W�L��w^]���/�v��B*�Un�*�]�m�_n��F����y鷴�7K�M9�gZ�+f���?yk��6���ܺ�u�"+����M���W��fsַԱ���3�9K��~>���G��{�Ø��Ę�e(������D��he�c|��!|z��u,�r��ƻ�kc<��P1v���n����T5M��⨯�C~_W/��u�����z؞�L>�n�}OZf��<��#o�%s٨��D.�=;���=��v;�U�GS̈�ë:,�r��"ݴ�E-��Gʚq\�����1�7�<��]�0/D�S�Kj %�$8yF����NsHq>р���n��q6��s�ߥ.h�n-y�;������Kzj)�Uz/�es�jK�>���;�	m�s>�v��0�f5�믷lzz�h�N㴝[l��u6"fVN����P@��~���}�-_I;{6q��3^�%�̌��Ӊ��!�^�cEeL?���v��M{2�mN�}=�g��A/�c�;(��S]���]\�C}V��7Gҗ�7L�Orb�T;���۽�����?`�k_����=���W��B�3��x6���7y&�e����{������=o��s��_>\]V�{����n�>��m��׷�〭V�iY��/Q��^�?F�9�1�:���Cra�~��+f�\�i������7mÿM̪���kڲ~1��U�mg�|+j��M��>Q�gW��w����h��L���?{o<�9k|�<�i��ݷryJ�_��H�!������]zC~�V�Ge䫾__X*w�7������Zn^�95>XE�s�}�w&+�>��v���s�Z�C6.n�O��n�t��1Zml��깎� j@�i�Y����Yw���5V��:�:�#&��/�T9�����t�A 5��¶4�A��6w��δ�K��Z�l�ꯪ�q4�z��?~wy�:-~hi�-�޼]A罴�.�9B;� �uO{+�e���qK���<O ��C.`�t��5H��]K��꾻�/=��(O���}]�}O��ײy;��s'����~�ί7��B�>�ֺ��l�wQ{�	m.��w�|��~��2�̾���s��\������t��q#e�{5��<9?b�8ooc�h�9	:Ε��p-�]��Jq�_�9~�y��b!�~#���ʧ��c����e���'^.�4�l.�	�N�bJ_nP�9�D����8�;�.��xTM��z��M����X�c�]������O|����u��g��L��N���_?]�5�?CJ�ˁ����_��n�Px���̛���z�߶��j����+�V�D=ў=����6����x��(�޼�=h��]O^T��v�9:�gt�����|}Ɔ?��4�:�\z�ʔ�#M{65��9��S�r>מ���=����A�p��t��{ƅd�j�v��Us.�.�&���ٵ���N���.�B�Sͺ��GS����W�UMN��}�x͉ٞ����B�O�X��\=�]^�l�q���y;����׋۰��Z�s�Q;�U��Z�Yk$<s�d��X�h��P���[�{ӫT"�L�{.�L�Q�n}{s��a(܌f&t���.�8��縌U��9�r� 3�z%��1r��K��T�u:�|�+t�o��nxJ�
{�]��Iӽ�y	{��T�Ů�b�^��͋ܘ;@G��0W(\?�CQ�3?k���J����u4���^��k��*�7����=^�k�:�ΜLf��Z�wS���.*��_�>6|�v3�}��Yʏ�V�E�Ի~~YY�ky�����W],X��f
E3w����o�_G�W�$q�}���c�~~�8*�3��u�y �t-~O�2>�zW�ʻ���\�Foi��Ω	5�IC%љ��=w�C� y��m�"��K34��j��90��OF����^8��fN��d\����M�f�Z�.����U�#um��S��Z�J׊7:3���=�}��4a� ��n.]�K�:e�]�E���Ѐ}��W�U�[��N�<'B_�4���z��ݒ��z�|�����r��$���y�^�ۏ*��j|�7Û���T������,�>����7�ڴ�v�N��/�r����Ơ76�ܛ��W7~>]�=�ES�w��Y���o��P�O�L�ʈ�g��L����m|��r�a�oǯ�wR��P���j�Q�lwk���iv����og{�ս�AZ��կH������!��f=tbjr�3fle/�k1���������r���;6�#�M�S�bc�n���?Z�FL��|6�T��ߊ7Wl譇io�vq8rC���rm��jy?�`�7�̈����_K�9o='$N��8s���:���W����E&��u!|ף�?_��������ק�&���a��M짒I�Ve�Ȼ[����Ľ4I�R���6o�x�+���.��1v,WB"e����J�O3>���ٱ�.�m$��Wn	@�Qh���3K+�Vps8Z�5հ��V�y�/�PX���5.>�0Tp��J{b�1�;��:p��1uaR~����*��oA"��n]�~�UMټ��Tח��Ό��vi��Sk|����E��o�:�ho-�0w�_�Q��*���-��Ŕ�t�w�<�Nj�7#<��|B��V�1���8�h��]]�x��e��&�I��ErW��x����O�{��Vhػh�Ա�}�`��Z��"Ͼ�Jc��;jf����r��!pi��o���~�nW6G�N�s�"�H���{�����)o�x�5n�m{����~���i��q�_���bu����y�{�ȜoiN��Y������>э��ɞ��|�~��u&k���xǝ�ǳ͍�izg|z�h�/�o�>���MK��էn F��ڍnѥҁ�񙼝޺�2����a|=�=��o���v��'�ӾB�3Kif��Y�US')����˥�֨RN��Y�B� J=\�n�_q�6S�Mu�VT��fSUN۳ܪn��l_]O��U2���\[zop薝f��U��$�m�b�\����x���Q[0�����W+�����d�Wh���d�Z޾�͡7���ZMD��\�«���U��_I]���k�|��2�l���5)o�����tn�87��Y6p���u�
{Iq˔�]IY�Y 䎷�w|�w0�Hgo+k��Y�Ee�gR�m����Z��:欫�N��w,�Xo-5rI;�d���m�����x�:�g�hZ��Bu�a5(վW:1�.��CO[���o.j��hszl��6�S���d9�eM`��S��7[؆�$v�Mqj�:Y��8r�ZH�7�1=�*�'�Y��P	�y��A͔)4���V�k6�K���ݘY���Q|�ScZS�L�r�s�6�Q�Z3�uӲ�mӕH����I�ֳ\�[�Oٹ�*킻�ra�mso.��Nb������/�W6��fk������G��hS�
c~�j�vj'&��2��B�ko$޷vI�Fx���^Z�Э�/-�>���D(z�r'F��S.�ژ68��o9�N����:�����O-��-j�&��[V�'�k�wH��6�&Y��a�{,��gv���+���5�5Ge*��kkpV+�cc9�n��<��^�Ң��'�_N�q���,���\��};��G>��%I��}m<�p�n�E�ӄ�xU30���8������Y��U�}#�_-�^���w͋�C�wD��}V:wmԘ����gX�V�5��6�M�I�.ՕrE$��"�r}���j_G�>�ӶvQ1�K�]B�ヰe���Ѕ�4�r�9��������K������JHSn-9���&[��[��{��EE;�#�����U9˸]�Wg�c�C�r*��,vWa��Fu���o��qK�����jP��j.]��FD윃�����(Z_Ni�rģ+8;8m(��D��M���;�Xf�/���Ŕr��V
���̳P樂��x�ZNWVI]-���`��Jt������q�&[���z�;�,����ͼ���rJu2+ж-Z����ۦ[V�wM3�Nt��'�O&Vw@��s��b���װ���u�ˌV�Vʟ]!��&qW(�u(������I�:���b��m���(��L�|�1�H�*�� �tS0�+.�\��������ҋ&RIV=ۻ�;%Y�`[��,��k)�dF<0
}��J�o���w%z ��BU�E�	A؍q}+{�9ǹ�;/T!�3���v�pC����&�����������ǡ�[�-|�H�6/w�n���DB��T�ŹJy����.D��{dȪu�u&8䜢�E�S��]B�Ʌ%r�Hy"H�9fz��Rv^Aq+��r("iӧ

�*8\��\��M֑�g��y��5�^e8�WrL�ePz4�J
*���YAs2��rvET�t���k*�;������sX�nd�\I�"���\)Շ�����X��#���\p圌��ʢ�E�*�֛�w���Rʪ�((�iY�0���X�((�	�.Y9�#�Iɥp������Bn)K��UQAr�ջ"�-B&�@Y�
�r�r�*�E:��
*3ws�I���9���BtE��*8GI$���kw݉ȩ	�] G$��#�MչĪ��w��i��L��E]�W�����븐�j(���nE�DW�UQ�H���w9H�y܂-hy��4�Q��Λ;)��P��_��׬���K�l��yH�ٙ���v��w��M����n]݅p�v2�+���pV�AgX����͜���9��G�}�:�$��q����H6�CaFk���B��#/}�󹊘U'|�\�ϘT�m��M���R9)��zG�o��q�N8P��{,Ĝ��[u�`�WW{*o=a��VO��yɣ^v��mb�=��n1W��5�(�ң������'nU�i����X=�T�z]�w��q�����y9��ϭ-}���-~hi�H��޼]L{���&\�Q�v=���z�w�y^����u�ܯK�w�mo�̜Q�}�WR�.<;����T�A]>5�x�>��u]��߭{��<����U<��]&������/Z��\�o�:Q���N��l]�j����|M��^��yk�w�^��o��ߏN�9k���t�~�}�N!�Ĺd�L�3�zR�uwf��;��W����:y�O�nE0�9Z�\����z9�(�ޭ��:�0�g1�p��bl�U�y��\(A�Uk[\��,"�M��]7�խ]���'a4J���-�<!��C�YM�ڵj�V��6��q�k��bAg�v:M����j�x��+9Q���4�etL+:��t]�I7߾������-�
������Թ���-���?/f��w��~�K;�wV�nwNU�������_�S�9�	�i��m����Wf�����������r7��jŝ{���5�g>�{ϻ����1�|ћ��M�}@o���f�5��|ŝz׋~*hl��e�ʍ��K��O`��:�c�3����a���K��fb:�{��E<��{5��S��u���վ��ѵ�)OޭVw�S�Tů�v���U��Q����u8×�5tw%���y�Ƽ"li[����Y���u�r���Y��V�A�מ��6���$mB{,��$��_=��RL.V{��K�{�l�^���pt�͌B]�� ��m�Q*�2��}G�sJ������ӱjfqd5)��9�^�\O�ǖf��=֙�wS,��x2��r0f��SV�B���ox ����"��[��]�7\��FWT��ND�Ȭ[\���@�CR����N'�JveX�m-W3mC����k���K-�j�J�����Z���@�T����g+y�tP�Q�ʗ�R�/b�����^��ZQ(�K�}���R��ӷ��_�Ԯ�l��b�^t�qis��i⿡��<��1�fU8��v��&���.��nYڋ_�Sv�R��RϟP����Sk����4�|������J^&n/��EQ��N�=�.�#�Fnia�4@�Y�߃�XK��D�yj���F��{�w��ͭ����tc�l��v��^�K7�h�ׁ����{fkG�_���Ǹ��eg�a�R��XY
�H�O��ۙ=��uY�T�˝ݎ�=�+Uv:�A�~�\��J�W����*����O��\�ޚve8�ҝ�k*������7q��k�l62W�{8�Q��-ãƷ�1�/�o�=��o	��]o�Ѝk5��$�}��}�y]�t�G�����yS��o�t=c+����t1���:�C-��z�+�'N������Nk(�n:�d��^���n�0����Y�gh�oP����}��� u���#��Qt�CJ�i�Ay�u��L�4��F��ΣǤ�f]C��s} �HWV����{-�(��Lw����NK���� ��Y��1}ik��V��M�ݾ�)S�!�:&�&��Ž]+��>^4�����k\�o{2������n}}×,�o$�����'`T=b�y �׼����{``�y&^����''��V!�j5�9�1&��({$��0�=C����q�?r��?o�+�.z��.��n�0��C�����9�1%k�+#*w��Y��m�$=H�ߗy���P��K�R�u�1�HOG�tz=~��Ǫ��ڧ.��e�����-|i,[T����,����wy�Lׇ�9X&r��:z��>!o��{,�k��]�/m.��ݙө���E ���}�C��óǟ�צ�Lm�͢��S�J+'\;��y�fFhr���e�lMܶq�x�y����5So����.)ʲh���i:a?f�kt���Qfi�=<i�s�TThɼ�=��Ʒ���y8�<����L�Y�"��ؐ�<��kͅG��o�=���h!�w1��R��c#��_CW���ݡfҊ$8��ƻ�-��+���kiob��}�[)�R��֫���I���� �ˏ�p��Xvn$���x�w���M��U(k{(�o�o�wC�ً#ft[^^��
��N|����0Þ�m?}����`�C�=��ݯ��g�<��a�Ȫ3lb�w7��W���k�s�ĳ���Ϳ9W0z7����aѤ.�:�����J��x?IL�zb��{�]v/6 F�#�O���Y�^�9�o����f?A��X��يv�f&1�f1��>�ʨ���.o�b��aW�f����W�k-d�q�K�~��.����Re*��,�+<�z�fU�q��ʃO�ٿ>��n0k\c�ě�Ƴ�j��Q�v�_��%@?13!䂶�^ܳ轰T^�3�CƱ��t+B�ǣۦ�[�^�z�:����s5A����Ļ�P�F+����zN�t���ޗ���w��K�w�mm?#H�ڢ�
�����n�9�^����9x�j� j�v�o/�b��5�fW7WO���
�j���cq��ثI4�K'�w�3Ó��i�|-W�PK���ĉ'}�=��[Z�ҹ<��(�C/s�W��b�E/^R�7��,'���0r����J�W�3��Ԟ��}3�V����̌<}��y\h���7�𱳕	@O:FN��?3�ߗR��寨};|6�����/�y�,1[�	�+�JTOo_�:{[�M��jW��N��=���,�qϯ����3���1,&h?F=�==�I�+:ܕ�g��ya��nD�]��ŕ��=����K��Ęu�hLi�9偀���k�~�[�r:��S��ޒ��d�,4�~Y:�	����.֪�e��!����L�>]%f�у�>���7+
e�6���"#f��ʩuP�0q�`g�V�9��b���A��\��t��Y�'��Oa��G�b;��:oT�,T٣�_UH�>���S.������ON�G���'��9�����a�OȎ����!]�ơ��\;9�g��PS��f���3�?-�	�=���-<��ܞF����\��\:�"������.e>��ĵN잁���W�^/L�D���7pa��ς�+Hg�^4<=鐡u�P�0G��W^��(�\(O ڣV:Έ���Y�z�{��:	]@�2P���]��YYē|���wD�{�}0�ݼ�*t���+�ǻ;ָ1���-�g,�\��T��O4X��lu�iVl�KZ�t6m�5���	���C"τ�BV�J��yf� ����	�]H
�l�;Q�㞜�:�Z7����]��Q�y�j4���S��*o����v��Gr� :�&9��*�I㢒�b�9�`���?y1�LOl�	�&c0<�^��,����jG7�Ɨ�����K5f�����n��m=���/W�u��d��h�F�L���p��'1�u061w�V�ʞ��R؋>��y�N~�L)e?״�،����ꙫ�֩ڟ��\1Td��d�\�2{��t�֨#�z���dIVf�ݾ��x{�X��W�r���NL=��h��hu}��L{0��S紺U�n����9��̓�P����q֎Rs��UäE�\��Օ�5�����</��+zmN%M��s�&�{�R꒺#�1~<�g�#��t��ޒX�w#��	�ۨvO����Z�Ý����Ie歞�7��|{ZC~��f�ˇ�����"��,5���M-��yo>S[��w����p{�����ou��	��<[/�\��;�7%���t�-�;�Q�(=7B�UA�k%��	�C���5-�)�7���t;�Y=^L�7�+ P�"�,֜�gN�C�,�Յ��%�4����M�\�a3�{���]Tg�jY^��U�[�Q�v��t���F�Ҫ˼��9Vt5r���\�Ծd�,ֵh�Cke��4	l;|ӛ{�5�����.eU�gj-P�1���٩���pet�G
�ٛ�K�ќj�~��;��(f�ؑ;�]���*�o�+�ᢓY����$�� ��ڒ���x���AX���GG�欐<��J�u� 5�Yj��<�����ҡ������p�.���m����>&����\t\-�\�3�S�@�7f�'l�Q�!y�S���z�X�]m,=�/KF�s��>�!M.D{fHzj#�N��NI
Z�2(�$z	�懶s"��tg�,7����1��ΨF���]��� L>�D
�`���
��������L�A���o���f�hb7�ß/��F�%��:ba�ʢ6T��w0��2��_�w�A��Da��[�ӫ����3v�*�ژ�����YV���j��F�Y�=ﻦGq�m�K����뀮)�^�~��{�3��3��c��ϽP�=s>5��⬖ �˅ƥ|D�2�c:Sv�!=��zzA���Gz�G0���#<j�"�ӕc���^.��p.��(1�j����=��'c+/�S��$�	4t�W9�:���9iu�y�U�-�Y�8-ݫ{���5V�ae��췙Ux�'[�����y�p��OzX�n���ޮ���p��a⏰N�R���X��1~�~�?>^z3��h��=�a�Z#p�V3��e��Q����B��n��_�37W�+A{��=�C��j��c=�+|��N�k�>o�"���{����z=�|v��B�~4Na}���H׉��N�Q�W��ϴ��șd\M�5��y&@�W��Rit�'(��-�d���45���G���nu��f�C5=
�I�N���vf��F�׈-E�}ж��M:�&�k5i0�����a��7��EG�9>���G{tj<���]Z/�����mTL��iH��;�u�Yj�Q�\�q�Nȝ�;ү���5uR��1��=九��pl(��t��h���!�Q�Y�����P:΅3H�ڮu�������3k<y��t��<]}}t@��:0�\�}��L�{�ƀ���9���	�c���w �s����g)(�5�Pg�y�mAR�� VHM�Y|E�o��$��ǟ�
��K����FsO�<'����|�MCyT-\�w]�y..�jVUǈ�Z���|M�5{̋'�4.eL�4&���H�n��1�.��龫ZpM׃:�ަ�ܯ��Z��ԉ���XQ\KU;G��$R�+�Z���`�������G}ܔ++��)�#!�nev�!���	����H�.�l�譚�l��d2˛��Z��:�
����fc�r�ǽ&���
�;$���W�&��?ݩ��~"���M�1����d��1�e���� ���nٿ�����C�Ƿ{^���Rx��Q��ߪǮy�~%O�ک`H�4
z�(n���{�y�3�g���a�hWm�AO���jrxa�M�fիqJk_�f_9^����޽��P��cS� [7�~�uWԤz#��'<n�=K��z��/��î���"Wm'�^�k[/R�'O}ڇ�``z6]@������ʣ��:k�w��W;�<��{�Wd;UB��f�f�k"�ޚgEǭe2���;Ւ��u<}�=�ު8��AM�~�F�=�G��_�W�1�������U����V�����u(1�Κ�e��P}��T�����ƨK�n������j;$KT���o���������o%��\{���@����I�~wx�}r�����`�z�;ْ��x�uh�mT	��Ղ�;�ʑ�L�YZ&k;θ���U	��i�m<5k��ƫ��[�!Ѩ<����H�Nl���������%u�V\u�j/v�Z(̒��|�g��1��jk�t�/:k�)� ������44�u�A&Ƽ�z<�-l����Gjݑt��V���f����J���Ș�C��s��QW%�
�vY�������E#���lKBܧv9.2n��l=���=�l�s�Z˩�U82�����J9��bf�J1�����(��"�­vm-��)���G!$�ǵ���$k��mZ�T+�]K2N��h�k�&h1$<�Mluc�nj\$��bݚ~�lXQ=%���:�=��u+�w��v��+wz���X���)��(]d��%_���rr�0��h������X}X��:�kH��6Iͮ��v#X��X%5�biJ�V*�[��++0/r���op�6�$���x�t�2S�
�L��A��*���rH�����(P�L���uCz2KY��:o2P�\���L�p,C�U��Z-\0�9fQ�jX�^j�Gp�n'�i�}���欶�~���ɴ�HK�3��Y�W@��i�޼�}���vW)k��j����7݆Ib���s�����-�M��� ������0�����v�	i�ǚ��}�ں���/2���̏r�P����_�#�'I��D	عMv�R�д�O�v�Ǆ]��Y�A�$nr�ڭL���� �2�m+��A.�3K~��v�An��#���v�m���z�(ߘ&����1U1:4ץ��ų�Z�xδ�g�"G�\П1���> ��
$־x..�@|�u[b�^)��j�y�)SO0�]�H���ff[�q��j<s]��Ztq�����P7a�3��&ûɬq���LS��j���F���8Q��^_Hf�Di�������[�M�JH�dK�;�t��[֗���;��t��T����p��x��$A�컾4x��N���΢�[��9�KR9�
��%�Wb�	.U�t���b��HP엱s��������S�^��9�FU+�5U�΁�\��:w�&�4-^ZB�.���%����/�gq�sx������2͌T��J�52�%�\�Φ]������&+R����+����3��1]��=`
���v�n�\�SK����ޅ��_�N�q+��	7�TDoàe��t�t2V1�k�>�If�;+���j��ڷw�n�����a����է�� ��ǜ��.��)�E��{ܕBw��+lfL<l�F���8�����y�$i����]�SJ�.����"�=��+d���dwe�h���]��ǃ��<m�p�z���A��{VV?5�e�V	+�R��V���+�*.1�k�Lau�Vk�6ާ'R;%$���wR��#�6����%4�v����=�-k���k���<NN�}���a1����j�3��4}�rq�k��Yw!��8��t��s�8UQr�)�p)�]�؜�9ՅJ2�+��$]�����BQ	��� ��{D�9$N����9^I0�*��h��RqT�Ȍ���ݖG�N!r��[�y]8����;�Ց4�-�vRt�VNNQRpN'i
=�V�#�'m5e�J��ʒ�`]�$T
靳�-
��L��;��=w4��ҵ֞N�dY N;���Խ��Γ����H���J��8QTT$�&Q��a9Nq	2(���s��bLH��.��v�9G(I��t��
�9	�sg��
��q �(HH��;N�rn���H�RD��G(�(/<�wpstp컜�0��"�$�.�ww�ɤ�:L�$
�\�qp9��̃��w�������cu6��L��>Ii�x��b���KN�if�_��,�dw�g0�G�%῞#�1�]Qײ��=`�fy��y7�a[hgX�^{�=B��2��]�d�z|4�Ã#�a�_?":k��!]�ơ��\U3jo�f<�͡]�|"�u��>e���xT.������,g�˙|f���@��T�G�}��r���D���-�$�*��Q�N�|K�w>���,�����p&ߦ��;|���-v)��#{�Ӯ����o�ӒGO�Sh���@ti�t�F��4E��E����2k���B�L���UFԞ:*!)�.�畃�o
�}���W�J����R僧����ԋQ?>�x�9�p�	��2��3�?��u�6s`? ={�Ľ��f�p�b=��1�`(����Z����ﯺht�]P���e���=�ţ�W��5й�o�Ua�tU�����@轚d
�\�Ou�I0���~�g1U�7<�O�h����=�p�|{&Gz��߽;Ǵ}�< ���@Q�W�OE�4A�z�H�G�F�fDq*�ߐu��&�.�8"�L��wV�m��2��"��$S�7����k�����7��c��P&��.�*�����o��{��ʄ�>����ȧd1�՚5��wM�)�gy�h�hunRe޼��Z���n�Z�s�u.���d�кp��!?�v���7��~�{.*ΟV�v�0�i{�G����</_�,/����N��Uk�۩�;�'���Q\[����t��������V�{u�/5
dˁ�)M�U[��|�#�ѝT4v��:[�T��ϡ�v��%�N�CW��XZuB�ɒ������6'��W�����.�Pn���,W����;�va֛��;�𞢒h�p��l�]9V�'D	��oV�;V�h�ܜ�ON\<��=��.{��e�'F�eff���#�����R,Rw Oթ�Uj7&�g0�ܜ�s%�Ȟ�������[�d�:2�ׅ�ə��h�^$��:��Wˮ��RϭC�^�5K�+�.��L�}C�غ�M���]oQ�I�h��x�����L��ڣ�Vj�!�t���~����osۻ�ܬ����O*��ţ:�u�}=�I�l�w"rH���d P��>����w�H�ё��a�E�
���y�[+�u�y�� ��=���h�r��h�Q��
�4�]d=�H[�v��e ��ү/w������Q�K��rw�֒����x��Gq.���v��*կ-ߕ.7O�U�r]�F�=�����r�ݓZ��c����/d�z�T������G�xt�d���X��:b^t��A�����@�O9��D)��s�z�rO!�̔uTQ�Pv}�q��ư>�8N�O$�<��2�����:,��޴o�nuߞ��2�\Ш�ve<���,��9�����|k��FK j�ëv��蝮z��s��5-G;�G���wq���	X~4�I]�ˇq����f���5����5{�}0=�Gz@QګH����5���n�xS�I�܅c�pꈹ�����-�'�f�{dO��nl'��ڇ�`!ߣ@����K�ծ�ˍ��x�:�.����v4j}�]&%E���߰Oغ���3괽��H~���Bc^�
���5��eG��Q�+t�5F6sx�ە1ޓм��[3@z)m���d���d�l�5Bo�p�ih{�/���qX��r{z2��j<���h�W�:ó��:�&�k5i0��R����~�8�|�n��.��/ؘ����q���y�A��x�6����OԵ�Uj���N%�SVhd�u��}��i�!Ҏڒ�����-�oT�[�↕YՄ�Wkp�FǪ��8.�~�@>����:�j�֗E�h�y�N�讹ɽ��0+gn��pƸ;�Ð�W��t��(�d��d�h5қ�ڱ���U�B�B�"�m�E�[{�5K4ߋì�͉s���M�D6j=���$_�9�]Z���5ƨՋ�X-���ߏE{������'K�x�_]1Ne������P�<�lf����ڙ��X�{l-^�/��b���k���,�B^�QPZ㊾�s�u����jy+�E��.����C��}����������Yˆe�����<+��q��2���ۛ�7���Ly���jnM�n�P99���~�u5Sh���Y,xO�l���#'�?9N�B��9���S#4�hDs��|�O�P�77�~��p{	YX�ߍ��d,��J�@���ج���2���|���B��()�<S��-z��ߗ���4w���8�]m�0�O���鍿��d
�#�o�x*}�Xx��Q���v��m݅�8}|٩����b|}�[YX
����������)Gz����,�o�����E�W�U��x���Us����YF��u��z�%���
�w��P_g�V�w8~̔�����-n�dV����>&��8��3�xͧՐ�h8Çc�N9Ltk[1�2��x]�P���unT�]v,�?]>w�U�Յ��@+��c}�)�`�N�붇E�ťԑ�7k6F��6�\�˺����,�n���ųD��)E3�T����^r���/�k�'zf}{R�E��5�u(1��#ׯi�:�&uѪ���;[״{Fw��Z�Flw�gM-V��:j,	���Qek6O��X���܎k�׵�6�ũcҏ`Ѹ}n�kk���lvH�L哩]�ݫG?w�k�w]�(ϬE��<m��F�}8���,���5�"j6��w ������Q�j�6�J}��~�5�F�iaW֟�T�l��nK�<G�{��:�M�"ş��A�k�\�dq31�[�Y�JL��کP��B���
�֌���m$�����dqR���
��U�$>^_D����"���B{����eD�H�P�M
�w�>�X����A��q�������>�O�w�S����O�嚁[�y��$�+���'�`~2o�W���?�O���(��p����$]�2�{�@]]j��.GL��;�(Q>�F~��{
yW3)�oI9~���Rz:B���$�l��sg���;��&�jO	L�w�+yM�����p˸��@B� 0x�%Z��"����0n
�)��z�pm�eۥAb�c�J����e޷��k��i�c8
��Vk�l2�ڴ&`���{�8-\�fD���5�D=b/ɏ��|X���,Z�Q۽�ջϷ��/^�H+w�+����=�خ��Z6�"v��Nmf�������S�x��AC�ԏ(�Џ�:����H�[(S��C9��g�F��<�7<���`���x�Ǖ���ư?G����8i@Ȇ���<gz�_�;�$�U"%F�<��"�C�3��1מSxX����5�&��,�?g\����W��&�����4���߲�ɽVjw����H3���w�*�{Ӵk� {/m�����q����W�F����rϻ�a	��^�=�Dg�����Z�y �b�@�Ln˹�Ls�{�ϴ۫ݚ�����@]�K*�j/K{��=�������]X0虠+ra�I�B�`�_)�]��ڭ�؞����竾:�:�Oѧ��+�Kx�l�Tz��;؀L�w,5Ujd���\��I!����[��9$~�^�X�i��A�LH�[s�7ܬ5�u�$�-������D��7����{�� n_����]D	�[�Yl�ڡ�cq`�����"����=��ط��ےjs��:&���mG�8�wWA�;/j�X.���Vcs"*}㠳�L}�x�;�>��e^g�j�p�Q��i\�(;��X��[I���K.�@��I�*�ؘa�:R*2r��׻6-��y6]�u�a�Ww�W�V���X��NY�bw����뛛WLo9%����jv-��8�%�w}��Y�O8���s���?n���HTGt�v<�j���IB����,�P��
k'�&��}���.�}-/�E��:,w������s-��7�(Z�\z�M9�W�����}y3~�d���Y�}�P�3��|Z4��ޤ)�ȏl�O[��w��}>A: �v�m� �ՙ������Q�tyj��� �����y�� tW�6pS5�uU�`�:��T�;��װ��X�f=�æ�'��T����LK�7�Fʑ���q�]M���G��x+�ѾH���ڨ��wgf�a߽=���W�=�S�u$�1�y�w4f$:p����O]7�����z^�_{Y�0�zٮg1,z|� S�l帹��vT�{4UOX�J�h,�_\�4��c�'gL��4�I]�ˇq�����a7n�{�g�N�^�n�7W����@1<E���Q{㩎�X.0}A_q�-s��u���*��s�+�b^x���5h{�:���-Oy!L����u��_o���)Etd�q��*�� �
���fR8�ޞ ����������,W2��qWD��تJ�9�6\�t�hAo`����t�vq�+��Owr�w>Sg4�e�W60�Ih�;�F�U����V',�����4�c��1.�]Y�K��(mk����{�����r�@{�HE��^�¾�K�l����H<��'|��H�8�^\nTm)Ȝ1{S�6)g����1���V�)��:�@��X����,old�l��(U��9�A���h���3��?��S>;�VF_tL�_Bi���[Qp&�H�r�j�a鿣)F�e��\��"z�3d��y2�V�Ύ�ႡoO
��tY�@#Z�]:�嵐S�~�u�V���������K�쭝�.��1�9���p��t/	��LO%ĽD6k�3�)����J���{'_� ��p.΅G|f�Fr����a:u�<zīM��3̧s[�fw����f�aCC=� {��lP��,�w ����pq>Z�Ů8�Z���P}:�g*�]\[
�[�b}�h��!s5�P�<��P��ܚƸfAb����;�:h��-~�}U�Ub�G�ٻ������_Z5`�����7���}6��~=5,xLl���dc|v󢳰*~�۞4{�@<e ��h�9�R
�Ԟ;_@JGY�ٿT;��#?x��v��w4����Z�Yi0�/ qo��^��}�.���G��fաX/Y����Ԭ�x���q\~<�?1�w��v���No'c�n޹�W;�+7R��e��$4�OZ0�eh��W�>4�;����j���e*Sz��
�����2z:�|4��͠}3î��]����xn.P������LeuʇX���pt�;�c�
V4�uQ�[ T>G��}3�>��������{}{ӿN[�˟W+�eD�[u�۳��}�L�.��O�}�=ʣS��.�P+f_�_R�S}�b7�q�W��������}(��uD\�����m�-��;ؘ\�	Ʈ��ή�����똢%2ene���\���KT?xN�׼N۪�fojX���Ư����3��`YO;L�o�yT��lz�:]ތ��N���%��Նv㦢�����+Y�K���ǳ޾1�zU�̷7|��;*�ӗ[u�������h��� K���\N�b��u�}�n5]N�N{��N!�;u^R�x�G��9�p�xi�up��rYǈ�'`�L��/;��خ&���ѓ�+�W4��e�g}�A��k}O��+����#�G��!��b�t	�]y�K�tx�H�2���ώ�Ъ֌�/�I��Qܰ�~Dw�ܴ-W�A���5�V���3=���iN�9�~U�p�L�d��^�V���d���a�e�͝�AU�q�W*��0�=�^fP���C���'3\���Ml�-�,���W��*=��b���T��K_U����e����W���P;��&;�g �,.=U#��R,��wp�1�0�P�'�8���kb�?P�^�W���g�O��ڂ'�3��*�@ob��B�O��Q/���;7�~>��ǨvM��s#�t_��t5���Qޠ&)�R ��@�Cx�rH銩�{n}ݣ�$m�\�n�nt��{�v����6i�� �ΐ:�\�/ˑR�O��{w�ʫ#�c`�z�eesў�
|�x�><;PP���1�#�q������R�C�gTd��ճjI�����I�}2�G���܏+��9`+Ɂd�G
ݒ��S�wM�1��Sg��~��y����yB��g����q�7��QV}�b���R��s�^�g´q������I7�y7sA���~��d'����ͯs{��y�=��O =�������ٺh�:;ʸ��|^63�ưm���Lak�|.צ����]��p�f�w\:Ǜ|�m�'��쀣Z�U|�b�����	��4����|\�x�����v3�#��v2�`�/;��\���J�u��o{�S�˻r6�TwW!�8G�Sh��v���\�g��K}�ړ�:�cg����]���f}�2u�Fs"�J�[Z%q��xq�`!]J���.���n���>P"U>���ʇRz��'W��A(u 0��b��nP��)Iܳ:;�
�o�me�)k�̦���v���{��ݚ��*�ݕ8�O��1;w��r���>e��N�b��n�<1�ɍO����+��������ǵ���m8���}u(A�v��@�+j��Z"͛�°&>"��.�Bd�S%2�:�P�9��z�� _n쩂�)P��]R�֩ z�;�����o)�_U��y��MFaԹa9�;���`�`�E���χ�T�a�쥉t����Î!QY���.S��5e;�l�qD��BVE�I�x��_q��*b�L@r������v`�/�e�1�b��Pe�[Γ.��c]�u.r���J�5l�9�A!�K���X"��sdT�8L���hEria��Ž�3���
cs�0�֎TRv����G�P�%.��z���Q���.Y�6�l�&�YH��<v�
&�s��t4�F&��i�Su靕�^��JF1�����F�Ԑ�[\U-
��a�f���[�2Jt�hiW9���ǨiJ�ZBmv>���&
���3���?m-X#<����@�P�v�t��X��������Ž]2�X� ]^�ﲯ�r4�]�1��wUٵ���KG��S��3I8:D0���7vV�����-��<ެ���5�|[ޫ*�
7�{kQ�Ά�EW,н�vJ4�H�h-�hR��Rn�Wi('�/�B��
�X���@��搛ܘ�n��O��IM�]M��w��I��V�
�6��^��>�)0���^���b�%��R��BD�;�K@����xA��2����µf09Vva7[��Y�N�_Su�xJ��o-'�\�5-��F��5�,|��Ϊb*b0��ma��Wy/�[Wc7F��6��PK���{R1��N����u���.�CY�djf�,kNs�N{��2�]��7R^L��[�4(>OJuʹ�ھ�)�/+��w�U���qp��
W��һ��9{OFh��N��W�1�4V̺�94�U���]�q9r٘�>p�x�f5�rmٵ��L�n}k2�õn�6���,E��g�ޑvo��Qg�w�[s�K��5Z@{8�y����+�gnf[���b��X׶�Y��$���H�Y�E\�ӁU��U�;���X3.�i�Rʝ�Ҭ������;�L��ƺ�o)�֊5��{��r`�F�"��� ��Q4�rsf�<�z�K9ʪ����]�����C�8��0��ptvwJĻfɎ��i>��^N�z�^>y>y��ǔTIޞMΝ!̆DQC�Ny�;wAÔSN�ʼ��2�99B{���^s͂Wbq�9�8��ŕ�(s�9ӕj^I	4�I&�gi���)$���a{�S�-6�Y'.mu���*ܔ��@����9��X�"!-O!Ֆw:�t���I�w�NdI�EU$+�Ws�l�^wt��$�f��S��p���gg*���T�"��I�ҹAn�:�++��9�Xu��#�MbLE.P;���A�:�$����Q]ԇ/\�B�u
#�P�M���������.�9'K��\:t�眸�#&� ���'��*���Z�˗���w!�2H��$��E9�G%J(J"�L0�.$Yn$�����T�� �4n���r�qK�	���͠L��)�,��r����-ve%g^B';Lmr:�|=�͊�Z\�TZ[���(7�2=����<q�ڌ���9]�+H��~���GQ��zFv�ƕ�J��`�-�&)n�i==q��u��	��<o���Nkj���%�g��H�;�E{�1�~��oo	�5����j���u�x�>��6���S��	��k1g!C|=�l/Fw����ڌ3c��̚�p;�2�	�� V��e�ܥ����4�׌ϗ��zO&y�cz㲈𘮧HWt�wȶ����R���2.	שK~mw��E1Ib[���ٱ��8z;2a�-dq�}�����NY#WJ����on������0�vUY����&{C�wٲz̷�K�:j �ţP��ޤ&)��"�ْ��b��trT*&L�AZ�7�G�oV��!DN��"���ˀX��cN��]#y\#�:Gl�s �{T�'��O�"�a�cn��x:���#1�:k'��#T���1?>Cy$�7�=�&$��m���;�k��P�%!o#ڨ���;7��ޞ�Q�`*~�K'�'Z�?�����~��ʧˏ�����fv����D��Z͚�;(�Z6�����20��E��bQ��q��>Cv!ɫݦ���ma�QtG'B�C{��q�`�u��(
���#v�r����Ҋ;.N��y(������g�i�z*fR���ׁ��g˽�o��iH���()�'O��*;���a�gƾ�|qgqU>�DE��3������onW��5�Lj`񘾹h�w��sẎ�#<j�"�ӕP��Snu�f�x��ѧ�����=1�ʸ����=��;�Ň�h���aX�����:Z_�#0��.^~��3->+����g��,u�i�$:y�^륅`\�Ժ�qsG�}[�����nՃ�2Eu��¾�K�ե�]�A�d�S	��Ng<�<�ae{�X]�oн��6�"e�M^����
;E�E���E�����l�B��g�}�k��f���Tux�vK���5Xu�֦�-mE���u Mr�j�a����X��S��W^�w��2�Y�rcr�Θ�_t�W�W%�cȶ���(Qu0/�fE�'�T��r�ޅ�z�}�7��z�;�a�K|{����5���ah��D6k�g)S�^��m��k=��+�\ت���U��1�Lm|�/q�'M?#��T��2�н�k�����~�z�,UX�1n��[�g��T��]ѝ��~O��W))mZ��w�.�T��O/V�C���59(C�G�c�{��y�&(��{q[��q"��-}[D&�\�yF�^.w|�A[���ٵ��N��2���L9s�"�mbNtq�e��R����l�?;TYf�k9ذu|�r��g�):�{��2�^m�S5����mĸ1�Ή K��񃃷=T(�Srk�k�d+ڸ��S�p�3���	����ӱ�'F��_oz�	��q�dv�R�w��Dt�M�?i~=8���n�
��1K֍��olx����1ݲu(w��z��=('=(��2:�9����Gb��}9��]6����sD�Q�=U:*5"����/�xu���E ��9�𕋇���ƪS���:N]����c}iY�Ɣ�h=Q��[ =�7�x.�#��O�ֹ������d����k�'�WB�Z=q��=q�b|k��1*���[.�N.�P+S�.�QӺ:.�g�];�vfo���6�;���^��������k=0~�M� ����C�Y, �]O{k	W�&�:��e��z���Lz��9�-r���u}������Z��Υ�+FM��1��=�B��;B=c����W��6:��u����tm��-T&�3��(}{u���K�ނ�t4P��3s�]^�
��ɪ�ӓ�c��>�P�>(B{�c�\[�I�/۱����싹�klaw�F�,ꢔ�z�D� d�:��k3�ns�᫰��1]4F�[�`��Ѕ�e�eg"�4��";���g'��on�K3�����sBt���ֆ)�mxM�9�vm=ep�.�E�ķ�D �v�D5�nV���:3Ӹk�(or���F:�?Y|sŲ�u�up��rYˇ�C��0=��R=��~�yK9��N��?=�\��@M-�«M���Tj�1�nK����uuGg��M���n�Ey�6ǂ�h�:�"'Г�5�
��o����^��#&�*Ǫ�O���2gz6����*O�����<���#	ܵv�1�0�+������e��w������ւ��޾��Q�1NY����j��خ=P���;�K�w��^�5�u�y�T=�Fo����3����˃U�)��>� f)�&�gk�ʆq�D��W�J7�\}���E�|s��u��9�㫐��y��������O���WyNd��^�`���V���>Oģ��{dL9͙<���7�q���� ����o����>�����/��gxE�������b}9`+Ɂq��*50'����[��l}�?K��F��)�[�wnPR����q��-�)�V����|�L~��N����3o��&�r΀*�v���N̳wj1��r�s,�q��+�5�Z��(���v�YYQa��m�&<b#-ٶ6u�ӥf�`�lGB�2�,tq%;�K���i]����݃��]����Ǩ�6�-�%���i�N���X1�2�q��|��s��yP�֨z9؜�\����\�aݬ��y�=�9i�lq��eoTս�� {�;��:U��;P�l!1n��Tn�N�N|<u\:D\��������w�][Y�g�w���%�՝ +�:��QZs��i��GL��!�ՋQË�e�ؘ��vlV����}�2-9�p��U	�����ʏ\7�<v��^��/�{�_<�Ϳ�c?�[��o���.�8�q�V���d7��LX��Y�������	�˹מ�^�{J�8S��U�6�t�/d�'j����Zw����20?�rp\���TM%��W�=G��<�z���cb��L�p;.6�E��q��Vcp<�ݥ�}�6�J��}Thr��x������]]Hz931�.�=VH��(o���Tn��<�L����/0y�%��{׽0ϗq����F�#���)�з]�G��b�x4�z������A�D:��X�P_iV櫡m����>|V������f�9��m�8��s]�	u�:_uEAK��pÃ��嫶��nn��r��u���ڮ��K
B�'�֫j�v=&$�y�WR��JB�4.���E[�����'6�q���7�_E�ت�}����e�LuB�Κ>O�E�@=��HQ=�I�"''�/���M�t.��Z��gr% a5�2*7�a�ٝ���.�Q_CyTF��3�=��J��Ws�*+�9���'�=�<H	��5L�]�u{\yX�g�xt�OLj�X��������j���e@���׷�yt<���ýP��(orGPF:�����w�F5����� ��9�*��1�{<�;�=cĝ#�d���dw��hWm�AO����}ӕ�q����+4}��rg�ǔ�����9�;o�]s����R�"����7�<�>�خ�2t��+�_'�E�s���/�%���΍�7�t_}����W�\Lk��"���5�˘V�W��{�#0�F>�L��(��+GX�������Qi{�Ty��0�>�sF����{�TGu�{�gw�!�~��������9I�6N���+~��gd�贼�E��]�A�.=�e������ĺ��3�+/B��c��ۋn��~���j�j㪬	��X��-f�&7�2h6^��:$/U%u\�մ���ov��]�����4x���|�g�Wy��ʗu��j�7Q��{*L�!�wl�}c.�ή�W�ht�[��M�<xQ�rP�gVQR����%]���ج�v���	���Nråc�v���%F��]�Jj[���kz����OO��P����b�Ձ�e�H��4�y�b�z���r�shC�˪R�מ���'�nOX�=�u�:�Y�oWˏm1����ِ˨��[U���_�JE�t9�䩳��{{�_@��O���Q����9�:s���.=м+���+�Eǉ�`CҖP��p{�^L�	W���]�����Y���o/Oac��.��n�����*2@�������㕙ԏ�A������T��ءGVY�vN'�Tx��L�wO73��Q�YwK�ݶWX��E5<���OMr�����@B�]M��{���,]��x{��c�Ҷ�-�V����mv��Gu�Nx�|���_BS1���u?ET�:�Nz��l�l���d���k�BG}���FL��ި�2;�v�<�H��<v	C�꫘qX��R;ܭ�:ufVjYԋ�WG�3���S·fW�@{��\'>{4;h���<��@z��Z�f�>��������%�`,�����qq�<>�XϣV}��[�Ti[g�b������R�&��!-	��v�9b`y�l罫�H�������/��wӛJ��o~7�\{�sm���s�U�ua�0i�wuR��4z�wN��pcV�#��L`��ę�Y���u�fee��-������-�X]M\�W��ۢ�f���ᒗl�3�^�X�2/�Da`+�w t��ݖ�b����C��jj�7B.3��g��WP^@������"���֩�������5�FK g��V@�Q4��������Wg1~�V�舂�7{�w��h �S�K�k�@k�_���{z����gl�����
�&����a\�s_�C�F�̡Z����MF�7�Pߌ��s�1VǦ��\��%��p��H��>�������v�9������/i�Y��C��x��co�
���[�U����0ߜ�w���F4��Bޞ�7E�ٱE�����ڿOc��;#���*b�in�
��gj�?f�a��nK�o�_r��Jn􄯽&��������p.�0;<�).���D=�c&�	�·w�g��߻�o�2�=Ho��]q��q�uf��7*�`.���I^u����A����W5��wWo��g-x�u�:���M9f�o#�o�{�_��P
��v��M<`ּN��:�l���T:�ۢr:c��ֹVU@��+Z� �}�qn�f)R�$H�b��Oy�V\���b�ox}4�6�D�s3��}\�!���ݲ�gp�r_q�Gc(My]�v��2aM`�ڦ�/&e���,���~�S�3���< ���?u��@i�Gæho��9Aplo�sig}��3s��]��d(s�d��x�l��܁1Χ�Q��g�B��sHu	[IOu8x~����J��e�a���x�3�9ԏ(�}��3û��g:���� ���'Ɔ�A�l,���3��+��g�����CP
�{u���mޔc26͟4Q�==�v"�|L��N����x�������y��0#ʷۓ%�
k�0w�����,
�2�uʇ"�UG;�6�>.m�a�*ox��S��U��:�q�u�z�ӕ�~<�l��h�Z�)���)�VF��ˈN|<u\:D\�(�T$�v�}y�w���x�</9��k*����.��z�i~�C~�8>���M����ϝ�{j�	�u��(�{�:w���֐��-�Q�MeG��zޙE�m�����ѿqg^���u�-�N�K��d�=���u��	��<TJȿ�`+Y�P���:o����:Yw�ڨ��8�T��vԮ�߫����i�X��XM�s��΍��r� ����m@�N�g�=�+���^�k!�vb�L
S1ًsp��O�\5������*��eŕ���̊�{d�٥>���rY���z�An@x�h	.HZ�����ڏzlh]��T��,��ʏoJZ��;����@������+Q�ȶ���U"�'r֧�z����[6���ў�^��+�0�k;��#�~��H
��<Kk#���)��r��;���ҥ�wm�p|��rVa���L:�O+���X�T8<���Z"������j��s�<5*��.�_�m�*:p��ڐ=1�dت��쁴_yGK%�h�9�i����Y�[�OX�U����v��#��j�Y�}9$(��̊�Z�9p1��P�-Q0s�U�RGۖ�5~�n��]j@��Ȁva�S0�����=~V1�^5<=��u���ִz27��t�P���CqS�!��� �$�.>�G�QS1�pvo����k�R��4�	��A<��W���uT�kIi�����n�
_1DU|���,��9����+g�ß���#~g�+z�{��U��e�
�R�"�S����#O�6+�G��2Fx��:�����K�s~����i�o�Tk����yr@����P�� �d�ِ���qT� &(���ݓ����Zzv�ڽ�o�֮��e�f`�o^c(����t.����Xؤ�5��7���3����Ֆ�p�V�8���#�Q⡥�*�Lp4�2[Y�t1>�\ޛÆč,M����V�F�a�u��Dᱺ��o{-�n4V�'�ٶ^>�I�w�-�G]~��p�4�DYs{���\N�A�ʝCk\���|l�w��Ui*���ȳ+5z���t�8�S����l�?G��-�(5�kjl'�9���{&dX������>R�աQ���:����u憱�V<��׾#�ƈJ صy��&X���z��ΡYR���=]Ώ]>�����omŐ,J��|V�]G)��;,W#�����
M����2S6�p��34M]W(0tB�a�Αe=WN�2��z�9v�o��;�v��,^��Ӳ/�z��R�^*���;�M}�+ �V�Hu9ڍ+j�G]KDʇI�H��n�[ƪ�.�:Nĺꜱ�j��g4[Je����J�*�nT����{���+��*CD��V�Ym>sV;�k%_X�#B��v��nt�M`�!0i�zjܶ���L�^�&H���VX_6z�c_V�&��[+���-�QI�G^��Y�p��|j̜��g
�L�v6�::����d��-��WO틣�*�&c��K�؍*we<�;L�iV�bq���v���RP��N�+C9Yb�=�_lwS�Ô�.�`q�k
�ۈ�f���V��.�v(�.B3_e��W�Y�ot��"�@���-㥱�I(��w2Ҧ��Q���p�aw -��x���.�7�|����S����@Fe����y����ĩB�K��0D��	N=X��Gc�C[%oL.b���3��6�Ng�Iͼ��o(r��i��#����.K�]�|�y�w}c���KY�$ k��a�i|�M4���_�{j��oe��ˁ�˕�i�Ed��`#3��v lqT�+��nJ����i�*V����`]�٦�;y�yru�F�0m�QL�*U�d�e}n��8�d�%��xR�יn�����o+Rn�.�\7܉��E�F��]M�����t�]�;
��c�L���k�nW0텒t�"�z���(����-fڦZ����"��Wk+7;OH2q=٣UbqZ+9��e�U��hV-�)����Dr����ȯR�;�fz�gW}ó�<���i�S+��ov��(N|�W=}��|.�����'/^����>x>\�8h��$�VD�;�x�N�=R�ڨm����3�u��U	:VE���s<���AR��p�"4�1=ܨ.�yYV��d99zAr�H�.j\�MN�����XU����E�r����TI���*��/2��"�)��N�p�9�T�����iz$uܫĵ��E�EbiJ��`z�fn��3:��bI#3Ze���)]�r��C".RV���3�:^��a�qi9�w74�S�ҳ(�t25����t)ʜ;��.^{��9�څE��.�'��T��K\�UįV����#�/7R�0�B֮�����D���r55	Zfy�ʴOt������~�����}�����-v\Un����%	G���Vo!x�J�冹H�36;�6��'m
�}$���!�:�X�Ѓ�q���_�+��������X\k@\F� ����ྨr��#�b���[�����Sˣ^ �]���y�n�[K��0�������
��@Q��$*�5)ro���3�~�[)�[R�y�x��.����"���b��9���]�$b�!����@��׼�OP]��Xi��F=GL{^dUi���Z��b��b��KY���޽�]:$x�h�~�!��9�g��*�}q�:�9���ƫ�/�D�P�`<�٨��;�+�x�mo��L�v�,姣���7��g�l��jcr�Θ��zxg�f�� �����Z�et�xVz6��k��{�W+�@�^�J�7�~�P�:sDx��~�^�匎W<�A�-`��>���|����mqg��×�2=I͊���T_��{�P�/G�t�C�<^�C��[,��C��|���vN���.��"캠2i͊VY���`�mj��T��.㌯i�l�U^�Iٚ�f�a�_z��SSȁ[!=5�(Z;/�@B�u7&�����-ɗ�s,r	�(T:z{ؔ�N��o����+�-.�P>�S%�o�n��[x.2��s��m彫���~�n6��2��ڏn�Q��ݞzf鍞t��=pQ8�[��� a�|8K������y)Who�:���-f�������v�.��n�ȮG�j)ş���̀�6��G����n �uƠC�d%�Q���#���Ź�),4���U5�#�wz����c�����2��Q�dw/��:�AWΤ�ڈ	H�&6޸;jj��}�5�ys��x��S��;U,V�x���??uW�@�ۥ ����ʾ�UؼO��ni�]��`�^���/O�x����1^Ψ��a�<f�e���z�C�]��M�oQ�v��K�_9�vW_ޙ�.������|�0�l��1���ѭ�ӑ��5s����ty���}��+��7�	_����<�?\���m�Q��{���]U^�(���\�������w���" �\��@��c`r��A�{)�E��:G1��v�dZ����ۖ֢</��Н{,*u6:����ѯMd&�i��:j,��\jܙ���-W��E�@��4���3X�#q]^Ά)n͊��,��%��d{��u%��j���7�	�ӊ�����4�yW�Po�I��1�	��獶�s]\|�	�����G��eJ`ݮ�B�ߟ������.�b�8#�WX����j�:+���n� �o�Y�A�ۢ]n�hYYLM�y��0��	���H]��ݺ��:uےP�!�.�;���5IPry9:�\�f����Qj�­�q�ý���\��/���3��.�74��w#$�r˝�_'4��Ql��ޛNa�;r�v�;P+zT���^�z	.��>��Qb����9��T��I١Pu΅V�eyxl�����mɪW�9�X���*���]N�
���P� �;��Z\z�G�'sB���w����n<y<�Y-g�c}�gvN�KG��́��}u��p�Gr�H�^�1y1�	�{�iex��sX��'4��Q�[���t�x5�p>�N�Pْ���|겦n�ʮ�8�b|}�K�:j�ќ=��n	vf#d(s�&LǷ�Ʒ�?�;�ω�ӭ"��qn�{6+;ȫ��N2�_<��/aSLx���z6D��O(�Џ�[�w���N�-n�oEp�H��W*�������=q�x��X���9`*c��Q��7����;�{�|@�r֮eO&Dos�4�a�}K���q�7��QVm�Ue���9����j���r� nR�=���ޛ&����G;_g��CA��a�?��N���v�B�m���Kn��"�Γ%%�*�;�.P6 !Q�Z2�� nf����*��2��z�y���WR�}W�%ˮ�1�I���L�a��L�����^ٸ��HLR�D]hͼ9�{(�j�Q�����
#Z�*���Oj��Ղ��ђ��xi���7�>ZN��ߤ��ً�Kګ���j1.�ΐ���u1zi���x�+Oh��c��2x�*��3A��1�O���uV��GTE�梾�K���(7Y�CGkH99Ǯ�,�&�TW�5��8��Hg:mLڵ���6�@��m�?R�,Y/Olb��d�C�ph��uF��0o�ד-W٧�S�]5���rY���z�m ��;V$��oQi���У��o�3���{,W����}��3�]Q��XuǑmU���"$���;�w�b+ܗW�ύ�a��ҹ��1S��a�k;��#�~��HW��ơǉmly 5�[�O�Y��39���OB˪ v���qu�L3��p��9_f�#�zU�S�h�{tH{w ��o b�������+$S;v���VM��$;fb/��w���|Z5�7{0tOF����îkb���r���2G9�7M}ʧ8�$�-U����r�.cdL<<�CP���sZ���7�7�ڝJ���Z�O /�����txS��ëj�%=v��ge
�wS6��l*��k�9��Ӷ���{Fiq�$�9wQn���%;:W�*�,�\�D�V���q��ewKOGB/c�nV��N���h�k�Vs�Ҽ��Ė���^��Wb��]�:���ɁU��)��D-��j
��w��=~V1�^5���"9��w��ʅ1����lwd���#���<z��`�JB�y�_�_��+�����$��,�L`=���{y��F	کѤ�G��z~��:R=�e<���,��5�4^�LŚ�`\���f���{.gƼy�U��
/k���\D�참�z���C��8o����q�I�z(�G�X䋭�e�\G��ʼX�X\N�}�����{M|����e)ɾ;��e\�ߵ���yh��9��GUv��^���*<��UP�Tc�
7����Y4�X��k�U�oo���Fu�?b8s�a:ͮ����.b-m*-/3V�iw�y.���(��.'OS��h<��?l�US�uNL_�����y,�i��(�(�e�{�Ӌ�h~����+�ٷ<?T>�f�������X�<�r	�M`��E���j\.�Ӳ+��+q¿p��{�I��e(ُl��ڞ��LxoMup�W%�"�h~θ�y�h��V]`˻zcz�3u�qT�i�T��Rb�VG8j�C����g�zu�-�k7�;k� ��s��{�h���/~��",�ӎ�U�᡿N�MA{�qU�����V�Z;w�p��يNG��Y�)n�������(�L�Z�*�꨺P�aϼ���=�K���1>���gY��O޽syҍt	�C�ك����I͊���t+/}^���/K�\{	�/��yM!���.�׋�q�΋ۢ)����<3P|����NlP��,��:�d��כ��;c�Y4^���2��������=�u}=�I+��<�h�Ϧ@�	�ܜg���$�B�!��&���{����|7�2���������&b�	�u��?yu�v�G�`������ecK:������N�@��%|�ި�ɪǏ�zPNzQ8����Y��W��z�jFnghTz.s�q��|�^�L>;2��H�|@<|�g�C�#�Z��@��/sܽ#t�����V&/����^�c�P��t�n�l�P�3�����OB㊶�w��sC����*�Y-���i�<��`�?e��`�
��P�ה��C�����Kp�1ٕ=O���@柱W���׻�b*#���DѽϝQ�S��{�(ך�C��z��������l]=�R/ҙ��*H4kBō��K�:���գ��hιã�������ۄYx�`�H^
:��@S��m�nѭ=�hD�'2�vFm9Bs��"���y|(a'-7��o�;B���0��@:s��K|�ѰT.�qujk��{���U^���-�PV׀�,-=gs�c���"
<��@;���ݤ��.;�ƞu���h{��P�V��'}��z7�2P���#^&�Sa�c�т��΍�y,�h3�����'��]:��s���;���Z\7��߱�	�Ni�^ﬆ*l�Tc�,�`s۪�t��}�3+�����3Ϋkj�M.֪��.a�s!}E����O�"H͙yS73]jNg� �;�>�"6O���B����R�<��ѐ�l��݁\,�&}�]�cmt���+���6zWTu��ny.�l�l��P�BN�
��Ъ-h͜�nM8�9�Ifg��Ҽ::é�<}�:ڄ*O������w4n� T�}��F�����/�X�^\�A��r��\����嚁�3�H�U�cB$��:8�3���{uB���
:���<+�i��x%���w]1N��TǶ����nb�t��ޓ�o�O�L���x�=dtjѿ���a��]�@ü�2f7��W :������4��47���k.y��{�(U�t�� >0C���[ھ���W\p������檎 ����_m�f�іx1l�/C5t+�{��u%��1�h��;v�SJ�T1W,5��h�^��L���x���Rx�%.q�+\y{
�&<R�c��&jG�b����u�z�_q�7>=��g��}ߪS(T?��9s9_��=3����#9`*~��*r->��{Y�·Y=;Ps~i����<f��V"�|L�1ڎ�Ɏ��)�,\z���@l�ۧ���q�=ݷ�CW\��L���͖OWd��/�P�t@��!톱�R��w�X{֔����=i���@{�'����
5�����v_���ӫ�1v�(?2�_�'n�!~�/��䮟ZY�J��k5�p�gH
/\�*�TV�z���D�Ry�;��u{׹�x��6�o�xX;]U�^���֗����Z�(7�24v4���|���T�4�s��_�G����ޢ��ݒ�]&ͪ�&���Ki==q��sYs��C�Db��#ϳg����9����;�o/Q���]&~4���L�
S�����������ot5����T�3#Fg��G�v���G������9�P<�j�<�e�T��������?�����XB�%֫�~�bt��h�N�=�����cG/;[h&�6�T9�ى���2�j���<J/�Ѿu0��F.�R�Bث��mv�4g?�F�A�$re,a�����:��/3����f�x<޸u�_�$o�������Q�K�:1r�5�v�l�}]X.9q�qr�j�w�#K�9u׹ylZ�'1T�=�.��O������>]� ��9_k�8:��<{�sŨ��n���w\�:"�'�
�r�R�"�بQ����Ɏ>KO��Ev�4}�J�)���4��=�?SuIZ�zg�j���g�do��a�W��΍v[����JVE<�8U��C-�NW@��u��r {尻H)C��ޯa��y����=�*{*���2/��$��1E���QC��@&y��N�J&ceG]}g�0ώ��}��������ӕ���۫AS�N�O
�ԋ"b�zc�dw����fPS���ֱ�N�Zf�{=][��8t{�~�ˏ\Ϗ��呒�g��jW�L9�R�_j������:�)P�י�ǋ8Md?���!׭䮳jӳ�x���s���E5��څ�:W֭/��F�NN]�l�p�*�����m8V=�2�͹�*��(��C�TaC�|���G��m85���=B܎~ź�^Sw����9}՗�S/i=.��H�hڍZ��y��u���Ӿ�Λ�m�똧P��WZK�X5j�s���G+�8�^j�=��N�_m8��]ܨ���G#��.��/�^s����{�s��i	nI�p*x���H~�9�U��u�W�>�/�OZ�w#����[E�'���^�V�pU�=�v�=7�u=����C��0��S��MeG��Zc�-/�M[-t��[e��;!h�?�9��΃mYd�y�d��j#�?_�������5Z�VFwBL�i���|U��*:�sX�`UR�����Z\����6��Y�ml����cÔ���b�:xޚZ��*�N�]��p'�����:���]ub��J�7�n�9Μ�^;���{�x,Y�:��xq���A�v'��Y=P<��k�3��2=P�ب΅E��{��'���Ң�.��0*���߆�_�I���?���$)�2��px.�<���P��6(QՖn�3�_L緷ޑ��	덙�/���֜U�tWި3�� J��Ͽ*\?m�R~���y�3T�<Y��="�/�ZO�Zft�ʞ��ê�	��3 �]�Д�k�����*�O=�w��Eu��3�<\�bƠX�%���j���H�E }]y�ņ=�)��6�s�^j�i��$��,��k����):nލAL;5�&��q.�b�i��+�B�H"k�v�����Թ/1��_@�ՔE)�\��V.�Uˮ�M�H�Z�F�$�ϵ��
�%[݈��T��A6�#�b#'S[Ƿ���{|��[��=0m�u����T[FSO.;i���9HV^��vN����;����n�N-%�:�K��8lw���>��;qH��\��K��w^S;̗Nk[�SVHd�a�ګ�9��'���z�po�s��)Z8en����)G��c��YN�w��Lx殾v���}�ҟ۳b�9��c��F�m+	�e��ͱu`��=�޵*-9QGv�
����[Z�pt��IPӗQ�R�f�F���j��M53�T1�w����c�j�����ͽU00��:�KV+����̰�k>��um�.�5�����6��1�2�J�d=�,"2��-�45\s���n��{(X �d�CB�,j�	&�����S��i�����Ǐ�L�nڨ�mCJ��]9�0�;���eG]Hb�t�{��+Eh�]��kټQ�l�����ݱ�ТUw�=�n�h��=�`��FKY�^^׽�Q-{o����`�od%%Xqs�1�H,���5�Ny,���V�f'��v����.x-۾���n#xNV,�V0l彚�!p���%;x�%X)d��ή��"�`�!K\juXI�#�Ɩ�/�x����w�`vv�t�Z�t�NZ�_MkOW"mٝ,�&�PgG��al�3{2�su�%��QὊ��Rd��p���a��Z�:Ɋ�e��m1�m.���x����+J��8��u�RK�ˎXh�8R�7K���Y%���U�(�LfԒ�h7L��67\�3�%ԡ���������Z��bg(���Oʏ���M,�-�E(tξ����\O/v�[ ��jg�U#Rs���`�;3;9�7��}��踹�.�,�)���TN� pU��IN}Ũ�i1f�?�l�+U旸g-b�Jd�u�$�@��}a���p�+�-�����69.�P5����u��)�J��4�|H{@&�;DܝՊmfh����+����Pw&��,ݾ������>3%��+Q1v��ԇ��2�M�dnX���!�ݺ�0.�씳�#�Uaf0n�v�T���%.sF'�/��{RE�JmR��c��G�n������*���XC���l�J����Ei��RT�1q�Ϻ��3���F}�����JU\U��t,��E�l��G�G'L}�kh�O�X#렁+e[ǣ�����z���7Eҏ��i�������j�����9E�3���M^'�)�a�N�9b��}�w��[A�]�8'Qf�Y+gZ�ҷ6�A&��Rn�!��0��4YN>�u�vc3��o�Z�J����V��������ܔ����J�랣=r�M�s��$Ȃ�"�\'=O0�3+R�����,��BYb܋�E�p�;��DN�4N�E���P��ds�v�QN&	S�Ny3-R��ADHve�$�V��V��e«�,Vr�"HT���e�<9y
�!uQZ�Vd!٭Il�K"$�r�3/8��3�QPE���Q�'ݹ(�#,�Y�TEW��$�	hEK��NNy䉱D5��(Ɖ��k��T( �9\��
�Nt����(�s9N�����p�q�1hM:gH9ʱb*�0�jv@Q  H�D��A*�����<�.��b���f�O�1��Z�s���o�{����җ��-^=S�˔K��8�^�e���ͬI��r�7�#��h�G�v�j&��5�03i�{�����H��q�}U§��0!Eh�)����ox1=af`�'���5�O��M�f�+qK|X
2z��J�@�8с
r�\��|s8�gǣ=3�WϽV;I8�r�ug�[OuA�O�����0z�m��C�6.X�s����ժ>���)Gy�z�FC�����e����<3�YE݀^��ҽa�33+�À��E�|�k��x{?1��v�~�D+����@t�����xAN7x5^���:"��k���"��#c^�
��u��#]�/�дmC̡Z���j�V�R�B����I޹��'�wP�,��Qip�7���	Ӛs׷Z�5����\��=<pe���Ǟ�Gtv��$	����+�V�V�@���}e�\FR��P���9�߽�7���w�uI߻*��j������5΀֑Gt�Yi��j�=kd��yg�,�R�+"n�h�=,�}���q؏�t��di��X�>	�P}�ˎ�b�^�=�������w���z����dgܫ�ˀ�u�֬�W��\����;v�o��;�WS���h����R�����WZ��������H�G��n�Wm�L�M�7��ä�-�̕t;M�-R����3�3��=z��Wo��gs\��١l�dg�	���:�.Á�ëa��]N�@���hO3f���H��x�o]�󋋝���ݼ��c���,<k0�P������9Z�u޸"�f`{zO5�=f���cO���+�����G�*d ٪���>����� � k�����j���9���kq7����<\4�k>D���3���@�߳�ɝ��9[��^=���H�z�~�O"�jO	L�w�+\{ӁO�)O�1�&wTo�1#�c.���vQ�V�>/�e�؁���)�*���K'�J���X��8�)�}GAx�ͽ��@w����7�Zg��w)5����e��㒗��/�>�f2.L��<q˳O�V��݋F*���,�?g\��==��jzlTs�9�k���F�f�#���W�,���wQ��XG��^T��܀�b���� /k������M�&-���(؅}��K���ON]�/'�k�ZrH�\����Kܫ�Y�ĸz��ֲ�L^��Ɍc��B,���O_o����:�R)h�->)��hс��W\����=(R��0qy�����
�/o�ߩ�z`Y;��w)�з�:�ʼu���(6��|�rα���=�C{F�8E<����apԾ���9J�K*}5�t�]����g�e��Y�c�;ҙ�Z!�.|<�uU�?^�C�K�EE������:�O���"�ߔ���J�|�\�HwZxjd��\�/~�%��0�mU�Gh��]������p�{���{�z���{E�V$V����m<-N�=�1��OQ�܀�l�\�t��޹�΍� z��uU��g-+�g���ƍÃ>�[/6�����pl�T	�ˠv//6�=�r�f,n�{��k�P�Wr�X���Q�5>��P�f�s��#º\����P⻫s���I�u�q�t
��w�H��6����d�ԫ�P����L:O+����rF�#�6��]���G�zt. ws�$qX�P����R��sb�����홎��^��[��v��l���ۧ����z��s<��ْ�2����KUfEk�����}��/ʏ<�C��ק�Q�Z�=��z�
�+�~O��4eCF��)��s�\�;����X��{���z#�Ǧ>�$�A�L>CyVʑ�q��rJB�y�PT�u�`�bK��:��j4{�-��uK��36j��dz���{�z�j��\�uX�M�JJ�^�,<����k�ZR��1n���v�I\9�dkx.uJ=xm���N��x�w)� �a<:�Ӷ���^̫���O#�0�<8٢�����&�y�������9`*}<8LmT��K#�s��oL��P�P|��
@x� Jͯ�~��}l~�=�����~T����qŉ�=��O
ԯ����]K��/��}��dڙ�!����ׁ7Uۢ���4Z?~f*���ׅ�]��jP�ƹF�!��jz��Z�dM�"���L'�w^�q��
�6z'��L�\ۚ¬�r�d[^u�~fgqR�<1��ۉ۝����}���/ܫ��=^륆�|�N�=j�܎�"���b��;�Ǟ��o��9���]�u��]�$3+'�z�NV2�f���z�鍧�L�#zZ����g���n�p�s��=�;:dY9��ZZ5�d�l�5Bo�p���C�5Z��VF\wH�����w`��~��������LE;�'�ռj-&��Q���5��a�&,o�;��7ղ���w�n�Wf�^�ϸr9ʍ���IB�?T	�Z�*��7���C���5�{��&<�p5k���_�{]��C�]u~�����_b��;�c"�(w��Z��3s��K�w��d�!ytVϧq���/e���dQOZ�V��|��_�'�ě^�hF��.�m�;I�C���~j�(���Э��[ݗ�	�������q�T�ݰ<���FAW�2�����ֺ��j�˦Vw>�i�(�ǖ'[�́ǹX�\8�������5�$��J��̴t_�x.f��-.!�v��U����<��Į���̈�J�v7�p�vd��ɨ�<��k�u}��vBzj9B��� ͟�*�^P��z]�R9�'��LfA�ZY<o��F��x�u N�3 �{���h+��;��5_�O�\����GGx��K��LN�J�_qzuL��6����BG\f��k�9|��8v�	H�7�~����#?}��J�L>3��KI�� �v'�k���*�Ko+��_`���MtRyp���_*���gG�R��`/�+�9������"O��o��]��ջ'G���ޫ�j$嚎��z�a�mU=��<W�?_���߳�*��;ίw<�麁�+��S�U�s5��؊�v'<yF�>�TE�zk���՗��o�f�ה{���C�FK -��%w��F����'m�[㐚����&��rJ�v�V�=�S��/i����Y(1�Κ�e�P�l:�֌�gF�審�`x��9��3� ���m>���q��r��]
ۧpV�(5QS��]q-����6�ʳ0������Y®��Jn	ci+�{h�QoW=;�Yb�1\�;f��(�v�kݠ������gG�w>\�ݮ�cwHc�Ɠ�������j~��^V4�sQ`M��u���<3��a�ٌ�5s�Es]~���q������_s��W��=�8˿� ��s�6�uX�P&+�Y���|�2�7X���g�����9ٔj���7��t�f���k���j�,弒��_ӵ"��~�[������qC�<s�zr�M��w���R�c��)��"��WTv|)4x�����+��m$����Y���/�e慵�G.?W�ë�I���p���GO�����5��2<��=��S/���aΎ~���="�-��D�Z��x9�X><��/��������W�B��2�8��K~έ0���Ɵ�� /�~�F�?l����w̾���N�-pj�O 5����ג*��G{*��Ws|쾢Ù:v�r��s�NIR��x�Ļ3�9Γ&fj�g�Y�w�u#�^8�l�O�a�@���S]H�e1uݕ��o
��v<X��ճ��}�13�щp�[��Q�tU�qGDvB:f1����?H�~�L�O���\L�~����;Ƈ�;��x���y��͕��&�M&�؉}��r��v?�g�{��C�:w���&��_��u�`�|�F}3L��Mvd��4������Z�b�����3����=��m[�ȋ\uwS<�F��t�1�lGK�g�;�xWnNN���y��@���]1��0%�<��>��]��~FP�7�����x�Q~��ߒǅ�)T�^��H%�1í��
��&%�zlt�}�_s�9�:+��K(ۣ�.35~�\,��څf��VTw�l��4��x�� (֫������̈́2;%+�s�"��[3�{yU�����r�]`�פ�\���ե�^���Vt���e.Ƃ�~x/�l�'n�M��d�=>�������=�E��χ���:������V����]:��k[R�&A�m��98[��}���x��Lz��<v�;$	d�L5�mU�Gh���XOf�k��܃�ѷ��u���鱼XC�Mϼm�xj��9҃1�|'���ˉڰ0i��|e�/��F��ͬ���Y�+�>;Qj���7'��>�y$z{��8\j�����<��Sq5Qg��M@w�U"��@]5�UE�ܚ�x�]ӺX�����	���%�Ч=3y��������5Gȍx��#Ǫd�Rص�׽0������s��o��E	ۦ�(ǉa��뵂��K�F�.�fp&���x.��}G��@��5ն�9}���Z�ܻ�(��s�(iV��7R3!
[v����6���֞b�v����@h�[<H��87�d�.���<tX���gg�5+�I��Z4ʬC+=�e��ytDәh���<X��=R��sb�xn�G�����k<��>'�av��=(��y[)ƀَ�&��"D=<eg<�KUfEk]���o��[d��{��Tz:B��Y-@do-G�wD� ���~[��3�:����:���8��>�Qܬiv�G��l��:=?F�%��͑�|��r�t�nT �}D���jQ�NvtR�|�n���k����Z�ư>�8N�O
ԋ!�'��ǣ��h_L�;�1wJ��i�I?Aje�����Ά�0��P�IY�x�8�2X�zxx��'vX\]�8�@bes��SW}���{3�b��a����:h�3y�������h
��"8{�lR�x��Ѿ��G4ǰ���}t�j�H�%��z�H����d��dy�沕gF��#>��SY�o�}ݓ?K֐���{�Q��T�3���|M�s��ٵ�X�Ɵ	�/���9կn8�w��%�^;ٓ��a9ZΩ���R�p�&Y,�-3/�6����ԍ�ڗwӸ�+1&�+/���в��]�R����y8��0��<��#J�T�C��CS�O[��<˰E\�
5�Xt�/�����}!���V��`�{����Ĺ��m�*��0Tp8`�q����C*@��~�ح��e�O3D��y45���y��t:�����>q��ܨ���<ܱ�١�f�ӯfH�ց��1PK�?W-f��a鿲�l�g0�K�:cL8��%M\ɜ}h���=鑇�Ķ��d�)�ub�_fշJ�t��:Ǧ�H�ڻ���-Q��؜秀�����"��24�BlgB�O���ެ���{=eT�+�P��=ЮwMqxN��x��9���<2<��Q�sb��.6Vw��y�㎼{����d%���8�5��_z��Wt�D���˦'Gm���CP>�������`G}[�����}�����|�M}��U+����S�5�}����e��gs��wД�c�Rn�UM�?i���c�vBbw��?>@oTj��p��&�lf�=�I\�:��u���X���2W����^a)�:���K������F��_���=�7�R^�@~��m�AN��xJ���M�Qj���Q������vq����LWJ�j�hg]��n��{x���0!O�YS��QtJ��Z��c>�7�κ�.Z(LnM�wj]��<2�t"��ҧ|T�W����_���L]�l�������Z�Yj�wk���:d`����� W�t]�E�44r{%��)}�c��r� |/Wep��n�;�����P>9�P����c�2���7W}��19�X��Q���v\�O��{�������ݢ��ҰP��?s��V��y�Wg��<��}��W�(w�%�5���v~c�{���u�G���9g��ӿ��t��Q����Pl�E��+�K�j/��2Pc���OS
bN���G���)F�;�+��ٹ��7����V�SmL=��O�Mp�7�0��њr��5)�/�[⽷G��C�X����Ign;$	a��ȝV�V�@���Ղ�㱗s�q�8\���6=}'ga��;��,;9�N�\b�:r�Hth�\�H�ԁt�O���z��6��^/_�wx��c�>fC�^��������Ҹ�4�&�d����E����Wf�_�aR�����~:;��K
�ϫ��g���ZZhw��B��Fߌ.�Ecǒ!s�'��}����e�db�Yn =�L
��H��2���9U+B*�Q�o�X��T�&&UU_��F��1�1������"�w���*�7K�E�e�n%��<	������.��8B�"�!6��}0��x<�;������� t*�� �fX�yK�7WJ#`�+9H{�e%PE� b4��1���
�_�_D�74��S�4�V��"����K�������Ӟc�F~Е���o���∨"�I��s�;�x1� ��zU_�@�UPE��z1	+C��������������'�:a�P:��2�V�$��z"�����Q��DUz����Ѐ���o�1dR1OY5�?���],�5ٸ�߷��iw*=�`�ӑ��,QPE�vZr���MTԂ�aU^ W� AUX�"!L*2P��7��)��R��U4�>�ʪ"�QT4o��/�M�w�˴{ϼ�C��\�����bi�_�����=�'���R/�m�I�PC"��-z�uK]��M-�?��`k�P�t�|�h�Y[��q�}\�tu���ը��׀zt�hs-�Ǽ���H��.����0���1��Ω�\(D�U����G@�Q�DT}��0��p��LJ�݁�.�BA2*>���� �`���0>CF�l���������Bԑ�y�7��ɼ���p�t�a?�}<������-!&S�Ի
��\��"��:���v"�M节,]�q�������O3���[L��������@N\wwK�
��9q{2�O���ٗ����EA����lmA��I�U������EAWΡn�0h}|���nG���Ԛ�7h44�F��R�D�Ý�
-#�����˻,B��$>��#���P��Pm+�[�Q^=F��~�i<.,�w^A�M�jz �C���Zw`T.Cԕ� �@����0/���tx��&���Z��C����vv��5�ep!
�NtyR�,�D�~d�ٖh嵽���H�
����