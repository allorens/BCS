BZh91AY&SYM���6߀`q���#� ?���bQ�}T        ��
)_fh�U���M(�"I����h(j�&5�*�LR4֛Yld���j2Y����ѱ�fj�E*
SF�1ZP
TH UW��"��&iA�b�m�֒B��V������cSZ�DR�kU��
���3iU�j�P�Զ$4��Z֝j�ƨi��

>n�lk,�i��m���m��ޙմ�������Ubڬ�XX3MVT��4�6���l�b&յL��^��E��h�J�������k�6km5-�vWmV�m4�G�@ gk�꭬hu�]̧w:��:wn�d��әk*Λ%�.����P	ڗj�Z�:ӕt+]��GJ�b�mۑ���� �rͭeMQ�Ʀ2mF6�4���   Z�[�܀��3�
�
N�� 
]��s�( ��Pѩ)s�pAC��r����Jw;f�+F�%�X�4�mg'.��9�h*dҬ�J)*�e���  �x�U�����E[�gT�B�+���E��ܫ�xA�K�VS��
P�G�zU)T�s�h/e��9�@W����PU%x*���[+5	�$���  �<<@UJ�����{Ώ6����҂wOx=*�GOu�y�P�����JR�u.���zx<���m盉
 ��ǻ�Jn;Vm�jUZ*��m��6�x  �l��ݩEWMsG�݆�@맞4=<���9μ��P�^���CJ��3�4*J*�h�:�
U�G����R�&�̫�(�,��ЩR�Gz��+V���&��lj�U7�  �ݺz(R�wi{���AB��^�N�����^�҅)�K��J��J-<���=�T���m�()[�v�lq]�WfN��Z� 4��JvSUZ�d��fmQ��  1�B�K��R]�9λ`R�g:9�҂�'8�ХP��� k�: ;q��qw�(��� ��M1�Rme�[Z"��)�  w��AM�� d0 5��c�u����� �7  ]tp (f���kd�:t�6�4Vڤ�ci��+M�%a�  ;���N���((�ή�+���M���@4,w j��]p*���t
�:� P.vۀhs����٦���6�L�^   \� 
�N:� ;Q1@
����lS��P���P���@ �h�@.W8:Ӫ���}�    (50T�P	�04ɓ	��S�4�)JP���!�F#d2O`��R��@ �  �O��MT�	�  4 &��"�LPzFA450�P�F�& ���z�)Q��     ����	gL�)g�1{�ؽ�Zy9�2��[[�,�S�R&[\�KcX�
+9ڕ9��������b �+�G�H�(�eP$�'��t���|�nπj�� �������pQ����3����(�^�|�S���Bu�$��ib���� :@t���IzK�^�!�/��^�����	zK��%��^�%����.� :K����'IN� :@t���^� :X���C�'H�%�Ht���C��H� :C�bC��H^�=$:Bt��	��=!�H����?HzK�zK�^����H�����%�/IzHt��H���^�%�/IzH}!�/HzK�^� :@t��	��� :Bt��� ��� �H������I�%:H%:@t���$:K��	z@t��IzC�/HzHt��IzK�^�����.���/H� =%:K��= :K�^���/H�􇤽!���=$:Jt��	�S�'H��(��!���H�����􇤽 :O�:C���I��t���%�!�^����8��$:K���H��HzHt��'���	�^�	��%�!�S��	�	���	�S���S�I��%��C��/HLH|%�'���S�*�!T�@)�UN���G��=$E����N��p�S�= �/HzJ����t����t�S�"$�
H@zJ��@N�t����%G��t�C��%D��IA=!P�'HT:@��N�"t���?HN�"�T��=!P�'IT:J�� N��t�C��� P� �IO	� �IP:H)�O���!P�
IU:B��� ��C���H����!P� �I:@���t�C��� �
�H�zJ��N�"t�C� �IP:H!�N��t�C�(�$�"�I�C� �!D� 'IQ:@�N��t�C�"$�*�HP:B!�EzJI�B�H:J/H��$W� �^��Ez@/IU� �I�(�!�
�H :@/I�*�!��Az@/I���􇤇I:K���%�!�^��:C����/IzC��􇤽!�/HN���t��� :I�_Hz@t��� :K�^����$GHzC��Iz@t���^�!:K�^�%� �� :@t��!��� :K��I�|$�)���HN� :Bt���C��"$:Ht��!��H�����%�/HzK�^���'IzK�C�I:K��zK�N����?H:C�^�􃤞�O��>���{��N�ݟ��a�A��6L��1y밎aA5f���6�q@�V�˺8Řj�x2yHڑ���hI�m6�\�w��������q�lZ�B��of㖤�Ⱦ�5�K��E^c(D �1�����l�TY�e/ڎ�T�EZj�Î�4芲����В�e'D`˨Xf9����*jŧ�/jG"30L���ܨ@�(��-;�������,�7�GYc!��)±p�:�$���� ٴ̹h�th��E�vLV&ޏ��m����<��A�:7*��h:*XB�7mIHxVR��U�="�7�v+p�䲲�5�	B�!lQ'y����Vt5jˬ�a�ɮ^b����D��é�ܪ'˂���,,��>ѡlFf�&�m��ŵ0,t0�3�`�2��abw.��ٻo^��TH�����t�h�72�����hB��I�S%mIq�1�W�����H|��c��ս(�<+���]{���@�z4�Y���"ν&��9e���/������dӮ\P�u`��h���V��#�����*�*Ǹ^պ�6���Y�2�`�l�5-Y.�N��R�c�{v>�udf����3Ism�A�N��̵u�ŭ�f�CC���tu����b��E-�N'd�n]�D#I&b6d,��7�u��P]������k����2x[�q��^\;xQ���闌7�)MJ�15M'm鮩���-__<��/�V7�"u�)x��tі�Ϥ��W��(�W{���!銦��w�A�NCI��i޸�"	,�B�� ����0`��U�wRaB C����-UÃI�qY��)+�o(����4��Z��q?��2�9)���𗙺�Z�^4�c�L�M�$�W4���iԫ���m���V �,�i^�[{i�5lb%Yj�Fb��'sA�Stk%U�[�AZJ��\��{z�A	"I��M�c(��A|�	;���y��D�@�)��-`�4�wef���/~nS
ފ��w5�G+^۽����[u!�V�!6�aO�C�f�+C�ֵZxQUۥ�Z;�4�r��QB��U�G3 �]x͛v�mL�F�F=�#5fjh� vU�;��db�ƙ�,@^�1��۽�M�yGI;���Uڷ�n�i�O�_�MRz0�}�N0�ծĨ��a�-��M{�Yj��F��V���=�:stހ�^c7i'�͖���_;��Y�oaI��G�Imu��%즊Ŧ]i�E`4J��x@���j�!���4����,F+#��d�,��^��$�BU�͡��li�9���b:��1�핮��_@{V;	�Sdؔ���	�We��閪8�H4��[T��*���ɥ�p��hm8�$0�iRӍ&��[��&*�jS1bݿ� �-�<��Xl�P��oqPE�
���]T�dŤ�fmȡ3���i[o17�d�����w��@q��cD`�4���j��k ��&���i�1Xl��1��w��&� ,��#5���9WS\�4^ӣ��A�����Z-ꆗZ�����Xf���"�]�*����wm�6& ��C ����n��:4躙�(Kxc8DY�A���M1V���q+��=�k�b���l���e�Kǵ���e-�M�b���N�]Tl`�ǥ��+8��`j�����]XtZtq浼�}�i5ar�M���ӉL�	|���ȑAҐ����J��nQ@�)�-�*���YA�u��5��QOu��V��v�|/F�D)T�P%�vq��5��u��!X�uU�;V�ss�+���`��dӵ�Z�e���5"V�N��7��+��aV��ID�o7p�s��3Ij��V�=pMS%��;���-6�:��,�W��ˡ�Q�dW�ݽ,ȕY�FEK��t�.UC�F�`-N����S2��]ө��̺��[�Ӭ�X���Z�L�o��h4�pՉXP��ǠhҲ��H��bH��:'C�&�l�hi�x�MV��!X/-Z���w
�6�sA8�iɠn�Oi���ׇF?�q���EF�Um�ޗ��	�QA7F�tj�B�Y�Sф%c7x��-�K-�n�J�x�zb�q���,wB�{��ŀ�f����
����!wT�����܌ŵ�^R�q����!��fQ�H�Y�e��۔cv�5�[.\�J�0j����$���9��j-坣VFK�M�У��cb�*���n*�5�NK�zb7�)'Q�.�L7QV5�b4�3E�X�;v�S����L��z��2h�(Kkw^�3o!nb��HV;4���34�ٻEk̟�8�(dl�N�R�ܱ�R#	�X35��[wjr�PC��hi�滑t�:������cۦ0�m����>), ��zX|:�],��*6�7u�F�%ݖ3H�I�;h�s�v��Gc����RJ̅ò���BT�v^K�c�������$Il�ё��� Ư*K�֊�%m�3�ܰt�2��j��#(!���꼤ⴱ�;�l���.�N�7\���(�)�2���AS���V�&mV��3Yhf~�����G��iL;n�.�bT�e3d��ZQ�,J7�z�T��B��@kɵ�+�#j���)a��vK5f�+� 6Bon�5TChPr���Lٷ��fU�蠔~�D��/{�&�J�[�Q���
�E�:�ܥ@)d�v�o�Y�ujQcq�B�b���x���l�vv�,Q�F:ڑ���0�0���|&=QR�$˱e6�|�K1л׈<'{R�J�*��-�YxN	T�!��餱t5`VՆm��i(�aԔ��S����h������z�
y�TwB^=�/(-w�f���ɀ잙.�7K�+`�"��l��U�޼S3�������m�Ik%,qʅG�n�nc��YFG4k�o# �/p�*�ˤ��"����o
̪�`%���n��ӱ�N��1����HEY��6<#n���_75�A�%tS��#T�G��4
)3W�J��c��X��A�XEuv}u������n*�ja[����7u┰��f�&ƞ��<�,�h��m��I���@ˋ׺,�tT!Y�۬��Bư�Ɍ�tj�(n��u��g&j׫X(�����ul�
�X�IS��Φ��ͽ
�$�n���r���H��e��H�;Q�U+��2��������TE�q�E�Z�Z5�,����T&��M�@����-����R��D=f5����K12V�-�COjũf٬v�zU�E��}6���f(bV赱*j����n�n���ĉU���s �7d`'ȋr��VWm��ݝ�V����N��i#�km}���Z�Q��.�,�,Y��)�̨nQ�m�m���Ejřmek�+^�
���حN�f�� P�"�i�F�{q�s6`ͱ�b�0/�́8V����i;���W)�'FG#�Zf�wi=��Z�3��Z�&��/h1/+3r��n��1C���Qj�ێ����٨�/Kʌ��w�GZ�����Qq��cd�O"�6ssF[���~�X�����7F�G��H�;"enY8��;Vmc`Z�jHͥ�qȑ�X��ื$�D��f�O���#��7]d�|ZśLee�e��f~6��k�{�����F�4�'Zh�c���Tq���պv��
�9�Z͌*h�j�y�h���5��I"�.�Y������ۧBȕ�F�!c.6�[�^��@�f�-B�^1�nF�N-yNcF�AR��%j�X��	��4UB��Q���zv���Z����z���2�a0c~�K,"�<or�V�G�m��qm�ճ����m�j4ԱhÏ^����-�jn�X���v���d�;Y�5�ܱE�����!�fV��ɳSǲ۽���9[Xέ��L��n�=���Ca�"�&Ȭ#�����YJ�j٫N�f��JhШ�7����!���QCa�{�Qkl��z)^�4tQ�x�3ˈ��5E+
���Mװ��YMЦ��Cn����,ǣ	�VV��\!��,��ܧ������E�U�P����)�ƝR֑.��^]i4^�@Шer�Y�cr�O�T���y�K[N�Z����˵�6� aҖ�\Oj��$FΡu�!e(y�7*�6hD��I0A)Br�l��6�R��7�pdY�D�W�>���Y��ԍ���' �=����y3Lz2��L��#*�XKV��U��:��{�����h7uE�8��oT'Tj[�Aʆڬ�df���,�%�t~�P�F�55f��X�"�q\ȡ�w�x�*�=l48�w��Ql�p�i1Iق]f9Vj�8rP�oI�Nm���8e*�D�/����"��~86�R��v�*X]�q�Q�-��c�0*�ݑ�{��s?&��͛�r51�����P{�tl�GH�4���m�nn��-��d�O�-�G�.#z��Je	tB�\��/$@PeЬ�wEQ�J��ʜ��{���{����G��Q����2�E��.9z��ۭi͚5RxY�ZyG틻;Q�D�X�d�x���V١��-@5n��f�i�O���-�:`�2�B7�1izQ���.�����{����cф�[,]@F���V�{��#5��Y�>;�le�*acF�w"8�G3,�[X�IY���ͦ{�v5���Fi�>�X�R��˭�ݕ�f��m�"!wM��鵇�a�[�v��+�խy[xM�Ê�$���1��՝XU��
�l�Vh��&7i�4
�ۢ�;�x�h�2���٣��70��)�M�v�Jy���r��R���䫤�!D8�e�z�b藯B�&U=w�`��Uɉh5�`��Hj@�׵
��U�K�@
�N����w6�9QI�,��ֆ0�qeM�[�:�/&��Q�? k|Nn��ba�h�ji�@�cI�'m��R�&�l�tm:ZŌ5 �LsU�1e�gf��TA�T0���K�+��F������4�gaT*�/#t.�[�)k֡����Ҡ�R�e�f������@�ю�+��ǯu�,*��',M�P5���P�Տ��f,��	y��G԰˚�r��C4`Fnf��X.Z�h��&�˪�DPZ�˳Y���	5l [m軱��EɆV�Q��U%�V�ӦZG!9���H������Hd��w�s0��6��pӸ���A�F�`[SL���t�c�Q1Vзw��a�aːڥ��-CsN�R��ڢ��6��F��`r���HM��:A;�3Z�8���h�)�%ѳ�8�V�S��ʢ��D��T��#�'��
Yp�x��JMy�e&��`����ցb*ӓ*���&�^���-&̒��rX��)5b��F2K�m��*�&�)����c�i�Rz��R�YZF�m�i���1w��&���ـ3+F���Ct�^�{z����P����ݸ.]I�p�Ō�Z�9f!w��(=�D��K���v���V��:+r�4� �4�)�.���'�7
vje��%	v8�%���TP��u� uSI�a_%kM6.e:���q�2v��0��ڳ,����TN=�ek,%��Sc0�+�Fa��m��A7�F��['j,H�C�'z)ݨ��%����˟]%n�#s�>27�N7��+1�W��)�t�b�Z>ݎ1{)L��+�L�i��d�A"cG����m�Mle\�[�kYZ*a˔����� �m��{MqĖa��m�K)�Z�X� ��`�}�QQ�yD����n@�ۥvr��A^Rx������v��3��4cX�q�u���z�{Z��e���~wWܺ�x��H
'�V�nT�d�4�M�փ{���z������2���&0]BFm��auy{������_).܂�m�����͂�W�U�q���^]CgoE뙮-�r�A5��u-�n��Y4�ةV���C[��6��r�4нbc,���7v�{٘0�r�K=H��Y�1���u�=t���o��D'�h�3wa.E�#�-,�%b9Y����V�O��a��ʬ�2��7�����R^mG�Յ
�C0PF�Y�����Ҁ�t��#@�L-����i7��m#��6�F�)��ǡI3h<����nU�$ï6��L�yB�;�9C-e�z�bx�]]�xn�ٷ��+�4�X�ʐm^P$���^��RY[g�M�^k�W�ɋ�Г��خ��٦P&��%���ͤ����c z���OYvf�]�������h�f�Db9)��9RM
�Hy6��1�A�o��J٣%�[[ c�Rl-��q�Ԥ��($��UM�̀���֙���:@���w�M�YW�Y�V��H˶�j��-�x�3��5��m�烇���2x�*�� qI7}�=9�D�4��
�FE��˴v�7vK*;5%�lve�<YGKF E�Y�4�n��3�K5i�DX��l��sM�gXɎ��#,�k�����`���E�ܷ.�;/2�?�4Y���p����=�p�n]j����(ir���"����r���0���Uv��(+qK����%˗��#7-;�.]RU�Ӛ�ViF�6Ye���t��NB�b�v�Ǯc�l��I$���(�K(�I$�I(�$���%�j�0�M��t�$ҷ%�a�aWMeɢ�x����(��$�IF�`�Nz����3�r���9G.�j��s
d��e�0�.�:'�CU�D�n����kviAc)���DîV-���2�;yi^�Ĕ�0�Ӎ^dA֍FT��*֛:I�K4I��0���IG�̠����A6m�w�.)O%J�ʶ��S����b8�E�w'��?�VO�Y�L��]�Bz��/�?�����S����y�{��?~~���gvw۲¯wzKNn鬤#s0A�s[��I@<pI�'��b}�4���pڝ��B�*?���k�����[*X'E]Kt&�2��7*�\�g��x�Zh�a��&E�`�C{Tj��"_4iՓ�c���=����O����&&~�{gV*dm�p}�]�S/$��M]�̼���
EUƸ��Ԃ�wt����y��j�kJ=ZV��!.O�q&�����d�J.����T�ݪ[tw���	B�
���V���:Q�e�������ZRk2�n��ٸ��W��d��lj:���ζ~܌�@sژ�7���lt�bЊ�<��M�Ւ�R1� ��0�4'��S4r̥7.�8��T�/l$�����.&Β�ˮWNc�JZ)ֹ�5���U;�9�,M@�V��^d��Vk{�6�U��]ګTFоē�|fӷyĺ��`�d{ci�J�\q�6�|]IXR�e��s�73+b�hu���"��P۹�X\��%:�E��֨JY'_i�]-�qn�����t�o�Ʊ)%��@Y���KO�mxHml��2��Hح���s��vx��F�7��Zib7|l������-%�|�f�M�"V��ݭ�]0�aɝF�.�+>C6�F��K�)��dpk�%J�U�Cw��� �Gv�n��VU���U����.��;Xln�.-yo&;�A�Z(�r�;ѻ;����qO��9��5�N`V��$����[�ɠU��V�����5��8 T�n�-F����Qft;J�l�v0d}�܆�*��5��t8Z�i��se�B��|\JՍ{+b���ޫ=��!m�-:	�]=Z*��7�5��-�H(-��G�O���.�Z��i�7�qwf����Nᄒ��G�زo(*���q,��s9R�%�Jm�h07����0�ą!}���	��ޙCE�`�rs�wԦ�+�]P��t���c��Īf-<!��խ�y0M��:���]�p�m�UN�[�����P!�����^i�Ρ5���Cv�$Z4h�6����7�E�������_wl�u]�/Z��e�d�ŢI�y�% ,�͠*^wRhd�d����Q'�)�Zəs.nU�c�|!��f녳!5טl�S-�[��Wi�W��	�]���Ӏ�4�p�j�(��c�w}[0�4�r�S|�1J-?�_f�zK�����lu�^õw�q��G ��́5���:�xq���qⶏ+�,�*8H����L2�kA[p7Na�\�gh-��Ĵ�0q�nU��\���Y�{4��"�Hv[��i�.�@�[bZ�=�v_�jzgq���˰�s�!�k	V��)�+FvSR�A����ӵw�tN�
ݤ�a5Ǔ��v�aX��5R��٨�A��)s���6Wa�hy�n"!���f�Y�ր�T�j��w��*N晫�aX�'
��R�l�8@��F���ur��f��{(\��I��RI ���8P��v|U	#�Z^�Ũ.���b�-:�|�$Sᚺ�۩S�Q�.��u¾^�B�fۡ��}.����"�9V��<�q��F��kt��D�]ݪ�u�H4)���qK�����YRiv�*���q�-����N�������h_.7�P��+���[��#w��J�*U��wË��G�
�=L�}]4�������ne :Z�	N��{�� ���֋B�(T�*��M�o2R�����,]��<�ُ��Y��hu3�UԱ�����^�9���7!�.�3/�ܚy�@�[��s8�c7�]��*�]p�sQ�<)n��m�W1��X��Q��f�Wu8�ǉʣѺḤ�~�dZ�A��ڰ�ȭ����wj�:�N��Z�4�����P������f��N#�٥9�� \�ib�D<�w��-F���j��J�p�٧6�-h�+E��k���!o"��}CJbaNB*�9��_4Nr��mhT���i�KO{�yN�h�=�A��!����U��V�_-�o�
��s�����̾5��С����[�$�j��8�v� �-j�G�%, 9���{-f��6���@a$3ّ���6%Y��kG:R.j�;��b��$�:�i�7��
���˻ܟ_�
��ڢ,����,ӳV�p�\�8�vr�{4Ȟ�V��u5�)��CЊ6&��X'f,�A��� vHޠ@�M�^7�%9��DI�Ť���g,i�Z5[W��-c����� ݼ�p_� *V)�(k��O�7Y]΅�u.I��H5k`����T�m�\�떜������NL)���p����1����hdGqa��;�;[�u��8��|��;hp�9Տ��t��_.^���vD�7[��++�,�cR�LKqhS�����޾G�e�J��������Mݬ�=��K0o׹��!���%(8��U���#&���J��t���@��Z�34U�l1z���]�h�Qum����"�[
rv����^�n)G(35�x{���j�ڊZBl�����ƪ�:��T<���c]fQkkv=l�N-�8#��C)ml�KzZǠ��wf�mlN�l��W|�]$q�M�/%)� ��'3D�"����t�YY�x���XZcJ.^<������*W9��{a{��ͬ��7����N���I��<���S(�1h�Z�D�L�&<�НI�gv��D3j�|�84/�4�����͵AO�8���E�ȉ�a�����P��C+Ntʷ)�u�5��D��2��}�ɭ\s�豾}�k�傱��ή�l�j[r�,&���b)��bsp8�:��r+n��B����fbKT�w/N����=�Tu�[Τ���L}}n��4�fY���u�t�N*K2��	����K�r
1�����@�������{�q��#��7>���O��ȝ����f�N�͙�hc��B����r�H��4����U��r�`t��Z嶬> [��F�
[+���p]��Y�#���o$%����c��h�ٖ
����&�'�oQ����+��]�� ��+}J�>�7��v%Wbg�u+bf�0^j���	��W8bg�<:��ղZ�k�zwu������:YB��8���wlcU(��)�Ʃ��5�J���u���R�Q[��qei�K|޴̽C#�{;vn#.G�q������{���u]<��2�i�b��:���-�n����ys+N������l�*S���Zىx��f@��ժ��k�0���Ц�
�oa�ZP����c	f�ֺ[e�%�a�H�nA�g$8c�!��������ܛ��N��԰`�*�ْItW�VY$�(�W,�>�)��屈��M�ta�Dqnk�g0#�]R��w_>}e.�У|IT%�y��PyF�
0h�+`R�-��q�pΕ��֦�����K��iy��|3���!f`gp)&�j��ox����1؞���u'�� �p�Y�9A��(:)&��P�
d�I��#��Xh�{oq�eဖnn�p����Zþ|���5iM_7}�&r�x���H�h��d�4�ܭ�z��h�D�_eM�D�dk�)���6ۺ&0E�����e�1�N�:���m�xQ�u� �N<��I���w&����-�1�m���+WQ�t�N��r恀n�z«�=q`����a r.��˾�\l���a�Q�1跓�F�eâr�dࡅ<'T�&b�9��v��BtZ��Ŧ��.II҈ώ����M��6����\�V���v2�0���e�W=<��ĒR�\��� �q��k%S�7�?�|��w�L�Bc��j�1�ViF�+w�4��.[��͖��b�X3s�3{����r��;����p�4�jtG��*U�ջS�^݃l�M�-=�\�z�Ԟ�C7#�x4�ʛ���K���k��9u�a�6���5=ϰ_�r��n.����}V-�G��5^^5y4=w|q��A�Smc����@�+��������*<B�@dv�e�{��fb
����`�i\avb��|t[��N@�����绁Kux�C���ذ��4�C������e�'-�. �\-
�lvs�<�մ��6�L�v�L;���,�k.�)�����	J�!��Ȩ��^�W�{-b_7��a����r�͐��j��L�
�G���[��P..�g���(��X,,]c�T��{"J�˿�	<��2�fj���k�%�˜B��X�؎I]ty���b��wj�Zd�tV,7�!
�QB�.n��5��)��-7 ɒ��Xᳪ�r\���l=�o.i��\���g��*ړS�۾�玄��j�Ԛ�u��:��5�^o_�de^ϲM���c������5͇�0<�mނ]�.�.W)���w�f��bt��Nd�zj��t�
B�%ډ�2�e^!�=r,&�Wd���uu����,�Di��L�{=�^��z��=�VX�0.iB����y���,>�R��t�st��Zj���i�KF�K�{t�yF��/*ec+Ol�MO�5��{{���u&�B�q�*Πf�J
��ح}�a��R��n�A���'6��d�fl"��M��9}�tN[��yǂ�v�S�i�j�Ky�7�ŊAѭ3�U�����0��`���|kR����-��"���\��/v�[(�]�W���G�sx�N�蛾60���X�5����==[�o��}At`́�.��^_+��L�y�Q,e�c��<�z]MvE'8)���g��
jc��*:6P2��|;fPT������R)C{Eem�3Z����I'RM��LW3vNN��tc���Zf�zѨ0p�٬y�u�Gz�[!<�l��"����&W_��8Yw�^K��]�O��Mއ���U���nfϷsu�]"v{%ZYP���=�;K&�ݐ�\�ݙ����[=-6ڰ��N���qZ[)�ýv��2���KAt��&t�M������Vu�S��wˁŮ�'ɶ1s&ըwn�����.4��K8}�@K=t����J�a	�����Rr"[[�_k��$^�v��hj}���et�.��L̥�z�A)y�����̱�9�&�>�֕um���%`��!��Q�C'mCMès�ƚf>A���:x���,�D�l��M���b����PaR�v���S���_P
�Թ���$��>�����[O#�q�:^,����B��y�gyQ�o��.���Iݕ�Kt���*���z;'%Vr�Q�E�|��pV=[1�4�X^+��:�:�2����Pq����'���V�,�7SC�wkJ#�݉h�7}lGry5�?n�����9F=5դr�kD[Y8�jT�J:�A�&v��9B��'���V���#�=�f$*�}�S�LGu
;Rm�p^�-3x[!��\�.�7�F��e-Sw"ۭ�me��t"r�=&>��O�Q.���K$qyF�t!���ܻ��۫7x����pz~SX�iҷ;�)5D����`���լ�k����T���a��h�Z�6+v���_ڇ6۳oj�}%�j�����3ppr��ר;�|:w��vU:L���mKZ��Y�uNm����0��5J�=Q��(�l�O�r��٧��byS�"�t2,�]��t�#���5u;����Ӹ��}�j�dt-o\F��b�Y2~�
��������(�JB]-��b�]6�s��
�N�9f�{n�U�r�w�q���a=rt�>;>��d�{1x��U�ܑ���؜��V��Mh��"�������x� �z,��\�|8�f�ോۻ�g\�f�s�4k�F�J�]���Wl�&~�̝��kD�u�Z���d6T�:��&���s����1��DM�	dp݁#�k�@qsT��@&�WiX8�o�b�z��b��X��+X[.�J}����<jHTgܽ�w����
�Q�LG�u������w�C2M2jУ�a�7����;��\�C/-�a��h�A����s'S ��ܩ�${��H����|�Vn�ˡ�:5�r�*;��5�ʹr�S9�94��8ٜx����~�6c�u$đ�YjI��zot�e�4��޷ǜ=�R��m�o-Ӏ_9�3�R��H�����8�"��վ&1��ަ9?JKt�nM�l�@J�ene��*<]7������U��r2m�T4�l2ɢ(\��-�5Z7��.��� �͈�n%	&f�c�� `�$�mA�&u%�|Ƌ���3\P�.�2�����c�L�Zk�M� |4�W}W�r��U�
�𕹮�H]KFR7Γ|���࿖�ZOnL�)����,;$���3+e��yH�	7��t#p�gG�7gpR����L�v���WB�e��.Rl8ڇ��Pl�%�ɏq�n���d�W�R�Vj�Z���#]O�y�2�b����frY��n�LI�٨X���M�B�2] f5�|��p�v��gz1f�ń�w�Dl�k�D�"H$IE�B�Rgkr����;2f���Vූd�Ze�j��^�N�@���QS`�DI6$%B�N��i� %��"�T���O*�v?,�h��,��#��'Y�w��!4�-�c,�\o.���3_��!�DCf��vE�A�АZN ���l�dN'�ʹ�D�C��Q���3�X.=����d�o!2��f�9GN�X��t>�e���bɤ���Vq�ƕ�  �![$/ԂK(Q}bx����_�'_������e�BF� ��R���ԡ̓L����%8����t�HH1���*P��V0l����PQ�aʺ�vG�Vi�k���>�t�;�H�
�6њ������.J2~��HS?�÷Tm"���i�'d0�	
���\V���MٮKb�ft+�e��?X���?��5訿���(�����C���f��+JʒρH�u�1lYe�ۜ՘�k>�u R�e�o�����8���s[� J���>嫎��j7f��>�%!
��#&�EY��g+{��ꙻȾE��+�'M�����L��^���3�R޺�ʌ��QF҆=\X�엘e�G�6�:�vQ�I]7H��	�W˕ޅ�����{��N�#�.ݴk,0f\�è5:𻤥�=�C���USTާ����엯Kem��w�}�F�f��+V�4q�ʎ�Vee.�ù.�zӁ������q7¤�K���cy��b5�L�f�)�*��t�s`|E�iQ�uki��/�>�э��QJ9����1��E���\[�zv��e�!J��:��7j/���S�:���tX_t®P�˔`B�)�7l�W�2L��K傶
�qG��ֺ4���D�N�Z!�*R;�]mj|��8(՞L{N ��.�����X�j�;��V�s( NG��� ��k�q�0w��*��y��|���u[cF��BLJ�h(��+q���b�7��9�Y��rF��/22��*��>�wnv�I����	���y,^�=��줫�[��
�6{y��ne�Hb�݊���'ugB�j�+/]���,7�NlfN�|a�#�A��G�Z�d�فc��`Iwk��u3�ҡR�J�*T�R�J��8p�Ç8p� ���Ç8`�Ç8p�Â8p�+�靲�D��u���sm���j���9���N�$��7v[�jl��)��=�V�5�YF�d\w`M��벲Wk|�e����j����۵��i
7���X��7�J��:�$�R��x5r��![@��r>�Ô��m�%�Ha��Z����Y�Ql�%�xE�J�Śc�C� �ͱZ�f�7/j�[?�b�88CYf<�UL	�+H��sΡ�l�q}�P�w��FI�UU��NL���_tVa١�KP�kx��}��v��g-������s:d+�E���/{���QV!n�P]�a�f��R�R1�,=Nb��Q���e����w:Y�\��l��C��((�t89ɍ�k�ڒ�OBe��d��I@7Av	
;���_)D�u��h���fj��ΥB)�*�f�$q�(B�K5��.#�b�S��Bn�{�a�\��%�S�����-ZQmݶ:���K�xy��Z2iB���1SzT��֐jR�X�WJ�*�멃�S�2����K�t�S�v�d�b-��aa'(�Q�UՊA]j��\vd-�	Z԰m��sUE�S�p[8�7�gs؜��(n��sF�:�C	�D�]qv�[*g%��3n�u�@�^ԃ�c ��|jb�be�z2�xr��5i�{�eu�Y��A���0�Tq����8H�cA#�8P�Ç8X�Çp�Å �8p��8p�C�8p�Ç�8WV��fw!����[�8PB��w���nn�o����#[$���\�+X��1�³b��;-ݽ���<|U���H�'��[�3)��9�0�d@��N�,�4TT�8Է�%̥0��+�P����Q:ᕁ�5X�֫F�:uX�&O��&sf �����L��v���&Q���^�&�Ž,,U�V_f�ͼoU�Q' 栥��tL��r��T�Ȋ"0���Q�r��K��B�s3�C��.ֲ�j^��vt��ó��L�n>;�{���kwE�H�!9��{��C�[�i���"kU�������G��۳ql�:�/ -�5l|��R�[�7J��,�H:�CimV��}$W���o>�fpk,He^S\l�r:�H��٢���0�(˭]m��;4���5f�nK�9ح�n�:�����Z���]���o�J�(XÔ���+���n�O46��2�&�J|�	�N��2�>�CJ�o9n(�rI�h�\Ƚ!����s~	u9k�9b�
�v���0r�D���XR����;D6�{0��BGwGw���Pm8�x��V�p��.��,0����	��O�8oY���lzq�}D�5^�ݮ���B��ЬBl�^Tܮ��I;3��
o:�HX+����O{64]���]2Nf���.�j��5��Q�J�J�*R�P!Ç8p�Ç�Ç(P�C�8p�c�p�Ç8p�Á�R�Jb�U�-F���n�G�U��So�n�k�%v�X/���>���EN`p�u�돪l?%�+��}���:J��Y������>�
Vo�G}��Oq����W|�ʾ2��sLָ���}j�v�[x�Mɇ�m�U��b����#�w*�{�@��!�B�>->x
��+[e^LkC�ݍW�k�kbWQuԋM�j��3� �hF<
��H���C\�l/Ǚ�����U�h`��o+fm��+M�lऄ���!@�-R�Ĝ��h�2��z�`���G��f91^���2�J���hI�}�b�q�9f�Qٴ�h\�٢�d��t��R�H��TB&o�X����ҫ5ҁ��ҩ�h*��2�2tt�R���2w}��e��݀��[�;#S*��G�{(&��j�s�+�yx�M�һ:Rꉹ����l����/E �5�nͥB����bʆU�陵0�YO���^*��\�^h��RR�;S,�j�17w�:�<�pЉ�V�`�OE�هgo3�֗|&��ga�bC�bL}Jj6��V8�u��8w��{q)��դx�s��b�?,;e��.���}Y�N��[w&�8��f=�T����Qo֒�اZ�녮�-�1��[/E�i�8�Zf��$$2K���ͽR�^Q!H�K�ӛ4�M*�Z����|�̬�@�,Xᣇ8p�8p�Ç8p�Ç8p��Ŋ �Ç8p�Â8p�Ç8p�Ã8D��s���S/���E�w����m.8M��51��EgȮ7 ���#ް�6؞���Φ�Z��`�qt���\*	��WL�tF%0G՝�����r���X�x����m�7M�_C�'��ov���F��uBo.��BnV��:c��d���E�fT���iky�ݚ'�T�<e�o[�p����c��3m't�]�X3D�{�ns��fU�V�1�C��pq[�K2�E�<�yIYv@��C��s(�!(��:��n�[mm�a��7���u_l����N����d)�˒�j����+�#$C1�6j	��g0"��f��C�v��Bo]��E���5�rU�B�/9Kx#�;-���'#�k);��;����sM[�
��5uw�fQ�X�=` �������pF�DR�����|������J�M�!f��E��M��Λ�J䶈 �Ҿw��{ N=�74��deZ7v	4r���ZͤV�;A+��ұ�JĽV�j�-M���t��\OS|CF�fZ�i�v�Ѐ��`=A__8q�}��ͫ.�H���YѼ)��Z�yJ:��Y57��W-9��0�X�lG65>�7���J�嬷K%@�<���;HF�wwM�����-�/�M����b��j�nT�]�'m��-�SD=�e�~�k:�V]��FX��G8p�Ç8p�Ç8p�Ä(P�b�8p�Ç8p�8p�êT�R�J�*T�ED�rq�s-�-n�!��]��i�\&�������x��XM�6�N�Q:��N� !��A�nR��M}�N�<�yZ��uy{Pm�MvVs�7����V��:���u�qt���e�O��b������ё��e_t6H�%��d�����)�|o@���&$����u�l
�T�	6Z��:�2�:#1rO�qN�����pv��:̈́Փ[��3A
�Uh�E�E>����@��F �sh�8캖�>��Ǭ>�&�q�D�)�Ӽm��"��o�Ǭo��s�g��=�(.l
�x�Z���)��$�͏t��2��T���Z���,q���T�b�,i�Yk��.�gT՛�-#F��+�o�72�Q�:*���ȣ�.���n���wi:JnW��r|�:㡋��{hKfG�F"�h55�!�N[��ʻ�/n5���&�e����¨�t�+)Q��ӵ��!Rn�N�D��ҎV����_�������g \Π�Ȉ/��$�fc�Ŋ^o<[*]4P�#x(�W0m��yNJH�9̺�TY`�/0�lNQ,�˕��BK�G���6�ܖ!�6K���p��/;8ǚt	w{�޸Wsx��ǡ��	֢1�1�!��3f�
��,����!���ː$M���ɸ�!_V�Z��|o	w�.p�×9|�� �d��>�}a-d9�S�ҍ�y�ۣVR��w�S��R�
5)T�R�J�*T�R�AÇ(p�Ç(P�C��8p��T�R�J�*P�R�J�*R�R�J�(<��#AxYr�t.�e�,Jݔ�^V���c�;%u�i����W:�>����Z�i�ŰH�I˯{�.t�c]��V	�F���
�޼?!R^��1�
�nY[7�ȅ�h����2��3��n�R͋�Y+����yG�c7mҾ�xq8���f��T���b��9��D�:d���l�TK$�e�~����ٕ9N�*m��k�09|�l�[g��t]���Nz$�+��ZGEQtn>�GZ�>/��%��坒��4E˫���F�&�G����4��^�}��)0�:�.
�t�2�`��.{�7lc��*��AuvͨL]�6�gyd٦�IïX���'�Ƌ�顈�UwU��|أ&s���;m��ۭ&�����|��;����2��%�3�N���,�E���:U�(c֚�b�m�9ڬqh@͝�ڜct�G47�P��-��GF]��ve���t�ff]��勉�}Ozhܝ�}�@��V��t�ͻ��GčǮ\��T7�6��No�Tt0"y˄� [r���:+��>�&՗R�z��2
�%�yd]t���锶�����Ls]Ez��3���p��7]`�9'Y+�N�네���̝�����������3�v,��b�e���J�m��2�Ɏi��F�]���BwV,8�Z�=m}�S�3>���N�Ъ��Բ��"��abŃ#0`��0`�S �Ç(P�B��8p�Ç�R�Jڕ*T�F�J�*VF�]˻S=�k*�XZ����GP���r�f�-L[U׷Ǎv��{�8�R~d ���0��+�o ���D\�Y�;z�z#����H�����.���:6���itR�2���c�]W�Q�u�e#�
�Q�`�μ�̺LL�-e%uUFQ��fݐ>�ᚪN�[�9#�B��e����Yu���Lmo�aܘ�TXt�*M�O
WyieE�����Ty�Q�5�f�֨ NU���N�vs�[����qɓ+N�[���*��ǹ��bN<��Z2K="��6Rʹ�2�����$�У?�;�Bz���ͫ&76��d�fw�yw�0�UmS��T`) �ۂ��֦M�s��7BIӺKw�M���9��C����-\ʪF*��F�>�q͑�MS�6*�m�h�Y���=fs�%��X�.�כ"4���h��B��i�$�ôcy&D�_�\2���-�eG!Ζ�I�_+�ԏ`�,㹐�Q-f���ܗW+�j�Q�����*)�R�IfӸ�r�eu�4*Rnf�Br ��0��3 �.���q�*C��F{qf�����[OY��=%6��e�m[��^A�$�!�O(ˈ����ViI����3*�wd�ݮ�}d��G�m����mf�̨ �v`�AF��yco{I����:c�5�;�Xދ��]���ތ�8p�Ç8p�Ç8h�G8p�B�
(p�G8p�Æ�8p�Å�81Ç'qȎ�=����ں��#t(����Ҷ�;\z]�R��W�쬜�Qrw�������1%�-E]���i<��M�H�xvRj���r9P�\��׎�{/�U��ޙiRޤ{�*��9U��k�'p�|��V\�l��Δ8.����H��
�v���J�z��.ή�UAS���J)�/�q�A-XA}�m�R�*� rY�����J4�N��ÎL܅�Y�����
Ug(>̨���tA
Yq-�M�:�H�����t���3xR�r�ȅq��o���Ҏ^8;}\	&�=N��|��s���t���l�W�js�a��Ux��{��W��t3�-�B��}��;� 2�M�n��Y����$W%G2�̙�H�8:z��_c�˰kB4Գ:+䕍���5hvl�������"�P�m��f�YIڇ����V�Z�]Z0Θg��R�B��fk�!�ݠ�e��Oi.�[gv��&�8��Z")�5�͆�V��Z[5�y\�}`� 	�vڽ\wB�wu�s�vv���h|�x"�2���s�3+�X�2c6�]t����y`c����X��Aϩ������v�="΀�i���.���hF��"Tb'�H���"��]ݣ�}�B��!|���c�m|h�3h�"�t�i���
GE�Xr�n�����'T�W�K���$�Eeif���1�5�b1r�����6�_M�����j��֍�$�UG��vkO�J�:uV:�s9�٣R-��������J�%]w���ra��a�7;�h�5���GJm\��>����͚Y�x[cj�d�Cmކ���|֥�j	�֓ �(fш�wtA�Ҫ�����ݣv\T�ؒ��8�j�_	�a�r��}Y�*�vpT�r�L�'%]��Z��!���'2Ӽ<�#3��o�)z�l*�qyM��791�%K*H�{�,���s+�[Npf�P�EW9�;C�u�i�a���}k1�ԷQ:(r�˚�f�~��܁��E�g{�,����eʼ0��k4��}�j�ݒ��k4ގ�H�qSo��i�BS�:��T�@ÂD��&k.���|ZǗ�s����w�~�77�ʄ61����Ş�l+���p�v��iV���v��#��a��3Q/6]�a��Z�����3q��B3w�k7`��+AV���4a��"�_�ݎpO��<�:�2�!�MG7����	ш�Ҳa/�  ��\�\8�Y�����ҝGۥ�����PR�ӽ#
'�RGf	3`7Ky��|�|��'�}~�f^�x�+���;��4gT[K�Z������r�*8)��@��RYq������J^� �Jl�Vs1Ѩ������OG����ޛWנ3��g���L�<���ob�'*��X��+ޘ�s	{gsQ��Xh@�M�#o��}ߎ���L�x7���h+�t��X!#5R�	���A��7[�y�i_IAVڳ��Y��c��u�t12h:�^�șe�rQ쪻ٜ�ٻ����-n�*ɩӥ�t��p"��٢��r�b�p�E�So4�$��}.a�U;���.�]&�&��j�)q-�^YBAm?�#�{�x�k��y[���	2c���b��%�7�I�۱@�c���Mj=\$+r��Y�-.��Z�j�R}}�q_*�P[�������<ZPL��ux�{�
��n�~u�T��q�sa$KEEu�8��˃��1a&���ݜK��.*���l[��F"�Q�P�7�*��μW�{*1t���;�1v.���mifa4�L�^�V2���Kn�BmT% ZH��=�����δ 
M>2�i�&���M��wa��u�7u��(po�uKNVV��(>�;Jqd;qj�5�PWKqy+���M�|/���Ա"�n�N<ں��7P�lj����b0�׹"D�<���ޠ�S�|[����s��G��6��3ۖ,�2��}�0z7 C�.�ώc���b)M\/[%4m�B�G�M4Nc�ٵHhJ�A����bDف$��/+"�Z@��Q	!ڨ�u!��[�B�.�w����9�v	���H���9�ъ�m4Z�34�ͬ�g5�4Qo9ʊ	�8p��~���Q4�V1�lki��Er�j�ح��h98r�����X�j��D�F���zzz{W�ڰm�;Ð�r��Z�lN���"�����4A4Ĕƌc���}==�M�" ��钍jcmL[b���ەɶ�v�X�*�Ɏb���AQ:t���z��$}9�A�c��`��6�!��G�$rl��l���i$����-�9<�pv8t�������v<��E�
b����7�ŴE��Es�fJ,o�o�*"�V��9���lΌs�mb,gD樠���?����m�լm�kfŔ��S��c�9�m�?#W���.�Zl,IM�F�5�sg�s�SV1d*�ǈ^y���b��F���`y�q-��&��G���?O��o��'�1���8r��p�.Y���9<yZ5�����snS�EU��ǔp[m�71��km!�rc�c�T�s��Ä}ǆ�y����ӧ�߫�Z���ǕO>�s��g�*-h(�n�xc���-rۏ9r��ハ�U�b�Z3��m�����ܹ�Xt�&����m�$���&17��s��8r�kTX6"��r����c��˕kr�u�$M�"A(6�ߴ��Ps��1���?��t���[����Z�̛��.�''A�ѽt��5.��-�F���	%�h�D��fݒ�}:���ka �pO������
����Vky���s�?3W��p�Gq\������So}�����e�f�4�s��|�*A����s�dι~��{�ּ���-�L�h�� n��@9ۓǼ34-����{�w9�R~~i���zK�����q�� �9�ׯ�7`��'�:���ͭ�d�{Z�{}^������ke��f��x_
�j���vn���!O�H��%��z߾�M��o?tL�C�sF�P�+�����؉6��1�N��$𫼶 f1FO�y;�;ô������V�ʀ��%����Hrou�bO �w�G�[��粏��0)<�k�ON���k��+�W΋V����ٺ�]�
,��Gj��T<-z���n,����x$Wf9� ��4l�l����6}ѭe�1��1�겮���1gÞ�%�y�����I�c���^mÎ_T �����n��>\�Kŏo!6�9X�?�۫m&^�A��@��hSn�z�F��V6�����+'"��Oi��/y��9�6�K�Q�Q@,i�I7�S�w't��-���F���\b67�E��d��}��Z���=U�F�糡�`�j�ȁ�d\�y��ށ e�o���D��ޘ8$�~�Y&#t��$���o0�>�ft}y����	�i³�G�7�|F��p����X8��up�U�ܒ�A}^�_;�����5y�%���{�I+���I,ԭ�xuz��{~�k,u
�� W%N��=31�՛��*��y�����ۼ����M9K����];=d�8���HFgZ~��ʺ;C��GK�%�1�A�82��Ƨ���77���=�]���R��t1w-�⻫p�g��M�=2�^�����m��p$�{�ŏޘ��@;�n�]@6������w3�sw��K�_z�4���6�F}N�W�?b���]��L+���T'�{��Ax����s���t��"��u~��y�}3���]�:����F";b�B5LUvBB'oi�]�/��K��l�9v`��[ﺺ�ܭ�f�"3�v�v�E�KU�9����`:�7f�����8D[B�9�AY���@��t�3�dtt�.DD.���l�pGv���]��ckqY�ۨtW9���K��)r�o�+���Z��oǬ70���OU���I�c%�K�4�z�ٞR7�PDb����������s�Rzx׃�".��=��n��b��N�_Y��������~�t�}�x_�׺V����B�=����zd4�d՛����u�oϮ�B⼿]9��f;�"lPlӯ:��;�6�NI�֖������	��ˍWJ6*l�<�i���U�I�rΪ��ws�dC��m�Syw��4&!����U�Nә�D	��l<2w4�3p&�O�a2.�_fS'���Ta�9�n��ͷ���{�U�{�x���ߎAԫmPB
���Qr����=Һ�W9G�}WdӬ��P�5zne��Pc}P����{,%[�U<�u���
R.v!�ئg�T�=ڹH��ו����D=�JXj���X{�Ė�9 o��It�[���l
�c++�B�!�e��kb�(A��לP����)>.	���]uf%�GDV�HH���F�}�3b4���ٝ�}�8�����x4�-��0�mp��VN k�87;��Z�7����,��=9 ���c ߝg�M��yD��y���=ԟ�'�PwE����Ou�븋w�}��x��jx׸���O0�U�]�o�x�>��C&G0��N�����P�CO������^}<�����z�73�f��aM�~���s��e|&��1�r��Hk��\����7��1ŉ:F�l<���j�Kd���|�>a��M����/�~��sȟ�G��P��k�=�X���z�`���Y����ɥ]asޝqv�߼7�w����G�ςլ��vD՚'����a�M�Wx&��]Wq��_�٪{�n��Ƭ�����s8�f���0���O��g0²{�kOe����,OHE6O�֡����N�^3�oշS�9��N�\���n���yQ�ٽ����������9�8�-�Ϻ��u;)gۦIg�t)�N�$��"�˃=S�o2+�L��1S�E,�P=<�a�=}�`�a����F*�*�v;�2�H���"�e�z��wd�GWofb��w�Y�)��t��~�)o��߮�|�P����@�ы�C����y��v�?|+��}{s�]"�#y��5;�ڋvF%�g,�^�x`�E���x|P;�����'�<���?l�o����[e����!�����#��u�=x/hHsj����T*}��߳{�ҥ�ך������9�s5���{�\��b8Ѝ4�]��3��C|K6�X��_	�y�y������̗�g��/+����}O�e>�&�Wz�u޹N�3�c���exzq�g5G���S|�NR�'��O"�����Y�}&^{�U��"��c��@��>��݃r+ۤ�=l�y/��9��b][���zze"��� 4���T��ٯu*~�����e�$��u����}�X|X� 7yp��xb�ژ��
r�!g;��������m� *�����-6���%^�c�2hn�&�|l�נ����|�e��'X�n�@U����|B�H����V��m]cu��*��S,���m�ۼ��	>��W�ZT�����r���gc�S�9b�����YW�j�Vk�]
6;�<Ƅy�ū�U���F���8��5���.�������4�Q�4u�:��jw�b�CU��E��g�S�w0�����~��zz}�h��&�n���-s�{�>���׵���R�%{:�7�Ͻ����������crF����
8#_��8�x�ם��U���̫�{���3�r����¥!�Ʒ3�#� �����P���Uf? ��x�/Ou?Y�Z��~��q�<�޷��5�ѹ>N�r�/-�ە;��l��o���n�d�x��_�s��?5�+[Sw*�5o_�`�*�=_mc^߲��@Y�D�#<�<缮�_^Վ>��7��'~5r�Im>2����k�ǴF�Iw�������7_[�j��Y�k���_�}��9Ik�3�ٳL�\��=ܡ;�~����aܕx��ޥ��2���l�F�0/�L�o�}�&m6}n��������U�{˜�Sޤ}�Kj�d�}�C�:r��\;ޣ}A��1�j7u||r��иc��R����5�u�7b��d.{���8Y��NJ��fY�[YC`�/��2���:�We�Y��*Qo�>��\���o�l��՞��w��m�3&���l�uwս�R��.�s e=��!����;ŕ�g���Uz�珩�K�x�x��jѧǢ��NNQ7�C��;-���j��Yx���dd�M����dwN��vOQ���]��9�#6�v��ґ�R�v���pS��6�I��-Gp.˾i�g���w^�7y�����Ҹ��އ�>ш.g8ğ�ء`�bW�^Ze��7�Cs���|�}�G��'}V/�������rc3~�����~����Z/3L�q� �r��Zlb"�e�;]ѕ'�w:��,�����3��ǀ�Sb<��'��@�Ή���$������;�^�i�N1���_o@�L��_�:	�zr���o�O��Z�����93����*Z���Ĉ�5���4"��} �����b�-�G$�i�:~��������N��Q�X�~/=G=4d�7>��Rq��[�q:t�ƍbR��w1���r�)V�ZVH�N�)�m��9�ofH9�&�\���W�7�4S���S�EiP��P��2^onn�ok��(��6�@�W\🊫���e�c�κ!,���w��:�@tK����K�b��U-íI&,N�V{�)s��hg{io�8�_m����7��5|�!H��֏��%L��=B�Z��*O*�����1c����ŏ�	n���~����˻w=cfJ�Py>�(����2Pz�D����Rrݫ�/�T��8{�nQ�{�(�;�[�ymg�=Z���y���^��%6�����ߗ9�R����z�4�Nf����e��T3�%�H�{�ɕ@�}^��� �@c���S���ޯ轝�Ot=<��({e�~kL�]�fͰ�8=�m��̏Tc"6��gh��,�a0.�m��Ƒy���g�񓳚K���Ƭ-Y$�i�\�#£:|���缺{���u�3�{�E�c��=�jN��g���\Tz��u>��vm^��F>ʹ�1�}&<�w�{�evC$T��Uv�)Q2��>�W�a��{ީ���y[��=�,6�%���֓aU�ͻ�������T��D�wl,��:�!;��'<-��yK�������w}L%�4��d�)��h1al�+��{��cX���wz��N����!-�g���,���s#Itr��Ov��f���{�����������6��Y0��:�5`��2)��|{r&�����g��s� �C�L�uw�G��F�q�Ic#�z��q��;vJ��տJ7���0d�Rj�(����E����[��{T�M�b?Di�{�zgz���|0���7Fva�d��)W���u͟�#��}�A;���'��F���U֥�5�R��J�Jʲ����7�^��Y�Ḵy�A� e�A�7�R
ڕ9�젧�,U�n)�=^�~����h7h���<z2�D�g�.GH�^��a1}y�g	��6y�w����s`�ӂ�������/����+Ʋ{���
���:Rw+��՟O�~#����'�����~Ă��F�u]�N��wf�nz���'����~�L�u�H;n�e�ں+bKd�K�����X�V�۔�B;�n�����A�8vt�{`[���]�|��;��ut��T $�lFk�h�ON�y6����X �GX{�g(��{��Q'�gi�p0�����dz�cjdy��6�={zٲ����1Թ�wh��;/6ދ���/���']TU#¸�>��;l�v�n�N:Aw�ϱż��g�n��n�w5�Tu����|�����b�]�垧Mמ�����!�>��oQ�$Jf�*�����2�#=m}��~�tgcs�����-;�I4I�l�U���[�X�u�3�����@N�R��#�[����ٝWn/U��s"O�+}�14�C�d}Y=kJ��$����>>r�����V՞�^��4�h�û�S�L���3����{};�߱>}v���k�(-����ϟt���������1�Q[<|�aR9i;�V]ߪ��U���{(��WYGо������J�����)ח<a��$zFU^-����{b��5�u)ا��V&Av�^�s�J��;ކ\T�G?YC=^�k�K�J��Bܼ�צ�>���{�����3Ǉw_rNF�<� ��4gx��XJ!`���~ ?c$��c�6�<�.~u�NS��j'�4�h�8���f�̤c���dp����@��˻���*T��)Մ��ܥڴ���!)�k��.P��|���/S���.��<�M`�Tk�@��t��¹̪;#�; B��7�d�ጶ+:�7��T��;:l�֧��J���5���ڌs�����}s�GE�\O
��{��[Wߛbż���ma{��M�O/8�t��!�u�z�X$ۣa�`�Ѭ�Hk(����<�;]���zRz�a�Եt�i��tք��d�e��͆ �$Cpm�ה�]��Yo�C.}0��+kv<�$5��[��o[�R�R��E�>|�s�V�����ǻq���s�=�q�S��}���0t�S�E�&l���� ��Tn���ɩ�`Ҕ��/&�0aO�����L���c���ţ1�vB�(��,]sG+T�M�r�j�)�0E
�)N�u���>j�ڢ�+���� ����(�u�������i9��d��\|upt�G�|��$���3"�Z^-��w}	�ڿ�S���fgTͧtt9ywc�ɘ�[̮�sqҤc��9h��bp�Z���j��#�D��YRn��f �j�Y��e�:O(Ӻ�}�W�r��KN����\��Y]�:�z�KUooN�E�9E���/4b��}�w|z�W{tPN��A�TL�o�f$;��c�!%cщO΂�,����3nr�v�m:��L�JA�,g��������FΚ(weu����d] �ͨ��-�{v�M�8d�,:Qv0�)wsЗѻ�&�.](�6��]��Cz�Y�g�P����bJ�έȻUt��n���lW�Ɣƹ�Zǌ�D���?M��+X��Sw<:��`�9��G
Ы%�����-�5��.�{g��&O���Jj�R��\��/nӥ8U�"3l��d^����fi��;D�����H낳s�J�
(�˧:�!����4K�͒ �.v�Z�ݩ�$�t3��c
�*���9�W������P���J�$�l+u����s0v#��,���ji��%�-�.�!7�m�fYU�)��.b$:���Ŝ2�������6WUm�h�/��LbH4���.��\������v�Y.�����Ŵ�M��A�$s�[���N���7dz8o;-!VŶ��Juf3kiP���D��ū8��1�
�������v���F��oo��w��'��ڝ�ɘ]�HWF���v�Z��r�Q�%b�@��b��I`�ݐ0>�hZ�<�{�'N]���$�-K��7�sݓ��$��%�P�n��8�lC��2�ntd>\Mq���"��kL�i��Vr�
�q���눱r�zu���p���t�N]ҙ�#;�X\�
Y�U�u5{�uu~2�$ 
�����H	!h����uǇPPm������L��͐@'�$�(`���+�I�M"B0�ZE�i��͢墪��[V�s�ss1^cy�W���^.mi�O����MJ��O#U��U�P^sr�"*b�Ø�Q[��Z5������ ���r�6�j�b
�y��kZh�3\�8�kcm��L\�L�����z|��|��l�U�r�M?cs:"��j�����M���ED[j#V���nX��������"+ېk�l��u<��L1DE[�ق��i+��VM������*����#҈���"
��b�5b*��;SEPF���M��D�Q�cq��m�#O�����m���xsb�o�b����kUg��ɮ�ᶴ���k�5��V5DG�A�	刭h$��}?����{���+cU�l�F�U�E5O�<��T�و���*�j��fj�?d�PDs��4lA�j �����kX��	���ѹ划�*���B�����>��D�\��F�7M93bۄlWBN�Λ������Vo.i]��E�=F�w�  �Yy|�#}4�o�f����+�$c�ֿt!>�	���+Ю���8B��(�3�,����{f����{������^���C/N��z��HJo����A�<7L�g����mZ@�%M�@��'k���)s���O�tჹ��XT��>&r1����	�oվ�����-�^|��{M�oEx%$6�����ǻA:�����M�9��/E��謨ס�N��<	���@�����/�oB�uJS^�ze��#&���mg}7;|�.`��������T7�!uJ��W�x2>��Ɯ���F�T���:��G�cqF�ڧ�O���J¬��������j٦M�L��W������L�H�"l�����/����#����DW]�����G�X�+H���������6qSx��g!��A�e�O�\�^Z$��j�Ս㻗r��{lo(�m�`�҃a~`�-pC��Z�T[���B������z��q!���oS�k.w0��W?�C����.����l&�9��VrW-`�EE`�2��O}�PE��0�m��v�bk�f�{ߣ��H�ߑ�o�F�*����o�=\���w9T�P&Qt������<������<���ъ��a\�fEI�>w2�ɳ0�i
��l��GD����	ٕ��ǆ79�  roZ��u����B�����OT��mSڲxT�e��[s���E���QV�ʴ%:�=������r��ۗ������Պ朜�ޞw�0������
����8la�N�A�K�s���*	��@(�����F]r����9���}�\~�444>���F�>Co���L�_T`��.�ȱ�tkV��/z(H�a�t���E��;<О����&��5���6?dG��<��X���CR�uS��t�֠%��Y	p-Ɣ�n>�N�#"�E*B	��������T+	�2cW_j��C����ݚ�:���o�Kd^��q����n�8�0�fˋ8"*Rb;ۙv;�^��P��{TK4�ar���~���f�������x���K�%!��;�������/�V�YοL�y�Q-� ��!���MUza	�9���r�<����-vǩ`��d77�#P�̽:���!�O3s�U�%];?(�C�6(�yן=�P����SS�X�2�ƮO��g=�F� �S6�gd�2���O}b
?{���Κg��#��l���v�nvR4r5!m}�-
�u�٩�q�_5��2磑E��[B���G���iw*kޙޛ���$庭��`ghh��,sW�T�����aa�yN:�?��u��,����;/���I�#w.`�#��؝+��\�TA�Lܶ��v�BR:�ƣוm�G���3�R�Iއ����|'|oth�k����x(����G��.����6;-��A`�ł迧�"����&5����-�y�"��)�p�{`��qo�c7�0����B"�i�T0\aۺ�=d w�i��{�	���u�������x�϶�.O'g���=x֢�NT^��ٴ2��(+
N\��þ�i�"BM�Cy�HA��3V��v�:�4W9f��|��6���F���)�?g���U���$��Ǩs�e�<F4�t˞��hǔ�V=�13T&v�ݎ�-d:*L�z�uR�����28����k��(���:�^��!�-���#g%f�,��מڷ�-�܂�^l�Uㆌ�9Jy����I�s[o�@���h�c7.����daq�ӯ��_<�)��-�1���{����0�Pd�}�	�֣�sJĖ������!?y�;��{���8���6(1i��~����z���}%�=ܕ�Ĥ��z����r:�o���i�ýv�-c9��<(�>�~�Q�DR��<]k���W㿵�<�tb�]��?�v;�4��1AAgן�-�lK�}.	�����Ʌ���>T"$x��a���Kw�_3�a�Т=n�9N��1j�L�il$N('s���9l��~,�eu%��U��n�Ч��ڷ'�s���N��+�2@��"I ٗs�]��>���4�ۘBv� k.�k�}M���{]ް�������B������s5��!�3J�3`�&�سmGN77�� jse�F�{�.1�)�/0��|�Z���`��ϐЎ����`�&�\^��<�K���u���ۻn9O��?tA�KH�৖�)�	����t��Bl���9�ڟ}�8gd���Gu�Bj-dX��R7v���z�?%��E�	���F�<�n�����s�L����xaG{�'@W�Vh<�i�G)u�"1+��6i�%\�Ʌx�Ec��?l�V+�ǽC�\K���*!��.���mm/�S�j��T"�@)��ǋH&Ug��C'��9*�F�|ك��9�S޽ J�l��YtP������C�?�;�[8��K�Ғ�b�	��k	�5z9	�����[}pю�$b�6��bsg�˟�]6�K.��OW02�uqA�Möd�L��n�fmr����ݙe����#w=��%�d��U)��*����u��$�C�;�!����*P�ػ[��!�{YzlAn�d`dӆ`�t����g�Dz��_���6�R���~� �ޒ�\�޳.2�^��EÁ:�?�'�0��s������������@�^��A.�R;]���������m�_]L�@mGo�dv���͚�dF��v�.�s���H���3,A;�u
�q���/��A�`�s�3��#B�S�N�G������/�D͹J��S��kSx4����J���ÍGŦ�2K��#+�a�0 �_v嘓=}ML�ώ��� ��������W��2�Xl��g�ば��2��f����g1oL"���~Z{4g No�cA�t���$0F�x�Λy������LS��nΗj�l�u<��:�Ӗ��`�����=_2�������@u��?~F3��j~�\�9GMlͫ�x;���8)�aI��=��(�b���H&�������D3lPXY���:�V܌m�/ܨ�0������a��������U&�Z��;����ufx���jŋܙ��uc�o)���V���V܃\&��q��z��#�͔j��f�N��m�x���P(�����Q��xh`dm�mﻳ��=�I��ߵ~�a��g *�3����c���͕�.�7��e��fݵ�hd� ��2�������H��>����C��O�"�ah;}���qv�A��Ħ������ ��62��{oO<f�ׅ��ͯ@��m��8�L���I_ʃXFނ�<���|�8�4�F�%�'��wN�C�I׼����ȖMZ�mS{o�ek]�S��׮�yJʯ�D�\��g�~�=�w��&+��I�QyD��ڰ��	;,T~�Yu��]�;�$�8�t�m�R[��-��pJT��G{Y���w�U�{ܪy+���Mۣ�R�[�Y2�^hV*]&^LQ>���y�ir�ӻ����x�/`��;KI�7���n������'�?W����^�Ȃϓ֊��;�s�"�~����
b��d
l�����S����zt�vV(�)��sn�u�B�;m�e����'��2�����B��2��5����M�sU�tn�f����o���F��#��~�PY�_O���J�,��Q����og�F|k��Z�u��B���$���a��L�!�\�x\�'���vM9����U��6i�n}�k|'��;�wk�S���e�� �:�O��q���ç㾩ÚK��k���4S�w�9L�2�&����-I��7Qe��}Z)�������y�so*<I㨈�Y�jF��y��aE	JEU�gg��b�����{�Fkg��x�/���w�U�k����o*��止�pقැ�TcN�F�\�%�a�F�5xZ��Uk׉��Q����,�V�t:bϬ�ٮ��|�d��kY�V�ΏvϷU������rc�J�ZX+3�wX���߉�ÊTp/
��֯����A0u5��Y�s�_�b�%�ϳ'ۦ1��9���Ih{�S����������p\�D&�w�.�Cw�~��͚@��w�(��ٮ

�X6e���{�f̾�q�^Jd���7��6�춏b��}u�N�T�jR�4<����+�^⭀eu�3�8�2���+�ț��%�bC�4����M:���ك��8����hi&皁�����.�i�N��Ƀ��v{��`d]��e�AuF%�!�:f^�3�L�f�%���*��w����O��ޖ�Z���n�Orϣ�q�43H���b�s]����S�@>��z�l ���iZ�0�wYޖ�=��U����K�g��fT-nڭ
Q�ی�"{�2b�O��U�5� �RԽ�E�,�'7��Պ�k��[��;X������Yn���ð�k��s��y�墿eO����n�#?wDȿ�f��NwԺ���CIqo�<�r�f�OGL*�Pr������=��i�����L�F9f�S�lc������m��a��n�	�������W�m U�a�k�H��E����c��D,��_�!�*���H40w��
�m�������LdU��НT����,��(�%g,�2�9C�h��0l]��V"�����w1Ͳ�\�[��cz|�A�
`�]Z2{�Z`,�&)��$�k�{����j��8z�b�OZ���f����g'�Sj�Ƚ{S�
��B��dÉ7j��/�G��d��9��d=��.$3�=�e���?�;lt/U�>�Ӵ��vi��4�mo��6W�fwU���o�_B����AJ\:+Il�׌�p��e�st+e<)[�o52�fS]�c�;�N�ɶ둞��m� �ͱ�r[�y��<!+�fDJ�����Hkbu����<��*"��Q�}� �S~����a> ���	��?7�s���U�L99�AͨOVc��8�%^,�C8�v�JΝx3���d�x;����� ��|�\F���]s�[��Uy�7�%=��:�=��N$b�n2��h�P���b[oG��=~��}6��L��6�7�/Y���澖�2�)P���n�\<�P�§��˘���w�~�߅�*���-�[8^��?0��%��s-�͹Ւ��ǢS�i->�灉��� c5��QR���KD?��y��;:��h�I�I�����C�i�+�u�TF�rw籑7���`���)�	��c��M�HSU�k��`aT�1@� k}��n��þXk��
2��0��4;"�V��!��e��\�5��2�����0�j�(S4O��w������\sT�S\�UM�y�Jh��mʷ�S��e>������:���<���쨅9R_��fͅ�K(������n~���=XZ�w��Zkܰ�,:�K����x���f���@�om��l]⑍�o�랝�u��X�½V��<Y�A]4�SnA��㝔]Y��s�L�)N��\)��sS<;N�����ŭO,S쒸k���rd�^=E�o��KL��R��G�p���]�
yQ�H���7݆�f���WBY��n�����UT:�I�]D�9ަ��Cze7��UL��(�7X;u�J�å�{2z��������(��d��M{�{������t��q�K���It�����
}M��rq����l��\M��r�Ҏ������ݙ��2}��l��I��d��&C��4��~sJ�uQ�Y6����Ֆ�R�%�E���,�2?��9E?�h������>�-S��^�^�v�4ٕ\��Apc��Č���%}��&�����=?��t�1����Ȱ~
*jTO����;���5؍M�x�ג{#h��Fނ�q�GB	F�[�PZBֹv�0��ƃK�X.�#ϾT"��hu:<n��)'l��i6�G:��Ȭ�Ǆz�)�9��dZ�3T�:��E˱�A�[� kC���>lj�v�
�SƞD�:b�N����d;f��Odǲ��2׍��~��K�u}��w+��FeT	��Y�[�����yYP/����mGUs)^�� ��`�Qs�1a��`�06�DͿ�Ow+W2���Q61ag�{'ƄC
��f�5�`;Gu�f�/ ���,l���M\�k�
2��0<⣟�0���%R��ܭ�5��5r�t�l؆��nPR�]��LG�]�챼ɠ/�y�/>�|>��պh�b,V%L38��3�W[����)��.�(�7�ä����*�y�_͕�K�§պ8K���~�:}�]��r�����OQ-1&r~L��yl�v�Wr略��_�/$<�^��p����u�l&4E��b� �C�?�:p`o�-
�w���ܧ�F����&��Z�o4�8����mO����<�-�x7�H��g���*J�I��u�2E5Ջv������Kw+y����ZY�\�K:�[�Ed�aK=Z�z�!��2�f�r��ޥ[[t���C��wk��A�=��[��N��&m:́-s���]�U���5y:�h]G*eGou�b��A�Ϧ)���;m�0f�:�<��&�r���'T��z�cS6{'K2�.{z�+��0��Qr���]�ay4�˲}W���4Yڎr���q��d��x���&5[��R�ޭ U�^X��X�YbZ���h���>e{S?�m3�+�SG���:J��g���9���f�s�y���>m�����lq��g����5�x�z�h��Տ����Ӓ�	i�ܪ�{P����� �3�T�M�;%�����dX7�0;� fw�4I�m���	_��d���]vU˥�ҵ��	ᭊ�Ö��#��JS;"��}�*d�H1��n�u����y�g�8.ugtS{,�I�˸�(c�y�ۑ$7�fh��l��:V��8��v�;n�]����'}��	yo=�aW����2Y����l�t�k��f����4�lT�L=��;��w3Kvue�cLa,uI�݃J�]��IbRc+�%�6��䰼�9�襓OM�ȳ��`�X��(OoS���o�ɧ�91���|���#��ջ�mΎ��=y$�E!�z��q�#��m��d�8��2f�w#�+�c�P4F����!�]vS��^:Pj$q'������u������ְ�9
r.��)����:�twvDK�xe�Z���Uf�h�;b�F��m�'��-p�a���&��DM@�D	�sUr\�'�k�!��ٯ:m��實� ����r���s�Z�\@�/�䠠-�Wv��[�oM�/���y8ChΔB3[ov�U-4�Q�������f�:�$�N�/���h}z�'M]�z�K�n�\(�/���(_U�2p��.�e� �H&"��r��7wwqC��c�)�*񺬝�������q�nk�'S8f��$n��d����C���G;��fkS��Yk �QQ���s��aFԓ"���րqp���K�W0���ζ٤�6æX�j�е�%�Q��U�C8Qދoom��L���ִGQۗ���ur$n� �H��Ġ�U�Q�)MD3��,Z�3m���� �*�N�U�6"�_`w�)����&��͆����F�/u�����i�T�L�6N���L�н�e&��n��s8�j�i��ͦb
�ԭ�՗��+����,MMs��k]��R�'ѻ�u���5r�k��*�N����.}��a�k&87i��4V�hFC�,�SP��l�l��Sgq�������Y���Z�K�#�&��;��,�ΰ����ԧ��Т*"�tD�뵄�j�QX�5�݋���pX�_���i�
�n�e�\;0N�xr)�jj��X02Uը����}�X�}�/��(^>;�ɴ�B���2�n�,�-pB�<��u^��ֺ	Z��v�Dx�:�aD�O��k��a9�����j��8�F��@Y��]��y���:$�h|�1iQe�h��ۤ��q���
)�t]d�o��䓢��J��@)c6<�V�Fǰ�z��p��t띛�5��e�R�v��m]%8.4.���"uuL�9ʶ�q4U��Q�Ҭ�ɉ8nm-��B�bK1J뮩�պ5qE�:ܸB���u�<;V��!4�8G��="��צ��Ý��w@�I�%�ѩ;�c|����Ip�쮵#�����m"B;ilP]_�;���7�K�r��*ޑM�#�h"k񪄚&�AV	��w@�/5�nV��[.�+!5!.�(ŭ�Ԅ1�p�C�Q�څ�j{���� �$�Yt�N�Հ�5SE7ȬUEAT���ruD�[���h)i��������S1�{�g5m�6�.DSD��W���W3�b��������j��ѓ�:}==������"�y��RRAAD�'MTGѴQE�d�
��Tܢ�i`���ӧ��u5LU$�5I��xN9;Co�Ȭ9�Z���u��1LES���,EW����>�O����pV�N�H�?9�DU��$��7��/v�>dĕ5�ؚ�&��h���|?S�*/m-Q$�T��UVڂ����QUIQE�bj"
h)��#���}==(�h(9�~�Q}�U�b��5��1L�_6h��Mj�cT�\�1��t�=}��-TRI��5R�7#Ulj"�Z��=�˔_,U6��D~�8�h��?����S{�QT�E%�Q5PMUL�1PEQU��&"��KS$N�(�֒�"֛X���Pk�YxC� ���eIpG���,��&�b=�nQ�7��d��NJf�Ě8�8#��vr�P�nJ�W�@��$D��p�~~#��W�ܩ�����E1{ү(���ޯ��l��խ�=��4�a��pf���ڹu��ll��:�P1k3��6�!����\1^Ǥ���#y�t��O��C��ǔ��I�``�w�����{�3���XH6|Ɗ|�����/b��?��zl�G�;x�w�j���ɚ��0j��/����������LMy�cѹ9�b��*��͌�f!^���� ��J�L�|�c�{���i��w�}�F��W+CߌŴ'�����Ou�d1��OǇ�.�+Ǣ��o�aUe�}����N؟�pS�69�c4�����V	��|:|ܢa�_6E��ᢕ�6�:���U.�R�\[U���>���!�=�Pn�Ժ*�r���2�KKm ��]^���ܘ܊�����ꍧ�s�F#+_9�e}�f�� �D�#X���{���������I�Q&�ͮ��n�2��~��֜�}]�쨼&��Ls.{[��g�����`w�����#-�u���T0�wc��oG���O��A����+�ƃ���GU��^Fm��(�ܽI��y��/-}�	����Yc{M����fm|�༂�����h�'q�����Eo�^��q��k�}�{[3yH������q4�,�&�u.i��A�TD�E�\�ێi�Ly������:�j�Z�KpTQ>
��,O��	 �	�3��g�{ѩ=���3�I�-���*�o+��#8GC�f��K�З@�7>=a����rR~�ɩ���Y��oe�fB�u*{�P�)��L��	O�Y��L�LP��j[ ��\�v�p�n����V���D�*Q���i0�#R���)��(4[�B��=,�S�÷�ȃ�����/��u
��/�WR9�{לy�л�yŝ�E��FK%�������4M��9sR�5�]q�lݕ�μ�)����Ӗ�:(�i�T{�^�C�Q��� \j>z���Z�rf��:��kOm+ɢ�y�C���}c����	�}t锈�-��gqX9���_�q����5����В��ff[[��Ar]�q������d<��L$�}q,����Ӳt�M6�n���+23:�2�3��O�HqTY���AzĠ��݀�y`h�kނ ��$��.:r�p�n!	����-�1V�y�����=`c4�+B�XQr��@tK>��D{cN5��V=Ll�!�>����B�����~�k���Qc��w׿tt��`ԌE0k�6П}�f��/{9�e۲hb����ʶ�U+�u��/z��:r&��Z3:�uL�"s�{��eu9����Uޘr��6��T:�}W"a�ޔN�B9F���-��F�<�<%H��GT�'	gq��݋���f3���� Tř� ����p�f�;���-���$ "}36{�/&�˗�!פ@�w��)���������>?G��gE�G1��llL�ٽ"zڦ�����?dh��Xw��uoB\sU(�;je���������sK:��^M�<(�u���ߴ+,ne��O�0�@���l�M	��C췠�7ߑ��S?�~����3`�~�A�x}~a[%�0�Ue��YQ>�����BTlƻ�\�[�YVd��}�W~�&`XN�d�ܮa^��-*�: �;�g�r�Pr�� 6=��lO��c[z�,���\&:F'nB`c.z�A�Y������It��U�Mݞ�� ���2��՚�����-�}�����Z\��P���	�Y3a���,qniQO�
"��.~odeX��Ue;;���]u0�֟	�9��1N� �y�|�������?KR[����Ur}ӭ�	�$ʥ�!gL#�և�HZ��1���w��%�k��!�6�xT�l�Ԗ�7
�z�c��-�{;����ڭ��I���A����A�������*��yh�M�Z(������0�y��kY�ݤ{�%h��9��mЎM���['>�S���x�E��I�ze׎�Oj��%��ō��l.�q������Ѻ�Cw!���H ��Ccak���S,��9�b��2�ɱw�;��H�bkGZ���D�]�5�������A� ����iW�eۙs[9Ȗ�oI�Ih����ɑA���v4c��w���`���v�V��R�T�]K��/X��c`cH�����3�ǰz���O���`;>�l{8%�W��Q�Zі�&���b�G>ю��W�F�?H�ֱ�ӥ��e��x��*��۷��LO���v��V��i�CB�-�h���~J�X��F���ܱ^�s��W�?�&�n{�۟V��>o:���W�D���3�|��|����ޟ����^��{~�;_��E��1̫}�����h<�06 �5��i>�u	���SW�_
6�k⏿U�>�2��E��ض�B~���t�
�Ոvg��d�d��ῷ�H�3��}�SY��-� U�,r��2���w+��1�	���\ԍ�u8۝2jYɶ��u�v+�j��q�44ۆ�I����>�E�`�q�V܃vH5)٭8-��M �烏]�I�:��VȦ��Sx�筥O8!�����f�[�暥׸÷XW�E6k6�
!4����}���H�R��eWk����Sݖ�I�>�.l���aY��Wt:��&ɗ�z�	��{���1ͮ_!!�p�1�:KcH9W:m�4s��䰆�D}�hcAN��Y��]��Jʘ�º�8Է�xL��)�)T�[�j���ղ�:Ѐ��;m[#�7�>�ݽ+,�Ǒ��n	"�Q�����ıKD1$By��;�������]�V���o�a���C���xE�QM>��,�q��ݜ��?2��0I��ʅ�M����y=��wt �(�n{��K�r��4��/�͑L�Q����K���o�Wb��sR������j�����j�7$���=���F�W�Glq�XkO�l�R���0��ػ��q�gakV�Y�O�]
ם�B���r�4��Q��q��Ɗl|pz�ڿ~��*�~^�H~����<�!���^�姝�ņ��[��9�9�.�=�U� !�Ú[�n�㌟FKI;3�c���6Ag`���%�a�iO�4��펤�r0%���ድ����#Z�p�fXෞ�K�IN�r��A���8��$N������/�~�p�X�������-�/��E��[w�+%�����U�⍈r���F�:��6/��:b��\�0�c(�t#� �uW��}����w�xa�������Pߢ8��\���/�9D��LMP,2"k�D7:LZ(�H���u��hlef[�k�g\�,����%����B9�q�gl�C~u�m|�'�凞R�Ҹ|hm�lL��S����PV�T��2L5x&�`]چjUmL[��F�΂+"���&�]%�sյ2t���m�=Mj��v�kd��μ+AP�v���ޙd}�bj|�h6pfb���gKO�ܪ�d}�I��� y�x0o�0o{¦nГ�����%�[P����U^����%6�2!��KiN���ڙ�h�>��vWe�Wb������G�^��pCn\y1L'uJװ3�P�E'�+hV�n��D';��������m��DHY�����ԥ~_��gʍ��,�q��������"���֪���i��o�^��Q�{Anн�=��B�o�����p���cӍ$[&k�8ź1����u�6�j��ld�e�J|���/�z��啲��Rg� ��k���&����S���X��6i�{Th�{�ߦJu��s���!Y�X�1Qq���OA�1� s�mjoz�o1^��*i�R���<��0�>9ԘP&�)�|QR�����څ?>/BVN��w����vh���in���u׃��`�<�7�YE��T���,�\��"K$�9�x�/�7���͟������φ,E?�,�+��S0�(7�u�B�O*2�l�P�ʌ�eo�Fd�	MM����[�)�y��/�Y�oo����j�z��Nn��>�oL���
.������]ͼ鑾�ó������<WDM�r���8{J��;��Ur��L���ˏ!Rnj�U������7�����Vv�Kb��k.%A,��;���>�۞�һ���n��G$�J����b�o���$�j^aK.����m$F:��_uH� bX� "F$"9n�UH)��C?)Q�V���tj���q�h/E�3�O�بC��8nl�ws�m���V+�ܚ�ms�m5&u�uyI�/M:L�{e���jsb]��6�vmzt`hI�����>u��Ͻv���ߢ:�D���l�4��o�z�01�*��b���tK>����u��Z��7��c���xߠpN�y
���|�j:��D�[��ߟ w!�|KH"ASl-��E�]v��7��b�9kK�3���{�Y���ME������ڦ�{�,a�rθ5�9�1?�L�v��Կm2i*�p�z�F�x���|5OE���-TC�@*)�DbWm��]��f�=ي�E�����4"Ы�s	e
ǵ��*�eD<��XbVl��m�u�>��}�ǚ���}�g��9��m�3l���~��i�_�է�c�ݿ�v�k�|��D�F�>{Uj[��N�^>�Ƕ�;��4��:�ఞ��p��E���u6���6`VkE'p���uf\ut��
�;.Y.�B`e�C�>𑏲}��ߟ�K�
�M��@	\6����l�9|�b^n�����k$���8=�;�奭��Ue+�+0֣>׉K�Ws3�l$�ֹ]�΍z�1\6qݳ���~F�XLR���pN"�|���Ew�
�=�Ji�]g��ݨs�v���1�i���+z�d��{������ww�{����!"%bF ��!W������~��Ͻ�!ST���ڧ���4�;SP�vd�L��.�))�(�O̲+�Sݝz���Z����SZ�k��0��@��.�Z9�_�dKjE���#���f]z�e\��b����W�z����x�k`&��l0m�-pn^9��"�nqb�E6޳[>�w8�F.����3�d*kd
S*�d(�1��c!Ai��q���@��X]�!��,��k>~����)�f���p݋��\���Ő��L��)�(�{�>f��[��v8v\3��!�݇�<d#C��v�e�t�9���ױ�=Z@��:��&}��z暚��r���%�:d�c�2��#m}Ƹ1���6�Z�D��z(
<���Ƕ��MWN�f/ }�iԃ��,��1K+���.{T]1a���nL�A�d�?M��C
*�f�>̠��˥Y��`�y�ȶ<��?S����0`�u�?}*��r�i��g?B��2%)M�Ƴݵꇼ���rN]��
���i�̄�=f]��x6���4�jF�Ӓ�屮	��)����͸y<F�OjO���7�<�x]z�J��P�դM�|�W,`Q��gP:�ސ;�z�Rc�D+z�T�L�"��?���ZD��k��φTk���F��N�)�IZy+��*%�����'�K���_h�Ѽ[�i������=�>lןO8^X�y������!X�b�R$H�"�P?�s����������Ǿ���3���z��}�O���r��iy�n~�I_Ȋ��|�}��OK�K�q���κ�8Oe�Kђ)���.jB�1+^�t ɨ,���V�6�YZת.��[6DH̼��۽�?ZɆ�k�>�k�Ͷ<_�FB�%c��N��.�Nyt�l�/�&�v;;Evl�e��CVh����vWA�Ϧ)���v�-F�mPyƇ�4����ڧ	O�5�[��bg�k�%"�\�l=s��v=Y@<c�5z��m�����Gk�=��/�w���9��}���h^�F��� �ʵ�!��(�i�/h����+ܰ���ʒ||�Z�·�c��Z�Zف}�M����.�'�w(�?F�ג�u��L�hg���[ ��~R�e����V�k���/:��H��j�����˔Ҟ�(����3���~��~����A��Ցu]Fm�i:�03�����a0��I�	y�&�VXa�@�7OYa�69�=[>{&y���-����������~,�ް���xK<�*����7,E��dv7AN3�41�,�{�K���T�D�T~[­�V�a�WM��^��2{p��:��s#&5ܾ�C9�<������Mڼ�Wp�!Apm_�-"�!�7tDgM�l��r����{!�/��l'��Nm�|��h�3ۏ� *V�U�W/�L�P�P4���y��h����?�ĈD(D*D
E�xy�x=�o  �9d�(h�Z����T�=��_-�p�$N�a�.Z�	���c��#u]74̾5q�����s}�-�H(�w�O
fb(�����T9D����:�����������������8Ȝ�L�ҽ�}���]�õ����b�-	�gEUUс�H�`�"L�Jj�w폯S��t���qN"ZˡX#�2��g���#yfגZ5�J�r(��{��j�ݯQ�YƟ���A�Ⱥ�+���S]8Gwk��>��a��,ii�@.��q�a�I�#x�oN��<��:����G��ŉ���b���c.�ZR��=����
�V�]k5!�tn�#�WC���ڧ����hn��s
lꈇ�P�>6`g6�nL�yOו4���p�ݼ������r~f���W6㤔�s��C^�UX\]��["�b�a��gN<"��1a5ۆ[���k��(B��ե�2z���;�:����țl^=��6�elXu!l1�z,Y������2fW?��f/��c�eN�O۝%��|��".���j�t60��Gz���z�����%{�!��EF���ug<��U� ᅐ�#��*O�k\[ə��S�v��A0�Ꚏt�L)Gʜ$ۮܦݼ�8!��)l�����Vr�*Hv���zka��k��|B�ʌ�U��B�T�!5V�wuo���H�QЏY�����<{�Շ2�VїȋX(Û��7���7E@@
�X<0˫��at�p����� �[����Z��x^�9�[}�x��P�Q䱝��vq���xoȸM��noc��ke�SE��kŝ�Jg��\|9�C�s:� ݾ\�+"A'�����ˡ���B��q�wz�~������n�Uz�Y�+��[X�����u��K�֦�1Չ�,d�êՐ��E�Ԧ��^u�}�K�C<v2�	Zu]��F�V*ݎT���]M᭗�pl]ˠx�8�� �(����8�=9��Pα|]�N��4<�FWh�mEe�;����+����'c��UP�#�4�'�H5�3e��e��٘&P�io*����f7�z���')buX6c��ƑSoP�k��=ӥ~�>��;/MI�P��\N-���:�e��'H*�*E�0%��	�I�ݽn�Ί�.��"����6�:�g�����,�{+�O,�giD�:���O�Ew%����1r�u�=Ek��I���Ѷ����nI�s����X�m�1)Ϯ���=�`����洨�^�Ꙧ�7.�em�dJW��[7�jҰ�Q�i����{�L�"�Zq�TB�we���h�w{OP��{�ќ���˂
j��Wt^P�6s��Q*[��xM�roz�_^��%|��;�2�yGN��|�Ynс���"��n�$���=xz��z��I�������$t3�:H��m�(��k]�G�S�ĝJ�&]�\L�CH��;���m��C]#���c��|��� ǲnR�gr�^Ƿztb���:Ҷ_E Z�����>�[Y�Ew%�Ma�ʴ��ü�av�x�մP]Eou�x_#�1�*�9�3Ln�0�!�� W����e%.]m�Yf�jn	�.���tw�M[�^VP���*���F�����L�i�Vd7eڧkcX�Y�ޑz���n��!QH��;$ݜ���{�qȠwR>�\�(.Ƴ#����=�2TPE�9r_����A�ۗ�����Æ�|ÏF�c8�3F'�WEجob=��ݦ�5��B�ck�T�7�5��)J}e܊mr�Y��*Z���EېH�0�NS(yD�.��4n^9ċ;�hs;��]��+��릣����_D�~�M!5s�CO*�Va��L�d�GVl\P�u�gS�汝�o;��WQL,�,e�:z��#zu�U��	_ڱ�7fS*��rB�-į*�O?�>�oe�ɽ���P�b��kS���4퀶��x�Ԃj���y����H?�H-t.L�8|��(��}y�66t�DQ_3���"&��χN�O���U�$c:�A���6*�!���X���5��wp��xt�����QT^�j�"b�#��H*�4�7���AQEMUT�<>���{�T�PQ[i�6��娪)�n����~�#�j+͛|���������>O�OC^cD��ሪ�`��MT�mIQU1�s�ERr�U��h1~sp��çN��ʃ��h�h;�5Q5QMW���b��(�����"h�������O_�]�����X�*f��}Ί&"h����N��֙���\���>����""�,[��DA^��5$SGvb���X�#�1HQ\؈��8t����xmp�mUE'��c��5U�b���*��[��uPUDDQ�qưTUS\�QT5M44�j*��k�mD_���6*
*j��-L�F��:}���t�؁Q��S"�ΰ�9�4��%rR2�����n̙��s��?����6��@��m�>;	�7I�DgX_��� ���# D�D�~BbQbU"C�����|�����o��|n�z����S�0;0�afa1OaEJe��y�ʕ�=�%���4�ȅW�!f�B�Pb��ߨ9�xM�~��z����#"�s�N/Ɣ��9��6uQ;]N���u^|tw����5k�@}� � I���q��	�y}`S���A/���C`�56�ؼL�{s�9�"_ϒJ98�	Ia>�-�Z�v�/D3�fO��&cS�+޺vT�̕��5Rh�4�����n���D�cs�052(Z�gіn�q�h/E�7026d1�!0w��]UfZ��KU!�L�l��:��1�d��i��^�tZ��b]��������y��G�D�f�-Po�#%jd��0XVz_����m�c>*���1�*����B��Q0��N�A�Ws�浟B�כ��V�%=�1����y��]��m�KH2��ai#�O�j�t{�W�A��K.���Z����/��1�S���ٙ!go_�沷�#z�s�C+�[zGtlt�h�����"���p�+�+>6��B�NL�S%��B���ֱQ��ӎ'Ow
�ys��lmm��\�5��}*EZ�>��u��{TKou��Fi[����Jʭ�id�4H�	)=�y�{1Ԝκ�#\Vo�V\�o����n͎��v���S)�sv�w��O���>\7��|���}��� D�B!�D(��x ��  ��[�R�Z�ߞ���/6WPLU@�|=�b��յ�Ӿ4��[K�6�:��B-��I��mu�b�vC�����lt�P�R����i�b�of�,�E�ʈ{lwZ����'Q�s�6�syy�ཇ
;�W����c������FoL�ZT�.~!t�m�X�Ɂ.[��848�w�]՜p�4\�{�@;�G�ܻeL��=�\��;�!��HX��g�R}`Tǵ�{�U��7��p��&,6rOC����Sm��5ŵ>�֟YR�Z���n��Y0��ieIO	�Uz�8�K�?d�vYꈙSoL��7���\zy�j=c뤟�^ZlNgWVP�h�*0ڎ����ԟ��S]U��!�W'�~S$�t�����g��D��pjP�,*"%���O:�
ego+ӧfa��5�����	�j ��,�,w!���r��6�8���C��M�-��gw�&����E5x���Y�����;���W���U��:*�v��ՠ��jמ��EM����Hy��z�����I�m	��cg��1��=!���ܨ�����l(��VK6����w���5Ҏ�*�\�I-��u�#��k�v��掵Y�]��6(&�I�绻uX�t���[��fgaS5��#�B}���23A>٪Q^�r.!i�� -�1�ϻ�	�-�I^vH��^d��bw_�d�[H��ܗ�w�����ϗ�TO�H� D��H~J�E�E�Uy��������Ѿ7���x�����<���y�<�"5��Q��������ơ����x��F�0웭�Dh{�M�j~���(m�&N0~_��p�}�@e4s�K}V���H����?S2�'��%�t���ؖ09�*��J�N��Bz�}fgl��|���PS��c���8b�X�u��f��z��SNb������e� �Y�N���T����XX��1���/�YҖ��&5���L�����
��Mz�j�lJ60}	d�=��v��o���>	pr�&ϗ7�o�!�$\��B��0;�njGW�l�����&�@,�d�`��6�s�NumKt�?��|�_i~���$k&��ۃ葫4�BN�8vM|�s�[��A�ɔђ�b�o�n�C�Sx�� �*�`-x~����~��¯�����>���'�tֹ��W8�x=��ًL���Un��YrsǕ��ɶ�7&^�ǲ��)��>��3
�iM9|7�*�5G��.q�������TI�R�u����l;���Α�B#a�&?xg�mp��\8W\Ham�[WwՖ�x�����&U0���=K)!l��2�}�}����ӭh��Z�;�f���J�G�;�,c���ʕ2�ԏ�H�2��喖�W#wܲ��"s�O�ɴ�����Z�zA�W��@,J D�($0�`� 0o{��Nb�IN�E�M��"]5��i�g��nQt���K��[��s����閴�1��o����)K��K�:6H�y�Z}������~(�e��})�n���Śy�l��ݞ�~�.�zD�����=kȌ2*�ܨ�Ӽ%����πֽ8{����ws��������ب[l�q�S�]���!|�����Oڶx�����(�|�ԇV?p��/#�����K��4�:�U��̶	u�hd{C6�?�����]Z/z�YT%wl��{��b$����\�|�[�&��E�z����D�Hx�h�F�\׬��4aY���<�7T���|��;荃 ��>4>n��;D��x����:_�L�N�8���@B��$��I�`,�f����(r��=�KF3O��t(W�Tp�Z"����ܭ�����?`�6�[\~�L��,�F� �ͻ�����<�2�dK8�}�vfB��7���zma���&C���xiߙ9��5}�Sy���@������/ڬg?�<W��7i�����XA���l�>��.��Hl����ξ4nv��h�h��n0���ϐ[��'(�
���E�y��ur�$�#r��3,<z���M� �=mֽSe\��Q{e̝i����I����fBN�/.f����o���ϟ��?>�P��D��"���?���%�_x0a���.��ev�*���"��-}���g�6��~oh�?�~*���2S�ݩ���:zq<X����c�M�5-���%�{н���z������W�-�nhcؗ)�E2��ܣ���u�eL�t�&��5�~~�)��^D���Ae��VTk���q,���g�Lq=Qՙ؆��v���PCx�l�,�f��T�����x�\��O�@Vr�ܙ�dœo�"�wF��Pk����\4�;�&�1���Vh~�S�~���SԦ)�(�L��aϯ��'+����u��8nMê��c}�^x�eB|�[�L�^�<���м0u��S�6���k�c%C��vm�h��m?����խ5��T�c	��E��ohy�)�EX�t��6-��/���J�LEt�٧F\b�Bz��2Ғ�F!r�|H��+�%�^{ʥ������`0�+����l��)��Ē�ڠ��7���j��Z��4�`�Y�k���km���UB�=�5Y6����F�[����n�c�Lc]=�\��!��v"=C�/�b�z��0�QF���M��n^̍�~"d�2�[�KE�`���|b����"n�m�OkV�M=xԤ���6�ܱb��	W��o�[炖�t�oM-X�#漽h�1#4qs���
�{��7��b&�H��������W͍�w�w������b@�R!�"U�<<7���-���͵F�v��	�E�J?-"���Pz\�yH��}kx��)���%S��M4�Z���MD�15���g�E���
թ~�>��=3�>ʽ�����]�`��%��������}�ӡ�[�s7�_O��������wW���Y�v�H��K�~��Dmg�*,d�>�����[%���ޗ\vC/j�M�g���=���`��	4���p��0�v�v�O�}�f�x��B&_�-w�k�MW7.q	���L���%4W��	����B�X�b��=�ڝ��f��}�T~��3��k��6qF��<��:�bk��;�ֱ*>��/�S��e��YM�-b[���l߫�ۭ?g��׫�+dԹU� ��]$3P��,(wL�ZT�.~+�V6�ܭ`J:�N�Լ[V�>��K���[O�ޚ�H�~C��R�?��^��1J�=��$�`,���Ѽސ�Rr�B,Sxs���8ԁ$Q�Y*rO�y�5Eab_�58?�٢�T
Gq�\F0X���0�gv�m�aҎc�X�����N�tG6����]��rg�PP�����v�ٸ�;,��޲�m�rZ��"�h>��&WA���6��ٖ�vҵvoOi���[`�|�.YǢ�L�o����n��)94�+����m�s�N��*��av�ڹ�0�΂�R�H��;F���W�k�'#۲��vQ�?�Bz_�G���ѩ{բج9$�U)��%���?��E'�~� ���P� D

�H��=���<<0��6U�A�Yt���,�A%\��F L)ʅC��'��-�+�?�C�WUԵj/���\I�z��ֽ@T�)�*��P�&����Tsr��T�����e�6����w!]=�(�/�հ���^�����P���|薽�%?b�-j|�2<L�p&ZG,ZZ���d�ʟ{;=�l[<A���}ט�/��_F='�2vF��E�ɟzzFŝ{p�v+Z��ʺ[ó���x��;����]H��ۆ�_�;X�+�[tl�����ρ�덑+iv�>�U�둡��͗�9��&��u�����?Od��C>��NO�,�&k�'Y�M6cGa�A�M�V��DC��- �p�w^3u	���[�d*�2����>�^]޿��U�tU��ς�N g��32]�D6�n�`�!����}E�}���%�,0qP��O�/Z~�yˉW���!,�#�К�mй�}U_��'�	O@c�ī�lՒ�4b�I�7��~���E�v��	�%�?��)Q��[e��@��L{�����0�kRȖM�
ڦ��o��2�8�|�a:��8��b�]�K�*ӻ���~҈5�!`���ԷsO�e ؄K�D���NR�S�U[�G���2zu����ÊY��@Tuu;�C��WMU���R,�q"T6���~}�χ��P�B��D��,B�Ĉ�����{����\J����p�,�ٍw#,\�[�e(	�^&���m�):�Ӗr^��3>.���F_s	�y�z�L	k@%7��<V�K��=:������h�dB���=8�}P+��A6����w
��ծ�`�c��ӓ�U�+kP&�%��e�F0�)���>ƾ���:��_*�ݸ�R�|T�=�fnZ��*���ԨzX��0�*�q\���ؚ�RCs$}�Yٻw�b��K�ki�\K�z�;vp���B�+��}��}l���bL�fw|���uY��YU]t�%�>z��_���Т�b�M\c��O��J~=� ϣy��Z������vW����p����~I�z	�i�lO9���讕r��ADg?O����:x�;8s�]c@2�<��y�TR��ޭ39�+��,��c$�|S�Y���+g��3�tz.����������^�ө���PƯZ�Ѧ�u���^�v'X+�#?,�����}4*ue<�_Q�]8�R�*=t�,�.�L�Ffˊm�K��بx;� �8@�"*(Q���b��b��ia�2���)��]ʩy���Õ%>��ލ�w����]Co~�M���4�(C�ME�:]wi�.iN��pbc(�P��}���4vA]i9�a��`}�Nd������bf�J�d��������D �� Ģ1((� 1 )�ߟ;����s����oW�@���Bp�3'�GL;c�����
�-@�[B~hw�RP��_3�;`���H�ڄ#]�"�T�Ľ����ͺ�Y�ͯ^E������\u����ٚ3��zK=��.�����xX����=�Qe�f����ST��~j�� �"�,�;q�wT�v��/phKC�׸t�<4��|u^���kP���p6�6�}s�F%+^6�D杺cT-� ��(����ߙ�0��:��;B���c�(���F�Mu� ��~�̡�@��ח�����v.%[b����-r�)?_���������ߵ5��v3E�2A񽃕�7�p>�}%8!鳞{q9�׷Sl�{]3`�j���aO6��U&�<��,B�����W9/m��ÓE�2�4�^;Q���{lM��t�<h��h�40�n�)��?L�� ]l��Q�F�g��	�������*�c��Ӡ��Ż�%�n硏)�ل�ze0�R��`Fx���W����]�\4r���]W�'V6/%'\
��%�+^�#�^t8M�����h��4QF\w�m��`�1�/$�~8X���\损V*ו����ƭ����1,�"����mtNw_.��s�ٶ�t٠�A�2�c�XA�i|�������N�]M|B����3^
�Y�n٦����jl���B���)CVcvx3���^`|T�Z���I|��AO�"�B#�D(� �B/��P"Q_������v��)�s�鰝-d�����ɵ���c6�zA��f	�@�k�LW:��eM*����تZ�'o��
B�T㷣S�Q��/ޟ?g�Ū���+�N��
�	>���:�����H�ݒ��u�,{�b��O�[ם�U�a�(1�V���U6�q�h.Y�q�k��c��9g}���3����M��L�q,XﶕsP~��({ϝб޼U��^@Y;�4=բ�!��}����yp�a|	�^h�>���-����,0����5�-�Ɍ������a�w5<���}�v��η=��_T)e������s �o�|�J����:��ݨV��w���0j�n���Z	�ֵ��h7�`��}0�>�e�P�֯$��8�"��b�����<��n/LU�r&�Y�쭍�y힞��콊z�/�v��_��\Ag{)�24s��}�m�B.�sp��-o7*��MNɦ��j�ېt�|�Ae@�+�cȬ���~�Ia�Y��ƭ�9��9�'m�2����ɯ&�Ц۹C'E�dsg[�!+6-�]D:�{�u[�~C��b���f�3��K�E̴��N��e���L)�4��r	t	��/��S�|W�;^�=��q��u'J����z�Z�`iv�� ���TȰN;��|a�g)��ۻvCnNԬ���o�W�̢�MF��9�WE�r����v���l�����e��6Y=�v�C��S�A��:N\���q�=m�ξ��*�� H���"7�ڛ�o����~���z�B˖�&��c}Ғ��Kch�J�\���}�\��hv�X�/�,�v��B�h��Gd�7\`Mǋ�9�|���Y:,Hu���W\�f��|3!+"�DJ���Sl_v�-8L�@�ul�\�ٓE�U��� 3�l=ϋ�'��,�;��in�0.(�\�l��zv�v��e�R�(-� ���|Y��;c��$��K�T1a[�`Ш��Ƥ���y�j�"8����R���!�U`��,�llS���Қ�F�N-������ǔ�|�*���[�yci�_qCz��v���b-�P�B��� �i�)Rb�������`�*�SDU�w�2�f�X$M�%��
�~p�Lk1�1��d�S��ܮz���,�Uz��<��z*��v� ��ҕ��P���z7:���- v�����y�\o����d�{�&�2�aeN7�B�̓�S�Vֳ�)i�`���XSUaR:<���)���ޅ���~̨h����+ޒ6��PԸ��w���3*ҋA�g�����.��Jm�={Ʋ�]>��tCN��gTP����T�g�eu����N][lC�zv�ަg�21&�̣ۙydޅ��ݘ%`��y.a9���&����֊����2��dK�-�嫱c�=m2�1��n��$�GT���Ќ݇uF�e�Iqhi0��-u	�r�'^w\�>�2q{e�N�����$�B�x8쩣���7�b�ձ�6*�M�D��.���8bSo�!�oc��DT.�;���⭩5��@0���(qfж�S���/�1Z:T˽�yb\� +J��U�?����I����v�p{ѝ��TX6��Hr]�ԁ�~��s�.�vuw��WR�G�^���q�qG�	z�9��ke���%�mk�]�Rr�yu�o�L\�\�W.����x�4 �d�Bc��ݿ�N](z��͟��I���?+"�]��&"��+iV楇�ޠT}�{:�օݗ&C�2��� S �*�����̂3	BV���WN�`4m��⹋B��ɽ�xm�8Foq.����&���syQd>v�o�����ړ8�EU���1�-5�qN�|'t���d������n��m�[
��Y��G+6��Y+!x���r���sbeP�J����P�|����P��pXV
1�8r[���,aXE�������	!a�MiR'�,�)�&"8��Ș˅�c`�rG��J
 ��УB2S	�A$M&m)���K�� �<E�"�9�ھڂ��_����*�
*���Dh�D��3�8t�zz{Q]�TDyh��.k1���Urq7�-4EW�qS� �Ç�ӧ����NBj)�c-S��q'�2<��*
v1��6����MkNO�����-��G�3AO3�j�6S�tyh))��Q%,O'�8��8��4����;�~�����79�\����`6ƍM����x���P�Umkh�Қi���(�)y8t�����(=��~�p���cQI�M��A� �*f+V�-ˑ�b���/3�\f�c�ӇOOGВ�$�4��8���4m���g�9r�U4��d�$P��ID��� ����AU��㋱�"�*$��5�J+���r䦹1ӧOOO��E���ZuMQ�����'��c�9�/9?'����Tr�D��m�k�����1���,�&���:N�l���N�6�����~ܩ��ą1QM_s�?7�������>��y���e�' +J<����;�y�&��%�l�U���ks��U��C�]wJN�f�HAc���ی ss��	���B!@�U� "D�B$� |�|��]GFpM�X����	f(Tl��1��v��*�����L�x��E� �m�T�8���W��e�=�bU0^��i�L����foc�����/��Ok��E�y�;�t��X��ٜ�e����D��9/i���c�g��G}���%}� �P�<z�1����.�o|Ǖ�v��J��]�]��򤩋R9�q?6.�淋q��>j>b��O�ѷ座#�3$�T��n��W����A�|	*-�;�M�J99Qϫ c#��TcsQ���b��u����D��Ö�:���ݣ+n�0
 ��G̵���SP�F��8
8�����rֹv��Lh3o\���٠�B�6_Wo*-�Ȑ�����Ѓ	tt��wzw�`�L�db�`w�9<�;Eʩ�jR�d�6�A��l���_��'�����|�='�F�Ɲ��r|�>�x�����A5��2o��,P�V���Q��o��
����!�`2���p�����;c��)��	��p��̡�7��pF�r��x��}�6_����/�����3�i��:45yd�qeCY5�4q��-��S�LU�㰒�m�{iU�;p0j}ڹ���8'3}��ޔ]�
�K-%,pgi�i6��J�>�B����[C�@��p�2��W}�����d�1�}��ҽ*n32J�;!v@��rx�yr"��[��e�t�٤V�ݙ_Ͼ���U��H�@4#���� B���J��!3]}�4���[6�<�A�����Siè����.���9Wɗ��\�W��!7�e��VO]�C��v�Ͽ[Ih�nx��^����0Ɛ5[Hء�.��~���;
.�w�4Z�VǭЮt��c��צ��T.m�16��gk
'|J�f簲%��Ք�.$R+��c��n�V!
b!zw��!��1V�
?���<��܃������"Y6�Z�z'b��y��vk��>��{�Zn��3-�8�b���5#.�V����GD�zqg��F�̱�\�(�8Lsĩ��t�Qsc�l)Nc���z��X_��tl����2	����ꇙ7�+U��[�2�˰ggf*X5��.�2�쨴��Y�+kP&�%�:D����a�� H�=H��mA|�Xw���q�{}U	��,�>�Qk`"XQ�uAs��j2��gu@��*���+��4-��/�	r5��k}���9N6�nW:���F,GF�RGl�W\��ON�	�Y���㡮�S/9����O
���"y�Z�-#o����4�����U�`�M�@�%ю�$K�,��a샲�.� Y�4��Gi�������>Q�.XF'���w\ñ5QU���2��u^�C�)�悸y�e�]��;����w�9�.��v��xi�4F�����4�l�p<ޣ�;���y��c�??=���ϕ���*$H	D�@R D�{�b��jh���>��|�L��;7����£���/<��z�Gpf4.��0��j�1�n���v�u(�v�L�h�A-������f��(Zvm䱿X���Cv�zO�4�����m�|[COV< P�R����ظ�*�硊03��`���͑�}�v�>)-�&'�f񁇽�\У��.��#��5�{$j��.�W��5�W���88�B(3��Z�t�������t��k��@�u�0y�	ͪ�U;c*������V>vp�O��b���|��+ �"�k�ྤ��T]�9>�"���8���6�/vI-9g�>%�ݜ*+�H�\i��}�}�@w�=�c���Cμ��"�rJz��qmW7>Louiw�Ǫ�0֩��5���֖.�Z���F��Z�R%��(VK�9'.vf��_�U�L~5��aTE�^F�`z��t��;*��2�]k�ĺǔ�VH�!��1\�<�n]���fy�A���ߦ��{�� �Sۛ���?P�k�[q8�˝2祑I���aCJ��~�Yp·cM�o�9Μ�[�4Mt4u^m^�A�K~��ׯ�e�ק��d�+��i�P D��YN^�z׫�N�K��pL�N�r�c���OЊ���vǷ'�V�vV���y��u,Fi���2��}���ƮlִN��;�)1;uc�g1�t��q�y��?��B@� D�(H,H�@�"w��������2E�o��x<
�L�z:������0���}§ț�]�5�E{(m�r�2��n���Ӫ�����p����R��%�O����0�Tv肜��L��=��p��&U�g�˳�z��6���;��6D�U|~j�c�?D��?ܠ�����8i0&a1N�6�Pܛ�Z&&![u�*M�-Jא�%G���F���o2�{#=�S���0L+~��HIGN��q�w3T�\!��sH�d���{�����SHh�Gyư�ߗ�=�Ě�kz�]8�_ss�Ru;V��F�a�P��Gs�_����P��]�oO�&7��	�vwq����}ٷ��U[+�����QL�6Kz}��X�	ԙȰ�����ci{h��]�qI�ʎ�k��5�V3�f��k�A��{�0?0�r��띷J,��`����6H1����U%�C�&������~���#��0Nj�G�hA��ߕ�|��,+?O��kcش�聉��6�&4�u�}ʬ��7��d~��_�T)w&U~��F}�OL�
��S޻k��Ɇ��6IL�ݞس�}w}�
N��� ����Ѱ��� �VeP��+��򢂳����ۺC`�׸�!B<2��/<>�ɘ�`���2ۦ���	;Ǎ\���yi�|�����p��I�2��/���]��6Q�"w5�$���T���b���8o<�y[Ʒ8y� �"D
D�D
D�R$B�@$H,�U��
Q�ͯ,�l ����b86�X���K���ޘ_�����ð"
�SQg"e���L�L]��b�σӔ�붋v	�(yA��7K�!�� ��?bg7�_yYuf���ϵ��;�x��:�5H��c#U65�5	M�Bm�Vؽ|����!��.��#lΔ��i�ݨ�)�D���ןb�a���pN��{�{0B�k�]-���2�S��Գ,Y��g=���jV�+D���j�� hת���q�W��+�k�0��B����nصU9wQ�z�y��˻F�],jH�c�Qp0^C���Py���j�	��s�?�h��EΫ4���:-h�UƬ����$^�[gޔr�d�^�>�V�b��Pe���:�ユ�	��c��B�˺d���y�؃��RNJ��;�}d�9��R�q~C���S��m�i��{1=}���ڒwb�CJ�/8��f-��'�A�;��w/���v�燍�$��h��3���
�H�F,ukz�F�^c�i[.(�x��M�����56�=R�(��Q�*9��0A��Z��T��8_2���"���Df�.��6�.N|0�4�Y�����r�'(]�y�_���]@��)V6����δ���g��[�W�C��,k���8�����ɺD���]�$��V��\�b���][��Nt�W�?�)�%% R%  B i!����~��s��:W�?���=�?���/<�K�kH���ԩ4r�-�B�z��s�u��Y���jQa����D��h�@��|�6��o�k�;��v���,�}l/&��V��ۄNƑ�]	FC队P���;Z��y��!�LSHO���펬 ����V��<�eQ��@t'�&-@�Zw�8����S����Em��vϟ�0I�,��l�W���ƌzŘ`�<Єe�(�z�����@��y����{�����g��M3(S�(��R_cZ7���3k)鐝��SQ�nǰ'��v��T�T��L;c��C�j]:�%��ڼ���ы�3�7w�d>��;�x�>u SH���SQ���t�S^>��O��mz	d�f�?3�*�;�Q�W^����0(`��[�;c�y"�2nF;�\�.�>�63���;5�q�xk������U��/�Tڕȝ�3���r���t�	>D�@M�Gj�����iֲ/��*h�:�	�:ה���
l���=YS�<���v��y��v���ly#���Ӗ��ꋊ���F)M�k0�K���J[�F߾λX�6���߸����M�G�SS�dv޼l=�bjoN�o��EP��s�:ݻM[��$�3o��z���a�1P�W�>�eD�dH(3��$5���l?�m�.Y�Ku���<=�`��Ubb"U"T"P"}� ]���j�HnǦ>�qoҩk璄��*�����xr��z ��벨����t������ehJ~Q_�OS��&C4ԫ����'yO��*����ȶq-dwgpW�Z�Wv�ʔ'Ph�������5�2�'P�jQt���A��l�n��f�\o��4����+H�� ��ܨE��VA9�Z�-;}=.½�t�4���`��;��m�9��:z���y9>��z���+�L��1,��G��9إ_/y_�_�2�W��.m	mL^=Ti���q�`�^����c�}f<������8�Y�??5}�V��~�ψ��*CU�tvoC�B�m
�()�Z]Bڅ���fc^�b�����-�;�h�vZ��a�T�a�SstB�sV�����b5룏X�1��^&y�3,,���"�|Iߞ�Փƪ{�������A�׃�g!A�A��f�sC#�74�7c>y�AT�l�b�����8w��7н^�Sy�N�м#LH���(?����z��qgT&f�s]}��h�,P���d�y�aD}��ڼ�8��3$��{k�����,�5ׁJ:rV�R�s&nP�ٸѢ;�f�]˃].B��ކ���w@P�J�ԅ���Q��;���y*me'j}��TV�X%��9��N�:�O#�\E#��JbO�?c���I���w�������t���wKQ��#��H�J� �B�?�>w�u����K7ܮ�N��?s��ƈB+����H�����nB���~�����ѧ'酧kg�3�y��t:���ƂR%���n/��R�F?���߿*o�g����H��KP�JgX^g.nDfDc3b���r�<�7`�P�6iYB�����1\�<��v������h�I즉�+��ֵ�ǝʑ�9�5��L���b��,���[�3VL06�ۖ�J}2.��4�1k�t�gN����\kO��$�)N1g���;�R~��|�[N�o�e�j������{B]RS�//�b�`|���\�5�h���[��=��)�˟�t�9���z�����'7l-�žD�6"��|}���}ʿ^.��XW���Y���DH�]y�o��R��%su����ޞ��?z"Ι��;~8��o`�ע�j��v�BLʎ�~�6��s	�q��G1)�
f�m�E��'C	`����o��}�wL�jy��o�"�##�Ǫ*ұwΤ��k��t�(��F�._^����d0��9J�}���MP!�ڭG���#�Y�-�E^��C��>�tu��D�jJY{w�>��[>��]���_��h�򴢆�EZ��Mz�(�B&f0�b'�y��4�c�Vɥ,+�q�`?c���F�Ζ�.��`g�c���ߍ^�w|��Iv�uWuC[�6A�N%[��sy����J�ĉB�)!����߽??{��k�*=������S��c1�^XȌ�oH�%XԠ��jC]j���4�h���Lzg=�}�g�6�������� p�`�G�?<0{����Xg|��W�/^wA�sGF<�G�}��|�6%۸X�����1�>VG�Ȃ³��0�l[aNZ�Z56�A˫�l�΄�>����w7,�1��z�~�꿿w��k�5��_�IQu=�=o����3EWk�h�﮺ ��-#��V0j1L���0���/Ť��2Wl2i�̸���=��.��T���[����J46ׇ�0\�Kh(z�Ǝ}bܣ�jʵZd��{Y�>]:ƦQ�q�֛�E1�*��z�M	@M�8�/^�v<��+����cyfrߘ��]-&��;� �Mf~R�0<�z	r�q�ޏ��
��OKbYjS��]�sS{R׎!��Ngە����	DBĞ��i��}�+�Tl���+��<X�lS�>"�t�+l�.�6�b]����'�cu��O-iT�pmG�f{5���i�v�p�c魟_���,:�b{�C��4<yx�?cP؟����N������_y9��ˇ�q���eiv�3�������/"��NV�gߒz�=�"X_�%����'M ��x�����n���P����+����VY+q�6�z�Β�u�]rv��D�}��2i��C:�=F����|����9���D�@� D$H)!����~o���ϾMZ��D�L-.����n�st_���_�B�B��'ވ���U]{g�̙�}k���9��B�u��\1Q���R}d��>rR���J��y���ǋ�L�߂.��w��x�˕v��FCy=���3�������̹��J��]��A�K����y��&��xZg�_!�(���M�1��Ce�ڦ�0X�x��屁�|%�d�@��ٹ���/�߱�sↃK��>�TS��,鷝(�[����hX�f_�{�h�������P��ױ��ѱ�����������T"��=������c"92ҧ6g�&:���.��/�.�[O�l���� wH�n��
:�+���Y�s�~�C�|�CO<n��W�κ�cJHR5��cl����Ѓ�7_#���Ďm�L�g��F���`y��
�Ŗw"k���e�q�;鱎�K2C�ni�v�g�x��'�/�WΣ��?�Yuyt�ܕ��^z�u�<�Q�ɞ��F�G���l�>����C4�iڊ���a�%[I�,X���2ܓO1�P�ZكU�r���=*vY����/�~�`�����Q��bt+H5�f�ȫ�E�[�4H�`�R�e�I�z�>�Ϥ�O����z���5J:���C��;z� �}�I}��������.��f�a,c�o-؟m����TeA�s���9ɻ��T����F\iۋ-����n�bz�gʦ��p��W�����[�A��<�V���
�f+=�z�Y�ج�F����Ɂ7�lPb�s�v��խ/�7ՈՎ�t_���l:Н���LҺ6�F�9kR��um����i�s+b�.̾	�fX+i/��n�{��rE�i�yO� ������Z���C��yA���We�jU�}����9�C�K�3yI&��ҹ��[�41*<>c��6^�1����bN�eE@@�C'�[9�0T5K,@�.	�
�HWE�-�EvR7�[k�݉)m+�(T�?��\�?�2+-ް��u���(8e�ݵ��Z���[Nڊ�ΘL,Y��m���	/in�o�v�].�7W���d�V	�)��Vk�r��5�d�.m���ukl�T�]�S�����]Y�f֊��(M�u&,R�ΐ���
���@��K69�#.���ʹ�:f�^'�T�E�'{hoJ�%���p��ur�_��J9�6{B��H��FͥJJ�"��2���*���J����wV�#ޠ%���a�.��H���z��6��ˎ�Y�i�ɧlY�5�1	��0ZX�W�ɫf�O"r�Q���]]��g�Gc����k/�+�f%u���� ��˶2�
���X�7�T���z�s|���ĝd�k��Wq���\�B��TN���tt�x�d��Q�9ˤ�"랷P �؉n9[��L��Ą0��+�t�h[q;�4V8�nc�SNe�ut���T�&�v6m3���9V��|D5�*�d��.暷.]����-�GIs#�.�����vY�ԙ��g������DOR��U!���*�6�!�z�����3�u��و3�g�`1t�.O�9[�Y[��J�:��Y�J��İ�k��P��BgmDVuVޜj����QL�� �:�	{�9P�ܭ�0�ky�Zi^b�\��+Ҹ�Xwj������}�;���TP;�WZ0�7�]GJt?&�F�\=��$qk K6�+��!G��{ocҽ�ĩ@��c��6V�����bqO��r�9N��ډ�����][��+/w��f�u2�jj���MQ�`<���A�t��Ϧ�u>7��܉f�&�u�&G�>�h�.]�Qd�wt;uyyϖh_�9�OT`,�9�Xp�Yg�m���	��8�Gz�uJ���N� ��9�>��B�.�(��r�gA��UoF�xe�\�r�S\���,V�h�I���J1TD^Z
��IA@k_������.ICM4QJW�DZ�xz~���{����4i����N�)�mE�����4|�D|�y& ��9,Q�OOOS����*��q���r*�����ͦ���&ъ���ւ�(�Z.Z*�m�y�1ӧOOOv1FڨѪ�t�%�15���yh9ݣ�TZ��#�|�h�
(y��çO���:v��?�o�|�|�T|�PyoF��I�m��b��?VZ���r.\�Q=:t����8\�9?y��(��j�F"j|�EA\�b�&�s��[9�UO,����zz�^ι��<���E:J4�PJV�Q~�����çN�=Oz�{��|�DˬA͎I�(�*���
)t��9�-�O5�Q��:zz�PѠ�@h�4AZ�i�c�ncU�p�RUDQW2j�&�Ѷ�DTִD�Q4j�\�9U[m6��7kj��d������>�v�ݟ��<�m1�V>���G�����NSɿwC|����%�����r�cCwF�H����0��H1(D�@Q1 ������J����ء;���оӴa��?5�E0��Z5~��^�̟��͎��C���;5�Y���K��ɋwuY�X�������S�ȵWB��-}SUm������U�w5	���������,����P�ϼa5����s&���u�g�;&瞶�f�{��k9i�s�jCj��)޻��O�tR~:�SerU���1����v�8��ۣ���E31�(ڂ{��-'RM��DU����X���N��~BnX��U�ʶ��啴�������q��Ց;}7���溶�4�|#����r����*��pR�	�>$�sw�Y�z�BG���h�uv����!�����x�@�ӟ�T_�~�ό�.�73���� ��-Q��U�@�4�j����X֑=b��thh�l}`�>5��V^=��j��!���"U�gF����gj�xK�nd�Jo%�9�?����~�$_����߄S��
~j6��i��ʺ�S:�i�
^�i0ӱ�	ϭl�虡�Pa������Ģph~?3Ǡ�U8���Kꭃ5l�*eB&����3ig'^����s[(
�DF[v�>�F�~���������4\�b����ٙGV](�v�Zr�KT����܍1p7 s�Y�O6�$O�cs����f���r॒����j��a��IhH��X�" 
{�� �nU���51�ע��=�S��hcP��L��a1�<;�k����l'9�G(3m]w����������>܉��sW&F*���lX&6�Ɏa�fl�cB����� ���������^�̰�Y����bg���� ;���]�����Q�̩b�'&��W>�����t1��Io�Z�@�/�.��|e��U��?ϳ��*-�sg:E���̾}u���Q��8��3mz����MF�b���<��U�Q�v�q����2��w�V��i�=���0���(7X0!�B�w�9M��c.��3�G��,��\��^��Vg]��u���a�Ǡ/�P��XҲ��X�\�?K�m�{k��G1�R0���v���|>�_�Y�yAq�#�%65��L���b���[Ck����r�$n!���ae�1�);M�6��@���$$!3H��d�]F�x����ؼw5`�� �e`ى�Ő�S~����)C�q|2	��3㽹���f�T$���Z�)���́z��c��7�i'N���c��{|�)[40<ƦJǨoOv-�zLo<jIջ&S�����hٻ\�ߪ]}��Q<��c�U����K�;�h��3w���k�5�O8��0�%7ݗ�.��x4�.p¬Ue�۪��0Q�(����<���4��������H�0��o�mf�+*6�aT���'�B�����	���%��3D:e�R�7s�&��MSF�r5jV�mwT�Y��]&���o�ʹ��+�mz�f��V�&�F����ǎ��J1��2��o��f�u�s��'`m��p�M��
3 �Hc=A�-�mj.� w��c�S=4�]yd�,��ܕ���Lj{���ػ�g+4�X#gS���-(��F5s+vn6��'�Q���/w=�c��~*�A#�ܬO��ɖ}b2y�;���#Q�V�H{�MS[A�p�y]��H�����"tLik�@�;
����=W5z!5�)���8��k\����E��xoT������hWX�c^��=��ő詐�����s�[*����������W��?.���ݻ�m�s�H�g��c4#TZ���w��Ϗ�G�<�ȉ���ؔ�����NU3x�;V���Z{p���U���σ[��}fx
��A��e�WF�D��)�9��]g�aPlYKl쫪����MF�E��4'��Z[���!l �A�s��p����0��T�A�� ��y�.�c�w|s��Qh�f����H�9(WR)�׻�ћ�q������ܚt)�J�M�F<�\1%峯��w��*�O���h�->��$���i����#Lf�J��X���#R�V���D� :�Õ�8	ګ�/�&$"&%�b(Oϟ?��M�7}�|ocLq�j���slMv���!6PJAm����5cH彺e^I�ix����ە�����%f��t�;i��\{��r�Y�����W�2�:���ȉ�B��gپ�L��H%�b�I��ڱ��5?R���e���]z~�}�Xp��.;k��vU�a��牃�؀F��ܺ)��M�)�0�uQ���Ի\8L���D�m�g)�ⴣ{��\c�zHo:�\��K�
�Mܔ(�����O�Th;3���xv�5e��d��= *kM�H��A�H���)Ӽ��Ԣ9�R���8xy��UMZ��b����֘��CO�C�l~h�d��۾�<ޝ�QB	����(�e���z	F1�v�lvqD�e����Z�7�-C�������C��	m��-��B�/��c(1��0�^�h<�F�v(tlS灡���P�`F�9x�P�Y��硫��}ٲ��}��u��)�4�=������K�lm���}�,D"�����oI��!Ym>�6a�T�إݍ�kn�_	�u�s��m�	�؟��o���b��;&�^�>�׋$O
��6��Y ��J����'����$�<��F�0��:���� F������#�Rw<<���of���O;R"��.Ҙ=fZ���֖3��~_�?��1!21	� >�H�"�ՠß�0d��:�\C�ad�W��y4��X������kC��Z'�~_)�%�@����-�o�@������]�z�׌���v
"���_�d�ԧ�\g�>��L��l#�&��N��W��%1ٰ�ez=�r���<�C�H�!)��b����{<.a���߽�Y�︦ϢXIF��b<̤�i1m�[�>�7wi�I�b�CwsDY�k9�4ۇ���n���ڦJj>��_eG��"w�TV��x��@��R*)�H���@^��x�h�w��3��ڮ:^6ek5?�t8�	b�"}�N���D�{�\��*4k�w㚢��3}�p��V�~���[�je��ɶ��U��A���b�׭3 }�Y��.���F~ߠ��y�0w]n�1ܲ��&����2�Z�{ؤSbQv�T\8��v\���v�0�`d^Ù�H��O����+�|Y��D;鲵�LM�y@,�z�ڇ+���)��#����ss4=���q�?0����8�-/���[��R���" ���ѻa+O�;��E{:��8֜Þ�q77�l�vּ�������K�K/(�9+��=�,��W�k�7cwIʫ-��Ohs_A|s���&��@	�R�L)�6'��1+��8޽ݜ\���PU`��nėoud��^Ͷ���w��c4.��� � �"H�bH� �~����<߾�'�|'��8����)\�])�kH�&��g)	�\�u?Nh�Nfwͷ�gqOlh�^ɨP��RGlP��w�|a�>u�:�/��.���'�ӈnz��w�	n��u��V��@g�׹\���{���G9bV2h���/=!yo�y$Bw��6�f�v�ّ5�w:�S"�Enve�>�6�C;g�D�4ّ>{g���1��kj͘d��cmBübj�V[�!.1�zO7:hWt���g�>�UU�^&1��s���
Ĝ���$��ֺCmt��*D�~��%f>���j���c�-���K���x$�s�r_�v��1;??���w�`�c�e�x�A��-�g�߫��üpE�|��[-~d7'TV�f䡽���ˍL47e�õ�Oհ� ���D;=�c�����dF��21#�W�����[�G�3���(�mz	4c4���O�^j/_?Ǽ����o�X��fRH}�Ip�)����^���h�Cе�'A�pŮ�NC�MðljbW�	�w�`��J�M��l��c�e!mI�쥷d_�K(�L�{0[��rG-L��`$-��7��:�;.s���R��ǘ�Bh���m}�5��7��a�%h�K��Ý{2�W�^B�����]�)[A�}G�1nt�]�f�V�m9��V���PD�I���?�ۿr߾Qy��c����5�1L'�Ok�:��{���h�)�C�}q��KR��u�t�b�6�L�<���1��� �q�>xR*�A/>Ɂ����q!�3��[�/�i~���l>V�~���]5U��dxw4whj�AAY{P�1��r�77=B�t�O����m�%�[�;�v2�茧@��2�_y�]Ĵ���i�|z�L���h�m��LV��wv��NVn�U��]Β�e�ؔ�g��X�}/#��](vg�Gګ���[�|�\4}b��=�D����c�y�kA��j6�X�R�˨u)��%�/�~~zYX�+M��?#��q��^�J��$�<�!�Z�[����PƮaf���k�0�,�lj.]�|�-��9.����Œ�9��ꖥ��Dj~��hȚʌ��sf�
�\m��}�\������5�m�A�{ZX2�I_�^8Q>_|�]kDP��N��IH��S�u-�Y�O���'��e#9�m�6Dr��Z�ѮE�`�g�Z��5x����;�#>ͪ>3���-{;�}z+%%�2�f.��"m����'���
29tU������K��	�i�{L��F�u��a���_�t/w�*wͩ!��,��]��;�?��Y���_cK7h���*c�!��)�e������]�w,.)��L�|�'�RҘ�yg�ʺ�<��W\�Dk3s�X������w���v4�۾	IgףU0A2%۫�'~S�E�q{�'��U���}�.�c�.�y4�����^u{����|_����=�_�(5&�.��c�NUzm��ϱj��x��J�Q~���n:�E�;zd�c�m�0ISlyM�+�w��]��5S?��6�%F���q��"^�Ű[��ۺ-cP�c)B���rMÇ�9]C";u�`jOur���Rv��[@nie���%�5ME7O���z@��A)	��VP�|(Ԣ��eSġ�� �K'�:��i󽵴��͵C�AT��kŨt)�2~��������!���V�RbX�i_��=�m�勱�ʒ7h�򟚻R�Mm>�<�t�ֶ�ͣHk�WsϕWj�⦖�^�2��S,��[R͔U�0���`P��W�i�v�ze��?��E����p5��׽��2)��"��MU>{�S��Jn䦛9d�i1P���ib�l����o6�|�ef��}�X��#΄ڸ	����׹J/L��<^��/�?yq��Ob���AJ�KO*����/��E'�ý�P�]9���$W[(#]u�[Q��3�|�hD�Bͦ��ӫ�r�KxVFm�S4-{1LA�Qե��g��ܫ������GF�7g(�S���u���hټW�h�Q�}/nCPZE�T�:�_UZ;�{>����m�Īy�T#���W����y �i{#�u���꭪�4�:_/��J�����l�02�gX�Wڇ�'�@��޿�!�~���j�A:�vJ+��d����މ�[$��0#�5��+`�}�/.�2�x�P����H�?5q<��9���ߓ�j0����y���i�.]�����;o@p][�sYy�W�i3Yk7ol�?
�P)�j�0���|��@�_l����p�Ԉ�a���c���q��7Hj�+O3k+�@�%��2:K����ӹ9���LEӐ�,3���j*-�׾�֎O�v4JJl���꾀���Z��F1��N�{t܍�� ��%�`��c����a��Xkn�����%f�%X�'_�՞����q�ݗi�i��6�Y�4eB�\w��e��z�
f�.T9�Oɉ��ӷ�N/҇��%����W�D��u�ei�Ur�5)�����3��tXSר��#}獸>T��#g��m�jЌo����j�j�o4�@�U{U��"�� >�όVNѫq�m�s�z���ݎ�z{qsm��I�s"V�����C^nj챷�q�������L����h���U�jhzM�v�ڽ����&Fanc���nG������;���,q�z�Y8��k
|seg�'�e���h.Y�t<M��n�.�)Ⱦ�,1�_�AdK&���ș���\21!���1�fɂ��Y5Įӱ�n-�ۊ^��Q�B:%c���	�=��jE���A%YϏ���G���k���Ki��xVa�k����=�~h-K4�nCR|`,>)�qoҩk�
3A:[�R+$t�8�3T��=��+;���*����O�=��E��?W�8i��a��T�P~�Q�/I�E�˳�Е�ު��B�I:�z�N�i��w�g�ݡ���P��xȷ�Kb�v�ͩԞFws�ن�kVo
����x�F.:Z�=��|H���XF�{ ���"*?�8A�m�p��"hA�vӑ8r�
d2ɥ/c*J�WO1Y�k�(-i��1����4=`eZ��鈫zz%��`������[s
��:�MґU��E�����kg�@��0����폳�f���%�%��{�i�H��4f�j�-�Ǥ�(P�BS�Ԍ�n�C�UZ佳�ފ�xS x.�;wp�c����(|/�itdL�~��##بn�F���?0�r� cl����t.nQ��j�6޺I��B�����`U���4��Q��k�C��&
��ѵ2��I�¸�i�_ŵ�˱�&\W�/�p�I�P�Ȍ�;�l�b�K7�wy�s�� Dk(Cl�s�f�<�>BQ���!yWz�v.;,WS-�Q��ѻ@u�7�ԛj���Jx�Ԝ�3��w82���󼫐��B���Ɔh�Y{XH��um�#kr�'a&���ǝ��W)+���E
��G+�u��?jy�<X(��pF�IV�;{��n�`/k�� �bj�u�;�v{�sj^���n,7�]��39e��s)�sԈ;�KF�s/%���w+q���eE�B�ƂK��ʴ}{��w���8ЫT_|�·�i�;K�T�u��}f��p���/��,��� ������7��3������� �*f�;��M˩c6��$�14�k���6G�,b���X{���Z���zrfeh�ĕf�@v�q��Լ�:�Ŗ���f�b�7�0Q��d����j��e7PD�f�6{���6kO�
�y���6�|S�k�(�G4�	w.�܋�x�e��R�^�=L�.7xm�A�o�/#�.�'6�,�mf����z�Wrf��ѧO��F'�K|
�Q�Fi����bSn�j��5=����N�a�sEP��������Af��̸�H��ғeK��᷂�n:n�A�y踏v�7��3^[��V��9��vZ嵺4�v*î�b�Kr�d3� �;Y$2�:��Σi�����;��R��]x�a��j+ܱ����;�^l��u`�'\EZB�e��ݵ6®pJ������BԨ��w��ä�u4p`}�\ ݼ�����Uy[�Kl�>�i�:
��PƔ��9�WP���bV^a�Z�b�2�+/X�҄�F%�y�ˡЊ��vfZR"���i�y�踧>M��i��!��%6�T�v.؄[�A\��S���m�m��ŷ&��孌γ�A!٘׺�	�̙ܬ�ƕ[",���X٣K��Ut�ٺ)���/c�s	v)��W��hBg�jd&"�s���Ud����1�*�tS�<����Y�y�H�G�:ZA�q�1�N6r�f��o�K�`ᮇ4�y/����*}T2�%�"���e[j��8\����}��̰g��aЧserV�S��P�N��ę)�82:��gv+sE���ȋJ���#�dWEi�|rP��"\�dml��xu���麉v(2[�0#������r�[k/���Э"2�9t�#l�-$(cw�T�)�G˜x��s+u^e�'zڨ����N+s�{4h���p���IR�t�\�W�t^���Cd>��Xp��bZ��-A�A���*��8e�o��L�y1.��u@�o�v���F�Js�6���-ڷK)����܋�����(����ne٢Ї~�BѸ���Uп�M��'�e�:�
�d����� ��.S��B�XThq���Yv]@��ʂ}�ga AE@$��?��ɩ�8�S��W�w5���[b�ڊ��������ߘ��.[��*ӝ�����h��?�U����!�U��E1�c���TW1��������$EU��T퍋bh�ꈂ"���*����TUV-**"��������cAS4Q�$��5LE�TU�7��G���Z� ���UQӧN����LQi�(�v�11,DDX�V�rh�*���">�O����$CELSF������"���'1��լbJ���������{j��(��4ykC���N�v��ڢ��AAI��G�sӧN�OA���SIUI��!�PV5��B��bmOc���ʯ�8�8~��������6� $����
����Z�DJP[4��ꨊ����?6)��#Z�M,DU��%�`�"�����`\�}E��t`�Y��B�r�p6�A�))�i��I������i�l��Ɣ縴��v�R��[˺�jJa��
#�߀]��p�����XkD��0u5��W����ɳ�_�Ac�o{8��u'�낒ʭ;M��s��zc���[D�s˾�q��`D(�;��m���x�4^-$����͆�9�����&q��s�>��y����4���u]mQ0��`>9OG%��]���]����S.�>S�lh|��'!��dKz�˦�ߔ_�s��؎���`��Y���'!�͵_�5����3�W�\�3�ت�����d�XW"mu�-�ShҶ��;s����.�3�ih�Mɞ�%�s�_�Z����R9�tBkjЙ'Z�md��Ller[����L��8�C	��e��m����F��0����W�߰,ΡC�����k�����H���Žq�2�ՒhT��ٗB�}u�Xk12 ���X��~>�C`� 3[��u�AY��ϖ7��s�rk0��$�x�OIE2�XS퐬卹����!t�V\^${]E����Z=�%��H��Ls*d
�;�l��0���(�Z�GK���)s�鈇�P��co~������7��~:�M�V�q���Y�i�wZ���V�]��xl���i�
�e���K{>Ц�(i�3X�e���O	�w݄�2׷WҝsM�7�,tH������b��ް<�3��lױ���ֲ�!�t��̎�-�#p��'��kQ���o��n�`kYz�?�<�R'�ɗ	�\��FKRN��a@'��-��؟�3��<��S����j�k2�d�w.�s�T{bѡT;�psb�Tw8���R�6G�Cm�3�Z���8���c���^��Nd�W�ڠk|�C��q�7"�g%&2)f7\��i�+��\��(5-�gs��T>D�Z�-~!��΋t�!F�<(a]�i�[��G'��ck���O(9F�׉�gנj�H&Ļu`��Oσ\���4Q>P�dn���n��ދy��������O����9CTG��<w@�iF�ũ�Դ:�Ϯ]��y�D�N����I��G%b���Y�� ���OC��ۻf?"5Ƀ6�f(5� ��=���=���u�m�eed�Y��y�n�/5�a>�Q�sq���ę�eh�!2a->�TCY����ý�,ք殍�r�Ƞ�*<�Tõ�xl�u!���.9�}w6�ILK��i�����u�.�"Ⲣ�������*V����ۆ	�q�9RVI�f�},��5�;��i�*�fG�N��T�0*f���M��=Հ�s�3�ζQ��8:���۰�o�O,5�,�z���pC�cz�~�,�4Ք��i�2c�9C2K�Z���?6���J���aA�fVjc)i��G�+2��2��h�a�X�5�EJ {:��������1-��Ek{h"�pf{n_�;�.�v�����\<ǋ�E��[g���y�n�Y*i0�r��"�����)������i� W����5���޻%z`��1��s����h��^�������<L8��^��v�7Q�c ���\c�����S�)����2��ڸ�3���)E�_����֔sm ��~d�k�u�&rjV�v��.B�p/��<������0����Tu���w�P���U�ӿ6��x=���Az�{�"�w�x~4>G�4�
A���}��|Dm��X2�=�1P��OrYL�����L���P%�ЂPY��G�5H��6&4�/l˾Y��S��߅.>�'D��7�19k
kwL�� �Zb�j��R	�i$\�O![� kC�A�Q{U�j!��#�*�Fc���u�E�$���$O'��3�i�!�'���p�ƿu�΢Ib�����-��[�w���8B^7`T��.��nu�z�ls􋼹�V�	^�Z���t<eX�뒼��M����
�Jq*w��T���v�U�D���h�c�5�X�rR�����{�U�ɑix���W�qz�3��:hr,�7[�l�I���W5��.����s�H7��"�V��e�����J���w}^��1¼5�/�L\F��r�;kF�9�w����zڙ��e�|����h`���v�9>m��g ����$��4;�!�c�һ�����U���x�TKL���*������;���?K\��s�,x��u��4���Uڻ�����)pmA)v�QƠ�j].Ċ�194m�/������n���To�ҘL�u]��}ky�֘D�N�Qv׵�ś^�Q-t5e;	�=�0NJ����ނ��o�+��6v�p�ܝX���Ӯ�u��m@�Ξ��t:iW.����n���P�U����.������`��[4�*�=Q7�1���R(5i�n�H\��ǿwBeε�>�R6/(�z�8���
�|,��}N�oc��F�ߋ������~���y��qoҩk�B���*���4����_/j��=����rpF�G�?xC���1�>[)�/��	wON'�)�j�r��;U�I��&��c�R�{ò�X���n�4���#|<Нs���$��xd�D˷P�⯮rQ��j嗔kMNE^��T��3��tke$v�~�c��ie��`�!�(�|�i��a�߽5a�!�zI��|�󫤾y)߮͸E��ID�hU�ݱ�㥓sE�R�i��j��tN�f��D�����a�G؛��DU����Jr�r��g5���nL6T�ŧY�/��7�
�ɟ�^ݖ�x�Z���\��Z�<wa��G��^��x.����"�>���CN?�3;���x��8")�*��m����e̗P�Q�]`cб��>P�8�iP-y�������?�����߾���J� Kͺ׿S�O�0&��v9�9���&c���[?���>�IPZ�@��zٷ���[.��
p�ݵ���8P����Jq�����\�UL�ӇU�jmZ��'�c����Ͽ(9
�1Y��][��y�kO�G�`��w����Z�r�݌�*:y��Ȱ���p��E����D�:����,<wʄ���Gkn�S�q�d�K�)L��mm�4f�bM�q/{�`?z?�|ݗ�\�[�Ɩ"VT��(�g`�S�66f֎�p���i:F� �>k
�b@�n�w~MQ�3�$K?[D�A�Uά��s�]�]����t.�fð�V�#	QY��������PC�{��fev#�J��v/mĶ�m���2�[6�T���φs�ؤ�=Ƨ��Y�N�sn*p�������Tb�����^eG�@�u�V����|�_{��1�cVTM�z����#WV�������c����)'�ZQ����hϻ|Y&��r��wViRFAt���s�eM�C�y�C��ܥ�-��*.��TGp�y�D��[��X՝Ga��.oR��:�j�b����7�EW��6���70��[ԓ���"n�d�^��ij=�ss(����5��|����q�����1{+�2� �0��&�|����A�ĭ"��^Iڸ��5!����c��d����י��1yk���e�|]+�7AT9I��%t�{�^��~y�S��wg/Ԟ\K;�3������D�������oL�<������'\����#�<��Y�G����l��=��r�+�h�D��Z��X%,��t�m��srn�ݏV.�3����1�*ײ���3rє(�5y�x�ڽ��j)�q�=ss����(�4��=GӢ�ϴa��jic�1��/}��Ed჏��<Ѿ �p�}�F�G���g�4��Kj�2�nRs&��u�8m��ۛ����A�⊺'Z�̞��z[L��d[l��XkZƴ�I��ݖ�g)hJ\�W��9����<�D��B�����`�������5[M׌���1���72Y8�f�}C�=�?{^�Y��Mʀ��a��WrYu����x
�R^X��+�m�*�D�Q�&�~�vp����zK��c���Z�+��8�z9�{d_q�<붻Q��B�s2��r^����N�'�82���n�8�r�l���B�M�����So5��b=ʓr�];2ѽCl=���M�s�>�C`i>k�")&�ׅ�`��d���/�SDl�կЮ�;��+NGy~�<Gu%+�3im��L7�,Ou������A>�����gLi��sz6%l8^J�r��Y�x��WK���P+���)��4���|�0�bB�W�v���x�L֎��s���%yT1[�P[���n�8�������4�h����'v��ju�� ;�-��u,���EZ�V>�2����ڙ%�S�Y������v���Y�#I�9��Ld����q���gxQ��3d��>J��`s��r=:�^�GrDr����V���qFM�������8`�����<�L%�LPجgԺ�9C�%rکg��YǷ���;����A*��lm#�j�C�w��`����cהg�ʜ��u�7~��q`�G��ڜL&�qfV]���s���1��*5xdM:��KâYԲSlY�+VP�r��R�Q�ko���E�r�a�X��6��"����໶rL����h��`Gx���n�N�#�(
����.�P��{��D�ri�&�a�(+�+�p�S�MѬC�[�}J���<�n-�-n����e�'�ou���.A;$Sw�[�y�dN1[�*�w��Y5{���qtc��G�H��V3<L�kΙ�@�d���E2�m���;�su�(_5J�Ĥ@Xd]�-���0Yn�X��ܶ�W�����5gа}�f�!�������A�]�Ἥ~;F_s{��=�Δ�豃�U�~�gP��0o�z��,,;���h��
W�	f�ʆގ�s��{�7X�6:Ie�
�h�:~�<d5�B3�(E]!��l�5&*mc#J-ݸ����'��6��7Z��}��#��l���/v{k.�].q�3,��G����)Q�bk��$V��al�rk�\���56��KH����7�^��(���������U}�mx�e`�~��u��ʆ_V~&%��:<�a�ɤ����yi
��`��Uf�!����a�(����؎J��W.��5�tF
�ͅ|��XRj��t��)m�նo!95��.��X������聜9�ر©�W%哝��%�^i�Zqʨ�����oFю?і�( �.�dK��o�<&������|��Q���X��oU�M~�
���t@2�)#���{ ��>��o�x�V�\�֕#q�vd�)���޾&�@ķ����d�od]���v҈$�y�ޤ��ߺ��y�Epg�K&<F���x��z�\*΋��<p���G:�m�rBG8Ty�Z��D��]3�e��>\=��$pZ�����n��J}�uu���cVO�!��<������)�*�K�mt�U�a�g�V�tAZ��	Y�@�_���WΆMJe�Gr'dhl����;q�xu
�f�>��J��WV��ţ���<�[���;�S���e��9�0S�)�#�v���==_��Q�J/�]�����Cwg���'����y�Z-cm�TD<���6�e@Lqw5+���K��S��B`��S�2^��a:DX2޸�$ ��C0x� ���ˢ�1�]�c9q-��\��L�]���)Q��*��f��c��^���ߎ�(@�~�i�(�8���0��ϰ���*��te��F��J\�Y�Ʈ���	����ϨVR�z�m�H�6ﾪ�P�7ʯ�Ŏ?�~�5�-�����*�j�Z�V���Xy<���/M��V��@�Que��1S�b/(����mu<��V���F E�ܽ��_tS�[n���t�"�DtǦv P��:�W �{��іϲ�ދ��yך8k:Z��b"q�:����g�f�-[��t���Et�˚:��YOO��Os��U��<l��2�1�k�@5p�CY`D�XZYS��6-L���z':�n�&*�q8(���,�d����W+�lh]��0��Y�7���bl��]�o��w(3=T����Kf�iO�	h�+v�+dgm9���T8��Y�	�2u���Im~��U<�	V��-��%P���Y�v	�3RY{�]$�U�����Z�宬�L����y�َ:;�v%Uفۇ��j+w�;��g(�u̞�:�T��3��YmO���.��ў�c���x�� /"E���1��c�OC�t���}�'"����&q�+2d08�oe�:������y[��@��}��bɶ�F��{9=x)�ELѷ��4��o0��%O��]��51	�5Mq2�i�8�t��T��hr�u���x[��DoS+��;\D�<�7�]������7�'Y9_bD��ir$�>[yw���(�vb�� �|�-�~:�H��n���,M��ʵx�tZP��qoS���(n�Jٰ�yKw�R���vĲf֩�����E��)w�;1&{�4`��1n�Z�k��8Ca^���`Ҕ���-�Ձ�th�2��0�
�ᔅ (M�1
�N�u �9j�E�]�eu�x�5's�<uA31S��X-��qd)�;��C�T�ӎ��q��K�j�n�٢P �T5n�9�21����K���G�����������\d��ٲr�9*�g���V��p־rB��5"�t�r���%��i+<�ڏv�T��� ��u����U��ٙ���eՃts�R'�uj�K�}����j���]1��<��I�;��Qe�nm�[�{5�b��'T���:u�=�1�D�xU���г���f�u"<M���ϒV�Ō�C2����4��c�sի���w��dR:�C)��]��<�f��XГc���(��i	�)����5�9[]�2Uh���*��6�*,����>����ݾ�f��.�6H\Er�7�Eb��1�Q�/D���Ԧ�ڀ��9P��*� �Z����{7����b����D�Q;�]>�T�����[��m��Q���.�t�=�z!�+�M.�vf>��sy��}q�v(�]$.�^|N�h��y.��I�>�	Ǯ����/b&X����fm9�P��olkW��$#h��x��s� �6�#ŧ��.�ż9<�s�]�i��f�P❎��m��uRԨs�����AM\+$�>�5u�gh:cG���I��'�6�m]���7L���[/��Q��:��!.\$�}�xJ�h���Z��;2�ܹ0՞d8i�z��D�')�:�UŢ	m\�����9M9ub�{�z�W�d#{�K��w�"�D�����a��ꗂ]�)-��śڙn�ZB�k�T H�B�8ۣ��6w���i�v�.���^<�cV18�nO��U$}W����eqn�W;Œ���(Rњ�K˷�򧰾������36<xl��;�q�����Ɋj;�`Ѣ.�]C,q]0�	p�5��v�;��%4��F��v���CoZ+��b��6m�3j�5�Wu|e�0�6g�̹y�_8:��"��[�c��¿&ȇp��ʹ��|�����#ՙC��ٮ5����8��1\2���{�:h"#aۚ�:V.̈�9���}�[Rq��sI�[���#2��b|Λ�(���e�\HǹINиlۭ�=��;��z�mIM�!g^#�-�d�UE-34:j�mi�R�ѣ$AW3�[Ə���~���j��9��у�"	":�����tN�Q4Dl�#gF��O�N����A�V�-Ug:
�EDD�A��6Ѿ�2�Tֱ6��#���}==Ҋ���ncU�
�m�bvU�i�4:�Ѡщ�-5�����}>�OO_Hh����Ce��BEliM'�˒Q��y�I��IF���>O����G��.Ks;f�����F����K���G$�\��R\Ƹ%�1���~=Rb�a]7��94m���m�TRX�Dt�ӧ����U}�P�����	F�&��J4�F��"kT;j�<��y�>O���4Pzlh�F��F�Ӊ��iq�� �Eb�Ū�X�n�U\�:ub��FlE7�r�Ju�b!�5�i:N����@�mE'зcE���{�8#��V�u5�6.��r:�{����Jt;��m�/dc;n݊�k�2���n�0'�f�FZR��_}�}.��x3�����
;>�`Gx��oH��>���T��y��;rR�^WUp�g�#I{��1ݑ��x�y�[�CbSo��k�Y�#m�fW^J0�(�;�V	ت�ٛ�`��6E��lqi�7�:�ʨ�(�]��&��t��Tؾ��܍Ϳ5�G���� �j�!��n��{�.��V��;�� ��������zT����Z���K\1U�<:�<]�3�x�[����6�ו��S�n�����աљ��/I��&��_!�;�M��9S�mi�l�u~�l3���`=r��J�P��^�$���e:�3���䒻�@ɺ���C��K�k��Ϟ��01烁��n,�oq��X�����d���`��mP�ZT7l*�=hQ�G/LU�S��ˮ-�N815ٴ��.J�&�Z��^E>[��"�s�:e�������OF�%5-PN����-��i���b!�92vmi�3�c[jW����ˣC]��,���fR����ҷ�.��2���q��Z��:��
-p���'w]�7��pX�ڳ#�t�aEE\g;=qkZ1����E����פ#�m\�}�(��Gm����j��d��	���\is�󸍭؉�:�]W��B-��#���4wYF�0�>/Fѡrz3��սW�l�oּOf���gK�0d�P�p�]I��?f��
�����>��Gzܢ��'k��1W�u��gCpZ�!��D-��&&[�d����s��L��Fx��:���{Sf��5�tv�o[>��Fkt刮��L&g�J�����g�'���f���9��*����կ�y��W�GY�r��[��8���������J��p1�]|���D�a��0���CV3r�,$�͋�j����ls�bz���)������ng���`2���>y��g���H�\�`��w�j��S��h��xZ �w/I�~�ιkx	�e��*�iS猏5�CBL��z��z��j=.�/ߙ5��[Y�.ar(�5�+�V�cIGy�ޣ���2�R��V�孀	h�c%`#;;��r.�d�]�e�_]ݾ�cª��k^u�Ɏ�y�熴6n����~7W����IH�4��\�S�6ONP�:|��v����JF��r����6(��z�^�)��e��쏄��Ew3b��%4?}���x�4�ΰ�A87ls��Ҳ|U�B4�xb���y��qp9(��xJ��c__^n[�vT�Q��5�E��T�V�G+w���/A:{
{n6�1۪5nhǙ�sC�Ղ!�]	��n+�٣9id��VN$�te�s=4���yl眢w!�5p�'ͱ2<�@��9+/R���Bʬ�O�f����1w+a�0�Vݳ�N4�˔�h���|���7AU�a��$�����S5�q3�]�&��H�pĞ���S����8��7�$cd�Ҙʕ�zg*�9���ݰ�*���u(��|+ΖȂ4����N�����َ�oG����I�`�\����G�;Z����~�S��ǦF�|�z�a���"$��خS"�;��R�W�6��=�����gR�j��S*�v��ӏF�!�TƒE	��IqZ�w�g��in��:f�Ş3M��?����)�ӽ��T�)]@��VL����l�Z>�^x0��3rT��!ףt)�s���Тr����t1{��{g'l��#t��d�/�)	��rN������������\�"����;H���}X�$����h
��<�`�������wJ�'R>���7��=<�'��I�vVgz��(w�C�����b�
�}]!�K�gY���s6��R֋�ӧ��v��4A�ۀ�Z[Heo7��d�M�`b���*`���|j�9>Y���[�FL�����W��E��v��<��g��rm<Na���W�C�u�62}��$��t>�"�m���e��z�6���V���q����{->��"F�(���lc�2�����DC۴��j�{U>������X��i�]��7g2z���l�G��w�����i��8:bUו-��X;ODlG���������y4-˪�:�x��k��������M�RS�7�w���M��'{�E"l-��+�0��X��13=�9�g��ƻT7]q�R�����tqoV -�X4ggt�L�ה�=���)��P�|��R�yJX��ۧx�T[�pJP�tX$���pɝZ�t饺�	�$�u�w��t��F��T)�%�O>�´9��xG4P�o�;4�|��;�ޟ���3H�)�5o�n�%X�'��A����PXU���C2�/:�S	������yf�7$*�.;A�_y*i~O+V�֔��qyڽ��b6�Wgٻ�e߁c3I����]�V�y�>��IB�h��e{�q�������LAw3���w]D�hpق<ݑ�!��.��F{���S:�����ھ#��txjfk�#���H�!M�\6k`��hN���=̯Q�b_n7h��o	
$����א�� g+�u!�1����KZ[��'�Q(������3a�t�ƶ���D� Ql�d��-C~;����\x�u^qOSY1���� 6Z�B�<-d}�֮l����\�f���J�,O�Ưa���e�G�u�S��X���l$n�Á4K[�~�\�*�.��,��Ӗ�:Y�!�\6�g�]��E�U�7Bˋ�h�gOdF��W�,�7�9��GL�<�~	��+��GVumh'�*�#}:���E��P�Nm���t��M���=��t�P;�x�پ*E�Đ��n�����s��enT�|O�Ng� 7<VK�6�UsX��h��b�4J)��3@ާ[2�<Ts�kK7t���f��#l�b�t��i{0p���R�)X鶏Z�}��ow��Ј�\��n�Y�cv����LG�t��܂uq�Ob�F�b�x`6����GZ�h��X����{[���q?s^���7<o�,���R�&��,*��:x�Fk�e��n��銜j��3��:Gk���-�!�� �u�K�Ҭ-x�Q�y%��<���#���5q��[���*���sH�n\\gnӷ;�;��Yǟ#f*R�)l��uzs�V���:��b�<����p��q.fļC,]k�jn=7���O/�h?!�IVh�%����jv�qyh�Ǎ��ԏa�x��9w�6hGU�3�uk[�m7ɳt>����
�B��Gw�*�j���*�2��;E�[l^:�V����:�6Se��_�c1�G�>��E~�u���IYxIU ��y�������/�p21�]"ku��9�����}9f���$^V2��n�\H��U8f;	E�5�vme=��>�!GpȢ�yrr�`�[�Щ��I+��e���t��6FvZ�M����_,�����UA���1��v`���ɹ/��w����(�X�5U6��-2vV]EՖ1ñ��7_���������i�t���#:���޻휺��Ds��F�e{��ڋ���by^Ѷ6Fa�ɭ���fr܌5���7x��ݠ�`���yu��ؽ��k�"D�U/3���]T�V�X�'4�wE%��0$��̳E+f�i���e¼�$r�ܑ���n���'��p=@,�������$1'��l�r�x�K!��{���gR���:^��6RQ�S�-�v�'�YW�K%mx�����s�Bڐ�a�/;�3N�F�˹�ݳOo��rR/Xs��	m��wM���R7=��I�u����j�j���`�Q!��������"�K��Q�ŕs�>��m�7�߻v�=��f�A�[C��H;�,��$F�l��Q�g��%c6��jkq������5�6�]���q�.e�.���Ӄ۟.}wvtތYW�;��H�L���؄��;&��ͭ���P07wl�\P�s��_A})B���i��B7eq]���{�ŕ�R|{�e��kd	n{�2lc�L6�8C�n�:Ir.�X+<z�j:M3���=;7"6�*���2�*˷	�^���bhs�o;+�s�z���:�/���\l��Ǒ�)��^'8@��T֮w+v�7<S���ot��h����r�R{��N��>t�;s��T�%kڬ�W�4�~���&{�v�����U��YC�5���m��C��iW�w{V��N�a��Ì�� �6Gp�}&�J���U���ݐn7r�)��\�$[������O{L��8U��!�Ѯ�L��fDn���b!��[\��Zf̆5����<���yYnCv⪛��`�ޱ�ʽ��yZ��:��2	����U(��h����h�f�]���E�x��`l��٥�<8��@� R�#U:��ȫ��֍�fo;�oǻߒy (n~�Wz~r��]��3>�5���FQ�LMhOUA�vTK�n�-ծYE4r�z�aW������)�{fsϓO������*?�Mw�	*�־��R�$���!�t`�8�d��;;�͟9��}n�	c����V�[�������S�Ѻ9�J�a��E�K�zn쫮�x��F�;6x����D5�^ϝ`�2*,��T�\�	{hgB�������I�������=�K�������ܺ^:��Pk��N	�-�A˘�5r��)��WU��K�ӎ��{�rk��z��ߡ4}D"}�7��9٭Y]�'k\��QF���b�����j����=�w��*�кsm�c��	���dD��Ѩ��(����[
��A7�s_]�v�[Lvuo.�|���T!�"��h��l���h�y;Kw!�h|�wSsL�����T�jOy��
�K���z�y��ѽ�%b��ȇ�O��-4a��b�����V�C3�`�T��c6��bM�0ӂ���^Ϊjɮ���'1e����Sl��|o�ˌ�u���Y}˷-�o3g�L7>�s�x��E�i8�p;�d�,W︃�G������g��ɶ����|D�sL|a�]���uـm�t
����j����R^w���Fu�W�������;b��gj��(%��9���̅}��Gς�f��)�s�e�7u�-�{Δ�l��QY��5І��U�+���j��*#p��1���'nx�d��=@�����	�[bň���q��"��mH81�f����Zx�	�!�5��-dsD�:r��odt<y�<�W/i�A�X`E6/��m���9��W��Gp�볺��ϕ3���m��β��]��5�~�K��W���~\籔���K3��( O�-X��L��f���� N�EH�I6ۦ.�7	٫�؋S���=Sd��8��R��w�N�6Z����[�x�OMZ[�Vb�'ne��N��в�܄,Yl��U�Ѽ-�lj�nP"+�ml���k^����
p.��}�>��KdT����z�s�%xC�FbM���38n1�#���3���V{�����?W���:Җ>eI�2��̫�>&́�DFP+&Cc�ր��
�z���w$gޠ=�z�kd35�v�X�'��5�t�˯dOQ$.�,��N��IӬk3U��.�����ΉAuEM��s6Ԯ�Kh��Ae	�9/hBv��v ��h��(�󬕔tcI�%��ҷ�O}����i�3:~��]^MrU���D�7�̲�{u�h)��L�����)9��W���n8�;��cM_e�r�t�E�ӻ��vv�ֻu��|��SH�FG)���{�i���]M=f��B2��@.g��[��,������o
y�]����>�,�!���yu�+2]�3J�[��-�)-O���&�{���5�q�7�+f���K��ً`�7�4��сM���z��NK{�>;븶� �P�9SM�p[�R�C(�U�vÐ�P�h�H��L3�ދ27�tw�����Awvm�Be�6d��w��XT�ׁ�2�:³)Y$��H���OX�Vdtq&)N4���s��k}FR�ٚqwo3�i�}�~��l�"C�^�5g��tB��ӵ�/�i��ג(�gGA�J�e�e��D���<�����O�W�>��fRܡ[�����IF�"���(��1K�Y� ��gl{a�tBN��S�v�j�$����M��u��8Ƣ�G�'?Gx�P��0�2�\9�7�9�4�;Y);7k�gw����@����a+S ��Y�u5�;�Yõ��P`��ԸVuhI๚G^��أUu�2��atu��qZ
���AA��N�]��L�Z��w��7R� NeQ=�	�}���HQTck��&\M>�dʸ��+����y�^bޠ[��zTkp �KH����`��1S���.�Jbr�Hi��>���J�ڷ��v���.�&]��F�E�m�"��R���g,�͢��f�7s�2��cr�����:�7Pb[\7���������l�C�TY���Ċ��Z�gnXR7N��.j»�)k�Y*u:��fXo�L6T��(���'s���+��"�����f
�P��w���h�c�D�l��+��s3T+Dj\�Pu9�tL�j���u���i�:!�d��Ӆ]s���,
�j��?�u�
,�5{v�$6>9-���Q���.څ�Zs [-��I;}N��}���  X��[�#������'&�{ri�ofɡ�6�U��H�^�ʝC.�X�,�UN�w�ۚ~��U��+-_HU����`L��A�3��]�ͼ{!-�ﻏ0�<�{<����M��։��Gecu3s�E�)c����]0�SDO��ODɴ$�a��̆7w�LMYv"�o1@�ͼxW� C�*vԚ�f:�-9��Sį^��nL��L���L@G.i��guJ�׼�B�9��윅"��w}�B�KK��M�?[�K�:��LF,��7��o2�x����h��`�Q8�IBӄ��e�	K�p&���-G#h���Q�(�?CM�!AFB�"$)�"�4�$_+��������^�c�^��6;�G �j��K��i�A���8\ԓ62V64c�������6��lh4��6յ� "��T_9�g�U�P�Z6�44����������Z��5@bqhш"
����-mo�8<�6�ZΜKL�A��:J1��}>�����`��0U5N�g��h�j��3g�(�m�Uh֛cm���C�}<>�O��^�Ѫ���hJ.����NG$�b�j�M!CC�6�N��V:t�������<""������R֫C��rѢ�&�΂�I��0�ѧ?���~�����P�&$�ꔡ��֨�-�h�Q�m5VڣT�������}>�����K��j�&�N���[cAT�[:)���&���c�������b���DUiш�X�٬S�ce����i��Zb4�`�G$"�����D[d���أI����;d��EP�b٣�oߝ�?|��A���+c'1ֆ�і���e����Q��c�+C1Φea�)Ⱥ&s����5c�F�-��]p9Y\D���1"cP��_�/��kꩡ�<��og?��X���IgT"��-"��g��~bS�#�{5�*<v��� �e#}��*^��s���ê��\s�ݦXd}�/�%����l�j����L��en���$��i���^�������a�_�Q�����Z{��~ii�9��+�׎��0� ��)�eEd�M�r1�vcfC�����F�fEʇÓ��˫ޅ�zJx~���~���J'��/��#�sܤ����o�wH�E��˳�q��n��.��{X�
|P:����Et��׬1���!���}ｃ�x��&�����s����r#���'H-c<�K��������x���L2�q���ӭ�&��/Kv��3;7�s#���6���^����Ԏ��=���=_I���òn��(ӏ3�pb�٭�^B�F�"*u[_*w,��=b�lm�8��:F�fŘ�,K�.�m��M�+����q�2ݔ��YS�h<1e�츖�z-1{���vB]�x�.�Z6Z��_(����z�fpكvᩎ��4��oM�5�V�3B���J�*f(_v',��k�Ἥ�׷)����g{xӽ���ۀǦCҫ�:�H�W jY\�%���\�R�<f}��=�|�I)f�7+3��ɷ�^&�T�H���N�R���|����5��YIfET�"�B�t�q�� �p�W�`��9��m�;k!����,箁'M5f�n���H;�-n0��!k��ɶT:���i���;{�$�'���Y���~�;?8E��<���[�I�O��.k"�P�7
����S��$"�=$S��F����;�F��ќ�����B�Ґ��T�2.6%3���II]<}�	��r��i��LK���G�E�~�gh�.ٜ5��Z�!��b����w�6J�i�`�W(���m������M�����p�
t���~[Y)�ԬӯU�k�< ˮ�lل"�6�J���|��6�=�0�]��`NW//�]��W+�p�^��Vt��ᵒ�L,�'��Gz2���1�!��T+{l%κ�l�6p�:3��	TY�獊-�Ff%w]��Z�:�Y���-����'xY����⺱M���]�7�m�&�'vJ:�f�LS���9gi熅�x����&��-<��۰k&{��6e�����w�w��<�;��`����.��.��#Z�t��ӛ\�Y͇�P�Юv�xP��Mm���I��1/���#昛�0��l�<GW�؀
��6�1���6�6�+.�C��6u��֚ʱ]v��ܝ��?A��z�K��9;��ؿn�dRDu���!v�X�<{�����`�)�����c��~�����)��}`��ƫ0�"*�9E�K')u�~Վ��
�������.�'�WvtJ�3~���8³�械��U��J��mԋ�]>k���c,��]������p��B�l����	e�)eu��򜉦��\��t�4��9fŋ {�f��
���5H<9ͅ�iwX��U�х���]�h�89�3ja��j��E���7{�P/�E�`'��TӳLth�m�ǭ�u����ٚ;b;��[�}�˶z��ȳoîv��/2�#3����㜾o�0n�H�� �:�u����L��YZlbM�{}�(�������<��Ɏ����e�ӛ�Y�ӊ8��=����>Q�!��	�#_��.e[׿^e�M�q�P���藾��N���MM7sw|�{=X��Ix߂����цgl� 2�w�a����h��A�}��SV��D���l����Xs\ר��B�I�n���Š\X�@�5�8�F�m�p�����%ey.{�(����Pt�0�jϵ�t�6�t���^s6R�@�2.Ly��dg#��el�3 ��뫅Q��Q�xs��th�����\33�T��ȁ�d\������m�6/j������|J�O��(�~���G�2i��.���`呠J�"3����ܰi&6��S�tFli�qh�'��{w�5e�;��]�	)&�[�\2�Q77��3����"��'�h%��Z3��k��C�@�0}w��Ux�x�a�E�M�G>^�F�	p�fd��x����h�\=D��e�1C�IT��%�ߒ�ͽ髢���,.�N���;%�{���3��h"lZwP�����N��Aq��Oqy�u��ʪ	�I�xs�r������}�j}�p.L
�����f]ʘY��A���f�vJ�����j����s���R��-�����+O�%"��JC <�yyy��~��ŭ�������Hpr����*ɵN���.NԀ�n͝�ّ8Z�<ʮ_ZV)a���C�R�J��ɼ��MqٹsW�ْGC�%�W�+'tD�{Z9���3�pDj[��y\U*V�<�}���m����W��RV����r_ ����Z��h��.l$�Z���f��Ă^./w������ԕ��/ �t���`�8k���7�L��e�i�~n�N�v��ʀO�h�%gW���#������-��l�y|��4��m�
jN�uzaEtG�����0��匱[M�'������y��ny��h�j1����fv� ��X��_x�>�1�z�*�B�$&T��ܥήڋ��"��
�d2-�3g����P���7��G��*��݇ʻ��eO52�gXe#��X=�"�3#����a�`Z�v��T����f��l�q�;�4��]Nλ[D�l��	��ڛ:�j�b�^�z���g��Vr���>�X7�jvT�����t��eD+�4����񣤆D���0��|4��W-�m|��'ZA�H��f��X����s9l�*s9 �9�q�b�t�66:\`M�s�+y���k��Yy;/��r�w{��F�&�l	B�1N����#�s�̬?�Ew�9��;�j������ZY��7x���^K-�v�����*m]��v�'r���}��?x��G�'����$2Qة�Nؽ�s	Mn�wZ���"�y���,�jm.5%t/P*����춗��+=��ޏށ?9j.��}�-ߓ2�=-v�
���KNdt�и+Քqb�iH.]�i󟫧�s�ڑ?{���[-��{��M���B�+�����]����gDZ�P����aGw���7ky͛]��{���~1H�ث��m�Y|cKU�Cݑ�wQD�,�K!W^rm@���hV+���e�Q�+��>����u�(�+߻s��oϢ�Ǽ]$[�ס#��x����1�7^TQ�Ǵ�wx]e.1����'
F� �w�T��Uu����=�o'y̫X��s6�1'2GLv7m�q>�z�ջ��2\3�[���u�3rnJ�1�c$�%YrF�*ͬ66�U��Ƨ�Xň��\G3���j�v�_m��5�������y���f�5�H�\�D.�j�`ZS#�;��r�[��̾�8�jz�a�v��٢?8��w�J@#=b<of��]�4+.[<����e�Bѩ�p�}�H��%����mW�;�#���ҩ�Z��g7;����a��k��x�Y^y�|�vA7sg��T)r���߈�q_z,���塚Fݑ�T�&�ܰ�M�i��3fCW6���R��6�J��۳fw��rz��Z�3&��]��ӛC���6 z�yS�6c��Jϝ�������{�c�S�����L�}�5�	f4����7�X�����z��/G1;�6:�~?a3�w<K�
�����3��[tk�	'��4��_�C,T�B���3v�(�-�*g�*2�6"9��$�#�M��7���ڪ�ȃ�2��]���-�7W����^�Ŗ�x����;�W]�A�������z�J��O �V|%֦u�f���޼ɔʵ�X�^u���$٣��%S�i�uH�\.fo4`�ﻦ�_wI;��y��n�ξ�N|�J�[��W��^4v]�4:�eF��KO�Хس4%wT,��W��]5s6\����w6,�{����Pq]���uҽ�{�M��^�N-��d�[�S��}�T�>߸���H����m{���I�"�qh�G��
��N��I^�˚#�Jz�;wQ���kbFT�O��ທQ-��k)Nŗ�iބ������37G���&�)�>�3O3����r"���)��6��^��*�	:�,H$��E��%��y�Dy��2"����u$���Z�A+��_ons=��e�����\wipH��)�ހ���:b^;Ӷ��vU9�$�ͻ|w&#�����t����؄���U�>�3U��yW�V�妙hj���ˡITc�U�r9�v��8fq�<aX���n�a�7Rk�k�}��Y��k4y���/�~������|��zNQ������e���8�v��&gR�4���݈��܄Q�b�qq�5��A��,9wGU��{���|��A����:V�jJ��t�����X�<z�l�U�k���OQͮL����&Gu�Ŕ;�If��XW�_g;��{;�D�+�P�E��W�ffN�^���ȩ]^Сo�NÝ���!�x��bʱ}���i]W`z�xhv�Us��f6�s��sX�)�S��m�{�5w:+M��'i�������m�~��"��0i-T1S44�F�a���2��L���Ϧ)*1�j��t�]��y�-W�ʨ�m�Y�xu>j&����`����ڭ���o��u$Ys�f�'�Ѽ��pr��«���N�2)�n^>��\��2����!%xl\l�t%���M��0x~L�T�1��ntqz��~~�1L�)���6�%ݤUnߙ�Ȅ��ٍGc*�za�wREY8��UNY&�hS�\IL�E�j�{9�#�����X�M^X�gwɆ�ٺ�K#rI9�K�WK=����fS>���S9`�
�2��zzu�N��P����m��+:��Y�g�_�	~y��֙bw*�9���e;�N�
��H��^���qj|�&G�v[`[��N��|\�老��n�g3�e}J��ӑD� �a�;f��r�-U�6nR\�M�r^� �����ǹ*���]����Q��&��k���q=Z1Z�y��� ����� �k����n	����f���+w�;౧.��d`h�nc&^��׻)��(��k��]�����L	��zt�NVJ�;���^nkr�h�`��?�skѶf�J����z[J�t[ʉU5��K[�s2�pwS��a�vy�8i�|G�}l=iLt/�-�t՘��$Q|�%��|-<�����o�Zǖ��W��}B���G�Z;áa��1�8:9k�г;Uf��<[%FX���lL�-�2�d��FlN�f��}p�W�~�Kw[v��U��7ح�9S�N\ۛg!񺓙m�$�8�!�c����S3�|gj��$�HH����ݘ�f����Z�� n�澗�nc2��q�D�$���
{�zmd���X֛�=9
�2���$���k�M�C��cQ�~���kx���k[m��V�ʹ�~��K1��)��{�]����+֧l��n�j�٘���,k}m��e�ܔ�;_6�T��bf�<6��D�3��X��L����=���G�ze���O�}&�Ad.���Ɨ���D�[yٓ,���+8ŖKuʍ�ζ��5v�u��[�2���vӵ�l[��T-��e�S��w��讏z�mY4w��o_ו�ufI�|n�ɉT=�G�6H\y͇��K�C�*�����U�Õт�_��8���Sj(5��V���]��5�RL�k(+��9K8��a�N[�sZj�r�ܲl��a+S��G`���͝��㻻<�䶰�!3�ku�mν��hVwZ�����L�F�-+�}13��MI��ym�y�JM�Y��8�ڌ�섻ӄ���a��4�A�Pա�o(��t���nݚzvkD��hY�.�K�٧�0>"�5�i=4z�-����=�������C9K��nh&�
$�j��ykx`�]�u���`Ȏ�6ڕ�^*��3�����V��U�5>T��f��/3�N�;&��<.�9K���{�j�YP�$���ޅ��V�$N	���s�[M!*V-�:kZq#W)s�8�<�̕r�=���eݒF��9���ޙך��.Z�R���z��s\�cxD�u���G-�!m��S��8��]�`�Z�	���4;w��<9i����"��
��P�z������w�ltd������2��v�O���h��m�����VC����o�,��Y����эٷd�6�<��Ur����ͬj���7X��b�yv47�$��Z�(�L�>��ˎ`���FUɹ��}]�z�d$�r�k �G�ň��NM�*#qfض���$:����@�gnٓfBZ#0l�^oXvE2mnwo8�����!`X���ͼ�Q5��pa�e�Ȱr�GQU��Z��4�oj��b�Vѵg`=İfT-ɰZ�I�S�:��N�_+�k��֝6T�bW{B�g\ؗM�����ۛ[u��q����*nogB&=]�g5EG��vr|������A�J�s�݅�����n��TI�3PX�K�j��}79l���4��J�{�Zz��k$��+�y����gc���&���m,��ŎO%�B��$����eM��_�3[��-s�x^I#P��	�W7V��U[j��.�>7�Xl�*��	I�!N�c���0���ʮ�	����"[X��r��X�b��6��Ri�3�!J�Т�9)�yԷ\{7�%������j2R���"s���^��9_gd�[��n�I]Ҿ-��36q�b
�;GoV
Ȯ⦉$a��ĸ�hVMiZ�h��
Xr,S�4�-ݕ3�0��pΥk�2�w9�^��*c��j�݂�����d��B�e�"���%u����#�f�;+aч�3���Yǒ�/M����1[���Q��6����Ůw��6�)�2���[L�TI���/ߨ�,�P���lh��!c���Ϊ�i��61lj�+f�kE1���~��l�S��EV�4�QE�8j
�����:��D%2�RE˵c�ӧOO����q6��[c�&�gUPDj�����E�6˶��<�*�"ּ�>�O�����ht�h?3���5IQ#L�9r��kh*�Zu��/0�0c���}==~��b��v5ch�ѣMi�j*��E��?6I�m�ETEi#����zzQ~}፝%��d��(�E3����k6$�+1h4j������z{�[m��F�"�j�5N�1�4f(���s��"�"�H�b��������}==��p�M% �A%E:��D��٤ߛ��DxX�)��c�N�=}��Q��d�ZDT��\�t5ES���Z��֍��mlZLU�:�v<�\�kU�mgkE����U&�"�Ԑ@�?� ���{ޝ[a�T��Y���I�vڍ�3����ݴ�C�����͖��[�ob��Z�"����P|����� �븉����G��X�7)_UoV�p1i�b���{X1l<���oV�S@�'z�ЖX	h���d��^�T���̆�A��]�x�XOm�<�B,�A�p|�
W8��f<��	dyW^Tu(���Q[[��0�_�z��p��`�Sr%O���3���Ƌ�`�ݷr�-�K\gwU���J��̗V��8,�<�|�ؤ�F�tO]%�j���mֈiƩ=y��3��
�0�5d�3;X1�� -�ʬ4+^/�xs��'����MK����}B��ܰ	0/6O3��-�خ����v���yц�3�}ϔ\�l��	�J���>��t���L�����lz1I��;zznn��="�S�67���v���U_�\ڔ��e���a����O�x��K�X�Ԟ#y=c����l��z�������j�J�'����;u3H:�����������س򱇴��D����㾱~���@V����@9���$E~�'�l�}~�z��@yf�T��J�M��L��nJb�h(���w)���$�*�P��A�yeӽ�Mĳ1�CYL������?@�Y�����/��^PM�"&�W����t�������o~Ks���������M��h5�{*ŋ��̊�/8	[K�~it5�'6N4��R��k�yyS5��WS�)}0�d9�UH{5":i���&����s��xU��5t��9�}R��1�v�V%�e�0=�������o��vD�����*H���vv�ޤ�Y+k�s
��{6꽻���.���M���;=�/5���g��%��V����+���ճ���v&��8w]�`��!Z���Zm�v}dW�mj<�ʅ/�{[9A��/f�;�i�;��m}.���zǦ:�(4����l�!�z���$ps荃��	#�!��0�<��'�hi��|��~fYQ�z�A���/�7h5��o���.~)-)��=[�J��<3��|p�5�w�9��|�E��U��㶀�7�s:�H�0��޶k��T�U]�#����_m+g�f8�0F��e�B�qLv=���b�9|Z{&T�^N<��.�˚j�C�{�.)*#���$m���j��u�nu�#U]�����`���F4���*��������V�=)@�Ҹ���x�GՖ1�B�d��؆��3}lx�D8	�T��"<`������{�Z�3�S�e�s7��Tt_ۼ�~���|=aׁ���P\c�$��x���geN��"7+�\]ݑۏR|M��?*8Y����g,_E��}�f'u��y|ط�0����1+h� ���C�C"��h«����<�)�bM��F��a�������N�*uá�=�]��Ț�g�I��oua�wg����p31H��KTT�`T*-�^7������L���3�4k��a�{�m!s"��ƭ�nByR��Y9CU��/ԗ,(��n)ޯ���z�w�@S.;6��ab"k�`�z�m��P T{λ�.���
���;���_=�;~�O�gW23a���\���^NN.��
�d��0TLPg��zkm[�3n�":���Xk�Z��� �խFe��/HH&W[u{�k�:��+�s���2�6C>ثm�rB����MN-�1�TQ���	�m�!��� �L�gT��p�Ele�L^e���`��������U}���J�T��j�m�>*E�МiM8v����V��Ϣ����93[�X��d˳R�ī���$wU��B
f��UF临���E�Q'����:�<�OMˍ�qX	v�Ig:/��d6HЏo4%j�Mњ� E�'�N���6qn�,�9�y�F�%|��<��ӎ�|v#ް��#lZ�����+�e���g��9��c.�9�s;EM�_D���bQc�Bi��Ӑ����>S�'�gw&T�A��I̯�����_~�avw����3r��:͊k;eW觍�5ʺ:��]�dw��C`Qψ�Vz!���ܹ����ӎ�<gvqu���I2]}^��}9��!�����f��oz�d�f���Ȝ��k���>�}��8�-�4�J�@R�仭�L�Z�Q�ٟ�c�f<��t�Y(��pn�1rl7Q�7�DP0lBŗ4��X�/+��l���+~�gX�۳Fx������3�'�o��Ǉ�9�pN�	ܰ��kZ��Й����Bt�����Y��}���o�<ru�>�V�`���� �-h�lNU@w�q��k���c7_M3zC��,�x�jU1h�MԁU#nњќϒC	�]��W�,�=��_퓀�����x8gT ��u�!��TL�,�ۄ��o�����X��	ӻE-�R�*w���]�cP܄���C��M�Kt��s�s5H�ַ�>���v��YA,ʠU����Z�L8��]wJ�owsۈ��	6�5pff�J���e�����^D��I���B�f��^F��ָ��b���3����B�ЖB���U��<�su�Vz"�.w���q��v���G4\*�k��04sR�����EO_/"r�:s�C1,�Eޡ��Z"��c�Z���خ�vt�혪m9���6V�Ϗ�����Z�$����5g@�kkf�R���"x��e��c�h��M
!.v�v���sM���w��:OR���Le���*���"���Y�o���o�nJ�v_�����=R��O���\��s���9�Q��\K�h#!���ǽW8%5�N�/��GVS�dܥ�B����y��6T̷SP���r&�D��<|��l�:�Rݺ&�vv��-�G{z=���Mn&�m��\@z��͓V�z��0���Ҳ�<��si��i�}��b#
�MSaZ�����0f}g�
q� 8�3Ið9���.�`��ճd��ι؇���u�,/��v���$��;��y�"�<��>�g?7~�k�����'�:��a��}p֝՗���@��Tϗ�ز&�I]!�����������ā�NgSj���a�)­���%�U���]'(�N<�=t�!�n����
�v�T��-�u�%��_f!E[��'�mَw�#%^����ި�ڪ�n�'����͠ε�ɭ��VϳR38�U�
�iKh,��ֳ����C��L&]�*�Eb혱LՂRڸ}Mr)f�Q�27a,�)kk�j��l4Q���%�g��	�/i�MO���ǒ�WRU�OI��:V�ݲ�(�.��w� �Q�a�wJ����v���)]��v^�T�+�[�Bq�X\�'Vv��sl�G�c�AWc�t�b;��ؗe�E�fK��4�H���yι�\��)sk������ݼ �E&̊����~�����>�bZi�J��[�Ċ�U!����'�V͐�|Zt�����;���<N�9u���o\��o{:��A���y��щ����h��ڼ���,���p��3�W�r�U��V��Љ�B;��^��Ͻ]��2��#}����"���{�	��:���'�{X4;f���t��U��b�sb��ہ4�;�ڔ�ɜ��$C^:�ݺ�����$3�m�m�����]��k��VJh�t���wU���J�.z����]�� �����j&��{#_��ʨS��(}p���%���V��r�=&�$�t^���Yw�������<Ց��t�q;��g��l�fE����*L�������~ڻ��|#-�;�=Z�{֞��(١^sA�]���v�^��͟+]-����n��4��aBR��0�@s����&��_�h=.�/e��.9[W�*iB�C��s���֭�H
-ov��Kv6�	�A�H4ʄ]˸�j���[��^�n�-#_!�B�	'Ǧvf����=��n:a�7�z��I��H�+h����^)���2���9���F�\<�����Sr���C1;ӎ]W��;bjOq=��^]٪�CF��KM�Tͦ]l5�K�z��:����mL�M�7�X�3�gT@�"�Ԯ/�`��.���Y�#�`�����&" �jS�d�k\��\�@�0r���̂Z��]u��>y#�f�Ѩ��w�~�Ȕ����U^n��>��	=,2�K���y���a�iF�Lenϻ��r8բ����7P�֪w���e3�؊?�}��7�̼��(6�IN
��c��������Sa��fn�+��8I��aa����/�(�n��ܸ�;ug�bJ� ����;%B�l�1�+�8Ѯ!/�DpQv ϩ_H��$�I�N�|���MS�k�j/�w�v5�d�5��.S���1�v�E-�;!B���8�O[�̳uf��7�Z;�ϰ���lM�����T�s=��m��7}�K�>����;��E����*Μ�".�u"�Tɋ�̸��y{7c �xt	雜Ag��}vMJ�he�8j���yk~GЯ�H�u�,�=34s7ׯ��R�hE���S�P�������lYr��3����%=��yP���������R����+���D%�5��Jj�:H��޼��6�C`O�j�;�9�!Mj|=���M~�[�����r�J���N7tF_��7H��?�h�����zq9��Y?fm���3���P����eks����g�|WO��1��ԆSߨ��&�ǻ�=�LOߖ]�[	H�`n�7������5*I��`=����s�˵�Ρ��~�(r�j��ʧ�=B�3���	�����	���5��8�K1i�6v<d5���Ji����W�s�_��3/�+�%�y�����;��xۼt��N��5н�'��W�=�m��NG�5 `��
��J�mS�je��\��n���+a�r����{�L���1���z�H�U�۹­�u�H�̼�d�Њi�ͷx���j���C��]����+�rk���+ްk^�����ʳ�Y�c��熱��d�-O=xerzFUutXf�����u�ΏK��޼�p�ǫr�gJ�����}�_4���O�zx�7!�mE���ܜAǐ�AM>}f�D��s��2���R�bv��{3He=(
�L��Wظ�����u�5�w �&�@Ҷ[IF�y;�%,i�M"F���A=]d�<��iC�o���e~�4܈V.;�=fr���a�a�6%�/^����="#g�^��;�5ŅGS��IfW�͇�9o
�:�����%;'mֲ[�\Тo:���~����$��7-cVH�fp��{P��F�*-�ܸn����{p����7�g�c�{O2"Ve��dSd�0m��o�mD��"F3���U�.@�h�����ՖO�e\�b6�6����݋��w�*e<���֍��)��#+g��#�6 ��NT��3�w��8�� ���;F�E����Z��>�2��UB�ٿs�ٴ9_�y�CB���g����ʜ����T0�g�a���xD�ژ�+g����1���Y��q��kE�G��Ѵ	l�#�,`-c ��9�V`EV��j=�}��7� ���PPA}O�����G�HPA��q��A 3�=��%"�&(��!HAD�%H�%T|� H�(	 B
*>�!�% ��|>a  B � H D  @   @���   �  	  � !� @@ �  �$ (@ � 9� r � !�! Z!@@ ���@!h�  P �U� @" �C�� D�	A( ABQ @�4$�	0 ,� B�
 np��H��J�D0�4PJ��C*	I 1 D04J�PP�@�f B%EH�  _��`�/�Q�:E�PD!�ѓ+�[����6���P�R��#��H�����&|e#�%��Q����g#\v" ��8��s��v� ���TW��@�F���	��kw��x�::��._#�.�&����OlI�@*���ʳ H2���D��D L+B,� BJ� 
�*����D�P�HH*�@�B R���R� R H� P�" R H?�D] D( �2 �  R ( A  L �B�( A* @B  ������JJ��2��K ���JH��0! 0��BH��ʰ2�2(���$� J�20 J��K*���2�� A(2�I�`�~������ 
D 
D�q�4-z�����C!�8��u�TAEy<�З����"����������(������:4�)�1((��DW�� <[T�HQ��ǂ((�F�������'��x�?��PҔ%��ƃADWI��n_���(��i)Y��l5���	���u0_��$(���r;Q^��,؀�=~`��bNA-�ۡK4߽����Q�j���pH����������Pc@�DAEw��f�r�"
+(��:vU�͐���d�MgD���f�A@��̟\��|��AT�"Q%HU�(� �R	��QD�R���*���U�U ���J���R����)T��$[�UUQ�((�J]k�%*�IIR�Q�ҔUT�)�
�F̡*��)DB�"��!A^�"����	P��QRUE*�JD��*��J�BJ)AD)	)$$J��UQE%$���)UI
T�JII�   �ש�Q�Z��9�8�i�۷vtn�v�U��2��6�
�cm�Vl���i���wMw:�$cN��Wm:u�]�6��T��'U1�i-t7R(��5@�H
�D��   �!B�l(P�"C��/cBE
.�B�#�B�
/c!B��W�z(��{ꌻ�MC�Z���:�U�M�f��w0��h)��ۙ7[��wSv�VV��n�]c
ٕATH��@UUT��   .�kE[+���t�mf�:Y��f��[nɻrnN��[��m���Ԛ�l`W@�ͦk �������1(�V�nؔ�1�����I6��   �zx5�tݨN�[�uJ�Ҵ��*ݝk1��M���+�@ZK QE�f45���A���B���"��0�R��ABPB��'x  �� �� �2�RҘيV��B�j�
+Z�%�UAl�5R�AeTe���5H�b%R�T��)HU ���  ��RT�%@(��U%0UHC4�64����&5QT��aTU2���C-6�1TU*J�����TRU	w�  ��
��YU5��aR [m5
e4UT lA@ �0�5e`  6S  [b� YJJ(B �
���U�  u� (��� �  
L i  ��((h� ��6��j�  ��  l��Q4iE
)%   g�� ̌�@� ��  R�  � (�  
�� -5 
fS �C�*���Z
�T%J��  e�  c, ��M�  �X� m%��b� @ά Ҁ#�(&�  a`  x���R� 2 S�0��� 2 M�OLP4�  E?�&�  O 4�P   �)PLUB  f�Y��a0S�J$�B�N6@�HAXށL*��L��TD���r%�z�� <<6�����1��������L`1������6��cl�`�llz�?���/��(�Q�4�A,����K��� q���@��L��p�&�n�Sp���Z�i�J����3r�*���� ��eی�5���WVl�L=�	u���:!�R�a��"9�u�V���ۉ� �K#(mI���,D���Tn��/c&�.�
PU ���O.��B�c4Z��qֶ6�TJ��;�R����� ��:R�l�,lK\Z2X�]�-h4�h��&1�(R��:\UotC�j���kA��r����Z Ae�$�5p��'BmE��C�RcL4�MR葦-�%���!.k��,�� m����"N�mӁ"&p���Jλ���"�_ch�B�/~���$�^*7�4|^��7WM[yw�hȚz�>q*����]d`#���kێP�k�𼣐��5X�ɋ	a�\���#m�cr�h���x���q#�R�4��ї��V�
�r�Q{�Gfܒ��+P[K"zu�klD�og�1^��K-�("�F��o!���{G4�9����S!�֦�ي<lک6�kov��6�PA���jB��a��r��v�Y�����M���(,-�v��w&�a`�Vem7,�a� Ɏ�Q�JY�p��c�EV�̦6Z5[V�Lf�c���ȵ����BY��2�0��,�)t�����1N֗x��0B2�Z���gZ��
Bf�R�b0�[�ov��ZmA-��k���r`@k��[of1��"�"Y۠U+/ ���e;�f���+��LE�fKQ
5-�6&ѡ�z�6oa�N�u`)�7Q"�^�wXm��D�rF4��=��7Qn��ʽ�5���h��^�t��	m�Э��цU��QQ�~6�IW��� �e�F��D�4i�2J�@2[�
X٢�U��N�ܚ��C@�u)U'*=�t�kI�̑���[�QG�k��d��vQDA��L�O1`	]�Te�sDH�.�
 ة+�@�ʲ�J��.�.������˰��qێ�BѦ�C�q��1�Gj�Xȼz��R��g09�/a)��b�m8�@$N]e�T�^�aP�8��ɉ;�̗�i�(Kכ(K�R��f���h��0bw(�����3�-u+�5�p*8n^�w����Lt�����{e�k!Ul�v��Skw�G,�=�F�M˟Ep�/6Cث+hM��n fT��Kbٻ��Y�-��Qv
ݢmb�
�mi���!n�.�X+V�)���u�÷���{5�/2��̲�Bز�h�v�Yu� |nZ6ݰ�
{{��+ݙtu���jh���l���Ԁ(+#�X��QfV:!e��FB����i�]��X�e��q��䗴��C9-�����	����{�Է�v�%�P�%��#�6J�fe�>�R&�;�t�Z)��;q�d����ejR�9wX����{5� �3"yN�#u�[Y&�ͺ�;�6�ը�*��z�\���Akkj�V%"��Z��^�ef����2^2q�i�E�w�*�{#�ecos7��YM�yd�j!N$�,�p�Uxv���n��a\�|	%�OJ[M^�f^O��6H{k����gi�b[�O�ڕ�����1�Kc'aŏ5��ځm(��I��oR�h��f
Nmn!�*�j}��ŪnmU�w�:Ğ^-�$���~�z^M¬n�d�BۛW��%DMN�W0�W+	p$��4G���uA���
�Џ�6��+1�	��t���&���T�,8v��Vw�X�ܸTkX(�N�c[���=D��7��tVF��YZa}a1�JD��ݻi�wcu;R�Df"�l�ce�ʳ�j��v��G5�*�H�;a��`��v�!s6��h$n0ݼOm�5m+ݴr�� V�6�<��D֩�h�N�����bf�rʽn<�[W�eɍF�E>������q�Fܹ��u�X�$�W��Y�w�MZj�݊�(����]�W{{1��ٺ�dˈ�Y�F8Uݬ����2��T~�� U-���0,#&l�y�t[��$�H��B<F�01���K�lC`=�F�0X�h�X�a;��Ɉ��j�S_Y@�ܹ�#��9wI���F��&&ȳ[`�v�IMO���l�*�5X4� ��-�v��{�p%y-��R���廏.���.A,�jjyE4�'B�b��&���tِP4pޜ�������4	�<&U��'�2`���\}X��&Aԙ]��=b�ἋU����z
c��N�$x���`�OP`k�"�b�k(�vЭ)�/1]�e����h�p'�⭦��.��D�����*�@čj���v��;0d�@q=P`9l��ܷ����vCa�:�V��:�Q/F��]��P�R���>l=Jܒ�M��Rr`+>9I�{�q�I!Qf]ʷm�ҏ�*T�̎����`6Jt�-X�4 ����,�ŀb���c�Mh��B)SP9AV䥷���Yr�@���d�׷N�5�L��n-��˷��^���2c�N�[B���G�����[��a��`�kh���ɢ�4�ZŴv���lYc&��ib76x�(Y��sn�lJ	�j^�y�D32c�jf���t�D������b��q<�k��,Á��{�2�F�+Ձn�,���m<���4���#e�Yv˕�I�f����Н�e�Q4��n�hF�E��Vy� ���-by/�-7SSx�!z���0�6ٔ1XZ�9bܡoE5F�[�:�����de[�j#��ѤA[�
]̴�m��°]hR�������Ɏ��B�n�;-��4�Z 9DV�B9�C�Y/>��l�R�D�j�e$fR�^���O��/��s���s��
U��&���c6h�ٔmKw��E^ͻ��LnMWFf���
���A��!���˻Mk�WL5�cD;��qnP3t�'$���� �V�B��Ԑ܈]���"��KN���̦N\���)i7�̥y�HAn=�
�{Ke*b���ff9Fۗ��/vH�n,�Zoe��t1�md�
�SZ¶�e
ۍX���n�6㵈��k^SS�� U��ªѫ����8�������3Dz���l�e�i������-$i���q��,����d�[�kS9��b��WvtLw�6�S�^��rf�7���kŷ�6̺]�K���s�^^	�u巑@F�(Z5R�9y�m�����a�;�X�ļv5�D��W�|5T�W
�3V�1�r�k͠P��n���y�v�����AY�l�KLN����6���%�����l�����R��r�ڒ���)�J��*"X�5�y��Y7��^�)7� �R�H�Z��J�mRU@��[;)ԗ��u�[_Jŏv�fej��[��ù��]+hR�*#��R�L�Z���\Y�ۃ���t0�eb��v���6��+����xa�d�D
fm�eû��fS*aӬ��~���Jf�#!�\�v�KD�ijL���f��Gq�dl�Ř�ȭfT���V,�����G1�+]�ܕ��/qd�8�:X� �.i���������l�@�"�u��a ��-C<zI�L��[n���Aw�'R�+��mnGX �M����!OvlL�w��c��h[��:c5E�`�:z7:oP)�Y��2�����G["L�R�l����Md��%�%��a�{�m�aMki;N����*6ޚE��V�hVDr�e㙮jXT ��ŧ+se �-QU���ͦ�u�nw-�;7�n����j���@`槙L��X��0�(�5�F�9zȱn�iJ�}v�1\���%zh
oe����.��R���[�v�RɌ�6KY&�5�ԗ���)ط��"y�Enn'��
��-9N�ǲz��u-
w�~z��Jx���nH�Y B3am�z%k�h7�Z��8��5m��w�z����m"�IJ�ն"8�:ാ-!l��n�ki�׆�/h�1Y�>�^5o7\��2l�����Y�+��nd�$o�A�p[G[�������4S�;� ו��Ʃ���v1�Iy@&Ӽ�4$飚�ȧ���)��4�B�ּ�ՙ�����W�c���LՁ�xT�p���S���@l�OC�&�a�Ϟ<�jeD�G6�f�ϩ+u�[Ӱ����$�F�@�OuЦ*V9 Ҳ����|�VC���B��WH-[p��]\�%��zh`/L�w"�mGFV�R�nVm�x��n�ҭt���Z�	a�2�n��e��cnё$/[��bZ�ۦ�ڣ�W��^:J�Y*)���7��n�P�[��陭32�-WMR�Gt�N���8��b�9p67s4��ZN2^ט�]��l�jyb�V�9U��Lʨ�c�r2�fu��($�w/��i��CC�	�h���wCi�f�����Y;�R	����m���k�B��U{1hiV��V`T��@Ȧ.,JZ�N�OD[yr��F�h2�d���JSe�,R2�LCfKo)�mT�X�m�}&Q˵F�f�����-ơ0M+]7&ˈ^kY@��swG�@�6��2�Z.�Z���P`l:7t�����1F�f-R�鎨4�*SŊ֊5�(��X6PS �-�KV����E��+.�ԁ`ֲ���h�LC]	��<I�a�pAqy���fK,�{&�ˊݒ V��:��{(^�h,橪�ڑ�m�'׋N:6n�hf;$�+Rj\��0���f]���7JR�^]�e:3$L�3{x�^���9��yC
��L�;�횹��)	&�ױ6��Ua2*�MZ��j���j��Ͱ��t��Xɵ/+c��sR�Ƒ��[K$�Qw��J���orl�CJ�L�M�^^�d�TcY嫘:���\�y��uA^���xU(.M�0+G�U�H�p{��F��K$۱�jM��S���ť���EQ�V�L��Nn����[����4_ɼg(�D��#Ջ4K%�l�y����%%��*6�\3˫P��Nb��F��Vo��l
ɓN��K��M�X�-�jݫۥ��ے���Cq������j�e�4�Ud|F��9���tb_FX��F[��⣔»̰ y�|wp���ܴ��}�i�x���1c���P�Q�	F��&|p"�m�~��e�j���.���[h�*�����IjWw`�7`L�-X���E�ٔiZ2�cۧ���(��#l]Y(���8t�tMӷ�X����y5�0j�tn�R$�&lHG�SN��X%�Y4���(&e��vǑ"m�̋�-u�.�(�*[�m��%J�J�HR�`��֍�AI-I�ə�ͳA/� ����h&C[������%����=f͗6�A�B���Af��k[ݧ�[�Zmn;E��7v�ҽ� �.#�Һ�x+)���;�xr!4*ŭB�,=j���l��̩dT�T���x�D�vhX����$��r'q�Zѵr�kٶn&��6�l�3��`�m��cP���Z凥k�8��0�����iE�ȶ����Ǵ)Y�v̕fd�������z��7�D��v����e �V�#�nh� ��u3yaʻ��:�GA�ˬ�p�cM)�^����m �F��;�h�g7TK	*����&*j��D]�e�X$��4��(0ܭ����c�wku�k�Z��MJv����bX�X7H�2�˵�<���e��n�V\����aYS"��I+��X��"����%q#��3�dӋ��Q��˳M[/��B$݉�w���l�ݰu�4[T���#.��tPͲ$�h�iJ�����R�����f����kh�����������-���D��M�;'ֱ�.����H��1S6F�GDhF*T�7�dp愮e1.� om�u�P�p��\�ejP�(O������Z�mCH�q�7R��H�@8��Il�ji�1�i�\nS�wEnÂ�P���t�h��J�v�Xc�V��Z�և7J��ڽD�^�i�Wx��]n�wO閍�TmL�CF\�Z!�#��T�ebyt�T謺f���T������cE�W�Qf�D*�i��E����*5 ܫ���eД�1Ҏ3�U)�XDU���P+eJե=mJ.,�Au7�e�i �a(�p�(�\{xa�-��x��!�GXv�q(JV7u��2WM��E�5t��C����kI��Te�rX	�j�O�(�����yy�Ɋ=�\�'a�6�ȇ���z6Y/�sTx�A���n	w���e=N+&O�U�Rm)��A�����²�0YZ�Rbq��
Ӷ�U⤐���Զ[����b��X��`��V��SLxM���8�Ղ*�BU�" P��(������F�n�M��`(�/6k<ZZ7�&$�i�[��F�#pl�n7#���H��/M�*��#��e^=��u���p풣��{�R�)���r}��wI/cHL��z�.	{�NM�a1KѶt6#hwq@̍���ަ�Q��֘ka�C*Mb����2���Ŷ]з^��Y�8v����@�:2�d�.�5��(� TC(��nm��ז�TB������ng�pԙ��c��vm�E-���ft^��O	 �7�TJ����~P��/-�r�݇�X��
Ž�`�mT��݊����s4lP*��q)-��ƭn[����Z��B�0jm��`c-�r���u0l�̔��ܤ,�{`�����!w١,ѭZ̦X²�}�q�v%���w^5��(>8�є^*�Ƌ��������\���&uuS&��V�]e�l�S-��#�F��Vvw`��{xt�T�L����3���b7k�'Q�����J-N�w4�w�OgTJ���q���L�{ڨKN��EV��7����I��2�iMF$w��]�=\��я�8�	JĦqwp�c~u�7����Q��R����Dq���Ր��z�:�}�y!��/�DWuk*J��ԛb���Y�䆫����j����j�r�-�(1��J�)��7�����yݥ�E�XA���oI۫�u�\�co��U����w}���T��9��^!u,�Z��B��i�e���ήT�vڼǧpF)WY���Ue 6��ē�Ɏ��w�pj���zn��%�o+$��tu.O
R�M�7�k�P��.����#�]��MZ��wLUԂ��.ةo�fVT��"�A��T��[_D�0�;�V���w
{@<�>��7�;E������������݁Q�����A�%_���leX��Q�R�!]���hYDn��k�,V�"{�V�M}ۜ��X�E�y�G�ݟk��]��s7>ی,lr�
�n�S��@ʐ��E� �Rmj�e�K)�F�V��П9���j�1�o��jXx@k4fh�Q��w�\J�����S��D�_6^�Mn�A[�x��R�X/U�,��t���j�jV��x`s5^Й�p��QK2��,V{o�Gם��]*��0���F�HL��h%j�ݺ�Z��E�P���у05��wl�=��[T�8�EXց��{��G/��9�����_˨ҹ��F)�af�;M��\Dv��������ǂiC��n�S��\w9�s�9VCc8AZ���0[��4v[C'pb}c�9.��[�À���;d��cY��g	��v��S+/�2�L��*��V���"��r����u���oQ�_K�]45�Xo��d��-��.�|ͬYu��䱕���5���7K��|�ze-�4u��e���UL���ꐅ��3x=���d���\��Q+7O)�Ǻ��-V��1V�={Y��&\�L���o<(*.��[�h��M�a�hn�$��kiF��i�nl��v�c���IZ+ȋ��98ٗ���O�L��a������#muN�{�OpM*DLM�,a)59�
�BK��HV�9G�;;�\9���hԮ!�prw�����\:����(���7�|D2�	�r��{���Mu�s3����5��+�c�=�<o$pЩ|�vˣ ǹ.���䝋�)J�W٠s���j
5�e�+a<eh���u�� ��;�	p[���$�S$�,�X �X��T�m
��f�+}�WX!l������*�n�D-Ҋ�s��V��3�=:�t�vǥ>|NV�`+u��:�g��2xN��I\8�ݬ�][�������b��{��L�KX1��n�78p�U�2=L���*&5��ʏFvu�S����eEd�=e�.³�j|Ƽ��^5��y�t�F�KAb�س���f�a����̷+���-����.�f�c�M3tWU�\$��#�M���;��%�ްrugu�'i���θd
󌖵��Q�؝[IBm�h����k s��˶XQ7ɩ�%��*P9������P�j��CL��q�")�zq��tr�Uʸ6\o���n�|�o+Dc��ak��W�t(�tP�� VͲx�4s�sk]Nz����Ѣ����1<9m�v�Č���M�_���U��ރ/�. ���N[J���%�}f4�8V=RU��Q�+��uk�$f%�o�;w�>�_c�����f��b���S����tF�\{&��k�ң�b9�}�i�ޕ6�k����8e}�2a���+Ӭ4�N�*[�Y'T�7P�֨_N!��˺��@���.�lo�/�V� �RO��u��%'{���P���v�~K�Ρ�뷯��@�
�5s��1Hx���5��y�I5[&����p}D���-�}��mVau	�);�Ю��_LÊ�y���;��O=5��p�O���7�f� n��`J�q0;�n�J��_r�t�̓E�2½��ϷD��T��{�sXԷ&V<b��?q��54u+�:�S�0�Kݤ�U�
���}aomw��kj_F�:�I|J�pp������#�#yF�Tü6�T���7���rXF�4�Η[���-q�T��Gc[�v�\��)�;R�we*"���ǎ�f�W�svh-�丸fS��v)V/��UȀy�q��O��;(��et��oH�S�uv�y[: m����.V>�7<��UCTڥf��vCӵ�0�J�jЩ*�v�V�Ӯ�Z�XӨ:*񉇳��ۼ��ۨ�Pjir|�r=�(.}\�� ��w���Y���A�ĕ�$�E�x�%V�Rp���f�&�Z�.�r���wd|���X<�������|����J��Q�8N�Z&F�H�j4JV�^���{�!a�m������c�
�1Y"�3����n�A�P�Q�*�.Μm٦�<nl��¸l�<ÛCF�V]�<��.ki�̓yOh��课U϶	k�d�VY�U����&�[-,q7Sxm�oJ��'d,�j0bܔ),\P�BOu�r�k���K6{sE�9�-��C���7$��Bu���G���1�l\nt�M�zh-we��!�d�W;]�Ǌ=j��ׄ*)R�m�N�uVl�ɛ�ٮ]��e)�+��������}lG���5�g:®%���Rt�;Y�i��~am�x֭O�w�o9>X)WfH��f��o�X��բKt�Qv�i�G��ѱ~�`�FI��̖�ʊ<�]�h�����YvO���x���6��.�X�a)͜U�1Af*�qٺ�ѫ7�t$�G��[� \.�^Q���=JW7��h��2��!rb-��GiIf�ڥJ�^Jo�C3N�'��a�=�r�Mԫ�v~�wCÎ��;���S)�.p���ȡ�j���s�`4����E��y��*��:BI}bwU�U�ټ��&+�R���a��hR�����g���ˠ��&���>ٙ��J�̮��BdO�F��2�.b�S�A竩���(�򻅞 
c�8��R�n�"	ԕq�{X��kt�����)ޙ;����Vӻ��qMi�R����6��Iik�6����c��#Em�_P���Vm�jvB������;��աV��@hP)�ՙ(��k{IB���m@��
�9a�U�S+Nsެ�z�v�ޠ��ܛ���ܩ�i,9R#h%�A�;[����}"���Ğ�z� �Vl���N��u�� ��Ȟ�+3z��P )��k ����+����)�U��o!2�J�����#���˛5&1=����7���ҙO3����%>� �N�9���[�����k���u�{o�o�<�KF�Y�o>���9M��bd]`�p�[��6h|*�T}}����G��^4����q�y[�rJ��ܕ-=�R��V�
f
�l�Iܰ�y�������k��+,E�2�R�p��"�=�)g0U9m]<Y(fj�Δ�o醱:S#2gX���Wb�8�����b]���?�ҁ��+�:�U�l������S�̫�PrqIxB��l�gq�mm� �1������t�1v�w������T�Ĭ�Z�^��<����oR�ڙ%!ڧ]����5+0ƍ;νU-����@K7Λ�K�����fv?�DTf>��<����k��e�+5՞��%Xm����T;�K������N�@.{[�[�-�2�k�ŝ�;���X�b��>q�`�y�`p��7�g��еbu��B��*���m+��r� �B֎C`H��:f.���h�+^^Q)�kz�����1�[s�)b��64,��u]�!�@n�2�X[�a��Y�k,T�w1Џ�tn��V*֘��NZGOn�+��FQ0e�3�۰�פ��.��Q���S�F��k}Z�	�mL]L�l�׳B���N�����nh��z&�m�ejz1��:�uq������V���r�e��u���ncp^[�QdoIǣ��>3ӝ� �\E�|�X�������Ք̐vJ� ���*�R޴�{��q�B������;R�gVw��o[�6��U�J<�}ʴ@��|D�z��6�u{�����W�(`����;���W�Qf��)�Ej�ʾ}(@p�Ak���͊U�ޗ���C�:�.��[j�2��ͣHaW�.��/����Sї6���+��Zv��+F�ﶲ�����.��a�;%[����tF�0kwVvf]�#��Yi���}���o.�e�yZ �� L��3�5w�p���9��2���w6���ի�]���Ivx�踭�����]]�|y�X����S��VB����H��N�yTv��y�n>C{���͡ɽ�s\�EwA�@/O��mæ/n�> �T�� {(�^��:�a�V��8�JV������F)�wX�}�u�ɗ#J@v��1�ulً����NF�IR�n�b�Lpm��.������C��SV�����;��ɀ��p�3�Vx�#}��m^��� �<��W�}��>�������Zkk�+��U�P:����Z���6�R��b/2�/+OE�{{�nֺ$	�� �M��j�.tt��\��W"W2��QldSOV���[;��F�\T�Ω��B[;f>G��h+V����[Y�s��]�5�Õڸ��)wh宅���8���S{�a|��4^��Dv4�fsv�j؉W�[��C��Qn�|.e"{`2���ԆkL���1֧[#�oi4�Gt���M�/yA�yWVc3#1��t��;�m��R'tn* g1Ʋ��@��9��[�T�uǖu-ޮ���[�&��l���
�˒l6���s=�:���di����t1���M��ވ�{�9�䣤v���D
[Д�s�cj�(�.��7Z}(��8ӈ^&��W]L�.�r�5�*�����:�0w@F⛶#<C�K�5�^�xjl ��o��9�J#���C���WWwi�>����\�ǝ��E�;&oR�QJv���'fhg�oXcl&�J�Z^�`Ճ�@�yŒ9�B�+�Ac�S�d6.�!܅�D�΋,՞w���hw��;NrpF���,	�-}cG6Ge�?Y�?cl��t(��oSa8���]�s�k�z��-��p��:t�U�Ɇ�K0������ގg�ͻ��D�Wy���R�Q���j�修94TO�N�W.<�M����NY��&�x]�:�m=�qu>WP�X�G>H�A��_n�j�B���@��o.���
@}�nNr�;5�w�Fsy�HIk�wmY�]+��z�O�3��C��R6��'Yۇ"K)�WL�v��f[� ylYu�-��&��Hz�Ad��x�_r�.0��<6L@��)N윹o�"��U����)#�-�X���Վ	�6�b�T�d[��
��P��Ch��	:��W�m]�=��[;ne7�M�i�|  +��JP��Փ���%�=y|�pw�|�+�E�(���k���I����FZ�L��}��fw �ث��ʰtB�b�'`�
2�,ң���n/�T�KS��2�[�t��=���S�X9��b��cU5`�e'���V���*��.�Ӄ�t�\�$�e�vʜ�m��vS�9m1������ܦp�U"U�=���K���ڭ�[�Z�t����䎜hE;/{{b؎��{����#� �}�y�brf��̸������ ���'��/;�[=��ƥvmѵ��	�w]"�Zd.^��v�!�G>�f]�x`�Fb=�#�5�՗��"�wp��U1�C���˧{%�R��g�s�q���x*}��{�I�1��a�b�Y+��z�'�o��z��/�M�ga%�8���n�k8S�.�(��Ϸ&�2�$�t\F�]�K��2�г2�eE:<Vvͥ�;Y�Y�{�=}v��[&��ѨKӅ=��_C�> j6xSwjO�	�G�-�/6�ېJb���U�0-�+1��I[X��a��l()Ne[�]�p2�t���|v�=��U/������wb͗nh��i7u��v���v�����d���Aaվ<���M�aS6��e�9k�x�vHG�gIB��v����㧻2���gq젳�A}yϤ�e/�$�D�6�m*�*V�M8/q����H�t�*qx�1�L��w֫����2�_(�C�$�;�'���p���$�����]*T�ٺ�j�936��]�k�����K�Jt��\\w�^θ�N����jX�]�&>铆�<��'q��r�,��X�s�#���6Wm����g�9:�9Ҷ8�/��� ;U;ʼ����y�o��˔냅�<�][H�X�4v�j5�L��c �ݤ��b�]��U��9P�O���Z�Z�� ��[&T5��Y#}�%���xAu��K�s���&e-���Q�"��V���_�:����|*Zde������K+6���HAw���fD�g���Qs���P�!�_K�'���0��"�F����o
�;�}��lZAD��"��t�(oBP��M����Ԭ��w�E�@��X�AգcXv��f����v���o/+)v�If��	�Cq|r��z�����i�-��ܱ'�'܃�)�pȕtB��3l�ӷ�/��푮ܤ�2�VmT"M��<I���+�]��2�x
�a�Ed����+���@�ͺ��w#9m����ö��y�����Ż��u����Gqu���p&�
��<���
�w.o�QL��l��-DgJ�^>4�`NN��R=�Ǘ�3,P){�	{�)��p<R}�3,7����'�ܳ�A��etz`T!�2H�l�w��z@yf��`m+��\��<������Clm�����}}���/�4}t�6�����o9�7qN\1�����@43[�`8r��e�Շ���G[x�556	Q\o��kX�����<��g��w�`cۦ��Y�(a���A����<�6��|~���J�n=WA:���\�����d3Mbט��C��%}����D�ʙ]v��4-��4J�(S�F�.��L��NQ/LhZh�4���lљ!�M�أ.��Y���.���5��Ց�����y��y�=4�ZiB�9�Ok:��V�U�:4/w�0wS��[�v�-��359z�e���ռ��w^1t`'��2h&:�i�o�]��8�ӧ���ˠ��z�V��n���ɱ%�5ڋT[�ٌ�f�����Q,�����ב�(�Ul�g{����y��B�&eA�dmv�*��)�GLu|�#�����%�Y���{يe�i�_ �0md�cX��k���	ʉ����cћ�#��v:���>�m)V�,�b둦gk�{E�+c5x-W
�ނ�.�\�
�txma�-S��w�Iuu���xn��W�Oz��m��)W��=vw��{���;�9a�����suw�E����R��oQ�)aLX�t�`��Ρn͠�:ݜW�bp�ơwǻ.��B-�ڻv�����u�[E��-�+�5+�86N�d��±�|�>���\�ɚ����ͧ�<�qt�T��B&kژk��-�Y}���IM՚���p��[0b�,:��d����ְSF���+��snVe4�+��k9^�nQcm<ʳS�o'9�	Vw�(hs�zG�H^�j�X⸤�i�y���v���C	|��t�<�Ly/O�Rs��ƹ�ݔ�u�y��m:t�іA�Ǵ���f���)ɥ�����jh�E�@��S��-���IG��뗢��S|�7;���^P��ʂk��{[�r�U��t*f����-b�[��yHL���9���j���q�9�k��A ���97���|	��c��T�-A[r�n!Y�����ci���.4�cu�9��&(2�G�F^��hg+ǯ/[�y�[��8e�l��U�8�GaE���ف��s���1�wʷM��e���fegP-)���oj-��a��̬��Ѱ��[�Ѽ����γ�}�Y4�$:Y*Ѣw���`��[{��+�k(GC叜�">�p�̀4�^!�m�1�B'�oTJ����S�d�v�p�]��{,�(�	�W+�HHm��[]WtnqT��ð���4�euG��opB���nɓ^:������A\h��Lp��T�������,X9����]���$���3wRtkAX�Nׂ���"@�Z`�]4�1�7���P�/���9����u.=o/q;�
��iyU��k������	.��a�͋�]MMry�l�X=J����r�kUw�k9Rv��˷˻+#����:�Q�� )��R��ٷ������3��5{t�o��uo,ōD�j�	V��s{A���-����h��OlAJ*w�h�4�4Ώ�Ȼc���� 6>vEIa�:�/jbOlru�^s�
��u� ^�hafL�6�+Ďq���$WQ�[e��L���&rl�Q�c����xQ�A�,+l�Kݓ�\�ݎ�ᦡ+�PL�e����ceI��g$�.�X��c�]��>�]]c����X�u@�3�K������n�	H�w�8�x�;�5׆���!�Ú�4v�}V+-�7*=yO��ޓp���-���g�e[��w��k/���	�u�v��x�/em�y[NW}1�i���׃�zj|�XMiw����M;���j�SD=AhVwJ�o:XM�:�ټ}�h;˰=�g��w-�F^ J�_ 8�>Z	h�k�4��%�ӻ�^���
ve9};���� �3�+B!��̲*�T�I3v���C�Б�R�����s�Y�Z�'�Y��#�΢%����-�2h;��np����C�f@۽�'X�nR�5`ڰ�:�`T�0��w���*�)��ڭV����Pڦ@�z'<�8<��ڃ%���Vk�����[b�ǝ ��G�#sr	��h�� :��y) ��e�3o����M2�iIT)���k�[����L���/:$���c�ʰU) �pR+v�[�*��&�J���G{��{�B�5V]h��ʡ����fh֣�(Z� ��5>:��c��ʠ;�7���N�޾��1m�K(I��􍯶[��R�\����<�YL�j�'�+ӝi���d\�2��8κ��^R�W�!��G2+SKղ2�����@��<�ˣͫy��&+���T��M0�w�����o!�}Eh�Ag�k��u
�r�y܎�v�h��[�������F�%��8(;�s�����؅1����r��9�z�%({�\8�b���漰"�
Yi�꒒;�w`O��S��*Cr�f�:ڡ&`W+9�	~i6.��v�1�t�����:C�CM���]�HIsU�n���4{)�|�ާ��N����>ϳ�Φ��r�Q�P�/�Kq�;����͊fظ��,��V�������]��і)_N���a|6k͒�������E9�[W��i��Q�)��kO3e��F�� u��j����hXh��sS��][{ȾĂ,C�j��;���B��ب2�����gVںx���.��r��=�,�X�6j�X�ot�7R�<`��*(Uۡ:&i��s������5��[�2sy�
V��.eY���\��{,ι �aKb�`��*nmj�ʍ��;r�uyO���O��k�wxWe��_s�ԫ�{Gegū*�+�U���NYz7@o�k�����j�I�rb�nu���v��-ԇ.�D;t�o�ՁVRW+z�T��'�6,%`[E3zk���+7�Rb��큪P��>/U��U��DƘ�m�d=�נv�u齽ʶ��y���������teò�ީc� ށ���0mҬ�a��zuf�fF��w�N��J�7i� )_Nos����-�U�Xc5�#�ci΍@����{.�s/�4U�W�۽|2�b�Qw�fU��^.�eC�9sуAD6�� K{jU�rΣ�m����eY
e�vF=��?��JZ�� Y
����T�^�f+�;�[ޭџ8��c|��Egc[��2����0j����r���W##W� u{:�m'[��Ԋ�owP7Y�����7f���Jzn2�[�u�Zz1�a�_b��&�U4ͭ�H<�G����C�0g38>�u�{���o�y�ٌ�ATN����+Z�kU���2bF�jI�e6:�yS���g��} ;֗6��K%�K��7@:�"�(݇�[����ԅf/���5�OGI����8�+7x�\� 	�0�h�^^9��u�
��M�I�E#n��[I��ހpp���vPז�gP��V��R�`��QV���9+��7[2�k���f���XM�v���B�NH_VSֳ�v�d��.d�l]����lPp���U�u��ꈆxLZg[��U�:�n��f����Fγ۴�q=y|8`���]�41�;��������5��z���[��*j�z�f���щ�""n�<�g% r������#1����Eo��Ee�R���P���v��K"��M�]d�� T��6�Ǖ�ϖ���g��*�EW�mF^<m�'�LvN���O���5�pܑ0�KꝮt0q�u��%��ū�6-hfe�5c��six�]�ܼt��U�wukqfI�9A�N��� P���� �u�B�:��y���B��Hp��x;�Z4���Ҡ ���٢�]Ȓ�t-���hIdWd`��u_hC@�unݟ��F���s�+8�F��S]�T��ғ;{j�hrDea+٪�D����UGR�F��$�2��R�t���:�M鑰��X �.�Cn,����b�	ᨀq��U�9��g$�9�%(�����ư0��|j�䝐�*;����ƒ�A���Db��x�T�o-��'+��H���n�4���Z��i��}ui��k
s]L��e�9@B��k��T�+q�L���Y쎮r�J�����R*��<]:�2�mt�[޴����GPI�P�=�ؘGV'�wp98�9�c�WKu��T����ӫ�,�Zb17�]�Ya�8n���ذR6����W}�B�R��֎��]�Y�+��ԝ��8̑�{.�9����ă�h�w����ྮ	���7M�%)�(u���:���ɼ$�G����f��c�1C�t����k9Ry*ƺ��)��������
8ĚY��;8��)��b�f�[*-t^�5�x�wu�fwFC��JZ�(��ܤ[V���\BF��n'4ۼgrUuM��ɪ����;p���K�}-�XY����pc��I;���w��v���[E��#�mP�Oe9�x�S��ٜɌڊSݮ��3m��6�iJ���˦/�\�rv�`FX���z���U�P��
��_m1���fr�ɰ�]M��CS�E;m���.� �p�y��zq�]һ���-d�,�+��eYPt���*�:��8�2qc6b�A{o/�{�Җ6ZɎLJ�����J��j:y��ۗX]E��J�j#��9Ws4��n��]g���Bծ�,��S+�xgqO,��qJB>���0S�NٺDX3q��͏��x�N�f,	bcT���C��0T&�f^�Q1)�"����6݆'P�7(�9f��6΁��e>Yʻ1()�yl�/޴��٫5V\��g��dh�=c]�=��@p9|oe^V`��N�D]�;�LJ�B����K3��[�r��Cn�Z��1��Gm��s9Z��Օ7��A�4�C�f��o����K:ؐ�
�A�Q��:8Nq=����d��K�w9����MAv�����!ބt�u������(�aI��a�|*L�،�*��J�]aw4�ɻ�9��'J�x��T�����sU������ f�۸l��dYfr;��F˧��f���8�㱈��A�6�v=n!�3�1\���z
�]�v3��$��q����1��?u3�ֵ���R�"ѣ&Q��(�Z�r��՟6��/v�z:e��ӂ�(�u7м�&��j��6�߈�e�V���۾�6�V�ۦ�gd ����y$&��:�ꥤ�����)��sM�ޛ���:�ѱ�8�wVo"�%�O%e^潺��n-����f�o,A�xm��*+����+�ʜ�Ӥ���i�w(ĞՕC'r7�W�K��� ��<��ΘHU0\�/�Lln��o��ӻ�I���f[�vNof�0.ڵ�MN�A��c@�tm�!E��8ŷ���Ya��dL��6LN��Y>�0T#�8vt%i��NY���QfT]A,�^N��(g. r�u�@�[�r�Z�{kr�
��0�]��w�+���Z�;����څ=��3̓S ��c�-��@��U��(7y���kn�X��t�*;c�Y34��Y@#}��KW7�ԤKcyų��RܵN�e̥�xj�-oqؑ�����gL��/�p�lNӜ�M�̜�MŮ���H�z�\4�J7���;v�� �4�-��Ζ�\.�����Z��;x��C�\��I��~�.r�F�� xj�V�������N���+��V�EZ.s�N���kFI�h����z�2Z<�Rܱ8c�hB04@I�.]��]�Q�=�'�$�uՙ���iU��벯d+H��6h �7��:v���WPV�h�nU�uX��r�p�� =�+��{��s���R �*�t�����S��6�S�X6�"V�t͙ш�v�rww��V�K���s�tdZ� 7��\:��Ip��%��k2�X;
fJ���Y�p�`U-N)Νb�:�f�KH��咞��׹�Q�^'��bWO��(�dH�jyr��F��S������{mM��b�E�(�5k+V�3B\n�]�\����[��x��C ju��gY7h;��A��m�Ս�2��_rSc����n�n|9z�=�r��[i#��is��`��L���h''�lS�Xw��Nw�eT͏�w�"��moB��D��:K8�.Ծ�@��{ ���r7�{3(k�j;{�;��;�e��a�5R��fG���L���uQ�Z�?*�(�|:(���⨅qf ����˾�$۽ܚV�D��qs�i����|�s�x.�X]û��mq�����J��[A�Yzx(��A�nIа��N�@q%us^iP3���)eǯ#-����J�gٗuѽ%��ʮ;���*L�Ёi�ڳB�蒔����P��F���Al-�ʪ�\��	{	�]�ٳ���͹�����8U���]�1��q/;{���7�5�\v���b5	y;J�4mG+_I�J<������6ޢ�Ɇ�6Y��V|;x�l��T��iQ��V�q��фZ*fd����u	,_-���jcB�C���r�^_Nە�3{�θ�����e�WEAC�{R�Շ�@	PR7n0�U�2N�!�3s(Eӝ�ٜ�+2-��m�.2:��"�I:��DW��c&��z-!����������b�.�� �v���磆Qu�v"�.��4X��2�-�ň �]{����Y��Tf��R�m�u�.q���7l|D�6��T6�����s��԰.�a�EU�����Q�Qwu���ѵ�a-�}϶�g��(9v&�M�.t]�s#��K�/��ɇ�փVYfv���,���vk�-qsuI����&m��)��f[��.��F�$ ��$Y%�Z��Z�ڿ��������_}Ԟ��@��iW*ͩ{t¥�[5v��X2Գ�H5������{���R�o;A����|���.f�Z*A���3"yG:�um����/ hw��֪񾾬mde@��\]Y��m[ϯ�}=8Rdi-u�
l st(��?������oJ�l]����Q�,v�ｂ��M]�^2�n�NSS8�w���k3vL�y�s���i�^�,����ݴ{C�����n�={1�D�Y�b�7IÃ@��xr�jkb�3���[�:mt[t��k�0�Vov�X���R�mjIl8c���wv�v�z��� �G�s3M�OD�]��]���v�F�Zv�� Ќw�1-6���kNS���^���f	y`�d5՝W��iU����8+����I<��:�D#0�|�΢����`��u����+���+�}�XOf�U}�A�4��vgv<RQ=E�z�m�n-�B�h�۰���,�RKOE�5����.S+{+E�fL޼9un�2/i5�YK��Ϲ�k��HqnlF��5���wr���]�xۚ��g5�ɊsxΨ�,&eΰW:U��+�j�ǃ,T���ǭ�	�RǼ�ۣ��v���v4�	cv8�������NN�Л��abt�E�λ�*��]���Q�[3�5�PK��.�`�Эf�_�#��;\.�wmZ��˺�k�!��5u���s�3*�||�	$�D,�\"����Tf'��ŧRJ�<qw4Y¢�̙j�Ȫ��H��ݚXF�PȊw(��T����d纑et�Т���6x��T
%F����Qz!Ȩ�	�u+9vj{�r�ͫJ<̅�RL��ԺKfI{��8Rj.�K��"(("�i����OVW�"!Ty�NT�' �EՒ�A��*��;=��q�L�qH��[�E[��D�EN�z�,$���P����i�ݹj.�,�ӕR)�(�nx���B.���#�a��K�a\,�s�#�25[�
��t�HJR�TJ���Г��܊��I���#0�G���ZAE\���r��1M�e��J�M����b�t�*W����am��"�U"�Y���RI͞��ws�8hZ躂e)���4$®���L
,�䜋�H��ADPEE\�:rL�J(�tu0���s��z��Bл5�;�rL��������^���iv󋐹�g)��EJd�[��μ���z�`�-g0b�e�U�\x�uz�p}-�s��KY�Ɯ�W��f���0�W��x��nMʡh3�f+Ee^�t��N���,�B��v�g���}��_�n����@�wT���[#�O<E���gr���R#|����MU�.�Q��5�7�E��9���qY$�R�[�e��P(1���|����Y��f�Tb���^=&y�`����}��b�D�ֱ�[�6TY!q��Y��B����x�x���V7����\8C]<�Nu;�6�����p��KM�rЅ>뼌�R�:�R-�c"�)�S��NE��G��0N���i 8J dG+{�@�N�W���EC}����Q"�y�[ʊ��k�J0q��>Gl����Cb����`���xU�KH�?��pJ#�G%�����}�u���Z+�Y�Q܈���f��u���1��F�9�Ξ����5��V��7q#�%�/���'�Z�(������nL��Y�E4z���9\2:�nb�ۼYi�e#��cBMK��C��c�-@U���5�@a����� �A'>���I�e\LL�w$�QA'F�_F���:��L�[ۮ}�6��V��g�[�Xyx��T���Z
C�yMj
'zyw�ZK��j�F;:�]�t+l�y�4�-ӫc��s	O��RJ��V�]���������.���V���tu��}7�KG8G��V�չ��n���J�G��)n�0�u)t�q35Zs�P�V�E������9�X�p��ӌ��)��tl¸��1�8).	PL�1�:Xr	��aw,��"�[����P"�� 1�K�o[�G����V�c�d�	ƙ�@�Vf;�����)���u�_Ҫ'1Yиd,�ݝ����%o{a$M|�FG���E�#<�g�i�5���S嘬$�FV�E\�����{}�ܟuMz׆��z�{R�^���(���ty�#NQU�p�¯��G��^^Z�E�v��m�:��
�r�J#\�T
�v�ԃ��$�W%��ӊ .e帹�i�5��yk��&�LOl��M���mP��W��L�"��;�T���	x�q×��9GO��+�]-W����T�\ ����+��"yC'j��"���3X������X��RW��@�=�@��ߴ��{����s��/�{θi;|�*�4D�r�-DA����nг�7du�Щ�8����%���W���g�)\�i�\بu܊���7���=�"�`0�̍�gv���a�\\p�5��׃L*L4�U��nI1���[bm�X9�ŊV�u	{"����dj�c�ǆ�z\OqGXV�P0P�6��->л�����Z� oA6y�,C�V�.���\u�sq�#��K��30�3��N�H��G�=DAG�k��_���^�t�ﭑ�mZ�CGG�N�O���*�Zߊ�D�7��;*�,Ã����h���=BM��w[�v�-L�#u1VD2n�|V��Y�|$�ٳ}��%Էd��eqy�����Zm����O(���1��2�b�u��c7k듉&�k���*��m��|q��GW������r�ګ��Ü	{�6��V�[��0�F�spLGe}�bR�&�2�u|��}p���F�S�2�_FTT|�rtMwlΝG�ˏr��&��%�JL��>�����C��y!�?w���
/x�2����Q����K��9���*������9�+/(vz
5W]q�9�FpEq�z�Sķ��<��Z��F��)ˡ�c���|��:�p��V�-'Ԩ.v���y���P�f:�7�dB��R�T�e��*��'s7�#���5���'"JFH�{���4���ϴ��vi��nE3A���
�Tu3�k�M�L�^���K@߮�5)��{r�bn
�1*��m{�zG��S3�:nXvZnu���l�r\�=�fۥ+���u�u1����LV��fN�\����)ʓ7�yNV�[���&))����2�b�!]��3��Н���9����!�+��;z�>��ݭ��ܰ��ԋo��"0�iu��㕊bT6���{��$�K�U�םk�8���* ���)q˥_*���;�l!H����e�J���p�X//6۾�4C��(G���&�u4�&�|��]zl:�����({�_il��r��^��T��o	�u7Q���Q;ܞ46�~�o(�jI1��pʉ�C0Ȏ�� �-�8<A��3��$Xv�z�e�¶o����j��ٰK
��\��**��pQ��w�jK܍��Y��Хt�aH�i�m@⦙B�f�� c]R��b �����7�Ú�(�u�\�1՜�'�$�S��Η����f5:����7�,B�����:�����GH��S)ks��V����_O���θk���D`�S����θ�{~��|e-�L<���Ӄy��'J�9�3(ƾ�cC���y["�W��}>+@�Hp�V3�vCp�(bh
��Kپ2v�؜�Hek ����޽֬�$�#
��0�,�J�V,��ownPu�كA0O�g�8\	O��';�oLK��"XR��\.^��ŏM�Pmn�F�hzN�)�i'1;5���4Nry�ս���:��رʓq��˺�g����Sg"5O�w�(C<���(�
�u�)�<�s�@�w�U���lc���郓}%�-\�{%������¤Ώ�K(G(f��C6bR"c�z�)��8
����ʙ�,�ǰ�A�.�X�Y���)�g�y<T�s k�����R���D�Ԩ|�v�����q10���14t<6J�zex��0�ȍ�+,N�����{7o���b�'DC��L���%t��0�t+�������M>�
��f�
�J��3q�@�0PZy`Z�R i�;j���9l��X�V��gr���U1u,�1�ak�i���A�v]��盱SᰒWyx�ˢ�+xk�[��TW�/�CZ��fמ��!����_��g��9��T=QS��on���Q�@� u�����0(=��ƨ���N�첟.����"��f�'{b�[��w����Fs!�=�y�%��ZI��[/����P�!�V=�;����p�9E� (�@�Om�ˇ��ӕ����ެ��N47G��7�'7{|pS�bN�ErY�l�YeqS��˗�����a�4<�����9ra�on���}���pr��"�8����;��.�}���ш�M�K��Xc�;f@�p�+_Gx:����E���u���|�>�v�q�������Ϫ��c,�[f�J j�!��r�q�c�/���.M�i�v�L�Y�h��о^���YĆ�N��K�H�\�kh��-�Py�vG���Oy*����b�Kf��+��U{~l:�.'��gN�k�K%�_�=+�L��6�ʣ<�sӼ�0Qq/ଅ(=6�eq��Q��F4\s�e� ��KP����o��>��z���	�����.#&Xv����KG�����@k���`7]t���"����-��'�k�Cn��n�)�<9��u�u��B��o":�i·#�7�!�������^�z�g(Y��\�e����xm �,��1��,9�wP��\p�J�w�P!�f}f+n%z��P�؃:��C|@t��4��W��}��oko��L��b����%8��"-w�̮+���$Ol#�p���#L��>^�j�|��ۭ��3���ܺl���Kӽºˌ�+�O����E�Srt7��0��.9st�[$yL�Xۡ�{����d�qj�Q�0��[bU�uy��ʀxT�DW˛Gs�:�5��P�X�(�Y�x���$�t��@�}�8+�ѽ���}sVl��ͭlR���'T��-ӝ�Vʽrb[�G��T�uA�o{�}�lºG7\����� ��_9��"�
�=�� @V�m�=ta�ۘ�Nަ/:h\/p͍՗�7#d���=�{�hY��zǣ�g�|OY��hЇc�����g�+�YΥ��Ս��#�-ă�Ud�l�Sڡ&*!�� ��]��G�<;��O�8����OQ��<;�A��� ����c"�DT9�JS;K5],�i�w���ݸ�������u�~���Z����Nm FD	싚���=����w��u.�l����}�M��;��PK�ZV��Z�D=ۑ���3�>��\�mr��D�s<浕|���0�H����=:r��V�l��jՂ:<����;d��=�����y0q�z���c�5�-�Eq��a�W���<P���P����#�qy�ڹ}��_�z*�E���&{�Ȟ���l�~��4wa��'�^7�Y��oc����N�O9@�
|m6��q�*�ҷ$��4p�uxX�U���ԯyxfU�X�p����ڕ��ΐ�E�ba�亝&#����@?JU���y����	V������p�xi����e̪��mZ�,�2�|�9W{�[n״s�[G�{�v�u�4e ��o��V�&���v/�����r_7`�uҌ�8����ӈ�J�9ZCk�^3�*�v�]0i:�}3CP�n��Y�p'��'��.H��gp�]J�é[{�6v]"z�۷{��jʆ�$����ПB��;�
�������V���C�c<sz5�:�緤����>��
�SԬ:�6!;��>��mP-k*`A��v�υ���:�]*�{�D��:�|�+��3���á�V;�6�R��1�j&&9����f8�{U�ld��0Q�R՚�\b糞HyaS�����36�GKd��=��)gl{w|���L��H�#<���XM*���W��2�.�S!\�[!�eI��݌�$@��cc/���{����E;�X5����E����;�s�GS9P�6Ta��I<���m[x�uf�TI��Fƈy�O�g.��/�^d�B�{UjB��L����]�Y���i)��gj�m�ْ�gB�����e7�?	�2����1����?����IE�S��>���G�[k�p��q��Y��C3��s��Z�kg����mZB̃�Mȋ�o�����,��=P\�~����[�Tλ��������\��q��@b�{����ڒ�Q��n$aK�'�����r7�B�*��Ԏ]^�]���&t�wR�]���H�yO����"|�o`�5�d�E�	�F�1@T�c����7Z��}�;i�#�+{�9�Oo	�{Q�"���u�ÒWkl3�;#���/h�V���Y�uV�x:�@_O�]�U� _��>1�l&�_<&:�GSxBd^~���ڄ`�}fX��T����g����ixW�_g���|��P(ENr�����k�*J�:�'�&��ѷ���F���,���Ɩ�OY:���j��fSuF}۲'��F5�k�8\Ou!p�m�>r�TV���<�Ω3�uo[01��d��*�ۧ��"��Wt�������.��������a@WGr�C�&q�[���y��������aY�i'i��
�9X�%�w���xY��[	�o����#�܃�"����xv��	-xk���|�<tO{�Y�,���R9m��O*����}a�Bl��gH�i���PI�/~\�"�ĩ��@���P�mFom-v�Ҍj3���;2�E}�qۉ���j�k�f�́W
Y�òK���}�����y9u��tm�X�W��j�H����7>����8GZ ^g=��LZ�$��Uٟm�+=@�8���3�k�TD�vS�����tLl���d�aa���i��k��o2���Ӟ�;8����ry%^�����p������!��V�P)V� ���s��v������:����$T ��@T�����M�5뗳r�os��Ҵ��}=<�U�˶�s,F�V	J̓,F��Pc����&�.�x�^j�A�v�.6ti��҃��3�f1��EN�on��@yG�� l$v�kbלwZ�f�{��;�Rc�õs��Vt�d�@dw[�c������2�	�l8~G����;�Q^ǹ��� ��#^�[�nB²�s�������'+ �G���=��g�]��_�Ez�r��J��5eW�'�8![���B��^s�Lf\��mZ�YO;��!J���\"����n��NKG�?�D�j�~�)xm��yi�>�u��y�ѯM�X��o0�L0��|������òP(�F�S=+��^��2��I��_�fa��ƢqՎρ��7)���9�.��AkhvI2��H��kkr�)��򰦴
5d8��P��&Pv�|�)l��q��¦�|�M��.���5{ÎrX�oZ�-Ye���T�Q3q69��(BV�E�����\Oq��>��c�/�jV �Ɗ�-e�X5�m��Y�� +�C9�'mR�6:
&�;���31T%:�Ȣ]v�}�a��J �)�`�����!����.\�&�v`�к�K~�J	�^���̋Ŗ�^��׵�| U#�TY��b#t9��u�\;�v�:�sZ�9p
�ۚ�,5uu��)��#�΁w�9�w^�"9:sX�{*VpolK*��1��f��L��)]<�k�n�����O����&���<�$[
ծT\+�=�
�a۵�NC��,%^�UZ�}x�����Q��P��϶eK�%',��h��ȻP����<r�nj��:�Q�7��Ll�U�K���g0�x��
SԮ:�RJ �{ь˴)ӗ��7��r��k��&#�-���!:�}7��:B�����N�{׌����s$Vnv���T�{�I��M�ګ����f�+�5��ɐc뤨b�[�̎Xα@hH���Ә� {z���-�wX���s_Z��#��>�l�¥u�˧)���Ǐ׺Ճ��E;�S�	�;(��<�<�c�|�EU�znP��h��Z�ڙ����7��釄��s�p�o�[q�˫N�! �Յ[Zd]�m�Sjl��y��[=CE-�N��zLk+������C�;�y�:��F*�KP�V'}1��^�-��q(���)�(�v�+^\��iնnReϺ-կx1��uo�v��]C_M#��$sњ�^j��^S��W��lZM�e%v܈��n(��bS'�\����b�u����z�:�Q��Tsv�
Z��0N��xn�\F�*fuMU6)�-�wQg_1Q�֦[��sܻ�|䥃��ne��9������)������A�q�eu�+)��v��.'*ĳ�mi=x�����( f��G4��-
���_@���[�K՜��y\E�]C�+��e8����/%\&D�-��H�kB�P��Be�P�r�m47�b����{�#@*S�ٮ�]�Z(I�Xd��̻�oP�42��-�ҹu�d9��	�;���$̏b]/
�up���}��ⷛ�=���3���,���^j�`�#Ջ�@݂�}u��'[�Q�wxmU��B�ë
��y:��7ڶV�Ŏ�6���v��Q�l�{����+�x��%1ǽ9��;��]�j��v����EW٭�	�#C[Wz(�7[W�'y}v�ޭ�\��WL\�V��f�چ�,Ple����8;�
��D���l��K��X���1m�v5ŭ#2\���.�[Jԩ��R�
M�NqҬ"��jô�T�H��g�.	/������KDow��˾���/��kF��t�:[;[=��-�}�&:�l��l���!��uϒ�'R=��kYƬ�r�ܬ��4}���=�&�����--�V�5RT޳w�\*mkNk�]OU�5��.�ët�=����*�vP[Jn3�f�u��+��n4;�nV��f/
4>4 �^�9���m�wr�ʮ�"z�$����3����)hV"�$�D��-@��=������(�U]s�0����U�sWw�#�Cj�i!,%c����Q��P�*�urn�bJQ�H�(�v�bܽ�Y�J�r"#]�ˢJy�y)!F�J����X�t1W<�)���"�]]��a%�����9,�3nqS��4(��wd�S)%�)[er���U2�^z,ĺT�<�� �P�B*6�C��u��gP���JĻL��*k+��b����.\�)X����G=��DC��z%B�A;�P^�C��DG*�	D�%"%ZQ��d�nS�%PU��a�	:�j'44.��V�G*5*�!3"(3
�DJ�UM���,#S#0��s�Siʢ-bI9�,ITwvQ�*��"Ȥ�H�&�C�*QT���I��UJ��a\(������=����?���:So�Q�N��0*La��SΛ�3���u��+�&�:��=w ���+-��	.��mwP���[�ו��[�ެJ���1@h�,D�WQ�}b>� <���}~��y�9�@Y��=c˾8�Y>;����?�ѹP��O�z������>}��w�Ј�D\7��!����q%���sײʋ���z�z4Dp��"$z6{)��;۵������xv����ό~y��]�����r�|(U�������|qχ�]}C�<���iɤ'}C�i��+�aTߝ>?x���C�>�k랏e��͛��#E����G�|yAw��nv���{O)�������߻�o�'NҾ}~��)�	ǒ���9����N�[�S���>{��ɾ�~����%p.;�����Ϸo߿E.���:�U楉Ĉ�E	�����xw���;�����aW��97�'�|��ϸ��y|8������O.ӧ}}�~�4����ܮ�������x�>�4.U�z��D�˜��s}��(h<r�y@J�F�H��#�e?���W������ۏ�s��������QɅ�\}���?�x};�a~����?��|{o������׀��q��?���~w!���$B���P5��{<�%��# >�#�~�P�_�|OG�yW{M }O>�p|M?��ۓΠ�����R>v<&���v��x����?&������|�~�{o	!��T�w�߼�p)����l�����b�V@[�3�#�|^pO�{��BO>��r�����}w!���pyL*��y�xC�{C���{���[rq����	9�����e7�'�������~�o�H�" �k�@�z�/yeO��??aC�������yv�xB����*�]����:���q�����ɿ��<q�0��oo>�~��®��A�<&�����~���!�Ј�6"!�#���S^)xEz./MW��׵:S�c}">" ��|�+�`���n����0�|v�#��7 {I<���ϝ�w����Nv�y]��G&���v����=�}M>�׻��arh����P�"v����F���]>��tp͵�~��|��{��A��C�����=;�Nv�^�N��r!��g���0�I���׀�����C���bW&���~���&���v��C�k�=������,m�>�����O�K�w��%�T��Z����3���W����p�=�	��~0p�aSb��<�ྸ�f-L�Cw��hi�/����Kʾ{kx0F8���IR��p+�!cS�T�η��e���v�u�#F�
v���P3����]N�"��v�iE�BJ�۵�Q��D���1Tb#�τ�����$��r����&޼��������ׄ>!�9>&�N~޾������r�{��S���r��s��/����m�S����; ������z>�#�,C���F� �c�m���o_`��\����!���Í�q���m���c�]�;۽����c����51���>q�G����_��<?߾���L/����O	�!!�Q�˷��|O	��>��;�[����HI����xC�k�[��)����z�����Sr���㝿3��N���D�cV��5���#I3��u��r~�{���?��1���G���'���<�|}��O	�>]ɼ�&7��<����@Y<'����|q��{=��|w�;�o���o)������#�F� ������j��̎��^:�o<+�&�~7��e<!�4�O���q�4���k���דS~Bw���x�c���;�'N>�_z9�����Wϋ&:���9���w�<���G��ň7���VzK���=K7��#��>��1DX����ԫ����v�?[�n$|~���97�$���}v�����v<��&����������4��>�>�V~��>���#{�^��g�׶�U��_<���<�[zw8M���ӹ��{�����y>���}OI��P����&��pz;�x@�I7�$�~��xgoi�}}�{�H�����>7�}|&��A�?|�"������Y�c�^�q�O��0�S�~������<~q�o��n���P����El����q�>|��z~8'~M�����v��<&UUG�,��>��Q��D@|�G���� �Ug�t�Su��ۿ�W��wߗ��/���zOs�8���x��~w�9>;׋�S�������������N���������=��	��!�?<p��I��?>��oo�)��X����
��Wɸ@/V���󟠻봒����S�����ˏ�'���o~C�s���x�'���|w�~x?��L)�z����Os�>�s�Ă�w�>��(�M��ł>��}�G��T��h��顶�Xp�e�{5ɷ[�uη�
�[����NN�q$�_��q7�W+��qd���{ֹ�y����u��Z����b��V�-w�n���!G�V#PYg��n��OX�E=Lm�xK��nYҺ�Ɏ�-�x�n��N�3v���9HG=�zq��@�~޽��\N'��k�q!�4��?'?7z�"��C��Hx�o��q���P�������!������xL.��v?�)�|���|��>��H�Q�}���wk�u׻6�����Ǥ9?>q����Ԝ{?G�xw��7&��q;~t��My��ߓzC�a#��bOzM&��
r.�ޜy<G�ߐ�㷷��
o�O�{��4}DC;V6q��k׋3�tWo�������xp~�s��_c||;�{���D?�_8��w���M���<>P�O�s�����߼��w�9<��׀�C�aT<��{�)�{C�=�x��*#�`�G��|F���VO��G������{�y{��xBC�?�<y���<�׋Ӄ�~�����C�����H?>������P<���{O��?�O>ϰ����~���|OI��P=���"D} �{�"��|�V�Jw���4�	�w��m��H.��},(M�<��y}�ro�O�pxq�_�����<8�O��>���H~C�����v�t�?���P��������#�O�V@��y/w��L_U,��>�B��8}DBB��B$G�{^��i��~��=,r�zI7������w�����'y�xw��nq���ߝ+�����/���Ʌ��Z����������s���3�+#�������u_<A>�a���� "4�~�>w�p)��?�z���8$>|���������۝;˵�7��x��p"q�����Ȧ���;�h�� ��"&�n1�(�eWY�7�˷�ݼ���G�� {A�{C�zǿ��}q��{��(�C�4�>������7�$=����I�\
o�G��˧k���ׄ>&�8��>טw�i$�c뼪aT�}������_�w�ۋy�}b>B0D����z�m�!������ߝ�<�~O�~w�>��9���xM�����{>��c�8�]����6��$�ۿ�<'?�7������W���c�N'�,w;��3fow�s�S�j��}�"�|DBO�#�y~;H�M���7��\r���ro�_ �}�����!��~���o��90�>~��_)������U��N?���yL/�oG�����Î@��P�/�q!�u�I�&�<�f��|$�b㥭�۾��w8���������'{^�ť"e������^��/ü�xc�/�$�u���.
ѻ�ףx�i]���%�`��8Z,�v',���m�,���}��U/JY����Z�w��x�3�4F�NP���WzOǈ<~��@�~��n����n���v������o�I�ǟ���������_|r�v���pI�?&��}�=w�ǇN׸��s�C׾~E,��Mb��=�� �׿~��0�S�y��w��)Ʌ�]�?�G���!Ʌ�y��~C��G[s��9]�$�!���߽����7�'���o�����֭���*��I����#�|d�7�����?�N�|}{����aw;I���<�r�C����|Nq���ż3�C���}v?:O	�������yC�8�7�H{Oh�&�D�]�u�w�-�>�g�`��DD!���|o�zOo�nM����N'�ݼ��&���������HI�=}���<��]!符�����y�xW c�d��_�d�;��U���uUFJ�+�wu����4T7_B�sf�@4s�U��D��ԲV��`�n۱�P�Պ�N��2���vl��cLΆ+��Ѫ`3�E��+�j��p�:ʵ�};<�
˭�S��Eh�}Bc�E$\���5��@O���ƫn!�6s�]��z�4������o��Y����Bm\lR�L�6bմH�
�2g�4��'�� n�٬������=j���(,ڻ����oF-�nK��2/&��; 1T.�}�ˬ�ke���k��1��Q/LZ;�ֈ殸hϡ����Z80���h��ۿ/���������>�(c�\|�n��*Y|�*���8w>K�33����-�NC��.�1��ޥx:�����v�:0�;Y��y�iA:�Z�_v�Oq�BB��6T�[Q`�"hY�/@�E7-�����).����j��9^�<z��s��*��Z��Qrz�e���:�0�����9CE��ǱuB�����n��<�nȮ�b��46qsG�D����#�
CW�'p��w'�uu!gJ�S՜�q��`>+9�*�R�k}%�<��7���~J ����v�
��G��v:Z82�R��̽5
�����9�K�Ў\����w1��Un��g�P�$<��8��̭��B&��B�j��q=�o�t%�Y��M[�\_* f�����mW���mO��]�����ڰ������]P�㄁k��ϥb�t�;u✝�/���.1�#Dhd7L�,�l�b�B�1��[.��)�!Em�SY����x�����9����f������T[� #>���y�ԕT��e/oK7�n-~p����B��=��v�����>�,��\��VPp����73����cY�O>g��
Y�_I����,�3AC(�Y�Wʙ���g��D���]M���Or�F}]����]��\%��5�n�eU����1P�D��(;�VK̕0ڑ&%��������<b;�;�cTMn#t��V����n�8U�i�w�l���]�B��t>��'231;��:k������i4�`��t�͕�w^�����uw}t���2!�[XU��9z�p��Vd��޵�Nu�^0�q;�Xa�d�R˃�]I78��]R�?��e	Cf�sB�`�O�E��Z�ub���T]��\��Q�t�� ���a��<�8���3�ݗݚ�]��!���=nbF
����=5�k�4�7�+��w��pK��;����\�;Z� �v@u���s��O*�Gtf}��b����-k5�!�7��x�>�z��T����S��ׄ����~�x�ZF���IӃ~��
�軛V�|����s�7�����/�@�����{\tX�5�x��}�x���VS��n��۽B�R����.��%|e��(�QBz3i���-Ϝ�\xp���-6�Z}��Z���H]���G��(*xu6�Mf��ʸt��}>8�O=,`К����Jk�Z���=�C'94p�U���>�|MV���E���Ûϥ�t՚����S��,�-s}SY�l&�÷Lv�:�7�dB�Z��%�JL���B�ua]�7��]M��:�͞��{�I��G3P/�~�R��7 G#c��n�H�ꠅq�@HBp|z�]�8��ĒZD�.c>
D]��:[-lc<z��i����~�W����,_��y�q��i^K(�ǔ�����/G��3��c�����6�n�B�ͫW2}��t�:{�9��9]L֌u�9���]��݌��7��VN�i�-�ƪ��ڤ��>=]<T�b4u�ܖ�,J����<�8!�g0���1J�I WB��B�8Q�̓w��)��T�����zk����b�B�=θ<��+s�Nf���p̠y�es����I�b�8̭%�rR9c������B��]�a|0Q�����6���^p�������X�?�w��_ԗ��j�r�a��,E��^N�g�>Q;�Q?n�P���;�V[5b�8&�j�}�Ug	� KBO
��e7�7��=��ʎUダԹ�uː���$n��a�Y
 �Bn�¹6y��Kg$�6^E�U@�V�U�|�j\��r	�Ui����f�΀#ճ�9�kR`wB�>9Y��j��"MXN�@���:�H�跫��2�"ys�r���x(n��g��\�����Vq�v!N�\�E:��;Uκ�wIgZ�cI�r@znK�a�˚��0�}�@ĺ�=��l@�1��%��ٍ*TgORZ�N�R9�u�[[e��i'/� >Ca3)SX=qC�,.P�B���~.��D�b��wb�����CQ \50�T��U=��L۸�o�"ɫ��K�\H���
�wY)�/J�%���`��jsη|���8�X}�)c�nf�Z���J��b�MnuK���\��	�u�Y��bL�ڽ���;��@��W�=�����^g{P�Ρϝ�o�u��O��)Mě	M���g]B����H�Ѽ0�����U�C%D�q�W�Xxo�s��c�cD���������`>��n$8 ��Q�?
�gq�ǉ���f���Oj�]6sO�n��(ECUo(gݓH��L�^�|)�v:����y[W@�UH���1c����8U�v����Kf���	����őY��W+�n;�Jу�b��2�mka��;f�*������S�ok��wm�k��+���+q�`���NQ1�Ĵ{>��["�� 	Xz�y'�]x�z]��\q��0,:(��U��}����a`������tC�x�xv��H�炥O���zۿ+�-D���ԧg���g��Q�}�¸Z}V��Ѕ ;[� կB(3^n���:����z������z�-���Je��c�Q�<�W��$�A%$X܄�y�rq��a�ݙ~�뭞qη���������E|S���ɮ�A�y����|�EN����U�hB=Ŵ>��t�����1K��ҭ�%i�L�4Z �=��m��7A��^�3��[j0��w@^m�;�v�:�GS!�����Iz�]�靵��_Eְ�,�V,3z��	�fST�J.�GZռ2$>��R=����5l%cI�#M��'�}}SY+����A+�[�H�eҳg�Y�/�㊉��(
�z�C�*"��:�y��#frs�����k'+^���)W��`���Y�\.��XV]���>���q�pDŲ��ŝR��IX���z#�_��6���@���-ߍ��&E��6M��̻�3�-�kUb�Bœz���u�%������?)�񼤬YĆ�e_I���z�M�H��zgY��<ë��R=<}��^X>�[ɛ=�h{&P�%'J�����g!X���[��[�8�ۅFL����v':�v�a�΋)�����1���ppi��V�N�f�k���rq�ːo��q�/i�R����w������=��|M�	�U,�7^f�ro���\+_��3�8��RC&�z�2�;���:4[M_�lr��[��q�j�T"j�3̑���3ao)���Q,Q`[��4����}넞�{������4o/�uop_'ԁ�@�P)�ܳP�l�c�Eq�����&���e��y���E̽���w�yu+�s�-Mgb�F�$�I�R=�XP�_3�0�)�'rP�2K�a����Y�f��8��c͕��N�-Ş��9^�y�|�-�p=�Q���I7F��_Z��4eJ�R�v�jI��jN�����7m�kn�7�t���'��YL6x�Zd7z ��wDW�IRF̾������5À���w�GO8��8���
Gt�ļ)1?'��-N>F��g��@OGDii:��f����^.Ɋ�F�q�C�1�~��8��+t��S��_3��R�@uˀZ�a�m��v��V/�7�IX\I�SU]��ՎuQxb.�p�B����y�|%3%LwQ]q�jƓN:�餮�q*k���l�_�,�)ӑc�΢�0�&��:�]B Byd�|�{ծ�q�i.#�v��vUyR*�h?K��5Y�����5���°��Eq�e��t��nl���Śd
��#���Ab�U�r&�:�hhK�Z�E�Z�fK���%�e�G��a��O|MƘ�F�K������|��W��cF��Q��{��}1��]>�$�Kv���F ��~�5O��V�7�Rd�+NM|�+�m(��O4T����y�GO�Պ��J(%�.*����q%�J'�(+�����T��@����*��ܘ} �䔝ݝojdUykh=NC����SHp;��^�{}���O�u=i��wn�ͤ�)�ZV�e^��-���%�����Б#���k�׷n�W)gW7L8WK��u�syw��e*��F��a��YOM��c�Ӛu�LWQU�ٟ2�d<f �NTȕ����[BJ�1���^�ۍ�Qi̬�L��EI�cC�x#�.b��N�8�F�n�|*�'�i-��@����J냔U�!(P��q٭�r�W
��^�
��})�����"�3�(�,�&q������oWRQ)���r��{�!h�~js���z.�i�Ud��'�%��%���v=�0�l�iAǠ�(���h���c2��� =s3M��Y����/�V� ��&�ͭ��!)��/x*��cK^nZ�Xʥ��+A�l<P�m%�K��%4<����#�#��
��+dV�:��\H�"�����aT��yJ�f�K"kui;2���/���ٙ]3�lNmM#�T�Q�jv�p�+��MK�gEv�9f�X�ݟ=)�.d�j�%��m�2�����k�.e�ѩ���ڔ�a�4�BW��Y�6��ա�c~��)2�{޷Ϣ�;�c�ԉ�T�iTR�A=Tn������B��_V%�ʔU��yU4�l�/7r[������(���n��{�:cU�����+�L�s��4��a�-k+ڎ��J�[����p�t�GE�Т�u|�ۭ9��������;�-R��l�@@(E��af��:O(ڎ�X�hּZv�`!Y�Db�ff,��ӯ���� +%ؐ	JV$hq�\^q�0�E6�۾���ס��+FjNJ���S�v���
'����t���+ S�7j���SW�,-���'�(ɯ,$xveI]��J��6��²b�TY1f�J�Pu��莒�ө���f�R�9A.w}������x�������Ze]��[����Ҥ�M%��v�l�b��Pt��U�ϴ�j�>	G�ݚ!��y�Yx�UmK �!��-�t=~>�28b-O]����\�ķ·�,LC��,̭���=�
bm\'��'V�#��Ni�Q꺱�z��\qi���_S�,�rP\8�ǽ�8�Rp��S;�*�g7�Ad�zn��������)fӇ_rfn��`�j�й�ãw+��\cm��sf�pj�+��z�p�ԑǳ,���	�o�@\N
T3�B�ڏ)mE+VF.ʂ`|�yػםF�����*��"�ne�SJ�o�邱����[!�O�-M��u��bޮ9�����.�:���9��䈼dc�X+uu��N�J�N�s����2�K�� [Ǫ�����ݛBu���\k5�{4�c ��ŝ�ʹ�E�a��%��n��'6��b��� ��j,�pry����; .�w�i ����=Y�7)�w/�H�!�I%(�r��/7����\���X��[�Z's'J��]J�.�˔��9��Q���PР��H���Pi��6MV�fj+4��s-H�L�$�R������9��W*RI�9XAr�r<�9l�	Yh���vK�heE.������T��=O&�DTTUȬ�s���E��:�Z��lYfYR��DGss�V�X�f'#4���I�\�	5,S�Gu=B����%��yy��іG�eBG��3��;�y�w(�N���ݓ�s��u����RԵ\�w9&���U��'5���D�r�O�=��<���(/3ΞI�5�6�e繂*VՉ�N�5u��7$�hD�z�3ιYh��\,SwwMJ���']ĊPӮK�U#32����b�e�jn{�J�RE�AA�j�����	G3[��΂^�`B7��3ku�좈�X���)���{)u������v���t��T"�����w!�WTN��їD�	�w�}�DDym󣯔���������!���R�Sө�7�&��na#yS��.(-���q��X�/;�
�ûn�Y�W_Y�i.����t�y���JS���Vgk	���ko�Wp��N�|C�շ0��q,n�0w���17TW���������.}����o�ūӹ����Ρ�P/�~�T�#���͜��p��By�.42�p���x8=^|�&絽_Y�~�j�GV�B�6̖�����)�+d3#�Cr0�ǖC�V�=Yq�N�j�ă��d��1�����S`��l��p�{臥yk�D��$��}��;x=̤��":3b�FFT�8fz$���EO�@�䄽��n;�i���+k�ҫ�1Iű��C��X_�]Ӓb�u��-1\�2�驅�[�����]}g�yE\��w�����Z��ɴ��8��cX�2!���9wci	 ��,C|�9eI|��$:��ڸ]4���SW-��A�vm�:#D�eBf�̶1:���X�m�������O���?�-�ٿ�1Z.�N��X�;qfPlj���BSJ:��C"��:�6���o���˳k�䩜a��m����,|�n�q�9/-Ι;-�35G)P��,�KA#'s��b��'b��ž���*\�t7�r�6D��[w���#-�&�uu��ѷ���q�18L�ʬ�7�|���(����?gm}P��:u�����鍸թb+�&$8ʜ�q�_;((n���)W��ٝ*�ϓ�`�+Ú0^a�2F�C�'r�븝o�@A[S����U�\"����*�u���և��[L����5˝��[��G.�{n�v|��>�E���n$ň��f��{��\
���Q׭_��4x��n���xa^�--�C]KЪ���
�غ�)��a)�����M������|�V�^�uT$o��|~�R���瑎ϝ�/�P���Gd9UA�zz*n�|5��l�{�%�̳���D��.�Ď��}P�9H�����P東�9E6��Իa���S�j%re�HEJ(�х�:�OI'���X�3�~�5�ԯZ�Mg^�J²*;"u.426�:E%���o-�i�b�%��Y���)�g��@�&֪�o{sq��z\j�5�U��E�Ո!�1�+Z���u��
8k�&=Y�_�hgʗ�����z�����n��A$7J��N�OH��Qy�}|@��U4k�=��K��gٱ,m�>�d��>v8r���$�U�պz��+U��5-��C���yJ�e��w��4��*_n�����sVP�/��\�U���Q������;�>�n6�1$%��4��{(��_[YX,�dq\t���&&�T��j��vLʪ��N_.ؑX���i�b��Crg,��y`W�j�ȁpa�ڃ?!�>��}0�T����رH.Td�Ӌ��@&ԛ[{�[���v�;���T k�q;�cz�fz�G9`ܾ}O���� �)-����fj2P�3Q}ԙ��/�"���8ZʨO�"y���/�ݵB��p0@
��,>��U�
X��58�u��2���=���t��\�>@#�ז�{�f�g�a�i��[�iB�	�Q�@�W��  �Е����ն�d� wn�GN���,M�OC�7H��r_1u��匘�%�_&z�wR";r����]"�:d�1l�Z!�N�	����fQGs�vn"�.�}�.Et�w}�/2�%��g�#6l(�"b��x���Y����e�(��6�o��{x�]��wu�s��=�v�{et�������W��GY�{˼t_��ƅ���������Ʀz�˴�;aK@ɒ�	ɣ(r8җ=�4���;YyG��L��T�6WG�u�c�[�֝i"� ̫�S���k"=QN��=��$�&� �,�A6��f2�wGYز^�Xq��[+�sy�.�Ν"��V��o���}�|&������8���q<@�ɔ��W/�q�T��u�_@/��
�8:���z{RJy�w�N3���/���p���̎ e�hy�\4��;�Yu��L+u����ã�CzAv����ؗ�C ^�o!�6�DX���֢���t��1��ۻ2������%YV��
!S��7(B�B���62 �o�U�d��ܼ)��z�{�=��dK\ՖN����	wTV��l��^V���w�
u=��"�P㢄qZ�M�ʹ�S�-����+>Qq���v�'i�3��jጂ�ٙ7�����7"U��8�K�I��[ι�UI;���鈨��z|���[��
f�-����z*r�bӴ�ު�f¾�֌0hd�K5q;gԍhƛ��V��8�1��N���jv�=kJ��?�bҏ���j�#�H�+����<�=�Q�e$wU��s��0��ú�A��_1(�����%���f�� {s��e��:�ĉ`�v��N�Ջ :Y��[rPֲU\ل"ҰN�
7{P�Y��ŝ,)��I��U�1Ju��w�;MInyՀ����Ȯ���L��Ma����Z.�G�tw�pE��]�.����v�}t&'g.��'k��
It��n���]j�C$�������C��Xۧ�^)�����Q�N���wv�����`�K Lru"�A��Nq����Y8c�b�����m8�v�rw�s�X�#\e;�y)\舶V��M���7p���)���}!W�N.g1ջNwQ�!��V��Ѯ�v}*��*��q�q}����ܷ��'��KG;�,Ҷ�ka��BK�r�6�`�����;u\��Ã�%|eZ^��K]1���?O1;�z�<��T�w���;�+Lً>�\��g|D�ؐ&Y2�Q3�2� g�G�_)p��7�6�#��~:Ք����^=<�ALbn��#�>��	Jx����Y�����KIt�[�9�:����C�]Bౙ������c�IEtR �9�/�����=���5ʔ��À�;�nmBF�_t�P��q���n1�Z/)Vn�L�F���YU9�X�]�d�\O�B�[�W�!�n�i3qڍG\A�٨.cp����?	V�D�[�)�vX����w�z�h��V��zJ|���>[f��n�hy�[����~�YT[;u�61@Q�n+���9}׋JR��s��;�� ��b^�r� Y�\�� ��79p6�@W��8Y��Bk*͢r@r��P�Gв��Ve@�:ޮ �Lg�wv#)��"scTwm�������_j;�Sq2'D�旴��Gyt8\
�F��>�����ů%��Z8ML�jbwP_�p��{��Q�����}��w��2�u�C���=y���'=*mxfY����Q\BR�LX�1:	/N(��]y9��]NjA�Z�y�6z5q���T�W�LXRa
mP�⪆3�L��t�2YPw����vy�ֻ[Kf���:i�c�;��+�N��8�P����в������Zq�h��:����/�
VL�~t�kf��(>��1��'5��w���m��Z��Y�1󼤯^�%C��d�VѢڷ�r�1Z�/f�3��Ҁ���N�U���CΚ�Z����뛕������3�'��8i׹�g��U�\"���*үW�����vЧՃY �%��9-HKN��*|a������kl�3H��b�mD�&c���1p��$�Q�:�􉞞��u��{�6#��=/T�p�-sU�Ik'G.�+����ߩ_��~�ʶQ�<">s��Z�^U�fӻ��9����:��u�X瑎�wLh�U}hd)�"6��Е��ۖi�
��a�b+=���i��'u֤3iBcd����)�#F���"��ʬ���N���5����q�V�{�F����Wr�'��z8�q���46�-A���ϋ�n�+d�΢*o
K����S�m=���ְ�47(�^�U�?D}��M��lU��\�9>��LEmDMg�Ď�_r}p�.[,���B&�[�3w��i�P��)J<mƙ���;&Hy*��_\�ы�R�&�'i�p�30$��ԗ9���|�}��	�t���lĤo����'�A���=rr��	��P۬IŸ]x�"d�k���;�<5�Ѐ��y ���נ@nEKHI�ԯ�=Q��X�=I�n.���p��*�'X��A�X���L������k0��-�S�K{�b��޺/�pݼ5"�	b�Oj�6 ]�P�Ԉa��t�{��jk�OFk�_`��B�;'t�.��S9"�;�-��.f�8
�'J��k���ͭ�ġ.D+&��B4P��U�|�"����CL�}�(5�3>�f10�EJ;#���h�-��|/P�k�p�B �]R=����ҍ]�uQXb���)�/$>U�ᬎ����ȼ|�S<���>��n;�5>�nH֋t����,+/��xV���_����{Xxn ��ʏkk�o1b�66��<^�\�
�0s��r�7�1��@t������8��e9�扲���n�d����@{���ݑ'ɼ��V6�b�2��OSUF�n�� R�<�i1��j@����I�z�^1��BHgd��G�f���e)o��S�d�����u�ݙ���������}�\�^������F�[�@gF���B�{��[Z+�䗇VU}bb�[�u�:� ���np��켸�� K�h!��L�"���N�E}]pя�WԱ^��Y��x<Ӌ���zJ;����ȷꢉ�H��*�}������=1؝1��4=�<v�L���׽]̭�@��&�L�����2�ۆ
7�F�<�g��1�v`��ò��seo��7d3����O"�@o�;�U��\d��|����z�W�<�lN=ٞs��c�g�5���g�트VJ���ʣ��M��IW&�YѴ�f���Qo��{�V��{�Þ�\8:�Y`a��\1�ӌ��$@�
�ꮣ��K������v)�5�]��֭�7�*�U.8H�N��7ԁ�@�_JdW��7�f*B�c{OpݜB�^b�m��j���RÐO#��'�%b�qW�6�+AX� "i�2�uF&�<E{ݺ��7��I�pAq�	�/F�Z�)��Vv��+ꏓ�4��ʲ��5N'9�6;l��vM�u�1�a��v� �rM�ST��v-uce�����Oatx�!����M��ʰ�O��$���ȃ(�!G]�J���v���$������g7�,�t5Y���]Y��]/�W�}UU�l^1�~�e]���'��U�T�$WB=>Cmz����+����k�ٽ<�V����ᔓV֎zq�Me�Qy�G�E�N@���IL�V#�t�B�ʌ
�'~`"{e�e��غ��8�v_��ߐ��[S��4���:�:�PYfR;�"���E�aa���P�Fq�MrC(x��T�ũ�Ds�d�9�7�_\�7s/��N�,)�Bǽ�Zv6�x�)��9�QYJ��?�=wj�ډ�.'!������!���������#��������v/K'�z�{�oLF3K��ۍ<퓐�[=��B~MgdSX)��v��nv�N�J�8SY�uJՂ#�΢vzZY�Y�q�8���Μ�{Ǵ���ڢ�~�����i����v�:exՊ�2�P�� �(a
��F���|VOTPN`,��-6��獍�ǷuG竅4u�zTOuF\6�'��\6�Vi���� ]O*��z�kin���|�ޚǫgb���|�=,`�q+�[r�ګ�
�@�F5��I���@车��iĸ'���Qb��.2�\��A[ٔ'_h�S���k|�����-jCB��<����z(�2�:vϷk��7
�V0�w����k]?���=[�ս�~�����r�QK�--C�9�Z�����wo.y���t�KP��]\�����ꯪ����y�b��q83�g������h9���9��=��:�����@�Z�o�L}gqF�|̓��4r�z�|*�cfz5Q�	�_t�P��q�n@�Gn��%s0�w$�?'ͮ�����TZ�A	�j��9�p�KV�
�����s#��|�'U;�ST�ӽX�V{��=�p�S�� N�Z1�U�u��*�(�m���}4{o\��a����o���Pv%��UZ��]NM��rJG�&��LR��� r7�l��rRZ���١���n񝂤=��hc���x-���:�o0��j�	=��q&��Z���/��O���r�LXRa
mP���|M��O@u�5/Y�8{�����]j-ڇFm>7��k*)]�	�E���h����au4z����v��K��H^���q&��X=q���get����p�9Mk(�nO<*�7����-b��~q۔p�ܤ�* 1��R���֘�qx;2��^�s�R��~�m�Ƨ��g;Kay�E�j�f�o0����B�Z�����uȝ6[�R���t3BNθ𯋗v�D�fV5�ي�vΠ`ԑ�X��/�\x�Μa�v�}��ǈ�Ѥ���m9po��R�Po��p��<�GM][��m
l��Gq��tc�qw<n�q��W��J�vW�p�Y{K=���w�Rh�Ƀ&(�����7I<���+�׭�j�{{rX�MIt�����:}sV�����6{��N˱���I��+" o%����:�E">ܣY�ۥ��|B�&R�e)��d�ƴ�ُ��k����E������lf�� Ь�ˬ�_C��!
�x�ͳ�F�1�R5�NI�}�q�6_(������I��72���.6�,��]x73�
�i�ד��i5��` �l+���K{���M�x��5����6�l�.������d����a�"�e����9qJ���J�5h�t�V�1������e#3q�}&�mVj4a�a���q�a�_nc��n�[���ڡ���79z,�z�9/]�.�M;mI��~ �7Z6 ��W�e,(�{��j��u>oi�z�}p��Q[1���6�S<��r6^	$.ʆ�o�\<:��!�����OFN)��2S)��3�S������c��՝o5d�+�?G ��,t�B$+��r�rp%��r��9�n�mD��Î��q�����z��I����q��m��V��LMAMوm�a3����/0���L��Zii���q�4��������t�~۪UKA�Ƙ��V�� �&tx������O*{O qp�Nse8�7�POdD�K�:Ԛ�ц�$m�h�1��9��/hq�PZ/xo����`����ف��h���Pw���ܦ��ptw����:ɢ%��[�N�rf'I
��"�jY]Vz�ak�yt�p�F��=��<W б��>���������l`��Z*魼'T?��BՊ��0Z}h=M��:�e�tn�fۗ�(�J�]o�'D��5�c�4]e�wh�tzp�Ek�s����^+!�ݎ.ohN��ֳ��+� ���w�fS�)���l��if� ���ZW�*+�[��}ծ���Z��j�2�^����7��b���Eci<���O8o4���H�����(*�#�+#�_��.���F��l���u:	Tx����c4XI���T�׆�2n��Ȭ�gZ��Q�C�*'2R����ʸ�y��]񩌃���Xx�xv�Ɵ �P�]�g\}i����_W;�X�;�H.<����x���1�fY�g���nn�@l]֍�m湛�ݝO� i�4���1 ��HZ�[:2Tl��` @?A0�e�J$iQ%�H��4�����:s:T.�^�wJ�rr�	\��z�9;tNDҢtt��twE��E]Ж���43�܇��*�^�:z�:��4��u���k���G���&UU�g몚����<�Of�]Z��u�n�K�$(�՚�"�����������TQ���8)�z^z!fKL�B�t������,����/q���m�=.���N:f+�.����*.V��U#m�����e�*JF�$��sH��\DE���w79S�g,�"Vg9Q��Ҍ�� �W=�a�ՙ��3 ,*Ѫ���D.�Ms�����4�SH�R�LJ�waI���z燜](BU*�e*�:�
ͣ=�r!ʋ�e��d�T�ʈ�2�*�Ri%t3T��$3:'"5��hU&�������j˚���2P�-.�.f�"�-ISQ$#j]CY����)*�kt�[���Y%R��w��Y:؄7�P~���9J���9m-af���Υ��Q8�j�K��/v�-`l�����:X��諭�����=�ڤ�-]��|�\��˕�+kݗm���J
��r�����@ċ�z�/L'7�����7xbm[E��b�ܡ��_Ϛ�(��
G��#jf4:�����㚣��o��a�17�����3�8hrc6;|_9��Pƪ��؞к*��6���S^xE���'o��u�^�㭄�"�*�������JK♍u,1J�o���¼�����M�q�ܧU��gyC'2(Jdǥ�%f�!Ş��֋��}��7M�9C���s��T�ҞH��P�p;Hi�Vp@m�m5�(4b��
xh��Rx��RC����|��$��V��^��
G�.3	�AkMȹ*B[�mZp8�,��(?<�14!iʞ�C�{�9K���9�iw�b"iJ&:��bZ=����~;�Vhw�w>_z��I�g��Vюp��w��K��P��Yހ�e��d2����N� �f2�b�c�Q��:+�z��nؘb'y�a>�e��(X���*ջ��Qf�[�g�Z�D�@L>;u�d)��v�Y�I�{�Tx�*���-�9��`}%
xQB��R������NuLx�K�W�Ҙ�n�8s�M�N.t'a�͸qK
E����4��w@f)9�sfY�$����!0e�f�Dg^�{1v�j�)���Ÿ�dT�7�OP�Sv�,������>����3�Dנ��uE��}[&��.��1��H��'f͵ 6lK���(�&��9!<ͷO�Q#rp������c�\��:��S��
Oupw�'��_��1�p�I1��*y�Tb���+����2��ah��uF��*�	h�d�@Tgn��r������ǨߪDZ�� ����F�tB
�f7z�j�3~�4lŨ�#N�5n�o���3����H
��2r{h@�j�u���E=�X/�kEw���ʯ�h�7����,�9f�]�ρ��/i���]�T�"��2m������o)�~�W�Qљ�pš7�t�����K��g:���_��}CxϤ�1���o��v9�0�r��u\H个)f�7���Ƈ������r��z���?T}f5�wz�P����e#�Z5�<��::�H�������:�g�� ���j���&�Hu������u�q�׉���m�lc�{yTt8����1+���ju�L����e�f��:��8��<��O]ںN0�o��Y�s\�dY���O{ji�WȌ�ECFH5��+(��ז^��m�]fʬ�[uu�ҝ�B<�;}X�-S2�,F�F���WK���h�J��jb��u�s�G�x�MiS�q�PȆ��J���XD�}-?�_UUW٦�{w��0G�Uh��7>��:ۧp��?;W]�hW�2`���l�A_�Z�B�j����C�W_Kk�y������9�}H��� `��L���f�g�d�W�!{N�̜ק��_W!�sohI���	h�����K��T6l���V��S�"ME#,��bJ�w����E�!Ǥ->Be���,�~Iږ�ϟt�6���K�(��t��utcQ���}����tF�EWiȣ�Ny�F����_�P��k�&���!t[~����Y+&����nu�@x*l���d�7H֌&��A�Qxb/����+�u@�y���m�Z1��%��b�t!kݞ̢����UueFO���x��č�������K�4�O����f��c�Xb᪩D[�D�7QBECX+�|$黙|v�٨]����m�˩g�fk�ԵV�x�������y�0�uF��i���8��A��a��e���U���Y@������gq�q���b�vɱ���n��_D9����	
�D*t��,�y�Att����[�)f�6�n�E�(�R�2��R�[��B�wN�tq�6�S����F�Tܫ��w��������;��cɲpկ�NU��U��G+�|{{�*r��t%�R`���興�]SK�>@v\W�X���df�V��GG�N�O���*��q�q}���CG�Q��y;�.T])�'J���4ү��6�`��Ҋ���QW�M��K�{�-�^/`��U�N�h}t���Σ�j_v��������\>Zu]7�/�� _�\»(��J���a�V�nК���(��bn.�S�Z��lc�����h�ti<�.�O�ÝY�.\~���+�/�y_p�V���Q�%�j��۽��׬�L:8t�)"��J�Ӕ�Wt��@+��0�D����NW��	G������ѣn+Z��;oț�1j��hV��@@�"�q�K��Y�)�����l�2!Sh*����;#G�3�aw��"�U) _�v��9����זfXW�\�c�st��V��5w�e��Y4�:bvf2��"-�+�{d`U=y�q��^N�|��mV8
�!�������{AW�:����E�Q��@F��2Y�=�s	H9�(Wk�U�F�v)g�5�u�Jb<{p�Z�4[�+n�5�hE �=�R�+9�IRNJ.��ެ�n.ɮ�wR꿤�������X�.�{MR��]b���[�6a��u\�
�umf�*�-
�1���Po*�t=ڙ}5���Z��������������z�.71o�x�n�s|�yPt�K�x�5�f�Z@u9S��=�U�Vs���V�3���F�c�J��ڤ8�z��r�Ϩ�)��V.�YV����^YK*;��c�����;:��[���5X�s2w�oQĐ8^���&�m�=�\HQ�b�Խ���q+N�P���:��mC����ͨ�ͮj����j�����^����1�4|];�nv�֡��jg��t��
!��p�Cw���r�	\��8	!{�r'���l�׺�����#��}��˛ۇ���oQ����w-��Tc�+���nAjq�t�8�ڌ�/�2�TE�j�'�իv�5�ݟ7�
{��+����8��N5�9>螨=���2�LV�U�m}��-,p�26��pntH�+�.��ʅ덚N�`�����Q%��R�Qi��ܯ�Eg%��.�qz �]W�W�kβ�J�Wv��j��� iR�"�,3�����I�]+/�3�
���_\���U2Ԭ��0�ݭ��of̧���"�*��聹��7��}�	V��Z�:�j�%�5���ƨ��p����W�_}_T&�+�+س�n�8��������VK�rʞ��s�έjղ��J-o%�%����u������
�b��v"i!��5�Mp�C4:�uv��%*N�^�ո���p9%���o���O!U��)f9v@����❕���A�e���e�Mg-�U���������;>n���4��Z�z�j�vh3�D��~��9��[QʆT.f���M8�VʘTy��sDq��n���exe.V2>���y�i�����(�]�݊d��U���P6���V-�
���8�E�+�v�-%�n��K��Ӝ�S��1V+NqE����k�e}���W�q���~����C�ܝȈ��:��O��u��\\f���[��MFh�O����r�U4��;�˂X[/R��X��_mTc�u���6�$��o����C��^�n�����+m�R	��K3��߮�~?��WP0ڋk%E�9	����Lq6����}��Q,
�lכc�^�ydV�/"��H�q+JM�K��1չ�������\a����G����e̙���U���0�թ+��xO51�ŗ�M����͵��}}�G���1���:*�nè����ug[�T{��}���ќ�^^�ꌅ�{��1��h�~�9ets��>�_:n[U�Z�ʈ�m����ȕ��W��J���Oc�� �~�=�f�i򾆼�;hJ�~ΡX�g���ibq�mWtN�.���3m�U�?��{��Z��b)U�:�GeD�0R�s2*���2*v��w��Vv����p���M+�qݷ�2[��]:b��c��'E�q���ičr�=/໮7�tb�W�5��p��̨r�×L��V�.��(�v�m�>��8�^��t]��vf\��S��@y�����7U�r�X�^���]����Q�����	�^���O%���DĨ'j�;�Ĵt�q/!C�Ō𢷨��a�Y�ŏn*����ҳ��g���^nz�cg�=�D@L4�e�}��T^b�zz��|k�վ���]�`l���GM�9��4�ڥ�ԝ]���*ט�;��ׅX��Q`��[,���QT'��0>v�;ؒy��	wp�#�����ɥa�8�g�6-S��Z�{���o�>�">��;z҇\�	שW���Zڂ��uP�mdܣ��񥻚=��������rs��Ǵ���q�}�M�5%EC�v�ʚkT>n��,�ܡ��OWg�U`��"c���mROM^����QQʞ.4��iH��W�����g϶��%~g������6��������Oz���x}�E�jpr��2��Ӻ隆36��{�V��ܞ�8�H^�]]�i������w��15.չ~k����+��u�&��x}��v���5~[D|��퓝�L\��������kr!���MvM�q�"z��h�\���Yރ�?�y�g矩��'����_Z���c]��oi*�7�+m������V��!�ɞ8�mL�V������v�O��)�p��T[�j�㽢r�R�J6�W��p֬X�i��t\�'Ể��yx�_��u�� 9Ԉڹ��H��2;���U��{wY�R�^��o����f�H4$�ս�5n��s������$�Npk��ݶ0.�j�^ث�邞�������=��Τ�m���ۛ���jK�s��0JF�pb�Oxn�ax��^d�鍮�\8�;�}���}�7X�]�Z��ͥI�+%���!�P�w���3�����Zջ��3.�V�)�bk��(]�9�p2���۶\��R�d�O�XҮ����{�=.��Q��I�T[�yU��7h�7�$�=S܎-��^�G��o'uoT>���K�-1��Y��o^T���J���y�^zo>�u:�����BW2������`J6/mWi,Z5�"8)�|i�����X�'[������J��x�f��i�x��Bڷo2�ZX:��__����F/	�Q?wS{�'&�
�:�.��e*�1��-Ы���We}*�vŹ�Qn��{��Êa,��OmoWe����Z-_J]�^����hx�j�����2�M���C�6�p�݌�}/o9����О�7|��&�^��Ù��L�g@z���2�DY����v�߳{sк|��c&v癓A�c��G�n�g�Y2w|�gyQ�����Sn�\;���*aձ��I���-�j��sh�ѝi���L����F��}7z�v��i��\�p�`�i<�I�}��}�G>�\��o��j>��_E�!�o!Oy�����z<�}<�u����{�DI��9κ�_��b�m��d��Kt���v�PQ��U􌓡��zܧ�����z��:�s�%ۤ������T��޺�~̩3��ݙ�8]ai�c�ݷp4)���ʒ��
��]E���qFU V�Ju�����m�������㺭����%l�*��	G+��ϭd��z�5|�y��E;���s�8z겟So��q��Oͺe|���ב][�R*�N����t��1�����0�������k��3�����q�O�+E���}��XW=�:\ռ��TA]Q���ș��{����hb�9�ȶ��������8��.x`mMҳmإ�s'w�q�Ĵ��;j�m;��=�ו����Ĩ���I���o-g�-�oFM�j
"�y$Wf�9������KR�)��#��E� /i�K(����BG�=���gf��T*��u��YWds�[n���2�;{�M�%.�	�\�6�ڥ�?��*��8�^�F8���+1����*��F0���c�|{��o@���1��K�����5Gl� b�q��^�4,d�v[��	J>6���Y�r��E;�tJ�N�&�T�}W��ػU.���J#76�lq�bw:ܮ��|���l�{���mݝ��Vv�����ī��;$��i��w
��q_$�,X1�x��5�̮ٶP]�*g�0t5�a=�˽����ъ�ܺ"����*��i���p�jy`���Ud���8��k�E����ʅQ����ق�tg��*K��7��jM���Q[*b3>ͫ
�e�I�1��Tӫ Ln#�wa�/��d�͘]+�X�b�+zV�7W'P�&��-X�-P]έ���+dw}�̨Q�O";��&k<���L��X}LU����#����8
�����w(svVb	�P}fZ&m3No�h�iq�f�o�[�-��7*dW[��Qe@�[]1:N��v�f]#Z�yd0C[��Y*'�r�y�a�Dڕ7׭�e�W���[��k�z�T���#����"���͡ԩ�絼��R��>�\i_U������_] ��.IV�dӅ��m"�n���qv���\:���:쒅^p���
�m[��ֻf�Uk��m�nK�ݩ�u_P��9I��а�Ը�8�T��,�;�/�uں��z�Ӛen��&ON4�\]�V��6��9�N_8o{�V .�j"�ԦH���\�.}ݝ�3�E*���o���\�[�
��ỹ8���4��[�n�63�`��V���������W;�;UXiS`;�UYJ��]�7�W:A��2��pq"���¬�Vs$J]<�Cΰ#7.t7�&*Ef��� ��vj�h�Z�R�yx�Q�[c��RVc��_Ҭ��.��B�Hp����:�n��
�Y�@�㩋�h�Y��w�J���4�O�b���Ԧ�W.�n�ӊv��$�K������m�����mu�6ucՠK�e �a�D(]�ev��ƹ�A�Vc6x�٦P�`'@]��m>C,��&���2��<ej�A��'FsI`��� ��5I���Fv��h٠�˙2n���d�j��)�T/xlʹ��V��P��v��e_��-J����l��G�n�SD�7F	쫺�9��R�ӫW���w|�S��EC�WJ�"�.�3Z����m����:Y�s-ݻ��]�Wϓ�ͱ��x&�
�J�!S2��sU�{��Y5�*r�����P��K<S�'�V���z�O����1q��;��Mtᦕ�ZUԆ�Y�'���\���ǁ(/���`�ő�+�L`�fL 9�m�n�#>׺iڤ����tr�bLa��V]�/�vz���iMli��a�A@E��/ F��(Dr���΢d�!GU)*�ADF��º��̍����+�V���MB�(�(�2��R*�O�C�a�a�t,�gV�KJ��VU��J�LJ)S�(rN��f$�e���Eb�$em)���R踧Z��I��F����4�Q2R̪,�R�����t�
��rL�B�:b�u���%@P�K%�gH�j'�k\��J*�"�C*�Q�!"�Ne��R�GVE�e���Ŧ�4"�*N�&ҩYP�]Ee��d�.���*�"�$�]R�QP��Tj�B�wK�UQb�����ShZ$Ea!�QQI�P9`l�!L���֢�Y�j��&�Au���pH���t(�L�SB�2�0�����z�_�Aa���^Xz�B��Ϋ.�I���o\�|� M�eĈ���'�h�ݗ�e�k��Ϸ��{;e\��4��""#ಚ��}=l���=��(�v^�\&�PV�}9��M[̑�����}5�x9IJ4ރSv�\S�mT�V/W�X�Z;\T�uРҫs��fN��vRy2y<Z��/�(��ڝ��׹���~ImW�[w4�fJ�^���X>�s�w�;c�U�{q�ب�K-��Wl#SMS�:��f�Υ��n`z*��Jsr���Q��]e�n�'�y;�ը�6��y�k���B���q�uC�J�pڕ+Z��_o����ש�F�!7j2�ӵ�vr�rn���:k:����Ī�ݕ�w�_%�);�H��ۧ��������O/.�m�D)�t�^CP���eK�����\�sY�1W݂�v�F>�oa�������,oL��'&;uCJ|�>���j뗰�'��x�]3����OzN4�K>�o��|E�KW�S	�k�x�O;nWPڤ�-.��G��֬��^,�Jj�3���H��LΎ�'x\��R�^��(Ӯ���B�*���]�s�ս��]4ˏ,���97z�'V1���Xn��*�WD��B��5p�G;���{��ۏϢ">��S�5,d�=�<89�{fG7wvn�kN(Z�B/4+ݺ3=#���8*��k�jz��"�O��A�~���y	���_so�������N�[��+Y78�[�nn9��,��j-��Ӷf/��j�pua��T�)/i�y��_'U�P�.�r a6:��Kj�:�+�d�Y���[ݝ%�i�z�r����Q�K��	������ӝ?�{3�,vo��T^v֭�guy�5u*c{�Zxs�۪�Uw�V�j��@�Ǖ:�-:�T����u�'��CCk�{ϥ:R�V�w�ħD�=R+[S���B�B���ϒ�^4��޲�<�=�-NE���b��-����J�u�y�d�]�B����=��j�˞���y�<�Яv�n�{cj;0w
���>��]SE�e��n��f�ri���û��Q���h8����Z%�fqe��^�;�F�	�A�έ���C�oJmVVf['�+!�5S�OC���V�J��K���R[tj's���T�ȅ�̥�#���+\͈6#�ea���U�N�u��[�U}��W�!�!�V�'}�W\�w��u�|��;{IQ��'|�KM����5�����>y;�T�:��֕��:�X����m�)�W���fr�u,]�BO�+	<�tU9��2���\��Д���ǻx��Tks�����.�����x!-�l\�Ln�����|r!'�4�Z�.�ڋn�V���#z2b�*n�Wa*������=��v���k�Ӭ���r�
�w��y8��pK縭��R�GB��"�����;�.�����Voq��>s��<B����M)g�����cQ~R���̙�ή�]ӎ�7���ٯ�Nj
������Y�c�;93f��c���y��g�Ϗ��L�N�Ϲ�T4��F�	��n�t8G�9gk�Jŀ�/!]A{�[��U�c1؝%g�{/�u�-%�v<���s����ǬV��J؋>�{�eL�P%ɀ��{K,,{�֍�w[�ĭ��C�8r �%�4��s�/xe��������;npR$ɭvzó �.�\�gf��m������U-����9��ՙ+�08����ve�f��3�}D}�6��S���W��+�;P���\���c������5�-7�0��_K��k/1�h��A�����]:��O(��#���e��n�����+7�F?��sR��_��e9�%�Uݱ_qN���5y^�i)��TE�P�En��^��O��:1T.����Z��{MvS���XQ�Imsku���S�z��ld�s�6���:�ʎ�ˈ\��C��㼘�lA��ɶ��1d�$��7/;�VM�\&
���,�;��.�Ԧ'w���D�HC*� �ה�4cE����~��C�-Ρ��&����O7����ع[ys/�܇�|��9��8�U�(��#�G�D��ºη<�%��y�/9��݅�O�U�ҷ�8�S�jS
�Nʷ�k&Nt�W�tS�����q����&������jgzy��T�K7�y��z�f��5ع��0L񡓦6���0ʺ�Δ{�_J�3�8"=ǶE�e-W��tăˊ��9�nz���.�r��>��n(J�����I��k��YwD2L�3q�)�`�PI���m�c����x�Ǔ������!�z�fE6.;����ꯆ�ڧq��g��D�+��z���.��<a\5
`S� P����*�Ar��SUa��`�+r�<ˀ�{�i��=櫅
���S�1�
5�\M:g����{)�[�2���8��KGuah�@̼�f�R�QԲlˌ��,�s�~Zi���Y�'�}�K���Iz���tmxˌƳ�y�vѾ躵��1q�F�V�oo@����zd��yh��}烙7u����Q�=+V]_�f��������Tǁc˾X�?p�o5�+�'���Q?_R��O���{[5�x3\��`ըy�ٞ�f�	��r�i���c΋{��y��e�z��p66&z~KR�˨�:�������6��{*�vh>=N@���{�G��`����S\�s��o{Ǚ��W9Wt����V�r�;mL�K=�\�g~�����R��e����vʖ���OD��۝�Uu�6�v�L�K'��r'����`�t������)S�V����;]}/yXS%w[sZ���墮�3�&�s����t7~y�����3��Y�cZ82[\n��ޠ��v���;�c�&����ﾁqO�ѵ�Y[��o������1�p��bPPbw��_gcW�S]z����}<���jyq�ko9M*�4;.9�Q��1T�G!9�5�Ԏek+���z�[O/L+{Q4��ܷ���h�o�=ު�EU�����:T�ϯ�Ol��i����y�+ԠZ����%�s�J���34'�:`GV鸁�݅�Q��]�Ju���o/�뚫y���7<�l�q���C>�(�t.����yu}�U��k4����=:��'x^���:��g�sq�ܩgG|Wm[V���f�:E������jH��=�O|6/�����U�{q\:��	i�����ԫs1x�

�(y?w������{O=��w��nR.:@���X�t)���O�D��ѪA^�Ҽ�󱚻����RTW�Q�o)����b�Y�s�'�tkĶmh��``�7j`τ�le"O0�{t�:U�����R	W{�}�]\�+y��B�t�G8�$���kS�>#r��8s�p�Vc��-������Lc*XI��;G��;�;����C[�Uv��ti������jw���D|�=M[��M���]�Pq][�W��������U�
M��7Og\wz���ݽ�\.a 3*Y_�N(|
]K��}O���ti��7ݩ�{^���<��y=�C3k���^�mߴǜs㋍�5��^�����{��-E�Up���V\g4*/R�oYu���]��B{���^�^֨�Y-���u��Ues�67��5���B�츏y\���q�'�j����9�[�8ˉ���,�W�Π��p7��ɭ��Ԫ���SA���`O.��Q�GN7bv�Ge}��L_%�+�'σJ�,�u�Z2�ǝU_7]/��4��3a��0�|:;*$��+�i��ʷ$��P+�f�)���Ř|�W���[��߽�|"�V��Ζ���l���^�]���ɋD���M�v��S�]5�}m�c�U�[�I��.�1�k� "�E	z�s]��LMx#�7�{9��C�a�S mՎ��Y����݇Aw.�� �D#}X���7�xv�<�$з�#�^8�\ɬ��%���ō9	}K-;��i�8֕�Q��/h+;\�n��,⮜"z�^Ln�
3 Èurg����n��C��zi�1;���c�XX�_�=�p32�E�V�p�N��ޥ�hG~0͏�Y󽤱Xl����q���8jQ��n���n�'���溼�oo.�7�z���A.^͓�]��&%��u1S[B8��ؗj�G�b�W@>L,�M>���x��,{S�V||.W�Εk��z�t"����窊�v��v�����_�Zʈ8�yob�r���`(Ŏ��l��t��LB��:���kG|�Ω��e>r�+���z�=��W��nnޟg'3�~��ި�B�N��V���Oz�\խ�+n��]x��i�E�@E��90�H�r�}kj��%���6S�����k��(���ٺ.o�iG`�pn©ޛ�U��u�
�S���z�bw�;fp����Kr����N����]_-�TkF�Z�}y;��Po]�\���x�Є��]��b>60���dڂr�"=��!T�9?(��X߻|�ӾL�:�S7-��#�wJV}�r�0ic�G�����L���k��R���� ��;��nʉ��cD���V�KF[��si��&��Շ^�W cxHs>�u�������c}���8��_�ݧ���]y�v�Qnur��ɧ'�t�Gف��׮ ٳ�-(}^��}�{S7�jn#*���Q%��.HQ�zqͩ6��Rם=Ϸ���i���v�c�n[�'Í!]�����[U��^7��o�N)S������]0�xMB��hW�e�5�R���73�R��]���5A����L��w��4�t�AZ݇z:��X����hS�i4Gf����"~}�Q���[�a<�U��>MUA��͜Iĸ�F�
]:\l�j��T΀�:�O�ٱ���_�[Ec�ka�O%U��fhv�sP�*��P1׿�hoM���G�������p�jJ���o���A�6�5��VS��W�C���)�qG�*gZ&gOc���"���Z���ۆ��z/"��]�)K�O��نl������$���}L����5�g�XSW[vt���߻�k����Zn"]���n��;���$7#�s{c1vB]J��{�[���-v}��u���\Pzٚ��]z�Q�AWL��V�(�5q�ӼK'ku�DˣG�|39�n�}��|{Rޯ{U`�[����m.��}Fu(������~��:��ъ�q��2���>}N�ī�?V�\v�(}1�.��\�k9�O-n�sa��p�MSj����t�}ב^�+l�m�Oe]�/j�o�Ux{�굦��E��LԼ�Hp������W�5�;,%���*V�VqE��ңt��v����y��e�qS��[i�t�S]�m����J�[ƾ��k��|qP>�_�EE�y�W�1I�F�US����q����б0����2��(U��)�Z�Ц�U��cr�"����ҭ뿂i\F8}����3K�n��կ�V[��X��91в��0���<���bU��P�k[�#A��l7=YַRՃZ�
�x�.�Y��t̾�&��&�{+������Ei�r����9S�f0���[�?R�b��]�c��,Vs�7藫沣�`�fÆ�ni��%*��ei�Atn��F��o�u;q����M�SVN��n+���w�X/��_6J���r�F���Vc�P)�x*]μ`U�7�������/k�y\R�JV./H�dOuS�ś�d�{Q�x�9�Ʉ�Z/&
���3��YI��}������T�h5����#<��3@cEz�w*�^se�ҮM�|���8_�7��1X�d�t�.:��y��� ��JK­0:��E��Yhd���U��3*���e��V��iZhu��0w1�̺�ؓ�5&�[�{�W)}y+��n�7���mK趮�t�;FCճ��Z�Pt�d��Y&w�T����Y��csq��s̬���:5Z��ņB���Z���<S����W�r�%9-�?B��߭���q6��B�K��u�h��a$�^�#�� �J�Z5��$�}��7(U1V3�ڽ���`����T���1�v�� oU�e�h����i[�d�s\��y>�-F��CU�:�i�E3�KtO�Tz_xm�6�3ƹ!��C'�iUIZ2�����@��܎���V��<T����vT���9٭6��@c:O�����S.����k9q{���9���ю�U+�Ի����1Vb���|�`�Z������}����-�ݏ*ѧ|$�o3������i�V��I�ﻕ�4cF�k8KM�V���LL�C/:t����w�46k]mv��!YN��8ؠ����q�bqn��-K���:CiV텊�y*v�c_}`(Mcwt��
�l �j��8����
p�ʭ���̻e��{� ��L@�0��T���;N7=PK0�]���`N�a�g�z]ɔ,7[�v۸��z2u�ui]oD���c|�2x��=%5F�p�ˀ��}�V���8�p%h�`_]a�)4����!��C�Y����hJ�|	'�Z�3��K�n�t������[�{�S���s�9� �@���.�)=tw\C�d쮕:��1lm�.�	e>�*L����
���������;�����Rv�]�j~�՛�-ޮL6�v�2H:.��7m�$ܙO���װ��+7y���kMM�4g7(���Q+����Ur�k�Q�q����{��9Gu�`�P9{j��u�v��B=���������.V>�5�qBĔK�O:���>�u�d�<�ғ1P��`r����)gf⬎Dŋ<���(G[{SL�@*ؒ3��=Վ�އU���33��sGm����h�����p=c��̻g�4��7��okpZ[���.�)���¡���}(�j�\#3�cT�Yi��;j�;��_%�y����v�ܼ��t�;�Ѭ\\lK96V��j��v�E���n��Y%]�ʛ6s��v�
奜��&�;a��^Ho�l�-r�Wuu8qa��E�-�x"q�V0R��1B�ĝ�2�-D�Q�(R^(�Nʾ�9�-mDi�(�٦����yhjIj)XRE�4%e�+$�,��J�i�"-ZY�J�!E�V�^�UI��Qd��Z��ˡ��R��'%ĻU
Ȳ���UDXj$jIH�Y�J��U'B+K�ˡ���X%r2gGA۩���"�\El�U���d��H٧MC��"�Y�w)Щ��I&%ʨ�U�T+�X�kE2��(�C�Yi�2�ZYEU�,�
i�HVS(�s�U�D1��]V��VVA�Qg!9v�r�h�)M�!�S"N�3E��L�Ze�EU ���D��PS"�Ȉ��l�@��� �4H��7�w�}���Y]��1`�H�L�[ٚ��f��uY:�+K³M�/x3���)[Svb���Xl�j�?��>��1��o����ZV�,�kV!�&8W�vQ���ǉ�(�U�Ҟ�H��ztl����:w�j�W��:�CBQ:�t[#|��S0�Us���ż�c�zg�x�s͏�PtԕO��p�25}onZ�'܇ q�yeJ���W�j j�j19����\s�t��=2�e�%x��W1�ٳ������j>]�b�����z�o�������l��UsK5^��[�/�9o=�M����]���h\t��*1F>��YXr���o���#�2�f��B�!�6��_M|��X7l�θ�8qs� ~)f=��9Zy`^R��Q}��sR���lO�\�䯸�m�3���$��I���w[Vs��=�j�й��w��o{*�5���ȹvH�}��XJ7%�\�A�ia�Q:�}g���cV�Ҟc庝��{�ڎ')،��E(!����<C8��Պj�\�Kk;z��-��4={�qQJ��ş�;���{)�j��񭻭:��y=�ui���!YI܃;e\v�������7�^�а[������(i���%Y�0���t��Ϙ����2�d�Ȇ������}K�n�i��'��1�P�J����Q*JLU�Ur����;�KHݫQ{0�`���y�p���&����o��*vܨ��#��{��tÓ�6ӭ4�y�w�ͽ���ږ��Kd�:JٶVK�rBW=���Dײ�չr;sfi]3����s��;K_T�B��:W_q�-�1�oT��s|��e�����ˁ��p�����v!֞B�c)K<)�N*k>���&�S�4�<��b{rj1=ۀ�{�}	�������V%�X��6���U�EC��WŬ�>�4��,s]�k��\�$��.��Lu�x��9�փ��T��\�F�T^b�+�)r��G�\p��V֣��NtYYO6�m����u�O_�����8�W���qN�f�$wv��������D�M�58�41�L�oT>p.��.4�I��c�MA�m<�W����}w�&+��Z��(i����V @Xz��b�IWv��|����ػ�sJ��2�\��{��f�ʓ%��eڼ��+�d���egi���S�����+CVc&��,�n�!A�V9�%Y��f>/\��w"�[1x��5Fg�E�}���9�ݰw�p���m�J}B�f�o�v~퉞�ٴ���t��bc;�A�_����S�r�S��Q}��--/g6)���y���n�ׯ<��o{�ϔ�N7.z�V��ݍ�N�U{��U��syP��ǩ�J�xh���v�~쾞�y}㋗�LA�Q��kUy;�'�T�y�W�b�Z+���s��t_W���]�|��������Vk�>9v&�wUY��:���k���n�VK�\�&�}��m�������[Q�W�c����`ȍ�g��������"�%��|�~�4�\wm㌖���0���Bt&�{c�2�ͫ8L-NL��p�խ_+/���}��N�h]l{HƩ�͜�m6�Vzc�\Y1]2���.iwN�Z��w���ʌU�N�wu8ư(��)�c#�mA�����<ˀ�{�oy����`�7��By؆���n���k���V��s4�cYY��%o�(��Be��Յ8�K�]��5{�"�	�!J3��Z��T���Y�+��y��Yg�I�w;w�Z�^$� ���Z�8�����"iN�ݿ���U7�ʆV�>Xq~�}�{�q�V,g���_[l=��3�,{޴i��t���mٕٷwx�(uCyU8}e\:
�i���8���]�y6/�Y/;���ڥ��K���O���5%6�浔� +_�PV��$�1I����J��f��]��O����՟C�����[���B�+'��6)u���R �<��<�
ū�ƗՆoV�N��j��oQy�xE��M&�'�̅��Y�)<�?�q�8���7iu/t�&���{6��T�g-���ovW��>��=6t׶5+�ݍ<�ڡo�G)���95s\�]9X�j�nu^%]�lk�f����T�h����*+E��q��4�N�JN�F9ꁍe�i��q�����CȞ�K�YBb��0�|#i���+��;*�&��y<��:�_�Sˌp�no{6q��+�����5�wK{]I�z��%�y)�+��� �EՓ+3��Z��4��3p�,)����2]�=Q�VN;�9jx�D9WK�7��ַ��]=n������~
%]�{��km;2Pl��̖���Y�b�<ak��6�;��p[w�UCf�7V� x8̨�R�W�e���,}6SJ�>ʴ�r���R������в��UBv#��6n\+�\��O����󹸮�gnN�v*Y�3�)J8ܲ�0�U��s�f}ve�bnʺc3}@�#�S�q��	�,��//����Tq��Pc��p1+^#	�$��V�R��k7�f񌶟>s����>�ް����(��/�)�)SHm��4�B�`5�8��5��s�AW'N�z��C�4�YX���˶.w�O��?�>��1_i�ǎW<��A�J�mC�*]cw�W��������]�_A����U�kV�;z��
��Rz\�3Xr;Xy�_s��U������z�R0�;T=��G˶�ū��}L���es�y��͌��l���{{5��h���8���P�_:6����V0k��ˇ�V���n�A����|Z���m�k� E�Y�^�F��'�Ъ�˚D��T�ީ���D���x�ۓ*u��lN�^�\���i1	��%��b�8w(��Mp��o�g����m0P����H\HȾY�.F��l)W_����r���7�?|16��*}}+ln��v˼�1Ք��䕝�j6x۱�ߔ���LE�\�:5Ž�x�}�F�K�5o�z�/#�Fг��R������Um���k�[�����WQ��fp���?�nuc�"'r�ժ����c��@XL�V�:꼫��r�z�k�am�Ī=���LU�N�.��o�}-�3l<zL��渔�:��.�c�0�CHT�L����zw*����t~���g l��9!��r�5�W�i��)����w1Y��j2�[+jX�v���{ѱ6qoO���WI�L�����q�1TE����.�R��NÛ�f1�6�Ѕ�#,��Ya�e��rI��z!�	�*����#)��%��Y�^�g)�b��e��")�[�i�pW;�:O��P�ӳ]�b��(�N�%�j3����$�{�����5�]��狦�%�v6-�ܫ9#D��T  n3Vh��u˕�����Zu;�v�t�]����t����2�.��"9��vi+\�Q`d���s��pr����
=bD�|��&�gi��0Iٮ�;umnw|<�I��X�mm���
5�\Sc���Q��^���Ŏk��[]�ƽJ�9I���W�T�4V��p9�� +���Pw�J]�W�.V#�^iV�ź��b\�Լ�m�OTߛ�v���%���ߴ��f��J�It:=o�W'�3���+��;�P�[�2�
Y�
�+V���ع��;��W�K���iz����3z���vz'�fr6o����?v&a�^��u���+ƫ!ώ.�>ڬQ���͇t�\rm��5F�)����>�w�DT&��f�����B����Ue�otOwf��l������{[�����2���3�Cγ����u~�"w�,��I��z�Dѐ�6�V�����Zⓟ�U�TsȞ������ށ�g�,�:�w:/)�l���>w��p�9���{l-�
zGdwU8!�M/E���mi�p�f��W�\b�t��05� 3w���d9b�%p�d�!��ʒЙ�� �V%/t�݁�W�t�WPSf=��m��PCxM����޹���r���wuA���q���+pE�!����]߸�o<&X�4O��^�<$����OÜ�����%ҭ��4���v�׻P庎��V=�:�(�Ky�h��x�P�\��>����w���M|��_��q�0�n��Ś�R��a��5�aeq�]�@Q#Lw�D����p�V�H�JE��X6F���e�B(����W+s!;.��=�[ݖ��t;��x�k��,n���W_7q1J��qv�[L>����H)�Q���oy3]���s�}e�&&a���\:
�����D��bg��4ޒ2ꔬ�Z���Ǿ��1�{}�T5%Sj�YN�+~|]`ފ��������]���o�I�(q���f"�D��M�WR��c]39d�Q^����Trl��x���P�h^;Gϴ�ʌOMEꉋ�Q_rx�f-�p J:������wsɕ�<�m{��hx����6-�V(�P�Ƙ��fSS71�SO/z'�Ʊ�Ŧ7�M�%s�d�}*��7�@�֨����,���q4Ȕ5��ِ�U{�O���<��^����j� ��H Mp�}�7t}7�^ s�lu��%���
;�ۨts��eM��ZE,�7'b�tf���y,��*b=�r������R�<��K��<�.qU�s!�΀J�lӵM1��l*鬃/zr���}m>�W�M��^��#}�luO/��=���Z\+Ҳ�F���gU+���i�(v���Z���=�FE������{��[Qs�����K����_��pu<p��[�y�X���T��*cF���u�*9f�/���R��\/���]0���X���q"0�=��$w��Ip9B5��7p͆�Q��}.d%��;��ҷ8˛޽��!��M��	�����ş��5J/%�#�T���>�]t�a���e���66��e��[�z9��v�D�B'�vW�;�Eoo<��|Oݞv{f�s���}˟'J��^�m�§�Qg@KΑ�)�G,fP�2�6z-����K&�1=�U�oP\��}T& md�Z���#����4��0Ń�Z�4L� Ww\l5{-XjkL*a�7GIO&J84��*�W��h�s&q���V�,L�Yv�AԽ|�@Y����:���v$���[\�gv��u=�o�M̀�N��Ƈ��_�/e�v���	B��q���G;Jet�v��v�XtF���;h�Kq��go ���^sTR�G�e.^����5;o��������f6_l�pefv�8ҳ+*��ۇj�5�P�����%�Ī����}K�MG��(������Z2�\{���?��lt}����������x�먷o0��S��YZ���]*��9ֆT}ކc�봶��h\t���8*�l<���2�o���E��Ҟ��v}�����m��+n��J#n����f��槩h�*^�YŊ-�˥��sb���>O��k��k�u�9_�tR�V�>�4N�vJS}N��*�/���[k����kq�Ъ�*�O�b��ꐹK��]P�%T�5��N�c����V��Jx3�Vo3�K]�=9�����m[�W�в��������I����p�A�R�5���W���W���Z̷���f����t���ѕTF6c�9��6���g[ϙW䨾��i/���%�K������O��άw+v�i�"u�}K,�Yn�\zڻ�,��6WeZk"]v��$��o5��&+v�g�H<y�� �n[w�ۣ��&vK�OWZ\��֐�G�IJ]���-��T�����D��3/�e⻴Ùټ'8���|ʻ`���v
��HT��vf��n�E�*b�VN�u�f_R�A�(�N<�>ᗿJ�kދa3��B��|֖%�f�Z��-B�'6T���nIn�*�����8\�U?����邓
�.��V��D�xv�6����2�-�ǻ��2�t�nqD��u��m��}L�@d|��ucU�P��������
��`��v��v�6�2�!��<w����a��"�-�IN=��K�wwm�"n�n�v�s
į3Hu�+Ml���e󝖭CCM$PV�'���%�8�ۥ��f�7tq�Ŕ��wp�ŝ)�QB*:
�K�[iqTgoi���g�"B��������=Ku�)�ӟb�=��48��~�Z��׮�o%�2Qt�u�f1]�m��[�#���ܢ����gRLJ��ΡB*���ܷѲ%b��yh�`��}�6����̥ڌ�O�#��n.�w%����0�YBq9Ձ�(��	N�3#V��2���噓9U�]I\���yVAYQ���0曵�&�Yp.P}�¬NöY���VW(	wα��^.Z�C�+oq�V>�/�W�͑fI ��\L�FEu�ݮ�t�mp�0u	��\�/g�m�c��N�6v��R�Ty�z&�Ե��sԢ��]>li�"s��fJ�O����y�B�r�J]ԝbeE�\+iV��x�zE %����݌!��ɿ�3nS�Y���p]���N+ N�AFU⨸9Q;��He����Qk�]�.N�b���4Js8�y�s����
����Uܳ+x����de�̖y�3��a���Y}JQj�bW�a���0l���t8-�b�G@�2�;����I��P�����L8,��Q/�U��wcqqG���|�c}���<�iw"��pN����0P!��r�"_10�v�G*u�-�7�ܻ<�;Έ6�ʒ�L;2��Nҡ�C�Rt'k'a��eY%�]l�u�5�4έr��i,��:�#/�rɍ	ŕ_�ߵۖ=�ޗ�*	��s�iS���S2vB�p��i�KV����3�].-0wi�+�J��:�/�k;VJ]!>��s	B@���M�H����zD�t3�Qh��]�"������g��q��.t��]�N|�Lw#AF��C�^�5K�>�n��;����@[�%��G�a�9Ki��fn�R�(�C���+۾<�ܵ-��O�1��y�Q�w)�CKY��ԙm�2��]�&�I�>0ve�аLt�'�e��٧�,�����]{8��v�b6�hZ{&4y��]�������*�.	mu���,��h���k0�����=8Q�|O�	z�D�	�	"̩V��+�QE�ӂM&�I"�+R�醂T�ȋ���bAu6TAE�8�H����$���H�J��(�
�&d�XFĐ���Q�r�Y�
"�"�M�i��aVp�H�feI�s:HHE	�����IRXT��T��M!*�N*�d���EɔamL�J�A*��դDYa��2#���E$���)�*�e��- �I-hjk�T�Z��T5��aBG��S��琓�˕J�9�B*�����Ҁ��KۓsVfUEDAAIj��!0�*U���I�V�:�В#**��`�0Ԏ�Up�RL��Ͽ��=y���y����.�d��H&�@�šoM��|v��&1pk`������dm�&�3�z�)z:Qg�PYN�Z��Y�I����+7V�����x�SIF8ֱ��:I�L��BS9'��mE���Ч���ݧ7��>���M|�_7���ql�V�p���i��Z{^H�+���L�Z�^LR��ypf\�.�p�+qhwBj��u:��E޾X����B��[4��[�Q���W?o0��s[���C)�;6��k��L��TBw��f�z=�h���!�.^�9z�s�0�l�����3V9�ơ�%��5��ǣ��E.Ҽ/"��X�M�{M�"9J��h�p�۽R=Pv�o)�V.��	e���8��]�F�;{��7��rN�r� g���M�mh膆�]��ޗ~�2z�0�񲠴�=ܽ���gL~ұmR�/m��=���=:zoI����t�m/��z�c�cE<���C�r���>{��v��2��~[�`e�d8v�����V%�4HF�����
�z��`KR���-S��En���l�9�8M�r��]r�#��;B��at�a_>��	Պ��$Vs36�Z���׫iX���-�΁�|ի��B[ط��QunQvL�P����hm��{������g���J���6��7��!{~>����Y�FE�;���!a�{�NS�-ڴ�E�������Cγ���c���i�1 R(�*�^5��e�R�p1���\��|��&���!�J���R����N���'9��	��w��y-�����k2#}]^�s�/o��2=���}�r���������M���Q|�\b�V�Zi/��v�8�n��to%T�/�W>n�oa�ޠU��u�&e\�&�����h�o~O��y�p�W�z���:�jQA?�ie���������?��u���;��;7�kY��5�FW��q{�G�ǞB�C")J1]�By\ҷ2�ap���7b�)%��{��c�l��5SP�3_9y	��Lh������΄Rһ��ny-o��%�'��׾�8�߷�L�CjYW��%�;.��Y�*E(�6���3�/���諁�ku� rB�����繋7�8�v�r�x#�1��\�̭[N��Q1��W�M��9\���0�ř�bޒ�N����CR�7�:���.oQKc��6��7X�9�zU��w}4+��0�N�g.T�f������n�����T}�QI��%.�xA���kɭvo_C\������m�*�{Q���M�RTT=GNKo
�yuؒ��\�tˎ�Q�������ϴ�[V��}B�oRX�|��L�n7�ݎ���H5\v���±�m��.;��6���.��J0�M�y\d�1b|���+�R���kޓk�fy�iX�Pn��D���e�����w	l�td>�l�݇�{��Dsbi�z��]��VXK����1�ѥЫ�1���ʴv��YΫ=�ΪV5���[���|����Zڡ������_8�Ը��be�Xj%Dꋧ�a��uj��w'�kq���FF	&�	����GVT�釵�ueF�)p����O�޻��FoQ�U��F��C�%��DU���N����J0%�:TK���
�\������ងM5��=7C<�ֱZ��%X�Ixm�.����T�f6h̻��`��z��&�ĳ� #qe<�ް�����b�a���ևm˸��-乡,|Y���2�ʕ�]� �����N!2`��<\��V�cr�9�����Nx��5�������N��nYX!.���}r�E�X���.�\�u�-�#�j{�L�������b�C)J1л6s�s�#+p�3�k�����a,ˈ���͞���e�p�ҥ,�nok<�˻�epi�E��O3�²�Π�9u8{q���>�Ia�Fu;��1bL������A}����u}oN,s���G*����Jv7:oy;q;�Jgf��v��unQ��-m���V�1X���٘Qٙ&M!�;r�+-]n;�8�i���t��c�>���z�Y���S�^m	���D�q��Է��.�ه��_7�+�ܢ�(�P+���/[R5G�y1�ԝ(_R����>�{ޛNG��~�m��9cW{��-���*U��蜹����1F*����9�P�>�w���휭��HU��Dۛ���Vۮ�{�ڰ2��~+λ��ul�j���1^��t���%߯d�A�\�$�u���ok<;:����w<�1o^��U�������r����yf��:�56���yPm8��y)�z�+P7{�̾�L�8�T;׷r���PѴ�n�1�Z�����4���&��{��o�g��>ǵ��e�w�*bo$4���{�rU;�E���k���y�W��dQ�	�>o`s�aW�H}�k��ٝ�����S\�8�Z��z;*"TJ�Z�;�z�Y���k�(��{�9�5g��5#�K�p�*5�˙ߺ�wܷ��X<=�LT�/.t��������:�>�W�4�J��r�.W&m�a��m8�>�32�ٯ}ɿ{[����Ùi���>�}ҏsJ =���Z�_����Ǥ`���k;�]��U�E|+�10�}H�����9�-�ǫ��#ឥW�m0S���ŏ9vwr��J1��0;�� ��W��r&Z=s >7�c)�m��{�L<5�¼���#��uv���ǩd���Xo�� �<�
u�$��͆:�h�W��5^�Q����H�Ȭ���י��������u�����sf��t�ϥ�`�;G��+A�����\fև]`�fjE�(��;�Q���ؤa#��ck�����V��2�׆7M����R��]8)��Xo�X�Ҙd��ru�LS6ҬQ�c_q�{W^n;dw+Xr9s�msf�g�ws��6[��f�.T�]2���E�Iܭ��cYb��A����4K�8�so����>��fk��Sϝ�ǭz����z*x���q���a�2��I�;����O}7�`��Ŀ�����s���?,w�}������J����Z��'J�vU����Θ9�+�&Uv����Z�JZH�>��;q�.#)�c4��5��ζbW����M��\]�	w77�cUg{y�-�<�Eh�{O}'�ueT<9;0�#=]`�e����v�\_>� k!6�PkZ����o.��Y�(�9�r�ǞZ2<�R�ݢ�b�L�<��;ɝ���}2�n�Ց�ꌏ+W���n>���?}�_���ʧ��Ǫ;�/7|3�E ��N��@��T�����𪃞ntk�����15�{s�GIH�'�Vu�9�K�h�ϴ�uj�r9�V{�
f�T���b%h>b|���M��?}sh�/����ږ?\yz��|����K���]za��z�1כ�Mv���>Y���ǝ���$/L�Q7W�܅�ø�����凾��=���O�e�z �=�r���Vz2���B����͓��ER�z�%��ͨj�ZF�ïRD�F�&�CK�{���خ������9YI�RV������R+�}��F����psψT�&s��,)���Uo0���obewd)����ોvtͷGLk��)���E�i�f:
���-���8�QDg��SF��Gz�:<,�W��W\7�V�f�z��r�4[�R7������r�d���4*��9�&��k̎Ȁz.}��=Д��6�_�����x~��箈�uNH�!����,z��?S�Ӽ��K1�׷佴q2ϼ�*=p�������N}��W�����ID|uM���������veM��.g��}��dV��{c*#�`�|��s�{�M�,z��$ל�����{�	�;Q�n�'W�����X���Y�$ֹ�f�[�����軋�=�Bzo�jǩ�!1Sö�z���*��}��7}�nv�޿�+tü��ޞz6�R�_�&�����)p>�gF��JnmO6{�v��`^Ѝ�D���V�4�6�����=l��ߴ�(?�=/�z��Z��۳����w�{�����h�{G�dL�f���3'jFO�ίF�	a[��?!�~ο`
�g��s����l�^�Ǒ*��|���������U!畳i���U{�z��6Z����󘿵HNn{�cr���S�\u��z�F������?��6�R� eX�]w�;��rVR ���Y�X��+hf-�;�W?R��v�l
�Qj�;�u���f}կ-v�7)^R�S��L`h�Qo2[�Q�{�[}Z���v��i��;�Ķ�k�����g8��',D�%��p������Gz!=�N����lߢ� ��|P�wǾɟ"�"y݇��x���x�ܿ�z�dy����v�Yۗ��ԣ�F��*��I�T̰3�D
���^}�P�g��c?^���b�Y�up����F�fe޽u��P��GUޏs��vC�Y��Pn&�����q�x�ن�y��Oy��Sf�7�ݰ�o�d����{�|8\G���j�,��	��k�B��H�%���<U=�s'�}�:�5Χ�wW�d���*�^��G�!�o�tT_�܁{��]ƙ� s9�J�y��ί<�f��V���Z��s׵�ӝҙq�Tuî�x��};ģ�{ޣ�ѵ67�2�_(/����"��75���t6�=rl�}JS:2��s�XʈKև�=T��}��3����ʂ��MUH���s��^����<���$�ǍL.߲�LM5[F�5χv|%���J�K�|G��9��ZN�S��xw��vAؤ	>G6&�_�[�竤��^�U���p��W�uE\Q�k5���s�em[�>�tC�"�z�Dy�Q��e��3a��Fn�;�ͯq���őU�ڙT�߄
��	AZ�sV��qGPe�&�G��pk�x�i���$a�s��J����YE����&����{^�ն���׺�e�����H<ԡ<��;Jn^Ŵ�����2�rx���}x�;�^9jnV�<���L/�t}ۙlc�]�#>�K�G�����M��Q˙�ZnvX��V�o�/OW���B�[���T`��{��>�X}3Ft�
�~���g�Q�'�{��*���ΛGǧA�C.���:�)�䄩��M3�P�;������`u���=Z���^��Z����Y�ߵ�~�+ٞY�������;�}2��}�Z|/&w����>�R=����C�>��\9���(n;�׮�\[Y(����l��E6r"Na=qUƱ]1q3��L�'��َƽ~�1U\�5��M��(��o�O���\?~�I���A>�.TD�	M�P����\;�2�yU���$<������p�h��v�(������]1�Mux?��{#ޠ)�@-�������7�ҍ/p~�\r��g=47���y\{�6s}#Ǹ�F�_Mz�:�^F��eH}܄{�n�zF�z�{{�!:��;ҩ"o��s��V����~�=�|��}^�p��)��#r��J��}�GZ��1�G�ٟI�_�Å���>	<V�[��3��E�o�|���++NL/v*��V����k7H�Tze;���^t���fF_8g����\{8<���IîIU��-�\��*d31��3_B��9��}�+��GVgy6�]�Nԩz/)tJq��:x5�2�^�i�Z�dӖ^\D�^�>%,��%!}�g�����yߢbaz��D�����%���%�St����w�u�q=sڹ�>��Ĩo�����\5��"e�����_��>���_�v	��V�p�(Gdd����z�w�C��V�:݅� �t�[�\�r&|_�l1כD:��V��h��G��Nou�]�{��G�W��^�Q��[f�����s�V�d@�V�q^?��Ϩ�ø���)�Rp������_�;���c�Ԅ��fit��O3#ؽT\���T����=��^�Ie�_�\`fT��e~�b�WOs������\:�wO�#'Ei��>j/m�_%�����ceC���S���X3���ھ[V�g���f/M�H�ه{��,f�Ì��Q�l
�[ 7���K����P�(�w�ٯ_�)���Y|(>�87�Ew���:�a�߲��秨�k�5��]��A��
1�}���U��'���I���	�/�p�3vK;q<0���P�}�����f�К���>�wTv-U�(�'��nG���s�/����t�/c��!Q�
w�_�L�E�yMiQ�'wl�RX��������ڭ��e˷i�����`�y�{���64f��X���'9.������3Vck��Yy��ފQ�a�{����[W�
�lq�@]l�C�M�nP�L���õh�l�$�9Ěw�����ҡu����׷�K��(���V�C+�!�6靺�Vw��k��2�W�_ʧ+�,���{"}��+;R#�itsXvo�9"�������;�n���n-�)�>�P㏏0�7]-��)�6vaz�B�%���4���.։�kH��Ì5P%fj�h�+1�18,�j��`�7D2P�R� |̗�SYD�>�uO��r��V�p��ⷰ�q,Y�7�Rme���3p�D!�=�BA�PK���k��\bFVA�Č��u�w8��:]�e-2��n݌+���J��wm��m;żc����Ib��m�-�5�bU��8�̮�,�v�y��e�6���weҤ��p�ݗ�v����蕝X2�!�4�[�u�@�KQoh�/��Qѵ2�h�X�g�F)*�`I�����t�rబ���h��ݥVnS�X�m�;���H
�kMd�Co���%s�zź�E>���g�F*.��u":�(R_N�0��+�����M$	�]%\H����J���L��/vS/7-�v�r)k�J���,�+���ˎ;���l^N�%ue�-������Δ��]��c�^��]Xd(�K+�>�cXp��YS���U�{�����l3~������y΄�.��0�x���[�lJ�<ȯ-�I݁�
	���pWwT��ZA�*|��*ث�cZ`�s-�E @�|�QS����;<�u�gT'�[l
wNB`��b�ڭ�m�"X�h	Z;h麑��=+.n@L��=<>K�eJ��t��xC��^Xh�lu�s%��ҹ�-�*�EMVZŵN����<�@���L�U����˰w(�V�<�+�g��m��ː5�e�]�:�\v������67��s�=��7,\h�:b��=O��a�����u�;!љ��W^�il1��o]�i�Lj�ĥh��m����l6\X��)\`������;��r�;��\���1��Jܮ+89�����-^��u��B�؏v��-tvؐ�iRTj�ڛ�'Ր�&)�O4nL��IB�w��n
S$���Cm�)���p�h��q�d5&�pw�3����nR��Pd�V��G�Q�[=�p�f�-��Q�z���SBQ���.��>Z*���ⷪ��79p\�#��d�����y9<����u��k��<�D���F�k���3*��6wY��1L�n\�9��.8�+�Ԕ��v�sE���f���C�Cȇ)8/F�3-^wVKK̱�$I`Z����Hͤ�7ݾ�1+*�	6�$ε&�hWkJ낏+MKT��Y��Ay���#R��΍�S�"S�yP<	 ���!� �)J,����Bq2K6"�e�.�*��$&S*��$���B��yݕ��`��aEY�N+*�N�aTYV$rֆl�«��9�QSI"*.Z�eQ�U.EA+�p��e]�ª��ʮr8�q�)8!VeHS���dD$��R&Ȃ��s��\�	Er�7q��g�B��:��A��(H�r̢-H���9�T�!U
 �W*��<R

*9W(K@���MS��"&EW
�p«�^,B�RL"��+��QU\��A���"
Iu�r�L�"M�9Q¨�J�f�wGj,�!$�T���Z��{�Z'���B���ó�D+NBt*��I�I� �� ��55z0C�[X��X)�,hhG��K�������%t{p�f�!j'�f��x.�C���{��>�(r�.�b�f�k��.�?�3�P��R������x����P�x�\sRY��)�NF���~\�nTo�� �������϶��\yz��D>gFF�.9�O���T{���b�1���iwerAӘs�~�═�&H�}2�D�^/�L*���!c!�����>Xv�D�[[��K�ne+�ͳp���٢T�Q���KA-fDmCU-#C��jpe�y�K��w^9��a�wux��E��H߽��y��r�����Ш/��r	h��������5������а�wO��x���U��[ ;��e�*"�2E|�2���c֤��4��DVc��s��myۉ9;���Z;�>%a�����+���q�Isr/���������UfW�GP'G]�m�rr^z9^Ѿ��!Yzdc����,er�p�:������y�Ĝ��������ř	g)]�r!�5��gML>�fއ�ä�w:�f���'VO��T}qq�:���U-�0�	�G�[���K /P�ے�B`J�q_�څ��+tø�����g�����_���+sdz�
^��ݼ����X�WK���M���r�b������j�w�� ��6�8�� ��
�V�w9�ve��nu*�Q'XȈ�����y�wm����W|�CՏ��� Ј�Ŭn&OdN�ZT����vo4�����+{��;����:L��((��qſ�E��7�OƠ7=�Z.<��9q3�t�ó��ꇛ3�~��zb}횣p{�z�'����� z#����zqr<��ݝt-�Eh����ș�Ly�G���j���r�/��J���vt`��)���z�M��g�~��>���"���A-V,V&����EhƯ�s������s^*�&u�^��sޫ��_���?�b�3^�+��[e��0(�pW�������ܠy\}98����g�rgY��gȼ�y݇�:}��y���W���]8��i�ٿYi"��[�u�A��>��nM�SqT��ȁ��L��j�z��>,g�<����'�����xKޕ՘�S�\�G�O{�N�:�U ũ��C�\�(�5��"o
�{�mCDŬx��F�KK=�V���E�u6r>�D�.���������r�/�n@@<���Т� i������7�^f�t�^����j5qԑ�>�<���	�^����s.O���9�yB'.[��=r�����®�D)��a����D<J��{�x����4��e�S��.k��t�~��z����yS�����vM��;��S �5�)	@i�Cu�(�M#����y�uJ��I�S�j��$��l�t8�⦤;�M����v>����� 7W
�t�����.�h6�h�N� *t���e;����|!��T�
�`7w������
�d�=��&b����>��`;;���lz��L\yK����u�9z]��E��w�ֶ���1�̮'���[:ja��x���h���û��ʬ��׊sׅY�d���3oˁ�>����]�Ey�R�g����>��0���t�O��j�8��W��~Wq毧m����]׎C�����C�!ù(����l?��ڇ�>�hG�L�ȧph�'�y�=\�x�3ﳮ>��xty�K#�,N��{n���>@�o�|���c�jF�_��s��w�B��x�az#z�H��ٞ�>m_�=��o�'iO��|���oʎ�N�^��3�"��z�:_O{��́��t�\d֟_�,V��H�M�K�;�*#=Z��NiＱ\V�/<72������^�;X;ƌ{�E{�D�aՕ^_d֖.2g|n5��ʻ�^�"�=����}����8޽��y��r�ӷz7���1��[7�IXO\UC�]1��=�>	��v*x�y���|�LS��5=oR�w���s�3����WhhϽ��}"\�6���`LWz��L���`F��H4#�����d��;��o6_19V�t�E�l�S�b���&�!>��ɘ����R���_�*9&K���4��u���oOk���F6^��"G\ �Ǹl�b���0�[g7��U�� M��\�7Y���Z����]Y��*֭�EQ�D�W�^���]���V���T�z�� �d0�������W�g�=f�:Tv�� }�l�.�&�����=���9����r7���z���r�/#L���-���]�y�"�羊�S�ț�c�������c9��������ڃ��}w�b��W�N0y���R�J�Xr��|��Ы��w���.{�^�]���=ٹò.5���_����G�^؋�LLS������w =P�$|=����۷�{�;$j@V��V���/<���7n4U��L�z�dƯ�bc}5�?1��J߅l{�g=5鿿��B����^6_�vAU�p�����(�|i�u����y>t��5�����8�*�����Lc��sg�r���U��Q&�<����ς�ihB߳���eE�`W���'Y�>�d�.�=k^�Ƕ���/\N�~��ǡܛ+�a^���[�[[�	r?��M3�$��o����������7��3_^�*�ǇG�k���� �=���4�����7(s\.��m�z V���Ӵ2P��6��QbҦtfn+~o�/��y�Y��w4��oN�c.�E-�19��ݏ��7ةp���f�X�eŃ�[�X�y�����J�����1�<�U����;u�moYߴ6��v�N�����sd1Fz�#���k����,\f�i�@�vu�1u[ 
;c'�x14tfe���gu<�^�O�ʘw���Z/�Ew�>ë*�᯲���g��� c���=\�=�'�-�b�{�{�|����~&���=��Ôy������{"g��(z��<���Ȕx{���
�^OO��Q��Tk^�i_w�?.��q�m�]�g)(�{@R���`���?A�lv�T�ڟp�/.:�g�X϶�x�sA��^ӑ�K�h�}��Z��yE���93��#��m�2��9���O������"��ȶsjX���c�J�3�=V����2�:�F���/�]���+Y�\B�EV�R1��K�8���H�D�exW���aS�_
��lt��(±��t>����B=x^􁞇��G�D)���d77�n"�Q��*�[��i{��L���c|��k�^�4=���x�u _�^�\�Q�~�#�n	ah�ϋ���m�f{/d�]�˥��U���GvgG�����}�����@�3�d[�rF��2��L=���c1G�%~�����<F�奯���]O��#{6�ھ�.���J��I�����ҳf:�]R��syQ[Sǈ���͈]l����T�ӗT�]&�Օ�E��,�i:�=Q.VX-pi(8��t�T�v�as�y�ͬ�)��N�j��S���*�J�taத-�(]�"�����9�%�Q�~W~8wլ�N���wTӺ��=J5��i�P��T�c���EI�}7^q�����F��wǰ��X�w	צ�.=�C�r\�l8�0�3M]�������X3ğoJ'�rO�뛨�������3�;�C�'��K�ʥ�S^��<�s-�;�T�#�~�{\���6�e#�r}Kw�V�L<������3_^� m�.|��V�ٞ��gk:��X�uT������ǽ�b��	��BO'����<7�w�ZrG�?!�b�ck=�{���v��Ɗ�k� �k=�d?N��y\j=��C��87�<gN�R_�ᔱx\�r�	�~j���~"|Vu8ѵ��^�UzΆzz�@��W��߶q���޸Hߞ+��v��p���v}�ד<.�ñ������s:3�5�����o�''��ϡs���Wg����oT-@�3X�rG�)�����w��rp���7=���γy3�^O;��O�tc�3�yN��<�rx��w�����G����n7!{l�>�ES7m7L
<�~���mL/\�ō/��=�����CJ�:�rՈo+�"��Պ��;���N�4$R8�� �+\��y�]�ָ�L��v��1��G*=t{G+&\]l�Rt�8�u�Ht�. �@�O�EZ[���a\�����C@��Zo1���.�	k��`,t�WS�ëV���^_�܎^�L���#�����Z������@-��p&��M�^/s�G{4d��W����ޅ�Ѽ�ǰzR8��n�k�4?W�¹U^��������v�v��xe��7����A��e�F�y��\U���s�zB)��7�:*/��E��UzKϴ�����Y����g���n�+>���s q�o��-9�l�o[ȼ�J�F�_�ǽ#K��Y��G}>��=j��j�0�`�l�=�_�\LL'QjȚs�:0�V��X�Kև��J�1�}��3Q����O����S�:Q�Fy�ގ[�o�}%�Ih���>���11MV��}�zc;UY,Zy��>����5�~=^�Vp���P����
������5�k�cB��ǁ_�����O5�ř�1�������U,��@�"�x�x(��1%��;A��v3v���k#ض����rջ�1�f��R�3q�ƛ̿�7w>#!*a#�?m�U�G}�$���,#��u�ϓu��qFؗc}��������o:X����e���׻:�=�}=��ڟ>�?yJ��<F�t��K:���3�g&�u���w����/���,��#Oxa&� vȰ��m!�(֩�E��j���|�#Q�Uv��mF��I
�+:i-Į9�,���s0�����\����g)��Ж#�7N��6�����0��:{��p�ѐ��X�n\�)�l��{����Jd���c�r�<>�d�Zn5��NOKzy���P<�>%���`�og���OԹt츿Q�k�<�Oi�>U1��ZX����\������_�H��Le%�;���u�(���ݹѩ�p�ym�b���l�I�:����c~ɝf�ɟ���g��]T���۸��٦�jW�=�>G}rǪ=��C�}�P뇴)I����z�����2j7��J�;㾅U��'��8����Je-��~.Z�2�{#ޠ)��Y>��ZBx��pFv���'H�����>E��4^��|�M�^����)�����U�YJTY��m�ܩ������J|��>�7n*�:�t�7,y���e�O��M�q�T���Dy]�H��c��`��j��Y��e8�O��K�4pu���N��(�����髆��*�g��ʡ�{Ӏ�ǿ{�z�Q����ލ���1��\D���r����W�����,{.�����E���~�尫kq�aCgf����)������_E��2��^㲩 =��S�T��^2s�J9���^7�3��U�����[��'�Ӎ�Ѩt�)>�]�"
sbX"�ډ�Ͻ؄�ku��>ݔ(JƦ0����;��A�a�4u�b^�E҅�*齛{]{��u�[��z>/i;��n�[�9b��<��v�7����]�{2Ͼ�^7�S^6|�{ �������w�NL�.��m�IT��ޓ�X*�x�
������fғZV�Fҗ�ӱQ�z����:�京�(�^s�^��x��ۨ��ή�y��6}�������;�=,i����S�����J��t������vJy�ֶ�P�h��t�$y�;_����>������f���%~���wb���*2�p�+�2��N�@2Ϣ7��R�Q��y=����v���y��,,٭7�@�\g[�:s�f�(�H�Y[�݋��< f�S�}�|�P������Ew�$������+j竬����i��gh/J;��ԘS�9zHCn1z�M��sǻ~~�ǞZ2<�RrK;�3�M�C���,��x̬ռ�'y��4ϙ���/�wq�z��>�K�}���6�����Ec����|�T����_��n=���}U�L[년�LvL�'�U�����x��>�K�j�\k�q�	��ۗں��5���T#q*@[uL	�*yW>E���,{�ԇ��O�Ѿ�=�xO3P����.L˕�������A�s��¤���)U w/LZk$\���5ƺ�=��ٛ��XX��0�{�zi��}�YC��D[yX�۔�Vћa�t�+	G�*�}�݂T1Χy��i�2�����;ݹQ;EB��t���\�<���q��<r��v��EARْ=�-�N�9��>�b1�g*�I����^G�j�U3>���{�lz@����gN3q��L������*1_�Xp���Պ�U�/I�>�&�y��z6���
��$s��@��������@���.��7���%4M��R�e���we)���x|O#��&4�Wp������� >�&�S�-He񞬰�����VD�k�����:j=�}�D�JV��S;�	xi/
�\?+����}%����:g�Lz���u��uָ=V/�&�0��D�xu稏TE��"����F�coU��p��s��bT��p�o��}ɭ<��,p6:���>%�>E_�7P��[��O�I��s��B�c֝Y>\��9�3�5U�n�wa]Veǳ]	����+���+���B�N����7��fz���g�g<�l��Ӟ�������2|C����{n���pTy	:r�|��N�<7�ꆧ�ĭgB�˾��v�g̤zo:� ��~���<W���^���`��x�L�f����7����_�<���.��cNp����6�Q/�;q�L�c#�����,!][-e�s*4�+��:αjg^�b9��k��V��y��6��� �YP�Mh��'w�����l�N:���NG�%�G�Y���8_|
q��u���]��K�u�&u�QAR��^�c3�:��u��V��ڡV�.��2�mM]%ӱ#=Y�\��iS3��hj���c��!�4޻�3_{/�m*�[8��hg&��eEQ��O6H���E�o:�Zc|�XЫ��H�4,�v�=8|5���v�f��>�Jhc��]�p���'s��w��	�)�ihbS4^�î��g�b_�2�pS���-L���f��R��v�V����i*�WS�!��^�w�Bs�`ƕ�q[;rȕ���hG^7�Q���j�� Ek�����݅F2���퓥M:\�m��[r xt��h�H^k���h��*��hUܛ�k��0슛{[���*��b4Fܘwθ���`��0���/�u:�i�AEt7{^�m�-Ns���5e���^������)���u"ڞ�:.�bB�똎2앹0^3˩�܋g�Gxn�HNA)/��p
 ���b>��Ⲑ	R�}4�ڝ��P����R�9f�\�p���
�!�D��gw����+y[%<�{��Y.^��M}�z:�,�Kw��Q�W���r]q���zn�W4c���ò�m�7XX��i�Z�{�̻�Ԫ*ɣ:�W�xw��O�{9�p�`���Ε����FY��(rj����B�z:w���Xȶ�U%��nL!���^:���*�1��v�^�*�(�P[�FM.CJZ�}�v����Ps�*����6�d�����V�YZ�(���DmB�>ì�(5���hj�����K��>�g�t��da�i�W���G�+��cy�:�#�9\W��Y�v�y�b��E�&�r/X�Z:����:��>�0�����JE7�h��e�a̺�8��]	B��Nb=%��p��5�]t��[��j��y�3�僗���plsF�
 �]lY㉧�B�閵R�����7{�WR����Ap�0�`4j�௣���\�y�K)0��4m�Ȟ�kK���[�	���85�T��M��].jmؼ�ٸ;(��1J���nqX-�Z�0Y?!uȬ�1=zh�#�2�w'���'-��XL���p��WҰ��@|f��w���w/�@���z��(�����4{jZ_ݛ��q���-�o`�#���F^m�{6��W��z9�̓{y����9eA6�δp��h50gh0��t^^Qj[F��)�+z�t�+� L�9�89��ord�}j���;�˥N���P��2�:�e������L�G�tEj*��$�����y�I(�E�Ձ�H�VUTh�s,�"Ћ6Y[!0�E�PE��V�(TD.u���H(.DQQQ�+�D����PW��Ty��EQw*DV%b^y�R��T9�T�yjj�'�Z!�((�A+β���;��^�
�UZ,PJdAr���QW�{�ԉ���tH�+Z"���AW�8G�ED]P�Gq�9r��A�#�V�"5'ZQUqչ��TWrKRj)٠\�*"�Q9����U+s�����:��V�D�DEUUziG(�(�(�B�D9r"9�AEɔDQ˞�Gdv�
�\,����A:�%L�s=@�#�W(�٨��J��B�;���r(�9�{�b�i�^NAxU0�RT���g(�"�$��w8�����"Y��.��wd"ds-3	$�23�(��%$Q^ ��\j��+�ꊹ�O��gW=2�]j���^ގVq���{F�뽮����]��3F^Jp������nfb������bH�ѕ�y)\�F�@����:����7���R)�����&sB<\��ir���r=�*ɳ`�U �&���g}1����is��L��gt�X��w�����ȱ3�5�v�]�6��^��[g�����M�����>�,���}{�ǧ�W�tꙉ�*dK�lG������S�����_��oG����R7&�SqL	�����)��U���Ȼ��u�7�ٻo���l�X=薏g�^�n��c�w��}rf�C�1�"L�(���c�W��m�9�W���*�F���,��~������E}�_��VYe�!���P�ux1�R���]g\��z��z@����{��x��[�ZG#ސ�g#}���n�\{�^��;>�d[��B��Uwͻ�� ���^;>�O����3���*��t�{�I�%��2��L)�Ŏ���~�~ {v� W������D�S��џJӹ ��z���z���������s��u�݃|�_��_�ېj-�zJ'>��뛨}��ci��:φ�|%�{O=j2Ne9�}B�pӏ\����j��u{Vm��{3���Wrk�-��F���̾��!Ȕm=�Ϋz2�lk/�c%��uGӷ�z�Y;:�H˃��:�t�[c��*��(�l�׃h �U ��S�c[%���Z��v��!̂�E�0%���Ι��2cJ�<p2�S���VU��C��V��:�rpW�=� W�~���|���C���0�3��T8�8��ؚ�}�����=^�CCt'�Z���y�A̋�Đ�Ĕr��c���~&߯�����<ĉ��ϗT��w��q�/�������y��uRȿu1<n=�������y	(��_F)�.s��N:^nG��>�\��S��rr{K霒�nr�Ǽ��Q�'�����#/���kjmz��O9��a���?�ϗ.?��}i��V��Y�ﳥ���@��u��'��[�w~v��[��t_$�>�9b���G�y����O��b�&��y3�7�v����_o������/��sR���@�$������]p}�Q�{��9���z��*�7��s�8yݭ�3�#��sڮ|�_�;������s�3����:�]��r=���NnM�Rfl��#������^����ߣL�+6�7��뇓�����I}=��a�����_� K�B���7W�Vn�9�Q��}p	���E�x��&��q	�\{>G��Ϸ�<{�F�_�U��5o�m��3���`&89�D��z�!v�2Q{��]����r�!��v�r(:�X��G��_x��}$9�|-���7�h��*��[a-t��K32���w�g/�A�x 3�!�e��#�oe���	{(�)�KP�X���N��rrV"�|������Ԭ_�9�2���b�G���߲X�;���v�AdC�6b��
�&O����W�R�e|��ǣ���ɉh��`��eI�W��^6�|D<V�{��&<j���v/���s��8=����>�H�=�U�f�xA�<`��H��}^ӐKGw��^��=[����i�9ST}R�Lz��{n�S�-�����	��lzU�7=.����]�;��E�ݐ&LO�?*�>t� ��������~�D��>�w.�..:�����V�ڌ��4w�Q���������6����i{+G�� �9�=q�nI����}�5VWw�Zԡ.Q�&s�e���q�Z�N��l��eqcܞfG�z�����⧍�w��ּ]��ǏM�_�=7(�_���$y�����y;�ד����_���i�)_�</�B0���x/�γ_RI*�B�s�z���8a��ؒ�ۉڇ��W��f�i�� o��Q��s�.�:��Y���HsX@�G��h��:��-
��|�Wq#�quT<5�׻���&�00�7J,��Z��j��;_KWt,s�Kb�+w*�S�r�N����k�SvKݠ~�dE�d�71�ox�M��R�f��љ�����g��t�=��z��d��;7�g6d�h-�*���I��D�Y���`盟����z�*�xv��x��Nx����W�y�p��޶3��,i<,����h=9#�և�GWq�U�ɝsq��L�D�ƽ~�{����e�q��w�<��**�+�/�4Ȗ�|���/�l0U�0/�G�&S�����o�Uagù[���V������͵�ZB��M��v��n�g��
f�z@[qL	���E\��FԱ����쀧����߷��o^�]�J�DD�x��q��_�=�#�Y�ϵ�;7T��d�d�exW���aW�mL�)��O�O)�Cv��������?E6W��W��l�/}d77�n�Q��*ϋ��X��8b�X�h�s������U���4-ש#�{�H��E��H��ơ`#�@Y�"v�L]��[���]��z��3�c�5�i\Q}^�Q�\
��z ���_[�rFsN�?O�{���勏����j��S�v��=2�����g���x�N*�Z�޾q��������V/�n��qa����1מ�=ei���|z��\;�N�71�Ϻ��?kY6۱����M���f�"'R#*m����N��u�z��+L�nJ��ywhvh���ы��ȶY�}S�{;myQV���J�%_,�o�*t�ŋq�S�ɧ��j��r���ۘ�dDj�X��a�����&[�%˾\��\�ri�h���Q���u��`��@�w���Ĵ�7C�$�Y=��I�=M�5q��^���A���ǻ-s�L^O�kW�։�a6=��ǜ�s~sC��H#=�Oa�+��N�/d�}�^�/<c�hN�f�;�ҒC��� =w���:�d_�������P��87�!'��p�ó����םB�ܭ+�lJĤk\��Gz3j��H��g[ VjǀdC�V5%�`qZ��\?h�y'���=Y�w3;�)$=9�"t�%����Z���3��O�v�W��Guǽp��<W��]�� yy~�^�c���v��998]S�ɭ.�g}1}΄��E��l�_Ze��p�멪��sj�W(�4|����%YD�M�\U0&�X�u�'�[��vj�8��]2��w��x��Tpys�3��qsJ�6#��>0��L�H�ت`Q�@ȿJe�_��>�g_��V{WO�����B�O{ף"=�������U�F�z�p��=SPO ��P�W��=�Ew�N��{����}��}�Q[�Q�j{�=���A|w��EG�~�S�Yznno��2R��|\����Y��!�h�yDoc�O�v'pN����]�Sg��p��<m�WR򍬜��N�����å�<A��{��]�Tz<�����c�, ���:��Iv+�Ϛ��s$����(Ĉ�=-n��]�t��5Qof�r���Vo-��� =�z �S��nF�4j!�Wn����meǠ��w��Ho��9�A�Y��ו]����~�L��o�0[;qJ�Qs�sai�/�CĮ*�u����w�D��Qq؏u���(���_V�P�����{�Y~�r@�PZ<`���"i����Ҵ�|Iz���=�Ց�����i{�f={��gc�8�2��N������n���W������q�ù�ɽ�w֗��]��7��d�^�׈��D��=@����(��#��m-lW)�K��?K�6������?Q���i��g�x �9������wc|w���"�ܔp�;č��^6'�w�cZ,�qc/����7��כ^���3׷��̿9�d(�S��ʨ�@yG	1�<rc7v,�{my��O�a�졘�����ic�3���}��߼gYD��k��X���c;�.�\�v8�.�8g��I�1~\2R��r��ҭ~x�������\�{};��"&*}��M�oJ�n�Ѫ���b���v��x'���a՟U1��ZX���dc(�W>���6@
�S}O�^���Ι�p~���)[�{:
�D��ۻ�Q�c�=DKr��	�F�5�b�Ho�nP����cޫΩ�+�:�[*���w�ۢ�V�En�7���R�KW;M��
�O	��C{��ҡ��B��vqM,]�{�o}��ms${υy�ѽ�����(�)��I�'�*���b�bnTv�s{A}�ދ��n�ӧ�2�����ޯi��י�\�k��{�)�����a)�����bk�[�Z�G켸��>e�mT/�}p�8����Je-�{ ��K��^�ћS�q~��Ԭo,��<
2}E�1M�
���Wl�H��y\z<R+����ol1s[`yl���{���=���U}zd����}U#�.�&�X�;���E?���b�϶�ˊ�r��Wj�T"�q�ܤi��n��x�zK1-��0P{uJ��Y��x�l�%W��˫:}6�c�k}�U�����3ޔ\�g�iW�.�K5�b|�ȉ���t���}^����X<�����U���Gw�t:�z�>�U~#�,��@y�#m׍�E��2�f,�ɿ|�nq͜��`�z-�Tt6wxL{v��ϗ�_�A���
�S�XG����[�����Ox�2���<�6�;ћD:�[&��O��R���بۆ�sf��t��uX<��r�[�1��r"�s���q�ʉ.�Y�
Fɸ�'$�tX���:�>�7ne����FLP�Y������Qη�4�h���e�m���c�T�nRG��5��4�k`�ϒ�/j<��n��[6u����Y���&�=���P`y~����8s���C�����8��=P�fG�wg�"3a��*kԫ+R�c��nUEz<����YxzO�۝��;�ד��޹��^�F���eV��p��8�qUv�V�Ǣ;�}�3ʎ�m�
o(�h	�7Z:kב�o�=g��XU�-�;Na���k;/�*�V���~ \?m&NC��J�C�{���!��r}�,�����B\H?v�(��ܝ{�:x�;ѝ^�z�w]�^��7���A_�yhp���H[ݢ�D�Ά���h�f�_�}��nd`�c��q�;���&O:��k��>�K�}�u�I�^xUɎ�ڏG�0�����]��Q��=�w�f��|}}�y2������zsޗ�ћ���|ì^��m\)]�T=�}�{q��E�^���� -����SȊ��"�ͩc�^�=Ccr::�U��M���5��{���j=m�)���\*���-q.� r�����&��E;�֪�{=�Kw��_;�B��팎�JG�}@m{��QϕxT;�!��'�=�Rc~�ḙ�'E��O��(��y�+�/z�W�.ho{9�P���{�,�uc��6Uic�"�C�fYJBǕ��W{�gތ6�ʒ�$��%]����w]$ʱs���5���F��0�4�Y�Tug������9�t�s.���y�`�jv�
�jf���Y�Zg��\���L���w���n�I�{�������^����<yO���f*�Ͻ��T.b����f�`���㪞�'�2���K�qW���x���\
�� F{,�o���9\*��ڷ�G�B/����RG}N{N���ӑ�)/�(���L�Ku�};�G]ﮗ��Q��w�m�W�IG �4xԱ۞�=ei��F���X�T*��T����&���sG\������9����5s�V���z�n������l�g�`Y误��������mY,\k����A������ ��C�Z�+�>Zد$��f�����?�9yn]s��3���3_^߀���2<ꥑq�'��7�Eh���;���u��/]�o�U���/O�]B�ͪӡ���g[ Tb�`Z~�e����~��������������~Y��hۉ��59:+뜨낺�t��.s�J�l�������C�
�}v�_��Ӯ��[����F�=�;�NN�T��2kK�w��w�����v�x��-1�*eܫ�#�����'�[ŀ���m�њ�j����m�6�Ჴ(s�hԭ`����)0O�	�`�Ґ���<u���M̰�ܨVr;�������gU�5���}�w���v�%m����f�z�R�e�[[s��n�{�1s�����)[���(�?��{��[���V�=�%������Sb�X���p�"�{��JΟ'6�N����]c��+Е&xdyϙ�\�=�������{���);T��ȁ^�jA����]���s}�&ݬ���B��;=^��|y��f�%����j�uv����~�  _z���W��zsCc��(�}o�����mCF���dz��>��W�và0L?_��7%Hd��6��_�w�TS�`{fAS��-n}�x��\:��r#ސ�g7�::{���=5�:|2���*�,��=�I/��POr� ��T��!t|j��qx���<J�;Y�>1]�.��?ۛ�P}D���;�ߪH��S��(-����ꏮ�3�tg�Ҵ������T��ܣյ��_�/GUu������
��5���#�����ϔu��J���>��Ͳ:���gs��]���k�w�D�s�׍�~�]9s�z=U dC�L��\�B�����ܩ���ʍ���{��RkK�꿚����:�g�r�9�~>/Q�$pO�R�]��y����Fv�7��s��J��jr6�J�!�z�{�_A�j�r"���z��uch[h�,�qC��6�]����1V1�oS,fK��[��F_�����º�Qy�����i�;�����:,anW4��V*f+��1LR[H<��nջ�`����n��ڙKQ��'@(HE�wLw	�o;	�5�C��8�oɜ��f�� ��d��Z�͹JblM���V�^FJu�-�9��Ɨj���>F�֋
V���czU�x�[�mk�:dH|E�9k��Iëq]������+W�y_<�.��f�0]1��Y�2�*)Ф2����J��)n�5I�����Q"�	:(�����EY�_9�eXX�.���*\q���*��Bե��k|ԉ뱘���ېќ7�fi�P�+o*�ΰ�Z�EҨiTXOjtgc:�ʚ썬�MC�z�b�E�Ս���Ǣ�ɪ��׬�֊��i5�V���i�4J�#ɶ����@B���'i���;6�<%�������;����n:噘��UkC�Ę�Қ�Vk�]E�8wZ�s��~�͔�NŕV�D�&��׻V�P�:��㎝�y.\�����3C�'!qu�s�o[}N�����w]���=n���#�uݍ,�.[ilƴ��]B܉f�n�0��CL�Y��f�daWy��(<5ƕ�v��{oa�
��98�Co���꽴�*�	��'';I��,��g{�kw���VQ�N v��V�\H�V��zJ��t"ʺ�������F;;J�]ê�\�x�j��X&�>��[9z2��G�t۰qǝi%Iͫ�,��hWA����(v��G�^���ދ��:��q���Y�1��T�Њ>"uf���N8rgm�g,���컗����z��]���&�Ժ���|��n}y�]�����|s7�w͡Q>|\�&.�5ڽ�Q�8�7{�D�`E�C�������X��ނӽ��G�;�V�z|�Jh���v��N
�nr����kS:�
���@q9��x�\'b�sy&�Ԗ9z������1��,�zw[q�VX����%{)j��:��b�}W�3�M*T�c<�ܭ˹�%ʺ�D �2�+���ht���.����y;���̢l8n�IF̭*,.����� �fĖPK�A����%�][�p�Wn<W�;��(��w[Vf��nQ�ï�U�l�B��]v����ʺ3� +H"��6kI�1]�Q�2�>ݾ�0�o���[C��k_d�l���CO	v&�7��g.�����G:R�3TS���,��w5����U�Na���s9��)�F�-�ʱ�N�k��-�ԣѠ��C�1�1έ]�C�`s����w�乪s#q��N����p�e���x�Wq�;���]�8tG]p-
��=Hc}o����^S��_
��.��)Ձ���Q��*�n�6��廓7Ow\�I(_r�G�뿕�&P%�0���S�]J��Dt��
�5=\�G:\�;��T�r(���Ui!D��(�\�K*�*���p�K�bQz��3YUNI����'+�<��I�d���Ù�p��S����Q�.\���HPE����=�ȮTEh��TT!	Q�z��pT�$���5*�3$�K�!�E��E:`��n��ITD�*���Dʹd�f���&-g�����E8���<�#T�N:X\'�'2sN�\�A�Ң��Zp��TK�DU�=kI.�E$*"��U]��Μ.���;��aB������NyN���9I�r�Q��="JI.RZAU*ˤ㩰��ӑ��TC�Q���I�n{����y%;�(s
��ηYHT�k*s��KJ�l�G�dU�
���$Pͤjw�78�,�����'�Kz����(�1���-�[�zS�c8QP���GMtK{-���\���Ex��ټ��>���������{\�}���&j�����^�xl?U��g��w����9k��e[Qc�=�$��(-7;,e�p:����Ƕf��/�����Z�$p#�^��P���ƫԧ�uI��ko*+�/m�7rON��Js��\FMiW��Zn5��Nq`n\7[�@�ɺ�{����.\�{��^��;��r7�Tu�.<��I��*��ɭ,^L�����g|��u�U~ף��}���${\����F����C��l�tSd��{~�����,���+�ս���/{�=3�n;j��gS�mz��=μ�l{=`uǽ�����\=�JFǮ�h��j�~����+G�UO���i��xex�ڨ^7Ϯqu�9���[�iS
������͞��~�:¥h��J��A�ِ�Ȋn�Y�W}�Aq���Y�ٽ��.�z��U��{��{8�9�{(znků��PT��d�dK���ǙŲ§��S����\�X
�+��+�zr}Xc���L�o�i��[�y��,i��F
n*�%x�9���UӚp��y$z��z� ٿ�����H�9�Μ6�Y,�;��S�	���rS7�WՊj�K�ˇoQ�{=���ėjv�QQ�ur,��o�}����짼ԕ��ë
�B���t4jJ�C�,�kQux����qu��y]�7��ǜ��s88��q��~��օ_ޥkō��(����� ����P���3�<ۤL=��`r�\GݯL�W9���y���nR>Ԫ�G�X)|�z��nAn�n�h������~�����ebKRZk�v�^��Jv��L�g�a���^���p����g 
��`/Ma��"c�몺w��~�'�<Y�vl���['4�>���:a�\ٿ��@yV::h�7u1Y���>� ���I���Ľ�i4|:�p;��}�ƙ�ŏt'����*c�IYW۝����)_{Lz#5EO�۸�9�߉e�Q'���ׇ�;���N��z��2;��j9�b�^�,���nS��Y��o��P:=�t�ܫp�����n"KE�{^F���ֆw���0�s�Z��/�M���.�5gW��U~ \'����e�B��+E�碻�D�a�8�IT�%m�mP^MO��Q�]z�\F*�7���WCò4�_���Nx���hu����-��];���5�ֺr��4o�80�d �>�w��g}7}3s��7>k��9{�����\wp�A�}�D�Tl��d��yVtd��Iv�Q�<-����9��E'_>h�|6b�M����-�������Ż�]t��ټ��J��^��<b�\붴s�k��t;��#T��궲�G�X�\�Z2���-�7�abȥ���Δ��|���H��U�)�!w����E��@^��u/sJ���ʧ֖��Y��w�8�,a[�ϫ6�Z����d�Cs�n"R���Yy��(��b*�<���"�ͩc�g.���>Uٯ�6�e_�_�O3�#}��ޟq�u~��#�Y�ȍqN͕ -���z�e��	�w��0��RVv�Tu5\�R���w��F�{/�fc�0Ķn	p���;-{��Ы���-RÄ�/6a�u�h7^��}�u ^o�~�r.=��t�JN����ݳ�y��T�	�l�ϊ��9�a��M��ϝ+��\}�M��\�G��D��|����(�=���>�s�Z�3�s�w~;�#�^�K£���Ƽ���:�7�J��-V��ܝ��9<�=���J��0�뛦:��G��i�Z��;c:yT������}��p�/}�j�c#��	鿙p=C��$��]��O�F����|:K7��V��(ݿw�W-C����a�{�d�_�t]��΄�ߜ���wDQ�{	�lN�/aQ�®@�����@��sd2�����wu��06.d�J�,Na_���Y��[n�����V�YN�Rd���]�{>I��s�u���� G2���z�T=gWSH���T��IӪ�>��,r�ÝI5՗���U����5á�׭ˏ�U�c��t#���K'�R]r�1ތ�\o�θ��� %+��g�UO��*tyC�]�	��	�{�v�bc�`�>�Ul�:���飥Lu�}��=q�U���Ǧ�3��1S�5?V���A��
)^�z���z;��W��RU�X�ݢ�dD�����2�+n�O���`o��ү@���>�l��X��꺞N��j����_\_��o��{'N	T�X;)���>�K?*��C�����y�cwR�v�A�ޡ�����W��rS=���>���w�QEC��[998\U0&�X���B�-��%�M��͎����|�ߧ���B*���|���}��n��c���ƺW��g��<�S~	�g�l����f��������VF�Bw��|XϏ?^���KG�ޯ��]��B�����:̕Kٹ��w�~�=oe�q���Q�&+��8��Pѧ��g������^o�Z4T{���Ǖ�����~���뭽C|�_�9��!�l�ٺ2$�\�Gض��_<J�׭#��HE2zʽk��3x����X�!�޷r-���^�e)���T>F�0����\S�5n���үh�ӷ~Ĭ�腩[��ڬˎ�<��q��[��V��	� IJ�A۲o;8S�ÙK[�2v�R4�mwkU�;�²bgvp,�]�X���U�%a�+�}]��VaZQrffgØ�eݦ�s@���,��S����P�xX�-�Y��s��f)�u��g|K9�����F�`�uNH
G{鉅�L��8JӨj
gS�1+p�t���x-;�d&v\�W-���8����ź�(�����S�+���Yr�0�}k�E����t|��݂X��VO�~��G·�r\����+�7>Gi��?W�WR~�X�e7�-z7�KL;�t������Â�b�?U2�ȿAX(�*x���]���5r��5ȁ�'=({A���ݨw��7��3_^�?������EǺ��#f�Ƀ��X���v�a^.P:}��G����\L�-7;,eǧ���ic��?)���O��_���c���52}��r}u^vQ>�)�ѫ�6߶Λ�Oi��Jq��\d֕q��Zo�r7ӫ��3�C�U{����� ?gv@�U��>s�'�q�5�Ȃ�y^F&�>U��[T�Xa����Țwq~�5y���m�x��P����W�/�;�+��������0�!M��9��o~Yw�wu���R��<}�e��&u%��vc��~��^g��^n��ў��Al+���|}b�w�oq�^�cWx�`�F��Uʞ.�{|خ��ʔ��e�^�a<Z��K�0RO���ikDtAЍ&���U:���R�x��"��d�ξ]K߬���_���͛�����$��y�e���<:v���`
���a��ý{�?��:���T�ҿX)�����&�'"'��O�e���Ttz2H�(����yo ��+�ʭ��� ��+@�R��
��(?��=-1�e/y\{>G���>���y^f�}�w��+����Qs��O��k����e?�����m�H�K����X�;�,,�b��M�5��΍�%��U��lǊ�i��e߳�`\�>�LKF��a쪑�J�XF����;k|s��g^%*�{���qн�V�\:��C��Eˈ�H�3ِE�f�w�1>e0��:V ��2f����¯"b�������~��H�gޥWㇽ��{=X�����s�P+oz��ꚯnEu~�}��F�V����G= {�}hLS��;��=�a���>��W�΀�au�c��A��s�ڙ�W�=Jz���M$���Q�y(�|����ؾJ�iSG>t&2��͕�ʉ>cՏk';��OA��}U��{+I�|\��ςF���^mhw�N��l�&M|�X��fNw@�=��*�l��WS6��~�ު>��|⧏��Q�(���YxT�3�;^�g���'P�̉��3-��o�
�ҏX	l�/�lA�}���-\+qe��3�a�]fc�����v윁�)��e���p��1����fB,�l�q�,jc�k
���I�b}�AI��qm�Z�DU��s��q+�^[�:>Gn�{m���̓�*sC�gѝh
��=�ᾜw��Q���X����� �S�\Rs\�k|/R���Ib���w���_b�d����D�y�
��-
����Eww�$\/N����6�2v�Q�k+j=q��� c殇�f�_�^���N�y;C���X���f�y_gW�X��72K:M�;2~�Wp�2g}8=2�y�Ƶ����~/�F{�MmKX1����woT�#���,W�"�(���3��%������zUZ]�S�K|o��V�z+������ݿ@�^=��i�)�����7�F�TY��)�� -�o�/���E���l���'?��L�7ʥ����������#b�zwK�q�����Ր��1��]���G�ٮ&C�S>]&0{۫q\�B��'�u��^
�y��B���2;�)Ϸ��{��S�7#L���~�ҙ�������[�q���U�b��SÐO��f�5P��f�C�Sg#ޔ�����v�B�Ks�~>�ڮqږ
��4���@xk榅��8KGw L?�Ҹ�����+�L��/v{S�U�4ۘ�p��T�{/��u���{�4�&m�i��H��/r�Z쓋Y"��u�Uyk��d�u	.�ķ�������)kU�1��0p��u����mNC�d�J�7Y�Gp��V>U'-��[��ߥv�?�5$pu�:�1,`�r�"��NH�!����$dS�Ӱ�a�%�K�n=q7����/'mG����N����ɿ��Q�e�Qn��Y�3��c��G��i�Z�|z}�$��u�ל�K����#z�G\/W��/�t<�"\�_��j#�|JӒ|�\M�5en�T.y�۞=���oX[ݞB���Rn:��Bud�Znϲ2=΂R�dO>�� z��<"����h�I���s�3�g�zد���9�f�m�)+��g�T�/�NO_��b�Ǟ��k $��+*�����-Hヿf?��{\�����{�=�L4�X��ӌ��� �#g��d����o{���*��䷯�=��ng���c2v�_������M�S�z�~'��Y���{~����5ůҧ?z���w	����Ȁ��E�,V!����5���e����<���43G��l�O��?@��`�L�;q�����=���5�Q-������7=�!�b�΀~������[��q�)�e�Pht��F}μ�z��\�Tg�Qf;�nM����܇��u�OW��+%3Ok�{KJ�\� m��&����[Am�D(�fb��ֲ9 �uq�-��OH�彾ǹؽ�ݏ^h�Ef�u:�ӕb�5�u6�KU>��H��(k��V�ɝ�P^1Nb`MB�>�Ϋwo1y�/ym�r�ʵo���n
�����r��~���*/���mL/\�Ō��ף{�-qU��Jt/V�d:NvC��vyF	^������|u��z׽H��+��G�PѨy��|�����ڷ��I��\��s-����u_�WL�_��!��'�{2��U��zZ>܅���J��׭#T���׽W>��xSuW��w�r�����ȏL�K�2D@l䩐�pNf���5�Ƕ�(f����l+�͔f��^��h����}�H��=�E[�r@���֨���=�V�޶�w�*m��Yفwg�
�@:2��?cؙU鋃�O�9��p~���5�(����S�h�I�3o�}^�×���{I�}o�Q�^����4K	�k��:�,��?	@���>�`Z��r��I�DM�yd�}��MDi��U�5~.!;�~j���<����l�t<ݺ������>�j����Y�|;4͏x�n�;ͯq�/����~7�_���dw��E�\˽�R���H�}�w {(�!%����vX���ODi~=&�Ζ�����Ԭ�݇��}��WǗ�~��5Ђ��D�FxKۺ>�\Z�K�(no���O����O��Z=8%����.9{Fy���
GT
b�/����C"ˢ�Pf����#i�ʹuvZ!%K�u���H��A̅��䳍j���޿E�����[��~���yQ��I;�O�;,]��]>�/V�Lz~^�0m��C��t��+�|�j� U��t�4�X�*����z+��aՑT�XV���J�w�����yFϔ��&|��5�5t=���$_�ב��W��{1��V��E6w�;b6��nۮ��gl=�o�U�J�;�q�>	��ᅱ���9�}��:�]���ֹ�2&�(y����h֨p���J�)�6�����1]�xe�ax��}p�����s})��Y��c=�'lwm�u\�<=�{~�9�,�D{�;�(�qE�?Sw�yd�\n��#ѽX�:�ّ�3�<r}V}����Z}4��zr�>�@l�*@[2G�%�D�d��w;L��p���5�K�����{բ�t��q�����5�w�=5�X�ىl�<�U**���(�����u*�����$s⑿F�
��*ỵ����}9�l΍N�دS7����o#��~��f��:^��*ɉ� ���D	�)Wqc!��6~���|�������?�cm��`1���0`1���q��6�0���c�m��0���8�co�1���`1���1��6��1��`�co��ckcm���`1���1��P�co�1����6��1�� ��zc��(+$�k?�6�iϻ�B ��������?�x|���V��@RU�����
�*I$*R��B�J �%)	" ����$��TQQ� b�U�Z�*JR��QRT(��EUEB�R�ER��R�TR@�	J�B��U4e���D=.F��JUM�$�fH�@*֩JB���Ģdd���"�K��(�HIU	U {�D�  �Ͷ�-��QBS06R�CSm [Q���*4V(-�MFe*Rjդ5tt��R��P��  WP -3@�` )��
)a۔��R�@��)E Q@�ܭ���Q@s���QJ�8�P4(-��4�)4�I6ȩD�G   ���֩c��(���� �)�R��� �SN�@tinq �pH�룠ֶ��v��!E-eE5�   ]��:�b�����5��A�D�����E�3����t
�V,r�ZQ�7-m����AEtf�"�T*�
�Tp  ����%*����U�V+��
�횹���
�V�t�f��v���;�!(�Zn���[[6�Ws]�)17A�e,�5F�(�DF�%8  .:v`5w�)l�m��:�m;�"픵�ݸ�%V����Fl�lb��F#MV���66�h�-�
F�T@�A� 3�UP�F����,����ll$-�����Tҳj���LѕMR֭��h�UVM��Z�h�F�٬��$ʊ�	$RJ  	���F5�����1�f���e�4[5f���0a����&�U��Kh�V�����P�V-Z�b����kT��P�p  �t�l����
VkhJ�i�)SCSU�mmlR�jUk�kB��`Р��JK
�U
��RTPm�2T	U+� ��������j��S hfQ���H�
�`�Z��� k�� E "� �  �~�e)RP&F  � 120 O�bJR��FL&��@h�� b�{ё���OP�      O��R��0     $CH	�=	�4��$d=f��� �IF��0ddm	�2	��������_r�3�F�6�_j�ųU�V��Ʊ�i*�l��TA������QPy��@h�
�j���o�����C��T�e�><8j}���������7�3�'��@Y!"�W4ʖ���y (�?�;��CDDL�"������1��q44�E�a����9��-�l�����m�m�m��l����m��m��m��6�m��m0�m��m��~y�k� � �I��@l�a mЀm	!�$�� mQD�EqV��"�"  b "����"��@6�!��� m�l$���Cl 6��@�6��!6��M��m � m��i$�HI� 6����I&�m��I6��l	6�$ ��@�H�6�@�BCl�@h m �m� 6��l@����$�BM�$�BM�I6� �M�H@	��Ch
b("�b." �H��H���m�����m@ �Qq\AWU���a	��6�'Lm�M��qEW1�Uq	XCh6�� �mCl  @��H�	:`���
��!��A���6�@� i	;@�$6��"���8��b
�6�m!!���mCL1  �J�!�DER𯪾��ɲH޶[m��6�m��m�m��a��m����m�m��m�m�m�ۦ�m��m�M��m��m��m��m�m����m��o[m��6�m��m�m��m���m��t�m��m�����m��kꪴ\(�_f쮗�ezbR�b
���X��F�(���!3.�e�a�'˝�ei2�\	�DF�np���S7T?�JV��r$�,��WuB�[�6Y4�3�mY���Gz� ֢�&^��Kڀ��E�eK�{	���Ԇ���u2X�&�5�j�"��1[vwe�2j��Tpӽ�nfX�!hѧe3IJ�ZT�Xٴs	@l�
J�f�Ǣݹ��ڵ
l�nӸ�Q�@�	] �f�������8���M�i*n�z�b;��΍�9��NB!���Kٴl6�yV/L��2��fV+aPj#�'�=X����yE%DG	53[U���M�;�ob�\$"E1ve�0j(N2��skl��E8��B�e+�乭�G5�ٕq6mfމ'{{��R��.�u��HZ��E&�{�A��Ͳ��Q̣�^Ǣ�8�9W�I��dN��ݚ���<5t(0�k�1�"�S17Y������E��4�٧ ���P�/tӲ�f(DL��[9�-6�5��80Hdݥz��׿f�X��"�ܤ1�5I�T�f�UC��Z?c����EB�yt���q�4�Ypʿ�0D@"ˣb��u��@��I ��YÊ�n� DV�)�9i�D����$��j-ʹ֎)� B��%��+(n���ݒ��XT���ֽ
����.��UeY��mß���~�lҫ�1�cEHɛ�����=j�f��7%�5�gdm� �KDp �Ɩ��V�Te���Z&�͚T�9�	��m��[�\��*Y6V�0�f��k�:.+~���	n�u"��̶�X���z�uAW�j�t��tr1��Y��A!�aq���M�^����t@��5���O���̈kI�����1`��S�RFD��%�ƭ��U�2�]�0��.�CO)3Y��#K�Y�����H�͗!�Z�4+v,��6��V���cO2�r�N6HW(b�+�F���A�i�Å�U��b�V�U��-�큖�+^�JTb=�����6Աm�Yy��4�`��s	�.1.X� �Dn��?��V0�VU��.�D�fZƑ�v�������r��d���[�jJ�K*n�YGX�ST�*�40j����MC� r��em:�e�7+o-�x��qۚ-DW{��4K4D6���O�����	5c�zG��
��!�%��
`�F �ݻ�f��u��BJ�F�U�DX�n�WYD�����W6��1�p��<�L��n�%��*;xN�u$ypQ�xo.V�j%�ox�M�ۧu6%J۸�u�Di`h�A�Q�u#��2l��-�V|A8Ȩ���owh�H�u!y�l�jjj1�tƖ*�tJ���0�["[b����f�wZ��I7,�Xrg�-�{eT��A *��`�r]%��_ŘdܱS�ج�,#��nKӉSn��YP�X���K)� Z]���ӽ��Y`^EW���k�f=#,�[���U�|�*I=+ ���2��J91V��*��sYО%[hқX�W{�t����Zڋj*=���"Ud�tV&�J�Å[v�CUrMZ�f��.����
T{�2n��)O�m��h�q�L�n^����"�[x�hٮ]XPec[�#�DhV���g׆�cԲu���m��J�k�ޛ�iEM�;�G��V�n�YR��.@�
c(�R�,
_76�Z��͵!��d�r
+&�mդ�̖�f�t^�����U�rL��a�J�jV=�Qs�&"`���b�Fn͙�dC+��R���G�k.���16��ש�9��]Ћ�/m@�;[0�37��LR�{�m8�D�F�a*�JRn���f�6��a�Aѭ��u���-�d��3���QmV�"GoKy!ӷ�`b����Df9�0lI��& y��U���<����BB)0�:���U�)ͨ�6�Vӻ�f��U��jy�������{t��OUjS#��MX��Ȗ�٧3(f��6&RL7[�y�5oF�W[�;Z�5CR M�6m��=CFc�Km���\��̏1J�e�3�������B�-yt§[�-Ԗ�;� Y�z����Y���5���d�Є���h�ƺR�*��%���{72�KnƉ�%Ư�V�BS�Nc��v\�6�y�Y�"�XS��ȀLj��Mʅ�77nT�zP���G�H�����l�,Ռ[�)���Kv��jQ�"#2;:	n�,�iSQYÚB��&)����ii���M
ʹ1_�ͺ!M�j������-e Ⱥw�a��J�*�'(�X��t4Iͼ�9��[a+�����6I�6c���\�"ywi��֯)i��f	�6š5Tcik:T���nSC3��.ﶃ�q�L�bU����V`��@���(��Á��@���1HՔ���Y��j\�M��*em��w���n�ଦ�P�8~���{V�)Q����,���6�-e�Cc��e��#E�SA�h9�����n�j�TV�<�j3���Y�p�9����Sd��(�eKY�<��>f\��
��2z�6����7���h1B���f�y���l���ٖ��v�ީr�V�5c�E-0a�H �X_p�� |�]�`����:z��B�Fں�q�ح�A�Anl۵���f���ղ՚���T�+Ȣ�I�e�s��m���hD�Nr��p�Ǵ��I�4%����/&��
��U��aJPy�	�d�V�jT�t�웻�]��=Mb&�]��t�ݬT��y�wa�U�
@;L��eml���H��ٶ�/Rśz��(H͸uv�]^\�S/Jtc�؞�t��
�k���u֩x�]�֬�t�[���U3�̚f��6�*ܷ
n�bօ��S�,d�5��S3M�N�ڕ�pf�-N�)>�Ե\wFǶt!�VBɳ�ѹ/A�%��WEhFvB�D.T��I4�9M��O^޳$e�������QH�~�hk96,d����cᆅ5SC�Z��2k��k��pIgf&4�hXt�P�Q(��զ#J�s%�۳�Y6����b��^%�u,�Y)x2��@�B��;��d82f����E�C)�V�Mb!RJ�hE�Zy��aq�����A�/`��me7KF](�e�!�ՖD���T��S
����Xb}�D���v[y1���W-�}j��S娰��4�ZѡR�OE]�̋��5��l��8�A�j1gi����d��¯( �:Ƕ�̔+*�3�[.��b��[hdJ�xFlz,9�YV1QX�-&�L�j؃�!��MI��T�e��Y�#
��bcLLt�(^�(�fט�<*ˣ&�2�W� R(�j��w��t@҃
ǫ#�ʴ.b��c
�-���e�pN��º�����e*-d{����l:��n�LO){��$��LX�v��{VZ��c�Y�5��f=��o�dT�lDj���S��E���p	nCTr8�ܩPD7`�Y�%�
��s�k]c�l�#��m�����(f"��-��L��Q=�\�u�
�X��2Sp�	�T�^��[2���+u���ݖ�la�Ԝ)}*ʭX`��i���@5kI���D��p�r�Vnk��	�Kqbvo����9��/n�E�up'M,����)&���IkVmm���C�μ�� Z/��/S&UKY���5�X���c��*�īOr��M�6ķb��N̰�`��awp�	CV��Pj�i��lM:.*���ܛ
a���.�ʴ�ʵk$��T�y54�b"
�!��Q^fn-�ȶ��2��3�wķ`Ʊ��2�@؇�+axCʂ�J���أlԀ��I��l����8��Ө��'� Z���ٛ�%�aK'd ��o]GL�X�V���S�l�2�-���d؞��X٭�/k\0I��4�Q7-���bՅ��o�"ʬ��m*��k7����@�e�osVҩ40�TRRl�Ő;��ଆ�/%�aԍ6� �.��j�&�e�����(���J	w6Dj��XH���Wq<
�Ƌ�$׊@Ci:��,�[�ޖ�eI����N��.n��yC56K�r�#!�< Seڸ����a HזQ�Q'���@��srm�ڭ�$:jQ��+���õ�1�հ4�h�3�DQLn�`i�׮��ܭ��j֠�P�V���t'7kx�ٹ+)�O@:���3b��++B,�s&^�&9V�c�nۻ ���Ԭ�X1��XE�.���t�wX°��$�-�֎�vQ�Z�`��6�P���Zܬ�Z{����p�u:�j̩���d䈧�����	��h�K��a�جC�Տ���%Г7C��ae��D���J���U��Q��ľm+-5�fA3r�b�pnM��a0V�W�n��#�v��f�fX�D-��v��h��!�U̵���V5��9�oN�y�kU�������r�����*hi"M��(	z�1�ÇJ�F(�sMa�Z��v&�P�m�	`��$����xt�]�(v4b����'�Tx(9���'t;���P:e����ڸ2]���h��Uu6#�)�ٕy�"�[+N^��)�*��]?�"�����!��������^��0/A!������å�A{���8qe���ˢ�/�cwP���T[��,��{J���1?��n��փ{�dq�q��9KN�P�@�+Ħ;���Z�Qhѷ�hȯq���TL]�݄�M�QXV��dn�NXb4/9t�:sq��l�i�Ku���17i�r����T�^�y���֙���u�;�^���9���ٺ{-+7�Z`���n�Hj�k3@k[�W/Y�HR�VL bJ�2Va��f�$��-�W�w3��"�S�T��-V}�/i�BrEQ��֯T6�\Ho�n��n��;���K�N��
ȭ8�襱T����m5��j9��&�Ө�B���Z.���	�u���Ir��e\�Rw-P��hj�ɚ�)Ml�T�l��(�M@�-��S��X�0I)��X�c:v��/Z��tN,����^<�0���W� ��e����F�*�n��h��2�%[)���Y�&���B�C�{sI[�*��,�mk��֢���%,�x��c��
����,�)�M7P���T��tf2X�%��Rx���)n���Ft��50�����kՕ0ĕB���0m�u��e���rjB�70eh-�DV���utk6��R�.� 32Ž�M���RZ�ҕ����GʭmZܤ>�,�f�St��2�02ƥY*��YO ���KY�%؍Uv��j��͜�FMX+��+Z��M��ύB��$�N�s	Y�V��lf]e�۷���u�
�E̚Ki�bd�Q��w@��Y�2U���YIۈ52�-��VU�6�3O5Z��yqĂQ��Z�ƉeR���-�6�T����Cj�C�|v�M7��,��[tfJ��t��hl�
�٢���T��./�y
���J�!sh��3D��^!��,��fF���t�=gQ;�ko%j�^*�X��]*��4��� ��-�D]�#�Q!�i��4h��E���ت����B��}uf�:�(
i"C�e�����)�QHEp!��/�Y� ��QR*�CY}�� �e���L�	�F���
+�W����_ƛ_Lb�w�[��I0�U�L�^*�i%R��s1T7q%�>꺖�S�4�Z��NM�p�:Z+B��N�-�����5�(S���3�`�F����V�K�ʴ��y��O��=��w��:Zӻ�Ge�uH1��M����֤(J0SI�B��r�n9Z�45�,��Ƙ5-c+�Aҧ\���5�]z��뻯y�6�k\�������/fK�!'dHE{׬���a$IMc��jr�a@����}��z���\�G���3Q�Xwj����z\`�P�I����uۛ�t{����י($��(V�vS�+{��d�N�qZ��$̬z�:y�`����&�}-7�{:�./���Z�Mø�D��k�Yڡ�zhY�W=�7$�P��E�ɕ�׬����8-z���h�o�o��xye�!�o�ؑ���:�ihI���"{�
Gp���`��tЦ�n�ֺG�5-�Rm��O&Y	I�s����Vx�]�	Ӌ�,f���m�K��z�wfj-^�cE<�����n�����Q1����ƍ[;��sn�I�Qo[f�����5/�T���*��z+��&dT%�8�g�N�hu5u���,�wABٙ�z�l�w���ؒ��[QdӠ�_�#��]��ݥ��b	���ҽ��E�m�3~��E�h0@5c������mnv�+)�j�j_��!e��YO:VS/v��0�lS���
q�dc�m:�����Uû.�$ݾ�ΰ���r����3Z��(d�����.���5�L��)��l��{�.���Ǖ�B���F�y��ء?,��H��y|�6ji�ۀ�<3�8s��/����x���sJQR|WedWԯ�L����R���J�)��!.�m^e;�����Wη����Qиʾ�*����C/6ZR��fﯫx	D��V���T��������2]�7�Ԯ{�a\ᘃŢ񱋻��$����Q���|5i�I!��~ݿ-�7T�$Iw_)i��xl�͙���zv,���ːlr�J�O6m�&Jc�MS9(�T�����s�u22u���|QnIH���Yڄ� Gv�^�M�R*ެu}�y�ږ�G[vq��`9ĹD�:5-A3H��X[�W��\�y��vm��I_2��7\	���Q��u��;���霕�T..8�[]��TJ��4�{�嬜x�l	{�G�2j�s�щ[W��F�GT˛�i�Ա�vpٻ̨�N�ƣ�/#}v�R�X����}w�uk�7��٠B��2��*8i	�+�+��&��Z�Y�VP�t����4k,�t}���Al|�ٽ��ɪ�x��A ���ݩ�r�I�]kr9|����.�s�tM��d�|ҫ���j�Ӵ�y�ok�S!U�׏t�s�I�us�˒�.n۫!�e�$�:�!N���}av��'�.qG�WgF,b�/T��+imv-�­����*n�GB��
�w.�����1�ս�GcyD����\��G�Rq,����k����|w��2Q�F�s1ڎ,G:<)���7�3*ֻo���+�4��`��K4"�ddԓs��8ke� �2�F-Vh�˴�U�pqQ��o�+�J���ኵ��{�}�]��x��R���o'��tV�MA�iIN�T�&ndΤ�]M�]N+�A�#��R��f�&�iX�걷K���ƷE)�8�����`��8L+�����6�YkJշ�*/�vEN�8���٬���c��S<o���(��;f��Y��W`���g�����g�emq8x�� q\6y:q�%ڬ��BS̹�m���p�u�n�ۺ�N��S��Ά=�=�tFQ��i^�r�q`�i���v�)� �oD���a�Hr�Ѿ��9i]p�}푆�
�S��f�rugKݦpAw/89�Qx;z��F�
�\Y{X�@�?��]^��ko�7LK���R����c�Nt���]�2��yχ+�֠s:��D+-�����^�3mW$���5znWA;}���@��U��:��NND�'_wo_],b��"�n���je0���M�H;;T��"�uضs�wZ��e�k�X�'˸@�<&^�N�Vvm:�k�2���Х��-�ݼ3���{��'�¥�7`��o�6�z�3�'tf_�k������r�]��$R��4�Iuy����SW5�[˕��/���kŭ�����N�۸�����;��g��2׻��Qjj�o
�������t2�In�N��ʼ�j�y������+���K�TE�=�㔊���	S�s��P3]�ATº��`�ڼ�:oq\`��ʵn]�0��*�=�D�7;\�Kڳ;��6�;�1'V�ܚ���wK����_^^����R�}r�Cύɐv�d!!�R�	��k��X� ���/���9�}F��\P�(gl��ۘ��ۭ��ќ,]�#f�hM���r\r�p;ʡ���j�uĩu���\�FR=���:�����˗���Ӫow>t�9�[5��*b�u�Jk+i�`:D�c����j�kǂ���.�=�����o��ʛ;l��R��|������r�Yc^���Pu����-�T�Ґ�W9Ԥ0enC���-*潦�PyR�pVo�J\�d��b�����K������w���)����5m*:	gW�.��]L�|�F(0�o�*��3z���6�u���1�лW�؄;ksO�ru%�*�N�٘����>\!̧�����b"wk6���tu-���Ub.r����t��։%wr���.a#I�U��ɗ��w�A����ne[&�v��S�׽����j�nn��Z����rv���	��������Q����.�l�Vоy#a:rm>�R��R�Q�v��û���ô��ё2���tk %�p{V�Jq㽡������椻������n��e6�r��걙\;��Щn��F�]�_�!#�������U&��E凭Z�{�a�IÑ��Ƿ�l���L��>�lNg�Ow$�llJ���7U�b�����kw*�>S�7�J��2�[�Q��{�t�&wVNr�o3�rB����%�WtE������w�"yu���@��؅��hG�w^��L�΁μ��E�U��[	�[���]L�KI���ٗ�l�"�\�+i�f�ñ�&m]ms���_m���N�\'T��vu�9�kN=�V�mj�a�'$(���N�+��+9i.l��9Cx��s}��;�]��6z�rcId�Z�)�s�ʏ����ʲ�dRV�e�ӏ[]�]ͱ}Y���謓��}Z�܁�C��\eM�(��t��T�ww*ݺǃ	�Y�2����e��ڏi�N�
3c`=e�`u��b��.&�:8����-���g.����JM�x�-ŝ�v�P|�_u�����!ӛq�E.����:3����drݰ�)Z9*����ܒ���B�ke�5�[�99r���ɋk���""XwjEݪ�T(��gCIN��C�V2�˖]���ܨ9�p���ua�xK�@�t��n�
�d��(G��G��ߔǵjj����e�6��@��dn7(t٩�l��R�h)Z��Q}F�o�b8:M�4�-��ZL�']t�lZ�h�:�,)U�8�[��X_vQt��ݛ͍�e�wIocN�m��u��8F���cX����ܘ�]�ktu*z�	�r�
��:�*�_؞�e0��|��	O�ǳ�:u�>��3�M�X�:��cS;rw�u�/�1ܫܒU��֞��:`Vo��X������d.�+P\_TӑR��R�j��symZ�=AX4�e_E��p�W�kc�P8����{�s���t%:�7�7y����wpc�08�q����Ϣ�n�c��.G�g�K� 6���1m�m��k:�*�$�ac����r��k���$t��a�sv�[f3v)��+�����0A�]^.�!�$u6P�I�-�:�&����h�������>�D
ݣΝ�Q��\	i��b�2���#�\�#����5����t�.�_��I��+��=Y'w]M1�\ctKLۄ.���TU����sR�Gt��r��CiQܷvu�+���IW%bpl���y��mB��ڕ����3u������k�KӬ�v��H�쫴�k�mV�޺�'p/Y̜0R���ƾHr4ԽxJ=���%3�a��v�xC:l��iuޞ����t�mե��p�.[v�JI���� ܷe�Ou۱��mZ��)��oe���o������˥����\�KI��e��u+�th��լ���&�ҍv�λbB�b�U��f�P����l���f�Z{�p��0����}Vzu������Y��:N��-A��8ĝ�:�쮏r��!�#QZ����f���egu@�9����1���i�f��-;�k������n��Ө��m�|�tJ���� �K*���Zs�Ɵ���mm�L�
�'.	��5W��R�l�(�2{J�,�k��v��Kj; h�+�3si;�j�1��Q��x�g��,�Ǧ\��R�95uJ���^�,;���f#�e	YJv���,fbPJ�����I+q��s ]��ek�ƦZ�W�w<�d��[=YVZ4چ��R��fcT��69k��H�-}�Saaա�S�Cmi�b`���O^]��:��<��C���9�J�R�t��[+� �o;t�����$����G8�q��BR��Ȱm��zl&��^����]JEX�0\�5ƶ� �e��U����0�$6S�v�wo�P���|
N�e��F�L�\3�e�3]��j{u��C�	�bH���Ӛ�Zs949;�Z�w7NҌIu�4^�[�k� ]�TDĈt�����i׍����k��NԈIS�kl�I�M�ȫx+͘������x�ozp��e�n��EP9{�h�;���_9����S�]����{����X����[S!}J[��&
 DX�T���=Gmܟ9��i�&��wBݒK��us��3�f<-�\���B��rdW�W#��E����m�$Ou��U�e��J|fau
������r��\�F*��ln�Mv�#r澾b�;ӏm)-<�.]r���uj)GuaM�T��d[��-]�S����Σ5_X$���^�\���,�F���OM���e��yN�}���#�b4�߸�S� �J^$n�T��Jڛ�T�":�v�̍�q��2�]��:���Kc���Uʧz���YX��Qŧvhh[rTR���B�S��e�{E����%o@.�m��S�7ϙ9]�����jf�5������6h���<֦P�.�wJ�[���-��׶���٬Y�w]�Χ�\�Ycw�DiwR��i�4�]���0ʜ6������3Σ/��T�����[G��GH�Y�Rƺ��ڝi�z��Hu��\����7R�������!A�a�̓9�)��@(�ү3%s̏�Wm�x�N��IL{w��MW���k��w8Z�����X�����7��ƶ�\�h��8�5�w�Z��8Ō��ʻ���FJ�c�|�^�����ƺ(�p�o��g>]a��ܢ��x����;z�&�ᬵǝp<�u���e��h��mΖ+a����#��x�(��<��|X�Ukfd�݇j҉4�`�ee�u�)}����r3��p=ȷ��>��]��}{u��V�ι�;�ҷ�<�U�RN*��� Дub�f�� ������}�*�ڭ�zv�����n�
��w><7��T@P��_iX�ў�
(�;�����4:#�v⚔QG��̕ P�C�G��v#����_w&&�ߚ�ڝ'0�յ{�
��]�%��671;A�������)��l��Gx>��v���]{q��.�w������;���Ǚ3�V�5�rV���lSm.��oe5��<�o�V�|d�:���k6-ܣ0:
�J��M
7J���V��3S��i��;�J��	��:7r��軉lط�5]mlXr�*7B�
V����|���I�&sr�<�Y��z8P�i�ǷG>x/��v,(Ђ��*����u�4�� �w�n���k��7V�.�.����F��
c��D��VǱ(/(wK��&V�X�r�5��T6u�n���mķ���/R\"Y����I*e�9��W%0���VBv���$�r�!8���i�έۇ�����򎚩��-t�Y˓#C��%�L��L�Z�bv���<�]�X�u4��n]�w4�CU�Y��<�v\�u{�����Cvv7*Gv�Ǵ���u�\�*� ˸��F�k�)d���4˲�c�شw1�����tN�ԗ�e$a��+�j]�xi�tu���ތ�#��:�m��mdbk0 ��1� �H
m�]r�M�v�z\�;RlCgvCMf�ݞ����Y��m�3�\��}w�:M�N^���YT�������F3V��V�'�̵i�/)��DL���pghK�y�eQX����Y�S+稷QfTU��_T�:0R�1�|��g�W*�@����g��]����z!K�P���M��eN���#yʾ[8}3��kb��×�u�\��g�t�S�v��k9y�K�>z�{e%.=ۊ
�_.{[���}.����]��{�����wZ�X)a�γ.�grp�q��o�crws�&�w�c�Ȕ5���=�}n����6��B�Z�{X[��7cfq�`�1���$�8���l���9*�;1hX�ğO#@��]�Y��-��}:L#(�������M�2E�[7W���pL��5�Y]����,��U�2�Rnr�{;�Z�&�e��(�d	B�1m�lv2�Lf�tKI��{�n���:��u!���=��l�Υ�.2�<�gf�L��Ͷ�7M��Y<(̸"9�i���#��*�P[Η��;�P��`�M��\R#}_�ww/��>�(��� O�H{�D+�<��N�����za�s�[�\I̼��9�͈�K�p4�%cŊ�t����7�;W�Ә>�8�'$:M/�Wϣ��76cYu�eE�o��s���"d�����}��S;�"N�kv��ȹ�!��u]7�2��͓�4�����i;Jk��7����0���Xq�$�_�o`� �K�N�wy�W+c�@
[Εt��B����X�M�ء��<����� �f��h��q��r�ܻ��Q��{�
V��t훁���4��[=h�̥�nڛЮ �q�']�Ķ��(�)��Y��֮���±l�*R�ܦFW�6&�������YES��7q�]Օ}r�)Kۮ��8�om�9K�Ek�Gϯ=�De
x@�!Ӭc�MV�M���9����̴�M��]!�`\�[�w3̲[F!����ӎ=�����@];o�ʲ���Z��.ź0&�5�JSUm�[�vk����n�:-���N��Ӱ>�6�p��0��8^\[_'�\:��+�*��r�muQַ.������jN���{��S3 (\ 6	����lb��s�2c{4���̙݌�_\U�1wT!��LQ�	]Nf9��ʲ.��v+Y<p��:�b�(pm��A�e�Os�K4ǭ�= �w����9�nVv��uq�g:�h-��z�7،ГU1���}�]�J��8�)�5���Yc.gu�w-� .��5��N.���\�_��!]���iZ�4q;X�qW�P�%ɚ��@�7N]��f�32-�Ԑs㠅��b�K�d���\$y�-�o�.����]V�e�������2�5Oe�]T��V���ݾ����*S��w�]��U�hۜz�H�e�oY��na��ʌ3�OH�O㪠T`��	�K<1�yBSwe��
FlV��MPk�1��S �b��Ov��k�m�Z2X��_&Or��:^M^��{@���r�Z�ΒS�rvq]��0Խ�°�4�[�N���nS���>�o)�jl�r�ٲ@EJ���j�/�䌽<��7cX���:��Y!մ�F(f�鳍�5���rV_!�`���S*S��6�S�jv۵�vh龥�^����=�["R.��$���� �*�� d������v�ܰ�'e�5�x�Л�@��ew9��N��31�ᢕu��7�ٲ�)���ޛ������oNe,3�O��Z�ͫ�{kr`�ʫ����8�������M��M/e�a �;��y�
���} Ȭ�����JW�(��	�WV�Q=6�ד�9��,�U�V�ڸ1������WPů��ʹ�������)�7�����+Ha�.��f��Ԭ-�NK+u��x��W`#�[�ɻ5���3C@���y}�=��+:���Z:�B��W@�ᮝM&-��,�.��}�n�k(���O�Nv��f�dtdl��d��$N-5�Wj����b;t�!��\'%6�wL;� ���&��}�>��R��ƶ�j[H�@�Wa룽Vyc���N�
ز̩�쵥"ŤI�oF�wk���U���7w�8��ҒF���e���Etn�l�U���I4������K]ܝml�P���(5r�6@��`VpWۑ�'�M�gq�}��S/ Tz�f[h�)ɝ֪�q���igw^��>,�7����C��f�U%j����okZaM���5� 2&USp` [9�Y�3Q�mZɛM^�А. [�T�tg\�7Ճ��mr��1,;Y8��Z�)mDt�7��F��{]YN�[���je9��3���P���{��hTv�ի��|veݷ��ƻ;�"��7(��G��Ȃ��c3 яҦf=��=�;��.b%�u�3���t���N-\
g�f	��o����
&��L�m��Zk^�&4H¼�[�&��9f:�[��U�y�5Vv���Iʾ��Н�^��*KkΘ�FN�u��­�⫰��/�����tI�U�Ow����n�XK,�*���U�1!�I{N�[�9���`��ս������.�ݦbgQ�})���F�`L+_^A���}��lU�Ԝ���Q�@�[��Éd�&ۺ�w_5�o+r�tY�*I5:ܣ��7d�8�*�����#���ONi�k]��:���I��4ݡ�i��vN���sX�**N�q�0��W���"V�]A��9�F�V��6U�Rn�+�qU�W��3F��JE�6��n�pK��Lj��Ai���с�����:ˬ� 9��k��Z�ѭ����h 0	ffU�  @�Κީ�9���8�X�V��r���QKd�Ǵ��e]v�G&����*T�ڑ]�p��r7�c����2�E����zv�͔�YO��SZ-r�[����ּ<@���s�p`��js/k6�O&`�WTʗ	J�c��&��X��Kgm�7Ջz�yu��"ӧˣt�F��Ż��}-T˙�$�>���f�ѡ��'��^ٲ����ќVC�m���rԅw3��)դR�WP'HH(X���6��|��d/�oN��B<	l[�aቫ��A�|�u�&f�NT�����Y�E�N�Cl��*�J����hj������J����]�]���k� ���+3�Jܵ�l@y�@���M`z��/U�p]��σ����7�j,m���z�=6�)�v�Z�@�]&�s����ki6(У֓�*&6� ��^䗚6���v�f�|룇vhJ=hQ��� *�V��*�vʉ�2	t�{)�Y�í��mB�9�icR�tU,�}�-�slS�:ؤ�ݝ�ԛI<Pb@�����)��]�U2 � ���X $���@���;y���w�B{�	��L�	��m�j�2+<�6D:լ�k��Q㻪������f9�V4���Ծ�{:!�/.uL�͝����8o�|��x�Ju/
,��/���le���TD���`Y�3x�kT�c	bS������R����̽�W�*�`#+�� �82
�V3��������CWK�R ���;�2+y�{f;x�9P���ە��Sݐ�F9ٛ1��^BUu_w^b��ZV��[��Y�cf��՝���T��{�7HP�\2#ٛO!IlV��{������Z�n���_T���T�z������ �s���ع5+��Q1�M��m���x�B�ȯ{���cz�@�پ�P�rr��u������@������K��c�"�.�ݛ��a�V&#�L	 ���g���V�=���ѷ����m�v���]K5�5<�Wr�[�D;�Cqή���{]�;g	S>w�]>6:�|�iojD1D�m��	6�:�,�1me�O�W%�d��x�ֲ�淝R�mv�p�k9��p4+�T@��r��}�ڨ_N��';R5�v�����غu�v(Y��_�©{�47D��YO{�}���8M����6 �
�c�;�]u o�����8�����.SGl��N�\)��Gf\Y�5p��@nn7��o��&��k%5I�0)fa�����ԯZ��s�N#�Mc�Z�#�N���˚T�9u.�V��Cwv�
�n�
Zjeo^��S��p}\�[#�v&�d�X�v����.�\P��!�gfV^�(w̞�c\��3��7*Ŭ�{g{�������yY%c��K9�Z7� ��mLy/v�>�V����f�3�լ1S�4GN+��-bk�����G�� �EE�b�s�'Y�o_Q�aR����	�WF�`;̷���)h�7�ھ��A��*�c�;RU���N�*y�o��%3�ogvVRt/��\�s�^1�J� (<��HQ���'04◽��ˮb����:���_RՍ�[��٣�����5ȭ��[w)���)��<�H}�}2�*��@t;gZw��\�nµF��m��	b�;���1G�S������f]Bw��mif�yh�oa�F��i�^f�V����K��9-�ԬKB��M:c7�h
}�>$N�Dv����q�2]����z�3���5�b�W$�IZ�j���z��xHj�W�b��.�K�d,]�A�eƑ��9�v��R�t|a�;[N�<���î&�K8�`�*w��ދq��wi
�4�Z]�O�P@ὼy�k��%E���C�Rn�b�%R(����Z�4��ܼ���
��R�F��
�"�tէvoN	���F�Yz����aJL�u��9�G�#0�.���M��ϵ�2�K.��k���o(����*�lgV��n�s�9�v�]bm��!����#����v����76�wvmY��w��`I[Y���Z��QqK�iT���Bb��+A*���l�yP��ŝ�ʗi#�MS�N����ڳ�2��ڮ�6٬���.�Be����],:���k�MH��x7;{��{�ݫ��Pm�C�;*����������,'-`,LE;��Î��k�]I��;z.�&�t+��m�&֧��6�/U�D��n�$xT�$�u�6��{�v#��Y@�M6�r����Y�o��;Br@� ֫f`8�e�gx�X;��\
g��+���?[b��U�SL�c+�|���ؾycMv�^�Qdb0�'p�����'�s���%�a�+G�C-����*h�M�]yqΩ�)�%�9��u����(�t�)Q�&�^�[���Z� �ԍ�uж�2v+9Do4jX��V&��B�֓q6�o:}���U���A2G�n�<���F�Ty���m�=P(1;f|42u-[&������gOHm�WH1oj�.����� �K�b:�+�V�GB}��dހ�\cκh[���4���ĥ��<�ڰº����K���e��#k��X�2�-Ut�kX-ݻE˰�A۰�gj��Y��}+%WXT4�1uj���t[�� c7.��T]L{��,F�ǔA훧]�6����R�+
ޙsea�ʅÕz�"�R���.�Z�u�;)�d��X�W^���6��RZ��;��*Revmw4�߬�;��_)B��R{X�
������$�,��@|#�֋��۾��ZՖz҅����v&�t����ݹ]s�I���p"�0���\�Y�-
ל
I�W��b{��6l�iV.�l���EܻOFf�O����kǒ���0M��)l�[�����̫���{A5�w��Q�hv9�t[`�b���e�ղz�b!�;\,^��=�:.��Cz�pU�Q����.��gg:%sU�{��lfJ��������i�ޖn�Tj�;�w���hU�s�������Oz�'9���TC+JemUPKJ	\��+-
�DAB�2�A�6���ib"�4��1��VP�2�B�-��+)n\\V��X�WZֵ���e�l��X�mb%s	D�XV�2ܣ`��T)�Q��5��V*�ep��2�DR�T�U�
�ƬY�Efy��4����*�L������b��nR�V���kZ��5QO2�***�����QX�bYhcY��iE2�Gf-�V���5��*��UTb�B�E�*�����EUGh9��������ֵ��PQ-�ʐ�PQ�X�"��Ŋ��R���W[���5�kZUm�DH�e�M6
"�p� �"����2�Q�W"
�f4Ƣ�QU2�T��\KG)e����jۉp�[����]�λ��m�I��}���M-gP�嗏�jjU�$���/�d�˹c�r9n��TΓ9�N�}��%���wEUT�t�$��=��?����nqW�%�C W|�	�&��W�C��&�U9�V�rY����lgR�Of�q���e<��@��^m��o:�����,����S=Os][���g�(�*�P9l���.�QC*L�M��+]����xu)�HWL���N)S�TX����x��3�6vl;	��Z���[�GS�j�q���-2Pz"��F:"�O�X��:�'E�y�ej�0���{J�i��it�����p˧91���{ji��h���>&)��[��[Pm�Z˙��}8�,M7��ކzs[��啁�r7A�lդ.�VMv�mt�8����0īhVs3��z�:Y��<�/HC�i�U�����e��H�@����R�H�C��r�RV�TBwK��Wf��.;�G-u�!��N�������5�q*�i	��S{��Du=�ͺ�Tk	�fd��_�)��+�ge��z�re7��,K�;
FquJR�D}K]}u�e�kY���s����FM}�Eu�w�Jux�^}[#V��֚����Yr��I-V��+p�Qq5w��v+Ou��u����\�e�ʇ��z���͉N�}j��{���ם_lb�3�J@�?�(��Sٻ �-�y��j［���TO�|�8��M�)��Y���J,R*S�;���ʍAP).���3U}<���=�̥8T����|^i�j���v}F��ε�̆'�ެ���{ε"+t�i�Y�l�4	���YJ�t���8�m�N�oB	(��О�1Lir%mg`�f�j��0�_s]Ѕ�l��Ԕ��"e�eI�}�1���'3�<�Wؕf�����-T5��\m�Y�į�5�&ĞLeU�j�ϱ���)lgU<�00nӕavv�Ή�C���ji`��vmr��q�햖���m�R���6�)ֈɆb��J�t�؜�%��`#D�s8sv�&���9����s�:��s��k2�u�}V�Z���YiC��lw�S�*�՗`h�R��ك��-�st�]Fk�Ԫ��:b1�L�\\H|L���(Lf(�����W*M��q]=�#-\�T���~q2�npL6٧���媦�AcEuX��#��p�቙�uF�γ͵�M�bX�N���g�FE¿�\Ȼ���o�<��S�s��'tw׶3�9yC�ۢ������Q&����u�<�Ӟ��q���Z��u�k#��د�d��:o�Bۅѷf��W<�*鰑٩�����w-��MrZ�Oyq��:��.rZ��c�U�����Zd��xr-��yo�����_�������R]�H�idgyW�Ux����V�����Ж�����r�[~;��,q7dG~YJ��Vz�z�����W�n�����+o@��(}n>E�z.vzɭPP���b�n�%��iE�����D��8��;_�4G:��W]Ќ�{C	�~.��G�����II ��{���W�D��_X�u��8Z�b���H�/�ۆ��c�����ԠG�-eϓ$N6v�9jN����V�w8��-@�Vgq���,�/0��<�̮��W�u�˟����R,G!V�IJGqPDM>��&�%�cx��E���Q�#�`4��q^�Xv�ʸ��-R�trwVzr�0�u�̛Y|5�P%�Yy��6kdg�OL��R��F�6���W�Ϛ��q��T�z�"����wr[ҧl<y���	ҮOZ��?yPu;i�͠�a&���m{���Qc��f�qbm��r����dPk2�]W�s��P��ɩ�(��Mf�ӓO���2�zv�k��6�)�!���\��	�gj�7m*"�
�n��l͔0,*bs'5*+�].A`�,�W"�9"J���m�9j��֔�.���F����s�{Ԗ�t�S�[(H�F��v���kp+WW@�m���9�Z��mF�k�LJg]�W�t�v��[��i,b���a�[<�yED�P����5�i\�v;wS�6���{`��q���u�{lٰ���D���7�u
/�J|��۳=٩oJ��2�uj��-"{��`G(��>��R�a;���w�KY��\�u]��mq�l�m.��F�������K #3���/����w�K�|w��{9�h�㐮u�-�ޕ����ҭ�!�f"���P�["�*��^=L��Qӛ�=���/:q���L�!�C\���3�ob���%p�7]�D[-���kL����]N�xF�v>�k��g�(�VϷ����ⱍ��S�~�ߕvF�R���Q�+V��U�*B�J;��{�V�y����+��̧q�h���;�Ω!ɯ��	0pL��������s�Bf����m��c�\�w�&�:C¡�p�$&aqpg���n��QW=�'5�;�x�+�{��(V���m��+]B|L5fz�|�+��W{�t�Y���ꚿʨ�MRn�}�bW7J�K�4��38֌���;�� �H�a��m���炸�󷛈A��:�V�j��<���z'q�T��4'�Lȵ�d�f�����n3t�sd��޿�Q���Jw���)��L�Ïj�W�w�12�\ƴ���K����>�
��,{S �$��EM�=�ձ^��l�����"ۧi@��ъ�v���_oʬT����Fqo5kWR��a��X������I:6Xޮ�����~s���t��Uq�}�iN��KyU%�1 Ň�V) �W]ϻ/\�Y;�2َ�����
tj��gVt�50e��z�1,�3�}��ǛY�:�4�C����T�r��T�]���C%l�}�ғq��k�ZViu�Fs*wa�^㪴\�q�t�� �y�vin!s{�>������[݋�z��)Պ��rC4;>�J"���̬�k���E�Au�R���Jΰ!mN뤮u���w>�Ə.8�;�@��)��p�1�̽��ٱ��x;n���hj�]E������A�Vʖ�%�_�q����쏹\ҳ6��6"88�:JR;��!��/t��<�x�6�y�X�u��	jW	�!�^*�fW�;�)X��u7	WJ��B���ꖴ�ڤ�5�#2��U�5B�<�]��/١OW�4��c�
`�\�:�v��K���T�(n���X�� ����pMQU��&����yڍ|�u���+tY��\�к�D�-���۲�J$���TS��C�6����5��@��g�����wo�b�ڗ3 ���E_N�|�g��;�7.��$v\{;���9�:n���\��R���Q�΍jB�U��]��;��Z��"u;t��7=��H��X�v�t��Mt������v����rX�9�{�����S���N�{����W�+��7Gu�ƃO5-��-����`�z�gz�)��Y���-,�����8+�R���F�9:ތ��L��^˾�t��/��w<|iv�Z�.���VՂvV3��Sk���7�����7E�%9��S���CZU�*��}�M�%��t��tw�;�=��]�阸6���Dr1ԡ�E>�ܾ�R�F2�ޅ�&!� Z�¥�7,�z����O����B9��A�����	ച��H(��eh1C[�u=��gs�1>4kvm�����	�����j����� �rfD("�i�4a�W��1�Vx�ov��)x[��y�	�C������ؗlP��՗8=R�ڵS��ܴv��6v�[�|5�₳Yt8j����}{R��̱׵�V����[����Q�b[�:ݜ� �wh9Qoa�N󷙈�Kӗ�V�Ɲ>q�bv۷SÓ�}�.��e��U����ɸ�/�L�-�x���(�w��]-&����W���u{v02����4g39�w-�os���9�47)��=E��4z"�{Ҷ��/�յg����&�¯ّ�aŪt{Q��ء��OԸͺ�в����⭾eqx|�jlG�Dop�E˪�\��0��:��%�{�]�/b����V�����ψ"{�!�_d��� ��n�>�yPv��$��=ϩt�VPєVŸ���U}����)*j�ܔn�i((�᥺^��q;u3l�ۙL��`��Fҳ-����}*,�+�:u������M�;:�w�m:�gd���wb �bNԛ�Q�s�6�Yt��ێ]���w��۽��quL����w��)U�Qq��=5܋ƫkf/Rz_��;�T����}ӽ<;��v�S�?9L]�*��>5u�;{��<�-{lR���O8�b�8��B���O��f���V|[�V6��Z�X��ab�_r&Zfa#��#2Dq���ȭ�̋���t�ف,X� 1�B��6��-��5LMn��Sn�M����n�1YeL�pЭ�Ŏu������1پVf]��;|��ǽ��Z��&�v"��M����^<�<r4`c��[\����u���^s���<hn�P�\w۰/�����ߎ�r���Vj71��B�5k��ۺ�E�����k==�'����0���+��:g{�{<?@ܐi�?�`{�l���}�Z�+�7�a	�ow�7��P�y�yf�:v
vd��Z��sZU��c�Txܸ�:%��=�6�	���tN�3�P�o:ϖ>R�T���{-We^9�@�Nt:�v�<ݥ[��s�V�`|7�\ݹ� 8���VR�\gD�����P����O
M�nҜ�Ǵ378�]�Ty�$Q��]��T:<��_4���x��`�����(	���f�W2M�#G>t��l,F��wE�G{�Y�y��0�i��s��_Uq<�Y�a�M��WVM�Y�hWi���ڄΙ(��\��ɝ�5��CC�@}t.�skd��.�ά����s�Z"�C���kB�u�����]���;�!�p�e%(^�����ӄc��u�n�נq������$��y�ؖ�9n͇dݣ�wSX���;�����d� qI4*���Z��K�SĬ��T�;�y�%\�܌V.t�M�頀�x+i���55V��4�s3�y2<��X"e
��X��]wam(XP��;z����{7n.��e7���ֽ����ej�����p���n�1�4�"�0�[�s��y�x�+7�y��م����]vjN���̗�ju)%�W���|<�17��S_NH��	��w�U�W���{�#�D��ԩ�УgEf:ɗ@�ݓwfI����]��.�T.���t�8.���O�"*�(��yo.�;Vq��K.5�d��Q���[{�1Q����|�
�@�F(v^к�X�Ƿ�i%�Il4��X�e����֥Y�R�Yv��՝7j1��CI�,��)��xN������0a���]'n���O;w+�3���Tj�®� �ːZ5m�?`^�j��]��[�H�Kc]X��R]8�騨L���a��Ԥ�ʊ�'8�۫)zt�ؚ��d!�7j]ECXiR��fJ���[����+(�U�-	$O��Z�u�l�x`�#�p�]n;�v�{��E��.�jű\�Z�Ⱂ}�t��]�wl�,�X�\�]��O �J����ѡ��b]B�m�ƥ���@R���U��5�T�<��&���+���T�s��ׂ�s�1G����B�����6Nqc���v"�ku'��4M�����w��o��֏��\�E���ܴՎ��[!.6D�Oi�2�i)O�v��|���?�eS�X�ՑQ1��G-KiR�31eJ5)P��������^�`xƕ3�KmATL�1�`�e����h72����l�r�-jV(��Vʏ~y�MElU]5�"($Uc�̪1A"0V[*\�*e(�j#{ֵ�鸔U��-,�)F�V��YjX�����UUX�c�ֵ��k+j�2�V*
�#J�%F��+X�b�(��PȎS�ZքԪ���֭�QUT2�m��n8�2���9�kZt[eUWMKmJ�IK,Vҵˊ�X�+�e�1֭�WKKl��lu�k]饈���V��\�J5cmJ)kK312��p�Y[3(8��QR�5�Tmu޵���nR��VҪ�"�m�UZ�V�l-�ҥJ��p[h�B��J�h��bU��T��lLK��[W)UL�b���e�ȶٔ������V�E[e�Z	R%�؞v���~	y�w�C\l�3x5��<zyU�7׍s�2����`�p����OR8:�`FZ]J)�B��Ej��o �}�
y��q�p�M��Kq1��sNz�k|�VwK����;i1�����d�u�U[�2î����>�۱�Wk4��!��y��m7T5o��Dp��0{�p{k.����A|�+1X�!易J�T.J�>~����<]��䛡��]_�dM�Ҿ�a����ђ��}Ra�+�:�m�u|��b'd%>�zn���\�č���c%u�}T)���Q���Λv���j�-����N���l93C��%��\�LQ���J//޹�W_(4{�����cy�*TSb]!��x��^F��T����wCv8���c�T��I�߽�!��Ӊ�o�g��,��)�R��~旀�ial;\�>q�6/�G��Yb=�S3�\<�\�5��.���_*w/=o�H����������t��^!�/3�7nt�V�=Afy�T��;�Cm��Y����Q]�o�t6��&<N�m����?��'{�I��io�����& ��h�G1��,d��O�������+�T!m����+c���(���ֿe{�����'\���������U]��f�m�U��ޙνIb����+�V9����k�evn����+�]ať���������c{E=x���~~]J\9Mߵ��K��~�ݞ�y�k�W������)�^N^�����JMW�ŉ0�U�dS���<�^/_��8��:��2c\�2U�G�G*�]>��΅����5�ё��W͆���rTUVzz*��s�ؿt5�4�^�?(���'&�j��W>��J�32ra�f�r9��}9��.����m����F�M�DW��-nw%��N�򽿣�P�8�_�>�d7�t��@.��_��˺��k��������7t�N<*�C]���(yW��<�ޭ���b�ث�Q��vl����ԏ oYD~�g_���R�VW�G
T����+��W+n�J㮋�a�%�7#ޱو��GZ���Bs���� t�\��ϝ�r�����뿺�bo�/I�.�8'��ġѮ��_K����n�%b|�X��R�~����c�,.��h����k<�*&�1�o�4�d"����G�9z���&>��z�{;y���4�{ı��c/*x��y��A��Q.<�{)Z��8g����\y���PC����O�ة]��>�S�BZ����^{ҳq�����~gi�dW�n�*:�;�g��I�����L�d����|+�z|SN9�����>�H���n�^	~�qɽ��*�^b��9���s�}��x��JO)ϽO�P�ۼ���'�r�-��=#t"#|3j鰬��{���~���N,�Mfc)Z>^��dS����������"|�_$o��3.��WX�;٥�_>d�/[���N�k���� �Pw=�E�@��B�.r�uB�J�
�]!�ܭᷠ�z�[�����:�f� ���w�i֜�ԅ�}
o.J��;�X�c2�d�Ϋ1(��q����x76T|����U��3a6��-��ޥ��������u~Tј��שEz����2ڍ�Tgֻú}B�^l����9$Ȯ�rm	�+=��o�jS[�U=U���BI��GW�<�	{t��.ע��gr���g�	�j���{�_%:�@J~�H~�H��r̏����W�����\yN��ą x0=�I�_P4��d��&�t�}�'���q��yHi�Hu2�$H� g� }� Q��=y�Cމ󋋇�s����WY�o��>�L�I������'�+���|��)<k	��4¦�1'<@�4\��0���!�j���>�@O��˳�[\�=�u\�2O��d�}�I�O�c�[� Vg�=Y'�8�'�'��!�Rc�'}P�����d:5Af���k�]r�����ow�P���� )��+$�:��!�,��	�%�:>�$>d�:�p_XO�=bä�	�� m��}���}���A3ރDZ��fs����}{æ�>I��uB�q�}d�OS'�*���=d�Ӥ�|�L�2���r �g���|���M���{��n���ӛ���B?폆�r��C�O���h����=E��$Rq0݇����2z�C^�$>a�I�򟀃�~��0��[SS�&|7���0��ی�~.���rN���1��ũ^rt�۲�;j�r�yz
[�[Y]*�)��E���nz��\1�<��{&��a&�%�m*ٜ[�'�ky�ٍj���x7QFgK/'V�����m�N�`�>���?2�`� G�9g���N���:<���d�Vi>a��6����e�c=I�O�>�ʹ�U{y�����a��O��=}�%Hd�&���КC�N�����d�T���	�'��w����|�}������^9"d�j�ʗ�XVL<a���C���̘��l�@;�}���3�a���ve��2u<Ϻ�m'̞��y�'��[u7����]��e1�����l��g�3�I'ht}g2{�z �1�=�$�$��C�<C��;�`i����)��ȏ���+���'���ҽĽ�ڀi�&�yl$���8�r�����~HM�g��9x�+':�m�x���"��C�v v�u��Z����cn����i���{�~�� 
�T V�q���ORwC��;~M��9��Bq�@��2I��S�#�~ B;X��b�?n�����'ﰒ�[8��&�aٔ��u���m��@ڡ8��C���~P���ć�'�0�7I��wx|痯{�k���|���*zσ��P��N"�yl;�Eh@�y���}�t��q4w�I�O���'H<N�Hp�>�����?Jɫ���o�G���>�!�CA�	���h��>a�{���	է6�MI�l�'Wy	�S�0�� �	�4���s��_ey������׼|�m�c>��|�3��:Hq���2TY�쇨}��=I論�I2e��N2vL�z��N�����~6Y��_�*������8��GQ�['��Z	J��㮤���-W,۔�򥭅g-�{�X�1{�htl椷z)>λ��n�58���\��>�-[��V�T��T�=���VG0�H��S��� ��o�;�m�Q|���i�0:�`���I�I�
��H�s!�N�1s�r@P���OXp9E�L'�FXIS��z�\;�~�>ˮk����O�#����@&v�vw`,�����i
�e$+Y=E��s$=d���i�bb��Q��r5ly�*�.�	��1�ɕx����I�ِ>d�N���IY�k �2��>H|�Ă�`z��+'��(|�$�>`z���TRcP�5���^df/[ O���B���#��t��<aā�����>f�i��$��I��#�{�E&�'�>d�5���<n��k�{�����P9l����|�t}�@���'���b�3�'ya;~�C��PﯲC�'SvLd�twd�'���j���u�uםk��<ח߹�ϡ
�a̳�C�7�����X�Iv�!����Xg��a*Ol��L'V�i�̝yC�<~HQ�̀���Li��*���v��<�N}��4œ���}i׶���X{Ր:���'o�N���bϾ�<d�{�x(J���d�>f̰�~1~�!lA����uI��3�� ������Y's�i;d��ߔ�a�֧~Їɜ�I�I��C�;~Bw��I�Rvr���Y��ξ���μy������s���i�iY�PdϹ��<I��=@6��'=��I��q�2`|���2S�q'�����M2H����g�.�v��^�|8�g	�}�C��d�:�6��N��������>���d�2q�֨q!���c���?W� D�v�e��fo)�3�L��v9cDZ�����r
�m����V�ֺ^���c�8̥��ai"�kH���	�,Q�	��y;^���E+WNujj����5��f���"����Ɍ]��%�sN�k@�r�;Wb�`��Ɲn]쓶������'��Bm�aַ�P�$�TY8�x[>I�&�'ya=`u~rI��{d�P�T�$���٫0<ݓ��9��<�����w�^_=�����8��'ք�!�V�i
�Ͻ��:>�"���<�|�x�Ψ@�'G5�]�C�3��q����xz���w��0,�G�0�����|yH|�gt�	�9d��w�d����
,��v}�E'�'A��q���� @#�w>T7U�mߺ�7�'��XJ��>��q�f��2N��w��x`?YP8�VJ�׻�OP���E@״Y<�����߸&y{�Z��^�~���OY*M$=a�|�I�G{�<B|�g�C�x��b�S�(�>`�_0:d���ߺ��>g車Eҟ� �����mmE��^{~���g�χ���,���e��%x��VN0<d�r���Tē�>�$����*fXC��l=d�G��a;��E�V��dk�^�I3&!�,��
�g�=XCh���I��I_�6P��gy	��_Y=H">���$I��2 �Uַ=/ǇkZ�^o���>�E��Ҥ�'�O��d�2e����!�C���|��(���$���4��Н����&<~�2>�ys1��3U]��oG/��N���IRi�!�,�g����t+'̘���ߺ�Sۤ�'̜E��'��'Hv��Y�s�^��o5�k���;�\�4�|j���&�@�'�:g��=fr��Y&3�,>d�Н�u!�M8�G��m�ɉ:���d+ԛt��gX�yK�u���xsUr�5����T��h�T>��O7*lx�/��E*��1�y��΋#FP .��(��w����Jdn]8e�V:!�������_T��-��Ď�bxz���S�-��{�桷=�[�Ŝ��
����������������P+$�VN$�N�@�OY>NϬ&�>f�Cצ��t�2{���?q�O�|4қ>T��������^	P>��=Hu�}��l�yg���fI�)'\����a�2}i߶H'�&�a�=I��A�N����~��}}�����OY�bO��I�$���܊û��C�ve �L��Y'�;���)%��O����0���������;m9BTF��~iިkw�bc	�n��2�^2N�����!�{�,�i0���&̤6��N�������>�Iǳ�'�����Z5�������'}�/|>�(�f��G��?�=a�!�'�(g����q�1�z�q�m;���!����I�Rw���z�W��� z���	t��=�w��w��`�'Ƭ�I�x���X�>I����g�N$�y�2N�9�P�aP��'}�(E	ճԜd�#�8|ED8���{�����G�����|�Y�'a�hݓ�4���I�;fٿ,XL�g��s$���O_9� ��>$�������?o�؅IKv�W{��֯>M"���2wi;�6�淐�`m�k܆���cX`o�>d��Ļ�����':���g;��r�>��:��J���"�@ÔY<��.�4��d�I�N���z$��,�2��j��`u2�$�� � E�K괟Y��^�By��$�/vd�&"ϧ���OP����$���)6��;aSl�Rz��'ow�gTv�m�l'�o�5s�)���종�LQ��ٲ��s��j�v�;�'+�}�;e[i��U,�E�Ő�ꬡNyҴ�0�F�Uw�:�r��7C�k��@E|ol!&v�Z�	�)>���X]f��H��*���m�Ň�mZW��H$I$�c�����ރ$�J��$�T1�X��=I�La�\��V�T2q�zRI=��+��w� m��w�Bm��5*�rc�|º��]��<"��큐���3VVI�u-Y=E��P��[C�hO�+C=�a>d��0��3 x��'&N��]o9|����IY�{�C��<Hq&�X
c�딑I�x��H�P���Bu9�J��&Z�H����� <�w%����ݯf�U��~�2>�a	�>���Xz�;z;���Y� j��'�6�� �OS7a�
�Y�|��������LB����3�9����ߞy��u���
��>�y�XC�)4��w��O���vã����N��c&�d������}Bi����X+�>W�m�Q�����j�����"�b��~a��4���@
O�E	�Ri�0�KBi>`u�`z�IN+$��O�=E�I'>����מ�]���u�}!��%g�a4�=��:J�}�4��&0���'��]����;Cl6��1��d�y�@6����=~$}�}ʋbZ��33��zS��dG�{)8��'��ϊ���4��iXq��C���Nَ��vM2N{��CI���
#�#�4��#��V煕���v�\ߢ�<I�k$�q���>��>d�=N�d8��9�?$���x�s����jo��'���Ȥ4������3�����ֹ��=E��RI�N�d� u�'��6����ORj��Rv��q��o-
1�ҫqw�UP%yt�c;J?
�W��XPXO�{U6�5�.�8��eNa����>��ql��=-E�"8)�^O���ko;�Rt���v�m��m���u������Rv��l��[�&��l������>���*�dY3��|���g����=0u�΋�tm�ޠ'����x��dk.��hI���I0[���a�#z�g�s�{�1�GO����մ7�
�����G��{�}8<�g�_9�;h�C٠#�%ձW�l��<��N���{*��ʹb�r;h)i�	*�;k���F�ܼ��ż��G��b�ũ��O۩@�	[�bTk�y@�����܎OINq�G:��Az[�?t���̙�ɞ��lt.�-��C�	j�f��BjE��C���t(N�n��6<�#{�C�*݇Y�[���?9�vr��e=7gn�s��w�!�6he8\KTwE�TS���	j~���s%S�����y�n��
�Ey��zbG�ĵ~������A���:W���@��@pﴅ+gӂv2�_�E�SӒ�^u�KN��O���δ^�Ү�|ɲ�T<�+ �]�����Wّn)ת�q'V� Ұ�K��J�<��7�E,�+\�N&�Ys3�[�@���pס,`��q�^�tM̺{7MX���w+'-(��loe�la�p
�dԵeZ ��"�0Z�7�����Q�Q.������8{2�]�Al��<��eq\FT<��G[�k�N�8�a��Il���X�#D;s2;���M�Z{WT�[u�jm�����ܣ��B��`0(�AWI̺��bX��T�-}�(�Ԟvi�+���u!���uEێi��	9�˸UNqEW*�b����F�%�����,Ĳ^���y�G&ˮ�{d�X�\��r��a�H�V1�DoW3�8�V6t:{�iV8J��Yy��_mmF ��5�8R�7+���;N}���f�ts8W%�I��3鵛I[�{�jVh�u��e�r����/��t�̻U�Y�  �]"�镗WRVW�l�O�*u��g/�3%�5^6KIrY��Q��#bv���&�Rz��E6�-�jI*[L��K�5Ck�X�⮥z�v;pE7�7�ims����k�M��Z�;͇bT;n�<l�3ss��c�l�;V�AD�$ I��M*�͹j�ԲO���l�1U�����Q�^���Fi�����r�U�n�D�:W]&���X�$�)�]�R�b���F�81:)潻 �7�G�u�՗���L:�5�\-
ʹ�=�l�{�`� 
$��Q(��H�h�Yw���M:�mĆʽ)b,�m�Ъ֚]-7�X @�Kfśj��6
X3*^]��J2�,(gN��)�g�<�4�*0%<ˠ�p�Kl���ƥ5�]�Yn����ˊ �l�$�XIj�cZ�D튴��]�ܝ�Y��}Y�3eA��*uaN��a��sY����q�������;�[D��h�)����-�o���0��,��9h�8]�H y
�o:�x�P���!)V,�N���qp����)�*�\���0��Mj�Wpt���\�����@�ٵ(��&�2F����d�&�aܽ=�z�n�΃��]K �wt��'r����j��t��ow��!v���ƕ���Sm,牍���%�*�b�=WV���;��SQ�1���8J��s3���\11�k�;)8���]��J(�:'la�{Ӝk�}���|� F��$EiT����_�h̴��ff�r�p�㖍hܦ5�L_�浦,�,�ժ��benZ�mlX��bb�+V�q�j���2U10Aֵ޴*i���
��9mJ*�+�r���aG.\��X��,R�Y����kZ�i�KF�̵\��PUV.m��3��(���Ҷ6�1i�j�9�kZ҈�U�0�5S���c�i,���Lh�m�"c�T��6V��k�kN�R�5T�k1)�AE���L(��G.,b��6�e��[�w��2#�C\�V"EL�!m��ETb��(�sZ�Z��5�EģX��l��\�V���V�BĮ&+�Q�T��z֜h���X�5���4�Js-rbJ�V�`�̣mE��e��َ9B�3(�"ܹm�4KL�ҊffAKU�-G\���r�&!�8��ۜ�|_:J�c�-��������ۏ�hm��oF���\Z�(������4�;O[��E4�q�:���ߛ����5�s�|���,X��#�O����'������5�3�3��\���~�ޟ\��龎�.�^��/ybI:�P��f���R=�p�<��VQ��oZ_ts_OJ��º�C�d�DFh�Ow��df�K9U�H�͑�OKQx�m䒏U��ӉU�)|r��M�1|��g�IΧ\�����&R�5��%�~K�Z����B	���Լ���j������/���voX+��̅�[	�}���_nk���z���ˢ,5���ߺE�!%K�ew�|���1�N��>w�g�s���l���}����y��}	�`���S
�Ȫi���(�o�B�c��[ڥb��C�gp5a봱z�t�|�K�x'(h�����оz-����
����v�3!�}C1l�*Y�ra�,�VVwn�k�H\=�'��A���f��T�K%����Zp~���:�]R�@�)Or��eb�/F�w��<���g{�FJ=4��/�W7���y����b�`,�E��\u����]ۿ.'G�+s��ÿ)����Q���}	���TU޻��c�]bx��x]�J+hni`��\M��rOIk6]��(11�4����)�/��1T������w����Z��Z�,�P歡A���m�����0M��	�Fk\���kM'��S�����=o�Zt�W#�wl���MW(���ȋ�V&4H����I�+�w�w���m�p�zbn;����[��#�C&�����5��\��c�z�3ft�:O��7�KE*����Pv�s����tI��3���2��kޞ�,Z�W���vo&��n�
�`�31��z��el��	宺�=�o�u������.��\iԯ����Em��S7س�
��uʴ)��d513f�0u-	s0M�ݺ1"T��S��Q̢u�uS���������cҶ��JIe�nJ�M1C��vz��և0X�a���]�)u��}����]���\9��k~s��E�YAdO� '���_���UK��9QE��9���*]o�t_C���GaV7���_K������"�+uKg�qVW�kx|�{I�u�;��ݪ8t>�b�!�o#�^!����v' �%-��ED��t�܅H	(�+�ll����Gl�*$W{|������:C��Qg�z���8Y��K���"��[&���yiC��ð��:JC6O���h�Y���ϳy�7JQ��u�b��#P������^7�υ�,I��*����Ri�[ Dԍp%.���¾�	Kh�v{$�ou���So�˳V�C�������~���oyՂ�z�^M�1�&ݻ��r��ʜ�7�w�B~���ɔ�TO0L�ϕ�VfM�e��Xt�6"�`�c����i���3�{��N�Ӫ�27&��Ww�Rt�T�,Oh�ܯ[�(��ҷ�ѝ!s��+f�u�׉�M�j�޾iq	�\�ߜ�]�~�|�AId� H�|3չ�?wB�?����⇊�T�=j��J?g󧴫�l���~\�%���T��v���v��T}��9W4�Ε����A쭠���ъW�:L�{��gdr���O+�B�Uj�
����N��dP��V�L�Ʒ�J���5`��m鮜�ơ��&�������y���1�r����"�/rݫ�}��C�V�y�
�<|��&`�\�4u��Q�پ��}�q]�I����������h��\� w�tm^c盉N��nDf�([=S�C�R	!�J>��޽ۗ~�Ѿ�O}�c�N��+(n�'BB�V)f{6�r�_R�B��*X��v+@�j�P��)	��}4���y������ݗ-�uD]��1yg��ܤ��:���ޘ��Ou�XF�*��W�n���L�:�u�u�2��u�9K����jų�`�#��ώu�����y�O����|�OЇ�H����	�ﾊ��K���$hтg�}Q�c�5W/>������XryR�r���gz<�wN���څp���Lӷ_z��C�b���܇�b֩�j/8�O�qP���V��2�uK]���o�>�}�zV�a���D'oy����h1�r���EV,�w�������������鞚�czU��x���z87Gr�]���)N%U8�W��ｉ�ؽjo���;���#T����n^2��%x-җQ�3��9����t�VcG��J�����d��s�BDb�H@��v��Ν�}�U�7�5�7�8�U������hq�n�b�����{]o�ϯ���V��=���4\���_n/�<�3�=�����+�o����Cw8fmd:eq m�}MG��sէ̞�μ�ˑ倍A�<���
w�"���������W�۠���`J��o}�.̝W��g�%N�ՙ�˹4�hmι����s�k�s�� ��,"�� �|	�|Z��(��O��u�m���خ�ԕ��{��Y�l':{�5�;�|
sMOմ�60����]S�D��AG�'MUj���E�e���ʠ�Q���n�%�����p!d���N�$�^<�����������A�H��7�n��b�}�5ۥ�o�~���P0�H�7�}2V��Q+s�jwo���1lB}�A晕$9�9&���ҥUF}[���M�j���y\�qE��:<-�cL�qp�6���W�[�8�2���l��/5�R��S�o��vy	�K�}�r��H>ֽ�z�� ^r��:*��n�h)h&�;�؊������u�p�r�R��7��.dZsS·�i��?$�t��Z�Pz�*�D������0��n�f�̈fv��t������m�!]�L,��8�O�����Ǌ�u��Z��\Q^*u(�G���mr�u�w6 ��N������A�u����y��s�� 2�XAd�� ��`Kޯ�/�����oo����N�z^ʪ��}YʄDbM�gn�<�#T-�����R�U���^�B��X�E1�*����ϕ�%��v��J�zy��ɮ�^�6+\N��YW�֌���)3�|��o*A���c�6�Sb$�RE���0������սK���CN�3ئ�Q�\�d��ǽ0?@�9Ǽ�W�},44H9FM{��AND���wFz�6ꫮ���	@T���Sh�����R�u L�!@}�V5YY`�	�l38�71��G�)7�1�@�Ԡ�+�0܉�,�u�V��׊���q��'儦PZ�B�Jj�R#�=�ͽ�Qv��ҵ���X����|�-�`��&L�L�!�yc����]v3��s�I��t�Pj�ǅ7G6�Yʐ�2����}���M҂�ζ�.ơ�Jf��\�����e���\�Q��黻흷=Y�w ��"p�vQ{��T��ݖ��Z=��t�,���\=�����Gx���P�@�:�仩gA����s���0?<2�u������9޷��� �����"���Hs���}���p�y��Ʉn�����Z\楣9w���]	�J�E��D��N'�~U2*���s�e���h9nnf%b�ơg\qb��Pl����x��M:�YN����}�WW��t>����]
�b�a� �+�´-�,��bc��+������5�
v��gz��Wj85�A���m<y��"������:�.�y��w�yu�D����]��Ė��ښ�t�6����}�R>�޿S�����]���T�{�B7��R��=�Mg��tW����eR�^����G�!�췑���bH�-Oàh���<\n�{��P-�jӷ|{��Ln)i�ccL���Hޜ�K�3����Y3n1e��"���Veq�nI�H��\�Vv�Ȭ��Vd�>2]�������:DR�f93�\n�&L���厡���[3�P��j;5#й]$����|X@�)�� �Hh������{�Uo���Ͻ�p�W��O��ǳK�6оk�]p�C�P�Ru7����E�l�	�P2�m�1\���&o���Q��o�1��J��{�br$<�q/��NJ>�C��.���)hET�t���u��q�f�,�^�KȖ#DW`�r#�]��V	E�o}�%����V��w�`�9.��8UI���R��q�R�mB��^���k��������B+�Tf0�b���5y+��X�T�Pj9�JjW[��w%a���3�4����9;U�U�2.�2ć^�em�
9K��tSyq4����J�_g����_�J�+}K���#I����SS*�z!`YSN���;]�������dzc��S�u�y�@�=���(eaBb���O��X���ŷk���b��S�(E��5ʚL�*��K�,��P�b[s�0�m��Vu����7��f=�fI�����@�H(aaBA?}������{޾T}{r�\�M��t�yw�gy���m��i�˦�ls�ٗ��?6{&��~�/���1OԄ�;O�uNv��rU�V�]�O5�|��$.�)v�[�>��]S��jg�;m&�.�ӌcr-F�R�{N�� �{R�A�ȼ;��V��_�u��}>����i`����W|��4����̨��ޕW]Nz�zâw��u=�۷Fd���kP�n0����U{=���H��u��Q����P-V�ܬ��G(뙪�55��lG18�[BUp�p�]�p�����7]P̌�z��4XSq/G��ΩdC#D�8}�A��C"�f���;\�l���ƅo�V��(Ai����p\��z�}� o���U��'64��u[��-��1lO��GqM׷��+�8(����\������$�oA��<����i�����g(�Q�Y��K�� �^��c8��|�>��"�������Lb:t-��kj�R�9���~Puh���<R|��M�w�k��te��Ah@��&������|�%>j��*\�{���Bv�خN�7԰�
4t+b=����dv�Q�㷥N�yΤ,���8�9�\n E��Dkb��u�_	o�ޓ\byJ�Bl���]YyCgr�)3��Ջ�#����r�wCo���Kۘ�_��T��֚u�3���~�{��R-�v]��D2���5l=�n���G�N�ru�	�����BΫU)�H���qP����ɱN���a�}�yEΒ��$����ԲIgjhĠ�raف�dދR���iPW�����3�{����.�W|a#1<t]�,,�XȽ��j�Q#8t�*Y��)n�=x��Rr=��-˜N�f�9�ϋ�{�A�`�������n�{�A5���㷙k��W�r>!c����L�ДZ��kB��١+�k$Y5�����W0��ύ\��M��7G!s\g_��נ�k\Ğ���Ӧk-�S�mw�$��W�H�f�р�p&��^��Yb�~sF�$�f�%�W�M[[�aq�2Z��f��Jr+�H@�N]�a�oMŔ����J˼�.�X��Y �@��tз��'D�Xp�c�l��u�ݸ�~�n�b���8m�ZA����E�3dZ�0��V;�3?a���چK�^��h�> ����*�W���=��X�Q]�ӎ�v
O���R�F�7d������̜`��V�t^6ɥ��[��X]F#��1�q�9�d��;v)��;&)$�`U�Tد�$w���*��lJ��ܡ + CN�n2s�+���4l�ՠ<Fl$p΃z��+M[ǈ{cls��K�q�'<Ș�X"b�:F��{W���qzm����G�&��az�6�譐�s0�
u��jd�a�6�:1��|9įXꋥ��Rb�_Oj�+���ܥwpv�ԃ�c�vv�	�<tٙ�m+�:l���]�u���������O�Ǭ�s^}? }���%W�ƌ�h��Z���a��ĦF���-�[��Eb*����-L�խ��1X(*,���EUq�**̦8�&%qmıjQr�K�.��mY��S.Lִֻ�QJ��4���*Vf\iYQJ��b-T̸�Ae���\s3Z�3Bh�zn4[���DT�*�Rۘ�1hѨ�3,�m���[V�*�k���sV�S�5mj)KV�ᒷ0m���8�EZ�X�ba�kDkZ�ڔ�:n�ާb��eV�Z�q���TAB�X��V�c��c��Kf��kZ��ed��KQ����
\�E���TD�G+G+u�Z�]c��L�+�-c�\�%F��i�q�\E�ۉr�mZ�Ҩ�Q���m�R�)�ֵ�j�-+��-�e.W
.%m
�D���F�Q���K�\�ۘe�eh�J.5̴�P��\0R�V"�+q�+Z�s0-�K��\Z��V�Z��Eq��1Uq���+YXQ�����eDqe��z���7�ѯ:9]�{0�yF��u�c���k'k�r�J�f�KqKc5Z�+�i��+��+U���� � E�"�E�I$Y 	�}��s�5�z&����c:���B��V������zk&L�s�;�lƷ5"�j�*�g�I��ć�d.����]u�<��,�"��5�T�j�n�K�Xѓ�*W������n-��Y뽵��<��:�cyL\ͨ��.ی�g�k,����ʷ;ϣ*/����l-[
�}�lN����t�Ǵzn���ȜI/j�VX��B�:�s�["�,��c�.l�|�C]]�{%��16L>3��'��ͺ}�ϗ�x�����Z����k���4}:dC����t}�d�Pf�Q�?�캕�.�7X�N��I̺�b�vD�W����U�S��sh�(i��5r籮+'ꖆ��� ��T.)�b{g�NϽ�v�dy�Bߘ8F�	+�[�����My}K�K���-�����nc�-�񱏥�춥���22���N�"Z�!�N��2�<��K���N$�}2S	�������
��gT���Rz�Xg^Q�pJA��N�G��P�Pb����kB)��F��~s�;�;�$'䄋 �E�"���A` �	/�y�_}��.�����[�z��y\r;ؾA��}u���e�z��|1@|�*5(:��?=`�g�Jʩć�v�pP'7��Oz�'Al�w?r�z�Q�u(�H��S��b��yχJ���M���P�_8��h-��O���0��ܽ�x��j�k=��*k8�:�B��|s0E(�U+��)�b�4��n�F��[�EA`_?i��ޑR5�yeD	�W�eT^�ʸ� \co%w�[d�m�J�[��m�.�Q��dh�N�_W������ޅw5I�1-����S�QWe�ОW΁f�JO�y��o7G���\=㫽�Ś�-�n���]=+u*�Ŏ���4��s���	�R+�O�ٟ���7�y��.��x��_�ʕu�v��)�z-�-�%���s:#x�����G�2]���K��iq��"��E=蛔/gWwR�,�����r������Wqڇo-�K��}��~���?HE�"��$XB) �ҟ=��.��2d���R}X���j���n�34{:���Xy_�����$�Og�w�5iKԃ�O/4�Tcv�囱{��i��G@�?�(G@�gi�N:q۔(��\�w�&R�kT��t�X�/W�R��,9c�$� ��Smf�S���mg^�J�M��?����/ �K����3����^�^�kF?��W��Ou�C�d�=�b��;9��*�(���*�zp�U=h�(g۩@ǹA�cT�
Ӱ�.�A�x'(h�:\y�fk�lm�OY��P�	v|m&%J��]�OU�."� ;=���(���3.�:ը�]�R_OqPd4 5�ДuAɰg'T	�����|*�1ۢ�6𸕝�>T��[���Ť�۵�sy�O4}Pzb�]Wf���u���RC�M=�o�D�W�$���lR�oD�8��Ӡ�mSVot�j�Zý�v�%�\YB3D�N�U���9�А��H�Y(B)$������|o�s~���٬��.�3aq}4ۃ����x�E*NfQ�������Dz�>&ʺ)=�X�Tؠ��E�R�w/Iд��qDZ�׆h5��,��楬���L���A�ĹE��(����}��y��f�|r���RO��(�����:ը�w*Y���m�P�s���X	������)=�ef�
�lH�㒣e�bk3�^)�:����%Q������Q�}Qo�l
�~�b�o��[Ws�V�ܧ����T����W0��m��u��O�3������u�HY�����1M���-Ey
����ħ4��������D����GG[Y�(S�O������$��>g�c��b\yNr�E��L�9�qY���� b6�;h����44uqŚ�Q���J�If�Q�R}���YP��}r_92����3�������+��p>��4l���N�ڐ�aN�>8,m��F�8j�0�7�n��7MR�:U�i�ZhMα��E�wO��W����@�"�RI  !'љ����X���~���*�++M�S�b=,�F�k"�*ci�o\�\�*�x��K5M�2.����I
�N1��8���؉U*6+����0)HqB$q��@�q���L�K�F�� ��VO6�'��H����9T�.�{�*#>nA3��Ht���M����B�]K���vk�����p(�v�Jn�k�f(�u�%�U��%D�`b'�	���aĖ�&N��Cr�b]<�۬�8�ǫ(�cJ�.�0V��[sE=�,����2DJ��E�9�
O\9�̈́���s,ti�lTo!��~+���8*7~A�(xM�hxi0/7u0�ħ�i�(�t
,�r�)��Q0el�SQY.��I�rʗ��M:|��ʚ�Q�XS�l�t���ӭ:�b~��t�q-1CN)w3݇1�OV�m_ZV`\v�F8U���u�۔h��ɰ��ئ���^�~̰������E������^]wb�+[�ۼqi��|�`#��#�{tט7�{y%��&�;���3{$�b[�}^��F�t�*f� [�`Yk�E��E�Y:Z��-�����a�]�|��s����*�r}�]\!��K��ԖO9��У��i�Z��OZ�wy���~s���	�	a$P(!H@3�k�ީs��ۂD�S�Hۅ�$~���p�=#�� �΅@P�c����1��l��g.�hHx�&YF�#�ܨ�"Le�>f��i�3p1��K
7F�X<V�T�/ӟX�'��W�t2��E�F}<�	Kʸyb�ڍ��oA���SN�6�OK������B#(�Dk���J)�.��/L;��4�ּ��sw�W��"�|Y�O����Ř�TA8A"�Q�.��\		Ky��o�o���/^��J�r�(�<��p����&���F�[z��z^�wT�%h����т��{�Y��z!��Ĩ���b�����;#�t���E*G	T ��=㇕x���H	Ppb�"��}^�K�<�4I��/�]7�A��K�XX=�\�tX8��7}3�B ��x"{��w�r!��u�U!���L1��mt�}�Y�/�"�eģ����]�D(�t��f�ۙ�0��b2�z[5}Mt�a����u���_]��w�|h��4pV�g�d��k�9:��y�[�|���湚�9��?0�,$@�� P,�� �x���wt��7z:���%2;�(�T$�Xe��t��e8wTȲ}�5Q��q�[��Y��Z*UD�NY�xA.�����H�ְ:&Ǽ�.�Jyt9�x�Sb�Y�����q����[}���"�<�o��>�	���������sE9�h�SƭK$�E��8��c�8�*��L]k5u:�giNu,#�3Q� �3���nYW��."��YV�K%��W-yU�u�'���D�+/�J¡D]/��9��|O~^�)F��L���i>�Қ��J<i��i�p�H�5(�A�+U?'X|�A���צ��.���o3�.3�O��I*e�1ب�h�x��L�N���FM�#�P���L��t���7�mET_��r//�D���QїV�`���:Z=���y��{y5�$<h�G��e3��!?��ռ���o�x�j�����Ѳ��J��=����܃�-�n�]j���:,tJ2�)�CEn-��h�����AN:��)}}\�*�듣���S�j�j]vWv�,����b���+�:���FLɼ﭅*f�{�'�y�{�~s��@��AI P�Id, � g\��s����θwaP�L(T2����b�t�����@����ӏ����a("} �!pih�t��~Z��T��Vl���.�҆�M�{7��u�W�����"L����Bhi3�:#w�*�d"1�FP�/{��满q�b�����2������P��@DQ��F�8gQ�����^RQ�UL��$����I�E�J�,��Y��z��ՙ��D�z��p�ў���i�#o'HA�ٛάm9Qt3u� �n�u�c������G�h�o�hu��b�����e�t���E�I��/kFd�5mi�M#ӧ.��{`e����
���+%�t���ߴ�x�v��N��8k<�d�)w��ɞP��{3�$��P#dS�M��q
��3�9�����ҫ�����N%�����cާ�Ү�#b�>���:'�d`Ir�+�V'�˻�5lyT����<nuu�^teV	�#u�0�����{�L4����މ�ү�w8�	1O^���KCԤ9��'5�lE̊3n��$�֮ö�(����5[��w|�9�Z�?�@?2I �H��,$�@�[��}�~�z�>�$g�WDP��wЋ)�x���nٜ��*Dq.=������u�2����L֊�;��g�q�����L�ʫ%�ۯ�����~~}6��i��r����o���:5��Q��_(�:޾��0J��^m?%��)��{��� K�=�ύMҿ�}3�Pھ�h���5����{�Kz�{���x�EFq���_hE��uq���f�4��6F\ӅP*��u;��,z0�������&x"��#�K��6*4���G�Nt�C͋��z�x}"��,�����#3���A!d��Ȋ����Y3w�*R	��X�F�����9�,��f�J�p�����n�E!\�y�/��\ׇO���}D5"��.�q1P�7�L��c����|�A����8��9Y�^�p}�4}y6?T� �G&Q�{J�-��r��v�B�i��)T�m�mU�y����dw���X���t���(Hx��+v�0��j���&��*�N��A)X�W/�O_r�6[0�Bth����
�(�t�Ϫ���
���0�,�!d�, >�/_�{���0?^N������W���͉� >�p3 �.'�h�o2x��5ϡ�d4��p�.�r,�RȬ���ߵ�B����Eb7�T�=F�� ,,��kf��'�z�X7���M�Գ���ՄP{��+�q�TH������4��-��@��|�R�C�`!�f$�Q�_mqf�.w�.��G>x�dڻå�Z��衂o^����Jj���Ζm�*r�����Ӕ�V�NNi��QF��Wopnu^�e�)���*��~�t_��(�QСTz��l�ᆰq��3�����G"�����B���t"š�O7�����|,S�����Uix�2�)\��~NXc[�B��Jd���N��|s��k_f��g^v4��TlC��P��K1],�b�U��R�1�tA���)���m�}z�[�����Z���m�8*/b�V���y��S������9UW+睊>�K����b��Y�����eo��_��b�^��d��Jջ��2����f<�Wtn�x댮��A��H�6a�{2��m�h
�"9�mQW.n�0�䊦�����{�V���-U����tIK[Z6��/JQ��Z��6oP��wS�pT�厰NLԮ˝]���u5�]&�
�h�W��I3���u�cKh��t�p�ӸB�P���|��gdq_�h���a����&�:���� ����/��wa��'iॎ��P�>k\Md]�N��� �wc5z!�k�9����C��f���7C�્s�`��]�Z֞�۾=�����-�U݆-A*��x+�߳I�5���4;�h�^t�Xu}�S��]:�;yM%*<[,j��l���}����l^oj�*�$��9.������:��a��M̀^D�\�&oZ���!w�06@z�Mw����8��U˻u?��=�n*�Y��}�u:\j)��
[�7��8�9��!�6ȏ�W}҃�i.�6�K�
��R�S�:Ιi:㋨��1���r=����ܦ��p�gU�d*O\��8�X0�u��
�i���=[������Z�,1�]i�{��w~3� ?���I�h4~$	
�(�2��I�'a���(��wVQ�=l=�@��=t^�z���M�������K:娗1�O7�S�9ʙ��V�.��u˛[0�#�1�v�Т�rm�4�f�n�*���7��-�ej�B�Ldk�Q.�N�dp9a��VDeֹ�)̩V��tR�� J*��+U�Wff�<�7o{)Z��F���(U�vq��`Tg�׌��������[������5W]�m�b�Om��A��t�TyE��E��T�i����G4c�Y#2��=n�j��w�(9r�-�\A��쮀`�ȶ�W_1�Fx�FZk��7w��@�ȎR�+�9�K>�^1��λE�.W��n���]=��k��pU�A4�U��J�Yoz�:Q�V6fZD�C��uu)nV+B�re��f��1�����B�q}�L���-��m�� ����'�[��<|����{�u�Y@P�\�����7��s雘�ZU��ц�N^Xv�yah�O.�U��n�d[ݲΠ�a�z�R�W���Ӭ���M�+3�ce��99����ܫ�2>�Q��E]�*���(�3�t���wF� Π���7�UT�B�`%���yr�`3E�0Ź�""�mIZ#Z�&J��K2�[R�̶���U�=��h�������Ɩ�C1���Į-�֕�esB���b�V�b�3*���m�mP�����ֵ���2��r�i��8ƍe�*�E���f6��ŎR�3)p�-�e�ak�S0�sY�kZ�[m�p�P�#�j�Z�VQ��)[Zc�	�3.eJܴqq̣m�e�ֵ�&���cی31L��2Z�-�����\E��P��1-�jcU��1S*浭j�jc2��
�G,�FL[B��Ķ��*��1����3Zִ���T,cZQĹJ��%I��F��[��k�3*���ֵ޴�]
�m�h1�EU1r�S33�Y���2����mJѕ��A13-ֵ�"MJ#Z����kY\�1G)\��e��8\C32��֍�,��E�&"U-���֍m�r̶�
�#Z�m1[�T�����30ʶ�m��s(��$L} ��J@��W�5��im�!���ck�V[.Wu�љњ���{;׽!]�"�.&�]�]���Nji��lU$@d d$UdV!&����9׼��=��gR��B�}�+]:\�w�.U����O�n�x���f�+r�^U-	�9(u��Q��Q$D��Y��ld�5�K3�:b����v�.lks�0<5�.*�Ra�Ix]u����x�Qp�~:=e:��rG���3��~� ���=r�֛A��x	�Ȯr(�x��,�#���}�rލZp�`d��l�Cr����׵�W�����r��~7~U���Y�Yy�<�m.I^Owa��Н��~�.,���D�O��oӧ�b➉��m`�tq/�R��Xܼ��rz�� ��Al������LY��ָ�;��)��X�`}<h�u�V!ф�B�4�nX43e�k#JF1@}�v2�^�9�1Ri��%��`ɇ����Q���F�&�l�(��qT�*��V~�L�۹����ll���#��W�5��V��j};��
G.C<7���R�ɣ.</
lh�hH�l�����a��
n�fF5�&�0J���z1�c�F���G8��<֯��T�(gP=mq��so��K���Vyn��V��L��&�帯��z�b����i\������
�E!"���I$P!5��Y��~��.�θ4 ��X��`\Y��Q����6��O��-����s	��m��%	Ô��&�;�N�}j�O~
)�tN�,��OGp�s��z5n��Ut�(`��ǧh<;nlj����E����,���"���Vm}|��*���,F�9g��B:Y0�."/�����w��>|�4$�R�ŗ��g�w�2�%�Df�x�bT�E����O��h��-	(�	�����]△�J�l� .I�&B�Oz��/�D�<2!���߲W�K�

���V�ꈃ8�Y�o��@k���ԝef��bKi��p��׋��Tw����虈;�Аw�N��<�:��/μ)�G��k%���zBsZ���IY�o�H�s(���ʇ���D�\|J��/���<,�c9d\��7
��6�l��?YOWeu�b���ܷ��u�|K���^o{)Y�I:Գ�Y=��Vp�h�vuԾ��eJ�wk��3/M���0[0�~�7�~�zn��0Լk�dI�F�n辮��:��j'|(��jZ�*]�r��W.WN��j۾x�s��^p���� ��H,!�B
HE��E�B��k߽�~�|y_ƴLU�Пե��M�3���|2,�L��qx�h!'E35Px��(Wѳ}8,sk��j���d(~��%�VѬ���xoK.,�1/3Vo{��.�4C�6Q�]�/zp�}J����'�ڦnbH@��t��&�۽�m�UqcUŔ_)�8��ǆ�V8�
����,�SX"
z�TϪ�+;�yٱ�*p�� ���[X�x�h5,Ҍ�iJ3��7�+����W�x�)�WvPi`��(
�g ���J�FO+��O5p��G�b��v�d�rC��W�\�t�O���:S[���8�։�3%�U����~|r�[�ԇlqcfI�����	�tB�9p����ZȮ�ŉ�r��Wj�i��}:���CT]x�
__|�q�����O���l,x�ļ�oj�n�7:C�v���˹�d2Y����g�~�$:��x�$l�C�:{��E3��N|][��,�B;@B�5]�f7��:���&�<���r�)�����M��ɛ��x.{���9��Qm=��r�����p��e>�9�2��3�_]s
A9���Z�?I	��`a �Y$�,	'{��{�Ͽk�s����s�ev��5f�+�pe.�����Z_yxm
b�z9�����ȝ��;�o)k�#�,OK5�Y�Q3a���$*�,�31��0h\pӹ8���4C<�U�h�.�*�ʶQ��DWQ�cu�v̻�9K9�场LC�Qe�r��>�2+"�C6k��lI��>,8%���P�c+�|����$C�l�����Q5�7&�f�70b�F���x	킗��]�yg\�k�R�i���J�đ&���Eg�
O�+�����_�q�ɰ�(T�-����sg�<l��ȥ�Kb��9�5D���������<*�_�7\�,�U*��q���l�1GDWG�v���˘X�dһ����+��w4ڍˉ���E��#cI�J%��`T/���!�j>���rέ�S��<���r�Fȷ�N��&�+G<�O'��T��}u��U]�u�Ndv��1
k�U��ǫ;���d��]�S�L���@�^�m�v�޴m̒�q�ZEi�}l�b��&�:@̵ָ��7�v,���W��q�Jc����Y�r�ʘ��rP�L�Y�aQ���m-������P�@(A`�C˝���{�v$��'#���@@�����t`7�N���r���6G�+
�Ơ����ogg2���(�C5q�Y[��(�*B� E��"9EY�b��M>�����wd,{��)��펤d_K,ئ�̔Y���� ���$�	���o]R�ї�MT����'�W���Ĵ?��Tz�x�US�5���/��<���#�U�Tg&0m�ËUa/�jq���*��(���=�D�ywv�=n��t���"^V�Y���ƛ�ס�z4���_F�yw�ܺk�;y��뀠ç."�f��})-3�o�0ǇtP�$�϶����>^���o�X�(p� �QA�CZl4"z�Ƞ9Ț����쭿e����޵�+ӽ|p�b�����0g�\E&�3}8a��#d�Q��`�)=��l���6�l��aŌ��\*GK���}�Ӆ�6<�\S�0p���������dBwo�Nwz�gM�÷^fxѮ������sa{��x��������|�T�uޚN���oW�i�����_uuiq��1�%�YW�I���j38�N[}e�����8�ߝ��~��`�B)���"��<׼��~�:�/}?��yױ=��` s &h��E}�6k��v���\w���:y�J�o�ᕮ�X&xѡ�xچ��MdiH�!���>S��ֵ�w5s�����S�2*�?@��xJX��Y��8��p��;W�,���"r�-ދZ�TSzٳ�L��Ⱥ������h�%��s԰9���=����A36E'���Gg��mx���xcqH��(�g��U�@�����j ��2��.)实����Ϊ���7�h��LʕL�c�Z�Y�P,v�B��Q������_a%�"��x���,�T���5�ο���p]�a��W��RY�d��w���six3kE��xS��X�|BO�z5B#k���suj�R�m_G7���w�#b�r�&�DlkLaY�F���eA�d�IϦ��3��N����,�:<c �A��3�*"�}iZB<;�d,0K~��<)Ga:�B�٘e��ɿh�3��:�Rk������N�lU�HǸ
�J�mȳy:�S�P^I[Ϩ_J�\�'��v#��R��o�ZP�WL�m�)ํ^�� �svz�c���>��U}�W�!�,��E	���j�ݽ���"�~�f��:d�x��N��V��4�[�#��BH���[B�(�^�ATk�0#˃��(�Pt!eAf�T鞃�.�s�ݾ���,�lî���eW���FE9�g�D!�|Kؼ�k �ׅt��g`�8�
c�u��Ġ�4�|�5�N�t ���}�O�且nY�˙;��{�yb�k�*��!3���V<r�{��t��M��p�;&^���|�-�5C
�!(÷R��_>�5��x?�Z+���5�~��ċܭg��.�|�eD�7p��g�*�S��*͆߳��������ʈ�W���%��z"�z�niN���<�SzjU'X_�ג�\�:%w���v_�v��;�>�Ϣ�e�Dnt��>�h��:^E[�h˩eK�p�'��8QV�Y=s��e�q#�DWE}qǭ�S���#aL��$�������d4k0]���`�����V[KB�k���ɭ��:~%���.�=�v$i����m�JѱܢѨuJ'5r���-n���Q�pq���Y�Pɑ��]kkOJĉ�e�ݵJn�o���y�� x���H  	 �E �wϷ�����LG�ͮ6>t%P�^�"��S�@h�u�:5LEmS ��sv��k�̘4�1�k��VJz�D��hZ�k���3�wot)�Y�{�Ǣ��?���^��W
���6M%�[z� �f�0];�U���ש6�q,��FCTC6p�f�2̊,�5HR��8?���qq���Չ��������;,�l����0�(ߢ�@�2޾�<���sd�7=:_V�=�5 �:x8G�A�v��
Ar����e	��{m���Q�z��g���U�X�tk!�ւ��r>��}`U���t��+W������ӜK˷v��1�ه���Ǎ|8F�J8@��|%B���lxz��fQJ{Qۓ@9�lQt�5�}�a ��h{�fx�?��f*o�iN����/���N�np�R�_�"�4�RȬ�[���!}�1�JG��}���ѐ-]h��mU�Q����2�yҶ��sۨj�吡Ą`�vyd�t���n��(�B���	>�Joq�Wi����E=۾��\z��o��LD	������}3���N�sO�^��9�s:�7����d"�"�> > ���$����7kG�fx�N(�<:�9Gڥ�4��c2VE[O�J�0*���e�3j�K�u��X�d3TС��g�	��1GEuqf��t����>��j�y��PC��d��h𞣣>�@V��w����*��[n�}Yq���nA͕؆�[u��� P���6�i���΋g�̜��>4/e��h�)u�i��A�z����wu���xۆR��\xT4]'�T6����(����#8��k_R�k/zv\�½I�F~�������f�>~�+����@jmۇ']�������\_�-B7J}�ށ}�*f�<|v��2l��H�Dk�I"�F\�\ɩZ�9k�\���Z��ɳ�٘]._`���Q𝉅KWG[�jQ�S�9��q$��R�Dk�Z1�yS"*�<�D�BT��JD��ӳ7x��WJ$:�fKA��O\�0D�s�l7��p'�p�=B�E]��K>פ�S�u߀�!���:�k�:����-�Ս|Y '�hJ��"�C9���R�����R�V��,O��k���#e.d�#�K����W?>b�Lc�����3u��mjY�| ��~ ��,"�(���^�������pМ�!A�*#�P���!:����R"�Yύf��S`��]ws���t2�8����0�"~ZeɊe���Mt�`L^Es�f76�!�k�v�j�_�P`��$����G���fk�ym��#���c��{��)�߭_���V:���U�A�<}P౬�0���8A+��qxq����Δ���A�3�=�7Ԉxtx��S�:~�]A՚����4ƣ����G�������^��QOdYA��Ύ/��<��t�_��:<I��G><3=�����:�-�v�f�E˦*�q�^��_{���JB����[,���Z��f��م[��=*�a����[�̜:t�
a=U��D�(Q�G8̣���*��)^W����r���P�[�!��Ⴣ�=���אo�x@��	F���|Mz+�#苺��w+�C���P�J�\�Y\xO|�x�Us����xyCp������G��	yϦ��f���PV�T��1���ϸe
��.0"f/m%&e,;����V���ǎ�:MNg<�	:�u;M����;>���T����"Z��������|y��G;��VN�Zک�iLG�g.mꛙ]��0�!�+\�Wp�8F�X,ެ�bݏ�r���#����["��v˶"I�0�\�����K;���l���r2�SJ�
k沣�2�������-���D���ǈ�mH��:�H������z�x�;�h�E�/���oy�Rr}2֗zj&����o ����r�X�GQ���uv
�q�m|P3�B �;�!�@[u-��+��3��ѩu]mr\��K��J���Κ/.����ݕ��;z�M
`�{�X���qj�3��ؠ�7�b��u�䵼�}g�i��T���A�
�Л�5�S7-ep��Pèk� ���V����P�"C��Zx5�P�����V�r°�`>;<:9���mf���F;Oid�lWR�[��M.*�c~C����> �ߺk�]�KC�i��g�V�En�d�����R�(��W.�d��e��{�RP9�3�q����{e�fg"��܏B��:��;�ǻ�o��@F��;���)$�� �J�'��η}&�z`�)�_Ǡ��q�^.B>��9vU���^5rVMQ��3��
]8�jST5K��4-S�d���[�9\�]�H��φ5��;����L{�S �ו�`z.��"Ʊ��4�=��+�yݤXȁ�P�#��蜕�ԉ}v7];��	��>��Z�+��\Sv�@)s���N�]����o\�Ȧ�ݼ)��ܧf�����U��iIӆWtI¦�z�7�L�WG�JYAV����[�9��U8l�h�*��h��7��W�C(���K�j���D�sp�3_s���Yr��SVj�>�єS$`80o�v�$�۷]fӧ|��2�.�D��+�"Rs�ަb�3 �r'ǖ�����%�[�jÅ3K:���#�inJT�`];�q
�q��L X��i5r��`�ȿ���2Rnv�Y}�g5�˦�ü���u���;�hZ�Nf9=����t�U&*���}^]s�����G�G�Y��H���,�\��V�wv�3m��H�&(�C�t����iYֈ�|p�>���3�,kx�[#���k�+�!�H7-w�%n�'CKC�o��#g��9��V\�y��!������a��J�<�ps��nS��Ws2���b�ġfR�iTRč�S2�-�-�$R6�-�u�ޫesR�W)���-Z�-�r�e3�[��Eq)Zbb0�n岕�Z֎��Z��"�2�(��[F�a[j����`��m�E
5��Y�6%j\ֵ�Ճn8��R��c��.+J�3.0��%j�L�`���eF�ۙa�ֵ�z��j#qhcrⱖ�ife�eq�h,��ѣ*�W�c*fck]�ua��U�-ˉ���pf%���Lk��S32�l��%)�`���jbȮkZֈꪚV���*5U�Z#��bR4���8��(5h(����R�����i�W2�2�kZևT�k5�-�T1X`�kR�)K*��pJJ[��qX���Z�B��m�c
�Ҏ7,*�D�E���aV�UeH�b��R�Zڊ+h����mG(����+B�U�bʍ����6o���_s�>��j�%��m@p����']��7��~.ܮ��w{���0.ߵwm(��R�k�d�w����	dAb�w���׺=7H�GJ �0t���aV��٧6���QP����C����e��]x�R�/�e�Ƅ)G B"NF��3��b�x�򤯲ߕAA{�[��O��m�X��j.�h������,{�O��D8�jt�s��vfB46�
����{�2)���'V/�ٕq�G��
4/劂��m,'��|o���\&�'ދm�!!���;�'p��P���]�e�]�L(�	Bhi3�:#!��jGm����i�Ҹ7(�HG�f-z`Ĉdd�f�d�1_z� ��,Ա��HS��$d��E��W�t�&N7+ M�dP꙱�D�+� ���L(��
��^3���0�'n���<hC+O�f�u�f����<�!��_s�qZ]l5�j;Sn��w�n}�3�&�p�L��S���Ƕc�p�J����㥭��ae�`j��ڛnt���Α�
�?\|�����|���`ݜs��W�%��4R�u;��H}�.�Ċє�����MbXt�v,�bs��Æ�����l[nou�I����;��������%�������8��]M-�s7G�g��8�s�޻�?B~B)�Ƞ) ��$}��o=˝G�oի�L�?��<\^��0�V�\2�,�
Q�؇�7:���'����4�y�{iF��N��t8��,�r����Mmq���ً�\��TN��K4���^.�K7�Lw@��	�@6����C:Y��W��l�o��ӯA�L��ڀ�E�o�C�t��$�]JKG�"�]#�X��=Ns�ž�O�1j�`���5�Ծ�06!�ԍ���s�,L��Z�F�+Z�}�_�f��p��.|=�g=��w�L��*�'�D��QNΜ!
�ZJ���Z��qaE�~�9֭X�[\i�W�*ZE�J���F��hN���L[8w��<=��~<9�_z4��ψ��y�28+V�Hx���V��d���F�aKS�Ձ��UR�x9k�^�:5��P��q��T�_`�T]X��ţs���QJ<�v!S�Ȭ�Pp͓��'1�8`�yN��Ϸ�|0�4
\�V���[S�|�"�Ew���tُLئ��E�v�5	�*��j�n7@$&�e��tξHtU�����/o�l�LS��L�gy��h̝�L"��մoP���Īo4j�8�oŖ��Q3%>T��obܼ�w������s�����)B)"�
9Ӌ��{9Fc��F1��#����R���ʏB�� Q$-��C*���u�$0[1 70�b(4fxa�����������&=!�������{7��-ӆ�$�s$D��D��e���A�7%�g���1H��fX"3���kJ�w��YՇA��x��1�j��Ͻ�늽T2��Q0^l�]��<��z�;�JT<��@]N�$���(�Se�R��ϵn��n��H�М����CX!���+�ӭw�
nz�dv�G��G)���Tm�i���ܞ[�FUM+�qgM�bQdM��­�#�l�c4��iQ������������Z�<s�
�.�;��ܶ.�Z88��J��z�1�o�U�� )��C�,V��~�K�.�u�E�TOCt%,U���|"���=�V5ӯ|�(Ï'��X��5�[�7�E�Ү��
�]s�_҅Y��Y�$�D�����@T/h�_i�Z�5m�H-��[��1�����]\�LUN�d���u�
�xN�3]s�]�s��;o{���~s�9�C�H�
 ��H, O�|	}�K����j�8�s<W�8�o�e죷�|Y��њ�Y��Dy�݃w�aJ���e)��,��:]����:��ONL�'�T�<)}�oB�L*}j���7;�x���u$�6��G�Jt`�[l�|k	K�V���o{��<�<��Ǩg���g«łϡ�"l�:Q��~y$���Gv�mr��Z��*�9B���nW���������u-|�o�m�^���{�)}��Z���އ��7���s�IL91��@��A�A�	H�#�y�#��L�uJ����l�6� <�p!{ߟ�g�PM}�Pc�*	>p��[]��(U��ndN/ڪ�o�>����O�A�5�'�����)������y����Q��(/#N}���,���c�0g����T%�&��}��%��{�la�'���N���z*�Ε�N}�xۆ�~�4{���_��L�5��
1�W8����U�yc��lX'^n�_+��`��Wǲo1JV��������g	YS-����_��ײ��|@�2�v��yr�ܼ�0_%ӧ[�%�J�s6�]�ڶ�+� �~ � |Y�AdH,I!�{�^o�~�w����9�8{=u�Vr��B.��BYA^���A�����"�嚰�efv�o!ŋ'�i�~X<�߃�������]t�Y+];�D:	�I^vs��������&��_���������c�%��L�(��b��o޼�̮������tB6;Ӟ�^�VdB��mu����.�*.D���'��Ǻ�X=AP�.� <!??���E��͍R3�i7�������S���[��G1�(����2�㰧OE�DQ$qAٯ	VsA�&	�(�vf9tI��I�ukP9�4)�����߈����T���2\/�9g��x\��^�ӻ�:X�e�Μ�@�)� ���:鴰����ߖ�'���{�򇖖I]L(�w�D�D̲���x��x�V����<U�Q��g��{8E��I�>~z/�
�B*�"
�]Dq��J5�g�*,z����W`�dz�.�8��s�����N�g�fo_cRb�
JaڲZi�4��gwg>����+�gS�����G�s�xU���N��y�L�1����Y֟]�/��[oc�/3���2�^r����oN�}���`E���E X
L����{�r����0��F�l�3��n꙰�h�E(��L(����ޅ��歔�GQ��0Y��8d�������G�(dY8�Q��}�4����saqb�H-U�|Mv��$F""�F�����XlL3��7{��7:SNߞ���E���������<
}#l_�&�G��16�w��-�9q
�ɫ�]Z���czYp��ϻ%�*�{8b�*��8I��gG՝o"J/~��"(Q�x�!É�)| ����",:���t�YC�z�eM�<�Vt��@4]�A��{K�;���V�nt��"�PΡ�Uy"�]�{��u~��Q�gc��G��#�J�B�&��O��~2�S^7�y�'b.��Z�ٔ0�U_+DH��g��(�K����:S[������7/���i��.��(�0�E�ߠ&0N�nUq؃JY߱�!�]��"W9b�o�;��$)uI��x���K�nݏQ�+{��x�6Һ�ۉ9��%�f���ϦP"�g+j�p�c�fF�h���Yx�u��b=V��m����U�a��ΫO�����/���%��pj�k��L^.�0l4�.��]z'K*�V��JL��$s�u��������rE߿X+�]x).����J5l�rՁ�9O����pՄ�WY)�d�s���ꜰp�f�ixT$��Ι�*Q�n��^En�{]�Ӽ\l���K���vR"��TN��dWM#&�#T#>�B���t���"��d�����+�ZM�j�YkE���Ya���$%��c�Q�j�W����;��xe���Y�2��\"�DeFLh!CX}�x+�@.�6���L+'�^��7� +]�y��w���B���G:J�.�?.�n�Z`���|��3W����#Y҃�^t�3ԑ����n`Ć�ܔsa����j�gI���ʙ]#_�&���h�o2Yv�������Y}	�SȮR.^�0^c+lUa8�;����B&��0�(�'�`�6�Y�\\`�p�R�5�sdPY��*��C"!nygKs���+���X��TxP�B�'=��F�P��:;]iF:z����g&���}�\��Xe�΄N�:x6<����Y���Wb��A���R��2�ߖ>ԝ��½[�������=.��$�ǥ�F��pMm-\�
�R�����5��h�k:Eϛ�ӝ�t+��Ĵ{�}m���n}p7(w�%�����Y}���&s�Kp3b��@�;C6D���4pDqGm�F�(��=8�"�Åӻݭj�A7��	��="5 >��%�'+ǅ\��C*��@� ��g{�}��9oK���,W�z����:��o�o��%O�s����c-������i8�]H乄��0�2�9�Z�^�R3�p�yVf�a}�.��Mf�w�5"2	c6�2>��]\��\����#����J"���i�so���wl4��FCR�H�IfP�
��Er(=Fq�_]2YV��)^l9��r�y��+�y���帑R�`ԱT̀�h�]�EX�.�e��*~�Y��rɣ]�=�B��=��u����>�h�1��G
�
����t�Jd�h��'�9%l0^�D��/ }�u�^�+�r�Չ��ӽ����#Wm����u�i���Z���`�ٷu�m�����Z ���4�8�f�ƐK
\��:;ۊv� Mvl�{�;;�t0:���u��f����&ͽ�
���2�o�g)ߪ�{9�M�ʭQ�ɢ\D�#�dQ�:I|<���e�����}O3�ǋ6�)�O����."����bS��*�����(��\*z]D�	�)U#��{y����<��Q�D��������b��#�!���GH�#"�㍦2f�����f,���\`ݖf��E�/f�	�"�}�xչ`��$�ۆ�u;W��l��r�Y	���2�BΡ�W#���zv᜞�<�r�Ǽ�ö]-=B�����/��'>��R ��nxe2�U~��c�X����Q����A{��⇺��|LǄ^� �V������< w��E����N9��4H*��ɊSC�r�#�0w�}��O���^"�v��ST�݉�1�����g%F�ŀ�p2!Βj#��>��m�5��uhU{>�|)t�vT�&��o{ޗ�LW�Î��>��r��\��V<%Px|��|�� ;K��bnc6k���V��8n�Rc�+�<ry؀�x�Ok��\2s"�(�Z�0>��쫣p{�a�u�f��u*�m����	C�:�����{ 2a��Kwz�f���sP!9�7w�5v����o����X����\���.�fT=��#��艗:Q�kA��،z��\g��&�qB��Y��_�(��B�����u]u���h>/���:�ծJ�E�c2Y���ƆFK8c�*�]��4<��%�(����K�+9��ӼX{$TB�2�l�{h��au�0���t.��%��wSn���9
!�*�͆*p��8v���N��z�|tlIb��}7�T�Kf��k��z^q=�Y�f�}�d�!����+ �u�"Gl�s�� oQ�WӯO{��-���ܣ�xc3�E��#�g���������/��ݓ��������8�ä�h��Р�ۛnt�e�������]i���H�9�j?fot�r�p�VZ�f��
l���!
��y9�,���=F!Q캎m�)�W\��bL��o���T8������S�a�����Zf@� *�;�q���Z=孾��<����|�wQ�9��oMM�*��G0�U��%m�	hV�R�im�N���u���M=IE|�7�Y�͑�s���2cZ�s%�@��9�qq�.���(�� ���ê*�	�=P�#�\�FW�u�]�bM��y	Yl����Ӯ 
�5V�g�fJ��ͺ,�B�H:�l���"�*�m�猭l��٪�0޵�N�F�t���}4gG�P8Wً{�λ�vWn�E��i,qlV�#2�Hk;�}s�n��犸_�:��Jp
|vwd��Y�(	kyP�<���Vs���PRe�Ơv�H���(
*�Av�"�`��ШT������4Z�0���k A���y�X*R4�_V"A�����^�gB�f\�z�#x�Z���m���,u4�s�e.�V��e>�.W;w�'[䶏rm�?;Z��KuB
#w��كHT��Y�"�n�M���rh\���oj������s.����WX�u��O.-�b
R� ��Q�q��{d)C�kN.�gcx�h����2���t��:3�Յ�ZN���f�-H�v�U�n��(�Gf�/��u{Ջy=���$�gQ*RM�h4�y�LYˁ��Y�So�rG����-�Rm� fn]J�oP�F΢�&�t,� 
s?����$i�\��F��IB��7^4��X�RV����Ω._M+�D"+�tj��MFX'ZL���iL�#P�Tv��y�M_�����]L�\�5�F�h���A� e�V'yH�c�ݪ2�&U��M��&�D�,�J%K�n�����m:YhjV��p:.�����%�6�mX�@�1� ��~��,� nF�%
1;a�Gb�J�LH6]�8.'����h@.��R��|�LKm:듀��-�J层�6�(����4�ʛ�j��:���_��5z�����Yb��&"��W�ݢi[#�F����GP���+Mf|��M��vJs��)j���e�ñ�csl�L1�J�ohX�ri[/�Uv�|M�K)$/�Q2z*�jBR[.���.���mm�4�M(t	@�n���	�o�F,���fHG�%�Q���uu4ԁ�ѹ���Q�^��k[jЗv-���7X��ij9���,���)f�3o_m%�s�GM������]��N��JZ�ui}�kd�٧ܞf.���([qEZ�����f���ikP���2i�rʄ�d���
��*��(Ķ��F�J$�3�ǝ��H�Ѭ�*[jb��j[DBօ[��e+m�kZֆ�V(�%B�k�h%V�aPR�Q��ֵ�i4�Z$V� ���@kk+���F�j�)UT�1J���w�H��� �Z��T[h�F�+Q���-E+m*�Zڲ�ֵޠ�I[mek)JhڍeX�Qlm����KEU%V��Z�z6ڰ�*
E*J�Ŋ,RV%�iPKTX����KZֵ��d�`���+(��*UB�m���Db
-E
�FЖ�Z�z6��+�
�Km��
��YXVګ�EX�Y*VV���X�P����ԩR��T
��¶��M�[q��=�{��ϝ��z� �:���s�r�.�>jX�v� o>�̴�+!�q�r�Q,�/�iɑ�/C��Y�6T�k�U�����[c1n�n!�|�r`%d�>ήz$Y���x��'�3b��#�4ۮ�^]��5s�侵���hf���ݵގ9�,�B6"�U��8��#�)C#[�5P�*�9t�7S�;R���U���!_�6"�Tͪ�.8؈E�S(��+����I}J;�L%?�K2Ҥl(P���z"����)@C�r"�J�ʙp���Ӯ�-��o"��r��pJZ��G�J��=x"�>��Q3��{U��΍�ꔒ֢���'�qxH��i����-r���I��iCƩz�d]uxĭ��/M��IWNn���5��,��ב���:2Fzp�WV�;?Cs���&!j�ث6z��O:��#������@(u��sDTE�>0l��7�C�.{�j�,j�w,�P�Y�"P�k�Q��Ɏ0w��"@s,���𭠣5�����$MȇpH�'��.�q1���Y�_�#JiS����;�BX�~��^���4�$��g��ѕ8N�门1�/E@���Ӌ�P
���[�n""�o�;+g���R���%��9�����T�������g���1�緁�7���?S�ϧ�2D8�09)�L�Ȇ��J3a��N�I��h
�E(�Y4P9p��8Z�18�,����MH��>�USy׽�����ΙL�9Ƒ>�Y�=A�{<\X�~��s�}�<ɭ�y����3򜯑�� p�^�p{n�����*"�3C�*-R:aWD��\wcw�f���EYc}>4�C&�Wxt�hN�μ�+���>�*g����Du1w1�2wu�<a@ʩ`�.B�x�ގP��J�cz���Y�s(�~�mH�����O�^?9�.�%z�`cx���#B���.��xU˫t3�y@/Z�Jzz�;�򛔵�U�%J-Ӧ��
�5s���%�1�$Z����6�����r}��^Q�҇#�'4����r��3�]��a����f�YFZ�2���~j�\ٜ���O��*�h��P�Z&?>�3������)��������܆�@���Ռ+Nn2����h`���cy˼�ݥl� ����kQ)�V;�╟)���z����5�sp�1v�}wkba��#y�!���yn��I�	��Z>��ȘE�$�(F�K�B
1��.���<�{�w���k9D�z��h�Cq"��0a��q��g���eӳ����@N����.S��OP���'��LB�@;�!A�j\EJL�{�x���k9�Ϣ�3ؒ��|#�\�f�F�p+�\���I�.LSR���upE��E�6�s�wĝ��U{ʓ4<V�� Ci��{�#�0��Z-��;�Q�<��d�As���c�}]�W��ߨS��3Lt>�aq��w���q����?�ȃ�E��M�/>�({d h-��wR�����T��Yk3s����Ǟ��2�1�R���G����2+�0H`{��Ց���g)x�6�f>O�P:�u9ŽCf:��(8�Bia>jc<W�ۀ��L��[�xJ,D`�
f�Ou�ܯ�Sg��l���*��`�'�`�D�b��
S�+���'����w�U�tF���E��j���h�A
Y�ϣ�@&5w�'n�����Ӈ3{��Ȼ�u�;���&(�ݰ�-1�vcr�'"��-��w-���o-i�5�I@��QQz)�*!p��(ټS�^�i{k��]H��y�½}(-���r�����#A�@q*hm�V�q��qōrʽ�
�����Z����o[�����0z��<XI�s�,��� w돮�シs8+��+�J�C���4?\������3�x�:Gc�(����1nT��X��ru�3ǔ7~�A�4`P}A�W��,��.t�b\�~(��0=s���;�f�S\����/�iP�c������u��h:����S�ЅN=��R��|�S�q���_J6NC6<Y���((��:t�wΧ4Gx��U��Pc�S���3��\��8��A�����0x�	�+���90O�_G��G���H<�,�ӟDQ���"9>c2Θ,8!sN��9nosi;�.,���fWL8Y𳃵(-�)|��=���$m%�����)+����y�n?���*5��:������o��!\�=�C�ROxP4�[�t����9;C�t67���6	� Ȍ�w���cL�-\JkthK���ot�f�%�s��,�\W��9��{��g7�j�!�;!��.��UPl����r�"G럜�~��� �9Q~�0g��G��g!ej�'y���k�}tP�ΆIf�r��nm����@>E�ȝ��V�� �=I��B;��@]N��dg�|}�"VK9>���b�H���G-S��{�\] t���,D�:ɮ��ޗ��Þ/*Z�s��<5�X��o*�r����t6�TN��x#�Q�}����]3����:E�u�]����ҖiV_@�ͻfpT�ƕ	�9g�3ŒG�V
�;dPֶ�'�y}�����~�!f�=��ɡ�y[8=BX'����:�
J���9�3_w&��0��4�?Qˍq�d�F�P���$�x��Ё��)}
!��R���v�-j�i]MҎ|=��Ŋ�:͋�r�"_��[ׂ�C!����4��͝�Y���0�t:"�J6��Z�>,t_E	�]���T0!J�遼���ɣ��S�O�Zw�L��ޕ���HNf0pI�V"\T�>�u��z��>��B�N*s3\8�]IiD$�(��M���cC ��Ns2�̲TzF㙽�n����T�]��n3V��kW�)�4ĭ�b�+�X_��8�3ᒼ�SB.Z܋��(�j�%M�D��Y�~� �A)��,'Κ@�T���B�p��Tg2�z3��}�������o�`�@�FY��E�2%	g�B�#p���^;���ұ��&^{���s�i��l���p��Ja��w�&��{G4���m������{�.aa�V��6�*�6P�D�?t�!�F.2�ڑ5�7'�>ӂ-�y��75���G����O��-bchK��{��ڼ�+�"�:�U�9OX�W$9,Z�㢱�L��H�/6�����b#@6�Y��Ū��3fI�|'�*}]X˲�V�Vr�;a�'�����z��B<1�P�=���ӟ^�1��CK�f��i�/�|�8Eڑs�w�Kb0�D�t����Bܒ:��*2m�يqv��U&O����F�����8jq���wh���Wppڪ�1s�ja���ӌ[E^"��ۡ�R��fA��� ��Kk���^�Ky'J�w'���<V�����nkr�6��em��٭qչ[��/��}:���q��-�s���K�Pp��Rӝ�V����twTR`�u=}ѥ�6�C��|Ys�ChF�S�y�`	���:��6�����3����B�S6%�/a#qJ��Dp�lX���R�G�T�o���}��~@�!�قUF^�q�sn�Jx��V5h�5��/\}��9<ӭ殤}�Y�A��sԀ���I5�+�U�T��pA����v#���4��YSv�:T�i�+��0�j�z�Pu%U.TF�\1����:vWA �+.���읆%Hq�P��2;���u��
���!]%��=�k=UD��)�;���?��?�  l�=}YV*Pl� �<L����v���Y~��r���QQU�b1�"OVBq�D�C�T��ԃOW*��������!*z�?;�r_M@FzT#`{&�:Is�K0}�q����y��8uX�k���H������joѿ
z�u��O�A��nǢ��<�a�g�'[��m�L�#lè�ӹv�/�N(�N=�>3λs��/ۭg
��p_<�om"{�r�:�0�\VJ��ه��m=���]���pYyҢnpj��K< �K��N����~���<UNtH���%c�p��)�^xi,g{[]УFQs����4�S�/�H͇#���2&,>K�8=-{ŝN��}~�M���v�k�-�D=�W� +���Cf,'�b���	��Dw�����{��J�E��mB*��e�P�YV1W�Ύ:�Y}�)�{�Nf�������c�����q޹q�:qY� ���c�e9���s�^�Q��X=�>q^�
��B9���c�g����$M|��z��ӽ@#ǘ؝1X�2<	q����D}L뙊�}�����Kx��=/�.�]]�x���S咷�D�5����x��:�GE��5�ɰ��Y��Vs ��{����f3��U��z#���#ğ�>�K�������0OP5a=
��5,�FihU�O�Ϟ�uQ��;a�.�����+z��u��@���ۛ{/8%�	"��r�0Y�1���M{+�/�$�&��@���e��ڵ����������Ob��d�wk�zA1�s��o_n�mF8���
��36��_!��^r� ��������T����,�|%aੑX!�6�L"��,�e�rl��1:ċ:���{uJ�0�D�Pk$+;h>TS��5�B[Ȃ+�h��q��;K�X
F�ƙ�!�eAg����5,�<
�O§Ғ� #�oiuzu�;b��ھ�ǥ}�}D�N� ��"�`��ՇD�Ju���G��>�综�����^F���8�<�(���F>3醄A�@��Di�2����|��� �n�v?� ���c�.��c�tx.8��&�.��Y�ꧾ-G��L&E�dw_���{��V
�U{Q����/��7�˄���(�*�g��l+72�ٰ��kѠ����lLI�P#$S��ޗ��Qg�aM��7���qٳ�
;{t��voMf����f�.�+z��xkfBpgK8�d���ܖ��ڋ�"Ntia�lu�
��wH�H���D�>�#�_��7�«_�d�{d���U��S�s�8<r��k����h�T��v��2�
V�u�X�pfv��%ooَ���b=��w&v��f�%C�Պ�a����NNU�k.�J����վ E���ީTVǆF��9�n��J42g�M�l��ሪ�;�4�!���Z:�V~�7�����D�o>+�ᵉ ����Z��i�ح1p�7P*C�yw���~yv\B�3�?g�Ɔ)�̫�6���#�TxT1wG�+�j��g�<ƺ\��_p|#ȡ��E��7a�37ե�q4���^`B���v��$�{%�wfr�
���/ʐ�>C�ڳ�S;f@�_X�G���daxp�s��\�[��� h�q�>K�WK�g�Ŋ��� ��6�pt/���`�oZ~!�F7#����(7�&bB��k��~OQ2Q�]���n��S��^��
�K��A��E�I2xI���f+qEC��e�fOi�P:XĩKͨ��]���f�|L:á{8uN�G )?/p4�zҞ�A�$�;�9O��{�� ����Z C��IĔg2h�9pT.p�R�&��8Y���� ����|T1`���>�Ή*�z�F��g8��K���x�T:�gֆ�����(`4���^ؾt��-�9����{n!�,���ޫe��R��'{':4��%6�Q�D>��˝K��M�\�~�KR�+dܫ���q����ڭ鶛��J�Q�>m=1�fG��0񈣽P��v��_D�F���Eڝ��o�KM��\�A�I���1 ��+E�|��ڑ���������܍�۵Y�rVܱ�k�'0&��=�l+X�,vq&�Z�e�4WS���h���R�A*1��b�v���q�	]-N쮺����1mj�:⻄K6J�*�	�X�A��U�}v�ڂa��:F�ԫ��^���2�).��]c=����w"Ĵ��L�7�n���*��to8J?Xa��BM�s�h�ұ4�Oy�[5:r'���Vt^��O�M�����ݣ��u��򓘦����RJ�^>��j����N�(jo���wyW:��LGq�9q3�okr�#��T<+�"�"�;ң�WB݌����	���v����DZ�K���s{���q�=ӥ�ղu+Αv࣎h}o2�:�f#vWR�
�Ӡ���T��.]�ӏa��(ľ�ں+;2ޑЗ�c�N���B��Bx��^��g����Ԯ�����C6�0h��V�&@�tа��a[�&t�z�8)�Ә�L�i�YJnVHj�1wZ�j,,�ʈ�L�*�s�}w�SȫGؑ8��l�i���x�Ӭ�9��o�( L������G}0M2��w���DE^��ӭ��F�^�6�LSg4�U���/m��3L��7�!�2s�g/~�Ð@
���b�r�Ѹb���c��lm���]�-��,�P� ņՖu�GV�I��	e�.��h��Q����j�e�z]��uoHL�����
t�X�U��Q�1<�6̒˫�8K�գN���J���Q8٭PG�Yd�ͤ�V#��N^��m�-M�"�)0��y(*]�%kώ���hO���<c55�'�f�
ޙ�(�x� �(�p��c{�`T����%�UN�Q%�3�wO�ؾ���Et&�-Y�)��˷sj��[tI4^+Ugo�\���n���%ֺ�y坥��Cu*F�t���ڷ�Jo�-�m;8��ӳ��۽� �N���K�*y;�k+k�oQ�1l�y5�1�x6C']��<{�M������(}@PS���	QA-�5��*(������.�m�FT�%)b�eH�TJՊ5��R�J�2���D�[�kZѡ���R�����lV�Z��"2����Z���ֵ��j5YZ��P�b��	m�[cj�%k*Ej��-l(��F�Zֻѫil*	R��(��J��6�+V֔QciU��ŭ�%imen��kRibR����-��m����*6ֲ%�*Q�V,�����E%ֵ�h�YVږرJ�����Y�-��Z
V���SZֻҚ�eB�V�شE�JQJ�Ĵ�e�m�V*тђ�FVֵ���j��J��T�ȭ�
��YTR#*%�+�E�KR��6�
Q����J�J�ieIml����}�o��ޟD_�a�&��6�9�Sv�2��-��;m��\�d��Y�s���bz�^%�� ��=~�{9>Ǒ��C+�D���k��6�\���nP5�g���#A�9m]�c�o�O6��=キ�Sج	W���"�x�8j��j�,�`i���@5s3B��2d ��R��0�鯻]in���dd��:X�1]��B�4"�9	�..z㸌��o�"��p�:S�ͷh�)�QFȻ�(V�UX�)amEK�W�u:�K�=��ۗ�dYG*��d@�u���ǅ��q>4r�'Y_��Gf�8�G�`$����o�2�}.Qw��"�H�r1������ݲ��f�gd	`��hk{q.���\����'X/�sL�<aE8eҞ:�V���e��5�I�սVo!b�* �XĒ$��`��@��/��J���f~�ӯxf�u� ؖ���R�> �8]u%	R ����X��Y��͝����j����b��R$9�wKq"�S0a��P8_}3�-+ڬ�;N�G�������E�\3aMnj��O.�e칫�z��u�X��z���,��N�}�8II�Ae:���oWfF���zoSԩłk������-�|Yu
2#:wn�}���O�o�z�nV�c�Q��Ft�p-zp�	B����@�@P�>&���<A��I̒=t������NDMm#F�<p<IZ2P*��A"{��0��9ރ�^m&��報���'�z�vn�ʓ5�io��8 꿣������a��j�
����g���/��N���O�ή6�)��(��.{o�U�[���Ba����Z�`��j ��)��TM�Ce4.����a=��c�.�$��N�Ⱦ,:��P�49�8rQ�n������v�Ł����к����L��P������$���DXP����ۀ�����c�-��.>����U7�1Wr��n\"���hO�,�,��zE��E�|6�_�3�E[�A�X�jI��uZ��zk� �1�\ni�u�����S��	��>ǣ��N�j����Xi��qy��
<w�N�'�Ȱh�K�OV�q��+�������6����ր�kAo�n	N�#&��f�����^k'�_�]�Z�3�'V��j�;��9՚�z]e�*�p�tz�w�Ԯ^�ʼ$�+@�:�X{'hi�������vSQ�$�P��8��{���v�&$��� �z?o�,�����T��`�9�I<VGL��O��+oީ<-t�$��oIUK�H�r�CZ��aۯ�C��x;�-�-e�X2��K:��U�^��g��|+�a𩎸�/���"mUxˉ03����fC��3��]��Q���MEO������Q��cҍAaR�ttbhD�" � ��TK���֔ҝ�;�:�^'�i>7O�C��@,��!&�EG����)����f�(���`��O���WjZ|�?**�d���1#�����o��{����p�`��FG��^�[#�V�X,L:�|)�<����_M����I7Ѥ�9ǒXh/��2
."~\e�}>���dx��N�L��"˭�|��37[��,e[�FŊ�\���y:OW%�E�l�A#:U��j���թ��bޑt�W��͜71��2�8t�_8��r��s�Η�8�Í�HW`�9!L����#�����ג5|[
b�m	;5����P(Wk�L�s��7��ىm�t�Zo�.΍��[��¢=�J��� �'t_Y�'��ͥڵE�^�����Bl��G�L��wV��N�;�L�U#�� ��Mb�4.����}�����r�(U��х�$-�h�ֶ#�j`�z�h��xZ(!�*���'٫Ŀ���<(��'\��u�*�,�Xմ��91�\��$�F�~�9P��P��W���U����T����ie7�.�9mu�ͨfT^E>T�޼�Q��<2g���8�0�7�	n���v����s��.��G~S?u�AwR.D K�7��n��V�&��(�Û�}��oAD����?1XK�Ӆ��xa$���/�^ɤ7lhO��fz��j��/	���Ka�(0}�=yB]l׹_��53<���y?��D�b0r���7ѥ��cc��<}@L�ǄWi46��y�r̓>��fE���*�HW?����S:2J|)�*�q�tC�i�t��[Ui0+&%X&x
�<S����4�APX敓�hT���Q�'�����*�՜��'����*����~���nO(�R�����̹y}��ȳ9�S��#k*u:��;���+���]3��C��7�۶���4+�����`hf�W}R�ܕ݃�ח.�p���1NĻS����=�`��僟+2��'G�>*P�!�:�1Ӹ��ؗrs4V��>�N���=A�^4)��T�o���|Q>�$fX��W��� ��bdR���Lm�d�� v{�_�K��ړU'#�w\�5�ι{�Ϸ��>9��|�ƾ�ʛ1��AԵå~V<뗙UU��ا�hշi8Wg�������+����*�<&6�����ӣ�Zdp��M+�]��e��;9ARG\SR;mQ��j���W^��ͽ5dV7߻�;�OL>�g��]���r�|�Pɰ��鶄顝4v���Î��W���~3���rΕ�j W<���mE�����6:7���(�Q��VЭ7.�{Qw9ir��yeΔQg~�Du��g��K!����_ݫ��|2���b����w~��Y��QdݙB-^�s|%/y����Y۪��T���h�/�a��Rߌ�A%�5�����{˻�1C�f��ʸ�َ�Vo�f��\�RS�C}ٖ�|`=Z�Y�,����3��T��R�K7t��u�u�gt�G(r��;hM��L���+3�U;��xO3|s��^ߨ�(Q����!_m��l(�إ:hk�{P&/�1P'���WV��5�.w�D3/(��BI�F0a5��:���~~1p�%W��z�t�}���?�/��: vG�S�p*Z��T���ʚ;p�|���q\N��uʊG�-�8bT���R��	Ċ��n(�T�h�,&�+p����s9<��r\�,�8h������,:0)@pc���O]w5a�uj�(=�g�D�`kʊv�TgÆ�CCt�T=@�U$��wVc�74�8�ɇ�@0��I�,������#��-��`#k^�}����-�V�oL5��	e����4<��XCeLߠ��x&Y��kn�WV*�I�B����,�Fۖh=2� �Ǫ��F�(\V�yU;���8�ޫo�����p���#A�="��T��nd�e9E��EA��gJw�]0���K���h]m��Ok���%s܂��w�zv$��/^��i�S��}�ٛ�W���L��/w�B��Z�am�uuY��H�d�D�u^%��R��̀�v�t{O3�n���;]h%��;������龚R}\�������@��$�Ɣ�_@s�N(z\�{C'�ג=�	��[��deF��4�<m�+!���*��TS4:��R����gtH?yNEY�ٔ��X�
#(]�ƾ�'M�8��	�Lۆ}p��0=Tmc�=������m\��	�N�J4���0��L�(;6��E�:/���+N��v�"�q�6Q�ͮ*���1X�3_"�&��"�B���L�ڹ�O�y���uT��eH��DQ�r�{̯7�>
z��Tyu�n#�j��n�c��!c��t~Ge��<'�t�3�&�"��Y��ً/��97���$��ӡЮ
��|j	+�y�).�ޮhW%�&�i>Q;�;+�}]���*��KI��u����Ŏ�O�c�t9�g�Bd$�!]'����[y���YC� ��-u7Ov�e%���jt��p��С��x-|��;Im�߅�Z[f��\��Y����l�J�&�<]�ig���DF�+MoK�{z�l�!���������d��Ğ�K�EB�l!�	�+��s�:+«�t��Fӧ�7k�P�G.��-ҧ-�[c~jp6�n>ݥur0sέ���*�C~��s� �x��������S{x�1�
9O�Fc���+&88T�d�7*��)��¡�#O�-XU��u�l�f��ċt�b �.#~\e����bO���F��w�0�L���[٨*�cO���U�g�C>Y�9�5��'�i�Xb$N�dg�ŻQ��M��;�(�%����eƩe�W�c�����Nt��ҝ7$�(�q5�1o=�4�yM��y|h����������|}���Df��d(���'|���4�p&y��K�a�Ы�y��ę��2��t�ΗZ����]�n�����k����1���ǻ9�S���$���X"��"����c���휹�ׅy{:���m�"��\:��͆��(t�"(�b�t����1���-�X=�Y�>S�i���듙�|O���i9�d�����㭄ߟw�����KG����CGe5�����+Wg�]��'����#H(��Gx+�pz]���ٍ�$� �66�x�l�� RX
#(�ˎP!"6o���oo�����凼�;Z�k}r���#;ٸ�S���w�P,s�",C�mC>�U�;����qgj��M���ɿ�nb���
;t�Q���YǤC#F�{�Hf�J���e^�|2j��0�/�\�yOy���[E"���ڢB{˂�x�y0�{+�h4�8��c��c!���3��d9��|��g��M�%�=A���:{Ђq�b���,'���nL+`�cݷ�M�i���rX����3�5�O��3�1��,�2B�Jd��_i̽����.���Sf�]BJ+>�&P�A"ޱRp�O�L(��l��/������X�]ҧhb?.b`������L��
,Η���p
�mG,�iL${�"�7��P���-2��p��"��-Uz�wu�_,��P�ͼ�qV��Y0d<�f���k�f�h�ۄ
�nȭ	\�Q��M��SVj��륜4��.VEkT8��j��IXn���E�H�Y��MSiȝ9������}Eʻ�os�%]�g��*;6|��] ;&Gd�󣴱N�n���s��61iz��y�TS��6O<�N��d�/�V�趹tۢy�:wYK�7qt�;f���1qҎn:�۔k�z�lળ��qڦ���\w�ϖ�ޭ��R�9b8�RH��h�|2�6��:ݢ�O(��W��w�*�x�����!㼅[	jbQ<4z�-�����Ppu|�_�X���q�7�杶�9>�9��'�kE
BQ>��:2/�.�b�<S��[�������s��8O7vH��X6O���^u��ФM�*Q;�j\2�j��mJ3��G]���-b�g;GQ{H��Yfښ4
,ũ ���D��l�Q5���#��θ,�V�o?y4;����&�|��/c|%S�p*Z��D�!�=R�AN#�;bq���'��� N��8`Yˋ�bT����H��|�^w�0t	b���� �w.���֯�K���Qt��Ѱ��,]T�A�˼d�b�f�n���>���T��Ih��r���1�۳��Y�pJ��/��� y�z��1{� ��t^X,�˻�:rI��-�B�o;av�B������F��Gd�r\id��P�ןp�F��b��N�;,ș�VP���*J�I`�(f'�jc�fYͭ��0IR�W-�,�-f�������:O**�{+�Z����.��7Ym��,j��nA�R��u�g�pmT�L;�_-?hZcKs$\5�c�3R���q3C*#i��E��`��j��Sf���W���*�c%a\_&�柮*/���w�5e��K7���D�iE��ܡ]�t��a�mܴ�<U�+D�\F��Q��ص�"r�<��t�[�F�7v4yj�إ۰q��qGnm�}��h�üCQd^:ٝE��%�NC��χiu�3I�z��[D9�)�s��9]r���B]_W��\��F- �xuv֣f))��2	Ac�e̍}TM�V]�/mpˆ�P?sd�t��Y��K�gTs��7���*���.�?��9a��B�ٗA\ȈDWr���\�F���fY��F������Z���v���k]��,��s�tl��K_u�YV�o�ά͵"�r�k�cD��S�u)��rK��=��48�Y����{{s�G�>U��JK��N�k���lr��ml^5�uMˋ���t���]�5I0�!�A�tӢR4��ҠC$%�"���b��.4}2�lZ�%c���1���'X� �V�],V	�YO��a�*�չ)˕�w		'��l�#Hn�=6\�ڝ�\XaS �[��V��ȑq�e�@iZ�ڔ �H�h�e"IiV�L���$�(��\]�VNH�ìb#1�<�eB�"nkt*Pߌ5�CX� E�T^K��p,+	w*�Dp�Jd��+ ̏�"�n��,iJ�ּP>���5���v����K:��OjG@_�3�\o��I����nb���&em^]��u���9+:k��1ю��3���u#��̩F��a�z�r��y�����fZW|N��AgT��C Ρ.ք���va�v�Uʧ��T���lYO�+\�	��ZS���4�l���Sۡ�S�5�[�VT�b���l���u�\�m]���ġ�άK-��}s�����:��	�0��g �y�pq<�W "��ê����΢�Zs��Z�s��y�P���_D|�Ud�2��*�d����^s��ЌЭ�KV�V6��*E!D�ch*�f�����J��JԢ֕D�\�°��F�EU��J���kZ֭&�ڍ�m����mXҕD���j�LE�إZ�	�kZ֪4���J"��Q�A�\h����V�cV�R�*���kZ�Rj��J��Tl�V��XV���qYQ�ZYiK-*V�T�:ֵ�M%[[F�DB����$X�F����)m�+R�]kZ֢jQac�P[j��Z�Z!m��F�£*�AUQu�kZ��Ƴ��*QX�dU�PD�\h��b%Bո̹��D�l�TJ�k��E���,R�(�,*[A����sϺ�W�A�[�n~|�E�A��b`�<R��Ϸ6����[f-&��]$;���,���JP�Ы��s����w�v��À&Y���i�=��&�Y����b_�Q���6d��c8����W�+�"��/ň�夿����o�p�N�������uH�[`�w�]kl���V�,�l��Q페�r�8���YN}\�ȸ����<ҋ����;̲�([�/`0f��-�luFqn<�S2�#�������4���gw��\�<O�>���^ ;8;��q�-�����;�q��B�{َ=�]��{��`c#�2*C6'f�BG�u�ˈ���J��ff��Z���7[ں�{��(���h���&�v)Т��D'M_K�F��,�h�(��h��\���3��/C>�Er�P�x�UE"���$uJ���1*�����ږ��]�R/2!^WS����
/���dr�5������m�{Q8��y��>5;CX��s��u�iDa�֧�;O�o_��Y�(��MvK�~������P�_���K���d��!z�"�.ң���U�9�Yxl��oY���]G����uus��g,���z���o)\�n>����5�+�:}f_I���GenR�P����q�9Gr�\d*؁H,ģ��M�7'�����!��)�<����j�#U�C�k�G!��m���Je�Q&�C�Qg"�<�t�4�r=�w�i�'˖��	�^��V0���_Gy�k�ͮ�������� ��-�����B4+�S�~�j�Y����n��K8c�6��g[w�S�JǼT��lY&g���BhR�Y#�L�9�R"�Q�t�ԑ.�9C�|�t.7���(�)g��3�2
ɂ�	�$�1���tS7=���.w���� Z��&���f�f�S��,�ᓥ���]pq+Oy��S;��G�f�k���b4�t|�����҈P��`|f
P�0�i7���k�+�B�;���hu��DjVZ��>�< G�ǧ�$J�nN��|櫚�O9Nu,�F�	�"��dsr����>>�����0S��Z�nW�l�=���^��}^�~�;q�p�ٟ0p�FH�R�ƹ~&�[J��gS�U�(�vu|9�"��K�P�v,vT�s���Loq�oZ�t̘U,���o_�Os[�Vm�m���R|��}\3T�yi][�*UJk7o��]���Zft�+#O�x����S�����`Z)��_*�p��3n��W��a�n��"�)gK,��XQ�Ҥf��<��H���e�ɽǮ�ON�d�4'����G�M�Uzxr���R�������ήQw��^�<�껡꣫��KGU9�4t����U�qխ
_>�t��g�a��]놲yq,m�!Sb���DJ<���>5A]�pJ������e�x�v�Sά��Oz-�r��<����k�s��Ճ�Û���L_f����Kp���"��~�R���+��DC�)� ��S���N�j����\�k+*-�X�F�4~>Ue�\<K�:ǂo_�s�����,'�h��[��Lu��[�����_d����
��Ra��	g��BY�oB$�ʪK\+�+���9�`�@��YW�L��,RNK���q1�5���z�h��2����19[G6��#c��U4+fyg7\�m�B�6RRe��������Y
�E6�eg�8�&�e"�7��7�u`�C��n��ݎܗų����.	]ݗ��7j�!͖�TȻ{�\}�	ۼ4��pq4��@1o˃���(1ë�u�ؤ(K�z�I�Y=H2we�i�)ݠ�`Վ,/o�%{����`�c���̚:�O�3I�Gz�o�n����O�QҚ�Y��Q0qf�V^~��˾��%,�׶FI�8zr,����p���͐��=��:r�Q"�e�gMMufu&�ޞYK�6p�5��1GGO{�M�4**�Ν	ӷq�f�n�멜MLO%��6�9�:i�.��e�dҙ�cuӹ��[��(&_���]o|���$�ĺ�3�&���>���r��Q�E��T*���t�P��o����=s{�珦�	��<*�պTO�wU��b\��B4D�R�5-�I�.z��n�ҕȱѥ��2���W�'\�����K�]��x�;AyU��r-�o�t�\�H{��"�||n��?"�o��]VX��8M{(��{��������L���V�X_��j���S�s"}���ʚ{E��Wnu#D�;��eN�T���3 
Ĥ7M��q��t�Vih�	�S@ެ�8�������S����!���u���9� �өg>=��J��.�놬�0�x|��yU�µfE��
(�TEP7<������Dp�g�e���o���#b*T��̰hwKq"T�7��V1�ba4�%�/�2�g�$��=04��J�J��V~��)W*��e��1���=��Tx�DECY�#���#�~+V�/��蠴��aD
�z��_b��z��I�M�ra��+/��ET��
�����B0��I��������C��#�߶����)})[Nx���p��A�U�9�]��z;��l4����=.��'�(ٰ�`���s�t��<"MԶ�i�]����)ӯb����x=u<_�QѕQ����箸V���lA��N��{������Xu�|�A��S$�#�f)ǉ��c.S���;+=�NyNJ��=YY^?h���V��`zGCl0\GoH��WY*�����kg*�VW�mp��ޮ��[c9m9�H��}&B��.�j�B���wuk�ʗӱ�Wݼ�ݼ܌Ԩ�=W[�,.�w�}��V��ŀ����TVd�Y.b�X�	�S��Ԋ������a�f�lgh�ԡ�r�Vɀ�
�Ko��:_j�9��zg�~g�]����U-�H��peM^'��/Ĺ�Ta�s�ԭ ��M��/+J6;g������+�E�_��zhvt]
���K'.o�W�'>�1����e-�D�خ*�҉F*1@f��a� rZ<�~ˎa�<O��V*����b��q���Jz�qĳ�?����%;�g=P��w.v��8�,��HY����>�"\&���Mo�����~m�.��YOz9�[�Lx_J5�:"D�҉��s�
��pt��H������
q��T*��{3շMb�!Oӄ@-y ��M���0��>/���e��G��धW%��筑���Ԕ�q��Z�K�:}�)���KO��~TUS�d^�^N�p�s��$�eh��w&��Y����aJ5�E31bC"+�,4D{�uO���[+/5$�i+1�{XE.�Ȓ�)čb`�\B��>�Q#�
�m_/_���fn132�s��d9��[�@m�ZxY�9�����"��ZF��݃NqQ���)7/y%9fn�G7����W�R�'wtO�	�S�dWں�h�]�y��ֈ8M;4��#B��ʃ�I҈�zᜨ��?w�f�P�p��&{ԕ�X���,�y5��.b��5MKR����������~��,���4�Ұ���(�.bE)�_[��t��gz�}�*P���O���D<}L�C�E�<��u�o�`�{T͉�2
d�t���Tz���g�r���Z�U\E�a�SS�a��A�����y; C���D��[�ڻ:�\$
����C�sŞJY)��rR����7�$.�n2����5���	�*k�!�\d`>>�"�W�_?]]s��z���go��D��Nt�':�p��%�z8�B,���lLQ�
���F�M/h���º�5�{��QD�sy�r�,V�A��!ZB�r"����+��z���%���-PeӧX ^��*���J�|�J9b��!��D���;l�k.<D�W��~��x��]bm��ȫ�Ɵ޺M��ɵ�5`��4F����ѽ�g�o6�iނ�3��g|�+�I�|S�4�/^]��@�Huw�:���:�}-m��.�pT�JGGa1�93]쏻L��A�rq�}�k�=뚔�!�����ѱ��f�^���t�g]� h�*�@�k�y��|�<��%D:s����)"QD� lP��u#��#�Q9
�a��8�E�T2�u[mFP쨄�HqJY��9g	��܂g��㮘6�Y��}��3Zf���6�M����?}�X�tj��k �Ap�2�R�Db$8A�˸��[�5G5��LC���^f�F�S"�(lӄwGeY��e
	Z�[5ۢUO�OS�Λ�2Dd$`0��=���A^���þ(}Ց0�}v��گ�jk+�]Y�E5.�\
(���,�jA�/!������Bz��d�����6L�ъ��r��|��t�+�A��eŪ��,�Ӭ"�ݧ�Y��=�I"+����=6��OE>ʕ$24�1C`�Ş�8h7<h<t2l+�:w�:�k���&�.��9�%��Q�#�ےGb��ڛ#OH�v���r�����%6�P�_���ݼ���t�cչ>�=��n�ǌUp��K�H$h�t!u�����ٝ/�,z��^�ζi� +�EuL9�x5v�Sz� D�f�]�Q[�1�ܣy��#�]P�kM�]�y�$�v��x��g�W,� ?�z�ۡXk�h๞,չF�ʈDIEZ�p�dw��wQn�g���r�K6Ǉ�wl�)T��C>'��nvxзT�˔]�dd�y���<�(u",}��]Y]���
��XQ.י�9���z���sϼ��셖.�q��_Z�o��;�C�8xċtA�bI�ǰ�_�)��i�
7Y���]R�4��F��}mƁq�.~���[3��{�R���� 8c��OV�h�U��­AdC�����+L��q�N*���X5�-ĉͦ;����pM8}�.Zg�Ip}G:KA�yb,XХ
8{��t��<��3��T�j��#����ǽ�W�)Ѫ��^�薌@џ5c�g��tP�B�/�Ǖi^�.tӨ����f�f�]����l+Bhtf�T�r8��x0t^���E_wjOzTf��(PIs��ω��P/j ��"����IO�z�N&wVrXC�N��qj���Uʕb���J����yd��f½QVZww1W��Mg\JSr�W�L{��.u~���
XS��'ںV���WT�ۑ�+����!M��	��oZ���U���AH9�w,O��ӝ]��)�ea��n#JΗQ&��Lٲ�Y�9yH�y�����w�1���Qu�G�
�����k�Xp�`s�qan�2/�����Xy�^7<��F��Dz�,�`a����P~����!@S�g�X�k:�Uӷ��+�g���#^�W�O��xJX�f���/�ˈ́EtQlYZint��.d�ͤh8{l�&<���@:���@���*�'M�Q��<u]ӳ�ε-��Uv�E�샶��Ña�p�| ��Dd)򓪠B�f���ZZ��(����3C\�ҭp�6�w3�N�)�68Zu;���N.�R,�R:7���X�w:jU���}�؍��,z�=��<�9}~�K}���C�
�.��c�b���	� ��������
�l�{�y���<�[!��j��Z�a�Cӳ�5j���~z�Bj��d����{S�$���cwS���|����۬Җo.����X��!��q��t�[�dWy�9��)�V�U�b�];Fݷ/3�v��ލ�9��"5��ũ��J>_����Yy؟n]ݙ)�U#pz\�qVe<��jEX�vÀr{������c��x+>Ȣn2��9�Wn`1i٢�k��/	"��ŤѼ�oׯz+�]|��o���A�u�M����41�sp�����ȭ����yX"��X�E�w)�5`{�\�Zi�Yo/js\H��3��"�����(p���gZ�Z��:_`�`gf��tm�u}p�6u���]3p�Ԃ�5qU���6A]�J���&���l\4�v����"t�,7d:�R��i�BV��Z�&�1��7�m�/6�<�y7;�g_unufg9Y�\�<�ݻsX���F3�nM�lV씧.���=����@�����P�Q��#�<S/_#h���#���J�>���^b�5��Q5~o!�ԕ����üN�>Wٌ-y�����"���]Yu¬S�8���s	���vN*�
��=���b�g]�#�oY�\u+�)f������A,����M��4Q�ׇ��DT�k����-]��{C���J4bGFS���7ب�'�ie��:�d��k�qM�,�"kB��.Qރ��|�gU�d�ڭ���7�{q�|i�9����M7%[��nfǸU;�3j�I/�]��g��Q�@�G[����V
ʗqU�1J/��֎N.G�{};�3���n�ޞ�)�#	\�-�x	jN�N�ޱ�
u��4>:����e9!`;�H8ÙSV�t ���xyR�D�|�"��W�ĉXaǄp��L�4��Yl.�
��Z5r�$�|�F�{�̳Z�gf9�#�+S�1 �������B�\�ZY�'��+�p/%s��b�_vt�PP����1}V/Sk�������_GH�K{h;���b�0,�.��&��
c6'	r�o�RK2�Z� ��3oŅػm=;k�y� ˢumӍE
��r�J�U�X3Pb��;��#�
j�u�Q�޻]����x�u3�:�����x�#��,�Ɏ�d���/D6�K:��-��H��b'J��1��T�ˋ-[0���v!�p��}A)[�(&���9*���/{w�v�.�d�q��@е-�=���Rww��~�B��$�I#�M@�s.ZT\[K�%dm�2)r�1-�u�kZ��F���e���WVlS1��B�Q��Le\ֻ̺օ�*J2�F�Ʊc��Q�P*
Jإ�+kZ֦�YP*)[mUf2��kUTAkbLV+3Z�z4i���0̫.fYE�Z�\¦ZL�Lb��T+��u�kZSV�ز�X,�F"U�.$�Z(�����E�[h�ֵ�2����.e`��"�լiP�2��q,�����K�.��h�k��mmF��r�ieUh+�[���V6�\ˆZ�R浭jw��QPXԨ�J�i\LLB�YmD��-

��Kh��G,)Y1�-(��F(�k�R�b&&a�-��1��iYX����ǎ��PR��y�.&�^H�J�]u,ɵ-s��n��h�Zm��9��>��_4����յ���obJ�.��X��8p+�	T8qS:\�%l�tо�sa}q�^ڦ�C��O�
�q�PS�aɱ<���
�Q�Љ�=�*�ԡ�Q�wB�ő<�����xGH)H�*���X\�g�z��=��S�%�q+�v#���(T����5�h���wjM�!-�[��&�oi�}Q)Nm��Z(5�"�G�;}7g_9?NRm�y�W�����aU�����`��"���ӥ�q��S��~Y�R���v�V�m�<�y�A�&��1N�k)Uz�睵����B��Y֔�}p�,�ld�id�!��h��z�wؕ�bs��֖��o�m4�Û�R��;���O�9�7���m�����'��[�?_+v�!r���
���v���^�G��t��P'YK/�˝t�wu�*��f���\���0�h;�!� �v�t�	�	[|�͑�Ε�k閧[́���a7j�Q�b2p�u�y�-�Х7��.�&3�R�{�2wl���.Nٖ�#ս��H�=~ǧ�zU>4udc��
��/a������w�Q�=��U+|1^��V9�}^����������&��^����0i�G�Y��udH�I��F#�֖��	����w�>K�����r��D��D5^�8���co7��Ajo���h�
���:�?|�9�#"+d��rn��`㑷G&�)�!+9<7��&J�{}��ٶ��+��ܻ�^!�.�Wv`V)��R,DrhvD$+�rw�qq`�e^�S�TX���"��2��OW��Kit���n�9�+�Y���{����N�5���+Q��W?S���jR]�����I=���o����>ى��B=b�+3z8��=�l���Z��(�U&���'ɋ`Q��U�+�.�
�Q��fN'�R��C�J�h�bA�X("�-���n�`��c��,Ȗ�a�Ki���y8
�Ω�GI�6�[*p��
,�p���K{�^�{�N�*v����ր����b�����P;Wg�U��E{8�l��w�����O��T��J��j�̧æ^T���䛚�t�)hy.�'�q������Y��aW\C�K��¶���u.`g�6���cs�n; H��OWh�E4�u��qH�Q�`IV�Vi��{"�^��sO����㱭�t+�V�NZ��N����������'�^X�#z����@�':37��,vsK;�٫i���q�o�R6�&��ffc�w1�+;�5��A���nK�QY�52�V81��(�|���LOȶ�q�ҕ��;���q�콿z��x�:������� �Km-w�{�x_R�}�:�J[��,\s��5�㕼- gkJ�U�k1��a��8�1�^�<wD���� �ڷr�7�}N�9WBn��1R��;�v#��󆓼����r'�0T��ݱ	S`��\��m΋a(f��s�����+�f�&.�φggC����_30Ī�.ĭ����r((��d*�V���V�oe�́LG�I�l4���+ܘ�g�-Vg4C��VCa�s�L�qPZ��p�U��ā����Q��܃��w;�K*&S�ㄆ}��ԏK����H��!ք�W�}��]�\���ʘ�8bE����R�m�j�͇����Ȝw���̥�T�w�~7ʆ��K4(f&e�Fo������V�i�%s9k���X��g#����Y��"�d�ڙ8���t��E����餅M�q���}֑ԞwK�[��ZzU^��Lj���Y�[}bE�qe!���ıf����b�=�~�Xi��y,}��]��8I[c��������wVC�]-s����=g�2y��Ӄ���F٩���|��WN���q+�i�̋C�׉ӔU^�I����җ�!s�@#Z��c�t;z�:����7��B�v�V�c���>��}����Z�ν���ّ9�	݅YG+f����vz���s�~s�d;��p��]�Gα��{��_I�͛+�W.��$X��Z[i���o*z�I�wU����S�މvn�ߣ�=-X�t����;T=׌!���K�X��&e��Z�2e����5(��BU}�=�q�}5��؂�z�sqY��<�Co�[x��x
���\FS��fQ.�fQC�L/�'KW�{���f�z��k&���wCL����\�����[}
���9F>�nc��p=���.!]S3�+1Mthz��w�x4w�W���\u�Ҟ��Ӊ<�8�m��1�m�{��������m��B�}�U�NZ��z؉�󵸐v�����.ݨ��Z�v�a�T.�ӗ38��0>QN�̑��ݭ]7Z2��s�:p�=�iֵ�Wv.��j\�e�졦w��mI�Q��7w�7�s�j��s�4��*5;i]�e�G%��/�}����s:�z]W�V)����!�j����%�%M,k���9�e%N�x�+�cb�a�re-5��4P���ڙ�z�v���NW��ֵr���o溔��qNF���n��T�7��Ox��u���%���ɥY�)�bW����;׷�b�k�Jz�q�g��]�^j��ON�ث\�嚖���W"4?�ͨ�5z�r�'��{���\T^��UM�>IL+��Ѿ�u�F|)|����F��G�l���t�.x�,+��E���k�U\xk:p��JB�/����T����M���;�u>�ȇn�@z'y�ϧQ���|��-te��O�Vv�m�nzJs��<-Ͷ� w@z���L��m�����z���Z7Ak���`Kl�A�t�"���^�Okb��\E�ݹww&����6�5}���' )
�CB�1c���_T�V7���ped�l!��UЛ�ևI���!�c�3'3�f�y�'�W5+ԊҬ�VT����Ӣ{�N�}6<h�t�R���f&�N��=�;�2�@�g}��G	��N��]�w.�'zE�_����h�k���S_�'��sp:�Ok��-���oBːŢ��6�����*�uZ�qʤ���n�NVJ��W��n��K�K��=)�T�S�r5/=��~�Ք*���W����Fﭡ5��ڧ�ٮ^<�H�R��n%�y��1�z���Vn˃t�Bf�i�{n�.q����I5������\��\�L�S�6~�T�F��=���F2���7���lG����N��lP��T��Vx�Xֆ��Ȝnr�U��]|��c�oP�gi��u�r�tY�[�Z7�/��C�eb�A�}}�O�m�n��;�)c2r����"vhqA5�2n.ҭ^�h:q�W�x�t}Rn�og}`�+�7y7!�١�>��a��#T�r�#ձ���_Vͬ��]��j�v���s�ĳέ���_�������88�$���[�;��r���`lA��s�Fue�AXK��i|��Țݭ�R�:��z��8yȭ�_D��kT皷�NI
~�T!���Sė��o���?��lʪ�����w���L�vO,�\��"��;�5�q��o�ΚAtf�f������(�E��1��K��(���z��&׼��*�y
ŭ����%�z�<g%���B����2s�5�%u���Zy}ǒ�~�^Oêz���b-3rE�u��ᜮ�/����w�*�+�MMoO�%]�,#�}4�����Ȑ�NUw�n��ι��>urmN.�U ,hV&z]��T�V��ϫ���΅��v��:l,��;����j�jZ�v-��z;�ݘ�R�f��^��.�F�wO�M��ö�5�\��ԫ���XK%4v�ͷE[O8���a�(�W�	W�:��Ջ�M��J񮫵����ֈ��v�\��\ۼ�l�i�(����^�Ŝ��j�S�%R�u,�����J.5�y���B	�p�Y�˷��9l0�{����t�l+m��W�������,���^��k��M�yʅ��e%�:GvhM#=)jz�ժ�)�g�Ӗ�OeR驪��"���8���ɹ����U����0I�ܹ�?R���]�8̮�J��{�.�1sN/�K������c(O]d�ǞЗٷ���[��t�I�[BS���!�#�k��U�8�����SV����F�a��T'RR,+��V0�K��u���<�6�<���Y"�XH�!#u(��fa�����7�{'�T�����@$�!ْ��elr'�:]H^�N��m�{]O6�$k8_���ҹT	��j72��j9�r���1�p�+���X׻�o�W�;z<�uĞd��u�nWk/�>}�rl�8��]��-Λ3��H�+������?$#1J���?4�
��8�n�p��[܃n�P��[�yCi�� \�B�xWx�b��P�Vd�}ᆣ&9��Ȩc8�4[�����^ȍ�R�߃P�M�QtWJx�w�a�6i������V�C�3����wS��V�ޅW.��	Ͻ���㹿���>�R\ȴ���7�4F����7yk�1k�fV�V8́�[���_�w-���8r�������WQܯGWh��^:��z����*ڏuf���I�ވ��ǩ�]����GGک����S�Φ濽Ƶ�:|H�zn�ϹN�}�mO'Y.{>����ۥB�ׯ#�&��Mr����>�Ȯ���P��5*����L����?������<�QбB�?�*�*H��$�YP���(2y�` 
���C� ط���!��.Z3,�4�q.�K�:���P��TL= @� 3 ��X��)T
���(��kH D ��@R��P)	��UȰ��##,���)@��,�
Z��YJ��X��@b@b "*b�@b&Ҁ� "2i(����� 0@@`�����X{�0$�ąO��B�����}:Ԣ��߶`h
K���w�z�TA�QHT���M"�a\'V2����m���iJ�
\�b�ԱQ���~���!���F�ꟽ�M���/f%-a��}��GH��,���3����V��*�Gg�x�z_���'�P�D� ��?��4�T~�AHD)xg��|A�Pa��?�b��\�u��w�O�C�?��<v:/hu/��(�}�
*��E>6���^�� �q��	p�=���.�y�L�&A��T�� �x}�������xFFEĪ̱�\��>��z�'s�X��mZy�Z�̤ ���g��L(��W�C�	�
@� ����@��IP� ��	D��B䙬�b�HfB�(v�m@�X2<O�2#q:�n�p�?C#y0 $ B�
 �
 �h@���@���0"�~���9�ݴ�v�N ��H|�2B�#j��
uS1�"����9)�J����I�$J���
�F�j��Ѹ�4����x-R�s�����G�w`���e��Ub�l��ݪ�wyt<M}��ɷ49���D%�]܍�{��X���{��>��gj����5�[ �KN�oA��������K��~ ��<�a�'VPA�/D���D�fG��
(NE��j{��`�d.�.to�4�-��=��o�

���O�2\
)I�)�~���QTX�E	���+(�z��I��|��Q-�Hځ��M��#��i�-�����W.Q�,��).�j
*
)�?-�w�I�n�G>���;�>��_TNލ)s���'�Կ�u;��< ���K~���!�x�'����u�P(C�o$�w��C�`s�,�d�g�vp`?�������=o<���4F!'�M(�^�MR>���r3Ұ�c�����!�>C��ڧw��lp���؎�������l�=��$���p�\(�At���>z���)���S]\�/��n�3�|��v��ca~L��øxf���������gz��,s9��\8�4�!��D���W���x�$ݔ6"ؤ�C2�f�B]Su����E�v� 9Eb
������[��Gn�}>��u���H (1<�@x)�"A�4���5�&f���hL�o]����F��$�=����Q�o8
��t�]��BA�2�