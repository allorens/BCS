BZh91AY&SY�0�B߀`q���"� ����b/�                �                �                :� �P�R�y��uN�Z}ގ'����   X �  �  �� (
`0� 	 �           (��(J�T�H�")H�$�@�
�J� �$%)RHJUUUIB��J�$��)T� ݂TD�����UE��y���6{ y�����0��U)�\�N��y���������Qu쐎�n�O,z�=`  g��(� 9
��U�_-K�5*Q��Q*p 6`z)A� �����@ uwx����^��u���  @ )��E( |tPT�*�T��٩U_ �}� ���� s��� ��}���G��p�>�G��7�p�1�g���}�B���|� r�  ���IH ���� ��}�$� H准��_ }� ��y� x�}�	E������ =z;� x   �Eve :�*�J�**�)Gv*| fϣ������ y�}� ����4�| l���=���|�=
ף� �9� �s����@ ��JR@`}� |��{�=>��P| -����>@�
|���\�$K��g���zz �  �   {۫�%� ��T�BT�B��(%�ܱ�� ��{@+�ETp ف��=�=��c��8Լ#� �]�Jx�s� ��<   ^(>�R���� 9�Ҫ������G�`|���===�Пx<�S��zz9;�]� ��he<�R� 7Ȕ�%QE*����"�G��y�ǰy����� �=�b^ 6Ǟ�������
{� ǝ*�� ��=�r�� |�J 8F�͛� g��
����m�;v{�ع��(����� �;��c�����    " �   � �R� &�0FLb)�L����2����@=�#�A�      l��B�#&�&�`�#	�M"@��@@ �  ���U=H�$ژ&I�����=	������ï��~�
J��r8 ���#��1����}���~�����@��`���*
 ��AQ_�@�?r�*+ӂ�������������~���

���\�����
���|!�Od�����������
�&��_�`Q� f�q�\aGE�Uq��1�\dG�q�\`�(���q�dS 1�\eA�U1�aGT�@�U��q�dSA�q��a�1�1�`�d�Ld�Le�a�Leƙq�q�1�1�q�1���<a1�q�q��La�i�1�q�q�e1��N3�0d�q�q�q�1�La�\e�q�e�Y�`1�e�\e�e�^8�`:�c.2�c��08��q�� c c c)���2�!�0ˌ&2���0�`1��!�2�c�2�Yq���0�c	�0��c!��2�	���2�!�&0ˌ&7q��C��2�c!��2��d1����c.0�c��ga�!�0�.0�c&0Ì���q�z�c0ˌ��c��q�a�\`1�q��`1�d�Ca�q�q�d�0��q�q�`1��c�q�`1�q��c!�\d�q�q�q�`1�q�a�a�\a��0�1��Le�e�\a�&La�\e�\a�Le�\d�q�q�q�q�1�q�d�1��\a�1�8��a�	�q��d1�q�1�Ɍ��Le�e�L`1�Leƙq�`�\`1�q�q������CCe�fe�La�Le�Le�`1��2c0d1�q�q�q�fq��Cd�\a�1�e�e�e�q�1��q��\e�e�\e�fa�q�e�g���^8�q���Ì�ˌ8ˌ8�Y1��.0��c�8ˌ7Xq��.2�.2�.0Ì��0̸�c.2��2�'X�C��0�!�2�	�ga:�c#��0�&30Ì�Ì��c2���c.0���Ì�Ì2��CN��.0��c0� �q�q�q�q�z��&e�a�1�q�q�q�e�La�e�e�La�\`�\d�g���\a�a�a�\e�La�x�0�Xq�a�`1�1��d�1�q�1�1��Ld�\q�1��a�e�a�a�1��1�q�q��\g&Ce�\d�\d�`Ƙq�1�q�q�q��q�q�q�q�1��X�^����`1�q�q��c'q�q�1�q�q�le�a�La�La�La�d�c'q�1�q�q�q�1��c'1�q�1�q�1��1�1�1�q�q�����u��q�1�q��fe�a�e�Cd�Iǀc���c.2�0�$�Ì�Ì28ˌ0�L8Ɍ�Ɍ�Ì8Ì�Ì�c��ˌ�d1�q��`8��1��.0��c2��2���0��d���08�c!�1�� c)��08Ì�&0�c�0�qǋ��Xd1�L`1���d1��a��q��C`q��Bld1��Cd1���I��L`1��8�0�u��Cbd1��a1��Ld1���'L`1�����dq��fa�`1��d1��	�d1��Cq��Ce�fd1�`1�����Xa1��^���`1��d1��1���u��Ca1��la1���&0n0�!��`1��q�!��2����ce�.2�c2�3��0���	��8�c	��2�N<L`q��Sx���2=e1���8�8ʘ�/YP:®2#���Q�x2���� 0��ʮ2c"2(2�c�0���� �����
��L� 0���
8�������(2 c(ea����0��(� 2� Ȯ0�c �2 q�1����.0+� ���'/�_�����$��_�#�w�Gsn^��d��;xb ��yuY�1�{���{��wva�-ӉW�ʠ�We�tE�x���P:΃��K,��5�t���e�WF�X��S%��n�*{	'd���W:�7�s�N��pI���C�p��@gݻ�k��8��;�����������5���H��1��C�l�Zm	�nc{{ 4��sY�&hH�����#
�œ�s�bQ��JNn���2k`�Gm��.v�,	���<��Q|�EاJc������^� 
o#-4]��^]��h��e�w sMz��n���V��-1Ĳ#b��8j�-;�s�(�.�rS��'�`Ӄ`���*���pu��_ۋ��c�Ŋ"(�Z�{�+t���G�(c��tv�uM�-9Q����mm�Npɵ���qo.�O�H���8�M6�����H��Wr���9�� H-k���I,
�4,a>�0Z;n��,+�嗞7���\Ž_V�Ɏ�eM�m;*����8v��������ؽ3SZ�s���v0B/�S(�`�/j��X��ݼ�w]�W驋i�~7
3@��ٱ��;{�J����a���aQD����M�����$\�3v�̱k�{6v:]����ӗ��4�4]����7�`LP��c8�N�e�MX�t�[;��߷7�q\㳎ot<�ca%�m�3�"����5����O*�u/�y�J�s�v^VX�%o��VG9�G/E�E���n���ރ+N#�]�E��n����)����P2
E/���t�Zwv�7�8s�НG�|/ݵK8�:k����bz��&��u���-Eѩ3���$��@1����d�Ymͅ�Z �v>@�U��^��d@��׹�{�{���Ý�ø��(w
����
WK�GW]u>wr�{:p��.��y�������M����r=�{�
��=��Y�4����@�,?i7!H�ܦ�Y{������U���n	�wR�L�e�ryS2 �F�QL��G�7���o��~�隰��`��q�=�N��O	ç�vu{�� p<��惢v�0�C�V����Ai��!�Վ�9R�o)K<M�*�2-+lv'�0�u�@[�1��.��(�ч7��g�R�eF�ݻ�<�/}��^ۡ�S�K׏�;�Y���N�tuTS�1�7yO�-y�qLlR��qޝ�p<�P����<ΰӆ6���f�z��{V�Q�Gm�W��`�>��.�tWr�zA<��]+�w���J�Y�s�ѝ_c k{��h���w����j��pf��W��"8���a�bc�]�<#���O�ܖ$
����L*7�f�Mĳ�"�L)��`��8a�L�}2Vcϕ���Ί�L�v]�8<m0Ob2^,��w�e�Fj�c��0��~9G`�0�3���3{G@�tCۛ�F�����,�P��M�];�2cO����1[ˍ���@�����ޗ��DHA��f�˱	�H�:��8�=�i�H�����j�xp��tL�8��n7�޴����-�J'O�����������y�Ȩ,d������7AwKBYЍ��� �}��Bfn�b*��Sn�NN;NKa�g'��P�w7��;V�1h��m�zn��4�)wc�i�wop�o$n��`/u,=��
����N�S�T}@�F�^ܺ(#�&<�d:n�C��v�;�D����z�ɇ-����������'�Bx�T��p�<�XՆ�ٸ']���Ϟ�����9�4wM{9�r�)�zqI���;:T\|��V'���Ky�"�{�Z�P�:@�M�K�ov��}��zȴ����8��Nr��@4vZ���{���f��77W����>��i"��^�s{���d�GMiȶe�u�էIZOK�D:6M$�ɷ�Vwn�����X�}{����'8uL�@���"�F������Z�N���F�Rc�m�æ2�}�Z�����xNF2��E��fɔ*&.lm�f�R���8ek��<7gl͹�&��%�po�S���e55��Sw�<�Y�q�&rŪb�\9�kݐ�l�ea��k�\�[$�Ԁw.��C�s{[��GL�d�:�Bq��W���ty�>�slm�����ň�����4v��s��a��ٖ�rg���)���ۅ|7��l@-��Φt8 'OI��/�ާY9��ۄ�]�a��!�yv&wrO�y��	��n��&����sS�5֠���d���}����Oq5�۫�\<��NM�g8l�L�;�*�:s�S[�#ZT>�*�A�"�o
�c�v%�Oww �\F����B���OJ4-�- ��t�S@�j��T��t���q�6�'b�Z�s�3_J1ʰ���9v#���<;��G��-`u�%����<W7�9gQ�-��3u@�g­��c�j�1��N�ӗI4$�n�U��p���8�r���9�N�R�ZuW������g�}�nI�n%ϝw�l�wnK�®K��owD�&�Hf�.&0�x�o����w9��l4���\]ïN�&7���~�3F4!�ڲ�<�[���|0�5ܾ켻�2�i�n̍p�1h))�̲�w�M� ǌE7�@����V�L���Gש��ՏIڕ�D98���+*a@5W>\�^���cE��w5���d�D�Avn>md����^�RƷ5����	yW��˸Ԝ�9��O_��=�G;vMz&u��;AQ*�2�c�jnoe������B/�@C�G�����W^w\44�$ q��ڮ��O���k���+{u������s`J�p���%�)����v nv��s������;���13Jc<gH�p���rާK';s�Ҿ�*�*�}�
�8b�6-ұ���[,�ٻ��=I���N��h�wcN�5�pf�ɶ��"��:^L�q% =P�-ĦśdVhRl�����Z��v����I��tͨ���`P�gF�����͇�:���0�������=�i�N]G;�T.�s~�N>M���ؔ�l���XXD�S���dVN��:EG]C@,��V��-��kݢ[z 8���І�f�e���y�v���͌m���:�x�'��)��ь�ׂ\��Q[S����B�P���Mڪ��8������مޣ�a�÷F�2m�*�f�s�ek� �Z�ck��2d	^�3�"[�Ӌ>肹�R��8�l���l ��k7.�x��/7�Q����$�2�*�q�vO��N�bJi�{��X��1tEʁ����V�>lV&��gf�vS2,���HR͍c�����Wc�L>�Cj$�S���"h�Ո`��hsvޣ\W�ׯC[�:��n&�0.uI�zs�����[�p�,�Ƕ�ԑ�K�98��280_.�/_Z�:��9t�ߣ��	��\���v���l<���.�w)t��f��s��κ�wp����&<�-�J�"�1��*�A!��ӢD�r�Fw2�V�����\�d�)�LF�Gr�8dy�]o{F7C�"F
��ҝý��E�M}Η��N�\^ߡȝK�
L�nH7;�ƶm(��91]!���P�t�N:zugk�3����uH�k|#�
쌕�5�1��.)�&�� ;f����]�O[˄�y�Ѕ&��@[�f����)o	��e�'8f��9�ȮȨw)���s��Fl�!�Ǐ��V�SM͸ �+]��i��vr�kr��9�9 Y�żk����Q%��K�����Dv�q� B{u^Tv&�etu��/H��٢5�� �Rk��J'4�c.�|74���^ܜ+��m�s�Fn89�ә�q.�1r�7;�d<NWٗ�'6v�N`���Os9õ}��W'M1�M�]ao[&�T��bôr\�%q�6�=�#���5���s�%��Њ��F�ȯ��Q�;X�C���yrwD�Oc��]���|0����h�˻f.���� �-�4g50��vf��p PI=�2c�>����1؃a����L��9�׉��l���wro8s���{�j-�t+�.�7;/G�rtC:��r=O�����ٲ��J�R=��5u�^�3�����u�n"�7�ñ<Ѳ$�kF8�͈Q9�RS\~>�2��Wڪ��bѠ�%;���y�8#ìt�[�g^�:�]Sgdu*6K#�2��;�q݀.ȷ��ˤY����'�8�Vy�'�m�f'�sq���z�B�$N��"5��;d��8^.�Y2٪�RTf�;�;���f��wvqҪ Wtʛ ����2��K�n1��Iѽ8Sl;/;+�Oۥ�xp{��%�s�;��`�o79��A�mˌ�tkG2*��2�5+���4���C�6��\���ve���+�N�E'ɓ���j��"9/\�i�XrN��\�k�á<A�;.Ly�b|�Q�dNG�C�0y��`��={L�5U�q�:�=���w�N��ťkC��t�0�'~T�W���8a���9m��@��VdD77��&�=��8�;��a�r�!-+�ߎ0t���w;�ԑ���}7ii=�}��o$Pњd;��z��$-T��@�;����W9
`t��1L������qj9�� �.�Z�5�x�+ᚏc��@൜��Q };5���]ݓ�w$��u��g8�,u� O7�KEVMK��UF{xH=�݋zK�������������$2�k6)�֬#d�Ol3�ˋ��p��<f3�;.$�M碔�G�74��u`��M��4`�*b<)�q�{��'��t��C�r�^�@��q�vi����`M���<�&�Q}�>7�̫}��}Nl�(�G{�:1�)7xk'%�L	Oq�|R
�!���Q�q��fj��6�p��I[��㏇ �t]	��|T���������\".��K�e���*ٻ�1��6�۸qe|�Vrl %�↎�3�3���J�^u\P�հ�q�zgu�EGPU�+nv�u/���{(��H�;���so��^d2�"%��k��{���2F��I���;�Y����Nԓ�*��b�w����pC���-$;�&%��f�I+d꬙�A�^��k�5���$�Ƶ��4y���;�,�4���j��z�j�_^�����s~q�#����g����vP�۽�Q�Os�$��e�J�B���[¨�-�Ͷ�����Ӄ\xDV>˭s���u����J�c|��s�����]���l�)�l<��y���ǹ�-��t"�p�ѷ&Iznl���v�v��-7����v�<46����������ld���_p�����٢�m˻�T$�Y����=X�L���Jx�	Uj�Q������Y���l��{<�
���鿧���)M�5c�ہhG����3��.����m�Ͻ7x�
?Ha9�����*U��[�w�c��s׺��`�ݱ�$tu������G���!&�����?�����&a'�؜H�xiWo�3��������_�h�/"��m��A����rF��J��]%�������&W����.%c"f��h�G��Wn[ڱ�׸�úM����w��(�)�R�5y��2�^��ޔ���8�$���+����Of��wu�<uU-9Du��y���=�����xś�.�[�F�wti	���̏��|}N�3�E�J����S<g��+c�;_G��G��#U�f�<a�����鄒1�L�?�m�����_q��7qа������x�$]w�gw���^&�I3ԕ���O7��	���������H7��{`|(��׹��h"l�3ۧ�/5�t�vh��j�K��J���r�X����Sx�3�e�I4��?��|:�+�=�\O8�J��%*S�^z��_�t���A��]2�^o��x������[��1O���oC���2{Mq�{V��nL�$����g�� 8�3n�z����������iPk�;~���_g��f��3^��|�Y��݌L���s�+�`N�i��+"�շ^�%��0r.��{��V�;�Zgܴ�t'�ߡ��qux�Хm�sO5W썥���4'S�v ��z�s����z��=�g�wg�oc�}���6���㞳?�S�p,[�p���n�q?���|�5�	��$�Ǟr���n �XP�u�Q��2����\���o�S��io𐉯��>#�8G_B�)\�\GzZ��e
�n����3���������7��Es��,Eo�����O�C�=�'��po�B6���Ҷ�o����d"Խ^�_n�ýf`|�um���ΦV��S;�?��|F��~���n��BI�ID���}�s��:R}�O�Ǐ/,]��|YN��3|*l�S�ݳ�h��p�V���p��w�/�:�����c�<<^�R��2n���_��B��3�=A��ǢH;	=�4�����z{���;�����Lc��MD�F���~����Y����se���Ս�Y��*}!(�	�G�o����glY�O��4a���EO�_\ܺđ����>�J�*�k�w�ڢ.�B��9�
��[��<���k�o=3Ҵ��z�ʗ��K�Uz���p)xl�3���/B�by���S������񶐏��ORUJ~x���ҭ}^L�C����~�|&���?��?v��y��ljB-�/������C�`�
��%���x������8do���\���=N��7����_�1v����C�^C�;�i�V����Z�yZ6t�w�)��G�r�ee�n�7����~��#v�?'����̏�����~���$@?�U�^J�%)y"�r
D� ��iJy
� iE ��AZDhP,����IP`�"�$䢅" ��J+H��9"P�(�@	P�$�  �$+$T ��� J� ��
���B��E��@JA��V��F�P&AI	XH V�	R�@ ��AF�hPB�DiA��@)
D
IX@���)T��I*HT@��
%(Q
��?��~#~�ԉ�3���y����{Fj,8���B�θ�h�����]��4l����Ai#ེ�z7�>��u���^�H}Vni���[��zc�̽�pJa��7Z"�bL7�2��Ƀ6�[�hma.kO~y�_5Ԥ�����9�3��c�z:����n��%]J����N�>�B���a ,^q�fP��aj�&eO���=e�/�X�"��h�K�딧�i/e�HA��<*:ؖ��|���~~�̠�{��[��=�Q�q��F�/�@�YD�����]��"@-H�JO<c_��s�FT�4#�o�U�x�f����~?��-[�t	�fLY��۾��
#C	3���Vp �$�7P�`2 (��7n���R��p��.ϔ!����d�qSL�e>�HPXz��ǉN��z#��>>��������I]���xP�Cx�/)��[������&�����TB����HjX��
��3jL_���ߟ��`�dH���2��� S�'!�hǪ��(L����;�1���;�y����滥ͺqNuz朂�%/�>st�qÚbec8
J]+u�w�U�[H�xw����Z��G���L/C��w�[c^r�׈a.�߆�?*�����>��3ǈ0/̖�\�]����ό6��T�J�1(���fc���������4�#T�>~��f��ƑAaw�A���+�t�Csa�i���0m�'X^X�e�S�<'��r�jj� �,�͆! a������ŚBn�hA��?#�n���Hoo�x6�zf�t�����]��&�b~���<E��ġb��s+e�^V�0��6�����g���֒�Z�~h[>���ڻC�w������鵈�40�tk��nݳ�{ӆf��9��_3����(���i����QU��~���O����T �@`�?����#�G�����O�����߯�<�D{�����9���g�Y�{������z�".+���w}��g/{$�v�=�r����"웦�����J�Lt�g�9�B�O��ڝ��}�<h������=!y��7�vl��NE^��r�{7�/�~+���IC� ��[������g�=pj4��~�{�KZ�������7w�+�ގ�7��V�{�xPs��qz/s:�̃a>��n��=��ݱ#0{çj��B�(1�����F�cQn杢�7.Q��p�p�=��]ό;М��<q�xg{w��%����^5_y�����<�m������{/�c���]��bK�xk'٥���j��טּ�C���{}�|�^���/�d�M�M{��XgE,���Wr�����bڷg{�yxk�M�@�[�\)4`����<7&-���n�z�����LVxm��o�tO|��|*T���!��y��w�^�d�Y}�X����9�fw�{7p�/s�vc�:�)�KΑ �;��,R����n��~k�v_�{/Y���]T� ��n(����e�����&xˇۇCO{n�*Ѭm<w�sTbB.��}��.z�u����z�=��6�E煬�3�����y�������^:뮺��]u㮺뮺�tu�]u�]u�G]u�]u�]tu�]u�]u��:뮺뮺�u�u㮺뮿]~�u�]u�_n���]u�]}:뮸뮺��]u�_n�κ뮺��]u㮺뮺�u�]z뮺믷]u㮺뮺�u�^:뮺��]u㮺뮺���]u�]}:뮸뮼u�]u�]~���뮾�u�\u�u�]u�_����Y�u��]u�]u�s���y}����{�~��no�ϳt���qx��͏���ot�u��M$�T�s���qr��~sɟ%h�2.3��S��U�X�>1��¨7��v���^_�Y+/,X��§h������/C��MR;u�k��x�{��Ǉ�Gi�vz��S=�fh�C�HD��;w4�s|���O�7z�]�_�#3��bO�O�<=����_�����T^�ӯa}�c#Ƕ{}�R�mN8-AV.�M��w~��E��8�'���[�R1F�fr�����!�������{<�r�}|Mij~|����*ҡl6v��x�`X���{�z10��ʱ(�7X��ޓ�:��Upv��&pM����i��Aϡ����^�G�������ݾ|��}b]��f�Z+;�(ǥ��ffa~�`�z���߉�ο2�}���#К��?�̼�R:vh�D�hf����/1��N��F���d�s�`�3�^�R<J�����R٭�����.��f�<�8/x������<��x��{��fg�gg�^���]d��[�鱎���ќ��I���V�v���&��t�Su�o�R����l�μ��<�7���6d�;��}~�/�����_n�뮺�u�]q�]u�_N��:뮽u�]u�ۮ���]u�]~:�:뮺뮿]u�u�]u�_���뮺뮺�뮺뮺���u�]u������]u�_N��:뮽u�]u�ۮ�뮾�u�\u�]u�Ӯ�뎺뮸뮺���]u�u�]}:뮺㮺믧]u㮺뮿]~�u�]z뮿]g_n��뮺���]z뮼u�]u�]~���:뮳��뮺�{���dUX������%� w0_g���,�GOz'C�����=MnQ�o3��o��ua!�K�'���.yg�u�´k���G��N�wQ���2v��oϵ���&�8��7j��L>=����"��6�|_L��e���4���sϲ�̼���}6�^���C*#�?����]���}|���g�0�a��w���CI)������b�d�&v�u>��ۓ}�wl#��z�v�
�x?g<�T�nq��/��\�K�>�X���7���ac���ao`
���<]��9�פd�y�Ӂx2^C�|ɝ��K�F�Ҡ�j���}�5g��?b,y�{6��[V��0�	���3�7A��<�8�_��<݅EN!T�q�vx�9,j���{a�{��`�-#wO��W��|��dI�l���<V���s�H߳���K���p�!PT݊��;]�E���[���}�8 O{l�vGs���'8zy��%����ϲ��z���|��뾒?j�}�}k���su�[��3V���n�t^[���}���i&��{����ח����ݱ�Q6b��k�/���n`\���go664��ڛ�뮺뮿u㮺뮺���^:뮺���]u�]u�\u�]u�뮺뎺뮾�u�^�뮺���]u뮺뮾�u�u�]u�_���뮺뮺�뮺뮾�u׮�뮺�g]u�Ӯ�뮺���^:뮺뮿u㮺뮺���^:뮺뮿u㮺뮺�u�^�뮽u�]u�ۣ��뮾�u�\u�u�]u�_����_n��:뮾�u��]u�]q�]u�}�9�s=_7G���=�$��A�6���w�2�yjPe�e���yg؇���sRe���]�*�綸7���.��^�Y�.Xhlw�>u���d����W�2=[F��`c������ĸ�N��D�s�"���>��ئP7F��a�>n�T:����s�����Ʉ�����^�i����l;�܄�kl�o��쫰f�:��xs�$�nm�Tقo�c}=��C� >X��1~���7��F���F���7�f�Q]�(��K��o,�0X2�й��x�K^��s����0w}����`ސ��p:ǚog������BVy��a3�@2
̋0�_Dc8�U4�����}ߎn�Z�R{4u��¹{g��uu�z�ۖ�ٗ]p�˚��7x���or��.�.���$����8+���KJ!��}��9��Wy�Cϥi��������}u{��8���u�o�_6k{x�����|u��u�+�Q|s�RN�Ĵ{'F<:��ܒVI�O���9�T��.��w<�Q�i� ��xA��弳��2G����~������ߟ2��������뮺:뮺뮺룮�뮺뮺:뮺뮺�u�u�]u�_����]u�]}��]u�]u�ۮ���]u�_N��:뮺㮺믧]u׮�뮺�u�u�]u�]~�:뮺뮺�u�u�]u�]u��]u�]u�]u��]u�]tu�]u�]u�G]u�]u�_�����:뮺�tu�]u�_n���]u׮�뮺�tu�]u�Ӯ�뎎��׎�u�]u�͌�n�a�Ӌ���U�2���e�����nN%t,fVb�$b7o[��e��6�������,r����I�ƇŰ�x��ˉ^)�ەw�^�qޯ�OA���u��A5/�1��x��������e(p*�ó\�/#�ֶj�]2��c���WA���Wy��4(��T��
Ԝ����_�G�f��ٺ}��??��\��Γ/-=�&h���m��^�ǈ�,�R=v*��{�Z��N��({�v�w�p����sQ;���q��������JY�͏u>{�����������k�劂��5���rˋ=�u�毕Km��{5n��<&=�r��X���,S37ޘJD�W���(�=�g��K�����	�-�l^�I�E�BOղ��d{ �|]���1��O�_�ӭ��	�>-!�;hx��ȥᵘ'�����v�ft�p���'Z��,p����	׷>����{��u��xvs�9H�\5���ɻ4[^pPz�v���|xƼ�4^z�:�{����߳�+PD��X�\�$��x�^]o,�6r�n}�8���dq��*+��s�`ﯼ���ź�d��v��>�(U�4q?g�G�k�4h��7��U�� U���[���c���.�~X����X�\���J�yc�Y�Lq��t�������`s<��1u�NB)f�����z_�ͤ�g#��m���Rހ�oX�X�F��k�t@�[���<`f.����|�e�����U4PF�qTy��,��>���Cـ9��G��(=�����w;���tS*ȏ�&��G<i.	7>�h�2A>�L�=y�����m=��ĲK'YvJ漧��s�
'�����UD'T�R�^KǐY.О�wv�^�yxh�͌YWU���i����3=���`�s^��[�Zc�k���3��ǘCQ�w�*&ӄ��h����=&=˺�n
�=ü����<,����<�x��)��ͅC�l|�����zcH0i��n�����K	�lP�yo�)���g7�uf�ה<�
=I�wI�H+C��ofӵ̷�v��x�30�ء�}�k��]d�@=��p����s{gz�sk!�`2+%,�;�:-���t\���yc�����8���g�]�9��9�[���3���\=��p�Έ�\Id�5��cn���.@:�/v�F��{03���8љt�2E�` ����*>s�ys>�ގ�=���"�R��Ҙ���W�{�v��V�j6����)U[;����7T������Y�^o���u�y;}�վ���{Z���,d��}�7�����$�1���n��LJ�x���Jϩ�g�W� �nxs����T��f�g�ƛޔ��7= >��k�U_}!�(��!��~�w���=��}��5-g>϶���Ζ�������;���Ք�>Yǧ�}K�v�%�G��T��|�8�>��e\�ӧJ���?�>��OK.�sź]�\��~=��x]������۬�$%��<�q�u6�>Ӹ��gVW�z�~��Rn���L�[�p�y��g��{��3�Y<�`@qc|y�f������,�ގ�2�'�M��/y�M\�qC����pmk�1w��8=�f��b�χ�����ݳh��8������.�<��0�{��g}&P�[��w7�,]���A{ݞ��]�7��9��A�S]�}�햬}��D�;�oLf�ۂ��'�v�i����7|��w/a��{3�7|쾞�3�fN�y+l�}b}���[��/=���{=>��z�s�݃dLxk��5�����d�<�Z�uڗ����H}�b~j���{z1�O{riǹ�K�k^��-���OY��9h΢��=��'{eQuےLYS�3ƠJ�U	���	���5w#��1�����͹�G��/Nd>�;�� �]ƹ��k�ږ�]��\��nLZi�>�����A���;z�U�$|�|r>���x�j�K>�7�d�@�Sa��{��#���S�p����V�g�y�ly�n��k�0�N7��>����w�KL{޺|�ۇ��������+�$�Dl��-�u��b��_��������Ѥ�����MW�t�[���m�Y�K���x�4�hXњ.tӕ���w��o���ȳ�>��w�<���?}�u��x�,枅����gk)8}�<�S<�y������6��x��}�ݐÅ�{��A����%��w#�uW<q��S���opɠ؉�DS߀Ͼ�K�񯳙�K/q��q����E��x���>Ϥ���ܷr(�'���G����AryY��w��|o�sK��h��WW�'�iR,�}x>�:��FqˀDr��WQ�����wC�Dk�[pz��S�>>���a=��wU�Ov�v0t��ҶkJ���n���@�a����}��F<����n�7I����K��i\,-{��.��c�e�����\����+D�䙇����9w�{�=����At���J餦��ȦG+���Jf�g���xR�w���Y�n���u�X0������@��>��|��� b�������yOSݷ�y�pl��kw�
���"{�{ظ���L*�yގ��h�3lc|��]�]�nC��-��j��i�+ow�z��L�'O"dc9=|yp\j�t��hV���Q9$Ģ��@]=�����]���|0��������@��{7���x�c�\��e-]4gL�e�
���y�ʠigOl��V_T7�t����'gzw�<�	��M���XlV��}�9�١�ϻ7pCz�K�r�v7H��lK)��4�ͨ�y�#|�J0n[�!���Qj~<��7��`�rѣ	�6'U�Ю,��/����:�yo���\~9V���y�w���}p�03o_t�gzj'��G�Һa�b_v.������x���x�9گ���M,�N���]��s�M��xmG�#$p�d���L��}��	띇R�����wo�[�(�|/N�{)�+v���V�fa�O{5�z��<_�f�=�뛽��d�+=��M��?y�/�CGݺ�0W�nZ�u�׷ۋ�#�~��EE��8�"�uo��K��R^6�!��DgH����|}�јp�ےw�wG���������ʦ	w�58N���2tS���._p���o���W��qZ=�����о���x.���K�o����\�~)*���_N�Z0O�$���T�P8�&��3/y��>�!V�B��+|�����g%s�po1S�ޗg� �����y���=���=5�w��޸��xu/M�@$�,�^l��ʹݽ����X���yV/g��=�W�:�n��F^�""�ǌ���6�#�y��yyx��5+�?b�\�ήCO�_d7��w��K����͜=�7׻���.��Y��6��A�{���`Gv�Y��߷8K�s��qh��2e�W���+���#�eK^>�sd�|Ok\dZ�E�fQ+�u
;
7)Y�g{m	��.�[.�xR�>N
剻�֋�9�w����i^��� �=N�_2�Z��r۾J,��<	��eh�Yd�_�r5Grvv++�>����q�4����x���W��M��L����l�yf{P�奾�'�0�mA�T��=*���}1p�/
}���;}�9���C����9)<��/� ր����ߟ���QEu���g������@G����?��#O��Җ��T���4�4��e�Lf"��d0]��u `���G	,ay�=b�"Lb>_j>�~����|�[?�}HC�M4)���������v����G@��ε�^fqtu�n�$�
��^Xr�c.6�LBKs,e2�4�X������f�\�t�2浦tR�,$�Bv��Ō�ErR���L�t�h�n���b���e�j����!�u���:�b��8��MMҥ�f�ap[].��.�6�Qk�%��{,X�����0�ՙ2��W�.�˴�!�̺C�����<��Z��膐At�M�t��nrY�&4���s��d ��-�ݜ�,6Yc���e��c��x�4��@mI�u��Z جMB�m�SZ�ŗm]�uUs0���:�W5�V�7���D��Wm{L�-�+y��:���J�iD1lJ��,�a��u]�X���k�DЁ[�Ů�#�`&M�;m�a�$ٺ�\j�GA-ʹ3r,�s���Z�3K�c���@Q�n�+P@��`�cq/][�u�ciKB�MQk
$�7V���)�0ͦ%v)kR�qF,�k��5*EX��76YI��ؙ�j,l��\��bJL�-�۴�YbT��� u�Җ(��&&�ױmW0/-ٰ�,-�6�m�g^MW1�&9�-�I��(aYqBlmE)dH��vBe&�mN;:*-�E]6)riN� m��M%&b�Fa3��M�e�6�SB.�	z��x���i�%x���M���q5t��l�U��M-֥x\;l�#��[��[hmMlH�RbP�Ҕ�I���4J��l���Meee���5�X��35sQ`DJ8�K6�h�6!��
�0��
�F�;��Źx+�6.GZWiKD3b��d�j��1!m�i��9D���a5�v�+��u[�2ز���l�)#�ܝ�/V�(�Kl��:�tf-�kv��X͵�7,,��%�&pW�i��w'�ƃpA��e%Ф�-�0��8�ݬ(�·!M,[/Qp�@).�	Z�h�fL!E�,o$#��{L��k]b]�a����C�p�K�(�4��Q�L�t �h�l0�I�(63cV͇��M`��M�c�h���b1��Gb�VR�Q3n�e�h��	��4+a�ͣ@��vk�6P6+3H�"�s��7nP�G ��DM[�wb4�-�:hir6e!(�Zf�`���s0��k\�P�!�S�5�7J�RhT����Viq����6��K���
1q�@�Xs�	S0��K1��	Y�磓Uc��ЫY�8��i���ι�e�<.����ԄYZ¤�f$4�`��Ѻ4o\��*�.��M�A��u���hb���f��o6��S��X�ss��&w`�A��L^eu�P�6(�wgK`��)C;2��D�{uЖ�YW1�T�vL[�� �fYE�&��rCRi�b�i,�9��dmJ� ����Abq��͜۳���e�[�X�{!a�v�#R*R5��jg�](�äZ��`�G3f����Ae�qp����-wV�3E	n��D5d�zܙI�����%�섩�0ٺBih�2҂S5�jk�!֪L7ԚX�$M5�W,i(`P^���$\�&��-��D�F��Cj�G�ҡ����1 CJ\ꍶ��Fl�&���sd����L�6F�b�1� �)e��m�6$Q�:[u���aŕ�.E��-���y0�H`VX�9f�L���	�qq�e��Y�ڰ� ��p�eY���<���%�c��t3C	IN�Yt��F���N�K`͐ND�B\�y^k�R�Z�!kY�#���G7rb�̹)�
"�Ҥͱ�5�F&2d��It	t�2�)�����Չ�Q����\��D�	7TP\,��l��t2��L����ג^�JB�)��%؛�I@�����#��K��b��@Ͷ�6lC[��-Z�p�6ڹ���3s�.�7[f8Y���(&I�X�F5/d�FU֖��u@�{0[zٵ�g0�\�eׇ���� C���B�ga��ÅͦW��iNEs�@���a��q	H���e����˕��]j�#���C7�k��b��:�� [x��h��U��C-�e���:W*�Iv�M�`d�Rf�PAInT�ٛ�-J�%�#	�RX�f��
q�Gpl1��3X�՗J*\4���״� X���!ڋ#j�Ғ��V�UW�t��Z�0y�[p2����iV�U�0���&�eՎ�З[�V�j&Hl�9�R=J���;F`%�.��3�\LV��nqx�.����gT�a6�-������6�̲�5��&��W�),n�Ј�Wi����2��a�k]�T$m,�,t3�*�Ԥ����3S[
-vtf�n e�%Ѧ\��T�Ąecp0��1��ڕ&ql�`�h�4ysFs0��jm���+H:ݰ�������@�6[x��6`�q.,�"mHR�H��.�L����jDЊhـD�bV'.��f��-�.^���l��J�&&#nt�,��;F�լK��	�49,�-mM6�˸�
��Ġaƹ�R�k�\�׃"QLh��f���ի��bk.��Р�+�J� ,�.��X̼s�׭�R�ƛK��6�읭[�v�-�&.x�i�e�d�"�H	3J�L�^�jL1��h�[r�f�q5K���0�6."vX�`2]dȶh��"`ĕe��(�r�L4���4X��RD20��\])�FZԚgh��+wWE�ms"�E�t���V��!���ڌق��D.e�U`�&66[mR����5�q��cQ)[�,��esVQX\��;%4�e�:M��k3���en�8F6SX1��.�5�R�T�RV��Gqf�����@�6�ebh�2��v�g���x�a,0]nYcN�d+r�����0l��E,�!in�*,k���`&06����͔eZ5����-���4����Y� ��5��d�4� cup��
��,ԆMsJ��5�6a�X̥�9��nJ��ő��ힼA�u���2K��a��q:d��
�m�c�jT.E�A��BV,԰�l!{b���a�p�y���v��],{��/%�[	\��9�8�΁F�v8*K����E��-�ƅ)�n�F[p� ���
ݲK�	V�L&�Ü�9�K,ƍ��"V�uyH�"��AF��1.��i[B��e��bYu�Zsl�:`K�D�\��7��K�Ƥ@pZXL�sիb�hТ6a�j��-21�f�ԍtLeLՎ�[��R�2GU��Y�� [m3D&+
%���TY��Ό�Q]��eJY`�6)�+�q4n��b�[fX�.9�%W6V[�(b�Rҩki��eKGV�e���9Ͱ6�����[5��;��u����u�X�1����u�,�ڥS=M��2Q 2�sL�Q+)�c(ddr�����Crf�7\�F�y��FgL�G�v��J�2.+�-��Pn5i�f��έ{B�1�Yx����:��l],JG�vl�p6�Ѧ�$45I��"ZQ3t�K�-���Vi�i\S����@1o���%Jhd�k)�i�����6]�bK"#��K�]Hm2��[��t4n��Ym���bZ7A2����X3Yvܒ��kM2���WXs�Ա�.�:�=��S5��b�iMDl�6�*^�º��Mc�˝{l9����W�ؙ���S�6��Dե�,���e\�e�l�W4�`�6Ķ+�E#3�Q.�"�n�a����D�:�L��en&s+���e��3@��6��(�hr�uݫb��r+�-%�^5%]Z��%�ɴ�V��J���)Q����І��3PK���]-�9�:�+8�2�戻[�I-7Ui�����E��\F�D�E+r1����U5]����*����c���;�Sa��l��r�̪k����Yn��j̪�e3U.S+�Kv����ʭU�UUUUUUUUUZR�G��na�����a`[Q����`��MB�o��B`���o4=P���-<��m�޾<L��6��~�>ᚶ��Ƥ� �x�ժԶ��u�ǌ��'��C��ؑO���{�z����ڒ�Oc�|�)n��.�9��'���LO�<��<����$�Չ�ɌF��*��T�˅N�۬��5�(����W_����u��뮺뮺룮�뮾�A�^��9�J�c-�l�C/2VI��c�6�a6��~���]~�뮺뮺:뮺����r}A�_������E����Ab�E�k䄶,�'������뮺뮺룮���ND��)P1R�+�1���+ޣ�ó�>������u�����]u�]u��]u�_O�h< 1HȇmW�C��=��Dc�����Ҋ.�K�+��3%�ݲ��XJ���֢8�X��8Z(��A�DX��a�%QEu*�@�,-̡"�"�QJ����5%��-��TA��FI�lc �TAV@m(�\�T@q̨gY������"RZ�5�7*�5�b�fb{kƢ0 ��l����c-�V��xc���(�����hb�KR�e�
ʔڢ��P']f��E@�Z�Td���l`-�5���48�Ԥ�ށ	�JSXXҔ��tK�@%����%�%�11N�̃mZ��0⠡ή"	�)����`[!H��Ƈ�%q��Sr�$��ۆ�R��M���J��ӛ��I�����*u�(��^B����^�t���g�d����C���p宖�Ԏݵ��ڀ�e���mf`��ʕ�e��6�	r�\\��v��av��	C���lQ�W����i�)hh�s+[0����A�mN�0��l�[\�b'm�k��T��UՎ\�ҩuvcGU��n����X�f]jk��3/$���h�H�Ԗ=q���Y�^��*�V�4���1v3V��[��ZBZ& Q6A��U��eX�k�t� ��!�C���&Kn�`4F!r�ֱ])��q	B���8�	����tp[r�lɥ�2X�6@p�i�3e�C��Y��� Z�(�(ˋ,1�hƹt�˙I���(i�m�fq�	V[ڹPZR	�#q���ZQ��̻R���i�X���\��Y���k@��l�hf�e-�Z�2�JVa�.��@��f��og[��݀k-Ђ�Td4E,,`�A��v�F���-i�QtM�kV�� T�h�P�{�DT�����ݢ:C90��:���[r͔�(e�Z��,�R��C���q�vV�:��m<�}�b�8*�%Ԧ(�qJ����G<a�ء�
�K`F#��fXCFK�Q5�lL�����a6i	L1sa;@&Z+oe�0����D�A3)Y���P�M�:9"ؘ���f�{/SJ)H��E+����9��bc�Ʀ���t�^�%Q�-��2��asIT�K�C�\;fh�(BƖ1#T�gS;mfC6Vڭ���PLGD�K�&�J=�2��m�E��6fA�
��\�M���46˫�ʪ�,p�6B1me��-�m�6�72�3+�,cbBI:v�8�w�W�
��5J�B"�UU��A�)ca�!V�6R��J޴z�:��V<��iV*saj�y,!X�ר-YT�0���x��)K�#D`u��%%ZVR��P����j�H����6��6�������X*T�QeP-VP�e��e�6��kU�߯���.����~9�匒ݼ���dre�fw��f5�wm��Q�H9�'B �E��kO��{�;��� ���SD;$ly�I �!���2H/�wu�h�F����9��x�h��� ߞ$�ݪ��o�J�{c�{_`�k\C������[�$�� T��;�@�#�(���c �k�T
��1ׁ0�g*���!DA|ke7�A�L�f<1���z3ڱ�oV�]��w",F���H�w��u~9�P8si��,XA�����H�r�0�&q-sstu�
��J�5�b C�"�#ٺ����i�����Y��=4�	$�p���D^zq�l�S���]��;spի��ߺ͉�cʿx�?��ȵ'��NL.��^>��u$;�R8��Q���C>��:i2 ޣD�w�Z��*s�����>�'��!��1$�y�QC���_֏��5GW����Lڕi����XIЅ Ï;R��u�
����d���oe����#����$n��Q�J(��Ԑ��K�/3+�W�}����i�2$�2,X�3S>3��{i	��ƽ����yP(��X���8�m�	�B�/^3Z�̒e��lFf�z���0D���� �Ng��dNn�*v"ܭ�EC��H��N�؄���x�.���l�u� ��6I����������6�wuϝ���C�e<�sE�߳ɬ���+j��>�ȘL�� i�8���`9��m��Yn�fq�;�$��+\C�� L��,A���(��I��}/ �B>�sd2��K�h���c��x!^C��)q��M8s�x��E�n�+�{���eŲ�':�u^m����^�O���؊ո�yo�zU�y�se�b 1�C�����Nz�	^l0���7�N�(�ڗ�̉|(T3B�İ%�n�keL���2ڈy7�I,���m�2�B�.�D
;SZY
�y��&h\M�z�5h�_q�Ar�	��f̓��K��ߧ��]"K�h�ՙ�u@K��U۶�rhK�9�4X�󛭢�BP@���I>e��h,H$n�1̓�\B��yNd7�l��:�"o��"���/�EdcQ[��f�[�**o4)�#��8�A7^��l�p���/��m˜w���x�T�K���`S�)�p�ϸ���K�u~y"u���{�X���,e�4�c�xq	 �
���=/g&��0"	U���� S!��PA;��h��Y��=T�C��?����6�?��O7�� �ٯ�}�W�@��wx>�t�}K�Gq����{z��WJ0c�1��|r$��^Ձ'B����.o����<*��~O�	>�4�.�,��>d��ߵ1����;���p$t��A+7��s�����Q�0CnС-��2+p�ڶ��??`O�B	����^�Gqn��J�N�ݱWݸ=�� �O���A�^)�ָ����#a��2LK[��l��H�ׂ�!1�Q��y3��'=ם#r�K��Ά�}f��|�:�|�_=�0�K>1�B����j��l�0��9�B�6l���KB�H麆sIR����ǂH�f�b���v!%���4�fgKÃ�xI���8��$�D3�1�2��Y6�D�i�A�H��k����L�R�!}P�d-�{Wk�ͯ��ߪ�z:~G��sW��dY��`���O^2�.{��ٴ+��R k���D|}uh�N0�Zh m?��A;]��ޒ�l���R�����GXKfԔ�ZO>��1��e�O�gI:qě�xY]1YDk��cB�7A��쒢]̱��T�$��b��]���l�Z�+�:S-�Vd�ĺX�[f�f��d �b(�#t���$`��Ҙ��ܡ�	�MuGL�5��6�+�7��o<�֩!�XiXˮ.��&"v[ny��X�fMGL^Z�2���Yl��p�[Zh��j�G+i�\m�R�օp]�\�b��fF�qvc;a���ЛJ6媗c���w�H�� �2=�ٿ@rZ�\L�YA�׌�Ax�5�(Ԛr��$������JL(.�Cl�A!]���է�|0��Hr�A�����}��dL�kպ��9.��0���,��lsT�cS�ȱF� @ ٽ�J�o�@�����Ay�w�0.�n�ض�OsDu�h�wDZ=�y�T�/6�>�xbBdz� ֥^d�)��:{c�!��q	�r�>� �ȹL��4N�����&��ooۇ4��s4Q_|�1n�N��w�̣W��E;���Mg;]s�Av�H���Y�L�W T�W6��6_�Ͽ�k��;t���$��p�}����F���l�^ռ/����%i�|2���~��Z0`@/�����U�ڥtR���q��p���nx���fg�x���6f�(���_�O/z�o�P{�-�7>�g]vw��aB�1�c$-{vZŃ�{54� �U����O7\[یmh��EyB�� DH> ���%�z�3��ޕsU �'w�LD�[������z��Jό־fR�[�U1�J��%1 �O��vp�ɖm>�������{v|����#l#�ϋ��q0nۊP��*��(j�,��؀@-������Q�\V�x꫺���`����˶���&�ؗ�&�V=tV���kCR��1@�JX��Yߟ|���z�^���P2f�8s�ykU�S�I�T�`$BJ��q��(D;��9l�y�ׁ$�3v����i�.2@Z�Rқv�2�uSq>�h�X/;i��'s��,�`��~8����� 请���j��0L��ΐ9���j�w���!�p[�b4�J;�)�S�^�뉸,;��@�%��!ͷ������9H��3����0ި�{h�.�ޱ(�'q Iآ�VMzZ�l'dʘ�V����h0;�i��~���fr��0�h��`�o1�"0�1paTTERv2�v<DkۮZY�K}��&'g+�YJ�($>k���6�#�ƚ������fL�N��.�%����L*]�b3>����ζUI7���y���qM��"�B>>�S�WT��gcF��qm�[LA�j��vZ-�^��P�{!�)�P� �I��	���VH���X���~ϔı@��Zg-l�޺�dےL߫��Lͧo�u�d�_��ME�|��T��slK�X����S�1˵���?S7�������p�����rǈ���$�؈$���
��D���>�������:YBg+S������y��^����A�g�%�{|���|ϲ����c�v+�� �=d�s��� DS-�HA'����>h���k�V˻@D�H�q �[�B�{�i�yڠ�'�,�R�=����Q��"�����h&d��mѺ�d��`���� ��6�p���D7�����k<И����'.�.�e�{cƟ^�6��_�`)�p��o�}���\9���y"A�q���#~�L`��.��Tﵯ�qϠk�#V��&Z�+r#Y&�q��c/MA/9��/M��E< c��Y� ��bX϶��8������"�v��,���������`G�0�t�\@�"�v�nlX�����H�0К��N뗇���5��	�C޷�n����L�:i�md��x0`�?!�n~�Z��yO�RuriuWwÇ����"}{�Qx7��kM�iV�/z	�oh�t�k���{�����ByF&Z�4\��J�gsZuG��ZVѵ�Z�.��Xа��)���Éx&�	|�#�1�&��8e���ii�	�RM3K�ۈ&����؊�LG����
7Z����,��ld]d4 ��(�a�+���Rb4�Ю�d���Km)�b����	�԰춬	eZ�̆�v.�8��k�p�+�6SZ�Jƒ�MZZ��5�њj�����YU�(L��tb�6���pqu���מ5\!�ĭ����86�B����VQ��s؛?~��P?M������O��ؠg���B�AS%�Nf`#ƕK[�S�$�"��[[b����wr��3^v[(��2��n[N�pE一I,v�፷���z�Q=�u7�7�/oo!$A�O}HLln?}_,��G�	�vw��V?�NFmF���0�#vv��xQX�	xJj�k�dZ�8ͼ@,I�c� q�%f��*�W>~��� �4��'�$Ͼ� �v��}̋�����L�	�p�	3��	c�����ii�30�db�d�"�0�=Y�Y�Wi�����bm��h�m�H镗V�G3H��;��� �����^�εw�@n��^c�E{�^�a�v�E�R@��В�	C�	Ś�tX�Hk�O[~����[�fI[_N�����T���;�W$1�6܋��8$$�y�x��۷��v�ﳺQ�;�c�:ϰ�!؇R�3��U�l�����8��E��_��������&�JѲ����qZ�^֍�ݷy�>�`�%l�Vc� r�<$��֔^(DA�"����Y��kNȷ��#3�X�˦�����B-��}���dҶ���;L�ӡ�^�܈v,�;��x��V�N�:�f���c�Cu�Ű����6^�?6��z��?hJ��pɖ
�r�aF�9خ#)�1s���o~~�j��t.q�?^v��y<����F��E���O��������=�g����� �����E�x��\�I��Ck$Ũ�݁����e�V�G�k��s�^&#K���ηy�^��b�D%��0o��ˠ�m�2�Q"}Bǈ�>���n�ޜ4{�y�#5
�T�+�9�����������/݋��5�}�XF.3��Q���z4T����%4]û_4ڶ�'��=����4�,ro�Y
�5^�蹱���kn��>�t���5y�|^��y��}��F��Iб��{֌#!�:� Z�Լ_u�|���#��ˉ����>�4v�}}��m]��>���#���#����������v���>��1���f�����r_M���s��{�{�za��5c�����o���=����\�e���sD���Wq�7��o��F�Ǿ�n�L���-�|%���F)WxY�������~�}�'�$����N%�����3÷���}h���)|������z����6p5���ZD�<4��e>�o��%��d<m�>*jݒ�@����f�b���>�?9������c�tx�2	s˱s�L�����Q^�e8��疭˃S���v����'���O��E�$�kY���O5�Rdj&K����;�_��ܧo�r��œV{�[��Y��E�@.x{4uY�M���~���0pf��DHt�hC1�-� �yB���p`ᒛ0!����#V�	u[�����m���dp�$�g�p�?0�������5Y��f�����~î���B�Q��R\kB�c2̞P��LqG-FT����z#`ɪ�D�zu�������_]u�\qל����젹o�@�|K�&e�u�Y�������e�Y�Bɬ@��A�n��u����_|u�&�8,@F,��ɨ�|Z,1��-��*3�����������믏���������8�r��}f$ĕ�z�&����XQZ��DTPDX�G�ԛ>�T�b�Og����}<��뮺믏�������8��s�O U*���qQ�[E/�gwTV"���iX��S%�H9a�����UڿQ<m�]N&3-��ڢ�>B����
�U8Ԙ�g�,f&y�'�8ǔm+
��
��E	���Z�!^[)E:Iۏ-��$�Y�U-hT��J,įI��T*[R�x�A�������T����r��Ĉ� ����\B�b��V(��yL��j�����n0YS��ћ��I,��,� O��������5���{�9� �!X~�݀����=��'���Y@
�q���rc�O�0��8�Ř"�~~��N!A���J������
��2Ƀ/��۬��>���@'h�>�h��w�ԇ��G�4Zf���5�_�݇��G���ߦ ���^���YsP�� �x�,!}��N���YD
�����
)̈`k�	!�a����V�r�w�����J���]�Srݿ��!���f�e����1�ڰΰB�2٩ѵn�[	�Wh��߂wrK�[CY`> s#��²Ì��d���߷H�:�XA�.CO�0CґalXte� ߀�'i&�O?y�9�A��,?�~�"��Z�^�Jֳ�(xSD� �0?fD3������|�� ����2q
$�8�'Ԙ�>�9�)8¤��Y����7?����� Q���h6�Y�i��#����$�k�ÿ�����s^�Hv5����Ñ��-��B�|��z�jB�;�,Θ�u���<C1-e��r�E�Αd8��Q%�����+
oʯ�~�[|]6�38xJ���Ny��L3�5�3_i�Y�����hY�0�n͌�i�LG~�/�y��
!�(�v,��8 @��\��{�>���.	B���	���Lz�ۺ���������F��v�=}�y��}��G�̩��<>
� N_�7�mhdɓ&Me�YK!60+ ��y�E?0)d��2L8u	����&,+��dAC�%O����2q'�}�/�u�C�²��Fs���F��=� � 5��6���m��9%�ÄH@6�:I��<��.����lv�w�cK���J9 ̅4r�����>���7�N�Jt~ooOd(ʐ���n������!Z�dI�0`T���C���Y��wϳ��$Y؟���J��d(���gr0��u�g��3��{��I�
�w� Ia%�f�ѝ�j郸��ių�:f0*T%J���ϳ5!����	!����P�,.%�`���U�?q��07���
��*X�xRw�h���p+ �R<��A@!���dXH�>���4�S����V%aY/�����'"�݊�k5�D�3����t���'&v~��n�׿E�_����}���~� x��92���R{�5턭+��ߴ���YXlI��:��?p�!�Z~�����C�C#&�
�9߹����U���ӳM�L�Ȥ�K���@� �",6ߡ�������Vث��H�T��:�H~�K���[a�d�D���Cʐ�S�Uh������w��b��4�٘���]hbQQ�F��ej�^�X7��ʹD߳}^�0�ߦn_#6�ӻ|1,��2���@ �4�mf��)<ק��ʰ0��Wʹ-�7]��4���lV4<��w�8�8���>������H)����@yɳcu���3J�:E�B1j���T.�-�&�:%6��Ey�E���CFj�L]�mql��0p�7I�X�{Rb�Z�$���L�kHLt�ѣ���mځ)�\@�T´�]�3,+c
��.�M�!Y]bX�GF!L�:��vs�}w�<��ٯ��;��>y&��2商�����8sq6Z�b���p��R~����¥�A�}LW��N���Q��TK������ƫ:�ݳ��ב(�I.ˑ,ZJ�O��<w��=��u���A���1 �|��%e�-%�s��d�aE��~���0��c�3��]��* ��y*�2[�Ӥ�ĺA �T�������6 |��o3�����u��	�gj�T�KZnҕ��1����,�]��\⩳��جh�w���p�0L�H$�fLH2Jd�ϒ��P.]��[�ބ�H4�Nx���	u@�(AXs\�^ ANdV`W��] �$�����A͜���(?T��I�[�ւLxy��$Y��[�/<��o������QbTܒm~��p��p�s�˂�*[�29,�!pGmtɮU��~����J��	t�%���:�Y Ht�D��w<��̉x#�ɼ��p(�9N\3���k=:y$���@�.�D:�xS�zT��k�N�`2����.�Q����#�2c|NFVN��-�\<
����s�±4��j/G�U^��~���:��J{?O%��Ye�,��$���ϣ��y��~�!'d�]��x&R����P���0`0 "���4��A��Hws��-��� �G�e Z�������9��@�Y�O`ݸ�0�'g^<�%��E�@ �o<�)3Vy;��A��@*����;]�����:�'�h�ʾ�fU9��<D��x��H�zFH쨷�Mvl<��>}�@2&4������9�0��	n[˴��̒̉ N�%�>I��zvI,�@��������k̤�'C�m���S�	A&}�'_�����5-���6�LM�N�	/��X�n�X�fi�LZ:�\)�� ���#ݧ��%�� M����H$3��+�z݆��-g�J��L�;��za�8���3v�� ;<�V�gxK6^w=	��
!H�8u@z*.Y��bn}����M�o?+�@:��%�/2����	�a�N�ē+E�W	a-�Ut,J�g��	��^a�J}�"Q)/v����bi��	��'K�AF��z�L��{��qG�\����^Q��>/��ex���3�#3Dy�<wq2�\yF<�M�z�l �Z� �2dɓ&L�0L�U�B��J�%놉	 IZ��DH�p�>�N!��|�U���&���$�KYV�隒	��A@D$�6D�I%K�y����b}�]�Nk�';^D�j��y�8!D}�����H;��7��$$uL��W�vְk��<4"�/���W�"ZQ$�guE ��o��Y�ݶ~����X'�t����F�Ԕtf�)��V��m��3Rms��������YCM�[v�<����0NF�bh�I$���i�V�{�k��s�Ds��V���($���$JV��$��S���}r�H%ޯq�P޵�6�OO�I$K�r&Y$�k3;��1(������&�-�Uw<�M�D* ��yK$W�ͲX_lKJI ���N��f{^ ��H-gv}�+Y8��q�oO/L�g�&}��
��,�;�U��?N�e��w����$|�fęI&Ir�R�H��?��C�Q??���v�����}����ꑐ,��)��Ԏ}um�2a�{/�T�i����,���ui��݈Zt�.��8��_%	b42dɓ&L�&MB�/V����^�TS����|3Wq!�I�F�I̑��iw%׼O<��>d�>�+��p��\<�IdVw<�՛��w4ΐEZmJ�%����e�qڊ"J���k�[*j�j�����|��A��:$%��ӻ#��Z)�:��4	��d�����oO~�"y�=���g-��Q�}$��T����d�{�rA*��ȭ��^��G��/F�4��ْ�g��I>��-�4Δ�fA���*�l��	����$��S�&��7+�H��P��uu�@J%s��1Z%���1� �Z]ML�I �s̥�l�䂡
p�G��3�LAk���d�E�l�$�M�H�@$�w<�@s��3�V;g=B�D�gw�엖@!4J	]{���;�1œϲ�D�:$�p��)^TP� ���ޗ&ڀ�C�]��N@%.���.�*�������d�'�dhq�/z���TE;��,���u�Ϸ v����\��/߰�8�f_�"|`(	�&B]l��X���E�3`��k����v��-p�:�y�W��np?NJYe�P�˛�*~~]+�G;6ʤ&3IYf@�SklBc	G#R���BݰJ��*ݨ*�bPچVkU�����
�-�ZU�7DY��T��1��P����tMH�l�2X�00Q�ێ c-�%�t��藿ØyB��-��l--�F0c	�6b�7Z��2��6a�q���%1�d���/������M�����Ҕ���s�f�m��ev4�<�]��"����ӹ�Z\��Ѐ$;��(��n�bd%�bU��,�3�K+y�%�$�;�{�uUv:w$(��68� ,g���s>�ܭ`��=u"@L���*��%��&QT��8H�^��&jBO\Ef*u��a�H�-�N=��% n�1�I��=�q�N ���z
��:A ���(���H��Hq�w���%��n��v�Wfw{3�,�ВH�KȔ�� �BI�vXL��IޘȰnm������׀ã$�S�Ti���H2�) �wD�Z��U��`5&n!���g�Ie�̤���tșLX�@�tĄ��� �{�=�&V0�_�950����hER�D���r���GFj�p�e�&W￿>�f\�O���~k� L��8e��s�u �ݸ~�8�����|l�2Gs�H�,�I�����b�=Q1��NL�H%=;op�'���[�7ǚZ�v]W�=��4vF�-�vk�xe )�uH���67'O{��Q�aN���dD����p�!�&b�L�dɒ��J�o������Dʙ����i�̕��*��k���K�Z@H$��`+] �xc~��_D�).gw�)%K� �>]�u�mv�4�e!�AOl�j���w#�"))�N��D�Ow�¤�OV��0����Qq �RC�;�g(�lŵ;�A/o8�����s�U�r�H*�K3�ܱ�%D)Ͻ�C����H߹�Vﰶ�1�$Qޑ$�H��`�d�*}�y9���J�M�D/ ���AO'o�����t̫���a�� �K�ٝ�>~�v���ZI�Tp L�N��
$��x���y8���7�;�x%[$\e��98�������O��$��qW�Uжy=Y����V�9���~��.�s�-e^hz/}Ys��4��<FM1�0��uT���2!%L��z5�	P��Z��+�C���I����2�1�D�s}��ɣ��^D��h��n��TD���~���F�~��;9s��0���Q�Y2d��Y��5�SR`Ny��m-����3��P��w�2���[�Oj��wC�i��""�7j$����I�+�y��I,��鳳г	�������:�r�,�(h%�o)/�RC���v<�K�ܟn�C)rdN��s�� Y9�yI$Mw<o5�I�Savw�u	L�d�;����(J����$b4�u(F��,D�8�c30+[n`(�q�Z݁��7߿�/�U�q��Ʈf)#~�����,�]��ҕ���l���� I1F��2����	�P�8uF�K�� �@L�����H�D� IU�̤�fwwޑ-(�J���C��c]�������u �P<�֔{^��/vă(%�p�<���C���`�7�n�zRL�=��I2�v󉔀Ɵp�>��ч^�Pz��<&������5;��x �3��;�D$�i�s�Ʈy\������{l�4W�E�X�C��S�E�}���	H)�=��rQ������6���ň�1�~�_ï^�x��ׯ^�e���� �q/����}����)������KK"� ;�0�pD����:YI%^��IB˹(���?u=%�K���U%�';��-%vٍ��cc�61�����[���X�ˇxr!�Ɉ�2�i~��B�\��<� L���e$J��/) oy��gA�}`��Y�S̪d���l	i�Ȍk���
�S��[��1�&	�L���uA��7�/�)$����RX���s����O��%Ė����Ť��7WHTB�	é�	���~�H�d�����"Ik 0-JA�@y� ��T��2D�ɁI3��$>$X�W�oJ;�x���/7ŏ{��_��^5��� �:��ڙ<�3�ϱ�QX(T�ְ	g� ��1H"�׃	؄BwFF���o�1& cے'[�O�a=��0	& ;C#�K= ;y�9<�V�H�̀Bo�Ӳ�������!MF��Psll��0{6&�V���(�=	@Z|�Y�����b��/d�������ڽ���5&/c{Y�h��&Y���ã�;�w���we���qʙ��ٺ˚x�����O�[���G�����큮~�s^��G^9��}����n<��[��u�W6�Ö̽KJ�wܸ?U��p�&Hs��xw��n�z�+5o�_d���F�zx�Z���<� �����Ԝ��YǍ�0�e�����O���|�����+ˇ��f�xR6�e�ǉ��}��bí
�ɔ�d�b����/w����v*
�(����w��R&��n=7w��#���ױA�qg��mz<�{�H}���p�:����m-�=������ݽ�s�>��zp�o���Vo{D����0ujx��N�_k�!�l=������ןb�V��3�8�g�B����չ.�RnjEg�' �7����[���O��v*�ǽ�����'���ʶ-��m���	�CF�8��jZ�{�;˝$X��~�����:��{����v�\c�Gb�<&N{���&eh�����wT7�z��=��$},�*^ܸ������Nk�����S;�^�8=x����)��C�'�Gjh�]SV��:`�%�,P���Y_�c[��I�jC����_�ۈL=��I�b:qg��6$���A��!�F��W�}K$� _ҡ� xs�4��&�WZ��T�s �ܼ_��.3^���4x����^!��	�ǘ��v։�s{�q�N���,(���﷗�u=���g���5���c�~{E����olOZ��e(���h�#���2���Z[��{���9-�i��7�������[��~6�
�<���f�	g��A��R�(*��|�[�>���3oO e:�s-�7-�+0�A�����~y3�g3�nv�yJ�=�=�3��8�F�E���L*���J�2�E+RҀ����[��=�O�S��~�뮺��_>>>>>�`�"*T�e8�QB��S%E�ܢ���80*?[��I�Q�/O�������u�]u�㮴�}>�O�S��2}�p��(��rc���\2�v��y����$��t��A6����w9;�O'����뮺��]g]u����e=s�ة�T)m���9f���QE�Z�ch�%A`�b�[;�Χs������]u�]u��뮺��^��ұa��)�b�2��K�E��gG9�9�xx�c%�6��ƒ�*	l��OY1>k;j(z�"�%x�|�2�Y6� ��C�j�TY�}�����T��E���偈ca
����fʤ�IӹQZ�TPR�t��i:�d:�:dԊ����%j;aSY��DYr��j�ŋ�E���^�eH��"-�;q'I*
��jDG�L^a�Rw����\��{�>��z�%G��o/��V%��5��M1wF�l	X�e�n%�rA�Եkt���2�]l�d%�Ib.�6:���	�L�M��4�f�:�A��P�І��S
�3��V��l���l��YN�l�j��k��3cfs�+��c��L8��2X�����u�+q6�8e�C,5b�-�7k�Y�MIbif��X"��k.�`]��B4e[�ae��Τ]�f���]���Ib*b�h�!��̸e�^�"ɢ��ݫY��u�T��R�K�kt�Ѷ�*��$�b ��/j�*�qz,n-a��Y�#,�d�\��-4n�F��5Ux +A�mRT��h;X�̢V��mе[�uiH�Y����[�5�9+��Dy�R�������m�L�F�`�:��4�K��mݭғ���<Au �&�R� 2�lm ]v�̩�I�����Rƻ��hE��͋�-�S8��Ή5��K4ܒ�f��r�kW�.��l���2�[�фáw-��b�we����f��%�̎�vr�dP��s�e��4��%.�X�H�PF�k�Q4�cq�v�n"��@t�(�Vr�˸��fm��e�A֍�c��36+e:�N Ǝ�K,v5A�F�I��f`Y��e�۵ը�lq�VR5�D�m�-ÙE�Hg��^rj��Jn��F+
2�*/3H�RV+).�4��&cF�B�D�i��g���]�m�\��B��F&�CZR%�CR^.����ɰK5�g�q����X8r�+�7-L��@e�qKq��+�1HP�̽vH\�����ٴ�Wer��6'��|��[��_1K��l��Q��O��z�
�^����G�uG�z�^�zz��z���)��~[>�B�qh�m�4*8HW5͘l41�˝�	FiH˥��Z]��"%l��2��Ը��li���V�+,J銭�60��L�)16�f�ln���]95 ກk��=(7ZڈF�ej���Gj����n�h���J\�M�M��Lɘg%���W:�[+yLK���\������g!m4\�cf�KLْ�c��aF���k�������p�%��>�Šǳv$�d�otSP�������@�JeM��4#���|��B�V��K�qd^����5�M���bX��ɐČd!wCH ��C��I�m��"�@���� �23�\���ld�g���h��Ž`1�p�p	�p�.deM�̗�:$Cz|5!q	BN���U�(�{u@��� N2[�>�X�(�ٝdCt���D\��0��p�%��$eO{��҈t����r:�q���f��K+�"T�|�� k�3�(�gL�k'�����9������oP�(N������;#7jh�F�]m#a�]uٚc+�f�d)��~}���@I;���Ѵ�!�"J���������8��.������t� �X���0���:A��h�s�bZU>C���66���}�:p��#.�{�FڟSG��C��?�ot��{�oW}G^�5�3�˴�Μ�>��~�a'_Ǡz��z��T'�^��Z��^#�s�~�:��̑-�}�� =�����rQ��� ���W:+ ����^+}r$�Hn��	$^˼3��㧛ʘ���	���@�t9bX��s�
�S�\7��6����Q5-slX0���䳰��Y۲^�y���ހ
zy\�}V����zZKdp���%	8w�9>Ba%��l��D�3�xd�#��8�[��4�葪b�a
=x|�^(Ӫ���-��nY�� �2J{X�R��֦{K�L\DF^�'u�˼r2�]�������q �	��)���R��2�0� A���cD��h۲����v 'wtb-?z0�Y�;?���v�O��=1�v[�$���$��+FN��b����G\��xcv�N���=۰�@9�7u�b�Q�[����Yr��zK\��� n.U��[���Y1J4j����r���A���_o-�2�{�1~zo��N�z��	����z�A�B+\�����)kϠI �z��D�O���[�9����P��0k+Ƞ�A�K� H5��K�Y�{l��s���q0 K%=�\�S�*k*c�P	�	���\
�;�{k@o1v;Vᵎ5g?L�e��uH"j�,�k�i9)"`�]"_ g���72�1֭�B��\J��lx����W:�����_�vmp�b���G��$y� L������l�w�tk��@,�O��d�wS���NS��G��ME�C��|`ʱ�dȃݽ I$f2���y�:I=q��zݽ�I�
s��(���#TM� 5��x��H��3���.��	��7��SH��;-ekzd� ���4�.�3��Q1H�{y��=o����`�[�B&n2df�� ����=8;o����|c���|��ǽ��g�Q�
b��H-�*���?p�{��O<����,?�����?|u�z�ׯ^�z�꽔��z+�A�ZEh�N�G������A ���I}�ċ�?�d9��q��):�L-�k���2e��f[�݄����Q ��れ��)0eз;K0.	ue37B��ĮT�kT&ҍ�l������a����~�&m�� S��A,s�刿d��;7 ���mjS��"�BE+�VC�x)þ��<��m���E�k���Hb�[�0[7���I.��I�3����MME[q�cu�n�
ܧ�b�w�@�#��I$
���l�p�FA����(��""���@N�#�=�Q8��ׅ����Y�H;��S�e�Mޑ������'��"H�QH��Y�rF �#1�p�Љ��w��7o���8& ci|��4	3 SK� �e�kS)�G���͗�#���ˠ�*G>�4�/m�R�{V�!i�x�ِ��>>}U������6��6���|.���Y�7�Ь�7�׏�]v+/�g��، :!,qk�Æ����#����gS�UN�O^�G�=z��ׯYӹ����~�i�Ba�]Q�l2̧]����N�ڕu��G(f�E��ܚ�F�,��m��֭% Z�(�\�t��e����ۦ��[�t����-t�m�M�����cGY�a��]�C�eZ����vR[[]mBh�Xav�a5u�ڠ���D�3�V�2�Eo]��nL��953�m4��
�h�4�3'9��"��V-&
L9�Β� �P�7����ɇk�H#s�.ҭ��އPf�ـ@�&X��Hk��b�H����\�� �;/�<��7ܯN/֋k�jd>d7^��,<��r`6���p�d/C�x)ýPL�|�q��,�����!�� ӏ��G7���u�3���,$
$��ws��xLoYV����+=�T����k:n�O{:d�k8r��Q>�'=��&3$�;���\�&"�<^�1��ff���s��w��1shy� $�A*�r�D�~�H;u�ռ�S�� �(I�C���P�%I�Jlv���-�(mi�a��AУ�E�_�~�~R�P��&�{[�d��b|^��� s)��^O����o�Lb
�s$�W:J��\C�v���bXT�q��ߴ@P�s�v,���Ӛ��_�U��Z���ھ���I��izkh����<���p�IG��)�wE�������oؽ�dy�0f�����Q�S�T@�Ǩ�^�z��ר�^�z!�0r0i��2,y�덉 KS'?{�u�g=�� � ��@�H��>A@�|ɽ���W"I9=� <+�z���tY9� Mvô�g@���	ޠ�O����A���g���?�o���&��,�`�[��2$K	�1q~��lhm=臜.��Q�t�0k`SH���]�����úr����i� ��Lz�}�q�<���+=1$�as�N�8�)G��`i�bG�j�8b?f�Q���k���5ԬKv2�����9vr"3,H7���1|�v2D���v��[!��_s�cCo���6�0k
s�A$�tSP�LXGC�ws�y���I�e��Kﾀq;�����)���þ��� c'�"��>�=o�)���C��(��Vc����#1خ��vw'����	o��)�k��
�r�ky�8L��X:���{Jyd�d�{Ż�"������܎���W�o6j`�(�xfU��F��?�����v`��'�^�dJP'�^��@��z�!�
)��}{��Ȋ �[{�_�&{��uA��_�j)��j��o[�%�eL���"	�7� z}�
�8��l���3����l��	�:�h���H>���8y`��=�cf�H9��� �Ι�͚�M^'�� ���81����������%���lɝ�JUZ��\/30 3\�`d����\�9E<�4ܯ�2$6��I�A���
#�5{Q��{�3�6��	v(�s��Z�6.����]1d�T���nja>솆�\Â$�L�)2_�����ㅢ�:kC�LF0j�gLT�&���Ȝװ@ �%m�: �!�I]|$ǧdL��@e=���F�Cc,��$!�buo	�F*�wNà���1͢H$kHg��02eW��%�V/Y$��tWfk�{�,,��X�U ד�K�O�W�����@�{<{�g��c��zs�i���d��0ݠLQ�ev�v����a[����~"�_O���ׯU^�z�T:���{P�)(����� @ p�ϐAwP ��g���,��;�5�@�yO��<;�mi���ZPvt̂�����b��-��($x��r��j?iJ���s��,4�3-k��L��-	c١�r���v���ӭf�v�Uă��;_>K���w�NL`�kpĒ`�������8}/D������Nm�(r�xqL�� �q,�Z��3���5�����u�	bA��ơL	�m�q`7z��l�L��͑�"�?OKp�[ˢ&�H5�*=�9��[@g�;j�d��fIb£�dނO��	~h'�6�l���z�`��0��K[����	$�{2�K:}���(~�`�H���9��p!�/Z�$��<�^r�#�����-SY�z�`�$>�u�� ��Α>b���e �P����SＧ��a���E�z�ǸCޘ&�7���^�����P��'��zE���]#�G5I�t��9=��pIOY<��~�[�Ox��K���C!�^��o��z���k\L�s�W�9nf]���� �g^�;
ׯDC�^�D�u�'t�_���4�͎
�&7�������6�Vf��AK���Z��ŀh�fN��a	CP�t8%��R����cH.��JF[�"�֔���5�)0��,�%��4�B!��2��	,�1�YKs(�WB���[��e��%��f�5z�0�h�h��.��剶v�j���9ޚSM-v�"��j���֎�ɂ�(N�Ò�0�w�~���" ���Y�5��7�>d��XE5�M��^�B3��z.�H�H1{㰠��N����^�O	ԽDa�p�z(��r"|��t�@�j� �"�f�{h����h��!'�t	���ۙ�A兄1�p�ή�v���$���%���C�$�p�C�1�`CG.�ٿdfE#pGGzXkV��0}Q���l�}ޚ�3o�;��E�H��tεvR%���W�#��,GglQ���=�/Y/�S ��D��� ����A���"Н��	����h����_yJJ�]��.u����L��(�� g��lBt!��DL�+�m�< �(s7���L�;�a̋ �wl�m�w�h��?�]4��"A�Y	�%�z��A�Dn�=s,H,�@�>l���I���De���4��Ъ0��mQʨ�x�k��q��f5�t8{�ye��Q�I�S���^���	��o�<(�*/��Q����P8�=EN�z��=z�D:���;"���;�� �	[�@�M����[���W��w=Ѡ'��5���������ө.W�ױ8�vX�X��Y�!�r�|ؾ��%��nt	��8X�BO�1���������z�����@��S�P�4�n�L�z!���[���s��A#�̘H��RJ����� b3��D��8�:f���Ž��%����vL����oCx�h��a�tQ,�v��[Z�q��l��@��-��J�.�4Ơ��L��]kC�b!p��,�	3v$�I���$�mfآ�"#����m��hd��� H&'���r��1PԶc��������ק����ĝ�&U���NX�A��LP>��՞�os�I�� ��Vn.� �����jd��t̰�Ah� jv�k��LI�tm�۴�7�X�{�+���p�v����m$��*i�Oq��j&�� ����?oUr��1J8�.[���&m�4�F^=ϷӶW�ɨn	�}�ovG;EsE�KZ|D�ù<Ǖ�r+�L�s���$���������Ӄw�����k����|��:^���g�M��p�_��9�8��݉���7��Io����:o��ąFt�tw����wӚǽ[�/xȯ�l�+��];����Ӏ��.��1�d��e�~�'�m�-�K��q��om�7/��λ��Ɂ>����{�H(6�7"��.�e]T�Oj�����H�nM���?jK��k�J����t�K� /���g�(6�}�9Ἧ�9\:��G�d���;�7�5��n�����1hFZ��5+��W���A�ZV'��Z����{Ɋ7�8�)�{����t�to�n�UPB;��ywy�\Z��93yr�m�������v�MA��1�C���{)�Z�����ly��?"q�x��/��m���=R�������tug�,tw-���_�����f�������Dn����o'��v� �����3FB��K��Q�G��=���/n�_�n���y�ӝÃ��ܾ�`��q���:�R�|j��9q�>*k4K�'��٪1G�[�b�0�	�2ѕ����=z��βv�P�^���E1%b�V�����R{�᧭�{rbzд5��{�ɖ��D�i�{³��t��|�2	/jr��i
����4E��^FO��I�8!P�d�P+�3
��EH�`��o�}z9uX�d��A˔Gy˼R�?��_u㮺뮺�u�u�]|}��8|�NAU�ʋ,���`۝�J�b%�Ϸ5Q^P�g�k+�S���z�u��u�]u�㮳������̝\�AbȢ�'N2bZbJʕ�۩��XԬ�mR�Q�9�^u��}������]u�_n�κ믧�=��p���n\
�C��,(M����U�l}��)n�l��^>�}?_u�]z뮺믷]u㮺�|c�>���˜�=af�5	�X�eQE��E�DUQX()��E�&0��X������ט�F[�WX���b|�1���5.L�1&+㉈*���8��U�9k�V"!�0�R��jW,�E�|J(��������Ԩ
�`����QX&[�f8�
r�H(,�/|��0�=��5�$f��,��-y�E[�Jµ�mQ�DUA�o�+&+`�y�Q\�oE��/n�O�����XcX9�ח�[��n� &����#�z�� ��ע�ׯ^��tT
��|�?�'i,�;l��Ɖ?T}>ҒJ����A0�]ө��r�&�lx����o�F I�vD�@!���2`{������ĉ��F�J;5s �@�B9E<	칒E��U���ĕ��` ��H�X��Ldn�r���6j����!�o
�W��k�[���ڍ��S�рѦ��]rA�ZC�8uS��$;� b$[guz�d��Aw+<�fX��2q���<�>n���x�d^̒� ���&�JA*��.�At�D-m��Q憘�,���J�{��j�]wHƉ�q�1FuQG8:���5��x�b�T9��oE_CI؍l+d"�{|�=6jf3�H=;��@�`�u��گ�
uC���r�*�xzA$�\�c,�3���`	 noO�xױN���A�UT�j��hU�:�{ϧa���/��_�bE��uA	J#M�_dNHk'�f�@s��Ç�
N?�D�^�P�z�z���N҈4
�XX}R$�TjD'N����&�u�nW���	���MA{����-�],$��წ�d�۝41�}�?��R��1	}�h4�b\-�afhYwe�͠��ˤ,b��DD(�A$��:6	�(���[��ِ�A ���&�,���4��:'ygG^���;����Z�c%��,�����Ս�Z�%��l��\����OU�H=�65=��[� ��ЫԈ��Xק�|՛I��
��5�Ћ�v�i� ���5;S�y{�>��A#��x�Q�4=�r!9EC���=H�P��ܒZ��2	+2|��ص�,��h�	��l�	�B%��\I����
uC��w�4�d.v������M;тX�}��6�z����<A�0��U�'�/s���INA|W9���2L���xt6o�I����z�K2V�`bg78�,�þ� �/�k��*M+�P�A�M�G%尾8����,e��{:]�]�}W{��Q=������ע�ٓ&!�&L�I& C���{ih�9f�]�\`��cs2W���1Av`�c�j�7c�\����\P�<��cA�B^�dv���2���d��Ʀ���*�)n��=i�X݂�ڐZ�t���ǒ�e��^�鰊FZ��HsFS1�����#,���H���b��.��.���l��*�[�`�Z�Vն;���-4�5x�b���.��v��8����?�@�N���zS&R�=� �IR[�&}<��􈗂Ù�wFŀH��I%��� �r��8�^�I
���GWk-bM?�$�X��H�[��rꋿ+�65����r�AD������$�<�.��iv֦x�k���~��ڽ�2�)� ���&ᱠA=�G5{)�� ��ŬZ�SU��s��d�K��	kd��� -���2L���*�x���o�H	���@�����T9�o�3�2I=�a��XD�6e_Q5p���>�$�F7ve��<�5I�.&($�+�УYcU���!�3�&�\;m�\���(&�ۖ��i� �O�t�WL�LQ}ə �$� �W$p.|���b/ �z�	� ����>~�:`��Ԋ� u+��L��捂��}�ީ�F
���3� ��dd]�O�8��$aQ[9��|�aJ��sF������ښ�~>���<|���z/�I=g�
�q$�A��Bv�n��T||��^�z�z����ע	�RI��g�����u-a��������w�$A�e�z�u������`�r��9w�]<s���j���Ar�s�>v�	w&���K���7�D�{ �"D�y�z��f�۽��F{h]�kYY
�p,�
ʌ	e*,�W�aŅh���-Tb[�Ik�,�[h����X
�Fе�l-P�-��:�y��v��I� g�+�}�C�6���:^�\Y��'��w�5м?!�6'U�`r|ɐ��'�udjG��D�	d��$��]�@٥وL$�wp��w^Z^L$�c�LJ��`����+P��5��а�m&0�Ϟ�z�[�*hU����� � ;{�	4��m���s��'�@%���j0��w�IN��q�����i�I����w�uw� ��{0q�&vH?u̝cNb��2,�S��7��<�Y�
 D'^
�C ���޹� ����5�iO���7�\ؚ���t���Y�@�E\Ҹ����b�e`��j������w�_v���E� 8��'^�z"�z��u�ת����<��?GY"w��Z~��J�IZy�Q��tn��
̤�a�^� �Q�Х�	��f�5"u�Q�,�{B��1�s���A7��]^ �} �"�}���$��;��rr�@��+�]��<2l�$���^/���OT�ˑn��-J�� ���v|�u�6ƌ�˕�����n&�*�J��"ک?��߳M�:̧��=~_��&^tH$s*tc��H��z�s���dyq�����lI#�E"Q��[����H��W�I�@^
�=+WFU+�h\9�ȗ�jL �z�|�z�[�W_��*�7}g���3���g_�]�C�d��k��@~}�q�|�V�yf̐1���)��3��^`B��@���%Yi�Ga��6���O��I�
۲�-�,3���A�'�p���"K������Z�U���7F��� �uz_g����Ƿc�c���� o��+\�C�6w�s^_ag��F=��� ����ׯ^�=z��ׯY� C3���F��H%��??"��:x��C�M�Qb9t+Q{yVr���p:�g����Z�s��@!ש��~���X�b'햖�!L�:�m�ҖUθJ�v*�[�Ι�L��>�&�{ �_�=
c�x�%=2$�s��"n�=צf�
��!���&OY �f/�Y�<�,@����K�_=�c���C7n#e��֮gDˢb��MW��Y$��� H�"��D �(s��y���,���c�$gd�Q�S�l@�b7�A�ފ2��$�Y�EJ��Y�膮�gOW�fc�M�/4�m�g������%s�����B��̲ni�Z8���b׼}p �A�����b�ue�`@�wӍH��p�n ��ɑ�����������3D�tR���c�{���k~��sz˛�z/m�;��v�k��d�;��{՘�2q �0-�:�*���V(�̈́˔�f趗�57[S�IO�稧^�z���ר�^�z ���|)>��k�K*�=FU�3!Y��1�c��j�B-I-#� ��`V��R4�����G^�fl�8���d�p�e��dz���r�����]�Qt1�[-�	��@�ۡA��DR�����9\i�bW��^�T���v�g��[]i,�@F�\5�b���lA�5,H�gmqH8ȣ�l�0fT��mJl&҆%�2�@�����ٍ����}��b�u]��*���>��w�s�'Y}�2�'��x�]�ee�	��C/]$:0��JޘÇ1�S�	�X��,H��%��
`\`��۾�\���w/�Y�4�Z�g<�!��^���%�we��=���2P�eĐ[,ވ�[�Q@�����%c��� ���F�&H�S�iX�on�H�^�[�p��䓡�*�aps��:(:P�[�\����'��{��E�F�E@�Xcq��cL����U�P�C�ox@�;�nMrKv���kn��ª��K2�,��lL���M͙��\��=�ϣ��;_�|c�<�� ��ˉd����Ǧ
��MU;X˻�.� ����wxxN]�O\�ˢ�����u?	��W�����C�ӑ��Ay�e�����Ӯ����v�T��םk�g1�by��x��ϟ3�y���C�^���Q�%=z��^�A�ׯA�����1���g��Q���H&'5���y鱆(f���0 �z߲�	d��Aw+s�a�2��}~ޚ��
q���vd	u�4���БI^��r����E�{2{�^�{�Q���id���dG{���ͬ�tC�>]�}�$�Y�cޤ�"T�v>�C�IC�������x=�<3ۏL�乮�bﾩ4�c�g��,h�F�@�u��"v؉����t�wOe;�%<`*��y�w�s��L�u�+�n+�;AB�_�Ͽ6�֬�{��s-m����)�3�}��!m�bD/u�m:ԉ �_t
C��]�q	ם��y�=8�_���ǽ-���}�S$H�����ή��[K-z#g�<�����ŏ�M�H-l��y �{ǽ|��V��z`�/JiU\{�.i?��x���	���"����:�_c������z`�������&�'Ǫ�z��^�zׯW`��fa��B����#��ēV�A0ǭ��nF�yF��KuT� �M�9b-����g�;&Iư4���Ɇ�R�r������������W�'����!�6���nO���\A,|ŷ���.�[�
�T��C��nа�\2�nHl�͎˭�Vl�1v���
��&��kG[��(s8me;{���A$��#=�S�z��n}�-2�*v���aD���FW�t���dS;]��� �l�c_�S���+�]�nx�B	���Hɔq{���ܫ�?���P� V4������l�vz$�����	��쮌��U�$e����ot�P�"R(n��㹁S�`��ˆ���x�#J3o�m�݋��0 L�U� Ie���?`l�e�����܆zL����}M�|�>9���l��Uܸb;����:��NH�w��^���k*\0Z����.R�߅�D�ר�z��^�z�ׯ^�����0�L|7>��A8�0Č}Q��I_m�;�k�j�]P@	2DOz�A�����ѵ�u�=}��^;�?��n0�T���[-�lVZ�F%3D�MV
��V��r ���+9����׊ke�K#{�X�h�+C3c<˪$]nȑ�	1Cq��At�9���W엷�!����p�$wn��PE���4�A�=n��/�V�|�Q�	�t��Q7~n��KK�d�)��謙���0<糘��a�d�P$@]��k�r�ú� ����N�G�u�ؐI�� �����-y=����b�S>d�Z�s��;ĵF��A��a�Q��~�HOz�;K,d4��hi ���!��( �0c���ڗ<{�iI�#�<��Q��}.��>$�;��{;�┉��zz�(�;X����s�"�_��_wk'v��r������<f��2G�W��a\S�ܜR�Mtt�8ѕ���d�lJ]��tz�qx�ꑗq�z>���o<�^�{��n��&n�L<1��g�3�ۃ�Nw'�h��mJ�������ā�u�)�8����okN��}�[P���>��M�$M��]>��0yN������{&z&/b?!*�ogZ���� ,�:� �Oo��[�|�q���qǧǧ�i �/FK�i�������熷�윱O����O�Rb����3�y]!��
�%��X�=���:��7���J��ի{&F�����Z8h���7������-Vjd�_��GK�����pxz��,@5>���oހ{|�����n�8�����,�P����{/#+�V�o�3xg�5#��K��dA�gh{�{��S��Z���������\�]��k�nm���u4��F芄bc+�#iP�c�R=�Z�;p?,O<���X�6�����񷃣�5�Α�3�C�������]
�}a�����ͫ^�|���N!OZ��X2c�f��f�6*�{�K:H؟���iMd�_B�0׋E�O2�3�'P'1�2`�&����X��fh��4�4�-DKԖ���Ë.�ލE�3Cd���_?h8���SM������s.DJǠ��kz*�m������`i& X�k���^����"�fժ�R
�^��p�ƾ#��LK|��� p�4`h�>���ɋmԯ����C|�f+r�5cue�±#ea]#��o���>nb?�3Ė~��2ў� j�tT�_ѧ�{uĭ$��F���֬�:Ž1-�wKH;6-�������ɥ�n�35�p~�����*`ı�?m	��O~�<�[5u<�<����6��Ļʆ�Ua����N���K�J2.%V���6�[�UQ�׻`��C���ɯ���������]u�]}��u���Q��	}�^YU��q��iLJ���L�J�T�$��b*�9j3Z����>�O�s�ӯ����]u�]u�뮼u�_A���R`ɍ�R0+�2�r�V�	e�=j4��5�Y�ݻ(+���:��~��u����뮺뮾�u׎���0���xp6�Z�����PR����c"�ێ��RQ��X�YmS��������~�>>>>>8뮺���]x믳�^%Oq�:�hVʍ)mQJ�Uf[Xa��X�Z�F5����kKmT
2���W2b#�b���6Z�,1X,X�(f8dƸ�Sי�V6�r�E�+Q`�K����2���J�
�"�1����U-� ��eL�Q�T�cW԰4j�X����,�c_\q��b-�TX=P�oV&SrS�X(����3aG��U30�Te�{����(���l6т�l[j�JQ�򕘗�����ׯ.�~ݼ��5�L�ݦ��$�e�l��,����rLj�G2��p	nuF�FJ�4�]*Eh!f4F���TSb�ˌ�ׇV�͠�50�w�7�7��|��H��Jg!�aX� �`f��BZ2�X%ucB�ԸC<����9Q�[F1����\�F��!.r�f.!Y�բbg+q[��.�W=��)雙�#:QuR�e�.f"0ݦ��\��6�	���3Pvi�h�](l�i�X:k�8�.��V�f��ڷ![���r��v��Xh�����+��Z�P�B:�K�� AU��rSlm��WQ�tqmH4��S�#������mL�4�Kc,K-�]k��4��ɦ��� X�eI����QrX�h![t��9���YR�����u�\2�[i��^]��ghV�ƅ��Sc[b�K��	F��m*&�ұ��^)Lmw��*$&U�feW6�ksz���	�/u��^Kiu��Κ8L�b��t5���[,�2��� Q�c� ia��������s3ph�nH�G
��4��h�ՕҗL7Z]�m�ީ"Tm	{�@]B�5�YhCݫ
kj��]-3�N��f�����%(Z(�Ѫ�k[nkR�WM����MvcK`-��kY���TӶ�ҭf@�&�m��1�SMsc4qK5 ӛ�����y��Y@�E�`�.v�fps`A���ˉ�]�,%cT�[��.Z�0�����CBgkB�k�t0��-�[�܀&n��c�*4�P΃n"�R��=}=�h�s�jk
������b�Ti��g�͗ ����y|I�K���6��ܮUU=l��D�[[uAf|�o��t��������=R��z��^�	�&L��D��T!3��y�֙puCMG'V鮺��qE�5�\a�Eq#�j�:X�^a���[����*m���]�u�I�
�jKH�Ԏ�%%Ý���qn��J��6�9�BMm�r&�H�L�͏lslk��r\᪉�kbًrm+�`B�T4
ۡlb���l�m����5,H�g`�V���� g�pEE���R`���i�Kq�1�ɕ�������� ��;���H���w��E�${z&>^���Y4��{:Ƕ�d�AL�>����7K�:Px�vƯ��*/N��|{�� �H^�� �,;��$��f�v��n��)}�P�Rl	m\I��@ ��]�z6Z9��$��C"]�����=�x'��8����?�;�?h��	�6s��BH,3��X�[�9ꓯ�{���ia@ǧ��Z8��r�ú�����$��Ĉu����o @-~���<ȿ@�L�;z$o����������j��k[̩�K�sE�ݡ5� �S=��5�Dٲ�Ŕ�,Vju:��~}��&�N�����/����n�v�H ^V<�&��v�O1@�̀����r���Iڮ�w ��8}Y����ݸ��(]q��%�z��y�>�s�� V+��x���i�͵y��.*�ۏS��'e8�#N�Ӿ{��%d�����u�^�W�^�A�ׯTJT.����!�ِ%�4��Coo�D�ֲ�e&�L�E���;��B
}���*)��vı �'c��9�[�����G� G�"[�zd�-���U>��ta����@o^�tvϥ�B`�d4���D^������ޡ�R�Nzǹ���F��@=LK�X5ܧ
�cf���I.��l Uf	�g�%�\�Sk)L�Cw6f���ޥo�Nt	dX�a�dã�$Ř�SA��-h����Q���n�}�>O�9O��H��~ir]��t
$�_o��g�I|��X��J�B%�� w�&@9{=n�;�P"��b@�Jf��p�_/C"	 &^��I����]��{Gk��%��P*���Z�!�E�4u<�$�A,��V�L�g8�۷��I@�6���?Ǉ�#�N
U��`٥/D����{�s_����r��q�So�%�T�r�M��,�AQ0��dg���z����z�Y�ת E��c�?g}�B~�����78����H<A���o6��tQ�s��$�U�$�D{z��u����Tz �w>���X+݋�����1��-�P�;�dK�o�'a�+��I�͙$1 ��29ˌK/;Ǽ]�B��D��5�h�j����H��1v*��us��]Yl$�ܴ,t�g�p����Xb�$H�!l�5��/O�O��]����H	c�g��'�}cL9O��P=Щ�jjmR�s�q�~m��%�#/&E�A��y�� /Ē��s�uNz4��W���g�a�:��\;�� & l���i��\�0�)������Ov�R >��,Z�q�%�����GY�'Q�.����.��ia�����d��(�~0H%����
õ��ks�=��6h�9���hb�)�tI?5���xC��F{c̕��K�����3�w��z�0t��s�ܿ��^�z�{$����;;;0a���E�_�2C��W;�`�d]��v�M*�2���G�J��b��ze�'���4�"�foN�%��Qww{���aV�k4���m�:Sfz��7v�(�pGB�9
m�	La���ߗ�l4�������d��]�2,�z"X�i\�;�N�㵓$;,���J�	�5j+]�P�#0cv{(
�H�ܬ�U��ޒݏ���xh�$���2@�Z�QF\�S�]����ִq�)�;�1�V`���Zu���ۭR��ށ`�Z�@�;7�E2C�U篜�0
O����X�����^�,m�E�wfI$���Ko���<���8� -z0^�N���N� S�d� �29�#ݒ^ߌ���;$��&�e���0����������$}{�{�W/z�^��}	^p�s�sw�۹X#�J51��R����s7N=:XVH�����������}�ͦ�jq�,���/���T���pg����r>V��*z���B�պ�1O2�'���뿻N�z���׏^�ׯ^���^�WÆs���ݢ���X�n,� �fu;6�+�R�V6��Q��F�@u�4��d7��K�P-i��ح(Mb@�vt\�6亳P��Z`v��D�ʚ�%��6�I�P;`�K��o3V<��"�2�Q�#�%�^mq.��f���Jp4[6���!]��;:��&���-�8��-�hb]&��d�5L��$]��\��[?�~��$�l�?���d�i�N�lI$	}��7.tue"-�Qβ��t�%��kU�OB&x�]�Nl�y�lnS��L-���@��:���@��\���,W$��\�;��d nc���#�hǳ$HZ���3�{�o7_D K��g���I�)�;���/K>H��ލT������ ���,� ����K�ٙ���D�q{*�˃���l,�M̖�r�)�tѧC0�& {��2	$��M2	 �?�3��k<{�5�>��h�uh��GM�r��Hm�8ݩ1��\��es�nm�!�ￒ�;%��o�cױ�-☁,�FncN���b����7�A�(�̰��bA35��D(p�����|�ro!�n�}s���=���p#��\�{n��.k����S��_G-��Ӂ�ݡ���=[�j�s�X&�'�x��
�|N�� �����z���z���:���W�<�=�ώ�D#�4�vA	j��� ���O]ˮ�#�Mg,P�0���ɐ	8˵iң�����Iw�`KH���Hc��`F��X$�R:5��(gvޟt��g��rLLT�������k�{�_��4deF�m瘞���<r�1<P����ꌄ�nH��e�14���TQ ��{ k$�0�*˷qBu=,���j1��52(��3)�͜�XE��${`��6t
er�������h30�@�pY]�� r��%� ���C�g%>� K�ߚ�+!��4zt$��	'���d�&B��5J���H�	d����$@!��t� �>�w�|�z;1z��&��>�B!C��5La�_d#̑Y�8�7�GYBO�sg�K��z�pFC	لp��[�v{�WM�G�F9��Ț�0��c�����r�Έ
E�
��k��g�$2dɂu�רu�ר�??3����������H��pNAxB0#�_��7���=,P v)�1�?��C���\�ǳ`�/`� ��d����w.���z���T@&�(���=�=����/&�/��H����B��bT0�u6�3��z�f�ԃbF�-��6��;\.	���0q6�Z)[��0�-�R����A��-�Lc�"v:@��g����6vt��_>�,�푒H7��r�C��k�{5�7�a����#���̝��$��bAȭ�Z����ts%��ޙ̼���`ts� �s���Q �H�����%�������E�k�$-�e�lQ�ؐI �oD�Q��C�}v��\x߶�O��`������ANj�stS��������{:N �[��xF��L���+p�>�����9�u?�?jD)�8?�5Vk�~YOB��Qp	ǌ�d����Ks;3���D�ׯP:���S�??>��G�g��:�wĿ4B�&n�qY�T1@��b�*�quW�K=� H6�1���m����Lln���p�xI���
�:��[tK�/-��2��Z��Z��x�7@={=�wr���˙ |�/�D�e��L��G�
geM�y�H�Q�؇Gze�; }�"S,`#=� ��Rw6[�cE��%�g�ǅ�\�Y[���@%���$�s��(M{�_��A��j��12º}�\B��G��@��ZK��d�{�AB~��삖I��MB��!��Bg��S�E�^)�� TxM�G�1��y��K7��%�d	"�/2{��S9�� Axpa̋�z�B%�gl	�0�+�g��X�d�i�-g	����t��2���VG����(��b�7˯Q���J���^�C�A�l��.��=�;�[�#�	�C�7���F���ǯ9��x��q�K�1�aM87��K�Q�)��#6�\B�#�ۥ�������Kx�Ǟy���<��3��{�h��0�m
�M.F��ˢ�Z�f���[2b ���x�4�fĦ����6�0Y�# k�JP��hCGܑ�V��밈VSj�F���L��Ks���5�!GLR�B]�-Ү�:��cq�(i��h�+�8l6
�����i�D�&�Yh3�f�e�LۦI.V�iJ�%��ں[��t��u�4��1m 6Bt!("���_���}���v��c��KK-�Ȇ z����1�Ų�QM �6v@�d�ѕ��N��u�U�;ѓ �س&w{M����usR�H�6:A�(WGL���8@*�����Kkc=�$GB(�;��(����Q�Ϡ�G�go�&H,����^|����H�(���L������!�;���Ӷ�2���\��Se5�G��ء�5,c�wv�� K����va�q�X�'�p 7:�{�
�oYj��1�1�s/�M*ب�Ký��d��S �7�1�^W����p
H��$�Tԕ�m4Ħ ��S��"f�%��8�qec1�� �����xgsÚ�x=��iDc�:%���3�/�,:�ŨqS�v5��C%�K���w��u�8��5�
jlt�i,���J����:��]~V�m�����.��	����AΞ\tr��9�mt=<8xB��C}⒛
yQ~~<~=N�z��ׯC�^�T����11v���쟑$�p	!��{����#�~��Ul0�N躆B*��W��L��u�Z'̓d�9�~��,�`����H�%���I
(�R��sD(Q	'G0�kM��}0Ph����H�M�\M�D�I����q4^��G�Dn+��t��ͯ,wQ���n�e��� �\)��}��1E���$��,q�%��ϗ���7�?/��? 6�ڃ-���3V�.�Tr=�1�ͭ��4�Ԇ�i2e~���K�c�¿d}���˙��3 	b[}�!�,���6�M�z⡊$?gCK�H5��\��a���[�$	�uuxg#:��Ib��@�N�>1@��"�KQ�U�D�j��4p�����i>d��C��A���X�%m�w��N ��<�ǽb�R����r�+�=�"��°��]��uÝ��u z��V�<E5xax��dW[>���P��"�!��E}�%�L{&�{wF���3v>J��(����=�5Q_nĖ��Oo�m��<�n"+cާ���+H��d=���nnC�3�=ɞ'���t.�ŷݹv�6����ٻ�%����3��y�h�x�i��
ٝ>@��v�� <gv�{���O���C}��;Ѝr`�O�c^U@3k�&�UY�(kwX�?=�q
�{�/R�ޝ��8�^�-�=���dq�ti�%Ӿ��Jwp�Z3e����L�x=�38=��z�tvC,�m6{|2�>�g�o#=i�X7;��G��Z=�Y�;|�4?�S���/v�oz(�|z��b0�=e�T��9���������~�+�,�Wf��xw��������޽Ïg�k�����q���~�U�4D\�z��i�}���q����C,Oh�9�٩�{`J�d����X�w�����
��g!Z���}��0��r�=�����4x�}<����w[N5��?�l��Q��Zk-��=��,�=���{�b��O{�]�p��U�;�Ȳ����qo��"^�?��q��_{�.��;�ձ�˫�^ws8���<zc�ѽ^����1�G�/r��=��v��}���D������D�q�ވ^t)�I�1��$� ޸�XX�������ۯQ�3�	"�%'0�q�d�$��^�] ��ܺ�]?�z���%5�~��z�R�A �b���F����T�-iV��QWZ�U�>�ϧS���}>�O��f�뮾�u׎���=G=�s�9S
�e��F���Me��ў�8�ĔlYgs���y<�O�����u�]}:�u�ӄMR��DV6�}�nm��
��4ӫ�-�0b���'Y(�e�G_���_��_|||q�]u�Ӯ��2{=��=r���DX��jcy:�
�}�LZ��ܡF܊��/q�}:����]|u�����]u�Ӯ���]}f��DP���Ŭf��eA�Kl�" ��TJ�S))��� �e��h�cYիu�>�1���)�'�EV׶�Sm���U#�n�m�e����*�̖*-/.'����Ե���5.�֊v�J(%kZ��z�`!�Lw,�QDX�ƭ���V*�-�E�X�*"�weMUb�FL�l<L�.�JZ�5,�X�jTDEE�����e����J�$����*�/��}=�z�:����ׯE�=��� 	~��;���ދN]ʀ��s�GGK��k��S1W��X�$�wa-���t��A.�Z]k[/ؚfYN>sA�0aF�[(���ĉΌ�c!���a7Űk+̟L�X����,H��3��v A�n�8�r"T B�PA&�\|v�Zz��l�\Xи��&��lT�	�3I��t�K����_���ίޟ`~y��i���F�@u�":.fA��e�R�ޖ�����C9$��{���@*.�z�Xc�̊~ގ�A`�2e��� Y���D�72��Y[����o����>���Ü�|C�dftHL�-��{��|�I����X�� y Ovt� �7d���Ç�G���\�|n*�Ƙ�k�Rnr�[���J��m�Q:/��{���/%�����ƴb����'N%%>7�<ob����l����5<�C��k|��-����f ̙,��ɓ&"#�����w���ۅܨX>�}2I �� uADy��^�I��&�$����+և�V�������(v����\2�g�2��v���H[j��W�ʠiu.�9��%>���;xB�29�ָ�yS�Ɋb@%��$cC;ؒ}�K�\b��޾�.��R��@xu1���ϐ4�|�Q����ǰH R΅�������֭[UF�{�}R��Ѿ�S�Q ��*j�dHzy��o�9��v��O
0ɑ���X�X�%9�2]�f�;�r���>�9�zη��d�wt�&X�̹�K%������!�'=� ���%m�8�4���i �c�����l����}�cL�3�������Ԣ6"�v���`Qd����������V���W+��x��+nũg{��X��i�E+�'������Ug���B]����
l[�d�b�C!Y�d3Rh<ЄԷ�)8wt����7"�S-'7s�/����zz��^�{ׯ^���_(���ߎC�)i����iǝ��+7h��h�(�T��F� l��l�I�LH�+h� �xu��,��+�����K-�Mj��`-&��lݦ�2��X�J޲�+�֎l̗�v��2�{*����F��fti1�TŃL�F�-������':�U���[
`&�7��J���63�20�Z���.�"˕tS7@m˧�����A���pc�-z��,���Ɨo"H���%��p���{��$��͙/u�С��IP����D5=�"�>r��2@�A2�s ����a�3�=�Ͻ�r�po1~��o�V'��P�������2
[��ɹ�xw�ژM�ȐX�ކ�a �g�O�YD����� D\.�bv��Z�#�B#+�tk�q� ��%u�P�d'ŉ���]�:P�Ù1@{��$��Z�X�^��bEC��kwp��Bi[�Ip�tA$�;���H]�GK��"\�r�������h���#��yˊ���7T\h	f,�]`���2��8q@�b��$�x�@�L��ޫjW���t���h^��:��E��Bg��Ȅ��lۢ� ��<�9�u�t������z$���{�Μ�m��̷��{)��~�o�;��Zw�kr������o���/����O�z��ׯ^�z�;;;;81�"l�@-��m.9���fA �an\l�g
���\���v4%C����6�?�F����SOC:{^�s=Y����V@�$�[��d�6I7������x�-�O_��|����}s��o���z�93���F�U�$�� ��0�^���W���A'�ez�=B�ݍ�R�Z��i��S�Q �-�SQ�̓�nt�������kpy��Fk&��:�h�A�3�s Nt^���%� P�
I�ܢ=.?��5<�F��^SKsR5Wf��E*�.�k6mJ���|9�ú��}��Q@';6d�Z�;�#�\'���� �^޸-RϐH>���p�!S������/?(�D�$�lKC$����X�1p	Nk��D[�7�gd!��7�0����@1�{n�	'̓PU}U$�����pZ�&fG���5G�gK�gM{����WDݫ������M�:���DD �S��c�rJ)�+���*Nڶ��N��􄊫�O��y��&L�2dɓ?�>Z2���XK)J��e%�ݭ	@��)��o�;~��wpQl�!gt4�v1~�iMZ�f��u3���eU�G��H�t�~L�x�/��o�O�_y`��c:����'���Y��A�t�[�� ,Ɇ@:���<��x"�3"�`���a��]i-Ԏ�8]*�-�]]^��l�-`�)�(t!�<��}�K��
�H�:��2HvJ͑'̐�@i�R�b�!���b��X�;�S�$�{Ü:�(@�2/��� t����&�Cl��(c&Bs4̲hgL��Z�2s*oÉ�/s�gC:QH��7�� �8�q���`%�5��p���<�G�4o>
�!c%]"l�Wv3ɆLz�����@1���=�5��큝�_	lcR��ȉd���Ngtp�i͞���!�g��a7�=<�B8����,ɠ�Ǥc�{�^��~kF��������ܽÔ�檮(] �ikdɓ&L�2d�},���_jD��I��ք�Au	XF��b ��}"��������:I0�$M��1�����$[�:d�ĿO����E��x&QY
]��Jc���:hC4-�&�bG4-��ٖ�cm�nW���{�B �B�aڲ��I�7��$?tI�q����4��	�sػbw����A'&�����C���f�|�� H�f�Ke�O�L��n����Q귃ёy� �=�8��9B9�}��&wve�����*g��w,�J�r�"�o�aK��H'��Y��;�G�����>��>
qdi�$�A�)���	cL����d���8���=*4�Y���N^ ��ƾ���H�ِ'yp�tVKb�*�A3��,@&2[�"go��u�.A�:%3���eAOޘ�����s���\�h�w#یf�5xw�q���f��]�؀��;*�S�]T�eM�˾oѣ��$��>�-�ǵ�Ɗ��e������;�8�8�ׯg�ן��׊#���3h�מP�1\�n��� ങ�5lv��:5m/kljMٚ�8�f%e�R[T�R�\r��fb�)��� X�QdHjF��tУ�+�jV�l���U��.n�m�H�4�ٵ���frM�0�ZR� [ʹR,u �fe�6k�+	v��"��w:�U�f�s�.VX�i��n�U���H�����0S�q�aey��,ʐ~��ͺ-vJF�9a��y�`�)�%�o���3�7�[�wU7��_+X���/d	%�//�z!�
.��9]�$�2�^���֤�z���9�/3���q�z�Z�s���K+��zW�Q9���.l�M'x���k�	�FwzD4����[,r�dOG��0	 ev@$�����C� C���]C�=�l�8>b�����N2Lg�5ULBgn�����S��d�<�W�ِe�=�I0TP��X.��)�!��b�s�-���toxdy�����2�tȖR�\dk��Uʍ�B��h�7mV+�\�՚S]�]a٘u�]0䚙��uGM�Pߞ�~�t��(�D{�dDWd�P$� ;o<�c��.&u����5�"��H�t�3�q�˩eJ�);SE��@r���R�}q�+ʉ�k�zm��d� ]�_����F��l����{ۛ��2���op�n���q<I;|gܳ���,��,���Ƀ�dX �e���5q� ���M7��z�:I���~�A����#.�H���t ���pWn����Ml�$���- �3_�G�6l��0a�Ӽx�t���xSۛ�2@�ײ[������$�{�ӽ��[~��#S�6|Ӗ+%P�|'W��o�a�BM��˽\�6Q�GD�HF�� C��2��9���ގI��Ĩq�z�jV6,�4i6�ƻ�F�se�f�d��!��[F����DC�K���$�P��<��?�E1a���y�ޙ%6��7+�����+ީ�8���i$��>�!9x�Dz�g�\H.��j�z��lG��H�~0@�&G��L�N4b�ͩ�eu̖��Z*�Zp�R,�ҲZ;&UW�.�D1�������r���_v*j�,�P�o7˱���q;�W9.K������ww-Y��N<�S֐��iĂa܈O�%�Ye�Ye��/r�s?��<Y�� �s=!���b)��wFc��N4���Ĵ,�R,N������� �c���6$�0�=�C=G�i$�g��a໼f��dă�2n�k��3�:6o�1��$.}6��W�fda�vt4�X�HS�}(A�t�%�	c-��7�Z̜��S)a."�ۈ�%����3�����D��P!�	�|$^v��y�bXN�cP��S��F�A�o<H:�T��LAJ�42w�X��I>�i�*���e��uV�g�� WWCI��N��~��Es�$y����@"=�~���fMn,�l���:e� ���'�y4k<�kBw/
sCaQh��@�׭���:ŖflK	��$;W��Ψ�?o��+�Tßc��Y�fc��}�n�?x����{�u�M���]9�}Fnibs���M�&�����^/5EC�6�dɓ &L�2���,�	��$��Ԓ �3r��(�b3�Fǲ�� oW�aO�z\����+����ia@���=����VR�ޟ8���}}�ξ;h�m)�m&��T5��(�2�T��`"�^"%�KW����w����l�, F{�O2E����e8g�b{Fa��Iid Ϸe��mOb��P](��dʹt�̙ �kkؼ6��[p�:"�2����%72pJ���%�V\�惪2%�'�g�b܎���P+��HY#ذ� �$���y�)�^��I ��ai�b���~2L_��	���[&|��ǮQ�����<ŀ�mgsL������i	2qލ뼍�4�]�o�s/9�Н:�A�(��������u�$Y��dɯL��{0Kjd���@�DgX�w�u��Ĺ��"U����P�z�jqߙ*?��y������k;���=�<��3؟��E.���Fwru�1��������|�h�q����;���I_�{����.{|O�a��
��cy�*����(	[�e��U�����]����rew'�ܣ=��i�x:�{F�c�9��{�WQ��X�+\1gB|4��m�vk�{�V�7G`F'F������+�{�ygH7M�8�r�)���\�ް�w&q`�	o�����O������5��wr��Vq@/�^;��z`D��p<��5�6?r�/�:�U��!N���3MJ�&|�;��Η�zMs"<V�+=�#�x���Bx��־;3Q���/m���>�})^rK�`=[��.�'�n���W�)Q_D�Պ�+y�� �����(��zxs�-��Y\�S�zuqmۛ9�:w|d��mo����5�Ur�또���d��c#�Ǻ�o���.��گ,9��N�o��{�n��S�������%�UB$s�+��؞���W���oֶ1�g��������=�������|_?+���.r�m�z�+���dz����Q�������(�z�:��Î"��
,��;�p��ӹ�2�KZ��	�)���aEdE��x��h�O����o`���_v��)"����(�/��1����A`���l,(��'�M{=�}�XD圜h��J?>a4L��Gn�f�2�`^1��{�P�_�D��ǮT����L9R��0X��n�ˡ���B�^O)ɼ�:��%���T�LI�j#|��0g���̟.4%qԡa&�v�p1�8YI\ ��nϡ�b��7�ͲeFxu�V�y��S頠쭁��x��II�X^),=x���G��̢�	��X�V�����Qb��b����TUz�w�r�~?���믎�>>>>�u�\u�]z믠�����#�1T��ҕQ.gd&�:�Eq(��+{z+���b�S�����_O���������]u�u�\��g!���ت�R�"��Ym���(�U�SS5���"+�A��QK<�O�s���}>�>>>>�u�\u�]z믧�TDq��-���m�{�T�6PEv�M�C[;krw;�O'�����>>>>�u�\u�]z믠�
�+V����N
��UQb3�Q��t�vʊ"�V�PUf*�6�EC���S\gv�cb�Q'An``�G��Vmj��.am�TF
cQEB�F VT:eb0t�䭴b�h�e\�F��L�Db��d��Y��!AM�2>��ġ�X[�`(�I�,`"�J�ǖ���`�T׬��q��F�(�eDAU�Zň�Ơ(��J�"��T�$�ES�Rz��x��)���y�j�!.�A`]�P]q�x�a1M6��KN�l�hQ,00�&�H�kY�l�SXJ6j�鈃e�q�ZGLe��J�2��u��b�0c=��Z#��˶�-��;f�(��+m9YFR�Vͻ%^K�`�n�Kc����m,���׉j�J�xZ�a	� 5X�,
h�a
[pU�j�΂�,&K7�/��9��	�k�c8�����*��8.%�wc4�!��^74mj�&Sh5�iV6k%�	�����IQת��Z���d2�j����ƶn&є��3�eRkA���n�\�Y���Dن���X�˓�*��,K��5C&m+y����::��3�j��ni3v,S+��UءpKiF�C��ƪ4n�R�n%�J],m�
MX3qH��f�%#)\:d[�͉WJkv�du7\����/7eTz�ɵDpi�wh�,Z6����jF�͢$�ҕ�e|�q
����h��6�S�[eʕ�M�XDmK����ce�Y�Wfr�G U�iG,`nt�@�xh�	��ږ�-�X�,�����&b���m^
�o`RY��U�"K����)��G�mM�:������`aFc1B���h�u���6��
-��������#�����}]e��u���4 ����fM��jY\#i�F6�����Yy^s���M+��Xk�;e�!�����3
�V�j% ���9�l��:;a;:�e�&�t������h���tCL�Е����b��٤Ζ�Z�[�Ѽm{S7�b��o'��-���\�j�;4�&��W+�ULM,l�}^rhSO&y����I�<y�KԘa��8�8�8�G>��HS3m[GZ����4�3gq)v*ڄ]�r$����,�p�!l�l�(�6K-Z�JU,u%���������ez�.�n��l#�[��*��b\��-�Ya&s���&uE1jL��٤Tˍ���J���c�-����z\4h�+6	��wTQ��rҷ5v6hm)�TGf��su��4"�,�I�H\������z�pK���x�o�@��-��,�$��H�6��LN�Du���J�
@I�hoz�M2֎��.��P�蛆H��� �Iw=�2��R��yZ{�������^s���P!̏0��� X�w��U��vW��M�v�D�Ś4�E�����GD�D�A�9� :�>�+��b#�kv��%�a+�36��I_uGt�t{A�Jk�!�	�$R��u�;���
{��${�=�󽙆��ώ�@=���-,�&Q��ӗ~�8-����;|��H~b����8y]۲M]pW[4�a�s�Z��]�[X%�8������ȗmM���?�;��\�F翷�p�Z���z �dl��՘'p�q ���ĒϠ���|xx`�����U�^	Ug>�O�W��3��TM^՛Y����si#��||W���c��4tD��II�yr��B�Y��$sKc dߎ��ɓ&�|���A��ٓ�Y��iv*YV��l�����=X�<A�	�(y��e��>�H�d�O���#к��2Ds�O�� *::d�v	�	�D�9�j��j��uD� 2a�c:%��c��<�S�j���l�A��d���;�r��oC�cC�۠��<;c[��LUe����[��F���*�Ƥ� �~��|������86.!�3*�Mq[.��M*�Qq���61��%V������l����>��	W�-$��qlz�z�2v���:*.�S$I^͐%淄��D@�]�q'�� ��bD�i�$Og�I`�H����U���'{u����S?z��<��"�s!r��P$�x4ν��,�OL��F�C����f��y����;�u	�]^�����&��Ψ�O!gX��^�hTNI.�u�f�c���~q4��vL�22dɓ ���n�]��So8�d���`N��O�<:�����6;b0H;�r$�)gCmd8s�Z�czO	��gD߽�`'lo��sk�{�	2�ɜ��]w{)�$v%��A$�_(M!��-!C�����8��D���x�:�2���u�z�n�3��Ĵf��3���l�}���o�@w�;�WVCI ��y"GotH�qk[��	�/��gc�|Ĵ3��c ��JC���O0w�α�$*#���9r�ޝb� �lA ��6��I�x+Dz���4Wf)�Ј5x����z�"X�����/}��V72[�2@��%�	}F����"űȻ���*�{{�`,�Ee< K ҼΎ���`Bdsx���mn�y�������P7�'�ʊ��k4�����k��Ӟ��Vx��	H�׼�w{��H�ֵ��[��s������/��Ie�Ye��-���<߹�s.��x���\�&X�-����]j��#�D�H�"՗wfK�dK�t��ყʬY	�;t����/
eC��L��i�mt+bMf	V�Gl�sjU^޿}ϟpT�uj���}ˡ
d���$@,�'���؏8]H��z�H� �t���l>"!@w�4OGm86w>�S  	 �ó&A$���,	��=�O��\yg/��O+���)��)�gl�6�5�w�w�]���A$���i>d����j���0�tD@�$U�z��Fk�F�7�s�g�-�����ʖ�q��7�y��d�O��C�$��ר�/
�_1ó���֋̬�g��z�*gQ�� �
��I�ܣ����L��.��~^޹��:���ܺ��C�O
y�'��&���X����;�\���(�KB��AS�A@a����\�'p7��S8�!� dl�B>Ϫ]��u>�ɼ����y�e��=m��~ya�Ul��w�8�8�8����)a~�},�;e�]�F��sn��B E!������״�v�9L��Ѡ�e�m�LX1K\K�	Q�d�����4�b&C=�]�-�2J�!]+,�ƌ)� p��I�4�ęƃ[�*��H�5^y��b0BhR�K�:gZ�ⱖ�b:SU5�!Er��/[B�mc(b�c2GFҐ�6�m�9�*;�2�U	�B�O}�o�"��D�k;�$�Um̔�d�С���wp��U�2H)��#:�*A����a��Pi���������4�4	.�GM�;@uɄs%�������n�1����r�͕��Y4�4 �㚠�	�I��G(���K��5�<o�0&�֗�PS��u?E��/���d��ԉ���@,f�O?x�wF��d��0
��.�tD@�$xS��2]��{�����$��u�KC� �Ѕ��� ���g�Y�,��	Q��_��E�s)k�A�k�e�%e&�ȴ�ً�Z�kr����~�k2�������=���$�tIvz�57��e��;�N�L1�.�搥���n	�������Ya�8���F�>B��*k��2*��	w�Kק���Y�t���i�S�&T"-�*{W*�{v0�W烲���:�/)L�D8�ɹ� �U0���ԡe�,��,�����9����-ݽ1N�������3�oD�7�U���N��A��,H=��$�Ƥ��Nc���5�0�y�yݽ2�l���0�I�ԯ�ȏ���Q���!����x0do���	�O��+F^�z]�Q �_Π��$�9�_�BO����-g@Lv�왒]z��a;Z��;���P	c�Ά}���Ո�KZ����_�5�F)8�"�1��՘ѵ�:ŕ�j[���h~}����n�V��z+�Ӭ�#�vpo��@'[��Ҙԋ��@9��y4W=��"[�o�)�C�?�߽�o�it}>z۳NI�J��d�隄��
�=B���X�eH��^ �O"�œ�c �d�e�A4�	�CઋBb��'�œ�y8�/7�Ƿ���~U���wMz9� ����b6�٠{��xu��{ ���t�'����u>�K,��,���>z����ْ/��H��j�PD'P���!��37Q  kk'�*陖 ��^����Do#1� ����|P�9w�2=L@}���T����!ۘ�L�zT�B2�1-�32ƚYܕ��,���](���)s�]�r|"�0�#1��VY��an�(.8�a�8�[�ݣ/�~���7����Pݷ��@$E���s8�Τ2�� ^��Կ\� �Α${��ݼ�$興H��03pΘ���f�N��cѤ�%�';��� P�:`Ӊ4ؠ"L��ڬ2��q�	��)%'�e y����LjZ!i�	�B�Cz34Қe�����@�k'�Z��54���Q�n������)4i�`�
!D1
����uȬ��w����d�h�Iӗa�O��U�Հ/\�y���	�Ao1Sk�)䛾O�; l2�n߿���:ם|a�vl2�WBH�C��ƦE.ވ]=�hHg��������~~j:E�{��vt9�t���{���T����LI�D�Q��yy��^�>Me2,'�`^ڛi�UFF0edb �H��
A1�Y�Xv���h�((�&$�&��ǥ�6rYe�Ye�YHd�d��Q�9��w�/N��>5� �� w�v<y����,Mt�dy�	��g~��o\�۹B����֒�QJ!"I%.PaQ�Έfg�v�J�(F�,]4�(B[�P�ʭ���㾨B�Þ`n7��N�ra�@��d��ϼ�P�57����朂%�=�Q�@�e��ec�
=ޛj��C��<t��9]v��?_��D�M1���N	�����y4b/� Āfj���%�73�YS�3�B���������6�	Їx{�l��˕Z8GCܝ�Bt�$���̂Ic���*��z�@-,�Q��GQ�Q;�O��\�$��"|j�/&+{*2��t-�m�@k['��� Sg�%�OEc�Y�K����w�w����
�t��Wp>������b~��{}��^G�����^;�ͱͭ��^ %�3�S���~�����
��'S��
��?9�Z���O ũ��d���:��8s�M:z�ܺ����K,���Ye���K~$+�5Ж���U����R�A�nҤ,ѡ��e�	[s)F�nV�Jb�-�m��h�k�B,��FR�4�ԩ�m�͋`xQ��T�Ga٬1(i�lK��ZZ@
 S8f�j�n�Y�)�R�p�-Xh��L$F��P�!]�VU[�h�V0�MS+�XQ�ٖd�9	*Y��RhkA�ìa�!X"Kk2�eM�5�46l��͟?}Ϸ�n�j��p��t�ݸ��'�K�=�L�3��y�=Q��1����K<�-��@���V��!:xFG���H�
ޚ�@�r.Or�D�� 	bI���SCU�}�f+�TV�B�pAP�D���z�ldA��vKI#�N��=JH ��W����%LfjtS�b!##� q��~�g9��%�כ��b��(��	�+Ok��T^���d�R<(�A��#CMvv�?v� p��-Hn�-��wL��ΐ�װ(�j}� �v��{����|o���A���ͮ ���bj�D��[4Kq(*��͆A�ɕ�|���)��w�<���9��Ω�I#�t=2kP4���2q�l��I�L��Ȗ��)`�b�;�b�o�J��޽:��f�H����*/��4΁��!�f�ˇ�S![��g�[��{�Ąk��G_QW�o�7sq��ޥ�7^���T̸�P*���,��̖Ye�Yaz��g?��xŶ���s�cqy]����	m�V��!:xFE�[���yL���vT=^d�Ge�Ib.����x���(�%k[��tg_�qF,I�H��bLO�y�(L�5g.���FO�9ݬ����t�L������BFǍB�d�WeEqї�n2��l�_NHI㖡آ	���1#���^����9H�cK�����nE�&G[f�ZC�Q��Ku�P�ۛt��ۨ������7sr$	4���,No\ɰ=��� �GH�9�-�T�<ޜ�F	x�P��ޮ��62��7'jk޾��	 �.� �{�2���k��G�P�=0M�9b�����Jh%�c��'!����;�Ӄ�����������JH��kd���a��A�>����o�G}����Fy��ބ��1/b��Y��t�5t�WSw�W�>8�e���W��۹�42���	=R�w_x��~ȧ�Ⳳ����i��F{���j��=�s�洫��/} �Ažw�^v7��p�Û�.����J�gnگ}�۽�t�񫴮�ya�q��&[����F��6�ա�w��ygi>Hv��v"�|3^�<�-��&{x���z{<�NŚ����y}]=+�WY�>'W�f���;�H�Ա�}�0g�Pq�<5�_I����Q��~Q��oۡl��C��+�t�����?{�+LZ{���_Dw��WK�w�Ƕ!�����k�i�r�g]�ٯ�Z�BI�zc]�o�\J?��������}��/��^ [�.y�p�Wy��]�n�3�VN�Ӑ��0\�؆��=�B�(9�*��ʴs�ٶ1��t�����g���xYS�g"����{�6eY���3I��h�cO^�V��Ǆ^~����Uq.�X��,4��?[������sr������{����Z���*����w��	�黺c>TJ�P����U�e��X�ڰ��C3�Ч�q�|8q9h.X���2�\���LI�i��E����()��W�!�N���'l	�I�q;HV�O�b�Z� PW�r��M� ��d0�q�C<�^��32�Xv�嘆�1�֯��+��N��y�F���ݿw�\}μ��{���*ENѴUQAb=5����1�.%�,�*�EZ�X+��g�������㯏�����]u뮺�������gv��P�k��Q�H��q��(�e񺓎D��';�# �\~�_o��>>:������u�^�뮺㯤�Q��;�v�*<��fR�jeU�����m���s���}>�Og�����ۮ���]u�}>�<�y�L'�멩[F�eUbZ�)b��)ӦҺ���4,�u>��||u������㮼u�]u�_Aއ�0���UeܦJ$��Kj�P�V%U�(1���E�Y�j/�UG)ET��-j*���ƽP�DR>ڮ�4�YO-EcQU�V�3*V^��ň�U�a�n��3���]k%N�udQU`�ŕ�j��Y���:f��"�V*�XW��X�N�6�!P��3lQ����X��Ŭ�)Ё�e�*x��d��&L�Yb�3���4�"��W��s��M�D�%9�ŏ����gt����P^��f� �0ʷz�i";�oV�r��r�P)�o�*��P���H�ˑ3>�Ǿ�5�l���A:���碈�Z�Ȁ�s80�+0vH|�JI�%���m�X��͗jY��k,z����
Y�]v3*Q������Ͽ>]K�+i��b��T9�@#����H�������yA�@)g�٣��wȂ�Aw�����7��,F6r��mn��!2�p3��y��(�Nֺ����B/
ŭ�޺�wb��D�&D��z\�E%~�@y�m�T�	 =wH����	ȇu打ݠ��Y��n2
�j�B&�����lc�r���Lgq�������?�����{m�7�o��>������('|i;�K�~�{�/ɣ�qÚ�N�p̍/��rYe�K,�e��~cՓ,	3����xN"�9�aG�$��v��ɧ�~3�L��xĀ�}"I ϻ��Ki�Rn�W^OW��ҡ˧F%u���HdvD\�J�ă��ʦp˜ԕc�9��9z�!�_i�BQJß} ��;�I��ysg�b#Eܚ�Gz(k �{�d��I��9:)���kR�QR%�Y�3�b�,;���}n�H�H�f�M �w�d��ǯ�9Y���OG;���C=Ȅ�AOa1�cI�x���L�ZJh�g�v�H3��i�{W%�0C������t��>��y�c�WH�	�>"��*^W,�K���cGY;�	ȇu��3�x�X�j��<�����m��A����T���������r���?�ɥ��ۃ�w�{7%����G��u�)�r?��3���O�n��Nً���0rG^|��/��m���'��R����6�"ɺ�ݷ2��]��z��̙2dɓ	�E�ޞ�ݱwv����6
�6fѰ�����&%k��t�[*KVjG��.���G����CjB�-�,�UV�1�f&��nل���"���.�3�\3=U�f)�3lb�Z�u6�#hl��锖iLt�ȗr��X��Z�	�īLM�(k�֋���Y��T���F���˜�l�4�~o֞z��i���٪T.
�(CcV��NFmM� GQ�N�ϔAq��-��{$I�Kʛ�"��f�[2���P+d�cpǼ�L�uĲ$=ӑ�&ڽ�tAP�D��uE�啞���y���H�l��C"d@#;�%�2��\�Fwo�7r=��G5V�'I:""
���XW},��:�y�w����X�{����2@2�=���AO��2=7^'���ƻcQ��f�=y1�A; !]�+z�<N�k��� ��)���DC�<>eo�d	jeq���d���=*pDCxc)�!/u��˙ѭ銩v8t�K���c-W�7��>Vj�gC�`.{E�Ë�mM�0�e�������AND(P�	�w�X�ٻ9��!Q�3~$��>3�#H�.� ��͉%W���AB;��&O;�$��
{늅�j51}���@ص�s�ad�4�9��U�0q_��91�ux�{�WKپ��� ��1�VyjǤ��E?g�v�����{��/�? ��zt:��g�^���z��0#��q,	�}�'�P5��2	ˠO�C�����%DA(H���%���T�_��x����É�fs̴�3�<�GL�ib�3���wHDAB�����dm�<;ćm�6ҷ=Q� #��hX`�aaNqr5�}�8zɂ�ȓ��(� ��t���D�L��B�0S�X�>ɹi���3Y�ѽ)�YlG�u2m����w�t4wL�;�����:§���жhK3�G�e�U�:���Ȍt��w5�����ϑ��˛���~�fȖ2�N���7GF1���3��)��2e�L��vq��X>�'�0��(P�s��xN�@J^����`m���A;�2H�Y�O>�����FDo1"��ix�AB;��lb{ cZ�Jd�Q��'��N��8^�����>;�Bʝ����g��;a?V}�s�$��P����PX�t��j�U��Oa��V~��('���؞�z'C�^�ׯ^��eN�Ē��2�H/�� ��$�U��8O�=�Rݘ�x����G��"q���c�z"�����#��SL�jt���(W�2�K�o7����ў��G������sy���҈5�� ��铵�{eA�N�r�a'I�7�*�v�R������c���бu���E��n�x�1�
x��6nD�}�$�w��u�Nn��}>��'�Q-� d7mNh��üCv��2q��֬Xn�כޖ�I���50=��$�V��狀�i�p���!B��Ek��6޲I��=�4H"��:)��&/͌�[%� �w���5g�3��(8�x�^;]�'���OD��� ���2g����\�����4@Ur��P��Mz�%3�棒aQ�I�^>����f��?���LSq�=OV(�� �X�<Z`q��ͰҲ��[�qׯ^��ׇI�ם����a_\���p�����_}��	#�"}{�كC�������L�
bs�D׸�=xu)��G���n͂�8"l��jf���.%ъY��1.�tF1�ƺ�^�=����i�\Y������IR
���I,HY�4m�o��k�� *g�� ��H3�s���X�-�WB��J~F�O�u�&Ad�;6D1�_}�H�b�ga����1��{�1��
xO��[r$	W�	�d��L���ͬ����jH/}�&@0m��R�Cx/���ѝ���M��d��"Y�^���$n�ϛW=Z�N76�s�d%��V�C���z �O^<�*�<����vN�2a�^�t	;�@�g���<������Ee��7�s�E�.i�E���q
����OL7x��$���`u
�}�-gv��<KޘMC����\p��^~b{4j�� ����g�lu�*�;=_c��������ć����<�[%�o}���g۶��JA�+!���K�� T�Gl���3�p,JČ0��0қfʴ�5(k�!Ĳ�T��#kn�a)!0�fי�Nƀ�`f�4+-����f6T��7a�����4IZ��uV\։.��YYi���*��+�:��GF�޹�*�����M2.�MjeQ�e�h.q�eR5
�4�l�4�"��ٰ�c�W63{T��4�\�~��>ƺ\������x��2��M@V�;4�W�*��x2+����lW�yBw�C�$]�x�y����ɼ�nY�s��н8�I=1���$g����Wy>�̫;e��6է�B0𠗈��ɸ�<�b�N6TM��׈�A?vN��o�u���$�N�pS�x����ʬ���/i�x���B��H'.k;Z�v5 �+MDˢ]���+l�g8��IЄb�kK��JH����h���j�奲�C/3��\�}�D{c���tHC9��cm<�5 �6�aMq�k�s��[fDɦ�е <13*�	����|����}�Ƙ� I�ǀKb���g��'s�t�r�~�֔�N���E���D(p�+Yz�rІ�޴n��b9��P.G���n������x����;�z#�Y�:�Uf%Q�S*j�/� ��Y���@Bvޫ���m��0�vp䳳���.3&K��a�y��1M����j����O���g�΄h+&i��=�K�M��$���E�{b.շ�C��)��q�j�H� ��w�h�������K�]f�o�&4GNc7O��u�����Y2%뺴�WD��,���{Z�<;�$�%?���m3���:�L �{ޛ��=N�$���hh��$��zf���rK���Q.�b!3c2��!4��iՖ��]�M�f��H�����S���g�� #��4��S$Ĉ�馨g��>Ѹ�4����{�&��6י�����:N&�~� ��b"�:D��Z��yuӐI�z�� �Ӎ0�>_v[��}��tmچ1��8OK+e��ˁ �E.�[. .������0��r�v-�}���ON5Q�[�/�=��rI@���sh۱��uҎ{�]ο��BY���%�Y��d��w�>�v)�"|ʚ��.�f�%BN	w��2Mx����A��t6@2���S�]�"IbF.�{L��#xU!�0[E��ɤ\ �H�7�'��^"叚���c'��n�����CD{�9�x��)��̱N�ǹIܟ`�5�;� �Eˢ�c�2���#ֹ�D�[�h��,��jԕ`�ɕ���n���<.�w2��Q��)���7)�Y��|B�k���$�����TI ״��t�B0 ]�=��{r��o��2"X��%�t�#��r�Pl�dЀw3�'e����f @�	��T����yA�%;<}�(�{u77���kw�$L��܋!�����p�=��s7b3e�tK]
���A�ڀ�]���1�j �p2�������5�#�9w�c��p���b�e�ܯ	�ѱ"4N��E{rt�zЯ>��ü�0�������)�3&L�`�ڑ+�d�i���	ܒ�	!�-J�`;�&)�˝�5���[22ds �d(<ɒ��Oz䨇�٧��MAVXw�C�:���vsNr���"e ��5�aakۛB�}}x�^#�� m��y����ӓ,����t�2�$�ёBN��n���j�b���;����C$�}��w��gR�[O�lx��sZ�ƦH�:�RH$4�t� �m�үD�~�ɍ��F�$�Uw�dr$fGbR,v�I)�*7���k0�vڙ$%|�K$	���]���"	0��*�\?�̟sb%L9cL��2F����cT�#r�%�g�zKøJZ鸆4��]�S쪵Z�޹5�,����K�:d�K�r�%�0B��o�{�&.��W�����˾F{�gK�{'^J��}%٥�A��xe�s���
�����K������5�7���7Y�O�K���|��Fk{ׇ%p���Ơ�7���I$�4���[D���-Ѯ]��Z���ADy�n�}�ϸ���@>���h�YO��|K����7�X�S=��j��Q�w���ڋ�~�H��{7��zn)���2k���7ح�홳=}����S��uv�����W������2z{���ت�=�^&��ay7�Q�c�}{�>�;���Z�֢:���o��Z�q37�������v	:��E�ӳ�]��z�����LٌN6.�R��#�8w!\ܧ�V�a�~�=����^;+��ɱ����M��n�<~-��IZqW�M7��y�1�&/�O�������=�NN�+����S���^�
"L:�}NRwb${�'�ˆ�a#E�W�O���?o)���*U�l���Dw�z<�����}��\Y]=�E�qq-H;�d��q�.��OL�j�7T��>��{��0w	�����B{�M~��;�����d�;L���Bjc��k�o���ܕ���E�r�u��	?S��췀���y(G���Y�*S�6�ՋU���sM,`�$�j��4���E�������E��������f��B�_wv,�X��`ıw\�#�J����;��/��D
$%Ed7���:�X����y87NOov�^�����)�1

��@��0�m�C�ޫ���V ����Кj����!㇂+�r� \�'��ژ,�UwN��Ȏ&��b�<L]Ř{3ki��x2�����o�¸�=GVd��]t
��Rz�o�X=�iu��ϒh<�$=u�k$#	��>�>�m%�釲&[ضn�4��6'�2z��8�-g�l�z8f���ܮv�s�*0�EAla[��'�g�(��DQe�v��������||||||~:��]u�\u�PK�9T�>R��+B���U����u��_||||||~:��]u�\}��'Yd�0:���a���+�QbմR*���j(-�NOn�>>>:�������u׎�뮸��b�E��UU���
DNs�L�SK\}��o�����_����]u�_O��Q��0R
",":�YQcDC֫LB��'�)�1=���M��R�æUb�
��",U"���9^�h���8ʀ���qܢ�r�֕'�G��T��#RwF�m�-feC����j(Ub���]Ir�'L8����D+Q�b%eCY1��R,U"Ȥ�YRt���"�d�+y�MdY��PM`�`�"
�,���}s�7,\�:�uǘ�5L	�q��Iv�9-%͖;�SYD�Xm���X�WbZ�-e���G7m*���M-���$�%Y�f�$v�����)\a���-�N��5e 6��u��08���ku�vJ�M)\Z��q�#�9��M�a5F�����ZC���sL3.K�ݬ� �r�!B�V�aeIqa��e@KXJc*Ձ��[��it�4U�ƚ���XJ��ionr�t0Z��
�8��HP���XŨk���˦���&�R`�l\U�.ZU\[Yn#t*QԵ3J�q��T��kP.p�]Qu
�S\E9!5�fc������41�% �,����@�U��lf���bZGW`c�4�vZܷ8v��ʰ�͖�l�]�Ǚ�;9�)��M6w%��^K��sAa�@��e���ke��jh$�챕����[Gh�)��)S75����m�(4�	�	i���L�3�Z�٘�0�����`UZ:�k��nh�� bZMvL�B ������&[hS]��M�u�	��ژe��T�c%t��۴�����-c�U7��˦iH;M��e�`���v$:��D�x�ڐvM���5k��k��a�LN��u��\R�� �M�7e�M	�E�sq^rM�K�X��	����gaġ2n�,c��e�#�R=V��"%B��ca	s�z��ݔڙb�7d�ru�͚��%�4J�����ƙ4u�#-֤�$�Ù�
)�5�#5��K�����%����VvfT�c�2�;�+`�-����%ж�TaUլE-ѱs5��ܮUU�cs��ǃ�q�L��!��ϛ���>h�����.��w9,���2d�,��=���n�V��Ghp�.���Z��öM��
�f�hs�ņS]/����B��a4�h`̰�Z�-&��FMR��LFܺmR�l`�h�.����A�Ud�a2F h�ƢX<�ʝA��	(;��-��9v��c����n��	���k(�n37h.q��m��V0���Gh���[n)��j�3K�9��2��VT�������@�������7Io�$-�$>wL��ͫ�Oj�r����O���gAE<(#�MĻ#�&��曢�F2G:�5K�z�)_��>�($s?N�p]�(*��ۑ""��2A,�_����vv�&k.$c ,_�fN� ϳ��0� Zke'�&�H���w�Q)�%���Zܒ\;[c�%>���M�d����jII+�́"	0��[�$9��y�sݹ�G2vq;=��%�w͙����y@6�SpXҊ$��
tA���`e�4��0�ڕ,��B��-v��;\u�*���=���C�;̧�<KCK;��2�I-��ݛ�ͭ
�hQ@�����i+aR���I�!D�kj�t�Mqʧ;���]�/tg����i��]m'0?d��~Jv�p�3�^.a>>�дy4r�����ϭ=$E;�A�]6���K,c?�	X�w�7�}��"C[W�($�x���~˲���Իa ���/&�r/��y�lnZ���Z��ǎv� ��l�:�[�p�	�wK��AP=�Ez�s�"�(��a4H�V�T@��I�h�~�ꮜ 
mĜ�͖��jI>~4.9�d�ÐX]�D���=�J���t�Y�SצJimh�d���R;�ɒ�OX�/��5䫘7a#�즬���ke��.�3USme����зF��]�q��~��b��{���j�b����&{�d̋�5���fz�A�Hb�P
h��.��P���xK�L�$s��]`�>'ܽ�nS��$�W����L�Oi�3~��	���I�!<�ֲZ���5�q$� ����"�w�t�e�G�2����`���J�8^`��h�d�����/�As�o[�{X/>��V��\��|�B�dQ�o�z�ߦ��,��-�5�93�����:������Yo�"SNR̈́��P#��}�e.��ׄ�(mUt�Xy�"ƽ���G���6�ڢ�oX��ؠ[$�=W�໨P�{��%�� �Dd��ovZ�x<Hl�u��ycl�sn�MHU��Oz~~���i�?r��a��
����|:�q�-���]k�fpf]�u6L�>~}?��!Ȅ^	�6ԟ>!����he$��-2{;Ǉ������5R�P�dȷ�2J���K�A�V���hmTn���.I ��Ēm�󺀖��#!Ƭ����/����j{p��H��=�[ �2�ݦ�	.�h�� Y�%yқ'7�H�@'��UX(^��wrO	!�Ǐ�X��z�yy�F�^"�T4�d���M�E�o%$t�8����w�^�O�Rp�����������{ �4=�^�n����{����t~B���V"������:S������ �e�����T��O���xl��JAD(��b��2C�}��{<?�	%F�T� ���g�G.�������0I�	�2
��
e��hYZf�ƶYQDi�Wel)n\�㛮!b��K����H�l�ɒ�u�e�Id��M,����G�[�O�� ;Z%�2d��I����9��20I��q��~3ǽ�#z��X�d�����i��K-g^nʨ�c}�B�.;d�,�հ��%� ��V�6�)�j�Ve��>r}�R�rI�ކ�c��}~0ĉrK�}�]C�a����/׃{Ll��m�m�w���IT�igM���@�%��4�ϼG9���<�"��1�˲�R���(2Uّ&=�z�,ӵ�wS,I#���H$wzfH� ��L\b�{͝��x�Ѹ�E��F5�R��޶��L<'�.:=��-�m��o���%���mk�߯=z�f�uEP�1ԅ�Sv+\�
d,���i�sZ����,c)e��7��k���]�����l�nc�A%i��6Ѩ�Q�X6��e�qsq1�}���hw�46n���5��M**mr�*�z��Mt/`�
[al��Y������V6�N��t�iXiD���Z^��f���+�J���\.�ɮB]3��"�b�um��1�����E����bU.T��JF�֍Q�[]v�kF�g�����\�+�?��_}��IYjV�N�t�O�
*1�y1��o[;'bC���6�����[{����&�s��_�9lÇ���w�w�X�{��Hn��H8������\f�fg�(�"x'Ŵ.�p.��"������v6�w���v�{{�N[E�t!���}`���<o�+M-�6w�$�I ����֦Q�(܎���ľ�Z��	�I�����Ѕ\H�z���9���+</��-C�����(]{&[;�H������-����D��L�f��]XG�Uk+nVa�èm+i��}���cu��;�7��$��J�2$�I
���\i�-P9�5��cx":wdH`�8}x%�!��:}�AR�{0�;x�dLY J�orb����r{W��8/N��jظ�⮯q�&{�ci�I��B�\�z�`�;B�����A� ��1��v� H%�]�L����������5����3��)ш*�>�E�$	/��Z'8M�k��}�I�Hf�̃�|ަ��ґKշ�TC�	�#�n��ݗ��sڲ=��jkgD�a��|�c;r������n���#�92O�b�6p�C��u���g��ᱤt��)i�*K��Ǽ���hF�d���я�A:z1�s���{P�D�QP!�~��զ��W ��cVa�Q�1q��ҍ��Ґ���u�:�%QǛ��G�d��̎j,P$�	��� �!������Z������̂)������A�^s�d�$^�=8��y4�OMeǺ�U�y���� � �g^�깻~ѴI/6v�(J!�C��<
깒H9���1\e�����K�U������W)r��<���y�p�	t�"�q����������m�;�{�z�V�'�,X?�����(���������D�$����.
tb
�#.�q/��mՎM��6�_DȒ칉�q$�����m�_7"��}3Y�JH*޾r�AN���oU�ld3y�$ͮy��.G2Uqr��N�س_�d����wȯ-�
�M`�'�u�F�e�l+��&sYs�a1�P̲����0 �w�8x!��6�����$�� �O2a��EG�#ou�m	�vo��<�v=��K%D^亇%BQ��,��KՉ��ͬ�Dd��I"� A1�{�`��������g_O)g{��[�Lsm��s���{r����w���A ��ĂIld�G��r�0)��H��Bb &K{�Q��I3����Q-���ӯ�)ue����$W�Ă[��dX�ޱ��R��߇Z��֎{:�6�R�$dhT"�)+jE��9���P���O��ȕ5�)��aI�
�(ء�+�l㙘7��6 �1Z@S�S{�M$����'F�5�FH^ϤuN]uw�[�z9Y��$	b�3b'�Ov�/�?�f�� ��4qXo4�\L#��m��w.�ƅ���o.6ͩ�~}���:�٧�@N�H7{�Lhb�wL�B��>ڇ�ͥy�m��^e,�z%���� �:xG[�_ݓ$Y�S�u��q�%����,���%m��`�7���ˉ3}Π8�� ��t[2�GnD� �Q���0l���,d���Ȑ	wtHQ5��]�x����r�쇝��w����9k8@f�Ē!�%��6Ɖ��޽����L��E��I3�W�`�Q �Y.��:�d���^��<�8���e�e�]�I$�}�-�� =�wٞ��3�*�u[v�µ�3�����1S����%~k��"��{�_�]��o���������)KG��ZX��7R��}�(�o�$�a�e��C���{��y,��l������t�}M�}�ׯ^��J�~K}~Q�q�n]]qhՂ��mv&2��+��0�o�l�i���k]M�.%-����[mlK48�R٢�Ie��c�0P�ˋ�V&R��jB��5�	�SX�#l�Ku#VŖ�p-b	�� a�ɊVD!��Ka�.�ݱ�AsH��T���n	�cq�&B���+D�ʛY�fu�$M�X1�e��Wm�I�冁�DD���>�qT�7=r�B ����UA=��������n�T�ęȹi"6�I*�g��]D�5�Ύe�Y��/��jd�Q�[[���0Ԋ���:��wsy�4M�.t��7���'�I��Q�5�6��w`�H*��A�q�n�8�� ��e��8vt��9�nXI;r�$cm|�hl��t�׻e@Β��Z�Y�v����]�x����9��D�$���LW�|V�g�b�HoV̆$Ŧ ���v:U��E��_�%Gf���-4~Mb�0cab��	`��x���A������ke*���s��~~�r��+2�H�/B�@"K�ِm����*��O�2�ųLTI59x0:%�9P%�`��vU��2�0�ؾ����;_�8��d��<����~J�r:H���wh9�KUↇ�wV̞��9�ݚ��7�~�>��ޛV���� �@�1�T��x��%�K�ۉ���.�;e�a{7��on�N7vO�("�T:��3�p�"o��IM��>�M��7�����$�������
���(<���*����>5-�`�"��y�$��,��%���şx=�͂O'�!�&{�@q��v5��H>d���#�Z�Ǎ��{�$[��#^��<���B�<��J�%٠�M.Z��\�щ\ꛫ��L�Ʊ�mb�p�w$v��!9��Q4�M̡�L�r	;�ȐI ;$��4Խ���m� ��B��]�P>�A�������͝-�i�D�F��=�;HdM�m��,dd���Y���6���8A҈ID_X��
�"��Uw<L2@�E�Ă�ckE3��5ܶ=����z�]������^ɋ���t�{=v�}r'E��2��Q�1h�B؉��Z'?�k�'�v�)�y?E������`���sw�ʖ��}��H��c���{�y��?n�vy��O��8n	B�#����{7n�h��g,����k�{,���(2�����ݸ|�����\�3���eqP�	׺��	��ܹ9��=}|�k~t�$��H?��5�"�Q����E�[��{	|�ޑ�AQ�˽7դ����OVw�_Yxw��������R�����w'�o���M2�^����2��Ι�j~����}�ճ���L(��}Ou8���NFw$i�c�kX�_v��Ϸ���Ϛƃcy�%�����珎]����kº���/>P8���*�����z�\�w�e7Oپ^���'������K�q ��V���~�x���>35�z,YۅL��,K�����9�b@wgg2�O��vٻ7�{pk�Ek𥃾ƺ��d��Ka>����h�������t��r�1��������wğu�µ�%E�	�5�Eޙ�����䷼H�vc��4����J�v>Y����W���{Kn/R�����9I�n���\��s4l��)�r{7���gfE4lȘ�x��wފ%�.�h���B@L3�%F��e�C���ˋ�Oi�m��O<��������8�J�����u�V��ᣚ��~��]�yT�J�XkF
AAE�*�3�}brh�r:�u��|~����������Y�]u�_O�O\�G9�.DC2TX�PS!�P��̓�$���������_����뮾�LoW`*��d��N�Rz�,�!�U�������|||u���������:��g���^��z�D�TU��UTF�̠���H��'�����}>u���������:뮺�����{{�5�9���<�N&�	Y�X��N�Y%�������+�1��\LMU��d�b�ҹˑ����ÖɩA`�媻I�����"�Lh�S����mY�$����Z1�]��v�$�E��sp+"�8��ȕ��dQ�VF��1q�1F1�;�--���kq�J��T8����11��������1�ed'��Y�y��.���&Y6�2X��>���w�C��s�rg�c����2�~�c@�2M�6Ǝ��^y�q��ǟz=A�$�3]�
;�"��sD�A����	�qC.z�J$� (�L� ��s-�������I��_0�YNRb��A�B��9w1mi�t�Q������5eҼl�ku����a�ﯢ8��@��=�,��y CH�E.�搩��S�^��=W-%��|ԡ���]�	�C�=�\g��ɕE.���遟U���r���/v���9D	2l~�&�+|�x/?N�3�,V�B��T{��ΫنH�Gܠ�mO;'!��-�g^e���j$�G.�H�$���`�.��d�9��>�!F�.F���	0� Kr�P-�� �������o7���罺�y�n��f\�N����_�����5 �v��c�xW�uc�e�S�\���E}믾?3�
@��&�`�@�l��������=�̕t��]���R	)�w������~���M|A�Rb�:�͚���D��[L�9��v��׵�ka�+�P���߲�"wx'�Uu�H'�8�(v�O��=J=�������y��O�%zi$BK���� ��3���T��}��M{=ޒ	<oi�e�;��J��Vxu,�d�zČi���tBrb�0ڧ���w�,J���}z����{w	:}�)���$�H ��;�D(xE�c�7��k��׌Z�3�g }��TH8ɔ{�}>!��Bjx�# =d�[�0�]��l� �Qo�>���I�׏���ys,�$�CKH����`��Q��8�pWZ��qDpE���(���x�z�p�pop�I��i�Kz�G�Ǭv��-+}ц�X��N5ȕx�������߇�Ŀ�_���˹G@�]F���@�R��� A��s�^�L.\��j�V�շ=pPV�������n����e�#hU�i�I����.Ωk/�Sub����H�A��T���;MmtIX��s,���n�!b�	��c0nLh���7�a3e���+���u(����e���-�E(VՍfG5��rcL�˂X���iv�j�J���%�$��y���`�jm��-L�1�Z׵Z�p�InI�v6L����ݢ�H��G��>l��HL�2~���<^s# yW$�/�ӍBY�x�vot"�A��3ۢJ�y�T���v�K�9bA����!v���2��ê���uc�q�4�}"�ю̉� j�#�fA|�r�d���6�������wHbs��	�(P�Q"�ic�,I���$	2�$[��]\�Q�y��+ovʑ�Ȥ�v�X�BO(��vn$}��9�zx��~8���lKI}�F��e���٭>��_+�/�(	g𼒚�9b�tlɇrY��Â��hN�����
�9P;��� �F2��$�{z�&������o�S�����A�91��9c���j�x�Ax����ؑ,�}rhꉈ�~���M٣$��<}����^ѳN+/���-�(Z�%��=0,x>Vy���F0伿�d����s)C���c�/��o{�*����s���'���2z�̠]�6Tw��!���x]t�FYC�p�1S�؟���Y8�R��UQ��O�j��ZKL�0�u�~�|+������f3�p`}c*Ŀ1J�e�A�BIy�H�m��ƚ���#7"�0#��-6ɢk���N"�#�c�O �K�����p�R�N��{�1%��˻>��d�w�bN�7��^D�Ek(1X~a�.ʲ�.�Q2"1�� 4�T�iB[MS��2�m�:� |%2K�_;��2{���#���Ar����#H��3[�;M��+�hͱ�Q.!��޹	��'TOS���Mq^��%���1���#�V��Y�z��%�5[<@�a<
�򮇆#�o{b��H�B����F�GU�Oe�r]�ѽZH����N�����}YW�L��z�;='W"�U�>ݴvZ�����p�FG��|�a�iy��O�c0c?��{�?�����2K}�3f�k1LA� U���T�%�%E�q�I$�u̱�(�or��^O�	��H�$�����
rbk����>>d���S'��oCCUF��A->�L�hgrWwLÈ�3t�:���	�h�4��k`�KsAk]��:d��٪��r:�L��M�r�����&ٻi����g�Wz�i�&;���j�Y�C��A7.Ep$�oXa�xIG��C�ٛ���hwўއd��ݘ�Z3zE�<��u��Ug�^�ס4,�� �P%���w�$�����w�#4y�H�n̒	1]��D\ys;��a<
�g���=�>"܎��%�(d'���� M�@�����3_�����zI�e�??h��^G���%�iӋ�O�y�$o�P�ce��wۏcj�c����p��4��+��«�lA�1���ꟷ�9�%���)9�=z~����U��I�^g,����n���_%�A%� ��fq���;�����*lx��N�^�����Ҳ��u�1��5�Sk�r+ʋap�P�ѼF�Uġq,�[�����;$���#����&}�ͬ�s��de뿮nE��Dd�i΋�L4�4WdBNC��wqTj9���2���&�,gwlX�J)���nĉkgr��@'̠'���d�p��!cw���b��\�$��q����OC�ud�ɭ楬��J���)��L� ϻFq�-F�:��-���pI��Ē	�����醩^�[V��Z�c��3�jʅ��9�h���L�B�f$�L�}�p��I�:�O�!��al�-��z��Ǝ�sx^������]�1�cZ��K��}�'t��}=_Y��?{��v��{m��ԯf�ryٍ����������0m���[�"�8����|��mBiC#�u���r�2�2�յ�����q!�wo�Ҕ��9�������.�K1��*�)X�azԥ�J�/WS]�Uטh����sl��Y��K�ƨ�c�˦(ưv�fk�m�h��u��b:����r�u�-��w!J��T���D��8�P�%�7�k��Y��i�+vt�LM��]-պ�E�6�m�iI�0�6Y��z�6�e�΂k��u��v-m��(� �,73�Ȓ�
w&��߅��j��1�1�F3�#��SH[��c��ૣNX3�Mb�
���|0�'& m�{�bA����^�~̓�����@4���n�L�}�����U��#+o�'!��;���;�x �7z�h�c4���@��%�21۽UNI.�����\���_��;�=+[cǳF���,g�\̆�wH��I����88�V܀��$kEoPx)C�xg���ۋ���{�1nwca6��+�m�/tI$����X0���o���)��&�h�EЈ�2a�Čۚf�bZ�Uו.Ω��>{�}�x�JA��W�$2�"@�A{�!���{F�oOP�]ֿ^O@�q�>�ɚe�/Vq\AN�y�wdM2��2��z}t
o���1�V���ـ�>��鮞@���tZ�{��1���g'��^��������7���,v��"ߥ�c�?�߽g�+��g���������@q �G^[�{
��{0����"���2I'�b	$�Nו��7��E�b�d7��	��l�˼(w+�W��h7����c[�E
` I�+�1-��{v�5*�p������g>�C��[�-�˃<=��zK&D;*�y4,�ٮ;����r� ������[׾1(���dd����8[Oi[Ι٫�6Hk��J�2i�n�d�3r���*O~�ہA�w]��{fCk$-��ò o&xvI�jށ�}�ȝW~���S��U�fg9��(� f��׀m�#���o�:�Z���+��-����$��� �s��K�{(xI"s�N�]�:$cf1�`A$��� �&[tk0��˄�,=>��dJ�O�1�9�ŕ��h]*[hk�Y�������uy����.�q>�^[�ת���0k�g� �1������?���i����5Z'����2r^;sL.y2&�Fu���9�bF=�v4�gt>WZ����F�}5�Evt�<N+�w��I,�����]¼z�K�C�1Y!��L�C>��[S){71	��� ��,�f��ì	cef�q0ܛ���1�V]�bl����r��ʁX�s% ��1��ǘ���u�ޮN3�ݿ��]�[du��Pa(wR��t�.�F�do
��}1�4!l���<�б�{��%��w��y]���?l�!���1i6 ����o��C��4r�b���P��1޼�c�g7�A"�G_��K�'B���@Xgڲ��y���  �9��a��B����:���yc�ħ�|�w���m�'λپ���{-[�`<`[�C��/ܫa��x,�o��!7�Lk,�������o������ۋ�9�A����*ĭ���$���>ߟLC��x7kk%���-�
v�7�YP֌��Kj�6$�O��G����ksh����`Ѣ ��GmKFe�V�r��8��<�h ����l�n�p`O�"�������eg�H�e���2�6�Z�-�� |._�ł5�c{9�M������@�P7,��"�p��x���4�`��	d�g$n޹�f�>�IU�0����	�YI%���
�
��5�s$��Ir�ٵo2��bۺ��^��|���H$�t4d���xE�5�o|v���@ɨ���jY�rbL2D����[$ټ�o�
�턲x��n�M2,�el�b�Tk:!�'cُ 9�]�:�����	�r}��}s[���ޙ�_�������_�s��PTW�� ��?���q�B  ���L- 3�W`$b1c��aT&!�EXdXaU���@	�f�Xi�@eUf��VdI 	
e@ i�Q�XUd)�@��� 	� $"aU�d &��Xha  `�aF� ��H�F�ŊF !�Ō �I#)h`IZBQ�� aHFP�� af	�� D�� dd�V����=p"@��0��@�2$�+@���� @�0�0�,�@��0�2�0�0�0�,��,++ @�0�2�!+ @0�,�+@�0�0�/�~��\�2�,�!@�0�0�!@�2�0�2�0�,! ���2�2�!@���2�0�@���2$!+ @����� @���0�0�	+ @2�2!@�2�2�+ @0��+ @�0��@���!"@�0�,!@��0�2 �2����� eQ `A e dQ `Q e a eA a;ޫ�DHHHha e ` dQ `E {�8��x��&������D��D��D�����D������@D�$%!���a����he&	PHHhdD$�i!c%� JD���b�#$ bŋ )@1	 b�` -4�
��C*�2��+����
���(���C! ��C"�����M2(0I#0�F �K@b�AVi�	�� �Bi���Vi��Ua��P��Y� !��U_����z�w���0�� ���A��������~���������g�y������#������ÿ�ޟ�Nq�?������G��j ����������(� ��� DTW����?B@�jL������?�D����0����}/R9������o������s�P ��
��bE`$�E` U�E`!�Ee�V�VB U�V%�$��VT�VY`� �!��V �ae`	RB	 ��d�H	�� XA # Y H���0�B�$*Ă�(	B* P%	�
�@��@� ��H�D(%"!	HI 	$��HI	�$ ���BB�K(��*�
, ����+ J+(B� ��"��
,��+(�)*,	*�ʋ"B+ 
Ȓ�̂��
��"�J� 0�Ȑ��B+*�+ �8��!�Q`%Ο�"����WOܟ� iP
 �
���������o�
��?�0�O����>��^�������H��g��=����~����

��������'��QE��C���?g�:�(���C�t$TW@����Ԝ��}B~��!��I�����Ä �(*+~�?S����0����O�;�>����������}�����?O�� �X|~�Et��N���E`�0���{
N.�����x�?�t����I��zE}'�jO���'?�`���~���'���QAx����"�//������_�C�'��(+$�k-�s2���0
 ��d��D�|@�  	U���@S�*T�R��*�����PM442��P�� 
 P��  CR��R����m����b����f�(�ʭj��-(�m��B�ٖ�]d�[mR���JV�����J����cO|                                      	       ���R���D�yc���� �QYj�\��1 �ڠ� �	iv� n�I5Ckh[�  *��튫�҇�׀��M�֡@\Ɓ�}��`*���� (�8 h�����{�t(���]`(Z���)J�ފ������   �         A����g=΂@^X)KϹ�R����e) / :��
��r�XUH)s �w�E���ﻭ�Gm)\ 	�ղ�����W[�u�iN����  yW�S�o������W�� y�S������.V���Z6�5J��כ=�i�� ���nw���a�jܺ�5�wv�e��i�[i�h� �P        =���6^���w6�g)��m�f��U9�� .�,��of�y��on��wvڶ�k��ER�\ �R�7u6ֶW-p^�5Ҍ�i��  �=_Z�;}�w��ڕ�p .�n�X���][-���M��7GL��� ��[W-w�ҭ7�+���y����e�ݵF�G�ES*+k/�  �        ��գns]��S�k�V���f%�붕Ln h�LM�a��U�Tr�ц˖u�V�w���-+����r��Z���1��_ �  �Ӌ���jK ͩ٥W 2�e���#UJw ���a��F�J��Rdj��J��d#�  x        ���0Ԫ�-�
�Ԥ�� uN �&"���"�j�Rͪ�'� �
ˮlҫ��Qʔ��TI�   <��^�r=#�� ���#Ue��U��D��T]k��Y�](�F�3U�}����T�!2�* �S���(2 h��S��%J��Ɉd=��L$T& hT���2�* �M$e*H �����?��p���3>g����f1Gfv�����@�$���w�p$�	&�! ���HB���$�	'���$�H@$$?���~7~�_����;�y���O4l�Cܻ��lʰV�W��ߥ������z��ʤ��໵���*é�r�/99��n��nAS�ȵ�:��L	�>C�É����Yȃ�,�p���rwר*����<D<2f�������y��ҷ ��M�{x��\�r�T߹��t-d�Ɏ�4�|5���ܟG�0�2���6`#�v�*��$'������{+׳�<�nLW�%>S�Ɍ�#wuET�gHC\�OInE:D��on+�d�H���˶�'4.��L�@:'N6���;�-	a��f��f+#��)5C��i�W��=�"�D��q�J�O�Q�;����E�h�[�Ǎk��[s���V;_-�T+�Bqvj��h!ƞ}]W��wtE{�k뜠���[تmY���jݜ��=�@qV�t��i
��1Ƶ�Y��HF��h�>�ۤ���g3�*_�nw�3���B�7m��k±�n�/��h鏸G� �q� �y-��໰��7ks��8�w���S]�±8��%~yl��8��5�F3.nַzJ����L����"4���8Xi�5űH*nC�Mـ�V/Z�yK��!�5��q��c�٩�XK�F-�>cd��bi)����;i}{p�)9�큼R�$�Nũ@�Mó ��ot�&=P��;9��봕�|��8���O/�ܢ�
%o��x��=ޢ\����n�ҡl��g=��#�@�"-���\����\��^��"aʓc_omX�)E�xV��C8��U��N��;_N4p��ވSy�/-�\�Ll�݋)cŜ�'{t�U�ȶ<j�z'2�=�/d�����0����n�ݗ�V�yw7_��U��Yhn��O��Rm/ ��%��U�%�f���sfE��{{�=�֘廅PA"n��7Rӗf3ϰ\n� k	��E7z{X���ݙ���(�(�1�D�N�"���CX�����O!�������<7���f@�Q
�%*��%+!^��Ź0�%��4gnۍqC�#�O%��j�m�x�YW��Y��MG6븴��(�u�_�Tz��=�T̺teu0� ��9�7����Y$�/ DF�/��r`\��h/�T'.��H���c]YnP�L�(���աHm��B�#�V[6P���ů�:�S��y���q��2��K΅��έ[3�����׸����R��֞��P>�G4��ۄ��E�1����~���	��q��T)M�׀Ŕ}�gtH(x�<:��	e���pvR2�gm�-��]���*�*q����h���WF���5Hk:
}��H���2Y�[<������-�Ȟ��X�g�2<x��ۂ���]!�J�:�_	��a�r*i8:����]�6Ӽ��ww���af�8��Q߸ڷ�vV��[�7��H��"=p>�9#4mü:jt���\M�P�59.����(��i	#�.]-�,XW��D'�M���v��"����+�*�_G�����8�N�������f���4�g��;��
�XE����t�]�(i.D�eM����52Uԗo��E�8/ ���,nme��Z���g�uL�w�G��6�{4h.�;�ƫ��gj#�����r(R�.L�Cv�9��9^��6X��]4�Y�asD8�@=+��.6��S�ΆdK�;/5rv�թ��M���9��%���Ԟ���S^�!v2�(=���ѐX����%9�Ю���Hr�\l�aM���F�x�wsj�B��}��l���x�X7L�u��9p��q��,dt��c�}L��g�5s�te�?
�r�4^��S6�˚�Х��Lj�gf�^�8�C�H�W�M��w]h�B%����aq�]]����Bf%���!*��v�=k$z�T8��ZC�`Pn�&�J��Y? U�oS�5b�ҥ+X] j�R��Ӻ��h��@wV3|Έ�����639��ַ��hхuFA�k���Ts]���u���4���h;�/nF��Y��9����Nc���G�l]�5�"z����8�ϫ�Y�m��'�ۑ8������5�3�T�@��7��!�wtە�K�BL�-RN�tdыvd['vGC�EF!4�L>�ԓ�K�M�9rXf���%8��w��:q��
�<�aQ�0��[��9<;B�&����5�4��0`���@�1���;�Eܶ�s�9�Ԓb3V�@TL��"˨�8��<r0
�8$�i�6���#y��r���ݿo+�ŧao���Z�E6�Yj����S����LcRd)K��w��aD֌��pu��1��y���M8lB�^Ȟ�=�m肁^�/	d�4֯�E��[b�3w��d�;�1׀n�LibQ>���1��;od�X��(ǭ���ڧ��Ey���˛��N{s*�1Ƅ�c��s��#
ͩ6	%"���0�A1i|8�2K�����D���E��j��h�$'.�Wy�%Y�@1Eiú�RJ&�Nb���tQ���f�oA6 �W�3��=t��+;fV�Yη�]�L��OT��ǖ%�y�+�u��
 �f������K���݅,�</$seڗ���b��v��!�'�`ŠX����ʸ���[�M�͆���"nqm�D$�tu�,Љ�Lx�oH˼L�_&��j�v��K�π��1���+����5�o
�Co�m���4�juY�B��:L4W����a��D�<�K9��pŘ�����źll����I;��kdp����tr/��՛'N�Ց��b겕�3�Yt�T:���$�`	��)�bC����I�4��'}�D�v�8��.�������(<}@[ ��<��ʑ=���ո�0�3�;�'wq�D��P�]�������ْ8 ۊ��v�`�u���{�O^��P����.K��u��tf݂��XI�����ddm�4�d�%�Mf��6��2(.��G�Iǵi��lK��(ފ5 j�!�O�S�&��S���Z�O�cN��֌��Hǻ8p�S��-N7n�{٧;5��r�)�~������)�gl�(�9q˃r)�(�Wߓ�>�`y	I5���1���<n=3C�!��m7�an�m�7�#4�^U�;�X�?��*���=84�^'���VÕ�������PP�T�Fʶ���Q�\F;�;����x�Qź�m���K�Fǥ�7M�U{��i"�1�g�j5Y�f�Šɔ�ᒩ�>3@��$Ě�w�q��'�4N��M�d�Ӎ�zm�P��E��fܿ�!e�#�y[ˣ��*b��8�`f�.�U�]�**8$�~aH��	7�j�l�e5�;����9[hB�7Q�0l7	��w���\���lFc������9�{�LD�nIl��7���ås����xB��Aۧ۹�[V*��o���v���Ӷ�9���બ�}��D!��(e{�c��!�*)�;q��/Q2=�f�I�1��aU�\Z4V�F�*��u�2�H�b����� �Z�h�̐�n��5��4������1,�,�(�r�IԶ
��~w A�f�;��n�D�����ri�l�n�.�@
\tv��;4�c���d�&,�q�8��:j���f�=L<�:�1�,�ui�-��T=�:�,%���w_r�8���#"���h�4�#hV-φ\|���X�y�{��#q�,knvv�V�pt�Hm��{�ͳ9P/\�4+��i�s��9��7��V�,��mt��
W����WWǵl���� �Z͂�w���6<�L».0���lܢlt�2L�s�����	�ꊅ:ةX	A�\�4�u{�%�v�nA@H��K��K%�^��b�ʨ���BZf���O�pG�'���ch�#h�q-	���́�{㎔w]e�M؞�����]l-�`��N�A�[ck�8���)bFL<֢ֺ��Y�05H�k\{A�T�����\�q��3�T9+H�]j�pDƭ9���d�m�Ct�6�Z����mCs�މ����t��N�������Nԕ)�C.i|��I֓��(��S�	�+Ń�w�-ԥ	j-�R�U�n�.i8��p�WC��U��v�'Q��J��KY�]���V�)��Q�����_a||�qy�	w�%X�
ũ�.M��id@�7W��nʆV���;y-��j#���uMKqk� ��S����
�j�N_Z�ذr����DA'$�h.�ܫ ��Ra߉H$�� =F�����{��<��-�yA��B�1��x��s��g�h*�Y7EH�&]�25���A,�JPdI�� eak�J�i]�P��z��T�bl����V�ɀ:)�N��Kሼ}���X(Vܧ�ѥD�y�I��D���K��8e8)��οH�5����ȷP��W�0Kzi(�xR'
Z�yn;J�֙#8K�����J=�%��y���j�;Vr�L�My�&�z��<4T����gn�Z[�;�=�1V��q�`}��	��˄`v�\pW��N�;yc#;5�9���M��SR�s4je�k���Qkn�;fv��ƹ�����:�D״���RR8ыԯ��4|D�Rעa��υZ����j�Ӏkz�noR���a�m���v�C�������Ʈ����tb1�0�;
\������q�GnG�<홛U<�a��^M閆je�@Ȑ�U�U�v�X�\�G{��н�ګTrЮY6\���wj��Q�KV�bN˅�B2ݡ 1�ѣ��Y��N���gs�x�Lzچt�*Զ6�9efc��*�ɲ=�{�;�����ZWD��4�K)݁>�Q0�w{Y���I�S>	HBm�*��;�s�T��ME�۳D�C��&Y1M�vr���G.�[�k.L���:N���s��Ӈ��(cz[�L�Ӓ
�H�ڋ�u2�vӦ���r�҉wM�1���ul�J
,�)��U�E���ȋ*�2k1�ݶ+��Vs�x��RN��:� �xin�n(͆�^���,F4��7�%q�P�)�9�7���J�Skx5f콣z"4X��q�)eD�H,�k�ZY�ώ��N;���\{�5��N���	��%��>w	��a���V^:���t�/mv\���t*
�S�[���0X�p�o�#�t�ϖE�M�݋N���Lj�U���n�24��ΜX5O���1�8Ș{opW��o�á<{k����`�&LԳnoH���s�,�Z~n<�������:ڢ�M�r�RԆ:�2�C��L��J����mdg���Ҕ�2�JL^����b��=�B�{h���x̭�{l���[ 0�"�W�`�q u�*-MB���fEM!��Ң!�]�$ck��8i�]�{:`<��39R����#��#_ww�7�j�%T�����"<���F$4�Aˏw�vRSv��n�	p�u䭻�ڲՑ#��[�`��M�⒣�¥eh��ڡ|q��$@k���sE�|�6��#s_@:&��E�x5j���`5A�*YVt�RK�0�VQ]A�86;ֆytK�
yr.c&�@d`�H���.wfTQn��C�ǈ)�N�
����܊��|՝A���T骷�]ʃM�m8z��-+���)�hB���H��W�`��m���`Z!yo^8J��q��!�wqf��� s����rZ��tՋz��j���w�lF|��LLpUԕ0�A�����5c},��OM���s���sz����i^b3��ʞ�PŒ�dA��^�G��;Ȥ�ӹ���{	���98ӆ����yu���P*�qm�������Ô��WaҞ!�rn�C�wC1V0�����-!��a�ఃǻn���N�&2K����c�����G6Ϧ�D�H�U�ޛ)�c}u������6Q+��rӳ�jY�S��\<��bYP�@�u|s��A��
����e9�ɿ�Cx����ev2F0�h���
v��,C���*˨(�> W7CD��2��dZ%+�hLj����:�z��yT�����˴�eɔ(�w��p�:۳������z� :�=͇�gw��fv3(���ۍ$�.��v[1s ��&r>Md��cX�5?�"32:YOgn�{�8,�g�cM�] %�qYd�f�^�k`��c��؜��Sf�,�$f}��M)0���7*l�����n=�wLw��w�A�����=w��p�e=��Y���p$:�8�����I'��$�x�M�s%X�7�u-���-`�p�
>Y�neթ͂�=���B��Vk*�����&�=�R�y��E; ]Jg����%�W2�_���ܷ���Պ�_w6�n���I���Y��yƊ��k�V4dh�J����f7om�eO"B�[�"�8$x
�����;��\A�p0�@�Q�{��R˖�!��g}c�7BZ�[�K}��sKޗ�ˬC��'���<�&�LWu�H^��r�n�J^�%Ѐ��WnW�t�K͖�e"nv:�a�H�%�&2]c�gy�h�q�?���H�E��BHRB�	@�HP!P	"���H�  IYa HBE�$$�   BIY	Y!"�) H)$$+!$��
@��a�E a$��
I!$��$+	"���$Y ) R��, H��E��X 

a �a �R��*�!"�� ( ��@�*�� $� �H��IHP��$�T�
�XD����d$
�@��$�Y$�H���d���B	,�B@+ V"��X�Y P�
BXI"�P E I�@��HH�B���޿��[���Ox�wf�]g,�ηf�]*Yf2{8��h�G�jǻ�!mܼK����U�]X�0s���{�-�7&��}�nݳ|66�Y5��U�Z��k�VvV�5.⮑��]��=��x>?n�x���=�I8���t�ȫ�/b����;r��kup:�b�Y
�����n��}�΃=����7���^��x(]�M�,��᱋p��@�6ȲGm�"����?w���"����}���ǝ�LNmf��m�����c��E��a�G�v:�i:s��Pˬ��`�$'�c[�@��Gv8��<�IL�ނi�,���.�����/��{h{Occ���]�&ܱ�#i����++�emc�o;9w[0d� /���ox� �jB<��{���?��p�$.g$Wk�� yg���{7����*�f��WWø;��|����)À�����6'�R��_v���'�Y�[k0t�=O�n*��Mtܭ��#w#J���_]]Q�˽�|$[r�ԗ����R��t������}���=�X��Lݣ�O��i�W)q�t$tu����t�<­C�T�{R@OO�t殱�"��w�.E}R$)�	[ݺ�H���v4�		x�L�Th9�!���}uL�KP����iYY�U�,��m�4�:39Y�VMU���T�����<�����yˏ�O,��qs
�R<��l�)��Xd�/��|�|�my�����8��{k���y��7���o�������vV�*z�j+��s��/8F�AG;�I��ܘٛ���m��fu�s%k�4�@�ޫ��+dR'�5d�+�O�֗�9�P��>Oۖ�ݔ/��20�I��L��k����\́�@�R�ͺ�PwV#e��;a9:����%Q̙:W�� �DX���Guř�r�v�]tQ�Be�z7d�[V�=��ڢB&����Z�ɮBP3��.e��]&-�u�H�hk���=���J�|A���c���5�@Zw`�	�r�s��n�-�߅!�NV�w6�u��z��R��jx�)�w��i���}+���⦥9-���u�4ڳ�Ə)1��$=�9�ksd�.�7���4X}ov&���vD|�%�srq9�:�޴(�8:�D�E�Ӑ�7\�&�� ��6��YkvD�����n��U�Ő�b8�v�:�{e��|] ��[/�PtƦAz�+5?f�O!�	Ƿ�:NJ!.�vE�b�v�%s��.���|��Ǘ�כ�Hp�mQ����KF����1��kc�v���X�6��Go\�[�bY��u�Lp4���{W޾;PN��iV��f��ѯ�4)���ud�����<���հ�{ٯ\�&�9��W�+�H�JQ,2�
���4H(��\�s�<�������?<�q�a��4x�+whJo��0�%(���[�*Mdp����R��u�	�$���������v��T��Ñ��r�dt��^��=�y�:��b��|\���$�r\�kw��밽��RP�͚F	#�����'g�-��(�]�V�<]n�E��P�0��×qHE)�}���z���N�
�H���짋+}��$W���ZO���`묮T_~k�=R�|�� +W���mu�ąuwq��+~���S�#^��Y�M���x�J���j�+�v���\U�[�S�`��,`�*m��f+XT���m��.>�"��=�
rؽ��X,���{��/q1ON	/?w�H���hC�S�.'���{�ʖb�q���9W|�7���D��Wl�C�'�wCA+3��2:�j��N!�>ȩ�s$3&�F����tV�`[��//::4p�S�W��+�Յxwr��O�G~��1w�)Np{ugo�(�4����`������{<������2�pq勵�Fz5�s���Ii���o܆�%BX��O������W��g�ĝ=}S�>�Ϫ.<�ˢ�Z�])��<M�~��7p���d�)���'��[y��^�<�[^//?*�z/#<��sQ9�b��I�z�{�.����PǯKۣ���崕����@Kd`#�Ҷ�����N�����5c��W�����������&���X� �.wBV��⌾��͚<��bI���yy�젵|]
>�}�t��s��wr���0���YWHjޮ�˶0_D�Ԏ�<
	��Fr��◜�U�|���"η=����"���Թ�jy��$	�w$�� +;�ޘ�l9�{%5(��+d��d�,�$]��@/��vՍs���Mo]^�[*5�3��oz�m�W�yv��ҪjF$c%;�ɝ|BTB�c��ǧPAI��G�:�K�23���+G"� �\U�^F��Lݫ���6��u듣����>�ڑ�?mu�����V;\��E�x�x�tY�\qr�َw�܏,t��hإR��ϛ��)��VF7��F�x��c���n�d)�7$��Vc�L}�F���G�s��� P��ۘ�V��`��}"7��h���+f=s��L��xN�f���Z�Z�����#`�����}�wQmW�K�j�N��R�qjL�:�b>yvR�]<]�Vv;��n�s���o�/�u7؋M@��ش{f-RгER�l�h]]&�c��r��ea}�X�/�qr�m�(�d>���X�.�k��qyk�-���O��0b��l_"���jW[8n�!>���t���gu��5����b��6q��с��~Ug���U�2,Q[p��L�7y�-m��3���Qg_	5�ߤ+5jՉ_܀���go�5�W�n9�3V}M��*Q�ͮP)�u��:h{7hDħk@+V��x�M��:��js�gɛU�JwzgnSR>+�맺�����y�0�뻏î���K/A��^,c�k6e=�	�:R~c U*SM����51�^����g'���w:K|a�u�pi�� :�3=�VV�T�4B��y�qX4vngn��M��|IY��y�k���K��w(C�w=wRojr=Ѧ���
�{�[��,�0Q�+[To]7�M[+;�ꜝ��6�k�Lދ%�p}��1U5Xn���7���,F���.�h���YUo=A��9-�ל͠9�v°_WKWϦ�����P����R�� �=�0����u۳�ogM �C��r��ұ�z���l��<�W��ra�����}F��%H�jN��va�Fo<\#�qg]��N/<֞~��G�Yݜ7c|d�����̶��wq=��2�*U�k���-j�h�YOGB�z9�b)�[�v{�ML3�?m=GW���r��V�\�S6��DV��m��z?p85�Ǉ����Qv�/�+<����Tp:���4��׮IB�I��l-��L�T)g��^�m	�9�}�kCf���{\�<�5�/�ۑ�Xr��Ż���c�F��ٔw`�5�n�"� ����@w�A��ۀ�Y+����z�|z� �10�4Y9��/f�;A�ryd/��ERH��[�gr�g����ɼ���b���S���{���)�^�x��������}I�01~�C3�75N�`�p�=�Ȳ�v������͹�MÀ�f�7;G�Y�`��AWb}��w�m^�|�G�Bm��o]l����i\���+c��uTi�^�;�
j�z{_��x{�k��n��؍'��7\���h���є~)��W���9=Oi��8�ل�]�yUkA���%�;�#�A�ǹ�yu�)V�y�s��;I|�Xs�B��0���wi�h�F��c�����w=��K}���8� ��
�+p�N�J���ǥ���h#پ9{���_<&�9�gT�\Hz�^˭�<�\��E�(z���{���V)h���U�(���q93B�*��vg>E�^e��f,������s����Xmu�:s+%�k)�ṕ��/i�*����K���gˇ�v��KF���V]����?�#ȸ<`��0-���LgK�[�Ч���ہ�𺃻}ǈ�/L&Uk��a�S�Y�p��E�@-o;�O������R����m�@�B�m*MG�s`���s�f>�HV�];q�eq��zv!�Fl�-D��J���jbE�e��8��F�e�Oc]n�t���]2��y� �HDɸYF�jh�8��ӹ	ܢ��8��DiR��7-q����p*uj���䩳f�B�҃]b��ES�x2I�:��)�绸O"���c:�����h����r��fgOCs�y��Y	�+W)��w��^�ے[�6�h���Io����z�Mvnp����n]JJ��Μ*��K��T��@��O���z�31]�
u,�m�Ȅ܉w����W��.�g�/G�0�>F]�i���$���E�a<l��+:>4��-�� abV^�aWo�)�Nr�&��_�Y��4�Q�=%����n���҃��n�y���$N6w
#�O���\�)�^V�*�oe�c;���:j��t�YӗS��ܷ�O����kc��_�RiS�峐�{�Ayew�}�I�D|;�/i���#��O$� W���_1�@3h��]]�+�Q�df-��a��;6A�0�HR祔E���專�<���yiJ�<j�����[��h���� �p2��HE��7�`��=�yL
&�U7�q�(�Pq��兵�X�0�<������	P�c���zo���a�{CSv)�y���
Ѳ�ޡ�Oȵ�u�<l�)r�jT�{��5�������ze�c����F����p՜�,3r��V�~p_�qg�;���!'���_n��k'�&�T�. 9�Fl",|�)=+E%�$��+6�ن�h�]�繰��Ѿ�X�e�%B	� �xMxGhA椥�2�V]_S7�p]�������K����w40�]�v:Wnpv:�8eq��f'�� �-���ub��ՆQ��>�
��4��%�o�v�q�~Q��"��0K˯D3УN!�^wf_�>�b<J����2�s]��yE��GV��pmΫ�Ӱ]�E-��,��W�G��+������л�/��WC*�f�f�8��IQ���-���F7[~�7ʛ��߅Q�\��n�J<}zk#�Ç?G�qC;x���R���؞�[@���I�u�A��{.g��:��n�ү�0k���Ґ͉���zGݰ������}�-�k�@��jR��3��-ы�<�k��q���9�l$wY!�}��c�\
S/��qԓ�B_��5>@�>n%��K����9�+G(ep$�^|��>Ɣ�3Mi��h�CsR����1��.8umӰ�2��9G"/�F����އ[�a�{ԝU�Y���3]%�@�=.�^�5ʌky r,O�\�!�RVY�oo��^y�d3T��.���9�r94�ս��P ��0���t��5�����x�/I��r|��ɸ���W>No�c�۠ݰ����*�
��ә�MS�MBA�"�/'�f����Ӟ���"�p��!���lU�q���9٢c��x�׏ �f5��D�u���ҥ���&mi��Gh��obx�S�[˕��F/ӫ���v]<ϵ*�f��/{'V�o�ɂ��6vڜ,��!�1��U�0�]:���:$vq.�53z��|@z�t��Қa��3jo����}�B�&`H㸱�U���u����Ksy��$6yu�R��5:�TY�1b�P]7���-�����z��e�wrp{�{�\������y�yG��Վ�m�ɕ���{�-��q��n��!-����x/u�>Tw3Բwz>���)>筣^��/������fNE>��=����Il�OHr1�[}�S�\2f��a�5���B\}��i�k	-S*޷)@�9U8�W���4��_����#���m� �ur�,ڭ���x2�S�^��<n|��\g&��g+�\�Z�w���crC#�R[�#�֛Z�#S���s���X�k6B �'�qQY��墔|��N'�N�t@5>�Ư9��0���q'�!E�JR���ya��̽������*��}z7C��	�ӇT5����8zr�e��g�!��א;qD�	o.*ޗ{��6����h���y������D$�*���Q�/N��$�$Ҭ�/t>�iFr��y|�B>�9�(��}�Q�������a�71٬X-���=:�0fY���墶�>�
�>*F��#�k�S�܌�����~���!��Ms{V<3�t��w7�̹������*��f�����|�v�|>�kK��H�x]��U,�sQ�٬�<4�B�ᤊw���ө0,�6��b�A
<�N�7ze��/��q�q�,��:�{ό���T���J|7����xď��>㚬�\�o��=�s��Oļ�8:����6���-�K�3���gU�z�Druq6қN�n���ʎ�X'N�w���X�C���^����QIg[�5��}��	�S|�G7=�W���ł��cۻ���5�iG+��<�]9�Ր�`Ǉ���=6@tx{���'�q�*b���ԯ�F�,��v1˶	���p���i�����������?>�����qx�t0������X�/j��Jm�F�[Ymu1�0N�R�%]��Rcx�u�FMXz�ź�V]�dP�frnV	Ԫ��p\�
�7�c�)on$�a�K�����;���&#�6����ed���B�c�[�rw{����&�J�:2�\d��[BP�
��G�~���@�~$�~���5uLӬM`ۚ�.n���nM�\�-l �@�Ҝ,���N�M���P�d���uQ��+.��{t�y�Z�<��s�t���F�\m;v�o�u�ݳq^�N��nֶ�g��wA����7�mŶM�;zb�ٮ�ݻN��M��0a�����n7e�nd�u\�1�g���x�ewC�k�q�^( �n�q׮��k>���������u��g���=�5���g��û]c�gu��㛮:��}s�g��c���c�1���A��D�.��W^�\u���&�f�1�n���'��v�kn�h�!����ݎ� .+M��n4Gu�ûW��=�
�`�2��i.ɛ�Wt�T:�l�����B��.���;���ٌL�����w7܎^��E��y^���ڋYM��y˝�Ws綠I��pp��!����t��ٌ�q���$��gc�M&����g-����/wi\���Q�n�Z�k]�f���غn�d��\h���q�#3v��n�tM�z���{e���W���[b'n�spI]vm'U�Q<:�G=r�����*v���޳�ex�Z(s�v=��&-{mј�hy�Љ&��]Ș���z�t�<�nٍ��c��6��[�v{j�q5C��+u�;�]��zڣ���tj��s�W;�X+I��@�Nݮ�ϋ�K���7u�睗%��w�n��w8,h����JK0n���]�\;�J�wJ���T"{q�ݝ����-x��x��%������W5�t��k���_g\q��"�&�ݰv�ᛋu��pG�������j.�۫�>W]�v4�QX�#]����X��9�l;u�&�m�㛜�<�y�܍��l����uc�3�7b���<s��B��d��&��%�WX��NGvS����"۫��rq7\=��>��xP냶֌/n�i^;^3UL�z��o0YƮ�lk�kp6�A�l�t�u+�!��V,�n�.׷D��\�9��n6�tO��׉7V����v��� ���g�ut>�o>��F��P��ۛ"�]�\�+/X1�8�T�ɹS��'Y���'6n�S���vv7d� 8ܽZ�9x8���@�:�:�ey���,��c�n5knm�3�q��{d���55��u�w>�ɸ���ΛW�X�����N:��/;�r];6:�����������ó�u��`�wۦ������nӘ��$�y��F��nh��<r�X2�n�U!�@�眝�;y�t0K�m>^δe�r��m=��vڹ�
Y���.��ka|�{ƕ�ޓ۟;z�y��,!v�l�
��ݳ�mgF[�w=3S�@�^�k��������`����6�����nxs��9{v��6����4�V�r��!��X8�]<�������kj㲼iOk9����[f���ڻ;Z�\p��g7k���K���s*�5���u؎b@���۞|��Űo�.ዠ9��軕;mO�*�G��6���tq�����q�h����=O�Z����ko:�nvm�ݚn�uc�Z�b����Oj��bݣ�4�0i���u�nI��1�NY���`�<�f�h���z�F�{kOd���-��F�vm�hO>k�q.���A���ɥ.�+�g[E��9�{��q^ϧ�.a��F�l��tu��װ��v�zz\��T�F�ۺ�s=����oe���{���fў}�7:ܦkZ.�mۅ���א�,n�g;���km�U�|�r�8ͮ�����v�(4��ۘ��L"�n!.���sX�j����c����g��e�	V\�ǐ��4��r��[�a�v����p�Ä���]���v2��q���uZ|O�헬v��l�6J��[4g�:ۍ��nc;�'n]ڎ�vڸ���f׮�ۮ��,ۮ�Z맬'<��gt&�y:d7m��0:��^�5�ǰ�Okm���n�3`���kui�պYL����u=��f��9��F�d㜛y�`�'a,hi�n4��ػj�W���mq�ݻu�r�t�:�9����������nƷ"�;ǰ���v�m�m�m��{sv�붡��l��.��ٵ� 犛��91c�������M=�=n5qQ��ų�N����[l�pQ�\�on�FM�b����&�=ˋ�#�>��;d磐.ݐ���5m[v�$*&�+0@q�L�2��[���۹=g��/n�ہ����`8�vr�kny�ml��2rX7n;,d��y��@�61�{l`���<s�$g��}��=&���Tk)���e'��wF�s��iv����k�=��_O��$�Lh�v.n(ۍ�/g&��s�-v.n�;s���z�Bۮ�k��-݁�Y�N��2����pk���n#/D��\��L��8m�Ȼ���1��ݺRNܽ������τ:+vGG&L]#άp&�an�&���9w:3E��m��oX��\�'/9�s�q]u`�b�v�sv����{=����]��D���õ�xwK��Q��
<Q���;�(>��x�&���c�g���Fx�Z�l���!�(usƳ&ٸ��J�kn5���(�99��v�r�������۝Y:4[p�6v�������s�nۖ[����UV�]z�7�N�:��ݸS%�.7�	q㰞89۳q�v<zM�K'�F�d�n=�^t{����q�%��h�8�4d� �˸�o6���%�e�._�m��-77
nռy�'^�n:�'tc��yz�z���n�v�d5<[����e��r���W=��(�u/�g��j복�]�k3�%�1�s�{��o%��JZ�m��8	�p۵�۔)�#���-�rtp��N9�Ǉ��v�klg�g�i�tA�q��`M�>%�Uw\@/V�#��c2�n���i��ƽ��͗��wb1׭��v��ˎ_\v�\�����E�xq�w���Δ�0�ay�c�i�k��ɜ���աEz���z�[N��[j��N�u'5��'��9�ʈ݉����pPqs`p�zأ�v�M᤺�Z��ۆ<,b�ۇen��t�Z۳��V%q���n{�#�!n���Nx�W���u�#��ۓa�;�-��y�Ů�@���w'"�U�������<�b�u��ً&�0rr��od굵�PK�vE:��x�[Γ���V9��ݸ���p�m�v�ɤm�m�^��5���3�#�6磝�wf�ѐӉw=�m�"��<�r��`��r���<X��V�P�����nn��;]���ƃ��\R��n�m5=n�@v](;\�j�>��=�����9�,���u��]v��L�fæƵٵ�uy^$*�'[�Q����)Ńmgqi��xx�<m�q/��[�ۭ��j�0���w�ün�Ζz�nݞ��g�Olm���n�0�烸6��;���z���/0;������p�aݗ������p��%�����}����]��֮�-�c�o`e�V�"�c�\�g(�M���I��W.zܧ<nS��'d�Ż�l����b�hy�<nHE�[;l��JR8wg��Rv��U�u���ۍv�Ͳ����k�S[d��w��ns�`Ә����5x�Tu܏$��ҏp�1�w`M�1��]��We��=[)nv��.��E�;YػcM����n���{�;pngv�3�nޖ�9�d ^��"1,�<��.��3k^�j#:��ػ`��j�7f�>Sm2=���E���&��땶���[=�F�guz��Ʀ�s�uOn�y����;r����昈.|l�n��
����Wj8wo���m9�����Dn����wl�[<����ݻ���b��o]�&����p��3Λ���Du�]�sq���{=����q�CD��m��{z:,�m/g$�3���<v�x_^��woT�3z���nٗ�쑘���kfƐld���FHn�L�sɽ ��lG�S�@v;l<�U���t���<�������a��m����e��#k�l׋<��� n:�v�8,6�㱭r��<a6�Y�n�]�vꮶ���:���qe�c���f�;���cs�F62�ݙGv�:o]I��۝P;%�J9�ۊ�c%��`�`"��G9�9�8�7k�>n7A^:2�sn��Cg�Z����u���)�ü�nb�Yvq;X�&��uY��7ulKӶv��SR�<�{^�uLӲvm.�=�޺������5�/��P��Xy��۝�p�P����x�;-ɜj�]��K���;˽[���v�+)s؇�aϤ|=��(�v޹�\Oc�K��x� ǝ{4�=t}v���h��z���ez#��(U������#۷.���7^1��������{GI��i׌aY��%�8ێ"碝ۄ�m���	�i�rܧA�kv�3u�,�V��v펼o1gE��Ok��Ӻ΍����Cn���(�������HX�vc���������h8N�uؼ��J	s�cn���Û��q۱�z�"v]�έ�����`��b�ɣ��7d�KÓgjl�'
,��)6�[�xک�S�&�9��L�C�j*�t��;u͋eͲ�u鶳�U�k�1Rn�[c�.9�{[��c8ᶸc\��kn�n�i�c���QŨyk��of;��2�bM�m�J�gl�<�8�iv�5����b�s��ے�ݝwc��;Y������[�6����֌��\8y���O6�ͻv-��q�zp�2���wf�z�q��<����u�)$��kZ^85v���)4ڼU3գ�=�����p�Ί�(�H����\�t��uh;qh�Ɗ�],�5�MKrU֭\��������c9cn�Փ�1ԃt�\�.n��e��#1ۣ=���ޞ���i���:ыZ����U�P�����e1�"�-��T�V�̥���̦\�b���+�`�D�Rc����Ԧ���
�ŌTb#YR �Z�n+Z�j6�-*3s �T�Z+��s*��+��"b\������2�-���U��Ш�(**�&aR�̰��Z�F����QL�"����`�]a\�u������KZ+�5�dAc��2�+��d�PU�e2*
,VEVV��2�e�"[X�V+[�QXj�Y�5�V���er㖣 ċ�e�E�S)\��m-�F�Q[T+X�����F�-����V*�4n[*��f1��A�fI���"�X�E�vm���x���O�p�s�6�;oa9E7�c�M�h�̹��*����V�70�Z��Tī�(�5����Tf�e�t�Tt��a���T���a��Um��J�ۙ��*�K�����Z��+b��$���浙��Љ�.�tsFòjrVh���8��W�N���>6?7a�9:Hgn:��mj�l�\��i����x�k�ۃ/nw�nl�f�-�Ϸn^ظ0�m{g��0n�ۆ�e]���9y���P��E:�����!.Q�jb���Ӯ|bۮ˃����8iN#Vnx���:���[x7/:A+�YJѸ\��9a�ؘA�=k��dI�d���tc�J��� ��<�nx�Ĺ���1�z�۷m� :���WD�R܎T����N�m�]����|��=��[��=��u-r�ngUܱ�C�>��W�w"'`̜r��؇q��v���[v\�K�;1�����V�Ħ�xg����������d�sx�v��c��wW75d]�6L�؋���)���7R�\9�j�=��6����:w�^d�k1j�Y�;[<{�qK�-vq�6]�W�7�1ä*��[#����v�vÞ�x��ƶ\��ۓ7>���s��;�m��t�'��	��� tP�� �ZۯN��`٧�	��H�#�-�L�흲��GY�����b��A۞s�����4v*�Îx�*I�q�E�����cϋ�]��;���|�y �v�����5�1�U����p!�ؙ��3���Xn��[u�v�z������<r�YL*�;uĥ�M��l�hd���ێ�����1ی[�
9KHt�:��̤�ٻ]��.���+qG�^�ܹ듃�X�I��u�n�k���ݦݦ��@#"��3�8�˓&�k��tp����b�<,��9�l�A��v�T;E^ٗ��뵼��z�/F���Nvwg,�Y�>wf�ȁ���\�<�V�"1;�8Nv�tݜ�G����ckm�V�q���e���k��wa|c���s���w��lv�q�[^G�]1�)�a�=v�ƹy��tn�C��uF0t֝�ۣ���jtk5u�3v��{��ݴeyq���yó�v���&Le]�c`2c�۝���n���*�ǹ���n<��y��^xÝ��c��c�x���4�Ɉ�aVզ4�1D.F�m���ʋ��-WA��8`��mɳ�m��)ȧ�z��W9N2v�˶�+Î/���`x93�6�G��;eA8ۃ���/�^9Q��6�\�p�2�LmiJ��Ɇr��SM����ġ�%#a����Q'�CS���B���߇:��5��=��_@��B��~L��b��zt�~>ut��k�:��q?gt��{�(�P��N]�)<��U�z$LI�L�vVΔH�k;eGb���]U� �s=������'�&Ѝ��Hz��J�����G�:Q?H��P�H'�mgX-��
�o�"��|H{e?�|J)H�'I��N����i�W�N��$�:P����J�A��u_�31��{Y����6��2"�ܖ5��4݌����1���OC��P^3tw������A��!G�^\�I?�l���Vu�ƟI�����zT�L�8A��A\.�d��%a���糮�?�2-\�U��=ݧ&�Y1�s���������,򡉃�ݨ���D�;��@z�?e*��.r+���G<;��+��w��	�6��Q?��I�s=��{��9W0�~�C,C�t(zv�� %�� .cKtf&�w�/OUK$��(�O�}�v"N[�"bl��d˲�t̬e���]BI�}(��?k�۲A?f�k���w��@���_<�Q��T0Đ'�U����z��>�-P/=�WēϳlX�gt���jW��.^i��"���:"�ڹx�<	۵�9�n�]l�M`��-������zR	H�5S%|H$~Ρ�zQ9W����m=�o}(I���ݛ7OQ$I
8���@�Υ�uz��V��I>y��$�gt�IޠǶwI��5��JK���]�.��$��|�ޕ� �]g������e�]sPJd���u����Ȥ�������T�P�o.�����V<{D�v���H��5d÷�����n���-�m�Ă=�ҁ
��e��Z�>�T�D�tLxH;:�œ�f쯉e�Iyh����޻��vbMN�%�=�����h�s���H�]�k\��C��߀�׽�<߭w`����s[�7]`��܇^�6tl���=�l�cg�q��
�F*�i1�\0ē�.v]��77eH$e�W���B����$fwJ���)�[�*@�٪�(�Y8*��ڕ꾭$���(����A�VL3`��g������$��j��\�H$��`�������<��${}ҁ ��vt�G��P���0���{;�m��������Cu��$��(��~~S޸��v��}��;}��t�G}�{�:�R/�d�J��I�*dm?V�s��`�P����!խO�n���wK���[T���&m 
�вɆM���J�G�fݬ��Ϋɛ�����*Q��Jq�u�r/y�T^�_niJO�zL8Xn@A��Q��.�;c�ۧ�.v��9�a'G�n�����?T�K����zP${:P�H8�:��N�8y�VQ��(I7�ҁ�<=�ā(d���vA��Ղd���y���mh���?%T(��7Ew^��LΛ�#�p��o� T�K��T�(w�:����BYÛU�ћ����X$����� �L꿉��@��IBJ�3�;�`��6*V~��&V��5@{��-Y ����D��%�a��X���� �o�Q��@�"�@�uB�'�3��$�o�	���xX�{��_[�֟y���v,�2�ް��%�u���f�{;�N&j�a���G����2(�^񘯴g%A걷}�5�9��oF��U�0�۶��5�kU������0ۑ��j���]�Xq�)����k=���{G�Бt�M��a�H�uv5�<��ҭoD�E�m�{v�C���'2;`�r�\w�mnϤx�\���=�z���8���L�{sql�7=-���0o&��ѳ�q���[�6�]�r,
m+sh�@�k��0�ؠ#�'-v�`;\�]��g�!^8��mΧ����1��h�2�������_���y�	��gT�I�lͿ��I'��w�ܝ����Qu�Q}�6�|H�VM}%F�]�7�ٙ��]�z�nz�`$�����==� �̑f�Y��/{0�1��h$	C$�^��� ��lU��<��H��h���%� '�J/F'�O�@��`�N�v�kr<'�_]������2�a��x�|���+��`�uM`$I	*8�ܹD�@|"�f�U�މ���7~�o�R w{�~#/�P�&���)iHCH��e#�^����wF�,�{6�<v��\p����ps�γ=��P���B��ǳ�n�$��M�B���[A?K����I��[����� �U��I������PQ|_z)�B8.�cʔ����:����;R���ȓ-
�Y����j�u���	�뙔`&>��tLǂP�&s[Vn�W��ِ��M (
ӳA#/�Q��w7��E���y,j�B�.6�2�~����/�(�H#�-ۻU3-�����w}�Wă��(��xz�Qā(d������oEm H!�d	=}�Q$��޶׊Ӿ՝
�^��;|1?�~i�
]�j�� ����kF��1�\�/)�Y�@|9>͠	#6w���C����啊�{'Yȋ��t'`��F�s����'�1���neM�/N��6y9Pğ���D����q�˂�}��$�;�f����!.����}� H���� �w���'
�������%ۻ�<pr�ē��m
$���z�[g�i"��-�d����p��(�c}�x~>}��$�j��{F�t����o6�b�����LV�=Z��;7w���޻�����ӧ��L��}��������QT5��K�z	е��<(_�Q��}޻��,j�B�.6�2쩽=�6���H/��A?c��������'O{���i �˔	�<6�QāF$��^� �F��P=�j��oVL���� ��/�_Ā}��F�gzجrwˏ���ϒ�N7�d5a{b��#�]��k�1��x[��tV�۶n������|��
P���'�ٶ,�� �}ҏ��d�θ���z���N=λ"���H�Tq�{.P'����!+C+zx�Y%@P��٠P.��lv7�tx]���&.�o��l�I�t�A �7�-V�� I7;6����J+�-'L1�F=��qr�w�{ʫyT�$�W�P��͠> 5�̞�W?eA��v�����U,O Ua7��9H��Jfʛ� ��9g.uIb�����&V��T�����/�yd;��5��y��u�sr���KQ��ć��7E��&]�7�'/�Q2��I�o����H�N��T���Xg��x�Ũ�+��p��������vۮxչ�X`�Ҽ8����rb$�	pD�a���0�1$	��}�+�;>߀�����}Hy򩢲��F�${��D�_�'�O�@��`�uA@�v}�*��_"7wrM��߀�T]�@������m�������|��AQȨ�r௉���� I'��R�r�vڔi�J�ĂOw�P'�N���@�wZ
0�Z����Kr�+��	M�J ���P�	'�[�&�����^@�w�J$��M'L1
�IGޛ(�	>��n��sxr9Dvzை�Δ~9u�w���)�CJ]�%K=�z/<Ɍ⊳ۊ�61\�t�G�"fܦ/PҲ�� $��T}M=T:�:�V����)��2��a�)�8�;�[$ۖ����s�S��w&3��=���ں�[��q��<`�����ĸ�puv�I@�mÍλW���h�c�����ck��j�f�Z��Ҿ:y�ǆ}�`ڼ=� �'V�s�>{J��L&@�<����d鼵d�ϱ���/�i�۴���Neݹw1�v�c�>�Ln� �
����n�j�dR뗋��v���.Ѩ냞�n�m���H$'��Y:F�����H�L&#i��S:WĒ^�I �ޫ/=����>�>t<��}Ҿ%����9�I���d��4�x/-���H����@9u�V	����^֫Ӂ>���le�
]�[u(�H;w���d*,�m����a�ۛ(�F]�]�uH���%�o]B�u.��x�^��H ����'�I�{�m��$$����uX
�0�Z�kݷ��A�t��������xK�]
�2���>�t�d����].��ǲB�'[a�:ļQ��:e$d�i���n�tZz��q�����o�ڛN�E��>��~�Sھ ==�T2�heǊ^�|�G�,�A$z�6�3f���	��f]�
��W�<��{��>:�'�T�ة/z!�E����_z��3Y�$\�Yƕ���>�sW?I���v�M{=����:C�֯�0�Xt�J���E�rN$ E�/��٠|;�~�yg�z�!?���JĐ9���V��A ��vVУL~�c���C2S�Z�W�(w�P;x1?�=H���uOeQ��2����$��H#kz]w��j�r㝣��ۻ �uH�F�$E(�T�\�H�v�ҁ>Hq���Y`�v��H'���~�ޔVP�.�!z�(���4Ľ��m����])�������qm�XzDq6���P�`�D׸�vزI��@�N����ҝv�{����̻ ����'�|���D$���_��k��:f�.o�����{� AkzQ޻�o�W��s�.t}��	�0s!Fb(��`ǽ(��>��@�elCΥ�4��<V(,n���r0���fs�ϕ#��緬QG��j���j���w
Nu^� ,������|�w7��<�q˾��}Zu�\��A]�:Π�R��^�l�]��c��⊾�=�3ËZ'��y��q,L��泸��s�����y��0a���9.r�x�op���3u�.��֝k�+N��k�$����QIy�c�>��O�'��;A�\E� 16n�E1�L�,�Tڼ|ge�>[囓��!�[}N(2��0�1�*��5����k���滕��tr9)r+n����)�Y��j�V7G���oY�����^� d#:�:="����CS��%kʡ�ǊA�!��Aӻ+�2�.�|˺N�,���]G���t���Yw���34JJq���T����g=�ŷP�Ci���Ǡ�R-��j������լ\�(�F���%��ᇼsu���L���� ���c��c�v�Se��
�=���Տ��-�*x#A2s�/׌ǰ��C��J�J���%�F�H�\eB+HZ���4���{��v5���;E^���9����S�t��ξ�@����X���Tì۴�[�o����n]o�T{^0^��La��
�6{x�+�_U����OSU]s�"i���]␛:�֝/Y�dy#�{�=8����&��kvc�t��O{_l�<.b� ���~\��i���pS��ٯ:ܤ��tp<8��z�����UÁas~�H���;S]ק���Od[kʪA �@$�&0�D��@����s��t�-��փJ+4��4��+P�ԶUGMQr�F#�6"0\���U�(����Z�X���2Պ�Z��#h��Z4Vl�%+R�-���L�k-��m��Z�I��YZŭTGV����T-�i���GL+-��Eծ ��D��-J�ҋ(�j�����̳Z5�څm�lE���qUQ��)[V��m-E)h9lr�c.#ec-�D�Q���(��Ŵc���dEm�UMSF�V�4Aj[ci\K��JQ�Pbȥs,\�V*Uh֩mK+TEJ�Z���H��6�e��F�R���A�����J�&R��[��3	Z"Ū��T2cSTl�V������2ڈ[X��5E*
�[Mf."*2bK0����#UX��)e�����֖�f"(�A�QeJ �eZɔ�V�b0�P�0̠��V��-��[G\���_�y�����_��S!� �	��䔾�C����� Vg<�  ;\�� ����3���%z_v�,l�]@^Y�u��#�*@��6O���m߷�Y�Ll�ϛ��� ޞ�� �ݛ��[�]�mw���ˇ)�V`Q4,#�O�q�R���6�`X�+�5��^k���&:�k�n�����AC@���R. �e�$��l�A$�����*��2ϩi��k�4P}2���-�T0 ��4Ս��o�A����՟�7�A'k�� H9u�B��s�Ġ������o�{]��'�t�pJ����*�~��m!n�k��p	[ҁ��[�`;�`�B�&�Q�.�3gM�F�l^uʂ�$�׺�Of��ΏP���^%�������T�ᣮЗ�T��[�_AP8`꽡�&��[YbJ��U�^4�?x'ɡ_1���n�x���MLڠ*���"�I�H�Um� ���B�*�d�/vW E�� �x+��ʈO�}(|�xV�Ǟ�눷�q�N���[]�t��I]���PL��Q���`<�%t"3Dw'|An�n���D�Fk�Q�W�P9[҈?������JixEE"���*0�`ɇ���@|Q*�szP$�w�*����N�O�.�R"��D�W`�n��d��ޔIzA��N����@5�%T Ͻ�@|8<���D$�w'K,��;I=���H/kz�G��
�����Q�z�Q���]v	��0�d$
��ɗ`͝+�I�vQ�0��u5��=ݡ`�����Ad���Y_w���N	P>����$��R��s��١�{f;8�A�K���⧪�-nj�@t�r��&�f{���y��Yp/V��Ƽ߱�w�u�g�^β��B�H�
A��;i�ԝ�g��y��V&{v��O98�>��t�5����m�-��ۍ�Y�]�,Cpv��v�=��=n1�v�@�DB���s�{<��B'n0n��q ���8-�j0n��cGT69{`����T���kv�c{m�Br��'#�Vk�+����:OY�q�:zy ��!�m��vH���c���y�G#�]�:�6�y���v��P:F\�7
Olg�ŝ{`�Y��g�������bSZ֝h�|i蕆��}����R
����i �`V�����8 T�^��;>���<e���7�u��D/~��C�IXS���ڮ}�2���!��+�����Ro�<�{��X�l��P}]��1��QUD �Ͻٴ����k��}������O�t��R��KߪC���].{��-�k\��ė�}ݛN VPd�������A��D�
$�?_��{�ַ�9��<��=�+T�/}�ݛI�
�Y(���>�����L��[� ��͌ !�_����~�����~��H(y͛H<�*Al�~~� )��+,O���7�d�wfV����nw�������U�Q�����Xp���̴�pɫ�k��+���{*K�*����͝u�[��8f{��%@�����D�
Ԃ��~��p- Ґ���}��ïX6����/�|<���[q0b��ج����rh����(u�=�=����܋u�����o��6�Z�װ=O���o�ͧ
��YFJ����gJ�IP�J��~��Ì:°�ۯoo�y�1���wf�~B�Q� �o�w�8%@���7�n%5�i�:�@�V��}�q��ԇ��H+�ǰiP�T��~�V-�'Tia�/!K����1{��Bi��>��b�@P��C��m�=�X�j?M��p �L�_��$���"���9N T�eO���ngY*A@���U��~�D#�~�yD��q�Z5�q�XW{���r0�*%������d�2�Q*o����}<���s@���cX����{��H4�-���}��׬
��9���1�Q� Ȳ>W��P�'r?���M~� ��Y��_?y�vq��*Aa}�?{�u �� =�߶m'}�9�]9�mܾ�1� �o���TN��=Ӣ��5\ǇR���퇰z��HYh}���!w��n�����~!ְ+f{��rN T�e��y���Y�2VVJ�B��~ٴ8�����w�y|��R]������摐!H0������sK�X^{3����$���*�Ke����}��a�����0�|޾�q�$�T��?w�����%R
/~��H,�>�����Ͽp翾� �{���)���ݯ��'m��d%
N92��K�7�ͧ"eJ�gu珻��>�Ͻ���z�� �����܇Xv0�%���l�N!Y++'����U��NN�{�y�8	�h����qִ�u�4�Ĭ5���a���!m�{�|�-�+X矾?}�?����o�w||�!*�S�3�S��畲����;g�`��W��^�����/U�Zk&�J4�j��Z�I�]g���^�
�D
�@���y��é�d�PB���l�IX{��v����n�kp��
�k��k�x����揹}��
Aa���72zʁbT{��p��
����}�k[כ�׻׷�sO]~ �HZ~�~�:�`V�9���1��u�� bpIy��ٴ�@� ������LC��>;��s��V}���:ì+
*J����f�'Y(���u���b���{���X}���>����q�Ɂ��ϫ�.�a��[�ٮsq��h�B)B|dj,_��b@C��[?H,=߾~�|=`Xԅ����f�HZR��_y��
�*w�s������矀��&���ngc%ed�T/}�ݛC�+8�<�M7������
��z�a��$�'�ϯ������?�k���:3��e@�P-��~�%H,
��{���H6����ν�����;����u|,��(z�yd�Y�ֱu�N�K��ͤpd������B���@D|���zws$�n{��~���+
¤�{��vm'*Ad��z�~��D`Aޮ��BfHS1؄"V�ϻ��_�ey�����
CV�����|�-)
�i�<����
�������ìu��y������5�1��T^Rx
t���ɸ<{X�Ŝ�9�CK�#.(��V�o��)���i�}*(���}�1�a��7��gu��V���V|�
!~�ٴ8$�;���G3���h���W{���q�IP�����v3��������k�ܺ��z%@��w�@�Vk����{����-���~�:�ZW��S`���(�#�ɂ�gv�^bT�f�C�'m�k�.��v�l�rZ����8��f�.�Z�'�K��ݛH)�d��w���RO���rH,5�}�͵��O!�&���{�i9� �~�ܜJ�O�����Z4f����Aa��y���z��H{�߳�����o���)e!Z����>� )��@�?w~��q�+(�P|8s�xi�w���͡蒰so���pɪ���W���{*J!RQ
��w��Ì��*A@�N5���|}��~6�Xư+_߿~��p��aHV�Ͼ�8��"��;��%(�q�ɗ�F�}�m;�[�;}���w��8�R�����%B��X�����Ϲ��0�(¤�|��m'6?y�[�~Y?������_}`�u~��Cp�[1؈J�_�϶�+RZ�ϽپR��۔�{��5�
�]ϵ����Y����ì�%e�%B��}B������ʀ�/u����O�y�����,��i��Y9��N��̹}�3'G:�y�T�n$���DVזa�֑,C4׬\&BꢡK�A�>��E�@��9		�S�m��G^�u����:�Q�©�F{uv�^{s�b�[���ٛ�1��=q���M�ƽ���ui���q�v����v��p�8�������l;�cq���c]�ۚ%��qs���8ݡv{N]�5��]�/�: �zk�����qj}m=@;�k�]Ѩ�ݑ�ٞAܸ�vG�ƾy���s����s����8��cp��C��Wm��ͱ���v�oU�m�nK2��Z%F�1�F�m�|�M�C9a7nٺ;����c���\��8��a]��sa�a�(�H,=�=�p�'c*J���l�A`e�������q�x��X|�w���� Ґ�����s���h.��\�䯀d�>�ͤx2Vgw�ww�~��'^f{�Ό�B��X�����Ϲ��¤�/�{�ͤ��d�+'w���tv��͎��o�_}��@�z��2U�xu ����a���P�{�*�|��@�|��n��#�8=�]k�u��}�(�YS����gY+,d�X���~ٴ�Ò�G��)��Da������V���2�zI�B��
�^o�tgY,e@�T/�{�h�Xk�}�>��s���篿���AH,<���p�A|���ض�2浭b�:�Is~��iȁYFJ��_?g�n!���~�<��������%af����a��aRQ/��{�i8!R
A}�<�rpM {��ϼ>�{�G�OZH6ڢ�mȃ2��Zޣm�Pp�����`�˟�a�n��<���N��sFc����V���a���!K@}���7�HT��o�kϹ�:o|��N��}z���s�é�*B���mD��=_<Z9�.[sNnaхw���#Ib'Mk���w�`_��J��'���ύYH`/E�yO�
�X�"x!���)�L�<\x��˄J'P>��{��{�߿z��w�72}R
����@�J��`Q��Ͼ�j�Q�#'���?w��Om�|4�? �+��3sK��Z�N$���6�+,+,+�s�vq�HT�
$�>����}�u�G�}�7�<a�aXQ�Ib_}��ͤ�B�VVJ����������R"ٱ�|	�uo�<OZOW;����@{�l�A�!Z��>����*Q�����ì��;���'�~*���f��JZ==r�n95]:�6�_�g��~a��B��
��w���O��v�}��������;��l��(Ԃ��}��sT��Xy�{��Ǭ
������������G[��l:�k�����DZч��`n��ӳr�=�YmښM��?���o��(�_@�u�6��d�����8ɤ*J��+
w���C�:°��������?C�=K�s�6������?#�����?moɴ��َ� �Xk�9�ñ��!��N���{���׻7�B�HT����߹
Ag"w���ì�%e*�w����x��wf��J��~_|Z9��-��9��»�{͇i%B��Ͻ��u���#�HV߿t��뭫^���O�1�7W�Ҭ�D�����gIc����1��y}�:ƌ���y;�utr��@��|��B�����A`5�c_���w��AH4��y���u�����s/�]4�3������~�P�)��������f�+(�_�ϼ���HX$������C�:0�+
�������OO�������Y(2���y�9H��#J@C��[60�0�~�u|-��5!K@{��6�s;�/~����{�?
Ӽ�<�N T��O�Ͼ�:βVVJ����vm ������޲�mx��ݗ�Dq�[N$!��0HG�Q���G�ۙƳ�A `��)�SrM燆��(7���װ��
��o�Ã$�%B���~�gY�JʐP)}��6��J��}��������0<k���n&� �����ۇ^�+f|���6�2�kZ��@�u��6��
�+6o~�Nw�}7�O]s>��2i
��RV���!Ԃì*J%�����Ad��ɇu��3CXϼz�~���! !�W�h5��ᤂ�?o~�`y�P~�ݛH<��H.�����+����{����o�7$|2T��{�hpIXS���-ϗ-��9��»����5<��߾����
��V׼�g`βQ� �[��ᴂ��X�����*���?3�d/ߞ��ʧ�*� ��ϩ�}�P�9s����C%_e�߰��l��-�%�a[��/W>������k�T��~5Ǐ������?�?�e�}{��a���ye�J&���俀d�ݛO"e+(�_{�_ہP�;�o�o������?ߧ���0�0V�@~���6��
�FVJ���O���ds��|BւI/F�bI���=\;q��v�t���r��mf�\g�J8�����ː�q���{s�Pp�)-�����)JB�������!�����/�W
� ������d���}ٴ8$�,�����Lɣ5u�m������T�B��Ǉ��Y�&��{���O�*J�e��}�	X�
��}�ہ̤!{�>��\5�����˞~�?=���z��f9��r�S�.���6�Y��YY+�~׻82b$�? G�{�?�ߗ�J����������Ęe3��ݛI��ĕ
��3��_nN����6}�=3+��sCf;���3��^?l��y|!/j�ןkߒu�$�0�LK����&�ĕ
�C����uN�b�@d~`�_o����3����V�� �}�3�1C<���hr&�����P-�-$�u~ 3}�+�d1%B��V����u%o7�s��׾Oq
���>�f�i
��RT+���ۇ���*J�a�~����_b�O~�����f�k�s��o^g��C�Aό����:z�'���T.�ކI�ٺ��.��Γ�y7�z=c�Rεc,J��$S�_o$�V���8��d�ё�틒���X�6]YʶҨ�v�ZuR�G�y���`;�'��-����m�8Xi�r����K�=v�y��tD��+Rbg�`
�ڮĚ�a)�������w"s�qY|�����ϋo�[Sh7��^�m8���qW�ȱFw19��wr��𮛠��RA��&�����fUvb���9�Hr��Ǟ:�{ކ*�x�g��At{�!�N�W��fG�kn�c�.�W7���.ɇ81L�H��]�,��)�6�5���z� �2��bo�v%Ʈ𦫤�'�w�\x3�{�D�&v×:Cb)[����!��Śr7

���.l�����{l�*/&�>�W	P%�~�IDAk������UR9���&��F�Jڛ\{+v�'+3�S{G1ssn�B�і���=�w���>�Ҋ�'^<�|�7���qm�or�:�"U%����-_^,�9��'´�ye�n3��ǜ��G�D��p ��㻾}%�����iP��J��睜`��x ��-��)yj��n�p�G�	ܔ{��9�Eƴ�{q��O��{�[;Ru��z�cǧ�z�:��.��$�v�+.�=�c�w�Tkr�.1ˢ[k��=�0�BϘPL��V��۪�̞�X��m��M��/���mZ'B�5�P�{Ke`��)��$�� ���ADV���[kS�E��%�JZ�����R�V�Z�"ԫiT��V��dQ"V"����r��)h��j�ihҍ��Q(��G32��mX���6b�i�̵�1���s+��b�-�s�T����Z�0*�2��R��
���SIADq*	R��!KT�ZZإk�X9L).�G-(��Fٌ�rT��KTW3c-��5�U����2�Zbe,�R+XڨU[(�(�inS1X��Z�iul�Z5*��*WT���D��ikc2�[iEE*��K)V�کU*��LqU�Sr��aKC�Dʫ`�ʢ[CIf:�c�JQ��,�Z�2�J��,V�V�-���Y�]U�e�,V��mj�j�ԴZ�*9f8֪���F[[�r�Q��jWL�q�������E���m4����+Df�����6�(Ĵ��Q-�t�U2��U��!YZ����EL̹U�Li�����ZڢZ+s1Y���j
��#�I]i�Pm(�nYU�R�(��k+L��.%{�cc�o����B]�9�mr���4SY��t�Cs��Kf7Kf5q �[�i6.8�x]���صc��.�b}K��z�
Ʊ��Ӷ걜N�=3x�n�Hdz����<s��C��[�ˮ<:$�2��1�[b���g�/B�V��z-�A��xMԕ�q�'<p�ƹ#l�qۣ9��.H[Wg�u��uh��7���1v���[�67�$��0m<���$zwq2:�'nrr��J{7mt]x��g]k�۴��N�1��#����7l��F�U�v�S�A���=��<P75C����$��=r���]��Q��9���3���M۶�B[�b���p!��eSv��e'���`:��퍞�q�;3ֵ�\=n������� $�7e��=��;нyK�t���ݹ��/s�@uȣ:��v� @�w=���n���\3�C��)���d��b��/�� :�5�>�m��c�t��Sc�����s ����"v1��sm�m�Ni�.[�X�#;.�.V��pgs�i˹�Ϸ	�x����+u�TG��㇞'�� S���d{;k�Ħr�-S�dyl�V,s�mn�l��x7Z����K\��y���ɷ!��� �.��*'@"��73�9�9�9��`D��M�la�Gr��j�vN�t��ׂ�U�v��݈�]�Ӽ��]3��f�=6�<Q���{a]֎N�+klۺʂ$+m=����vϲ�=���:#���ۗ۱f�����޵�uԭkn�#m3!ˏ;�v��랠K��J��׉^��Cs�����yS�N=�j�Kx[69^sm�g��i������8���{t\݇�n���:ׁ\s�n���ǎضG���8��E��ۧ<;��}ԵIu&�v���h�ٰm���p䮶�wGkl��̝����[wcBh��gd77�{i�,��U\ۻd��LX�p����7\�D�ݹu�uكv��v].��v.t���Lt�ǰS9��)���fdծ��\���.��wwwv����V�݌X#�ظqІ"�b�v���tsn�H�k���F�Ň۝=�Ӟ`d훳��{ۘ�x�]���f+mc��{]Y�����f��u9�+������Y瘼��퍼Z{����[�5����\0�e���۷,���ژ8;v�un۸:ۚ�d����=�/�����Q��ۚ�6}wc7o�9ں��7f��3q����nv���n6k�H���'h�{0�zz�Y��p�����g�3�ι�_ﻈi?���s͛N!�1��C��1��y���4�bb�	�c�w��s�<a�8�0���>[w���}��!��2����6����+�Ę�1�������m&&���q�hLњ�cé6�!������������ OT5{])=��u.��l�e&�ĕ
��ǿg��!��
��1��w��o�<g���3b�0��c�f���xm5�}�
 ~"���7�hB�b◄0�c�y��c�6���2C{�}���&8Ę�������.߾Ϗ3���i4�DĘ�IY�=�<�p�IP����e�������8 ���(��q�ҿ� a"�P�3���������q������1��c���͝gP�&!�`��0�����<C�8�$�T�/���6�z��~~ٳ=�">DG������_#Ğ��|E���3�G�@G�*��u���Lf8��*_��vo���������8��~��� ~8~��Sί��4��10C�b~���o�<g���3�b&&{�{�hpM��/�����u*�����1��Q��} o��>��b;
���rĞ�h��s�sV'����}������Hz�����{�q$�T�2�0�Ͽ{��3Ę�1&&	�12g���I��bLc��{�xcu��������y��Èy�LB�I�c<����|~�������*2�'%�0��@d?��� #�����z��%�2#�/N�\����w��"9��찆H��5�m�d3�o_�����|����[�4�=���w���~���>��~C��^���4�	�b��0�Ͽo�u��!�0qI�)����6�����g�G��uk<x�(����O�����N}���sZ5�����M�X}��?o��|I�T�2���{�|
M��Rb�a�c�~y��}���~CT*~C�`�y������C�1C=Ͻٴ8&��]l��hD���◄?�@fv��7_��Xg{�����?����{���RW���bf~׾��M'c0q&!_}�_nC��=���￉�_ғ�,;��<߈x��_4k�������\��T:���}�ͧ����b�f!�߼׻;�4��ו�i��������?}�<Cĕ
��ę��s�vm't1%pf$�{�?W��ψ�|�\3<5A��j���:���a��cͩ��S�];`�ts�/�$�n�=g�OH��1C���X-%	��G�G����~ߌ��&3#�1&Rb_}׻7�I�1%B�1}��}�qIP�۞��5��9�����|����C��1%K���f��M!�3��/+W0�շg4�Xtq~�u�Èa"#���~=�q�J��Xx��>�*J���3�w����bLB��W�|�ۇ�1
��|׿�e|<�Y��mq��� 3��/�E��0=\ַ!����5ݛI�Vr3�c1|��}�qC��b��0g�~�/��'�_�>zո�e���c�=����'t6��/twc��w����]���N��I\�ř\��������`��UAMLZe��~�W�8��}���o|���?0�qa��bL�L��{�i9����1��}���C�q%M�����q�f�����n��W��3�_N>���A���#�"h|�]s�o��C2��b�y�p�N�b��Y�y�}�񌓼�|���|��&������J��h���9nfe��ư��}���!m!m����Y����������}d}�0�G̙���ᴘ�IY�Ę�q���jC��LB�I�c;�o�u�!�����߽e��)�?gšf2�3� H�U%�q�
Gg��\���̝a�у&�\��߿߽�prg��2�
��*]{��m%B��b�f!�߼�GY�:�	�b��0��|��x��*��{����7����I�S9����NeI\bLq����u��>DX�m�Q����#�#�!��vw���RVx�LCX��믴o��8�w{7�LC2�ĕ
���{�u�P�10C�dO����3�b̌d@�ϵ�~�~�Æޭ�@������Z(��b;�?��y�C�*'r�0��}���RW���Ę��g6����m%O1&3I����{���;�LB��1��<����1|��Ja������!"~��D>�l_�Ꝡ2#�@D�
��y��C�bb��Xa��~��!�#�c��bL2��of�!�[X���*���U'�?H煫��i8//=���NV��k_��=k']�̅M�焼kU뽪�~^�^�fǶ��t����NlG�����z/��}�_%ĺ��bLpf?y���é�4�;����Й��ǇRm:������~!ԕ�Gbe&%�����J��?y��s3��}��I�T+Ͽ~�܇P���&!�c0O|���3�b��bJ����Q�!��w��߽����Y��̌�٠<�.���n�m�y�A�Q�y�\�N@X{�=�6�h���?�@��� c�?}��G�bL��3(c�y�����c�1&&&$���߹�i*pL#�~������׼G�~��V���a*���e��y���b����ѦWk5��p�q;��y��m8�!��b��}<��N�u>��w�q
�Sĕ
��<��x��<qa��bL2��of�T*J�I^w��ZQ�����~�U|<F�C#�C��d�r��4\u�4��V���}g����*e&%��w�|)1IP�F���}��ów�+'� 2&!�c2'�<���C�x�C��C�13�~�͡�1a�~�^V�a��l�p��ဲ5�2��Y���]n(�}˨����@2>D~������c�1&&&$ľ~�{6��Ę�q&!_}���8��0���ޓh^Rb����~!����'�޹�S4���\ֹ���&s��fӂ�3�bJ�}�߷��gP�>ז��������?}����&!�3�����y�CfS<����NeI\�1`����_ ">Dܻo�]�h�c�+�
B�/��5~�0��q��/k�!{��;y{�:%��K������j}�<�t뜦�Z?��������\s�.՘�<��Ŏ��t��;��}�u��<c��oj�Ƨ���ٺ��Z��ݛ���x��S�-ۖ�Gn:�
�.��p<�<hӉ=��q�:�;��e̊k;��z;n�n�Է7�$\X�oV��S��F����م{w[��A��'mN;(g�mTvu]�z�Hqev��g���:��s';U�svn �x�e�Aɮ�V���ۀ,��������벃ڰtW^�Ma��[��5�f�Ts�ěO��w�}ߌ�|I��b%K�of���e&!�C����rB�P�1{��EV��'�8�`��ί<GȁY�f!�`����w�hq1a��<ߛj$c�9������@q�"a�1'�>�����u�o�u%B���bd�=��6��c28�������C�Rb
LC5���� �|:J�^ x����
�$q�]¡��L��ofӈb�f!�*�����uC�1LC3�{��پ}�}�� #��,��a��=�{6��RW�Ę��}��op�tLI�����w1��Y�0�p�N�bc�����o�w�t��*J�IR����|���e&!�1~��p�:!�bb�3�����O��k����b3��1%K����IP�,V�V���$َ����]��I�C`ea�}���x�{2�������G�F�C#�C~��b���Ę�q&3}����u��+TG��~��U1�b�ƾ@����~P🳾��3�B�w=u�p���טU7n��zx^M�ƼrƵ�]��Cy��"d�NO� D�C9�w�i�1IP�*��u�γ�iĕ
�?y�s�<a�,����~��̬�4����ߪ���Pĕ��I�W�{�w'SI13��,��5!5c����vo��|G���d|���R�r�����h^f���:�������WfL�yʉM)���/�٧�k��C��&?9��c��7��׻�{�Ē@7�N������Rb���8��>�������b�!�c1?y����C�x3�`�C���|>�ϯ��}�of�T+K�����EB#��,����@p8@�L2�$�(c�y����<I�3b!��#'v���|������2>hT���������1%B��V��V0�?@e���@��R4���@d>��B��a����xO����f!�*�?k�γ�i��bJ�a�y���<a�bJ�IR���ٴ�믝{�x�<$�FbLB�{�_nN��LL���{��Q�ˣ^I�+{�}���|I��q&!�Rb_>�{h|�N�P�����@�g�����_�P���&b�O<�����1f3�113�~�ͤ�V����3��m{]��Y�ǾD0̂!E�"k%:r�,vۃv6�j8�h�2)v��?7��`E��Y�Y�����w]�t����1&C{����Fx��111&&g���IS��1�~�^��߽�=�N���}��:�$�^�b�y�o�<|�1_;��Uև�����4��bg>��m%B���1�^��}��"���o_l�3�iLCȘ�0ϼ����x��CfS<����J@D|�����?�=��'�}�ߟu|=O�m&&K���k˭&\�:�hV�����=��1�8�̤ľ{��o���aI�c�C��5��ֽ���p��շ�:��n���]\ܮ�N��'#�o���ұ:��6���Z���MK�=��[��ʅ�ϱ����f�߰�!�w^C�i?��&!�c|���:�#1IP�bbg��of��b�/<��esMi�\ֵΡ�Co?}���i��o�CT*J�a�y�����$�bLL�bLL3�~����Ę�q&3}���èk?w.���������/)1���>���Cĕ
}�ܐ(�JH��� a"W�D�b��c1��>_��Ό�C����C�y�=��>�x���1�!�*_=�{6��CT*J_��uv~��(���۵��������9��@T���W;�m�a����(�,�gic[���P�IAug�����G�O�o�w��g��Lf8�ɔ��Ͻ����1%B�0�1���~�:���}=�Q���@���#�gmy�1f3�2&&y�ٴ�
Ó�/+n[��35��a��1����u�I�CZ{|�~���>��=a��y�}|g�1
��&$����y�i*%B��W���nC��&!r�|�c�Y�ʣ|wO|��V@��~��^���L��r_��C��Tm%B���1%B����gFu!�d@��?~��{S^�r����=IP�=CfS<����NeI\f$�c��߷�S�12���L��������߻-�/���C��u���G�m�  ���w� %���ʞ{r�¦ee��hy޷E{r?��9Z ���<���6-�o��TW_�3�.oikE-�c-k�]:���Y��p�~��N�ד�w��%�_|�����h����(��]X	q�uK	$��^,2o{�v���~z�P
�ÔX$�������,��ޥ�{5��Fі�k���fl��������\�i7Kn�����HdEQ���WGH �ȭ�WG�/VwfbAsr�)���8��_��H �T������ڕ�كK���Z�`�=����� ��n� z�{3 �;Պ�|�{�ۈ�� ��(�3.f��q]v��������Fg�˻�r� $p��_i�55�Ϳ�!�+�@����a+�A�OFt��b&��B ��ّ��oIr��s�Тo!�$���!|
�0Ar�U-w��,�I$szB]=�<p��c�_��E�Y�w�������V������aV��n�Od&�wQ�W�9DZ�W�K��B��R�nԎ��Y��+���~�v�Ԩ��W`i����u��7| ������AH�d1�#��^�.�:��=s��t=��;nN�^q��i�Z��.��v�u�s��b�7Q�=��\r��%m��n鬭���Y��x5�N�g�Jp+��u+��L]Ƭ�v���
�u�%��m��͔颬8pE�v˝�Ss��3m��h6Y-��N�xq=����r��ܠ����G�r�m�Sgg�v���9�;�0�*�;svn��Uۈ��h:�p<��+Da���/JF�Ӷ��u�k���B��7�K�p����.={wD���o]�$@,ިI�}\��NvI�C���D uf�f �W��"f$c���{}� �����}m��@�T�� egvf  A�����{��Q��{�4����$&�F6Ap��Ysk����� �b�bs�^�uk��ά��ĉIf����"�i�j4�vE�����ޤ������v&y����"7i�  G�޻��낡�[� >�V{3 Q�pq	����m����h��<�XYҗ��r�����t f�t �Q�v�t��e��B��q�u�t�S\[�]��:@�c��G�`������wqr����1�3�ۙ����) �w�m��Ƶ~ו�������F]j�nL���3K��õ�I}W1��ۺ%wܰ_�R�G텹��I�-鷇���V�F��(�N���f�5�혹��
Ꮖ�_h{[yս���v��������j���%��Dw�q@ �]��r��Oe���)��\��$c��A���� ��j�����^�̐�_{� g��A��vJq�jJ4�FLR˞��WS9������"#���� @>��� �_v`�w���ԉ������H6��3vF��l@/�j�n��g�U�Q��F� I9��~��٘����!~)����h�Y��uq��.̜/E�v3�ٳ��6�M=Y����7G|���L�D庞�n�Oj����&j�6��-W;���s� '6�" ��i�W �@�D�p�e�z?s2��у�g��l�3�I��H ���1 �ȭ�X{.��$��>��JFB�lI�'5V�|�޼�%~��O��T�9&��ȝ\x3ܥe��d׬i��=���}iw�,�)g�z6��z,B�ݑ:ť^�z
��71Y�:ܕ�{7��<]�mW�܃�(�t�^�:���P���n]`⳥��.6�=s,7�m�@�c���&�"ZX�%�7�[]��Wt��]�f���I�
�K�ⅵW}��agˮ�z_�=���u�B��8�N����(q��\�i	�
9F�����'|�s=��H�Jg�nr\>�7}_���B ��Gl�G�Nw=2u]�2.��/u�9[�z�fd�_&,͝W�z'���pL����b{�k�Ox<z�7y湍_-��'�[��i����Z"�<�U����[�^�w���w�1��0�e嶆��#�;ι���\劀�}���smub�
���#后)L�`k&Ζk�v�Ѿ��;��/����:B����%� �=��<J��<ʻ���`���Km����+�k���:7��y҂�V�B&� �n�Wn�Souz�8)�~
�W��F�q��:ݢ���ۻS;�gqM۝ohnWxEj���B3D�{l�`�����M�۬:��: h�jE��zs�Z	�ŋ�:q���93i��p�l	@��ښ�l�w����M�V���=�U���h�%Sկ�Z{2��`���V�?u���t9@e��w��Y�H[���V���c�Z'�1�eT�Θ��7Q��VW#�ɻ��	�o��e����mmΛ���j�A<o����V(	��R%"�Q�ukS-�*c*�U�Te-[l�)V7�s0-��©F�\p2Ю5ilKR��kY�����MZ(�Xj�8��J�K+kR��Z.e�.j��Tt�Zت"*e�Ri����EAm(����Q�U�ժV\�J�)W`�c��q�p2�W-a�PQ�̸�ը�rʂ��s1pim*�R�Z([EU�ZҖ,KkR�����V�m��QTUʲ���Q�2Ҹ%nQ�*�F�,9s%UUƩ�mEV�KJԪ�9���ֲڊ")R���̮B��c�D��J�� ����u�PB�,X1YKb��+�DcL���Q�)-�ФX�mEFT�-
����Z�F
*5���D�Ub�h�V�čh�DV�Dm��Ѷ�EQUkD)ib1AcTX֤E�\���h�"�XYQ�J�ijҤF%��0WY�V���F�" �`��)��bm2�����"�e��5�$�s|��~-�u�붊IWg��q�<5"���Cv�k�R��q����|U=j� @u{73  ���J��<���b ޷�4�Q�Dh�BP��R�ݘ0>gkt�{�G��{�LC���� K�s��"PK7�%�}��}�d�kZM#�h�gE�s��y؞E9����h�����q$*1{�5�Qm�j�{�*�wb�@ ���ϰ H��qH9a�~��<����S뿚$�vu�$�7���
je�n��
�n"�i�kQ�y4�=r ^ͻ��7����߭�r}=xZ��d�����,f
��b=:sİ#}��@$q=����ל��@z�72#����V� Ƣ,�R��}Ѝ�/7�kI�n�A�H�f 6�5G__�����>ɂ�*�4'3��i�2�1۩zs��F�qg+����OG��PDP��O�u�k����^��C��-K�r���_�� �����{7?f`I��Ȅ',Q2����{��H Vt�*�]��*	^'���z%%��($IAe�붲z�ÈwoC\`-��I�S�VV�`g�g��ז�4�,1,م�C_DI� �>��a.5w�uYٟ`|A�n�OĀ~k�ȁ�Y=�붽����]�w�/�'��)%�a��)6�5q;������S���z�Ӣ9���d� ��� ����"!M��)�Q�s�罝�$�8�B�l�TR]:�'>I%���"S�+��U�[�.z� H�;[� �����C���L�"i�9���\.�59�ao� F��� ���X z�ݙ4�>��P�f�{�����X!Č��Lc���޹�V���<�Wһ�8΃��^�ՠw@ͧz�v�Iz�ݙ���S���N�zv�$�틈�v*J����/�ʊ��q��+�v�hNn�z؏s��޻�vc��a��'<�#s�0{,C]�랩{�|����q RF�Cr
p�y�v�+ֺe@��;��ӝ�v�z![��7�u�:c�m�s����Yډ�����\vy���m�m;y��[BS�C��\�c=���E���B���ݕ���$�x�Ok��{^�]F��nr�:w\\9�m!ڀ}[6���k��uʼr��'�Y6�p�u�ʳ��QX��^9v��sݭ�.��S��^��#tw^����㫥
�<���ݺ6������i�Z�t`���F��\��2�� ��t�WN��� �]��������#>�n	���=�ni��(��%�]�U��;�e�WUuM�U��| uz}E���vf|�	
Y��{�Bq��@>@�����f�>���a =�~��xSv��\p #���䈃վ���$�8xB�bF�2]XJ����"������v�Hl��^��g� �7���G��̧OȊH_+�Y?:����ee���Q����$ ��n�-�h�}f�zw~@,�~�Q&�?=��d�@}��&�O��X�-����_�3lЯa��_<�v`ץ�Eص���Q,;wU�t-�M�X~�ӨZ���QOW��=w'���u�� oS�:��n/�{��a��[[�'bxjD �)���%��RH%�C�ϥ���3��կr���'�����l=[2^�)���Q�4�'��R ���|o�"&R��H}�s+mr'`j�<��_Io�����b�i�������[K{����	u^93{K�2���Or���&a�5uhu[٘ gkt��w��ah�^��""1�u� ޒ�Ja��)>e ۊY..����컗<�#�h���R'�@%>��$�pNݛ�^;l{:�gĬ�$�@���-�$m�%Մ�nJ	$����䲟q����Ѱ|Hݙ�H 2�뿙�_�yUo���d��vz�����Y�n-�����kaG���k���Ln��S4"0��p]����"No7H  YS�s�o�"iEgo�������'D�Bh^�@�с�b����W�����N|3�bK�"�y(�Ԁ3�N(2���m��gս�w�����1����6�i������ ��vڶ$ C��};e�d�g]Z�o	%��N�~ݾu���㆖��dJ���Vl{ɆUF��<n�ܺ_j��ӑ�e��w�f9�������;w� �>�n�	F��`�yR�B��
P�ڪ��4U�냻����)�*{no����}p?��]0{������<�s,wi�n��C���ŷ���8�`|<�q�Q$�T}��`"rt�L�J%�rU]1%��d��!�BJ-�0������o^,��I��p���������~���ߝg�����r�n� �h�]���}�q�U{ϞTTGv�K�t �3�l��P�Y�;��s�3)V�F�ݽ�}N%��� DS�����'C�@����g� opZ���;�z���o^, >	��x���u'��� ��gl��ٽw� �����#Lݥ�}qV*����n�@|��̈��y�0< s�{�{{�����>��;��ׂ���G9�wu���1�n0��5.��C�N���9mw7�f�U�ι�g� Hy�~/��=�V�߮��Kf�1K�U��,�I#|�W�QyW:��Or#Pw�6����̈������7��7���m1�"�A
q$v۳<ܘ��\�Tn?�rn�{� mTB;m�WG}�����A��	&Y5���հ"���` ���=��-�-�#n.�}vD�3=ل�9��#�bGui_;�&V]� )�ZX\�Yw��m��?=~��% �6yԐv�V�^μS�$�[�XB��1�۳���� ���JAAauW�3�(�/}]�7�x"����@ >��_H(��c�L�D��-��={��C^ұY G=��2 �Fvӈ���o^D�����/�J]�fbK��h<QI��b$��[]!4� �;m[�7|���w��@+�{3"3�>�n�A���l��d�i�'�U�����{`���-E&7ʭ ~�嶝�p,�{����sF��awbՍ���� ����נ��|3�^��|`W�d �_��3�t��Z��v���+�pG���b�\���aR�
u=macz9�7��'i�{ �a��N�k[����:xm��n�գ��pKgqnn-��q��u����'�[��:h�Dm�{d�F�M�ۙ�e���N������'We^;��:i`y��<m��v�r�:�fc>��\m���;�mЅ�`C��*�Ǜ�t�StD�T���vCa��.�ZSv��X����p��?�����I!�5~�����A�� Q�Saq:�y��[��yw��� >�3���8Ϡ���&I7hwl�-Wf'��ي׽x����q@ z�뿙��e���>�ȅV����Sc���p^�t��	���_�K�K��n�y�D�H���3f΅C��Y��ܭ��e�k���'&�) ��)_yZ�@���j>���ߝ���u�}b�(6bib�V��_X� �՛ט>������6"N�l�ē�X *��́WB�/w�;��Ω�����l#������0��&�����g��v�0���%I$����t(��m1f�'�Τ A�nڶ z�����/�r�.i��㯤�,�`���G31P�v:��ŀ�y��jn��B��kQ�|����,�����u�5x �<��W�ǵ�C���牧���t���R�Ќ�\i���VF�{�J�O�$�K�S����,������g�٘���zj|�u��O�� �/8��e�BS��Fݥl���� H7�����3��|�w��M�/�3 I�o���Ċ1�Du�83\l������l�f_nf@�}͗<��FZ�~�݆�9��"@<D2�	Bc�k�۹���$��� ���&��ch�빰2���3�>�7_ ~��a9w�4�{q�B�N�&rW��g���7g�Zsss��,�ԅ��ۥ��j&��)u�.�{S`|�޼�@ o��Do�Wru�{j�/�� ��Yݙ�|J�(Z �$Ja1v��7@$#ʷH�Ϲ���~䭈�]Y��� }��ȐI�����U��Bdr������\J���;��[}���A�n"�I�q��յ��#�˶��pn�:�w�R������Y�IȺkLAZ�cv��7.�\�AS~��/��м�7n��ެ�v���|��$�/�?�՟��I��!:(xL�sMH�LF�Ҕu�ȹ��o��~���;�X6� �`]��~V�>��n�4�����)���ۦ�A�~�T��g۹�ld��l�� ���H!$�oz�R��%�e���>e�g";����3�k���0u�c����B��@�w��Y�Y0�&<���ۖp$�#}��"�����7-�j�3.wj�/�~���	N����ͻ*4�Q4�8qh&��i�Wk{p�Ba{<��2h� �{i�| ����5��oثϻ}�Ur��������=�� �}�uNw_m\�����R ����@�G������V���K�C�í��^��Q�F{}��@ ��7H"����� �of[]u�vuŘa!���6#N�����3ǝ��T6���gd�c�"��X:�i߈r/M%&k7�RY1U��O�� ��| w�n��K����&bXI)��@�WT$�w�oF+w��l~{��t��M$un��$�"�W�@y&H�.��{1zz�����)�!�ce� l"�;�W��f�ݷo2v��䎭H۳�7G}�~m��xu�)��w��m�� �ؿm�� �7����"�,��+�&�fi E�=w�$��"�p��2\���ۙ�$b�k��:y�A ��z�����55���=���[�R�b����6H�p�u��v�  �f�� �:\ɝՐ�� ��u�m$=Y���"�� u�M1��{�[B�q�~�l ��$��� �4OOfTꚼ�Rk�eh���%U����ޡg	�%�Ysk��(${�!5|)�{��^�o�m۴k;s3�Do��B�e�2˵�ʝ�ϭ�y$�y��2�aNyF�hϷu#ٽs^�Xu��ܽx�c�{s�{I�Qab�ʊ����PK���f�wH%���I���=�1��7o��{;˔Pb�:ĻJ;6�!m�7��"�3!%"�����ʁ<��DY�B)��Lgc8�깴,T�j�������\�@�ܜ��7�:�g��gϩ��ڙ�����7��9S��ų:e{d�յ���= Y�7)��Cd�ȠF��s�������y.d����2���h���
�囙P�-y�Q
:�#��}���]���E���s����V�;�yvqӮ����}������M�J$�w������I{|��ތj� U<1i�U4*�yf�������ݡ��y��&�;�H�r�<V{]�g��Q���?l�>��OhB���:��!]m`d%7;{��x��2@F釚��W���b���Zj_���G�aZzy�{��KM��
��g��R���.�Z-��wma��tm�ܻ_r�j|�^v3�K.���OOw����^cs�2-l�ݖQ��췒�M*�����Ʋ�U�#��a|˺I�Ŏ����g��&�Of�3��5bN�-�@���SM�����84b���]�%%/5����e�������^CV��ߌ!	g�@��rw,��/Aӭd��j���[W��sV9�=��7��b�\@S`�i
��b��7���P��DU(����Z�m��U�H�FUE��65��J1��jJ���(�E��VհTQX�kU�j*��Ib�b�ҵih�����`��Kus-V����Bҵ��ڋm*�E����APPh��j-�������Aj�iU���DQ)j+�����:"�6�ĭF֕�QB�)[���&Dq*�Z����l��b
�DQV�mkelkV+Yc[E�mZ��[�*(҅KlH�[QJ-�R��J�4n�qmFS�(���J։m��4e�V�mm*�˙j�0m�Q*���+R��Q�X��q��R��T*�����=����������ZZUQFT*Q+Ej�"5t��V��ܸ�+eR��)F�L0��j�P���c��m�KR�PJѬA��+[QJ�r�6խ��*ZY[ZPU���1cS�0{n����mW�v���nx�M�����)���z���:�|7l*n�>٩�rw0{Z���<�\�.�q�7,:ӂ�T�f#���*�V�R{v�䡱�;�;
�d��\�qq�K�9��t7&��u6�n2<�ۡ2X`�S6��5]. ;g>z�֌��Mx������9m��n��1����ʳyy�]�s���.爍kG`��uv6�vr'a���n�In,���2��h��.װ��k=\�p8N[=��U���e�̢=˼�6������M��fݞ�@&{sn�b�h��vm]����ט��0֡�����:���Iϕ�n��u�R��+ًv�{u�M ���a��^<�m�h����Cv����7l���`�E���s��:W�7/3%�N�\Xk&d����⧃���s<���6�]V�2�e�n'�{��:�sl\t�0�L�u�W 6v�q�㮡�\��p�s�\��/n�w|��]��m�j��{Wv����N�NMvaw��+v��ɛ��)M��էu��`t)��Y(�4n�"�v]�(T���ͼ:�1\�kFv�������%m����b���qٶ��^{v�`!6˞���c�$Get��<��xN�Ն�/�|��p�Ev�s{�e�ͮ`Ӌ3�I���w�����h�&ݝ�v�Mt�,�v~\�����-VK�v۔6�	R6�������YG��\�yx����۞70&Ѳ�\�7��.A	�u[��:�^���7%��]��5��rݭnl�#�
��oS��ol�� V�n��;^���"+�tgQ�ݍB���.W7d��Λ���N�L6@�&#�&[<�^Ɠ�<v��$d��Ѫ%԰�u�r�|�ӷ�{[3�s��$��njύh:�n5��^�۞��=Uk��s<�`�0@�ۮ�Ƴ)��8��8��)����@q�eF�'�=q<�qώ��unb���!�����ֈ8�Z��]�v�g��<R�T9�c�cv�{����|z3�>]
�kΝ�gc=E�q�ێ;����K�"�<7k����<�1	�4s�oOYku�'�`�ۆ�@j1�;f��CfB�V
�x{6�����ű*�p�^;��[����Cq��F����x����^�V��� �h�scgx��xm��/gok��E˝nѶ��- �����y�.6�p\g/͸�5�7fc��#ؓb�X͸��z�npX2��sGh�nȯ=��QQ��ѣ��/�l��LF��e����F�v�,�#}��@��:�9u�u�\&�Ck7�1%��<��-C#��K�ܦ�O�}��x�ʚ��,��]� �y��s�7Qy���ڃspR@ޣL�,�
%�޽��Ԑ	��A�I�5}���^Uv�	 ��f�f ���ͫC�I!�����TD�ȫ��� �g���Iy�D�G����΃����:�L��-%�ݙ���	Мi�"P֥5��� �w[�sY����巙ّ���� �E�]����'�?|v�~s�λ��};o6Ӭv�.E�uፉS<ط*PYi&4�{O��E���/�e�b�����2 �����`���ߧ��,���{31  H8��`�xL��m�[LF��J�t�V�{W��z����b )SeovjJ�X���_�$֌�ݡ�X�7:].���o���̄`TR��u�G��wZ��u��'�$U�����Fg^u�XD >�1߷ TO�T.�����2���D��8��K�F#wD꺘"%%�����wF����� Aǵ� �z/z�z�2p2$(L�-o��5f.��V��������  ���[�>�޻����ux�j�� I|�*7��s2H�p�uh:=}j�@�o^a:�f�a�{�I�ŗ� At�k#�6ɮm��{vc��?U���6�M����Ӥ]�t�m�E+��ָ�g����ލDB�K�ILo/���L��� ��ݙ���z�y fy��M�ݫ��v�.\!(R��Z���dr��>x����I4���D���y�5��� �Yي��z���T�8�%9��+n�ЀAu��� �.=5닃��uuS����պ�r�����Di%��ڷ~l�x�:k���TW�^��R��ɪ��D����{�So������5�z?�/�<o�U�H��׻�f|��k��%�#��K�[r㳣;s@\om;uݹ� 4�o��==���g��߀����qY�i��� a$�j��r��:��+�$�w2�cn��q����]n�� � 4�t�����p�z�!�g̕/�I݇�7;�v<�,�2e���ۇ�]�s�<�a������eƒ�E=\�_X�%%u��π �|�A�T���9c^�Q~��D����f`I'��4'i��	���m���7�j�~e1�JZh"y~�Ȍ��$ T욅���W���E/W��%�%�Q�U��L�I#��7� `�ܕ���g�W������#���5e���sO��rݡ��x( uD����&�(q�( ���R덇� �'}ؽW�x����(��`���5�Y%s�[�e��V���9�b6Ě'��U��PU�h�����}}���gcج����~����~���~��V��(ȑCcm9��ɶE�m��v���Z�՝[ٛ��� ruԑ|m��Ϝ�fK���UtTZ>�H��*%0#1@X�cv4��:�q�:(���HC��4�c=�����`a�$�ʻݹ�bIwJ��PIm�u���q���j�tg��3>  ܝt�>��dL̩� ��uh7���g/�лV���N�/0�c�Pz׺�$�-��|E�����@I'G~_p%�$�.���J@�,ݻ`5u���'���� d󯤁 >=g��E��Ip��@��a9��l�]��v�����ǲ /�^�ι���ٝ��S�^�r"I��	�+��<XjG$ħ3v��V����q�8��f�v{q��}N+� 6�똋@}�~�̢W޲*��r���]8˙#7o����o}�U,��p�G|��p&2��[NY���0�([�}���CC�yb�8E뛾�g����Zh2�CFzGvت�]��<�s�X<�M��уT����M���)ۺ�8�7�I0���ۋ����,�<�C��;"��9t��n;j�����Ą׎v۬x��5۶�7�ۻMM�s����7g��0��|ݴu(�q���Y�n��wN�d���n����v��V�n6]�l烗F��x�vm��4γ�-��ͳe�������vʔ	=]e]��mzt��B�k���/%�;�}�-�pF����? �)-���D�MNSͺ�Z�p[M��ـ�>2���Έ��	b�*SM۳{}��AJu�b�=.k~@ ����+Q&���l�D��e���h����� ��6@11�Xo��V�9O'L�OĿ��1�X�@]�� �v[$�K�$��>_x'-��7a)�s/8B���C>$���T��I�O�Nm�h�:{0��}�x�M�M��'qg���kMq.\ �R�I[ٟbI�n�7��^w�ߴk1 =s�s ��}~��@F��������Js�.z�-�����l�X���=i��]�ς`�Ǳ|ӷS��n��	�D=���8��Q�X���.�q�������$S���z�{ov}d"��$�`/ !�B��V\�ZA�m��{�+�E��:��R��K;�A�Ƌe��}���`[	��R�&��Nw1l�咎����z}{�s�X������~W"~�u�F �}��w'�f���m>��՟YN �A%C����̟���#�� I��Z먔�����@ 7�ݙ� �7@}�ՐL� ����\�~�o�l��c�p	{{/ w��P #/�ב���O>��b_w�3�!j%�)����y�@�e������Qg.����d�O���f�H?KR�!��^n�{p}�pE,;�"I$&��J�������^��U��3ۛ�$�C����?v�A.y�n�٘D�n� ��yDޛ���++��{m�~$	=�}XL�ņ��2�n�)Z����T��y�蚺���0 ���+ &ͻ��X�g��~��^ B����n� ܶ�(~��r �u����*��&_���WTuoO��>i�<�:��vaq�
y��Fi� o���R�N=�+.���^�z�����Q�TO����QQf�q�{�}G��$����g�H����A�~��m/�i5���@�\���ۂ�#ƹ�QT���pD�7I ���e�A��ve���Rk~����g��&e&;��?N�Ȁn{��TG� _y����&��}�I���}�o����G��bJi�n�	��a�7WU���%�g�1˶�8*��3�ϯ߳q��K&�/���@�;\�=�<�&�r�ǋg��>[O�{�1Q �R
���4��v�,B� �R�)+{.0<\W,�ݜ����v�|�sX�4I��y�D��|� ��gQHV�<<�-��lD��S��"m-���ɢMQ-�iZ�oo��` �W4��^��fg�}���%29 ��X	v[e�;��љmm�� ���r}�$��9ͲI t�f��/�V�e3�Z�q�$3�Ël�o:yw�oe���Y,�Cܹ��)���q�A������4&G4��W��٠N	���>�|����[HZ�7j2�@�M۳o�3 ���uܺ���mD������/-����Ā@|�l�X+�����BB$�.�NV��^��aLϙ�^z�ձ����Og�%go����(p�11�r���r �۞��" ��t��K�A��(�/Ϯ�h���{�ۙ��>%��}�&�L9]��n� _�6�.���v{g-\� 3sݙ�$�n�A�8�;}�A�����ӴKF����jJ���	$�y쯤> 2���*��gY� >n�3 I$N��F��&`�lƃb'v�so��+���}ퟀ
����@���P #=��&�:ʊ�q(��f`"0v�&G$��v�Dq"w������mS�ޙ��ȓ��n� 	/��M,�>�A���6�lL)�3sk�e��?_.A:S�D�uW��oۮ��SN]�n	�/
�O��b6�Ļ�.��v��{����r�}���ߋi���n�(7��v�u;����\�(n�=�]�у�x��<qv�<m۸����.��t�Pܞ�,�)y�n��6�\=����h�l�q�n����� 	�K���nݺ�Y��8�C�c���V%�gr+�����f��a^N�������i�S.��%��<ciݍJ/l�ϵ�l��q��X�rh��x^�Ǜf�Slmsr�-i{(�<�n��Yx��]�rq�p��˞��8[/�q���!I����w3��O:R �c�-v�OWo���7.�s0 �<�)=W�ƈЎ]_�my��A(����Jܽu}vx y�(�=잢"��O����~؍D׈"66��.��Τ A�������g:�g*�����Do�J���>�>�iu��х8Ap(�����-:��f���"�>t� ^��/� ^�{�#��ױ)�C¾ :��|����ٍ�N�)���H�9:�c��\�ُ�;�G�{�I'���}d�3�y�D�i��>J���>�>�.r�0��s���`��:��wolY�e��,	�1	"��h���J������t�>�'o똀=��]�
����nH��N���6�?~>�~J���bˁ�r�Ԧ��]���A�7��<hȝz�娾���+}=�fsʜg�zu`��s�@��r6%�Ѻ�ƌ�J�^�kp��tͪCB�FP���?�$�ʌ���@���/������I������-2^d�j���BcC�9wV^��"�پ�� >K �w���ޖd���$J�_c��0{;ݙ��ne��h=�wb�'Tz`�4HĬ�$��'6��K�t+��פ��;������P�.��W_�$Iǲ�A�z��^B�mO��dEh�������H��Қ'v�o�O�^�M?&�Q V���:�t���cnK\&f�:�M�T��.N�bz�'�9�[1�؉��[��I�}9?�4I$���X�����"��։�����0��p�!FL��
u^H:��} �*��J�ob���W1_��3 ��Τ�&�+��gx��g�r
ΰ����R�n�>�z�`DnO:�A �ƾ7��7�U{\��yW�n�c=��ʋ[���*XS��v+^N�V#�s�g�0�2�=^92���o�r��{/��[�BULZPU��m��S���T�ך���o1���>'������.C���߯�J
��g��`li����U�1�hU��+�pHGt�HPb΁���N��Fʼ��x'Gp�`���f����f���.݋��?^,��D�J���/x�B=
þӯ��U�Ce
;��謉��*Q�͛��ɮ]kxT�z�:iXU�K����6���Vwg�C7as�3+�7�3�e��6<��T�}�u��Hʸ��I��^����u�oZ ��r��*4��g�gm.#ݠw9�v�	y�W���-j���N��23Y;ie�?9k�����s��xf�M.��6���\#��L���S�N�X�vx�)�����:�����Rm��԰�oo���g�'��˻�lQ`���O=!�����N2���#�/p����k��8a�`��ʀ�=�Y�I��O�3zbR�
�Tf�Ӵ���;in_f�S�y���J���|YV�Z+m�;calzl���^���7��%i��:�c��r���on���;���	���V�X���U=���S�ŭG��_7:��J��z�1�k�C�>暇����D��J�Q�����q�lu��p�������F(8�`uɳ2i�ŵ�u���Q��ph1�kc��wU�>�C�;�F�y�wNs��Ѓ�G��<g��V<T���YXQ��V1����̦*ĶŉD�)V�"(ԦR�ʌr�֍(���D��0-���(bhѕ����lUULn\Q��̸ �YUPA+X�qXb���Yr�m�B�`�-*����j�A2�"(�m5�"�k*���3*����k�����K+mQQP�ll�qkTX���T`�Z�WUE*"����TZP�lTU�-5��eKd��KA�6��W2bV�ō���Ekf44WTu�"�R.5�j�G3V(*"�(�ʵ�]Y���S2��Eb1�[��-����+U��Q13��H�m�%�j#b��b �T������"�UFKe�R�0�ڍ�U��mTQEYa�QA�3�*�0��cA5�cU�EZ�Qs.F´T��"�#�LLAb�X�*��*�6��[`QU2�1��!#������K�o��  ܟξ��Ԭ� Li��w�U�/�v
w[+��O����� ��_ ���p���o+s�ty����bހ�-�.���A�D�c��^~�r�uma�;���~��@�vO:RDA��I\�aݭ��Xȉ)��0 @�����̭�a;@z	nD�-!"4��Ǵ�TM����.j��`�F��"� 7rz�Q<���V�ݘN|�K��P!Za��e2n��7E���gg2,�� 7�� w'�ԑ�=W+ �����/�p�(�Lm�
uV�[�A��	o���$��1�*7R� A��<ȊA�=DZVm��hr�Ԧ������FQwas>@w�)��}e�>@+�of]:�F栭�u���"�vY������yu�a/�=U�`�_�����&(��dO���^��6�X������%����%����ӎ��JȒƜ�1x�|O�_���&�\��l��}�S�R�fDnH�픂 FnNݩ @}~���I�^�5��"&�~MD���ێC)���|�<sq�̈́6��g.?8���A�'o�RցN-�6"vq�� ��۹/��w�'tٛ��[<�I 	�>�-u��	Q�A�#%�e�fb'9oη�<F,�d��` �Y` �7��MW��-��n�iW���Ml8�(�Di��_S��H����J�؝�^;�7;Y�π@�>�R@�7�0$�8fc&6�;��.�s�9�UnyC 32}j�H /sݙ���<�D���0#��*���ΰ�d@�\3���ĂD��ҾiZ�zv���[��_�$��� �7/�A�^z����DӘh׮h}�-�:���5���{�ޱY�}�8�}m襰�Z>�p��f�i�zkH~U3O��,z_����}��-��M�e@Q�;�ۻ/�k�������l�\Vwq�����lR�vv�NG F�q��k�.�u��nn[h.�kpcüR{F:��;9:Õ�m�oD�\��'[�#�[��7YݜE�r�\/>:{!���=h/�����Mt<����c�'�O<��\۵��aw�'p��v8ls��j���S�kj����v�^��PL"���F�e��;�Qaz�S^��앞ۈ8�a�8,=�q�b(E!n!'��K+Ϭ[%%{�׋ ���Dn��֭��۶�#ד�r@���n�O��(�2���'g��VEQ�u�gN� @%{}ٙ� ��DW����jOk���w�iz���	��A�#%�[.�3�A��| U����Y�~������n���xGA$��2�7htژ�a�O��y����o>����qH ������K���ٙ���+^W��3f[pM��v� ��<��|�C�ӫ%�y_���s`?�>��$OǗ_��8�u��J��a�I�sp*�᜸֦{q�����lq�4z4)��De�$�4�c}�I����$�������H��7�@?˯�@�j��u�<)4�__fbF�_��H��n!%U�����tہ$�lx[<��o��x�FՅ���o�Kr�Z�p��˜�����x�s��kU���*Q�+^�%�f�?|>�>���� �s��  6�]� 
��F��f������Ԁ'ވ6eNT��1v���E /�m\��I�)��������H�͐�I�}H���,0� FJ>u]g�$���-̠������_=��	 ��ݙ�7,��k�V�5�%%^%�r	��-���)\�ŲRW��y�h��=�v�VI��$�'��/�� ��m?k�U��rZe��%��!
(6�4�]Sg���i����=��x���?;��]��g.�m�;QT�����W'�+��fbͥ��]s�Ɓ�7_D����)ga��\	�M7n�[����yM���b��7n6y�� �������fDb�n|�˶�����2\ĹM�Xo�z���޻�ݏ�2�)Z�h�gr��6W%K(�j����k�q�ۚU����x'��Z�0t�����R�����Z�+["��i4��us�?/�w�?  ?_��� ����f|�O�%ka(#96Kސ��Q6~.m�� v�ʖ� ��{�tH�79�'��;�r_�c�ge�`��rDC�g�j!�����>�vk{Dږ��-����u�5h�IQNm��A-Β�:����/LW�9�x<A���^��1�c�n�97�&͹��[{C�߽��H��'2���Uwl 6�v�,$��&�On 4L�YA�F�L�W�B��")%�vf�#xL�ܐ�uh:�H�}�i�w+���ޓ;�� n�s1 ��7� �ʟ)�eW�E��i��{+i�R�n�z�޽X�������ʹ����lے�_^���tH=������!�dhm�uh3L���=�3P �;o0��� ��u�=�뙈��y��F=:��}&�xY��{���
P����3ne�"ί�Ev-/��\�f7�)�+�\�ͤSs�IwG|���2#	�Pq(l4�L݄����H$Mb�»�k��vfb ����"�+���b�2�j�=_j�͚Q�&B�rF�d4s3]�k��{U��7=U�ۇ�	$�߯����i#�(�󉮿f}��A�n� �W���Q=��g��B~����Oğ����^O�$�8���v���l@qS�ȫ�[��{^����n) ^7��d,����6�,Ý������JrF��;�dn�_$�^9�iGg�s�n�Ż=]{܀@{����+�
��Sp�	�M7m|zzs(�ّ9�I���ٛ�&� �+�V&oO%��{�RY���b��G�{5�A<l�!a�-�N���R�D���ɳ�L]�h���=���gm�d�]�̈�#�\gۋ?��;�[_�m���2T B����U�ȥ
�a�S�)o�g�0S}�v��]�q���f�"n>LY������ U���)T-�-����8N2\K��۳����=un�6�q��o0�nR���nO8�֎��}��cq�[��®�۰��&��]�v���Yn̬���@q��r�Ƣ�'��8���}������������ۇ�>��v��{h���vWu�8vvϝ��B�7�������c��{X�^�l䓅G��p'���i8����:�m����#�-N8�� ��Zu��U�Јk�u�u�����Sf����������i�Ip����DFY�Sh��vf������+��N�t��oU�u{K�1F|Ƣ������ �c�U��E]�@|nsnl �w�3@%,�w�԰Tސ������$�8���v��V� ��m�D`O�}�~\S�MxI%�q~����p�'�x����"N����\����x+�2��lM�qR�D�~��瘀��7��!��=�Μ��K�ē6���J��}�d�N�I�%u�ؤu�̢�T�������o�J	{���}�����J�%!Rgf��#��m�v����İ�#v�<b많��%Ov���(���%�	wc۶�'k}׋  ��q�꼍�Y���TDx$�W����	��Zى��NՒ��!$�g��V���_ev ":M7��v�x�����T�������`�~��}�B�<C���j�����5ޒn���˜���T��jy���>������ ��{�3��}������GW��x�/-��u]��dƢ�(	��:����$�H��BI��u4��������Ȍ@ �st�VD8��4Ѕ�"�a)��*�5M�[U��������ń@��qIf��G3�s.��6�A�âMy'd����D���n�6��@�o�z�����W�q4� �U�1 �}��,�}h�����
�I����0rF� ��<��k%��N��ɻ!��܉9�ʐ4�0������Ω0� �'|�����D��HM�Y�:�:ۥ����w��N�[�n��I�9@KLm;v~�����̝��l��3:��  #��� ,�}h�K'��9U뼹כ�I'�
�0������N�~�3�v� ��'����s��Ik �(�XH_Hߩ����[���,5�<�̃A u��������k5��uGI�Fq��~Ͼ����Ě'��f� ���VMo�,�dȢ�(	��:��5pN�h�����@|���R �{e��z�ݘ�%o6{�)�p%w�PIV�["؊]��[���K���x16�(��3/��A�n(�E�O]� A��u�$�����m��*�&�0�Gǝ�]�q��d�r��n%L f��c�R���f�����P�ld�&j�6�| ��ۻ$�~���tK��ߢ7���_[�ng�$�����_Z�)2nD�%�$�`-�{s0>A<��U��,���[� G}�L]<���I󹎺K��V7mK�o�D�\�PR�Nݠ��z��A���ŀ 
n�QY�P�z���MQ\�%���.�l�O^��*IM�݃�n��M��ע>�����]{��π��sdvY��Ό��ձ�E�����}Fxdʅ��I�򻮁��xCj׮k��&�#.���X��}/8M��qN͠�W���N{�����o�2dF�w�u[�3�w��r�)8�{]�h ����h ^��0�n���2��R�����^�����A2�@blI���dܞ��Ţ;SыuB�m�pvi�����;��e��L9{�����H"6��w�|o�po���@W:�f�ON���j�kӒt_@���A9�$�ե�RNwb����+ ̛ې~�]��| o��	:��'���P�Z�VP��0���M7N=��^��st����ޣ�2�8�����I��<ۢ@? �st���܎PR�N��~��֧ W��{F��#~	��^," �ӊ� ܞ�;������x��b�,���Ē�Akp�A�$n�{�y �fݾ�>��y�ښ߃^���`;�� |��:�Yn[`��]��N����a�����}�mZ5�5R�nm]Э[�B�m��܉���1������e�3�5�\�mv������h��˵i���ځ����5���$���Vk�$K�(�ٱ�{DoEL���wt)�:��M$��f��`�Y��+�u,��.YZq&��1��>��.�w��8ͅ�;x�MZ[�fV[�9<f��v��]8<媚�pK@�=9A,��VO��I�}�H�f�I��h+�� +���.��;�K���۬�H�Eѭ�5�����'	;�J�+z�=8�9�8E��;Mc�"����Dh�v�n6=Q��MY$\����n!Ƽ�o��Rk��s����]As�,�[�:�z���U�����@7�t��'wܶs*K��M�;u�����vt��w��]7��iU��a[$u�X��s�%���&,7�;��X�:�{փ��[U�mls�-�`=�Ww�^�p	��R=�1�@w��6޿z�!V�B���)���b��S�p^mWV������f9kz��
��b��̕H�'�y>*e�����Ƀu:�v��l9��/��a�٘7�b���(y�$X�r���S���/?��1�6�ngdG���M����Ɂ�j&��p3!޳<�����h�<k3���R,n�kR�ͣ�T,\����!��T혤���ng��۾����%0vo�|o1:ӕ$0�A7to�fUh���u��[ֺٓ)�k���A4g��h��jh����5�h�~R�QQB��,R�k*�*J�[+m�-��*���Z
*#i\��1pJ�m�m
��D��"F��DDR�V��ZU�������Q!JQ��ҡZ��R�UUDejZ6Q4ʣj��b
*��	j�#j�#KX���0TP,�mժ�Z��P*���Cb0m�KKB�*�,`������,EbJ�dDF%�4�tଈ&%"�R"��[Z���*�,���DX0EX�Pr�����e�TDb%j�QJ"*T�Ƶ-��UkA�DV*���`*�DKLqD5��4
0\-D�Pb"�$V%J(�TXԬY�J���+E�X�)Z*�0T��Q���Q���3.��*ԣk��c���
"�m�U""80����,��媨**�J��l�����5u��F1�m�dЊ�q��"���"*�
�X�S2[l�mF<u��y.;0
>.D'=Q��ַb9�u�:�\�z�!S���C��=lv�m����7Z�S���ڸ^Ʈ���i��,p[��<��v6h�玑m�����tx�;cd�[k�2�U2�Nn�W!��nƬ@�/k��m�ZQ}c��1-�}O���O����Rf�<;�y��#���\�ןn�u�]�C�-�8���
��w\>K���{v��z�;,�.1ۋ�����XD�p�^��,���s��۹d8���qٶ�]v.��/n�t���T�d�n��On�f�x�n����Vl����[�|�%��;��ḵ�q�Fmtz5�����!t�v���v�3�.�(�=�cQ{]�ŷح�DCAog�8Gf��Cn�m���p��(�]Kڧ�9����^L��;���ۤ��BL�v�zٛ{1�fx0�z��[����=b�pj��j�e8��v�A�m�c]��nּ)F�%N�v�@���'����tިԕ���kq���[��u�6��^�I9Ԗe�[xsf.��,8�.y�4v�Z�:6�n�V�۶8�^N-������\���\�6�xL���f��F��t�<�]�=��糇��������͊�Ն�gW/3��X���h��!M�v��m�*&onz�lu�Xq�{s8{>E��c�o���ݶ��3��#v�B�����ͣ�\�;�<�]vz\���엨5�KW=�s�����m\lvoh��:�ArzΣb�]�v!X�'Jg˔�=W
�t�g�]�MgmAh��{NM�:�v��N�Ψ{z5�ù{nv�tS�c'R�f�NG�87v[�=ٺ���ْp\�����7+�����z�g%c�n�v���齶ax6�9+��3�5��q�T�(����凍�����v8��6�w�;��^����]�=�gm�"I��s<��p۞0n6yt�91�8��g���s�W;��������⵹2�2p���
{%�n�בut�h���Pu]�����Sh�h�#���|m��sp��G0l���j��f.�<{s�<.�Gb2�2�<v�Y�nM%1�x:w��­��x��պiǶ��u�@q�^�<��9�>�����@���h�c�5ʽ�-�8sS�n{g�#�W�\�Nn�kz�խc�j��w	F�����On��mѷ6ܥ�^nm����i���e����r���gp�q�T-�^'X�'Y�\��zn��i-������\��[5A���s]�����<�F��ί��MVv\`�n�  Xnu����[d����n��	2v`��5�~L2"0�.҇����K:�n�i���%���d�� G�?%��I�j=>p����	`�=��D�C�k@��c�Mh��- �L�t�����u~�� ��kt ��λT
���F�H�X�K�߻r�O Yd�mst�@ >��v�ٝقi�����G��:�� �k9@KP�N��z/�N�Dnf���"n�d��o��F�n 4�`� TI��ͺ'_�r���'1�d���6	�&$�6Z˄;[=�����軍��][q��u�.9K�����{�[6KI)�������>����v�ٝ٘�+�ogty�AuM���ݪ�j0�b%�3%Z{wٟI,�P$�퓽n>��î]���M鬌��#ӈ�l|N�eOF@�u<=wuT���v;���(�U�d�s;�T�~�fX�Kކ����@}���v����I�'ʵ�c�@��0�ˆ����9w0���� ܾ��~��s^��}�+1��@#l�]�@%���s'��A9�6��=$��e�,�|� K+-[�>ܾ��@�o��2u*��f0��z�o�m���b	*Z��w0bI$����q�]]
�W�#Ps�shٗ��� }��A3SG�kݾ������#]��x6w%���y1�7�9��l����Y:��K�"s��l� 5-Cm?W ��6�޼� "o��R����u;���O�{
��́ ���`�Ť�H�fa���{��y��ӆ����[�v^�f �}��E ��Fl��=</�к����Jg���P�2]�N��bX�G{[�� ����{�}����!�E��cf���c�qͼ*�mUv���V�!4:<TGt�2�N�k���z���b��T����d�]"��}�e����~�������$�|iC�H��9v��׵������l ���ϖ ��S��#l޻�����FQ&�N��$�2y�' RHӺ���	$��}�o�fi��{�;]h��ٙ����  ���a�b/���j�x�����r�mNCIQ���Bc�H[I��[�b��\������}~���!a��d��۹g>	$����� �.�"����*�y��WN^l� w�JI|�W�L�.$���c�Of���z6Sכ[wq� ��q_A��rDAU:.������V�� �Ť�D�fa���y��2�v�D�$^Fv��5�-S�I�@��  i��֍����Ɇ�f;����[/.�ݖomF{~�/�> 2�햀��׽�ج���q�B�n�e�M³7���� 9}ᷳ&֘�&�c�`��,�:��)��{�&H����wMhK�8T�`�W�V��I���H��������.��������m�uS��t�߀GmS�@���J��|��6p��5�w6P7�b�]l�Cc��l7�;ä v�n8����nň�J���pH RH��&䓂@ ���	����0�:=����k�	u䄚	 ���ѻW����X��*;���2I��h���u�s�Fe�� ߧ�Z@ �^��@gcr`�Y�rbA�k���i�d�U_�o�v�H��y� z���T�}>q� w��ܑ}~���~ZL�d8�jF엽%߽�ݧ��5��	 �u�]Ȃ W�ݙ��nsf{*�qj̬��H�y�#s{��d�L3�5��f Gf�A�>���E��y [�/�׻���s���OW�]HǺT�L��	��Qk����q����R��u鄽I[�֞_�#R�_-�6p�p��w�}Q�e���e�Q��-L��?���X>���<��H�:���i8[;n��:�V��[\�)k�ߕ����m3��% v�=Ԝ4���Lz�W�;�ѭA�'��cr��e�`���q��.:�c������n��k�u��Y�t��[��ᣏ]���خ��sf<{'F�3mǅغy⽋���z���q<���M�Rc�rz31wl�p��x����Kq�T#�۹�{hotɬ�5Ȼ�x�wϖݻ6w&�)�����kohz{z?t/�>'��9u�@���ݼ�A$�T4�m�.CC<ϝ���s�jH ����@X�;1�m9m�n�:�� �623�����1 ��{�x� ���DGo��d�^���`ij�XN�m�JIr�U���� 79�H�g���'}��b@ ��ّ�H79���'+��P9����wV����룫5f^O ��x���S�A|m���dJֈ�]e�����$�����F@�r7Z�=��DF_Nг|�c~��9�0���DGf�_����Rf�/���˛���ح=t5KS�;�3v�g�vm{W]���U�:�D�>��w�;Q�Ss�9��1` >����@-�}e���z�����vdF$�n�J��#��ل@��U�����'�뽿K����-�i�g����父w.WW����p�c���M�8�iw�.;�炳�wZ#��QX��t6�g*�V`z�	k}�A]pr�	������U�S��{�� ���DEn��$D_��"W���g�K�@��	�I"�D��bH$������PH��x��՚�{�y�$I=�%$IJ�_]�ҥzXN�m�R0Ir�o�sk�y�U��"NOG@ >��X
��f(U8��퇹�3� W��3*�P9�0�m;�H3�=i\� ����ݟ7繰/&���>:��R��Ξ�"��}٘=��ΪA��f� ��(�#-݌q���c�h�;�v�yn��G���Z��^������`�m2������+6v��A���V���]�P��TH$������iM��q����f;��w٘�\�:vܲ/5�|��"�u������ĉ��m�V��Ԅ�a�Ga���8r�«��� �+o��, 
I�j.�[�z;Vf�]Y=�1�S4[5�,�ld�#��_0E�N�U��Lrn#���sd��^��}Yr0HJ��L��K?|�Y��q� ^��ܐ�z�~�'�yf��I�]Z]U s���`�"���W1 ��fb �s�ױ��^�{���^��i
W��n�m���p����X�F�7A*�׏?uz��=������+o�3 H��|?m{}���k�9G@��	�?�YS�<�h�e����N5��2Ƈ���J�����NF��,w]�ozv�Ȑ[{�p�4H�����|7E^���m�@����s0��I��a273vy��Kζ;8�xT��5�<��� �>���I-���mGY�s������$�!��ݞw}����� �"�D�Eߧ�"�y�� �/w3  79��uB��ҥ��×v������� y>Q�	$����I�����������mC���k�<�V���S�=����Y�/�N��/ol�{��m����F�7O:c�=:��Mp�<~�M�'�>F|��^�������y�%��7uk��t� �Dm�����S�윛v$�Y����٭�D�����C�����eQ$�)��Y���c����v|k�}��C���\��<(��|R`�ew�V{�0bA"N�7_ o_Ya�}����N�V�5��31  �n��z�7)�܍�N^-TOI~_+4N�u�P�?.�MQ% �Χ��m����@�iO�}뷱�g$�O�ۉD�-�#wiM�( _N�W1knc7���@�7A ��]����~c���c�[.�3kz�w�J�zJ	��� ����� /׽�v�0��9y���,�����k?1"8c�iJ�v-�{}�q�!�N�K�S}�uN)�M/_%d ��$��E����k����:�6�����^E�y��Vmu����S��%�:S�m.B�F��6�=N)��37K�[In��#����cs�	��-�ƾ�(\d�LB��ѹ�����E�\�v�����w�9�� 8;'v�Ǔr�rv87�����'M��A^;uQͪ(b�`K=���ꋞrv�X} ��V���p��An��=�ݳ�l<Gy�.Y��ݭ�� �ݫ�i烞}�v6]��\�ޜ��`M�k=lM���*����,�P���2� 8�{�85 �GsF�}��u�*=-�*kwl#�a�i�h���n��������2F܎�U��n"��N�`|E�m�7tB�\�s����	k׶�ھ,&��($�3}޽�H�����^q]���o'�XD/e�fb ˮ3�݅v7��g]��1�2�D�wV�Nڹ�n^��� �.*�F���PD���$ /]�f�'�ۉD�-��Wa)�#G"�q̞��ۄ�Դ��I-/so�I$��&������*��$��w^i	�\�-��
&��'��8D���A%)�Oz��q%�Ċ�@5�lD��ل�g�2�k[뢛	�)���
j#5��u��b۞B5h-n8sg�N1���������߽߉��a���J�ՀH;w�V��o��hJ^�7C���E"K�(���<L��5�U��_Mz< ��Uʝ[�g��,k� 7n���(��ڑ]6_Z�B�β��o���הo\SՏ�Y�Ձ��R5A�*5R:���/=v�6y�y�?�s����AO�Ͼ���O٢����-��W/�:����	�%0�
	%z�޿����$��Ľ�{_e� u�u�$���J����q����JR]���꩹����iz�&��u`�N��B�?7s��ݞH�E/$����v	+�5���[qF��zP$�fvmӪ����^�q"��.�ݾ��D�α]yRo��5�s"%np�a<���Qs���(���4��g[X��s]��v�9��e�ʮ�`�s}���;���=��Wmw�%�5�*  �;6��t#������k,TBt�~=u�1�V�H'w�B� �7s�� �^8�/	!q�=��/��/<Q�&��C!�`��AD�f�u��>}�K�/���;�PDy%�g�����!�.-q��(mL�Y��(��W�t���+�����K��2I�*����G���x�{ό>�����<:�]�\�\+r��9A��d��c"^^#(��c�C���5Nòܸ��&q�uç�[�e���wc��O�f��=�v��/>HG�ؽ\�;�m$ξ�^rd��6��^P�<�~��KjOr����ԼKL�<� �(���*�&AӸ�p��Ͼ;������|�Apn�+V�y�Y&kݐ]�x'�&ӏ�Ĳ��쯕Wyu2�=U�I>�P�;��L�VJ۰���f�����%'+�����+��%��t�����)Շ���p�\�t���v��Doum�a,�Z�2͏x����q�ճq83����i���ə�����`�ѡR=r��u+r���R�W<��IE��2� �#C��z��<��W��v�]�}�_a��Å��o7�%B$]*W%b�O���Uk�1�`s��? 9�ḙ������e�X�f*�/���hq��&r�$y|Wu�컈r��J0����.��b"1.]}�a�{��i����)��Y��9׼������J[��R�M^��'<?!A節�ݛ��+]�lA�6w�j@{�+5����׆ ��h7	��y�]F�_3�m=�-T;�v�f�Dǧ�����rl�׍1�;�02��O����~�Y�˹����˅l��uG�8%r���������i���8�ze!-�l�a�+ <��_rYy!+��`Rq�7���T�eK̰��KQb-�����f2�X�֠Ń�)�*���k5�&	X������DX�#�d�1�b���[D��a��"�f5��V�cZ)[�2�hR�b�mb�*"�U�-�b�T����ʵ��۹���k�9h����V��ҴmR�(�h��nY��"Ȫ��cm�cq���\q�k1��.�V*�,�33!U��0���QPS����b�������R-�ji�M1e��U5L�U�Kb��-fYX��b�bѥV���q̩���DV�ێ��Ј�̴Zep�ֳB�D��*T�iZT��Ū�mi�c+r�ښ��I�X&5�㋤�2�mR�5�.�F�֨��QQ���ň���-�U2�L�t��U�X�+�ʍ+P�*-MXS���Z�mUբ�)J�ePb*c*֩-����?y����Jf�uX$R�h���($��׻��������IΙ(H$d�����{ʹ��=�7ۈ
J%W��n2�r�ngo�~$��z���y��N�u
33��>�ޡ
�h�ev�ϯ>�q�-�:�֩�9n�gms6��qۢ=�0��m��\p��.v������`��6��zw�~"gfՒ�����o~�靍����Е���m�|���#��j۫��I
��e� ���;������K��_3�1� ��VW�������Q�v��'n��`	5��!�玷� 
���
�{�[<�&&���!��}U����yߚ����ؐ y)�T�}Bt�X�V���_��B�'�]��]���yo���qjw��Zj�U�B-����I'�����YX0�y,���z��n�i_�%T-0�
	%}��u�?w}�v�8��	�7��?~ۿm�?{}Ҍ|/ָWo���{A�o���J��6��$�Ȩ�͉9�n;E�Ӻ��pR��9ՙx2���$��$�_!@�����'Omm���U�W��>���*B�ƶ⍷
N�|voJ�t���6�y�{��Q��|�K� (:{4P�e�k���񫪰fu���(�fU���vI �{e���4T�¢�����A��vA��"k?(D08c�>�7���S�D�߲��$��� v���gWz�w�>�5P�(�M� p˳}U(�'k3�^����[�:'�T(P};6� ;y�*Sm��G�{72���7�޵��X��ݳ�xh�5�7�
��l�;�O?���{o�{��m*��n40�V-��>�u�<p}1� L@� cV�n���n-�	�b��2�VP���"c�[sWce������r"v�S��Ӡ3a�i�ʽu���
�[�e�H�i��8��eJ���.#g���5suFv��[)χ�R��y��7l��6��]��v�|�^Π�l��e�v�מ�$�&[b��z�Oo=�Qu�n6�%W���� ]!�c"�d�	�m�۷Nw��a��i�M�P�����ց[L0��Ië��d�I��A_H��뿋6hJ^��]���O�w�(��{.ĎDҎ��K��O*@[5��7�]ģ|u����H>�t��$mnu�$o+���Tі�vp$^:ۊ6�*8"TM�(r�6Ń�<�<������W�F��]�3mi���D�2�-��v�qK[��e��_#�3�,�=��k3�q���h i�APf5��B1��$> sSچ]v�l�7��{1�h�S�@PS}�q\YN���P�Ҧ#v�����vX�Z؞ �\tvv坞nF���.6�$�y#�LM7��7��T� �v��� ��ʤ�o�����L�~=W�V	�z�*���P9+鹝v~ƺp�e�f�3�^�{^wMYh�}i9���S������fdXE��N�N��;��@^k�Jf/zP�x�|�<�a��Gs���}�`M�w]�@=�w��W4�w�]N&��bG"i7E<K�#�_/��{W�(W��No�w�v�O��'�λ�H���K�:ӆ6�1�"C_t4.��	����^�_�����v��P P��D�C��5@U=�d��ֶ$�@�a�v�����wf���@
����
��%@|G���A�����y���k��^h~�߂?)!;u:��:	���s�]3��>xq�o��!����ln��==ÿ��!�08c����W�����I?{{hQ{U����`$��[�=|��F&��� ��o�J$U�0�]&u�޲	>�ޫ�o�Q<��knu{ڭhP��D����3n����P'�~.��s�<�O�T�"�8���?H��1�n��çz_��#'�{qG*i�gP�uZ[�L��Bu��(��Y}�R�4��s�1���Y^���m��t�}yvn&�rM��'��cEZ��B�he��_B�Oem��yM{ԑ~��@
�l��*��m�p���{����w9�/���Yד�E�� zN��P�.��w���y�[g�BsX 6O�!�`���Ȥ��n�x�m7@xM^���e4I�~�>���ZA�L30�\ ��l�A'mw� ����I��vmP��
~d#�r�~��IyٓV{M{�e�e�}�;}�(A;w�v	 �����o|��/����bi��	w��͠ ����Ln�B�;�.5���}�l�A���{�E���T$,4J��_mgzᣁ�-�Ӄ~+�h (�D����;X������Y�����Yb�pm�̫��Ǟ|�$ۥ'AH����a<��u�d�%�����<]GVY�E)ρb�A���>k.ĉ�cJB�rǧ��eoU���mr��+�ٺ(,��СM)�Q�W���a�g��PS�b%�4L%��p�k����$-���X��9ڋ�GUr������2�dđA�rgJ$O��n�ē��kە�µ�w{=bCT�$u�z����-!$&�vN�5Y�`�H��ب (��@UG��T9�[}��<w�0�7��d#�r����Y$P��T�PS��x�-cͩT Ju� �+z��F�,kQ�p�%پ���H�-��A--��{�Qn�>�{:��}�u�eW*�q�=�vU�O֫%P���*%����'�N��(�7����`���T(}��� t�Q��wRm������bW�r���*���he}x�W��o'"�NW�Z�dan]��R(�r9��ֳÃ����o${}���v� L�`m��Q�u<��:�T��LN{k��zh����ͳȩ �3��^��L���vfwn{<�Rj��nk�r�we,�OWm��퓱�x��j�q!�Y7�{W�n-,c�<)�����!��ܻ� �v]kv�T��t>J���t��}=�y1�s��4�y1�zk����v�.m�q�s���6̜qXт��޹��НZ���6���[�c��:5Yq���y�O=[;%goϿ��Ω�"������w�ł����'�A#w�_<�}�+|`�u�uGݾJ�{�m u�[qF�r"Tٽ(�X�Gz�L�۳N���C�{;i| �=��@s����wU�}��m�-!$&�kj���͛� ���EI�k��y��w��lY?o�WĈ7��e�p'�m�x��[��6m (
~��o÷��N��/�zn��=�	�^�r$�Q��]�o��A �gQ��U��������g�@Wo?*�噔)I��Z�n�t�;�@uqma+��v6���m�1&��.Z���<���Z$04J����;�`H;�t�H�6�:�'�i3�V����m�$��w�W���$qҐ���;�gX���i<�܍�vk�ݍ�w��[x�r1�,���;z��[�f8٘srM4�{tV#��vħ�E�x�z������gWps&U{�	�{`���]���=I��W�IU�@���!��9�OI�ٷ��H0���wjUN���{`���d��oIi	 10̻j��7@�>^O]�$�gJ��A ]vm�$�/z������6p$��_@�>BkH�1H[�\ݻA���Tw<@��Pymm
[�H�5� �^�{3}:g}��j�y�m�Y�������)�����o�k=s�\�l�${f��_G�=E@�mE���UJ$A��m�$e�U�P�䙕�]1��x�۟Q"�3�d�V��Q%���f�~>�Bu!�^eqO�3�U@v�����ƽ�N޷v�a��zp'�̻G�("&�!�>� �w���zz������"֟a�r�Wu�^�����ǝ6�Q�/e��^ �^���Lֵ�W;;��uv��w�I�%����(<���A���I�չ���/z�Y���P��04���}7JL`�/��|i��ŐI#2��@	���j���>�T~�u ��%v	�g��$�$b$�2�mW]�9���'p�:�@U�^H
�]�  ����҂��)4����j"!@�n�X����j�@�t�m��Ű��z��o�����1H[���W� �_m�=���}�R���:��\��P�^�B4}wl�Fڊ	Bt�	>���=v�ʺ�߬�H$v_u� �o�P �r7}��û�-���oċW���X��˒������Gä�m�����q,Ҿ���{ڨ�A���{.�F`j	
r����굫d����	��O��u
��:��]�/u��A�U;�tU���BM^k���gy�!��z32�� Q[E���9۸%^��x\\uK��wv�[y�K:t�{=�E=*�sЀ#�($��ӺWē��vm�5����Z��-k`}�[J����߅ *�nu�ڳ��0W��R4$E��"���f�n��Yk	uc�Uzp����$gY�w������-	�0��S+��$sw`�O�չ�d�4��V�B�uذI��������I�$)��۱d������ܬ�B�}��� 	��� b����W$q��FLm���'98����������K�g{� �٢��M]�J�\/HnB�F&�����נ��vA�](�N����$��u����Ϭ]U�=�W�3pHT�`��V	��o��*�qd�D�>���.��[�MS���y�䪇����XgOi�
"�5,��X��o�}/���X�>���^+���틻ff�o`�T������4��I�>GAg������<���6!R��G���d�|�g��>{'�n��,�����r9��'��c'K\���8f�v8BX@c����1S��x����j�ѽ�']�鹨�������j�w����SQ䣾����h?�'��Mg�{���)���w�9 .n���ϯ��q��U r�<���'Y&�Y-oH41cE���ѹ8d<��}w�Oz=���V&gl�Z���0��>zj7��{�RƔF+�9�[�7���^���8�c;k�kN�B)nӛ�]t%윆��[�����`��w���y��s�6��YI�iu(����G�Ʊ5�^�a��l��k���j̸���W
qPhQ��`bھg�R��\��o�~+;�{��}���W��`�|���/#�*��Y8m�8QՓo�'��)�汚�)�3�q�gz�r�o��f��rr�!�j�/�3���z�\�*���	|��g:�޷���~¯��hR=;řm��W]%���qE[@��ǻ��kj65.u�o�v��������?nt;^ ��u\�u|3sS�J9�-;�s���� �S^�F����"M~�}����y���f���A�ai��Mo:����Yф�W9F�8��\Ke�����5��,:t��,����͛���o��� ��@ q��Uq�m����2Ȉ(�S�`�-X�f\E�TQA�q1�UZֶڨ,F��F#P�Q�Z�Z�����DTEh����DQV�����Qm*�.�#ȥr�0��b���[+Ee�([E�6�*���.+TV�#n%�?Z�Ŵl��WU�WT.YAb"�)m.:�ЦR�����D[n�3h"�ke�TUqJV�
�m5n+Z�6�GM"���b��AUGm\�q1m6ʙV��6�5B�VZ��GW�V�A��
خ5�bm���`Z�r����m��MF�*(3V[t�0j#CM`�f5n���LJ���j�&���J�dRUZX�VcG
�Z�n���� �[eFZ)Uբ��WQQ���s²�,q�`�{ol��|~��.�;9e�>�W��w,�5�t�������xv�^-��l]r�!�ݝ��6۶�<r��5��������z��2�:nM�����r�]G<ˁ����0:�񐻬Q"�ml۲œ��;vȻ\�[uhģM�2��ݫc���m�%gnw"m���[gOy뷶}��%������mZ�����3TNsǥ�$� �No����y�8��ݎ૨�l.u���7<��득�����q�m����;gn'z�Fit0B��E��j�c�a�#;p��7;����7+;q\v3�7I���D�"�n�qZ]{rl�1۷	�rZ�X6 �����:��xƎ]s����uƲ'A��s��#ݎ�A�v�gT*�uumQ�^��\>ہ�]��b�3��k��p�Gl�&}n3�;����׈�lc���d�z��6�Ca��n��sq����m�u�[���S��ŋ5��5�ڶj-&���qű��줽�#F^�|�cЁ�e�u�1���1�k'a�v�η�އ7��v3���{X��]�r��.r�6#�ϝ�!����+ۨ�;�r��|��Iw�c<<-�]���^ǖ�t��^���ըwl��1�(���F�Cc^�z���L�\ٹ�v��Lr��v@���6�u���z�� g��M�xm�-�;n�8�D�.wj�K�y;uts��Z�����lcI�c{u�"�t�؝#nǜ\m������ZԺ��+��R�k�n:�7g��3Y9�=ٗ��#㞞���b+���c�\��6v��Ʒ�O4����G�S���(�n�3NH*�Q���ݲ���x����G2�ۍd�e5���A[���7n89�=������vԚ;l��������nNGv��lFvx\�%P_8�W<=D��u�uƻk��Y���2�d�B̐[n5=��2N��v����;,�:P67c�ܙ^��/�s/��^�e�듞��1�ޝ�:�07UnX�r�tSŹ��qk��W��n�>Ֆμ��2��NL�sף��u�v���8�v�\��i�V��d�%Ñ��nrq�>7Z6��V�%�t�#�ے��x�ݳ���(��zʷ�����ۣ;;+y��@Q������W	�����x��D����"6p��k��^¬,�b�Gphn1�ΰ㇟U�6���뷨v#^����N
�Cv�tW����+O���9�s�(�tTtg�mp�鵦㎌G�,��A�b@����m@ɿf�D�N.�t�A'�}�d�w��	��;�`�U�?�y���[�Hh1�	D;�����.]�̾���);�~r��v��œ�}��F�2&�-:��4D�t�4���d�IE�mذhL��@ 
��g��G>t��� I?d�u��1r~��"d���Y�X�y�yΝH@SΞT�N�f(���E�쮻ھt�nB�
����/�
��ݚ2p��K�T�{&�C�'%�Bw�6�5�ٻ��L��~v_�I\�e���tA�(�}1�n.ϲ3ۢ���E1"	H�O{9�0�`."��sٝV	>��U�?olv/@款��VnV�A?eo��S���	��5Ggt�A�����dz�T��+�E=���mE��ٝOo�q<�bĲ`8�Z�4l�g�<��;+)��yx{�"5g��z��B��[�!T(Wl��� '{�E�+=W��F)*��_��$4�$�2��&��$��_H"�H,z���"tͥS��ӵP��٠c'��HfHT���{Q�2��9I���{���	��GI�s'`�k��,X̰��$	��F]�k�ADP�߶_�=�g���5 *wv}� 7s:�续�n��<���"˒�sm���{&vͣ	����Ҩ�a%t��a�z������0������'	��]�I=���H w7�&7P�MS���i|>}�J�U��f��).�����ae�Ok��Z]��VH�Goz�Iw3��"���`�l�{��O�^�����zP��fm�d�S�C��*���%�TSm���6��M�����|Q����+�e��5��gx����ס��	#�)�y��)�q{G��U��nl�č�λ��Y��2(�˱�������I�L:E�T�I�Ρ~��Dy�W�en$���T��	�5�
���@�j��$��mX+j�C���P�%綴P�$Pg��zp�\4��;M�@�bE|B���t��v%l�}\s¶�n0����4��h������� 9�gz�[��
��򥳼���������ԣ��s����ڌ&�j�I�n.�H
����JW�^��@Sy�"I���~=�a?r���̖�H(N�E��ERV��۲	7=�V	 ��f�g��J~������D��
{����� �(�`�ƨ��H*�s}[B�N�H1�m�$�E��݀Oğm�_ʻ�����A[���B`�u�v�l��RL�32U����v�Ӹ�oP3��%ʇ�&�D�g��We�DC~��v^j΀��qƘFU���|���߂=�7}�~�k��*Wfȕ�=�J�� N^�
m�ϓ�T�bG�7[�X���q�1�f�Z<�������o���[!����M(d�+���ߜ�ܴ�E=���.�v��O���
|�;�}3�*�/n�$��ڿ���&��N#*�]T��&��>�95wJβ	$;�m�Ē}�҈?���Ir��eh6k�M��	B����}vI ��J�p��kn���{~���wj�$����a��1ERU��gUWn�`ܙ�����U�� ��{B���H�޳:[�R�}3J��U�JU�!2�e��EEo�Q$����5wW��G�QK�@C��߅
���|};%js���a��T�\;�9W!�4��7s����uՑT����~�{�1	����v�ٓ{�л�����hQ/��љQHB�M<v:5'��nۥK��/#���{C�����;Iv����y@�x��;�˖t6�j��<�0T�z���z�wξ��S��kjӷk�y�u���xrS8�N��3�3�c.�j6����=��.���M�sd���Ձ˳[��/c�q���)�%n��5rFխ�U��mso	���'�tW��#���S۸y뒢0�l�7N4�8��-��;hX��&1h��F���{zPBGa��J�� �޽�� �}W�v<y�í��$˻'�7�e]�TH��H$�_���!�]_�ua?�ξ���{�d�Ό'V���46�e5�Jqvv�F����&��Wjɓ�Q�������*��j�%AΌ6�f�I�s{)��W�E	 �z�|P���"�Z��c����|�`:{�@�˵a��GRU�v��v.��W��r�R�;���$m_zŗy�V�[��wm{b��" [� �(BYa�3�G�u<��]ح�T�����c���}�~~�9�P��⳽(��۲w��'��2�D���@�n�:�̀�P�ƘFU�vo��>�m�~���f�wͻsW`h;;�w�&>�ߐ�~ɚ��V���-����aP^,7�J� Nn�$��5�U@�2���o��8H'�{�Hw��/�k�`�́�;���x#�)$�	 ^�Y��sݵ� ��χ�����>Iz$�,~�_�Ղ����R%.�5ҧe�P� �ٹ�ċ�޻w{"������Hꝷd�U0�j�'%}/�%����m>^MS����+蒠 Y=�`�}���˫qE�v�XH��
"���z�������G8�Ơz8��>n�z�%b���Ԏ5�I|{��v.��W�od�͢[�/x���v	%���Z[~A2�qA!iD5v��R̯o��hΓ�PԞK�(;�4P��Vf�oK���m�>��C���(�i�e؛+��$��@�I��K�ޡ�݂�N�بlgT����tk�� ��9v�`TۧJ��ΚO���R��3H�_٫�)�ެ2Y�23����K���H��TH��6$���V����]� �ud�	�����{���y@�����]��V�6{*��N%C{w4 j�T�NZ���\fԏ��K˰H$m��A ��W�b�l��1Tȴ_*�@"�Fx� �� �A@�Y��r�Q5θy�(1D����~~<&�F�NNY޻ �w�҉����K����܀x<���)� (?.͠:�a�#�G!RX�Vuh#G�Dk��p������N^����w���c%�{v��1�V�[z�e��BҊ�?t�H��m�$]�5��+�I;���$]�XXz�"�J9eZ&��2+�8&ž\�@���
 D�j*�Ou��3�I}u(�G�g.i�|uu�g|R���K���3%�fi��gK���kԇ�Iv�'x�g9�B9�]W�x������u�$�ʂ��.UI�dM�%��{�V���쳶H��ڭiNHP�S�J���l��a^�+��1�z�q����=���-�7gCd�O��!��V����*D�	�N ��;w��B��jg�����{Wf� �~T�J�����.��vE-�zy�Xٞ����^�T j{�|)_�(����5ҥ���݅�5$�Iw�����;ھ  k��E��*�{~�t �}�d�]��쐗��&X�H"1(�u�e�u7!�$ܜ �j� �]�H
�ܽ�
VӭA�f�Q>���Q��(��6W]�I �^�lg��~��w��|��_Xw��`�H;�ҁ_}b��<*�l�t����7�2��+#�x��k�������i��Ck3�����u�n�]jw�5gA�����{U�e�
��@�f(#-K2��ΎLk�q2�ne���Gc[�v8�r�nzമ�/7�u�F��1��÷��Mp�)�F����6pV��v-0wiۢ6����z�V��{!go:{sc�\�Z|V�G��vΧ��q/;�Fy��H�;���q9v_l��`������:.-{U�uSsB�:�h�7<����ea[<tsb�˔ݛv�d��u�W��ԙ[��n�'s\��{��qn����-��O@���q�~��Dؒq}Yv,�{j�$�7o�P��i���v�%T(b}䪀���(��R%,N�a&窭���۽U��_���گ�$���A=P���`n3�a6���A8 Q���'�*��r�W���U�Y�s��$��u
����_��
G$����gk=�묏�*�BM��D�	��}B������B��߆��L>�yTQ��,C$�U���͠> E�ʕks��������
�Ϩ}}�v}��,�/
��"=%���v��i1�zۭ�]�4�X�	�C�7b58p�9{���E[���@�A���> 
�zcr���e/ϝ��6 �g�d��ʣ	6ᅱ$��]Ճg7"?.���;_3kKJ�KG��4ʻ3���^9��g�r}�<,@�� ��-�N+�kF ʆr�*�=R�*�A ���P�I z�:�B���s���t1�v��Oޭ&�e�	�G�[�[T �ʐ����OP~�Ӿ���} �V�]�1Ma ����NJ��VT���z.�ytʻ\I��
Q8��)�m�<2��¾�Z�h�+V������;�� �y�+� >�ogR�Ψ��o�>o� )�A>g���s�	�s�0C0�RF-8�a�l��YF�v$r�-q�.�z1�����_���&�H(���J$�3lY��B����g�
��{��t#�� q�$a�	%$I�e^��@��Ӟ���d T��@|~�և�5��wu�:�� ���/S�4ۆ̒�� ���(	�ū=D��8�y:�C�_zn:�s��LU����졣�P��b�2g�IM˭9*����7f���m ��s��Q���ͼ�yhk�����y���]��{r"���j]h�n�\�8ˍu�M�x[,m�L���m=]�j�7|Pa~���A�Rc����]Ee��:n�=dZ��u.��/h�j~:��������#Yt@c9�%����嗲J�J�����ל�1WT�ze�Z��Y�'e�����<�
���R��e�i�C�� _�yŽ�v�S*�u���)N@QN�̬�q�m�M�.@�k��o:���TH���,����/{�Rg+My�_�C����_zQ�{W.��v�{�8�GL[�Pb�=NҨm�Ć�{�1O���E�a=�9|3���6�-N_
���	�D�'�\�P8�^����X;�0����OwqY՜�wM����i�ի�����L:פ�J4��C�I]��vn��̖����])�XR�f����>���'�q���@���c��j�1�Z��awC�����1Z��.$-�,��Ws6���F�27��|�~��9� �M^ڃ�n��<��#g8P�&��{�u����aӂU�ʼ]�tY/�ZYr��V;�hg[����5n,�����FYrQv�Ey=��&��H��>)�}����cȣ\suWa̬7���}m�!w�XOGG�΢��,���Un����gJ�p��:�'_)�
������=ߔ���ĐI��W���T�ޮ*����.R�@�c�̖��0�Vc���V�Qq�5Q+Q-��5-��Z��-*$]�Z������W
��Ġ��+[�a�h��SyD��Z��]���3z����4�L�W{�"�DWF\`��bHͦ �F"�Dr�LJ9M8���4UPP�������ꕊ,ձ5j,V�-�%��*#k*b*n�����VU��J+�.*Z#�1�:KDTM�b���Qh�Z�6�V�)���J�V(�"��̪
1�]�3J�mE���E14�M�!R��ժ
�QMZ²�I��(��bdLR�\݆m��Qe�L���F �b;�(+ ��Z�E�3-H�ATDE2�*1kX����lm�!�Z*�ڙaF�Drرբ*����.B�iR�R�����4J0m��V���*VX��*".6�UAQ��b�UV2�UT����ة�(e���"�-)cڢ-M^l�X��9;�7��I�o�@��`�UE�ZeG�/m:��W_�A$���A ���Բ����X뵸o岽�.�SX(��j0S��\�H$ft��ncQ:y��^λ���_���|_��Vd��P��N�`~�e�[<�>�m��u�g�vvG���l��lq�aLH�R&��;�Bj9��|s�T+��{4 (	��+=ΰ��]�s��d�~����3M��"QP\�V�z���r]�di� �ݻ���ΟQo~�e	�W~;ϯG�f��E)M#.�Ϊ	9ٰP"�W;��v�u^�$7;����Ҁ$MнN0�rS2J/���ۯL�łqw���J�H�͡D��yװ����ct��f�"����U3����=Z7aU���C�o�e&�5b}��G���kOKFO^99��:�4yVG�^\B=
��/+�.7~�(�7~�<��[�H$�2��]U(�^u�����hwmR�d�P���UC|����xa��:�m�%$�h����$\WcV�ܠYEgW,�s�0��O?~��ǃ��20���켡Dnf�'�μ볝c����f�qO�mU	;=(흳a5��U����K/���3]ܨ((/��6�;�;�9^�?g�M�}z0$��&H(���(��^m�'�F��y�vו�]]�߸	��gJ?�o:쟾���C$de4��
��R�g����m  sN$(O{�ڗ��g�2|H9�R����N@�fI@����������v��/�h&;�[T �9��>���F��qɠe,��yc���g����F>�X�gc�b��:��=[�H��Y����&���[VGds�KR�_u�[�Mi{Fs��^^���'E#��#��I�	�cj{t^��B.��������qd�ޝ\O`K$�u.\s�^��ۂ���sY�;f��	�v8��=̹�t���W9�yݹ;3דg�n
ރ� �O=�{�gV\ �	�]Ux����]��<��[g�3g���[��r�@�wcMF�Yz�Y�.,�p�.{[���c�a-,n�v���6���=���%Ŕ�E����Ω�Q��'6�s�k�<�yX�x�`1�b����߯9RA'��YU(�N��� �}��_��gاj�U��<(UK��|ӝd��%nM깄���Z��km����(��|��P:{kGp9ѧ��_��[���n�Y��RDԂ,u��~@$���	��|}�Ъ:��כv	'�����w�aE$�U���J��7�@�^8�����
�� 4�����7z��=���22�FY[�
~}�1��q��p��T�m������UI�Ε�3{�zJy�S��7]��z�����^��nA���n�϶Q:��us���)�{�S�"��~�˻ ����$N�:�<{Ϫ�Gp�
�]�`�@��U|O�~'e�I�F]��U(P����i^�s�K��t�n��Q��5�n�<���eL2�����h8���>���?/m��7j=~�F�S$&��t�\+38�}�?N[���ꯉ$�t��V�w��tq�����Py�pB�m�[��D�O�߳���0�׹c{�d���U H$�t����	�$M8`���������Cg��'vo��J?mh^~KӸ�6����Q);�eH��T
�l��>�ͨg}�5t̨A�*yv��٢�����&o��:���'�Rb!r"�29I쒫�c���n�!Ŗ�%�5�x�b^���[}������	M�=����$�{ٰQ$��~Hb/�パ����<�hP�?f��G�l3����s��Y2��(\ÞQb�( +��kh
����2$���X쬲Eޓ��ߒA)�:��An?$ �-����;��|>�>���)NȻOV����!�"��[���6-=��I�<�3g�&>y=k��ٝ��^��BG��k��P#j`���(�roU�:��8��	/Vm�(�� T���-�˗�x��}=(tk��iIN&���۲O�t�o�7����S4��yvրy7���o���˞�����<	���
,(U����6�j�u�.�pWk�'/��͉����������04��'?^�Ղ~'���۹~�=Y�B�=��B��M�  ���$�M6��Oz���}�{�e���Ĩ�ب  �����On��R��I�(���T��r���8p�}��Y#���$���x�eaE�1�@˟���h
�����h��`�ʞ,���ң�T�a IS�lY$��Т�b/u�<�5Tz�"+�׋Trs���ʔ�Px�T��/�%)θu�^���+l��n���]b~̙bĔ��4�\BL���q�່�N���&��u�� �nI_u�P$3��6����T����=3}w�����H;���9�˗08z�p(�Gn#��C�6`0=���x��;]m�+��0�յ���-A�4&T�#a��~���:{6�P�+����%xz�+k����9:�w�rD(���C�"�gFM�]��A'w�(�F��+�	�'G� ξ�ټ�H�1��2��N'�@��@| 3��sY�Cݱ�>�ݠ*����W�o���8\D�d���2��4�1g7�|3��߀�(�6� >k��w��v] +�=��@�wp�D�QĪ�,Y� Q�'�5dy��҉�w� A'.���ҐZzrwy�q��g�G�x��,/A����c��=.B=v$�E�������H��ཫU�ge�W�eͳ.�Uq�4И錗d��8�d6ـ��)}`ۜHe�9˳m���֋O:�h���]{c��^�	��8�ƭ]c�n�մB7Y��v^���W9{9��+�@�vv�;��vPN��h�[���y�q�\]ۮt�1�<���&�G>wm��h�#�7�;|���(�q�/��suv�M�Q�S��x}`+;d\�Gj��۷T�eS�v�`<��<=:��'p��u���֎��ۍ��,��1304�$�{Y�	1��i� ����Ĝ����?�}�e���{�Wz{�H�o��f�	�$H�n�㾿u� ���I=�}zC��D� :mh���� n�o��]գ�m��%+�HA�$@�Ҋ�]�(A?]�� |�hn��]��vW���&}�4��ˇ�� Cl��hʿ�Ozz��折Nͪ��y��K���A�{7ϼ��w%���f˔v��H��a.� \�]���=��5�;�+��Źph �I�/� >�͡�Aў��XG�;rW��{s�̇8յ�m���q�b��݈+�&F%A��y���J@�wǮ\�Hۿm� �~9��@�--��%�m|o��Iw����\ei1 �$��w0�w��K�9#<3�K>�V�nÄ�}�1ec��
űw��ӟyH���j�T3+4�]C=�Ѧχd�*dw6����^D�Y�Vx[(�oվ�����}�d�I�ނ�ɕ�]Wx�����̲PjF
��ݎ�f��?��͡�U�ɋ�Z���]@Py)�
 ��)+�$ � `iEEol�,���D��ٷ`���A;��ev�u\�A7ۻb�9�eF[FX:�{�	��4f3ޞK_��sZ�^}٠}@U��G�^P����h0��	)	���ݺv�۪旳wg���,e����6��?�ݿ!� f�p.v]�?�;`�I��A@q��*��y��	��n�'��i���J@��=r�A�{�����[&��B�sٿP ��>0��+zݛ�ڸ��
��
)����@�I�w�@$�o���:;e��UOU��"�_:�
o<�1���^`��nDQ���dӗ�V��o�VjV����W��y�}���|��gwX1צ|�2�|H��� ��J$p��%�a)݃��sn���	!��D�A����������Q9��+��4cT)�J*:�`�I�vm�V��H�P�y� =3h|>���^�L��Tc+�a%�"P2�D@bE�<�Aֶ&*����rZV���];�k��7����'6��m��A9��� �����Ҩ�]%���'	7��@դ��d8C�8d��s����͠�Ue_��}�x>&�:��'���,玅������ċ����|���>��#���u�P�I`������.�����}�O'�K�w*���@QNF6����^�e�H*^J��w/:��H>��kҟU$�W���ϳ�e>Q�;ڏf�{Z�gq\On:�k�Zeu�'s��|_�_#���v�H�Dk���q��ÝuW������P����ݍ��h��$�f���ikZ{��cQ;7hU@{�D���}���}��u��Io�κ-�l=7Z��\�n�&&��pk�2s�ړF�]<�&�M�>�w.H�,�=(�������`�~>��E��7���P �ח�d�GwbD��Q�їel��:��F<ؽ�a$�u��'ٽ�%;炊u�{��0�N'�&Y�8��9@�ۺ��H$맇QG}.��>�:�P$������ �;�����O �;�u�㖫W����_uAޝud�A���D��t�����V���˰l��}$$t}}r�'�[�~�uY�ED�-�H��TH$�����ߝ����$�	'��IO�HB���$�	%!$ I?�	!I��$�	'�`IO�IE�����$��	!I�xB���IO`IJBH@�p�$ I?���$�0$�	'���$��H@��B�� IN��$��1AY&SY?��٫ـ`P��3'� b#o��)%HE���""Q"EIu�B
%Q@��%%@IT�"��)ER�	*(� �R"�T �AP� }AW�t �:R�H
 )J (R�m@�$)%
 JQEu�
*��@(  �J�b� RT^�                                     �     �  #�}�)[�v�����.j�swm�94��/� 8��7!S���p����B��NE�m\ ���w�isP���@�>   ��|��V�g	� ;��\��e2nw��S�!�j���ڦ�n 7SM;n����y��m�8���9ؠ����҃��  �        =2��r��MR����T �X�P��5UL�to8����z7�x iJ)*fԽ2�5B���RJ��    ���W�ӈ�U!S��:U((�ӈ5O�y��`R�H���1�媀�� �
�0wU{hw�ĥ�HS��eiO;Q�4}�/�"�   �        :��R���U��>�UyjC�.m"� 5�Hdh�0(d�RE��` @��U@��A"�   1�!��Š
�� s����*)���T��fЪ+ ���&��� ��*�̀R�)I(��         � �ET�ʨ�mU����
�&�TX Y���YQ@��
I��^�� hP�k�l+{��bhH���� z <�r=�c��[ef� ��is�+W��-l����u�p ,����B\ڄ�V��*�.�B�h
H�
�  <         y��M�s����rƮf�FҜ�t֖8 85�N,�VT�й���.�c����p 9��ng:jU����j��A �  ݙ�t���v�#p 6�ж����5��vF�Yͪ��'.���� 9�+�ܱ�4�7-]%���n��6�r�J�����Pz	� "��L�R� 0�~	=U"S�� "{T���� 4 j���T��hL�i)��ʔ��z���}��_�1�Q�>�����,/<*1�O�f�[�$ I<�?g��IO �BC� IO��$ I?�	!H�������'��/��?����|������!�;�~dk�"|����y޼��?�C���z�3a�h6,ܢa�D��0� ���;��&�J-�&q����ӱZ��`��c*r�}q�!�.�K�hGu<�IX�����]i�8��MC4���eb�r�2�4iwO	�m��M|6m);�n/�,ʆG�*��[����)j�����'2�ǈㇴ�횅$!�-=2��u���웼ض��1G������"�"�A6�w�K��Uyo2���8,��^w@��JqX�)2�k��9b�R�
�lh��Ln�-���H��Gr���>�S�{l�T�-x��{5@v��Ȱ�s/b�%��H�����韜��2��^�y�6��]��32媪�� �W�#X��f1���h��ڮ����m�[�s�BgaO�V�E%�n;�35BM�c��v��۝��������&:v2��MP7Lqؐ���𖥡�ͯ�˓�������s��;;�gQ�Ov�n���4�w	x�O��x;�Lu$a�n��jo*
m�L.�b(7��v�Wn�����[��xz�$��qw��`U7�a��6Jr�W�f��Y�뉭�$���v5@�ݼ�s�d�] K�H��+�J��n�Er}��l_q��;ܓwd��D�-x��#�np5���RtE��,*�Zx���A	S��P�Ƣ�{��:�Y�ݽ�0��&0��xooH��������^d&GN	A����=����SXM��s��E���+c��3��A!ͦ���>���:w��x���g
\0	���˕���3��3�y�y����N=�O;~�y���yʍ��?6�C��y���Wq�6Z�/��T��͛�Áܝ��jDZ�Hx"zP�d�)�#w�����Ķ�a{�M9|;Y����V��<�a�đ��Q��x�E{{9\'h�A�|�vN�@�۪+��L��i�W�����BV8R��H���]��	}w�U[�8�A�Y&��]&�Ó�B�;���pN� �^����(Ϩ���"{��Y��|.!���7K��4�a`�����!���{;���KD�k�όx!��YP��Fǯ%t��@��/7D�K���W$J,w�;r����#�H,�:�Z��J��{��u�V�V铇�ႛ���ɖߜ�H���Jc��k�����/`�隞ܙ��<�-���㻰jN.�t���=�� �-˔u��HT���FMۧM֩�f�n�F����[ܟ^(7�:R�]�|�%�UN��8'n�P �Cm_ui��s���j���8�����0y W{��(w�Sx�e�J=�E�P_me�������X���C����qp��M����;���x��r�HE9�<����峕��(
S�<G�aqm!ڻ͈}�~�i��������"uۦ��S�D��g*on�_�5�m�,K�ѡM�&��G4�wX2�r������-�+��z�g#�"v�r�t7?ot5�aYM��]�g��fɯ���Zz�����"D�ðA��7]���.��+��<2��&^�+�W�%��lhq.7�C<vj�2��O�
yd ��+z/r�]���ro�ݰ+-�(�ۼ��-�Ol��;+��hR���	I�d�݀k��K��5D�k#4��Z9�q���s��E��{�rףd�ה��CO^
���B���\��sw��Jl���%�I&��~W)�M��9a�;�{�}=�-_^Zuˌ�Q�|��Bǉ�u���5k����h}c�so�vq���C�ʢ�ˉu�|����p˚3z�b9R�����󾔮�d{�X�l%���l�ѕ������4�����N
��5w�7~�E���&���VN�dBC݀S�����;�����=͔�~�;��"��(f��R������c�P��n0��y^S&i�����S8��,��Lj��@��]SY#;�gY4Dk���3|�jpH�97ۥeX�䶼��"xʺh�E�{^�������ޘK!��FJrݏr�����V�H8;$�g������a��T�����:fTVᙲ`������<�������(�
G�A�i�a�b]ݥ���m��v(�`�w�%�w�sÒ�8IP�����Z^��t`��C�_��:��Y�}T��l>�<5݋:#
IS��^�V�w��ԓT���Չޒ��f��7��<ccqٲvoC6+���Q��
�C��
��S���Z�안s'����]v�85����X�(a�ʎ�.0G�c�f���2q��x+�oF��p�i�w9Ó�f�vՔ�OmNP��Ƿ��뾛`�W{kWW3����Be�:[�xb��7��[������ZW�m4�Qi��N��QH��÷�y-�!#w #He���}�K���m4\�\�
vޝ��W`�{7�yҾ�C3f� &�e�A��k��V��v��.�9ٽ�yTi�#%�Ŧ�ޞ�o�,�Ǔ�;�[���D'1l��xIn��@Gٽ���<I9E[Ǌ�T��8nn�)�|�֨i��W��f=���]N��eA�P���t�-#�l��Hm��nEI��%���G��Xz���t*�JtR�ɹ1'hY��Å6�{˩ř�FYɭZ2��q�c߫4�-bʣk���(���₻5�������N.�����u��\tƧV�SD�16Wq��ۃMg��[�okDl�v����	�-ȗb#d�n�6���C�0�2�X����(��z�Ya�7��AJ��ו�]\xu�o޻m��F�x\�a[4��H�|oU�'k�n�$G"ݨ��ݼ/�� >ܛz���{��*b,޿��YSAk�qQ]������	�u���9S]/ C�M.�М��?{���[g/	zl7z\=vn��F݅
�,Μx��m �50��5eǫq3$d`Q6d�l�/�w���L�:���Z���>�����鸣�GT�X�h.�voa�m9m�veZ/<�Ւ��I��T�����!gm�+-w:����R�t���vȦ+���U��fn���v�2�ZR`� �A	xoe5���B=P�ۼ���Z"�kVM�wH����^��d7n1n>ʓ'w4G�1w!�e�@��(
٠w0��,����w,�hD}��.S�u�����f��m���ݛ���F��%�4�������X�����Oq��&R�Ӈm(�ߪ鷦]=ϋ�{��p+���8NM�����z��Y�s5gR{��V��=�)P��{�8�q�i�:�zj��P����Ch��=��p�GZ��d��`~8���y����ʝ�S�� ��
Sz�\����� ��
��f���M�ʪ�vp������fO_��V�t��s}�լ�$ܥ���7�\���t�ɥ�0���HQ�m�%F����3���4i�L������VP��"^�=ҙ~���>��س�k3��ܰ��;.o��s��u�М��T�Ҏx����z���+�
-p���Og'=ۭ�x#@�7��Dr�������F��{@8��d[�bqk���/z��w�>)=�',{N{���Ͳ����vα�%=����k�Ҷ�����i��]/�s�	΃�ƽ���xz_-y��'wN6I�)/��:���Ž|�ۺ�0K�k	9�,���*u���m(E~VW��h;踕7Q4��p:2t����,�D�������ÉW��G���#�{5���H�e�Z����ܞ�xp)�^����֏���־�[z�I; (����yI�	vb�F.0�{1��eJ	KV��H�t�a,�w�j�E��*FKxraOb�:w��ñ���䷏�ң�q��'����{�6�b�}�73�4������z�kpl����n´�l��R�S?��z�0�2�䝬���pظ�;��T��;�Q��C6U�n����w�r�6ٱ��E6�ǲc׫5�v7ņ�yT��X�Dk���|V&�<��2�15NrY���a��+U�n_�c�8���� X׽��P!%�g�������)��N���I1�k֐�`�`�$X�2�k�eZ%3c�)�Qٱ=���w*�%l���<�2���vI���eO��e�L'q��E�n3��[���םWp�34&�9SEȊ�s���.�?r<ٜ���,��w��ֶ�f6r�M��{��2�7��{�%����S�r��N�-�Nyu�{�yQ���N+���v���j�`�$#�x�{�g �I�F���Dt��,t���MEKHh67t�V��]=;��O��Wi.�������]��*��a���CyM��SW�d{�;�0Z{�����g`�D���֏p����ӭL��NO���o����/@�uEY��
E��>@FD�KYBg���/���;�(����S�e.��=}���-UUu��}�Z�Y
=�&�Tb0�uer�Lk�R;"�"g���}�<6�;}�������$K	]�)�?i�	�+�����yy��w�:~���o����%\��mM۴�J]���5�I����m{�����#��,����eNBR%��
�F����VǸ����<n�AHf���FˣۇF���)�d{��h/ꏽp�d|��U+��˩]�zb]���O��4T�B������֡W�]�V�x�� ��)��{L���s]�Y��:oh�<�e���!ۇyc�)_���X2_aT��}"*�}E+Xl����(��ov�Uk��g��3G,)*�nW�Iǃ>HL���|J��C"3X��������`�����1�M�V�{_9�kͱ�Bݏ�l��\7�c��
Rʓ�����e�)v�{_��u���x�N��]�.KV"�}}�$���D�/>|��É'�q�nl�%~F�m�E�m���ϫ�a3^˜BW��λ��JGf��o:Y��p8y�1=6(1xv�W���W*�w�]ec��i	�`1��q�j^����l2z�7D�8XS��;zk}���&�Z\�D���r��a�'>�ܞ8:�4BgU6p��2����.�ͣ�f���ۭ5�:��x�].��� �vr�R��ٰ-��r @͎"1��7���{���%@�mw�m��RB��{�^��5#Һ�h&wlDA;v`�6��7e��+�N��*�z�P��*=�ٶM^�hf�a��>�n�O�ÓD�.��Ԭ�LL�۷�7t��(��p2���Z��yj�л{Ok�P�+�݆��4�j]J��q`o2,N2y:�lފ駎�.~��9�&�\�ix#��9�	{���9D�n�א�i]Ֆ�1�s��L�n�o<�#���l�_���w����L@�~(>��{Ϙ�z�y�W9��'����]�w��	Tͥw>�y����]�H�12��%��������������ɲX颫,Sh�`����3��КA�FE`ܔ�	�3�=��i}�kg��q�Q���oB�fn����X��N{�Y�7%.RD�e��J�r��'w��0��*�	�=��Wj�*�Y V=B%�q=:�W��]N���Ǩ�ݘD�TЛ�;cE�e*��ɮ<6��n�l��*ΨF�u�g-�V���H���|1������*�;8*٫�5�;��q�F4Q-��yCv��I���� ;����Pcg!�A���s�^�h�Ty�Y�3�E5���7t㮗����S�`�{����FKؤ\�W�mj7]ڎp��]���b=j��l�
U ���]�9H�i�ۜ��ŽF��6tI��4t�X�8;��w���u��n0C��nɽ���0hd���6.aVt��u�pMU/�����1�x��1�>&�Ғ�yg�uoy�Y���sq���)������K;��>��.؎{�n����u����Y4/x`T�v�ۯ�-��-~�z[ͩ�¯�h���5Ne�A��*���(rx���@5�����@�J�s.h��b��cd	g��)N���Ω g���e��"��l��K�[����#���'7�����Ϧ.�������ؘ��*����҈����_,�]n=8f{��s���օJ�l�}����9�7�,RfZ���1����'C����p�ҝb'ʛ!��Z���I��@C�E����:�9츠3+Y&�?�y�CU���v m�=V* f�;R<М#���V�I!o=�9�z�?�<�JU���,�Y&]�{j�M>T�ѭ�/�U�9�o�oJI¨K�5oR���^�4#�^�3�3j�����ԏ�gf��Pl�`;wy-<�xl@6��IP���K�r�EvMj��S�١�JH|Uw�ʙ=�bE�7a�,�I�=����'�]'��͠Ȏ��a��)�zj[���6#[�Hk���G�zmyvQ���g-����
ǈD�o7h�:kƺ�s��G"������pzr���;r�10���:����$$�$R�Ha!!�$�
%d��RBE���d$`I
�@�d�P"�J�J�
�RAI�P��HV�B �$I!Y%d�� 
�T ,��@X  ) �BJ�)$ �B(T�H ���)!�E�,���
E	X@�d�� ,�"�H� � V�+ ��P��	d��"�
�T�"�Y$X(@YE�YP�I$a B�%B�@"� �
@	d��VI!@	+
�J�E��
��"�$	RE B,!$X@� �HTVHT�(�$ ���@�HH�BB��:ޟ�.��o�������������&�tCqk"m]|Gz���85!�p�3��d�?*�
*�Tl�`�hYbI8��1�]{�������)�{^��	X��1&�k<��5b$a
LP��E��{�xw��2�x�����'��]��&i��+(`ҩ�e�ј�;�Q3�:*��3��;RC��&��ײNkyQ1�g�<�l��#���^�ye�-y���5'�1
}wf��=�\�M5��3�!��wN]|�l{ڻ�zAـNx���Ǣ�ǰN n�:���������BF�3��'kwa�����f�� 4w0�:�	����
Λ�D�z�p�|���<��l������T:"�e�pM�:�����!�.^�dr�3�;���f,��XV~�=������h�G<�1�� �o��P�n^|)���C6`��3�n��ď2����7(��r�NF�]��B:YѦ�<��e5K���QS�� /x�ʽ��E�	�\-L�h�m�����TȒuz���pI��Z��z�X"o�q���~o����7�4�6�M�P�'��sy;9{Gf�����Ǌ���<����G
L�����zKoĆ=hww�o��P8����E�-S��{���k2��s�@Gm�����g"MDr���N�՗��ǎE�}Iw_������B<�ұ[Àö����y����Y}8�y�g��.�+Sc�{��;�׊%k�0Nl�lX�N�)�jU3E��	�n�$h�O5�p-��L�)6hpX}��3{\V���^��B���H�z��N�'���69N{�ǚv��'Eg�ۤw��z����M����J���Kl�"E�_m
����}�x[�А�.�w�	���iÌi���y�����{'����n�E۝��f՚HЄ�ى��7q�0d����gM�i�F�h��Ϭ��d%B���ú�?�4�~��,��J�I`�(���[$B���8T��R`<{#����	����O��|�X;$��bf�9�nn<��,Dq��a��^o�������.7�=�=	y!�zv��?��~c�� �{��Y��ÙZ�B�%n"�M���A�BM^K8W�Sa�k��[�D�����ޯ��ow� 5i�u�]�o�|�z�	D���g��l��s[|��k>^m;�V�475ķO�Z��S��Ŭ�r�D�8<�gyIf^Ri�jz�:8==�ۜ;��]�DC�p��79�h��l�F�dָ1f	�Y�M��On{p�ÔCH˹�jR�N�h�9�N�1Il��m��R���f1��,����{i��-~��Þ/G7��~�sʮuWk\���X-�Lܾ��+�{���ݧ�b�]���mk�2�\p�Y��}���񩀣%��[�X�3r֮۫�'�*)�x��<1We[u�1��w"MZ/(a����X���X�w��+/�®�,|F-�TOx%�d~M��|�r�a��k��ʠ{J�/��������۝@^'���ogG�C�U)�O������w
(>�A�w����F�}7C�
�O��[���F���LV�%O�����Y�b���M�m9w�K�-��������$��=�w��']���݋��[&馌þ{�U�$|�\�Z֏�=�:�-/Y�1�g�v��w�C$Mf���Ӏ�X���?�ӽW`���c�U{bO�ԃ`M�*����<3�vo�(�E|OtN��g�
U'��:�xg�2N%τ�U{���};M�� 5��h�"�]	�����6�;0��Y�F,������F�^���'��	-��Ȯ�=�C ���z�p���p:K�� ����{w��m�%X�"�$F�ƵI^ĺl�=�`�[\�:�^_y{�Z���mLd'�g�q�:�,��+� L���5u��:xe���2Ӳ�* 1Le���U*��c��4F) �0�WI0�l�ѴQ���\�&���Έ�ќ����\A�P���Y�2�9��A�f�{+,:�ډy_`����Ge�ג�;]�=g8��3د,Q�މ��坛7UY���wpǀo29�s/�
I�\��t)����~�b�s\��SW�p�w�2+�^_W�q�ޞ��9�q�N,�(�9����t����o|භa���ܞq�k:zbg#�G9tx�;��{���s'C�)}=�S쉸�mcҢXײ ���ES�����۾�vs�����rD�w����s�{�U=r�Y8�|��$;۸�Ա{V�����*�n�;�u������v0���M(ۼz������1���3ހށ"g�^�ޭ/�{`����hin��V�z���פ����������9k��oh� ��Ky�c>�iӇ����W���)�`�!鑬�M����e��Y�2�瞔|�g �h�_�w�2x���${�<P��-�Ak���t���o��V��1T��t�&um��X�q�`�N'�E�����G���&y���]�l;��\;�������72�����bC����I��d|����v���A����[��8�Q;��7(oqb@�U�^&*���j�kz��FS���'���U�;M���;^��UD�4lĆ���˧v�i�7Ow|^��x���9�a���>I�InW|@Y���"x���bܳ��w�hsV~v�Q����g?5�=c�%�l���+|��ǫ�a�.�V�c���(��i��207��W����jf���{�.�c\�6��s^^J늍&�o.!��&��D��iZ�������6%��,�cY=�5�r�����Y�33M��R�j,J��
�At�n&V�E�q�`kc7S����^l�8�.�^��ܘ���DW��zL0<��AK<��M��ꍑ�Sf�N�9�cj0�B7c3v���{M��^ַYu#87!��p��SC4�o{oYw�6��9�*�=��X�Oפ�O�]m�v�1�.�����7Y�j>9S厱���o=���^�{#M��ڙ.�kS�8qЄZ��6����x���'V9B��Əe��FySva������'GB;Ԗ�W�����q�56��Q+L5C+CC����~�XC�4��7\M���p��Z�X��$�F���}�I��4{�j�	jɝae����_3d��*B\�x/{�:�M��3V���j��F�l�{
��q�J�X��q~YrͶ���hkvfY<yAx�e��iZ|g���[��ˎ�DC#[V� ��8��wZz]U��1aӡ�?������xgC,-�BJ�¨t�N���c4ȿ1tٱ�����6�v�I;�}���f������lB
��ؘ�^|q]קޢ?'#��r>���{�W7�7Ó�����u{:Ǿ��H�@�����/?j:���&u��aJfZ�j���2\;��.�g��4K�//i=�\=L��r7�{��6�q7�% �յ�t�=70��ʕ�H�b�T���
�W�;�u@'q=��AQˊ��=p�^�y��s�ս��{��~�|:x�ʣ^�A��=��,6�oӡNFCA%��@��i�G���^��2�_f��ȗ���ι�����#�ΐ0�S��OMۇ��oh�����'YIf�&j�'M
g+����X��62F��.ŷ��g3��BQ����fw)����L�(юk����Y<�{rՄ<	&�O��J�gh�O�����&�6bn�×��\ļ����7Lŵ��%���3ӱs���+1�"����U��M�x�hN�순/q�tV���6{�����l=+}fM>uv7OQ���V�)�9�̼��5�v�k]7AD��l8ܛsP]��8��B����5P0��Y��>�_{۫��-:"9&sةP/k�P׌�I̷�1�r�N��7X��]��`i� m��{��{'/A�����>V�s��5w|���Ț���H���'���I��Z�/h?�<-=��a�湼��
t�Q&޺�w���o	�Yd/��޾��9)B�m��Ŀ.��8��w���#�(��u����j�/��1de	���ag7 5~��~��f�6A�f1#�g���uQ���{q��y���?"*�W��;��3�A�:�aI�b�����{�T6��%�r�#�[�c�Ie�5��F����۷�;\��G��B�\�ϋ��ʞ�̝�S�uLNѠ�^<��Ъ��c��e����q�4����V�~�-E?E�^�\}�B��}W����xZ�݈p�m�.�V�5���w�M�x��Z��B�x�g�W|��y�W���s%�}�~\��،j����;Ȱk(M�Ab/<Dɫqr�՝n��-#��]�_U�XZ��vy����\k��xK9�>K��S�wݯ�Bh�˻=�'�y�N-'��Ȗ�K�X��*�P����9&'6�N�u�<��q#�mþ=ݞ9D��}Ǥ��ӛ����N.ECbr�1�P,���.���/����͛�B�Ǎy�t-��`��uI�VZ+eeн��:'lnj�2�nN��Īn�غ����{����Yp+��E�R���9��~�?JGNC�dV&zF����ی���{��mGDg�% i�IYE��?D5{���'��(��
(3��S���9���v�xE+�x�8�L�w=�E^Z�
�0���P��I�<mp9�Ǜ6�X�yਾ�K�)�[��{{ވ�OjM�/Fc�&a�v��Y��wJ�h�q�jW&!֚	��4po7�����{��������Fn���Re�*\d�q�80	�Ic{�#ѽQ�a��]Ịx���	2j�X�`3؁�:�������@g�����\:�k�{ۚ���7�b�ڳ܈J��9�T��{��O���c^��^����3��=�r�w��j{Q�u�ۏ��������jZ�ʵն�gv-x)]������L����U���xF��Cjՠ�!R�}(��Q�^y�CWw�������*�6�Ǔ;�����O%��|G�ܗ�f�fߢ�P�	�Dm�r6�X�e�4(`x����V`@C����V�<;����g���Rh������m�/�	�;k�e�������~�<���b��z;N�I���.���U��^T����(&��!�w{��
�_ۉF�q^��0M��ews]~��&Jx{�^�a��%�g�rɮ/L�{ ���mꖹ��ky/ew�S�F������E]ƫ��ږ�;��C����-�G��q	�����sV�z����p�cԏ1n�����-���<|9^�6�ŧ�/��x�ףsQ:7�X;��5�j��>����9��/�!w������!�C9�{�`��p��sޕ���r�|2|��=+[Fع8��a=1o�Y�x;�m�X���h��8F��Nb]��ۻ{}&�'=W�k} �Zў���EŻ��b���F�v��y(�ɫ��5+J�P��;����1��I7�z�&s�ofm��'�r�X�\�F�E�kc<,��ѻ�R��}��/�YwVSz�׹���~ۡ��`�{�y5�r�Yf(�b��-B�^��vuG���n�=��@�����~֎6�����;�:bJ��\�b���cpmM-ԱH4�ʫ�Tc/T���ɛ�zj��v��7|�w�t���Op����7�Ť+������zO�	l�#��Ƹj��$��q���uM>�O���i��%'�ŉ'�O	p,6W���}�U��1�'�gs^���Y��C����-���$ݹg]����@�ǆ�w�\��־�nF£9���.K]Ӻ}�O��Fyw܏{w�5�R�V��>!rZd����9q��&lf��B��B�F��{��L䡕3)lRy�i�K\D��!eo�� �a�ÑZ�هn�D�K��%���"��������B�z����vU���f��Ž��Ns�a�p���C�띂-���F�=����ٯ�8Fm%�V��i�^1��XUnM�����~�B0у[��f�M��;e{��}f��tC�v��L@aԌ���i+����w3wZ&�!x٢�^V��h��2N�q�ʩ��ƥ:XW�I��`�?{w{.���;;v�e7��_��1MMJ8����X7l��	i�}�v���8����+w�zZ.�\;ˠ}�c��σ
��:&�����͋ͱ�j��5"�e8��?]^œ�~��[ ��f����xrn����ӃMPg�X{^+��7���<�}�5l��wk�zuӋ�Lk��8/�"�%{�����F�Ӯe�i��f�d�����'0��ِK:d��k	�tb���f��x0���I��:ƽ�����V��Z�v�Ci�uo�;d����6��}כx�%y' ��VOk^Tf�i�;gd{���o��1�r��ؽ۾8�����7e����>]����h1��HW^��7�w�xvr�=y�v����8�4[.�V�vݩq�u�V�;���?�y{�~S�����mؚ��g����N�7���]�=���@>eh��
�mo��I<gAک��}�O{�U��K��O�y9��^�x��,��C����Pީ��V�6m~h�0�K+T=�KA��t4M8[j(l8\�E�U�>������'�Frx�.��ND�Kf�뽕�����S��[��8��ȇit�����Y0e]��38+n�mI�Ig���WA׽ix��K�_.�g4z��>8���w:���0�ق"�2�A��)�h���2���/3� ��{F�=��{o�}��<��mT?Ttz~�+;�;;|3Ss�x�g��8�Vg��-�<���;��,UZ�+�".v�h�����$�$�|o���<1�||�/��p`����������ۮ�ݛ�q�	֬��f5��ٻt!�����=���8�ݜe��8n��d��g<�z�N�+%���O#G2M�VXӧ��F.� �7Om�[kpH<��nh�J����Sxi��n�������U�ގ9�N�v�ݞ���\�8m�u�.P8ެ[��]��]�n:���-���'b�7u���d�|�����G��p`3���g2��p��v�n��okv�1cm�L�ٞ`6w=��I\�v�WG;Vlcj��N�4��WWO(�IBgpg��e��O]���Z�R�2X�۰ݪ��������`uq�uǻۋ��n�Y;]k�1��WnN�$㮎��܎{t�y{i�cn;v��p�ۆ�n%3[��T���TH�+�`�@�w\���un�&Pⷳպ2���і�v���c{7Y��zty(�s�<s��&ݬ۔��u y�<��q:��(q��ԥ�0s˲�[K'4om���V��z;V�o8��x�k���[ۃk�.R��l����j�f���H��N�9�kEC����ꝧ�nz�᭸l����v�nw)���Wg	۷F�x(�=��̼'OlG2��jw/&�����<8�"l�;71ņ��8w<�۶E7f�co=�0�ɸ��޸�}:c��ufx�X7'pv+��:�yn;���a�N]kz'b\<���k�m=�8D9��s��S��{ J�r8{u&Q!M�L�M����ۀ�m[��k]ny�.}2����n�	�n���"�w��%|xm���`��y�m:�tkc��nm�xp����m�۶wF�'�c�N�m�]�n��F�]��N���m\�V�9�!{gux�p�5�q<Y��qOm�p�E��K-��ۧ��nܣ⎷m�{�&5غ]t=]9�Y����N���s@v��xq�]ZD�v�ń����kۄ����s�\��.w@� �l�����;.(���'B�u<�kh�ӵ�rg���q����"k-�lG:�3�1C�KH<cНn�n8���@�8[��M�LF5��Tv��d.y���\�¤��Z9����4f�+[s;uH�e�N�;v.����4;n�M٨.�q�w18\V�أ�\���vvu���t���'�^Ĉ+B^�ݮ�E���%�n1Q\��8�FH�#��+n[y٤5(��&!�kW����U�p���)y29��tv�ts��z�犱�n�e���Qm{3�l��4�n8y�h���V�#Z�4A�מL�X	W`]��*�G��1�s�90��<�v�v�T.���v��<�]���붺��Oq�{v�=��[�������pd��'�N+������
=sOnR�����,�7���p��^�����q���@'6����9��3���g�����C�ۛf���Ϝc��.���j�5xg�ѻ\��xL;mf1��nwn6����v��w��v�v|AS�w�Nz�vW��"{`6�v���<u�;{	��-�����Y���]�3�^W�=nM�ׄxس���ճ��bۓ��5�:��k��u=Ѹ��1��M��nK�u<����ks���
Z��|��m�l��{>�Pyt[<[�A��im�kkL��l�8E���]ۮ����C�R��%��
	x�ռf#�"F�kp+[��.�7���:��}�E���9�<�79a�:��Q����:<�g������^��&����m�[�
�7=��\�Un[x��.��ܐng��q6�y�b`��{U����ͣ�eݍq%ѝ�����ۭ�k��]{\e#�;Z��i�d�sF��xk�V���'r{n��9�h�Zt��g��=F��\��kf���s]��; P�̹v8��;�v�\�tt%B]��Z���m��@�G5�*'�zN�`"�Ɏ9�K��y��`��*!�u������n�^�F����g4�\�7!�s�wc^�v�y��8s�s�#Z]�k9�p�um���Y^��+��V�K�ݔ{D]�x.�����<u���I'n�i"sۅ+k4���mR�z��<�ӌu�*\V�nAu�ʉ2\���+n۳�X�,�̝O$T�pq���{1��x�0��{g��z���Xꣶ�Q{1rWC�*뇞�a�Ɏ0v)�m�q��{�Xx�W\�gp�n�[[+�譻r�x��
9����3ӼpTN-mWn,�8��3vw/BUY7Y\�<t�sr���s[Fy�iц���잖����y��C܋iS��zϩX�v�cn�g�oW�3۱�nm�{n;6V�U��qqv��xc���F�:�c��9��Շڌ����a��b���/9g��ut����"��[68Eu��1�ӂ-gyRp�ۆ:X��� ڻr��\���ݼ��C>��q�rj�#78�u��prk(�;mJ�]`����]��{�u���r�6��pIH�gz !��qػ��q�
p&ݳqΗnî=�N��D�i���0k��8u"�scv�b����m�|�p%H<-�Q��ː�� �)8�q�\�4A�/)>]os�{X;i����u�2uyΎ�;1ۗ���=���ۃ+���J�c�����q4`��y�q]S��7=N��n��E�n�j�C��Ր;��vm�q�,��_V�k�n���Ǣ{uM��#5�Bt�b������D����d��cEu
�����qX�y璲�&�}h\��ch����S/8;�n���nr�l��ľnݽt����'D]�ŀ�cV�Ƕݎ�%g�2��s�Ln�u�$��A����ӌ���qu�����N%4.�D�Y�v仏&rv�N)޽�:�ղ�e�R���=nxp�\VKG;n]��uv����,��ɗmF�W��=�\�����A��&x�z�X�Q��*�F9�>.I��{��s�N��L�u�q�Z������\���[�vl�Kq����Z8J2 ����䗞`���f�l�r֝hO��mqf8�; ��=v��t]n�D��>�#�}�m�sue{n5uj�5�s�&ۇ${�8��k�<=�7
��a���l�g�l�����Q���L�]u���7�7o7bz�����B�1��^Nxp���I���!�ptun��7EE�
���۶��c���0n:�t�l<�.ڝ	�y���q�f���; m�5G^7g���Ccp㍱��������vE�҈S�dq�E�.�RÎ9���}�B�����.K�[����f�̃�2�^��{2��kĝ����6ss�ݛ�

\�S�+��#�;����@ls�=�m���ssźS���Qk9,&��&����m��q�WR�:��Lv^����V��յ�/Q=��vS�zui�^�8�p;`瑮�4��;tgPb_nAOn����2єz�aۮ ��=�gǎf��N��ռ��mup6��!�I�ۮ8��[u*�=���Bnm�۝�]��;��N�t=k��s����1q����ˁ�n'Fv|��EZ�M���M�\�j�rpv9v�݉�ʇ�3d�o\,&8�4��ں���ݴ�%(\Y㓸��lw<�ǎ�m��3��d�{b{rGG%Z���lQx�0�<�kghgU�%��ۄ���,;�9	�qa'=�d����mu� u�u���F��rrn�����1�͍e�9⤑9�-���sK�G0�=N���g��kOg����.�������9`^����7���Z=��{rvn�,�\���<�zݰ��ƲV��-Ǟ��P#�n3\�<v�v�4Y�B�{v��q�9�_H󎬻�h'�r��\�\l`�����+����[�;T�{uݢ��s�ŷ�wc�]&�P�:\�+�G�uN�^rm�v�u�P<D;���3���	,�oWn�	�����q�����.���ov���9�$Zs�E��8{�����Ǣ�;v��km�;]zͷ\��:��ǰ��v��-�ZK���]�w�Þ�qۋcM�t�mZ�K�r��H�Ư+��جƔ�]y���w�q'նw� ;r��a��ݷk[v����d����m�#H�s�̦8Ը\p��硡<�TWwh��۱��Gn���&���v��J��ѹ7k��:q��gI�덶��홎��b�\����l�d���0u��s��u������.��n;tErl�����t�vq�5�6\��q�;��n���<�g5������yC�z�q�6�M�/;Y�1s��ֲl�-鮝9��$*f3�>ϙƝVf�&�nY�#^;r�ֱ�����Z8۞�$Ȼ�kk���N���y�q���l�٧t@�v{B]qj�&�P���msn�=�����u����b6��{k��g�<Qd�m@�U"�nW'8	��%�c��6M�SI��N	�Cγ�q5�Kgթ�r༗\�۫�������ŗ�۳x0��d�����9�W$u����&�� d�\p�$ZtZ�΃��WF����>^M�ˇ�lb���笽k+��5�Vl�ٮ��k\f����MȀY9һX�#l�F�k�U���'�\[fܙ��ҡ*�΀c�����n$�&m�vh��c�XͰpk;�O4K��֑��匽���O��v��1�ش80֍�,\<��ۣn�<�y�Qr�a{;��F�(\�95I�8�{vٰ)׌޴<��[���m�՜�m�g(�Ӛ�3��n�FP���:�{y9ր9�glǞs��L����Gm�{V�i;��Ѻs��q�b�u7;yx1մ]�����#x�4ν���٘饭���Es�k\QE�ţs*u��k�nLV��=;nguƸ��\��Vvu!��M��=r���c5ٯݽ��m��֣V%����4���m�l����6Ƭ���.R�(�ir�̶Ա��%ih�c��V.R�2����\��f51�UPJ�l���R�l�B�����ZRڕ�,�Үa�5����Qe**ʖ"��m���؉m�F����JEQT�Z5-*f8�Ȣڅ�JҊ��mP����m�j�2�,l�m��UF��km�(6����F�mUĘ�X����PV�Ѵ���ը�,��V۔�L�����E�6Ҋ�т�DJ�kE--e�e�Zڲ�-Kc��ʴJ�V��IQ`�Q�9��l�%��V՘�E\�Ue�֔lVض��T+j�J���JZXQ�Ah�Ue-���,qH����ZKD[K[,�E�5��­L�\�����Z���ZS0�,�)DT��*ڕ�mJYTQiJ4EX�[j,Eijʭ�jեKlh���am(�1���j*����{���7G�s��ocr�E��
m��]�t�w�;O���]��8�����K'�y��.�%��\�f�ܚ�Y3u�{A6���k3��s�;N1��݌հ�Yy8J� 퍪ܘ��֣y7[pjyۃ�S�Cn���ƪk�{�뇏nk��uv-g�Hw�v��(ܻ�����"]�݃Gc�SK��-����W3��K���մ���1Ѽ�v}f[�G��K�F�1�����,�c�v��۞�EN#q�n@Mq�q�u���n���h�ZN��u�z$	H��L��m&��$��c�Э��}z�<ñ�[�r"s�9�z�'�sv��x�ق�0!��ꗡn��麺��:�P�i�e�U��u\G�Iͷ;��z��§;��������b��7H�rpnh�˷*&U�.6���JX��[n����Ò:��t����vM&|t�î�vmv7歿?7\���5ь�ixމ^���r�6��dѴԖ�糁);8�97Z�knJb鞻t�g=<�g�q����Xl$+�;\�bq�H�	b���n�N5��.�ឋrbz�\�ã͢�u r^:8��u����ƣm��p�3=9�:�<�u��;�K�Ŷ�nw<��[��t=:x�)\Ӻ�`�k��ZGq��{TFpN���Yy�.;k�urہ�����4�mVs���[N+A�n�h�윏k2���Zf�����J�8�%����%�ۜO��
�Fp�lo*bWX�6�&��mv����\�*���4=Z}��aݹ}�w<(�bg:�mf���u����v���z��W��4ny��rRpR�!9��ێ�Rnb����1tNj�v�����Km�pm��n��G&۶0H���g�� qgsX-vݒЁ�X��ݣ�ϻPE��nG݋�Ѷ9ݯ&�W��SWn�\���]�U�۰�f���f��{����yr��L­\�k�+A��;x���l����Ȧ�����8��7v�r�������=�\�a��`콶\T��L���ʗL���<gl'����0��#n�
�9�TRˈbۃh6��QKU���0ƍ�f�h��<&Cl.πC���9.��'9;�C���p�U9q��+ɇ�'���@�G����m��d<��޷��>�S�YtDV��	���<�D�����d��O�y_�!�Ʈ&��[NC�7�2[����"��[��y�=��� v�q� nNc��բs���yo|����'�cw�$bʘQSB%��������A�DNWNź�\zj��� ��̀�9���@�a��Zy�����X�����4�w�� ���}�9�Z ���x��j&o�go�J��z�,�KK�1��;�����o��v�[�!�pfTR;��`|�砒moo<�b��T�Q��Y�!C�&$D�gm��vۧ[�n.qܔq�qv��;�Ʒ�,)G���ILD�(-9��IcW�2 ��z�M��I��1dW����!������K׾�����5���{�/0bA(ʲt���s�׸7���ں�]��F��n^{�͛��_�&��}��/�0Ne���P&�nc����\Ow�oǇ¦�6�ㇿ�Щ�R�=��H���b�vM�� _gmڲ�2��h����u����1
�h�D�g��mQ ���v [�K��:�a��@fM� ��3�I�fR"��`(�]Gfr��+�}�V��D{=� �@}���v�@#6����w[Vz-�wSc����UTR�����^� oOsB/+w��uB�a$"�v�$����=���3k�ls���:	�3'>��L���
k�ZxŎ�:��m�x9���4u�<���:��&���)�&L�1'O�P�����n��@l�aJU����A�g�[uճ֬$J����Hm�6H�"`ē2���7�X��jd����9�5 fv���͞������E�]k*���ٕ!uAE
j)��=ۗw`���r�s2'8���쉟b�Uvjz1�/`X�l�V�hO5��N亇��.V���'*������_�wDx]�!o)��W@�����"|}���2� ��n"�3g�i�Z�XIK m����w�]>�π4ߋx��׊��z{O0n]c&�O�_*���[���M�]�4�L�D��%MJ%�籩b��y�;t�{y��U �{;n��>ݞ�� �.��	~T���ѓ�nc	&Bl�Õ�4�Ɲ�7S�
��n<g�J�s�mz�F��?L|�*��$��^�.�_Y|��� �ܝ�N�����e��&�m�Ey$���d'4��	ic����C��"I�p{U7��^�z�nՑ�v��>�N�&Ҍ�¢�Os�b]e�H�"`�2��t�h ����Ey��Wz9�U{3@@#����r��{�����5D��˹S���GL���� A�;�K @}�u� /��Y���|���hۗ����RQ*{k7isz�TEmz噆�mV#e�s_G>��(rc��߽�'�ޡ�m�^X �u��u�k M������6�> 73�ڳ���*���N���]׸m �	wM�� ^�mڳ�eݺ/��*e<6E1�
>�DL!ڞ7'�
�֫3x`:�;;>����ɣG������aQ5(�pk��. �7K�5@ 
�;n�^tߥ&���t�}M�2�c���h6D��A0�w��Ph���k�S~��k�Zy7�X�;n�˯V����{g�*��Lh�~�}~�z\���3:fɩ;|�$��3n-"R��y�īI�#d��&�V��*��������ڈ�5��|nv��$���W�+/��<Ǥ��ۆ�,%O�$��*hS40��m����\ײZ~R�o�o��3�v�Y-sܨ�JLӋ���r�n�Ԩ�9���՝�5��uv6��-jm�4�L!�-T���7��mv��R>�4(��>�)OvB��q^�ř��Q	�O����ch'n��az��8���8�k�9xx�����I��-��۝�厡�8�)Ț:�z�0g�8�<��'6��mƤ���a�wk���n}�h��ۮI#�/	lY9���-ד�<���ۭۄ}=g��:��x�n;;��n�ۿ�_��ߘy��c��s�����C��s��]�n�p�z�zz8���`V�NKD���t����k7������y3:�w@z4tvn���f�&�DMUI?MdV~�� 73�ڰH��6���_�2�]����٩���ӡ#��m��x��P*E}DԢ[s��:{}��7�|u��Dyۙ�H��;��h�%W��lu�i=U��B��	T��2���f��k�3$����Z	/��;[Q��c2	%���3� ��6x��PTJ�Q5:�k]��.�P���v� �῀�;�L[�{����4��1�ye��3�L3Ra*�αJ	g����z�{D����~��.~$}�ܬZ(%ڳj	�!]]":"��[D���qu	�wn��^8��2h��\A�=��G�l�`�}���E�q&KC;�;��nՇ�l�h �/=,4�x������י�j�ή�ѭs�*�S�E~OC���5'��*�v������>4�/,Gŝ�K|����w���n�\^pܒ�:�Kݯ�؄
�<|�Z�p�'�ns����N�g� �����o�06���>!�}{��~��zw�`���7�I�O��� ����T ��MG�G�c���n�p� _M��v��A�2���f���v���R^?tv$|�8�iy�`�o�o���q�Q?�NƘ/[�
�)R�"����ǵ�?�o�]�f�����@nWh�n���H�}�v����o���v�o��q-R����l�@F$we[�Q�u��:�n�P&�6W���~}߽���y�
�`���7�\A�n�t׷�m���s�2e[�:�Or�@;��7P4)�
�M�{�.�}`������U��>��=� ݛ�,�/���E�n׵�՞3=wǩ�����R�x�M��'���2�z\��1c�y�o6y��z��.cM�2b(���Dg��{���S���yZ!�8����ʳ4�Ec�j����N�h��Z��q�7��VpH���ݸ�H0߯޷2���;�0C�� ��݆��\J)�D:/<� H���	�A7=��ܽ&1EХ��OM������N���7�C���X) oOq�W�U��Ԁ�Os�/o��Y���?���Bº.�B�9��x���Q��JF�y5d��=g���nN����� �S����$dH�F&F���@� ��GSEF���E^WG�\��盖�@׻v��"�RB��U01��KxS�b����٣��@Ǜ�q��v���>���<�v�	�{�}��]@T�"%)�,μ�ш�[��%$�[��U�}v6���^x�	���DE���?�m�򲨩�MQ3��f��z�lkެ��Q��Pz��  ݮ� �X��M(���+.�wЩ�q�٢��S�P�e�\�CxͧӸ�s�/"���Q���^ʳ�59=$��l�����:�ZqT�Sv�&Z��䗓�{����߰2C���=��ي p���R)�����:�3������=�
�3�W�/�r��؆�4��^�����=��9s���Ѭ��b���x�*9o~��SEE)�������ۻ�7���. H��<��S��;drV�y9���D�����HPS�R�&��bdY�|�n��7��z{e��3��z�X@���� _fW������c��_��`���raI1E!���]s�`��^h1���N�1��r�$�r�Z+�,�ڳi!x��)Je�H���r=�H�=��	��O�'f�ǘ��8ho{^k�<��f�{�1��e��VU|MQ3�ךF��ly��N�>���������6 ^fy�@ __mڳ���+�.��Lm��Rb�!}:{��UX�{����W�����znt��n>�7)1
��.��m�P�G��4LZ�V��A��<>YRШ�"7�m�XV�-�;d��7���aݬ�\�ӄ8;�t��s�i����z'�Y!l���wN�-��s�Z;����yL\nA��N�������:��qn;Z�{��q��I�Y���Z�T�@����t
r�<�s����XoY6�<;q�v���Y�\�93�iӷ	�=��էs��8��Z3I�]���	F�;mA�g	=�����7Q�]n�|�n���![ƌ!v[�ۿ~�;ADҘ��)�A�k���$J��0�$�,Ƀڢ/����4I9�{`�������2������z���j���흯Z��Xƀ���n� �����8�������}��E�I��ߪ�I�_zZNA��"���ܳ�Tz# Y�X�@"��n��ęR)"�&(�xa��6>����G����$��݀Fo{��zg�k�"@���2!��W��SD���țG�r�� H7z�����������Y�5/���>H�۵d7��d3�t}�O�L��s9��~Eh!��'��V|ԯ�W����tg��{.�/;a�q�;M�vW���r�
���g鬌�鈎��n/� Y�����d�5�}["Μ�-A�;/��Z���QAJiHMIM����Z	9����#Wml+""���N��an2��ҕO�l��Ƿ���H��������	�)�ⷡ�&�A�O=ӽyb�g��桎���
m��7u?8�jw�{��@ ��������i� #]��{����Ā��p��*�E)�NF߻������� ��;8p�Z�j9"R׍�I���J����L"�bw��'>�]��<�n-�����{7�}ќ)ږC��INs8�"��$[�[2)"�&(�1���� �/<�]�v��'�]�篮� �F�{��@�mA:��A���7�<.��QP�(&��=n�۔#X�sɇ�3��H��0�$N.��?v5l�MSS"qY��X w����+ټr�(�ݧL�[�V@�3���	u�y\�W�QU?�|m�(>�.F֢���\k�++پ��Ȁ��C`$�祠*��oe�M�{�r��>���`d��0�&˓0�O�40 �/<��il[�ݿ{WUώڵ>{�I���旰I�|�z���+�3f'�wޥG;�%�ZΑ42�nx�o5��Wlf]�'�o��;3������M>;���1%�8;f��P�35�;%����e���j9��{;^q��`���Ć��}c|'M�+=����#=�n��R*M��B��ʌ{%�=iq&���ܦx�5�}���G[�S^�yb��v^֪;�wo�{fvo��ɫ���}�7�N����x���l���b@�q��h*i�(M��fb<h� �zt��TN\U��+�j^v~��C��Gj�P^�n?z�zv��=��N��*B(߬��V��^ۋFx���<^�zY�F��p�Њg�4�W���R�}�ad95���i*�kn,��7�3��w�M�A𺙉ׇr�H.ز��݅�Y~]ֱ]��G'({eo�ta��������ye�\{���6��y��mն9�y7�vF�2"v�e&\Su
،�D�i7�~��V�������3���2w���Óh���.1{1��l����un���x��>"��OX��s|�`1�{��S;%����uKG��_�ϛ�9{�9��돽�8�����0�gOZ��7�g,�>���v����(*�YR#b�-b�A�W��A%�&7�m{��a�?��C�u��b*��S��.�� IE��p^� S�9Uf�U���6�T��bhm�N��l۬5�k):3E㛅���զ���Soc���xٌ��W�D�)'B��&cMpxҪ�[��3z,la޼.���ʭ-�[j����0�`"/��5����[e�XԪ%-m%UDq.V�U�X�-��J�l�����m���Q-��Z��F�6�31majP���[D��j��[B���F�(�-�V�Ds.��Rն"V�m.8�F��X�h�EJ(�b�)Z��)Um�ˆQKZKh�l��*�#e
0�«+KL��,��qm������ER�Tk,eն��-*��AcT������klF����E��[J��6���Җ��QmY[R��h�4�m�KJԴ��m��-��E���mF��KE"���kcl(��R�cj����kaF�UډDTmmZR��(���J�е�Z����,Q��R���)Ukj�"ִVX�TQ��X[K(�U"5���Z�6�R�FYhі�ƪ��Pc*-�id����Ɩ��h�"��)K[J%��UQmh-���#J)m-E[E����D��(���Q����QF�ʍ�Z�-cVZ5EmKE��D$Q)!F����%���i/c�ۈOLߑ-���e��h��~��29�=�� 1�[C�fM�����9��E��I6�c���c�7iS1\eDȅ �BR�ڮX�ĢPK;�=��;̬���K��d6� +�r�� ^߽o�U��{$fw�Ǹ��[E,e��m���L{q��Δ�>�.�ۓ��5����ȓ��߿_�=(�IE#N�=�[h�皠s�'�������Ѵc:x�Z($s�W���߸nT�-2�i�rL;���V�B��oλ>�iy�h {��Y {�#}��w�:/�7��E}T����=��j� �s;]�` ?tKE��E.�3gq=��r�;��S�'	�����z} d��cC��A��*�3���u�A�c��K�$���I��́j6�f�1�McM�^RS�����9� �sY��U(�ՠ�/)##_��NÙ��Am뗸���W>��S�� �Q����Z����$�*f���m���Y|�;����}���fn��7��)f����H,�mQ=}��qj��������Q��m\���ۍ��F�\ܱg��F��u?ɐ�icE�x��H4a�}�~��BA"q�wgK�-sܬ��2zz��iv�rrդJoo<�1m�l�U)E"J)���,�~n��q}Fv����@+�ݻ�� 3k�i���uȈ{o�߀�o�$�T�1550�+w2�X v{�D0�Quu:�����R~H�޷vI'\sT{��(dI���"&<f�*n6��5Dë��� $�{��� ��8���&��w������n��omݫ��(")J��5E6���5,H �/<��_{ѷ�ono�S^�����DA�ܛ�,* a�����L��>�oa�e��(���<m�b�f��=3uq/�в*u:��/k�
��\D��T�{zz�\�;Ѳƪ6& T�bbD�R�$����;if}���/ο71u6���8#n�l���ᶔ۷٥۬'nݺw+^5�.��c�eYk�:�G��;!�n���ا���{Inub^�:���\Z%␭zm�N1�֚-��]��5#�0pFp��6ܩ�Ұ
��y��>2m�<��[�j��۞۶i��zGiwbˈɕMv���t��m̒����<Y��[��5�6�ʇ�Z�{+���=��l��ֺ�ޱ�����J��(^��_��Ť������M�t��yt�TVw37�.�� ���?d'M;�&�6j	����K����qKdif(�re�;щ�A��VM���͸$������F7����ꚪ�E"&��ƃ�u��y�@����)����D��t8A�Ng�^�	�}� ���(&�K$>�˷��+|z�� <������9i�	"��n]��ɅE�'{�`��y\�PR��5_E6k7��I'���A�
�͈$ǯ:��6Z���� ��Jŋ�����2fB�S�'{r���,�ݳ��&��KpW��z{\^Ǭ���˵G��؊
ULLUM{�_VG���j� ��Hgg<�rnK3�M��I�[�v�82t�9h�5�=ETIA�Y����줒��<F��gP2��}|<�{};�о�ԛ���[v_e�e������9�s�曊��Ʊ�Ǚ�`�ޝ4A�g���@h���p��[�s
_�aS?���Ve����7�_� ����
+���郈�ۋa����a���-A��D �=�ԀU;�s��Χ~�Ј��9` ^�mڰ�}�*�%���C{��`�f^�F���$K�n�JI��<�I���q�!���3�D�X��	�wN�EMUS2�=��w`��7z�<�ɻ�<�<�����7,y{�Ր$H�|�>�e!C�1U��a����]=f����bX�Xe#;����[!��v���h��L�"L�����=�6�I�s� o{���_bhXU��N̗����3ov��.��U@MD�j���5�c�noU��~���.���h���wh���4�>A1V�"���F3۵�3~@�-�Xm�2}g�[���=��qzy���os`p�Qd>��.�i�C;�0{��=&}���Ć$!�n9�b�߮-cvVtk�U�kk2��u���Vp����ymW��| m�ݯ������g��dD�̙�fL)�6���_p)]�5�N��>��wd@۵�6�@^��=7хޓ�m�	��so:�LɁ0B��C>�楈"7�5F���|�%�S����H�ʉ�$��m��&�wX���rh�0�D�D̉"JF|>�zxѸ;pskAN13�퇞��%jz��������X�&����V�]݀Dv�s�  W��qa*5n&u�1Y[�,w�0{@$�n{��C�E����"$�6]+u�Q�91�D�+�݂�"�k�o� ���/�lz�t�b��}wۻ{�����5PT�H���ޞ�� g�j��;!o�*��sk�^�@oOq�!&�����?�d��S�m�2}��k�2Q���D(����<ږ|ޜ�- �E���r�`�^�̟fz2/b�s4�T���O�1�e�B�U���\��Gvw��UP����V���¼�E�[F�<�j�IW�,Z?{�{*ل�k��D��@i��l�ry[(���n�b�ݬ����:�Sϯ K�[È`+��r� ����[w�����}6�&�m"���L��u�#O)�f�a�5���ԨxzS�f>>~���Ӹj)p>���F�醀@[�ۻJGNTЀ�֥��s��D�kv�����K`�)���0������~zkr�>� ��9��e��VA�[� �.��r��Hv��2�L!D�e�x{�@|󵸈�*�_���Z�V��5���:7n	����w�ɭ�b��	��MQM���ytz��@ ���$w^�ݠݮ�TDC�.s��)���}�k)�q���'�ݖI�%��:(�e;��N�Ʒ/��7o��� @|n�p�L�^�]��yQ'�al�p1��Y2eP�u	\g�)5q���N*ΐȆ�t�y�N��$onnй�~��/e`���9��|����>k�_�8��gl�v�w�v�^���\�Xn�o8�ѹ��/�=u!c`�.yv�9�͌;�q��:��=�K<s���K�g��wg�·+���ݤw�B^m���e�=����ڛ�v�κc�:�1:ۖ6B�a��셞���s��À�Նd7=�^]nû>�@��S�W���m8�h׶�'%*�^�s\ݞ�Yw!>������O;k�h���	�	/K��G�]�$⡵��g�؝���-������M���bV��K]�~�I8����I��W~	E3���wW34#b���% �gz�O�_�Zm��)��L�_�(�D�w��l��( r�n�,���=~'��l�7�w���Lk��6
@��.ey�Wn]�V��԰�9;o�EzO'[yu�h"#2�]� ��?Z]�@�L%IP$���v���D�9� +��ݑuw��^�����9�����S@"�w�iX]s�����l�0�����@��B��|��$��n��ͮ�A�������P�=�ǳ'�r��DT���3�P4�ֽ�˙��a��b�I�O8� <�e6�����ٞ���iQ"�����~�� �3���0"���ŀ�Wi���v���m�;�x$�;��0Q�q%QPR��48h�7�(�� P6���55F��ۋ�z�(���2Q']b���Y����w�y�����wz���6�&,�Ǹ� ���kfO���=��o�I$^}\n���`$>��;��b����y�險��DME!�]s��fy� 0��W�����o7��3��� >���/�Ϋc
*f*&���v����V*)�V�'B]�.��$�\�v��H���<{����b�e,r��N��2�v�Sd�� �`9�c�6@$�9�S�h�p����^�d7�y9�X "��n��V��I���Q�<"	B�e@RH�oX��lV��-��m���ʱ�Ńd�-�J۾�?�S�X�U)��1�c�q f��t"���f�=ɣ/��KՙPK�x""�!�q���>����I`�A�>W>&�����r� "�v���I��\<Ӣ�S�y�Y��QT�eL�8h�7�� �u�����+җ�m������2nJ���m	��4F�v�Տ��؞V��
��|�j��ão!�����E
�v�j*'k-���~�/��_O��~]�C�Y���﯋m��8S�}W�n��n�2�"�]��	oy���	�Yp�����5�QD�[��6c)BQ�2baL@�חvI �8t���c��{g�0��wv��:	�r� bk?������iLn^n
�[ƣO�!�	�s�ݛ��V��ۤ�nL�9|v�S�~}�����3����ٻu�����vA$��吶'�skau:�@#�[�Y�*	*JS"��5�q��0{BwU8���	� ���ݒw�k݃6��LfE�ڮ��_V�ɉ���D�"�Y�b�'Z�B�uT	�����@$Aw�ׯ�zU�H0%�Kga�c7��M�&P3rIȚF	>1Wb�'����Ƞm��A��#��+:�ߐgy���G|���ɍ��E��SJ�VY"���:g.l4����s;���;�1��l`��gI���ދ���O�/��|�����}��|MUD�&��b���$��B��揲��=���b�m�5��ܱ�;��I�v�#�'B�e��9^�<���=��Z����cQԌF�l�/��_�8�H0�-,�.��  �׉�>�ۗg)��{y�,���I�,�}��L�JP$��y������uIݨ�Y{�X	'y�4	$[�˰D��Gێ}/��[,�w,2��2f�}q�$��ʿ$�@�Ŝ�ݽd���K"��r���0�&&R�T�U����Ú��T>5�H�����~>��a��f���#|Hȹ�����BT�B"$���d�2����핦
�Vdq�	{۶,�r�����&���<��r%��uGQd���P��n�(1B��mdX'4�8��U�.&&��4mjzw��Ex�ӯwWg`��ӛ�Q��4i_��ܲ��f�UZ&��$�X[��E��&�%(&K5Oxd�\�I��<m��>���~��8�v��c�ؤO;"��&�9�6Iq�)�²�XR۹�Ahۡ�nv\~m�����}��Vg��0|-�w��C۽���#=��MR�����6�:&��wZ��5��Gn�hm����H��⫻��tk4�5�����]i�Sr�]ŝ�#T�&�DT"ۭ�${Z�C�D�ݨ��J���\f6�ڂ��j��Nva��r�է�Spgy����z����8nD�Y����R]�m���/�i�x�����'�M�.��k<���IQ5�:?p*�/{٢BLIۅSwޞ	f�D��='�
N^坞0�'j�t^=�|�BKk1k�6l6Q����W���B�����a9�-ˡh{K[�����Ϗx��;�v��&E�3_zv�{dŚ<����,�gYu�x����x7�o�1P�E�����NP�*E;�q�(W�Z�yw�b��b>|/�sb�8���s��4�ٸ˸w3
Z6�1�v"p�hL���jf2�ps
=�X���-�Gbp���T�Û��F�݊�SX50/([���^�DHm����i�|\S^�B�;���zf�Й5��d��#�0[��|��wB���܀>N�?m��,ܦ&ŀ&��R?7����=����n�_<���x�Ȓ<&^|:�mt�ԢV�U�Z�ij�km�mQ�mB����h���,ET��m��UEJ�Z(�E,b*�+Dj�F�ƕ
��J[ZP�1akB���D�A|_ �� $ �[Z��Q�֍��D��m�
%�U*ҥkimJ%��ke��J���TJ�Z�Ѵ���ʨ�2�Dڕ�b�XQ�U-��K+X-keh�ؕ���,�e�km��Q�k-�Z��c+cem�,�V�����*6�(�խ�
"�Ud��єKim������T��҉+[K+YF�mm��[Q�����)mXѤ[m��*���Dm�RѡaR*�J�b
�ȱ���"VڍV[V-��"�D��T�iV%J"�kF((�ZT�"��6�"��H�R�E-�j,��#%T�b��-J��hՠ�iJ�Y*��eZ���%b���[YUe��Z�h�eZ[*"[e�-Z���$QAQQkR#*KV�kJ�AUEU����j�,�*��j
6�c�U���&����nAηF��4�n���Ln����%q��;Zz��)m�܁㮱�&ݧv�ċ�Ńm�<�^DFk�V1jǧN���In:�pn�/=qGVx��ˣc��2��k�Q�x�-�P1F� �;m�3n����c���r)�v��M#�pq�VQ�Z�0p���C���c&�x:�Glrݝ����6����݅u�v������u�X�i�]��k]޸�P�ɗW=bGmՎg����fOC�c�km�=n�[��i���ܾݫ)�5m՝G%a�nm���1�d��<�Bkom:��NW�TT�n��e#�q؝�絕l	���A��aq���v������<�v6ܓD��6ݵ��]��g��ʆ;^ ]l�8[�o[�CB�C'<㎖t;<c&P;qӓ����Α���R�������x.[z����M�&�[�.1<zÇsd���fw$�i��ۗUa)���y�l�a�����v�ƻCHc>܄9p����6<Y����v����s�h�WcsvM�[hQp�v��\�ڬkny���8����宮-��T�����8��^��n�8���6�f8Z���=F@�V.R1U��6{q��v�Ʋ�-�Q��v�b7,O3�ƌ�]l�>j® ���0�v�E����N��m�u�J�9��.l�g�;yw+�װ�S�=���v�Nҝ�ƥ�cF{o<Dn��n�z�q��j6���e���f���֞9+�,�E�h��m�Aq�ۧ9��ynv��6��m⎡��Ml`���4��rn�;U.+���g[En�vS��{b�zN�R�{g�9��Дm�Y8���s�F�Pi���Ź��=����<�����Z�מ�����J.�#���y�ܣ��Ywl=v�`w���c�.w]�8h�=n̻�.��@t��܍����=��q�y�ĉq۱�r��[F{�r`�A)����������G'7Cw>��a����{����_�vC�Od�wh�[�{l�A�
��=s��(m�C��n��U����\gw�7������9Q���x�$md�1ɗeV�=u��N䭹��Nx�4S��8K�r)n x��^|���N��*Ƙ�z���z�v���:���3��x���6�]���F-5���s��t�����v��w[�����f�(�I�����Ba���[�@��iN�K�����3��K�niG�=�������{q{K��^D.�����5/d'�܇^D�^n�X$�2�;d��i�6�	["kzYH�{�~$Z����B��h���Y2f�2�_�����$��n�#-�X �OjD�,L�5��D�Q0d�I�w���$�{���5x�vz0� ��nݒO�_s�����a��,m����UF�>WޤgM��$��;���gokm\Z�7ѕ�;U�W�GM�10T"�H"���wX�	{�����lL�ؑs�(���$]�;�A#w�����q�g!LI�r��W1�v�wJ.۔$�=����ţt���g]`3C�T��ϒS(J�(DD�����$��݁d	�,�7��`˳��tZ{W9L�O�_7b�S�Q3*eDd+�}���1]�N��&X����"�T���f����쟷}W�����z,rr��&jr�]���$���!�S�y&ü����ܫ�L�GR��xx	��t>$���w`�w~�hRٮyÉ3�L~F��Ƃ��h4�B�٘ ��xP$L�HW7zI o���wzY�������`�*�v��o�:q��`&cX��I�,׉6�v���Q���T�`w�3 Ȯ���a��,m��:�e"H�n՚rVX�-&	��$�=r�x��j��� ���F*�'9��v�YxdMƶ�3��ïj��C��+���T�|��阘(�R$C*���O��C4	$<�۰h*U�pFb��w�B��Yd^RJe	R���s��I��eos�����eFk� ������˿}��Z���Ξ��~)�[-aL�Uf�#�owhY%�
�\��jc"��QӳI��v������嗖ɮm@��=�����k���p��z��o]8�C��X��"��6r�=�.}3�\�4ះ�=�����w��h3���O� �}̜h,L��K7�C�`�[�t�%����wv������+&�nHzx��.P��Q�{v �ǴF�a�H���[�۲I���ts+D۾�ւ*�NRILn�+m�}�6��bo�2���m�Ӗ�]�>~�O�J�J$2g��FP@���ՂH9���pLHm��"��M I;ۻvOe![M�H=/�H0;����@mmX���4� $s{�`@9���������]�(y�I-�e�q$�o��.�$fswdq7&:D*f�>&�n����bϺ�r��Ra2d+��u��E������ ��_}� zY��u9,Ҁ�cRbfN��0�g-v�[�h���_"���Z<���otȿ�U��M����b�U�x��$g`��o�z&��;S�p�/�g� Q����A{�:Yе�V�3��T���2��'���|��z4��'�xS�?�����v�[sr��Yf��y��Cb#�!��9�lY
Ah�k������;�8n.���ާon�$��w��oC4l�/*���d�?�u� ̋ڎ��S��&����@ת���&VI�}�4H��w`�H�Y�|G���+�u۞$8�����*R$c����H;�� ���}p4��������b�����$<�Ikd<a$�o���卛�t�+0�w.'�6��_����^��<��k���Ng��1�o�ٗ~�(�laL<2����D��ݫ6tmvℳ �uuY'5�>y]���"�=�U���r�qY�R|�Ua��ج�g=
J�y�LĤM��Yyz.�ME�����ِ�g7����� ��G2#�(K���oI�lmv�:��c4�-�wX�pE��j��^�.������]ّ�9��pQ�WY�;�J	�;8,��I���kg����[�)F�������]A
�v=�5k����WO\z1�v�����W�z���n{nݽu;m�����6u���^{{^�x�gp$v�[&��ݷ<[7A��etf|��"����4sz6����$�ǃսZ�
m��=�<α�>�<�c�����"`��S3* |g�]�$��äA>�����Z��,�ջ@���O��f��2&
�
D(RMKy���'���3ю�<��},� 痝v	�\G��z��Z�2�-�������H/o:�Ă;k��z��i���$s\�D�痝w�}Ӂ1s10`�2$a��![ot�YQ� �}�y�d�s;��r�_H�Z3H�1p��"�R�$ʔd�L��kz�s9��@�uWg�% �����&�d'���s��g����]�5��F�ڃ�Spq�^�K�����m����Ju���~~��5�e����7��&��ՂI�'1��vl嚹7����|�~����~l���i�m��p1��v0�u{:�@�:�1�c�����A칢uB�4w��aީ����\��{;.M^�չd=�s{�]���-7�v]���0�3�{�xx�����v	$�}��^v���N���'7���"B�*"I��v�����z�t�6X�6�j�� ��۲I9������Xe��=>W>;�k��0�GMnՂI��ՀAo���x�����u���E�Ĉ�L�E�7���C�(���}j�8��}b� �>t,����#gp�rB Ȕe%2�Ȝ�n�9���srLqgJ�f7Q�.���9���Ko����JeJ2b&}�=}b��9�����У9
N�۶:�P��Tӻ���|���ꉙPdIQ&B�]}:H2���s[O2��_S�� �	y�ݒ	�t(Vի��A<����`�R�j"b�S2f Q�yu`���P�������<�۹��]�&@�]Ż{�z�k��k����ӎ������΋��t�Fn�'NH~{�l�c���Ǔ��n,�æ��1|��Ϟp�A�;�v	!���3��v�I�h$��=u���-J�<	 �����I#y�
$���g`A��<~���9&A��j�1�Oa����E�3�gB�r�dfF�4��ɜڲ;[�@�C�λ=����V�����8��4�ʯ���#={+�b\�b�z#Yޖ;E���Q4W�z�R�U���E)�QU��ł�l� ��Ρ��S�\�FWA�5�1;�b�Gwm
�����*Pa&�yv�� \RH�f��M� ׾��^fu��i\�1��o���;�DL�2$��!X���� �y�V	� ޳F��ة��I#��
$���v	�:p�L�������?D/�B���/�~�<��q'A
�c+����ѕ����^���ڐR����4�������ӻ~�8���9oO_-�YwEڕ=���+���2�0{|Gj>�F���z�G�պ�\})>��k��n_�HBG�␬?���֠����?�1��c���m6�]���m6 VVJ�2T�?����}���V��� ��
��}�ﻣl�ed�*AO��y�lM�:��,sR�l�	Q��	L���/agGf㋭@�ɸ�;f�v3H!�m�"�t������������������a�����HXZB���}��+Fh��O��y�M�T|�yg��`,�L�}�PR
ĕ���=a��ag=������p�x��6�q�N{���l�J@G�K�^O�o���Y��7*����H�S�}�}6���jB��}��@��Hx"kz�k�2�_S��'A��BwI��%TL� ,�o>�i�����2T���捉6�R�5��ϯ:�|���
��*�}�tzɶVKVJʟ}��D�&��W��D�1"LD�
���~�c��_M��1�;#���6�n���`V�
��|�=i�@�D
�'9�{�,�ݼi�<�~�B��X������Z��!���B�SU5U2�Kc
�~�7��IP��?w���2�j��g{�{��%@��߻��q�
5!m>�{���
Aa�w�^�>���b��6�/�Ym"����}���_N�Æ���]q%[�+�\�������JO-^�:�2��NȺ����<<=�{�d	��`�R7[�Ɠs�C�70a�&�r�ss�=\�9�g�{��G[&�tn����򛩹���.�9���̡����p��3ɷM�<�K��I��8�����r3��Zx�a�'���9�k�i)4nݹ��k�wg��[4��k��ݺv�m�y��rwg���[�݂;/����c��=X��i9�{},�E��B���y6L��"���ݳ[�P��S���&���"�=[��������t�
�~~���c��o�fx?�~O�'=���m6�R,d����Ѵ�B�+
0�?s�֠H�${e�|��|N/���I{��{VJ��FT���h�M�Xo�g�<��g�\��}4���=�~փ�jB���l/��dؒ� }/����<@ ���y������@�beO��=�z2T*J�w.�s���}�nf����<��|0|�^|&T��D�E���*w����&Ь�Xw��d��Ĩ}�ƽ���w����jB��7���7H4�+D?s����	X�d�I��*&E�	 O?{����W\y������+(�S]����M��Ý��+c
��R<�����zn]���������I�>�ȏ�����@i�ҙ2T�1d+H,;���B���@�����vR���vN��߱}�>�u^��@ ��;�sP��2T��C|��Ѷ�+_p��ޝ�˗���<�c��yȩkt��2�t<�<��7
ۇ��y�P�\�u��?��[J&bfL�w�>�����6��R�w�h�3
J�f����><Q�����A��5�H����t� �����5
���~�~[���x[ᙞ�m6�����6�@��%|��ϗZG#�Q{�BB���W�Nk����q��[B~�<>��=h!�n9k@�dli��d�!;���[��}���tt3-�Tś�=�<=�ނ;��ހ�� �����=�a�
��*K|���6ɸ��c+'�����������$O��YMPF����1Ѧ�a�sϵ
����>���h_"�"�"Ϟ��^?;¤Q=Y�y�����Q9�뚅g��P�J�C|��Ѵ��g=����\1��/�������@K����k`=d
�YXy���Y=eH(�7�}6��E��Cs�� }�4埾ʖ<�
�^��H)�_O;��<|m��燠)�$�?o�6�*Aed���w�7m9���;���l(0�;�|�X{T�B��}���d�+%ed�>Dn}�P�0�&���WT���-�����~b�N��=:��q�����rp�pk�C����<�xr!w����Θ�������tk�}�4�$�-�o��=ܤ+X�
�o���6 T����x���pO|޽�+=*IP������R�ʘ�&"fL�_�>|����}�U�լ���ߞ��f2VT
%@�����ư(ԅ->�{���)
���Ns}�/�ї�_^W�? �Cw���"#�3<@�n$�s���m����9���%aF��۝x��vj��ݞ˷q�i�?Y*m�`�#���m����n}*�`Uf:X܈�^N��\C�Of�<�4g�KzvG�۱_n�����z������0�'��~@T�vxN[7��r�:���s/�B�VݡX�j��[��C�vj�h�NK��A�9]�a ���)���]tw��>��
VK$�g��H�m��r��y���7�|4�&J��xD�C�y�<޾5w{s^ym��^$��3E���ř��)�17���� :9ڽ�xt��Ît�g�v�5���FUU^�HUf㚉���y����OO�w�ˬsV�v~w�`,��`�ܜ[��2�s630E旾�UJV��a�G)C�^��f�IÜ"�C�C�/<�7�/t�{<uN��B���ryzvF�UJD���B��҆K���4䂙ٺ�e��2�� 7J�b�8��3<�Rp(l�6<��n�<��Y2&;�j���Ꙫ�גw��T��6��r��Jf��ˆ�f�1{8�/k2�Y�e|�c���ap�������t����n��;ޅ�^�]�3��p����m�Q����y���w�W]al��3�� ��v�`��_���⥱�8-ɩQ`��\�V�0ڈ'ەv����V(w�M�M�Ws�0c�{��(��my{,�L�鷸\�/?�AA���x���~֑���vY�}Z�߽�|�K��V�$�:痎����ށL�'ؒm�H*�ǲ�˸�K2t]�la��:��Np�_2�jZc�R�ֶ�[j�T���VQ�Vص��
m���(�[[kD�T��������KT��i*X��QTb��[V�(�J�����j-E-�km�+*��`ŉ��J1m����QU#-Z�X�����6�V�V�Y-�*��4FX���VҶڅ��[E(-�DAX��KPkkV�U��(��J��+j�Z؊V�ֱZ��!Z�6UVұ[J��R�Yb5U��*�Ej"-Z؊�m*XЭe�m���ڶ*�)mk�[U(ƴb�+iTc[e�*2��j�R�Y�b(,ĕ-�(1�TQ�
+�̪�R�m�(�5��"��[ZX�eī[j�EkJ��R����*� ��mh�D�J�Qb �f80c"*�l�\V`��`�9�m��˙Z�DZ�cl-���bV�Dd�mm��bZ�L�&#*T���
%J�"��� cD*bTU-(��%kE�W,DTTWʊ��

��iJ"0kY��1b�Fڌ��FՌ�UZ\�2�3���H���{��?�T�B��?wsF�6��c+%S��~��6�@����%�Ď�-��|Q�w��5�~��~�{�RZw�����!Z��;���� ��eO�V}�p��o廊~IP�y�^�F�laXS��ft�.L�-��6�S��h8m �VV�|�Fc'�|���}����1�T
���M�6Ԃ�S���t�t�j��sP������|�j���~��_��t�z���Ԇ��㞄c[��L��۳����"߿{�Ͻ���5���]��h�l@���YY*}�߹�q&Щ+
0�)?s�簬=T���>���{��@�5��=d�2�VT��o���lM�S�w�x��p�����M�7ÿ}�t������y����{���}������;�s���؁R�e����5
�A��D���%a6ӣxʟ�3�>�%���W̸g��xe��,=�*y�|ހ� �lea�;�4z3
A@���~5���s���m �8Ԃ��{���
AP w}]^�>��̕�""DDH6 � ���G٫��kPz�����2T����@z��J�XY�9�{
�=`��;w�}��{�}[#0����EڍC=~�6�3KS�ߏ՟�C�������{ݪ��9�e�j�y��5���P���7�K���&OBe��  O��'�eH)����i���_Îa��<sM0=�a��ϴ��Q�� on��x�G� n��Z~�S����� T�a���g�%Bĕ
!�}�tm��V�����y������;�~�������Y�	�1��u�:ϦFx�ݝ8h����lb��������\'a���k���u��
�X~�|�Fc%e@�P.�����A`~�;��q��[�>x�S��������j}]^���B^�1&JR$�� $ZMs���i�����}���}�{"������J+>�u�aR
OD*J���wF�6��FVO��������a�������@W��DĕLDym��q�7߼��
B�>����x"���D�5��
ɉq��| d� T���;�5
�c%B��X@�����O�,��"LDȅ7�O������e]��H҈]��0,�|<@L���o�}�ј�A��@�������q�
�o���������O��+A߾��
���g9��~�33��\�}h����S�@�����Dv}�P�G�����5z��'��0��Zﰬ=aRPB�w�}��L����ȍ���{� ˊs�*T_m�:�/�n3Jc0��x	���p�CT��.��5�`���"6����e ��s�����w���ݺ~ W��>��{������u�ٿ!|G3<���-���S��;�P��.^�nJ�Uی67R�>�649�1��>��n���]�Sm�y88������m�I[�����:��˶[���n{u���.���H�E���k�����j��p�	x���l=��y�npT\1�ڻ���-K��{`sq�9�c�#L�Su����6F歮�����kq��.���9͂��!��7m��n9�(կc��d�u���y���	�����g��3��<�����k{�>�{H)-�}�4{�B�`V�K���z �0#~���s��Y�>�β�=d�T�
!�>�����
þ{vp�rfao����9����Nww8�SQ��q�uӔ7��}�|�߾��=`m�
ԅ��|�4��
<	�*��ck@�;��GA��P����|������&��}Ѵ�e*AO���ѱ&б%aXVk���|��}��]e�&~�G�A�DyI��}�F�&�Y,eO���D؛@��w��g���3<��m���7߼�s�������v�ĆZA@��o��vR �`T���hSh ��;�5
�ۿw���~Cq%B�~�ﻣi�r��D���
k��|��0��)��ea���d�ǻ����\���q�P.��s�lư(ԅ->�;��� �B�s��_A�S���������[&�`�2�$�t�tv���E���b۴�FTf֞tE>���}��+Xnnx=iؓ���4m �c%ed�������%aF�9��簬=aRL�z[a�`q��>��{����2Xʟ���@z��[�ޮ9��y��S=4�Xs]�z�H|ZA	����<�ǧ�h?ֻ�_�r�h�%@���E�A�&w�����^?�^�-���r�ӹ��\}�8����'�=�j~:n�'.{��HBg�޽��k�`T�>����M�
�Xs��<���2T��o[�{��}�y�����y�a�°����2ܙ�[�g�����{�h6!���FV��xz3�KP(� g�g���߾���>�#����o?�����a�w�CI=�����>�RTL�  �w� ��;��J�;֧!`_�{�D�2w���4�S���5˯�����<�+'VJʧ�����W	!/��hUPJ�&h�>����|_R
B���ߴ{�B���<���
}}/�o��i�@��s�CID�
�?}�tm���G�k���/��)}2$LI&b$J�W^�ݫ���n}��nէr�m�7o*=1��q�^n>�~�:+�g��xe�XtaS�o�h6!��
�FV��y2zʐP)��}�M�����g�� ���h�H4�+Po}��dx,v�ɍ�����A��&��?h�n VVJǺ�z���M�RV0�(s�y�z�хIb%�s��wF�
Ad�o�߼�\я�5�/���
z��@
�v(�32��4�M0=�������B��}�����
сZ�����'㿳/5��#����Cs{B��Ń��@ݼfAz���F˱��y�� �o7E�ۇ.�v�G�Vtݹ�駳|��k���$�}����?���{�5
�P�*C����F�f��cr�f�f���*s���=N��?y��H)�5�>ѶbA@�P)����M�6��HYi�����f�闚�A�HV�k���B��*R��32faDI��6 $Yv�ha/2VQ���~���i|�G?�OyV�w\���
�P7ϻ�G��H�$x7~P��W:�e+�
�ƿ��s�7\�&�څ��v7N�u�ͳ��#g�}:ݩ���|��WXX�~�w��7߼�R�HP���ߴz�]�l`T�������M�<淭s���m���u�څg��T����=H�\��ʕ"b&A��|/��/� Y����z[��?A��]x#�ѕ�T����z�XjB��o�� f!�PC���q;¹��+ﾯp�B�o2cf"&eD�(�l�`k�}�H)�*s���%aF�y����5���{�T���%O�}����n2�VVJʟ}��D؛@�p-6$���A��;������-���=Y�VdB��	K����_ �0*YϹ�z�q�@�8���|�ڿ����[]�)�*�ؚ���.�y�%z���Vh l�F������ީ훾�pS圁��çz�cڏ7�|s���O� ?��$�T5�~��l6°������r�f�3�m��T����t�m%B�Q�����h�3�?p�k�Y�@�"<	 Ge�>A�
ԅ-9�{��t�JB�C��]^�>�6#��k�2/��"L�8
�6y�gk7@�9��v���i�Ӗ�c��<��E$����bD�(�11'�#�<�ﶆ�
��YY*}�9��6�V|����x"<	ۄn�6��d�`ZLOk�ѶM��Q��������&�|/�j"eD)* �60��G�>�����B�C��۫�����~����
сR�}����؁YS���j��J��J���ޗ�f��>{߾�Ԃ��_|�����y��y��������J!Y++~���1���*��|w����{����Z������� C���j�`w|�٘Q3*&!D�`#���F�m��i`
>�}�G�"+~��hQ%aXV���°�aR
<���ި3[�#*���y�#� ʞo�6�g��}���y��x��M$���|8���)h������B�|��_a�����0*Y�u�z�
l@��s��5
�Y*%B���x��Y�����]tfS)N�9�������ދ7_{ƗC`������
n�}�@݄˷��!_k"i�;�.jy�g$uˌ��
ڟ� x��{�vF^�1�;�En����u՟BI��"�v㶶_dfݶ�-�{a�'x0�>Ҭ��\��Í�g�����9��%��h�l�h������g���֮f�s���\u�ˮ��<��U�T����;m�9���d�β�B;��B��f�
�"��0�=��۶;j���u㰽��7=7nºl�Ɔ����ˮ5tJ�1��-WIж�Y�/�WsM�t�kxs'3��cuA0D��n���DD	P�xY���#����&Ь�2�����B�D�o�w�����wOL��HnZ~�������s��5
���K�6|y��73���
����� �s�^�>ߚw&����4tI�*J+��\���
��T�|���m�c+%ed����713;��O��@��w�ٙ�3�.b�zm���7߼���AHYh��ߴz�]�
�G�󿹩�-�Դ� 2<	"uux"<(z��P�>��a���������&"&��|,�"!��@d��7�d�H)�y�9���d�� �}�߿h��0�<	�����T��Zg�0_x#�[��x#~>�m��0�fTy��y_@�m'=��h�m������7��@z����w�&�0�V��u�aXz0�%���F�7Y(�yx���u`#�u��m��Nw6�<�N�y;7V�̅�������u����Fۣk��m߿��xE��c��~oq�ko�}��ą- �o�?~��Av0+FO���@z��>�k�Ϸ��j���?0�w�u
�Y*%B�}����l6°���g�fe�\|�Y�6�l*s߻��IA
�����x~מU�����|�ĸ�4���|��ݒ��Qn*��z����*p�,�6M�cDc���������
be�˄V�r�i2���y���<=�x}�>����}(ʐP/;�߽6��k� ����P1��F^�:>$)�������(����"DB32��"�#���m �m����9�=H,6°����L��Zld�������D��߿h�Ad�+%eO���D�m����D���F �,�(�_�?P��Y�����!|� _!K���'b�D
сS�~�4��@�beO߾��|��Ͼ��ոg���G� P N���l60�-�����|�˙�y������@z��+%ea��|�Y/M|}|�Mn|�P6y��ޛH,�!B����4�t�JB�߻�j �~�����1��߈%1���L�H$�H2�MF�1���ka�v�i݄�ӨAO�����hf����:	5���M�T��S�w�Ѵ�H,,aX_߻�{
��¤��9�i�\�s���=��V�a��|��$v��P�0�+v�D(�33D�B�����ϧh0G��C��^�X�
����g�9�~�R�k����y�M�(�YS��뚅g�%B�y>��D�������2��C��x�#���g�32�.yn5Xm�N����lCi*��������
�~�� �b>(G]Oބ�;6^N@�p��BS�Q��eN]M����W���ͨ�v��)�ʝIh�Wkh�%�v�m����%��[�Ԫ�������O���
5 �~�y�6n�iHV�~������P�Ę�!B32��"��gݴ0�+b1��	�} ����T�{��m&ТJ
��s�V��*%�w��d��u�w}�����2z��FT��@�9�o���������w~wA�Ă������^<u0�߬M���t�B'������
�@�?w�sP����A%B�s��F�laX{��\�����������bܻ9�n�9�t������rnF�:3�I.wF�a^���u��?>�?q=<睂ã
�����M����?~��*A@�%@������q��EF�����#�����u 3�+�x(%����G����aQD��55SJ,�`#�۽C�'����8����f���~��$�%aXV���=�a�
��T�9����i�q���5URk�>?E��$(y� � �]�p`�|���s��=4�X~��oA�i(������_"�"�"�!3w�~�|��5�߀�~*X�Xs�<�Y��P�*��w����
Ú���s-�DJ���q��B��y,��~?p�����Ğ�VJ2���=f2VT����~���ư+R������.�zܘN�����{>�e��Q�}��}��q���@!uH��7$���np38���U\�������FC��̿g5�����	_�JB��~�z�G�"�E��"D�dL�F��#���؁R
AO����6�h~�s��5����Aa�}�_��a�¤}���=d���YY+*}���&�h�ÿ�������˿@���N��ޝv�ڎ8�m�������3ݸo�&\]��߻��$Y2��ӌ�����c�ih��~���B��Z
���������=/�i��9��{���Y���D���C�'�<�v>FB��&��XT����Ci*����y߿:����|��ј�FT��w�������HR��������/s�+�$��x�#����,����7��Ĝ�﹣i�
��R
s}�4lI��°�=Λ�˯�u����R
O�T�>���ѶM�VKR
}�w� � �۹��RE�@�S�Q�~���@nh(��9VI�HVe�<*Ak����4���R(��u��G�u=�+�ٚ�._�d#Ȁ�@���i����y�s-�_.V��l60��{���m �VV��9�јɿ�h��oq@�*�w���l�`PjB�N������a�w�j���G�R�}����	4"�"c���WZs:�����%�(�)�ɗ���?w�}�g��z�r���}x����5s<A�g�u�3��G��:�X��$�#�^p�Vx�xz۳�d�:��U��՜�{LG93�ü��9<)�gy��q�z�0A:��[�=Lɰ;�i�&UdA��M�q�l7�\i7c�����,�q�23�3�{^�b�����A����C�����(c;[K�T�<}/��	�^�J>1��5������GvA�����Y�\�^�����p7�wf����ꩽ�X��&m�`� {�Zƀwu��yqɽ����u_z�ۈM�,D~�����U�ǫX6���w��"K��C����R�h�}��I)�tH3R��{8-=�M�UL����"�e��W��'0���`̈˪�E{�_kZ�O�D�{^�ce���!��\�s5S���2�쳚	����ܷ3�9��w��p�upн:�݆�`�B�oo�o��ݞ�dѸ7^�*�:Q$�4w(l��WP����e���8�]
�&��ֵ��]�[31I���V!�(��/l�����H�kjt�C�����0�mvP8��8W���w�N�N$�c; �}��nzE�r���#]."�����c��^��ZU�mŗ	7<n�s����ZU� �3l�=�|����K��W������������)zs5n�c�{<�����T��P����u���tf����
{F�ٞ�1��W��F��t� +��ª��̥��)eD�X��kAb�)��3A�R�X*+R�#r��(aib�
6��HƵ���QX��FҊe�嬨Q���QQb"��E���m�De�F����b5�V[TjX��W*��ܸ������Q˙*��J��-��ֲ��*�h���P�Z�R,U��4jU�����J�h��W@Q��X%Jɖ�TDX�`���!�-����1���Tq�*��"�J�b*(�bU,ƪ&P�j�QT̸ŶV�ł2���-DUD�!Z
媕*a�����Pab���c��*�����`�`�ōh��-[`T+LT�m1��9j*J���V5+\�兊Lq1Q"�LL���EḅIXbc�&9�T��(�������q�X�(�ַc�elX�G-*�T�#����D���0�JȪ��(�[R��Z��Ę�Drږ9j�R��ܘ*��`����f*QD\�X�PS2��h�TC.&���|�����[��z�5����d;q�g�@��?�?��ǍJ<�;�mr���;�5�X��;<��8��{f|ll��5Rz�3ra�n��(\����zlu��v�h���.�;m��͌bz�9�ֻk,�t�ee��ۘ�۵%��x�rF�q@���'�^��F�v�m\��D%�{z�7��պ��vn�.�[��5u�[��%�-�;6��l�6��((s�v9ι��'$vz����,�6���qݶ�^w9�%�2S"+�u��wI��5Rn7j&,\:2p���U3�͹��bn;Z���%J�y9�g�Pk��b6��W���u���Np�/���~Bpe]�]��=�.����{�d�oLT�[�l��v�)i"�la������{f���Uc(�퍖�b��cCq�Cq�[���56:��]����]�޸c÷���t%@U�%zK�BW��6�Y�s�~~��9yҠ�6��T�1crnK��۵n%ű�@.B�ڇ\a��x�;%\�켹�:��Xnt�n�${;l�\;Y,v�ۮ5���Av���=�H[r.[�@���Y�<^��k���.:S��/b�kZ]�vq���vJ�[����]Zcm���ֽ�>y�nm\k���#�<k��眏e�m�p��7Dv��9��4c�n7��;��gs\��^yh��ݎ�3�[1��Mݚ�����*��e猯l�	�t=s��.��/]r��{�j�^u��m�R�l����k�n�-�6wAU��7I�>��e6BWA;V��vݶmqj�����ٷ![�-�sxnݮ��v������p�x����ӺzC��s����4X�b�����ls���x9�kO[�:1����su�ŭ�
~.�?��Z�P��q�Ը���3l-�.wn<��[]N��܉�����)���Ϫ6Ug$��b��]��x�Ęw��\�`�a�k��������e�0g�!�ʆ��皸&�M��&���7B���W�;�k�:�<�%��={�>����������Z���;��:�|F����ً��F{d7-q�lͭ����^��g��<ܷ;�ϱNl8��rr�!	ƻ[	b"\V瞍�\3p�{OOi�Vw'k����q+����(Ok�ld��Y��'��h�ӽ��j����]��^8�=�[��jD:��n���k��c	/�N���۶H�v��v�ڼ�`�lLƺ螣i��+Un�k���^�	+�=�S���j�!-��Ɂ�;'#1�C�[������-lk�� ������4m6�Yc%H)��s�6�hX$�(°�9�s�V��;�(}�N�|vƉ0��#��%��P�<,�����?~����l:~������0�@2,a�Q�~�,�	!�u��{�" m�:�C���^>K�~�=i��@�9���B��J�IP�>�W�;��y�ގ��0��pѐ����*b�	����e���T�ß��4z�JʁD�eby%�fH�߸|||>���� �+P��뚅}!y��j�*&&"bb$E�0�#�|�#���L�� ��>�>^>�">{� ���(0�?w�sP�=aRT*E�1��C�*m��5Ⱦ7޳�a�>�>DWםC��0���ՈQ
dē2$E�0=����څH{i-�o���r�#5�ߢO�sc7�2<	�; aSh�߻�5
�A��RT(��?y\|�Gȏ�}>y&׸��1~8UDԪ�bM�Y���a�δۀ��:\��Z�<�`T���F`�"$ʄP������t��q�����j��ʁR�{���>
>��'~��6bw��������@ot�i
�?w��R	Cz"d�dL�F�����#+(�Y�v}^^ޜ�}�2�������H8������m�Y��E��\oa+B3��4-^��ރ�e�fza3�Aؤ육�W����P��xx}�a���?�mV�a����j ����￿h�&�VKY8y��vf�ͤD���@�u��!LB��@2,a�k{���{H)|���=�R�
�L�z>�_�w����H)���?w\�*AC�%B�?}�ߴm���#�_.��сF"nH}�'���!��(��g>�.Y#�dz����|;�}�ј�FT
�����zm �
#��������s��c�<!���[^���i�*&&"bTH�i�I�7�4m6 VPd�9���{�G�q�אԱ�>|��zn�X{T�B������F�62�Q���"7��P��S2�ډ��k��~��ݝ�C�<���p=ۇk76�l�L%[m��WY�&D������ədH���(����څH)|��h���+X $-����x�E�X2'����Y*AB�}����6�l+
s��}_�������������tCi,��üQOc��L݀�$�ovł|s��݂qڙ��F%�3z�>�8JR0?DL����H���ŀI��wdF@a3�Օ�D�쁑k)X��')����w9,�餠7�l���86��Q�-]Z'o��p��
d�4t�^��ϳMa��<<op��gm'�/�ps�"&!D�b�L�du���j�+"�/j�$��:�H%�K"�\��[�M�˷���ͻ�����0%DL�S�+o��~{���'eqᗘsƛn���^o;�KޖDg�?��8����%ÏL�	H,�8�7�3=��u+M/l��Uk��qt�[��~�I�L�"��c��$<���z4��n�T����Y� ����v�x��"fA�"h}^D�'l�Q3*�2��|O�;������̸숄�lZ�`�Z��DDH3��������>$��Ǧ�9�q��t���п��
�>JE��DH(ș���{�s=%�.,�[���I#w�A�}��Y�j�V`�����U��!�D�{��;��]J���$}�b=q(-�Y�O<����_�����J�Y\Me�@{xx ����c��[0b$��Eٯ����x������'���9��,���P$�gmX(�k�F\���3��04�l[u�3�۱mcf���۳Ͷ����z�g���O�v����
`w����`��nh�㹝�#��b.iD���{��Ľ�^��.H�fe)�S2�]��g*�Ga!����ɺ� ���
$���$�A
3N�Y�`ˠ�!H��f��/�FK���$<LD8���j��w�'_9����~�V�= ����������+��ɾ��$�[�ۿ|s�{��D
n&;���O��P�R�c}
�fe"(u�˲H���2���8�b� �q]B���$����ﲜ��êP�:�[4���f&-z7z"Xs��x��&n�5W�i{����:�/��;�]\9���yF,1O!�� m���n���u���j�;rt�s]�#������v1��m��]s����w�������q������n;vgnǱ�}x�5�8Hay�nθ�\��?���6Ǵ�w]B絨ˋ��[��\�>ݲqI����]��`{\r9mnN<\j��l��ÊN�4m!�lY��/W���X8S�9���g`��z�m[=�Xݖ�8�:�{5���TB�lz����/����e.^7����ُDT��w�W�(�L!����4	[��,���~;4mH=��nF	yon�EB�&B�0���k�Y�Czk6�q��Y>���{�`�A�����gA���g���w4�c��)�w�y��|�ޱdA�t[Ӕ0��4��?_���I��;�n�x���<Opoz�\O^��N ��ـ��n�X$��!��s�RE�3&�ro��ڽ��
B�"_�Ws�Y$��5�:�]L�خj��;�,�����}���)��d=d�۪W�C��$ȉ&p6gj�q���v0��s����!k���y	�BI�㣽&!�(���I��v,�N>�h�/)�=��y`;��|PKd���"�C��"T�4�a��g��x�C�� y�U��'#������f�S��EY���\���ŋFaQ����`�?��g��� �Hx������k��b�h�&��J�*�d)�&"e#(�n�>�H�AY�&1d�v�=��ݾ�Gc�w�}���2��L��S2��<�n9D��2*��Uq&�kn�$��'ć��lcO�=��=>#^�U�t�2&d�"&�5�A_m�V���K+�g�j�� ����I/����힪3�������H�����B�m�������=M/WgR�؉��x��_����??��������L_��vA#ǟC��$��۲���y3���ن��X�I���A�����(�(�u��d��b��N�M�w7U���f�$���]�|[�2;%)��Y�,�C�l�10D@2,u\v�A&��$��m
���؟�$m��؍1@����]A��T��df�ǳ;�~씬A�=����X�������qUF<��꘭��+�pn�[��^T����h����O�OF�"b��$%�O�M�s;W�w��s�v����ͻ����={b*#���#&����}@S&TL(�4��V�I ��w�f�Ů�M9Vt��2(;��$��9߬��U$r�n2��%B�&H���z�خm����XЙ��e]�m�;]\�{��~�%�`H��}A�c�$x��9����s'�UN��,A����e@�+h� �Ӿ��o�g͑[5���dOyHy���I ��w~��'~��}$-@ē�B)�Fk�vH$��;�Ddv��s��M�����H��zA�w�X	41,dI�yghٸbfV�X�I9�V	���n�ĂCq�=�H�<�wn/�f�v��#Os��K�5J�t�痃Qݽ	�z�u���i�PP'�!?N��fΆ��丌�$���7/>����=_e߉�����IQ���Uo�vI��ЋW���-�1��b���㚠0��uj���	��a4���i�E�^�66�K�Z7#���r�3�m�u9S�����gb���Q7�w��d�{���#ĂCq�P$$�݈ �����|w��kFURd6�5����~�����t���;�./k	u�w`�|�sTIb+ӛ0{e��7�T�"`�ݗ]�B��\�=I��.�L`�-����׭݂Hn9�$)�zHQ%Q0Q���*�uO4�&>1=�b�$��mQ$�y�rN����d�=����%l����w�\��/3X>��o.z0��쭻$��Q�:�8�C��T	��I�n�ʾ�G?��g��(}N��x���B�e�&w?�k����V���Y��2��+�we\H�;b��h�P~��N@)3���$���ͳ� St/'|n	�Z�m���^yݸͻ\U���g`��B���m�ݷ<b�lB���-���Mn��Hw.w��/�H#�����۩�:��<�<����)��-�x�vwm�Z����k^���۵�B��Ű�����fp��ζ�y��,8��¦�^m����p]&�1�Z���՟Y�����ԝ#���/I�<xZ�^񑶬Wn�D)��)�)ڝt���������ی@�V[�I;��A�-�uٷ�`t)���>$oCj����L�L��Q.ü{vUqWG��;]�I8㚠	��g]�I��S��ZU�u��KT�2�`)�"$m.�I�y��,l�/�vU�!����q�Q%�gU�鵡HP"f�0M_�u��#TVL��B�>���9����q���.�@�0q�D�Fb&�C�o��}��ز��7��وA��9@�N3U H$nf;�H�|��2m[�w�����I����8�ة�"��v]�J��/����L����~l}�j0�%�}o1ՐA>�|�����f�8���|ss6��c/��IR�������O�E�O�_YN�>_N��X�UtUTS�\�uAE��u�ɢD��z�h|C���������_���\=���=��/g�Rz�
?��w�_ٟU��s>�ؿ=���\}���r�h����l6�R.�<{w�I/;ARjiL�0U9p޶�2`߾�Ȼ*�Ja�XJe��uЫʹS�V{��d�	������y[v��P]Vu�/fօ!@��bD�7`���H;˝@����7�{VH#s�݂Hn9�Ɋ�%=��w��Ѫq�zsC����sl��N.�m�.qP[����F;T<E�~~��x�n�,�s����>$�6��O�!��-8�5�T+�G�.��I�m��%d�0�0i��,����Ξ�� �}����H%�樓ӂ��lM�F�3!H�T�H����� �\У���m�������{.U���\
�!�;�]`�W��b���ؚ�^G�G�C�r����RG<��}��&�����j �Hӣ�r��0@�{ũ;=ȜS܄�_x�mM����=:~�yn�vm�s���N�kW��;�t�Wt���Z}ts�n��AX=�V�]����W�|�����Md�n8F�Fr��[��k=�|��S���Z����jX��n�
jW}ܩ[�9�����nj�`�.#��0'M8-N�6���'��Y쾼7���0������E�Iz��S<Qބ=���-�vq�y��Ow���=��A�M~ًn��_�5�UֳG������{ݷ�Bː�zn�����qbK}���D���W5 z����仼�x���	� {���f�5�o)���)��a ��ӆ��7��j}��SP�'g,�Y�oH��N\zw�Q\j�˖<��)�D�����ŻQ���5��Ы����X96"�C��6��_w{��_�d�7v�<�&U��������T/���;縻Ygʯό��/TM�znm�|�qҶ�w��;�8�h�=��V�����]X��4���3������;p�U�y֡Xa��ڭT�;rk��Τh톲��-���H��������xe �3j��[�z{ޫU��#�sĬ�=�v~�,~r�1+������{�s|�9qynk��WÆ� �v�Z��jq�TL��9p�j_#�ŧQBNUN>��`�O  ��,բɈQLTF
G-��kVڌb�T�����1R&ZV�"������JƔET�*�H��U�AUbD��B�£����e((.ZZQ�DUb,U�"����Tb��s2�+�Kh*#)r�"�b-h��.3�U���ѩF,�e-��B�,�iV�b0bDE�3H�+Q̸�*1Q-�"ƅ��A�ʅUŵ�V��TEDh�TQQEW,��h-j6��1c��r���*(-�A2���`�J�����2���(�1EQQ�r�UU1�As(�Ze���J"� ���L���d�L&-�bʖ,�*�V����آ �%�jX�Tb(�ѭT���5�-(,Q\�YiLF�Prј�-�+�j"�����Z(��J���ۗ2�30��V��Ki�UX�iE`�ĩk�
�Y�AQ���)Q�zBo_���(����ł	n>j��{I����J"E˷�(�n��l�-0�'ǝ�߬��ڠ	�fu���:��W�&�*�hɢJǏ ��y�;��`��߶`�w|gfE�������x�w3:���k���WG������w\�X�Z���D�I�G@���n��m.��:�����~~�qp�[V���ݾ�$o-�|O���v��+0+�[�v�n7�x��PQ%%1(�;]Z|ŧjU�˳k $��� H��λ����)��V�9��ޒ��S �Z`�  ����_�H5�X�$v���λ�1!L���$Poe��n�f����T>$[�v,A�|��`���&���2>Ryt��Su�Ԃ{=���2���i�Z�GcK���4��ݳ��5�;��}�p}xF"!Zs��\�Aɼx^o��#�Ֆ����$B��L�(�]��d�o�~�m�bzi�j�ڠH'ϳ�$��Z	K���p�7����6�nm�a7[nm�lf�sas��4�>:7�cjwO]���~��6ӭ�F��m_Tz�c����w~9�������<w�Zw���_��4
Ğ����c���PGD;��h@$�2�n�Am�`�(�6�Tc��H���((���!J�ݷb� ��w~Qώ�ٖ�+�*-0A�6łA��wg�p��VɅ������]�`�p�j��&o*�>$��n�H��G(���FH���誽������fAFd�(�캰H8����k�/\z�w�/n�$��:���@�{���}w��r�E��ӛ�x�7���.�<��Og��g�m�<��4�F����l�JEnOW�6�*!�=����__A೓C~{��^��B7�@!��1�#v�wY��+WG[X� qܧ�c5��ok��۞�r��x+G�l:9ku��k9��Z�&l�;�r#�7��f��Y{`�=n��{s�pp�B�5���$���=si<莰L�:�,�nu�t��ڤi��%#��0ͧ<OB�t��bb6�<��Ӯ:|q��[uٱVۙ�����l��uZd
��~i�{ٝvp�2���x�6k�mpEZ�l��(�,�����~�v�qu1
"E��۲	v�ز#\sTЧ����n�����C��Ő#FH�f@m�I��������J�@z�����I����$k�k��l�wy�'\�*D�"&B��]����A'�G[�ެ��H!��b�$7��2�! �&HJT�(C����;���&�/�Y$�p��E�κ��/j�_7�����,��z�y�� �Z�����=m���^`�[�I���H��f�&�gX�Ŭ*��u���Q��OҊ��D�Dsxש�ݍt�����Mی\��=�����������j�'Фq������p�I���`���>Gye�i�۰O7����"`�1	D�u����W�L:w� �Ozv��~}��K��]��3�7݌����*;ϰ��̮�R���CS����C��3ӱ��F܋7f��Ki� �q�hP6�:��;g��ng;7��4��m�m4��������I$��Ȅ�n��u��ܹ��$�y�w��j&
� ȉ���w}�hOaw�֭�|s��$�٘��$�����s�Q�{:�Y�f�ߎ�~u#�&��B�k]߉e�wp�m��y�.j6�x�ٙ�g�}κ��"՞E!�f�P�Ա�����)�f�\n�K�d�X�u�z"O)�3�)�SDAS8������B�#-�]����H�RV��Q;�|ӓ�	�T���k�+�:���(�b���qd���PI��ͱd��޻�|�wۢ����)���^R	���]�A �{�,���n�l�J"�z�����=�}�ZR:��=|���R����o��x��Nwo�
���vګi�J�f;��1݃�b�^i��8�h���߽}���"h� �u9u`��{��=�r�擑�6t�I�e��S@�I�x�� ���A�{;�V�Mф؆ja\�N�޻�N_o]�H-�5
���r�+;��ؿ"dͶ����n:���ܴ�B#���bz7Ku���H	!!��	��()�*P�t��v,�	��h'�6�����]��A�����p��V�SDAS���A��ܲ�#:�n�$�Ovo]�|O�>qDHj_���j�L���=Q2$L�B'Ч˜�$�/�W�6���2�;�2AouذI����=���
B��D����}K�N�t�����0H;�nŒZ�W�w�i����پ���T� �;�O|}�]ܷ��^��'{H���5#�L`��*�:�4k'C�a��j��.���C&iι��hEAåp$�u�>��Hl�����?M@��ی�:��; ������ ����B�m���'0gQATx?4�����{[�U^�������qZ�.���~qo�߉������*D�0fDPuX���Gj�B	�{6�`v�,�R	��2`;���*�Z@DȄ̕(Pu�.�Y�"���례�&Р^�m_�ҝ1Y�q��Z*nfŌ�`�(J0����B6��X�M
����N�پ�TA{vdG�Jo7�����C����~�����@&��lY'3�������S�>���pχ���V47���b�/���{��|,�.�D���۷d�NgoX�ٜ�82c6���2�V�*P�	��0tf<}�u��\A<��/U*ˉ\�5;�R۝t�~�U�}:޼B�`��4�.&@((!	0|�L{��vK�#[I`ݛY��v���q]�kz���=�^�Xz����֍K�{Y�@�����r�k2�s���[��1&wJ܎�]���7W��M�c��t��eR}��$g)��Սv�n���<p\N���+��s\whvqնL֡�ndm��(vx���f��]�^�b�<��8=0ҷ��Zg�DA-��'\�Ő�뭊�8Z�\�κ\�y�EH[`��%�`��#��l?���Bf�<5֨��۵`��;z��L'ӽ��ٌ�^$�۷`���Q&�aH='��_x��S�`���I���>�W�6���:��T"TȄ̕(P��wd�Ngk� �[6A]�0.���n'�������Ncޱg�<h�dʄL�������{�*""X!^VвIx��Y;�,�1G'���B@~�̘��SoxRaO7ެ�,�sz�kp�=� ]V��$����,��ȧ����˪qW|�B�����f�i�Ӹ�v	n-��m�ɬ��3��l��	s�ل$(�L�xS�˿	 �=�A$�w�� ����rvlP�9�y>vI� :�z~��W�C`6�2�4��D�z���^ځ��xf���#Mw���&P.A�:���=Җ��ء�F��}O]�Je��j���۾�w�}t#����6h���x��Ҽ���q>'�uݒwz�H>��$��;ą}6�2^��@���ZRv��{zH<�C�Fi�� ^=��FoK5�F\��Fb$�LJy�:��w
T�2L�yW�I�},�$���}Gi���}�EP��:�����a-D��2j�VGR�c͡�Ep:S:��<졤���E}�Vd��K�a�o�7Aό�tm��H����s�&j��vg۰�.C��"�<g9���m�	&��(�o�I��t���ͫ�9Y���6���'��5�Dp����A2�)u�n�Ĝ�(��D���v7��I��f� �n߰���jD<�z����$Z3$���H���E�E�n���������u�n
)�v­���%�xE��׹���>RuF14��d͚�5xպF(���m��s�v.�Ӎe�Vq>$k�f� ���/z�ĕb$)P�"�y���d�.��d�^@����vH$��ˋ��r_0�fb�p%mM�'�K�F"$11�L�V���rl���q��f@3��=���H�A�����5LL���<A��G�|�Sh޺�y�a+�����x�V۵<�'k���8n��dȑ
Q%�3�H���B�>$�}vLH��Ct�>ܫ��d����
L������=>Îb��خ� ��ͫ$��}b��fnš���߲0f�HHQ �P���w���K�}b� ɬ�|�e[|�����u߉$�g} >���e��i�y��_�]3���>���$���*�'Ă}��ݒN�tf<~�.�������p߱�_w��{|�ei8�Sޘ���&�g6�1�����שeverN�o�5��W��7������i1��)�e������$��J:�0��Zݗ���_�����f��qC�c*dV
\�c��Ѫ��znŉ<ݽ��iݹ/M����[qq��m,,���}�!&�,M��ϳ���㙍ݒ�΅dmE�p����8�^f���V�"D	�$Mٞ�����B��؃|��� �	��w]�@$k�f�;�[�W�5tvT8Y�X	��3 �1$����� ���'�o�:(��u��O�;��v$k�dP�ڒ"$*�w\�m󼗮��H�X�����H�r�A>n�YH�q� �>�ޟ�=C�1�Kl&�ƴ��t�>//:��k�M)Իtx��n�Ēr�Hn������Q�����]fti�e����}���Uzj*�ֶ��\�6q��N�M�U��f�>��H�<���<}�Bw�Y���j^
x%�~���򠽥�z�<�8#Q�s;�x_5}&�9#C9�e�U����^t�(�_�-���t��#�����tM@z���,�`̳�e<dB���q��s;�%���˪� �ϗ�M�2��=���p��î�iǳ3��u[��Y��N9��G݆��G��x������l��;Z$}�2{���r9,$�@��I��^7�4j�Y�Ǯp,�&�=d����]�0Q H׌s<�zv��������� t�����i�ڮY�h<p�'�7���AQK ��	�.$#Y�p�0f��u0����4��1>')ۧ�Y�Oo�Q
�^]Ȧ����}�羢Uw���'�!���^���t�jz�a���Z���zH���;,��^�tg�̚�������X�(�4ҋ�u�� �Ͷ�!+��R��;��90h��s&��T�s�m.��./Y��hj`K�y���_R��UF|9���ԟ}�3�ȹw���P���l��z�b1�Ѯ{V���[�6d&,\t�ѹ���^4�Y��{9�:�dL�WC��޾�{V���{�Ug���-ܡ��5�Cq��ӽ�b�N��,K�)0����R�ZG.��z����䒦/�����9�!���W�H��e���Z\����W�͕2���O�Z7���z���`��zjVL��D۰@$�|H ��@�/Ԩ���%T�X���be�n5Kj�Fa���A�� �*�PQ�e�LL���jVc�X1
(���XPTQTQD�R��±�m�%Y���̔��"���bԲ�e�
�iZbT
�TX��Z �J�"��,ĵ�ʨ5��m�X��Lmh�[��UTʈUPF%h�(��%�h9k�D*R�q��E���+Z�J�JŌX�(�AD`�������Ն%��⸸[m+Z�,h��E�dF�X�BڶmV"�ZV*�DU�1TĢ���m��q�V�Tn\r���KFJ�SV�UaPi`���+r�̶9E+Z�E�.+�G.8�R�-kl�XQڲ�*
��b(,Ɖ�m,Tq�2ehQKUr�E��A`�*5�XxX�{��L�.V�Ճz��q�c�7��q�m�dy:7K�WF�V����I�k�A�nnF��\D<�N:;��^e�q��z1��u�<�iyR��0�p��[Ȟ[�����Ct�B�w]�,iNT�yѬ���ƴ�[�z{*�L۝H�r�� �k�벮�t]�b�ʑ�ȏdm;��5�[�gu�K��76{&'vX�ᗵq���v�nG\k��>��..���f��J��{��og��7G#��oں`�v�d��qO�����s�y���(��!g�j�٬uš�ɶ;k0d��۝�NA�[;��5�*��!Y��uq�'ߝ�ߙ=rQ��{sE!v�8�W���=6��l�;N��[�]��c�;�K�����r]�gvi�u�l���q�nz�k*Au���N��Iok�ļ���غ�cl/6wn=��t��mOv�{�:�r���;�kx�e���I0�[c=��Z����
�n�u듰Z��9��]m�)�h8uΛ��un^ۜ�3���-ѽ��;��&0W7������&���i��pR�Ξ۱iћJon�t<Z�e6W�6{y��{U��y�sڷ��s�л����Cl��&8��C&���ǭ��Ӹ�C�Bhx��[t�q���kFB��۷Y�d�4r��u\q��ۊ�d��:y���˺��[����ne�����ܥh�-�;ii�.�sM.����Z����@�]p�g6��l�<�>�G`��m�Y�t�ې���$w]\�MS����r�y�3<�r۷��Gb�IƱ�m����>s�R�T8�=�"��e�<��ݬ��cGp\\b'k�:V��7�ړ��Ӎ�
���.z�u�=uv��uu$���F�n2n�wP��,̽��ۥ3�q��d�<���ǫh�n�k�d�Ƈk�9�6�=�|is�=s����65���Akgꊉ��M�`������k���3qt�q��v'�qu�i�B����N��=v��ռ����hV;�㓴s�;�!������oE�U����c�i�*�uw읏n��n��m���Ș���h�\vu�v�t.�(���oAq��L�i|�y��Rێ���m#
9������γ�R�wctv��t�jE6�q�G"0O�<�hm�<4o9���]�����1�C��n��y��-���z�,����ó�E��6.eܾ���,&�b��O6Y	�9&�@v-e�65K��1�$[��Z��:��~�߽��"H�P�"�x��u��$�t:D�緝v1����kR��շ`�FwK4O�S��I�m&s{w�I�uʉ�=���$���C��$�m�dt���Y�C��ȑd�Sw�g�:�@��[ڲA"TE���9��I�? _O�f ���m�,%�����0&�����7Q�;lY ���t~JO��w�;S`S/e#$�Q�j�[ݻ$v���p�?T�t-�0����w�������o��t�_�l�n�o����2Y��$��� ��b��Z�@;e��jz9�ûm���?�?L}�a.W]G[�u�I6�Y$�@����0�oO+8g+�Y�I���Eh�2� ���ZRI�'�� w�ߗuz�.�}���w��_vmA��9AoDf<�5�eT��k`R�Cl�wU��a�z�(�_ �[��it�	����>9o��%9�ç0���z����9���±6Zk7�����ސ`�݋r��-�M���]������\A�" Ϧ&��Z���י���{Uh�۽�`�Az݋$7����#k	��%/�`�]ɶ�R����>�ܲH8�5�r*:��K����y}v	���:�5@�*oDq�Ŕ�i+EGe��>X�OE[&�PM��b�1��ԯ<&:�-��l����1�O eD�='�@;|�ψ#\sT[��g:܊�ۻ���zd]Qq4�/A�X�~ڀ�q�R��v��P�Iw��� �\�+��H���Ү���?ea��x�E��u�u=��z	 �5;ZF��+�iV�0�O=�UrNx�<��Y^QԪ^A�p˭�����a�o۠�Qx�����º!X��6gt����zw�܀~�/�w �;���±6Zk7�}0g��75�V ��r$�����}��|H�y�Y8��`ٲ.{�X��`[B�
}16:�v�	%�� ��V��|-�m�'��j�O��:���g(Y�>��69�Z�,�]��^�.������;��Qʼ�'k�4V,O��"���Kϰo�d�Iƛ�$�n�vθ͋*bf�UwX�A-�j�c�v���$J�(Շv�����]�i9G'�X�H�mP �w� �����$8�3w�D���H�J��<��@&��P�Q������� ����y�w�Eh��`*"b.�w}��+�5U�|/rs+����Q$�73n�$�r���H�X j)x�v��3G�h���-o�+7o}�"ML����4���E��@���w=( 5=�L
T�0���4���瀉N;�f}����Q��Y���������D9yr��<�hV���A{���$�����̂��(�)!(̗��lm�q��᭔��<s�=λ;S��ŝ�=��������
�L���ryPI�c�$	o�ߊN#��v���֨�os:���kSk6�'���v��r���t���A��V���{y�ٱ���c 1��!""I��%�u�۰H��|��"�l4��j�E^�a�hw�ǘ�� g��u`���L�����ѷrK��G�����f�X$I�gs�� ��#}��{�ȫ��v<O���W�S��M)3�}�� /��jvN땹�b5��'�v�Y ������㚠o%�ƶgת�o|�a�/�����L��H*i�KZ�;8���m#U�}�����MN	�Ʃr�8��R��={��u�!>5��m�L"�D�
XU�C���cg�(�s=���
b�Н�6�[����M8��q���m��m��j6�rۅ|͢�c���v'{�)��9��x��j��؅Nn�r�����,]��D�opn���m�ѓ��vr霮mq�������1dt%�=���J�Xۧ��T�
w�v���y�[�6պ�,3��5��2GS�un�(M�� �R�HՂ�y�Y�:����~�~[U(�`�L���H9���An9�/��@8��qnr�x���س�x�Q!)}36'�v�[9���!��W|H'1�b�-�kΆ�_�`�ܜ`�8Y0�>RH���]`竝 �g`�{�S{�;5�I;��`���j�ûJBDD�%DJ7t���s�7���'��X�	�8㚢Iy���zr���7�,^;���l�A�n��o�/3:�u�����Iw7t,�sT	'=m�Lb��ʁ��H��)��^ QݝF9�lr
���m1��.$Mi�6����6?�?�������
$D�����]�$�.hP%�g]��y�K
!;�Uv�`�{���71���-�5��ޟI��GB�1o��������C�g�S�n�4���LG����uZy��[3{���X�a���U�`��-��B%� �u�m��	$>�Я�3��".��\��[i��Ѧb��
T�����q��� �}o�'�0F��K����pk�� �3���A#s3���=��3�R�DH�s˭�Y��seY&mNЃ�I�����~���R)[�E�� 覝�c�=I	
$�
"Q��u�� ����s���4�Y�Q"�7n�� ��wy�L�{���K3�)"�`� ��Kۮ*����i��nm�܍�mѻdѪ������|�S!L$$Lq�]u���~ ���Vo!���o�Ϡ5:t -��g�'�e����2�JA�}2����\�����E�n݂|F<�b�/��ħ��-�30�&YM4Z`4�o������� ��2�eP����Hҧ���sݶ�Τ"��Gh���8VⲲ�XQ����5��@WY��`2`bͼ�ԅ2&.~M_t��킾Z��),�����{~�<�bϷ�,�L�FB33vk�ul�&�..o,�b'X$�C��vH�8�Ǆ��������݂�DL"eHFQ�#|k�e�$��ν���L������t,��P/&Ƈ|2��ȈuDʙ1"$()D��On��������6����a�Y��]�߉!p��'{��:�y�;A69�##��[���� ��_� S+p������5�H���x3�b�tu�e?	%�7v	$fƙ"	���]H]dv�Eὃ��Q0d��:k����t�mJf�{��+�$���_���f�r�e��e�Mg?�4樞p_Oz@0n��D��ͣz��O+��[������L*�hʲ���C�f������=�/��o��3ڱ�eE���8^ tZ�{5�cg}��Y'����,m�^ ۫����$�o6�l�Q�7&2:C��v	�#[�h}�ٷ`���%ۍ��d{�_@�02C!26�4
.��/=�Y���b�3��א�:s�h-���߇œh�ѝ ����$ކhN�f�����t��L�U�����#�>%	
$�	L�s�n�qnFX�G�"wq�u���Hz��7{6�t�'�b-���˻�3�`n�6#5�}�4u��� ���TА_a��b�z'��,�$�:��u�jD��IA�罼�׸z0s��ImŚ�v<۲A �n�H
�@���^A��(�`&�Ζ��A��wb+����S�vzl�$�n�'��]͚�U��[yyr��ͫ������&��|Y��k^�K]ӽ�����gv����n�|S}3�n���2�Ȃ�&lȖ����{����}�����T�a�㞘�n
��;os����7\���q�����*��+֗;k�S��޸��غ���ug��YM�z���/y�n�;L���r�g��n�6W����B�q��\o\W�u��v��-��,�4�{=lmG��;n6�Qik�-�M���F7�,`+v������8�]G[9�����e�8�ٶ��36��n�q��ָ�u��b:�h�-m�;K�.�9u�v�t'�ߝ����鸜��|]GRo6��=ޫ��ow,@
���F{�ѿ��;�^�/�D� 2�2���տYx���έ.Q1:���6�Ēv�_��y�q��:��bps&�)�I�َ���w��.��"v��]M�$���n� ��w} �3+p�������m]�m	��l�g'�_�>$�uؿ���]9��v��}t����zz�`H�R�L#a�>vI�<�:%D��Q�F�GvoX��q����'sB!�燅�}��������e�pb����#��ٜ�ep�8k$�gp���T<E�~~�5fT�ڥw�Y�އ� �3g� ����- Vε��cVv;��/`�)8�qv���d�L��E*�p�G3�� -�[3������S{ܥ��}
�l����~�}�,^i��ߦ�I�t8 e�)���g�a3r��W*�Z�ʹ��ݲ|uU6��hu�g@^c{`��.��	,q���	��'�`;.���WyI�/z&��$���� @�_����g�v; �3e�� ��{\��r�DJ�MP ��^��ץ����8u 9��!��=�_�}�ݾ�*䊘��6s��Ԁ5}�L���h
i��/����'� $���Y��YĦ��\G�0�fU�o�@$��wߒ-�;�WB���:Eߟm��
mq�p�`H%��9Z��a��q71���ԛkl�^����|���� ���|>��3����T�	k�y��f�;�\��)�W{I7y}�Gϰ�)�ڂa���� zd5Y8�vW��LA�n�_� �����
�zMnϦ@�s���H�SJ��US���s�����j� /ߴ�}����@�8t�a�zPf�V�dO�>N{��w]��͉qݾ��*���@ٵ�y�\-jv�;e0���ށ��j��,��z 5��}�"Xǵvo���Yl��Qy�&�ܻ��`>KȘ��7_%f����w�so�=̤��k~|�G�s|�sŨ=��ǯjW8�X����n��\"T�	�7Y�Z���0xu57뻄�g�^Â�j`Ct�v(Lk9�j��fr�Ky"�Ͳ��,Nfd�5r�i'K5eY�m�TAHg^=���r��ʹǯhV�7�E�m�Z&m�A{16èw7���C�V��Z��l���Wz��u����nw��o���rI:{Lv)�5�>�p^9�-�{�,:�����T��
kd �P��� ��u2��u5��m��a�lE;S��l�u�Sh�7���:i�ܣ$]l�����r�]��.x�����-���.f��l9�'��\CY&��TC���oyUIO-#�a�G�C�Dz2��)�9��jj��
*��-�A�>���t�p��5����	kd��Y�[:��'��H�}�� -:��,��^�[��~ly�|z�Z��	���<xn�T� æ��ϨFj@�p�*�K�v�*�;s5SkId�����۹��J��x���pf� �[!����s�{]�>��O���W����jg4��>��{1�F.�ب�� 7�:��� Zq4��#���Z��[�ě�{��������.�jX�+�����NC���5�%�N��Ytq�2���p��iP�őb*�m(�*DV�-�F9L�U�)EAAAE�-�R����Ub��J,Q"�jj�-�P-�2�-�Yf8�(V.2�l��(�l��11�T�+QDk*Em�+Z���2���mC2�f-�ƴ[iBҵ�"���+���Pb�(���V*�m��ѕ���ʎ"�DҊ�֢"eR�Z�T�mZ�e���3od2�p{n;�m�ù�K�T�mj�9q�DU�5nZ��[ڭ�)���)J��b9q�T�K(8�2�CZT�q�XQ-��3-m�U�Ur�Ҹ���cF�-r��VT̠�eʵ�*ƕKk)em-k���PjQ�ڔ��JVұ���"�Z�m�ڢ�%AF
�6���Z[ZE�-m��iF�ҬcilUZ�#G)�-V��B> �B��u�� t�� ���ݫ	Ψ2h"(�(��Nx�s݇Nj�����	f+ڂM���s��@#'3���:�nw�(��"�t�r���k��H��AJ�q=�� �L�j��e�uߪ�U^ݯ���y��h���V@�NgKLœ����61�{/�؜rջ3�m�]��{����'nN�x��ێ�Q_T�PImj�d�"TOԪs��[t�v_k� d�t�����>���.�����oM㖀H��nՂ�p�e"� Ʉ��}1Ä�1�I�ޕ��}�ꂍ�����h �Ζ� A��g]vS�i��U4S1Jb*�}�oeڰ 0�֩�";��.��m���λ� ��ݷh#΋��9�蠠)�(�	��~]j��\ўS�e����h".��ڰ@�y��,���;�t6Y�/�Ga�BГur�ôo�
a�'����~oEQg�AGq���_��6N�����%��I�)<��/�'v{�Rrwj��)
*aS��x�mS ӷ�P]��;8UD>כw`iy�� ���r����gv���x���[��56)�ܕ�M��ŭ]lq�K����L�bd���A���!D�AL���uw�j�^s��@�o��Eڛ�������V@�2o:_�%��CS$�LD�J��������7*+��{��Ӹޫ/:|��l���k��6 ���=?���Rs'�Юd���`l4{�S��;|� D?E�^�d6�;K� �f��Z$�\�	U�ؓ$4�����v�_���>�A=�,��T�	fOk���ͼ�ڍ�ZU�Y��@|Lֹi0[�{>D�m�
�a��Ld�$����$�~�>l����w\��3o:�6��R����]M��*u��n̊y�ׯ4�E��n՝���7sU�r%��5��s�]b>�
��.{^�����/jrm��'f6�[t�PD��OKN�Ֆ�V��i�ͳ;����tQT��C8����H�G\GW1ק��K�@���N�q�U%�՝���<T7k��S�7�����Q/F����\v��s��]Ѻ8�c9��5�<�:�b]Bc�s����c�[�^�89����6xҌ;&ԅ��c8N�ru������]�NɞC���%ɶ�q��:3����v��,��/a���X�(v�^�bG��^y�Ͳ�����ON쁻��H�탦�"�B�EW�x�mS i��J%$���f%RA�b�Wds�OC�V�&���,%U�iL�&!O�����bA'ϧ�VӞ�ۗ����%� �gu�f�s�d��~C�>���<F���vBT�n�	��_�7 ��n��/o9ڰ@zU��=��<3���>A�n�X #6�Սl�@`�H����}8��ky�t���|���@r������]S��D:������J/'�DP%}*������봬> 0�֩�U�v�Q�D��r\�9` �λ�PH���i��\b�/\�xty�wX:��G.ۧ�H�����Ly��ƍ��S�n��aTԮ�:y���"j+G3��@�滰 �Ζ��nWt<�E?Vk��Krm�h�y���U��"��d�f��'yiB�Nv�����zO�5�>�R���{�g�V��VM�̏�D.o�Y��+��o
�?��{՞�)Z��F������I��J� /o:�"�FNgO�@��Md�֫�^U�?_C"�"j�T�_6��n/�>A�g:`Dv�S]U�9�X���LF�ۙ�Y ���2^E!�4?Roa�?Y�9�>i����a -�� �A����-��sؼ����Uu�#��^b^��)`�L�2LLAVKT�)��3��5Csٯ��VxY��e�˻�	��FoEM���5/�i�g٣���|kea!A�
��eְ�sE�DG5��Q�e�yMs��w���ߜ�K�L�o���" ��]1 �t�������)�xZ���vF��H��|���B~�~[��m�IL8f���2��FT(����w��D������s�h�l�wu��o{/�w*4�QB��8h<m�T� n�j��V���ҩ�������[v&���@瞜�`�1�yI�V�N�4��v� �^���]�^���W����ןut�#޷;¢d,�M��EW���H��&ێw䐺�6��
&R�뵾{����zg���h	-������PI6=����Ee�u: 4IA5�U?Bc��!�4P���?S�#$����b��2g�J����9l �7}- /s:�X�ӝ˯k��2�d��m�p���]���͢�h����8+�ڮu�W�@x�r�\r�"�M)*H=���>q��D@��3���rפݣ�oL]�U\�̀��r��]b�� ���H�?��}v�g�x���s�ns� �o�!����wd7;S���od�
�Ο"�UJ ��c�� �{������E�5�KIgG8��@8o������gŃ���8�8 �[�3n6�dy� ]�������$�p�yR�1��L�����gƐ�y��/V"qAصo���60��T�v������˞�$�=�r��%�S���:K2������?�]d�ݑ�)R&�*&f��F��]�`/��ON��߸���9`|���Y� ��햾d���S2�x��M@\<�+{l��V;\m�m��C�:w����b5��MZe<�}�A�SE �<n|z�X@/s9݇� 2o�[��o{���zfM����wc[+ũ"*������ ��?�������e�t�� �@}{��q��Ϣ�c��N-Q���N����S1H(��J*A��n5 ��j��4,����׾5A񻙷+ �&���gꊔTI)(�6��_Tu�U�i�j�D�J��;V-�͖�A�Ӿ3�Mz/�
�ϭ�O�}�3�����#� ��� nt�z���l�n�݀�y��d�լk���㨢)Z7ѯӋ��ͼ�G�ȟУP�
�x��	��aμ��3�79�!?�K�7�a�������1��o��aY~�g;�t�������l�㣙n�m�\l�ݝ�š	�#�>Cg�Ձ��ml[�{���7=�6-�6����׋j'�Ӱvn����Ѧ�쭩�N�ɀs��y�9�.�9��;>'A�F�n�n���Z����`��6�kZ�1��^����z��8�P��vn�cc-'q�n�r���6{[ޏ�FQÐʖ���n��:�.zp\��y%T�9�D`����ȍ��u��q��6y����k�d�\��,oD��g�x�$�a$�p羯��/9�>�լa[J=�T"Q�fuڲ�M�KL��@�5"~x���򰉄��rf�ӈ��ө( 6o:[ ޭdCA=^����v�5��Z�"����G��b ���?� �;�;�r���� GM�KL��լ`O��L�ET)(�q���e��)F��� ��v�g�I �v��K^�g:��9ԫ��M �����L�%LI)(�4�tî���3]����M����ӽ��v�� �3s:�d�/�2��(�����;8&���^�����'��T�b�Ą��N��Ř��O��A�5%"LL��&VU�� $�;� �f�u݇z2���t#�7v�EU�a$;\�Dغ|-M�O����}��$����H�f��vY���c��bd.��e�q���ee<��/��A|�u��4�����C+���K�J.����X���Bs�ҵ�0"yլ` �λV@�fu�<����EП�0>�aE���xԟ�m� ��wd@[�>�R�޹؎Ν���f�u���T9����34{Kޚ�}pԕ��Ґ@|�K��n�@d�t�'�z�TRNm��b��A�KE� �}�����ގ,86zu^��~$�ߜ� ��ͻ��FM�O��9���Y���n�lvF�h| ^�z]\6�kd���4c\�n�F�bJ~����	L.#ѯo؀ ܼ�v  ������=z�r=��MgĀL������x���p-ez|�͍۶"�#��}�7�>�3/:�� ��Ζ� zn�?g6O�8���ȥJfjb�fk���ܻ�X ^sT�/q����u:O�����D�����	[�v疃���a���wM��א�w���
E�7��1Z�f�64��QO�ݺ\@��^����	�{�!8��!�V�i�]f*̡�x����$��v�]�	 ���k�&�C_K�o/^�V���A�O�.��1pڑ$'�$� ��Mc�%��:�B펁�z�f�L��r�� 2o6Zd�oV��Y����]�~k���y�k�ˣ�nI�&-�R��j�ó��X��ڷ�ծ�o��߇ޔ�٢������� ��g�ޭc��u��}�h�}�?��nR ?�+�Z��<����Q5Ǝ����6I���
��oMS��l�l� n�����ȋ���;���J�{5Q�@��DԠ�cA�]Ϣ^��t |�n7��wSE�n���/:[ @f�s@L��d��a���&�ׯ���U��̄E���L�vNk�� ��xx�&h+t+��ځ�h��� xN��	I�r��nYqu��ڕ���6��S����_N�����N��fJ�1�=���aQ�����`�j�9�2Q*�T����j� ܼ�X���Q��q�߀O_Kh"�9�b��wg��L��G���!��g��5Irv"�����:v���GV�8.o=�ڔzx��������P3u��Ͼ��/��`�gza��n�u�E8g"6��G;Ъ�]�J�z��Bj4�ŅcM��,A���Rp�;��^��;�鋣=ܩ��9�Z@ n�}nR�\�G��_����<e��Ȁ������� ����Y z�n�gb��/� K�s��> ݼ�oTP(��h �c�(�n�zv}3��~t�[��w`#g3���95�s�p9��ˤS�&>�&���$��Է��1$�kw�M��췹l��(>�>�,"�3�Ր ��Ζ��yAߊ���D�%��sd�]s9N||0���ș;#c4�w2��K:L��/�<�M��ְdc`39h�)�<�.R/Q�3���6�v��������C�(�4���-<}��;t������zv��D��v5{����;�������'^�#�{�Ex�x�)�n��U���]&l�T��Ʒ\��;'4�ނ�������-�6�6�n4ht��D�,�� �=������F��m@ȁΗ��@ %C练��.��]�㬓�R��"����;���[Kv��r�r��Jeײ<�75㛙����sV{�ڝ��57H�j�1^L�D�x�<�Ǻ��[����s�뚁���R�ON��/���D��{D>�s�bYGc'a�"u��6浙Z�Žt�9�$`k����g�.Cy�ɽ(�ۂ��m��~�&�t���%~1�"�ا�Of� �K��1iiwT��o]�{F��4�p�2�=}�mc&�Z0��82t��#ݾ���y���l�,�u0}|^za�]��*���xu����xH��%�x?�{D�j&���a���t\J�	U+��Fz�19wE��Oz罉��I:�8=Lm���y�?m�H'ڏE�f����|���M`�����[��t\BNM����{f0�]>�Kq�0��H�y�����1}������zv�H�fr�䭛}�7����C���s�[/���h�0*󨚎-�X�s<]���u�s{]y{���-��ޢN^��]y������[��U����Q�kZ�9�-m�J�R%j��������Z-E�ar�%-�KTT���-�*cDZ���զ[1iH���-�Te�Z��,�Z�V�b�[b���Z���`�D��P���Ȍ1ZZ��̮aPʅW32��Z�R�jJ����6�e+-U�)bֈ���U\j���F ڱ���,j[P�D�je���e��[U���b��D�*�U�-�)����Q��G)�m1Z%V�Z4��c�ҍ�)h�1�-(��BШR���D��X�������e�F���f-m��iUJ幖�V�ډFZ�J(���kEZ�Yj��F�h���j)R��,���,��DE)X�)J�TJ[e�e��˟c�o3>nT�.v$m��s/d,l����l�7Sby�bC+>�wav�c�8S�^M�-]�1��܉-����z�jݱ��`[�{"�Yvp7"�ɸ�m:�u&���h`�S��a�吶�M�h��Cq��N�msU�Q����\�y����v����\q��K�pWK�[Gmذ<<���N$��d�D�[���j(�"iփ��Z-��R��[��p:��X�9�����m�'n�m�[wL��\Ap��:�%�$���Z�1rc:jۃGu"��;�6�h�:�]<-�bێ녇��g��ku�an{p�[k&^�n�s�q�ݷN�ø��\�vw�Wn��d�q��
�]�z[��2�pt��ֺ޷%Oh�����^x;#�^�lm��c5v�ۦ��򒸻p�B�.����Z��X}�=��w"�s���q��<��􅡝�:��WA9�:��o>y������k�kT�%}����5G:��lĭo+��Ǭ�㲶��ˋnk�pȝ���1�Ƽ�q՟m�.Ɩ��m���Q��ɚԆ�C���<�-�0;Qu�F����Kl�w<�w:�M�S��O
�.Ƽ]�9]��7R11�W�̝Cľ�ݹ�a����VZ�r��+6���Y�Ds�ݍ���B7�<=��n)�c���N�m�Ls����j��m���� W[��խ��N���Z�,�f����^���`�����c�����ؽ����-ps�۟e��n��s��=`]�prE�;a�v�m�����ɤA\���^Q�[��x�]i�Ƕ���on2��v�'$m۷s���o.5�����].�Fb�1�n��.2=Y��$flc�h�]c�Onг�uD�)<���M]����C�nx�;vY��2�R֢��%<m�s�8�m��Vq��x�m��sې�P�!7;`pG7(qDn�)��m���z��]�6���ѵ��\�+��-e��k�a-���u��{]�Mv!;\ʽ��n;q��{vx˺�&U�fM�Wlp�
\g�糸�ly�q�ur�Lp<����m�4�m���pqϜ`G����۷={t�uӝ�լ�3��w=<4�n6��C�x�;�OmǷN�I��G�5]�q����nÜ���vc\yɭ�ی�m���]�;�l�TC*f6R�8��nxĻ-ۇ<3�ĖC-m.l���+>�����)�W�����A�n��k^��	��ϼ]�����s�6�ͪ ���a� l�t��/�w�w��/ڽ��r�	 ��λVM��D�H��������{g�ܥ�o_s��ޘ� ��ۻ@|6s:Zd���Y����K@W��uR�U5QIP��o]� =��,A��{j
���d��Th	 �]ٯ,�p'Ǘ��.�U5Hj+�C�[��_�� '����D�i^@|��9�Sm�t�������y�g6�L-���T�EJc
6�>�_y�D�{ى���Dk�u�� ����x�y7�XOS|�߇���nd. �/Dj���XLe�Ŷ�M�9bL�4�Σ��߿���TA4�����|�ݼ��@ �;�� ���1u�C���>�ۻ �����	�h6c�b�
�*[��6�F8Ҧ��tH��ld(Ʋk�7�Z�f��t����DA�F_R�cN��3���|=�၍9�rh��B�ٸ�y����!9���B�m��ڨޝ��)?@�oO{��>���/�]VMuã�3��\ȇ��"�xl���Ͻ> Az^�b!��ڊ�U8zzg�3�����x�y7�XW��qR�U3$&ͅ.�c�+L>�ù��H$M��> }�7�X ��μyM9�s��d��'��?^*�XI�N��0�H� }��A�H�9}J��_fZ����)�θ$�7�ٞ�S�®�Lzc���ݿ�&�ҝ4����v����gg�=�v.�4{nK�w	������O�v�Q������>�,��T ��]���0�7%;g���f��	�54��iU3_6w���� w�.���{�,�S������7o:�E�i���2Qr��^	�h2c�b�
*[GX��@ ^�s�"v#9o�ʈ�����Z�����9u�o86h����!�n�����}ܻ��'^��F_��x���v��T��>���4C��]هs�@&�����[v��A$�c�` n�u�V20nfI��EUA�GǄo���> &��5A�/�5��7�gtw{�[���;'�mK�@'◱�X�`"�8��� R|n�}3��YT�SoK�/� �ξ۴�I��~;�l�m���3��0&[I`�}��k;N�8+B�K@�����O�sY��fmB���D�V������w`-����,�Q3�9�E9���[�L$o��m>� �A���c��(�+�.��Z�:=>)�c@�����H��g*�I���E�E���Ƥ�}^�QDJh�k����˻�A���� _uϫy��Y7o:���Ƚ���'q���m�I��"HJH3v�uR2��:�O�I&*��bA"Pʫ� ���qU ��&DȻ��=.Sc�]/�o�>�f��V;���.,��֪�N�{��ɥ�K����&=1!s�!v�|/�^ �b�w�>��P>)��[���;E���'f����H"/K�5Dպp�]5���]�<��s4������(M����@�I+�4����d�L#�x�-��Z-�t:H�����d#��Ů��lu�k�7]��~?\IER��*=V{z�X ^�)��r�E	o��vp]Q7���
I>W�W��&�*�����^�����ztkgg;����}�zz#� �o����z�v�L�;�݉;�&������*�
6�>> 2��5@� ��r�5����:��.� 7Ǿ��<��)�����0�)�e��h�����`�x�>�Z� 
6�>>�}�a�<�k���a� ��8��ړB6�%�|)�AP���e������������Q.�Ͷ�e�� ��}�@7�����5tz�αW�r.B�W�G2�~��[���[�ݪs�-=�/�$�y��\۲�����?}3��,��~�_k>vMC(-b�1���H��6'm,�Y��=a�z�pS��q�ʾ�u��K.��I�t�|�Xy�R�h�q�Cn���p��"�e��}�[sXW�۞Y���v/n�lq��I���=���w]��֎ru��� �h@����=�������l�x8]>�N�į��u�M��D��r������c�����[x�V����eb�#����[g�&��#u����#7�i��S6x����jaQ�=P(/���LM"*�=�������/|����sUQU�G��Ӷyx� \�9 ���d�ԔU(����+}�wa�wn��2����@�N���|7o��Y
�s���+BC�?;�ǧ���1� ��L{��P ���X$ w����^�o2�Y$�܌ۋH���9�b^w�L91@TULAP��Q��}>�+�;�O~�`|����@�|l�Z=�s��}�~$�|�E?m��x�)��9�e�V |_z}���;�")T0�<��>#z�n��>F��P{���������ϩ�͘���v:� ���u'f;� 6����,7&�In� �o^v�ql�{�> /o���f���+��d��zn�>�f� �_�m$�|�) �!0�'�|gŁ>װɂi�>^�-�D�Y۠�*�����FCE�j����\9cw�5k�}٘��U�a�Q-���؟Dzniʻ���D����DZ6s�x�$�q�_��ḂX�	bh�`L�HD��auWve�4�� ��m?t��QY�y�$o�z�/�I���?^j�X�Ph�8a�I���<,� V�{)8 d����zjP�Z�U�g�����I����h�@!��g�qi�!�m��j��F�{�2j� S[�w`|��{� +ɾrõ�U_e�ߦ'�s�~�i����!H�q��U�Mح/�8�4���R�A���)T�4�)T���޼�g{�� +ɾr�/N�wMG7:}gn��k��� 9��x�{Y�~W�P���m���@�Q�f�z����@,���y7�X7+��~��+י��ůd��M*��(@�A��)�D^��j���oEߊ��W6��@.��藽9{�MRqӓ&���ͧ�f��j̫L�"���{q��r��ٮ�ʔ����>؆� :sO%���9�u���UT�T�4����\��;����q�����n����6�O������@#g�T8�4T)��j�x�{�m��	���ˋ�5v�؀]>����ޛ�-|םn!��sۓ�V`?"������ �q��㙈ح�u��<�[U�8S�W�n����~l�鐴]��9ey e�� }�y�v�{�C���2oǗ� @%�7�X/�ڊ�����iI_6{�����������ig^}> [�z�!�3�:�+ ��L�X)!���	�%$�����`$���޻$�Ӎ�� Ь���ɼs� μ�q���E4��i�&L'�|T�}� ��� yQ�N�y���� �q����S�E9Uܟf�~��W�qi0�֧Y��%�O��T���uWD���E�����ٻ	ОuXu
e�S���9���f��	 9�;��HM2��H�3*�8k�k��v |f�}��xq\ۻ�y�` �ͷi ���{��k��yT:��r�J�	*��SS3��s�/K��f���ȼ�;����ݴgV�����b���j�29ӛP|�{y�Հ %��{�^�yysJ�����n�z\��|�]�4,��fa,��夙Y�G�w]�_����3o6����8��s˓�΢���R�ݧ<������*�f��RWͣݷ�v >3�>�� �ec�r�V�\`H��7� �P	$�yI�.�d�Lϔǌ�ߓ�}q7�{9��o0�u�n� �f��G�W�|���ö�+��]�`�k���fjh@�8�g���{��u{�Q��w[��n�A^���&��A�|<'�����v��윛��q}�Fu�}�o�v�vͷ��uK�zrgj6�46��o��}x����]�k"Y���� �,cv��;�s��6�0�[�۳�s��v��'kS5��<���mX����u¨F��O9�k�V��uqu�z��S��X�H#Ӹ�.��kn����q�a61'8n�m�N������&^�m.,;�磸��0������7�]�q��(�6��ݜ��v�*t��<f{uQG�s������k�Q ;[�c�ђz��!�-��.�3�d����`s�6�.�]�'b�'@�i���]r�y�uk�Y�-��zJU3D��UK��c��Da{�> |�o���^^�u�-B��#޾۴�	'��w4��r����)� ��Z%ˊ�4�d^�2��]�I��-�E��hu���a;��>�uDN���(�������7�L0>r�0��S�^^�XN�Kd ,���~�������O��}�{z�ǽ���|���9�Z #�s�K�a]�M4qـ�]�/֐�2������܇��D ����zZSϭeީJ}^���_�[@�9�_��9�X=v;oMV�ws��=*@�����iឧڱA�a�q���-��.���JCa,��BI����<�S����T  ׹�0W�q^Qo"���5�.I=��	�4^�Kmf�>{�������w�y}���9�U9c�v�� A.5w%�l�{sٞ�*;�|�-؞ݜ�N��}ڽ��D�M�վ=���U��ig�oyǬ��|����@|g_mݐ$S�/�|~漟۱h���T�h2�b�i�n� ���[�H�^��ۘ�����s� �r�f�k�}@.ƚ�^� #��w��{��@���f��� >�ۻH���z��؞���.�P����e��O�f��W=��D��o��3롶|my$K�- ��m�Z ���i�Q���ջ�O��ħ�,k�e�lug�n��*<�	��Bx��v�ϔ�0t��O����o��b*~���l�o�"";/�ڰ �ޖ�H����Y �훉�w%��)9[>0�S%�c	��~[0�����׷��7�� �;o�� {�?d ��^W��τ�� *���u<M4�"������@�}�p�$	��72����|�x���d����ǃ)?[U�1�w0/n�ز<s{�����J��<��wώ�ѻ�ŗ�:zdU����Rv1�V��ˢȊp���g{��I�r�}�I'Aؽ��5��pٗ-],�Ӧ�+��q`�Sb��I�{�%,�܏J`��F�'UC�خ��m]�|�Ǿ�r�;�$x��^c�v�g���}�����7:n�ݎ�+��)jH�i�~�k��wu��O2�޽01�z��s����:��#�{%�-�}nT�#�Y�:��Y �nTf0���{�2�TSəg��v�ٛ4���u/sF�g�(�̓/ �[����#�/)'n/Z1��jM�7L����n(�C<��b�����>���r3v�%-�������جu��8�?�9����|g��c�\�{
We�5���F�ч�[��z��W����������FPɯ'�k�� }�4�y��i�Mz�n�<ǈ�]wa�
��{���%��Jq�&!��z�F�\V˺U����AR������e�N�=��1=f�>��c����NH;��<~�Y��t%��P��8���B�}��pE�M�9�WaC��[�pй��o��vb�M��q�9����N	�=7n�~�xƟ*��[�d�2[.��X�|�$�'��fcCǃa�P&[�)�%kH��o/�F�����g�pdOjÔn�f;�4�����s�QqM=��WnFh~�{�sCS��~�?�*���ׇe:�ؽ�<Re	�^��r��:��Pᓦ����wV��jK��#	���yT��a(���H��Z���j�Q�Gĩ�U*�V��
���jL�J�E�������ZZV�J�iVZ�ZV��%Z̲���B�����(�Vڣ-,�Yc��m��[��V�6��5
���VXѪ��2�+�UE[���)Z9j�I��E���5m���(���j���m�Z*P�Q���UKm�[-��j�F�X���U.R���JR�U�k�piU�QAR��,���F�-������,YB�#Q�k�F��m����ZڢU�ƈ�*��Q�R�����-��smh�̨�"V�ZUk[e��J�cR�ch��ٙ�im�kkm
�J�UJڮ9��T��R�փKZZ�,��T�V���Ыr����B��M۞� �Ge���d a���L��=ʦZ8q��i�&a�K=6w"sT>���&�n��I"P���l"��su=������#ۛwj�.}Q���(��i��"7]��,�ؕ�?��.a ��Z /�X�,��DGe��f���y���kl�)��{tN��sé�*pᵝ73�Z�:������J�+����e݂ 4���@��幈��zi^�켻������~����x�A�*TyL�v�kA�U�{�j�6����X ����l ��`|�ov��}�.�}�CXSc����GI��P ���l��N_�������T$�ϹOM%���	�����9q��^#�� W��LHd�`|3�6�{Ǯ�k��'*&��*��L�m��Zz0ݤr�
�.�eP�c�8g'���A!��k>Mw��F6�4��DdK����ӻv���)�}��:��HN3�U2�ÍSL�2Ӫ�N�,���uƨ�9�-]�>i�fN[�� ��ۻ<���������^A�&��� ��v��8���h�]�ǭ�%��d#}�����B5pTa�F�?�� �2�0� ��ۻ@�j)b%��ٿt�� ��g-�@z�cm��lcƃ�'�_u��&>'��d[�D�e0�Μ�- �3�6�b($��f�u8��r&��il��x�ALV��v��I'��z@$)O%>��������r� ��ͻV��e�!�q�	�����7m�� ��fy�|��n��g7�b�;�-���K�^[�ziMML��UI�6��݇���7�j*�^dϩ �^9h >/�6�E�i���U�#-�Zu/�}����.-�C ���e^.��=j�j�k �M�XS�\�xW|3���F_zq���°���wh���P1VM.����H���!����ہ�kI�sfvcnZ{G#\Z�cv��*��\�Hv�%�Y��˰]4�66��n9�-�+��<�pf�|�&q�v�m\�;��p���Ź��9yqqmO�ĉ��7 �kW#s��c�Q��k�%;��v�m��#�#�\M�gl�}v���2�Iu���n)�\��yb絎rN%�z{�����*dc7:�N�+�YЀ^  ��磁na� q�5>��I�5����&�&e4��zI�4�R��ݜ	־����)�;i뽍�.�fO{�������=���%�%�@�ݛ�z�9ƵKC\j]`�JIv��݁�����CA;����f�qg���$����-��`4�����H�o5L@�u2�Ocvr�����n�#Mޖ�|���: �
���"��m��r�}��  ���v	 ���m ��s����{dO�P?_����ճ>A��	[ԟ��E~�d���ڱ*��ӳ�o�_��J�^�fZ@|�[�dy9�b߻Ь��O�~wXRj��@��{N�sZx�06�����ι�����!65�����
H)>z��`�#;k�È ���,'��S�r����i����&�TK��bCG����?=��3��k���:���9q<��;[����ܼ
zX��4{=1������09����	�'���[u[��i�^F�̺wYvy$��t6� fNc� Fo�Yн0⽾�J�w��3@U �cA]Ս��3�P -��bvz�׈�Fn��� ��]�Bz���-��`4ퟎ�n���M���D>�Ɔ ��zs�x-�בD����l^�AԒ�t�Ȓ�6 ��&��*�Hz^�@�A�ٮ�ڬ��S�D��O=��	 �'1� ��ͻ���U���듢dN��u�������9x|$3Z������;=�����y��߄ѻ�U2AU
���[���2�Q$����	9P�t��o���v�ز	'����\�r-<e��������v��-�WX��ܗ�2����~��'1��ݛv��ટL�w�K;;�_������ibaSLA3��H�$�����k[�)����o��3C���[��F�����o�O�I��4(�9�V�2�-��U���Z�MKﺑ��j���������e�OK�������1�@|�ٷv
w��h��*�T1�wVN��y���v� �ߝ ��f�����:��/���xx�>W�'��m6��DL�|�Ƕ�nҰ@ �����tU_�_NB��	+q�pI6}���ċnx��Y����;�U� �������
9��]k��A*k%;��t��tgc�܍[�tvn�߿�<T$ER������ s�[�p$�u��$i�s�A��QM5���#��mť~�xPEQ(*�L��N�zՓ�,]��E'U��I!�����F����@o#_�P�'@^^�=3J���QUI�:������hb �^Ng)}\V{e�@����j� F�����ƙsL������p�i���..�Ǘ��޷��?��o�	�{�gL��;��58�ӃTB������OpzΩ��t��q�3��߲�p���]D��7���B�=��S-U���Η��+!x)��n-WtE,��b��AP��Yh ���pܯ��bm�J�=m$�$�o� �3��ﳴ���L�fl��X�g��άv�q�p�9Y�n{��'�C�!���USU%*�&b��=��w��Dq�Θ�@+��r�Dq�^ˊ=^�g9ji���PH��E�H<���1I� �3eҷ[)$���y�˪�qҵU���P	 �wz[�Y��� e��M��ϷR_Aٕ��,��	a-�JD��}>h ���T4�GV�v8��) �>�w7�:��S fdY�滳�^뚨x�eQ��-Wm�L�f:i@����3%1g���	8u}�O��Ԃ���L&���L`}{�Ҳ�}����}y���ܶ�3��A���FQ�7�
.�UOXy��5\n��M���w��]��7��
�Jmb�^/��|��uuV�b!��.�����������m���߂�n���v�K�Π궄ۅ����	˽qn��y�Oh4&�G��N�x� ��e���c7[�4k;��%�h3=�4��n��!-�c[��Dm��q7ik���{���y��)Ap`L���%Ϭ���6xj�]��s�E�����ۜ�q�T�������״�$�,��svy;{3������:�Z�����y.���:{Eά;��Cg����OG�7O\��ۭ��<�l:�gr�W����?�|X��ӂ��j��Dn�t�;ۻr	�9�3��Oc�L��7&�����[m�^&JA�����r�/���kK��1���֩� �/=/� 3��� �'�-���;7V���������&T(�� �����n� ܾ�X$ UW�ӧR����2o���y��C�Hl���!>2�;h�@b���o�� �ѹ�A�D6���A#�����`�`)g4Iq1��$�N�Ԟ2��4�	�}��ܤ 8��G/�*ݚΩ��|��M�h�7o6�Y I-��ie�M�ܺs���� ̈2����k�җ�95d
�zϣJ���;�n�gn��w�-�T��fB����T�:Ѱ�I�kw�� 2w:[	݉�͓�z���u��`��v���{*[�LЂi�
;�|�VÛ����/��WPvr�h�`$�w�4�Fo��s��!�TP%:���;{���9��;B�:*�+��1>y���S�N�o�!� ��:�� ��Ζ�[sZ��֨V���Wل��_i���/% �Hs�˴� 79�>A|�����N2��ٓh������#'s��[}��	x1��a	�����L)��d���݂A�gO��7�|zBG�3q��J+[�9tf����1 ��D�;��iy��芳M���Y��m�n�#vs�� ͛�1�8��7��?�,!����,Tg�����9:��kx����s;�δ]��	o��~���O
D��G�W�ްR@�}$�{�����QR�s\c=0��VA��w�d'H��-,Oxbw��L�@&�'d��fw7�l A�9ǟ� ln�_�Ib�	9��r�k�]s��W*[�LР��&�A]=��g� �3=0� �M��s��y�3�>���qY��˵NUeK��y6A���`[���-�bK��u�FL��BG<����qBؿ����M��r wV|fB =��$�_i���/e�I�=������qn���\�� S�jX���r���ε�Ν���}�$���3!=}�$K@c)���Z�w)$N<޻=gH�H�6'+�/�W�m �Y��������S�F#�6`5��P)���M�I,�h�j�V�V�u�b:1m�a޷�魝f;��~�5�^�T"_9�r� �3=0�@v�uݠ���S�Fԯ{�i�X��>�3����~�<e2E��L+�ﭤ���7sEz��tv\Y$���qi/$�o7����_e��jӡ���%���^���w�����^���I3;G�K���xw�{9�bGm�7�����gl"����bx=P;>߭d�o��%�5�� ��� K�3�yZU�%Pz�/x(�w}cO���ٰ��}Z9����w	��{A�{��#v��#؊�8F��0�-F�ҩ��Ge��>�Kk�@O�~�m�_��!����Ȁ7g8�΢�~uQS��;�1�/'ٯ0b)"�o+�nM;4f2KG�����c���Vϩӻn��8Lཝ$m�&"^۞w8�Hk`���?$�@c)���F����;�@�YÈ�tLr̾�V8�k���h �y�iX���ō3�l'�_�(}O��=�o�7ب	 �o:�""��� A���_��f��?.$������H<i�8h���ݑA�9�K> ���X����h�y��- ���s�-,l2�5�w��]��\�Y�N�����"���7��9�n}ۙ��������}v�>��o�3B�����_^�P��{���|��b������ tޞ��e����$�	'�$ I?�$��	'���$�HH@��B����$����BB��$��H@��	!I��$�	'�$ I8��$�BB��	!I��IO�H@��B����$����$��B�`IO�����)���]���l�0(���1w�            
 �  (     �(    +�       �  �(R� QA@P�E�dJR  )T�RP@��)PR���U

J� UJP
�

(P�             �             
 (      � �  @   v;e�@ � ;��A;�� � 	   H s�  l�&��( P%� �:���W0 ��  2 d�Q�X!� c � ɮ���9;�5��j�VH P=�  |         ��Ui�R��˝���)�eJ����oe��Ǽ x�S6<�R�f��j�ԺT�痻jզ{���)��V�NMt�T��  ���c)=�yiJ�a� -PJ͇!�k��r�ӧ"\�t�J�d� v�"Yc�T��(�UWL�\l��*�� ���  ��        � �i�eUto{A{�(uJG��zδ(h���x�B��X�h
C@sd�se) .6��gAAJR�x �m� ����hz4��BP  � ((/>�ג�cK�p@R�� w
9RAK��{̥(�0��:�u�Gze;��JP^\ 5��R���锩�euj���!�S�v�ʰh�	_  �     =   .�#�.�0e�N�Ū]��Vcsj�*�rU)��6�6�m5)�T��m��uE�  -�@+�1@
�P .�z(2 ���@wc�  $ � 8�  -a� Ԩd �T�RD��  >�        �@9�7`rv �na� ���W09 �u�� h&��2�(
�{�  `y zs� :2�u���3����� ���@t� �d |�T�"b��L�F@OɄ��$1 ��ʩFT& hT���
R�  OT���@ � 	55MJ�� jw������l*�?»����|~L�b��9���:_s;���B��	���$ I9!����IO�$ I?���$HB!!��w<?����u�45�?����ܻ�O���w��=s@/Ik�����\鑜��C��3���ʎ���@��*��@u�B^�Xz�@�fӔ7��+�٣���7i�s��V�X#y�چF���۽N(���N%��P$��~�{w�:�1�Oz���X�u<z��8,2�Vk
M�qo'^������r�BE���j[Ϊ�6k3L���n��咳]! ����U��؁�8t�^\t$����,��2D�܆���>对֨0�l�R,�]��
,z�75���C��v�ܢ��.<#�� 3�ul5��v��vd��Xu�I�+�{�����wR���%pCw��݊� �>���(H&U�x��,Ӕ>�b�*�� (��!���i�Wݑ��u��N�7�EW��s�SI��"�g0�tR��^��[���X��������H��O7ƴ�W�ە-�_H��3��ʱ�h3w�m�0(�5�U�M�0ol/��e..`n��)ݼ�e�<V\���QW%��r^=��S&w41����ʎhͭ�����G^:[Ðc�9ѻ��x�K*\����y��'s��*�ś��޸�k��ˮ���Qx�W*Ý���Y�K�nΦ�ͻ�6�ރV�P͚+��!��6��b�W���e��Qk��0a��	f�Y�)G�[��}�U�\a���-����5��)t������,'����k �&e��w�"3�.]�Q�8��w{{d��i�յlcr�����5����\����2&�M�����1�a�pH�x�T���Y������V{\x��.�oU�l�ܚ������0��T�����ۋ��B�l�8���d[^��rU�à�������7b��v�ȕ�+^��)�Q�r���̝����e�*ʆ��0c�{��ug���vq�r4�!bg5r����R���!|�p�
;��p������KĻ��`��S�Yۋ�'A��U��˓�6
�oL՛:Ж��:a��Is�����fi]Yc7Xd�wf�`ȨS�����S��k��Oj��.nv�s�X�w=ˏ�_m��q��e���7vlA�s&�.�:���eɃq٣owE�
	�M�e�q�R��^�;�]j(K����Sчx\�>ː���zU��F���'!���Ox+e-�h��R�֊h6wQ���p�a����� �[gH����c�f��/)�� l��'�d`�t��q�#��/Kk�d޽�1qn�{����/��2LCh��vkO�k�۝z3�kws�.U�ڹT��pf�Nwz�Fl؎p"� Jv�ޘ��E��f��#VE�}��ܢ��x�d�T���e�A7�;�34�m��w4M���g(�5�F�;S���{v����L��=VL=dc��J�V%���ټ�)62��p����^����YXZ�M�ú(�!�҆8x�ω��T(}�q�;�������H�Mt�7�z��/{{�윻^�p��(�i>�7����8Ak�l��4�Lo�qq�\����2�a��r�T����+���ô3���n��@�;��x���b��:A�븇1���U�.����$vhwa��Ns���&�y-to'�v��n���@j�� ���w�3H}���"v����Ǧ.�RG��=���Huỽ&�ڦ�K˧!�Y��w*�x\uu0'����r�vo)L�睗N�V�A�§iX#�u�ݡ���:�1�$@˵�X[�u#ʖB
�]P;��F��*��0b����mFU���̓�N���-�f��(��c�w�4���F2�ޅ�˻~jhǥBz�Μ�]"�nEj��֩�&��H�
"�����+�z�ص�= �Z�h<�{�)�oh*�;PuhǶ`f�s�ћԭώ��Xe�2D��67J��{���v���uZ�� z��&X����H;@������!3w�],P�}��J�P��=qt�`d
ECa��t��������=�>�^ ����4ź�/:��L۽�sȎ�N�H�N���5 �~N>��sIf!:a<0J;:�U�V7�ύ�D��V�X������;�=�{�tc7�i���Գ/�A�F�;wp�2LvE`9�r�7Wq9�2kn�`Nۇ�t}򛳻�_t� �݋s�q
�w4��#nXN�D3��滪�V2-l���a��gi�&���4�]���MX�wʃn�X�4���e�T{s���O�'�����D���Z�mط`��:&|���ư ]W'�hؗgX[��W�#���a��-�ͷ@ቼ��n�0�'׹�q�a����G�9o�\��7�:P��Ѳjҕ��8�2�4��Jq�;��-�:���Tp2�"t3�}��;e���ğKZ�q���ɳ�=9�j��a�7z��������cu����_iZk�L`i�]���O��u�-�����Fln��xD,I�����؃��Ј��O)�C��L	k��wF��NZ���^�}VV㷱;��;�Pd�U�}������k�K�Y�c���.
`���:z��j��л�ш8�:�ޓ��z�)��n�%�8ǔvF��� Eu5X��92X/uNV�\�ϊܦ�y�)��E�I�,�oWi��W�7%D����'��M@�K��f��@q��~I�yv�Zb9�O�u�JWGՍjR��Dú6��LgIt�\��w���d�粍�(�L%˛ouZr=-'.��-IcΓ��ػ 8�o�2���r�0����Yi ��4��9�S($�ZE}�<��VB�X\��_$��)'VM�Yu%�-1�Y6�X�I����0W�-�����_^�V�����"L�wa�u+��A�X j��{�;Gf�I��"�n��!��{�7�w�|�֏k��4%���oB�Ô;GD6�庹n#�]OV�ù��ޝ7m��u=���_9��z��z�;ѩ�e�C��9�cxT�Q������Z����,rn�ٝ�c�v��3��҃�ѡ�������E�N���Օ��MTy/N���a�Lo>����}�ð�m�^�^�>����07J� Yǁ�����w)�A�8��āx�Z�\� w�.��` ]�8u/^�ͫl �;�Xq���B!��A\}�H��3h���ߦB�m�dx��4.������G ��]�U�XԲ�1v���.)��S��?����t��l 5)��+;p���M�<=�$-���\%�n
�^wdIM��V���RS ��%�wMc0a��FF }���=������b�Ɗu��a�*���v�}�S,�P�"��8c�{}��㐳׷����#�u���؈�w��UهGdb�XT��)гcg!�C�^	���(y.� �RG�΁ X�@��˽]w�}����̯�|���n ��k�{� h2�b�ڰ��aYO�"�{'W+;�%;�F�.7Gu\�-_o("�{�r;�T�Q̛\O�u�swg$ޘoK ��I�PwJ�Q28<P㠤/n�	�wf��p�2�D�d�x�ٸ��-�;�*�V-�bG�:��O���8{���
-;�wS+�]�a�H��O�Q��WS90���/�����X�ys�+��F�#e|Q�z�`��m�:�T���;�.�������Ƿ��-�w�$��ǹͼ( �xCoUo��V���1�֖kѻ���bէ�(���	��Dn�ձa�����
x,�Ms�c(&;gPsb1�^�z�&nn����+��Y|Gs�G�q�O#�`'�N�Bd�:f��Kȁu�Mo`��V�f�&A�́�U�v.:�����<e`c��V>5vv�EV�է���.��#�,+\B���I�M����f�Z��
=��ݣ�䄌�:�*�rH�Ҳ��,�ʷYE���������'uNwm�����V-ףj��+;�Ϭ��7a�K�6ѢJt�-|����������4��B�ɹ`�tU7�{�ϙ��ug_6Hz�7u�`�i�/grcv����7D�{��
j�2
��@"&���pe��R�*:Gn3�L2��9=�k���Wǒ���Kq���kL"(�獢�tЊ�3eԘRq.��.�H�o��\��Vt�Y	y��1�̵��i�g�x�-j�wj�d<1��x� ]��]��'�����2�	9�O�@�A�Y�.�����y��FU�x�f^)�?*!������!,E! ����7ܝ�L�q.�7C�R1wu�����r�u�WqQ�;�b,�6#x�*��U��+㻁��SzM����Z�6����;�:���%ּ|\�Mph�J,vQ�;�����sW�Gd+ն�o�w#���5��N��:�ӆv�ZE��_r�9C�4��uꝝ�7��F�k4�^t�}��|�y.�7�)�ٽ����6�c;���DX�F�y;�.^��c�d{�X�/m��f�>kh����0"l3�˷x�����`��<,[CP�Y޻� x��4��B�1�ۣ˦3d��]��p�U��QOg�t	��|���%S���
ùΔݘ���Ɓ��"r[�b��C�1���^���G�&����Ǖ��ըV�p�Y�_�����6�W؅��\)%���qweT�ֻ��]�;�^�'���+W�gMJvB���	�:w 9GR��o-��x��nh=�h�{�	X��6�݆�%8ȒUu%zk���rs��
o�,L��3ƕԻl20쿈)c��T�@Y��@rX	�c�ٿOuLw#����}۸^�OBh�wd��|�t�h�q�f+��6�k��8��[�x�ܱaJ@&�)�\tl{�ؠ%{���9�0Z(z�D���6j��2Vg���>lS���i(6�[�Q+�y!=�B_p�^����y�p^���dG��1���BUR-�j�&�:uҟqM6zԖ<黧m8��n��f����k:�X�\��(���U��e�u7f
����:v
��pT��X��*���x�1����P%-����l6o\�<
R����pU�477(��9�\��x\����5�[�{-�%�{5c����'Nn��YƬ�зz�B�����^�0�&���j�Tef�]��4�����p4���/ܹ ,b_Q19yd$Y�V&CG�dp؎�(�o	�����t[Zp��5�2�8+q��n)�sHH��ab��ce[T���Fdx��!
Scc���Լ��Ĝ8�Svx�ܓA'���:�sq9�����k��B%��h7�>��sH�e�Y�x<<@Ν�O>��wv^!^N���q+b��w0oWl�p^�iq��[�gk�c�.�ɘ�i�fѭl�x��gn'G';��eX9Z�A��٩NTݝ���h%ѝ�s�zrCN���`yl���*<�m�w��96�=�wP�*O�ɑ�ΐ�^t���i(.�i8�v�;E�d%E���!i�<䂄	_�V�u`���%��H��K\����XOc�;o�����T�zn3��Y�;�h�i9|���݀bt�3 �:�屽Z�}]]vR� Ń�H����݁�9�;�\#P#�y&Q]��=&,Q�����%`�UA��.�r��q�1�� �l:¹��'|��o7��n?*���H�0I��U�A�oK��b<��t}���G�r��`�G�>��f�z���='Q��b��a���53�ɐ3^�g.��sZq��36�H��Ր��f��,���:vO%�n^�O�˶���c&u{ v��b��{�p&2�#���GN�]WRpM�2����foI�㡷�h�gAz�ox�;�p��0i���h2�R幸�e�l��U��ydLb�e-vͯ�0`���K�s!S����n�n=�i��g[�dɉn��Ų���c&��g<��h�hЖ
��f���o(��˺v	����6`n�Ņ�bO�^���JY,I�W)�Yv���K��G]2��wzQ8ۣ-GdGQ�ۀ��f$��QR�CHI|.�{�*���K�X�9�e�ix�u�Ct[�5N�����ϒ��@ݗ����ʣ�#V�[,�rݏ7�]ñ��[/7�뙷�/<�ziW��3ݣ� g|'<I��ǅ�3G�]���A�Z�ǜ�B&�ӥ��P`��;x'y��]'�p-�۔�ĺ!��y�P��p��,Pٸ�ٻ*������[��ݗ7a�R���+R�:�i��ǹ��F��{�l9�.���U:�4��*a����jY:��Dpt�f⽀����>J���⒘	���w/�<��E1-Gv�̷:�b_�7�p%�L�N����nI��Mݣ#i����r���uЦ(ۃ��9�n�A{:ut�p��/�, �8B ����ss�X�N���A�]`�X;�6,�-�Y��q�*�a�([|�t7r��rmF,W��MM�Z��LԻJ���+�*%H�����9w��!���V9�ȧU�E",��0�^�&<�J��F.��\0C�P��RMf������UX������VƵ��Ur�ح[���\��Ekm�-��Uʵ�[jŶ�ڨ���-�����Qjܪ��F���ڪ-��Z�ZڹmX�kcmTm��[X����j�Vض�lV�+b��r�6�5j*�mm��Z6��r�-UmsUk�V���F���V��Z�-��U�[cm������U�j��mnkm�[Z5��m�Z�ִ[h�j��m�Z�5j5Tj��V*ƭEV�ʭ�kmmʪ���6�s[k��mF�AV5sk���cm��lm�n[[�h�[�ֹ��ի��U��խ�{Z�mm^����.;�~����*H�Y����j�eyo��t�_��y9N��{���^���K9g�tÌ�6 ���,v�|�$
�y]"_�yz�BF�ts;�U�'R���`�%wn.���a!�b��: ����Qҏe��;N��X<2׆��mKK�V�7m���҉Mbې�猾�G��nu����L�È~y�H�0?z�zs�]�μ��.M�qz�vT�DC�=ʇ{�����<�1��ɛ�/��QK�7����*��;~LL�ź��L̏o�OD�G0�~�.x�l�x�����e�hɋ�;jѤ�5 TO&�x6ާ\���-�{���9���mn�_Z����w��ݨ.ra����d�f�1%`�S���ѤK���eH�jN-�`�|�X��sVj��됬��u?Y�T�pc\��vOl�����m�����j�ܒ�t���vov�>�(���w>kiF����ݚ��Z2�/k�ߟ)�����<��]��9�燇��o}k/?q�un_y��ӂ�{�������=�z���3{�)p�������i������= �8����W��q�ڜ���;���ys���|�=�|3}�p�+�y$gf��'Gm���k���?��*j���됂/lf�rL�Ru�� 3φ�W���e�!��g�3h?V��������[yf���=�AZ2�{���$���.s�^�",�bn�|!�vЬ��Y�Ī�nw���{�=2|^��3{��ȼu�pn���Ҹ��5'ּ��цv>�܆�3|��G����Nd���ٴ�<��9�a_����Z���:�u	��e�lz,�����'��X��� ��o�SڑM�-����{'��sί�v�����{^XCr��^���U=uVQ��6�%tL��F�BL穸3�<������y���$�,�u�A�p�;ml�j��Cv{���5�U����\v���_��51����� #9����[�靱`�{��+�}]�.�c�n��P���f׾�Q޼�ݽ�>ѿm�8|L!<�nz�B�d�m����e���˙�$	�fW��@���ܒp�d8�}�L��v]=���<�?"M��^J������D܈�ȭ�9=�2������9���g�ܥ���g���:�ǜ�X�6�y�^��F�{~�;Qh8|uz����y1_�{no���Ԡ�gW׳Ug`x�e�6������3�P������<�x �{�΄�N�8��PcڷFLc�����5�ּ�s/L�2hƱ(�!��w5a<����l�ܦt-T�m��wm�c띞(`��g�~p��
�����A�Ĕ�U9�w+sܵ����cG������]Gf>�щ.mM"�R��6����pml4ߜ���z��O�9�T���q��A����m)gxL��{Bv�G[u��e^]y�>g�Չ�=�����ԍ��ޔ�/ۻq��z���vu�E\ %�;���O���I�s��2����� ���w�C��b�Eo���<�q�:��Q�w$��m�f�NǓ+t���W8w��6��fN���N��v��h�3��O�u�y�I�xx[��[�^���L9:�#������^�fk�{D��թ�o�#���ȩlz���2N���ڽ��Ɓ���M=G�7�{�zՏ���ǔ�9������:�~�1��q]y��^r�3תH�״�$�"��͚!��nh�@�nST�o=h��m��!�p�O���e|]��riM�<���<��x��f���]����^뾾>����4��vn�G �/F��v�T��;�.ZE�6̬����J����$�r:-�%<�{�}o�cWݗr����b��^xe���ܛ����� g0�y����E���a���4J��ݙ:N�Wc��;nt)v�o��\�"�1'Y{Hd/1���ǡ��,��=�*b�PO�Y��=C7bxn���#Ŷ�������L��z�;&/�Q�����j�om�7ܢ��:s_�}���vz�z=9��Y��y,�g9�<�knϽ;�}�%_x{-�������Y�y���o���~M���ܙt=s�aW��;����ޗ����si��{ޗ�@F�	��x<>�n�5O_ ��u����G�,��p����q~*w�c'�7�0�u�$JwW�Ji��>��ܒH,�gz��<�M�U9ټYGQ����L2�{�	]�g���9yoV]�����9Af�׶��ͅ��q-~�nt&l�<�+>,/qJx�]���S��;�@�>��n�p��k{DF-�o��E��qÏ�ӚibB���yc�%û�!W��������̠�hg��CO�*������ſ{�%��8�w�3Ж����Q�h�)KX�t��[Ssm�M��R�bV��K����ADcɧ��%�'��
o�cv�sZ�swU{9���3�������Z�ĘZt �<&ɳ�yt�0;+�n?6|�{���Ѿ{���)�G�P�߰Xb^mfP�1��t�4���kƾg�R����ƨz�ry��X#�~�dx��Lע�sĲG�,�oAݩ�}u�-�'�D�U>7p���2ξİSw��<)�OZ���!�XloN�˨{�ǅ�N�r界�Q�.edB�v+���ᡲyu���q�ްnUV3ӟ���H~y�,إ�]%+��+������Ng���bK��E_�\X�뜮�^���ڤ�������-��q��m&t{��n��>'��\�h�.N}޾R�2`6^��E;�����P���h煒3yt��5�Q�r���=<�D�M��-�vh�]��9{�*ۃp$FL� f��Q��}�^��'Zͷ��=�Z���� �$�s��^���r�=e3�&;�k��Ŷ7PyO%��cD�<X��W^�� �aLƣ�6n:�4T����{/>蛰&���8_��^(+E����}��oxP�拑y�z^H��2��{�Q�e2_Q��u�*�I�8����\��]"���#�j�}�r\}����[�l�K�׺8wo����}�<��n����u�wwOn���=��=�X�4�n�����ag.�^Is<���1�;�F���O��o�}��l��?c������������)P��2Rp�d���4L���xC��&� ={���j�փYDb���@|ץ'I���.���.��{���UJ��ph�h�r����n;;��.P���&�5�w=���3h��c�qn��-W�{fmi����'�}��qy������\�(+6f�Vؕ/���|��i�z-=�{��n>�C�:3�==T�ާ��g@���ܜO����Y����+���<�n�Ո�ޒ��y�E[�Ek����x���z�1����?7ZK�מ��83�	�����Oz��>�fǢ}imb�65���$�!T���o3�kV��^փ ���&��*��m�=04c^sξu��^�qf��1*F"���1`�4Em��^���E�u�ػ���Ԯ��@Т��r�S�S�3Gܳ��z|n�zm�|%�-Ó������ ��.�r��>�ԕЙC����F�}8�[�8�7q�~��fb�Ax܂e�X��-�3�L9r���x��a͛�Wg��DːQ�,'�6���o� /.L�:>�����E��*N������������Ҏ��[������ִ#T<�Y5��~�^{�f���FIx��y�3@��9�Ĉۂ=��u�{�r��p�=��nC��vpI׹�p:�o##�f�����E�Y�3�f͙���`E+ۦ�$�����̙���/Ti�o�f��_�u��wE g��q��w���L<�G���U�:<��ԟ\�朞�6����4I����>Y��o�����l�����vw�~��vi�<��r#��i�NT�o������D�E=�=��b�yV7H�Y���=a�����ok�w)��m}�O�/O"�}�k׿D	�[a�`�Oi�6S��1ǺM�ڼ�n
�I~\�Qfn V}��%�6̽�T�r�������f[��Fޞyp�ѽ��,nr�Y�L�ċ��ɬ=���-�n�{}yi����tս�`��{\�r��yL�{Cx��=qJz}���A�/1-�]Zy!��}������w�O?���\"X�����.W��x�^�{@e�y��w��e��ڙ�O��~�	�e�wV%�t�:�Rt�S{�R��[��Lz�}�`JnH���{i��+s��d��yiyQҮ�:��Z���sh B��O%�J�O�!�:�u��6{o!����z=��;�2�G���b�rӴk��|C�?4��~N���9��O��L����BtA-��Փp㾨�d���@i��j�p�(������p�w.��zΈ��vO-�+�[;g/wx�0Z��<�`�=n�u��˸�L�,�K���`Hf��%����{Զn"�¼�vuiz��	�Ij�>#��$�7�����̧��U|d��cȶ[�N"���-l��q=�dF�����A%zb]7{�����}������t	�=�,�3]`�髆�f���������Ø%	яx�����ټ��c�i<�#�|�MU���㺎߼ކ3����5�<_Q����b?y���'�<�ۈΆ��������
1Q4xF�2�A�'z��3�bx`+�b���n�=]���lJL�����+ཌྷj��gT�V���rX�ڬ'UW_g'�c�'	CY��N���@ǻ����r��G��9���1=u�|=�����9����D�l���aT�8u�;��-�S*w��'N��N��=]�yh��E����Ռ;��B��^����?����Z�}l[��ѽѺ��`X؇��B��t��X~�kt��a���/[�ŋ�ǽ���t�H���^I�7��m�9��jNo��d�}��x��{�mʵD��
!�FL݋um ��mů��9<�h��Q�C&��7y�㮲m�
�H}��=y{e�ܳ��\G�K����h�z�f���ZrL�����=����zk�bm�$�����eq���i�\x}�<w��m{֞Kku��5��a�|lLΞ�.i[�8C\�.�|���^�Fw�������{�,��������(��j{����i�w��V��y��;a������<�>&�z�xٶ� �%Ȟ=і��`����y���5�N�{��p�v�r�`݂=��g�Y�w/z�R�2�ř;f�Zy����9e��1���j�^��]�'�����-=�_{�G���]�Bl��s���p��C\�4��0+������:���������՝��2�o{f.C�>���f˦����f�����>�Ƹ\�E�/�f��7w�i�7S΂礆�]�ܧ�yy��K����ţ��nX絊6�*O��������8�������v�ΰ�2�c�,�0g�J3���,G�XV�搞T���\Դ{L�������[N���,���mB'p�	,��3�zA��;�/'�U}{��I�;CSuE���:��V�Z���iTUe=��e@��k���x��d<�x$Y�z��S:��e�����O�{��A|O<x��V�o!���릥��&��{�;����g��ݗ�R~P���f���Ҫ�z݌mɇ{Ge��*��Ű�.�W�:�E��Xg=����N��X�u��7�Ì��)�Ǫ\���l����7p������$(o�D�Z-�8<�e3��L��O
U҇�2W��ճ�Bm�o==},m��>�a���σ�ط%����Q;�����T�a<���.��[�~e�����o˷�VI�ث��r�k�L��.<]d��@�n�`;׾��PNn9��������3MqU�ZG��|K�Ͻ�[mu���j�	�џjo�p$SGb�a�w��w ��ϖ��r5n���<�,����žY��{�z�7���c�t��U�/�f�͇���voH	jF���Gyv�����v�ta[�������dxy��8�%wܽ�5�Zd�6��^`ר0�i���+*����=9�=-\ϻ��8��Nu��7+%�����VŰ4bH����O�E�
�v{��4��{�S(��ͧ2���3.`�D��V��Ue�����sm����V
�{����G{��;��;�Q�Y��O{"�"9�xo	e	l�#����G��ܽ<����k�kO�Էhژ����|�F��ף�qs+[�����M> $���B^��눡���0�13כY)�Iv�.]���%�1A���gfދ�s D*�Ρ�#�@�8�.;��ޠ�A�/s�}�tX�Û���m��@4�.��eRe�_=^R!�
G�b��2zvI��˝�U���pR�v�������1Q�����W�c=�;^�;9�^��V�<�on[g5���E�"́L )�7P�����b��?gy��A��{���_m�m6���#귳ezrZ�ݔ�s7΁B;�sL�Nd������G�D���.\����ǧ�K:J�z$8��3��N�bs��pT������^�OC��n������ڏ�pKv5�1C��U��f �u7{2Sv+*�Vc,����.̃/���1q�Q}���=���y���V�s� j�ٶ��0��X����}�{a`�����;�b��+��	�vc�H9J{�p� wMi�؛w��|S���{��FL����ggzwj�
�E�lf��K�o�ԋ���lbnh��
�ӁZ����+�	�o1|S��F�f��ׇp�O{r����i��|�|>�{��{��~v���������Ҙ�g��)-i�t��w]n�n�nM�7.�%�^n�,%�ݱ�zKv��n��2��n6������q���hƺ�k��8��(����]O<U�`��rK��϶�&���g�ڃgi�v�Ik4
�í�Pt�l�:��pYϬݞ99�i�Z��6�P�˥��x���j�[r۩5�t^^n���V��!i��xx]c��WM����nϚ��;����qUkv�k�l��l���$�*ƕ��݇���y��z��tX�fϩw;#gSF�n��&�g\�S�Ȃ2� ���Ӯ�c����һoZ�;�v������ݖ�p�vN���\�n.�;�Z�틶�� �f��S���hvz����]v\r�/G5�uj�-���:��8��lq-�ᰜ��d�9��q��hݻg�u۶�i+�$���z�-T��n�m�]�1����l��p���oU�;m�k�^»Y�*�K\y#�m�F4g���RI��s�cZ�u�p���� �����.���x�BL���w[�������9�s���uUt郗��8#�;g#M���q��ڸz��η+��9�Yv�F3�9'�C����KzG��:ִÈ�{�+����9���V2<v�q'���f-5ׯO;��"m6,.��T];�t��%����8�kgZ�g꬧�V�=��p��Y6��wT�&�\gv����cb��mG�]���8�v�y"6�W�q�=s<�r����]L�e��������ˣ"�X�������H[��a�{���z����p��m�+�\�6�ez���9�M�n�f���k�P�=Y{$��/b�c�7���5=m�}��rTI�����`�gN�O�q�W�H%���p�5nm�u�Ҹ���z�U�59����P�v���a�mڝ�������/k8���8s[[pk��T^ն6ۺ+�=q��"H�\��Mpd-��U�6��xv�ǅ�mK㵴�92�5TA��hLg�<�����v���;����ܾγh�	��۰��=<�V�%���=�]:F���ݍ[��n�m���מ�zy�q�r�[�<�<�0"�:e�F6�癸]��vӊ�v���bc*��ļ�s�C�:-�� g�i;<<�����m��1m&l��Ku��z�$���b廑�/���-�m�˚�����m�:q�E��y�7O+����s���%�wWm�'��� �5U�Ί�%� ���#�gxr�85q�%�f6��qv�%������vɜ��ݷK��.!�<����腶���L$�<T��늆��`�n$�{��Q�ۋ�]��{on8�_ns���m ��y�b4����r�1-���n7a��u�F�v����U��*��ඩ�Ǎ�:��]F3۞B��k��R��7�T�����<�o�����{C\�x��p�{���[m���\Y�s��g�!�6��gF����\Q�۹��ɲ�q�'��=�7-l���e`�/.�v��9N�wcX�+���6X}3�Y�F�y�fu'.�g��}+ۮ�M'k��l;��v�<Zݸ�^�q�6����������-sv�-�-�	�;N�bg���=c�;q���՛��v�aܙ�Ħp՞�K��[1qu'�csn�<U�<�]���\�2;\� Y:^oJ����{��u���,ןk`�c�\��հ���y�	���l{qf^
%��v]����мY���t�m�G��u��f��:�:�������9;���1���%�N���FwN��=��c��0n뗟=	�Ԝ�n7.��^:�n�I����W 2@�7���r��֜���ZsQ��n㶹���	�ۮ ��ݏ��Q
�&��])C���/���M��V�u��+�c��V��5���q���������	��D]�	q(�쯎xSZ1�e�#gv�!����Lv��%�sPq{��l`�+$'�D��Z��t��룶�x�����o@b[�_lp�����[���]d��
ˎc����8�Ɲz��k�c�Y��d����㪜xR1�=��l�8�I��:�#xI�Unu8Q����#;[q�z�ҶM̝E�m��[�$��]���z�$3ۤf��v.��:ӥu��}���]�5]���q�VݺVN.��x^+�u����\�������ۦȩ���; ۞���mήzq��烷'n�W�]wۮ��(��t���O5�<�n�lBk���ӱ��XS!秪r�v��#�+���%���6�{c �1�N�V=/Yv6�]���Y��.:۳��,��d'q���<`�6��ĩ<5�����^�,��u�N}׶�k�Mq�t�5v��\�sĚkWo\yݯ���Us�s��g\@Z��o.|\��\�眩�Gl�.�+��]�=Z���s˲�w��]�8��.�ev��6�;:���ƍI�W[wIڅ�CS��#O�<c��M͸ݞ�cۮta��8̧kU�8���5�x�Qc���s�<�3�v��`v�[��p�<���7�5t��B���\��gH��Om�6�L�m����:��z�����\4���rD\=u�A�[t.^�S�3��N�oM�#b�M%�E�-�<�=K@�;���]ˌ��"v�"�w�[�������;�t���vw\F"��c'�BW^�q��l�{v�\���A��`�������ol�k;��̸��}n.�;]��z���5��8x⛷a�W��������N�ͳ��lγ�ظ�m�]��<��y۳B+�I"��;<��n��W=v�ҽonqq��R�'��lq+B��7<s.[	��n�y�Y����9w��-ϴ���ɲ�ն��nx�C��ႃ�6B�[��Ci�擷Yue�͹{��;%�vO:8=��ᮋO\�qq��قG\��
.�7b켚2=��n�ɳ����G5�ɑ�rj���n��1�;�ڤ�ƫ�/b5�m�9��7=�f�f�z�mu�m'l�.��mÛ\�:N}��T�H��nn�KU�/�ף���7uYx���6�8�O9v��Ym�E���w���i,�v�䵛vbͧ���.�Oi� 0��׬��ۚ޽���q��q6���^z_���]�ȩ�;۪�U���:����^����u��ۋ���n9m�]��%���*�p���=��m�F����+�9�cqjQ�Y�[����+�#�:.P���nO9���u��O\ܫ��5���L�ƍ��7ѝ���,�;�7c�%<��Ev4�Â�	�h��(���4f�F,N��h�"�枡,���mT�,5��Q�[�H� �#��caԎ��+�]>��#��s�6g��e��g���S�<r������u��c�7uƲ����m�Fv�GWS��qt�����pr� �x�	J�nx��s�A���]`�۷Y[�j��<��F�j#�[�x��{�����'/qo!�#�V�\��#�;�xW���^�Gq��8��k���r$t��=��*U���)ư%@�ubs�c��Ksl%vy9]�O�z���r;�����͚�����n�{{1ˆ���6��R������cڞ@,�n9�l�-m�t��W^l���l���ҫϣ�sʗ���u�C�x��7Q����zr��9^t*�Q�hC��ƚ䛰1��C��DQg�[l�9sY��l�	̡۠1�Ur�,xx�=��������o.):����m��ᖣ�v��Cu=g�MȊ��� ��JA`'! ��AL��`�ܲ��m�t�>)�kn9�vf��Fv�/YA<�y�j�t,�ˈ�X6�����M��v��{ ���BJc��M․��2�r�[��.K�tm�s�5�9�B���o��4⭞��c�u�/��;;�t<OS�;�{fB�j�e��t���ݹ1���m��'V�mtm�n�=�"�a\�h*e�P� t*��Gg8HG�͖Tw�s�ps��湇�n�}(@s�v��*s��������xI��{e����QɤA�i����p�����簮�ۮҹy��0\��l<x���<��ݪ�P�k\�=vz�>������2Cݸ��%�맶4�1ώ�ݛ��-�<���mQZ�����k�>P1�z.��u�n����^]�]ѝ�u���q��/n+��x��j�A==���Lxoa^y����Ւ��t�9@��u��&���nՎ:�Ok��H������'C�q��ɂx'��W:Z�g����. @]����p-]sͷkq����+�i�cp�ln��N5��E��6M�<m\��tsӸ�{9�N�'3��d]Ygn�t
�ɺ^ufh�d4��ov��<p����ܵ�4�ٵ��֣v9���nw/�hu=ö�<�7.�m��5���nm���u|<rQ�]s��	�s���}��am�-�1�\�т�\3����Ѻ,�nN�[.7:we�b�{�wFϋm<9�7��˨5�n����gfw)�l�=��S�=G&��Ÿ�Wo['�.{rvn}���3�S��ưw`�=4�+��4/0�I���h�����k�^�sb�:��ڣ�����Om�!-�u�\�.��l���q��Z�\�{�]��x�g���h�����i+l�_n^�;ͬ�c=�)pns����b���+�z9�SU���{�Ob磰A�t9k���S�8��v�Qkl��X^׎�[k�=$n�L\�目ܺ渻px��%�j�U�� �����Cm�npp
��G��D�ض�d4�ؼb���ѽ�8lsɍ���W>`����r��X�`t=CB^�]p����n3�f�Ws��i+j��f5\5άOM4�5g8���f�X�=7j'����Iu�a�FZ����pje�9nS0\��vF�_��F4Rm0��͎[�n��ͮ_<<���I��9\+��r���U��n����9wtQ�n����wy����u�s�r�r�r��ȷ2cc�,k��".wqs1]�k���wu��=���,cr�1����ƞwv�77Ms�����ѹ\�#�]�����4�r��NWH��\�p�ҋ���������t�+��̻w\㎹c��n>���$\ō���ܺ�K����wWt�w]��Dr�z^�ˡ���:�msE\��N�^�:�J��E�tr㻛���u�N��Hl:	˞o+��nH��&* .f()�I7��/3�7Oi����n�5X!�맱����b��q�nzе��f7'+m쮬�D�#��v9Ŏ���6�-��h�8�8�c���ըzy!{q��r�N�ڱ��s�/��]/5�y�Pr�᱆�n��^�-r)�������Sg`c�U�ؚ��]��M����x��6i+v��n���e�5�������v�Wk�8���\�[��"�2s���p��>8��nݺ�B��uթ�m\g�[��J����B���ԭ3&�zr�q�u��.,qڰ�u�l����!
D�YR+n�/XwY�g;�������p��gt\س��sS���U�0�ƽj-��pe��� ��:��-��ey9ۍ�9`s��3\{N�pE���vn��6�L�����h��D5d�X��*�R��T�I7m�g�wH������<��q���!�'m�=��h�f�v8�ͻys���m���HQp��������wk�=n�v퍥3O����+��<����g�u�+솳�Ǝ[�'^t,jwn=s��W���oܘ�t����[	c�R8��^��9ބ���g���m�s���J�ۖw &��h�3��Ǜ��n5�L��Cv뷳�g�;��trs��q�mf�����9�1g2#��ڴ{�D�l�]��&�����ü�q�i/l���L|'�;|qt��<�gun�<�[��ԸA�	�6��@^{bxn ஢��|%ϳuݽq�z���{;Jk�����N��OV(���<.`�P�X9{c'/��Ǎ۵�t�(́qS���Xm�gk��<��뽴oU��=4���/'���[)z|5��yt�����k��@�����@ǰ� ��E�:,3�F,�v��ֈӵ��~82nքݪN2:�ݶT���!�֬�N�G�O�"��1�614�BU�f6��*���b:����uvL��6��f�b�3��d�3�=�{�|���9�N��N���c)�ô�t����zs��{��S+L2�%�d�
\�չp����'��xvvP�w;n7#�v�v���2+�;l�'ayre��n�1ݽ�Ey�8�@�Ϗ��� `�nF���0���k�9L�cnf�r\y#�g��v7c��8|m�/;�G��r(v�'g�092�ٕ+cq�p���\�����|ia8�	���G~�D�-�� �I+=41�ߺƥtsw*NH ������Ͱ������^��Dߡ���ᵖ�f�d���(�?�}A}�β
��h���||��H��TAE�t���W��Hʞ[�:�+�A�l�H$�}At���-�՜�]��֡�W��G��Q ��g$&��ݚ��=W��O���Q&��QDRp��z������5xu��I��(�H+�}_ K޽�K�6\��u�B1�X�)ӱ�G�Hg�F�su�6�pr��1�1<h�&	S��\a��B(p��� ���h"	���팋%����~$����>ߐ��XM�e��V>=U�;t��P�xq
s��bq8��Y���}�wB{k1��ˬ�z�߆�={gEl�r�E��ή5W<�&��g�����x����+���Ē��n�u�}�vɸz�	:��B��
��3e� ���A �����K9��,U�� �^�������<�H%A$����z�k��H%�/,_��}�n�;[<�S\H6��	f�ى�ڂ:{U��$/5�$R��Z�iQ�� �~��$�������{8.�,6;@����<��:@v��[�vZ�m۲Lk]�:"L7	Rni�.����Q� �J_z���H'�Oy��:�m>W���_	!��]��j�0dE�w|����p;����O^�1���,�_e��?�g1@�0�l��]�k�' F9�|����n����|w��ĂA̞B���֓˥�*��7w�i�E����]����lY��r>�zף��?_��z5��f�ӷ��[��}ʟWo�oM�����jb��^�������V�:'����!6C�Fn˛�g껔v���?I�X'Ou0�E�tE�Ɏ���%��$b��2�R	PI|��:f�J93�^��5g��x3�Yw��]��A��(jGr��g��,L����y�x�K��|t�Bt��NٴkV}gg��Z�	'v��mD�e���}�sj}_���
��o��Nmw�vo��	vԢMi�j(�d��Q: �ʔI}^�����bˬ�$fuJ$�n��Iս��[}�:��Ԝ���1������wg_�(�I�oJ��}��z���H=�R�"��Q?u������n(��ޏu����w���PN�\��}��ٱ`~�E��[��թ���/U'��ޡ��PЖ�t�_ٙ�Ϗ��5v��N�rS>��<�>�zp�� �uJv�Y�%=�>ɛS.K��e�o:�#V�d���ut����e߫^�C}t=�W�A?钁���˰�Q�&�]t��k�9+��ڝi�h�;��y��m��68s���w��pnQ���~��,��mH�U�8�Gd�(�����`�AR���{x͛( �͕� l��bm��A�"���u���Vz�c��ʀxnN�D�F�{.�$��x���*��Zyr�)H�N�?T�~�����_�}��e�S_��| '/'��	�mw���j"eC1��uܐ"�1%�5��~'�=�m��:mAӯ"�jN�ܢ9���� K��P5�6ŒA��V���u��6�TN�m�$wN���܌�Ȟ�����j�g�e�{��WZ���K���gG( ������9��s�	��}��Y��{<��J��q�ک��8��6�R[�+`˶�r�՛�V�Ѹ�p��y}.F^;���k�P��6�.����h�\��m���{bi6���&q��,�����+�gEu<nY[o\�tnƍ���%kq[u��e4��&�$����؞�Q�y.�d;g�Kj�Y]�g���_f����uw/[[��nڻ�e\8ö�����eŶ`���RJ�� C���8^��\=-O8�KzG��u����_Oxm6��\���	"^�(Y �N�
����&�wn��3%L��U�u_�),%n�!lZN{~�m>s5���Xm{f	��=��	;ӥ\�++������a,��J2�pEvo��X$v͂��u7+`��V^����X�A�(��i=�9e��Q:;�R���n�0�R��G�t�I�����^�;��D�o��:�!�jn/��ǉ>�@�����S�{Ҳ�O�Nu�}Ҏ^\���˶"�p��Gu&�vKSqefۜ���jޝ�"'�j:�gv�K=�_y�#�(H�7�i�u_ă�ӝ|H$���P������M�wN_���$��t�D�l��h��Fһ���(��={Á/��UE�⧍�s~n�ҭ�����t��v�B��M��U䗅l�֌c4�*��|��J�d�7/N�nm����n՝u���n���H�MtA6��	�٫I��=��{�}[��	�e��1Ƙ�Fۍ�w��N��@� �����l�3�;��;��~'�f��O����~ڴW�D�Q��]�s�w�ݳ;�j���p��75� �̡D����b�yx���Q�'��#��X�'@瘟|A*��w�'�Ht�{������'�o6P �����[�}�읷U�h��dOᧄ1�X�Ξ�[��NW�קu���m���ݫu�IpI�E&nb"B`i��v'�tA�zQ$����f�I�"�f3d�yξ �o:Q!���E�$vnY�n�g^��oA �F��H/{�V	7ݕ���q�7�~*8ɲbm�ciU�3e	���,�I�8q��n��kἦE�]I�������R�=�7���k>��%��%�۪�V�>&��ND2�B��屋'w}#�?~�@�!�{.ɮg�c��m��{�a�{���/5�A��<���	�NalS}.��Y��5z�2���Fp%c6�a�]R�����a'�1P$W{�b��ӝ|z�{ػ+�G����c�"d�Q$���ocF����u��Z���:5��V_ϯ�??�"���U|�Ă�=���Oںs���k��/'�>){��J�{lX�5Y���4�R��:�����}�X�w��'�B��X�	�s�ǵ�^��ʑ^y�
���i��D7�
�ͱd��Ә��{��1V{��R��{��=9�Ĩl��A�$�Ұ�����F����� �k2��yl�@�H���g}�X�ݗg�õb�ؼ�RC�:�n�SAuU_Bg���b�����)eOb�z�5�^\R��'�x��O,q.�vŋ�>�i�$m�ؠ�{�~Z�W�ޯi=%d�$VL��ă��:�mv�r���wn�
�P�$��U��n���������G<�m��3v�=2����$}�'��
 ��,���݋ �;5�$A6�j���G�̉@�ٵ������k�.H�,&#��;�UA�y	
f]�U��$j�΁$�m��(_f߻��{;�`��U��hAN/M��A�v�$�F�d���z�߭y׼H$b�Ή��m��927��CpI��z���¶���+]A ����+�O>��ݰ��Jt
g�H#�UfE�L�?{)�x��j��[~P>k��`�5��즶��ݩw����W�ڼ���C�A�v�pg��jH7n����<��������O��"��!�F�ܫk]SS�ɦ���u��u���(-;�#���g���:�vݻm'��d�l9�xw8��fZ�#�pi-Ĉ��vlɭ�-p���]Lt��m����Vkmzw]�����A����V�[��D�Ds�c�d��q�_���[��b�R8�3ps��9�Ύ�F9���v��u�*���3��GiPlY�@���۹��w
�b��7�ʹ�8�������,/1�4�.�y�q ���yn~;��+ۏ��\5������_߳z'
b�N?5{��$k^�D�u�����{<V�[���Ô�t~�ʧ�&p��	]�ٗv,�5�<hv��*�� �M������ڲ@!H�^��S����j��$R4S����U|���m���H�w�h���y�'��{(0~:��V	�\�b(Z��ӁK�^�����V���Oj�W��H8��VI<�s.�<���ܱ>>��A��y���pH��I��>�_Y�FgP���ϻ�ꯉ����O>�@�_��i�'�ׄF䖦�Q����P��D�ی��oJm�<�G�����l|�k-9/����?��H�J�����~s���A��(�����p��[O�o��`��|�8TFp�@}�P��9ٷ�MK��^>9N��+��-�P�����l�ͼ���߷�}��'/C&���Z��ߋLyJ�j���~$�o��d�5�J����UwU=�Uq�8X�0Å�J�컫��vQ ��UvQ�U��w�q �g��A��(��h=�I�$đ:}D+��'�W���=�d��:Q$��}��Ъs3n��x��Yc�Jf$ф�ۀ��u��|A�����=O�P�ۿ���>�m���*<��7z*�|�m9*�-�0�����Պ��7tPvu�[^�N.��٫kS���2#s��n	8y�$��(�A"�N5�F��6׫�o��z���΂�.��,E!V@�N�Oho��ެWh�O������+�I����Qy��o�"Y���r� V���B������/�Ҁ �~{AN|,L���y\�k�J���U�����zf3�fq�
z��k����mj˛��I��x��kc��i��d��@D�r�v���<�h	�	# �w�������k�n��,;`�+�wY��-w��׬[�)�����{�C�pT�:�+3��.�}=�4��J�T�5<2>������`�:4\��ٺH��j𶴊��C��+��^R��r(h=������$���#�a���@���ɽ���F�;T����q�������9�fz�[D��8���<��h�Gp��W+8S����.7�y-�c�%�,o�!t�Ӽ=���S�b:�^y訔�Ax�n��8��6g>n!����|7���m"'_˭�}Jӝ���8�I�Σ�H���.uo��t�V�[�p����	�|fLo�z0Y�h�$�?�Z���6�ºy\9�R��2���ZQ���f��ů"�yN�$o�J_jJ�o��Y�Ɔ�5�q(�N^�����݉��C���N�,vK�p����=�i<���r�x�PaΤ����
�Y-n�ݔ�Э��hzgpޣ�Q�O��X[8s.��'� ��v��{�5���}�}��nR(��OM1L��疷�f�s����+%���@0���w�ǘ~����)*��K'�]�+UݹR9������{�w���g�0m|wBD����.��v���Α��3��Y���9,/b5�CO0j���A���m��J�.�ZCܮ!�h�����X�������H��$9���wg�Ӹ����W$�snqݳwm�s�yh���!��E��׮W.Z�r���ܣI��.��'wG;}��n&_w4�7��=�͓�n;�����a�Ɲܒ�p�h�hǝ��0b�.!;�.�D������.��͂�������4\M����˒�b2�"�̀�7M�WL���țݺP�q��rD���wrF�6R,_5͋�z).��c��I%LH��8����vM˱�]݅��\� ��0`�i�(#<�9��zl�I6��)�O�D���˳��qm���웳�$y��D�V���;6��:�_�9y����T�H�L9������a���d�����G߶���>|E|O˻�c=��ˋ:���
JBrM�θ��粑��6�u���W��� ��<O��<J���j$ф�ۀ����'��D�H]�˳�Q�/o�]x@}�R��z����l!�>/�����ٶ,��k��z`��,��6�q��'���$���2��K|�;ɫz�.�X�!V��v��@���ʲA�%�j����M�{K����]�~����bh��}�-����W�d��}A���m�?{�I�C^��J�����c�r��bhf���i�퇳s���r�s;�EN�ٺ4أr÷u�1�!{�p�W�w����U)+N�$��.�魫G�D�V�Q�=�ٙ�����~[[��6��b k���Ă~]�ۿ�$���p��JLX�֠�	�V�X��	�*�!	�M�;R�r=�y������l���������#S�\�|�:�A }�$��@�̳[Sxq��V��Vo��9��q&�&�]���(.��oմk����Q��IY�˿�$�N�	'���+���ws��qϽ)����$�Os��{�J�~<���k/}�D_"�۴{�o��Aޝ(�����Q����.s��Jc�zl�Y&��.�$����@��6��W��D׮��[�]Y>��2���[�
�Q ��������;	�g_���d��7l_��wgJ��I��(ܯn�^S�pQ�s�ґ˥ֵؾz����oS�7A��J��.��n&ׇf_pk���]���[���{�3XU:�x���({��g�<�t�[�ͩ���btn��ZbTU�1֒�S;�l3[8���it��'
.n�N̚���G�n����y֡�[ں�hp[�c�vnz�N{o͸�Ry�<���]q�ƫ�n�:�x�ٶ�X<g=��{s�"=�q�춬ݘ�լz.��9�9^7
ucҼ����`��]=�W&<��O[��q�榋�y��8%�V�׍��m����.�1�6An�m���u)�+�,�F�'F-���>��s�\��b�U"�m��o���j���U���wW�$n͔$�ޯ��t��f��}�H#�6P$Zi��#	@�.�;�R� ��&��<���� �Fd�_I��(��wv���R���#��IB`m�e��'���(�2��+7�KF��e��$�yҾ$��D��϶4��PI@����]+	u�������	#�z�	}��}Y����k �J�)=8ŸTm2D���\킁%�����'Z]��w�@�U ��a/��vs�Q��;�{�	�D��EX7���k&�0�"�����9��$h�b�p�#��v��c)HZe�g�o'A �ܔH������Ǖ�̓u}(�q��j���`�F�컱a��>�ޮ��U�{�}���+Bڪ��ǲ��/M3���O,ݲc{���T��x-���Iz���$5��6Kpb�x2�N��A��������_�]�;]޺�4��c.H�Q
�'�%_{�� �KN�fRѼ/�<��D�I�(�Ww���W",(L	��=r���f��go�����~$��ʰI��K�{�.�]���U�%�ϖ��	�PIF���]�n{�}���uR�8�A_	[�u�'�y�J.�-7y^��Y�x����McX��^�룍q�s덺�t�gX���n*��ìs�F�HZ�.fJ���+}쿅�'�t���B�(ve���W�	+��vO��Fd��!i��+�I�v_;A?e�t�M$�Vw���~$}҉%va��g�t�G�4]ߚ�&h�<�����N"�~����i���I_��2�<���>�Q��&��At��_�.p�_T�к�6��=�����:�`ׂ�׍������qJ�]��P�t�������`�O>�DV�� m�ѥ ��I`�����~�߀]��?y�A@�}�w��zw�$e{nŌw�؁�	�7�:�����E��[�ݫ��'���X�N��_�?}�!����l�^�}�Th�����,�,;g�òu������ݥ���i ���߻ߎ�:Q_��N�o_�Oޝ�Q$����m#/2�g����	'�](�0��p��WfN�D�<ܹ�[�{]��{2��{+�	_t�ū��j�u�T�^w���2\�&[�
��Δ ����A�����T��O��](�H*��6��dA("7gݕ~�Qz>�Y�Ѡ�3�J'�J�t%wg�`���1�,�\���M��V����m�>sO�c���2]ȷ�w ��\�N�/j�jg^�f��K�w,��1����A[�+�N�;�ڍ5	��}$�$+���Y�V��
�\�OĀWn� �	[��{_�b���8��L;����O�܄X������N�bw��p�:8R_���
n�yԜ$���+�I+{2��'�������J�q����ZʉF'�A%]7o�d��o��z�h'�~&��}D�����,��v�Ss~��{z�~S�;.�!�!j�y�> �U�eX$��nUO*��l�O�d�� ��ʲGxؙ a�Ji�`��:V^w�WӴM$NlA^�˲I��u�*�_��9w���^���������}� x�k�z�6��=��{�fWP�B�ܫ�O.�t���:y�#�[菞�Ѧ�����^���8�w����ֆ���{�`'vI�7{7���5���ѹ�
���]�Xvg����\�w?�qû�C�|ݫ�ݷA��n����a���r�.����#����h��p�,�]�]>��/����2-�n{\��;F�&�ћ/\9��]�7��u�s�^$v��%�����'Z��Q��Q,�y�c�'%6�K�ɧ�v��70�����oA��ź^�]��s�5�]m�a�N�T���cv��h��l���쪼&Q9�팼f���[u�A;`�;v|8�u��@]Tv�8Dэ��UZ6���~�
���;�|޵t������$��us�{yvP{l!��f�eI
��v	��w	�@`-��)t�Q��Tv*��M���+ٹV	$r��D{��\�%�Pg���eDcS栒����d�|z����e��-`ބ���B�ܫ$��tHS�Q��15w�s�T��g�9���^���G-�P6��\���!�L$)�w3���@�eC�9�$u�eX���u�ā���O�W1_��+��gw�jq�ٕ���W_6�BI d�ЧM��r��X��I����z9�倎yK���~��u�D�#�{�Wb�$�k]|H'�o�P���<'Z���p������	��Ή;g=(���;�۽_��A�l\��&��y�=l���:{�d�4�_K�{,�N��e���_�?a��'R���1b#�T�G�-sC�E�;1���GD��� 3zwW��]\�M��(����� �*cɩ8{�Ak���`�\�+�R����:P��5���q�	|��9(h$b��D�A��M�%���jT�ƺn�I��A��׫�$5��I�vΡD�~[ٗ����&��]v�~>�-FC�D��g�U�e�d�ߚ]�V	���� �s�J �B�̻&�nkqW|�����,L6�,���mۊM퓌S�;7��o���[���[��f�ѽ l�l�`���	;鲁 H]ٖ)_�����*����	��Ӡ���ͼ%AHb6=}+>�+Ω�7�];�o�7��	'�e
���.�3*zofr�����Ȓe����|zz�@$���k���c���6�c�`!~��r���M: C�χ��6��v�}�</�(�YDd�r�z~�l����<����-���%fe�>��x5� ��o��O��wg�@($�~�6N�Si$���N��Ν:�e�}���	<��K��"_t�V�==;<�;��6�@"�2���C�ʋ-q�Y����u�@ ���w�-���f�'��{VI���L5`$�I|���MKy�[]v��[y"} ����&6�]�۹���F����5𘴤�X�w�W}�p��Z�'|yۘ���İl��|sk�7;���s�˙�3�ma�%���-�($	�T2ͨ����-5��ݐ�V��*WN�I �+`vzviA�]qQw���x{l�n�\̲E�[
�G��ۺ|���vvi@�x�F����g_P9�m� 	���P�t��V����3�W�#
��7[����$��H ���h >=�z�"櫸��f�����<P�}�d�wN�����N	��{�Awg�C=��;t)�r0\ó#�uo8�?zN�=�᣽g����Ay��O�| �Q$���Xl���~��	�r���N�4�H%�+���A�����u�| �����g�{z���N����^8��P�`�A6 ��RD�z��z��m�<�v�u�'ku�*��k)o����%Rڬ
��$e�������@������
�+�����D��$�z���9g*�P8�Ѵ���- �↛Ow�2⸰���tZ%$���j�I$�t�	|��WR3y�E�p7�x�oxS������n��o��V�6�	s���[�f��ɵ<oBD�����@#=�\o��5�[
Ј�8$�{����^���~'��k�RH^WU�	$�{Ն�\��`���t�M�@{Óւ�+�3�ue˴JI�L7j�z���ȝ�_�t4� ��˘�	�k�07�O]���lf��~<�_1�H�9��8(��Xa�|�u���/xo�������.y��(��Q��as<ݣx��:��389�nm8�ai�%V�8��4$�`$͞��0�e"�w*�;��v�T����5'������[L��-yo�ڸ��Z/yy���m��2���#1#��;������h�Y�F�aK��tԧ��zz�{�=��)������L[<�.b�q�.����&�w7�E~w� 7�ڵ�X�sӰ���a�.U���[�_���%lG���>w�^�w�h:�>�G���"�°���pT�u� ��4ȧ��O˟4)��9$
u�W}E��Q��[ǯǂ�Y����'M����{���<�]��-~{�j��H�d�����]��)1��I{��e]��v�q�Wz�[!��S�<��`�c�sۗƮԻ���>X���0�W:��ޒP8�������]�+Ec�����6�����4���N&{V޻��m���p�o�����݂��{�=&��>Z/b��n�h�5}���Y�P��f��}3�M�kޗ�F�q�h���L/z�7ݼ]ع��co�<�/3XܧS*�H��y���=N�z3o�����tϽ/K�O7!koI];��u��C�0׶�F���Z�k��6�n�O jS	��z*3�;ذg
F��IA����h>6�:��o�bn���,��b���n/J&�\ͤ&���{_2s����Sɮ��̓o��ce�3{������Dx�,E�n��b]��c��\�����oӯwD�n���g�F$��%����s��)wgv�gv��AG�xzM�r���̋���	%��ˣ19pwO8��]�ɉݸfB;�D���;��w��DwK�].p�;�w]���]��Jd^��P7;3$B���"@`\�9rfwn2)4���AD^\�"��
$����iFDb),
Q��)�@�tC0�F$��i�#�O���fƈ�F�N���{�6HJs�(�n�&I"/ϟ�����}��ڵ��X��vm��0��s��u�g����g��y`XuvSO�k���7����`{.��g\��l��q�@�޼�P��!�&)�8�ut9y�Ӻ{$Y��a۰���n��J]�;�'k,��:���0��W]l�\q�s��k�`�ܮ<�=s��rʗn��7��y�۱��n���\�aÓ�4��t����CՋ-��jx�cg!�s�y֛�\-��ۍ�����u�q6�G\Ruω�dȡ�m���ǋ���`�u��qoI�������UT�;[�2S�������U��.���롇0F7�:���V��
�mۖm�v��\�.vy�h���٬xܻ��z+��G��<�{9�!v����9)�H0�qض�2p1���[��U�!Ǻ\�mE�8��z3�q��F�;W;��l��]6�Ƿc���S�'=�l�s[��s�
���m�P���s��I�ܐ�7 �؀덕z�!�%���/��[c�7��U�N���v���ԍ��q��[^�9=1������۶�`M��ގl���3�nx�3۝j��@�ybɲ󻱭��Z��ػ�Rwl�qx�݇v�y�)Ѽ��ɣ�8���S�[d�s�:)���G��;!α8���N��G���ry�Lx��\��)θV��5̹7�	�k�'���@t�)tlk�Nۆc�u�.�=c���I�����a�c6�x����1���[f.�)��gG���t����'$
V����rᨱ'�:�����۰tOj㮓\<,�qr��&y��m��4"[��.�fsv��W�3�ٮۚ�Ɍ�K��[.Qޘ�t&yKkF��ݺ�Ü�3x��ڻ��v't��N��P�/NV펎}m�1�]�u��t�F�ۘsE
ܮ`N�������e������}���n�����\�Ơ7	-�lݺHn�b���i&���&��~�w����:���]��$�T���gsp��Ǳq��uۍ�nc�m����g&�t�q2�nq���ݛ���{tq8�=�����ݭs��;$Xz����z���Z��S�u����X饵n=�u����6.���<ݳͻl{�^�|m�T탍�p��1�7W!�]sr<u�����h[��q��l!fێ�Tyy}��y�&[��d��Of�n�:1����<�j=f:MqCt�6z{]Q���cr�2�uw�������s�njjj 7�v���}x��b�wpfnuy߼���:h�	 �ke�WUu�҂;5�i�I!��:�ٚ��> lY�sX� �S��b DWL���ٶ��?=���끆�+�����v��  �����v+���3�jf��;�r�n{׏X�q��(1�T2���Gɟc��Gz�Y���]|@ ���,��)�k��tz��o|H����[�ԏ
����B����{��� �'M(]���x:�].m��$�{��ɰ��=T�G�s{��s��-�bm2��]��ي��Z�Xz� "�U��U6�n��[-�:zv֊!�����fg�o׏0'y�J�W�
��2�%]���%<�������1�DENUk���f����;���2e�ޗj�܇�ߧ������\:k����nz�}�1U�q`\j���tW]�/.�à���͌i
L��Xw�Zվڛ]�u/OT���}�[�ߖ@ '�k�1 l���΃m���>z����꣍��PGf��8- ��/s|��W�N�����;�uH@N�\y���	K�yTDU[a4������^<�1�I���F���������",�O�Xۮ醬$��z5��&2��Y�:>T�$+���H�]��~�_n�$�f �F�g�(1�޸��=��d��V��,]�<WC�흄�"�)��D�:J�g�]��*U�J']�\�S]E*K`m��J4y"w[�A�I+��f���#�����d�I/tz�������xBѦl��t�d'	��m���~Lz� ���i 2��0�.,����o}ه�%�y]�PL(�B�������z� 4�Wl��1�߶s�'$��c��Y��y�w�۞�
P�-����Lj{�����Gh=�&�N��޽ξ�v������O� @�^x��g���qv�_޹�}t��Uac*�a����ռY��g��iysƍ�K�eY��I|����p�ޜd��ؽGS�)��E ���ez�����A�>W��Wo���J?O5C�I �+e�l�ެ7a,����e������D�[�)���u��T�.ݻs���W0��v�^d�(�t��x�h�u@+�~,���� A��06N�\y�*�^'�ƍ{%?:Nz�U���^2�R4��^�6��B��&뛶�׿@� ��.� l�{���@ ��0�õ~���b��"1�c-[��/.,�	�^<�`���w7��������@�}�@��������cA12��:c�ߧm�x�����`$�)��0�H�������ʬ޵���r�ϳ�=��l��r���^��hn���(��XU]���5[��9�&���q��[�/�J/�[��wƎ�6<��}	!	q������qy�~�(�NUK ULϑ���� ?OJsͬ���m�W�)�%�^�6�I�Xn�I%��ϝ���`�1g����ʝ��^`��g��;�Gױ�sc�]:��Y�� UKy���B�Z�vI���'�0شJ�$9��Y�!;�X��C��␐I9�τf~�sy[�u@+�����#�ަ2Nj�`|A=�Ǭ|��M}F$>,Dj����a'.pp,
In�!��v�K�-�B$'+����J�L^�g�H����D��5�٠kV>����1y�v��"|��ظ�� A��������H ����3M>��X�~�a'-n	0�tx��;��$Q;����Q �/ut���W�9�<�4��q�$ �9٥F g�됕�/��v[[����]k���}�r{C�o-�6���M���C/{9�ݶ��l����������o�	����/�ηN��ٻ��I$��f{�3vz�=�gdG�'�ͳ����Sr�q
��b�4t+$s��@�m��,u��������dŦ�{BS�=Tq������ܥ�3f��){{����L�������q�"��m$q���8�`�r�q�-9�<��[�5��Z�\�t����[pH��/bn������sɑ"9�#�N���m��)����甤�\�M��l�/#m�s��wg��#ُR�����}������U�G*���޵� �ޚ� }�c���Ǩd��\ Iy���|��&���a��%��D���/��Yw8شJ	!���A$���*�D�����>Ύ�@{���+ ���y�,=鯕�A۾�6l�ě�S&߻��bD�K�Ј���\�$����(�`RHڲ}}(�<6��~�7@����A˾]<H��6H����Tmw� ��󨑯#����s�c��eŀ	�^<�M��pY@�Icu��I�M�W�E$�{Ն�|��ga�7�y��]�����;s՛�[[�n���[�s�I���IDu<�j�n��w�b��vғ^G!�H�%�KӺ_֒H$�����6�ܑ��d������4�W3e�HMڰ���m�vk�Ӗ�K�z�J�Cj��<�w���^���5zv^#d�}���?!���B�������E�C���6B��릫e�J��-D������� }�׸�t�C���u� ��k�0H%WWS�_-4NtV"@;�/ĦT���d�ܾ�� &�x����Zn���*�����^��v�I ��`{s�+�*8+�\�����G���> .��`d�ǘ�@�\_r��j�U�PW���/~]N�-�4��O�` ���H�a���͠>���� ���<�l=s��zj���y��}"d�L��$E�س�q��nTݎ�뇥:M�]N
ȤU�Q�A���}�}b��ϝ�9<�w��0 	�^=<I ������V{eo���K$�9�q� >�}5�1[`崄�=i�$�y{6�<�Q�G]���$�A�V���$���ɠ��E��5�yg��JoKˁ��pGW����M�$�]͚�"e%v���{!�2Y�n����$,��;����&�_��j��$F�V;�{8�r��4�v��xK;O>^��kQ�����>Ͼ̲t���D���7i��sf����ː��1�v��,kx���6=[A$���7h�W�o��	/�7;�{��Іe����ko1 ����2*�e��p=�D�ٹ(��x��<���BHU�Y�� �w�_*6�^��>�;��Rmo.mzw�wZ����M��l�s��Vyz|�ff�ģ	�)�.�U�x x;٥C�/}�x�]r3�����@��v�I.kyЉGWkbBU>v0Ɂ�̸�%斏8��]<� ���I��@#9�\� �b��;l.�BmnԐ�NVP�i�:vO���� _?�d$�O�����:O�K���M$����M���08҂D�p+����nTPfh�ž�~H��P�N~�O�_8! z~\{���U�Xs�ϯg��i���+;W�x7_,�$�m��ϴ�,ogk���3r��M^�F������z��=���HH7��0η�3f������n��#mݥ:�Q�����h�~�I�]�w�Ma4�@޽s>��Ǭ	.����}��Y�񋞊L"�D�i�u����on��R���><������V3uB�__|�����Yb��\�*�uˋ������68��P�3�BI��R�׆"R���F�W�Vn�	*��7�f�iwH��{g� l��ǈ��_	>$���$2[{}����:=��{�VIT���& ��\�����<�"[�1�8w���I$�ϔ��I���ij'k
bNH�uaquJw����=n�7�I'���!'�W�L$�������K[{p��%+n]����`vV�%Fa�޺���O=S�a�/�wy��R{%I$��Xl�N�|v+DR~����3��ǼG=���w���6--]�Z���	��G4M;f��sťW����8Z�8r�Џ��n����=߾���̥����ϦuC�{�v�^�%�j�8a�����od}=��6��Y��M7m0Gk����q�O�;���0�m�g¯kgz-�wW��l�4���&��N���;�ov�ѱ�<�s�m��7m�ۘ7f�������
���s����l�u�}�l��O'bϦ�6�y�tݤ.ꃓn{kM�`��!��D8Nl��;nyp��W��gi�1[�Z��^ϫ��'��E�OHx�B�DD(����H�MGd�^���?6FZ�vI��^�., {��y�?O9������]#��.b ��q�y��mH�"��Y^WӍD��پ�wM��g֐I|����d�H-=8�E|�����,�T̥�7�$�S��JL��8��[�Vh�a.:��A%�A��7���ɶ�g��m$_��7a"O|j!Gsb6�$T��e˭�]�I=�4�Ii祓_$��t��-�m�5�I_ei�Iso�ڌ�Z�m!3�]=P@ �5��m ��	��%��\l�I��j"�H߫�_�S]����M@d��ls��)�P���u�X���N^M�J�':�����%�����%��d����>�H}�z��H�׵���.OT���?	0�I<?/��ho tX��F�XJe��i%1d����m�;s29���6c���I��I#_�G��|�Oy��:j�ά�����7����y#���]�v:4jb��Pe�|>����ng7v�, �������oA���j���jn����a�-�$*8mXP���4[�����H�V;��Ml������%��ӍDPI~��$��O�H�!��j�j�du�J�[�������B$I.�ʳi$��0�jl�9e���DI��č��0[ ӵF�9���A�n��UޮL{Fu3�l$�\���>��W�E$��Xn�W��sk޷ΛG�J�/�h:Qu��j���[g��k���1�ԯni-x0.'����}wT"�j2�^5(Љ����7�D���Xn�I!F�O2���&tMu��׮g�;��d� �VJ�����F�K|M,pg��F�J�W������~�����j�!��G�$�Q����%�&�m݄�_K�D��0ݤIO�d���ێ:�Y[��R�<^�h�;�� ���.\+7�9�Ww���������>�JI��3S+�c&܍�xّy�Zq����WN֑7�j�t��{ۯE��
��E )k�N���y�|���1inp��>�0����gݕ�oN��{c�}\�K�;p�k3�t{OW�r{OT0{n�=��*�{}���O�i�'���E�x+�u���s5Q��5�~~�(lH!T�R��Hoyfk÷�do�?������{d�b_�hKҔs8GI��NX����B=�^<�j�)e��d��Bת­ɋk~��Õ�f�{�n��hOF&Y�'b��3TiL�@]J�w��x)+��mVyR0�n�y�6ˬ�y���3��9W��d���ON=��Jv�zI�宻�|!�
�ga����|O���n�}��2g���z%����g�|��X'"8�ӧt5�Ρw7E�/n��7q��طAa��������ё�!y�
%{�8[w��,�o{f)�����I�u�oby����k�İ�irn�v�>�;�z�~\�d��)f��L�-�lQ˓2;�ct���c}1=���C� &��;��jé�8T@e�+�������t��w�]Q��.���h��Κ���y]��M�~���iR���X.m�w��:{�|j��S^]_Y��j�Fེ�j���h�s\@���3���yY�N��A�Q�|$9^��W����c������vߪ���I�{��Pn���� � Hl����7��j$��2-"��wQ�X��A�4/u�>��ɢRBR|�ibfM�)d���4�LY���&6̦9v��nQE�ęH��э(�J�ܥ&%��H�6A�h2����"Ѐi�����Y&�d��q{�P�R`G����$;���@2!�f�]ܡ&�)FL�B	���"{����l2�6#%K2���b�IǺ����"d�1")E��ۥ0Q ���j"�L������e��"0y���%b�H`�&} BI��s�}��1̧�a�J��Ն�$����cq
���<흐�oF�&IԀA�vo2%uma�H�����M����<�^��]��ɿ5���ݖc�9�c���OM|��I�|�D��ڿ�A-���� {��҄�o��͕��46�ƶ/b��-(�d�S]Xȵ��:딷����	�f_0�� �"h� k%�v-���Ɇ� �+���@$ss<6o=ꙺ��װԧ�`4W�.��7i!���,���9�����(_wLw!�ͬ� ����� w��҃��o2��R�G�=�dۑ���7��sN, {����>l�v)�{s�|��h� w\�b@$�'���̮u�p(��V�����x��q����Ɖ$��U������V��~]K�������|9L�*�Oiw�����ot&��=��[X؈o��Y�����S޾���\�IQ�k�Ut���o� 	�ٙ<������9�)OKhZ�+��E�Ǥ v�sE��ooz��o	}�Xn�@$}���_$��}w���up�k���C�c�Ԫ�V rV�Zzs�)h�u�A֗kRuK�����i�+��>�{(�E�m��7�c�� s��҃m�\�։�/9���0�	�U����$r�zP~;֘� ۵C&y��0=#-��ff�v��b��^�@$�]�RB�:�p�&<��v�7-��R���sįp> 7{=����E�mynS��|�}/^�����<�=�\�F܂7���Ӛu��.̷�y�h�z��]�a�|���nG??՘�.�O�zN����XGI3]�� z��ņ?N6<L۞�}}@����@8j=� ���݄���U��~D{�u)rښ6x�����M�{�Vy_6��3~�r���n�����
��&��I:7z��6g��o�j��]Θ/E:w����|���zH\'̰DpH����\gZ:��
v���Kv�ۄ:�[8��箣�n�(�d����Km�nw
ǣ�uw�ϰh��� Nь�^�g���]���c�#���V����9��m>z��(���1�����bo;�S;OX�guqA�v�J�ϭ܍������z͍l��ۛ�ڎ7p#ڦ���pp�&�+'��� 
'e�rl�8�5u��D�s��\�Uz'�(j.���ܦ��z.$�Y[��w}����Y_O��zk�I.�r��JIuua�	@��~8Dke������PK�'9�B�c�ɬ�G-7��Qc/�U"|w� ��27��{\y� �ѽ���w��]��ح(��CS>A���+`{\�y� ����5<��i� ���7�/k����(�̅s�
Q��_L��Ku�]���7�L@����v�	%ܧ���7�F���D�u�lC#NA�]��ޭ4m$�b|i(��|ֳ{�zZ�}�=̘�@}�ua�I$��h4+\U��A�cݻ�
�d}�x[��v�=������I�"���κ���ŕU-��t`嬐��i�LߖDI/V�4I���Q>�r�{�~��K�)�:�"�Kճ|��A�3J8mX]Jq��χ�T��U���Y�feЗw緇2�Rξ�}�������k���������r&�{�y�=���ƅF�ro�
ً��n��6*Xq�&��w�����}Z�i�	����A$~S�|�@%}j�M���#�/mp�`���2ԅ�a^mY�D���
�R^�ً˼�K1ogs�s]�7��z���w�m�+��x��?��²u����I%-����%��i@ ��K���E��G����MZK�n[�?�-��.�m*��|�K�gSi�R�6������@t���{��3H ���&"�OS�t��bS��׫n�!%C
@T�+˹:��#���E�{1���9�r�Ӯ��]��<X���O\e�#p,7W4��P	{�AM �J��S��{��M���i�e�zo� �����kP���BAJ���)K:���H�n��=|5�IF��A�ڍ FS�̣ ���v�y����
/+c%-�H�=�� |勄���z4��X�yawk7vo�t�ʺ&�[q�>���w���;S3��w'�ք9���װ@4�\e��mn�a�U��ۤ��T(�� �K�������-}�e9�1P��9x�,0Ԇ�j��n?�9��t�J�T�I$2=�w�I%����8���3fii(	�gz:D�#�L���}�>\�������ꤜ���i �s��b{^�b�y���;��Ʊ�3n�*���҅b(�t����ͱ����5�W*��&BւWB�-�s��>*�YG4�KW��{�}�[ ]׵ǘe}|a��b9��w��Y�؉|���b�r�
�]�9h�=�Y}�vP����L@|<���X�ñl߃�ZJ޵E�v
W&g�tsژ���׏0 A��M�����O��V��+�Ն�%�줘��2Dd�թ˫�i�<�,�x=~�b��g�[>��� @��/\-�^�%��N��[9�{��'�D@�����O�ݖjB������7����盚=Mֿn9�42�c]*��[�d�2w�����I���v"C��%���ܖMgJ9h���[�[��fޜ��O����Iuma�	�]˴����=��ꐘ�LQ�vX��<
h��=;�H;�P
ڭAG]$�cr�{��B6_�Vrx;�Y�@w\�y��Ϩ*Is�(�ޏ5����E�Wk�3�;�2�ERK(�a|kKP&�o�a�^�p�+� ����9��=��Z�ՙ�.ri�k�ϨN�,��U�RTf��ן`~�� �x�#���Xa���N~����`#����fj�E��W&`]-���y�oI_���b�I|���@�I$�ŝp�#{ݑ3e�I�ͮ7`�1���X����\�v-��\�K�:����1%7�f�$��n�A"�Iqg]��7t]ck˖bݏ��gGB1��ٝ�<OԜPp{��kG�Qw��?,W'w��~o*����k$+����8�j�9\�?a�����W�t�ß��}� ���REc��緷|дv��Ga�yܜc��5V��l���m���gw,�$�� ��V*��v�97��լu������+%s����X���mw^n�a�ƥ�����^�+�c��t��8yW�y�`���=M�(뷄j�m������y9q���x�����;#n����;ov�Gwn�=��kv��ɳ˹�Zq<j�Z��!N9���������q���h������AIK6����'E��-���5�>��9�pP	 A$ǝl��O�g�t�/�"��q�$ ��4��^�zP���H�v�-9W`] �A��U7�Rc��GR�@ >�=t����y��A��滞~�]��쳚��Oe��(��R���t)%�I/�wH$�Kh"��t�*v���o廮�$P	%fg]�I���|��ڝ�M?f^�kh����f���k�  ��e�l���<̚�֑�����xo�4��Nf����H�m݀�5�wK�K�������y�g�K��M$��v)�醬%�wwy�=�-
�#�X�!B�9e�[[�����홶�3|�vca-i��d�&������I(������� A�{�\��]]Xn�^չ�P�ϗET+�	%ff݊\/���D��LΔr�K���4W#M����i�g��OW�x�Pu���d�'l��w�j�xZ�ʕ��v�^>���0{=t�۲yڸ���"�Ē�|�&W� ���V�]_���R+�[}{��T+��z��)�H�,vd�|�fh@��ǘq�[�EIi?A"PXf��l�WV<�=�2�
�[��W|u�p9��{����/�B@ ��k�0�.���LU�~��������_W}I7[7��1����ӟI"{AM�v�X﬚���{�,$��ن�$I��-A �-�g,��kb2����.���5n�)���h{5 �J¸�'�HZD�j;$��|��-N�����^��� ��ǋ }=�h�=��ŧ9�x�;�]�D�WV��_u�Y#N⑙ �au.�����z��aS�`��W�����������UU�����b�~ؘ,1n�aVuY�$Oj�)�D���Yֳ��|�6�q�"I����S �Pf�\OOmg��>����ӑ��ލ��q�.X34�ʛkuڭ;b�C��%�S;����	�z����Ҁ����c��q���KqU��v�؝y \�����j4� �o�${�1{��j�ZJ���ɵ��[���e9ks3��5��  �9��/�=}�g4q|��Zn�%-�)�J�\^븞�9Ώf�
�J�eQ�R4;\��Y��s�$�y�)@�*��K}��Uenʦx�o\y��@$�ꇠf�n������4�<��d�,մ)�Ц40c�E����,�v���^����ݼ��~����t� ˹�ϔ'����ex��v50�vJ�c�G�ST�A�Iُ,[Iy�+�����^�5������J�˹�F�{�#��\�L�k�l3w�y���Z'����/0π��q�������h3�`݆Gܺxz�zl��2G��T�ٻ�J��v�*�]���c��c��=1�����2���J��>�=Zo��N���|���%���?{���¢(K��sS4b�e��.c۾jＱ�A�lG��� π��Xn�H�:��ra�߆՗�b?D��{rm���	֬u��D��,窭����C��^y�m~u�s����Z�ߑ������{v�_$�����Y��~��;5�+y2j@|���f}[ޑ��U���]~�4IOpDR\�G~I|���R��	.�7$H�^���k���>
\z��'me+�ɍ���,�7�lZI ���ﻘ/�b�u��w��$�w9��f��ژr�eD�TYV�z-�w�۹y��̝ő����b ��ޚ��Yr�D0���fC�{�B��ʙn�$k��<��D�[����w��':��d�PIwT�X@/w5Ǚ� Cޚ��ﾝ�y<��5�%���/�r�C(]}�oNvj�ٵOY��0X����ko���Z��HI��̒{Q3[�+U���R=fn�&�b��9��[�K��W70� _��g�w��|��a{��.��U|y{�;�Y�|�x''g���Csw�>~�=a�ܞ���h.�~��z��g7���W��L�á#��y@˻3����,Rm1�+�y��O���{�`���o<<�P�����{�]�f��z��z�G�� ܲ"��*P�����$V�KZ�M�5P�i�zZ3e/��l����M�{_r~���/zn�w�ʎ�	�������ʮ���� <��i��V�,�)ݜ���o^�h�x�g'ܬ�7��rwk8�����}�t>�6Fp@��~�~��_�����/ج��Ꜽ(aS�~����x�o,�?~���&��=��x������s^gם�U��݁�S	������|�������T��A������F��a�R��1��w�7��,�B��z�>&��b��~�v�t�����Py�E=ڵj��>	Z���Y��cs��a�4u�,��Kf��__;��w,"{�&�(�T
�ޔd4�gk����_I�ޖ�Q��^����nn�4�
Z-�1>Ô�xc�OQ�t��7/y{�����sj�n�z��(��F:�귎ᳵ��ֺzg^1�Tܔ/f��+h�^�G���;�ۜR��}�L>?���;�/�׭?SW[x�1�޵�$߷��L1`��;sX�2���҈�nEL�#I�+�F,��h�6wj��a�IF��~�r�>뻻H$(1��Cfd��.�4��F��R	5���#�<n�n�p����owA$���޼�\+��d��]DC#s��u�ݹ����w}�}�oc�]��J�y�wsL�r�U����s�"��ܹ{�H��{�M�4E&�(���ًݮ�����¤r�/8���w;�,b��\��!E�s��wb<�xQ����]"�Т��޻�;9�+wn"C&D=��sb
wm�)6��1ؒSyv�E��H�W`Pf�	.\��s�/+�B"(���q��8kN��f���**���BMiMABD�&��0][���O�j��\j�
70Z܉���R�;rl۔u�n��N.:�ƞa���D6��e��>�ݱv�q�t2�<F]5H]��:��#q��d�x��s�x귌Wi��[���3�!�0�.&���;��pG7n�n�g��O=�[=<���,�j �qƸ����M���p��Dm�#YW�M���r�1��lW6|i�˰��z�[�\mk�`;z��VI���{l힣yن�����v�N�^���%����I��kuw�'k����݌G[u�J")>L�:-q�m\=������skuu�xԆP���9�<���ˍzm��:�4c��9{m�\��uvx��u�t���q{Baqf�m�Б�b����ݙ����[� N�-=���]R]��3��"�>K�m��:��8�J��ݍ�(籺7b%��N���n��{-+ɶp��Y��ń8��׳�9�m�c����9��Vl����s�c ��<vM��7T�8˒y{m�4ȸ�����\Bh���n�w]�.�v��rvݰcq�����g]	ZN7ck�]���t�a�&+9�ѫ<�C���ќ����WX4�OV�n�mg�����D�a �mɲù{�"�=/`�U)I:��K����<U�{gG>�q���:쏑��t�������8G����f�.���N�&�p��G�cpm�9�[D���V��GY�,�ϲ��ŕ��]��!�����= =�:�p\8��4�=�9Ng�j8�z9�s�s����;<��u``�ryw!��77iM��[b3�7H��=�b�wTn�q/':��#�;v-2������x)��&�!�t����X��c��u�{m��v"lqk����;���ٴqٮ��c�)m��ݛ�.��_1�|�c��{@B�1��������u�v���M���R����|��\���VF�Z1��r8��q��ͭ�ϖ-M
��9糞���f�Z���
Q�������v����>�y���7R���͌�}Y;v鬽����u�u��(�u��&�[��gs�l[ٷ+��,�i�Le��s�j�jեz�q�(���4/7(u��5gsɇ��n����N1�ٛ�;۹l�;�)�c�����e�sqwMA�۰��s�<�e��A�y:(�v6|�]Av�f�p�؀<'���=���9���~?�8�q�8Nn�ۆ�t��˴Wt[�q֛Ƴ��v�c���n׎����������+%��2O��w��� ��s.�`؀]�ޓHR�m�fm��h���<j�Hkr�L��rZ���o�	����Ǣo�{i�[%���xݤ�Ak]͓A,����zg�q��n��T��k��Fc�k�޸���>��#� 3	���n���p�6/wz��� >;zj���>����W&7y�����}�3��<� �����M�{6gy6���׀%�k[y�]̜��T��vU�"5��$�I漤�����$��Zl�my��B"�E�ϩ>�\��+�4r��m��@i��6����pv`v6�]�[7��q�Ԋ"�����J@��=�ʳv�� �w�T> ����n����ꦚϒ%.k���V���a������p���9����A籉����t?8�� w~�i�|8�����"�7��N{�fC�p͍%g�3l�`����+&�?�I,oy�i$�/~�����zn�;��u^�w>I�?s-#r�rZ����5��6|���D��kgs���� �=�F�_'���誷S4�Hc2@���z��z޽�y��8�� ]�P��S>���e�^ߧd��X��pyQﭥ$+�ɍޝ�,���y�0�ᘮ��FIT�sd�I<[�q�[},��>m���<un�����T:��{l�nVn'm�Um��ӟJ��j,t����nʤ�����ryP@�b� o��X޲۽@���$=믨��f[7����J@��LΔr�6����t�9��*g��o�M�RbхB��u��C�i:!P�P�VQ>������1�eB�q�����4Ӯ�<M}|�f��B�������ir꺼�aѨW��}��z��R�T�\
�������+FT�I��翿_]~l��7պ�y��:iГ`�7,��䥷t�~�q�Ӫ�k{�a�����vxc�x�CK�ӰX�Ik��H������6�I��%e���u������XJ�$�2���s��:�ǧ��oM4��ۭ/!�:�>��ͧn��|�=�_*����1eeB��T+�kݝ�4��T**�����1��P�+P�)p�_�ٴ}�b�T�� �|��#�Y��ӷ�D�J��w�^��i֝kG$�u+�y�w���%ejJ��J������m��[�����9�1F
��5���*LC�
ʞ���!�teB��*
�/��m&�����οX�~������o[e�������!u���mW���޿T�l+�C�Dʀ���W�Ͽ]kW�sM�Hq&!��滰�z��[�R[�Xy���x��IZʒ�J��}~�f�i8%IY���=��5�I�u��s_���a*L%B܇������(Ҏ~˲u;,r��g�m*��*]߾ٴ�Cb��y����s�ǳ�>u�5ݟ�:��b��{���C�:5
�T��_�ٴ��I�RW߷��{{���ߵ�����IP��YG�(Hʐ%��#��»�Ոq&3�IP��Tϯ��7�&Щ� #�w���*�j��߅�@hT�T+*~��;�C��eB��1
%K���C��+�>�-�.��8�w�#�@G%N�f���B�!�?��5Fu%leIR�IR�5��6�Iȕ%e���ן{��x���N�%�F�q��ߨ�B�T�xf*��)�)/b�u$�1������.�s��\X�o��+<=��Sp���=�����1���S87��dv��<?�ﰿ�����V{�}�C�1{���٪WZ[u��4�S�/לٴ��Ь��VQ�
���~��u!��6��yh�8�@gῦz�����+
5
��/���6�HbLxʒ�eu���p�tM$����_M{��߻�z���n��	�$V�u��Tr�U���u\n{�9\=�)P���E�����X�]�~4��1�y���g��J�5%Cbg��o�h[0�
�¡[5�������@dGg�ܓ��W���?O��w�ۨu�eB��T*LL���f�Ϛ�J?�J�l��)l+,2���[�B���wp�&!�/�����N}�u�����׼�|u%k*J�J��/�~��i4�J���%ek�>׻�P�1��zw��oz��}}u��Q�3t����[ �|��Z�h��m="B���Y`ʅu�����B�B��1����>���َ��^y�}��C�5
�Ĕ�_o�l�M!�1�*J�W^}�w�SI*|o�>�P���*JGȏ�¿Wz���Q�F��5�wi*��.�j���h[��T��7^y�9���*(�B�����u�x뇺��ǝ�C�teB�bT���f��M�X';�[��\�.����tj��{�B�����V{��u$�^�������;<IRĩ*Y~�y�i4�$�1&3�u��p��J�$�2���{��^��W$�w���O�oާ^e���G���,��%~^���q0�v�W����3�˞����`>���E�dl^���ۿ�> |��h�g��j���d]��Lh�[���q�g�QλN[k��đrE�G�	��qـ-����c+��u'R7(��uݸ��,˙�cY��tcSڵ��^)gKC�@�:��6n�t�}��ᵺ5\m�;wRrv�m�m;�&-���s�A�]��tmɻC���N:���VƄ`&���*&��"xr�����.ڮ3r���ٓ��ŧ�ֳ�v�ɼ�n�:Q���:����j^������G����Тp��eB���W_}�{:ΡRb����{���j�>��>���Rx��6m'&�*Lk*J��3�mW��x����w���jB����I:�0���\g�ԕ��*aw�Ӿ��9�f>��w����h[��V��V�w�y�uI�bLC�>���P�:ʅeP�p��_~��w��&�df��B��?%+:�5�sW9�:������B��1%���<�����J�T�(�%FI����S?�W�I��q����op93 .$1��s���01�����4�m����#�;��n���������:ϙP��*�=�����&!�T�V����P��B��B�����I������5����L}eIPǟ}�{��T�/����3kN].k\:��Xo���Y��%e�IP?�2?7�B� '7�~�*�w~�>Dk
�{�}���1&!��*����ʅI�bLO����!��~�ou���~��̼�jm�b�*r����6�by�y��`�7���ǧ�ql���ѹ�����I�#��
?��9w�_Cv�T�\
���cѕ%J�%K�Z��I�1&3�מ���t�u�v�Hc���Èt�J�S	P�!��O<|~����� � ����C�1>�{٤�!�*LC�|�r��@�g�N����X�\�=�>G��?z���_iA4��`G��z�f�iV9<Ƕ͊|z{�D�̥�g��!�����?og�:�BĨT(�
o��C�:�*LCR������$��I�bLo������>oﷸu?	RT�����u�n�֍kG$�tJ����w��ԕ�jJ��J�[��5ɇ�@d|���dq�I��{����5�~��1<�T*T*�>�������
�2�P�*~���C�m
��gs��sZ曫��a֡^}���^t������I�bLC}�7���gRV��*T�*S�k߸i&��RVV��c�>�{�����x����o��1&!�>߻�x�H¡W��l�-��m&⿇��"����$���VPeB������ΡP�}߿y��~�5�����BĨV���s��
B����_�l�N��1I�������N�RT̻������
�R�#M�<��P;���ݭ��t\lj��d`"�K������y�Q��5��Rb|%a�>�w��=IYZ��K�����ٮM�i��T��7^}�9���*;�3����_�������>���gFT+,eB�R����� Y@g��B��}�q�pH��a��+���{�P�1I�x��_{����<�w���:��eIR�IR��k�i&��RVV���u���p����%B���7���[|���7�C��¡_(���3Z4:֋�T8��T���l�M!�1gP�����tgP�Q*
�
ý�i��~�j�wְ��f��N!Oq�/W��֑�Mu~|���?c��5��`��t�osg�V�p�y��aCzT�h���3A(�����b�5
µ
����٤��I�bLk+�?�����T�݁�&"�2����?_�i������u�"4>dsw�%��!i��V��W_}��!��*(�B����s��:�u����_����<CL��T(�>��6i&��G���Zp�Y��a��+Ͽw{�P�1Ie��<���x��I^{�;�>��p��*J�J��7�}���iI�bLg�����uI�bLC;�������T+�ϛ��߾��u���ý\��scW\5�m���%k�Ɖ�f7j��pޮnT�&{9���m����@�~ 2oW��4�Hc8ʅeP�����!�1C�T+��}�!�j���{��|��a��hlu�!B#�lʒ��׿�op�u*J��~��n��u�k\:��V����c:5% U_�_�5_��7+7Ç�G7�B{�>��J�h0�V����9��1N�T+('�o���teB��* *���oY�"c��!��?/���8�m8$ud
?��_�<|B����1a���Fu%CbQ*J���f�~����/����$�|%IPĘ���}���:\%CbL���wP��
���ױ2�њ�o!P�v!S�^sf����s?p��<PĘ�3L�W~w��!�tJ�BĨV�ם�C�;�aZ�I���~���ol����߯ν���˂���Ⲍ��M�����>�G���x�%�LZ������L?�O�GY�C����X�>՝��!��e��g���|�Ę�A�������R��B��?b. ���G��?�Y���z��Ƥ�R�*yo��4�Ha���ת����?A߇�@�>Dxfg�� "v!P�1eϷ盨u&!��*
%O�~�f���B��:���y��_?�}o��(�g�Yu�g��g>ݨ�rs�$ҝOF���f�ZL��e ����RV�)(+�?�P�>��8�$���1a����׬�Jѕ%J�%O���I��3���;u����s#���,�~ꯇ�t�J�S	P�2~�o��
��wt�z]R��g!�4�V���$��`ʅg>�u���y�������͞��B�P�Q*��|ߛ�8ñ�T��$�ڿ}�I9�
�������v�s���W�H�"�#E��F�Z�t��l�LN�Xw�����+(ԕI����ٮM�n�ZF
�o�������y�?!S�B�Rb���7��$�1�eB�bT����4�hVx�L�̵���@���dr�z�۾uX@�k��)p+��o��+c*J�*J��Z��$�r%IPĘ�:��}�,�;����]ג8>���̀��f���C�F
��}/L\�Ӛ�o!P�t��W�٤��Ь��VQ���͟�x�� :ŝ������Ɛ�ĨV���7P��B���*J\=����$��*Lk*Jє�d�_�!2#�|�.?�����&�qKp{=�:��K�8��.yy����5^n�7WZ�{Zc/ް��"�;y%��V8�����Y˦L����ϻ�7�|�]���<�
��z�ϙ��a�K�7�(C2����x������9�z��q/M��kq������0�g*�2�;r���m�-{sk���@v�׃����sks�Is�l��\r.k7W�J�:��u�;���]u�]^���n4me���Jm�n�ۇ[�1���pR��~b'�`�֋lc����c����n��f�t%f���p����Jx�[����<��1��sڠT@�4�\����:�UX������c9�����=IYcRT,�J�[���hZa*�*�|�ۇ��*8on�s>���g��=g�w����gFT+(ʅB�O5}��Hq6�aMl���n��u��!��y�~�à�
��
�߮>w�gz��k�7P�LCb�����$�|%IPĘ��}�èt�J�\>d�0p��z�{~���d#�@G�n�9AT�Jk�*�ZQ�ߴ�_T1�T*LC����!�v%B�2?w��)�m���ٻ́���XX�*Kp����ʓ��*Lk*J�W����N�RT�Ǟm�G-�7	rX�"<C?~��3��N�/ӗ�)=g�IPĘ���/0�B�	P�aP�����!�1:�B��1�>�}�u����nwG�o�[�g�i�eB�D�����4�0�:���ˬ�m���P�ơ_��w�qI�bN�
��u�w^��+�=����x�=I�1&%���xT�N	RVXԕ�k�����;.��	P�?}����a�w�/t����`*C�$�
nFy��uW!�<5J��ے�������������\�u��s�T<I�ܻ�ʟ!�+,eB��1��ogc:�I�bJ�a}��ʇXvB���hk��ߟ=Cğ���k�6T����1�*J�W�ݪ�x�|C#�C��3�	Abu:���ߟ�Yש++RT<���߀����m_T?���]�lCҌ�og/_f�I�v��/n�Kۻ�����Ib����N��O��Z_*�K{�w���?��zkw���?���^���a6���Z0�V�w��9���
�K�VQ>��}�C��ʅe��R�3�_���K.�2>�~��{�n��u��!�j�?~�ñ�&!�).a��ﻨq&=RT1&&�WG<����f���*M'�RVQ�+(��������*f�nC��o��-�����{���ѕ�L�u$��_��S���������:���ʅe��W�}���gP�PJ�I�c��Ｈu�F�XQ�T��e��Gݓ��oi�`G�����,�ϳ�����J����iφۭf���[8��V���ΏRT1&!n��}���gMw�Z�~m$���������:�'D*&!��?{����Yѕ
�ʅBĩ�5��*M�3�:e,�߄�|�,�I2+�9MN۩�]��Ӯ�]����qqt��%�.905�~��ؓ�6ڂG�H~� 3�~��Y;p*LC}���ѝIPĘ�J���u��*M'"T�������%ٛ;��!�����Cۄ�e�J��>�}�C�XT+~����0q�u]9�T:��T�5�l�4�3�eB�2�ϯ7�*�߻��7�����7���&!�1ag���y�u�cP�+P�)p����'&�*LCc������m��op�=��|��N��t]5�8i'S�X~���gG�++RT,�J�e�험M�n�Z¡T�=��n�}so������q���a�{��ǄW6��w�~� <����|�;�
E�����[��u궰o�?ֻ[�6S�����L�{Fٲ*����0��i7��K����@��8������x�=��v��M��bZ�E�'ݳ�y��`������G��ۀ��s�=��ǖ���1�ش��*0d9*�:a�[k�(i�E�J��.��ԃԽU�z�Ě/�I��^{�Q|�᫧�i��Zm���?P�{=�ij���r�ʝ�}9_�Oj�qwL�+���KA�����72�7+hcM������v�����'N<�\�sh������gh8�|�=����ꏟ���<�W"�^�os3�Uo���_J���_��|K�7���>�|W�κd���aQw�2�kB�zzOT�x�f�]WŰ��>Z��au�9Y�h4�	cw��k�.�"�����{-w�j�4n�xt{v���+��*�,��}�C�yg��FT���λ{c�R�ǉj���{r����m9��o��K��3����#)^�Sy'J�Ē}�/sW�;�U�@�v�ٲAT�~4�7����"��%�>^w�yS�^���it�
.�1quE^>Ь�m�ذg�TÚ����<3w6��u��W��I-��p���{F���N����H�s�:�[��z�Dξi�UK��|8g�*��J��N���.S7wp��a���%\oLx���/�",Q�da�\���G��]�ur-vi1Ir� ��u�v�{��
lwut��X�71��4�r.n�+��B�I<�L؈�r�2D��o�\�FA0���91���t�b��b
+�f�5��{����S��G����G���c!�m�[�j�3&F1�331A��;�rE�H(e��/��I
{�]���E�;��؉C��ܓ��&}�r�W(����&��s�F6"�v���ݹ�w9I��-����]{��ۥ̑�s�r+]�%��4�q4cDl���Es�ID�αEo.h�-����E��sk�ȸ�9��,�&
?�?�u�vC�
�I�c*~�=�!Ԙ�3��T*T�5��ʇhV����ؙu��\ x�< 3/U��p��Zh�~P�'�RR�Vߛ�x�gRV��*Q*J�����*M!�1�G̀���U|,�UܿE��e�&�~�fC�}���:�aP�=��4�tf����C�i:�M�}����2�YYP����{:ΡP��>�׿����Ͼy��!��V�;Ϲ�u&!�:5
��_�l�9�
�ʒ���/�W��x�G̅�K��`����#�:��v�R��nwi|a���q�.:�h�4v����7K.o��B[*��o�ƾ��������tz���%B�%O�}���	�*LC¡^�Ϸ�qN�T*?�(8�C�0�>�/zs#2���I�bJ�f��eI�1�&���$�M���߈~���U���� ">w������!�~�Ք�I��eIPĘ�����*M' �%Cc(׾s��C�p��J���xw.~�~߯ԈGȀ���i~q�sF��*N�*~�s�*p���
�FT+��{:ΡRb��d~�y{���q���D#�@��B�������*NM�T��ʒ����{�PĘ���xt�.��tkY���u:���󟷌����7Rq��RT-�T�_���a6���Rb��>���1:!P�P�VT����x�����z�.C���#k�"�_�~��}�g��/Dă���a;��v�W]����:��#�Y�d .�:�>�8=��f�|�s.��O��?�T**f���P�m
��l���Z3-�g4�Xv5
�����8�$�p*L@��?������|ɠ�o�f��~�>D`%IR�]}��I������+)��>���;p���i���9���|~����~3�ˇ�����hB�f�uۧi�pب�۶�
z;O�B�;���V嶣��|�8�'QQ����J����|���"B���YYP�߹��v3�T*T*LC_�����B���;��3���;p�5߶T�7�RcFT��+��{�éԩ*_�;��L��Y�Un�é1:%a߿s��u�J�ԕ��|��?o�I�\����a6�I�cXT+O߹�9��؅B��1�>��{�C��*�eB�u~�������7�s��Wm@�@g�E�Ѧ'
�5���D|���u@h���Ȗ��1����w�Yԕ��*T�*sW�����>��w�I��	RVQ�++_}���Cb�%B��߷��=aP��>~oLisUӛ�C��
�j�4�w�t�������C�m�P���W_��{:ΡP�P�Q*�?w�=�!��aF�RR����B�����9��_{��(����̏�c+�|�{�S�*J�}�Ә��tj捚I�1������=IYZ��e��F7��	a��������-7��x���aP���s����T��B���~��:��T+(ʅBĩ�W�i	�+w���}�ߵ���O8��n���6g��w��ޫ�A[&w�3�[$�Wõo��+�5�X+ ��{EU�=37Z��+�SV_�s���e�m7'?��>^p�����]n�^N݉�,n��W�f�\-�q��:��D�6�{&g�=�}<ų�i��s����m���b��=\wg��GL�۬w�e��-��#�����p�<Էm�۸�΂�y7��p�nnW\�l�\�3���8�ni���Kk���֎����#�P���;͹�u���nwe�c�q��k�n�^V_/$�c1�p�m۵���;EDn@vd��U<�����uR�����R�RP�V�0��B���7���*J\
��
���߻ǰgRT1&%J�����f�i8�%f�N����{��$�65�>��èv�*�ː����:�0�VϺ݃���TG%3嶕km(֬��J��B���V}���y�ֶ�����>n��{>u
��(�
���~��C�1a֡Rb~���4����1��|�/���W\����UW�H�C#�C��]%�8�0FK�ǈ��g�鿽Q$�1&!��*}o��k�hT�@E��dr�����~�w�_����� $�
�!P�=����ѕ
�2�P��?j��f��M�XS:oߡp��PH��
?|Y��ڠ?a4L�{���#�@D}@3��Fu%k*J�$��߿l�M'"T���+(׿{��C�w���<�|�y�<מ���*�7���z¡[/�����2�Z��r�A
��y͚ND6�e��T��=��w������?f�~@d2?�=�:ãP�,j%.j���$��*Lk*J�W�{��N�RT��y�k�Wrd��o���P�Q1��r0K:3'\s����a��$LE�:���>��~}^�DѦ���OS�+5�>ޙש++RT(\%O-��I�1&!�#
�{�����1:�B�����y�}�x�Y��^���Yѕ
�P�X�<���J��5��(����[������B�����8�$�\
��7���x��|����R�<z��Wba��N�(O�L�F��	���7�f�Ҝ^�}�d{>�G<��&�1��)�w_���_�~ޟ�IZ2��D�*_�k��$�r%IYF���{��w�u ���C�@s���;=�����I�c��{�Zz:3FV�g!�4�B��~�f��m
�P��*��?opY� "�d~��5e��y~�[��o�}�:�֡XQ�T�����I�x&5�%C��w�q:�%K��R�S1�h�,x�� �~������O3�O�s������=f��*��}�f���&!�T+o�y�uN�T*Q
�a����Hq���{�|���ҡ�Q�
�J����C�m
��=����]f��ѭ^u��j���{�B��p*K�X}}���x������tO>D}Dx����L�bi9���RVX׻���C�	PĘ�S!����z¡^}��-}�]��K=޲;D��c�����X�g����z��LYr]ZQԡ�6�m��������������B�����'6�eP���
�}��gP�1B�P�/�}�y�:íB��w������r���!�J\7���4�HbLyRV�+����éԩ*P�����hˣW4p�N�bVk�~ޙ��%ejJ��o���u��鞓�ݿsf����*�
�ow���:�'b
�!P�>�s��� #�����\������e9�ͤ�����0���ŷY��aѨW\���:=B����1a����OYԕ�ʒ�������ϻ��8��z�����Ѭm?�U˒�S¡�XtI�ɮ���ko�5�[������^Y�v���9u՛K�������Y��]^�s������m&��J���RVX���op��	P�a*����w�:��B���o���[u��B>D(�~�D~��o�r�Uo�GȆ$�1�w{��=J�B�P�,����4�Xu�V�T��_���6���yޚ4��T��%leu�?op�[j5�j}����d�R����kiXw_{��$�tjJ��J������C� ;r���VU�/9ʫ�'��T+f���:�$�1&!��O����Hu&!��*&&~�~ٴ�CgV~���w�OV)��r����}M��Fwr��eص�t`lUQ����$�h���|��JHU�_�Ci1u�����
����1���<ޞ��+FT�,J�������i4��RVy����~��I�x׻���:�e�T2�%B����7�8��B��|��Ц\u��3��u:!R�y͛ND6�I�c>���?k�_�����7��6zΡ�*T*�Xy~��aѨV5
�>�~ٴ�7�RcFT����o<�~糯y湸x�I*Y��};��W.�\��I:���]���΃ԕ��*�J����I�3���T��>�:�����3�k�x�I�b{�VT�^������VVT*����f�ia�{{��[䡕����q��n�I~�8�O/vz��CԜ�%.a���zC�1�ʒ��RT��k��6�Iȕ%e�����k�èRO���������'�V	&�{:�|ΡB��(�^�N!�۞�}�-�'G�[XǷ[|�݄��S>cE�e���*�6x3K�+t�kQy�S����H��/��gT x�ǻ���oˬsFV�g!�4��T��l�q�Rb�ʅ{���u� x�j��0m��j�b��4" i�X_��~���P�+P�)p�_�ٴ�Cc��%h���=�:�b��l��|.�����q���P�ࠡ�d�*��q��v���Qsd`�K���߯���.���s�|z��+��{�!Ę�Ƥ�[���_l�0�B�%B�0�V�y�ۇP�t�T���c^y��gS�s�7�:Ό�VPeB�R����f��&Ь{��uq�k-�����
����v=C�,.I�ܖ��؎K3@����������*T�*g���6�I�*J�$�V�y�ڇP�LC;��Y'w��=�����S�ͭ�~��#�8|�; ��FB��!��oz�i�#1 �����`�d ��!��X�[U�e[޿�C䘆0�j%.���I�1&<��+Y_���C��N��C��>���E8#PX�}�<C?�3���v^�OZ��e�T���vo�h[0�
�¡^�ߵ!���T���#���P����X�/�w���"?C*
%K�϶m&Ь.�����uE��Y��aѨW�����P�K.IB�V]����gRWϮ���Ϲ�"�Ę�/u�8m&��RVXԕ�������:w	P�a*��_�������u��ym���Db޼_4�F'��!���ť�{���1T��ڬYs��o�xwKsB~^W�L���b�e��Yݒ��~�����b�}ۏ��xSq[1���9����8�d���n�
�u�[
��[��xw[Bq�h����;�<r�Ϛ��C.:�Jd��1+ݮ1�''l�\��/�:�������q"`=�n�cE�0�ю��ky��	��',��sИ9v1 u������;U�=X6l�v�(vciUk�;���]��vr�����69M��k�n�\�GTKE�ENKX`6��=Of�q����?s\ڹ5���&�������F�����q��T��~ٴ�!�*LCYP�w��u�B��1
�
�ϵ�����x@g��~K����>��@�>�\/�}ٴ��T��$ƌ��w��i|5��wgXKdv�r�[k᭵;�>��νIPĘ�߮��os�W��J����I�3�J�I�c|�����T�T+(����ސ�:ʅ~`���X����ͯu�78x�o��0� 3�a�k0�I���@���j����ñ�%���1��~��=ԕ��*T�*o������ߎk�M���Ę�5��~���;.��1����ސ�хB��|��陏�l�B�� 2�WB���Of��m
Ͳ�Rb���~��Ρ�,J�BĨV{���4�RbãP0���D}ه��v�a~>��y&;��+FW�<�w�D�J����8j�r���4��Ԭ>מ~ސ�LgA�*�*g���7�	�/�O���﮹�?!��B��{��Kۙ���{ya"I忥E�R���P���Z�y��b*����F뮍�]�86�C����y$z7e�ۻ\�2A^s`��\��"J�槳�@!N�b��$AsΎ�\ɾ���w�����A��2� Z��S�u��e���J-�C��7�����^��z�<����B��q��4��7�w�7l嬘��h��XŊ�#�"�����=W�!���� ~�_~�	 K����~9���0)�ݭ�=��w�7�2y����[��oڼX~;۪%�U�F�&�Fz��{&�	$�͹X�s�J�o9�]��*�j�^vd��776�i��ܸ� � �Ott�I���YV'v�k��x���n� {`w+�'Ņ���<]]PHuy��~ݸxUջ���ԗ�z�]��'�t��H�y�Xi�2��`d֦G��8���.�S�� �O`n9g7dN5;]��&J�%�6��"ђ�
���s{�� ���m���n�A��˕	�g�����ӝ����]o+LD�&Z]t�퓾}��]�ަ��˜- �$�5�Kຼ��7�_uŢ�ɞ�mc�����Jdς��� +^ض�I�[��(k��ɩ�Z=���y�4Q���.�+)�`R�<g�:^��{��W��%��i�J:�ĳ ��RJ� �0o��BL�⿳�ou|�� p�믨���nw�{Nd�@��$jPBe��g1�\����˥C�{]�ш=}�4�k7��8j�D��J�w��P�
iA#��y防 �̘���������S��@|���s� �/�3>��w]�cj�4v�+�� NB1"��g�Oi�φ�ݭ�*���n"�I��|k���������<M�˫�A >o'tg�|e��bH�:��3F�	R˕I ����0^�|�++d�©��M�Ou{y�}�t���gt����[�D�|��3>����x�v��z�/Ay�mJ1P��.N�Făg���6ݪ:K�K�)��$J]������D؜,�[Ԋ6[�݀�[�6P��9ᕓ�C�l=%|�z����$ŵ�W�I$5��sq�{d�LY�<����v���k}�.�Tͭ]�nA^����F�]�+�Ƭ����x]^�u�^�;�SJ�HUYڴ�o���|x�#�ɼ��N����D[t��Os%�D��%��*Sˮ�?M�$��Y�$��������Ҧ����^}q�y���v�B��HY#+R�DA8�<���qu��ݪ�pD��-�߽�v��[9}�]�f,���5�0  �����]���f���g�{Ё0�~�K�H�H9p���G�<���m-�o��ۀ �ۭ��x9�o܆���߷�.a�:�s'��p���2��;�G	 S�ɢI$�^�����[����Ē�r�f7��z�P�u�mJ#�;'�=�d�kU+]����Ww4Ѱ�I/=��$=�yV2��R�C��ԀJ{z��^��g����L�wJ������7�m-�[�&S�Xm�@�z�@${[���-��w>���6w�����~^˂iEy�%>��t��{,&?�$�$�5��Mxo�1�CG���A�2ژZ�J�OwQ�{qj�<��Xyؗ���|��nv�|��:%vA���N���ZC�� p��m�+}w��݈хg���ob4�S���G ���|��3.�'ov���z�e�ļ�7	ѹ�ڐ���b�}�ߚ��4���ւ2�[��[��L����&G�r^��^�(э���m4n�<�U��'k�.��f��������!�yI�Nw��:��	ɹ��'�����ڧz�!��D�u+NM�L��6�����Հ���)n��m�g_{��C�<��:i��l����4���}B~���~�w�k�8�O��ͪy�e/3א��f�q�����<�n�����bX�����jjwա/{+}6��j~�2X�`��N�onTY�%z�̞�֟�|�?V�NwMu�T5I�&/>�)��$���ޢU�쎬Zv'����� p�	67��S:zy�:Tفrd�g�'��������b�pW�g���I���e��ވ�r�(c����2 ت������yf�{����+���>���x���D�n���{Oh(82�{�Q-���c��}U��/{޽��ux��G��7}�ӥ��k&`�N�|^��$qyw��O6�ڗBP��C�$�G���|o<o�@���rݹ�����yٓH�+To;�qp���vnL�Z��g����y{Y����/Rܰ��ʬܘ���U��j(5 d�r7wnj-���ͮ��F�h�Fwn����b�=�P�&�#cc]݊���(��guE���<��(�N��p��sm��#F����N�nUJL�k��rǚ�KF�4b���t�q}ޞ+�Ԓ\���᰻��fZ�yp�;���wE(�ֺ���NWJ���IŤ�4hf��Ε|�d����\���sj��F�m�4ƹnZ.b��t堇u�R[�s[�_r�W�t^G������lh؍G�Y-=�5r�c���^W���_6�#E�������+���c�67MsO�����}�!���a����2��Lm�!��I�>q�Sڎ۶t�c��,G�I:-ƈ�1{XN�)h�Z7m��^��Ls�tt��<v�7X��l�u�m˸�屶��,jh�J��7O 4�-�ݭ��937�֪|���8���W$����$q��1g���z��7=H-nphǏX�ݮ���]���L�Du�sƸ��\�׳����<�ΘS�.^0�jMn3u�7�*<��BN^fۇ�=]u��ll�g��in;wY{��)�8�:��5�-���۷6�s�A��Ol��Y����ۯ.Ciy��Ϝ��gv�^�ssں�{Kی;��`Bpm6w�lo��8U��ѹ�^�G>ޜ[��^͹J.l�n�95ŉ�1ۂ�A���-�m����K<�ѝoj�W<;`���s:��,]�.��R�n��ϕ��;�;woǺ7;�Oc���z]��j�7��=�#�3�u�n9G2���3�:�{'�|�zT:Ϧ���5��Rc7�>wφ�ݙ�k�%-ݸv�XxK��7F�O/Uج'T�Ԏ�q�����xN�<�Y3�σ�v�vɤ���(�で��a!��n+��m��L�v�βJ�s�i����YԞx^e��7���U�Yϗ�۝��I$��a�<9�Nɶ�:�+����0��Rʅ�3<�uݱ�FԘIZ�AY��݆�uہ�75�c��<�dZ�����v�.,��mbny�\��1�v�[�yspk�S�����ٻ�]e�6odM���1����^���Kp��;\�7\�]	:�e�sf7�H���<0���*�
UdE!T�h�i�S������,n�
[�֣<l�Y�q����OnΎ�n�k�'8{�t��,N�[d�"b�	�[��A��w7g<��a�QE��u�um'��g:�Ů����Ti2�m���V^\�3�'5hV�T�M@Y�m[d�yv���gvz�6���#C�.����s��u���kj���n�nٸ��2q�����`�8��r�@wh��G;\�
/���rBvHf�k�]aA�B�s¸��ܻ�x9�G��m�r���>��RA��9��:�n�k�i�9C�64[ӻQ�7Y걹���Ks��kp��q�7\�6��\��.�z578Nt�7]�v�#ȭ;lqUύ�Xע+\�گN�M�z�����cC�v۶�x��9��y,ܧIe:�.�vͨ���0���5�Vm�۴/��e�`96�]W]4�E��Gj����~���bV+mm����u�0 ӽ���K��m�V���z-�{���M�D��ǽuA5����,�P�ٗ�3�h% ����k}u,�Đ	 �����I��mks�7�E_�~դ�͌�W�_�,���.�z���=��I��^��ǯ���	O�쨊I.�=�i�KBS��wk�=�����uT}�K[�H |=��A�5��0m�	��sӵc�s��p�.�u�mJ IB�sS�� �wC!�Sw'�z˄�·�Z$���b����k|�i�њ�&����!����u�n�W`���ls�su�Y�n���X��x��
�#�/��ѳ�0*��N�Û��H���N�%}�u�'�=�=U�\��p��oHf�{1P�3�J�m�,�l*��W��׏}]��)˫�.��n�n��˖����-֨v饿&/a�y�h�ˀ�ҟNCޭe�9W��tz{e8����Ys���ޞ��{}���_>���� .�{�L�>�����^5�-��^u����5��c�%��U�.$��S�z�a����)�ٿ{^����h�s(Ā��0wc9��/���.����yە=��	$�+۸JI�e����$\���{�E�{{=�5�?a��*�Ѵյ2UT��û��	$O�&��?P�Wwl�ل��/[�3 ���]*rfy�y�k2��o�l���[�N�gGdpB;<Z��b��.�VF�b2��U-�>����(���׃\5�L���f����Y����7�1��[v")%�u����V����0*��L1 �}t����ֵ�'�|�4���~�  ݽ�1�5oFM�{�����?[7
��'2�Ym��5��3� ��n� o�������E�b�Gn�4����ut�;�'��w�}� lG�-Mn!����y{��M���d{�رb}?�^��|���{�` ��X����i�܊D��ܰ�R��=;�S+&wh՝٦�$��Y�@����xe����%�Iٜ��K�Em�w�e"s3��uu��A|oز�k������%���1�NvꍱǶ�E�y�]�s>��BDB4�(nKnn��	�V^����cuF7T�3�A؁�s�:���J���7��y���ꍶ_M�& �&���*f��/8f|��z�PR�[�ԣa
05�^Ŕo���]ޮ�{��3�?�@ ��H�?��U�[?_N3ėr,$rN2�9i�=믕 >�{�E���K����Sm�9�0���.����
ARJ&y�%Z��mn��?�@|�{���}�UC�v%l�.k�ཬq�9�2i�T�>$�����[(ݳ���"��B�����ߴi�*�;���yoX�{&�w����� 6~�u���ǉ$���;f�|צbY�s�5n�.������Lݚ�w���-��]���|�ݿ.�[���Z��H�F4Q�"GRk�2n����n_j]nk�;U�pu���[�xgz�j�[)��p��� ��Ԭ$����Z]µ��n�t���z�Q� �{��Ϡ/^��jZ�UT����z{�H$E�=Z2W+��ʤgR���g��}�g�$
y��{����Z��D�:��d�)5�Lz�>� ��3�[�oފ���XN�jL >/7;��g�������|��c���aa�M��N;���󓙐@ >�ٙ�6|z��,�:z�.��@���y�1�$��-"-����Tq$�]E���~�۸=��/Va=Y��`��y�0=�G��x��\�:	l�C�l�=��l�V��8���˝��=������������b��:}/{�|3v_��l�~���u�_o���m;<rH��s��^rs�L���X{v�F{.GV��n�v�@8Wm�[��\�焂�{q.מŹ�5�1g1M�^^�it�Ƅg���]]��.c����)q�8aɶ�� ?��u�ɻq�a�;]��pL<���k��@�z���m����/n����F�
�l����<v��a�]:�.V�ms�kˋ���<m���ꗍ�V��.ŭt)��0���<3�/ɶ�2Fّ�{N��  �ٟ`  ��Շrj���Of(1�}���j�5l�Nk>\ԧB$��റU�����	��ʉ��As[΢)!�9��
������Ե�����L�ŀ��令�Kk7�����M����%�Kd�W`$��w�T%xu��R��(\ςk�=��=��	��W�J}ʍ��	rY��I$���8�Ҫ���C�PK���`kk"p�F妌,;館���F�Ջ~Hugb�kC$�Wi �X��(+��v��{��&�W���ӳ1��ډ��%Y�p�0�q��[�\3ێ�:���ܣr:�����Y
+c����#^�����G�l�gu�/.��2�U��{_��$������82��{u&\�6dw/䶶�	ee��}��z�9e��j������VE��^�5���vf�T��*�ͺ�F���Uz���[6�~��<�ҥcwK.؛㶳�ﾷ�9���I����������H}����<ځ"[Ǯ{h��!#�js�Y�o=s��O�k��&�6{`�=viQ�#�����5`HHp'J�[�W)�����'��צ� ��szǟ �f�ش�Y��t3>#����%|�M�Q���A���X /�z�ًWW}]�k�Ԛ@ o����b���c=g�J�h��&S�$.DX&ی�4D��;q�z�r������:��3�Zx�������G
�nZh�Xo�T��wq`|	%�;��*ɕ����5�l�	 ����w4�RV�+e�������7߷�3Z&��J���;�� �~�BO����J����h��/�3�I�9m�;f\�/�ۋ  ��6i���0.�Ng=�������K[�^x[������m_�����[^����̯{�a?	����f�+�xn"��V�hv�*d���V�KBc���7��O�|�]`6����3 ��m�Y􄸜�v��M��*Rc���ڒ�^��>@ ��X���=5Mrwk�n=�p��]`sS�+T%D��-��*6�	y-�B-�{�M����k��^�sX��}�b ��y4���ʕ{dϵ�ɍ�$T�L��|+v�/�m�ge�r�u���&c��8&S-	|{�#�.�$�^�A�{wO A�Oa��|�����I+B��$vV~�X)$\�Y�{T�+*�r�E�}#o�Nu{;]Q��VWVS�D��ʘh�	 ��k�_%d[^�wQ���=��ߒWsm���t��ۧ��{�}� x;�x��NΗ��%��pv~'��а�z�Ҡ�������+g.ƷĬRVA͊��D�9���%|Z�ku�I$���싧�+�B&f�o��G1���=6o}HI<����v����r�U�9M�b��6���*��%�7y�����|�����3�$=Ӽ���m��ա%��;���R=| u�r���[D���<������p����Q���%����R�9��v���B3�|/gh�g�Oksy���m�:��g��r֑��b�Uio=�A]RJ�Tx�߱ݤ��/%��%�$��˻#V>�g2{��׮� �ݨ���q�q�@�ue��V���G�q�r����I#�{��!�g�� ��(ez@��]z���C����N�r*�a��?�o�Y �c�N�Uӿ�����L^vz����6�&�1�\�TY��k� ���B�~2=��Y0���o�����u��z�Ẅ=�+�E��KB[3����|3�7���_��l9�b�$<�������}n�>�"���X�Kj^e�s����l��G�<��,'��ά����%k�!���c�Q�EIӁ���q{�wf{��G�������w�����g��[k�dMDR+����';1㡛hN��ʗ\vݸ�pPs���u����u��:Cnܝb�!�����A@8qr�M9n��m\�E�d#��QdB^��bm����6��cvVw5,���o�6��U/F�K4��g��G;�۵��{;q���=gv��;V��w������=EtJJb� <�]�`�>wq�;kss�;VV��l���U� ��;=��4���y:.y�n�Չ��m]�Bmƿ>��~�H�7"2@g񳒨C�?���g�~'U��w3U[�Þ��@A??{=v�����7N��^<���r�[�wkQ����g��#������r����'�VFB��Q$Z����YVH>7�蟉=g��U�ˬ)v<��@w���$�W�蟺���q��	�Wf������/� $�wz����(���B3�y�J�U�	�뻰OO"�К��	rAB,�t	�{V��u태;Zs��$un]�����H�-�پ��������_"0��1+�L��Xg��1���㘊�Ij�R��$v;8��3��rHԏ�S���A�yn�$���5�Y���Y0;�3��U�X$r��@�VJ�(ӑ 0v��
����ׯ��s
��~�<wn��{��#֟
o�AN��m�O5]�')Q���kt�,[����[˺�z����W��"G~�?�#���O����v��yZl�-#~R_����#�x�M�ۀ��W�	'�y��"EV���V����I�������Aޅ��E��P3z�|곳2�a������k�_C��X�̞��8߁1_����r7�Ȋp$L�Xo�'���̆r�٥%�5��J��ǹ�� oc�Hy��}�BV�!�r����~�)�P���ֱ����k�[������EG�$F'/p�cB�$���:$su�A�g���m%�ޱ�o�wS�~$�=,{��'�F�u���A�T}�x�/	W���v>�D�C��]�A}�M�<��r��$j���p�\h��{���}��H+��@�k��#���W��^��������M{i� �ؕEL�����!W�ꇚ��e�~��ø}��%�͇��i�DQ��[	��5<b��/�{9�ߞ����4x�s��^�L�q>�n1�=����Ny�wݔ��)ӾS�.�f��X{g6?L�=���%x��4�8��H��ah�F0�R4r�B���v�%2��Nv��}�G�={��V�g����:�p��ُHd=�O��:;F<��ξFm[���߷�W��pN���s����}�%93��_s~�pU��nMo�=�z�>�l׽��Y�R:����!�����*���s7v;�UVr
�h�y��#a�E=��ϰ��]��C�f� G�~���wsKf�r��s�?!�5��f�}�X3ҁ��C�!�2��m��(��o��b{�x���R���,��h�cև��A�ƯM�-��o�x��|Z�x�������d����ݫ˵C2n5�m�&���2�o��d�ǳƏ_Y��s������O�\�m���|��Z���)}�~z'�}����M�w��"�V�[nl�(����f-��w�E���=G�*�sx���=�/^!�(�T]�{��4�MO{O{-�5�Q��zp���_w��C��1���+�xlJ�v���c�.n������Vq��fP�	������V.{W�J���e�t%�
����0e�~Sv�'{ @D���3��]�U{���j����R,X�B�
	�a@�Q�f]ۚ���h��	�$Rk-ĸeLI��u��Q\�#��r��G��D[����9r�׻��o5�cC˙5�ݛr�4X��W#��c�h��d���]9�sn͏��]}��s�d�r���0�~7�h�{�|���u��F�建���E��;d�\5��gݾyU��1�b�wqXkF2�^�Y*1���n]5�F�8W���k�ʍ��)��;����w\����-����:��S�(�������7�u��/.���.���n3`��qr ���\���s��ȚJ�C�(5�]6>s�b���5~+�^~77��wWw�\�4�[��TH")�0����o�$�gP`�_nz��C�m�#p��.�r�c�0k�L���$�*�dHw��A#Uu����^��w�u���	�����4� Rq�% ��]n��Z#��f�-z�'�NR�K�o�X<k�����{;;]��e�r��v�����]�]l�ݺn�؆�^ݰv�:2�4c��7��D��
H��2-����b�$�_�����U� �-� �w��H�QQ�
(L�#׺�I��׎��2!�w��$9W[�Iә\ۇ�����Ȃ��k%8����Ƀ��� ?�X�������M]��!�w�� ��W[�N�:�#aF��@��Pv�:�A'r��,�H�D�[ݖ��q�A����$6��k�� ,#ȵ���;��X;��u�q�Ϸ�`�b	ш���9����1
'"]�f�}"���������y��Q����W�ŽA�w\�䵇�LwyvH$b�n��{�z�:o�|�}]�X�ax§D7�v�{/o������̔��/aV]�s=�cPb�W��?	#B�0K��8�L���'�m� �;���#{��
��;��fn��$��m�$uy@�%$W`ɯ��~]�y�I*��$��6�I�k��dλuy�.���f608�@d�S^�tO�v��D�ﻜrf`$�)����Ԍ�KY)��)�96�r��^ ��u�@4z����oN4H%��מ��c~Q[ԏ�嗮�'��7L��Q���͎�A ��z�y]�<�V�N�$/�w��ĂO{��@�{}vgb��I��*���\�2����;2Otg�5�;�s�b���C�fz�1j��d��qC���M�`sT��<��B��}���o��V���� J�@:K��F[����g��;�|��R􋶲�
l�&}��tm�u���d�ipq�g��A�^^�vt�Ы���KS�V��M��=�׌(��ז�u���9�6��!�!ӣ�'
��]-���.M�\j�ܾL|`ݭ�Dpc�g�kn8�ݚ�wYS�:�fa��Ө�rdK���Am�8���y�l&y�7.�f�z;��O�n�!�g��1�n�Nzz�L$Gյ* 4�;����$0���y_��F�R �_{}v	<����eݏ^�tH#�R7 �H���� pJ5Ӳ���sx���l�s�`�[��c����� ��Oz�g�o}��n�@�%$WfN|E�s��=N��U)w��	w��{n�;�cc�A$H�|׺�С������O�U=4$�{��c�yN�T9)"�*t,��}H�.�d�#�(�v1���I�1Yut�xf��TOć��]���_�s�H�Y+�K�BR�n��24k=n�V�9�TVA���M[���%�[����
0����甥_K�w��?j�����|�n�V��_e�_�����28����_�$߼s���LT�\��8:�23��{�'������z��ԅ0M�o4��P}���$����X�}q5b���.A�~Ө��j��$�^U�����=꣡���2I�"((#$H�l�Ւ��	�8��Hy��d�/��-`V#��K
H��2-��&������\s� Y�Y��G'�	=kyS�^�s�AS������,_������F �1_���{V�|Ҫ��x��i#;s�d'�ǭoS��ʮ���;����!�gF1\7��|s=�ts�5���7O��K������O��Y)��9p>��$ix��A;oyQ��V8A������m�rz��꣬��4a�C�9��=�v��<��f��$�O$���A���]}�h�b��=��O��m�� .�j�!?��B�5^⼛w��]x�c�s��'O,�Qw�}�"}.Բ�FM/ok��h�FïW���Uo�*��f�\�����5,�����SZa��JR�u�5�����BA'mwS#^�H�
��k��zJ�Wf�¢��h�Ǽ�$���	z��R����Y�=�=�^��؍Fb,)"�uA ��˽=w�������?��S��^��k׊`��ƈaH_�0��ۭ��WS��佷:���7F'5E��I��]#����3�1��w��F�ͦ~$����'Iν���^K<� �{��������#�>��ݟ�����}��!�V,$H�}�� ���n�b�*wR��R�ZW���e��c
H�ܪ��]��OƬc��Y�Q�څu��%�nB���w}o��]n{3�ݣ
jmI��~��`9�4��۷�L�?Z���駗�x3#�ݧFܗ�q��cfa2�<�d�w��jy{�|��O�mkN�D�+��/_�lx�RS��$�R�2��R
$�)@�Om�'�q�6�sn����*$������|G�ywqO���i�T�*��H,��B�	\����o���O�p�ߥT"%V������Į�QdU��0~*�����$�o�#�c���n{�ϻ�  yyB��Y���bC"
�H���u���g��Eν�d�o������ =D)	��bf�)A�������k'�O�"��W�[}O����U�� �|a?j��C�RP���*���]��ǋ��P�O�^ߪ���o'�4߻r��Yޙ^{�&N���%�rD��4�W{o�|Io:�4cem�U��^�g�Y y�3�~#M��I��)�.��g���{H��o�d:������*�L]EԷ�N��lo��q��ѿ����G��G���|Uc{�]��	z�|�L�{cz1��<^�!����"K]m�}%������\q�)����`�n�8ю���۶�83���l�3���'nwc�X���k������0�N�"u��g3��{y:���ǎQ<�W�m��\�t:�b�A1g:��9�q�<;c����G����7/[���h����\.�;��t4�n�:����>�'��G������ n]q�'1���;:K��67np��܃rp�.�W���߷�U�i#���?F�U���L����?|�$�9_�ѳ���\7��%��z��H���GY��N�eI�^v	�7Ǭu�
9;o�d�N7�� �s�����&�}/w��x���~��!q
��;�_BO�窷`���K�ǚ�> ����!�oA����Gw�=7׼�����z�� R� $�����Ou^���Qc�w�-�������	����)(dFA=*���=�}��>3����	#�s�@~-w���fm3���=��HC�*��!Z���o7 ��ρ�\'-N���6�m#��Ks�����'i���ߌ'�Mި	?wU�����LuY�[�	$7��v�HW��������d�M�|i=�k��4��ǳ}����y]Q�[��^�V;R`�vQ��F���q����l�c�cK6�vů�	G�^�s8�_�4~�A ���]A�ڰE]�_����0]׾��q�n�lH�e�نwT��W���	���q�GU_��F{��W�`�x���10�q
}�6����;${�Psj���~$oH9M�J��K^�VH�����v#�($���^�ş���{`��M˞��zg�O��*����n{�_��wOl�KEg����u�*+�l��Ǧ㈰/��������:ۍ/�o��"8�.�����Q���e{j�$����~'է`��D�T(G���/�.am��M��Yb�	캫���\�H��e{��?o8DX|�rcl��|7��B��"������v����0��PX��K���.1악5I���{/��c�����_��9,�|3#���T��h���t&?I�E�F;�w��N�U�<�A��8��z�����_�ɑ�u�4�2ᅶu$d�������B�c��� .�2 	$g8D��v׻��+G���Y���h����$�՛N�<;�sԯ��Oww��$�� ����P~�CMbǖ�OH�mH�$��D�khۨ�����DKl��
OMuЖ(ݝ�I'���p<�ĔH����u`��A$���ʁ#�����y傺������ ���6��2(Jb*���T��ȱ��s���n��	��~}H|=D�E������t]7{�G1����3 M���n\���� |*�V�]İz��ē�>��?�>4ꢩ41������nU;c�P$���I$z�0� �꽾�L��_����z�#�SYH������џ�i���X!���~�T�a6�{�:�^�w݈���ʮ����zF�̳q3-ڟp�d�^ԭ���M8�N}_"O���.��ٽ�ov2w2A�^R|Ou{n��[}�=���BH��'�;���k�l�\]]C�w����72{U�7����e�(KF���A�Ǵ� �W�Ƴ�i�X��o�o��k���DP��8�ĔH��}���D��?�F�4I?�ߧG���dn�y#�~�L���>$�y4�(H�-����T �W�łz��g�6qC�E潯�$�W�ōcեϤ0�e�R��=]�&X���O~�� �WH 㿉��v}GG�P3��~�����E,	��ߤ�(��`f�������>mN"��u�?��~y]��Zw�i7��4U�{W��)�c��OuNk�Eoi|��bZ_���n�#<�m�^��g�����_��z离C�n�����x�R�.z�}��t{56�BcFcY�W�6���\�a��h�[��a�v� ^��wk����<���p�Zb��>jO�/4�[*h�?!sp[�Ƥ�{�w��j���Vu��9Kϟv�����_�s}u��̞�C8����?/j|1y�"��m�7�����k�ִ�.��5?+���fw-8�>�[�r��oZw=��4)y�۽�_l����6-��H��f��n�1��kv2�ԙ��F�שf���瓞��q�s˾@]�[��S�	n�OwL���ϭ��z
g�Rm�Zq����
S~&OI�uu���8�ޯx{-�<�ʾ��O�����߽1�]�����-�^/p�.M��oxx7*�%7?_ ��9�Է��i/Y�QѨ�:�o�W��kx�ln��^��I	��ۧ��qlLZi�s|��ze\����T�/YxA�-
���/A/��{7wL�e=�V**�i��x�6�/��w�jؤV��;����,o}��mԲ���ˑUX�\=���k�xV�
�,��J��{��F���2�b^B��<���|ua��SN��5%r�Wng��y�N��-x�o\[~��
���y��/�	׮J�~I�V���g	��z]��v%��@y|읎�Ą�NCqL��I]�*����WL�p������3��'��.ˎ����=���E�}����z2ʱ�<���]c8g�|�BjH�?:����,l/-ٮW/<���߮�_;�\���Q�q�&���w��U�����}ۛo�r1�/������s�Y���5���o7)2��sA�F�nX���
9#�KҒ6ܧ���ܷ+�%��u����y�r�n�λ`�����[�u���r��o+�8y�WM����W�#�nh<�|��G9PE湩.\�G�j��wh�F����-����+�p۟*�ǚ�y]6F��;����-r�v�cQ6��ъ6���^Y6�ѫͯ,Z��_-�W�ulEy]�.G5�U��9\ܡ�pؑ�d�4T���+�5���r���ܢ��6��^m�ܨ�Z7�s[ϕ����9\�ܫ�^V��7G0��M0˘�d�Y+���\�Ϛ[�Xm�+t簽��/Wj�y:g���h��ۧp�.�V3�d�v��\�<ڧ�2k�Yˎ�q�����7��ln-۵��*8�Þ��qݖ�c�l�p�m�h�l�2�.��� �'=���ҷ���'lXH-f��F�;����u�`�v�-���dƸ���I���ʡ�[m���y�5���S.���Ɍ
��3�+s���[����Ǟ���e{uΣ�l�WF=�gu����:�\�wGc��v۳�mM�7�w���%1��1���3���y���n1]ٲu��rW+7ŉ[&��:�w+�ɂ� \���u��,�%�Ж7dg�Wi���L��֋y%�u��k���"��:�Q����\x�ݎ1�y��ۏnywn�.�^�l�A��eoks$q��b��m۷i�(�i��@r@��:�!��z�lg���'X�9�ipE�.�{t�y5������6c�/d��S/k�j�粗A�K1��u-c˲��wV]���V���ήc����s����[qf�s��d7)<�ʹU����ۨ�xCaT�7iH �ȼ�6�u�ʲ]{m���B�����jy��kŴm�M�������׵�N�3��^�g&�u��4�Z6�;1�z�=�u�V$N�8���tr���:�oT�ls�ꭌ�@k������[���h�b��Kv{n��A�M�к9�y�V���w#g�hۇ�.z�6�tPl�z���/XÛ�y*��y����=��^��؞���۠34pcg��J�r�ֵnݞ�n[�{;-�kv�M�9�f�9�Ѯ��+]�79���[{Q\��Cb��K��}�î���s����s�-m��&�5s�gm��g�7���N1�͓�<n[��[���U�m3&���[����a�[j7"��]g�(���:Kg�b͛�=�n��s�5�P�d��[�ܙ�F�n�s�i�����/�̮��n۶�R�3q��\f�P���gm�c���KnI1خN��Ar�\��]�<��}]�lq��k�<�1�
�����l�8KnL]
Y������.��gG�e��[��=,��.�壱���#ugn���6�٠;D�n�u�!��"�y���Ȃs��y�@]2[i0���sk5��!8��;��[V��ru��G�<q�]p����i��ۆ����N��wZ,��V���vݳaB�2�Tm�[M�iQ�ȋk#��Ç~nm�����'�}~˰I��O);s	��t���l_U��@bP���=?�X����㓡>˼i����e�.�j� �Oo�3H�Ү���~�0h��$��Gv{��A ��_@|A[��۸��8� {יv$���_^&�;&Kf*}>���b�a������I�]5���A���l��Z��ח�y��>��M�zn��>ߗ=C�_��y�sۗ��>z	�oPG�ǏI�o	ǻ
1�Ȱs)�L<ݸ��҇gk��9����Ӵ�n7GQ���c�L(b9�\�]�㳝A���|	�g�G4/wnvg���$�]9��i�7�6Ԇ�5�/��V_e��(G�l���x�q�'�6χ�~%H����}шo��$㯷��a�ܻ�\���8a��ڥl�@�z�Kw\,�	�kI����x�|5_Яh,u�Ty��;w[�B\e8�;�x	$�Ǵ�^>��0�Y�x���X'�t��@�~6��|��\0cGR$����]V|�Z�5�=@�x���$�o'G�{krLsr���_���i<���Չ�N�D���� ;�� �zg��҃Α�yfs�>|��_l�m_��0���\ݵ�d"P�(�ͨ#0G,Aٰʗf��޵�h'>��Ҧ(�'!dM|���2�M���~�@I��h I;�c<���9g�Y	>�D���� ����E&ʁF#�G�gX�z;2�
*��r췏1��D�ӽ�[��[ִ�W�<��}F�N7	m�x��k�A ��e�`�<m�)a��������[s�5��CW�3�5�(�*1J��Î8�8��k��z;-��g�,���yo���8�����H�ٗd��m���*2�b�����u�N-���n���=�X;��l�ڷ=5ﲛ�G�/�Df#!�K��ί_�el�r�m�ÝyEy�_WN���~=�ҁ�ˬݡ��ľ����/Llܷ�z�1ţ�M].�4⣥M���]�F[�{�퀉h��'9��;, 	��WJ("k��f]����732���5�|Æ �m]���P'��}x�zJ�#���x��ʰA��
8$�Cֵ	I�錇qi��r�@e];n�?{���$��>�$��7��U,��ܫ �F�t�HXO�Xe�)�!��އڪ�`<�eq��%��X�$��	�kyf�t(qք�ye;k2���n/;��}�w���7���* �w��E���������g�3y��z�³�<��Τ�c>-�8N���Z�y=�m���*2�b�+s�ֳh7lՠ���O�$�](I���]�qs�híQJ�")e�eR{�C���`;i��6����L��Uף��ޫ�~w���$�I3��mz�����$�H���|N�˳w0�][��f݂~$et�Oǯ�턙`��7���HW�z��>[Z�A����r�t��� ����J��.h�H�@#�gM�"�ͼ����g���g��Uk���w�$j��Dm��M��EA$N0������\����I4o|�	�>�h�C�̿F����{�=���{�k�1Ax�J4"��Ԇ��h"	������\gfU{�ޱ�\Oئ���ה��ʰkGb��5^�%l1Ҫ�|�U��k}<�zn|����iR�I��\
��hy�˓7D�9���1m��xc��~' 5�U�m�m���?�!Ӻ6�j�6����׾c��I�TE���<@���v�w��0���0�v�V���R�±�c�����s������17������,vCr�lv�ݺktir��X�=����3rr��cr�S�v���Ɛ������-���q�W.�b4�m
k��f�7Z��*�ptA)���#�p��w��s��َu���	��o9�([sT�̦S��j��x3��\�}��5���b"�ٜ��z&���mC�q�'�O5�H/��vs����f����P�k�A�,�$@�2$���U��h���ת�Ͻ��v$�N��T	'�{.�-��W�ws�S��vu�焃Y���BL�S���J�~$��m�d
�-�~�e�+��|��H��?�N�]�5�-0F�p6J����|lh��TS�Hm{�0N=�U��Ӟ��y��I��^�A=��PI�) 2�ڙ�`�����s��z��;1��k���{.�$j�΍��[��:v����)�5Ҹ���9�w�u�l&�ߴ|��E��l��S�����B�QTHJ��7�A ��e�˧1J���EO@v�Ry�����m�$(���$����f^e���k��ֲ�+g��O�̯{%�h�1<޹��\5#��
Ӷy��{�+��8��_�{�1��}��CZ�Kv�'}� �y����Oܟs�A�6V`5��Y�8�-@�2I&}d��o{q��rމ[������F���k����I��JqP7��z����^�S�O��αd���: �U����n�_Uɷ���ޭ�'��EU���#A��7�O�{_OH+�������e|H��˲I��]|I
�u1֦�����%i���nT���X�̛v�[&ٻp%���h9����?����}��]ih9 3��\�x��D�I?+}ʈ����X}��t4�O9�g�;r6"&ӂ��0_�*����Y�y>�@�B��_0~&���._cw�ʛ���o�F�$��:$��{h2Iܼ"��$te��{�T�*����J��]�Rݥ����	��o�[�7���ˑ �����Xּ�����ٖQ�HV����A�ץ�Ē<��A%yoS���#�)�U�r��,�G�ݩ�zUY'��tI?����$��ox-�5�������&��/��L�S���A��}^�	�G��-z��$
՛_?�WmX=��w���kP��ʚh�c��֯9"�*��f|�7��f�F����Q:8Re��Lp4�J�j�!Zޯ���������&�(N���^���SӤ�!JG�Fw����n�ٶ%�0Ύ��~�r����۲~,?fzd��W[�B��ܑ3�6�`ȳk�A �����$L�nu��'����:����`� �/e0~���v���l(˒A_5}�M��B� �X�n�r�I�;��~<_see�5ʷ��{����Z��´�H�6�É��l�7%7��)F����\����]l�*�Y�%�y^�,��ȓ�,��.Z|�[`�-K����udiHd���۱d���;�z�Ӎy�`�^�//6�O'���Ş��f�����$��&V�թ��#$I�B\���F��E���V�s�+�����w�\���Jy甪�O���n�:�s��}�βiy;b��ԅ2g���n1!��o��+�?��L�OfQ��7�&��'�};�v<�ssiU���#)����
��2B�����;�O��b����{qR�l�i��$��>�+��Ż-G%�\eż}g���;�]�̽� ��#��t �m���ݨ7�yݗ`��m�/��08ゃW��~Z�PyOʭ�k�x�zM�4��D�H6�r?�O�L�GSJ��{�*����ܜ0���޷�J}:�G'�����U^��o[ݣ��9�ZkC�!x�z�_q��d���ww�F���Ga�v�]�]RF5�t�#Ś��n�;r��� 6WXn�ܬvۭ�<\�<�1�`���`�;�5��
;�`�� b�ۜ�;u�-8Kq�9A�x�-�e3� �5����<�y�m�X����q��X#X�J��'�zSgZ��!����3���\����xf��7���pb�Xz��콇���m�3&!�j��u�v-�"�ٌ��uӵn�j��Ӥ�gaJ'E�hԔ�6�2I�3��b���]|A�����G����|�/����u�$�kG��F�cԦ_­��>�_֫Ϋ��'��t	�mgS�u��뺱N��&Ug�%d܂H�r"��]���LQ �[�?�#�w�Ύ�3�A<�k���/:�+`�d�$��]�3y���|���A���_�?i�:$��e�4r��/�i<�@����5l��pXMn�$�s��+��|�4I�َ�?N� ������l�j���=��Q9D���"YK�]Ut"mutb����.��3����Z5����>�y�ɴ�>�{��������x�{ͅ�ta�{X#W�|H�~y_.�s�:�:R	$���A�`H��w�/6�JA�܄y�'��o�W�&w�-T�8�;'�s�������UB_���f��#����w@�A�v��(�횪|I$��Ɓ?���]�	=~ܡ�`yT�=�D�k��bBYh�������{hY�闸�d
��S=�i?z������-l�A$L�!l"��/z����r�����'3�+�A ���ł~�ӝ���{��5v�A��&HBN8T��tλ$��ӝ�3��jc�3M풍I��v?j�΀&,�/8�*�-��?�����s����1��]�q��ҝ��=;z�,���/�Qz�N2�i(7����ė}���.���]���^Y�O��l{H^����+x"&�8঻��y�t���e^[�|�%���,=9����v�p�KVU��k�Dz��:�qD�G.���]�$95� ���\4i�E*�B��:Y�5Q�/��Ou����/#�h�W��g*o�Z�]�3�oqz�>U_<�a�jݪܲ�pݒn�p�����4o�J�R��G���e�a��Ml�=HmK�u�&(U����Ӯ��#Yl�B#��|���Ͳ?����t��b��{t��g��3}�S�M���Nw��7e�����h%���U�g�|4�4�;֗l�۷ �s��1$���`ynyR�eq�m4|��&�H̢+��
�)ķ�ʡ���$6�V�B���޹\^˛�sD�iP��1�2�{�S�́V:$�^�ye>�I������FR��g��|N*C����;�,�]�b�z�`�Wj>��4݆úl�\ć��fOq�8����{�|5�L��?o�76��8�5ը�e�%��.�|��yJc�$��of;�[���8���NT�����їy"���6��ߐ���QbJ:=F�����>����I�]��潍��T���[�ز�{]��<*�\G���$c��85w���
G �Fv2c]�w|�b]c���^��š�'���a��{��i^�z����i>�ޞy`ۅۣ��C���3����WVW�M�D���-w���WE�������s��/w�x�E�K�l�Y���&v{�(��\�ζ{_�����7=��]JM1k�v�Y�;_h�q-�^x��/�r��E.C/!�Y5S�.[:��7�sɄrg�U;���M�_f��Wr㛨��KAX�ʑ�L2�aq����o����oZ�J�pYpE� ��ʍs�\��5{�׻\�k��-ck�ܾo,xh���u^\�W��둨9��v�k������;٧u���o��5�U�p�^W�|�W��W#]9c`�F7}ה[��,\��1nsE|���Kr��u�x��nV弭�������+�u�s\��wj�&/-�+��.�ҋ���d�+�\^r�wQE��wA#���W8\��T��%I�v��׺���Z���s�KynN�+I|��|�7+�ܹ1����S��*9����]w%s�4W9���r�����-���^]�������z�{�"�i�b�U��sbM͓Ep�[��+����|I#�B(�CJa�A/��vA�ӟӗ����q��GX��S�Y�� �K�A �]5���H7��5���b��uؠA޺���]3��"&8c��^�1D�}�� �:�[���[�da�΁�{RoX����pq��9(HnL�؎y�S	 �q�X�}]wZI��I8�i͋WϿ���d�%#H�fOe>;9�����>�)5Wx�{�ϗ��v	OMt	
Y�m���PXo_8������Ї���$���:�m����]���[q���d��'���Q(ZbpW�_s�H��#�xxԙs7G��*���|I8�s�A&޾����I��'�9]�>v!Ӏ�x��@�A��	�{o����m�q�䞺k��ߖ�"Tq*����߽�}�������{%R0E��Y��=n/	���9���o/�g��\�H������\l�'ņxx�UB>"w��w[��+�E�+�@"�N�3{�V��7�j��&�����Q�$��;����������1�s�y����q����<��~��/U�RP������H>;5�$���;¶���~��΁ �}�2��i2Sq��P3�u����t�:����c���?g9��$�7��/㕷��Z3�fk��6E�ǔ$�� �1�jwC������@7Z����p�ˇ��c���A쏨 I��۲G/+x�P��.5 ������b$<髹cjb��\���D��݂A#��7Y<|�d��}K���7nH�r�N�Ϭ�8��G�yV�OQ/�0�$��]�	�s�gyV�ƬuxU>5�*�����[%���9.��z���|K,�:`��:��V��}Q^��]9�����������k���S���_��'@�ߏ�7m�m0h����P�d�0��^���5p�p#��7�
�6:�@=�����b��ٶ��q��xvۤ�Gn�v���`� ck�S�7l<�\��;�l��A�|vr�F�n{:��5۰-�k�����s�H��?�����x��^�Mc��y��]��]v�k�`�Rn<��LCoC�'Qvv�{c�ɇ������ޭ�Q�x��k�ٽ.�d��DN�5��Ͷ��0z#<�4���>�� ��6��"Hw��,�A#S�c�Ӕ2'��ڒ��`���M�7��1�v�m�h�]+���7�D�{��m�����5����?H~�m� �}΁%��m��<_�{)� �+��Sq��P3&m����_I���1�w=�x���]�I#��u�dXqe$�`@*�N�S���s]q�oמ��r{ξ'�@7��������t�/���>^V�D�i�dAI_s�A;��#��5�|<�UذH�}Ή��o_PA�f���ePI�0�a��C�#��MѺ��N�62sz�a�u���_9=`�I�Tr4ԙ��}w��4��� �o������*���e����O^��p��D�k��!� Q�;���9@.�����7����9�*������[��"�Lt�(ڕ����g �.��z�YR����&�v�e��u7}I��{!u~� ��󘯉޾���13�M�w������h$,��D��.&���~$�����	'��j�<�a ���: �z��G�%�n@Ӏ���@���fzP�<H6rk�I?��k�ON�є�;�҆�ھ�C�&�h��Y$��Vc���>����7='������*'�=���������th��@/���DȤ�,�v�˞��㱪0���Wv�0����v��8�^�]�F�-�[A�;}��$�P@�:��vv�0+�n�7|�Fd}Au�Xq&�Q��RU��w��Η�|���x	�a���eX$�n�R�{<�Ex�;f3	��΍|O��{�B�#��18S�z��=�R�����,S��&�����Y���ג�-|��~�;D�k����A9��Q��3
��G6f�bI쏩H��e�[5�J���u`w���_���~$��)I�����I�rUZ'V��o?pDpq.�r�P�gX�O�ܧ*%�g�kr���.Ϟ�f��@��=�`�O��r�r�*�s�%��S�NnZ�\E��y�p��
��{k���#�[k^�l<��T��\=����7���.��X?;��_�X�%l����/��{.��j�j8Ɍ@ؒ
|�ʈ�9���~�N�9��A?<�u� ���*��1:��t����F�ө7
�F��A��H �~�X���-����7ڹ����ۿ�yNT	5Ǚz�3�����V9�HJ���n� ��s�~"��Ы3��N*{�њ<I��/>�r��^qFQ��M�.f�t);;P��;��'�{5��ԓ�vr8��y�s)��z��]�sK��Y��_U�J���Ha*�e݁�~�@�|��^�v��W��ݎr��&�ޯ�_��owG���%(�)2�M���l�m��7qڜ��K
6�֕������
�������Ow���ܧ*��H���C2H&��:M�I {\�D�ijJ�q�j3v�yQ�q�{�|��~	#1�TH$k:��Oa,��y5�ě���[aH�"����q|�l�2�$�}���6��/ޛv4��g: �k:�=@�I��q�ԗ`������a7�tOĂV=�+�ӯ(fq�b�f���.�b�Y���C!)� �)T�����m٩���Nn�d����s߿~s���i�8yb���I��~���xT�.�hf
���.�h{!g/��u;;��@�u߶�J�<�wgf'�%���_�GF���]9�P>�g��<u81��v�qg�L>IwGa�`xvWål<�4m��om�3��Q�s�Kr#�;Y�5�ƌ�mV������5�N�湝�y(G7m������[Uـ�{�Ӻ��zݹ�4�n:��ė���
�=j.r���t��d<Ho��y����uԹ�%w5��n�7A�uqi�{s�l���tqۉ�]�ָ���)�����k����!v�ocj�/-�X��m�ci�l� ݌5�5��ەU��QKs}��UZH�}�{��$��_2H$oU��7/�����*��}���d�H$�/m~t�D�'$�7�y׶��g_�Lv%�M�I!y�*��F�^]�Tu��!�)���,���
�XX����i<������X7M�^u�JŻL��yw�<ig��&$�.�E3�J�J�'�E�A�I꾻${�C���/�v�"�{U}��ԛ�GFIvݻ� ��6��9:g���Oi
���u^XϦ�T����˭�η�P�	���r�������\㳆-n@+m���h`�����_�5	��	m�7��"I�U�X$�����~����OP�H���|�80�9뿊��D�ID˫��H�c���d�����?~/��x�:��dr�������j%ę�G��F�w�nxg�û}��cumg<�H��*���=�ド22Do�I�٫�a��e]:@A��N�H1�p/�o_�"�>���p&�2���I�҉�S�ެSq/_�@'�/n�'�Aޝ(#�7Չ�mK#�z���[����e�]�	�(�%o�g��f%FA>'�ꮱcW�x9��I��t�~��yATr��>1K�2�A�(	������f�W��YO{���$bD���ĽLh�1'����a�v��.��.�r�R�=���$ي(�nOwǽ�ud�Gd�_�%o�8��
r��n��땷d�t�@�\u�bF&8n��thU����{������~�(�?x�����S[t,����Bُ�B�iD˻;�T �_`�={d?�ɓr�Ӌ�$8��'V[�{�G~�N���A��'���4yE�����3=���v뾜����F)��^\T����NOz�S�#뢉��}�jٮ�!^>�N����REn+��=�%�h�{n�T�t��I��醉$t��KB�plz;-z����<($�%��5�澯�?�yF�M�}�(�Vs�(��u��"�m���q.�f�)a$u�[@�����1m���=��9%��״�Őz��4g7������\u�	 �^� �H+q�|�ēӯ,gYI�yg� �H�r���Ϩ#�ecĘp���b���#3ϻ�Gf��lA�0���ӯ.� ��=��$��MW7�H�m���:�A ���_����he��zxI[����:���Bٯ��L�˻���w
V�3��<O��?R��z��H�tѿ+��:�P?{�+z���V-������S�Y�B9M��p�����\>�ʆ���xk'�ݰ���d�t���?	Y~q���!�}�4T�0���j{��$�t�.P������?�=4	�son���t���{=�����}^4Uӱq�pg�x�4�u"��ڶ,�`s�<�^<��E�\�3/�B�%.7��yAI�חd	�t���]UZ�.�>�tE��^]�O�U����0�����0�b�Q9���3j �ON��$ޝ Z�+ݕ��[�D]Y^xS���,VmVY�Gl�D���<�z���>8?�ח���҈��AF"�	�_��K��N�.�
���?A͛|B�|������5���{k��'ՄH$6"����%{_PZ=}�o]��D������d�I?�o>�$ I?�H@���$ I?�H@�d	!I�@�$��H@�����m�ڵU����ֵ�z�։'� IO���$��H@�}H@�d	!I���$�XB����$��H@��	!I�`IO�H@�t	!I���e5���\�9�� ?�s2}p"����
�%(��)JP�PJ	" (Q!I	H�P%
	P4�I%P $( �$�� ncHD�ѭ+6�Y%M��B٢@�Lʛj��Vb����I)6�HT��Ji�����m��Z�5M4��d��$���Rӷ�                                    �         H�__Ay��g����(]�/A��7� �������)s=�j�-u�\���z{d/ ��Mͮ֠��#]mSУJ4h]� @V��l(��y����x �5��pW���G�d�1���yj�g�^ ��o�w�g�E�ם�Vۓ�^R��d���@         ���\ϻ{d���f�<[�k��姫a�x ק��^���z�[c���m�ΏfK� op�ox}9O|�9_Ԧ�m���|   ���}V���� �}� }�������s����pϬ��j��� ���\�����=�(I�7/�g�3{K푕k)EZ��           �X��o�o��ϋG}���9׬������ �^����o}��|�K��騇��W� ����L�ż��Y�J����G� s���t0\�ZTOx �ձ��I]�;�ݺ�\��q�/ ����}��P����0�������J��/�6�*�՜  �        :(}�3���W0���C�=���Ξ� � � �������^�^`:x��g@�g�G�:P^� <� X��� :<�ty ��lccn   �>�� 8��h�z� 8:�/�{�t�^���Һ�;�y���m� �j$����[���8�H�g��Km���  �        ��2�N��i�*���ǐ w\  �x�krw�����������À��w1����y��<]��K1Z|  9��ruX��hw�x �{m�'^�OZx���=/6���۞A�<�^ ��7��wMk���:�-��[Ǵ����T��ҥ)   E?!�)J@  S�"R�4��ت�m%)   5Oځ2�J�40�I1J�� f'���?����f����'C6�.��C}��r���/]I	M<���$ I4 �	!I���$��$$ I! ����o�������ޮ������u�?UNΜ�6��ȔKNZ�2
�i;Y-^J��ژ�xX� �f@�.�}���7D7��W��e�������c&���E�ft�,Y�4����uXʰd寷.n��HNKG�2a�<1a�B�m�N�r:زͻ�z����fC���K�&�B+.��t�� �u�b`X�������%��章:1�"ƛ��K�K��;e��]1���٫h�qhJlgZtf�X,�
�	�3CAF��P�1=��8����֥m��V
1�#{����b����d##9����Ƒu�K�!ٝl�3Z{���j0-�dj2����I:I���L˃]0�sM=����Ј��-t�08(w�1��
�ͳ�V�Z�Ӵ���d��z�PF Y��뽑u��g*_�,��ۤN����n��L�N�\�WV���kڇ<�p^a����$�	��𙏆r�<U+�7-gn��4������9B%�H��e;��e�/(	�&�p�L3u���&�,h�;q>Og��m��W"h���pH��((
)2����ϐM:�P�32�۬N��[����"��9&����J9�l�-�q�<D��5�v�9���&c�1�M�����1��og�w�I�f�5r�׍>�;�9s�k ��g5�S%����Q�w7V�V����d \�0��z�;�!�gdz7Yϩx�%,JxK�ԍ��k�u�p/)Q�MCGzٻ	���5:.� �<g8;����*ᇧѰ�;�h���|Kz���]���5��.�{۔Ǘi�#�kE���"�8�A2Y�k_'�"	47C3a {��#Qo��W�[���o�50P�b��`�p)����9�T�`ٴ����;k]Y��?y'��}3{
Bj(c�02p���幌��n!d�:�aYn�gg�Y�ګnݹ�@ىe�!\�w%sF���øzc;l���I8���n	�-��j�����X)F�����[�W����׿�kc�tP��QPMZh��$ D���d$��cz��b�nq�aܮE6<�X#��ێs*V,��_\gs�v7���	ͺ��na#u�`�#a��G�pI3�5L+�y�F�����Աt����gb�n9�ɩ�Ή���W{R��p0��gQgR��/z��2ckbT�Gh�g� �����ݹ��m�'��l�<�
�6b�d��vt]��npK[d������-�`�~#&Y��j�hn���r�XO��!������;b��u+�h;�Q��J��1�US�u���任�r9��7����_�6����S�\r�e�.J�d׃�Y�`��뀧�S�Im����F@�;I�8n��'J��$ފ73o_�<nn����\里���f��Jm�E&n`���LQK]8�1�w�b���l��p�7��/[L��C.��z�UcL50W�%V:�:�!�UB���a�s���gV��
g��(}��X�v�a�nf�4�{�	�]�K�q�)P�gCʍ�e��[����2mް��hXD#xE�NrX�S^�ʙ���ܗ�G�Z4�ݛ���#fL�,�^Mm4I���.��%j��6�t�IS���sn�2�9�Y1�a��I�E�M]>Jc,C�ٹ�v�ݭ���H���@�T�5�,�3�n�����^�:w�;EO�U�>+OhX�cB�\���/�(a�ZY{D����.��s
=�n�f�
OC��H���c'�#����tk� b��ҋ��*,ۤ�@��%ۑ�YAs�4!#K
,2���s���Ϭ��[q�%MW�t�jA$nnY�B�5�ۙ6<pA%�.�w1K�I�8���a�\�����J�9��:8w�"�n�ܔ��y7DE޿(�".���`����g�9�c��L��yt���*̟ ����r�98�%���.��j�@��Sq�ۆs�`�;j�/������BeLc`3)jK�^��'1#4�r�ܽ*"hΑ����2ʀDܐ.d�N���fǢ@[3U�<�s��`o䑽cC5�g7c�34��w��%sf�h�,)�7��J*����H�I�|�w.M�[\�ˁڽ������|�Cs�ne�̚IT t[�Ҧ�u}.���v����N���x1ꤛr�^�3 =0�9�VW�to<Y}���֖<#MLǇ5�����N
����)��ؘ��ә�"�"#�}�YE�[�?��2�e��l���44�Mcx�`��L��!��J�^>��|{	�m�4�DM&	WJG<��fU�%��(��E����j�2��ZZ0Z-���̧M���NKdZ�-P���0�va�
^��r�e���$����E��R��cXE����u%̟*���^f�1%�JK����b�mM�/`�2�r9����ѝ�l`:��ڪw\��X���)��HwZ���=�M9Ӻ;�.��ݳ���'���q��џmԧ:q-y�^Hۙ|�M4���0�����pz|F�B�u)�D���z\����l�/Wϵ��D���leY�ǜGpLz�^�΃��{�+qi�#މ�h{+D̘4Q�Ʒ���Nn1���f����*�gs�(��\�t-�Ӈ:�%MNrH]�H�^9�����K4�m��H�!���r��H��T̹��Pф��d)k�)�f�:�J���ޛ�w&����c��mg�D��|�G�k%!c����������L'��W�&��&Na۸*���`�F������A���sl="$rK���Ss/P#�kP[���I����ǘEӒ�Ѥb���X7�+\匬��vX���{Rѷ����<6ա�c�����v��(��.��t��c3{�'i��V|S���Ɏ+ٮ�d��x^�=��R�c7��r�)��R��p8JID��zx�
�|����S+s#���z6�{�P̙�2Xz�MU�w%�����o��$ϗ����يZ�Q�V�N�Dc�Z�UMҁlV�.�Y(�	[�ͅ�b�L�c	�8k��^X���#�fd���sOj﹙9�¨�6�#�ge��X��rP���0�8�;"����O��F���Aˀ���2�%�qK����@@�Z�)��~�!l��&%�f�n-�n�Ԩ��e(h�ۃ>��Q��t ��;��I)��c��9��0�+EBݫv�7^��r%�7s8�#��W9�����9�<[/ue���Y&���i��:c���o-��Sⷈ�EZ����"�Ϧ�f��-��G9��2 [�m=N;�͉$0�[��H����w�ۯ�ע�����Ý��`���O�����6v5�a+f��3r����ۙ��V��l<0l�P�vf�����8>�iR��>T���N�Y)��i���sov�.H�����u��َ3����kn���3��Iy�	�K3N�v����L���ٓ�
��:V\������J�����]]�k���6���D=sCo���&B%/wl8�G�jH��n���*U�?)�H�`I�DU�J;��a�-]'ڦ�Y�.�"�:���ۯ�S�u�bm۫.f���7�^�3w�gە�5q�w#�1��a���~,e�j�7WE�V���@ķZ�X�li�u�q� $�ٌxpF�iOxm�س+��u�]pgD!��5ԴyI��6'4ͼ�;���=�f%TE�z+I7�>l��y�����h���5Ŗ��D�6eAqVX:�Va�AGgq'z̳]� �u(�Z[t��<��5��72bim�B<�]��/{Cl�ZČNj˙V�Je�R�1���R�$ ���Z��1�#l���my�������F�Ǵ,viJX룃Dg�S4�S�uSP�F�i��y�pR��ߊ[��2�p�4v���2���D14�I�r���A�Z��l�,��a[���'�}a2�"\��@i)ø�f8�eC�x��a֖f	�n<rrDM�)s:qxk��G�l�b\�n�\+��ٟ ��V�qދ \HKݍ^@�V.ުkC�Y�����)��;]�I�����6[l�S<�A�Ժ��wi8z�ǽ�Zj��
���I7��\LB�>��)��.��5߭ o�t��Ü/^M�{^n�pq�7���	�Xr�sff��/�wZ��iØ��CrR��X�ň��O���/���s���`�-�#Ǝb}I�!D�DsT!��kM[ ��&]14���8��ZgiT-i���M*h]8��Jb�_|D���ֵ���n�a�5�� �y�K&͡�:H=�j&�hT'M��c���y�V�c�c7N�BK�3�\��
�=�����F�;�8kP�FM�r�M?�n6�Ś���]]q�Q�y¤�˷5�'J��D�t�]F��ö�|��j����^)���x����-8��tY�Հ�o;+�|�2���5vn�-�.
0棥͑��L�����s7��ki񅇶i�yP3 [��S�	J�����-[�n"��0/�V.�%YFݙ9�ں��9ghav�t�����ϸ5�^	�^U�+Â#�m�,�'c�_p�pn�ʚ-j�c��E�M�t����F����^���f`���eL�v�i�j��mm]x�ZŘa�a�w1��杝�ӜXz�qm��sbk%�Avl��\;��r��چ.̥�U����rM�עiL[�1�}`�G�]���ق�q����VG�6���58��38�wk8ɢ��a-om�4�؜�w[�67k*;�*�MJw>}�����j�9��i7���<rM��n#�ޝk۶2-{�b�����	��ђ�ٲ��Kd�ˣ����!�jR�V�ރG+�H����8+��
�='y�㙁`Ą�՚]\8%�XkLg+D'�gS��x-0]��c��D�.�ԄD2pۭ�,/��T�.�t��uj��[���$�!�rU��Y}x-hkKx����32�k�x�%%V.����8��<��w����v?��fa9جaE�g�Gv1_+j��e�:QO���j�j��7Q�����Y�v��0�� ��%���KWr׳��؜�-{1�+��˻ *�#(��o���f�8+���8�]�+t:N>�PǱГQ��̉{wkGM��I9�#IW�k	�%-�m��}�vLȵsk�^��u��!13ts��N�i�����._���FyE%Lc���S5h�r��E���07p��t��L�l��S
K�
���
_2�ŋv�3�-H<�^��'q�Ȕ���-`�Q,Y�XOov�ڎ9��X�Y�2vb�`F��Ka���aL�bˠ�lS{.�*��lИ�GBҨ�LZ~�v-y6$�i�X���0��z"��𼰽4�ǧ+�����=r�mV����rP؝��l�e!�A���d^3j�9�mH�OG��#;�n��B�MT ;�9�agbκ�m*nvΨ�˴2X�>ȝ�e��%M-�1�w��aaq���9����k�-�x��8G�Vf�ɧ�F��RӃ9i�&w�[�5.˨ۛ��[�B���'5x��w�S6$�(寚O��y�>��{�V'yk��9^��<�>A�Pm�ҙ^-89!�~�r����;�VE��vh��}��/�]q�U�h쩭Bu����Y��uޯ[��y���ItB4V�i��2��3�sa8�l���u[�5%�� ʚ�=2b�*�n�T"U��f�dm�6��bUX�*D�%��`]0�y����F��Ni׬�!�_�Y�st�zcd�ϡhօwR�@�c t�H�a|]."R����`�!;����Y��/�����6�Q1co��M� �Uk�����I��w{��Ar�Mѹ���͏Y�.���.R�f}�e�t�	�)Z�6×�٤�'121���	����[Ƽ0+e�㘍'F�ٸNw��ڏHdv=��.v�ůyA��^p��A�����c�5�dx�� p�6�fл.��uLŘ��)����F�y�ƞ�M\�Q����7�h���{�vNI�����c��s�ܽ��e���q���=�A`�I�����LxK��s���\A��B�RCV��Zl��;�&�!�9M�F�T�ǻ�A���.t��ǜp�պYsf&E���}u��>ɷ�Tg}&׹*�@xf�F���B����f��Va+��s��2���!�D�Ξ�A�#���Ŝ9q;^՚�i��A3��$�&k�[����Tp�!5(#A��WBYLE��{J�B�&v<C����W�n�[!.�p��zā�r;L�{�T���W{��)y����ز.��/r-j��n`���%`(��tKm�w>!�	uv��l:.��܏p��90�F�fvr�-	M8��a���6.x-��m8G-�[;�j��±��2�G y���o�Ћ �A���3V�cT�.����;����d������f�u��vdl��l}�1E�I����r���y@m����k��,�	u�;�ZsV3��6����MB�l|"T5��ӫ��ma�R�p^���BSM��:{7q��I�J!̣�]�J��l�K��hg.�Y��?~g^an��C� � AB�$?�!J����+a$P *B@�I � �,!I A@d EAd$��BP Y B� ���I , J�I �I R 
�B
�) ,	$ XH�IP�H�!
�$�� �	%d�( �T��$P�,�T���Y"��
@�(@ ��XH$��	!Y,�aa�
�J�H��I ,$�@X$ �+I*$XB�%d���!, ��*HRI�� Aa	
�KlH@P XBEP V@�!(��H� I  @ R+$�V�?�$���H@�}��.�>:��۽��8�4��A��$��_���W�uˆ=X�	r?!�{٨x�Mo��熡��l3�j�[��py�:UA<I�$�>���2��3w�Ej��n��T�ڏNQ�O��y�4! �}W����Yݶ)�@��s��QC��GK�k
ҝ-��]�Wڳ��Ȟ$�eA����{**�r�T��a_xx�Z|�>�f���l&߆vr��>�w|�њici�x���^�A�s�n����5���e�[z7�v��"	�m�9�(���8",n>�iM�̣5��{Pc�3�?&P���s:�F��������=�&���/� {0yB^�`[�i}�7���۸�u)�9���nꝒ e]���ٍM=2�;}޲���
m[{�A8�[ �*�}aZ�����QB����p�Ɇ�T��>�}��ہ���96�8�Ƚ7�fU������x����1bNh�;����`}�ۻ��d)�`�E�	�x�w����u�ᕈ'�����V�W�UɮRt1^��G�u�ak7�)^�>�)�y0E�L�q/Z/h;��:�ZGZ��_ ��w����j�I�T�&�1��2䇝��|�O7JMLY+;���֢PS����<Ǯt�M�+��˳f�o��T�v_j�z�68.�L�\�#���M�p��Q7���tvQ���b��ݜxh=�1zـ�i�J����)�ܸ���1�߫�M� \�o�*׾��7�]� D�빽|��Ӵ��+y�f����>��usd(�o�Wm��gD�M�5B�N�� ��2�[��Vٮ���e���*�Ϥ����#�紘��_+�5%rz�:�����'!ͷ��EaQ��:���po/Gǣ���zX;㘞�ׇ��3p��<����<A�4m"���c!�tUe*���ڞ�3M�{⌋�/\;������y�+�Vq�n�ʼ�y�ƛ�qʅRγP
D�ΨV�/kֱ�ec�;�T�K�H�4�m[��	FJ�|���5�M�)������	�S^��q^7����g���7�$M��x(Ң��.�
x`D�O����t���$.���Z�XsN���L��ܫ�"�ɿn����#�oxn�V�;����u��Pv��y��/v7�,g�����c�{)�G�\�{�e���)dᘺv�4#��<^��� �D���{��N�&^Nw�]�z�L��/�$��^��\��켜qm������[�]|rU���zz���f�▷��Ԙ1�i�jHu�����F�7��C����8^�}�h��T�=�&�"]cli�^��(\��J�����՞����0�ϳ�kxV���8�|⓮��jN����j�݀�@"�j /"��gS��i�Y�2�5�n6&��2e2��u�����,R��^�Y���z��[��ߑ��^�뚌6��*:�8rJӖ2mX�fi{�Z�mmU+���o	pCjW�����90�޾���έ&G�+��q����A�>͞�^8Έ�ia=tr���eq�=��,�tP�A�h:���X_��.�z�a�{cB�hcU��ŝ�����'eb�_Oj��c5�&���G�퉨�>�5F��k캆��;�<5�≊=���ށK�f�E��V��3�1��S�:���;_���T���x���k͵l�:���7+w��u�b�c�FY�,�h�>����Yx?fͪ��|z��y,T�|�=��2	�q0}�q6{�a�XW����������*���&W_:�Ʃp�7���m�$�r2m�.K��N���&L;��ٞ�؟���4O�`��ND=*�|�iS�A���=���I��{��Y���}C�ރ-q�JG�cE�I���y%�ǯ��Ցo,�cT��l���5�v��^^���)�\x��D�RG��zw�Q��Ro%�0W��8��I�������w��,�>��wlp�-��-\���|��'�3{8T|�93w$�)�����x�3�k�90��KF�/�vN'v�v�"�j�o&�헅���Y���i��^^u8��q8gY�2��T`�7�R�N��z�\Ja���_"��Ƹ"�:_K��Qi�͛ݝ{}D�3�<�}jm�w�ar�x�c�1�}�n��U��a���|!
�C��U�S}A�z�ʊ����u.�������5w��=��]c�Ww؋���12�����x��'�9Q��{7R�͙7��F�=�Ν��]b��S����G#=�lp\�kV�1m7�ә��=X��Fh/�:8Qk��Xu���_oB�<��S:�\�1�E:d|�M���;�&���>=�ɤ>�If��.��Ls�D��+{��7Ak�G"���Ϸ}*���3�̴!V�nT#�:��n�F��n�Ҡ�}Sj5�Ef�	���	�iv�q��V����g�(��F:Oq�z%^�&ڸr��0-�EMɂx�qeL�r0.{1�G�Ax��r�\�������sw��qtD���]"����i�YQ%�^&���͂ヱ�X����N�mF�B���z�.,q(]��Z��e��J~{=H{���S�mQ��/S{��$;R��r�s&�Z���I�j#Ӂ:�n�N!����n�!�#�|���Um��V�v)3����ʽ�)�냚ݩ�WZ0f�/oN�x�'�['�gC��Ӯ�:x�-�l����=��{��!��U<��w��/�����kA���� ��̘�b��&5�f�d��m��q�>�%y�=z;<����4I/L:\��3�
��[[�9T����u*P�>��%O�,=���E;��"�􁱛F=r��7"���S�-�yV��=�T�'aE��e�饶��Eo�[��������<���}&�[XI��e�"u��7M��K߇WJ͚[��-F��Y��.�"`�{�q:/��=w1�h�/X�~��fK#�+Fm�9!�k;��QVǦu'z���ȯYF+��!c?lԳI��b^:w8֣���®m-ý��)��
I��;��jW]E���ެ��*Vd�����g_rO����x?l�������k&dW7:^)y�/k�+�֣0�%��z��̽���id��A(:ꝛ�ͣ���z�~�TJ�zg��+�\Ssw,ɯ4�7e�X��OB��݈����.��/:mMn{V���"�g���.ط��\�!�8s�*-B��=�\�ƫ�dZ�gv���Ho�o]"pV;�-�v63�D6<Eץ�j��K*�X*vVo=��L�զb��;�b�j��}����<$���qr�q�W�tpqz�	��k���!���자hy��
�s�f�F�;Q�]�S՗��1 }�#~�Uoޓ�r��d@����gX=�FȲ���&�@�ޫ!L=L�#�����_3�PxIRj�y�:��B~�j�v~��Ręt(>U��P���t���4��˥���n�y�����-�PPvמ�m�q��h�N���OOA���8V&1��z��H�qy���+T�P_o"c����\:⋥2���t�Z�Y��P�V4{J��=D�����=E���f�=��5��夰��gm�eC�9lB����p!4��X܏��z�wY�fG�k��Y�i{-aC�l0a>�Z�ó��Ƿ�C�^�"]v��ۧ4�n-@h�~av(�6�[����2;�z���IS��e�kC.�.�z1�n�niK��͗��{/��ݮ뚳��d�l)}u�U�u�3Z�l����{=[]��o�d��U���buu�Yz���h���"���,��v;�������t�ګXfp��%
��X�y`��w%̸Vp�TE�b|�5wYӻ3Y�=�6�N�=o�3Ͻ7'�ɸ�1�`����w���"�,����[�c������� ���^�z���{.ռ�R��X����2��� =Р�=xyAw`�o��;��q>������Me+�������X�������^]���>V�����f{Z�=-fk��)�����{V�ҀpP7�F�,v{+���}����r��bՑ�LN��2��X���0,����[��ж<f����V;r����w;p�nV�D�ɏ1e�TԲ��Bph�s�+�Z_lxݓpj	d��<�h�7��K���=|��J��N��n��]^N~덺���ʳݷx�x�rqF��d3 7�$��<%�ڒOGL�[����ib�	������8	K�"�N)�Ex�����ѫ_ph�)v��05v2H�>XvA��v�]֭KqRy7\����gL�Um��Ҍ}����Pی�k/��Q�KZ>X3C��{��]D7��S�"�B�n&1� ¶�K7P�J@c�U�븨�(�;��e)	w	m��+$54�؇�j�S��Y|v���1s��8��%�ɃV1�eh�[/pN��s:<���Y���ϵ��;����"���z�4�]h:t!��2��MV/�=l˗�!H\��w��U�w�Z�7T}E�����V�c2yz�T�%lb�"���(��X���Хܜm0�F�ju��ֈ~6Փ��չ�U��!�ϪC2������V�����+�`@A}ʈr�+�8\J���%1G郙Mv�6M��%�H�~>��WR/����8�l7�N��)N>�j�Ժ�7��̰/OM��n}ƴ��Gl泱��x������>���$�*��n�^��PW|s�n�3��ܘ�b�����Jħbb)�|���t=�%�����5y�v[��ef��.-Z�W�&�24�TF!���H�=ӗ9V����	/����2�k;A��ğNS��tط�����۝Sd�n�hY��2���/�!�Y��J�~��J����1Z�֢���G"9(5��X�����B���/Q�RVrȯ]�o��f��Tm� �w���$�}|�Y����0��v'#�!��c���]��z�hNY��tq}j�!��g��t��;�ѕ�d��2$�ֻ7�5��)���왷νh�,�����d�G:��m*&�Z(l����A��^��&�^�裡�)�n<c\��Y鱔�'����so�¦i[�许P:��bWg*�,�9}a��C�Ǜϲ����`,���J.,!wu�D�ݦ*<V�K]0{@����T�k�t�$ekE�d�!omV&�õ���s`��&��0�l�Be��S������jip�E�.��Y�`�;U�Y�L`T�Vٛ�x裂@�{C
� �37�� S�s��I�B^}t�W����v�#ur�LiÏ=���?Yf��m6��u�fd�
��o�+�p/���GP��{5�5g8�ʽ��3����I��^�4u+�\2_B���7+���=	I@�x�QD�Kp�u��Bģ<�\*�W���x�e=��g%Y�4[�P�w�j#�8�rΞ���o����t7�.�^�`k
J�4���D���W�Z8zؽ�q�0��B����Y�d\w�*�.�u �2�yh'-�]�K휥;����\��[��FK�ks#;Q�����Vf^��[
72���*����u���kGzܻ�����|z�_T�@U1��zFR���B3����Ew'�h�,�t�(Q%�z�kK�P�E���}�̘�B3)}�e����Ġ�a�I#�.'��ufl�&X�4N����;�-[����)�ls�����u^$VkO�Eڍ"�Bp{:��o/+��3�c�=^���+R�a���P��&�����t�� ��������Y��,�Z��!5���#F�L�Z���6��͵�)�;�S�������Z{o������6[��ޛ�����=<��z����w�q���+�g���f���&���c
��3b�_I0͎U>��������ڸvv����6��lr�f�k�+$m58��c5������?y&��C����r�9f������/�?W�����|�{�q�h��t�0�L�0c��]�!�W�b��i���5x^<�ff�I�1�odaO{w.�P���<\fQ7$�	��2�(�ȞT���r|l��ҁm���陗�}�U�	SZұ���޾jaYi,�U�CAnuw&:䨷�r:��/�����Ə��8b`�Q����i���11�]Sw)�J��g6g;]%���Vs��<)s����ئ:�e,����fN<%�����8k������ؙ�'�I|�,��Ot���i�,`��k�`��e+z+�g]���k��,��,�c����d�DO�E�]\�箝�ӷ�j3K�V��|�/ W' �G���=6w؅��o��΄İ��������e�a�)���r��>���p<\C�E�����j��Co�8MA�x�*�d�:r�0��q��v�C��#HiB�)xr&���Ŋ,����(��:��Y��Vi��n<�>�l��@�����>�a��.¥w
}��繬ԫZ!����h�R9����٧h���<��~��E�p����q�v����~<��3ۼ���;�է�sE��òT2v���2�;�-˰5�y���jhg},��U��?VXfNg�)�������++N'r�ܷNiRI��mR�jߢ�z����j�+��;s-�ܢsYLN��h��[�M�yx�踋;��0:m�fm�e��t�׀���G���A��U�Л����"fck)��ӦI[xi�M�q�^�n�ѻ����{����{���~�ٮF�ƍI�Y�����Kz�8��d�bZ6��K�Oc:��^m����*C�d��v�v��+�g5�c��\�5(᠞�r���v���֢��S�Ԃv�6�;���D�[B\9ݞ�R��������8��� ��[�u�Z�kj��=��6���li-]<Հ��WW�;;<7m����-C�[�����XѷER����<f۞�u�:�m;�Ϯy��k;{��n$�s���U���;:7Wy���2��vv�<u�c�jOU��s�����CsXkd�f��ۡ4h�c]#Yˬ[����5U�Bc��&<vm�뱞�3�on=zk [p��E�km�;�W��.ܼtg��{X@�ܪ�{��
=vN3���M�E�=lY�ck�|Q����n�x8���X�uۮ͂\�n����cg��yՔ��ó�R��g�:}u�C��s�x���.{y�=�sI���gg�M˗����M�)]r�\s���1��\�y�CB�y-�v���nm��܏��'�����qtr�'CwJ����a�:4�&��t�+u��;Иv��׮[��;:{)���`���͊�A� s%j-�ɵ�$ۇ) b�b꺸��-�^�mТd�pg��<e���ny��>C��O
�S�U�җ ]�:<e�R��n�,ܒ���=z�u�ge^�y�;M�p�nN�{\�gN�Ve�P��m����qgy��-�C7)�v�Ź煹�����Mѕ�;F��.�v�s�5��3� c���:{[����.WQt�5:$��d����.�rc	n���Kh�s��!푹���[y���sl�N��WN;scV��m��t�]@�Xݣ�c��{lͳ�@v6ͻv��ϳG��ɘԜl��lۗ�����q��Di�۔Qzp�e��tgp�a.�Y��unA�j��1Xs��n�����7��&r뗭�l��9wYm�pAۍŰny_U�s[����[��Q�!hj�����en��!s��Fx�n�݃h�c��m�u�f���u�Ge�qu#�}<�9��zݦΘ�<�^����u�9�p�Ø�Avݬݰ m�瀫��뎻q�8c�K�"vv�؋Rǵݦ1���q��Z�v����Gx� P��4��e��>��:[r�)��F�sr]=K�N�]�wG>�O�j�e�[mƶ��kբ�g0�Q�T�M�BR�*b���z���՗�zC1NN�x�wFz��#�g���q-rb��F��n��%������F�zmgf��Oc�}�V�����i��-n*�R��;���!��띟Y�:���絞�skl6�����D�΋��N���[���I͵��{d�s�Ź6�ې|��/=u�4�G	]�۷8�c�u�ۗ��՘M�u=�\n��m�X��դa��=��-�dd2Obe�/l�{s�bh�ݱfB�=���BwY�lq���v8*�5�)�wHJ�3Χ�C�i��K/S��q`ل}�5����SF�]�5���u�iN�Bνchsuj��!7s��n1�^��Y뙻��6)x�:������n�[5۞��ҏ��6�t�h����0�m�
/��<M�g�qz�lg:K���rfy.x�;n��ƺ��^{k��n�&�"1�����b��óƗ��������ێrxE�I�ǵq)�ݝ�ͬ텈�L�Wv]Q�+\��[m��vx:�e9�>��v�p�=���LF�1ym�5���t3u�/n7�R�/�e�����Y�	rv��Op���آ�y3�ϴ=���-�Ź�).��۷]��\�t�p;�͎Y�vX퍀�2<7�p1��Y,+�S�r��<m���,����PX��jz�s���i���[�q��Dw9^Kq���1��Y;KS�^�l�n_c]��.<�#z�;q�ݞ�xc��i��vbLkm�F'&��yp���5�\v�uՃk`݋�+kBk�G���v'Y0������2>z���\`�n��6��=����s�ٞi�U�W��2�Udy�2j�:�j���f���㱋��k�z��z�2lI��cv�Y[���^I�[)����nx�X�]=����H�Ӏ�[^P'dS�f�j"v:wbn����;z��[cl�-�Q�xѭ���ك�����q��x�2wfؘ���u���P6��k4Ψ{;U�];�qt�v�N�gv��m�Î�^���s/\����J������,��f�muر��.��p��]��.�n��������[�[���o/k�-��V^rw/m������X���Jb���\#����=�o*��;u���x�z�ŵ�-@�ۚ����ڲ<��Q��Rһ�g��k <���7��z�n��t��:���í�c�ݞ��ۄ��&�d]���<��v!Nދq�����vM�ێv�4q�)�8wE������\koM�`���z������q����9����y��Qw��z�C��O]ree.M\�;�Om��ۗ�n�v6��#�;������lF��ݗ�q��,s��G����v	��ݵ�q�ݎ�ֻ���	Vzܼ���)O dʖz1ў
�:3��P�m�'���l��.�t������e�u&�C���˼P���jLc�C�� m�
b��['5!���9����Z���zڐ�._&����ni�>��wv����y���7�F�>s:�����	ލշ=�Q��u<�ս�����Зgm���td�:�#�v�5475��v�W�wv��t^�c��uÕ�:r��g�dѦ܄Q׶ۧ�nsG��q�J�wn�=�e�᜖�܉�$�����7��ѧqV�]GS�r�0s��'WG`y��{k�Ƭ���G@�r�͟n��P��7��M��݉wGUs8�C^��6BCJ=�ޝ��j�\t^�ۣ ���&ɭ��0���V0��0g��q�n��9����X�)�hz��{�zʧ4]�Ss��k����Z�kĽi�n��Й_n���K�.:@x�Ų�v��w�������x�I��&���<�6�'�cRqq+��L��r��k��U+dg��kp�{z�FݎH|m#j��u]�d����\8���ق�o-�,"���'Yۍ���:[�e���k�6�ޫ2���k;������V6�.���b�6��9PѪ�ѵhl��nXl�[Q�c� �m28�8��G�������+Ѣ��K�i�zI�q�n��y�hׇ����/k���Ѷ��#��<`+8s�=���v%Ϊtc�GN���qs�&��n%��n���u���k���T��Ӓ�֬un�n���uͺ���\�6��ps��8ēڤ{Fg���!9֎� 2vڔ��ށv7Z��2�r��p�'XtJ\�;�]m��s�sy���O[a��
Y��*����ݍ��t>(��/fpݮ��kY6X۪�y�M����ue�X�ҡz㭛���c���1����r!�
[\���v���D�z��@�1�p6=C΃�K��/�L\.5��wF���.��m��˂Y�5�v��f���r8:�k��b�[K=�v����Q�g�\Vϐ7r����/m�;'m���ޝ�'v��»�&���v�k��9ݻg�n:�۷Vv���\
sr���ӗe6��݋h�8�i�����ڊ�����.h-M�S���x�精ؐݴ��ۺݧV�s�'7m�d�ӸhޮδoGUu]�:�[��p�ѻ+r&u� �u�O=�Ʊ�ݭ�p눈z����y�lp���5����c��܋c��p<���:�{U��R�m��ѕݭ�r��n�M ���b��δ<�s��^���;.;=�'z�;�=b�/
�mA�z��붗��Lr�x���I�=�LE�y�^y8�6U�n�\R�]Z�涛t��s*n�ƍ�^ۇ8;��"t��n���e��=tX��e��:��xS��!�k��NZ3�[c�GS��\�4�=��������q���j96 �x{p<;�c�/��%���k�^���n���=]K�pgm�lY�Y����7�^6�]s�J�g�.x�8�؃m]Z�I�=e�r=/���eS	�����]3�kZ��n�vy�qwc��q�5�j�t�z�l�[v��Uue�u��ۜ)lg�:�۷���h��҂J\܉�ee��u$\�v�h�"��%��M{J��cR�/[�6cq971��F��Q����<�v�Ҽ\���f�G��nޝxp��t��8yu����[������h�ٴ>�^'����5�Q�<��mh'=��",�5>J�Nm��Onr�c<��d|[tE�gٍ���$
:����h-c5��Q]��a��e�Eȧ]��=���v��%��W1����n�uA+�v�.��l���'%�)�-�U]��(Pg���2j�,���D[�.�f�m��snx����G�Dpvt�`�S� ����r[OlqS9�d�j���[V� ���WX5ʻs���&��N�Gi��\ۭ=��Z^;\j���Q��k�0ݡn�bԖ \�p���֎t�5�N瞺�VJu�L��ծMY)��:�vz���]u�j(�����N7=sv�ud�苋L�=IЫ�\��Z���r�n�{/7<WC��N`{>z�R�Ѯ��h�2-���r]&�í=�p���1��W��р�4��nln�uρ�>:��m�k���v'��`�ˍ��:�lXWl<@���{cQ�V՗����읥��㱶��bC��Ff�q�y����N�Z�N�z�=���6�u�n�v�5�;��[�pC�n:�0��`{rx1�C˷��6�U�j�b:l�1t�-۠�g j�8]s�1ėigwh/M��lV�l=ߛonݷm�U��=��9lQUz�4TQV
�aTUH�N��������Z"1��AAH���r��0FETT��T��-E��,m�((,����eE�QE`T���Vڨ��-
V屉�&P��9[+�TU5�0��(�R��Tq���f!U��ڔ���EV(�Qtj�rZ�Kj7)�������f*�QB�Ш�.P�B�Ԣ��1PS2�-J"�QQ��s-�KX���PU�B�+FcZ؈�@�(�(�Z�1��7���c���Z�b-K�iUU� �Ib����Lee�EEXֶ��UiJ�b�+&5�D(�֪�ciQLq1DX�0ũ*-d�V���K
�Z�-�
bL��ۍn2�h-V�@S.fe"*

�eb��AC+����V�Y1�E�-q��7W-�WY��5%D`#]=��{���������� �򐖎��c�g��%�ۚ �f<�r��"����>v��6Y��]��� Ε��gC��p�v.� �6��,�{��X�8%��χ���	�6M����+M�s������ ���csg���:�9��j.{5��ئw@�wl�6���`����_tԆ����6���6�;x�L>[��3�Nݚu��nXZ^g�˳�u�}�ɸ��u�{]��º7]���y���x=��q�o<SCPq���:�� ���]��p�f��Ɍa�77z	�K������������d�f���*��/k��0����G�ݱ��wF���E�lv�ظ+H8�_���8ݳ�b��c���ہ�`듢��jMŐ0{R������Yc�
��8�w�d�x��ώ7=]�ַ�^88�l�q���2�v���u��"�C�wh7\v˫�:�ݛv���Rᖶ 8J�N繺�m��>y�=<�u�����m�n6�����;�'���9ۣ���׮6�ނ�0��v��vK����ÖK��Y���2�ưupv']e��ڴ�x��݊�Jg,�^.wE����w]{;���q���U�䭬ue�v݄�r�lpɜ�/i7��b�Y�q2���;5�Yλy��l{m�����=�.S���2mʜ�]s����t�:0�r���;Lv��n�X��m��ݺs�n��_Gmզ�d��!���Ӱ�\p�֢y�����.��u��ӳ�ѣt��F]���Am���Ob�g,Q��n����o9�ofR��t���1p������K�ή<�Y7n��,����R=�E��|�k)���s�g�!���Hn������Qڷ	Q�b���ײ3�ٜ�yw��Z�N͵ۦ�y�c�RE]�o���վ�i۴��z˔��Rlu/��V�x`n��5 ^�����g�����"���Cw��z���l�{/(q��78s��&)Lp���VdJ�Z&fa�!r���[r�p���[J��ûM���9糞y�yq��m���l�� _v^s� �)�!�{m��e�r��O��x�aNCaL�q����`s����l<��ۅ9y��n9��˽��re��*�����v��n�N�s�G�{'g�S����;=��rep*������8Hj7W��~?�`�z%( 	׶���E�W5����{3 _����q�)�S,��M#�6�I�ӯi�C�>�ݝ��6|�U��: �o�����8�����8����U�t� f]���ѓJ 6��� ��}�щ÷��ϒA$��h��_����VfS�H�"~sw�=�܅���{��OJ����@��l� ��� �����]ׇD�O�*���>3&�E���LD�P��=�v� �+w����=���#� 	�o��
���|��1�u;_i��TR�tl�!P���ir��K��cpݭl-�љ�W�޹6:wq�+}�����Ή�����8+cf�{}T�g��ۙ�6a^��{�m����힒�1 �tZ�$������k1j<��tɢ}B��)�ܳ3�#2��t�A�S�˷�#�}�w�����V��)9m�;iɫ)H��;ǚ2g�bo�5�+�~;��VL��L��d ~�Z�$�������2Ms�ATr�]i+����)�%� �������n�`�N�,�}Q��������P	�=��Ł���P�+��nf ����Փ������J�Y~�Z�H�s��x���GI�2moBy�9羿]Z	%>ȑB�ȟ�բw7s>��t҂zOy��ŝ�uh4��I$���n���Q�6�m������}����C��^�\��5.:�]�ƈ�5�,�9��x�W���[z)��Ә��ɉ�
5s�W+�	��^,�}>�������t���Tߪ�>��bX����2HA12�`�D�~Ͳ�쿜�_�Y=��4I$���f mϣ����=5�8��&�^֠vΒC �%D�3u���X6�l�P6 �ͭ���AN1�dz��غ^��)�c��t���ܒ��~eӝ%&՞�<s�ᣙ�r�.��$�F�P��[4.��3p^�=vp��o��}=% ����`�1"�YhU�v4��{kc�-���x���� �O������1zf�P:��X]j�µ
F�b�����P]�ʧPY���������@{�ݙ� z6J geՇ/f}Y���:�<鮋�b��d})��"%�-��Q.Ѻ���(\��r�`��-�>����ݿ~��Pv"~s\�����c��l� �;.�$�^�Y��/܆s�m���	 �\��Dx�(�D�3*�]]�N��P*��ڿff���\l����޷�$c���8��U�Lߵ/��Ƈ$�9���>���۾��� ���'����\���6|u��@�gz����gI!�9�d�3uh��f)��2}\��}��o��
 ��{�M����o�n,�E��m0_�����+;�1��z�$���;2�OS�	�̝�n;ytD�k���w.��h�z/�.��Ix �=Lng�ɦ�V�C]�o��숢�޸�fX�I"�X���g�� ݾ�XR��Ga5ۛ�wL�P�o�u`�;�췙���7���½$�10�J~�!2ۉ��+���M��ͮ}��`Ճ��ΞW�r ��������t�����6�2� -�z�� N�{wR�@�^�m�v˦��PI6z���Or$P�F��{���!��Q}�Y�|�<�z�� ���b���5��Ƕ/"�ʀJ#�b��9�P(w��������� <� �lê�$1 ��>�z���wz&ț�Q�0�2�,�'e߽5�~�]���vתՀ[��� ?\G���v(ز��>���':8�AI�^������	�K�%��2�N��u` >+������1�B�uZ�=ڮ�r�dz��9AEoXr�����|�[��c����|$���r,�{��Ƈ�~�-Sf�b�W���:�7oϼc6�֭k��snɄ闍su�Om;�&���q�<�ulqg�����v�k���g������S�[�;tg�����_:��96���2�m�c���pt��0�M�]e9���8{E��΋<^țvqk%��X�Ӎv������%ש�۫�����-�w7n\�S6���x��f٨�\۝��/,yh�$BS�e���	ŇF�'	9v�W���W��q�㗋�<ȝ����=��Ʊ��7�������`��?$*����A[�뷀|���Pv�l�*}�h��r)?w��� 뻽x�>��n�c��AV�j#�+܌�����)D�U<H +=��� ?eW&"�I���O�j[�#ē��ØR�F��q��{�m��pR %��ʓf�_Ov� lEg��m���a���-�&TB�X.����Y��}Ȼ��ܻx-���� |��-s1�{U����D���4�_����6��g��h�~$w{�Ƿ`���6����1 :.:*������+mFV޵\(���.Hsbe�=�v���k���CV�W����ٓVܢk��lV�?~�.���Z��yU������S��w�ua�q֎.������ب��\l4XL� ��W�v�ol�~������n�`��ia��Q㫵%��.�Y�wV���}�L�����~ ���ӵ�q9���x0�rB�r]�]�,�H8��(��oD��=ޥS�����a߳%�@�����"��*2�� ݾ����N����'[ެ� >.6+��}��ՠ*7�b[S-O�n����S�ٓٱ1���L� �w�V�|>���&g���p���j�o��J���*ƥ&TB�v/m�݀	n��>�ݲ]�Ua��|�gDP��]7`=���U2n[�����7F�t~5k,q�Y]%J�E-��z����R�J���8�??|�Jr���s0{�
26� m{�괬l���f`o�f
���Q�`	�{����s�%�I&�x��z���K~���/���]�} ���� oo�>�� ��*brc [�.<�XK�Y
�n��]����H9�lmygߪ�y�)�7yT�rR�������VI��k�9�\�P6�s��5U7U�c�yQ���\��-y�g}^w�C��>���� :�tM���.��' &�.�uŬ����W5����@�{�iXeww�1 l%�e�Z�7+	���I�}C=�Z�$�Q�_�2��h"~svO�w1`|:攁�����XB�>��I�n�Z W�}��Hz:�)�c���*3��<�g%�i;#<NMAؤ렇-��u]����È���"'������p�Q
p��- "s��$�I��� �r��(��ޭ�� D��ٟ`��ܡJ�"j�bMt�$�#���9��D`�x�@�>��f ?sA��\��R�f�x�����/
E&�`J�����i �4غS 	J�ڝ�=�j#Ӱo�\���m�G���vK5@Zd������X�=�?�>��{�j��� 8ظ) ϻ޺�W6���m�Fï���� K]zn鉨��
B�'s]��Fh��Aה�����[���q(\���ŋ��o��I�3��I�ẕ�ș�����.��ZVj��c�e'p��ݷm����}lI�{�VO؝SxSA=�I�槤��E�jwk���;��ū��t��y�J]��J�I<��]��_��+�&�	 t])��}�����8U�U��j8��vbX1 ll\Tǌb�C�Éd(wz��X���3ϊźu�o0 @tl��	�{�V�AJe����d���&���v�j���^e�TJ:6�Y����d]g�
��<���� ��������=���I��J�}o�ڟ髑X[9���Vt�NE�*$���Յ���{����z2+��rY���L��",�+���k��wט�:�2*�����&������ɫ�1ǯl������RBٵ6�v^�j�Uن:Ɲ��5s�N��uJZ�٤lɂ��׌h5�M/�h�b��WL�Q�o�����ݻ����`L��>��KdL"�������u�t��]�Z�l���aX��������f�g[9qLA��sӕx�v4�K��H�[��]X3u���Q9����j�5�p��m�a.���|�6���D�b:��G@3�^].a.�8��뵳a��Vw<�F��nw�Ѵ�Ռ=a<�u��[��]�ۇё��uļsы��y�rюH�����v��93[��L���:�%�*��;Hf�&�knvy��<<��f2ߟ�����T
S�W�����^��]� ��n�O05��~��9�8�ں�t��������w�̦�Z��ݤOo�1`��(q��]I��0|�w޺�W��2	=ݓ}����U�������6���Q�'8ى�w�~�I=�-[��e)[>��/�v瀞��/}����ޖl$(U*��I�k�UI:��nW� w������7��� �G[�~c�^��� �MIj$�����$�D]_���f,�62yo6��<�w]X6�}��X6ϏGFE%I�g�,̜��&D�U�mP*ŃD�kOk�< nݷ��v��qwg�8�����V�����58)�E�w�w`����]������D�z�u�Wy�� K;�ۣ]�'���L�Ն� �����,�_ԟ�T�V�U�ݩ,of���K���&��@�0���R:q[�����&Z��Ȭ@W	x����g`��Xg�fn��;ꮱ��ѶI$�~�{Ud�o��)���UY��9cSڙh"~sn;soV�J`@��L�;�>U�\_�'k��E�� �tzS1��H!�B�w�nn;�ݞ��N�� ����ŀ�@z:} >��]P��{���q�NI���$�w�c(,JfB�(���o�՗�TET Y6�d����m�H�����&��n��EՓԧ��9S�PIB�ԥ�e�|�GM�.ݫ5���l�֜l�^ܛ��Ө}�-_��[1�@(�W�e_�-�7����D�@=�z����m�Oǲir��Gz��� :�T���f�$c�a1e���"lo��f�r�n���t�2~$�#}H�{��ՠ���u�2��$J�1e-b�I�k��6kg�@[��a�'슌dAX5o��쪵,:�A�>t��X��eq�u�g+�:c����s�X���������G�
��ʻ��������u��V�g�k�>南|:�б��&p1��g�Ɋ�!�(�Dh9ǯ5͹� $V���|;���ϧ��tf��LA`��B���1�i���LYCKS�!��8�c-�50�;��`�X7w�ڝ����}�I�N�8<s���9I�<��T_+�D� �"Da�}�mi��oa�ǭ=�Fƽî��m-����`+ūY���`�+��eЧy:���w�ͫ��{=�y^�*�U�!��R��_A�H���7�V��
s�p�\h�|��Ƿ�v�s���A����u����j�j��^]ʹ�m�ک;7��M�\�w+s�A�1�c�Kބ�9��.���-!wo�ru�h�x���>6)D+%��K����i	����;w�n��uXU�-�P�������h��>�;�b�U�ˇg�Kđ�&g���N��{w��q�y��ȹ�O[�b�V��-2�.+`��*��g0�м���x��j�Yߓ@�w<U/�a"����g)��J�����vHh.�hv/	0�{���er5
g>���ь�E�w�d������̰�`7O�A\2elys���nV^�㭸�tU�O[��^��z�S�-X��Gӄu��vA"��0�g��GQ�{p=��S�=�+�fmL����uҧ� �5	�",r�-ah6�l*���*T*[V
�ڥ2�,��ƴ��r�!p����ʙ��b���FJ*c-h���"�\n[�V��YeJVU"��:,��-T��ApK�J�
��Ff6�l�Ecrۙ�ڥQ�T�`��fQLq�9Eu�a�I1E�,m�l�eQ�ܖ��A��.9���-V��º�N"T��GM�[KPZ���\��Kk���0FfSZѵ��`�em,��,��9R��,���%�Z�)��R�h4JU�-*,
�ZJȥeq3X����c���7C����!��1`[X�mj�q��31F"ؘʬLU��5գ5V�.TSljT��7)h��3-�
�hť
��ej���[Me(ʹr�Z�U�Y�C��m[LB�[R�V�y�⛭̅fb�V���DT[IE*1��*�m�3%�+r��2��S7f)�+�3,h�8:f��ZT1��Mh���ֲ�R�X��qˌr�*c�lkh��v��8n<d��^��pcQew���(Ѡ��֔L�3�`t��M���x��l�D�[�m-(��2��Z�?e�߹��;�R3�����T�_�+0Q7�J�ONn̬�7����@|�2 �w{�V�H^o{d�+.2H<��Q��;�W�IMՄ����Q'�T�D��Lm�i�+�����go��� E�������㣟��
*f��\��7A��3�/cr�=v�L=u�k����wq�+|��߿�\`M��a/��3�����Ԉ Oލ��/wܶB�OA^���>�z��Ozu��H E՛Wٖ�3r{�ꢩ�vT�`}޺�>���X6��l����{ޚ�7$�{�{��NH�2��EK�T�$=�:d� W�|-���\�UtE����u /;���*/��T)��L͆�]lC��'�z�z0�.��]� }��f ��V�ot#�!�i+�d5k}��]I3���:�\�]F��mz�{/�)j�h!"���w�q�������˕>��o�����_B��̍L�ȟ���N�n[��w�f����x]j���M|���c�nEI1�S���Q���~��'��ev'i��m��:��uz�����aN���<ϙm�����Hd��Ag~{��Ս� �oz�` �K���̗{~�ɛ� �w���4I��ލTf�:�~�&d.�PwR��q�|��B޾�V �۾���;�R0	��o(�C�P�:�̜�����+�U@��͚�f}� ho�)� �gul_Y~˚ʭ ���Ń>��E} ��� ���9h��%�Z�2����]8l��]� ��DP ����{f�C +�;3W�!�J�?8��T������U�em�j�4�3����nf �6�R����Ua	�*�k��i�l�	�]%���0������7|������z .��cr�e����fM����m�������#j��|wǇ���CmW+\�z7;kfs[���À��]�]j�ɓz���6���������3�p][���6���ɵ�D�^+/l(ۮk���5�pr�1͍�v&^Xxם¡�������YՋ�k*�]${T����hDۍaBsŒ}��"����OL���;�S�&�u]9؂����X�{q�h�S];[��rA9�nf��f� rjܴ�Lpg���m�'&��m��i@��i�u��-�>�������{t^��g�4������ ��T�`	�{�V�?b���oѶA$����X4�/�Rj�D�$��w�>Wwk/u�]��6 ��D7H�޺�mM�Ũ�h��z�m����D�"DL�]�����>骑4H
�AIgƦ���{����W�0�z����N�����HUc�v�fv����i��$M����m�}޺n�	�ۙ~ʘ�)z] 1�QP�,�p2~d˒"�B�˻V��۷���]����2�TL��;���� �ۘ�q-�H29_~����N���׮��f��� �����V���L��hݺD4r���Ʌ������~�덚qs��E�_k�ޫV  /7�3>
�U�zyzȨ�<����P1�{�W����Ng�R�3�O�71,�*/8�ꛁJ��EU��u�S�_�����w[!00�ނ6��k�E�)������\�׽��2�1�#��Q[�Z7z�Qu�'Ě$�$Z����O�@[���	ׅ�,V�
X��nՂ����π@��݈%۞���mI�97@D����w�2+0�&߉���qI��=gm��[a�6+��f7��ԙ�MK��{	&�;�1�H_���n��5T���c}�����إb���~�G�<�˫������z7yu�5��|�g
t^C�P�[�m��(���D�Z�Mu�n'q�涎�Y9�cِo�1��d�ɗ$F�w�v�> ����"RH{�Z$���R�[�{t�&< ����[ĝ�"�J��e���sP;��D-/z���0,몧� wo�3��NIH�Ai������k{DP��+ 9�H��A�L��b�I�`ڹB\�����7u͕�����A  ��U�q����!$�4e�yK4�^�=P%�i�F�Y���~����e�fQ�"u�Z�u�N�k�6$W���� G�rF�Lx�[r�$
d��]׷���f��n��`J'd�6I'�O���4������Kp��&zF�̉�OX�F��F�0�h+�dt����Z�h�����v�_��� N����I4=��]�������~ݭ6y�^������sm�NV��x��;Odrk�ح�����wi!ʇ/��Uz�� �rjA �O�޺���.*�dOǧ;ٟ`Ā=�vHj"~sIcS[U���E�x�ݮ��ܸ���$����,m�{�-D���J5�	^�ç3¨�ҫ�D����r.k�.��S�@�"��}�����6����9% `s�z����q�ә�T�L���v����a|_3������I ���s` ��w���}Y�UJ}c�w�l{����r��0�]��,�X�=źW���j;l��T)g����l�>��>��5���vWs��ٙ�d_h�$�ɇI�;Īr�52B�Vs�ۿ�+w�x�����
o�}3=C�>�w�o� 	��f`�����6�����2��f3�IV�b��e����W�/+�u�����Tfw�rr��2�+#�P�Ui$�O���ۢ^�0�&s�=�d䔁�}�w�l�J֜A$8��}Fj�n�5D�&[�6ⷒ�$�~�}�@ Vo{3|�/�����9����O��)�R�����H$�{�׋ ���v��N=�ۮ~�g{�6�@���X:�Q�I��a22彸����,Y8�;�9@ ��7 
�5�z6�?L�L6��?OkfnW�<�<�c0�1w�]��7��Pb�'y��~D(�_���6|W�}���}#|t�jɏ\�e��VR�#�ɕ�F2�tMw1OX݊�ޚj=��\^��'�>m�E�mH�o��yL%B��ui巠&�z2�Dy�ss���bU�S#04���X����\i8�q��x\g==��;=t�.�t�=f��7�x��8�`�ʌ�!�-���q�v��mq�6�(�v�cc�Z�糬뎉���c�]�rlknj�Yt^K���L���n	���J�E�i��/rLO�?>F�&=<��98�s�n:�`���r�f��g�����n�sF: �ѷf�:Kcg%ɞk> m˭=K�+r:!y�bS�����+WGD`�s�ۘ�'9�Nra��:�y���P| W��x� Ht��A�{a\sd]��R]ù]��ŀ�W�59Ch��%��d�IqZ�f���ɸ;�HV�z� �����)d�5�z�L��$��c�X�X�$%fs�����ݏM@ w��t�՞u�՗8�H��ٟ`���K����C�O�Dě�V��+1�N�g���=��
��D~$wm�������)�#���oc��R.�+��Z)���։]<ĠUz-iV,��=���G�\,GW{�i�qЭE�=6�dS�S�`��Aҗ<<��c��)�h���u�j^���[��~��{f}�`e��(���P.�i ���$#K�av�z�}@�kJ�k��U�P�I��RuF�:�&a��Z��c<nۖ�����HWm�qQ�w������|�y��˻�|����/���69��W�{=k1��9���)}���C9��q���"g\,OW{ـ�`�y�I�~_ڸ�(�]�O�~���H�zy�Ēo8I�Wfr#����L�Yuw�@{#�/}wd�J���6����{����2�H� �\�J�����r���P2��L����x@��McK'��[A �Λ�e�c�����94S�$[�e�WO<�	�ݭ��.뾾�.o�w��������"<q�F0���I�w>�=�bź{n9�vgm�����[�����?�Uɘ�����ֈ��<������c/۴!9?W�fyo�
o�cO����Q!�>Ie9���0�n���� +��3>$�ogk񦇡~w��3	Gڰ�0���v-)��*�+ᓼ�n����{���p�izF���yI��z2�x��%�_{�8`�n���v+SX
�`˯tH��`_�&rR�|n8^t�{F8>1`��>w=�c���S��hԄBh��
N{c��_��pA��+�< �E�M���H�ۆ�����B{����f|v��jՊ5TP�x}o����%�V�c�{<�_ ��i�#f6���eR5%h�TJ�b��$u��;���v���:��n�fcoc���~�~�!jH�s��۵m��ܻm����з6��B<k!�M$(P��I
�z�qr2�q#.�z򲥽0/�/ �wS��A�附�~��)�H04�_^��&ܰ�w������f�g�a ��vAZ��T��]T� ���L��)�?]o�a������]ش���x9����i ��y���Sz�$����<o��U�]�>��u�ܚ��а��x�L��z���l���n��ͧ�jؚ��ki��P�Y�S.:��������O�<5!�"fAC��}-����j⳩�vY-��w����c�d�Wv��R��o���:(�M(п��{[[q�t�m��v�]-V{�DOnָMɶ�:�W�Ww�~��j��(U{�m�3$�1d	]���jP��Z������V�k΅]�!��H�0�!��7[k��W�^osRڞ�/ZC� �c������I�zAn��揰��)��#V��<u��]�C5�Uy��7����߁=�A��]��r�`��2���1��R�(��r����≇@�{�IM�1��{ݓ�y�faz�`�>�I��UF�}S��A&�;3�滮>���|Ku�0ARo�( (=�-?}^DG�x���b���7B���:\�����ro�mDԝ��n�f���H��8�����*�!��/�Ĭ�G	�]ܵ�8/?�Lx�
߶��7�J�Ãf'|�[F���]��}�!;��ã�R���q����&������0�8F�F�uC�:�H��M�8"W���6��g�,<w
8��Yw!�#Y�mc��{�����{Jg'Iw]L5ی�nCԐ.���9.��=���]/�Ȅ
<K|K{Cwq��1P�*`���Y�E��������˯u�b��<�dݻ����,ph��Y�����/�`�G���Xo�Y׳G!�M���S��d�;��	����n�p̭��Ncy�`��i��f`��y����C��Y��k ��cިWu4�Z�÷b3nu��B!�d�:�v۬�W�y�{}��m˿�{,� H�֬˪M�n�d,��m���&�>;89�+���9��.��&�!�g[]tp0T��6�ъp��X�sF��y]iqp'Lu�U�!]����NZ����]�ug�+P<xޜ�)�"j;���{~�:)���8�%|E�WjH\7T�F��1�>�C��0�5�&
}6��Y�s�Wb�ԭRLj^�t���=�ds�ʊ�W������'���]&��S'�{��0Aؓ�[�Z�c��/��.T�(��fm�5n��ʜll�u��_p�/vq�
�2o��f��ֈ�V]�پ�B�+���7a�͵qY�6��55�t!�1���_'כo.�볆��6�E�9h�ƥb1�f%�����V8��*Z�Z�^S2���KV�im�V��"R��GAQ���d�Ɉ֊�.Es.5�1h�,R"+U12�W͍�nN;a�8�{6�1-`�2Z��(ev�Z�El�`��k)��n���s�w��F��2�5�F��ܸ�2c*��U,��jUˉ��ci[h��2�k\il����HQq����j#\�V9��cJ��r�K0�VP��d�m(�e�ѷ.QL��㋌�er�]\�-Mb�li,ᘣ2�f8ZV�Ъ0��1
��X��#YF)U�������b"��Qm�ʈܱ�ln.-��ࣷ5[uh�ʕL�X�B�*�KJ[M�,R��3W0mkD�UXbUD0�A��������V�[��m�֬ۘ���1DF��q2`����*ks2�%EYupQ]\�b��әUV&j�
�[N#��"�*��F�\�q�*[��e1Q�6�Un��ݱGmwJ"�*��m�.Q˽C��h���wo���<���F�J���x���gv��И���Y�qŝj��y�n�TV�3K��zŋFb���Q�⵹F���x��;v�;�M�L��$�G�q�]��ٌ��}u��!8��UGWFI{�uϔ%�ˮ܎�/i�G[���1ԛc�p��r�=�]�.�qŞ,79��9�hj�g�w�g�F��	��v��n�=J���6�:��������d��N�tv�ꞧv	�cQXV`��91���6��l��;ۨ�r�C��f��]����'�;/=����e�c��6��aR�k�s��"��]nֆ["��=rq���X���㭞:�ݞ3��d�+�O*��>|�_mۋ w2�5�>�1�e�\����eu�cn�4���d����^�70���q�3�_n��4�udm۰p'%v�:��&4�ӧv��i��[g`x�lt����tا���{;]���&yݧ���MLcT\uژ�n��!3֮G8M�{]Q��s��җf]t;	eк�'`��=�6s�]nv�ռ��ҧ&�npa�їi{ܸ^��ny�v��3�݈x�J��j��7!����8O<���rR�ۺ�R������5Ƒ٪w\����#ӋDr\N�a6����q�]t�cv�nr=�v׊dĻ�thyN��T��:��,	ϻz�s���g8j�!<��/5��3Q[i��7�3q��lKZ�)��y�v����¼gtZ�c�4!�0��`�mV:6�����Bo&���6x�ɻ���՞�a�巌�'�I���[D쭹��pu�.8^8ۖ@L�]�<5�wc�D�{��X9@Ipur)��r[��z�]��8ͺ�Wl�5�x��M�6#v��R��q]4󑇋J���E�^�0��E�
{qe.�{q�p�rXF�v8�g[Zѫ�ky8��=Q.�R��v���՞ȷ7W���S�Xu��]`|�&9�ˣf%� nu׃�����p���]��Y̚.#�1�+��E�Oq�{��7�ŋ�P�`-n��\�8���&��Y���Kr��tۍ9J��s�k���\�{FH	���F-R����W;a�;q��Z�sΪ�Fݝ��v\r�8�8�vɌqq�g��.���q�^��q��p�1beF�ٽ4M�E2�օ��.:і���β"��fܸ�L�th��ۜ����6���	�8۪��ۗ���v����Wjz�mp��S��q�;�![������햠�v��vՀ��W�P =��T�Ηխ?\g~S}���+��*�݃b�\�l@wk��k�I����yľ���č�B�Ry)�]�RU�.����d��6�K ��Z30t��n�!w�p�d�m篾7� ����ACh#��6��͛��7���|�^H�����JE��W��O�K��fˢ��Y� ��3Gg�T�| ���q6��կG 
��i ϧ���B���/]��~��#T���D��V��ik�h�=wU��.�7�sk���s�ފ��~�����V
9c�=����/%J� ϧ�ho���4fT?���~^Z�>������
N_oW��٦_���&������`�Qj�W\FE(�X�P �lB��絤y�w�OTY�r�,�2Ɛ���(�>�۰7Lz����H�I���0�t�ަI�y3L����=�%x r��]�6/U�䪐 p��@�^Rr�l.�K�g���|;�-�]�L��JWUT.�]Z����3O�KaVUN?n`�H'˶S$�|�p��u2p'>I��]]Z�˫"������@�϶��bs�
��|(q�ئ�:��k���y�Z6\A�a�v�<�W��Ӯy��͞i�����}����@�&���d��w����|{y�$.��6����<r辽˞c�����"���B��*����v�|I���[�����I3��� �Κ��<v��p���\��T�Py��p�)U�$�"�F�k����~"����f�>��{b;]�N�ij�c6�r����s��pC}��1��CB��H6e��eB�ޯ=�ġ�On�1�27&U�7pK�������&w�X_�����J�]�wb�S���95����S��dks�� �I���>��I2�v�m'�~�M�~�1D8�V2��`�~5��B�=3sd���;�A�޶	�f�}���0f��{;\Y�}�|�o�Ϻ�Լ󫱺����i��:7G�m�yu�n�4���<�[���{����y�8���� �����nv1]�oxo^�.��T�m&�e�]���N0L���ez=�|��1�Uɯ��}�)no}��(y�0�6�f`&�����O�]T����°Q7��ȴ���H >;� ˶���Vɏoē�vof	;}�j��'�匐�
�JI���k��m]xB�{�@#�ݏ ��������O��_��6�͇��^��^���W$6闬��qld�,Jxu�oM�}�4�v�PU��As��uԽe�a�������>̟�Ͼ���?f��B��J�=���۾Kg���cMd�r@Mov?��w�b��iq�FgQ��fț�N}<Z��L�pnz�O��\��j8��fR��l*wT�U����޻ə�$�^� |)��(F��^d^w�ߖ�� _{���(St)�S�"n�qB\�(��׻|ƂI���$�w��� ��=�8=�\?=D�8��Zp���L�#��$=��`�\��s5�����ouݧ�m�w�B�~����%���b��b�s�;��7[T#�i
��9����7�.c%�vP��N�ɟao��yY��������2	מ�X�l�z?;�L�I{�lO^w���(�\���4N�1��B�P��y2�M����&��Fp#����c4��s~n��&��6��t�y��h�F���d!훭�np�v������=�]cv�����x��I��kv���N�|X��tD��^�K�n}�iͰ:�V�N;\k�㵃WG��� Ou���n�wC3��j�Y�6�=�{`�n4�Q�x��۴g��^C�`{�睲���4��/b;<��5�{ ݽX�_X�P�
�6���&����n�n97\�q�!R�՜/*$9
��S���6�jњ��׍��k�Ӣޫ�h5�<�A�#8�f�s���9 ����H8�J��T������O6A �^w��u���_|i��ψ2w��{����Z)"�m�"�}h����6�\x�����=l^w���3Z{N�u�}mV߆���@#.��˥I�ӝ�A;b�a��D��g��d�[#�;�d��Hٺ ���������wwf�x�h �z%B�y�F���l]J�e�O�,ɟd%VER5��1�Oă띙�-�7�����lA"]�ݶ�O'��\��L��uG��\���y��n��k�R9y��z1�.��v�B���'0c��O����7g±t͠�;U� <������㫽&,��,�)Z��g���eb/�HF=�����qan��+��]�h�{b,�E�p�$6hB��E�˾ܻ�˺Z���׎��٧o���+���)�k@��\��r�
͗�Ϫ/~�ᕛ�0I���` {�J�u<^�=��r�����BB"	S33
�\����i�{nն�����R�a���UBZ�j��yn�Ȫ�L]�$��O��
��̷{G���@P��IP�T�d1���^2W�(Z�~�f|��4`G5�
���~�UB����PI�g�*7�%T &O$� �f�[��Y+=��"�e�H0u�,���[��[]��6#�x������4����2�}���!*�*���K�pgă띙�����l�u^�ׯ}�H$������"�p�Cs$AwM9�辎"������	\��I'w��I;�%c�pzL
�c��l�eѻ��ǾIP�s��Hu:�@ϢĢ���<����wSm��d*K<)���׆��F�SM�"O���i���ļ����՚�M��]^�i���W�� ���'�����IO3�ʮ엱!!�&f}7���j�(
����T(S~���?o�8�z�x����٘3r#UJ�]�$��Y����� ��sϏ��������Y��|I'�%���y�;���.���~X5��OIl�Be�j�{@�n]sq��)֫u�6��l�,e�������5�l>���_ >�=� �����y�9��y)��� ψ2{�1b�{>"�J���k3�]���A�d�es�`�^w����-�H+�y�'��)\g=���dL��۪&�v��#ݜ�?����IcX������q?2Ia�^�g����Y�_֑��=|����m����`$�'0�'�@]ϳ ���Y�U�M݄uew^V�N�gc��̰����Z#�sr���cZ��宥�h�Fwf��������++��|�\+J�����$���X�λ�i�ީ�BB�s3	_�k��s�Ji܂��T�em��0v_n�v7�|���ՙ��7m��<zź�
�]�j���[�4�1�]����-�\3��AW� "#�ˁ�#7�t�r)�Wy�0�#e��=|J�5�`k�|)oz�$�?fS�$�6lP*��`��� ��g�U��Y�>�����{bTz�p`&i�3
Uz��S��Ƙ$(��l��ȪF�y����ʝ��O��Y"��u��/Ў�����A �{����>$n4
1���/܍����� 7�j� �����l��^gjPZ�����t}��������Th:n��TW�89�������0~�/�6NگK\=G��^z�����o�7��cͿV&�k��y�S{0��p�;ts4N���Z���jQ^��D&�^���#�HX�y�{+]~����?���s^ݤ�ϥ��kn�7n�\�7l�z�1��:��ڷc�b��p^�uW��&��2ȉ�A�1��c��qn��Gxz��t�غ�5�g)�&�����q���r]���N���<�<����x��ֵlu���k��sv|$��B�i��s���eq��cs&Z�`^��M�<�A��Ɨ�2��Df���넋�n8�	����ǒ��\iln�+c���Go��coc�����ϻ������w,�i|��s�({fxm���Fv[���wm����e_ӹ�D\9p2$k0r���U5���{V��I=S�� �~�/�N�{T�ָG��>����XI�lؠU}t=Q����y���$���^Ζ���$��&g�	?s��d�(��I��"����̪�q��4vT��|�y�$�����u��ǇLޱ;�|E�ٟaG�_mЪMڪL�{4��fwm(�.�o.�7^�����s�����`�%��\Z��y����Ϡz�����~Gd���r]N������/l����H������'�!0���9�z��d���'�J����c�����X���FΝ�3?z<�d�Qm�hA[��Bs���"�/8}�1���g��.>��g:��f�i�q�{���ʥ��R�3\�(�s�YF�}κ�*zS;�&'��m]Β��<��I����y�/�$$3�o��8�)���f�e�]��6�߳˚�YpE��k��vv�e]����@| >��_�-�9E3޼ܬO'��A:��0I!u������i6(_]?����}WY���|IwٛT
�� >���t�Լ�C+�\�,Q餃d%VER5��q�>2�faH��q��F&���	%e�� �z=�^'S�g����[A0�C%�
~���z᫧����M]�n�)�����U���߾ǿdU
&�U.{%����xH�@��fav�9M������H.{3���)���RR���}o������q�zX�@%m����z�cs��|}�k����ʵt���UWwA��na �z�f �ܿmNI��H���u���̰��-Ի�D�!�ڛ9u�;Б[z�{E�5�Tm����B^�Ʌ��b>"X��}��%c;a�#�w~��uwm�as�<��?b郾U$3dǭ�u�f�����ݙ���w�5L��5_w(����P���c���ʇmc�3Kޞ	����'r���e���ܘD
�Ի�wW����N^��U�!j���q�ƃ��`S99ᵢʾL1DVnC��o+}M��M�7&�o�-[�.�ba��Hq�1y��y�\Mٻ�.)<�!���r&�Z6@�ț{B���DK�e�rC��lC��d7Vs�8��T�/Iwܥ������<^?=P���啣�z���*���d���l�),�py,����Cm3��g;>W�/���3���:|H@���׷��Mxsfxp�P;���%�ʓS��]��z����ފ����\�i�|�F��׭��X�}�g�ËN�&����s��^�7Kl��J��w�B&��y��9on�/
�׼\Oj�i���o%�e榉2n���J5S����cv�;[C��F�g-4 |���4@n��=�e�+�m�t/��;�5��5�B6n�jfEX��A�n���bP]:�.͛'^���J�9OUچt�AK��ls�K�Kس0�j�u��MF���)��mQl�Wd@8���Dl�ǘ��ò�.M�G��Y���\h%$l!wÊ-H�IZ�N]��Yt�3F��2V��8̈́g� �昋�Y�)��v_�Li�l �TJ
�"� �0QX�:�A2-�nZ��xb.�Q��i(�K��`����j"ƍ���*f�#J*�%�&9K�hɻ.��i���\�-*�L�9��
��e�m*6�Jԙ��TM5k��b��F.Q����Q�,�T,m�S)G5Lިb6Үaq�TED��1ȴh��V1ڪ"��J�QR"�jJDE��6bV�j������l��f`�TV"#4�1G�T7e��(�퀢�-J"#�UF�*cTTV
+�H���b;eAQ�]Z��l�KKl���PcZ�%���EDD�DU-�Z���e��-���"�����;a�ufe�UDVD4�Dc��D��A�TEWT���e�QDUTZ�V��ٷ+r��
�[Z��EթiP�Q"�+���������,X����DE�QQX,J�ITD2��PG[��wh(�]3#Z(�����a[Y�~�HI���g���|>�s|���Ap�Q2�h����
�-e�� �s�I#�٘	�}�`����w��;,��L�%>���Dٱ@������Āo�[7C�g��b=^��s���A ʝ���s��*�r�[U�{f��~��s����bX����g��n��;"���˷�����s�m�4���￟�v�nS3�}�%N�A$�/��3��Ay=�uj��T ��K���"�]0�Cy��M-:$�4�7���;H��$G���k��ݸ	o?�1�!�q��h�0>���ff�V�c�9]�f��I'jv`�{�����&���m��B��.N���?wN��sц	����-S[�`�7�a�VHSsەֲ�2�:ڏ8��-�&��>�=~^�W�5���`�ľV`N�^m�2��(�_Ѷ_�������efڷ��j���[�3(.�q_�� �����ƫna�$�fgē���o�}wl��ޮs-tT�l��7���[g$A�e5��\������S�>�������(A�nѠU}u���#�A��lIR$�����u�w�K�����2�.`Q��"��}�3�2X�݇��n�  �s����� xMz��c.�����h�i�ѱc���{4
 K��>$�����=C�[��@	�K�OT�<${��(�
�͡ky�ܙ���	3u�$�V���G;e������6}�O��{#�y�뻤l�]��A�d��H��paY1�+�?�$mw�* 
�檑ñ�W�Y���u��MK��ޜ�T���J�Ҿ�X��$!o{����~q[�U����o��:�tf%�.7Sw8����Ň��x�e5�9��~����׷y_t��*��{D��ǭ�Nݻ@sI�<�Ԃ//��62�y��	6"�����ԡ��=OU�{�kY��Yyϰv����Z�v��i��v8]ɨ\���5��X�8wtm�n�Ӂ�x�r�Dm��v��Yn+v�g�ے�JǺ�P'?��|�����,N�ݸC�˩}�u���V���gqny�A����� ��V�-���^VC��֨:�t<u���Nݶ����e87m"2v� DJ�����	�����M���c	&9ۘf��]z��d�\��#���>7�A�Ɖ�J�U�����{EB�q�?Y]�j����$mwf`�A�v��A׸��d��خPo�YJ스k0K�3	��ϰ�H-�v5;�xIY� ��S�0�O9���0�Cn��F՚���β�I��څ�C� ��瀃�#��� ��F6��<}dv�}3	��R���lV��;�~���W��,�M�� �I��s>"�ч�C�_X���ߝ}��Y�Y�@�W���%�0�G�n��l[;�5gd�������)��Z;��&fI1ɹ�H��a��Ǎ ��O�RD�
 =�5Hdd��Z7���9�)�3���!�V0�nL����m%�y�[���֣w�����eA�wXw�r8z8�y��4x�f �6H�v��>f��ծ~��~���w�}�}�8���k�qA�<�y\I/��	�a�Ɖ�*�U��\�f��h���ˡ�W���]0i'\ܻM7����7*,�m5,&Z�]�u�E����_�M�R K���=W:5�Ӌ!7��v�<�1�Ɂ�N��+�� 2oj�x$���c�$(}���@�
>�P��-HB����~q�h
�u^�X��H'��[�$�E����bDN@'�@�u��p9B��Lo|�׷�I�� ���0���x��À���	����tb��l��f����gӯ}�h6]A�y�> d��E�ؕAl�����Oo�5���+l�`Xl��r��I]�<�H+"�����f��s��*��f����7j��q����m��[�m�M-�Jf��$Cxdڗ��C�p �W�����������~����_;F���s��[�G28����}t�_g�������Y��#� k���Ds��,�r#��h!?,�����4�E���T�fWI���I�y*Y��3O:J��g��Fv� s��tn�WT�ǫՎ�tQ�j��Zɨ��Zi4�+>ˑ�P�.G-y��Z�|w@V�q�t�PC�\A�<ˍ�6�=�ڶ�����$�\��w�e]z̢�h�K{ʔ�JM0�Bb�9�����N��^h����\�	���	��y��0�o�K��呿tvb��l�eU݌n���~9������%����}�	$�;3�r9J�ɫ*�,�L��>L�=Îg��N�5P�W�rT��~����LQw���ˏu�h��X���B)�G�@�R��NwiK���=���U��c_N��v�eo��U��g�V�2�U��s���k���� X&��f H��_R����_��?O��Vn"��`��q (W��K�M9Ύt��kU�[�͔���)��)q���e�R�S\�<���{f�\Y�Gr�s��|�ădvB�i�OM���O�9ـ` ��q�X\��Z�v�Y�3	�{�jץxd��C�AO+���&vP�J�;U��x~$y��0�{�łOp�OY=N�����C�*a��s�gf`&��G�A;W��>�����F���E�_	���l�eU݇��gA�G0=�؆\�A$���Y ����鎝gP\%��~>�����
��+�b�+4�����ݑ�o+��������
$�v͔�$+�JP�/�7��E���TM��S�+��:�3Tux��g�*Ef�/?;�����]΄Q��Y^�J�3�z���� �/m�t\�Mu���[�Qkը�%���m��\���dY��up���2ɭ�i�㶯d�m��L�H��Vݱ� �^�]�ŶZ����;�䖙��\�������)�nx�m��'F^1���/)��nn�ݮ�ut�,�7oWK;���\ᶝ1���3ځ��<5�s��tF5�)�v�����vv
��٬�M�v�zGd�P�u���k���J���n�8�vb��n�~���w=Vo��C�(��N�i Gܢ����1�oz��2y�`?{�łE
��&�
+�-{��AgZ����7����M�_	'�ݞ�!Ծ�X��|����u�ҵ�^��s����CMj� �s�eA�u�t�k�B�L��(���B{ ���`�de�5ysR���՚7����vLω"�vu=¶����޶X����ݓeP��yyZ�o��{ܒ���� �%����d�$�rvf>Z�V7~n��IK���۝6�hל�u�;�%�ܻ\[��7l�۔o�("o�>�蘕*`rA��n1�m��@"��y���}�p.��}��`���0-�'+���렧?1Ap��~M<��]TmcG�go�gC4^_%������Ew��~��ۡԮ�U���lﵳ��z4t��Aui�cZb�O��B����Ҋ�����Pu�︕���-z�`7~��i
U�����
ŕH�g�$��� oӳhn�\_����B�q	g9�>�~��0�3�@��62��Om�_��)k�.�A�n<�~�Ǆ�����N՛.�q�$��W
5F�v��`>��J������W����i
t����HA���H}��˝��� ǎfr�~�N�@^�x�4�B�`7cU�0(E88y{n{q�:O�"I$����̷,�*b&%u��ڶ(g��R
�K�к{�x�c2�b��$���y�9QʫV.�J�0r����2Mu�~ů�c�[K�7�<+F��a�Lr�i�
�]�f���}�/�?ҹ�4	�������n۬FvU��>�mӶ��/(�� ��k`t�|W,���vn�Tf^�Q��$�d���+��Z�~����������J���xh�0F h�ȽUݓ�s�$��`�	��,����2u�4�s���A�&g�~=x��le�]��<��@���ߚ.��em<�$�k�·�>��D��Wo3���
W?..��ۂ�1w�8@��m�V��v����+����s�tK7���}�����F\���E����� >>�I�1*��ǋGFn���fH��C�Ī�*��ua��&fA�����7<A���@����
�}�
��^��W��>���YRe��c%+~�<��3�=��-.�vi����k���K��C%w{3	���F�V��렧?e�n�t���,�� 5��>��iP��bڸs(bU~��g�W�3j�܋$%���J�SJ\1����z:p&���ʤt�u�@�@Q���A�;��f�:�7s�@$'��Ms�u�.���$�@�U#X��pEz~��=[��6ȷ�xX$�٘	���v����ڲ�������1��q0#�.D��"��K-�-���<�/qģ?�}�m�q&�5K�L�Y%t��?�w��z�������{�0~��ࠤ��������}t��y�L��D�_�l|�%@|*�*e��dpvE����;�&�U�t��1�����~7:D� /����d��Q�@�tI| 2{�Rʼl+�9YYg	�H^����ǞyO_j�,Rw1���{>Ϟ�����#���̾������E�!,��je��T�6z�;��In_E%u+kʕ��3������z���v��a�ޟY�F=��J�҉�pb$��.��t�cvv�
)�e(8	�mu�� S�jB�#s,�6,�z�Y��3P��s��ȢM�ch�C��)s�!9�9�X=i��༒F�w�VC-�c�1��T�`������q9��Uzsb�3�)Gwc����چo��<�89)�^�S|��w
2�C&dYSf�t�1�d��Gvn
�E��0N���X2�]
�q<F.J��j�ԋlff�֏](��1��Ϯ���o��3�	��FϽ7`�・4L|���d�wS���,�˼{Xnh����O��뒟��Cw{����/m@�C�uZEu���je�6xh���UK~a�%�˷=Z"���9�_	G5X�z�)c�޼�ԋ���a�[�+�{9�=	��I�x�/2���/�ޡ�m�ad��gW�֤��������v�B���6�j��㺶�,��y�3�:?+;��,6�{ >6��ɳ�^پ�k��ǾY�Q����٣tb�J��3E���֖��k�Dnᇂ�}��ܽr��������z�{�������my=��	��=�Kgi�qm�Tf�>:cۘCU�����Wճ� ����%l[<U�0���H����Oy�s�~.��ȪR]E��h��� ��+"�<�.7�(���DҞ#w\��v��b�]B���.3v!:�]�/6�x�,d�C�q�Q��<��<�o�c�C�{]yš*�	����j�c%��o��-4�r��UN�EQ�R�Y/��1ݡ�SL�1E�-Ps�+T[ac"Ժh����QYZ��*��`�EUL������AM6�oUƂ�mbV�k��@���`:J�IA��X-j(������]R���q�1E�jV*���4t��V&R��EA�E�AU`��:-Vi,ESU��%����4�&%L]�(i�M�����`fUV;��3F �K�+�AV(�b��+F5�M[�(�#��F%IET+TUT&���*��Y�Ե��QX�LӌUPPPբ�����UX�(�r�PF%��+1`#T��X[ETER
�G-X5��b(���E�QE��L����Ŗ5����%������U�EH��-���*AE��]\�.g�T�{6�]��[[���s���o��W �흃��GB�0HWg����ur'Y�>�O>`S�c>7+cyۡ�N�ϓ=��&���)�������ۥ6�ưsm�Ls��e`�!٢�c<�n\s��g�H���d���mŜe�O�`N�l����۵�<G9��V8{<�<�ޞn�N�_=��#�m���Rl�H����	϶��.�c��K�LǶ6�a6��6h��8�G:��ː�<`�V5B]�0j6NSk��s����%��[�F';�x����%�U�q�m\�eywE�N�|s����{�:�u�:��s�r�o<��I�u����C�h�v.�]k0���1���%�_9����n���!��bvx,��۲ulL�!<a�ܺǍ�#Ƕ�mtp�;sz�zנ��sѽVT����7a�!���C<�]�,u��qnݵn��ͷnɹm�O<vg�����.��q���/;]��ݧ�����N�/|Oko��v�uO`.70޳1*�l]t��M��x�pÉ������s�7!y<79�Ίk�l���(�v�����u/5��|v�\��q��>ݪ6B��M�k����s�$��s�{<L���lu�<7�2���RvMڑN��%����\�[��	��ݫ��g�K��N�����e��lX�li�$���]�����-��|#�� hn�tU�w��V��e��0C��q���n�ml�X�;�A�.��	n>g%����I^'���7gn<��-�����a�E�b�]#*s�W'2t�A���6�����F;f�F�6���/Ϗ�|r�;l],3�k<ro]��6A��ׂ�:�l;��K�F�7<\�7��[{v)$���ζL]r�T�v8u���v/Skۮ��qvǋ��vy�lOS������i��e7�.��]Q$V�[uգtb8z�ԙ��&�/]\h�#�9�x���x�ng���[���j��p�R��?���w�޾3�����������y�nUn3#�{vG���D
p^�V��cV�h�9Kc���l���v�X3��ֆ@�kg�Y�r��F�{0��h�m�v=�J�{���=���]��]�t��d㇍ոuڥ�sq���Ht�<V.��0u��{Y����ᮌ�����ۗ�5�=��e{t$�Avr�#v$:4BS�i�[\�10^�v&�]�'��Y���ˣ�6�[�T7�K�6��k��܇~$�@�*��������<�{0� ���~���<�(1��M@ ;gzշ��x�HHq'���Cyuנ���EK֞����营=~՞$c^�9�����~٣�p���B����/�٘HΕ$��]s�Wnn۹���I����3�|X&v\UWd�#V-+��-+}�׺Ɗ ^) �g ��aN�B�
��ԕRM�l,�9V*��T�B?
�9�����p��Kt-����$�<7��)䟰����t�uzbZ��p� B���7��g���Lt����r��'[�;S�>�������߱�
$���9<���m��GP�o��7�Tb�ų�}}R�g��@.�����RxP*W�߭��^�����Y�]�4��z����зz=�ҥ�b�\��:��8�֨g�v�l����WVA�1���q]��M�;���!$&�y���?}�]���}�(�W^k&:&8yS�mƴ���$$8���c���|>�_  �����z�w����P�� ��B{`�ɼ�k3(e�/,��n��\#-o�t ��T�
����ʸ��D}:G
�n|DL�HD��+;s�鹕T{������s��S��\���K�v�]U{��~�oO��j���=�+u!n7g�uɻ��GN�j9�����;i2���u����;�E�)����Y�����瀒/Ӽ��p����[j|��~�o�ٔT|
$���)�u��}��5M{��v��B��� ����s#ѕ6��ZjZ�B���ʠ��w���;��IG>����]�㹤�A ��a��`YL�u��{�8��p���C9&�ڕo��=��*�l�L�h���Nx�����|¹����m���M�o�U�����$%�Η��R�� A|�F0�/��/��`����Nr��L�Ds �o%��z����
�
�0ǝ�0�g�w�m���0*���@P1��T(`����>
вQ�ō�ƋIp�%b@�F������+��nK�님��c��H�����군�`��c����rO`�	$߻��j{�GGwl�3*�rf`���"�qVf����ݤ*�����\}��G���|7��f|H$�ζ	��'��+%דiOL���P�$D}1N=]�V�M��s�d�_�8�ot�^{0@	7��`�;٠�Ut0�7��W}=��뻎ǅd�W �i|� *v�6��1s��8U%�_�VW����=q{U����Rx�u���K��*׌uUrF*��+��
���ԡˮ��w�+�o��?I$�;��7�����}���Uuq̻��͐H.{c�亭���m]�f|Io�hP�\���="��:۬$����G�����tr���xBx�O: {]�N@/phd��w�ƨ��(��~�˵m��s���$��w�>6�V9�L6�H3�Xs�����F�X&����lh"t˶)[�y��|ƂL��`^N��A�:%c�Hqs_���*���i����0�筐{;�$m���2O^z	��� �������L�B��UTE�5s��{�h�A���$���$];�*��\u>���)�j���
�*��Ϯ��`�����#z���Nml�`�Hs{ـ�~5��?WWu�ܤpAV˻�՚�ʱƒ�gg�J�J���/+k�{��P�-%u>�Mh}B^��ʭ�P@��k �Yv��:ƺ�{�jr��ww�������۫tkZ]6:Zn�v8&���#�#|��9��l�C����r3��]�m�̽��'��m�m�U��ܚ&|������zN��(�<�q
��N����g(��sa!�s�z��z-Oq{9ڼO�/6����Hs��ծQi�:[k1���ONyέ�K=(`��݀h�l�\�F}	�ꎹ^e�c+�2Fh���lR8��۵vٲv�p�כb�N�r�$ cD�.8mo&}���~��=���6��F���a�K�y��];ن�J|��(o����AI��C����%1�ca5nt������%��_{[$=��	5'{0	y���οU�o�]�E��/V�&��
����0�A�� �l�J�}�~!���&�9�2.��̫�p������ƚ�2'7s^|OăRw�~3ݷ;G|fn�M��fݶ��FSP(N`�Pn��~~$'k�=�ɾ�:�^e��VN�'�MI���g�m��E�TC�����Z-��]���u�T� ��{g�v�n�a��!6�G5��>Br �q���ݦ5'y�'�L�m��\����6��V{�M�㻽j�/?�%�$8���W۞�}(C\��_��GR�vR�����YM� rOTػ;�bx4�C��w4xF�zBR��	��H�q�;���������¨.}���r+�ﻭ�MBd��ݗݳ3�^��W�X*�ث��|�H�5�Oz��*�a�v�^�{0'M�?Nv�����X�pemNm#s֪�Z6�?��M
���`�𼝹sٌP�ك�����.d(VUՋ�AYUY��ی3����4�}�=/���TH
���o­w��ڱw-�G�?��p���m�����!<��ת�n���QoJ��6�
X���n������Ȓn�P�t׼0�v��$�+'na��$�}oАc~��;�x����2����{��(*��@P]-MjvL���lEd����i2U%�u<6�o�hq��_��j�Rf��}9�(tq۠��/�%�TZi]���س��̋����]84Ν�6Gu�Y���"���4�\ޡ�(�/��WZ�q]�6��~  _f�����m?�"�~��@}�#PU`��WY��㒟�Nu�������I W����{۬Y��=�0h&��S'��K����X�T,d���H��=��r⽘>�����w[@�4�������^Q�豳��J�,��*��s���Ws�d.�;s�w��yyӧk����v���ǳp8�@j�yyC*��n��L^� .y�>7=�xfu�%]v�t+gk�O���)f<i�A��^������z�h���~
on`���7���`&�[:��H��O����vn���W�1| C'z*@�X
��/|�z��@�s	${;ل��>K��n�U&��I^���(�س�P�;ڀ���K��~������~�"DC1u�ޖ�A��Y4u��A��ܣ�U��C�𺈄�7p�^U���/���,ӧVn�������_�6��0��~�5���4�]�����0�6Rz�VD�3��M律�y{z�&�X���ӥ���7��.��+n�l,��v}�`�qXyp�(�s�w`B����"��>�~���g9�vnfa �O<$/oS ����a�:�H���![��ի��VU�1���jSâ�[�$@Vt� ������niW}jh�L}���v�UU"-Z�3Rg�	'����
6�'�����m��(P�EJ�;��C���B��#O@�����Л�ߦ�sT*��z���/'�F�umG�G���o�a��%�X7T*� �]ɒj{#���������X�`$o��a$��`�ɜ�F6h���Wf:��)���f�_p���}mE�Z`pY[q�ތF/v�zR�!/�+f�L����
�"�߃J-M��!��� g_N��k`�kZˆ����Y�Ed0�*�{<���|~?���p���&�u��#��ڎW�y5��'n9�퇉i���Cx.p�7m�+�pe�1t�ݶ��n�8�]\�3�tu��;v�Q��8�_��<u�qgA�=Q׏3�֎6�n՘�]�ط];e��Oc%Vqy������u��;���19��/l^td���0��:�p:��O|�7|�>.�,�6�n.יsmv�k�>���Ǻ	�������٭	]ys�"Q*C�S�M����y*���W)�7v�4���_&��S�R����|�/�V{<$@1���� ��5�Z��Vq�wwsQ�w���@j�]X6(�*��|�����`$�^�>�&V���I�uw��k'n��[WwdP�]�i�;�9�	ݲ	$V��0���x*g(r�+�2~���DDݛ�kN�BM�w�a��1cޜ{]=L��;�0�O����3"b=8�{�+�<>�D�A�ܓg�YJ�ƞ�sլM-�3Og�Qыp;����ￛ�{q��
�6���~5ޚ�I"���8qUǪ+_ -���+zB/�����Rj�I�p0��wRӷh>֬�9W�g[�;ua�YND �Ӿ:�3sk5�zY�"��ʒ�nm'}hr��ɉ	{�;�
�W���+� ����A ԓ^A��{>�~(S�\�;յ7�0H�\���9 &~ji,컴�ݹ����%�:Ėc�zyi@Ui��@C�����(VUՃb�����r����~�H>�x�M�w�~�Wj���ρ!F��	��E��U� �����T>��x���c�m�$�B��t����x��R�eɈ�����䟉�6wbm�M�t�mϞ[�tq��]+�=�.|���Xk���=DDݛ�jp����Rw���|�3����3��������?�
[�@�N�ɽs~{�Oo��pI��ل�Oz�S�� ��b��O��Џ`�y��ʼ��M^J��
�=��B}+[0X�Az�TMxu"�)��`��<�3���4��;�C�q��-N��������	�F���g�u���O8�X��Rj�egL�����)�ϵ��u:�++:�&Ӡ��c|�N��02v�
��:��YT�����6NCṗ�֧)�;�:'L��j)��������5^ ��5a�ޜ<�w�{���*�g�Z�6sxu�ř[��i0��{5�<���������]Ѿ���c��-{ωף��6���HR�bI�A�5�;*�}Õ�DX5������V��9��}懰g�^��]ރ�/�C{F��6N�oh1�/emvorw��5o�Iw6�͓}���.{����{Nk�^洐z�gS��ym��%6H�峆��l��]ݎ��]�1���0_n��Ʀ��R���w��5
��`�a��lu<�cM�!h.'���Z��CC�>��y��M��w+ZK�Nj����$���ٜ�����#�u��]f��|�8�N]��Yyj�hw;�v;r=6����G�ڙ�/w�"���rm�Ӕ6v�MG٦��At_s2�~����k�q�TV����:�]��ֹB c��E@\�J��a�v]h��,����"wo(1r�����k�Tv��*��`)۝�4��h'X�b�;��>�h�Տo�<�GD>��g,��̓�'z�f�)�w4-�!�ҭ�L�.j��(���9�i�/\�߮�r�n�
���f@ǵ�݋��U�3�z��������低yZ�����7u��6gnN"�?ZVUE�Ƶ"����faYX��*���Qb�cT��e`�E+XQ? VE,�Z�j��D��QEV#4�LKA`f 1kH(��i��dĪ�ċ�1AE"�$X1���L���2��,-l*�71J�,Z��J��3)E�C-4��b* c%Ab�VB�Pի
�`���l��+%J�²���E��mTP+(�4�4�ҡX)&��VT%kQ��Q�Z��Q"�E���PP����(0��" �h����-��ch�0�r�M$1�ĕ��+>$>��|A �~���I�~�v�H��Z�0�M�Y��u�`�����
(w�5HP T��;@^^ӺM�Y�2+T'�����\LJr��dE�N�˨`�k{9�-��S�L�^y�@���3�x�5�ڋ����Fn�*��Ç B��wc:�i���[M��p�p�vzSػ"x��لo�������*!]�M���g�@$�v�D�K���7ؗ�lfp5CI/�>�@T�DA*��	�o�����`D<���0�H﫼�'�k;;3�Kg+}G�ѵa����y��)n`Q>���I�21�mܞ�j�W�]=�{�<�?+;;0���FY&��*��WX5�yx=x��s�|E����vL�	��V�z��z��Tn��9��C�U��5m�V1}M��E����ec�տ?�I�͔�ut�-�,�?�(f�*��������z�`��Ö�ﾯ����W;�w���(�M�Y��n���>~�[�,��X��9@i��P���D��A[;�3e�Jm^�K��Vj� �UU���u���θ�^�V�ݶ�z^��N8;b��ݮ!o�QU]b����布5�9� �_z%B>s�~[��鳽~�~��_ͣ��:QPɖ��G���]1>��{;}�=�pX�LR�[��P /�R�fTث�ơ>�b(�D��*�~���@��HP�)o�%��ڙW=�����@[� (ދ�� 
4jɺB����b�ž��'��{瀂 =ފ��z_�X;6���~I*�7a��`��%Uv*����>�y����φ�|�cp�w{3�;��L��UǴm����F�nN1��q$����!����UwN��]A��LP^�g	5�,=Nm�a[Y�ҝ�t�]sN��ox?��<�9��p��Zf�\ݵqф�)wgFe��u�ϟ��qn�^[��yq{v���D��0ڽ�vy��UJ�������=`�>B.7e;9HH�y:�s�T��uwC�\�v^���6t>����t
f��=G���v��î#NV�YM����X��^��3�Ys�tz�ٲv�����kq:B�GGn����#48�.m�&���9>\Ӵ��3�8z}]Z�[�rl�of�����<��%+���H��������$�	P�E�=��I �<��;��kk�f�!�OW�x���� 
��"�U��YV(�*�3���O��]G��g�����I�����~'�ޮ�`�S���YެOI�D!C&Znc\o_�$t]�(��;��OowEZ%m_C�޻M6���)��]?XƠRɁ��}<�y�R鶲�7��P TSe	Y�ؐu�/e���fhC#�"l��*�<\���IRdy�����֙n���}�|��L������簓�p�r�I!9j\�%)����>��^��΃����{^�ъ����}�޻T��3����|{c���ۙ��5Dn�x|���gUy�]�{|yv�
�.�"�U��~��3 �/!��6��ˍ/H<ĕs�z�d+��k�AS�r_;֞�.nK�;-�������6U��+�jJ-0Ӽ�^�o2�>�}����?�	�y~��� ��ۘE{B춣��w�y�Cb�6�Y�r��V�� ��� 0�����Ay|��|3�-�J����)��A
*�n�7<��A<Z+�n-�(VM���{�U���.7�T��i��t�mZ�}c�XWHڬW���w�+��ثN�]+��A{m@z4��?z%�J�ӱ�fo�۷��fɷA�k7^z�n]�۝c���wVL�ۮ}��(�JFL��X�mp��rj�y�H5=5�$�M�w�^��Ӹ{�G��P�4���A:��2ɻ��iK�!��v�3y:�{4 -�=@Q&�w� �|�~�4��6��V���,R�/�᝙�0�~���X�/�QZ-�o֮�,���[n�۞f[��i`]��G߭m'Q_�j�+ݽ�Ni�N<���w�ʐ3�u�n�y�\+��B9�y��.w�{�*k�����[k���r��d��j�.Lw��N��T �X�� ( �鏬)����e���{&a?Z�J,U�+�	�`�v{0�*{�w:i�q^��1o�3��~_�駒,�a=�S����1��0
i���ٺ��4�vc����6���DG�|�vc-����}������&����S��U��o;:X2�r��ԅ˭�fE��fC����VM�I�}9��ۖ*nz�f[~ �	�w{0	;���'������㸟m�.C���wIUY���fvf	I��� �ZUz������H\���I{z�}�*]���J�������{t,�U� (6��T���Ew���U����/5 ��؁S�?c�:5��u��RR
ӳ48����v�:����czg]�y�r�d��U|~��~W_�i�!�,��k��i4f��_͟h�q�=9*�E�f�� މ
�Q|�*���3�Å.�S�:�P��.a��5��q�R�֪x8����������A}J�j��[���A��$,�����|l�`�}�;��@#rK�m?$�گ��6�Ύ�Uz��H�s�� ̝1Y;ـ��b�׷�)*���M'�k2[�AI59�M��t�@���C�y�EP������މP��:���2���˴����dΙK7�P�n,�B��D��
=�_!�����o������`�����~aX�po�IPC;�&�߮�M���򞘾���{�_@�藨xC�����CzG�M�Q����aJ�]�7�D�e#��ʝ n�1sUӴ1f�=LLCi�/�pק���4���&�Ʒ��w����?�p}��p���q�Pi1tL����.�zrsݯ$l�@^H{I��8�u����ѱ�7�%<� f��T���� 'pv�D>�-;Y�ݻn+�N�6w]w[�n���X曞M��9��K��&�琶u�Ʋݩ�0m�g�ݯ&�B��.Z�nF��1����\�;��њ3��M�mWm�М��P�F�w:���]ɛ���̉���Bl�0ýu��9�s���Ɣ�/k�Jq��3�ǳl�������R0� a9s�ok�s��� �'z%�kN�����^��(
���s&�AF�j��g�a*fV��֏{H���(�I�(���B��{6�^:[�>'�Zq.�}u`٬�s�*����*�N����*]e�佐
'�K�B�N�J���J��j�}Ru\���s���r��	7#�ω$�.N�$��ھ/�|H�n��K�}P"�U�T��V�?a'�'�0���'g���G��I��h(��$?Oр:v�m!Z!{���o9�~?}O��1�F/,�V�)��F|A`�Be�\��ۂ�f���b��S<��k���?�Ͽy��=vWO@�|$��{ݝN��2VQ�����6tI�*J������na�¤�}�;��k�<@�����$OVJ2����6N�u�{��w+��]Ŭ%������J�v���ݬ��/�
_���%v�������\-��+�J�?��K��/N�͝Π��|��穷�#\1�;�'��#�.�-WjV��������<��;���)
�h��w��y�:�*Q�{��p�8�P�*����^�\���߾���������¹Mi9��aS^{�6�Ad��=���3��@���������)߸a~�(��	������A��j����6�R�O/�U�Ճf��o���;�1�f�B�e�g@�62VQ��}���;u
���+
_|��Cl8¤�T�&���l�%羞����ﵿb�YY+*o�����G���.�YL��X:��<HP��-~��9�B�0��<����}����R�V�{��pd�Q%B�����:ì+�s^�|�t�O'�:��� ���t(��eP�.�J�@�untj��Ӛ�G"p�>[���-������b94�g�?0��*y��݇`�RQ
�FV�{��N�J�����8�X,�~�Ӽ���|?$/�0�:�������oK�~ٞ楚2��p�'������YFJ�;�/����s�9���y'S�o�l�$�%aXV���9��¤�%M�߼�Ԃϟ�>#��u�s�#���
b���:����ʮ��p��`���w�9i
Z�{��9�B��Z
�k�����'��F 1j=6�3`���g�/3�%�3K���{�����RL�Ͳ��XzQw�/3��S�o.On����W�O���;��>O�
�YR���ng*$�T7���Ԃ÷~�q�W)�J�!�5���a�Ǿ_��ס���VJ����ݜg)R
����8u �:5!e��}��}�;��kw��.�~ ��^}��x
��|x�)�\4�N�S�&�����t@��%e��7�y��N������	Ԃ�����l;T����|�͝d���YY(ʛ���l k_z��}�f���f���q-p���N��ӹ6,\�k���^�;T��n�x�Q�~��~m�ݎ-��>1��5���}��x����7�����)
�l`T����p�P*p�������}�_=y���/������D�
�����:ñ�aN}�|�]e3Zn���C�:§����u�G��9�|�c�&�?��83��e@�J�w�yì�XjB�o��y�;;O�_!�G&=��~y�ks����Ϗ�"P�|ٞ楚2�jp�y�{ݝN�VX�YY*kϽ�gD�B�+V��~O/����ߵ��y���F%����6q �u�����������9�O�ö��Uպ�H,{�l;�-Z���{�z~��|�_ W�}�������{� �t@��K�߼~���0�=x�O��c���.Vn;}�i�Ox��mP���}#�l����t�_,��N��W@���(ޙ���<ͻ������6�T~����0�
��y�)�0�SF��Cl9T����a؇R
A`����9�K�Z��������e@�*o�~��F�+R�^}����AH,���᷌
�����R��g�B��!tj�ȲUб]]�\�l\𽮡��uN��7'K�t�wkO����7��֮sC�_�o��l�|�YY++%My��l�N��aK�߼�6Ò�#���wQ~��� �>�s������ed�����͓��S��<].���1������<H[Hky|�>��΁~�~��i
�Z��f���8S��R��Ŀ����l�%B��ҽU��c�ܵ,��Ա���C���=5n%ѫ�fg!�aS����:u �X����|��q���J���/J��ǳ'����^c�!�|�
}ݴgi��_���ᴂ�9��3��_X�E_� d`#�ۺƐ��{�aI=���@�td��%Mo�;��N�����}�!�aRQ
�����8ɼ8����7��=R
k�y�v'P)�x����ʮ��p��`���v$,��-��͜�!_��o���l��~@��)�~��Ԃ�+*_~���l�%B�*o�}�ΰ�aX0��}ߣ2ފ0��_�X�O����c�&+S/�ONq��.<,�u�+:һ��k�zRA��,u���ɓfQ8%\ڕ-f5�`�.4��nC���O�����0�����'u���Ar�1��Xܔ^n=\�n���&��rŀ�����cy��|7�_}:r'&��+��&�W�Ѓ4��9�p���)=��Q�y0�t�1��}u��^���۾����A����4yM��>�y�����L��,���׶��U+Dٱ�r��Y�i�����j����T`�W�j�~�둉��Dyx��BFq���Ȅ��T
��-Vt��/K�&��/�i��,Z�PA�l��fX�}{I��ס7��+��=��^����i�����Y0��Q��j�+@욣�Sd|��.���V��|":���SkV��>8ȋ���A�㊪c�z{E��-��x-���4	�t�z6��O�:+�|��E_,���ׂ��y�{�?X���yI�o��Ѵu����˴�1�t�_�8���Yz.f�Y}e����|#�˕���}�p�����*.�Xz3^���'gf9ϕ>��-���{e��5�8�M۝�2�R�E��u�/6�����ә�.��2�oS����of7Ոh[\:�:\�������ews]�	ər��+O�i��5.��3F��������7�ɕ���EA�[/��k��S���/:w��N��g�U�R0<�3��݉�@`.��dϱ�v�����p����C/<|���+���C}9�����v�ֺW�'D�Ȉz����1Mer���FA`�Ȣ�5 �IY�+%cl�H�]$�$\HV���1Փ�`��ť�H�Y
�J(�ªALJ�eJ��B�u30�5��A��Ku��֪�)�WH
ҖءEd���UP,PAeb��L\LTY�1dSIPQ�
�L�dR(�R�b�4�E��6�m�ZC�T
�����TPE�*��\�b*VV)�+DZ�0�帀�T̲`�� БDf
�\f8�E�U
��J��Q�QH����d�dm���P��B�T�4�CZ�j���edժ��Rl�U%je�f�1
°�bc%�0�"ҥ9B�ְ*�4�DUam���C�r�",Z«ELT�V^�� ���{�حb��<�]�@�Lxf#�^�V�٬�F)4d�k��l�tap�K oXy�[
b�N�����:3�u��ݒ�m����&G�W��b��۞ل���1����H棴����lu���e�㬑��:�ڻV�������;r���Lp{V{���<n=n�󌻈�"n;&���4L�Cgi����Ñ����U=s������8������[���Z��c�����'O`pn�`����l���式k*d��t�[`bQ��&�{	�l���6ې�獞�vTN�#��=���W2�o^ٞ����x�ݸ�=B�N�8θ�������;�����ݲ���m�\<�a^�9�m��2��[݂�zon����-��Ƶr�:���n�V��>;v�llX�<�A�q����;^��PB��oݻ:�����d��e�����ח�����z��)>��xG�\㹻�l�p�����x���p9|�Ac�C�[v��.<Z��0댃Yo&�]�E�XճҼ���[�W�/��S&�&�ϗH�\��@p���].��C�6��t�`N��r�e�[t&n�{F��<f8kv�8�&�
.u� �x0v����/l�N�k'��� p��pnx�mi�.)h�x=�k�sI���Ye��@z��9C��o�|����!�:n��m��e����q��K=� vt^��	c76������񹝳�q�!&�+n�kC�Σsn�`K�d.k7�y�l�MZq��7]�!�r�H��m`��|�Bvݫ=����we�� /�]��`
��k���&�.ۏ磭�����b.�S����&����a��Ęv��dTظnQ;]x����Aԝ���Oc�l���GGe�A�Hݶ���-Ʈg9��f"��)ΰ�n���_��㚹�u�Ѻ�7]�������^*�-�9�n��v��;gi�[��u>�Ǘe�|�*��Z^��{�H�[��
Q��]\�e�F�H��Չt�L��qs��k����u��gq7=���l�Z�S�Az����;6��\���9��ݝ�m��t�����t��n�d�����\S���>�m�tK����%=r\�<�s	X�q^��d��h��Rny�x�f�`C��u����og��g<'-�z��^ntan*ɳZ��v�g���.soc���i�ݮ�x�Q��X�nM���ls���ٌ��߿��.2u�����¦�{�v�H,����y��8�YP*T
���p��`y��o9�g���Hv���}݁��A������g�"�,a�
�B�X6o :�k���ΧP++%c�翽����߿�OS�~�g���Q%ac
������a�%B����}�βu�����_����\�[��u���#��c�� �W�<W����)���߾����!m!m~{�8�^�
�S��w����.�s�����T�}���l��P�J�C}��6u�c
�{o��I*ID_��6����N��p����bAd�2�k�l�g+*�P.���8u�ѩ!KMy��l�����m�=���= �R����6�(s��3�ԳFT�N��O=�{���
�YFJ���|��$��m����|'���_~���0�}��8����FVJ2��{�������ߔ��^��������k>�J�(�v��ݔ�5�k�ݺ�,�l��t%���3u����2����un��������8�!KH(���l�e!Z
�Jk��y�:�Q!�j���'C�~������T,C~���:à°���^-Ը�4�ra��My�|�v!ԕ
�ߟ�������Sq��\�ݬG{?^�~��s8-Kh���$�t�<�����a�7����Q�݇&�h�g9���8���+{g�%y�����|G�2r�t�2Q��@�ߟ}��:���i��y�;;H6����~}�\uy���~����K�|)��t�N�S�Ms�}���@��%ed��=�͝I�*J�Xkӽ��߻�=�/3���m ��&�{��:��T��S_��͓��G�⧅.���1����������*��ɑ����H��?1���
�K~��8S�*e���7�Z�n�ϔ��/�I�=T*�������a�<������֓37$���"IA
�A�������_���������}퟿`Ԃ�R����|���)
�������"��--�O�wڲ��7k�vDO[f���*9}�tW;[�\�\�ϴ�Vw�U�w���}��hʙ��@��9͜O�
��YY*k�}�gD�B��+
�����6Ì*O7�뫧���֯���?'�{��:�Y:ʐS��͓���z���V�.�u�:��X>��w�8ZCﶞ�����}��R�
�K������*Q��}�����J�P�9�����>5�C�y�vq�F�.�8qn��ST\�6ÐaS_}�6�u%B�Pe`���l�g(ʀEUO�{߼W\R���f�"Q��yK/셻��
������wM�����g	I�Tj�+.�[�sKM�y�G��w	\μp��<�����WO�1_PQ�5!KM�����i �}�᷃�;��
f�9�Ӯ�߿{���Ow���t�v2T�s�l�IԂ°�)|��9��¤�&��э?}��{��BZ�$����~D|	?~���:�K���S�YL���X;��$,���{�l�A}?h���s���w�=`T�~ߝ�H)����7���
��P�}�͝a�!��S�~��G<z/��ڄ��\v�Y�북��s��A�������k�뵹6_g��k��տ�U�t:�fg���хO;߻��C�* �~��6q�d��*�}��`tk3ӟh�����yԇ����<�H=�+P�<��᧌
����=�K4eL��N$��vu:�YFJ>��?]���/���Qy&����
���~���*J!RT����:��VJ�ɜ|��g���������|���>�@�����uk��Q�p�Aa�����;HP��-?{��8�^���z�#?e�O��_�������J��{���p�8�P�%B����6u�F��~�8�R殚W9��
��ٴ�>[��T�K���H|'��X~�ۆ�9P(%@���yì��E�$?w���!a�Z�n�%��{���A�%�6���
[YS��9�vu2:�ɸ׵��'��j@��u��\	��)���׸�Ӭ.E޾�s�>s��HV���nH)��r��f�5Mit�u;k��{������~��#G�@�M��g����~�ď��w>�p�AI�*J&w���N��Q���T��~�d�u������������r����j�p���4D�10��n�tmֻj	;^��EʦhTu��Ɂ��Z���⧥.������7{��iih�������`T����p��韹|�o~o�k��S����i���T�߼�Ăá��V�z���֓39��§����tC���y~�?s���an��g��%P(�>��6q�������`w���]s{ٟ�\����q�,��#3�b�U�H�U3S�m8��s��Ԃ�Y�J���|��'P�+
0�<���|ޫ罹����>��a����>���d�ed��7�߼�:�@������uk�i�p��X}{��sz��y�k�$;i]��l�JB�`V�K�}����J�YS���ۆ���������==��x$�Q�����:0�-���.�.kXR��m�Tןw͇bIP��ea����83l�fk<���?]���ҠS����:�X�ߞ����i��1���߫�.��v~&����MA�.C_�����)b�R���G=&����Z����uҎ�����[W]�/�s�=6��˹Z0�>]�{������I�5�Mg�mݞKn�͋�"K*.�m�j������;��)�ع��z��Mֽmi��\�ڞ�����\�E���麹R��\�;�v�E����7�v�ηNgk�y㣱�9�T<vtu9�p=���G��.���8�I�r�x.t㙞 ��m���L/���^�<+��ѲV��Z1V�.�֋�18���qcc��Shc&�)D��\1���&zݪ¦\�/�n�e�ߦ��x��a�.���y��� T��S~}��:��T���+�}��CL8¤����{���'��w�d�ed�+%S}����?/��t��fp��w�~�r���{��^]i߿<����� ���%��N���
�YS���ۆ��J�IP�ϝw���5,�~�.-!����9sNCC�&fra�=�߻��R
Ab�w����5�m|�I_{m����,�j�A`~jB�o߾�`t;H6��<�~�p��0*Y�~ٟf������i�'}�;���?{�?~��~Y+(�S�~�݁�:$�,aXS���܆�paRT*J��}���O����_�f2q�������v:s~���i�kX��8u ���}�~v�R�3����Ρ�G�ۍ������x�!ߟ���P*T
ʟg߾�4�%H(XҎ��R����C�M_��2��`~�1����z��Q{[�k�z9��O��^�uR���3G|��O�f��}���M~��l$�d�+/�����d��J�L���u ���k����$?Zw��@p� ��}�w��I8k���S.�XkK�\��I�{��:�_��#蠂�y^74"A:�(���m������Q��i��b{6���|6��&�АjLMв���&6ܭ��f�C,�9|Ip��㏿�W�Ͼ������$�IXV�?����i��IP�*g�~���N��Q��3{z��s9�5�x���4Obq��������)��_��a㴅����g�{��C�����"$�3�'�\�wy�O*T
ʞg?}�i�d�X�i	���K�7����>r��Q�u�XT��~�j��/��{�}�B��
�`����pf�+*A@�w�����R
ANy��^���~��7��ў_?�B�CY��nx��Ny���4Xᘙ��6�I�����v VVJ�2T�}��I�;����xk���s�~H,;5��܆�q�IP�*g��{���Y++%S�}�������������?W���&'3>pܹrI.7
9�ƻ����Mx�����g��[�fٯϿ�����۶�����￶v���)h�Δ�h��`T���
k���w�g����o��c?	�=���L��P�%B�g���gXtaX[�wS����N��ra�5�>�r!Ă��2���w�k�ӌ=���>f�+*A@ϼ���$cR-9��hNR�+�9��x9w�۟�?���~%
WZ�Z]:�@�9��8���d���9��h�N!D���+�;������#��ߝ�� w�fd4t-�=��)�X�-�= �R[�7�I�G����k=��Bg>[�Vxf�Re�-?v���;���Bw���:��%B��g�~�gY:2�R2�Xʜ�����
]_����K��g`r5��}����/�FIze��$|@���f�����`T���}�8�� ����}�q��s�;~���~C�%B���߾��aXS�o��V�u���C�:*{߿h8�%ea�=�P�'|��oMj��%@��S����:`PjB�sϾ�H)���{��ǌ
���l���;6�?�B�N`���cC�I\����v��3ۘHùL��M��j��߿��f�3ZO��|$��yݝN������9��h�N!RV0�/�{������D}�����T|���p@&�d���YY(2�=�������3晬Du��`tk�s����B��a9�wϟ���ށ����β
Ad��d7�w�{�6���s��������~��A`��Tޗ+u�F����
g��A�Ib ���~��g(ʤ���[��;�}��c������K�%Z��iϾ�@p� �HV���ڇ0*S�o�.u��Z]:�NĚ��}���������Nt���YY*{�sG�B�*Aag~ﻇpaRQ@~��0����~�y]b�J�>g���h%_��=5���;�R����8���d%�ڳ�=�+C�Å��7������HҲFVJʝ�}�8�@t|�~�[].���1 ���϶#�H� ~�tc4!�E~~��j=��>���������p@�be��{�73��P�%B�7�y��;V�9������f���E2V�Օ�Q��.��:)mV�y�	9g�-�n�����?}���K��3�x��<�|�q$�VJ�=�w��L�P,J���y���������ߎ�_�|?�����&��N�~j�Y1�,��a��߶q�z���=�>�3ZMÌ�ta����ퟓ���dC��F�|��9�s��YS���B�ht����a���~��m�S���������O߬�K��d̾3���r{�Y;���0���5���Xj�9�d����������&3�c0�&<�Ͻ��œ�1Ę�q��}b�
����^o�_�ҷ�Q~*��3++0������6�YP�1��Fc�>�ݟ�~�1�_�v�t�]c�5uj���#�+?bʭ��:^�!!1��xJ���c&L�{|�8Ͳ^�1�Ld�'<��x~d���d��1�;��+3����?y���:�������?]�����ؓ��w����Y�5�ӮCl�u�;�������V~C��1���_h�1�C�����_|��Y��0�w�u�d��:�1&AǞ{�?2~?Y��%�ɘY��w��^	�L_���~�z�,1zJ[~&�V�j��-M�c��Bʒ��
�cl����]G^�Y����쮟K!�9���L�z�<�>&����_���$)LSM��H�.C"�ݶy-�.b8�ϱɮq����79�>�^ݱ��w�;^(�g�[D�us	;t� ;Ib9{T��&�1�m��u�m�jې����#S�<�lc�\�[:u���=E���mne�c��7L�`�-���p�:ܸ���\��0\�m��a԰������Y �6�홮L!u�Me���`�+S��'fĄ��ۣ��p�u��q<)[�.(�
�Y�k��r�8�o���ߧ����)��O�����gY�JΙd�a�Ly��{������D��d���u��Y�������������9~��f�+*f3�c��}���?D��a����35n��F�gXu1���_h8�8�f2o��ϵ��<9�������~�g=�����\Ld�y������?G128Ɍ̧}�څgY1�,��}���*��홺�5�1��t����ݼ~�8f&���Y��}�߿l���V~C���;����c8��c�c�o�{�}����9��m���Ę3`���{��̟�~�.Y���bw���W��Lsy��k5MG5ì�������'��=y��y��w�1��&3�c�;���,���	1������n�N0�bcf3��~��m����S�y�돭/��4�Fc1��}�������%�;���a�3�Y�������Y��f2d�1���~����L�]��{q�p�G����_�c&?y���:���8Ɍ���;��+8rɌ�g�~��՝��?3����DfN��Q���缅�>w���!X�k�u˭r0Y݋c���vt$����d�0�'Oqb�����}��=[i���=d���l�|0��fc1��3���f3�`3����w9��4���H���x�u�9��U��\�̏�q�{�?2u����_Ř��j��d���~�����YL͘���8×��l�v<d�VJ��߻�|��i�M}��o~���Q3r�\�Q�u]��b3x�d�����˽�l����f(�p�Yu4��
�jH���4��}�P�'^s�߶u������I�����+6�a��J�̉���:ͳ��d���?t���סJ(ϸ{6~�c����lz_���u�u�1�a�c1=��pq�d�������{��,�&`Y���LdǼ�����gw�Zׇ����2bc����w���Vm���Lf9��l�8�&3;����Q�15��:�'F�Ͽ~��3�}w}��������n!��d�bo�wG �g++�0�s��:�0��d��28��~�g�G9��~���{����<d�,�L�f'�o�B�N2c���Ϯ�5MTG5���:0~���:��Y1���&Y1߾}���,��������>��������~z�	�N1��YX?��8�2VT:�f!��^}��?0����7�~�r��?o��sK���8W\�I�̷�R�at-����gfb�&����g��b��p��ٸ[����#��<N'XgǬ�%eM~�48�$�q�ɆY���ݜ�d�VJ��Ɏ����}�>>��<X��qW�8��#�5�B�l�����o�q�|c10���AQ�ut.ɳy�g�#O�~�<G����f1�ɼ�;�?�u<�\��1�Cc1�&3e��yì��3dq��y�������f2\,�L��x�S�듩�kz�f�+�5�~���].���1���<���:���̙d�fY1ן}����~f8$�c�1����)�N��_�CF�e#|��	X��Y�?p�w�W�ܻ��nm��d�c�Ѽ���Z�%� ���9�\�r���E䞠���[��[�]A��u�65z/0��4.{�;�t����T�6��Tp�u�#۩A8,�_;��X)�Z�[���3����jvz-��6|$�^�{�7O:=S�}���;7�%��ge`�0J�l�L�{�2��g���N��%>1�����$;�v�Ϧ����o��'���K�i>V�5�}�y�0���-lyΞk�bڕ(��]�L>7��V�9mr��L�m�4.o�6r�p�Ł�M�U�m��֕Ӓ���bʶ��}�rq�VV�x�]������F���u'��=u^�U��~PuM�XCl����;�0hO�ˬ��N�r�|���jaCt�{�vv�������L�(�C���^��.�{����ݸv�#����(�Z�:�	Иft�g��^gG���u���+K.���@űU�Gpއ�}���Aخk�4�_�\n���]Yban��?
J�ݰ\MͧvO<��{��K	<��@v�t�x�"�+�^�}���^|�R.�('A����BE���4�f�y�1����U�pC�8K=O�U�R���j.n��4���l���4Q[��$c�a%�շ3Xlb"K�YX�N�̺���C34"�~�Z����q����7�e�6��y?n�@�Q�� �Y��S��FEҫ�D��X6°��R��m�����4��+m�,-������*���J��+*V�H��]P�EVER(T�m�����FT�-���(�
[Q`��ĢUAJ²���e	�)1R�*
�U��q̘ȸ�1	XVV,�XVJ�ƴt�qk$���Ze�d�eq�4�DP0��Am�Z�
AX�U���KIR�TY�AƢi�@�@�"��`�#l�h��%�VJ�
6�*8Ұ�I��&!UP�4+�(�2�3.D1!Q2�AJ�%[a���d�*�Xc]Z*�"��i�B�Z�U�I��j�+�1%a�K�Qk2cR-[h��PUE1
��J���mV�������khX��H��Tr�Eq������
���1����ȗ�y����:!��1��C�����g���1���3�fi�Y���ΰ�L~�;o�����kLK���ɇ�G�����UY�=��g/e�Ɏ	����}�gY:��d��1�e;���+=�{}��u߻{�N2�VVw�l�8�c12w﷍�E3ZNC��ta��}�����0��fD1��YS�k���ֵ��^�M��������g���Ę8�I��~��?2~�f2\,�L�1;����vտ���������\��K� ���<�=\h�<��뗋����C����7��f�����=�0�4Q\��Y*|0}���:��Y1��Lfe���l��'�c�1��I��þ��³���3����~�߿m�?C������3���b3�`�w��>������a�����^�c�N�g����5����g++'~��N}������������3���1�Y+���>����~q�Y+*w�}�Vm���c1��������?g5��3��I�����;�SFk5�Z]:�6Χcw��>������!��dC��u��Y�8�f2VVk���>����}�|x�0�Lf$��bLw��>�����f2VVK�bw���Vm���u?~£WK��gd�v8���~���<�;Z�����|Y4��d�d2ɏ��~���O����r$�bd��p��q�3++�=�g���� �[t?g��΄�cl+��症31x�8�	�T���=�g�)�2ld��$���K�w4�Zt�^��o}��kf�7�5��$!��C���d�߻��ΰ����38{�����n�U�1�d���5���q�I���L�f0.��g�>���q�9�|G�}����_�?'�11�LfN��5�9d�\�Lf8!s߶u�z���7��u������ѵn��p�����Uq��ݬnםl��ز�Vw�Fo�������.����u�d������|0��f!��`�3���Af��1��1��/�{���:&3}r�xc�i�zͲW=���:��~�.K1�0��{�Ax�d�5��9�ц����u��c����ΧG��|G���h�K�nY�&K����@��͝��~f8$�c�Lf&wϹ�,�q�3 ��Ŀ���:�3�c1c1~W}?h����|�߶~a�?3g��٘�3��h�gtLf&����2VVJ����~�Ζu�2Y���c&;�.�v�s�}��O��q�1�N��5���b\�h�߿sWğ׺�YW��Y�`�B����`C��Y��y�GT�N��'ջuh��}�):%�<o������潐��9n`Qث7��l	�{�0�]x�:�`��UҦ���v�X6��f|��Nz�x���x��ͪ�|VrY�n���N,+:�y��ך�i�l��dZ:�Q�3 �oB�)El/].M�i�&�?Ϫ�ﾴ�+�\nޘ����9G��v��nTy�c`z��[��|A������dص���O"��Ϸ1�=�������{�<�9���<�P+�E���������f��[���XY���� ]�vGxױ���u��KZ�-Ϯ"��
yG��]u�[���n�:[�ov��ζ��C�����Gl�l�ٺ���֒�z�7\�6yy�9g=��U�÷!y��V2r�5Þ�DJ���� ��s�#��9o~�>�a1#L����_k��V�l	����|�Nƞ�#�u�:T1 ��V���#~���UW������I5������u�| 	�w]X ��f,��>��\n���}/�q�-x�G�D�4 ���-�˵a�7;�u�ρ�k:��j�Q$v�-|H���^8��WbQ
fa�ՠ����d�n2P_]]�� �{�0�<痳���z[����_�Un�D�K�r)�q����I�y߿���mf��=)u~��9*�� $Nw�1`π7'���=��s��?~G�N'vMx��T�	�s��u��S���ON�:�n�>|�E3~?7}�x����3�{v�+	�{������`��K
�2�FϱO~��A$��$�	ه��	��οd�F)j���n���z�OVW!�辮�Ȯ����{a���y9��|�;�N��2]��і��R����g�=��� >�;�/�@$��=۸@�#���������Q3Q������nCR��Z=]y���vF�( n1�.�}��#+f&n�� O�ۙ�>�% ��>%6�m8�v���݌tm���IΜI%�sٺ� ^ͪn� ��޺���u�}�� ��ݹ�qz�̡,`��X����������՗��M]s�'5u��ۙ��sj]|���޺�~�����;���� �p��\5�n�QCYi7-�OQ�.�h�_.ݘ����s������\��{s 7��4��/z���vlEN緁�G�ݹ�0vmK�s�\!4"G0(��U��v<�yL�'��wo� f�7I �e�UZ ([��I;�vK���2h�	ه��2�d���L��.�m_�{�}�D�b/,�;Xk�ut��=S�U�Wga͹J
13ՆY���uv�Iq�լ�[2�^���#�Q�p�ޞ�;8��$����~@|��.�������]V�&�Q,�ϗ�f�V?_�_v���7a������� ��a$>�
%���n�DfT���
8%6�~8�~B鼻�H �����"�m��^�2�|��'�M�6|�^z��6|G�ݘ���PG�z+{}�G�.b\�Tk�R���
�>�\uԾ���E�.8äݵjy�����!�QQ
"`6�=Y3@؁e�U�~$�����@l��Wy.�]���� ��6�H�pTLB��"��D�v�}��݈���:fy  ;���� d�� vk�����Rn��6���B$��.Ы7�Շ�|����	÷�z<�M�2�L�I<H:��Հ}����M�>�L&Sl��':��ѯ��>�~�'�Hz�l�I 'w}�� nuK��r+Wt��}�1M��\G3M�w������)l�.�$s�Y��S��U=׃o`�^r��g�P�3�{��-"=�0-�.,����/��N�N?u�괈p��.��z���� �ٚH"�Uf�Fn{��������f%� ���e��a�ڏ���w�qRʪ�
��8���=q�Q�Yy�u��FԝB��q��3�q��+�tQ��mL��q8�
;2��ςw��ϰ @nuSt��&jY�w�/G��u�u`۞����Q�Cv���Q]Xud� ��&9��kzn�����o�3�>�R�g)��{5�`�TLD��"�������Ι�@�S��+��onm7�"w��İ`�vI*�7( BJꈪXF�ϋݬ_�K����|�Jg�3@Ԓ%v�d�	��]A���<�<����t��JdD��K��V��t -�mZ��eg�_���{s0�76�� 5CWyh��V��I`|�]�t��f�!��ͽ�r6̞yB��*"�3�d�A��e��D$k6�'��~ Ӌ+%�%̦�_N�+���ckF,�P��ݳ\�l�N	���m���c�T�$�s�^:v6�/]�睰�*�f�
�؎4=��lu����s�\��gak��.ݥ�E���b:yqD�hu��6�y1ȦA��uq�Ѭk���pc�^�]���`z�����s��ɗ�u�螠^��ʳ̖^6�ch#B6x�kA۵�=1�o���gv��X�ݯ#1';<�ѷ3[;tjgk5ö]���nnһ�������8θ���=��� ��VKxpa��F{��?�Ͽ]��s�Gҥ�q���ϰ�͙��Ht��W��W+�(�W�^��}��S G��]|&jg��hQ��v��Ȍ'!����v� �j��:��,�B��K��~��ꌂ�D�B�������n�f�Z� &}n�L���[z;6��6�������`H�b̹M_��v⒏{+:]w��s�3@|�׻n� �Oz;�C��Z���vU�D�~���H�5�LrC����,�uӰ}����˂�@�jꛯ�@:�����{٘_QS�4�S%��O�>mO|F�e�[�+�q(Up:z�Y��Sת�7tu������Js0�$�s�3��@�}��D�H�'z6��(��� ����#>:����ʷfĈnӗt��IFI.��^u�f1Yx�����&�>���w�gc�.nX$��ը�
�I���멇7V��E7��i��j�˚����|� :���� �o{3 �T�e6�e_S��xγ�F� χ��j���D�~':z&� x{�n���[�D�M�W�H��F��ɇ��S�Qúo��E/	���tn����V#��fb�s�[{0諹ʇ 9��ՠ�dD;��LK�D��N�nf�7:f�TD�)]̓@'9�t����b�� oz��(��}	�_z���9�c&$����ѳz���]im�+�H=h
{t�L/le��>�������C���
�m�nҰ��vu���2� ��}K��`��u�S_ �~�s�ǽEH��M�J�]��J�̢6��f�L�&s�1$�_V�f���()�vI/����"����wo7� �]��g�.���]�o�o�ibA��NWZ��o��m�X�}�	wl��ٔ#���E�L�W��gP$�,�C˝�x2�r�.6���P�_��c��%W���޻����}Y��w���� 'w;-����T�[У��ڙ���4
>Kk_�n����3=#���������$:y�Ii/�����qxo��f,��pݎe��L;���e�@|
�z�˶���NX��n�3 |�w�] b�o]7���r���^s$[��u��-�!�!bwJ�壮m�񓭑
9x��g���Kh��x���{�sI!��@c���t/d�<�Y�� v����x�!�08s0�Av���t����.������� ��� u��V���ǥ��E��}�&҈�&+2ɳ� 8t�fp	 
�v���A�^�A�:��oA��e�6�������Cؑ	Ą��l��̾/qzיOv�{؀	��  I���V f��*�E�(�q6��
�Y�U��ĭ�sxvBI�U�D]��C6���ei��g-�e\͢�7�o{X�p(��j��D���[~e �{aF��53���ۿ��yv� A�=���1F�T���GI;���6�?P�I���{���_�͸AX_C��*����s�h^;N��M��������uv�g��wv.r9gs��������Rwߟ�ȹ� ��V��(�������\"�jJ؞���v��q��r�f%Tr?sA���wR��:8�3��"@��ު���ۙ�>
��%�8�Ňh��@���`X̱WgQ�~�Ъ�4M�{�dMm�p�]]�X��懠|�κ��"3�r�|e��h�b&[d� ����5�ꋭLX� QWuj���ۙ� oO��eފ��8H���NgK�Ut7h��f�ѕٙ� lzk�	ޓ'0q�Yyɨ��˫@ ���`�{��) ����n9����O����&�������Ԝ��N�8J�g�iv���J��ӐZ�*l	>z�ek�f���Ԍ���q����y�x�w=���v�n�ޛ!�a�	�����sйz>�AO<^-��9Iޤz?U�p��}��
�=r�ḙRNܾ\�a��@n�Ͱ+;2���Xծ3d�q-��c3;w�wG�z�
�]��`��S��f��n�6���Ǘ\Vtv㇕��l��ܼ뮓ojL)n�5�]�F��̡��xI��L-��w5mm�ǡ\ת�"5�k�P^�	ޮX�b�DS��k��R�㓳z�fG�k��M2��Z2�`kj��HM����-�4ܧ���j�\bn�J�_��+t�t�v˭��Dw��{;m߶����=3{G5S�v��@Lz�v��;t3�,k,5��<u�=�[�Z��Ǜ�KM�צK����c����x�rGİ�y�o�yﭜܼ��d=�%�a\x�,X��o^+��>v	�q['�BʹU.��E��򚦨�0�)���-�tn����h��Ղ�eL��Es���]�0��n�+���]Љ�i��#v�-f�`�A�z�th93ˤw)�>�R��D�-����-�s��*΋�_yGr���J�l�0�o��#��H������1�\�fV�Y���ƺj�t�%�'J�3���6��NݍL�{I��k|ޒD�H����_�]`yu��t�v�еx�bB�L[V8K�%�|n�{�{�ݛö�m��=|�j��-Xi啽�>���\7�'CL%E*]ZVȫO)��T��0��kj6�T���DX��m�"SM2ŭd�R��iR0d��1jT��Z��H��KR���QUkm����	VVD�A`�h��*�TĢ#V�1TQ�K\q��)j�CSV,Y(��RVA����e-J���"�#��&�MIQt*X�VTӎV��d��l�U!Z���b��Q���\aP�`�&R�!YUQj\��MZ�Z�Չ(ҵdm(��Ķ�*F�
�*6��*��Z���Q*�1%H��QY��4*-b]SV�P�T�I�,P�N�t�+%�chZ�"+#i5�LB��SHi�dD�**��eʈ��:LV�j�Q��b,QH�X��5h�Jֈ�bD����ł��uV���otj�b�g�{T�Y��{y�m���01n�.��vY|��7h���m�y�;E����at�D�v��(�؃scG��q�����\��:�:��km�Ѽ��lg^f4�<��z�@t\i�ۗ\��0r3]�:�Ŗ�m�mSE�h��ٞ������Y��w\q��9�c3gՃ���[G*�xֹ�Q��t���zE�n�k7��|uڐq�;v�X���.��:4�]�8�;�^�:��.� ����C���������{F6&Ĺ��p���zLn���,\��6���6:�����-��'ɩ�I��m��k����Nus��/G1ug�����{`ڵ�pj�;C��mh�e�]�̼��;n!�B�O`7<�;0�xg&�秷U�:Z���6w'9��ˆ�ڵ���\����U=�s�ܜ�t�]��nϬ�j� �t�o6��v��:��o[��\�J&\�!G��$;���j�Á��u�`��Rv$�@�I{���u&��[+�{�����q燍��A\�Z��M[����I��Cq��]p��>Ŭۧ��n�j���v�cr����'a:u��=\�5�k�����GS�E��6x]��`��n��q��4x�˻.�;��{=����9�Dr��N��n��]�p��t6�Vl��.�%���vw#Y���n{,�v[q�A3�;T]�zƁI��"]	p��݁.�<L�4tmZN �4��mn��9(��>79�y��>3�ρN�ڃB�����[�s�W]�8��M�W<<	�n�=nګt�i!����b��=���p��n�u/Z�]ƶ3s=��ojt�R��7��͒Fƺ�z�Xh5Z啫����m]M�����&u���>���穗��x4�Gf��ݞ���G��U�xݜ�<�Y���P�t����y����f�LӮ�d�$�@s�桭Lkj�������s�'��+���0�E���'S´o.9�F�-�#��R�Cs�q��z�ɻd��c����3c]��vG����n����-Yh˞ĽV�y[�:�v�\19�sn�<<";٨N{[���C��:�O#k�ޓDn��k��i�ctq�Iq���uϣ��sj{u�3n^�X#��Vt�K�V����=�٨�"Qnlk� v����|�tI>��/{&��ۤ燱Hnf�{@Z;In��N7e)P� �J��k(pԡR����ug��k�unv� ݂�F�xL�����y�.{t���o�o.���ϰlz}@�r��Զ����@TI�����d�ia`��`�H��Rj���Ks�G�u���^]yX  J;�s1 7��W���E��#�7���Հ���dba˅2���=���` oz=5 �QT�_�У��M�����X1 oO��	ǎ�R��a��ڜ�M�����$����2h�D��F�I�����1�ߚ����$��ݖ�	��l���_H ov�ԏT¯��H�Q6�~$�����Y����^�V�`�rܱO���I��ɏ�Reqfv�:�,���k{$������D����<����ϰ�7��@|������D�V��6���f`���/sP'� �����'2�<��RI�L�7���S)m�}W�z���R�Z�]hpS�{j3ꕾ���Z�����xW^�Y�d�V!��|�f��h���o�� �x�L6�w�uk�n궳�a����_rXz�B�� %�	�TޗS @���Հ�w�]o\��| ��LR ����(|M#utn��"�0+���n��{�I��m�y=  ׾����3{r�����.�D3�|WLP��dK6<�vP�s��?I��rl�\���:�	�T8�lX�ިu� ���gv�}���Ν"���.��v�
1t�n�h�xù=q���N�ӗj���8�m�˱��S"Un��ja&[d��(�R ]{�iX|�3{s1���?O�
��z=�@ρe������4��K%�"��̮��K"����w������z�� ����V�|Fong�|��F��bc�c ����*S??�b�biR r{���$�{�8���w�h`jW� ���z��M�H��L����kD�p�۵ZH�9!�6kL�a\u���}�5�3~;�҇�I�7�6$���W� ������^PP��3�����@�x�9vw/�@�������w�oN��ea�뛭��:����m�Z군�$d��S7���X6|�N�ґ���mv��N��$}ٷM��$F{�3�lw�(r�~��q�%��9���99�p�c[a���[�!W8�2Fw:�v�>{���~��v�J��f�3���۵`��۷��+�谓o�zM��k����I$����2��p��	��%�
;��6I��Y��O �ݻ� ���E[���{�v���G0�b�r)*o�+�3>��o��l��:ƺ�׽̬s^��$���M�~H�޺%��T:ѢM���W��O;�-�wsB�z�n�zo�|�����D�N�*^�F���������C���N��٘L�m�(uu]X�L6ϷϸL#1zb�V�ߔ_>y�5�@@�Nm�M]FۉD�a�Xi�4� �_uS���jp���[�� Ѿ��@$������Sʜ�6)Q!ȁLI@�kv�47K�r7c;���Ny�\Q�_.ݘ�~��?v10��e�k�>��� iޚ���������2U�x���x�@#�ޘ�'7s*69�j �B��V27r_G�}髾�� �_ �]�UX{mT�5u�+�tr����-v˗	�0�m�]�wMH$ -�ڻ�A����_Gw{��}1@�W}�V�_zTlH��\�K�2��%�苵;xP�gd�R>~��դ�gv�K��'g�n[�|WLP*�d�pә��ɷ�����=۷�l*���^�Y+�uP� oz�� �ۙ���^�x���J�nHք.*}ߍ]ro�9�z_Zc#R�QqcN
2�2�)�T�ݞ,~����欋�r�F99{�A�zM[��N�����]�]g[�%�"q3��Kn��h��N�v3:ݷ6�{�8n���e���1�{m�Ǵ]���N��g<��y�	�3�;0��M6雭mXs:�l�z3gqx^�d��1\kp���<]<��[�#�8n���3v��*�������;r/>l��I�ƧO��K��sc�v�3[���˛���Ms��;�7�7T�r7B��ųש烋�S��8�P�k�1@�%o��mG7��$�k�i�4� �^�Z�H����A����^Yqșނ�%���]�UX�U̓��bs2�d����`�Q2X.�LԀ_uU� #7�3�8]����etMLj���ʆ69�p�݊�v��{{n�h��ޝ�,k�.�ɇ`|ϯv��Fonf)lj�	�0�)�U��������}��6�����@ ������ޘ*h!Afo���geSv�:TtH��d��ɮ��餤]��/��@	��]X ����x���� ����ۜ��x C��(@���L�W��" ��ŀݞ�OO����#�f��>����;W�̛|��o.Ղ@n��,  ޟP�q��:�o���>����Jn�J�\I%Շd\�� ڿB�ޚ4j7�p28Ã�ʃ��О�2���z;������HY;}RooZqd�r_VJ�l�%(�/3<��痾�kK�O=4I����@$���m� ޟIK�b��W�R�ɓWW�9uK9��'1?V����,���P�6:&0~{ﷺ�2'��� {{s�z}#n<�p��3:Ͼf����3g� ��˷� �M#I4I	w��gr�ʴ|��<��{ۣQ��RȲn�+�y�O���D�]n��%������I�I?�����3��=�Qq��]9�]���]��<܂�����5��[i���X܏3̉�ۓKq8p9H(��Yڠ�p�51#S<z��3���Ҁ ��uՠԫ�d{c���+=&p�RIz_����`�����/��)$�$��1�o_^ݿ ��  Or���	oyq1�y~��ǒ�	�9Q0�I.� ����@��_U�|�����_�bSKG"H�|ؼ���V^�bz+��k�g�9_������@/w{c#Jk�C�J`���.{}f�h|�T��[o�=ӒR ��κ��H�t���Q���B�ϗw��^K�AM�\t����uh�E�يt���U�V�$�:F�=pE���L1�J�H��"h��+�萕��um�n� 뛡� {ު������[~��=�dD���2l��n��q,e�*��x&6&K���\v#��{&}���y��[J�T�0{�Y��@�}�N�=���T��kS�������@πI��]ZWz[��9M-������fb�H"z���xukؙ�>=�m�$�h���̀=�%ӯj��'gK�r�̴|ɷh[9�N� ����� ��o#6.v��{3�2� [~ګ �n�}��V��sBrIu`�.W���SN<�� }�W`I��}ܓ�@��ӿj�_D�*N�Y�1�j7��q�^��}��]�Nn������~��ϠS�����ZN����^�//�s$��k3� W;�M�%��j�n��Y�+��p��#;-�f�"�b�T��'�����s4���khO*7����a�6����L�q�8k3���[3\�R@�s�ۙUU��*�%Z�(�d_���$ԓ�̀~$w�`�v-M/d0�[My��"@�ۘ���-Ks
	R��v�f���z���i��]���X�
d黡"RS�턊�-�'�M�zk�O^�%N�/��fY����m�����D��/�����s�
k=�l'�w3 oz�h��@(�,��Yig2�S�:�D|���@ �۩t�@'w�u{���wv���M��"ws-�ڲQwbHNI.�칤� ^�Z�t�ʉu��.�H	g{ٙ� ��s4�6�w�ua�U�K�������t���4�J=u�/{�6�75�d�>�.ӕ�?�N��8��g�L���5�e\sn�t՞�V���i�νY7&�qo�Ɵ�����Ӛ�vw\{3ƺbٟC��	�=Z�'n5GE�K�p\]u�\ �=���љW�7��v�Y�]���.�];�N��N���[���[��]6k�th�\���n��aS��q�=����=Eۨ�%m���n�.ݻqj�$���zݶ��s�v�j9�ppN��ſ�>n��vٷn[��V:�c�و�n��- c����-�]Oa�\�f���KJ��h�x��l����!2"K��\�I�s������=���
�z��\r�J�S��˶���N<q`�ɑÇw�7�ՀVg�~��J�9i��m��  ��_ �	��]X�9k��*���K��<��K"ɺ�X7K3��}-��m�jұ� ���:zb#�� ���h��z黽��&`r��[S76{�3'���+� V̺@ �uՀ��v��m޺�~叩Sm��s4�hy�1��,��Yh]9�X|�9۷�a�r.�>� |��T��đ�E���	�{��r��އ!�ke7S��'��v[�dx����1���x���k��^Q�8��=��7��� d��J@ WY�N�N���ތ��nlA�S4�3��:��ꖉ�)���J�/w6ɢpx�j%�
�~�cj`9�is��3]����5�ٴ�����`�=�O�f{�#Q����fX��h=�zb���r�r}�oX0z_�g� �y�V�=۷�0�j|�{}s6�D���l�`;"��d��W��7RI%w8藍ݕs�u��x 	��]X�n�`�|�e�rB��)���r�V�B���(�ڻ 
��s3����ܭ�#��`<�˫@}{�zI!)�e�2��m�I&���Xyu)��#�ӱŅ��']�uh 
���X6�c�b�}�:Ѿ��W�V�8�%�0`m����� ���TGcq�\��;g����7_?>���(c�nX��-�˻ Vom�  -���I�uj���0s9�V���������@%B���o���GfF�WfVA�u�VX >@*�n�`��ˢI'���>�ט�ԗɖ�����ӈ�����Հ:澐A$�'��uOVm,s.nw)����J'�躐5�5���b��*����i�9�ܲҞ-�gT\~"����`�Zg_u~A/��!�'5��w�9��
�y\�j3�w��9b�Ջ҂��#�5��I����f���J2#n^	~�Qn���f�l��)*�L�����$ߟ�?L\y�+�zF����Ǽ�v��#
U�hM�lG�)�+.3�J}]��.���}�鸦�s)��^rU�1�+nn����\�s뗕N��A;��?7��fB,�#�^����Xi��hʳ�Ft�&�P�/T7��s��r�YK��k���F��O5��ҩ�
��㪳N�I����TJ9�v�[jb�0>4�9�B�n��L�V��.7󹧮9�B[�һ�}�5[r��,Dh<&�.��G�֋���a^���B��,����ivL)�9۱7[Tgg�OX��c;<B��v �r&8r��N�e�e�ub��3i�pʎ�Z�ŷ�(�"cė�A�|vCVy�=�-GY1>P0K��Y���"�����ug#�OJ
�lŉx&S;h[�����d���/9�3��cL��"�2�t��["^��]�	C��Ie_{��tS�4�����{�|����{x0M��:s%+��A��M�u;�,<��wf��֦��@�[z���!�C���:� ��!.�24�����6�p�d�f�76̩Ҭ�ۮl���9�l�eM���V!���}��n��'��|9�mΏtpy�@8E�Q��lSV�
�%q��EQA�TQF���5eՅGV�T���l�ж�PF,EPEQU`�.6#Y�t�Ҳ#�QEQd�����Ud]%uh��Q\I���b�+*�jP�̶��̶)P�����e�ɉQtܲ��(k3#iuM3I�E�4�LJ�0X�r�D�*�&�+&&+��j��� ��P\E�A��1T]!�b���Q�[1�*��Ԛ����+�궍eE\�R�4*�m���P��4����Ll��Aq���%mkh-�"�L`�*Q�(�naY\r�T�U�	uj��Z�#b�q
�լ��Ԡ�UX���\������P�TDĩA��Z��DƂ&Ke�[`����Y\"�ݹm� �똠8���1.�S���)�_�=�H�މH��l�D����p�1��T��7_�����f��yC,�D��lI%�B{c��[3�o3��
�pI{;t�uJ�a"�C&�x��^��q����m�mˁS�$ն4�9f���ϡvG�Y����KU��-_�����!�[u~_������ �niH| �:���Ԏ5;L��sܣ@:$������O�U�.��$e��s֕"�����s�|� 4�t���]_��?]E����w_�����HLUy���J�!�y���$�����<��9�'כ��z6�) w��VN��U�U�U��1^t��T��G�բ]�ɻ-m���R���n� >+��p�#l���I\�K��5�p��\�Ŵ7gz���3�o�������	��1f
Z�HJx]�[��b�뼽b(��"c�1HN5����x	�	�9$I o��M�\Pt&�y{���+��a"P;��d�H��f��n��O���#�C�	D�q�!K�����vc�nvղ��E[���ݵɱӻ�![������z&b&fS�3��l�R ��W����s��%�R��V{,l�e��HNΪ���{0�r�-���F�ff` �חy���ͩ�  �sn� �+{�3c=�7�G��J�0<�C)��LYbܬ��@ ���ŀ��%K��J����@��j��
���Xu�
!����HDUZ	��]O4j*��8
��W���|�����> ���������!��	��]X�U�Ɉ�M8����M�w-��;�4�]llv�Z�Cb~�˫@ O�w3�H��M��ש�P�N��)t�]7遾��o�~trv�{��.��$��Z9G&)��yז=���^h�]�-��M�5ߵ�v1�o��X{^���h��^Oj#&�˛�:%5~���D�$"g���v.snu�� {Wu�)U�m�Mb-O>�[�"qz�:��vjٺ7�/:����ʂ�h�p��y
�旓e��t�Y6�=1��k�n6�p��Ѡ���ܮ����v�������z:2��=�i	_�a���7j�Xy��L�<]0#\cմ������v�ݸ����Ὀ���[�tpt��r�6ק
t��+����d�nơ-a<��=m�o���߄3���`��ջv�>�����ϐ };�M�{JF�D�>�v_���	 ����I�p^Y�I��`�m��� ��b��E�}T�{������T�@���=Y�:��TOM�~�0{ ���Õ�f,Tg�mD���v�I$����ު�P�=��I=޼� OuK��pk�p��!1e��R��C���!���b�N�$�o��,$�HT�m�{_����TK��v�%����P�v70�HD]XM��|�ڍ�U3v";z$�E�	nW�3 ��2��	��]Z\_���Kj9���'��]n�Yf6-����KYsÌ<���G�HȜ���9�	M8����N��b� '�f� ����]7~����m��}�
ۢ��� �I��ۃI5��5�3��`���,�� ������ܖi�o�#7�K�o-�Խ���3U�u��Jz�b�+9]����Ϸ&Z�gXU��.�Y���=%�����'�2� lN7�u`��˜�|:���>��du~�De�7��rʰ�d�b�w��R����+=P5q1�z��}�.��'޺l�,Һ)X��ݝ}��3�����HS4�|�n� >+{�.��p�I88��sۃI3,q�#Y��r�(�ۻ�A]��ϰ���.�A�7�-�I�ͪn�ove��w�\�~�������il��t��oX�Fנѫ�Sٷ<tt�]�%�GYc��w���~���6��Dz��L� |
{���@[ݙ� ��U ]�뷥^ώOn��I42=���;[�� ��"~qn:�opDj�h�u��3&l>���7h����?=�j��-Z�t���Ě�|+Hf 	��
����������	��*7�)>3]����v������?xN�'�h��� 5G��"�����l�Ӳ�yK�=��X�¯ ��/���-� |�}�W� $Wwfb�F�!�A�ĄL�&����1�p�c�_�!�u��|חW`�@*�M�'BI\�f>��UuR���Ƨ����t��.a��蛛6�31`��3A׆�ȭ�xu�U����fg�PW9�&�Kz��M��3!K�� �N��l�\��@�-]��&�r֑-��<��q��ُN��$)�� ���on���M�;�K�u�,$d�&�=�4���ՠ������ʈabs �".��L� ���Zj"�Mtױ��5��U;_��%y����w�]]���3���\[{�� ��"~qn:�o~�@ ��� �w�^�k���ݫޭ�V �v�����t�i�: ��j�Tk��;X�=��Z��"�2�������z�t���ؼ��9V�+T��YI��2��H<����9N�������I�����1�\���wT���Ŋ�hb���d鹚���W�?��h3&��G�)�F�OU��H$�6w�j�*g�]�䀩����=;% {]��2��/��;�1�L�((�Gd8�ݸ���c�kr<�B��d��9ɮ�Ģ&]fy��	sa��9/+n����z6i@ �{]��2���{q���zV�ۙ��vzJ�����"g�a��s{w`����VoMm� ���t 	�w���]q^3K�.;�}ڗ��lU$���E]UV2jV^����W����s��kr.�.���` N�I_-��U�ŷ�9�	M2'�d�v�3�[����Z�t�� $���W�6�ٝ��wU|�*i�?SR7H�kE�d�K�5��$OĒW{�:dvgy�]� �OĚW�l ��-TI�I^��l�O�3���a�Vߪ�ѷwpBpϝǕ�Z��w�xu�~ȽX5�ݫΞzd��	��:V>^�+�r.����"����4�Nb텏W^B^3�R�K�$ԥ�V��i+�R��\S��v�vs�ٶ}��ƣ�tRn7P&�s��3�k�D^G���l�jq�ktru���ܻ�;��O;Z�{�5�ֺ����+�.�s��|�w7<f��X�m��s��\�y�۱��٭����,=��	g�4[�\����D;�)ͬ�B�����	!m�����K���s3�c�5�q������>X�n6��F5�ص�u���c��F�>�H��	�9۪9��&"&e�|/�R ���;�v]�Gf/dEil�ka�1� �>�۫Gl���TLH��͛}����<�}�WET���]X_wfbX0=AR���vGLx���4&L�, ����Ӵ
��H2I?rU��.����jk������y}nT@	�n&""��I�59�o�O3��E��N�U� >����� ����g�5��o�'e�@|�۷W��`�4ȟ�ێ��԰> (ޚRv�{޹'ސ�˺�� �������:�36t�3ej?9������hB�J��۫��,��x�I\���և#�H���k�2b%��\/n���	 ��{/��7���z<UE�B�5����I$/O4��=]y`�YI�F�x��d��}�����mv7�;��/:�uw�أ\�{nF��묜��{ԛ��$Ozr]����D:�����W�8�녑3yOv���Ʊ[�-��sͳ�$���n�$u:��C���9~�j��Sy��mr����J�����m�ff��ݖ �wl:y92׷z���$�:7�ѽ1H�|l�ML˖���HW;���^�"��>�g�0 _Q�贉@������>���i �y麰>��*�9m��D]XI�5�]�R2Zr�<�4��\����6�£�0۠[��V��c}3~t"y��$��J�TkF�Y�%�t��'�u�w
���H�A2�5���$i�?9�D��s���_H|���Sr�͑���X1 ��t�|#�`�1��`��5�<� 3S���t�zO$'�t�e�4�C���D�&��������y�޵a�$�2���<_M) ,�ڴ�=��z��B�{���nYS(�.Sقa��0�i�G��z�����P =�8F�/]��oYY&j۾����J�tͷ�C���� �����PI7;8�Y�h��5uh���6���d[&=M��@�JFπI�_]Z _onV�Ӧ���pK�P����>`�Bl��M_M��b�ݼ�>������SQ�q�P�	Fv{9�E���r�}�C�fd�~�[8GX��n��VEv,�#���&�s����sy�c���߼���hٕ>~�#���I#|���I''M�k���-�*7f) `	��]Z�o]��Ă���bUG=������}�c���xΟ|�6����[���0!��yh���L� >��P�m,;��=�@|��{o�\EK��uq>� d�.Z�I��s2OD�l5!13(�-�Tt�({��>"Ȭ����uZ�@|{�s0�l��*y�7a曢9WmW��|���¯s���E�� ���i���0�P;�F��r�n��F����:I/3���ޛ�$I���I����
h����t�^m�I?��ͳ��By6m~��y<I��4j$�����m�ǝ+�T���㸶%su�̳��xlq�6��k'`;h��x���tS���f������n�Qn�
���X V��� 7[#n�|&�xlmW�7��ϒ/zLѩgi�@ұ���"��z2k�1ѥ�os`jX�b�onf �:��+�`l�GUu�����5�8i�e�j�D���w��o[4�>�Ҍ���8������� ����Q%'/�4�B�� .�V5Q���s����诀A��� 	tl����]*�cjZ��]X���{�Ѡ�Ȫ��+ZM6�6��~p"A$=���Kg��/@UY��πF� �{j[�HH@����$��I	O� �$�	!I� IO��$��$ I?�	!I��!!I��B���!!I�BB��$�	%H@�rI	O��$��$$ I?�HH@�Đ��$��!!I�@�$�H@���d�Mg1� ?~�Ad����v@�����6�����)��P�h;�     昙2h�`��` ���T��J�� 4�    jx�$���P �     �ґ�2h��4i�F���4di��&�&	��0`��"I2&Dɤ�FL���i�M#���OЧ����5Db�%��~ph@��A[e��J������s�������h��P��`�q@bQ �C�B��,�$�e�@q�ۊ�r�����o����P:�݂�D�*�o�8������fvHxW�p^�1�k���ڶ�<�b�	x��4��
�-�7�Ȩ	D�̛��j�ţyD��;��b\�dfd��*Lc�p�1r3&3!T�A�&�uv2q�*��&f*�Ɩ�먟Y�Ш����OVt�a �Ϫn���A�uIʩ�v����堠��P��u�y��Sur1�.�|�Pkd�/m1�N��}��T|��Q�#��q$!�ĒD�H�!	I QX���pۀm�"@\1H��jΓ� @ D	 ! -b#	!I��@`B@d�$5CI,�Qtڬ���"ڨ�.g�����	#q��e�������@�Zu���f)#��"��X�1V��!KR�B����(Ԩ�-Q�m� M#xƘJn���Qk-�jR����Va�	
������~rNDU��Ù�cwA�@1w���m�Wn�|�V�x�WKr�uct�ϘC[[���'Vn��P#.c��
>y��+<�uM�퍶�1���ԋmJ,���p�"���e]/$�9�&+�MQ��WNϸş�ўql����勒��	 �����R���⡺����N�0 x�2<b�"��X����n�,M9q�x�#�`�<�F�zAN! - &�C��Fsw�jm�r���3���ں�9z�HBYCùz*�,V@����]᜴%Q�/��I�\8X�,j�GE���靎��dz4<�\y�������Wݝ3��;�6Hv�PD��.�r6��j9r�YjFcs�(Y���Y{-VV�{��fC��JF8h�w<����+Ʋ���)Na�7>��D]�����4[�`Z�7�HY��4�L�NO`r,�j�s��s;�k�G�xgP����(Y͐B˄�1ң�H�f�b71I�sa�S��NfFw�B�Ѳ�v4k6ẁi�'�L������+�R�)djZ(q��]났�CU.=�˸��5�f��F\yE�K��g7'lP�(s�p�dH!\C&P�I2L��;��MG ��*2h����i��7']���S#��"Ξ�!!~Bʶ�|��r�P�2 L�Z.�Mw���*M����ڶ�C�'�i��
�#�/���r�(6����a"����&z��{���|�'��,�:E�̘2M�i5��dqt؆x;��p��,��[��	D(��U��"B�kJ����l������Aj��(�6|�"8�2C>{Q�EP�]ͤ�����T�b��b�.��6Gj�#����ט%���i���N�f-&�{�D�{��T
�>\���:�;��-�1�&�N��"tI̦�Tޥi�.R��.[hSLb�@'�*���;�"������(�T�F$#�oD�pɦ�3�m+HRe1_Pu��2Ԇ��z,9E�հC+c2����S!�/`�w���П4�;�冧
�\)k}'�q�h��N8��WT�/�����C`:�����(�-��p��1#l�t2C0��cB�<�lXѢ��i3\�.X6�.�7 �Q���-�]u}`0\��Q�sG��$�Kc�9������a����C�v�����,���7{C�ޣ(��(��)���`w!;]Ka� �Q.tL>�h��8��nC�(�h�_�YW������;�,a�o����4ZN��r���U�ub_u���i��!`����D]̼� n��b�ἣ8�`�_��a������26=���\)�H�u���Ls9����(]*Ќ�^�w%È}P9�B_a�d����G��?��|>�+L�8����cB ��4�԰��D?ȝ;���,`�(�C�1ʋ�R����W�oy��[ђ��n���=Z����q��g�����{H��s�����7�44n�!�
_��
#T&\�,�����B�\���(N�Ö��4�OF
8W�L,�� q� H� �6lN4,��x2f-$[�7���g0��r��[SU��T�4�4��Wi�B�U	����ѳ&v��;���{TN�9�2	�;�������W���?���Cy�#x���X`�HX���Z�2������OV����ޞ�y'2�:������J��y_��rU$�B��^�/��$��K��c���}����|>�R�@68	�垨g�4c���C��`�)i҃��A���_�v��5#�>��7��F�L�q�eȜ=o����9�|%������p��Mx�C�7<9)հ�D�;�3��u�\L���%�={�Q��l��䆐�=C��aӊ�=�ܜR& ���7�0к1�om��`N	#C�C���߱�GnNo�rE8P�3N�