BZh91AY&SYѼ���_�`q����� ����b2�            �                                    ��  {���Pt<�(  0�  �  L�  A5F  
 P             (  �EP��T�J)UJ� I@��P�Q
�T�$ ��TT*�)(��U*���!
�*�U��J�H:��T�UER�
�C����]��K��8��*΁J�B���P.��*�vw�;�ԷR%S �ʁf�   �Jt� �)|�%
^m�4�4�.7�DI��)EU��cP���� ��� =�^T!� D� � �@�1�  
( b��OJ x�!Q��TDQG�TUO �y�������<��� �y�R
� l�r ;�Џ}p@��� o/%Q< X�� w�   :}� #z}��Xy� W{�J�| 6a��Z7�א=� ��;� x{�����Ϙ�9�\���>��%  P��I}P�*�ERP$�U%IW�:�S��|��n��0=� ���� <���� ���@n�Cv �y�U 6c����   C��* 0<�<�@�R -c�G��u��p��Ԋ��� ����<�0�@ �>})�� {�$�THP��P�� ��1 wX�7` "�`ꨮ "8� ���!\�����`��<�����@�Ѐ  ���)+` @���8��"$� [@����`T�B)p69 �������   �s�ҟL� }�D
R)EPT�OMR�`����!V� r�{��wI% 	�2@d�ǽ�V���� Y��   ��I4P `�0>�3���ި�� { r]�� ���\ l� ��2 ��`�  �    �  O *HF� L &�0�~	���� �&� 1   �Ѫ�1IJ a4CA��2�l�"i�T       %?R�J�L `   LMA�QLLCS!�S���O)�}��~i������S��-����P��vw>�o� Q�p)���^  T��*"�c�<?��&*�"�����C�G�?o�?�}O�t!��	�����U��,�I>h@Q��G�'� *�������x�H JU[J���#��@0�p��� 	�t@V�U"�4UG��*��Q0���Q\ #p�.E�(�nQ� B�Ep��8AFh���U �*�ERҪQ�Q �
3EEp��ªW(\*�h�-ªE�(a[�Q ��QZ*�a�T Ep��8A�	����G3EL"�+�-"�Q�%¦f��E�h�A&�#4Q�ᠴ��I��.0�4T�7
8Fh���XP�h��K�L M0��8h4D�+ip�¦&�D�P��C
�G	p��¸D�(a�C�EL#p�i��h��K� M0�&�D�aSD��.0�4P�¦h�iS
D�(a�A�a�SDK� �0�p��֊��G
�A�*a�GE) �
D�(a�GE \*c��� \(ah���L"M�p��h���tG�֊�A�U��W�
�@�f�8E�T��S�
8Bh�iS�
8D�(��GF&t@�Q�$�G�
�D֋�p�p��I��.0�4Z@�&�����n0�4T�¦h� JQ�&��D�T�ц�.p�4P�¡�I���RҦf�8@�Q��G���E\ \-�\"Mp�p�h�H��p�p����!�\"M �(@&��0��p�4T�¦&��aXT��C7
D�*a�\�JD���K�L"M0�p��I��n0�4P�&��D�RҸD�*a�GEL"\*ah��u�L �0�p��I��.��	J�D�T��C�
�G�(h�p��	��&5�"M0�h-(�h��K�L"�!�:¦�E\ \(�h���$�RҦ.0�4T�0���
�A�(a�SE�*aZ*ah��K�L Mp��:®��EL \*ah�����J�E�T��S
�D�.!�G�EL"\*ah�4\ kE"Mp�p��	��.�0�4T�%¦&��A�P�$�!S7
8E�*�Z*L*h�F�].0�4W
�@�*a�KJah���L#4T�&���C$�S�(ah��� M0��8ht@�*a�S�EL"\(ah���L Mp�p��	���P���I��D�P��S�(�I��.0�4W
�@�(a�CE-)�K� M0�p�&�@�T�

: �*���  �0��"\(�&� ��U0���P�*	�u��8@ �(a�p���UJ@0������(�nT�3EDp���Bh���Ap�8Ah�U�P(�L ��\*�Pf��K�p��QL"�p�Mh�&�T�
���8D�D �4Q
E"�(��f� �B�Q"�4T�QI�tDRh��T�U �� 7
+�(a�PtD�E #4US��*��E5���UG�\*�� f����0��@ #p��H@Fh��Q�QS*MA�"7
�a��8Ah��
 芤�T"p��A�*��P� 4A 0�.� �*��Tf�
�B�DJ �I���A�A\"�4U
�*&P�	���@F�P��E��
#���Ic�<�'8�����/����p�{6~�{R���z�0������8�n3�Ts���^�Æ	�z�Ӽu��*�N�8�Pb�	�Ġ��zY�C�� ᴢ��5En��������;D�x,�m�ٺ]��u�;F⧨���vl��:��u��a��{�+3�ћ~;����Y��pc���2܇���J�9 D�{#0�O.��J�.������8���b�(/=W5s��{#����*��*�X;�/
:�u��54�άu�O+���achM���7;�3&�8������
�Xٙ�8����J� )a��?�fr�[�F��=�]ɩe:6�z�H�
��.����␍ ���>g������hz����s�;�3Bz1Z�9�.���ږP�ވqٲY�A���F�EدdQ����	�VG\�����ln���:��S���`���l�,�`q�c+�7�!ث&=������2��Q��n`����8p�n�拻��ۤ�"m�b�c����{�w;U�Mb���q��ur��&7�۲�FT��ʼ��{�fM;*;a���۶5j������x��P��	�P�DשF;"�����RG]�9�����n0�Q�����4ݽ��*H^��bP�9���(Z�r[� ��q����\C0�GOt�n�w*���`����j��1`��im%}�̅�@2�4�t���j�,Pr�ҐMu[��U������K#\���F�b���c�wL�b�!�{���u���wfq<�����	;�c�t�܊�l�8)>�ew7�4ez+ެ;���Itb�gG��ì���kze_w�;[!�|�����3�ȗ��L�3����\-[:�&�tn�[�xX���a.���n"�b�^V'��Ō�q��l�uw��x�XH�4�:a6��5���9�r�U��Ҵi܌�]%;z��.�V[�e��}����zK�q�9�!.t�͵n�I;�(A�.r�����O���
l	)yN�7����pcF<w���p��1�����P%=�UE�]x��O��P��9)�_n�w��j���Kp��]`����L�z���^�2�S܆0��x�.��^ ��!m�����rsJ;6��V�$hֻ�iޫj�T��r�M	^�I��ua�F�4ŧ6�����Q�a0�� �j��˝\u��zܽ�+�7��#�5ΔF����"� 6�;��.��q!��s�p����z���D�уwB �3���s����}�+��`,�r����ra�G`�ώ^�l7�Xz�9'��|B�3~�'k<&B�i���mk^ww5E���gr�� �8b�~��ɭk;�h����t4��f�pY�w��2@����7����80�2K�����:��ی�a%+�`Y�������˹rܝ{�;mV[�A�:��0�������á�V�8������T�;����p L}] ��-+7��9�9N�.f���>�؄��f�[��:�ո�y�7zv���I'e]Nc�j�"42e���'��-�F�;T�Ds^�u=\y`�١ъ�3r��+�k�I�!�{�����"��ܼ�K�":(��@��qk� ��^ƪ���z��곆��(믖>�k�u �t��n��VOA{r�^й��F�"���ã�:��M���-���	�sd�p�K�Ú7�6�u;2��sf� �:1^���КjO�;���w��I着�\SZ����s��&�8�{[7�]�;��Ֆ-16��r���*�^�:�hcc�p�)����Es�]	�ts�͚�g[��R���k�[�ۑe�9�8�l�s�4&q�j�z}uoy�t��<0����d;��'hI����V�r�05/�5v��z&t��F	�&[��:1q���/s�]�$�.ⰻ�}V1^#�}k�\�*��z�s�vo�2�
�I��o��+��3��ٺ��qr�Ml�۪����ջ��:۪�.\X�\�N<�f^u��w��\��*삆��.�L���ţ-��]ׅ��W��M�!?5�w&h�)
H�o�wö��UF��pe��'wL��T8vU�v��I��4&��c�t�/�lR��[��g@+����]���l]�Q��;�)p�vn[�l��6�M�\�N��NQ���-��F&�N�#蹮�{N�	cx������q��-��vL����<�����P}�B�w�wv�6�1J���]�9̑��k)�r�]�F�|��7:�EW���Z/�1P�˯;�*�w����6r��̓�.�'�ZX-�����X��L8�N���{q;�{�i�Z��v��H�w뛇�=�ti��j� ���鲌䨫r�t�ݷ.��}��̅���P�wE�Gu<�OCp���\XW�l���Ӛ.^'�U�S�N
����w^���n�5�;���Qj}�Y��5�&u�Pn<�0��[��]�#:��;TlV�W|�nh�i|RK������2W�]w�w�nK�p�L^j�>EB�1iҳ����GO#�v��$4Z�g{4BwC��Š�ʶ�kuu�X�֍gt�U;�pn�J9��ܽP��n�{��gbP�|ui�7�(tGM㳓uX��S�x�jQf�6�wu.������@}5���,hkb���'K��Bkt�"����N3O*97z�i݋V��P;��h&yݖ��NE�{nU��͜sA@�Aެ�=��x�\:�\&��4wnr��b�KZ��VSZn�:��bw7�%=��0�M}�]��U,�%w�p�N5vTEK:���[��a��x{�m|{"���w���/k;�غ�ǜc�Z#-j}xKj�5A�Bb�yb�%�j�wL�x�v���U��gM&k�w��'�o ����m<D�b�ُY���h}������n���p\{��N�
�'ےC�<ΰ��Y�2lk7�\��J�H��
���x�׋�getAݸ���%Jp���4N��٫B�L�-r����R��!�6��bR�~���f>|�z�vgj���^��9o
F%X=�Fv�cG+su����,C����[1� ���M�My���)x���Z:�ߴ�U;���]k!v��*\�6rz`JZF�B؎�ҶX�Z+e��&�f������XLk���&JE"j���s^�X2gN1�6d��r�Hx1^p�\$�#�&gN�B���#�K�s�(sc�H΁i|���W��c����#��5b��.�'K�˸�.Ωh��ܱ=�7�v���V,��9��ef|M����ν�	�={�����\���p�b�}{/=��:��x��/���]��>�U��n�E�i�(=P9��l�b4��c�;�p��(��)���ٗb��;���ͧ(�8=|`:�wbҞ��d����ө�w��ɰ�R��v�;=tָӂm�3��8������\�G)<Wj��y��~X0p��Nڟ+ֿ�v��ѽf��x%��ud����A2~l��`�*�=q�1/�l<�
ޭ͐��<@�[��|_܈�i��+\�`�8]���d���j���4��qp^Y^�g|�Tf��e���YǫO{�B�x�Ⱥ7�P=9�u�5v��O�X3�b
������2���z��zMdl��r���ɹw�g㓠[�|Sn��A�N��V��1�fj peS�\�e����$��=��Ȃ�֎7Qov4��+ J�M0=��<]�Fq��J�}v�����\X���g�r�3�;Y��Wa��۹.
mx��\����p���Ç��������*J �A�V٬U�t�\[N��E�4�����e�
�	]��\j.  mUZAx���r��h
���� u|���-8��{ɏ�㧅E@3y\<�E����<�w�g�����Y�b�1�qF'��� �� ���8s#{^�(�\���nkx�׆���{�f�
�m�κ:sa7D��+-,��aU�+,!S��i�v*�R�`v�x��b��/CA��̜�H3uL���EM�;��4�e3����0����a�<4��{vu���@��s{�u�˗	�j"�5�1�����j�w	/x�t�5�215���6Ɠ�S���(�QG\}Q�sZ�R�PBoZ6C0�Wg�10q�pjُ��仍�br�F��ԋn�!�i��Y�#�!d8�n�U���g=��ww;K*�;�4kFy%@�r��jd�K��v����;���8�҆ȷ4��^���W�ηz�L��~=�vd�IA������e������f�͵>����vF4���vu�`�z��֬���(Э��t�[�w^3�O���{��˚�\�>lb����7)}�G��K��h�e���A7mɢ�Um:�.��x�pj]0+�p�}�̍F`����k�n�ٹ�99�&�y@/\��v��r����q�{h�ŀ]v7M܂=�O<�rg[)�YV�î;x=�RU�=Nl�U�%tL�n�M����Of���������#�/><���'8��;��*��ӣ��r��@貼��b{�y�z�r���o  B<9���K�����ﹷ8�9p�+���K���B1ߍ�K��RCJ]�37q�'��[&n����n�z�PZ;��N#rY�&��90N���(��u�����|���Ӛ2��J<s��Ϗv�ӻ�`}{�9����9=f��D�H�����@g���k�N>�u��ASL�3�q�W�B�n�Ho:�Pkɽ�1��:-ƈ@��fh͂m�;��ܠjA�国q-��'M�k$���q��-!f�U��l�nB�-���)�0<�j��M���$J���p	NUWy�Ɗ�ӦT����ܛ�6�1�Lovb�Piʺ����_�w��s���x�����3�r��ٴ�)��Zjj��I��*bYoVygo�lg4��6��2����s��=(�#F�ơ]�E���;9m���dx�,bgvMH��B10�9�{��@8�89��ڛ؈�2���7V����]�	���5�h!%/4�q��K���r����gJ�[:�r����BD�:��r�wj��띝�Ǝ%��Ǯo\�v�]���Ë{;�e��������{�F�[�ǋ9��ݑe�w���v�s�V�.):�c:l���ъ�1w�*����43�WV3X����[vY����~>@3�Vh�˞���'m�Yjڸ�n��Jb��{�Z�'����)��{��KOћ���ҍ-m��� �����v.,744Y[����]'��r�';���fN�{_wS��[X(��Hmw�l��/$㤡$͎ks%��3��p�%�%�b�wm����`�5佒�1��+�c��Ϛ�y�q�%s��c�r�w9D��B۳:����&�g7��0w0�m�Նb��ő��h�V�	�e�BT1łc��Mu�3�w%U����F�dcA!����٩��~�Ģ�sn�k�����/i��Ъ�%�&���+��5܁��vo�d�ΨTx/�.�ב᪽�M�:oN�=��& �ʃ�r�Y��#t�7ۣ7��@�un��wFj�l��;&����G@jL�Y2�!�~�b������f��8��R�8�ܖ�M��%:�r�$ayզn�	���j��!�����p\pj�
�˅G��h��Z�>��e<�q����Ӊl۷����[tm����� t�{����|-�ʬ��>��q�/p��U4��.������w|鴅	k�o�m|^I��zᘶnn�t�c����d��k7������<�h[{��x��=�/�2��ۏ�u7��3��}9�̈́.��xea�'�����{LS�'��7���v��P`�S�l��4��͓���0����L^w\~hl��%b>�x�Դ�����n�����x"��V�$�RzW;���=��=�	��vv���!\���iq{�a}�nZ���`c�,�f�����������d˳����<0����n�r:�\0�{L:�����j$��m}#a���~2c�d��T�=���w�E^��[k����̅��[���inz�^#�d�$�>�>����G�A����q���hC8{��d�^��TL�}~�H�͉.��Կ�������T1��E�~��/.�i|o�z�q��I��J���b^y��P�R��u�0_߽����:=�����������c:�������t��B����Z����3�˪ }�u�3�y�^��a��N���/���_��C��f%��Q����-����a-�<�k�+�{�߱��ZD�������4�s_�����i��}�7�u�K���z��AY孁=����_3�ުp�]�#��i�l��&0�??>�<��Z��|��!�]�he���1{����@��4����V ���3[a|�te�]a�d��Q5�>��M���CC����8��ߟ���ޤ�%9�x�Gl>�#�V������M�.�?
�=���z�i�gN�b�w��d⫠�S�'hVY�L��v��Z?_T���Ʊ��/�=`�چ�XON��@�jb�	fq:D����Nb�(Nb�7Wf4.���s>�Ŏ�3Q�e�I�	���m#���ʫ�W��?y�ɻ����
lQI$U�U$Q�D>؂6*"H����؈#"�"���� ��B"��#"2
�"$�H�"���*`�( X�	 
�
$�(X�ب�
 X(X$��"����# ��(�b�� ���X��(X � ��H�"����*H��"`�����"���H)"�2*��� �* X
H� �"H � 2(��$���$�H������b%�"���� ��H�H*�
!"*H�!`+" 

  ��! ��3����AOO��+
[�������D�_Q�&���a������9�Ƶ#�f �-۬u_�3�^��)��X
��!
S��	nl�^�ɃF��8xxb�D���8�O&A<G7K�ͅ�L:(C�b������kM�5��cp�Y,�8\�r<SX~/��r�[v��ya@���Σ��V�l���	(�i�=}��{)#Ӣ�>�$O�0�m{�2��aH��OӖI�r���u�8�h��c��i��1Td�d�w���ǻ�{�yz�G����8 �a ��3�a�pqn��э�c_<J>��|7g���S�<��x�$S�"�%=HwRG#?�s;s5��L�O#*|||{�#�����m�j"R}*C��!h��g4-��_�@(��zň<97�Nр`�mf���&٦�{���Z%,#Q��j�1�r�"z=��ý�B;�s=�q��À�1wI��
xy����U��e�&2ḢL��PH�)�)�;V+p��G�9�����H�E�8��Ʌ[��x�p�Q"��� �p2H�H�)b,����� �Cda��8D#�H3oU�׊3ؘ��?<���Y��iq��(z���[X�֔�����D2���9�ݽ��QG�����b
��}<����A?��? >(��{�����8����~�����?�(L�QD���]���Q&���n��:��n/@W�����s�������-�=����[ �{�(��,����]����ޔ�Ra}	�ˌ�|�?p��j��z��=��ڻ��QK�L���ܒ���b�wq�U8r�,H��uo��SV^]�'/2���cm��di�J��mי�=��G�3�>��Q9L�ؒK�ѭ��I��L{����sa�>G}�N˺-K����.��fq�f��|x��9�w���;��x�d���~�[Ǯx�c���2�z�s�9z@{�ނ��|'����13G�cS$�O�n�W��!K�q�9�r���ݼ��E+�wy-��z{����� ��u���r��xi���X�|�K6�y,�L^��l/Viǲ!���w%Z�5��[�HU����'�f�#,�/��Ñ*��c��隷�1�0�V-�n���/�`�w���=E�O�#�z�pɬ�˺��W*;nY_��^p��x�<zv�ڷ5���,[�Uջ��f/`gNy�5 ��q��Yvz��^�n��s��K�?R�K'd}���@�L^�m�~[oxo^:�g����R��ϩ�)��;�n�6lm�oU�sU�_c(��g?���pr�����۷�Smv��M�nݻv���m�m�ݻv��˴۷f�ݻv�۳�;$۷nݻ9&ݚ�k�nݺ6�v�ێݰ۶�۷nݻ:`m۷nݻv�m�Cnݽv׃nݚ�k�nݺ6�v�ێݰ۷n��nݻyv�zv�nݻv���m۷[v�������÷f�ݻq۷m6�v�۷�i�~�6{=��g��+���S� S�J/�5����� ��A����ީi��Z;w��KĵJ�u#�g!��7;s�V4�)���"��<���y�;=���9��1�*{]�!��=�^^n
�<��3ލ�m[��E��xq�u+Ju.��|�����:�<���td��?����xh>z��n{�絢B�
���:�}���������/^;��{�U1yY3}�����w=��g�&\�[�m���|=�zj�#qO��O*[4b>;%�˾�c��{�f�WrX;ԫ�|��}�=���ۻ���T��s�r���_>�I��V篓H�/v�2���ӳ�L��~�����N+х��.@c�IX�����N������)�ė/5��x���U)��x���J�g:�ʵ����vY#	�Y��ql�X9��nb�=��Y���w��i�H�}��&�~>$=V�L��I�����=�����'9�ɶ�Ԡn�R�˅sR#* N��~����hn��������wy��}s�)�ճ�ċ�M6�Gxede�x���F<ڟ,�0>�f$`ݴP���d���ĵ=��F���fN��`�����&Q�s�n{�������G���i<z�s�W��0lw��}3�#3�R�_\�}ȁ�<��\'����c���۝=�{{6��l۷n��v�ɶ�v�6h�v�۷��۷m6�۷6�ۧi�nݹ�nݽ�yk�m۷n�M�v��۷gnv��ɷn��ݻv��nݻq�m۷fM�v����]�,۷n�M�v��۷nݘM�&ݻy��{vh�v�۳���v�٢m۷9yy,����ɷnݸv�۳	�nݼm�ݻvh���{=���y��հik���,��6\C��~��Do�����q%C����O0��Ft�E^I�����uX�q��s���ɻ�����{�{pz��Yi���G����o��y��,K��������������)�/6�h�{��@;�J9V�t�@K˜.@�K����^�pq�1;�a�p�����4���o�,�>f�/>����:��$��9��h�a���X5�ȃ�e����6+�^���e��Ife���<�!������b�2�o��}��{��g���7ؙeP��-~�Ǻ]���x�|��wz�M�{o�x��e�ϳɡ��Z;tصS��J�{�M�v�ͪ�(�ł6n�v�S�Q�k�zts�qK��v����8���_��F_)�@��I�&��'��*���Ȕ<��ᚑXd{�@���CVr{o���q����o=@3���g���3d�|�n4�C �Kpy��5��s��ڶS�z?G㺦z��8}��Jd���B�?Z���:�8Q��<�Q~�}�h+�;�����W�د!��(n��[��^�a��.�t�g��z�yxҩv��Opq��rW�7�����⳽�#��ٔ}�.l�4���qwg-�v_w��{`�/+��dS%E�@�b�
0`��F`��0`���0`q��6plٲ�6Sf͛6pl6lٳf͛:6l�͛6l���f͘lٲ�6l��
0�0`�c ��0`��0`��0`q�0@��0`���$@����0H��0`��08����!��;�(*{w7�;/۫#8.�:��W�z��n[�L�g;wY�F��x��O��;��h�G��#^�9Ǎ���gx!�L��?|��%���Y��&l���w���yq�Y�P�LC'��ﱚ��`\N�9V�'\�����ͭ�s�|�`՛��Ͻt�Q���F?f�6/5A�r'��5��6W�x�{��]���\^7��2��׳�e3�E�2��ݝ�O����
�{�w��cSS���L��o����P�T��v��'`�z/�o��K��Q�s�_�[O(~����{�}4��;G��NP�7C�+_�9�w�e۾}�_��%�Pm����q��}���������4<��c�A��|�p��}���j��ns�/��x�;`�F\[�J��{���ޝ�d��j���)��u۳��g�sݣ�'���}3�9|6œn<��5�#W�Jߵ)9�}'Q{��Gy�P��hW:�b���vh7����~��j��ϳ�C�:�G ՘(W����OY;kZ�a�u-�\ÌީB�!\칤U���^�	6��2��Nl���ED<s�h�uv��ٺ�"9��:��Y�1q�'ђ�Ů�"Ad����%Ña����gb��=�5%}�L�Z�0)ݚ���G�]�8�f��Q��Oa�N����$@�"�0`#0`�c0`��0X�F0`��F`���6lٳg͐ٳf͛6l��lن�0P��0`��08��6lٳf�M�!�f͛6l�ٰٳf0`�c0`��0`C0`�"D�$H�#,`0`��,`#0`���`2$9	��2ψ�[�8.�|�ۣ�?y{��x6t��G�{s��i��Y��5�b�h��0V�8��Wqɛҡ�g�1�A`=��u�{�C�fI���Ņ�"˂r�Ӄn��|<W�j5w�)R>~�<�>���̇��#/��>%p�qܓ�������wl��߰c8�������d�2:������;���x�y�F���n� ��q�s���]U��|��X���X��v�X�s��E�����ɭg5�q�0u�o�x���3�&������n�4Q�$��Q�,��w��w�n���H����j�9�����Batg��%��ඌо�������L����2�_h{��� �F�ht�O�,�<�ONRnz~^w۾�ٟn�*�\w��Y�x��Q�t�)�G0z,�͊�{���_r<- �X�KB����N~|; ���Q�Ԟ���?#t^����?A�NXd����o��bb�$�r��~@j�Gl!��8E�0�(j|�@d�1��a��Vz�<���T|'��I�x��E5�)�l���d}�E�
���1���%r�S7;/ ��F�oh�jO/�z�����а��=�s���!�}�t���x�B{l�U������0_D����d�W��p\��	��w�O>��V���'�{w�#�,M.��tmo���Kwn�9᷹�m�ۙ�A3Ǉ��ioH剎AL*"eH,��ƺ�V�3���y^�7(��gI���3���"uۧ����ܦ��ƘKs����N���\K�=��Y��==�8�-HF��{u.\;�g�ϗQ0�d����+V�$=��	�
|r���_m�ws3�g8�����2�l|�\�m��_�H��h�Tj��<d������v{�Y��Ҙ�x�#��/�y���K��Z2ڬu����ܼ��I)p�sS��S����h�izEz��ྛ��̠�������}j����n�\�j��g>#h�������<6�OW���7����I0�OR����n���ٯC����o��*�Wtr�x�m�}�B�͛�|&���B̈U���Zϵmv�15c��Uw�㼉�u��? �Dǲf�=���w�i�<�͙/�q�_o�����d��d\��6:3�{9{4hFxM�#ϻ�x٣��I����Nе���`i{_�[��7w�9ǲ,��^1��P\�^o ik3C���آn��.��zzN�KM�b���Q�:�񊊍|�.Y5.|���<�@ov�v�0�yw��pol]��Ӂrf{��n��OM�g�m��� ۂ����[�[�]���g�5�-�����t�L�r��fŒ��@���W�!}p���_��ZXwU͉Y־�<.�cY�m�z�{E|��x۾ha�/f�]p�[pg������\w垧R���|���=��p0Ksب=�:�9ϱ7y�=�rI�}M�O�F�15�-�R��z������jcSw3�v�}���!����h[�gr4y���1-�{����}�C<�G]���D�=�9�Njd2IK���f5OQD�|#��x6{�����9yj�x�	���=Q������m�+�E)�%�b�ꑢs&�ݟq�mD�}��vvu�Jb�(�m}�w�>>�7}�p�Jwr/�R<5Q�޵뀀�����[���Nl�,;�jjֵ՘]��W�(�{�h{�x_Z}$m/�+�;���"�t^ M�F	������݌���nu�8�	:����W���پ{���j�B�� �Y`��Ɍ(`c� Ķ&�ir-�#��x��9�#2�5W���D&���(��C�5O?�`u��n7�T�K8���{8���@qo��zk�����YM�`�-�̓��O~1=���%��e�~���qvɤdszW~���X�F��9	b�w^�PC�a޸(N&s2���:gu�>��L�'ـ}�d�z`�>�}(�6/q����y�FF�N�f�Հz���7g}���m>>���7�l��|{k�,��`�r��{�[I�w.j�2i�}F�Z�t����xz�^�C�{�����V�Qk=�6s��SW�W�p�<j�{�y|�K�;����#�S�W�7�Z9���[��c G>��
G7J(s�سw��{���}��ҳp�zc���u#����X<$����������T- ��/��f�f��C��?�٧�G��g��{�'�E��/_F�;zcVx{����Ѿ�a>�[�C$�c����!9�A��s��	�ñj�C��ǩ�_.�{P�8zv��6����������i��O�-�[��;ܰM�ΎSO�n)�{.�'�~����K׊ﴱ6�-3�篳�|1��%�<<���}�b���;ؚ)囖���=3(Y�����ûZ&5��}�{�+�H=w=c��� �<:{SI��{��}�,6!K�V���V�yLJ��T0h]ȟ�~����%^ʃr�5�Gj��B��
��ۛ�&6y���R=��H����-�}��j"h�:��w�������??'Ӷ��}̡��\�^��{NlS�`��gm֜�1��o��L��q�O��#��1o*:Om�/���V����̿�>\�@!�<��S�L�px�_���bY��} �,<VU��Z�ܤ�0z��XA����G��~�:V�yv!�ܼz��x�f��u�%|�/h��(�|�����ݝ���<�/�,��͞*{8'��_���|z���>��n�}8`��Or�k���+���) y�=�W��q��}�|��g��}��O�>��ׄW�>�������V�*LRo�73����\���߷�;��K'n��Ӊa� �c-0��wbׅ��uG���)�#���(��y3�/}_{u������ �����R4�L�{%m0����ﷄ'�����1���}E�\x�����(N��2~�����"��f��~xGw��fR��^������[�ƛl�;E�y�{yt�(o��w�Af�v��j���wP}����m��a��d\����/�N���?n�ꕂMX6,��Rka#{�f�ws�N��X*p����b�tpl
�9�Q�fՀ[��������T��a���{�ɻټC��;�x�:�'=÷��K�7���އ�n�H��|�	㥣��F��������g�u_�g�̫G�� {݋(kt-v�'��w�U=��xq}5��O�-����7@�s�mg�{W	�4��xsu���g�����7aگ7=�۾^V�L�Y�/��yx��ї���^���qU���Q��I�=�#���N��b������CHF�x��M�<�j]�_z��'��0	yݞ���]��.i��}�.xi<�g��e<.{BM�T��:E��teLQ/���+79��oqa�/D�#����&u���iA�M�f���� �:
��,=��c&Y���9��NgW���/݅i�kޜ.�9TCXkzEv>&�b�(o��������e�������<�gp�e9�|�]>�L���B��xf���r'�Fxg��tɷ;rh�h=N�S��jw��=l�Ɏ��z�h�qZ����\��ܢ�Fvr��s��W���/Y��£�f��d��ƴ},�&���\d^on�i�6�ܜѽ�K����^�rE�`�v:�,��������.cx����v�,էf9�9�{��+��B�\:��Gt�k�u�����oh��y>�vd�S�,��;�f#����F����`�w��y�����G6��7{w�][�t�����>��~�cH��W������q�k�kp�{L7�4��Ͻ��p+]����M(M]U^����x�������	޲�ƍ�釳�u��P<'��Gp�9º=^{{���� rN~� t���ҍ^>S������=�@�y��/M�؎����:�%�8¢�˴�''*��%��~��=�xxxW�d?g�����~����� /��}���ݮu55�����-6��lq�%FP���f��6&S	b�Q�0<��>�!#�
��K��h��iàl�˩*Z�Z-��k^�	�r���f	�MH�W!6�m��#� ݦ�`����(���5�܍,mqF*� ��eC�]�-�k�Z�hۗb9��0A�,�.��l�hKh�%�k�F`�ۍػG�QیY�� ,�����1-��6V�Q��8Ĵ14ninI�s�`�-sc-����K6b�3@�)��[���SM	`�.de�)t[�JaB݋F�$&��3-�����LL��\�U�Ͱ�w��WC���#*�]0h��\���9h۳%#-f�.��:�Yl
�j�֤�� �0�ݠ���(��Ɍ�ͷ[�X&�j��R3G�fuF&��t���]�����W` Р��X9ڨM�n-�l$�e��.��a�]\�r��MQ���i
��3AX�[n&�^��s�К41xQ5t�EC6�Q��ش���^ƕr�dX�I��������h���%��iFݚ�ek\]�{U�F��c+"Z��RX�t�:e�P�p��&���^چ�@ы.��1���mUr	
�.�S.�ͺ�ׂ=��F����P�cf̄ �RLb�[�����1��^���ݰ���PC�Y4�3B��3<9c�b�Du�1��HYw�kt��Ml&\,eu�j��k.&Kte�3U���Kq6�3���ɘ���ʹF�f�GIa)-t.�`�J�؂�&�,i�pU�LY���n�1,���&
,WBl8��Lqu!�^����9Mt �fAl�4�k�x�^���
h����--[x¸�dU�{;k`�,��m^��J�D��հ�ْ]�������Ȯ⋢�x��RjXd\m--ηkY��l#�%#��ւ�&���F�-1��41�32�ѶʹQ��Fı��q�	�T�J�i�LK*cLF���֘�-)�H��
�Mj]d�M��vQ�fv���M�L��X)����m[t �)�L������@[�H2��̭*`�I�mis�2��6��ѻ0� Jc]i[�f)	`W6��(�¬XV���0��e"��bָ�eƆԺ�5�{4rCXTۖ�m�niT��u��(�n�D\a9�h����f8KG��W'SV[R�5�^���1��
l����:���GK�kFKU�\j�f;�6m9�GR6�
9Ń)	���l��Qm�f�Z$�Lj��j�hG���]\I����W�7W�D�m�`:��ƫt+gFR5�V��'R��F�Z�n���ݴ,\c�n��/*��Nvњk³]i�-.U�F�8���gL�3!5t`YLLP��A�Wb��9"�&l��ɥ��a,��"�M�ܮL��:�oR.&��<���g�ˑ&�h�b0��e9ZY�ۥ�RY��ZW$�Af�b2띓�h�:kjv,������q�*�ɊK�eI��ҳF�gX�����!��)l��]F�9��J[���ы\b�D�� h��E�fЙ��F��$0�Z;:�t+�G��Kbb��&�Q��V�3��Ynb�H+WlĆ����umF�93�c1�e0V�ڋv��+c,�:�v��T5X$#���3a�ƹPb,�gm���Rj],M)J�R�[A��.ї<*:���adh�R���e��b�mt:��'<%�˴�$&�4f�M1�W��f[���D��]��G5L\Fi��m��f8:i��̖6]fX�ݎ�pm�cC�6(�Qr�`wcV�9�V�)���K�������R�b�ړ\^rF�%	�[���X�F��+Gdka*SG3E���Ma7]��#��H�q�`t6�j2���s��S`�*��&n!ƳZ=T�k6��]QD��J\�mJ��D��YK��$ \nx�)e���[M*3[���@��c7�J̡CB��Md���R���/
�&E��l�K��!Z]fU�eW�:��-Q�T�ʱ�GM�[�sF4��f��X͊E�A�*�,r7j�4J�&՚Tt���me�.��a�4��WSX�]-���eiinv�!6�nҮ�۸��qK����;qL��#�Ah;��$�i��U� ���,%�c5&۫K�]"��e��4�����s�ݍ�hV4^\�=�K^M5G*W�,�6��U͉�-��]���0���h���K��h\&��f��b)s+��nfk�vs��+`��w��`(l����M�M�mHj�G%�a��&���sB�᥸�i����4q�]쵐l¡�e�t���+l,fښṚ,�*nv����)Ƴbf�a�h,�b��Yp�c\�ᙤJ],phܛR�s	E����t�Ɏj5ƖTE#�^s04L�Օ�d�i�r,���oiJ)Al�VՍ�����붘�8��Ì��N�&m���]f�q��JsڨM, "�<�Gf�J��2�pZ�]r��l��3]1PKe&��s�kl#0K�T	�fRb��u�`ݫL�L[E��WY���3lp��.®�j�lm��[��&cYmI��㋉sR�8%���CM`荵v$5������;*�v���ƴZ[�h\u��&$���*ʱ�#��S]a�ي�ZƽS�f U��M�˚�D��V���n�e�X"��mi�A�kF=�١�V����@�[QbRZRn҉������a6#��[�]�0k�jsR��a��JMb��"Qa03\=sqx4+`��+-��6uXռMi��iM-(��v��HAu�(�\]�i.E�R��y���!�fGVZ��X9H���3d
=��snƊ7����M�#Sl'RUmBE,ټ�e���XV����(my1n
�JGl��F�M���-�f�i�b�7E���f"�8�lf���6d�e�G3Uf�˰ŚME�ݍ��C��4���ͮ�ԑ��(D���պ �8��,�A3H��#X)b����.meeХ��"7m���n�]5�5lU����n�q \X��6�,8���(��lc+`�ˢ�Z2�u
���.J���U!Kie�Q��G$uv�c\�B�`Z��Cv!��lػ�N�IM ��`1��5���S�u�"{k��Uy�ܫ֗9���5�ܛ��0��3���bM1PKz�u;:���61�0It%�HꊁqP�Ң�a�;i�X��@�+v�[�Gem��cKD$&�����&%����2�S	���I��u`�׌�	)�dtzW6j�
E����]*F�0�P�̴�nj三t�L �^���l�P�b�M�����V�#�t�f�n��ĦtBP[]m)���%�3[r�`�Bm�Z#m�5�P����\0�&�m!j�n�Ne�ِ���D��L�#���4�S�:ݲS��ز�mq)\T�`�#t���X��Z���ii���@��+t6�mLE�%�,��%f�hjlb�X.bC��b�tк�m�aI�^�,fDF*��Fa� �Cj�^��	�W�k�uJiQ�Ѕ!���A�ɠuҡ��,�Y��#��L�$rڤ7-�TR�ݮ�ë��h��Ʀ�m�f��r˔pGE`�m�	�ݝ�Xb�p�m �4[L�v�dv��*�!m� c���kΙwa����ڰH��ųR���ڕ�Mb�a��cT�6mL\Mv��r�@٩�&�*�Z��]e�����(������噬�%D�r��a7;[�f�:v��jZv����� !t#���n ��1NL�Mv�ŏ��X�M����y�d����\����+���78�a��bD���	2��[MԺPuƸк�Mk�V��b�٩(ECca�B!����;Y��fh��ή�VgYk�Suɴ+F�G,eq�ʰa�6�2ͨ�"��x�3l�lcF[���KA��j`�s��qEI)�BWb#�Ka���!D�f- �Aˊ�-u���M5T.��nw��YW(vY�1�	�8l�,��j�	��=H).aJj�ԫ�Kɒ��6ڰaV	zY�f��&r�pTLU�ft����QG�*B�:�Vhk)v���J�L�0��83�hF���a2'g(ZVX*Kl�ll�h4(�u�խRb�{;M�j�k#h���$V0��[,���ҝte+�Q�H�k�!ee���6da��faFe�5 fb��j�g#t!4���&R�ؖU��6A��k�Sm
J��L�;\�!@`e���f�z�L�37u��B�ͪR�U�h�D�cg^˕z���yV��m�t���E�k���/U)YKn��5�j���ķ-L�M6��4A:��j=��:�J#L6g���7Gm��EX�6
�\m�-Lk��L���4��(��ʪ������\�uc����ZyS-�)5	B.��U��F���/�G׌�З�70&�̺�O��5ѷ)J<45.�琾�o2.�k����6���-�q�*����5�l�g1�<�<��,.���&��.����]�x"ٝ���[�jy��u���e����8�ᓳ�@qI�R���{V�Fٳo�h��p�>��晫|w�{����ooo��۷�oOOM�B�U�q�f�yyx��mi�vd[��{������$�$�1�����^ݻv��˷�����f(��mX�{wy�^����:��|�F0;G,�����ɲ��6l�ɳ�����9v�X+4��/�/V���ЃIW��[x����y��MVrͭ�Ih�%B����^���(�im���L8/?/����o�_�͞6l�����<�B�[l%A�OEo^�ޛ���׫��a�q�ԕ�{X=�eT�����+#K�㳎�׉uIh��B>-��F�V��Eu�MM@��[G2���	5C{d��-m�6�oy�O:��ӻ���;kv��di�3vq]2�z�[j��D����ٷf���yt%��׽��\�'l^���כ�{�y��_O{�o��M$Y)H�V�Jt���nFZR�	3nk�S��w�׭kYe�ݻC@�<z�ٚ���L��۰�ok��,��P�T����I	��l���w�=��dA��p�秫��I��tu�'}�����k��K-<�/kZ*�%�i���w�RG�Q�"D����fB\����m����[�'H>�۳��BD���z]n���n]�L٣nt]���	u,����Y�mob�e%u�7�r���BXX4h��]bP�� k�Z�4�	i�5LR�WB��1e�iaLXա�2\̙�mRR&���,j���β�ڢ�1
�
�uۈM]�eÝl̮i�L���F"���f�ڎe�,�m�����Fc������,K���2�d��u/K�`��F���{J�_;��h�K0.h�H�2ԕ�YW�!��Z9��\�4bXb�s+Fӭ����&�K�Qj\�u(Lk��`��Q���$m��(�5U)�����H�3"Ŵ�R�lI��%��I(G!�B1�4��Ֆie"��X���K�F�)le�),GPcJ*R����h�Z$�5�@�YZ]st9��8���k��)�2�CIf-�k�%�5a�z�00۰q7j��&�f����T�6���:�B�;X�4�ha�vS6']����e�0n�#�����p�����[I+E,�w3G(é,.�	��Ye�M��M��p��B.ժi	C%�5�:37+)Ӵ ��c�
�2�T�j�����7��!nfe��TÃ��e��ۮ ����-�Pۃv�5��R8q��ΈٮPtb��n��	��R��[A�clj����C]i��:�ٵ�6�ؠ��5�	
��ѓ0i���K(�&�t[P�m�6Ѕp�	���@�`L,�{2ͦvg�'�-���1,M64��abk�9�f٠)0M�i��(�5�B[�J�8BU!)��A17ZsC�mƉAU�n�8Ψj��R����`L�L.�6SWmikJ��m)z�b�)f���K��[T�X��]�tWZ"8��s� V�XK�F��}���'w��: XkThUB��,��z��-IHT�R�D��R����-K�<v�{1�O+)�ډ�RXƲ�mT���J�X�ڡͯR��Q�"�愼p�J��F��ʱ�ZF�e���hЕaj��A�X��m�V�*���-*$`���[��$mB���+j���H�U �xc(����a]p��i�O����'"��A ��p��mRtf�[Am���������	gom6 X�N��^/oO �>:Mr���.���K��{5� }�Z���̲��@S�a\^e����l ��C:ݟ_����/�m��`����PҬ$J���Iܭ�@����[�m R.h�~��?˻�]�}��y��؂	� �Uǣ���3O�!��-p	)�C�T�BvtK�٬�� �Y��ɇWM�x�k�v��'o\9��ӻ�����0Iٚ��D+�`��Z�0^8:��Ii�.����JFO�u�㳷�3�]�N���< #�X�>�k�9Be��8SG.�$�^@�I�Y>�-�#���',˰,ѭ��{U"6����W{�{FU.��iK���	�;�	4ﻆ[}��W=�{�9g�ԛ=���l���Ȥ��w�C�L�S@��>�HZ����Vk�y�^������=�R���,if���O"|� �[�&"�tS��3���#V�$ʷ	'�z��-�X�������)ة��`�k^A��y�j�s�׎b����m��$V�6���@���c�&�뿤�O��=��PS�� #un�'c`F���y�$�䧹�ƪ�G�a ;r�ik0��J�j-nE�0vgf �V�Bvp��ٴuN ��`�$�	h؀��)�2�6�`��� ���o&gD�P�����4S2��:��'}�� !AS��;�I�5��\{֐�3�L��g((��� �����q�^��q#k�*gj��2`^���r���c���==_�^������C;����vs���b�v.�l�7����4ۗL�$��6i��<��f`��"�b H2�8 �=?L������,id����w�Ce��!�D���$�h
���$O��nB�w����:�;�M��l Y�� ��� �kCǁj@��ƚ-y�<@���W1�����n�DI=�j�H��N �c	L�Ƙ%����n�4J�%�T����#y�3G&Le���c'���ܸWrS1x�����@�n/"�Q *ہ#|��"*���T�k9���+�LYN����@f�� 1�dֶ��xa���6YiI0�q>�%�
�]�>65��{�C�a�	�o&gD�U r�@'k-��3�9��&��Hh}q ���	����p軧	ɐ����1��[�L�w�჎�����U���Im����#��E{Nܗ�sS^s4��Z1$��r�Z}�5�������l6�!�h�{�}՞�,�<�?��Ԩ/�c�|��6��7�U`b�#<�v^@;�7�H��z06����X�p�I"'7H�E]����_Ʋ��M��;�I�RY��~Σ�C���͊ӨD�Ŗ��T��&�D��S�)H^�ԋ��K;�����k�1m�q E3is��}��"�ȱ� E���7��0���U�6AH;n��q���y�wo����[o@Gm�� ����X�K<��JN����zY:�I&�irA$=Ќl��N�##2�x��g.Ha:�So�X�5��������&P;�qf��'ĂE�Ypc�ș��m�I3d<�U��;�� L�;�dW���	ݜ'$�ӂ<�$�*=f$��pH}������f9�����ws����Qܛ��{n�`�f�W�yp��Fr�~]4�]�qZ�A�UG�Bv�e�Ed��~��r��rӄ����)����v��M'�����7,��wWWL�t�D�˥����y�s5q�4-�9"Se%��02�3��v������l���dE��7i�Xm	p[�ٳĬ��0kF��Ֆ�mU�v�C��-PeL �;1���&�{�8H��K�X)���z�s
b�3,���2bU�[�����i1u�]&I��h�،��J*�V�F
�K5Ү��b8M�L����m35��gB4�ZEj����^i�ZKt��W���H+����$�/��4<S0��s�M� m`��G#I� 6���������"�5V��Ō��	��O��!Tl@�A���z�.��D0O$����靉NK�X"���$���j/;����&��V��浟�k^Y��^��x��Ů���閬��L�&0 �F��K	��3]Ņ�e����o;�$6��(���p���0p]���4l ��[��Z�a�b�G���i��׊�W5�
�n S@$[�cx$����ޠ8D�qt-��u�qi�cG&��R�`�F'{Mmk����7�X�;;8LN�5��c&��sm�R���U�03SQpI3�}�=����0�I������#t� b��'�5�LKO�,�����u�D�m̫���> U���S(nњ�s���S�lmʳ��5^��d'�ZN�ze1���sv�A@�ʶ�r��#�v�rSN�`?`����'km�Ɉ�t��e�����A��q���x� 5�[hgt��NK�h�y"�v��Y���"�y}�	G��ہ$�6���`�,��A>-�Q���O���:�gr��;
m��I4-.V���6�`�L�ωo%�ܸ��r�Kߖ�پ�{�^�XPX/0��X�Uέ��t��Ř�Kj:�O��@a��b�??e����)���b���M: ��x� �6�K����q>U}^@;�t�`�V��Za1��- Y�g�؈k��1l��Q[���$���I �#V)ձ�t���`A�Nd�kAӺ�]��-Q����/k���>Q�WoԦ\(]�D+/WM��bZ�nл���Se3jȺ��"�PZ~�z�}L ���ܵ�/ះ�	�Ң֏x3�8�;��<�D���Ã��'�m�8[��?t���ظ <���RS���&�S���6#`g�m�Ǐ��[C��v%78aÐ@7Q�C��'����ͱP"'۸���J���N�'��2�t��ZY��fr�Ү	���#�3���
���-�;4���?a�o����i��	���`��lk��kY����#zv��A$�6�h����_��n�RT� tmn��� |�|#�Z�C	�	 />u��YYȯ�D�?��b]��ɘ[����&,�p����|I��x�M�����A�X\h��>�+t��d��U���(#]��ݖ8�F���� ����A9�p��"��Y�r.VMoRh0��1.*ܝ���ް]~Z�c/g�<lo���gd�����OSza�m������	~�����a��Ԋm��_A�-qH��x�Ƨ���e��d�XF�<�ݜ�ݏ3�]��A��1&v<�)	}���mS��$��X%�(��mA��K-��e�"�<�����6n�	���ߦ�t$h1��@ ���D�w�L��i.
񶍏A�%ɲ��$Ą��HY;�gٹ��SW��Eӝ ��� �B�f|U{N�Q��`1��ɓ��"�����o
3/�X�1LWH8D��O�6�A>R��g%Ӕ��Զ�d�^E�IWq���z���j _�Qz�=��.����h�8��_�]X圱@j�1� �N^\1�^�5O	���/[�j�HV���y/�GhM��f���Қ���p��]����v���hl�4L���>2� `9❩"
)/�k<��|,�p*�Ho2����"����9�ou�F���fŦ5)���k&)[1�Mv�+�Z��� F�%`��!���lc�e�/9�AK�4��m�b-E��3S���6��V(]�Q���
��cpb�7c-ĴB<��c�ɂ��L�l4гn�e�	E-a�2��X:Fl�K14��Q\Yc�*M��Vd����2�.�F\�T5K\�M6+,�ʦ����X��߾�}�쨰���'���Z%�'q���ƪ�meМ�2���{P�-��	"j`t�� ��L:^����5'���Ql�6-9�7B�)�㳈
}�!x`��O���E�ѹ2k�p׾���PN�� �N�%Ƌ�D��A�H0��y�3�F�4�!y H�p |H�z��:��;&S8.���73&m�����tT�H$��<`H�I��pP"�Uش�X �m�O���,�b��A@�l�$O���K	���XviFz��U@�4�-Aب�CG���|��~��=: �a�:����4�L.�[[��L��B�]���q?>~���LU����� 2�-i� �q�b|w��_n
�����X�i�
R�.ĸ�wQ	���w�Z��F���3lL��)��[�����=�Ӳ�@Nr6��,�v�y`R���A>��j��0=;QZ�
l�^����Q���.r'b�v2i�g���f��D;�El^,8�5��S)��{֡MV��]�rN(�ǚ�"�Ll��+��d��9tCy;Il֨WW��k�'�2���%H4fDz�ղ��Pud��/OY�S�����;��L����u���	 ����i�KV�Y�0�֪��	-��
�ف�7��}ߑ�a�~H#O���M��Je5w<ʒ�m��uz�`^%�e��-9��̓���tag%قwE�^'�H���r�\C�X#Lg��*���u!����9b�ӊ��Ǐ�"-�h�l�
(RkX`O�"$�͘�������ȴѢ�'xp<X���� ���9�3�HSS�D=��5���z�W�d�����ⵚ�a�݌�r����N���p�=����qǬ�;�x������C��}�K����W��́�=�<���y��k�l��^�S�1��p�3MmK%/�o�qg�o�S@��7b��{}���nL+�^��.ٚ��l��x�� �e���}ܼf���~~U�/��W&���s��m�U��Q��]1]���;�)�w<��N�6L�tM�S�o�=��Onw����^.��GH�w_:V�o��8y{�/@!{㻨Q��=�yg,��v<������&�~�+�qr[~e�z���"�5Dۉ��^�$�GZ��+[˝'ğ�kr���=������*�����j	��|���㱅�˸lf%8�����ls��\�Z{��N���綷����*g$g����^{�B�Q�����9V���xus����r>ط�#u��;���1oSř������&u�j���{G��7�:;7� ��p�&�s����w�VNd���>�~�x�b���^�]�7u��y��5���>�6�Э�ɜCa��=ؗ�6V{��u�=�б?Z��\�˃�_�ͻ�����7-���Dut�;q�IN�8�0��t)��p�\N�I,w��`�����?�$6�Ý��u�aW=�nЉ�潎�4y�uwb���(��<�/c^���|l9�q5��̧V͏��m�/�ֳԬu��((V�6F(t�|.NPIHJ�Y�v[w���7:�ep~��٬`~^�{��>�-�i]��j{��oo�Y蔎��L�d�5���y���$����b2�sV&�����>=:�����o����Ή:zzt��HB22I�Oթ�'"䧙�H)S��r���~w��O��|�;v����������T$�%�c��r^v(�(t�&'h�v�N�r�+,h���0hѣF�(P`�� ��A�]�~<�ЊJ�8�c.�v��r��� �|
D��,X�cF#E�4hѣ����{�B���ĭ�v���n�:۶vD�	�W6㮒�D��l��e����޷Vu����s�Y�ݠ-���M���˷'�Okrȳ*È�N���8�PQ$v��9�N���	۫��\A�9EmnB�Y��c�:�unGvV��Gڲs�(�(���+>���[�>����tE��T����V;k8�@�;2
*̈�I(�!:R̶ݖgd���'PfgZU�-��B���5��	�,��ii�����T���=�C��
\��F��d�����FKˣ�ތ{���v����� ��	T�C�/0���߻�D�`׈yx��|�t}�{�9�..�{ډ�6!aa�kؼ�9�W=Þd<.L,�s�I��^���D��y��X��x<6��> #�p�S�B��qי<�SUC^gy�C���$����� H�l;a�.�X>�{�'�>����/��x��<۷�wtw����W�h�u��(`�ԶYKGG��X�ö��H]�g8j��� Y�w��#�$5Ci� ����#�XR>����ȇD,R�(A/}�X'�&�g�#�S�Nw޺�s�G�Y�`�h���|�2)!/�ɱŜ��ء~��R���a��ŏ�x�"�F��r���dsI�E$NC����w�p2,K�,[7��p@��]�ߛ���ƭ��{�E�zAG��X�س�)�8���� �����)mR���z�Y��A���i�Xqיw��5�:�!�7 욎��a�}�<��[�K��no,RD���sz��`�v%�x��>�#�ZH��b����ń	��|q��u�,D,]�̰N%�Yb��޹ױN�met�i#��:�C[a��y���Kҹ8��3-՜|�N�㶾�s��[��%�� �0pc��g��	�o����s���a��ؤ��K)=g�&n���Wh�w(�pȳ��=l��<�q�� �a�W�i��]��3�Y�o��� �)��g^�`H���^.���������X��3q~�M��$�3�gD�am"4Y\*�F�-���G&T���F�>bߚ}�;�ti��d�bgZ����I�N��p�,���,)�Z�ڧ14��9�y=��1��F�;�;��RE$`��u�D���<�}���Ma3]���`|S�	>}�}�������X�P����k�x}�D+�(A/��8��,Lbh��R�ί�99���G7yU�!�Y���@�@�B�[��ե��Y���ē|��;��'Lv X�a�W���8bsN;4� '��}g�q�Ox�]޻���,D�M��d^�cb!a�W�j��QṦ�ᜆvr�h�(�t��,<�Yϗ^��,گ�JZ���/Z���/�Q5���k���	��>Dw?\1Y��u��鑍*�<D��(A���N ؝�;���Z�I��8�%��]�W�'1l}��V�\x�B�"�
�p3KG`��pB�o�{�E$M�lRC��;���y%�`�S�yǾp:�Q"W��z�4�\�)�1ƅr��ῗ������&��k�?�\��aP;��w}�O���]��T�{�%;p���(���r�0�M����z�����|6ts��`楙�8��i�Qn���pZ6��*���ňGZfD�4��- ���м^��r���ڒh�Fh�2J�e�ۍ���Ytc�;"HH����e�P��!F�4��u@�WS��#]�4�S`�Y�6�f��c��3�)+�#�eR�t�v��ܨf�� m�i��A���e\��kz-���<�ƱF,�n�T��������
�&�3��1�y.�������JL��k�O!��/���X��A0uD[ι�Hq��R��s����>�S��T�벧��g��>��e���,lB������$*�t
�F3�b�Oϡ(�F��xIb=���4=�ه�[��p{�a3Z�,RE$�����|�s�� �<���욁�E�,[�3��Ǘ}��w�X�`ؗg\{ԗy&L�.����T�9��t9"s�,B��=�^����#��
����LYޔ�My�b<�(K������$RJ@��x�XSZ�e�eN]8B| ��Zxl��M̎� 1I��Ǵ��RD�lKߞq�#`�D�hİw�r����^<��q��{#���l��>�wP�<6�Mb	�9�썊���(�N��xs5������N������#Iձâ0��H`|#!v/xA⅍ 6��;�lH��`����G�� �s7@�0����Y��|��5rb�kv��0���
�d�]�׉�]�TXC��߿.	�l������I���49"s��Ut@��|޼�$r#!�]NِMw����X'{�o~��x�M�<�7�����D��!����n�b(���&���&,��xI t��$ ���<����dY��;��P򱣮�&_���5kƨ�2[Fm��w�Oh:(m+�2Z���������ڑ�^*Q}j}Gm¸]^f�<גXi=c����٨w��Ӳ/0.��̊H�����GPX���5Q���X�,RD0�Q��1>���t'�<$�#A &	��u���g<A:	b{ν�	�2)"��Fks� ��P#�$���Rs�@�� z%S���f8:k�;�L�$˵������"]æ�T|cZc)�5��g��H�u7K�z�|,�Tx$J�~1	�uyI����U�xA4Hzy�ey��H:�ċ���N��pgO� �Iyu4�y�����K���|�҉���H$��}0!8L��4r���eC���|ewJX�}�}��8�h�`�R��eBͷZ��(���X���4KCK'��������5�Z��v� �%��\�HKC6��)�%QŢ���;�l�z���`t�[����"�K�&��/��IUQfB���_�=|/�4L3��B���%���p��[l��Ҥ&�����R ����X^J�M��fgE�5���b#�`�z�2Ҽ�|�9�tC�B\�lSu�Z.�E42�8%��q�Fq���x�����M>���X�پ/A�W���/X��/��_���/��N�H��r�mkJR�V {����$�H.��I ���^�Z��#�f^N�!t.�!t��;v<���9���S$�޹L���o5��X�6�l����=�%�q����W�_IZ�w���1m0��R	Wk\H�탺�>˽���A�f��Co������D��>C7�r�%�T�ڣ�����O�!��f�.�WF�)C`έ�ʑd�6֩-v.F��B�|�pX�/
!V�v�]$��`�ۓ[�	 �Ki�倔%{w��+�UN��m<ٞ���r��g�M����r��0r�����!GKdHd��44�*��\���!�NBB��w�5���Zֹ���i�j�}By�g����0�BG��u�)��S��H�U�l��2>@��k��I
f�H�+y�CK'q^\Qra$�^m>�|�K;��H^KpM�K�fwI�U ��N<���Z�/Z ���m�i��
��^eHI$|��~:͌��Jh�C��q�*�%4e>�=Iy�ѣzIbi7�$���,fV�'�Kic���G��%�]�l��e�O��mkiHB��%���H�:٪e)�l�J�v,̼���!揞�Y$������̓��堪��s=(�A%{�r���y�8f:��<!k��<�=�!=�؁D�;� A*|eqb$Mq.d�a	^4��]�x�0�ըm.q%s/����X�-��]6���z|Ҽ��V�\K"W�vt'M�yv>�Gʛ����2d��� Rᙇi�I�%;�`�u���A-�Qz�Fg������G�y�`W�oos�)	Y�"����Ke�K ���Ŵr����p�N�����bB:_"|��^����E�����:�b�e�!����^��M��@$w9�D�$�>�`�`��xߒ�k�����4���h�e$��^@�	/$��y���7�{�Ē���2�@����Vs�K�gg	�]���^Iy*ƞ����ћ۰�F�{ޢPg��RA ��u��B+���Pm?^nV5�)"�����v�Y\�L���u�N;9��,bV�ͷY��Ͻ�`�����C���;�{��7Vo�=��� ��-�]rv�����Rq�qfq�σ��d��iJ!JUR��9:���d�{F�,f��ZRe�óHź�Q-�lIu�����,�	a`m�4l���l8i\�E�\=���Sh��+nva��]�0��B�1�T�rR��YR�U����3 ��X��]X�p�v����pQ�h;\��F�]b�m%0�ଦWj��vmrXn�թ���|��4���{ek�r��fZ?�;�O/�bxƺ�l��!�B9��(����]Z�e&�8�{�����f!m�%�{��Pdk�#`?��3$����	+ˊ�d�w�*�����v�ԢH�Ro 9lA��\��g.����Q�<�h������
͝�1L��� �z8��3y"Cb�S*<��VWb1`{�saX��2�ĝ"S�L�+K���2]MW!�/"Zo�^�o�"zz@@X	 �y�[>�i�y.��R%!��l��������7)n�)�3�S����RA'��B<Y���z�$�ws\)/.󸉯x2��C׃�ưE0t�p^L��[%zL�H0�;��lPe�f�a>��-�.1�h�bKy���%��T)��|P7��n6g���������7����9-���S��X��R牋Z�	^K6
2�v]fֺ__>�6�b�g��p`6�B^�fK9�$7�&��_5�  ˤ��<籸ϡ�k��V�a4A�vI3!�|�O���H%kE�l�T�w�st��6�nCB-A�f1�iQttX��v(c>[̪g��Q8�~�-�w�ۓl��T��q�;��x�^���Oƣ@#�R�R�@�@VDdB�c����dm�S(����p�$�����GK�4��=[�bpc,�2vt�U䣚vCJH�|���&�����ʱ�o�_�A#vӪD�|}��p���`T���;����l����jrQ#�+�ܕ�n�iI�W|�*@J|�������٫rjk������y�M����!ݦ�-���ٌ��n�d�K�R�P} x���bo���P�g����dF��%ʥ���O�}L��V�3`vg�xd�Y�3�اpQj����kh�X��ѹ�j��,&"v�Ժ:�>|��>�)��]�} ���l��$�U��CA$5��B@&���ϱ����e�b�A��|�f��[�wQ�r�gr�ý
<�����&ƭc�/���+�a$�_6E�D��G����U�����>���ọ���y�QY�"�X�j��s!���k�D%�䒚���4)j.�kzb`#��qv�,@�B�`�m��dPʋ��̄�d��B�9ʰ�EDU�>������N}'5��?xx}�����)E)J6)"+"�<5��K�
7�����o8we���=��rȦN�=Q;^B>!�Z������^I%��6��"�\��f@d�*w�Q�}hVB��E�
�*A����R���MiLQ(��(KJ�;�P! �K�O4ډ/RCմC*������>�>H$]K[^���ə%z��M�f7k��������Іc-�Vh�S�6F�5k�������v�f���t�1��"�:wf1��bc�$���8׊@��I%�מRD��4�v�i2�߼%v5���	-m~��0��\5�)���z��>�w���CJI���Z1�._Ow�"!f@�&�3$6b�}W��n��'��b�az�Ǉe��jH0�X���w�,�N0�W�����ZR%��f�3��WL#�L7Wc�x߻��g�Q���y�"W'4�&�fe�A���תЫ���J�xYI��G���ffKu�����?���H5�^��&R���|g������EF��E��=]�(0zFf��Խ�u�Ο��7��%>�;���G�*Jo��W:�S��9��'ߊ�B?
ֵ�( R�J! �T�^m�޻�rG���'��2j�h˕�%���V�"/�׀��{rf���ǅ�IKN�����s�b�^(%���6H&�2�h�A��]��L��z�K��ܒ�Tծ���,�GK�E7:D��v��%V�u{�1ɝ�n�v}P I�N�ܴ���]���Jy���d,o�5�6J��$�i�3����!ӺaJ9L# �s,��}�"ǆSK!/$@+5���\a���祙K�V� ��������:ǫ��t�l%�2	A"\m�D�'�(r�6ڲZ�ǅEr�$�!g4�H9s�InM㐂gd�:�7��R�T��	�y�aM���H%pي%$�K��zC2Inx�p���l���Au�J�JZ-���8A�/:�et�I�n��ϊn�����6y+�P�K�WͰ� I͜�П�)���<���C�KkTSdUݦ{�<�k޿�;�
��z^՛&wowm}�AL�Қ=�3��L�~a6F��F\^��zvI��y�,}��{���4����q^����r���}�{�L�0L�y�Ώ�'�����_1�w���O����__1V�����|������j����T6�����ԯ��0�Μ=��_5�\�]��yw#w{��h7�?M�f�zl]�����g� O������F�ީ�Yʒ��y���������x5�i���b�����Ӭ���◼��Fǫ��g�sx�"מ�����xk��Ȝ��]98�eȥR��^5���H�=.�����t7�_�Kz(��sU�š�����CX��١�������I�s�f� � �GI�M/JNK�%���2��єT�D�a�c��z���5�>��,��y��'{��v�u����1��'sD�Z���q|���7	�n�_!�7�.��L���8���C�m�A�r��μ�#<�v�>�����$���qÞס��M��]&�5'���IЇx��>3�Э�{�`�{豔�|�ib;	h�g�v��F�c�y�/a���ۼ|��׾��=^�8fS=��H����v*|��
��HV4=��J���cΞ�}|WOX�������s���}�=��@�(<����Qf��y�zzs��/��vg�S�`�x#�F����8�j��˦�����n�6� �ON}΍����Mur��`U�� �2Z����z_т_�O�a�;X���b���C&��=����X����K:?)���\�m���c�G9��x��ĄCzae�D��F��a���R��-�Y��Y�J�P�����#�ݗgtS����$�������d�"꺁6�����zzv�x����Ƿ����z����qH_�yd�������g9"J��u�v�����zz{v�����ۮ����;�k�e_:ܤQIgb�q�����G�D!�ѣE��0`���,Xo30�����M���ӎ++me'D��A-�:ŋ4h(X��4X�a8$�A�H��W�n�u�\'g[7q<���V���f\GI�Fٵ�g-9�,Ă(��Ye��G^�ݒD�Y��,��$Ⲱ�=m�d.�	��f.���v�kmm���V)��㡷nP�PGE��ݝgbY��e�B��)���YtP'�� �$蠊/�k�v	��Y�qx�-�fuZkc�M�5�b�3V,l��� *�CM]5�!Rڒ��.�!ftƎuR��c̗*�(9�6سgfZ\� �%�m�-5��r,�H��
��GTS"�k���Zl3@%��#�f�Wb`��LR�b�D��l��4�B������b5�7,���M��XJ\	1���vi4�%�9��#G��.n2�3u���ā�h��b%� :������f�h���J�X�TIR�e�$.�ڃ�Յn�l\J���B*��LB
u��[�U�)v�l�W�6������4)]*�`1LK�C�E�qqF%)6�LAs��M�VhC��y���-y)m��(KYF�J�W	Q��H[�A�]ei�YLA�t.�\L-�k,�˪�胮rՒ�)	I\ ��\��]��M��Ձ��jVX:rm#4&�E��0�e��i,S/f��/V< T�Ms�����,n�� ��L�0h��⮇2-�D�sS���-\�k�8-�	b�!5��3aM�,�Nktk�ٰ��q=�����#n�	���J$m9CUM)�h�SeLuZ�e�	qF�-�kkZ�x�DF	i*��Jkqn�y�1�n 3m�"���ʗTZ(���m�!^v��yΙ��x�a�vL��g�z8�]`�MQ�mvv�V� Q�f�]3s.qu��f��kEv�mx&V<��l�fm+�%&6b��՘1!4�����٧i��Պi�-�Y�WB��M�!�u֛����vհI������ ���Ŧ�Q�1a��M�7:"m��Ɇ]�®�N�͘1�[lԙ5��r*��L�1�m-�D��u�T�sv��xueIX�uAqJ���j�Z�Gk�)�l�QՆ�%6f2�#0\if�8뙣r��3srk���4#g��e��ƶ��X�+���(����Gm ����`�E[#Z�X
TP�*��"� H��+՜r]k�d2BZ�,d��I��k\��٨�y�M5��0�^�3B[��,S�n�B3V�X&�7U��[t�um��h��2%��Itt 4kci�`]e+�f�iVP��b�!Ks��fcK�"��� KvȖja����A�u��B�l�&m�nh�e%3P���1Pf��n��k�{l��H��шa�j������G���x+�λ�+\�0�jE1�J�+��	�e�;sl0!n�6�y��'��Z��w���<}|g�&�L��G����A$�C=��p���ܫ�|�+M��B|��Nr�Cl(I�@-՘S	grABզm� I)���W3ŝVfSn�iA$����&<KZ�?����c���x	it��d��bI#/H�+���	��ѱ���W��0�	�R�mXg��)��|�ֺ��+��k�',ă�5�I���m(湣j��!�
�^I&u��	$�U��	�$s�yx��N�Vu'��	�=;B&=2I�x�$Cg�b���2�$�ƞ�ޚ�e�:v��%�oo\I$�
^q��"�D��<�S\8�/���U2�6�|a�yMM�k��L�L�5��,�-66T�u�Z�i
���.�L��{���>Љ[1=��N4I�RUͥ�$�Ky痦R4ŉ8��i�%̗s��7���D���fŞ���i�$4��"�k5|S1�C�8�b�I��iTX�y��qP⥬��:3h��q��7U��U\w��ۖS���:>�>�t��������io�=~5Q+Z�  H0�UJR� �H!nq,��W�o4y���>�U��y?=|�J�A&�:ٛ<�q9�p璑a]u�]�P�l@ng9�o2$�k�[z�I�R�l���'���S���,B-O�!��B�j�C{�HT-��������3ǧ/k/��۵��Y^I%�b�I�6dG)����火��s�o2RH-�lq��ӂ�$����/13���h���V��O3U�Z�zB7����0�Ǳ�P*fY��`%��1V��/�n���ɶ����<�b���l��`h�*if���sd�$atun�X������$��1��'����D�ӳ�T3ws�$�v���duش��j$kͩ�,�1���8A�^V��gļ�QM�$vWzF�=���f���z�$�	��D $�{O{k)��$ߠ��`�6�ŋ�g�wiG5t���2U�����Ļ�������8�ۄ����§��d�H�#��+R xyV��s��Ǟ�dw��=�|���u=�a��]�/���w�N��}K�|�~5[AF5�`+"�DJR�� �"��t��r|֤���R%y��m��	/m��|	�r��P�@R�\6����V�$���>JI$�a@J<�M��lq^pVz#.`�47@�)�!Zfo&-3!s��� �Ir�%���w�V�b��H�-t}�a��[q�O��K����֭[���q�����;k�A���I�� �@�??>{��I���{�l�L�� ���g����!��`�9�w_����e�C�r�d<��<	.�k��`�ë>7t�]������s�6=U���Ko	$�!�T�\��2i���3���P}��c��91p�,]Ux(űݘ/"@�n1�	y$���W70[����RE�f	.օ�D����R:gI�� ̝�=ݤ��X�|T�d�b���GǞ�'��S�#��K5������~%��Mͧ��8�.�� �.9�v�v��N�8��+}OM��S^é�۳��:�?	c�-~:#�x�"G�U�V5��(�AR��`!"������μK�$��:`K��P�� �n��,����54ɻ�Dn��o� ��q4d$�	�@ra%ෟ�Nz���K��}�
��'Ā�9t̙��V\�7;R�����nr���h�V5���VlLm�����g.� ��,�h��I���z@)	7i�5�����J�9�f��,�⼗�z�2M�!/\O=j8�M�`��}~t��%-Ǽ�y�MҲ.��o�$�r%��H	�!�Ʈ{�;
��a����I�x�&r\2��`;S �D�J�����^o7�;��b��dm�\OO�2A{o�@���Su)���$�!t��jb�&�2x�b�����c�F���̚��!$�����L�|{���n�G���G�� c�s���� ��Y�=U�(�^�d%׬𕌎�s���� ��v6! �*�%_����XoL���:Y����s(�����o��pų_B��Z|�ɍ�L�]��-	\�5��X��:"�<+�_�m�����0Ɇh��,��!Md�R��"r�jִP)J(��x�q91���2�]t�� N!u;3<��H��u5�.2BP��h5͘�:Z[h�A�&u�
V�4�3X��A,Lj�#jb�lBS6��310�fǘ5wjZB�ah�[1(�R�M�يD�@�ZX�2�g+H����)������`�*M-�u,�5tIh�`��%���^Ή��AZ]B��&�mp�s�\�2��kJ��t��T�5�a*p�pM�j��\F(y���������%|c���$��]KM�Nw3�H*��X{�h�w,(���'����H8��)�3�r��W�ݷM�ϒ �B��n��y�M�H����RL��o<�D��,'�>��C��j�4o|���y�:��	d�솕����f��xI+�y�ҩ~�3c���	$���~�2��"ß�	1�ړZ��w_���y0�gۼ�c�m7R��*�^	 ��������fA���C�)��a��jb�&�sv�u��N��L»ODl&�~rh窐�@I��s	 �]O�<�����?	�o��� sij�lp�H��!���Ƽ6�R�q�E�_$+�����|�,�ř�>I��) ����rI��7����L:6��h}��h	�SI^����O潫�0.��,)PM��!$�l���Z&�k���5�Ky����a��驔>W<NSӫ�yV��jc�SE�h�,�=ũ��Ǹ�f�a	����D�	��u�i ��HDy��	4|B ���0e.��Zנ���kTB��JUK�U$	�j�A �J��|I�����$H��s�쾻])h�sGc��9v�33��V��"PNm�Ȁ���ul�N����z�W����U�<	@`̼�vC�؄�ǼGRL�;佒z��rÂHb�֐A�qٔo3�Ov �o� $�7���9R��&"�wd$\e�� �l�\��ø-B��C��$��J�����=��ݓ1��G�h$}N����G5�ȏ[pgd�cܩ����Yy���M �T�͎]2Lb�D�.꒗m"s��(v`n��XM��!������]%ρp���I����"ĳz�3�����e�A��;w�5md��c�,o$k|�"?��cq&�Nј���0$��g5$3SbO,��R%v����H����	�PQ��[�Y�D?C���������v`]3�XK�����$�;M���@��Cj�tf���:mᔈ��޹��=�v'����7�x�.��9r�EJ�����%p�9H�z'��n6ʙ�-���g1Pfh��cV�u���ƍ�!��	 Z�ݗwR�캻��.9U�D	 �����2|-�_1Z�P�b�	.n��}+����c:r嘻��]Tгt.v�c��u� ���$47y�~OR�+g�����;<�\� ג��4��d5V��&�;��ϩ��m�PJc��w'��	��fg�����0ߧ�Ȕ�ւ�fl
T����!�m؃��d��;�LZ��
6Z7K��k)��xtJ���Vͭv��~��~B)8p�v�Dpm蹄��S���,I$;���"�"0�B��m�0�^S�!@Kg�})
�8��&%�`�U����J��q�.�D�g6�����2-�g�i���{�g@g� 4k��k��L^����O���/Ēz(��(3;g�'y{��5��4��)���K� ���߰�T/.LrA/ ��y/O����[��H�$�u�.���`శ��_Vk�Q�E�+�C߹���*��� $����

,������OK�j�@�7Md4�Y4~z�Z8�$/؏�#�r��m���HKCcjo<{SDɚ�KSb���r��3�32�����PF�#Z�4�AR��"�H��+ �H��	�fj��3��<�;�'��9r�]��,/��#�$���G�6��]�T���^Jq�ʐ|���s	*�1�~(:�9ub��Ct��^2�3V�5�Gi`��XR��D˥	�I��)���,�G�Fi?>{�/����Cw��[-Ԁ��V�^�<?���	)����PBݝ�ɢ«bih���T,��rFx�r�Ar���
���LB 5�O����R��R`���%��b E$��d���JN08��&�`��C�g3�I��+���fI���]�����-�����	$^UOƤK.�&� �2v,�UI���Бs6ޠ
�[Hn�h�$I�c�M�`C�z���e�P��e$�v<��zۑt�t��aMI��ǳ�̑,��Z��Փ�R�H^��$�s�c�%ͽM>��&�����bZ�^e[�x{�N��3�@�n���n�/�kO7E��	����9�/[�ך����_�R�}�;޺p��8լ����(�o�9���u�"���?�;�_��$�j�`##
U�D�*��H �"�q�5�m�T��u�ͳմ�c)�-��9+u����k��n*Das��릭��h&��u���w2����c4��\��9�av0��T{iJh�k�[�ºܙi��3Ԋ���f	�@0��&��mmfZ9�^��]����[-0��!�unա]�Mi6ahX@s�,2u�6h�YM��pW�U��U�=��Ŗ�kZD4X�tR�c��b%�!�#�q���^p�QN�h�ggN\�.�{�.�n>d[��Cu�	/$��)�"_�|շ��#�R���6w�^w��K ̲�K�1C�$�g`\���j��JKz�9~уi��n53�9 rH$�{L/%��M2��3^�l*�ӧ����y ���:�8w�U�n5��BI����_D��&�znY�5;դ��D�)���Ҫ<|�%�=�"R\fF��t|��g��t �P���I����"]o/9����BZ��e$��n�DI��n�N��!��hh�g��]��<��@.��,��!��b� l�Y��i y�����>��ɒM��~i�.h��x�q?>�3]�QƷf٣ �ˢb�i�&X�=tm-�a@���%_�_~�-�.�4����f$�y�]4R	������Y�*�mySm��0IsoSK	`I��k�wNS�q�jT�:�4�o<�m�a8�/��T��Ei�x�׆T�ᝯ�U����o���/��L�ö�+`�q�L�`�t��-/���K,#��{��Q#�@�D#Z�b) H#
R�D�(*�"Ȣ����2���n��׃Z�G���zy���;�Hw����M[h;]g��y0��M`�)�r^K��.Md<��IW.#`feu3!k�u�Y� ��7m4
��v�X���m+�] �ø-v	�5J���xbR�7��0K��5@�
A8mK]2P0	���\.�f���{݄�����2����p�ã�gT[�>3y�fZ3Z}Q�K���w����+w�G����y���ǡG�Ϸ~����3�[,���2���
��v�-zY([J���K�MH�[�V�,�O��a�}�AFL�:�%3����3s�<$]0��ߣ�Ǹ36n�S��S:���YC\�L��4���x1�9J��,Jl~>�I-&L��W,���`wk9�A$cوD�5x��E.o��,����Y��X5�3��Fbꦆ>�D�N�Y�	/$��� zگ�9.h���hr�}7Y��r��w�#S��I�9g�P==��uK��4�\����������>/vf��T�e���5,�c�ahI��G/���^Y�R��蒭������fy&|�\�oQ�f����7{RE�e'��w_y7:,��>N���M�(�u�t�|�=��#�{��?�S��Ś�s�^�>Z��e�z�s�R'U=��p�=U^���]�	�̕�p{�a�n��7`oJ5x՛��%�6����3N?%���Cn��S�5Ϯ�����~{��=�G�K����ݜ7l]Ğ=�CwGr'݋�P[��^ܾ��|�׷f6�:���9�~���o7޼g,p��7�z��!њZ@�����5��S��;}�\HqQ�ܾ�n�_�z<w7h�~
�����s�3{}�;<�ED���5�?w51V�[��dj�@|�>\ .#�PQ79X�>�W�Ok����t�Z���L�%�>�7:d�tz�K�Ζ$���8�/{IY���{���3�ۛ6�{;�R���[�J-ˊ:�?��k`�Wsɮt�A�ջ@�/Wz���sOxT�~!_x+���f�]ͳ�P}�邾p�ݫ)����F;�����L1_,��<4n�S�|e]��{��	��Tǳ�T�Q_�N��ok�0�˛=�@���cY��_qzp?b��.�U]�N���|�ɼ|{�Mm�l�@2D���� ]���A�kAy�X!�b31��Ш�K�i�0�@�3(L/z��,0���^��BƵ��%NC���,��0,O��=�A�	����d�����:�1�3Q!����/A��@�O�$��BTt\�9�I�z�$# |{v��<�=�v�۷�׷��������b�l�"H�ǎ"���������^��_�N��v�۷�öv��BIN��.N�;G/�np��?w�9't޿l4P(`��4X�a��is�����q���8�����;��"�C������o��N�͛6l�����٬A�V�X4�HE'G@�N%�Q�!�QD!�t��$��q$t]DqI��%yc���~��wƴ�t��I�J�"��]ićI�rq���w"���a���ե}��ܵ�mZGG1��o�z���[e�]r��G{q�γ�u�H�B�>���a�R�d$R��
B�JDY	dY`,�P=�y�~�o�^��� @��$�M��\5N�l$���I{���Y���q�Zq���Ws9 BJ�3���GƵ�����;��Ky���^ $������H8p�X�殊3��'|�&���j��/�D��J"�^v��φ�"�FWW0+�hqea�1��5���3�5V�khQ��`�B�]Dj�	�ne�eXԱ�Š��j����wW��4@���y��K�@I ����N�-���qo�O�I����6`�r�ٓ=T��W('�[wv9�	� YO���x� H
����s��g��r��p�wM�I����U��(9`��Y���'�2^K���4�⼖66-��k�}:�@$�_Lz��[�|�2��lKit�.⪂ꦎݷ�BH$�Is$��z�2�aa��;y��ʃ�_�ܧ�j	��m�cUx���cmTNFV&|QN���u�pFեj�w"�V�Fcw���UP�mMHqF�.�����5�w\�N�H��[��v�VWQ��w]��AVA�YHA�P�B@� KG����<0_z@�v���K�8c�y;�S�&��o���H%s< �
�M�<!xО#dD/"|�s֩�,�W���4��>�	�>���e)����٬�G�ڗG4��%�U��S����#X�T0%�j3������o���A��W�0��@%\��:b�p���;��Xݣ� Y	=�V���B>J�M�Z�)>l�J�`\:>gu�w3�I���Rm�5�3�<��������J�7�!���^QWa��ޗ�18��e�A�N �t�ɟ3|j�J���\����/$�f�͕0��3BK<�>�U�	�$�o<�?�즴K��XS���r��̒H��f�JH�.�x0�I��%�olA�^lH�5�^�Y`�I0�.�r�*�L���3c��vk�z4�^s6'�X�%��A$�yI} ��k��^1u?5I��C;�c�5���7I	5`�,��NC�i"=X�%X��@�aj�b�nJ(3�4���O��8��M�h�)n�,�\��M��[��JR!��J��1���k`!!
TB��vWEW��GE��$� wo��~k�CM�F�s��)��ĵ�]]f��\PaG8�%�qS�D7]�Pe]���0�V���Ք̺Z�/,Қ��M��"L�lY�\�e�b����F��i�[a3��A�p]tDh�J5��k6���Z1��I�%U��M,s��%]����s,%.�`�J�])ˤL�Ef���F���sp�a[+i��k�I����i,v`�-�)3��2�hb��PeE������jSu̥�?�=@c⬒���׀H�/�!�<\[�d\6���j� �����2Ănyp��ؗ��Ldg	Y����b�v�m�`	7/��H�����_�!l�Y�xʵ��d���Kb�>gz,�GkD|�� g=����wsir�u��{ @$���0M �p��ށ��zr��EH p@&��c�W=�Hg4�4�9�C��2�co����͟G�!��6�ıA�9%��^��O@�	 ���m��{��uOMa�ޱ��؂����O)�v�[����޿}���|5
Y�h����Ri�2U�1��Z�j��;8���~O�r�M�\(a�w���=a-�c���V��p,5�;,����#��Ws� `حȢ�L�$�@Ԭ�y��� M�l����4\Ë��
*�K'$V>c��G�z�ծC�>]�-�@�������0	�`=������0���߂�
�N����݋�tt����R^4�&����d?# H$kT�BA!J%�0�l$EI  ��gy�($8/S�SO�Aw&:^�/���:��p��ؗ�H4��S�_�t��1 �jw=�4��Z8P^ �FǠ{9O(%������)�!��Z�w�x �BՋs�t�s˙���3�� ��Zy�=o<�v�(�6�KmFT�0,���,	ph�{=>�cy,;�Nô8��W��Wǆ�3��|\���H[���t�N7S�<g�	72� ��ٓ�X*�� ����O�۲�Q�Ke�G� ����x{s�<3�����������<��{�a}���Ѯ�/Z�b\M�k���v����L��2Pa���߿>o�B"���)�<H�Qp��@s��|s�!�a�P�f��k��tш�"�ʴi�mr\&.�����D����wm�H�m!������	��.�����5�&@"��s"�y3��̝��H����> GDUV�l0�k�Ц+��ĭ,82b�2�2�;}���q3ݸ�c��R��U�NrUd�R��P�_1Sż�Je|�D�+��n!"��F�	 �5�X�#
QK!J"6 �����H�����|~�>x S��a��tY�z��R����Rdɋd����Hw�'�ß��K��
}{��9�>㾯@9D����K;����V<�xCy �lD��[s4������J�wnDKx�u� o�`�nl��M���IH�^#����L��8� ���儍��3�����<�m�>|����Bp���x7������k����A<��$	^PN;�:�4��ֳ �A@f?G�������%�9%��e=lT����	��o�%�Q'����݈�o%����%0���;�Ӭ 2t)C�p����ݨ��H<�pм@%��}��$��w{jXd!\� �~������-��O2}Үf�9��F(�]VǠ"js�$|P����Q�������7�2C!/,�J�ZگFR�w�/i��J���ط)�#�xD4����n+��{x�w���wn������̧ofh�bR-��Y�9�x
��A�B5����)QiJ�bȣ"��������(V��;�|�.ٓ��KȐ~ȦX��0�=���#q�q/Oz�ʈ>��ayo4raѮ�b@  Iд����b4���`�Qp�1�4�`e�*���X�:�_�?��]�v$�g�����)���	 M�G  ��yV�Cf[F讘���^Q`�Sn{�� �]2w�U�}A`@�����M ���zϗ�u�� 7�-y��|�Cf�
u2Ku]]�]�I園�g�v�?��u+�c�yDC�zb���C�o\�)��=��@9&�0u�	���5-�5�lhj g�=q �\�TA$���;)nHar*<@^<۱�z���-�gI'���s���ᜬ{�,Kf޴t���wM�<g�A8�����@#�}zïf���B+M�2T]����'3��v��f8~�w���,W��)/?wJ�$�T��]�t��^oczX��y��2���z�0���d_��V��<>Y��6İ!��j����U�j�"��ΪZ�u�Q�A�t�Vz[/](Ʀ"ᔺ����r�aM6��uK�0��X�me���2���a��Z�q5�ұ��#nc86㴫�j۰1�S�i��������kS�M��lcp4�kF.nR`�t������*F9�;��k��j���Er�6��c�ܗ1�F�vi�٧:&66.���pVZ�UK�f�7�i@�F顱fi1)��%�B�й��U��;��/��]�rY�~�~񺝀 o�֟oK���_4A��=|�ڬ�O��=1錦l)�;2$;<��~�!�3m�{�Q׷o��$��okтEy!����`����ծ��sb��E�` �K�w��Y�pq����@�Y�Ϣ�������I"{�A>�ވ�A<�\���IB�my2)�qA����b�� �%��\��d��˙H&��t�a�	&���;'	�8����B�^�.���%�M�����<�`�k��D �;]��`����������jJQNg�jcvV�a�nu��u`M��\�U��JYf`T��m/��ϼ~�[���O��L5Ǒ#j���}~(���N���<W�u��{1�-��i�p�.Θ&r^D�����yb�Y�jZ�^^Bv��"��L%�韥ia.(X�d��d/_k�T��Wߗ-�u!���@�:�]��a~Am��;ئ4����DI�hء 
а�����I� ��KgȀk��[n��|I�����_4�[{=�ϮG	|�m,��3������\n� A�>.�a��7��3�|O�;�=!O_\{%zEU
�Aؗb�5~A7scov�c�Aه�������	}p�#���w�ύ��/{s��CN��5�!�� Uk�z �[�yw��	��-f�cl��3�м���x$�.�b��\�L��>pP!A�M`�h�k1X*�Y�%�rdi����	q�5�Y� wY'<�;'	�8ފ� ��uM��su�;ܪ�Mf��	���}XA���Kyø)���Q�����;Q�^����By��C'� �+[�G�3"w�7K�@��l�Y'E�g%��ٍ����]r�
'��<���5˛�b�9i?��|��n_-Z�q�"�_n�hb����ͽ�}=l��{Y��~3P���e�f���Hk\�>I�ơa;v��Z�եK[��:���$R@�����ߝp�BJ|��R�Hi����9,��^�莈�-�0���$U� 7�Ϲ���>+/�"����O5��=f�S�^$��x��D�@A8.�ޫ�b� ��	ok���";�-�4WEO�p #]����xv��C�=��@�B@��I��]Q�a�/$��3YP^t��Z<kfŌ��WK���k�!L� �x��PH�+�bA�ހ���2oLwSCbP���T�=4�Vѿ*�IӆgN h��6�Φ|k���*"��Dz�~y>�uvDx�l:�;{�ӾPI`仂���S���O���ǉ'�\F"^��:أ�`�4w1�ǈ>뾁�N���'	�9/^訄˅X��g��(�B���GƎ�y���O~A�#>j?C�\3T�_,L�l�g���L~')�dU��#����Ζ'.��sWnw�k>$w����������޵�<�o.�ï��D�ѢV�,z��e���.��
�*���Hؗ�
U[�郰-�O2uߢ6�����-�ȸ��:��U��w�Q�I}����n�F[��U�pQ?~~~����8ZCm�Z��7BD,u�e&���F�m()�w1(%ڴ'c�E�v.��\X݊1<�$MO\z�a�ԙF-��o���Ȉ�lv�)��⨪����C5b�P�a��:�oDx��x��D.�f�q�5u��?��ڿ$Qe^M�e�O��ry�Uy'�ᐞ�*�d�wk���vD	;S�>Ǜ��Y:��'�S�")���)�Iخ�$���LLם�ѣa&S�"B]d�ܵ)�p�Kذ�K�'ƹl�b��C��i�W�=���� �g@�}<�Ď�zPx<< �����9�LA�w#j�U�uȇ��P�_�����9��Y��7<^sF}��f���H��x�a`�n������0L�N�%d�_S���o;M==��vK����.��M��kϡ���{���������n�>�Ƕ`����O$����9�R�F5���ۗ����7׬O���q������h	,��l���J���nY�V5b}%�)�{#�y���g�]�%�l�����w�sֽ;��a8u�&�k���䷘��. �B��C�$�-�����O �Y�{}�������~���D9R鞉l��ûS�PMs���;<_g��-3��.�U�ң�ͳ���G��f����7��T��/�w�ٸ������2�(7y�z�Ц�� ��J��ǔ:x��'v�������>�#D=�rgn�l�ݞ�+l-%��Xq����d�z��O7�]��7�7X��^�?g�i\��?M�#q���|��GY�<�{��s���Jo���&��i�(�f
U7;�j�P.q�檆l{��;f�o�g`;��v��nl̅m+�3��6x����Ǐ�`�X����N��c˞W�3ܵrNnY��NI�����$R*�)��1|��:�����9�{�6�vw^�8�'���ޠ�����+�]���w��������8a�{ �$��V�满�`�-I��P�����)Pz��	X6�h�<�� �OVG;M@��L&( h�gV�Ð}�Ӄ�5��n�HK����/	Հ�<��S76c$h-��f��[<-���,G߇���S��.Ȱ�V(N����&b@��o�Vy7��6�������?�e���Ο;BB+�������ݻv�������������$J
?U�|+����<q$��Z#!$$�>>>=;ycӷnݻv������	�I!v�#�u@�@q�~�8)Hs�� ����(H"��0`�b����褪.R��H��H$X�bƍ��0X����ÂG�E9�ͻ!OmG�R�')��d. ���/Ź!D!|:��������gO�grH��"Bpq/��G9}m�ݲR�s�H�9%{X��ZqQ!G9��������Dq(䎊: �r�/��x��h�lvc`����J��de����	��!�̶d
s�SL��FRn�\�B�zg6`�rmͣ.f���5�X:X�I�Ǝ�Q���YX�4�j:kp��I�lոQ����5��v"bWSj�sWg2���lfڎ)���A�im�3b��p��[�.�B&ٛ0s3\V�a�D/J�m��k5�ᔔ�s�����Қ��7�0a*GA��l�F�m0�[�aP�h�M��R�h�te�ZB왎XKa+Ĺ����B�,����%��l�۱``�̌2.�ĘY��Ue/;l�63#�o&�	��i��rl(y��pO����v�8i�U����2͠M�,! ���m�����S��$�a渪MYbRf&Z�SPf�XJ!�%�5Y�k-f��\6�[-z��F�j���2�G�F�R�����am4�0��d�b��3XL�-��
�\��p���S-�n�F%�T�#���%t�m����.b�bhY]j9-B���]�bc
�0�0���9�-tbG#��WJ���\���E�(�#�a�����X�+��(�lYL��b�d@#c�Q���TIl���6"_�M�t�+�hM�2�Jꨱ��Q��X�,`Kv��4V8�.����9�C�ɐn�E�f:�w`tؕ��]W)*�es�D(BJT�i�s5�9ݶ�SU�u0��Ĵ��W�""a���g,rh�h�#3��+��F��Ym�Ɩ�2�%��5s+b�\� �l��R�c-���X��;76&�)���5sffR&��+V��71aM�Whˣ���	�Zҳ X6�2�ir��L���G���X�,L�X�֊Q^5W)�[��y��9��&���lŵ�(f�EΈ"W ��Եr��.r�]�2jy.n���fb�f���=D2�x��ļe���$H�jX�,kVŭݕ�[���s�.:��@O}�V�`v1�6Ƅ��,�if&B���P�\�C�U�f�H�њ�^5�ر��JTfslu�`ыu��*W:�Mn�\��ø�e�]b�ns0љ[�h<+K(:&�Қ�ִ!4�k�Y��d1l�0�\�JA�u�������c�.��	V��k5lР��vL8��v�m��bm1SLm)"o9�E�l\�l�Xs֍d��a�Z��+f���*��.0fgh@��[��3�Hwo��L����=H�n��]ο=���d[� ����g��1��]�J=��)e'�j{�}�bu�<O�o$&+��'�3��ZI��j��;�0}~�^3?�{]�)�g$���L��=�7s�!]�h<�z*&:n 'Ğ����⼂^��-'äЂڙ0N��	�Θ�l��6g����2�=�+��)�f��H�ލ����r�t�F��B��ˉd�pS̞3��$q�x�u�E�~����"3�8ώ��h${/�<o�Ѷ]�4�#��^(A�,i��E�C9�liojM*�"�G�u[�&Z��C"�z�j,S�᜖��:*= ^@�؏9�v����f�#�P ����f�B�⏠h1tWk�f8!;@��� ��Oi��SN����vb�^��g��l:��{���[�n��z����?L� �шg��h�;�釩kaB�Z�����N�h!��x,~6�5��
Q)JXȌ#	Uk��k[�P	���y�\v:5�zVV�DP��C��N����n��DWk� �m��nΎ��A7v�cĒv�O�R`��L����	p&�O�<`����RN�)�$I�˾��$�ޜ�վ�������VK�C	�7D7�8t���0��bH=��q�_8���#=��^�	}[�'��9���e��ٙ*Q��`�7�
L#t�u"���ĭ�*[S2m�h[���%B�@>{���pd�pS�{�T�$��ׂH'%�oV<H^ET5p�L��7\�`w�<O����b�S�r^�J���l�p9-P�{�\�^�|�Wl!L/���9�P�cA��׆Im���0)�	�dl>�>4�� ��ܙ5ҋ�Ҁ������Ȏ��7���ܰI;����~�nh(��:�O�����}�Ѥ�r��u��y~�ł^��&���$~5,�m�)R��bȐ���bB��y�ϔ��o��p�,�>��.t��ՖV�!������ ���b��b-x�kz�7�!>d$f�y`�^b�N�Eq��"|�#�^[;,];�X���"Q ͏P�E���Hh����:���,#��H3�ٗ�9 �I@�1d����M��Eٺ��2h�5m�ʻU�R���y�w|�2fp�øF��x��Vr� �A;\�`�4���^���q��W��}�d!���NুT���퐉Tǖ:�����z�	���ws�yI�+�6m��A���ˇޔ�y�8�,\2p���ޥyUI ��y��1=�{�/�[9�_C���:�H�ϝm3y�ǋ\�陁g'ir�o)̀�w�}�J��ԉ3ZaA OgDc��n��w
S��S2�eOS4�[%dվ�9�wX�h�z��xaG�w�5�/plL��>�a��Һ�7�q�V狶�u-�X� BṜg����~U%�bȸNΞ</�nf��W��x<:V��D�Bu�A�ֈ�NA`�����.�AJ����2d���Ğ.0��R���4�G��V�p2�%l���J�Ֆ������o3�b;�%
��=y�;���ח�׼�g����uƄ�`��s ���y�ǁ��;��Y�3�L*���O�.�[��\���<{V<�W��^>���: 4L[n0�vFTu9$+%݈N����#�ھ��D��nab���v�z�����1H&|�;�����	���'	�zr�5+��UM�I���D{ޕ�dCk�A�� �\7�|
zlŶz�`P��#���_@ @$yz^����pBO�a��|C�ty���n�m�u���]z��k�E��:���\�\(�ֲ,���/�0E�ܣ��mH"s(\ikiǛ�˼��|׮�{�ܥ�;>�H9��w��;�7s[����c��}���@FG������0�ĘqlOX���'��#���ͪ�C
е�R�[K���n`�5��h�0�-ɛ �L7@��ZQ����*]i-]F2�k	sn\�:SaT6�k# lk@.��Rn�u��mö�ۢ�L٫��F��H��0J������J���b�QҺ2����P��M�*m��h�����3o��ĉ��$u��Ĳ��aԆ�bV�,
%������3��j�Y��#�B����X��<����3"]� A�7���YE��P��>�@� ��s�'ľ�Dȋ/6��d�����m�`�3Ե�b;�%�1�v�	Fr�D��׾���'�n�D I ��@�Ak�;l�h�zݕ���_��2ft�Hm��_��A�l5��mv|f�X���7��A蝁K8*�셤��Ί|�6#P�6ٜ٨?�U����A>���S����=���F�H�����ٸN.8NȣӵЗ����m[�T0T|O�o�	'�����A���x8��Wk�=GÒ��@�a�)�z�H��)tk��Ų�`���5�JZ:��VK4F���ҳK�"Y�d��_��y��l��	�#���[х��$q«� 	�P����o��U��,����]��/}�� ��{hf��Gm�n=A�]f�������~����4g�Ź�zc�O>��q��h+o�����і�C��6��x����'���G@%oU��� B޸��/�� ��3�_a�G��r�!�`���&A]��<0%~]�� �|S�[���h$���H ���	H�~m�3:t��d8��� �-�S�:/��J����	������ō��w�������z��j�q.�˳�MRE<\xA ��U|�a'�iݪɯzρ��x��f�`A$�oDM<Ν�:�2KH ��lpXwu�h�^.�E�i�lk�*C-Ȇ��M�[*�������v,�ܗ���NǦW���G���t�dgk��T0@7k��@�WC���EgfD���=P�q!���	0�FHay��Aޫވ!�j��푗Q�ҥw�d]gM5�1�� �v�
/�����Lts=�E
^I��긌Aj�	�e�4�\�>_��6����~�Po4q.�F��Gb��r�����A6eE'�[=�K�H�|||A�*���Pf$�����7tH����X�1ܐ�U���ͤ�+b�?v�x��]���TT�����Dw��\�xEt�1�t�Ι0�cR�	��2�܀ ����^޻��UD���kr"<���.O����Sӻd�Ԙ��؛dl`�K�t1	bF�Ks�%Lr�6&�:�$ �E'����fv��n�Im��>$��sd3�"Ckf����$P�ix6
�{�fdח�c#I�3�g���Us鎾��{�%O?���ȏH�Aj�^��%��Ł ����n.Y�����8�eg:fbY�d��:,J>${����!�'8�g-����ߢ@=ⅻ�G������+<�$�r� �n�/GW�8����Iv����i�iEoS�۞G�:��Hk1�����_mi�����}�Ka�cZ�Q=㫝��=��W�l�p��V�A���e�]�=��b�V`�o��� ����󇝈>!޵s��0wpJ%gLA���u���C�v��CU�A�s�����z44KK[5Ҳ���W�(V3O^c],��$M3C%�l�.�����+c�%���N�WbA�L���5uDx�(k� �^"���y��s�մ���&:�
��[Ưn �mJ�if.�ً���Ӑ#�8�.�8�ވ��K�b#ƴ3O�w;�>$�O�\^�cV�M��h}�����]�p�KP�vg`$���\�� �Cڱ���B)�pH5�W"A#v��tV�f,�A潯���F��'̋T�z#�"	3�� ��GDޣ��t�-�W�M�q�n����r��Qy��׃���C���س6/��,Z�oH��3ʕ*4�����R�3ɟU=�L�537\vP��O��K����7���ǔ�nn�7Ak3��E^5����H�&�C�� G�~YNaފB����w�{z�g �0\0�,�X�O��r�L�G�a�K�N9��˚��L�db����b�*����!+�Mv^
GE�Ʀ��a��U.�ab)#�`c���]q(�GkR���#��4�.4J�H���#rl�u��=����:����c-���l�7X�&c�F,�Mb�J+Jඬ��5��0\4�!��Yf�]m[�Q��& f�������R���w6#�g�y �y�-��FWW����[�\B�Z�{T��0�	5,d��v�������HC~+2^	����$�:��>���B��.ю�� �W<��i!��ftɅW���A���>�p�yL?�.n��Q ��� ���[�,�[�v��ވ�ة�^�Kw�5YnL��2`�U@B/n`_���z�A܀I����5�πA�����灞���t3�)ù-zx��[��$�e����A�$����wuU,�Fc"۷����+d��L���,��y�<c�Wu�B�9[�<ձp��H2׏^�M�ْ$�w���m����|+o�籮�3L(#��"qb����]Z��$�����:�u�~y���|������'�O�$I�&�u��|OV�@)T��qjEb���/r���1��MWص�b;�!¾�x�$�k\c���&�v*�k�����E�#��|7�ik�������oyv��]O��;Z�_{���W�����������*�3���x� ���q t��5^L�I�;�Q����e�QP�1�9�6\���tY�$�dޘ�@�$[�&�	7Kr̸}iך����O��c��m@�c���d嘰t�� �]U0KY����C�fS��	o� �Ȍ/v/��������	j��l�r�8w%�O�D�����6T0�
�����!���\%��	��|j�v�$Iu���7�[sx��&\:�R�L��˅�bV�-è:�Es�������`Y��z�r/��C�j�q �����
d���K��j�	���u�A��	Gx��0v`��͘GK���!��I~���:��<|I<��|�]sq�L���󲽏7��z�c��0vpB?`�I�ِ�A��wx�q@��i�kL��T�M5s�����?r�d���'ޞ�yz�ӎ��͝��c�By7U���
�+x�Y����f�U[���ǁ��Y��O<�Y�ڽu�#W� �txo0��Ǭ��ΣhT��z|�і�+/�t�פ����>E�*����>�O+g����~��yvylΪ���WGy��ZѼNw�'�gCb�Ty��n�v���'�]��g�+<]�~�=��3=���P��5��2�	ͷ\gq��f���xGN�s�3�'��,������K;K�	��]�{�d�W����֭i���s���_���A�&{���	��;�I�/�\B�y���j��KPsQ����1)Y5/���5�|��k��WOy籀R�W�
o�_{�vK��8Q��Ӄ>��2���D=���%���y�7��V{��fŒ�����[@��7À3���Q��hB�&�������^�od�l��~��B�ܲܐz��mz����V@���݇Ĕ)��-�V��|��N���}l��f�a�����멳�j˞�W�qF|�&����m��Fi;�~6��/vz�ޞ��b�n^�N�z���l��r�����m1�Ə�I���ˇد�|�=����vX�,@=���(v���u�纡1�|}X�>Ӏb�e�Y�<�pc5Q��E���q����'<Y��r�f�,��� ��!E��@��)�R�E���ĔB���!5Q��G&�%�ž�ԉ�7o�ѯt�^��aHN\���&w�%@7,rp�j�A79�ÉJ㋣��:_z)'�~��|��}��C�x��۷oooO�nd�a$`BD��N$B$E�;?���Q��#$<|q����鯎ݻv������̇p,I$���	B2�B1IN�ƨ�[@��ɳó����6lٳ���ó��!9%	B�r���tDIϋ��������xlٳf��Ώ�8��"n��[e~�l��N۰����ܜD��r���{����DK��R�mk2�;����.��ZpW�vV���mh�8o�^�E�[MTf|;;�B��<��?��<ͱ�k1�H������<˃,���GaY[j(�I.)�c7@i�m���	(㈁N�߼��I+�����λ��'��Ď�b��n�Γ1�w1X淚�
�A�ُx �e?[A$���|K��2����8d�S]0 ��9�A�$0A�U��]8��z�$ .�9�6vȳ^��̷os�B�@��Ə>����O\s�:

�D0Y�D��Q�-ְ8y��@��C7EP�&��6��Z�M=~W��gr�{+�XH�ւI]�m��#���N|`Ɋ��Υa����Jt�'I�=ؑq=2	�L>�i�B���h���2��P�-�'holƺءF�<�vb���@i�����x��U�O#;sI'�̻<O��ވ/�6ܣ�	� �
����׵���"`�t7���@o+ַ�	�m���m��/M
�4
�R�KCM0��r�r`���fc��6�p�nۿ�w����AO}K�?
J�{Gv���j��ӓj$+6�"��@_����|A�2�($怒WĿ�I7ΊgI�նܼ|�G뺇���Ж��*yh$�k '{m�E�nm�h��<D���~�\Rmu�kAP�P�(�@p3V;��n�e�<�A#�Pwx�b��t�M���䓷��A$om<]�(�c�<���(�sp$��� �a4���w.�@pz�y3o5������� �O��	� �mG�p�psy�	�
���
r��獈��x�LA�$gn@�P���m��~H�v�Ć� �catC�XE6i��� ���ݔ�0ݻUy�y]o
ʷ�B0-�ݸ��ARn�]}7��+��������ħtJw�ەI>k3�^t�6p�e%�G>h79o�5{Q���)�
`ukN���%�Y��f�W�<ӫ�B�M7��w�yh���1�]�6{�xv�?����.��״VT���<|KP��G�w޽z�,��'�G�*8E�EA�mu[s�; �-6���+��f�.�L-6j3������7+�a�36%�t@d��\k+�3]%6SQ)�`������uɵ�wR��3Je�I�h�Sl��J+����#���K\Gh�����N<����Jj7�Mb
�k5i�"´++�!,��h�ir��e�V0&ߞy���	Q��	��2]�6�aaYZ��gV\��(,������\���˾�1�$�v�A�}���g�w�_b@κ���sz�zX���Ȃ��������{Az�z+]������֗�t Q��	 ˸Vwl�tC�z���)^��&�ټ��Rj3�&�D|w�l��c��禞<�3�q �{��� �!nS�������b:"���>�@����H$^;�A]Пi��I;�˧���^��hN1;1wwe�쮦�D���~� �E1a;�^CU��<պ&@ ��|1~Kƛy�_uo��|�7�>�<�Ɉ���1�I�x� ��T���	t%�hs�m�J0�����|���+�%	�rl��0My��+bI��Lf�5��aN�ǶB'z��0A�i��ΊgL̰fzA���Ǒ���=��ǣ����D-i��sw�zl��+���E�d�R%���>�]��ma�za'.��{k�p�&o:��!��t��ח�6$� ��� {~!y��`D���"Q��41������{"@"T��rN���)��0jO/� ���K�q�Ē�kb��l}S��:��W��CD��۾��#D^�-��"���U�j�W���������֝C��rD'<�9k`y�}��/D�̸��-�h堖�y�Fz'����E��{^� �7������C�[�k�	�ym�>-����^�ۈ�������������KML�+Ut�ҹ�Wi�����]��'��M��1���|��c������)��A���^�A$�l���*z�Ĵ΍�ݜ���^]�!����%;�P�+� A6�^s��I��s�/�bۙ�\$A޸��M:!ݧ<��v�&A}�M�S8I�ٙ�U�ND O����y�R�żZ��D
�ބ[�<�m�s�,�݇^���-A��3�ƪ�-�'7��D�K�0OF���:����.����x}}����� �.sm��J��IﲠF���Ȃ��������\����;\TT؉�$�聾H��3ܴ��Ñ�x�Y;S�ݡ��:�;�����Yit&p��o�CN��$p�Dy/]�m�)g$�dy�=1q ���;�8k٘��^�e�AS~�lF���B���g��m�U5C:�FQr�P��ݬ �#�#���v���]����@�y�Q$_���$�elsE�E��F8ڮ��}7����"q�NY���)q>\y�J��n�t�����v#���w�p%mx;���A�o]ѓm�9@����y�N��AJ����d��y� ���;D6D�*���	 w:�/�imsA4㙼�O	M�������T4���������#�VϜ. ��~��
��u���1i�r������Ҟ�{K<�|���?����n��&815Rp�h_e�5�-`hƼ4��'���v�N7���HIX��d�Fq���<�h�x��(?�4�c��䓕����8�9މ>荈�>$Q]� 	U��M��߽�~��1Cs�@E�����@���ńVMcyt(hM��[Y��U�O=|����_�;3� ���л!����@>��k$]b�M�Ol@�C�-��Ā�x��I�Ab�C_� �c�҆]�[��P��|�� ���ao���*ݘ��R��n�L	�H:f.��t&�7�Y��	$�"�Vys�	`�<Uj�d%����#q�!��vA-�s~���>�l=�H6��"k2 �7��eo9ũv��Zc���g;�&c'�^}�G�ё�ҹV�V`y�þ/�d.ߡ�޻��5c��;���[�9���m>���=��޺�yV�3Y���J�=/{�=���gN����!�y���[�b�/�Ke@
�+집�g�-�4aD�3I���>> x��>P*�%��p���rb%�hҰ�f�B8+�M���ҸXƎ�#t�b��C9⅓�a�SG]Kx���@fK��y4��
����hX[���D��eVᎣ��Y���	��K����7kv��1ݰ�7-�u�+،{V�M�m�-(
Q&]��-#k,@ή��2�X�Z턱sP��[`V��!4�� _7���a��t[��-�m�B#��w	S9�'\�T5�Gy)��~��`�A������	/��S}�� ��툀�w�Ŗ'�����xu�L�^�`��ýĸ6��F��zuH�u���Us�Б5�޾~��k��^�@�NTl=3y������Ho4pUd����b�G_f �I��$�s:)����!u-�=b� [s�� ,y.W �q���3��@��>[��ޡ���8@� ?���x�|J�ڙ��9���I�>6UL�RL���.�:U�M}2�(n�1�""�7}p�`GVL�'w�ͭ]Ո($�Ֆz�r�jh[sG���]ق���3U��r�Hk%��j�<jߟ�]�b�]v��a����#o.D�p��2 ϛu�a�;������N�� �6� ��VCkJ�U�?�9���mo��������$*f����N�)�8fe.���Xf@PKA�7���
f�%D�dɫk��Qt���)�_<U�@Am]��	x�U���X�u��@$�
�r��)���R`�Jt��!Xf��r��W�!o��۲LgNk�r�"� O�z����J^p�y���+&�TF��C�D�L@$��G���ȸ熺v�F�Xb�� ��m�L������q �Ufs��X!x�;S�Z=.��r��A$���k�����.%6+���vwf	�uˑMB`ѕ�.�ƷZaΣ�n�4�E��l��i����d\���������)�I}��*W/K�[���M�D�EB��S8)�:-B��<�9G: �c��}o0Ey"}�� ����O�9.ɳ$WUs��������L���`�z�	'�_Oa
���9H��/H1H��߷�nw5����Q���K�[G��Y׷b�/ޤm�X�A���ߦ+�O=�ɮ4fd��#�J=�}τ���v�A'��3�0��X�\0N�j")��շO��F�������>G�sOr:���� U^8�}�ef�R�9%�������$����4r��yB�BB�:$�yf���	=�� �)�D�?G������3Qf�T����LہX��� �ؼ¬R���_����˨�s�����O�����w�|	��5��-1��vz���3���t:^g����dL6����R�����.|s�<���sbD�!f2�Bێo@�K��-���9���CS�kE3���p�r9�$�>\��$���qՅON�9%ݱ �T�AQ��wo�鈗f�v�RYzǯ���|k'�<H����a��ዕ��`��*k�����3/��2����q�ϒ�B�`^h��x�d�L�;�����f�i��hM�O��k�~��?ľ!�A/�Ց �>��X�\0OP"F��z�$�ܧ�zkye�?�	l�	�����M��A#{���(�g{���8|>$/��Ol�E��X3,�^"kK�:�$]-hcj�8�b���=O����D�%��|��I7ӱ�$���=�U���C^!0�����A��x��;9wv)�֋�����æ�z�pM�s�o�q&c-����$! �zӥ<p��Ѭ�v�K��pZ�������\+de�UEBS�(I�ΏA'Čޘ�'�\�
g��p��e���r�g	--DK��{�Gz<��y�.h�@�ރ�-����^b+�*.���⋄]4I�1�O���=!n���zi4����*�\A<BW��7������g~i@����fڽ=2�X����c�^����精|oL���3��a��*�?���[U|�������:#�[�����I�����޶R�U�<��!���;=�ѫ-?wzn�S����ZYR�N��w�J)ݼ_d����bܞ����S$nM�se�S^�ǳ<}{���ͻظ��\X����s�~*�re�ظj,]Z�~���x[�v��<�([˙�p��bΜ��
~=�Gyz�c��R	��#}�z od돋���<����|�e�/k[={ǈ�&(
Nǥ���yyٞg��{�9�ɬ,G DS�Jg$�U�XҰO�a���!��͏��×�M�;�{�����'yzH����}�{h:��f�{tj�Ob�CÖ�@�5�sEb������=�Ov�=�o���/Lg�w�/�nz-�}�8{�d��f����z�G���f�Ή�y�*v�u���rk;�F�}�
�ӻ����c��M+,����^	ټ���|��x�W<;ͨ�x,�5v���34�h�Y���ո��5�t�u�j\�����_8{o�G�>%d<�>O�Y��(�2_;�=���~Y��	�����l6���m��{��ULz���^]��ˬ�j[��[�wX���^B^�$�G��b7}�h����Aj���w/s2
�<v�ry�A��}}z5r�(@�}q󮹬�/{�7^hg�_�+��܃85�М�|X�o>�7"/�h��g�5�Q� G ���2.^ǀN�`-�F�i`�X�� 8��|�$�!�00>������`�jq��nOճ{��<�?�<��saֲƟ���7�CE����ʈɿ<x�ӈ�xX�r5��L���w��jox�^a��d��H�6M�30��wǵm���HN	82�e�nY�% �Q{xv������ݻv����v�d㜣���mi�wk9�w��C��;�вm���"�חޞ��x��v����麑���\	�aV�d|],��m-��Nm����8�>�����(`�bō4`���(5�%����E���gY|��\���A��g-�R(��I�GF
0h�BƆ0`����/������6ѝ���V6�e~;���8��6�˲ͷr�wʳ��[6��}oJ��{yY��i�ݛ���;.Ҷ����ue��{u���*+lڕ�\eY[7dm���O[3 ʳ���Փm��Y�o��'�km:���V���8��+�����,��fOk�ϖw�kM,�_~�q�qy��5�Z[wM����+m�Ś�>���v�[nB�m���8.������:�I@
C��T�����e�4p�7b��ٴ��Ŷ�/A��GHA�:��R݁R�\cAZG(�Du���Q�%�v��f��0[Z�������	�M�B���Ůn��\�P�?�/���k�-��
�\�L6b3bWL�V�e�k4�1�^,�Z@���H�k�b�2�[�#���6b>lOSBA�:
,ts3q��f�(m�vH��fSKI�lF���[�c3�f�٩�2���V�(C)+nH.!+�땹�#SQLӛ�ɻ]�"��]���j�	�&��bBm�����؉�7��bm�!�㣠cT�R�"��暊ۋ�1���5e+.��sa��Z��hf,5	E����h8�	�Ś9y�J뵬B� p%��1�6��Xh�)�m��n[
�b��
��h۷5�Ci�u�V�0�-
+LGD��*���R03Z6d�6Zf��Aj�Mu�-�*,\[\T�D!&���r��P[v[�rM�X,��]#5����.���0��T�M+�,��+�#��9�]e���G`m�0��{0M���r��m�I��hAVC0ٴҵ��H�b4��GL0��U�P�\f��[�bAj�jʸ�7\�T���W\��1v��%�Y�˚�:X:.�:�Q�l�/Lq��ڢ���٠������u+b�(KB��[4VS�������S��Ԃ��H���ݖT-��(Z�;�q�B�q@�-�+��O)�)l#,jV2틈�C\����aSb�4mE���ħ[��V��36/��M����K]�����t[)�҅jgV�F9�2�yɴ�b�9XSa[���ûB�8vmNh\%��$KF[�����[:�]���Ep1��	��L��斖K�uv�0���M�@Z�ܓV2뛵GkCMh*��+1�4��]���^�B���瞛.6��c�ŷj�f(�[2�����n�.�]k
��a��ܮBZk
1��Z�奖�L����^{F!�i����Y�iLE� 4*��S6ۣ�[�n��߆�nv��p9�j!5�6+����\n�٦�2��`K2hG��p1�	�m\$̤�h�:$ggP]f!�E�Й��vp&�R�u1[���Ję[3-f1�X0"K������[i
�������<@xw�{R����7���<y*�2��7��tǣ��ͨ�ȉ;���D�w��GT8�-a��ЖNFf�H�C����A ��uwG��}���Z�K��
�A�W�ٝ�:)����P$=����dy�a��%�ǲ�(�5t��>^G�: ���m:^w,���6�3�{�gb���e[�y�պ�x$|TW[e��	�q� �h,υ'������s?��ͽ�NȻ�cˠ{�܃����x$���YOYC8L����������$���I$��	b���b�L�P5fW��B^�Z�J��S��({��w����Swx�w< H$�ǀ`ǋkWDl�5T9���i�66��+{b8�I]n�lȮ&&���ɋ��%s�x����q���������Ḙ�e�7��Z���q��^p�G_e���Vo����}s����Uv���w�|||A�[��a�	�{��A$���� �}}��
�bDlo����'l�Y�v%�����3�%�=���mqk9MY�	��ȀI'��(dN'fwvr����{��D�-m�n<��vO�GS�$&����(wcɫ�zER�:�b!�bt��X'	�J}�Ey
�i���mNC�S���㱙��7���AlF�\:�Dgz�)�_�5�s�M�lr��#kM��e3���b܃�Ƙk��}|�֎�t4~�?=|���0E5�G���3���w<��=���I>��w�[�M�vY�'I��h���"��#��_U��I����3x���#�.���cv�����|��LZ�x���"l��@���x���d�WCK��M���c3�P�xS�Y
�çp��$������.9�ۓ��}�.^�G-1�bG�/��v=��������>>> ��#Lt0�W��n��>�Lx�@��K0��v%��s�ąqc�:��^*7�A �|}9o&�"Ogt;q��� Q�P�T�B.'S�m�H��<���Q����>��\I�ݶ��p�j H�ף�6H.#���H6�YYu"��Y���v4ZG��ٵ�;�`���%aA��heJ���3�����}��/8NK��T?	�h0	�=]�O�����(��Fb�
>K6C�$n�р*�%�L�fL�ٜ'2�@�I��ԓ��������UO��O[тo�}��I�U�&fQY^���{��������<�9]� ��<�T?�ZZ#���O���z0	ymo<����6������:b��V�]\)��x�E��H������PЭ�\�l�s	��&s�=���HCn��S�m(VC�Be���dQ���ޚYnb�m��'/U��YqqbJ�#�@ �
��;�F���r�8t�g^� NgS��������3=1�+܌���<��W���gz��'6�6M�q�H~���h�m�X��(V�-�R�QI�,���y<o�b��ާ����j���_���~o^R���y��+�Ge	�	����Q�����c����;v@�ځ���\8M3��	���Qʩ��k:�L{��ޫ.i��:�=]n���1�n\�k33�fp�6���؃�똂>=�[QqÙ�L�|�!VtG�Ot��V	$=�/k���t�}���-�DwK�d�&~q'֒���o��|77v���o-�,�����v�����ٶ��Nc����
`�i����Ƨ� �H9q� ��{"��i�lF��[����i�@0�%8�Ӝ :�q���\T�4�VN?t�|�1�=�&v��w�c~�vm��~O�q���0���u�Q4���w�8�!/�^~q��XD�ͥ�b;k��[�GhuI�)�6��%V�;�I��
Ɓ{@�4���u�з�Xİ
W1�#[Qi�P(Y���b6-���8fmFZJ�`n�ƖjB�.e�'`�6��Jk7i��������Z��ka���;6��,,&mA&�a�l���
�.ɉR�RT:�BR�g ��(�a���um��K&-IԮ�(��Ibj�n,3i��~�>���ck��|�� b<�1�DH$ws�yI�8j튉�[�̹�U��A �U=s>o.9�gwE:d�����<��ˡ��{��H=��y7y|{��lU*z��1�#��$8N&�<ѝ_�z�>D2VrP��g�1�t��G�r= �;��m5���˳8N��&��b��J#CƟp�3f����@7x�`}����f�e��aj��U��m�&#����ıvh�~D�r�'Q����l=F� ��؀I>��Bw� Mc�\ҭ�5�<�e�ߪ��l��Ѯ�kflΡ�֭��(T9I�lef�bU�̷�ߟ���ϕs��5�  ǒ���	oz��ki�F n�w��ݏ���3�]�ד&p�=P�ځ�(��b��ID�z���[���� ��>����)~�p^g��2�$M�7�p�tM�N�jq^3<`6p�!�r�]�{}	�I?�L`|�� ����|$q�7�]�d$���<@!zq�g�n��8)�S���d��-�D��fs�$c��͓��l'r�{`:
�{"	��$@����.Rw%����;�!��=��}m�*��&/�;6f$�5=�m�ؗ�<�Bk[Ǹ#ú�)K�^G633�vg	�`�f�� �=7��H�j�-Q��?����>'�]�~1�&���w<��N���<�S�ع�\V넖�P� �����-��m,3�]z�)�B$��Mв3���.ͽ��Ѓy,�ǀH��> cuXX�w�fA$���'þ�?x{KN���P�Y Z������`�DsnFzV�y��̉��G����>ُ!��.��3�I���	nN����37����uWr�3|���\���xO-pX��_C�󉫀�L�m�����`��=pyT���U���7�� ��6$�H�t@� I����hs�')��ɓ̂��7=[�R��(O�ӯ$�@>˛�$��{��M^�ֲ�6�^I��[�G��}��g%��yO�&	���N8Bpv;�D�I9������cŵ���ܿ���}޾KY[�AXʩ��Ms.쮉���jڋba�œ�<6�Y����ӄổODx�(�MǠ�I��`��S��5`)���$��<��K���-g�.]�d�l3�
}�.�g�*2)�����T�;U�{�H��H:#�z&Ŭ�ft��0�K�o��Kҿ����o��^����ر�	���IK����H-��[��q�Y5������������&v`��� w���[�B/m����������l{$��G��usقv"��%�N���<
����f*(sL�3�GwDA�+��Д@:��9|f�k�=k�*�r���n���˲�;���7���]T��6A���R�R���,��Dj}�۾��|[oNuϜ0IHF@I$ܮ���"�]VTw_[u���Gƴ�m)iJ�I�\o�Χ�nf2)���/���}9>���F�S	�E\����'��� ^7��GW������U��i@|���L��A-�35�b�))�:��YX�0ɷ3e�BC�ߟ%�ˣ��
Oh?A�Ƹ�0M���9���nqӈ�EU���7�v,�"CU˙�;�p�6����^��ɫ����|w=�e�H�&˥�pNR�����S����)ل�L�h��yu�< {�Y���F=�m�L�ǈ#��{>��w����3)�҆t�3ă7���FW�*y� �2BXݮ �J�7E�u���.^"�-���%�0M�.BvgY�6�)y�INtd���+Z�K粌��f,ؿ"��"c� �ˎ�Ѧ�8Ou�#�Y3�r�ĥ䑽#ɓnC>:��&u�wo���r]�4��œ�L��Y3�~Mo2;Na�qXGs�%�i��ϖ��g7��|s:���L�z�1�)ZR��׮�Ռ"a��٥��cD(�FcX�.m��i�EssXA�'V8��ka�5�ژ5V���)v�,����@]0LA��0bZ��bk�62���Q�31�ji���\��eX�	��X�V��ւ�eM7Y�K�
�QڐA+Y�����v]��a�A��g=��q�`�����\E�5f:�S�5�;CiX�\;�Vʲ���\�6n�m*��;ZY��L���{ǝ'w,3'���L5B� ���x�	(�E��=�-ɂ{�g��旃�m�=�!�.ɐg�2r�+�o]����������Kw�  ��o?������U`]9�A��3�wwE8h�i]O�2�m���@��ˑ==p`����p���A��<�Z��ĺN�@���DS27Ȟ�׀H��~��$7����^�0�^���l��=���l�	E9q������#��q��"�L�m�	R��uT��p�C�ǻ���+���RE�qr	�f�$ԪքLɥ��e�\a	���k��1B�݅�X��]���}�3f�	���	�� ߚ:k��{�]q �=�A�ىdJ��'S�vLf/�q���7Z����U���g��{w5Y�.:N?z{�yW$"��c�f���v��No/=�	#�����_���_�L���W����Q��'�}�>> ���u����4�C�����Н�����eݫ`MvuCU@V�:f!�˴�%� ��@���G��� k�q���;dfGD7�ћ�^~'o�u;wtS��8�q�j�yA��O�>�{<I$f��I���4l4���$�T���O2v!�t���[��8��^A���4��m��~�y"�Zȑ+�_v��UZ0gu?���K� ez*j8n���,�YKc$n�sj鄁5����,I���ì��P�3&��c:�B��ky��HM��!�y�k9���,�_|3~��	��)|O��JM7��t�G�Xؖk%E�ĳszD0^D��Y�|Nm�@$ɾw��<�2�" ���*�vt�f/��k\��灁-��z)�#��K!�䋐�=��2ɧ�/0o���̛�l�/�Q~�f�HPq�t����"���'�w�y��?|�H�	�x��яM��`F�w}S9�{i��G��ˣ������xr����Xs��3���U9����O�{�����y8��b5������ȆtO8��'�}rﲖ�5�~�E�ާ&ۋi˞��j�C,�ϴ�罉��3ώ
D�#@��e�|�Ӹ�Da�,,c'���4��Lю�����G���׵E��(;S��8�M�}�16��g���׾���>�r�Yf;�۾�v;H�n-@�.jӬ�ْ)��d�u�.�7�����Ew�x]�7�e��u��D��e�M�B�ɿy_M� ]�������<0�I���D��z?g���!�}��	|p[�R�6�a�2q��|��7�؟�	�_*��3��<���7F�����M���y9�c�Iޯ��z�	�ٷ�=�1���`6���e�����iV��B��wA���^�Y�sT��9r�zx�w�-i�:�o]�)=�q�׹���֝n�3��=���^���ҙc�N�a�[�7�}�*]�˞3��A`;�w���/x��X>��d����L�%�8=ꂞ��!�vf��jߟ�MN�3�^���yfD�d��'g�úiH?�b��s):�}"d7��^]��eY����0�Id��O��VtE�A)"������33Js��K�2'R@H��I �J"̆?!��A������_nm�[�W���lr�����>�n�_[^Av��J[!i#{�԰,,6�����۷�o���v����ɪ7]I�W�Qw$V�࢙��n-�:�ۮ�S,�|{����������۷�G��۷ooom7����݅�[Te��6�+f�Cs::�}����H�FYI$HZ���6xvvl���f͝����d�>;���3��ݜ�+|�jY�@��,
[{8<6l����48у,S2H�|��+6�w[n�;mGv��vVVeG%�M�2�ѭՙY���U�l�촲99;;����e�ӎ��GOn/�]���훭�ci5�!pGSf��F�;q���o�^���u��e���vۭ�u�w�Vu���Y	VA�-�|.�JC����GaYv���^g���v�����;�E�m����k~>^qY���ſ5�;��u��³����"���;�μ�(R���]�w��A�R����]��ސ�!��"t�ސ��t�C;�j��ndb�*���l0H6��	3����vf�����%��ڈ���w�;���5��O]A�3�p#D���@��w�O�;">'�v9�r�c����H�I�x���h�bf��!-�ݠ��[bh�W�V!c�2Y���&(����`�C"�;pa������2$o����(��5�[��o���,��?@������kJ!���[*=�M>�॑��3�y�|�WoD�L�t@&���e��c��-b&gfr�z&,H2:.B����˳K�+� p�@7�� ���;:v	3�=�ՙ��
��M۴D����G@�{���������N7^%h�5I����=�?x��ȝ���^8~��pD4�`��8�m�v��SJ|,7u�X>5Ik�3�U�H�Y�����/AŽ����zH��C�Lgr�u�7�$�s\-�z*�
<��輈3��AƎ`���x0P/,f��m�(,����L�	Di\U��&K55�Z�۝-�"�Z���_����>�v��Vo����$����4$
�k0��1�kO^��v��E���ӕ�Y�w �t��A�^U�����c%�?���I$��Gۼ�DxN�HL�0J�zsF2,�TC&-~1�Q�;��(���.��#{�0^S��#�n�ـ4$�oR�!�fvg.�*�����b���F0��P �@;q��;8���ފ�՚��.v������q'gN�&b�7]�����EHT�Լ,O�.�O�tTA�Wn>�gD��$i�۪&E��,��>y�MQd��S�@��C���[�_�.�������cx�O�ɉ��uޣ�������>$��Z�g�>����F�����׬��^zg8uJa�]A��`�f4H�{�y��_4�����P��KXc<h<l�ؘ����F]��f.�K��� �+�]1����9�:�X4a��ٝK���q+��b�b���:5wYM���̑�#�ۢK-�`%h��C+�alf��V���C#�k�Uds�Th�h�%ݒ�t�����,Z�ti�vK�a��X��A��kRY,	� ��-��̆��#�~�����Q�&�L�}A�� ��k�AC�:��Y�֩��8R�O�������ē���ݝ᪼��$�v"*�ٌE	��sq+����|O�s�^��몠hZ��� FOaf!�Ń�����l�A�ǒ	�cY��9�H�n���fԖ�;�aZL�TC3��S�|�nq�:�f��#�0H_��z�xI�~�#���<�x��Ag(�$p�g���IXb]2vg.�&���- I͞��Q�rl������LA7ְ��=O��*Cvl%C\�>)蒓�rL�tJ;0�]��4n���2��`�K��G�6�\*��������;������ �j�^	9�îz(XMp��!��6���O��́��sœ:,L��P+f����3�Q�����u~S���G��|sz��F,��H���?<7��#�C?v�P���yK���-��őiΧ��L'����x� �;P��^f!�r ��y*���kܾ1P��8����g���ӱN�	��	���6�I������A�^Ac���=s �7����,'k��<� ��������O�����������$��@�EW=��#�ގO4�\pO�ڸ1�Ѳ����f�T�FzQ���
��7�/����bk��! H���"|Go=���öb�r��cP���E��`�h��� ���CE��ֳl �h!A��8w.�hb]2vg.�����	���@�o5��W��Q��)��1] ���= U��mI�ݘ�>a톨D���
�׆Y�I� ���^�j�]�f+�����k�� �qœb�N��z�Q�,H���� �^Zؽi^�v]�%Th��NP���^bɋ�(4����,F3�t犑�gg���;U�7#!�Φ���\���Q]8��.c�!�����d�~w�a�!��"����8�p�˱v-f���b��LЋë�Os� �MV=�/z-��Os�y{8��j��%y���'���'�o��k�DHV$�D0^��d���!O���n��H>smnﵚ,Q�"�Ys�]�ő͂ގ1kA\���2�܁�i���Djd�C�Qbx�=G�J��k�|l ����<�qycE�^�zdNy:& ��G؀e������Q!�u��9�o($�{2 �7�K�kŨn�[�я7q+��vwf&(��lk3� $��lT0y���O��q�L��yG��^]��|׽�z1E�L�p�w.�3�z}�*zCTe`F��aM����|��6
�yG�WRvS�5�T6�g�|Bu�*��m�`r�|��t�~�d.o����)�u���p}{�r�/�vU��-t��;��sU���C�͋�@�>ޟA��2NS^��.h�໇bᚩ5t�>=Qp!>�����ã`����@$���!v�s1��<[�,����V�4x K�.� )e����`hY��{j�KJ��Ͽ�ϲ�1�?9���1ncǌ��h�7
5��أB
����|�����p�$p[Yr �{fZ�n�:��em�s7^	�;�Oq�:�t��v�W�*�1L���;3�{^'����H�}���J:�Y��U��$H�.d�<B�ʱٙӰE0y���Q2�Wd��I ��<x�O��62 y�ة6X����$(6d�bƀe�n{&i����+��T��͕V"{��>$�ǲ'ۼ�BEơ�e��_��A�V{��=��yF����3-�N��3vL�h�(Rw�w�z^��j6r^��
|��ww�����nL�+�m�a�$� �T����-�suSY��||{�/ޞ��8���盜9��Y�f�G�*K�R0UԦ��c:�i�Ɩ`��Q��3�KV��&;SK��6`��k]��к��D��v��*�k*uxY�֣\e{,��RMs[���K��6[�e��CW-��v�̣5MZ5i�&G B�%���K+T���q,�PNnE�YY�k�հѸR�k�U#)��T��J,`+�r�]����nF�J���R�N:s���pYñpͼ����O�8��f�I�@��Lc��4/Q~{�$r�����6r��<�薸��=�+)B�۽< �E��{y��R�9���.���S������p�7�+)�ZF��NoNt:i��5����F�>�� XK��M�592v`��*���ֽ	�qs�CY�=> ��ȳ$�Gv�Klk'����%�m�H�\��]�1LF��_���n�<pV�6Qލ羰O��b<O�W5�$����=S�ߟ����߲��fRʍ�2�3:k)�n�F8�����kZ4M�{AM?>T�3n1��e�}|�"���E���y5}`��"Ѿ����`L�=�A/;O0C\r�\3L�Έ!���g����ȪY7M���(��xz�r��k�6��R$���뾝{�r�M^�/��؇�cg�g������|A@�k�	�ֽ�+���`����i�´v����$���9p�b��t5� �K;1��U6�v�׷=��Dx���$���"� ]L;�b���:��lڨN�׋ݠ��=6<��g��\?�șާt�l�1F B<�`��0t�ك4�Eh�$����}�6�W�9��0ecـH'�ױ��ޘ�=�=m>|��FU���m���I��@�<��[���b�#)ê⩧�����M�'��.�l�� �v<B�=Ւ,z"�G�>]�s�$X��|'͕hBbX�^�2�4�X�����!���ȏO�wTz���'�"���3|Xr]˹p͇[��>'��]@���[���ŰB[���ꪜ����˹����~���y�a�7��[�ǯ�[�{G�ܣ���}�ٳ�sǻܸH�w����� �/u�'�� &{���H�o	�H9`�b���-��N�����f��o8M�,�����;��P�t�v$Tb!T�@$KE-��b92��h�j�L��$�j�#�WUO]���"c/����x����p�7tHy.�x0FԻI�~~G���Ǒ��m��̲гe�!5J% ���J���&�dʹ4�ѹ�}�~kE�ߺ�* �	�	��7���W[0�t@�+n�D=aU���݃2d�&�z9�5���˫}��]Q�w�"|������ak�̂�%;���+���	��l�	�N]9N� �� �}mP�/-P�o?s�x��y; �vS�'����ZXr]ˇp�%c�%��C�u�$��?G��	+���F�tv2�A瀹@+�Z�s���݌��*���߭�����=铔�0�7�{��-@ɾ#Ȳ>9ۑp�EK��������x�݇k��A�X;�' 1��V���Ad8;��*O4k����F	����f�
���}��߄�3<��_�Q��� �45�	i�b]^b:@�JbK	��'�罉��[�~�}L�DIӹP�}�},P>fMⵀ؝�/lzf�G���q3͎Y�,Θ���uTv��ܵ-Y;{�B��z��&���tG�)	����w`D��dO�4��d���$��G\[�B$��L��D�����g�"��u��z�#ų�C� ��'h�7T?Z{j��,1 �Y/|�G�� C*�T�cВ;z�>�ϘP��ӧ�h��� �=r���\����|�^13/ �H�΋>��Ta�^��i��5��?�?�i0��}bv�=.1�����'���N �=��l`�{����X-�4�u-KcW.�{�v��"�I�J�_`�U�b�M�^.4qY����m��z�ˎ�z�t��tr)��(G�s�A��_��R=��.�����- �x��/�;��(`[�;L�a�J�H+޿i����'L�wv���/	���N���g�.��3RCx�ǧ�Gg_G�μ��zÐ`�X<v�������[�Z�n�|vt���;�/n"\�x�7�@���(�Bx2t�S_�$$��{_��U����i³���⯡�����H���rsL�M��U�i�]��6F3D�g�����e%a|�2B��^�/�O<�e��tu�S{FN���%G{ʢ$ӎ�3J}�K���&��<C�ӊ?��w�+,x ����#{�n	w�¡j��k}f�>�wOo���F��a~A^g �o�L+{�'lᳫ�t<����׬��j��Ů����N^�m٣��ݺ���W���3}���3��3����-���ܞ�ń��
�\�5��9;5y���(0�R�O��򳦟z��{<.���=�=
N�q�
2V�ozsݱ�_��Ts�ژ����O�u��9��鏴���#�>t�o���׊A\���V��ָq�� �|��x^�&[�⋉�,HhA` ՠ�ɜX���M�'H�:4��} �B4|z,�I۱;���~����@�p"
��h'v��D��=z
�f�3�#�8H�a�B�"�X�
Ȣ���[y��k|��x�a���ׯ�~��ql��"�W�mt�<�V[��{���vw�wK�mv���c��vqfG��շ�y��j��������_^�ݾ>8�����ӷI��Y�˲㠲��#�olm�ڎ����d{j���8�8v������۷��	6����2{gggX]	n_^����ZE�=��m��A�sk��H��$"�,Xѣ�48у
w׎��i�l�������8G;.��8wwgq�j2�-��MGP���������ٳ���:::9�e���K�����ۭ�gYE��޽�����KB�8��);lYe�eg%i�ͭ�����u��m���A�%�Ӊf\��ϰ���Z�u���r��s�gq��dܶt���C�rfrIAݶ��>ioM�6�M��ͻ	Y���ѕ�ۭ+2-�A�[�~�>-��r9�:w����f��FZ')�4�����-,vc޽����i�����j�O�n�3j�[���u��m�`A�yٚEk��9�ok�me铇GtE�}�y}OI5�f���4-ʳ8��0943�0�ź�m��qKD�	��.�l��b��%�D-f�m�K����qR	��ZHՖ"36G,�ez��\MK6G�ȃW��e���,�$�������5Tvf�����l��׈ǣ���2 D�L�!�����%b*鄮ź��V�%�:4�uu�5,%�P���Vʣ�e2�fl��֮ƅ:�,�m�,Ѹ"Ux-��6�EioQ3I�k1\�lٔa�`JV�J����٬5�]VڬB)�X`nv�2�^#-���6\ �:�k�fiH��.v`Sj���(����� �j��u�[[��n֤�ֱS	� ��w ��䦚�V��6��5����YFQ�0�[�@׶�L��M���Т7,+-�.�i��5�
�%p��f6ѹSmAچ�5�9β�hIy j�(���7-�L�Ti����e��.�ah��-溎^��Ŕ�45)Xm�.�XhVU��LGW�Pкm�qQ���:�t��([e����sf6�U,	�j�4%K�9����k�2����Q\,&���¼�ٵ���,�Ù�sT�R�V5��,��o[Z�FL�6��ծ����jfͪikX�Q��\�"�J�e��k��0+i�a����Hݬ��ś]p[�u��B�t�l��(�*VۯVXj��)�f�⌛��+a�\\��Sj ������շfbh�@$Zb�Q��;JY�:�%f�`cJ�s�X��نf2�h�1���m�,.R�C[M"�P��k�����$2蚢�q���iI@��͚�)��ˊ�Wg��j�q�iWQ��MG��q)9b����Қ,t��#f��T6Yj0m�-��ԎP��dH�b\��d��ք.VR勝��r�s��m��S�1�J@2]aZ���(�0 3�x����B	�I����a���j�[���T�41�-�ͬ30&0WF���02\���vt���5�%[��4�m�j�������a��q��с�P�H�V[L3��-�aq�ږ��4�Va��0��Kjk�&)�&͈��B��a��Vք3]��,&���4�K��@�,����+`�@�Hj1�.�� .�n��a���c5q3A �iu����me���{�,`��~7�O��u��D�eD���k\L���a��]�	y�ce'$�v�hp�WN@�r�����+�m�hWW0I���	-���@&��;H/Q���kb�gLY݄��y�� ��9���M�nfcԜh�]\�a�����	���V�&�&OZMX#g�s2�KV�k��w�'�1���	�0 N�[�|U^���(GFL��5��`����26ӑ PdE�dF;�5o�VNz;�g���U��7z���=���\�0����([@�x�&l6��G::��VV�chݖ�\�kR�69gvI�3�Y��x͙��>>9{Q���]����%�Jw��u�Q ߗ�2�.��bI�N�A�X8d�`����c�v=8<�Gjtm�TTTɶ=t���`�ޟ��w��I�?S��G ^G����=�ow��ixL~=��s�oQs�SL��C{%����5�S�$hH�
ט�/ �o[D����g��"��`���6Rr]$�0|ɸ$�=�A��&�ZS!�]��<|NDプf0�:ͬ�"�]���s�cf��_Nc4�c���<��O���mv�F�^�Y���fBF��b�\o�̘3�,Y�ٱ��I9�� ��1U�H���qa O�s>�I$��ȏ�~�,�z������mM��.����r���^%�#��6����4&��=�v�ݜ&!wH�OmA �۸r}�^�v��"cHҡ����eyqƶ�H��C��gb��9u`x؀�*�o4\u-�	 �U��	=�μB��M�Y�[{=y��I,`�̃� ?�� $@H_����f�q�����L :)�ܦ��3nي�����RO����{a�x�eS���G�g�e�}�������
[��m]��j�vA����d9�1R�<||Ad7�;:�
�H�y�;�WfD�<��e��H�QP�c����!.���/�������Un�$���v���5s�N&�h'&�W���i6�}�6}�?�H�{L�`ٸ��1t�@$��B�<��1��!��n�� �I ;�c ����5[AL�����M-	��p)(6����Q��E]�ߞ����Y8,ɟ�:_.HJ����5�o �e���V���aRѨ�F�h�7�p��A�b�wt��QƎ� ��cKf
���PYy� ��>4����4]vu1�����PX|�'vfw	˨�j�<gL�Ao%|����%�ҽc�e�]��A7�� N�9�Fp����	�p��_{�2����ܥ�t�o/+~w�jI%1 �ɸ�O���]�W�6"7���J�6p�$v#��y�=������e��Y>��<'[,�����$��b��8*2�'W5A�Es,������Fh����a���íu�<�G��l���ˤ]����fޢ$�����=��
���h����3q� ���C��d;������I-�rN����Ε5�b�ʊ�&�v(6�lK��l(,�ń��绽�\3�����p���*Æs���I=��`ͤa#)퓛8]Ӱ��"of:� ��Ӥ����H"�$S����������kzY��	��D�R�	�͆ �T5��|�P8$s�l��ѥ�d�wt�3	�y�
<�ƾ�@�5��դN�4�9��[O��<W�;��`)����ݙ��gFUy�:co:��R�������kȭ�iq���ێ��<*\���j��g�(�`��d�Kd/wf<ꭱ^ܳ7fGGD@$���f{?�'��%���?�3���$N�n��ռ/���Q��>ޞ�[�
�o�8A�"Yv������2�<pV=u/L��:~Y>V�����,Й$h�]lhJ�;�8��3�5��C[0-M�`֎h���immR������Q��$�]^�5qK�I��ʼ�-�Z�m^Q�c��1�h.����Y��ڃf�)�f�Ut��`��$���C���p��3%s�tQƃK爋�i��5֕˕��lج%e,��X
:�u�jJ6eu4jC]HfF��\V[�faMD�͕t��G*W�t����P�Ė���DN�b�%��t�r�~�|��ڧ.�v�}���i��sc()�y�O�c��{w���Y �oDO�1�ǉ�znO6�A��ިu�D�f���=PI�5\�} ���H/]r�i]3�{*��q����L��̙�Z�.�l� |o;^$$�ΪWn�q��\� ���k�	/*��aP����2;�E�D���m0C�$&E�7�&��#Ȓ	���3�ʜ;K�dL���K��Bp�N���.*���8� $g&�C�W]l�T�л�Zy�ǉ��zgc�CYy���AI"��X�&���F E,��Z[WG���H�1�� ��!�X�ă��`�'�Q"{1�A�[<D�{˕g71T/=q�&  ��؀H�U�兓�@�
Q>i�=��A+h���1����$��$��KLI��������4����N�=��������a�o�^�I�'���0�3L�l#���pý� A��yIͼ�|�$�<�A�3dz���z�~sm��Eû�w���\z'�.zDA������ ��[�y� �c���b�3:�5���s�O����+�:$B@�&�&d�ͅ�vXј4<L��'�����dwt�4~)��@��f�c5r��I��\$���w5,��̌�����w����dX�4�^ ��1l��&uP3��e�1��y���t��t�.��;���ω�¾m� �'��ׄ���wnϓQumP�s�WNHb�NYE�y0p���-��H����lgn��$5_�k�� ��of|��Y���f��*��,,���Z�~�#yPa��pǽw��^��+o,�Q|�_�|wVV���E�V"�*VM�ճ踬~L�����������3!Bd.2N!�U,�E�e�L�I��W���� ��֧�A�ˎqw�ȁ!f2@�r��g���q{�\�oR$����	=��`��y��vt����i�vmk�r2�O�yކ[c�΂L��I�9�|�"I��x;q���7�I��x ��{0I#7:$HN�U;Q�"���6B�06�n:V��T�{2�1����`�	gSم� ��i3ɡ� .���"%��㧅sX��Y!pvw_��]d��i✳���8�O��H`F���xCfo�2Dsy����>}�#ǹޫĂfQ��Ȏz�p����!0tS̗�l�;�%ُ ��y=�v�D�c�{��<�V�}�;�����O��$�.�T)3�I��M�斨D�����!z�?]�LAA,xCp���1t~/ǡ4l�16�v����m��[�Y�Kf�3v�g�ϱ�|4��杰�q9���cB�!��g��/ܳKu�$��p��A�f;�E	l&��t��s��#���� ���I��젦���岄�[%̝زL��%�*K�a��ڲ�a��e/\�Z�l��?>�����I��涨�W��$/!�/��g^ (��و�]�Dx��:X"�9t�3U����!�y�.�ݦ<���ٰL��
�ݳ3P�q�yfA>T'��`��d'��� h��($��y�mj��4� ��#�:�$�9/q���&�vD&�z�k�T����D� ��%��I���{y�Ċ����3ϊ|N ����.��HVz�מ	��!jek�u�����#%� �@����^[�DO��^�o���ߗ	Ė:��9Є�'ʜefI����z�
hP$�2}{s���z�[���M�/����&qm�^���v�Rx�ݝ>lz�lw5�H�v�޸�B�ׯ/��Tqk��n1e&�k�[匬,�X%M�գk3���պ�� �ٕ����G#��s�i�FkSr�����hE��.���5�M-f���#�\��e&LRY�ufk�SCk)T�Y�+����蘆`���	���%�d�\�� FF�m"�,�%��jTc���T�3��(f9���-{6��H�c�v���2j͛G4*�3�aGX��������\�BRmMPZ����~��%�4�{��+"�&�6=O����1�l"�a�H���$I�~�B�����vbS$DIn��|nL��U	E0>�ɗ�I8�[7Bd?��[�dO�%����l�@Ν���˦I�f�t��A�j�A$��
o]2ה�}��-S��%w=�*Di����tI��A���@��sH�� ��C���g!�nKi$�gDVA�.]�,��O~�3���c�pfYN�T���0��s�e�D�ߓ������K��[�⭻
K�A�nil�)(�V-F�'� C3�C"�ْU���X�Xs�56�>t�V5B��͈0ڜF�Ơ�Ɂ ��F	jO`b�t�ô�O[��,��0��S��<��x��]T��B��&���7��♦񝖇ڨ�����& �l���ǲ1��2|���H�l��VGz||||Av�'���^�}����[�����s[
�[�%�0L��Mwj��%
��p|s�A\�Tv�P:���@�vgC��t�XA���$� ��M���-�&�Z�������$��SZ���)�x"D�=�n�ˊr��t\A1�[��D��=�f�z/c(�h1�A Vv��n�ELz�s%D*]	�l�)-����amte��8;f�qYsFm
���,x&������fK]3��K�Kt((�n<A#nz ���u�Z�"&ߌ#sr f+bqt�v���z� %4�m����Cn�>!GnlA��]��TV�mJ�#p1�V��\�t���}�����jU�4Ĵ<�C�gS[1 uS!�i�&m ��*���fM1�6nkZv�&tt�:����f���U��ы�t���&<�QB�E8��<#ٕ���S_���ּ����w�l�y�;�;s�%㎯-��,��i�nt��Ņm����vG'{��ś��[������g��Pޜ��ơs%x�>^}_�^�s��֗+�& �.qS� �!�3AѡN��\�����z��cIg'��g��3���,*�7�>>Θ9�o'�A~Uy���1{����{��..�,�pa�M=��X��T,�j �<p�������_h��5깯�Ͻ�Ge�r�5�.�9���=+}|:���N���}���oN���~��{�{��hч$���X�7��O='(��Ӑ8��\<��߿!Ǩ���߈ԥ3%��q�Wϳrh쪪�w��@����J7I�_d�{�_v��F�����f���X�����O=���NF�����~�텼*��݊�8��wԧ�����.;��[��1��ހ_��9��;�n����|�Яp���;�������T��L�u�.F�/��N
��#}��s�R��Ⴋ.&�*��E����s��#�z�rжr
W�㆑֬�E��#�y6,����ws��d��$��@������ޏ})1x���8[��>����~ۢ8�������;�*�e��ě���|J[�yS[����U��jb�����J��	���.�3spw #2���g��t�K&�$@+����i��8(��'��gv�mn�o�ݽ��|||x|v����h�n���m���m��im��'H�²;�bqȄL�0�HH<=>=�>=��|||x|v�����*R%�R[m���2!ϛZq��@�3�m$�I�6�Y�;䏙"E�4(H�CF�0hѢ�����>�P#�pY�-�V֎Y���n��.5���J�:G�Z�7_��0X�B�4@т�
A$�A%^�"�l)��	��ېڰ.v�8��_���j"��t+29B3rv6(F���)=�,�F6���ȣ��	û�r�ksmG��u�����m�R�A
m��
H�����AGRڳLq�YH�k׭��m����ۢڴgZ6°�:	��۝�e���-)�����P�,��q¯[��$��d�Du��mZI۰��NIf)J$��P>s�B��oG�'�
��A�]2|�F�r]�d�gǛ���fCu��J��|Z��A$�NDo5�pj�ki��o;��8TwHA���$�.3�5O@�WcT�m�N.@�	��ZdH����7�&&�����/�a���ϸ��T�2����e,��p�keX#� f���5��+Q�1l�_����]UA�q���ɟW�<���"8$L�]fU��"��̾�� �m�"p����;tC0.��t��$�_k�\��/�h$��ȀH�<�5�:
���j�����L�9�a�'NQ.���S�	|�}T�y��b<|A���E��-�π�s.l�?bi������r����T�D�C��>���^F��.��e:,.���i]&��>e�t��c)�g6�W��[x�c��ۯ{���:7��;�[���Ml�̘ó�5�����
zX �w����A��gBY3�Cl�dy�w���M����#�Vv�x�=�t��� �u �Uu@G��#�z#Ƕ����?��ƾ�4�Pk�6:]m��-�j &�u�1Z&�{4�߾6�����X�eg��+d�A����ӈ
�1�މ�stYǷw��w]���?����L���겝����U,�$�{�û�:F%��yR�|���$��xa��Ɉ�=2�דP ��:�9�:ô�#�� ��F��@$��0��������'}���xА�x-:r�
c|��:tΝ�yj\@2����D	��m��༉���$t�S��z�ІɌ6�.��]�Mt@$H���p�)��-1/��,َ �	��($E<=-��g#�����wP��/e�����.��=�Z�Ϛ�w�8�ds�6�(�_l�Ecʻf���dFJ�R�iʬ���0s$r�g������AfRR,lY����u�ip�<�������ILM�4\,r�Ƶ��Zf����5֚�l�\0�VR���,��)KW�X�$Ĳ�v�ݐ����wa�����!d�tsrŲ�6�dԁ��XCh��fг]�{.�[�6�PԕKmD%s4�]M�G�uH�hb�h�rb1r)&4��vI� .�g�1r[E�[ͥ���Y����L��3̥0]\�Ͳ�c4����SG)W��mJd9�#�����y�]gg
{Ȍ9.ᘱu�4��$Vn�A�s�2dSM����9b}x�S��1� �~�̰��b��&j�����Y"�cݻ��;[� �j7�(���M3�#��x�(s:vg`�@oM?l@�j;"������a�3ݼ+�2!��/�=:r"d��W��v]�ڬ��h%��]�lr@=��������x��\����!���N��*^Mf@ai����Q?d���>���#�ύ;�\!7�0&Bn��}==	ms7z�ץ�>y�p�1P�ڪA8�M	�����1��P[��e��8f�����t[nt��&�����ǉл��A��6_������ I �OD?�h �:ȶ��3W`��{�Z��.6����)u=�/���6�]���_����;�ZϦ�3��O]T�;v��k������޵%׬`F0� �{��Fd�zy�|���׆�=r	ݕ�Ȗ.�f�xZ��bH,;;Q%w@���v�$8i����	+c���P �p����;�Ğ�yaIL8x�|{. K�Y��F|�ݒ	U�%3�����/v�ׂ�6�A��$�Wir���v��y�ǉj��K�J���OEDA.��쾨	;}�1��ڰ��9�1��I�K�O��ӂ\D�0��׀�1���,�4���b&�)������K�J�.�x��@I�Z�/����:n1�k\o��*���Է�F���&r�&z��l^�]�I�0.�]�z<���9m��9}� ��{�[3S�~�j"yZY�"�2��������v�B�����ła���t2ɦ̩e�5ّ�\c�~C�f��g�<�0~�q��OoE$*X�>�ͻ��R���R��tY+�R�R�	ua���aB��=��m� ~��&ngyܤ��~����a }.���|x ��8Q��b�.	�~��s(ՆZr�Ν3�LL��2$H��7�U��cD�P�+<g��_DI����k�j'v/��Ŭ�)�W9)ڬ2��]c5 ��kfk�"U��m�Ap'�99	˒�u�rT� ����F�tW�^G��1Q�M��x���ݰ-�frv`����핤�+e4�$ufDW�y�X����_\x��v퍓�\۞HW��P�:N�L�ޙ�p �+g^������[�eO��$v������D��.)�"��1����\n���	�h�s_� $�H���'�zP;�tĿMv�'�g��Q��wV����r�nN�*X���i���T��kff�m�}�!��BN���王ǚ�n����������;ĉi��uY��$;�H�M���x%���tqɋr�Y�O�Äw��R'ğ}S�C������8�a� ����#��4ii����2r.��l���u�T�ǯ��gN��& w ��	m�DA#c�<�S��z#W��ȶ�2 �V@��NB�����U8�K�s;C��N��o$���<�E�l�͵ު�q���H���39;0\O�6S�&�y�M��"y�!���mvǫ�x��k���>�tD��XH.�:)3��u��P�+9����p$�O�[��2y(�����X�n%��"^��Z��k{Px�����ŕ���"�"�BS����Uf�@7�>ݜ��=T�˻u7!�+%�c�fy�z=M{�x������g�~�r�}�ө���c$C��X���Vٶz�[��,8q]�#X�����5�xcO�f�51�[��a7���BYe}oO���t���#x�r�剚�I])��U%�@	��aj��&%F�,5n]��CZ�I� ��4�a3B�k�a�V�+n�%�Z�U����Y�J�P�:�HJ$��t��Bm��l]�<�YeYV�R��a�f%j��7�#��Lk�A�7�M,�$l�)�ں��.504�2�*6� LLi�oYx�P�a��\�Įe��ҋŁ0�&!��Y�íᡓ8b�ǆ����$;�H�G�:=���[L𽵼�
�e�+�#�񛸁 ��M�G��JΝ3�f.&A:^yO��i\�y;}ѷ0 k�i�Ĥ��2-�WW�^�n���rwE��_�(4�v�M�0=y�o�Fw4C7F`:m���#�� sn�`�����2�ʯ0s��
�P��cē���@�o���0���1�Dy��Kb$�.�g�S��i����^���4�F�3A�SɄN^k�'���D&�����篳z���!�&�s�l���.h@ �V@v���S$�]%�+L�>�~_z]�2�H߾x�&���ׂg�/WWDg��=��2�'�;9���A$��؏�s��@�wIi�q��A�i6p�����a��v������/`�/f��r����"�x��e}�F�����!���E�E]ˤ�ȹ���(h���> �����2�"	��� H�U[dB�5�mZ�	����t靃1qT�� ���E��;Sئ���;żY�� �A��q�:����v9�/M/�:�f!��A U�<��BBD��W�3��S>2��G�I�|�'�N��3�� �Ą!d�	��q�����WZ��ﺀ$	���B��=����nb/5���~��%����9(��L�5v�vťб�"]����Xb�l톨k'�����G5Gk�[�a2�x$���Pm��j�����.��A�UX&�Y�󪣭\�Bêc�*�@��ǠX�Ge�A$��IN���z��HS�aQ�,�NBwt��PZ5�=8��,aZ���	�g�"nc)I���5�ޞIӱ����x���K�X�ܥWV�
��y�i�(3�U,�� ���~�!�z��4HM�}��>i�Hs;�gp�\`�v��ӹ9:�t��y�� �&��� #���V��'A%�. ����X� Γ�.�0؍ۉ'��vs�9����P b��ξ	]�D H$NSق|k{�3��u]4�E�1$�f���݃;Yc�\��ũYk�H�z������E�[�Ȗw���1�P �N�6�k{�\ѳ��0�����7�������\��1��;ɝ��=�A׉��Rũ����O]�$��:���b޻���ӰD/L�V[&w%��3�M�> Vv�<K����R��ϳAv�`�ށ磴�v�gt��
�l��`��-���B�L����&��5��l5��i��<x��Q�R9��Q�y���q��tL��<��V�\r$�'S��T:���#6t�䘖���y�)*m|e-��#�=���KU�F��&w��
�ͳ	"zn#�/�������5��U^DIvz"�t~��u?B�@�!���x�4c括�^ܠ�SB�0-6PQn]�<�m�����|�#:N��
v_��^�
5����jN�t�ht�@�#�zxk^[��&&`Ɏʏ8��o76[?�h�x$��ǂA��>�|o[J�;e��E���7�:)���5��	���@�(Dn��v=q�E����z��p'�eI\�]&w%��S��g�w�%>sS\~����y'ē�9�;k�u\�kh��h�	+�(O��'���;�����h`��o�A����x�٦g���3�l�Bw�}���߽i�������Z�� (���AD����?֠��3���Ѣ����Ɓ," �(�B
,a(�dX"��
�dX���
�"�A���+BB"�dX�� �+E��
�"�(����"*��
�a�"�a(� �]���I�U8�u�NNH�]�㜉UR�㜉Ut�IWw8�ws��U�s�%�8�)�r��s�w8��8�%�ˈ��.���'wt�]ӎ$�T�%�8�u)�K�]J��ҢwwN:'u9;�t듊]r�w].��8�t�]ҢwR��%t��N8�u.�r�]ԺU.�ӎ)u8�WK�%\�wR�].�ӎ�T��t�uK�R�T��t�wR�WK�T�uK�t��R�].�K�uZ��K�A"� A"0 A �(A" A"(A ��<�8	�
A �H ���"A 
�H �*)��A "���H$ R	T�D �EH$��B�J$QX$X$E\ց4��H�H��H��H��H��H��H"�MPU�D�D�+�+�+���+���(�H��H��H��H�Z�
� *�"�� �� 
� 
� *� ��"
� *ډTV	 V	V	V	V	V�V	V	V @Uִ�`�E`�``�Ec# E� E�DU�D� @���"�dd"��� �� ��!��H��	"�H��	"���C��q�
s?7��A	U�@DH��������������w�?��u���:~���A�����G�BZ��������� Q�O���?��EU��*
"�������
@����"��s���B�"+��?Hy���I��Bt���"w�_����RO��� ,"0dYVcVb�c V,X`�`����X�c V$AX	VAX	 V,AX1E`,XTY V@�����AE���$QX�F �"�B# 0(� D,@�� "�E!"E(��B,�P�r�w.����W;�+�:���u;��;�.��wK��:�J����ʣ��dU�dVD $DV0dVdAYV@U�QYVE`@�dY VD�X���V}�@V�b@�EsG��~���t}���"(��
! *2� �$���|_������	���`~'_����U�~T?Ǔ?y��gf��O��8?�����0��&c���U�>�?$�}~�>��PE~�TDW��������1ن�T^?0~�
"�_������s���������a��G��NC �*�"�����?I�!���TDW�������=7�������a���"�����
"�����O�?o�*�"��z���!�H���q�G���~��}����S��%:�xUDEt��N���*������:_R��T_�x`P��("���o��? �~t���
�2��,["�0V� ���9�>���`    4= Ud  ( � 6�cA� l 
 Ph F�h Ѡ�( �%��'��@ITQE)IB�I���*�UQP��R!UU(�"��B�TPUU��!����PERR�E!$|                                   ��   @     #||�[����y�th7Y���6��� �Y�ΥK[��B�;:��7Yҭep 6��Nwr�mg6:R��T*��  �u���(��i� \V��{l��{ ;� (�  �� �`�3`�� ������`(��締 dR�R�*�/�  >   �      �  M�ϰ =�� w��7X
(. `�"� ��L �� u9ؠ <{� q�z���z`�7WMDR%J%K�  ����k�zí�m�5�Ѯn���淬�lm���*�{��ކ�M� ���R��wX����ڧ����=��
�*��{� �        ��}��-N}�:�6�u���Km�n��cp 9���;��m�i�R�b���M2���IQ3p Yt�sw
�)tҧT��=�  L>�eZW����c,� ]np❶��;js`\խ��]4�� �+��N��W#�v���v�KmɩUڦ� BD��           y����aKs���sr
����&�6p�����Yv-�m��S��˭�lf��]r�-8�w2�\��$6���L��!U$O� �{�/��Re��ꄹ�p N�iG.��2e�]��F�v��ju�T�N t�ƝqԵ5��\*ѹ�ͭ�[��[ �)UAR��  ;�        ԧ�.sp�i���m��ҕ�屪� \ʎv�T���Qs�[hU��J�� F�ª�;�(T���E*�   ���6Ԯwu"T� vt*n�T�ػ�:#l�۫Z�W7��9]��GKm9���/[�u����OJ�T����Jz�2 S�1�(� ?L���J@  S��h)J@  	Oԥ)��@  	
1&R��yA��w�������ĀM��k��yƋ|x����HH@�����HH@�� ?�!!K��$�	/�$�@$$w�������۬zYW_ǜ,rj�Q������&����[5Y��f=h+��rH]��+W{���A��y�aa��lf�˩OhDo�U2Y�
�ʰb�W�C���{�c�v�WZ���CmV�{�.=��WH!�l�<���)��0@ӼDh9�X���P�y0!()�1�L���Zȋ�,"��a�Jʏ- �T�[B#�DDF�h'2��M�I��5G�z�fh#Y�u��ⵦ��PSP��tm�K������:���[��2]��{���⻻J��u�pe*�c�[zm���ׅ9�+*<����ct��Qъ�2Rź�-��&Jɖ���Y�2Y�d$ٳN:�c�jT��4���*J��EUܴ�9��V�7p�)���:�Ah�X��dzk0�x!FC�Na���3eQw��A�Z�X�4\�;��n,=P� �8�2�f�Z��kM�٬�`�5kp���5maN��A�IɗZ�(ݖF<Q��n��V:fTr�AM�W�j[���i��ڂ2db"��{���Gדv�p^b��T���"֛OKw��� �A�DT;��sjKE�"E@^��U�Gȭh.����P�p���Y:���)�#x\�Vl�ҶZ�����tk��0�@���3~�
�Uj�qm0�r�զ�Y&��ȴ֍�T 6y��, ����VP��s�d˨��Z �(��'U����sfm٭Ҏ�s2��h�&jW�e����f����bɬ�lHk2���8�jx!P����cUc�(�]G/Uh�Ѣ(�@�"���fLZ���{���:��J�j�*������83�L�����ys�>zmB3[�[tA�De��4�:�Ke�wO�3L�yB���Q��:@i"��1a�U��]��L��x5&3��k,7����_c�w�L<���U��+Ub)�@W���,���6�Lf�j��[�(��{�ln?�!DS:V�J�˛�܏Xͨ"��ݱ���h� a�{�MZt_�q��T��xLoWt��m���tv�Y�Ǯ���w4V
���c�d޷�屄�Բ��j�:�,rGY�
�)}�W�Z|>��K���b�q����/r=�j�*�4��K�����V�̊=�	�(�V��cq����5�y-lҤ�f�Z��[YZ��p�c7me�U��]e�b�L�2� ��Z�2�N�ׄ,��QJ9�:�Z���oY�P]\oB�H��2��V�ʃ�v.5��ٛNl�o�zcQ�X;��7��ZfI�.R"��� h�]�W��.j4��a��*�f��"���4����[��uZ�;[wE��n���f��YF��k-��,�a�B���ʬ.��p��mhf�1��F#�+&]�-�Mۼ�c9Or�]��Do�����$9�#/�yyw�}�&�ͳt6�8^��eǨ:��ua<��k`����Ӕ�P�ٚG�E[J�h�ͽͬxjLVqP����G`Wy� �рV>��D��T1v ����-���el��*
��bnF����c&��BV��⳦�k�MCi'wc��"��vig�R�lh.-�ņ�|��퓈d�I[j�2نZ
�V┤�f�Gbڲ�j�M�v�,�y@p�h^e$&�q<�%�2�!Wy����ݐ-[���̼��:ځ���T�aˆU��cVX�
Ζ
�r\\�Y�ÑY�e�hz��f�n'Fj(�Їf(D��+.�7���F����]�1ʻס*��]��0����ef˼[5le3z��x^G���7%+�l4!����	 ޷��#tkhDֽZ�
���+ yGa
�+&�au��iJ�bAU��w\�7Ϲ�޵uC0[u�M�Y��b݊.��y��Z�v�ְ�wy6�c+0��T�#r��)��#q�L,n�aܴ����
\��wL�cbX/,�%���a���M�+�ޓ�͍Ǵds5G�r6e�U��G2��&Ea@�c�]m���Gjj��t��{-V)��F$��eX�Zw�o����d`X,֍�R�ت�8��V0�J�6R�d[�l:����F��ʎK������X��˛G<�i�&��£���|m�2����>7ȴ�`�ݴ+�lȈU7dں���u���{�r���Fٙl*w�Fn�ī߉'34ؔ˽j�^�t�c'C�w�m����Ήe������f�]�UL!�D7Y�f�%���MU�#TL��nJ�n�������;��l�ē�X�P;���ً#D��gv�heL�<є!���fc8O�sVM&�/�TsqP�\�B�>��wwh��oC2���KXV�XT	g/-]��, �7�mmZ;2�.�8��;a�:�ҩV&,Ҁ��%�pY�2�E̽��:57,ʛx�ĝ`����)�v�]�I�n�㊦�QJ&�]n�2Y�Y���W�6 �6<��N�Ѽ�ڹ�\���rė�X�57.��gPe��w�L$�����O^���B�����4n3�:۫����2�*Sf��9�TlA��wFn6efLw�{�-��U�1�Y�b4�k�nRh��J:�5ݳ�S4Į�☖#vv���֍L��fKr�V�s�T#�d�=�q�D�L�B2n�/�kh �+i�f@U��t|'oT�V�4(e],��.n��V�-|2Kбn��Z���9�V �I��Csf�뼵O�ն����.E�E#�ni��4c1T�C,;��&V�Y6���kՕ�#6���9N�ym�̱uxhF��U���5��3C5�/j�5b �L�Ǐ]����v���$�Ǩ�3�ƍ[6XHs�6;)b;{�i��=��<p�`=
Lqg6;2YS{�w&aTYѮ�H��V�	%�r�K�=ˋFmiRq�Wd����E���YO5ˠ�b��((4�Ak�n�m��@��5f��{[@YYFk��y�+�պnV��.�,T��y�4@�V�$��K���tYx�1���[�5�å��J�B�CE�M�]�,�:�b<��,b`Ո�]a��1��ud��H��U� ���rһَ�`��3SH�[j�a�ɩ1e�Y-��n��[��|����P�:�Xպ2+-djT���2ز�ELX��h)����±�+��q[���'Fc�ǴU�'f��׃*�8\y��|���9������ݬr�(����6i�:��V�˭x�@�xaYWd�أ�����������ށ�����$�'�����h�#�����Ѯ��5vnM;��P�̶�Բ�K>qZ6��a3HK��ղ���t��(QB%�sj3-�h<�nb����.��C��Dû��-�J�bic���]Zkmd;D��o���*�Nj
�T{�b���f����[J�i��JѸ��ܺ�{�[x3�F���,k���!]��HX�E��	<�-O42=��&'R�<[���1yֆ��N����7g��P�eIN-�B��a�&�wR���˵H���ܣ�]�J�7s&�ʌ�N�*8c��ɴ\�vY��ss6��P�)0�%��3�+m<ݲ�jPO.ehܣ�u	.V�ĳ+Z7���8���jaD�'q��-9��Ue��!��Ŗp�2�*�^'w6�jz݈�uaм�@���H�A��+-�'�����J�5��/>˻{F�n�FsV�5x6B�\7a�g���Fm��@b{�WaS��m�G6M�"�ٗe�yd;ekZ����͛�ZH�Ӹv^���p�B��T;��ݑڠu|�\Lm�]�,뙔�Y��3f�w��AQH�2�ǣI�WwP0+6'��k$�����4="���{ud����+�\݇m�-���q���1g�6f�M��Z�h�W{�`h*�/,�&1��zԣAVQ�Zv�Bdu���Z۸��t�r�)Ijӊ�W��ɰ^ӫ�r���ֶ��N��KYf����U�"-�O/-/�ekS�ei���@�$�W����L���3�)�2�%B���k�ajl�F�h�&���Q܀�7Cv�GyS2��I�m�uc��R�X�@\ �y��ѪT����ߤ8��q]\�fi̗Y4;V�GM�ܱ��(�������%�]��AL*�� F]a�f�E�Kzr��UҺY�ۛ����Y��k]��`��ӫ1\
��EeRݑ[��������.�Ք�"ŭഖ�C�R��@+K;[�D�Ew�Y�W�H�D���j�ss��]�����Pfe�F��o�x�R���<@P�F��8�u-����(��-G#�[��f���1�*f���"�('���� �ݧn*AXw����Y��lfb'n�]m�0�)�
T���?�A&��A�aL��Q=F��m%��X�5`��)(=�����1l��ɵ�b���X�X&R�F)�Ǩ�v'�obj��ᵥ�vmFj�e݆ɹ����V�QT\�le�5�ݙ"��*�@֚I�T�o3
$����d��.���M���N�hf[5�d&���Վ�F|#l�r�9�Gqu%vX���J���h�)�t�]����o��Lc�x�7��A�t2�ޚ��2d�k1�!6e֬��[�Q�IT�"����*R�ȅ �PU�em�r��U���5��%m3-U֘^�/��2�j9oL�%��X7q�Ð��/j��5"؀�S��r<��+lŶ3fV]]����۠����
֘�V�J�;6��U��`�Kj��s"v��Q��]:�����hWn�7�� ��n�`�R^ӥ�*p�i�he@�TÏ.�fR����'�l����\H�͉f�ݰ��R	���*4)���*B�M�*���X�UF�5�8!�~R�4��YN;��ׅGM�t�D���w+T"�N�xu�^X6�.�����i����k�s~���)�ȳ>�n�,ɩx�����KS^�˷[hIQ��o�dq���[�dyua����ĊF���n(��vB2k;Z�S7��h2��-#(� ^��f��X7�'Boz$��f����hfQ;����UMb����1��n��m�'�ɱ�)e�c��On�k�h��Kb+-��]�s-�f+m���87����,��t���Q"!�*9��-��r��E���з����=�/)���6����W�Ӓ��w>U.8~��{B�\*�����Z 5�@��x.�AÛ7{�T�J�4/3Yunլ�y�L��ӊ�C��J,-�b�W���f;EZ�R���ѬV�[�sr�m㹮:�J�I���$Q5%ǥ�,k�\�:��hV��XV����Y��n"�p�sr|�׉�`�ʑ:���[r���ujX5�(M!i�2�j<��ݙZ���
iie\$�B���V�ڵBB�)�4spP�ے3�0�c�B��f����+^��J�E�si,cv�`�#@R�=zoP�sky�9$�-��G��T�bZ@P8�5��2fڐ���q��TW����fV�-��!b�V�41��n��qQ�kf�n�m��r���]M�G�x��|�[�\k�����Xss�7,�L�!�0�0
�v�ŽLØ��������¨�yq��Z�K�;��K�(�>'+)���W������X
�w�=
�`�6��-�U��j�M�Y 2�Eeo�,,�awL+�X+���}]I�Hm���&�\�/����(�5o6��$�q��9����1�X��u�xY�ff��p	R�%F�YZCu�w6�3`��X���Jcq+��=��e�(��٬Ca֢�
���ڸL������ �-a˲ð�ܩJ��Ù#"P��\��YE�ܩ���1�W�E;˦2����}Z2ȫw����,�ʩШ���
��D��	wJ�jfБ�b��,f]Ks&ՠ��@3�V����	�����i���ӓ��`��S���e�J�K0\ūv:�Yn�����ݛ�ݾ�d�w�ר�[�C�dɪn��;Zp��nbA�ԥtoXf�ɒJM^hُ17�[QҼ4��Ti[�R+�{D=��
R�Մ�t��c��-�]M�n�Č���ڰI�v�4��f�u,���Q�2m6��&M܋ndۼ���/#5q`�d�T�E�;�
�+.��i�6���^彻sH��}�j����c.���� /�1�-& � Ck6��������{wr��^ٴr���R�V��jga�H��4(e6L ��tF��5�0^���"�=�m�(�4�{W4)��iK��ŭ���]��XNT�{������Ue�1��z�mm+z]�@Y2����U3��w-����X��幛AM�fR�q�z���Xrb�T�z��4���+^Փ���٫U��2�ZWx�\�ޝ��D�~9JV�Y ���^��̛�v
v������|��+Oc�՜\ŵ��e���K�Y���y�u��kD�Rka���B�o9�l��&Bn4�%���\9u���ը�Z��-L�`���+[yW��Ǔ,�Mx`�r�ڸ����[u��3k
�RZ��f��֩)'���NR�:�'w3d�A�
�RH
51�aʷn�_A�0��.|�kF5ZL;�ȉ֨��f��v�$w�]0ŉ�P�]n�ḍP�=.|��1).�5(7a�Z��Yrn=h��k%��,�R���զѧɺ�M�K99�a�t��5�%�X�2�Z����	�6�YL���*㠋�M�*��Y����w��`� ��9t�87���l&5j�5�Ņbe;�[Y�'Y�*�,iV������j�,Ab��1uĨ�yv�o�ӕ
;�P�n��&��yPVE�n^8.�(e�Sb?����������+��:�:���;��b�㸮����.��㫺:��.�**������컎��:������:���겮�;�M�M�DbJ4�	�M�U���q����wu��X]U�wE�WYwq�w\]�w]wEU�]�gY���u�wwt]weTu�EWGwu�UeqWwYu���Quu�E]q�u��uu�u]eW\u�\uU��U����Q��p$hHhHm��Ā.�諸ꪎ���:��:��㺋��ή�:�ʪ:�:�+�.�.����:��:��ChH� $� Di!����@�HH� �$���l�~���7��G�(sr�U)R�H�GpuTڻM]�����Vq�)��,Ax��v�q����܀��lܸ�d�e�w�Ws��F�N�4�z�K3��uo&�g#���;�H"��+�]�u��'�s��4��EX�T�>���j�g]`�Z��PLK�s�_)�hEԞ %��j���N��1����6-�9X���EX�_iY��r1%ˊ��=��u����ݾ �!'�qX������]RΧ*�/b�sr����"������&����e�@�Vh2<0���lwE�MgiQ�+�ݡ����S�-�ic�������NE�T1��@☮�)O5=�r���<��c����{�w�3+4$��:��\�"S����U0B]ø0`X$Z6�y��ٻ!tް5�$1fR�Ai�r���j=��m7�r4�Z�!�K.��
�>Ő>囐�v\����D���7c����S8�̜�J�i�Q�Ѻ=l��qΓ��i���Y�V�D6f��cEȱ|+3i�#o2��b+�z��(��w��)N��j=6Ej�8��5b839�4�_w=��u��v_�ر�6��q}k.aH�=�ow"�s2^�Y��R��W�w6�Ͼ�]���o,?UT5��eQ[v6ȭ�A�Nx��L��;)�IWu��s\�ᙼF�ₕ�2�b:�g��4�)��X��Myu�̙j!��],��%V�1�t�	��
��2�A������J(����֮i��7���ʻ��LZ�����八�o�3R]	X]��j�=W����?��`�o{�ݞ�+��o^�?g	y�V�n��Z`�l�X���S���,2�.�U��@nb7�r
�����\�B�	�ޠNeLߢ�����7��3����sD�9x{nN��1ݷv쁘�y��۩��Kҹv+�GU]L �J����+p�P6��0a��}U]�I�K#��/�پ={��r�]M��wr��}�\���Cw3��b��Z���X0Z|�U�\�������ʩi��q^��\71Q'%��*·b2�rU�s⚙X{��I.Sp��	r�O_n9������H�n��T֚A᮶���t�k��Y�*	O3E\6�K�޲�-l��2U��TPNrŸ8��,��J�@囯:d�kJ�"�����v#&��M��oiѤD�jKi^�@M�5 ���&�q�QI�fsK�v�c|�$tnkޥ\*�W3�DX15wcx�ɺ����P̀˗��+x4�f!��8
��o�e:T�M�]��b�P�zP�[!�
�Z �1�[2�<iY	�ff�,n�o�6>��MIY�*��n>x�m�ŉ�r��él�)�T�	[s��jl���}t�m9=��\fb��cf5.o]���2�+�,܏�Y��� ٯd�,+��P�x��R1].$���d��!��a��W�e�e�]�v�y��k�^�8p��YoP�޳8r�u[G+gRo/�B�ӏ��2P��f!jnr=1�pY\�6�>�QY���tX�8�(u�u�/m��Z6���&�l��5i��2��>&h �n��Å\�W/x2Vo��D	錍t/�<�ALYb0���鹐�[�j�\���Q�kL�뭛؜f���nٯq�`�ű�{��tF��ͩ��+����ڂ�41��wղ�&DOh�����q�%�X'X�4�S���Xɛ|6�45��noqn����F����/*r�3�:���[y��}�r��G/q�7	�V%_��ik�s%-����ʹ�=�;�8Y},1�L2e^Yy��W`���JͶ�fՓrc��+�c�n��󮷝�7�fn�P�&0��c|����l��ڴqvE	1(-��*�:�X�)�ۚw2��+-��6))��c��|l��x��UJ��nnæ� f����X�Qj�|�T`���ՌP���ʺ�)�zí�M��MX/��}�}�*p�3f��]�e�OuV[�o��B�<�82K�ξݺ�|��JXf�`��\���)x-����MR�DH�w]�n(��IC8��(V��UHp$bic�0k�:�wS���Z.��xsq!l��Ĕ�z�6R:*�ɋ�=����ȥ;�ԛP���'$}r����wR��@�e�k���9�����y���f�xwذ���m.c%�z�]�u�T��gfl�r]��[L���Q_n�J�����o���M,�8�n�]Q��C1��S��̬��j�L�k6�w��
���!sGk<lwnΚgbǪ���cE�_}�.�N�#���T^�G��Zn��kbÄ�cdu���2+��e�W9�a�j�8�v�/Z���٥p&��^�w�b�5u6��^�j��O�q譞�Ǚ)Em7�Oo �	�x�^�mnnYRc7v��۲�H���k�P�1�mKG[��u�K��"��1W�;xLRkSľ�ġu]��=O-�bpy��E��eu%��8�E��Pڧ[2dӲk�{{h�w�ӎ��������\�*.���lt�Wa*۲�}��ݦ>��Nb�$]v�'$���n�m�������nG�u"uu�n����lG����DwR}��K�b,]�Y�)ի�8�ݼ�wk���u0�0
������T��4֙F,8�lF��۹Ẋh�i��^�z�@�1�Y�)[���Rv�um��G>ǝϳC�5�	��K��-hQ�;n���܋G��*X���v�+�h �oc�(GS't�+��yN��[�+����U��sD9�f���n�M]u6�r���sO<��b�h��j��	{������:u�+BHE�\z�\����l^�͎X�Fs5��IV�����̷����g�Deg5O��lZ�[�z��*ͬۢ��7vc�k��Ť1���q��P����R�]Lj��Oo�s ���:�=��Z9��6��q��\˴0L�%eq�;��JM�d4;6���Y�L�(V�y*p�3�\[��%w��-W+�W�)tUg"�]��ͩ�[%�ݪS�i�1)�/��H/^��!��h����3G\1lR���]�au´y�.�n�n��ѪS�QZS��۪�Q���ۊ1����c��*WW(�9�.�\rf�����U_���X�_U�\ެ�*�Ik-tu&�j��+C��0m��L��R��7;�O.����F0A;޳-[���sj�_����8;+Zr1�V��#GF���'jE]�wm}�Ǿf��)&����_,��Z��.��MӰu��@�N���K�I&���d�v{;�n%��n��I��N�5�rw�r�K�n���3kT�M��r��\�+�o�L���8��3o��u�����;jX�|z��ڹ�ۚ�V��h����gT���w�^u�TT7���.�eZ�`'[u�9���T
L0��y�6���bΫ-�Ɣ���Z�Wl��Q*��v����ˬ
��j��?�WUk�`�e�T��{��I�zTh�,�2�ܷVk�n͚H�Ec�U�����7d�}v����R=Fݔ��ܧ�]+�n������V�����ߖMb��u�sv��E-�+��N{f�m�Y8SW`���%L&� h�%�0D���*��mX�-���ZPƣ��⬽/����a�t�$8әZ�v�^W1���x�U5�6��׀���H��r�u�WB����:M<�5ꉩ�M1�lu��F���XBq��ح���D�ն���j>qs�7,Z׍PB��R;uO\��}z��<,��ڳȂ6���wX�pg)��ɶ�t�fd���Q4��n��+ٕw5�Dt�|�g�X�qVPP���<sr�#4�ܝ\.��r��m���SĔN���W.E�wVr�c4��x���:�K��l���_Hi����u�M.e��	��jӁ,bw\�u�f4s#:��ՁKWQU��8�6:�m�x��O���-��]� �k:�t�� c���FsՖ�c>ӕ�|u�J�¡K&jZ�EL���D"`op�-w�o���GF3H�ȫ�!��/�D�wg���&�vi����P��KB��J٩�R{ϫQo�@�A�B���s��̽r���a�F���nT�ӅH+�ɣ�-��o������Q�7zUw�$'�1*��_k��ebG&;���nt�-Jt��!uQV%e��-�cT9D;v��_U��Y�Kf'�R�q�6�=�J�aYB;��:흭�Us�6Iq��S�wT�dK�K:G�<�:�7��da@B9b��SNV3��ڨl3�O�hu�7�v9�V�;�!=d\�Y����l]�4�Q��X��3z�o4GV�Oj�8]���=l[����OGN�eL�����1Qvf��`��D�5oiH]�ޖ�X$'�K'y}�b�cחgv���
��
�
��/#�Dp����� �عX��`�d11^�wJAtљB�������S��VZ���鴷{7[ycw���㳦^8��F�M�&s�]��)La��5Ķ��	c�'hG ��l� ���;ĺ}W[jP�{h�ð��!9�WP'&n%(�0TGvR5�q#2�v�;���|��[*��6U�/��ѩ�:�C3:�+�T�&���o�Nw5�[�����n�7ΒL�7bqt�Rw�(��=�4�@��|e%���P^
�~F��uf�v�tJ�*l
��V�];Cv�6q�eDԒ�X�.|{���<q��v�]�P�ondV�5���jAA�93噥&��UCO��bT)v�6E��T.ˑ��w�vU.\yD�Y7�{l�'�<�ٜc���]&�1�����]fg�<T�K�K-y��{Y{���+�v�q����4:H���y̝�z۹%�.HiG�讎%����7���΅BT���.MÏ��Yy;�D%By��;�0m�P�P�Υ��=rŘ�P-Z��{��Z���<f�>�Ĭ��*V�&v��6��;�?��X7�MVko��k�5�t�sQ۫Bũ�j*��*=Ἲ;;yRCF�胭d�
]
��B7�T��y[�^`��8�1���ܼ�r�Р��ae`9���Ăm��n5��^ҩ/*1�����{���օ��w+�7#v���֞��LK�J�&�͐m9�u�ˌ���C�ح�A�1�U8��	���-��3�,�(lyb��wT�;.W�el��Ѓ�W�Cw�Ԥ+��lQ��&�o�kpi�f�qP���f��*�n���X�m�A#��M���Y�Ә��wn��W�m���������CM+�n���W�n-�d���e�/��q��W^t$SJ%&��ه�
�Q�o�ʝ�L��a���bٴ�ee�����{%�-�w��F�h�c�k>������������JM�t�:K��5z��k��
d�Xz��4Gu��ӡ��Ї����I�J�0�@�yx�Au����p�df�;���P��c<�뻏1�ZlQ�FXt,���:���vb�V�p�{xK���(�vu�ξz֣0���j���4^.iK�I�q��{�uVH~�K�,`��+q��	Vw3�%ʥ���{����v�A����z�q��Ou�%9�X���l��x漡a��+e��d�w��s��3�h�Wu;���we��Sph͝�h�MI�$�]�c1o^Q�]��fc|�{]|mU�f�򮻸�ܷ&�֗�
����%U�De�@�K���΅��l*I]�n)XF,��x�έQUז��X�\�5a&����ywSVi�U�k�4]��
帯o����ӑ�Bi�ʽ�_p��M�[4uo�.>�z<�V
�1)����;��b\3�2̮ͼ��*��!VQ��QR�$����T�$�E�C�P����b�V��v]"��Z�/������q6�d���1I����q8kQ�&Se%:�r��7*]S�p5�A8��� �cb8�^R�/���sb��v�Mm�}�Rv��ba2-��`����eeZ���)q-�o�'��U�k�#ʋ������c��\����f�V�4
�o��K�[��)u+j�r��f䉕,)�֭�OU�I>��*ŔV��- W^ ��`��_gF�)N��|&���V5�t��ʸ6�����0�eL��}1w�\.�ypZ��
ڻ�U"-]������d
Z�\����.	�@��%��"����Z�ٵ�V�0�AVU�V2;ǉeQ����4pWkMhIV@�b��%0�o\���rcY i�_;S`/��4ɟ>�n��S��OJf��q�]!RwP�# 84P�s!��J�-wiY�]0���.�m�V�8�u,�~�3�^K�����W�W+<Y��n�.Yp�g�uܲ��c�z�l�a釜jٹJ�V�'+\sp���<GP}v�ms�V΂�w��꽱�f�Z5��i=i���6�M%l�ug`�	�9�Y�*򘓶�]
x�"j�#�&T��3T��n貭UT�/-�ԝ|���.���g\�YF[�����A��,w�ZX�{�b��̐��q`co5$T��V�q��)��sk�6'�D|S	��X�l,��a��:�a�w.k�UVL�	��!���/wa�;Ra}u�+o��p�+*�k��.f��k[��ʙ��/m��)4�3�z�� �F#�sFc�M�Q��Z�K�����x�r�*���Vj|���j�Cr�[��*�4.X4{ڥ���[���r�F��O�ɽد�ǅt <��ч��3�	�1]�m�WX��ꛚ,a6��\�y��f��E�-#�ir���e�x:X��z�{�7��J*:F�i���;_C2��t�#�����f�#��7b�Q��H�|D������6�]S3o
2Tu,̒f-��׭�����>5�pB��������\��r�qs��:�]e�ړmsau��u���r7�qۛY��1oT�ѮD'�l�Є�:�k��Dq�#ryn���u�S�I|��&�L������vѪ�e��q�xv�����©�L�]]�a6��}QXs��ǋ��J���0�y0-mx˻zSP�{�l����݋��Kzn��j�u�`��n��J�v6*ع��.x�z��t*S�vID:9�O<��=�����h
4s�籕�:��9.��"�T��qu�o]���p޹ŊwGav��8���)b�;s'X&Yp-��:���4�N�=�Zܻ��cN%M��9�xwfʌ�S�q΂1ض���v<Zb湦ub�ɺ���k���s��@ۨ��;=Es�BK���F�>۫<w;��V�ո�ي���P#��OQ�v�.�w1a�v�v�� �1J�ȯ8x��$�'����9�`����VV˱�����1�DGN<u�m!Z��q'�'F�ζ�+q;
��3�F��tWg��Oe֎5��Š��q��m���q�".�F�ݷIx�v����9���s�]g�3���{����=��mvy�۲�v��^�`�
sֺҡ��S��&���ێ�.,��.�tn:�d�=�n2^+���t�˘糝F�n=�Qnv�;&�%xxG[�Kt���=�n�ZN
:{OerTe:|��65�>��.�ŴuC��O9ƻ\���������v7a��2�r����l�f�+����j7is�u����3�6g�\��n��l���ȧ\n�.�y�x;l&�m6&�AK�:�q��7NӃqn8����p�X�p�Y�[ް��.�6���ݕb^lvN۱K�M��:��,z���̝��j�])Oݭ�����ͣpn��;�h�5r�i���!��e��'t&�ɹ{a%��W�ћ-5���]��6����M��:���e�#���][;��q�ݶt�)�՞�l�@�6D�ǫ�5��RS��lygL�v�1���<s]�<=��О4�{vL�K��E�yw�M�ڭvɝ'v��M�a;w��z$qm�m� ����c��Gmo\���v�;N�}��7hSN{u�=�]�wLMv�9֞:;kz;p�7h���:�歚�0����q�-��[ٸ^���v8�Ok9�8M��nz��zW7�"����ƣ`fyk9�]�Hz��p�uC�a7W!�vq����v��h�&�\v9v�{�/8�O��p�	��o9w\;.m�[>wc�m�s\�q����`��=���q�g�K�}�.�A��Ğ٠�!u��n�ۡ�d�t��7<���B6b��5F,��]�4�^V)ݸx����v���0�E��s�Տ�\��t<2E�k�:�g��=�v�����m�47e�3��[R�s-���;�����3�	M��v�â$1�n�M�9�nz�hW��"kή|r��^mʽ�g�n�!�u�덎\+��v�pOn�A������v�A�6�e	�:x��:���\�w6�Qt�7(�F�+�x6ۜnyܪ��FG���K����Q����c�T��9�m��Ƃ,��n�[��+�sږd6�v�d:��{�qp��-�ð)�v^�p�Gp�0�:�������cx��6��軈iX���	vZ�ȍ�Ц�ϷQpUċn�Q����e�u�b��Mh�e�5e6y��c�q��"��>wM�nΎq�iS�݋��J�����{����N<�S[�́./l�����՞p�Ć����꼝Ʊ�����q�a�;�+��Q\�)�
v.��[D��3ۗ����[s7}����7r:yd.$�+u��/=<C�C ][�v{vm��tyZ�t]��������s��W����|�f7#��ۍӇ�ݐ�K5������K���.;i^d�3a�ɽt\!��N䭶u�V��n�h�֗�����[�ǀNgs�n�x��e={vڑ�2@۝O�mZ۱ݍ�8�ݠ�Uc��h��vй�x�{��,��:�kZ��]��.��c�б��Gg�fu�F杲N�f׎�юL��n=�����5�n4�s���L�WY�>����p���Cg�����O�j���ßK�ջ�Q�$��kQ��e6]/�v�󐻋�v��E0.�z����^�u�㫱\�b�y�@�Z���m˶9q����ƎN��O;'�s\Jg�[qn��n8Ƶ�f�qp�)i�Y�:'u�;Mg\qb�(s&����"X�%�e�]r���Ǳ�m�3]�}݃��8�͹h�&��������n�`�;T��s�����{��.�7P��=��=���bt�^��T����u�u�m�;Hgv(ڸ�#{ۗ�����v�l/e]��Y�V��;wJ;��lo#�X�^��6�4���r��t�n
鮂^uF����trKj���C��q�lu�g���[�P��;�����b�ob�<��Y�燫t{y�N��X�[�8�[�m���W�T��xۮ��� �2z���v��s7snХϵ�ۮ۪듊'�w.�X�kg��ݕ�<��lt[s����!�'Z1��=
�k�6=q��t��n�6���3�V�l��%� �ўt9�*�#�ݸW�j����<=�6wZ�	�۵���`���,���������Q���N�\�9�����cl�/]���<m 4ۜv�7[�(��vݞݳ̀ہ�>n:��n�ѱ�����0�^u�h̸7ֶ+�����l���Ŏ��8v��ݗ�aSCój�hw;\s�F�=�V��`�ɯ=Z+���%�ŜNͲ�f0�m���v��p���r�M�O�gۀ��-n��'\z�MS�{Mle7�ڷV{���I\7�<��8��Ş��:�l��g���ö-�Z]�tܘ�s/-��k�'GZ���4�/�t5�b�f�c�c�-�p������c��n{dXl{0lT������������׊f�8���:����r�'F_d�;n�ݷz㱡Ƥ�麰�^V:����8�,��c�����Uٍ'��0��NXݸѸ�]���<[gF��z�v�箎W��ol�G\m͜�l�r��ۼ=�ukyy���8qu��DJ�=��݁�A���;�3�c����T��6���1���m��0�}�]�a���z�۰�'5Nrs���<��ֽ��ܜuW"�nwt<Ae{����gn�s�.���v�eݴ�9n��K/N�uY]�x�r�"�=���G%�Aq�ێIA��:�n��*�v3Le������1�C'5���#������	͋�p>�L����؝�M��V�v���Dr��ɸ')[��ۇ�*���z�ή���x\V����1��N�ݒ�sr{�;C���;�Gڋ;�k������[d�:�.6��<�����
�R�t{-�rv�Plr� 4/<z�NOY�n�=���h��S��݉�M���֜l����^;h�]S�ۊòn��A�+q��suN��H�kd�ƤVy{]��ye�ˮݸ����u�m��g�����ؖ.�@��Kf,��.�(l�5���X�:�3�8�z9ϳ��n9(Lb�ˮƞnR�B��a�z�ϒx����S��kE�rMl'[xڸw��v��\��r����
�Xwk�P��k]n��ݎ��q���f^y���{RX���]����)�P�̇j����8��l��[�n�]�s�z�<�D��p"��ԝ��;:���{qhq�mh{v�m����9�g���-k�屜oc��дt�M�iۍL���K�g�`��ݍ�ˬ�S�3�`8-��M�pn�۲�69�`%{2uҾ���7�5;���3��F�y�8˶M�\3��Yۭ��/��67'mAXݳp��m!�Ä�kLWl[��㞎q{nv�,e���ΆvmA��f�&�琻��c��{z{�<]͢�o��NNw�p��pxw�r8w6��h�٤� v7E��b^+=�������nۡ#������)v�:Kn���;U�%�Eq�Z�Ӷ�n�`�>n*ŭ;�� {s��n{!��gY6��n�n�[m>(�z�mvwV��]b�to ;6��r���sΎ�R�m��[j��uе��.�v�������֫vK�O�֭ǖ�;yu��m�˺Tf^[��ZK���n�m�p�2��yI��&p��q��(+��9+�7wN긩k�E�۵�u��i�n͚��<.�!����7D�@����h:��B��f�3��n8�X2�s���c�Y��C�����C�7I�`��٭٘��i7m�q�x��wAӡ�H�:�n���X���k��DŘ�j] B���e��VǍ̡҈��Kn�2����y��\�X
 �/{<���vod�\JYax6����m��r�F��t�����ݕ�E�;/.�	Pv�{C`���Gf*�[�`�8�Z�N�/Y�8�3�:ˣoM���Fk��ݞ��%�����s�8�n���c4r`�\ݙli�]p۳���a�˸��Kq�i����/lki�W.=�5���v7�e��d�9�'] ��y�����G�B[�sn�,q��v���\�7�y���^\ѷN|'"�s���nܜ�)��軬X�x˖���c������\i��qq��L)�u��n:և/[��nU��z�D+b>&v�Q���>�����H9�&ݼ���c7 ����0��0���fn+]<1�Ok�z��u��)��k�6��8xm�{M�<�����/L���-��lƵ�y�tb��8J=����=v��qW�׎^.tbl�3[7�v������[�ÁA�sfm]Y�Պ���;7j��gpy�gduE�	f�)�}��;���k�-�f�8t(kvQ�I�  ��ۼ��!�Q�!�P�kj���X��=��*I�hX���;8�;��#�8�FY�X��9B�vv�\��Q9�'�cn#���
N8����e����ܜw'Nt��%8�q�XD	�l��GPu$�Iӹ�V�E+-QG%rP�$Ht�G%�D$@�vG#���m�tI�{bNC��;���۱Gq5XEe�Duee��%ÂQ"\�VU���
B�ma��vv)H ��pG6Ȕ胡C����$���{YI�\�9�rqv�:H"�H;4���=�C�Ģ���:"IÂ�n;�B��N��K̃��	*8�9����﷾�F}�v[K�[�
&ި�/��Ռqh�u��ks����;e�s�v�B)r^p����k����F8,V��.��k�<vic��:�{��4�.9�ђ�7N��ps���E�H�#Gb�r����-ݶ���2�Qۅ��mգ��v�ʽ{�p����ێ�^�QX�콍��;��;n����(�iq�ay^燮ݖ.8�3��x��4��wl�pa"@�l�׷/F\��^�^,��G��Mø��s���'=�'n�aKl��6���n�^�˕a=z���Y���WuY;vh���d\ۭ�1�;��&����u��������m���8���cw�8�B���w&z6���pc8��[#Ǥ��s�|űH���Y�|����a�:7kQ��(�U�C.{����n��G�!�������og�c�5��tc<k-̀M���4����/�w3��:8�7m#���x݊.7�;1��r�ۍ��Zy�ŧ�k���W����ݖx�1nm�t�1���2��Iדg���ϟ;o���c�ICe��Ȣ�;�˦��!b��p�P�K�*��[�:;#k!�Bv;%�a^�<�M���^�wAl����=X��Dp�ԡ��v�<��ٶ�v�kƶۙ�{88C8�kuNu�}�]ۻ����|jP�g�����h]����Y旎�8B���3EQj[lLܟ!X����V�Qa��9��cny�D��c9��+����{v��ۓ�8�K��,`N�1�[�=Epx����尅���;2n���]ҧGQ�]v��s�!����Ls�knn;8��
z�η��cm�v��k���HƁ��6��y;m��m�-,��<�,-or�kn�mg��=u���o<�ٍtcd�7j�G��=8�*<�{[v�r۠�9܉�H8�k_9�>��OJ
��ċ�s��[W�/mA�gg�ގ.ny�5ζ�����[��{Ǧ9��Í�G#˰���yό83�AUǻ<pg�we7a��
�g�'o�3�ώ|�;;�nxT�����Sw)� Õ���^4�zmA��O^����-�ݲ7���m���zc,m6e�g��ޗ���罡��d�]�kvx}�"��wo;p�ɞ@ʢ(��W{w8샲q���|�{r�!
|2'�H�8�~�HD�]�EW_��fv<y��?�{���(�2컕������$&L߈�A��Pwg��g�~>w(ѷS�q�LP�U=�́�+��T����̓<���T�e] �Xi�鱍���׀a$��R�*�հ���	���.l s~Hd�wa�8o>��y�l���1b�����~�T >��%w3۵���W�y����h�p�TW,U�&�����o{���i���#�_e��S��5�@S��z�p�6d6^Q+s��h��Eѽm�q����+�o=�	�e����B��Jё�W�(Z�����޶�����6�wU��4̺�SC/�ܫ��Y9��k�.�kb����K�a�lٔlg-:'���-Wr^�E��(ZtO��_h`^SRk\�x�C3�D3]I��8A�ݏf��Ԗ�͘�1�em�U8�qr�%�&c\����
�nǞ$�Iɾ�$��o��!��Wdo�a ؿ\}	 �D�3E
�����W{�����I� ���gN�	�2o�'}�����%����E���۞��i��}� 	{���O���n�|=��/X��u
\���L����B�+Uc>3�ݺI��ߦh��0���A�~��&�n�O�~���vF\�p95u��98�-�N�EE`�ڃR�:�h��9�v�v�,�6|rj�F}����ߪ����:E��!�y��ݳۧ�H${���{n
=�5�}�G+{�P��n�
�	|��EX4Uҳ�o��#�8}dyɴ��\�v~$���$�����:7Ƥͽ��ӭ\�ϴ��E�E	��8Y��w�k�󙤂7�x�n����	��p��SF�e��Q�v�n�=�l�f����̡��9���{|M$��U��I�ѻ��u�S��2(t�4:�9���x��f�I�?n����"�|M���E���$ڲ^^�.��4�	��A$�n�X=Bvu����v�=�	��T5�ACto{^�$~y�6�w�g[���#�=�:��h$����2�I����6��Ha���X�V��I	l�d���zr��v{;�Qh|㉲2|-�X��9�z�j�4.����&n���7��~ ��^�mz��v�{+�1��GTst=\V#^����`���
�ؐ���1�����{^{I �M�߉�-�0`%�sH�)����� L���V��h�5k�O�� P��YHi�94J��7
^ߥK��i�y�ii�oF�	��NY�M�ܛ�sk��x
��L (.�� ��ɳ^�nc-gc��W�iN�q�ۺ�7Wk���/�V��[�v1������a�r���1R��Gl�x�_��v�9G}VHB�&���U;�_���{^�מ�@U��t���j�U�����R\���>�m)5��Ki#M��w]<pO)a�`<<�\�G�mh��ρ���Ʊ,��;�v@�O����> !٫(Mw�����듆x=ᘽ���!���
R߰���r�R�"c���������]�[�Oڞ:	��t{6�@ѽ�7q���m}1������d����/W� ��� P��{��Z{y� ����5�s&��s4�����SE����c~������'㸣ϫ�����Oҽ�m�*7��$�x�k��i��N�Sw��i/93~5��>8��d�ע���#�6���Ɍ˳r�]�,W���	��	�A��Ӝ��휗�7�3y/o-"�����f}ͻm�u/9�I�-m����r�$�K)f����&�7��Чۛ{NKe8�V!�A���+���m<�]4����N�����y�X9��R�맵Fn�uv:n�j�.�y^�$�ѧ����C������%i�M�K�'n6Z�]z��7��_k�x��k�ev�qɳ���!Mm�lp���m��nKv�d<�cP�k��؀��77�o\����K��ܒV�m����>Cc��r�oG:�8�:賽UZ�]{7$Vw��1����ֻ���8��F%]�߅APR<ξ��VЯ��k�v��� s�l �{[������7�Խ���ɣ~��
PD�$����y�ѧ�tU3n��>W�(�	~�7@!O{S�({ֹW�ޚ��cJ���[�9f�n+­>w7�,�����M��O��bw�yԵv�������L�����A���s�UUV2�1=�g�r?>r�"�Y��_�I �����I���s������kɵ6��󎎧�QV_v�>B/,���C���Й�j��� ���� (!��I�0އ7R�㕊~>��W[����QZ�]��a��q�k<P@����X�>=���r>�+�w��s��7����X��ϲ�������A��߉!E�$!uvE�J��l�,��:6�W�Қ���*��ߊ7��HTꝹ�eY�X:�1�N�e�,64^�̹=>������	��v��'U1� Q�tt����
����#~����"��8/W�*D�4�k@ /��������6d��}{��J�ٺH�������Z�B��*ѺV0���S�~���(��� ���}k��՞Rt��Mg3o�F�g���셳�kb�N����Ӽ�bٮ��g�0>�+U]  ��������з$Sf�"����H�����66��	��孃����>�-�̤d9�8+���ZqѪ�W)뗾�m6��wJ6 �Oy��n���⽃3ӛ� �f��+�]��$�8
/y��-8{��v����z��m�( 9Os�Y͇��[�x�B�THB�"���7k�
��:b����9��nK5	��[��<r��l�B�h^S�.�<�^q�\�?����F�X��'�� �O�s*bͼ�mc�gW3I�Y�(��~$qo��fw��$X��(�B���M�~z�O��6��%�B�Ғ� ���w�w��5CXt��5?5T*��5��]v8��aV�}��,i�����{ݫ�f��TH~�~�6MH����H�f����Z�D�(�Q�vm����[oh�t�sݱA��[c
�t�#���S��~|��moy�f4�i{�ͱ���;���{)P�-����f7:�Zi�P�\�����|�kw�����+ ���T��so�s#����A}Ǖ����h�TQ��T��-N�M�4�PX�fZ��^0
 ?o��'��s~$�����,��Ö���E��X=�x���t�I��t
k=[��g����5�g)��$˭f�$��Ջd�l�:����Dk��j-ݻ�����z^��*������]�أ ����#��7����������So��`P����hc��L�)��jb����� PZ_��.\����>r}�c/݃#N�V�lN�d")����͂��gX�+!��Ԕ��Q������Z�e��Ϲ����	��S�A���`nռ�4��<�� >�{�`Uy��9c(�R��ߋ�ה<65=��ف�y�n��|_�]
g6y6��7S��LQ8(��_{�`P�� 4&����y� �H�~�v-�
>�Ĩ*��J��lL~�iS-��~E��πnni ��|�/��c&yw(W��s�٘���G�&��-zI�F��� ������B�F]�(�����~�_��=�T��Я�!Zk%�7�nǪc�$X�;�=�L�\�>-�h�c>u�+�X�(���5��=��|�wfn�7Y1�N�v(ہ_^"��30��R�p6c]����`��V�x��2ۭ���n���qc��8���7���K��a-����뗧=�Lv;&�
�g��v�Y:�2bcm�톥��g�s�»ne���AqsY����*�v�#ss���91K�!r4���5X�=#�9����l1̓�%�J�B̫�����ce���n��RY��@�uSG3�m�OgS�zD�;�%E���rlv�n�����m��K�Y6x^�J�D�������H$��Ub��2w���Ok˰�yg�� �����KFb�K\L��U�y��I��C:��z\�|A���,$�}�M�FJA�Q�ؑ�/kr0�҉R�h�]�e��*mX��{͊�^��$����VVw�I �[�	"��7I(���QV�v�W��g_Y��y�G,�$֬k ޞ� �g�۽4$|���� z%V+lJ*�ѻ�7gb5�cH$����<9i;��Aj�@H&�{۠�g�ۺw����*��RUL�M�3�8�Y^��q��{[�v}�&��k��M0����s�5� �Z��֍�Q���;��P�z4��/�+�{ �F��6{��`zR�!Hn���׺	����j�区�D�:�qT/�w��1fE��mG����ʗw2��*K�}��S)�,د�G��F�ԩ]+��AU=ޭ��:�^k}(�M�&�=�m�*va�.wf���u�Ja���	V,��^����@>~����4n9�vy�𠏙t�gw�� ���m�y��#�E�����Y��]��v���˯f,$�_�ۻ� E�M^��u�-�b�/�o|œҏm1�2�JW��w�����B�s"�>�h5d����Ӡ �tm� )q~W�:V\��t/${��l����pT��d��0��F�<ϣɬr��ĔTvee���"$��$u��>��X�B{�T����=���K���n��ލ����i�9�˼��$g���5�@�7y�>` =�6�\_�_�f�xԜ�)�۞�E ��UU ��n���|� �X���ʔ��(���\������N�ו)��h��V�"�b�3X��Y����#��1E�y��'��,1X�m��zZjmD/�Ä���i�fn.Ɲ���b��0ە��6X˪�u)|,�#���P��5�k������&�;�J�;�+s#�v�2#���R��&Ħ�\s�J���8n9��Q�l�y�l�G��7��qZ�݃;mۋ�ay�r���j),:���w�����+�]�n��s]W��s���u��y8�	����N�OZq*Z�b��V+������)�&r�����[��I���S��lZ.�2�I���&��Q����3%s���C}��c�Y/C�����E.��b"٥��&�T3CWq2^KR�]Kq�b��ۊK�c����5�P�٘n<;w�PYݾy2EB��[��R]O��slR��㺹<�r]ި&����q^ս��R���烜�WD�-�fѕ��[ŕ��)��rmr �r�R�3�����wV�թΨ��oRXr�_�|j�HN;����cM)eI��]>Ǝ��a���#wz��v�r��ӂiL��l~���!���S~�n�������C�3�U�kvp@����B�<u/���a"��[��nV�e�J�]:�,���N��_<���̳�d�}�W�@(�fu�7���]F������iG�G�0p=����Gk�T��qe>�t�OovW2�y8�ӷ-������u6��՚@��y;z�$�&�b�G5�g��v�AB�{K�f�D��׿7����m�"-��]����h��"��mC����v����,ġ��5�)e�H���mI8t;5ygA�Gm�:��!�dyv\q�p�:qyݒE6��8���' 9()(#�N��@Qͺ�	Ȧ���6�Gq�'Ds�$���16�M�kpPD�ttpH�H���e�ۅN�s��������P�2�U�vgM��B��"Skr'm�q-���iȣ�vMl�D���8H�s�mÎN8�)�8N�	��)�8(�,����f��(��;��NNk@E%�ۑ�֝$q��.(���9�3s���n����Z��I�$Y�i�ps�prqEwp$&��r�U����WE���ӹF�]勠J��"�է}��{�dy����4�~$d�r�I?\�[�Y�]o�m�oy��^���%
��Kfb|񽯬UC�͞A<�+��=�D�� �{r�7�9�z͜i�uk�d�̤M�VE�{K�\��^�.Ӷ���s�;vu��ݠy:��'[���{��h���R��wZ�3k筞�G� }���P���<2zg�k��>�>�3Rul�A�:&R:���=�ıo��e�f���ݚI��{VH�y��I�mE�S����*�/�d9���WkϨ�o�&�4��<���Wmk߈ �/n}@�/�st@y�R� ��n���ƃ~�1��C��|�d����������'�s;�2MXU6�N�z8�2�tͱ����Nh���w���V�M	��\��X����� �;bm�G�%n��Fy�eg�
�c!̓.�&��u�2��?6��P��4�;��/y�R�_�ՀH6�y��	�<�_���W��kد_&�R߅F���4@g�X�fŮܽ�-�;c��5�_����B����<�B�`�̵����C�:c�>���zd�V�g/�p�{|�O�{~Ҟ �5db(�Z��{3��ăӽ�R��jp��I ^���$O^M�A6)7p�^�V��^����g��>�Gz�`�H��1�݇\,�����M��z�n�x�� e��X�����MU�/G�M��Lo�4��٤�D�f��yh �]�th���I k�w�����$G�ط�4\����	����4��=�A �^�Ǩx��A��jLf����W�����,��6�|��4��W���N_cFugq^mW����x!�oء�޻Wasx��s�^�L���%��M�FX��l"�i���`���]�k�I��:��3ړ'b���m˶��L��:\�T�V�6��6�6�<u����=�8�H�k�ˊW.�ݓr{.����xF�S��룡��d�]S��sl����N1j7@���A���,u۝\�ח��g��ƭ�[f��Lݼ0��L���cu��8���������i(q�:i�lI\�y��Z�p��c���ʼ��qӹ۞y�]���R�q�\����%Bn�����f���i��^�   u����	�r����Y�N�(�m��^�o�)vt-R�-�15�ʫX��1�zH�{� G���$�%z��y>�	ι�&ԲxZF�W�Z����O�^���I�5&�����̙�5�]w1����h��A��adu�=�W��/��2�@���piS��~���M���=;h
̛��¨C\l�2��Utp��U�M�c���xA���i�bY/�ۿo�J���GN�6�ޭ����߇���lg��& n0Y��c�{p����c��m���d"n�]�|�'>v���s5�(}׹�Vw��dUԨ&��u�o;��o�9-͕��&�n�>��u���9��̹l\oۗ4O�Jn�o[���3xI�lH�
�\n��MYʦ��@Od'�yU+2�w]$BQΰ�S39��럒\���^��u�m3~�r�7�H���Qu�.�U�G�.�,�e��G�o�$��t���  K� ��n]_�ߺ[���6�߶��AA(�������wn�nG�in==�Z��r�E����\��~Ɣj4�u\�M*a��+>���bF&��{�~�������ם{��!����{w��i#��D8�VG^-��24s=��[A�1�z�^A�=;�se�/|�!��ˤe�6�*���1�M(�Q�{�~��o�����&~�Jk�w�6�]Q������::��<��]�A�w��R%��M�����ߟ���t��|��M��Կ?��Pa�a+�ߩ������z��[���a9�ns���}4_1����ݠ��� ���=�F<h#�çNu��M�l���W�E��j(ԿOF}���[���>k�y��֕0�a�D��ݴc؆Ń=�Q�X�F�j4��+Ͽy�\|��s����U�����M��� �h,+����1@=�ߨ� ��6!�_���^�W��kg�u{�Vk��#��bM\hq�p��;k۾��\��s��A�Z§f��D5���Ρ^=w�M��Ud�٧� ����m��������HưiF�J0����~����U����ѽ�o{ܤ[����}�����\��ֳ�F!�|0���h��iD�b�w,�24q�m�������u�c�v�O�`�#������9�����OP�z{z�����F3j(�M(�+�(iS�v���}���ݯ��F!�l�>��F4cDh����ܢر0�CiF�}�m*Ll�s_��~�7�>��'��e��0e�+���q�VmW:띝�M�tn��C��4�GWv��k�Oo�X>��h1<h#�DR�gr���AƂ8��� �)�x�5�V��s8�9��)�&�j(�>�w�cLQ�S�>֛��ַ�Db{�l84Sa��d�r�ϫ��6�{����Ɣ�20=��(�!��Ae{h4�: ��s��g�fy�c��kyܤq�oʃ�NԐ���h1��,��h�`0#؆�+�����1F�߾��v����<�Ѣ1��s���0�I��oƿ_��%�g5��ABRbldh�v�A�m��ڮ�g�m���$��e�D��#�A�}�e�6�ew��#���(���ۏ�N�f5/5ܿe���)ky[v������vt�+M�W��t�j���=��9����r}�F�~䭈l<¹߿Q�1�4x��;���l��ޝ"�0h��3aM��0�y��0k\����g�����.�##����21��7���UA("DDW��R1�Au�.f��3��#��z���M�Ȇ�8�1ȼ�+C�����[�'�]v{uv��s������n==�yg�ŗ�r�bX�Q�m����T�1FQ��s֌h�4F��|s����(��}�Q�X�4�Q��~�m*e0!�^���wnI76��24r��PcƂ8�o}�^f�[����ˢ�A����m���m�sԋkQ�l/��[ߝ}�O����8�6���i��kM͍�Z��1����F(�F��~��Ɣj0"d`M鿇��l��������dh#�o�ݠ��!���sԋx��<gG�I	��m��ك{3�c==��&�05M(�6򽲆�1��D���Z1�� ����{�����g7�WlCi[Q���A��V����CZ�ލj���dh�z�A�Ƃ1�}�r��N��}���Y��!��rv�H6�L�0#Q&W~�i�4��Dþ�9F0�1F��9�~2��lq�-��&^��t�]���h��u�L^�3��}KNe
|��vj�cfWX̎�[9XC}l&��;���r��r���QZܓ�I%zf�qjoZ7��t����C��U����6���a-�Om�֧÷7��8�=�\�����[�mx�\�)X;%ΓіE�(=ɭ�hu�5�t��m�C�e��=���S�5⽲X�h�m�3�izk��E�(h��j{��Sr;!Ź�'\�d壜NW�iݢ��E�s�:������n �$qC�h�*?��F���j��������5H����r����&�s'I�/s�*����Ы��K�h�7kC����p�7��?�1���CE1�#E^wԋi`�`A��������o�=7��ͳ����mG�{h(*r�"�����A׊�����Cq����FX��gܣ���J5�}\y���%��^���L#a(�{�h�!���{����iA����}���oS�qmɯm�}���2h�m�i��lChʯ���x�D8�6=�r�bA��G�]�k==U��k�g����s��cXҌC`w��(��"֭>�}����$�|����C���+��$R���o>M��F!�U�r�k���#{�s�c�h#�����/�J��j�oM���} �G9�~�cƂ8Ptχ�9��m���{3�c10#Q4�Q�����[a	�u���gELCh��޴cF4F�4F(Ͻ�eŌ#J5Pj>���i��{�^�ת��ѷ�s��� ͹vU�<��F�u��]��g��Ҳ��WDu�����í�B�~M����s(1�A� }�e�D��Cp�ԃL�e�ye������z��F5�(�Q�w�ܣ`�!⯚���p�6ozv�h��������?�{5p��x�U�cj��x�wá&P��|6s�雙�R�C�z��pN��h�|�a�ʵ6�c�|�>b���6��t^�������aS�H<4s��)�������w=�c��A��_��LC��T}[��z�W���[����Esz�lzof�4�e�__=�1�0#Q(�Q�W�SKl"b� �5�}/y��}�g���y4F�&��s��Q�X�F��(�}��L��t;֙wm�{t[F�U��֊;�����h48�@���-�yG�8}�� �)����}�#�����eog�8g�u�J0������a�h��ף�ڎloz��-h��L�6��#E}�}F5�,����h�q|�6��z�`u���1�g���A("4W;��S�޼]�|��aJ��ZH�1��,�7&�y�l�F�l�ȝ�8���O������8'��<��y�.��1���F�j(�s�Ҧ!���4B��}h�!�w���>��z�Ȧ-3�s�Q�X0�CiD�o��ҦSyZ^��M�ǧ�j��6�}���T}�y��h��W��h�Db�p��R��dC5\ﾤcX(�6}�׫��������y��É�4C�yɩ�6CD٭�Z1�#}���S��Y��"؆��F��}�o{:w��eS۴�������#�"f�b�:b�;κl�c��Q�֑���#�c�i���=�k��h�{}+�2s�L�N۫N�Sӛq��w��rW�HO}��0:21�m�=�PCb��~��#4�Ӣ�7$����oZ-`{�̢�<}˿N}]����|�6�ҍ�+e*b�+���6�M��s�F1U{z�]������5Q5��iS)�q#�D!N��h�����~v{ �񠃌DRϳ�E��q\�Ǡh#�W�A�P���5W��ԌkJ5Q��粋bFs�x�6!^�jOV�������d9�Tq�^'g�퉻ljX��Yh�_5����@�M�-?|�G�#u�l(h�(�F(#E}߾����C`Ow=�1��#AF�v����+z��{��n7��h6�6!�W�z���:c�}���{���bʿv�f�6�W�0g�x���7�a�(�1F�^�zьChƈ���F1cҍF�͕]��9��o\_73����G��ug�Td,��I`�ѿz�H��� �w�[��#�|j�=I�|����l���Cj2��z��CkQ�a��F0��!�yɩ�l��٭�Z1��߯.�4��>�k��{;�oȌCb�F��{�`5�(�bv��Y�Ch1ƂP y�������ƈT�hs?^c[�2��P�g-��X�U�\S��:���v)�+ORÝ���n0���ft�|6�����V��r�Y��W�H<!�����1��G͹6=7�Sz-e�^�~�1���ҌCo��Ԃ�k�_{ܟ<��S1F����Z1�����ﳼ��aPj4�j7���+L����{5)�K>�W�����ѓ�mq�0Qk�ڌOXݶ�݋�Z^J��-,�	j����G�v�A8����ɿ�j��"؆�6ye�?A���}��߷�,�� �uK�]����9�b1�Q�l"a�gyF1�K]�d�m���or������g�AcE1A�b��ݖOn�}ϟ��;���>kQ5��;��,�&F��C}��R�!���^�;Kz5^���g��G���8�>��=kR�ٵh1���fv�bX�Q�oҾ� �b� 1F���U����uh����>�w�c�X5Pj>���+e0!y���7�i�k[֬lCh�v����������������"�w>��ADb�گv�m�0#"���sԌk�Y�g��_���+kCJ0��7�z�a�h�S���Cd5�krэ�ee��[�����4�3�����N�u[�����c���������E��F<h#`����gsax��K�E�vb�Fn�csZS�I�Y�C��S�])��� �r�]Rj�yk�06B"Ȣ+�;�ݠ��1]>SFs˰��R��P^+i�jep
�6"�.��*Fv�N�����ZWg�2'��۳3�õ�G�:ܚ����ucy��ެ�&�F�x�;�| ���ٰ-�Wd�""��C	�1ki-�����қ�r߃���OG}k6����:Q'eK�i�*��R+��}/�ɏ*�\�xRi��U���\�$�N��V�]v��f�C�/����^m�I�GSi�|��ɗZb��j]��X1*��V�A|��8n�qUb�]!���ٽ\�"�wO��^��w\h��n�MYET��T
�ai�71�,�;�u\�x�r:�ۤũ�[��Q�ъv�]�ʔ"버�2�l�H����� �Y��c�˒e� �X��0��F�5˹�.��
v����i���fB�k�6����8�y�J�� �u�}k̠�-���:㙈���+;yr�gJ�s�gH]�Lf��N�@�naw�i@�H/u��C*�|�O�c�9�:�Ph�b��yXGu���fY�*}>̰���>�����H�&n�5�O ��# �D�K��WY�'p���ۃ@nH/��U������p�r��Bo�έ�P7���X4����oK{/)�ۄT�9��|�Խ �9OKYӏ�.���F���/z��RA�����R��YroR�JŘș�e
�f;��V�)S�I[���T��
p�}�GPM�É+�~5���\��]���{h�K�.:RN��pu�rq�ڶ�trtD�p�Gq9$Q%���Gq�ӎ�9ʟ7_=j$����+7>2(����i�B�NT�D|ZT'�q9Nr�tA�A�q�O0q�|Y�A���N��8���;��3�(䯛p�q]��;:Ȏ98�:K����.$�⒃���;�9�	ɷaY��IP�)P��d\E�ܙ�����2�(N��s�lۨ�9����:;��Ol^�hQ��q�[�8�I�qJ��;��B)8��.*!':�)� �8"��B6�Q'�Q؜v��o��{�vL:�wh�*�
�t`�mY�ݤ��\�8��vҹ+��8�j�nt�ؗI��ó�eD��e�d펫��t]m�]���랍cR��ǁ�Y���x�[�ܛc[Ip���ێ�ɝ���;o[ٽ�rgۯM�'�p;Z�[����+��ݹ�%L07�S�놛��/'n狛��wO3�vs-:���=�U����W����th�i���A�����ី��8K'�2{>���v�'�N�a:�m�0���u��!+]�N��}�S��<'��|�V�Wa׃=���l�"n��^9�gG.�[�v�K���ܹ��l�����bx�Bm�5����ѷ\��ֻ4N��&��AKV*�Z�i���z;d�@�"�<�n����=��{;���Z��BS.�c�����{pms�m�@�dP��(�r��F�m���Pq::GC6Cnc9Ǯ��6���<s�^���m��͉��f�����k�.���\N�l��Yq��ۍ�뵚!�;g��v�{C�rJf.�|����]�w<&v�pr7޷f1��A�`�v��@%@,m�JvV��6콱�z�ڮ����<�<GO!�-��1�����ɍ���xQz:��^�&���^r�c���c����� ���/tq۱�*Od�hawnC�pV�Gg��nܬ���xkGi�:b����ۜ�[�u=��u�;W×��]�]����.�7:�Isz�網c/�%]Dj��읬��2G\+��;s�ū�������n̽+��b�mxy�n��X�n�t��bE�@X˺zb(9��$9�N�����\K���8:C���׆n�P�֮�{\U�Gf�a�m�r��;;�E������n��+�Y�=�ۃ�1��ֻ���lnK��l'g����w'��L�3���`�.]��y��<�˭�c�)�L�x�Gr�K'��W�[uXxqJ��n���X�uSE����{���:���U��L�۟g�/��ό �W���gg���!�tn^n��gײ���R:�g��ɏ=�F��]�f.n�m���H�t�@�6ݹ��[y��v{ruǮu��8-�v���V@�th��2�t�B��u�q��s�;6En�+磓khԌ;�9-�&�ݚ��TA�K�`;a����p�`�g�n-�]A�v��5;��,s׫f\���)�ָ�8G�b���nN�2��/���~�u��B�O�����}�c1��(�M(�+ޢ�J���6�_+��cF&���c�~}��[�q1t��v�b�0�CiD�J�i+L�o���s�͏M�ܳ�9W��0x�D����׿���ȩ��>�W��!��Aگv�m������W=HưiF�J0�/o\�������%�F2N���or��!���h<4Sa��}���X�6d`f<��ѿo���ڢs*��`c#Ah"}����9HD_+�R1�o�q��Zԃ5�mZf^���c9��s�����1�mu�J��m*aa�D��޴cF�4F(���e�yW�r��Ϸ�z�^<���iA��*�S_=
�nܚrk[֬lL��s(0x�G� ���^A�������>t4�z�]��-0#ډ��wԌkQ�(���̢�`�>�N;��o����w��Y��m�I���v���u�S�/mˮ��uٞ�Z�0l���~��q��GJ�c���[G�#�V]�E1F�#E�>�5�C`FF��̳�ݿ������;��[A����}H,*r������1�owR�ǹ&�h٩���7�}t[>L�Q�W���/Hv|��N�'���h��`>=L=닃̱9u��6�tS���6�V�I��b�d'/r��ȢWÓC���������̭h����z�������{>�a�b�Ch�����hƈ���~��e�6�F�ڳ��Y{�늟�}T����.}�����1�����z�4�""@=�y�^AAƂ=ξ���k���U_ �80#�/~��&�j(�ﻙE���������ַ�h�E���ޠ�.K�o׻��>#lQ�b�a.�yF5�(��C`C��e������Ƃ'�ԃXo������W�=�D�G7�}HǃA�s�kZ�����A��/r��1�0#Q��߾��m+a���:��jWw�����6���cF4F���Ͻ��1��4��iD�o��RV�lׯ}���M>G�vzo[����`��6b�vB�s�x[�N��^{g ;ۦ��������d���M��4?����E�8�6=��/"EG�8N�=h)�����9��g<�}��Ϸ����cJ5Ҍw��[�3��&�ٸޣޞ��э�e]�[L#^{�{��w&hϹ~��cJ&��}��-����lCo��R.qA��_��w�s�_�I�}�Wԏ�4Õs������٩���ث���c0`F!��o��Qm+a�1F��J�5�={��z��#��s(�L�>�u;�q�� )�wY鷌�	�K��d6ln��%�=z1�|�����w�rϫ������_ߑ�!�|��>�^�1�m,j4��}�~�V2��A�nM}G!��-��#G/���w��y����h4�@5��h� �"84�޾�e�#"`F�/~�Ԍi�n��}�{�=,��Hmr��I[H��M�M�5�=��*�waM!� ��}E�#�ݹ�p»�}����#{�v�``��G8����Z�!�"H��s�F<�����^)�����mK �(�DcgI��t��1����ٖQ�ZGa"uE ��]���$�Vאc<�����c0`F!�����M+b�"�W>�cF�;ɟ�}X��q����F1baQ�҃Q���he�!y�W��oroZ�77c`Zdh����4q��:�rps+�_H"H"8�G9�v�[,`FA�/�ϩ�4�PiF��_����_�}�.4����͛�������m4G��
b�+���|�4�j0 ���p���{/��&F!�q����]�AE���#4���ɢ޵��٩����{�e�T��ڙ�m|ҍDҏ��l�Ҷ�1�^W~�cF�!�1A��o(�>�����Y�{{�F/�n��K�t�TK�_�C�W�<�{6�o<\Y�/!�Ո2e�(��V+���?>Wσ�h���$��-��j1��z�So�du5?3Q�or�bF~�e"؆�6�}WE� ��S��kEg;]}o�p��e��!����_�ݤcX4�PQ�a�v�a�C�s�5���k9�?��8կ�a�%�Za���]�w>G�XY%�ҁ\v7����ˏ��L��f���yh�Dn��R
b��!�h��v�Ɣj0##w޼���x�}�m��y����pD�E��#4�A�tֵ&�{[V��W���c10#PiF�����oܫ��V�6!�K�}��1�4F����yE�����ܹu����]u���z��/��4�o�����X��m%�4?�̿PcƂ8�B@=��(��#��[>����[�os�}AL����_}H��4�Q4������6�f�E;Ur�!u�ƾM���IeZ��+��3�i�ba�Ѿ{�Q��iF��w��Y�Ch1Ƃ7��ԁװ�p���؇dG7�v���G�yǢ����٩����{�e�`F�J1�g}E���l����=ꮊ�pb�����cF�!�1A�w��c#JF�j7��ԕ��ݝ���+-m�w`^�?��_Y��]A�ͺ�j�n�ˆ�aW�����~e7��MU��\޾I͛��Y�s����V�|�yEs�� ���4�֪S����d6pm/L$�v2�,;�::]�Б������OpoU���^�\���p�m�ϧ�c���\��nwrܖ�{�K��@�q�g�;Vn^	p��n�铵v�V���Ͷ#,�v��Sʹ����U�+����#�9��3��kq�/=�۱�8Վ�Zb8�y�S��Ӈ���3P�\a�Ga}�5e����gu��%nh��qc#q�W��Wʼκ�.1�`�G�h��z?4���M���wt��q��@9��(�PD�h#����2�����>U^���j�_�ϩ�(�iF��z�a�Q�j���1Λlֵ��F�,h��;�A�+C�ݾ�Q|�^��\�1���9H�!�8������c�q�o�>� ���9�WL��_��sA��y�Z�r=��A��+���c�Ɣj!��w�XҦ�1�������~�ԫ���4cDh��3��eŉ�iA�ҍGٟz�m�w���;@�J���K�Y������<��/��b����[�A�h#��{փl�����~�v�mk�ϻ�����.1����_ܣch���v�6�rB��m|��K�|�k�&�0����`�4���^�s����	{������mN>��i�ࠉ"/���1��G�����;�o�g�>>H���bbo�D��
�>��@"28��N �@�N�1�Z*(�UP�O8��:ԕ��޴yg��;�r�f0#ڃJ>L���Ҧ�0�h���mуDh}��k�9�{����|�1�F��C~���+L���c#���H�7�f00dh篼�Ǎq��=es`��=�R�%�ͳ�R�mevJ��-�s-fǊ�����5:af�`�4��j}�EEf�=F�
���>���H K�|�z���� ��7u�Z��������#Ɣj!�e�;�gs����竹GXq1F�k{}r6���k[ܴi��#����Sأ�y��"؆�6����s*ʞ��:[��q������ ���$Q�gi�h#�A�}�ֵ&�{[V������������>VW��Ƹ4�Q��_��[a(��y�F4cDh��1F{}�(�-���z��w���1�CQ�����%l�3�E�u�`U!K���4?�������1�"�z��QyO�g8����������-�����}H�!��J0=]�(�!�s���zkîn��`ә��Y(���iUAk�Sˋf�m�qv�L�����Dn���s�}�X۵���֏&��*���E1@a�a/���15�(�`A���ﾢ���?��镮}�|��?M�i�9I}��R1����<9�d��pٽ�E�l��｜���6��sټ�z����{�A��A�4K�~�э�"h�Pgk���bK�.OO}��{}�+��OS�]%є����1��y���۳��y�O8�I y?<��H|G��R�Z�{�wS"��Q�i����iI~�2�Ylm�{�7]x�^�����b�����@�X�����'*��:����|>��? �?0#ڌ��w�F1�Q�z���c�DZ��	rumMk{��1��=A��fn�<}�6��b�#F_��5�C`A��>���1�m'8�>�Rw��{�߻��tC�!���HǍp�v��z�ޣokj�c1������4�Q��s�XҦOw��=\���6�}��э4F�4F(���F1ba�ҍG��z���`ogط[}�9�S�ӭ�;�6g��Z���k3���\��k�[uY[Eڇ�UA����ҹl
���ɴ����߹A�Ƃ1@>���^AAƂ8w_g��l��Wޟf���tk����R1�iF�Ҍ ���r�a��4J=�9��6����=�1�D~�WAm�F.��Y7m�����·>���E���`D������c8�A���z�m�wM��=;{�V����ԏ>�p�9�f���6noE�l��߻|���6!�Nߩ�u�1��̱�ǽ�f���#�уD`}]�(�,F�j4�j>��ԕ�)�5��m��u���۳���w��w��o����ݝ���҈�$��y�xA("84ϵv�m����#?<�q�K�Uv.���J��T�{|&V�pl�(1�ope�m�"�[���m:`�d��^h8niɽB����cm�[|`Bom�/j�E}� �%�!���g���c�DZߪ6��ښ��-h���g���LQ0�PF��w�bkY��+o~�euq�c#����؆�`��e�Ԃ�r�"���C{�_�OS�Y��ﲻ�>�u��ΐ"��zq\�ݮӹ�v���x�7�����UG߱��J�n�~��]k�J���1�mbiF�J>��h�Ҧ!��Q�+�;�F4cDh����˴m���s9F1`0�(5Pj>ϳԕ���>����[��wi,M�s=�1�Ϻ���ϻWu�\�@�}}��"B�$�G��v�m�����e�����`ҌCa��q˜��}����(�G8ru�O{z֞�уD~�WAm�F!�_���15�(Fd`C]�g��z�E������F!��w=H.��"Ey��HǍs�����zn77��6X��|���!3=���鿀�V4�Q��ՔXҦ!��_=�֌bر����1���o����p4Ҥ�iA��9ۤ`^�c����I��f00dh���)�`� ���/ ���/���ˬ�o����G3^�Z��d`F�/����`ҍ@iFa�_��e
�����t������������Yu]�B%G*�7��l�%J㋜�`����:��nה���F�M���%6gb��SA���t\6��ڮ?��}���c|O�2K�ލj=K�ػu�=�wl��2[��vص�HD��^�j��U[����[Glx7���Y�g.��:mc̑�aۻ[_!�Uخ���ȝ���l6m8��i��(�i���z����ݼ��8@��F��=�q�&wZ-���+��۴k�v��][a�u�֦ݸ�.[e�P�d����ٺ�W�]����)���nB��a�{��C�E����K��u�'�맘�^8�K#�%�N3qѤ�^6�����~�뗯5G�{��4Gs9�h�(�1A�h�s�Q�X҃Q�l	�_����_2��x����}�T����6�=�]��/=Ϡ�@g��/��t+�#�#km-m���ς���^����5t�����N_w���oT���I]ZsZ�1ck��s��7ֶ�B�tx�o��s��_���bu{k9��I)�I�]j&t�sw! �70h'�����?�ن��,��Qw�x�7�]�1��������*��F� ><��g��hKO�J�[nn�'��N��	?Ol���˔�B�Y�I��e���=�[-��Mqb����X:��]���Wnֱ�X���{m�7ϼ��
���o��b{�L
��w�eh�
Yy.W�ܹ���f�٥�1��ETvXI�{���q�4���Ug����U�3jg-ۛ������7�w@�l�ŒK��]z�,m�xj��q�8�ϲ����$���2����|�?� �s7wty>{��m�3�\��{XO��r����H�����j͒,Y#t�s���I{,`=��딖o$��? w�#`�ϗ�R{�a^]��]��_�q:�e����� ��S�( ({_bེҾ��z?8:�9-o�+��tr��yY�������Ϳ\d�Z�O�y������֟�f���.x�5�O�;�����Ϫ�y8�v�W*g�jt��ڮ����-�5����>�~o�(�2������S��
�[xjW<�_VU���7A ��g�E�A /�,����zt1B��U��ƕ��7'�H'��Հ��x�~�:��:ky�]������؀|����4����?���I%
2s��x�"Ueb�b�Q�8�-��炦�������G��q�q��[�xN��@����	/�v����Xz��"�w��d)�y�����V	�ҮWO��嵨KK�Ծ$��}v��ǘ���+V��Rבյ��9���Xy���K��]��p����n��"��uɐ�b��i�R5���wV+.�:ذ�2���*���v����gs�'CNM�K� W^�k���1��w��O��Ւ^�!����%QG'^=���E��Z�<����bg�L#"F�b��m��
���m�t3
�p,��QJ�q�_�9����-��iu=��U�g��k33��F����5q��S�&�A�˵*Tŉɡ�쉆iu�ݕ��Ov�K���9}cd7�cW�����9��|��b<4I��oe�ط���z-����l^!9��Z5jϡÔe���e���1ڲ5��,ǉ����\�������"]]1R�+ۙ�%�8�z,�(���W�x'}���3�+�8���"bt��o�c��4�m�}��ԭ�z�yJ(&�`5�#�XC�k>��N�J�B�4%�v��M��qeDr��;�B����O`3\M�n�t,\��4�������t�d�Lf�w�W�~�����\7�}j�A�V�*�Z�9����ES�6a(f�7Nk{�D�@��Y����:��*�V3�]a�w=��_N�%BHdk�>e���7|�&��� �M�6�1��YptA�	�S�'%�9wE!qw��v�헅���Q r!�AE�t�R�em������p �3;�ó��.#���"H ��m�E�ͻ(��.��8���@�8R��;��#�{Y�9�e�o{]��Ok:mݗq@�A�b�(�)�J9��N��\�ͳ˵�g�yfX��ywe�#��us�B�@UG'I!DuY�NIf�D�ΜpD�VZr�y�De�VYp�p��DEJ^���(r��;����;����n�򳂓�:�phm��ƛ$���H7�̿i�����T�mk�9��ڿz�;BGYP�)�^S[Z�ӳN���8����� >^���{�^�B���R�z@�W�f/�q�#�]�"���T-.�O��]�:G������P�6:^���=��~�����1`yz�d���	vԝ�#��M���3�h����d����lSf�����O�
���uc<w{�~$~}�I3ˢt�>7�X�(S����{��AѳR:�tn��{�����֧�ڼ���Ύ���k�.
���GK�f���$�s�T���=<�t�_����Q��I}�x$����$G����Wj�uGe����}�}��t��_Ěo��$��ǺH$���Ν�]��3�i�'A-E#�̬�:�*��'���8������Ùf�rD�2����f���s�+#YYP�����������A������z_l�~�M��0�M?ϛ���inQď�xg6o��4���{��H�݃����p�w|�}����V�s�젥�kf0��ky;<8���G%���
�q8�����T���7ۤ�^�y��H�c�^G��Cv{��O��O=�	�ɺ%X�jŪ��y^p�������,���H'�k��o������r��;7��0舅�c0ҝ���Aދ��mf�e�=�_{���F������]��z����[緛Qe1Ms�����{��`W�^>�� 	���4m,�4�5����bD[����M��*
N�Hz�;�Eʝ���Oâm ����׀2M?o�HK>l^N}K���8U�����K�P�׸J{3�.
u�K%.�h��#3O:�tiǖ�2�P����Idլ�e~�|��|b��D��;c�X�c���r��x8�uOn�Id�٦Cs(�r�I���uۃ�N������ٸ��s>dM�d�ccl�[�Jx�3���yw]�ۭ��8��Z78��t��lt�|�\q����Rۋ��ɸ��0��WWkmv�v�[c��c۱��= Ar�mN��:���ػg8ء�lc����S�vNyM�C����$1P�'N��2H�4�7dwZ0sڙ8v�3ǟ\�J��J[(Y�F(	�m��ެ"������Y�s1` >�﹚>@$��?N�	d�gY(`�Jd�z?����X1 �>﹟h3|5�;%��F�2�7�F%Q&�~z��}ԯl��?kN�<d�%�}̀*��_%+�y��N>�7c���U3��y�3��6! j�^dd���vV0�g� !$�󛸉(������{��b�&�0�{�cO�xCK���H�Jc�����I5F�z7ᒋ��D�8;�t���|("I�c{Ѿ�潽b�D�=�����{2���$$�I��y�ٿK��������7uv��e�$OZ����{��=�9�}gv���`� �Q����#�
U)hnx1����%�[��xrI @�on}�.?��m����������ƫ9��*�n�V�C��wR�&=t��G��Ԇ�����d�gt7J� ��;V��}]��l/�s}Ok�;Y���7�n�|i�������3X�U�$�g)�/�RHI署 ���8� ������ \ɴ����`�\zsZ糛 >�kz�	 d�\��S'�2Mi�gH��^�޴�U깵�Z�f`y�[j��R��9H$���u$@����$�9/���̄�;��L�I��g����'0�A����d���w�^���L{��bB_�����$!߻0�I(q�3�Fgss����D)�$�v�E8u��v�4��N�ڬ+�+�!	�D�eh�>|IB}䒵F�>�?M}ܗ�=s�@ԂD���oR��J�1�7��'w$�A�o3L]�d�J�-�������e�xz8�9zV7��^{	�$�Z�v�:�P���"L���W�^���(�g}BG\R�M?<�5_>������&�Ym��7)2熕d�;H_�DTe�g�N���'E��Vάѝ�_@黲����l>�F����q�s;Ψ�Y�Q(6���r~ �{���䁰����}��/��g�����Y��	�oމ}�� �ω4J�N�D�MC��I4����K�z��@#�]�b�W"�ԮrTJ��]��|���������k��$׌Q�$�e�NyǺI��+4Y�A�S�*m�-������<%8�<�]B�����:�c�P�qlk���-`ܦ��E~�fh>�0y������_��ID�=M�N��Ȁ	�ϛDҬ߈�Ȓp������B�2����&��D�'�L<��D�osr��2J��}a{;ԉ��t�ʥ%L~�f�߻��D�Q�Nsy�Y�6� �h��w3Cg���{@}��G;Y#���*ۣ��L̯j���D�ps�ѢI'��$$�<����O�*!{-ee׀̗�	����v�b� [�+�t)q߈;�.{�3SW�bK7:7Z]c��mW�6���)g?Q�'P����/_MQ�B@������]� _{=l޴�t�,C��3�w����bZ<�4�Uc:,�j���HH���msI��l����|����(Ǧ;
K��W^���,�e,p���T*�L�6�$�:� E�L_��~v�A�Q*��{��4؃=��6�6���hoT�Զ��h�k��h����rY�Ȅ�ت�I#V��OُQ<��λ����M$�iｲJ$�~4��� �=��k�V{�ﰜ���O�I9wXtgOI* ������ h�}�u��g����Oğ���HI$�P��Š�]���)*)(�b��o'G�-��O<I�&r�؟ICz,�$�;��S�#֛�L�쓻�K���UQ�b��+c�1 A/d��mff�/���	��Ě׻�J$P�G�2O�ym��)����e�����M�"��^�F���t�%&�n��T�=3��U�$�{��&V\L�퀸��NT�������Wp�濋���|EV�pۮ�<9�k�v弘o*%�;n;�W�s��S����'^�����Ϙ%DIx�n��ݢ�;v)ݞݹr�cFcRq�炎���o�����c���ȋ�q���N�ὣg������+<y�f�_k>��xr�v��mՎJF���mMB�x`�vr�Q��4�B�p���۬;]��=�����Y9|��n�M��[�k�s�[��S[/ggۍ�]ey�d�5FI�I�qt��{���:H�J"�<�"����� ��I�Oܷ<����S�}���v�9Ν��K���Ĭz�3v)R*�ʶ�EqӰ=ǝ�jfE5�Q&��G���$��� 2w�Rz�םx���lŪ�+ �Ǉs3���W�jD�e�^b�������<� �@i����ClH�r{1B�顱g�ˬ:3Ӥ�Jt��]��� ��XĚ$���Y$�O��b�si�� >��^}k��F����Ɂs���?Q&�sݮ}`=�}����I�/��$�$��� 2O���$'{��o��"�i;�*m;,j"�_��ݓ=k�4r�k��kd�B���EUI�����P��E�W�|��$�<����~�I%
�2"���^�Q�ǭ�	"=�Nɧ4���v0��.�n�?n�!6���V./9��l.K�ח5ʽ[��:͉��l��n�D�!ǳOՋ�z��$:I��3�!+u�IĠ/�C�i�b=��\��U~I	.L�s��n@���׼� ?�}$$�~C2����wv��ly�\�~�P����fvo5��s;�9$�\k�fJo��y�ׂK��^�b�=��f�Om���U%bd���>lN��d59aR�$��}��$9�`J$����}q�<Oq�$�|f������$�600��)�Bw�sQռ�V��z�� {\�w$�I+���Cƛ=�MP�3�IJ1��z7��`���5����ɝ#ϋv�'%u�ȁ!{���O��*,��F�����DI%��l ��+炳N���}mn�\=���,�{��{Vh]s��HR*��9���9�J�0�#�����v����g=���/�fg�`{��SF���C۾+��'��}��v0��.�n���7���/f������d�������X�ډ%������7�#�>sp!o;#CC욈|3s��s}�g�N�#+�EW{C����9r��Y�Y���.����~���0��7�ۼ��^�|�P����c~yqkY{3����$�����Y����$�|��}���OO�/����Nl�ک+/1d>m�I'B�6�����-�xy^\�A���f�^��6�u��Ѽ�ë���ݯ|m�~���&�O��KY�a�:��l� ��WUE%�Uʠ�%R�O�]���Y{o�y��� �sYF���|���{x���)n>����&��m��!>�E����=�سB��eJ��z���Ò	$������$�9<� �2z>�e���I(���
�f]�EF�bF?g2�@���K4| e֖n+����$�_+/ۺ1>Dp^��E�>�V]��9tr��9�z#��Z�������>��츀��6_7=�C�K�f�����V1S��q测�؁��X��NX�jN�g�\��p7�Xrs�Ns��^��X&W(�K>���_MIy׾�*B���z�Yl$s3����>�y�\�ml=r���׌�I<��D�O��}#a�'���wZ�����#�Q�>�7�.��ێY�s�u��ڗq��''^�gT�������RV(Kx�q������{W3�|�${�.�>��O��c&�� ��f��hC�ZdU�{���v�m-qh�L�����U�� ��� *~^�%���<�h���k�w�*��P3�2�d���Μ�� �{��� 4-�=���u�+�gc~ �M�2�������`X��>�cE,j������U��{ޥ�Ǹ�p��e ս$��i�K�ͳY~J!�I6�o1PY����(�A�s[�g66��X��g��{B#�]~�j;d�$��o�U~7�ͼ7_?��{gy�vZ��w�5���;�`L�X�br�F�;H*U�.��0��57d.�NẨ���h˰�3�R�P�/��U�3:��ۊ-<��;k�P��滏7�WL��vƫcm*��1V=YX�&�;{���S�����<b<x|��s����=S��75�o�m:�,�n�?�ʣYZ�����M>̺��cqh������%\=N���]�yx��nlt�$m� 6�ެ}2��2�2�+%�>�a׋ik�at�Qܭ3��!�8�^'/O��8{�5��}e�qtZV�y�1���w7u�X�]z&ܺ��v�\�jݽ����`��vs���5Z;�w�����u�Ḻx���w��j��K�bW�pǬU���t�&���뷐J� J�:ܝ���V���3�o`�P!�]�8^U��,�����U]Ԓ��	��[+:m.��+���|'c�`�H�C���O�0�.�Y�ɢ$�M4+f��/p���k���ᣨS�G�/�u>w���e���Dn	�{6�s&���@�M*�ܽ�=4�:��#�a����	s��[��k��b��4l�$d#-��0:���u�%�muh�%�I���U��b�Wd�݊DڣQܓ�]Cxp����P��O�Vp�cՙ�Ղ��EP��K���r�m��e�s�5X��(����Y��y�q^+�2��;
(u���CČ�Z���e��q�!>�,^��+q2�k�Шޥs�����i�fιG>�-�O�n�oT�����!�pm��8�裢����.<�ɶ=��[iD�D�tN�g$GP����y�㢎����#��g$^vvچց"pyXy�8DM�N��ӄ�	!y�(�JD�8�R'�'���O-\#�2�g�PB=�
rJ���I�E'��`f�Mj@�'a� El��4:H� 	<�ݷi�;0\��+;V��"�u��(�0���s�NciPs�Vu�Nt�J�քy�GIg��9#�;�.$#��#�p���8�Vd�����}�(x�Qh�z+��k6�;�����D]�����mۖ7k��h�q�i����g�{v�tl�l����۷mыv���㗆l�=�[.+���5zL+7'eݸ��nHSv�v����e��v3�;=Zm�qGZ�n�u.������\�=��ہ��=�x���p�Y��.�=��ѯ.^�`�+�;q��g��\�bl���8���1�q�C��Ǝ��ҟ�ַ�=��t�/[���Lj�
v
��{=ˮ��<��2m�۵և�Ꮋv�{[����L����C���m	�$�[]0�s��r��R즧�z{#������8b�\@4�����&t�=s�Sr�x�M��=T�i罍Q��S6�;��/
�[h�q�8 Ļ�`�(��	�Y��|�����˾t���e�ի6�g�n�2���8�|���nݙ�N	�p
�X�'G���=g��S7=���糱��s���o�8�e41��s��\u�U.q[�h�1�e��a�ul��=�y�7/�(0N]�n�K�ON�v��I��ɓ؃pr��Z⩓u�_v�]��(j�'sۍ��mds�׳�4P�!�d-����{EMn;N��>�m��덝ˌ�܎ۈf1�ه`��+��ػc4p]rv��0l��y�˺�7V����&ݷl��֓ux:�mLr>�ܯc<��"����.�퇶�/{�s읝��j�n��;8uqs�dM�sj����ձ�{E���v�q��'������u�7lq��{bۈ�\^�kf�v�ڈ�e$c�)���c�s�{8�b;wMzpk����=ن�e���΁�I=�Bj[v�v�n����y��/5v�����l��d�]�.�n���A;��.6I㔥��I���sf0��۞��<�V�rz嫋�l�^�=�9�j����+���ՏrAp�{������[C�B�ɝƸ�t{��f��D�i[]n�p��;$���|�ѰZ;cZx�9h��2ss��ݑ��LH�6&�;��/]'�;��nR�ri��`�,�o����ө:�q�u�t�2۞���R�#��5�����ۧ�km$=�+���8݂W�힓��;Yn\>x���:ݎܯN��a�'�k�fq�Q�r�gpki��=�!۶��1�o;���v�6qܮ�좮�çvA�D�7n'�v۟�\r%z��۱Q��xș�ї	��n�M��������Ռ��,�\5jM\�m�.{d�wih
�֝����8"��$s_ϐw�}�s^�o����V�1��5��=����/��a����RU,�)e���oz��e�Թ�[t�3��I�ž�|I��Tw����N�g=��_v�52��	t@D��:3��J�I V�l�I���0ftɞ��W�H$��ӻ�%�s����w�cvJ�LA���Y��|�v����;�f�� |��5� �ظ���0�;=YP`��$�I�k�9�F8:�j���3���]�]����}�$���wp	$�P�ݲ��;���$�~����[�6IS���G<�Vs.9M�"q��:�<��N���/��{}�yY��J��w7�� ���Y'R@OG�u*�)Uoz�
R�=��	 y�Y��K^ug%�Ȭ�I�	{{o	%�ҽ�?42�]����qR��U$�B.����S�lxn����5�y�^)ם5!��Y���,����������8���Ama�F��Dqv�_� ;���.߉"����ڒI	��ۘ	�r�Zs���s}́�$��\R�t==�z�� ���\� 4���V�ݩ6?v�I>ʹA��G��@%ʰlx54��*��7�w�&��Λ�%�x���@ ��c��g����r�_�-��I${wF$4Y�M�;S�Udϐf�� �o\�oe�ꐮ�4�|qǌ�TI��{��~$�-�%Q)�'�K>�F����Be���n������)�.��{=�/��nL���$��(:�j�<���Z��l�@/�zID�׎�X�y��VL��H��bN��@�&��7����OIP��p%8R)��溙 ���I4�����%��2��+쾥���ŝ�'"�RH�b����H�k�ʄ�I&d8��(�1�U�zmT���,�,��Y�<Eʒ����콧#�?x�S�R����-P��T���M���0˧��.���}'�ǀ����n5ĒMߟ�` �������+Ẽ7��ӝ��X�h w�Ϊd�I�����I>$Tk�����O'�{���H�V���O�V���i��HW�����'����J�S  �qo��I$U��2��.��"�$��"�H��l
�d�;n���n��ygq���뮋c*�Dr�߾�u5=V�h���;�� ���9	�Mh{9��'<�q:���s�z���1���\}��4@�o������E}�f� ��%<��V�V�	"�+����RBFs�uw	3L����E�vo7w�s��(�X<�\��������f� �坞�r���~;�m~%��n}D�MQ��m<�:����Y(H���a����������@���Ģ@47�4�?�o׸��n{�����)
|Cww�rYC؁Q ��'r�yf�����$v�����J�	��+A�~��DJ����ahÝ�bWG���?�B�ߟoh����S*vY#�\����s3 	;��.��׳;"���D�V��%�H!靻���Q�^�V�S���=ɳ��`"��Z��
'j��W9YC+:��SeE7��lE���V�qy�b�@Y>�^?M}�rI/��ٺ�I!�o٧B[�_�����Ov�߉4I�^�����:��bj��Y1w����]5�
�n���@����k @#��b|\�nwY�M{���/j?J�$+���+��4� �;s  ��>��Z�L��� ������=sf�{e;d���"�{�׻Ʊ>v_S����hԂD����N��(o�'tb���x�jg����~���� ��;�cd�$���l,
vƉ�m��6�@:$�����A�_��ܢn��ȼVS��K�NZ���r�G/oV�E�3k\Y�;�ybl�rr��1st���,]���R׹W���^��9U���{q�S�z�ֿ%��蝝����T���l^n�جV����zq�N����7-Kl�0���
��tZl�v�m�'�wb�6�u�����;�,s�l�m��U�n�I�[</<u�1�3�)Q���6y�yӎܠZջO\�К�\uϓ�1�WWjy�8�{�n��P);DZ6{k�G�a7%/W��n������pB�ۣ�p��s���<���<�y������+�s��<���ͻ>tn�e�7��ɳ��5�"�+�ר�]���}����M;.�]��F��[������ �/��nQ9�$�νu�߯3��4�[l�I�9����-# ��P�\0߷����Il��W<�Y��2$���0� �y��x%���y��ԅ�lX4��,�����g���߹����E�Bx]��nK�̹� #9��Ϡ���Z������I
���wZ�[ZǞ�޹��l�����{F ��s���'�q��b�=Z��CO�V�=G<{�p�w�`4��/{d��5�:f�}��t�������de�~$Ӟ�I*�?Q"�Ѥ6G�,K��U�~��]#r��;/u�k��[̮���&�$v� q�]�m��b����qI)��?�������o}��ݹ��ʔ��ۗ�k����@gy��{L���H�B�Ԏ�yt[L�}��nG����2FC�3s�d����)�-��Lŧz�[ڶ�����ٱ�=��T�𙘳e�lr��v�cE�eK�>�>q��6�A�v��IߣO�A�j���݇�z�l��K$i�UH��>7��w�� A��7�H$�	x:G}������٘�i��� ��z6�_r�k(���&w��j��>�`2�ͭ�Q5�'�&�'�o�ot�\�5�DG�>�����~��el��U]ƽs���H%��7�Mz��B,΍W��o��| �����;��f({��]�����h'QS�� ڵQ�TN&O�k���ٛ=m���U��G`:��^\�{H�d�Q���'�O�$�[ͤ$��3́����z�ffx ���������$�n�%�}��vI��d�q����D��M� g�_���4M��dM���x�����⊔�V�υ�s��� �w=�m$��q�w�������u~��s��
��}�ONד��i�\5��eM���u�$��g7,�6�.]v�L��Y��.��K峌�ꬂ�| ����$I�<Ѩ���N�۴��FU�C,$�Q�B�|{)�t��2�W��$�E�����3�uD��.Ot�q[��"ҙ�3�O �/{�y�}ŪAOnW\Y1{�ِ 3��{7���ߵ���h���<�$�hΗ���4Iy�w{�	��=s8*��*1�9U��A��[���O;�y�su�!A�.�s�ri�>{���$v�E8�\���̂@$��ܗ���%զ����RIw����[���V��G�0�����lW��/�$����Y{�̚$��/Ȁ���#{�7��$kT���i�kά��rJD�p��;w7�d H3=���6 �qHu����L�-�L�E|��s��V���I'e+V�b��g��~��En�:�	왋!� fs��� 5�k5�{�o=��p�MXt��9���ނ���agnދ�ӴX2���㺽y)n��:w�75��Iqk��={/0=Xҿ��_}��?Uh�.7d�A�>qj�E�\0�ﹽ� ���5�t�.�����>D�s�̲I-�s`O�5F�ɷ�>|׃��� 	�Yf���'ag�{{g�.y��q���*���#SE���{n��VÿOС��7��YͿor@$�I=��H��7P�q��=�'�>� ��=�������H���V�Ƴ�[d;���\�������������3>��7�����g���/����m�q��>3��J�MysH2MQ)ev��z���o_�x�I%�ޒ �^i�ɪu�ِd����0=�M�Ŝ��w���D��w#�}	�Ođ��@2M�~}z�����u�� ��緽���'#�n�(�ɂ�7�� ������z�wI���=���^׳3��w�����=<��B�!򦽲���+Y�*�$�lQ�d��0�fA�tiEc3*���L1;u�Yu%T��(ݫ����]�O}���c�ӕS�q�w����Fe�}F���KJ0��7kv{�����y��a�av�t;sx1�r�˲����l��pn�Lc���lqq����ϛ�{a��G�k�we�:�\���s^���k��ϭ�6���7C��^��vY���[����plV�-v��n��UN�i���z5�爴&8���'��y4���9;(�v8��۷L�y�.眛s��cSz�q��/���7�.�ݺN.�۟`�7Z�B�*�P�J	��~	��@�#�?��o��r_$�=��RI�J�"F%�+�&�]j��o��%M�Ծ���H��� �v{@;����94l�/��B$��6� ���@d�b*�c�ǯ[��������k��{�����C��ݛ4��s���}��D���̃D��t�7e�g��X 呕b���~��SsB �$�Ry�� Mn��.�4I��{���mM���]j;��.湙�r-��2K"v8S'�.7f�$���!�w^�u ʡ<��I$������ ~���$.�W�1w���N��c;��Kx���vO1�:�l6�Ӟ!�)}x"*��P%s����G$N�\v�y ���H$�IͯbВIo�ӻ�e�w<��.����l�D������MkA��@��61�g�������3Ld�)�A�}1���7��U���/4�j��N�8�<�p�̒����Gz�^ea�UH�\���5��mD��;ڠ�2�������W�:�8�� w��I/��Q(�WY9(�W�w,��0q_�(��L1w�ز�7�w7� 736�m��=�'ĒI�w��I~��Bs�\�E����V�����NiIeI��Ν���{��~$��¥6��p���zs2���"��VX�������$�N��9f��v	������<��,�K��ܢM<�uH���{^���is{�j:�*�U���"�l �&����e:Ĭ����br�B�ޖu{���,����ަ�!���{7� �x�$�h�~�7��$�n� ����{1��DH;Z��S��f�|�ܐ)�����C�>f���{ kލ <��K���>9�t���E�R�U�]�s;��� �w���UV�����zz<��i'ؚ�&���Ҁ}�44Ŭr��x�w���Y*�`�U��i��%�+:l��oD���*`[���1�)�v�}���e1jձU�U�ֻ�l$G)��yJ��'B�ņ��;��G�j�9�&S��W^U�����2Pe�ܐ`J����-���>Jᷲ!Pm��B�^��%�l�v���92�Md�af�%�$f���X�RfX̾�ֺ�ɥ��Ե�og��;W��19(��:x>��S�P}O!��Er���M_��:WN�˨�Բ;�㝓^�n.�a2��51p�{�m���=�Us�<���]��FV��#�H3�\%�fG"m�Q���B��Y����˷���f��T*��IҦ��LW�mL"�|\斺��ZH�5Y�]c���M��r�S��w4K�,1-�vQ�w]h=֗`�𳍱lt�j)�b�f���ɜS�u�Bs]'5�u5���)W]>�*HX�)�(��ގ� o�E1>��$�/�ǟkM�j�z��n%g��^kln�ӕd�ʫ��˭�uhw��Ni����g1��D��(��X��:����3ꨭ�=;#{&$޼k��������M�˾�Oe�>��}��;�lg�(�.���X;OTy�.�;���4$]�:�y���Kc��'�	�5+ܺ�2�k�Hd�%�XBH:�kN׳���~��6�6(sjs�,�7!R,�;%�i�ɮM����7V5`��܇5u��m�`N���|���#666���8莎N�#.��m���v\�u�A����S��JYi�\qp9 Ry�NrDyn(q!�$�:�#�㎜���G�㗝���+�Җ�Zm���;8�kYٔwؖh�qv�8�3�"N$��؎6���X�q��@�/+B�;���;L��؇��d�-�s�!΋fpD����3�h�t��e�Z۳�:�3�mFA$�*8���퍬���ۓ��:�&X���NU�I��Υ�β�-��Et�γ#���	f��kGIy��N#��%�Q��Z�i��@�ӃM����o.zF�����I{�ww%�6�mIƞXYd����V*\���D�zzG*D�M��tI$�����QI�- v�������`������Vٯ)��h�<��ӻ#f�)b��D�X�I	4H��i�2 '�ߛ����gq�������},���k�ݴJ+]mp=�Ax&ۮ0�R��E$i���3��|Eh���<q�l��$
�F�S$��'��x�7����o�_w�H �n�ߴz��9"�f����z�盦������Υ�@��5�� >;�OfA���x�������{�ܒoŔ�*����p]�s4���'�d��S3������U���$�Hzn�E|��ב�f�w��Z$�yl3<����K���ge<Y�I$37s���$����I;��;�n���Q�+Ӂ��-��N�⨒ffD�B�r��{��\��<4=���T�+�BVN�n8+7����fg�.6��]}r"�����;�mʲ�%����$���6'f9�ddj��J$�蹧TH���V~$�M�6�nǶ�*���q��`�*!'n��R��[n��8�˶�K�[��푈����������X����e��������s+bD��������RY$
�5����?t�s��^x�4Ո��b.g}�{�%�s�ƍ�1���R	 ���ք�K��s��H%|o�RP���>բP���X+!&����b������H%���lN�L�%��6�۶�+��I(���hسf���31c����~�����Q8<㦉&�;7z@%~�^�]�]�F�!&�(f��U�\�H���<G��w{[ �kz�"������<﷫� ��s��� �Q�sF�^��o֑ ��|_�">V�\ʚօd��QϪ&�x��K	E�3x���e�*�U��`�kV9VJ����ϙ��}�-GuZ���M�E|@���ݎ���V��L��4=D9GX�"��w/��E;N�g�s��*�̝�wc.���8%��llv��;�C[n�A�|a�oA��ۛ��K�Q���e��Kۗk۝�"��ۃZ��n�æ�X�d�����2n�.�`x�m�w>��G;=��$O7On9T��6v�K1�������esF�Ʀ2�nN,/]˥�v��[v��+�{z���-�1����T.yz�>������8�6~H1��ϖi���{8r_$�I|}~���#����=7��_�[��Cl]߹�� ��ꨎK3+���փ&���7�O�Y(�OOos6�@!O{y��+��).����#��=�Ϲ}�(�V"��X��f> mN{zİ �ĝ��7�3f�˴�H3}�s6 S��b�ם[�1�d$l������I3���'�I$_z4�?O�{�e��%�z�Mc��BO���Fś6/>���:kh���N��mi�Wk]���D�[�$�����vo؊�#�f��Ã|ܬm�o���;�]q����.�cs�6���;��Q'Q�)'"�"֝h�ן}�S�KN�#��;�������x�@t���>{uD���7�]�ft�D~�fh��5��tr�1 ��{3B朋��7�y��~i�,�θw��̶���w�S�]4�%8mMD�\6���N<��/����K=#������3��3�a� }w2���oٚ�x�C��Ac�G�5,�f��b�/2������D�t��@%y#��ǥt�ߕ�}�A$���H���o}=�ȣMX��f;�o�g%װ�d�����D�I>;9���l��߻�����J\n=ы����B��ZtO����~�́E�:��F����$��o&�&�O6�4I^��!6٢W�uk�Z=$�p!GD��qy��v3��l5<�.3��yY���Gj�������^���캾H������||߱,�b�zo�����kiDI��gj�A�G��MN�s�V.�Q'0����@�7K2�%��I5\zy�$�_��I�$�{�s�J�d�*��ω�.�b����Y��f��f6��ܲL�u=N�{��ud�=Eo]����$n�i� a�"7[�嫳�U2!e9��� �� ]s��}��7�NZ��p���4�|6y�A$�M����*ABlQUuv/4�<��y���wf�_*p�<�up��ٛH>#�����N��oc��h�lo���_�;�}u�c�Zϑs����@|���D;�;�@��^;5�Oė'z@!&���n�#�����"a����vG�]�.�k�X�7cܑ$�Q�Z�7J� �m�0۟�g����[�V9'?��j����>�D�l���N
��˴�pk�iI??Oz@'��m��wf��Ve�B8�J�\YV$�tѢI/ӼܢMQ'�c���~&u����M@�v�&�إb��saa��� 云 ����&W`Q����I{7�B@?">�3��~��:�J��y�J^#�x3�D͑�r%�B����H�/���j���aZ9�g_�zþ��U��2�#�%u����͇2ǚU;�!�vj٩��<ͤ.����a����iM~�	WHgH��%����z�2�H}�q,��kw�{�M"z�qM�Q � �$�}��&�F7+遝6��uWV���!1۷O ���k�d����ie�Ʃm�X�T&�����}��H����7�o�	}�j���vy�{��;�x*{��O�$�c���]���X"�&��y��,�Fû��1^������%����f\��<:y�A��������Vm�l�MR+ۄn8F_����o7�|� c�t�D�H�����}�<�(|�ɻ�$�7�W~��qJ�+���7�w��	|�w���� z�j�@ �{}ˀg���NZ�X�?�'D�m�eW!Y�8�J���b��3|�oe~/�Z}���
�ˈ ���1h`��J'�}$}�,%Kh�ۺ۶%Ov�F��K�(�^Y���>�5m��H��f�`�¥�'U��k�OO�ҽm癮�n�����X�T-
D� �Uڮ��@���8�n=��9\X���9�'��n^�N�f�-�MB깇8��ϫ6S��:ܶ:�m�<�Fgle�=�;�ZP�s�vNgq�b˽�@���g�]���l[=���t��^4tܞܦv.�ǣ��s��-�oY�O<l
Ѹ�_9�e�95��u�N�I�Z�Yʰ��㋳�w��-ٕ�P�m�1�L���{d�x�!���*);�gm��K��yDܛ��lkk�����������)j�zw;��h��﹚ @~n{�J$YoMF����t/sh�I��t������W�c�Sts���	$H4+�Ŕu�gG�W"I$�vy�$�sޒh�oy��nwg�)��sy���Z󫜴Lr�93y��3@	g=���NZ��d�<���� 8���hbfo�����r�ڊY9��x����w���� VN��I�K}�� %���<�m�:�%�o����qG�-+ǈ����{��މ�5.��W����l$M'�$ܛ��Q��,��ݡJغ������5{cO=��!��ݦJ�U��\�2v�9'��������	+�<7�b� A��{7���������mIk��o�� �&g=��h��z�6��jR�s~�eo�qJ�k�}*��J���p����Qv�`]�`���������aLk͓�v/����咺_F��3�`�؟J)M�|���I����Q$���tE$䧅�^����j[��`�5Z�m�"�{���� �>{5�h'x��R��v�%���Ikw��I$���+��z�(��Y	�z���]�v�%����o7� ��f\ ����{q�q>bO�ğ�ǽ$���>s�6� _����o�3�C�m�=�9�,�/��оf�1�ޒ~$_�5a�@$u�=����/��g,�g�������<��v2�mˮe번�b��j9�|��f��X�i��qz(�:��������nx�k($�]�ш00���'q�/Q�ﻛ�����3����Ss�WB��s�z}��I���sԬuV���"D���̘ �=�x�U��+3�3��8��}����[E-W1�9�h����߶�I)�����Z&��X�f+b�V��o[$L��+�*z��eU}�Uᶊ+�Z���; m��A��}���g��<�7w���$�M��f}F|���=��}7��D�V��m�]=N���W�����_'��'�MO<� :$�M��W��}����?��T�|�@�,��A�no2I�_�s�Ίt�kث]Q&�_Gl��ojf�E ���n�Q�<]w�|j��9�8���c7d
��0n̎Y��䎷"u�mi�r=�rv9\�y��B"/��y|�a�f* |�Oh�=�{{�9華��Q�1Ѿ�o =���3�,��N���p0��wt` ��tc:�'|s���H6�	���wrK��d��!L��Ng=M*׾�è��Pш3��n�ğ�sw�B&���M����O/cx�G{���=�{{�O��bhw��^^U��~3\۔�l�֐��I5ٽ�@g��o{ {�xs��&�,z��PӖ߄�;�$�!R���tfgd�àaJ��[ϲ@&`�W���'���\�����г��O�]�)-��( l]�A;��g�� {��f��b�ʵ�(��ל�=�w{���=��w��ï�������9���a�nSn荵�n[�	�g�	\c��ze���v2������D�+$�^���(�3��sk`�@)�]�*e�;v��癜���Z)��&���w���͜��'~�ۗ>F�ә�>�|�f�h��Z��&�/���I'���d'��b�ˏ�d/���] 2F:Q�XW���{��퍟����@�h���/c�o��$�i���B@4}}7��U��ۇT��P�:sӻO��yc�/I�'\�r� ��F�В
5����a�Ț��=�Đ�Oo{�
}o�~�ZZ�g���b���E�v���w7����$����� #�5�Ĩ��߳3��筋-]�-�N]�.�7e��%�.�!������〆�՛��u�,nf3����2��0+B�*>'u�:'eoU:���6X��,�V�U:��(�̺MT��!�/�M6�hf73j�f��2���5 �9hf  �b7�U�t �E<������6;z��sF vƼ��'{��q]���ݩW��j��3�Sթ^_L�9o��
�3�kyM�6:��Sn�#pq��$�"�7/%��tU��D�Z�tR��IR�<� �G������4�#�!����p˓!��>��N^jyE�#�kD�4PJ��i��[C/c�#&]N�M*&��//;�d=ټZ�&:�N}Yb�\k'f�&�cOp	WBJ���T�s�;����Wm�v.��K�2+B�\hS'�"�|�ʷ������hU@Ⴕ���D��ՙyq^�	[��kC\�9n�s���Y] [��9kn�8�]:���3�μ*�p��ˣWg+	��k)�t{d���WS3�g�d=����������w�kX]j�<n���Ի?w��Z���^k����]1����!F����ne�@r6�Wa���7��n��؋�{��W��c&B�&oCtF���Z4]O��%��hI�i��e4���0�j��:7*d� }L]�X��+�W�M��Y!�Z�XȖ����7��b`0me�����aə�r��&Xc�[�k�
�qn(
�'^�9 �dj�j��~���
6�r��zZ�:	Z��DT���v�Â�w�qVeh���ll�cm�6�dH��l��nv������5{ݣ��"�����"䎃-ó�NvomI�n��gjge���{m�d���(�:�9����io{�{Z)�5�����y��a�c�u��[h�p&Y̛�3�:�+k]�n��:/*�2ô���S�aL�qI	ʹ�@����e�`�":w��=��6�j+;(��n��(��[3�n�䈲��������"��Y���E�E̛��u��8[]���&v+�D�=�%j���K;6��Ѣ��5;.��/++,쬬����ݝ6��ۥ��m�{���۷ w��G���U�r��p�^^1�]h���v�h6�*���8z��ŵ������"�+���=\�/�Y�]�ŎB*����?�|���=�z��n��n��)�t�v9.xn��a����n\j��Ps�g�h%9힐����S����#�g�ȅ˦�O��9����Ռ�ݍ>���nv��lUe��aζ��畵\n=�-��ݰ�㭵崝���N��v�[��;N4f;un�+����:�KX�����d�b^ۡ\Õ	�.ݵ۝W�m�jN�D�n�l�v;��6`��K3눺m�[��L獔�.5S1���;�t�*��/N��G[J�OO49�&����_���|��n���,{5�lb�N���y�7�����pH�&Ք�	q��]&;s��Ľlm�Wm�{;h�"S;u��������p��`���#vq�x��\bZ��ø`��1���c9��nW==����b�\+]�K�ɇ�t��Ͱ9x{�����gѵۖ�N�d�S�-N@uhѡ��9x�[G=Eȝ͝����ƻN�zƩ`8�'.�i96��<���fX-��|Y�]�m��r#VC�i�F�^w�J�ƭ�I����5ٷe�J1ivv�tr�b�۞�;[#�v�Dx9�l[���R�˺n��M8zt�ݓ�^[��M�.ێۀ̯ 8ls�u+�<n����5���{&�n���sك���Qv��:q�v6;sOU�R]��O1���O�k��k�����qlA���=b�x�k����v ؽ�Lk�F�:��:�6ڭq΄SO�ɸq��$\&��6i�y���K�t�<�Er���͍n�j�M�q�����x�ù�m��쉻Llƭ����O+�hCm�n	��P�Gqu���r�U��l�ۧo[��Rks���\lw�*�k`�D�k�$k�ܗg����|��11�Čh��q�3��3k����7n���Ds�r������M�8)�; Ս�-Lٶ��-֭���9�v����8����n��]���M���E�7:;t�kn3���6ݳtqɧk���Ƹݺ6.c��9��q>�l�n}��w�>����Oa�wm�OGe�.y��^�2b!��Ύ15���n�q�g�5����l��Ļ�wkR���ԏ�On�����:�;;[�wQ�ŕ䇞C�\;�cvv�� �3q9�dMU�v��0e��I>��z��poC�.�=�����d8D9�d������>m�+M7�����BI5�:<�h�$�j�ny�'wۅٯ_��&�$h��+�����.XW!&�����2�/���k���}���@t��\��3�Ϩ�׷��7����� ^���S �߫��ύ=���@�A����+`O��q���[����y[o��Ϩs��L��Yn�tg��?w��]��|I�pgD�4I�N��;j�4���\QwO"�z�������G���8�%"��|�|�xI5D���!�"�o����a�QK.��Б)z-���$7��w �ټ���^����l�U_p4�J��o���mGH��j^�����.-�UD�VϋF'Ϸ�(!?}~��<�3���C�w�w2��f��n�5T�*�$o����0��a�!s[��[��R� E�H'fOk�	n�U�y��>�g]C�=e�Y�X6�u>��v����t=�t��ÂbK��c{r�]����k2#f�]%�VI`'�����V<H���� )���� ��7w�U�"��:r�t۫|�al�vf ��P�9�w7��=���fY���W��rl���6ś�=����nrJ�2'~�۫����=9+ۜ��	P�t���������<{�"���A��� �l�s��Zo=2�Ye�#~�{����	7��V;��q{ϰ-�?qێ� 9�7y$��/<߭O5ǯj7����dvlr2gdⵙ6
n�rK�^.��A�ٌ�M��V6�W_S��=�ȡ���=��$�o��rA$�yy�]죵����F�{��`g;��{A>��O�_�-A2ǧ7T�&�=�8؏�o�{Ntx%���I'�c�� tN#�1w-L�Sޢ�ߥ�(�B��I;��g�O$�v���MQ7��O<��,ɸ�H���y�1}Q]97.e]�oa��srP�Cv���y��4;���d�*�U1%n���,�����%{�߹��i����b�kέ���2��tO��V���M~�b�D�^�+`��C��\ �7�3;Y:uq
���!&��yvH�>�9�����Ȓ@�g��*{�����TN��7	 ���� �#��'���O�Jܶ���5m��-��w3Gl3�nBx,�w�=����vۚ*���_qm>���c,����sݝܒK��<ш��:�mW5�>���^7��$�HQG��b��4uG%�C��Oh��=�`N{'n�3k` N�s& �Gy���1�ٚ�=!���޻��S�x����j����G��%A~��qd Ay���|z�Co۞�7�ǹ�F �s�<�>�.UP��`�wU��p>�ړ�M����j�@$;��1 >�߹��8#i1u�^��(�Ý�w;��[WaAO�ِҮͪl#2�P�˶f�0�tA���U�r���i�z:.�R�b�3.	�fu�8c���~�al�vfu��� g=���o\�O��I}d�ԒI7��ߩC{������Sκ�T�T�[�kx�Sm{&�n�Z�Pvu�ۆ��7-�.�HO��_e��߭%��<��fhlA�K�vI$�n��N	�s�ߘ��F���C G=��w�X�~,-�cĻ�N�M�-��h�L�����b_$���ش$�I�~���	.���dP��w�[ǿo��@�������E�y=Ր@�o��ml���k<���%�Zs&�e� ?�4���%j��B�ꭩKS����s7���-No� ��o�g�@4�w��D�$���1"��w���-��d��N�H�*e�'�������&����HՑ㇍��,��6Y&�?-��'Ā~6;Ѻ�o��ʹײۋf���t*Ϩq�{8��T��ձ�������Z�LA���̶nsV���N�9�U���5�N.�k����i�Wp%8��䱱9>v Ƿ.U�X����V��@���:��r:`���������[�=��n7�[�v�{66�3�\��m��m���w:�Y�Vl��[�ڷ<㜸���{��:�jf��W=&5�۴�r�r.x�:�F{t������_����yP.�s۲���֮�#�c��q�X��sp��&0q: 	�-���+�`��*6Ur�[=��wϟ=ne��S�n�Oz�H�]���cq0���ߟg�~~�4�Wa'��?d�{��mllC��\%K����������4���!'�W�d��;���߳z��~��w~յ.#�I$���%I5F�z7H�N8��=�wz��� �`#F_��+WwA�=ۭ�$�M��MD�NxnR��ǳ {���������E�� �5WT)bߒ���<������%���yϡ?I��E��$�:_��a;FFyg�I/{��$�阩�7`|�~ĂI'������z+�r�2I$�D�h��F��ߓ�K����eɬס׉?cP�����'�V�Ӷ9�"�pI�ù�Sr����D�&����|�d�Y�}t�O�%T&�4N�$�{�e�O�����ܞ��Βh���A�Q�V[k+�I�����!�w��a�a�^�Zk�%�d%���`hX��+0*�mX�����i��!w#�kf:�\Ebk\O-�EQa|��fk�B�@����M~�Ԑ	%��۴�J��Oe���p%Q�Aȝ��]F��޴� w9=����s�^'�ݢ@?�z7� �~1���IN�XBD���Ӡ/8�-���]ug��$
s� �?kϳ�d���7X�3B~�fX�yhI �<��E�¨v8�p���s�Y���ob�RI��X[��0oUG�֙$�����D���wrS�x<�s\�h$OE��^w\=�nSv_Jm�U��s_;�Q��!p������X���=�5�ח���7d��9=�n|M�e:���vK�� =���(^i��A+ke�'�Z~��Bj�������bѢ���r�߷}�y��{����&�y`�/wߖ��|r�[\��&b{sz0I'��{�K��o�0��-�e��Ƨ��?^(:s�q}]�5���b,�]L�k
��4�^!*V�j�y�ʹ v�m<ߐEw�o$�SϫV������Qq&�'�/���Q��$$��̱�'~���\�s;�շY4�^n{F��%�H�����I!s�f��r�]��~@$o57��}�'��4+�ڰ?��ތJ$
����G
�:ٺ�n�5�g�I4���%~$����'�p޶{Kj&>v)�eD�Em֬���Mq�t�N=eɔ���- GD�q��p�%#���ާd�ﹰ$�3��:%3�O�ߨQz��-.n��"�I��wp~����[S�
绚x��}<d��WA#�_Ě�zn��$�h�o�����=��o����ei�ʙ ����c�v�_����o{�}�k>�� �^�r=vE�j󹳩 �Z����`| �}�ϰ>��s�VKl)\�+��<�7�jW�M$�O��rD�j�wkN�4I3����H+ڱ�A_���f��-b������	�G�j�G��7���[��<�-%�x1��Zw���W���O]��G�;=�E�.6Ex]Z��~@Nk|���\���"D�в���f, w��ϲ/8�tߤ�)��$2wN��$A�{��	%ӫٟAm�׺���DH�1�O����bY�l���
\�R�vn^�Zg��������N�+�ڶ��{���� W���L�<�w^�=��P�\�b�I(� +��3��U�R;`�p粉rC�(1��7x��I �<�	/�K��n�E�KM��[c}"J��a����R��M{������}Ŕ@$���<5]�w��H_����$����0���Vs�A���җi��� ~�]�'�Mk�睲I*{���5u�f$���X��EIe���H5�{Ŕ���1��Y��! A�F�ĀN�o ��t���ш���{J�lz��^9���t�ڥ�;h�W�ŭ��lu�>�PȽ�հ{��/��K��b����)S4�7H�^�G<!�s���;=���'.��N�Kd.�k�6-�R�籱���0N:���0�&��txe��뤝4�8��`av�H��ֵ�%�v��G�N���.;v��	��]�q��G�k��"g���
�����ѱ��A��	���svΩT���u�Pn��%���!��<d���]����[������[&MT��D�wW!�u�����n�5�<G�Qș�Ɨ��0�'ģ+��=��DH��K/�\z�u �	F��6��$�w�;�%����5��m�>�<�a5�0~6��33)����!4H�e��u�r���;7�� k~�w��oVwk׍oW�Ņ�Z�R;h�Μ�e$�^�ʄ�I�o-r��c�󋨒K��X��o�����vjN߅`!ҷ�B���U�[��Ƽ kg{�e6��'q<H!s�l�yus��i$��fg�3��s��B�_���k��%���_w��X�{���ML\8z{�1 %��wrH$E�<�5_��{�Y��uC��}N(-v��gm��G�=x^;u9U���8f�v}UL�V��p;�!l�VC^A�7�$��r��&�#;���^��ӋG��g�wF"���7I���j�U#TM�uuz� ��tj_%Y�������)�Ό2Mk�ҴԷ�Xκ��%b��W-E���v>�-�1vڮi�l��9S�4X��S�9��[WZsO[��	/�Cc���I$�绨��C��,�w1l"~�n���Yt2�e0'���T k;ڐd�$/vH�c�ޱ}�տ$J='w��3�4b_L��V%�R5F�Q�ND���ڛΪ��L$K{�orI$���:F5����8"��o"ޛ%�7�wpI_����]2�<Ċ����h�o��R�{��V�>yȩD�{u�D�0w�:DI�7�F�:#[wP��u헇e���
W��3�؞�[H�wF�y�k&9	�k�9D}"����G�^_RV_�k3f��(��<߰�I=�<��+�a�6uH��Yo������ϴ��87$-���f$�{ŕ���^�.�	�{�Զ6ة�sl�Lk=�L*����o���I����9�Ye�=w�� o}3ز�$��x��ͼo�^�gR��9��k��O�k+��&�n7�uLh{�:k��R¢>�X���\:sA��6���N�a�!ï%����]�Q2���W!\��4^,����Cc��2�jy��L��䥎���?�tVM�qh�]B�K��_d`<ƺe݅9�|Sܨ���:!��&�n���]���]e����r�23*��gP�����4�9N��PϬ�7Y0f�/`����e,��ב��S1�t�#�+1se��8S�S����Gg.(�)��z�6v*��
���i�8��x)���/1��S�m�ȥ��ؕf���-�EږV.G����K͡��_e�;�̛�����ݑ�����9�����{�
�9�z��/�V�|�طw��Ӈ,�%�;
�c��:qn�v�K[�C �Q:	m��$��'.�V�7p0�C��7�9�c#M�-q6JnM錜j�;��}3��.��o]c��n�&i��W[��U�V��<Xx5��ѩ@��6��0�l�E+ڲ7V��2�n���k��hIU�s!��gE5.�^��y���r3�$	�N�0mw�j�[�`�h�t��v�|T��QPbJ���n�<��5����A̽uz5�c�]����v�^m�~�8=X�����{�M�����s��JΣeeԔ��V�]��{�a��)��t^bJ�c���e��8�S�0k��J�kL�+��v��U�¥�trt{X^^�v���;P�B+�Щ���꾎��f�T�����J��cz��	����{���Puyxp���H;kYRe�3w�𠋍,ö�D�3h
:��⽶U�Ia��n��Ҳα�k.�T|��86���l��<z2=-��F�����i�f�8�'yztw��'5�+{yם�f�M4�D�d����#+m̘:w�oY��bGzY�sb��G$F��mcl��Vkn��K�v����E��[T���y�jΎ���+ �͞�^��e�ݬ�۶�Y�%�{Ǜa�k[n���7�U��Lɧ[n���S���8�y��X	����Y�g�)�fy���K�Z�Y�N�mI��K�ԃl�-�V,�mZ��ͩ�4u�{��$6���7L��ۑ�6�dΰ�X��21�������dg9YW}@|_��š�xg���sXψ��t��w�ޛ8�A�ڱ���y���&�D�{��D�K�����w�yךѻ�� ���3�Ϟ�W��r:.� .��=D�%��9��Ű�T��v$�w]�� �i{}�B`�Ӟ�����h���H��:+]������:�;�cpq�Щ����H�biF'���z�6�he�y���2<;���A ��k��d��.{A�I��z��4{]��&�W���!4���y��i&a�x߹���V@4O�ߑI4��� ��s�����h�'s�pnH[e6[�WKm�����!$��;�oo�zjf������r{1A�g���hs/-�A����.�kә���xwˉ�</`���&��.7d�D���$�@?�\{���n��ĞE��/v�1�=���C���F�z�Ul{�*�C�Mtg}��	�L<�-X�`��ZeA��OD��W�!$�+����X�8��:�#��{����ٴ����ؠ�ZV.l+�Mt��.�$󞛼D��ޮ���{-�Qn�r�ΡB�����pV{N���;ۖ6-d�X���O6��1��6�����d���$ߧs!�M����$��\E�O�����v����������~'{J�v�2�Aw�=/Y�Ȯ�a��8r�5ki�{��w�� H�zo1A����v���ַKU��PuV'��Y��� ���x {��qss��P }������	 g�o1PV/rq�$�[��,�D��w@e\��0���Knk�	�M__Gl�����s�����k,�$�߷���L��W�-�,�S���H$��k�>����<�Y�$�z�w|�	��4R)$��{tR��^��4�^��'A�+�:5���L�\̋��C�u�:��G� �ȯ<��������[��m��1�&<�/�������o�{�~�Q����#������[^]���`Ҵv��cY���z=�@��
����)� Spͦ�)��W���f���k΁��i�Ǔ>��K�a���.];]�xl	��=���]�1���r�V�/e豽�%7ZN��&r�71�!��q����n�cq���m�w�r�%i�Qz�;K��۶��Z��J�<�����k�6Û�����t嗲j�W���͋y�؝����jkYҦ�ʥ
*(7WՃMX�m;lW������N�j�����{�����voY @s���	vk�d���|���v$�Ig=7��u��l���c����=�d�:+�"�릩�I�^�� 2D�~N�$��֬�96��I^�WSp��h�9�Nk�9ܝő�%��c#]�ީ��	/�Io�]��"�F��ي���rtE*�i��oہ���������ɚ��Oh���;��.&*���$~�7i!t;��rB�*�ɘ�]��dlg;��eZ^���$�-��x7�|s�=��>{=��{�7�L��˫s�F@��P�++Pa�sڸDy]�o*���*�pY��۲ر֯n?>��j�(��[t���ә�@H����dMg�� 4���I;���K)����z{2�����N+�Z������ e.�^������a����T;!Š�\�J������H�}U��н��lv]�}2n��r^�̜�'�YW�����uR+�c�NfmC��1-�w���I$�g2 =�� ���<��[�I����ӳ�v(B�����,������ ��X�����M]�ލ��$AL�Mߩ���;���O%�$R��Vl��~�z9�����VH;�Ng� ��w��������[g���k�W�7{31@�j���B�A��s��D��^��v{��鶏uC��K��e� ��h�g�{�P��'k����C�������]V���U$kv'uQ7*n�l{#�PI��ӣ~}��O6�
�Uv�~���@׽���I��޸�'5��;7r�3z�ݐ~���{���7hナ�e��o\�I%E�=ދ#��n�/�A%���Ě$Aމ��4K��+���vMTj��H�N�jǄ�=����$|���D�H�� }�J�֫�`K��3����u��#z��
�<���%�X�������+�����w>E�pU�B��I���a��8SJ�I&�z��I����(���m���_,���d	����+�^����$�9��6�����zI$��������
�@�$�%ywI	3���������{^I���|��7�|����j��IQ'�~����I��o�A��V������~�[9��(�m���(5DTB�e{n�2`��k�9{ �2[kQ��M
 k�k��xD��$P~����} A��M�n�hI���]à]�{��$Aq��tQf�Td�e��f`gw7�do����|uנ�޼�`rI ���l�	n��H���N��������y���ܲn�R9[E��ϑ���b� �[��,�@ y�Z{y���i����6}�3��w�ِl��Z�rզ���B0�W?_���5D�ED�I[똴�_M~}��9�:=����'.veQ�w�뾍��̧��2q�}ɓ8���.��)��ӯ���%ֻ��
������*���_�"kW_�d��V�{��� =��3kg2��~�7h�̍�M��@�=�����d|O�����97TTJ�"���&�@�VH�hR�(��M.FvzWG߿>�kUB��)[�+����@|�gs!�I&�o�@�ٱ^��[h��"5��f(
�V�:�q�*������}��7\��·�\J|��I+�~E�H��d|N�H`w�%<��k
�]v�n��46�7�s:�6 [|��� }~��	 я���d js�I(�k�M�
G*l��<8�����}W��a��P $�e;$�$�y����M;�����ggS��$�um���THd�eF�Ɲ�z�'i�_%��f�����9�d�T���oڴ$�IG�;��� ��s��xq�U���?y�=v�K�AY�*������k����K�q�����C�fj�n���r�ر�����2a]z�����釯(�@��ع�'`���ݻeѹ׮Oa#�%v��/N��{>��c��si[h��ɜ�M���o.����{>C�S�g���9x�)=pl�x,q��mn��m�3��q��^ɑ�Q݇�1��!j}�KV�pr{���<�g5˲	��x΍�� &w#q<�3h�ZMp�W�<�z��-�s�5�!�ٳ۝L�q�xЧ�\�:��<=ɸ5���X��V���v�cd�o�o|��ru
*B�j����=�����ձ�  �=6�-��r��aa{�SQ$�������r��Y>%+y��{ٔ ��-�ݞ�� ��;�� ;������x�F8�S�b/�����)X�_����$��{��&�^��&���ډ���q<@)��tZ_n�'�]PRJW,�wsy~u��d@=��6�� �Ow& =�ڒ�M�(Z���;����ɺ�#�6Yn<���*7X@$���ӱ+��Nv���� ��̣���ϡ������in�n"D�ƇE�T��&Z�caѳ�^��;�ns��4��l�K*i��@�%q�9j�|ݏ}��I����I$ۿjԥ�`�_����ؑ&j�7�i|��2�h�v.ƭ	l��Z����r�U{l��ki�	D�8MF%_3�3�
��{ƻmɽ�h�d"P�9��*`8���ڮ�I,��B����edSr�Uo�I}cĀk]���MN�ߛ� ��z��=^G�Ɇ{���
��B����)[�5���Tl�;�N�Y���{�fʺ����#�ReN�ۯn�Z=[��T�2���3�f{~�Ի�#�����K����x���r� ��wIw�����nIy;�D�����xS�~9-��XY��sz1 �{��c��z�my$*Wn�:�N:��R$����ܒ���탡Y��j���h��n���[�b�y�q�I��np�+j n�D0�")I�p䝬QI~r����|5��> 7�Ob��f���!*��{��༕a�$�gK�C�bzt!$"��7�s3���&u�Z�}d$��'�@=��e�~$�{�I���UW9�vc�cg�e�H�F�]�Z[%{F�$��7��RG=�/A���tv��@ن��""���.�kd��u�mP(D�7�λ����4���bR� xw�#2�D���_$���j'R]�I��$3꒶��7c�8��C�������o{�}7�70�u0 ���l�>���_n�i�1O[��GWhTI������gG�Wv(�fA�-�z1(��>g�:��r�7�������q�tI'��́	?��w�^�~�����-���X%
b2���H���v�z�$L�㫎:�p������~���
S^=oy�h@/���{��A,��+R!Ī���x�6g�LE �rI��y򪮴�W�WxK2�Ȁ��z����ق_�_y�4 �o���H���n��TOw�OI�\�<��MX�<4+"����y��a��=�`�J	JB��	(���q�)zm�N�'{��3�y��3�{O���V�C��P�	�ΐ�d�~���M{}���,�vU��?8:��/j��E��&˒z�ϲW�W���#OJu�]�I��W.���7@݊�_^ܮ�{e�D�r��z�uz��Tz,���H��}�閦�Q�Y[�<k��� u�GML������8�f/t��$����E�����rt��ǎ�9���k\.��V�3ñ��^dtt�����u�c��:ع�~�����=�D�S��U�O��gs������  {yp.��_-�yn+}[G��Iy���$�O\N������˻,���<���z�J������I$���DHѾ��I��#ȧ�{s��o�䛠���Gm��z�f   ��h�~$CE��}��x��#���b�>㏜�b�ʰM�Ed�Wc��rt���{�z!L�I �[���$�>1̽I$���eK�w˫�}�����55�EGb�a����}�l�g���h�&��*a%�de� ���F"�K�ɻ�/|��(�Wc���ųE�u�����N���PS���SG9Ks���O1<��k]�7M��v*�'s�|�JdS��u���:U�;�%�dV��UV(c'����8�Z�B��g
V�me>��˻t��� �j���X������#Iڳ���rdS�&T=���X!��u�xc{�X�S{e���[ڲ�����k]U6����'^�Ɣ1Mn��6��&�0:���R����^sD\�3�)��9��3%���c�v�c�-��xr��5h�b���_c�S��fK��+,a�sX}�Y�oaӗn!�yL$\{{����AZ�cJ�Sd�X(0��1�cy͕�{�vQ}Y��
-���Ve5-�X�2�+[{6�L�`x62�n�$5{��t��Ȃ&�)A�}��n��>�h�����7�kp��e�t�Ϲ_�c,�4�m�5�+oR�4�͐��"oEݽ��1+�I2���3�o�]w;*	/��U�w��X�n��kfB�)�A�Y�Q��O)ptN�qf���w��u�*�Z�q�qr�}ͬ�.�B0�����]fȰ�a��`gP�����M��Q;�PwnmĠd�jn�����vkM�-k�3���ّ_(���BC|�mu�5t[җTs�J�3e�*�sn��TS1K�]��>���d�$�o/�jV[=7����.�7SYn�e����+��ʪ�c̣���CJ�b�z�İE&+<j�p�k2���\�[Miq�]�l�֙�X�a�/�ҘBCb���7fe2�-p;;o�綸m��`�+E�f͔s��m������l�!�Nٲ۴r�b���9������;�:9;׵�l;0ٵ�����$�.�;�G�x��L9m�g�k	��'yn=��݈]�Acv�;o)�3�'m`���Y�	m{z�Fh-������yx�ݧ6Z�)���[�mإ����$��č�,�ݨ3k6�X��Y�M��nm���-��m�H�3�3Y�+k]�iC�'kV���ƒ�16��lK����c`k���C�V��m���K#���	ܤ�im�����6����%�[4"��e5h2����v݋m��gn�I7���iM��Sm���$�X6қq��Y�4�O�i�1�sUNRu�k	�On���Wm98�v�^�^'�-�:�l����5v"�V9�X|�F^^�pۘ�x����#��g:���M�q/v6����4�3���7E�>���ǎ�l�Nz�^�'b7r��� �]]i�=���]��� U��atnce:�h�4;l.��
=����m٤�K{m�ݐ��v����M��+ct�.��U�ݴ��ޫvy����'�w�yz:��U��kAM���ɼ�����Ug	�Qy��{A-�p�/�]���c�s���y8��-�m&�h��3�02{a�"��yz��F��7����gF��5]���������6ύ�h�n�7M8�i�۶*�x�ҭd�Ø�^pgÎ�6�e�#+���G=�[L�;��m�"��u�\y�q��y0�j���l[�6s������9�lAq܅��gx��9L�s�܌�ܼvͻ>�3��:�����g��������Ƨuv��QKv$�ŶO4k�A��9��q#م�8�Ue2��u렎`m܄�v��G�K·�=j�rxq����������sp�9�zwMg��H��v��t���.5�9kuˊd�dx���<���zyp���q/��Ů�"G>����;f�x�۞x��5�t�fG����XxF#�Q`J��r�3�R�uֽi�e��t���li�:۞I����/l�9���0��1�؀Ϸ2q9�uہ�<kkm����sxf�Xc!�X�`�"�Nl���kv����5>��;�ܞ���;g�8�ţ]�ËRɶ7��sY�F��n\��g͎���Nx��s���Z�Z����2;�]��W!�s۵�v�J��չ��&�
z�L/Cc�8�8[ơ�q�h���/GkOB]���t��jSj��ۄJ7[�c��7�탃x�o#�vy<�n]��7������@G����᎝�v�Jyn�$Y�e^
.&3uU��,o*���:�[��v�@�oa8�|��C��J��յ�q�ؽ���-�
�vy�
7E�i�6��l��:���v�^4OMկ.�f�����=Y9���tm�6v �L���q�[����x�vrt�Ԭz�Z^b8.ͽ'�cdl����s�ʫ���1�om�ԇ`qv��b;v�G;=pcmgYRKPN�l�gu�{n�rvwZ9�v�<�i���pu�z��v��=\GX�h��u<�x;W�Y�<1:2s)����gemX����5�9����C�В	z97y,ũ'2��:�e.����~粼�=Fq�T���hA�Y��w}�%�nQ�@������ʹ�I$<��{�H�����I!O=�����{a����^?Im� �k��:����I%����H$xV��ɷ��8f�W��	/�Ax�7~�W�%�����HE��b`6E��w��3�z?mϻb��:�^m$�w��I=��{��5}�g��HǞ̯&�	�4*�P5v4���<IO'ٿZ�OF������$<��oRA%���'�Jy>�4��g�xs�s4��7�VZ�v(+lz�� �< ��W0�,V�x�N�Ur���㾾�tvKeBڳğ����>�I���<d��<d��m� ����O���<� ��1�+y���s+���fnmفW9��n��ex)�Û�8]1�^�r�KC����@���Ԫ��6t9�/��tѮ�t��4ȼ���TڼM	[�"���n/�A/G&�$�AC����:�ï�;�/gv3���'ΫGM�9��}������u{}�o]�)�����16�o�=�WJ>���@
>�ct��߉F7t(�{ɀ�}��ڠA=��~�n����'뷾���ǐ���ύ�n��`���^V-��t�P����$>g�;w���y�e������ɉ����O�ENY[���k����9r�`�\�ʱ���5-��g�|J������ހ�LP$��~�}A�h��X�o9z���֬L�xs�lae7GnOn�WQ}��?NuM�d���g	�SVA?toۤ��/q�m��2|�X���ڑF8Z5!����m>g=�I �z��z/!1s�td<1#��wa����s9q���ûQF��4���"�gK����Z���Z�7oQ��3:"/]��Ͷ�慛*�����H$�SpP ����A�b)�,Dh���ޚ<���w�瞩��5��XH$	�M�~��� |.Q��p�<��HxrJ���_�g�_g���/k��ڵ~�p��򦻼������zi���_;����-��W � 8�e�h�{(n��]�6��k`���t$�D�ξ���G/Ĕ��|���	=���$��w�Cn�W��g��\��ZM�k��,�+߰����q��1Q�'�/Ufz�$�����k`�)z���P��ޤ;>8�4pef�n�u�ݣA>n<�	z�]:s^��Jz�@&l��$<��'D"�+$]آ,����hV5��: j�n�����$�{utR�<�M��2=��g�hoO*�sc�yƮ���g�%�nw����[唲���f������.P�,�����]>r��E��P�'�n��|���4)����� W������a�2���]@q� ������]<��[}n]r�NeX#��_#��Ğ^�2��l\�=�e����#�ev��!���_��J�R1�U�������sX�M�~˯�s9�[<�(<�Qj�����T����3,���8�½�/�������/�����n�@���h$����s�o��{3[*}��F�$j��ߞ�?C�n}�>�o1S�j�o�P W�z7@P�����u�ӦQ
���y�9�o��ֳ������I���HN{y�?:s��i���Z����B������x����UD#J�]���}������gN�� �ĵ�� �]<ҡ@}S����3�_�ɫ^}d=]�X��@�R�k���E���d��VH�cl1��/�;v��>�&�X�e��X�]���+4�,Y���k�nXo�[�(�ЅD	Kd��/c�������E�c��a{h��͗,8ɸ��"m�g��&u�M��r'k\�h�h^D�]<f��3ړۛ�=]v�:v�ca��8�zлw\N܅�h7k��u�#>x��y��i;zӻ#�>�<ɕ\f�s���uˡ1��f5�>B�����yʣ.۫InJSV����'8:V-������t�ښh�]�������e��q�<�O�G;V�6_�2�&80k���7<�	��k?y�����kT��S�|�K+���{8+����ر��7ܲ��rJ�Q@,�����;\'��'��״�<��Gs��A#���7が5, j�̣=�|J�<`2��Í�
�q  ���T�9��y��ر����� 9�R� w��t�0L�5���H����vx�+��@W{�@P�G�6(W{z?(�X����(Dޙ�����U��՝�vzv�y��e?w�fy���$��^O�M�I O8�O������TY�g�k�G=n�1`��F�x�� �ٻX���v������mN[�R�4���9�Ѥ�t�ڙ+����(��,V{��bM�G:�Ѭϗ�7���7����$y���iƸk�LuX�1�Дh�Ϙ��Z3������/���|ƈ.Z�Tu(�]�s2�͞}]�Õ/)�R������A"{{��(,*-��y<1r�IU��ʼ��Wc���F�A�90i'su��w��P�L�ٿo�yɺ{�i]�X��B��|�c����oF��=�́@=�-���O)4i|���	�4�0���9�s16�����ʞv����m����@
c��`�P����.&�l�D��t�GX��ݟ>N���z������Z�
�%g�ߚ��,����MZ�MY�+zxi�|�y����k	���\=�ʻΪ.��������=�H���Y ݒ(^e�BǔYJ���fTj�v� ;{[�P{��(P�{�cE��[(=��=d١�0
^I��@1<��(T��sީ��a�{�uۡ�WV�9WI�_^c�}n�귎v-��k�/6b�!����b���9��3r�`%�hM��.~=i.� �}�?��Ǧ�2�ʪ�V	�U���y��d7�=���|3���� 1�v��
�[���8���>n���<`U�|/0ccB�j��"�6��:�!�ޠ��ɻ���p���?h�P3�f�}D�Y~EC�}A�����q3��T�%�O+і焞�Y!�M=���h�m��L���A �p_ǯ����Ycϯ}�����R��[�x�x���:��}t�A���ʞ�A��ma�?n��w)�$�����[Y�����6��X_P��,�w&��Ў{�yg:���x��������#|uU*���aߛ����(W���"�  }�wΟ�w������=ܐ��Q�l`��A��7mN�0
p�:i;K�m<���`Q��}|L~�~lK��ZfX���+�t���ͯAӲU�G���'( �	C�ѶOo4�����'��g�nzL�I�n�o�P��פ�{�W�B
|
2��M�v�ݎ\���x1㧱��D��e'��8����e#���׫ )�:t{y�T5RK�\��,�X%����ܪ%K.�(�Y�yǺI�wjH�v3��I3��'�>�o6��5�n���=�3�[�'��x�x/y�n�L ��J�@�̿<��I/<��"y��'D"� &�/2�3�$޷ƶ?y��(�$��ۺH$3�kA��*�����K����9F���i:�s[ S־����T�e���Lm� ��m�@P���C�[:\���z���m�]x����6�D���u.�몛�n�w&8^d�ND3o�[�^���؛���*ɳ���m�!ױ�hD�O�G�wg>�+n���x�3к��!֛�Q88�q:pv������c���U�Xy���=����s�I1���mz�n����%i�X�����/��+D�^��s��o4Gױq���Wk�^ݐ����'D��n�+��kɈ�l��'u�=N`�Y�9���b!ݞ:�kqUr�x0�wn*��t��M�s�W�z�M����h��ȯJ��vG�齞��]�p����p
T���(��,�x<:�n��>w�`�	3����0'��'�/��;t�D�F�G���AUѳGt�>���!���o��� ��7t�I}���v�fxrX�I{*Y�^��ܪ*���+�����t�I}�Fk�F��~���@$���I ����:D)ZA�I�x����oͿ:(���K�0 �
��^/�T~�%�����qΠcكs�jRb�	���~�I/;�@�>�Gi��(o������2{�`$�OM�_�n[��M��.웪�j�]%����s�:��yL�x�ɢ�}	F!��t���3�ʪ��4(���vn�O��{w��nG�`��ax���//kb�EU��Uo����,�n�!����,��~ul;~��Ӽw��W���cFDz�xdt�ձd�Y�H��K��횀�SM]B����t���|Q�p��Qusyح��� h}-| ����j��7�/)V私;���
���;�f���4#��ӠkQo��9@B�}��;g��&f�RD%YIj��g�G�pXwFPB�X ���}���
����[<ᘕb����݋�I�x���Θ�>��?��NRǍ;.e��%hP��w6^�slS{���^�^��n��;�ܵ�^�B�kX�ݓ2�n����Vv�Y	�KQ�7߸��|�cM���5��ϰ�DޓF�O�&�q�F��(��ҥ��?o���{3*쁕xM7����
跼����{�{�B?{�=���񭳘��w��mދ��
�n���Q��+}������ɹ�%���Jߝ�����^]L�HV���EB;��U��ʷ��ё��$����[	9wL:���a������ۑ��a�R:����3�":R9��1VUN�)({����t%<R�SKބ7��غG4��F��s�f��[`�$�u#j�M�N�4�ޘ�7���`��r��� ���L�k:]��z������X9T���{�Z{xhu>ŧ���\�R��v;�Ě�����/n޼��M�}���C�����B\w�2����s�2���eu[CΔ�]vfկ�ַgF���e�d��)u ��]QO�>�ve��MwR��A�u8cu�대��wǹ���\�˱��&:5Xn��4n�ˢ�T2\��ң�س���T��E*���.�]R��*��U��ɒ�"��iڮRf�ꗗ]����5&��i�Ҏhse�י&�����]+׏���]=A�nӷ�۟A$�\�Ǻ���S7KV]�����w�`��9��Qq�b��7#�ۦ5����7�\��%k�r��fV լ:X�6�q�{�k����=wn�mg��@��	)�4h.*��8�켬����us�f��!����9�*�d�^�qQ��4�Pꯌo��6�ӊ»�q�Ed��O\�6���=��X0�M3 ���#���۴�KG$�4ܧ��{�UB*fnt�+�g=����e�"j��hs�svν���C(9�Mӈn�X��,���IN��m�����ݗ;�޸�6���>l.WZ�mGl-�<�WfI$�E�?��3S2��p�m�N�N�m��E��Q��7^מ�&�ی۱;5�����N�H{dAH�	:s+I�ӠG6���өma�h�[^�pソ�Cm@s�m�pm�A&a!��r���NQ��
m���2,����I��ggGm�s.�&����:K��6�[�k;-���f9D6��1�6ٓ��퐓�T�y�֒�mvD�T��PD'Y�m8��:	(�pR۔m�܁"�!$p�pDr8����YHGHm���8�����'JF�a�p�H����Hٻ#����i��i.=�r(58ٙȇ����%!��	�9�[v
m��G	__���!���=�7t���]dR�����;�?kj��O�(7�ݺH OI��@�ޛ$#\��I�
��y��<�H��@ٻ��; �Go�3ZNY���bj6 o�Ͱ(
��*r��5����#�UD���:�Ӳ���q�=u�H&��Z��r]k�ud���#o؟����j�Y���i'�{�nh$�&o����ƺ��-��`�=�M���
 �Q����u��a#Q�W0�0L���Ǫl����'�ͺ�(��t�����ڃ��T�bk�v)"n��3~��A ����C��+���A>���%6�^{zU���{N"�jjB�&s=���ӷxG���&  }P�KT�)ޚ
h�o�6��y5�u��9�.�s��^�QǜF#LT5�=���[u2�>#���@̮��NB��[{�*n62Ot��S{3���DJ��T�U�������U`����J�N��'�)��n�D:���=7A�mz_����C���=�m�K'/4家0�.�0�.��B�@+��R�)-W]��ܝln�ؽ���n��X ������v��ww�3>��MO����,��ϒSh�J���ֽ��Ôf,�fI\}���y"��0��M�O�nA'5y�^��s�H���U���3<�8��}��k7�~��jj߅W�EK���w��W�����@�7O�k�J|�^F0>�"B����l +��o�$��0���� �~���O�غ"��VA~��8�4���ִA&޻ω�7�l
����>�lƸL��낑g.����֬ȕ�=�}�n�]:%�@��R����:[��x������԰��VW]�Mi7[�2�"݉�_��q�S�HS��u�nۓs=���T��CU&[t����iV���#��sɣ^��۲��H��3��nب����u�͇���h�i�q�Ok̋�u��s��uS/4vܳ���\r���;M��Gvq>��e�����K��n�=��q��2���g���m�:�j�[n�Ɍ�oh���3Պ;��s�b@��qX]�W	/Z��{��lx�˦��˗��۞n�m�k�g����mp���O7��O(�GkU���w�ڥC��:`
��kl^z7���we��Q* �w�������P$a�˯_�c�O�gT�VO�nL$�H�{�4�{[t �������{�.]�:�|I�c,�7gt5�� ݭS����W�僲�c� �&��>�{�۠W]$�
'/,!IOQ旗���3���8�t	�����]sǫlq����U)�����0M�Mo� ��ɗV�O)5^݇�=ѿߞ��O�M�`�}CK�Ug�s�����VRW�KT��,@��)���M��$5���vv|hk9}9��}O��cUG$+�������~繚�H$A���3�����^��?=;��OΉەc.��f
���G�
cCDS�M�fyGY^�v�P��;�C�C�7���JN�s
��d�yf��_\�fn�LiUy�3�zM� �z�<���{����l�n�L�i�O��n�$�~T�aT{���{g�O'�&��Ʈ�8�淽������f]��hg	Y(�>��=��A�M��������c�$s��F������;�ٷ��Y�|��@߱P��O{=�3�Y�j:τ$�P^`�IN�s����̰cv-�ߧf��x3�o�7Ow8og�;�����imR&������[�#��y�N�g�-����*u�&]�{=�%j��5���>�\ޤ>�(��lU��_�]���СB�z�C�R ee�tE*Vp[���ΒT�#������5W��@P�~�T*>�'@P�}�i/O7J*'�wwW�+��&*�~�:� ���գ\�,^��Y�Ǿ6���eJ��m��5�覱ʺ�D����kڻ8��mi2�$Ѻ����:!�L�lnu	���ґ�ï'��o�����5��F)(�Y-�_/_w��)>S��5B��HP_���=��t����=���A�3��&�(��B��J�4~�n��=�74)�[֜��H� >��t��{�t9!w����w7'}W�^���=^���K�Wuc+�=9�{s�6�A��j���7���,���k�ϵ{{��
��6�V?f2��H�P�N�,	����dUVA�(6�&�t'b��=���v�0yu`�
�{4�}�M���>;h��MQ������OCv�*�	j������o��s_b9�{��h�ש�u3�gā5�ۤ��sl�D��g.���5����`��e�u���.�{4�H����	�wÝ�s\�C��W���K�������Z��W,��ǋ��W�__P&Ӝ��}�9+�yj�CNv��:F�����̊�Y�P�5����Ϸۿ=w�Q��F��ڵ���16�Oo3���s�7Xj�\���$:I�7�~0��>��D9W���*�g5:������3�;��nG�rp�1���u��7k���֌s��~�'��U�i]O�=7A�����A&-�VW�Mk�w��+�۠(
����@|�	��G�2�������A>�b�����n��~�@�M핽�#�L�J�JѲ�����	>;����6�O-�UU�#��D;��g�ށ+0Y�f��φ��j�o��{���5:��>����{���R������z��6r���X�  N{Νvv�7v�ע~�9S�y�@P����|<����b���ֳ�w_��[�����^k�����L�훅:�L�`�b�u&.� *��Ӌ�gK��Wp,l����[6�5�h�ي�&��k��!qe�l��2�ѱ�\<�&�����O�]����f��v��&��}Z�[P�v�gvsî�m�u�.���Nz�4F���tjm�q���mۊ�ۺ���ُ[ay]�@{v�Nr8�wqю��v�q��wd�=�ܞm�nbQ��n6��Gd�3�9B�v�mv�ω͋t��b�]�5��\�o����w��"G�y	(�@��cTA��սrQ��V�=dc^u�ָ㜔�F�D$U���sp~����ٟa�G�zn����v-|�����A�3��$,R��YF���5��ѣ��[��|[T�>��f쿺o�@󏲼����7�W��A x`���
�9  �M�LPA���'�e�v�P �ߖQ�����\L� ��hd}���2��(�t��A��L���k�����܊��zj�{�"�A�Q�v3���n���>~��/����U�؀���$���t}�M�����׽������x�{hĪ��@egv���̼���;Jԍ�Oo�=ډA��}y�����j{��@}�{�t��K�ݽ��ꦛ[��ى7�r
29��2����F��dgX5w��~�s��g�^CW�r��k���M];g6��^>���{~���� 0����bc��o�����[���f�������U�����(y��ӡ�{�`|$W������f?���QG�2�m�Z���b��nz��
���=����$�7d��M{��b���X�ǢN�k�j�~�*R�x�a@��� ��7L}�������[po�� >���萡�]�A6a�ߣ�� y�J���V����lt�{�� }��-��V���VI��V��c�c�<1�	v4���¦�rݷ��3n��`; �FՕM���Kt�*��W�~���O���:��s~�6�� ��5�#����?5ν��� ���̣F����O�ޡo��g]�����4�H$G�5�י贝�t���=.{k|� �&��QWwC w�ۤ�I��� �z�a�Sn���Q�	���>rmnzRƪ�񐔋o�p*&�'.���F��5J�*�/��.:�����U}�޼�b�8H�M��;��g�3h�J�eW[�{��������(UB��}@P{�VE;м�_*��ٝ��v�tu��]MHǹ���`�
�����=5�F�7_E����ϰ���ޛ����7��>��v�7�f�5�ۧ3�9��v:��x8�g���9�]n�jn�]{o��4�#j���7��cP���HP G����G\\�ת�۾�7�5�g��3����@*��V�|��]��,>+�fkZ��i�lU�e<~�'�\Hw��S�E���4k/���'��n{͊�w�>}� �w~�k�*�y�*_��o�;1٫h��f]/����jz����)��77�:��sqۡ�8�!5���Q~�^��<�b�3��w�l��W�5�6����J$�gn;w�vf$o��
�B�C�'l��{��=�Z�C��A���=y�x���7;� ��J�|+r�<w�	��́@}��7^���J�J�u�2kl�e��^��q:l���n�n�ӫ���7[5(��z���<Bz%F��wg�Vw�$���t(}�{���?xo���
�s) ��Η��vU�@����Q{�Q'mT�f?TN�a���H{��� ����.�a����|�i�z#����8o)^�:�{|�S�'Vߩ�+��Vߵ��}�b����$߷�D����YO���MgJ�Z��t���� O%�� W�˛�(W7�ur��sfx��*�Z�o��j=J݉�Ybק������o3�K���M�9Ө��PMZ�  �o��$$ I���%�)$$ I�$$ I@B��$ I����%��B��$ I�$$ I���%�	!!K����	.��$�	!J�HH@��	!!K�$��	/�$��HH@��I!!K�H@��B���PVI��c�H������@���y�d���O���                 
  X  ѭ h��  ��PP  UU QA�n�D�J�
�QB�JAB���AJ��%Q	
�(*��� �*
�*�����Eoc��_w�\w���n�Ӓ�c���Qקi���
| ���5�Ǐt��l=P����A�`Z&��Q"���
�R��
�Sω����ݍ�kT���){�;�t�_Fv���[���F��I` la�����	�t���)ѡ �(��y t	��� ݀&�lm�aY��@/�y��J�w�;>��4{���	�zE�<�h9� {0lE��E�UY�ۧ�(I���_`}[�>���^��:t�k��!��/xY��\ㅽ�=��K�$o��}�E))H���5lh��+��Н�FC�w�A��v=:��
 {� �}��Y�`i���݇.�w����5�^���^� � |$�U�R�(|}��K���^��W��������FE�T��R�=Wl����B�� ��Ze/n}R�vy�Wl�{j<ܜ�]��:oZ�f����e|      OL���(�4�`  L4Њ~�$�J��` #   #L5?F�M2�* 1 ��  ��UJOF�� �   T�D�2��4�      &� )#Bb22���P�=M�I��>���zϯ[>�~�|�y�^>��~�N��!H@4I�P��P��!!! ������	! ��  $�d�q��H@7${��?�?�?��?��w�P�AQA$����0�a�$���0��%`�	! �!���-�Y��A?���>���DH@:��;����\�p�K������s���?�~�ἅ
X$_G�y��>O���)�.�֎��˭��7�:?�<�̥{_Bo�����lk"琥�1s��iYn����o�W�H�i���֟����H���a�����R�����Y\(���Y{�އb��ni�c5��w4	1��������9��t}�g�ۋ��p6��b��x�vwcB�E�<9S{�N��z�Y� tD$`��H�����X�T��6<���5�P횕�A�V�܃D���@ 7�c�K��f56Y��V;F.��|�8��;-#�3BSx���!����vZU[�ƎDic�\b>,0��6�zdA�8��H]���b�@ˋ��iY������]��.�+�w�����l���'Ձ�����ۗ{N\��{��bY5�r~��t���k�LU�d�\݄�N�ڵFz��at$1�i�Y;��5���ר���\�_�y��4i��-�aS�����;F[3m]�uP��	�x&��Lc��S;�A!���^9�qq��*ܢMt���'�ś ��9X����o]��\�\G�Nx��n�s�sغŃ�k�tٜ.P��g1����Dnŉ�ይȸ��A���6�r�����C�j;�Jg�fo!5m=��-ݽH���l����K���&كq�"����6���s(őI�!h��W'�~N^��:���7���+��jÅ���S��ϑⵛ�A�
��pyn*���:����'���zd�N�/4�!gl�S�[���Pb�nr�{u��i�e��d�-}���kL��y�ut:.�ǖ���2�:�~����2����p�sk��y��4�zMa�oNk5��|�n���ކ䜥쓱Y�`��b�2BlYY�spc�X�"�DS1n+I����ӻK�.�b����]��u���'�`h3vb��5������囙." �6�q�T�#(��j��Y۲Mz[΂hK���r�Meۋt)�؞\�vv0�]�Ԫ1�]�Mҍ�j0X�,�Y�8U�nl裛�m眠bl�)+:���zpQ��MS 팹�>	�o�3��tLO��Y��%�u��9q$�LT�͙��q�f<4�'![���ь4x_�Atz�ᩀ�Ѡp-�Tm�5^������C��mK�vP�Q'�`]g�oc��9���ߎ��"��܇n���_l_h�7{�f���a�o�]�q�V��������Jqʥ9�X7D0N�$� �X��\;��$��?�Q�1u	5i<�q���qJ���l���=k��Oz�%7l(��f�WG��ܜ-d���"u�5����� �]kn�Y� ��;J�^H7��D�yZ�2̝��e�N�nV'](p���v��k9B���X������[^�9����+5X2=�g��'�sl�˲���4��lZ0�"�,�{/)�D������5�r�[��k�]	�귥*C�Q]�1BQ`��r�&��f����=7�D�ձu�(�φ��G��"i�ri<���p����t((����#:-�}{�2��HgǤ<(v%�ԲU�AɅv����iB�]P3ow,��@�{OB��~c$l]<����9h/d%�tM|��+ur�QI��q�Ud�H�{�ع����@�(�v�<�=�wc�LD����!<=i;c9O�o#�#��E恤v���n&�3m�u	LbY�І_����v��:,��"	�Z4��f;^���;6���c��ϧ�s�6���g�������z&���m����(5��;Oh] ە�看��q�:3]�9�m�{'57s�|�����>x:*�M��vշCp$/7m%��=wx``)<e�N�ױ�a+bN���+�	"4��q�
��X^l�c�)z"�f�ݩ�s�.�����8b�cfqG���n�5Y}J�Av��r�w�8C��k�80�e(]����u����ir��g\[��)[Yu�����܃Ii�t7���I�>����HV�����R�ڙ`XN�r����t������d�f�6^r�D�'n����H�%�;���V��Ӈ
�,�YU�J��w7�@ kѻ��l�S�q�ቭɚ;����ft�{cY����@(7��g'z�����P��T�.�w0���<;��>0]��4�Ր����%O�����m�Bw
#܄�w��CGFY׍0�&αԻϻ�F�^�d2��BP@���7�P6�uL�,/u:v�����K�c��3�7Sݘ�qT���cyy�FDw=Ȝ x�GL�YS��v�v���AW',���qEq�wv�.l�p��F;�np(H*B���R���91�1���4c+a����;Y�7DI������Wي����ӓ<�U%괔.];��z�R ��n��=i��2�����
z�D��Ӽu�P�pN��4v�eG�`�v�Z�Z����[z,sb�Iش���ؾAE��e��7�A�Q�̒��
�ڻ.�S�R�U�=+l���=oQ�!5)�w���{	۝75�)� T�I'��ֹ(��Z�5"�Z���PwE͌�9������M.D'·u܍�ݎU�e����-k�D��6��{#Qh�oF��ϳ�\
h犩������XY���C�*�@���f�Җ�����;qvp�!�^4Ƒ��m;�3P��f͸��L�y�V�o�d�\�Ex>�yG�gnv�}���aU�7!c78�V�٨�@����l��2����c��JBrcZ6� Ƴzm��p��:q��@�]Ɯ�S�����3xƥ�/k���\��Kq\��V���wp7�;��[8��xhi�6����@5o���jLw6Ot�fv.@��sn�5v�������ˈ^N�:��l�G�y��0vm\�0����7�`��Dv��^�<�/Ġ�ꙋ:�Poeߕ	�Rei'��Ѣp���f��.�4h�vW�Y����� ��%����;i�)z�o�,�	Ek�݂:���NE�]�f����)�N�̦5������T�):^���'��`�8ʪy���E�.�#xw�y���I��;Mu�������������ۃl����+ͣ��<Q�=���٭�P���~�\���y��6k�w������vL�~�v�y`P�m��V]ZA���u^�r�*��G>���My�^�0�11��m�V�I��ڎT�}C��zN�j7�n��^K���͡윘��dC9�`��&)>�lעm�r:o@�1�d&*��І\U+owS�6:��.���3�3�r�Zy�����hʠ��Q�s����΁��=W���4���j���U��F#�@K��q��Tz֦��tТAǻY�t���'k�И�9�:�=s��n82Ⱥb�n��cMvaӨ�X�hɏN��d����C	�y8���`�%���&� 7�� 4��d9����^nB�]����n0)�!�uٕ���� L���ITvjfC�Ww��9�za����S�w��Im�m]�7t,�[�5�X������^q'��v�.�w�k4�����K���
[�w���=݌��T�ʷ��f��Q��k8y�z1so`Z��B�8���9�ۗ��1�'��V\��ά�@���ݵ�rzG/�t�{@�qt�Κ��ɣ4tb0l�f�1��yX�"��|�ywN��ƃ�T[�"18�x����s�����<ðˢ�6,O�q��5BˀY��,�|<?�?��D;�(���:�N`��>�>G�<Ϗ@Nm�ӫL�G��q���==Ԅ�I Ad$P(@�@����H�H� � � AB���H��$� �(H`!$ � "��� �@+! ���(@�!
��! V�B,	�H������,@Y ���!%H��H�$Y$E BAI 
��a!��� V ��I$�@�$�`� !O����3��O������>����H��I		�	���l����$'�C��T����~a��j�Ĩ�_���1�T�i�l� ��0�u��ע��v,䇓"<���6�4Ov��.��[q�ݧ�U�q��/=����_�O#/3E���>K#6�ւ.�K"61�yX���h��k���"b����h���\� M{T�y�/+��?k�<�j�.>F�{q�n`ۢ�z'�2Y��f�G�-�٣�<��_j=�d[���7��j���Þ�1=�3���t���#���.�r�c���D+Ø�m�st�l�{/���	z�?d��p�\΃��fڸ���v-�8{XX���Q��LA@���C��^6h�jp"�є���p��I��1�;خ������W���t���5��� �ԟ{�2��w���|�N�ob��v��
]�F�Ɨܝ�b��bb����"Wk(�Z8v���z���U���[
�P�xfv5l��8?{%�_��<z����Nw1{�Fo���o�{Ƚ�~��W�y�������yӭ����޽X�����t�R��lD�.����p#��ڈ5������t�6V�,ޢ�q����7�F���U��xy�-L�۱{w�ј�1�8���ﭲ�2O.�<���6�*�F�m����a���7�]8��7A��o8[gɧ�Q�x���^T��֘[�=�d^�h�ݤ��r���3Nj�k}�E�2���q�Nn�x���@a�]�� �HR/�d��ｭ��'��o�W1;�K�w��{َi�=���$��˻��9�oJ�΂o�� vhm�?+�9���vw��}n,X�N�zQ�ר����[�n���wv��mʦ#^́���3Ų��xeL����5��5��ba��x�or��{}��,[�ul�u��s�O���أΛs����c,u���;�	dȨ�������a{�>y�C���9�*t���7��۸���[�-<�pCtBsa"��jz2�xq�;G�t�O��B�g��aǢ�C�����1F�ĕ+(Ѕ��9I��4�8b�u2�D𖍣�,�<���&zW�n�A�$���u�C'�1��r>CH�N	�j<^�|�ȕ�2�s�z�8�snmÀx�R���ny�"�v�����O���,=�a��]2\~W�״�A���!hPbܹ�REE	9��פ���Q���m�3���V���N<����\���� �ጭ�`-�����v��/{�eū�-X̑��]�Y"Z�����-�ꁌ�N�B�����y����z�R��M�`Q��Iiru�����r��u�f)���i��Is�Q;�wol����3Y܏��Ȟa�0�x��c�L{�{�kW�#��&E��I{��b�x���Zr}�����>�t\ٚ���h�COzۺ}�]�c�C�����I���E\�*-����zQhE�Z�;�i�kr�h�h�@��H�ǻ��a{�^������W �O��.��w�����y	{k_,�Ҽ����F�9��\�����;�e�`zw���e��[ϟ3�އ�}=}RSp���0yD�e��U�m[8��i��Q���u���9�Ո�lV5�ވw���"͸3�^ܡ�<L�svP�,�K�E��s��_;<�՜ ~��oJF	��u-�T�bמM�Ie��E�2�`a����,�&��]���;���Η[7���w4W�nW�������$F��6)��r����/}ӛ �]�S��RR޾���o"t�T�ҠeR��>QO.:3oa��С�N�,����Y۶��it�+`Q=O'���̞������;�p��^�׷#an)�1$P=�\������u��qv�=���K�9��c�7��>��,���k����}fyĦ�77���)�uh����Fy$�%�M;�=Oɞ*2@��1����0�l�^ݝ|��D;���{�����FG��"�Ĳ�-4'v.�^�7bli��×+Y���[{b��D}�Oxv/yߗ* � :y=��z:6�s��	⧖��~�>��i�9�}�vG�c4�&i��z �V�^m�m�������=�n���L%�,����	�Ž����_k����ǟp��{�c���Vn�.n�͙f{۽E~^r]cz�I�6{��ђ���7s��S`����Rwk�O��P3֑yPnV����:�������e�g��Τ�e�޲J�.�Q*.�R|���Kzq�@�z���+�	�p]�y-\�N̈́i�#�w���ԯvl��A�=�7�9����>�`�=��K�]����z�����zߗ9��D���X�A8m:3���\�c��Do�~B���|<�ܰL���`=6v��%�Kۛ��=٥eJ,��-Z��� ��H��S&�۞ↇ�8�ò-��'v
� �l��[�������m�|Gı�SV���+�Q�o��=ޑ����uA��pk>��~~hI�a�ݔ絇q�-�!Y�ָh���i�������0��sI'=�.����Y{/����wx�ӯѾ�Pm�V�]��Nvj&i�fO0��y����d�^�I�����ٓ���������ݷa�x�M�E�=ۇ���Q���l�xk�SL���������S�{ Y�Mh(��h �,'X�N�i�:��w�ܫv��W8_N�8�gޣ��ec����z���{���f�0��Y���͡_�WA����"+�;̏ZBr����E���ᯰ�e؋�ylW.Q��+��}�(=<�2����
2�^5�-�q��E�Z�=P,;̍�M"E�pY�%wLmT����c��S}��䬡w/A{{;��7"�1���r�j459#B��4o�����{l�˻�΅�8.���Z�v`L��N��'�~�[�g)|֥�w�Ѿ��x����m�\U��"�ݸy�Zނ��&NdO���N7���]$f�8J����@���x)��?�{[�s��=�9܏W�=�s��0��k�x&��b��������u��`�#b�QS����,tp;��y��`�c�m�����>�j;�+ey4@�Q���̀f�&j<p;q��� �vn6O"�O^��k՞یs"��2��������i��[���~�͞�m���bl&CY#N�n����X*+#UH�)��� `��/<%`�n��~=��bwdlTBp`ך32#M��Т��no|��e�å���S��^�'��ҳ���(��j�س�Y��6d	��sث�t`<��)�2 ����P�����s��(܇O�p۝��7$�˓����8���{��`�X�9��|9tEw��v��]k��'ww�u�L��7Ԭ��K��<��Q�g4�h괿xι�.��7���JjZ����J�v�`���e}�d{�	��@"�DF�{�Fy�w�2����o�(���j�x�}_h�=R^�v��*�����D�wB�ۗ.��bmk�Op���NlF6.�2����.��wQ���.g6�L��kA�P�a�eF5{yF`��(S�Jc5����a��"&v��J��g�ވ�3�Z.���J�v�a���b,��zc�Յ����v�^ѹH)���=�Rݛ�8��`2'pl�a�R�W���)�ʜ�j�-��VEV?Yr�M�L� �gh^x�N���Lozy� �6�f���(s}��;�P�3�F|6����9؇?>~�okã+�2H0�4|����.���^�
懦Nஉp�Tbq��0G�5���vЎ���Ny�[�5|������!��ߒC���3� �/�2+&��qu��ܯ��d��&��{��d�/�O��Y3�H�s�o{�o�Z��k۾�7�\e�>#��B3ͣ��AUM�'v�j�׫��'9��
nݞ��`옡��ʗ�T�]�{2F_����xx �,"���t�`Q���0���Ӗ�&�;�_�GQFYyq�[Ա������̝����i�'�Nv��	��f4Sx���l��fzy�s���{�\&���Ź�@*�pǉ�X�q��5�Ό�][��D�Ɂ�����r�nr�<qv��^N]7��
耷J;��g��a�nC�M�����\/n���4Y�2Q��8�l1�"tZ���sN�{:Ě�$a��f�*���C6��U�kl��4����	i��,+�L.��0]�J\��`�+�����O����}�:HQ��� ;�Z*M�;�m���Aa�a��s��P��ÓaW��3��i�;�6&z<O�j�2Ɇ�q��д�e@,�X>9�p�;q]0��E�� .���7EFhq,�Ɖ�4P)�.��yf�������6�#��+�k:7&�a����uh�M��/���m��ض� ��6�.'�-�J�ں^�gs�<�{��@��1�z�J�A�ܮ�-4�"kxJ8��6ly��]F4r<�aרJ�!k`��;�1q��&7�S�k�\VossKh��g ��/
�����u<��O)`ݶ FqU����Q�K�^���{�IVbw��X1P��͐�J�k�4��P�k*�![Ml$�+ŷ)賴d�yѮ
V�t�*��d;!��L��p6xψ��:�8-Ї���]�p;����ŉd��$ꮺ}X��[���`�È�"�6h]j����u=&�t��+=�vW��Wpq�a���f��<Ž%��u��&�GX�e�髅�Ai����זڳ���]�P��pr��g���8�Lm��X����H��ܼ�o=���ey�Vt{t6�n8���
�mi�����4��̓�V}��m!�;�AщL����r]��sٻ���y�����-a�ʑ0�K��<�z��h�m�++����$����n�wcG�:{gq#�p=��t���]�ݞyIi��������M���ն���	l$#���b�}��\G*�8�r��&��rJE�ɋ�tt�g������3����X�P㡌0
��$��/Jx}�ٞ��ۚ�<�<�V��g��+׸�ʏ���rsd�*u�n^�gv�=�=� ㅠ�4]H:�쒮�L������s�%��s���9�Ϡ�%=q�v9��Z�s���u-�{�{��1V�+��/j{��ۢ�m͔��Lq���3j$V!����ۆֹ�kt�w��,nB���p%���0�D��=�5۳{bȺ�:��b%H&�&�����К.,jx�S�H���9�"5��p)���l�+����u���F��u��l�@"A�ķX7m����Խ&W,\�=ZB�=쎷7��:���-�P��&-cV��[�f�� ��v�(W-����p�n4��XSEց
r�K�2q�dۃ�۞aM�-�����GZ�6����*9����s%�MƞD�ˇ^��Ճ5�Oc�Lg��������o&�2&74�g�r���iCFf$a4��l�6�NT1���Dы깋n��.����Ր�琳BcYq����Z�f���\:k^φ��ݹ�6��؛g8"� I��*X�Sk��p��\�9FM�p-�c�w���s�t+����Od|e܊��NI��45$%��lVås��5eA۫Nxݎ:�p]`Ui7:�3@D��bkl �`*63<!X�9���,kK�,�ٝ�a۰lt��B)�\@�!���1Og��a�{��G/V��ӻF��5��Z���̴4�!.R[k�e�T�%+jC���Qq0�r.��c9k@�-N��DV��#��)ql�Ҩ12����	���`�˔4cG�!hhB���e�	��+]M�3�k��.J��A���T���Pb[Q���v�����(�H��h��Z�d�W����`��=T�]x0PW>m�0	k)�JF3HFV`�һP�9v��2$fCt��k�d�
��=k�Y�g!��ݪ����[���ۍ�@��m���s�m�O�M��r��뵍�S��i�3�Gmp��ױ�p�4P�`K����
A$���Y���!Ҵ�Ѧ��,	���M��E�y�[���1��)-�r�͒�Cv���]�:L�wf�',D\qp�A�u�k�_)������l�MY*�(١b6i�9�.y�Բ�uv�\�-�v�6$l�jU�y��p��� G^f�,4�+��m��0-�6xM��F(���\�p�t9:�Wuݱ^����ؙ�vl�	�]��xQ�+\G<����oO;�0#�`�^p`4f�s�z �8KE�x1�0q���jbԶJ$�`QFnc!�F�1urY��IU�D���S�5��i��F�n����%�lL{%��oE�0a��Kִ�/`_k[����S\i�7��f\���b���ܙ�M^3qつX��n��͌X��@��Z�Q�:Z�������UUUUUUJ�UUUUUU:刢��..�8��r��K�W�];cx�uI�;t�8d醇V����Y/oqg��'�n����Zuŵ�T#�n�m�fc��IT���`M���5%�-u��f�+�)f�&�+5��
$@�
F,�F�5�Y�fؐ��{+�Z��Y��ݥc��J��5��5��. ��U�p�:�0`5�ٲ��Z���R���/@U f vͅ�	5c</nر/,Ř�ź��`�U6�M�9㶴�#�d�҉c��"G�N۹z1�����5�j��fjͲ�_��x�ug�9b0X��
DH�:`V@U���"�.Y
 �*EP����H���T�ˈcR�d�.3�X��ƹ���CL�2#�YY&"�Ԙۻ��R-��PDP�I���H�l�AJ�B�d�Q1M���*,��`���Lf2b�Q��(����T�HIV�DUKjE��dHp�`�m�Q`�0QH,"�:h�-�AF�
¡ib�PX[E���YPX��A`,�+P*E��P��C�P��,�E��H("�*�4�VZ��;ݿ���gɫ�ј�YjyK1�P��ɮ�cƷ���1�6�N�<Z�J����x<�Q/f����8P�������Y��gZw6�@9�p���ާɽv�=s��Lr�j��w3�Xږ�k0�fͩ���+����vK۲�<n_-�c�xunN_W\�י��ֵ�q*M�,�n��;s�q�8�:H���ۋk,�+QS�͋��A��3�b�0rю!�n׈X�t�e{/��XX�XP�^�ShF],cM2MP�Lnjmb�Q�M�88�����y�n	�gl���`.��Xb��6�f7_ü?>gx5vx�\�����ts����8�6d�gig���yZ;K����u��m���1�/>n�*�m�6nMX[��gJ��P�
 bb�1\rq��b��v+���ہ�(Y�41��5H�5�Me�����d��<;�n��tyQd4e���z�üpWD�um�0���p�"�wE��ɭ����b��Z�ㄧ�ћ<^��5�SV�{vMa�n�1����C�9v���<c�k���ݼtƎ0I'&E��bh^iKy������Ϟ˜.�_<9@��6�MK14��
`�Юxy���x6�*!��{L�e9�܏����˃��˅�G�s�<��|	�{;��s� a�*������vߗ�r�l?�.��Z��W���w�:�B�&r�B��4�"n_�E�*�� G���� !�����>�)�u	����� 9�/Vc��G���䁖qw�ܕvfu̽�۴���j��	f�LFv3�G
o�P
��]�/d���� ݐܕ�ι��������u`9�c���p&�^L&P�mBot���O}3��� ��J�^WESSs��pB��tDl�������'�ߜV�7f>����Cv�sJ�lE�'�Qɨ\�x��c6�lfr$���E�O&,��nX:wu�eϪ�O^GH2(	�Z�ۨHG�f'�K���'m(�6��=뻛۰�7Z�|g4�I�T���M% ��U!A7����R�q��k�U8�O�%��2�#-e�.Ź\U���B��씉!�&}��yq{=M�Ԓ ��+±k*IW�9p2�}�~����T.�{�_	�qC�m�8bK�l7` j�Q%nq��<A�s�`l]�,�NU�q��"%�nDF�7�\��||�W�ބc�DB�aĭ����K>�=4�p�f}���~@L�4F�0�1��	�E���ܠm��n� O�mw�Ф[�j�ʘ�fTe{%�sr]8e�������RiȽ���P��C����� ��$m�'i����I��&ig/X3Ј7�#VT]<kѹ=��QP��k}�g3y]�>�j ݟt�&�}U��|���*��[�� !wsXC	2[�FT@�S-�#gr\M�ڛ��$*ѕd+Qo"r�*��h�D�@wZ74;��!f�T���k�� 4���&��愢��؅	��YP�t.,�tKL�Z�;���a$b=9	��"}w�N�m)��Fp��gd��M:Ռ��N]�d�I=�m��oRR�7`�T4�l��ΦF��}���p�E��Q~=�YRJ�E��g��. ;o�O��O�=UV��wR$�8�?7j�ê/X;Fe���Ak�\a�f����
����瞪Q����|[�?/�h0�|D^��[AxvST��ۨb�1�CX67�ehVݘ6U���?>tGt@ڶ��k���8{g׹ة�xG���t�,h�mD�b��cefP�z�װv�Y9�]j�L�����Jr󧱆�H�ڎ,�6��7e��ڎ)�ΖЭLF��3���%:�T#���ۚ��
� =�(G_�glZ�Uέ� G7�YC�NA�|i��NV7@���<�@H�^��c��QRz���F+�n��	;6���!] w	P�s�����bZ��҈#1-��Q�d5M���rI*�kOڧu��mR ��jF$�f�b�q�=��pKi���,�Ζ\F��͹�������x��͓��y�����Ļ�[���a*�$B��+y&N����;�
��34�Od�����t�	�U�\�,=��.����OE�.��r�' ���3�'Wڿq��e��e��.mWU9U\�3<��U���d����v��;�0����7�(�DΩ<��{OTzf='��Y���f	H'��y��5��GL�UM*��ʒW4Wn|k� ��2�w�!�u��p^U�K�9���|��r ��O����뛍��t�\Y �M��a(�XV־�r\�c��C}��뺶����_��!��-��w�Y53�Z��N�A��	��U\1	ߧ�:o��׹��` �?b���@��<O	�Ts���M$�f�I.�Ӏ�{���z�_\���a��sqt�ȴg��46��w�P�|:R�:�� �B°�LH/1<��zI:�*�`2.�r���ʤ �8����}���U�.�ҡ��8�7/�x�܊&�D*Uzu`��||Z����Nb�[2���k����٘�x��b�w���eүA1�efʗ;�١;͆rJ�l���^E�va/w�@n z.p�bv
1ʁL��뮵:���.�r�s����x8M���bd�5��S�vZI��	�@������^�V-��$��D�z�)��t�w*����s��j"��-^U���n�:�p����B���w;����>v({�qo7ښ�� Ek���9�����YΦ�=���Q'� ��][�E�
0�<�����p*���g��mY���m�\)�{�z�����x���w�::漢ơg��i��%en�x�K�v��;5�\.�&�]�h�0qKS��LS�%,[q��[�aRh��B�\�cU�p;V�4\���+rf G3�l���:x8�)�1ۤ��7\]qj�F��Z�ƻ(��j���TvS]_���<Cc^y��|�8|w�K�S��t�q�p�`Xp�s@�c�d�k��Qaw�F�0�.�_":�^���7#�y�e�G�G���X.�C�ݪ�ጨ���A����v�$�Gٜ��d�*��{ 1!I(�\��I�*����zE�H����}��EP�9F{�X8��yM���`�#���4��_#`Ë�Ԁ$��I� ��pӤ}�`)Y���@���bGl�FSgi��Ùv��1�e(21��:�Y<�Zst� �E@g�U��S+��Ζ�*%$��r�0�8H�dpHӽ�� dT���w����VS���|d<��T�F���V^��wiW��ƒs^"�/�g,tOW6H#����{��޻������W:ѳQ�u�ͻl/��[��|�'��C��]�v �qFD�V9��X`�7 /%�-���2D/T���&�<��p܂*��{y<�z>�(N2a΋��D�!������|�:k�]�LD�_��^���p�.�ڃ:��P�d`ipz^������ϑ����e=Mu�p-%�d=�(zۻ�zBV��p���o���5�$��0��A��"V��"w[𵱛����q^=���BE���I��8)����1�2o����ȶF��g��t�E�=�ӥ��j�'/P����?i�����]��G�[Q:w��#i��`�=}���n�(jњf.���7V�R���P����rx��� P�����:���=E;7��F;�}|7������>L��{�f�Q��.a��Z7kw9�<s��0M�ݞ��m]��m��i��jK�B�4ζ��+��:�p{�y�OB�W�]��gv�P��x���+��nY񇽐���0�)��~���>C����	���-�l:��<>ޖ /O� ��$�A`,&%@�Pb!(�16��X�`bE��a+
��J�Q	m�`,��+X�U��:�$ED`"��R�6�Rn�R#�������U��D`(�$�TD@XT�e��U�#$�Da��M0���(�E�� �pq��|+�tǿi���o&�u@��h]X D���C���_�(/Y��������S���!�$��
I}Ă�$��nk��{�B"T7�fH�����77++176oOAi'~��Hw���[ ��D����>�c�a�ζA�zXaj@��ԁ��*{�us��0�8��A�M�H4�w�м����i��
=�o0��Sv��#<A&v��$�Ȱ"�`J�x�@r��j֛b����2��rj$=���y��
X���G��ۡ�Z�h���x�ܐ'ăӔ�,��U���zs$��j���liV°�,�1�[���;�oe���ē�UɟwG�oV��+�S^�m�M�7|^�i'5�*���n����b ���Y��o�fJ��,][�CI����/oV���)��IVߴx��4j֟���='ލ, F��d��Oe�<��"��#��ԙ��P�R+�p=��!�͵MV����Rv/�g��:7ު �g��9���ͭ�1;��db7��V��D���ٮ��n\10�w"��sn��ge#.Q����X�[9�$e��,RmV1�.nX%1]���h�Va�j�s.�U�CLe����,B���JjM��ۮ���퉩H�v�)G"��3��P�Q	��w�q1�m��^���i I�ʡN�9=�a�W.��n Yd[<�p���~����z��	9P�>$ws��.��v�w$��1�����t�|n������b�"�
����}�HT��\�$v���p�+�����%�a�К��A=��1��������ݝ�!��G{e'C��Ϫ���t+��س#��V�]�ϳ�ͳ�+�v�A�mPwNs7��)� �}̀HU����m���)��)�8�6��j)n���-[x��	��#��CZv#6S8^unwPZ�L%(1�9���d����0L]^ս��p*d���	�n}�l0	3\���R���$�^f�Xf���Q'TDЇk-,ɛD�Z��H��>;��u4�#F��Q����$ܓ��d�Ԙ>����ƹ�����bw�N\�ᑌ�j�1�k�a����;��~��gMk��O�sapZ��m�NP����IBEQ��K�nyR�I9��������FX�L��r/oXQ���6�+�;��]�e;ʛnE\|{��6I{��re��܏���\헱�2��AwPd��B&��3	�nGu��G�l�<$ƶs! H9�����s]�$��}�ΎFN��!Φ�1�y�]��=�'�_��
|�ϭB�k�����f�(��i�N!��I��P�:�#z<�v�M���j&����A���$�8�\��<T�wv�IP�����l��85��JH�����)7��&WK�3Ё_sV$[-�܍��`�a�#�z�33�k�ѽ���K��lH��ye抜kv.���ilh�U{J�څj�3|��L�FIVNW�?�����?���CI8M�����ˡ����D�l27u��멜�YL�Cd�oS�U��)ƪi�9���a�]��I.yI���jSD�P(�^�ps(b�S�E�nWe�e�v �S��a���,�w)��Z�!�P���':�"�$�L����d�M��P���{�3�UUlH$�jd�Dֶ'vʪ��"pHЛp܌��A��fS�35��͒D��� �������a]�3163k���Y��b2b�3nj��ѭ��o`̮��~���3o4.���6V	��ֻv�;p;��GoQ�\]���fg579]�-��7c�ǝ̝��5�<]���k. ��\��zhೞ�H]-ݐ��hM��Jo'j���j�V��vkn%��sz�fcg��u�V�U��X�~y�ߎvj�w�O�ֶA�F�c���O�����s4�d�Np��|�%��H'���+�C���'�a�l\�1%N6#z=3V���I�`��5�
��q4&��a�<.mR�A���wk/4��Z�mrs%	AIG�m;�	Z����x	{ʡ��=�GLLDͤ�6ύpK���c��ʲ��t%ˆZy�ۆ�]���A��/�����Ot��bm'���$܍��.	��k���Yu.������x���~ܝ�d�����}�`z�
�͝�� {��s��I"��?~��M���1��*,D4����PdX���ڻ$�u���؈��
�/��l�!� Gu��9ݜD��(zd¶�U	�oĂOu�޵R�;1�L?o5ay��Q�]���ztj<��G3��zyΕ"��Q�+Vuc19#�1�.P|,�L�=�����_see�n��Z�+���>����/l'&v,���n-��VA3\���Z;��#E(��s�����fvV��7�Zh��ب�-�#cu��'!���<<�7n=�k�$}���͈�
u��&aX�	Φ�ְ3aˬ�p`߹�sb#$��S��ɋ�`�ws]m����W-)���~NٵcK�.d�Zr��;-���k��<6񶷿z���õ��H�{�bY����j|%*Ԓ?�_Qq���n����%�����Z�S��B�m�t7ma$MB�$%[�r�>�� �v���wa5э�l����[;sdf�g�ݰ���قryM�6�I���rl;C�fOY���e�q������c�v&�a�S�4~���=�_�|f��_�"8(i�ǜ�Co�dd����{��r`Ȭ_�C�wy��]m�+a�\��U�7X�W;Ͼ[=�՟�뷌!=�t��G=��Vz��T O��L*J!�P���9�v�u*��CI7��'����lƌ�z���I�p۟R=�~Ρ1c>3P���%U�n�;�cf>Z>� 3�T}�����^��\FΚ��l��z��f��g�m��^i ���$��d�wy���:�$n������H�9a�Ib��}^��]�@���-W;nM����P䛩>Sx��F�6����#65T��Yd��X.���:չ��8��_+���ӗy���L��'I݌�F��M���f��8���v���7�[�2_m�=�/Ç���V�Y<�20��w��9�^�z�I���k����j�8�BaeMH�sX�1w�y��Utݾ����t�^=v�ɪij��������ؚ��_�PУ꼧{}���ri�l�Bƛ�յQ�t����I�4��Ʋ�p;�;��A	�$��6�[5�C$���0lA;�\Ym�r���zz�POj�шsѯ۸W/4n=���i���e��.��׷w�z��-ʁ��qd��L���ޏ#�=|�ٻ��Xl���rv�èf�z�K���Öp��.|f��k�Yϧ��'z��ԇ"'6T��>�X
(�c=eUk
Ņ��Q���\B�aU�UEE����YR-`�5�֬2�dER,
�H�I1%dM0�H��d�]2T�0*HT����2��Bi	��n�	�J�@P�%ea�Xi���
�	STS
Ȫ��J�U@�] �+
�
�=y~}�6�!5c)�]��5�8�C0DIU�g-��n� ��[6�P�Ŷ���b�0kbd6�W�@�.B{��9j���H1�[����em��zS��J<˄�����N:M	Y�3!y�98�:s�Ž���o,�lTL7���ٰh�85��cR�l-z�q.W���X�i�����B$h��iJ닊Ć�j��t�`���d,�i&�	�']s>���\�-�febͰ�+B��`�p'�ݹ�S'#w-�ss9x�rYp�`�6�1cb+5��É�\�IItt�Wn����n2>�^w�;��:I�jcl6sp<�rN:�������+;��n8�y:�g�&䌧mo9
3E��#����J �,8�[����9�(�s:�C�E7\�//���dp;;]4�0���)f�h�n-�u���!.�:��:�rY9X9��Ӯ9�y�.��ڡ��C�	�M�Cip��̠�h�ϡ��&�v���}7�!p�S9ct%���[UUUUPk��n��5�ge��@�%ԋ�l��lCs Yh'i�V��q��ہT��%E�p~ܓ��9ʶĲ�����^v�;W&�ܱ�qu��lB�=�ǂ�˛[r���&<�v�k���n8�5�s�u���x����;bVZ5���t��8N~��s�~d 2Ce1PW.��Ղ�K.u������m/N�����	�ljۍCQ��9r���~A��i��!�GĂ����A#﹌��P1Ј5��&��} �H*y�j~�weF�U �][���s��dmӺ�g~ FgiP��`*^k��!_2W�{&�mҵ$�Ż�����,fs`�I݆��^D��B3D�	�	�ݵ��T��:�����I�v��ހ�ߟ|Ͽ,�ώ�+ʙİ��X�*��nfI�r�9��=˜9����H������w3����	�v����% ��%n�O�C��K��/}������6k�d����}��g�vdH��b��N�B���7����x.�_���P�E|f�hݫ"��~�C�$8� �� �m�K0J�`�;-�7�R�.6���yPox1Bs��U#�f���iQw):�̛M��T�;B̀���;��Y�;�2Ml"I���N�:��~o�ډeK[�p�f�.��jʰ����מ�g�V�SϽ�$��$�3[7�ON���`^@��r1���Ho�̬�Fn��!��n��w���gWQT����1�6��)\�u}��tF���܀w�7�U?�;�/�����4��E�#����w��Ef�������Ē{c˾��@;���8BJ�7
j{�H$
=�j�'3G���9��"	2�lLLT˞a�s���S쏂̸�fK����1��y#�46�:9r0�i+�,��j�9�u�C�=B��,˔��l�o-;xn��@D��lvhZ-�nh�b$�<�Fz3���D�z�$�rQ]1����� ��w[g�\��i��.�<�������cCp���4-�}9+��a�7c�>�I���;02�4�`�o$O�!�N�^ZQ�Eh�+�WV:5<w���b7�G�&��x �d�^����:�`-�$w�ٮ�9:�#��R�^��u�0U��K�����0�x�V-r3f��kǭ�O��ʠ{;(>������c#U������J(BJ=ݞBR{hܖ��mW�� �Yv�6�wmN#`��㻌0H��E�HZ���� ;{T�FkS���Q��sw���T��@��� Y�����<�)�Q������LΡT��n�Os~�Ё>';XV�5�3gg�����8.���緳�nڼ�vp���y=�t8ٚ= BK]��kL�)M�փM�a���9K]2u7(@R�����v` -8ې�U��ZݲA��mg���bq҆���k�q4�J�iE-��1e�
��dj17U�]T�Kd�]MY����棝�8��خyh�n�!�u�1��V��/�����Mt�*u�O��A>��4r��*m�˦��kT^U`ܜ�w�B��3=t �Y֢���A�;/qI���*L�!%�3� ��^f!B��(��D��7vhZ-�n�����Yʅ�K$m �[�?y�L�P$�Bl@܆����g�\�����B#bE��]*>�Ԝ`�:'xt��F܎]ۭi�)�ӂà�J*��_}�k�=q}�u׹�A�dtnX�'��p1�P��1��*��jy�M��J'$�m���ڥ�=Ӟ�Wqsǣ��x|�?e�}�r�o�ʅ9ƴZ�08!!�1	N���$��A����8�g[�s�>=Ò;NH����Y��ݕ@��� sr	z;i�s`�������L��'f��u���ϫ9�;�x��S}}�obQ�XB�ZЪ�U �f��u�Nl4���i ���B7*m�����#��|h-�4D�*�p�:��Y��?�����h��d�	*y2A���`ΐ�+.Պ����A�,�k��}��{9r{.ͺʒ������֑mțH�F��������	U�`���h�&!*��r�?lM��	̀���:�>S�!�6*L��9#����ĳ�i�r���� -��|UIjn��>m
�Tc#�����KD����]	r����y���ۆ�㹈0ERD�J��m���'�f8v�wj9Jݹ��{�8�+Ӂ�����+�������5L�U*�\����k��,�t��X��
8��6�\��r�}t�S� ;��GoF�IT���9b�9 ����C�v6%�S�k����=���_7�{� 
�B�b��1	T���$u|�7l^����<�33R�D��=�j�,.��3�Flr�0\4�H�?iģ�$��#�yu ���Q��u@�B�=͗��\�7#+���̜90I$9��㻭��Ùnai��9(M9��I��$wq��1U0,5M��A���gB�Ki�2������$�݈2Ntŀ�#[~�B9�!eu6O��uE�jre�X�o�$�k5y��^9�2����6��9`���V�B�0PK�(�ݛ��UF���\�xS�_{����0E�
~���)\/0�ҘQ�����<ɇ��5��ӻ7��^�I ����1Tֺ�(B]�)�jк�k1���$�4,[q0���+�5�U�X�r�юH��:�b�w6�iA�[-9b��7-������~O}���o������6]Y�j�����4��*AH)ǝ�@ܽ��y.fpbA`��N�
Cz�����4�^c��R�y��AH,�_}�b@H�$
����B��>ìd�ַsT���$� �y�!�IP9���n�gZ�Rӟ<�6�R��t0*uy:��&�$W���bFGDtg#4 �<��k�9m
���1��%B��{�m��|�<�:�]M2v��FT�ް�hw�L�Z�l��X<q�Ć�!K@�p�As{�p8H)�<�@m ��d1��T*J�<@��$�I����uk�u.�&��z�j��])�M5��y�]�ny �o�I=��e`���JʁD���`m��}��^9Hu-8�8�H6���_<�c��S�}��s6q�N�)�z�=���&"I|Zx��S�f���hj�b�i�v�7Z���Ym��B��L
�����K�U�� ~�����:I��°�,�{�c0�(�IS�>0�&�*Ad燐���<��H�ۼx�eى��x�
B����h0*u�y��q�@m8@�D
ʗ���P�J��a��O�	��2
l�>|,#�Pj��>�r��!Y(���43I �_x�F�mH)׾�����)��r���o\��F�.k\��'����h ���8��6�hs�������g=v°����40�(�@�p�&�R
AN��	��\����z�Ϟ��kxuWS8q����`���]\�{￳y���xrO��04�B�H[@�a���R
l��4�bN<{�@m��
�FJ�P8�4�l+���խ��a���� �{�W]?#y�|.|�+*�sǸi�������0�m!^z�y���8.��R�6pw��3�9@�a��Ι*AN�� ���aX2K�޺z�ݷ�]p���<N���׷=�����[7��))��(-	$^07�H$?_g��'��XS��|�1Ǎ�}n�x������ ��9g��j7]�c��=�B��X��;7��9�Uo�v\e�����<1]~����L��������d�����O����k|�VOe�����|;�xn��5��z7$�[�J��و����W8�����~���l�s��n���{U��Ca8w}�F�װi���17��]o�D{���ś�C�����j�	��W�U��U�ۀwBk6l�!{����-
��l�?��K�Fʔx�n^�·����2����h}尮��#��`�V����>�My���J��E%���+W����1Z���+b��F�1�-i����+D1�1��c�4���5���ֹ�h����ZV�<�n�[���W{1>��t'Q��_^`̍F�$n�� �LP��$Remf8�Q�1��*IY�T1�
\�b�$�m��8�ֵ���ED]j�2�
�ăZ11"��J�ҵ��Rn����$KaP�j�P�cb�"�#R
AE�jPĬ�2��.Pm5���\Ȱ���P�R(�̵`VJ��Zҋ�*@��-���j"�0*CH_�BC�3x��
��P9���I�l���<�{�i�7w^k�vc���p9��t�R�A@߽��B�`V�
�u����+*w�d+<��s�8�HhIP5�p��
�]�v�\֝kp�#
�����ɶV�p�1���M�y�6�XjB�O<� �� �C��!R
e���ʲ�k)	aKXQrm�p �B*p�N��/�4S| � ��i ���q�������܅H)9���a�M'���6ʐR
u�M��כ��1��k��-a��!R��w�<��y���4�R
AM��i6�Xw|�Vhd�T�^S���ǜa�Aa�tg��[nq ������T����f2VT��gl���~�,�#��&��79 't�i
�s܅t��{6xs��3�9NbN9����=�z����YY*{טlI�*J�XY�{�VT���������&�i�_F|^�5t+�3�>�5�7��Mbj�v���.���T�;^�|$�c'�+%eN����M�+�s/08ko�
�R
��8k�B��Z��g]��6��(�YS��!R
T<�0I���;4'/�Ң�+F,���N�4���nA�.b�������5�Z�0��O=�hm%��7��H(�S��Ѵ������ �y�I�B��̅H(���z]c����t��z�i�+8��/}xq')�{�BM�bJ�X^3�B��¤��2m����y�;��z����;i  X���pӡg�Y��qXq!m!K@�a���k���x�^r	�J VQ<β ��%@��0�Aa���߫m� ��M��{���a�AH,=���1 �
o�tm��� �^y�uק�vpAH/�k=�WC�96tw�ۙ��)8�6�@��������mz��8"�Xy}�V��(�Ibo�p�AH,�S���4����}�<��w����ZnR]:{�sNxTrQ&4b�Q+�Ðw(�-�Ż?S��'S߄�-����RݛX:��9�aܩ��re�;����^�uL]f���-c�S�M
')��q�u�x���WYᶹG�N���{1�1��u�h��}�42�f��t�iŮ#uύycq�ѕ����Mm�YX3 ��]��ϳ��_��$��û��HYi�y�[�+c�`T�p&�*o޺������������T(����m�a��zkWZ�8H)�`v��T+&{ϥ�',;��+&�P*T
�ލ�Ƥ)iמ�7H6��\y��׼7���R��<	>��CE7@	 ��daYY+(2T�ް!�� ��=�ۧ��z�a�%B�{ϸi�l���������؛@�yφy���\�]�7�w���P9׸k�B�������
m���{����7'	{�0�aX_��ն�R
w�09�m ��p�1������<�;�@Ĩ�޴m ���8��It�jg�
�`T�}��{��wO��n��0K�6�Pk��b,72�n4g����#�=W�IY�J�S���bM�RT�û�B�$y���,=s�|� Ͻ�>�<);��&�h���k�x1 ��>@`(���]� �.k�Yu#�5���'^���s��w�$V� If]x���Q�^���������������oxk�+X ��ύ���Y��|Xi�d�3����3�C��;a�°�����ֵu�!�AN=� �N�+%Xs͆2i��@�B�k���
#���H�Y� ��;�+<��C����i�k`m8I�a�d:��N}�a��p�Aa��I�u׹���ni �sS�w�i|�Ϧy���\�n�.�
B� ��0< �5?$�.�x,�#~� �l@��O=��4�P�J�C���i��ޯE����=)�Y��j�P��D�k�,���������m������H)���bA@�J�}��`lk~��ַ�C�O}� ٺA��a�V�0*vo��P��(�#�!$H #��)��z&U��g�a��H,(°�a�¤�T�:��6�R#�>��<��w5���ɉ�{�i��;.�r�^H,;��N�
B���HV�+X<����-��5H&��h��'�d��!J��%MN�Ѵ��U=�ѕ�%���{�W���
�@�:�
�P�J����a��5���Cu�Z���aS�<��q��a�Ad镇w��d�e@�P<�4��jAH[N�� �λ��g���d*AN��gy�ZsZ��w�8i:@� �����m���s�~tN�x°�gZ�a�%B��;��6ɶT��S���4��7Ϛ��ӎ���=r��)����i换&m�i�f�.|(�|*%�(�[H[@�a�� ��w��AO7��W�u�3��g�
��
��D8��6�Xnu۫�VۜAH)������VO5���q1���:� �_}�F��+R
{��
x�/$�^d�"(p��J)P���N�*AH)Ǟa��H)���߯��{�°�aR
J��6ɶT��A�:��H��|�s/�O���3;k�T��#��� �P{�*AH)z����Y�=�r��ʟ���]��	9�0t���9{
�����*	$K.�B�=������y��	�'�D9�6�l+5��ףu�Z���0�ǿ�J�d��9��+'���s���@�T�yѴ���RZ{�x�H)���D䔛��;���پ$LXʴ�BVٜKss�1K��>�{��j��k�6������AH)<�I�C
���B�����u����*N���ᴂɶVJʜ{�i�;���]f�p�Xqw��!��������`T��瞴�h(�YA<�2 �����9]q�{�p��V���Km��H)�x���J����B�heH(o�������)i�^`� Ґ�;�d)�$e�R �,�BHƎ�/��L��d��ḓi�V��P�40�(�IS�=�l�p�y}�z��Y8S�{�i|��{�2�c��������=��4�_;��:�
o�z�M�T�����f�J�P�{�m��Vu{�|�vʸ�x_�>�+%FL+v�7-�n�%Yk`��F�w(^�.�z�7���O��|�>�0�b%Mu�eѥK���ZJ���Z�������
�#]� �w1nl��(K�6e���֑a�S�5��"Fa.�Ȗ�D����9	'�M,�TD�Y�C���ς���7�%lc)�Aιx�34���-���O��B���'�'�����6��T+%ea��!R
A@��1'�H0|��\':a��P���B�3܅u){�����Ӛ� m�y�I�H,�u��u���M��a��!R
M!RT��p�&�Y(��q�y���&����@�q�o���\�9Û��H)h��5����
��ם�u���
Afӌ�!Y�J�IP�{�H,7ך��km�R
k�07��$�
�X{}�VM��=�L�H)i�~�k��9��}tAH/1g9
�S��}<W́�u����j��_�lX$/���A����Ӗ���o��IϏ9E9):�TP��Bd&�5�]3�g���n��z{�':�d�3��{"�w3(����7L7�E\D6aU�͍Y�%�3�����ô��1F4���h�/�2b酰jz������ .�@$�ߛw�A��]�.UI�A��nfs�l0H3��$�ő�؋o�$��l�I��۝4�4g'\e�?d���*��N�5'͝�L�D5�b!�/)���ǔp���R��*�l�㝏�<P˵��r�^ϚmYe�F#m�����"�QZ�}��>�[������oe���̜��Ц]&�n���	�B�o�����24�EJ��[d.{��L{�$4���� �4`�s]c����hm<�%�r�/�^�5G����2�iY'4�R�<=]��>�������m�l�n�u�i����m�	袉��ٷc.��l�U���C�0b~8���=�@P@�{2Q�οZÜR�F���d�6u@N���$t�MT�����n�28����쌲(�M�N�1y{�ۍˮd�9��9U��k�����{u�;E�3��#|:lLv�G�|�]�;� v}3r�z�}ޢ�r�s9��<�20V��;�.� �mçVWcj`(�zp^:�ʓ�e��гf����ZDI�L�Vec�c>��>�����M�m�}m�	��\n\�:��������w��ȥU�U&9���LjX"�P�i�������J	m	's�g���hg��O#��M�n��䳘�Ҋ�� ��@n�*�c��X�Ӻb~?\�(<Y-�w��¸��y���k�PdT�$���˘��$�rdM]��2�8X��S6������,�z�Ycl���VfW�<"=��{���f�7̥��맬gw+F\�k�����[�rCoM�=�3�r��W�>W����|�~�j�=ǃg��\}����O�1ɇ��s-965�ڙ�%Wv��6���q� x�Ѻ�%�y�0�������s�P=f7�o����v���f�����<.�WY�/���r���u�G`ΓS�v�{-���S!;���g/J=_���C��n+�v�F���'q+�Fh琭ż�X����v˽�׹�»��	��a�L�ݨ��e���K�y����|�=�Hn�o�Zg������5k�z�ơ.�=2�gX����7|���U���j�C�4�[��`�}�����$��w�ҕ�&y�j��	�ם9m�Ҭ��+�����}
L^�c��\k���t�K�4n���	��m񼯹���roN��gk���2%~A
�B���!~&+1$�@���� )YaP4�H)]!�N��P��iY%Led[H�H��Km��M$Qi��Vb,+
�������.�%T��ib�&�Z���۔kL�+Z�m���aQBҪ2[dZ�X���W����c�4��eg�趲٘���Z�j��x	��0�u4,z칒��nc۔����B�yfs�[����\�m�\3�,BJ<q���w2�B\�9�.�6�ٮ{nP�n�=I�n�hr��,��F4BSY�������d4;;=�v���g]�&�!v7I�O@�����A����Xf��yV�
��*���b0q���q�p���{uV{rнs+g]SA"�k
Y��t�\!��GV����@W��x��ÓNx9xݓ��7�����v�\�ɭ�>�WX��u&當��c�k�۞a��%r�R�,8��P�]0�0l�x
�ڨ�s���$k�I���b%�K,xL��-V��|j�,@u�=�;9뛱��������������"F�bㄵ��V]+,�Ď-�3�]���%�Eu`Q�'+e��怭Զ)wm��:n��4�ɥn�nD)J�,���Y�\D�4b,H�髆����W�Ý`WU 8x9mێz�)��E�%��鄘�UUU5;�0��$oj�$$�;��_\��F1��`��n��aA��/g�|�?6����8<������NH�tS�c�y�]�$�!+[���vU���01
m�����s�0qۋy��\��=0z��b�X��TnǩÇ��l!�Z僎��֢��g�P�y%����Ve���ų��+E&.U����R0�sn�6c:]nu�_�����-�Uy��ԒMu�=�(���2p^f�3�m�RU�,�vz�����.�P ^�!��yҦ:3N,Ecp�/=�D�<B�'�X���J86�҄��s��x�m*@k������� ��dgY#kǺ�-ۈ��=���pw6�q����^^�����L�a�5�����o#q��vDi��R2u"�"O���3�ʈg��������6a��Ը�����n=0�x8�ٛw:��zehs���1��Q�hK9��
�������@5�$o��'�+df=��v�Uш��N���:�$bUd�,�j<�u�5c?6�P��=]g68��I6�&j� ����m�9JI���J��͡d��E�J���p$������:3,����T��R.�̥�Bњ�H0�i(N��(�e�x��^`�j��-���1��}��A��E�مTz��V���]I�	��yyP�:0$��c)���@uR�O��́�w7�}��X&M�e�gbk�!9��7�Ñ�0�d>�<]�^���r�����Ϸ�a���b46��L�cm�'-��	���T�lk&]�M��k?&�p���a��K7/`uY���	$�U [�=�󎔝A��)��F�WGKv���ř�#2>�po(J
Κ��gu�O�9��l���W0�=\�A(1PR��������]��6m2	#���Ј�[�<�B�ӈ�bqo7h@�v���{�>��W��p��`�a�>�.J�"Z[��ׁ�	5P�$�}�5�㸈��G�m:��q1#Nӹ"04���+�;E�犫'9�ĥ�>���	�Yo�G�s��fy0wq���X�ă�����w߁���m�x4�ҥ����b̮͹�^w>��U�{���}��{�3�''���^��`�M�$�˗��k��H[f�6X 3\B��xw/x��m��[���7��]�͸���Y7{@ۈ��A^��u:�˳����E^��\T������I���*"�bs�o��[��d��@�j��I��̍��+n]#�	��C�s��~NA٥�s��<^4I�l��_{��+}>�h�h����mل�9�;�I�c���γ��� 8��%L�9.f��e�T��X(M�"���c@5#dȥ7i���*Wh�;��,TTCZ�����ݥ��v�N�C�q�2Cp�F:dAZ�W?|��_d4��D�D�W�9���M����L�ZkP�/.�d�|*�������a�o7��TI8/j�J
����^��~�:��&:[�>=�XqR-H���P�玠G7% 7�G��c�����,	����CS�?r�2C�ws�	<P �_�nw���%���D�cF�[���+u�6a8L�wq�����a�gm3��E��,�<���[;s�cD4�y�"^�Խ���xC��?������q#�f��&Ya�4�.2'NѶ*7uȜ��{e���@'3X�z<�X&>�E�&:U�L�,�`�����RK��j}ǫ���+ER��*�Uk�^s��35��<�$�������a����8�.|䀷n/ys.�:�������غL�����ܟ:j��_�z��E�M��uuKL�
������ه_�a�}UE�v��3X{� ��8
�����:�ݸ�k0�yI��̥_��fJ�s��IW@����L�+��d�Ips�$�Y�����/Z˻r�l�/Uэ3nq��~�jk�	�H'w��"��Ci�$����(NU�r#9"A��ϻw2�;k�z�nM
�	U3��W75��^^}UZ���n΢^�Quw=Rv˭�g\S�E8�s�߼�z���#�r� {r��Un���5f]R�pv��QN��jfn&�rF(�d�`�3u�9��{%�3�L0�yԬL��V+��!C#��$��~t�QZ!�戚�;��fOĂN֯?ؠs��7o!�L��D�:&w����V�c�2I���u�,�0u�e�3���Q? �ՠ��>��,IR�}�[��D�M�'o���Z�՗|�KϦE%"12�((�JJ���]a2�j������v��U����ϳax��W Ȯ3y뺥H��K��1����ܮN�W����� Z� �k����+��q�:�U�6�!\O�=޽]Cײd�A ��ǈU��0�s��z*�/e�9Xd�QGۺ�V��"�"'���:
�'T�!�O��ܾزOf0�q��n�>y�	��%smo܏�S�811��3��۱:�z/y+��{�n���6=��,��s�x���g��� �����n�i��v�\�/a�Q�㪂�y�]�һ"ܚ6�x�������&��E�j�0�e2[1ۤ�._a�l���H��x-���&����2�D�;�3͞�
���=��{#K�keL���*����/�\��r��	��wse������qD��˻��r���*]c��[egS��o��-t��H�|G�F!fܠ Vx՗�y���"E�	{U	X��t�v�M{0P"R��T�p��-
�,�q���	�#z� �:���� �G�<�y��>��d���݌�1b�a��걱u��W�=��]�=�\�`�й�,-�9�l�4��i���t����朲��G^Z�T|�k&�rC�g!�F"�߀��@�E���F�͂���.t�p��U5�0D�&F�s<�ɮȲ|OW?3{���D�?�_?��� ��lU�wOW��4�s�)pI�����H��ѵ2ʒH���#v��q_F����(�.�m��8-��YXI�\\ۊ���˨̯�{팀{�i�	ށ#�w- ��cn����sDr��3���E�9�~� ;�(���j����T�J�m�Ğ�L�Gt FO��-h��B��2��ϰ��;1��n�tlV�ޝ��||`��3�k|��Gg�^釮vN����G�q���cB=5��-��:��Ι�!��?g�3��;���B����R�Fzẕ>��q��&],���g�^g5����^5���=ުzFo9�F9�9ٹWwL}�i~��yhN^
�&ʜ��r�Y���ӻ�5�&��Z��W׳��iG�M��H�_�sCmL=�ʢ�@Z����6��U����)4���z��󣎭���n2Ծ���8��yyg �C;Fk�+�֡m�|�/9��9��}�*��;������o<m�}]�?h����C�Z�����1@�fڇ[�l����Yg.:��f���5���t���\z��vD=�^o�}��X'J�^3%X�?�0��g_kZo�s`�ݮʧwگ4�Us���̀����R2��sN�4#�vf�6'9D@5�"JB��x	�P-��ц"�ar�+�Q�Ysxk.�M�e��*[WD��µX�R�4уl1�k�eb�2��o(m�n+,kuZej�ƍmf���kJ�b���TueJ��j�լ�-��D�M#m��)��Zn�7q�*��+�F���e3�� ��W�����$�B�/`��J�k\����ti��H��7�=��K�n7�Ua�8��t=ԃ=j���W].y�_9��j�0S+��[�p-:M"�VM@/<SL�R��R-~�>�L�!��U$I'3�3ְ��LY]l0H��^ƫ��۞�~؊�tZ��d�o�"w5��+�]ؗ^AV!��AQ�TO�|w:zO��H���c��4�~�;w"�Ă:���\� �����y�/r�7V�<�Lj8a֔�4��c^�m[�v{�=���	Ιl�=��A��܈�- ���0ȝ��t`� 3�G�� =�H�W����i,�ـzƭ�.��=�$i�H���u1�mǻ�C�[1�9�3ՙ� �j[��Ve:9a}��@Ȱ�$�rg��߲ffMAb�㬴��c��`��m�A�n��v��d�3)P�^c2��Uت��λ��A���w-	;����kf��jl�>=T�$wC�ν���j�D��a�g1�l m��x�e����m�T�آ�����rxƸ;�:[��Et�@�1]�v~��>������!���������et�����v���|�n�̭�1�K�(ц����?z�z��pi�����;p�6.�����lX���h7c�6�4U-QZ������\��.���� [�mɈ�&�lFQ��ݑ�?^���.�}�|��Z��l"뱜�2���[9�.|B�q�Jn԰���f8=�ˋ���M<��h�a� z��	]� ������<�}��W��j_f������;[!N�Msl�	n<����-Ťv�vFv��r���8p`oS����I�tyws~9�U�F,J<]tag�/.F�ˮnf�q�[��CM�8�Rd�3�Gw6NK�=�3f�t48����Y���	S�B��q��'�9W(�˶�*��3hY��7�Q��[�I���o;ʡ�vc]Kʉ��R��T7��n�����ڥB��'Q��/wR`�|'�NmA� >�F��C�� �����2g���ex���s�72V-�>��z�"uQ�p�m�ζϺ����a��^`�j7{��t�ʎ�C �	�ü�4���sgfDW����Ѭ�iϔ��Pd_rg��wd�"j�$n=�p���4ω_q�bW����A7����-�1�d��1T[A*s���=���:h����3{����X����#BW��͇�3qn�����s�ʏ�$����o7�Qɤ`ǻg8��6h�>���B��{l�z�֬��X�f׌�6R
-TNT�a�~ ��@f��0 o'o	�g���՛��ӄsO4`[�6o���\&o���|FݶI#z��N��\� ��a�]��:�B�jwP���l�3a틑մ�'�q�Ç���Q���\wD��;�0IFc�b�vJ�O����VFbmr��@�/u���0�aq�R���b�DNvdi�7�$$m�|;�����/v~����L�3$�0c���	�?�t�R�-�`�N� H9���_OT�O�,mN5�����z��M���$AM�-����|�f|{-�"�H7��V��=��>#�"q��0�{�P��}��|#u�F�e>j�o7mA��9�:�N;@s�|6o#ې}�ݭ���aÆ��̊P�����$�~g�^MW(r�P��E4�����u�c:�:�Mty�l	7������VSU1b�P�t�N_Ě�항��o��a��J��j�}�{S�O�9�]�����XۦQ�-�0a���huu��o[��Nq�Ngcn҇l�&�:��Ŗ<��v��pa3����WgP�n��Y��& �iۖ�����;jjV��i���Ѣ�9crr���dX��>Nj�۶y��\�Ҿ��������'�~f��E�ޭ�@ݥK����J!��m����@��Lͷ�հ����؍�a��ݥ�k�`���0K�a�;��)n��(i��a�,Е�i�I���782.���M�*��ӧTR�\ڤ$,�m�(���\n?z����k����x(�ƠJQCs.v��G5E���|�ΉgUc~$��i�	̈́��U󊲟sJ���������}�ڣ�u���}�5\(Vt��ؓj��us����ѵ�]�����1�����f!���$�?�����8Tx%`CIպ����I'螻�1�NAǻd���Z��m�u�E.5��|\�duB �s�	ъbE��ݽ���9�S~o����K5�2���$<K�}�����k�l5��\��踭l��;X�Uw^�畭Q��}��}>���v��T>��� �Ƣ�]wdtIww��Y�ӯm}HB�j�ڡWGk�g{9�������1��ꀷm2;���c`�vHɜT�J��&��]9�Uc`UgړSV�m&f���Uޓ_@D���3�M+�C���r� �P�I��'ss�u�t�}Ę�D���V��*�r�P�^��7�JTMpݔ�{�ą���wt���c;W��4�!����5W����/�$�_�:�Dͦ>9���Ղ���_-p��e�z��ͺg`5`"D�&I'{��R��=Q$��tU(�aU	�l�k�!��mkp��@��l����oH���J#��B>7���/o�$<�v2����X��/�U��DNΊ��{�����|O�5�M}Pi}
�Tz�Uuy?]v� ��bt#��f�n���P*)6�D�A����YR|08`q_���������Ţ������Vl���A���o�%�CN��TMP��z���#v=�O�v�^��p�ę�A�����]�z&��;$e�	��sEERn�9|��|\٨]��ϧf*> 9�Csg���⢯iWݠ�]|뀌۔sD����̺L�O\ Gn�"�#�z���|{�]��1g������w��������<,]�7{�r��� ��go�;�Q{{���n�1F��2{Vo^����wy����}��8���{{����7O���<<�C+6�n��5R=�����؏cI�r]ڗ�����[�z�/�9״{+�yr	/f��B��O1���W�}�q��wO���V&*�<����"���׋$��z��U܅�oIayp�~^Ҡ{�ּ��X�8�{�s;��Sc���h����%���.y�r`'�zm�l�%j�,�y��2B�	%��<}ʂ�w�%|���鷺l\ok=�d�tk��R�xjïfzgN�[ ��>bk|��w�����I�z#5�L'b�z��&q��כ����M ���4䜸��e���;���a���K�\������x�3���H4������d���=�~�9�F���U}n(ۨ�C��B�]4u�̙e���V���(+V*.�qt�T��Z�̂m,�YE("�V��-��&�FUq�bYU,�]�&F�V�"��Q[K[U�1�Z!�5����`;��_�Cd�w�x	6ʝ�&��G�{[V��Z�܊UQ�F�5+iU]��)l�E��l��m�0�ŖեeE˃Z��9*ѵF�jJ[n�ނ�҃����~q{�7P���a���Z���	e�Օ6lݧ�R,�ɠLV�#ͪ5ܦ���046�.��ud��7�i��٭�0vƵb|u�����&�8�X�)�a5 3���g\�S�w�i�v��K�U|طm<r]vvE��Y��v�5&;[t���-�i��a�&��m�N{\��8�؆xM\�g��w<�A�; ;ѧ�t� �-ɋ)�2�*�R�X�d��3x���<��]d�F�m��=L�Ϧ��eq&�͙1y���5�gp�j�:B�Q�vk+R��۞R� �.�y����XJ���SF�i�Z�*ls7�j�Ɓ)�.�0�u�; �2���t[^�۸%�V���ѻ;�=u����P�nN�`q�E�F�[�����V��G����4żhckNL,dь������x�M���l�u��,7:���;|��Y&���qTs��C��@jy���mK�-��K�����5q뱹s�ڃ�7�1[����Պt��Ҫ���t�4K`˺�������5ɷv΋(��a����-���lH��4ճp���e%�h�!P�6����T�buA૳�f��7h��*�����v�q	��j�6�<����x���8�vp���6�8k��ڇN��&�e(�/QKv����;�ۂ�S�hR����^�ڝ㞍�a�2�-�x�qY:z뗝�����R$�o�~�C��K�$���r���Ssg�X`���^'Ƹ���m�޶�0�cL�Gt A���!"�v�]��v��Z
i��Φ>�Oy���o��څf��p�ę�9�{�`���h?��c__C|p�Ht9w�ʤ#��������6<p;��fk}�ձ�Y�*œ���Dx�4c�C8�&�8��E2���/I�y�c��^D��L^r`�i�7Ǌ �k�f�C���*���L�K������M��:]�w0IQ�&�.�FmW�{�����~`�r�r�zP!٥���m�u�}U͒@7*�l<h���2|w9�kt%����G:�uu���+�g�(>xW�m���D�[f�ۇ,Hg~��6.��q�vt ��R4�����uE���5�w�n9]#�Y�#.�8��pSq�23Q�agUcv�2H8t���8/�dƭ����{͒1� �(ĝ<D������O� o[d���+ą�w�Cw�A��d��GWh��Q�Y�u���])��-���Yp�4�R�l':!R���w�J�zSs1:}������?>�6��ц�u.�9��wdZ32R \zD�d=\Ng�����\U�-4�"�=3�����l���Lu���>�䱻��|rLn*Q��Rt�9A�m�94뙖������8l�������^����խka��iD�`8UU:�2L�c�
N�`p�!w2P#�[]��od�v���k���͸��}�ᯎ��� #}�;����Z�Cv��U�'u�$�HG���H���W��x>���Z��7��&�$��/��_{<�e���}���8F�Ξ���_��g٦�Ah�oU�V�lf���B'/�׼��e��PO�;>Q�ܣ�< �(�ef�6�1j�j����C9��'Z��u���I �~�s]
��ve:t�]+�J�!���]���*3)R=�Zr��*�]|v��.sb[���LI�n��gv�A;��&`�e{#^B��t���^}Q�($wsd���B���n���Z�-�U;P:���NU�	#��.�k8*kt�JLqf�j�C�Y��U�����}	N�u%��� <F�A�<04��R��eN!-�fmx�M��Ե��ZU�42 �m@�AJЦ]�ܳ<B��W��n#��$�s��z���V�-�w���\��&$���q=�JꪦRb�"'ywkcp4��n!�W%���2����Nl�}���N��îߟ�ֶI�q@�ˍ齻Ǚ.��F�i*}�R%:�[��/ T�ȥgƯ[$��6N�F�\ӂ�e�>ZO��_�G(UT����^g�9��b�
��Q�5w:I},2'�&��f)���Ia�i�:L��1(�3�3n)�x��=��V�Z�g�Qv;�Xo�=�	��S����u���l�t�V��Ze������ߘ���|�$ѥ>��!���:ߨ�D��x�0��`]P���7,���\g!�ȼ[�T�T:��`��9�QMTt�!A7Mx���������o�3?���8��`�h�D�W6P�\�3-Rv@A�{(=ޕ0Zl�%�WnW��x��$_[�o��v���^ TqF�@�
T�=��蚚�`���?�S�*;��wޱ��l0��^7VC�G�fek��W�������B{�&�g6F��*����l�(%h#��̀e9tf�����I�[�t�v�]����!��{��L� ��c{:fw�0�=۽؞���io4]��z�����{��7٨s�զ4YYh�������v���ߓ�܃���!S��?��C �� <<մ2�#vP{�NM���nz�eY"{j�#�ب�,����>��q�Q�r�2���ղ�H�sZb�}@��8Y.��A��F�y���1��f��6}�͐GI���x��uv��VO�3��> ���ąt%(�aF뽘�WΧ7n�����"�u���n}�O����ͺ��1] �3�yP;Q95��H�;�^^��C��B�'}�����^�Z aß�7ʡ|*���}���ڶk��fs�kz�P9�@�3Psjf#S&�	 �m���7II�Ӯ��U�[Q'orE�2:A��툔b.G���|�.�Ӄ��X�3 �0el{:P$LTU��d{�x��1(�0�wg*�</e�ݚ���V,��N
nE� ���f���9��sނ�/~���c_��4nY����&?�B���1���Ҟl��Q�����0`�H�pI"1v����gx��z%�=���M͹i��qv��(=��`��v��۲&�$��������ƴV[J��[jH�<�=��\J��v�b��#T����I��G��� z܁]Ψ��Q�J%�u��L�n�9U���b�8p�;v����ՙ/q��XL&˰�P�-����r��vy{���'�����5���UQ+'d�7�f��ż8�t1��l{ĸ�%�s�Ê�����1(��s%{�1�{��ܭ��U.�^�Q3���P1�	E��!�A��^g����~}~����2�VR<�����[��\	|��Ř�,D�O��9��:X�rûQP�5=P��ްA��m�U*S�K��G�٫ͼt0g������b�{라i�-HO��	��9�G�uCڤ/k/g4{v=���C���X`�
�����z�J�SJb���X:f F�VF�צ�5����؝�;�V����T"�(0Ziq��l���kT�;�~��'���}����j�*u	���!�	9���y*��Bך��*Q0Ӟpz����}���흄"~�	����Z�A𼵻��@.�V�N�~���.{÷� I"#���>����i�咲��v1R�*��8)��z��z��p��M�+2���crf�Z��+�m�C)m�I����f�=��w�D��u˷�s���#��(`=�����Ő!KI�8�!aA���b���5��8t�[;*�-��g�62�]���R���]#m;w�m��a:W������:U?������nxB�1�"`��,���cw$�;��l�s�l���	��gy��։)H��Q���v��.�w}D!Z��v��6�}__7!>�1��Ő��o�e���_{�.f[{��>�~�����G7�����+I�.��^9j� ziu�L9s��s�'^z6��n���ot��za��C�F�}�Ș�8�ȣ@�4�cor�ˌ��Spn%�ZV13
eZ���UƊV�����J"�T�wu��l����Fժ-j8�Q��e�.Z�F�q��r�+1��K���-�T-���m���lc�*e�e��,f�6ֲ��+[PYKb6�5iS2[*Q,dƠ�-��m+�5j�6��wp�JZکb�Ѧ��Yq����d̂��˙q��[�P�ڢ64[iV֖�Z��жƋt�eR�N5�Ҫ�UV ���֪)30YYeVʕ�h���0ݣ�-h+e�m��eK
¢��ۡd2��y�~/�y���	��L����X u*�3�0�؝$��!M��H�uO4��w�u	��ۙ�WP�ѳ���P�S��1��E���{��e�)�z@U��������t�WDD��8�b,pL�3��ݝ��EЇQ(I���:��-�} 	�@Wr�X#0Ӎ��uYz=��ݐl���H�u��x(��7��Hݮ��A+d�zD�Q&��B��;����o�f2'nh@t��
|�{�*/xSチ��@��6_1w]^�=G\$t�M�P7��(u�ܥ�{�^ә�{�9�@�B���Ի+ն�3b,�ei��q�(��9�ز�!�U�O/Ȫ��Jr7k��v�����f`I�=Z#Q0ӌ��]ԧ�^ځ��+7*k#���}u(ߥ3�N#�t�IeC��׹�$�J�'.�]�D��8kTy�k3���?%�4��Fհ�/M�+�Y۰�[v;6\-��1��a��L�C1�/\�@wQ���e�ƽn�\A�P���a�εky8VM�&+')��ၼkn'Y����Ri�2�Ͱ�3��Fo��L��iyW&Vu�$k��N"������{?�cٻA]�*�˒��m��.��8R�;�>fW�mǽ��WbqTj�p�t�P!h�6�{vVoF,���;�GdD�,C�׺2'���3W�qw��=���m$�Λ�)��]|�w/c��7�N�2߉.�+e��KGm���V�?{�����pޠgF��Ft��l��u��-��,��/6y���*���ҏ	�rǜ����	���ű,�0^��?vj��}�Wqܪ�ry�k��y*l������P��ze�!P�#]�ov��X���7-Z�ȩ��Ԫ�u�I�y��ԣ�����V����O'���|6�:�Er9�M�e.�n���8�������}��A� 7`e)\d�{k�q،CN5�E�T^�؝�������쬷�Op)���{�6[��b���XIԣBrkv.y[�WGg�Z.����87�n��œ�?j�f��2���/Gp{��M�7C��}�e�!`�8��:u�M����/��^n��&���-�*�*���o�T\^��p��i����n�~J��|�E^��{a��ֽ���劐�I'#v���^/w}�ݘ�{5у�_;�iϗG�� )HJ;ӳ�����;`��{7Y�1� uKٙيZ�1�����<����$�=zo����q�۽�x{� ��HrtH?1d��7�%�7�
T�:D�����UyZ=squ�cRA��#��U�T�0ه2�yG���� nJ���N�rЫ ��d�
���@���	�[{}0,�]QoF�M$���^}K��M��	��fb�y	�:�	�{AV�:�C&��O���g�OR���l����K��������5�yVٛ�V�&4Ћ�&�sH���U��l�;K/1�:�ݳ�S��E�Q!
䯽w�����ƭ�]0�R3&�Y
p��w5��N��:책1`]�P�Rh�5I�f�n��Bq̵�����]&3uזj�m�Ƃ�i��]�1)�,< h��Cec�w\��jM-���M�����\�<��%�t����%x�Da�mBl����7��F	�Cg����4k3���<q��Zg���R�Y+0;ջȸ��}Y�W)B�0�y���mJ���X�7`uت	��s�[\b���T2�xu��̓KDo��>��ӑ��g*_�z�� e����a5O�jZ��W2�b�,Z�6�N�߁���5I�{wP�0���W���%P�(�\=�|�$�;�suwx�L�ȇ�.ڝYY��7G�6�Ś"(�|�[�^!S�4��-
���W�R�Vހ@���"QU#Ɉ��Y�f�Z��w6��6����=�A4�N{iy�=ʒi����꽓����}����㳺ɛ<�A?6�8I�5��	�������1���7�ղ��7`�O�en�Ԟr��Ļ큓�Ck0'�Ue���������:ʹ4g���Z�Jj���w�KNcΖ���r{��'T����3��D*el�:|Z��^��^��%�ɩ��u��0��_�c8yY3.%�yn�����"m��N�!�Hy9�5�F���ߟ|ʒss��/f��rZ%�uJ�Yd�A4�Om�ջ��^�8��	�w�6\�S�������^E�*�AF�;>Zb��W��z�z&�m�[�՝�]�ʥ�u�EH>{aL��2�b{bcJs6U���J��DB�V�l�H�ef��mnA�pyp��6�0R9�����pZ�6���q�F�
;�/{&=�!��#0:��b�&�I��ɇ�1�dΉ��橱��i����	���|�����nEn�[�6\�v��lfc�A��Y���0���j�ֲ�%m�6&�c��~�C.W�u	��f��h��ۤwam�d�e�g��}�{��x�c�ܣ=F��F<�8�P���bE�u���Y%�U�34|{�dU�w��9oު��`��]t��L�t��<bs��,�u�7�'a����p?{��Hnw<��o�q���
ێ�l���ӆu-�;�QD�*�ߦ���_n�|�������|J�2�Ԇ�����ۻ��G�$
��+�T0Ҥ�=�Ӷ�s��P*y�]>rm�:6Q��B���g������ҏ��͖�C��6�,9�0��}��4=8/{A���v)�6a�������9)�� ���w��zk�}�?a�>f�t/��Ӧs�/$�B1ү��Z���Q���+���^xzc�qɶr�owwmy����]��Ãw<B��zb׹���;�e�"���ً�F��3�̹��\ԧg!8��P�j4Ѽ�;6!�q�1zst����1*��9���%�")+YR����p��(���-�h���j�K�X`5*(V]4DX�D�ʪ��Q�J�[�c����R"6ƕJ�Uk.9�ZR�J�l��m�V�E�B�JT��Ur�r��R��\�[Q�I�Lm��V�L������#�X�bVTQ`����\L�h,fZ��
�ic�+��fe1mĎ�@�b,2�X�PPEm�\r�ݬQf:@�� m��)mU��Z�cq�@�,�J�i�4���ef[*�E�jbcY�Ԫe�T
ʋX[f���H�VB�kmH�U��]3��� �)������į<�i��\���	��F��s�<-v�	�<�����uyW�j�6B��:�y�d�G��$��m����h���n�e������62-ˢ�R�@.bں뀲>���;v�B�1d=[��	��B�N|�7dw��3c�J)3�F�q����.A���9���9:����m��XQwA3편��*	Z�vR��uc����Nv�ݱ�K�i�Sl�p�c��Ц��M�F����5�ϑᙸ�[�a�4�2+�;�X�B×���{st�E�F�]��pjv������F���.qw@89�(�[6ڎ�E�)�!v��c!�`M�n��g<�d�Xx�v[��sg*� ���Wckh��狮׎��z��f�N��
l��æ�B�K�����Nۄz\���`6��m�5H��Ξ��\�rY��ۊf�X���Z�,�0p.���j	7/\y����z��c�ۀwd��G��k�Δ��!(,'�gQ���UUUr���g3h�cv<�jU�j�7*�3��Æ������Ffى�ō�5�2Gs&��N@�G+������ŋ���Jns�c��@\v���;v�2o�<rn[���rd�s�G��7gF�\�3B.Ωf-��4:$�c��d*�=�ϛ��d/:q�����R� ��$nZ�^�L٥&�a���� �ŗ�T7c��.c>҇��yv��f�W��b��Q@��_/
C��W�G���	�<k��	��v7)=�볇q�������A4�]غ�R�կfZ��h<c��of��[�~ݵ�n��ճ�/��p�������[q�����h��m4�,��Y��p�Źӌ^���Z�FI�
���ЬOnL(%㸭����aC�j�b��^`˨Df��N9Yf�%�*��BG-��l���W��m7N=D��dh3� ��4
�t�t:(�,�Wz��rU��O3+;B�0E�D^���ϸ��B��sa^[ �c~X�IG�K�n��t���E@bp��`�I�W�%��trc�.���r��V���3�"JU��5���#3%ys��V����R!�/7�T���\��d��"� As�`�U]�ϲH��C�0!p�v� I'���I4i���z*�{V�	ǻb�bȋ�ȅ*aȶ�暽�27�P��o�E��]p�H�]���e��>#��q�U����iR~\pd��{�ݢ�㫳3��M�:{c>M"=<ߎG_j���B|��u���v�k�k�-D�!6�i�^��t�q8� �!��t�^窟ty���r� �q���9�`�{�!�����5�9
p����lt����(��U|-~ >��-B�g%N;М跭	��'٪�u���G��ԽO�84��2T;W��{�\�)d��-��]��{�g�c+��qn�N��P�@��ܦD��[#���H�\�'o������[j(꣇���A�c������{�c�^�>��@踘�fH��u�Uq��.���dE��p �n^��vru��N�"M�,Đ!g�&VJ~��"JUv�e���ρo��ݳk,Zx���=�'M� ��Z=1/Ǐ�z���q��{N�b�P'9t���.>>_r��\��{�X���8�{�&��@l�O;)܋�������E�y���qal�-��g6��Q 8cC��c�HHN��':;��b�a+t�ڲg8�ܜ\�3s�Ƌu"��)�����f ;)��i�y�;g����K�Ml�]�v�6�S�Ŵq��R���us�[��������7�d�u�F.�i����%�ԣ����<���-Rs2,�r�.���QWg����R���=��5�_�*�u��;��<0pA���/#3�2I�U��W^�@m������b%QWe�t���W�׈A���k���ֽ����MϪ�t�F�oѺ^mZ���������\�j�F�Bz�ֱ���0ձp�k����N�@��ݬ�����k<ךj�H�
̪�;%�EH���;��k���hQ�{��������H��Ѷ8�tg5άݵ�=B~���M2���,���q�ƹ�y]�v�bw҆�Y��ˑ��<���.�}_�t�с�w�dg[Wfn&��s9�I9n ,��7B���<����QWhWn!V8��^�V�}�j#u��0���}��о�Sl��sƒ�&�]C(��/~y=�ɛw��	�s|�WON�Pc碡r���r����x6�^['ӱ�z�Qs;UCm�f�YT�-(�/R�� ���)��*�GZ�urI��3k/�]��46C�s��cpnNa���PPw�Rw|Ar �؂�6([����K�B�Ȓ-�A���z_}s��ڀr�A�嫪'R�)��ʧo��5�|n���(������줰�|�	0Cl��Օ�6�������q�\�<ER@��$�L���gm�TnaZD��-�BA�ɕ@�7j2hj��j�"�X~�CvV�y�\TY��f�Z�� 3n�@]��F;��D fe*�;%�j�|aG[�_P!�	�ru��؎XnOr�tT[�fj����f)t�'����hj�l��8�1�*��w��X3UČ���:([1���hP�޸�k����7}T�f�k�î���}����B�0strSY+3���.�u�����}�y<�W/�޴Љ�A�3�dv�[J�"I���{%T�W
��9�\m�#3% �桜Q�{L�؆�Apęv�$���An;j���������.�'c��AKzѳf�d�(I�i��ERp(�dX$�t�f�~'���j��%�xw9�z�T����e�E�[���a~N���z�G�u�v}�ߏV^�^��ۻ.aų,фV%ȷ/nv�g�۝�.x[�N�"�ճ�V�9�aS$�]F:`V�Nqێ[���t�����Ce
�ͣt�k��wZ�FhX�Ef�T�z;8[��T%2@p�!vv�6�t�:���&��H���s��:����\��~ySU|��$���5#�=�ϴV���	d H�Q��z� ��V��&�i����<6�eN�:�p�ΑT�%�"���{/�ʷ� 3�ܐ���be:Re�9/z-� �0#� I{V;.b��-�=�r��W�n\yȼ��F6�����uřQ��Â���W+���U�������
3E�"���Ƣ�K�e�"c�#m Mٺ�P۪���xvL�uo3�yIT@��#.�5�;"�Y�}H3�O�+Ƿ�+|���� ��׾��|�7G�;&���b�Ԫ�����l��̑�,3^7��c㬧9�Tz�j�Xfz$��a�;au-��l�؂.��ȳ`�����O�R������!�@��6	�;�j�<��p�N�76��r�Ҝ.ijm�(�s^��`��w��� y���p.��v}Y��[�d�QN>#M";ޞ�˙Y�Q��j�4P�LDOUOrd圠m��Ԇ4���9�`7~5�)���u��wR�E@�#�����G��g�5��a�K��m.v�oٵ�9���f�>hN]���S���	�[��uŜHSX�g��w�fN!���̓�����9	��}K�(���'q1=ǚ3�]{� �n�o��E�����m8�"{�87{+c�B�o��I���aҠ���==�4�u��������׋�Ǐd�s���7���s�ڲ�N?:s��G�*줥��0���m]���sK�����xߠ�N�F|͡�Q�z�=l��9&��>b���o$�M[��||�6����tY[��Q������532cɋђ3f3�HC��K)�tc�x��%$x��Zdy�w�[�*;^��v�q��S��}��W��o�&���u��s��̍��`P�*.�S���j/v��P����=��s����7I��ڮ-�z[Q��5�`�J��!��)9�Fmch�Y��Y��cij ��bI��� �J�`�Ī����T]%H,Y�%b��j��
��d6�I�!EdY����d�V,Xh�4əaF�m"�UE�Q,�X,XM0(��*��,R)���EH��PX��Z��b�`;�\ed�%`)1E�
��dU�+X(�I�e4��6�ek�Jԋ(�b�
�T"�����(
LCl1@f�)Y6�P��Xq�=|{M�ogH�i�q2�����L�>�(�/S�&(̻�J^��1Ju*��`�+<��c�H$6|���c���)��,��-��Z]���i��q5f5h����2�q�N�ד�=4�/oyHA��=�M�g&���|�p�wh@��D.��'Ƚ�L�d�(��<����-�%��x4Q�I�oN��U]��V�Z���f� ���A�{_��{^�b��v썍i�	H�����wpM�M�t��rqe��6���n�}oV�u*���@G9�J�4��A�^F���N��	��	+�.�G �p�[�7%�����Q�8I�x��D;�I��R��\���{cL5�
�'�_6&��P�� o'���}w\��[Ź�=�8�w]���T	�����Xz�B>7���!ʏnӄHFg�Q�K�b���Kj���ئ�zָ㪫�f��
��u���(	VH\�������/�/l�u�Q]g&�F�a	Y�k��5��Л�Z}��~�Zf(�+�;~무��B��r���>�H��mڃ��s���);v��oZ2ٺ,��N�:���1o
¦��].�46$*ZwN�8D�9�9� ��1Xܚj���M�&�h���
�Jl������\���E�m����v�mf��bܮ*����y��{o���&'�<�dƼ�H�ժ�!�N}3���v�:�MD��6��F�Q�
������x7Z��.�� ��}L�U=느y�Q=Î'pe�d��	"���H/k�Zћ�o�����[*�>[c�^[u���;�|����{���GT�t�úW�{%�:�p�U�ߟ���P��<s�0EB=��6��@���}1DNDp�L4ݽH�t�7��	��a�ݫ�&�;@�۾�%��y��Վ�v��#A�Õ^�_�� ���rf\�O^�NJ�,��+ ������l�;�@�/AQH/��zy;]�bA�Γ�o� E���b��(����`�>Hv����\�y෤@��U��C��T��OK�����>69�z�����|l����选'�z�=�N�l��FvDU��㪫Y�<���q��X#} �訩/��=t�F�ZM�Rgh0OUC�q>�kj&�ķu1�K]�O����
1b����Nd������q��I����4/l��U�64C���2�0����֯;�=���|�#��D1Fg���Q]�9�2wE�.� �7)�a�$ȳ�n��v@�UZp�e�6���-:�T�׷ƨ����� eҠv0��kK��Dv��}uM�TH0Ț��p�u�I�/2P��|���X|nG5
s�=��$�4Q'*'�X0$V �M�f�8b%���!�hQ���5QumVc]]5��f��I�p����&����Ef�>r��7�`�W�g근F�%H ��X�Ү�y�����S��qq��;��|�{ozQ��ZĘ�-]��m��)�k�gt��kY���D�cA�h'�\����r��d�ѩ�p�ڭ�m)0f��� z(k���r��:q�T=b=1�WNc��):p�f �����&��=U44�Ȁ�q �ٽ�_�h�{c���VS�Ig���2��Q�� ����Y��qND+���ͭ�Q8���hZ%�L���\^D��Lܚ�_d��V��e=���_�kz��IP�4ф}�ڳQږX�XR�1�eU���V�q\�e�j��m�����Gٛ�bqɹ�mP�],`jM��2�-5��=��q�9�!�i�mpػ(e� �	:�H�cYkM'φo�;����\�m�9z:g:���}}���!id�	/� O��[�۬qe��P��jt��sk���~'Z� ;�RT�i�;k�W%@����}f]R��}{�喁ݐAy��|��(�G���j�b�j /1H��y{qL�@@v���M���A�4T���Iz���[�p����������
�En�8�M5���iф�2�^F�a���:� ���gRQΗ|�$Ojb���P�vYd/��z����s�J�5ϸ�ya=�ۃ4�ْ]�&�d�`��������{oD�j��{@M��O��l�TC�wL�f�]j�o\�z˽_Q�p�8�V�]��}\ur��3.Q$nB$��2-t׺����*-���<uA#�lN[̎���LV@^$^�]�t��.��3��Z�9)�P�ᗚ�ͣ��:���<��7ew�o-�M(	�H��y<T@u6�4t�9�pD4܁��!���.�}!����As��VK���QԒ��e��Џ�/"-ϳm���R9���%�8^@��d>s~�y/t�+��D`��dT�$�#O�cב̕���.��}]ĂE�D���v����p�O��FW@ӡ��額t["L/�w���m�P�d�H��]���S�͹+l�Y��}���Q��@���W�%u59��G���.m��a�z���<��60��D�l4��TŸ64D4�8��L�w9UJ6 #[�71�k`�ZI�U}<�b�0;aA3z���ٝ����N����H��TyyW{*b=��p�S���3�/���(J��7Cj8��$��$��d��+uk�"rFz9 �98� �wa�u�����+��`�4�KIH\�Ըl�(�s^���]<�;�>i��r���W15��� �UN��T$#���k��[��f��|-�>7��5���"����Q�� |i���a�Iڦ�"��B4`P�z���:��r*@s\B�]n���-uҪ+GAi'8ER^}�F݂���M=�QN{������!��`��ҵX*��dH@����	���); BB�j��F���l43rgW�P,4��}��D����,����lf��&M�!$X���fX�7�	�"r���_�!C�3\J����nK��ϥ��X$ ��~��'�ߥ������=�����zТ&N$ٰ�4!���h�Ѣ���s�(s�dσ���~�2s�ف��s�f��	H@?�!����Ϸ��"I��$!! �`d�I�`}p��ɇ����_���C��B�?"�r�����C!������}���$i�~�$ ��/����" {�C���Cg�?bhHs0%8����{!��lĐ��B��gD7��G����/���0?g �Jb�O��H��'GѲ�"M���?�\��HIɰ�Ϲ��N�ک�	f69`\�'�뙢3�/I�sG��H��|��C���S������>� �I���.#���vM��ɇ�>��O��}��=6P~���)�_�~x����O��FRB��3� }A�H|�������G�ÃAO�O�8��	�!C������~�����a�E�>rl'���G@ �|I?���?�r}'�@������=}��?x�d��6����oD(�d5�$�� ���	������	�;?�	�6-!����J$����(H|��~�8>X@$�����	<&�I�s�|��HI! �d�d�9$>��$��;<�y�Z������	���qĳ�@I�-!������_�փ���y0?a����\��@���?���?�	$C�?���O������3����>��A>d0$?�T���?R!��>�����矋��Bg��C_��|C�k�?�R$ a�Ϟ�����"����~���� BBd�;?X=L?�?��a�C���>�!�>`L>D?w�τ9����O���C	��C�>B�?����g�'�!����ؿ���d9'g����������~�Y���ϯ�#��wt'��(�@v/�O��a�0�9�x�WF�jC��d���J����#$�&O����v�����������HBB�����8$����w�I�oq�)'Q��s�dۙ���"C��I������9����"�(H� 