BZh91AY&SYG�o�� ߀@q���"� ����b;��    ��JJ�m�A6�R-���څF�"4զ�w9��j��*6���T�Ʀ��!)�w7*��$�Җ��j����-_a�`��jڴ��bֵ�D�ƶVKb�X����h��Km��j�����KZ��[em��ff�l,m5�T�cV�"�4R�Qs��M�mA���j�kY�j�6�j��2�Y��2حm��m&��k-�c6@�kh�Ka�mTe��6�&��V��iR�m�͉Z�p�;6k05�l .�B���sUU��p��Ti�vN�v9]e�Ҵ�[B�����V���ݵ[j�Y:]�U�[\��}�w���f�5�f�*�lQ�[[mfo� s��P�Bԣ��h8{���(���z

�Us��(<���'��k�^��J��A��( �����o3۽	R�=>�ϵm�2�CkeV��kU�Zo  ,�|+�B�狸�@=����@�w=^�����)��}�|[R������y妆CF��}�|��}��}��ڗ���Oz�����>�U  ����0�hEL�Z�*��M� ��(�m�����}
���
 燎��妕�>�� ҟO��>���C�.���AT����W���}v�_|J�����ި�Y{j�w�RVZI�����3Q�e>  ���
F�ˀ�9��=)A�Vt�N={�R� ZwzkC�ҍ�P����z�����{\�)]��=���jv���=��	k31��)[mm�43� ���@�7���Ƞyr��A��[���A3�A��@]�ٽ*V�����^���^��V�WM=<0v������AF������Q�U��Y�խ�֚���� h���)��Cݺ c��OT�ޛ���(=�wOUݝj�M�鮃]�c�B���=wM�p�\T
v�q@smm6�Mh!)l6�m�� (�������@Y�p@;�`Ab���������[���of�@=�zxP s]�Z��m���ض��m3� ��� :��� �K �����  {y^� {{�� hn���g��� :5۶:����ӽ�tu��=�Qfl�ea� 6�� 
;��� ;�+� ��  � �3��A;��@��  3%� ;tq�4��    �  S eJUC �    �{F��(� �44��JT� 4�   j��	J�z�2h@  S�UID~�    B��$M���4�L�	���������5����	��Կ�oS۬9���E���zק���|�:;=sz�;��  *�J��  "�� U��	UU�ÀO�?�:����������UU�h@ U�a*I���w��Ք?D�Y	���S���S��l��[*m�v��6�e�&�l	��m�;cl��P�pț`M�0�dM�&�l�l�0��l	�D�6dM���l���l��D�"m�:`M�&�Sl)�6�;`��Wl	��(x�a����Cl��� m�6�d��� � m����l��@� m�v�#���A�A��"#�(#���*��DGl*��Q��>2;d&v�(�A� #�l*���;dv �Wl���Dl�P�;ev����� �`q����l(.�E�*�evʠv�)�UGl��A^T]��dUv�"�@6� �UGl
�P� ��QS�QCl!�� i���Cl!�@�(m�6�2�Cl��� p��l���
m�6��&�l	�SL�l��
m�6`Ol��q�6��e���l��D�8����:�׾�"�����|r�˿�k�u��9*c����i�6����u���"Y2�pC�b�g��"$�X���GP�ٿYBcw�\�A�i�L�bf^h*�oeh�j(�wB&�x�fm���j��͡����Cm�Q_Y��JkLq��Y�:�6�m+�9RẰ"W�)p�	����Nme��e��Y�x���$�7T��X2��z��5{VM���Q7w����Mao�}H���o��Ү݂��sdݻ cU�� �+6:	��.�o�7���W):yw@���R_e�u�x��7D����S��bPQ�R �cn�eݧCY���Դ������g[͂�e:ǫM��n��)�U�&�+,��tŨ�GJU���#l^����Rȳ��%��ǗW��!��
/��;���!%^��Ԗ�VL4�c�4��@�-T���;��E�n�����fCE���]K�F���]���*���$�̼r,e�[!*�2��2�6��#V�ܱ�ӆ$V��nM3]�#eJ�"�dcXXT�7�()�j��a�'~'"�Nڲ$밴Y�٫p�t݂t�Yt�ɛ��	%�� X)�Yj�i�f�4#�n�V	�����-�q�=��bfęJ�k3o&'����K&� ȣ�0K���Sܲs�\��Z|���X�G��sX���F�nS�����B^��2�cj-�!��0��S56�MdЭXז�E��u37ih�P�iF�Q�f<ط�c�6��uR�S6Ĩp�Y���.JeJ��s����3��1	
1��-©�L�� ���z�M9�5m͵�D�s��{�D˹�n9mC�[��f���e�R�T���Ƴ@�1SӦ��37�x�2��&��,b�W`���r8�0U���H��!q�L�؅m<�nBd�9`; X��Y�7*=��ú�U�"��F�+r�Y�����ƛ�ˣOn�����5�/j2���tm���46�m�wQ�V��wZ�ln����� ���E�)��f�S^�J+�GNjӑ��z��d�*k9UI�W��/c��@ҡj�" R�n�@:-�@ӻz�!�P[Ws���M+(I�#����5m	�[�֨�T�d5���!�Z����M�NęjHr��1k�D�Z�i)WW��1TF�r�������N�V��j�bW�D��`ó^	�ݨ���-
�.m�{�u"�z��3%�{��HN�5�b�8�^�QKHt�#���ϵ%�Ԥ5�r/C�Y�HeYqa���̫��+Aڏb$��k�����
}J��l�cy�W�+,hW�ܵ��BFنس �ڽ{[(�Q�gE���j��'n�;%G�D!y�:�4bI��D����1*̊w4$)�I
�W�eH��/p7O%� U��)L����K�@�i)Y��F��N�����$��ڭd.Vr���u���JT��X�[b��u�eZ��X �5	��UЅ�cX"2�,�n
﹀���I��E��P�߹��v�\�ot����[r)�d����
memqޅ��|s\�s��:W͑���ɫ`��>�*�kq*Ģ� Bn��B���b�x�&��̊��X��������5A��j�W 4�b�3¯e�@љ�Pk!���!��X���dW�f�3YjȘ�#��UeB0(o3�n�ʗ�q�&2�w�����e ���MI+�
��6�M���P ��hx'�L��Dc�f���%�V��n�aT6���|�����0&Ft���\�m���r�*B�j������ݻR&���]�>�t�iB�*�9r)��刞 � �bX0j��lݡ�B*8\5�ۻz����Rl}���$um�m�d�>�N�ͣ�d���u2Y��T�,�}��%�:ʠ^�<F�i%�.��Q`�Ƨ_׍P�����
]$�f�*޷�������t���x�@bf'�5|��Ysh�p�M���l�{{1U�<�6dD̼���PՃB �m8�*��QQr-�2��m>���t8&0*�7��uT���0��͠��B;V��4�$`�j�[�F١��U��De�s���聤��Ǵ���`Hh��<�ܨKyWa��v�UT��"� ���F���y�e���U�oLՒ���B�!;�Xê�
o4It^]"&��/Q�8�,���=��sKe���2�P�F��Ȗ���Mu��+7ڎU��Kݭ֘ՙ�Dց�nf�5����+8aW�(,"�y�Ⲧ���ЖI[�X�����62eQt#*�71,D�j���6�h�p�4�ՑW�h9	T�a�S��
T+�b�̩H��J��1K*JsF�r�f۰wq�ҐJ�.b'���6F,R�/f�� =E+u���uazp��}tq��I�@̀�e5�׬��+l2��7���o�R}�v4f�q�)������A�u�*�����v��Ri�ot!�
�͛t�@�(��M]"($!	�6���l�Q�&3�"����o*v�1�Қ p���SpN�� ���5��hʽLdhQ��.�Y�oX۹F��0]ڀ�_���A���J�����W�W[R6�h�-�[6��#h�|�n�%��X�*¯^]�lkt�U����\PVm��2�3]�Щyk#�;`�V���1�]��i%f�wh��i�;g��g	:�9YN[�y[�w/p���pf�v�y����6���ѷNQ�� �܅*yEP��&4bkl���["!����k0#d�PխҫE\v4=o�D\�P7[D���&��X��xra��뺡X�Fɻ����<�cJ��Qn�U�f�v��	#0�h������x��M������e.�����!Dm�ӼF�iv����l%f[T�WcCl���Ū�̛�1A�j��a�l�P�^+��4Yt�P)$Z�����Se��ZҞ�jК�w����ޚ�b����z��m�V�+hcwo��c��]5=�Y�o:��ٕD�v�Gb�4�f��Y�����r�[y� �Y:��J�vJ�pR��a�u�鼻��N�l�����6mR��F�f��w-���W��F3v��������mc�C�T�����<�ur\�.�Y�3��m9;w*U`#�ҭ	Vj���cr�;��ǎ�c�v=���{A���║�&X%��Q;�'W`���i�p-zcX-X%	����c��fnl�F1�hjX��4��HY�����Ps~XAx�U�!b{�A�ùG�v1���FS�*��PB�&�)u�3O�ŒM��Sx�*V��86��Ī�)d�![Gľ;�`n�Q�L*�z4��Ż8١�J� rf�x�m�gjCS2�#um2�!	F��ި�7�n��L�S&�6�Vfi��o*X8�
am�d�cjLj��i�I�P�qM����F�XF�<Ѡ��6Kn#Y �,�Z�xs1�W��ji/)m�T&�r�&��T�Cj �@Q�F=Cv��{�4i�!���� �I[��e�X0m�Ӿz8�_����ƍ*l�5��ZL�XHR�^�tޡ;�v�\��ʊ:.�.�L.����ܺ�d"$�\�\�+u�O�X��V�5|�l�}���*9zL���I��:��[f���mV�&e�eMyCj�f-�G0�
�r=��&㵛`�Y�#Qƞ=W���8�ґHa��b`qX�7f��f����`�doZvѥoV^���_l��
5`ذ�5wR�
`y+D�4--Q���?�vb��j�B�l��&�h��A�R��|oRv(���S��j`�#��b�C0�$؊;��H�kW!�HT3еP�kwJ�[�<�"���F�y/^C�X�l��h�an�Y�aA�E1��Մ��Օ�����5Ŧ�x�8��	&�=3���$�S�l�4�C3՛vrT��jgcM�z�SE+���X�6%/����$[�tt�U��&�FD�1��5B�%ٵ"ԭb�z�J��sMm�.�r3�aʷ�q��+ji22��"�� ��]S��	$�%��	�rf��h[w�^Ai����i��:��4F]�9�р�I�y�h5�X�2��0�[:� ��$͇t���v��R�V1��yw�.��T�s4C�+kra��P�r�����{���z"F�%D��w.��!i+Pa1��gb�6���k2b�G�j/���րT-�:)<�9sU��!Ӥ��9rҳ�w��Sm,T]a�4t�$������yx�:�^���4�
�X���W�	��$Aу` ����M6��Z݂�aǕ��]=�j��(�jh$��q'�k��u��F��i�����b�Hʩ.+�Y#m�����т԰�7�eniK`��6���V ��zS�k������tپU�K#���3EZ̢t1y��8f�z4�	)�<� r����fEX�Y�i�ZY���6�B���x-&��E�p�k���%-��:�V�a��T�[16�^5��x���l�|��Mн��VJ
]�����Ww��F�[���¦L�	��KKmk�yz��P���Uݩ3na.���`,��I�{�kr(�\�U�ƛVA@����Fi9!F0��7��[Zpˬ��2�L�ښu	J=�,쭰Nau�'�����a��U��p�,�$QuOJ�,E�e�J�#P+T�tp�Ҩ-�E�@h���\�)��*�jdf�g�W�YQh�t1�7�:2��x^C{�lha��u�^�A'{+p���F�D�̛H
�N:�{�Y�:lL7L��K����CT��[-�)�Z��f��t�Z&�:-i�#ߓ`���l�3g��*�(�NΧ�0:��z�������pP[��8��@24��zܻ�{(^�b�\��#ji-�\�%��/F��S!������i1ެa�o*�]��,�ڰ���+U<���F�j=um͗f�61����:Ů��GV�]v�%.{V1�؝����3�q�eͫ�XN��a#3&��{�ދܹ0��N�A�C��q_
�d72�J́������o�#A�j�E�L�?�}M�<Hm����7b��R�Z�6�	>�{��U��i�ٮŇ�����BZ�e�;��m,�4�v7P�ġ�2�C��jXkp�XN�Y�ÍV��hf���2�)tW��V���]�Ҵ�P���r�C#�e�j��)5i�K�aj]��j:��C`ek�X�J�q��7[J�8t[������A��Z��L�{�mM���`�����ޓ�(�*������n�YVs����d�${(�qE��Øh|uS�0͵�35����i���,ͽ�r��:wf��e��q-ܽHkך��F
B����D�l �i�X �zH�� ���tR���R�2L7V�TU�����x�7a@���,���ݺ�$��Yx��i0�n���`{AKv���s)M	�b�2���F�p)��73(���t������3{��7a�.5Y���h�z:f[�x��ٵ-�79)v��w�0b(��@��aҙ��)-5d����o@l!���bYO�b�hӋ*�ld.��e��� c�/��Л�Cm��R!X�m<��.��
яb���^9��)�2k�I�Y����eY!������}w\�u\��E��f�b��w���L��m�X6����j����N(6	�!Z�ܕB@h��۽:��f6D��S��p3G핵� ��{b�\i��*�dZ֪�R���՝�4�¶kˑ��p��1�a��h���r�/l��i;�a�kGjP/%j�j�geh��-f�rS���ڒ�w.����8��4�X7��URu�L<�Fl��5��W*U��B���"�f��X,�(���d���*��Uܷ��ܥhݽun-�LK�C�]Y6�e�3J;f=�wA]�5&țۺ?Jn(�i��f��7r�"���"w�[�&i%�)��h<�w�m�	��yzN>Ҟ�A����o��IJ'};s#��8�RÜ�勶�/�iY���5� �[,�)��zO/�(�1�n��Աvo1<4}�'��6�[5.�F�����Z:�ܪ�CV�2��Σ�r�X�f��z٫��Ԙrbء�eL���6n貞KW�[)�K�����!��Ĭ�&fLI���%��q;�vJ�f��2�Su�N�Ѫɹ��T)�y�J��f��<���k	��&Rʦ���AkY,��nh.���ǅU�T�Y��	�Yvp�ǔ�i̗��1aGm֙a`������+��G,<۩�f�
�pi�\���l7�Fi��+C�h��*7ov��ӵ��Rɬ<�\Gy��7�t$D� ��V7w,�dJ�)�Y�4ua7�4���Z�u���um�	e\�!E��&�I���U�Ade��ɕ���J�C��zA����c�*D�ҁ�]2j�ZbJ��Sg��٠t�l�"m��ՋIt�B�"�Y����V��&��n��J[F;�%Zdk�$pmc��5	 ff�x������%b�{m��h��6��Č�&IA�-U�h�k)#s�9Zt	��<?l���aX���wT�MI�W�83fM���j�e�CkI�a@�n^��Ap�+e٢��RPź�	�r��X�}�F��O]�?!D���S��P�<ݴ�9�Ens��)4�$8V�8M�lo����Y�&%�T�32�ӥڪ(�DA�_3��F�l�5��V*-��h���[ �V{��p�Z&͂.���(f"�8�h\�M-Z�nkj$Z\�Q��j�^.�j�ڜ�l.���Ρڃ���ir�Uٓ8;`ΰ�h�;u�e)+��,rd95ֺ�Ѓ ڼ@`p���X�D��h�7\z-���&�B�8R�4�n�!P��u���`y��� �.��?�r??傜�����?K��_����>=�����r�3����-mH����R��7�^�,�j�Ew�R�|��Y����]��wxo�Uy
����_V�eg1Lr]1��\�c�o%[��D*�VYYO1���"c�	�r�{�Rl��Qs�zfv�	����B����h�(��O��Ұ�a-L]�ݨ�-h|*aQY�i�GERj�֚�ϵ��}����)(��T��q�cS`�7E���,]�u�m�W�����.[EV��EI����l�p������Vw �+9��诉��X���a]��-� ����f�$ѡ�u�>܄�,�PG�S�f`쾻<��qѳ.��;I��5�<K+&ss6���v�]ŵ���pŊj��WI�Ŝ���Eg�}In���O)i�r۾.R����O~�	�+s�g�p<�軜�aG��U���;�sb��s.�v�FwM��Y��\���T=ʱ�J���r��WrT�71�����c�;O/�)V�ܹZXVA�]tY�2���Gp��UmC5�� (JO��o���%�oj�x�4v\�uP����Q=x�E:�VZ ������-&Ʋ��{
��y�&��(V��18`T&QN����QBoK]��ť�����	�2�V��X�R���ݧ+1�����;m��Y��+h^��[Y\.�Ǽ���Z{
�V��8oH׋C�	T�EΪo��y;k,M�J�H`����su����3mRV�]���gU��C�yJ���K�&���S�wrH�녽
h�{uHS�sLZ���h��mN͖�ִ.,�(�\�NB��r�7٘F�齸0���W��G.��.5�o��f�V����s�{o��`yRj��P�G�����edj�d�N��Z�ˍ-���2�\�[|���\r��sv�-=���|o7QbRl1l�.���#�f�҄nM/2��죝c��Iy�����¡Tp4J�#;i���t$�{p�;˺���_�>u�E$���bcJ��4��7����*aӟM/�c�rB�>�a�|�v���7���I2m�X7�'�>
��am#w���'i�ȕ�#���8�6�+��(a=�װMc8%�e�L)�b�v�͎�:�j�R�~u����2�f��>Z�RJP��A(�+x%�9{B���-��ϐ5{{���&�����dh��r���vn�N�+W�m
�,�2�V�Ȳ�V(�e-�ْ�I����Ӽޥ�@���:g3�hT �EM��̾�P��'���ԊI�ǌ�̦�v��tڒ��S�&��Y�7/�ģ[h��m�΄��S��F}�b��~��ҡxj�Xx3��z�<�!��;X��f#*j��ա�؄��[�],�v���O�:����(�j�V2v���K�N�C����"cs�e��ST"NQ�l]m���d!%���r��a��qf��Μ5�%o_%�1NsH|s����L����{ټ�1D�))"�ޖ��9��Dg��2[�˰�Cu��x������31��Z�LVN,��O&�n��%�7��w)�2\�g�°mA��� �l�{�jugMbhjc�C�BĚt��V-���ZQ[�8-��V�i�*�d����Y�[[])]�7m�y�X�e�C�雴�5K�Q��pu�/����kdOQW�,A����7�{X!Η`�v^F�ɤ���I1O�@�9��W�u�SX�jWB�u���9L=����43^�n�!�s�M�sv��������=N��s7��X#�v_+�ns��+�Y�M��BV&�d��,��y{���f������UyS-^��vz�>����d����Fvkt)>�l���t�r�άo���JJ-��A��;S9Sh�c��g�
^���3N�n��ej�gK��� ~�p���q̏��7N1��x�5.�:���e�ؽ�[OU�2m�������Wb�T'
@з!�XD��,#�N[���6e�S#�Gm&�XfW��v�j� ��0<r�J���V��+���e��(�.�8%�gX;�i�ޣ�:VY��ٷ7�7uS���&�"�p��Pl+�WönG����-`
���p&B�`���N��J
�<�+��E]��Դ�w����7���06����:�,���m*3B:�+䯷���>�j#�g�BԨe���X����h]��g)t��t�ܮ�ԫ�g�#�w�:Z��5�����W�G��S��V2�z(j�+$y��t��^��Xnl��tà�Ԯ��ߓ

�i[f�w]}�7pK��'e�Zo�#]Օ6K�Co���%�tQ��I�L�̈́l�B�=>]4K��U�����w���>�+�췖�5:��N������XQh���ރ4���pM�)�=}�����Xos^B2�v2T`��+j��y՜+�̓!D�RdJ��̈VQޅ>��E�B\��tǈu��k���u�w����3CX+�opQK�A��Э�m32��dE��#`�X:&�5�U]S������I�zf�C_6��Ѹ���0^���c��N�(�/'TZ��J	[=NWnv�ED#�Q���)sљ�Tq�c*��s�cN��xJ��xo�ͻ�r�s��&�:9��e�q�L������U�������Dj��)��oG7����7y���V�4u���',���-�{o�E���:"�#WK࡙ZB��7��9km8���/�����y2 Ȭ�v
!����=��֜2�^$r�x�)�vS����N%ko��8���7ӂ�:r���o�x��L\�z�aD;�y���3���v�#%s��4ORU��H��΂��I�Hpa�I���aܽ��vn	�n�^Zhah����������h>�ia�[��h�[2 #Uƭ7�]������Up��kEG�Ei�}�3#�r)W2�ޝ�.��ִi��;,:��]\㻂`�3�qÊ����k���:&+�h�K� ��
OfWLA�9�����j���i)q��e���+2�'Wr�Z�o�r��� ��q��r���N��J��lk���ԓ��;�γ׆q�2��2�7MhIլ�b.}g�]g�O�cŴ��X��(R�?��+ʎ�ۑ+N�d�-�] �y����(w�oȰS�.��0��rd����נ��[�H,�ޙmM����;�uhP��`���-{V΂��۷sWb7Ǳ͍���ָ]���:i�{�E�/%vEo��;���lYf�.��8����u�e}f^at��;��E�R��9�T/'aQ
�����xj��G\K�}�r}�����5#��7��p���8��Oi?��uq��l���r��Nؓ���-tp\O�<#���}d-WO�J��ֹ�3T��n�zL���뇚[�jŊP�tڃmLL��u}PV\��oR�	
�5�*X�f�oʌ�CH̷�u/�U �WG��b՚D�Hӗ6`Wgo_uXO��;H�s�_u������L���(�{dէ�_u��wQg��G�n�u��o3H aT��soQ�k_@qe�Zɚ�ڗq�"��A�zFe C�ѫ��xn�w�N;�L�\�ko�e�Փ�ϻCx���s���;uU�5�5Y�ݤ�}F�L����f.fv2q@�Z�T4tĬQgl��u62��m?��s�q�o��'�`BY�n��|ޒ�ߏ{>�
���hY�8Z1�p��(M�ئ��=7rmAs&�n����9Շ@��0.{�m\�4v���
-u!!���Ow��:�(�^��wٔ���*ͨ�J����E	$����k�뾚 �x��)=���lǒ�7}�nk�Eʚ�(�7u�����5���p����1M�́_v��T��on�ܚ��}�z���ar7��1ofc�\��;-�l�6��wnԩ����SZ�i�b��Z��`˝A�%�s���X��sǉ�2�'x:7΂k���q"��h/Y(�f.�VN㓔�E�#	�����I+'�n0����� ��˾�yK���6t{�3�c7UH��|F4��ƽb�+�[��{���}Ss��ٱı 6�v>A�*u���\wB��L�}Pl�lW�t[�2va��Emc��6�ҐUQ�G[Ɖ%u���P��֋�����;�^<���;��.��b�Z���`ϋ�e�'k;8t������V�I���ۊ��R�7�Yv��n���R��*��.�;��ǠWU���'K)P_72���]��C�|�gM�cqe4r;���q�����+�!� �=�S��3#�h�;59���N[�	d��*�>ؓ��Bwhi4��_P�N��c�b�x��%jȻ�6�M缭�������T��{tB �F�����1�v���um��kp��-_U1�$=7m�[��4+d��8��6ɥ���`�R�8kt�áO����|(��!��&f�P�d��1"U��iL����E���
�7���Z_3d�˩�-Г��-��헽����i�8�ˤ��S]�Z�N��t�[�xFY�H�\���[��$�t��^ͮ|�Ѣ�A�˕ fE\�]��ZY�{MnJ)0���m���V�):�ͺ{�;�m�>#i;��J5���ic����]�	c
�Kft�6��v{u}���qH�_Vj��WcP�Z�у��'�xd�����U��Ϯ(Qh�#�Y4�e�k(�.��<Qa���֪J��G5���Y��c�Ԩ
��\&�Z��MA:�M�܏u�:v-μ��Q��)p=u��;$��wF�ރk�%v�n��t�-�I;����(��o��^𧦭���Ni�6Fw5������q�(F�7GJ�&s�p�n�4t�-�K;[aJ�I�FJ�*ݒ�7V1��`�GM뒬���ű�N��5ލ�Olq�MW�e���B��CL;f=+8n�S�^�6_��eꧬ�^�4�|]�(k�Y�:Z�l9̂h�ZWl9Oe^J�	S���>QҮ��Z��.�B'��Yj��}Ҹ�^�1(���*쪰�c��L]��fRU�6�(�[�dt:Go'H�\�U����7N����%R���:�3A*w9��Na+��iW����ۻ�|�r�OhyZ���q�U�7*sй�<_��uz��{���q�cBJ�YX�+3{dF��аΞT�7tzb�/'2��S۹]��`C�S���8Xn��1Q��h��w(���R,�7C�6.����Od�k!6MF�Ӥ���T�+j2�h���뮸-v�E�;"�&�U��Z�^�7���{K�����$N�x�(=��Z���i��E��#6�[(�a,�����IX��+_0��Tm�3��:���N"'���빓5��[F�xh�� �I��A]�k��L��Wc��oJ�r�/%��n0�����v.�q}��"\�n��liM���k�Q3x��9`����1�{T�
�}ߑ͙p-�_&��X�4�u�.�<�3�N���6 �N���I�-ewU�]���Bl�fB�2��蔽�X1��k �E`�Ss�F�ru՛�L�AJB�[r�!譏qT��2�d�w�����4o,��nn��lV]�=MS�ud�+^7 �u��㸃�-�;��JAj�\�ӝ@�W�0H�=s��.��1
%��A�>�YlO��¤��v�b�Qܤ�e��S��wc�Ξ��A]8��yкu3F�ڴ���`��d��f��� �u�yK�L�����B,��a��1�9��v8ըVi�cK��t����{���8dw��E�]��I�[��Y�*�_f�'�t�=�7����6���쐮Lvt{S��¸8�w�^*V$�.��|��w{�0x��}f����1�	룶�WL�\D��]���2 !20j��MH��.V������/��n�9�&���+lZ��%a"�ލ�@�b����ݝ���bF�t�E7�(fh�������X�1��8������J64_;Nq���ڷ�YȖf�b]�B̭��Szv��,��%'"8������[L<�v��ܢQ�, �I+M�5�"�����I�(z��\�k��dΜ��DA��N�컱���`�H�cl�9�lt��.���p��up\y]�b�L��kl����xH̲�oq�q�6�d�+���.�e]��i�s��7�Ɋ��הw�{Mr5�e��%����w}l�:�wX�sw)�G-�LT�ͻ�m��O#�X�4$���!��
�F�����̳�\�7����v���*�q1�'����+�!�s�� ���=� Z�)��#�Fu\�7@�kx'�$����J��t�*V���b�&ͬ`M��崑�;39���v�'a%�2NҌYۊə�����)�n���;.��@�,��t���B\�I}I�\j�vg��� #R׵,�;��i��,3���x��+�7,R�
��{�v����l������u�;m�='(w���$��I��Gt�� =W������9ޭP�(0fA�u��7��6�!�\u��X1�3�p�!�2�D�4��a�i��U=��]�i�w�.�MD�eㇸv�v
��<�U�·�x#۝�xrQܑ���r��MJ�9U'v=}M��)o%�zk`�uxx���%���r��R9V�$�I�IP`��.�S1!�_l�9�5)�7G7u�d��A��]k֞a:�CK#���G�r00�� <B�'M[!qI 2F$��G�?2/�5<�B\�jh8�w��΃�ȩD����?�/��⛍� �`�Â����O����1��
:������
*/�����Q @>;���������=���������}���5�u��y�TY��<��T	�����깆T��e�0��L��{����[ˮO1Mh���Ά���`�*N�A y�����&�m��&t���S����=Ķ��Z��H]���슋Q��LY�ԗ��e ��vGb�1X����WE0�"�j6o$���VNsr�D�̶n�o^�oJ73�p�D���AQ��z�0�G��*�\��̗'-3)'	u��J[���BP�9xm.��;�M��y.EŠ�N��±�i�Ew`��Xo��� 3#p5�ܷ��:��%��-��F�F���%��;���Ñ�4>�܀��S94K��1Hd�8Z3���
X�S?X	�;>���V��r�1�S:�mv�f=�LR�eq7�o�`�-��[�J|��+XN��ܻ-l̊�L�C�!�;�l<�Ôۈ^�{=��-�Âj}$�5)mn���6.�ť,�7k��8��~�|M+_%a��[�W}3�pcz��M��ݬ%G�	g�j�q����IW�k���X7��Y(�뗅-��*��2�' �[ ��6w�Ȏ��6uh��b�r"���J'�y��C�/Z{&�NU6ct���4*Vwx�ݒa�H�j�3XW��y�hRH"g�W�v��C���]f����$0�4�S;�=e#���sq��ՙ�m�j��y�����1���3���Kc�|����EM�[�XsdV5��i,a�E�x���o诓N��]��)T{��4!��*Շ�i��t�(�q�4�����՜�9ԛ��ռ1
M
�f5���
�Ӽ!�ݿ���N.F�+we\�K�m
s*s6�ܥ�)���g�P+lwے�w��q�=�t)U��*V�P\M��,�"<+M����w�î��3t�e���Cf��t�"�\�z2Z̺�+^������c˃\�ц[T%�ٟY�4��ϔ4v=9�86ĺ�ވ%%�<]l1Z(���o�0��Xʃ�N�XV�����[{h�ɡ�:�k�B��Df9H��%r�(��V^�c�|w�xj�e��R%�y��t9xkT�����Y�L�!�=ou��J9�����:Ko����9�}��\�e*��|z��d����#b5d�9J��]�Њ���U�i�]��`�z�I�2��\���g${��+-�j�R�ET|�s� �Ǥ�=�%�r�qu���}&��#M��3�O.�J��������g�^]�P!/D��4��ݾ/�jqAX^dS&Zz��Q�f�9,AW��yʺS�����N��� x���".QS��"V�˩�"$coU�u.Zt�OS	�P��`s{G]�lk(Ѳ���_�$��t���Ɔ���������|���S��*������m�J��);en��p���2c�)[ٟ@g6Rl��P�3;�����w��ƶ��hOp���]NزL=8* T���u$�h����2����얹q���vm�ES�Gu퀀(]\�'uɣP&.VeuZ������WÙ.k�5�:��Sާ�WM�o�c��Љ}�<�V�j���pJ��s��WT2�=��B<-��a��B5T��#D�jE�׼l��W`b},R�=�%�,"H�z��[H�Fm��q|K$g\���ך�ŗ����&��kp�+N���r��q����_&˶��]��͜v��-Xg
9���]�\�2�D����C˲�[ÁvU�h�woMY�Y�tK�������;����W�x��iTz�eo3ʅ:0���s�r�Wu��G9�p��m۴��-X��6�ƷM%گ��V_Y�!�z�)cL�ٺN������]q�?V��i٣�S7�1$q�����ksv����J�^�����odY�%32/�Sx��ċ��P(�yhS��q�vlY5�-�
����ɯ���[��3�ط�R!;(�e��:s7L�z���H��>�w��h��P�d�w�a��8��+�o��7���M���}(��n�Zк���~�cG�[Vө�2�Z��XA:��'=��r���7��s1N��b(d����!8�}'A�k��I�V!�Q�ӣb�آˤ{��$ro�����j�Mm#s�M�u�����NΣl�c.�HiƑ��eo	L��2����DX�:�� ��QA�Gf_ee�}սE:��2ٚ2�WI�������{hQ�<N�v,��Vsu%B��;�Ӷ�.���uk5ھ�B�'U$�
�����\�G�Q>x/L4�{�y0�Q�{h��ums�ECZ�p�4�4����BM��m7���r��L(�4ө�Yu��s,u-�
�b��՜㙖��R�p��D�m`�(�!�n���"맊�)���fotkOE}��y`)4���0!Dm��WH�'��/���Lu˗�� ����%�i���.$�5.M��áX:�XL�|��[4�yӂF�6�%cU��J��_nl&g���,?���\���m��"��k��3)��-|f�4{'O�
�%cS5����4ii]�urȂ��sg����L��z���K2���B��!r[qh� ����e
R�b�	YE��`��	�q��ll��T��"��̵����'Wz�G9�yF�g�xZ�K������:�
����c�P�����)'m��^�x�����O�'a+OB1'[fL��̔`+l\�"�=D�k�x~���݈ͪͮ�{Be� Lp7ͻW"˺ː6��sY8����rM�+�������U�bYYU;���޾]v��xz<�aFx�;H2,]m_`�6�*t�&G-]�N�����6�ldnֱT���8��}��!:�]�g�l��
]����ۙ|��K
a��Ge֕Hww]>�a���R�1x�Qհ�c��Z���ySR����;k�2>�+o�	hӣj�V|v�['�&��E�q�Ͳo�W ���	�@ˡ9�Ӈ+˶*�a�*��n�N����}>�M*����z<������5Ԣ�d�m<�y���S����/Qk���C�� F��w�7��s�7��4,f4�mr��f$�jvc}yϠ�,=�\9YoT�u5R���s�$v>X:��'!J|.Q�U���5D�c0ȹ:�0����X����+b�)�YoP[Yl��Q��[L��҆(�"2C/��J��g�G4�]Vf��hi�z��`e��	z+:�.��'ʮDR��z_dDԎ�laiV����olǻ�cKW�r搢��)w��Xk;Vp���"K��Y��f����RHy������u�ڙ�AtF�*�މ�i��V�N��5ӯP�"ˮS5�s�Lv�kK����aI�^Q]_�g�v��څ���\�g�{ʐ�q�b��U�98M��Q��ØE������
 rW��Ή8(]�.z��� @��q�������)�V͒Һ���B�t��5�J��ۈ��`�UM�n�,�0����z���F'q����6f�:�}xt���GsTp]���]�����)�7;m*w��.���sXP{�VZ��d�N�����ފY�ɔ�M��u�ڳ^�=���H-�Lڝ���oK�<��ݒ^E0�0���j�J��m�]D��e�+
Q�,��3�-�㜑�U�b�1�ņIm�u�Q�;U��
R��ul����!x�J��v�9W�T��r��T�a	��&��,"�^��Z��ͻ�E�,�˛��@��0��XV�j�rO��|2�wL��v7w�A����V��GO�WNQ� �5L��+��]/w��Xg6.��[���*����ov�@_K�ԥcy��e���#�-�/)���G֐1��r�F]�L�*�]uy�F7����J���݅�Z)�L�a�݊�l��gu�S3D}�8�f�M׍�7�ŋ�#r<<�����lPC3���gyu9W]j���@��ل�_V��zUQ1\s �:�TB� F����So*lѱ�aN|��8p��	�n+���K�b����r��%�u��:�@����1c�o5��r=���U��H��8��� � �A˧��)X��0%�i롢D:�'2��)&W�*��ś�v7f"rI7�vՂK���6_qm��Z䘪�bY��s�W&a�����(멵f��iE�ՙ���T�Gp۲��n�g^�
�u�1�T�GY��1�QD�ۮ�N����@ӝ�Hq��ـ9YQsy�x�Y��[.M�;��nmX�.O��0땬��}5鬓8>B?�
�e�)E�+�v���O��R���uQ��q��R��;�{|m.��䙯:s��+�����ze*���[�RZY��%�*8��s9mF�B��W����ed�z,�{�y��I7w���X`&F�˳}t(R���F�XU|nY��c<&HY�\8,��q;I�f�r��gtG��V����n.2��+���Ua�$��!KT���w!]�dя^QRƻ�Q���BX��1Y���F*��-;\�x;h_u10����l�Ȇ����Gˈb��3_v\E-�c��.W��'n �͆;.�-����M�zM	��Y���(��2��hCH`[^:$���R�h�Y��=Ñ`�(��ޠTla��ލ[��쉁gt}7:��wQ.\�+%��u��q�U�!.c�����c9\޶2�d3[OtFa�9��M�c;:���h�^BՒN�6��c�r�3�I}��eܒWZ���Pt����.�\�/&`�!��d�*�w]�HZY������)PO�nt�Z��d�����`ֻtQ��&X�0��BN�\��R������6	[�J.t�K��=���#�v����j*�'ۥ�&ܼV���
4^y�,��m�i�)��te@;*�3'p�j]3����B��_vK�N9�g&>��l�M�.[��sM�pWi �� �Q�3�/_�p�j:ut�Qc����ixL;y�es�������W�Iť�]��YC��Mfv�i7�Y|�=�R�x~}�'�f-�Փ�kT13ӓ;غ��eb�LQ5o�M�N��Kj��|Ƃ(�G��� ܮ�Wk<}��Z������[8v3�Ih�V� �|�(�Ѥ�nYW�dy��8��m_^Е�np�|ѻ��Յ�]�������e��t���Ԝ�ޣp�:(9�c"��vqF��᷇;nf7.�U��w۰���xqE�uk��B��U� �UPu���0�1nW8���c�4��s(͐�X�.�s�^5yH��gh���L��Ԇ���.�:���r
�*��O����.;[AI{�G��8�T�w4�λϥ���a�s�4Ӄf�K����E��1��������v[϶+2^�Mi�v�;wiݕ�Ǯ�v�n�d��ј�C#���r�j��9��Ґ��.�W��f�G����3��rc2��ʾͅ`$Cj��L�� )�
5�	�G$�#���k�WTq�^EI�<[��̽�9�.���s�W�0KFh����Xu�r�!��y�:h�3{`�)ժ��@��|��x�̍m-�CR$i�L�������]9�T]P��j�/~;R���i-�ݘ�e��x!,�+>,s�J��#>�7Ju��e��f� 
�b�.�sخԍD���u���v��hM�i��Ul�:4�e����Q�Z��sX�D\��:��K��ڍ����yn,[f�kx&���Z�Y�v��j�p�u0d���:�	�c�	�+Bs,�wm�2|�%�1AJ�����U�"���:r��N��76�����g�b�ňGY�ʅ�`�e�ӻ�1�2�8EP��W�J����D��Yp�Xyw1�ZʁU�LS9w� ��ַR8�'i�7������������ed&Y=���7����E�N�-���E�Å��i`��*�ݵ�J�e�w>�N� T��^�7��L�O\�A�,�-��풬4�oP۝���ț���h���c�n'��Ag��_3{O7&qqIv0�]hޞ��^����T\٫���7t�V�0-��ȝ��tΕ��K
�uϪ���2�W2��5g1.��۝�]KM�(����1��¦]R[�=W0�
2𿋶�'oZ��k>=+i�r�.B�d9۹<I;q�V��I���nܥp���AB�,R�+b�G!޺��c�M+�WLr׋Jx�s�%�Ϋ�~�T²��}Ͼ��h��7-8Ur�q�l5�xH/��^�Q��J��ж��(����pM�Ӛ$T%�Kz*K��>���._;7�Vۻ�y=�S#=6�[�l�Tqk�^(��B��p_e��
�W]��u��-���T��Ǥ��gW�v�hȥ�lr�\��E�lgX���ӆn�Z�e�D+�J.��5k��*��,k,��Mm��f�z������p�Ί�p��S�I�,�bvel�T��Q�H��Vz�}bw`
N��΀weΰ�ݠ1_[�,
��҃wե�B�#��(�daOE�����y���2j(�/4,Ybn3Q�2wk���m����E6V�,�	�eY��\�NNoɪ.�j���/T�n`�(e����A�'\HR��i���js�+���G��;!�o$�����/U��Q��U�qR-4k#ݹ5�%+}��s�8��Ft��e��n^Q��E�$���f���Î.�Z7wi#s�*�a�ue6����ћ���m�}���C�G29w�-.cl
*jV�թNp�s(*KS�N���̢�=Ķ��[�����E���jca,0��*��3Ұ�W�&q�I;h\	G.tlT�^�|��]Bsm���ɥv�wC�t4o\}D�HB�IX|qG��,��I
ŕ{��32���N�˓�����|��>���G�UU�P~�����������O����?s�?s�=��������?��-���Ah���p��ɐ�i��BCM��U6h�
N�J8�q�o��%9d����!����1[�
��"Mp7����^�y��o^�4l㗸8em`���҂����E]�Zp��Y�Π�-^�l�X9t��[�N�ֵ��X]˩�D;�T�����
찪�U̵6���530gC�R(Q�͛bs�w�\�d>r�G+�sC��fl9�Un�o�CQ�C�X�X�b���T���ns��i�Êl3�aPC�CB��{����WM�{ӱI6�7�r#j��3��r<X�k<�Q8vV��V��`�R���)�J��&鐲g׹ɻ�Ť�.���S&��=�&ᢖ��U�`HE�m�]:�,��UKL4���r,M1�nv�ĳ.�-���];í$�����m_��	��֬Դ��c}�)-Ǔ�|���� ܑ��U�&�.P9$�vN����
��!�y�m���3����੢�C@V;.����l �����Y!ֶ��.;�I��83]4+��ݼ�� ��0G�m�6*����ݫ�/�`����C|�^ڰ��UK�p6�ʯM���:Y--\*_���J��mgL�+��W{�&�4���G����@���]���|Ja8JU�X�|^�&I��Z�v�EkԳGNY�6<�����BOt;tf����-���Դ����݈�qxh��B��d�w�\4j !|���'�P�D�0� ��6) �E�SaSq��a}RA�$M��#���̦��StC�m�t0��6-���@"�O��-��(A��%��%(�F�X�"%3��!(.�r
��h �JiiըiCVH� 䋨$��B�H*�!��PC@�j����`�d	��Bd�YP�"d�Ӑ��a*�b���:�����J��ʩrV�L��u-��H fc@eMPӕ"QJR�d��KG6�T�CH��!�Xe��d�@�Sj2]FU�U	�dB��=:9�3��9�J��4#I_Ä���-Ư��8r�nr��]�Ad��W�K%m��{�yR�}��m:�ցǰ�FY�]pK���nA$��b� \j�E8���J-�(��`���R���Y;��%kǟǹڤ[Eʛ8�5$w�'�`�}�oW��l-S�IΘW���[.�y�l ��69��2k�w*�s.%����/�;h���Ӻ�@7��r#�@����9��x�ĞxИւgx���a�ݲ�H�{ٺ~5l��n׉B��:�Qs���{�zxz�~�s��w<�*�2d�;����${~K*W��{*mEy�3�oPZ��y�F3����:=�y�&��k���{)�� ��>��#O5;�rs_�s7|�zBa�|Խ�w�i��3�my���u���?��*��a�0�������w�}����gHu9�4����߸��n��
"<^J��O:�J�,WV���;��ͯF�zrn}�NWꊓ�U㴒�����M9��!Eyz�~��;L�-��P��4��/�|^�&V�)��;����fJ���ln�c�N�^:�Y)����d�7dG%.$i�j8ָN���Ap����d-�9Yc7/�bb���0�U�̵���-�kX:oJ��s�g�0r;��	N��7�ն收49�ծ�j �Nb�_sS����¡���)Ե^��.���~{U��|�Ѿ*YHSYV�pqo�TPek��~̨�f��'��6�����x4j2�,ƶu6Y6; �nly���ĒH�qb :��+�b]�W^��ͥ��^�p����9gE፣Yc;b�ȉ��7>>�<����`�a���kz��[`�=��Sҹ�V����k"��|A���OcM��~1�1|����wǳ۫��֫L}Cy�4X�õ3x�$g$��WpP߯{Ҕ��v����~��g��q�6UU���� ܈$Enp�;�A;t�v�zq�Q��/��|������4v�~�6k���ꈏy}���A�N�׮5��7��+;��u��%��zA$���re���;(߽Im�y���X��b��9��y�(�΂N��O���;�����T{���6�ק<\���*8��`���,)c��x6��(2�Wk��C<è���{�U ��~��jҜ�9�-J�y��GM�
��a�k��&�mĮNf�įU\�U�\1����D=x�X4s!��~���-�TbѬ'L�xz����)��;('��<J�]9�
��_��;�T��vzz�G�f߼(��W�[��=.�Abw{�lX�58x9��i��1O�v�jv�N�z�>P:�m�����;�4�c�wy@�yd���������y���C�}�&���^Mg�!&���\�ԭ�J����G����n?m!��Dc���>��A��c���>��ֳ԰H�=BN^w}��rS�}<�Ɏ-��{V�����ة^��]��Ƭx��]�{}/"_+L���x�A�-�>&#���=A�]�`�y�KA��<j'S���U���q'��'��(�6M��T�r^EFk�%my]ml�yQ�^����b��;���4�^�b�����#���z� �C��<Z9m���S����^̕���#4���ח�[���U��lJ�zOr��S�˘�#�i�N�^��|{��G`,�.#ǒۧ�*.��N�X�\M�Wm��^L��Ń�m%��������b��>�%�I���]�����i0� ��C��u,mu^_�J��f�f&�ok�{��V��r��W����y�L�4ݳ�󶚾�4��*Z��c`�ľ�.A����:�)$0-��hfut�i}�}��^����]�(����^f��+��=*x�>�44�4_.���2�r��&�4��yפ{~��2��������������{��5��[�#\����MT}�w�}��g��Fzz-���G�]o{w�p���xtg���Гa��'a�u=|�xDk��ʝ�ۆ{j*k��F?�lA��޾�5ţ�I��G���7��f�/9�wKt�r-K[�m�Ϯ��ȉM�=�9��Om��u*y��c�sz�>yy�:���J�������8�k��� `v�鍝1��� ��Β>~��G}�zo������ۦ(��Y��t��x9
~���D�ys�8e͞����|����<rFl�����0$�{������S 8:f1�O�{f�����Yc��'�c���ڊ�m�Wc�`��b���ن2TѮ>\FX޽1g-�V�����������@!�כš.��4.�#��`U���.�T8�C�~��ii�(V��"�V_p�f�]7���0k���Vn򙺝s������b��o/ Y��K8��]�|����J��~�R�^������S��%(~ߡ�F���f��Hf{ֲ���,�^`y�}�+'Q��2��6柮,��X�(|x���+�d�e/c��le'+�;����N�w��}r{�E8�'o���A�% 1)	��l���^~��x�~xG���n����ٙ�W�/��'��}YGz���'gj�.N����	Ɍ�{ZFoe�6�m�%'<d��	��io���f�>9zj26}��ޒx2j�Wk�
����t�wlw���pz��t�{ �$]o�u�'���wM��{��a8g�^���C����˸宀U�m{��\=>�<+z��1��p�A�w���#_;2p��$��tT������ײ�V=�����xC鋣��~���Ow�}�w�V�ݳ�#"!��A��y����mV� �'\s��Q-���3$umzg p* .J�p�n�pvm%�u��<��U�}�]p�5�v�xX�8�X�PA�ק�J���&ig��JƮC��ޝU�;�.��o��]�����L�?6�s ���q��»$|�]H�5=��u-���N��>>fzM�󁟽�\��)�i/(+q�s1OYj�x:��{!��t�=wz(	;�����}-�!�n���F��
``W@`]�͟d��P��4�܁�NW��TT��t�3q�Gol@�l�,8�F�y�{l���4�<[`�w��bu,^�#�V�����d�ה5s*?�
�)W�]دϕ�M�C�I]�f�oii���s�{�=[�������W�,���\�#B��9{����WK���Լ0��^Y�$�-��:݂ik�Ǫa�����>��c�G��K���tsr��"8m��"|{��$�ic���2��+�A�gA�7�_��a h<�p^fގ0�M��=����m�B��)��N7��/|0�������0�D�6M���+I��~��{w$I�Z��P��W�[F�&����l�,��9�� ����7^�y�*�ESW��-��c=8vҐ7�"�`��L�e�f���Ғ�N�ip�y��@֢�#���i�H9gs���j�s�Wh���<�G���R���U��<��%�������x��Q��<����a����	��l�qWE�>�\���t>���'�3��AcF��<�[���ۯ�t?x�A~�:��o8�*rFY����R/�̳>/��Oxaپ��M�o�󺕧�J)���֠�3o#� �c�-�I�y<oͳ�~o~�;��L��|�9����7C�`o��|��ړB����:h��k�4��&��^�e�X��2=bt�&/	G��_�v�8���ͽ��_{��~���<�^a���������z��2�^��������P�@���z�Vѕ��b�r��4l������������ڍ����r����쑙�x*9����FVx����=�o�����9/�{Qu<�o�NįN��-~^�Xx��ᣪ�.H��"��Ⱦ'��48�����{E��5���ڹJ�x��,l�bkP�U�>�@�l̊�Eu;�>�lO{W�[�Nb�#�����c7�%�<$@���Ɇ��U�[���8�(�޻�$g���V�$�a����]�H�%Ir����q�����B8`f���#ef�ݝ���)�#2����xJF\�]N��F����ğ�LPz������*9.ul�w����V;^P��mN|���J���V�x$Ѝ����W\"Fwh�6A#(ƣON5:�"�&Tg�^�=�-�]R �p����ؼ��p����*o�{^?NA�M�gח�װ�nǼW���z7�P~�*�%�.GTc����&߰q�n٫�ʷ5�,�B:�[}l��bjΝ���2)^JM��7r�ʫL�^8d�3�>9W;4�@�l���L3����˩{G��+~*�e�z=��&�<j���M5wb��#&�!�dz����u�D)^ߟ\�����7��U�O��Ipo2{�Lk���@~�!��=��"����7�f��zv����������=����eԞ��Nٯ��Z���xn����;@��rs�戴�ٗ�*u��bK�Aĉw�n
L�|�&
��[ZY�=k��[��J�[�f�Ⱦ�����,�}�8(d^V��zC���'u�D���Xۤ*?�def�ӧF���X[�$>��ݦl�#��:�S�BS�7rHl��dۄ�˽�S�.� �s������z4=Ǳ���/<v����:&��K
��;��-P-����ws�[G��s�++"���Ч�שJ��U��̛5V�z���&�o�97��7�<����ݾ��O�T;f�wx���ӽ��N�V�� �8$�c����g��T�x��1�W�wJ� ���؏!vH��vhm=a�6�i��+@{bM�E�)̞����.����!,�G+7��e��]6�b3�l`�'�*��=���o=w.�Q^�7�!}6��Sյ=���/�W��],s��W~��K.�S�V0��/�G�"<�g��M��>����W^�]/A���q@>�Y�+{ٳ~�=����T=g�I��7S��OkO�x�fW��{}�fΊ��'���ǟ d���;,�������n��#��Mn;��۟y �6a�P��z㸰J޹����ۤnp2��K�_#��7.�l#U�n�vOS����(l=����ý5p��]LS�F�b�q���ߣz槔���K�{��}G�e��e�h��NTq+����>K%:��7˄enK���nʒ�7y��E{fȩ��M3���.D V��Ӳ�θrA�6���y��=��Ӄݭz�w��$_Vd��k��ꐎ�-��p���c"r�McL�.ս[�:X�&��;������^�1�_/{f�n�M���z�/���2_wFq��2N�<H�:|=��|;gO��"/e׫���]gq���7�'�&lԚŦGYؚ5�����o-�t�/���f�_'^õ�iZ��/�U]w�� Y�+!�]'�ߨ������m{���!������ձ�yM��<>��A�����G�g����;�·��}�����-���(`����L�@�g��#|�h�#z���˚ͣ^���b�:�����Y�&OG�}1��P<~|�+�����x}�rt��q�O<���}����4^8?p��聘'���a��/�xW���^�w����>ϟ������x}�7⦂�R2���=e��ɼK ݱhEj���(ʀ�5բed����iR��pu�ُ����P4L[OV]� (+���K
Y����S �C�*QQ��>P�YH�D����b���'���B�+Au��V�gӊ&)�PN�ɮ��AZ�t��h[���6=:b{:TVTL�j)H�zW9����J�w�s���0����x��g,���ܴ픰�y��+�[��I:��g:��ޢ�6�7�5 
ws�ݫ��7R�*c��ӹ��:l�c	�!ηٻ�d�z�C&̮�Uy�����.�G|�z���Nv*�f�g�Ԭ�\gi������ӵ2��1��s04�%�^<�˽F�u�y&�"��'^�h�m^�l�V0f�h��v��2�:��]!�{�(�{V�fEh��F&�1�%�
�)r2��Q�VN��Ph"!(m�GY0��aWf���:�l��GE1|�Z��Y{˹�P��R��ȫ!u�*G��g��wz�����$��[�3��;d�K��[:�&�`�S��N}|�Xj�X���ꗂ&P���}³&����n9ݝI���r�r����;D��W.[���2������o�\d�Ψ)hO����U��d�4粯�U���Odf�j�u�g{LBS�� ��滈��ܦ���LB�����0�y7U�&�s�ܚ�:.�n��.#�������@�,�Bf�C��Ĭf-�1a���ko�w�^iB��O[O75�-���#\ݕE�E�Ȱ��fg�~�O���^������g_�ߦAk"�ܡZԩ�b¥ _�37ND�ol6wu�Y��=O,�١�Q�k��çE��f�1`��+�8d�*u�>�rT�	�f`�y�U�;�Y;�J�����&7kBawV-�Y5J=49yZ���{E�����KB����8��1 d��u��>.�`�ux��f^�XٕG�tռ�6�u8@��u�֥?��L���,���@��O��ts�j� UƊ�����E�/1V�2uT`��U��6�nI����m�}��W3M���h�1'!�s�_0@bΝa���B֭�.(w)�Ao{wg] ������.Z-�m^����5��@���Ń��lؓ�wT��⸗/��n��k=�at=y}y0�	��(ed]��)GXVϭC{��V���IK!�=Yj��A80^�Ѧ��h��o2yo%b�ζ^e�c(^�8��N�dD�ʖ֮M�|x&�,��K�װ��c s	�����
���J�E��K[��X\���f����#�u�������'q�.�|i�ب�\"�4�BÊ��/*v_WQ�ڷT�������/PN�EΎf�q�k�r�k�;ƃG�̚I���ט4_9(  8z�o)-��*����ƶӧ�=��]�{��9b�rv���o�]�2�u�aw��t���y�)�z����> )�P�K0K1� �*���K0 (�%"@��2S"�Ȥ� ��%rhb�������
W,�C!�
ZZ��%:�LA��ɥ�2b�R����3X���բb�R���jֱ����	���f&�����4NK�ֳ�5�D���2L�	�fj0� �
�Q���Դd6bd�Ɠ#3���2f��(ri0�"2i�$����2b+2�3$�jf��6FVe�Fa�Y�XT�efQk1�c��Y��Y�XY�2�dі0�Vju�k2a�Y�ɵ�deDZ�k,̚"��0��s0����*�3���?|H���?wٚ^,��s~�ʗ�8�v/��)C7L�:b��OMr���:�]Lb�_F��j��J���P�Re��|~���v:��d��;���it��9�����$�hH����/�6��i,�xU���>�a��n����B�Bi��=P�z/���摛������v����Y�;��伙�o]J�k��7�iᥡ�X	i��Қ�Nbc�_/f@ƥ�S7^A��l3����w���Ve\��W�{v_�2Y^��(��p�0z̅k��C���J��3|'�#�Y �\��"�x�t��D?��b�<>u��({U�_Y�+Ƭ�P��9)�ΦGp7���rN��*�]�m����b���8��Y�$��\�I������Ο=N|ҡ$8��x�\}Ss�t�>SY7��GWf�`PZA咋��N��s�^��RT�ۄvN�y�-��te�4��>3zY=�����L������A�f
�W�@>�J���NV7H��y�5\	=n��Kln��R��h7���+�!�� �#��Am�N��覔�0�vA�M�����#���NR�y�q�=շI�3H�B�f�D����c,s;��q�,����m���\�~0�ğ�דM�������_�_����Kv�q4�=�n�6���i�v�׷�J�wTH^���1�Y{yԎtξ�KoR�g�F�Ì�
!��ݼ�y�T�������T���C4'&H��K�
�L�&����6��.Z�a��@������[��w�"�ybC��H���_à!w$O�{'P�urdS�ޭ��U
h���aTu�i���{�M�s�R��|�U@	��*#1���#��<��� p��9t��dԭ����}s��+��M��Ʋǿr�7��_-���q������9�P~���T�糍<'U�Lm������ݎ�;ϵ�hGVI���i����ԔT�M��^ÿ����6�Х<�s:�s|`��ap��r�3���w<�p�_O��s���'�w���l��m5PוY�(�bO^Dy��3eg�D��c=��LL$��=8�nply�WF��:8�7�������,�ܘW���6��2�M��hr���킒x<ğ���g���W>��ح`�U�7-n-��%�q����#/�a���	\�ԑ�g�f�2��l��$б��]�	E�P:>�8z��e�b�}� ��Ƣ���]�d	c^(��@���5��sn� �[z�7�vq��J'ct��R]�ڄD�i ��,���D ���tB�B��U�^�����z},6mK-ge��\[�<���	Z)�U��k:�����`C�+��<�'7l���%k	����&1��0'{�r�[�𭝽�qS��P%YKUɗ;j ���#B����	g��6k`�(»{YI�c�(�����a�*B�=;YyʂF_���n_�כ�
AV����`����&���5�3p�_Jb�:!2N]�9�R�j�QO�m�l�fqz8��%m�u�n��u�d[BQ�쐄cL:A��ˮ�n�2��I�.��nZ7����k2����Ce��P6#�˴���H�p0 �k"��:�xK*U; �J�^��so��v���:fT�#OH.�b�g��q��X��@+� ����!�T����z)9of�
s�4D#�[�z�_5��q^�wYaw�w�U��RX�Gi@�$�k&� ��F��g2"�渫��������!�\ǒ�zMв���U�]<�ly]k	OvZ��À� ���^g�CW��}�y����[8.X��9��C8ȵ~Q+rn��S����T"�]by�g�V����Qq��й��k}�8?��AAi���\Н�d��:Kj~O�X�9C�����cZ�px*�].Szk'oj􎶦E@����s&D����ȉ!0���~��vI��z]�Iopb��T��3��A���Q.��e�c�H̻H�`���\d�B�	��3������x��U�T�n��Y�v�0�0jND�-Yi�h��/6����dZ�<�w�h�7�񉛡v
̞�D��Zt�pP�R�(�e���ݕ9�(�%o{��ɘ�X��|����-h�����k���QU�4��+%��`NPf�#sJ��뚻{��y/���]�扐Hz@A��K���-��*���DE�<�#���B2��}u1�R=:VuB�t&���as�ٰPyja�W!
�y��L� 鋇U�goM�lŰ�VZ5��_k�eX/P~�軚Ǳ5Բf��!7��� ʖ]
6�����x=�ӝ����C�UWS����v*����~bW@���_���-�^�"Se�,R%8�t[�����+�Fڻ�mr-
C�w\
�=[�M=��	��L ����HM�x��_)��B&����Y�Aˬ�ͩ[=hہH.�`���c����߹�^з�x��A�]ICÍk_�ʡR{�����m��������9yb�I�Q,���Lk�*L^y�=��p+_Z��1	���*��ӫf�u�;p�b�"D��I�s���UJ.��	c�z�������ձ�B���f��'�kԂ%���U%�G,c�;���4�Rq¾���������L?5'��{�6ȋ�f�*�v�E��a���AngA��'f��f�����*�=��s2��_|~�O����bۨ/��7ˮ��1<���m��ws
�p�s(�tRr]��{r���6vŭ�$��n����ݒ���P�ͭ�6��)�%�L�vK}��VY�	YaMY5U�t��
�A�]1W�F.I�'4�L���5�\�j���bP;V���}���wY�H~���.���
�tz:�����j��-l�G�[[��פ���ʥ��f��,���+_�u	�������/�q{�mpO�!�q�׽6ɽR���@�f�7����n�yk�>�}fz<�=��v
>�y�	\<�z�.jr� +Nyp�ȡ!�Uj�S��׹����!�ϖI/����!� ��a�h�`X����x�A�xG)8ޅU;Sf欭�g����S�"zV=��k��4�����E4x!#�S����tEC���[.K�!�5;M��S��p��tkL=�O^Tg5�h�C�	�n*f��Xux���#&;y_3b���ц�Զ��~�q��Ì�Q#�VDč]�/�:*��ϝm��n�3:o����"C�*���O/}iȞ\�Yz�m��/ƙ�+�dQ+��_X w���}::e�K%�{'ӕŪ3�vf����
Z���ɩb�Oj���¼z/��[�z��xA@���+�! �H�* �+L;��)x��Rd�q���%�t�K#(�k�";���ɲ����A��������9����uהp�-�=ߤs���,��K~8T;��:栯����O3[��!R�R.��"������Z�:Y��:O
4��-����<��W�D���]�@|{T/V��s�O��[˰t��o@�oU��-pj#�e9]���:8�.O�C�u��]�1N͈K�`k�� We�눔�8��4�7�8�=�&��#ry��.7���&/��U�ۭzt�@�f�b|�3tlǇ�e�+0�ƙR��b)9C�I�b�o`3	[�s����k�λ�r�ϑ�>{aA#��Bm�;<�:m��Z�.�Bn���-?'���وR�i�L�v�У���灩t�=�����i���(GD�/f�i��U�m��5w+T��pL߻��"��m�#]�k�$o�&+S��#�!����쟍zz�s��oĩ�v�tn�lW�oU��*R~k�o6�� j��+�v�;�
�c�w�=W��|�y��Eu����i��]NC��¨Z��S��5�?.�Nq��b�a��B v� ���	�&}/�8�{0s���i�oM��	�t�C4Ў� $���i�H@;�%Z���:` a{�M�v�v��[�������	�D�??e?>i0���WP�~ޯ�aΡ5�f����1`����\����V���0�
���A�p!@`���+��vq�������3Kz��,xF�A�R��c�Tڛ���4C��*wl����\C%E���9Q�ڛD0y�|�gI�w��N��wn��Pr9����0w%sB��^�����ͦ��/��]�O7NÊ��n:���`��;!�2]��V�
o��3/�hO^�����ф��<#���v^Ju�0�*'�l>1��M�ղ(��&|�@�F=�}\��iT���p���۝��b�C�N��rCRFu��G����px��h��� ��q�I�Ԏ5p��S��{Ʃ�S]^��V5�'���'+ K�����o�YQp��3*�����l�6�O��ݠ�_陋������-�2=tB��RukU
V>�7���<��;��Ό$�3}����H��>)����	�?ߑ��a<%��-]�'�)͔�Z]­�qU�z��������&Er�p$sW���q�A��{f�C*��CH�2�#M*L��S�LtD�����k�!��� �Z�y�H�@�Ef�xa��hAƘr�zzA��`K&��ڳ�2��������5<^m)�M��Ӌ�F������� ���!�T��܀ow=SI{]Z��o5^�Rn�08�0��+��\��~Ib��0�����C����sZ/,luD�a����q��О�.`Ԋ;�2q��RX]<�m]k	Ovl�R���)�y߬�c�~�siC��1E!�,J0t��L�Vf	GZo���b�͗����Ę���=[��0w�H�����/��B�W�~(�wm꼥���l��*Gٺ��I��shp[J�K��S��M/d�im5��0IG�bc;,A�P�>r�����;"������5����i�W��4�|��s8NX߲��7V�i�+qܟ�kߊ�^���k��c�'1�u>p[��B�þϔ?���lsL��;.�k:�j���&�*���ӽ�e���SQ�VZ�N�KK�z'���dרT<���}�Px��뜗d�Xޗnol�BgT�C��a�b�9c�S�{��v=x��iD[��_Z�t>�yO��oZ�r9��z�I�߶��g��sCU;�d<�H~*��].�C�.x��8��q�w����ҹ�qr�oQ����/E�\�5�m~͎硛	��0�z ���y��ϛj2�Л��7�[eA��w�{��Ԧ�n�\�A��!�q1w5����=�R����B�a�RˡY�]s�oJ�呱w/p�����?w5��K0��,�| �4��M0�Ɇ�.�lV'jc��]Jm�1o)ig�ku�&���(����u-ï%	�^��B�Fc�M<6��;@@ߥ�S�!�Bo��4�)���}7ʻEFU�z�U���^'��R�tR�u��_a�WPW� ����=��<8���zq���w3J��T7�����y�V�A�~>`Ъ��d䮸K�]*��[臹��Hu��>ζ)��(c�{�A�Zd��3n��t�QnY؄B�ďrGNJvE�B.��a&����Q�,��|eC,��z�*��֞��4m
��2LPΈi����j����V��q�U5y#��N)��`�YY�x�5�&���!>{_Z��ޓ.����Ȋ�α�^tچ���1C�*��w��酎U(��x�4�Cq]����dB��#�?���z�
�;x'd��d�G7P���װ�
7�4��W�*�z���&rĮ��$r��7������mg�xM } @_r�ZD!�S�E�ɛ`Z�+R�Vɇ�����*j�56���}N��7p�[4�>'���@q�
�@���X��("�FĶ������*���O7^1��~�jձ�`ޭ��a��).����/)�|���!ot��x>�4u~1�Gq �M0�FP�&ߗv�������B;��Γ?S��N�1�ۖcF,3������p:y�/�]�zCsf&/H��9�T�n��?9��ސͳ�$�X/��"��"�t<�l��dtK�I���Ge�r��b�Q١[�q1*m=���~X8�s9���P�z)�!#�S���>�f�y��.�)����F��)���� �1��՟ߕNw�����i�h�,:�YA���zY2�m���e��6:_�	+OL������f�zL�{ב��#� ի퇽	�d��q��Jv�2�	�sKdb�ȣ"���Ya
�ϭl��>H� dX4��DU�(�{�V��&l0]\��.��`L`ˋ8��N;(���2��E�����*�v��(e�f?öo�}�6Td(4,-��=��o�^b�~�z�8��R�noI�9��c��<�4���lW��g�=[®�N�ŵ�E�3�>�V�I�5��Is3�U�pfN+5/��}��x@ؼ
�2���:�r�Ֆ���hYd�8r��s?aƕ^��ڵ���i��#x?�k24P�5�^���(�E�%4��(�k����\2,�@]���1���;$N���c��N��WO��`�D�I/])�r�	��"��F�[>�s/r8N>-!���z�T׷$w�|@C�5��K6����a�`�̧q#L�����S�A�`5�����\�$C���u�=�T�L�J��k��p8G�9�hN��覒�.�rt��EHN�F[['�$�Fs�o=��y=./#�t����y�c,7�݈�#bYs�Ϫi��:�;N̲�E&�2s�����O�A����}ʿ,Hw�H���a��<ò~3U9����:����k�뮡loЍ[^�$�ֺ:�P
���k�+�|�Y�������^��OOo�߷����}��o����(N�����1s��n0�:�d�0Q֮9/�B$�ƺ�:L0��ՙ��$��2��ݼO4@�X�/;r٘��u�zpa�W�b"����Y�WM��u4"TbŻ��YS�Z�=��i��6�9$"�a����컲JqKv�o�l'�PţXc�<h�$o]js�O�R-=�� �88�T1X��Ի����"��P��rh�o�ť=ڸ+7y�p=�\����u�Wu	ِ򗽂���.�#ɰB�����E<�Sr���m`�h�H�1�A�c�6��
�ڽ6���j�X̭<C��n��9o4(����疓���ll
[��*j�d7u�%�Hi.��.1��UJZGB�<�qϛ�:�t76�i9�z�,ՙCN��%�[��mv���Uܭ�mb�Њ����ե�E�s�$���G^e�P^��Î�@)��(ٓ��K�b�j;F>WK��Tb��7_�z��F��s",�����2�@�9�`���8�E�K�)�3�3&r�6��jݛŽ�Kv^�M�Odҁ��V^�V�=;������]I��j�G]f	�*�,�Vr8��#�5e�q�;2хPs]2h�{���I6+������O�e����F^r,wB�2j�n���e(���<K�����k�(�=˒���+M���M�b��o��>8Y�Ciis���5� S�RN�����	\�,���W�K�4���C�z�����ݭ���8N�$���������K�Vb��
��yK��FX�a�V͢����ǂ<���'��a��s�'�#^�Q��`�S��.жS�FTwc\7K���grV-hV�e�����ףQ��t�Aɓ�A��jn�J��6�Oz�S+t-�5rڹ��]����&��T.f[c����EO�m곣[j`G.�0�
�Vux����x�)v�}([�[ �q��p���;��te�8�7c�ۋ�ר���%0	����}�a�=Wa��!�g3�c��*b��wx�M�Gp��R�1�u2N��\�%�����92����.�`}w �i��1�N�,��;�h����w�sP��]��t���[rJͷhQvFO�mqt"���*������ʷO����n�o�:�vvW=&�Jn#i��wl��k>�خ�Th�i����9x�k;O������75:�Z{�f��ٰ^l�w�a۽O4Wh�h�}�u�DK[�m�gwOk�6�~(��\�����b�;���6Ti�/�U�$�����r�z�5�[s%n�bsH�gK5�;_3[���%j\��]3����ڏ$΅ö��n����hY߶�+m�ln�c����O�GǷn��6�Eo�}f,�+k�[�l�t,���C�})���Vo:���,�����j�'yQ�Me,8�����\a%�*���2���e���.J���I%�$�C�),��2]A�U�r���*2Ժ�e�Xf��44ICTfeM��A��i�eMQa�6bdSA������f1k�������TU�ʪ����f�PY�R�U%%)MEQD�EDP�F�Ȣ�)���*�&
��RdE4APIIN�%�9QEQ��A��afU	LE�3!LEA4A$Y�5�AKM5@EHDD�ET��aIQ%:����(&5�U��S5D�EVe�UTD�5RUD���Q3dh�T��IM�1T�PP�Q�L�F�>h1����F�A�^���X�v��Ͳ�J\�>�.noWo�RK����hr��"���u˗��Z�Y	,f��}FZ�Wo6 t&-�a-6 �E%2���� ������ʎr}��:X��͸P�\����⸞9�z��D��,}�}Zf}�[,?��C�\�k��6P�#��I��L@~gA���קa��q��Gp�I86��0VBA�	EO�F������q��"�r;��!x�<��r�y�9��_��?<�Ρ$ėn����ݎ�$�a�[��O$����_��t�S�K<%}�^��$������q�'e�Y�j��s��<e�ct7^�Jf�8.�N�T�p��{�bE���CL�^�$�y	��&��["�a��Ļ���ƒ��v�^����:� Ũ�����g���U�\2�%X���?;�Z���ӛ4*.�>k����6���zO�~�'X��(ֳ׌u�6K�9�w"�]��[]{=q�{uj��
��'�d<k��N�j�����2���):��P�j����=a.[n�z��&�㾺V�U���ޅ^�L�B^v��n})�s�d��D�>J�r{Uf����׽�Hm���v�@p'Z�][.}
G�q #�}ruñ޾2�^o��ɬ�"��R��u���N�dtq<6nK�\ug9į�$4nl��]m�٤�����'�t��GE��كx�Q
gGƪo^�!�3x%�����d�G'�Y�i�t�;]�d��LV�s4)u���P'`u׀�������uޥ���Ћs*�m1�����3�o7�8�{U7q�N�	���q�o�������td!�9	�:��od�l��=������5��K��^t�1�#���lH���5���:d�p��p������-{�Uܜ�9�P��^K���K��̮xj���^l%�y�a#S�vi�Ǌfj�E�U$�u��֔�N�2O�z(��&�Yc�V�*�
���f�J�����ܜ¹RSF�1|��j�8u.3���^bŬ@P���9��q�j�J�`'�Z�T�ȧ�9�\r �OZ7Ԣ�a��G2OAܗ8?���i�����춆u�0�@��F�g2N3C[.޹�&���).�C��/T<k��yx�+���p�
�����om�2�t�����=ͯqY��ӻ������.�	�nǠL˴�l[���9�߂gDau�'c��3]�w'�vV���F����N�=y��2	E@A�r�v�l��ohlk��W��ɶ�:�+G!K�#����<�5�my���f�A�Y�׊�r3�ی�M���?�N�/ñ�D��e�n�u�!�w7���n��|�>�A2&ZzqC�9�/`�RP3����+#��#q8�e�D�n
ٱ�Q�G��&݄�}&:��_��ۡ�+�/�KO���V��%��,�s�
jC�u�֞N�G27RJ��X�o�;��SD[c�����饉'j喌s��?�g�`���~P�$�K�OnUKcR�!s�t��Q��0U1Q��ʻ˝��5��� 5ڡW���p����|����ѳ��D&�=�Π���4͕f�[tX�S���K��]��O���eb��\Oʘ�=��P��i՚�Oh�������'�/��2�&��`FKf��+�,�9�G��O��]1�&7ތ����]Ih}iW�T�N�<2.P���6Q�¼��(=��z��ή'^k���M�Y@���TA`�ѨA�"D�2��S��@r�E�s� Ɩ����-�o�j1<���oq��A��C�i(f��Btt�F�F������z_�����T3,v�d�]�uΊ��7l�ĸx`>ϘG����z8F�Fė[&m�l&�V�*�>�9�^fR׺��q�-�U���[R�^Y]yZ���>,_4�]@M�w��Z�OWD^�����&Ţ���)`���{	A/r�UԳm�l���P(x-�a�ϣ�'L�qV����Y�����
�@'A2��C��ގ�s�*,�E��ZG'��xH/c4P Q�8�wo�h7ېky-8��T�y�Lx�q9�V���=��j��xL����a�&���ٙ7h�tQ^NDk��0�&b�3Vq�w�8��m��4�Y����x|����q+w<���É�eb9Rc`'����ӯ�#��C1 ņv2`3?�A��
����d�g��R����`�?!��A
{B�Ũ�Yx���H�v��x�yb�X�c�IZ|gB��Vݾ�]ugG0��Bæ�a�θ��e�^��#�3���
^��^)�!>����ې�;LM�z�N�S.!���r���_p]��D���q�����編sNn�k�K���h�$���6�F��L��Q���:a�_xo?�``�(|9tHM:>���t��ˇ�8�����i�����Z�Zֈ�s��]���K��h�{"�_0E�����Z�x)"������y�p������HJm�2b)��t�
��z��x/^��t�̢�a���U��շ�K�鐈{; ��:�:!�D�/a%5b{��v���b���#�v7�S2mM�*Q���us���Q)ٲ��&���$vI/])�r�	�(ܒ4�۸NF�ѻ��ո�v2����������cT%,�^�����6e;�2�'��NUz=U;Ӫ�-�#�#/�mv{�#}-r�y�,(�d�u
�Ɓ�X���q��������>� ���K��G7>���[�.Ր�aւ�8LD��'
Y�>�/%��I?]-j�ak<�%Tkfm��������'c�VS�22����k\�}�]��}���p���j��ֻ�\��ߚ��}��+4��� lWy_��9?@W���,�3����h��{>˅�{)�G"�.�ؾrp'�K���9tK�������G4Ñ�$k�.w��b���ĥ�[�����R���ZcO�����/���$X���?c��2�U��(�O�4뺴Z�΄jxK�I��@�j�����׈ɷ�Q��bb�b2F(j��%�`L�����Z�
��;'%����Ȥ��S�1�e�c�O�l�W2	���f��9v\N9'�<�b�c$������tz%��Bv>��4#�$�1,y! �K�ת�t����T�V��[���5��`[�r�y�19##�6Aӿ?=�*���D�t��[UnlF��콦Y�O(����v9V'��"O�A��|c��z���>K�rE��M�m��{3O���i�k���j�S��W#.����3ez�H�W�y	��8>�}B�*z�q�|�5�l_C�mA����_R���ֺ
-?-�\����=��U�-��������ݔ*6DoAnL�\��H�R�0S��P�Ik�4��9/�Z�V��_�mA������B�L�'':�v���ce� ��vܨU��y_F䘞e��l��@$BR�:�lk������}0���hųS��I�9+�ѹ��N\c���}�*8��w<���
�#��'����]��@oA	�� ��@�4Q�g������5�4���:&�w1yG�=�����!ԩ��9��45.����XZ�R�E��;��7g�Uw���B!�;na詯`��0 ��(2�t%�'j��n})�W�D&I�Av�i���S�k7k�;e�a2��u7�*�"�d�5���6\}#����p"V/��v!���{z�ͻ��ew����J���y�\h�t�vl����A�v!?[EԿt�D��4ɫ˜�]��h.�L	c^���Fa�I�Sm��y�0g�0o��O��\�4|�j���~��Jnk�ܣ��v����x�9џA�G(Q�4�Uz̮xj�r�͂�����0���ͫ�k��V��wm�;��;��:nD@M��z+�A�t9��.��,(Z��3`R�a��Y`�ft�YK67#�&��d�'�#���b�(Lc�sn�8д�����9&m5D�H�r~ث���^�	���X�l,�9�`0 y����s@N˲���><}�����ח��GLr�U!ߒB�՘enK�m���]p�R��ww�x�m�AG��*`e'��ʒ��rˤ�Z��W�aܕ	�Q�-�1�D���аa�mӭh�{n����|�-��3��� �䦞�a�1�/�y�����>����� �@���(��^�����w�h�����;N�&����/E�3�끀���N��w99*�c�Ѭ���-2�V��1%ډ�c�^̻O���5�l��k˼ O�R�|�B=%�����4�K�#nq�`��/�y��<����D[*�x�'�`9k�;�7�[��l�n���hL����7>��5��4w��_��W!
��;�
���mjɞ�sF5�5���mr�S
��:�Ϛ9��Ô�D]��|i�U-�^\�.{�2|��R��)�n�y�\.���.���ٲ�N:�G�5T8.���!�Ǳ8�NTda�P,I�Mً������mp4ր]#���B�ܮ�`��z����v���iO~j!��Hg^�^� �%�����99��5���:
dJe`�Jsc�=��]�r٬8��VY*A�k�GN����]y���J�zH/����v4'�ƽ�!'\Ĳ.���LJ2�s�W8k����مpd�H�R�+e�j=��H�f��B`y�c�@��i;���Rt��ʥX9��z��<�wV�y�M��yͽ7�&[{�����eh�=<M�@�붎J>�7g��eW��^ߴKG/��l�@�����2��8��{;��뗄d�R��es��{������<����K�s!2R�̰t]<��;f7�)aU�w-#�J�`X�s"iƸ�`���}��~ �� D
�B*� �J�f���N�f-u�yo�������!-�'�&40�
7�4��Q�]/V���,�g�Nə0V�b��|�O�>ZԻ�Ö��\:��G�-�"8F�P��.��L���'(\4'�&��i��q��ֈ�3����R;����E����qHG0>��8u��;4ڙnR����������-lP����Z�ߟ��+�ό~���s�N���s	�#��X�w��+-��5i�񐍇d^ʊeނ�1����~�>�z�3�@��1���}>��mgmAw��n�OGf�z�ve��؜G��y �H�����ID�x��Ǚ��VY$64�H�֪+���v�89Fp�$��\9�/����A�l�/���S@CKML)��{��x+]�z��?H�T�����/D��k�!��Bu[7�ݧr�5�w�<�ڝx֏h̀j_�e�r����c�r�A��N�*$a�(X|a�������/8�|���"��7]�ר[��H�7-��ȅ��PH�A�4�+��D�‰{������)�q�S��o(�"bgo��,`Y��*ECO'���ߠ'��R�h���N��'�HnM֕�$���t�d"	��D��}f���ƇKs�o'��qF�frk;d�z�g���=��X�#��c:�ֹ[*.���4ݽ�^u�{<�>�5���5�]Z/���D
JF�B�B�B���B�Q)�9������5{��y[��3r�����o�QR��7���|�L�D��]:��վz���-�܀y��v�����*PǺ�!hX�`��G�}������!�y8�d_�Y4��(�k�����	]��rV��\<u1����I?~� [K;�F�a��щ��"B��-���	�~1�j�,f��W)���ץ�ݍ����E���} �5��ۢvx2�2�ٔ�$i�Z�/12/&�z�l�u��s��y�e"����b��|�>��x���o@r!6���覒�W=j��b̮�����.�o'e�c��J-?,O ��j-#�.�a�?p��8�`|����\7U����C3$e^uʤM���曯	�k��Qx��F��n���?yI0��0�;�S����c�S�P��ʍ�%�ɑLk�M[]������FM�ߕϠ�f�طvmt�����Ⱦr�n��[ܘ2����C�r^��?>��4-'�ø1�e�c�N�����W5�)LQ��V��	�C��p�/��t9?2
A��}l/Bv>��4#�a��Nf�r��hq�����c3�%��FͲf��(��`�ybɖ+w9�/�V���ΓWK�����B�r��C;�[�ғvl��h�*��0�P2��R��mb��Y�r.fP�ҳ�f�����k�yFj'�j뒔�퓘<�A�������<���֜q�Z�<��ξJ�� �
�J�R-Ĩ�R
- R�������Qx��[�	��QE�?t�<l�T0-�q�_�W3��rFGu���o��W=i�k�����{�dJJi;R2�ZG�q �/��sdK��Y��D�����k�<�)��YYS�o�9kq{CT�/,�4״��j*q�j��\dW�l�P�Jc�OK~%�T��Ebm�͜�'�,����ϫo6+Z�a �,�X��AFu���6ʽ�-�;Ү,��pz�+�K�Ů�-�/p�^D>c�~��	XڊƯoA	���a�@�5�k:'�����g�l�5�wS=�k^i�����͸f��X�N2�'��˧Y3�}�,{�(���s�����Wn�͔&��,)��[`���sB���D�yA�k�%�'j��n})����M,5%�Q�Z��_��_�IP�bU��b�u�4.���	F4äLl�F}*���U�>�����|/:]��Re���_<�/@�4�M��\0�ǖ�B1�m߅��kܙ\��2��w�8�SꞐ�z`K*���lԤ�c��"�<�4�4���\���Ͼ��|��[�����������������Ѯ�n�;+�]i�{��+D56�HTs*p�MB�s&k��%嗣�����go;=B5�M�m��*6���b@䝙.���&���go7�qv�����\q��[YYvt�h��PtV�<�,������ͧz��V���0dnԭG�R�S]�\�^%�`/�8A�G>��;gCS"�VwH��Y�a��WN��{/rܩz����QU�R�D>�W2�*n-D)J��Ӳ1�"I��%5�\G��/.���;�퇬+��w��'3��{1��N�����&˔x����\ru�ή;�e�
��4k
������b(����A�n�~Z�u12��S �@*�T���Mέkwdz����E�ִw�Y|u
��sW���3��p� 3w7h�M�oYI�Y��!)�yF�0,A��wJ>(��f���E��d+:���a���	4{=X2��B5ks�{�*pF'k��Sj��U�7W�i`źW7����>����5�k�{�m�ߵ+�s�A��Cۜ�'�4d�9������θx��>G]��NL�ٛ�C �?	,AE�x�)�h��1��E�$�;kuͣ���]�7^�l�؞��cU�M�,K��c�QQ���}mI�.��F�tuJ�!ɹx�w��!����֔��H��=���y%sx]s��h�R�WWa,^�����Kͬ	h#�v���f��kr�,�g_���8�Ѡ�4����T�;�+֪:�ɟc|�g�����!=�GJԮ�(�~�s�g�<���|n�`��%�)ݲ��؉�}ћ�`��`�t^���'z�u���\9o1:/+�R!LY�[�[7�9���t�a�n�7�ܳ�w3n_X1h +b�(u���cU0�[�gjL��`���n�ܮ�uu2f�:t�5�U�m"�����ԙg��r��)�x:+���G��F1�8�9A$�):�|���WP�(�V.�okO\�S�hy��G��e��h��\��y5yU�5{Mfp�b�%f�i��o2�?ǖ��!Or���vz���O�;ۛBȎ�v`�&6��M�����t)F�Eq�Y��NؚlS��$im���	Β��}�{u �^����s���hζ���)��қn�oe�+Vi���2�	�c!cauh��H�6�n�m�uvG��҂b�{rЈ.��w�T��$9o}�N�i@]�����ʥ����6i4qjXz�&[�56kU�b�v�X��6P��ˣ�;��=�Ɯ���u�����CX�e:n���!�Ϣ�K��ܦ� 뵽�
T:1���~���kK'��e�H�Ra���04���p�p�vyG�V=]2���|Bޔi<St�p����kR��}D=W[�9:��a��(&)
�}i䏰U� �RӲ\��ݎ4]`��k������n����ʝY( @$��E����((b���"�3( ��������� �(jj�(���
 �` �*&��J"*��������j*�"&(�	������&��ʢ
������������b����"�$������*�"�����)&�(��l�&������I"��12"�"&jH���()����
�	&"&&�������"��b�)�����**���8K$�Q1fQK��Ya1�UMc�e���cSfbEQA,�dME	EAEEEQQURLG�H>��+#�װ��R�kVY��Y���ǽZ��s{4���]j�!�
�BG/1cq|�ፓ٦TR��y��5�sמ����\�!>!U�Q�@�X�Qh�
DQ�ZZg���~͝�~p^E�/�!�_�T������H��&B̮xj�r�����6�V�cq	n<�{V�h������MyDЅ�Aqx�u�n��s']�����c2�f�:�i�39����t�ϕ�\�Ó_~V�|�OA��������t�C8еn�c��f}��m������������Alr{k����Q{�"��(~��~^�6#�s}�C�^�s_*6�ޚ`Y��
���=�i��5-����z/a��2%��:aOcF�扳���Y*��2�����t��,+�7��Q2�q��̻O���<���חu<J��lr�l���,�HR����yO�*6���v/"�y� ��Pi�]��D[*j�m��rKʌ���+6�քAc�O~!���&���+_�l$Zˠ_�W!
%�T���껃6�����20m�PS���!o�`��ni�%��:��oH�>�q=[�D^�^�M���HjA�H�:��oL"ڍzƺ)����h>F~����Xt;4eھ�j�j���L�L�T#?94<u �Fh怚s�uǕ7JR�E�����w|�է��
�;���R�p�P�����r͵Ȭvs���]�(�~O1�[�÷���73��h�����g�l#Vi3N�%�%h�)Ў�R1�=���着��T�@�H�(����
(P҃B����1+J�@�@����G�5��^��r�-��5��!2����i��K�1��{gb�&C�Vt�8K)m��\pV��܆��^��LX�>��%5�xNx�LP�U�FNc־��z��w<+w��zn=�ϫl!��C�/�z��hH�5�1	:��d]g<S�F�
�\�W9˘�Ǌ;{�f��ƽ72���$D&���1��H�^�I���:a��Q���w���|�ml�ٓa�w8�}��=	�jÇ(��ѵ��ƀ�t(��I�UU����f�i�c]{KDu�Y�zd�ʗI�栜K��v�s ����zz��+���K#�*ԫ�X�їI��n�L����J�4�̟R������{p�9{�@�����@p�_������^�d�s-��M�OW5��!*���esߖ�/r�T�6w��~��0A\9�S�}�����w���aM:��Y�ݻ/L��I�����c��u��so�ܳ,3��|~ǒn-ڤ�ɷD�؜<�2������|��O�3d;l�J/ş�C�v1^>o��ib��L��û���Mu�oQ��X�#��k+�	�kIO��|���^�f���^o!x.#zOom���Pnt���ҩg�&��&ݕ�Ӄ[�,���l�t�[*�C~Kt�n7d&�����:h
�aP[���-8t����Ϛ�gg]�|� 4+@����!@�"P-!H�H�"4H�E")M(2J�JH��������6��{�� �5 �����~����!�"T�{���Ksg�ʟ�Qh>Z�Ŵ�l�jȽ��]̄�3���N?Oؕ#��68/D����D�q�j��m>-�C����7őSUy��F�=W��K��,y��0a��E'�y���y����1<9tH�4���;c��7��jk;n�}�㎆��1IK6�����'z+��@��%񯙫+��D�"�wǋ�P����b�ݝ����BU�;�mEz}�����MK�{UӬ(�ǫz���\E�'�U|&bҼ����\�!@��"%�� ����Ed���_�O��$��\�I��b7z�i�:��ȩ�=�~��<��TT�d����%ٲ�SI��� �$��g=WN��xO���
�\�u`�nGb"��܆�.�I����b��X����`�f����p�0SfS�YtrBԢ�6��K2��=�s;Uc�G}	o�Ȼ�U�9�^�#ϲ�-� �z�	��'g�s��C_�}�췷�Y7�>�m.�L�O�Bn�����	�������L"A��ь�
9�޿?��8M�ul=�.��q~S2�\�xT�^M�Ra��.�?N��`F�.� ݽ���P�����oW���H���v��h�~���|%nԳßpHĳ�g�V��6w�ѺM�$��[i�;���:������֜o:�m���#WѨ1�VԚ{���)Bґ
R�R,ʔ$E �#B*4�(�	E�]w��}k�^{���%�{5sLo8�5�^)@��~/�����<�E�xQg�����4������=�1	�au�Ҏ�<�D��ɚj�����O*���f������[��"^�׵k�ٶ]� C�:O"��z���C8д���5���]>���0r������il�:<��h���n�P�����1��W����:x�!��|·^�E���R�!u.T��㡞���#`��`��^��3�䌎�/�P�"��tw^8܍S��9t3�hMy)��C�����3���ʀ�-?V��Fh���l��|�+�v(�veh~��̻ױ�L�e�oG��,�Zd�8�5r2�m�I�m�ײE��{s;�g��n�8��7����C�[v��5s�C6'c�u�A�QW$5�ƹ����-�zI��Tk�v�b��z�p�>=��%g��9-�a�0	����Ͷ�!?5��YX�M��S}�䓗�}�e��Ǡ�u��9�B ���\�
@���:b{g#��Mv�ԸG3Gё>���&{\(�<Zmft�j���n��Ηco�)>k���$�6�\n����JΩ]u�y>��+9{�%�<}J za'��[���d�մ��pѫf��1�tu;��.ֹr�|��s*b�v�]�%΁X;.�>����<yϝ�+�V��ZE��J ��P�<ߣ�{�^���l����˺�%2�Ko���WT\:�q��"zf���$�{�
�Ye�0�6kea�{�O��KC"��1ޚO�V%QN.���a>�a��*�p�H"1� �1�v˚��؞M�٫C8˱iEzM)LP	�*��"�׊�^�t�z�o4c�+��Q4
�W��mt���d�	�T�ʬ�v�Y�I���m�^��1��#4����ܜ�!U5h���T�.���!�.�w?OE'6$�
60�Zaw�S|��-\��T9�v����ȃ�W�&*xwf��\>2���t�qz�6]d��i�+q[�Qa3�Z䷻�j"&���cs���ux���-5��L@����!ksL	�	��t��QpT�H��|����4�]��˃͑��(%�T"�X�bh%�`��X��00����=&N�IHVkm������wW0-@bJ���5�c�;N�5-�yŗ�^��¯)�#�%יZ ���w檳�������C��.� �Qa\bK�,���iD[�����>
���$�]��@N�VN�S)�:��w\��d�\p�饕���Z���s�-�ʈW��X9{��fs]�H\����/�q�������N�>�g�-��(fy�ީ+m��RZ�����j�=#��J�P�wN�mZ�Տ7�ֳU��(�bgu�]=��x� ��+@�"�!H a�x
K��n�������O:��y�������#��}6CՍ2	\� �ˤkV���a����&
lDKlp�*3���&x+���T��Q�s�̈́��U�@��	e�ٵ-7qC�{(��Z����댷-C�.W�E3����~Bw+�ņv�����#�H��V:%�A�lٱ��U��C*.���͋a޹��:�΃���`�,����c�EM�:��x��ƾp��:�jY5Jl�R*X�R{��B��i�b�~�vk�����
r���'s�����Vk�4��<�Є�Vħ%B`��EP�Ȼ}l����� �d��V-��l��;�	y�:A�����/�{LBN��K"�=�ģ)�%<n�7[5}9̽����$2�W�q�BB�l��`��c@a%Pi;�<�L4r�E�^gh޻���m���A3���Υ\�G�D�5�(��.���d&40�
8e;�8rꢝKTN��׫���~UN����mkJ���&��{90ڠ��B�Պ|z�?0��r�b�/6�h���y/`�i��SX=���m���"�*[�j�Aכ�@2��)a^��n_�N��4!�L��p#�yiB��.�N��:Q��m`��5��w���$����f�	[�g�a�o��_>��!�]�ux�Q�!r5Zh�A������C�z�U���}_y0�{��x3�֌m,إ���hk��i��T��n\���BaF^�Gs��]Ct�4/Mx�}��p[�WȽ�����F#��,b�)��94�ܚMl�Еc
�ҵ�%�^��4��f���|M���;4�0�����v`�
����O�!�q�z)�T��~���>�z�3�^;r�ld�&(;V�M!��ŝc;�B#�3�w�����'�o�$��d��`�zHrC���۳���3�����1-ָ}�oQ��	�iD�	a��Se�ӱ��gsg)s'f�Α������މ��g o��т��1*GYPl�1 pk�(�w��ǲ�d�*0�5e]Ns�=��[Wn�4��0�
�W��}{6���6�Ӫaq`���q�TNr3=*�`?�gvN���Jq�MO�^�"�⩛��2#�'�$v��ŧ�z��]"��u����2�d����%��>뽿�����j+�7����d�,SI�WN��,:s_��wG~�ek/�dv9#����`eT���K���y��E�\�:!�(�E�Q,�=���ռ:���?J�v���Y+�
n]���3�嘜�
�L��0��2��eh�����r�v���jR��=W ~����('C~�2�{ �V��}�K�`�WmT`Gs�U6��,����+�F�䡡�+^ޝ�XJDc��������H�F�hJS\tw�s��g���(�f�"���}F�R9�x�7%tB�H#�	})�z#���z���&(��}����z� Q��Ϸ��9�Ǟ�kg�۞�����,�g��Ԙ���̂��+�p�R�];�r�n�F����5 LYz���=���C�	��r^9���$���s�ǳ5hb��j/x��I�M���-?,e �����F%� y�л#�xz����e-�+pO2��AxFķs�깦�ʹ��E��c��@'�q��ݪn�`å���mﻕ��Cld��R��ʯOW�s����ɚj�zR~k��y�+�_�rjNe��7�?� ptg���ȷvc#�`����C��/^�����4-X�.)06�%��Nq���~�"����_�-�d_p?�#b]��9g�4Bb��}l/S����q�����i��l�[���e^g��S��J�H=~J(�y9�g��T��a9z$)\ώ�l����OL�U�={��1�����Y�'�IG{��|��yqt����~3���3͊�>�P.��Z-������n�2�����t�+-U����RoY�q���m�N�x#�!�9L��t\)��t"�:��vƤ��;S����%�3�؄�p3��sF������������Z1'\էk���ō#s�������(�H��% 4�JDSD��ըn��l��M�L�sӍ��z=ז��kL�v�8�5{��i�Z��<����1?ncM��z��;n���3�{�b��}]��l$U�A�W��!���r�Dq�].�O�5�9Ǹr�F�%����E�P*&�~ʊƥ�B~ka�خx4FYzxNd(x�$�0Eb҇�uk=(���_�Ѵ}dD`9�aN��T�ՑрFB�"Z�,��L��4���D5[��\�֪�֮�j�˜jꋇV�ϒ ���f�𓲭lK�;i��]p�k:ݓC13���j��=��Nl�Z�TS����"������<:�@���ٸu�����2�b�ñ�J�,���LW4	/��4����O&�Ý����g'�����d��9�C���= ������*���jRy�Sl���AmE�v�g'�M�Y�f�u��VJ�vjg�^�m!�a�n�=���t-W*��\���W(�ڮ�����6j��g�*]�]ߴ�ތ���i�� Aa�7;��_==ήMгa̜q��<�\ɾ��W�=���07����R�-��DRJ��w�h���qs�A�f�廫5��6�Ů�}��S�,��pq����D>�ڻd�+��i��wTk�"R��n��4��ґ�Q h�'o.�/0G������ �SyM�-s�}u��)�
��J=vo����[��'�����3��*���>�q�d�p����Ѕ��y�>��q�7z����X����{����Cdm��I�V���7?:���m�g�� �\��j���>R�#�jb�ֻt��Ǥ'eۍ v�j~O�X���ں��bԺ'�^�9�dK�֔�C�v�75��6d�`�?Dp��R�=r��i�͓#���Wy�#Cބ�ޑ�=���&�1䈁�}s�k�/�O��g��+CBg�	�B|ab6��v�Ȳt�$9Ni�g�Q��ˬM�]�z�:�ƪO�f:���Bx�&縩4�Cxv���PV���?v��g�~U����x���2qn�ݒ�5曌�M������az��"�Ws^6&���.�{�d��P��8���;]b�W�]
7��5\�ʤ}X�
�K��=�$�`�p�ݒ��!���5��U�LZ�a	���&T*�d��Ӻ�1��}F��%��$Q�3B��9�~p"x�F��|���Ly�� �LP�yP����4{=>�_����������o�������a���k:�Cힱ[m#�@�tNc�0��{1�;%�铠���\co;Q"u��AL�;0���mBj�ysOJ�K" �#� vC/g��v��r����:+
H婒S��ԡ��%�[�8�����y� GL��q��̉j�t���f����e��gRd=�Etm������`�s&�!epت�9�y��0*�*F�q�FjOf�Kv��f#��r�ܐܮ�������[��z�|���r%w�3yuʗ*W�`�nB�2��<�8�CG��)�f��49��[[�zy��G<b}2	�k���"�%δ��-��[�M�S9S^k�T�dQ���JRz]�^e�M���!�mʁomq9pōS��n��ڭ���o�^���4Ã��B�Y� ��$�Q�"��"2r���4ň�,��d�4�֔�B{&eM��6q��;�\B����_$��OV�a���a���r�s�޶pѾM��V�T���9cnI���ͤ�(�R;Y�"䢑1H���Μ�ћMPu7�5ۥSL���X�îv5UWy܍��~7Г�M�|pݷB���f�V�!��J�� -�t:k�+�@��u�;Ļ�%�b�X�����n�	�݅��Wَ�����j�\�Ģ.��J�qՓ�[ٓ����a�lx��q=��&��6.��UnvMAr�/C�܋T��O��r�r��{L�L�P+���j���j��}jm]J���,b+�,1�dL�o-P��or�nX���o�T=j�1N�ʺz���ݐX��4%�։��nͬ-�J��A�uG�ɻ�o����u;7V�$E�7+xkS��و%�����Y�h*:�S�DV�,�&)�����Q7�}���ڳ�ÁkII*���ԷwQЩ���zd��g�ίDMV.&�1W�]vw���k����uiδ�^�YM_>��W@p5S6�r�P]@G���6�Q�y1��lgm�N�uꕙ����]���K�]\&�̎�qeXԴØM��nC�=8,U-늻dI�DV���ģD�4���!�G��}0��q��:�g����FV�c��O8�����E�ς�ACܣZ�
�˻%.���_Ĥ��Vv�v�� �
2�Mƴ=ވh�P��I�}�d���
��O�!�8�����K׋I�6�`|N�T�EW
���u'\֩�fuu��"��%�y�Z�o�>oN�����7�Z�ɟ�1��x��4X�4k
egk�ܒ��5Ǯ{�C	 �T�iSU'm0i\��;z��v]L���.��G���h��ڣ��8���է��36�	�^wn�;���wd=q�麓���(�qvhY̧��8r�QEK73.���$u�.t:�v��uP�{�9�M�C��:��"�ַ{�Nvo@U�I��|H �3��
�����������h��� ���fZ����2����#3"����f$�j���frq�"���*b�!��
*&�b*�*��h�ɢ`�j�h�d�̢���"�"�����f��2���UIISI�(�3(�b�
�0Ȩ�j��"J������*"h����,"�����"�&"�
b"b����	
�	$�������0(�(�)�32(�����ʆJ�2(��(�i"�)�0Ċ��������(�L��������$�j,�&��ť������������&�(�&��bUDMfc�QR4USQD�0PAQPUY�HTU^?vz��4YI�� ���]|�%�Φ�R���V�}��/�Z�5S���Y��1�V�Z�v2UR9G�p�vf�3gi��7

��ɸ�o��_&����J�eO�L~@}�G��Gc寵Ӧ�+������G�|w�$8��rC�/ ��;/�z}�e'X^%�u���/5�
���F�"��5�0Nb����O�_ZAvl���s�Tư���w�yN�R./cP����t'��]oɔS*�ިn�`Ӗ�p���PP͍"8Bn�=!1���Qm�n��|��{�����
KiKը�����4�L?5�\<{����ZDp�n}�P�٣{�3����\�$Ͱ-�܊�*�=��s$R��k�<h����
' n?.�X[OW%�cuS�>N��ؖ&:SS%	V0�]+^�%8�_)�T[o�\�m�`�Ci�ڧ̉�s;Suwk]o`�4
p��E��!�9i�d;n=^��+�I�����~%W��ʙ,�6]��Ǌc���J�7�}L��a��v3�|����y�����z�GX����(�X/�BӢg�sE㌨��+�KK��ٝ��ZW�ED�Tz(m�c�Q5���_�+���{�H��65���ELZt��6���a��d�����=N�_E���P���9hd-�l��7�vC69i��x�@�1y��G�wg�~Lde{{������	rKc��v��#���]KD�W�3�w�X�r�w���ôm�jmY����ye^ޖ�\�M��&XF�:Y���� ��#(�Garۘ�Y�1�w2lΔ�Mô75�>���y�{��\l�I�?���s�r�͛�Y�}�%�rЌ�p�{6��)�����sK%�s�K�������vtJ,�!S퉩�����j�S7Y�A�ȶ���z͜O^�o\���dL��|a����l:Ën�����38�.��W���Jm�2b)���]:á��A�)���]�}�,��x/m��`xav"!��v�#!O6��A8�Q,�ƶ1N�����g2����Y���;��pKYqCM��nG�r9O�C�+�u��F��Iz����e�3{ͭ{��q���սZ�=s��%:�R)�$i5��ܞfǨu��]�ڽ	K6Н���L˹�4���!�\'o�g]ĕJ�|1��n�G�n&,�>G�|�B=F廌���bz�z�:q���=(2��X֟4�v�㐙���-:�l����uf�p�D限�*�MU�-�ـ�L.H��@��ؖ\�U�7X�U�v0�/-H�0�?s��q���<6�`��+���B��o�������6��y�vOƄ�
�W�&="��3mZvR~lD���~�c>R$�U@.�b�،{����tq���x�37�B,��� eZ�m�-|�`j�3�ʏ0��d�df�V�|��N�e[����ζ�^�3���ficr�w1��&oI��d�kv���bGՓ����pvK�������|�nK�G�{;y���ΪY�(�vn�l0g�!������z���C8д��t�qi��	���p�õCIt��ն�+������Nd�qO����֜򯦵�j�6�.&���[�6�nJsgu�^Nf�P����q����yXH>L����sCH���y�sMC��{��ʭ{^���M��χ:D���C��㾎����(��@lX�>��W��F���\Є������GE�S��輳L�^�'����A�r2�6�֝#E�feTeN��~���,��D����L��8f��5s���ZԶ,�[��!���q���[WJf�X�B�u�6˽cdcG��G��a���q�[5�f�{�2���9	���8��Dr���T�s��dt�.��ƼI�g�c��eEÚ�"�9�
|C�����j��茙���z�j.h���F�����< �^��):���%2XKo���P��9�dk<�-��,ױ��k�+���j�O]�t�#��D�Ԧ-C�$�D�6R�j��"�w�"�{�������IuST����.~�nT���_T^��ݣ�+#Ob9x�*���C0�R��sב{�q徯_�D����wo�����y�I���6�V$�V"5:�!��&\���M�sR����wJ�gi�����B����g1����aԟTŤu�n�����m��rÏ�}�r��/~��{e؆�;.�4Ҥ�x	��%�ޑ�GM�s���f�9��͘��3 ��!�O��= ��0��T,�+�������d]c���3���]����bf��\W(���?j�5�{�	Χ��=t+�0�aT�\��8��w5l&-�;J�9�n��z��ΟGW��x�b4Y���&�	��	�ubMг5v���Hd_0�Kt�^�2�T������d��k		]��+A=@���Zz��y�>�DC`ݓ�r��������Ԭq���{A/mbTs	hN�5~΀���f����F���b��=s&I�|`̭���_(N˷ol��0�@��t�>�0�;^&����/>�b9=�꙲)��{�*��I�A��k�DB`���������t��E�1%ځ2�q��2ƷC�u�,67,���o7���kj��伻�Bg~2�.|\��fɁ����2	l��x�F��U��m�_w�	��I���W�T�Q��Ay	�o�4���V�Ň�"���?VD�Z��B]��\C][�ڣ=F\*�[W�����U8���!�� �S�Įhv(yg)K�-x���2˕�����7|moa�Wun%fas:)C�5X_P���l}-`p��m9�+(�ܬVd�q����s�;�K������M��}�='8�tU���_-E��%r��ךE�[�������� ���8�sE͙c�����B˓��Ͷ���C��WUKc�-{.���Q�����O��Sxg��&փ�E�!�O����]�Ұ{N���YaK�1�Iv��s�	�G)	�,T)=��g�1��L�5,�&_����y���^0y��G�q�����9�t!)�g���SΊ�H!î��O q᪫23F��r�-v&gԭ&��^�WB&8yYY��,��~?x�|
�~.�H��Gf\��m\�;�5,�I�>�s���O���3d�&���c��*̧y�P���5>��[��h�Ǒ�.�,���-�sjQ�NZ��kÇ��3cH����&1<��Th�q9�,1&�s](v�wAb���Z�O�iAb�?7'��ݰ|��2mj������z��g4�e���@Nҧf��f������C�}�f�*�K sO�Ӈ��o3�,�4����ܖ�TB�q������Ò�f�z稵��%8×@@��˪~eU�6k;qY�O8M6C��ےwlgO�x��q��=�fg�j�����C��U�k�cH�J���3((�	��ڷut�X��ӽ�R��M^ώ䆟gG}ѐ5_>8� �H��FU�m����d�N�߻�Սь�b��{�'E>�oj���T�~��
໌�cD�ьf�6n:�=I������=�ͻvU8뻵st��\*m5ڐa�������ȇ�õ��!����8���E�_�Zӽ�6F6��w*���^���m1^��)�W�a��P�}`/���_�q<=�{����MJr�{d��A���!�rC�$@"G�i/���툨~��,����2>*R�:f��eh~��-��z-=�ז��Od�EdPA�2a�U5O��\�͇\�}������k�֮���}a�B�G4�FS��O��E��j�S7�J���PH�͋Nޖ��]u]żu��qekr�Uȧx���,>���j��[/>�"b�(2j��4�C&|)b
k�0����U�B�YZj�'Èv?$=��d@d���'d�Lp�v9����`��S���]:��L�J4��Dv>57�E�r<���|b����������10g=�7��+8��tD�%��'Y�E2�Q���nO5 ���b�ki���_��^��e�5~�kh#���mXK��`N� Z�|N�gf��?v�A)=}=t����9g�7�!�>�f���������c`���j�p�D6j�|a�rӠ�]J*��]X+K���]��nXǝL����բpmen��᪨��zk�ݒw��&���C�Q2��R�č4�'�b)9C�Iኸ�>�-K�?-��dR�,LԹɟ�F��� ��	�tYc:m����e1�6����e ����uk��w^�_ �C�Q�tE�A���
H�C�H��e�c���o��<���a�^(Z��a��xWz6�9��v���|��ת%ݡF3��r!P`伈vNU	��nL�cPM[]����*�@�'o8�Z��z���?��ڨNV�H��k �0��qwf�E�OC���B�R�6:���p{����)�k-{+�շ�Q\�����9���x���֜���]c:_�.1{�G7S�3���I86��0��Ŏ���uƇ�^>4&Sاu�i\U鋮��i�Lj|��ܹ�B^P֚��>j{��s�^T�B��L�v)����>ŷ\��O	(���"cK���m�;����f��'����r2��t�R�f�e�xw!I������"�@1�L��,�w��C��3b���a ��[|�t\�����?uݶ'��v;c��S5�q߿[��S-C��-���9]l����3�䤞��.)�ewk��j�$Y�?kG4�@�L�M��Ǭ/.G'%ђ+,X5j��6����Γ���`I���a�i̥��웵�(�5:��:���	?�ΧVgOO#:
��5����z���4J<��q�#0;�TU�Le���2�{�zyn�E��D�6��.��Ɗ5�����T[^�	�?![��<�4�;�̜Nܢ��*�m��VŪ.4�Q6����X��B��U��8�/P�=q���-�M���)�
��7|I���Ǵ͈K�.���f"E��-C�$�b%9�
>V2.U��6q�c�B�<�W&�����٧W7�� ������A��v!�_v���&X�LU�y^�\h������Ҕ�M�o��e�<	vT	 B
|ӍB� �}�YPU;M���o��"��Iՙ��6�f��m���!��-#k˧�l�����=� p����z��N`ԉ:0�aW�^r�n���Lі�+C��e�*;�P*KGjOLBƋ0!�}�!Ѿ5:�Oc�zb=���D���:[#m�$�k��˯դO��-49ZH ��� i㗧�6���f��7Eh�m(NHLk�UV�X�?JװT��%G0�Нj��9�/����7�����\_��D��{[Gp�p#t����x�j��*�k����~֨��Ҷ��|����B4X����W���x1)�q����|��T�E5�y���΄9�MioWlj
�t�=�ӊ;͗I2�j�U��o��E��ho,vܮ`��F��õ�s^f^��m"�:�N˲��XsaJA!?Mc�v��j[��@��@�vl�zz����u�:\�
�.��t�������'G����ܢ¸ėba���j轝md���*����w��P��q��\d���L�	��3���s��{z����)�TN<����v�!^�@�[����\z]��XD��z���c�L�
�D�����5�a\�S�!�gQ���1�@Y����f/I\�(r5曌�MC�.W�)�0Aa'[&���4s&I�t��]�P��MG5vL�[.0�aT]
6�psU�w*��U�>�5!��pe����֦�`��G;,�n\'j[�����d�Ȓ�ʻj��ǧ5�[�֥ռ�����R*:˃+�D�BP�}^!��|�ڽЄ�\]�JtB�L#=���tz=�mH����3�?�V`t4�|�x�2\�.�=��P��Z��>�����t�����ۛ�y~խ���x�44�6��{������3C6;����40����.Y�F�b�l���B��:QҪY=����f�ėV#8�Xc:��/��/�1����&}�Н"��(�"�Z:��]��Z��U�mƅ�}4MhVt��T��jeFzr�S�ZK��6�nil��-�ī����Mv�ۺwz+�r�QwCTQr�ҩE�y���~ާ.�?Z�$W��fA̜+��x�����=���s��s5c�R'��qH�/e�?2O���t�~d�=��� /��W�e;�Fy�n���GSK(��N�7&m�j�r�߸�0�-D������Գ^(
��T�W]�K��˼�;�
�z`r�v�94�o��Z�_�*�9t�{*	{��q���Ċ����S���\�:Dr:ǐ�/0�c!�q�׽6�ħ��ټ���m6]�ej7�w���ӎ�=3ƽ�	�C��G���y��?�Q��<�q;_<�c.]�ꨙ�#k�]�x��r�O�� ��+�{D��V!�Ϻ%�XG�>
,�����8�s�������}����r��skCN� ��	�=N��_E���EC�dK:Z���p�k.mFpWf67�ps3�l��W=	�{Y�C�sqS4�d�@�C�yyp^M��TTr������mE�Z��ݻ97������1:9z%4���O�����5.J��� ��d������v��÷�������������v����3WV��1^ާ|OV�x7���ےM�Wq��atqLk�h㴬�ݘ�l!�;]�O���@�oS�]jY�%�����J�Le	�!r�[�+JވCVL4:�I6q�-Ʈ��[�]v[իA2R�l�a[��bm��O�8m!���]�-�x_F�5�p��;h&P��;��`���T��X����{��Yt��fI��1)P�%gI&����.+���Xƙ����{��;�/j��}]0��`
Y�IqH6�aiK��r���p��몜񷆤(��s�Qپ�󝌦k��핬��
A]�T�(;��V��[�b��5�;�j¶*����>u�]q��tܨ�Zä�(�JV�E7n�/�:�>C,^��OD��Ff��!��+x��l�ұ*��4{9m�%�H�!����U�Q��{]�[b��Z�38�ڧG�D7�n�	<Bi�٦0���S�:�ʜM�g�+�i١�X����y�p�����8+�0j:���ioz��,_G���ێ�;(�v[$�7�*\U��t�?t�F�y:���ȍ����-�,������%�;/�խ�ȘZ%M�<��l���N� ��)��5rׯ3M&	*S�`���+�8��	l]j�vz�݄�C���MmfѪ�1�f�3�
�1�R[��] ,<@���D��݃�{�8�&���Y���x��v.A�V��B﫶[7���j��e)�bМa]�	Jbfs�f�վVr�ͧ# i׏mɨ�H+2󥫷�l�ʀ5x�8+SZ����t�e�}����<�?<G?aE�,~> �U��פ��-޻�xc��t�
��`�e��ݮO�gǛ����q��j���B��\HM&�Ǧ�8���x.�ݧ��<�����v��g�6Q�ʧ%�J'n��*��V���WB�]%7���@oMCgJ�3uY�r��9Qq�xGE�2��12jV���W@�Sv�#�"��+��\Z�F��z�tv;}�M�Z����c�˵kU�#�b9ue�A���L8*����p�P� p�h0��aZ�|+157���U�u�F�)�
Q�,�+�f�Z&�V١Qu��}��jfQ[�^��7���Β;�Q��Λɮ��a�e��eB/K%�F����w��H��ۨsr��4������{�l0Гh�6s)3|+��,6�<�7�+�μ�����{�UFP��a���Z;$5��Z�[ZI�v��5�\82�tf��fS��	�pu���6��k�7��-���d%H���/h�2HnVM����S,��l(�t����[%��^���&.�VX3�ΐ��l��T�Xq���0���<��@P4���a2�TD�Wu������]����x��+����tSYu�
�T��\6@�,3b���Rε��'\��WDb���KP0P��lm�nU�:N�I�`�)�j�ogEp�� �;��fk�:�wř�r�RPUQT�%T�1DQGAT�!U!IEEEdUSDUTUD�Q�M%DYaLI@��ITT�fD��d�DS�aE��(U9cIP��SSAMPT��CA4�D�QLM(U,DEA0��Q	EE%P�AJPD�%TPT��@R�JQ�"(�R��&I���Z��ii
�)�� �������hi�ZJ&�����i)$�h(h��(���(�*������B�$)*������")����(i
B�(����������z|�=L�K7� W^�y����ݮ�����I�V��j����C#�I�9�N�}�m<yF)�@ݞ5|�<�~��߁�5�����)�.=<(*�`��Ezw���~�(2f�6�@�j��`��mB�MS����}�l��+��J��9aL������J�g����B84h����7���2����
SL�ҍ&��Gc�W��<��������|b	+�wo9�ڛ�`��B������5���g��Q�'�D�:�K	Mm`F��P��\:��<��j��MK]a��cx�/�M�hSR�,0��2���I9w���=fu�� ���#ϰ��k�_>E������"6pN�H�d[c`�7pΛjOc
�i��mO\�����A3�j-#���0�u]�v�nN?_ud�`;̽y��l�1�0�s�6%�=���n�����a�^(Z��a�U�(�;�oq�k�����߮/ܼ����,xQ���B�P4����
�P`K&i�\^N�1!8���;��n�#O��V�a\�T�exl[�;5�|<y"u~����k�ϥt!s��Q�r:�{7r��D��S���O�l�W5������Cs9��G�*��������X5)ʦ��q�v�z(�%{R������olH
�I�y�N���j��В��dRMb;kɿdW��tLʔEL�<x�g}9P�̪�R�
��a1]��Kю+)�v�mNwW��Ɵv�bkheH��Zd[��2�����d�'�+����O��5�*�ua��N�a^��;hb���r�^ø���_rmLzK�ն:�[��;H��xsnP������Ar�gA;�r>菌��=���i�z��\�FT�k��Y��p�yꗲD����}��ä�:-�����/,�4��-���T� �3$�:���]�i��۷�;slW�3eu�D��#�p6�;�M/�[�Y���[Dt�����泖GO(,��Hj$γ�l�*�Ξ|��6�7D����M�È�vQ�\x^T����̱A�� ���-�5�k�Yq_:V��Ј p�.@���<�O�9��YrĦ���e�%�W� ��D��&�Rt�H�URaMKnq�^��=�Х}�ZݼS��v��ܱGf�,-o/T)f���iv�^�7	�S��L�و���R�<\R6q�L���5k(�Ι�r��ݠb��W%�!�v$l�C*��bo��N�M�L����בE�&��rb/k(�ќ���Ϝ���m;6S���Ag�]��N���Az��ʗj3	<ϟ�'KĎ\�ǣ��6K��ڊ6��f�W#���*ޙ�w�V�Y:s��L���K�w�;�I{i��A�9R:��tMԔU|\u���{i����a��[5�m���e|F4�v'�;0��+S�J:4�.���N�	WX��F���w�h����c[j�	��'���/W�����W*K��
���@�=ʽ=�ܛ�GD�5]/s+���4]�i,
*u<5W(��JKGj&wvjq�Q�a��c��/s�V���UY[����7l�*�(zz�Ye�V�TXP��I�i��t��h'�W�O<�v]ܵ�������4�aSS(�	���C9P�n�c���+\�%錨��'Z��;��9@�X+��;���Zw7n+{�`��̐PZDI�N˲��Ú���~�+�ô� MN���&u�I��1S������H�Cy��ϲ�K�8y�l��Yۗ&;�X͓?{r�
�]��$������D�ݝ��4�Ĕy�Q��\d���L�	����>0�F��#���N��OF�p�
��o{q�;��l�)t��ג��H���p�z�ʏa� pW�k���~!��n�`�N�yo9d5F��G���G9U ��ךE�ۦ���u]�`�D)�R����]���\�����h�B0�kؚ�j�U-�]�B�0��T�)Ok�͋aP����gQp�t݌�F5gay��]�����8�o\�[�SB%q-��cH���S�� ���^nL[�Vwuw+]�f8���0LG,�2��Q�W��,�CRqa	v��"�d���2+�sݘ���x]��$MJ�:������*�3pM��:�Q����fG]@Y�.�0�����c���׾��4�q�'g�v����Ȕ�<�&K�Oʻh\U�*ffޱF��8mﵪ:���YQ4n.�$q�](w��\�[�B�_�ħ/�������������mw����*��t�=}Ǆ����1d����׻|k��'ȷ��i��:�V��}A<K$� �c^(�aO�\��a>�� �6G��)�箨 �;!�΄aĭ�~ҟwBs'�׭E'L9L"�7E1�-���Nh�$F58�8��Ӓid���ʯ^��?^�4ڄ�ʱ]
Xe;�㊺^��~n	Ab�?7�\<��$�v��x��^Nmk8g^�<�ib��NlI�`Z����Uz���s2�w?�؝�chj}�+���>�
�@G0Rã�k��;4ڣ��2��J��]+^ʂ^��2�w��km��m�ޘ�L�\��`�GH`�à<y��ͮ��d;n=z��m�*����N��\w[R�F\���׮S<�j��ņv2P�#G�+���N#�@������6_��.Y����('�2[Mc�|���&���DV18ռ�T�6eL[��
�w��5;�b\�̺6��ϲ.ٽȉ5+:o]�׉W��}r�$Ⱥ��\,�ؠ�e��wf�ĸ=�xӽ#	U�YY6�%Ϲ��V��t[�h�*'��+�K���Ӻ��Ǥ��D�/>8X��;^�� 円���d-H&[��0h쭙Yo��ܽƃ�ͬa i�C׉�ǩ<�;jT�V8W�6�D��Ξ��b-hE���tv�<�'����ޡ͛���5�a�����a�4=��}�tS���݊��Ք�ʞY�`��҇Bg��s�}��Ơ�*f㰃"�q�j���|#�<ާ�j祈�q������Y^��"�A�.,Gx���Ӣ����N��q�Ō<a�Џk��RYP�k^�>[t��f��81|O��+2�K�	�4P]�����xw"_d]��T�ڋk���Y���e�j�B�\Pn�d�A��>1����-w�٭-H��f�`P<$6����'�b%9�R�ޒ4���nO5y�.P��+|��5])��f��;	�;a�6�����T�A�f}fS��4�'.��Q����5x����sX4�P\ut����]y�Ϭ!�Bmzvx7Vt�R|*�[����Qi�`�� �?�&�e\p��*ِ�E�pxfʅ��yZ����ej���M\�ohӂ��7 ��(����/�\���r"��G�j�u�I�ل���r�do7"�>c,�=��w�d�dꔉm,���B�k�Iܸ/84llY���`Q��>Х�5mL휻���_�~^�u���]�����!����V:�Q�ʹ���/E�˻4J��v^ɊQ���n��xƿk�*�ćA�/�x[A~�@B�S��ީ�+���!��|����;9��U=y���Jx�5�X�y�s�6����i��4<��]�>h�E�4M<����F�U�'�@�n'�9�"��u1���r��i��m�}����#=\�*�╙^���Ŝ:U���_����v��u�;ϵ�hGP�I8)�K󞽨��߄�=g���UM���C3ݗ��wڃ@���Ʊ��;#O�6�}�9�+����9i�yO�k�D�o���C��2�t��C��h�q�10����m�9�>��4�44�����αՐ�4���Ζ��q"b1�r/Ɔ����I,x���@NY�=�5s���bd��̻�^ٷ��Z�����i�����!�gY�fͲ��.�D�A���E�P.��2em%y���w:���S��[�A���&5�k=�|jʋ�4./����^�Kʿ����m��ny�g~�,Խ�^#~V�����["~Ү�	h�j��`��,-#4�$���+�����:��q�]�y�ۦR�dyՃ��V��+����6��s"糪Z�}b�o}�F0"�CV��.Fw3uH��c:{�n�Ѹ_(����	L>"�Q��wNGE|��5�p��l:yN�L�0�^[s�^ꋇEu/-\�ΔMl��=�W3�r�F�]K��`(^�7	Ҙ��L�߁���"���)Ŧ���e�ǔo���n���O\�������8�.�A���9.�4�YR�#Ozզ��&)��z�����ltw�����6^���H܁!�=B~����o��N����F̽U-�&y�˩�.�b�`>c����s���� ���ڣ^@va�<��vA^�	���_�~~6�����J疡j��JKGj&wvm@pB���C�ȹּ�sѹ]�����2�N�'W&�Y�9��/��ƷJ�Z�B{������\0fJk�%���ۭ0-iA��[8.X���͹�E.u+u��+^�PK�B~a��	�9�Ltq��U2��=w6�m[�p������4 �������m;-���)P6����Ì;N��5o��5Z譓g(��M��@�z	�A�H�V��	`] R�;b\��={���w(�>oI�*�a��W�������z��u�Sm��c�貉�wX��l�hy�|���%��j���~l�����}�~��f��x��Z"�貐H79mt�	}���H��YxvP���ǅ�v1��	�:76+=�,� zF�B�ᙏ4��=�~,+�[�����d�;s�Go�ӷ�fX�
����-�8�r�0�+��%	��3����.;�\v�o�㧂����N�z�7C� ����=�0<¸������ՈD��ߍq��ܜ�$_����'��;���N$9�kM�r-W�G=r�r5曍�M�鋗ZS>^9;5:���O�r��Oe���A�R�I�u���;}#�����,�m*<����C�v�w�r!YN��{����>�7��`��!�bN�2Q�ͣ��M��&Eb�I�iHd�9&����=O�Wr���i�b�Oma8�*`$&��CH�S�΄&S\#Za��]�_r��B�Prx[m�yl����+��a�W�K�����OC��T�]�)�>�-��t^.�9]����e)�Hpx�%L9�+��w�Z��<�Ŀ���D��R�_*�59Ygo�hb�$еI�E�Rt��*�]`�LV��q~��>w����.e=.����gu�`�������4�8��j�wqOK���',H��a�Zq.|����#�p�u��3X t��f�vXxK:e��h��մ;|w���Q���Lȱs��9��F�|��b^�����cA���p�v�)߶�{wtK��QG.M	�
���;1�]mJ�uSG:��ʣ%,9,*�b#&J�-��Q�t�踱v;L5U՚#���J�#��M�P�kuN�W&m�j�r��*����̚T;�.q˧��ɴu��^ �f����͸p�����u��f�U�Qkep�c
�J�^�]���=����M\dG]��r���:����]@A\9��.�D��o�X-�k�޿�.���u�?�H�}��8�GS킧ӏC��5�,ƌXg>��$�<�z�(�՞Y��ԨmZ�U�Nf��mg����!�ȴޞ/�x���Š�1^�tE1j��dtK� 兑����t�6�ڶ�7zS�ұ�v3_�4��0��0Hz$@"x�;I}��lEC�l�����Gq\n#7;Yܡ��C/hQ��lS��x�s�z���C6�3M{�K����dÇ���5���E=�LW:<;�/��������(~��	 �i���11���{3�K��n��aO���]����6��֊�듉g�MO���5ez�E�G�~��`��5��d�0K�������<B�i}ۮ*�,��RԼ�x2e�%:��`OE���o���ёÐ����U�{����3�
�v��Q}�g=�ʙ��F#���4�ʀ�k�ct��s�������ma��d�l���D��yޒ��W��]�����g9���񨃍P�f±M�s� wІ��p�X��躳�]��)���RS��nwY�x3+��:Gf�6�u�#�l�&��N(r�MGx���*�U�E�Kl��7��7BA������Y75Ze��/w�X�ݛ�&�|$7�K߬t�'I�lD�7�E1��&����O�p��=K�ouʓ�ؚ������7P����v
E�N�F�T��yNR�t�4*����\I�n�2=�y������pЂ�(Bm����Y�mE�aR�6�=�%�[-c�q�|}{��"D���y�Cx���#4�@=�|�-��0Q�0�s���eC�n)�]�������Z�/s�n���89�F^ݐX��U��{O���%݋�;5�h`�Ͼ�0����
�WUN��7��T��E�^�n�!lP�궻JR~k�d�ͫ�*�f�zwf���`�C�?�a���r(յy�L�����.��:sC
�i<&��k-{����/<�_p?�u�Ndy�_awm�8�]��4������~G��XJ�0����I���i�-�����1�t�Ŝ)��2�Ѯ����
�@�vu�#�<����X�6���z���Α:8�j=o��z��ӷǧ���������������[��4!���D�l���i��!���;�����v���q'����F���.ݾ����k%@:L�ۡέ�3�YOP�����"�֗H��nN�z4ډi%�����Y���W#�M,� s ����+]�}HEyr
YU���;x�,��/�9��"�8����4��u�d��|���܆���m��Gs�r)5��0JΣ]��'@j\�g���M`�0U��nQ!���of�[֝�N�8|G l��|�3�t��Ya��z���{�f�qr>ު:5�G:���I��(�hB/Ce�*p+@ՎN��eK��yd��r�)"���S�УYۏq�&�����'{���Fnj/�z��5C���������a�{�Hr�JIx�ڷ�ضJ�bR7	�OtZ�h�2�Ӡ���cY�w��_c�X��'(;,�&��S�n}���Y�X���Oo�e�Sř/5r.�5� ���^����9����
���z��ħQt%'1��7B�Ջn[w���5g�$w����˦��M�{/���[&���U�]����Z:o`�v�f"6��Zʦ��k����JU�
�ø���ǖ[�D�'n�)�4���ۧeQ�Z��#���J���wy�(2�_֣�9���x����Ѹ y����]bՎ͛���9Y�e2N"e�|r��:n�F�����R43��#^ͻ���e5���˹�@���w���`j��0���AX�՝� ]+�O.+���N��@K���]\�&�Z�������5���>�<�,>�N��Ū�f.c����>���l�����zP�O<�96;�r�<����{��Z%p��B^V�]�J�e\�v[��v#�=��2`��Bo֟F	��9#w��	�������k��q|�v���P���Rv�_
�ʵ�\ywyOz�We���I��γ3(�&�.�c\�J慅hIE�30�/7F��a�`��Q<\��ۘ2
Ѽ�2�m�4]/�kx��&h(k �2��Y�O��X�.�򢍜��]z�d�,��+��֐���h M �֌7a��nn楖��wۗK������7�J,�dn�F���|qW��](J�K3&�Yq'�>�9��%�F�P�6�	Y�ۡcy*ekűKX�4ޜɷЩg5�¹�q�YYp-�!�������:�l��D�J�a$���v9	��l
�1���6��y�/�M�ޡE� ��Jwb�7z�Pl�F��ի��;:�=���{-�{�eV=������/��M�L������%�:L��8"�ۓPJ�=�9��l)��'����+f
�Ҥ�8���Tλ��p+�q��V�t/�v�� �7]�[�#�{&�d�PIk"����I���7�BV�7{�5,�;0&�| �]�j�ީ�v��橛�ݒ�,}A����Pd�`_:|h��
�����8�sh��FAV�%&���ZQ�{���+��:˾��9�*
X����)i"B����
��#Օ4SI@�@D��T�PD)�I@A��5JUUCIKEQATіMPLSD��,�LAICJ2MSI@@Q@SH�4�P��B4)CE P�%--	MT�IATUPR�@RRPPR��QBQLM%.A����4%4J�EVI�TP4� P�UKJDKE ��AQ���4-%UR��5E P�4)BR�	AHr�>��&J��n��<^
?P�A
!��.Є�ƫ*�,�XԴ��`V�(q2�h��ɺ(���:�b[ٳ&W^"�w+��HtY�EB�%�>�&�ͣ�����j^NA9���~_w��48͕�"I_x��"a'W=8�nw��/,�4К���pӉ�[��n�;j%�8�1&�����aQ^`d�%?���� mZ������W43�ZۭF�|r�^�z;���{"W�7�-@���Fu���Ռ��3�-3�	ĜS�����,�w�ٹkg����S���ڽ��At����N��1��k9~����=Ûp͛)�A�+HX�l\�C����8�jby�ON�j�d.z�,{�N&Ӭr�Z�K	e�v~�[�=n{�m��l�k-i_��O��f���f"�ވL�ߌD�6
T-1��ۺ�U����8�"�,,6q�ع��	F4�t���lʀ�b�öi�I��P��m۝k2�q���k�E��A}��!�-ᄁ�F4Ð��zA�	eyb��LDt�D�Ǟ-�}��P�U6n)(�[�Bx~�Pmt�U�\W(
��$!�V7!��M��x��o�<�[w:m��*MУ�S	�2��Z�E����5�v��LEcE� �����H����˝/R�<�՞��Qs���B{*���q��K�'���C��>�sc���cWc�-0Wb	�O�oҸ��q��W$��[�M�{���Bg\�&���71��|��V�{���y��I�^t���\jK�M���Ӹl�$�z���ӗ��[��h� s�=\ߤ�,`ۊ��QaV�z��)����ͭ�N��H�6C�ȼ׫�`ˤE����} ���ͺi�j�J�a?JװT�П�1��%3��\G w�6��Y�NB��$bؐ�||����,9��s�X8��k�7_=�p�є�3wf2��'i��U,Z�z'���g�D�Ǹ��w�~��vI�@�c2��}/=�wy���,`��N��Y�=q���Ϲ
+����<ăC�(�?~*�ua"d����C�ʚ����E��9�J��ȲkL�C�Jˡ���*��0!X�N���.�dE��:u1��
i2��ME��f�6�BA�_A�
�r3��덷MC�.Kk��IU@ֆp���.r����V��Ŭ�Dk�E����{��j�U-�^\�.w�2>[t(�Tyàܩ�����?v�s_|1��)���yg�>[|0L&v��b�.v����%6X�!2�W45�5!�r�Թ���u�4�w$RY�8��E=��[&C�L��W�i�y�^owA=J�f�E������=
��yˣ���L�خ��^'�Ձ;�ˬ�Bw���'�g&���9Xo%&C�(S7D��s�:Tǧw�+��ymԳ08�r��}�!�r]Km��`;{�|�[X���t�/�s�וL��ŏ��7n��Di����~x�O9��0蠻�B�We��W��R���� �����b����U�m�l��y�^ͪ�����xd]k<�/O�0����s��}h�a�7l\�뙚/rOb�xf�0�}�!�D�Ve;�<�	�*�]>�g+z���r��k���vYUO��d�N�N�GC2i�#���&:0�
8e;�㊺^��~d����0�ݼC�7C����%W
u������9���q��F�T��uf������	Te�Z��2�e,�`��[��{�t8��O�h�� ��[���R�w�N�;4جOQ�=�t�Vp�d5ك_d��݈Ъ��t�
{�T�ڮ�k����hp���:�x��]�yn{�뽙�;�#q�Zsw![��̭�u>߇)�b���q��'��`���%��&�EԚ�<����rjwG��`��-�����>��_��zHzZo�
��4@��>�d�_�jl�����?f�l���$D���'c5�g��s9��!��!�8ol�O��h�����M��Z+�n\�~��:k���/�óJ}�'"��QCS-ظKqT�@�����\<�D�6��2�����
��+s~���F8�==��<7��3]q4�	�ɴ9�fS��`��"��tn�Y!�f��ݱ��o?�gNs��㷷����q,��ZZB���|��ǳ�z�4��4�=�Xw��%׫�}�Z��+Z��a��P�׍��ZW�13-B������~8<��>��\[`��nt9�RŚ�Ŗ��@i�Wc���@�W��+�l�%� �p�C�����U�2��ҋJ��z�.��Q��^C	�ҡLV)��z1��Vv�Y^4,�WA�T��aαSզ��S�rC�n�d���'9D�.��d|��k�����l��S۹�.�r�ܼ�7�"���r�ħf4%�*�H"|/�����'�b%9��E1��&���͙���t j�e��]≣���US��Ǡ'f����hN�T˰R,�w��$�b)9X�Q��y�=�K7������Pw��|a��?�+a#��Bm��������K����/�1=Ɠ3P&�K�F��B�s�o=��)=j-#���0���,"�kL9�DlK.{깦��Q>vA�7kE�U�BNv�(��Ũ����M�㋁�ó���!��n�vO����c��ߩd�aՍ�Pf��Kz�+Z!q]�5ȵQ7v���"=d��y�d,zu�[�gA+����M��?
䣊���]|��З�dzt�;�Օ۝�p([�[*�挠��2�h;�ud"uf���X����2�K�:CR�]).�/s�taj�p�VK����X�t	m�Е[]锟��O*�W�+�f���H���+��l//��%���͟��f�|�a]���S�w���"�Q)����ǧ	��j��z�;v�On3��YE�N;/k��ށ� ��.�D�z��:}�2#�$��Nf�qg�	��n����d��=UZ[��<F��D���G3��[���d����t���~�Y�����r�I�f~O\���}���'���qt��`�~#4[� ���XӍ����Qjۖev�nn9�b����,҂�)ڀ*q�j�e�m����l�bK!`��mTw��]����YY1i������b���`��ˠŸ���Fu��f�V@�t���B����Z��GY����+w�cA��ׯ,�{��>ʊƮ�A?5� ���ƒ5��c��j.�z�Z��e<�N�m�1�NﳄG9
��N��Xb���tW�5�t���<�'�)UO����q�뚖�d�՞�~�QS^�o
@���y�l���ײ���ވL�و���*2*b#��k���H��u�M8���٧Eg���}B6����w��T��4fK�Qܮ嶍��-v�8�'�A]Bf�ɖ�n��9j��N��`���Jq�U��_U1x�����g���s�,���M�u7� �EH�cAײT��ڳfRǻZ�p��^:v��?v\dt�c�_��=E8��l�	��p�c����Nw,,^����b<}|eڡ$���vn�L׆��Sr�O2W�y\�2�W9�[�	܁!�!�O�:�A�n�v�']&�;��o[�w8C��i�i�Ry� S"�09�-�׺W*�%�r�+,�ڲ�g���c"%󯺧�_�^�Z�OE'W*�R���
���\��iIcH�C		��F2Y+[�H{|d�9�FnD�c�'�p]�b]	�srn��s']�*�]����w��bz ��? &��3ގ0e�YO�9b��
���dRAԭq��eK^�PK�\�B��>�L'���]y��[U�MCù����Y�����i�l;-��E�5aJ��̙����[

��}�K���b�5-�G�?6 ��"k����)e��.]�u��P�v���ȸF�u;;�����#[�Q/���ϫ�����adh�.�n)�olA��ݔ9Z��!s�{=�N����d��yt�I�ʇD����̀����i2F�DA�����dճ����u=q�2�+;Y���"۪�E�)j��q|.\�J�X�;Zb���f�K�C�˜x�\ЮÊƎ
�[i�`�/HO\�*<�anVķj&z��WD��{xkK,�'V5�۱�*�����X1�ۊi����%��n���G|.����љ'���Ƕ��֟^A!�_A�W!
�k�7n��7:ށ/����q�eu�kܡ_���Ņߐ��W��)᮱�Q��r���a�PYt(�ǽѹ�g�qG���b���������}#��-�d�ӵ-�\D&��_`��ʰ��0��쭴)��^���`��{�ᦞ���֜I|�L��W�e�����ƚ�SY��E�BX�O��R�tW˽�,�v^eq�e��p���8o;��9t�;[��P�_y�pV�zt̤��"�x�%Lu���O����yuO3�(��X#;h:f��	z55�pg�����,4�r[������G74��M����`d�T�Tծ�ڃK��(f-0�&��	��la���TqWKе����5��U�7nֲc1������Ѝ�YJ�@��P�@i�p�n�٢��Sۄ���˚�w]�z!މ��Vw��z�sԪ���tyR	���s���W\�GX����?�6џf�t��f�߶�3�ņDp�;=k���h��B���>�����;iPTg�t�t��yG��E�Z���3��d}`���v��m[������.#D��y
�5�g�[c�r龘���%��$M�HmJ{�l9�r��"bs6�b_P���������oOq���G3{�X~q��{�PKܽ�\sO�ܓ��;!t�t����GW�_�h�'�Zj2��h������M���Rcl����O���g��grY�x���>0�@���z~���	��^��	���C�!�f�Q~���!��Ťv�,}���{�C�{5��Jj�W��5��٬7Gy;�������/����9��!�I"|H"8�S<�m{8:8=�haidS��AD,ͥ^���Y�dDo��������զYm��g��ݏ�v�m��N�ڨ�ك�Kr��ϊ�*.x�]��d}_��׭�f�\�B�Q��v�GsmH��S��,�N[20d�3�it��s�_fC�
AN��R��1��>��ɷ2*��
�^�3cvE�M1';�t����Ј�t��;#]�B))O�ڽT�)t�5�9��2�6]Fon��z<n�▌!����ts��U��/�Q1Jq�;Nf��U����eg#�n�ʊ9:���ٻ邈\����or>�}f]?�^�j��8o�����|}i���S�۫v!yLbl�3���h����ќ�}�������B��u)y����G�EZU7况�H`���叽O��o�����7�]�|��A�1���*}e4i���y\n����.����7t_ChÆ�dfԍ�l���ah!t�-~���ޮ�6���Ӹ�g��L��Ą�NF�Ҥ�t0� 0[r7��]�M-��͋ܮ��Ɯ�+w_x���Y<��+LPwJ�~��+Y_�̺�!~�����2"�s���@��j9Qbjs�R����UC7}S�W���f ���%/ބЌ��y�*�#)��sv^�Z`��:��t�x�t�v��M�0���9L䂎lކ�>�lA�u�kѬ����]��J�-�/���ri����5�Y°��e�����8��Yō��2j�p�[cg���66s;���*Q�tQ��s#!�/��P�߿V�ڝi�ݾ]�O<��j�Jg��j	���O��y�Զ��s��,�������<0�wa�u��[���N��y�n<.k�b7<�䚐m����3{��"����ܮݮ
C&�=
��Z�4a�޾Ĉ9�nd)���;K�|;�l�:��n�d.����^o<�Z��Zr��
ށ7+ZϺ�mI�}�|�{=ܶ��*�3^'�φtjҁ�7���]m���6������1l/tҋх�9粇I��{�T"oU��qj��mAԎ���ٝ]ڄG���f��v==ۤ�g�ml2����q��΂��(��%���q|�LО�4�l)^��NdU���A>��V�+Vȑ�RUp�J_��c�[8�zd�;�n���v[��� ��H[����+���-�w!W�����6g�Yt��y%q�}�.oq3���+}�}�O!4���������]��8��&�&�FR��q��j5��&Csl0�׋m�[u5�87���O���t�BOU�Ues��R1IwH=��(j��c�v�-�0�~����C{ﮋϮ����Q�ʽ�ל���ʭw����w�27)��x����,�0p
`�j��7{k�Ҡ�fד�ͯ{|��W����{���o������|�|�+��["��k��X��]n0�bÑ^'��3��*���:����ÜӴI8��o(w31�S
ZO:�^]��R���
�K;���a�Ǝ�vk}�S�gh�v���>����lqk^�r�b?6>�[b��(����;���`+&��B�VX��8^�A����(���Nǥ��7D�
K��,K�[n�Q��QoC�������ägK�GU�:�[)�;!3F'+6Kf�	���:Lx-�-X9KN���t���5�������M�ͭ�J�I��*Î�u��GKZ$��V;-Y��V=ـ�K�H�����R��p�N�M��}MrыV�B�y㕹�͙�Yβ�Em�X�z[3�ս����Xrλ��]CyX�Q��5��U%D���9k��j��Τ�Z �6~Ͷ芾��S$=��A՞lMh.�&�:����������E��Ǘts��P�&4��B_\��No�w�gn|7�Z�����G!7yy��	��l�D`����ԖJ�ݖc3�4ɐ��K��fV��Aҋ[:��)�
�pQ�YY�����﫥p-ܜV��l1�x��`�]Ւ���/�U�#��S�<��ܫT�����[�.i�D�pLkl��4j���������u��r�e�y�2�u*��n.����q<�+��D�3���S�e�S��s/���s��Ǹ�e�)�|�&�e�^��S8��7s**���!d�<5��]k_Dn���z�|֭�8c����#���8����xk fk����f��F^�A	p;�>s�c�%�(ͬ�ԊnbI�q�1�ҫ寶��".���s�PԨ�A�����~��+�RfĲ=��,<XȞ���1]�_ﳺ:2��uh�F�T`�Z_VhP����[�wARۮ�\O*�{�۷ȐU��.�Ytr��.ed�^���
fV��<fu��f�V��[�n�ڷ���z�28!,q���%:�<2�fŽ�YnΓ�9�S�|��lu -u������Sņ�NF`Z3���X���ߢ7MQ��wCu��.��9��}��I��[o�a�#{�[r�-KzCu9�\%�6�1ed��f۹b�E�w�����te����"� ̹VU�ĽTt+���F���X:qA%o,RŔ�)��Y�\�����t��LUs�<�t62�N���6Y�qD��wZ��2hk���cT����s�z�K�*�Zm����j�q�/*r�v�K�,��JT8�����!�Uۻ�]aj�U�PVP�6�<55n�s�̣O:�'�g,9�U�=�d7��P�jt���*���B�7H$����Wu���7J:Z���K�g�ei�o'�R�C�%�q��6�1�Ӥ�.�*�lXw�T�D�\�^�=l�:Wش�\.����-�lU�j�yE�,�Q����e1�*�8��{ø���JZ)�()�2���)rȪF�(J�B����)
ZiJ��Z��b$�h��$�)(
��
H�!Jj��ՉN���hiJ��
���rJ$"(
B������B��������R�������
Z)J	@R��P��D�@d�4�R��4
J��B���S@VNQS@R���JZ��hMHa#H��P��AJP�+B%%d�	�d�R%d-��((�5��:zz߮���q߮�}_�'w�o<k. Bݫ�<i�5�y5����EҜ��q��W�"��ۗI�/lj�Q.nV�s���ZyW���������vo�S���j�|��R��s(RFDc,��ym������dQ���tn������-=ѽ�Λ`�>c��������]����'���rsN��|�u���8w��r;v�s�쁉�WU�a�u��9��v�/M'���o9X�n��#4�'�$9sg�
\�>��w�o�k������Q��aɐ���m��ʡW]y����W�ʈ�<�Q�O��ҳ��s�[g�̆�c�xX)���M�U�\�Ev0�s5K�������5Оژ�î�n�ĺ��p�� ǟ��k��X�k&�^b��n��M��|�l�V�K.
{*��H��3V����1��&�ލ���oȋ�+��J���8��UA��r�M6hqZ�eM]��z�E�r:}��#ռ�i����"�^zx�T�]^��n��\��y��p��mѫN����w6�K�R�6��!��j�����?�j_q�,]	s�%z򥚙P�DxnG�j��!^'���*+1�U�i&���J�
\��sj��yGW�nZx��Y}�ãbg
N�Øvչ���4r�����3�'�3���G���F��9��ql�SE4WI*�*E[t�5��B/��Utg�62��&��c)�C#΁�7�����M��2u!qw�is��.���|��}�7y�J�����-��>������'k�T�5���ć70Ĝ8�B�:���^��mv�L;!����y�ޑ:�5�;��j Ŝ�[���o"��͵Ir��&�®ڑ�����̈́q��`�q�=�A;1�3���E�#��1G����Q{�:|v����vqlUZ������k�t[@�/�F1���}�|�P/�Eqn��>;j2������̖����ކ�v p�C:³^��Ky��,ā��H!g5d��ƎQ��h�l�Z�u߷���E"���aͥB:�(�w�(M��0��>��qx����'�%�=YJv)��e�X耂Mw㣻���9�a^	z��*Z�yK��l�5��]s��IK�\�E���p����4�#��x ķ�ְn�hY=Φ�;�Z��-ՅAs����C���`t��)=�T̼�v����t1v�NL�R����U\u��k��ծZ����.��(���|�HGs�3�4eu��p� �i#� fڸ�W�X7�l�8�ww����ga���a;ܲcgx���H)
̚3�����7V��O=�E�nE[>����u���T9J4R�����qܼ=��ϳN�l�&��Ow'|�d e�Q�ݑY|��g�����PsB��C�226���7�����k�/�	�.!��v1Z,��2���g�؁�������ć�����zE��&��|���.������?���z�+�εӺ=�}}�ǹi�J�+�t�\� �����|����>�~����������sS�NN�z+LpwJ�~���<�odSQdm�Ƴ�]\Gjj��PC��#�ӽB9Q�&괥������O��m��,5}깛��#n���!$0D�svO��^0WPc�hrI��_� ���/�G�[�3e8�++(k�JY�I�:gN$��,@�v���q>=R�]��멶�;�ևDԻ�D[����Ά�o5K�\o-î�Z�rU�T� �v�,����JZ��9g
ŷ��ժ@�<�
��=�)�ӥd[��pm#��u��e<����J�{��MZ�/p怂,wF����}���\�#쉡�L�ui<me�s/M/b��R2�k�²�u,���u��3�lQ�}�u{�pA2D�n\y��>�22������	)�y�u�Y�r�_vvoQ¯,��'��dO��E-��Npl����p�3*��/Of�c0���]Q5uל�J,�d� ���^R�N����T��0:�0�^���[�*x`��w=_)�k�1k�Y��r	��:ڰ���ͪ�m�S=�-y��5��h͊|"�8@��DGq�]<�+����Df�����M��&$�;�R��駁4�����E$_w���ȥA�^�槨ޭ;:�^8גJ\�{�>ܷS�̉ :B�Ѥ%�6j����t|e�b���($�?Ȯh:W�����# ����g�i���惾���D�Ao%8mj�K?�~�p_��C˺��*�em:�bϒ�3-Iw�̧m�����35t��~7ۮ;ˌ�)��cX)di��9+i�Dv��R�&k.���7�NR��"�:T�����e�o���u�V�Gr;����FR�2�ߛQ��� ��f�nN�dE�y��;�� @Z���r3�5=^�J���T�%�'y���{i�'h��xg�3F�un01-����K{l�Bz���B�q��	��<�]5`-M�6q��K�,+q��7���.|�Z;M*t��mV���ۘ�Y����+��9���)x����So��z��-��A�k[+�~��A�����.6��n䣛��)9��r��Ll�v,&�p-���a�:�y�%�F��L���x��ˌ�����I���=�߱ܧ��*�kHxɃG�}�*�?JQ��oy�嘝$��˚
��!��
N�Vg�5�{:�-���>�,��SW]~���DO�TD;Ռ���1q�٦�&�1ބ�w=�)�a�P�BMw��d\�-Eq�z�����u�AٿĚ���4�������{�ɼ�=hm'�3�HZݜ�z�gZ?:����Zӛj�Ljw��3*~|kj_�X���ג���^������e�]��~���7�J۳�5f�1����8{ ��f��>y�a�X�;�xYj�0�w,�cZ��W�W�����:�-�¼��[q�v�]�B�O_Swi��n���ԱR�<��e])ϖ���<�r9�f�I�}�9�ddE^gX������l��r��8��UO�{,�	��uY���y��Z�:���QAH��q��lD��3�RV^�S�x���7M��Q��2<�}TNt�wl;�����T��"�P(���%r�Rn��j��{ot��b�o]���v���,�}R��Lf�Ψ4Sq���\S[�v+��Is���S�����!qw�J4���a}�lo9[�^��N��n�uor�6��goF!�y�s�� ] ��gCzoC��v����^'�����d���sԴ��
 ��6ȹ�l�:|��.��0���5
s��,@C���ݙzh�r�v�iS��:N�c�;>�x���j��_�f��}R�S�`a�U���=Q:;���)I��dEb�ͺ\�b}��d�����z��4ÔCZ������v�4�Ƴ,[�5��R��YX�ح�eE2��Gl'6t�ֵIw���VdN��Y�Ui#���Uʹ�m��vI�mՃ���0�ζf���gs�^�ٞ�Ù�#ͩ�roK��#�Ϻ���t�L�V��;���O���f�/S�A˱�#�xVkѸ���}f4��Ci���no��W�Vz�+Ȩ�ߋ�n�wWG��T#�(����>��h�������@�;5*+!���b��K>c� ��T��H����O_cc���}���JևO��5䎴�ڛ��(z�a��*�R�B\���`}��:'����7VwVLl� ��()Wǭ��\әjMy4Э����D�i���à��}��V���t
�R�x���ߗ����B�h�Lp���c��έB��V�j��D�p��v�Tz��'Y#��z�FdS6�vF�E�#3GX�]hWSmX먄�^t�g��n\/�8�^���74[|_��/ܣ��	�S�<�2	�>lǁ���!lB��}���3o�6e��+����'�t��y�����r��c!�?]�"�fַ����g%^�U�G���U���Q[�q�"��#�8t�/%��En=����iл�_)\ɎM6v�,L\Dg�z�9h��І4����AU��,a	ڷ[�5�sMA��'G�����b�������l��T���Y�@��S�"a�E�o�����e*jM_��rF(ܻv6��S���5�w,��i8���O�abM�Κ�Tiɺ�:R�-wtW�(UC-��3�kٔ��K�#M�^�1�1BÄ������\���V���u>���צ�Ę�&�^M� �n�h�5���������=6��W��9�y�7'6H�7�	e�?a�2:���`�8GV�W�ݎ ��%{CYP���k�2N���q��A��#5��O4����1�������P�P���;#+%����E�c�lǏ�f��Bz?#��Փ�F�v�b��:�մ�y��j&��׋V�(Q
��S�����<5ih�6)����s��`�h=T�D���L\�Ko�&�vz<`H}�.|&qXqj�נѣ�J�p�/[au�h.��^�(v����ae�XW���;Jz�]��Mv�R�U�l-CM	ҰT��{|����7k`n��؃�P��F~T;h�S�X��:���J'(>�;xo;��BL�蛕�м|�����W���9Ù&��xR����,����U��n喍@����,�w��ε��W�K�7?q}����쟾�MW�[4�L�Р��HV�d.�ˠ��R�mu�-Gu{��+6�%%�x�=�ܧ]w_y��iF��Pȷ��/:Y_f���"���$�$R�d�Cd�S���/��m��sp�����K�3���إU��FR��Wmt]o>����U4��Qu�=&�DQ�Xc��#>�A<��dY����UB��R�h%��o^�E�4�g��^��G��P�D4t���*�2,��o.J��s��������+w�*`�r��[>�`���o{e�u�gj��iM��"��@w��'v7E�foA���'����[#z[�|������+L���g�=ZԸv^�k{�n�^ԑ�'�Td�F�a�h1�a���|~����N-].��Q�.�9��3�w�q�.�]f���j�)iѹ��U��U��kc�7qcǧJ��C��6��d3Fr�Ɨг�t�M��P�9�j6 ���t���\�2u576pͫ��fXn��>P�S��d`��Y��I��!]J��P�����+X+Wd������'�ӖI��J^s�Y�3�������x�O����t^Y�$�I! r�*{#��)<�d<�����,�y|�rg��zJfu�uכ�\���3�c�)g4p�~��}<�Õ'm���ֽبż�z��d0̣q1��ص3����m�����f�O)��tR�l��%��`Ui�8��!�H\��U��'���}��"6#��iIPX�(����K�m!B��ӭURf���f��l`�1D@��M���AH��q)P�US�܍�U�֝�5�+��n-�wX�]!���1�H�4�YxF�)���V�۳�����G29s�=�k�%�`9KkӼ�e�hΒU�WM=8��1.�EC;�0잾�2m� ���,���:��Mcܽ�^�w�����{=��g�������n���f�n1ܛ�R��pYR
���f�5+������yЭ�14���[:�1V�"��t�����T���n4��jv��_��b	H鎸_ѵ�b"^ %U�A�S�G���SFiVm���W�������g��7vS�W�t������`ʈ���63P�u
��Yk�L�o_V]܍��蒣���;��h�D��A����D*6��o���b�V\S�VO��Ě.L�����z���R�`Z��ɣ��a�{�sɼ��%�m� �>�e7x�bl�!����[K�@��.�jMa�o9]�!���J���5��MJ��d�G�E���֒7��z͞����>��aGv�R��0Ȩ�@�����tf�Uf�E�:Ih����w<�����]�b���m��S"�z+=p���#�.s�qIZU�el%�>�fʇ$��j4�yf?c×η}L��|Z�-�/l��^v֬�\�S��kk���q�]'G��lQ���g����:軔F>.n�ž���fQ{���[\�ee�f5�"��s	�cNM(8���S*���$�:�=��S�:�O7��7J��X��[�R�X�x�o ��!"����_gA��U��wv'A��rb� :Kn�ؒ�g�4D��$�a�X{8#�SJ�o�+.+7�c]��n�zK+��G�n����8k�e��ֱk3+W%L��{x.�Nv���
����N����V�q�ܬXi� lv��X������JS���N�&f�Ǵ��`8vҵҸ��S�f��;5�{ ����-�c.Eu��Ym��=F����ƍ}���'+*H����}%��E:4\>�7˻���mZc�]��s-t�3C�i�T��WPxm(�Z�޽�moPFv���;q/-�����r�e��[Q�Pxv�9����U��m�WpQ�o��#�R���E�Q:�f{vi�ka{�fQ�B*��feL�+��8L�9�t�k"�b=�E[VL8ni{Vn���yOX�9���F��U�]ٗ�[�=�/�ӏ�%�B��W��<
��O^Nj�����\�}[��+�0S9��aЕ����f�c��u���1,�vR��\[Ꜵ�Ff���ۢ�E]]-�
���f�"�o+r�-���՘or뭣z�H��Mj�/f��X�]��6�H�s,����Ep��TH�tu�o<�kɝ`Ԓփ[}��%+ct���:ͧ�.�n\Y#�� �Ѳ#!�gڹZ��6��Q����u�h
H�Y;!)��WO�z�޺gD8,SsR�N�1�D+�+��^P�T��)�G�E�^�wle6-�O*�a�Oo�o\�ԝ+��CK�WJks���I�g�M�o�9۶%������:�B��od���ʙK���Cb��C�UqK~J8,k-[�.�34�ː�E+BR�B�M#E+�r��(�
)��&�hJ��bZZ����hi(��h�������
i�)�
b
���i
���)�

J�(&
��
Z��z��Q���hhD�R�%4DR4�KT-15MA��%*P�d)�44��d"�4�RjS5�@��BRДHS�8@QKA�%+���!KJ	I���!AANB�d�HQHБ#�S!�iJ@d)CC�S��5HҵM%��ƺ��<}"W�M�'ʾ�=��%�Ӝp�xbUy&���|�T�:j�1=R�"���K]!O�}��$�X��ȴ�.!!�����zr���k)��(Y-�r�u�%R��~��2��HF^���-�?��(�Sfve�퉕`��N���sV�+w��v�/>���� ����(oC馔5>�r�M�VJ�n���.	�1��Դ����S`�s��g��ਉ#!�@i�3j�e90a2�8<�5�&��S���ޕ��'h3}��ʰ�R�p"wb�1�����t��3�/K��x�A�-�&��@�����;�莮��V �3�]����f��ĳ[w�}�1�`�L������ȟ1�������W��9����?H�B��%�:�(�6n1P�jr���g�4���;�u�J%�Ք���rZ�<���<������l�O��Sz�U��:�Z�m	i��YX�l���i�;�y��.{^NPR�Cv�z�g*1��B����`�ب9aׇ��7f.��3͍Ms�:j��.W#�q��)ط�[��&���k9�t8 ��q^Jޛ:n�f嚽V�(�#˔�M-|ƾ�E��;�l.4r�J�(����]�Ss�Ⓩa�T�ђw[��8��	^_GvMt��dP�F�gc��]��K����ȮƬP*dev��ov����B��G�j�����T9J%(�*�nb*��;6	���Gf�e� 5[�l�����tU��\�_�J_�9T���Ȥ��kˈW|�z�J���S>�uө^���m��s�������2�����"̓�\���㫨�2�u��1ń.����ih��W7����=���Gtt�Ǝ��׹R�~d�k[+�T�7C2���_�&�N��%4�Z<Oۏd54������|��}ܻ���ЈM��=�{Zb�[�t�b��Y��:�>��Uh�59�)���F�U �f�lƧ�q9����<�-
����z�|��;�}zr�r��ղZ�m��2�]�SW}�����>;Cdu��6�����Yl�㹎�<��D5�*����:%�*���~�+�y�΅ԧ�A��q��}��+��zg}�h�:+���7�ο%�vz���}H	t�K�$  a��:��)���[������<7U�uS:p�U����Ìw�e��Mj��ۘ4�ΐ���Oa�
��Y��Eq�i�=�z�3��&���G��5��k�\}45eɣH��lm��`�2��V�E���Lp�o8}$�Y�Fz�㴀���{;����w�D�Wod>��'�e���5vm�O(�u�Öڮ�s��cZ�u�����u���������'Pfl����Z�5e%Q\+]9��W�k�1�H�� ng�-c��P�S�z��W%���y�챷8E��pӭG9ȼU*��J늉s8Yv�w�/��/���6��������M�+LI��fMU��٦@�r+$�����{/7�3�[�1���W�At�,��[��Q[��O����hH�z-����N�<���΋y	��G.�"+�H���}⸌���No��AS�W�Z��뱓ͬ�>s��ú�#�)�FR�2��mF|��[ �6��2��:���5�_l�d�ᄾ��$:�G#"�OU�UVV�����~�,.Y�}�1�4��Ɂ6�*�Det���p��#�gd�-)��HzH�b���c��{��R�1�v���)򻞸��	4VJB�7�W7e�!�umf}ʒzj�cq�&�:QTu�Ƌ���[̝�*�R��Q�/��,��.����㮦x)pH�ټ�Vz\F�l0�`�V�F�T ёg��[hLsN�k'�l��#�z�%EJݐ��z�8�`���5�����Պ�^����*�-�/z�s"� �� ����$Ұ'�<�F�S�5�0ў�#���kw����NongwS����۳����7Z�'�6{�k��*#n�B��6#�n�b$ZgV�1�^6f��$�H9 q�� ���f�F)�g�:ۖk��b��vC�8B���F��u��$��J�tjO�֢�vx里�w.7�����L�}B����6���v/	L㵪�C�f�v�p��}��3ja�ɧ׶���5��P���q%�Lrb����Ęړץ�`�����<�^$�]��/-H��2�8A��+�
���˲r7a����B��hF@�B�ҒX�r�s쫚�>����������Hr���s@����D�x�R�;�6�=����L]]�,�I�LK��&A�K�tS��lo'l�{
���V+C���d1��+6�ml����Ϯ�d��:W��b�	�`f�E�so
�tk=����Wa�L�Ҫ����ڵS�o\>��8x֦0�+��+\�+V�t�]�L%���|��
1�	�ٚ��_V�s5�1���w[[�L$W��41N����پaC���y\[w��~ː�N��P���q�z}e���K^2��yh�&�^����74���ٻ=��&��
p��H����̊�B�!����l�O�����ӯ�A4u_�&W�F^<u�_ym?FqL]�F>�e�3�i�ݜ��H׆%�^�ϩg<����Q�;���ieB�{���|�%'�F�x��y.��t��wL 83"�)>͖��sY[*�u��>q8A�pJ���^�,V�vҢ�q���shų��}#u��d�pAg>�홌e�z_d_#���&�3�ĥ5*���ܳ��i��3��5��� ���ˠ��O8��9�!C�h�Mj�5�^}�ݷ,0r���	g�I�L��L�,�I��S_1:<�ʬ�؆������p���.�ˡ|�/����Ҷ���V�v���]��%�tۜ�A�u�m��X�w���o+f:���R�Wk�m'V�0j�_>�}�w���ʒC)�����nr�ȩf��n�'F�?H�gA�
����}�Nd��u���7ݽ��p�]p��]��BQ1��lS�%��:/,�a,q	q�������"w���;B�2}ܐ������$��i`�e˻H�m��G]n	~�ٌD�\��l=��ī�1���6hE*�q�M��i�b�,�y=�
h��O�#�V��]p�}��T9J;��q3c�Ę��]���1$t������ճ�ӑS�����>��ȿ�6�����q0�Z��2C����T�}��ucK�\HC����o3�^��z8Tb��j�A�.�RXܸכg�q��M�l��`�a25��S��ΜOB�E�qDiE��-֓yN�V�Xe�-kd��R=��̲x-�mڗ�Q�y��f�n0,Ñ�ceuWG
��u�#
�]����#�l��a��\�/J��e�V���CvU�, Ut��_e�4-Uu���Rv�_�:�W�7��Od
쬈Q5��W^\&��[�<�`�-h��'9��vs(�+�KR�&�ك['z�k���5C���d��d��|1�X�o��8�8j����������u��5dq�NM֔�Էz/�9ݯ���9���K�ZdrL)�g���Cz$g�ݗ�V�u4�˱b���L�n���R�ڼv������o�� {�hF����I�^�i<�Q�{rx���G&�c�����0+]@�2~�h1��xF�u�9Ok{���tY���;�O4x�?/�ߍV�ڢ:^��kũ�zym�m��ХPއ�J4�y��L[ڄDw�#N۰嶃��]Ut�F5�k:�)��k҅�=�5蚺�ò�Y@�$+3�n"�Zg_v�m�͙n�wd�+s t��"�P�S�{F���V��Lf`ʝ��zOSuv{X�k�G"�����)>���8s��Y��#����c�	�3����}mݼG?��dٓ^���̞�y�� zg��MJ�����kC��7+�U��I������s�#*��ւ�j'CTog��~���E�JZ|m� ��Y鏸5yxy�/� ���s�K8v�'f�V��X�f�΀t	����$�'GI��-\���o]=���;Z��=�$5oΔ�y��������)_��5⒐�Pߚ#�a>ɓr����G��b~}A��B�\�v1\`gB&�Α\�t�['^�u�f-���S�=��4xkgHQr���;=�eYM�ҕ2��D����%fQ�z�Ύ�{͎���%��K�8�#bM�оJ���]m���>��m�U�����;�A�u (`㱲_��V�z6J��i�L�+*�����I������yW�w�[��u�:�8�`F�y���K�=:���:�r�D�Nv����x��F�j�ի8�J>���l����8����ܐ�j�?^*��fm(�X�!��>6�g#eA?G��3�s��6l1|[� ��J������c�����<5��*E�dm�5�d��#�~�Ŵ�`�|f���_�gb�=]=f�#�ߋ��`<*5x��7E��H���Ȟ�k�UQ����Vz���eJ���}b���\_�%+���X��SN@Ôt���]����gj�Zvd�j�K6�3��ӎc���F����ҫ-`�]�[O������3.pfl#5�i-�}/V]��yQ��p�+���}>�������_(
���*��M�?��-I>�L&�[�N�^��\�J��~�eg���x���H��>��g�����.:�!١�����K.f����gٰ��X�+�)v4���Ĺ�l
�E(��љGd�ݧvtO2}wguȌ�׊F|l�1׀-��SNv�햙Ԣ&���]��z�����VT$"��_.�t�P����T��ۜ����mF'ݣF���0�8��ḢJG[�C�yƘIXc	gx���j�p=�'0�O���N���*<譩��TSWu��p/#r�n�u��3�R��)X�Vn������
p��H���<���mﲻ��?��)�+�;�'
�jx��CӗOz&=�X"��F��0z����䷹��޸���M#��7�<����vG��~�@ k��������m�ZR/+��;ǩg�ܧ�B��� 䞞ŕ(�걪�Ë���;g���������^�Vx�KzׄU��B����+�ᵇ��)�8��&�	,vC[�;���b%�%h�yp<9�u�[km;[��������1��i���W!��H*�n%]��ۆ�N��?��`�*9z��B�>rij+8ME*>�{���7
'�H����{���?������	0�oѭ�"��S����iS�M�䓵�3b�����w�@2`jg9�F����oK��z�xz��q�8�ξQ(n��_��=~��·\`F<�Ѝģ�I���Ʒ�2�n V�(�$����`�;�#!� ��U��B:����!�����U��]!w��	�%�%^�9����o}�����&����X�A����nﶢT�^�O�$$�;�"�c�Uf�Jʻ��wlSX���&�:а�����Ĳw�X��
U�`�s��vO9��"��\9޻�m����B�#�D�`�[:�f��\f���i�E\�績�bY&/��ϖ��!����&E�: ��yo�����yy{=��g�����߻�}��W�z�,��cȹn��2��Md�⯇7S�.,m⽠�! ͩRi͊��(/��#qQ��W�b3F��*��e�w�K�5;]G-�e�8s�a+ikʚ(
,q��5��J�w����}0��d`�w�[T1�1)�aSa&4f�i�S�.]6"�y�f�^�Z[T.�x��^�����Ռ�����YQ��r�':�i]�Q�U�Z�e	���m���*��r-͚4e`X��� ���FԎw"y_e�:֛��P��ҽ(�SgȢ��q{s�N(�*Q�V�Ι+e����.���3�Xu����a��n)���Ŭ�L��*՗�Y�R�� hd-łJh�����x,�ba�z��1ظ8��E��u�/��pe�u-G�d�!��S��n�Kq�Y�dE#�l��"3f���MV�.�L�*Ӡ^�CCZ��v$ڹ�[�P㷖�j��Tü�ǰL�����ee��O��@R��oF���李�L���]�p&��y]; �VQ�z)X_��úfF3$�]yy7enu:���� ��c�)�e�Q\��\z��ub=��}����˫�4�W��؏#���,N�oF���s���׺����n����Bor�P.'�΅vv0����>ugh)��##��]�Sd�:��B�wmq���*�������vX��� �#	�.1|{��۰�a���:7��@�]n���W��G8�]�*������]�X-lz[��*�n��,"hk5�L��P]�|7D���C�Ӽ�B/��*-��u^��u���^�rE��q�z�aKN>f�^v5^���pYk�Y{yI���ɷ-���	;7�N:W��$�m��n*�#�d�S"��x Z�&V�@-w4��.��Z��g�A���7	-��/�MJQw�9�f5�5Ys�$�*�MRI�1��ށ���<��T�w,n�i���l���\nT��Z��r��;�JN�.rj���,H�qJ���m��1���om*'iC\q��\��f��/�������c><�˼;��"Ɨa݀��"�w,,�2N�0=�`��u��+c+��/�]�����vw*�w3�^��̫�J�b\���i�˖�x���ڼ4Z�ițlKZ�
���ı���+��yF��t�QJֱ*-�1L�/O��ͭ9b�}�-������ʏ�{8سv�
\��ӣz�*�5�М2�Fa����Èo��gͅ��ʃ2.�7)7HEH�`����r�+���k^��l�SEh�.a���y��xn#,�Ϻգb����&��v���(������f�ǳ|E�r�ΡV��<R�nm����pn�k#Q����q�4���]�ҷ��Ԛ��)g�v](u�0�A�9�c���u2fu��ΐ�3-���gVj���D��j��v���ڧG�z�K����2�p��\�X�ɨ,q�&]k��\u���(Z�r
F�V�JA����u.�)
P�(�(rr��!�&��4��E)@dd
"P<FIIB�S$[12MY(R�HP94-.Cf&�!u
�ffT%&Jd4�����-AF��j�uJ�j
JG$���!i�*���G!bD�(r�(�b���KMjD�2ZJ@�1%dB4&�2u �S!R��kX�Y)0d	��o�˿-^7�rr����yj����}Sq�\�����|�**��j����O\^�ė�m�V�׌9Һ�Wu[���'%��ݴ7�僚{��;Ŝ��?Q���-m���<-������L�L���Շbt�_f���ͤѦRVr�M��8���6Fc��w�䕈5�Q���qGi�:lt��H)��2#�2/��hYM Ħ�R�`2ص����X�n����������D��G��S=���L�-y�H�����a�)Y�&��7���+��Pw��1�.n��;}���6u?,MIҖ>�]���{�ZtW`;]�pj\m(U���=#6�
6#�&�Ҋᑯ%�j��_33M4Y��E�4�%�U�,6�׺�tg��|�!t?b6���|T����|�m�vf�o����z����I~;Gz��g��b*R�Л���-��u�N��}=t�q^�tY�oi�;���zXیY�:�:�v_{n�a�cDh쇍M�V�{4ǯ�	�H�q�[<���_V酇Up���+�.�Ť�Qm5���=�{!�`;�̏u"�r��y��6HU�~�y\�,b=���ž�{y,�<t��Θ7�Ɲe8��Rť�iR��v�`ǘ�^�Q��[�v �\�̻A��dH0Z�k�GR�ۻ���X5M��e+��D�w+KO��v�D��^�� h
��$;�0���.< �-��3)�^�-�Q����u#��j��tM��z���-�t����U`�i���3��&�:Ǫ�%���sA߅�J�wZ3�2���ns�W%��R�u�Hɳ&��;�=4�5~tC�~uT��sU��V=�B�o���W��`�#^))sƚ�`������"\Z�Ά�ٽ��������b"��΄M�W6Ir��[G_>7�sO�F���u>8�!��t�d���eYM=	-2���1�t7�q��K3��n��]=,1�K�
���\��f����OT�E9ʳTνg��Dm��'�A�xM��Î��+��2�s[�)1��Z��Z���5�ϛz�s6����1R�d+���7��oS������>Q��v�hU�2���Z���,F�53ta�G�ۆ�%I��q����[�x���X��O�
^s�^�{�Ԟk/��f�K���L��f{���c�`Vb/.<��=F�����.���v�����\�)��moG��;�=ӳ.�-j{sU�̺��Տ��S�U�J�j���J®[#o��=�d�鷕����	��L�"�.���yܳ�'��n�FH��6Q�"�AA��`�g�uP�vw}z�A�8Y~��y}O
R/ m�4L�H6e��	�|W"-ٌMI툍î�����ד9�j�e�Q|�G�����A���j���*�,����նw^�y��ח�d�c�IH:�����=�T0O֧uu���Y�D
��}�8���H���/Ca�
�$Rp��m3d��U�N����ׇ�Ǣw��PR����\ә�hݛ��r�����lGe H̀�8H[��8�D)%�)�;5�w�\�'Z�N^rNm=���0�m���Zx9���
�"}|�y�R5B��%-��0χ����lF�pp=�rC�܍��p��Dd�t�����3�RM����A���Cn�6��dK@�ݽ@�V�r�WS}��U����U�"6ͻ�:ǖ�0�̆�V�#����S�3��C�Y[5A���i�啺����m�
ia}��#�l��C��ڜ�՗RƿCA��.V�X���xh�7�9m�-	b��[8�JJx���^�$q'����u~�pE2+zy�Dd�oDs�V>kW,i��2nN_o1�'���m�d,���,�aN����cȦշPҙ������v��ZP�rhZM �؝4uYD���̌�m�ú��_�]���b7��pK�@��[4����{�/>����;��O�0j1�(��Aڪڎ��"��X+zDl�*C�QҖqD�W�[��Nh��h�}��Wb�����ͭbϪ��0s�0b3ۓ{Ԩ9Z;ah��n��ط���v.���G��hGHm�����琂-�_^��设���E�V2��I��:&�n�w2��n��1�E���w^a�Y����7�T�s�(��sw�g7E��$$i��(��?Ld���6i�M[�ƚ�1ݳ�$��]Qה�:������V!4�y��tS��yv�����s�?j��#Z���K���N�\��qoqZË�"�o�˴y���C��n����Y�ʒ��`b��X�o�n�dsô��a��Ļ`掓<A�J�{�V)]�j��ݟCB���%8 г�|G��X�˹���l�]v�L�iN�y����X�ջ<��(^�O�$'��q�i#���!cDd6FUE[��{���n��qA\@{�4�d>��!my���݌�|l�:���VD{��^H��3A�UlOeA"ޛ��ݷYA3��w��i����Ғ��
zd�^�u���p�S�yH��֞��ɕç��svV`�}y�K�k��ҍ���EOێ�u#K� �^�ؙ��n�ZW�6����Î�#"��2�|�\�d�u z���l��Rk�5�Dt���0&#1z4��}
k�u��yR�a�ŭl����sD�ܿ��&;'o��qM7 [�v����MO_(�X�W$`"xAdq��38toT-E�'`�m��o�2��^]��f���0��	�����oC�����IT�����x��oG���ݕ��V��#��ꮒ���JX��/*5���;c���g�e�;�%�lJ�Ash��{���U`�B�Lp`��1x��T9X2p�P�PnG.I+�i�vs��qݖ���g%�i��Ap]`�R�ہ���L�^���h�G7-��(�VՌ�:L�+.�nv�F����vD��?��V����ǏQ�=A�{|��3-w���8]ȉ��ܯߵ#[��+f�=@��%1ԟ��ڑ�@��N�t�΁�~����ji@�}�hЋH����7Ӧ8H�L��E�P/ߴ�Zv�OfF{2>�v���_����Z9��,��'��A��3�����'nz���Lfk�oC]j���H�`�!F�����;#$����Kmj�6T�@n�7�E]T�K=��P�S�g�����3���
:��H�ݵd�mA�$u����ÚY�����5]��6�f���X�?p�������B�X��2\���Ήx�S�d]�۰��5d��e�J��� V�[��%`�#@����=��D=ذ�E]rc��9�O����u0� �o��*��B@�1���c��G}靳���f
W��c]�Y�Ōtl���9R^���������j�8��ZN�)��f�Y��[Bz]��Jus,݅�����Y���u������Z� �"2XYI6�,yj��&_^<I�n�J$G`��Q�[[C�6F�@9��
�δ��c���^���]چ���ዧ7l��/DU�$T��f?�p�t�`���*�����I75Bj�戓Bs��n�m�Ǝ��nmi�b��}�z{�^a.+%�.��dY��;O�"ok$��wݼ�	j�����R��ce0�@��\]�o�x���[�[���/�^�\�g��x�]�(Jݔ�����a>CL��цh&��Z�};������DbF���S�s�Z��Ǻ����[Cg��n��w������յ�v�֞�p��F<�lnk;�1�n�ъ3��u^��|͸��"���e^EƑ�����J�#O|��o� m�$��p}w�����5�GaN���� �A�=>�ndt3��}a�Q�x����v�R.]�%g=��]:f��o�;w�%!˛
�k���tG���&yk]ɠ�Q�*tl���䆭��":��Yy5e.�Z�;���y�-�f�����	�s��bO^��A��.�iu^Y=h������G2�|��;BE�o�;AA���8��v�fmu��R�Ӵ6��b��/b��tj�d��tI֥^uh��]��n�QA�2H�ܨH�f�͝�=���Ld��.F�K���O$�E婹�.b����.;3e����"D��z<�8ĸFDg����,R�u��7��A�c�6�kA%��m0y�:m�[Z���BB=]�O��H�AH���f'�n�̞;M�v�t�@GT���1�%�O��"2a��b6��֝�©�� E���yڴ��Ύ~���	%P}�.�X8"�Ίڝ���}gچ���*��q�U�ʡ:N7_�|l�Kl0������Xr�1�[v{��������%��P���č4uYD���eζ�v�j�3��Ѻ�=�0�/0��C�#Cf��9mP�ȥ���vM�&�
�k4%}s�bsku��h���-������QҖqD�mSKo7kn[���z6y��:M'��s����_��o�*�����6�K+��B?ח~h���~��[P��~��j�b>��+b�6��)V:H�Cf�k�#`Q[E�͙���������֋���y�_`�nX�"�V��r�3,�Z�GVa&Do53,^��ې�Y��oC-�������͠_bD�gK�p���v��6[�"��򺩓�G�Y��:A����h�B0�fDc,��|~�۹�q��{>u�۪�~�ų�Ɏ��3��5��
`��Qo�Tm�N��Ѡ������^�m���	=��=�(��?H�fv�%��*��eq٢�����	��67������8��	D�VR��dE�H�Ӣ/.���Y��P�h0��5R/����ևOD<�=�W�qj����z)��o�]7F�=v���^U�VLl�x��vimwVj��_�q�1��`A���[�z�ni����UA��]��>N����"�6難wo����h�)GA���n�U��.��X'��W@�%�o��K�f�(�"-#:����Q��UO�t�F�;!0q �k���"v�q�?�ïm����a%�7.5�=<yu����m�M��+��L_��(!�S���5˒�}�WGQ�GRY�|�� 3aph�yRl�;�}=Q�˰WP������[b�*C�q�{6�Fw��Κ��*���H)���gJ۴^�N]�qL�^�_3��޼�eIR��]u����盾�ݗ��t��`��.����}
@�M�IO*�.E�{��S�U���UN^Z�1��f�T�������އW�g��S�o�h��g/BNvku�w_��5(+�>=� `��kC7˷θϣgUG-[Y
6ᒋQTwlə7�ѧ�w�Q��P��H�`��#4��
,��h&Q:ƺ�aF�cs8��u+�j��.�A<vF����2�fwr�T�R1�"�o[�n!|v}e�_eW&�����rC�S�l���M��-p�KN�VR��Ý�~�������[F�����'��i⼢�p5;�	��r���B��}xJC�Z6��)��"w����R��粕�z��-�{���?�lzs��a:(�ݢ�76��<�K�ĵ���}�X/�m/@c����������(hH��������?�����'���@ � Q�������(��~��4gLOF��0e�f &�eY�f�ed`Y�f &�FdY�	�f�U�eY�fQ� �Ve�f� &Q�`Y�fU�e�fU��eY�f�e�f�VV``Y�f &� �a`X`e�fSa�f�0�1�a�f�a�f�d�fA��Fd�f�`�f�a�fA�`�fA�A�����u˂�  O8��2��( L 0��   L*&0 ���0�Ȃ �L�2 �L�2 ��� c�U\` 	�U�PeUf �Y�U�UY� 0��*�2 � *�2��*�2��*��:�
�0�ʪ�*���� 0��02���0,ȳ*�0�ȳ"̀L��u:E�V`Y�f� �V`Y�f��� �`Y�f &�F`Y���?��_O����@+0����`�O�s����?��?���K���9���������~I����q��_�UU����~����PEy�ʪ��@���>�O�_�?q�C���1UTW�?,?`}?�z�@g�w������O8?��}��a@@V$@
U�UbP $�U��U�� $d Y � %BVA� !%U`$ !  RVa �U�Q��*�#��E������?�TEE�J

 �>�ϙ��V|�AA����}�;�_  �����C��?�x�$~|�����:c��N��UUEvj�>����O% W�*����>��䢠���~�� z��L���gC�Z0 �����|�G?����8�8UUEo����說����P}z������>���A���$���?��  
�}������UQ_�.��>�!�R}W����N���X��?��<x�y�I��ʪ�+�uA}�T��pӸ4ϵ��=m~H*��x}��Ǯ@T\���N�����bz��d�Mf=��99f�A@��̟\�ؽ�������ё4Ԧ��H�R"J�IU%U*HRBJ(��%U&�֡Q�hjJ$�)%RR	E� TmY^�ݶ�2K[kVj�mJ���PLՙki1M6YJ�cZͪ�uݥ��m3�f�Z�Z�ف�٬�6ҭ��D���V�f�[j͓-�,�K�L�׷vM(�u�ն�R3n�9IQ�̵kSR�I-U-�[$mf�ٕ��ь�۵j�-�խ�e*-�m�j�2�Q26kmc[�����im���m֬��m��}�� �m�]ۮ��B6�˽{�]�ޗjn��z�s�z�=z�n��m�@t�+�����A�v��uMԯ{۩���޴���[ڝ:�)�z�h���ٽ\��+OC{�k�dT�&��["�k5�� ��СB�
A��/�=>�
(P���P� P�B��{�xz(P��g׷�vz����M=ۻ���v�O4�筻{���c��ځl������ӽ�חn�z䧭뱚�5J�M4�b�hlْ�  s�}w`����ӆ�:������ת����nN�{����k��g�z�کJ����ܫv:=V^�q��S����ҷS���=�Ot���wz�y�)���OM������5�MdY��m�  ��}:�l����w���zum��h[zu�G����{���8�����n��7t�C��N�G�vU4ۭ8�ր���t:̌ �j[DƶR֨��j�eZW� �z�cMs��A�Y:pU�ge9Z�Ӫ�{��Ͷ��wsS�6B�5 �V��ON�o:(h³� ��Y����m�fHJ����� �{:��ZM��:���kj���5�l#CER���k�1u� :�7u�J���W-�t]�keV�N����V٦�Y���b�X�d� �x���ە;J 3v˺뵀-v�
:4�Y����G�L��S[QY@�b��  ;�7�����P�:S��Vյ*�̉��2BZj)�� s��} s�n  ���@n��[����^��� t����4�@@��� �z�x��t� N��^i�Q��h��j�5��x  >ﷸ� ���  �v� ��u�@;�7���Ѫz���  z��� [��� �Ӏ  �u34�V�հj�[1K��y�  x�� +� i�w�� ��� ����z
��  n��ւ���z Q�:�� ��"��JT�5  S�d�)J�  ���%)P  � ԥSQ���"oH*Pb @�"&5T� �O������*?��?�?����7�����B��Y��m�UG�Jv�Yn5~��{�f�{ފɝ;�T_DU��W��T_悠�¢*�y���\�:��2����=�2,�w
���hF�<˺����ݖ�J��!ɡh(+�5��5t���a�Y(�62mѡ��w0��v�f�5X/&l��P�����)�36ed�+�$�Ò�E��d��P�p�G�{c]c�Z\����w%�J�*�K�-�ʛ�a˔Y�߮-�(T�3ocj�G��%(4�R��ņT�e����+MզӘ�B�1���QƆ�T݈�m�Ҝ�	0^�ª�h���w�*����N��������m�&���a( ᩉHnӠ��G��+
WHyp������s�Av�ZA�-�uc4���/��Eb�N��bQ��3X[Ij��*ټ�M	m�-h���X����6�9��%7���NL�[y���b�]<,�Z����c��1g�e�E�qUB&�7$k�ƭ.;��]�Td�(kU���өf��{R��$�Εmf⣃2iͭ����i� �5�c�A4ঋ;�J݀�k��"V��t����l�n�ɹD�fTc3@-��.�mP�4P;x�3�� ۫(��I=����0�72�J5��T�Ա�F�p���컥�%ME�?y�P��S8�w�g�.9��S�)bo���c�j��SQ�7��5�'vk(L̛�J�u�0ig��xQ%g�@��sa�0E`1�(�Z� yn��'*�1P`h4�R��_\F�l	�73ti�v����X �&�O+/#ܵVCʺ�	�,�FHPڒ��Iޢq�+d��ls32I ݬ��gN�v��`	����*�1Q��5
�H�ip:TX�L�u��.o���5�
y �A��,ȵJBe�gT��� ^]����q�4��W`�L��'VU�q�쭑�30D��[-և%^��i�4Z-6 e:�)�6�Y���F�>�QAR��Y�n:F���*aZr�w.
n���mDɊ���#+4�<�t�,ݪ�I��ҫ7��i�*E�ۋ���G0�q�إ�YH2�ل�	�љSZh|V������bf\0������c-ږ^֘�)�ț,��d봆hv��#�b5P�3S{Y��FM��l�+S�����)��-�;��͔�TlW�J1�0����	Ttv���ޤ���!eK�t�	Zeԍ�0\wfT�V.�y�b� 9`�Z{�9
�f���T6!WX�X�B;9�Zv�L�fw�Vj��L�ʴ��d�	�U�ER�h(لj���6��5����2q^
ĥ�A��C��`*��h(ɖ��9,�lm'ZM�kM5N�R��A�X�4>�2�/s%K4p;���-*�Ө������
� �K��j��Ea�u����x���K�c�M�hF���J�"��0bMLsh:j�Ħ�f]Ҍ��.�y���(�B�Ҭ�-���Y[���{[L�%�*�-�e�X�*G]�-��L�f�^�y��w��7˅i�)HE�Y��)n�c��\m��H���2J,y�4F���@`���]�ܴFS�sl뀻�n�fl�&�x���ʱDV"���KT,:1�ۺeS�Ob�JY��jk�M����'*��.A	ӭ��[�AT���:�a�� 6/�0��n�:�G)��o*��hx.]Tgiӳ�li8�!W�hHul$/��6��Ԡ�U���0��µQ����1!1o�b Yuz���{��^���m�FΛ�[Qmk�rJ��Z���;0:�tfꨍ�����wiQ�j�k:^E�������na�ڻ8N�*T������
<=Q�"��w��ʗ���m)y��K��=�4Kt%�+�f�1b���-Pk��kX����T!]k�mF�%�*M�nA{S>v������%C�uҠ�Ȝܭ1�1�	9Q���6��6lP���.;�B��!ԕɩ��FųJr���7J;���`��4g�ڡT"f̴����1���t�����kwMc�J�&��V��W�Һ8�������f\��@GJfҖ�̋M1(�<��ܲ�i�n��@ ڼ��;�%�A�m�jB�76�1檑�@�y>5	�[ò]J�d�\mQ�@(^}��T&��U#fbۋ]O��Qֿ�Ҋ���mZ�Kv��[S�ǩXe�(`�\� ���R� ��
ur��É�Yf���ŊG�eI6��Z�0@/>K��\�����6ث�n˅XS`�N7u���k2��&���fңw��}I5���2X^���P���X��W�Ϭ���-���3+/nh�1C��E��U������%�G5�%�P;P��tA�kM�0,i��x��ۆ���\��V��
��{�Z#Qݿ��bb�e��C/+(c(#L����2F'X��U��%id��ݕ�Ni� lF`�or�m�޻�2�rB����
W&L�d.�'�4̂�k>�SӍ:̑-ܘq�L����n�%7IFh![�����iH�� m3E���c7��OMdn�K9��K�dC�.Xf�:y�*6n���W�7u�K����@ZTt݊�̌�	�Տ1�T$��(s֦�����8�K5+B�P��=�Ϸ+0�W��)p^h2�Mӕ2�C��^&[t+��76�!B�CQ� 7
V�X��ь�jJ�e֔4�n[�G�J��űu`2z"��Y+b��V�uV��_��Q��:��(jX�#6��l�Byov�d�D�F^c*�n�s4c)]dy�3W�R�"�D2$�F��1Kɴ�T7�)���%jP��[8���)�4���u���D���U����H�^iZ4�Q����u��2�� �J�u��"mk��� �ݦ�0C墣�n��ˁ�IU�۽C��/��f҄�+p�*(B@�9S,�X"�tl�2�&!`E��lzhYߍ�%����BDh�&S͔Nh"D@��N��qò�Z�gt�b+.]�B��妅���,kuulij���$a����IO�|܇*��m�
�eH���d�U`��,�W���)�&H��/2�a�{u�"�9�`�WVn��^iù�Y.|M8�,�5��t�7L��Zsh=��K3Sr*��zмIF��.�r��%��y1n*z�&/V��ܳ�i�i�
E�%eʕ1q�wf�=*�Q����i�������A;���F��:	"�ű�.��i2	�6��%R�����Y*�2oX������=�J���n�
��;gI��X���YN\�e� GE��oe����/�lJ��ӕ�so�u+8�!M����&\.��g/)�������%n�ͽ��P�ݳ&aPTɄM�*V:��!�qKȶK�4�e�S2ޖ�D��F�Ae���X���[t� ��^��+$���&�ݣN�Ki��I�f̤��E�̲�̐[[e�*J�[Lk����r�z�H@ے�m1��Séfn��&��$�+͂T�f�lS�4[8*"��iG�Ț n��T���M>l�pմ�%�àՊtܔ�Zr�]�w5��W��Z��f�ʶ������6��X���ȱ["؄o�a�����+)B��U�J�Җ
RM���ô�
� `Xε�$��G�R��V9��׎D�6�4��w�6��S��V�,��r��E��L�5)��e��˹O�>��R��=QP�x����Q�n�մvcww��Ac�(eK [r��Ć[ɗ��,3ZK�ݺ���x�W���t���"���'�3w+L��ǒ��[%\8��H���8�)y�*4�#�Tvm�(XY 7��E���-%mJN���ݝV��6��NEZ�+Ȩ�n��3tf9,��-�@y(L_\rꄦ��fE��P���sE�0���p�:'S��j�-�YU�����#^�>ĔlƎ<O1��qKv�7�'͋��j�3�VsJ�y��A)��$���U�v��,��-��\�JO��'c]��gmw��$��M�iӡon��@5��dJ����هwfܙ�*373"P�r��}tNL9v�`623�����.Hoh����.�-��+rdZ�B�8S�Y�.�1[b�Aoh�1�Z��܁��nl��jXϳh�!�%;VG���S�T�|���Q1��(̊*��U��mպmЕͳ�L��|)�.��Y���°��6�����K&0�L1�q�&��:��|F����i.�w�`�0L��l
�h������*e���"�V^h��N������"��qD��6�Pv�6����^�W��Bm\�����I��V�C�r;�m�7`|� 74k��r�f��j��<ʷ
�ږF�1�T�8A�5T�' ���B��H�J��]�b��&l���5ֺ,�iPORWz��mg�"�C�� �Av�d��L�������^fX���Pf�U�%E"�I���H��Da˕�*e�df 	��\S�'[�w����:y��%Y��GW�ceHY��ƒ��ᠴ��IZ����{1@U�cf�46^Pt�n��T��n���K-8P���Y6�6��4kN5��u�36��P�:$�
W3!1�u��bfG�v6�YS>�V��D�e52=�v]C�vM�5�W����$���[OS?5�6���AIt�tU��Ȳ�j�C���suе2�ޡ�Ŵ�AW��FI�&[�I�E�mn�Y+w�S!J�:ŀIY�j�4���6��ݧ�B�Ѵ����ĢsC��cC�8]�/��陛��[g���e˲^|�=.�(�+�M��d�
�2J'(Xj�Mܢ)��E��S�K�Y��ѨЗ�.�L�F)V݊.��l�bʼ�5X�ܣw�[�+�j�؂�2�3L�v��oc�yn��0�輼��0܇C4@�k�.nSݙV	y@=:�l��7hc{���l��N\b=,F�)�!*�W�[F���ᰝ��Nkr,�e���P��`1�2a+S ��2�&e��+D�/�-���A[1B"Z����6��D�TV%e3,���
�n�
���mǮѽmr���Z7r���`�eY�T��dn#7"7��� �jA��\��Ùn�`i�2�����&��0ƈ'trm��@Ֆ�7ZxN=0��lH��1<����V�4#˩��ۂ�4�leXڈJ"�=Iq��X��]�L�ʘ7 �h�؞�Ie�N�Y����jk�[��ˊC��1ല�DJ�S<k�w	ւ�"��$U��+�8NX�ȧL+���bƮ]��0��:S�ތ#��N|+E�ؑ�r�}5
zf��;�<�֧���՛41�Tu4Sɳ%oj��[���̙���U��#�FR�4.�8�xt�9�z�0L����Ȋ�ک�]�or��dȬ*j�G������,Ve�
������J���j���9�IrHpcXZƂ:���:��c�$YӍ)���5WYD��.�i*Ͳ$�t�2�[)�n��KU�aiGQZ6�.�c�He�v�Vo$�-�5h��$hӥm3Gtl٬���K�������s&�&�l*�V)Yv*���Gr��I��"A�eH@���������e����d-�f�w
��
k)��8����Um!��� t��nQ`���3)��\&�?��J������-e=ܭ��W�2�C�2��x�f�Se&��qK�A^f-O���!Hed{��hͼ��٦.MעQ��=Y%��ȯ-�V>6�F�u�u{*XZYd\u!���jN`�YF�����2���GZ؉�M+�0b�`:��&��hX�WFi��qΫ͵ۚAk )��R}�
7�PN�iv�d��a�d�Թ2���
:�@SJ���ݍW��]G.(2��e����D,J�l4�e �J�9q�v���/30L�y#te�(SƑ��c�+2@���+ի5Xq7e<�&6�P�X�<����TƼ[5��j����SUlC����.�ӹ�U<����j����(5Q��r���0nI0����֮[8T���IL�X��r�Z�j��� i�6�7xo2�&�#�j���.����<�/d��$�}��SV�DHN��X@֙�q]",�����/+N3!��
�M
 
���L�xB�o>� 
r��i�|�5[.	�e1{���C���Zu�J�,���W`�0h�7|��0�eYуw@J�\e+��6����"�{�P-ɢ�7  �F�e�-x�^R�Ŗ�f� p�BnfB^�{D*J�@�n����n�B��Y�VB��6�K.����LX��죹�/Y�n�hN}�0P�ib%�ԙ�I���KT\7.H^N��W�L��g}� ^rWMU�{dm+�B��ҡ�n"�2 e��z5���9d��p\F��eL�,�M�Į��j��Iq�[���j�\���ͰF�96^V�SMj74�3M`�I���H r�@�*TX.�Xl�X:/\ou�&���K��W��Sdd(E�r�0Y�`,��p�x�WL��yN𽿆b-�L�m-,G�+ql����c�ͻ��*N!A6��y0�Hi�MyTi}r�S7g�m�:�Snn6�!�#w�k�+{�S!�/���t1M��&&f��-,c4��Qm=���Ќ�����&��Z���7$��0�zf�jhm�Ρ�U���t9��WPfP����B�B�6� ]�Y%ۙ�A�k�&�˖[�a���ּ��ט��
ԕ�S��.K�3UJb�
	�@�kh�i��M���B�̀(�7);4�FK�!�iKiU���W�,���I��iD�,�b�*f�(g�R���{˨��~�/�<�&���^ہ:X^.Gd�ӳ1�*�l4\wMp-N�@ũE��iޗ]�����5Ɠ'j��������5sq��,���Y��V&�|�`�����,�Z�Y�"[�5ں]���8~��p9�´���Sp|hF�z�D���	=�sV^ �'մ��K(�6�
ֈ��.��X#�}ODԜO8�˦��0v�7Y�s�A(��7 �#�Y%�WY�-u�7@O��X"l���7����k�
��[G����U-�mJB�6Q!p�M��sz9ø��U��{! hA�iL�m%*"����3���ܻ>j�����?=�}V Y�L��Ԇ��g����uk��1�NR��ݳ������G�b-��=��|:�.ZFf��&Jx�e15�Pa+f�9�S�J��K��Uكg�'M��S#v�r����+��5��C�i�۹f�
SZ��ij*���_1t�u������óY�u���oFp���p���J�㋀�/H�jZqv�"�a�C#���z
�n��e���88w}1�&��J�Q)@�55�W�tw{W��")be/�;dSOkM `P��6����MC���k�ڭ�RTܔʦ�	�����i�˙ӱVǿe(f�q�e���vc��[A���󔢾ʈާ�Fq��u<m���Tn�j�q����ڤ��<���횪��܄���ن�X��R��^{���Xހ;m��%����V�Q��Vb]\'Dt؇���v͗G)���Y�ȯm�[��Gʤ��m�;;K㋺��У��ʱ�#�C}����
.�:���vXݚ�>N�w!�\���n�hډT�h�6N�|�g\�;�7rʝ�ĥw@S)a��`�	�t��:v�Ö��R�ʎ
&V���mG(�!
Ur[��ku��7����6^�����9�7��ȼ�զ��G�U�b�	�:�&�ɤ0���I7/�x�=���X�+�����׮[.]!���ww�	�n�s���)*&o�e��9%E���N�sr�NgY�H�+DI��m�5:�K}P�v2F�u�,s��/1�X5ð��$�iu����D%�->�.A7w{)�x �'^t��gV����4{ko9��R��5�J3�u%B��M���{�(r���>/33�.[���8�o�����z0�jg`N���E4�ǡ�,��uvG۰7���7��}5�̺�n�@����/{�+�vk�1]w$�s)G�H��;[R�g�%X��+w4Q��hȺ��u�f�����w��.D�E΅�
�h��H`�֏?���9��!"��[��\y$�w�6�i���ܸ�S��|�	�
T�H�SeAܚ=Yr�J�ud髠�+&H��
yϮ�kYX�s���+�����v7(�U�+/Mʔ���m�c���@�pg+�p����8�{3�����]��˱�B��S�([5&�G�ؘ��8� �[p��R̳����9��]F�tʜ��JΥ�S�.��}JMr���>��OV.�?m#�0��WR�:���ہl�k�u�-XH�w5�ت^�IX������Q&���u��i�h9d�}�{���i��D��Ll����3�^���l�F�c�;���'cb�Y{���w3�CaΒr�7-��/+7�iS9:i����fZ����>�f����8���H�ɓj�rjȹ ��98��ڍgaP�����@������0�r$5�[J��W+��4~�Ŧ��ѐky�*�%��f'��Z�4�e�*��"���\���t ��!P�c�.�U9d]�sx��e�ݎٓ{s_Es��C5�RN��x,��[q�9�9��f�K	��}�S���O�so7�+3PD������LrFj�4]C����r5���+f�Б��T��b�t��C�������S����Yj:�6�D8ZR�w�N��[�e9h�c%�)�7r��R�rc�U6�|1,L�E�K�7D]ݩ�� �euEM���;�V�-���B���!����x=��VIs�.�Q�v@h��R���JW�S�;�9���Z"��LNū���9�&}�m&Ur��[����ݷ�;�����Y�N�� ���"��
���	�-8�����r������MSEg(z�^i�姕�Rs v�w Ux�hw'Ó���S�]����R��o�.�)܌��.V�(rw'D7��&'2�ZY�G��1�٧_�$���f�b*��D�;^�"��#�N����U�N���zj�Ǖ+��.��ck^���e<�d�+|�VtX����1�r��hln�uШ�HEZ�Wc�e��ꮝe�G[0�>��_�n8���[wy�ޥ�s	<8슶�m�=7��]3\�'M*,�
��F{��OitP��] \rl����yu� �j��r�ܼ2mX!��.)6a0Nq�i.�@뻦�<eJ�lM��{������Z�n�D֔
Yv5��C�<rZEu�J�@ݷ��E���� `ٌ�],�a�5�JS<�qL����ٗ��(����;Im(���`�Q����-��V��q
L&�j&l8�D����6���et�Њ�_���ȻOEQ$�wV"}A��7wիa�q�D�`cd�u�����@ᦥ��x�Q?���O^��C�u�0A���X{%u��ˮ�"�d"�IgX5·��$:ե��vf
�\Ãm�t__m;u�f̹�'m5�G^��JEm��gM"0�$#2�/�Z�����*�Y85V�Ӧ���ɶ�]�2��Й{�����R�\9(��WaP�(19{w��G@��Luee�`����)	��.F�7W0�*J���O S�O5/�2���x��6���i'/C<�eɸb�:�����4﬙9��<����)]�2�%Y�l|zUk�o,ک���<W%"j�4��#�kKj�3�����>�Aw[��mnƮ�,ݨ�4�L2p�9������^����:<Ĩ��sm޻<E�Xw��t�:c\����z�:S[t��{7�!Ȯ���j��S���p]@d���f�$o��;��Fl�7u��X�޼��'gl��|Dz��Cxuue���U�0�yһ�`���U̓�-y����;y��6(yU���fSy<����:`2y2�aв�s�}1[��# �Pժgn�����Am���'���Z[�)�~H��e����,���Ⱥwmi��U\5e������(�S��)Aݤ��R�u��r��FD$����S).�X��ֵ4J�z�p�������`lhY�-�>�f)���i�w�4f]�i %��H6�,���+5�)�'�EZܡٹa��s)mI���d�u��V	���".Tu��;���[���f�*�s��W&�*���qm���3p�oe�jw8C芓+
U2��5����V��o��!�N�\�(��'f�t�.���95-Z�'N:��b�)���;V���itW�F�����WЧ�hB%>W{��ڶ��N&c:cjw*\fh=�h���̅>�ҷ�4��-b�V�}��T��	���e��0���*����λ2a3{n Z��8�}��T'9���Z���oH�-�/,}�3�Gv�l���V�w��򤪒���P蔜I�a�Ay�A>��9����kقi r5&��Ufde��l2J�5��̨��o{A�u��1)Ն��f�i�b��cE�;��t4��5��A;+�f	�ce�x�����U�Վ���P��b� X�";��Z�JE}���G��L���n�]#t��Jh�t��Q499���_:��5���^�FU��;dFF�F�)��qq�[w(�Xt�C����4�h���'�A�q܈6Z�'���Yor�]�8�)H�xP�Ғ��**��B��)���"����z4�T����Q>l�F�}���<�8���SL@1�9L��ə�ܩKȷl&��[ܱ��n� kF�'� �nq�8���G��z���x%<X�g$r%������̖c�9�'37-��������n�M���b��CI�g�<�2QT���ۓk�Yt��[��e�P�˕���B�4J.�AL�c�ڭ��V�+er6�v�J�7�}i��s�I�l��JJ�l�^C�!o�n�{Lwd�x*D���:��*�9��B3 uv�����:������blM��C`6�YT��z�vt��:�Va���z�%��~��=����g�x���Kk��8���`d�;�(�YQ�s�J2��phyد�Q7F���god�8�%���� Hu�#���W��Q�G��c���63165�N���QT�Gp���w�1j(��V�˼��
,�4��I�[�ݚ�|<�/"��-WZ�Fv��F�^49+�9�T��E�Զ��AP��FH���,­R3�9���OT��n����9�n��Y�|��-@P�!��2,��:׉�Yp�N��-��2��_n�������Ǧ��p�VH�rĭ���xv,�9E�)�N���,.y}`!n菞����6m�Xn֥�9.b���W�P��bЎ66Y�om�ƒe�gi��<ntJ�K�MZ��������_0_n�Ф�s���;�vO�B!�\l�ޫ�tE�����U�j�IN�o�x^��Kk�}�nio5��Y�ʹ0���.w�aG.PC�O$���X霪�,
��K�L��g��'ŉ�{Ͳ�zesżi��}\yeP\��6L�w>�q|�Uol[ԝvA72Y�s��p���g1j�p�x���9kt:�c���k{Xg��9�ALW`�{4��Tm�;e���P-Ψg�(�.�X�),X�Q��[�xs����_=�;(`Eɵ�X���Jg]K;Z�������°@u����2/t.��ܺ8��dɪT��K��8�-]&��m�u�۱(R�7�ΰ���G*�.�9�U�A�����|�v����5��-+J�;T���j��#x�N�oM��H����ޝ�=�ĤԲ���JxVI��@l|1%sљ�57�ٛg��1nјJN�c=LjcӨ�A��ԛD�h����*��{moC�̶��Uxgӡ(�S=�V�������ƽz+�a�p qǢ0��U�\�����k*@����t��A�E�h���G��X�aVu�H	�u%As��:�fƦt�j���=��)؜���	�dz��	�کM嵃�w�qVN��%t�Q���ux^s9`�6jJ��	�j��YIӓ�)C���ԉ�R�a�8CYr��FN;D`��onN�κ+C�`�+��e�����;u�0ke�*�ъ�(�	.a֗-���'�u ����L;�j�^�k��Y�	�%e0�>"RH��S��]7��"�2�e՗ѹIhy!{�%,��-em�C��s8���-B]h7��"�.b&���)�]C���TH�+|�&��2p�E��"G&bG/-�Ux���yڅ�;���C	��r�vC�/ ��yY�m0�PZơ���
�o�(є��``�z��Y2��E��j�������<uY�oQ�����ĳ�@'Jۼ�|gJpL�5+�xw�lCy�������EH�� <��R��0��S�3�'�bѕMEs�
c<rT�I�8c!��ڻ�l>�)x��e�X��Skm6;�"�xwG!��M�lT�ͼ�
*�>���+��W�^ �����)��D	��v%֖���^	,ީ.%��oX3U��ۧ%���45Hr4�V�e�Ԓ!��]��i.�E�����gj�.4���P����B�dr��f�L�k��7X���SBz1��m,�.����=r������]� �"?N�RS�4�ƕ^_�z�=S+1l\�٥�g{^�dk/7;��C
�L��3����j�E�����Ӯ�Z��f�d웒��UY��jH^E:��4����D����V
�t�H���1Sj�[����	:�^8��0���	uu�q���ځ�;x��Z�e6+P�{��.��q��싷a�a�M10�7[AGY���@��]l���1��mJ0�{�h;��P̈́���Z4t���4��QD����8CĚ�ϱn�gurlR��*;:�l�Yilާ$s]kZ�7�c�����D�ތ9�#=FfJ�C��c��'�kP[���̈́J��v\[��;)V�ӝ}��lO2Dp��A�;-MA�F���"�']W;tA��UYJ�����pu���ʜb�����Y�oz!���C�g9NW"�e�It�ʴ�]>���e�V���	�&/�x7�d���Gbr�ܴ��VuJmY����6sPg=��
3yb>�ޛ�a�M��� �++H�N�r�R0L��I��+��V^�Ƚ�sz�>��)�sA��)u���N���1ޫ��K9LFV��͛2��!��b��s2�Ǡ���&ǵ.�W�pEyϤ�U��T�:u���t��3Ar�[��;�%!9�6�:�)su�ڨ�Cf)Oe�91:̫yҾ&��s���fKW]X��YDq]��Y�\�&��\�GB��l�T�$>��θ�\E��u��k��ѥ�>�+�����S�Q�'2K��Nt�[S�Ɋ�-�8���e�4�������+k)�c��|Ј{�'V����ܝ��	W5Vc�{{\L�nF���
���ȯ�ٳ���;҄5L�D�"��N����sq���Wp�:�`pފO�o�����o�sf�֔�x%BY�.���w��u�F��7�*�<�\�
朡�c
�o��=���1��p��MZ�����dJ-S&l���7���7���1{�NXV���i٠Cݫ�m�f�p�v��:�A���;�.L2I׉L�w��?�EQO�PEw���w��w�܂�Y����T�T��둭�����2;��ݞ�j�����J�	R��x]`:�]��]�]2)=]X"�Z��ױP]��R�Ɂl�C�g(����7u@���`%;=;�ͬ�r�%��+b��Nn���*d{2V�l���5�jd�ӫ!��
�[N�b�Ғ���,�=�Yd�SP�A9";�;WZV�`i�'n�j�3L�U��)n�{V��V���8���k�z%r��G�p���H�޸����5EmF^��^jF&`�i`�mRr^]L���^u( ����:%y��CSos\����:��]J�t�Y�6�!X�����O��hʜ���������ժ"S@V$P�4�&�)�nek��j��v��C葥5�v��um�0��\�!�:�Z>����̇�����UgY[E.�3��\K%��T��ݒ#����X&]]q]	KQ�p�r�Y�}[e	a���9�t�Ɯ/6㬬��#N��j����#&��]���H�6��M����ͣZ/�R�R�UG�9N���y
�F���l�����ݽ�u��]�7�H��%E�^��1�Ӟ,�A�n��[s�ar�2�U�\�����%��L����b�/*�~�,.��^�d�bۗg0�w����yvSY��j-�a��[���c�X�7D�;;���o0��%�0]���%�euF�Lٺ�\w9֡�frS��|���LJ�a�M�ś��´����Ek�A�6�Ψ��#�P)^��)�}�pw�jY�:b�2��7%���];0P�sT ^����
u���i�!Ҏ�W��W�3���p�c_W;����W��]���÷�0�.T��c=EmmLm�s�x�I}�\��Z�UoxIf�wJ� �6��e��#�n��d�Y�B����������pQ��n��,)ϣA�w����:�!�g��f.ŰdX�me*�V�+sz�I�;��꺋N�j���7Wi�҆:���ǥ�%��7��A"Qh����=c����+-텴Z��]:ʗS� �T�s6�%J#-�G@�RSS�v$�4kJ�ن�m��ɣS��\x��leN]fej��uZ�YbYbU6�c�&���ә�\�^N�壍N]&`[ێ��s8/�q媷^�:�nf��%Ҟk$�WB�/v�w��[f
h� (�¡ܭ�{qF�hT�����٥Wgө����z<�|���D�D������X��厚W;��e����R���h��i���y�kRM�{tEP'�;��rR�j�n����Z�ɻWY5��{4.ٌeM�$*3�LZ,=Jf������\b��wZ���Cyi� ��L�1�d�쬋5ܳ
�yk,� v��t��w��f����Q��u:�+ǍZ��U�At�	�]��P��ut��o�v�0�f�ZrFN��Y��Ĥ�u4;~��Z�H�,�p��6�A��res(q5ʲ�꽛3�Qu�k�4���?rD��� gTAz,e�%�+����Y6-��p&W-��#sw�{w�]5�*�Z��,�����L�g�n�0M��%޳E��:�W|_P̵dt@������t*�hJ�������=Xiq�%�!Z���G
jA�Zx���;Xut�r����]z`�獑
F�(�I�뺊+-[�s���E�l����Ka��opV�]�Є�6�3%'�:�a�:�)�ua]h��Ғ�|�����Α �uo=pSI�,w�]�$�SX3�da�� ��E�U%�y�Y�j�J��r#;btnX�M��Q�ӑ�aٻP��]+��V�t�Yŵ�U�z��}�mN咒�&l�d������{�!h��oi.�b��-��;}�h����[9�5�-��Νֶ�8�U9N��|�un뚲��}��� 1��Êg+=�S?�ERb>љ��5��SanU�94k՝\�"���k)�&:�Tά�Ӡ�EAz7\`-�uv�Y�@	�/WJUq�:9����z���q��v��Xފ�����wx��!��_Nf.�u.}X:� O��vr�-��$�HE�N�jY2�M�)�]x�\�;��c�O���$�1�\.,�����*�;6���+�2۫hY����!��z7&ظe-���a�s���F̱(�k����59�ɑ�V,��sl�������$�/	\�ȳt��D�8o�^�H���z�XF�R�?>,��d��Vw�MF�����̃�L7U;::�MM���,0W�p�� H�>�}�cb�QT�'����5)�U�ˋ��ξ3e:v�''�_�ڵ��5jn]0{z�q���	��qVn().;���h$�FٷY1_N8���N0d�&ռ�|	M�	��(M��=��C��M�V����u�\uʦ3�����P��JƢ6���Cz��VeN]L�7�Iv2J�B��w3k�fQᲶbԱ�%�ŖwuSu>����S[�F�_K��z�Gel�M��O{��-jň�F�`�Nج��p����j�������b��1SL���f'�0Pt��p�[�Z4o=�f�5�wQ�*^���ݻ�ݪUA:9��&��@`{!�MV9'sY�Ryǻ�wY�Qr�W��+Y�[#�"�y::�r����� �8�sm;5�nE�zr�	������.�}�M"(\�ʻsy}y@�����i2��HMA�i��tx)#z9��A>[�s \�̠Kg2�s%m@�u�aQ�,��Ȩ@r��c<�%��-��'@�M�[�%�N7a2��Wt)�^7��(a�U1��U��钲�mt��9��>ш�t��GkW3�+#���.XCu�M+;�ti\%9q�����/q
\��5����VC���z^J���u�J���@�fof�,C3]c�%���ڜf��V�a&�L��֥�ۼW����u]��R!������}�:���{V�ۮ��謬�8�.���n�)hAQ՚�{���6�}q�H�R��r����Mh���7T�z%�$�PJ�����\i������Ktv�r�W�(z�n�m s+BSU�h)gu�k(o����+���е��I8��G�p�G�)��[Y�9�(�WG�E�I��쒶R�vC�If���H�E��6��TB��1����v�t��x����|���b�b�0���b�,5��	m�nnWP�7�&�����е��(f.���`Ҵ�4�bo%�8�`zrc����!��#'^l�)�1G�X��U�<�,d�U�9���4:�����n>ں�C�m�w�e��������R'1�r��t�4�s/��W��hZ�1ڱ8�s �C�)Gòj�&-]��ɘ9���x�j�ۀ,���w���84���JQD��Q�e坔��}����Љ�Q9�U��f�LVl�G.�?���V[�ӫa;����>3&v�>u�s�ԫ�����^�5�����b�A흛ϵ�Eȍ�g�� �˗Vl�Y�6$�I���e����ӻ����֝T�Aד%���V���ݖ�/���!�'|�:F�Ƃ"ͥ)�C�>k���V�NYx�8�."�i�.b�eKrn��ofb��w�u)MrT�L��c`�"�H��t����F��T�̢9L=vmu���MbKw,�Eev�B�ޡ�b�vl��]�̅���y9�ʜ��D�R!��4��2�p��鴽��b|��֎��;c�)�IYs��q��i��d�z{Smɂ�1Q˩SZwvq�A�J��% 䮋/�V��n�; �D&�����7|e8�sY�l�$��Ν�t��G)M1X����1��S�=�H�������91N�k�ڮ'��'����-ꑼ������:���S�*W��gC�R��8������,�f2����V�J}L���r�_փ�i���.@�<A�f�Ej��qΌ��o�Bh	��Jx��Wa�2u=��x�EϤW��*47rFs��m`��|�V�3�N���܌�'img)gNs73VV>�;��H�$�8+  횹b���J���zuY�Jwi�����+�+h�%�V��(7N(]���u,ͩR�<��W%���(Q�V�'�T�.��]�d�4���4�^f�W�#LelJ�En�۵[B�՞D��(�?p=yMR�	�u��"���x,ߡ��	�Kt�����H�^�a�H��/�oM'�+6�D8���
+�Z�v�Ra���5��&Pz��oGЗS{	WW�W[�t0��Ь��EyX�w	�VC�M�B��ƹX(�����C��3N�P�ve>�Ge�[ΐ���#�����5�gkк*�uiR�C{f�7(r�ԪN3��v�m��)��4e#�"�
�V,G���4`YCv��z	�Ϋ�'XRL�ۡǙn'��|�q֨�Ur�1/�ɭ����w:wj��L�c���3ƋE��f� P�#4�]p�ˌ�"sLz� ҅<UQ��,%F�����6�j�\Z�:>�p�՝N�W��{��Mya�^g1�9��V���Ц�q�t�Js�zy�|'Ӡԫ_$���A[�6��p i;z��WP��eE�fB�d�����&
!L��;�-���p�t�-��E&$K�F�j*�(h��wv����Ws�.v�=P���ϡq�B'�̓��^���\vv����H��'(�>4�������c]^ͮ���ad��1�y$K2�o�P���+Q+�B��	=��oT��b��&�wkX�rN���C�w;��(E�zt�ov�I=E��%fM�@�Y��a��B	O"��,Eb���j��8��عm�c����.si���-D5�Т�]�[���B�G̼LRy�t噋��.bM̒P�5G)���ۦ�|�o�e�"=�����q3�u7_;Γ�F�&ɩ�[7y4�j�#�aW�ue.�x1,RG]^,D�o>z	�o_ �e�3vRd1@5�������]J�L�����6�pa�泺���2u5�C��K����IpM�hWP�����x+����PB��N��V���v�U
n�t����U��KW����ֳ!��]K�G�emZ��x�I��U��$]C��	��z���G)�Q��Uck5�)^���}4�k��L�gk�aZj��nlo)�t���_ʘس4b��2G����nZGv�ۜI�ԭcD�M��I�ƙ��-t�MV�B�-����1�]
�������ʧ�E�5v�S�q^�蠈�ͥ� dU�J�829��:�I<w���c�tÇ-�_dw��^�M1уk��u�������΢j�"��1�5��n
�:�
��-TRc� ���܎H��	�u'0)q8tE�2�Û�蹩ԩ�R�໎U��i���V�g:�^36�eS�e�T�d}t�#�{\"�J2V�v�FO?��{��ur���qwd.�k�l��F�WsڕxLtk�"E�2�SN�=���4���V��8_=t5�0՜Jy��*Vs%A�$*`�qm�.,z�w��>p�`�m+�D�64�Ew���,9c�n鬤5Z. KO],v&С|����K�`IĊ#�r��{
и!M7;��=�gv�R�&��-;�a�ܘ�ʒ��c�&/�q�JX]��*�ޖFfS*��i�ǲq̣�T�q���o3rˮg�F%J�N��N�묷	ͥ��BB�G�[�kv�m��#e�0�;k�ƆW���km$�c�M�b�%��I���Ow]��6�T}\�U�Mr�_m��Bby/�.zj�+� OZb��u��#�N�!��V��ykJ0�o�֧�#�@�C�QZ��bd�ځ�	�MY1��i�I��������x`!N�ڊ�smd�b�r���ѭ��z��P@�>�ͼt9�v�m�+S��Z*�)���-��rT�W<�WnB7/�cүWh5׬c
���:T��\�l˶o�L܋S��T���:�3/�u�R�/�L�Ԟ5�A[7t�ؙ������b�r��C9�e�ժR�
�SYcz�)�7�vL�}��,�(EA�u)��v�&]�$�ӄt;;Fa�K��(b�I���*��(�P��Ȇ�T���]�v��-0�7����2��1��}��".��yDn���I&K�fD�i[�[��%f�Z�q�+�������o6��Vd��H��t3k)']$6/���Me;Ml�+6�H�#f-��n�*_agm��Ȇd˰WVƍ� ��KF�F�:h>�iTI���Y�K�4�1J�j�w�ri�:!��wG)��	�5�/\�/�h:��zS��B�GK���$pY��#�z�J���1���|��2q�7)|�W*,Zty��'��Ta#hv�u۔��Uy0n�G:�̒��O��t8�}��u�miaNv�]�Ĥ���q�x�X�}X@�o��R�q�
t�yGf�YL��#�� V�jߢ取�	�-���B�qܬ
[��V��=8s��oI�m���>�XN]����dԷXU��U�4�#����I�D����v$�����7�L��Lh�du|%�͹1�m�Y7���]kПe�'���n�^"�,7�i�{2�ui_.�g����As�q.B�t"�����5�p�teU�.��]t�l�l���t�r�^b��)�7;^mf]��o{
�B�=ӕ���8��CcP	B)Bѝ¬Vo"�b)�emuq�S�Z�Gl� f�Ø7MmJ�n�.ș��VM��l9'^g�#[d��e���Ñ5)\���*�q�C%&V�j�;�wf�T�E�"%쿝
�c>��9Nqٖ�;l �W�������9�VL+K����tV���PE{\����g�����o{�hٿ<4�7�`ۛ]O��XVT�:D,tU��Ŗg'�,�u�/+�v�6�+�cY��c�3n�ZP�ph$���j⏂U�x7ps��t+[ܼw��ɪ@%X�k�N���ںlCԋ���K+
�}��]2�X�;�������yINTYSU��ɴ��,ܭ�wl+�fq�ى��s��w.}R�d���8gC]R�L�DA���ӊ�ѩ�΍.:��R]��ۖ���R�]��7��]M� �3+p/��X�oeeJKV]��̙K&H��m�ޜ6A��oH�D�,�cw@b����tu�E�:h=*Lφ�;�s,�ݘ��Ӄ)��Y��62�?X+͏P]WW�$5�Wo$ؕ����O����)h4!ײe
%��l���u�>��[�.�a�CzgBCQg2�`+T�s9e4\��ӫ���v���&m�ח1�G��}����P8�
D�{�]�TNl����bc��,2����Y�EZHI7c�!ꎝ��[dԧ���{ھ\�c&k� ��Ye�y)b�A:�k�;�S�,��R�=]�RI|��ȳ6������.�;��Ub��3�-rlɐ[��lY2��%��;o����B�[q��_Wrڣ�����t:�5]�#���-�L�^Չ�O��8�U�PxO�aFz%���҉YJ�E/l,��HG���PN��?vw{����k�:�C�
i���)h���(ZJ �)
B�h)J���i����hj�)"(�
��bV��
T�)
B��JJ
B�*�R�hJ*���"(
(�)iJ
i��� �
(b�(J�����()�%)(�)j����&F���b%&
��������
)j&� �"����ZB"��%�)(����
)��Z�h
�����"�
��B�����*���b
JJ�"�ų�~���׽y�w����d�,I%���םPAvl<;�N`ފj�F���&(��劗�z.(bX�֩�n�J���G�'nq;1�n]�����FgqHb5�Z�K�NsT���T�]ܺ�\F��B�^�x�i���\�<���qX�u�onW��#+��}2��P���T,�ZOOajt�86��M�a��]�F�+E�w�X��*��&��'Rؘ;UFfC"��R��$_˯���NW��S�eͧ�T"�u��i����GǏ��F��{��a��''.;k��J�.����qϛ���Y���W��N�T�j�Pon�[I��gU�a��U ���g.���=�_Z��h����;n�LY浾��IF7�w(�D�3?X��tC����R�9ݏ�d�G��O)��X�*���K��b���!���~�ۤ2�BN��B��u�W�uZj/����1�/�@�yC��.��_+�Ễ�\�Lm�Ɏ�(v�P�|�]u�xeKT|SR��U��`죺��B](P���㜤2���~Cm�B�4��l= 0��:y�]�b�a�MαݡJ
�X��jjOk��݁�Η2����H�����@���pij@u �+(�f����I�ke�"�Y�Ⱥ�Xrf묺�VB����%�(R{0�ƋH�ar�+c����X2�㨴��y�g2y�Lp�\�0�=�I9�FWrQkp��Uk9I�ƾr��=v��FQ���NaT*J5�@����S6:V�-���A���&W)�GDw؝p���@y���']������	g�{�-hh��6���j֮(��R>f��p���'}��z]"b�7�*d�.�7ĵ�WV]��w�F�y���[N���G�!+���h�m��C�kd�;��C�f�&�mz[���� �P02�7N��'�@}��/#n)�|C��-�ڲPQj�Lc�C{�%+���THxy�G��@o��6V�d�ۮ;b��W��e{�ҝ���w�Kjo���8/|xvZ�.Drwh�k��5%�ۄ�l�qxV��@r�t��=��>Iݯq���c�UKW[�_��&�����߭N>�[<��j���a�]�k8��,0��EFu�t]3�e9���Cl�m��/:��]C�8��:�(jhn�)=��ea���ۯ.�n�m��F�3J��H�,ՀL�;Ȉ ]���e8��;u��)��'������*]�9@
Go
�Ba;]� �7�T��K͵�τF�"n���9���c|r\�N�Q0��WGXrw�W��h6�vs�x�Wk W�,����ۥ�G¦�.)���:�Q���ޢο��t���Ĭ�M�fK+�I��g/v�˥Qc��n
��� �3RD"��Ge��8[Z 
�N.�*�rW�d�Ei���>��;����M�(���@bI���#n����c���:s˴��a.���t��,^�g�*����1���h9W�k�-���.���]yr�{ࠫ�߭�ɘ�7�KT�u9�[����g[Ux�3�D
�BS!��r���Jw��Ww�X�grB�a#x���n�H�U,`��ь�r0�	\��@U�L�vܥ<&cy��C3��W�����XO�|�j��c���**�|�_��p�{lk�ĉ׻"��cI��Q��o�BL\ �y��1��ط�d;^ոG�[�m�.�;OgZ�]�\As�9�`7	��.��QQ"g-H@�,O��W�X���]�jx���1���EMu�-��"�/>
�eL��F�7u�cT���v�d�
Y��v�X�Lo��:���
�'FO|��k���-t�#7a9,���j��Urw��:x5�K��'�:�u�R��ѝ�t�h%\��6���w�s���4p����!�hF�'B@����f����&u(I����N�p��c�1BK�N-����h���V5Vi�feC�oJu���,+��HYT��z���6���ݚ2*�k�ac+e��_'w"�`)��KF�ϔ#S9�-�&��JSa����XN��u�[��J,�}r�>ަ0(�VX�����C5�5-gM���w�VY�ʾ����ĉ�j�(|L@��]�]r��J���so����cN�/�H��We2��ٗ�|Ѹ���v��z*#�0E�KTf|�ʟf*"��>t����XC=Zs���\z!�{p��s,�1������l�![f�{�Y�{@}(+R&i<h���CW=��<�A9ò�Wj��S̰r�g�*xF�¬���C�l({*�>t*�����#���,]"�k�"� k�>��*-C�!2��>2�4f�[�W����� κ}�=8Ϫ�Z>�l�p^�|��]����S~����e����mds�Q�3��X�wd����#a�^c��6�m���t�o�}��~�נ�H�][W���p��Q�3w_s�-�����	� ��%�za"�M�cq<�/���Gr�e��ģ���'�� ��f����3��A=�(��z�ۡ���PI}��L��DY��z�\�[U^��ӄ�_D�zN��w:u����\��(���S�<�on
+�ܾ���K�(��̘�P��9.�Ĭ��绫]�Bq��^����g��-*a�ӟBrm|�܌���3Jd[@i�~D_�ܾeIpZ:�f�SO��	ܲ�85�W�N�1��R!����9:�dR�)M���-&�V�!T�2��Me���9�m��7����W.�Ϝ�e��c*ï�1/^vh���[��[�Jbf;��0F���]��}ԃ�j�1pT�Q�2^@r�כ��i��c8n�go�}PE/N�	�KU��=ӕ���U�m�Q�屍��:b�n3V��O<q�:�^ 48ܝKςʱ��:Y=P�I������Y�{���w1l�F����Ű��5JD'��NB�@:s�6��OѰ�O��
��	qw��җ9��~�<�bRzr� z{=�5��]�^b�Ӽg�:�J�TΰxR���8�0��<"�k��nK��Oo:���J��|'O����Ʋ.UC�N#�ҹ6�pQ���`a�)F-�]�IޒnsQ�L�h���_U�a��@1q���s�'��y���/�h�_�nU�I�x+.������/��i����^�_��pN�5Vbf�C�ɾ�E�j�T(D{�lL5­���˵�a�,R���v:�;PgIy�uI���&30��Qu��t�mD��_K�m��n�L{�y�,���1�v�X��tfUl��ԕ�;2������ �
�X�;J@K�s�^�}���0H;S��憆���=I�t}���Jc�p��zV�`��7�����nF�L Q�J�2.��Q��zܜ�)��U���yq��3�1�9Z:�&8 I�J ��R�ۆ�3�n���3t�y�A��n�PQC���T��r|t|�?k��\2��WQ�Q0+�سl��"�7�)�m]�y��굜����|�.9봏20��c�sB�RQ����a�5З|(Ԩ����D=$^̦�v )������͔59�&ۨ8^��VE�fs��x���{�~��~�gV�ldc�k��Ψ#�MZ�D���1}Ne�R累�9=��!	[.�|���@�к:�T��3��u������.�=�aU�ws�s{��m(�-�
���@�ʍ�S�P��"x����f�!<4��jڦrt}akn����F����Q"�Y<ɢې5��۱|b�3�L#���x!���Ll���z��u���H؎��+N����B4F�
=٠r�R��v��#��_f��Kt�hϴd�R�e⥫m�S�M��~��k�4��	�;�p�7���ѧ@s}[��_^i���f���.��X�T��i�g��s�ǲ_K0n,���!��A�9����i�ا��aYח9;�c5�̚�y,N�w�x;3gc����1�˧}�L�j?g-5}F��4�௺�i1�PxdXa����1�Wǫ*�X�U��I�a�-�9�j���=���y�+�aTOu5��]C�2�#9	�3�D-Q.�WU��"����c��KӰ�Ķ-�aT���?��X3�� ;�w�QR�OwW�*q��1+X��˞)�e�!��mR ���)�p�9=3�n�W#�'F:���X�h����2�c�}ϯ�5W&��i�(��i�&~`ДM��c�t=�c����L8�t$�B�_+�e���i�e:u�q��<Ѓ8Z��F��,�̞��w�x*�cZel���]t�_Wo��ν����gjW��b6��w�UuMFr���x��`X/�Ⱦ��������U,`����F5�g]U����#�سY�rLZ���(�<�m�&�%*�l̬Ȅk����n���"����
N��:��'�kT���-��L%ͧ�{���m����<�s�P��t�D/���]K�|�f<��Q
��n���C#x�mY;���9�M�Zo���y�����:|�Rs��놊����]�m^M1�YJ�[�F;���\3Q+d��Rq�W�����ڨ�~n�F'\@ҡ��2=rY�[�]����u���g?74ͱϹbG���H�.tCg ���7z�Պ*�$L�e���¯7��ۨŕ����Eێ���h��9�R�����.�F�nc�0�K� �SJfEB04��w��;�o�~�	�{R�}5ƃ�na�g�i��:���
��vd�b1�UQ���7Fns�Z��(U����9�o0I�Pw�*Y�~�P8���dAІ�F�����r,3I�M�ݲ{q,�����>^٢_cLi�(5{��A���f�Uuצ��nւ���T�%R[���k�����8տ��a�e�˥��MXW<��\�9M51�0\gJdl	�m�*�N;�U{q)K�C�2^�����U19����
m�~�,��9�(�C0q�l���o{�d�'K��"{\<U\�&$[8�Wھ�?:1�>�'��R}�r�b���;���w��߬���,��l����`�L�EOݸU�h�V4�sz.،sW�NJW���d���B:��a�#�:�kd�s�׾ 8�p	��T.&����0�~>�b��;P�G���x�ܮt
q3�����rf��"��%�-+݇��kf��5P��Kʾ�f��Vs^E>�Y�Qn�X�F�'|-�3�\�����|W��WL�k�C+|��o��W֡�')�ȧ\u�6��n�<�x�����*��8*�d=i�a��@�?*���,��ތ�\L!�ym�-��~����)�l��}X��Uk#a��<��l3\�鵹2ˉg���:I��r�������$��C���Mo��u^�hm����d��j0T"�"��ET��_Ê���qF�E��q7Y�7�1�q95��摞���P�!��p�//��~d.٬<�v[�����xF7�b���:l�������P��9pꙐ�)O+kY��M	ܶ�R3?la!�o���Z�cr��9��r�aWQE��P��U�C�Q8�x���sm��z%�D�@�����:�����wR�֮C=|jw�1&������[�!�CΧ��:����TEh�9��_��R��[Mez�*֫���j��l�||yVA�����t�� 1_',/ʱg�6.�=�C��Z:.�k��v��j��zd�3Rm������f��Zܛ��f��ޏ`	�.�p���+��L7�\�*�+�72��6	9�[��k��(���`�c�ճ��b�j.�.n0��M�v�!�jn�m��˯�m�qt�լ�gM�ǵs#F�(]gg+�\u^���PG8������˝ ��D���yv/��,��ׅpF�uC��b��p�]"̜�#(5�����:�<sz[7���ٕ�*w��N�y*S:�]*c��I��*���b��c�f��Ӿ�����Q�������H
�k!��t���u8��x��apR�}�^ʕ�/��p��f(`�.��U�
�>�xn���P�I�I;�[�L��ζ�5�ܷﻶ�6}��⮡Y2`nȽ.�-�a�1RkmP	`�v>���"&�8��06\,�	s���B+7zSyLG9�gD�}�R���hC#8�ǭȫ\�*�uԼ3���knq� ��[Sӟi����O���i���&�	:�(��t���qփ�D�|�(��0��,�"�	�\����!��#O�m}o��i`�t�� xy��HNq!`�n�\�]h�ٛ�2���3�M�Ɯ���=v��r4���W�aU{ٵ�O_8��].9�tD�I���;<���S�*1:��U�6P܄븑����k�ߗ�7B`�[q�kC-�%�]<u�K|�L��]
r\I�Fz�`��c����TH�֋2��0"�"4J��9
�a�v>�6�3���)h9�+�̺�Ih�tNF��G%n�w��C-��5�>�p�<����y��U��,�K���m_*!��4�۝J+8���9�C��.��f��t�z���� ��9�SZ#<k���]�S�ٕw�}o;�}S��Q:Z��5��kW�MÄ��+! �p��N���E*�]��z֢�6/�XS!f	sM�:2�op ��ޤ����:H�Z��-;�ä��᮹/(M�h]�7Ty�I��:063�h�L��m��,.�����^�[Ez�z���b�,�\f]�>�w�\���ň&k˒�@Բ�齒C��;Y�����ƥ��
]I+����	`����mL���s.����iD�ۜ�����{�jz�f����0�\�Њf�쾳�T�t�XWh��s3�6k�Z� Tu�:�U�:�J��~݃��%C��>��x`���t�ſnd��|mM�b��o��jJ�f���L�i��<ܬ��M��zʽ356��M�VF���|�v�v�C+���t����@4g35�-;�yuL枢���� k�c��TW_U��u5+��f�fi%l���T��^b��zO3/H�&ǐ���%r��*�j�wԠq��G5we
�N'�C0_ �6`)䝽u�Y�/AU3���+߳��n���v-���'��'Z(*���戹׿[�P5����s+�M�� �Bm+��ޏZR�_X��s�W��9u̜h���۸侌 �,�:�D�[z��-I����֓����=�:��"��g#
�
N�/A�u�/�S�֑�,.���V;6���;��Zvn,fPO\Y�8�K��v�Y��PC4-;7���tm�w�m���Y�e
�+gWɊr�3 �ڹ�:�@,�m��MNh�g1�;��]�:�B�7ʥ1	?YVa�����٣�M��ٔĭ��q��`��n�;Fgʜ7 ;gz���C`���7\-����9�/jd�5+�������Wm��rJͤ�@�k�u��&Ǝ��jh��"�O�;n�.�9�]�*��[�w���8K�f���X�ٍeG��_wQ��}<����D��4��]r]J��o�f!��=Y��Jߋ:Ms�ZP^��]�����Բ�ū�)���E7՜A8sk��غdH��?*�rSΏ<N�Vu��;f�%��[�5'�>\���|�U��Z��S��,f��u��1��*�$�K�اp�tE�kd&R���v���B�P�Mv����x��s��uW[Οv@�'����I���]2K̬&" ۻ3�YD�j�hi�eM[��9�}�f��ԩ���k��L=��C¦L�:��J㾳:�	i��hj����Y�
f)����h(�b�����*���� (��!��J��)�*���h�����"�*d�

"�ZX��"hj�
)*��hb"f"��
B���J*���j�d� �(��"b��(i�&��bh�j!(��*���"��&"����J)��%��i)����J��&"�����(&(�h �H�i���j`������&(��(��������J�&*ff���(���**���&&������(w�5�����y���r[{0�|G�J�S;1��@���ީIXʑ+̚��xOw^u�g7z���#�5Z���fc�����/}������I�5����5	Ty&EG�j`��2~����w��5	[���pz�Pw�z�{.s��f��K�>��>�t�\��2:��mX��|DC���p�?g� V(�Q�W~<���u�n��{�/e�k��΄�|�3�`wr;��qѬKX<�4�'Fa�����]��w�'n���G!�5g��7?G�j=���78#� �#�ȯJu#!�◹�^��B^�q=���r7.�����u>˚ǐ�3��A��繗y���{�#'`uu������pZ�%%�K���OF��Mԅ&��G�X��1��]{)o���}�o�;���A�j����{:��~��`��;s�P�����߸<�Q��uw�iyI�d{r���ywpd�����]F���j�5/�����"!�0>�����n���9����������NN��{�u��b�uRO�<�.���Ƽ���-I������S����I�����9���A�럴��	�����_��5}�{�M�D�7pǫ�Z����:˻���k���.}��ø7	~��;�7S�\��:4a쿭O�r:}�A�:��Q���<�n�˒�����L�K�{�]//c�%?���^��SO��<�"�DJ1������K�e��/=�p�Թ�ˇ0�?I�nѨ;|����Q�f�*���������%��a�k�亃�kA�d��5��;?{��~�'%Ύ��]HP����'L|�D��BO֫}���˸�g���n��~�������RS��4nz�!�<�~<�~�u!Os�u�p�X=��n~�S�<���P��s�����P�N��5�2�����^C�����2L�#���}ϻ�{ʷ�w�;��y������w��8u�u�^F���7����K�o�i�]�yG��'s��\���������:�P�:� ��������=�s�u�bɏ��`�#�<�It܀�9�{����]{����Z(=����sHo�'�3�\�Q�~�O����>O��P�G��s\�{�/0�y�}�%��<��r����;;���K��F���}�.A�8l���u��kVu�4�s������'�b���YESR��n��g��0?م��Q��Y�a�թ�W.j&���͖�;�=���њ�{SUk�ۚ�Ϭem4����V���u�w�4���������p�.���p�O��91<�ٵ6����x��d�'w���yu���w����;�4���6�BP���6O%�b���䚎C�5}�CS�rMG����r�(<��ܞA�Ϲ�02Ӷ�����o��\��UB�6>�G��t�r}��bKC����?oF���?K���{WW���t�r7�m~�:~�I��>���	A��Ǉ�h����͎֥�J���rl���#/5Ws�;����pd>��w{��5��'P�I�q�h��[�pdw����5'��pu	k9/}s�?O���>�iy9=˓���s��}{��`c��O�����ߢ$G�}�D}�s��}�d�֮�p:�GP��w���������(��{9j����}}W��5fkC��1u������%>˟y͏�u	u�=�}��0 �ջp܋��3��O����#��ޟ��r^Z�$�>採���Q�y�5�˸��'Q��&N篰7�]_F�:�NK�������!(4k���|�5�ߚ�n~�d�r-u���]J�ݩ���2�u)���� ��1�Lp��v��J������K�\ӿ02�r]~�6��K���g%��d�rMu�d:����n]Z��5w�:�p_Z��a�)�r��}�o��z9�v�g�p��r}"G�c�#�>����r5���i� ���5��Q�JA׿{�����;y�n`�yGf��7��j5r?g�N�?FI���;���ݸw}�e��>���rwU������s{�s�`��	w�A����K�o�%�rw.]�' �qN��}����P�}͇[�2y|߻�:�ơ+��NGRj��ל���#�y���.�w���Go��j{k���%����} �p���X�����n� ��u�pj��=�u=˓��ZO���Z�����d?A���y�{;������^����>��ms1~��[��7��kʡ=��)Jz�|_e�5?�����ڸO���J��'��u;�5�����Ԛ�d�ѨJ~�d���?A�J<��w�?A�;}�I��2�{'��tw���\��u��u ����߻��w�oÚ���ۓԮ�2��M���5q��B��ў�[�2�}ٗ8��pT9G��D��:�2�����-C &���[.�Eƙ��\\P.�:�� ��lF�k�;y�a��8)B�2�϶^m^�w��n��o1�r�}p��ET�Adͪ5Խ�؉D{��K�]`��u����^Z�IN��<�GQ�7&T�����Aܞ�k�'�9:�� �7	O׽c�z�O�j^�u�u'�2�g|���+��u`��j�B��[1�#�r�C��$����Q��?[�q����%\��5�>��P����N��.C��9%���'^a�~�5��u]�����Ðo�	������\��s
3��7Wz��>�h�Dz&��>�F������@n���~��g�w	s��i�}��K����Bd��.�ÿ����*�c��M�����0��r������j^�O��/}�����߷�.�s�^yמ���A��q3��B����ֺ�/q�0L�&����f//�p~5�s�s0~�3ζ��r�=�5����\�� ��I��x��>�BS�y��Q�`�%��z�y���;�7���;��|���|��9jO���1n`d5�>��bn���N�o%�?A�gZѹs���u��:���_`�3�l:�����y��%%9.]=����Ԝ�*{>�p��A���k��B�ȨS=��A����}|�G����j����?OS����2��2/�Ƅ����kF�e����7&�ۨynOL�]��J����h���K��=�ב��.O��89^��^��W1�7�-���}�쟧�9���9��w�k�����j��'po�'۰�N�ɩ�5/A�:���jM_ON�p�KE�9��K�N��I��}���޴u	N�����*��u�pT�Ϻ�W��"(G� �_iw�pj}��y�%�O�w��:����Z�9�e������Q�HP�A���k�C���乘����F�O��`o0����r��}r�R
`Y�K3��E��#��#�>�u]Gѓ�>�Qï���;��q�k|�j=��5��U<�/d����y��ב�������|����u����\�d�{%FK�p5�}��}������:�3���K/Ѣ!��}���� ��INC��Z�<�cR}&U}�d?������c׸&O�~�������K��Opy:���5�U'pd�}�r�-`���a�ur]@n33&w���{�{�:�\�p�"����M1��g]k �v�b��3����韮3!�&��*�B}6AOCc&�C,J�'
�}�_o\ѱ^���T�%�#��i�Er�C4�����Y�F�Q#a7��u=�UǱE���X�ne3�g!Ej2�<*v���STcp�nxk��%^�Q��:� 5�}/���\���/��/''����;��g1{��ە!C��������g�&G5���5<�I�kIO�>�I!�ʹj�Ԕ��^#��]~��} ��.<�n<��Kx��.��P����q�Jy�'y�����+�z������;�K���]T�}�pFG%��u��\��2�sݯQ����o�Z��ω��Z��}9�B#}"'��p3�;�e�����gZ�)�\�7�.��K��q5����I��x&O���֎C�:���h�N��<�R~�&�y^I����;����@����G�;w<I��B"�>���mz�˨{?k���>̀��kp����\��}��Sܹy�˻RRS�m����jO`��
���~���x&O��u�'�<�������0H���;�su����}���zA������I�=��pn��ￍ�q�亀�}�6u&I�˨yn�擸5	W��s���=���{��g��7?���P�%�r6���?��D�z��k�L���;̩ս���>U!C�����<�?`�����a�Ԛ�cQ��t�r5'�u����}�{�A��B]��:���:��=擸��{�g�~��@ta����5�V,�f⟠ ~hmB�O�>]����Ժ���hё�)�jK��?��ߥ�5Ru��{�K�����Y�y������q����v�����bT�*c��+t��0�T�� l���<�څ���������ĥ����@7}KyC6�^}e��ew^�Y�ת��V�꺅d������-6���VW���>�o�fBYM:|����"EÒ-����������hT���Fp�O�r�HX�Փ[x���xK����es��K�-8�Zb�v�3w�/P�R�MCȮռ�Y�1�E:��.�[�*�h ���S�5�E�"=*�ouH{ ��BLNmU��HfjҪdi��Y�Ãmȹ�꺹V�]��5�t�NՑ|'=�K�X�:�Yٴ���@�����ʡ�~ӑ~a�:��(������� �1�N�PY�վ�[��gS���g�]S0�;�,�2�	�\����!��4��*~�\�����A��3L�5y�.������p�iW�t?^GZ�}M�ƾr��]�w�r4��d��Tիl��2D�f�q|��Ds%�����
������ދv�E��yp�����{(e�X.��ΦNYZ�sך�&bë�X�]i���M���yՁYY<a�������P�~9t�t����u͗�ki]XG�1�Q	��.�~�L��t�u�M~g������*&c���G��ϐ|��e��C�M��^@t�!
R�5҉�l_x>=i��&�ČK�c��h&Ntz�S�C�7Ҹ�ܟ_�ک�y�F�@s���_�L��=2����q×�b	�/�g��+�b*W���/c𬃡i��yp���F3\��xX�ߡ;�:�f�Ƅ�]���W���:��p��.a�����<63�ZL\n�l������b����C�4�.fu��m���.��*���f{n�TV��q�al�gf��.���>x��*�A2�x�R��Ӈ5jpl���h�[�%���T�8S:�������,>l��y��]6�ҷ�%�"3�/���V{�c���ͭ��}�Oww|g��AVlW ?v�2����0Τ ��P�ך �YR���E@��ûCc=S�xR�a��C漡<ϱh]țh~��	z��c;ZŎwOI�9��7p���d�f%��n{��2�E��i�Vgh?f��x�u��h������{|���s���A\A,�j�e����V_ݷQ�^�G�q~�J��1���^�v�����#���b��T$�-u򿆺`�.�')������/d��
S&z�T��裧�Q] � �o���f9F�LP4��_σ�3�zL9�(��⫐��H��[+�\3'ןa�y�P�=�H_%R�m�^^��B#�b$N"��Qz��R[���0�t�;TU��q�R�Z0��{�P	�@w����6F]��]�����6ҥ�)JuÍ��=�󃉺��#<�"F'�?1��A+b���N3�8��ݬ|�^Y]���q��!'I.tCd;��P,Q�u�=��W�cK��o�-�(�HR�u%K�X/yL����#<�3��j!.{�Z�Li�%vi�an�V$���\u)�y��T��D:��s���}���9q�s���:ݧ��s�F����B��A��:P*�k�HnM������uX�T�;#�a�;�-��ʸ��mY�1d6�[�m� �ab+*W����c+�[�q�pb��K�
�eLȆ8	������r��d�6u�s	5ܿE<y�(�"���i����C�<*LW�'fJ��ʧ��{K�C�Ԋ���.��>|,�ܮD�ƆC=/[>�ҷ!��j�#��^˿����)No�~B�9�r�n�ޏ��s3Pۼ����X/<"]v��^a�_�B�]�l��_� �V'9s���tf���Rh>�!k��w}�L>C�5b�<L�����1W5��9���F2�^qe��yт���H��S
L��g"��6��N��u�u�6k�50l����жh�m�y�'y�b0�144{�zỽ��y�놫���b`�u�+m�=u۪\V�u�y˲���(�c ���ڥgFt�;,p6����O2��t����4��ې7��>
2)qq��7f8P<\�S�P]�
��u�0o��;P�7���,��LHZy���Wњ�^���(;}Eg�iC�hOyA�.~R���?��b�����Y�a�M����P6�Ew�墟OK���,�,����G���6�X2�x�-:���_���W�����0Q���A���'y��$�9K6�׹�q��ޤ-��N����ܝ{��]L�Y�8^�+�,ˑT��]d�h��ս�ۺ���0Y�T�N�K3�p|�a��� �[�}�K)V��Sa�l�3���.C%]S�'^�9����3�J]��.��!��r��z�mª�P4OW � �s$N�7�pnfƧ����9q��oMTJ2�q���8��O��sH�$2�1��9:[����� a��AN~g�B3���]\;"%;l��"�.cn`���<p�vΫ��1k��29��l���d��<�hu)�3�a۞mG.��s�gƒ)ߟwV[��&��N�{��r���c̱l2�\���β��E�"=w+�N��ֵr��Wm�9�̓.p��x��s��钰9`kȁ_X�A� ������9ж5��[�ؐ���=ԨB�vZ���q��L�0�W4g�œ��?-4rlv�Z����Y�2�Y|�wY+�e"��
/r�_�;�9�����l���ؿ���˃G=�|;5����j���	�ϡ�eꨏ�8;������+�R��<9��T"gXr���fK��d�
�t-��#b�)��m�+�Dt�G��n�i�Q�E�K-ێ�T���-a�l�Ȕ��M��k��'��m���{�ڍe^����r��Sjo�Vp��2gj�}��r���i\����x��"hצć��i9�������}��:�d��(�k}j)��S:Â��iQz�C��WFK�g�22,��1$�7�S�ZK�
����gN���ʨ>�*�1�Ն���+i�"z�*+7�����&���ɜ&�?=7�š��Zn�'�����������JsԮ;�mX�*;q���C�"E��Χ��u��1�u��mԌ��:vO3PeW��cNy�qW j���M���������@�ON��v��p�����Rǣ���iq���e�KB������ק@p-T;�n��AQ��H���9�9�:>c:�\!pM"���0Ҭ;�Xƾ'R�KC׻`�p���
�����)�V���|j���=v��r4��S���;������5����g�4au;��H��@�ދ:���������M�1O:6&u�nUd��m��&�;���K?O��Fx��	�H�����>Ï	ëN�=����7_<J��;a�(�P��M� ��J0Y����&Vӣ��GuD�{Y� �2�,�I��XR�����Q����'�����[/)H��/�s!m�2�jf��	ʲC��Mn�u�]c���E͝b�!I�I/�mܶ��NKӁS�����ǝ.��@34�}���C����Q��*��z"#�A��=����^n�b�Z5iT95��^L��!`OʩIN�Bj��=y�^Z�F�T��o{T?{�Q������N�?O{�Y�ܞ �M��<�"�%���Uj1m���y����.�!�u�����pv��-��ь�s�&�K�Æ���E�!G��=��J����# t��}bc�
��ZLn�;G��C�/ �lgdN��j����Lfl�5�U��f�&@~�!��^ÔOs_ ��m���퇺��с�q�nu�^�P�ez�zzx�B���D1��R����T�gM��L�}|��� M��e{�*�|��T�t�,vS��D�ת�;C�("y[7�]��uwG��m�p��Ѹ�s�X\K,����}���a\�7\�����	�.�G:;8͎�~ w�}��Kk�ə����I��~]]0n���9L�v��6���x��Jv�`v�Y�)�Z6 ��H;�T|����f5����\폮!�t�?�����@�Yظ�	�+��{&��U�X�KE�PP��7���l�E�N�sN[����ۖ�gX�����^i���1v9�j���q�O�ʝ��򾴀~�C׹��ذ _W&��)�Y�,�U�,3�E���Va�D=�2M�v�r�>�%���F��1+W8.��C���F5�澦MtL��,����4gb����O:;Du]u�
�lj���[ڱ�s
�uzNHy�\ze���S)��jɔ�����n`��ۏ�w&�Gv����ci�Y�p�߆�R.����[w��%B�f�8XI�������8�Xߺ�}a���;��2R=]
�I@SE�Q��67��[�>jT��O�9'��`����zqs$4�5��nMhU�q��O}O:�"���`����4cH�����ZYW��ĵ��HкΚ��"25�̖��	�o"�9S*vA;+ekȻ��\�lb����lʾ��R�zkr־pH(�M�o�CWf�q�#�e�\C812�d6�� ��ڊ�s��y���s�/�$����,��Ls�aO�%����]WMR�J�[��4�s�6����W��WU��o$�."�f^��խM�H����6�W5�b j&8a�z����.Y�x*mh�Yg3*`���yz�l�y���iv�`�G9[�v3�V��TY�/ʹ�E��΄ǧ��k2pN/���i\��o�c{}Hl�̺]2��a���>�V��+�î�iej�����9(y�3N���36�9�;�tÑ^Юh
����l�-;p�y�T�y�D��2��,���+�b�7���T6BAΉ�&���/WH�7���1ZV�� 7�鼺�Q��Kz��$�����\7�6j�����=ك��� hQ��]i�;(1R�A��ʊ�=oJ�s��c>޹�P�R�+p
ɝ�>$I�;L|�ݳWn�"�T��x�"Y�]3�A�	7/4�y���Z$��}@!�N_v�E������"U4��AjF��Y9����;�
N[�z	�ұ�Ѭ��M]\J�	L'[�V�]YVJ�YU�s�^�Uכ�:�n�MD�f�@N���tWE�u���nPN�,-��ee�[���]���X���c�}�~�(D��Ǒe�`b��4+����J�X�e�Dh��&]7��]��Y��!��4GO�n���>����!D���Q�,i����K�i�}4+İ�'��2KÍ�g.�����O��;�bL` [c")�v�*� �qMZbTͭ�D*d���dpm��Yv[ݚ�p-fM�q%Jӡ2]��,Ό
����ɪ�Z�l���cU�G2L{c��N�]�P��*/:�G�����B;|��b4�:F����Z���Q�R�p�/���jxsu��g�跏���i\�݃��ky�N�hʝ�����û}j��)*b�����*��b(����jf��fh�"�`&*$���"�"�"���h*������&*���"(���"*	��jh�f��
%���
��$�j����&i��I&���*��"h(��*
�(��
*��&&h"(��(���hb��j�b
H���&
	�"��
����"������
(����b"�*�H��
�"*(j��f*"�"*j(�@���"�"f"(���h���"���������H��*�** �)������$�*�

*����d�p�RU��t7�5�*?r�cNκ��r�����.�ږs�X�Nف˃~6V�t�s$�A�O=�r]�~�ﾏ�����Ɋ�M~x�;��~�B8Lqd��(	��̎&+*b[�o8H��"�v(�E���:E���-|<��[�b�ٯ(��ؘM��ذ�G2��6�Ù�؝{a>.��C�z���������88��ڨ�u��N$z�i q�&;����*�nG�g��q�En�'��X���9H��D6p���w�_�pA�S$�;9�a�Q{y�u}kZ5t��� �g�TuJ�c�f3A�q˭Ѷ�8C\�%�XNn�y�K�B[�32���	���c%�1�~C�1JL�S��/d�����hz@���ce����r��jVe�e�ꑙ�%��s�W�)gC[kO0t;CkU��8IΣps7k"���{��K���"��`��[�h���ኧ_����3+]�hb^���yҧK{BF�!�h�|���Z�3K"E�����dE�NW���F�������"�ғɃ����-��]m���Z�c���|Ѷ��v�e��Lu,0��z5�fl�ԆΧ7ZU	�����r���u,n�:$��*,�g��E�Ow���9�53���:u��0[�7bZ]7���9�4��)�gX$^<.a"J��LХbSz���9o[<3s~'6�������I.�[�`g.,�\�r���އU�����ﾤ�!'��G����X������8m�Y7�C�U̲rgnW�q�#�Y����WT8��W@�8NN��ѐO�fU�T����Q�F�e���3ù�����q��
�K�V�X�:�6B�T�`w@�0_���O\b�]XY5��owu���ծr��1i�yS���1���n�22�E�3�D���~{���Yn�E<�̥�#!%Xk��2��o�����G\�ǂ$�~���¼p�+f~���������_i~���O���l���g~�!��r����F�*��@4OTGH��q��L�Hw-@sf�-����J��*�Ս�I���,��1�z�#^:�{iPkU�;R��/scW4,^�D>k̅���<`���y9��N�1�ޔ�f,E�V��M��}'-�V�4Osޣ��|PrFEe���T�>�֪�9���ܺ�B
V+�T�=j5����ɌD�
��T��bиgI����oȉ��2����o1���(��Ry��0�)�ڐ���m+������̽���nθ>��������Z�R���O� �=d:�86���J������=���N�W���1�y��FDk������*KQ��2���	�{�S2�J�	���v1u}�}e��l>\�,����S�|��K�偯}`JuD�qD�|���/**"WV[�*;�J�Tf�s�W1aNuB������\� �Br�����^Y�O:�.�g=�cy�es+ܥ�S(�5ɚ�����
�e6;d4m՛Ϻ]�؀���}��l=3�SM�'o+�]���8B��v2~��Q���@�;�Ѯ_*����x�u=w��)�R��n�ԥ�����X6k�PV��\�W�|/O��� ��!��T12�����
,�2�a���;���n��[:,� �5��+�x/���%Hla�\�cv.�h����{��ї�����{�i��aWn;:��
M�f�ׂݶ=k�td���b�Der������mP���2E��Ψy^��h��Um}u�Ո�p��&���!I�ej]|_݂���a5=��ON}��^;��\D�LnNV��D��w֕t�7�lfò�L�V���H�
�PBD��-.9�gE����mƉ�����Q^}n��Bsq��-|nV�2��e��j�U��#z��E\�tz�;�-�_�_��.�f�� _�S����o��'Ğc�X���reN�$�i�簣�kQ��&��pE��̶�79vά�]5��C��(�Cf�\�M��\�~ɝ�
�}}���	
��<�Yg��6�@���_�T�묎������_9c���!�ʊºG;�h�T�.��<pq�V.c�^�/����������Z�z-�p��φ����S�k63��%W����Bu�I�wKK:��F}1��k�u`ɖtdQeK�����ʚ���ڝ�3:T�j��I�C!ˤLXc&�7Z��e6G�����Dtb�T���꾐��d�]���>w�Ѩ��*�&�u����8XB��T��t�~͑�M���p�O#�d`��Y�P'�A��n7�q��_֚�"�d�MM���lbT�CFگP6�G�����$�2�F^��!�u�����pv���u\a}�~d��UY�H��3#�r�����w�PVf��:E�.���_xv�T\X�^u�|
�r�ꙸ�ȫ��A�I<9N�W���|+���sJ�|�JJ�B�E�^r�m���d0kӔ�4pA���g8CO �a��z3���vW���4��y�šw"i��G��U�v�L�����䢧߆�p�{�_�`z;������-
&Ƀ�QEW��Ok�j��2:�ϒs;�N7��,� ���X�� �,A�y[Po�ۋ'f-��:�\�rM�.�c����
����fm�Y�ュ>�{q��Ǧ�W8�gS�>�J��ﾪ�3y��RE��gFKS��U����w^���O^�M���֧���9*�&�!��%���wr;]Wik�K�ŖQfUF�:�;�1����JGYZ�_� ��f��Um�Y2�O�b�8ݮP���#�&�:<�	h�O[�U}q�i��_(�,��xn�ʘ��:��:5�3�Q��L�w��-���h9Nk�8�![U�L�ݙR�Ҙ�is�>a��:`v����O+���	�;Pڸ}��=xv�M�8�]ә���$ۤ�˥�P]���ײ3�8�!�[��w��T��,��-r0�*U
(�s��{�U2='���yJ��J��mn��c���? �Z��;���v!:C��j�1���$b|@��o��MkE&Y��ʹ�9��8;������`O�Ʊq��r�EΈl����� ���GMC��ҙ��/Cɣ�'Y*�� a��+�W��3p7����u�7�s!�.q��ͮ� iE�4�)�HW�Đ���M{�C�J*�A�f��+N�2s¤��kj�(����{�\�nxd����j�52w56�{���m��j0�3�G�y��5�(V���E����/*�r�TZ��]+� -��fV�uoYR���h��>|�ޫ��ʈ5�e��Y�x˭7�NS��p���֢V�l�2N��j0nT�p�ǽ�������w���o��#��Lײϰ�k�Ahd3��ǜ�j��r�0p�B��<2z����h��iO�=l��Br��P������i瀆�+������P.y��օ�q�@��ɓu����ݪ�P���LE��A�Y���Qĉ�wR"�
'*��;�D��}=!M���)2��/����/:[7�}l@��Cu�F�Uy�k�4B�~_���h��q�Ny�*m���T�1QI84�b�2l��W2��C��}���q��W㽡��e���f�rp�(\�lmS�� Ҡ���`+��EG)�X;m�S�<��';�P>���+� C��� �B$�#v�V|5Յ3����S����\��O�8�p���3�N�>�3�b�eJ4 ܃�e�z�/)�XcE[ܼ~���[���j�F�n�k�]�c�����GE�+�$�k�S��ɬ�+�5.�:�7�I���%���|�Sßs��m�s2�W��@�t�U���©]�ڽ�5��x`x���M��@,+�Il�e�\6�7G^�9ǖ=��Q�,s�n�]` ;�wS۽H�� ��}x�qRS:S2w,��9օ���cu��r�tV�xg��jΫ�-͏u���x"�̋��������jg��bj�D}������Y�"[g���}&��cDV��U���o�M\M�g��Sv���ڶ�Dn�GZ��E�|��A6&W��@����
���괩�A�4�ڴl�^~���4{�Lx7˥��{YN�Լ�P�g���_F5G{���P�_�����ǙA43�RZ{�����E�Bey}YQGI��	Wz�.�N���]ܮ17ӒhE����*D��|9�v�O�M\�!����S%�,hW��PDO'6;��*�l_��.��u�OJ�\�����d�͸B+�O-�MUɼ, �',/ʱ��#�����9\�e);gne=w�J/�sc.�n��n_�F0/�g$�V�\�Npm���o-^��Hb����,��y΋1�+�~�+%�{�\�^ɍ��o�s��<1���2��ܕ��O��J�yf�5��w\p�����id�TA��'����|'�'/���d11�K��T��J���	�Ӻo����6�pQ�=�i���3QU�W����xn��N]L���^!�.��V�!�z������@����/)'t�m֮�u�U�+��P�G����5�L`p�9t6+�&�=�t�n8���m^�϶���r��$s�vfI���0�Μz�J����R�ܩ��p���g��S�Ni��3�lo7�ƿUW�}G���Jŉ =��ӯ�uI���͎A۪קHp�C>W�;���\�^C��=�+�I�R���}q��EE������U����n��۩��8K�%��G��_{r��2��'#Lp(��w>�����;��_��1��Gs��NT^�#���Ka:ܲcF�N9�wL,�F�s��e�P�[�s���~ceoS	_Obڲ��kc�	l~�q��K�G�� ����΂���Uk9M�Ɯ�� 1��k�C3Њlg,޴d\�;O�CNQ�����I��!��2lfy��
xETќ l�0H����i^�'\�(js�OF7ptؖ~B*��x�����!��¤�f��9�ذ��Q��5\��T�*x�a���7Z�Q:`�@��5"^�
����M��1���C�ݧF��՟r��֌��%P��n��� p���*�I�EU���'4:GV�v���"��?I{X*��Ѹޕ��'���j���2h��v���ˤ|1&J�c�4= �����] ��
��$iQ�üԘ���Y�f.ف0'���[��9�eE]��㉯TaN�+��x�z�s�5�����ŘNs$���l�uJ�S��mi��fatl�P)u$z�uٖijǴl���P���6�򪾯�﫱���ַy��7 .M�()s��kв�G�9�Y�������%³���#�g�$��>�>�y�;ƽɠ���Р���n�к���0-|��s/���t}�Q��kc1��3�m���#5�ê&_o��^'1���@�k����Si��5Z:�k��}���{�� �y��e�Fq:�bᩡ�v��n�E�J']��;�Ð�(<ɋ&(�3ß}�QV�E-�{) ����2��^�7������eҨ���<�v�->yed���k|�դ�!be6a$z�ʯp_��v9O2�a���Y|cw3�V�%�VP���4o�uc���D�TO�Z%�o�U�\au7��t7����>�~�Z������k�\������C�)a�x�qu� _�P=o��ϫdWŮ�@���=^����<�X1c�t��m�r�LfA`3����q���>l8�]ל��[m�vx���N7UIB����N��$_ʥ��i�Y��;yW��K�h����{�U�>��L�@���]u��W�l�[�}��/��$>�"��0	��	�YB�6(���I��B�U��AWwl�@{E^�Z˻�P�ɭ�k(�1�d�?,����������K�8��gBŁgw^�i�y{Ȱ:�GO��n�[N���W�U}_WQ����:h�@!2���R��p��p�9O��<4�a�.%�z�F/;�v	h�I��9�:�0F��<�A��+����\k��'I�l�s`�mހ*�_T��&˩qԸf�4 �2K�f�� ����+��߇Jf���er�t[1��F�T�ɫ�j��{�4�a� ����hiE*�_Þ���;M_�ܦ��S��U��ь�ښ���P���P�7z��H%�y3_6���� �41���tceuF�/r�n'$䃌22�+\0��}U��	;���e�N�S��f��NY����q��Ο�T�1k���k�SԺˈW:#�z����VX�J�����4���a����D^NFp�sJ+���t��پ�����yԷ�Ce��.3�3�]L(<S6�|Ѹj�'n#�^��Fi�s������K�3cW��@j#K��XYW�'�9uW��k�����LH�sE\]�Ds�']��ձ��S�;l�Ol�QA�,��\GIoF�� ��چ"c�N�j(����ʫ2�`ʎ=ꝱ���c*�{��(�UI�HY��<��Pn�6����c�1������\|K�`l��"Ռ�P���ݦ�M��[%�b����}�["�gh�+��,����@g#�]LN%5k� ���"@���6�2�$\v$q(����B�����+2�����:S'we�Zn\�J�����H��[�Ю��/�빍����Q�Wq�+[ؕ�w`��GE:�c*X��.
��״Y&2jl�:�]K�u�d����i>,>EV�"���Jkm_�{����A��\�R��G'fPuS�
Y)q҅���I!J��-�u0۬��5��s6�G��rss2U�p�[�Ѧr��3S���Ґ�х��i����S�iM4���Ή�ƺ�]��p�l�BN�u�qu,mh�+(��e7Ě��p*����,ՠ���!��$Ѧ���}P�)L|㬼L�_h���cW�b�=�
_CcM^t秥���1�$���=u&�uf!ŶQ��5Q�1�%��{]�.��qi�����e�S��^�4��(ʌ�6�gl����&��F�ug1h#D\J���QL쏖��E`v��-f-�k���vuɪ�{��p�7>#���}9S��zm\��8�3�5YsY����ZR�MwU�I;jw_m��I�x�'9�j��t��V�����ԏ �t�G�z���@�Ɍ�k/�*wfG.�0���m;�ӫ"��]+��ŎJٯ��QG��d����q�>&��2��ѝkw)�zI�-/Kuuk��I6UÀjݙ����W:�tt�F�����MJnoy^�h����Sw(w��6	7]�'p��֡������F��t��\�ub�Q�镶U��Pt�5�f1�W��j�p7�
��ԩ��ztv�V��vk��Rǁ�q���f�٣Uo8R��X�e��_+��#qc��m�y@�+����cD��nn'�e��s5�lj"i�#Տo�4Vۥ�u��S��m����9E"2Psq(�ڼ�j��%N�<�{]w��q�+���3oV�6���¼}�S�E�4����u ���T��Ț=ւ� +��Z�02�TrLW�ca��Jz���w���@��V�쮁�@O1G��Q����̾�{J�5h�
����3M�Rf���&e�w�W`E�X�������:�h�v�&���rVg�W]�dnVҮs���R�Љ�l	����u�;^��C%����-�+����N�\Ս�ë̬�A�w��6я��`WJ���Y���f�w�K�h����<�`��#,
�xOq�%��א�������CJ1}�F�+-�ԫ�mu�i�X!���iCZ\a����c ���P������#D�4���<3���6hk)O��;��2�m_a�VU9W/{� ��6J�c.Ĭ_��UTETSQ4DAP��Q�AQTMS5D�U!�5KMP�DCTSCAPUU,M1#TTQR�TEQ5MU	HD�U�ET�DKM4�-M	LMD�@DSKEP�QDBQ�P�SLCATRP�IUMU	QP̕E-PP��1)U4�ST5DL@�MC1@P@QIQ%R%SUM"QJP��L$DDQ,M)E$�TP�%P�4�@�T�SIE%4@UU$�AR��Q@P�1D��D1EM4�AP4T�U%4�����ee����3�U��+�m(��Z�'�it�5���f�Z�դ*t�����{u���-X�Uڤ���>��K��
�{��n�ϋ�[�_��`�t*
�2��@�0Xh�S���\�����U��_]�d.��qj1�r��u��0�ܔ��4��֏obו��ڛ(���;*X�?"�P��9�ё�&ˈ�@=�n�znnttQ<x"J�B���ƭT���=W�p��Q�К�P���D)T��!�Ŏ�zn�HۅO�ړ����7*�W����œ|@�Ė3E鄊[43�E&�&��=�!^��w��_+�~�bk|݅�	SR����3�r~)�@�_uǝ(�T�2��f���;l�d�[�<M���pn��u�0EG'Pr�S2D��#�ʡ���=�Ls��3�^��.&EkW�4��(��<�5�}��o�\�d⁫Ce�<ɵl2�Zt�:�B��;�����4����/ӊ�%�L=j�0�ꟹ�d��5௬SΈ���&�xqhvI��)���Q�5r��ۘ�{�EF���&���F B����eX����"&=��J���G�ĩ������iV���G1&��M]/���Y��]�j�U־:E	;��U)O4;wlwU΂b��ŤJ56�[��8VڅE�lq\V�ɸ ������w:
󶕚��΄;ެ4�����r*�Xz���,|�l�*y������Qm�����ߙ�N��ߌ-��Y�{���)�a]s��$��:Ӝg�Ϊ�p��W6]���x�>�y��컏�Z+E�w�_�_ܭ����s;�}��^�Z��Ց�Bz�K��'��\'�%B*gX?p�aLBk����k��\|N_k�t��2�gX��O�-�ֹF����,�9��c6}�4ҩ��@H�����0++	�7B)�g��\�[�_-�1�LDv+L�Ȥ��/�T�숥_n���g�zq���C>V���<"l��7í��,T��j�K;�����7:����s���tM���R3\_ՕE�u�Ћ��֞�E�2:�atzjc�֘`��UB���ϴ����p������d�ddr
'�pj���OP6M*�']% _	Υ��xeKTY�X�4�[�̆^�ݑ<6��mΝq�@����Z<K�<r���`tϋ8S��魈�:9yT۸э*ڑz+P�֔�	r�mda������
��F]D�T|�T�M$:Թ�ҷ��mU	p�������R%�ގ��������%=����շ���&zzz��#Wݴ�gJ����G����`)�C��|��Ix!����g�ke_s��������B�#�"���@�^�S����6rE��S �j�p��$j�r�}�����:�b��f����Щ��w��w��q7��7�	g�(CW$t�����7=����o�ej��Q}s-ϑ��z��P�V�9t����M|��Ө��0Y�}VL{�\=��ݜͽIM}(�$9�]F�R=\��kF�/����-@t�,A`\�\�gOM�<}RrI�(U܁P��3�Us���s:U�辸MT��MZ��#�v`n(���Y�`G���zi�t׎�g�e9+�~R��4,=�.��f��`�I9v*�w��������O%���;�7��<(�joX#�^Á�Ǥ�aP�y���MP�������C$���>��N���_Q0���W������6k���4�I)��T/%�S�6�|�b�'/:�Qz��FY�g!:�b��m����/#���7X4�O-���x��f9J~D��
�̶Od��ع䌈�0�7~��q�p����Y��a�n�E\���I�%ڲLHDط3�G�p�9;3�Jf�%��ϲ��6nOO#������{%/\�����aga�Ṝ&�@"ﻳ*1�-� �XG+����t�$�x�c�}��z4������VWT�si�in��U#�kik6Q��7��#O� �nQ&�Y7x�庹��H�2�ڙ������\09���^k�V*��FM0Lډ��TDDG�9�r_G7˄Vl�
�Rlz"ܒh�Z"Լ�o\as|��C|�0���W��S��//g� �}���6��}r4ذ�c�C���u�9�F��S=w2���k����;Zq��Q@���c��T:C3��gi�p�>3��P�
���O2�
���_g:�Q�\�=�9��WO��n�]/�R9v����ւ�s�]D/��4Y��rs����jn����`�Ȁ_7�����-}qN]G��S㺝!��=�#*R���X�(frF%�_5�fx 4À��)�t�����_RN�8\������H;w2`,`~ȶ�1�v�r�a7� �%�_i,�3����;uxz������x��kĄ�主J�P� �Nq*�ʙ��F�E*�X�����;M_��i^j=�7P�&�Ÿ�rĲB}<*L4�=�F���.��v@������P�m������~F�z�������R�N6�]������q��Br��U^���e���k��j����|&qV����"8�E�m91�õN�|.K�`t��md�׻�9�J��	�fVK�1�j4�L���T�y�¾[!�ՕD8����Ẻ0V^����\jU�]K;H�ƽ�DF
���˛���ΉJcd�ͦ����{���G+W|_Vt*��'��bdw[.0�/䪘�Z�3K!�X:i��1��DMC�_g_OX�o[������x����Δ]��ALI��/6��ȓ!�ϛ��-T��gH�jp��riE�������z`���� *!�	UDY$,�4�-3/NvKu3lFq�Չtg��KW�Cj̕;e���}LL�F��˕W|"�j��8!\���Q�`,G�d��U8�6�Lq��/�Ί��(R��k�nڬ������+�t�b��c�b��}R���'�48����
����gTS�����O���7Vh
�T~�7ۨK��&>HG�I>�/%�끳�*���vn�dk��3���鹹��.O�2�כhCUؗ���ĝ�a#_F�r+>]w͊{?T)T��!�Ŏ�zo�R6��|���'��SN
b�4��/��P,�b H��]���ˌ�pg{�gP�	��^�Ų9=v����.y>S[ZS��Y}4��B�G@{%�)W´�e��=���sw)ձ��F�즜��v�B�B� �ɦՙ��]Բ�ʦ\�KU�I�lR�S~�z}ň���>�Y+�h�y�;iMP�Fes�\I�BGdfok�-�����2�B@�!B	�Z9V���r�T����ײk��h��$�ۿϾ���;����:�z �E���`�S�ts�x��2+����D${ܘ��P��g^� �EIi��.����>چ��C�e��c*�:�%J��(���<�&���E���\U�֭���%�F\�17��z��b�>�����KϠ9`kυ}`JuD����5�g6��c3�i�=}&���h�{�c~k+��n�����\��Rr���ʰ�J����Ee�5�G��sd��NAɱҧp���P�Ɗ���
�wzqs�9�O� �k�N���Br�����]�U�r�?�xV���_ܪ������t�F��{iW� �e*��/9x�wq�W2����Y���l�D����}�B�=�����Z6�&�e$����t�z���\1���{!���Ӝc�T鿑�3(�!��J�$͡��ܩfq�U�x\t�1�Lv;�lE���~K�vR��at�
dW��<KD�"]����g7C���G�?�B/'+U �@�v>�-�*-�7=�򘎷F_��؏���XO���`���B�v4��nUɽ{���i�g�\�J�ܙ��VXŐo�ȳ�Od��Y�X$��+6��ҟe))�=]{}��u�Z�uwB��o�S�-��̫���W�,9\ʬo7�+kEb���)�5y+�!���ט�A�������{����k�N\�}��XG��Ck��6���L Q����s��i����¬y�҉�iƵ���H`~�^�4���&�	:Ҁ!�u/��k�%�>5�Bir�ř�������)*�lY�/�~���&�P(9$��˼V�!��#{��_{dl��|bW�l����%��;�i��c�f��0� ;���
�������#���tU8.R���J�:!�u�F|���<�Cr��n#�:`��B0�Jf���Q���Ty��շ��i��~�����i&��2�;��yYǃ�(��,�ܛ���B�Jp��7Իf�y:�Z9P�9���^�R"�g^R*�z5�S�a%�Ѳ*��?A[�Qu�f�ymB��5D��I��'P��n�4K���a]W���:E���OfTe-sq��-M==�,)��ݮR����؜2�3��Uk�u�H��N__��ޅ�k�`;���SFvi����u/�l}B�,�P.����Y�Q��VKH_ q^���#���#��m�����9���)���$���)����}�]ݩ7[,�o^Gx8���!������w���?��'FcY��j3�	���R��ﾯ�y�M\�\�U��F���ڷp����c��GUq�fTpB��ڡ:���Wo;\	�y�&��2�O���v��x��񹙜
�m����/��YW�&� �;c
�����ғb�ս�k��WXA� ��肵F�}|�쪤P7�i��k�k����˛�!F-���mʗ���Z��{�󾘽��L���T�KW��r�uS|��:��Ì9���b�{I�Αj[m>���ٽ��Q�}��:g&x�z��ox�՚�J�n�N�y�ᬼp������Q#��0Tm��s�����P��)��u�zSW��.�[�JS��vk��|/T��Jo���ܘ�q-�����ދ�Қ̀�����/��}��h���c7��k�h��;[c�̖�s�送����+�`[Ջ�RM(w��w9���a�͛�rÔ��,��í��K��=	��*A]W����+�����
�Ν1�vGJc��ou��@>�Ցe��5P��W6 �?f����E3���O*�E��绰d��W\�H5�DB����V;���ں�+���r��}�@m�9����u��7)�\0	�AH�h4g�>s�pt���ȵ	�Z6�>v1>�[J�l+w�WJ(J��P=��&�u�ڴ�	x�;,��ܠ%ө�ҩ���䘚mƸU������3~D\��W���',I�'��g5�}�դ�j8sP����V�#5����%���z�)�K���.ֻ�L^�J̮�������ԥ���U����t�F�x)�[v���N�q�m�ȽQv�m�D�Q��^�;*^#��z�'�Eb��,�f53'�A��.ʝ�#={�ye��8�Oד�ţ�>S�ѩr�:��㹜�:�ڛ:�:l�B�{����9�]�AW0�m:����vfQ����'bU�f��QO��sa:OmWnھ���ĸ{G*���חP�NwI�G�<���Q��j�p1�Q�����O4ϣB�n����5�����k��om��+u�n�+�c�+�W#j��)�;�k.����F_
m�H�w*���
�3/r���3zw����o2	}��-\B!�s�Z�Y�wv�w�S�lEj����Y�>d����������a�-@B�G��*�a�����DNN��벪R�p9��Z�[O8��N�OfӌHV�YI��hc�Ip`w=���t]C��JSˎp�㇆6�T\0��L�ؔ�mKؐ��|W�&+�)+���S����Q/L�[Ө"���S�6�ˣ6�1����]�vA`�KEiMd,�M�+::�C�=��`u�D����jy�5,�<�P��9��R����ӝ�)�HQ�K�)�j��5ֹ�"���˚�e�w�
ø�(�v��6`�F�C���͜b��Imqf��]>ٸ�n���!����&���a\'$I�͚�i��f�kG;#�5��W%�fKy9�ڞ�Ԟ���Bn5����Lcx�:�s.�����̪��ިsۧO?M��L�*��nՌ[�>�ߠ�{��skmȌ��%������P��[�U��c�g{���1y`֢�����SLX�����.f����A��^:ޢ�HA�����J�cMg_P�f���8��l�z�)T�\�}�bٓ�r���Mgp��+�-l�Ӎ�Xqs��Zݙ��i���|q=D�t��u
f�!�sЉk��n<gI�[u���l�X��:�;8��޻pγ)�����fU�;Q��E�R|��j��TY���H���64�����k��׭��d�$����Ye[���pʖ�=ωW���n(O=�s��˹r�MJZQ�5.�o�V�y�z�ݔۨ,�v���b��E� �q��I$���2m<i���mYl���H<0#�d�L@Nڃ�R43��X��cpނ��n��{�+��me!W7Q셱�6��1��D���_Z}�H��w:��*!M�&Q#�������V�o&�3>4��%egd�`,��-�$7å<�)�TD��B��wP�u� w�wPd���-d��cɘG�&ݡv��M�q�<ąp̫��3jpҰ��aLD�HE
�@�u(�4N�un�s���{}/ �"J����8�t�K��Q�ݤ��0eN[�7���U���¹3{zR��ћ��+�!�B�Q8�J&>T�y�U�ڬ�H>L�Z�>=I����#�S졻�[S�b���u�s�X�.�kE8�8�#$��~59�&��F1�yU�Pqﮔ���	d�2�MC[�š��tec�N�c���#�1L=@�[�Dt�d�t�F�SOU�����0�A����tn����Qr:x_r�r��������ӆ��SB5Y��Z�^s�'W��91fԗr-WN�M܀�UUв��K&���'��P��}��-�`)+
�e��)���Mחj�l����7�Ez�i�3������a�l�޲i#٥3�G�hC"�M;�&��A�b��KT��Ac���5�6B���#r��;�r��u>�)��#@b�F�Qc4�S���[��Enl=s����rM��6U֑zb���Vݱn>j�����|���R�2�r�{�Iݕ�mipi�;Nj����{�����{lu��f��ۣ�*iא>W����iG���9)ҩ����`+��HWc1�|Z�d�L�Ճ/*'\��C�_N�Y�/��%onk�u7]ze��l��J�.�%���>J�؎�ʉ����I,���b*u[��2�r�D6���-��-<�2���6��8n��wnH���xf�,�t�:����N��)D�J�b�B������Ѽ�I"�(A��9+�\t�*�E�n�ʍ���+� :�
�����I��3���kiF�Kt݌�ރi<I���� �{�wV���Y-�-��t
��dP��n�i��vI9�ҟ�nt��Ty�)�Q�بۜ����pwȍ��nb�:ď��i��^L��.[���y��T�r)�e�����(��wכ:�GYk��h��b
*��i

"i(
����JH��"����(JH��H�h
Zij�Z"�
Z����J)(i(B%�������!"(���(B�������������hbJ"E��Z
�h
j����h)�(

"*�
R�)@��(()�(i*���(B���jb������h�"T��
J
J���j���H��&�"F��)bhj����R����"�JR�(������H�
)
wu��מ���o��m����>��0�ݤ�n݇�e.�\nQ�=��;)�;5gr{���6�Q��U�q>TW)`��я0wXХ\��ĥ%���{i8�>}Gj2���3��I���t[�r#u����d���WX�ڙ��K���f�F��[���!�PU��or�LVO�d�R4�|糱��Rm�?���\{޵��k:6��yI���w0�Z+]�i���=(�Z�{^�sQ�����[��!�}n��fu�NGwl��_!�mR�YUH��`U�Թ�PV�T� kyq��9y�M^E����J�:��!Ƕu�����o>*ʾڔ�D+��:���f�_jr�W����ӎ#�7��վ[pi*����ʌ����L��9c�iP�s�Y8rؔ�K�/���vF�ͯ���R���p`G;��]A@]X�彃��`{��'��I��!=�Qm����(�\�goH)�㘜v���8���Ǟ�}���B:�1q��&��/����wL�h�{�FD�����E�0��r��ޥY;(#QG9W��A��}a6;c;	91�X���i�?\7�K�ޢ���N7+���G`V��E˩܃���|NN届ֻm�̠��eYb}ه�j��;Ӄ7Y[]�s�ͫ.A4��YS�<��Qط��i0�	�Q�����u�<�}8���o�qs�=��o
ѵ5�wB������W(J���T��u��7��{U����s֤����f�̃�m����6��n5�WU��:`Z�t�]��K\�Sܗ�crU��q�$i8�W��bp�x��'�_k�u�L]_� ���6�n�i����?s��GV�m��T^��]��uS�Y��5UGw�e��$Sm����]#D�����c5����m��ՕX�ڙx�D'�\5[���b�\
�5��K}Ǝo�z�w#g2�:1GZ�_ʹ�q��鉼�˞�A8]!��O��4�^Q27h��#�}a�L��ίt�k�Q���ң{�r�E�3q�٩�֟9�͇}7�r���[;,�+b��}�TO^[�	��b��7�	��=�j�yQ�3�ގ���vi��Z.[<G�����H�9��Q�Ů������m0c�P,���3t��Pl�|�J,طD�MN��TTDٛy�}��Q�*�F୛�l�,�ާ�u�2���C�����H,�A�� "��'J���g�ĹOJ��ͮ7��<�8��a;ݥ9_+#i�������U5�����Yc���z)�:~�t���8:��J�a���F���uޚR�\G=k�5�mE��X&��O�Mw�.}@��� �KFƞk!g,{-��b�gB}�s[�w+��{�z1��(s�iGJ3�t��C-�s�Y�b�4���!�6f�p�Pu^����v$�+�l�"W�R���S鮥۱ɪ��]�ϻ��"�Ӂ�sZ�8]�i7��xð�%J&~�Cdu�`��<�8�0������Q��i���[Z�t�T�ܓQ��a\k�/�فs}������|�)Ųr��߲��W�jU�I���jpv�ʨ�dG4^�B��=-uN�ڦ�SjM��*#�k��{Q�X�)}-p�=���a[�)�Z12��d��=3}�A��ϭo!'��=�oy<[��ω�k�+V�HK��xK�)� <�]b�AOl�H������YSi�٘򣢱��[±��G�f�7��f��6�j<��F��nP���l��mE4ż�`[u#�$k���(JA�SؖW#3$ltC�D�ta�t	�[ԳD��b#��q�t�糈n��띠��l�^rF��c2����Q79P'�;�8��\gj�b�r��;���g[�rkw��׈��J|9e������({�,�Ŭ=�nL$�>�����͇)��J�b��:p{�~]̸;}R��	��~ués]J������DZ���M>��<��<�ߠ𣓗���K�7���烹�V�N�u�U�JT�sy����iꟌpX�^�٬����މ	�����^Ԥ�]N��}
Sˎp֎�R��c�jW�E3����)+�8�>�l�|�J�&4$�嵽q)���֬��ﺏf�֔�N0��N/:�P��EU�w#�L�4OK�Π:�:Ss׮9�WZ;i�\��RҰ�RϠ<�P����_T"s
GCF�`���\�.gJ�H��q�˵�h��5p����<�,��E��^e���2���1����ۘzMl�&�n��z�x:�9:�u��G��8�F�a��"���-#s��s[�����gY���)Gٖ�;����(��m���w:��3�V�|�wDnoS�*��`�Ѵ\ޝM,4;s��H���tS!N�!s�Y޶�t��������އD�v�w�V��&v�䣇^WB]TC|6lua[�y\�oun���Tic���k�bGP�J���?P�Ku�u]�*�s5z�����?9RsOoe0�ӽN(˦7�:I�w)c�J�{gj�[�Z���W�N/�o���5�:�}��P�� s��|�3M9��t���[�If��c0��eZ��y�R����B{Wd]r|���c;z;����L�c%����U�.������OW����_�����|���79QT>��k-Rl\C���v�ל
�9$�!�R��]�S�1P5�m:��uBW]+�ب���|�Py��i΍�YR�VIzť�v�4�ݶq@7(�@�u�y=r�H��p!��s��VW#3[�����&�_Γ��+.)�o}���s��ȏpz1�S�������0"� a�:T�(���,͠��ED쿕=je�Ajwtv�H��z)�5E������Y�#އ��q�{��M��c�Ԓrwv��98!�Ѽ�󡼷�c�۝$}/X���yC(�C��754ðv�`Z�� GlN���f����ճ�3g�b0f�.�R�{����[�R�C��}0W����N�R�Ԯ�,�ڙ�iFe����*}5_e�=k�5�mE�2�����.n]D�d�`���������;�V�2���:��ެ�=�Qm��,��sٱ6�v�iܥ�5kV�ڦ
[5K��B:��\u&�e�w�-����#�����t����3x�} �P�`�s]K�o���5��s���vsr�jлͩ.��:�]	t�(FT�y���C|�4g�*�9���[ґ�@�q�k�J}�F�x���cப5��`�����Ν�A(�Ƨ3ZN�΅�s\�&��Kj>�V�9:�N��8:�κ5��H�ӎ ���("��ƻGo�qQ{�~�Uv־�����5���k��s1���)���Җ��N���U��6�c��{B^��X�ڙx�|�5mV�uX����^�����i�{뱲ӻ�6�d�4&%{��]��H�;d��k��N�6`�X��<i��1N�5�i�S1�]{t���bRsn�pi��5+�-��;���<)on����i[l(��Fnp�ԕN����O�թ��Chv1�ا���u�f3-P�+X����{3p��/�y���j���p�pu�N�������b/l�E0�*���k�N������N����Y�-0��<�7��������6��(��z������t���R��d+�;vd�Ys[j��kb��7��i�Ĵ����ѡ	뷃��o�v�y�6?l��X�K�UEl*U+�΍p�_���|�{pm��C�,>s��w����:���0��:9.�mRޚ�R�_=k��q�V�d)�3Gb �V�l�<'\
s椨!-���z�k�/����T��UQ.n�n�R�۝���fQ
{䡀��ҹ�,�\s8�7'\�u�1�:��p&������3�!u@���r�;2e���:���2�����p��9��q��+�R��7 uC^K'���}���Y2T���d��L� �	^N^(L���Z�گ"�G�.�Ļ���g��;�@�meCw��*��Ch����E&�=cuG��	Z�k
�Z�m�O�yÁ�ç$w����6¼��jЧ��\NS���������˹�!��fueM��]��엕�f�;��je�}SQ�15ۍp�3]?rH�r�����*�E���:��e���y2T�r��<ӥ���浕;gl8�c�j݀�q�����d�����U�:V�ﻞ�M�J_Km�rҪTL� 8{�K�W6j��5ù��x��Q��m�D	X2󓽞le��[��ѩ���-Z�һ8j�~R}�����H���ӕ���{�i(z+I[z �ԓ��\1�k�ne61֮��t��/!�z�OÖU�٫�u?r���ul%�/�_�\r���:�خ\ظt����W״rPz�M�w�P�k��p
u�;5�Е��J�6*�7��z/�^�8�:i�x�]�c���`0uLʢvx��+e*W����5����v����9괳�%ǭ��� ;>*���)%R[t�j���n*��[��o,^PR��q]f9��f��(�wɎ���G�ȫ�֫%���̻[J��XL�Vhd���t�qlݻgx��s
}M�Nۍ+Z�2d�vC�sfݎ�"�U*�vbp�ѨCs:ZߗT��r��T����Fh����3�@H3�����/n\�X̈́s�j����l�7����/��r�2����)+�����S��;<sP|4˼XZ)iq-�����Bq�Qm��r�����X1�KA��櫾����7�s)�1WK\�X��Դ�<Գ��BleC�`���yP̥ϫy�<��x<w<�c��n��ڄ��������
��s_f�)Yj�.��c�ϦJ���;��ME���ִ]|�T�rL;��c4��=���Ho}�v�?�Q�mrV�_�g�&���y�W{���{_�<�v��ܩ���ث�6^�ƸU:�cT[_����_e-}��^�r�ĝ��hfF��g%*S�][k\9Wl�CyU��Dk?@��3}6�(�[%�b��X&λ�=��OZU���������w+3��f�5��b9ח�عP<k7I��Wܜ�ځ;�.;TLV>v�y�^=��cɗO���s#�P���·�Q���>\PW�I{ub��C��;{���BMJ��q�8[���zK��wY\u7�`NG\9�s9έ;ژ�P���3WP��1i�\.=逛z2��A��>�*5�p�7m>��c�p�r�5@�lrG���I�ۘuDM�P��0���̩M��ۉ]��@qݤ��N�I{�K�w�.{��uNs�2�;����l�+OmY�;�&�J��νj]�Y�%9��Q����l���5}G����Z�z��j�}1S|��]�a�w�%�ӯ\7����=�5�B�O܀�*ʣjRz񒚁le+��7[�G�|�T�o7��ۈ�j-����U(t�|�~*���'��щ{�e�t\iM\F:�C��N_g<kq���T9J��5r�J�d#wc�*E5n����oEiMf#�����y�s��E}m��:�Un��'-Bŵe�!�F|�~����Q���B:���i[/�V��;�d6�IT�\�ܬ�{�]H�ȳ� �_��J읭�羇<fըq�Bi{��-I݉m+����q��
�M� �VV�v�ڽ�[ؚC��V�	`�pqq��)���Xl�[/&U�[nQ�	��[���6(挂9]�#���y,��v�Y��ەǮ�|&Q�y���%\��v ����Zyy]���r�*զj��]I�\�{�5���䬠0*��v��M��F�k�#'3UE{S9H+-s��sk�d��K0���`��`��Y:�˩�%c�d���؅KlQ� ��Up�<7q�ATUwr�j���qu�'7i��Ξ�m}��w���B���9NT��*�o��UcQ˔v�E�Z3��1Ų�a�fN�v`%Ɇ�6�!�s�Bw,$h0�
�/��m���D+aj�w��yAc7��{K���������4�p1Z�em,bC����A�7�w�o$��YS	�aKBT�C���<�y3,ᦨ�!Ӹh0"[@JꝻN�.nf����C`��*��ֺٗ�Qi֎C��6����ZBc4���ʾ�ή:b�˓"�	��!��G/��
eT�������\�A��j�|����FbT���-��R�fֱv>g:�@v��,c�p��d�M�ؖ�ʅأ�rJ�%��7wHd���B�A�d�#�k�Q)�po*Ս- `9���b�+�u^�6-�:�/��з��.;�-�Y��3U`ݺ�&��ǅC�.�=�����n��YO �eJ��u�ʲ��ԡ��tu�2�l��*�#8��%�]7*��َP�pg-* iLc��Q�q�u���I�S/*V�r���6y0��=��f�ҖS��|I���1I��w9�v�y�u_7�탕�n3�^%b�7��Y�b��V��uk����Q����ՊĔ߮.h�[Q�W��s��J�Fh�Ǣ�j�V*�#�B�"��[]G��G���&���n,7P�w�́C՚�ؼ���\]�L�o㱎��btVsI��O/����R|��il�3@�(u�S"S�f��³zGm��d�����w�Am�:&�����:B�����m1N�R�(�f��L�Z�^]�GE�4��Ҵ�fN�,>z3���Q�ubT�ٴ%�R���f��Œ#�V��U���+Ul����T��v����	����o�X��H�k�x�U�D&< �ٳ���i���ǰ周]*בM������{���n��٥��@��vi��ok 쐷.ƅ���XW҈���Y���8ڹ��
#���dܷ,�j/�'v8�	M\P$�"Kz ���M��-&7pH���*���Ж���%)�K�Aܳ���,!�2i��uc�H���̱�����z�d�:fU����
p�S�����]�}�%��@�!�X/�oeZ�m���j�;�G|��B�N�p���=���W4����TP/��$���WӒu]�r���a@:����
�;;z��\�Rș
��}Pč	IC@��%P����% �M+B�@R4KIU+@PP��,T%P�A@�4!B�S4,B�)M �PD�#B4�IJR�QM	CLIICIBR�B�*�E	KE	CT�
PҔE!CH@�!T% �@U(SU@R�B��T�#EA@P  RD� R� P�4%%E%%T�T ��4�C@��P�R% }_�T�(�k��b������//۫�����a�(ޥ&���07n�=ݼ+��P4�<�O.�w�{�&�b�cYX;36��=�����+ɸ��"y����Ad�u(��{���{X�o5�j�W�u�pϧ����2�xl�a�y2��^�d���Jb�j%fWRѹ����w�R�k�|��dE�$��G���o�MS�ޚQ~���uFcț{`��Q1������|�nV��1����Bs-oWU�jmY��3(���9�%1�1Gb�9�N��ct����?-�]���j�t���'G��hr���ǝ^����sQ{k�a���q�xT5��D;o��n۾�����5��ֽ�н�o�Ґ���s��.#)�T�R�ب���i��^h'���q}�������^�i�eN�uQ[
�J���Y�t6��h^�nn��
��OE5�1�w � �!���$S���y�������G�Z8SK5=���Mװ��S��T��%ԑ���n����p�Kz�}�����ˑT�u�y�s��6%d���,9fd�n�
1�]��Ot��]0�q�N��� ��s� (�:W�&�;�fV�C���W��*�Z�gz
�gJ�υ�Wg�:c�\PKEi�wB��P��u��e�	���h�U\wm��ʇ(��w�H`�KEi\�>z��rh�����탺�bG�\��y����
m�:�ʄNt����#���~M�u�KCۥ������&����j|�xÿ�����1�lc�g�^�*�4v��x���M�quݳq�kS-��߹&&���+��tE4��po*es�n�}����]�s�e�S{9�:!uZ��J�y7E��B(¶z�s#�.E�[�t�{dL>?{��/2��k����nV;�J_f_�
C��1.hn�*��*b�͠�Y�O�#[״���w�/C�/99��ؙ�Qf&b�C�mR�g����7��q~s}�M�;�~�����DE��mE�AC���˱X�6_.w
e61֮��]�{6��}�fW�]7����������v�xr����5�#�w4��y��A
ub�;"3��Z�j�{H�1�X	 Q����i�]�H6r�1oQ�7��ϡ��K� Z�ڽ��p���CB�շ��:�|���S4F9,'������ٽ\�[E�n�HݼAvU����N�ĨJ�c����S޾�Ǽ���C]Cq�O�Wo�����^� ��Z�ֵ��%��5lZ��O���s+j�t�g_E�ɫ��p_���pUG������l�����p�D����*4�f�*���c6�{�;l���.�r��?tu�I2!]P���3��oM�]�-Ϋj��ܡ��p������_
1�>���I��).�V�(T+�s!vv�Y���W#J_u���>N3k�leC�P���,S7ڃ��26�{}a���zn�󕋻mKJ�<԰<�_&�TC�g�B]0�¹[�=��|���z����\�=�E���6�.i���V�"��ۜ��=I�ʦK��9@�����z��vN�'Z�t�T�G$Ý���r7��J�<T5Or�-�q�$sg@v�>�}���s����Й�w6J�'��<d}%�,j��ș�o���L����+k�8�����MҲ�K<�Ӎ�4
7�؈�C=���z�+ �ٔ0�=29����w��r��ϒ�AZ
*b�լS� ��6�,��Z�w�u�|��	�v/�)6d�Ȱ�����\U�i�Х��]�uZ�c�Z���y�K_c��O�n���'�X�9:ۅ���(�+��U���3�]^�f��%�FܥRn��F���~�����<�3�N�Ovס���
���-JY\����]��W5;��S�_M�P��.#�Ec�Цy�����Y��淵)���Xa-
X^�S�1�_��ܪnr��}�F�.f�T��=͟��q^u���ͭ��Θ����pUpǯ�5����j�VdT�e�}^-���7T�t^��r�E^3�P/*44���y��d�ͥ7�-���r��E]�<��Cyq�>�I�����*��:O%<��"�[Q�ڶ��
�MB����m�8{Qo�٤�P���q`٭�}��Ţ�Y{[f��q�:}4��\sֻ5�k�ob�2!��<�^���Y�E8��<=�;��8�{3��.SJ'f< m�wR��������'N�Aa��`R�^�Uj�m��T���uC�
����[‮*�8�:��6������v�$����R���؈���ݔP�7�$����z���{�Z.4�Y���'��9i\��!=с�RB�LLv���l'����q�t��%(���\�X��O����v*�(
���ca59�ޠ��B�<�t���=,�k���;���B[휍[Z4����س�ܵ#�w9��t=��Tu�BUt���Fn&�k�5�*���:��Wsjw{�5'�&&�7�)��DO!�����zš3jl�T��uЧ[R��Ǖ�e=�׵�����^'��k���vn6l��R����]>��/�����݂j�|�|�����K�Z�Zϵ��v�uK������.ww��8�j�����ő6���e�r��|�.і��쩳��U������l�T�P��^��*�8�)��Jc�(��M\h���ż-s�]~���ּw��nTOCI����>�᯶�I�1�	��e	KTL!�7�n/h�-��g|�
�ό����E
J��ʊ�BqY�\+K{�%���nm5s��_a5
�A���Mk�٨űH�\����fR�u0�{�5]7�vX*5���㥳��7
[y ����r��6p<�i�	����,ɎP�5�lW.os�m����y���K���iF�������0�1�ó\B�R�J��*-�yp�}q-=�{?v��r�j�bFW)i�{�h	��0ڍ��w�eT*U+��p��B���+2��v�[fj��JpJb��@)����;�b9�uޚ�)��ָ�@��{W��ebh^�m;heGKU��dAP`%��O5��B��~��Զ�����U�V��m�{U��&��
\8{ Ϯ��W���1'k��+���.En�槱����&���[��&�)�U��
G�ѫ5��v;%_��|��K��{��M��{˜�Co��xz�T���#����D�u���x��ҋ�R�}��w-�������bk��k�����lY���׳ox��n���Q�,t�Z{�5���W.�=��f�uJm�絛B`�"$q
ܩ�k��r�W�����g�u�>��������"j�=�T�5������T���9I����f���I�پ��HHK�9W���7��䋿N�3
�1[2WC��d�QC�P������7�.ǐ�Zz��D�u�U�ҞTq`���_fJ3�OD�u��6P}�I����_C��~�̽;�3*��5��,t�m�]+qƵU����]�.+����AX/~T�*ٲ"��]��A$�:�_�K�p�.��Ckד������=k"��
�})�T����^18�^��ϡL��:��	���vr���Ӫ|�4.���l����r��X�C�.l9O;�U۶��у�)C���Ļl��1���UmK��P�k�خ���&�l�ȝ���u�m�%���偁5�<�'g�F������˺P�df���;\m�c"�8n�i����A�] �FQ��$h���9s�Ӈ�U\��.��
V҆��=y���Hu�}�_F��wÌ�}Xoz{9�}�E女��|j���<}��fն1�r���f�B�7ð�%ꭧ�a��kP#^��ǲ����)�j�vmN$��TyS+��n<׺fm��t��F5ے�ţ��j��DfS�8�P+̚&��^�ƺ�m��v�Z�'wX�FR��.H�w]��TGQ�����8��8T��EX^k����
e�=#;y���;���Y��۵|���;Ԑy�6-�u�g�՚�Q8�%�+��z��OJ��-��IsW�����DЌ�i�PB���.�>��W���S:�u2����T��T���އ� ����촩��c:5_�\'$_��l�
�upS�UZg�&��sv:�z�ST�㷵6���R�ouM})��k����vD�1�-mD�//ZH�{r�ٹ��^��m,��b�K��\9��r�eTj�uT��U��ezx�d�sD��ؽ����2���L���N9��s�2�c��5;w�gL{<��;k����լt1��&+;�3͌�����6J�֒O�25����N�N˨�c0:���Q79P%C�*&;3p�6�W{o(���*ۮ�����6��i��G��~��&|p��%�\����T��Τ/�m���7��j�n�:.T}��c�rB��d�A�.���Vf�G�'2�NR7�#)��pa��Wh�fm���׸W'�`t���e��P����OV���#�ɪj8�U�+�{�\o6��dR��t�MS�f3v+�]%��9��N��Z���W��x�4ʨ����=�@�zז�X����#r&���s�����j���\c����S���jm��G�ڳ���T���=�r�:�XUnJiԖ�̸\��k���1י^���j��j[�B�����m^g>:���k��n4�W�*�����q�Z���˻v�⺞޵��1|���=�Ϛ��Z4sW��Tb}̴��vz���h/��A�߻��Լ횙�*w�!���jk�����8㗸����WիOgZ�Whr��)7�P附Y�R���V���]�oq�SO�{H���K|�y���8�9��n7�T%Ҩ�*�@�?�Y�_p�h�E�/�x�7ʏt���{�W<}�&�����&�]�S:��7F���o(9v�=�}�:�^ɺkO��k�i�\��x���^89�'�NS�`:ܶ��e	��´H�%�>2�"�29��ګ�^C�WR�%m�|,4��v��7G�F�n�8��RC�ݺ(��	Jl	����o^s#U7*s�@qRӝٵ��-�c��(+T���^ᔓ�����v�WN�ʵݢ�ٯ6��Gä�NW��^��|sۦv�k��j�E�-q�1�gd��[Rfv��RK���wf���|w�I��2���굏�EU�3�!�=�=�R���j�)��Ǐȧ[�EG��o*�r�xj��,�d� ��.�ǡ�z)N�.bj�t�'�����MUnF���v��Z�Y�#t5�o�_�N9X�c~���5�EY�گl��44�z햟���{e�8D�u0���=��vt���-t�[ἸM>-<�z,J\1����Q�9�uX�(��굮^����N�{ۮ���6�-��z�L�,�6��m�

y��T�cw_:.��5��!m�v1���{9Y�^'�ݵ1S��A����/��BM�=�3��N��N
��JJV���5�����q�q��0���]���vI8R�ةO�n`���"�������o�:���|�Yo����
G��tvcרwa��k�,Gܴ�r�Wq�`��0y&���Đ����B6�!t�m�,�O��$�!tW�5�e�T#4N���"��zC�r��tí`qR���m=��{H�t9�Ӕ/�V.ٔ��_)st���W��O`�t��r�i�˘3���ۊt:�Y�$cC.G �W[ӑ�qYW��7��tެ��PFu�Y��l�7"������Δ��t�O*Ğ�eԖs+_T]��h�h@���p	̮���q�ʒ�I��8�,ki&��|IXz��}RM������rs�oƶK�`v$�2�h��fNPU����NRTտۗ��j��j�f��J��[:�Xϴ�~���Y�c��6�!�y��nH���v�q<��nىF����v}5�p����t�Ƌ���ZA��ˁ�I���ޭs����e��ܘ+�jl=��/�ej�([��3�D�[�j�ˀ�w��p�7:��Җ��ڇn�=��y�]��=[>��jnU��M2J�,묺
�W)��q��@)d��ȥ�صB�	����G{���a�9O�tӘ��k�����f�Z2�n��֡��h��JAt�u�����@���:�E�]AJ[y�����\��L�v?�d1������+���<t,�R
���u,)�q��#{	�$�ݤr����K��N�W�D;���cm_�ݝ���ٕ+�V��L��g��X�륗Ox�
����E�C��k�&����j�I�'w>�hr��§���(��N�ҋ�6��/5�.{�?)�ר�iM�+�	|Gl0T�@K;�cŽ��$qˋ$BU⏃��h��J�9xr���ζ���J�;IBY��j�ӑ�|���^��-4c���y���4J�O2���_`K�%�Κ��7��z�
}�N�s���J�=�{���WI�y��Ͳ5����r=���7��)��/"I��鷃	d[]���e۱�%�S��5���_��im��#ZC���(�$�_JM�%n���fS�������K��Yr[��̹k^�_��u_�j�ֽl�`dz*v.�ql��/�kQ$6�j]R#��/C�	Rwby�;��OvА:��1溽ckBѥgE�A�3jFܿ�`��ܦ�9�v�M)SP���1S$���ۃ%v�F��C8̡��$z��D�}i�ρ��9W��8���ἦ8M�*��r��%��CA"n�Co"�Mu%�YK�nܡv����Ү����]#}]�A���z5��gG��m��=�;��K��8���qq0�@�+$�;�����C�׷�ԇj9�u���n6]#	sr���ح�]sa�t�h�|�oH������Z����ٴ WS'GmPy���g&9c��:��E
�*�YX�o4���U�j5�aA�&�v�Iz>�}���k����~��uZ�ME��BDR�CB�B�RP��@P�(B�!��CBP�QM+H�%	BRҋAB�R��4�B��(1 RP-C��DД�SI@��HEKB��)T�� R��E5B P�JP �#H-*�R�*� �W�~w�|��ug�^��ע�a'd�W"��^5A��Ɩ�҆�L�CP׸�0�`z˾L���$�n�K;*s��T�����9K�@�U��RM(w���&�)�3��R5���
͍�Y�m�g1�FR�܁ͽ�|�ˈm�w�xÅQ�B�:�ʇ�#��zȞ�Q�HN݇W�{�r�'�b�S.��I��mư�)�g8f���v�7�D�6E��Au��R{9�:s�ry�Y�`�Ӭ��7����r��gk�g��>�$�U~�}���}��*�}��������-��)M>�}p�Õol�;��f��Πf*�W��z���6Έ��0j�=$����w���x9��R-z�5��fQwn�Ι��x�	 gJ��;$���ˋ�
'����S)���u�k��v-��9q9Rwg<�Ճy?7�g�����ʱg���k�c������6-�{j�v22�3P{_����t߻��=C�}Y���j\�҄��W��o%�V���*����d���Q36��h�Ζѵ�F���aS��4����]�ƧD0���p	���u��1a��^^⟵��/��~t�f����w3 .�V� >̗z*�FJ6V�B��{[�E�֞là,�o&�A���� N�
y�nN8uJ�:��}��h��Ǯ�U�UX�~ǐ�"��M�kc������g��5���\7�������t�] �Te�"��a���������w<S�K�����b�=�y�*�:���C���ps!�G�U������:w���z�Oq~O��<}��fն2�r��!f��Y�FZ{`%�E�_f�8	OEi���݈���y�d@y��61U����f�яݔ����9t��K��B-���4�Л**wN�{��4ks�{���q?t�?qgk��m�z"�v��rz�q;z�ǣvb���q��}�ҺU�ć8ƻ���/�Cd���V�\esٖ�WX�}Ǧ�-�s=���v���B�
i7�ப#]�1�t���2��-��m�y�r�OV������.o�N�������i���i��(U����5Z����zj�������ܐ�n�\�Vv�co�
�JG4<��W(��v3q]l��!����*�.=X]]�n}ψ���דtw:����dS&�s4�a�.�Y%g����\R�=�C�vc�!x��ki�dܮ�q��AV��Х�e�/�2�>3{֤
)�����������98�Q���m�����[�]4ٞ��A�M�U���^�G[�W����K��)	5a�������c���w�g*��q�A�̵C�+X�P���\�S=����(�gP�Յi�w�ft\cj�<�47:��9eX|Y�O岤b����ϱ���"���	@�s�/z/�g��^F���n�r��4-�S�FF&1�B�e�8)j��5������>r�	͉܀�3���Gt�$Bx�>��bӯ����t]D:u4�=�p��8{Qo��K/ ��k�������Uӗщuk�A��Ғ��Z�[�_9}����q�$S�ڇwK��Y��ÜV1Aw��KEF�k3�w�"1>�r�ʙ�� �<�P�7h'*�Vۍ[��1����1�%?��f��y��I��/�'�I�[��tʌޞv��f��m�Z����H�&}�k ���j�<8�-��l�7#��r��8駭�3��z��0����F�����ά��H��/�s��]L�i�6hS�5�s�no`i�īV�չ��� WW'Vܝ��{���l���M�S�g�Y�R���V�Ü�+dN�ұ��R�&��{	s���q�FB�L�1 �[pi����k'W���,չ���ٽ嫞>MQ����Mƻ�)�����r��F�,{�O!s֓�3~ɺ~��ص�5O���u��iメ>!���e���)o�]���훥ä[ꁘ��y�+Fo٩�^ջ���,��5l��gjX�g�P�Q���e��Dw�$���/��z.;�g���dW^�u%K��L�g!>jڬۍ��F��C2����TM�C�6�mƀu��|��b����\��k��S�E���z��r�f�a�;m�U��&��N:��P��p�b�s{����%����8��rv]e���
J)ݢvÀw���֮.��1�t��ثp�&�����Y�J��+��짎�fz���r��~��Ʒ�<��\���7��Hg���@�vV�WN.~#\Tˡ�	`L+.��FR��1���ęV~����Ӕ9�+����+*h��4.7�%ؖV�	�axzc�R�چw�����8B�-��յ+n�J޼]�G�f.=FQ����vR�3�.om�k"^q�wA�"�T�ˮ�ʍ�l��.ۃmT
1��*�MFfKgAл��`{YJ����y>��:m���\^w��eB��P]�삠��C�ޙ�"��0�W<��aw=Qr�R������'�3z��B��c}�7_c�k;#E�\vk�\r�i\��@y��y��B�[���ު��y�����]����{��y��ö|��Ș�}VP�3/X���/�z^��Ume?aG��'3��[}3˘��d�}WSD�s!�y�n�ʲ�B/*z�.u��M�Z{��f�Ɖ;����G���*�o�&z���n�5�Z��X�kk���*:���8c�ӗ�l<��+N7k+y>����s]�Ț��9�΢b�;ۛ+�y<'���;�i���.�I�񑩱k�8}���K~{w�@ed�RT�!����@i��
	��^$gkۥM㼂뜘��YỜ%"��鰮���}`���i2��h+m�s��2� ��Gj����I�9{ف\���GF}�A&h�1ԓ_v���xG��+���T��狮1Pʏ^sF���L�Mf�$]���g{f���V����+~�|��61֮o3~��<��������ܴ^�S��e|h��uJ�
��c����%͋t���3�F�Uѱ����no5h�U=]��{�ֹRV�H�����d����'2�B*�8�x�5�/*�C>λܪ�n,y�i��#r9a"�]���A+�yq�ˌo[O;�{�(t� ����ò�һ�+����_�ov�u�u���rw�᭼p��y�JҨ;�}�1�A�yw�I�3ݩ�e��9Ű�_gz��5>�N3j�P�b죧#o2p9ۋ�Y����{�O������`vmFs�-(�잻m*eo��t%=J9[����s�cH�J`h1��_m.{���/��.�D�|�{�ɛ�f30򚷣y/[|�W\1c9�r�ąt��=�����vRč�R�t��d�f���H��HZ-��ev� ��һSNK�ZE[K:h��Y|a��sw1$� ��ܾ�Wa��gd�u����u�Ɠ�^�K����ɐ���خ8-�%�;�pO�Iu7\a��=�4Л����q��@��rv�5<2*9��z�q��k�I�a��q*@;�'�yë+pӒ =�ȳ6����;Wl�o�:���v'5���Q�Ȟ�0+����/�c����n'TFS޸�yX��N��k�5O+��Vn����OO]>�/Uu�QI����{+������R�㓎k>}Gr͆�ǽ����X�^!S�x��]&k���O3�<�_ݪ&+4Kc+�+��8 �%{�M7�q6�^��E���j�YW�śC��>��]�4 ��|�*���$�ވ���x�����x�p��9_�͗빯q��3�p���k2c�����Ks�m���u�={� 6`�P�o+���ަ��(���T�JTv�W[��Bi��Oo�[�4{��/Զ~p�5h� ���{��BI��R��_J�Ά�L�e�s]]$bF N�~1%�)�+�K4�%w�tT�Yu)m$��� O�s���1�d��o$��e��S�v��겅mJ�OF|�^X�f�Y+�P�p�
L��̇nW(��v
�d1꾜y^���?�d���ER�SQ��놔[���ѽ1f�{d��j�:��
9	IP`w3Q�%b�ӿB����u	秶:�f�K�`\�6�m��x.~�}P(t�˧��ѣ���TF'�k��)�<s'��a\�*��{������9�#����GJ�p��h�||�J=�̨���Օ�K�g�����m��L����O��~����s$�3)���G�|�`qN*f���5��^�WKǆG9������M_���ȟ���σ��s21zd�\��	y-c:�oy�_��dب�/���S�\��_5�\C���f�����'Ԇ%7�o��.��wՊ�e�'��ꁓ�J�=���-W�k7���wx�O�qo}A���B��Wg��U'��J�zﾍ�h�%�"���U�A�0�ӘR����޶<.3�/��s7U�s�3�b���^Z}�C����0p��-�~����fP5ߊ�"�:R>�|B�%���c�X�wpG�k�|��1듔���;O6���՜rXu�ݱ���tM\S!�e8xǗ�dSU"���3���'��m񚐛!�IwpS*jlNGf݁v�y3-L}3�쮽�o�-rĆ�u��9���j� 7���6Z������Pw�/^��U^�3��B�;�덺��7&�KN��/L>���&�lEW�.fj��r��iq���e@��\\)�e���;Л�K"g�d�r|w����G7�'��c!���>���y�A��
�O���t�|3�\�ǥ�F��䓭�S��/�QTn���~�}dUxz��g��uW��[���M��#�����O�{b��f0�L�&*g���	��Xq�GnT�A�{L�|�����W�]�K�v��\5�^�M��F����ѻէ2�`�/��P����qϧ&
�ƾ��fk:�l4\-�k���/�MݷvW�$d�N�?��;.�7>g�}@{��UHۇTðl�� �MI@L����#��Dڵ�a�"�觾/�Tw������H����ӣ�����e�9
F�nħ}Hb���촧<�^x�D�W���L�X���F�����m��>޶��ӺM��덿�7�#v�q��gc�b�е��>51��z�!q�ԧ�u|���ܬ��m_�_��g��|K�s����[�%�l�Z�M���L�W�.p����(GA�*���ΆuL����v�u�f#�6�ܭ�j��oL��������uS�1g+s���^n�����X����)�|�q^���k_n���{�nJ�{Ks����\7�-m�Җ��vt?����Y���3w������\����A�?\�yUP��UA.���o_����>[<�� ���K'�|k�먨�պr6�u�N��W�(��Z�c�=ϳ�IUѿo�U�_���sC�s ��<����U>��괡�|o+}G����W��/��_��ۋ�/W��}����s��l��������ur�W���B(�3���{׿���>��M'NV���:�ǋ3�1�Ӭ��]��&��#�g��UL������u�d0��gC�b�(迍*�6�X��<���T�<��ѹ�[�t��Q�<���~�1��Y����b�|P���_4�<���)o�������*2�َ�a�['5q��ߧL�\�gH�M�*&O��6���k�O��[���P�Yם�ޫq�Z��g�M,Ο���Ͻ����R��nT'O�YM�o�0�gъ>D�L�٨\M3�OtV�]zG����^Ӿ#���\{��μ;>��
��UB�	 07�t�~���)��
��ث���С��
ը����o��%�꣔I<�-pV?l:1�̷�db��3G<���u�%�R��M� 鸫����
Kf�Ղ��즠O:�eۣ�3�Kc�@;t��Gc��4� ��TՏ��F�pu�t�s���r`ɐ��0(F]��[�*�d�F�S|XdG��7��Y�DgJ��K������.(;�łjɗ�;�n�S�J�'�o\��ϭF�]WK�y���[���p���p���ǫt��sWN�1>�Z�$�,�<$F؅]�q�9���	�̽=]a��kG��ݙR��YLw5�P�z���c]�6[8C&.�\��$ЁB�nY�t0�hQ��q�EH�4�lV��9��{��zuTE`.��y�m��Hܨ����ɯVM�`���DR�ٝ�[LX[��]5w��E�2�œ��q�D:k�:9FSW���p��PJ�Y=u1��l���L�X&�g;��O7���(��&t߯;(N���P1Y��x��e�ҊN���ǘ�b���.Y\KO9kt@2�*V���ڡ�ܳ� ͥ���F�=0�#Z�K�z������K}Ϧ�殬t��#in�ެtl�����RU2h�U,#�8*U˸2Q��<W	�
�ʈ��:����[�<�*b�U�/�I��1Q׷����'n��˫nW<=��(�V/�z>�~y[�
ʹ��?S���c��^T�O!�����'���NN[�I�����z��^�D]M�d��,�U\#]�ۃ
Cn�d�����Vm#�2D5�� D�\.��1m�[Oژ�P�;X��} �m�bM��.��Z��G��� rU�%��l
��:Ѻǻ��K��T�g^[����H=WՍ�h�]1��Nq��^��ȫWu�8G[K��A����
u�pf�ŗ@H����ðJ����<�yO�]]N[��"xU>ʸ�gj�W;�]��Ƽ��≍�k��s.����e�H2�/r�bۨ��[y�~oQ�:����*��ҨxJ'�ˠ�"m��� �t��5'��>4��w����N\�2�1�w%��b��ONn�pc�ɰ��!2́�LV��c����KK�2\JD���X�<�k�|z_%�n`�ۼ@4-/�Ζ��7Qu#�٧����n����\
;���y��M�<�]Y�ˤNv$d�.�QRu/v���H+v���t�<EF��-�yPS�;+G˸�Cw�1ya:V�������оD�u6̦E>՛��.i&V�iٖ��,�I�jNv�벜��E�F��L��<�'�,�C����q��L�7��k���X���fn����S+�TN���"�eJ]I�*W2�t��cg-���K��a�Z|�E2�^t�7���j��#P+�'wV�'�Yw��e\4WXU�U��wm�F޽"�v�kdɾ�=���yn	��ν@VV�Ə�2��sI��xW�v���Gv�PB�����
�Q�JiZ)R��B�(�J��)T�)J
��*�
E�JF���hB��hT��(�* J�)R��R��R�J ����(�)��"	����)J�iB*F��F��)Z�:�U���y�����dd���
����oWAu����T���,U��'^WAG�X!���1��κR�[;;��[E�mK�iuG��
�E��~�6#�u>7^�A��w�9�<_������m�2��Q]�K��a�ٽ��-�'u[p4����2�F���ȧ�Bo��B.!{}k��H�מ���^�dU������b��"D�;
�o��yܟ��u�%��8�#|��^�8c�;c>��[o�w޳f;Y9Uz�R���q>��\6��K��n��L���'�+��/�n�u�o����,M��7��)�+z��`�ޗ^%�N��l��;���˙�/�8��Q�r��^O�37�6��,�{�Ѭ��������mׁ�z| �(�
m�W(N�E)����O3k�-�ok�7��U��G����|v�������=��;�6�|�{�zU����輝�ڜ<⯫��n���'�KӢ���ᑽ/M�����7�c>}�Q���k��,����<2d�=f���߯z_w����'��Q'�*_���n��ޖ<��<-:�dd'���o��#��t�wP>iy	�G�r��7���	��1�Mϴ�U�w!u��xn�n�W��u;�1�	e9�c�mAc�.�l\[���0���M
�݅�i�\�#n��ݷ��c}�N����'�o:=��啝éV�ŝ�YO#�-��χ�v�pEfa��ӤDޡ�h7Z��KBnJ+E�U�#�V�Wb����+�ڲ�K=��ʻ�{�C4�l��R)N`0��A�T+���A����ۘF���gg�C��c�<�>/ޒ��Q�7���xtgNI۹d�T�ѝ�Q��jiFP���w-�{GЮ}28��>�M�e�����ȯ+����Ӓt\[�O]+�#�'�3�e9���3�������*V����W��zG������Ey�{��qzsK�L����ʗ�=����,	"��ҿWu,�;ub��~2<�����y�ǤT�k�ɟ]�
�q�-�A��q�,�"�`L��Gۜu1�O�|$_Ο�GxG��D�@�r����N��<�؎�!�z��A�P�T+�rQ�"�A��y��o�W����j9�U�'L/P��֩-�{�+��|�k���ԇq�����0�J� �O��������r�793q^�~���{���f���֍G\7�l�ޙ��>��7���.=7�5d�fR<_&���6���9�������ۦ��S���5i���ޟ"|r�ý��^��̿I<�鿡y���9]�K��#Z�P��u�|��_O!�((Q�^t������dDJ`�ȃ��,�Ʌ�}}o+�8��-[��~�^�OQR;�T�8������+:��%��ݡy;`����\�.�6H͇�O��+l������Yڻ��.ƭn�znp����R�c���X���{�dr���k���w&.��ѿz|ϟ6�;SQ�$���|]\e�s���2,�����1��X/-W�k�X���0����ߙw5U����7s�U�0�}�<�Ǟh�޹��q�*��>��a\W�t�+���c«��@ϣ^	q��ۜ�)�CU^���<Vzh>��4){*Fid�^+�P�'�hӷb9���Ȳ���yq6}r�}�_�:�����z�y�y�W^���,G./�m/a�U�~��*q��-�&9�'����%��8�m�Vk��œ��m\�{w	gʳ�a�pv���������՛mE���3�&P��f:}#�F�O���+����x�S���A0�%}��
-���佘c�r�����Pp;讪����A�}�� o������֩׻�hN\X[5[��(��F���Zc#�*x�D��3I�/��W�>Y��)���������'Wc�����Cb}㹾�=��1�+�ɅH�<<I�*�GZ��k E�
ʷm�_�O�Q�6��ٯ1fF"cd�ڻ��p[�kn<}ٱ�ug�hR�=�Y��w	�1c�Qk�s��P�c�X�.�����}ٺ������P�M�� B�r�^�]����qe�(9y�2��͛�Dq;� ���T�MY��r�Q7z65r�މg��&�z�����}��=��ڪF�Ω�`�3�����w����UO���P>�~/7���*�_z�i>��\v�G\{}r6�=4̲Ad��]�	�"{�����j�i#�/ՠޙ�|7C�F�Z�ۆ�m�Φ���%7Q�~���DB��������O�|���!7�/�:Ga"��w�hRǯܬ�mW�(������A񎽓���>馫�����s�F@���hm>�:M�1r5.��
�(Vّ���R<-z��=I���^�Vz��}��6�>}��~��W�)d�|r ��*_V�϶�x�^�A�='�"��{Wj���}���o�TS�P���{�*�����O�T���"���}2j.6l�=�M��Y����>�q�m���o�h���R��Q=oۖ-d�_O�F��~�+ו��L�ok�|�K
rP�W^�x�t�εq�5�1�ޮ�{�=�4�p�~P��mVt�Ы��^w����:vv����·'$��������,�uK��v=u̩���᱀A1�/}����8�,ƍ~��[w�fn�ܰpGƝdǈ�(��A��yi��<��޺-���۱o��e+١��mIyrdpY��Տ� ���qU��GK,ҽo'+��G)�_=���ؑ|�U|���+��L:��}av�e��Ŏ��&��`�K���Z�c��(2s��|��㆝�>�o�x�[`b�u�۝�C�Y��a���L�wHw��U�N0o�~�2����k�/��� ߩ�Ď��J�t[��G��g�S�/�z{c�^Y�Cò&�|�*E�J�0�F�G������iߞ�2�	_>F�敍�I�,J>�n�@�W���x���g�|4�����K�N����3���P�}-��|1�{jg�XO.���ޫq�߸���z\o�3���\>�8ˑ��֫�Y"2��O��kGj�X8|���A�0�f��e��u�9�Rq����>^�[G{�4�����7�����e�h�1��|��c��f����&K}$_L�9݀炸��C�G���4 b�kl�WFAU�;������T���냦�^��fK4���b�z���\�}��s]:��z�qt�Ên���=	�_�}��"}�=:<K�� �_�&���eX27��"e�z���t:���[Rkv�>U~X]y;�x����m_��{ޤ�z� �C�]S�4����I@�uy�-jgtpҷ���L�s�؆�Vɳ�s��v��9��2K�\)^`������wH����V���&r�02�#�	����`u72�] ���M�z�a�a��Z������	�a�m:�/���̴%0la-٣��vRU��Au:���[�Ӕ�W,W���s��<��Q�;�6�W��~����b㏲dÌ&)�@�>y[;c5gO��>���������ߣm��VDoS�s��y�~�F2!���F��τ���O��n{����Y�J�Շ�����J�1�8T�N��n���<����זE��r�&=2{������-xb�����){*p�d���;�����8v� <��B��勉��3�˭w�tˬf}�R�y�V;�Dv�
�eH�x*�M�C1��t�DX��͉�o��5��ܻ<���е�d�e��\z�3�8������YӒv�'�6e�s�y�@�{�>�Q�^���m�C�z�wF�ˀ�ϏO�����Jex�_�ˏx�����m�_Tۖpw�-��t���dR�*/�6��9�J�DφP�C�:�L\u��������Fz��������q���&�#�y�������=��3�gƙ ��e� �X��W^*�e��۫qz�8g�C�Ƽ��׼��ZW{6n��!W�q�����*�nh)���s�sw�[��W�P}u�g	6������Pq�����ޛ�Jۍ-����he i�%��N3�
���0�$��V�Kl(4�;
@����^qڝ��Eˌ�K� �缜m��6�n�'U��8�mQ�a�!��h�_7W]|@E�+�u��,������;�:��#y)ޟ`�'��ޑ�}��p�S	���D" yQ�bbu��t��{�5q�z/\���k���\�1�6���μ�s��{cޤ8��z���SP�K��@��!,�����\Tx�]u�����u��j9h�o7�l�zgx��O����^�q��2KE���w���W�w���ש���D�R�Z:7���{�j6�W�7���N��g��4���'`S�=��X\%ީ���vj�5X*}=�C)��]��Dzߕܘ�^~�GW_��C��qքأ�r�=�7=���Dͧ���݌}#S.ۛ{�_YJ;����wz��&tؘ�5UWE׷�<��#�o�T���	�;�C{�RGO�U&\	�0��[�Q|}��竱Y�.*�\/C�޼������<i���>�#;�R3K'6��l��;k~�qѵ��W"�K����٧�jw���|�����c��s���;�_�wQ=q�z;���t�t�ּ�>Ւ���(>�՞L�΍�ʭ"Kd��e���W'�Y.���7}�۵�X/z�s�BigϢ�I]Ąȱ�M0b�G6���yR���J�4#&9������]������o �oc`���:z�e�}���6���+�f�W-Hi^���{�+HHn�g�h�fIǏu>��+\!��+9g,?8�oJ޴�؃U���&���?Iӷ3�*�_�t���4�y�� �z�Bt�|�}�q���*�d�PHJq��]��:����vQ-Y�2���Ϥ�9��V�x/�s(�:=�^qJ&{4�_&"b��NS=��!��9�\�4�a�ѕL_�uJ�8�*%�.� *++�Ts);���z�gτ�����z��g��%�,���8ʡ����
���s=ͨ�n���%�S�\M�:w�+�yν��7�R6�S��U) yMm+�v;���2�h�����`�-�ՎG"����W�#�Ӿ+����4���#;�M31��cnи������%@�DO���끾2�X��9�o�֩�u�l�A���t�t����f�T�q��l��8�W�'�&?,DLI�dt��za�=�#RT����'}K�Gznz�\�nwix�㳬9�4�ߺ:F��t�~�YC��.�Z�J���<=��p/Ơ7ѐ�rĜ�<���m��>���Q`8���S���~�O�<�"�6
�޵��UvMe=~��Ѽ~�y�29����S�S�!k@w8�;|��f�������@��N�\�6���N�,9O���wY複��$+�^�*�k)R׻G��nu�OW^���$�'IH5�:�ڃ\}�Vo3κ����ꎯ��ӑr���g��CW�p׺�3�utm�U�_����_���O�U �|w+1�߬�g��b��gI�kN��Y������������7�{p�]��>��s�~ܱh�&q�Y���Uwz�[�� Y�|rpz4��VRB�|O��gZ��D��i��N���T�m's�7�)��"�����W����~>�grsbe�T��*r��*���_F�G�C�^�� ��������Y��������&�����a}��6����?^~��\�\s�4�<���*�`�m�9�O�@�{.K��������X��.��2�Y,�p}�&�!���9?L�S��F_ܦ<�A\�{�b3IeπO���B��Q�y���^Y����쏦�.ʑ�r�<j$���VЌ�>���t]Z
�w��^�p�X�u��k�ޯi��}#�������^u��9\�6J�;g,5���ޮ�\��h_�l	u�2��'�S�u�U��n��";�<_�}!��j�}eC�o՞�w�W�-�x�^�lv ������e��u�9�Rq���������`��8���۞�W^�cf���Q������,�x�9�9~��W6Ó:g=xoktm(��޵�ws���$m�S�hx]]�S=#KMj�
��Ac�V]�ҥ����sC�A�#�Bwc��#4)S��W��oZ�Za��&>k1���%Jŝ���q���]���ñrYP KO����I�+�wC�
��~�8_yyw��%�n�I{�gW:J���tƧ=��=냧���fK4���b�W���\�}�۟=��eu���{K�~�k$pOΘ�sĿ@���7���.=~��s>�V���Efm�jF| �����=����Ս\{Ǽ���j�G���|�z� �`u�9�&r�x-���^�U/y˭�X��L��ਉj�U�]y��Ƚ+�~�{Ϊ���F��P�n�f����S
�G�%*stu���.�\��za�����wR���}~����;ˇ����}�Q���p��W��<�\��`��YGȬ3���U�j�ևT�N��n����=�U��e=���=7�>Ļ�Ԏr��V2*gl�����Щ� ��ew���:Au���*�ܻ���<�fj�7O�ؽ�ឪ����/��c���ip]�	��>�n��e���m�_�\�W��z�٧���+D��w�G����箣=Ӑ���+�Ft䝻�O���/C�V�)ژ5��~���AT*�㮅�T*ܬug"�1�3hJ�\�`c�������j!g�[(�ت�u����_`FMp3�J������g��L���|7=����WTW���2��a��[b4���y]�6�Efo[���\�(��w�f����y+��]:�ػ��sf�w���d���7��e�ɋ0 \����te�xMQ�Y�>!脞�|�B1c�K�*c�[	r��wq{ʠ�(�,,J����625xԻ�n=m#C-��,vv,2�73r�w,���eJ�S/��5� �u'Xfp�w����uG�^�u�]v+�	=,d�3�2�2�`������X{�����|%�y�-��Q7m�7��9lK��>&��B�ل&eI�1���"[���h�q�`�n��:��Y���76d\28��M�os�h����o_=��9�)��+t�������y��ډb<�Ӄ�p�	�gI������wvrV�;K;�^����mng)��NH��d�
�]nҥu�Y��7���3vӫ�iQ�%��Q��O)�Ժ�����l]�u����ɽ0��
ׇ����p֬�m} �wo�5��,�j��n}0_k�wR.3�C�U��Ӵ�M����u�݊]jb�k����/ve5vW[p�՝�Z�^-Qҙ���m�t��;��ކs��C���c���N�TR�@�-��������ذ��7����e\�����ꖄQg�}��;u�v�I&�a^6�ݡ���E�(�����y�ta*eƌ�$�+��ؾn�r���}��앜 �mn�g��?w]�xi�ι�k��Λvk�tN���c/M�Ǚ���ջ3F0�6����ka��1���,j�t�i�g]*����zs�ɱb��I�]���q�j���W%9�mH�cq#o���:S�+x
�5�*8*;4�ۦ���h�����lZ�o�@i����$C�����ܱ\ �u�!��V1��4V�m)��ܽ�e�LH�p�z4���X�e�:�Z�ĺ��/_g
NJt2pDY�Yٻ;��J�+�ͦ��wZT�Ȼ&�ٻI<P
[]�z��8���s�3vܭrL
v
B�e�W��h�+%��A�⾻���� ��߳&�'f�_aD%A���"��
�����:B��9w�c��
�#L
H�
�E�,/�Fﲌ�3dK/wSN���!y��}y4��*�gV�[�Ep��N�����m�[{W�^���l0T��Ś���`u�y�2�}f�����n0.������-PW^��C�3NGk��2��vWn���o]�v]D��f�|hr�/Q�*D�ͼ��ux^a�Q+g֑���cL��7��c�i^j�Ԝ��;��&���c[�j�[���P�a�7�� �ZA������n쩠�)�^�6�݀p�H��#�Oi�k���?����T(R�hB�Z
( �(Q
)�2�\�
@L��2bZ) )R�!��A�L�r��Q�@���h% W$�"T��Q�Zir�X�h��rb�������_��l�8S�/���$mN�{,�57��5�B���wT��}�o����w2E���4�D��Y��
���~��}r�y�����O���r�}޺�x�+��m�J+$�6�/j���
�o�K��J����'���Ltu���z�8�O�Q�>ӏ��U��V��q�7g-zV�H���9���a�i���ȱq�J��eK6�Պ�k��¥�7;s>�sR�{���%���Pg��w�3�0��EP,/L���mκ�>B��r}��ˣf^S��R�=��^��|�>�=�'|��;%��D*3L�n��gLq�̧�yA�]�E���|�Gx�k�O����y���'�鑽�&��sP���=���s0�B�y{��K/<G���ƙh�ߙ��u�1�߭��s��Y�V�q�z��Ӟ3�5��Z�����\�.I�2Ϡ��7���1>t�*����
_����W�7��>D��������Э��C�v�n�v%]~�=魙�^<zj�{�V
�=�C)��]��k�G��ܘLvߟN{��n�[��J�5�>��XϟS?C\b�D�pdy�7cHԻZw�5���\u������ѵw�;f��������㒋��Z�QekF��V$N��n�?4u;sG	0� c����`��O�B`�4�.�-V腝a�iZ��v���[��J����G)Ӥ��|���L�m�譵��Vm��)�̚8;�x��v1u����{�%�{�J�E��So��'����T�Q��U�}tNa�޹zt 3»,ϻܯ}V^{�lp�μ�n��q��x���^���B��R2�e���f���Oт���}����y5+Iӑ�}�}���>uU�s;�T/9���r�Tw�$���OnEϧ�5����[��k��{�=�x�[�Zn	^%9.�:�'T�|O����Ka��z���Z�������L�_zN���c+�3�uO���N���� �4���'K���.��+���x��+���"��ٕ�^��
����s�3�u�|���A�������﫸��{���Y����z�܏z���J�s�R�F�OT��FU1quJ�3rτu�|��ލ�n�z%{�����z27�>gs}@{�޶=�"''��%E�U��%�̲�o��C���Jez=�q>7^�\M��ߴ��:�7�����R6�S��W���=W'HGS���͔����8�z��+�����#���*�^��|};��?H������)S��W���"}���/��O�2��Eצ��Ԧ�4�nf_�^��p�}!��s�;e�#s�	+��]c=��J�m^{��E����!����ʶ�̎�\�d,��2��t��o�},䨰ӵ�"2K�0�wuӮV� {�JSDoU�n�޹ɾAo�?�̃�["�"]2�p<�cs�޵Hs�Sfo[f���ϣ��g���^���x����>�=�T�25̖��L7c�������t�{b�{��-�Y�}WQ�W!��*u{G���9���y��:��,��a{ Oa��}^�q�-t�ތő������'뇴?|��C�+��������w?]�4���|r����Ώ�}C�^��4�����������������p������g��X���T�P�Ĩ��G{���Wn^��s-k�p�}'�S��q�>��u)|o����7�rz��9�\��C��Q~]NpeQ�^��S��\��Ӡ�J
�l���exmº|O��_��ڸ�D��q�^�w�J3�{'��X���Ƨ3�仜�~�e�͝��go��gC��t	S��K����q�ݤ�fd����}+��>�u�+=��Ӝb�s8T"����"ūھ8i�j�ª�>#��{/s�x/0=��22+���r=t�VE:C��=��3�b�'���0�ў�l7�P@�PU��jҞ���WZ��n���~*���y��N
˽�V��_��=2���"�اf]�y��S��1���������(�d�|ఖ;9]Wt�e0�͇�py�6�Ky����;��F��]+~��ꇦ�M���`���B�?�~��2i|������P	��v!�i�����z{~�W��z�Ϧ��E�t�S������^=����V���u����7�(K7����ޯiȍ����~S>s�"r�&+�A���ٟO.�:�Y;�(z�|�J��]Ss���|n+ޫq�߸���z^�C=�9�܍��e�X��&qZ�T���o�犁@�����Pe�0��[,-w]��Rz�hh�H��8z�[���Ω=8���{�tz��qD�� ������-��q2��t9��Ndڥ�su��Ȟ�V�����z�2=;��lC�.&�=냧��`�T"t'�����3�G�j%:��G��w�yak��s�k$p�o��Ͻ>�O�����_�8}����9�L�6v7���ݠ��n�����ݯQ���h�%Q��3�W�7���� ;����9
�);�PYT���-�g�<fo��8�tV�׼z�"�����G�����^&�ǽ���(%��m�gvG�ng!�}�����Lx���O�_�Ӂ�Zpe=�
[���;ˆ���ť����T��Ε�T}��C��N�u0�.�t6^�wCْ�c���:�������eh<1�U���S�n���V��K�*�m�M���6�Ѽ�X+h��U�C�$���b�sՒ��.��E�GYpWe7"ހ��$�3�
��G@ȗgeC�Ý������_-�p.��l��G���{β�Y�*#��U&���}�B�<N�u1��ⵀꀻ��Gn/J^������}��^�;���Az�l�d�w�az釿VW��e�j�<2��x*��w<��ڮ z����U��g~~���άn���Ъ~��u]~'1��C5�SC��^C9�Λ����o�ʙ��O"VF�`
ZײFS��I���g�s�7H,��³�$﷧��Y�{2_�K�:�%5�X�}3�5UG\u��7r�y�����O�ĦW������ϫ�� �9Rj��=�Ńۉ���{9%��$���@��ﮫ�1}n����z�<��7�>�6�z<X{{:[�k5�j�Xm�o�7�;����2���!́s�o9���1�M��<���\�?~6����i�K���=�W��xＪ��9���rQ�|I@�,�28�܉]�π�u2���t.B��\��=
��н��y��i�l�8z!Өw�P���Pf��:e�-�S�p�Z�[�;�'�
e�����_yTR�W�!�9��=��!��{}R:�T�ǹ#�w�ڸ��f�U��)�%�����ݧ�Wg�[��3
��S��xn��8{`����ٱ@�=l�K ��r-Z{�4�gxI�}�V����q��5�� ƺ�rM6��/o��u�7
�/�����3�n�t-��#h��e]f.���.���Z���C� �F�=+���h�v��oZ57�l�w��G�p{Հg۠,�ּ>��7J��/g�pQ���Y�C��ѯ�ѽK��#Q���Q�z|���6��YYs�~�y�烬�ә�H����^�
�T��n��T��5�#��az�.��ڋ�AQ��*q{�ǣ��Y�q�O�w�:����Y�k�Y=P2a����koFӟi��{��9&�v�Ϯ�0���/��������y�������Ī0���\�Ş��Uf������������-��μ��n��s��C�^���t���[�+���+s<x$���Q�X*�-����_�L��WYI'�N�R�{iW�uU�s;�T/9���r�n�>T�����x8۱��^��I�Cr�,��[D��b�,��4��3�ߝǱ�/����tT�e:��dyUe���Cs�o���!��J�}��.YKBg�����\�9_� ��>���.�)NW�u���;b+�O�L�{�7<_
;4�
���P�^��k�o��e���Mȱb&$�c�+h�N��tw�̷o����[q��o�ʉ��:���;9Ӹ-&չ�ڙ�À+d	�,��ٲ>�
�.��r��H�$=�f!,�\�*��P��QnK�����C},����> �}y�z��`3�ܝ��R�����)��u�F8��b��~*}({T�rR��N M�-�wa�q�9|A��g/(��S�neD����<�޽�3��ڣ޶=�"''��%%1��G��d��/�Ҽ�tu�ۯ"���q>7�W���װ���<���P�~�R6�S`K:'\�U��gۡ��Y9���&�^㌶^k��C�+��W�"<s�i_?H���W��zf;j�:<����B����Ae@�䎉n��/ō�瑸�j��>��t���ҽ�N�v��-_[���g�zwI�O�o�^2)̖����w��"d�)�p������Խ��ןnV�	̙�������^M_��G��ώA��x=Q�*:�E����=f2_W���g��*�s�����k�*���yz�=q�w#��UT;��x�`���q�W��r|��� �|^�I~�=�ygs�QJ�>�}���i͹h�wT=)�u�d{ή��������`yV.;�RG6�ȣ��ٽ�����Y�%� ���
T��n_"�z\Gm����v��H�.=�Q<������vP�a��jQ���mv4%I�is�n=���n�Uu
c2w���}��l�Ͳ�ʶ@ġf������|��-�>J�p�pS#�Dx�h5=��G�ɹ�%L��y;�����K'.-Ү -����u.o/8����R͒dYX$���~3���6Y��{K�۸X��6�-�;a�K�W��g/�(h䰯᳡�exmº|O��~7��=�����#�'����q{��R�3ގWpz��f�g�3�����|?o�gC��tlU���]L��q�>��gf�w˜`�}*���w�Z�����v6E����B�t໑7T:�N}�Q�e?:kݑ#�5�;����� ߼i_-v�de7��9�������ι�;Y>Wa�>n����;��Tm������tm۠��P����Y���}r��~����o����}���G�|���)ʫ��6; ��2>��6NJ��}��u�[����F�G�܍���:��l8�4GҦ��L�z�н �>��'�e�!���2��;��E{�bn#��q��H�|T�>�����q�,�Kh�e��_1���w� �x��lj<��^3�q������ȯz���Eqwγ�����j{�����{�a՞����S0��f�P@J����#�^s��`� �c+��s�U.���V��^v�A�����]��g�pt�ޯTK��"t�u����#��70��e�1�-�5Qs���U�j=b.�hMn�W`�g�8���m���u��}Y$��s
��dH�����$�X�m�1(����4��.7eؽ��׏�A �Ü��/NJSJ��X`4b����t�?��9���Rv=�9�S��:wE �spn��&�2qv w�Q�
�2���j5����:c���ӣĿzp���Y>�R.��n�j�����W�t�Ϡ��2�J�¹cf������oCj�F��R�=^ w��� ����!���'x��e8K����Z�%�>���ȷ�j�ߌ�4�*9��<�ϊ{+�їLh�#"L{$(�^�q��݋�VL�S*jK6��m��
��|n9�\7��^�]p��GM-�r��ǣ��F���=?^ٸ��3�㏉T2a�Z�i�����<�<.|�":6G>�Mﻮ�1�זF|����X�ٱ!z�l�icv���D	�0�/d��-����YRz{��]��>�[^sU�D^�_�|�z���/�uc��ݓ£=�#.�wx~����x�ex�#�·x���	�|o�u�Zl��Ĭ�MxP��d�e��\z�3�9���x?�Ɏ��F�������E���IN.@���a�*�=r�1qXU]2R)�N�+�{:fc�F="�O��Iz/�o�8ܝ��2��3��]W�b��	so�V@�W�C���7��{᰽,��c��;��j�H��-��Vm�U�.e���n�-�����&:*�һ����5���G;��Ȁ���:���oLq��ͩ>�ՁQ�c���˛\�����e�F*z�(u'E��^nU��Ȟ��O=�Ժ��M^�B��{��VEy�{��9ơ�(ݹ �}X �.:�]x�,ʖiec�N-�"n��JW�W�}���4=Lno�x���=�>3�0�\�j�%Q��
^��v���꯯m���5/ͨ�n9���]?g	��FB�W�[ޡ���HN��t��.K4���&��z�V��.{څ��ߣ��mx��fZ/v��m���_��g'���ޤ8������z�����#0O��l^99�����|������p<Gآ��oZ5m��>'8��{gj=˹�Ǻ�������Ö��=߬zq�Ih�?�H/�¼��<;`)~7�F�nW�;�/Zy�z��.�Bw~l�}gQ/ :��3#!zh����U���xм�K�gܩ�Sg��¡xz��U��5��?$�����+�z}���eGO��5�"�ꁓ��T����xj��[����w�2��s��[5�j���w��O�r-�:�~�=�x(w�d��Ta���ݎ�P�s�'w�;����U��讯i�s�-o���8gUׇ7U�8��<i����x�̌�eH�����{.'P&^9:$�f��_�p澠���I���ھ�U�Ū�ႥG��6+�E� 諗^9\\!X����C�J����Z%���˔�9\iV_:.�%�,Q��I2�;{r��)�z��iS�f�8L�!��:�¯Q��`���	��t�p�8�kΰ0��Vz���)�_X�x$�TG�bC
�n��3,S�Cw7x�eZ-�ػ��#��IU��:���uEJ�Į�
ǫ��1��Vv���:T��iY�l;fS�y��JO��eԼ��
�w��z�gu�̹F�X`n����1Q3b�Tk3)��[��u�u�Pr��"���R=	M�rgU����Zn�N[�ֻL��)9��{k�;2�|�liK�<KWӑ�$LG�U����;��9��ڴsk�ځ$�WaJ�:�\A�0�����|yҊ�-&�\�uٱ�Yβ�ʉ�8���Օnca�KtQk�l�	�S��gT�iTM)�Ʀ�y[p*oe�5Z����\�=����
�x2i��`�@�6�a�;��2Ύ7�[i㛔�f���츍X/�<N��'[�8�*�-:�AJ�6�R�ș�z�v$��ls}G3+v�6�W�Z�f�=G��u�ʑ����A[p���q7e�<Tbۦ�ޝ\R;��	�k&^��r��$��Bf�˸%ܾ��|&��&$�˖q�ٮla��L�6oV��7�/b�ݙٛ�{���]�!\E<(�W���Ye��/�Ǉ�����ׁ�����^�ŏ�q<t���;&Q��K�]v ,�>�c�m��uwDӸG6U�XӋ!ŚC���T�Ò�ӧ����rڽU��S��T�e:ܿ�	�lݬ�]X�X��A�e�s������V�*�ukDպ#��seq}N���Rx�ħ׼u��+(f��E��EJ�V^Qi���ÙJ�W��MR.�7x}�{UD9������y3*ȷ Oum�d|�/�����g�Vړ,��@1E��0M�ܣ�ݨ��{��t��{�8Q@���S��e���c`lv�kKpsv�[7>��nl�4)B�3#�y�.M��s{�n��>ggQ�y%��u�.�9�2�@d��7q�P�J�ۏ�+��ץ�0\�"J;3�D;P����h%�id�?�=�rw�!���5����>���� �ڮ1�H�'��QBv��$�x�,��:sd�{�;�����=S:�2�8+u9�E3G1��]7u��cRP����U�����'q��T��x;"֩r��t�ǹ��:Vm.+3�0s���Yqsô#�to�1׻������y%4λ�n��QI�D�fu��U�-�v�O|��<�mz��2�d�=uŁ})QЧC�*c6e
	��,l9�e���f���=z�ሧ�{v�#���0��T�7޻�����C35D���$�8�'����ݙ�~y���޶n����2()A��2 )Q��D�22QJF�
R���
V�Zi����i%V�D���Z����((
F�������
���Z�
�
D��)�W�Wݭj<
�j��y��{���Ӯ*�Ni9`�\7*Vq�\��*�i���Ec�͑m,���/D�|fr�ʀꉝ;��q���jׇ�6k��h����ϵK��WᎪ��g}��9wQ=R {]�*������/���H���r˓�^9[��*#	b�>���\{>uK���[���"]�ο9N)�K;�J��\%��8�ay3��zN�%��<�׬�ύ:s�g�%X����~�����_w�o��|}�x�SW��Q��;*t�E�O�,^|�b⺫�G���$����×���,q~ua`�W������VEz��|cavT�vY'��0�u?��S�m��U�*�|�ԥ��K�o,C�޽���;���q���99<��(�!���[�Qs��|�<T|Z����}U���r��W���o�q�j��m��?eFl���e)��w�%T}� nj$�&u�o��^k��S��z�8};��J�~������{�[~m�T���k�î�(!Q�������_��yjP܆�+��=V���dNoC[�痳x�]����wI~�A�L��nd�7���A�hb�Kǭ��U�g���-�˱U۳Sd7:|rk�2N�vܒ���[K�(u.^��c���ˬ��_��,0k��B�볰� j`r�f��%�k��#���Ϙ�ֶwM�2������wd7:��]�GV���*n�V�2Ʃ.�wK*/�-UX����]�֏{C���5yW���g�"�|K�ꌁ_C�Q4���&az��cS�y/�W��w�cuf�{�G�r��YW����G��������o���0
~��Qd����gь9@�R���ޱL���KU�r6���g�������utm�S�x>A�X�{��gcX���r������9N���
��鿣n_#�%/���{p��W��)��lJ�5A��+�8��G�r�&o~��(�,(Á�exm�
��<sz_��vڸ����x��w����/�F=�t�^�z�\~��P��g�>;;q3���l�w9G@�?�Ϳ�����w�>��&���->@z{�<3��/g��N3�ޫ�[�3�3�aN홇�'ȱQ>ی�Q~=bw�>U��>���4���ߌ��o��s����Y�:C����Y�S��|��F��ǗY=��:罾�Ϡ˨������Py�v!����g��}�,��hxv}7\�t���HyYM��e���
��9*>�[%1,����<����H�{���~R���׿�|��%�֗(́R�μ�\S�\�7AD�����n����c�mee{7���Q�6����c�" o��41?���x��Xܡ�j�JĝE[2��+��G�b�[����Դ��븁�6kLu�^E4kz�q�UK6��\|���^R�'�`X�w�]Ss���V*���������s`�Zx��Y�5!����A�e�@6
* @�8)^3q�[,k��Z}>�H��Fs_�����|���>o�m�uF{�n=T�;�%�P@HzH���I���t�E���t�Լ�W��^������н^v��u1��~��o=냦��z�j��B 6��2�Q���ˌv�g�������ۖ��j9޵�8\7�ldz}H�g�ӣĿzp���g�}�߂矮�bm;3�2p/��N���^�F����3�F�\�z���y��o��}������G����1=9�9q���g�'������b[Ě���o�t�z�G)|n9��=��;�=1���]g����uv���n���wGы��@{v/�>ɓJa�4rX���*V����+7��51��ާ�y	���r)O���j��}�Q�l�O_��{g��͝�>%PɆ�mhw>ӣ"�¯���X����=&��L>ڬ�u呟>��{�V'�6�P^��9���fa{^�����-y~�k6�
���B���/z��0�خ�N���!gh�P�����5L����sJ��gtI�6�+3��Q���i'NV��oQ۵\g&��l=�6�=�N
�qR�/�z���{YF���+(ghB.�i=�I�6,�6����<��͒�y_�1���^DJ�65[ T^�_�:�^�;Լ^G�X�9�<+=�#���)�ӵ�7�s|�yߌ�asb��M��~%g�i�*��,�zK�]F{�#��	@}�;���u���ln�+�f�\�|6�^3�
�����:���9z|��x��nW����?nz2$T973�c<�^�Ge:��{m
Μ����I�C�O�3���t%;�Xkۜ���w_�[о�K3�@����=�~++��݆s�#�e�rA�2��ȱuҺ���Z��v�y�>���U+ҏ�n�W/W��p����P��y�{��qD��P,L��ꏓC���ߜ�^�\��_�㩂�E{��E�~��>g���z�����:�K#7�ca�s���:�ҿ�3'��W}2�^�5����ybv��o��!����T��R����X��Κ�;{c���	��O���<�2Eķ\��11�^�j:�[g#�;�߁�Ġ���k}�ؠww�����h�`�=�z��f��-�Rٿ�I�P�R�Ѫ )~7�j5!�=�95~�����<�����~v뗶�FF�������l闯p.�������kM�(Q}6=��h�WcV��U,2�*oE�:g2�u���fWl��L�I&����|3NA��"�O�*)�;����Sֺ��N=�,&�T�qQw���[K�E�l�}Ӿ'��u�3.fFB,�љ��Sc>�=�B�-��Y'ݾ�"����s�G���B}R����fM�����*:}fI�Y=C&A���Y����fV����击�6�^��uxu�;�'�	�:�����w�������ĥ���j_�N�j�Me����O�'8�K�ÿ+�q�߹_�μ�����}�4��bt��hWC��zhW�V"z�՛>Yƽ#�s� ��o�Q���"K�p�R�n;m_�C��s��z�yͺ��Nf�k�'�ٟ=]��{-��ɾ,9��O�C�ʮ7�x�p���+�d�{{*�j�����z���i�}�\�=���K"g��J�w�Yr�=0c�B�|��(����{G�V����7��h�~Z�Η������즮;��1��S���'���P�c6_�$CگEV:q�YϤ��Pe��Vo����=^���V}�Cݐg8��Gl�O:�ޑ=�-��
i]]�>�.�/n��NB̨�qM�x�z3��O�܍��z���rx&�4t�
�:<KyB���f��ڕ?��!&��uf�v�0�N���0V\cD�X��;b�5��J��v��GTP�r�M�I/�{e� ��]��ի �z��ꎃcK�6�+*e�t�spt+(�H[��р���U�F���,�Ϧ�m���z�s_��I����	-Tz��l���q>7�u��:w�9�<�7����<f�6��9�^��q��:��D�>R ��n���ȍuc��~W~�ZE�Eu"��M�V�{�]���}H��}r6���3P�Ae@���1-�q�_���.��)ښ��^8��O{�%��+��a���|��{屢�/��bt7kZ|�M�Ec.�f�����#\����dkj��}E�A��x=Q�+�N�j!K'�L��ʇh��{pu����sk�o���J�=}�r</����M׉�DO��dq�W��r��=�ޑ74�Ƭ���ϧ��<Y��싲��}���P����y�QQ������}����=9��W������2�҉U �����]z�M�ܾ>E"���ۇ���]���3�]��9aYڍ�VO���*'�,!왽��(�����++�m]>'�F��]�g}5`Lǹ���)'�M{�c~���;�pz�?��4��g�>;;s>�N�&��������E#
����^����w��+��^�eY��O�#��N�س����6LB���W�NK9���7A|z�뤈���9/t1�������ӚN^���"n�;�iK���Ij�)t�v�����d�ճ��-��@�غ�t^婋�Edb�Z����/R�q���z��]k+=��Ӝb�s8T"�ݿ������Hρ�.ESޅ�w��⇢����P	f�`-t�d(��~=t�VE:C��=���:z=Z�ۿ[��r|�x���c�hʨ���]ѿ����ýv!�zȸ��z{c�^^�C�z�/`�����#���C���^�d�5S5UC���Q��%�������W����/|9���^ˤ{b�{)y���5s����pP(��X$�,�yT;�����חS���Ш����:�辵���ޭ>��x��}���^y\>�6˿��*�,	
W��}�[,Ty^O����O�6*�.��o��DW�1.}H`^�R���H���\��S0� \�iA*��"�F�
���T�u��\��IS>�߇�����C�z����cS�wy�\7��D�K2v�9������ƫ,	�D	�`�OQ�떏�a��w�H�i��>�O��'�ޭRc+rbӱv��<��З̾��bW>q?�I�u��G�Kl��V|�����u�ڿQ�{ԁ�{�m`��_�z������-�dhP��mc� l;y� v��U�-*�K�e���FS�{Q�/kG���I����.�N�N��I& qm,�*'دl���"v�Z49�dА������j�9Z���+Ŕ�h(�'��q���hs�@�`
eɜ�S�xQ�~7T�/�Ele���9�_���q;��dmZ>���)��Q�[&���P���_dɥ0ʑ���Oa��m��Wz�/��r�D�j�z.���[=�u�����I~��~���}�p��|J�0Ս�w�Oɚ�xx(yn�]��V�'}�^�����u呏�Az^��V'�k뙳�id�����g�{���_�$�?/�=��p����|]����+��3��e|�K��X�9�<<_��]VVrq�C!wao�פoNg����{YU��K�+#M0|��d��/ޓ���t��"&�Ύ�fע����ܰ-�'�`��{)
���;qr�co闄!�r~��rW3��x�����|4�,c9>��I��,�<�����y\w{O\�fni{ ���J���)UE�%˜ԧ{=y�*A��Y]��W��:�8�x�
~�Ⲽ�=���_#�e�$���&�,]�ݯ��^�[{fG�J�>j3��ϣs*Y�V��5��Т<���Ϸ�<z��q��9���EVA�<6w�O���5��''coh��S�kHh��Y�� ۜ��5׳��-�I	����rNW�l��(��=5s�n0�l�ز��!�7��;�E��9��]ϕ\��{�ؑl�͖3U>\D�F������Cod��5�d�(��]�����vT�$��B���ٟ'9�����-�����2�#�CO{e	����23��¢sޜ5�*�5�V̔@���q<J�x���o��+��h3��;��C����A)`�x�9�ԣs��H�D:�	���.j y�DI-���}���GZ3ߩ#ޯg�A����cl8}�c)���n��zk�CrA�I���K��x�َ�-�K�[��{���Ba5�R>��W�6�>D���>A�P�̊�E���3Ц�K��v��G���oc������kЕ>7�R=?+�1��FJ���;�FWO��5�z0��7Fw�n��r�u��^������ͿR�Y�^|��1���C�Hu*��O_�h�޹�Nc��0�+�5q��uc�_�1���W�t�/��G+��W^�W��>�y��a���{�]�3����������!=N��)��b�����%�]aez�_��m��s3�s;{���-I���y��bS�����ܛ��Á�Gӡ�eW�R�J9e�ﾗ���KE�~&�����yƲ�`�0[��5�#5ְ���kWM�̚����y���R"��N���rD�Eh,7yTm�fYP_��;U���1���,KiT_:�X����"�`�f�]�YB�2Z�ֱhLAfX�e^��B��»���F{��?Q���q&Ty����%�~'m%�%�]W[�g�.�t�窅W�;6f�}�W�r|�A�����N����]?�j�#�Z�TgeN�� X�#��
<�n�����l7Ǉ��^���hw�����/�����~++ԇ�"���eJ:y�[�S�'�@|n
c��:>�;�7�@�1�bzqfTK����<���ћ�3���=��[��{ڤ5��ɪY��t>���֟|z��w�]0�k���{�%˯a^#�u���S�u�p�_s���/��*��Y����X�q�[/#]X�r�����s�O���kwe�};����e�L�:����,ι�Y�����Q�p7e���?[Ȩ�Z#���=h�}ڦ;!׭�}�m����&���}3�#b�jl��w���^��P�Ճ�ܗ��s�4=
�y�����djj��}E��"W�z� 9s��>/y��U0}0�N��ʎe�y�H���]F�.R餦�Z�\7U"�*d��>���gU��"��"���ʂ������+�*��PE�
�+�B*��PE�
�+��*��APE�
�+���+�*�j
�+�T_䂠��1W� �"��A��W���+��(+$�k+O�!@\�B �������"Cx||�A%(R T� ��!T
PP�����%UUJI  HP((H��w�tH�Q�H�IT��H�E*UJ�"%T���)M��
� �U��S6*j�5���I&՘	*��
����+��E�C*#�M�  f�  �@h ]�ca�f�%�����m$Uh��m��!AD�hŭ�Q�ȔP�*�"�tbD�TQS`�S�R�̊*��C�BWL� ��J�h6�U$͔J�fPS6�-B�2��(�;��ӥR*�UQK�wnq��Yf`�4�BJI2�f�%T�h���Ѷ��I � m���V�X�̐��D�4�-�6 S@Q�X�e U(�p  �%d1(��3PB����Z4��i)R���p PL�U�ڪ��d���a��IQ�D�*��*���,��Ʀ�l�4������A)�3�Ƞ    Sh�J��F��i�&��a��
R�Th#C 0�4 L4�{Jh���4 F@  ��@��� �     T�dm&C$����mL�hf�$i$*�       �D&�lql6(���R	Z�  �`j�rD����RYIGBI Ir0�)�U�x$�"�׋������O����
H�TTH�	*,���V��$�Q���*�¢$ʑǿ.6َ#��ggv>���@I~)5f�i|�r�#��;譔�?*���Y�Uk�5B�,/�~��}�����[;b��#4�z�*4�*���;h�8��`���]F�!V�H�e Y�Q�1`��Eks�D-v���JXp�:@d������P���}ԅ�J�Y����9��0���u�L]/�<�ۤ��36]�nf��K����Ynf�O�M�V�J�"۵o(��^�K��7FUUTw �NĜ:��;R��:襚$�mi��@������Z]��LՕ�	�yM�(��Q%L�7Z�mL/�:�-V�Q��;�U&��rVN�<!�fN$ݧw�LVaą�{Z�h�VQ��1�ڵ�ǩ��X�3Lg6�4\?i�KT�P�Qc�9	��8�^n*mŹz�	O*����-]��fm��/N]���3�n��*�TjG3�7x��� �r{��;M�W�mk[������6C���N�l�L���н�6uV�lQ�(��֍<�b�Ў�rMYY�vзq�
w2��Q�ͯ����aK��w�#BZ��@��UmRbD��rk�t\Yf%3`r�{�pW�:�Nv��`��"@�[�yn��c��9����G����*�6Ze���h�Yp�B��u(��b�Y��a:Ǳ��*n�f�X�L^%7�j�9יW�M�٪����e[.���cEf���:#F3��X5�ʹ)�]���^P�Q̪�T�F�ـ޼x���V�ƋZ��Z� k~�x��tQv�6�ֱH2�7����m�a��է3N��-G�Pj,�t��8��<52�x!��{owA��'/4�Ƥǈ�Vn��k�=K�	V2�]}[Zu��dfֱ���Ź�Ff+Q����j�V�����ZAtb�wB5T��\p��������E��7RG�yl4κ�,�����L�)�h�g��M=��r�i�e5A�{`t�2�~]{v�a�cڨ*�"�B�ïkH�Ӭ,)LjX�T���Vywl]�Bʚ�A�7lc�Č,�x�T�Z���t�����^n�gP�5[������U��h�va��#�����"-6v������0�̅n�nj'r�F/-mɌM�l���A�˺��B�P�����w��U[+tDwX��ڹq&Qn���i4NA��0T�T���G��j�ea�)mV�a�#�L�F������F;Q���a��\ZR��Ok\	��͛1h�-��5s[o-eq��OEޠ��r�Y�Lc{���㝇@����"^Y���F팬���A'n�aI�3WwV�-[
uh�YQ�۵M����Uv�JA�v�{Zʰ�[�t�J��Te�-ތ����Xic5�0�i���ݶUj�e�(�5=N\�{��������SI:�Ԇ�ڋ0D�SZ ��2�o	 v�5����/^���ݭ��(,������f�k�e��E� 3]��X����k�v�炏,�0�M��w���gK/V���l�t�G6��4b����2PW��{Z��EL�I��u4]�&-���_=�p.$��Y����,`�;\'��H}�-�%����u��Uh�����Wa����V�"b0ȱS�Zd2̥b��7l'K[&A{���`�HMYhZ�%C.�0���0ZA����P�BV�KMJ��@ݢ�J��Y�暂�0�<X�%�������5�y�=Gq�q�2�ȽL�02�'s֗u�3RU��hc���k2΍�˫j�b�2}��M�TB_IF[Y�Y��F�Z���Az6�("���zP;�eX�*;N4(U�M��M�:j�;&����区�N��[���n�h=֚��U[!�K�5�GMCa�{���h��ĕ�`ŘT奤�Yq�����4;��D"�aI<�5Q�O�.b�,▰�eb`��f�W�uv��{�Ui�N�ū�Z���͛�V�*��4��Ogj����UNL��x�QԦ%�Қ����mKX�72ӕ�2�fP�N��͔�0�Y���؃�m�!�=&�0-9��##!nK��Yx�vat �j,�y�6��6ê5Wk^T�f��TL܎�+55M��Vjŧ�������iIb���n��-�ffǯ [1�,n�uȼ���O<�e�b�J��c@�j�U��7Pcs���wd�d+HNάJ��;�a�Fཚ%e��>�HԷ_ǳYL�"������hf*�K)�Y�Zr�`o�&�є��0�[N�^̬R �b	Ë�Y�LB���ʘ�hf�u
�v[��`��x��?��+.��5��ߎn��/\52MU�K/]V�tTo��3�v��ݶ�$2��e�J�uQKS���e��(����7Q޽R��Ǭ3��)�2�/2�ک�m:�J��wl�lRB�J�
ۧ�+,n�Kf�+F%FV��QT�l�k�t�i����S�ַ�<,�K��B� of��uk�tya[cA�]�\jb�e�Tel챪�ř�n��gnc��ݱ�Tt�j�T(���6ʬ��J2S5�S�7D�"��6ur��"h:���BTœ6j�ju�v�#�p��nU�M��(WvfkN@���#�<������p��5���Xi�ㅜ�շˬ7w��M�}��=gN���.Q�۬IC6�[��E�ՃV=qe��Յ�/��t�+[�i��Ջ�q;D#BJ�p��w��gj�{x����E��'QffʂQĜ�D��r�0n12�\�Ȳ��,X��`��^^`Z#�4��=c	4�X0�W}�v���rЈ�I���1hH��`�r�ۭT3`g7�ܻծHẠ����Z殐mpƈL��{�����wc��F�e���Ù��8����zN��Y-��YH[�����B�yn�٢����*�Pه,��Us�5����]�UAd�UyJ������v�̊�nT���(�Bhf�7�[Te���J�]��|��޴����ӡ���v+�otmcuf��]��31�"#X6eY{��IuPZ�5�˲�2�9�.��T�5��[	���k����P\��w�7"?J�NM���8���-A����.��D���W[�j���;,<b���m��Hs]lfPY��A۳Kc�� ��ВУo�y	Ȳ�����Yh3d�8��D�i��$�+7��ݥwD�S��\�i'�-Vh4�+f̩H���Y���������T�T��Y����K�3�J��Tmp�{��T�4��Q"`A���#���>�=Ky.�:�(�ɦ�;q�˙�$BQW��+D:��	�(a��s����ga{K�� �g�N�µR<��
ھ˻���C��m���	�\�}��(�X{#+e��(]�)mc5���بf�/�P�S���&�n��hc)YKn��5�����C�۫ݭ� �����dUL���YAC�83�5���:xլ�xu�F�3io7SzC�Ӌ�@֍[6u�\��q��ǽy�v,-θaK��L���֩��I��E�*�ԭ{}y;�J��J��S-�%[��\�f�ތ�zl�)������n^�����Q{�Q��)���`�X�	�ޑ�ݻ��pk�^�C���Ti\�S�zg>X�^�o���tU�6���n�7��S���>�	� wT;��z/���sM*�c�BֻҰ��Yk�r-�]�,�u6m��f�w��b�I`Dڛ�m�Xn�}�^:N03f��j̮��N�K�L�ĕ��H�e��iЫ��`J�R�oz���if�h(Eu���X�R�v�b2 �6��$:��f�b�1�|��R-��]�,���<WL�6B���I�cے�ɓ]��R�d��5݋�3еղn}s�.�3twn]�N���Ƭ��¬�����`=�%4R�W�I]y�͍5�
���b��V]=�{��w�
9��rz���q��rI���v��9�����|GHe�]\��8��&ML�u��S�7�6庆���0��e�r �G|v�յ&P�p��O{�]vJ���7/�f>�$H�ō�%��\�0�%�/��j�0�\!��Q��f����mpb�J��kG	k�n�Q
7���w�P&���*�n���`��N���d�vokY�<a���z��iR������T���,���c4'���	w`9n�0�T�9���(����)Ѥ:̐S��D��9u��\w��F���[Ъ�]gYyͥ�j�IY�:A[��9jP�'çV�n�x��9����YȠ�z��٠�-� �c��%f�>&V����2�d0h	��mG�R��'�/���Ռꬡc3h�����o'�jua�Q2�*���[:�L���-���m�H*-3irc͇6�k�=�!��l��#����Y�y��YR�ɺy��E2L]��N̾�pS;��Yk���o��q�ř�v�n�-�;ng���R`�񓆃��n������)����9n#��2�����Β�L�5��cC�kպO�ŧ S���MC6�\��F��/3X�Y��4#ɍ[���V)h�ZPo^C�<TdL^ݽ9aP\!�I�y����*�B]�sV؃�|)Vj��b���GDu]8�i�����b��e ��mY�Os��ۜ94�^Z��R�@,��p��M�Sܧq
��4�'7F�@��#�'$�}�jӻ��q=��&N	U��H�x�4���]3Qee�9�(s3��dԫu���{	�ݞ�W��;�u��{Z��;�aU8����
R�y�jb���=��Y�}hm� �����4e�@��[W�nAu��å�&�7t��@�wh�ӈ�
��Y�N	G���E�1���\����.��U�7�)`�ո�lX� �}���/�K�c
7LF�8ī����+��e�%_�lr��ԝ�ᱚ�aա��n��T�Ơ���Q�38� �M�N/�䬷m<�Ԝt}�ēp7&.��Ky��[�V3�a:y�V~yZ���`�}�XH� ?5�1��{�3M��i�3Z�����/�BO��8���p���n�싵c�b�W&�����/F�dJߎ-J����)�ү2�+H�}Ж�oV�(�&,�|�;���������g]��a�/�Vqa�Vlc�t8'N����!��@�$G��ԉ�k:�0�¤喙�1�Z�)y[�7��*��a��
�����U��s��.�!]AC!ڀb2�*J�%�ഃ�Q����]È�2T�.��*�R$��́�wc��N��Q����TS8��}�2�#�5�ufZ��/ND�w��h#�ݸKF��om	Ԇ
XD�^�o'f�9��x�n6q�1��n`���ˣ�,�x�R���`�p����=���m���O�P�K��+�q�/*�����^�~��e�{�֖���r:S$� �F5�3���;�V_�8�ݛ_mɯ1�ՁE��݋��zwq*SS��f`*�������d�zOi��Ȑ����{f��.�BeP�p�x�F�`_�!�"�bϮ�J��A�u���v�z�:�T��mn�>�c���Sd�0u�ٛ{M��:�O�5פԨG��ߘ�uܣ�I�k�X���7�ǅX�1��qq�۰��o�2�0�m�6���f4���R��u����\I1���Q\��ܷ��W(zT}�"1fr3�ł����F�t:]�[��b�b�tT�5�sX�|ݣ��}���8�.�W����
��R�:˽Dސ�R��Z]�a���^�{��;pʘ�n���5ê-d�w��,��k2�I+�h�R��E}�U����&Dۢ�w��(��D�Ui*	N�c�plw@v�kU^���$�z1v�i݂�t+m�q�B��w�m1�g-&mӎ]��&�W�Q����o��!un^3WۄoI�m�{���(�y�;0��p.�pC�����C�d5�r�6��1ϣ����W�2�^�&�qQ�nVb�#�Ё-�kw�O��9�N"�8��������dr�!Vc5��ء	0������J%�Qr�Ù��wK��)�nʔeJ��@$rI*I$�I$�I$�I$�I$�I$�I�I$rT����|�Br�}{���f5��jl
�^c��Y��Ond�.�mt�u�v.p̉e�������n���wʣ���%�>�J�q�ξ�#�8�EH�vҚ+���vϵ@����3v�m���zw�+���׺���h*30Cyw�2�z qu�4�"ֻ��W�U,�]L��ֵ4l6�k2	.�c�0l��*���t�k�5zjK8�la��;O>��p�q�.�K��V�f���F$œ�gTוɎ�!��Fn�,�gm�u \��
 ��wA��\�ݙlsxݼZ�fԸK��|�]w$�PI+'�|7rv�"s"E����6 �/V �{��w�RnSx�{b��!զ8禚�i�ǿ��T߭�e�oe�=�/�H�_d5��!!O��xI	��9����R	'K�SS=�ﻚ�n��cz��t*���2���D%jo`I&y�]+�s���nJ�F�,�%��z�O��59e�)ҤKz!�S���8�{�i�U�jO���<y)���r�U]$I]���AWo9\a��65���_R��iB�4��x�*�tV��EK;r�����JVV�,��P�[Be�qM��թq�vj]A�
�Ջ*ѭ(Z+{�4`0^�V����q�&.�vm^,�v���W�8�:Xd;���7�LQR���6�Y�b�v9��4��	��<x3�X(��Z��ڤ��%��@����=[��4gK4�y[�MيU�K�k����"�۸m��m�]��dlh�Y*�9W���s`d�����0�����o#��hۂ �#Zs ǆ�m�B��X��"�]�(UP}W)_5�l���/@䄫�c��w��
���I?X� �p�R.�W��
ٓ�.�'�,�C׽]"�R�;%qN���@V}��ǭ�uS��m4�Y4�N��*蕤�V�.V6����G�,����l��(�>�[��yJ��F]�B����C2 )�rj+�Z��lwu��}�h�����r�cGHG6�pG!��)�)��]�5����]X�٠8��KK�.Տ�7a�wB>I�l���b�9�3kQ�f �FO���םG��_.�L�l��ln�ti`\��of�mΜZ��u���|њ�v�k��Y�i�Cn�+����h�V�� ՠf�iu
���ֵq����C�SD[�Z�#��ݙ�Lg�7*�F�0�w�+�4hh=�����Z����)�j�i���wvQ�=x6t�[��.<B�_�˷���]�NTӇ.�ޕ���Rs}��L��p�t�nav����8ْ��Xa�����c~b���E=�)r*l�G�D���0���<�;�	c&N:�m��jɤ�6E��1�a�H�Y�S�{S��U�c��&�q|��k��OE۾� �t{h������36;}YncX�4,�VNQ�h4�ȣV���,�xO7�>qf���z��,;�R;і]^�ڰh=�y�a��V0M\��r�*����)��rv�
�j�SS��2��NrM�Xx��]���nb��엥^�8!h�.�$��@F@���4��|��{)�buZ��"��F��`p�`$FtVN�]�����I�VF�V+ţP������T�z�$v$)�Z'��}���6����1k�'	Ƕ����N�蕺-ju}�s��.��H���:�"L���B��o���Ϩ]�����H�O0�e�r��=ȱo_:h�����?u��ϯ_1ݛ�so��������2那v ��r���T�,���i���J]mLF�*1A���yV�,&��|�*�61�",9mԬ:*�:7t��e��Zc	X9�6�����Q/z���X�*�I+h��YP�gS�5��\�|�V��M����b�v�T7u�(0([�v�ͫ/Q��t�J�x�Js��?_WAe��Q���)n�xM��e(�l���)u�5��+��zjT�Vǉ�����y��\���a����
�hgRX�cg0T�|�"J����,b��%l+y0+uC�U�c72��vu
��-
����w7u>p����w�7��!�(]�������;�*��J�'~�{՜����-+�r�x
Ke=Ӧ�vѬ���26Y�}�K�YZ,� �ŇMDH�z��l;��JZ2��j�{�/�����c�ؘ=�v��W`-Yc�3
�+��>g�xu��[�2;$>o��,k��vT����u]MY���Y�e�j�r���9P��,�%��q�qRG9p��)�����j3^M����5&>uj\��c���Pӏp۲'Z�f�vvo1{�ZD�D�@�q��o5��u	Xp������"�-�[��O�2cF���]��E5g�d,U��=9�Z�K 9�7wa�r<[�K��,S�t]d������'DȸN1nvd Bwe�W�O��S:V�`�,.8��Y��V�خ?;����ў���BG&-�g�5&V�8gv������`�b9�|��x�e�- c�8��N)D�§u]���lSu[y���Y,欮W�a��Ƀ7�6���l�َSbs�u��DW��s����Q�P��P���v92�'K�W۠��%���U��hJux��N����Z�����%V�pkgAՆ��V��+\��Z:����5J.i��%PG7�^[�tZonA6)�p����rH���a������}tE
]�����1qk� �ɹ��*�\R��Ո�q��R��j۲`7:�D�]I�U֑=��k�ʂ�.��_i����M�1��j�TZ誗]�8��u�5���ϧLo�s�>�6�GG"؄l.=vh�5Ģ)]�鑱v��\zg��9�&ޤ�=b��؛62�K�]-\5������;��N8z�YN��C*Ó/V�LP.�f?��wZE���7"9��ު���m!+B�i
I��m\f��"����[+/tn���Yַ �2muqէrS����Zi�O��
R�`��ͬ[Q�F�.���!���Yո*e����%(v����u�*�VT��jX��ډ���yD�Q��&��q�~)�����y��>�ʻc��%љ�S��҆� ��7z�w��.����*����[� �
}��}�N�jmA0�ܫl�$��WeaF��ҥW���O]v�(��Ѩ*�V���G�7y��(T�;���}�Q8ir�D^����_^�
8���m���8n�U���CJ��\�x�zκK����Ur�8��w�ҭ%���5ad�D�C��j�(;�b⤘����h��a�`�U�1�T�i|���V��ðK��ne|�f'I��O�r�KgN&s��Ј<)Z���n=�[`�OB��,�K�A!1L���j$�"�j��n��s|e��Ԋ�e����O�ҝp�U_3��]��麕o�UFl �
=/�M�3o�t�������
��.����;����urᑧe���T�I)�d;�+4�1{�B$��i�*�Z@vk/�&p���.�������/�;]��qt�η�!źenȭutz�<v*1n�t�T�=y�^�`T�-��R��%�x:^Fq��{+r�v�� $��Q*��ԋ�RK*+������#�@��5�?-�oc�wv#s:oIo.�]
��#Bc�����6ݦ�z;�ά�xe64��w��Şó�W�Y��W3��=����x�x�F�kڤ������)o]�&���=��3���c�$t�O�T�)R�Wm��q���m%����IU�O�AP�q鬪���g_(x�JR4.�;���P��]��-��\_TZ�G��9�N������:��U!�wx������м���wsf����\h�ҹ�Y6<�4u�Ɣt%:]\xµ؝��V�N͑9xT�$�{h	��Ͱa�s���r��쭘��e�����ͮZ����!Y]��:B�da�Q�u�с�+�T+�j\�mmT�D�q�̷�,r��Ɨ-�`�m��������1+�"�X,��W���S�8�	\�� �	+�PY�����R�k+R�Q�K-�e)��o���u׿o����K�F/����/e\�A��EwK��h�Kq}U��e�����*���܂fRDK�\���.:��^sP_$�,X�P�=5�ݾ �bN.�aKJw����iޢ
H��b����ĝ�R�D�@�w��-|0�(��=������-�� Y�4n��g�^)/Jc!�5�����=�t�ث�*ǌ]���E<ǔ�zzRŕW���P��M�vɾ�A�n�{ؒ�8�n�{�?=�t��#��7�
�	W���H[|�`�Ok�v����-n��8��'�>��*u��d{�0��)���s6��׹10��*o��U�zz[�Wn�m����Z�7Y7q�ݾe�'��3k��|l�>u��_h���/H�U.;o�n?E,t����1��	��h������4�2��(>x����SZ�j��Y����9��'|	~�P=w�-\uni�Źܝ�v���hz������-��;��B� �SR:8���s��Q>W�3�)ϡ�	���03ST���&p������W�����{n'����S��R`Ր����L}�3�y���E��{`f��Ubat�|�gtNsd�]�*zyN�v�v *ۨdVLl���Sj���}x���<(�p-�'�u�|9�P.����o��%�u�A7���o*�5w95t4�P�
0������Q��B�SΥ� �y�sp������מR�^�ɲ��z)��GV�}����_'R��K�bk3��/�Hx������8�>8��#_��r��d&�{H^[[�]��xA�������Fl(*�P��	�v�ƫ
��i����k:�t��}����(m��)�;$������K�Y�}CGy��ާ�Wx���uϥ�z̷�A����.��I��[D6g�r�	�o���ҥq��x��%��Sm��yfi6s$.�'�y9�}��/m�E��3fv����R��ޜ$Wk�Չn�3�wP�o%���z`x�����vc������ch����ˮK��-r߰�� ��s3`"H��豱�K4�9
M��y��s܇sa2M���]E�髾�6����#]}�]�ky�D�"�l����3��s8x���gN4<�Ϯ��aI^-M�\�v�Fܼ0/^�Ƕ�>�r)���}ѷ�r�\oPcT��T9�n��-���4��8�'��x1\cHq�HZՄ�[˸ꒇv��y5˅��ʬ}!4��*�6l�-���6���:͒�9��v�G+�n�뺝E���Y�]�s���솔���3����,i<X6��l��źS�5�`j�!�<�kV�qLRG��r���B�]Rd��5��ra��I��hx�t���P�����ۮg��h#x�#��Jj�����dc�[{9�w���@�d�o&݆G��c����g��t���skْ����[j�hroF��ϲp]��ѲRO-U�1e�s������mqv�����MLy7�����v�r
�uv��G��1�Ox�M�ᯩu�=��0/�Ưs��s��Jʣ��%��K�ɹ���p=�1P9�'�ު�,m���wUNb���c�h�藆��P�̌`9�7[ܮs�gR�����3BNn0�V�d\�-��}���KJ��Vq�r/`��·X�s�^�MC���輩���{İr��箹�5h���E�/4%����]��M�O����sewGIN��G�en�����Dw��
����U>��ɦk=� ӄ�����u�;�w��$�ͩ��c=�oc�$a�k&����t����9������q̻��
E.��lS���o{<3���mt�W�y3�0(�Ѭ�EO�dCy�`�P�%�4���o��=�>�V����?{~{XuuH����z�0\��i��(��E]C{bamd�g�|��o�+L{BWLW�T�q9�''v�C��tEj�7Z�i���B�q�ݷw�z�n�Kk��G��j�	�{4Z��[�x��#J��\R���񽪒��N�۝�̩�bu�[�Ǻ-� �bp�p�m�Nzi���ڡ^�K G��G�ۖ��V9����;b���2���gH�'N�p�����aӮ��}�9-*��'��<��"�lsn!*e��w��Z֫��h���K���S�ǳ+)\:j�`������a�i�4�Z�h�(ݖh��O��=�)�{\�@����i2�Wvއ�eX��Y�y�T*u����A>�VDL��{ܺG�(��z��M	������߀������l�rnG���2�<Ub�g���*y����k�wq%��&0��9C��z���&�z�PW¦Z��ʩ�Z�Ҫh�"��"D�(.��|�-C`�rqiJU�Y����/hs�B=�������Sw˔̎��4]br���1���h�3�&5EX�"��:z��>�5�(��Z��y�c�x`n���eFe�9����5��EWJ��~�O7^��Ԓ����צ^k�@f�z�W4��mdC�8���S�:����	�^Y�V�U�Yƺ�[��_���U��{Uf�ln�}C����G���f1~�<[���,�LʛL3(�X{��&�Wkct
�Ң�OQ�yn�VXh�w��Kzվ7�[�:͹�iT���Ͷ3Y��\6Z��RY]]�a%p5
�����\�df��V�i]��F�u$Ãm\���D���u+r4��Y�qK�.�{���L^uә\C��G��S�Qʌׁ4�����݃��M%�O&G�B�+8!��MN�dl�@��]�q.��(��BVZMl��a��K9_Χ��^�Êf���=�h�q��q�XwW�GI�xm;@���0s5:�r�Ħԕ�D���;�;�7y�0���PUE�s�ݚ㈤uc��pM"���hj�Wq��)[R��[�2������%���_�D����~q8��'>5'M��Rf���ȗ;r�reJ�$]7��j�<��p���Z3���I�U�+m���%�1CcRryK�#�e�%��_hHcܹ�e1/�V�o�����*\&�bV��qt�,含i���҄%�>s�Y�vڦ��  aη2�d���^:8���.�{�����&�-�V�V�D+!��Bβ�t[��@�B�Suy�a zx3N��Ć�i��37����ԮHs@)����l!�ᏕД/w�#��4*�|uE}���bNȥ2@��;:F�� �P���WZo:�%;�5�F�Qj�;�}���ׯ������,t�[q��ZU��Ӌ[4�`�GV��)��mEq�6�)�+ke1�����(�4TQV(Zk-�X��H�RWU0��Z�#V1�b*��Xň���V)�����F,T4��� �(9j+�"�.�(1Q����`���k�_�߫�RUs�],���qE��.�o%�m��Ԟ����3k��Ydui[�R?����QE֦/)������D{�1��_��c����T|�A[(mB�
�ܹ'�/��Ǭ��D��V��V,Bf3�A��C�f&w����m=.ϯ`�O`���{u#63�$:kF���4֭q�a<����\C��5O.���hh�;����l���rq�,�w������Y�OhW����Ay��@�)4��p��`堸^�1���9�qvQ) M���c���sڸ�]*�L�e�6�Z}�<}^�o~}z����z��C�D롖��<gV5����c��FU@�Ƀ�9��m�9Є�uo]ػ7[���鯽���ۡ���L)�ж�67RR�����s�1�g���m�uJ�U��Ί�-�^0��A��zfq�G����c`�_�<b�&C��Z*��}��-�?&�OB�VCr�����Wi%{ʸ=T��*��%k�]��u�u�3,fjcB���ע>�lNm�[p�Qʨ���'p��i*r�� �˒M���˼�T��M��6�>��馊Z�Ŭ^�W���O��өS��9OoϹy�]�V�������p�mY2�7�ۏ����(t+�H*"r����r��+���2E��yߑ��Ǒcy�P>H�s���%!�� �ϝ
��j���?@������K��$�QΞ�%��f:����9�%:�fŜ�Ѥb=	mH��s�
�I�OBX�ژ%�N/�����>�	�a���Wi��A���$mSP�SI�=$E����p�
s�M�;��3M+��˫���x^q����2n��u}�g�ڼ����+F���珞�Q�2��ɮ�y1��Sѭ���c�mj�a^��隗�݅n9EU�d�4q��w����06��6=��z����C�ה'��j���z�~k޶�3���>d>���3�)�|�q�ć�'�&�6��m�{�I�� x�Mm����9�����!�Xq	�M�4����>C�`wO�C�bM�!���Đ�}��7���p�8����q��$)��H�d=|�'Hqr��=`(L���{�Ǽ��ߞ|&~qjb>���kF�ugի��X�b�15��7Xh����l�R�vog����ղ���c�O.�Q;��������}k{��x�M0�'�'�iI�t��	�*@��'Hz��T��n�&��m�8x�o5�:�����o�I��>0�������2�q	�CHN�q������Hi;@��:I<d�|����1��ca���x�4������}�ﯷ�~{�q'�>;�Xm�xöHvr�=zd�'L��H`����XM���z�~�������C���8r����Y�>a�m�;���y�����	�C*���5���߾� T1��l!��%d�52��6��!��O;@��	����0�@�=�|�[�k�x��i��-$������tn�
e m�P�$�2C�oL!XBx�ǝ�}��s�;Ld�$�P���|�v���P���P���Y!y`=!��<a>̽w�^�����l!�N��	P�Y'�l�$+'l��I8��a<d�h��`��!��=zߙ���g�L8yI��	�G�$�2��N�!�I+���OY�ğ{����˅ԿQ�1.���!~-Z����0e���:의��jdr#�i�e֣��vn��ꜵ����I����_wq��/�@�>�H�}�'�I�rɶI�وC=�P�!�k����<I�	:@����U���}�4�t���
e�� k��C5v�*VIVm!�C_XI=H)6�P�{׻���w���|��d�hC�hM�j��9`i�d5� |�ěd�:�B}`m��~�޹�<����� VO�&�)�&$�`(v�|���'Ox�VCɪI�8Ì�N������sg��ߔ4ä�B�%������I��BO:�<a0Ն$ݓ�8�{��W���|�߾�@��������v��I�z������M%M{d��wϼ��k~{�i!��КBt��;aR�t��6��$��$�2N��3���o���o{�C�o�L��RL����6�l:;�=a>@;a:@;������﮹���}��8�x�wI1���C�|����ĝ��I�o�8�3��zkg��B��x���u^7�x6@��0���
q�>J�>jÉ��6�L��LN!���2�',���U���,=y���7��Y �y�cA���}Y�&�����7wM��*�/@�-��A��������ē���0�$�3,�����i0���:I�u��R�C�@���}�|���Ϸ���W�i'�:Ձē>����M	 �d<Bc=C���0�ӿ�C�<���=�^k�<�ô$@�`x�|�!�d�>a6�j�cz����t�cޟ�#�G�բ�wд��v������L�d>f�'���$;O��`|��'~P���Cl����s�^k���ԛ@9:��@�XOX0� w� �!3T����'bV�}`m!�k��N��~��z��y ě`,'̞�I��Hu��$���4�qO���T�!���<�Y�������	���$���@�l!��!�!�6�6���O�A��{��5�w�7)�t��8�Y'm��H>Y=a'�['����(|��'�k����̈́�!êI�V�������s�V/Wr�)�ݦ����R��J*�x ����N�_'f)o[~,���:1)t�d��|1�/f�ݕ�]o%���b��ϳ�%�\�w�$r?��Vf���VGdP=s�#�+z��ڱ���\�f�+C�#Y���I����'��yk����_�!�v��{od��a�p����ѥ��|��@���xp��#Q<�p+�8�X{J�ݠE-��L�@M�|N��tlL˩�r���:��[ʉ�vWշ�gGNPY�х��z݌ɡ:鼧�*{��)Z��lo�LN��4&q�n'5&H}O��mR�Y'3F�I��W_�_��H����\��TjJ瘍��_$k�b�D�?���	QJ?�]�=K���x���Q]5߻�!05(s[Re*x��x���f��s���&{�T�� �kN�e���f[�Ѽ�@JNf>��w /��Cg����5~��t�}�n�Q���I�/ju���Q�0����u�LO��&����F����8�ϲ�A7��U�YZ=��+z�/�,��˓R��(�	uQY>���e�4�(U��^���ۇ�:�X��J"�����3IA�^�-���˘Ԣ^���,m�e�r��b�4R�-�?�}��\L�1�/\Ƌ���h	[[*�ד��9�\�yj� i{+%E��x�d���M�������X��v�C�xL��{Ϊ�Xm���.��MeVg�\Zz�ʗ���h��ݽxR�V����/��,�V'b
��j�u�Dk5���s��Jg��.T�������HÃ���2f݉�΄�݇�s�����=��G��SI��X��\�yn�x�J�t1��Ca� n�_����{���.Bt1nn\��/r�,������\����fMtn�e��؞�-(��A�o��&sZ7��ު�S9��semhQ�+6�Z���om�-g�_);���Y��D�F�R�3�%� �Zszv>�[��#Oge�������W ]���	lr��MB6�֙8e��4�C&�\�ɓ7�����͌�tN���>��B7���	t�X�\�:�7����yy�:iӯ�R���+��7�x��+�ё�%C_U^ �2��ۥ�۵����t���j�6��wӊ�ww��C�uoLs�W�J|K�y��l���d��5�*�>���A.���I
�jj6�H�Y̥��%e�ʾW��x_�����~�0nSgT ��,�Lc�b�ɗ{����U�噏��[6�p�چ��+�N[��jJ�]�O�ur�M��ɿ,��KC:�R됎yv�E>T��3���s�޴��c�L��B�v��)u�����ӓљeD�t�J�1[Sj\��m�aO0��-�Y�UÖ��eNs����9��'|"Pq��;���%He�hn�|^Ą�d���|�T[ƺ��{X�>�f�4y7Nm4�.Rv���������*|>�طd+R�o��P}vJX�n	��P��i�$d��G.NqQA^��� ��!v7[�d؅�Wk����i����x~�O��U�E>j֨���"�
��ֈ����A�� ����PX,QDDVEE���TPUuCHcX�DA�:ZJ��,QQX�Ib��*ňȠ�*�jȰ$+�V�*���������������5�?�F9"����[VaJ�l|�Ϋ��s�}�}��5���~m����f!B�?�z���Nf����v��d�Ve�{\�P�S�Ctбe"ѵ��pl�X��S���y<Z�4�	��[����j�R��)�G7���}�y^�S�j�a�ʋ.��:-��m�PU�<����+t�ȃs+9=��~5�E/�~��WOcr2Léݥ�[���^g����4p�E�o�81����=�ސЇYY�Q�Y���d�b/�;�S=S[��ꩫ$`�Ϝ�o�	�4��։)�U�޾����Յ����w������"�WDh���w��*o�oM�@��k�w�
�'������&m��.R���f��uؚɧ5���}._P@' rz���:q:���w<��Z���a��/D�[���hno��y��uc�־��B��ғ����j���fq���=��aև������o�
�Ie��k�}k>�S�������''���:ۿJ��R���c�C��G2B��?�2��{��;�Ì��C����ż+U	ξ).&��%��{�S�oU?��f�`�u��x�� Df�y����F��=��{d�IJ����ћ�Hy]bej�暴��iOF��Z|'j�Ü�2��7sU.�s�z����h��7;g#yCx�gT�����GGokViNZy�����I�ˍ�xv��T��Y�����7�5]*=�'nng���Y�ϝ�ﷆn.b�����O�)�E����3a +�v�k�(W��3=�N��h<�YmKզ
��h�ܮ�|�Gy�4�K�^���Sh�M�Lk͙*���~ =� *�KR��*/�{&7�r����i������..޺�����&�gݸ�{;�c��V�UЮ(���G��<;Y2�}����3eV��n�x�щ�s*uV��s��d��;t���;�4���ɐ��m��&}e�
?|�M:�1��-�e4�b��Y6�f8ݺck���ۛم`���%�eǴ̴gb�햻7C�$�����c���B��=���,��|���x�75Ǔ�a6�ˁf��T�%�:ʅV�����W��'~�����&�o��!��?M��.�l������r�6E�a��8��h�Z������n�2���ͩ�����G鳙|�hL1������N�������Q�N�p�#G�{	�G�(�k|��D<:����;,�Lʳ�v*��=�8J*wp�� Ψ+!��{�_���O�p#ܟ�6���a���+.gH������26���QF'�]�{%Z�E��U{��'�����Xma�+sY�z��i���M�;2a�A+;��ť��̽�9%����5Mf���g��gEbꓳ�X�'����Ls
+��Z�3x�6�빆���i��Ȯ�ǒׇ�9R˶g(s"���'�)�v�J���kWi�sYϞ�W��+AŅd�'ڵ�i��1����~>�l�u^����2�"���7(*��&�5h�+��*�u�����+V�i��)~v��@�^!^��ζ�+������3�׉� R�y�٩�0iE6��cy��vY��U���#�4̤���=\1�nY썌v�[A)?}_UW�TУ�JG�خ�˿�6����g�ĚRqL�ޮ��[�]=�6);Սf��XZ�7�7��{�W�����ן��g�nQ�F\ƒ��8�\���>RW�ٱ�^����_U�t�n�Oq��������<��5�(��Έ��T�ߓ�N������΋y��bP����j�S�msV�gzlƮ�A��7,{�k��zuA����=�<���	��w��w4we�ԩr���xR�˯:6,�\P�:|�\���r U-Ծ������j�nˌ��/�֙�<	o��y+r��Vs�dC�c(5W��)��]y��U5�����eumUA}ek���Q��6��s��O���me�m�yU��L��Zy	��6ltp�۾��7�4XJm>ܹ+�	��E�_��=�k'�ѐ����򜶐����z�m�Nx�vI��j=+�'�G��C=�w%s�;ʒ�4�E���e��d��U.��b7/��ʐV(����v���ɏ�a�2�Wv��;J#��r_� �ķQ����c����,@k��4M�6�-��|��>q�ۢ�
��-��E����4woU�B*Y�����V(���=�`UK�N����n#x�r�/������ku�션G0�sdLE���,���}oq�S�^�8�����;�+������q$y����0��s��ݢ�������c�l{s�Ga�^�*�SZ��U��AV9E����t�3�޺F��^ő�%��gc�C�ҁفm%�i�jD+��ȗU��B]��L��/���𚤗t_�]�3^�b��,�ڤ���ۀ���e�3j��:�?�l��\=�\���8S��U޲}Ea���~���8�&�?�����8������J�"s����$�q�t�Z�̐�\��	v��k�t�I�j���� �K��>�5���Q]���{d�#����9c�̸@�Z��ػr�oTnV[��U����׵�g�NU�B+V�����B�{�L#ޫ�u<Q�On�U%�Gna���X{�:h=�����C%��\�Ӎa����Ǟ�0d�N�J�Z�����ڕNn���+Q;��#%���Xb�'��ޚ�7�~��ݘ�k�(�+5��������^��St�� ��]�(�L���rRb������Xe����v���3�7�a}�g|��sh޴���e�r�욵dN	0_0����R�{*��I��-`Ʉ�t.'�Z�����%���y'��*EJê�)�u�9�3�{�Z�飺�N�� ���R�p�]��IY�y^Б�{��	Y��TL
s)2ﺈ�Q�t�>)��$��\��m=�ij���%�z,J�\�,�y��6�b��G(gS�x9�\p���8}�2@O+yY�u���Y��!W����%�-�Y��[�opK��ٜK컯�4\ɊX�*���LE�63�eۜ.e共��ʔ��n�m���������u���t����8�h�A\/v�ws���ܶ�����A*&���]lsyr� ����>��u+��XyU��n����tNwl��: ���9�ի���������zP�=#��i� ���t�Lc4�%�N��wi�Bζ"���]s�)ZU�su��#UƮ��Pi@������FG&�9O`�sPC#F�Ԃ�?�.ү	P˭Uq�*�YŻ���V�c�� ���dP�*
�,��X��AAb0D"��(��`����UƊ��TUk
��X�E��@Q`�TXT��"*0QdR
�Ula1��J��U�E�
�P�T�`��"+��HQ$�"�Y��$�dU"�BT�(� �3X#"�X�,�x�u���>�{�ֻ�f����h*"\��AN��1^�#s�}U_}T�nF���o�2�^ǟ�$��z��ٗ��_�,xf�k|��qw����ҷ�׽c;Lx#p��������Q!uk���r�>j��'�,�@�Lm�]ՏkCw������h����m�l[<��֫Xi��˻�w�fy������q��]\k/]r���pB�ﭽ/�C3���p��μkF���<ǆ�YO�A.��$^�<k�7o�^R�+[�g+���:�s�>�^x��M�W��%(�*�L�v�VpĻ������KW}Y�|l�6=v���u�d��s��dCM^�_L����ٚ[�֪w�CB�S+��t)oH����{^���s^X7��NRo�?7=@����o�����;��妛�et��z"����{�Z�.�X<�+�m��R� tc��}W�]3<��g��<��(�}�I��S||{��3RE�k.VkR��&�Mq�7j{͞r�I��`q�Eu��`�5������M�^s������;&�%�Ȁ�@yv3۽N9�l>�I;rظ��}��<?W۟g��g�w��f��"mK�컍M�ɼZ�yf#3dFr9��T����������Dmd��"���5�=�=V����P�H`��"��X���-Ԃ�qu{��X[��b{�D������;�w�������$����tw,؞Ӛ��àTVgc��ȇ�g))2�5��(ns=�K�و��'#�@�=^u��Ee9U����-��Y�C��܆#��حxx��=�<=`��[��T]��\�S"<Í�[�\�-,����I?�U}�Q�S���td����㸼���.�0I.�дT�X��-�Z�Dv�U�ىpbS[q]���V�R{"t��uTۣ4�kS��ͣ5j*1�h��y0��x�;��ҧR���P��^��94I�w�kYG���e��ë[�N6�b{2����n[��p�{���Rb�����	9����&��U�f.!�E�ϵ�1k�i��@���p�U����v�����%^�߼pQ�z�훒�0H��:�^V�����g%:U��7���xoR��yo;�ßA���ݪw���A#�l��*<��������S�\gzJ�tB��V��L2�R������r�M7��n�J]i�I����cy�2��h�n�#Zd[n��\0l1���z���oQ�ybe
Vd�*��u���<�;�����\�mK8崶FN��$���g��&e
��C�^^E���ʄ����"�-��I�5^�W���mfF��(�8/���:���}_U��#W�����[.�E\��4��¬>�S�N�>ǂ�����@��lf�@�t��5�x^��=38�h����K+J|�JFt�����E,��#÷^F�7u�ґg�;�[�G푻w;�V�[��|��H/U2�T��"��%m���Ks�D���1��:�{��)��&��Ɉ�"��tM���dW*&&�
z�%J���ɧ��O��ms�{L�<�j�R�h;�H��s��37�����#O������>�l�|�s�}�W͇��k�c�w�V~����[p{���=\rf���w��� I2�^�5����(��=�p-���u�e��ns"�f�k�g�е��Ѥ���yYz�d��@�r@�q�h���c`�8Q��;q�!�G۾�<F���E������k*��)3����lb�����?a�fϮ1i�C5;�Tu��B�;ǰ#|�kV��m_z�ҽ���Z��;��,��バ�>>(����}�F��I���&@yl��A�z;v�!�.��������[3�z^�D��A�֡}�k\�R[e�'ﾯ�,"l�=�0n��*c*$d�|����<�.y#ꌆH��f�4񢗭w^�W��5a���$����AUyV��>+m�i�ɝ���GNX�0�i-|0�/��*>��Q�闾ϸM�J7�@U�ltzat�g=^&��\�n즹!ǎ���Q1���"�5�����3w��ɕ�xIq�B����b#]��J�`�~"�tX?��1�ᘴ�t���{Y'M�x8�P�ȳ����B)!{��x�L�ۺ��dl��
'O#�FD@|��������qs]��u ���8Tܒ`'�݌ںq:����V����T�Ț0�ê� ���m�Ţ�p������dF(�߇�n��E���Xh���oO�u-Z�^m���H�^a���-ʘj/�Ej�i��c^5�ѽQ�PX ��6H|d�QQ�o�HgQQ��X{�wkw;Ly�s�$�v��6���,��(�+�}���a�6E�\���l;ZSo��������Mͱ~C��8���5�� ��>��{s���^�i�@����qcB�m$~e�����U�E���x�U\�8A��$��dg�y+�.�Ө��Ӛ�E�c`�ȅ����<_Һӻ�m5[�ai����!#�4Y�C�`�=��.��p�;���{�l)��.bы�u�E��.k�ƽ쬓|��5A��S8@�u���������~������E�?� �j���?������ξ"h����g��DC����H�2F|��7գ�z"jr:��P�8�Z}p3���B�q����Ƒ����UHq�-7�B6��j�����^�p�z��טԅ���#Hf��(�/b#
�~�c�}������������f������9aL�) ��p�l���$�{N�o�2����z�o��$h�YG�����D�7�����y�E"�(��XB�,�0rҦ�Ǖ�/;8i�;���g������vz����0O�vS.�v��Yܝ*��{�WaS�]j-H�νz�ԼV�&�JYal��W0�En�v�&K����{F^�Ba�ur���(�O�DI�D��\ ���eN����j�RRh^rbvm"������z��X��nI�;�iV�&E�뷤��Ы׻�)�_ H��ܳ�R��WWj&�[����	JH�4�K{��z�W��ڙMׂ'M�ݲ�u���331��,��UFDm|��JZ�pk�Z�Y���`W;/%��p�I��˹l�t�ڪ�A��̀��^���u��4����[����I�=N�s�H�u�zgnHr�PD���`�����}ik�����Ou�;��f�>�׮���H�H��]X������|6�i͵�9 ;�Y]hge��EJ��켱���oO���4�Fdܚ�_M��#GtD������Ol����U�4M�ȢoN�6R��LÜp}va�9��y���l�ʼJ|�<�Z܀]�4]��OK;fN����}QStgUE{��}�3�2����p�B�2֜jF�	,��R�+;�U�܂w ���[�+��K�2�T��c,Q}��_����\d��#�[J���KR�:�f@�X'r�%㩭�"�-��S��Mǹ"�^�3�CڦO-�r�+8,�m�mJ�o~��מw��w�OGm�~��3�"�����$PF(� *�HUDB,X�P��$%AE�*��R�"�"*E4�a�X�I�Y��������,q��$��Ad��4���D`��$��PR����QH����i��� �T�t��<�����sx�{���������k�>er�5k�/���
�_4�cc$���#�9q"Ȇ[#	�i����ܕP�8X?u�-���&�kP(Sj���Ng���i�}<zy��>�qp��p�=Ή�6վ��0����Db_LşV�).�Z���f�8�����:ƿ��Bx��?R˷���DHK�!�H�+�q�־�Ŏ���5yN��8� �21�r������~�x�N�/�t��#-Y踸��4t�W�1+���8�z��5dx Ů/��)�$���h��.��H#��0��d;��hHk�gL~b}sߗ귖��3Sﺸ܏�a�)	�ڢ�,���F�� �;�x�86k��U�N�A}�k%ot�.�!�/�}U�wnuq�A:�q���X����B��3��V߳~�����ƴ����ńY��o+U]]{�!���5�4���������ӧJt�����r���[�'���C�B�a��g�<��k��&{8H���4E) 4ݣ�z����cͽ�yһ�Il��/�R���arq�f�	���^�H�cC�
3�B�#��D8Jv6�:2������'j|~�/ek�Ia|H��S�/w��Wmq�[��<8QȄ�Z'�i��gd��fn^�>��"F�K��#"s�C�K\t��'�׌��v7��;٫e��x�9��q��� �}І6K)t[�i�gY���7��j�r\a^�������Kz��d���y¦�Μ�c�b�����zx���:�+<@%�M!ذ�^#)i>��]�d�ik�C�ȣx�����/���]L�xԨ�}=,�e@�q8y."�	9a\��[���íbd�W�z��Y�GF���Hrb�3��z�3�Y�H�1��C�����/�i�vA��]ü�F�ņGD�����=���gڃ�8�?_-��2֖Q�5}	>o�$7Q1��Μ��y,md���V�������لdt�ؐ��=i���@�qr�!�t��A�8���Q����b�[v͹��ܩ��ݬ��5�!;y��mj�r�,�Yl��s���M����r�+g��Mf2������S?�֯�ݕ���:'�Q�:"<0>�WS}��!���c��P�`� �1da&���ʩ������U�A�X�(G���#�r�\갇
�$�!K�2�45�=��Y��e__�������?Q���G�c�%5�ӗ��D_$aé�UC���6��̘^R�i q��؉7	�>�T8.t��NjKI9�˦"�Hޑ":�3b�Q)=3�B���{6�_m�(�Gq��8��S�=�d(gl�ldor�i�=t}F�"���H�}��?!����O��S��d�
{�G�q�{2[�P��	:=���^sJ7�/��r�1*�g'�[J��5�Wm�����2k����\DG������D���Z�W�|3���>�R;����2�3��4�g�tZu~����a���:t,��ư�16wH�ҕ��]�d�υ!�45O�#�
C�
B���W��u���|I�5�t���Q1K��z���$��_Q�P��>b�x�5����s7~��z���0����H�G��Dϫ��z���R������F�ƚaS����=���"��txr���LD��c��ƈ��qs��m�p���"$�Qԋ2���Ǣ��ˍ��^�k}�T�y:eռKq>
�*K4�dSw��a��',;����f��B�s;�|����C�O�}�vڶG�DdD}�썅
 �w�����}~t�V�]������B�#�<.�����z&=��R���a�ǅ��8��;H1���j��=��@��G����i�h����wkt�¬���d�;��k���G����,��ݴ=�w]�+���?���v��9�e����$��3uq�C9�|G�1�eRxC_x�$F������
Ο��c�>��5凌B����"�*�sҍ�~\GU�!��IG�|�>>��5���4��"F�����8k����34|�Hae����h)JFfZ���� 6�R���oF�|F��1#Wkn��kx��3�9]ɛ�T"U����H�7����v�v�Q��$���q�(�"�F�y�����o��)��̼��!�Jң��1l��6F>������l�����b!5V���=0�%g���{ҧ�mh�ʒ4p���Fe1������y�˔��ҍ�'�`�(N�ә�q�gR�}c��m�o�ΐ. d�`�	fA#��N�A�H��OB{O{wg�D��C��6p��;0�RB��5߮^g��d�%d9r�d8���nq	W�/�"��G�4-��i�ش�Kix�8a�)f�郍e(�$B�a!�O?u�;��@�7���)���ev(F�HjeA�5K����0v�M)V�LXνGK�=��Kj�*a%(��Y��'?P$o�n~��ڰ��??!�v�C,ٽ�#�U����F�Y�L�څ h��\i!�k%����k��h�.hm����x��"j��,�T�L;&���L]�Yh�4��Ƒ�A�9��ng�,�zxy|����<t���4�����{r����<��4<��5��U�� Ut	�76���[8��:~�a�/���D2���DD���y�a�>�p�`�)ȫ3�<0�C͎�|�]�:l@��|���T@�����\6��o�����_=2��H�@u.��g���A�]Vˣl�*��m����e�)�_�%f�T���v�hn��.��w �[�;r*������nE���"�~�ޛ��@2��儸��/�_>3�++��B�˼��c�@���� �#P:;Qh��7*μs�T�H��N��@�9

�i�ƫK�`2' �eY�!�H��v�6�<2+��N�Ke��q��d�#��gbds"\�3;��Y2jTgő�:f&�2C��N�c�eK�p)^/&�M�ӎ�_��>'G��͚�^�s��ʉ$t8�(�>Q��R$T(
On]=�v�'^|b >G�d�����ɏy�-�A��X�fo�TG�<|<���U�.N����5�zc���^������� uc�E٘�m:ڪM\���o�R��4�=꽘��vi��Ff�H�8�Q9��E�j�+o���0���<���G)�^=����Z�=;/ٞ4Fw=6|Ez>q�1|)�dş[w����_�7�22����}�I�;z��V�~��6}����C�xCH8Ơg�j*�kl��j3#)}ĝ$�1�r��'-<��ƶ�eoyo�87�=,�6y�qi��t�����Uf������)ĺC���a���s��S��ߙ���Bv��*՘QsU$2f�lE��qG��t����������k�m�'h��S=�󽱒F�?���3�ځ9~va�X�cg��ȫ��ߴ�(Cڅ;�ڥ�9%w�;V�s9��<CY��T�D�7M��?�����vb�ͨ��ݼ'�<�٬X��Ȳ�e��N�F�2n�KA��`�K�N�-4����A/�#�`���u@�ު4��/���5�j��������i�+�
�,�=�.�Vﳎ>��i�uif�'���,z�ʴ���\+���v�F) �J�o�;[C�T)��-j7��2�X��%B�V#�{'�%@����t��ٮk\�����ɕ��ʸN�n�|�>�d[�v��|�>��5�*�1�Y|��6	��~�{�l�������9=�`��4���³���-�Pdq���I<U�R�*L:�^��w��Z�qd�6�~�w�x;�}`Ѣ+��RMpY�4G�:nr�|�%N�
�C
 �.���)�
W;땹}��h�7�_azuZN�=�vԕ��gy׭1��A9$
w�"�v�j��:��a��^�'� v=07Zr�������S���q7���Q���,��ev^� �xY�R��.��3�Xl˽EfV�2���r�t�z��L��II���jY-ʺ'S�ǥ\�,����[ݕ�5�rߴLv{E�t�!��$O�wg[Nt����v�2<���^L��قm����"�dq˛���q����l뫳�w��C����P��!+�Y"�$�DC#+�E��I
�*IRA��AM$+C�(Q K�AF�Vդ����%Q���Z$�)��IP	Xc������!
����!�
*�%@��L��d�$Lq Dxz"b ���݃��/oۮ��ܾ����K�79CX��r$���v߼<����zg��Jq��y��F�t��YN[�f����l#�����K�>���<���!c�2���.٢��ؾ�D�j�`ZҒ��|��\��ٻ��F�;m��"F�:h��������[���f��@Q�m��KN<oQ<�Aj��-��w�iG���}/u�;F�'WČ6nyu�����N�'[0�E���ʶK���W���tb���#Ǝ����4��E�}�~�#�C�D�dq4�X�>9�����v{<�QCñ�EZ �f:���U��u�������%��r�ʲ�w;�[Cx��j_4�+��U�3jX[��>6P�%XI��*�wy}�Yڙ������r���H���U��E��}ȅ�>8b{=d&\\V�G��+շk���vǩi��i�й�W.;)�!GiW��{�n���
�(bX�.2��Ar%��.���m��-me�vz�&|��Ӈ��A��Ƈj$C�<;��{>����/3��}k���d�\uÞ��W^�c�� �r&�@� �>�##���<�kk����>1�\
"�i�1�haZ�lM�w~��YD���Ql��Cs�!F��
�fP�q��B8���EՆr<��rޑ�M�S�ʵ��J��zd9ɼ��7�����N%^��mC�`l^��J�vI�S�n.݊�E���^���{����˸lG�#�@�������K#��F�q���w����2*z<0�$4r.�j5CDk��;�E���A�~1�a�k�
j������oU���N�Ӗ��6] :�j�!��z���o��0��@-Hq�n>�R��NB=[x�7��D)&$8��I�5dt$z3H�fAt뷴9?C(�yc����H�]��y�ާ���C�z��}1}�Vx�2����dy��/ظ��)����	�i���5��-��Pg��"�>#�}A�5��dB�v]��0i�W��H�x��Z,��²�v�ntzq�_8�Ou�Wz�<�̅�#-����{�M/�*��I���=��h��ۣ ���d066=]Kq�K�q��$�Z�A�j��釘~\y�|�]��Y��t��i=L_/������6���ݗ��ѥ�a&����1�������۱��V�"�L�:t��c���\pI�+�p�ۧ�-���(J{r����b���{����	�*.���}�b7���΂~��W��8��Bm;"�a�D��H�u�x��b����J�]}�W��a'Ě��^\Y��1h{�q���7��ُᑿ���$�Ň>���g�L��
�X��]MH���1�Չ,�R�+�ՌY�OshV>So:�}�n���6_7�Rs*3�������f��S���\�=��~�2�~AҟR:B�����|���nm�ިI�_/��s�E��?U�6T�Y�*4�=��C���:B���Șg�1�8����F0����{/gx%������=zb�_v�֜�veV㶕��q�Pq,���ț��y�ݜ�7ϕ�0=*%�c"���!�|p��Q��TV^�zq��L���F�U�!�Ғ��;�x^�׻�Ԭ�^6��H�x��/Ζ�k]����߷,xD��#K�Ey|p�./Q<�>�g8<cj���a��*�G�
5G'�Ţ,3�|@�m��J���xv�Ʊŗ�ئ���QZJ�eznY��U�k���M�c����]��g6�[дuEZ��V<oz��G�a�_~u�Y��3{]g��7o[��<U����#�)a�q�e�p�<�ٞ�,����"	����
��<r���{�x�-991~@K@���>1���F�{Qו�k�w��\(���DS��C�ȣx�R����ݕ�ߒ��"��*.���
27����Up�n�|F!�#J"��;�ȇbM_):f�{�r��!�6��n$Di�e���|�K���ziȑ�bC#�Aő���UrsM,X.=k��c�9qș�f��4I��$����^�p�����/��8
[[�﷦-��WX(��ٖ=��l�h*�R"(��vȤ��u���x8�'��V�Y?�G���k��H�0�T�	)��m����4@�XF��iL�;�i_���{�P��5W"~������
6���7��D�1�MY���",#L�"#`D[�f���y��pI�GH���a�\E�1�"�Ӹ��sSp;ٲ'�D�H�B��l�)�����+��l+#��< N��Z��ST@7;2�����@͜5���hk��'���"��~���xxߓX�a VdV㳳��ˍ!�V��O����/�5$�,��c��F�]!��iफ़�E�:�'7y�2s!�Rq/r��Y";^B�Q���U�Z�����Jg:�gP;"���%���rě�I}�仠T
O�#q"������C�ضx�A���&T���VF�=/g�#!�6B����gL�}@!\��л�Gդb_m�9a���.m��4�,�D������|Q�ǷH����'�������C���mi�Y�YF����l�G+���0��`�儑��yLS����A�殺�U��2�(�1ꋇ&��de���λq>ʝ[����'�<ZVX�� uy.B�w�[76�g%��G@�!B��L�1i���i�zV�o��3iȸ��p�#aG�E��^�b����Kk��H�j��X�j�<�&	�D�l�Um�W�#W����ǛI<�w�S�a{w�
�~�'��H7?}����!�C����N����i��Ϸv����D�Rȉ �P�[��2��l��uߍ?CG݌3�%���x�ETL{굑��Ŏ�Y�^�^��L(Y$lǆ7��fVv_���>���pq
�R�K�,�8��V'������Ğ?F��n�Ȣ��H[�0`d��\��fL@|Ld)R%
�0�o04�'��7v��8��t%�H����zN����P#�4��Tn�/�/����?Q����3%��*����=0iݏk�_CQsB����<�dY�00�u��5����*[� �"��Ɩ�嬈jv�v�Of�MTe��-f79�^��J�l���]�B�Ȅz�b�$�?U&jyX��*R�c�m��3�d�!�ZR_{.m��Oz�aȍ!�J˘�N�;��j��߰b�^%�TYQE������i����eJ�oU{%�Y�tb�Rt�_q\���(��* og�u?-�q�L�"�"��']0�ؙD' 2�[�����M5�E�9l��*Hq���c����������
>�#TB���Ȅm}�i2�V���-�a2<#=o�iX�i^PyN�^ ����ꖻ�,���e�&/��*�b4E?V���'z����D2B��D��-**�.C���σ�"�¡������*�p�w �y��En+��%+W��%a�Y��M���-�P���dYn�G�)�ˉgR��D�8�x�n>܏�����75L"=��?i<�m�q�=X���a��̍ia�����S[�>�e*��nT�r-G&#�t���U��I��BQ3�S�Gl�z�rZ�]�϶GQg[��i�T9ݓ����xA�S�0����P�!�.�˻������ѝ�5����VpN�$eB8��6K�����b�U��GP�O[b�G�t)W��7�֬5��	�h���mg
Xɛi�̭��4��ݦu�zh"7|K�c,�79*Z���й[VdZ]f��\Fe;�V�fվܡ�n���]H�kcz�Ή��UӓZ2��3k�(r���/2�#� �k�<Ou�t@}�P�o��e+y�n�d.Z̡�bS;bq7a.ԃ�9�6k��w��]�#�����4V[�=�*��=b�.��ީӸ�8*�#��|�y@gfS�E-_�uu�9�4�v��YM����@Y��%���K�z�t��C�Oe`�5m��!�'V ���JՍWa9���;��nZ��I��f����$��lTqj�w��c���v�|k�R�fH�̏rX���w�VL�_sKjQ��Cm^8u�
DN�_9UK����%AB+P���I�T��X��IYP��X�,+%dm%b��VR��aX%T+ -�#�6�
�Ad��b��m��Q@ӎ*���R�(((DJ�,�QA`���ecj��(��*,
�[iIZ��ՁQTZմm��d�R�+!XbW)UJ�J��HV#題++m*,UD�IG�[N��s���W�3��ɤR�u&W�œ W�Zn_�G��wu.� ��h[���zC���g�w�Z�4������E��K㖄&�7���[�?x����9��Z����;����h���gy6�D��k�." �)ۺ��\.�<��4��"y�6F#H�_x����y����E9��g�LQP��s`K=�s��1�o�1�����{�l[>4D)t���rh��]x�l^&<^��P�"Q�3h����7�;2�q\(�FǞ;��A�#���wn��"Gm����/��<t� [D�d����
�fHᬡ��ۺ��"'YE�O$@�K�����+>����S���T�Ѹ2[�#p�\�٫��Y n����17?W�t-A/�m�YN�P�����@�|l�xɸ1�s7�O�zR�cc!ZӶ��1�D	��U.l3���{�z�Ӕ\� 5}�&㳼��\su�uw�����>�DC$d	{"c�9���g������������E��~!�i
���:!�ue�K�8
�� ��eQ��[�׆���x��#җ���<*�j�~*1t���z��E�6�wUM�����.K��$9�����5������E�;t�!��<�Ȝ>�!�e'�"�:�<eU(���
.��#OD�72�������W����٧�����I���T�I�=af\5*,�� �,�%�o+{3�8�A��v�c��vЍ��Q��F~C�־�HEGZ��ԅֿ�V.�owـ�ﶘb�����4���?QVo�g�U�
/(�E�	5(��[w��1���#��N��n꾽�K�J͙�႐��M�#�p#����+&[��G���1�	hJZr�>�?�Q3WȌ�����D0�	�R�q�"33�b�ϵ������8�Z|�<NX�x�<Dijʪ��ߔP�o��Ծf�B�Hy�xn��vt���
Zp8o��ձ�(��G�] �x��W�o�q�;цp�<�A�=�`B,?L�ݔ6�h��UB�K+��Jy솖h��:ҩ�	*�}Q����u���'
��U�cV!n��<z౥]mu�$�������z���)���c`�˅d\��F�Q�k�F��z�I?p�8���+����I�*/�mA�#t�ӽ����?A�Y�Q��l8��uCwd�ԚO,�a2`8�=�Ȃ�{#�t�������P�Q�9^5�����D�jȳ�nz��^�s#�<g�t�|xж��HӇMk�	�+r����a�y8�qx�S�B��><lD�^ml�ojfャۤ8Z��Q��5xzZ"zŤ�˿n����8�/��Q���u�n!99��]�{��#��͜9ʒ],1!ec�T��i�U�7�R� ��:ElZ�J��2�%�9u�&�|J�v]��²&��v�A�a�c�%Vg%���Ԗ���H؞"��d3��@#m}�8S�$�FN���#��Ɍa`R��(U��V�|BM���V3��'���e��莩�vV�����j��U��<��Ǣ(�۟\��J�QVBe��p�;����7w��z��"J��4й�P�㴴��*�
�����KÆ}F�C�l�)cl���^�<B�:�Tg���Ơ@ӑ���ti�㫷1�`;+Ċ�Twc�r�B&~�B��H�w9���]粡䇘�K#�rDW!�<����{(�W���'A������ڇ��X	�ʅc��3�1ƪ�ە�YGv�lN�ˇ=r6��L�|I�U�������"���|�i����F� R����f�y|�ib�΢�t|0p��a�����b��D9t�e��u��̶�0�¢�$��5�!F���Aʼ�#{�O=���O���~�ma��ç !=e@��\���"���f�&E���G�?B-�}t�)�J��F��2�5ha�({�L����q��j�o0G���e�q�=����ָ���Y�\N]�q6�l�}zl� n/s��wz5\�J}�������r=���Z�i�,��(��#kƔ�Vj�-8C#'�f�p�8�>h+�Q�V���8<��`9�m��F�����_2��!�a���Y�,^����V�GN��`)# RJ�9u���s��fLwf#��oU�$����J��C~ɘ� ><�G��5���ID�N����ܺ�G��AþA<N!�Ń־o����mՠw�����B�����tЈ!�2���Ǎ�OM��US�a������0�69x����E�^�����{>|q��L��>���J�_R��@��f��vn��1_!�m���t�8��������߄�>����}դ9���,��*��Hc��d]D�����_ȍ�(��OD��Hv-*����0�2�! �s�٫BNn<h�7>��جL���/���K~��R�ۛ��G�}�� �ȑ���`��9m��nX�����{��x$��s��&>�����
gq��$wc6fb������j��VS��ۑv�[A)?}U_W�zGKVW�~<Yx��L0|I��!���j{k7ˈK�6�=>�,���,Ѷ���O-��7��YP�\8���ئ��dP?]+;'yk�{Y��k�����_3g���������/��ð�Da�*X��8`~a���Դ�^:s����*�Bmn�x�L7��,����\��:���!�{�-�s���xd��?Y�!,y����b�z9��C�i����ւ7�N���X}�@��Ocy=}�i����r:>;([ ������$�, ߮6='�ѕ����W��(��ư��HӇM}ק��%i�3�5R�;�cY{(ﯺ�٧{�G�z*���#`v&px�a5�|������`�"R~�������G"�H��<f�G�et�2�!K����8������Kp��f�=c�!t�o)�W:��T�+(�!K������C�0t���d�"���q�^�^]���i��T��G���n�9�F�y�]��·�АO�9Vk<�[��Z7�݂���/U2��^��X鞈�]�NB�3��ߡ��{�5Vz:�K��ý̩�%<S���9x��C�����Y`�R��(�Di4���WV����Sѻ���xq&�M�I�%��L�66ԫ]Ѱ�H�U�ڗ�xU���
�~�3�,��،;�x�S��)[�bN����l̛��Q#�[I�:5��צ-s���D�3[�&t�eꖰEBNM��k�9m ���W���!�I���xc7v��͡2�Ⱦ[][��!z8M7/��;��7h�f�&�kBU䚪r��C�yiCFuov���V�j����m��cYuh(�R+��쵔sy���6��]_�.�t�4��H�Zc�5����V�pi��^��_)���E���������/w}��f�+�KT���׌�Ցe�PJ���W����c+:e]q��U��=w3�M��&��g���9�p�3�j�6��|%�K�$m,�b�V�XF����#&��~��`�Ӹ��w*���xp��q8��}�,u��������Z�F�:-�/��op�ãzw7���2T�w@7��+w�3��᮸to:�1���V�_Bm��`;y��� U�GjQ���B;�����N4^+��d9i�N��n�cq���qҦ�q�+hhz	o�fš z��);�Rn���n��47����3x����@�r��f��+�fLP�piA.�����
����,k��z�2�g	N۩a��o1�'�-w*�;/ݐi�Әޛ�G:f��(���h�j��v̬&G��������jЁ��N�����!2	.h�.�<���%Y�fw��[J
�ܤ��4��1Ʉ���b����+C���`��㛬-	t������T^��.��*t�K/�.z �;����A�j����`-����2%B�)Q�;�)w%�D331A[+E`��X9���T��y�vgo�}�w��O^{�8�Ѕcj5�BVVT*#T(ł�H��FV���XV(UTJ�ĭBQIiV�mTmlm\��ŐƴQ]�1Tr�5lL̮"�����V�ii[iYm��1�IPm(�WY����[m�VJ�[KU��ԥ�k��)X������3k-����[h�"�
Q�6�-lZ"+jV�%��J؀)Z�k*(�cJ*Ŷ���5�lch��"K�cCa�U�Lcim��uz�;����v��J�fM���],��� ���h�?���Fr����ӟ�t�[_�G.3ٯݩ�����Fo�a�Y�U�ۑ�G���8�]���]%/�1x�mIެ�Iloh:��KU휼��K=Y��Y�~	�x�eH���C<�wxjz��ב���Am&�X<\9�tW]7K!����_�p��ޓRu����.��]8��*Y[2'�����< �I�9�|Ūm�yer���xV_\hx�q���[�`���,�(� N��Q���@�M�F
����TTb�k+�J
@3�rG?}��wF�N~��(k�U��m~��!sG��.��3%���U2)�EL��q<ƾ��	pX�R�[Xv�XUniT�u]���6\N��)�I�\�m���ٞ�Z�a��.��c5�*�`z5:x��(�|#�,[�;+�^@��4�⫝̸���b�lqOq��o�hV�Պ|�Y����k����P�0�d�G�lC���7��7���tA�`�U���9.߉�A�e^��} �>�^�;Kr�7��A�wELv�DGrt8�Ի�{|�l���ʗV^�I�(G����0�#s�m���;�H�#��O�!�wX�D�����t>y|�;~1��ۻ�c���Ѱ��oopo����>�u���M������ʆ��3��ؠ�(:\UY��k_��j�G��gM�O��V�=b6ٰ#�g��<�&A�ʅ�-C����BV=�Ԉ��/�N�Uu$�y�9�u�M�7�\��wm�qW�~�νw�����������y�W^w5*G/pq���VjcJ�c�6��OL+@zwӻ��9l���-�Ĕ� ����e�ĵAʳC�ǣ{Op�^��85t���׋�Z|�'ݾ8��nd2�uPmd�ُ:xD�6�s)u�Ue탽�Ev����*@3x�|ʫ(�Rr>]=��@NZ2��N�Z.�:�n�U4m�g�w0�����"�;5�9ƄL{��Ѣ�ύ�������@(��}��`p�w�b���\ZqF��ɨ^���mfVOEy��+_`�7hc@�c�����_j'��]���VCG���T�G3Q)c�+z����E���+;��{ȳݧE:�7��'��Z�⯟�hz�#���fu{emH���S淽�����9Z44{���*��nG������|Enc�����;�z���e�{�Ϫ?����TS:Pe{�{�V�}c��Y�(z����9�Wmp}G�p�q���6ek�<'͞�oZ$߯��EM����Y�Vq���]͛����[v��EsXF��*�xEWJ�c>���!��I0a�t�8�S+{��t��:��2�9��T���S)�SQ�*�����ZF��X|W]7K!���|�ǻyD�>s�:3T#nF��0��Y:ϝI� ~��':#AyEU��zY�ӷ�eN��1d�Gv��h��6��$әո�i��6�e�4uUV�Q][�M�l��{j��tRf��<j�NV׌�T���J66f7q�jlU�:Y\rЕד��[VռC4�3l���0��VHJG�ͳ��ǟ�WX��jV^�[��|�غLXk�����\����v��r&�.\����-դ�f�	��W\S8�q�tQ��u�7��{B�\��Y��&�dR�����&9��:
ɼg���qO.
����髱mz>O���uyp�<�>��@�w�Mʈ7�;�M��<s6����,�vR2�� �+���םs��3���P_�{�<��k�����TR����)�I�g|����PA���Rڥ�'�;���S7����Y#;��tC,��;V����nX�Ǹ��?x�`왊��F�v�F��0=Kl_��5� �˻㯣D�����7]Z#.'EO�4R%���k�����i��Y>�fKg��%Uw�l���n��r�;�=�[�eon���u��տB�c��qQTs���4���:����m��}�:zu�}/W>�bf��������fR�֙�6����A�ܙ4��>5i��u���=�2��o<���H�B�1ߢ�b/���]y/'�wӣ:=��V���!zD��W��,1�۝��G�D���'�AՇ:	A�l�Ϸl��z�K�4��4�/K��NOq�z��΢qW�����iH����pR�-�7�m���#ڿ:]�+ћ���d����JG�p��y2E����(CŲ{«(�k+jB��sӨ/pɵ+���R��s�77�0��M��Y��'���׽���} [J;�Tԫ]���$-���n��X���2nowW)��k�r��m�]H2��w��W6������/���`�'��5�MwkA�[*�Pv�8��1C�����wG0<1=����ӎ�݉��.�S��x��B�,��ꓡo���@�L�%ȧcu�U����٥�Ǻf�[��ź �������L^G�-�ڵ�Oi>c{A��I�,e�]���|�����x'���ZS~�* m��z��=�U��T��|���8�1����X�a��nB��w|��2С=6�Q�Y\��mˁ9���eDκM̖b�KhrW;�x�,��kJ�U�&�=�+����ɿp�Y�{����~���jO^��ě.� 
軨��ky�%,���4:���g"�=�n�e'e��oԙx�)_oM�g`��l@�cn�ŏ��ml�L��.�lk�Z�#�4w#@;v� ia1X�-,�{M��k���v-=W*e�{t����*��H��(\W�]>��noJ����M�.�P��e*����J�h]`�F�J���:|��If�n��*�#�j�Yk��M�kӶ:�N����'7�i�(FIW�Yo�nȅ_����Ю֯�����I��U��7�I��GpʄS	���#t�*��D���ؘ�&e	}�Cm�ӊܱ�z=�+S�G+_Yz���j_%�Q�{\~
�r� 
�M�֙�w_m`;��0s���]���J�.��P�B��M��8v\�w;+�����o��`o�_P����].|:^3�	��hq]�v�q�R�k�A�cq�#U}T^��֥�݆_;����W�oa��� �tL����y��Z��rM�:�j��tU��Ú"�؎Q�K��:_u�kxymۖ�5x7C/���Zܸ5f,�v:R39g"�1Pwc�R<�HC�S��1��Ȟ�n�@;�l��Y'9m�S��<箳P78�O���[�x����Sjk�m���� ͑9�)��k�ć�r����.��M<���:��w�����^*(*���#-�E��6��*0V-)TUAc��B�*Z�-�2	嘘����#b*,V��eB�eEb�ԕ�Q�h0AUkEQTUU���TcylQ2��X���F*��Ѷ�E�+"��b��E��U�m\�ب���V,�
j���Q&1FбDU�X�#Պ��E��"��z�3T��h�[X�,UĢ5lW)UFZ���QE����� �����D�	��${=,P��]wU�#����}�`A�u���F�������Cz�NW�w��m_+V�Ｇ����?k���[��>���8�f�ޫ�����w�Q{j��m�7��9��t#�6�wGx�1s�9筎*����^l��J�Q���H���<t�x����E�E�A�$F �v�/SC0���w�GuÈ���ϼ^ i�>�V�x�]O�C�ȴ{|��H�0����+܋���/:�zC�o�����6/,;5�������\�;���x�V�M�-M��
 �(]�`�ݦM��H��/z؝�fs�8�:��p��~���+��6S$f�AʢU�fk�a�{p����"Ո��2�sף�����e���=%mDt��9Y�q�x1[�����]��2z�kW��*��[�v��+f\����s�!L�o42����F�z�c+���.�2nPtc�DYpRv��N���Pd�����@��^��k�[��j��WZ�MB�������쯄��X��0�~�@��+�hZF�۠�]��L'��Vv�}@��K�&ɉ�͏�&���Ήru�f�ڏ�Q�@p��|�.O�#5�=��e��U���9An�u���l�m�]SM�ؙ��"�8�<����^o�+��g�B;���y���q�s>��%�[R�ی���SW������6.�|c
��r�Cj�[���,�}��%G�n�Z��J�u�1j������2��Qo�
�3��xV����+*ppx4���;���u����{+��_"d���$9.�=Z����m�?Q��,Qcr���qkkE,{�夢;Z��hP��5�q��ws1���ii��{z|��:j�{#�AP4s�Yw�cn|]x.�JM,�aҊOWod�pO]���Q@�BE���y��g-r���p�u�;7�(J<�j�hW<��M�Qh��x�8������6�nY�8,m΋̩U�*>�s�l��SS��9��6�D3��p��;6��j�����H��;WJ%K�s׷��1SHMc����1��ٓ�,�������x뉾�����N���vM$��RNc�#�� s�3w����&e�܋^�ZB���~{^Udģݙt�R�;mhwL���4wN�.{
JG��������0��{u�-��7��<�]:ܹ�k^���qV�0T"�h7՝g�v	�6�h|=YO}��ex+u^�0����Or���1��Z��L�o���ʛm�<�pF�?@u[Y�C$�뮷�Uo�SyV�JT�j O_��o3tW�*���L������<�F���6�����d_(ٝ����m=*�I��C�A;ՃԯL�%�]�m.��iU���5ݾҗ!�pʹ�k}���n�qS�p��kՑ"%`��_h'1��܇z�se��j�E�Y��g��y��a�}�V���}��	��p��]�-v�q[�eA˾S<�rs��n�Q�_]v�MZ��4#=��aU��%�??7���������=���}h���j�:�X ���E�nhpB�h������}-�]��a�˰b.RZ��1A�6H�����o"�FV���n�Lֺ`:S�E���ȣ%ASG:�:���+iͺsjbg��͑)N��r�w������T[R��|�:%�E����Yfg�=~�{	���B�^kU�Ӥ�ur�I��8UݏkR�@D[��9涨���1��٦لm�)��ӡ�9:n����������{j(�����8��壅�{�t�3:�n]Fu�X��}�-c�:Y{t�l`o77f��2ݫ�_M[R\��2�v�q#kԛUݝ�]��\���5C[-9�{��WarvͰ/���ƙ�u5��hւK�1�J��˪zz'��.gK��1�k��m{ޘ1S(�>޲��Sg{�}����W5�i3�w����<�9�+(uL�/����EkS���LR��u�ڥ��Q���u��d���
��=�uS�;��6/�O�����"��W�g��P����o
��*�h1�c��4���P����Č���>�^�~�n*�:y�R��0.�����=�&e�<�mLx��o8T��Qݥ2���o02�a:�r�q�����QU��3Qrn�ҙ��*�����W���{��?�׍�y=�'k)�^����޽>	�|��'HݢC�B��y��֙�P�m�*Ar��/��D�s�U��9�*�1�\^az֑�k�F����Sj�Gt(���e�:ꬸV^��j��@*����y�8�����w=�%�|_eRY�U\z6�^L�	���/���C��v�`�����}���T5��Ù]&X��hf�C̪��BD@y�����~)w+rc�g۝-N��x/�}��|��L7����i>��6�2��c[t��67�.x{Ҏ����d���
<L�fi~/g�������U���Ӷ����uI�k]�Q5r��\t,B�{%���*r�����K�О�=����Ѯ���M:��V�嬋v��ڳ��#��W}���{µ��ӕ���>�j�.���f.���Y�k�b�8����wϯ-�]�q!�X	��f-��F�/�b�'��=��kw�QU��һ�s�rKshni�{� 9D��M]����	��2�]���%VV*ˋz�f]�UC�7/�eڷ@Izj�ɔwV�W�}n�9���N����5b�6�Wk���6�[��"�jk�5�1�3huvk�h���,�e]��J�\,��]G� _cM���p��)VT�$쩊Ғ�<���'�k�,�1Pל��G)�͋���B�o���'�iTU�L����c��rVbc�����n�J9������D3�,_\s�{�a:�����M��ڇ�ɐJ��2�JU^%��
��(�wI���)^��a9/���\�U �Z��7t���#e�7G��_����3+�X�y������bD�\J-�vd�ޕ`��G�׼u���J��.ܰ�;u�PS��|qS;Z����uELO��R�qԭ3�:�x���n�0��Ȧ8Z�X��������n9�%ն�����6���ux��$�\�)��딎W;��NɁp�!��p��iK7a�.��5}��g5�h�������	��p"�������es0f��f5�q��[�y:
m*ᇥU�&q�J���SM�hf+��'4 Of�q���ӺM�o-�vl���)�OQ��a��O"f�t���e=�f�p�����{����T�K=j �V۽b�V��Ձn��R�K�*Z�eq1��T�z�#�鉙�̥Kh�%��e�[d遬,X�Ҧ"��t�(�H�+�4jbFՖ��\��T��kY��1W-T�P�3�(�hL[j\�FV��G-'OZ)����"T1���&8�m�O��S+�uU^�x�z���m���ݦN���n��r5���<��ܯ�Aǭ��"�M�3�U����^�ʅ��i{�r��es���&�S
z���֌��lD������b5�g�E��+�S�*Ff;Y.k1�L[��{��{pW��:ډ�aڷ��."\�ܭ��uХ��Ɲ�V���b�i�f)�[K�Ke[�}�/=lS��p�#&Oh�C}�o�!���=��Z�����R�^|7���z�7���G�Rtg��֌q=	�I��~s��7��0�nl.�܏Ƣ6��V+c�pNm��}+Z��q����Et��{r(�u2������^�r��DV>+u����U���}�6�c�F�/j�:X%[��$e����ڷf31݃�ቈ�)2���*���xS�"p�:�k=��^[�2�{|��I�>+,"��ׁ�R���Ԟo'���-w"��#sr�T��#%��U3M�l����W4.���0�<�.z���Solv��n���J�$�{��o�л���햦����Rൿ�����O�����f��j��{jv.�M^�!8�r��{��(I/s��l���/�{��X�L�Z(xIS��X���D}��y[�y�S}t'�yZ��]۬z���/GgJеؘ��CDM���ٔ���X������l��V?G�sSh�U�%1���ʎ"/[w4�i���!�S뇶�zp�sW��B*�	����} ��t�g�]�h�A�]N8���g[ڤ�0��Q��F���Y��ޑtM�o���z�ڥ���3Lq�u���.�5�:m���3��E��͎$�M̩[�*Y;���Ε{f��{;�FI�[+^�3!9؎7=4�7����W����u��{��!��q�j����Y�LE���lU=��HO,�&g�vkk�w����H�1��G�6.�:J1�	�mEpw�����u��7��/׾�ة��}�湁��v��\��TC��3,�w���p˓���9�f��
f
��f�yi����+ӏ�n{!�Q��o�䠅{x���Dә
ǫo!��YV���]����^#5����%�퓷W[���e�ر�VC�tk�lz�@���.qB�{k.W��RU�C󷚧��o���=�1�^�n�͎QP(]��e��4�Xw��>�:��2K��'�r���H�R�W�D�%U�#o(R���*Ի�]tz�'H�/����/s�Y�ػ�߹��x�����t�Zv�ٻ'����q[��^����W��o=��m1�m��[�c�%�����}��{���+G0lQ�쵚��yKUs�㨐�kТz�tj�_a5)�B�f�w���hu7�M��n �e��c�V�����>��D*w
����������6��Cުץ
���g0tߒk�5Ny ��fp��y�F�e����s"/f1ĈE��5���dԻŋ��m����Q[}��oG
Ά����o:�w[�����y�K"�vw�vv�]0�.����Z
��0�KygN�1v�^��Þ�6h2���Y�k<��w����@��[�aJ�y�;���|�>���7���[�F�zg
��٤�k�7�,Hl��EOl����a��ݛ�k�C�l����e�O۽*#&\��dS��X2�=����ˣ��^��q�qm��hBQ��o�L��M9��T�ͪ}i��wu�����O6�6�L�Ŕ-s��X��z�c�ۙV�ɜkRdG1��~��0���Z�&��J>Ϳv�v�I޲+�Q3�^�]~L%��ϒ�gέqڷA.���pv<���WK-��٫�6zy���L��IOɃ��s�l�bE&tl���ǖ���v4D���2���#��CI���!&�?G�.=��������I�}��Ʈo�˰��T�ʪ�9�2�b����{�L�<���s0�z���_��n�{�i�;V��C��rh��!��f-��z��w���xO_7�X�[�S��נ���G����H���.��~r��}���c�Ŏ=ɾ/��K���c���V�L�>��w�w��׍c�ji����Z2����x�0�`����W����ܓ(��#��C1��[k@�]�U�KW�T��.�}�7�������_��O��9	�S�B��O���n�^��WW��6y���HnmV��X����n�S�ݏ��/L����8�
��]%Z�αԨln�-��C�.�����zx;d�vg��bN�N���v"���#E,�ݻ���亡�Aӊ}�X�"#q��G<Z��LH�w�*�壘*�}-}3ɣ{�Ra3[�&�&�j���.��{��_y^��w"�Z�n�Hi�S��T<�8�8G�}svz��W���"
�ż��I�A{#	)�"�ГոҬ���9&xD�c{�>����g�Vz��FN\]z��'�w�y=­rS˫�*!��
\�q��t��y���?-�3_{S�צ�"0}�aT�L�o1z��f��oLզ�(n)�<�YTk̎z�m�������
Ñ�
���<\�D{{UT�e��UUUUG�*�@Iz���	=^(�jBM�����L�8��ݕ����aY[�o`��1Ɇ�5����I�$�d$$��H0�lΆ7�溏�fB��X���B����C���rպ��1i-����/P@Iप�Y�5V��;���=��%���貔�)1bs��_�#3�i�vZ<�2g�a�R�����'��
�܇A�9���@I��_��ڿO\���RLâH���*L�@��<ETZK�#�����c�����'�LV~�ni�����9LN�q�IVu����C�#��;�b����3=��t����
Fr�/ֹ�db�ԏj�W��}�a�j�I(Ǜ������k��sёL����R}�VBJhߊ�\��U�v4�z��J`��G�^:�	$�V5UHj�-.���fu\��'�L�#�!�b~�]�@I�L�d�UU%�YÁ1���i7��1�^�+�v�jLM綣��#��>X��lb�9=�g���g�2�l�ؕ,�&=�i*k^O9�;����7��Ɂg�M�\,�k��X̏ob��\�tv�r��&$�����_l��������ngroJ��ӟ�ҔQ�=m���M�Ox���:�E�-in��$��=@I�>���ME1}TN괪�8�0��KpI��Mŉ���2n�dd9�J*��Mb���J>Mt��"@��Rb���b�8�̤�a穯
�*2��Ԗ<J�^D�^I�R��
K�Z��3����U����"Mr���x6$s���`��ؕ�z~�$�q����R}��Z�����<}�����;��2mad����]\���v�}�Q�TsH��Ŷ4�>ς�@I��8c��\Uz�k,���ލ"�Ѐ��ybe�V������p6㗳ZoF��K�#�឴f�h�8*^)���J.K�]���|}A��Sm�H֣���Um���^3MMg;��7d����G:2�;#>~x���ז*���YM�wo�UQ�f}Y[��Q�=��Gn��T�'�J�y��1q�����^s���5t�8IvI��NI�`m2���&F8�ȲM%C��;�|YH�R�Q�O���6�l�3��]��BAlo