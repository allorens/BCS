BZh91AY&SYw�:���_�@qg���c� ����bD�           ����Y5U���i[5JT��T�2R5F���S3V�fT
[hKMm������fōR� -�A*hV�Ui�֛f�U��2��l�Z�i���Z�5�5��T6͆�M��5R�lm3i�E�V���1��ih���Se����d�m��� �   f�V�ڥ�n ��j�2f����MJ��. .�Ք�fC-�ѥ�5�֭��V��kf���3-U��Z�me[T��Z�khj�ڴ��i���l)i���k�)H C�����PAj�UV�=:P=�v
�Kqlڝ*�H j�wZ��[i����t*�u��"D�ܥ�uiA�2�Z�͕�0�Z���3�R {� ���l)A��{ƽ�������(S���
r-��=���+�q�� U�;� �W�����u���{�( �zf��%���&�mh5��[*hy������A�V�%f�à�j�d��v�[((����������������	S�Y�z
���ҽǝ�$��e��G�D�� �����Z��6��MmR%[i���H�{�.cEh���{�R��wI��*
����^�m/=4��;��e �l�-��J��P
��v�ր�U�gtt�I�]V�*�V�`��֩��ɨ<D�(P	>�� �ht�KW=�R�kz����r5;��Қn�pP.��wW t(�q�4�AB{�����Pc�Y���jm���P٣F� ��z }	�7tV�So{N�Tu�s���жPZs��MV��֎V��s�;�����֚ݶ�Nw:nS:@.�T�P�*��M���j�� ��I	�ύ ��Ӏ��]�.�hӮ�s@ su����  �si��w� ��m��4u���[-m�����fִ7�� ��A�}wf�]��g�6� �`;gC�>��� 9���@:��ˀ��� �˚t �9.�B�#[U��U�Z� ��� (�� ���� �� ����	�sN�GE��� o+  'W\ i���{�G����af�-��L���MR�f־})  �@�]ƊT����I�c�v��к;�P�04+�j��;�\�6�k π �JAH ��2���4�  ��   �=��)QR4`	��10d`�j�������&@h�   ���SR�P��4��  0z�!T Ѡ C@  $P?T�SG������4�4�M�����E'�����#���b^7���.��;�՞y;�|��w����� *��TV ���@~�䊀��<}�?w���>����3�S�����I$���P U�H��B*~0EE���_���غ���b�X:���MdbkX:��.�u��`�X���q��b�X����b�Y��5��]b���u�kbF�SX��5��b�X��`�X:�5��X:��.�u��q��q��X��5�k ��X��5��Mb���!�X�0u��c��]b�5�kX��1`����CX��M��`�5�kX��b���k ��`�5��X�u���!�CX��`��5�kX��k�!�]b�5�k15�kX��u��SX��Mc�X�5�k �!�X�b���]`�5�kX���`��5�k ��]f�#�1��X:�5�k �	�X&�db��!�X����X�X��5�kX�b�5��]f15��CX:�5�kX�����`��.�u�kc����b�X:��.�5���5��]`�X���&1�.0`�X����]`� �&��Mb�X�`���bk��.�u��`����&�q��`�������`�5��]`��.3X�1u��]b�X�tb�X���.�M`��.0�!�X����b�X��:�1�k �.�`��.�u��c:�5��]b�X:��.:��X�u��b�X:��:��b�X:��.�u��]bk#X���.�u�kX:�5����.�u�kX�u�kX�����X:�5�k �!�9���.�u��]`�X��5��5�cX:�5��]bk �.��:�1�kX�b��.��]b:�5�k��CX�&�u�k�!�CX�`�b��5�k�!�]`��5���5�k��CX��5���	�b�5�k �!�Y�SX�0b�5�k��5�c�	�GX����X:�5�kX���5��\f�q��T5��`(kCX� � ��T5���&�@5���@b�kX��@� .�SX �
��5�!�A` �CX � �
��*��D5���b��Eu���@M`�kX ����&�T5�.�@5���@5���Qu�!�1���� &�5���b�kX��P�8�u��05���@5�!�u���U�
�D5��`��X�� �"�@5���@5��E5�1��` k X*� X �@�(��@5��1��� �*�P5�!�P` kX��@�(���(� ��5���P`�kX"��T� ��@5���� ` kX��X��]`��$c�]b� �.�`�X�u�k�C�u�kX����]`�X���X�u�k �.�`���`k�b� ��b����]`�X:��.�u��#X���.�b�X�u��H�X��u�kX����`��!����5��X����Mb� ��0u�kX��u�kX&�f�#X:���]`���u�k#X�u��CX�bk �k1u��`� ��X��u��#X��5��]b�X:���]q��.3_��L�}��r���go�/�$��ecr�Kb�l���zj]�)�n�&m��/e���z�3o%]e�$;�mG�2�-ʱ�t�e�2�n,a�ʷ7T�1,�7�[�i����K��n��`A�[�ժ�`ms��(�U��ۺ{�(6�I� �NU�(�.�˗�r�̹,� ����4�AA�o*X�h�$��n���^$4�a���j��o%�{WU��6��c�Z3�ݺ�J���b�0��WH����b�C&��oEr�����UV�P6ʛ���~�!���o.4�mKڙGM��2H�4[۪��w����+RmF��zD�IR���jZjNRT�Y�Ei�.ə�-yqW�&����0�-^�T�p^M��2�u�<
Yt�'א#��]`ɛ���f���e0�nk6/4*)�Ne̢��/rM��^43�.bJ�l�3֦�c�,��Y`����Y&˙l��e�����3V7�{&�Į̃�P܊@�S8�!�Q��ߜ��	�V��r���iך�%ɥ���P�)c��˘�cv�kew5\�$qd��{����le�S���|
��Nm���5dk	�f�+�k\��՛�����[q&�Lm1m[�cZ4�h���(}5e�J�Q�x�E�B�����b�l1藁ے؆�FZ �)h���7���{n�kYnl��R��NnV�v�=@� BD*�
��Zʧ�1JV����[7SȞޘ�U�4ˣ.�l��ˬ�-��f9h��Z�t�}D��؍�{v�,�:���M��m����e�jaGN�Z:Ò�9��I�y�H�e�%�2��3-��.��m�j��nb�B�fQ&�w���6��K���5+�V�`�.V��{��"RCr�GK*oEA��ǆ�J���{A�D���vMm�f6�XkJ�C�k)YF�V��d<� �mU'l`Gwv��G�)Iݶ�c@��+Rb��iO��u�u{ʎ�tS��v�V�� ��9��l>V�*�֭ٴݬ�=�6�H�H�}|y�U���hM���v��
*d�.�lhѰ��1kǘ�f�*-�ٳ*��c0����pZ	(Q�~y�I �x,������3 ׶j)��u,:�D^"��mJ���j�f����	�uy���iec�L��G�a*h�b��-��o9-m;b�sBͬ�X���Q�ٲަ�X��3Z�ffJ�Wuc2�X��7�)��Y4Cu(�)��M�coD��f��+G	id�q�w��5��X5�d��Y����KC��d���i�V2�x��1�(Zj��0�w��"�eT{�P��-�]K ���l�1�Qi@�h��E�"�Rxwe�Y�壕�ʽQ�ך�1r]9%��E,	�n����Yinhh2�h���E���5�_����w,9�2�R-�F�C-����W�c�+)�,=�(�3j�ǁ�g0��5�^n�����Sn��{��ʌ�uoh��Oj��R�m�gn1�e'LY����5�u���X�4j�A����wZ,�Xb�V쇘`�g�پ�L��;r,H׭��C(�zq�dG2�nlx1=�u�0�%�կ�w�S̹uZ.��eV=�2�ѡo6����a��J�X��p�Աt0*��:/r٪.���T�A�p��.�C�Yϗu��5;M�#<��PݯbU^a�M�hnFk1Y�Q�QH5�l��*mn�N���Z�CA��QD&(+[��ڹd�0�˼�'�奐e`��ɷ�j�-�*`�*]�%!��۸sZh�r@�d)BD�Y�N3�]��kf���a
�홙C���M3�qb����p�/eJ^G�6���Y�:�l�h�!5��h1x���ה���rۯ���XV^'��Zv��)�VЪ�܌� v�,.n%��r�X�o��J�&3��/or�Efk&,.v%�j��r���*�LztK��2KM�J��Nc�P�ꛛ�I[�J��7RY�]l�/HףSc*���4��7[���kal�7��y���)�Y"��5�U��n�#�jp�rn����Q��K��i	��ʩQ��k*����B3^-M*4N7�ݻ���y%��}7N ٛR�N�/\�Аy�u�m�.�g]u0�5��Ⱥ�6�P��/LƞǙHV��%:��S�Z�f�&+�K�p��\�fq���R�ْY̘E��6���^�D��x5ɕ�e��	m1������%]��on\�&�a(�n�YnPf���gU����vi�0�pdk7�L&�wd��0R��� ��%H��WIi�պ���c����ո��Sr��:̓7pV1.��mj��EUkӋ��qQѵ�����H��LJ���)�Fh�n��%�ֲ�Q�UI'�q#+�<�m�Jj�Z�ʎe�)Gʙ����ybճ�V�'(��<��m���Yr!ЙZM=����vƫY�e�Lo[��ރh]�W.�0��V��x7M�zh�N���a�����*�kFe����Y	Q��[����׫.��jE�h�c"��1Uܻ�t6��Qn�d#F����n�B�A�o"�+e:9[#�N��[4]�YsoA�O��b71ݱV�7�� �bc���0C��,���$jT��D�����=�1����fY��MZwui5�ޱw��3DR���f�i�;��t�#~:�֝lͱ�F�vH�EQ�{2YiE��uHT��\vn�±���ҷ�f	b�ddQ�+R�-)�BhY�m�I�v�f�ql������%�+ަ�u�d0r��3MK��&Sj��k�r�Ѯ�2q���s2�XU�7���	e�2U(mb����Su�YԜoe��F<�h���XBW�8B��$�d�o^*�(���P�.�[R�( ��H$15����N�UU.�����U��I�,=Ė���u�US8��qR�E���6��F�q�m�F�'r8����Zݦ�X�%�gڵ��i'��fd�J#�zH�n�T�J{�[Q`��T��QI�wM���T���	�J
r%F:��u��MkJ�i�_�X�]�*V�hK�s4�"�����쫣��$I㺪כD��+�b�؉�ui�^��ԯj^F謗� ei����l�9Q�����I��p1�ͭ�ȣ�T+"͙�I���i+�F�V7�m-;�l��Ze���2CˮOR ��Ck.���1s2�#`�k$XǏK�aK�S^]\[V.����1a���bv��ł��d{bв3H�f@r���jP� �jf��&͐�f��a+wU(�j��Ǜ�U;���B�}�'E\�+e��w��j��0���ꨂo[xCَ<��5��Z�f�t*��ZsM��4��Lĉ�e�ˎ��PpX'f�,J�gsԲV1y��f^i䅹��b
��V�&�l5�㔷sUh�6$�F%��<����h�X�;b�t�9)�{W�yl�)e�)ث�<�K$i�����7Ic�X���I���3��ӻ�ek"W��E�{��n�$��m�u�UP��1�([BnItB���i�KS'
�T٢�����Y�,#�������n�BA�Zx�Nc`�G�:x�����L�X�$�>�pk�,$؏2
�k��t�FE�]HMa7W���-���)��tG3Hǹ�3Gstf�i����&�Nq�m=a������V7.<�bZ����iۺ"u+$M���	�i��������"VRc��͠�Mv�V�����m"�н{x�O̃Duhf%:�'kth�W�c�gc��v�09R�����1�����r���",��呖�n�]^*Pn��]Ju+n����/�楋a�{�^�Z2�:�)p���A#�&l���Ի�3S�B(�2e�b��c_�8�M��T����|�(2�A��QT��8i퐣+nb{&�����!�ZܺIn�s��	�PŹOe����mY�c6�d�K�N^J{�KU${T�͈T��<�m7���������V�w\�0��j��%��0�W��{gK��f�d<\i���wR�L�� 2�?<X-��M����z)�/ύ�̍V���D�j�Э��)
�:�5��c�b9~���ay���N�j���p�NE�J^�����i���3V��"�]c3*�	�W�9h�l��yI+�Ɯǖ)H�ؽ�h03F5k*e�oI�[Sb�N9g����P�2��N^��m�{W�NmL8�G&�Z�H�
�t�c���ݺW&'�UMVr0i�C���#e�ud9�*VG�E\�sb�u�e�TS�(/�m���h�1L���[�@ۀ������;Z��L�yK!29t馭��d;q7b�{0%�����3(�;�^Jk(;�=J�m�$�8_�35M-�6��u�56;��ǒ�&��ֲ�V!�W5f�m�Z8��w�<��3`���+/Y���xͱt�)
vq^<�j��\�[������ƐSژ��2��z��ӥذm�Z3�6�tG�&NML�r�Y[��N�ʹ�e���$P��\Y���l�m렎�Sv��Y�x!��Qtq�2�-=:7dG�\�6)�[
��nظ̌�e��ӧ(��W27�^UV�u���e��d�eTx�"PMݬ%�*a��H"�:��7
�Dm��/�C�ޭf���nڽj��X���5R��q]�v^�
�b$%�U�u�Lh�z+���6�r�$؛���55�D��M�T/ː��mXͰ�{F�|�͵���4qZ��}���5Xsb�e٦����U�WA��]��ų
�k(,ڰ��]�^���{�j�m::$��2�+K�lS�$;�t;�Ajtj�`!���[�j��������iB%���(S�̫���je!�̧xm�L���B��mء���#�m��M��V�A+tZ��w#�懘��֭�Z�ȪVɧ�36�դ�9�c��i�h�$��rJ�n�U�L��ފ�q��fSW�P�R3o=H� 2�&՜��h�78�e%��UQ-.�GN��,F�܆h�v�
jY�XGrjh^���8��J/k)l�W�����6���Q̹g�t�������`��c)nm37�:���U��E,�ʕ&��km�9-��ˆ�E��u5��uTH*�U�-	k�)�܂�QL%&�z9�p7�{���7���9��R�ö`�ia%����0�㼖F�ɺoi/n�[R�e��[͡ZI���Ë����{R�3s6J�äb�Pj��w0Vs$��ķAxKʔ��4�dH��n���#S.��j�/&F��Y��zQ�mmY��ͫcvφdJ�2Z�7�W�y+5��F%�}s��W���K0��:�OFәSn�l� ̋F�Gd_�E�􌍼����w%�B�3"'$���[ԉ�q�(�v��p���*�z�Fc�������ߨ���W�V]�ҷt��PG)R���+�#2 ViCT��MȖ��I�2<�b�~؅e��ej4�S,��E�/e"cɕ���C�{�N1PjW(��,cmeE����A�s#��[1Ӭ��2̚�f���cZ�����ۺ�Ĭ����������%�	o�%��H�:�w�m���;{�(3���خ$��y�!4���u72���b�[qI+5m1��$.�R�MFq�ý�w�,��jk0���7xq�sA�6N<9�1�3�F;o,e83t[t�z$���ؓ�v�����/.n%�C[%n�5��N^+�or��N�����[֭c0����k�+V+�JW�D��m3B�BW��%�ލ��i�Fc%
4�IS^J��tpJYg�t,�fI�ִ�"j��M�ì,{�Q�C�w%UV�K�`�ųFCP�.�#eQ7�h�H�u2��T�[��C&����`���CO
���P�A=�w��"�⋡��h�c-���ԫ|גFu�/+.%����-�J��r�-����5օj!ѧ��%���t-8n�$HT�J�J;�-�%MM2L�%.��������(�#5q�d�"�*"����!ӺG)'\r�Tf�	�]qP�͂��f��$^��Wzݙ���LO�6�Wnf�;��xӳ���]]Ygr��O�ST��]���;K)*x�͂�1+�����0�㝩�S���X�EZ�����]�b�\�"�[�`�ZIź,�5�ɄS.ٷ�.�]V�.�[���,�[XڤڻJ�Ԗ, �X��\���Ŋ�r�`�M5iڨ�깆�����F��BJJĄd�U�n%�4��5I�IkV�E�*ő&�3��4����79�VmpܫQ�����h2�6�i=Z�Pa�v�G,�ѕ��y���k�%���F*��F�g.L2�U3�gs&Աr�f�y_y�y���s)i�DvZz�]c/�fn-�Q��54J�wY��ԩ8l�,�=}�GHs2v&�2ْ+�T�Q�TƯ�{,�h���)�^�x�+NM�w_�yP���@�)�Qe��v���Øgs���AZK9MR⋒�C�e彪�pi҉%oKhM�֧Ԉ��ur�J})�(nO��{b۫Q
����J�ڳ�����̚����.A�><���ܮ-�[�Ί
��i�\!{�Ɇ�D>VGgu��cg&�rY@�DSJ�G�K��1隋�'WI�1�]�,�Y�-������,i�HQ�6�� ���w� v�+N��`q7��qʊ�j��U���>"�e���RQ��H�CF�Vy��:k��b^�?����|��,��;HE���˛�f��l�M�$a	�i��Neԥ�[X����� �]���*"�[-ԫ	���LO�����i%R�.ja(�d�f7����R�q<-�;]�L72�y�w�;S�X�,���*�Đ�[*��\,��*��I�Β�i�ںP���Q\�n6��]	�J��)�1׹��-�Y]�n�t�����}��OF��T�I]��v�̍#�����H��o-N+B��]�{:,�	��urZ©9�V����INݪ(:�nH��������������������0l#3��?�����$�I$�I$�I$�U6)�JAF�y9�}�� ]�n�7Wj{Z��R�m�!I��(79i�ˆ���\W/w1l�G��|��O��ҝG%��	L꺉YZgCu0v�s�;V^����lQb�Ҳ˲͡o���yh6¨i�PX��Yq��T��z��T62Q�(h���w���wQ9�,P#5� ��s9Hr2jU"���w������J�묬�*�/�,����U]���$�6�Kކ�F��S�7��=Ɋ��m&�\�*���Y��Y�����WFwtF71�CP$���.7�b��zIO�Wۅ���݄���{s�Kw���:�>y�V�n�^��D�q�%Ó���V��2���Xcf�mM�D!��H.��3����>�W�6@��[(�^�n��z1lAv>���Fdj�t�����*����u�W<��^�-�̄�la��}ִ�uV�(j��^D�>��&m�y:��z�[�#�gp��zs�j�2���6�ʾ�YR�\;:C>T�r�[��5{�do��jH�jA,��\��fX����$wb̕J��I��T8gf^W�Vd��SA�2���u݇JI����^c��Z�qJU����{R9\�/q�vҫi�/�[��Ʌ���[�tǴS�nk|Dw�����>�z�.v����9��rV7�6�[/P�C��^�ww�9��n�BOF4�v�t9Q�*h�*��Q͠�62e�7�m��g�,�jb�2D�W�AO�q���UUc\�9�+.ؕe�M8a1����\�m���E�����R�����ĭ��ž��6�z��Ո]�}�[}de�p�O�ݒ�r̝U�:S}K�5!T�rٽ*=��]�3��FxM=�P��8�V":�M�n�P�)e��J_o|g�������#�g�;e�,]�lD�C��̬4j��kU�m<�km��C��/w��m�^c�t���i�k�.]Uw+�YJ;�Q3}��Z�I�>������^��t�:̭��B���w�u�{M�-୾����F�wr���g)��^��F�u}�$[9��6�/q��J�	�.�n����c��t����&smi�u�9h��Hs��3Y�,&&
$�a6�C����u޴��Od���I��[{̙���jX1-9Q�6�U`U�S�0`S��ηk�ަnf;�O�-*�p��q�%>+4kt�+��*��{%��1�q��j�V���k�w,�VKMh8n�C�γyl�u<��M��$1�ߗkј���Dw�Ӟ��#.Wu^w.���R}8�OCVU2��+��[��Tܚ�N�־�%�w�;���UB$�[�T�<y��#�������ţ�c҆R�eӫ�A]�T�F_J�Y5�So&���W�[X������]Jۧ����T8�N%Y�D�c�'8�=:TUJ��f�&A�rm�!g�&��Z��dB���kY��r�ه{����P�uXD��ɳK�}�伥��&���{bro��\���}�[z�+�R%AX����ʡiܓ�(-��F�U�r[w�t��[��F���.u�D��bfSgb�Z{��$�3���5������]�6k�);��$sx��0p4�8jI�/�s(�n�k�w�zLaI��ಂ;X�^����ł��Q��<�w.��৹%ű��U�u���Ӡ��s�=�oNUE�S�w%�(�؎���n�ָ��0*Sm���6�qE�D�ۏsqjr� ��=p�UR�)������4��h�gs�G�in���EsЏT�T�ER��٤����9���-�aT5Fc��d�ʒ)�4n�V˪Pː�Kw**�J�	zy)�o�j[�a��Mg��p���}%'.���3��Y�tf>9z��_Tc����8��r�vWCבu�S���;��i8�fU�3�ҡ4��]�٪|�ջ�3#��ƅ�4[ښr��n�cO,���5y�Oe�l���]=��<�TE"o$����+T����!=!���b���܄��eJ�}��37��Љsn�$�v�-p�ȓ���c�9�Mpށ-{,A[})5)�p{l�U>��;���U�ٽ1�w2��Lc���֋#LĆ62�z[|Nzý\8X�^�G`��@��Źr�u��<��F��*��tՀ�\"NWa���w3�׊p���3\URV�k�N�۔��[y�rԴ�R���xcRT�Y�I���u��L��WvZ����{�����r�;���)39v��C�)|JDvm��K�w�	����RQ����hqΒ>Q��r�PM$S��i�¶�Q�Ug�e��=G;vT��\��I��|��I֞<�Ζm��i�f���M�3���Ή��t�`� ۗ�Z���]U}����Om�#�}z8:���$Ỏ��su�Y���>��9e�S��t����7s�܆H��uS�q��v]��q�۞+Ǣu:ťT7+ݭz�L^��ӦynN�v������B����b�<qƐk�R�]��J;P@y&Sz�֋ˢ���`}�jJ7|�(�����aޔُ9W�Ul��_h��i��#wxiT2;�5��-]hH1�n�{��S� ��黉ѼO�>��s���4�c{w���C|��Լ]�_:%j��9ӵWwe�4!R��u
�M�t�o\�3�
GIc\��;���[SK�P]��3�+j�N٘���*�^=�C-�Zu�o8mQ8Fg��y*=S��+�	��35����:b�����������m��{Fv��B͆�e�uwe��%�&b�V�����v[f4�K��"Եm��y��Gl^G�.������/�Zдj�9Ph��V6'C(�yD�4�eӭR���8���R��G��8�K�Yv�r��Y5!�Az��~��VچX5/�[;1�%ײQ�z�IL�ɥ$��-���
��te�olуΚ{I���7��.6r��;�ٶ�<S2��U�wr��th�����`��
y�ֹ�;J�wS�u�h��y�2Ѫk��!u�VHGY�F���]�ڣ�u޹�Q��R�DM�Y�b��z[\�a�30�֬9BpAh���ݜ��nݳ�կW�u���}ʇ����t�z���h�1�L9H�YskSZ�.U��d�F�B$�j��oB�{ܣ2��9F�K��S*y�h��8;f
���m��۫����:*��v�iSRy3�i�7U�U�N��(����nK�9�jX��wzV�NỆ�޼��y.����.�+�O;Ei��91�0��Q�v���R}�M�q�ʯ��E��ҝr��{ҭ)r�'unn��3�O��rs�5t`�.��7pp�iD�4��"��{�U�v��L�}���L9}k%ȩK��G��*1�z��M�s�!�a�/�'�)�锶�H]��ϳ�e���敔�or�o���$	�/{��њ3�`!�6��yH�l>�x�j�DoS�����I+���(����Ð� 좢�:|�7 ����@��}���)����n����V�5%h;�J=�n�ܶdu%�]�u�1����;���YT��,��dJ�����u����Y[�n����9g��3�B�]�:��IW5������k�>�Q{�/s�m5�6��q�t�]=U{����ӘNU�i"�Y�,n�J��۝F��ncZ���Үgwc��[�]SD)̢�0�˭q`��Q�1hζ����M&��[ĸ�Y� #�g��$�۸��s*�yn�ihj�R�1�����*N�=u>(1����9��j:�Y��&�-���4187�b��}F��oD��Uxq64)0oA���r�lb�~��K4]>�Ӄ�ӎۦ��n@�V�:.��yj��X*'n�D���c��� �
7�fsfWf�w���WC(gD�RM
������s�1$GYV^���M��{S}�2��f��g�"��X�6��үT�Ū��r�1*ll��W*�ޑrZP�Zn�}��Ou92H���Duf>׵iAh[�4^�r[:%܋���؛�X�ݍHw�N4Z{l�Ի�-w����9b��mg6dǸCo�#4ٕ9]&�� ����o�W�4)�z�K{t�r�ӡN���-���v�H`�׽�^t}��Q�.I�VtUّ�9�f�U�%�8\��&��{B����v��o���2��۹˒Wa04�7h��nKyԟ4t���C�i��t�l�����s������o���eѳ�b�.��Mݻn�ydu�}���r���Mcb]�Uݝk���"�;�u��b,O��vƙ�7�Y[����j���x���*-Y��9���.�Wf�Yz�{��jj_!]���ޙ"|:�l�5}o��3Be'��YKUX�kq�ki�Ή\����c�y���b��*��h��s��o�RVv�Rp������ɰ�s������W�K���XM�i4������X�ٝ��5ph_R��zd��٣mÁK�VI��}@�]fX}֞��9��uִ8��x"۳��f9�KF��}���퀩��Z����� ׽Bq�!L�r��\��,�Oj���� ��&p[y�GL�U�˰L��;cK�e�wg(ar�J�TF۾D�r�a檪�>d�u��3oVHQ�.�٣rpyv'qܪ��?�S��5��<z���Ǻ�K��iӀ���́޴����vv�&;���Y�;o&�NWw��,��J��@�Ur�f�;u��Cl�	�p7��7Y�^��l�f�u�+����|�]���
�؂	jlm=�$s��Mvq]Y:�4�{/�Յ�)��ⶖ��{]A!�T�ʆI�{K�ĩmmv�j��\�
��t�m3Ǣz�N�"�w^�hh���x�sFv�7&Ն�T�(|Dє������oF��ֻ�s�]rɼ/3�'(��8&�5bЏ.%H���ٗU��R�2��$I��+`�5��dr���屙�s0��"�\���.�ʫY&�*���Rj�{�r;��T:Ҍnl⒃IJ�ŸY�)i˘by��)"�
���6�އZY���h8ԇl��6��_ZMl����{����
�[��:�)�U+E@�<���C�9ѩsk�����N��oӪHDՓ�m,:o)��<��w^_T+�]Z�}��+q�VěAe
��5����1��˶ٙo��O]�=ӭUh2�a�$n�q,�ʨ��Z1�ʶ����]�A��������˴N�[�1�<�L]��m��o��\:(_:��,���x�۰O`w'nWK�B^A�&�f��s홮�[2��]"v���,%�n��h�6�4�)Ъv+����:Չ�!|���T�p![���Ew6�x&�V�Mj��f�[n�7��k]��frӗn��Dz����{9����_.᣻3�ecA��H��;u�����~�K*�D�e9��r;e:n^EM7v�5�A;�=�\�J}NB�+�ʐL���^.�)��P�Nc���8W;�Y���xL"�qc�^�Ӥ��y�Dw�K��ߴuV�9�c���k{��G4�,�Պ:cSZP��o�����C�nJ�U�$S��8^���iÊ��QX����d,#9fiN�ڽUq��;t��έ�H��M�:D*TtF�JLT�����9��s�Ng[�H�&�\[y����1q��IUx"ξ�����c
�+�t�'rN�t��������ɇB���[�XŮ�ڝГ:�v���-���Q�ciՙ�/�0���Z�^B��Q_UN��x��W}L�\�5b˻��[b�0.��3��t�nXY�n��t�n�s/w�jǑ��r�q�pNWF�16�R��@�ܒV9��v�dBDy[�̒�9ɵ��we�o�P��W:��b���S^�l�ձ�Pc��|*n�:	�G:��r�I$�I$�I$�I$�I$�I$�I$�I$�vji��]$rG$�I$�I$�I$�I$�I$��Q6-m�}�M���mBd(`��ߧ�v���O��J-�4Si�A(�ɥi*��$�Y�����p�N�i%��E"���
(��( )�H�#�m��O��#q�+�wa��%��EE�`�0�"�Ŗ�qd� I�RF�%ڨ�T~2@� ��"��3��P�D8_T�E�PdB̠ٓ�(���΢��&x0�V*7E�BP$�N���A�Ijg`���0�ل����f�%'Ey�UN2�A�v���#j��#nȢ(�	�17KhXM$��*Dߐ^�I
6mJ��a¡�tO�ECULP$B�4��Q�wH�ID�RFS&!%�ID�8�l�DmH�q7�"�ㄻvT��H����$� �^�6�u�I"㠈%T񒋨��7DF֩�!�6�!B[F$I
a��zy��L�JR%����aU�HЅ �j9E�&ҁ"�� 4)�!��Kb�e����$��n4�~A�����h@��D1>�p�D�=!�"�F���w���\e���%)�N��t*�L�%��Ji*L�#��Tt	*5.UUH�15�3��,���q��Lb�D-����6�tXC�].�,x1�"����0A$&��4�5T`��-8�n��Ri��YM�P��Q�2�f@����Lq����x�w�����_�����AAP���K�=�����>��? � #�����������������J�U�������������;[�n�������ku6i!�y�R�_cP���X0eK��Oj6��P>Q;��T�}�޺��1q��\;]�G
r�j�̣}�L<�uw
���|-ųpS��g9���۸�)�mn�����2�,�$-y�e�+Y�P�rH�C4�ƮT�B�9�ܺ��w�u����`�$��=�V���6���S�S.��rc-�Nju�bB��.:��Ƕ��z�1I؏GmUv���+��WK�����T�Ku��Jb��ѥw��ԃM99��9>Fދ�<��GlmsZ�B-6�<�Fa웯~sks�K�R��Cat潮�Ql��D��U�����	b^R�A�����q�݋�BO�
�a{�.�!ci��-��+Vkm^wuVHp@�D�O��n��W�8�'�IX�����mǐr��+w(�dtb�T�+��s������m�x��F$v���/jltt+�L�jڒ��WJF`Q�1�FUԏ�ͮ-T�F8b�-n�Z���_<ףK�G2�v�V�Ȑ����`��q�P�YkQmS�㡆����Gn`�������k�/Tl��-��z�q�ί5�����ֽ��q�kZֽ��q�k�Z�^�5�kZֵ�kZֵ�Mk]kZּ5�k^Zֵָ�k^��5�kZ־4kZֵ�k�Xֵ�k^�ֵֺ�k�Zּ5�k^�ֺז��u�kZצ�kZֵ�mk�k\qƵ�Zֵ�kZѭkZֵ�hֵ�kZּ5�����kZ�ֵ�ykZ�Zֵ�zkZּ5�k^Zֵָ�k^��ե�&�9�μ�:�9�%|>�ͱ�&�F���k��kS[���a�ɘ�k8d̺�!�|1c�_J�&�X��3�b^��4/������[5�p\l�[�Ӫ���V�7�4��r�8�b�r��dk%���ν'm��eZ������|,W|����2Q�r�����	\���H���6$��y�3�k6�*(xn�+x��Nx�C�y\i�X1�[l�x/4���p���Wϲ�.�#��ΕU�;��T� T(�Q�]�l���(�,�����9��}�>۝[���x��6꺺�NV	�3K-]�w������DU�z�[�I`���vH��lH��l˨������f�)�h]�{g
�-\e���כ���(��%ҳ�M�j�g^5Z��8�c�VJ�nV4�t���Dd�9ףxͽ����Le�K3Gff��b��]@_�s�����O��o��e&{&��3��l�-�N٩8�y�h�	������s=��'
� b��3�w[��`�a����U-6�WկJ���$���F�s��MgL��*'1>�����c�s]-aŇ�Z�-�rI��:t��y+
YCx�ݦ��#e�� ��\�2�+��%yT�WiK��'�����O�����ֵ�k^Zֵ�kZז��xkZ�Zֵ�{kXֵ�kZ�ѯMk]kZ�ֵָ�k�Zּ5�k^ֵ�-kZ�Zֵ�Mֵ�kZ֍kZֵ�|kֵ�k^��ֵ�ykZ׆��5�kZ׶�k�]uƼ5�k^ֵ�-kZ�Zֵ�MkZ�Zֵ�OycZֵ�k_Ƶ�kZ׶�Ƶ�kZ�ֵֵ�k^Zֵ����%��3�{�wyѼ8��\=��38Ƶ�6��[�-����ø5] ba�u�	P�\GH���m���`�G��+7��ϻ%͕��ч>w��JYk���!�����b@��cz���NN�׹���d�˹�.v��CH�ӥfbaf�#���������c��k�>�x�t����$����)B�ÄeI2;a�&d�P�y�^dlPܭ08%�/G#sU�{���Wu*j.��u���M�΋%�=�L�w�T����k���S&5{�<�e��aj̃#Li=׶�;&��uX�9K��;q|��J�����s|ѝ\E�E|��on�6�GU9˜/\�}VB������w��V��+A[�o4��r;�Qj����kj�%o�t]b��#8TSE�O.���1�b<���_^��u]��"�t.VRW
f�7ʲ�qG{;�SM;���h��$[�ӽMJn�ͺ�\�w��-ʎlov�tUJ����*�+�>*=�� ��������I�L�0�o�����*Muf\��Jb���.��U�s��]��<ޥy�k%��Αއ+�֣�[C6�����{�.�4,�9��m�ިGi7��egp���G9d�ݘ���)�[�d�g������~�ƴkZֵ�kZ5�kZֽ��5�kZצ����k�kZֽ5�q�kZֽ�kZֵ�k�Xֵ�kZ�ָ֍kZ�ֵ�kZ�Zֵ�Mk\kZֵ�mkֵ�k_5�kZֽ��5�kZ�ֵ�k�\q�kZֵ�{k\kZֵ�{k\kZֵ�Mk]xxxxxkXֵ�kZ�ֱ�kZֵ�Zֵ�kZѭkZֵ�h�q�y:8���9<���@{���t��J�Ʀ_�X��[QD�H�3˛6�-T��1/�)�6�ӹ�0>��J.�$�.����*e�B������{δ@�^Vc�<B�-K|,IO���U^��a8�����=���'E���K�w��N�%�]��ޱ�N��J�1��P�I
�Mೈ%Y�{�Mv�Ƕ�r��s4S��� ?�=K��2���{hH�-�ZM�#��#�{���l�l	���n�.Q�bb��w�ۻ۸��\�ډp�kJ�m;��1�=���}�EX�����MyF�bĻ�$�,t��è	��,��A��ˣ�`������E˶�D�Vc;>����7A!.F�&BS�{l�G'f�o��ѓFI�ʼ6D�:x����Q���tǻ#�R$w��CU���Efc�ˢų�xp�����a���
�]�E�$��~�[@�������3����b�ɹ�r����c������ӝ�H�ͨ�90�:���,e�qb$�vڗ��.��"�N��@F��-�-��}���-��q׸�(3Z�2,�>rfҽs�:��<�`ѤB�Z��)�K�v��㲾8��7H�����4[u���G�N��J'9��vC�;E��U(S������Lc�F<;�#�P�nc�noT���z���87r4�Q�j���e^uv�	Q��!v�3���6�(V�Fd�fkk:��Oom^h�
�n���lU-�Y��xLȧ��>��k��у��Mu!W�����Nn6�*����,v��5oy�q>�ʬ�SS|ļ�ȝQ�u�an�8S�ݶqj��tԣJ6�dq���,RgL+EsI>� #�u���z�7��i5XY���:.�9j�Y��l�E4˾A�^���A0�ڍVru�!���8�
Y�o^�D�����5 \q+��I�c�QV;�UkFk�z��On>4^^]�j��)Iu�l6��ά�;��<�	�<�2b�
ѭ%B9:\1�K�u�5��`죋��2�Y��ۙG�����:yUdj��6��3�`x��{6�2���s�+j��%s�
Dx�wd�:�Wջ��t4�F��o	8c̉��Z���N����x�3kc���gt�tu�+���oR�i��o��@�d��o�YPd�(�oZ�2�C��>y鵥�N.��m_^G��uu6��� �>n��v �#�����tm��3�s8�iܽ�Ku���@��Z�v�'n:����[�]����T%U>cr���RTڬ�ٝ([z�|r��(�K��;7Gl"r*4l��a�[l��?��+$�u$��uL�ٙ�MD�i��;w+�d�Zk��n�8R�P=}��7t�䱘��Tpe,\���"��8��q�6��.č��EM9���ӎ]�iG6Z�M谫�)X��U쬝v렬�a��b�Nۺ3��������*W�x�j�ˁr۷&q��u)
8��׍�/5P� �J닯�vs8�Ɯ�|Mz�^
l��0��z���p<�[$b��JWH��8�՛���smRִ����~��쪨��Tw��E	��e+.�s�S�jF�L��oX���scn��d�P�S��ێK��heΗT;�y(�e�;��� N����aU2�����,���ǏCޓ�/��C6~������'P�n��&3ŋ��V5�S{)Pªn>vc���'��tt��t�{����V��t�h���1Y���>�z������E�̪��Z��F47W:���vSv��33`�-�J�a(�yS���_'1K���p}��XX^�.�F�m�=���*�E�����d�|}�
�d*�
��vͪ�h��b�]����X̭:�'N���{����v]�;~��b=�H��\#������˕�LdY�׽ᖎ"�vb�d�����U��<����̾�`�Ɋ�cٶbё+t>�a�\���m�;���,T��V��3K]�s��c3��#]�
�l��\;�ǭV�}��t�o��/����1Y�;D��S�y���X؈6��Gv�R��gv�j����XC��8������Λ|�=V����Y���&�<�e�n�Фv鯍ZTݯ�çգ��q>�O���F�n��}w�9'/�_��E���� 4�k&�h����WT��{yUE#ts������ {^l�.��)�<�՜_]Mq�����c���;�Շ�g[�M�N���f��������E�:���C�ȕ���]7���u����%�B�C����=M\Ah̳��2\[C8�e��R}��4�3�nɥZx���)��U��YCD��7�`3��Rʹ�k�r��˝�^m=���|�����ܴ�  q+iR�\���^�׫�^��F�����4����(�!�{w�7����j�ޮ�O�ǰm�G�0�A�+�m���1��ra�f��7�)�J"������lug�KP�d��*�W0 4�z)��f�	���3�$1m��	��Z)h�n�����c�!��v<�X�Knj !�6\;Œ
W0*ǻ��Hl�.mN��|��\��&�(������t�4J+��\i�сM-I�X����{>)	kY{e��,(��b�ԽX��p:�r�|�%%��Χ3#e24��Q��$:�l�en<m�v��y_|�~���r�4N#��8�˚��꙱*l���Mt�n�|�vs�X}Y5,[v�4��˅��e�����y^g��- mv�Aj돰����R�۷q.��(�vЦ��N���Y����|f���g�n�}���Ꮫ��n���N�����5�^IwO�4�t]m�hC�X&J�5۲�Y��S��4�\��1�Qʤ% ���gmE����I�����Y�y�W^a�11����ǅ(eJ #���X����9*ĺ^�H��ӈH�|�OC]wC�ô��Fk+�P`��8f���o�4;�&��V�!�Ct_3��a��1�����`l۞�Í���0�hQ�w'��]WY���J�qܖh�m��-z{�U�/y���]��|.H:.YN�_quą��N���:�c ʔ��:�k7Plf�*LQ��Z�KY����q�v�Iܕnh���Hy��l�0�k��Z;xB����f�P��;(�#쳛��)�.�;3%umИ����D�j��+<�p8@�\MS�]Eτ�Ǌ֍엏�1i��H��-�{ڼ���fV��|qc�ޔW��)�D��6��k�'���e\���3=<[��-��;�n6a��Xgc�KFZٶ��{���qg.��2^�C4�S�Ƚ�ҟ%T) �
cT��_a���=2����RR]A�gJMܓОˇeae^t��l��#pV��G�=�v���y����R�D=������"��a�/�FhVm�R�sT�v��9��vWQ4ܗ���9vu|YXI�0���Rb�t��Wp���䦖&���/X���H�}��N�2�ݪݼ�,��D���[��O:�c ��]����l^��:N��C�I�m�\Ş��[�V���Xx.rfqo�0*��������SJLĢ{��*�p:��.eJ��������	Zt�N���n99���؄�7�J�l�\k������#�B�Y�����}�Y����6�[������*�O]�n��ۆ1��]�s)����Pَe��Wo��ʮ[�� -�����wB��|�u}U��O��fY�˻�V����A�.ٌ�=/	 '/���q��G5.E�t���ʼV���{h�-tXf9���
�X��kJ�s�ﵱ�YX�5I�>�L؁�9�p�jhC����D�ݕ׶@O�|2^o8(���`6Y|#n�7X�eVEޏ�5��$�ʲ�m����I�t�:qb�j�gf��� �t�ɡ�v�ƑL�v�� L�]�lo,����uN��Nɢ�M��3!�^�L�o+��aW����r���-1 ��V���;m�4�R:���g;FQzhӚj\뱝W�&��Jj'6�z
���Zn�Ǜ���]�$���z9��K�^+0��3Fa���f1�zLdK��Qf���3t�T�?]�3���r�nb�oNR�yM���p�K'�9��z���@�s�Ts�K�[S�j
�Nr;Ux��9��+ ILj{3lg7]�#9�j�q��b2�7���@�+ss&�C�-��h�4˄Y�{�y���۹��,"�;����GV�W:� XT�]�(᝖E�[�Z!E�S��#������9W� S8�7F��7!�;}�J���j��M�E�t���$pd����O���LN��^L��y\U(1fcR�W\�rTdǆi�Dʕ�`�	V�'Wwc�K=�6r]�1�gR��k-��$;�%K�i�/����]Az.bE8�cM�[;zTd�^u�Gej��f���,�q�΅\�sf��x��Hh��o�>����d?o���������/�����?����l�-���F�%�R:�DDJ9�O:�QRD�G0aY��Cwr$p�N5B�U茐��a�6�4�J���?��y�oOo\�2E��M^���m�ga�Ɯ��SZdlөŧ�i	
��y��<b�+�ȋ����7t.�_=��q	�a9r�Si�:��=ި�Ҝ�iG�&��Ԇfi0P�v��z�eK}O)+�,�A�����t�V[�y6�!�t`}��G�3����>Z���Ve����4��j�
x���u!9�N�j�M�r�7���-Ь
��/a��
�|��{ȋ�Au�6��[7m��}Cc��:�;�.��W9}�0w^��_%��F�,�������k�׵}��!ޛq[�l=w���=�tw0[�I�M��s����SכV�!q��E�9k-�Y���ځB�D��w��u��f�l�²�H�C	�^])��4g����K��6,Jc;���uS(�'.�QD�>Qϫ8��=�V��Ik�d��g`;�R�`�kp�R�
�S�5N�Ń3e����E��SNs��"I���L��fL��m��b=9`阂�P3.��}�Z$�å�{Hx2������I�צ�����T�4��-�/��)L�OEm����{r�h����i�BD�p�F�3���7k)��K���IJ�RI$�O.��:p�e�?]��($��@�$!�㤪��".#
8[;�sbjC��^%@ąU�jQ���n3
�%#H��r�?N�WPR@�T
�I
�HH�.�����A
��/�LF LK6\P�܆@DF$)`$�	�H��2�@���YC��I�q�Bk��������kZֵ�||xk�˯/D�|.,b����Xd$D�"Ø�!	F���OM|{{k�kZֵ�||xk�˯.�BO12H��^��:ܠ�IP�4!$	 B��5�oOmq�kZֵ���yyu��90$�P��I! ��U��>۟��_s�No�.���wK�b����9]'w#����o׊75��߮���뛤����������Һo!^��^�tn뙲�d�D�k��7.r��y�T"��wmwp���R��r$��1:w����uݫ:���.���myӘ&�];Z�9�����=wz_<ּ����.w:w[䎝Z�9Z���|�.U<��]�������D���Wx�5Gwm.nKe�<r[wy(�ӽw��juw���N��u�5 �������+��܎�G��N컥]�{���!0�������L��2$�!�`�F$:ܳ��u�ha�9����iM&��\����}/3^wt�vr�����/�.s��I:u^.��ז����/Ϋ�I|^���zm� ��Y?'�RH��R�,��gG��8�X�\�#P6\�R]��D�:���jm��,��vk�O1�۷��Pi��٬�݈�)"S`�d�MٌɺN7M�3!8�wǆ1�`�<Q4���3�g%�E��6!y�+8t��s8&:�u��~��㲩Ƚuz=$��L�n�&�3]�ΜI�g�Gm{�F޻�����wOp��/xOP�pc����E��f��&�'��4U{W��0�����;z�MSgS���n	=����R�I�Idey-�~�!F�[���J{�V阨zǸ9Ԅ�?^��<Vu_;㓽�^�#X���������t�����x�Pb���(aX��i]a���������}��|�x�<��>�=j����7'{	���ļ��[�����cT�'�Ϸ���t3ݟ>��h>�s�U�&�G�����$r�9�E�]�Ϯ��m�����ze�eC�h}_=�~�Z����;A
XR�gF���g<�_Z�B�w*�����CM��J��f�}���]&�tm:�=,��:{���T-�vJ�o�a��g3�ޚ���{�닎1@���z��8�i�}q�U�ca�}�BXj���/v�<�KP�:c�9�f���>ߏ��~?��b-�rv�o�~�Fm�+��=Բu�C҃ �R��j>�Fn���ñ�9��vK��U��l\N�k�;��π�9�œP�c��q3WB����'b��c<���I�	rC��G�cjᜉ�A�؟eI���&�잉o�������� ϣf�lg��J�q1���|������c}�n��}~d:����w���e���&�8��g�� �Q�b�t�Rt~�Ϻ�#=����G��������Xmʏ�J4E�ۆ{w�����+꜃>�rö�?W��9��@����?�p\���(+!�n���ϯ�����m|�)�@q?/�����!����Ûݯ6����e{Q�=S��޷���B��^��3�##��{+zfv�~�:ox$��g�pٝ�a�︎�'s��}^��˃s-�H�����J��2CT�z|4t�C�ۻi���c�YKv�Q��)�"-�38UU�1p�q:8u��<��N��jѣ��U�S!��p����/9}s���󃳪ʑZˬ�!�r�ʶ�PKe^ofu'�oSι�w��J�1#:ͧb
8�/>�~�3�.�{��\�y������;�"�L6�^���*⻿s�z����e��c���F2�Gu�	��]�y���ll���5���#�����pj{F_��7FH��73}�����gs,ܹ;�~փ�:�l��S=��8�G�g�=
]����N��f1g�=�bqbC����];^o0KO���?�_�Z�P��~���d�'�/�=�<�;BA8����M��������9�W�����>t�q�+s=}=�8��f7�49R������;Ԍ��ޫ����K�}�&���տs�ՙ���
�}�	+��*݈V�5*����t��?u���
%�h��W�c0�7�2(W��x&P�(}�Wޯ����i��U���l�V9�����~j�B{�(��9�,l���ׁy��.�?.�I3M�VU{Ϭ�`����XL�fu\M�1�8��+��mkE�Y��v�旐"ۆ!ٍ��lN�U����ޜX�+~�x:_c�W�wm˽b�ё��2��L�ڻ�T��n��3I~�W�ᵥ��JD�5FᾹ=6�d&���R�}��pG�:&ދv	xٝ���|>��^H�=�'ݏ���j��zM��sQ��i[,���Gs;�=���_y/���̗��`O,�]�?}o���sl3��B�%�d������Ǿ8o|wgg{;����Z���_,_/� �N��h"j��*��h%����'}<�G��*ܾ}y=�S��SOt�}��w�׍�˱���zt/:�R
�]y�+��}�/^��-衄V��>����l��֝�1��91U��{/�{�`��5�ǪF��]]R?P�ТI��}���>v�ۮKA�N3�Wa{·���<|�}�אS�P�9|��iٙ~󇽚x���2P���FL��=�oA;�f�Q���X�m�|�잢Fk�}�7�d�QkrM����5d-�~���ڏ�|�@G7�e��ߙ�]=�{���k;n�R��R�4���Pn�]%D�׹wƅ�4$8��l�b�������t�B��T	�0�*�Æɴ%^P���,��65�bsm;&r�ݻ�T�;e�X+��6K�$n+�unӪ�upǣ7%fǯ��}	
��&�E��`�i��e������dЭݾ�3;�f�%.?0��8<���y����M����>��3�*����嚾�h�ǼV�:9`�O�ͦ����m_5G��3#��]����4�xOJ��G���%�t@�g�w8�R�w����{�s�{��ϝ��i�6{�" ��;�����m|~�����z����ܗ5�m�������^#��>�fk��.��=���}ǯ���=z�M~@e�h9�t�o��L�`�U��OGP��G}�\]����C�����UT��3ݵ�������M�Y���������){��mKͫ�ӳ�����l!+��{�f�W��?n�~������,~1�N���j>�y��P��>;�-TnN�0��f�<[��<�w����= d͐;���0f���4��ϴ`���
�}���|{bWƑ��.iI
�s�óz��+�����!5�ip7R�Nn=�˳rʤ��\x1�(�,'0E-��7�VM�
�N^�����s�K�c�Kp��⼝�Hks��f5ë�*�����||<��fmKq�H_���ϝ�Ѻ�f�?N�@=<fu��+¥��0�<�}��]�$�u�`kStI�u���M��r�msk��[�bj=�0��(#C�����`���i�o�zT�ح�Ý�'_����y�`ݤ��zܼ�^_Pa��e��!m�������WX��'W��xzߓyC<��I��*�
:>�WL��Ѻ��芿E�}��=������h}�6�B���2(�<�{�7�;�s<��xg�)?~36�ؿ��2nW��$�BHnp��Gκ>��F�V]u~�돨G�����MI�j�/9� �<'÷^+#��b�B'���~�/��'6J����Eך�A�t���n"���4g�[5˘�{��������Vݞ�i}DH��/�o�i�����{��;�)�ݬ"�K��
�\��j�i��ml�壖�ޑ��K����������[��q
7NI$�����]�萛KbzfӘ���*��b:�#�N�ƞ��_r}}��*c	�d����Q=���������r�;Ν����2Uծ�xy�b�|�k���;���vY�l�&rD�0o��L�ڿ[V������G=�y`Lu��M�~���NE�&�}�=�@�nz���u\t	�s-{=���4��3���=}J���Kg�.)��_?km߽�fzx;���0d��-�gՙ]�p���y��*v{�Ep�,#��� >#g���c/H�����c�����y2H:-���-��i>����{>��뿶{j�?��Z���1�/�c�w���3���U��3��ל�v��j�OW���Wm,�xKp�/���9��Ǣ�'��SW���Y�B��=�k�쐥fQ�{J�^�$��+�Ҝ�%�}��R����6��¯Ux�]U��+r�T�	��}�E�w������̈E��ǒ`�F��{��vg�U1�Vv���ty����Ou�}�j�kX ����Y��>�q�!P&��[ݔ�j�����uu+�Ψ�>���F��)؟V<�8�:�'Yˠ���_���ٹL��U�a4�-Yݶ�\��[���� �@�sj��������Z����퍙'*[�8\�2zVk�}��p�k��q�{��S	@��_�u��N��B�걘��{�Y��|�����P�V�$ʓ��F�J�@��ne�5�0�����^݌Þ�}}��Y����?9�>do^�$�0���c�e�uq�|��|��W��3�r��T��/y�� ��̞�X{co�����b�p�b�]��^)�r��>x{@��{�r��/޷pD��=���Q��nC�/)����|���$���A�x�xϤ��U�u^�V�{�eW���(T�.G5���|�5�"�� �[o7��6��{j�$W{���9ܱ��+t�q��<����������%vS���u�H��x
n�L��c����V+O��<���]kv����>Α���6JB��>7�����O�i.���<�\�S��f��_
ڲB>��x����Wcf�̙���ܦLU<0�T,��D�
&S�&�o �r��S�y�1�n��񃇀·#��cM'�ד^�c�o��N��櫤̽�6��I0����.��)�P�a��,�;�������ˬ[;������`G���M�������J������W��y�0̮������(��wM; m�U����y�c5'3�;�]`_T��t�� ΂���π�Y</~s�q#�#�[�I�h�;�S�n�߰�$ٲٶN��z����pn&��|���9^��i}�ۂoz�l4�"�A��'��@3"<�:p,�����|�����۹zߍ	�p'Ns~�H[׵/�u�聿f�����P�D��37�Ά>�٥������Z���W[�3��X3DDum.z[��� Uv=a��"|r=�k(��<�z֔�v�Wcx������;~^{�Q�B��W��������͚��Ճ���v�wC�'��oD�A�;�`����du7�f���7���L��Rc�;��;M<�8���7h6�ZB��D䮊���Ң��й��ۇ.7N�̃9�W�Ȯ�*�3/��(��b�Ы8����O����۪��.giy���;Wi�*�)NT�7ۂe��r�vԡ�AW{��4��U)#�̅�Ӿ��>>>>>��8�p�ڻ��I�x:�ꃝ����y���l!�d����;�4gu��*k|(�����t�K�z�����+����ײ�`t��ɫ ���'���T�(8��P�B�u�����c��;���E�ǪLQ��x�l����}!�;K�ʑ7NǓ���<-��e�6@������������ݩ����g8M�v(Yj�<��}C��}���/�����RzY���X���=���'�l
B�{=�9���H�
%r@�{�¾�h��vn
����i�~���6�=n����g�8�)�e���_T;��/`!vu����s�[󧯻�4��S�}/3?vH�����P�â��]0_�ݴ9RK�L�:��/���_���֪ɪ�x6����khh�ÀB�ݠ����.����y�j{���{�qU�4Ы��;���%t��JF�Q6V"�B^�y�C$S��oEx2,tCR��0�g\���_)��!YY'`v��V�<:,_nb��]N2�'k��rЎ$P�Ju���h��,��1eJډ��𹄕i�Sc��qa�@ދY�є�)B��%r�ԕ��܍,��gv�l����9N�n��34��s��*sVI�or���)�a5g=�������3�m�v�LF�.=ݢ��c˥K�]qo7:���Iվ9)59�����TWn͢�����7y7ίW:�(ǯm���޷����gj_9���\�7}���w:�]H-ꨯDӴc����[Xs�D��31��_VS�^��z�j��=j]#ׯ�����1��ԈBĭ�fU�̺D�
Dܸ���g���(�es��е����i^��;�B���O�m6�d�"�;7��&ӣgp0��Sm��O4����J���nP�rԻ��S�� ��w��������ʢ��k��^�,	�ۡ=�r橓8hӖ��3E�&m��Ӫ��t�ki�Tـ��q]E�gI���(����d��M���ܤQ�E��d��;{����.ѹWj,���r_sV�1uS5VV֪Ζ��6������M;3�S;�73h[���WAH@��j�4��f�l1����+#-�-&��I�DM{m���V��;s[�/�᯷ݷ���!ؑ���]�+)0�6���^u��n��;1̨1U% �ÚP�$k����b޺[��w�ӗ�yֳ��rub��>��
{]VWI�b�Jޣk������9��n�ws����1ƞ�M�c��}z�&�g�c���M笙�g\���8^Wr�**=��+X���r�t�e�����7_ť�r���N�ўת���솹c��]-���u1�ͦ���Sէ�(n&ڊ�Ek	��dŽ��Q�5��k��r�#O=�2:�Y{�Vc=��!��2U|�b�v��(H��^�����G�<��g<@�E�&�ṋ8���D�B���I;�!?J��/ 3����U��o=a�&�:��������E>��Ƈ�_l�� `�$�E�s�����*EqVB�)nv�B�����x@��Sd���B�6���oz�t"��Ԭ`2�nh�f��Xc�x�8���L'e/=\�V ��0�k�Ï��;���n��&��K\m�}h��)^9WI�ǯ29v��+0��,sm�=�.��oo><�T�r���}���}t��i�Bd�Jꭉ��I��d������^�!ѷ b�U��?C�;�[�����&_�W���22��v$������־�5��>����||{{}}}zzu�8���iX�o_K~�~��N}NG�s�+2����{[�$���}z|k�믯�������o���ON9	 �$I	 �w6MIQl��휨Ą������������__^____Z�Ƕ���=8dg8�9����N�V� �5�~?��I���������)�6��wa"�f�F"���o�;�u!�h���|X����A^�6",��I���W�����D���k���,O]�(����(���aM���Dc~�PR����h!&o������Hlz�����cy�S�M�@b�џ}�"�˜������ҷ���~Z[�왽����{Y�:�ˇ��I�1��y6ؾ��Pn`��=\�^wi��)^u5�:(��//!��g�\�N�i<}�����}PX����0v�~.I�3>&]��8����j���xg�cj��[b����q��x�x�0A�%��-����p*^��_�O�]�W�W�d����y�F ;��f-=:�#3ڒ�[�����hp!�yg�b9��'��\�ǀ�y�щ*} ʽ�Tܸ�'����"8F?1jj���I2�����V:��+�O��O<��~@o��L������3"!5OK�[��S,��pi���3�����X��g�u��#@o>z����w�p�\دM0��B��*9k�jt���U�y{��������%�=�f��H��@8ͬ+��'"��Ϧ����.,i9�[.��룈��k`���ޚs~ȯ9�eo~~�oV��eE*Mmp��}�Wld:�`z"6�|}��T���d;w�����N}$O�XF�����E�k�����|�LU�H��I�c���}�fj��g��{rx��y���\���3�����A��l�.Ҁ9�ۑ͞U�����N�����aw��r�j ��*<:ͯx|����6i�$�=���v�81����S������ܟx(�����F�s��ӣ8�<�X���T+G�W�[�	n	sy�ٽ�O�q�J���I�I�7Q��%��z=���r��uI�N�y�H����B!p��b��L �	J-����Jw5�2B�O9����s�o}u��3��n.1�Æ��޵���8~
��g�yQ���$S����t/�O5ǿT����[@Z��5t��+�n����nh\��	�����dz:�FPp)��v����cG��u�7�|��n�g���W� ��A�	o�f���h\�^:�=��~g��ϷG����{�m�����ਥ�K�p!�5�����dŝ�����n|�����۟��0�m���$�_��I~�-@ߡ�y�=�6�������v��&�{��	L������|�	�\O�c�Y���$��0�Zxð�̇�s��hWzq���>� 
�VWA���b���b��1�1�^�������.�hEn��i숙,�c�f���Y�A��.���Q|�x�`3_�/~"A�?���'��~���+�=Uo}���ddHWT�fV6��21V���-A}r�c�� �D��v�4�zw�a������B0.��(�f����������`��U���MmB�>��&ˉ�~�7Zϯ��0�}������ܯS!��WBoz���a��c���u�O���oCd|�~�����$�Ta~��q�=�bA��q��SB��-b�0�}n*h^ 颮��pw���#7�y}���ږv��M!|���-^�H�#H@��A~�@ id�B��4��z':�K�����P�i3�J�U��h�GM�g!��o6�s������gF;��u�{��e�@BI�ȁ�'�$0�m��i.'�&��s�38�x`�c��u@�u�4�0f@y��{oe�ċ�L�����_ ��}�f�ݤh'��ov�m�͙D���WJ� ������^�6a�6�,3���F�����C�\�s�32Bs����	�h�o5O��g�74i���=��`J����K��~5A��+g�؛�7�_i�q��U�	�E��	�o(6�t�@P�HM*,|�����������K*ʺ1�~�5�E���O� ��7�S��U�'�X�BO�( ��J���4��`,D������6�;Gk�?T�r#J�������E��L���<_��ĩ��z���X�������\0eCz8�\)���f�W���si���6�7!05�ٳ"��������'�zc/���\�{����g�껭�x 3X���}���Y�"W�]���7��=5�`�������W�Y9��Dw�we�#m�~�1	��8�T
�t�@cG�.�(&��d)v`
��c�dWc���8�9G���H5��5���x-���7��|��{@���Y_)�_���|	$~�
�$_�Ȕ�fގP>�����0�=���K5[�Qt��%w"/:���n�gkP��K�~����jo��vmC�C;2�(ZP�&���Y����?Puu�ûr�}���_O�Yz�\F>K����6F�+�Η,auNG����j���m�y��\ޘ�{������y��;�`.k2�袗��fi�g��#S�\`�	2އ��-�����@dg!��Z��ҁE�<�]�x��}���TZ��m����3�^Bj�7�E���o4��i�P鋇�m�)��f�w
�1l�1�Y>C����>k���ǯ7��J��
m�'*Go�����z����}<�a���w�ڷ�YΗ��x���ρ�/|��
%���:,'e��%5ؓ���g��	�
O+��!�| ,��N�$���q�n?[�Z��h�J�/G0,�C7m�ߠ�ԟ����j�Z{A��}Ï�<����L���J�o�M����<�;�𶀝�p��cÅ�[f�ĩل=�	�l]�.����x.<�U\��xd�L����G�����y/�ϸ�t�˹9/k<�L5�"��Vj���Fu�XlAd��%��wEL-�]ctS*W<X7��~kZ!o�+	B�`]�7��G�NP�����4s��Ƅ��'u��N�{�s��}�~�O��(,h.��IĶ,i�h��@���]��x��|�AT;�y�Z�#Za��������4}O�T�r-@�(����l9O4̑�	�w�f]O�}XԶ�zp��^��/Q�u@���>��D�ٷ.b�����9k�q�CF8A>$�@F�����mD�����[O�r��ĵ�`J��}WLhz�՝���A �Vʹ��1����q�����y}ݟ�����|��v����8k�N�%J�\S|)�����V�0X_��Pp�_�LKb���`8f�����μ�Y8�#�b���yx�c�՘��jdet[����p��~�.��GW�4NZ�������>�u�z�˖�{;���P/��u�t�_�H����iݘ巚��gb_����!������Ѥ'��V�C���5<����pS�9���;���<�C����cI�� 8��w���+��D�J~�k����cL�x���\!d��/���|#�����v	z�A2�|�d<��0)���^a[��ם���`��/��t���v�@?A���*�S�L�e�����??ut8~ጛ�PU4єw�;�%瞚)��Y�X���0�Ӗ�7��ZZ�R��f�Cjp�51���'^�c!{��ͧ��b�z����V _h@�yOTO�|�؇�B���76!�����Z�|j�x��Mxc�s �%��cz��Ui�UhW��.}��2S�"�߈~r��)�:�c{��y��s59�a��ȹ�V*�Q���9�=5���H0���j��`�[SU<�L弽�$�̼�C��|��Q=^Wwi�Z��o2Hw��ޭy�{����볊�R	�2�����d��ѱc���T186UPƸ��fM�s��;�e2���aZznqՊ��V�vt{�A^s;bV�=sK�^u�7�����0cPȬ�q������m�TKxEtW���4��1/a�=>f=	D	e��I���<3ò.tOD��dE�x���|���H���ب�
@���0��J�|�LU���T�Ia���ni��*�Pט�ung�.Z-%�x��x����=�!�~��zǨ��Al?��|`�|�_}� �Z>���^f9=�ꅵ7}})x
�ݖ�
�uz�f���s��, 0��$L#���?j|��{;>�V{>{�+�3��1��]�4K�yf�-��������� �cU��cg����42n;2'�f���b��q�j�>�#��cxsJ��M|_Г��=����O�D��-�����,#�>������y�f��6��;J��_%ץ�`�^�"��^�a�V�ط{�H*^�8快�ZDGX���gL伜����l|�|!��!��=K�y6H�;�ڌ��u�� Q"8y��m��m�"����uR�ow�����]��S�8��/
="��	��Hlx�>,+�$�q�n�x�GOb�` -�,�y���p�Xy�l!�
��xE�x�!b�q��*j���?� �`�B���7z�p���Z�/&��ME��F�0�1�D`=��p͔(�ɯ���/��-"STu]�����C{^K�%�$]��xކ.l�X�s�k��,]�Sa�Swh��e�.v�3x������p���w��L!�)�U1 I"�jp�R3�|L3���'�X�1�8#c��E X�����ߟ\��w m�M/}�?5����y ;Ip5�=sͼ��(E��=�z��9 K7�7]�"9rdM�e�<�w/�콦4��Y��o/5��A��!��i�{��[D?4��c�=a�|�A?��.~v{P���/ Zu����ג��֔�}ύs��A=⁞�-�y��g�Lu��y�ý����5g
�ڵ�t6�+�OL��!5�&/mq�榺󁞋���w9iW��$��	d��f�L�u��,X`���l���u�z8�Uxe�Ry�"�0��	����Jui�J���g�H����G�x�2�}r�ȶ�] cz|ڽ�?��rH����}�ϓ&%��#L�� �w��}��x.9��rn�z�r1�a��/�;�P�f��~�B/�5A��+��l�5�Lr�^��fcy�QL������~�o*_�W*K��iQc~a�|�!���L+�a�*q�@�{�ec�/�����Ĕ�oq�L'NN�������ԥ�jxw���|p$;��];��7���ڗ���sB�֞��Rdt���qq�	�&�l�8f�eg���B{mniwdԸ�2S���u���d���^�\ڈ+"Uo�-���7�G�����q���1Sk�U�I����֚�pI��k�q��vpG�	��v�+*��Ɗ�SnL9�[�i!!�|�č⽪��)TkK��eդr+��y:�� }���q�"ヂ��d;�il,X��-����͔������f|+���ӂ	�Z�ZPK�_�G0�:�I<�s���BzW��02�����y�A�8lN�2��`[���Y��}+����v{D�O���.{�"e�	����h�恞� ��>�M���O��L�K���+��#�N���j����f5��z�,��Ş�LDS k�[9y�ߢ�� `�Xl/p�ay�6���9�o [�����Y���0>̐��k&p�j�f��V�[�<1��f�\C��B��j̶�Ɗ�ۇoSYu/V��-퀋�I١z�3����W����累ƺ;>gbɃ_Տ�.בOu���w��)$Ixy��@��ܯ��}*xQ��E���Ɓ����� 8���W�vn����ϣ���w���ª&b�_��xY�~B�>! _��[���0cǤ&G�7EeW;9���������巙��1@�F���o��N-�D@8��'�I�Ѽu��˗�n�Ҽ��-�/�S�f	�q�
Q�x�5�<�p-�C`('E�ǂj�az˅��V���愞J�����Df:dT-�m+�/9�r�5r�te�6�6���_�{��g���T�a�ٕ~V������ږξ5��'�T�%>�V�ŕ��i�������f��m���f��I7��j4S.�����'�qD�LDG"���<=�{�O��4��~9>�LzY89�X���)�z�2�P~���r'�� D�#�9��r��M����xb�����A�
n %�(�aa�w��4E2�-4#�`˖C�mv�V:�(z~k̕����������#���0"-��J�Qq�c����5���=�[��{���0�ץײd��aE��U�/�����0>��>g돏�{^�E=o�ћEQ�����4�,�U|!� i4w���yo{+i2R)&���#Q,m��8��*I�����O}?	�/~>~An :�#�>l2׳k����L����z�p=-���b<*��)��_0��V�썚�?i$1^��D��9�e����T����#gŁ��7�c`Ǣߋ���0<z���5��4t�!W�{Ѹ�m--3��ڏ�,[yץؿO�5�Ɨw�=-�u�H���-^6!�ׇ|���qz�த"�{yxX������X�X�2| �[i݄�C�Mza�<�q����s/se> ��9AD����A�C��d��ϭ��sc$g�2�o�-�͂�}j�����3I5���$��)eo�"�tN���-c���G��^P˷Ҝ���9'�k�����ܾO�I�?����O��V���H-I�	@�}o��9�Ko������>��e����r减���h*@�3j�+�ъp��h�S���sx�<�y�V��������v�w*�-��+j*���hՊ�ccQQcQ�	>$�!���������\ׄ�]�߀U�� _�v>�F�?����?��=OM�)��-A�e����/��ޱf�]s�^��mC��jH�x=ٷ�t1Y_A�R@;Y~�������}=���8�Յn��@i�]Z�xnO�344/�Ꮷˤ�����hL�3���1�4�[{��[�z��3����X�aq����'3U�s���,/]���|f����e��	c�`�4��Jg`��0( ��Q{g�p-ޥa�8K��m39/ E�A<c�mxLk𬁢j8�1�_����S�L�R���r7SլkRWf�q���z�̰l�mB˜L?3�`�\s{�wI����LU��|(�=��.~���:���B�3��Z���t����?�������՞�&�ضR���̉�]'r�J��{:�x�;� A��c��7C�)���vG������F�¢�R�����=[��M��5QwQ֏/ M@�r���h��%���;�r���~vFx�7�*�v@�`���n9ya�����:��Oj`KkzDi��c�Jp���Ũ������4��ZA�D��i�x���
���<s~�_�
����g��uv��ڼ�ȶ�U�wah�:�j�Ի�t+�gk�5�ޖ劉����`ɗ�ۺMH_��L�V�Ƣ�<s�M=��
Iw�ɕ~ܝP��doj�GI��Nř�\r�D;YWR���g�ࣽ��&v�m&])��sj����X
���-�1��z�Czо�R#p���\�E4���:�U�Ԓ���KR�:]�f�ŹKb�]ICv�����V]�fHꃡ|�S7Ej6.AlXˮ��k+�#uPmmZ�Nq��u�*	�Y0L����ޘ��ں����|���l�:���ϬI�F���YIN��/F�(�u�2T�6�W.c�|֐�r�틻1B嚧C�b4�k�o��+^i�;�#����)�����ggM���uN���5�A��*�A�S��v�RF��2�����$9���Ϧr�v�}�l]�A�
: }1֩2!U�1ͷ%�ب�/LQݾۣ�k��W:7�',/z�hl�Z�lz`�Yp�Yxıۑtb޵Z���W���x�dk�s�wd�Ot�̷,Է>��U�X\&�nR�}Z�OIxU��w0���	��E�mw$�@fd�H�{Gf�Uء`܄Ul�hCKf��ϰ�UT�+�ttL��֠&�aor�p/z���.��Rz3AG*E��(Cl(�3*�Cʃ�x��kR�n�Vc��P�I$FT���p]*Vc{0�J�Y���atS�M�.���h��2|�0Z�d¤�(�Hi�q����|����O�z����Ct��د`��Wܔcl\����.;X�٭h���7���i��<Jq�_G��ŉ�Da�*���Ι���������e���'��i��ծ���\mE��ve��P-�ٯ��v+2�Ʋ1C]�û�'8V�C����V����DȪ�+3��W�6�Cd�ږ��UA�v��M����'ېG.c��bms�m m*r�kM�o0�/k�n�v
�z�Lef�e���2��L�t�u�36��N��l^M��e$vA��i�d�%��v�h)urot��r�E˧쓝7j�\VmAF�Πo�Iv��J�Մ���p���Kut�WV�WJ�o��E���e�������L]�645{�x�B�s��2wcN����\��G7]Wm%��%��9Q�C[�R2]dTC�����;pv�S�gJ"�꽾�zb����%f���j�M��ר^�q������EO�I���1ꮮ�!׃.1Is��jE]��'�p�7=��d���x��g[ي�빯��0n��\�.��[�����e�|g<��bı�}��eP�6��am��r��ʣ�6k�Ӏټ��Xx�2�E�I'd>�Nl�D"��$0U0Lb2�h�	!	�i�$Ai��%��&Ze��Ѯ��0XF����^4O��%䅂�"��ʒ0�m���b��Q��16Z�'D��-�D#TI�@'�n(�e.��Xf�DK��h���҂��p�Z@D�$�����>8[���X��ߛ�|ߚ�=�5�������k_�_^��Y���rH5��(����uEcEx�4O���}��z�����ֵֺ�}kZ��������+�k��:�μcQES��oѼo�������l��Oa�<zk���^�ּ5�k�Zּ>��=8���K��� �<���ͽ5�ߚ��b�,j"Ƕ��P-	���L�sc~9����04h��wZ�F�*5͹b4X�F�X��-{vh̦m��Q�w���ʼ���F*"Ɗ4W���r/MpB�=��،E6���x��WZ�o��ƹ�ۗ㤆Clk��)
Q���@\��#r�"������*faBQ�**"����U� � C��q$ҁ!���(7]�Ř���=@��q��X�cz�ݾ�j'�7i�$��[T5����N륷Z�ʊ&ZLא�O6aloq��8�&l̇���G! pq@D�z�����y�|Nx3><a�C�����-�-W�2�o�8ۯ����`��V��z,�yy���w��oV� X�8g�L��"�̟)�XG�B�p��N2�_��0�������~�w=��,h�b�s!OA�@ǆv�靰�3nX�����B��	/������[���	;��ؑ�ٰ���(�%Z�@a_����!�1�08��A� _����=|-a�Mq����4�ȅ�@<�P�H�e�`$ִ��6�k�>���Y��xH����]���9x�1��rY"����� �����&*�AFCH��@���Y_(9RO�??���~UI�ޢ�U�����}��T/G����@��R{,g�P��G~�Xʛ=�T���q5l*n\��#��[6���{h��4���~��#@?���2�ǡ����cKxR�TXS�Ƌ�������e��~5u�;j�A���~"��8�7�3�+)���?�����-鱀��M���蕞B��b�̲E�mS�XX����^�#Ðɜ�~��a���x}�o�? >�~/������a"�pdÖ�]B�����E��ûTk�v��i���ZBFJ�.��?�:B�pދ�9
sY9(�̒
�9�-ь��#�ꄻ#3�D:wh���gr�_6[߷��]x]JשئmeG� ��z����ܾQMȦ��<��>�ϕA��pEq��E�00��͵o�8W$�n��g�e1V�>��D��?=s��T�́�a�l��`=T��-;t���#k%M��KJ���'ZG&�p�I>x����}o~�/��,���C�J�$��>-�솽m,�,�k�Ў"ˡ/�l�����xU{�O<���:O�-J���z&n8O�4�leϑ)2����{����;��U�>	p&��l
�=����*�,)gO ʬu�����\CI�.=]��w������ ��qЛ��.1�ّI�8���zV�������O�f��=>��{V�e��V� }9׊�O�ᯈ����]2~�%�1�݈��ΠT��C��F��y	I��.!��"4x�o�������;���y?(
}P��PU���
YR&��cX�8���
I�@3NvͰ�x ��0�נL��ǟ�漻ǐ1�/х��t�f��)���1��P��C0�w�+v�	z*>D�0ߴ;0N�~]X�	�sEҜ�����i9������$fA3�{�E��з��� ��B�O*��!h��NGS��xO,%�,W`�Yӎ�;��M4�E�4�T9��K�J�%G��u��I��m��]�t���e�	��pM+p�2�i�sj�r�/guY�nd��hFqlbeގ���M�c+v=c�W)�owםw|���=���c��*�q������:�x�[W�2�������T������ѿ���0о�ux���+*�onNf��[Zx��:���"��N���(��D,A��B�_�d�'ϻ�SX�N�O$�QMDfޟ9��b�>��τ��6Qb�+~W���3ߐ�}�$���#c��')FP��}Vݼ�!S'��H��D�`�G�l�x��l����C�oW�Bty��!;Z/�E�>���忹� �
s{�3 ���3<��<K7���2��&��+�w0�
��|�י��5tU�X�գ��^���v���� ے�;��œ�L��t��^[9i�`:�`�t;l�"3]��'bZrr�0�٥�6������`�<�o�lS��<@��2Qq ��}��# X�̊-L����.Mo"�մ�?2�Zs>�<�������0�4&9����<�z`%Uˀ��19�1��(��c۫����@���܀��o�a~u�ܞ�٦��#�G�ͻ�ާ	����9=ݲ���\�ay(�{oK](�1���ql6v� ���wf����)���Ӏ�	�GU<kIp��.�)���#ٮ:y�KQ��g��-�Ov�xK��V�9��哲�u6��*R�I�$�Y�,���{r��}j�q�8$w#6-��7w���c�n�J�*��KIi�4�Q�'TJ�����'�"���88��88���7�۬�.@3T�S�_�M���M����+6�Y�r����c�
=cj|Q���<K5�B�4$og.����
e-�@��Ÿo��cޡlOp��%��I[K���,K��y[�+���~���x��.�'�����@l�ʶۮK��� ����7�wf;7=9�Z������ �{��,�8@��. �Y'��x�sdz�D^��^��ޙ���ˣ{En��<�0+9�ʀ���f !N��a������x�-}\����5z��^����݉Ar�P�yٚ��̚�[��6+��VWӠ���!fz���Z�]Ǳ�9��֓��uS	��#���$�ߏJ���%����xQȼz��x/CN��L4�&<3�㳗El�;]��@�}���#X}��b���q~�V*������BzّGi�I�y;�4?�5��ô�/�ސ��|6xp�o���zĻ������)ȥ)���*;3X{[�[Qq�vuT�!Y����@~͑T���2��o�q��{�RO�a1Z�˻�z�����=��/�+��E
�n��큶��;���6K�z��إ�V�X�SJ$��2��Fi݄�(B!����Au�%�W/"���:0�DMc���g]�8�Q��<8�6(�B÷o�Y�i�׻x5ܵo:UC�ҹͩ��Nwq�1������O�dHR���7A97訾�A��GEPvɽ�������~*���)������gX�����v�z���7���������n�dxO�EJ�|�;ܔ��;x��Ee1��R�.������|9�o<��zi��w@~�a��o>���k�ٲ¤w_��q��GdN�v����4�(�z�,g ���=1/l� ,��:�4�5�R�6D	����Gv"�fZB�H�5�ڮ`/�p�}�y_¾�ߩ���x����f}��AbIv�:0H>��v����_[$Y�@*��Ϭ���O��BkH�ge�b�b�"b�ym�"F�NՎBÆp0Ey?0"=Ƚ˳y5͙��rRv�u�����zs$^�9�Ƃ0m��U�h��T�S)��G���I·�pY.'���vf�J���g9C�ov���o{ZAP�;�;z�-�����Pk��|S_�V���K
;P�w������n�p�7X/ c��a�NS���\��O�|kOC�m���`0&Bl'۶��i��,-7���4��mǊB������{�r�W-N�ϾX8ͶV@�t�ӽtwn�l��)���-;[�\V`��>��O��\U�2�!
ʿD*eS�lѓ�A����V�]ՁU�N�tɒ��Z�RĬ�IY�\u�d�F9zxӑ��;2���z|�˹�����ٻ��xd�N�w���s� �?#���  �q�����Y�:�����>kȇ��E��q+nm�ҺScP�oF��,���=6Ϧ:�4�ۨ��+�xZ=�oz��1]���z��7���0D��	�<�K�pͭ����;k���k����\���K��u��J��#�����Z�"«��(R.�y����Oc	M�A�qy��D��rn�jH����Q&���Rqo�L0nE�.�od����w����o!�� �AF{d�_���誷��5�$?FO6��,�����I�����}w�xa;~��֑���V�ۅ�uVj�׸[GP������Rd�����qQmE��=���c_��"A�d�9��[�HC\K��,h��;	R���0���/��)x �Ǵȝ�r�
����TG��J�;��
�;0�K�Z�w:�>:w�>��7����0:=������),���Uj�XT��j1�z¥]����-F��A�B����1�|cK���R�����nzV��o�<��r;cp���f������#�DR)*�s�~d��@p~%��(�_� �S��q��_�r���_)K)`Kk(�ˢap[*L��'q ���]C:�V#46��3��祆ݩ�E��
��Y^���<� k���s\]������Tx�JmNV5��� Uk�>��U"-��;�[�7u��vu�^���|>5�@ppPq��DS�/=w�9�%�����ײ��/�8��Lm�@@W��X'� �M@����诳��Z�`�]���.��R�W��eb�a^�OD�w��ܘ��7c�cW��o.�{����.�G#�6��&*ޘW���+�f*��鶊vAǮ0bLCg����yxn������ЅR����|�2C(]��MAD�,�L�������Zb�r��g��E=��S���K���4�v�ga�6��&2��� ��t�L]��q"�SG��"���1Yy'Y�U0, W(�Ǩ;Gb՛;���6Gdt���E<Yv;�DQ^'�|���d�wg""�������56!�AcK<�|bP~~����ȜTl5
����F �KO��A-�s'c���e�ؽ!�7�����{�)ՍRX&�%P��x����AJ�~#�gS��1�}��>�Ǎ�N>)�m���^�\װtM1Oh�2�i��ט2�58�?\ƺ�?�0��(��U���V~B'hub�����uC"��<�L�\�H���%�D��a_S[_��`a�.�F(��7D�qLj>��111[4����rX���5�okH��_G׸|�����xE��p�|.�ξ���/�󔊹�.]�_V�u�ܲ�U�4��x��ݽmqqDk!iG�S:�Y�es��}�(���8����*c������i����yo��^|��q��D��7f02%nM�;����j�:�MM��dT;�Ն���a���ah^��|���qp^�=�����SDZ	����lY�a�$"�@�%f���i�K�����X��x�6@}����S�Z�S�[�*,a��f�Cu�l���Ҳv�xqP�����|��le�y�S)Z!�{�c��?���w��"�M��v�4�/��͸�R�eQ�Ck����1~P�	�N=1�'�|'��ۤliM,�q͕kCM�[2Zx2����^�w�#k`�	��/�?5|������z��������)�_��S�{��C��2�ݢ�[�\��E��|d�fvU�v����z$@<�VJ�55�?q�ٽ�U|��`���YX�L��
��4���E_a�6{2�@�o�}�Ӥ����]J㜩�ީ�6�
g�Ľw�S�����
b���>a�w��p:���W�խL�"Z�{X��<���흝!Y���U�)�7!�ٳi���D����
k����=Z�yl���~���&��2�y�-�e�ը����������<��5�ǲY�V#��8��)�*Lsy�V���V����h0(�q�f�$�Q6�gW�pЯ�\�KE�c��[��gj�x=�]կ��^�ӡ`q���Z����m�C[���[�WBѩ���6\ow�݇�a���(<�#�	�{�x/!��� *��|�.������"�J��k���>�%0�2c�)����5�c�z��z��4�u�lH�=$G/{n�5���)!ᅻ������S��}���,��Fi��R�T���ӆP�g
/���Y����HP#�ׄ�����o��\^<�P�����X	P�M�1ْWm)� �W�g;��������2.]oG�t�#р�Cf�k7�;�J@<�O"�T;�u��}[O�X�.n���"��Qa�D����Ƕ-� ��|/�=˿�/GX�ɛ2��.�^�_�M�YQ�e������R9�o<��zi��@~��l|�O�}>y���`>���pda��muz���x�ܾ�)d�y���Т�5?~�y�JQ�F҅H൳����hj- 6�!0%��g����I�,�����7�[��Q�d[�pr�����3��(��Ǚ��>��`ϙ�.�K(>�vmt�Z�Y�J�$a�9�Yk�����3s�vG
���3	��u�հ�����Dz1���uB%/E��˃ ܟ|����ٿ3u>��̣�elʙ?v^���������V����<O)e�}W3w�B8������[m�t�'/��o_e�E��3.�d��D A$��������ډ���&%ս��s��@��e�5��g��k�RL�]�gt�k?q�S�w��I's����}�������E��y��z{����|q�KX!k���.��Uבּ���~��[|��ms��͎��R�J��N��j'^P,�b��a�A�^��[A���T<��(\sLL�Y|��Į����&vw�I��%��r�~F7�3.dE��I�6�xv�ִ��6�h]�w�5Ǜ<�B��:#�\�v$E�$z��,�T5�'�;�yj�t$�9�1n*��
2��Y�mu��l��y�sc�r��F?q��/߆Шj�JD�}de��	{�<���׮A~�[��Mc9�jd7q�������e¨��K���3� `W��	���i�_?+:r#�Mc�X
�_��f-�����`�϶�����+�Ey�$P��A^��|=_���C/��xX������r�N`Vza��H�T&Ʒ�O��'l���=b�UZ��t�$�YF���Rqv�Yێ���ޘ|�2~?|�=��|���7�ۚ}����@�
c���>�sǁd��)�ƃs�>;ݼ0���kN�R�x�ʛ9h�8�8�C0`#��S+��tZ�uI/|b�C�ු����<�����{���P�����Vqj��Ie�54>��^{-�6�i]z9�w.х��4R��cfm�t�T�X�R�չM���c�����ք�Sum�ֆ�R���g3i�q���r5�M��&պ���U+]�u����Y�h�Ҧ���,�ѭ��n#L�]��E+�+�>V�(Jk�I܂�wz��nI�X�XG[Q�J"�Շ7���}p���wV
��T׳7�[uZG0ASE׬m�݄�7ǡ�8����w\g�r�L�w�Fk��q��c�Ϗu]>�Z�t�8D�F�ȗ�jr0_�ۓ.'�*N0S͝�Jڍ�k�;���<�.�C���_�Rk �{.���%Ya]��Q�S!���&*�faSmU:*u� \-S��NJ��l��t�:uT�0WlGz��W��㲪��:��y(�2Ve���f��v���"�V�"�5ǫ��@]VT�r�KZ��6�����O������&�Y�j0o�|��"/(�F�5��k�w���ń!�.���6��v���kW#�]�L�y*�EG��[�nS-X�K�][�Ց_V�F��?LwU�}^�Vs���O3h9�W+���l�%���4a}r��}���wF<(�%nؽb����խ��])��s�|̈́̓��n����vZ�tL��Y}��&I�zi=�}S���J�U��g���ʲ+�f`V�B:���J��!joUaX��7�<�%�cEBN��`�([b�˅[���Z�];��!�F�:�6̧y�-k�����+�&Sx��"��REٵ��/��^�i��xZǑ���"�7zz�Z�{�X��:�u�]k�L�o�^�.-�|���{1Nv���W�&1�|��3ϧ[Ő��*����E,��K(�,1s��Ŗ�^�A�Ő`�O$��]�7����͵[��o��Հ�!��=]/_)U���Օ��ɟ����̾�`�$"�/�W�h���շo�!�E��6ÙW}��:9��3��]gN�5�%N���G�I������ߪ�T05�����]u����6��k�>��4�'h�jm�˨,N쓠��JgF�X��1k��k�;|��4zm�jU/��ΫQp�wK������� ���ݾ��m��v3m!�%f,72�Wh%�H����V��I��$�>$�O޼ju�M����r��h��F��CS#�M6^Y�ۃ&����F]c�^�2��4���&��,S�w������*�v��ru�HECY�Y��)c�>{l���\n���k7�m�΁�N��m��*.�6�.ӽ����(���+{'Q��^�:jU6Gͺ�vq�lm�}�"*�;=Ֆ�$��GfY"7�]fKB��̴��ݺ�þP8�l���I{������~��׊�MRZ}'\�o�]-w���Mx���$BI8�������믏�k^ֵ���k���ON��		<@�I$֍�]�XB�x�h��	 {��><<��>��ֵ�kZ��ֵ��ק�! ���lQ���K�L�*����w�U͈�[�׷���^�ֵ�k��Z�_Z����� l^b�2I�n.n���;Bt!$:�A�=���y;��\ۚ�1k뺼Qnh��j����ͣW+��b�U���瞘~u�_�/ܫ���F)-znF.��ңfoOZk�W����5�[�\�+�\�\ܢ*5��:�v��n��.x�7���A�-�\��1���Z��71o�1L���睶����Q���F���O}���7����zouA��	 ���ǂ�2B�T�����:�_��i�e���8��暚�u��O<ͭ����sb���SLxH�]��9����A��p�LpqD�����J�7�����/���N��̉��L'}�'�Z�r�'��:��	֦z�Q�ޖ��mW���E0�����3�Ј��	�I�ݑ��h%QaAgO2�ډU�x~���s+%{�z�T8ljiW؃���M��� �	����SfE&���b�j�Ԫ��Os=L��;�Ъ�oA����+�c�/K��@�¯���00���D�g��.��w�}���%-y>:�v��&�g~DQ�탾�J�`�lqq;�������Hf~�L[o��q��u��<�}����������Qa]�%��^��$�o1(B���}U-�o7������[��G� Cg9�ލasq�j��f�w��CvB.S�Q3t=5�B|d�r�d�����r��(�3�{<	�iāK�~O�N&\Pԕ�T\����xP�UU�_E
�sVCG�筝=R+9y����Cc���S��	��/�AU9�dA�@���E�S�e���*_�i�6�7Ci):��6m���9ז|B�����}=	����mq�;w�U`�u�Ք�E���D��e'�N�M$�p����ȸ���8�j8reoc�`�T���Åqy��R��	�"��]z
�<t�f4]�ʷ%el����滦e���>�:
�[5n7:��޻Ϟu�Ӭ���;Ϟ����	��E�_�<���Ϋ�%�O��xIl� �o�����o�h���S�;B-�8���9�T�v���������1��D��oD�V��	�"�"��T+��J���������]Y����bx��ii����"W=�}�T�����a�E�sıN���&��k�,8�_ ��m�36�-��QN�2ȈL1�C)=![���L�{aa��0��)������̬��!�[�\h|�ar��c���w�-�a7Nd�5�r����z6)��Q����v3X��Y	�J/��w~n�q-z�� �s!|p���?�ꏈә�e@��U�UK���g�:�R�j5�633ZV'�k�m/O^�܀��_��;�;�^�\�+S��3a�=����%���y��ډ4XwG��~*
�FSແ ��Z��U[�B������0��mW��i���:폍0��o>���$N�僱�Z}��ӏ\��OT����7O�9G{�`�(^�#�����<X�ǟrwH��?-�`��|����vPޯ?�\�^w��B���XN��U	�.����#�'&C�YD٬��]�}�u���{0N����t��T}p���m�H�Pي����6��a�b�k,�J:/��mJhq��T��^���xN[Cigr�@�S	[�eK��W6;lv�������E�l��H�&�&��&ppGw���p��U���88��AD7���)�>s�^�q���4�Qɜ>���T?�~M'����_� �����J�Hl�vU�v�n�+�IZĶ�%X��,w����Ȏ�z�7M~�p��a�������~��EU��c'�hW^�TtNEgD�%��R=ЬU�w�KL�1
v�~�w�)�z�9�����ct!�ܽ����ǨP���+�S�j7!�6n��ڙ�t�w�-�ʆ�8��";�.��3�	�� ''Տl��קy	Mg��L�"S�Fu��Nk�Ǭx.��<��,�x���-��S������׏��/�Cu�ko1�%)��
�

�d�Pg��4}���]��,+���8?3���!t��a"r�s��u	�v���Zepu�(v����8��C�5��\����<<b�Y�������ݑ��܄��#���e<Z��[�(C3;�q,4Ҍt� M�t	Z��1���xضQ�r!6��3ܧ�ygE���l�oH�#�u9�d2�!�1�OȲ�̷�茂�!�:ᅊ��l+�>5x-\���{����(v�`x{mͪ:�K�qm���k��>�{���C�B{}�Z��|�y������sźt��ם��./������ð�1�j�}bhE�d�L�($�"�fĩ���%㧂M9��jE{U�8ﻞg=s��6I���8)�"� <q�f�A,Dk�����z��cCpЪ�����M�U�Q�����|kg`ɕ��H��ղ}���˨~n-��ȍuS[d�>�ٞ&V8����ի�<�U܍���V��R�*�����q���74���Eݘ���%���	X:'���G�x�̋�;��xRu�7U�|?��ɯ����k��)"�_��9��yZ���.Fd�㲺�G1B�_��L�~mz�1n9i,D8ѯ���#��BqA���0$�[vY�Եc7�Nѽ݋<�N�nSy���)w�5����H��E>O�)}׬4���
1�ѵ7�|�����n�Ϸ
`�"jR��
�q}!�r��=u������S��C�65'C�m���fS�ƛ�R��Ǚ�8��/��8;!�u�Y��1���Z$�����Ŋ�A��!�}�=L��Jca�����TGtB��~��N��a�wj�� ��h]	��\�,#�����\<�u���͇�K�Ӽ�����b�$�K�h���Hy)W+�Y��XN-�#3�����Q��мͦ�S=}��Y������ɧ��k軩>�N������#��t3��A+��,�D1�	h#�[/wΪ�V�0P\�;�}}X
���w}݇���I�]�JuGB��!��˻κ4�L��9s��<�w�|(k�8�88���0���L��6ٟ3o�U�v�}���5G
�g�q�ʘ��|��8~�Gu��ɚNz۷�KS'0���=��.��%U�
%(L��3(Ͱ:�Ѹ:q������q�J~��ow��l6%�ˍ��'���*<,&���W=���\��Ȝ���2�{������w�:9^��O���9�1��jَNG�F�s�ܸ�����L&�ͭ�o`��X��wp�W0�!��4ph��Ǟ����l�y��ö�
9�,n�ҋ��nY���ú���N�v[ø����z��Amw	��='�Nꄙ��;jK�%IaQ'��Ҿ�/E��������\�_���"�,<`���+��,�/	�Ʀ��Z�]���nj�f�x��2�j�:�PK�Z��vz�[=�@9��?�Ok�ϒ���ے�v�nv\y3T��a�>8U�=5�K���C�|@->/A��j�`<�M���ڟ��u�A<`��w�#�T�ry�f�7��WtJz&��/�m<"ؗώ���7���������jDs�\�Ƚ����{uѤ��i���7�'�{���=A{Ҹ>��e!rX�[��d`WYɔs2�ڗ�L�ռѼ��Hh��7�������˯t��^gQ�1^��s���Y�9{}��\���/yy!��x{�[V��+yK���R'�y�����@��i��ڲ��r��C��ުit��bfY]-�ל����Z��8s������NyPصeݿڙ�z�Ig芸'-���I���)�[����%�������v�ql\s����ǬG0�C�^�%�\GH��k�M�N<�k���4м�5���!��]
��5��T7���.�k�E��R���b��?9��<i��V��=Z3�pIk��zBeK
OaQڟ5x�e=[ռ4��;B}8��nrj� �+6zw�ڄ@������{l|By�z%:����2kT����x��l���j�{��=-�;��;�Àe�|���*��8P��F���s��,S����rYI�u�d��pψ��$vu)�	��*K��^h�.@�L1�|��
���]0��J.�8�y�Z0�W*�����wh*9jw��Uy�n���6ف���s�B�0 b�׃�������T�OE�a�S�'ˤ��R	n�~/B�i��遧�|Ώ̢*\�?cf�Vux�{���M�ҡ�F�xݲ����-b�Aԩe]俒��q�e�)�{��`��m�9�oo���T�D��>,���V�U�"�Homٱ��ӗ����9��&	p�Yʍ�VlqF����y�@�Z:��BLFb������L|�֜r2�i˅���$�6\eƏ�����������yx�8��ͤ�7�~�wgm�*aM����{O�a)�mƷ4����F���y�O�Ջ"���U<��}|M���ʘ�,dF�s
�R��r^�ΌlO��~�c����9׊ٔ>����>���	n0�?~��P��5K��L�T������&G�p�������S��a��ȝ�[u[]˔v�:3�7��|ԭ�9�TG����@N1�>ռW����[����_h�X9���fiʥ����&����s�A���>���~��׀@m�ʲ��,a�O�L�jYʹ֑R�nk���ފw��D�z$!"�{`�$��O$��;���hs�:�b�Ӧ�i�a��H"�OE��>ŗ��Zg*�>0�~=��vR�e~R�+�l�1�Zzs���OM�iu'͸bC*�SlnC�l�|jg]�v���ctzZ/�_�<�yYk8��$�bg�(R�{E�*��0�$Jl���d�<�%=��
��p.�7Z#�ژ���]Z�x�na��=�␱�� w<���	��>|�‽�b^�3L�_!�ɽ�w�OT�x
��+3%����졑J�?bt���uW�Ė�h匩�U�r�
4es�lk�y�,�C�u����噖�S�����G����Z^�ݵ�nѩ:�'�Ϙ���x>�Z�#�WX��$y�����/!��<��e�����Bs}�N��W�ퟞ���H0#��L��µ��F�˨LK���h�Ysywש�wGg��	�M�	�Ϯ	��m}^��?!f�}�G�O��7���<��!���R�)j��U���P���y�k|;+���^��y�b�j`�=a�Bn�G�����N���!�T�&�_�)/"��~e/��Z~X���j\^GW��c�np����p��v���/7Yp8`���a�}�<6sО�m�n+�\��$&R���X� �;�Q��xc���rr�6�s��e�������_��x���V��Y��qI=�ێ/R�ٴ\�mD5�TF�֢Pd�[b�6C�%~	$3�p�p}aH>���:ǡ.��"̊U��C�5��w6�4;N����{&�\J�ό�RǐH�� � ���8֙�:?��%���5�y`����w����*�74B����Ť��z�z�W�Agm�����}���N�V�{�����G.�)�v3���@8�Z�c�'�~�D�+���ܤ�B�hRO�B�<���S��1�2ӱ����+��[����+sVn$;[If�F֫l��;��ҨFI�Ah(�jcv�̶��֟�%ϋ�˺��x��/]�[cm���sڤT�N���b��x2�(��m�{]S��{�y/!��<��5kgGC��j5s���z�<�t�En�/@�4���iXF�'��8�y�\�<�f���_�fHd	����{�m@=����Ŵz���pb�T �t�X�c:���s`�wyS����5�+�X<������f&C�C�����c�cU�h.�!�M��)�Jy�ܷ����օ����G��x� i�'�Mm�Oe36�lu7����tf�$@��݃+x�T�XhRS%�����k댇�{g�#[˽F7�][��R�Kd������[a�Ѓ��`���4 �Wi8ܒm�?f��{hG�Ӎ�m��>��J�,N�<j�m��>���`�}v�<�"�t�OIq�O/��~�Z����,�|_�h%�no��.�
�h2�5��9�ʌ����q�d]p[����ӏ��Z�^�Lf���r�;���;�@���1y���@�"z��I�W��;���,j�'�X�T�����^�k�ϙ��uI�����޽~}���L� &�z��������xh�b�o�����x�)�է.�L����`���Sz�Ufv��D�YX}�[Ho��-ZT�z���*��͓�Z���hd;j@/t&8?4h!B�� ń.���Z͎o���oe�k/\����q�n�n���.T'9.�'��k&�Ʀ=#\�u����{`��w�o0�y��G�2���*a�ޏL\��zE���ia��鿎��z�uz`c)�3m2��'�Y�6�&��d�WJ�oXJI�E���9��'�y��ۤt�<��lsZZִ��{#3�b[�}V��3���K��-~�h����w9P�u�=Wo`��Ʒ��@���ŵ�3���әKkA��)�&9pd#XG�#-�;2/���|�RXh	p'ła���q�EzY�n��^�`^*4P�����9�<-ꁁ���=����**����v.���2A�����I�7<�e"����v9����o�T�`ex~B�<�R�ߓ�L�5.< �r��vq�[i��D� ��ީ�6
G��##)�t=C�זx/��$�8���n�{.0K�#�����d��=O8w�d{d[_>�]�C�2u��͛a>���5�L��h���y8M��md�����E�v~c�O�w���,�&K:��~�j����OS����
:�M�xa���.�pIĶ;�&<Co�F4�<��JuiI`���B�b����Yߖ	��{���ώ�gn=�66���an5�1���}&�|���h��g=�%�m�R�7v��m�؉���U����E�f�|)]��l��^
��',Ul��>vOu>��`j��W�6HD9Їr��0��
��`H���:�-��_f�H�3�R@��7GS�����r��;u�������t���[7��L�['$�3��L���0q�W���kM}WJsz�=�v�Z\29��g7#��Զ�uQ㓱�W]Dz�����j���q=>[b�(�=햮Ny��\r�C���'��:��T��F��Ѻe=WX��e;W��P=�L�	U����>M���w]RVa��(¥%v�t���3*ʎ8��M��B
�yV��o��u{�GzhK�F���۴w�]כ�m�/��ҝ�A���`h�8V2���1�'�Q�{.;�J�v�C�.�汢�U�ʏ��Ds�1�Ee�x�q[,��s�C���c���w���v��UC�уi�	؁�*�7���.�K�ݹ*̹�?��ө�}C��^��iUZ���J�u��ے	pˍ��2�wvuk�2=r��˛]��ۢ��m�
�����(d�yr��¦������o��\u������zTm�Xo�]͠����8P�:uʮF=,���&IY�R�0��;,کZ�MU�:�m�d94'B�lZ���7%���%5�k^���Ze`m���I�H���LK6Yv,X|�^L�\m���d}�y�˫]����ad/z�$�[%\�PZ��ԆV<P�jr1:]��u9���d��ЃgwCK�:�.�k�����o%έX���7y�mI)��i2�)���lU�˝�o/�.����>���,����]����N�2Vs��������WY�=�Yy��}1V$,n��Ff��A����hq��N�3����Q����\�������V�F_CR����o���ꛊ���fM���B_m��h@��=����yS�_\ꌝ#p�t���3OWs�H�쌜�z2��Sg^�A0v�ru��s%�=7<�*;Dɜ�+��3|V�ƫB�nuZ혞�:R&��:�b;��Ky��u>��i	)�Z��ݬCq��&2[
�8�d�.�A]͞O�q��S=�s�j�7w��͈��$��=��%J�n����z��yKoo�}�u͡�+C�]cA��N�*5�SDu�6���-�7�4Z���*�v=�{�jRl��[�w�N����dOL`��Vޡ��1]����$oi+ +%c�f�>E��i�R}��g(��JԸ�n̨g)�(igud�g�B;V�{��^��r��!+���xܪ�/l�9�0�_cT:aVH�s�x-;.Ոܗ�d���F�����l���9yj��A���K�Zd��R9����AL�i�P��{�-�s�I:�V�5���UP#%�r���jU$�D�j�H�T�^ay��9!��PT�FPi�l�%B�5<��@�&�K�&Ԇ#蓅60�m4QmBA6�m�H�*��6Q	�˥�x�	&f/�:�r2%��6I�S"�O�Ǧ���ֵ�-k_���ֽ=8���$��'S$��C B,��L�dd�{}|{|q��k^Z־>>��>����Ȓ[�ܓ�������"�b? �}����2r���������Zֵ�||}k\}|zzsئM&G$��G"��3� >�22$.z$]j(�W�n�[�W+�\�����k��ŴcQ��+ѭ��_���_�x��5͋r�*ō��oo������-�kƫ��V"��]�h��ir6�7��_mr�Ź|Ur��n��7�O!�8�"�"'Q#�T㩷��(�R2�P&�r	F�,e-b�+�Ur,���7Ƿn�u6��[4-U5�czg����ĖU����IT�����w���ނu!����jB�*I�¡a��(�����<|G���F�s��ϗœ�ړ ���_��8��o��~ܹ	�:���(�_�<K�4S,��*E""�fS���-~e���qA��O\����-'��g䄅 _
�;�A��y����r�����dqޠ����;܉r��72;�r����f�A?�����M�}7���츑�s}}M�9j��b�2�9'��֔'��Z�<�lv�� |z�_1�zr�Z��v�X���&�r`����Ү��EQ��Q�b���>��^��#f��y��q�
�N��O5��|���Naᷢ6���+�<�k�PKܼ�jde_�q���<�w�V�3w ���<,=�vd��D����,�5P�n�O�L�q��c�j�;0�K,�	U#:P^����;���E�[�2|�\k˄_w��4�P|����o���+�~;�� �
��__ڞ#4(����W�5D���m��.e񒬐�V�I��t�ٵx����v��_�����b�%|v����H���
j�A���,���,�eP�V;�Qщ�����V��t4�^�je%�	x*m�C�D�����[�J�F��~�w��T��e,S[�6���Ȭs81���J]�7Cw��i�[��c��v�p�&5\2a����Ü{_j%�lN�[��\�S51�?��;�ǟ����ZRCܺ޻�g�.�hE{vS	�����qz��Ayǆֆ{Z	X�s��4fc�ΣC�O�x��W�4�y���ۉH�}2*)�̛���A�·Q�?�#����Wj����چ;��ٮ�����`j�.}��MDt ɊȔ�Q�a5� �������ᱰ;�qA��4��<�fA�KȀ�����m�h�Dp��ĽUP+j�_.V5�sn��E�9"W�u�5P�+���*mA�0~U�	KH�(h����Y�:���ǲ�lR�T�n�D��*E2)L�;�z:�O�"��ty� ���	Hv���ͼ4���駲�z���w�&Y������⮤�<� LP�����%�C���tcC#�9���M2D�=�1@Lpc"ᇚϫ��F�s)~/I�^���T��zi�������`b(aS��̵��s�6p���OD���T�j�vJ�9!2�)���c8B���OZ�p��j*vwZ� ��/�;>����C�* F�d��ٍ��,���T��U �f�
3=�ٶ���xAO;Y�jV�[ّ�}3-���'�c/�`�Cu����Iu�-v"p!�se��E@�f���;ҩ��9ҫ��3��y��a��VtJ�R�3ծ>2QX��8����Kv]�lR̜^3���P��7���8��ǜxa��݊r����� ��i1x �8-��}�`���m�е~�a�:Q<i���l�������q�1�B�H�N=��ll0g���!74C�"�C2|�-4�L���N��uC�N�6��
�"���8�����T�SWk����+`�ɚ}uǝq�A��-вCc����5��)=x�;�a�<ݡ�=�l�#`�T��n���l�&�b��~ŚA����,~vg�|��ע��~?^?/���ׂ_�Tyv-�I�础��}�k������JCo���=����'}Y�V��N֜ӌ���P�g������pYR�Ӛj���t,��5�"�<'��x�`Xd�ک���<�`ecG��5�uͽ��\୤9g,��@�ڞ��%���-�t�Å�T:���0.lD��x琞�32Th�/�������oa�A�pco����cȒfy��;s��ߣ�XY[W�JO�o����?"�Rљض2���5pͮ�x��B���5�;s�u�	D$�6m�$nE�*�^�o�/�w�}Vܪ�h�K�l �۫�#�{B�y̝n�vߠƉ�W�7Ց���F0Og*9�L��yj.�G:�w�	\���!a\��I���wU��:q���jS�E�u�j_K�<��0��m^�PLE�ovmSf����x���88c���
H.�ײvy�X4�K��v���Q��� h���M���%~n�I�I�
~������Ur�1ݲoٻS���!�;��E�3�|u!�\�vSѯ��ٞ=�d]ct�Տ�~��"�X����7�;}d��!��(���׎r$D���/ؠ�~���S�(�dNQ�L*�J�K�6�X���"@q3cS�\]	�J����q���^m��a	��n������[Y���*���K�UK�C��t�*�u�<a����@��p�-"��Ƕ����>�!V����\�4�r+(^�;>�./ƺV��-�y<�Oz-�\}s�^��g��!Ļ�e��w�몙�Wϫ�e����ݔ.��ڻ=c��fk^Ɂ9�[�� ��X���n�*9a���{[��3!32�40E�gsnna�s����w�$v*�����0\�
چ�]U!�eY�~��e���S>:�ix~A��#�ߒ6��3���GIL��� �L�E����=��7���w�_{`vf�I��1��l~b@>�!��З�zj���=ʗ��B�s�F�ʹ+��5/�)��~2�����:u}✿�X��>ݒ6�%��ؼ���+�n�=|e)��v���'��Hc��X2Ŗ�@�ڪe�DU�����+O���V�SHN��Rl�X��WJΜ��*�K�����W#��1�m9W��eu��K��H(D(B/ӌ��p�g�pH�q>^_��Lpp{�V���I��n�x�'���(M(Ԃ�{��o��t���זx#��8z�����bi�Y��4f����%�z2���Go:�빇V0�zc��B4;�k��f����zg�r�P�5�������&�&B�>g���[B���}B���"Wm����*�
�1�)�,�,D	Rg�4
@Ex�^�O5Ȓ�Ғ�5)*��<�O**�jv�y�ˈ��Ji驜�ZiW�2���G��Ǎ44P��������0�ъY������Y3�����jJ��-cٓ��?��W��`���@0-��|�����
n	x�}�G!2ƶ͓��'7�N���U)���z���۠� 㖧z�>���G�Q��l9d��Z��V�Ƥ���E�׾��B����e���zb��XJ���PN%��솏7�<�cI�~ٓlN	xpe��,0l�	�C�?C�������%Tx�е k��|��~U�KӼ{r���k�E�3�Gmm��,\��y�G�6����l5�,�vy���Jױ�	{���<L�5Xb����oʦ�S��fX��s���W�#���u#�5f�m�ޙ��`�՞)�
��T�0�;e�j�QL��V�Ci���Ɗ�[�13�h���+���ü��6�K4j���a}o�g;4��m��ۗ�۞����伇��3F�Y�f��������ѯEz#��Dթ��G�y��6�'�,�g�=5�5�y��r]���V�z���'�M���p͡8t'vƾu.���3]��E����dO�5j�"����}[_���?��U�$��\��$�Z�+$!,4�{��J���� tu(�v����=a��!��O^� &]�6	P�魬s|�����?vy1��߄��pl؈��'Oy^��t%�޲�|���o@����/C33E��X�xi��eռ���0ǚ�॥��^�ؘ�'�S�@ĕw��Dژ6�X��Fubw����l�����fe;%l���BQ@�F~����!���u�ތ�L���p=��(����ɪ�JsYc[��&b4dd��d=�]��������������'ލ {���a�?6��fsr��\���֔2�[��7c�I��9U2%>��w=��<��P?0�O���{��^���W|��s2�I�v��n|n܄�\MYJ|)���:����;"��{�� ���	M���C�����[b�z/��MN|"�Z�`[&��7+��/,�[7{�Kei��0ɪ�i�\��L]e`���n�X���|Q��f�����M-Wϳlv+���ʺ�r�uB�{�[�Ѽn�[U���O���G���d�U�����<���-c�AP�Xl/l3�\wI����b���)RTXsP��a�轌a���c��ۤ�,h�+ �����&�*cp��}��^�ŧ偔�i�S�zi�lZ������ӓu՜�p� ���5�+�=>�4�تq�R�ߠ���i����)}O��#F�b�s���eZ�J�}�*yw�r����7P`企���!�=;�-��Z���^�y\�������j��5�s��y�[� c�g���9���z_['�=fE+9�c"��>�=�X9���]>Y�e,�tg-��;5��h �_Q����qJW������x����gd�ۺi� ��i~bŤ;��S=<�؄�g�o,ߴw���Ǹ��U�k~��P�/\aش�a�r!�z��X��	]�{/�Y��?'����W�1�o�~H�ϕ?+��v~t�ٚBC��mxZ�a�v�B�xj���]�o�i禿M��C����`I������%�m�QM����Ů�ɞ�~���J�u���d��u6��WC(�ڙ�}d�:�7�$ħd$g*]j��l�RA�OvՈ3��sN��Ǎl�.����G��g9��əكi�ʆ�:*om,B�7��i���;��+���t?�}���>#��Z��efT�+�l����utg/>��\ ����=�{�V�1�<,	�Ul1�.��9�[PG=P%����r�N0Y��y����(6"K��
3�$�C��Q�p̧Ix�	O�e.��cS/'��0���k�%a�J�QaLt
�l�T\<����r���y�0�i����GzP�1��-��lf�M���@N�'�!L���GM�y��1�Vb�۷oxeG4��E�cy 孳�_��e"�[�M��R���J�t�N��n�����yU�"OεR����	����u����=���
y�1��潘���)�t�=�n�����E���8�2{1X���Ʉ��K7��5�p?��X��&�l��º�(:�������}�ܦ�Y{z���Ac�K��]�k���q�`5���!7��u=��J�"G������f��վ��9*��<ʭ[�<aӜ�U��P5�퐡���ɜ�r��wvX҄����Wy\6��Z�䠗��Q��i�O��[+�U��y0����v��~�ب���x9���������X�;�nU�c��S�LΜ<�d���J�N�P��*�>�HT.6��%a
�����WÅY�V��A���/#�mٵ��o�#��5�י��|I�^�i�I��om%�j�y��1!h�U�����S�v�Y��2�$
�(����t$ls8l�vf��eG0M;�P�z'A0'8���zm��{���4��r�V|:OX���Ƈ�7���|����TXP�/^&��Dsܼ�f�k%,�*�Ub)�qL���܄��|/0��<�z�Ύ��`�qL��O��M�\�!S|A3+����2�t�b��0%���z?Kս5Tu�}7Fl��ή8���Ɨ��^�m�r��_��w�����P���~��ς����+�4���NnmԾmi����|�@�@.2-��^����c���Ah͸E˧K�h]
������{s�'�yb5����I�Wk
�tȗN�HL�a��Z�F��(�^>�Y�p�$uE����v�D�73���Aq-s�>!��cK��[�)�PX&���w�k�aj����ҁK����������+��j%_XC���Ƒ��Lծ8X����$��Äл��E٭���}�e�����@�>��͐cK�~ܩ�������a���k��]�gWz�gVELC���{�,��}Ѡ��1�	:�lj�؍�6,\s8�M[�9�������M��c���C!:!��i�';/��������{���ǎ��;Ӭ�FRx�F��^�o���:e���ݩӕIҶ���A+d���}��>?��L�b�4^�ο0�R��nq˼���9j��ޚQ�� M�6C��ݐ�{���V&��8��L�����3��8ŧ�%�.�̘CX��`�<�b���.M��0!����D[L<?�:�9����d�2�j5�PJ�rc� ��8���W�Sٞ3Ҫ����;=��X���^���j��S��1-��`�R��%�^ÊR0>��|f���Icz�ql:v~���Y`�����L;7[Ȣ}6���qg�{{��1Y�v������ks����}ު���%5x����k����'�~S�i�ʽ�d�]�7+'��?2ޘ�4��*X+��C���I��:�z��C��PI�cù�+��bT�~N��7ן����v���ʶӻ'$8$ñ��׵*j�c�|G?v��n�����r�ʙC�bz��zV2|�]ҧ�E{vS	�R�oC�e���xl։Z�<�;�9�7�����ڧ�3Zμ�sKN�@=�����	/B��q)�C.QL"�Pw��m������Z�&�F>Dk]�����`�T�$j���F`W�������W��9ɕn}Sh����AX�V�5[�j����p��W�1(v�oX��d�Ɂg(����S��KO6��i�!v�v�u����Z"�
�Fc�S2��>��T���h,y-����Y�nH�嶵�3z�dY�L�Vm߲[�@��l��)9�[�8�26Y�S�59�*sy5��=8"�x̽�-v�8��Q�x��RE�Ƿ6V9wmoI�،�Ӕd�\��S0օO(�}J��;.Uӥ;�U�uKd9��q�>-0u�F��>yDjT-��ڷF�e+��ɨu�`���t�Tfн*q�b��0u��å�������T]�tg6�No�s�U����T-]:ew�s~zA�K�V�2.�y��ǒҸ��7�t�s�O���fB+Q�Œ3�����C����I�)�8�5mN�*]G�K;V�S)��㵮�ⓛ�u�����9�p���j��	�b]��6�Q�q�r�ynX^����6i�ʦS��B<���XB�L��.C4�][�oJ劃P�%�A��YD�2��%���/v�mҡ��B��ڻۨ��Q�Ƣ��Ok1�ɃI��W�"�.�9<�;k���4"n�-����.�n6H�y��ت��m�����8���a�a�m��<�:Pą�*�yqV���/N��M�CHIYG5M$P�y!��k,~Y/�o�t#��[��]K�v�6o;�]�}Xʦ_q0�j��G�o�Iٝڦn�͋"����qE,�d��$��6�X��:��*��N:��=�&wO�mڌ�6�6<����Q�.��C�[�fm�Ȑ�r��Ysv��+eT=����̯��w���Q�}OS�lw5��F�i#Mb��l�n��Bp��neV�=�QC._,Dɩ�0��"�<R'6��sz�:T(6]8�L�\r֋�/s^���ҡ�jVCd���2���õc+=r} ��t��̶�D���,[����R��ٶ��l����ub�nB����a�*i��W�q&L�]xF�};Sޥ�$Vޭ� �X&a���v�,��Q�)�˷�Չ�xa���L��=,Z�WR�M�]'H�nsy;�L�o��x��Skkϩ�X�-k�-�zݝ���IHr[�\��i�YLlv=���;8^�	Jw����;F�k�fj@f�g����r�x�s��Xt�.ݕ	\�X؏*�6;�!vwuVN*��e�q�ԏr��o.���ۜ/�dWr����O
hg`�}�[	�u˅\���M̢��Vo5�8��E�I%ӟ33><JG�d"�dM ȒH!�;���@O]x{yk�mkZֽ5����k���ON��.D���FDd@��������o�kZצ������}|zzpN� vw�$��L��|}}zkX��ֵ�zk_Z��ǧ�	��\��c\�ҹ������W9�{_M�yYoC���u~���Kr�M�k��E��~����ҕ��W��#x�o��sh�V-�.r���p�F��z^(���}�u�W��鯵x���o��M~6�y�\��*5_M������J7�w[��D2�r�66D8�Dȭ{ΟQ�m�����������t*�t��k�8�Sas5u�)��K�Jel�jj���%�l��Ex}��������\���B��<��x?�ȷ{-�Ô��Ql	��>�'vb)6e��ɻ)�X~��c��/��ӵ�,ȼ{j�3�|�fA8�����XQ� �ƯEr!��K];��9Q')P�^��Ji����䉵�
����&��&�w��U]u2������ o<��b]���F�+���I��:�����W�x�Z�MU�˟.ޱ=��z����7��B�d�Q��o?��R���LP��*,9�{.�����*kjYK�_v����p�G��A�;��T�m�p!='���9�{�q:�c#�B�yp'1���Ej��F��֭������ΰ�p~h�g�
��\�7�^�4*�%s���_��MN�.��O5�{o�µg��?��Ɵ��ƴ�DX�X�B���BdN���-��<պ���w�P���E�}=���-�(�J�a���4��3!��m���Fz�E�_�f6䮔�0a��7���C�lI`h�c�dﺽv�N0˩Ou��k ����?��U~��G쟥su�Ym��V��:V�L���So�7����跴2$&��O��r���>����뽑�av�N���d��'(nS7ҎmeI)]�p����\ܘ�f�;��ɣǤ�JHj�\�ֺ�+���x��@�v�qV1st�ޗb�"Ԍ���>����#�����=�}��ύ�T(j���GDn�&l+�ge�6y�6�Ю�&+`6?]o7���0��,K�;D_��kk^Ƣ��*�1�\���-C�Q�2�cV4bS�.�88��.O�Ԕ�M���.�En�/@��u;S2
5�E���n�w{�?K���>�l�|��+aN�zd_f��F)��$�MةL�y��S,��:s��\nt5�ߙ�6i�t+�*�7,~a�z*�g�!�۽U/`���ڬ��]{�[�S!7�/�G�3�,��s¼�������mW�<�X"��ȝ�Q-3
��4�n�/���}h}���v�cK
V��
c��+�\�<��=��L3�=:W�EZx+o%#*cK�Bli�|���a�%:�I¿��N.�6�+��FGS�T�GYn�_e���=>��+�)����)��e�	��Ҵ�=� �C�JsAU��m��Ȫ�f�ׯ������I]�D��gŏ���Hp� �Ҁ��^��x�ߓ��l �~�e����X���t�*�փ�Q�Wǡ��ov>���>$h�1�{iR�^���4�~��"���S��"U!eu7
4)וw�����<��Z�b-v༏�7�`��˶���*뜷�3]�+_IEu��Zj�wve�>��$X�Cl��a�L��I�����q�b��"�zQ����Z�k�Xß��F����3�̐Z�%E���Ń�,��n�fD�4��6��󷮟w;����^�E<�˔�ZPX�R�5<;�0<�g1ݒ%��LaӅ�P��i���*���*FvBO~k���RΙ�W![�<a����@��O�I��/�v��[n��'ʆV0wfz�P'����Z���1U�A�j��(�#�{��:�;�`��g�
�� ?'�C�+��`�E�T8���%Ċz�C��Sm�v��q���I��9���3�?�ʼ]h��z^.��/�*��ײ�`�N���!���쇉Yz˛z����^0�C���Y_��Q�Z��8>��)�EE�7��'���
�w���1�5vr�u�Aׯr�Cb7Ϡ��i�Ou�� `L�\�NB�QyB�~�����{7�d�NSS��6Eܠ�����.�9��]��t��UHA�6�ֿ�����qϏ�Dl��Ο��|���>��N�1����[fJ�e����3|��K �p~�j	�ۄ\�p��N˯'D^^E��h��`�1d�ڠ_�8�WJ)��s3�ì�NPmM��&8:��&gCr��>s5=+�KU\̀�4Ҥ	�����T;��*p���-]�Wo���6���2QYT�nM�%�3���|��mA�u�^�7�o?�y��qu}Ӂ+)�j���M�F��q	��������SY�	�XhRu'$(�xq���C3�r���Ե�{Tӫz���@=���l�A��	������)��+�^�O5��M�k��J�ї�|;zo�Gw�x��fZ�j�<�׽���ز/{0T���A7��kܺ���u��@|�yU�|L�Y��)�$�� ����5���z�!W�0�����6ې�U�]m�5(�9�y�מ1I�F�X��c,κ���ܶ�p����'�d��2�����=��S�͙���g��q�]�f��zKb����W�+kG�Y}�<��"�Ԧ���E̰�s�W�-4c���栺�1�5��d��Q Z�c	H�~��ֲ�m�>���#����t.?�O��A~��#��������0�ܥ_��r����lb�9�IO����3k��M0U�3�.�}.��C�U�����W�n�Oˣ�ӭWX�WKj��4���ӯC�wy�r|$���G@f�\<�!����K�|֓7�<�	RV|F��K�����+���X�;�o\�	|٩W�j4�M�,���{zM8��8m`F&H>$�)z�t�M�c�.�y�kU:\WC3Z\�u3�j�\;p�XИK��ޑ8�R�.n���s�I�B��W������~c��|sť>>��|��p�g�ߧb�$��5=G�!׃z�����Q�C�4p���=^B���� ����g9��[u�O>��R����<;*�;O�`��H�I�k��O��DT>�Ȗ|��]^=S���ʆa?��p�(����-=��N'�p��z�z�PݒÔ�yy��r�w3�����1܅7�7$���g2�u,"Y��#��|
;���^����L�T/��\
�`�zk̵�%�Xhl���n�vf`��Q v��{y��+��ҡ�K�\zd(��Ϝj"S\�2�5ښ�w:g���$gz��[ռ�6;>(�P�����lv1��͑�W���[)ӊ���{LD�7�JJi��T)ǫ�v���<�ۼ	zD�xN.fb���z6E��\��WDȦz����׏o�%��)^f����57G\�Ǩu���׀���,�75p�(�큔����q=ԩ'��:���,������n�4�� O�K���߼�q~?`�<~�\n��v�[��,��9e^Q���|Y�R9��1�j��i`�|��.���\sV�Ur����v�� ��m�Є��N'���K�[���4*Q�<��F]�;2��Q��Ń.qEݩT��Rg-Wr�׋����W��f=�u���g.:��&��d�YtqM;��ۚ�;;����x���/!��qreJ�y�긖{���N�gT��4cHNCw�\�$Ķ��U�'�]Q,�Ź�RF�lf�kw�5��~��~�Lq�c�jy���/��Ll/�O5��͇���c�[j�otUW��Fj4�,$;33�~׆lVнJy8Y���S��Fji	���t��[��#�?�>��������
c�ʚP7"��㪘m�D�-_����O��ߒr^����D+�Q�f�E����?.�2���z�`fxnJN:���
�+�sI~c�z.�����M������5>�>{�:Ńv�vD�1־��R�r�J�~{x}��=�/lcn6��n*��}P#�q���㙼�=��Z>��Ϭ �/��'g�y��a�����G�3����̈�Zo�xr��ղ�Qx?12�c��Eצ�ӷ۴wi��M�Aɞ�\{�Ӎ/������Q��={6m�dgO>�x��;���r�gKݴ3�:{Wg�
��h�t��ty�k��3X����Op�3�P,س��Ω���{RT�.��y��Ԝq�(]�aG�9�V�Ҙ����T��G5%��l���8��֜t��SM�CF�s��h"9O��#�&��8w0�5�>�r�/����]��ܱ�G��;������qt�%��,(o/:}�����7������r ۞A�H����}�<|G���#n��}(����a��
�{c�Oj���XXX����Ɩ��a-�nq��:�����3[C�<�U/5��U�%[9M�q��k�����9ll�v�w���|�&Td�x*S)8�M�3��v}����Gfі�2�1�L����=VFÉ��!���n"�nɤ�<?��R��q�Kb���Fq(�:�z��0��z�o1R���E���0�]~͙+�$�ǘIg*b+8�b�t�d@t9�l[�#h��>����L��jA�3sA��	~nV�`����&�V���#%b�aU�'�X�BO�Ac@j�&v	��n;��w�M��b��J�۫]�xr�m:��<ޞ��5������&��Q�^ukr�����sK�	�^ga�i<3r��걩ݔ�6������|��*���ڑ�9��	�X����W�辽'+�q�}�K.�\���r�?6W�E~����z��+�9ٞag��+���^�C��Mc�&�ö*A�i�v�H�RMmV㛚C:��3�����'aV���<�ݚ�m�,#�_�[)y�s*)`�>��X[�SY{�u
ȓif�]+�Ŀl�L{{���V�ݻ�#�N��ܪ��wf00� �}9aq��:w����4�$�%mT���]K���k2��A�}����>p_./<�=�x����x����vV�`�)o*/���|��3Dz��@�r��yw�0 h|.�	텈��G�|��4�g;�g,L��=��F�����b-m#^)�dg ��Ue�a�|U�v�f`�Gc-�Γڶ�	z�2�Q8��>�^���S�,x?{��bV��|���������4I��~��4��c[�<�5����=�q
�<���׏��R4���5���l1�vC.��> �����7�!�x�3�v�B�ό�uL�|����@{w�"|o�@L��B��;Qӥ�Zr.�U;ٞBb��}��E�Q���?��%P��W�?ь�DsW�H�f�Vl�|�xVf�����;;8�p��P=<��)P��x�U�򂧝�<($l����'Q�����
�,�M�֛�K������/�ıO`.�eI(>�����߳*e�p��`\�&ӷPf�L�c.�Sܬ6/ 2GH�%��K��.r���-2;�`�f��,g\���R]������s�^O�&�9���(C {L�ۄ�u��s�-?2NX��L?5'���*y����]�[[X����kS��{��Yc>�셻7�5ݹnf��Es�����ރ/�v���U��Y:��◨��k��	���Z�p�ݾ���5�* �,��R�>r���g5H�h�l�ڹY�������V,�d�F��������o?��튾K��+�>�~�Vs�*�a遧�������={��d�3P�i��s*�#��L.��ն�Q�߅�RO?0��=�~�/~��36�n�0��+\	T9��cY�(:���rwT�����#�de�a��2����v�M"�-�WE1��ti��6f��{�:ϼ��T�u�~�>��9�W���`��������3���s�L�1w�b2�w\����u��?-O��������^$:=�C��ߞ�}e��R4*K����S�}~R�#��yn���`ⴏ�*�}�IE�@�7~�>�`h�E?�"*�e�.�2�Mq<�N�R��	��G3�~b��T�/K#��u݂�}ʤ^�<�,����z�W���ݻ��;�����`�5"e�#CD&���Ǆ=����Ǡ�4��S���e��P�jی�r�>)a��n��پO+��P��բ�}{?�=Z.|��x����꣒7�5��E�֢S�(�0��x�oV�^�ٝ溁���g��b���q�o0�����ɍ<W����{[j:�m���	���zg6��Y����G�3e�S����� ��(�-Gi�����|�·�h���pCV�X���A�T�$�{�*l����!��k�^c�٬��[�m����>o;y�����)�ǌ��B�5�·C��`�eoc�O�4��*�kR|���\X�}c�1��-R��*jtf{���}iz��r��7A�ad��%4�q� uS��ɉ����L������ôYM#��,��Nj��v�IX���8	���ڼ؀�[9j��;MdN����n�������E��5�[]����Z�m�8��v�~��Sy��Ӛ@�;�^Y���C'���?<-��l�a!p�J��:�xg�N���vQ�`;�jƀ]���^�F)�3���~�޺��&����a[d[��.�|2�&�:Q@59;L��^L<۽^@��x�S<�O�����h�mպ9�e{��U{c/h6���a
xĎ�s"/�5w�U��+�CSs��SvɠH9�=�x�~���f�+]6� ۣ��7�G8d�0�C������~��y�;}�w1ʞ�����T0q��gʬ�z�)��`�q�S��I���݇"�.9˪rA��h�?v�o��a�2�me�%Ib�Ȣ�Na��,���Z׷�k ���]X������D���9��ı�eeu�:�2�i�ô�kFt�Q�ղ>,7gkH���F�7��67h�;ӰS4��S�3o�.�
�#R�0��yճ�����a�MMY�f��0/]��d���Н�qT���mcV��������&)��1X�M˪��d1[Ξ�\�.�H0Cio-�w��̍��3����jg9�FX��V�)3��G�A�PVbIGg��!�Y��
����P���	xP�iÝ��Y
�8�Ŏ*9z�m�6�94˪�{SOWۤ�<�|/�����۩����%Wf>�8�YTk��TNc����ܟV�s�L;�]�4cʬ�8vtm�έ�9��U���b��z��r�r��0�"8ȡ�z-�[��J��r�p��Y��gfuh]�V�<9(ˋ�fWUhV��F�:�ɉ�kfE�/v�1�M-�����2�mȫ����2�Ao*Z�{wU���G��2��q;dCy��,�i�YX��+y���
�졛\�M���,���
��VwX�9c��[�g�U�8Ŏ���[�4T��]�A��B"Y�F���ԪT�E�JXL�C�b!�҃s]�=�X�)�J�����%r*�1�:&-S�ؒ����f���VH{�BPE�]���ܪ��p�9��c���:܄#FW(p9��a�	B��9:�f%7�s*T����!���������-J�ӥ��ꩨΎ�rxt���G�Z6+g7;����c�LW"w)N~���K^U�8��^�
3#.��';+�y�kn>4���a�Q��<��itV�����yުz�L.��R!��S^"��W{��g������\�ڛ��͎m`����Ԗ_[Y����#��`t��a|��������.�.7[�Yhⲕ��ލR�f��*�I�w;nq�h!�H�<4=��*P��.�X�d�7�;3�7�sX�2���E�\�����29��R�+m�H��S�#j���#�/8Y�:*��Z��l�Qk
Z�JJ��y�e��38���4�Lv*�ȬU}���1)n�Y�:�T���w���:p��<l�o:]�bu"9��v�>�.l�\�bB36�U�1v"����:�7o ʖy�곍V�;K*�y'R�|�Q����"�%�3�rl��:��p���pS�OZ�.oU��n���KL|;��r32�=�.�4���T�J�J�0s�ap�R�w����bY�t��;|*������'bB�hA$M���@,�Q0�1�����ת�`�FcB�B3"QFH�Ai3�Qm(�d�Pm#�J�!	!BW�&�pB�(AQg��^�7$��H�XS&�������LZ���6� \N0��C�Ϯ��}�5�c���-c�A�\���dd�Ǧ��>1��kZ׶�>>?����ޜD�d�#�#��sr,{^�ܬ^�n=���>=����kZ׶�>>>��|�����8ر��uۺ���u_�׫ʞ���^9k��"�s��ק�ס��kZ׶�>>>��O/.�7��`���9	�s]�������x�7wo��ɹ�Tr�|\���h�ܫ���ǥ�]����w��|{}�kڮ\��ۅ�\���Ѣ�b�G913�&�� ��l,9�͊�$7Ȧ��/K\ֽ5��b�t#���-�+�?�د��7�V��[�F��b��m��\ŀ���71��gѳ�94����WM٣N�R��;�u\��I��ɺT�r�<��!�; j�W��aYύ�J���f����8��u�C�"�1�Sa�RG"q��)�JF~x�����$4�|MVs���8a#u6����@�0_3��4�绮���Q��`�ّ�;�:t�`�<��mW�-��a`��P���{n���X����o�g�4�)���#�̨Y��l
�7}������w�PI�MF�B�����U�рjQ��U�q���{I�IƓ��xSTK�,l��bsY��n��6�h�ߣ�T�G��E�r�IW�LG�Qscζ�8JM��Fz�=�l�`�<��\�J=\%X�]��*H��=F��M	�{��o�C�)��z�WB�l��]zQ[��<���g_���N�q~z[u(G�I��L��m>��5�Ԍ���a�da��x��$NNʦ��ϴ��Ϟ�>78_Ն�lFB�}�����(]���z�.ٓX����m��VA1�6ʪ���Г�xw>Svf�J�kd7m�*�_��9�T�F�X�����M�ò�ށ��jm�3j���H�\��޺�şb�B|�˺|��\p^��N�䁛�b5�/�H�	���Wv��N
����青=҂q�I\�r��B��*�G+?��n�~��wUu�Ę�m��螽v��oy������ò� ��`���m;��=�MP�\����iV�ކ>�{�fb��Ԩ�SvL�or`�uǎ���h�g�1L̪�Aݛ2���=�(�J®�EN�	J{����D�U�3͡3�F���̪==�|{Yٙ;�u=T�O��SQ���wp�ӛEٍ�d`{��т�/;��
�B�#E�E�M�S��ތK���	ѵ���.jt���d�8𨬧�#��t��h�{M�G��c�y(�D����Z��W͞���\E�κ�n�r2%��]˳���Y��~�o�E˗"~�`=�A��27����{��=�����J3&�lH�3{�#2�DAx�|�c��Ö <6�*�������'Y���|��Q��}1.�?�t-��K
,���?lU�Q��;��9���7��qk��o�"�s��u���j�Y���J�[0b1O�+zv7���n^f�~��닍����p�gL�qc��^����rM�s�#�®���]kG�r�P݊Q����\����n�o;�f1{yHM�OJ�y7���o�~�LE9o�^��]L㺵8bR�/vA6H��}�2R<�N�e���o7��o~���)W%9"Y��{�JR�٭�Z"XSĎ�)ݘ�B�2�v�m^�ȉ5Np�t��=�q���hK�T��RI&��7+�)��84i���pؚ{Փ՝ݜ�h�cǳ�|��XK�<ާ��*­�T�gl�_W��n�N����c���v�A�	8`����vxY� R=gczV$�2��2��ޣ�� ���%����`�e��@~�?c0n��1S�}�ʄwkzE�2���(���ߺ�t9wʆ;F��ƞ��zn����@�g3��zCO~�V�&T����\��ʹn��l���Tw8�K�t��R��?��7p��uCxy��=TjF	�2��Y�ٷ�z3��ܧ�v��>�u���9��0Ew�=����ҋ�^�,G������T��{{{C냈��ӟ�du�x�Sf�[�Z�y�O#Lx<e�(E��E�ۮ{�ω3�4Zh�H�kp���~��,@�h���-H�	hk&i��p�	 Zj;u�]d�v4�ӆ�Cu����K�B��w����nY���� �[��H��M��v{�#W���o�A�w��o�������J�oy&Ɨ���d����������>#���������?7T?~ �=�q��0�Ɂ�H������^w|�h�y�>s`Z*���G�s����i��M�CP��U#q��8�ΓY;���^7*�����nt4D��$�vZ>6�֝�ٺe�,�ń`{���U���S�1�b��:j��������aJ=`#�x;V{$߰!�>�t#5�ܣs(�ub�f��m�`���&d��N���ۜsLb���ሡ��|��++�-E��<5�i*�0)!L����Y���
n�������:�C33f\�J}��J�=Ғ��%�]����<n��k֫�/}:x��;��C��I}^�1�0>�N�2Z�FY*Y��AXҨ~὚�&[w��������[��!�{��y/����v�tt�����*m;���ZF0m%=令{V3�<a�کf�����"�N�(/�2�hc�R�M+�-�Ĭ��X]{���g�D;��q����,�{ڪ2,�����IZd@e2[���6��tID���3xV����3Wb���U����鱓��G�"��ʼ�i+!��˩�aB �ŧuvI�訕ȍ}��#��x����(��/����4~���?z�����J�:c��^K,�1����S�%:��9����8α�9	o��s�}'u�s��E:�{��k��|��w�$�uȸ�,�z6�-�;&�!���q� �kn��U@}���$�[�TG��4&q�;:�׬�V����v�v�-�Y��o\�<0���B^��a���� ��g�@�`��)��vkdo��!���|ܔ����NtS�=�Ĉy���w�}8�G!���nN%�7]"�{\�㣹R4���7Ȫ��H��j�S��,�s�L2!��冺�I{�Ogj_ݪ��l�F�'%��@��15���qK4Ȋ7-��A��|����G�X��u����f��>&�t� �T�qK,�����&����^���4����W���k�4�݌��,�:�Cɞؑ�D˵]U�TM�X�kt�'�xl<�[Ӯ�e�z�zS%G����s�r�����U'6;��o�2�#ɲ����T�}gZ6(�"���̾�e�YZ��Ş���.�׮�"ɜ���
w�Sh�Nw~�����a��x<��(�*r����_��F_��O�2$YJ�PoC0��eת(F-|����Vd���gH���������ݹ��2�~��q�����)wz�8�Rl׮�h2��G��x����a����mF�r��i+��U���uC�4��2:ʪ�����<��p�R����������b\�5�;���u�P�*Fwf7:j�ܹU��
wtz5��ώ��EFV�+ͮ�d��-�wO�B3�;��2���}E�|��WῊ�����)��c���9��HZA��Md��hT�ޏ8��z�Wޚ1��r�n��l/!k�˖�{�d�fצ��oGj2h3x��.�����1H�_dZ��}40e8 �m�ҤI/�'��m��2tYJLcKh���Ϙ��G�wM0m�f[@�&x�$K��Z��@�� ���?1�<�x�e���3�S�P��h�����5���ʫ2�[�e�$���B�S�x.�K��Zڙya��;�����'� �M"|C$��:L]�G��<'k��Id�ٖ�`6�R�L]�����4�[n`���Ŵjb�{3�΋��y�����(�2%p��|4?G��f&��n.�<��-�x-,��pε)�խ�'�� �aF'�1�Ӻ�_33TH��=�(��ʨ~��Q�<-�x�P�M�B9�s����3;��Mcz��s��X5o�����p
�$�� �E�Ņ�9��v{�\�՜�W�Fz����u���{�[Y.mYZ\n*��@l6����"�3c
��c��8�'��ܩD�}���P&����>��z�-���Du6n�ΛO(g��pZҼ�JN���VT��u��	�u�nEp�Uhѻ��xx>{Q���jI��3�.	�]q��7�^��Z�S�4u���Gj�s���	ɍ[}�� ���]gc�W����%\�������jյϦ���jP<���_�ùR#�^���%"����v�d"�z:��;���>��U��Ϲtx�������#�"ne��֜���t�c��tq����8f����2�Bd����'�VK��
}��sڙ�����Oi���gHǮ�
���D���7lk�mÞ�p�߀�wvE_U.x�m�\&IvJ��1�:��r}�gJ[&d�����x��پ٧(���W�$MD+�&/%W�ۃ|Gz�,13#�2����,˻��q79������<���ޞy>�5��(�Z���+�0|
�/1wω$�H=��H��v~�K�y�32A8Ԡ7!h��(.z�XW��kdr��	�����W^�Jl[�p���a{%c�R
 <��╹���]?H�j��~�on�5p�!|�R�4U����WE��]�1c4y�j����N[���{��խ�?�e�>���/���U5�iɨs��=���b@:tl�4�q�ee�(�g�n �`ȶdKL���;j�Z�Zl���LI��Cq��
iA�/��ǯ2���
�c�x�qr�z'��h��ѽ�n��g%�2py����L�ʹ�o�[��	m'8Z��-5r�Mz@�a8�#5���G 2G��9P%R���@��]�]��0��iٶ_a#lRo�ٱ���[��<��c�qk.�Ƌ���8���$[�M�G�N������d�˄Q){wj0��`���ک.;3E�ɶFp��(]�=���Z���jo\j��L�ZY;�X�IT��v�l��5��Y�(1�N�A"�B0�P�H!��^.^ׯ������ 1��)Q�w
��;��;;3{�l+�f��J��	����}>iR������{�9�zr��J��^������	�hZ�&_�sж2��1�ٺ���{�MI����`,������5�C"7�е־���J�t��Gd	�kz}�4;SA�Ս �e�����[>���n軖�������"6��*����WrW�Y�fy�ض�` Mb���X����N^�v���2t���0�wN�j�'���v�=�2]��J�wZ�k����y��vb5dxQ�im�^$�7\�@֪���{ͳ-�r��z��6C-x|�x`.���8�pc��q�k���I���:"��G}�p1*��}�ӏ~�~�8+���2�GD`�g-垼*��&^�d=
�O�����Hi���H�y�[j��247��(���ÿ�i����-Р��Ua�M�Fϣ�Ō>��Gmp�K#%]��l��3��b6�WN�XQw�;�"��L��e+<�|�bY��@�!@��h��:�������Bp[��۟E�ǃ�2���+:��T�X��z!kz��S\�j�^�^^>>>���T줺F��"��ϩ�V��	R��d�U����M��8�u�}=ÃzH!;��lQk?�i���^6{&�q������+�.j�?V���N�`W#��"!R5x٠�v�'Ƽ�����~��ƈ���&�yr��fעi�i���r����xJ��z�w�aa�iJ��4�Bs�m��c�roՑ-P���8�p�D��χ�[~�mU���;<2���]����V�).:^��U96�w~sW���*N���jǻ]a޿��=~ў͵�LQ�T4��a��y�A��ey�Uu��8g\�#��$�P��fD/r�Z���5�z�E��JV�3�������j�u�j��޺�w=����-�U�t��&Jrd��w.U�]�(*ݹe�`A9�����l��
'� Ῐ#�b3��SfT��'�ݫ${����y����ۚ�켮�4��n�;KWM�7�I����{�F0D�%�Ye�VFj�w����m.�jcL�J��mE]XqA���ɒo�m �S�y԰u�I�-Q"��׋Z܌i�I}�����S�g�M@��/U���ʈT��4[A.�����zBkUZ�Q�al�d��7�V���Z��[��R�3ԏy46���A�J}u��i3e�0b����ιѓU�I�l��ݩ�g]vco {��Y��,T�\9 �E�P��Q;5y�,��eUTڨ�8�o�h��N3rf�9kD��y;���w8����-	[E��٧6�3MnK���u�4�n���gRW���\o0ֵ���2��a^F�3\�̼j�>�f�\�WYBnK�Hҳ}�Kmf9%Ƶ�:i��	�^����F�4,�o�OS�k��G���02s���Z��d�[$Ţel�WT�E>�]0��?�m��A�1���&=�Y���Or��˫v�T)hxq�	C-��l%n�1J{\��&�U���j��;Y���z�!+ks`��'3z`K1丫��P��b-s�6�<}��F��u(��q}��M�Q��8�[�UV�#3[ʳk]�Kq,+w���9p��<x�N��-�Ww���Tu��lu����}}�0�?��O�;�gW<����IV-�AK�\C�0��?b
��?,oyW�m��j\��jav�����n�� )6�Q��y�2��$Sp��)�nD�{��-){�p���۪T�v������l>[XS�=ZM#[�a[ەٷ�E��[���R�V�X$�-��ׂ���*�}��}!�o�(1�Wq6���=l�ӰL�GeZ���9����%���&q4���P�O���pN
���2��c^�ȡo�N�Ś��hq�y��i\�)�gW�u�5���n#���i�Og�e�֯d����,��Jۮo�Z��u��fk��/�����r��ݐE#D��~�rnj�{w�s.��B�U���Y��Q̖6d�R����	A�v4t�����'��g���A]�εɗ��DTs��բFέ}���W1v�bXn���%��m\�����w;/e�F����XS��L�3�
Q�±�u����y�(.a)�������a^��3���L�����ӶS���i���m�k�[��6���]�P`�3js����3&���/z�.��{���ٺM���Z��|n%&(��L��5r�V��Ф�i�,����f��K���0�	4�T�u��89��{���q�5��_] H�@$H>�������4�����}o[ƽ�o�kZֽ�����}zyysb�����&�jkߝ�Bǳ#$ )!�ǧ^__^ǷƵ�k^�����>�<���P2$$�!�&ܮ P��s"��$�o����c��Zֵ�||||}}c��ˏ0�H2B2��_n�A5�,��1m���{�#DQzn��]B�5}��K�gH���1�o�5��o���A�7Uv�h�ME�����C����mp>9dѾ������K�/��)z����"
4X1�\F2i���!��D4h�ɣI��۲(�1�S�]�b�$A!�W˷y�9�0�|�ɺv�TuqˍJ��ݓą��Ua��c1���JR�l�qڶ��@�ݗv�ߟ���y��w�-��1��ݑ���5����+�����@4�^�1v���]1�i�������\b�{c�!��`�`\��٣B%�|��yW	�4[��3O�JA.��?�Z@�:�@��bev��l��4:�D{�9���J���t�3;��8�	/�=c��2����?���i���99�04|�??�sџ_�o@�N���ݾym���\'�K%P�A�5{�ط�vwF�˙�h���>@���NT?D�z1#����xPQt{+�~��V�ﲪ9'����h�ߩυа�y�:U�"ס��ڜ�nw�
�8�H�8[Țk����U����R���7d܇'<iޥ�;򙽗�kZqH^�t�9�l%D�T�*m���P�0��L�TtPNH����տc0m�s" ���0�ypc(���rA��M�����B	����[���GT�ʳ�D���k�Y�����z��B��b[u�����*�=/�RrҚ�Y}[U��!�_`{&�4ve�u�n7����N�T�:�ǣ3l��ܮ;�Wg���u0�c)V(�n=6�?+���:�y�������i�炉M?x��K&8g�wWD��$��+�Җv����玹��w7U��=�[���Y6�kz	؃��o�Ȥz���Z��EF��,�S��^�Ew�J�}�N�\����~���	��������w�J��!)a�9y~n�;�;��k�mƙ)ݛ���q\dDd"����h���ݣ��=�|=��xU�-����]/u��۾"/�Gl�f�z�p�����r����J\m�T��g�Pҧhz�@m�������+c��gwb̀��BA�Mw���tg�`��=�A�=������n�H9���5V���ZS��\���H4����������i}�o�p�����x�A(�lx?R�~�]�3�/�<�k�=Q%��T�vwz��� �?�d�ا��g��!
�H�tpƧA��#O��׷�],�q�(��6�O�1W0��9\�(Zʩ�U�Q��F\tF��T�����Тn�a�Zl�im+)�J�1�]�k�G52o��˺}f�nu^Ʋ��f���ķ�ٶ
��%������i�T�Co�uva��Q�00m��(
7��������.��˥R���(��f��}=�W���IP(�fʣ�
u��gŌ,����ģ꣯���/�,HW@AM(2/���3�{�L�m�9�^�*�ov�d�Y"���\��o�o�c�N�%2���NM�C�u�T(e��t�w��/��tG�{?pC"��
9 2G��-�Ru��=*+9�*}���V��c������ϱ�g�5��,e��g�5h��t���W^4��}ܧ�����!���O.&�x�c� �l���O��ӶI=�o�Mj�l�W?��J� �\㍌��S���r�G������Y��*L[u,x�X���3ط�^�=ޚ9�漗t��v�k�M�Y;z�U_u���v�܌��$� ��DF����zpw�t�IPNHֳ֧�nhV��Jo����:1G�])���p(ߏ�ֱ@,�ٙe�p�SϞL�&�T���+��bP�huA�m����>i��lY#�ũ�i��z�Sx,�l�Hڛ���V_(�g�G,��pFXf����]��{D!����Ჵ�3~��rԻ:q�=W��7�}�U�"�Ź�w�6��s�0/G�?����<J�*s���6}�����^e�g#��%�ӲN�$E-b�uy��r�-��"ـ��=�C�2���q��� `O�uWB�X2!�2{`��UP]Fs*�t������nTE��O�Y���C�\h�~x�j�ו���+{��u��u�>��Qc����������ϐҶ�]c^�C������Uv��.��xK�J���U��p�T�p��ݍ�M��w#��g�w S��N*^���ʓ^(�#���!O��N5�ٯ�a��!��l�)�.ޞ��L���ܥq�����tw0�i�g_�Ό�w��/ۿF�L]�9V+�����@�S���7�"ܨɉz�._n�Ҫ�U��s��t��S�`:�̉l��Bf�g�b�ZX���O꾚|$�� m�vzOE��SyXnx�(HԶ��U9�������^.��6�O=:n��w�̘�����L��T�eIg�����x�Cd-�=!o�w+��c���GȄ @@�u�乕pd�K�/��uC�f��On��f!��}��*�#��N�b}l�f����'R�Rۺε����?��x��lI4%��<�GN�
E_m�%��S�j\�������9�c�_����q��Gtw:�^��}�grP��T�t�%�
���gSќ�S��0u1�k���1�v��ރ�����׭w�8�"�7/�&^\�3di���9l8f�a��.��lǥ7qYM��~�����Ĉ|G�Y�VY���"Uh⁙�����>c�u����㣊��b��R�-��:��Mѣf '�������ol�L�686��x|�-�z�c߲�jg}��/���G�teo*�H7�����s����m٣07��wpV�"O$gG��Uzk8��`����	/Ew�1�����/�ع�z�
��O��JS�\�'�A�������c�
�:3vgz���i���O�{�x �̕^�12�߽7һ�W��T�j�d#���D�;H���p�괮Yy�1Yĳ^�\��f��5b�㞛�}�ڼ^՚�~K����콌�wt��}ǎ���%����"Y�kM]4�p�C�fd�{��گ��]%0Z=§tLe5}�ŉ��,�m���W�~>>>>>��싣�/��ΡZ��צ�ڮS�z\��`�z��0�!ZQ=��H}G6����9�Ҋ��*���W�^\K�,����;.O<����'����+9�Ä���V��va��Q%	w��ޞ͕�$U�8~������n;�x.ޘ����b�o�<�%R�S�x��.�,�)��]N�Yx�|X8�� �}
�{|��ǽ�<��imҡ��U-�"�:��ٽ��Wz�M�l ]�,��]C\�H�g`pw�`�\�#Kv�w.��y��^�m���o�Ϟ�w*c�B]s͡�r3�u9y���L�oB�~΂{�<7����4�xη�[��p���x�)��v��������L�_;�w�u��1z�V:b�7ֺ�y�/�t��0-X�{_��j�2 u�g�ad�����^��0SR�@�֮�z����\A��,f�7���9��{k���<��{kk�՟���B��#r�����t;���j��&�E�o#	����&SН��i�$���_y�`�gp"���ɦZ2o��p�F�p��(��^_S��q��X���S�C�F�B�l��L����C�*	>�������>U���(Wﯻw�2�fy���c�;a罆�07֛,vq�u�]�/@�Xa�ԴCPd�*��J��q�Pkf�V{����Jo��E�s������O��*n��
:~[W��v�
��Q t���Ry�8-�D�{�����y�fa�s�_;Sqq<��[T_��ϲY�tA	�U#T0����� �ō=c��{�ޭAh�IW�9~|�W,���P�X��T�� �6�g�Q�>�/ʷp��s�tH*�x�K��\Ә��[��Go;;�`�'��*T��ъ<݆���ov��T��J�A��-�n�\���=��ٖC��G���'z������"i�
���2k���3D�]�{�ƦILb�+��e:�W��U��J�P��r�H}�w�����rj�v��d�]D��x�p��!m��w���o��'"����_�r:��u+�'��W�CR@F�����o_P�eˍ��;d|�
�8�.v���>�P�[e�����dK�׵ֶK��>#��؜O0I�]t/�N�i�k���l���zX+���� ���r1wPעU������\�3F�{M1�7���T����`�kL����s��i�ƍ���XKl�y�z6�϶�������ՌK�x�����Mw��ss�>�-�oϻ�"4Ͻ
zv4�w +�3]&��,Ȫ�ʝ�SU��]m��}�`�:|�"��"6〈�v��e{��GDo0~�R�l��c��r����n��k ���7��8"9��dz��in���v�?
�n'�%`�~�@w���C�g9�)�:���=��kq!*ꝣu`w��!�G�{R�t,�����i�2�聂��W�L�� F\�>Y�{�w5^P��gt{������=�9`
��Vs����f��k~=�#&��y�U]�.v��~�{�+��/."�_UߚUXfE�FEN���u;�CP�AU=Qg�]8�H�#���<C�_y�H��L�����U����k���Q�7����8��Yw�23f[w���óX�s�;�=�ƱA	�N�Y��Z�{�b�����ӑ̓e�v�ǖ�<Y5Q�n�t�$�V]CE���7�SM��v�����x�����V���䢅oCMK{�y~��3�n=b7)G��j�k�8�U�V��ݝ�=�2L03ʨ���=n��^��:	�g��4W���Y�/Yl�lIn\z��U䊠a�&��Ԏ�u �@�i+Ss� 5eE'������o|+��c�ϥ+Ғ�͵��Ng1�]�	3�,��Hj7�Dvm`���ïhF�vTr΅^�J�\��PFK������n쳝����[^�����"uW�m��؆dr6�8�%IwT���$7m�<�յΕC8��3337�d1p�Dt�;��B��}�� �s�v�A�'v3`���ﱰt�[3p0����oso�V�7�WO`B��s7.i�{��}'O�a�cҺ<��������X6��B\[9��u��p�=K,���=7G�z-�y�H}&A����Y����u�r�.�
��aͽ�M�q�-���>'e
��\�86�v�>�������4c��xfs7�w�[��m�xq$�2��c^|���]`M���+�ow6��7\��eLٻ[v�Q�KR��v+]UA����f�V�{:O�����||���=+᚜����hUe"{��I�buyzWR۬�R��\1�j���w��<!��������g?�g�H��̠��|R^�RI�Q1`�ր�&����7U!��3C�É������ɯ�A`y�~�C���{����V�˕����՜��zr�U�e{]�-策��G����ܚ��~��8��wgQ|�܅�܈�WF}Ǳ�^Q��;�Bv-���(ڤ��3N�{fZk�w�bH��:�Ԓ����٫4�j�����+.�1+ �5=�=ڛ�[�6��"��������)QG�)J��;7^m[Z�vnwz���M�!y�1��D�b�x�AT�M��TM�B]N����gTd�Q���#�6x���`#�N�rIEM�S��.��7�
�q鬅<���G��E~�@hd��-�ճ}i�)�[�D������R��0Ң�yXQ���)�4��Y��1ݺ��Ziwm퐻r[��0Ess ��_X��k{�5�����oN"뮡u����Yv�̇��M8�7�j���Ft���=�lݝ�N�݊#��.�CcU9,���ȶ֊7����\QͮO$�MY��9�M�X;�rǝ���gv�E5���2�W�m#�a�s���="ւ�TrQ�ƻ(����c�S{�]Y�8��J��d�ݡ"�^r���.��,ٷ�����2�Pq��,�]��,��Ɏa��\�|,�WOk+U�[�]��gق�#/.�hgU9��N�]��:�(*Zs�[|��-w�X�k�i��9�r���K��a`ʋ�n�	��y��l��q��;aΓ���������6駡۾����m.LGKW�#8g70e�2���<v�]n�<՝Ed��)z�'WTq��u�T��oU&#���g@�GN=���kWu��1]�]p��Oi����Eì��C������ܛxF��oj�Ժ‑Zb��j�\��TpYwXm�	&���2���V���?-z����Җ;:�� ���zR�]�J�[K6μvL���
��7:<x�Fky��5�om+Ud����Τ��4��xz�<�g�k�ӓ�8�Y��7�p_T�R:g�S�w�rL��s�^_^��q:	�d�EE$	�(�Ͷӳu����6��c���u��%����_We������Ι �e6h�K��n �/2�̢�-��~#)�F�iά=�j[$��_bԗ�u��7�2��#C8��f9n���-�u���"Ҫ<�snZ[;�^OH{&f
�FY������\��OYO�U���*f��/;�ܛA��a��rE��KƇ\O{��<�^��M����`�n Wn����,	�F��s3
���U�8�ZDws�����:���5{otVd,��6�/e�[�^�-��O�k�3j����5�Ӕ�-)5P,�j�:Ddd���Zkm�p+.��ژg��:,��F�PS�� 9��Dٱ0��`5��J�:��R�_PC�a�R\�x��Y�t����3屷����w������3�W�B�z��'g�'s��]���$)��;�T���n,�A�tA��S䨠�nŐ�Wى��G:��edUp�s����O�I{�s1+8"�����3{����b��}(�_V���ݧ�o���S3qԲ��u�cw/��*�c�u#|��E����9��C&b&So�Ӻ���;r��]>Ψ�+�v��]�*(h.%�|�;+�s�	�|�4�e��8�\F��K3蹈'e^F�M��2b0��1QpJ�]k�)�YCVҬڠ��v��܎[[󏔝����䍈Sp���$B�H���$��>�!	0DУ�Hd��$�A��Fd�KD�Soʞ�sƜ�@�0�D&�N0��&Dm2�-6�	bb�0�'a:�Bd��?x�A�Av6,On�S�Qb(وH�� p�ק�ױ����kZ��������///����<���$���!}���WS�A�a	$���^��^ǷƵ�kZ������Ǘ���y�I$d	�ɠ�|��2"	/��i$�c2�y�w���wC�Zֵ�k������ˏ/.�
�ۑ�Q�f��R��m&Hɐ���FL�F��$ h�������d�i��ϵ���	h1�26=�`�)����7'��Ā%�W�]E˘1�I�M$L /��Ba�H0�!C{�2e�;v2II�$�&I�Fe��`be#@LaD�oݥ��﫲T&%��3F($�g��HD��]��Mҁ(�!��&
^���&%�@,�O�	$�ڵ8�;wQ�ې��*�fjBG{u`�-�}�ݦ�S^�v��|�'m]�9p;�x��Ω��Ǜ��uծn����:u^�J��<��t۹t�-T~A�{���01̀�$�M;穇zN'��\_��F�<d4cQ�'��?ǯ�{���^E9��a�[d��K��)���'Β^w$\��n3�!�ez����[�$���I��o����)��e�K��~s���$�n�GC�j�w%�Eq
�b���o�:f��KO-v��7����c���]*vH�ŕ�� mO���V��"j�^jͻ��s�����g��c϶\w�e�\�w��=�+ݒ<"!
&�잂ע�=�I	�=����Va�Y���X�ۮs����l7�s:i����ޝ=��K>ؕ9�����t�E%,�����������s`�]�<�r���瑝�z���U"՝��y��fM�s~�}��7}Щ�f���U�s{��Z"�mw
.�����񤨣��+=t�6[�+��?�9���󎅈��{�����V �Ԡ׫�b&����}Kg�fÔ�'z���53D�me���Rk82�w�ʋV����o,��Ӆ��h��Љ�T���"���b�*a|��*VY��\��7r�Α��|:w�0
\��8O{t����H�M˽������/���0��J(���^>��!\�W���(�� ���4���Qm��-��wew_	�ɩ��ߪ������ѿVm4��d�	MC4I����;GgN���}~I*c&��@��Ǽ�@�yx�U�,��p?-3Ԍ��h�˦������j���bh��������xۏ/Kp�s|AR�OKA��}����i�EO��f.S@sK���Yϑ�6V{���RK�R�lگEH�c5G`�q���:�#mluϒU�"dj���!���\�G��:3�K_�l��/5�T��>s�67��rR�t�Gm���%�R�8�R��*��~l�o[���yw�"���;��Vmæ�3f�lU��G6�����v�����#���e�� ,��1k��dܫ���[�����ޅ�+�����8f�=�鎐�\��~��3��t�Շ�%�ή\,zKK�u���!�ۆ��%��S�5�\�LL@���(�ʱv3�PG�tQ�>:�
�б�MF��r4�]t��]���s%��ܾ��{�Fӵ���92�W��{�|�y��3�>c��9�3$�L���ׄ�����5�Ҟ�R7���C�	��z�8�$/��_�������ɲI]?X�c���^.�扯Z{�O;��(�����Գ�ſ=�5���[,�h��ȥwʁ�g�w����z���	w�Y����ވ4�Y����i[�-c��P�S��=9@,SB�����bx�40��#.8�M׆hx��G���1�a�R0�
�X�ߕ#��[�gm53�+�Q��6G�0�I�I�\�����t��[?�݅�+�
�e0�ȋU�&�_3N@#�ݵ�=��	P�T�&��R7-��c�="�7+Bk�.-�4H��xӽI�nu����t�5�Ĥ&��=O�2�NXfX��W&0��Z:Zl�;{�~ r�"���7+�E�)[ϸ�Q4�&���3��}u�t-�Z#�M"Q}��j�{��2U�"��Cڧ�n$�m	�����fM��}#���P��.{�������7��l�[|�Ve*,�B�%� C��_5}v�i�U&ܳ�S�'\�w-�i1����/֞��O���=6���do�rfnq��]7^�����������xN~�z�}�NN�ݐ|㡟q�\09�yܬ���f�)�8Vf�^��;�+w�BU�&����{�`�ox���p�H�Đ-*���"i�5��\�[�������t��u")�������gC{0�v!�&�Ka݃q�\r��:��� z.kG3�l��k}^6��sg:�{���lݤ�f �P���h	�t
�į@��H6Ov	禎���V\��H���m�W����j*Y�J�{�h�=�� �.}hkeW,�m�V]�8*<5��E�p8(�,�%>�(�6#dz����������^)�'jV�t�ٱ��1	��{FG:Lk*�k���v�Xk�N����J�ד��g������=�9��JxY�i���u#���8���ez�e�:��]��3�m�
i��R��ʥ' �������Պ��/=��w�,g��=��#jeu�ؒ��%s��-�l�çL�����'v����uY~�?.^SWu����-sS�Q7*����U@�d�H#��yq�`�%�e�?��!��n�Q�"�pޏV��Mv�&��0W�I�wħ�DU$�n��i�������IV��5�z��'�#D��Mz.�"9_�� O�'�UY.n��l_�t��4�w�i���S��9�#-l����%AJT�5��A���k7�o�5�cA�g�%��O��L�Сp�.�ו��� �_m
�>1ƣ	�ބ��l����q��\9�6Lh+��''^y(�/�4��̪c��;��la�ٛ���Y6�N.�pY>�����3�=PVpșoks6���l����GO�:I�aw��t;N�/�"��G����\��f��w�l��9wU�|�W~>�r��4��%���ƚ��h������ۃ���o	m��S��;�azV?rH�ya]�
Tz5��e-�}����x�Tn,=�4cУ	N2���)�������z�^��ᗜ�zBff�H�B�����3���6�w�D�>x��}�"��h�9�|4�c'�-���5��DB�Q�'��63G�&x��@ ���1��=Q��W,AزRC򨢿3͎�����J�M�l:���#���r3������\]����S>��|�>��s�և;��-�u��Z���6v�;�T�\N���>�2U��9����j����{yy��ޞ>>>>H{ĕ����%�	���łorf=�T�S�q��[�s�����U/Vҹv���$lWU���=��|uo��"(��80f��'�<�eS�n�P��V]>�q��iG��T
8�3iX˚7!
(,?�&�s�:����RPGOz�W��Vy4���o�hhێ�k9�K�:��74�B��б��������B����0�5�w-��6����L�UΫj��'4�ج�G6Mhp���c?e����q\l���#H������Q))���N��K��&�-�ӌ�	ۯ.�i��g)K:8�J�ܸ�l�'�_���fp���9��z�;'�����n��b�����P~���ϣ-r�^�!w� [Ϡ�y���lt�ֶ!�Z�nl��DB��OL�����2v'�e)�%�#V5:\�-a+��f{4cy��ÖH��A���%�2#�	�Y(߱)�1;��t�{��jl5�`��_6�2?\ڵ��0==n޺!�c��H��ɸf�]��vMs���h7>���[׫%���(�n��4q���}_;�|b1�s	-��x����;������}�댈���kk{zxwo�Yܤ�`�-��mݝ�:�i�U쪹��.^��$�����F闶]�,$���������߽���9�BP5U*�T��_�k3����1�Wiq���ѝ˭�*ēٓ����Φ�^$��t���g���BIC]C�������z݃7����ek�1�m��Ol�l2H��6��cxC�-�����pP�<oHy�U�/�E�{�%AI���ܺѡэ,⩘ʌ֣�/r�y�����8F�P�d��]G�)t/x*����	ڱj$7T����D��V��+���ǃ���UGX�<�ח*w���[��՛�ҰiΡ���H��xr_ �Ü0½&�Ym!߰C�y]�� ��m`�Y$�U��2����ff�r��:���������yd���;CA������&������1v8�sΙ�\�A�_��3�n$��k�c
�A^���oj��`�zb�TX*j��Md�Ȍ�f�ֶ�$�8��Ф����<��q��X;U�`�U��`�תޗ@_�?����y�x�Y���R꿻D��}��v�zuXId�&��܀�v��fK�\/;Kv��;Wp�tSV׸H�y�K���mҒ�2s���EYwv��-o:I�N�t�kgv}���[�܀lᅬ31e��nyV�\l6�hm�j� ��Xٽ�}"�v|b�?�P�<�q�uI��V�W�a��N�T� �Y[�{x���t�Nո���cj�oC��uon'��U��UJ����N�<Un'��[�o`t�[3s�5���͛���ce�i����2j3}���D�겜sQ�G�G�gzz���0~��4��;.�ecE_?.��j��q�6� �K�������O92h1���ʫr�%���0k�<u�SK��eb�Q��3�w��ٍ窪�����i���r��]�X4Y��U��o�-�z�
�B�ym�S��+iS윳��5Rk��{�wy�U*���F����'o�U��H��.��gHڮ Y��	'"�0}AuN�VĬ�$Ƃ��&�F�^R�����M���Ш�Y����Z3/7z,%�m���S��*E䊨�bI;�R�b��R"Lm�'��Si&≴��������Ֆ��@���4;��ɈfX>�W<x�>�s"��b`=%15=B�n�J�~&'b;�.x�3�D��j����E��=z�l�=ܮN����^tmNα�{�6�-�_��*4k�z�E���e[��gS����6�z��aծ�����k���a��� ���Mx�d�-���r��Vs�}�v��mp�e䅐#*m�\�o�&�ǛH��H�����D)��~����c��o\L�Y�h
�6�3G	���إ9�f���3,��ԕI�OtL�� ϫ������(��	�aR�^�B�}4�K�]S�ӻ�K�+�Җv�u�-����<��߷ 0����(7�1W��(	%*D'6��m�č�p����t�v�ߚ߭ǃ���E���c�-�3m���Cߣv�Q�&d��>7�$����3�p�_|��[��3���������I[iOj?;���Wo�]�`���$�}j����)MJղ�S�0:���~�)B@Bƅw��J�ݩ��Ԟ�{`�e>Z�aԔО��7;. �o�K��������x��Bm��bϿ�+�|�	7���~,��~;�����L<�i�1�b.�ww%�Q5�O�w��6��_5vo�c�[�8S�I�\{z�#2uQ���-��m�*{Y���e�ghk�홊�j����1�L�Й[k|kۣ��D�W�[���r��7O�K-�������{E螟uq��GvY�o��m�u��hdVe�N���#����G1�<��zM��z��@"�Je7}&Wӌ��7��s�޳6��*��|q) ϧ���%]�>g�Vu��MW�n��A'��=g�3
'ĂR\�(*��o�̨P�U8Ĕ֐��o��G!�f��y�_(�|,���ۭ���#�ٜ�e�+�as]�d�c8n�p�Ae#�M%�W��rz�3)�Ɨ�td���(��Hyyq.lPoj��z��B�WA���IGX�2�.�6�J-|[��l�t��U��k�S}�5���N���'�\ela��*؁��ܹy'L֗}+W��\ۗ�$i>{�pe�E���<�R��63t��h�f�T\�s���Q�;�E��{�T�����JSVP�W��9��X_;hs�:�MV<4���{ozMU��c�݇"�ݺ�4SE�雦�d�:���ntk�S0d�:��b�h�H9��y+:�C	Ci����[#T��x�SB�Z�ۺ���]�����/6Rt��sr�ˣ�L��K�49�	r�iX�Wj��~�p(�ף��n�*�lG�E����fN������R��M�J�ٗM�}	M�R�N���ߓ#1�:o%R�����ݪi��=|۫������n��-��\](�mN#du����.�+�P���ǝ�e��)W.ł�׻t��'u��n���r0ݤ�J�܏�6�l��tG!�I�ǂ���Ll�5m��+L�*mM���WM%]��2�xf�۪�N��fZYGD1��\)�}M�����C�t�y�^�Ce��k��,p��+���/��|S���N�x�t�:���sh+�s��{�[�����9�'b8f�u��87������e��t��t��L̷c
|S���F%5��U��R�dѹå�Z�5�C'N����])��mt���Hf�����-�.^�{��[�u��I�z�YƜ]�&�@�q��wv�Q˰�ZF���}X��%AsJ��V`.�q��4��ޙVo��
M�[j�l���Ur>�+N��m����1�5X�������{�(�dZ�����<'.�P��X���ҐT|R��L���]L�=�Ąu��:��g+�7�\���m,���竃�^Gj�w��}�����/�]{Q۾����oJ���k^ѝ���#t(ɣ[Ew�����JU>*qS��+�%��t�ZZZ��dň���C/P�<Z���J	Q�ȷ����9 ��GEWԎчQ��j�x<K&���{�\/Q��Ί��$�yc^.�pJv#�eM�n`�Xl��߮�/wU���Pͤ���i��zn�уm�W1ܔ���'��
{:����D�����n�zo�Mo׺i���s;�o�N���ǩ�d����c��y!����EI1�^2����]U�a�-,�Wr��G.;����$F�]��]D����.��	�jGn�+�L���$]��C��ú5�o�¹�h��qN,�/{f[�3`�o�	��U�ڲ>�c���)G��{�m�c��=1��M�'�br掰���T*j��f���+tE��}��;r�V5N3]ֻZÙ�_I��@�WM&gt����������tL(���{�uN��N�)n;���)�^�E�M��D���-G�Q��V�G-�M�B������e=��1ze�kK����Χ��0�cw�rgR��Z� �q�I,�Q�u��� ���`�;��n�3,	���j$d�z{k�����ֵ�k_�חw����i��$čA$���C}�?_m�iA�dH{9zu�����kZֵ�|~���߻���{ޯD�d��3"!��S$HFF0������������kZֵ������/.��q�8&���MFY!4��u�L~뮂A�m��4 �/NC?WH��ܒ�����1Lf�,iF�ݸR�/}��`"���^5�N�D�$'wD�& ��2B�%2d�6"I
�̄�Tc)�"o;n�	F��I�FY"2�����40=�]Ѿu��]"����ݹϥ̟uK���]��z^A�$�>���,BQu��$d���N̆h�X=}���]������y��u�Z78T���8�/��0g�>���U��œ;:J�c��[�X�[�p.�����2��� � ��:��證��;߽㊕��)������t�5�jq�F=s��Q�Bɰ�VA�7��d�\8Fc��4�FΑ�b�X�ۻ!U�,�P0)�=3������4R�l�k���]���e�:"��⁓�|-�2��S*��ѳ��{[e)��vK�N�>��l��F�U%g�/�8w2��#D�;�p�|���2"1Hggcz�w%U��Vc:ӵ��ٱ�'iuN/`�g��
>�L�����eх}z�	=4�I΄P����+�����6�=�����.�1��I��^�2�W5J�^@7�+��JH+�˗�,2@�m@���H]ӓP�g��m���<8��UB«?]�>�n2	��+��Mݪ�({��/��s�����(���C�#}^ƺ瑺L�D{O6z��C��E��[;�e�������>����f;��W��ܧ]];"T�O"��L-=N>ǜE�G���͋�2eyz⻋�f+<������dM��c�:��+����{�lk���nK3�)5�[3j6��[j	�i��c�>չ�ݔ?��^>>>>>�fm����zL��̽�,ϥ0k�{�"&�j����2yK��!���&;_3����X;�#ײdr���zBT�S���T��;�ߔ��J_�8�Qn\���e�É���Q�6h��i��SÚ��
zÿ��w,��4f�X�̦��v�"��W��,��<�p�gfqo#��6��W�u�$"p�S�>���.�<�qx�a�V�%�;�+�tQrg�%��h0�6�F��S�fi���@�H ^���+�fB]z䷣ʐ��#ɮo�7�|o7����c�2]��W���!d:�������o&)����͟�]7���r"L��b��}!�/5HA=p[л���D�,6s��ۀY��3�����#6�xϻ��tF7���O���S��\>j�w=�^X���o#g�χV��i^E�i~	nɽ������ހã��Jݛ/��:\s	�sXk��:[�Mm\���n����UWA̹C�Ǥ<׭���Q��أǦ"굡h�%6�*���L2k��0���R
蟴߯��Þ�gpo+�Pr��r�Q܂sT��ۼ��,8�n�b��[�w�;�3�q�D0�ذ�' B	E��a-�cD"|��i��/������ک~oԅ�]��v����s���Y��u+���f��cj�C�M�5��]�v����C:nG����roS{N��f
���H�Uk0l6B!��Ec��T��C�5 t0���
 |�oL,�H�z`�H9ED����[��+��y�f�����ߞl5��G�Ǖf��Fm�|��Lͬ�N4qn�m�U;ݝ:���H� tTk���pt+���SSԂ�񼋛{�|�4�V�Xâ����y�{�gR�����gA
�&a�l�T����ݲ?LM���u�g����/(>��9��͕���8:5FW�!��y������=��3a�@��T1p5@v��,�%�v�d�ŮLȻ0��=ϥy�k�m��	%�EU~��
�vM�s�ה���A��w��H�I�ӝk�(�ؘM*Fo���^�n�&��t��4��fU�"��bah�4�����?gIw$�l.����b�Ŝn
g�u�^�[
e��R�#���������GtA�V��~vM��~��>�پ쨝�۹�#f��FQ�Y/N����Ky�-�>P�}5K��������8e� J��r4����߾��¼�7�o 6����%�un~�$��~�t�u������]X��pF��e��g�f����6t&�yxg��R�v����@5�8AC���&kqQBp�=m�{U�	�$��Q�oU-X����WL�/��V���;K.�����a�L�0b�1���L�.��F'�wM���Ț��""��gb�c�>�ar¾������u�,%Hs;��p(��KК�ݝ��֒cz&e_�g���ˁ�=��偕�t�C��6�����Q% y��M��O`8�N����5���HYuoM�Sa��ʆ=54����ӮG:��hz�3���t#����9�s�����Z0�}{�)�ǋw��?X�z����O�sd���I�|���gv5%�O��R�!�;U�UU@	�n~����Ϸ�k������];��sn]b���-W쭟E�H�;M��\��w��f��Mr���⢒hѩ�˒)w��.���ѥ=Rfxz�um
#�	�<��_���w����K=Q��7�������r�^���޼�Uy�Q�J�k��(TU�٢b
���S������o7��=���1�Jn�$P��p�?�^l�"����o�.��54�޺7k[Ӓ�Wٰw�4�z�ϲY�a?�|�sab2*���^#�E0��ɪ��6:��/���{r��맇U��A]X����d,�t��,!�sσE��n�����$ah��W�u�r0����ٙ��'7"�4��&]7�j�˹���W^.&^(!Ӱ�ݴhMx���
J�>��v�F�����1����g�΢����#Y�{	���kn��oSu�p�w�:�_=����f��!�6�AL�Jܾ����@ba!o>���XWy����m�o���TQ.GtA��ك;jf���aJe���%�㭶&r����i�k�}�>íot���L�;;��6���K���;%����=4i���^����GS]>��. ���8~�ǖ�Y(�{6�"���ӕ+-�>T��R�q�����Q�2Ft�y�����v�ո�-WKܨ����P$�u�g9+*���Aa�Z�÷�j�+��m^����?!�^x��uJB[�sB�^��r�'he���UO���������h�7�?>p
}�NQ=�^�5��M��4���o�p��P�u��_�zr[,��陛`l�I� u���&���<t�Hc}K �V�q�g<�g=k6q=`7����E��)�YD�����2L��_�x�]9샮��]A0e�w4�v��z=����摠�a��;��>-�S���g�p[X��d�w:�Ҷ�������zE⢽UH�x��쭴���3�ޥ�[q�1�j�^�T	��5
�C=BT�S��<d�me�W�/܎1���ׯw���w���Ѹ�:Z�Rwf`����-є�t�x���$�>O=��%�ofhUC��
�M� �\��xi�t��U�
�:�5�G#�)��]��X+˯�"x��T�>�ц�o��U������ǳ\�4�"����JEi��\�,��).�:��FM��B�Roݶ0�.@�:U����Wf%Rqvf�$U)��SF�x�"�z7����X��f�I��0�ɷA�JdJ'�Z�(C�h����!�z�u�׎���&^��;�F5�.�k,�Ng6vU���̻O��l)�+w�8������=~KBl�Lq�("	�7⢅��p��)�",%>���������l��_Գ�׻V�eWG��o���a�˕����=�Y��i]׻<���ȴ��NK6h1�ћ-��www��w�|z��^iq	�;�*~��f��C7\M׌�c�{������J��wQ���=�T]����;I��u��q�)� �uYCV�%����򱋱����̩�5G����uu��X�'O�K�0��ϧ�c{�,�˺�,Xd��W[��T��\�&o������+��O�
��Tޭ��WG�����_.�7!��p�Y����n�	��.�����U��%�R<�w��;k�e{����	y�V�·g�0EzDLQ�����b��ߚ����
_��n�_�o�i$h��|�[�� ���Q���氃�WC��m�v�J*r���8'��ԭUGO��r��`�uH�a�\����C������>�����׶éa�A���,,�j���z���5fS{�Kf�DM/:����Qal�yW}9"�[����휭�o0��8���nܾ�δ�R���朓Jg(Q:)pr���(fbw�^���������o7�{�0 �9�P�eYv˘���*j��<z|}qU�Lk�U2SW32R6�-��6EY��&�}��Uԕyd)�5�3V�<{��D���B�~uG��ϝ�QI����Ka�%�9��#:&u�x��;k��U z����S@ H�m�,�4P�γ���{��x�m6+����mq�#�(�Xr�H�p� ~1��t������0�Ӝ'6	��oI)P�).�����Pگ?|>{�{��wq�����w��>LKCL�ao�}+W{_r�������K�.ෟd��m��5F4��y��I�A0�7=1O��dn)��s�6�I9�i��wm%7u3R���]l�e�3o��9�w�~�P���;��G�����́�u��P��^CjW��V�y;�: #L8(|��szL�afXx�^VnNf�>*q����%G<�:�N��P�ffm!�#���-��i^�V�V�D����/�y��-;�a�v�Hnm��l������Ո9T�n�Ӹ��y����#�s7�Tv�Ń\�x���\E��+s���zx�|||G��8��x��CuO��Hk�m��;E�ӪM����Xn24g��c>��F����Z�9�ɣ�*�<&��C��/�9,��t�k��-��绶.��Jl�t@,`qm�%�=��2+F/]�;k�5��<�����"�q����8�����W}��i#��ە��H����L�a�e�$N����0@����E�ڧ.}q�L���*O�[wByv�y�}"j2.#S����m7l5b�1�uAa��%t�XCM[�N˲�\���c�$���ަ�:ޟ=ň��jd�v6o"��d�W{$j���B��%F�vUΛy��
cODD���Oov6�ޓԒ�&��}��2��JR
[T���^�o.��ͤ��� 7oc5��\4��3π߫VH��t�ҹy�R��=|�?�A|wɳ4��5�E'��=��y�J�4ncMGTk�,�L���ׂ����gi�%͓u�[Z�'���ui��$�
�>'aI$�ɃMk�@�����]�7q���Vؑ�ڭ��=U�.�����
݆�v�)�����l���u��{|@>>>���nr;��v���;�ha�f�ĭ��ܸ��Y)�i�	�#{��C�q����髕<5�R �]>��+�v�m,_U����쫡C۾���<�I}��ID�b->��j�=�j� )��`���LS��>ط�Tuĝ�]���M*f�Ny��#g��vغ�f�k'a�f���_1'�6[�Ms�yyu�Ou��ɽ��l`�6{|�A�f~ko�
z��;O���$8�'�m���XQ�'$q�:c�!�[A�U�G+�	�B[��w�A9�H��[BR,[�#<�7F����5;-��9��ۚ��
��v^�C��Hy�j���y�n�P�\ɧn���Ӑ]��oZ]9�p��(�Z�x�����f+����z�a=�d��D�z���x�
�KUE~��}ߏ+����pW4�c�_�@����# ���4� P`so���Vo}��kfK-T�e���[55Yc5�Եe��MMk55iV2֙��jjkSSkMJ�ԭMM�jZ�Rښ���2�T�֦��jkSR�5+SSZ�����MMjmf�55SSmMKT��u�jkSRښ���U55�����j����ڦ��55��������MMT��TԶ���jkSRښ���ڦ��jZ���6�ښ����MMjjV���5-���MJ�Զ��[SSmMMjj[SSZ����֦��56��V�Y����ԫMJ��զ��jm���MKjjV��kSRښ����MMjjV��jjU���5%��xE8"�@!&��5*�R�5-��Z"P�0@�U�b
&�ִ�*��e�%�u��U-Kj�jU����T����� A("�jV�KSZ�Z�j�jU����T�+UKSk n�!��B �A�-Mj�jV�KR��Z��RԶ���Z�jU�����j��Z�VK5j������mT�5����TA�" ���l5+R�eZV,�KR֖��-J��2ڙ�[SR�MMZ�K,�jYL�i���c+i���MZeLf՘������k^Zc6�c�f�����,f�5-Y���[56�c�X	�w22Z��2e�6��SUL�ml��k5-lԶ�m�b�j������J����ǭj�H��F��'��3�����_��y������������������@����?Jf?������I�?X� ��O�??��F����Ċ�����~�� 1��O�������~�@W��vx{����ԋ���N����O8>�>��&~'�pQ�D"b!"	"!�� �f�6Z��V���M�*kS-SKj5�6����2�%j�U���kU !�$Q"���*��ڪ-Z�VحL���%ZKT��)�M��Rڛ-RʴԵKMZVkSij�M�,ڥ����Z�5���T��J��m5�(�B+�)#*�U-Sk5����֖��J���jV�T��Ե@B(�B"��?@B`����i�O���(����)  $���@����������>��4�w��@@\ׁ���N?���q����H}@��!O��i��?*��ʇޟo�>��qD U� bR? ����*
"���v� h7�L���:�����p|�G׀�8�@V|�����C�~n?2� ��
�������>��?g�}�ǔ>�������C�A�� ���)��� 
�@8�8>ސ�$Oμ}ɇ�	��~��}�A��=O<��NU ^S�#��~t���wC�;__����E�����QAD]���o�/�}��~t���
�2��4�5������9�>� ���UR�T�IQU*�UTD"B�BR
��T�J$�(�R���PDR��HI")$R�$*�)U
�HR�������=�B�"�����
)D�BGcD
�Q"R"�V�DZ1H�E"�%UEEQT�*�%+�!�EIB�!��R$T!*�%Q	EAJ���*�)U J
�H�%IT)$�@�@�
�UPTUR��BT�P/�  ,U�����nTun�iv�[U��'k�m�K�eWB����jl�֮؊���+�\�J�I�����j���5�u�ݱ������Ws��;�Ԗ��J%EHUD��  ��ȑ�hPȡ"����lP�Хhhw��:�

۴���s��6�ѹWWWn�\�I��K��kW��J���ݫ*iew6��v�l\��9ws���]��$�TIJ**�^   #��m���]�;���sU�@;�m̫�ka���ݴ�����l�MCl��]Ym�2�WA�e�n�ըn�M����Wk��l�Uv�:L�MtU�UR��$*J�e	�  ^篛m�j���ո�����6��U\e2�XݷP2�[mu�gm�V�jؤ�B���تٍ�.n���w+RR���#cJJ"JB��  1�zеC�L�b�ړ��ҩ�W]UV���c��kv� ��2�Ԧ�9t��X9��e���M�U�*m:��v�K�$	 
J�� ^�EE��\r�u��Z�t�j�wgt�"S�V�kfګ�E�&7U��G:���6)�;��0`\`㚫���VۡӠwRUR�Q"*E$R�� g� 
��q`��]�0t�L���� :S:�P�(rX
n܎�V �-�9�(r7(  �R���@J"��I�  �4 �}�<h@nˎ�Ag+�:
-�i0   l
 7T� �SE���wn�䶎�   V*	H�T�%�$��  ����	n��Ӡ�, +��֜  �ʶ�w`n�C���( uV=�� �5t2n�p��"�OY
!BJ�U*��  �t:h�J@\L t���� :6����N�p R�N��@�7@�7$� Kq8   �~BfJ�(���$��@ h ����4ʪ��I�mF O��*   �MT�S�� ��)6UTڀ O���/�=�އ�?-���qu>-�dE�3n�����s곰6	6�ȟ�x{�����u�C���ֵ����Um��mmk[o��mk[o���ֶ�mUV���������w���鉻k4���^�)�1ZJ��-cr��3Q��Sj�Nm곺&T ����a�g�.����l'��Y���F��Cv�6�Z1ٓD�*��\G@�k��OkU�WE�a�*ӱb6-��DK6����z)�*;��צi��S�����lOj��AL/���C
O[�chnfX�(�)/��-��!`��^$i,��o�Vo-3u��J�a�X7]e^�aU���P^h��n�ɫwuc�PHڭs~	�����E-,��U�ed�e�64�2��h#�a��M��8���R]��9w)����$�NH��w)BƌY��k��"�����z^�VX�p��^&�Vp�輹v>Y"�>���,�k�NR���$���ۻ�ڼ-V`��sw�]�rPHY5��y�S/T��5�
1J64hg#x�@�s�*���`���#�Հ),:�	�r� �Ux��6Ld�>���f�%��I8so.=SÐ�:���B\�ۛl��0h�Ҝ�aْ�����"�D�حci��۹ylCx�t(͡����F ��{�!�ך��bT�v�G��{0L��E�W4�:�`'q,[H�P+�+�2VPf4eH&=�B��l�ctrٻ�(3s�ӕ�UƳ4=�1�h֊p)��v���GO%@��w��s5&��ʵZ[5��r�m��x�t�X��'�j$��6��;qdK و1���SQ��baif�jA�n�^"�4Z��k׳TT"�hcVhV[CM������m���g,����Ǒ��v�6���*΀�E��P�ys��^֊`�(MZE�b8+/J��*�3S���F[�/7�ge��k�S���E��Z����fZ)� �<ݛz�D�(��٩3�%���qj�����ZQd�͖-�nK�$E�C{�Ǻ�07B���W�Y�1&$ͪ�`T�M�R��ű����ɹF(��ͺ@��־q�dXj�%wU�l������x��eH�Q������3ڊGQ;-V�a(d�@F֐f؊�6��c�ސU��g"-�O/e����$fL�a�)�,7���H҂����;�ҩ`�!��u%�[�Z ]T�Zr����lnA��Mقd�L��X�|%�6j̣�n̈,���� ��L�
.�`B���3,�3�r̶Z��6���_3uy3T�q;������\��DU�eЖ�[�oo`r1�@mn�ę�,�[�\N�y-h$Z�4�j\׷�wV�M`cl(-��t��0jaD���7��lJn0kH6�%O�=t*F���[�VbcSצ�(h�d��B򂛛�I��ڹD �,� ���'RlWj�A32��]�Ս�x[uv��v5���%�lh���;�5��hSa-�@����]
���yZ,���x6�k3�F�c¨�h����r�\i5v�l'Q�2��r^b�u�ۙ)ٹ��.�V82���9+,f෥�ܓF�,M��R���R�ܽ���R&K��7hӂ�)j�K���$>�JW(Z��J�|�3t��[Jׂͭmrm!��{(��v���X�ћR�w`���!N�0nwbOb��M�n�i�Oqm��
7���0�C�Z�0���i���K�pyR�)D^jŤ��ʼ���D
ה&��#�/ ���OV��4tڲ�[ �	��[t�bJi�ŏ6�LheǦ�1V�1�x�n�kc(�d(K6A�n��n�B��vv�&���t km+O���w��� <�r��a��0�C+k&�bl�S�,�XۧK]f���^��i(+A�#ی�$�z�C�V	�3B�Ŧ�Qc���xu4%��YV	P' ב[6&5�n4�w� �ٵ/d�H��j���4ŗ%��2��6t�(君��j���-(�[^ɐ=���$se)A��sf�פօre���]m���v4�I9�a���hQ�n��.��^hc.i�*�n�4�⽙l�i����3b黄3�ڷn�P	R�5�*�p�6u�<�� �u�ܘ�áM7ôuZ4R7R�ƕ���7��1���6��0^�QJ�sha�PXV����;%GE
���[(��R5#E�\�Ÿ^�k&���n�;ܩ���uzΗV�;b���R�fuv�k]�u%�bjlm]hza�� �k�ة*`�4S�J�;��".`�Z�n�;�4�����ocݒ��Y��6L���&�d���`"�g��4�s$��7\FL�/,ք��\�\Q�&<�;E���T+Dõ�l�";����x�b�X��ה����®�1-�&Uv��]��e3,^-;1,[+Xx�%ii��]��6
V�
�Ȳ��#+�b�(5XɃ]�x.�ڎ��Ej�7/�j�:�	��p�k̉%�o
�@J5�=9U9F�F��Q�MJm	P%J³Nh�^���4�rKʳ��c�Ӹe�/��t�]�2��b��+u[z���h�6�V�C�f˩X0��y�����e! ܢ1�Rm��TY���CH[WX[Dj�Y��a������Ub�;ݸ��9{d�IJ�d���tc+kDu���z����W��ɓU�^Cx6m	�"[3>r���Z�ś�@�R*Zb�Ji�.Im��kS��`%�8��mGw�,:� 7.�]�mT0g�7cS9QDۊM`;wQ�[��ˇ@v� ���Yq K��@U��t���)�գb7���������!;6�Ƭj"���`2�=%�U���;�ǔ�"2�V�V��[Pa��B��a�F�X@�On�� )g��)��V�(^ۗ�ݖ1fX7�U�u!T��G1�b풃ۭ��XV=m�7�@�哎��h<��� U^Kt)٬�Q�cVX�-Men�� l<Cc��3ڊ�Y��,�Cr_�7�����HͶ��e
�(�mԠ��*_�6�"F⛻ݫ������̎Tޠ�ll�BP�nw����g8�Kݫ�qX朧M�3	�f+Z��b˗F'�tS��2�h�reL�{J�+n,c�U�wt�t嚖�8�r�V���,�h�S�lil���qɣ�aj����kW�8��^7RPdڊ�`z Ц�د-�[;��KYY,�Q�9oH�CwtV�B�� "+t���3ab���wZΠ�$�@�~���J��9���u��Xڇm�X��iݨd.��r����Y��i��I�K�.4�e�G���UuO/AU��\ܴ�XP+vj,�D����N��l����CU�,���d�`��+C����Id�wfBE��%���V�@F�Z򞰬=�L)A*�3��Zn�ҵ��uVV��̩��,�m^��a���Ȕ��"��� �P�i�f!�ԫ�t[Y�Ib7 �j�Y@QŪ�G[4kt%n
mD�{aj]]��q5�Y���j\tRϥ+5�[��fUʊ�ul�%1���C��;7GJ�k'��#v����b�l��I-i����Z��$��NbyvZԅ���U�3Y2��N�Эz7Z�R�����O6 ��ߕ�R�km9�0SB����q���ˮ��˗(�h��6윚���,��wB�\�����(�+i;$�m��,v6�����vY*�ia���wF�[�e ۨ
�
�̬YH��U�ݽ1Jb��Y�ٵV��k�� \Wwpb���Z�(X��O98)p��v��7Pn�9���[ugTQU���P`<YB��56�J��"a��Q���̹OZ�2;t�BT�C4�P�7u+1Lʔsi��b�m�ɛ*ƽlE�$v���[ZD˖[M��B�p=�O��T�ܫ��Fg�:[�J�8����:,���L%7�1I��m�d�I����^z��Kg�V0Ȗ��Y�^��U�YwF���+h�N�m)���%�$�VC�],���ї�VG `�YP�b�T5��(�v�F+tR�K�HX�Pښ rf�dl�j���{�����u���m��Z�j�駻3����E�BC�1P�j����+���MnT��Ѳ�b����f-T���TM���|�lՖs6=�)M���^���4�İ4�Jc)��	J�]�K]�)"f���E�E�KXYt.Da)�q��d݀�z���-���iZ�������%%�n�F��y	IkCVݗV%���/1�xH��Yt���&��p֐	J��p��"7���Nc0l9J]�R'��b$�[�7{a+�#i�ʶ:�6��2�ZMh��	��K1$f�$��R�Y2K��ik��Ln��9S*&ZYHݹ�ᡃ%�32l�'�gjd����j��l�#c`��8���r��N�۬ORoFܭ�10���w��-R�_�d�"%YR�]�@�L���J�&\�GT��;�n�Te��*�lF�,Q�lZ�)0"���&΢�
]f�oj�B��܂錄�t&R���U)"�����0�0�'5f4Q�F��56��٨j��
��HAV:�ȅE��f�N�U�{���jbVv���da�q�ڼV���7�hf�U�V�2���-{�%$8��:��ՠ-܀浙hEr�Ӂҏl��X��V��̻�p�u5*YoFR�2Cy�Bq���i�aW��̷���{�%
�ي�,�%���HU�Hm�a:kf;�6B������WJ
��m���頵��^��P6�@P����ӳf�[p|��o8���ثI!��T��Q]��J�=M�� 7ʂ�ia`�����;��Dk.�'V�5���Z�Z�J�Q/n��*����A��F�{{����i���%E�*���ŵni�kh���VkE�qU�v��+c	4B̈́Y�5hܸ���e�O	��`�W�f	`���YǧF+ȴ���JU�^�����Jc+H�	�Yk4ٶ��YMFq���6��̸��=4p�5=�5�,j6�XH�81���X{KpСJI�����We��ʭ������Q9���AZlҪj��l���5�riVkoF5��cEb�1��Jّg��ٺdYa��Kj5+I�2��&U��~�ۧJ�wbm�Dl[��j4��ف@�FF�+��B�!hE��)�	m� y��K�{���˛�]�&]�6(�V��'Ko6fޕN��3�+f��Ie�XEc��M-E�L$��X��Ei�-�Fͬ)��nC�;��U5���^(����[8�+����`��NT���6����ct�7j��/i=jJVT�k#���ɤ*v��9�� Q��̆���O�Z���Z)5�(ŧF�D2��ec���fk�
��^��%Dސ����r�	o,k�����L����4n*9ha��R����,��Zã���0Ju�n���ehR�+��1��ଗ�ցwR� XT��j:͒@۬�q�!yYWb���!��P9��k)�Z=�wi]�kCG2�R��`&n�/fe]��<ݦ��mۦ�Ol�š@����qLF�O�u�j̺��`�%J,k�E��dC�Q�Jl̙VA��ob6��0�]0����D��G �b�/s3v�%��bkU���t����-���i�Aԙ 5;&�F� �J{�~vL�{.��*R�3ku�������re�mmj�;N&pùm�x��9�-�«WZ��cu� ^=m�4^��	v��Ƿ��˶([ �Z!+_X��� �ٚw��8Mi
�-�jL�w�ykmسxȵ��sn"����šг�X�2S�'{d1C@˰���@�f�d��iE�D˿�,!�l�Θ�@N�4����.��^f�MF�I �W[r�C�]�[gK�ɴ��Wcr��D&v[o+	�*�V闀1��	-����[tb�35LtV7�f�R��f�KHɆ���<M_�M�p�/oY	]n��F�Y@;��ے�̨�5th��<!1��,�"BM
m�(B3&�<�B�`n
"����L`ҳr�̀�ͭ܂�l����7w ua��/��;�Z����(����˓d�"&���k��
��^<Xr���)�D�P,K�I�<mX�a-藙#�Bf�3p���6�f�i�Y�Z�"���Pc�M��H�N�*�����R�6�%hT�:�c��YI�b'�Q��]�f���Y��à�*�hV�B�5��I׈R�oʷ�����vV�ne���
��۽l�XҨ�U�����I7��S~��$@��=!� Qxi&��nf���(sfY�.f�mPS�h��Z��`KW5	��I�1k)2�f��v��+,��V�^�ۅ�
���{Hm;v�؞(�%D;�l�mꗒ�M]+�0�q]���	�ǵz̄nɶw�lYɗY�kc̬U��^�^��j�h2`�!�E����{[�1�en�㠯K̥) ���G-օC!ځ]<��5���1X���0+��F����5�l�݀E
,?�*��E�wu"<�m���,���ǎh.�*� J(��J�jS�x7-�{u����z��J�97qظdF���`#�s:J��^
�K@��VM"���%��@
�\;.��5�s#�F�b�
�z-� �e��{hFs
6X՗��`F�ר�6��,�.b�%Nk.�?K��ֹ:�X�s��[r0�T�Lt.`��^ѩ�7����iKlcQ�M*ٮ �VuZ7f�9���kX�#uhn�S��֒t�����1U0D�%���AR,(�yNS�K������T�J��$5vrٷ�6� r�m8���J�:vi�m�iZ��xCh�ꚦb��n����ϣ;@<����w�Y	�%�%fi�e!j�Ȝ�Tc�*V�t��%�bt�v�:S�6�պ����}q��G�d���k_t�R�w�wW �Q>��-�e˭)��<\u]�Bp�� �q|��uzh.�kP��
�ԣ����Wa��{����tC�d��'=P.eYHq��9e��ۍ�6�fTg�6N�Wme>����k>� ��˩ŋ�[8k=T6r�哈�;1[}`l�,�3��bS���ڮ�b
�uV����o���jz��@�����7�a�5J����-�/U�+:�==��� �Cೲm&��S��Q0�@��g�]�� �f�^,[}��mpߏ}V��<T3�^�\����`�vn����˖������S��+`�'�e���w�R���%2"��A�k��#�}ӫ�Qҗ��eK�˝]s�e�Sn����N��aH�R�����zb�z/�:w��8�������<��*R�j�U����OSn���Q�Q�w��ov%����Vx�\�e���Shu��*٘�i�p��g��WRR��V�)5@��hg_n�5����,�������Y*Ax]���5|��� �A�t�ln.]���{J�l��)�K�O�ɤ���S�x��)G}�JRú��KBS��8����\Fin�sۏ-�RH�"=B�r-��'79rY;AԬ��J���o�;�^�R�]-�	�W{ؾ�d�⛚(�fub�*��+�u�6�陱gp����p�Q8U��mX�ծ����t�f�p�LPVց4<�oB���c,���xZ/�Zd����x,�i��'�u�J�VU���X��aqec9�7�ɺ;��\�ɮ\�\�޵S��=�Ʃ͵v�|���۽V)H�0���C;u��NX9oUo1��;,+������Le�i��%���e�ً:9���*<ч�.B������r�ľ�Ћ���G#%���az�6��"[���D�m,�;uj�n� �v��!A����G|hP���7�*e�Ǹ��}�r�;�9�1]G[A�� �� 5��]V��ư��Z�֣D�B�J�9����ƙJ�^��VZ�0]=��#6�z���o�J�D����Ǉ�q+jb��Z��N��Gv���`�|�״�۾K��ݲ`��Ũ��K�wyb�=�/�������<ui���n�w�:3��c�R����姳Vr�*��Y˷��-tIe-3Fg��'(�v�LY-���MjR����e2��/�\���'y��9�PwץJ��}J�Y�v2+�j;���Y�貨:�VfSUsc�{Ն*86�۸4*�襗�u��4x4_o.�n�\Z��}�m�)A�vw4齸LfY�f��՚w�f�ҁ��AV�IU�����DJM��@0+K�6�]i��o���g$�h<;-�Rv$�w̘$�BhW�Q*�K���0g
�׀s��ka��5�=f�i斧NH�V���z��Os̔8�Ԃ��}�,_b�t�f�K��+Tg�V��9���V�ҰL�񵛄,(�$(m������.���{0�k1l%gTƏ-��eYQ�r5+{wJ������J��mJR��y��
��8Lޢ�x3�o��,��5�p[�K��b�*6L��M$���$^�"M��r�:��r�d��O�+�S��g���,9!;�)����_kҷb��"�BΧ��b7�mY�]�*`qأ�ڀ��X��qVG�P�h�����|O^����a��
įc��ΗҖr��vU����bיX�k>��P9�zT��ke����@�JP��tθ]�Gٸ��:Շ/+E*�wW�u�M��v_r"<v�<����i���fÄ��'c;��^�3����̺�k����I�����ɴQ|����C;y3|���y����%�{Kö�
=W�G�J�7x	xp��O+���GP!�b��4s��_V�K���onl�������B�%�nr��j��r�p�,��eR�[�j�	��N�r��ֽ䈾�Z��n�;a���2�v�&� ;��bOI��8�����wep�j��G7]q89cZ1'
Iu�9��j)u�ՕɅw���sw��]hVbe]�]|.k�ܻ��(k+eB���ڱ�S��/w-l�_nǬ�IV��8��3��.��(|��&����Bp��J�n�R��F��3]Bnr�l�@��*���b�zt��5Z����:T�ܩ���%o;z�m��G�me�+F8ºt�W��(B��GmYȎ�V����,��E����u;����.���}�c�:#��u�DvV=O= ���U��l�(����;Mt��`�t��*NV�3�k�e�:����Z��y�ƻ5ܬ��"�_Z��]��o5f��̴rpw�ߕ³��f�t��J�	3%JB�i��,V���:|�4�ZC��^�7}��p���p��m����[��������2����+l�2��w@dߌ��$Wr��V�K�;w[y��>�h[Y�K���j��]�4﯂tT��Qn&s.������㦳7H��/��K3WZ��k�.�Q�G5��H2�&�\}�Jx�����X�TkWv5n�)+�)��ň���4jܵ����hP�6Y}��{p�B;�7s����W�Gz6Y!x��(q]�=i#|+7����v�Һp�}��@�T�G�G�ۺinʐ
����3���4|'N0J9zjla��W7!{��c�{ץm?����T"^j���W�X��i�[��*����*iV�|��۪0e�@�_TȤ��Y�$ڟ,ٿ:v�NinL�C�|)wT���x�lI�����ߝ��r߶V(��5�%3�7N����͐ B�ExŢF�:d'�����Ů��<��m^)�u
�QbYSc�G�����2��GzF0�oe>�^����pJ��wȷ}�b� Ŏy'U�9��e�"����P���o@�\�M��f���kl�Iթ�[r�������W�}�:]�W�{�����#��P�*��V��ٹ��dWǞћ|x]�[;��sA��VsE��<�>2j��W��Nu�Teb=0Xx��W��μ�0f'o�/,���[}��:�4�'�-X��ɫ;)Q�7��J䌍�U�j��Bk����d�fV��⠻6v1�\Q�:�AXU��ݘ��E��e�i��Ts�!j��9�V��1U��lv���[��,���)
T���B�ܝ΍ƃw���Շ����D"1@��v����˳���].��-tr�����u�'�!��-vպLph��H�6M�S��{|K�(�*�d�ά�lvlH8}}.W>��n+v��e�J�;㩻v�"cUc�T����J�`�R����G��仕Ҥ�4�1�|��\�*J�N�����,�xaXmحk�[Jme�M��ze7� Wq:�}��\�v��4�Я\����v���>��A�H^v.��vt�N���y:MwB�գ����pAƳ�r} �1�ur�1�2�9�1�%t� ���G����<h���^��^�mm�T���Z*&��ə�f[�����J�`hU��}|�7W��(��t�-���Ӕ� ����pv�	�1N�Q�j�*U�r���}w	"�ï7�f�W7���]�Ѐо�*,�QLK�V�	Jқy��6�a}��WG(��%kEv��/C��F�QX��Me�-ս�	��E,��>k8���XL�ʲn�����k;;(�ډ΋��o]��WA,��5p�CY�+V;z�>��vv�� v��1+#�����<Z�$�i��!{�GB4�����5a��0�B�l�|��+�jaͽʒ�(6�A��me]l��
8[��`8�G�<�T�u��,�We,�C���@����|��c���v���_�Z��2�E��A��-�8� ɛ���! �-��\�i9�{;\��ңgj�6Ṛw�Ÿ��������i�ˆ,YKb�`��w�z�G��w�N��+��dt�֥\���oƅ���N
e:�l>�+9�gQ;BFW:y�|���w�m�z.r��4�=u͋U�#�@�9}���Oy���u�+���ܬz��vg�b�N[% ���əYYSF�yc
t����'���!J⬱��Lw-]���g"ݠ�a���i��X֣�^��&�\Ш��b}�+&�g���VS#dG9�w�/7Ua��Ղ�9V�<{L}�uΤx�N��]i����eeY�C��!�!�rڽ�"͈^sXs���dި�KN�X�/��6�J͝Dp3)�-���u��8��	Uu�yݳj}z$Cݍ�Ԯ�)�Ȃ�쫆��ø��X�ԣq��E��[�8%Wϊ�W�]�Q�x��(>�����L����/Y����6p���2���i�r�S�"�x8��*\[�����c4��]��N`gd(�q�5�:C������咠�f1�	iX�1�ʣ�ae��3+75*}�:����;KSZ��j���8]Y@n��_6�d���:����tR	��iTν��|�-7]�\�q`?p��;�Z�x#���Z����I]7�h�b������>�[�����q�R���r���rl����&�u�M��R�#t7m��{�-��kz��Oi񃝺����-�Id6�e����K�th��o\��E��cc�w1%F��䭫F�Sh���<�&�,	׾;��Y��N��z�:��R�f����:�����W����e�!X:��K�Ҝ�+�wJ��f_r�Yxչۑ<�]-*�c) ý�W%��;ќ/i<N���V6��W]���:�Z�8�Y�����|��͕H$u2z\��V
k��w�M�映��]ڶ_[�H<�fj�-Q�H��&��1���ݔ�.˭۹�0��(*pv%�M�].P�[Ϻt��S�> D��6X������z���@Y�f��ס�u!���*�U�V ͜ob���	��it*d�]8�ז��N[��ʙ�\�5ȡ����M�RTP��,M�jbyΞE\�Z�)��}�C�3��:����U��D�̈́8�\�t(%�lE35
�!�$VQ�������C8����;) ��7�ԗ[�J�իC��Ld�.%�DT�:��s^:9��f[�WZܙ+z��D�ڬ����D;�����b���T:�2s�W8j��+s�m`�%^m�����|�{(�en��t'lHq�#���՟j��M��}wMs
a�bY���}|�׻C´P�Ij�u5-���M��m/�֣y���m�V�8�r�����M<p��Ǹ��@�OQj�́���AϮ
M�H��\��!�W�O�m�ܝ���@m���:�!��qڎRG�E��r��r�{)��^u^իYYN9l���2Rq�կg"�h��v�<qϝ��E�����N1A:F/7�W�McɲL���Pv\�!x��7��Fs�g�YX���dV {׬��C�4��ssh�W��N��u,Q̈́C�4fbb��P��ڙW�>��
C�l]�I˾.���;O�P4vr����@��tEࠈuڴr�����i��%�����n��[ä/��z�,��]�is�^� ���-�������~n�2��r9c�)�C��s�KR�v��T[�I_>iH�$�K$�f�����m�^2��0❽+��]��5�($W��l���0��h[��F�޹2���]@��3���M�����ϰ�7�ʪ]��&�Me�(��>��b
e�h{x(��g���[���A�{f�9o�4��C����5_��훁�!Ν[�ӊ;n����fRά�ҹ3��Bf��E�e3@�ѡ7L����"!�/�yMEX6�p��آE.*���*pMa[��
���}�:�^�\�Ç\�%����Ϻ����N�96ڂ̷:���y�/�K�g���-�|�����VS9+Ov�N���U�Q@]��l&�8%
5���;�������1��}�y��:n�/������Α
���R����� $N�h�0^�	��9ې�T˱'�1��ݻ���ӷ�
�x��q��{��u�6j�c�˻��v���&ZH���-<6����n룷!z�Wo.t����1�!5��9�S�xi��E��"����s�m���(ej������p�C]뱟v����ۼG[�H�M��2��"r����+�}��T�e�����b���z��/�[�kc��q�ItJp:�(�V����f����7[+�Vv�cN��л��:�#�; dv���\��Cq(G��Z�j�򬮻��]�0ډծ�e��&uf�b���;s�k�SV)��3�S��+��k�<��x)�W\�\�]��ɠa��׹�������A�0�4�pu-��K�l���k[��f��}2�`����x��tS���Z�uAwZ�ul���\�ϻ1�q4��&f��jt�9,Kxkd���/���5�
��:���}���"#��d����;��_����R�+6�>aؕ�ua͗M�_B*a�ul�E��"Ŏ�%j鷖9���`�w\/eq���*Ek����x�i�%�:���L���iC��4R&�:u� ���|�]����(�+ϧ�P������pZP��rFe`���D�Z|�������W��nT+��E�c���B!%{��BD��K�D��F�n�$�I�s�չس�C�M邊|�7y���A�7:��u�G'w�쁅���y��v�����������oGp�$rҽ���.g�s�C3]7�*M�d��r����gK{uݺx˜D����n����$u�]7Y|�f;����]E�p��.�wZOov0Os���vo	9����{}���{�  �����������L��*�e�%D��n�X2#�n��V�S.��Ĭ���]s�JH�Y��7)$�T��뷙��j��s�<,��te���m��*Հl,��^b��u�3;iO�$n��]��-�.��7��ƻ�;p�6+;I��E���<K��$���媜���P���ãt�6�+\l1�*+;S�*�\�]�P8�婗�;B4�]n�uf�b�;����Q
���Y�.������O�O>R-�a\�p�A�l;���J��s���^��{�\�&B�{�6�Jz-JŴu+7u6ƫ��6[��Q%�v���\�])m��>�r=�C�������ud<�?b+u�1�����8���i��X��͎" n����]��T� �"�Q���k!{�n�P�ۛ�Y��wq�*_(�'c�,u{S �Z��IŨڣe�f_Zv5Z;2�(�@/�{�o8e�n���Y���4�����g`��r�pDt��F���קV��;.�����e>��8��a���W�(U����,��9ȹ�/�XWZ�4)M�v����9�g<ڎ*v�9\�p�ŧtN�E?�U�ʦ�l�XZ�������է��q�k�0�zo��G%g#����&�OZ5L�9
]}F�A�Y�B(̦��V��Y���7i�����i�a�%����M�Qv��5.���e�`qs[�U�Mˣ}3&�Q�H 鍃��"��d�������^�0hˮ��Z�Y����3���+�Z�A�`ɽY�Pr�f�+P�oh�r�Dl�[�GU��b8��+�Lm, +i87�m�9Gh��Pn�s.��ս,%-�����<��Hh����6;a�ߠ�䥵/�%wQ ��4�ɖ��4�zWL�m�Ӿ�q�T�hW�5��K?:+6ѣƴAb")YKe���{V������
�k1�ݦp�
F���u>������w#��Y�ʝ"X8@�i3��J�=�R���ZYv�q����57D����.J�}��qP�yIWQ�b�*�r�h7ch��� y$�6b3D��74���;�أ��7�#�ݺIR���� �hS�:�P� k���:���G�lK>�m�ˋ��@c�۔�m�6��6oJ.���ѻ��s��j�n����5��GV̐�u�cKDk��P����@�	\�uWh�=U���T�p�C=S6���/�5d��.V�X���G��j5����oIͥ&Pu�����L\�W4=��^������حki��m<]�U#$ڈGAV��N|9q�_�g�P�z�VdH��ם��Zkc,��_M?tl�8�����;����%Č���X'����m�UK�ug^E���Fkc�=s5�6��2��=""��]��Ct<�<�2�5�z�n�L�`[qڥ�q�.��`u,�#���L��I�;���pZ6�c��(;�m�=�e����B0��Fť�';ś��Z���0+(���$R`U�œX� ��{A�t���&7� �]���k��v ;�b��R�1�$�Rג`*��,��SzܓwN-�b|�b��^��fhs:�&������m7{�ʃԮ��=Cg9�}j�ݤdR�w��ѭ�&X+��Z,�-.�K�h[7d�!P-�����R*M>�]��gq��3Ig�f�I���{�+(׳�w��ʺQ��,���U$��I��]�Bz,/�;�{"x;��{O*��5 ��X���F�5At��#y���㖱u]6���ǅŦ�n�ć�cXf�D̶���[�WG��e�5�nd�E(mκ���Di�ڲ;4 }�Ƈv�4�fc�\"s��@t�ʾ΁ve�u���gb�K��؎�p��*7��4R�n�ʫy,̽��kҸ�Zͻ�U�(����L�3xfvU9m��b��{����3�R�hG9�;�{21��{k/q:��Lu�.�?m����8�˔��G,j.^�/\I��S84�5��{]��&9Z��y$��z�
�����{�#k��نa�+��&����dHI���Y8���ף6�f)�q�	q�VN�n�O�����h�'mM�zl$L�E-��%�fN�j�Hoi��{|->T��t���+�|�]�z:��wT$_ȫ([�^�H�ݣ�g%|��N@�=�dsy�D�GZ���3�$;��&	�b���)B���Z�l8�Fm蛶���yF�T��`�8;]e��C�B��vv��OV���<��G�Ds-J�Ӟ��+.�3j�:hUʆ��C���D�n]cڙQ�z+(�B':irθp�� =�U��л�����.���z-Յ>/5�@���i.�qZ���N�tWK�5BsVu��:�J�:�=ڊ-uh��#l���s��b	�Z���3	e�OU�.U��r���+�ݺ��M�����u�6���sr��me1�CaV8�e֛p�.������_Y��b�Ѽ/h`��%�g�^�N7��.�;"I�V`���y��R�Û��е���R잎QY�������gR{Ye��&�/��ɥ8J���*��!d������0vf �1�d%��}k/�H�{tT������#[o�&|�s$���b�e�5%EYMS��ִ��S&��ޫ`���J/���w���f�?=��SZIHǪ9N�;ө��R���k��T2�ȑwnt=���6C��6r�˅CY���tA���¥{�|;�Y�p�o$Y8l��Z�\�^r��A��8~3,�X�uڸ�/�vh 1�U�f��F�
v)�������@�h��;w]ϊtm�K8;i����/�־��sL����؄Նފ\j���WQ�q\G)L�ɚ�:��;U]�<��v�`.T�5�]�m�jq��/f�(���r���6#)�7�n��$�.��|VX;���Zj0
��u<�7����0zkX�|��Ύ�ܭ%.� h�����oP��Mk��H�+��0p���n@St.b�#&�^��[\wu��V�O-�-�;�ϻ7Su&c2����µ�u����D r�"R		�#w���� Em�o;m\��Eu��o-)��uL١�[��h�e�6�wW�5wR��0gu�x`����5)��N��\�uwN��go:����
�*�_v�FU:��v���\-���05�7�ul+Me^��-G��g��5^��Ex���������f�2��T�&*xȅ����X�}˦M�Y�q���!܍�v�D�u8��ݿM�4Y��a=��oݪr/�KwZ�8�5�˻Z��K�*� ��;f)J��(l�M�8���ȥx)s���A����wޙ�$u��*#%	����z�W^
�C&�rw�S�\�mvr^���2��'k�B�XO��s��x���j}4cGm�MR�H:�#a��.e��ue�ͩ���NWU�K�����9&Fk-��J��ᓊ9`G2;%iN��~5�H� �\��yii�A&�}�s��oEɱ����wX�.��P���vi�[/58|o]i��yxԂ�d�Q��7*��7����!ݫ��wI`�)�b�����9d�@u	F���:�d}ݙq)R��PV���f�T3b�T�Q	���o{k����Bs.�w.F)��!�N�4.��-�@�v��̈́�A�}��vp�k��ҕ5��T婼�g-��)e%7�Sm��wF�c�dP�ڋ,��bN%�
�Z6���Ad��/���+��˶�k�������q�����x�wi�tV��}�l+�M��ۘt9�;Gr��BβBS���&D!�)��Vsy�ݵǺ�@�S��^�]���JR[DA�����f��p���cH���UǑ� ��9s�mk�;�8���L�)��i���v��)�V���^���ꇁT����6%�&��M0�-�f���8�k����l�s��k�E�Q����`�t��r�N�5��a��j��kz��d�տYטd��3�]Ӽ��\��v��!>#Qi�GT�Wb�+bYֆ�qfV�v3u-�.���s��w%�N�(Ǖj���ηxqĮgt�ٵ5X	o\(�d��m�pWY����B���ʷt��읿3"�r��Q���z�%�IT�	�X�K��OP/��]�d�r�B�[��n�R�x�0�m�ř�m]���Ω�����x�W�R��89�xn3Â�0��Ϝpmνߠ#2��E����KrR�cN Y�n�f[-ev�h��yL�p(z�N�Į�Q�Yِ��R0�2.�Ww���f*�^��c*Cݰ���;W|��*���V�77�>�n�{7��1.��ܙV"Y���:��m��(���
�C���Lʔ�X�k��{�e�O���TX���x��ɬ�J9{��\�Gس����h���l���,:�\.Z�gY��-Q ��Z-����=$��/B}���ԈD־`�u:`��zL��h��V���SٝݪZ߃wn�N�"꺐�$+���q}ٷyL4����/��ܾ�sp�F� �\ʊ�|s:��L)��9�M+�'���Vԃ,\v��r��2��.��xc��άw��B��7�&��^#[�`���D�Z��is�q�N��wЫ�W�>喕����m��o�T��)�A"2d�΅n��'��׭R��H"_M�}{+Ѝ����U��_�9W�N����̍�m�dU�R��f �Z�̡��xWY4x*�M˵��]��\|Ĥ��m�Qx��N]7�F�J�c�Y;U�դ��~����O��w+}�`:U��1�E֮�ՠ�vW:��v�M��E��{���κn5�Ѽsu���z֣O4_c�k�W�u��kEX��>�Q_wur�V8cY0�đ���;�>���"�s:� vt���hh��ɉ8��V���C�v�!��Y���8s��>
�u@�Xr'���u4vwo�H���� ��� ���WͫB�/{䨱VX��ˢ�V
��4�e*,s��T}>��ih!�UZ��b�H���x�u����*�|�pL�[�0���A�o�û��I�i쮰���e�}[t��|��nlեc��]�ڽ&mھBپ�P�Z���7�KڏZ��o�dq��@ޞ�o�CF�RSb<Ď�6>�cHf-`�\G&@d�`�65���-wm�+�.�cu�s�ݸ�p�����Yx�u��䆳͡�i�c�Uosy��0e�Hn�R=�ԏ%ݏ�)+����}&`������C1ƹ�
�7�>.�|4q�]�f���:⭮�X<VI(G�w7��Q�����(���ң��_:�5�KF�F�H��[R��ne�Ot�e�J�;�̃2R����E���5�B�/���N���ý�Җ�[�z�`�8�Һc�`՚�pď�*�L�՜{;OWV��� �̺�g�|W>����t�s��W�,EI�uk�a6m.v�P�]����B��w��I��f*Ku�T�X��q���0鮣�����ss
u��#�ՠ�,�\'�I]��e�Q��_m�k�hN�M˰�rU�kZ�B^��9�G���j��V)���+��Q�u}�K�⫵2Ɏ�^x�l�}�\��Hk��Lok�W@�l���V�C�&R=���F�4к�H��+��̆���R`0-���Ք�ުy۩��@s�XCb�*#�[�;F��PssZ:Au#���Z.K=�Ν�M��hS�2�uKQ�A��_����χK��}.�c�ۈ�rl�{�7�=�����GBt�1��m��,;�����b��R�c�cR�c.�^ú��=�n�&��i*��b��@��tn�A�ٮ����R����j�#mג�bE��}��9��j�]sc���#$�ь�"*ҕ���,��E��)+'���r��8(��v�S0�K�f��-pƝ��բ��F�.t�A���"�TEݭG;Y��:��ے�R�߲f�	u�A,̢���KJ��i9�����#�����)��)<+(�I޼�I��|3Gc�^D��*��}��:��Q��˨ڶ��`�8�k8��ľݣ2�m8xPʔ6�s�Hfa��쿴�f�S����e��im�u*��7#�-239�����3��Z�'j�V�N�0�
�tN�xU򐾷Ag���˺�
5'$��r	}Ҥs6�媱5I��1j�*)�K38���7��u��xDۛ��DA��v�$S��K�η�&���"�eY�{B��SdҔ5,��(��6;{�	o`xGt4 �6y���>VL��ݸ��7=˫���ܺ]�I�������C�=*(i����G�+Uƅu�Xre����W�9˖�K�j8�u�kD�֮��ݜ�9�v�ʕ�4/�lU!�ys���J��J\w'
��ŝ�����5fj{��D�F��ho�eb6��fR:M���u�(+nZ�ݮ�CwOnq(��R|2�f�1P�;��1Zk�/U���弔�	�m�G*�l:����B�AA�tK���3�
mG�.����V!��	c0�z��IW.G�v�w��q���9�L�ٚ�CN�؎�F�풞��<�b&�-%t�&L�F��;\�h/�?��5��oWgu����g%BWCҭoB�e$T}��)'�F��%��z�k�"�U�Ac���%J�b��Cn� X��=���B鬂���tu�I����̴@���V:N����$��핫C�J�<�Oce���ЫoC��փ���}$9���$�扦���¨pG��<+!Q����4_ �]�ܵ�$\wr����Y����;io3);(�$�##�8�W�mg&un�H��/�* �Ңb㠳��;�K2�sX�T�v�]Sz�c#A"���[��V�� �a�̼�r�G�t\��ѽ��CVH4o��]���
hC�we`(M�b'0��B�G�j}��TI;,�	I<����:2U������ow%���ʋ$�NH��n��V�x{�������+Ӫ���ҵ��H�m�뵪�e�̉s�c��K\��9$&V�T�1F�.2�S<L��{y}O�r������S�4�s.� %;�F�u�i�f��9�V������/��˚+`/��n��y�Һ^�[E8�r6z�$ݾ����˝6���S�6� �Vb���N[����f`rw]��)����$.�R��.I�T;e�+���=]��h�l葻Hs�g��@�p}'t*p?����xmrŸ���~�Jx��/����'5�L����N���YQM%w��&�y�[srO��T�X�xY�.��a�tC��	$�.ue2dފ��8(B����L���goa��W��!�����#.��S���m<��q��oh���7�[׻�;��Fe(;L��Θ��
j�W�j��"�	Ј�Tq���֤Ɉ��t�׻G�����恤3��]�4a�U��f����r(4&(�}ȁYϮ��3*�g\���[��Z�O`üA|�N�/]��X��[�t�-�r���`إ@L�nv�O�X���U�o;�h=g2+�O_S�7)��VrZ�:����<�]Sq>A`����HX�M�E9Z��'�Uf<�5\��%�k�9'���%��1�W�2+��m���P�֨�tP�-��e�Yt�L6��*����3�t�}�jc�����ݺQ����b2f�(v�Ib"��w	�c� ��tf�L�11����xݥb�Rn\K�� CH�1K��<x`a��e����7H�$��3CL�LRD��#!�<�TD �.]	3���I��be��0d�4���+�#��d��%�D]�/��"멄�&���p$��˩"Y$��J9��	Lœ��fYι@���6i�N܄�#Qwn���f�"LdPh�s��!7/<�4F�˝&b�s��INn�l]v���7u�3L�$�Zr�$��JI(��E
�(����S�e��T�om^̇�>�R·����ހȮr����7H��m��;h�|�H�N!��H	��5ou�m��Xܳg������ɳ��(���/㊕�lϙ��V�I�4d���;��h�Ֆ����0���#��7,{�S>�,��U�{>�J95���H��"�of�qp���(j��O '٥jt�~,Q�6.g�Ġ�
ц.>���\��b�_��^�*�l��李�U���
>��Ga|�Ⱦr�w��LKr*� �u��X���O6�����'n�k����7g"0+����J�Ի�&o��w�k���U3F��A��$iʴ4��vӖ��^`:#�ӣ�8��OW
ˈ�m�l:�Ўжv�m{4ּ�g��x�����e5A��<E 9ʢ��Q8+]K|���~ R�_f���'.q��X���y7{�xRQ:��������m��t�{��+_���B���9xl�<��}D	�o=�q�u��O!�=�!
�?_J�5){���c�뷟3Hh$�%�!�u��i���,��v�x{���XF2L�x밾%���C)�pŕ>e�ᓂQ���D�
����s�aNr��5���~ŨU����O�<}fE�]ݵi��qh�Dk \�RPU缟��U��a�ma�tP{�3}hݱV�4F0�!��5�A�![1�d���(�S���ɯ��!��u�uֆNL5�/��::d�R-���4�����-���+gPگ4���{���p�7���s��0�xޟZ�p�R�����%�z����/�(�� #���²�ZȘ�Ov���^���4�Н5	t�
�)��}�-o��e�s�ӻ�1u~ʁ `��_\	��ڂI�h
�8�Inv`La��}���k/D� �k��s�(!�����0��z�g���l���A���7��r��.l�P���^4k��Н�L�R3�`v�����'
�������p�f�4*A�Dv���p��L�&��ZܦL�܁�C5�V����}��b��7�����(��v��i?;�"�Wl&6{
�t��U$U���r��k;l�m�w��s-es�qi�>��=�B_�J�� ߵ��F������2k���*rm	���)Y���y'16�Nԯ1�n�#A2��(Hj��n������C���C�i�9ܞ��fc���������Ot^����iܹ�s�wn���3Ś���;)W M����׀a�s�Ccң�#a0*�b�oxD�R����x�[/S`�õ1��Y�Wk7���{6r�jr�k�g�����(�*X�C�n����}،��W+��ʢ�F4Z��7d�M�������K�8�tFk왺��m 9��= ���ykV��y���LŝkgZ���������Fq���H���g�h�Q�'�V���Y�uWڲx1žO�\�d^S�����u-4��KF��Q%k۬f<����4@�b�g�����F�r��O��G���s�%���0u���o6k�r��q��P�=IG���ޛҠu-8�<��.Ñq����Y���5�M�:6��\�/�(��E`
���D��%�}N����5�|E[�g)��6bm���&�]�7j�أ�9�b�k��A��$�(�|�������ޔ�>��U��8���8Nq{���謹�d;����Lx.�K�  A}��@�)��0��G������^��^����l7��Y���7�g�`��F:ub$�6I[8Hb焺�z�oe�Y��Z�y��$c�=���r6��s4���+"5l�>�n�z��c�-CjۥM�_��j��Fw�N��C�mTsE��K�os�͇2��/��1�Z"�%o�y2�t.f�`7G�\���8�,�����m���+&��T7��h����
+���U�m
�]�.�J��*����_8�ҝ�����5ͮ̕�8\��:�W`�hi��:æ�h��7e�UglὌ��*��t��V�t8_4��,3�8��1)���G���_���Y��Eˬ�F�Z����wt�.d)����?x�Ċ�η+� &��>q��ABˣ'�#wNY��tm�����	��K�1��*vhǝ��{�p
$8Z����{�u�@�P0{L9��Z��f�U����7~���g+��F<�-���մ!~uLN�#�}���z�u |b�v���c������t���m�5mÙ�w��tu� 1���XjV�r\c4K�B�c5*�ȡ���.-FO�3�eX����mۃ+�E�8<�Ճ��ǣ��ֵ�'�s/����9ȝ5�+w� f!���������x�,(U�\��.T=�Fu�}:ˁ,�9�5��_P�PV�N��fvz�����.�斖(����|gS�
e�.����ccn*��.��8{j{��m�y]�;�#�U���X����ಸ�'`�/C�9g��S.7�ј���g Ic.~��н{��׳C�y�:�]��O �R�O�+
�zr o'H�!��[xk�x�D�쫅�l�诞��0#	W���vT;�V,_ M���I���V���>�ok55�Cv�9�.p����=�ވZ�:]�Z�θ0侾���vn���;(,�O�B�b	qT��`M�S���_a��������K	����' �>��ܠ�2L��t�	�0��$G���m�Z+��	P��*�d��@�GB=�lV�1��f��C�-�dY5��߃r2�"oU2���)�\
���	��I��W���<�%SSz�Cj��RN�Cŵe��8ۿ�4�,���Gm:ս���7�^L��>
5Zpr(vWV�y���8J�:ϗ����ˈ��;z��TD�����Zr�����������]�B�"�u¯=���d{�����딆M�8�\�_��nG�sJ��J95���H��"�&�6��s�뎩x�#�-����s�Y��׼ؼ���> V�bᲅ�����N�{�u�\x�'�i�<�ᵕu�ݑ�E_0���4�O_�	��Px/������q,��3�Y��ו��7�n�.VMʵ�/��n�Z��}+��<�o��U<y����+f�;JG$;�s�k�tD�\
�<�ُ���e?^��E��O���sa��4Ą3��e���A'�Ye�r�j�o�Z���5<���5�o2�}@�i4t�ז]uE\V9Z�J캘�kJ>����v�[�c/���2��Oun�L7�a.�7RD���8��cc�Q>Ԕ;n�\����:��FZ0tK�9D��=�h�+P����P�`��Ov��pՓ��BpV�ഺ|������y�9�=�Ӷ#1y������m�՞X �W{g�ζ���i'K�{�+_����o2�p9�96�t-`�*y測Z(�!W�w�-K���-S�ֳ���,k��!������wVLO�q�:�J5̡|���Yxoтʆ���S�_�8%JH"I�=�13��:s���.b�����F������5��\��z}k��pz2Գ��u��ݍ��g��W px ճX
1z���Ko���:1��'^;���5�j�WV���u/k���O��
��������Qċ\@�Y�!�ր�8��G�9�a�)�l��?':����9�W~��ʶŋᢀ�:H¨����i����_M��Q�C�E�T����T�z��ZJ�=~.ǁ�Հ��x�ߚ��"�K8�'�8U�/N#��c�uT��X��$Ԗ-����&���2hsj#]��!�� ��=W�T�5|H����2��b�P�ݴ�{{�T�WI[7`�4e�q=�9Oc��y����I��X�K^���I˩G5�����)et��v/z3՞�jtSQ�;��b,f�hZj�'p3ǥ����+�P��v�l��u�ͬm���M�R��o+��
��w^�<�n�k���1\+;gm]��ꤊ���M�ro�7�a�i��=�vͿ�uyG��z}]�
�s��ٰ��_�`�E��{b�sQ9St�����1rm��/3׽o0�������@ݚ����X�`۫|<���X3����M�}���j�m�153[ �c�/sT�*����fC���^^R.��"
�Fz^�E[90͖�r��<�XN��-��e���qyk�G�l���y,(U{	Sӂ����k1��lqT`&
 Kn��_!�3���{�3��Z:h}A,�����nv���nWH~W1Yp�Do�G�H쭯��=��9B%���H:�-4R[|NLԏc[���s�\�P�\�$V�ص4!\at���-9��T6��N�kֹOTJWA�w�BSO�˭�T8I�@�O���p$�o�w^'ܥ��xk���ɜ������7s7|9�t��Ͼ�̕�7���EVP�|��'�=�K��ҴVQޟZ�%~��e.���B�.����t����˺Ҕ6/pӂ��8ҜK;�p;+�;J��|�!uY��jpx�$�[�X/�]���{���ƨ�!x[�zT�v�����=:5"�D(�.���AD
�|���9%�ev��{�����D^{~(p]䓕�  ��� J`P�L�xL-7UGK.�[w���E=Y3��ɕ���o.lWq��`�{�����O�� k:#l$Z�����Z�2�@>�C��*���|l#`8d�OhedB歕HL/lɎӕ�;1�64Ý���g0܃�XB�t5v}����GNZ#{�,�����Y��3Me�NVv�{�X3�����ˢ���k������L�2�@��)�I&�Nv�M�+�5�;��w];^���PYg��~v�g�{&>.w�
�lJ���ۙc+�����P��+^�9P�j`/c�'T���b^V�B�ҽBxk�|���P���}[�~�2w��t1~uLN������A��C��*�,��{�zW��<ÚO�p�4_��}5�CvL��\c4K�^�X�zU��C�)×2��J��{�3!zvO<�_K��GӐ�p 1eh���Zȋι��j��4��9�s;Ѓ�~�<��O���Rd[ڴ���<���6��#��Q����1jdsU%Z�O�=�;�ZX(m1�Y
�<A���*vn���>�r�S�����=�9hi����5�Ɏ�
Ӕ-}�����`(�]aX2�\�C�N�f)����*.��4�K�&N���O���}0���X��|T���\P���ۏM�1\QS���g:���'��E��:|��q�"�
�-�<EZ��ݤ\'�/i\@����g�,v�^ӽ��N�I+��1��A!wn��v;D��:I��H��e#u2ƣ�2>[���c�mµ��$��q�J1��x^l��%���#��j@�����0�?���|�j���[|�|��՛���	fY�5�!�i��b���Ͻ��<�!N���Β7�|�Qcu_u���ub���}[�!ؖ�"��nF@v�M㪦TP�\Y�7���Dӱ9E���j��(��'�W�п��!���~U	;A-�lA�d�u�;���]�������L�L�\��"=� (֜E�{�s����1�Ѭ��N�&ػ�Kk$��d�=�J�vu��KGF�%�v�B{V#^D8�B�����_&�}G��e2Q��3�`4z�4�`x��'#��rU���G&ǣטP�>g;=Wnt%R*'L�/�jt�9]V	V� ;`v�F��j�qME��=| ��C\��ػ� [������
��t{��J��no	�#̜r��վy:�6�.���mk=�;�p�{[6�N*)P�.E���%[���	v*Y-�ꢚ�Kh=<���2>�,����;ݚ����(+;�o���C�Bˈ��6�]j2f���xu�k>�K�3�)l�U������p��*�ջ!�/�X��I���c�yT��<�5f�u���=L׻��P��r�Q�?b�dܪ��;��p�<�ǫ��c7�S;��u�F��C�$fa<8ik��\�T73 ��m�](:֜�3��[�:���b����`i�=EzU�ķU�Y������a�ʔTY��(��D�g�Z[��c��� 
���ݻO���6��1\�Ж�.2�}��vTƣ��:$�gW����@���"NZx�jz^���Y�ŕ@G�hOa�����+Ճsg(£���g"'��Ϧ�'�u�v��ξ2�($_�	Fj<��>jK/�`�1�P��T��ᓂQ�JH#p�L�^F7��ޣ�J�����*�"���.��OC��v�i�b�3z}|�8�&�E�ݫ�n���U��%O�� j�:� ���jt8VM���]�>�P��.��r}_g�h��s��ĥ���o/3���n^|+6��X� @�N�"vN[Y�Fq�IK�*���u�Gݎ�9lØn�q�V���ٸ��j�
�����F�eڦ��^�֫�o��]�$�W�[^]7n�R�Eu�u�����>tu�K�}WQj>���a��Hl�UYʏrfP�а�Ij���Ѽ�4Ѧ��#��|�;M��yu�]k�[�2q�{��7�E��u�>�褬�GA_)�'e���"��n,�a1��X��4���܇�{G2w��6�<�zs%mg���fU�D��J��X�o.yK��vSwǭr�&n��U��t��h��s�
��V{p���A�O1�a��u(_)7F0���'�W����b�f[���$\�v��(��0� �t`��f�r-1V�V���]NLq/�).N��wd���R�z���aϴ�!Q��ɩ�B��i_bVŋS6Fn�8���p7t
�:���L�8���ܧہ=�8ŗ]�R��(fd��ء��H��.�y2�.��5� yR��L��f�����V��͔/P�ս��Lh>n��/�����仡��UrPwTn^�z:�e�VwaS�v���P�7o+��k�ޝ��l%Ŗ�ngN	���$G�+ae�|�q}�we��#�Dj޸���7�|��c�Ss	T����5Ԉ4[�����Da��BM���X�|���C���m�9�$�Y��W��d�k����-��%��/XpC��`�z��>��f��V�o���9�b���e꠻�!I�$��$@�ek_
����:J����+G&z�^��I0�,�%^���YwՕ��l�t��S�,u,Q	E��+D^p<���41�����yu�9� A<�gh�_Z�M�tp�Y�pIT�yW��U�=��oH�^�
�YF���d�Y�D�h�D�7�LwMH���<�p��z*&p��!�]{d��i)v�P2V\��
�NV�F�63)���ʦ�<��7{9H!|k����%gNd�nV��zV���I_�w��"'�K���z�3A��fe�Q�&�n��O%m['+[��+[�CL�+빵��}a<�9}��ڗ���[2���S��q�]�D�d#��� ˌ�*����S=��'����������P��X��v��Ĥ�x����'��u42`��e�1f���3m?��-���`5c��t�U�)A�c����Ŝ�N�7��5g}:�N�k[�Y2T��s#�M۱�h��[6F����c
��M#�,���v�|��*�z���E�G�&�{ ��y����AB���bߏD;�R��[���pº�0e����S����B�����u3vK�;N=c�p�����e�5�t��p�x�tw�s����Bi�-N�GR��Ԍ.�K��� ��;[P��G�e(��'�v7��W�������}B�Tc@@&1�\uК_���d�jݺ��6e��F�"e�̊X��dHf6(�vDP�M�n(S�x�B�I�@fh�ݮH��%�nk�Bl&����vh�\��Cx�Y���J2cQDdF�1�3����ԄcH�R�AU˒H^u��vs�Ζ+��׎YH�22c�Rl�$QXd�;\��.mͦi2T�I�E�S�I�\#ۉ�����&�r`���w\;���Pwv�s��\��;����:E612םt��wn%7L�2a�li�M�_�������מ~��#}J*պͮ�(��6<x#��@�K�ؒ��;rWMɢvǙӤۛ�Wo��9���5tL�~�Y�?�9������~~�{����hޚ�^�{�^��zZ����zEx��Ž�:�����_��*�Ϳ��[ξ|�������m�z޿���i��o{���Ѽm�!�"-���c��>���u1�y<*]ؔ���"�!��D�#�3���0m������^��ۻ��]_���h����^k�v���W��s�������j�W��z�����k�okſ/}^7��Ԉ�h�hG� p���W���ݝ�%tc�V�2{��>����u �H��{�}����ͻ��V����~�o������<���s|�����Z��_�=���վ��-?3���m����������l
�>��D��o^�_Z�������}������^��x��ڼo����7���"#���( ǀ��27�x�zm����;�ms\��_�|����+�������������j�[����!#"O��P��`}:�j��oqU��������������?W����x5<�~���ߊ�}�x��x�������W�Ѿ5�|���k�/��߾�lE|^+����z�����~_�|��^�6�/.�?}""�#��F΂|I�8�������<�����W����u�^������ס�[r���}m��r����/O��W��?ݯ��~��y�����Z��ۿ7��߽����ѿo�Ͼ��ݷ<\�H
" N���ˆ#����3���«r
�a��p2<*@���_wߞ[�r��E��Z���w�ֿU���^��W�oW���ۼ������گ���n�������<���a=0:�04)���W��������<��k�o���W��^7��6��ן~����cQ��~����W�������������+�_�׋F����������{Z��W�~�������[�^G@����c�ǁ�7J�?e<��UO��u'���`��=Q��;�nWջ�6�/_~��[zU�]/��|�����nk����{�v�����|���o�zx��]���]��~����u���ѿ���x(�����2јլ);7x��~��������]�����w�=[�r�޿��=om����W<�ޖ�������|��x����ߗ߾W��sow��>/k�����m߿�U��<m��D
}�� � ��u>�D���P�s�kj~����U-��;(]�&�d��]��[�e�!0�|�Dr���-ކ�+���Z�b����;��5����>Qh��p��P��!ۺD����ķ��«�A��0n��{v���xstwn[Gmn��S�]߀:�ξ���Tdx�G��!#�~�/KG����޻�������x���{��ӻW��oּ_V��~}��M�}k��z���{Z+��ן<��k�^5{���_:�c������o�?}����9��s���#���t$���_��_��|���^���������*��{��|���W���/�-�=���G��r:=�8`b�z�~]Mf�͚۞c�G�H��D�X�">B.W�u���x�������W�s\׫w�__ͼU�r����oO�\׏⿖����������͹W�ߗ�~z��p��������D}9�3��ȏyosv��@�lL\�H�#�Ǧ�%����~7���o����+����/(���_�-?{cr�y����+ߝ�����񷧋ž+��۴W}C� \D<D��]=B�xg�������7�nk���������7����^.�/?5���ץ�W?W���׵�:�7����׮������|����ݷ>.z��j�9^y�ϝ^֝���������G�7Ƶ!k�C�7��L�����ѽ/Mx�ߟ>�����W�>���ƾ+�ߵ��7�ޮX��6�����W��߭�ο>���o�^�7������r�/ߝz^�x��Z��׶ޗ�|=7��{�1����{",��$�������VG�~��_w��o��^+�n����^7�7��~���^/��^�ϟ޷�}k�����W-�\�5�וz��}W������5�W�s\��Ͼok����������
<�p���p���̽��}Qw�W�w��W���{o�ܫ�����m���6��.��[��m�|o���@T��c���r1�Q�`xDW95�~5�}^+�o_����ok@���E�.��i�܃:�o2ҥ�>#��*����k�7���ƾ7�żW7�_uݼ�u��ŧ�|�ͽ�ۛ��v�/K�o׍�~y�*��������W��o������[~/�}k���}m�v�����^��޸���~��O�(�G�I���ߞy�h�����4�����Ƕ�zk������zZ7����޼��~���믫z~�����}�>ur���k��u�W���۽ߝ���m⯋�����s;��1���vR�e�8)�aL�iI�X��f�t+OI��۳`>��N��bF��!�����Deo-&LU�]F(f��aЇ8:�ܬ�J���7��N�����w�ht�r�=3��݈�f��/]9�	�U0��E��Ⴋ38U�������ޘ'���1�-�g�Ϟ����z�<����/�z���~���{m�{���?z�צ�k����z[���4w�Z������:�+����������ֿ��ߗ��~�`{ #�:{������|<5�� J������ߊ��k��z����o|���ҹn>�����ս�ھ�޻�~ｯ��o�ܷ�����6�Z����{U˼�[��皼[�<W�y��~��o���f��!�P���1�[���A��Gڼj��o���x������W�b+���/�>����~�om�����w���s~��_�~�ok��U��_��k��[�^*���~u����ͻ���U����#�;0{o|mq��{ܦU�|�DH�~5���^���Ǐ�ޗ��k��﯍�wm��^����7��ݷ���߯��AW����^�����Ӻ���;���׋���^o��F�_���ok�o����H��O`�={���[��`v��F禿��}��������y������h�����*��������}�F���z\�����~�zom�}[����͹���6��׍}k��������"����z�+���v��Ů*�O}�]k��_��y�¿U�x�^�|�������^5�o�׃\�[��yش���W���^�ͽ����/}zk���m�_��|^��q��~��oJ�-����?/y���G�c�o'��Q�[3�DH���?��~�Ϻ��6�nom����W�������5���|�~+��Z��wk��x������׋Ƽo���h6"�n���W�O��{�^7�����#�S>���|���N�ؙ��;���]����+�����޿�ߊ�o���^u�������������o��������گ�������_�Qo�����O��/>v�ϝ鹷wm���/w����m���'�A� |#�����U���;}����������Z�7��������p<"<�X�ׄ��Ȟd}Kt�]��uh�g�Dd(#Js���yd�V���:� ��c���ǅJ�UMk!ܷM�`���m����U2�+�:�.�D�VW��l�nw07��Y�Mn����X\j�6�ΐ��h\�Jq��ws1�G��Q�|��PS��1	���/(�5��B5gT�3���q��֫��LW�a�З\݅�6�I�_k��$���5��(�Y���P��c��Uؿys��}�k3 34z=���M}Ja�X(m��v�-�,��s4E6�F���󛗴��^�2S��=FV�Gt�py�a���:��G	U�|~ˎ��Y�����x�{|��u�-=�z#�`\D��q��Md����
{V#H�*��WB�.exRz{%[&����Ѹ���ܰ0�#42���"u����J�ɨt՘U`-'H�������u�}���a�	�]B��ު�c;��в� b��J.��ɚ���&�R<T�ѽ˶��?	�}�"wU�[��`��YG�&W����V�O��.�D_yT	��]�g^��u`O��I�w���&�V��V25|~t�����M��AJ����u��1�3��xn���s��'�	�W������݊�WKO�ٟ>^:��*��A���t%s"d���˺Z�5
�8Ƶ��C^-�m�>�%`?Pcr��� =�b#����j���取��o�Ӂ�-l\e��אy�Sb�I:P��Q�^0��f��r��bqa�l�gNw���.;_V#�u��}���c��s�(���;Z��D���L0e���>�i�w����e�Mi�㚱��Z�J�F��Oq���ҧ�;�mf��6\[]�������׮7:{Y�ԅ���R�UD�f�l~aR���(gaT|<� �۸l���1��Yz'o=f���$뤰q������Z��pff-�L�B�@BQ�'O��,���}A��e�7�]���3����j�����L��"I��Ϗ{���ƻk���1�k�ޏ�z�y��*�5��<�:�G�z�W\�g�p� 5�@� Pru�ׁB&��'˻g҇O-�:]��@�(����woTT��ޫ��b��ɘ,� =P$R�*�`sg���Π8�^���8��}/�އ��#�½tl�������t�A��@v�Hy�1����.z�=E��	Y��x����~�%sk`�e\81\E�H�T��%mH�A��W���`���z3��zh�l^��O�ÔoÚ���mHH�L�M��`gھ�/��=\z���ד��Us}���@2�}��RŖ~��v��^l�ڝܘ�9��p��wC'"��Wjr��nQv�c��'�6 �P*c2�
�s��Y��+�&Q�`�3_����#>��4����okz��=���E�X⢫s2d���37غϖ���`=Gd��hѷ��p�cE��hm��/�ӧX|NfZ88��r!�=j�c��D����}��H�ui1|�h��#W]�Ce��=�m4�]%���	L�+���V޲r�����BFFfW�"#%c�����ǁ��;�����f��`�Qs�Pn��
C�:.X�*�C�D���쬭Sl��y���j��:̈8m�~j��[�u�wA���&��zN�t�N:	�uْ�l^�� ����a��<�}�h��lP�k���^	���g�!8Q
V�����ɷQ��$���<#k�Pc5ֲ
�!�P]��7P����2��
�m>�M����D��x��b&\\��Fy9��B�q��y@�ˣpܶT�_`B��/Pr�-�̷��f<�@ؤϩ� ��\5�(WIk���}jhB�号���9��^��z[n�6���bU�����C��$��P���J�?�Z7ϺXC�������v]N5	�v#��of8�#`�N�C���(}��d	)P\�n�P� H��Y{X�zV���#Z2L�K�m�ܽ>nH��[�4����� �P�=΁�˝�����Sd����#x�}�^�k��5���ڸ4u#c󂋣���G�b2�����~Yc��Hwub�q�8��V�zGWgbN��8�u�vZ-վؐ(��|=MW_���^�2���o}҉�DŨ#[��ތ�N�V	�٧�f�d�Ym�;���(�5�楓�Q�݈��4t�!�}�:�굝�[�����c������,U����%D����!'��]��^p����O���l8�3L��^ ��;�c��FA�f'\��ot�6 v��֑Չ��ʸ ��N�x���GqБ����>7^J���d<�.'�y��2��S��!�����[C��X�.^���}>�wt�nF��f��֧�U!qm�i��Ddˍs�l��š]ѓ�T��r��	svk���1�u$.a ��,t�ZȽ��O��m�fh
�fb��X�	�L]��V�q2:���oZͥ\{qr�M=f}��xK�~o�d�^n�1t5��d/�=�{b�eL8E%��r���qf!��+��V3\���1%�3^m'o�5�qVFDL�[�I��z-׫�ŭ�Ϫ������Ԥ=�Y:>��u֢�M��]�������Nh�5K���r�?����#w�t�BY��RۏM��W ye��5ⱁ�Gg6W���1���Mt>�d^�ϭ-:(���~�*���SK�e>@W:�����Ä)#�rz����.�A��s6RZ����tU���u���v�I�JwE㶥�&�Q����:����i�`<ŗ��\Q˷���&ˮ��m�F�9Wû[Y�Ѵ&5�s��0Q܇9̭T�8޼�|A���T��v����W����{�7J[��$���Ba[�a����^���i$�?S��5͕�Z���w�{;�3����@�#|�Yp�K1������<�CK���b�zW �#@�+��lN���sՉ��<���A�ٱ]�B`��8���0-�Så\z��D�Ԅ^�$�/jXT.�mv�=B�C~� 9|;
�v@�2+Z�w-�d_��=�ۑ���K0v�<S)��}h�Cٽ7�]<P��6��@�@���&%>U�p���RN�C�Ֆu�a3W%A��[�����S�S�9����Ԉ��U�ȶ{'k��5������Mc�;My\�Z8~���u�2���#�O�ӏ!�I�Zd����@��#���U�j���U�ekgm��P�u�a�T�Y�����f�[��c]C����&��l�|pU�_[���K����/Cc�)^|���Nx�>����]�c��3�bR +D>�n��kO���>��/�h�P����b�]��a�S*�����_0���4�O_�	����������Ҕ�Y�����y!��؝�{\}VI>���{���1j<�IwKl��\�v\���&o!xg���E�!%���1�Z�b�����D(�w���a�5��fJ��)ok�6\y]�Эu:f��B�C[��u!+����<=�]�����a(LN���0H��\5|-X�����K��s�\�l�K�x|��2+�~�s�e��hz��Rk|s=]��~�����3!U��^���ϟ/,p7��ڴ1�{�v�w�����j�������8��gӡ�
���{%�
�*�|����z��@�Bs�'J�v�LD�!�;�WS�]CY햭�t?my�9qQ� �_pT3W�c�s2aE.��<X�B;�������(yA��w�-K���-R�V[�7B���6���ߙ[�.��E0�c !'�xף�x��Nξ����Wͫ�,��-�����66֪[�/��V&˅�A�8�s��iLI1��J�5�<.5㴎}�F�(��A�Պ7*�wG*V%&���#-O�� o:��p[�N�
ʛ���|�\n�S�ǽ=�l�V;վ{��x�N��%��9�,�0!�1{��R���(e���E%��5�Y�[3���0ﶺ,�YE���%y߮���4P�gy�$�����/VӼYॡ� �Qq&��G��s �]�/ ;&�/�ekSUx@*�9`-�q;*�� d:���ѣG8ժ�ߗ_Y\��w�;x�#� V��O��G���S�9M��wJ�,v ���9���F�B����ڏm�#���r�_ꯪ���5U��1S7E_�>��(:�A��6��UÃ�\D�pkܕ�"����)P��fq����z�c��5�q�X}�5��>KjBE2d�ɺ_���6~�,��5�����t�˳:y}�=@俲v��Kj�P=�{6��o4�����M�q9�����`���n��*М��c�0Q�U�X�^���^i�����Y�7�P��f�YV�ig�>��.�Y�N��xְg�:�f	�G٢�^R�#����H��⦢���*�ֻ�q2tl1;7�x熹P�w>mR��ֶN�!�G1yMM�ʘ}�R����ns8��F��0�/V��UP��(1�ߧo��_��k��6/�+��/^Dķ���e����i����J��4GDEf��ŉ��8�h����B�,G`%�ۋ%�q�����~�G8&�Й�����b6C�B/���%�����	�{g��n2&�Jx���I�r���n�kQY\5��p%�D�׷����t���<�=��G�ʝ]�6�A��f���*�O�2�"�uv���� ѵ�iק�v��n�Z��dn$���E��`-���X�m�$�ϭusV�����׹ث��q\����0ܠ��t�9O!v���f�=.���7i���k��Q�j�]�窲����3��W�H6�!�M->R��|2���<���RѳY��'
�s�uL[!U�"w̌�y��r�nYY��ˇ�6�o.�4���>����=��{-�����Kmc s��.�����
.�:��p��rI�7�vZ��OҗfW=PV%\�[�]uy�t���;�V�@�������Z�3��[p��k$�5�Y9�wsVV`��*HFmj[�Dw�*W�N%Ւ�=v?�x�|[+�Q�w����d�6h��7Η��(�܍`��
�X��d<\4���5�[͌��m���Li��4^�9ï�5�3m$�8�m� ��X��w���E��`W!9]�Lb��Hw,�"��M�6/�"�c�4�:)Rt�2�%�G�J�Zu'v7��Z7��SE�X�ר�fqG8_9М��D�(;Ś&�t�S��&>��Z���u�n��5�+U*U�VE7B[12t�\��[]+���xQ��t�!/f�|�m���k���`0��r�c�Z�(�q�ţ(��ܰ�AK}Z�,��C����̴��PSٴ��@R%Y��J��a�Z�Q>�VlsnwR�̴��p�ok{-\4�,<�	ꕈKx�Q���Q��Hq�mm����g[ה2b�F�`�k�^�J���a�1�;�r����Qu4�>�*)����Y�eİ�V������B�h��V��	N�z4ʋV��f�.��SR]�c-ҕ�/��XT����^n��wn��.��Of(�U�uaW4
�Z8���t*���)5=S��{��K�����#�밓��	�gR�����%��� n�i�]��O��W��Q��W���!�-SA���3�Mal�P���\��wBE�4M�9�=��K�v\���:��,"���x��7�p�$6c�JrvB��Ǣ>�{{i�X��]7m�:gm��m��]�nu���|e1�ESYu��o:<l�ق�o.����M�>�Y�%<���/1N8�&�>�ŕ�,�u3�wi�&\e-2�@�t���Y��hcnL�v�S��E��V����O{0���B=�^�D����ͼ4d���F��#��b�uگ0R���˙1LŨ'W�F���=+���ti�yJ��s�
�PLP��:�7��]�w�&ohJPY2�[�6ä�Ƭ]�/�T��<�Y�2��8��Y��
ܹ:����,������upM�J4��Y��wX��A�z���c����2�C�ct���e�K|sB���ʘ4��YoaM�3Q�.�y���:��3hv��W;�]\�ch�(�don�y���\�sW
��c�K�0E�&I�H��7�v�J�F2!]ۦjR42��ZI�Nj& ���w^-���DF��W:�.]#r�h��.W9rNn\��˚�FѶ"9�4�]�č�LI��T�9s&�$�	��b���%�1Q�����˳��F��G.\�Cwq��u��vm��X���s�.�TY"���fF("Jr�&�&.rK�0��`��b�6L	���^�Qa+���i),�F�S��@�;�)(ƱcHc����;��9���mr���""�9!bC�̚����,�#Q\�N�+��s%��ll\����������8jN���$=ǝ��ӷ��-�dM�B���U��{;�q�ٹ+��}��'�-��S��e�6`�1�6-Z��{��}j��M٘e/3R.�|>?0n����wyV=YiW�$�o���x��[�&7D�&{i-"M
lN��!�f49	۸~�(�ڰ�d	)P\�b�|�73.���i���;�5�N�����rb��x��~LpN�ͯ)� �}��s:�.z�vq\3�z$�������6�t��k���wf�wsj��m��˕ أ��˭�c�z9��}����a�H C�C����׎	-��f0B��%1>L�Y�]���Z���-�*I	�I�����q0�tm��g�CsQ����$-�tY��xx�;��kqi��=���U����ҩ�d]΋��$EmF�b�3���\��W��xR5Y��v�H������5� zq_X�TT/}p���v�Yg�T���g�{�B��P��.��*����m��C�|-7V"��f�A�KfDg����<�:�i��d���W��]cSX��3�T;=��bq�;+��!��:�'v_����<�@6cd\�� H�¡�mO�]�������|��خ�m�n��ew	(�ȷ-�
�iM�AVm�j�D@��&��Z�GR����n�	������R6����4T��Xu(N�4�G��Qt���"�@��w
%��������(��x̱h�Mà�,3�ٸ&�P����A��s=5�n�K�e!�.�^���g�&48Օ8p�&_sJ3bS�=�}��U��|�;�5<�w�lj�N�l��g5�u%b��;�^�9`Zg ���\%����b��,��?[�Wy^4��t�
Hױ��\�&	�7t�i���d^���R�b�� v� ή�%���8[O#r7��u|39�;Q��ؐ���p��u禧�lu��<z4���H�U��m�#vi�;z��/�{^�$�H�#DtB�]���c�����6��K���[Ń�]���͵�KTy����@0P����e3Iz�v��7��������^9h����ל@��a�>��?x�t$C�#�Xn�W�Ƴ�Â���r�6E�X{�# u�C�'���^�.X���)�qbsmx�� F����5���R�c�
Gp��v��_P�t:7^�-��ӻ�����M%�{��yOJqr~FjDwQE��Ⱥg��Z���S�E.�A�b.�Gk4Ek2PΕ�'&��X2�gp�@N��đ��A�߅l��}�k�2yU��]���
Ϊ�1�G��1v/������h��ч�Qb���O�"��:����w�hh��q��!6x�G�q"���*�z�>��:ǝ�l���>�����sB�qzɓ&*?{���ͭ%�2�1�0.#�����I�Zd���v�S�r�e��)@���̯U�w���8�|���ᡂ5�`a~�f�_�G�	փ���>z_���ہu;�H�ĳ��g;�	Z*�n��?��lҝ�|� �U��uW�Z\��SJ��7�&�y���@L`�|-}����ƽ�ᕇYB����C�7��,gˉښY�8#���p�w��İ�F�L.F�Z�������dܫ\�l�K����i�>$�b����p�M�ac�;پ�����J�*"�QU����8���0E}�&���4��'6��y��ɔ9�}b.Z�[�^�lS�ڞ6��~�u/� n��� {��g�T��FR D�� f���[�#o�u���t?o�3��7p6$��;�X3cgkm-��lB��EiB̡s,n d#9n���j��D����V˪�{�J0-�[�WJ@��L���wS#D��ey;x|Ԗ|,xF�R[p����_Unu���hq$�4׷+q�mo��� v�34�W$����W���2�.���-�ݧP+��Q�/�n_�j����w۪���z���r}�2�( j�ݜ77B�w�=O!}VH�>׼7J�����W埇��� /��_7�z�Vϊ���o䤂$�`l�0S�T�k2��r>R��;H��˝����R���TQf�����8}j|gQxP5�G�S�xR���^I��]E�	|~>��竔�K^K^mn��8v���9��>B&#"Os i�V��a~����D����W	�-�1���WE��YE����aP3i� La�l�շ]����G����գ�m^},�2��r��mla�p��"�'���%~j�X���45߶��B ����Q̦*K��9V�g�bB�)�F�t�����&����w=]{˭p^1�������1ym��Ի�Ö�k���;�ࢽ�p�,$H�9EOP(�t��c;��i���F�.�*���^A^�b�}e�Z���nlO��iNH���kW��u\=J�"ل���5���0N(��� ݑ���t\�|'G��Ǜ
�{t�y	�B��7����� �o�n��.Ƶ�wl�v]����\.p۴��k���F�tU|�G
C�8������
�ǱW��Fj]�첞�C�(�{S�^r6ㅜ9�-� %\�Z|&�v輤xS���'��.�M�z�W9��6�)��R�!�j�{�4H�h�c�uX��%T
�w��82�wB�]������wr�����|c@z�����`<�{�e��y���ע�v<޵�>�.��k�<�*��:�İ� n�,���DH�kY�y86"��Ѱ%��=z��I�m�XUE�:i��K�4���>@hvk�j�PĲ进���/vY�
͕��Ɛ����?Q�|{�
^;OQ]��P�-z#k���rb�V?�8\8�/+���K)�Mቅ��Dq�Ϩ=�7��U�
�뎒y�V �i�U��KF��}D�u|]%����"yD��b�/��s�#`�^�N��F�5� ���1��J���x��>�.���e����;Ԅ��Zzq�1xSɂ<̄'�BuR��D ��s�ջy7o�3������t�.�΍v����z�5�l��������۩���@(N8� D��K-�����IP�I���6tA��an�=,�����a�S޾3��B�}�cr�eߜ����4�;*��x!��N����sY�BF�O��"��-(4��z�+.H	�jncwv!+ʹYލ�$e�/㩗�M���/x��.L�Ⱥ"8�^�[���n�q������4W;�n��{���v����`�V��Ţ�^��يzGO�/[��,��� �wݽI�3BV�xOgR{�1�;�^���c+Gs�YUGO�t��,/��Y}��H��3Mv:�*�/Yp��5�sY����i\W�N��Y�+y%Cf:e7."q�\/c�k�0Gg+�����Dz�k�M��]��9�/E'�<#����_y�|9ɠܨ�ũ���0N�5ON������w[�ɏ�~7�:�����E+�+ţQ~��= �ⓐ!��bw����/��{��~���)��>��M�0�'��sq��ia�_����yC�	�[�"ė�s.<{N�%�oAR�MM�/o�}ȗ8z 1~1��*p�e�F��(͈�j���U]�GΎ��^�jf��n׺9y��E���a�Ӟ����ޙ��g��
��Y\#a�)�0���r��I�[�dU�󋗺� �'C�z�9�v���}fE��e-7DD���&utW��҄2��ݫ���;�?0��J�2��5�u�GcN��О��� �+��v��\O���Z=��}x��:����}M/�~�1�����{%��#��4�����X�͘����pt"�m��^�g�p�J/�iZ1��4�w�^��{+ �h��g
��� xթt�ϡB���I[J��ܚ&e���P^ ��{�̜�+Ng-�[��Q�a��Y��c��2��#[�vD��Ԯ�//��#n��"�7�*�t��a�m��<W8�}G�0b")O�N�O��q�PFt�7]�Bh�k��=}�Jyx�d��Y����營G��D���b��=�4�HT;�o����kZ�e��X{�v˷nz�^�nq�3�k{z�I�p�Br�����m�2���1P;�LJ|���pܣ�~Z�1W�c�:V�EhA�ݖ|�J��e4��NM{fLwTLFē��C��UHg���K&)!�h��Ya{�o��-�g���-}�2���#�Jt���{B�0@hC����-S45�<v8���ԭ���^�	��;�R4=㡂*��f�[��u�9+sQ�c]��M�T5
����v��<=���׆a�h��.$^�@�֖�j!ɸq/<�QjRx�B7�5
=������{cx	.��h����^v.5�N�YG�Ney�]���u�|�2���fL�dM�4&1и�5�`�h�1j�F���K��r� ��+�����,-�JM�����~�՜lc���k��+�%�fw��(��T*��n'f>^R�N~ʴ<g�a�4����,�>n�^g�g3o�9+����� ���ھ�k�Ɍ�D_�L�Δ�>͞�G]�yY!N�Z_3�������:@��ս���MT���%���7�pemΚ�L��Ck���Unl���凗�}Sbd��&Ů�ýp'b�d��{�  zv���7�&Hm�\Ki��]G��|��8��gӡ�
��3�ύ��|r��R�]r����L_�S�tD	��#7��+ ���-l\e���>g.*9 iV���;���#�wXY������F�˙q�0�^��:כ��/���OelE�e��7���a��]чG'	�,-�RH��K� 8c]����aU[��i!�˗���uj�t�������1`^=Ă0������R��.��OC��ce��U�S��N�-$�{�lu�>/���Jmx�� o�J� �-��t
�op�5�2+|�����$8���a۝����&�:��.�!�Ag�>"��g(����^�Q"�Dw�z�^����}]�u�̋�%y��"�ן��!�� -%d��~�襩h�W,OEwU�^E��~��D��(uw ɤ�h/�3^�X�N탛%\�/����o���� ֵ�4���Q�|R��40���W��D��<�F�6�7ڴ�{+EdW�̪9�� ���`)ݥK��`�ACw�j�0,.�5���A&�9��yʅj5z�ӭ��)m7ˡ�=妻֛�)z���I��:�b'��!�{�窀ʵ���so�!���; 7�r\)c��v����wӯ.���Q���~���.���yz'&#���V�^�υe*\��Ǽ�p��T�F�N�8*�����ܯ�m����}5�%�c�s�����b��cXj�'�U�uF�f�|�Ʀ����Y�]�k���^����xh��%_r ç#��hM�uiQ�k�'\�W��:����G�c�M*rޭ䩃pe�Y
��ب��=���r�5�x�n�S�$Ǎ�u�ρU�5�=�I�'z5_�Z��cO;��6���U/y^��p�|z>H��*���_�9�����x=��/��׬G>xZ�8.�E{ܩ�T�m�Դ����r_m[�X=�xv�{�|$V�7"h߯�brb3%ӭ�)D��奷�S^���l�{ ꨑ&�fzq���2[Ǚ�,���T~� 놂^��eD6�#z�0�U@Rrz�J�o3����*�j��L�i�k�-�k��l<AޛC�n�,���!a��ꝵ���<�˺w�ɫy�qT�Z)�D��֥���ڧ�q�oB=s0����"�y���R��{�����Lo*չ�VegWq��ڛr��V�K�NY��)D�p��u-Y�7+�����A�\W��a}�r�h���l�Jn�C�Fwꯪ���E��ϝ�t>�vc�b޲�On�������m4�W��w1���Z�Z���s�<������6�o�os�4�;Ę���2uj�K��}Ad�����[j
,��VH[_�5앎�ٽ֐oCMëE*�GA~��w=���i�p�Z�S.V��Q�|{�'���#sc��Jb�е{��Z�N��͎�X�\lsV�i��1��w)w�Mc°�xK���R����g|+��c3k� k�;YΎ�P�q#'������%̌ۛ�]Cu��|�(SL� ��Ŕ��F���q5����F���S]hO\Z�s�k:��C��t-�;@~�-��w�n~bC�䜹2�n	��U���}j�zjl늮;��;;�9�Xg4��a��j���^un��ϩx�}��l�S���.�k����PƷ�Oȝ���J�N!Y��h��;G+ڋz��˳��jli���s!bq+�J�a�3΂ϋ�5���%�kCWci�qf���9�me-S�#�4�1�"+���$˓���śx��/l�i��'^	fW�{�@�Z�<�K��awWR��I44x� �@QX�j�
α��Ԝ�W5.Z/������	K�;r��MU.ё���[����0=�aՖ�e3���}�I`��/E�vhDi�@㬚�m,C�ؗZ攁��0.�7�A	^޲
���j�]�ۅ��c/��fd����.�)GG���n���_��gW*�����W���6�=K�ܡ��;�{��eZ2��b�ǭ�[���-�|٧q�M}k�P�ׇu�0���V
bN�Y�^|1v3Y��۵����p���+Ub��n��w�emw�׻Q�w*�`����(��f2*���{n����>�l�-�u�֯����%4��')�Dn�Х��U���q�Lm ��(e�WE�G�aS���8�Hg����}�i-Ї>�@9�o)��
r�V�#B�����ɫN�Z�޺ h�{�s���O{��Ǒ��)ڮ�Vj�!�bN7mjݧԨ��n�t�t�O,������H���:�-hjyCy�d�]hݼ�*��Ul��.����֎��Yz�;GB#�ՙaҦ��a��p����N�)Z���mɷ:m�l��%�,ز�]j����$5r2���0����-_,�jQ7���oJ%��^:��8�]
���i>��i-���X��
����
�铡ZT�XT����HS���q�l>ݫlWwW[z�غ�T���Ջ��8jV�����i4�V�[K�L���u�XR}�Q�lD��L�[h$y氐����K	��d��+�}*f,��Lc�uԍ,�˶9[@�L��V�s�Ӽ�c�&w#%��7�#�S;Se�pU���d`�M�ڔ��W)(C�_}�Ig#�}Dwo^.����6��:��yL�YM��fJ�S.�m\V�UӚ��w��嘃o�6�%�VG$WN�W���q1 �-U��R�1�\�f�}�I[���n;�:�t��.�<s�rq��a�:�a7�Ww�t�!�d�@���K�r1�9��{aeÌ�qk�L�a��TN�2��Z�X֌�/�,ł:��4M ľY�/^H5F��u���n�D5MWt *�o]v��Jm��uS��`�ևD��:���t}A3�vV�30�w=�x>q�5VYu
�Zu��mO7���B�wF��z=����I�6eK�Ћ���³�)զ.V'\q�c��\��YJ��;C���6�Jt�R�{`Ӻ�R�:�Z��0f�ך�z����p�v�U�2�Z���_l	�}W�csoz��n�E}��H��b8򹝧.�7ų�e���c�é;�,�B�M�>��3�35LW�j�/`�j��Q=u҃!��$�,d�M�����C9�4�D"3X��weQƇw)#;�˚4$��4T$D���&XD�mб�"L��M3\����v�gwhьIP��c�I��RĘ�E�;�KE�� ���sBck���2<�F�F36J"�M�	 1I34e#F� �Fܫ�TW.��(H�����u��r��b6�5�b����#`��,wq×Z1ΕQ�l�;�]�i�ܛ&�i1�urq�ْ��`ĕ��ē9s�%����ɱ��.�� �E|hW�R��13�j�]�k5�;��[\e�U��u�:I%҅T��'�m���_e�:����Ĝ{qMl�͍�1_wZv��zw������zϣ+�тL��gw���U���U��L�+=�k:�y(܌&[�󺽅OWGռ#�b��oS�E4��^�
�=��f ��u-˟���sk��E[��(�-b��_U��t�|��z��2�!�۹ܑ�	wR�e������VO�J5䟞���xS���gc(mK�k-��q�n
)�}�|s�aC�1�續��������j'�Xr?y��V*�m+��m�������׳^d޼w��&)ϓ>L%,�ϝ��nٹW|Ƽ�A�8�I��L�[��`ד����K���7��6ty�fI���oPe�:f�&�术�P���2��;�P��:�"���oWU���o���f�M�l8��ƺA��5�=�N1][�->���w|y��,������*�\ط�f�{�������צXA��#�q�̴:
ݫ�����U2�Y(�Q��{�0)fɽ����Vozr Xc����ŋ����u��T�;�M|o�����X�i�|Fm::��G�m5�M|`3j������+2�C�&&&�}�@���{����^5�����������9Zv����^�����Zھa�)�Ś��w�����ϵ�6��"jXlY]�4'�|�ݩ�B�ʵ]C6^g���.��ʥ{w޷��\ ~��{�+	~�J������kWV [%���Z9�O3ޏ�ĝ�N�W�x�c��~Ƕ�U��9�̆�E�/MM�x�t���uY��	��~�V�����+ǝ��w�Z�Py�v�\�2	-��s'�E5^��log�;&�a���|'7�����z^�P}���æ,ޯc^Y�W���	 (�lW����{,�B�	��m�/�+�d^#姱�O{L�@���yƶ]��:Wڪ$��J(��o���׎�y�+7�2��=���//8�×�j���t.K�"7^E%����N���&�=���Ĕ�o71z�w��曨�-��e1�Hf�U�R�����[v�˦����x�/�h-U
ѫx�7����v2��g[�]i����F�d`�<����=�^;�\9^S�G�]\��e�JJ���q-��c�q���BCuhCb�U뢳Y�YB��d�-��aku˫n�M�s��ﾯy-�ޝQδ�?
�9�莧�`7�l��ҹ�k����p�K��T[䗫	�U���f1ϻ�Ư��ʼn�y����=y�8X��T�����n��6�i�f9�����Nop����M�:f�:l"t\�2�E&�wv�քT74� �=^�R^9/jl_\�3��ڥos���NV1���z������>�ڛ���Bw��ס=B2�ۺ��_^R�xQ�w̓)3��U���:3�v�W�b1sk� c�:�v!|]��[��^����]�Y�i1z�c�e_0�������cA<]��,�l��y�'tm��X'1�z�о�s�4�Gw<u�r�з��uf����oN>5s�x���2�B`FV�&�М��lV�u�ӬP<��w�^ך���3w�i6,�GK�	Ϭ9���uz�-udf�qe4�b=�6�ܜt:Te��ξ�m(m�\Z��E������w�*�@c��1D�(ʂ֊����x"Zv����N�6`��&NZV��;�k�w}��Z�Ӵ^}�=��3v�3�AM�<�V�.��镣0�v�Ŋ���5Gm!�`�şx{��N���V&�>���UK'n*��U`�BK�'�m���Os�qq�t_E��ql������t�s�ЎS~�s�d����'�Vg�{�萺j	3ǥG:(���a�w^��e6�Z�j�6|�#������^�3�;yt�=Sޓ�������(�Cz�v�S#��ģ�eT���Uµ��e���Uz���s;�����{����i���iVpS$��=�m;��?P�*���}醯�� �b
�&.�՞q��Qsk�n�y[�9ե�hl�ڄ>�{(Oc����y�wOwn��wh��ef0ݜ����KԪ5魇^f�4���.P��F)=�P�f����~Y��᜽g��:����fKze���b�6$s'����=��9��t�+B���[ʟ�+�rfy����{���W1���^�6�ŉ�PtOb��H��g�w9|R8u"�@F���5��X+)�U(gջ`Ѭ��S���G
�KTT&�1���)%a�x�A�z3�S����2u��Ա��0Rw�M�+lGt�u�Y�/%`��VT��=H��pLfg+ѽ�)BnK���\pkΫ������}��U�M����oN�Ս-���O��R{a�]�ʦ���ŬYX�u���`TL��u��]���&�Ի�^�B��jfywz�����>��es�������7������p.� ���*�n|w���&�!ꄙ�^�S&��f����-^+���dx�֧o�qnuzm.��l�;�gV*v��R�%Qq�ע%�f���d�nMs����L�UL��/vҥ�Sn��˨R<���[��߂|����=z�9�N�[�{N�5
=BGK˧������
iɭ^�������~���{q-=�+ڣ,��0,��f���ӹ�ڧ 2�T'�F��G�ҟ.*����}�#�]�d�\�-Q	Us�o�Z|��U����n��4�N�)Yu��N^��l��oF?,����b��ď�U5��!}�La	D��{6e���fmh�ԕ����3��=;S���Q��B��(s6T��WRIp�+��-dj񬇫n�d�DnT���{y�΁@qeÁ���;���X�aQ�xk 1�ڟ2��漰��w]-����Ÿ�޵Y0oB�gf+����׻ۈ�޽o���`�T7��$��#+{-��A�8�I�z����5���ݜ������s���6p^�M+e�vϘm�1͹���kH[B2����M��J'��Z��dK6�zdr�j���9��L�n�ؑΜ/tӜ�W�qN�o������pԜ˔'��z����P��(Wk��lc�3o	H�:��b�9��n-�(�y[.�.ы��d��W�74���ޯ�5�s�鉤[�:1TK����p���n��|�ݯO\Z��է�]f��/�*E��'z�J�S�vپj�[T�{1w��O���5�D�ެwq�ov�@ךA�c>I�r�O�o�A�0�9jwʊ�WJ���!��Q�	�~���/�����b�;�߳u�v,;t�VhNl !Z��$�:����7:�<;U��"�f��=���K������y,c�+Ȃ+ekghd��y�g
��S��X��R����l�goj�+�jE�G#�	W��q�_r�^��a�\E�(/�D��Ճ�<{z��[������Vlr�� 楪��+r�;T�xDzM��e%y���j���bc%D�(�蚮�� ����fX���,�r{"5�/T��V^�G�������z����/'+F�JV��fў�x�˹o�Nx$��N5���n�z�VNP�ڤ���baRw��ϟ����a�K@Xr�����&�{['n�#I�cϡ%���M��b�ޚ�i����׻��p����G^��J�5�Ujݗ��?V�j���s�7�;git��KC����\@����[��cV��p/"~��&/p�I�W��7~f�oiʑY5�N�ò�����,�>f�L߳�G��a�v��g��|�8x�T��uf>S���7f�ji��Q��k�j�]fxs��Z����J��U>C���pW Y�Wޯ1B}�������W�<�W��]�x�/�~�tϝ����Ww+�{��T��lF/sk�#A��E�/g�k��ٯ�}*j��}NR���k�'���L�U�^��%ۭ��'x��3&�ˈu.r���R��xв��� D��)�!�u��n��i|�l��tk4�9�j	}�� 7nB��Ԯ��3��RKs����U!�W{YJ[����u�9�y�v�K��U_E����0w%}yj�m����T�9M�/�XK�Z�>����B�^:��v���Z�`��Ƞ�e/{V>t&r�]�~~/5��W�nx�O4�X{ޘ'�p.�c=R"��ڗѷ��^��o�;�l�#�C�<�Φ �4�z��?r�9��C���9k�>s��(�G)��ͭ���1V��P�[���!o�v���G�}9Izxv����#p;�z�I�sK�`�p$��Al�i�z�+�	��Kb6Kك������,r�/8V+oq��t&�k����<���o�m<�S�Wl%�,��5Z�S�-T�^�uM1%ه��uD��n�C�a�ޛ^曬7���Kd噌B�����S:��>��Rw�u���۴#��[qx��o^H��f.p�`��z�oZ�ܷ�r�~�&0������Y{�����_t<�Y��1o��'���QN�;����r�_��kR��+r�)��q�ܶzqፊ��	@ә��O�uۖ7�/�I�U��D4�Ꚇ��ndգ��]��Y����I�6iS
R)X�.H��n3|6�,���u����Ӭ;����}t��(N�:Wj�x {�{M����|��)�������d��p�En��N�u!jOJ��Q�a$�l+�}���2��}6�?b�貎Ob�h�o7/����4[���(os�A�-׸؞b���blb2��`��b6U�rk{�j�bs.U��޷]ܥ
�8���\f�{$k6%��� �J)������Ɩ�K��3��W_�Z��2��q�s�X�: �� �{�����(�[�Y鶗�������s�k:�e�w1����7w��΋I�qW3�6��\�uŮ�w�A��#a,��m.�>}5N�e�U��ǮjO�8X+�#P�{<�~�W���A'C�-NSShO��S���p�gWv���o���y�������U�����G�Ft�`���.�1�	\P�w;��V�nej�/^�{�����4�_L��ݛ"^��ќnmʈk-ۦ�mJ�'���z��We����]��P�fh�Z�ze���.s~i��)��Z�m]�u9v���)-m�8NDw,v<�B��˸5d��C5}���D��3P�ڴ�&!��Q�8w��&ӡ7c���9����)v�c�WLE`�_I�<7��wP��ۍn�7��/���zj&��N��myr^�_X�����B��o�R��/UҔj<���e�.�Щ�>��m��X���v�FQx=�ތ��\>��;���C{:+���p{T�nM�+{�W��Vöm��`�e�����z3^��Y������ ���mm%2L����üY���>�T�L��-�F����܌��cE�N�S�]Ͱ#]n�4�z��)��_9�!t�bCďw�����ډ!�Nueo���mVw,�Y��j�u7��.<��}	��s��図PM�_�g5����dg:��M7r�������v�\cʇ(B�̓�F{ݜ��X��5ﻏg�}6���Kk9{5rS7���CQ^�瘸J�0Gъ��Db��1k�٢.�K�S�֩�UV%����U���v?2y�ȕp���X��[���o����z��>S"ؒ�2�+��K�m~��iˡ�C���F�pçy|0�MP��\��%�@�Uכ�y%�P�v�FV����Q�͔��R�<�ͱ���Z�@�)�;ӳ�6��$C��l9�)U���
���4��k�բX��-kؙ1gT�3b�E�ݾ��(��C.�ؓ��'���^���6h�q���*Y��-���րF�Ḅ�3� ���}øov��s�K�?��RF�&��t�z:JT-N��X�Kp<w�Q�|�r�2�`nv%�d�8��X���*wR�_CF:As�^�_|�7��#�t�a���&P�P�a��HZp���ՏO۔D�Sڈ-7��dE�"�Ÿ�n�6Yܜ��6�hZ6�w�{9a㣜/�2�aŊ���9�*���]o~����Y4��5'�n����SVvt��cY�k�:�����bp�7s�����Q��*oP���Œ�] jPlf�������=��`{b�
����H�7���}4ҼT�8E�׋Jb���\��&�MA�/�=��S�g��Z�^�˷v�۹�Z��h���e��k�;�3�j	�ugWHɡ���؈7a�N\Y9����eqٛJ� �����K��V�D���Zu�#�L�M��4����	�x�քH�䃾為Q��R�����/ja�D��l*�����)Ex²9uʅ�എ��,���=Z]F��嘗Z,��OǮC/�9>�d���IwB��i�
�t�v�zI�J�v돊�q�Gq��H{F.���;{���\�S�܂|�1��riz����j��p���cw(7E΀7�7�Dn˙��ۺ�4���-�psȨb������}�])����[϶��[o���,����$��r�p�<���\w���o���P��i���s[{���!������R��,�+�����sTN��|񳼅����z;��Ch���t鹝���Q��)_@��]ա�3�";�Ķ��Y���G�<ٔ�v]h�u3��b��YO{�%>�ms �`�ە+Ήu� �K��E��Z�o�5�\�l�.t�vFj���D���@㊘�����d�uN�u	�$]Q�N���n���a�a�4�ԓԬn�D�۟.H���+�<�mU�Uv>�ES�y�T�f�[��aR�j7��c�rؕ[��S����V��FeŴ��p� Es��;JuJΔ�p�������u��t)-sy���wG@Yr��1���Ρ�����,��@TI�-�F���K�܎�$Uŕ��p�ᖲ���OW�P�7Ҁ�޻7��mQ h�ڝfjtI�ע��]ࡷ�N��"����a)ڜ�x�XT��J;�kv�b4�s�݅��I�}��q���	9Euk'9Y'+E -s��}�\��5�9�_'/M�&N7S��g�_���~_��(Nr�r�#I.��+"��r9s&�\���h0b�k�D��@͢��;�M�7
#Inx�7�D�1P!�wv)61Hb�E�"�RX���*)��Y�%�ۻ��ڌl\�1#HF�m���c�(�X��;�wRi(�jI,�r��[F�(љ��:E�c���F��ŋ��Qͺ��Q��ƊbU&M�- Th�4I�ch�Hٛ7u�Tl�1h��"&��nX��,i�X�(��nW
�m�Db�b��܃F4`�5��ɵ�͈(*6����D|��(���6��Y�d��3�6B�\�V͜t��1gw�pL�|Zh��=�Q�L��!�O@ooxK��2�;ݷ�s�T��W�<=���떰����{+���Bܳ�nqusT1��E���yiϑ��7�ms�LL\M���c�L�g����*~�|��w�yeܱE�ԭ��c�sʁ�/��ìnG���hOOQ��]{���'�1=2���}O2��e�v�.ن",޳U A�S�7����ꔺ�9���t�~��f�iQ�E';���4'��w0tʰ�_�Ωڇ���g_{���F�J���R��'^XG՞rS�Y�e�����r<�oP]<m+s��V`^��t^p��2Ri^��e6�\����Z��`n��}�\eTv���ۊ�m�_�P���;4��[X���xm'M��K�Rr.��^;y�fi��SkU�u��.��x�gor�̄�q���9.3�+9g!���ޫ��]��.☁�Ѷ&�5��{=���C�n�7p�x"��$��cS�z�)U�X�f�\��c�3RLx��]<��x@C��<�+����|ܨ�����ʵ/v�ɮ��\ǆd����n=�⺕�Z�4�Cvb�]a-�Vf��������Nd2�<����V�>�2�����faEp�Y� z�=7�]�nT��M����0�=�'���ոy�g���0L��u�֮T�Y�g�Gh΄�G�:�
�Snt�2��%���{1�r<T��84��n���Z	;-nh�m�;AV?Q��x�6o��9C�G;�&#�݌:�x+3�o	����EW1�،Z���,cPv�v��q��啅����ڥ���S���P͹V��켫�B��g�ǳ�a5O�kz�	2��\�Q�רC+fyNֺŻ�*v���'w�ҟ��/#^��D[�.m��zs��>w�MM��|,V�u�ӬP<��FeN#���녝��QRN&1�_*��;��P�FmK�^�W��τ_�,�3�g]=葓ыxs�x�}��K��f܎����_����;��=���í�ی-6/���o�ץ������}���j��T�!��IqN5pņ�6�K³��)��5.��\����;�P����Rl���tK�j�${�o�{�w
�>a9O�t���x��V��t�!:,��-'��BlV�fp�fl8P�a���ǦRX^ֽ7E\\��IՁ-�an�n���[���磌=+%�x��2����)J�v�V�7���9^���@���G4(ք1��Zo8gR���^��$l�tC�^S��w�ހ�����tC���*z�������bN�PZ�������qx�00oJ��\����
���P͒����1�%1=�Y�^�+)�j��R�7ו7���UC��)i�:d�1ڄ>�{(Oc��'HP��r�⽜�z��4ז���w�6¶}	ӕ�.P�����r�˫ۙ2���!���2�1LnhT��֤�aŽG�<�	���{�z&�]�����)&s.�Nmʾ��v�wr�\���_�_ӀL�K&��r]�_��ӻBz�W���WX�ko�g��sg&�@�fI���[�t���{Ԇ�{��Y�Is���d�MZ���+��Y�/7Η_u��x��aӜ��vx���g�}06���(��%Q���v���k,ǩ�cR�Yo����@�z*�FG���M+��X�/�p�&��V��wi,KF��R�����q�,�ٶ3�4�uh]M=i�"�;�p%\m�G&ʟU�w�G��Lz��Yɸ�y9�s�Lx�괴~�iv�ŵ�����k�O��b�nS}������Qn�7/6���ⱞ�ߵU��XqFf�X��um�F�S�����a�b��ϯ���ɫ��7%��rw�yփ��	)y󶠮�'�P����·�����z^�j�)��s��4��V&��7ݼ<bG2�Cf��,�e������C�6}C?H����`��U�:h=���VDR�|������P�}��N��ə���R�^�o}9QϷC�h�zS�VP���B�·f�z��1&����=���l�.�����FGw�^�,ӗ���Ν0�{V���W�����o�VK�Y��`�k��{wٵك�}�>�l;B5���D�}W|
����y{��W�{��6�/9�(�k�:��V��)���8�Y�9�c����*�QZ�A�Fnإz���g[��K��&1k�hS5�Ϟ��br\T-6�W:��7�'v]�֠�6�j�Z�T�^�� �_v[0F�o�#�V;y(W`����3(q3��5hQ��DYkg? -/^�RuP���f9S�r��͎C�\�s{�,[�8�u��-��b�%�}����k��n�b�˕<�5���?+IT��	� �k0�X~ūf5��608��E��T'��Nݩ��.+�4�~SN�5J�<��3�v�7�qB���͡�ZX�l���"�g�N��}���T;t��Ŵ4�N�v-3�q]�!�����7WU���E�ة��w��&�QV�'���'�-�d��3����?���ʯ2�� �? ���0����� u��Q[��5ۃz�TA׮v�[�n�k�r�O�ϚsY��ti7A����}�Xsk;&��^���"�f���{{��N��L���{Ө�������	6]�3���Ĩ�_�eC[Y
�ԇ� 6]�˥��.�nn9i�W��rUց�r��� ���G�[;yq/Gc&�D�r���b<��N�w �*-ܺ�^b�q4)�n�m��yv����'I��]0�{+�����T��K��ǥ�H�,�H7s�+�p.��H��]�
���u�.�|��M���ަ1W,c����uZB`�j�\�za|�߫��n��Y�(��ؗ��k��,m?m<*�j�]�Pt>�,�SCԯs�z�:�|�3��LI��[�P��t�n1Y�ޛ\�c(��oN��B����Ù���[���S�q�++�=�^���~o2�����$���qZ5Ò��s��2� �c=���ر�/+�*�iC�m��8~�5���9���wV�{b�of�d���ڄ1�e	컨�5�y�f��!.W�GI��p�H_�Ƹ�z�Ϣb�M9Zc��'��������.l���`�l����ٙ"�TέB\&����(N�r�=B2�����G&��Ŭ���ʾ�2�m�⮬�EW1�6�b���,N:��c��Zռp�����X�f�;vr��ʵ]�]���M3����Z����
}�k{܎A��;j�7�򵫽�?��Vk�������v���]LNz�)���G��[F���=]�4���)��H.��{�&��N��乫��I����Z5]�Sj�VJW��U�e�Ht�ƹ�����;r=��K2j����2Y��X�O���ޘ�-��yeB:&9-ʥ�_�������զ��vk6$���5�a�8�Z]������u
3����}\�=o��c�zGϻ���_9~Ǎus��n��j���z�|4͊��-d����^KHb�>[�%����'iTn��r^���.�T='OkeX���w�����D�{A^�ץ�h%�֥���"���]��SLI�S=�^]=�����#�|����5ا��y5�D���ɬsg�(��8SjN�N�����}����zmS'v�I���b,vFј�H�^=d.�
�{���_ue��k��vQY���Wce�%��f^�z��֢b)1���$�rZ�oIDw{9�w�>1�7���T�U6�+2�����/E��ޥ�}��>s.R�*�d-��a��{+����p�d:�+!<;��VsC�3�z�jŰ��f�VϢa;sJgٰ_M���>z�4pдl;LF�+y���װ�J�[y�y)�I���ҥi&��l��"cW�B�:�s;yM�d�f=N5m�BVJj��vʽ��e�Mܦ�<�q[̽u��2�����-�7@m�';K�y��X�b��4 ڋ'\��r�޻��w�wﾯ�jw�N�6+k'�۹@[�͇�wj�7�ï2źlO1BF�sg1)�SX�-�fu��w������G��X���<��ِ���Cn1�#>��Yn-Q�h����W�͎ڽom9�r�4�e#���f�0��GJN`dT@D��nn>H�YLs�M�+�	���/M;S�z��� ��.��Bp�H��ޏfm��O�[��Y��]��ށwǶ=�h����`�#7�]���έ�"��}���X�t��ϜO�j�X�w�l�<r�����Ξj=�fQ��	�~��_��@z����r��{�j�<�M�^sC6:�ULu;͢�FX��&�K�r�_����w�����0�nP6��L5�s��.�"��Y佑�:В�O�,�--����{�̭I���6�}^���s�FYx����b�B^��])F��^NǨ��[~��"�n�\�W�c#;u$�����/q�uGV��\�!)r4+B���۲z��Z}F��3��~�с's�ي��\Um��&1�ۢ�JV 1�\�
����/�Թ��zNw���a-ɷ2E���Řr��E]~��C՛4q7�X�]�<���mף,��oH8�ؘ}�I�v�W[cm]���Yn��d^�h�(��	�Z�*�;f�K�:/{zH����gfő;ٌV�1�H�u���^�o2�q4���<��v��3��u0����c�&*+Ŕ�����i\2�6-�m�Ni�$�,�]nƯ6��ؓ��/\�)��Y�';�BZ�7����kꜷGb�{��'{`nVezB��.�h�Re���B����wt̉�Kw�3���v����U�z1�3k�bƴ�Bz�)���O[���{&è�a�w[��"�}�m��Sb1���-c��4���wp���"��,�BN�;��Z\K�^�V�hn�����ܳ�-�.�XMS�Z[��4c�E���{�H	Eݙn��k���z�оi�Q���o�<󊟢��()�-
��(�'��-�n���3{fCp�7i��I��׽O-<�t�h��)Mer�wU��:��%8l�ww�Hѡ,�rg+�ħ��(ʔ�YCIޣ�E(zJ�ꆪ��ê�d��5�V���TY�ҝ]�t�[�*ZO����b����Бf?���^��^��P���#^��<����5�o/�z]3�S OOs5��e�������z�ll�����wc;K��	ٳ�b��1Q9o���眼-���r
ـqTI{_J�^aRV�I����>z2�a��ٯ6�Ծ{@�\���w�Ы���%�Ή^����vj�Q)jk������>�y��yB�/x�¾ޗ}�fg�B�����������	/z�����wA�>��@;�|��e�k#k=c���6�"�k���>T�:�lL=�:�=�۵or�̄�K�oseH������^u�OTQ�^'�~j~�%1c���b�
I������m8U��)��.>�'Qђ��^�9>H��;]P�����.�P�M��1"�x^����7�J��p�I ��a�lO�ӎ)͍1ڄb���Kۗ�׽�[ڔ�x�Pe�0L�,u��/.��ht�5J�������R�s�sut&�a$��2n&q.���;66�sEw=��b�Ƿ@V�Å�u<�]��\���3��֬�7cq�:�T,���x��9�fQU�t;��p]mr��i�`"*�$�Y�4���#�C�7�X��y�C�@<*��yv2	2m��Mϓ#Y;Q�ۼ��l��Θ_io륐VgL��2�ȫ^[*�=�:��à�o2hh�fӓv�vq�6�eYO]f��;��AD�X�9P��2��p�5Ot�1���օ��c���Pձqd��ŷ]ί�oј�\h5Y&fuͽ�ME������lR�(��V�N>�v4pW����R�5�x�@��̺f�z�Y��ʋ���ꗖ2�>�v�6n�4ukt%#&��,�F�Ǩջ]3�Cc�[�ǐ��/m�W��n%���/�	��R[ݗ��q�KSp^�cT�E�yg&b��g��	|��M�d9*]�}��u018T�V���I�V�;:�ٓ��\ys5�7�	Ә�1r`Y�˙$�B�f���z��t����WȥC�$K�E���\s8�����Y��M�*��nu� �ݖ��}.N����,蹮�;(���F��Ai�A�ۋYy���x��u�������4�e���VK��A_"�b��A]�t����U.B�p��� [��*�HtLl�@�/��v�R�w<��n�z���H���ϋf�9�y3p5ܹ�ˠ�e��]I��Ԧ��q��pF|�(�����W�4�<�sw�N�u�%�kC#��H��6R���۳i՜��ƈ]ó���'Y�(Ư��>����vT�û��Ss�v�TF��8$l�X��i����Pۆ�МX+���1�W�Z�w�EL�R�\�k/o�j-L5W+H�[Ba�7�m�s��V��"�̜��lӺę��n=ڮG�%�����r���t7+�ܗ���������v��" ܣ)4�i����o�3ʗX
�j��b��2x��:D�35���ƥ�
 ��|(�:RӺ��]�'�v��Np#�#�U*����:*�n�rf-�[:�Nbq[��ؔl���ΖWf�ӫ/w�\ʗ�Τ�.
�u�7��4�79L2��_N�Rs�GM��n���"m=��꽧��o4��㾧W(mSk]�A�"!��GA&n�[3�\spc�20������J*U���u���-p��31-q]�ظs��u�#X`���}�j	)ջJ�^�af�'��'	v����Ww}��$^]�M�Lp�{�.�.Tjj��F�,m�s�kc#��g���Jrj�C������g#y�lq�=B�iıkt����(lAr��'"�8��W;j�w(���k�q�c�{�Ccq�Q��-S�E.�{h���ǖt��d��j}W�u+F�^>`;���o����u�E��Q��������]��^�������w]��r�6�sqɊ�����Lk�5�QcQ���M�:`���1m�li+F�cQX�k�kF�r�tֈ��sG+������d�*��nV6��O:�+Ex��H�Z�nk��+��m�v׍n�*�1b��wW�^7��-�x܍rܫ�x��m�j��ܢƼW6��ڹ]5�m��Rx��4mͼo7�Q��EP_���Lx�R�У2����!.���ބF�7�����u��7M���gə�J���V�y1���v��/���i�8�ua�?[�ީ[��W61��bF1CZs��De��������y=:�j^�mf�������R���b1k�@c'Aյ�S�v6$�8}x۹�Q��9;v]��됭Wn�z/�eSL�79�u;[��g�w9��9�Ϫ��O�Mθ�|�+Y��\P�x�Q4[9
8����ï���PF��l���k-�뚺����{�8�s)�>:�j�L�~�ⱞ�5@����g�ק���q�V�7"U\b����`p�ݛV�r��p�*��d��V7j
��M˅�i�ή�a�%s���W;�-���|�{G�W>�t�#^����1 ���ݿPy�#�{]�>|���[���P�,���S�[�Xg<�������f�Yc/3	�ȇ'��	=�I�wJ������󇉳B���!ó�3~bc{�� Q#60���>��`ڭ�{�4�u�8���x�9�`Y��ގ�雛�m�&����^����-�gnx��Q�dk7�j��Ҭ��46l�5���b�^��Ӹm�����'���GkF]_i�}�-gN k��w�Vf<������e�+����9Q1�RueֿR�Z�B���Z�E���f���qx��i��̗���]ԭ���u�E�vCF�S����˺d�L����qU6�&��=�'���#{*�{z`�{~leځ�?�)��--i�6)���&�(�>��p^�8�|k9=�竔)u�r�=�*��г䶦�&-�p�8������NI�E�ȅ��|��OÚC�8�r��o��v��)�1��NT�-(�=֛�W�jXދ�PtK�u�]���z}uj�7]l	�FnSC�m�6�-!���i���貱��OT]�V+9Z�<׹Z�;h:d�'�x͝Z��&v�5�,���ɗ����~�w�jo��1P�d���s��{I�e���kM���G��˼яmz�\�xs(��,L[n�%=�(�����gsq�z��I9�;�m��(�KE�Z^^�B;ɥ��7N��{��WU�l�Ӿ\�F�K�@��{֎���W,g+iە�Q��ni��;s�Ӑô"{OE��/�.��*��#.���B��$�k+��V��L�\�5�c{=�t��|���b�>}r��o5[Y:"f�s��ik�W���7s ���'�j/P��"�����=�z���]CZ
YR���p����ю;.�v��%���wPZ^ۍo��)�g�t������	{<�4<�S#�t��p{�;�I{Ժx�/����iF���bII���S��@;���ug��Nσ�K��v�\r�h��l��'l4��\������<���m4��C�׻����]v]����כ��]�7A�;�3ս�������d �A���#��Yfjng��?v�P�����{]����I4�z��1M��)i�n2t�Ijy]�[�,�g����9S�r��r769{�\�oä�e-��Oe<�gL�����pU��_�u�{]c�ծ��}j�=|��qk�ssrW���g���{)��u�����N�vGFkj�>ʷ���vb����N̋��E����
 �e`�46��*�("�;��+흆��*'� 깉��
͸��<��+���ٺ�Ja7}]Fċ�ص֨'r�%�(��y��8�K L�Ϝ��^��A��C}���Bz�e3�V'����U���n�Ӹ���1]�YC�[W�2�M���XŤ1����.��,��1�Vb�;d���c>�V��s}$�3K�OƗ��^ǽⰗ괥t��<T3/^��,D'Z��b��šlM<����񟟳�?2��Ŗ+{��{#3�˚j�����6GS�C�p�O��{Bzz����挣J���S�Rv���:���Q��j�A�@Oӧ������M͵u89fun���Ł�{:s9�&}ϗ�d���e�o�`����:�#^�dΞlfo�أ�E7�oK�^���˹�B�8������;aT�7 �q3m\R�j<���ըx6��
��XW�.��T5k��Ws���>�_9~��פ�tu�:y�y�>�b�|�M�i�fY���IԻJ��4ZwOE7殠��4��Bс�5�]ͷ|���< ��W�n���+��u���qe���U�	Oz�h��L��w޽��'MGfd@8��J0��uz�31+P"]�iƣ찳���s�^�3+�"Go=��B�^������q��ۇ����_�Γ���5�������hG/F���iV�Ea�꙾�ꋵ�=�쬨�)�J��-����v9{Z�ow���W��.6��֎��~����s~��l�j0�=��컨��_�(��'�Ǩ��3 �c��{�øG�)����pe�}����&�����в؍��2�s69{�T���%xsc6$c'�����JUt��g��*r������k,��i�R{q
�8�،Z���,1&��Z�;�S����0S���^�v����3�B�]@n�����M3�yV�:���o:��s�{��w�=^�XM{��}g�ե��r�X�W�N�t:��Ӽ��dЭ;i���x���XS�|��"�.��(#<�f��Z\K잹���uo&���OI绎�d����Cu��^g[�[���w	��sgÎr��Zc�Y�%���c��/9�@[ѻ6� s�T�����+
,�ء�p����H`��>+0�L��v���6Ej�2�	�[�J��q���3�:��K;���љ��u*����}��h����m��m� Sw0�s7�蛳��˗aI��f�y:����1|$f��^<��˫�o9z�d�*��R��n��ZEN���y��j
�rkT��\��"�MoCr�<�/^�=z�>y���"L3RDt�����xn��D��2�])J�����^x��מwj+�0��pw�y�����ޗ�=[�99��BYw]�+:ݴ�$���{�0R.7���R>�sgo�XW��oI�Dw	�܀����'�㓸iS��4�u�v~�I�ե�{vf���)
�>s�kb�f���zx���¤�\�h}�:���7p�gI��$y��v���}�G����W;޳�����/ӗ�P�@���������^ӎ�͉Nܢ\��t��^�>�"�<�V�N$��r����<��� ;�J{�:�n����̐�*�W�K+v���@��҃1��b��W<�o��]���(W1�:pUޫ6�Y��u��(�
4�X .��g�R>�˱�xFC�#/Y�K���q�8�� À㫘;A�aX�Vk\��wl#���YB����?���u[}eS�x��;m��X46�u7�:��<;��w`3
��x���ɀft�X&�G���m�Y[��}�m�#z�����%ݩ�yC:��t��Cik^�	��^�{��]�;Ӻ��SL�78�E��1")�.�ӫ��O����N��!�U��y�q�fr4��w�,����]���ػG���\XX[Z���&��9�O\Z����@���O[��x�պ��vn�0�d�A�N��N�w{��o�qo���iz��hOOQ��iO�q��/���kڛKr�<L���k��A�Q.t�[e�! V��6�=d������>�x�E����J$�g/���;Kb6@=��;�K�<7�7r�X{�Uz�j���z��t��-ZZy�{U��U@ك�`=U%r���1*���ŕ��*�75�rK�����<���{�E�ug�{zA�.KP�\yLg����}����oݝ�C{m��x��A��B��އQ�+j"�ys��=0�(Fb�Q���w�$ma�U�MYp���j�c��K�إF�R�+*ί^�{����6�@j�k�yD����d*�i�[*�p��XhrR�<mIbQe�a�A8�ޱX�	�i]�3�i@�Wz�O����l3}���͔���D����'�m)�����-�a�,�7���q����n�5w�3�ݽ���4��d����^k`-��)&��^�p�����H��őx���J/k�0��:t�#X䬹�G���
��;���^�ǣ�ޯ���B�v7E�.'l.�r���#��\��r����*/!4z�$����:�d�|Ԫz���^�6�ŉ�Nz�'�2���ܓ�#p�ϵ�p��G�3��7��7�7��U6#no��b4gm�.۹��Î�����/��S�dK~�V���5i�Rg�]�~^R�=����$<����q�{-����I1������V>"g+=�~~O4Т���8�o��� �A�{�l�C�Z��qnw�o˨������ݓ������~:���/K~�'O)�;�Q��T#6���<��کb��N(�����xF����!�+7�v2���v�	�]�}r��SCm׮�yy!��� ']��q��zW&{(��dH�F\�c���+uֶ(��i��d˾����O`����P�v�Ԭ�|t�J7`��켷�ɉ��t����%wkΡ����{����k;ɟs��yl��C�X}�=-/:4�۵k^�ұS
\F�
=��	�m�z��{Vo�N��ύ����b9�z\�roj&V����^M��j����w���Xn8�԰,*e�ۚk�`����}�}y	;��u����>��a���(^���YG!��NQ�=d.�U�9���Gp��e됱����ڎ���r���>|�q�s��z�+�Ny'+���y���;���J�U���)8=��^�+��������+��E}m�$�F�[B0��J˰�\�<�ۛ�v�]����>/͝OY�އpͰ�Btǔ۝n��ԡD�] 8wW�kl���B�Չ,����{����8�͌u���5�:��G[����������~9�m!�t�e)���R���b1ss��Q���خ13c.�k�7sQ�(N*�d��.��Q5��m�F�|g+��6�^��6�B%�wV<�ouf ��л�9@h��T��:�U��.>v�mZy5[��53�G���-�K�:F��h�f���*.����z\���ǼE�t0����C�s�u�1�Ӫ>��^�3c��[�Jmg%���Vu��]Cv^U����Ƣ��-��z�����2})����P����<99�:V��A�ᡅ�Uem856Jϫ�(^{Ӂ�9ؖ"	����gzg�N��'f���_W~�yU�����ia���gh�����Z,�a_k�މ��s�g�� )}Y��ި��Y�Ft�5���kN�%b��r��a�݅�
�X��ӧGDW�=���Q��j��0���O]G�b;�Y���HвR띭ڒ�����{q*�ހg���S=��2�2hr�u Zc��wu>+�WR�=��Nd�AQ�J4�����]Z��G�'��4k�*��������ۺ?i�Gh�g=�D=����4��u˜�Ցݪ���Q�~�8w�6�ƃ<IpF��ʡ��e�$���[�A�J���o�O]�����C���>��E����ܨ�ئG����F��]�9 '5'@��
�t�n(�/JX��3��_��c��2L�Ou+\|zs���O�(�둗ul��<v!����6~�}���D����W��x��q�ڛ�*38���þ0�Z8T�}��)�=J��ë��W���;nJ���N�t���c;k�Hٰ.�zou0�8֍Z��	��&��!TB�b��͓�v�N��\$�|�#��0�\jT_wol
�j㖢̜h,䩍���^�k�Gv�����T}C[�R'�[R�#��T;]51S�r�۶IAlx���N|%v㻮�p��2֑�s�}ە�a��Բ�[��}�n�l�q�
�6�xVS�F��b����u�N��kG�����E��:eY��8T+��Q���N �J9��#�Y�`� �w��ټ��\���SyZU�l�kJYӴ�y�nm��&���4)Px�),�́6�"�Q.0GmB�tm��iC]:�u�����}�,�]��%G��Q�]ʖp���3meA��+�m���a�@r��q*��1�T��gZ�`���r��(�/�=�]>3i$4�c��Ȏȧє����ϳ���oӭ���)�f�띪'	���{�Fj�Ъ�����i�[�,�#�8Z]�x�*�)F�}|�e\������+A���;�Qܠ����P�(wC�Ub-;t��PȃCZx��Ol��_tI�v�*�Xާ��ky9��tΨ���v;�pV̌cBS��:�cՙz�}��n�ȹJ��$i����wUڋ��mc��{�Xi�z0+]{���������,Z�Gs� �Bp��OX�t㼲%��n�����z˖�\n�೻77�z=�*L�G�G�w&�Z]-�ٝ�{:�).wy��6����U��/�E�����i`���V8����lF���L��:�p��H[�ӑ�C2� �ʓ�H4_
K���kk���fɽ%�êޗ��iV�b;C�����ͫH
ӌ�v�^k DVl��l���c�EZ�Dk
Ǐ2����K��R᷀;=�\�am�nom;�	n:�	"��L�1t>w��ܣ���]�7kp�\���S?�$���Y�p��i@�h;ת�n���_*	rG���p�!�5H�n�y򤯎jN�qNt+AӊQ f�	v�.SX�ʥ'�\��xi��O���%P�/T��'4�����>����7�+:nk�X�.�F�n�J������s��Q�/j�j"�8��ʜ�ci��j1s��[���S"�Bar����!�
�uq��z��r�{��R���S�*r[㱘3��7)�GRoa\��H�.��n���ʽ4$YZ���f�W�7�gU�8��2�B6Z�vnU�[`��̜�s�9>�t7�Cf-����Ji����e�:')MSf�I�k_#�f�չ��
��|�4��ѫ�ɚU[�6���Sܘ�ϝ���0K�XΣl!����l�܉P=��b����_1%�@�sһa	��%.�+F�V��ʚ��6����@��d�t�\@�p�H�C�i�}��K�m+����Z��h+�Ruqi�����U�Ʈ����ڹ�kW+5x�m�m/:�Ʃ�h����K+ū�η5\"�x��c��;����nHh]��h�ۚ���Qgv��&�U�<�󮷍�ΎW.V�Z���on&���E�x�⹷5FѢ�[���Z�Z��<u��s�U�x�%s����y��TV��[.��I^#[�9�v�E���cN�\(�u\Ưwm�76�ͻμ��E��q����#�/�����Տf<�MD�!:�X�mhTᙺ����a�쮻Y	��n��1��
@��>ߒ&!*S�q�wgk%v�[!r���\#�̛��W�����6a���g:g0���ێ��4/�URͪ�Ǻ�c�:��Ϯ�Y�������M�r��D�Tym�w�j�1�ܬ��tϸ��c�2!������̯MtI�����h�܂���#���iѸ��Mac�m�[UCR�%��g�����l�h��^A�٘�Μ���P�z�W�z��d�DmL�����C�X�/�nj��n�F'}�\��V[����2k���ր���r�	ux̫�l=7'��WVa�/i�ixOޣ�\�.0[���P(��z�FwP&��u�w��g9>���F��x+����z�a��G;�GCM/z�*�#ㄣ�ӌ�VV���)���w���\%{�_�G���3���H99s?�jˢ
����[sY|~�w}��N��<Y7e�M�\0�U'��}yǸ�սk^w��KP�z��gL�\�5���'��f�N"�צ�� r��б�ˮ�k����q�b���?�,��mm�N[j��Tx��w7�\}gĥpf;��~��FY��ʡ�F9ӝ�n
z��-�C�������[��E�l�J��5|ҧ��q�wO,T�(:Q�S\hp��Y��Xv���1�FP�SflQ'[�aW+my;l�{k�W�rdti�a��������ՍN�Y�Wy�O�o��.*#=Qٮ�#�ȃ����[�6��v����m���p�G�Hlw=��(��T�أ<��3FL��>8sf��Oy�Ţ���K)���O��p^������.ܠIU:r�rKs�=<,����_�fϺ��r�H�3я�����/O��K;qخ�Vq�D��Âut�O�,>�M&3r�չ�pk�;&/�}�Mτ�u������r9I÷���UL���<E���Ly�gE{�c��q��+��mMzcj#˯G��{�lnGun�q����PxMm����gy/k�a�_{�*p��/D�lH�S�^~W��C�;c�=H��]���߻b�&�X��y��f����ﹺ�۸��u]3h�-���K��2�VFT>4�B���Ϟ����.��ڶWlI?j?6��8� 3������۪�T�$򝃳b�^�
����r|��/@��5ˎ������ݗﻝ���ɾ�7��P���"�W�S�G�߆χN� 8i�R��J�w��?k
�k{����c_k�w]��'�� �w]ޑ�Cx�v�U�ǻ��;	L�i���qa oc˴��= |xT�?��ܨ�>�����Nl&�x>�8�����5�t�۱��uMQ����J��Ƈ�4����Ep31�a�M��H['.��ڠ8 š���!��mXAɕ�K`o!˘��ߞ.#���C�K��f��	��?P���V��8N^JW�~%=�}#��fw��+N�owl��/3u/k�fsԏk�Ne�����Wi��8d�}^�=��w��!����t9�զo6���R*�!��ϕ`����r3ϫd�g 9J��H����DM��1"�O�k�?x��{v���A=ZGD�щNGvV���h^s���n�K�xѝ�W�H�p9�1����6\��f��S0yH�I��E:����}q���b�m=��$���	�:${�����z;t�s�zCsxeq��y;,�Gt��w��u���Zi�DZ�
�~��פ��%����o�~�?P9����=	������ა�c϶�;}��9��;G[�/���o1��D�<�$�� r$\�̒����E�:}x9��:�z����y��+�^{90���=bl�r��^��R��"tf6 n@�;+��
߾B[O������&/�q��g�Wa�}�_.�M�uHێ��*�UOK s��3�n�P�zz�a�I1}��.���A���ٔ��0E�ڣ;h�XN�������A{�F��ϸ_	���8�2ڂ��eݪٹ[j{\���)��o	x��+��5m����`=ƥH���ڥl]
��8ŀs�ՕK{"|Y�n�l�y��G�L�x�f�>���l��fIq}�i��i�9ӕ��u`3|iê�,_ʤ�6H0RHn�վ���պ�eZ���C: f���u�j�M��y��3�'��`��ć7=G"�ey���v�OT��%Z���;;�����W��k�ޢ�ڻ�	��F����7���f�&��a5�������O|�Vy���5؝��+�"+���䱕���B]wB�Ϩ9�� �¨<�3���z�W�'��z#��!�#�0���h"���51��Ī�N/���bOn�����9W�L��XS����]��{z�9@�r72��W���/	Á�Z�{�+�2n��ӽ�z���d�!ӵK	����U�W�;}���Y'=�D��L����AZXZˑ��Y:�(ί��j��p�t(����u4���ռ}ި��mg�ʝ��ؙ��{���=��/k�;���GE�H�7���@�ռ`8������\f����c9�R9v����]zw����}|=@Ζ.*e�t�2�&�+� ��c��wK�+�P�I�J����៷X���]���7����KQ�g<�{�{��>�|w�ztQ�FmƲ�ܶ9ѕ�����-Xw���v5�0r�(��gotb��-5n�S;8ǘ*�2�Z��.��ǅNs����󑐞NT3��7���;���}b�`6����+-�ɚ��o��<IUa�FU1qS)����I-���=D�9����W��`��5���K�G��סi�VR�}E���Itf6 �0�F[7�L��ӹ�����O Gj�K^�ZD��=��;�Π;M�v*����z4�����N�!��P:[ �丫�7���6���Zo���{�}�p�#��8�9�p��u�Ω�kU	�qE�L�����ByL�H�ݧ�]�����w2P�M�����t��g������A�̳��a�o�Ӟʜ�Jj�dW���ޚӼs�Q�!�����g�g�K����;��{�=W�u��͊5�]S]F���Љ���7E�����:�Z��.!5w"�u��Z�9*�V�qԆ���-�7|�]@s��d��׎�
^��a��C*]��Ψ�=-_�Wfm_yoA'��j�S}��i�C3C.>�2�R���
�&���h"����~��.��<��b�[�P9I��>�}�>�:M���N���o9>��� �P}<a����XU�E�KN��c3�:�dP�x�IR���$�<�SVe�WOR�����e��r'�[4�� `�S\��k*��uf*&�i�c��/(�V�v>������1g{aL}�k�5a��:P�h!/Y}\]^�ZHV�E*�����ꗄ��ѫ�ێ���N�gUp�����_�O��?�Ng�?W]Waɫ���1����+��V�	T�x����	���ϟ�z%��DwMq՟oZ�w�ɟpw�'������T�#�����?T	�X����r+�`J�hr�w�{�uϥ�_�[��l���fֽw&��g�����.=�6Ot�ٝAח�q���>�eP�c��G~�3�9�x��1Q^j�^���fMt[��u���C�eH�(��D��|eT9��.eӰ��L�"w/&��Ff��r3�UX�%ݕ���θ/}/-᳒]Ô	(��rA�����{�7������v�~
mw[�fn1����r����l�v�\=���=�8%�p@M9�V7���2�G,B�A��)`��鋊����n�K�Hxl'�m�Rp��g\N\uݳ����/X;\*S��~�z|{`�����q�;+�׾��.�s��{�lnwV�&�ʶ�E/�髿���iʟV���l�����2΁�0w�uH!��a����������q)����O������Ҟ��,�l+`�G@A��k��yB���m��.��K,K05sS�]]$ �Z�L�A�WY�_n�KJC�xe��ek|�!�8�1�Y&��0�hO.���sM5�}�P�n
gki��';=�KqV�Z�oRf��uq�emd�ň���J�3�p��@���z(���@��0���{�/NU�T>.P�le���ǆnǼ��&H辇�ԗ�(|k�ކk �޾�W��.��6vlW���Wz�ڽaF�)旗���ѧp⹆��Q_yK�d�wu��j�oH���:���^v��z^���;��`h+�[�駟����߉�KEt��O��#ٽC����*٨��q4I�K�;MIY#�7�.c6�e`ۈ�xp_�ӄ��JQyw��S�p�PޟgMq�0�}e��33���P�}��2�Dw^R�~9�s ����+_i�'92X"��l.�	���O$2.�z}��$���_9����ܵ�ǁ��sk����>g�l�������o�3w:	��:������N����ζ��K����dt�3Ʒ;p�	9o�VM|�D��\r�D!��|f����O�3}�|��9�P��$��ap��!@wZ�Ϸ����c{�����0�q]@��vY�>������Qڢ�@�gA�����>��K�p��坅t�;Z���{QKm����1��"UF�n4�Z0��+(3�'g ����n�`S��17�������x0<)έҫ�:�z�Kڴ�]B ;/3��h�J�®��d��Q�r �`o��-���D������4ޫاl�_�
�2���x\T�!uRӚfC���ა�cݒQ��w��F{�y 9 ��K5,ۭ��|�QeI�3�@H�g��T�����-����'���H�|r���{]ٻ�b7ю�N�N��7*x��Ȁ�1�.tA�\f�������U<rw�&.��f�<�$����q����gT��b�L�Kd�j ��`�P+�/OV��qz�xg|��2�/i����|j6��l�7����r����@��Y���p�KSpH�P<ҕq�g��O��(��h��Xpg��k�MC�m_I����'���}���2W��n�]DU��tL���w�������|X���4/��Xk���!������Y�>����f�>��V�A�f��:�Ԣ�I����ݢ'l��?vVE�9�
���gUXc��]wB�����r��Z{�ge(�j~ȃ_s���c����ꊐ���Va������y~�ir�<�ʬ/#�o{H'�=����{��Nϣ�hm���]��('���d��Z��^�c1{ɟ�,C�����pVfU�����]J|�44��-Z��>U�:���d~+���;�K�2�A��4���Ƀ|9f	ٹ�f�l���j!��z����u�d͔��c|ޫ�ć��utA��cF��/i�l�C(�(	�JҮ�������yxy\��P���h�ʍ�n�ҁ�Ov۶==T�|�p�>ު�+ѝ��}ެ��]Z'N���98����a�
�O�j������E�(�~��\s�+�
"_V��wz�7g�m��N�N�=��o�B�ϫ�$��@<�3��ENQ�t�%7��T1�]K��K�|VDWz�7���3��n��]"��cz�/2���G�����@3����#qNC*�&�+�c�����^�Ǎ��BF��pݼ��UTK�������AV���hʦ.*e#uS�?]HA\a�~~�u;.�y��>T�#��~RB·��is�A�,��������*�te�qS(.>�;[�F_l:��~��(�ފ3�{k�i�wI�;�Π;Ob���|;�i�%��@	�D�~�
��vrZ,>��IS����A����-��(M���G��qZs�N�ιuճV��O "�/x��r�P4ly�d{:ǜO}�P(7,W���gCR��0:��/�s	��Ϊ�4.���lQu�۸��0�g�H�t	d�4%��툀x*��nC��W���g���q/��~�A��W��$57�9��;����T�yx��Ruvqт���۫����Lv�{S9�f�In���h,<i�րǬRd�:�Ɏ���AL��2����;+�.��ʘui�������J������v��`�����_<�.����4_\���Qk]�K���h_#6���+��L>��H׫�i�k�U�Ŧ��{ݻ捻�ߘW@��/��cB��ĭ@��7|�=p�}u�5�2O�h����6U�<:g/�
+D�~=���G{c�7��W�����C..��`�zo������'w%eCS"��w�k�����V�]CI�ic���{��N�T��trf�z�(�
F,������-{��=���7�R�q/	�xy��ڇ���{��)q�uW	^���+������?�Bw�}�NK��6Gs�,:����T��	���d�+ݷ:��ל}�5�U}�p��3U[�99]���w'�~��˯����d���3���u�7N@�q����;@��u�J�7-]���[t�����{;���|�i�{t��ωJ���;P� 5�#�:��Ig��:gֳ֧�Xz��y�s���c�����и�{r��D�Hh����s*���s�r�q��P��
�F��W�V.!d�{���g���/-᳒]��J'@_F��&��F����^������N��^���6j�䠁�H���dMiv\L��b=|�h�
��-��Z��W[��F�)\"��[r�Q]���ӥCq˶�>�DU�k�v���voe�툙�ᙑA7%��;�ǵ zu����#-Y��V��y�Li�8HT4�v=�Wr���{R���v�6��%N�OOah�����U�­Kd�:�y7��{r��j���"SZ���'����va;r�N�dJ!91]���Gu�8
kj�;3/���"B#�͖�ݼR��Z�͛�z6�{��w
�k4�YQ��g��'c+%#a[�����6ʙՙ"NR��5VJ<�(K��%�L/\��x��Ce�(6E��*��Z�����Q���:�][K��ԛ�5��ys,���U]�xm���E �jB�`�Mۭ@D;�Mm�\ڛ�.�;
s���5m��ᱮ{���i�ݓ{�k�XO�v�������r&7k/r�F-tj�X���r��A�Gl_
J�����ú���6[�
DqL��Z��j���]Z�)pܼ�5j�fP���&R��#<�1a�$?hT�]f�էnh�%!��t��8��F��&=�؜�6�t�V^��-��Q����Xiۈ�1���^�nB[ޙ�k)0���m��́Ӯ��j�Υ�p�2�n:`�n�J)�&�� ��(�'\��*#G*D���_+Ϻ����"�g�����N��ۄ�@ı��<��F��q�)ރ�;����N�vS���)����ݔ�*�6>u�ZZi����zs�1gP+%ʜ��_*�W)����,��VXWe�2e����B/]���l�X���x:��ƻ����1��X�� �����d����!6�fѣ۶E�p?��̥8�d�wF�G�By�iR.��4p:]u�[��ㅊ�r�ݘ
M��vGP��a;|�U���Q<��\Ϳ��\�v�^M;�ΓC�A;�
��gn�efhy:���j���C�
;�݋�\�
��Mmm�J��%��s߇'��0���<�:�Yۏ�q�m��\�wz���|e㍨�eG��!��r���,
��v�v�2��8�X�|7�R�����&�ը���z�y�4��D�o�NSǄ\�m+uj9�0n����ck%�F�f��W�`tޭ��J�PS*�p0i�ј�!t	&ܤn��;�D�6�Kb��OUȌ��h�M�����ʊ.�lۻ�4�رbQ�p��c��'�Wl�`��x��k���q�r"�}��VhJQ���^!齈����3M���0D啓��=��ًu�f厸����q��R[�oDb���U���/�3eo-�;���6�Z�󫛑��V�4(�c�å�W�Պ<+��]�z�c[J��"{M���/1]Y���mj�F:��w)[JV��|��E�oz�ϝq��_
�P$ �x��so�nm]����î�F�5�g���x�x��snW4�^<��o%��5�[�.[��t��[��u��W����ȼXh۞4�������\ۺ�[��ۖ���ۘ��Aw��x9S�<ם��9r��\
*���6(�)$���u�-���r5˜��c�,E���7���%�����!x��Pj 5��Ic\����Һ�&wGyۥ�-�J�-�k.��ۺ�ts�w]�t�FFX�`ъ1`12'���Px�љ�^q\��A�]�,��x�<�wX"J۲Gu����ƌ���9E@|4( ( E 8��ǀ���꣥�W�XՖ�u�t�
��wR�v����uG�R⭋���k�-au�����g{yK����NN�շ��=�"�{&$��v��3q��a�O��v�gn;��D����l��u�ܽB�qso���p�t���hNbIO�c�n�M�v�B{����w��'�m�i��]0(S?��g�1^��ǹ� 'Pd����k���yu����lx����q�i�p�_l�[�Qrz����'M��qW�:��n� h�+�ED����L5Q[�x'�b�)1���|y��Q�CJ�J`�2{��@���z(����d���#L���n(�9S�^����}��v�+FyD��/����p�����p;��`���۪�T�<�i�ml/��*�J�>5�G��
��Q�=��^\sn����L���z��Q���FC�W'4�fl�����z�]`g1�:|���EvSy/F+���j�c��+��{������]�=�p_S�=ǣTX����%p2�u�Oa�qNp���Pꈼ��cЕv�=����h�G;�߈��+ѫ7s<�Ϻ\V���]x�7��fc�	�!ҵ��NrV'����˰,z~v�2�WP*�ٕ���ރeǢ�d;;��Y���X5*0�D�GF�:`绬2���#���5�Z�Mn]��Ɯ��P*�t].�c,S�2�.B����W*ԋ�����h�z:+��p��+�|������E5嘝l[]:�&��+Og,��8Xޱ����Ϸ��j���X.;}�#<��N��x�U��Xn(�%8�����b_���I�Q<@ڢ;���z%�j_zpj]��~��{�y�>%vYZ�m!;�}���q�	x̋����\�jt�Ϣ�Bg}O�3}�|�s����RIX�jf;.�ϱ�J����K�S=��t����W��
�'e�����+��s���X�X n�>\�^@�Vz�H<��b�*U!qU<��2������:���,�q���特s�|�=��^%��|�U��x��#�8�ƙ�K@΁ �H�=-���z��	�^��g;b� �C�ޡZ����fԏ�)	�o��;�7*x�"tf6�[�*��6<8{җl��Og�CH�3�=ԗ���8���i7�gT�����*�UOK s��2[����K� F��z�,���0�w�aq���Q��}m��i�9ӕ��wu��^�W���q
��8��bF���޽����2lWEKgxf���P�}&�}<�����!��)�{���c��^f�V(��o���C����(������pg:��~q�o33��[��8j�� L��FF�u�^ݻ�%�0⡖�[��pk=MoV��Ζ����I�bQ���]Vԥ����=5w�tj�ZQg.�d-C���1�5����g��Q�#��.u�Ұ��d�;�$=m]ы�}f�����b����v�G(Irr�g�'���� R^�EQ�[v�R�+"Y��ђ�uUÎ�Q�wlFu�'D�徻/m*hd����@������B�td�EH{B'0�?NY�x{vX����BrТ*��z�w��\�v�=>���}�C�'c�hm��z����|9�0���r)�]���ʽޮ۫px�4z4�5y{hzUS�}��3�uFv��z�NzV�Ӿ��]��Ӗ`���y�g��]��"��L��Gp�9\w����%:�>��Fo�5�񿳧�S��&<�P^�N����p���|=_	�
�]���r��P�p*#WZ����=u��,q�r'��Ѝ�V�z��'�D|��Lߨ�=�eň:X�y�!�d��� ��c��Mw����Kܯm�#�O���k�z�|�$�3�*X��2����	�"�Bр��Z�p�>�$���&��r��}�D=��c���R6�Y؆Q%����t��ac�ޫW�9D_���&�������(���ǝ���{;3�pm�;�-��ީ��F� �U�J�M�ѭ���re����n��te�����n)���{RNXm�{�p�ɞP�;�D(2��O':�eД��lӚ��z�Eշk�y��sV����³[s�;|}���gP��;Hˇ�|;Ѧp�q@	��)9�x�G��iV_A����z���}�\M�v��9�i�n;:�e�ճW��<q��C^ѻ>=8Y�D�0T
��r�zz|�t5/���i����{��s��їW��sӾͽ��E9�C���p��o�
�4.���<�ԇ�ھ�G��7ъd�����f�]�N��P���
���4:d���J�#^���-d�9f�_O����e=IR�- �r9��K�xr�n0
��뀺����<�������}E���M�*��E�Ӿ螏I�;��z;�]���upy|��ˎC..��`�zo�p���_Ƥs�'ﷴ]�����g��/O�JÞ��y	u�>��I���\'}�Cmu���z�(��xk����Y�)yb4�r=��q�c.*^��
�QY[A��+�"���_D���U�~�U�Vg��3�_Ǟ�5��/�L�����y�"^�,�[8#�����w�n�=��O�����׈ۍ�{u©����˩h�#%7B���ЬX��+��d&�"�}J�U�09�����b�8曗oc�4ЫW��E�Z�{�[\�i��kG�i+бn�-��0�P�3�+���|O;9+��c)9��twu^Ao8�yt駫�s�:hT*O,;���οUi�};'w�f;�q.+�Xn���%��,v���6�j����Ff>�-[��9�:]kr�3OvJ9��>��R�3ƌ�C��n)�'9Gt�~��Rҍ�(�bC聮���u'�Y��)�C���������/\�J5Z4eT=�S$`���B�Y���z(�f�ɔ�갰�{�*ٖ��藖���g$�r�%R�͇��K�νԲ��;ኣ�S=�=K���37��Dr����l�v��WGO����eZ�=��^��3��6v ���@�sS)��"۬��	�Rӌ�:sG�:��k9�W^��D�G]�^*x� '�@ـ[ +���,m}�ף����lV�^�����9�^�����|��I�θ�7�}qV�jY�D���.�������Q@m�s3g��93��d��[��D��8�&�����z*��t��2KF�d���F��7�B�z�z���(�5]���&;a5}&�u {��ܙ������U]�?v.��H��E��MB��+ׇ^�I]��r��� �y[Z­z��3��ͻ�)�q�m=I3YO�m�u�3�睋ڻ7�'��K&D���n�)Kz/+\p�v|�n�.�/�VW*��4w`��wH�i�}j�S�B��;��sV�c�^��gr[:���ݭ'Q������j���9\L���{��Pˍ�B��kX��Yn��斨�o���:C�O��ς���K����د�ں��c讓que��8���=��bR+|'�+��C����H����Ч�9���9^���VU\8�9Wo�qx!Q�S=э��c6z7��������Ug#zA9��,�a�W���S�.2���:��9|�
�e�j��w���W����z}�oM�9ʰvߪG���N�#�1�!ⴰ�w�	��W�\�Ow�֢x�/�0��Ցq�.#�.�cS���/D.�B�m�u�X�L��T֝f9G�����F�,�itT��2����:�:\g�S�L\f�����u�PE)��jw.���d��L�PN�詖�.�����x]@����z����\�9쌶5�w�{����׍����;���H+`΁0E���T����~�4���࣐�c3�ǲ��Wu��̶�dqÝ�p��]g�F��Ͳ�.�3�O�
D��Kf���z����W�V����ʾG\F�]�yd1�ܾ��`��.�bχ!��7�b�d��+�Z��eH��Z�T�X@ڲ���2pk̙ph�,�]-¹,�F�U��z^�+t:�B­틇I�P�]����6�O1� �n�0\rs=��uؤ��Js���4�t|��eoH������@ܩ�l�	���0[�*��&�t[��sԶE篧(.�5�R{�>Wn�y|^W#�գI��ΩuݱW���� s�$i�$tfc�ٳ1������q7}���U�0��yi�v�[dq�=���`7�נ\uW�պ�����c	ۓ=�ѳ�O���۰/�zx����W/N�@/�G���m��6�y��3�'��=���s����kW��Nl�����d�W�ڰx�]+a~;�$7ڻ��o��ƪ*��Х(2���'Kp��V}��i��5b�|�xuH���"ľ�ȴ��*�z���U���g���5���P�g��u��֨)������Ea��ʁ[޳#���Cxد����1��QM�u�^Tu.ݺp9	�m���ꧧ����uX���wM��{=Cލ��@>�̘}�&*EU�\�O�/p�xN_����T��:�p�>�����6;�Y'N	Ù"�sF �x�fb3=�����;�Ua�:�F����;b$�� �=�wZ����>He�\�ʱ? gm�?Z�[�S;����^U��6�-�=�8�X5�խ�#M�7�[Q��e\&�Q�Z�]�v���wř,R�u;f��q����7-q�YZ��<�!U54w-03�X�����Κ�uǛͺ	Q�'Q��f���e��y�h�{�����ؖ�T��u�KGJk����~�a`*�j�\`{�}o�����;������D���޽f/�on���|JVe�T@3�����n��U�MV1��c�9 �z��{�$�炼�Qފ�C��.���n���(Pf9�ʦ.*e#uS�6V���?{ճ5�����HΈ�N�;A||�h���lv�>��m�Ik�F���C���H���϶�ο�=�d�	��P�_q�9<�}�u�{�����ލ3��r N}��]=j�g��/�tm@���d^���C�N�>.s�ӑ�'�vu�ˎ��k�������1U����{��P�=�F�S lwL_J�zk�kC����x���9�9v���T�?�o⃦���ѩ6c�ER���Ƥ��թ��TC|P��x����HX����l�����3��F�ճe��Ww��֒����������]F��_�hDƽ��Qk&�%��W�*p�����fN�<E��U#�:�{��x�*<C���]u�r�y��QR��D�mY{1w����b���)b���J�<���k���j8=8jnct�3��E�ԡ�i�����뢨��Ș�\|_�(U�ע�xR�2�f`�L;+N��F�sW���l�x��M�s>ۺv�Xo,�A��oTmRH���G����@3{1�]W�i�Ɍ��o�m�Ѹ����_���2W�(?��O���]8b��o����.�X���k0��w
��=�=WP�.�G�c��ߺ�ﻮ��.��7���m�F�8�s|�kT��Ȣ�����
�FI�	��|P�����Ҿ�-��o}�U�T�l�Bcl�����Қ�Vg�����x>7�p� �}��
�d�w�M��@.���{%�H�Ë�\�F��f��ѝ���x�7��������՛ְ�u��N���;�3���q^��,�����a��j^�;�Y�����N�~�螮}/+��4�;����HвR�3ƾ�;P�=���8=Mi9����b����!�:��.鬾�9OR5K�B��{rID��{O����7�7ns6ϔ
��g�n(�	�%�z�\,��w���O����yh8��.�GeEwRǎ�=�N@���P�Q�2�b���L�2��F7}���O���%����� �ݎ-���s��Z��
��}N	e@v��~
P471$�ӱm�	�Ӯ����|{�W%���{�5�NV*:�*(6ɭ�ങŜ�}\�Xۢ���{���7:Z:�:��{fu�ҨA��sC&�F=(�G���3���V�t�:e�l�(�cuxf��n'�������n�#��o�� ǐ,vOn�owP�/�:H���H�|�Ac�kw���?|;*x��	���d
;+�ׁck�.��[��K���k���C��'9��V��wV�7�q:n:�*��Գ" 5P$tȸ���%t���]�U/C�3�3�}�->vǺz�=�3�����6:�ފ��U�6��Ѹ$i�]�w�O�'ym�e���+U���bF��&���>�@��� 3��`���۪�T��zs���_��}��{�vE�y=zlTN�`���r�㑛�p���7r��=� g12<�;_�;��Eyn��έ��j�W	#�k�WO��
4�yR��y\*�^�~�~�]v�{Et���r�Tlmg�[�׳\�=�rwC.��Ʋ	[�ن�ᕁ�Oa�t�	ˌ�:�����=��I����x���u8ղ1OgMq������Ug7��pf9T	�0���v)���6��R���X��W�ۧ�y�@�U�{�뷧x������Go��g��ղw}G�W�r�QW�R�*moܤ��Z��On��/	ی� ����.WR��{/�r7]����5���Y%Ơ�sW%� �
1�㐡�c67|'QؘU8��%����<u��M�q�S.�mwRu��0�M�%�񅃭���~v:	�µ;��q7M�ڛA��+x���Մ�X����}��ӎ=p��3��G
K�tu�8����z�%���K۾×���@iv�u�����T��un�;���Z[ʻ����Vi�h�upX�9"���brŗo��*�>*�<ܹՆ���e�F-�Qz{SC	H��w)w{u�[Dn�k��RC3���l��P=*+�z�4�� /n4m|��.���X�ST3�p�svc�/�7V��:�v�VurBg-����I.%j\���	�9��˳�JO���{غ1��>׎ưD�����获���ͩ�=�YE���q����=C�8Ol��p��e���^�s�T�;��t!�
Q��z]�j�B��]6Ăe�$����P!�yS�X�6���UqVN�� T4~S��"7����L�:�6���Yp��;^+.�{�^�*=u\��}v˚��쏷&q9,6�M�a�u��e��Ha�W��ujMm����ґ�ɫ��D���W;v�[�t�1�"Qs�wxk~s� �0%Q�<�q�;�T�T�X�k(]H/w�Y����8�y�����:�r�bb:���y�0TF�Y��5ţ��}��v�BVS�1�M�-�D3�.Gzܔ0�'V�f�����VA�Bփ;��ͮ��ʶ����c�:�\"�F�W�Iͫ�s
��}��A�Rs_j肙�^t@����֭Zd�$w
᫏ui���/�����.vd\�t��;��\Z��B3�����] ��w[�æ����w���0s��mŷsyi	ؗGdq������;H�q8e�IL�����������"�A�>S3eBo\ڃ��z|AmS����]#Q�W�;kK��ٰ<�C]����[�hb��eMu��_���v]v�l}tj}��p�t^u�_s$3k�i���F�L-܋��rR����J�{��_+����rA\�j}}B��Cz�u�s���0��&Sj�u�ڵ��V��7D�ޤS��Ւ��S������]�me��vTI-9�;���@a��Ob��;���$�������뭃�cʐxG�-���!؊�P��^�5��0���CN��FR���zgg`M즴��d�g�b��v:˫hmS�N�	��ewGm\-�:��I�8�w�.�n���c��Nv1�=ڈ;Dֽs��6Э4,��^�pZ񘼷�),�{�{���c��Z����P�a���9��{!�����fP΃y�m2��s/vv��ȍ��kwۍ�������ݕu��_B��N6{gj)!�M���s+����r[]�Jb�����GS��b=���rh�۬E�l���j�j��>,ՂP��\�ʳ��`�w�֋5��ra]�;EΧ���UP��ur���wt�eΝ۲�%�0�4���bA�$�S"�#4���bhy�ݮ<�ʓly�ƊJM16��#)np������$%�WK1�(�']$�';��1cL��df��C���;D�咊H
���&u���]�I;�C�����p�\�2"�RX��I���!��˩��<��i/:�Ε�g8���aD�	�ۥ�"�H-��L���Q���s�0��3�匄W�tƼm͊�.�ŉ3��vx�<똹t�׊��&�#�ɔ��h�
4.T��d�QI4���D�ba
 P ������:孂��h)�Ѝ`�
����"F�hX7�׋#�3��0���"ȩÜ�O�=��5��t̥g@�8�r5�n��`�k��r��Ѽ=W�Q���2�8���o<�7f.�t�}���sI�m�xuQB��_D�_	�qS<�.�����<U�P+�'e��ﻧ��M>��)�����!uq4�}�kzV�I�_��,_�*������[�o�}�=1|q����Ș�{�=��"���v�|�;l9Y�Xmhx�׌�D�=��?Kf���E��m��;r�VZ���(��#�W+���\���w�P�}}q��<o�D��l	��@v!3��r�]�ib�V�O{�`F�֛���My���wV�'��Fo�wlU���� �����5�C�(���/��-��(���\�Z�D���(:�?��~�?|s�Ők��@����iO�j}�M)���v{����t��茩8���6~	�u/N���yi�vھ���'��q=�[�W�YF�R�}�3i�`~��w��\��3�!�V*"\��t�5q����������(ޮ��O��2�^ƮB�wƏ'*���FF� yw���1�D���2)�a��c;�s����f��U�[���뒼3W]��h��sR���ƝFe��QpocY®���»�mֈ|�M�O8b7��RB�`�9�VƏU֝Y��P���yq��$��jC{{+�TV�L.�F.,p�ō]�yR V�Y�NS�M�ֶVoq�whnJ^"�!����t/����O w��6w�r#��td�D=Ȝ�/�a�|�����.3�h�w��ո���V��t�BUON>��_��ӳ�df��z���	��G��wY�e�����7�}Ig�'���em8�'�xM��Ѽw�xN����;�}'��=�@����՗.L��������g���c�̔k��YΣ������oGw�3c��'G���c�d�i=:z9ϲ����ִ�b��->k�8%?!����9��H�Z�Dj�>]�飻6w�qB��仨�s��b�9��>��R���Ζ.�y�!��G+��w&���W�s�=���O@�sЯ}�O���ԇ/|]b0��WI���k�*�����Bw�Ee�4=|���t&�XWRC�;��=��v�o���>��R�}R��2�.�3 m�e
��[o2��jz=�g��L�L�-��ҥ}Ǚ<�=���تF[����p��i��~��B�_A��=%0T
��3 ���E�ˉ�N�!�qX{����둔ؚΓ������;�;��нy��eU���Y��K�h����tS��$鉸����u��u�(9X��*r�+U���ׂU��d	[�j�^}x�Ufov���q���1,�a��"X�_q
��JC1[�NR���u;���z�k&r�ٷ�:S���bAa�O~���T=�A���
���>[:}I�=�Ͻ�)���S���oE���{�N�v���4.UK7
���� l�h{�s�s�^[rg�zlys�K�J�{@���-�,�:g�K���_>�\S�=G�\	�����tZɪ^����釋�g����	�޲4[�w"�M�����������������$�Ƽv����'�l�k8�Y���a�#�qV!����HןPn;����fhg!ꀺl���R��^5*������`v�����;���Q�=�C��������}�����9��Cf��)�F�Z���^�ъ	�\� Q����pv�z�e�T�'��q��ۇ�S]�<�Eo*����|.jG%���s;�'��_��_�����'�Y���t��Ȟ?���K��m�Prxi1�����\�{�"	��+o�C�;���+��9�~ɂEC+�����uf�t�K�r���{2�Y^>�n����Gg[\�'��\�^WW�i�v��n�أd�W��exΠ�{�U#�~p��v��Jξ��v�B��5�w��1i�&�l�]e:�k�;�nS<c���;śf]�NM��%U�����]vt�X�ԏs�g��E���Z�̦�>��
x�#E[ڻ=��р�\�u�2�A���;�*�'CK�Nĭ�k�{ל��z�N�?�������TW^N�t�}��/Eu��z%�}�nB��$�d�ffio���e����<gj=DQ��C���(j�=V.IG���qܦy�/աj�]`zݣ5����z�ޜ��`5P�*e������3,��w�}�O���s×p"��p5缓Q�u��^�4�|6pO ��:�(���S�؋n�M�v���Jۍ����P�����݌�s��o��'.:�ه�;	��l��vW)�@,o,����WV�!�ɜ;�E$d��c���<{�ln}�[��vu��ꮨ�u5,� 5�$WT���=jb��Y����j�5�c_G��Go�����ގ3�����6:�ފ.d�}��%iYN�{eߵ����;kҢxY胻^�!��Ɏf��MC�m_I�}ԁ�q���k �޾���@Uꍮ��[5�#�T��d��9*�N)�������!�j�eq2Twu�/�{�y�s�^�r�K�_�~�y�!�;�Y�����#�l_Ժ�U�d�5��p����f.�"k���u���Yo�#���N`9�U|��uլ�T'gl�!Mn�i����CjQ���T�Ӱr�6�#Zu��l��Iж�/�8�v �)�� �u�]F���W:f�woV�Wo�z�͗�K�8���V�{��Q̒�a:yh�ͼ�Hd�=��Ҡ��C/z������X�{~k���rV.����2�b��:)�*�U�(�a��=�{���o�5�w���������@1ʄ���^��}K��N�qhLT�ڭ�pG`5�P��ym�T��-�c�ޚ��3��/���\�}9'3~3㏕������MێǞttOD�V����@��pJ��[=�Z�v�Ӓu�$NX����Y�̂�����'�I�=u�&�/Ib>�VX�Q���.�ؗ#�"��~4�"�֍�lS����_�`�-��(u����aP���*g��Ӑ�Dx��P=�����{	�h�'�ϛ��:Ď�>﫪�ǫ�m9Zi�D���l�"��J�&O';nh2�-��;���D�f)Q�Q2_���l:c=�Y��w��sX!������_� r1q=-�2Mk���k�Go�Uu�}o��E���3���Ge!8m���{�R+�DU���N�7�����p}|��Q��_^���-Z
 ��Gr;�3M���#o*���S��q����F�P�Fh��պD�V�δ�F+]LfV�X� �2�Ld|Ap�͝�B��@6T� gk��w�
�DLn���Z��b�{:�L�j.�q�Yt�>��9L�X�w�u�;�劕��]]��y���W@-�\�e�V���Q�W* ,�0�^����z�a鯼�����g��[<}>~�덋�79��u�~t��r+��wUT�
Ij@6N���Xxg�ƣ�MC����Ȟ>S��k�����J�[�z�Q�d��k ���jy[����O����ŉL���ߍn�֋\i�j2���;ִyQ���Y�=;��FED>��.�u�c����)�a������X�����#z�\���᣻��(��f���ۈ]qXn7�*.��*�0����]���T�y�G_�Vg�����Sz��e2~��?t�2��c�g��45w�EoH']ؗ�|�r����⧄}q6~�AZp���6�����B����nx.>�:���go�x���l�J�����5���]RW|�AÔ&_Ð�+K��H���;�� {�}[���QZ*��g�X�-�P�=|���>ʝ	��ؙ���Ю*z��r9M�a`L,w �å�+��1����s�$��0:^�e�Ew�3{�_o���P�;���i�K���|����<z����B�������Sk����[.� �Gݎ�=ݰ��φu
#��j&|�?�*YU��Ն�+;M�x�ՁK/J$��t8K=�PWW�Y9nS�0h���*P�ϧn�Յq�k�9{�8�k���$�=8%��v�cR�ʜ�c�Է���dn��%p�p{��	�wS��u!�Ŭ�)���R:I���:�,�.;/|�z�9�38���ʐ����������=��c��:�A������I�5Vq�����*N�w�����h]�F{��L�\}����Wq�ry��3��qت1���W���Y�\��<v�y��� �:�:`H�H�Ҹ�-v\Mçh\'9�i��8w��Q�ɃgVw�v�Su�~��kǾ�8'��!_L����@�a�oV���ً=ܺ
�/6�e�1�v�\���'7��uU,�"T$��f���;�=��mu�:���zrg������Ǡ�+<x��v#�� WϽ�r�M���?k��.�CD�,����+�g�k�t:��ȍZ�F���'��x�D3q�T>���]��7�2O"���j��&Ur�.�]�tt�ւ5��~;��lzut|�*;����Ϲ���t�QTG_����XGL��hf�9>q]Y�C��~��|��%�h����QH3�G�E����wSX�<��s�+�'��^'�q��������h4�/ry��˴MZn��t��.����җ-����3�y7D��}|�ɉ�U5��Cg;ý��?������R~�"�ٲ��WY[7;F�²u/�}�:�U|�	Z�̼Twڳ5P��?�+�wPɛ�n�(���C���u�$�'��qW�P�䦻o��wb���,���Xɸ������^y�+����O2��.��Fo��At�'(�MܬIe��<�%>]�����C���p.;����7�a��[����x_�ʃ����c�mS{9 ���+.�𗒀�;@��뀢]w�3O��i�׷(�"ωT;)��-n���8.�Z��y�@��S:z�@�qP¡����:]�Y�_S�քm�<�.;�܅�>Ǳ�^`y���6 �$��I�j�:�/M�Q����=P��{�u�r��<5;t�쏨C�W,��~ٯ=c���jP$�tT;��F+鞭G֦���_a�O2���z�^�����8���Tnqu�{�g��	��$)@�@<�����RU�9��
�ݺyqsY���t�=b�5��9��;}����~�<\ �3����k_,�3U�4�r��鮡=�ք\���~�cr;�t��θ�7�u�̳�" 5_	G���I��<1T6V����������#\HQU,~�X��q��Ɖpg��`�f�?B�7~؋l`]�n��#�W��[�Q��zJ�S:�*�l�����I��_��:�7����rY7�JK�1׿`�&]κ,�:{����eX'9�����SL��%�D���4�W� М��ז�C�;c�t���Dq�M�uh�W�Zs۠?y�߂jR���#���������ݮ�q�,f|wV��ڮ��}ԁ�G�����'M���<��5ޗYo�^��\ͺ��:F=��IG�{7�l�-���;7c���<z2�}WmAZ/�>�->5M���x~|��_�O���b>��+���r��w��Z���-��ѭE)7���u��ޡ�+�����nVqS�p\Q�������ؽP���J!=�~{������>�<g;�'^R�{��bG�YhGE�[��>Q"�:3Ŭ���9�9X�·���<��-�gK����;k���r3ϫd��u�euGdȧܒÏ������*���񑨝ܮ O�+�+�q�=�ݕ�.�C� �hә�<�n�3w=w�ĝz�G�?��U�����z�:�z���I�K�L���7�Gu,M�z�愞��Yhv7[E}d"��aA:�*g�E�B��v�g����������Xl����P��(.�4�yܞ�]��R�{��(5��Z��n��װa����7p�
_�����TtsP�t�f��1�.�tl��`)��ksU�캝}����!�S̝L�d�h�����ܔe�6����}��7�t�;�s�V�[2O>��u��uGm�^�p�V�g�jH*����X�J�/���\ǟ�̓�YKf�{�af���W�R;�u1����;q��;}k;�tQ�t���:�<�wV��6���~fה��Tσt��H�O��]<��#:���)	�p���r�T" j��t�ޙ[�1~Pz=��h
���n(��{�Q;󦼇�/+�܎��q��#n:�إX'2JX�M���K\��ў�:g'�� �$�3��W�%3��0�ז�4��#��H��9X	~�^��N÷C�ӫ����[�V�	SԪ�<��N�H#�D�T�<3� �5Zj������]�+���롑�܅��ģ�gȞ��)�{�[�WQ���XڰY�43�;�5��q�z��lH\�;�ٶ���/���[��E�����j2+��<@�ޮ�h�*�b�%�^bjsU{�]ҫֆ,�(�F�f=�Ua������f�x�����*B�Y���=�V�䡵矟�a~7������hlt���o/����q�3}4��t��]� ʪ�y��w;��	�?��%@Vf�5��<�+��Mܩ�s �X�V	�h3X��{��YY|�,ogV�H.	��+�:*s/����,�Y���ؕ�	��n�Y�6��M;ת��:�Μ���T��GJ�ZU&�\������\�U�Ag>�ǈ���4+mȶ�R�N�L���oi.�[������E0��Ķ;�ʻuqTe0M�*������b�dT�����A�1��/��f�ɷb�R�:{t���ԨV�f�[J���\�����r��7��K�ݺ-&)v��ə� Oa�I�����n�e8�9�����y�;֖�׈�u1�����)�c�a�4
�b�\�^�p��v�98Q��0�{J4N��ƒe�YZ�V��`��]�"��lC{����`����^]�I7�+�sg8,x�b�u��M	�.�${��wJ ��b���[Y�o����w#�&�]��j�����-�f��ob��j� hR�p�{%-��9�����H�E�0��	�+3S#.|�]�&e>��񅋺�mu7���B���G�L^-']�g��"sn�i����A�{�z�^ѱ�Af�ܠ�3F���t�4���.�e�j����|C�(�F~a��4Gf�b���ׄ�0�!9�q�g}͇�-�ޑL�j�6�hP)�$�gХ,ff��XL�����+5[���"6�Sl�udmv��n���ˆS���jf:�����]�*M���(�ƾap���8�����@:��L���XEl�u]�@R)_f`|��z�H4�᭵���`���u�5E�n>jl�f���fM{͙2	����:�ݹa�������YH�o�1���Kkf��1���C���/�L�{���h=���Z�:WcC�F�6��R؅������rfVp��˵��;�_f�R�_�;���X��mv3�|
I1�����k-��r�wU� �O���Ǯ�X�"}�;������P+l�GV��{�W ��;��n�Ďz���[��K8]n0:,�\^EN����W2s�5��n�e����(��ֻW3��Ž'�F��4n_M���[r���ϊx�7t�7�O!��r�S�WYUղ6�v��r����Ë��ˬ�J��*�=��Ձ��i�����ݫ[ŭ��M�2:ٯ�yy��	��Z�(XyzUP�� N/o"j�.���\@�t����� ��2�4/�P��W#w5�z�=�+�����t��u�q��ɞO�9�9�ʎc]�z���:�������S{�,�Oz����N&o� 9N�;�%-G�8�A_[n�P��Ӵ�z�!�1ռ���Vs�r+X�)��n�"s���¨���:���}�򄽲x���ݮ�¢�>�m�X�ve�u`��Y��6�,�4Э��7(��*Q�/M�onc�ܞ2�B�S���*�m)�)�B�M��6�v����mp�@DU�)d2%ݹr�:�r�fE�\�7XA�s�J(�c�4$�RG:aD$E4�w��F�[�wIR�&�L�4��`"K�ٺDtb��݀�YA�;�.n��I�D�݋�30�I���h��u�H�&%��k���R.���e�$���s�N�B�w]:��F�#	wr"w;�.�n���#���b]�b�c��B�JB�������d5N����Hr���#��]�NWQ�Wa˜�Q,ɓ�����̗6�J���ff��LE��w'u���1�v��<��<<x��w��®w��ݻ��wt�y�x��x��;�Jo��0c�#����X��k����cR��tf�V-���՘��$WS5��}bs5%w��ej#�m��w+z�kZ9��.�y��M�8py�ϾǸʣ��U��?��e}g��_�U]������\%`��H�{U����nğ�>Z�94�_���t������^.����B����Ab��2H���]uo0d�{OF��m�^q���T�]�8s~����S�pK#��0$��dG��V]u���pd��w���Ou�/7�4����.�~�vD $��W�c ��������93��tL׼�VʱS�K�!o@�p}���O���认9x��Ey���PGI;==<���*����ݣ�R�:�|��a;ʐ�����<�K㞎ڇ���#�YH?�K9m0��<�m�V��X�ԁ�I�c`I���:̒��n`,U�w�ry��3��qت1�me�1>:z�m�nk̴,����Ht�I�!:R��:WZ츗.��Ns�Ӝ�G����\�U����U	|o�S�C��6�pO�pB,�6��Aߎ�ׄ¯~[��k�VԮ�7���~��P�L��{Hwt�q�q;�UƆC��e � l�+�h\S�㜉�Dv���ř�}GB�6A���D�O1Xʔp5��v��*����pF���*юX�,�#��zZ���N͵����T�F5P4��r���pR�h������n���W��C
��V'����<�k���o�w���o�iY�;�ݽ9�fr'���m����g��:g�M�wu������Y���!� E:<)��(}�습IE��ё���FOKU�Ŧ��_Ϻ�����3�����w��:�����=���[u���:���xa�N��i�*�o�Lz!�WF��5\�u�{�342�m���v�ܔ����<�P�wmyT�����Ar�4x~F�������G����9���3���Sf�s��7���\7C&n����XW'���q/	�a\j��p�x��c�6Ռ����p�+Z-3���}�U�W���l~�7�x�~�rp��g�'��~:/�s��ϧ��-����z�i�j������?C��pv��>ޚ�z��o����ɂE����>�}g�x������X:�r5A/t�9�3�,,v�+�zs����X5|�i�׷(�,����&�����F{+.���=z��+*�����+�
��
��wMg���/DWZ7���5ݻ�{�32{�vj�[��g�zzB���z$�5v��(�#Qp73�^@T,��wuGvʸ�KZ�׷5J6lBI����"[5շw#(WF��A7�+�կ�Z�vr�������s����'�.��zI^|�݌N��jړ�Pu���le#:��^���M0���}w�N.��ѫ�C�0ww|�F]����J�o����gj�})��)�/Kg���9�C�z�h�	+bg@�S�S)L\Uu&i�fv1���9+zOw�w��7�4u%�_Y�%�|�;}�q���D�������.*e.��ٟ�{������4OP�uֆ>޶�F�;}��r�}w�;�ʞ6���:��Ǹ2�d\h�m�x�"��@��\����rڴ=����Wݝq:o��qW���=*b�3b��׵ϫ0sV<�x����Z��a�܆5�vǢ:r��dq�OwN�^�	��P4i!08��u�{_]n�����q���*�ә���Q妡�|ھ���ύxp=}��㽻�8�Օ�M/k�73i�`~������j�$}�Pl����axVo�A��F�E	�Ⱥ�k���q��5����2u쁏����"����_�A�å��p[��ϲ^�lt:�>4��'ƻ4/J^��·�w&.=���t����e�P�oH%F{�+��À�OZ��O:�Z���}�N�����CЕ=�{P�q�3�����]x�#zA9C�����>�=/�r�nd
{2�TB��v�Pv�9�I�fs�)3-�+t����˽�X���3�9�v=���@%���^v@�4�rn��`��{R{(;���8���z�ǽZVФ�)֘�f�0\�ܭ�o�����es���fu]�7�n��r��A]�����afWy{l{�T��7]�;�GNϻ'�����컋޷7�;{'8�2;�����3&W����Jܦ ���|�_��{[�g���C��P�V�$��gᄗ���v����;s7e�:����Qp9��
�Ը�����f#["�Y��Zr^�{:o���[E_���e�T	����S�9M�����.�\^N������I=�QGh�wOq^��q���#q��4�l�X��*������)��wnݪ}j���������,{�J9�w;��g��Q��Y�Q%��/oB�U~���n{{���`���詞�qS<���.>���<��:��'�__\w�nT�޲6.��ܨ���>����%eG�3$�Õ���@?Oi��a��ꑖ5g��|&������J���+�j�e r@�����a��ݨj_[g��>��%C�/zz��yoouEі��N�m���TK�KSpH0RqR���|#^Zjz��E�;ו�A��<�&ve�f6Mn5":,��-I�����e�̖n�մ��C{@"��YY�0����ҺL���|�SoE
B\��zU7Ξ���&b����+o7ATj�lʁΚ�.Mtg�7��3��eg��C;��=���I�emR�$�G���g��%�5�S��'�m�f}��\���,J~]����|�M�L�tu_\�ӞQ=�=�Dm�+�1i��ǉ��&=�Y��ޮ�p�c����|��p��z���7����v�Ӹk2xebw���wt<�C�]��o/Z����_~:0w�����Ki9����z��;���7���荦0U����%�z}���Ma�ٯ�����t�j��cYK��}��*��h�̨����}E�8p.;y{lzUv|�P��/V�wVs��8����>�o�_ϽY'=��8r�"0�ss:r(�'+ݷ�=�i��ט����I=z@�z����C6���hg�x�b�ڧNؙ�-xb��m_?!���BO7�{���5��j'����o���D����Wz�7��Q�n��Y�)Y�= �c��V�b��7���z�!��	X�p}Mw�V_S�]Hr�u������4%2{F�RK��W�z�}���A����zn���I-���=�=�磶�r����#�u����XTwde&�Ȩ���P��餻z0-˟r��vD�z:Q���\��W�U�>�r���%�U&�V@~	4�o����|3{5�Xi���w�.�C�m&:S��7k0U�%'X�7uc_u�@���N�0V�\��u\bWX��ge��r��{Qv����΃?M�$��24D>��e�^S?ϭ�A�X���'��@xv�E�L�o������p���5�{�e�^�L�=p� ��D��7��qFQ|}�\M�����_LJ��Y�<s��Vr�����yt�;q��#/����8'�Âu l����
�/OT�5E@�w���s���.��D��{���z{�a+�θ������s3,� =P$�v��m9��f�t���˵ݔs�G�܎���`w*<x�d�wu����u�\���p�Hi���ʛ�49��Bx�fר��[ɫ����j���]r-�R'���3��7C�w�Ǝ��Z���m��ngl�ʏ��$�i%��i�8�b
7�<۫�~j����4�΃�����~����Şԩ�W�'�V���םK�c��;7P�a����4�gU�v7��F��7�O�g�c#����U�'�:]��3w�@j��p2p;��v�ny��c��^�<����d�-�{Z�]�����;������J�߿]
��o���/�N�(��{S��Gv�U�5����j�3?5x�F������iJԻ5�Дe���n��vB��Fu�sa��0���n���וu/��B ���n̝V�]�K�ʖ_'��JG#�{c3g]d��6mI����U��8\���6�FJ�t�"}@�ݨ(��u	Q��Ş��y���r�	�W��V�b��Ї�S�A�}{���\ug�ְ��8��߲`����j���g�����s�@��BQ�=Jxq��X�2%r�@��볥wO�iK����{r�X�v����X�e���":a8��{Ơ��+�uH�9��pW�Z�.鬾�9z����z�����D�����Q.�k[r�.Q%�KD�~�<��Qp7�L�X��J=ӑ�[��x�z�z�P��9��]����Z�V�~��	*�gb&>�3�"��s7NS3c��,`����%ݞ��(�>��K;q��;}]g����RAu�`)@�<�ñ{޼N`�W^���m��\�[��7��`���h�oH÷خ'-���ʞ6���|g@�D�On,k<���P{<@�;=�k��'z$\��}�����&�:�t�S��}5<T!��P{���oG��^�����o��/(
�������-�k|�GNV������K��a���Vw2x\�+/u��Q���ꪜ�$���Ԩ��3�&��MC��W�_t�{F��B
��ח2qgK�V�e*#uh�j!�l3f��R� ��C1�3t��c�_i)^9ߤ��z���V�]�=�n<�hZ�\�&v�tuv��1��5�����GTiK��]3˕]�q96E�)��h+r��q|�^ܬ��֙�oG�;�Bz��5�R~���uL\)�����}
O�m^o�����%>���}��ʏDk�Dɾ�7����<EB���S�7<���r������R��ȬR�r�ʪ�/�\��OFu��}�}���mu���z�+����sᕁ�Wt��b���Q�z�z��ud�;��C*"��ÂS�p�1���t���ÿ.�]x�����o������K�}��º�4e�ٔ�
������w���ޝ�#�e}����~��]��I<�˫�ߖfd���:�;�3�fL9�����e0�*�\��%�j]y�v�^�������k��Cߡ~��C>���NƓT`��/�a�X���8~���cv�b����ZKp�z���P��Ew\f��|����h����U̱hz&v)��E'0�h6�}';�H٬���Q\�����,�}�=�z+�� ���>����$�t�[�[��U�5�)������}U>�>�4�����Lg���;w;��C��a�O���$��{��?�<D�8Ѯi�5ZsT�h!n�<�as����s���XlfT�T�6<��G�?]����þ���YD����v9t�����b���Z,�Z־q:��2Գ���"u �éѳP�Rg���X]\,�VJW)˕ں���z�63i�����\=��[���P{ �3�u3�n"�x.���-�����<��:���Bp���{�w����\���Mt��D@ޣ1�$��+�=-�&�-Z
��w#���#XZ|����z�M��H�ww��UT��2 Nk�#L��|6_^�L=5�����K�l�'��|�}��йe�:�B}���B����\����W�aI-N��]HT�����I�� �RZ��o�/Y�'��;L�O"x�:g�K�q���{��U]F��F��񡕷:�Cq.g*�}7����g�w��l�5��D;�����}g��g�g11���<@��z���S��V�*���j�r'�ؾ�1�D����l�5y,f.�ۻ����q`c�n+�z`n�����w�WmwZ�Y �}�3`�ܮ��qE���c�c�����MaQ��q��uX����b�z��X���V/pO`�|2�*��A<��>5㘃�k�4/	�q�q����<��������P�����97�f��z��Y�~���9�P_��2rrii�{�p�#@y�$�,�
!S�e��X���@*���K^:v�Uy�kIz{��#���X�W\��r�^n���KE���	At#M��X�ò����ʋ������s%oW^ݐ�un-A���k#!^�Qs�N�%DR��t���������5*�V�Jp�L��D�V��wUFo��{��:}�:<�jt�g��d��*}G ށ��7y~�Yn&�K�����zħk�D����Wz�7��z�^sۤ}gĥcʍ��W��כ�Y�^�X��T[4:��3�q^2�� �&��+>���z�������*���fU)�>�_]��J ;$��1h��z�]L�7N@N�*B:�����×����NW�:��fzi��O=�Xl���T��$���l	-T9�K�	�E��+w�yNt�� �z��7��<|�tgK����{@	�}'@��A��Kf⌢���ˉݮ���a\�{ٱۤ�ViZz9I÷��#/����ӂxۂd����_��
�Z1�@u�f�]+�9צ����R���1���z{�a*;:�v��uU,ڂT$��{���>�c�;YY�+���dМ>���Q�!���r���tϸ��덁q��5�b#Z!��BG��T��W�̧F�ܚ�ɇ��B��	��ZfXp�<��6����V�������km����kmֶ����umk[o�Z�ֶ����ֶ�����m�����m�����m�����m��kkZ�|���m��ֵ��ڶ�����mk[o���ֶ�󵵭m��kkZ���ֵ����m�W�mmmo���km���
�2��<$p	c&� ���9�>�9�x�*)BJ�*�Q�U J���H��J�P%(�H�QBI��(J�R���UI$(J�D�D)P�EP������JN���
U"[eJ**���D�DJ�J�f��J��"�T��Fڐ�[�R��UF��T�H����$����QUH$A%
�B�! �������J��TR!��B�R�U*U
�T*��H���J���!#�  	�����d�@*���TѪ�J�0P�� Dʕ��f	��4*6�@ R�[k�v,���j�B�T(��U.�   ;��Uh(��Z���k
��c� �@wNn(��( �6��   袋:8�    wh�@QE��Q����Uâ����@{ڡBU
��T
*�V�  ��*�Uf�E(l����F2�kMV������ڊ��X
�[Cj������m��%�u��ZJ$%B�U"�P�W�  l��z ��65��ZF�(vݳ�����V�S�+Y�Xkn��T�Ҵ�k�d��YQ��u�"��j��P���0%"�"����i�UDo   3��V����+�Km��ݱp��i6��bƆ�c�i�U�Z�ڴ�@�fѶ�J�`ɛJV��e-l �mٮ-�J%!E+f�QR�J��   '��{j6��&���WJ�e0퀪bm)RkU�B��
��Z�4�h�M6[Cl:�C�v�*�j�л��8�n��
�RUJJIU�A)AQ��  �7���YT����6�m2�U�v�S�cm��0 4:��mm�!�ff֛��p��+N�rYt�6���B��c%�5P�a*AJD��  ;�^:[R����n�қc����]���j��5�kl��e�)��n�tR�+UX@뻻w)��T��mT��bڃb�kT)V�����HU+x  �{x��ι*���iY�tꃡeL�Aӡ���Z��q�v�N��i4�;n��JP�
��δ�0��vH��P�UIAv�R@�  �xV���w��VT����v �K�3Y����ӊ�%ٳf-�.Νm(�V�ӻr�����PR�̣
V�O 5O�&ʥ)   E=�	)I@ hE=4�MCL@�O��I��T��&*�h&F@	4�M�T� ؒ�aB#2k��$�f*
�m02TF�
�^߷��o��ˌo�k�BH@�w�!$ I0I����$��!$ I?�	!H�!@���I! ���3�P3����4�?�5 ���;����nݍ���hҬ���	Q��f]�){��h��6
7ͨ�i�卛��{�jl Qp5��b�RKf��@ʆY�ͬ�E`�ǔ��tK�fb%�-�n(Xæ�`!��Lf��XB#hId��3� �Ր��+������QR����7�M��aGtԅ��Mջ�ݱ#��&�2����Ƅwg/�O �p������QQ�QzwsE��F�N r��jae��Tt�fE�rP�H�¼��i��XHoZsāVי)4(i��6F�Y[w2Ņz�&Ii���/�B��{�K��^لjX۫������V�b,v��jlT:E��z�bf�D���1�(�R�&�6��-�R�\������7��٭Ԡ�1�\�wM[�ckaƖ�1�a�(]a�Ymmm%�3cmJc5Y�v ܼU���Q˲�I�C`�K5g6�l���52֌S���LJ�5gM�t�I�Nmϑ�oH 8U0���^��O1���I����nѭ��K�M�	'�V�H�mH�)�Vg��6��+4�[���$�*�{���{��g�H�FȕyH��夐�A�g&婎}�] 
�/l�DǬ�6Q�%��G�6J�YaPX.T�5��M�m�b�cM-+:��guQ�®+!R�g��I�d�`PTӷw����8�:9ĭ		[�+CX�a�uf�ڲ�ᙀ�C���P�[�[���B��8N�H�W��Fa�Nx�𝵳"x�Tı�j���v��G��cUL
QZ�5g.	��Sk^�t���d�sks�1k�
n;��lJq�Ԇᡩ�ǻYV,8�Al�:����X��ݸ�U���&A�+JU��F�1�ԩ�llTE4�T�Le��YR:�u(9Y��iT&+˂<�۫-aK31W8.Ruo�W!�a����/N�K �.���5��*����Wr5���*�,�f�H��r�f�J'Y�&��D��5�C72��qT&:b�Y���c�	LM�Z�{�r��9�0���GlEIV����vor��"x'�H�
[���8�r[��ҍq�{��-�6TQ;�L˼:"�aBʊ�U��C�i"�r�1�-����b�8XTˀ`�oj��n�Z[ړ�g�m�t���S,�B��2�V��J�Cz	gTw�	�u223GNn�e�qb�P��E`���֒������oj�ݣ#[n�b{�;��5�a
x^aÀVFn�Z�F3��Ma8��S0�����rC`e�V��Ub�V�]��ʡkT�D�L�-�!2b�h��p��/R�F��V�	�g����J(�i��
��*B�����AQ�E�1�&�3[���'R�Y�P�Faځ���b$ٕ3���q&����VDp-v�k	��օ�P�&�ѻ����ݍ	��BV�����2j����MjˉZŋ�-��*Kʋ��ga�I�H�]�ř�fL�2�j] ׃6�V�m�5,�G·uf�o���YR=�[�4�X�P[�U��Z9j1�>81֍"�Ea�����fB�+[�0��˗d�Mt�&���0 E����r�7VbǺ�jĘ�B.�E��.��@[xkj�E�2>�z/]e,�J�W*�U(��X�ieШ���,6m��2��fR���F t��Э���7k%Ә��`B�Ңۆ&�kJV������-U���w�,�Z.h*�ϖ���d�u�7F[Xڛ�*Q6v�d�7�|��2�V��Q���"
�!Em�d�Y�ۚ�7W2��M<X6.B���h�ҏ2�:�b
�c�S��U���k62u����zA���q��3�Σ���ne��E$qZH��V�1Y@���	�\ū2�bY@��tulڗ2  �f�-e�-;;l�����C�{��1���M#w�� J�+dU��<ϭvPI�xW}`ڤK^B��:ra����x�m�G#p��l��O��(Q�WKw%X��A专3d��G��-?^^0�ga� da���y�d�h+��)4�!a��60m�wi��4d��]�̛�A����{�����L�m�Q���iS�[)�)�-InJG��Vl��ʒ]�2i �]�ʂ�����d����ػo]]�s)�^`��bQ����V㲾�b�h�!(i�W)2X!�M��ΠH�c�Xn�Ù���xRցڑ�J�������tf�5�,�+)Ԥ�C�<�T[0�D7Aێ�(`�k0�im	�4%e���x�nͦ��1�4ǟ�v���U;�ҽ��_�d0�;��,]&�.-�3"%�wBVI̰fǌ^[�gp��w �5^cm�t�kb�y�m,�S.�d�ǳZ�-�Ż�1x����b�2���F���a�tX'wT���h�{i�&��XOJ:��L<v2(�9DX�U�2:4��L��飅f�LA���o&Mʻ�(F�b�*5u)�,[��1Z����1��0 �wk� _0r��]�Ӣr�0*;�Z��2�BU�����W4ꊐ�߳wF76�1�ej�D��(ʎ��U.��v���b�D�����15pm9Ic�`Nl#*�C�X�vk�6�*����� �QC4a+Y�N�*ִvƤ鬣���m��ɼ��Y�]<(e�[Y��]��v��
jb�tU�-�9F`�O� ��ೃu�n4Z�P�F�;XsN��- kEx�0�T!lLb���ۦ��4�[Z�W�*��+E�Oat���&%��4�;WY>��\�4��b����y�"��̀U�r5.�5�m͵)n|�
c�,n��xR��~���t��;*����oo��7��TAڹ�"��Z�%G�LK^��C:n� �q�́���I�ry>;&���⦑ג�a���WK
S����#f�N�Z�߱ڴ��4Cų����-V�2U���ş��$��Ɋ1�	y�q ;��}��V�謋2��&bkS8��bfC�2��I-�ɢv�3sB�Z%b���"��賬%&^� �!�)��ך���'�������qfYu��5xun�6!aڄf6���޺��` �p�p3o��0S��b����#gw/v�����f$H&��٘赣KR6��t��A������"XH�ݕx]<$- a[VjF��`�Ry���b���Q�zcCP��[՗���]-�,�C��bI,[��cL�12�֑�.����tD���VbҺ0+����eh0�X*eKbX�#�����:;�ln[�T�v��d+��X��3)^�t�RV�F�Ʌ#��V��6��YV&sf@�0sV�+FI���[[��טJ�=R�Y�t����/��Te��)�R_F�s-�2�\�"3c�ѵx�����)Yƶa�N�2�#��kV��Ϡ��j�:h�3�f\�j�M� Y��d�	����7	/w%A&���!�e]��(��򒹀ȲUӸ6��1%�.-/DVה�ks1�@ڽ�Lj������%y�����6l�ج��M2�Q��$ڻ����;�U��^&�R�Y"�-ÄX*��բ����6ƇK �[ {TCyc�P��d�.�/]U��P�@�ݬփ3F��Y�E��&��,I�*�9����7�a,�9+L�+[�8�B1��X1c�	�����RKa�O4d�n���	�~��r)�qcr�Lj�P��V6 �]^Ԥ�n���*̛)a��Z�Y
U��֫v>j^���ō�1$�aTRZ�V��v�2�
�=JJ�Q�h�N�.�����8�9N�$�ˬ�ҡR�$�����4M��o#����l�����"AQByk1��)�T�Ӕ��1!��w{���S�+]%�fk�\��M�j֡R7��"����>u(V�.�B��Yi�.�v�ĳ�M�jfѹ��'1R��YB���O���z䣒�ƍ��be�ZB�Udj�A�X���bHثe�oiV�r�x�Ǔo[�kS9
p��Z�\�;N�0����ǀ�B��	�a�E�!���c�F6�f�%��S4|��6�̤�%L�w��c���)P���5���I��&tݵ�A��12o`vrY*��V)SHm���jŻq���TH��5W�xM�R��X���R-�d��FF%"��n�Ca3^}sȩ����%7�ݧcJ/6��KYp���4O7���S ���у��Y'Y�i{h<IU�p�R�V]Vh$������*EpQ�r��Ҥ��O�j�u��һ��Wz)�6�U-���aګ��=`�4�{y��֛	�e�ix���$.�c
:a5З2�*�h�n�D�6N�[�V�j$R�M4���/t�X�u�r�@�m���r��6��޻4ڸ��+z �-;mɣ.R��`�32�T�)�/�n5k˫A��hP��'E�\iՕ��ћI@��u�a�L�*�k���2���������7O]ak���;�(@IH'ڲ�_;�!�`(ѭF�1C&�;k.A.�;!Xe�J�Nһ��k˭PL���h(2�ؐ�M串�e]Zݨ.�%���#�u
����C��{1���k�*�0Zi)��6�M�w�bkH����6�z�NV��v�6�]ake6Ƅҫ�9.;1nFn��Q�A:@1�� �*2��\.���@�T�p��*8ޫ��tr�l0��%�ԣJ�<��Z4-�����(�hJ���(�H^�S]�B���c�	�>�+uL�KnQxwn���i�E�昵���t#�gN���6�e廠��-�%��*�!������X5�sWN�xC��)��l�6�J��y���U��
ʛV�-����)���˲��j�E*��4���5��&�[��k4`�4h^��4�J�.-���<v���PsY"Cz���e�1(쭸��ڗ�2��/Sۧ�d��4L��p^:4�)�ş[s0=u�f�Z����ցJ�*d{�Cv�"V����M)A�j[�����X�l��
�X+Z���L��K/粮�2��Uر90%n#�Y�S�.S��Y�3+���7�m��.1wR��ڕtƒUF�����*�+�ʳ�e��*�>{������FeXak	svL4�	��Y5�3or���u��1��l�*n���\.Be��uG���{E��&Mi]��@xFf�w��V[��M�LM�O E�j��a䣕 6u�e�@U�iV�ܕ�AH5���m)�b���5�N�Ks���X��p�)�.���%̮0�n��6�5`)��1Ҙ�:r7����Z�C+Sw�Pۃ/F&�����t�̷�3bMDi��ۺZ:rԐe�c�[�D�q`DG�u���c`̂�6�C�4f�I=]h#l۠bC0�2&�����m�4�LɶD��ZC�L��b��U�m����AH�K��Ø�Jҋˣ�h3p�)�����ځ7y��Ry�e�P�u�"
�{Vm(��h��D&f8n,�%F7	�g�96�k	�ƚM��C�7�b1[�wf�v�KYu��� 7��Q�6�5K&����/�ç�A^��Li�zi�$,c��W�~Ö!�)���$!�Bu�H^U�h
�oJ��gN��N��qR��{,]
Col8,�wE�U��Ȧ�Ґ�ilơQ��;)�[E�s+*��k�%̧b>ӭ�&�WJV2�!&�I�y���rímE%z�*������l �d"��O+B1�y�oS��.�׌#Ie�n��8���xM���u����6���q=�Z�l�TfCg2�n]��z�V37�M��ԡI6�(Ś7��t	
 �>��8�C�.��>�f�t��^�wZ�[��$�Ѵ�Ӵ�]dЊ�#.!{�`���f�aS[�[hS�6Բ�ʨ��4&ի(*6ߝ�c�&�7o*'�f���R�&���B��L,���d=�����cx/XV��brb��������b�F�ڬy���{GZ6U�hlt�^]�l7�\u�r
��d��0���-�"�cd�w-����F�n���-JԨ^EwW��^�n�,�W��"�g57fa%�-�&5�Z��)�`nQ2��{Z��J���̬[ �RY6nv&���@ۧ�cűi��r3T�#���oiG� ����@�H��EѦ *�[�o@wR���z"h���Ze�O$�Г��$�1v�#4�5�`l��9.,���#6(j-&�35ݴ��ȞǑ#h����t�<Ӵ�
]\Wh�U�z�'�kf���B'��l*��GVrL
iaW�m-�x�#r�Ԡ�l� ��r���vS����S�S���j��LQ;�����j�-X�x�yJ�T�AMUeٚ���f�\@�.�,�S��J]��I���>�e���Ku�jX��,TMle^�yX�7�)�".T6�Ƞ�JE�j���Q3_��D�C3th���%��Y��(��й�y)���F�z����<�4�ǌ�;;�7�=�o-Ѧ��[n���QJҾ�]wGtm$X�U�Mwf���A<cQ��f:�RƤ5�:�ɑa����4�7v�,ųU��H͛2�;��I�I;�� �0ԙ�Hr���.�뷒I�1q���I&-0�[ ��vj�cRyh+4wM���{���R�%j��I(�J��.)�p�ۢ(i����;�4�Op]6�zib԰ᩐr8�/.Fqw���FN}�Xvoh������	}�\�����cޙvLEl.��:�#I�����eB��W˕F2�4�dN��fG׬B��RvR��gXi����+���jΣF���Ȍ��t��.V��]n�V97gf.r���:=���[K�NeJ0�ԧ�vֲs���ws��mVtTy��H��Ӭd�?���m���b���	[RWu��Gw-��ep�r��1k�z�+��P�v\��-Gѻ����*o�X�]C��pԴ�ٚ���\������-�n�2�f��A��\��5P���շG.�v�0a����A���q���s�r=�7\W�u��nm�Q������o�h��BVK���9��J̡ĉ��-�LW�79�KE�H���e����Ʋ���R��O���S�n���o]��p�q��n�;W��]@e)�c��=���{Ø��݃�]�v[�R#|�wY�\���2��;&Z�uvw��9��ud��LQU���۵�X�:�],Nq��t���-���f�跺=�w6��k0;:_-���R���NW;���7�[�T$�H��J���	`O�6�(�'�T��y�7��>�SG~ fi
"T��/va��j�n�\��-�Vŭ�:Z��qƎwmuJW����]��,��E��+=O6�l�F�V>4�q�\tk���;��$Bvq�z�"H��[��V���g�yLHV�����P���!E�Y����V�itzU&;4[��q���8��+v;���;jp��1�T��.e���uu[��޳�[X�P��"�&��n�N�n���h�pu���'���<'d�kh��wn̔_�a�sQ�6�J�NȮ�45�O�<]W�S�㛂�l��8���&�ߧ[p,f�}*��z�s��j��{CR�{�4k3�m�[�	Z�"�n-�t��U�C��i�mlF�s.��=-3��ā<[���,+�u�Y�@+�=�'S�lg.t٫��U�,X�wǸ:��Mr��e�Ko�����|j]%�С�n��z!�Bn*��+������G��0��E�O������a�s��U���-�J���tLW��� {�ك�L��v��ћ�1�lpV������JU!w��V�v�|��-%�w�[)��Ӿ���f�,�9;b|RhZ�����fe��Oih<����zu 'Y<qR}�Rp��m_��a��d�;�-�]�;��B���dvr^�W<4=��-�3q�T��$�	@0��ޚ9��K5ռ��go(��j�z$r���V�ӷ��{�D���#X5y֫>�C�<˶��2�E�A��r���(���q�q뾣|#ǎ���!ιu=�[SL�Trge�{��#^2���qm�3�*aֺζ/���S%�� M�˯~�oi�Y������
��$�Y��{ӧJ탹B�Rb��-Z�)������[f���K���
������LW�J�liq���#7n�/r�'Z&5���^n7iu�t���� ���9N$ZȐ��ݝ�-��,�pZ��Tr��36Tս��<�=�J�H6b�
5<Zn7�k&\��tR����@����91W5����⬌8��$�͢M�
㘞I�� t�K��Խ��`[�w�M��֫cB:�s|���Ǖ<���,�
���F�7�>x��'7~䳐v�Ջ�]������Y�d:(�/#AU��&S�����
�����K�َ���������Aا��B�6�nK��Lyx�n*xbZ	+�����q3ݙ�Fjh�G�!LW!���{Qkz��ُZ�ޚ:��D�:a�s1E�����/m<-���aw9�4�U�.pHs���9̌5y�����6t]��xh���!�j��K�֢�IvG��!�lP����x{��Ei�1�dL�i����՜V�˥Y ��{�F� s+J��2�eD�U�\��\���W�OAC_K���N�2�rrt�5�����ݜ�f�6�t�0���]�!u��i6�f�)���o9�&^Y����j^%��+�z����v�HN3`뜨�ɂpit��Z9G���Y�����KQ�������YW�s���4�N������3��\�c$H�ᄒz��jL��(L��9C���l��Q��X��7�f���	�~ۏz3En�S����<<.Ƃ0�#��o����{%-7����wjȳ,X΢�N���o�i38���;ѷ}8b~g�G��:[�p�������h�<�V=��N��_u�L�V���b���Ϸ%.�ڝ���4��}*����\���7NRfp�T��k�V�f�`����&CF>p�Gq���|�ӏ����y�-D�Z�]���:֍�(<I&+����Yۓ;lJ�]�٘�Yv�U��yt�UfM�ow8�؁6�9cf'�����w�JH;�l����vC�V���G�+B��f��A�!�9K�I���ZoA9#l&�4x�5���oD#�7mE�W�]���U�-�e��l#��e屝Q�ȶ�������k
egC�V�_M���>#���� X��Lxqr]h��X�H�=��cKŖ^��&�݌$��V�+g(�@�]���l�AY��Wt�[+(]��hg3� K+:��M�ɩ�&v��)w=E�R��i�jlˮ꽺TQ��T��n��vf�j!�u�8N|�=Z�̎%.�N(��"�N�,p���� ]����^tlή��f��I�u�Wr�}�XI�է��"$2���.m#�kL�P�z���'��N,Y]���y�BA�i���"i�=�8�Z����or�����[�c��1�;�r�dA@�K���#pk�x��p�t����4kz��]Z묂v�tf�+�;<
��|����5��Z�5N�`�
] o6��J��t��H����+���+f'��>Ga��a&f���@w�����s7�c�˫�y\��6�@2�'�o+s�t�5��>��aΜlNA��R���IQ%�{S��s:�����T���UnL�&��=��.X�պ	H-����cn��.E��U��7��|�v 63]cy��J_X�'d�K�3��є�uj)[�����Ǣ���6y��އg'��U׉Ic0�[y���F��uB�	��*�ZcCt#ݘ�Ŝ�|�e)�)g�T�֭�b��L�ڞ�:QO���K�S/k�	�d��!�Ψ�<e<��[9X��4n�Y*��ejO�¢�C��m.�t���˂�U3�7_!�m�D���%:����j���#��p�Y�x	���Y��Z��v)e�ʝe�n�L�����9QtbZo�T�=d n�(Cs8+7�Ȩ��YR��ۨ�I�_s��c����d��
���a����z�q�{E�V���9��"���\aoI�-� �7G�[�! >�hf4OY��p�/�p5�����oӧ�Rr���yKw/Vlp��c���j���jc׮����۹Ś��4M-)Q��z�#�4���3]=	g#�-����}V�����rBIy!e|y�ۧ�+��4&�Qk��Ր8�7;n�p�?\I ۾=�L&����u�kkӲ��Mp�,�	Yu��ɪ�Ύ��r�dJ�!������5�)T�4	����ɕnen�ne;�������ݠ��S�b�]8G��ꓛz�D��*�U���������E�Tx��'�eS�X��z��|6��Ϲ&���ZN��)������=��U�19Q*p!��FZ���}X:�q�w���)͚�[5��u.e��&0����Q�^��4��*7��M�\������\�z�g4Qn���C��x���3Ih�e8�yj��ٝ�L��L��p5�]�r�`7W���]�v9��F�-����%+e��FA���U�x�\g]��:�B��8�W3��&�E\���IX4i���`TNq?::���ɽ��'��3�tQ�y�{Ì�"o���m��=ځ�^c�����Ed��N�����R�E�j�`ҙu�|�X:�۷z�	తjh�Y��:M%O��V]�V�{����ѫWwE���v�1U�j�R�)�t��D��2*]��a�V9��{��}֣��/n�J�bv;�ܹ"�-R
��7�[�j��AX�.ƻE��ݪ���6L�%�k��]X襬eY�i�wz�|���c�fzp�����Gt�ܴ�M�br����<	o9)ҤN�w��w�ͽ�o��/hA�:N�a���Np@V����M�.,X5TC,��p�t��O����M�47�O3�nZ��N���Sx.dg�����K����u�]M#C�3Ћe��Nj��4������kO:�ـmo ��d�2�Ŷq�KmV�Җ��Eވ�R��5Fڀ(&���FJ�j����$���uŷ���Kd��+�AU�/!�W��۬�x$W��)���YE�h�7mVV����8��4+��V#�4Fq㪢x�;櫸�!�e+5�f��ٴ���J�-�uY�9 �է	�����B�X�U� ���V��U�X�f��:�Ec(İ4��onX[��+�#��P�I�b�Z�\+^
ȷ#c���E�B����^�R=�Z�COJ)im.���e�Du�"�a8&Ó��I!<���Ių�n'����I#�+^�Tjj7��d�NTЖ�yȫbϊ�����N�iާbݤx��&�
��i�ǏUh�l�1�\�N���٭1wy�j�����!)ܩ[in��V��c��#�].�t	89禸��vh���z�S�qU���t�4j�]��3��Z�Vm�]��H��cn��ѳ�P\{o:
;���{��ڂ��+� ��}�W#5��7w�uN\4�*�k�|�iF;���i����^�欩�'}ɼC��u��噫
m�]Y9�+����x��բ�zR���20`�����g]�rynne�3R�{9�T쀓]�L��)��;^�IF�}=O���m�96����4j�Z�k����& ����h�x+�!���fV�\�)��#�H!�1ͼ��m��ڐ�n����1Q��4�^�:[ko.y��/��P����3�Jt��g��E��M�+��Q�{�]�3O@���J���}��RZ����:��n��[�ѫu��6D�o��B�k�t)��n���L��xw�����L=�_u�K�U��2ȃZ�s�W7LU{H[���$R�{a=�-ͼ�x��˜vtż�DL��
��+_+��|��ح����u�/z�{��͜�b��{�!Օ�IVl\�K��k��`�,�0`kǶ�rg+�[�ml4����hgU[�S��>#o����lXJ����񁩮P�� ��:=�ؠ�t-M\���Ҽ3�� ���ͦ\'7M?-�qm6'm�Z3v��'� :x���4U;���L�p�2q�M�]�X�i� }����ܺۻ���f�e���	��Fe3��˺�,L�j�]N9��z�h��6�1њJ)%onRК�g�q�57��(�������:*�K|�==s$w�
W/�r,��g쎳�<�|�,qq9�۔�����q�����L������������뜨��Rass~�7&>��%_,�T��Z��'�^�,2/!�r]�nc筪8oJ q_U��'nǬ��FGp�a�8���F���%��j5���U�����fҍ�M�v�������oF�'��>�Ό����][s4Ztk�WSz�_.��jr��[W�^+:+$����;`���ҹp��ͬ耐�f����;�ۣL��X]Kd�=/H�n>(�U!}��;oH��0]�;��\U�H�6CyeX{��b����Mq���u4�%f������n�̍���n^���\NK,���H�/���Ģ,q�3(k䖸�"��#Rt�u��Q�^�������r�}�t���3ղ���s1e�ì�x.펈P)E��nW}d��Ps6sY�1|��le�;Ӫ$$yb4�UΨ#8u��QW\nk�W���>���N.Q��S'y����8���Z���+|���6�����<��w��P��̝[ EN�++E�=�������s,u7�;��e�4pQ����L��]H�\��S{h_.+GSj�������rյ�b����tTv���w);[���O��`8QYY�]_G�n���?MP�%�5բC͵%���YՒ�7{v�P��n��ځt�GX
]`�����s�9�(��se�r��}��Llh�F0]�g���u����ia9z7��S��o���n��m����-ܸ`N�p��ϭܰ)J�9�i�@�{07�:��	��hgvS�����x �ү��WmL�6���b�K*ͤ蜣ء���PF�8�i4��L'��릓���e��X婋�j��(�����&�U[�;�4�kU�y�uP�h'S��|
�H�bջ}����dk�w	�u��|U�)*A��Xr����ǳ$�Ȯ��]����_q΋�t;���{b�5�{v��6#0骽�V
��T��*�w��P;��v:��31�����_tV����F��;�X�[얖ӇN��YZ8U��:����vf��R�OV'�{ ]�U �N�4:�a\�ѡwO�f����V�;BH[�u�e����Y���V���^Ψ3q�K�j����s^q���S�ڇӝ��{�ʲ�nv�R\ڕ�98�稿;���.�:V6Ḫ��6��W:���p,�Ԭw.Ѵ�Ed������\7�s�\ԍ�9��R�x��[�+�-�k�W:�|�N��֎��B����s�Ϸ��5�}��		�	!I�~�<���۠5�>eM�̰�aPyj������6mcX`t���m�w��m"����[�t-DR���l�k"���MeL��)Q��/:���ݙ�v��9}H0��gtmv��J$�ݾ�p/;��P=�w wP�I�&��w9�M�v4Ȏ��X��8rW-�Y��{pTo�f�[��64�R���a!�h���gd=+/)'n��sEڡf�T��wO"��7�D��%��c[}U�աV��ǄN�>�ҫ�9�����% ʮ�棳�擳GLW@���f��0R\I��$�!aθ��݆���Gf��f�7	ibO����"s�,=�,�ۂ�ΐLVY�bi� ۑ�p���>�vwl�KH�,�ޣp��R6$�}+hk1�)i��Ŷ^7u��E�r����9a/IOU����H	qɳ�9G�f{���b7��ط6#���+�.v.�(D��3���;Ʒ���WZ
��.���h����6���r(AY�l։(�f���a�;�.�
*�
�')���n�5�'���6= ��u�
;vm��k&�96)2�Sy{�Dሉ6wG;�+��s���iC�r�Ԥ/+��9�PU��Y��W���:"r�j�y����o)�캺�^`q;���e-��Z�����K��B�-G���f y��h�:�8���֣]f����n-̲�Tc���=��5��]�@��Vt⭷-'�i���n�n���
Y`j�]�.��b�Z{&�s����h�gi��l��;vv���|)hC��Ks��\��H�'�;�
�ϐ����x���DB���F3z���[:����Skx_���b����s���f�1��m�A�ټ���C�����|���z6��Ǌs!����b�)]u��+:V�b������n)C_�=+�_Q1LO4�ZyM�3���\�i��b�c�]A�x��y�&����z�z��]JE��	>�d�j˔���AQ�&P�o�e�	���ƮgrL�^2�K|��&��GS��xu�M-���8G� �Q�Xg�(X�]�9��f��
j^RH�}�-�4��.��ʖׯ�ӯ����G
WB���BU��t*�ϕa��SݟMݛή�^LU���g`ajGS7��8%f��e��OZ��w�,�:�ʈ6DY�0�9��Gv�7�@��L���:F����V�K.�Y[:���twb�4s�	�2��:6Qxh�z��dԎ�]ht�)�[�M�zQ�Y+��0�(G7\�� Ď�2	3��Z�N1��^P!h���cO�;�����á8��GX�#��d�S.��.D�N��Zu#ZFb��^���Tocq`�n,�.�b�۸�q�7ư6۝-V��|>iS�JV�ʌU�ʱ��C�mB@g�8-	�F-GI<����)>u��*]�6-�;�C��Z
�`�\��f`�<����%����Z��f�)��1���[�\��dܱն�oJ�vm��#b�y���ƅl
��
���o�\�tN�x����Au�g��e��I5�&����w�uvm�NN�V-"�ǳs`��OK���|�ZY��N���b��2s�*�5�wT3��ȳ{d�:'�f��&�+�����w�s����NsUнY�N��#������4�"��%�r���2���T�2u����(�N���	�r�ثʗ¶��l
fV�'*�<��穧�y���`�e.À���j�05e� ��K��լKOr�ؿ��9g-�����jr�����T��u���{�jx'!�H�a])T�`�W��b�����G�Τ��Ѥ��t
y��P�ΐ<�cgZ��a7����� �`x�M���h��lv���Κ6�*ʆ$�7�/��A�2�M+�u��
��ٖ�t�N�E��r4ƀ�Lͥj�����7:�5�rڳ���y
u1�;	�5���\�W݃��Kn1��3�}�L�TK���_v��ݹ//V8٠�l��ۆ�����[��}�/��|&�x���M;�X��ؖ���}gR�ʲN;+�mA����Myo�A���L�D�^���_Pt�O�HS��9��i��Y�kt��X4�ncN�;n!܏��E;��{v7��,�b�\���gN�.�Ћɼ:u�$*��Y�bl5[,uef<�q6����b�Lɛ��*�!k��ck�{�+cr�(+2�Y5x�cB��)���yy����iDnI�*a�#
7��I�%d���7��YI9�/L}���ڵxCJ�N��efFƞ]�Z��[�h^�U&����sr���]{5��/���>j��������p���F)���e�^�v�����W9�|�ҫ���a]�>����_bm�Ǽ:əy���b�s������4�oTξn�K��sET�n>�O�a)��^�nY׀uZ�޻�w�~c�j6���M�5>�v6")5Y9h�ރT�w'X�Y��>�3�y6���ғ\C�j��&�Z������H*U��G5A��Y���d��фS�c�unJ�)�YWՂN
�k�\R���o�OV�ʂ���y'r��a���Y��=*�Z�ޣK�w`���\�(Hl��Y���7w}2�U�%fū���A!|�A�[�%�,
%�2U����7M�E�;�ӻ�f�nvw��
���J�q����Ҹ���Yw����\�z��+�jq��T@�`��Y���,y	�������$�]�r��54���L���7S�|�j;0HIUlݻ�y����n�������џ�6"�%iy��Xe+PL�4�`�-��	=��Z��;^�b*�J�6����uʒ�U���u��)�LE��(7T�,�����dy�����h`� @I�i�����i���Zv��a`�E�������T��i���qd���o�HiǛ,�[�GK���+����j%�����{�boQ۵Y�����:��y�3��3���2#�"�kH��s��<�o_ev�ĩ9���$��.&vJ1p�Ew��v<'�^��Ud�\�]R�6�6J�C^����=�v-�����.�����]i���Y��	�I�|��cj�׷�:ݺ7y\������n�b3*���d�{|F�Gk
XD�.gY�:��Z��o��Aκ*Q�C�ֺ�`�p��Nl�Q��Ie���+��x
�4vĸ�Z�EֵVu5���J��%�S��)��
���Y��cpLA�:Cy��t��՛lvm!�+��n��[D��%'WZ� 6s�&/��t�z#Ս-�z�z�<�=x�3�!��3]7�� �&RT�9��=��{�����:�5�����&��ǲS$guCs��V���2]�����yW��^�l�2���gL���l�8r��ڙ�{J�۠Mr�p���GH��s�<ܼZ�K\�s��w)��sڭ�6wa�]�(ÖgdnL4�sG�j3�����b��-U�M�O�9�|�b+��{��Kv���DHކ�����on���X~Me��*���ǚk�HXsLֵ����	�GN�i8@i��!������Pnd�3ӷo E�m�y�F�|*g\��J�V���f}����� �+��ǪfGJQ=B��緧66>��.�d�\"OT�!�3�H5�̚�_>��[Oe˥ʬ�M[u�^@����L��j���
WCk.P�֧�K�8{��[S�ҹ�KW֚.�R��<��,9��ͼ��*e���Z�A,�RN�Ѿ���d�A�r��B;Ib|�=3Y��U΃��#��J�dC�� !��uM�V�Ѵ��˨K����Ŋ7cw��Lh�q�����i3��ۉf����U�4�8�lT��ȋ����6�]Fn�Z��1�Xr�m ����:Pov���ք��Uz�w�;��PG����dؓ��I�9�[=�T��(�Е�Z���c���Z�x��lg_.T�U�����RB���Bn�(0��d4l�Ǚ]ʒ�0F �wҲ���u"��
��<��ݓtř����������(�fbm�a�`��%�)�u���e+ۜ�,���UɩUYN[�iǣ�u]7(${���1�z3�eن��������*�,E0nI��Iu��Z/F�b������d�(\뤭��:ق#��xs�n����9>#�Z���K�g3S0f�h��&r���_-"v�d�xY�m�Ъp�D��\�S�h^��V��d9����J�2�,�36I(�,�����Rp�༤/x��r|/6�r�t��Q�fWZ�dz�*0�v�9P��|�u���[üi�Nv��&�DV ���t�(��.
l����,v�75A��	'-y`��Ω���ΆKT�Y�q�8���!�ef�l��y���Wc��6)%�toNg��RΐEw�A��m}۱�g/<<�n�V�����+�G4�n�q^�Z�$��s^9Y���y�M-dG�FX����
���Js<�𭳷S��_r����r�fB�ༀJ�@�s�P�Wp�%��k���a9�l��X6�5��vb��� ��U�]q�v@�A���ɶ�b��e;w�]It*�}��[к����k8^��x�Z+
;ٮ&�_T�A+�s�=;6�u�u)�T!��ٻ����#0�giܼ��k�8�Z�*<��|��}'	h���ur<���sy)�Vع�Wؓ��a�Ǘ]�F&"Э7�˸�C��s���N��*o�A��Ua�[�*��q��Z�x��.�� ��9�0V��DbN�S�g����j���+w1�/E��T���J-����L�� ���t�w�btvMFw(�|�D��
�|s*�U������f� �"���d��À���F��H�U�0L��
뉻�0a�Þ��K��3����]����(^C��Pĺ�ή��t���;���Jhw�+�ڔIR`ev�ENF��H��\8�[��U.�{�[���V�;�u����:R��;8�[�>��G�o.�N���hn=����y��f�U���NX�[pr�_oك3���N5��OR7YJ��\V��*f�W�>[���Vl��v-�o����"��뢥�lu�8���Vba0�t��h��ת-[�u�t��7,}ػX��8M�^G��6��>�]]l��u�X�҃0��%�c{�,C��/;����w6�j��6��(ƮU�2�O:�(G.�&��n�X�*�"�L�Ц�i����Ҽ����{ʋwѕ�Ⱥ��dva��\-����,4��0p�"����l��צ�/w,:�U��hr��kԻ�-_s�u����3�\�\=xn��*Ċ�ujuq�f1�\5bs�y���������Z�Ǖ��m7ΝI�4���R�����Aة3�����:ۗ;�:�6�#T��:TV����g*�V=��y��qS� �X�8��
Z����r�-u�u�m�@�-J�oqϊ%!nwA��<S��ӆWu�9��v�)�F��w��}���,`�&[�ĸ�Y����ۣ/ŵ ��ىc9=�	7���T�-���Z5շku3vt+�x�f�GaWmk3)�}\N �jP�sO=���%�6f9Z�DѶ�͡�"M�cj�J�""�{4��7�ov줹�x� A�84wfu��yn���r�����Y��y��۸�7�9YN:��R����"�,�յ\,�T��,��P�z�VSYK��!4��I�\P�y��9���I��y�[*�}}P��ˡ�lݥ��b˫6���΃�����@����捦�K5 ���6b��GM��n�v�[��,�A�LX�y��їa �jv#0���\�p�f}yIf���I�����_T������7����]P��c�p9z��o�9	��%�K�M�F]ɵđܳ�9��Pq�,_!MP����#X��}��i��5J��z/�}B_-{2��YM��zjF��ysE���6G��Y�cm+�];�.}��Ff��c�5��]��O	Eba�����.:�?fą�7y�3"ǯ�m�4��`�6�]�Q�6��Y��H���X4^�
ŕ�܉	��H�S�{%<��9��^�S" �l�j�N�f��j2֪�|�"�������Ǻ�:ߡtr�|�j���6����ő�O�@��W���ݚ���L������N�&��Eջj41�_>����%��0�w&�y��U����C�}w��b����܃�M���s�%a��E,[��]�z6.�t'l(<B�ۓx�S���4��4/N�����N\�r�հ�b���VK�*+ͼ��5x�ۨ�iɵ3�X����e0P�����]���!)������h��u����]gN�-R��m���+P2.�c1��&%ۋ{^�Ut��
U�#�۬�cC�FZ�3�EX��,���3>!ܝŽ��mM�CD�CH��%��b�@�z���Д,7��r�Jw�B3H1����`�GZG�@kY�$��p�W��h'74V:G3��{۲�[Yx%6�R���x�Y�gg-P0���O��HrG_���5�WoD�=ڧ[02�����.�NX�V�۽�.�%]�$}D�]�[X�sj���'ذ}O�g,��B3j�^�V��S�����[��w��ѬQ��g�JN�ٴ�qm�A���*7b��Ӑ<�t�|`���Q�_=4�Y�Y�N�
�t�L��F�S�p[o�H�ї2���jb�;�����k�&���l��aT��/:�Hq�ڜ*�^M��n���}_}�}U��*�yK�/�F��L�������&����˸ħ�V�E��^a��;�\�[ߌ3����:��n����[KN�O L1/�O �Zvnq�V2ے�x0�Q���Q��������|XA��-U� �W%�.��w�*�- �	g%�h��o 裘�b�},2�h�l�W�J��&�ǜ).�v��k���Z)�ۤv���^�qc�ga�u�j,��{�Ͱp-�2���x������ w*�H�r���ά]xb�΢G������4N;��;�����r����8����Gυ�}�I���W�Z�E��7OW1-��^u_tM�Bcg��gE��\���{��9�����m�΢�k�c5ټ&8�ѩ-4Z �^Z�:�i����0�B�M���,��l|�6���V��G:���9,��T��2���]=��.t5c$�ZUd�+p^g'�Lac����Lً`�U��|GR����|�^v>μ3���M�j��8��g�a[ֹmg�{�q�Ո�9w���ovo��=�Jz�P���Ǘ6�m����ӡ�XIR�{(CĪ��
���z�o��K�c�x0�7�\���z����r�4�xCJ�XY���o�L����]2�㢬�6�3 z�5:�*T�����T�6+ǻ��m�Ԧ��JNY�pQ�2��O����կ˨�{݄z��}���ڊ1�#X�Jʣ%�EdTE��YJ�R�
*�H�ʬ��U"�
"T�"�(���(��(��R
T��"�EV�
�Zʪ1V#-����j0kb���U����(�Ŷ�QTQ"�AT�����Pm��Dckh�V��D(������eT�V�����*��+���-*�DE�j�Z����B��Ke�-Z���,[J�[[VR++caZE�U�´���[h���*V�(�"��*,UQJ�e�ږ�kX�(�QA���-[�UQEE5�ŭE�Qb�iQe�m�Z%QEm�T[j�YYmTb�*�iR"�Z�,X1V(�����AETTb*,V�+�0DEQ�lU[J�D�UE�J��R��*6�
�X�TDb��`��Z[(�U�U*Ueh�����l��䡢u�����/�� ������AV��a�jr�6���G��z�]�#3 �
{��n؀&�΂I��qܓ*��m�;�����q�kzn��g"+>}t>�ਯny/CY��+�a76o�opOz�R�>��S}���s���{)���v��}��Q���ciJٚeC�楾���?HV�I=J����s��)����7�O��F��u�����i����H���p=��-��v �ź��Nv��Rg[��T8=
?S�w��nԱ�Bk������W���-�{wޛ��]Ż�iי����kw�74+e��1N�b;��΄�%�V=�l&9W�t�x�SͿrJ*��|���<`��A͊�[.z��n�}M�ii��럺Ϗ�q<���5O�fh3������V�﯇k�Vy٣1�����d\�:�����Gꙻ���a.ݯ.���{�sI���,.�@[���n*x����o�����6��H��i�����{8V�/]I�|+Gm��@w�ǌ�<�k�1��Ҿ���8���)[JT[N��g���!��m�a���4d�͐�pf-+�V���z�G�e�e��E�Ge;{�]���LD�Y3�9:�ڻ��&/����:�lt5�����/�b�������J�t榏zb�Xj��yn_��Vs����H���j���Qw'ƾΏl�_��8��͸�.��>r��ߠ��ػ��,�{�o_�V��;�'�+1F_o@���T�o	�纬;���;�;\��_s<+���+~���!�EKZ�,��4R�*X]0syܞ�9�	q�����D��_e��}.������V1{z���t/۶���sR� ��[�L�^�D�젵��fk~���;ڍ�<k�=ԟ�!w�to����T��Yr�jYI�O�^-���:ww�X��:��{+ԻUG|�7/���u��g��̉�W�9��l�𿹇�r��˙�Z���b��d��Jrb��;�ݳ5�3�>d���ǜ����9�������@t*��9����R�Uf_M�o��Tz-�V>�����"�Qg|�d��_���O���Ѕr����!��9�N�J��oA1����:�'R}5u��5�[�ئ�do������-�1R/�kgA]8���y�vk��{8��y�����!d8�r�Ʀd��mM��{�41�6��F}Cf1�T�w_�G�&xz�97Y�}��Tw\�t/i��SW4>��ўɯ�ߤ�-ك����y�]��T�t|���^�ߺ��zv�{LX͌_�|�.���g�����Se�L����<}�ռ�=��2Ǵ�]�����F/5��pUm�[�y�暩��<�y� q��s���l6kl�ϴ'�igxh���W$�Kr��r��Ύ\��q����I=��;������P��S��5�}�,�OtG�ç����Xt�z9�6	����]�ۗ)1��v5ׁQg� ]�$�f\I��֟��u��=�a��H��ڭ�Q�|n���<���OZ���u�ί�ڝ�7۾~�&��\yrO3�y�W���T���z��c�YS�/>�����j{���Vy�y�P|��.�՚�<��y��Jj�J����k{����pԙ�e��m��x��yo�]�_	g�;}� R	m���m<N5S��|�����cQ��)�V'p��J��PƧP'�� ��D���V�]lwa�9 }���Ƴ�6f���{=�^�O��y:����/9��s>�U���V@�dT�Ώ�������}=�%�ʓ�N���U�0�#׵��+��^vA2�%ӡ�lO��NƩ���'��Ws�e���C��������[4fK͈�oH�Kb����6����E�g:�V�X[~���>��	
9㕻��,��~v�U�����v�X����������[��ǩ����u��Q��՞�u(|��>�L�F�A�xo�OO��e��7s�o��ry�(�{7��u{LX͌{��I�i�T��c��\��O�ͮ)�w�e����:�+}�i��Sq.y���l�Q?^�߄�'���^�s[�Fk9-�ƣ�Y���T:��E���{�r�GՉ��gFu��9�q�l��d��
x��)$��2��#�k�^}73�-v\���]��aR_���v=��DX|��e^L�(��j\�QQ�Յ1_(�$�vU6�n�!u��S+����sBS�!��Y�^��y��[���nЎ�M�,��62��T]������N�������V#��v���1�n�l�æ�L�x6	�}�WC˥$�[�W�m�O}�]f
/���J�	�=�a��S6Aޡ�o��W�:{�3���v}��k�<4���9о���e����X��MO�m(%�7Y������:�����OZ約���@�u�:P��̮�SҲ��-6o��>٩�'=��2_^L�s���_��'�J�M��GC�x��ۆ��0��(:B������fU�ѻ��o���GǻZ���x���2��ٟ-�WS՚e|.��j[읁�~�!�O?	�;�f5�!�;-�?MI�Z�s=��c�}Yz�L��ѯ��RS{�ɺ�˖�k)�:O/s��S�����Z�`��I�n
r����Svw�)�v':�-?#�tF����0=�����3��{.�����<^��e�X� B��Q����g
�4���+or5�v�Z/{�)3W�P�G�{K�ű\u�|F&�ff��=ѫ9��Gij�q]�i��Ǔ�m�wu�M�G@�����9�㜔ܓ7��Gntj�Z˕���3s�z��qf����\=-���ܝA�"��y�;Gmy�s�V���{^��f��~0 �VU���Է���a���_Z>�;�E}/�uny�o�<��||��sg�g��37NP䭜��]^��~��qM7��Ō���v:��|�~͒?h���8����O^zzy+����-���Mb����rӗ3�ӷ��gkOzͺnm����l�lƶ�S��,SW�7�ٿ������eo�,^{u�kOB��\�.�P׽!���m�)�^j.���M��ja�%��U4���=ٞa�&OTs�����u�-Kz�Ϸz�Ǻ7��~>�u�u����=�\��>=�a��nh;��b�օg�[Bc^��ꄍ��j��9�wr��_��/���h	�9Չq�����D��gyi��I�4AS$�$'��AOu�%����g�ohOz���[�z���o7���S�wk��X�m�^o��ۧw�R�����^�.���WՂ_:��j�F6�*�6�EG���!Ae昻���@Y�!<��Ƭ6_Qg�>��`[e��ڽ;#ad�9z��f��ObR	�#/��O8]�:�R�g�2f2�N�}�"��9����)Z�l��4�W��U<9=����~���v���b���ڦ?6+���X���>��?J�}Yz�d>��n����l'�ғ�5�=���S�~�k�2�8����A?fஇ���B���v���D�O�=w���5�� �b�p?��9��b��o;�	�q�]	|7����ܮU�o;joM;��;��_���x��u�z6߻�<=��Ŕ�&��S���n{��y��c����O�m��1�Y�߮���k{=U��6�)��:������v�^���ZS��7�=��^��M�f6���_&�y�e�iOtr��?V?ui]�N�X�B���u���T��&��-��?o�'{>w��XmO)��!��Ͱ�eb������w����Nt<�'���$��}O�Ƕ�S�%oAw�k�)B�Ǭ����}r��Q��i�9Rfr]�׳�Ή��
	>��y�Z�����(py���\3�"\���V�%�RmC���[��$���h����b�`11��ڵ�ӱ�,�	�ymg�)ǖ�W���}p��H��.��1F;y]R��/�Ώ=�������`�ӰI]�?@��?q3�O��|�N�g�=Q��+������pk��uXw=�$�2E�{������W����G�u�C��@���ί���vY��ty�X�ή�;V��0����w��Y�^�8S�zС���Ҹ������n�0�S�����=�/@�{�y/�.K�*ÿ��+ ����~���ދ�u��H�Ɖ�7��7��<�*{�K�'�U�a�F�ω~�IN5�w�9T��{�:�8��Z��'2�����ϢoӍ�����}���b��o��͔)@�%_�ݕ�~̗c5�CzEbKb�Ǡ�T��c�*&+�av�x���VzT�:k8��"<���Ϋ���Y���~9�s��\�ߟ{S�=Y��(X���u^��f�V����~Qy{efq��bGы+'--���#�����e.��v|���6�u��Z�����MH���<r�	�P7v��(a����mެ��[3:[�`���t���f�=y6t_X�!2��2vq�d��F���xvVtA�j&�;�D���}}R���u�G~�˝�������O3e���9^��x{�n����U���x��7>�6��{�x�_������t����nOk\������0���lf�z_˝�����?h�;�)���+�4�5���o�
�[r.ہHh[
��sf��i΁ǝ�����v�a�s�5V�����Y>0�mm;K�u[���|9�:g��}�[,_K��y�u��ߟ�t�>>�y��y��S�C{�X|�]�)���'�6η=ܽ�k�=�fX~��a�G�-u}]`)�gr2�I{�c�롨����ڗ%��#��7�\�{�6Gv'bw�+��_�RAGۦS�o6c�n}��9��=�'=��^�:�����+��.
��urZ�u���n\C҅�u~;C|�~Ozڗ�����V\إ����a'�4����ʝ�v�R�G���Z��n���ܢ�oA#>�z�%�ϝY����Œ�z�de�t�Ml������f��+o5��U�S�6T$�s3P���!Ңj��g%J�7l����n�:���ۺ��D�N4Z�Z�Q?cE�.�Q}��3'r`_���yC�ͪ~���.���K}��Od+A�0f_U��l������=���i�-�Ϳ/d���<������O��7�	��~�yO{y�g	�c�9���˘Փ8q�У��ż��dB��Tg7"������{����r3�˫5oR�^���]F��>
�17f=���!{'mA{��� �q�&�=���W�ͧ�.[
e��E�x�)�Nk�o��i<�j��]=���^�/6��ߧ�z���Ѽ�a&�v�*�z�T�w����u}Lf�;o��;�n?l���A��|T�	�e����_����Z�j�U���8lnXN\�F|-u��G�/���{�sם2���H����c���񭵔�%�t����˝~��u
�^c��I\2ܘ����`rK�LR�>>�Qs'9������<ٮ\������H�Ҿ��}n�pW������X7 A3��ū=�ye[���7�d�{BEJ&��n�q]aJG��m��f9��j;Y��Jͺ%B�鼹t�@��;�lo,��.9eSLmkWX���V�wd��ܣ�b�X��boe��j�
�zT��v;�|��nV�1Ri
��n�;f���G�Ë�6�������b�D��p�礼xc�w˄Ź���K��]���-�,��x�u.�H卍u���;��"�AQ�n>zӾ�ة�t3[�r�y��G�v��e�1�H�9��x�d�u3�l�c33�B��7D�쾊ԏ5s[�S��;"�\����m�>~ᙨmb���i䡛hsFR6w�G��4EÔ��/��gPk��|��s2��0�ߐ�Rc\�AKQ���m��8;(pi�_ǫz�E��dl�2�h�]�f2���Q�;.ֵ.>F'֬��Z�ʸ̺U���b�xR�{�eS��YA�&��ec�ġuǸ*�nuH8�V1j�9���9Yce�Y�(Տ�E�k�`s.�;:�uy[�[Z�X\k�w=q�ht�y�v��8�S�����|#��NOoN��R�z,ev<k���VtO9�v�=�ķ���kk�`hZ3c6�u�JTE�����|ޥ��r�P[1�!,���%sf�  "�S��@��5�R�7�ڧss�_k<y�$F�g6X����0��w-���:S�]���e�74�n���U&�]�������G]W�����ۉ�|���Zo9��S��P��;���9o!U���/���ܾ���s�sj��*�p;_�2��Z����޵�y�K�Ĵ�(� �Y��K),��J�7��0kýri+�Q�֪������h�e.���s���k:vBZ/b̔nlS/M�ybsaz����k�Y��)JWu��3o��rE@��fCj�`hKn���Z&sb4�ܴ1������|l��%�"t�&å����2�����܌�֋���W9�ݸ6�e	��!3�)�$i��M(�y@u�8>|�.b�"��`��A:�GH�kѹ/���b-���=����{�p���__<�\36pMi�k�'Z�E�;���q�r�6x]ϙ�k�F�8h�ԭlW��j{ 5��|�:T�x��ǎ�8"��s��<k{4`�� �1��)ˬ��;*�/�}�H#��;.N��c]�.�ql.�9����9�Kựq�Jb����u�݅l�%�+���k��֦.��JG��:l�5�%E����CRCJ�du<��R�Ȭ����c$\�Q�o}��R�m��[�/6<��
�]c��e=���G��m$��^ly��ބ��j�v:�@M�{��4��#����껰U���{ͽꜧN*����yx{H��Q���v�Z�v^�o�i��|�	4�+UUPUm,T�PUKe������H��(�b��VR�ATUkQED�#%*�-��Ԫ���F�b���QUDc�kk[E��E��+DEF��V�m���P�"�[T[J#m+iQQ�TKZ	F�e-b,�KlcU+�R�m�VҪ �TTYm�����QU���T�TAcTX�X#TQDJ�QQ��QFDD��J�m���T��m�U���K�TE����EF(#TD�,-*��ZQUU�*,QUV�EUQ�**�����,Q[EFUej�Z�Q�"��*�hVU�5
�����-�Z�DA`�������P"(��U���Tm��-*+RԥV��eJ����H��""0m��E���T���H�(��FQ�P��b+UEVڃmE�X�T�[-F��ek
*-j�QVEPRҊ[UAe��V
�""��b[X�Q~��Vf>l��9;{QY7�80�ݙ�<V7�<��w݋H�G���4��'R��/�M�6��/7bF��8뫒y�K4F����~m�)]��9����v��-K0�{�՚:w���;�1+��R�ʺ��;\��/�`�y��v��U{ݻ^�M��Eg�{�	�M��g��W�γҰ���� ��g�ǟg�Oe�':��Ǘ�=tF�u��L�~��+������n!<�Ou�����t/ۣ�(r���X��C1�C��K�J����.��뾬��ht<i?u'��;��ߔ'����^b��+��.���ju-M�V	`5�י�Z~�b�W�z�]�Ė�o9�10�ٙ�09��H��v��$/��;_9�1�Fp�П�A�s��]�ͩ�?R�s�1���k��7��;Ne�5l�,F�������̊�wn}^���R�������8ۘ�c:oԖ�;��TJۅl���r�?jڰ͢�����1�sC�=oџ�˯Ɍ���Kl�:Zx�I���nr.�Q��Ytf�b�]
XF��Y�ޖE��b�I)�I;P��w�d���ng:��)��C���fM��Rr��w|�ѝ����{:5:uA2q�2%�F��L�y�㵎v ��N;�l��]J���Ғ��$��ו8]�Ӹ�:f��T�7����%i[��	�����_��[޺�[�A���W� =����VoNo!K�&��J��v��W�\�:_S�z um���� ��as�:vpq��'{��l��9��+ۉ-��:<A7}�'���`���0�� �/{$��
x��x���]��c{:�+u��Yd����-���5�A��s�o`�w��zw��%��	��~��%��WZ|kM��7��u7�!w���f���߶�<���u���B�C�Ks��v�{�'��]Y�ۆ��G
�G�����^G+f7����f�o�f�[�OG'�S$W�r��y͋m_eou���\�8ݿ���2_^}r]ʰ�9�t<w���`S�8{�&M�)��w�W���%pl>��Oqw����`'��7�^>�w��W1�__³\��Y慙�!\�B��AK,8�����̭:�׽~\���`�|%��"�r��^Պ��5
.*��n�7B�h�p�i�X�:9Kk2E���yT�t�䔏 ������o}��R\&q��J:S��v�N��7����f�=Fs���?ٿd>�jy�NϚ�/��'�U��eS��~�l:�鎷�O��8;�V*:z��^4}�"�%�a��a(��s0�mzǥ�(�ӡ��l�, }+X�sWEM�t�����B$~�VCǝ�zK'�n��qn�T�yT�XڞALg��ݫu��G����Z<���F�$'w������[�f�M~9&�Ǧr��}U��~/e�؃�l-�	����U���|uGv�75�����~����s��S��ߔ���Z'��{��:�/՚��4g�=B�\,f�V��\�0�� ��k���?g$���ݰ��k뱦=�gx&��R����b� ߳�65�iΘ�sg?>(q� �8�u�F��|ݷnoWyz��K��u���hy>͇PXN:aԞe`i�u��S���Ad���x�<��<����w9=L_o{ן����������O�ONw
|��o���'Y}�I�H|[�d����I�jb�m�y0�8����+'�d�'_��������������x3�d�~���9j݂��l���P��wd�o�mG�u�~�fxse羉l.�C�5���yB�<5f �B�#fc�:�%)���R�=+nI&�LW�V�4t�W��n|�u��e�D譋�"���e�������{���� �|���|�e�^�$���߰��N2j}��%I6�N�Y�8�j��VN �ͤ8��<�0Y'u�C��I���8����9��w��ӌ���+'5d�q�l�!�,�C����d�i��x������',��?d�a:��oY�(L��P��Aa�@�M�q5}���s��۞����w��e������<�a�O~�^`:�ԟ<a��q��׽��R|�h{�$�i��4�Մ�2�g}�Ad�C^�ٓ(M�}˽������3��o^���9�e%I�T��i>d�Q��&��k$�i��W�C����|�����N�O2i��v���&�Yú�O!���{�iϻ���o�n���������L���bL%I=�ĕ'Y2LRu�l�r�6�O�|��2��W�!����	��4��}�.U?}È���+��/%���DZ{�������s�T:ɔx�0hm����O0���2a*I�ޤ���`k�d�'���	�?�i���~��J��Hj~�d�JÙ��;�~�~9��}�c7G߾�?sw��m��s�e���wP�&�Y���
��L���M2O0���0�{a�H�s��Ru��4���:��gT4���N����}�{�ke����^�����q�g�0�d��1�IYP����IS���:���i'|ʇg��&�3��ɦ,��̘~d��I�l��q'��{bk������]��e,���d�~��c��������C�?n��2��S�`��<����Y%L��d�T&�{�I�T?� m�l���q$�ϻ�I��(�Oq]_k[����g���{͞�I��a����g�CI:��|�2u��~d�2u���'�:���ɦI�wt�'R�;�؟$�&�I��b�8ɽ���m0���N��{��6��Y�AYRO�۸�:CNr��Y-V�`�o�u�1��M��S��-�h�$��R�{��>���&���9hu�WP���>����[o��8���$���Ҷ�����F�D�ɐesV.Z��� O=��ػ��׼����dw����保a?07��N�a2���"���M&�u�|��C�:��j��u�G�'�y��.��q'P�,�e�~g{O?|Ϗ���د���g;w=y���������5�O��2m&����I���`�p�I>eB|�d�Vu�~eNj�PY&3��:�ɯԜIԞeO�Bu'���x��[~g�������~����8��~�Y<�oY>5�I�$����'�C�8�ɖ!��!�2���)�I�<�C�,��3�Y<����ϧ3�����F���?�GЏ�����bAd���<I<���'�u�����@�O�2~�'�O&��ٓ	<��hm��l>CF,!�N��)�I�!f�����÷�z�g�c��Dx���Q�|����$�'P��q �u�S��L����y'����8�猟���a�I���k2a'�<�d���jΩ��{�ݫ����?}�~�0�u'�8�d�jd�AC��d��~�Y8�ӿ���&Y4wX<�o|�����N��5=�ن'�?��������7���������0���:�d���ց�I�h�I8���VL��f�6���!�y��'R|�����4{��ԓ,���O3���i������e�k����|I��'����8��7�I�&yg���Jə�Rm'���L�VjI�i��|�d>����|��w>a8{��\z�Na��g��M����qa ~P�����0��P�C,��dI�4w�fL%a2r�aY8��&(I�Nf�3a:ɴ���a:���$�̇���8s���0~מo�g��<m�Ԝv����:�;����N������m��!�6��k ��I�q�2a*I�ް�� kN�m�٦�l'Y8�����u��Wߝ�S���Mb��A��v��s����ڵ�}�p���2d�'��j�k����L��Ǿ����K��H���\p�d���M��)��s�ս��7�����G�u��{���E�/�5ق5����ob1�֋��p���UQ�Z���k�y߿�N!�I_�e��]�L%a�Ӭ:�9����N��=�
�Y>Af�{*O�w���I䝿�&��v�dۤ߹��gv�߳�c��cG�;ޟ��}�?2i&]'�Л@�4̿$�C���y�Hk��IR���0u�W=�'�u!��P�&Ұ׻�'�3�~��	�M|����<��9���~�5��\�>Ǥô���E&��ŇI��?f��!����&�u����'����'�Vr�Ad�:w�d�VC]��d�Vw_������s��O����;�
���߻�&5�}�0��e8Ȥ��C�$���l4ì&MS��'�u'﬛C,�A���'�<�]� ��C���x�]N���/�ۏ�λ�~�N�d=��>a�M�I�9�@�'59��ԓ�>��&ܤ�MrȤ���L�,�$�*i��u���>fRuA���d�1��߳q�7����ƌ����}���4��8̤������'R��N�y�o�9��̛I���o$�@ީ6�$�o����d�hŝd�%L�è)&)�Oc�}�|}u}���a'P=�'�m��Y����I�4c�:�0�`�d����:���<{�$��6��d��P�VL$��
_|4�g�P�����:;/}�r~�Ұ�B���AI1��d�V�Rq�Y:�����O!�wܲO0�{�̝~a=���O��{�N�>I����~����^#$�4��v<�����u�����~I�{���'SS�I�8����ua�N%`~I�d��ϻ���fw�'�d�a����z�o��+�?��#��������.˕�y�x�d�O�&q�ա�T�Aa��Cl�M�N$�h�3)'��'�2~��N2y���Ă~����ő��G�!�/��f;��EU��� ��+��Y��k7����gzX[M�Omf[�f�n>WՖ�2�=j��[�I� ����9n ��O�h �I��	%�����z����� ��a��/���6v+�euf��٦�񝲚��p�����1�\�������?$��$�Nt�'��O��B�M�~�$�
���T�AI�`q�y(�8����q�a:�����>�t G���Ǳ��b��g��>?i��u�`a����8�$�MwX���O�4�Vl�&�;�a��k��d�
����Y>��6���$�O&CV�I�~����&�oھ�g�������VN?$=/18��O�!��q��4�8���@�{�$�i��4��'��&��d��k��2a	�_$��Jə�Xm��[��9˿is�k����}����;�>�&�0�a�d�g�P�J��d>�'�I��}1��y�w��,�a����y�I�~3��d��� ��I۬�&.�o����Z1�`�����}�cߒVM%d�?2~d��3a<ɴ��_�O!��I]�3?}��&�;�4�̓���2����{�u&�Y���O!�Lc7�����g��/����g��~��|u�~I�x�$�+	�s,� T�@�O��ٲ`y2~��䓨h�`~O2i���c�&P��y��L&��d�
A�f���;�u�߷�g_~�~�`��L�C��$2d�?d�$�O�q�d��$�,�' lŇXI��?�`~M!�̚aԟ}`|�d��<�m
�����w8˟;?w���n�m$����l�AHw�i'Y>J�~�Vd���gl����ٓY'��i���3l<��O���f��u�Ω�e��:��5�����x]{��{;�}�M ���!��0u��4wx�I�VC_���N�m+z����M���x�0ɯ��I�)&S\�R~~`f[��3��8�����֟~�0���+���?&Y>Ad���y'�_�I4��w��e�|·w��ed?z�d�'��8w� �i4w߳�l���N9I2���;�ݘ=�~���L2-�v����rN���[p�-l�vu���5(�M��2�X{�Ŵ�.[ ׋	BȺ[3�?��V�NX/&���Vw}3�����CX��ڑ瑫(|�-Y"r��4����>+����� ���Ә)��]B���w��$'�|5���]w��!���I��$�2�ua�a2k��u�S��:�䩬��N0�c�:�d���w��d��'ｃ��d봙������>��5b�=z�pw~�Z�}�ڗ��~��>�M0�ز&Y8���'��AI1�d�
�I�N�M}�Bu��h�py�$�׸<�߬&2f�Uw���E���۷_�:�Ï�B>����$�i6��_d�IԂÉY8��b�|̤�5��I�?�����~ՇRy�����u��S_������X���n����mi��T�}�����������P<�猟���:�u�1�fL0�Aa���Aa�i!��f�\2M���&'�Xu'X�`Lj���ѻ���� ��?}�߻��P:�N���l&Y5���N=a?o�XN�4{�IRM�]޳&q��Zy
�����'�F$���C�o],�V-��K�#O�}��R�~2o��ա�O2y��ݰ<����8���'�M���O�?''��N��=�`�a:�緬Ʉ&yN�Y8�Ð���q���x�N��o��5�6�L�O`�N��3�k$�i��=��}/0d�O�0�c����h��q�O�m�߱'�L�a����N3I5�}�Y'���e4�����7��)��@$�r�>�>eIP<�l�O���&ٙ�k$�gVI_�Ϸ��$��Lw>a9��̚a����N��8��/{���ߎ�Ѫ�ou�����d}�;��8���a*I���J����'�6��/ٰ�@�d�C氜a�<��2�gXL'�st�O$�q����{��~�yǯ��׷O\��4�����|,�Af�;��Cl�=�d�$��q�d�T�3w�+'?X'Y6��.�Bu����_�N����W̚Cx���� ����Л�[B��y&nȫo[Sz�󻄽��1��w�{�5W�G��W.���]َ�[�w�|�-كKz�[���k��-��q;��3��J����k�loKtJ��C7rK,��Vs�u>�x�\z�XK����W���v�p���� �|8nß�Jc��Zd�J���`�N0�N��d�}� ��M��^�T�2w���I�wfL?�'�s,��`T�d�M?'�hN�<�5�쟝�����_�i�w��Ä�I�&���C���2Jʆg���IS���:���i'|ʇ}��6ɟo�M0�d��}�0��=���G�x�o�?=f�Z�=����7��4�N���2����&�u'����'�_�I?!�7��Y%L�~��N%Bj{؟$�M����l�~�Z�_|�Un�ҕg�حpۛ<�X��L���E'��Ka�i�jn��u	�T��d�$�}d�d����I����ɦI�~;�d�T&����'�7�LyG���뻼���~�[�3�`i�,��X�	���o$�)��I���O�y�|���$�0��d�&�Y>C̞Au���:���g����{��~/��5ñ�-����׍2u�	����N�wt�� |ɴ�I��$�`h��ni'��1B|�d�hŝd�2�uC�,��̝Ad��N$�O2��������m=M���x����w��I��pu4�u���d��	�w�:��z��bO q&�Ӻ�$�05�ed������'S�S����h@'��Ʊ���(8�����3����'�6�i>I�T���Ad�v�x�y��<����K�?;d�}�<�y4c߳&y!���+&�|��XC,�N\9�y���̘�u�<��?x�$�OL�y2�<��2y+?�8�̝��ﻉ��;��v�e'�g�m�	���$��'��>�0�8����Q~#��W���h�s����m�ν?!Y? ���<�̝Mb�a<����q2�8�1C̜2-�q�ߨ~���Y:ÿ��$�d��y&�$�i���>������>b�F���Uz�e��1��_Vh��Xn�hI�\1G)�Tb���(�7ecgt#���L
-bz�A޽<�UxR���J7�ս\��ھ���36��Z(.�c�9G~J�5�卲;]vmk� b��[��i�V ��;I=�JsN��$5q���=����w��a�m��9��(N3�VN ��Z�m'����q'S&�8�a:ʆ�<����N������0���ǩ&Y3�{_o��1�7�W����M�a�>��?}���{�O&�59߲$����0����:�d�VL��u&�q�0XN�y3Xq�'Y���������<��1����S?,�]��SI�=g�����ۃl�I���0O3L�a��`'��&����u�ٓ	XL�aY8��8�u&�9�k6��L��<���I1�|���Oa�O~J�_���fC���|���4ì�����N�����(e�h,�}�!�M{?�	��?fL%I37z²m���Y:ɶOf�����~��ݸ汬gzw�~�&�0�r�>I6��I]����d�J�'9��<�;��):��׽�T:ɴj�T�$�}�3I'�~�>̘J�x��#�5�����[~|=��>'�� &O̚I����fuf��N������2i��d�+��Ad����y'PR�� ��M�a�w*O��4gߞC�ͿÐ����o�>������9��&�M��Y� dŇXI��?f��!�4�<ɤ�a���2��4}�y�������,��N�������a�����ɿ�L���9o,OqJ;@�2�н��o����;����P3J����:�>�g�$���ߧ���:�e��.:�����ͽ<�
sF�G-���������m����z��x{k��P�~��W-�;�"�R��	N�� ]�UΣχr��:c�w'8-�D���Y���D&� ��Q����vwu�������)���Y`�+�@C��gZ�h3��7wHi��}V���r�e�Z�ivNɳt�цT���uf��B!8�{#�&��Jq�e�]f[QzC2���j�üT[���R�΄n�[{N��'M^��8j�CLʺ��'a�'�i,[�|�X뎈��7��o17��d��.�曙��Q��v���p�,����9ә���s��Ht#�@��L��_^���\����a[2ڴi0��A���:3�e�tͧK��fYt��tSwt�{��M�|��X��r�,ھ��A0 ����Xb�w%��'�me����[��J�Yh��G��R�k�s����jMC-���n�CRpe�ѩ�3��r��Ւ�^E<k�H���OW���^@����۹���u���^z�8���Lr�RA�=��� �-[.�nn]�ǭ
��b�L*
fj��AS�W��2��Өt�����e��sWH���V�6�C�v�����4X�1����\.���������7a.*�rl��P�=�`W@5���뮋QբK��=ɧy�Ԝg:��T��ޟ]ݑ�WZ
�|�"���rj��M����Fr�!�B��7�	�b9���5�����-g_t��|�!�y˧c]�9���63m8s��W#�v�>Lc��]�q�-�5��w�p�Tq,C}�Th_^e��1q)�+�� vm	|��WϹ+������3�niX�;Gus ��t걗˳�o�������a��:�D^��P���un�h8�=��3Yx���KND�ˎ����'S
߱d���/�Ç��[�/�6�&kR�y�Y�r��72n��"մ]���W7,��m_w-�np���CO��u��<!��
�sưX}V��T�6��1��Ҭ�S�{�#���kpG����ŷH:[�7�h�W8�&����+��<��]-����&�����B�+.V�=I�n�t�\�&���E|�i�FRz�U�ru�so�n���Y�z��)�}�2��JL��R��{�1b�k�X.u�n����tc't32X´Wh�`@Q��1�pk-�U�,Ի���ghZ�'*�$ӭ�;o�V�,9�emM�z�u�\)�b�ip� z�X��P��{���m`�XH��n�2:{B������Ra��oq�\�>�?
�1�o���:��uU��F��z��.�!��yܚ�)ȼ���]�"�����p�9hw<@��e,��gX"oV�N��7xPƀ�72���k�oV�N�;"�,ݡ�]�Y�`����I�vS��������[Kp#�:�,��BmKRE��NX��zm���Y�P����ۺ+O*S�����Rg�ٛK8�+ʄs�nsV<��ͬ��+q5�i�6��m��6�kH�"�Ŭ�*)R��b��`�b�UP�TEPU��-EY+TU��D����m�,R�Z��"�U���j4���EjҩPYDDU	RT�,�*UdX�����F��b�ZPX1"ŊT��EX��T������m��A-�UjE`�1��UZ�ִ�R�J*�cEU+
��PT�ED�+mE��R���%Eh�b԰QbZB���("�V�U�K֋�����Ak*�#T���D
�����XZQQij��+Z�TkVE����X�Qm����֊
�EE`�Ub�ض�E�TF��m�,Q�j%�E���V�U���V���T�,�%E""2҈�Z�[IX���*(�
���� ��V��O�3�is�^�2���~�c}�m�h�v�u���x$� k���_|�j�{z��8�WL��o@{������zՕ�<��n�j���������ӷ>q��'{��f���'u�sen#C˝xz���-�-�^���l��ܰ��y�x��{͋�����E�6��H��a��t�/;P��:<��ç����.F�^�xfc���v�����)�x�{��K�k=��^���W97u��|Vڝ��W�u���0����_t<+�ޖ�<ٝ�л]�{Kc����:�V�ǃ��纤���g��=Rz��g��֫}]Pe�"=8�X����:O�_hOv�}7�2_^\�bU�|�C��.&�+���cv�z����쪟W���_�9��<�>����KႤ��*ǆ&CBlv2�Wy@��(��ׄ��O�W�?V^�C�֥��'cTą諷+=�	��vF��+�,g�l^��JŨ���{kk�e��w��ޑD.�n,�����_'�6�*�o@:�W"�=��?'�^z�w��z.�#��t�<�j��B��w3�,��ۡ�+�Kt1=�f�OK��ȍ�=wR%�̋)��x{
�i�򵰶�eN�&���c<:[y�eW")�Ԇ��{��� ��Η+���6���6=�a���\g�p��5;�w1��J^�X���ͮA��wɅ듲����@g6,9��#>�~Z:j���O^u[�[l���L-��jײ�PX��`{���q��><�������ry�R�S��i�A��?Q�o�V�/k��/o��[?s�^�}�m}�>�ž~���L����MW5�uS�����(_S���v;�}�c��dY�����<�z
���W�����lezAc9�c[���]���;�]����#�g�Ӻ)��y����<{l-�O�c��p�ser���R����S�F����I� y�}҇�{m۬�>�|�=�Ȃ��W�f�@�۔x�?M��+����z�,��ֺ���ޞ��I���c7���J���7���Jw����}�Ky����rGSֺOZ��&��.�K,�gmت�4�P�Lq�g.�%����kp�ƅ<vd����@���'R*[�A����z9e%n����	S�9Z��������Fg
a���X�֣�4�|�1NG;��쭙Hv�7!7�4�'G���rŹf��gg~������;�������A��.��l�{�{,I�}�d��:���݆F7<�>`Vz�B��hyͪ�}|�]��7ػ}�UϾ*�q���*���z���*��^�����T{55تX�N�*���9�'�8J�n/@˖��I�w05�י쿓����z�D�r�V����핶��kh�s�ĖŸ��v�s.cZ�`;���G�\�C��y|�����G��l�\�<���tb�s�g}=�W�M[!�*�=���w~��}��e۟W/�]��Ǿ������bM~=7ez�l9��d��	���%�?j��ږ�vs�*v�����[��|�Wg����~4u�-�.s�k���w�s�u{4���K/N�u��1y�|�Wݘ2�V���V\���#q�����ƽ��̱�����c�WfI=�uȒ咷S,27�떛�ը��N=/fs�;Æ-8�#��jM�=��J��-;Zv���\���y�kC�e6y�������ZЇ���G#K��9֚����,���֤�����f�g�ړ��!ӽ��]4��F5&��3�������6:�M�:r��}���O���y�;��v��[,�a/Fۉ	���g�r��%�>ݞ63ћ�%G:v����,)�X>>�ۚ��kk��,�PzL���E˵>9�熰���G�����B^{7<>ZܺAp����%�Y�E���s\�B��_L�a��3S��ۃ/m������2�d�l�n�~��hW�
/����}N�^�o{G��fW��5�Sٶw#}�=PMl���:�B�u˾r�6_kD�({5}2��ʧrc������G^�y.�`w�sQ��񠟺����z��T8A�˗�c[D����o���<���H+��rz���_�b5�}�{�\JW����c߮�zP��y��lG�G�S���2�E^���}g,j��*f��C�U�{%��M�:����{�wF,�L�Մ��~}�rU�c�;
u��6��v5��`u&�%�����y�*��
����KƮ��ι�WZ�p��uƜ�%�fj�m��} �[��)g(�5���
�V�w.w��	�f<��ӽju�0:�&���~��]��:���ս�������
~�5��8�����΍M�)�
5����,�Ҟv��$��{}4��v-�!J���x�Xߧ �jQYU|O�oeV�� �S���H���*K����=|��O�7�''���y��b�����Xy�ų�rC����!ݺz�~��l�=��w{�~>�F�y6{��,{h��Y�ry��yh��������һ׫goÝ�ӳ�q��;��7���X`7������Kb�Zr��ӵ�j�U��6o�n_�Θ�rx��Uֽ3'�*������;�[v�غ�=�S�����t�WWq�����^v��a�q�N��ϟj�)Oǅ��+��MF7y�m�����x��>�O��׳��С��z�~���m��:���Oa�n�\>}7G����W.<��޳�b5u�4#ٽ��f�]��v9?w>\��D�\��I���,ٽ:#����;v�0�r��d"��W�(X`�s%F}���ԛEoB�J��׌z�5�o��@WNe�aMW�8�o_9�U�s��䖪6�юZ�ľ���2�Yb[��b�ĺr�8�t}�(�����꯾{��)�0~��T������������m���/��qPnb���p+�y3���g��Tl��ub��c.��y��	�xT�$��*O]��wW�Gg�J-��o��/�x9�h���/{!��Q��;�gp��Ͷo_V��L���M/T��_��P��[�Q�9<�K�)�l����\���_/y@�~9��t_9�05�&pメC�V�~�(���x����x�Zw'?�����1a�~9�����V��Qy���=�ע��a�T�'�U#��Y�P���z��{Gǝ��:~0j��4V�tD�!����g��>K�Z^߽n���3cV�Ҷ?Flds���|�9I�qϦ{��ξ~`qmvf�����J��,����>�x�7~�eP������j>�s�����F8�\X�h,��@[
� �3�7��%���ǁ*�}�L�y����j�]�DX��B��k����%�)�-�y����s*�G�"��f��=�F#�gtO�]�����N1Ľ�Ef��Wt5$-���ΰ2or�m����w�҅��)�[��c�uf0NI�Vw�g����  �w��n�\����<�pk��'�����i��/K�:�5Tm-�ck��9�W�5X;Ů���%	'L.s��M��nԵ/�|}��Լ�G��'�t��^���x�G}�8��a��w�����_�0�߭u�xj�����:7�4�Y�M-�e����O��/�f�.or���7���g�6��^^5me�{��!�p@��~�.��M���j{7ޜ����6�v�âC�C��n>)��7R{GX�j3Ɠ��P�㵾s܇)��ϩ�WD�=�+-{��Wt��z�`nb;�CƂ��O��i���S|���tu�3�F[z��|�w2���xXOEU45������^��V+9��.v�>��v�z��� ����W#]�+Ka��{����e�j�ìz�3�q��J���#�gs}�ٺ�ڗ�Bw�:�b���3�˨,�!�'i�dz�+��`�h�;WQׁγ;#v�Y�D�i_��<�}<�xO3Rhy��{����f] iY��|��:;��}A�|F̌L��yj��YS�՘.�Na�������G�B�rW��Υ��{��Z#�˅��X�%�+��~��_o�|> pZ�����ǁ��R�ʹ
U��Ƣέ��t���Ě�|1s+����ɱ��������|�ᴢ%jU|��z'�[[x�J��B�݆=���+�^t��c�ۜ��x�_���4f��{��:���fb���m��:�gd�]��z�z�?s[���7���������/�B�Wy��3G�.�˄��o[�����n�=��|kme6����]����Rb[�s�=�1+��L ��6��IaKP�z&�����9���<�N\R����~Ώu��'���s�A��#�[�Yp�\e�������Yg��v�u���_L��꾫uT�X���������9˱;ORχ�hs�}L�^�o{�൜Nȼ����z�/FۧQ��g��	淋
�x���͗�;�Y���U�-DP�~ə��-N���O�j���j���U:�	���*uw���&�����Κ<�l.x�M#7<,�w+��o"����.�h�tD���鯀[�Kd����O;��b��vSí	"B�ñ#WM���{���ﾯ���m;�(����j{�ʽ��>y.+\�z:����@y9�P���\缠��Ѿ~�ОG�S��A^���`��X�MẊ;�6��>ol�O�뫩��^��}y�wH�詋�!Ϟ�^��JXG9^w�>��`|���3dc�ب�%�[���y��ߙ��Zf4O�8T��1�+�y�/r��OPL���E��r��dXk�Զ˪^\//��++^V�?TG�x+���K��
�;�g-�(ϵ�b9�z���#�E��g��rS���tO�]'<i�n��C.�u\=Uw�M��r�5�<��`��������{�����Wof�,�}�^(O%w�nk.�le�!����yC>�� ���v7��-+�����ǌէ�C�E:Ǘ2�em�8��b�y`.k=^�� [Z:-�+�w��؃��h�/�{t���քv�
�xS��&N��fA�
0���쥯Aqz���G�k�͗���K��B����t�YN�zI��e$�a�B���[���.-�ng�����_X3�.�g�"J5�*/SW�z�>��yա2��O���r�vtL<�$���z;��՞vr�Il]'54���Ⱥ�W��r@�nf����rY���7-��N;�jS?�|�}�Ftkzܺ:���a��`��M�?rO�P��w�`c���u��= ��\�>mK��^��ה���w�T�������\k����i�X.�e;���`�uu�^~^Ms��̝0�f�<&P�,
g�e����+&�r�Dx�G��wWl�74S�g�����(����!�bZ���o<��L�F^}3�g�����r�J��84嚃�2��D�2L~9�Ȃ�З��VT/�I�;����߄ژi���|�*�nzR�99J�nX����Cۈ�%����|߆��P���lY�S�Z)���+�}�C-p/j�iC���q�T��|���U��ʤ��2��K�G�o�l�<2�+�|����A�O*��$��t�����L�ߪu���xc�ͱ^����im��i����\9�H����.��1�3'�S$�t)O�c�E�,8)�,�;G�Z����L�=��=��,�B��WQ�v��4���^�B�����U�W'K�z������G�����/`���F��Z�y������Lm��Q����tTn1"�)w:ٕ�Q���:M��,
��f�^��Sx�P�u�oVܾ�.Q��_d/�劦جON�C\�'@��t!b���<�4+����{m��~���#�}ϰgN�u��O�ϥ�wC�q�S����<�_�PV<w�9�E�λ������@�[�YA���CKU���-=�#�f�t��]�
��Q�3��Z"�C
�]��ucɛ՜0ᢚ�����4't0���I@�zv�ѝl�7w����˲��Qye��v_]%K�����HG���0��uZJ�ǡ��!��Y�
��X�餃E�;
����ˬ��Yԛ�/��G[&�s�o�P�yЧoy��#-ε�k��xFu�lSD�YMI[*8�:�h��BC+C�6��%�5�l���i4�1f/�R�9¸�y%Y :Lo5n-����A��m�HP���6V����9���\�*�gyrʅ�C2����t2U��_,����N�hL��K }�e�7��Ѹ������v�.՞�Yw���n��~�`ƅ��M�E�ݒ�ݎ1��u>����
ܻ��]�oD�ٙ�Ԁe'`����)�k1\�heʒ��i�aM�[%��ۨ�ա`��[�)v�ej�7*]�sF�}�+,ˁv�s����W�#�cdS���3Jj0փ��ꖶwc��X�����[�&Ȇ�d��I1�5�m�agn����{ff�u�ӡ1k�#��N(�o:u��kVŋ�Y�q��5 Z�iv�N���JJ���6����\W�L;�^���N�폩;�S���^L�׷@���t�:�֐�L�;�#p�v�¥�[�Q+�{���i�ٸJ�Pm%}�w����7�-�|4�Z��^_i��
�aJ�v��ܺ�y��.��3��:�V`ꏎ0�V˭9����gkH���g+�#��;2�W[��pր�==�".���i�6��Y�0
�qf*	^ɴ���:��;N�$�w�K [��Yt��ہEpJ��U=���Xރ����*�u�5D��֣���1�{Ozu��Sf�1ʄ�ٳ���)�hNT��h�,����<)�)N����F�������읝��1��Z�B7Nnv�H�!�X�(r4���F��w�Y�+�U�N���-�x�`q?#Z����C�˙2��h�cO.v�a]>'Y�=�I�ξt�*���@�����ْ������
�8@���Pκ;]}O5���YjK�xj4���Yt�	�7z��*j���p�x��;�&B�)N����� �ބ�\�v'�i�K�h�x������و;��)C��|���{��ݴ��>�}��mj)��
�	Qm��5��uhF9�v	y(�;�5��xK�*6���a���5�}��(6d4P�v݁o�ޡ�{\�)^�}��酌\�3��s�k�)i�m_��)*Q���Z�Kh�Z�k
��TmXR�UX�V�`��+T�T�*
T�ֶ���+URV��D�+h��J�XQ��[m-%b �)b[h�*��m���E�ږ�)j�J����"�(Ьb�`�ҠUT�*-em��*AE�(��KZ��aDYE-�[Ub"���(�VQ�b�6�QEUUl��R�
�V+��Tm��%j����aQk
"�F#iQE��UX�#*k+
+AH�kX�����J�
��AA(�E��H�F���T�X�6�a*��lUPR*�B�)��X[T��I+*(V�D
��,P+*���mH����ңj��E�
��Z� #Q�J"+��[PX���`֪ŭO�o�k�	��:�=��+O5Z�V�$w�r�.�����4�<�2��H�ޡ��z�4A�pw�]E� cՖ���U��U��Y}���z.D���,�}��Y��;�sմ�.����`J�V�~~P��Jy��ݱ�m͎�3����QAV6VG��b|D���"}����!W�w�2��/�X�V^b����|�,��m�d��T���٣l��v�������ʲ��7��Y~�br��U	�ͽ�f��G8>{�3:e�m	$���({�7����?@�����������5��ح��C<"����Q�9)ۊRXӀl�~O�.��g�p&i�g�^�0R��X�(u�D�k��h�t��c;%��O/j���s��{����Le�������#`�z-�ųX���]�gU��ٺH�*��z������5��PdXنǟ��y����*�����u���
��e��ݖ��CBu�h3sy�u��u0"����n����R��s��L�=Q��ly4�R��)�c)�/+��.v�ru�1+���;˨��YŮ���Y��9;nbm��R~]�)�E�|�p��}{�	�xk0�5[���r�&�h��aU2��4�vV5��yY=+�#�x襸�����rm�Ɠt�*S�b�4o8�P������nT�Rt��%�]kz�+ni�_,p��Y�1�yOk�}�pn���H=;���b��B�b������}�MAy�=�w�j����.���K"b$N����<���>V7ƙ�ն;(j��Ls����ࠗ���E\��-�CVx`P���^fw�^V��Ga#�<�8�~�d{�z�����p)�;6��f�X��(B�I��q�8Ih��t���n�@^�;��������_q@Q��C�֍rd��Xτ��%X����+�[.]�uw��sA��޳��֕���^N��A��Zg�z����4�鄫���$9����� \��g_�S΀���i��Ҕ��W��-�1>4�ؔ�o���-����j\���)z�Z�Lc�ߪ{�E�^{M�S���ʥ���a�B�f���+�,2/��>7]x}%@�<�j���D/��]o������#�r���W�l��Pi������6��eK|���jm炎��u)!J�mp�K��N��K~ZcP���2���4�ϩZ����J�2�U����|V���$�zS����&�ql����'�-�Ϛء6Uo))��x��o��o�݊��[�f�ɭW*1�|��D �[m9;UeI� ��ɵ��b���[��Bn����|�'A�Q�+E>��j"$�������Kv*��8WF��Z|������s(]Z,f"�<��qZN�?WQ�z��|>�|�}=�yRJ�{Rj�Eqn��yUF��z�k�[��/��':/3�ja<T-n��z뚱O���?+�!��\	=�\[��g*SՁJdf}��w���Q��Nγ�d�7~6}|�4�
e�m���"�Lp����>��V��=i��by�J�m9���7��޵����K��Nwf\�Ő	��0:�L7=�ɰ9�$���(8�*�}����R���=/�X��>~R�C�Ń�6���n����ŀ�:2��s�/��z����_M��Ӌ3���`z"�rJ6�3�,NX�/�r]x@����OZn�3�Ƀ�y��e.Z)?���ŎE�	y�����+�}%"<{�hyq/xx=�����i��ܩA����r�&X=��R���j$�5�t�K����ٴ���-k����޿z�M����&6+ě�H���t�W���v��3�۸E�
kG-g�o)�a�B��\������������u��u�/k,�a����O4$���W����]E����Ջ�Vf��r�zkU(�&�ޥd*�{����ɜ.�&et��� �V�^|���0��P^�\L�Vn��|�n��'Ax��-��.�}:�k�;���I%ݱ�]���[�b�Q���ޑj��[�\9��:ԛ�������GV`�~��Z���r��3rƵ�@|m�[&_����:����h"�1��P�Rv����s��ŗN9Ά�����Q{�G����
�=��-+����~�=�)����^����7}�֩ăK��bϫ��X��"8��O�����x��-� �~D}5~F���B�WO{^�c:�\�(W
VH�������\�63���k����91�A<���o*����(,�υ��h`\hi�:�EJ��M+j�7|{K��v��*��x�@݈aϔ���7��釼C?����5�JS�+"g�e�K��ő�5n�r[����y�0؛�,�CܸH)���G�>�d۔� ��t/����(�b�bٸ�_�`�f�H9�u�G�i�|�a����ʄe����exo��P��#/�w_M/M�c�I(;�?iIB5��-�/uģ#����X��wֽ1���=-վ�]�knl�=Hp���@�:E�T�.����K��KM�槺�ʅ��>���}�VqF�-�
g��Яn>qܠ��^�s�w��h���j�2m��r&{��5�'����n��l/y�V;�&�jY�%�3���f�tB�s*๧��K\0r��L������xc�w��|�T/����]L7�H��.�IѱY��������y����-��bit��:u���&�g��:<���]�f�R��잩�)9Hs��Lp�{9x����"q�O�ϥ}r��l:�lL+�_ԟ/]S0��Bq�rO��T�쏽��7T��N����R��qQ���Rq�>���f��'��Zh����.�i��wjÂ��nO>��}f��rf��^�/ޖ<�{���ˀ�XY��#�~��DLC�x���s�8巛������@ػ�	�p�����u�,{����4�,��C�K��8:�G��Ζ{ys,�}#�h�*�T�3>�[9�MZdGn���ϟ��?3��s�L>S4E����M;��������%��
���v��:��q*��`����w�OiU폳���#�������J������o+�-�����xW��e]���b�Q��I~l��Zt����sg[�~�%�ݿL��	e3�^�C���v�4w'���u#Gۺ�,�a3���]�� \�>N_5�����9S�y.V�h3bϚ�o�z�9ܑ��2ʓqc�=k(vO�7�4{�N闘MRSp��p��*>���33c��MU��]C�{��y�ꗉMf����sr�,�N�ń��%η��i�(˔Ǹ��ek�a�Y�_���>�  ޢ�xˊL�9��2�#���VC���tZz�����g��ȱ��3��V���fj����{���|�#�eC�e��T_��bC�yeu�����x읍p���Ķ��uɣ��H�A�̠o�K���qqR���tT��}gqs�䌎5�����}��G�%���>�[��t�ޔ&�9��7�R��~���*�!��aj�/z�g����>�?P����-a�L�#���엸K"b$oJ\UҞ]yv%G�=-��xs�24M�.V=��β!��~[!�<3�8��6QC�l7&rcسu�G]�X��Xm�3��깒�-a�=)�|B�����-p�-�-C_{iv��������$�� S6�5��Rd��=^�wKIy�AzKV5�����)��{��uf��(ˍ��6�M@����PgEmLL��h��2Ǻa(���9�w���t���yoa$@��v'��Y���}VXc�R��7��Z>񗉎�O�HIϰ3c�<�/ud��S*VY���[�wh�Op�_��{�����Vc,)��
�d$�w����.}���M�G]8\���iΒ�iM�3���Xz)��㋻e+�v+�jR|��l���뽺�E��Y׃F�V����b��}��}�ɫ��a�I]�w�\՟��9��X�������Ұg�S���R�/��w`���7"��&�9|���o����u�^:\O��p�h�z}�G��o+��Ic>�<M#I�T�W��l��3ތ���(W���\�YL��NfC�t�������_�����JmJ�WK�[(�Z֫�P�YU\^\�k�ꄛ�Ų��tb��!3��/@��BjG;&:�}^w�Ӿr��rQ��YQ�/i}qyr�Q�o]� �D����|כ��i�,�ž�5tL��ӫ#������:E�C���<p�{鍓]}c㮷E�5y�L� �T�%���Y�d6rd�;�v�eQ�N̠E�GI?(���֙��cK�]�F�ݷg{T���ei�����L��f�6��:�L7=�ɱΑ&�!�w5�=Ş=&i��&�.o�R�(8;��.����KEC5c�1u蛐ᕂ���jH%�P@�b�]���x�Y$حG�+�3bb���ݔ���خƜ���2�îж�Rɂ�����F����tn�����4��C�'�f�:�Z�5��|���oA�����fc[J+U�Zؽ*\ֲU��оɲX��r9Ǻd��T������a�ծ�b_�GAm�epyE=u�)�wjӐ������}_}TF\랣���L~�m�H�O�.�9��(wΩ.����]�s^*�=���	��U���ߎ4E�u-W��s���%��^Z//��S
���e���T�@lk�ĺk�q���[9{�Qi~D��d�����ͼ�����ߘ�Ԣg=�t琶�v=ob��O<�ӗ��A)�{����G�᚟���[3�(��������I��}�>��M�n�Z�Z��Mʡ�}�֠��0>��[K�[�^u�C�|��ב��x�i�-Ckz��硏��d���g(}�������jp5���U]��O�}rG�ˎ=O}絿<���0ߩ��!
އ�d�x��"8��O}�\Z�Vr�W�罧�k�ɐ�=�)��=U˶\\Vx�ȽH�)��_�)�|�H�R%6\#�V>�ed�u�o���@��C~�j{�A�{-��C>�6GRwIVz7�ӗ;�t!�w3�R����\s 0�bm�K�l��*y�{��c���'�5�f�wB���n�4�3י�?t~���^R�
�5�ۊYX�u�VW!��W���[����y��7�:�q�f�M������3����b-����o������o��z��u}�	�����A��WVGh�6��%�N
��Y�P�i�F�����.e��_N���{ sz>��*�����Ko{���v��T�%�C7����s�2��`
g��q9�}�ɷ)4^'�ibqpJ+	���,6H#��u!,T��y6������wg�u�74L�ر�+g)�E�#{ݸ��\h۝7�(�K��K�x�G�*��W?�g�3�óV.X2Q��7�^��[i�$.��3������ѽ�����@��iz�qw�]��6�.��-6|��V�ۅ���S�A��U���b�97�V�<}K��n���N�8�DӬഖ�h�K�avxm�z��Yzߪ�����ȼo_�Ggΰ��j��pHi�8%}bU�X���+�]'�חl���/Cهf-f�{K��W�:W����J��$Tp�L�O�ϫ����P�H�^��m�������ҹ�����:s�h�ZO��z)�PԼ��
�̀�ag�#�|lzoe�ǧ�=!_OL�VI^�<s���
�ۊ�\������	��S��:�}���^��KN��d�֯"�^V��BVn=e�5R��c��G��1> ��~�Ϋ��2�+�����컧�vQ7X0��1Vv�0����C����F�u�E�#���wP���OE̔�VǓ���������e0��U*�m��w��%�8Z��E�ĳ:���k_ZV�����},��݊�v8�����%�qY�Q�%S��&ќ?|>�}��o�W�����P�$�;��׹B����=e����Lp�){�f�:����,��v_pH>��=��Z�r����?!�c���({����y^ym/Z�<�KU�*��7�TG����=+h���Xf];��.PÓ�ڹ�{�g�q3L�/R�
q�����:���Y��!0��.1*�D�}�	f˝P�N_5��W��=1�r�+�o���G�e����Y�PUW�TGX�|U�OV�Z�9�qsY���,�C%�!HSu�?B�����a��)�
R,YL�Hg��v^
�؅��t��̿o��[�y�.h�v=y�d�v٘�ƶ�5�ު���41961�}&���Z*�;Ϭ��X�ck�,n���ᶏ��֟���:m�B`Bzz�PrW�'���L����4+��wl��{=]uҍ.P{���Н��j�-:"f�]�J�	���)}�GAh����t=N����u5���9S�ג�����W<9��5SWHj��C�K���FW��:�Dz37��s{R��4G �R}f��X�nuiT���Kz��}�J�a��t�{�cgޔ��镣WA�#�]"f�w�Wm2�|��63�P�@��n�*�2pۻ9kA�X>�7�����ΤC��v���}����*CX�k�	u����9����PZ�6	o#�3��)�޴�n�On��E-���^
TH�*u��;Z-��e�F ��Mw�]���b��]�-M����t�K
��pݛ��8�u5��e���u�8L���)�\���gT��j�	��p|��|p���|s���_�:�E��Q�r����x ��;�����w�YUk��4�	�X���pm`sVXr]�y�[|W R�{����飕=��IY7o��J4M\�����b�!�3�@R���V��c8�SԫYYd���d �JLwHkow�א������g,Щm�5��ak��ӱ`�@�;s�]�K�GL�n��������U3]c�K��O��kx�/�`��Qv3��U_;}���WQn���`ֳ�p0�۳�W)F����3T��˓S��mG�v�d��!Fov1���#�_7;S�t��8�ËM�ٷBb�VXٓ�sE�G��Њ��YQ_n֞k~�������-�͎�-=m��b�T���
�E"�mvU��dS �k2��.�w�q�����ZN
�o*N�b��>��(w�������y2eK<�t��i�wv�ۑ������UՍ�V��C����ɘHV �]��{���Au/���`Mp�u֊BM�]���i#��o8c��G�+xյ�!�6�g:��̌��w���^�Ch(f�Ժ!֥ 
�~T��w��+��J�p�vj E�2�����#ml���`�ԌZ���j�3���v/�w}5Ӧ����m%J�.�w]v��Km�E��leh#�o �(��_Lɭ�ҎM��.�;d��n�MjCP])���-vW;νx흠�v���*��k����Z�,lښ�������g���.+�����^�97f�N�����Y˝md��DT��(��e[U�WL쭽�+�F����CTa��[̬��X��Y����z���̗G��nm�u�O(T˿�9�:�WC���ѭ��b|Ӭ{��'w�J��3�K�J:���j��&�	������G`s��=��m��>h�P7�ӭ��fa���̷�b��]�mD��8k��\����_[�0.W]@s��vU��c�j�+Q�	٣`ت��`k�b�-gz��Q@k��C-���맳n7`�������Y�aCle�	f$˵�ҡQνi,��{o6u����x�U���X���z9Հ¬����E6��w4��^�N��\��NK2��5y6�n����-c�gس���c;W���~�$|A%%��6ȭ*#h)*

Z�U��U�T��Ŋ((�AeB�[kXE�F�XV�Tb2ڪ,���-�kBڶؤQRՕ	mF,E`��U�("*�(D�eJ VF�F"�5�X�1X�VU`�H�ڠ�-��TF1PF-J"�X����DVD��,U*,�cՂ�b֨�X,E`T���[X�DQ�Kj�R(*0(��1X���ֱ�T��kb�,Q��Q`�"�J�YUVU�mXDTJªY(��[`�����H�k*TX�R�""�X�,b�bEc����EPj �Ȩ�V��X��Db�E�
5�+[h"ŊH��Q�Q� �1b���IDY���UdPTb*�,dX�¦G�X"*�(%��DX)�*���J��PBТZX։c���+���ŗM�h

Q����J66��^m� �]o1T��|�f�gf,��P0m�oR�i��U�>Ͼ}�l:Όפ�"�#�:��k�m����k�Vf�`��7P�bL�����Ih�β�9�ݘ���zlĚ��n�����f��yɒ�_ر�	[�d�pXRP`��-r����nE��w-�a>��t�������/��A�[S=��=�e,c�ߓ�}�{p����k��%@5�E����Q����t�=�ac�L8|�h�������h9�m�ug�F�t��Ύ���ܨ��<���{�S˕KSӰ֕��	�m4|�9ھ�Ylym�m�.aD�߁�6&,n_���>������r���l�QA��j�wd��ZJۏ�M���9"���U���B�����>�C����ut��#P�\�~Ѽ��}C���	;�����Yȕ�ē����}P�x��V}��BN�8-�y��ɔ�5��+�|Տ2�F���,(��v�jc�+GJ~lt��ćWʺ̫��V6#3̯ͫa�V�ft����ew�}�Q�ȵ��V��s�pbs�g��#GO��x�qM��c���cї��*��Ò
�c�6�݉L�&Z>���D�(l��|��"˿xW?�X�:���#��_��`���[�
8u���\Wm��0�D�sN�v�p���4R)N��{nt�ef�]�&���<��}_UPڸ<������"�;%��ﳍ�y9���s������*�
� vZ�[ܐX��F-׸���A ���vl����0�?�>x~���e�x����a&	�VM�t�9������2��B���g<n�B����h;οyb�p��/����P�R(�OG��)K�z��}���6��=�����$�m�d�Kµ����u�Ogޕ���DWcN	(��CJQ��;3�3�/|��߽����Ul�`
�`fR��Rt�e��/PJ���+/�X�+}��ٙ/�����`�^N~͂����^�0�Q�c�Dp�e��>y����:�vLkg������"���.-�m�L�GH�6�V���CڔL�w��$��zP�K���ȩj���y�S>*��Fߣ�p�O�`��6g�Q����/>�i����_��j�H��=�u�}�`��=v��Ppܱ�cP�M.��g��ΰhu[堅/�Sb�M�<���K|uv���^)+�a/���b^��pWU�[��^L�/�{��c�% �]#3%��u�ⷳh�@Pa2,�۽���]*���2��@bj����gd6b���?+���V`�f�ý]1<�f���U�y����� ����=ջCk&�MD�Ƚ���u�M {t�N��e����gz�+�hI������ô[���y�[n�
�1L	�V�+�s�O�FU� ;kGE��v�ط'��`�8=[�����.��B4��l�=���|l�/R;J)^+��`�'>�D�Y�~�[�%xnZ���@��&�Q���5=�!�w���C \hi�:��J��]�x�9�)������/��rS���y�1ͱ� ��g~�<�D~�/�(�x�R����,�b�U?2��e��˰��V5�3���bo<�-r�3�'nQ�>�f�����wyq��:,�)������C�A��T�Ձu6���x�7�ٗ�fO�`�[=����o/e>�����oOR[fݗ@��I�uP�Y�xR��W
�EgW�f����)fgF(,E�\1���0V߾��3MXx粁q"��J��>���h�rZt[��0VM��q�c��Q�z��o�r���̥�x��V,Lkn�<�rMr����Uja���?g�wʦ�v%-�o�w%�Z���yՆ���&�4��	BJ�"u�ؙ»R/��D4�VJ����)��k����s
p�'q:��U���y�I����O��=�=nF��؆�f��];u��*�c��<���9��{'����q���ˊ���u^es��-w2q1R�ނ���W6���d菾��]n��VggF��]��8�����W�TӋs�ü��Z�^?���Ff�`�����LpS�X#�}jb�IZE�W���M��J���v��w��͓����<W�a��,y,�b�k��|��t�z�������P.�69rL�[B����xm�S���,g�'��<�S����s���|���(|��I��60?�ob�=�Yp�K*�+�VG��O�+���:���t/�3�4o��K���FN�C ��w/M�r�r��O_Z������Wr+Ϋ,^b����,\��N۶ޥ]\\�3�A�c��?�~ˬ�S���4�*����pi�3W͕�OǦ���sS<���bu9C��p�o��%�ݳ=��YL�ggl��fkLj��
rS~Y*��(q�%�����,�s�	�柨|\�����^��ڝ���JOQ9���g�$t9L�W����Q��C�����O_]� ���(�]=S
��~��6�쮊�g��lG�k��X��貂f^;��v!i�M������/��s]kkf�s���4x� ��i����Y�7���S��/�I>J�wswH F+S��`Y��e���������ݸ�8�R�37����Q��j�vl���7z�t���jo%:�u���0E�w�}V��W��o��l������.j����ޒ��/�e��ڼAڱ:��(�\�<�tT�y�����x�u1o�n�!׸��-w&�O�ʗ�0	\֟fgٶ�`3B�Ѐ��rZ)?IB�x�d�KȜYo2<>^�0f��6�;+��6/ǃ�'G�Q���j$P+�bS������c��{d-���W�x:�G�7�Cy_�w����5g�(a��y�a��%!�D���k�K&PR�Y�ᎪK��p�؟�6��>���W8\
���<�N>��TR������B���1[Vz�P��ܦ�y�&Ku��d�YާG|%���,���Ozۭ�ﻔa��`����
�52�1�;>(�u�>g����y&��\�h�rm�6�F�n_9>|�?[$�ͽkDu�3}})O��'Q�.��X�)��E7h"����|�X���T`����tn�?qiy�6�;��\�\����D��hh�B�6���L���
T���n_���x�q?,���/O������n\�}X:����lgc{D6&�1�Xz��8i�U/�$�q�-�l.�����R��J,:Ϡ��=Y^������3P,��z�_S���/*j"�v�ۚ�c��r3^A�(�M�_>��jr��g
�%���[ �]�B�咰�K��T�y*+.���;w�}�|9oL4�M{N$�4��_�
/�0p�Qu2V)��t.���ơ�6�z�i���z��q���&~pu�i��Y�IX|e$�zS�������F+���$&�N3�Gv�c[�1̬�j8)�5�(|f�V�%ڰWU�����r�Q�o�t�+K��b������Q;�4^J���W{�D~V)hCa(�iw��J���v�������L�N=������-�J�3z���8�σ��|w�B�\�=:�,��I�OQ�Wj��e]>�4]m:Lϩ�Չˇ��K����s�2[՚>�|sh��,�(�a����O3�S����S&㬄#[�h<���.w����EC5d�1vL�l�My`ɦ���J��=�
����^�0&#��>���per�_�gޕ�Sف�WcJ2MB�����g^����ū�� �EÂV�%�f}K�E&�X����%u�;�P胄�HZ�����^��k�5w�[H��JZ�I��o�m�P����Z��y7VxO�"�{�,��)�x����g�����N�7��8�VB�jp��=�P8V߯�A5������Z�MPlV�<��u�:��]�6Yx�mJ��<'����9A��z�l��9o��=����p�ⴘ	�Kn��PO�~�����b�ۖ����U�s�U���n
d�:Gl9������Cڮ�3��f�9)�v7����!!���f���^����v���,��6g�Q�lZ�ێ�{a�O]��M����Um|3�b��Lf卋������Y��[�{iܺ�$eM^⮶3F���#��̞fNl?r�JK�痃�ߨO��mP�]3���iy�z�]Rx�w�d���#�`����;wLh6�<u�c�h_T��׌$�u��ui��_�p��3����'g��O�rߖ����߯�F�K� c�;1g��AϢ�	�q#\�6}B�ZfUoiN���jS�.);֪?P�Ƨ��a���{��<UAb� �{so����'����G���_�z����c�c�Nv3��W�����ht�`�t-�~9����3��L�"�H��}v;>�|��g�za0��ve��O�3�=7��n?}��W�,[���`�KȂ���.���ڱu6���/f�=3��²��˕��2�e;9���¸��15y�8�=�C��r��%E#'=u;9�_�ԑrɂ��]�u���Q��7�Vɟj�96��U�59�k`b�,L:��Y�W��>ޥ3<�ɳt��G�C�bYE�w>+{�V�C|ϻ�皯Z��<[����]��ۙ�&���_��+ge�6�&��C� Y
�e�v�~Ypz�L����6D�E	��&fI�Ajt²z+o�s�{*��dT;Ď'>^Z9��5ڠ95���>mc?I[��P��;n#�h�}�>����P�U�[t���� Y�/ۙ�}I{&����ò�1�|�eQ~u�ϝ[D�S�b��K�"�>�]�{�[��0�Cف�M��Y�h�w۲�{�"��i<wEzX���Qό���������Z���3Eu�3j,�������������ͬ�x�G�����[�~�`:��\�E��)*�r��ie���^��<��!V]�B�V=9q�>x���]�<����x��Ac�I�%�XDK��9n�@X`K6������˔j��yX���9���x��_ޫܥ���),���Z�2�E�X�R�x�yc���~{4m�B]n��B��A�G׽~�R�Sqr���(�>��mqpS��c��6;���d�_m�h���K
�=s�&��YI�lə~L�����'�Cue��}�������lC�j��#��y��ָ7z4��]0�ȋ;mw*��#(���\$v�o�	�/���˷s�2���ak��ʄJ���+�:ʳ֍f�%'ʟ|��]]�EW9w��2�zy�=��`��վ�}�P����N�(t'6��^��s>�\�����hi�e�-�WVs�:�TN#�EV�t�J��xx�<�^�l����[�+��h`�=��eV��)�+�W�ȃE��3�#���Vq=Y��V��Y��e���j���qg)�S0���c����k>N�b�L�Hg�ݗ�U�Z;'�G���WgjTh��\�o�t�E���[����u"�=�@�ip>�:��P�e�4�)�vY=���0g[�Wι�|��j��~3%sZ|fK��]i��	=A7��J�?.��u�z�$�#�{����+Ơ��%�t��{�����O2��0�^G���Yd�j$-��9��/ˇS�+w����+*}Ku;˱9o���%/+�{�񳃝lA��]�-�՞0�=��a�i��^����c�G�
�Z>�3�]̕Ҫ�,���IXn�
��`��^��H9 �o�T�7:�]^",{Lg�r����P g�n�3,f{4�-��)$
|˷�uy[��撱�Y��jf�$5���<�F���7f�pob&�0m�����XZ��z�ηi�t妡��f��ݍ�Tg��@�?�ꊁ�g���O|������-T��ٺf�`8�5O�$:����^TT�v۔��;}}RI��thE������r�ۙgҵL�'|�:�5v��&p�*;]��ȯ�ݮx��iw�xJ���$��̷�G^僦�����=A1�خZJ��ά~��K�	0�tg���2�1��GcҎ�����ȓhn�:W�`5���άX��jɯK][,̿qs���*X�ȫ��Acr�����/�������r���E=��X�<�ݐ�^zy�'���Y�U�O*��W�P�}A�x����+�d;�]-�|'t�)jMg6����1��Ӈ�+���rRV���T���ꄜ<[+1�r��W>�sN�sw��������g�C���
"y.Ĵ�ڊ���ĽĀ�����(�3M�.]3�3(�bl��P��g���V����Z��I�Q���ԗ�e7X��b� �]�>N��]��=�q��'=������G�ve/�Y8�*�/.�67�˘����,��}]SV|��|����bNyf\��8M�9�:�L3�aa痛�+����*�ɩ�;QL_p·��WX�
V�ڳn�<��;��Ũ�nɧ�y�}�e*�w����p��]o��{\s;~J�R���*+�umv���,�"��� GÌuڥ�b�Y���E���e;+8��������ec��&��[ލ�9�@	oEގ�tޜ� p����G�P\/��nax�:� ���k%>�2t��)
�n���ػBW��\W*�jp:UK��*;k8�ZujcS�gD>kl:w;f�MZr�n4��e2\&*��G���2�[G#�1�l��Ur�V�S�] ��6�f���� �TQ]��'-*Z��������SY;U�������z3�����[�%S�k��2�͕qhW�3��*�Bp�U�]��NAs�wX�q�Y��.�8�H/��<,+!��M�S���h�i���
$��Wk.}�)'��.��\��%Zs�e]�m>�:z�ܬ�%��R��-���D�N�DM�f��F��T/�	��6�z<!Tݍ������kQ*���x��x^`T;v$�gi�{¥��7���������o�(P�+_J��F���'��.!Y�z8�[T�R�R�]=��zc�{�enESNs�u��sz�G3:p�f�rm�n�Mލ� � �d4��Y��}u���7���e����4�M����{*���j���p��%sl��D�/<;��S͑�Te��&3.N�1��6�q��x��#SUX�ăy]v* j�D�;�w&t+�Z�yw̶	��ʩ��]e��4*��Z-��pM3���w��1ϳ⦘)Gξ�}�O��GR�w�U�Z�<ӕ��T�ɝ��1��Z�4�'��ÉN�ۘ�3�0/��(3iCB���n�u�/�S�¦S,��;�F&��ɮ�^Kz��o#����^�i�X�+6/���f��㋭���;�W{��:=BP6�.!��p����j,[��{)�E�,�z����W+8V�H�P܌F�c�f<v>T�+˻J�Q��ݑ�Vj��A,�ʷ �ȇ-��g'I�f|,V*;����I�5�:ue�K��9z�$g.��n�/fCj_#}�ӌ:�aWΒ��elN�UpC�$ڡ��Yk���y���'m��FE�.֖��Ϭs���ݵ�
���C`3:p�(����^l2�� �Ye�.-�9�ީvɜ�StYi$��S5R�	Z�����vX\�p����2�j����K�u��Q�U,wR�2��mL�o�^m��w�N͉z�ؕfJ/
�և+}]%����D�[�_lY��c6�澣�;�����X�v#uc
n��q4*N�u-�I<�Wk9eb�[n�
��$6E�.I�%X�!f��]��n��V��ࠋ���'�ɮ�
[����D�3X�n��D�����i�n����{f��f.���s���9ϴ�QcE�+���ᠠ8J��UPR)h��b�H��
"�c"�Z[*DT�ZR,���1naQDQD����["�DTDb�1���PL5QDQE�`c����XԨ��Ep�VU� ��
�Q-�Yib�ڊ*�AE+C	QSZ��AkQjX�Ak
*�%�`�APk1���5(6�QVj$TV���),*U�������UD�EUU�VҌ���E���V�akTU��*�V*0�j��+l�,QUc��X(���Q`��Q�@QV�EDA��-*�PXւ��X�E
,���T�%��*�������V(,��VZU���"��[A�EJ��""�,TH��WT\5UFT�#T�TQ$U�(����*�ҥD������������.�}Y�����>�p����⢕.s�_>�E#�ݺ��L"�X�}����S�R���t�gE���%d���I����B-8�w�~������R�|^�C5d�1vKtyW�!��Y3DE�_em�N_tڜt��f��t�
�X����8�p��_�v�	�g�(��k.m�nT�:���ѵ�7br����*�jϪWWT�Z���T^�9w;����%}s���^�5�RP�\{Wl�JDxR�nn`��pY���{%���맏�V��X�hr��m#�� �]�2�;��1�l8)�n:Gmͼ�t�W����M�J�z�Iu=�'{:�������5�)O}����
6��s�5?%"=�=�����x���^�r�K�\���gq�U�B��]�pj��3��|���?o W��ȶ���@Z��2P�V�{L!����W���+P�R%��/w�f�w]Z�jp5����Öx��T�;�I��;~���w�S���O��z��%� =�A镘jJb�rT�l�%�����DO�D�=}.`�8S�E��^z�.�4�.:"�p�<�oJܻ�t��=r�Ts���}@5T7�-�vwaC/�kc�]�wxtvI��sVƕ��.��m���gDǸ��IF]��O�ɺ���ȶ��cX��dú�'B����\�7�5���Q�w���ͧ�~�>��v����������Y���s�M���6q�����q9����r���6^��'�,�C��7�Q+�P�h�L�C�	��tz
�u��t^	VQ�f�����f}��w{-IZk�%v"5b���|��g��	���yg>�CܰIK��O^��z��,^'�"����۴Ky����׎D,{)��:r�27�0�w��~�p���j�(H����������g���@�r�J�沂d_�=6�(^�.&���R������{��=>M��-jbe�k��Xy��ċK�+������K`c�d����� �M��9�=^p�B�Z�s����#9T��3\���G�ߖ�So��§��{{ﺲ.?o���wFc�0�|�[D䆟#�}.�Z�hG"ͯU>�[|o���GԎY����/�yyґw��(ᖘ.�/Gh���~����:%�^�^��� u���S3.,�ǩ���&lZ�����%��X��@}$��m&�"��p_s�7�X�SC�R���7*�{1��:S�TՃ����4BŜ��޿`��=�X��{v�Þ������W����
[ų�)Ӏ��IOݵo������D��uK��:�,��H"�\1}���Mf����ţ���>{ژ�ϳam�BY��̠|6�&xeLo����֠8<��X�L�Y�ǯ���X6V��h�O��M죃��֯5PN���f�z���͇�N�֌Z�6���e�=u������2��gq��Ü�o��NI.���5�A]�=��#9v��z�՘�����&U�ٙNf���2u>�L���39U��z$k���ix����.�A�8 �K���2ר3;�w9C�',i͝o��%�ܮ�ɯ�n���fAk=yR8g���Uz��T8��(qf%����k�Y�\���;���9�{�CW�$��s�q�*b�p.����C�$��HV�K�+�z���9{�MX�v�KL��������a֣Y�+�#>��c��.0�#���|gʏNHvRU��f���X��r�e�hݧNY�̨Y�M��׽պ�Aڱ:�z��ɥ����B����=�wf�gC�J�ڄi>u1w
w�2W5��@�38��v��	bz�WC\��.��s=uf�+y���|��Sb����ɯu�tS��.aߎ�Ŕ^�2�()֤;�6�;T��8�A�����ep�����<��
���9~OL ��z
W����7£c����R�mp
�6���;�7�.�����D�S�w��u����Z�b58�q����_���~�01�{~qP�W*��艛�p<�}�K�%�F��)j�Y}{H��$
�m�`��u�u�^��9���K�g�ȃEw<�
��Y�3�N֬T��)5>w���}^V�+a#�j3�]̕ҭa��ґ-�Bܰ�<͆w=��szmc`Ϥ�ˆ|��҅���<�x�ط�92X�Ō�^[�o'T4�+����o��%>������Ƽ���r���l>���.�/�ʥ\ɑU�����Ǿ),0z��j��� �(I9��Tk|�3�Vͺ�f|��#�/_�]1>��Z�oÆ
W�`���O6�E�W�O�f����唐u=���<'9?=���Y9rE*�^�Z.u�"�X\uS������`�Z�;�q?-��z����+�'�_��]�d�wkѳJbɴ{R��\�*T���.j,�C��9�
�$f�t哘�G���8Wp�������{QC��o>J��Z=)���� :;�P�c{^�����y��e��w���7�eF]�1]ֽ e[�/V�ml>}�1!��+�8�X%^?I�⧹.#�IR��X� ������%9��hXQ0��V���oP�pX���o�\�>e��}}v��r��:v���+�p�j��o-�g��B	)��AL�����<�b߫�)��?6:e�ʄ�i̺ڏ����ޡ5`ޢ]�����Bs��z
�uj��+h�9A���g���>[
�<S�ez���7.��pS���ȿvK��8�Ǔ���P�W;n�gӳ(�5�@]Wg{R�Y7%�u�`0%�O(Po+�3�]SQr���
_��$�p}2[՚��e�������O�vLWS}�~H�F��d��I�!�ZW�q��ڽ��p��Zt��J�͉�ts��d�e��fG���ދ�"�gA��Ai�~��+h���-~��F;�fR�]rb��{�c��Ɯ�'�-�]�tڞu�s�(8�P|՝-�J�h/�S޿]ǉ'V`��IY�y�$�G��,Z��ڤ���z��q��hg���h�1\^8p�W�-~鄫LƉ����ȋ}�r��dXkכ>�i�;|��by����,V��ݖ�h���i-�0uC��G���8f��;D_�m{<�+	����囆\�ZNSr�(��wI����qr�u����c��%RX�zE��6��x�A{}�;���4Ƀ�C-7Y��c�Q��W�x�ǉ�;���� ��wH��.3ݝ�h�蕚S����Hs���>;h�J+����,wo.`N�0N���G}V�;�E^D3�A�j��3���>6�-�|�#Q��ݼ�G����}ΰh�:ʿ^F�1<��y+�P��T������sM�������!�������gU{$��᥵�L�}r���a���0=��gc�����"/��x.���M�8S�wL�&���\���(C��0&����s��E��[j)\Rn�WRg)�ڋg�K�uw�0oT�`�p��X���A����0���0���u��Iq9Y�:P�o|�P�ꦭ%ަw5�.�{3as�q`��s�]�a6.���Y@���+9��(��+��I��$G5w.��w�^�f{@��a�7�Y�f�M�uw�G��$��w��:�7<�gb�o�)4l�8��u/�M����*�	�uY���㏸������y��9����t�I�uP�YA2*��dzel�w����������޼�}�*W��N��S�,�ʘ�`��۠_�R-%~����Ε;��SN*ϧx{��a���:�%�a��Ζ���b�9i�aH�Aq�8�:^D°V��I�ǖs�:w6�z�AsK��R����;����Ͳ��=u>]�i�9���.��%���JlWS��=��ʾMm�\J�,\����o.}F�'+6���Z�^#ܦ�w���z"���2��*bV>kn�erNvo����W>�:��9����������@f���w�U�NHi�8%}r�ȇn׫������m���rx-���hn��g��\��>�X*O�:R.�'�P�3�z�a/=���*fp�����^9&f+�\8���ţ���L=߲�^�X����~�)�w���6�x���#zkC�ՏJ�!���+��f��]�<��W��ܥP����K��;�(l��d^J:_ޛ�G���^j��i��H�ьwq㜻a�R]�r0ux�G=��GTF����^��,p��FܥB]iCݏ#̦1º��e'{�#����11����K/���Nf���3��}^*�7��'�e꾄䓦q&�qO�K@��`���,oS-z�3�����9���7�+�T��^M��^�ܛ��z�w���,h�,ύ|.i��o��T/ή�����rK�c����yZ�VƧ$���r:)�Ż����b�����L삅"�s)չ��)X8�t��cdg�E��ǽep���^u���¦C�n	�T�4z�l�K��YG*m�\6�S��urkd�ZT�]�Y�K�����ZBh�ۜ�s`r������ў��`�3�qJ"1�Yj#q�oFysB����!B;�;�Ψ�2�5�C�lvOfSE�X��3�`�����䷷;Ўv.dO�vݑք	צ֞,��o=�/�׵z �_ө�{2����K^,]zvJ*�߶c�غi�Z�z=f��%,e24��oW{�w�3�\֟fg�NИ�OX@��=xv���ҟz?Zr��%)w��b�Kf`cj�������!Z���,����]]vzpwт��^���o�л�Y��.��:Үӕx��8]f��c>�[p�MAM9�|�TV�=Vo%�ם�pu�:0c�$\���[G�y��<5�s%u�>O~���J�w��]�!�*��־^�
|���ps�����x�|%r���H�p�f�\<�L�;8p^�b���G��ή����������r��%���;.��kJ����/����7�;��ʑz���*�̩����q�2Ǻa+]BH�e��7�=5���l��#U�G|*Ð�=>Vmɽ�+�׺ -�H�ǘ��u�����>�~î���*�*��OQ�Yd:�'����\����}J���.:겮�؀�Бb��E����,$c�Vgc�>Ϝم�3ko��UI|�f�9��<�����{���ۇ�qX�|X�G�e�c�����f����5T���
{�:�6��������0�Vͣ��*X�ȫ�����y]o�q=Z%����*���%�K���dzw��Z�_��i��G��Q���(S��9_Q�p2@�~'ܯ!���p����}�y�.����>{�!�β�J��V�i%�{�Mꄝ�*�����0Tt)N�U̖�x��+��2u	��~^�3���?>�=(���"^��W��$y��َn�spw!�7�I{I�W���0�v��(Nt0z
�ul~V��>	D�+v�L��t�o��u�s=��
T�Ϯ��s��b����]��ﳍ�'rv��=}���\5�h�s3���O'���Jyv
9�u&W)������/��Nyg�oVU�e�����ss{���7�	>3��ɱґ'�}� �v��\�k�#yx_q����ydN*מ~y뵏d��֠n�f��p�E�8΃b5��Z���d��"��U������=���{Dp��c�=[���>�NҲW\H\�NRț��0�Eu�@��gjwKj�/-��x7�BR5{�p��%��u9ʛB��x�d�!s����]Q�%L�=Y��rD�;�Oc���2�I�݋����Qo!<4�'[\K�XN˕�8�;��՞\i�WcNIF׆|��%�rV�%c�#ڰ
��U�3�O]s�n��J�C�p��Ήz��Xpo��.0��+�I^O�(��uK�i��KQ�m[����y�cރs��Ἢ�Z�P��-fʢ��xJ���n
d��9�m୚l`��Y+9׫��l���I�s�P�ឡ�f��0uC��G���8�����@��ϛ�)o�v�.���Yg�q�iϵ��~)��Ln�O��=R�:����5��<�5V��:�Ɣ����u�C�-:���aϫP�R%� �>�^�{��4��궲s����.���J\��r��b���jm4�dwr�z4z���Cc��u9��5�
�z�=������F:��M��\fW;��-�h�8���&�������"�e-�$����5��^��ٮ�t��V&���u"Y����~j���Ouo�}췻M
�E�+*zPڹ�mmw+����|����}CC��������	���0��9���=O:����㱢=�����'��j�{��2K���ifcW�f�H|��W���H�k:1�(�c�Tlʰ�OO�X���=J��7�Y�s0�8
��hڌ�&�wq�a�AX�m��-��	*�]h�z�9��d�iǏU*��Bn�	Z;Ga�0Z!IC��{���ɷ���μ[ɗ��N4@�]?�:�el�:K��t���9ۘ�l�,
���͙8_*t8��Q9��TOQ���9ct,PعO6��q�����tj�&�s��5ϳ�T��^�	(fڂ�-��J����c%�&��]��z�]��PF�})a�6Y�ܯN���buS]�[V����WG.��P@��y�\��4a!�!�w�CgB�;oTۭ�BK�Nȳ�u�����V�wndrC�Ʀ��5;�]��w܌����Ӗ#y��7g`��1���E�r��'��I2��S�����&�|��{(*̗����ق&���]��6��B�4y��Ea̭;�b�D��dJ
<�z���ս	]7�}P��$z,��ރn���,Q�Ѳb��hW����r�{����G�"��v�7�pЦN{�g
0P	a�+b�f���z���7�@ڭ��ȭ�WW������OPX%ܿ��/QZ.�g|�s�G�UKA<$r�X|1�����CI�R�({�7�;lZ7^�`r(p[ܝn�VU��Uk� �L�l�␰����;Z�r��Nstd)�N��h�D�Y+��;O=\�q	�K�� �a�U�aCgx�g��f)n��p�Gj�H�هL��V.���<=����9MW��'na��EeK˝
�é��Թ�cP��;Ň3���ؔ���/�,s�S�%ܲ^��|"��D{V��u;%��=���;XxTwtjVs��9E��w_r��1�o�s8
=̋��s��,�Hr�[�/�Nnܵy-r����<�[�]��_b���v��4��*e�HV��z��!�Gv��ynm�ٹfZ�,�F�-�a�G�2ec;��U�nG(�;f�Uh8tՎ�N�w0�p,�ʍ깹wNi�F�Q�y�v΀X�GZ i2�v.���q����)@:*�F�݌�XE���'Q���	_!ݗ���Kw��KE�v+��gTΜ;x�ر��a����
�Ҍ@��ƀ$��[���v+��rt���v;D�I�ն��f�}Euv��@�]��y",]�Ē־�ۼP�ps�k��S8&��I�m#,9.�;��r��諻7�;zJȣѝ�c4�N�1H��c[��-��v�ssv�
w��Op�еY)t���t	Qd��6u<T[�e�-�����u�a�1���,R�U�ئ��ݢ�>��3:�U���b�3��v`�u�X�9���"/3'iξ�AFw�*Lr�v�L]�Ȭ _L��z5�p���(i�/����]0+Z�8es�ܸ�2�����5cِ�bt�P��	C�>�Z�w9w^��[�?=諟W�UY���)iQd��"+mDDb�im(2�
�l>J��E�V,b#���P���ʈ��TT"��`���,X��#DUVF"*�ł"1,XT�F+K[
-lU�,V�(��+X�1�,Xʖ*�!����`Ȃ
0Um�R�m��bֱjUdD*Q�b���UU"*
�DQ�"���U�Պ��iP�TDKj�EE��f��&��U���	YQE�*V�bE��
,X��J�"��Em���X����H",�Q��[j��$H�CkX��*���* ���1�DTEE8@��Ŗ�PFE`�-�EU���c	R�0��DERV,+�(0DA�cZዅE���q����
�*.1�p؊�����(��Y
 �\6�`���&�K��QE-��J�O��>�����c\վ�뜞:y��5��8]k93}�W=b�I��`���Ap�G8���X��<�$��^���ƪ�ϝ����VQ�`(k����i�T��������M�\\�;
��76�����ծy�4`���\5O�/�Hox0z�x�Bǲ��iєY��o��[^|<=��\�y��Y����0v,s��τ�ܤұU5�"��4ؼz�ܗ���=֟������u>�^>��V�lژ��jZ���Xnm�>�E�u+���7ٙ��t�kOӸg?>5�L��ӧ�Ou'�b+�|a����V>kn���{/�:v��a]b�t�ø���{���6�� �xf��3��C��Um�CO��(C��RYU)
�ӯ��^����Hu����h�N8���~�`�*󠥾�2��=W8���Offc�<��'՚��v<'ܑ���lDp�k~�ַ�|W�a警�����W�䞝��5�NI��:U���ʾ�}h?�Ќ={�Y���C����ę�S�p�Z�-��W�΁f��v��5�Ε�/�ŏg��4���rZ"��~��Fgc�\�U,��ǵ;�D	hX��L�ApE����Ӝ(�;(�u�@�ݨ�e�̸tV��B�"XϷX�Q�`Ɯ�Y+���K��-,l�+4zfz�N&Տxo��X{�o/�i�D5Nht��3��	�Þ����"�
�Hw��=�[����:���\��nM�G�
 ������f�h;��gU������FPcc�ܦ-�������V|����"~�"^�\�G��M�|*ʦ�r�����K>�[3)�ú#���lwW�T/����/wx��}��a�{Z��ߩzе�9]@W��sz�k��)����6�G&��p���ۯ߿V�[[���w��F	�g�U�S*Baߓ1*����,��1�e{7�f�সma��,�	��
��>P����9�'�|��)��1�Y��'w��+gTM�>Wj}�F+z�,�..k��,��M�����'H�e3�`��fCkr���y��[�Q�z}>��-:�kAfsy�u��u1v��Ԉw=�@�ܚ\Y���X�3-�ޯ/A��w ��SJ^W��;z�:�"�,:`�38�ͷ���S;����s�y���|�Ox֥b���L��^'���p��|�Ϳ�;>���w޽�8�?oQ��{�j�7 ��'��@��GAh���v�Ux	�p�f���5݋»�WK����9��:�-`Ǻ9u�,������
q!�W��O��7_󍠛�'��rxa���EK���اn;���ob��k�;����*b¦�e�}V�3{�t�_S[#s���d�ש�}�����5\o/z]�d��M�������t��b�6*�	�}*��:��ѿ�dv'T��R���+�Z��(���5�]<s4��w�I@�q	���Qk�Ih��Yju�Z���F�Z�L���9Ob�X}+�5��3��c<%n�I_��$��q[Z������̳��+T�:��.:<���2X��{�1�w��+�q�w��8=CL�K%c�I̾v�Ƕ�ю�i�g�U�i>/r��=�o:�h�"��d��YC�r5|~�m���"�/=���g��y�,�`��^V�kF��.U.s��ޥ��
�<�e�E�S~#b��/���x�lF�mv�q���b���v�RIl�h�j�¯t�f�(4�Y�G�g��}B�l����sQm���$��t��\:���:����g~M���cP���2��;���J7�X|I:<���׳+ϖ_w�V��a;���D��.>�kF.N�0�o�}3�(|f\��'��K�Q��������J��3T�4?|���K�H��ō���/%	Ά�+����5��\���oJЧSg�*�޸1�gs�!�n*�{�\Y��Af���O:+��)����3X�5�ܳuՖ̀ݹ��t��5Rrs+Nn��dģ���/��]]�R|�1�㡔�1vyU�y��j|��L}�JvU�\�٦�"u��7�ú:i����(.�ӟ:����v'�:��`�5�eLjy^�9���������G�[���b>^ܽ�ϭ]�ٔ�Y���B�;��L�uMY�r���
_����������D���-��9��=���i&��d�:D�3�!��A�u���p���ԝ����[���2g���G�Ѫ� �Sdˆ�K�p�Z�4:R�]%µ+�O]��W�
׎F.�����.����ޕ��`z"�pIF׆ ���}+n���^��qQ�=�{�(�Nǚ͹�;��[�9�8�]%�_Ev��)�lIKU�5����ˈ�I�{kǇ����6��Z�~KEc.�
c�ܿ4�ހ�LƉ�2M�#�Wa�Sټ)�''{Bw6bM�����;Cڮ�3�۸t�z�5�Vڜ�ҽ�
6�#~`�⸣/�ˆx�{{�h��h�ϔ,�Y��a�Nj��O�]'<i��넫8��cb��Ko���1����l�n���\����\�-�����2��['>�^�S�2<�Y����� ����J��w�3.Xt��>�3��3��RZN�S(���Ƚ"�F�cX�}��iy�rt���"���ΑY����O;�n\Rt�K���YMb��oX7|5�|����DS�V�֮��r̳�ܝA�"��_r���l�S2���M4;À>���''�����T��q[ �c�l�	w�k/��Em��g��w#��{n��������q?-�/�;��(�+i�P�ޮ�G���y\�=q�ڮT�U���#�H�.i��7�?P�8��P����p{3����u�@����!�wJ����c]C=�za2��0�s���u�4�������:�m�O��љ*�0�+�'�|#��r�vS�KZfo��^��-��KeS�vvt�r^�=h?)����G�ج�h����.��R�VUoY0�����T�����L�nK�ָ9�l���r�J�����A2�y㠽y��7ᑴ�v�/-�X�`����7�zס�'��3����粁���ZY��X�])�ڶ'a�6���w�5].K����O*�Wp�B�Z�reB/�X,Ks;4j���6|�񊪎o���iZ���ڨ{�mg�84O�^�>����4o��ᇤ˦���]�h���^�-ҳv�U�㯚��R�|��`̑g��U�R�R T����|�\�
S��V�Z����\�Q�X��{��sp��W̉ҟQLݥ7`ה�V����vs�QW|O<�*�{���tT��_"6����[P/V6�`���u�im�=�\<:�?	W�Iyґw��(v2�PA�p���Gk��}�l�Wu,�g�̌t}�H�^�ji���WL�'��_0�}���hr��:gC�H�P�5̀�e�^���κ"bc�ч᷉3��3w��.J�پ���}�K<v�Z���#z
ߦ4�z�%�n��C�i�٣H�(/W�{S�>�;׈)ޜ�q�����X;�J��L��?Te69���m{�E��}�.�0���i͌��<W��\��>��H�Wn+�:��w�ĝ�ٙ�3�A��{��3{g�1���*�:��t�w���g�����V�eA���t*�ˀ�ަZ�g}N�(M�a{���y9�r�t������T>��F�g|*�je*E�b�bZ1sMLO|u��]�)�pWs��t��L���k}}������GH`�o�Ih�i
׃/���Q�-���O�~SV�1s��d8���x��M��=�M`N�b�)�����S~����B�M������'�o����;ɦ���L��m�k���z�;-n�3r�s���*>���8s�;DN�����k�]�3k[J�0q��1;�՝��
PL���F��	�v-N�
 <FEs�<\)m�8�V����u�#�1s�����Ɖ�9!�ֳCNt^<<������j�9�KV'R!��ٔ/k>>[U����Z���[;:�t�- ��b
i�-x�7Ѓ�~��pV�W���W����R��+{e�n59��B���
��r��<��K�����9������~<�l�+�����i�Aيƙ�~���G�cѓop�p��C�.*�)�ׂ�>V7ƙߏ�1�{e폛TR�x5�T��<�D�A�r�Y�a�e]م�����f�G�y�8n\u��=v���	x��3n۽I�ou�K�2w|Qk�Ih���e�p:ۭSz�C=k_�\=�C�7�^ؽ��9
���b�,��h�j��,O4����^̎p�='��K/&�y�_�__��Q���AV�(tw��9�e���]�Hr��^���N]����f����z�Nו�gx_Ǖ��ЫG�2�1ՍA�G|X���"7�zB�us/�ֶ���/��ǳ��tt炵u~,r��Ⱦ�`��|[�^�S�`�{y�;�mb�%7�.�_��񣉜�ʹ�2Rɪ^�W���\�ĵ����k�1��c���:�6�D��y���[��j�Q�r��	��혬B*���n�w��U����j�Y�����t�-����D�U�h-����N�S���:j|���/v���j�¯t�f^�_�c>�xa.z�*z��U��_��t�mo�R��w-R�+��̇~]/�������O�ܱ;Qg'�X|g�-��$�$i[�ϕ��� z/����V�B`.[��AL��a�*PMD�.Օ*��H�qw�h�2�N"��n켪�#z�=X�%�{;E��':�v��G�a��3�<�Hi���K<�y!�>I���O��\^�i��M=�tO˶��L��?q���Y����a���̆�Ҁ?m�x;�(f��O�`�C�WRgº��N\>~R�~�oOu���ךX�/m:K/��x���n|�I0؞�d�:D�!�u�A��hU�VY�v�~E��מlT�2�^�����@���f�������GGJ\���GR��6�ݽ5�{W��s8����9z8�J��Γ�a��ӒQ��9br�%�pJۤ�${���;��\�z�Axc��dT����ʋՇ7��+�.����䥪���3v=Hh���{]�5w�O]%馁T]^��KJ��,�e��.���]�V��#e���\��z�{����z<9B�^kۿ"M����u��3!RS������D�_Z�s2�w���@�;�Z��@�4_<KG >=O&q��ˢtC��M�� ߝ��d��n�+�W���2Ռ�tU�s�U��h�
d�>u<ߨ��^�5,�1��K�F�H���+ʫ�"U�δ�=f�yG����9�/#�(+Ϯ�6]�P����I�{ضA~��A�N�u�Ś�59�k`���iyVi��k����Գ�pӽ�����:�T�w�7Ti��o���~��w+ΰhu�Z�Ll<�/%�%qC°�+�ꚙgS�j���X۱�`���ڜM+#�{�����+t��0f��l��r�^>�3����e�y�����O�� U����p=.[�؃��l�|{^nx�}K]7�~d�~��:FZ������b`辧9���,.i��Q���=ՂS�q{�{��ɷ�v�6�ٕ�"�������C�E�����V5�3��˛c��l�US6s�Y{��ɳcg�]�R?]�J��6��a.!�H�j�P�|��������UH�xp{l)��"t���,���
g��7㏱Y6���;�A.�]H>��ʪ��E�!q�*.iΌ�ճw`�B����镝X�#��C�u6M�B���^��`dd�km��=:sA��cG�3Y7���* 㙼gq;fWs�e���W��Y:�m��
�d�\D����|��I�:�����`�>����V�����θF���ذ9�l���@�r�I(y���]L��&���W�_����u<s~]P�ux
u���>��S�,��*b��]޶�c�[Yh�mG��o���rP�O�,)/uʾk	��gf����`j\>0�^Z�vV��y�}�8��x�cەI9��.3p]��6�Y���<�j�>a���:�3\A���^�[[�Y�h��<}c��pZ�����.��>r���o����})�{��t"x�8�w��#�!��<���⣤|e�0���<���y\-q��d̈́�ѯ\Qk�{R��9o4�����,Sr�=�XY�����F�3�%V�?�᷉o�4|���ᦣ���������P�t,=��{�Ux;w����4��^T�ľ�b�7�N�Ԑ�X���w�h�����^��GvG�?\e�/�N-�^W��.���`ys�<�Xgw�Z���Y��5g����H�_����a�:�5�}ո�\\�/��F�V�bca	k&~��F�7DWX�s�Wc��ڭ�M5O�@ԭغ�|z��}�c7�E�m���P����oCZ�i�s�Wo;FP��P���D^�}T�A0[��e���_S�⹿�"����F���JU�PǛ٭�on��(��]EE�<ts��49݄��:�v�ܖZ��9Zk-$#V��Ǖ�rU��#b�`�H�΃v6P$�R���6�feb�2��z� �n��1�(	!�q���A��kƩ�;�4��K�wn[ձ�����5�#	3��9X�J���o���֎�H7��F��s:���J:�3Nl��b	Γh�['��wi��$Ih�vh�p���k�j�B���W�\���6bU�8��[�w�ʊ���R��_�VTTu����T�ýB��{����|�r��Um��}}��_Sz�����]��W�ai5�E���5�J�S|&��y��?
8�7���������v��콅�V9e�a�Y�La��MԧW�*�ޅ���w��ȝ,�ZX�yj=�b�TBV"C�,�8MK�\��$2��7L��l�q��������s*����X�B��Zv�����t�R
ۆρݱ�<�R�UXWx�J�Fu�|���Q����3�
����PI�m��v���bt4A��`��>�ڢ���x����Y���hv-mLӑ3\gQ��3i�j�]>��B��u���f.��V�|����̜��;s�5X؞/VG͘��dJ�m�\ιP�a���k�ŷ5���Y�6�}K:)㕷ա|��A�Ӈ�	%�Q�Z��ʴKu�1'p9:^ �_3cKx=�z�l�]����8m����o<�/�#֌��&��V�l�m�.�.�\��1��U��־8p��	�|��	�|+]3Z�;�ʰU�FIi�|�R�l�N�ul�Jñ�[)��#���U��U�t۫l���:|v
�{{;w���5>ś�u������so&x���_ E�y�Э�ymy_Z`]�f?��!P�T�n�R�^Vl��f��Vt8Ìk��VG%��A�����!��e)����J�ﶰn���B>GyˑBC��2�\������!���%4U_8�� ��>��
i���q��wAqވn:�<���h�1��F���jt�R���X�q�1&���u[�����
x_:�W $*S�޹+�*|�owP	s�/��L�ۂ���2A�HJ� �j�N�]�恹�p��k3:bY�Л^\�-�ݥC+�S:��X��o��Q�Cw��
!{�[��'xۍQ�m�6)����d�yq��y�%���n���k c�=f��m�:S��>������֔D�?2C��7���0�͸�mjd�5��}βV�����8�# ­��9Y�"S�t�flX�(�b:�Yb�m��p�[U����T<<�<)�����Z	X�V�EU+U#�QV�����5��aZZPŅV5��Ee�1!�Uja
��"���DA�U\1kE,0�L6Т-�p�R�a� �Ä�-\b��%Ha�ءL$�3BԲ�����J±����"�
2�`-lE���U�I0�QEP�*E�qh�Q�*"��J��,j,����0�)"�R�#��#`�J�R�j�X6�%��Q-��ѴQX�Ř�[IX* �,�H�F8� ��UX�%`Q
�qjL�kYX��\Y���$*�k%H�D�k!Y��lX�D0�Um�QB)+m���8�Y�hVa&" .Z�H��Y
���T�c+!R�Z�?P| r���w|��gaR<���x{{^椱(���X�*�n���k���x=��q9����Ԡ�__>)Q�ӃQy8]�����9�f~>ʌ׻ּ�u�5����)6����辝N��/��u��*�I���y^�SЇlϗ��89��'�\/�g�L�[JwԨq	��1*�E��J��.����^��t�a�d�������g�/�UGH�-�݄H*q�o���x�GH���*��V3����d8���+��,���̦����>�?�a��-U��ɦL�;�RfX�v^
�؅��րY����u�^j��3ԭ�3���=8y0���x�+�A3<2����a��;z��S��J洉qߎѹ+�իg�i�Xʓ��tR4)����]g҃0D����/�4�������;z�R@o��F�kM��7�q�Y�ʇ�/p�p�
���#cU�n���8B�V�y�ò�\=rk�2'�V4���*>0����!�Z���=��3�u��b�Qz�kg�Zk�{�T���I��<v�o�
JۨD�L9E�$�|a�P�ܭ��
b��CNϱ�S��g�A\�6�t8׊��T���E���Z+=r�F7�Q�l3cΉd|.�m��ywx$B���}an���<�$�av+�h����53�#*�^�{���v���ɲ8 /��5Z`\t]ܮxú=�QK\;k��u�1��ݶ随��opo��j�e��{�$��8,)(0\\u&t���Ȝ�l����
 ��ĳ�v<��{�@`~RR���t^�~3�5c��t�U�5�$���2ߊ��Dނ~l�2�yOl�Tgư�S��6�WPLm�f���;JJ��R�M��g����vm^��c��V����v�v��Po,7�����j��!|���X_��
d�~��s��v�q�����r�8䮷��Am3`dw��������;y]:A~89�'���7uF���{��x�K�8��+�#�\��=+�3�����*��bV�,�J��@�&qҺW���Z��vq��5 �dпWl}��e`�P�:��\�徂��[>)�����*��}N�^k���&��|���Ehx.Xv2�H�A�Ɖm���΃�`��R�wP·�`����t��ے;^�d���8Y���<�`���p�*��κ�h`{<d�z܏�g�����x�Y�X��G�};2�#����.�u�������]�[���	� �����*�ms/����!�nZ农�_Z�iyG�g�
�i*u�*-��q�C�:�u����N��瑻Q�����{dD�rg���I	>��W���ݢ���8�#�����=����j��J.�]�֛d���̵֭җ���]q�����|Kz�D��a���VM�I��۪4��S��i9�����u�"���gy��/��D/�Z�L���㯸�P�����5������옍�;+2��t_���Pt6(Zkj�_�h�����"�����
fJۤ��5�Ky
��R�^���zD8�R%���Y�/*/V�R��(ay����7��������Y⟴m�θ��5'�~Ӎ�u�ז�'� ��2�_nX�<h__�]����E5:���,�/#��0wQ;}�x:mV!81OU����n��c��Z�����[��h]Wko�_-�(����?%#N��5�g�f�޼��٧´����dc0�Z��j\�Y���r��t�� �/=�m[��v/W&v��2��s)xP����8sV��_x��g1U�/�6�Ca��.&��#�{�ͯ>�ê�*�VAo62䦹��w�h�O*}�b��H�mx�M����:�ܮ�!���>�X1�O<�"��9�����	�C����.�w�;ڥ���4��؂�i��$^��I��ہ����\�s�짾g��#]~�ğM|�X�x���Pp�F%�3�t���j�V.g����wQ��ǝz!#.�$����u·���G�r����	�}h|�������(���jq�p����E���K��A�V�!oG���:�oj a��g��i���6E�Ԩl�.�>7�Q+�P�,�����
�멕#γ���g���ΏASη��a�c�)����5���Q��y�y��C�q{�w\���̝0�lMwFD=ˀ�S=��q8b�9I��/E
���㙯�"'���O����qe��mO��{���M�e�}w�0v,�oY�;�{����9�Њ�x��e9�H2<~9�

|P�����;=^��3>O�o��-=r�ۘ,?mH�<q�˽��:�d'ِ?�F=y����5=մ��cR��R�.�cݽ$��<�$�ۼ��LJ^�M<ഖJ�/�=mx��[�wF5f��$=�I��۫w�t�,S�u���\=\��O(�-��)��c�x��~c�{�N���9`q��r�z���t�>pS��#�
b� �!0ri�5��=~�f��:��Bv�Ǖ�͏�+s�?M��^Y��[�b�l� &L��Z�e};b"�e��k��-���D���*�i�H�\�}zk�BcvWJ rFbt�O�\��kޕ}�+�(M��hu� ��0@S/�L|�������7�ս�v�ф����%ݪ5�B����7ނ�XndXY���x���ۢ%�fo�G����0�鷘z��E�H��N���Xρ�<��_�er]%z.Kb��齔5�pS/��9nO3�b��S�0��gz���w�4Ϋ��ݻt�=�X���l[U��z�p/ N�N�}�f��X�t~C¡K�rbch^x�:d�a�wy<rU���y�r���Xm$��W��C�&��3ʯW
^�-:���/oU�%�'E�me���m�nu������q7c�OW1��}�=���g��W�DP�7�b���M�w�W����<vO%�q5 ��Y�\ꄹL��}���e��p��\���<����W`5�T��;�/�Z��4�y���"�c:�.��g�����+��>نǜ���=����|=�/9��5�|�
P��v^U�,']6��<�]9]��Y��d��#�l������RDA޻�ly4���qyB��2���W��\����LbW5�����u�X:|����k�uh��K��SS֒��Ѫ���M�i��d��mgF����`]��◾۩o+�z8�XW)>}ZrƩ�� �xsT�7�[ڒ��k)�m8qpwV�.�2��*]u��������:6+5���G�S��$�l�l��|A��P�o�{B�F#�	A�z�F>��r�#����b�㯘�\�������b��0{���v��/p�s�5+�.*����v�p��\:������Q�klb���rZ���'��"DWo�dg���<'+,�8VBG�QV:�i�}F��^W|:M���`�mru���`����IT���Qk����E��k*���9��ո\�}�t/����YVi��2KIX�±%���K��yc��|�|��7��4��o^��kJ�����N���֩k�j���i���a*��&�z��^���ȇ����2����>�\ly�`�s�^Vp0���R��S_ZQ��Y��3�~�{��x�gޘ�m��B,�{M�^�;�������Jr��%R�/��&�P��OR����3�6���h�/�]N֟|\L�Gr�-�V��<v��(Ǎfz�uHe�9kw<n�z��uzG���S�s����o�A�B��۟u�i��V�J�>܍Ĳ�v�H\����t�K8WQ<fG�+0<7�O)�Zd:�E��ŕjи��ɽݬtY���Y����+$��K*��')0F9]��#�I�o�8\���%״:��橒�M�ɽ�rcּ= 6ܬp�/��/#��JJ�h�ٚ]��^H���O���:q�9^��U�q~������&���Vu�:��\��N4Ϛء�K,�>�b��<�ʎW �O��{Rj��*��\��eF��t��oghȄ�C�3�87��;w��Պ}�#��!$����R��.��TL�e23�%�['nL�W{�m�nK:����ϯ�f�-�����xG_"�J��5>��QHe��iq���^���o�v/��Nyg&Kz�eq�u�Csڬ��~gݡ
�]���-���7ö3(�����y�:ڗ��"�E-{&L�K�pÉ�K��"���;��c���ER��Y�ş-��8�J�{08j�(?)/E�G�U4�j��I{z��O�ǖ�D��6t��E�Ào�E�_��9%"<	/SMm��bǛ�4���{$�owkܖ�t�a�?��M�:}$��@��}(���VEny×=�a��s�M�������Bk�X�L調��N�EI��8��],�Ƽ׺a
 9��ϒ��$�ŻX�~�-%�ø�.`ď-��H�-q���4�>T�/xQ/��\�T��1����w	sv�oD�Du��ݷ-�zV�S)�J��a�wSOnm;5�|�n���p��#�$#��GyZ���#M�)��Ѳ�z�lO7������6_�Q�:y{r9�%����!���k��5kM&ѳK��,�A�҄�cZƠ>6�-��g���CO��W��\���S-<.�δg�,�.�з��L�X׌�����c}�q4�#�{��{���Zs�������8��Xx[>Z�9�z��%� Z\_�uX��/��q?!c�J㲝Ir��^TϞVT�s�g�e�1�-v
��p:/�D0u"X=.\�s[o��m��[���t9�ިa��]"�CA�7�Dr�U_�}C��K��v���ͭ����	��k��x���ß);�
oS��JҌ6����\ �y�����^zy�*�/���V0:��|ӆ��J��)0~�A㏱X��#@�>&��d�ޓ;�U�0X�P$Bmz#�ܦ�����,��:��r�Z��rv]���ߡ�%zvz̕��@����	�Wƃ���ڵ�;}K�_�f�&��,�ʳ�pn��5�폱�ᇤ䐣�4�Ǆ��S�=DIb�������[��3q����+8���,� ��K���լ�W���M�n�-ޮ��ߟe��lB��M��v�UК
RtRb����S%�NRSWO�۷h7J���;Q3q\�nN[a�������o��9W8�����/���p�2�q�j���g�|�3��$�Rv��s��m_M�Bit1�K=�O8-%��h��k�X�@��:�%�1FUe^ay�M1�k���Uj�w���>�TD:�Q�~!t�����us�$�k��vW�/$��ێ��淂����2����o�<��k��Cm4k%���s{2�׾ٱ\���ԏ���z+~o�W{�zܸ������v���C�A��r�u�w;ς>WZwem�
�v��W�@p:����|��``zի�bٖ��i��v��	�.`KC�ۍ�5NTyX�kFT��g�p{�����ݑ��Bwj��5%If�X��sz}��L�3N	Y�z����F*q�=Vx�T�/��Bͦ&�WVC��Udo����,?!���ᒇ{>��<pM�y増�N���V�`�?a�.��f*}�z��6u@�3�a��c9���ʇ��=���3L�W�x��uhz�w���L_�-dɄ��r�P=��u:ؗpsޢ��+2��y�&��j������ *�������ât��=ύʙ�������	�uãr�Zyu�Ί�Rܓ���.�uo�(��B�
���{;�d�r�z��:�P7����է(��vF�:�|-lM`��a��T9�r�͂��g�c,�j���\�	��t����C�ԙVs���H��T����[�G�l�^���?l�C��y,<7�A�:�bձ��������T=�3/�we�P�@��+Ő�<�h���Y��=iT�:����Kޞ�;e�(��<��
����W��gb���m��B�c��m���Yc��<��9��XЄ��\��[g'ʖ�8�O���!W�u�V�~�Ԏ�ה�����z)z{>��-;7�>yP�;�p�B^��61?����nǕbB�k�N&��җ+��/��β �Ev��AVx`�C�^`��V��G� ��,oiz2g��f��hJ{�f�R�7�%m�"�`�r�\0{̌�c>�l
椣���97�$���E�ϭn�B�f{4�ڶ({�$�y�a\�.&u/
�_�IE�`�1��f��Q�eȄ�`����G��O�eV���Gz�,��i��d����c���7�52W{ݩ�>U�ďK����u����w�Y��:�ھ�"<����v�멏;N.��:�Ѐ2��	�i�^�ϛ����AP�nY¯u�}�Fmm�;��ڝ@�<E[���t5z�o�u�p��F��J
6�
�:���+Z�{}����) 5�zN@�ۖ�|�ɝ���e]����꒱S����]i	������5V�Dvش�h15��3�X�]d�Z*�
43��Ag.��5�(i
��ۑ�Ļv�d�{�z�VZV6o$p�O$n��&����2��ڟ	Ɔ����X�!jgjٮ�p`�Mm>�T.��ܾ���_f����-/f�LƢЧ��B�(�e�=���LR �5�yrp6��o�'�P:�B��C�IK��G;b^��-�*K��[��� ����L&*�6�+���և$��rܛko��'�B9��[�s[��i��
^wE��Z����̐���`�!N�tr�=y��M1�.�60�q�����
�\`�0ި� *^E���)H��}��Ӹ�����e��M�T#�-%H�� w,�����LI:��`�B�4wwN��Ց��]3jh>T����{n��EKRu�w������P|.�dR�,D!C���Pɑ�$�����̛�����\��ګ6�n
�v�̮S ��d_]�3Ҵf�j�g8VwL��M�PQ���I��Co��Ȩɫ��,mꡨ�v�m�ט�dS޴��`���J���.��y����)��Y��� `��K3j��\k�U�H�&E*�!�wqj��p#j�u,�0�5ӄ�7��&�i,�u܂����ӫz������w^�X��g��)��;��X��`���>�l:9t(��+�ś@�Ů�.�dq��ҷi���Qr�c+��5�<��EDm��h�i)�Y��fd[I��[y����fm��Z���ZҼv�@�cIЖ�>=�ںk���b���w<����7;�p,���K�:��;��q"�Մ���ʫz��>J�r��>��k��>U�y:�;�sw��/�p�]��l�Fϯ>��	rz�B1��K�.Z7�w���ʏ�"�5GN��)�N؍�������u�p��\��0I W�֜�(ݩ�-r��Rӊ��W�i��9#�t7y˅���9�aػ�Sz�CV�b�U�r����C2�ta=�S�hd\w��䜡#lVY���Ն��N��gF5R�.��8�r����X����ۗ�H3r-a�v4P��$+�� �|��]M���le;��;>.�m"6/�Ѐ��sr��j�d�9��#��x;�W��N��qn�4�Nbs��s�;�ybUSo�"��jK�>�֜x���MkeL*���oI��K6��B�],��6E�`"�dNr�w���Po@g_����}���;КoG�GH���+Q�VV"V)PYU�k	�Z�
�����,F��P�e1jS��6�J�p�Y\b���!�X#��ER�¤�L` ��jKim*�
 ������V,�VKj���E
�i-Z�F,Q�+"6�
��J���aZ�b�*V���b�J��Ь���-�b��ZQ(�j*1����Qeb���,)U��ieb�h�Q�أ[(�[J�F��FA���R�,b�T�m+j��ej����m���ё�6�$�)m��m�*�X�iE��`ձaJ�U��j4�+kT�Tb���U
��	T���N��\�='�m��Ê�W!����z��6f��{ǟ���gγz�WU�
����'c٦�|+[Ǽ��7�� W��0���zl�7�Q�]%����m6iI5Pv�~�x�>�$���G�Y읲+^�;���A�6zǼ�J�����l::�����!L��ݵ���-Q���ܿ���/�͌����O��:����6hǧ@J�t|���wI؁�mJ��_�p7���W�X�y����3���p��י�=�v{M1�c��כ}G�kZ�
�n,�R��d�k�ꄛ�Ų��u�:�ϋ���N4Ϛ���QZ��X�]�+��lQ�G�j^TyŰ.Xv2�H޺Vk�]��U�o@v������\�2�:�{�[�̤!���I���R��u-3��3{)���{E�=�m�C��1�d�G���9��bv��ٔ�u�N>}?B����,oK������g{�vw�@��3~�~?X��Yɒެ�\o��"��d�H���}ٴ�z�:�5t'�����x �	y�<������R�|dB�zJ��.\6z^�Z�?L�q��P��v�9a�Wy��c�h�%����s�6�(:��"�Yq����u�v�X�v�5����s��Sb��#�,h�z,�2=��Ƙ�Vَ������iY���v�?�q��wy�=>�*�ͯ%�+��(���.|��T�}��4َ�i����-���[�=��v4����g�X��
Z�me�Uf��3�{��@�]���lcP�h�o(��g�o�E`r��+�:.+�{�U��)ӿ_��)P�0f6�ZD��]G������p�ˇ��y�R��}�^�b����{�U�ku���#���7҉�m��:z�P��=V*S;�p�u�4���YX�I��;�^�g/y��$�|W��(��<f����Cf{��u��LL�~[� ey[���i��Ѐn݆pj���cbƠ>6�/���|6�ʬ`u�Xwב�a�w�V�O�r��2p㾫HcW������u�t�4�� ���؜�˖��9�6ͺa��gg>`��L�+dJZ�U9�z��%Z���kGE��N�o1=C��Z> 2Q�a��b�޸�z�(H���s�\[A=^�|����� �{l�y+{M׽'g����~���<�A�{-��Co�h��>o�`sW��
�B �R�<��ٸū��DL�cH>[i^�յ�]r!-���v�T{MҠ�n�N�E"�\�[J,��t���0���\��c0��3�%e6�.�g �N��ԏ������ݻ�L,	��|��9K��X����8�a�����rp}�6zg�K�3ɼ��~���,	,xÉ��w��*yֈ�a���o�Ƹ.!������M���e�����S���`j����s	�滣"� \}��<q�+��^�4�!Or�M�]��oLXl�f�ȶ$Aڿ_7o�3~;�mM��d�/y�s8UK��Z��Y@���s�)B5�S�Ƚ����3}+|�)hY����],O�����3_=�d�s�P.$ZJ/���\T&���}z�EY���V]C r9�6�c�k=�s��֘8T"�`�c}mO�ഖ�h�7��X88hY�n��x��ˇ������ޣ��=�U�2CO��BJ�"����+��^]�P�3�k�o�o��y����J�Ε�����w�EG��.�{�O�LVa��!3���oޗa��^C�a��Mu#9����h��x�T��V=�`��+�̀�e�^�>6�=+�,��G��WVI^�<ru^�W�V�yB�]�7��Pu�/�t,=��g�W�䧩��y���R�*h<a�գ{�K�a�)��b�)vHDsnI�v�P-`G������]�iU�J��8���P�fF�Rݪn[g&���&��,�ݽ�J�c\��:��z�n�_S�-O%�e:���Y\��j�y8:
��,�����.5�S$w'g\�Sy^>}�_��\r�S�r��X���i�=���z�,�dG=��dwd{��'����a�{���#��e	'kaW{����h�UC����p���<o�D�������z��Gݒ�r�pW<���=A�wW�P�d���Iu�5���J6kS\�T˫���^A���Y]/�p0��z�1:���s��;�y���.3L�/R��ٻlއ��U2/�t�>�(Pťg�r���:����s`���$�Y�S°�Y��,۱���ܲ�n�D��}�KGJi
֗h?xk75;~����.k��?y���bIz����㴘p7�M�c��z$�3���i�4']*���.��t����������g�ڣBZ��R#�OfP694���̼�j`��0�\����~�˯}��{Az��>��kM��y�4M�� 3B�����䶓��L��iC0�ŐN\E�V���{�[df/�z����U1i����/p�p�D��qJ�16������=���]�K�X��ݝ6F�&3۫Kx�n��u��EV��Ů�wV��jt,So2�G��j�:�!W�C'>�j\j\x8�����Y��Jc[}ɝ��'�:��+OT�Vv,)9�K<n�xZ��Z��N5��_N���p��PTNu��L8k�D����_:�dA��]�-�U�0�ļ�a��U��pub��^ɡf�b�>�l_5)�����'/ΑM��<�+�9E�$�|p��^����9�^�5&��=[t�����C�[��2�g�K߽^��i+�¿����[X��w��*�L�:^�L��@p=�r!���@e��}.*�U�C�l�~�`Y���K��1��7غ�T{|I�[�[.W齂��eyYϘI��Vm`� =�ɩ]^���#�TU�/��<�/��~���zǼ�{���ʲߔͭ���Y�3.��6���{}E�!���A�6&/���2��/.&���;�{mޟyhs���W�g�u��.��8����U�X�-O��hf���Ft�|�/�.��=�*����������N�>9�ȳ�+��\�S�OW����X5Ӌ��&�#�3�[�������Ot��������a���TdKyJ�̹d�*4��/}��~��</��`�5#���ݷk8����M[m������D�-��[�#;5V�W��\�k�Xf�`��5D#�t��6i�$���Oݐ�O���y>(���W(�������{9r�v����sx�l�ҠVr�a���9D䚈΂*g�S�Ƕ�1��M?X��e/P�y>����t���'!�6��jc��Q��¾"���5��_�k�GtE?g2]���6p����j��=:�,����
得ˮm;u���1ޭZS^�;���t�?\�yg�oT�[�'+x?d,�@ڪ�F�Ew��xw_�xgLn�B��8�<u�,	ˇ��_��	��ٕ1vhɐ��%�hV���mV؋ӼMӏ|�'q,J}U�VC>���z��3=ԞK��Ɯ��.���H/��ֵq��Yt��r{�_�m�V
��V�%`s�y+_��D��,X�Qx�}y�x���h7��Ƅ��{}��sd���`�H�|�yd��C^�Ja=J.>�]�(b�u��	���cJ�W�Z�x������k>L�D�pS$��D����	�5�ׯ�u����ym�X-��>iw���m$=��)t�q�^ꀣ�q�8f`v���{Ys�-�Ae�8\�W�mAy&k;�^r��]�t�(=�c�`���-��g��[,i��\Q���~������K�����i<y� `����w3=��~�����y�N-|��.�&�٘q���
Ⱥ�2q��R�A`�a� �����&Z�z�ps��K��ۡ��{e*��E�L��%�+��'>�4񃂭�y!�/#,G�諀�K���;s ���i{�k܅�.���ɍ���8+���c��0v��J������qߏ�E��>���<2r�3Uj)�X6〿/�����x ���Җ󕊟���M�F�H��g<��ԈF���y��v�`c;3�m�E�AquOW�'>�R$e�W)����+����+����}|A�v2���w:W�}췻M�q���IإC�.�<^��Ѿ�씽�<2c��J�^1`ׄ�(q�������[�~�f�iF�p$��+��+�j����N�5�ǴGR�\�uD����߽0�o�5�YϤ��z϶e�w����jz�A��O��O-���� �Y�w¥����<�9x�bo<�/����0<H=~u�z������/�*a<�ѧ��	�Q�,�/uĉ�|�?��ߍN��v~J��wK}�L\����B�y;S�ދv��G�u壢��ꊀ��a���Ն0����]k��kC��{�g�U���Z���P�VͺHt+�u+��p������hX��|��-'�@��ۿe��A���>��;��;�,,�B	/.����V\����UP���z�|��,ᗇ����IN:�L�բ7�ΰ��=�w��el�֛fw"2������J��n����c{v��goU���<�n(�����}��ua������!��pJ���vD-b4<��.��K'���j'R�ީt��M�3�/��".�͘)X�� �L
~G��
b�IZ�o?o�>��8����~づ�t]�[<9�I��߼�h_�,$���*�s 9|�<Gǻ���8��S�
�S�5�O���B�J�!�@��ę�<��G�6��
���XOe�Z�����W���-�ٍb>Ӄlօ�Ҳ��T�����k���c�q��e钯:sq�!��T�����2>�22�C�L�^W5�5��O����%]��VZ����ٔ/c�D�9�0��5��z���0;���%��0��긴��{��ʯT�3C�Y�Ƅ��~圞%�o,��;�FgV� �T-`��bu-C��ƗM\�\/���|c*��Ogm��Wp�%1]қ��PdJb�E�\�Y��&Ψp'-�h���I�§I�t���잂�u�LR�/eT7K���TG_�O���x�5�i���5����Nti#�2�3Z=�euG���t6mY�E/[7O)�zbX��	�z�x���=ydmN�;^���۞muE�ʜb�pz�c-q���;��P��8�k�r>z��5�`�ۣ��'�(޷̼���w>�%��kU��sZ�x�w��Մ�#�bc��)/�S=}UL����i�]2���K;ZMdwr�9䳾ޝ����ݖ�j�Aڿ�R#���-/����31:S�UqY��'3�W�|6r[�Z��gҼe�+��g>��iɔ�	�G�"��%`R~]�P�fy��m��Mcz��;  ����	��v���1i����{����D���.(���$�;�C�7��Cw2�,u���{����D5OW	Y�}r�	����c�U�y]8]W��%�än+��]Qg�7=��Qufo�
J�ug�ޫ���W��pq�5Rs۵S�9�aXhس'0�Lz��Ch��I����l�� k�m Կo��@�lZs�7�c�����Y�:^V��8ҵL��-r�\�\�ס�{���}O4��g]�y� ���=��z�����e�A���PP��EY)T�FמA��ሻ���|il�<��L���DO���#�=c�Z$�Κ�Q�L�)Ϲ�� ��wB�����̳}ScH���̧���i�FՋ����[�v��cS4+`=&XU֨Љ^�<R(�s��ܺ$(贗�kh���JV�wl[jZ��]aY��:3�����E���%
�U��W��qiC���uj�|�k��@�l+�vX�������A{��ஹ��@.&�����w��Z��E*"�W3�Z�����R$״�S�g�L�+
���ŭE�U��.wl�t���=|�^�[�)��ʋ���_��I�>�"�D�>'ǁʞ`*z� u��]8���na��q�{���r�$ʪ�9w8��-.9���S��%Xa�
U�e�%�ʍ#z�=Mj��y�~�T����'�|7+���>sDߊ�*W�;��|J�:EͼN��c����0��'ň�������\��oY2��g9���||�s���;2�Y �yJ:/�cy�c���N{����h���-B����r�~��~����92[՛����J0؞�d��ἶ��vק{ms��I���V3�c:�r���R�|dt3W	�1vnI��"���p�!�E������`�>�R�UB:�����+���37�������.�o+n���ӷ���+Z�êR��$Nq#	���H��r���������֪#����1��v�0]��sL�2��>VZ�v �1򽕰GCP���,�5:f�����U��}G���j�Nr]Ovs����s*��� ]�������rZϩ�Y47�!I�2.��V=�z��7��x}����v]�k�ؘ+�*X/���}�G$���ˤƜ������6QQ���ub�P���{�gJ�3�eZ�^Kha䣊+!��U�o0�w���}Ԩ�����<�u�n��V�#]��J�� pԦ���::�����|��+�y�k��G�l>5��[�gԨ��zݕs`'@�Z�0r�p�V;�,U����3�Zu[V�z&ݘ�d�>t���'p_.�ܕ�� a6��F�X�� �e�	C-㦦U�#tц6N�D��!/�3��`辮����zqߓu�9��wu��vWv�֫~8gf*˙pN�S�j��3�BB���jcf��Y�v�n��Q��nU��@�W�~����o1�VSyF��P��,X�U�p�0iR��Gn�%+�gZY�s����$E⭢4F(����"�9�t�V�΢f���0�[�� �W8a��fK�6b�ПL�,ش�'V�J��/��y|д����wʘ��o�����5�ѰӣxgwWZ�5��ԓ���a������{k9�@�y��7�:��w������ͣ�#a�5��ݷ�(�:r��6�fB����wG��ݡ�`�����BX㯓ц��r1�����r93�tJ���Xt@�����7�m��4$$Ҏ��Uw�)�x�&���f�e��i_��S����a�ާ�>�����[�ڋ�E��}-��)�|�\G�vs3{�����4���D� ����J��'�Z֪��o�1ɻ�E�~vɄ�����P����b�E:h�]���K��3�:y�"�
4��w3r�4������Pͥ�3$з����͢�.�:�K�<6>ܛ{�(��iͱ&����uk��n�R:$���+�n3N*�i=%X�Y�L����c5�.JU�wQ���rV�֛٦ȣ�&�$�ӏ�d�()x;V����S��t����Ѽ�����oR���$}�^nX�2�}�6�_RF�G����Á&p�qu�8 �-U�9)F�=f��Y�ӭ�+y�5tn��7z����	G2cɼ�X�MkxU�s ҈$s��{�ȵ�Ob$r�����DuT[�����.�--�q���x�Co�fV���ⶦ0�,�=���2������#e��ǥ��ƥ:H�U��4�/���on�m��T��׆��ʮ�4�$)G���U\��������iV�b�;��2�N�Sgc�ft��d�*�ǋZw	��Ae�����uĂ��������t����7oc�^l���N�2��]�Z !+��vH����8ڌ(��=v!�7����mke*����j�0Vص�m���J�U�k*���T+e�kF�+V���Q�k�-
��j�ڈ�[R��փh�R��ȱj���У[l�Җ����6�jըZR�QZ�j���(�[h6�����j�m��Ĵ
�-(Um�
*+R������Z�V��V�$[ej%���X�QRʂJ�J��[l�ŋVV�����TD���ڈ-����DP�m
�V���E�TQ*�m�Z�H�ڡU
ʅKZ�F-�b�Qd���dPZ����j�
�TE��ѰTPkUiiJ�Y*�*��5
1U�DT[j$�Z���m*��"�J���Т��Uk#h�,X���(��VU��(���Q6�I��cDM��g�r�<�}��c��5V��.��YJ!�u3鬽]`�w��z� v��Y����v�A�����Z���WSqu�f��� n����0Mz�(q��X�\}x�"�^�`Fڐ��6��T�Y/���O���V=�!�4K�q%�҉�m���^��&�)꺔��㳷�k[ES��G�o��˶�Ί�=_ �L���u�Q�5Ǆ�3�Q�##�Hg�ۯ#���y8���)���޳�ч�D��j�����5m�0oX�\`:}������yl��Ǟ_=g]�&�4J�z��(��ٖm����T>��Cc=w�^!��m�Ʊ����4��?xW��"ǽ��	��]x�A�V�E3c��u<�ӓ�� ]��`������þ�*�����72@���c}�v�]�[��`Z<~��V&�T��(E��z/u_�ګ~*WK��R�9p��I�&�]G���t�0�ԧn�EF8V���J^���ә��whҹ+ިb�d�(x����ނ��o���U�l.5��5{�i�����-�L�"�#�@/��'\���3�����fD=��3�鸆�g��y��ʦ�ց������t-���3s��"���w@����s��,��͝��)ߜ�.U��� d(y��"a탒Aw����_A�l�5-��Φ4���"t�Qozݽ��qJ��6gg^�XA�NI�j��h3�z�yw)9��S�0�`b�����Bǯe���+�#t�Xy��͖<�`�	����}�8bSޣ�5��/��g�Z���g�Ě>C�eȧ�W3Y�N�����,�?��w���ٛh���/!��B+l�od ��mz}^܊��"8������K�]E@rk	��5��j�k���C�)�q�:<�}�Z����R�2�"J�a��{)!Ц��+��p�A/i���x�}�#"i&`�[�t[Va�U���F!ʪ"�Q�c��j�ѧ.w�����h���4H���Zמ�����^5J����+,pS�9�v���F�Q�����>w�ǽ�}2����̿ٞ͋|�hX�������Mˀ��,
���A׺:e��s�`����?jf���S=�����3�i@g�u�,{����e�g�em����yc��=3�n�	����o�nZ嘆�R���,�1?^-�wj�2U��[����]�; n�g���C>���;�x�3N	�Ǭ�.��o�¬��+�{ަ7k6��c):O:��'<Ɗ�E���̻V�ƞI�*g6�4{xY1��,���ٜ�5���Ma��ӣ��@�A�V���0�23�3�3.L�03B��sxud�])䣙�]�j��y}��M��-��2��S���������F���'l9r���_�yl��;���$���}�\}^�^=��h�?T0ia`z>�����y'	>]؁��C�P��+}|�f,��eӹ���8w<���p�ߦ{G���y��L�;�u���]K��C��LW�j%�\�Z�C��brߖ�
�xA�0){5e_yN4� U�;zK�&���<Xk�:"1�Yq��8�={Iݝ�r��u"U�ў%���[m�x��^�t��U��3*,
R,X��z,T��we�C�N�mn�z��{M�Pp�)2$���^<�ν�� �X��=�@��\	k��
fbt��.��髙�&Ew%�#�s��=N�fJ��i͛}�>/B���"�3\��O˸5�޿Oa�w�eb�<+ƧTJ��X�_���eKX`���x��̎� ��+k��Q=��>��`���>���f�����t�<w��"���g�(a��0�Ю�K�;��5aDxh���<3��3�m�ʫ^]Y�邒��B��4�/*��ᶎc�'�j��=.Ɲ�J|`y�/h�Ja�Nߑ�f4��<�D�d����p����I����nh[���>�Ǣ`�Z����҂[ݒ>O9�FuGBi*�{,��D�k������t��_	/]u+�e�c��VG7��&�������$�β�W��<=�r����@Tp�nSZ=:�~0L�2O�
����X��[9xhQ�ǁ���GK�Û�GҵL�'ڬS��PgEmLL�|ƅv��:�tN��(d���;��Os�U�w	"Ùo�F��齂��=��xG��9n�DBH����x���<U
��x��S#��w������_{��O5�)��5�U�D�+��������Bb���X]G\);o�O�ؘ��|^W\���������񥐕7����e�~~I��5C�o�ϒᄿ��Rz��8o���1[�����t'���v�)����$�HH�wӞ����>�\��J7�X~'ǁϧ��ꄛ�Ų�k�J�NW^u=���p���:s�y��/[���8?��v�ʋ�ԫ��D�}�G����u�#_AUZ1I��1y�\�;Dߊ�
�G{"���+k�t������3ƌ��L٩v꾝#=�7ɘpz�����x����w��g9��'=����Q��2�S�xV�Ԭl��_����Ù��] %.����\��wtlj�i�TT7k��k�ե4*Q����47h#t��|�d���]�mF ������!��:���K��.��)m4K%�}j��[
�ĉ�F��*g(���eu�V��o���d��L��r�y0�N7%W:��9j�A̮��SՉ˅��3��&��92[՛����(�튷*ux�Qmt:/���+&JD�C�!ks�c:�|��|����;�*b�5v����(������p1��=! ]o#���V����u΢ӋfoW
{01������4W�fd�Y�ϫ|,����^X��^��>��I_ü��]R��I�%�,k��I����q�M�нǛ)<o_��@�Ǳ��%"<�S�%�`�׮��>'��J��d�
e�Fw��t��[T��p������g�h�d���aͼG�z�P�����6�&]�3D�W7���`��"���G�|,����`xz�g��J�2R~x}�AD(��xT�R"a�ǁ�/}�jf�_&�LB��a������E���I���y-���<��mp�zk:;�f��e���9�j��[��ߨJ����ݣ���5;�B@}���j�"`��3شpLv��'��_��f���!���׊���uq�k�Ny��Q��Ϭ+�w.�SA���X��w�� �V��d�h�&*u`g��i��=<�۬�!Fŏ�Cќ�x=��iy.ݪ�oi7rT��m�̳���si�*�(4�BGɡ��b�.���r�|���33�	�1�$9�9�醸	-"��gsº�����9>�/�d䘮��{e�\YwYn�X��10z�cGT��޹~�r&|�tK��-9�&�Q�����B�;�{��<Pÿ��z��,wG9�cK�Ӛ�gK�r��TJƺ�,0�rX�	s����<�c�bVQ���Ó��y����-s�5���!�H�r�wc�S�KZ�oza0ؚ�,�P�}�)�ApRy��:�E��B�=�`�~���F��O^;�Bǲd&:r�FF��8酉�����Ȋ�4��ϛ�JY���v���?b�2v]9I�`�y�C�[Ы�g������������p=��{���6�|�=��Y˕؜�Bwӽ��)�����P���K���ѦV�Ƿ;��%���gc�Ϛ��t&]�T"�`���e$,t4Һ�����!�����,O\
s�x��q�@꡾wFgΰ���Umx���8%}*��u֣c=�wM�{��^lMR�{Ɏ���s�o�x�%�)eKx)_vH���������&دU��٣�]7��¤��l�rӅTUq��>�i`��Xx���tJ����1y���M���/d���b¢��f�"�S�E�g`:*��v)]��nS]֮v��v�0͂%E��y�]�!ն���vE���E���!�٧`7(�m����8�Ⱦ�~�y��p\8��'��G_��ex&�~�^��Ŋ��@t��!��V��6�<{ژ���"�dm�Y���8��o�m3_��3]z��i��� ���ᾚ�x0�rg$�ؼ�5��~��	�v5���f�,�YS�����5�+2/K�ڧ��Ǘ��wd{+���Q��� u����0;??=�6�*ZE�L�W�|1,ly�]a�o�\ĹOz�����٘��}�X~C�o�c>�r{�ӹQA��i����c�pu�K���W�0w��f,��e�N�(ut��w<��\/�Gn!�k�/w(9��©�U�&2%l�Uh��C�Q+��5��l:�����+�zT���p�+�r+�~w��v��FA���q������b7)��l4�/�����s�zѝ�^��1��u��z
��0N�c��ʈċ �)%�ҟ6:RU��d�۴×� o�ho|.�d^��]3S�~ι	��v.��B��xW��XC���n�3�z�����Ҥ��E[����ѼЕ�Y0e˲u�E�hu�s�m�CO�}��\�Y�7��Yv��@}һm�����9��R��s�@w�4Qc�PW}��vA��x���u�mR��vu÷�gG�&���]�t� r�p�g2|��y��	쿤�W���������e�_o�Y*k��a����<u��C�7.!�W�пn���oj{�R�7^����;���c�.'�GQ�ҩ&�#>�:h|������_������G
y%Y!�ݐ��N�!�yx{��iy�F��>�=+�S���c!���h���e�a\����K�C�޵<���u7[U:�{sʸ!~�5|9�r{7Wi>�8�$|���->���`�46,?W;�u���ѿO �)�
?gx�,��鲈�U���qR�O�m;�~6=�s���X������V��V�0B����~�p��]�W��������o������_�&��L���~�4���$���Ut^�U۰�оu{Lf�;���K��,ds������婼4Y�������̱
xǕ���*���\;\�;l�o����~�SǷ���3H�gg]GL��T:/� ۶"JŘF���&Զ�5}Eod��v��`��"���F�kg0�G�lcŇ������k��ȍi�ᘝrDp� 3�d1�Cc��w0�T�-�+˾-L�e�Y	�g�kͭμ�|�}�&N�;Ͷ�i�5N5l/��͐�.$���=ּ�J��7#�펜�d{�O��$��S����3�ߖz��^�o@�8Y#��w�g������ρs�}�M읫��-K<xQ�<�=r܅��k�o�W[yWPT�k������{����`�>�=�����k,��o�P�Z�vz�:Â|f�B:����;,�}�<�.o:�.<�~�fJc;�'��^����Ee>�yC�ht��������w���}7�%�u�'�9����k:��V��C�����_l���8�m�ά0? D�G�z�ۃ��I��U�a�F�ύ�ٹ�*��ӥ���0���$����%�m;�;T��_��'��*�cZ���^�T"�u�=;��Q�ԧ�.{-���w�^�Ka�����s.`kVO�ӄ��@����,˶Ӟ$M����Ĉ�9A�d�e��$���BZ��
�i��%SVM�}�_N�Wu,�V\���δ���o)Z�7��-;�h\!�\;B�ށ�v"o"cb<l�
F󸨹��rMʈj"�6���K�d�@���zs�7uw[]°z�'�Ϸa�K=��޹�g����v~�[�=s$1U�-���\�~վ�3�_f�{{Q�&=��ǺX~���k���n���]��:�كݾ�vr����U��6�{/����͌p��Z�2�ꂪ��k!�1���������iN��3��\�OM�\���Y����7��,!���4�}�
�v��`}�c��'��w�n��h,����V9{;w�Vsip �nm�ݞ���nR�燛�9�˛�O6]�/K�o�M	R3����D������9͟c��09��&���瞄L%�K��������~�������}R��|hc�u��<�U�9���/^H�n�x�����Kf��^`w�u�
�,!��v��g������R�llt+�2f�27z�c��WL�dM�z+*:q=�]�Z�~��ﾯ����BH@��BH@�􄐁$�$�	'�!$ I?�	!I��$�	'�!$ I?䄐�$��B���IO�BH@�t���$�$�	'����$��$�	'�!$ I?�	!I��IO�BH@��	!I�	!I�F(+$�k5e�Ӡ>���B �������8'�@��}  �J�@ U -�@@(@  ( �@ k@ �{��m�_v95��4)E[6�l�� Em��X�n�D�3U)K��CXԫ3]�v��i%T�K3F>;�WJ�*VڱR������Y��L���[��H��6Ѭ̱���j���m"�m��i���6����}�^mZ��  ��C��� v��tv�fv�M볛��P郛��8�`�"��f�d� *Tn�;(ʭ[�v���fw�   :�l  �e����@	�p q�4U,���Z���D��w B�*k[`;��Ti^  � z(Q@��{�  
P
,�P
( ^��  t��p� �@l�mz �u����R�[Ն�N�@(3��]�ͭ�拴��  ����;�����3�P�f��� \�g0�P�ۨj�t�F�]����)ۺ����U�T�5�f��� � )e��A�6�tE��3 ���GTn0��mtn�vt� Q�6�[�cB�f��kL5�<  �C��]�0�"2����;r�w;F��l`'l� �7lV��pPq�ٖ��l*Yb�i*�  6z�9��SA��� B�JZ`���w7P�1Z�Zf�k@�u]�T�ڲjD��!�  G�5@����\ ݧB(�i�5��Un�C�����6�٭Zq�i(�Z�Ɖ�<  �@�^��[nn�@'L홫-h4��Ύ(�w��U����-0 ;*�6(54�,���  �S��@�1��ـ����J��0��XN�Xh�.p�Jam��ϑ� � ��T�MQ0 �0  ��OhaJ��  �    �~JUQ��     S�F��J{Td@FFh����h�a#MF&�4�cA� �I�UJ�5L2F Nxp�C��S���ה��x��g$1��[�*�/��~~�L��׹Z��, I!!�i�]C�����EU8� 
����Ȕ�B�����%v���H~?��������R0�("��(@3D΂����)T�,�C*�^	���i���!�wr��;�Y�"���WEʅ޵
��q@a��Rd�ƞ'�����~&��Iw�]w���#ul�Ӭh�W��7T�-��~��/�+�ՂͷA�GǺ��C,�D�Δ�VC8w4�+�{�4�޷��b搮ӫ�X!�Hܝ��dG��*1�;���Yv��iXQ)
j��}�3L���^k�Yɼ�CFQ9^7j���fĳz�YD�u����F��}�a�3`�9	A�����[��廃Wf�Y'4�+1�P��;V��ޕ����go�����k���7`f�{C[��D�|���)���}�i�͙p��:l���sԖX�u�l|s�n�p�e�<<�Q\劎�ހ[���k��%W��(����F�ֲmGri��/`p�/��E��Û2'�"nr�<{@e�h���t��þ�T����	.����X�P����筌ٗA=9�W]��0�y�u���p|����v�t�- �R��D㪄w�Y�^v�B�j�J�k
f�A�_VW��\&�A5��&mY`9j��(��:b��Lم%4�ۚ5e"pr|��\�^� v�H�Ԯ6��EP�[��xC��y�-�m�1�l�
�K�S�2���qMs$E]�x�Z����i`f����H�@�'8]�/I�Mc�t�H��U�fj����$wU�s��t��C����d��/U��\�܈lp�O:�	��q�U���s]�pq�ÚZh��n�Lї��[ki�]��]Յʋ�L���dn-Ǳn�k#~�,�T� �Sك\��l�{K���ʓƻ+���ٱ��Rԕk�t�0����g.�pZɰ���FY�h��s��\O"-3���xs��Ի�ֽW���b��$r1�1�3��f��ac��!�51u��l(��M��T��vӝ��_4
/�UI�X�L
�R���(�fP:jҎ��
�t�s7"ܼҗ!n�Х3����sh uYJ�1�!���˺�;M�A�n�A����'��gnGͮ����Y�A�z�gr,-'{s[��PŜ��e|"��«ۇ:�8A����7��Y(�݇�N�5cQ�/sfz��	)QH^��nh܄�4"v~=G��Dq���H� �YSʠi�ɚ���
# o q�8N\:���ѹ�?i<�Y�vM��̚�ϔ�d�=��j�]^�-WVuGz!�8N����%�n�\��|c�7c����@�z��a�;���X5�KOr��J��$�����н6a�W�!�5�K����㍛wp�t���&��BS����U����XC�S-١��)͈];�)�n��h)�@6[ñio���\���K˼�tÚ��N�����MRD)T'qaSc�ady������e���JNj��W��Qt�.���0��e��v�+x^)[� q�n@r9�4d�����q�(u�wdźYYX�7�48�X!-�79�EΙ�uڙ�'n>����Qd��D֭�.�k*�k��`�.]�z2Y�y���A���p�jd0��£��ጬ��|����g.#uE�k�娱�+�����!*��6#p�(���PL���UT������������P�t����?B�6ܹ�Ab�G[0ĩwP��VwIs��G�owݡ�y&�q�U9ph�c:5����γI˹r_�C׳�9�c����®s'��4�ނ^quۑ��(7+�j����ӹt!^N�.�֛�$j%4奮.�om�n��ss���1�ڞsz	-g*4����V����u��R=�wr�¢�๱��ʣ�� �[ټY�q�{z�ǳO �V.Gԫ�Ż�=j~�f�sX�i�N�=���lI�2�;�-}�+,�' ࣥ�?]5X^���r5���n,�c���oR�z�4{vJ��w%���At)K]4,z����	�씳U�ݯ7mp��'=l1\�x��U�q���]���.�n�##��7��d��r�4ݛ܂�Qۧ��X������J����N��A���T|C�خ�7g���s��P��Y�*�a�^.w����n�Mk���)<\���mA-&,k6u���^N�e�
H�w���-�Y���`R��{Kr-��M�^�d�ܓ��P�Ep��f��� (ZnLl�w
��'2NF�s`�^6^%���rպb���)�t�@�2��K�Y�A;�1b�T������ӹ��5>�ke�V^�%o[\��y#�=�L"t⳶C�r���a�'\u�2��p�q�˰ͣ�k�x����bL�DpS�r@�U|�U�x�ooJ������2asN-�R#��F�p�Y�)�]�"��kWST�ǟ����/E��4-1�B�Po;��+�����ф��ۉ��4T)�08��sPL�Ốb���s�́�L�Yb��I��JR�5�(w;	n���-ÝYwv����$z3]H�6o[6)�v͙��N���۵��KE����x+��`�������$Sq��{6�/Nvt�vygӢ��n�ٵ��fm]��*ִ>>�C{�2���N��tlao�oܭ��Lf`m�ñ�am\:�"U�B�̝C�m�S�a/���m�3���[z�I/C� 2\ ��n�u�ݫ~��dA�:4�+pq��J�}��朚z���a��4k[�|%��n�e4��n�	�q����N���3*Pv�v뽗J���#��^p��i�u��9���e�5f�<�E�0J��u�v�"���^�!���D�rb9^�T1���L�؁ۓ%�q��2Ul�o< �:'�Cg_=S	��TZ4p�i��.���,B��1�^#P�L�g]�ݐd�uR��W�s�\CǦ[h�xsy��iL�3�u�q�vv�Q`���y=�?���gk74�F�&C4U���ps캒�&�e��]����5���mJ�M�۷����*�·N�gC��E�Cx�:�c��&����jwf�#���V�6K����;�M�^����ov&{7�j��7�ws�+b����r����w.�e�:U�f��]�7�S�L2���=�ܥ6�x�w�� �Y2�7�z�sӤ��E_^fg"�`m�0rk �v��œ�E�3tW���[���ٔ�,ە]�[v�R7˂`՛��.�pi�B�"�S[݃rD.5ܢOF�.��"o�֤I�Aks �671�Zg)�0�W�����e�v�r����5�G�m)��_D�.Hॵn�ň�M�f�y��r	�q�nڹ�?]���;��0�ywuH9�&7��ܳnH�{��E`��h1ɏ�+g��vv>�l���74�Rk��J�M'�i 4${��JP�v�	+:�0&��dy�*ww�x�F��I���W�֊)׃Hv���p�����r��hѨ����)o��v�N�̶�lԢ=�3t$�D�s�X/�t}k��k��S+��۩����{��B��5L� ���
k�l��ݪk�����G�Հ��ޑ���hz�.D���`/4s��۪���������e�t�;�[��<;3�[��K=�A=s��e$����"
�rbq�N���uך.�w�6G�d�u�+��dyH�J�ᒖ�\���9�q��֬'=ǃM��3��Clú�^�!".o��Y�o=ɩ�;7;Ӡ��.
���b�=��E8�q�sx�g���yc2v��8,�qV�#��ϞDT��y/n�)vn-��'62�G7+�!7�=�z+ط�@][2���t��:�8�e�nLto7ۯF�[R!�11:;�Դ|�,�&���o�{�P�1���3����[ͽ�ѕ��f���J�;vÄ&O3��ڇZk��<�^�������ҩ8jW#ݹq	����n`�9nDsV�̎d�2,���Q�����V���>�UG�n��Q��q� I�+{�2����Go�c��C;�ŝ�4�K�h�#w��vM\��sp���.v��D��멍n��ْg\�1edfK�wAe��=�R�j��f�M˹�sPθ �t��=Ch��n7��>�n�� b��'�y-�w+���A�
18�E��qm��r멍� �l���S{��gV���p����lѠ�q�x�/G��p��%.���gwY�ڇfnc�D�{�<{G`�g�ͭ���uL�r,��E�����)o�����N�j+4ɂC�������B��vVW'd]Ki���}M@YR�jTz �ۜ��d ��x�d��ޡ�*��fnh�ݛ�fm�F�����R=mu\�b�n⶚��0���eR��;� n�N�j�˰�s�z�w�����r0sC)�֮��,V1\S}�i��;���������b��ӇZpp�c���Ժ^6D�EC��pw]C�9,�V��J��XZ��n���h�xn�V�כY�6t�Q�rn�l�pYS��onM���ޯc+B�M+�E�����A�>�V� ����R�����˂�r�mʏ:X�j!��Ck%�1hS
��rܭ�-.ԏ=ǹcKVx�7hY�Fo���Boe!F�Vw�b�ֱo0��'d�x���鈙�p@'`�Zq3AGF:�i�v8�{/e�{k,��HOAm`=�G��=��se�쐾�HM�9�sJ^�7����P�D!���B��hU��m<�篍ks�`�^�eG��^�2�.a�6�V-GW;�����I ��H�:�4u���g@�	f�-�l��{�l�Pȴ�4�4��v"%���~��K��1��l�),Q8
��sg.�ܚ5k�{s�ާ�r��S���6��9=ʽ��M1p!����ͨ���v��q<��K�+j޽��a�-I�էw�-�ve6�3���`�׭Ǧ�d0'���gr��;A=�դ��8��Dͣi��ȷ'pLq������C�J+$N�9v]���b��c�IV��h������f���n�\}vi�'�w��R=8�(a��Uhb�cW����Q �[����?��1�g��?�7�}��{.�뒞f��EU�K�[��tf@}�}�����+��=���>��1�Ե~Y�ԑ���A%�w�1�]ey�,E]a4�#a\Rj�����"dv�`�hd��D26�6���+��Svq9ۂ�(��������шt4YX3���rt	��|l�y/2�u�_;�W�N�v]iDҿ��M38��=#]a����^�Vۛڙ\|cx�×l5�ZƋ� �Mt]�.���/�� ���e��s�@�{6Z�\u��(��(z ��F���3c�#2���W��P����/[׼ v�<{�ݧ�R����cj�f�(;AW%qy)����]�垫Y��P�)Ɖ-�X!�Ĭ)�Ǖu��Y� �tWuva��7b�X��Se;Q����$&{Qz&[n*�ȑbNTX����&s�?�e�Ć�؏�݆՞K��`.Ɩ���OZ�Tw�p_�^ݣs"sU],���� hVU�O6�	��H�z{+Mj�J�c����𝝐�k�Itf��F���)��Sǅ��߅f�xд���E����v��+R�Ƞ�S��R���>��	Ϳ�[}֝C�I˜�����se
U���eΤn�N��Nn5���"��{UR˜]G����v�ݎ��M<r�v�N����A-HWh�UǇ�ڑ����$�Z�F�ק�B\�ip�ޣ˛ݝ5M��o�T����y�=!At_Of:�,&qK0'�=�Q�-v�z��G{�psl���6m�	lu�B�@�r�Pjr�M��F�j��Nv��.]�VX&nT���@P4��T���]pb�����x�u1PĮi����I��2��"2n\:=���^P��`�{�E3�܋�}4��u]XQ8����glŗ�H��v/�*�W�lM�Kڊ���u���@Ӭ�.we@کت]�W(ط����>�mܱҲ�k�%����s�#)�9�r���oz��� �|��8�)Y%�t�_=m������_κ�3gR읪�����d�0^�������(B�f�$h��Z����/J��>���6�p-"솹Vv�݁���T��=+2��[�a\c��r��x%iB녭be���Yy��{(A��p`�緷;�=iS<n-|�Vh=��5�\t��SNN��:9 ����s����^��Nx���s��/��Jc��b��r�c�T���%�ы����c+���)�d�ݲ�뫛��se����7$${�hm��������|�}����Q�A�յ�Jyɮ�ris���X��6��=�rW�a�7�G���xg
[�_�媩;�.r�-��家�n��d�������<�\N��}����-d����qd<�O��킇=��F{�$��cdמY�H��Zϳ�0$np��X�����oZ��������z��1� Ǽ��&E���O�ލ:�����H2��궋@mJ;�>u�v�9-���ڹ2K�f��66�<z�����¶�Y�(C�'om�c�f�X4���N�+��յb��(F����o�w����u�H3p|;��c+��A��T%�����]�pZ��J�j��W�I�L��J�n$V�Jeh=���*s��e��	��-Fͬ=;hQ��x��47R"{���1�?Ltx�St��C�s��[Cv���C �YB���t�����L��og*Y(�ns���M����m�Һi�[����/�U��U�q��xm�WU��6�����p��Y|�v���U t���ηU������P�7/�kX�8zΫ4��l�#\m�kx�j�ذ.��n��x���6�ʺҨNO'.��<���W�+hah�kT�w���Y�kH�ٖ�w�9�Qn�$�V+�|*�]>�b9N�@%M�S1*.��\5��ɾ�*lţ����0f9i��aJ�n��Á�r[(����8[u�UgaY��F#�U�(��{�ʠ�d��0��9���X<[3"�����O/�(Б��tȗ�Fe�=!.��y�t]ָ{u��/MZ����ʞv�zڏ֢�D�Us�j�J�Uֱ�^꒵�.���]��<�H{/��O/1[k=�N�۾-/�鸞�¡�U��C�X:V���fz�cQ�3,RU����"/L���~~��_�l|���Cq��@����(�a�.{��<sSjϞ��݅���a$1�D4�c�����	����tm���c�Š̚�N�G^��{��^�|p��y����~�ˡ�­I�:�b�A�xU�јX��آm�d
��em�������M5ծ������:���V]�����>:�m�ü��d��k���o$faeű��ˇe046���2u����}6.�奀��:}o�}�x��j�*�p����̸�UEr�ݧ�I���` T��;6�>~O ���C#w�t4�7.�4�h,቟\�!r;Vl��,]�p0Vv�؊�z9A�"�
С!�"��ĮW�-�W�C�̏�ڥ���-p���λu1��o(�Y02�{x^���с<��{�<J�X3}�*���l�x�]]m-V1h �F���IsX�Q+]�t�73�����wb�;�L�\�gPN���J����]�X�*u�eTX]��T�����!;)J�j3��'��6��O�+����3uWCt/e�e�;կ�ܬ�� G�Y�t'�k��U*�]�;��7�G�Q�_�A����������Y������v�:�u.���^V�:�t̺�+on�R<b�4����jC�k��uшq̢��3G�Jߤ��h�j��3�����#FtH{ާ�{���dB��ٗr�I��G��`�i�_G/���h�U1R��v��[J]�\��Ȝr�h`�\��Q���׍G�i�G*%C�3�}v:��~�LL����ˌ�{�A�І�
�˶L�'w�����@�n\��ö���(�-se�K�U`�JBoQO�}L�CU.N�6��-6y�#v�H�elmV43��ާR�Eېq�Q�mE��u����L�)nWk8u�gAt�G�������Y�R�{-�!ǎi9��hЃ�G/��k�o&:�h��f��r���cV(U�a�	HLB�$�}8�:�=��FV�Q����"BͽA��FVghOHPV��j��!�)�%�h�6j\�;�]c�ڨ�arl]�������f���֮5�c:�1�P��ֽ!�hej<�y{}rɣypj2(p�^K�o Fє�c�Q+(Ф�otR�v�W4r�/h�2�VЮU���M?
y����/�1W7L�m"�M��=��'>,^����A�έ��E���=��Z�N���SM�c3U�xR=u�O�����j��Q����.(5,4.��v�@/*v�����vf�J^�0����M�x"���%pݷ�m�Մ5���=՗�P+hun��SX�nv+㮀Շ��bԋ)�/��n�p�W�z�G�g�$��6.�t�T��:M�r�e��T�rk�Q������M�&#�ǍK� #:T��W���r
�%t��nv�����?R&����9�#�Z�nkM���_D+6��\{I�줄��}ۼ�Ak�}91EK�^Rn��,Q�Ւ�>]wY��1�iDB����o��Ӻ=��Ԓ[���'E�2���5�k�}���S�R��O!֭t��\8w;N��][�����ݪ�4oc
�[G�.	�h��֝T#L7�0�N���A�!m��O>���0�|�\Z�	�=�р�G�z�?`���Ԋ��!���4�V=ۜ�"��4�0*���.����ᳵ{+���'�<!�zrA��p���i�}��U�*�6>Y�,��Y�nE��5��ֶFJۣru�+�<��"�r�N7���S��ީR�'k�T�[����c�w��&yL�����w��4]�X�mo�:ՆxƘ�P�ˎ��\�Չ!�5U��X���@d�������?E\���Ӹ���ړ�՚	�3�Q����\���4F�0�	A�)es8rvZd��3(��V-ѻ�up�����	�5��t�J�8~�6��ޞ�^R�[�c�׃t9�w��@���-��0֋���|c!�CU�w������AVU��Ewd�ݝw��y3�DF�7H������o��z9�L��a�y����*���dCJ�?a�/+Ŗ
2���0�ۦ�Ż�h�L��m�vH�V�Ӊ�.�l��1H�6N.�D�oz�vh�&WL���,��*<uV�oY[�|)۫���H�B�}���@��;V�Z.%�B��k�����L��<�sl�f#:d���w`��2V �ڷf0�3�:yj�[��E���8�;.�ٴ�6���8N��9g�{^IiЮ`s,��;���'RvݻOⲷDw!�=�Z�uS�.Q��͜,�ؚ6������	�Ej��mL:b��"�zTh�'����M���(��"����V�s�ڬ�كM��OI��j�}7m��D�\�n1������!/�����;d�.\��P����ȕjU�����Q�+k��8�Y9��չ݇�&�c����A�1ӡƳ��-��*�b0A����[Z�T��蹥�'�16i����E�N�1>�u���r��� r�e��n�WSVԎPoQΫ�ëz[[R�B��2���f��qw����1��6����o���Fu��#���<snWw\��9-SX�Kt�OFޅϐ\a��Rhu��,���p���"�n�F�6`�CR0]��8ۓ�4v�=pfͥӵ'�6Ǟ��Ä�#�Ὥ6�Pm��)M�J���ǳ�C�\��-��gH��\���nl��I�gL��0)�UfK����b�ÇL	����8-�Ҵ�_�_���"�8� �k��V#mR��d�I.Z��m�FvT�q�����D"-޺x"��?���K�~=.5�t)w��r(�*x8x�r���R����_F: ���_Xo����:�И�I)�s*%.(�Ju�ɰ=�&�:E�����m	R�+��5I.tM�@�&9]��թ*��%�)%*�M�^�
dĨv;�fE�V��r���ܫ�cY��73�e2��/�~�NWY���N��1���TTR�R¹�PT�|ꈽJh�L���;��E�x�ٳ=:��j@�*1������x+�=�gE��C����t����h����$�\��gBXM8T�ז���İ��K��+�.�C�>���qa�w��=��d�W��#HLi��R�7�sƬ�(V���D;G`�)���;�'�cIs�r��[��&�\7O)pjS�,S�3���7���H�y5�L{��O���zc�$�n�Re�':q�̤���2�a"���:�L�(��1
�1���ֈ��4Gd ��ǣ̇3����z-ㄞ�#�R|�i�i���@Y}���~�8V�����/��e�ν������V7�w�h]D���()uG,uqgu����ҡ��q�=�z~�9ڦq�崱��R�Ը���66�︺��w��j*��n���"���m�tk"G�1�z>�%�{Α��;U�vur����2�d\aZ���5�O���WEjU�E�3Hm��9��vt���\jI7�v�����Ⱦm���7A�)��v���s���hq�U��l���Hĺ�2M9c���c�N�Ur��3/�=��9àu��e:o��^>�`��W���9|��q�Z�<[RAz�B.�u�cZ��9��՘�)���Q�v��؄Wм(� ^8��wvc�5����ebK���V��h7z�0{�;`k�����]�yI5aة7$\�g��D��.�z�q��Io�u�f����x�"g�"���e�;y]y�8��\�{]�Y)b)��XAnm�:�TiЭ;�����o�[{�h��u'�3�Yᛅ�3UBp��]ʠp�}�:���j3|76PY����T�*=��V���8�a��q��A"^���q�;|ȹ7��=�*Q�7:�J�y6����;���XN�w���܄D{[����˚[N���||(�_{\B�ٳcO+���1��-^��l����pfKzOL;��Z�[C���c�o�F�.Ce������|��m��-3E@ w��-"�1:�Ҝ��)NX5V�9uM8���zC��m��"寝ܼD�7PJh���Ę�Rx)N�[̓qOVv��}�ʀ�F�9[8���.�H��{�cX~��^w��5yk�s���;q����#m{�K�k���ں��f��H.iA�q4��{��j�����X�T���#D]2�K�u�NM�q�1��hST�����8�A�w�	z;�)��k�*'�LG)�e��&�k2�pp�WZ����q�"�j�Շ��ԕqSidHe�W��d�����s�-
b@J��M�Q:����J��q$�V(Iu)�2b�A�y���9���pF�z�lmW�rڜR�B�&�{â{Ŧӏϝ,)꼊@��'9[��*��޼0�/Դp��<9�7�n�^�e�C�{u���Nk]��`r�{�@~�*pZ�|4Z (�Q�N���ՎÒ��YX(P"XN꽓.;YWXjl�5��!ae�^9�x��Us)�3����$���@�ۓ�c��7�F/yb��1eX"=}��t4͹[�Tq�u�; ��*�^,�q�;&�ɠa1Ɗ�hYەЇY�P�	I�v�Z���'ul�b���^5!�l��=��ƈ]�ʻ�u]�/E^�s$��&Ax~"�L|����e����p4:rOt�ӳې07z{x�-Q� ̂�XN��ل�h_ٷ��M��9��s�<�c�AH-o#ĥ�7�S�))L�0a�x4=�׹��+Ā��ז��p���:�6MH���9xvu��%ǵh�E�wn�o���B�+��U�Fj'd�$�\�8�`�:f.d9x+��{]c�C�R��N�H6�bX��Ψ�]Cu����r�:�f�֦��{�$�N<���S3�PG�\�b�\�gm<��R`n�4��+s�Ǘ��I����N�X�ۇ��N�Ly�@�^L)�11bK�K6g&W�1ڎ٣D��t�3�9��Նp2Z�u��V,�m%��䝯�d��5>Șpw,�p�}�\%�Б��_=��k�p��[��6��҃����<���/-��Xq'���GnTd^���u�_#�k��O w��q־Ԧ�;+D�v�,��JM*u8���#6.X@���Q�mŘ��ވʓ��u��;ÕhnoQ~{�o�$%��e{{�����Us�X�d�[+M�]�}L�������h����\:����ښ7w�u:���YP���X�:���??�
���F�Y��YJ�>���}�Zm�9�X� �1x�U'�Su�8����=�PѷZ��|ɣR)�*�]�M��v��T�*��ԹW��fus&��V&��&��+�ѫ��������"���V�bɎ�#��;n��Пn�Z��諲��Q;��jQ�B��vv�T�N��f�F';�y(��2���^]P>�8�T�{�Tc��?7~6��Mr�'X��1������1M�cDU5KZ��ۙ|�%K��>��&��B�:����[����b&u櫕R�uLf��bK�=����s�^��\��u��9�#�̈́��<�9�J����뭆5�\8�����	�|���������}YGCx���B��BAfZ��9���˝ƻ�4�˥��F��8���&����h%l�*;�6��#����-r��[sh	O6�� _gn�/{�է��wgn��B��Ѝ�y3v5�o ��.��cz���D��x�H4:�����:iN�m�yM�8�p�ŚC�h���72\�6R�e��\��^l�OUin1��nN�M�#G7�q(jGV#utPBD7% ���2�,�gl��P0+�[V�3M^=�B�FC��}>,v��l�
�J���Ql�{��k��0LYK0/{׽���pP=�t��ӭдr��x�o�v�E��X"��g'y�k�Y�3�|�>&��@;U�"��~�x��݇Kpw+�Y'�[~�:�u�wC\�.(�2�E�Yk����pk"ŵ2�ٸ�vßdNliY������s���OD�n��sRP�<Z4@��I��ԁ�㣡{w!�r<]۷�0��!�M���[z�)�7����@�����]�����3��W��oW���`k8&���wm��-��St�+dz��	�ǵ�)c.���:�M��oWq���|!�fκ����]��'vJ}\i��!�o��K�n֩@�Z�[ܼ����J-�F���t7�슺�[VKռ�����sН�=ݵG���r���Vx��D��N��Sa�N�V;`	��p�J{�p@i�,j�������K�FtA���� ��`���Oi��-�2�wݓ}rmy>�(�ч�c�Il�u�:;��j�[��
���#3y ��7�jzP*�pϓ��F���Ulu��IMW���u��࡫WtK<��r�D���][]����Z.�;�����R,���Wu^y�|��h�Tؕ�3��3���ٲ5ROF<�;�ZW�׸��B�~������x��H�ˮs�̕�7��I.7M+�-��'��#1�yP���d��U��&��L����V��������p�����B���=�~�n�d��I�����0�v��ib�kwx�,
�%��Ʊ?��	�#{��r�tbK6q��ŦP��f)��٢��`�)�"�a�:\�O���������ʜ�fs�x�<����Ѭpb4��Cv>[�]��F��JDJ"��M���Ԋ��--r3�����7ԛ_k�b���_Pȋ;[Ugh��,��&�l"a�� �<�ϼu��=��Ge����(0�4x��xdb�V�%�̽�s3T%S������5>A.�.��	g��m�����j�u��v����6%��������b�GiT�6+R�7�T��j�:�ސL�.�������çs�qi�K��T͵F�:KlM�(��to�Ǣ]\\쪩dG.[&��)��:]Y|��2g+�\q %��.�N��W�P���Ɓ�SW�%OJ�{�X�m.[)�O�3-�5��fm��6[�dq��N�r�V=�]�S{r7$ou�6��p��D{*�F͋��y]Ff#L�xGd�uˑ�9N�QΪqg&c��m��TփeQ�.�
�ڂ�.�.�\$�PCd�gk��*��ݸXШ�E榻f��k�]B	�[ژ4tYXLV�[��e�Y�ڋ:�azp�8-������_X����^B����20���^�oy�܌��L���
��%k�c�ݷ�V��*B��nX�֥gL��M�]QK�FbP��ΙO���
�A�x�L�#B�ؙ,���ծ�{D����Z�
Q47��lk��H�d�3r���������wV`-��4�-\��O��0���b���:�䤬.rR"V9�%��+�n���ix�cs�eѫ�'v���,��Pt�K�*B2q}P�3h�)L��f�QS;`}�eb/�X�¥�Ĺ�`��b�[��˨8먞� `ˏf�E_-�H���nJ!��5�/��A�k����sz�O���CD��B@�1�
hh%W:���6{(h7��uIAce����{�.�r�,
����J\�%�b�K.��+��-���s}�1lE�b�Д����u�)gYd�Pj8���ʱ�mq\�C�0�t��>Dt�[���۬m�-�� �ԉrѕڪCp7�'1mp�8i�1���H�,d>d����4��0-ٖh���R�����/Rx��4U�y@����!|��og��Y\:�ө��ZM��Q+ۍU=�p��v��:�4����ϰ�,����B͜�o6�&�(�ԓ��}Zs_9V?QN�ٴc�ߞ�wi���;V���7�I�a�.�����:��)��5(iN�
�Vww6{E���n1�4�楲��'���*&t*�P�6mb4��l�>����b�O���Iv�eк�T]�=�� �q�ɥy�G��Z@��幎� mGv$�*k]uœKYY�h��'���[� ��jvn nw�f�u�Mn:��fǧ�继��6��4�P�2�����y�F�ו�;���^����W5�d�i�D�yV���j��8p�y_�b�6iQ�unԐ g��2�~�ꯐ���!3�?p A[����[:t��o��7E�<��'�2�ڊ�:����:�����6���$?GZ�*)'�Q��"KM�>�M��&���o��w����dQhS�4Ht�n�E����9�*�9t��<k���˂� �j�|)����1n��l0ʭz�Gډ����w��+�D�pUa{GMIF��yXj��QQ����,+�9Z#�ՠY�=w�&P2h|$��,���N
ۊ�&�^!��і��n���4gav�!a��s�:efʅj�EQ�I��=�չ�k���a�Q��Q��\�otO�W;L\�o.�-�w�4�G��ۏ��v�2^���B�K���<f��Ƕ�Zۦy0"��l�AMIa�x#T�3���I�W]�9��S&Yv�uj��J�p��k
�����w����`3�+�[��O,yܨ����9�-N���m\�D],g<�G"�����p������@ݙuvS)��r�sj��)!�4��ǪI�ܯ4�9������{��w�y�^u{������!�Ai�vkв1]�9!۫����AF�i5���~��罪�i
������CS�ݝ�8]Ml\�M��fC������Oօmh�Pb�*��(��[K�d\ej%3+��l��Q��Z�ih�3�3+iF�ъ�e��@j����+KJ��V����)ib�JV�Z��KQ.����Vڤ�k)-��*�Ѳ�TDm���[Z�T�+h�ј�Z�V�Q��`��b�J�TU`�)(�Ų������V*�4�\��X�ʶ֒������SQ)�[m
\k���&&LeJ�Xҡh�b��V*U��U��Jҭ�b���q�մh�mc���+j1U�mib�h)Ecs.J�F[j�V�!`�h�Ńʯ����?�eN��+�WWe&2o.)��n���W?llJ��.lL�O�����3��t.*�J5���w�����].=4�S�칦~���ϭ�\/Q�c�l��p�n ��H�!x�D1���!�����L�ޑ�5T�Ǚnw��]�7Φ,s+H�\��ɧ��"i�I>�;ˆʞ�,=�=�N|ϝR��4ȡ��T`@�=1�DF�>����g���Z��1� ^�����zd��!r�k�!@؈��#�JM8���I�c�-�F��"�k�Ԃ�M�E�Bt���D9ƭǥ[x��Ҳ�:G���d\󮉋ڑ9��� 9�H�u�,ql�̑9Bc�Nִ5�#�[�� z0@�n���O,��p��٦��  ��cn���o^<��_J�Mȩ5���a�����W��Ό#�L<䬦q5k���%��K#`�����J��x}d�!�?
���4w?p���)�o��k�q�˫Y�v]l����^�K�]�n�~����k��;������vAbz�MVQ����;���F���䫒R������*|o�iB�?�`{7�^�mM�9\K�܎,qUҷf���z'gG�Ί�
������E^��svE%��'��y��]��Q��c>�t�竓�U_G��͡]{��y����Ý��aC��퉥#`w ���T3O@8R�ool+N"���^�Y�I�b��@�s��8�=���V��2�v�t��@~Dn�I��4�H�	p�t�b�ۂ��s���+&b�]�o�Ș���9E�*��t@�!	�3r}�[B˾�ʑ�o"V�����7Q�]n��M�P�Urm�ph�"���&W<��ԭs�s[ �|��2l�Of��%��0G9P�!FJtEbe>]j�es"ɸ|r*�t�*Bdʖ�"X�JC���t7U㧘��b#��J�G�$\�*�8���5�!�C��\��"#w�w�7�f��R��_w
��SvSҌ��JE��؍=�����{���ޑq����,m0�a��Ov�s���s��|xRton�{���i�Y�uF.�]�E6����:�fD���#v�b#$���#`��C��Ϩ�����e�xtt��"�0�,^��׶@B:(vɇ%��'�L�M@��
��i8���֣n3�A������/b!v��qe��/��P)覐�jM�i�/c���.p����dl&f,#�9��#��N�Ы��e9}ʄFΓ
:��莁o����s�ƪ��[ʅ��渴���Z�>�P<�����49�]^Q�w�3����O��үS��wK���'͋�\١$L5b�Lu3�p�w'�\�tR��ѱ�Yo��W(���L�3y˒�@���*��(�;5�of-���.�H���Nr'N#��d�;��#��HA��S:���쭗;�$v}P��fx�셅�5���aL�TDl�5���h��џjўw[�}.9�Ղh��;�+9�:YA�ɫ].2pk�gZ���c��)���gb���[��%h��V�o��Yoo�N<V��tŀ�y}
����%ۻ�eOS�zt��Ϣ�f��ͫ�S��F/��
��Q\D��!�1/]����޶���3�$8�#��:%aq`Q	��l��6c-���J�[H��"��>0�"(�>l�za�D�l�.:��éH�X�XFK���o~�q������5r��"��!�H�-�2
�Q)]�O'����U���B�$ʌ*�u�)#뻃�
�K����D���^��F�x�U�3��p��t��p!D������^75��f�G5�/��: ͺL�CH�� O�#��绌�x^�ȷ^���_��z�n2�(dU�^��$a�X��	�J-��rN�諾�3� �,:��$c�Y��Q+��gڿ�Rǃ�0B)��+��Բ��D0Ԋ�C�k���#-sK�e{ʓ&U��u��;V��~��۪�**���*C3P�|총�U��t�Ŝ̎U{�'��7�j�#��i"���CMt�+&����&ˮso)��{6��L�:4kEo��è)
��sʻWo=�u^zl�nO��d"ep�$�Yl�����������x��yu�����⣢��t�l��}�$8����Ή9�l�J�K(�dO��U��n��-W�K�@)X/�C(6^�{o�V�]d��	�/�g���TH�a�"��W������@��'9���9���i��D�� E��R��Nz+�+�W�hY�~���e�i�$ך�)wO�~]=�V�@�h�"�#��061�����O��j��ȍ�u���ئ�Y<��T��/�/�a�ܑ!����r疬/y<�q����'��S��4ϭ(����""0�|��es,J�Ɩ�!�9�z)ߝzd��"��@Й
DGD�.	��<���#��a�DM�G�>��[��'K���C��_N����B͗�nu�^dujݍ闒�	/�[W]�.�s�76@M���.�m>=��xf�3���#:ۣQ]m�q������b嗔�\���V��`���9����	�|�֘��g+ԔE�yC���=2/�����%�(i�zD3#X��c�S1sw5�j�>Gq��-;�W	Q02�*�qv�S�Q\2i���ᮥj����u(��� ��w��=�� �룣�Z\~l�xhf̫���Zܙ�6���ח{u,?��C|Q�Mt�.�#뾂�+��v��w8W�f��70m9�|�Z~cFp1�¾��i�7�+l�ERz�SBn��$�JF�.�6S9]���iUŁ�B�U�6�K����M���f���&6T{#}NF��8Ȟ��R��E�nn�mn-�)(��^;��` �8\�@�v1��'�����n�u�P�ڛ��!�))%#8 D8B.H��b��S��7�/�{�/(w�l(z�l�	J�$Z#�H�	�HLԟp�uD(syx#��&����x�OK���?�<t�9���uq=-*�Gy�f�uu����G�^2����VfٖC�y�,}�)�7 �8��̜#���)�f;�p����Y{���Թ)�H�p�;�׶zm��\��K�GS�:��mň�����|Г��0��3�PmPZm2[)0D�t��E�n��{�\FÏ8�\ltNB�O���A���A�lsz���)�(���BFǡ�=�� *r�O��8���5�!�\F�xTa�/�W;���:tE ܇&��D� �3g�L���XW��u/#�8
�T��~�=:�ۅ�1\���.;I�'H�'�L�u=2�D���9��j<vP�Sf�P�y���}�b!}����m.�&WtLdn������}t�Y�0�H�1�^��E�W�d�<��y�\�E���������{*�(X���} V5C��;\���F��;e!wQg���5�9G��"����ri�}f�
��٧c���D�ճ���Hڧ�aϓI�VtE�hU�]�¶��X���*�Uӈ���ZqV��$��9ݜW�љ]6���.�fM3���#2�E�q`�;�ܨ�e�\�.wQ(ԇp/�Pa.�tS���t3�I]P�냑P�7'�{ hFV[�Ab����J��
V�>`s.O2�v��3A��Tn�������je��Ul/,7���ܵ�?c��Y���2����rso{��
�|�"����E3�\mL�U���<��U���VS�`� Y
2ۯO�v�`�u�R�1�R��p�ls޴�֜y��@���(�m	�9#����R�d����L�m	`��2�{�8��E��PBs������3� (�qL��㬿gp��N�7Q.U{])�t�D��,�F��E2ٽ:���H���+>����Q�z*�PB �I����8H�8}�����qv�5�"$���;��P�,G`�H]�!u+�B��P����~�Yv����`��M��.9�)����.�UJe]p��i���N�����v�BP�)Wbq���.إ��h�E�ܮ4C�p�:�n����L�rm=U��oc��Z��eݥս�t2k���j[9����ʈ�>��۱ �mn�F(���P��Rj.�E�r�K!�D��>4����J�*�eg�IR"�L
��Tܨ��r3FˏdL(څ�^Z]�6���ZN9C�
�Q�EI��9���2�4�6i{ʘ�֢�I�ؠ7�[c6�3�������S�tM"*�Dϗ	�@�e��Q�S��_Uݜ�ݭ>^�����:���(
+6�
w��Q�/7�����ζ������N3OU�(�}B�q�l�hT$l)��w���=��Ԟ$��&��6������1�6'�*NY��^�B�T��#j�t�j#r6k�.cH�A�HL�zY�����Y��ˣ�?}������Q��Ϲ����DA�㠡	����
;1N7�9�skq�H�"�d�� 
�;y�6�V�1Qm�5ݡ-�@�Ӷ��{���~4���*aR�7OB뺦���g�W!�g�'Hnq;�Xޓ)�7qW}N5	���B�{�>�3F�|�P�L�E@1�9rh?�D@�&�fv'�����JS�����64��gϦ\b2ϫ��0%J����2���,�{\�Tiv}3"Q��YQJïL���!r�I
����S��s��G9�e����(�ps�a��A�� �q�m�2c-C�G16Xj�
���D��.&+*D��l���fi����㸁����P��d%~�F���ʟ��[�x@��<=j��{{�i��1f!i�W�&Nz6=24H#�q�~�%��f䴼�C'��v��G�7�k���5��b	to�!v��R��x@P+V����a��͢�."E�t����˩�٪��Z*XP�u4U�S���f�	V���QdE����
Dn@�,�k�t���\X�r�G�<@1�����sg~���g�K�ݬ� ���[ՑN��uo���ݽ�Z�a1J�3|7�Y�΃}g*�uͷ�ߦ.���qos7KMZ;����p�+@�u�u���-2m佻: �l*��*�/p��4j0��}��ʋ9Y[�uv��s;t����u�<�xq�Pr��z Ϧ�p���!af�,��Z����>�OD�n��� �ӺG�+ofm֧�t{�j	0�w�r���ޭӣS��v�[�,9Ă�j͂��5�R�:`J�LM�O(e֖�(�~ݦȵ
�OF� ��]����1s�Q��w��GVN�{�ɱ��� �
	�T���OvmtW{|bݓ�r������I�ѳ������]�	n�O	5�(W|��ە`�`7M��|"�	�:�+����I��1V��A�ܺ��a�k��m���hV�g7��pcm^s������l���hTRrZ��!����8�epמ���vv��Gms&=����ɱ�f͌r���v�i�f��w���z�V6��e�*qq�+d]��h��I|�����;���鵏8"���38�=����G�����T>���fvEDwP˦��~$w�Th��=��׻R�j9�.Dw��h�*������H�N	q}�`�i�<��	��������*�΀�ԖX�up	�M[���Mq�^��aA����B�v�eU�"F_Eu�N^�������͐I�l�����H�i�^�s�Or��u�qq)j���V��A<=|!D�㙵+������qO'I�H��]a=]�y#�$խ����,]Ф�\�k�+�̣"]�����A��}��o���J���G^$�v�v�l�x��]q;Aa5��b���u[|w��VBw�_h�����cS�Y�E�)�j��G���XN����s]oP\"9Y]���g��1��x�K{����Y�o�+����r���De}��mĞ��N{�oz�yĩP	{g)���k�.$�e:r\qwD��Q4�L\�p����yo{���c��|M�01Bd՞S�Ө� Tdw/���QL�+���gWh���k
��$����Ef����މ�" �;eQ�RԵ��jDU�f%��QB��e�f4�X��F�X����B��UD��-�6�ƌF"
hT�V�ҋ[V*"����QknSkm�T`�Z(�U)U��mU�L�2�E+��-�6��D�TQDX�nYD\iچR�"
�
+���"1EAUUX��X֫"e���A*#V�DjY�pbV���U�T�QXZTDT�#U�m��EV"�T�AdV. Ҋ�*����l�#E#�b��-�F��aVVJ1Kk"��2��(�����"
����""��P[k"��
�V6��OI"DDG�{�M�Bq��;2�?�M�u�d�ߨ�#�Nuq�K�(��}Y1؏ �	4����,D�m[���/A'�*�(���L�2�I��>ؚR6��C"{dS�SU`����䮤��9 ��Cg̃�jL�
����ѣ�>��Dl(�0�v��[�����P5��@��&B_	
�D�x����$t�հ&s�~�������&�4}pӑ�z:x9�4�HP:��'D���4�����^O6����qb�CV��=6��.1�W%2�c�h=7�w�遏�+MI�3(�v���f��%��"-Ѷ,�_W%�*": ��&r$2�����,�	��F3R�Y�!H<&��v��3�CjF�\z8���.T
�.4ѯa�l��]��E�sz�8�p�
�<"��!ɯ7>�H�,G�5�7����� �N�N���و�k��) p��&��O�do��/���z׭�{	]��ב�*��p�,)���)S�֍�ޛ��Ç�LZ{{h��)��/����c��rtl���c9�-�H�l��\����F���[:�(��Ņ*�|8�o��	Z�-�u�d~�0��i�C�F�t�Fp&/ݲb�|L!ݹY���; �aBϮEut�&�7�>�E>���;�-��x�:�$`�b�qPp�����(X��#��� ��ԸZ�;ܜi*�1\f�Aa��>�,��+ENE[���[�2���l�w'�K��bC�s]�8�U���l3GP���H�Jd�q�ˍdE��Q��}�>O'aEy���DO��i��\����`��Hp��Q�8w[�o5$�`x_c${>u휅�DB����JB}���yR!7[w)f�\�1$t�u��fQ�!YH� �je��L8*��]�{9ֺ���^�1�.z��Gg�$�4�+��SH��Sn�^�|�4l
AFll\i>�N��N�	+�Bftp}z4���ӊ�+��������Բ͡���+�̕nj2���r<����[����D����2c���Vf�.
�V�7���l��앝�=���YVȚ�c#w�;WfvEq�3/���8�6�k��
_BgŞ�H�-��S�+22h��-�h��tT:��m!�qLȍ�)#���� ��<�s^�f�<���h�V7ث�����r��=9F��g�ܧu�6]g>)��� �VXEE#q��{,GT�WD���Q��*�F��7�w?@P��
�5g��J�3j�7�a
��bql̾�*�q���DG���b62-��7^̡�iϦ�q�i�8�jclIu]|�q��*����NE���ԑq]`U7t�#%��.=GDW/�%�e�O��&�q)�
��H�T��(�#�NE+�W�7���s��\�ӁFH���\��VP��t�4EX4��!+��PB|`f��,��T/S�{����޽��~*�LT�h��W��;��`���K�C��i���7S�^Ňך
��Ȅ,�� ��u�ꈌ�+x�b��ʻ�*��*vR�i^�N�,u 	O�)�I�
���5��s��,x�Wnt���6mFR8_!TuIw@a����ggT=;/�RHlQ�Y@L��"h�}B�q�,6n\bT̥a;�u����}Ew�ނ�	Q�BFH�\z��Ŵ�V�q�}ֶ잶�y��떪Gajg �f��� E��!K��M9���[�L�$�Dڂ��{���I��;����f^
�_}J�V���@�Һ�W�R#��R��Y2*)�j;NTmvP��l�E@0�rX~ �1�H$v�jU#���^kK&�8�Ƞ��#zF�+�2:�ƣ,��Eǫ�T����1י�s2��L$DE��c�(����:�ψl�Kk�v�vo'Vl��v���a�D7J=\��oz��b=�ʚ��ɴ��y�!㑓^N�x8�Dȼr�c�М-��L@q��Χ��PDac8HQ�GG�}^��zCuU�M��z������խ��g#�&�Ei�Ȩ�d$�j�D�7[n����5Z��AwV�Es���T3�\�>��*}���y���������Gx�Q��:�խ�]��6|j�)ܵ`enc7�8��:�mAv�y�I�4_�G�n,4���/�!n�����\񥩾���;���^ː�f�F���O@3��M-�����q�+����m�>d�5�52��F��u\lzb���g��
��F3TJ3Mk�L����Q�Ӭ���)����e3X|���v�\IV:ȋ�tt�Q7�:�e�E�C����(䝇g�����:��M\e%3�Yi���B�r��v+>�A�&p' `�;;^�n�LZ������Ĩp2%d9���ȯ%#��"A	�B*H��\��7d�ͷ���ܨ��Q��}#(��T�l�JT9!@��	�.��W�.��t��1J�A㱂�CV��#�ѡ�pҚ��N\H=<jQ}7C7�vl�c��T'�"dFϥDT����PR6mS�l�S8(��@������A^�e�]e��]IJ�S�{;o+6|U����,��Ը�bն_��x{��_���^4r�Ȭ�?nNDr5�t8�00ȥ��}�+!�.�<�fM!Λ\6����V
����R����5�C����뎙��������,�	��F3b��z_[;��chi6!"ʏA�=� ���E[���N�j��l��
#`Y�쎡
X��94�D�$i�=~�'���C���mاܻ�ޞ]E��Qv6b%������0��]"�X�8}�˱64d�.�(�|���0��0����4�<|�8�YY㵷d5̩ҧ���h�2���}r)�d\B&�p�{d)������pM���<Њ�`<��aة��6$�u���V:B+���:b'di�ٳݳؘu�2C�V ���9n��rVJ�s�l��w��[]Sq�z��O���۩u���(F��ю�7���׭�VH��I��9�Ll�eN�E;"��i��\�d@������+ªzn��+�ĝ:9�7ew{X#�1K8v�!)_.�7�׽r����N��H��o����=v��mr������1�3�W��
����!���(]L��W;UaMG]vOd��f������}U�[O���-~�����C�����k��q4��Z�Y�'����Τ��s�b(I��aq,�5{!aH��WS,����rg���BFϺb �!Ag���/�:�TA�*Yc��"��X��$ŭ�7=G����C�Q�O� GA���AӡRV1�Kx�&�+9b<6�����o�\��$/F�����=�
:*�c��Du>��䓹���t�vn�éu�D8�])�`R��}�h!�nkwH��>y����~�dK���y�-���Ӑ�a�
Q�go�$���lr��	�2fBEÉD��ACe��B������pD,��Ņ35�z҈��:u�(����ʐۦ͍3Q�� S��L���W�|�m�G�&�B��eI���iצ��'2��,C�ٳ�G��\�ti�ܱa��Gr�����{Aȱ�1���<#��;�	WQ}�K`�.���yh���)y��u��:���D��X����Rf+]�xT�谪U\�MF.�{L�yv�DP�<=�;��6��>��s��h* �8�I�!UJ���#R4\�B�q��71�0�8qQ��iș(.���ڌ�ȥ3��=�Y�����}
�53�2��
f��T.�wj�\)1\�G�U�~p˸�	���zצN�1�����dt��7N����}����X����'�$@4c�=!EˡfD�L����V�W.A��<K"�{�*�뽣at�X�;$d�%G��"�*0Λ�P�n^��E�Hw��f��Pz�ux��"H6#*d6z=t碿�!>ߢ~OiFLr���i�k5�>sn�>�f^B�az=\������4+G��Ki4�Ѱ��������\mvP�-���*�N\�����E�l��o;��,N$L�;P��i�O�T��M2*-_ÇY�;��+i�����<8�s;5�C���L�	rz�H+]j�f�#�qy6�_����*]}�¿6���Z���$�7{���cr@;@E�@_j��]�]��P�=�5��i]�K�HW�x ���m�F�fL3#��}
F�@|rʊV��$6D��#������.�,̇Y����Ro��*�>��Ҽ~w~��Fa:�^+�v򵫜"<��"Cr�V�Ty���D��.&:��Md�G�nM<	v��qq�H�d>$qLף�̵^�F��~T���|��b�cFL>[�7���ת�Zhw���o�:�a�B����
Xn��m�p����1s8�A��.C��q�= ���ZBW��^�f������d6D��e�XG:�޼C�)�N�i�3�,r�(M���bH`��,I�NF�p�	S5�>]��ܧ�S��n�l�6���+��v�y���m
r�v��荿Zc�·�6M�bp�y��������\��AX��r�&c�L�	�;�R/٤�`�:�L�����|�%H���;������&a�/^�+az��Ād��w���Pf)���g��jfX�[p��a=2�aE@齝tQ���޲���e�_o�"�E������Rn�O��6v&��ZC�=������Ht��	%�����F^.o��(�>r.}�!􌢣�S��A)P���(�Up*�DC������Gć�Ǿ�#Gb��	}>��j��Urm=���'��QD�>S�4���2#gҌ�t�ꠤl�>�3�;�5���4o��LܨQ�
��3�,��Ϭp�p.>7%]��}s��YbVPD�	����!�z'O�H�P*ܸ��Y�8n�k5�d���f�����刡�C�^n}�h�?{� }�:j���.�\��﷖��d{� 
(o�&:~@�O̬�Ý�+
�d�S�P1���Y�1U ��?[1!Ƥ>�.�8�&3�}�i �i����כ}�}���y�}��I�f$�.���?r�a�������s��aS��c����Sߩ4°����`VbM�t���Sϊ$2�z~�fw�����>�����$x��i�Q��Ğ8��Qg��b~d�6~̂�P57�6ý�Ă��LJ�*J�~��Y:ʝE7�$��d�aV&p��^{N��|o{�G6r�]�,҅G%�z*�U��0��geh�F��Ãc#�-AE-�Q�͘��MEX+E�6�i9��A�w��eEg*����[��V���ʍ�]s��RɎ�٣!�e���S�)��;E��{t�e��ܞ}�!�{���d���g�AK�R~a!�r�2�kyd���m.�P�GrA�휻���6�|1\ۣv�}��k�$2�&����F�Rɝm�y���U'<���ԫ�P2V��.<.sK�R�(��VU}Ӕ�̲-��]f�W�$���5�v���r��E�]2�y�V��in�X3;⍤���]}|�+�4��C<�d�r3��{�lyu��vF�"����)��e#3�ќ	����j��h�=v�����QÎ�M<���,���|^�����Mn�Q��t���BF+BR9Ǻ��+V�S�m��L��Bu�ԩL<Y�)�1bߗ>ݧn-��FZ�%a����[�WS���e<����}E	\��V�#���\�rԘ�U���!�B��[w�r�Ew5zc�Ƭ�e������"$=Q�S�n��1�ք�;�G��:N��BO�n���c(�v�3��9c�m���^���b�Lړ���,����䕑{/Rܭ��JW /Y�&h��6��x�Cj\�wQ�\E��ьy+���u3��C<�����.J�;�^�yR��d�]����l��T�dQo��~9���r��^��*ݽ����7�	��&@y�[oJ���ˣMFJ�OپȅZ����p�w�U��W���Ҥj
-r�=<��Ml\i���֋��R�݊e=LIw��BYעX'.e�&�.�]'e��Y�z����	|FA}+J*=O�ı˿➛�h`|��@Kz/_W�6�s< �l����|K�͖5h�R�a�� V��"�_�aӵ��^�eKa�%-¾X��wq�B��۽���o�s7���c����~�t�&�i��-�-�E䲈�k,�%����Q'P��4��r�bU�,V�Pˊlɘ9nJe|mk���Ns��هJ�Rv��l���M�1��P�.92j{s!R
���z���UH��ik*���E��e�Ub�0j-AcZ���m(���UEb�5�[QKj���T�"���k��TAc�+EJ�Y�+S��"�)-�A`�����UJ±�6�صe�Q%�b���Z�Ŷ���
9�m+\I����H��U�����"���P�*#R��(�����*��Aj��"�Pb*�ʥ9B���Um�E�f4TbH�"
�������T�#�Q�UUTDTS-��B���Lj,QAq*�	��1km��A�
�#�Tb,EPAU�Tc�E���o����~�5��������o�o�1�㺯{^x'y4��&�E69{���c�?ā}�z}���t�� ��П����cv�& T��3
�㜤*oVx�O���~Ն3�J����S��ђu� �f�,�݇
�e��q�O�~ۍ|�׹��}�zqE �?_��H(o���0�w�06�P���Sl����"���ĕ��5��>٦0��&�wz ��J���&�R
x�����no����>|�<���|��P;�3�B��:�$��Ӛ�u6����*c3</�T����t{�
~a������3_�����T�,���G�D'�����U<ߚ��1���`�Ԙ����<�H
/���>������4]�9������8��i*?��膓��q���
<#��2"G�a��lE���M�ϐ��~9��gʒ�Փd��8�?fI�l���La��t�R
a��ɤ��=��x�Y8ʞ2qϩ[0���Lg��c=d���vŨj�����9˻3~C�F<"���H����.0<ՇU
�ڲbAgY�P��MO��H/��Շb�XbAC���4�8Ɉ��`��
 �����x���> 8�ę�d;���8³��|���aRUT���2Ȱ8�;a�R���a���]�0�4���ڲbi��7��~�T���o�ޛ��ߞi�M0Ă����7���hb,4¦r��H,1��P+�T��|`V|�5a�����6k�h��!Y���Rk��f��~��3����^�f$�ğ%�*AO̜q���|���8�a��bO�sHJ�V>�mE�SALH(z��?2cS�՚H)���@�ۤ����_������+T���P:{M0�
���3���3�J�6jû��S�6r��N��ka�R�*�o�I��>���Ra�J��1����=ط��F�&h��޳P@V�^ٛ����u���U�O;�	i��l.\��2�
�[�Wg�Ϙ���1��V�ޞiУ��_��i��E��S����[���j� ���o�x{�[ϥ��ޤa�O��g�4�P�Ԙ�>d�OKTP�%t��R:ɬ��@��Vm6jû�q��:���}�4�Ƴ�_d��!XcOw~�=w�\�{â�H(��|����,Jì�>IR�oZȳ��`l�ĝB�|�b~-"�aS��Xm ��z��
����
�}<v��/��������d�E�:w�Ө��A�!_>���Y�,�ͤ��O;LE �2y���,��_��M��l1Ǵ�����a�(
,�M���ߵϹ�v����y�o�=����&"���(�=d��9
�Y3�d�1��)�� T��G�LO̝s��a��W�M�y��<d��s$��ӳ�&�N���۽3��{�Z�=�t=���,=V~q ���Y�����I��q�2ns�H;��7��°�0��L|N2c���P���~a�j�G�{�3-��1��c���i��*1���s�y��O5H,�;�'UT��+濧�~�*<�gɴ��e��|�����AM0�1?N}�i ��ŋ=N0�LeI��g޼_}5���W���� D���4�Xo,3�(��w�i �0.���&�^���M'�
��s)t�i�2�_Oِq&8�`D���cg�w�Xq:KN���`�X-P=La�l1?n��J�;?fH
,�嘜E%Hy�0���d�ߖz�I��+=d��)�M�_�
��=s�?g������۟�^��q{'|ºawE*Ag�;�i�����/�:ʆ�#�!̰��`i �6�q�CS��O��a�,1 �É��6���_"��uO�}�+��	��ǽ1ERWY��C�Af0�`��!X|¿�E��R>٬�I�J��YC�
��y� �HW�q�M$<���2!#sכ��=����u���nb�n�`�z?M�u0Z�w��x��nRT�_��� ���3�߶�
\4�\�:P��5x�L���i	���[�lˮ��WE���V���Є��Q��܁�<���ھM�~�$�&�$��?��1g��a�XbN�Y�P��d�Aa�5����1 ������Xy�Y$���4ϙ*Au��'����w�g�kw��?vM�uI����m��`q��$���,>CI8�0���s&�@�cv�ˤ���S�ʪLH,3�,���J�YR�u��^-$-_W�z����쟼.�� y���!Đ�'�RN$����I�5�Ì�d5��|�+}��C�����j��p�}ѹ����@��30��3���RX?Xc0�N��J�:ɟ�p�!�J���VE �����p�a�8��2w)�rC�z`}�+*�X��ܯ����&��
�����t³�Ă����1��
i��ri �=���g��@�8�f�N��Aa��S��bA��y睿��s^}�������/a�r�g{�:�i�5��d��S���}`y���I�+�'�PĂʓ~ͤ� ��,�t�`��ԙhLa߈���j��Q������@`}�>q%H,�hxʟ"��׿d4�{f�w������:�Y�Y1<@��6j��
~dם����4»��I�.�G�,�9S�Z����}{򏇔d{�&2t��J�FN��]$H}�׶qP�Aa��1�gP�M�f$�1�y� �Y��,4Ì+[W���6�P����uw����e��������$w�rM��!Xm�P�6�̰=k6�S��_>�1*Cl8� ��c3����f�6�I���� ���h�I����>�6}�}���}�����g���E ��
�7�jM����P1��c0�Q@��m�$��&3l�'���S>q!�����i��*H1�l�L�1�q;����4���HW��sV��S��┃��:�~��"$��y7|6P߄$R�C��8|��ə��^�}������N��1���pV�F�ī����aU���UP�<���}�s��I�Ag�?��.�q*)�~d��72���La����$�g%@S�$�*q���ɉ�:��Cl?0�=�$m��z����7���纽�I���'�i4�S�{�w���>C���Y6��SF_Y4��ܢ��Rbx�FMo�4�}�/[* ��+8Ρ�>�Y���>f�����]��g�s5��{ץH)���q��~aY���%z�3���P�9��k�H/免k_��Cz�0�6�ܤ�5C�%N���f)=@���8� �A��>�x{μ���,1�Ld�bAf�q6wx�AL�y�����l3�%b�O����AI�W\����h
,��������L/Ԉ��Q����0<"-����1JJ�5�|��_;��%C��N0�i!�`h����4ùOP*Ag�x�'R����2)�N��a�f~�i1���H,5�)��RT��o?w��~���l�eOQI^��1 �f�|�6ì*M��bAg�4~�@QO�+���$�+7�B��{;f�Y?&09ˌ�%zɬ��� #�&��̗��;�y}��(�O�ʅHw3,��C�V�AN�S~�6�P57LՇXcXWL
�W���4����Ϩi��
�����|��z���^{�=�w��ߗ����&��ܤ�|�SL;�UH)�e��R��a�|��T��a����s0�1 �z�g�JŜO���m ��o��W��n���{�gO��Y1E�a���!���,4��5�06Ì+g.5�Y�J���E����h�&�['YyHVa�^�D��>���@0"<��K3�ȯ�'g��=q��J�~�q3��{��o�M3�����0�,�eLE��*AH6��&0��Cԕ ��xeE8ɝ�N T��9�{����U�Ū>��g�j��iڼ4�b[�_�A���
���G%Pj�/0#18ݮ�A˸?}�h9�d�ǂ7����,��57��5���qQ���aP�
؁}|O4�����������$���g���{�*ǵa�̛Ld���ed�9���
z�D�2ì�A��e��:�T��$u�C7��"�R��H)3���1�@�ퟶ�g���$�J��� �;/0�Ɉ
(jo�M;}@�O�Y��&���L+
�2w)��2�T�5��UH)�[1�Ƥ4{�����o�d�H,�y��}5����y�?y��;��g���3��3vJŚ<���AI���\�b�~��L*w�{`c0���>��
²a��Y�4}t���S|�����u�O=;�:�����R��gluH)<̞$�ĜJ�1���8�� SL;�H*�R��IY�N�� D��
���' =}{��8������k��d�a^�`bAep�0�@QLa��2m1�5�aY<ϲB�3��ɴ�j��%~d��`�����'YR�o�'wa�B���y�����{����y�t�����M�(�'׬���
$�a��O�����0��͵?2b�o�)1��CVxɬ�I�c�+4ɾ�,�N��;�w~��y�{�{�x��S���0?5iR��gF�R)�d8�@QI�1�����%b���$>���~�bM�#£����z��?}f�;����Aa��t�00�
����Y���
/���=@��7�=�+v�A@���L�O\I�����!��&�fù��H>�y=��>�}������E>a��1��W4��*J�5d�Y:ʝM��	��ɣvgl�&0�H)<?_Y4�}����^�����Y�!���֭.��ꉠ}�� ir�\��Ϧ;��2��
�JD}+F��{��'�ړq���qqtwճ�.�� ue��_]��pkj�js�e�]�,���y!�Ω��鵑j��D�G/[�)Q�&v�u�����\������`�);/� xz�s�MʸZ~gIv	��(Tp��m�_�_k��T�����y���۬��q���"�/f���Tp����G4��3�ū8��u�է�o&jC����D$k��m�f��j�u��LY�EvF�kQxݾO&LqP�7��ʎ�tvs����3"6����w�����ZLl��VH�R��ȕYA�v:z(�C�5r�z��x�!A�B�g̘G`EL��A���P��b;���<���6�-���O�r�H��MY�s�>�6鳰a	<vkz��S�Ӏ2��&� g�r#�8*g��bȲ��zyR��*���1;����p�E�r#�]"�*Db&D�U�����+��q�kQ���o/��;9�R���D.������=������zL�yZ�|� h6��~�lqZR�������ě��l�,�����5���#c����\`oqu�3�Sd`M��eU*�=;�|����r�z��RU3w�K/���=��Ǐ��aLv����B�xFa76|���CR.�M".'k4Ԝ���V{3��`o���;
f`è>�r�W��f�l�����:��c�Z��nў��GٵWY���,��b<�fEBg��=Ɔ(�Ȁ�Wn����3!�Q��s#`��]��v(�n��v�n]+��CU��5��z�Ou)��>>M}�zP����5���nz=�ޠg�^;\�ڨ�Ft����1��!)L�
A���"�-هb��6+���ޝlp=�:98���[+C�C��al�E@0��&��A�L���e����lܑ2#�b�Pٿi�|�����#L9>�vN��0sB��Ӱ��C��>��"t]�cxK���>}�U�w�x'eZ��	l�H�nH�0��"&�ǮW���$���v&����q��`G!nV��$]k�nn�s��%�4���I����R�u���b�U�����O��by�subn�+
���+Ḝ[���b1M�kUḩ�2+5���Bʈ������&���rq1g��(K<#��P�H�!�5n@p}�d*�8�����{�~�d���-H�2�dQ��~�"�bD�l�ty�j�\
����O`�=92S�	�+�<�V�U��;=�nCF�֯��w�� �zO`���|���^��L��1�2�Zj4i
�qMu��Qw�%-�����~bzE��E#�"EL���p9������������u/���Pݢ�g�1DI��E�9E9^�$YL���E�-���D���_���__k���jا@m��s|;�^��\%L���Gּ�y;�7b�f���6�#)Ь��o��
�O�r�I��j��V� �W�څ˚Xj`1{=Gh��@�v�=��6F��t�t��|:��� ���m@� 2z,E	!ҝ����8��2�QШ9�)H+���H�ʐ��/8���K��������S3"[�q�t���</J�=h�[��i���_'�����6Tm��w*����R_=�<�9�Y�u:"��E��0�V�NW�v�mh�
� xn>ƝZb@��#�����1���FYؘP�:���`�
�tT�T�^�R/��]�ro�ˉ������2�ׄ�#O��� �@\oM�<�b��i����}��:
����r�=q��8Q!�sQ�5���]���#��K�HpE��z'H��m�b�j�:f�>Y`:ͮ������r:����%��HH�-�*��vc��ص%9��">�Y4͌.��Y�k��AQ�L)0+�^��g�j�������&�H�%Vf7�a
�LF([cj�w\��m��t<BLJrb�xs�rm��UҦϢ��ዣ�Y��s�e�����;���� �A�2D�������"뢦�6��(5���܁C9<�|U���� ��.�EG���E}9�,LjPO}�t虠�?q�e�s������V4�bV��k�^�o�'�`:���jwS�..�f�ȭl�p�>=6Č'Z�8�t�[��M���)�;#Ȱ�zo����6����W�P���J�O�P�� _�%D�9�ǔ����/n���MR��u�^�GkZ�ִĉ�ɐcX�9�;C'�*v:(qۥ��������{�U�=�͎���`�`8[fD��v�}z}�nZ;U}��LK�{�DTd��r�h1>�>�\��N�"�qfQ�{!{02�vn�5��C¢�d�Wc`�	 t��8�Z/��ꝯq�(��k���6$Y�EZ�F��������#�g�A\�'y�lo6�!ѓ���(��G���P�5�O/����[v��I.�S`��zue:9��ؐ��z\u���.���8�])�(�c��U[p��5�o��F C;�`�)��Y!�{��U�tAp��fUQ����Q
L9�pX#`��a� ����q(����%�߆������ğ�J������.�"OPtA��@�e�fN%u��In�(����#^���+���K�i����~�rE���I�
oM�(���IQ�4q�l�C��g8V>8\�Y�RRdT�V����2�֍�����l�bں����یAȇt;����Uudt���I���LS�sz�s$JN��;yۈ�{1j��8����	�3�p���"�u��䎱�0.���]�V��3�cB���d͹0U�9���t �Wܭ$����ݴEޔ�m����8m��5H��;v+�ʔ�[��v���;���+�J��PjK�_>�%�@�t#���3�V���Ȣ�*M��=��x���XX��A))Ë��-��sî��Q�;s����;�h�G��G��d�Tu�`�%j������wzD�"jU�)�ڂXNa��u�Nb�V]�JY��+[n��l�a��O�\U�Nx�qp��|��q��Э�z�[����!�׹!K���,���T+�ul�6��T8{Ly-k�MX�Y=���Aڥy%U��r~}�N�e����ٲ���/+w����T7-%3����T�3�_&/��	��&�b��칸��N�4����N�i1���}7:��������Q�g"�c�.���t�[��Yƞ�`�p����K�k+jh�*3����xH�N��-^��3��ǔ�bQ!���.��H�-I�h�-Do���L�s/��Y��6�ծ�_'J�����n����-1N.�֮�W]�����s',�=-�
U�����S�t�D9�b�Y��d�l5��Ǒ
����+Ν�m՜~d�ӻH����K%;���\Ôq��|�g%�a�ݮ�X���Ў���D�Ϸzt�WfZ븪,�M�]�9�J�C�%P�+	puȖ�Y���^��g?.��r��νƼ���ѯrU�&f�2nl�V�|�ɉ
���&��2`��C�;w�$E|�{u�9������C���{�R=5C.>�j�w�T��p�&ef�ubx�b�w����rD+#�`�u��i-�p,�REm�W�/���Dz#H��m�Eb�-�*�)ZT(�Q�mDT��"�(墱1b,U#QJ�,UPDTAV
(�(*���1F+UAQb*�"��1��[j�QQ`���,EX� ��EQQ�1�Lh��
1-("�AE�b���b���(��"����"Ŋ.2�,`�*�eVEEkX�,TQTX
#�m�d��Tb�\J�
�J��E��Q�L���T*�֣D�X�h��S������e�PF1A��-���A"2(�RU�U�Eb���/�^w������_e�*�r)�=�o`6拙�&�uFA�}�S2��W%,u��{+k����u��Q���#�O�t��(��G� �M�������wV��D\hd�	�F#�ˤ�Z@ਫ਼>���Z������}׼Kj<e}�yF��6]O><>��x(�T"#RE�p=N�B--Y��a!;T�"�V��*=>�P�b��.�#��r*Myt�
\GED�u�	 ,�'b�K�g��T��o*�ׯ4}���4�B���B�U���3�yK�>T���aHߨ�*��}NP��9��팊����Uj8�>����� y���L^�X9!�ʫ2$QL����ƪyO-��J�\���C=	
dl�v�b�:,H�NǬ���l�e�ٔ��o������X��d.8:eA뎯1�X ،�Ӻ��w�p���쫏1�*+��VM3C��ϧΆ}^��3/#������߆3�ޚ��Z���b��Yʳ���-�$^�!��ESqsu'Y���t�wi�5%F�����S�T1f�V�,:p��zZtr��DV��v��Y�/�� x��Rm�$G����g`T
:=h�\f܍^�l���POn�H_m_ukQ�נtE��!�0GN�\6li�|�U8�RU���Z�\��D8h�z�ʊ�tƑ>&0ϙ�Ei��YQJ�gF�Gf���/|+��U�9PD�].�9Ok2��*�v��,�)Kn�2zq~cq|����1�s��p(G��d"E�&�;�2�T�簖D�6�Md�"��="��H�l���3>_��Pfݙ�[Pk��s�ms��3�7>&Z�+������}�h��_l4�H�C���^x\Y��{���P�pwI8�S��A��rl�N���Z85���Y�޹��]��4܎�zo�-�S(@�e�C��#o��.�7�S{��[���º�QP=��ǦТβ,I�NF�p�-���(��\s��+��V]���CJ�w�Ў�x3	w���yQz�T�g��,$��<�����s�%��2b�l�G]����Y�Z-a���z��lj��z�:�P^Kx�G�E
x �޼pܦ��9��׶��X�u���y�B��]��x?�����j[������9�5dOV�JFi�;����Q,��١��m�`�C.813�)
:�OD�D��=���	�N�N\��R��yg'��: H'!��!H�[ܹ�D�t��	������O�d+N"�2H~d(�R���$&E���ۤ:���ہ���p�>R���K:OE&���N\M�@�W�$i�3,�OG��`�)��p��uA˛G��f���#��Q�
�&�Q\���V�;�խ�S��0l�
R"���Ж�W��A)������=�	[����RP�s�'ս[��40�&z��\��r�j!����[��ə�z�:����묚g!�]�,������5�*s�V��񁊰�Ϳp�mF-�Ie�������q���]��f4f\�:�2�+�r��o%�4�w�z�G91д�.�T@=��d
���\�8��Y3�=����{��mc	��E�?y�'�L��j�xC�DU����UY��~�ϻ_g�<`�>���ai164H#ap/�m��])l�!	B����J�]m�G�ŋ!�_��>�/?��ȠSª�3��O���O����oD��Ѻ(u]SR��2��^�o/G�hc��/2��Z�K�b��1PqH�vTTlw�@r��8�5�����^!�2n�7����[�h\���ȳѴ6|���E;"��+L�d=�ק��]��\��P�'lԙ�"���WUh~�U
�4�����)'5V�:ɍ��A9�B}�쁶%�BHK�愂�0xe��Z^��;�!�|�B(v+��2�V	��<$t���6|B�=
���j<&2iݖ�ɚ�?I�4#�E��([�F������qLGD��C߳>��`��[}���SA6�)m�<�����y*����g��1� <�P�t��]��hh��jڔ�(�:7����vp%)7���6�}��}eN���W8���m���)h�v�~���[Ӽ�{"���m
{
������M�F`��^1+�[��eۈv�r�i	�6�ψ�B�f�w�fca�>���k�3"&�^�'����"A���$�F|Ԋe���Y!�{��T%�L��v�S��i�� Z������F���g`Fzd>.J D7q�r���g��(Uܡ��B��|_J��B���	�8ό� �cܾt�<���+3����(8�� H��Q�]&�葆�V*n0B��11�Ʊ����^�#�e������Ѡ�E
�]*�����!ɝ��,�V�>��e�^P�����8��8��;���� i�{߈x�׏�F��7���ʘ���9��U��4�t��I�o˯5�s��1�i-��O���[7�3
���2�`G3^͟=ݸ��¬��$��sA�t�������;_�m���s�ZsN����r�⼰l�o,�C�E!�jz���lLî���7���MwYeԹ̼����3��Ѕ�zc`v%ѱ������M������3��D���>��TeW�Ț)�ʪ�{�1�В$���J�[��#jdl���v'��D����z�'`HyUS�IH�-;;��n���^�`L|y��Tʌ0%������B��P곋}���vQ��;�T�k���R�9
�M3C��ϧ�>�bR�����sJj�f5��^x�H�F\	�6�֊�.6��C��|���6�8�JQ�1�T���0� ��jH��;.7�lR�'κԵ��3p��S�75�T_(����iLa�Ϥ26"�TE>�r��$:�����s���D��U�2�.�n��e��f��թ$���m7�x�y�GO��"��	��z����8ո�q�.�
�-tļS6�JXds�Yj�N�Ȉ����'�f��̵^�S�N7�!��v��W
�ѫyvO#v���v��m�7ƅX(Sѯ�K��F�^=�^\��}�~��T׶&����+�UѲި�$�����L�/��W��M�P!���'tNŋ�۽Y2_�  �j�6~�@Q6��I�O7��O������ �,+�q|n��Bd��bA����>P}T���l��2�*ٸ�gq������YX��p���!o�O@��>��r"EL���DƎ��l�I��Њ����Eu�	�UɦЫѬ�9JA�j���˱OFLЫ�!���v����9�5lR��K���g�;��������P���+H�5��F-UC*Y�]s΅�~ʆ�S�O'3���.L�T�b�!GVOG�
64� =����9o:SS���q*K���0@�\1$t��lP��s��ex��M�E�v��[P����iJ��-����	�HLГ�[BEGbaBYZ�&�e��]N�kNx��.�qA%W%2�x�"� uzeq��k>s0�3Ǵ}%��WR�o7���-59T� 
x�nWT�v�m�s�mpe��/��黥#�+�#�|�u��Rdz���YRɻ��bj��9���i`����-Z]�ǐ����@5"���^��o'*���\�T:}�l���lߑO:QH�(���r#d�n��H]����)���.T���#�n�2�$C�4��p=��4��\q㾽lG� �7kga�Ѭ1���0�uz��N.ܽ[��1р��9`L�!�鬚F�*��D�\b��P��<ݺ։Q�L\��U�}�p�����8(�,�6li�C�낧x��+�DC��eO�3A1�LN7�s
�bM�@Y�ϩSg��΅xS50��q(���������K�⺲"���v^3�n���'���ϡ_��.�xC��@�j�2��p%Qg� �((��
�pɼ}[�:q��jF�2�K����lG�ʯ���m];�ЏJ��zK���R��k�D�wT&3�^��k'�@s��ѱ��V�6@�2�x<���]�t�ėomIVV�ϸ�C�]v�sHEh6�R��Pe`�)��S%�ʣ�կ�B���.�͉��6U�n|&��v� 9|�e���⇶��T�:�����䯟6%���3�zM"�BvɃE�!«2*9�ђ��pu�,f���;�8܆0�."l��=HO�|}�6D�B*HR)ת;���9�DGf^M����czC�̍gb��Y+���#�����6HPY�V�s�;&�
�x�߬��ɞ4�/��ji��*U_�W-��'�)�3=D���z���T��]@���E��>�r��SPEs��GbfgwC�����FǨGGD�l�.:�z�á.���3��J{2"��p�qi��CO��b#A��AW!�k���: mMf�*^Y[��� 0�Q����H#L��D#�#&C��ģ!@ɨ�P�t�����˞�8�.��.�t�&��9����P������� ^�b64�p�;,@�ųH�x��.���vo����
�w��xدt��c��[-E�ze��M�;�/��y&-���+�h`�U�oPOoW�����#���;iM�:Z��t���˖��W�Iʍ���R)��p�M����x�Ng>A��}��[>�#��4����L�B-�I��U��f�6���nIrGE)�����)P��q�����T�=1Q;%[����#�Io$(��b�V�zbE7B���"^�M��v2�l������Z��٧��VC&{��PB|@��[7FaP�>�S�"��9����؎��v���>��a��x�~	��7���?���I՝�����-���li�V��C��[cg��.[5�������e��؞�MY���Z�0Κ}.�u�5^5�(OX�����V>��}碚������ziOG�!hɯ�|C�Y���}^���e��5����=�۷|�0u��b(���060"tz�L�͹\*�����y�/9��D5��Rr�@��0���lI0�aÆ�{Hإ�r�&��ߺZ�7X��0i���Ǿ������y�����P��@�N h�Z���޸���/B vu#�:'����݅��4s1i�A����.qA|R��Jw�a4��|�Lo��}F�s)���U�@�Wz!ߛ�$�n�V)'$�	�g^����(�B�3�o�b��,+k�4f��Y��]���Xs!=ݜ>����N�R'r᧠�T��+4��͕ʳ�F%up$�u��3�v�A�č-���}.(z�ޭ�+6ܖTu7�ɦW��N+��"%���)�x]v�o��7�[�ⴖ�yo�=.�V�����M=����s���[eg^�Ҽ��z���轈tnz;S�֞�� ���L J�����Xf���{,)L��j}Y"�-���aOZ�WjH��3��T��앾9���zk�[�W�xD����5����ͬ�]"���'b�v�#gw��"�=���vԳr��Q���I�vS�K�q�."I��S����kڴ[2S�/�.�(^4��? �k��PJu�3V�"�(��:ʤyd������-�W_���ܖ�	��v��؎.�oz�/)�R�!�n�*qN�Uv�������b��vG�F�+�:��t�a���J�ʼ����;��萞~��앱�q��.�ź�֖p�V�=]�4�3Y�6#;��K���k�W�(�(Wg�	��[��H){�{K��j�>ۡu-uH��&���:�ok���9�\��ݴ�U�GU5�������i�Vʒ��(�I%�B+'N�/R����L�Rܩ2��4�)�0��#&�t�?QO�b�j3j�x��Ӟ�07O� �1�o�בn�5��-��+)�y�px��x�$��۩�L�ʹ@���vF�v�.��J麵Et������RS�!,.H�m�j�rģ�,��W�,t��A)N��7����/�S_�	�-.�/�&/��x}�=�v써ý�G ���ul�۲S*��KU���댎мa���`bv�ho�v�:znx9"��o]j��˼�b7C��y�os���u2=����)[������A��p�I-�*�%��@�D@����TX���������DUPD[��E������E��1�T�Ѫ�,QX�R(�Dm��P*AF*$Eb�-F�VJ*���QU��H�E"�+mQ��-��QQ R��X�a�6��J*�2"
���UPX�(�ATXe�KlUr�AA������� �PYUb¤�ԕ��2��l,A��+VE���B���X�����[P��m�*,mm�UA�ˈ��Y�J"��V���*EDE�b�\k����U�,[d��j̸��{�tW���Ǘ��Rnt�@�l*oc�W�u�`gljs�!v$��*=%�zO"�rO��n��6��Z���5�֋�l�QA���$��,�f���R�6�m��sQ�����ό�D�r�hL�x�tn�&aTy�	���{"nr<�TF��P��b="1�s�[�B<��WD�W���I�x�D�c�8��/n��L���fF�"@�٨��*N�ۘEhW����Gzމq���^��r0[�QW�L�T8�q�:�J����ך��ōR*Hq�V`w^���	r�U2}���k�PM���%P�O�b��(2�uUɧ�p�� ����!�3�2�z��#:QQ�p&��Ղ��y;����R���������뻐�K��g���j�]{��h��ߞ��f۹q3;�;o�*�K��Dkz��=C�6��bx��;��z���>�t(oJ�v��o�K��)f~q��7�9ɝ����@���'�:ζ�]����Y�a��aQ�(-�P�F�q�%�d9VxvtH%v%~���Ҭ��^w�`n�DM����#��e�v1���g𯾯���6��~ �f' O�F����←�ˀ0��̍�Ȫ�N�8�VC�!Ic��K� ��[�>ٹ�D���-boZLK䐸16v�	ʇ$(B)BpD@L��`��>�(�=]las���w�3���9�hK�iU�L����D)�^�\hI��ʽV��YI�?i�"����y�h|�O�p�b���\.����cܒ��/�w�i�Q�.��=��8	#�n�)�"�R^*=�h���������|}��M)q������r82�`x%cٮ�;�s�d�>�ă�l�̇���H�9+��D���VM��
�FϺ�z��~�kb��ϔ"�5ST*J"����v�.��W���p\d�_x/�b!v���$?�j3��нǗF<�pC~��j�m]�}׿�� ���&����8#���B�tȹ�fd�����d�,�ԥ�8�$#A���nt� ݡ�2�*�U���6�Vc0�Zs�k|�J'��oz�_W.7Y�|?v��2/��ϖ�_={=y�~cH�p��}�31AFt��I��z��+�T�,e��.�^�#`eb�"���P��Q��@�U}V��9�DY�8�\�nKv��S��?*�O�V*��,e�_����P�E��Q�E�%`*!��0wL��g"�e��O����E;
`�8�c-=��֮������\�d@��0�Y�"�3����{��.�j�޴�צ���=`�q�k��h'� � lˤ"����z���zV�+-������<k��*�H��B�d�&6:�b �(��&a�������{������,�"єt%"���b�[�C���[��9����.�ц�(:t,.4
!3\}�峣�&rJ��Zf�36�8����Ŝ�3��Q�,�/K���vK�k�\�&�I��&.%��Ε\��Ѻ�l.[J`��x��̼�910z�__qq;�kyn(X�� �w�b{j����XV)�F�J�w��!�k�s�l͜�I�%t�į� WϮ�l�Q�>��DK"3��b,�"��D�rٸ�D��乑"	�2�=�7���[���;���=*p��p�"�"��<��펺�U��R3Q|@�X�	���p��ơ>3��[��e�ڻ��)Lfw�b�M�+���PE�&v!�vX�<[4�G��06":&�=���v�b�	���7Y�2-t�td�0�,_�|a3��it�9�F�v�K�o/�3 1@�jH��~�n�#%H��ˏN���] �ǉ��ҡXE�%��t{Y�9�|b�C��r��>���a��uZך_��/Q��"�q+��HO��ٺ3
���Ӕ ��g;����j)��Qcz}>gc`(���8�9Q=�b��>�!ǵ��8m�a���o)w&��~����Q�a�v6.)L���9�2�WGE����~�#�=��lӠ�'ST.��T�~�6�ߟqv�hк��t��6X��]��CU�)]����'�I�
&�3��IR��OpKEp�w�YЪ:��J�&�d^�*B��b�����Mka�:���(�ɺ0Κ��W>�r���������{��|��Ѥ|AB:���B���+���,2�~!顟O�����͘������`v�A�3�H0ߏ�E��H�@���Q��}h�\la��2�S�WQ��,����-ˀa2��~#�0���rH��;ˆ�xwMʳ= ��7��%/T+�*�¨�,�و.
>��y}m��5=�" U���֫�>!�'�e��ʁ�2	b:$nH��&�5�n�:N"4�s���AO��"��	��#���!�T�et��S#+*5�^���4�S"��D�mH��L�����C3�H�l��D�[�;����߫���	�^��EӪQV:i��p���1��NdL�+�'�&(:Vȩ#c�A��>�>Pj�z�l��1���/5�9U�aʞf�Eqm����Y���=.,���5}�BM/p��'�>�l��ΆL�����q�Oef�k�V�xʂ�J�=N��U�k�i)�W� �/z^4�,ny�Q�dl��}��M�{��	��P��xS��㢹)���3�s=="�]+vj��5�~C�)��{C���1DF�dvFD�j���˟�f��E�{:GУ��١�˫��Jj,qP��_��uC#l��ݹ����wa�٭&8�>ؑJF��8մ�T+6z�V�MD۞�]
�DP0݇^�Y0aJ�O���s��xQ�����Y֥W���S�j@�!�#��"`�D�B(I>�[g�g�-���\�u>�"X*6yN�H�rG":�B�'I!2���Z�a�-��\Őow��aټ��>�M�P�)�:���>	��2�4p�!r���ol��G�z~>*�6��M��s-���'�(Q�e���wvcJ{�M��ı>�.T��0-���PS,E�8#T�ܪ˘
_�~�ۛ ��G`ƺ��E�VT�T7�5�;n]��qXNf�T��mH1a�)�&��͘�)�Fᒶ;6�^�/��6�;�Q��_VX��m�:���;/������i4�G������@L�*�8B6N�Cg�l�r:pXU��l�U�&j��H�[>��4x��Cg�+&����V6b%���W<ș;�I(،~�L��aɧ�*�O��8Ej��T8�D��G�ֹ��g�0� �pdt��H����m?��C��׽?
����н����E�1�.�3dl&f,>�^��|E����N�~��%�\�K\*��B�(X��N}��V�)�vR��9��Qr�#�x�C���~U���U���\�j��S��6�eͺo\�3�X���%�t8A�bH�j�P����ȯYq�2|���y�҂�=)mcu]��M�1!9zf2�� l�	�&!$8U�2*9�&�ٵ�[~����}�՘�.Z��������]i>]V���c@Z�Mf�S���㵙!m�+e�g)��t�+��5��4�(d�'��U��]��[6zf���]&�Tp5h�=����;��(�P�)��E���8�s���V�ˈ���Y/v!�_�U\��~��Ͽk��R`�����)}ᶠ|O�������7."�X9J�&��b���^���T��^Dt\.#��R"`��t����}�Qq�d�0C��:/Ν�Bf���6�a�	*�w�8��#����i�;S>,�zaGD�l��q�f6×��n�(��*7ɩ)�3"/ԤD�1fA"��&��o��]�����A�M�c8��S�Ap�4^��aЮC�@�ջ�B�|��z���zz)"��'K� �5	�Ԣ��}մAȋ|E.��\�<0�z��E: ϭ�f��!DvX�#�eDG�t��Q��s�r�܄�(zV�&�32�E�>�!Č4����L�B-a&F(ܭ�2�D�*D@a��H��甏��y�W����<i��Kc�<�f���wm��+�ܡ���=�ڬuk�7#2;)s����a��D	uD����!vv���[:�r��C�/�Y�w
-�<4IyX�Y�wѭ�*[[��R���������-o+��"|Ԋ��B���Uzb���\���
5��������^zXɸ�"��4��Y���`B|`f͊3
��j��:�^�%ا�zCCh��>A^R��vX(�e��]"���������|B��FV�C�,��^��ҡ#aL�����v'��Kٶάy��K*ʭ�M("\�G��a@ؖ�
gMǊ�u�!q��P{/q��8�����'Ŋ�� E�˙
\�z����B��f�!�3���]g��J2��I�7��;�x)����L�Ok:M:�Hq��{驳�gܟ����:������!mLѝ�xk��=O&��t�������l�!�(@��
�	��T�=��|�s�-��[�"�r��T�;w݉i�)w2��X����6fMOt�s��۝x:�uwmS�������9s�=�ʕg���7�=Nx.�V�`q��]Lc�����iX�=Y�kI��^������е�Ee�����������A��$k0؝L�s��[�Y�]�U7������0l�h�I�m����%<�'�}\ٵ�Zs�X�n��ȻSNTйr2�zv7ms���[X�l�퉟h��]`J"�]\��H�.�nn��M���Q��=�C�X�F�7�@ڌ��.�R﷟B��8.��	�DC":`*X�Je�4�G5������}Y�سҟOg�c}K&�s��Mu�Ic�H�0�Ҩn�e��{s��xJ$by�S����[���*�vg�����
�e!���w�ɳ�I�[4�;�3BO/kvW��.6�zU�?�s�٨=E�Ej]Ni����K�[�8���I|��1��=������?c��RI8f�^� b�Æ_y@�!�L�I��.���� F�=��EʸkSu��,�'9��P�z�ޣ���RY��9��q]QՏ�1�;�D�<���jWFC��S����sp��C�����e��(�t@�]3Vi�iYF�r�:o�wH}�a��BXQ�ջ�`]�.G��-L���sϱ����x���V�2�]���a6����X�H���1�`�r��]��n�Al�u7�����>H���#}N�P�囫9���L.�s����i����Jޡ.25�����8���\���0�՗k�;��fX;�!���]bi]|�d՘n��W -���BRSF
ۄ8./_r����({^��k��b�����7sE�/��҆�h���ʡ�v]�� c�!��	ws�	Gka��GZ(���$wO9�x�x�W7wZ�Cj+��J����;�Ū��d۔H��g�i�`<��xe:���>��qe�M@�~^�P9�TOOEz��4���8�dUխ���c^�;>����^��	�7����k��zņݸ��z�,�Q���jK-�M�9���e�7r�@�/6wYd���^�3q��rN�3;$u)]zV��y�}�w=�Ip��n��(�|p�5�u��Г���Or��Y�A������4�c�s �.�!�;��J2.�v�Sz��:�7�%
;o�������1sL�CW��t�!�O��q
��-�vK�c��mF&it�������횼2֨ˉm��[�>[p�.�r�#c2`����e�%W��a�&��^u|��-1*޻u1�]��I�wЦm*����\	���qP��u���[��b�5C��X�)T�r�~���3��9;��ߞ�Au�5(㜉�C�����Z�74v����S�&d���U�6P�z��+l�]t�z��y�ui)f��V��[�]�-�;}wАi���R!���z�>��I/6�]3������j��T�[�i-j[Jѥm�1EQ`�h�m(*�*Ŗ؈�QAb�R[lE�*�QE�
��"X1QJ�`�EV�+q������*,F�UGM�(�EAb��1��&���2��P��a�!��1*.���QDEYUb�E�Z:����DU�+
�PEdQ�)mDY�Aq�I�+Fc+X#V",bkV`Ŋ" �"(
�������UU�����DQ`�e��"���c���1XV�J1`��CDF+*�`�(*�Q`�Qhh��QƦ�TQ`��TUA�AEW-@TEUYm����QE"������y������??vm�B]wA|�ǂSl�a�ܒ9��c8��݂�c��P����
H+}@���x�7	�	�r�ogI�~G�B�J?Om��on�*>K�܁m�����T�}�y�ߒ������MWe&�c$,�=%[�F��r��F{�f�
(nb���~�4;�CzB��N�N9�$3��*���t^�n!i���8��T�t�L��n�eV��]IlKu���A��|��B4�C�����c�fks/7T�K���_?z�/�L3��]:;M�MH	�K��ƨΥ�|���Vy��V}aH][Vmݾ���V:���<	,�V���XP����L��#:��ȼ'�+�V��po/Y�يR��r���#��@Ƨ�)�\������B�޽�"[n�r����ފ�h��2��ɱ��殆�M���J���ǎ��eѭ���ȏoQ�s!v�6�!���V��S�pQ1�e=J��:�Lr��m.�/.����u�<J��9lD|
��ч�{7�����qo^�k�z	��D����8��6S5R�!�s�"�/a��D��yK;r�SUe�*�GsӼٗ�rJ5@Y��cc�v�bi�j{%����a��~c%5����Mٓ��\���r���Kf�H�s�\��uy
��b}æc:"`�Y�sJ���4���I�%��[�Ԫ%Ec����׷M�A�>���3�*\+k}I���9ݑx�Z�O��=�M���p������z��U�jx�Y�z��x��}�H�J�/�|��o5q��y���E<�슾{���apl-P�(��0��!oy�oH �h"/�G�8��±�=�{by�B�6y#��K���%<��=�c������*�[I�T�:��+%:�S����'+�{8)���E-3s����VNO-�n:�}����i���W��z��{����8#~\����r##\�譮���O�Ԍ�N���iBx25�9��˾���1�|�D�L;n��E��jw%�;9������\��[1!8ю��u�Y�Weݾ2�\��#����M�O9H�#U��X�F̷�x^mP��n;��n�i�y��;Nx��yp�HI�f6aG=��e�G$&9.rj�\�qX�ׯ�U���Բ�.�t�/�5-nke�6�~>��6�"b&FX�.~����|<���3�7#��Ol�Ҹ��l��x�;ݭS~�f��9t�Eűi�c!Sާ���)����3j���N.�5[�6�2y��!��źk�l�sp}�"��^M]�j�xI�E�9��A��O}/���ࣺrR��.qb�Τfb��Mg$g+	��nƹ]��.������tv؜#�.������e����(��3�B�.�B�p�sӦsd9]q�0��9u}�٫L;���J�l�~���;l +]r��q�7����ei�}�4��x��x�=ƺ�J��n�����1�+]Z�OfAnQbW(�yFp�ݙ&�W�a�k��! �:���ox��t�b�F��$�b0��Xg�8ٚ�3m��88��|�(�J�=�x��0,�㌄�x-��j��M9SB��Y��o����Uz��+q��e5y����y�Mٱ5�ʰ���X�Wո{<_�Sv�C
�/�c�G}��60������wIH�c�^��k��kX�ݫ�z\��$b.6��]n�ʓ�L��&={;J>�,���5���3�(����//v��WV�lQ-@�װ5�j�k;S�����5�g�.<<F���Iv����H�:��گ���I�o����w92)��BE�x���C�����y-�]�MDin���y4��؍sy���d�c�7X�w���wRZ�ӷ�PU�VO	���y!����~��a�#ѹ�̷�O����c(���K�������{�MM~O/���I2�l/ ��^��_�-�],�xi<�$�<ַ�Z�^y�F�lϟ���X�dڳ� n:�$��.T�ֺ��v�Ӗ�d��uHsr������kB�1��)������ɣpq\Mn�W��2�|���#o��@h����A������u�qV��1�;�g�N$#�o��lج�>u�Fٜ���f�P<4L^�{�С~.��<j]�ǃ�;��2e5 M<��5��kX�Z��[�N�����\���ڶ��p]1鋒�%5PZ�f�*	Ǭ�ͽ	d�2+��U�Rۊ��r��q��6�����Y]�������K<�·��ɡr��-F.��h��,�p�]O�B��b��%p�Kc�WFt����Q���}\�sf"F���V�����<i���9��/;�s�a����lWP�.|rQ�t�E>X��s��sE�x��/�(L:V�5�mhH-/��WnU��􆟝��'���/rŷ͙�d!� �$�S��L���5���;�A\��Ή��A��H�Y���;�0��>�Uzܱ\��4܋*Ej�\��hE®;#��!LcR�����V4d'��q��BeH}���V�6G-�Mm����8��W[��i�S!�Ȏ�ԕm����v�۩�Lϵ�먫�B�+T4FR�*.U�'q�J�@A��>�� ��絝 ʗ˞��吭H��f;aX+~��9��v�F�ϡ�~(��⭫��d�Z��
&.�ӹ�)��9b�[�9"�Z/d��D.�m��-ɷ�od�l����ը��NEJ�;E�X}Z����z�=S�84��P�/�(�yD����w�M�K�BD�9Դ�hFm�co�Ʊ��d.VjwvB�ٻ����sZ��*3i�P�X��nr8�͔�C��"!��Cr�3\.�S�%�9�8�+e�^;�'���s���+R��y���]4�u�m+��O.����F�2�hՀ�Bni�b�r'�5��X�O2+�����&k�:�e`�}�9��Cx�C���eC�ob��~>�Ha_D�p�'a��0��~ypg�1(��'�8��Y��BK�~˪� סb���3��e�^�+L�)������9iK\*��Œ�)�ި]����9�����y���5�$ZSy��v�볶��U�]�[<��oӬ���W�{˛_3�A���h,�9�v���n����I�zҨ�«`dS��:�w�-T�t\s�ϸo�e�ާ�$����3�ޗ�ܾ��]��u$�|!A�����q�6�C�귴��5Nqk[Ք�v��~�Y��1���ܹ������W�du=E��NE	I_[/oz����z����w[+^̂چ,.PbgDQu�6�^�+��(���!����3�}�<�˹�Y����F�c	�>8����VQ���/@d*��[ϳ�2���6��ܰ{��2�2���d������r��:�4W�zm�2	�W���=�^f�iG��vy1�|�L�P�3�"mR���ѣ��u5�B�ݝ��6�2�'�w���$�G�B��z\�x&�nԊr��f�66�'ٝR�[�*z��d��Xߠ�+s˫��p8}<�%�8��C��s��'FV-�b��5&����u���nh�um	�rQ�ui�uѡ[�׼��6`e�#/��+���s��ݥJ郍�*k�(xxp|��[�Cs��A��GVȾ�O*�\oj��ql^)M���r��V3@J40�zz7R�*��^��%W��}��٠�C�c!���)�U"j�����W���M�OgI�a��0_e�f��]-��oi\���7�\�n]y�F�gt��{r�n�
o/^�呝���v��rIԺ�]\������w�T�n�Ǐ�av�Y��}C��ί;�+9�� 5)�ĩY7���s�v�,҉�J%���{]p��i���6GV�+/xX��.y�I�J�񝀹�#5��u������e-���UtoG4#~���єԇ\)�����d"7&�w:�݊	j!�P<8���M�����yyI��%��g'ncz�&8Ɯ!^�}^,�[9(UV�}sV�{��5��oԪ�ypSW}b�����ݫ·�
Lcɧ.h\�^҄���Գ�X퉚�s&�u:�w�9/<޵sn}wsM:�66�2�*��,n��dl�"�w�f���t�|.^V4'�uST��ȒVn=k+�fR��)W�J�p�ɥ�^��8t��F��~��O�!ҡ����r��Ϲ������ԝ,��=���t�~w\q�,�t���>��`�D��Uق/j^��i,��EX7�"z� ]�"�s��L�*�>'s^��G��ギ!0^�;K8aN�,�j�D���xL3q�/�R��ҎؔN6_lF�Hq��Y4�_(x��:]��9&,p���Y��ź0�6zxF������"�O�y]�1/��p��Ӻ��>����"n��*�:8�5�k��(�OFI�i��ǃ�2�Ux;���v���j���� �G�@	^�1id3�l��֖Q��ҵ��j�B���U6���Ff��Xxb��qTׄmD���@t�G�3-�����[��9s�D��gEw��rE]wOe$�D�Yu"��:-�n���s�ݓ5�+py�=�)�����T����^��=��Ѿ9Q��C���{O��o��tO�pj��F���4�p ��!76VU��6�����E��O)l����+P�o)�Bz
���v��Bݧ9ú�I�0K�\���������jfp��)����o�a�2fk&c�_cRQS�a=�mM�8��g���.x����%� w/�to�����(ܐ���{����֚M*���kyPn��-�U;��+c�ޜ0um;B=X�U��1#�Ja+Y�چF~Ti=�)ax5�u���N�YK��tw�#<_{Yy ~��Y�$5@����΍�2�9B��G�X7�0%�G9��6��g_�uZ�Ӕ
�J��g,P�˧[�쥖'�fl�LΆ��1* �]q�٠��4��V�|�M+�D���ˋ�HǶcM�����jx���Mt�.z��&�߄Cۏ�r�@��Q�7GzcC\�ꝁJ۷/;�H���$��6�dC���v8Z�X��\�z0�;0�G�&�/r�3�Gg,J���w<�� �m
�>�vy^�I�jR� eoE�["ћ�ɡ�%���x���(���]�(J-�����E/(%O�L�$�>lL�'%�v_�vj�X���5�ԓ9lۦ�24j���#=f%��/�A��܆U�ք�YA��-kH���0����N9#QţL��ڥV�䗧��89;�~7�}���{U,"�"���DO[EL����0���j",F��%J�,�AT�Ŋ�`����d�TƱYՕ,PQ���EX
����A`�*�XjثUUU�EU��Q��V�`#$*�R��X(Lea��Eb*EUQAD`�ACD����(�(�(��!E`��".�X
����������FЬYiD���1*m���R���kZ�,E�KF�QZ�m("H�
F*ET�5Y"�������E�*�U��Uh�2�0�?|�!��q���u���Pn{��;��[�˹.�8�$�(�+�:�2��W��=�nm�3+�W�nNs;?
Yig�8b���Zʔ� ���O;����O"��bKR�ߑǬD5�2�g��.Vi��� �zĂ�l��.kU�Z���p�b�78���c�B&����~PQ������}����O����X]�U�p��ײy�T�O���E3�ޟ7��Kg��3�Ot˧��W+=^y�q�׋tS�VL��7�]&���җ#�9%CE�C�ӥDf_	X���V!�ƚ�R�N��`.Q �tW;y|{��s��S����Tܬގ'X�FpEN�J��}zۈ�4&r�j�2��ۭ(pw�c:�p*;n���q>���N��k<��yn�E�^��ݨJ�<�N,}̎��ە����9�R<EQi��v��(NmN�(��4�{¥����jv��d0u�ΩS:�o�қL�	��-�5UYI����e6ڛ����[�{�Vt�LH[�1H7u��UJ���{P������mA���r����8񑮊�5H9(����-Q{}z��V��U|��J*�\- ^��tN��[bgp����c��3�ć�_2��ʐ��wa����&H.�����:�2���N;��x�{�p��.��s��:��USU
ͼ�{�����~Zy�~���(�|�v��*8v�4����ޚ}�Q}�p�_k�}uqڜ$�����y$˸PB��rw7���O�����֑ݳ�����׶ۤ���2���l��f)Cڪ��
�⳶#�v�#2�p<��tef󶟆�&]�F|k���"�n�V�9ն?l����C���"$9+/MX5g���ם���I"�nh���˸���(�[9���V)�=E�Zr(JY�lר�$�EOb�潯B0ސ�E>�jS��a!he�:��V�-hN!C:�X��H!p4��sa���2�[��6u;�:�m� �⊱���6-��o��@�Ѳܽj��_N�C-w3uK/�4�8�o�k�Y��t]Z��q�VBM����8|����o�/��v�a���ߋ�>n�/h�`C�<퓵v���,�Ur)��*�m�Y�Cg��LW9��os�C��"���#3���{M��.�psz˖m���[�.N���-2�W�����ggԶ}}Ѱ[Ƚ���-i@伂�2I�3��Q���Z{1�j�%AF6���t[A��}V͌��cy!sT��e����܍�Vչ�AVq!p/�Re]����onP�U�y��؍݇����*�I�V�kӼ�H��F\��A�%����Ů�Od��m�V���ql�\e0,d4.����Lkǆ{7y�
������>ɵʞ�I��c�@�⯪�9Γk�8W �L�Om	iW��j�m))� �bv7g{�qϱ��}`�#6T�=k�R#il�#����-ټ�ͩ�H��9𾓅��C�Me�\QJor:��[x�k�\�SG�rdl�G#o��CG�m�vJݼ%����vE[�Ϩ=�\8��HCb����ns�y�ũm7Ь��1�.��\��"�l"�ގ{��!�"r��H"�o�NTйn�BV:�-I�]Z�Yod�~���#���/3�t���_V��G�uW��$�)-�./�](iԈb��WS�h��Db��+�B�M��l�;�Z�[�u}�	��2v��K/+f�>ϗIq�}
��z�rF"�0�ҹ�wV)7����ަe�]�*�V*�C;9������wT��5�r򱡉�[C��5l�-�n�R�3��KQe2�|�����4�7�����=�LLZ�RnZ1���%	���mGn��W�Ɩ�p�����ԥ��o:�w�'�S��c�P)��dkyrq�7q��r���5:�i�\�t�5�YdnF12,���j��G6���9�Cϼ�3��Z����#��C�5�Iݩ� >«/#���|��E�<���C���������g�o���%�����n�-7B����^�{G�W%ݎ�t58�6����쑕�(_vM���i��h �-=�yT�zb�kC�m;���,:Ss�a�*|��+_'m��	S��\�R�L7���ۇ덒KOr0`�XO%$�1�Ry�1mX[�
_Zr4J�8�3;�+;b���k�R��lN�׾?P�.�fX�ą�$Q2w�p��6㗞�|"�g��^�[�$kU��P+Q/��,>l;��j��NM�m֔$p�=y�����͸���'�㱪�����Smw���}VT��354�O��	�M.0�ж�{��z��.�A��.;�������}���k�+��� �{�q�w��.k�����&৛���x���J|f��f�=�����|kd�����Ic��^GV�ʣ��m5����6��Զ�����������@pt��-9�wN��\���w�Y9!Y�M�7����%���z���ؑ��B)y|�+^p�:�Ewoqಚ)�:�lj��[�r���l���$���P��tz��9��X0`�i�]�"������� �6���Ӝ$��ZWTlYs���w�ܟP���e�~����U�Q����ͨ��mJ���ڞ~�����}|�{>�I2^����u5����/[Kf���m��{�m�III�!���ĸ��`��c:��d�}�4��WJͥ���Zs�f+Xj�,J�b9��!��|��24R��Sْ�x�טgj	��u�{�A༷�|R�8�t���F�2($��̸�U;9҇i(���3��M<A�ӊ.�5�p��#kg9Em�Z�U��\5�ݮ�e���)kU����f�j��o�vL;�N�K<��5aU�����f�G���lvjْ�jK�w�yϬk�8���K�9j6U�>�����,݀�?a��s5��3ibt�����ov@��s䐽��E�H9��t��L�m��f7� 2���4���;���}IsL�*�(��rp�/\�R�'[�]�ݭ�m��,r�o*����QB�[B}�稌�wSR��׺�7����FcG
{>���w���yt=٪)�u�>K� 1�ڲ�=�l�=;W�bdઑ��[%<)��)��O֦�Z(� �;�(=o�Wx��ϟ$ribx���Og�\u>�`���/^m(�/����U�VOlG��y��x�o�zql[r�y2�1^���N��_�����B����/`Y;��m��/_~G�:A]$�Fk.�=k�A��,MI����oq�VH|����}ML�|)�u�"��ԧ5^z!���Zt�������	���1U6W]��+�c�=v ۛx��*>��k�]�	Z���פ�C�|9#��7�Ru�?�7����u��;l@�5�.�p�.V�s&�r��ڊLm�|�����ardT�}Î�@T��S�pbE�c�mj��cGL�Iv�/��Ĵ�B48��q��8�xN�=���,]Ǖe:�:}���wn���;c��=�"&��*s�-֔$p����U���b7�2��LҪ���B��nD7�݇����ެ�%��-QY/��֎{��=��S�a��Ľ�z<#qB�)b=�k%�;;3����/n����O>NOi�]�zG��(;�j�S5("��g9��8}I�#��ei9��D��Z9b���8�Z��]Ӊ?N�lIM�Y跐�tO�"{��W���-t�Og
8X���9�;���$Ww)ύ�lƑf(����;D6�hs�.m9�֌MV+�%�Kh:<�Fe�Βds+��軘�v2�(.,����A¯.gEYW9T�9˼ڊA�[Q�Ew\+�R/z.�j
wZV�j����d>}��O��W;���x��W+�{���]���n��PW��m�q�;�/XG��8�M��Q�Z���׳m���/���OlH�E\�Fn=k&$]0�b�WZ�甹iȩJ%szn�rz��m'��u��.z�Z�6�Ab@\�acµ����hB�02�6�g�IPAʬ���v_+�n*vm�V�y�,�Mp\mi������m��"Y^��n�%p+:{�������5sv���R]����nfb�O9E[�LPB7������&F��1F{�O	�]jaԳ��7�O��Ǧ�}hI���=��X��.�.��[�)΀�Hau�F��/`i��h���vz嚁0m�ޝܬ���Y��J��Ui+	��2�ӛ��[��{k�}�.�ͻ�k7���.W2�7��Miԥ��;�pɇe��ټn�=.볛�\�CMmj�;3.��Ǚ�N�줞^�!'<T�	n_|9����x�WY�����O�h�]F�:{��,rx�!λ������=�*͠��~�V[�.Hn,��Z&�������#�9;4����+��joL��W�xA뺏s�Tҫ	��� 4O��.�VoYn�ۤ�/��#5e���fu�Gp�	3�=�ec^ĽM��Yx� �n[��:��}��9�>�K��:^��b+�{|����]I���j=���#e��ק+��M���-B��D�l�7~3H��?%I�Avp=�@���Qt;n�X)����<z����*�L�Epł���[����w-@��W�B�R�]�>��*�u���]w�6v��̉����&c�*�=�C͞��Վ�T�з�V7�w�	�땱V<���K�D	V�M켻�aS'eZ��r�vT�(rR����b��:���l�\t��'�Upi�
�^T�D� ^nh�V�9[�r�T��Ax��)�-�ʻ�^15 3��Щ�����y�s���Z�Pf\tH�;��F=/��h�x`�\ܾnp!�k�;�0��]w[�n��MS�iZ���ϕpo��Yu�ٗ���O�7�Y�^����BV7�O��ʳz*�DZ���25cPܽa�R�\9�V����u���bZ�����>��袔2Ρ�h\�d;�\��݌<�j��n�1w8#��+�z�o�:�V��L��U6�׫/x4Ua؀�<��!��
�tfХ���\�4�3>��C2T���%k�����$+j��yY,�ڵ���[b�V)�h��~4)��C���c�盞���p�=�7�mY!]��oV�h�.M:�B=e�1��=U?syv�Y�ae�:�����Q�3�m?�g�r��:�;�1:�kz�W�U�I�p�JU2ebź2[�L��6һ�(��Q�9\�;P�'I2��=��֖b:lƠ6��ar�2��VZV�T��Q�Ab�l�FZ�#UZ*�%������(��Db�#e2��P��Ah�((�
�Db����F�h��F����Uk*cEAUj��DX���ڨ�(��Z�kEQ---`)Qb1V��U�lı��-��KK*U�
���E�L�XX����"�jR��E�"�T�1�*�+*Z�X����4����,+Z*�mb��h*bUk`���DUT�fU�kij�%E���&Z[�*(�R�*�*V$Ĩ��-�kU��EX�m�%mR�mKZT�R�۔�h�R�[QZ�q0R��R��-�J���6�-���}Ͽ_�_��W�d��3� -��0&�ʃ�r�o��*��Ȧ,��m��f��R�"���Dj�:þ�Zc1����S��Vc)�u�����j[HT�x��x�RR��7�F=��C���,�\N7EV����H���NK��hp���u�C�C}`s�b��6�7u�i���]gY�/N��ə�O��ʞ�����y���M��o��v׈����u���=#�aQI)�L�q�o��캷��8�U��(q�c$xi�y��W��#��.��?r���6��&]�\W��0Ub6�bAu��LF�l���OuM�M쎵�1Ӵ��M��W��\DM]�`S��"3g�R+'�d�N[��%��'G4sB�;���~#!�
sz{}ڳ�{�b+��V-�K����k.ќE��J&U��{���/���Gg�y�yiӢ{`�Č��KB�$�|8�zM�d���uo0o]Y̓�8���{u%��)�ރ���M;2$#��h
��W^�9n��T>�M����cgE1[�<�@�T����	�L����Fζ^H�6㧹�|�{��3�<Ƃ�-c��ܮ�e��N(J��yV8�o-<)<y4��\�^۔8X����,]s�gU(t��I��k��sv�S�C.���3����T��Ik��A�"ʨ�3_�eE����������f�t�)��Sʳ��pҎ�+�J��H��{ SC+G+"H,,�i_�k���x}YC�}b{t�J>7-X����tjn;�j������v�<�;�2���6���;�,�fd�y������쾗[�^���Ԡ?uMa���5S*���P߲�u�jh׭sk
�2��e���hF�a9%^]���B��p"�t��Z�CJQOQ��{ɉk}pc��sR�Uf�#�B8.��9�l6���P�'���A���2��v�%��M�T��Be�w'�=�K��LH��O�s��k���S+�ۮB�v^�u��S}-v�W��gY]F�9s⭤��[�y�b[Y��x�p�VH��y�p�3P���NvL+���ȫ�U	�	�)bk�"�8q���)����y��D�B�x��}p�\��Jq(uUp��y�\�$�)��J*n�eX��F1���a<{�rh!vv���F�:�6iʜ�Ku�(O�!����]]�;Jo�� �:�����܁I���$e6.'cB����C��p��Y�zM�l��ڌ�o��0����� /�.!��I���b�㡪/�TSD�A��X4���iW��v��z�m�t�Z�^�?���׆�s=��ء��B:��7_=�H9Aʃ��<ϖ���6���mh�-I�K��S���0t}6�d�rQ���w�>�x���Uk��*WT�ek���R��7��uy�n͊J�dZ��V�9��D����}�x\ro�;'2"��Ǎ.�=V��˛�$h|�wr־��|��r�H^����/a���O�RSgkJ�
B�T�R������S�Tu;�zA6K/��t��转�p�t�NL�V��x��n��PW����y��=.b��Ӛ�=�'z��N^�^�oE�DP	�!���T��۶]^�L�#q���{ҝz�����/JQ�أ}�~����'|.z�J�����b�@�Aˌ�\�*h�Ԏ��چ�jc����
:V��d�v�j��:���{���OJ�w�_#�0�<�mIŶoh���;i,ɲ����{�
��Y�GI텀�ܕ���|u����i�V!���LY)�sW00H\4�ܸ.6���fvM6���q�u������J萘|9;��D�V6۩��V��v"�m�|�WOf��NH�\8X�̄����Ѝ"u��s ����V�7=]'oa�]/��q��uџ-Z'��D){V�\�e��w�ɦ�QB��^j�jt�z�����9�Y��F�B��$f%����ϩ�"�ƛ�g�N���^���
]<���o�����fJ<x=>����j��eV�/N�8>T;h��'�ix3*j��Yׅ���2vm�[v�a�ô�8�2A᭞w�mV�v�z	�n��p�8d�}@X�v�{wP��&�(�j����:#U}�E��mw5��=�fa;&�y�q�qM��R����w�����gκ�<%S7�p�v��ռ��Kᚧ��}r��{Y��Pͩ	&]��!yD�6�;��i�~!�W�RsR��M��m�Nң]�j�f�sQ��3a��3i�T%eu�;KjC�1\��f�&mK֪E- ��t��ȆxSUiӨ�]�E��+��Lj8_r���n�@T9D�y�kd9Q{��Yl`��N�L652ӄ�=8��ʺ�f�2���kaYb��m:
�X��C8��N�5:b\��{�"�����x�L�ʵ��N��UN��Q
b,J�#�O�l�]��snn�Yop�r����m�Tvð������!ڣ>n6}�T�ʋYM�.�1:	�@���7�#wjs�C�f }~KS�\��N/�K�',��P5]u�Qe#x	5��M�o�wOy�����6.i�e�j��&��Fq����}aZH����Αڻcb/��|����Q�P_
U�fPKga��;�GL��ݜ��s�O�W�O��{=��t̠��vU0�L�gR�/��=%�潟r�^X�Yq��au6�Y�b�s̆��|�!5��E���C֫Ⱦ5万�t�zJ�T��=�FϪ�!Ɠ93�ΎyO��n����2��qGCa!�l����X�	�^�w�?p(�z<^=M�V!���,��]'�cz\����7+`v�M�ΧX�;]C%����#�^W��N��6mC���J{^�͡�h��5ɑ^�8u�78,���9�����a��2]`r�v̗��ɝ�⇚z���u-M���7$n�$v	tdI5t�&�MMi�9s�;5c��^N��6ٙ�A��:X�r��1���e������y��C���X{���ѥ�0Y�Ꮚ&ʼ����Z��v�|�3$+�=�%	y�+`;�f�6V��	X���Q˛�j"0�Ω�zvbjq�"�)�ލ(O�j�5���?_��ϲ`GܮB� ��3��f5sy"��76U���f++K���1���F��=S�e)�"�h̡ݯ���ܨeJzg�F�S������{��\��Z�c�2.>��t�<��:x���D����l�)�6S씆�i���ϼ/�������t�ٽN(�}�J�2��9�vD�jR����=�p�ږQX��_#~uy_sWP��wNߓFE����Z��{!��������{�G�s�^|ֽc�ݫ.��4����s[�\ߴ%`�s���cָ������,$\E�x�w�#Y��c��,2�Ll��Z��	V���8_��=Nׇ\Ρ�bc[3�I£����������-V]%�(OO���r�VV��L7!̪~������h6谣<��cl�ݬ���T�0̥���;ܟ9�R����^Ͷ�֕A6_��gI�����O���NL�)v�=�µɧ��/�9�Hj�5J_N��LGC��e@ƍC\,�"�=�m\�{�3;��ykFPZ���p�7�p�MRU��C� W6�B�������x":qQ��1� V�sNr�o]&�^�y�'�9ꬡ�5��9����dp[m�Յ�#5EbӘ�}
���١��Sb�L�MH]1!lL�8��'�����=HQ�bz�UY�l�#h��=<dk��xl(�1vgZ���S��A��brg���B���zj�)�P�������]^��8HN��X+�!T�J��͙]�x����|�myS��-t��嫝[A�Cz���l�~{-=��/%u(_bg���E�:����a	����IEM��;Kb�h��ٲ��ϩ�6���Z����V]���j.�����Hʱ{^�Y��!��Lj�I�m$841M!���p	�&}^"���4?X�Mh��v�h��c���٥��%_K^>�l����؆���
�f�bT��w�I��Ys�Ͼ��j|�eߡqzDN)eƋ���性��r[�ޟT����?'����q�ۗ}�z+s_����7\�:+5x���Q��sOS���c*���q���c{���$p΁��K�1����n�uS��1���.WN����E�M�, ����S�cX���E��ن8612�ӉA�:q@��ѷ/zh�`������ Ŵ�3v�y�
)���l5ul��GG`�=*�>�o!ބ)��L��F�Gf�)�(�ui��rˉR�֩����Fr]��n.���i�������]c�w��5�RU�Ge���@Ѭ�\ȯO8�&�T<h�t!�3|^�������mݖ�W��E��s�����&B��v՚����[W
��~�"�5���w�I�ֶ�  �g}{�aF�"��\`Av��0� ��i���L>�ĀO{|c{f�˗/^V���Mn�gf����b`w�t��m���x��[�\��+��\����e����j1�{#�#�ڪ�	ܵ�t�#��ҜmT�b��$�b�tI��1�:�s�8Y} ��|Abd�����b�J�W����ۮuq^vN�s)Ģ{X���kͪ��"�:��~�����1F�@{	��ػ���p��;6O�u��4.�:�_$��:�g/�zf��k(sv",��2�ծپ�Z �|%��>�����4N�A��Zy��NVr������]ɇr<W!G��m�^���
�P	*�m\qC��S�P���Ϝ�	i��4�fE|�W::9[}���kK�Z{A0i�Ѣ�� ����߃PQI�zj�"_6./��9>I�w&j��@oi%W����yK-Q��me��&�{@>OcF��qI�_�\7ƿo�Yf��6�g��E@���o�9�t��{kREw�$ݎ��|F�Z�G$��]��.����ʫt�<���ZY[����,Ns(ҫ�3n��r�B���g�܊�{���s� �m*�]� Fg%�o�u���[�(!��(��J�ٴ��jV��\��n.(˩ۜ�V�|�h��e���KCR���a��;��2��1D1Ƴ*�i䠂�$�B��� m<�oB�R��Wk�CH��Ԝ�jR�^��K(����a�	$�RV�E��G�C6�Rr{��%ZTP#7�&oh ]�=�={*>VuQdc���G�3�\�\w��R�x��lL�I�"���4�7��|�p>��dެ���V�b�o+�-�x�0(ȴ�/���vo�Z��U�IQ�>���h֦�M�}���{3;�qPN�Nv�'90��Ͼ�ѵ��(�[*Q��l�f*ɍ�U�-�ѭ�E��j�ִ��Q�+b����0�"��F�J��j)YZ��,,*hёŭ���Q*[TU�ET(�
V�.YW* �%�[PUAA�[l-���1��3&V��Z���T�E�eeTb(UAd���`��L�bU�
���*��([Kj�P��ĕ*T��(`�*TYX�@�*H��)��I�QQ@�PZ��8(ȥB�����
��,��J5��KeU`�6Ղ!Kb�kl�Er�aH�Q���U��²��Չ+
�'�L ��LU��<�wyr�_mj�5dJVR��f�^�w�r�:i�Rj���rI�vn\�-竳�n	|�~V�٬T�C��k0��e��Q�bJvr�k��~Ll�F�v��SE�r�5A���Kݾy�����1 ��2�]�4��e��
(Xʛ���i>Z����mQYF.9�^6���P�C+C:W�E,3��O��#��t�J/���5���~Ù�@����ԭ'<���j&x��&1;S�We:|=.�vs-w��������jY]A��΢�;͗C�u��vo�N�~�`�R�8���ҫq=iC�{��j�ui8�mDH��X(ҿz��yf�ȇ���f�.*X��n�)�ƏiV�`�N�{�(�D��Ç�������^��}����kQ�mN@h���^���M�i�<�f����T��6��5��od۷��IN�����'�$ѣ|�v 7[/,m\��3���d�WK��\p�k�K�$������Y�
��Q����с����y3L�e-�}���09����bH/R��sMdĸː��ų��|[��+� �Çu0�X�1���ۼ���F,���2V^�ِ_L6%rd��<sjYYU�}|؎�����ރ7]M����c^�嵳yJsmZH�qE���}Ӳ"j}��)���B4}��se�[Cru���s�۷6ɭ�+3;�xj�f�{Ć҈0�
�\T_n�7b�a��FSFiM_3(wk��.-<� ���z;��=�Wc�Ln��2�骲w�q��)�m������(m��.꿩_�8`?�ǽf� p��Q�OR}9ku�yк�F�q8�){��5D�E��AQ�rQ�͋ʉ��'�c��%1�m�b�S�z{Ů3'�;�Dm]^�PWc[]7&��k�|	Xo_Ng�\'������Y���-+]P�C7W+�}Omo3D�r�}Fz�1�]!�%
Z�'Ҟ��Nt��
�zjyʩOS�v���;|���3a��U>��wwr���[�ැI��v��ަ%�jˤ�W���?-�-3'�6]�mzg�5��n:tۢ����c`v��P:K�y!��Yc���cr�z��z-*"�g�(��[cz�cS�U�N������=�,.q7�M��S�C�u�����.z�J���\���ٛ�e.w1�"�	�G(�È�ί�4�������vwR�|���t����>����F�q���ux��X}�ܸ�m�u}ېp˱�0iܺ˕��K�;M��@������CX��J����������ŕ���q'r^����l7���f|\�8`ୖ���|�L(e<�r(���Ţ8pX���t2��۽�=�l��Z�凕��n��X2�,jfSR�`��9���Sk:r�*{���g���t�yw����av�
���ޯ{���HczM�#�[�(]_�]P�DѺ�����&9��I��I36V�:W����O�t�I�&ǲz'�՜9F���S�s��Qda��Lo(K���bq��&3�/Q>DQ�-A����r��X�(�[��^>۔��"��:y��y��1��(Ǽ'}W�L�o[S���sN�c�K�~J}s���k>���mJI��j�wU_1��a���5���o���c�Kٵu��Vyk>�7�H
��u�|jz�xS�8�|gb�Z1r�&lM+R��O�ۛ\©��.�R���y��(d��zv�͚Y>����M�V�ᓦn���7Gy�wpT��R]X��)����Q�Jo���E�����΅�I�.Z�J��]�Y��=X�b��z:�R�
��:H����UW�:d�Z���&i9�8<;Ǉ��뫝r��B+�K�N(���[Y�cflrt;fK0ؑ��8���E��I�S8@���S�r�C��c�v�.�D���W��D���8���v�8.[��B�F�&j-������+no��/��謻}snE�ʹn���,�0t�����
��j5I���h� �UR)�����<�ÐҴ�8�r�9U��f��V�&�.�J�.}�#�}Q�:T*EL�y&��CM���AIV__,�F�3 Q�Wx���f�|h��rt[{��B�2�|�c���������*6�o&�n�G�ѱ��+mu�Շgo:$B���2����LsyŮ�����ޠf~1S~�4���Wnҿg-;}�;-738�go��.X#nA,H9�G.���qKֆ�'(5x�-��EYxѐ�l��a�e/k��%_`v6��Lo6�y��&_z2T�ip���k��B��D�G�2iF�et��9jmJ�$�����Vt��8������sY�=�u���)�[�-�<ԅ�G��WlJ�u܆�Y#�оt1�T��8W&EzP��B�N�Y�S���t���M*�/p�_L6%ݮJ�䨚����QI��G��QTT�seX��F ��
���۸��/�q�S��ى�h˕=�����`��;�D�~�O�Q�)=��xz}t:v�:�ٹ��{8��k��sX��%�MG8��ɓ��3�Zu�NÙ(̸���.�[gk#��
rP#�h�Ƿ����ɛs�]��4�/�{j�*��������*b�>�Y�;�Q�1�}V�B��/,eg�ᣑ�tje4sU�x1I�����u�Ӎ�Ɠ�P�ܬHd��zՄQ�TWR�_V�މ������vY�b��������_l�iZ�7�B����&��bn0�ahr}\2�<�˃lM���ݼ���N��݉��8�m�9*��pS��De���D4��o5T]��������fa�Q�ذ���<�׀K�hy&�E���c�9��x�����#��2G(_N�6�sxi^s�s��e�U��L��/wA%l��(m,�ԁ�T��uM�M�^��ZT\�a�b���C����)��o�/@�9�VcPX��Ό�󜷢���J��t��[8�NZ����'�1��C*.�����kq,�1�N�t��-]B6g��`��.��p��;P�����(�]z���A$B�m�{+�����O�D��w]܍,]������d>5崺/��h+\E���;�[^�YM����wS]�E�ܼ��ˣ��6����>���:a3���G����C���^�������=�G�W;� ksk����	I�����ζ�~�Lgn�V�y�vC��]_�Xq�Yn&��]t����E�j�"�UQma�7Jq
�è�$���j��I�e�G��?mo����e!�Ӕ���0���޿��	ۦQ�]�Eu}�\��=�h�)DU��M��y;.�ܖ��*c�
����gt��G��NF�]�z2�1��V	�`��;���)��)TE�.���q��F� ]Vx�r�H����pr܋W�ǅ�-dn����St�7dN�`K���Ǟt�����u9$	y)��g��D�{No8*�m2��y��o�ѿ!\#�2zz4��,�ǬO���ƽ��'fk�/@�rP#8�l��\���m�C�]�7n�cm��Í�H`�	��֌nI7�y3#]�~�;����Gy),6��XY�WI&3d9r�ce����L�u:e��[вH������ܢp)�[U.��V������s��"���H�����;���8�y;ۈdȰ��0���:���U�|�R׾�D����L�j�FR�-V����Z��,>�C��LMKjiʛ-�!�6�1R�O���eM�M��hVg�q�,��x�>9�;����{U�l���I�g)�x�Z�j(�8����+�񽢌��II��c��J�q�r���/v][��ED�d�oSlB�44]���ڻ���B�n���M�o����zg�1ɡ�3��l�H��=rX9/z��O��b|�c]6�⎨��R�TYJ���B�R�߾}�<����ᘲ����>��+�Cp�us��8���rT���o5v�+�ZtXQ����6����8�*����bNt�>\������n��q0�f�+���a�I�;d3d�*��]��*v�DB��3	�����K�����E®;8q�g��H�Zz�ɶ峯�L�?	���/�=nUy%EX�/q���pE+/�l޽ofؽ�s�zҺNG^�omLk��,h��T��!C*}^H����G,g7|���^��e��j��6���hö��#�GΕ��0N�Ң�.��<�;8f��{��)�̋�ޏ����{ڶаl=��S�cׂùF��T�FG�Ι���P}����r==eqx(��)NҤ��
ټFd&�.���A,d�E��`[� ���mʲ^"_gw��C��5#ٛ�z������ѴI��Q��{K�d�R���E�� �8U��qx����;ЬT���*lc����|����s��	�_JTε�*�o<N��ݭ��^��J����+&�m�
Λ�vڦ��pNf[+���2�k�Xז>��#��u�����g7XB�8��]�Nd�<���6�.�+q,-ކ��l̤w�H�_m�
�ς��V�����&��]�3v��Fm�`��.	g��[Z�
b��0�0�Yo��6�BWV*�r_=	Yկx�m�n��:��W.Ɩ����8�"�ZJt��jX���#b�o{e��W�k$�^u�S�߯c��2�mm^k��(������\���Ǩ�H�z�F��j�jݧzp�a3�؈[ޤ����r���틹.	`'�����I�Swf�9��'�ޮm��@B��5�W�#~�e4��v�����̽Ջ�$�t��w���!vx>��<H�p��6�����\*�0g"�8F��cMz`�J$�%K9ΐ�n��z1=Jfm��t�k�Vr�8��ű�9fT�t,��k!Ĥ���`��4�Z�,���hж���
l7��+�F<�e�;���m9)[���J9�%Y�'N��7�^-CWA6�~��hֳ}"f�ﳶ��z/t~獻����5�n![� �&K5��v�]�f�f�.�z�r��I��goLN�7M�o*s�*_g>�Ɯ��6Huk�
oB��戀�P�0�MN�j�)�Ty�=�-֚G=�U7)��A�Ө:�!�p���ր5(�v��u��#�ھF�t&�:au;c`ns����u�	�R���[ײ��G�:�L�Ot�fvmK�Ku����C�.��=DH��{sUq���QI+��+&({b#��nI" ��ikAb�ABډP�d2�P�\k���J�Z�1
�kVUJ�VZ�Z���B�TX�[eV6ťj��*V*�T��%q�T�*����%E�T����lQ@m�[bőcl*DE��
��)*E�i-�Dj-mܰ�KYn[��E�%h��R�m*�Xն��"VE1�Z�)D+Z���˖�+XVX�)UR�����R���¥E�EU���[R���dmiR�ڔ-.[��-ZR�����TKj�m�X"+j���+P��V��3#���Z[R�R�l}s�����{Nߤ�m�Q�������X�[T9 !Ǹ_(���T�Һ�A�.�ٍ`--]b��vL�)v�{�N9 ���.k�"�^s�qVuf� 9xY��fShaZ1ˡ�2_k�͹:�9��iA�q�o`;��Sr�n&�&Uˮ��IEގ~ݰ;\�䈚�h�:&�"��$�'z�U��!����~�3��[T&����:V6�\:��QǇ}�jx9���|�̱<i�c$+�j���$Ŝ��J�\�b�s�cv��c��ͩZ���/=�R���7MTp����Y�Z����}�k;�Qsz���Cb�y	��[G$W
�o7wXV7���O=:�|��R/=+Y.�֪���K�h�3y����j+�kF���|J��{;הrv2k�R�xw
�<����s�LYV]^n���3����97�F��\��c"69Y��Z���K�f�ڢ��mmJ�)J��[ZV�9-�.u�ܚ���fF�/!�E�A�����7�4v]����VM�n�f�u�W����پR�9���Ȥ�vz�KY"�*��RL�FNY��Y�9�{�
y��9�m�/����^�m3�H�!PNur�F�c�/�+c�I"�m�Ǵ��q�/:nB�Φ7�
r]�R�����tR��v�D]�F:���g9?[�ԡҎ^/1H���<������1�qLk=J�uIz�\�����B;Iv=f��g�osA���4g��T=���]�I]
c��2�ߓՌ��zW)�a�VT���:x�r���tڳ��O�Ru��NZ�.�!C��^&&�ek�#j�h<,�T�U�ޥ��sn�f����^�P�{Z�"k��qe��KI>y[�Z;��@h�ri����HW�0B���\��B	n�d1w��T��z0�W�d��;w2U���a/�Tdv-��pڦ�^���
�=��}�z����shǔG�O�a��/)�Ydd�~fc5��W�,��
�peN�uy���C�ߵ��'x�f��}�E�SAu?X����Ɋ�{�{�]b�Ղ�=���WD��ql��ٞP�9�Ib�z�QlI�%��~�ɶ�o^���Yu��s�J�zV�	�ޑZ}%mJKd�/��-�g&�X��I*4p���gB��͂^va�;<S|�f�/��qOi�u�G4����1���uQ�^�X	]1�z���\����
:6��'� ��?�t���V��/t���9��b�]����mz�̖��.�3�b�Ak�H�08��$���%���8���\�LK��W:�W��ܢąɐP�ö��A��32^�o��db�}�ɛ��lϋ�čLڙ��P[t�Y���(�ټ�^�lVR��U`.t3�c����n�ۼ�Z�]qG���g�	��*l��P����ꬶN���W�3Dؙ�wk�m]Ԧ�u�7��
u�\�.^uv9^��pGe�_3b���v�9�{���=$w
ӗy��sOuB�+�J�h���72'��6���E�YO���y�C�9ICƖ���d-x[��=�p�������Z�ꎼ�\�*���ʚJ�jih��*οb�*��qP8���=��W,f�N�6��{��t����B�j�܍M� �IS|z���ʟY�m-�ջ�4��p��z��E)S���99�����yg�3j(w5�ʝu�l69����L�A��
��^ݹSj�rJ-ڷL�49q�!�6�BJ5�Z�Ɵ��+�g����irN�0���F��8��ƽH�r��z�����o�Ԫ�J��C������f�v�B6%��= �j����-�V��h��Z7n�&���y�w:m{T��0��a��9D- �CpS��!��c�]�{��\�;�F-z6ĎN#�X�oh�t@4���c��.�.��P/�Bѡ>�Er�t�U��w���QQ���5猂��S�`�k�-tL��2��zEm��zw��\�91��S�5앒����&�[�D�0z��}�^�v݆v�T+F3��y�n�2]���Y�5i�+2�+.��v��/66?	�}����g'zL�f�J�0`Cs�S�[����������G8DV�sj�����<|���=(��:K�5��"M�՚	x�}<�Yn��Qel�ϩ����Z�՝nޓLERŝ�򣚛�I���7�ܕ4ri�7�F���y.�������_���Z��k.�s���~���Ḯ��:Lg=I���x�>��@�����tIZb��c>Np��ವg��~1���
�ҏ��Oc����߈/Ɩ;��wM˖��+r��Y�WX/9l\m%�������oӛ*_W�ү7�{!mt���7T�ZmR�uM�~���Ol@[a�����e��tյ�W��Rr�������;}���qF�ڊ�B��֍��F���WO]��պ�}���mu�M�s^�ՅL�G�<�P��]��T�s�]�'H��+��I�+)K�wz��խ�L����I�[�D�C�e�'s4��l1{I�w��O�Y�N�O�wQ<��~̕�WC8�#�u?>�c�����y�(:#d���u׺�EE�E��2-5Z��`������7��Dg�Vu�Hļ��u5wo9SW.FSB�j��}�mv���qԛ7���ވ˷�,��t.[����!��@��mm\��d7O�+�,�T��Xo*��܊(\"e�M;�l���N��3�n,c]�X��wG+b^�'�C��½%�􎳔�1뵓uȷ�pN�uyG�3���dSG�
~���@��W��7-�gfQM�u�8s�a:�^)��)�呷 ��3�'�ӱL�Y= tJ5�){N=}aR��*�zrI�Ep}Ft|�''��ҞiK �_{��lG5����Ȣu��t�F\[+�;0�ҕ�ᔻ>��7a�R]O)�3�'j�A	�Of���.q���1НB$m��.�8W�>ʘi��$$�EI4�b�>��t�����QoD��|.M����H�Ȏ�>@���		���t���"�h�,�y�r3��s�nm��%�ܙ���>��.�D�8Kq�{ɔ����<E	*9���>d�Z"`�r�DB��\vE8pեM8]�v*�t�C=��A���B��IHpD(�[�l��Vc����q�U�q~@�����b+m�_	y����5��#��\}1#`<Hq�>�ɤo���w�Co{R�9}��q k�q#���4;�Up�l""`&�l8�E3�B+h�������똂�<~�{��7m?��l?@X�bf�r{��z�Hb`�B�6AS(?�̼�+3�!R)��VO��jD��i�=���j)���T���/'��j�X��!Y-ZO���8�t�e�޵m����D[�P���[da�PM3$\Ss.^�]�Mf`dAK���8J��'ZYO���w;@�J��Lk�ex\�������'#��P�(Ωt�n�|��}��6�%��.�r*��j@�.2�Gq���W��eSn'oz�8��D�݋��7���a~�P���~���p�� ��E��y]I#����K�A�6P��^�0�T��U�(�;�����GcIqo�F������w~��?c��>F���(A��
u�r\ꈑon�
瓽�d.܅Y)A���je����<��uK>.�Y�t.���d��}s���v}~�<i�"��(Z�F������qL����Dbާ+�1�g�b���Щ+��48�m�gqMAc#�FU����a׈(Ŝ���GE��e�ˎ�b��.}��#_5w�Ѡ����D]9���ř�F@}"i�f�}B�?3����C��_u�\���{�b�	��I�����d��p�{S���qlϯ��n��v*Tj��A���S*?n�k�9Wd�Akk��q��6��p��|��cE<�{0v���;X�Q����t�󯽜��љ��E����Ň4�~d��|{V�aᮋ��W8����0�� ��uu.+�{/iЩx�m]����J.2�6����� ��#�c� 3��	[4������#����ga�V�&	��j1�Pȯ]^�!D�2�d&}!��(���ػ�2O,��0"�P��S��ױ�/-��[~���}{j/W��E�J6�jW*Ei�L���|�i|l�yR�%^*�]{��:;ۛK9M[�pT;r-�D`G!p�*B|3f`¨>��r�3�;��f;�¼���(�6v'HQq\s���J&�@����ȯ_��/]�ثJ��;YS���|��5�"]mll(H�o��@�ldm�Wm75�V����6�̟t�}��]��p�O0�|��|���x������'���*5+UUE�����Ɵ��EE=~JPsEE4�OF$#t�JR�Z��\i��
&����o�	�>KI�����b2��m�H�BHH�		 �B@�!$�6'����B�� L`��E2�MLp�I����h�lkQO��1�ϝ7�}���4��*���=
�[�b��^�3E���<��yJ~��aJO���O?�K�!�Ca���8��S�)��<u��\��\P;QQO� �
����$J-NI��L�j(���\�=,P�uT2����~�F��Ӛ,��y"���Om>eS�r"�M6R��{P�t0 ����i�4"YI��⅊�J}�`4�i[��w�"m^p����s�w]!v�d�A��P!	! ��ɲ�FM���?���D:�
d�(
$�P�a$��hԠX51�R�P�C�,L�\MzG�05�DTSZ�K�$�ho.����5��=�JV�Om���=�w�Ѷ�������Ǵ:
>߸�+1�K�45��Q�1���TM�榲�%?@ytCgΥ����}�*:��LQ=܊z���ڝ��]�Y�9&̀�����z7�^�ܘ�Nj���:ȱ&\=}C'�z�V\��ɐT�> P�ג�#J��ETR$*������@�!�KDG��IA7��h�5`.^i� e�<���������m� H� ��I����.�LPUQJ$[ÈSy�.�!��>9��~�Ԕ������U��=�A��7-c&�'�,�.���hj���iT�TR`�� �*�������>�C���F�P�����`�R�N�޺�(3�uBI���Hrtt��Ob�|Sj�|w�L���(���q:;���7 2y)JD9�}Bd�Ԡ��Q}����2j!�'����Jt�h]�jw ��'�:��dD�B5H����"U��3Y���O�P.��D�>�2j���U1����;S]�QJ������T5Ӳ�"dC����k܎�2'�"j(c�zoȰ�(P=�eN�#�#QQO������x�S8 �o���Ϩ���w$[��.=����˥Ɉ[��Ukb��I@�����4��t�q���)��/l�