BZh91AY&SY.D��ߔpy����߰����  a��I�      >��  �@ � ���
@   �    Cs 4)
�
P@�@f�      q` \N�3�m��8��i�ӻk�ps��ֻs�Z����9N�;���m������U.Ǝ�{5!@��hB�x��ْJ[v�v�T��$N �1���T�ݲ��[j�����h�f�٥L�w*9��3�8Ί��u]����;���EM�Tk�t��ʫc%4 .   wUkv�v�f�[jI��GM]��dˣ�p7%�C���9�Y�ƹ��U�G]���݁���ˎ��v�3��     wFݻ�r�Z��pwF�rV��vҊ�L�+v��'�����q�G;k����;]��hh5m�`�  " �s���N��q��6�u�;�a��iv8 f��\�mW8�v2���j����GKcJ��W�        P           P�*    �J��g�R�!3@b`C ��h`�?ЈRURz  �&�  2i���i��4�0LL��S� ���!�Fh4�F4� �
���4���A�x��z#�6$g�=O�Q@BT�yL�`� �&#F�4����qq���ے�r���I�r���̕����¾�$���jcS��>vٛf���zLfټ������.8p�|s�6͛ỳg�����ˆ����J�g���ՂAI��"D�ʎ����\a�Z��M"I�7E�x43���*���l�V�,c�c������K��|�]>�fގ���	�������J?��_�&>'�1��,�G�D����$�鄱=���{0�t��w8x��1	�\'KL<p��p��ç�'��IH�c�1��<UD�1�P�$�"��QD�1e�N�Ϧ:#�'%��0�Y��"��f8C�Lt��L$���pN��,鞄�;0�p�Ҏ�HH��K��$�/&I2p��za<#ۘL0��=���c���X�va�,��G���,��%�8QʒlF�O	r�x�F#����L""�	�w�1B	��X�xN�&A%��c��,D/&0��dŞ8<�� F*a(��â	�*:'�Ј��3	���A��:�Ğ��#p�������Naۈ8#|&F�����b" �<'��"�{pF���:D�d?C�:v���DNz&��x��L�,�Bx��~��1=�G!0�	�L:Wy�Ye���K8K�?IF#>'�A�|�93�:�bDK�LW��F���3�Bt�$�u���$�$����=�Ŗy�2$�K1��RJ&y��0�f1����zO���"8pA��)"I�Q �ɉ(&#��Q�>��"� ¢"c������"cُ#1���'������\��ވ�%s�	�}eT"_�0�5	�#�#�DL˘������E�2"���+���BYC˘O	G���aBTGDF�a��ơ'����"p�A�>�D��@�33��"#1���.LaBz�������.;0��=�B"��,���J'}1D�ʙK9���D��#����	��;��#qd��>(F!0Kb~�J���"J�D�l���(��xO%��ct�8�OD<#�D��G�&�H}��ħK;�$j%+�&1��u҄��D��Aǉ��N��a�B&=1G��H+2%:Y��И"xb",�G�Hj%8"u�J"v��: �@��1%�BP�"'^DЉ�G��'�BtO5��y	$D$��'��"1p~�A�D|�Ώb�'	؈KH��DȒA�\$	<bd�(N��K=��X��x$��'��%$��?B'L��5�'G>�	⇜'���a�$�$�<Q�"4�{I�?p��#Ј��8Nrٙ<"�%�	�-�J`�.D�a��0��'�x�gl����|��9�&͚�-h�H�tk�H�(Z��O&
����N�}0���6̦f_�0���"y�/�#����'.<�~aD�E�Q?Yd�DB#p�LAf@�|��d�pD����N�ff���̥v$�<�Ja�ߡ0y���e�DQ�?{�bRH�L�bĐK@�E����}rW��Y_U�%C�Z�|�||�y���ϥ�*8pG�BpN93��ř�������pD��>�nfp�ވ��AӌĢ[Ȕ�j'�F���q(�lO��&,JAlth���Lb#�ȓ�Q(�BIo�d0�/bQ���bx@��<,Y"=�OȐ�>(N�b$�����ra=BQLD'�E��J=�0F�e<tä����CȔ��Dr&�$��=��tN���\bx@P��"p�s=�,M���L�����ڙJ0{�py11�#�JX�=u�bǾ��b~�+��y��=	����>�����,���`�9��X�"|'��DGb8%#2�A�N@��D$��b!(Kď��-Ģp��`��Β��> ����'��A�IDL䒘`�<@�8%��zQ�z�(OS1�v��|�@���	(���Nߦ��a�2!0L�`a,��D�U���Y���=�2YԈ�ga���y3"q��\%�M����:#�E��:[�zA1Ϧ�jX"�騔�ĥ�/N9�e:p�>������,��OG~����m5ժrS��*ݦ�-Y�GIY�0�fd�}	E3�:q���$���C��ETH�|��r:!�<���~�L�}�fe$I�J���Ɠ��o���~?�>�	���lDG#	>�DN�73)�a~��P����ɔ���ǹ38p�}p}�X��P����~��N�a<#�$�%�(OL"=�r&��bzpG��~����?<�Dn/����F?G��D���'�8%��O<ȟ�~�B'��D���舉"a^Ģy�J`��&ı̉�1<,����H' A����&؟8q��u�J_#�ŉ���,o�=�Ȉ�$g��&�ĹH�f�vrN��3 ���]B'{#p�s�#�q10��<91�ta��M��%}ƾ:��C���k�>��Ĥ�/"lN���v�����R�X���������DG�K&�;�=�#,���#��<pz*(�N�D����x�bH,��$��:�Q��!8_K:3q҄�s��QT'��LN�#��x���&��(�f(I��/�Q�'Lx�E��:q8O�;�v�-$E��1f0{a��O�f>G"DǓ
c��Q���xJ"=$�DO��Bc�n$I����'�E��'&J(J HI|�Q,I��#�LtJ:'F#�t[���D�0�pJD��d�#Ѕ,���Nra(N�f,�1��˘�{pM4��)҄�$�<f$�Dn$D���>���tL�&	���D�"`�'{	ӂQ��A�s������2�:�by���H�fs&>K�c�c1'7̋9���Ou�#3C=���eE��@�>���A*#��ǆ�0�na�?s#�"G�ʬ��A?�Հ�u5ۆ�<w[񒾾�Ş����]���A���,���S�����g92C�~;�Xݳ'�w��ݢ��f�o�4�gr�VX~�\���>g2�ۓ~�G�Dl�ݗN��û�80/
>����:�zt�NM|�3���N�MM��T�5Z޼)o�\`��'�2�r�a�;�5z�?������-c�V��O�fw?��LOs�Ә[�W����~��^�{��X�U�L��{�g�u�u��jg��n�M0O���������?s��5�Y�õ�y�O�zR��3�{oG�+��_����Zof��?��s��������9�]OO��=�!����;��$�V���*|�N��y6>zC��Ó�#C��^�F��K�M8}��=�|��~7�O��������E��S���1�9��yo7�/e��9��x�tf0�L����b\!�9?Q�&��q��%ޓ�&ɜ���r��ַbv��}��y�	���W�w�o�ג��x���m���m�2�2Y/��rw�r����~�τ����8m���q�7�3���n3��]��A'��I��l��6lZ7�?vL���e�#=z_��N^O��/ ������?�;tD�
(/ƙ��8�x�������	���#������e�s��}oܪ���nU����7���-�n���NCSs�3E�~�]��Op��?���=ѷ�/<�J.�&�N����=����3�Qs9���#�ҟ�#M�Wgo�nul�������}W�� �f�3���7]��{�����S�q�����G}�����'-k�妟/ǋ�	�oXu����s�7Y���y��s�{:U�9y_��_���|�8v�)\���2�~ghh���w��cX2�ӡW���'d>	����֩����罪��e����Ts8���Ŝ�������o��n\w�ߝ�{}^x��)���֖z'��f���B
7����&�\�f�q�)U�v��Y�h���&�}��a|���YŃ�V�i�&��бg�|k���.A���>ظ�2���ox��}�����fJ/�.o{���l�-ֽ�?�ɝ��KL������yg�>���_��*_���\��͜�c\��o��_�9{��}:Af����"�.U�ƅ�vn�a=]g�ym�?=N���������wy73_�fd��חk��S�륿4߹�v�sc�=i��^�ӷ���K���m�$mv�2k�+�Z�A�'33��e����q^sw��8U��4���N�N{;�Ǽ��n��5�b��b��{�d���d�6qD��3f��u�W��+旜5s���s}�9�o_;RՎ{�齠�9⋃Z�ofF]�i9|�����Ы�s���x�n?<�1��4�p��I�W��eOK��n�lm����~>\��m�~ބ�.��=!���϶�+����^��,@�͏��0�˄>P�/B�nY�=�i��<~�f��]�M)�w97)��nzr��Z��͟����9:��On�1�l��x�璝��s��_�0�,�g�b�#�o�g�_<��NE?o�I�t����iR�K�c8w"sW��~��7��S�V���d�M�q�?d:d��M��{�5��g|�M�#��.���ݜ7{�����5�3��̓9��d^�G��Dj����Of�� ͂]��u����[��.���z���g5Y�7�c���o������9F}��<_�����H�����qFN�N-<��x�t۷ҍq���^xQqfN,�ÛH3���w��]��H��|�B���՟����?w2�"�[�0�����gW��.Y�pJ��d�*���|��Xl7=��VM�G�nO;���gO������=ќ�/�}Ț�����uo(��r���ޭ�s>��Sg�����=��m�?�P�.v���7\.O�;� �ϝw2�x~̏��Qu���I+���z���V~}��b�,�����M�g|b�:�e�3y���\���8mZp���õ'7�ي3wyl��;ɝW8�yx>'����j[0];j����X(�n����e�7T�7�)��ŏ7��t��z_����$0�Yo�����=7����ޜ&syO�ۺ����/�������ѷ&q�>^��t�h����;�͚\V������ɪ=�t�Q�=Z�$�x�{J�b�g�s0۸}��dsi��4�Vz3��p}~�QuuQW�/׹���� �Ս[���3#�&\�zp�2o.ݽ?gg{g	6Rh�ɷ�6sKD�7y{�pd�܈��?�켶7$��wl�� ��n�Þ}���|Or'K��|m�o�γ^\�'����9E��y�ܩ�{�����^����t�1/�|3Z���+�s�[��4=�i�'������������_�����\��H��ч�/�ͩ�����n0g��f�yqݑ��})��8�;�٣�%��Ӧ`v^��{�7���>z��N���W4��,��Nn�����zsS��,���,]�8�g�/��<{+Xd�S3�pe�s��zkxo9�.i\��8=��w8�8�:>���G���3ل���޽���5ࡿ�<{|~O��|<O�=xnc1�I��9��6s�<m�����;�1ְ���ӛ% ?˛�uo;!��0�ɓ���p���W](���M���������$�3n��Fm��(d����]G:?�0�b��&?���t?q��sƚl���<t`o��縹9�Z*+94ޗk��=q
{Gy����'���r~?�N��O�g7���ޜe(��_k0��a�Ǘ{ܛ��x\G�mT�%���o���w��\�'G����ȴ����=зrE���6�l�����rk�z�����LWk���߿H2�do�{م���nW��t̒fW���G}�ɟ�y�#:������K�h��Ç;������fg�������f��v����ӊ}�䥽�g�J�����fB�f�s2g�0��J �0�<XY���������߮�� 碄�g9�e(^��gk�z~��7����OfUrrB0�;���|��	g�yw���vd��I�䞟��3���~�9,�y���!�L�nC��$��{3ݻ���;]�}V3�$}�W���3f"�~�ژ��Q�+�}y].�x�#�ϡ_��y.Ofa"*��J~&������~���
aJi���)L�RGi�s;���/~\�|����=�����?�f`�;�-�����:ݿ�m��;�el���o��
�����
F����"��"�}�oO��xgf[ۿwg���盶�<�>J���kg�W)����{z��ux��������ӗNt�4��@ʪ
�D�R�4(�DO�Ed+�i�����5pTc�+���pb�*$AT�i��*�J���U�k���k�RX1�[���2������$c�O��J@o��A�D�p�@�g��4�c��J�MѲ�O�%��lV�V���}d��M���:}�1�@X��?
ܟ
>����دմ�8Ir�����(��q�jͤ���Me4�^�k7�^�W�9s���~�ZF��j �Bo�!͑�u�Gc�}Z�G���NBIp��ƚ�'���uڠG��nm���i�������v��[R���h��l�7Q`؆8�&���S�/���Bt�0N�DEh�NW	S�[>����-�]��EW��h1�����˗�Ϭ��4n�5��r�pkN��ZK�HM�����!���Ѫ;�52��nR���VI��(��6B�
K�`PG�=����q(dF(�	W!��풔�Z¡����5~��W�#��thJD��譣��V��,���mR֐�Q�ߣv�"tN�va�Y��xd���'��*ڎ�iT�B�+g�6^��/���QAX�ò|���g�Ue�Dh�Q�IUCE!k�U��m�\M��p\݉����i�$��	#,�;c%���`5b���(��!��PV����
���]���*L�������<Y�&��o�#�e��o�kJ�j�{\1FJ1�[�f�z�N�D�ado,:�x�K�S&Z�hNJ��M8�,����} ċa,��BQf.����~����إa9�>1�qa�g���)	,�Z?��hB]�u娏��fQUkL�ъܑ6���ݼ�.mq�n �~���@��뺓P���;��V�k�TG/Ŭ����q4�E���F��/97f�kv�B%(��7b�!!��L�S�j�(&5^���X��7$o�� ��H�����u��������ņ0�ENEb#�����>Y�	�u��Kv��J8�MCD�c�ꏐ֮�C��6�h:�w9��A�1��Y/Y@��5B�K�ﲷ����+���,/%gyt�i�n�;��k�/].��\N}��oWhG���^4�m��q�4%�M��mC�<��;�m�&�e�5���x���wn����w.�}�g��=��'$��x��������)���ه���v��N-�}A�?��og������lVcV�ֆ����*�k����^��U��eU[VUU�UUTUU�����q�UWUU��W��U�UmUUUUUmdUU��U�H�����$-"�=�|�W��U|�*�Ux��U겪��*��wswj����������ZUx��YUVՕUmaUWUUQU�����>���>� "���>�^qEUUEUWUU��*�|�*�Ux��W33.�j�U�U򲪭�*��*��iUz��W��UiU|���j����D}�@D�A��������U��U\EUUEU[YUU��YUm����|�*�Ux��U겪�����*��ʪ�V�W��Ux�����}�$�X�VI"��"1m�4�x�y��6l٢�)J��ϟ�������Ǆ�y�O77777���p�Д@�$�H�BX��'�&"xA0�0L��Y'�<'��	��DDO"I"Q"@�B!��"`�e ��^��==�ۖ�ٶ�[== �D$I(DDDČI$AD�(N'DO$tD��,L,K��b$&,O	��:'N�'��N�xDL<tO	$	���K�	BQB'�bxI,D�0D�Ǯ��֟I:����{..d\U������VV;e���;>��j�G+d��~����4'�*'[p� ��TʠF�Сn;���xʓo��Tݭ���(�#ܹ��L3����_�ؖ ds*j��B�I�4̃�G+ByF�_���*��V�l�#nX�Qh݄��ʥ���a�PB�5�,�0dC�k�Cs���޵31��(�Zg�$�-.D��VY�`�W��[Yc��U>NI+�V�����h��V?���E	>cu@)�d\��n	�NS�T���?�pţV��pV���y/ѺTڒ�h�r�(!��ڨ
[F}�c�`Q�!]j�����$����jG��+��@�����D���I�T ~�bLpRX#$�㈘��}[���b`��@'ֺ��⮢�B���m+��ml�(�(�O��eVVV�N�U��4�>�B#��H�A�J8��R|%b��+���VHJVV87dm�Ҭ�C)[ F�&�+vN���cr�&�ei�jv�lrK,��%$Q�Z�r��o�LX�1���b,ȡ���lM
�[,U�cd�D�r�	l�R8�H´LCV���Ȭ����-
*�?I��!��܊�X�d�����r�$��H��rV)��
F�T�((��q(몴'V;ZcA]E$���}�����7hݵ��25M�o���"dm")h#n��]CM��FC�%�;�}Q�T�N1B�Z�vTr<�P�*NR���_�U����󎉩D�N�V":�Q��YM�B�F��J�A�����vEh�)i/�XV�/�����4ُ>��"��X�W�$AI,�;?�u�K����r�v�#�6�s�	����Dib��kd����2(65%���X�AͱEF��cacҹJ�l��-������Q���r�I14�,�G�U�K,B�"���i�d�&b�F�<vD
�����X1":�M7$���Q����%}�+�V��M��mMؚ%T����W]!~G�Dso�4֟F�MO�u�+\-��5)*�߫��*������qY�ڎ�A�n���I�ab��j������4*T8&VƮJrHKF�X7e�k��*��g��������w��>�www.���tt�������ܻ�������wwwr����G~>�����M<if�Y��%�%�%�:h���٬���,��;�.�\RKkM8�D��6���PA;S��F���B��@�#CM�`�ԓ��V�l(F�ߑ]�TM�g�;�mA��2|&1W\qVr�~xw Gq��K!l�(J5"���j�WG��$��Q��H�qW`�}ڷM>r#��mL��2GN�!�V�)�僑D���Y��K�`>d���_���7	�$18��ۭ̟��G#45��qAbR)]-� ��O�BW|�Rw2�:���F��od\֕��]y�Y�����Nc��,��.��.�:'���۟b�n�r���l��J�trk#I^!�X�L�Ӥ��>O��T۫/#��m��p����k�N����G�vo�\3�����}�eu&�Z�.��t��LM7���$]jS�Stg7��.�&����~�f���i��$D���:`�>�^��[�FZ���.��T9ı�n�~�`����%�t�j�IɼQM��	_pg�1��3=�8�q�n�����yw|�_�N�47cwhcYd^�I¥�5E��$�Ԑ�Gm�æQ���_��9s�;g�I�����a�%�$D���:`��R0�TG�M&}�;ST��1T�1ء�MV��hجl�鹪�����g$$�!�M2��u�W�kW׮�k�ǑNc���\qElUx���9Ip>:Y��{� Y�_Q0��E9��h�r'c��g��y��2�9�Z�	:h�ݜ�d�r�Ѻ�ӥ�I&>(Ox�M�"@�BQ�:|l�6G[#m,�L7 ɪ�F���D���`f)�ϡQ1w2d�Ł�[��p�8aTY"��v���tHe�Wz>�ŕ�l��Ŕ�v�!�3Vj��K���Q�iS���I��9�0�Đ��D�GN��<'� D�(��'�<rYy<���g���8鏈�Y��w�d��+�r�Q<|�wǫ^E�w3��́s7*Q6���(�eu�'����9{���/�o�������`|����n�ә1t:�Qw��6�.-�\����e�N.���Û�._���	A��/�:��2��R�����M���[���s�J"ӑ�DV&�p�w3	L�y�����!��%��2��
Q���գ��L�3��+�eҜ�ұ�d�ن�J�G]m��0��� D���:`��\6\�--*�X�E�KE)I���%R��mQr��k�^��T7B4�h��)Ֆg�!s/&a�Z�}0w~{#��ί#׳��V�,�O]��2�ר��@r���s�]e����r���U��� `�̸̛\���֠�l�Vڝo�|�g��+�|�T�W�U^�,b2☏���}�t����"��#�L����=z���%	Ft�<'�&��b�&"��e�&�r���\^Vq��t�U*�m���+�<�3F��d��0l˰��d2�\l2H�=��8��~�~�W�f+ݮ���9�n:�I���諆��Q�ީ����h�9G�:�Z���N��:Ԉ�`��:�M<'� D�(��'��P���nZ���]U)�Z��Is�P���v�<��T��Gw*�����W2�e�0���w	t��P�J&k���e�Ôh�𛻖DU9\�ku+D ��,P�cD��mlh,�UU¾4h�f�|I���=�]Q����*�;�]�^��th��(J���}蔢7K��<p�f�x頉%	Ft�<'�=o�g%���Kp��ت���_�ܩ��p��RR�}S-�1�5_.Z���F`1��J[6�'҈&!����Y�ci����c�Wb���]IB޹g��.MN�1vr�E�=�	����i�j7V�s�93�f�֮f��pY�����r��������>���-��	��p��!�r�������f�ZY/S�kEB
�,���BU��H]V�Nr�y{4ܿ�ʮ����w��9ϖ2���i��\eꝭ��Ε��ݜ:J����@>�V27r6&x+P�[`�j�%�F�?-hiӁ9�����>%f���g�ވ��Â%�4�M<tAJ�:�uyj��(^h_a��SQ(L��&���>�QU<wgKW�c�]�)�e�m�՚�-ÒS��R���r�D�fX�׈n��.�c��Ì��l�,wuV������Gh�
��0����,��WV`��p�D��e0H8�{��tC����<���DD�g�Z{Տ���Z���Ymy�l�C�Y�$Sf��h����o�˃� �َ�UV�O&�'Ɠ��t�t�I4�"�Bp�Rt�t�4Ұ�l�'D�TF�I�Jӧ��<x�<\<OKH>ǉ���G��j<<_���������x�<>! �=��v(�Q��X�أ�_�	��:3ŉ<H��'�Ǣ�|><N�,�Y<���|Y?/�h�M�������K�F�%I��iBi8t�L4�� H�0�
����0�<N�&g��e���x�<h��&��t�|O���l|p�}D}QO�CŒ�O	���:?/ı��?'��
�Y%�<
L��H�	��O���/�/���.�￿����R
L��a�\!��\���IN�t�"ŭ�g�׷J�����J�z��s�q����3�x���zE������DN��E���ĶtcW�5�r+����?5ˏ�:s�̇�W�Kv{��c��w7/�̙/��joW�����Wh�}���/�d\��|�&�L|�s~����߶6~67wws.���G~7wy����w{��ۻ�����̽���4�h�x頚i,����8xؙ�ԋ-UQ�|R@0�,�-�x���ِb��� ⛋'�02�!j4�L6�0ȘF�s��ڎ��eb9P���V��~����$�(�w*�YJ��<r`��ޮ_�ڧb������>BB��{�[VK(�"S�RY���3����O~ČAG��V*3a���F���3�bx�U9d��qT|�a�vL�K&��I�5'�Xڤ2W�R�6ITZ��yL�$�9���%*2��2M�-��0z���!�X�,eX�?[^/�bܮ4]�$uUY�K*�Fj�ԅV1����LLHp�~Oǎ��i&�Q�N���&G9��T�Jӭ|���
�"TrY*��3,aC��-�1�ԭŶ�9Jd��n5����$�H���FV$�Ouk,����K(���'3�ݷ�v�B��֝h�ə�G&���phު��	��u[���9�q�ے�I]�#K,IM�ő��g]Τ��8!��!$��( �4��$�,�q���2Y��$�aUGZ��_��2�|@0LJ0j��]L�q��%�f�\��jY6�������"��K#��mJ�l�����m�0��U2w�+
�Z̩+a0UzԵ�¼���E�b2�����ȫ�_#.�M�a��ňt2Qd�D�ST��F���Ecn�'��r�Y+\~z�����$iF�Q�N�K4�$����cN<���_��n��y�nF,̸�
֮6b�4+$��h��j�'��P��(Y�klN2?��Ue�Y1�b�PJ��Ҫp,t�؋J���+�*}b��D4 >�����\���E�����.�ǀ��y�y�O���U�+sru�P�Ňzs��jjv�ͳ3;�_=W�ƥ�=?z��Y�UY�������c��o}7�UV� ����T����a�����#�7Ge����eU�a1*��|���k80~�MQ����h����b0�*BPz/��n�t4j���Ȱ§�#i�UM�zBIWF�CBW(�U�]��DNT�o3����>���):�
��UJ�n�a��
u����KR�ݸFl-eUF�3Rņ1�b��S8b��GbI�U~{o�[?]�'0r,���e��ˑ?eU���"_�ސ�d����[	Q͕��n����𩺣�%},>��11'U+�T�s�0�2V�\#fX~��v���)8�`�Y1��&��ņ�`��G?~���G�#M$�J4��gǎ6N_��Z�=���������$��qM@��Ҝ�3+*�$����z�̍X��`��g��f�*uYY2�)0��a?x�nr	�0�ō*aY�P���H�	e�X���BY�a��L�#-L��R׻�,�uӡtY[��nUa
�5?,bzÊ�d�����&
v�Y��EaUb0�L`�Tı��B���=CAb!��$�I���tY<_���)�ds-���R��T��+jŊ�$���LF��K���d��n��Ud�)�,~��R�V,3���k"%�����%��
���+?i�Ւ�[J�SVKW
��5k�����m$�2�*�>S�f,�Tв{)���4L?�M4�M(ӧM�8x�h��-X�=4�����'\z�*��i�a�uS+-EU�&TŊ����I��Y0�a���C�p(�lD�*��(������֝&qe&��9rqUTԯ����1S(�*79M2E�7�a��`���������9��=�̻1MQ�!���bC1O�1b�Ѩ����}F��P��A5PN�^=�-Ļ�6V�7[%��9U֊CtB���^�c���u�FJ��eUϩ��O�}�j^�ܨ�d�F�J~j���J��T,�)UU=��LGTa�ّ�%�
A�R�:|"ݕ�`Y��*�j�iJs��.jK,�9�e��W�ʞ,?Eg-�S62��F�0���b�EZ��0~Y��Ͳ�XF�+L�U~�#S�Y>m�U?2�*��I�M�[V�ǹ�`��NSȰ�����񆟏�x速�$�J4���if�8mͷ/�˒���]kƇ��$��Jp�����vrs�9B����g$V(K(�GE�XY0��őp�)��K��9���'���%����)O4�a�I(�':GK_�C��黚��3e?��{Y�����O��Y3��ȵ�`�x�M)�cR�J�_��)J��R��{ҳ���A�ɚ.o��f5_K$�x�<��M�ƫ�}'���q%Utj�H��,�X�"w?Q���"N�K!%�D ~��)U�|a45>)��iB2��B�㌿=չm��eJU�KV� AE �t]�<h�3쑎eT$�Ui(��O�`Y�!W�Sc&Sɟz����JZ�O���?�ǎ�	��i�t���4��j�8��D
l���`�9��lpV�Nƫx��d�&Z�Dۉ	=��Y�������i�n������vF��E(��qAR|�F�U@`�c�Y� ����Ş��*�$k\{�lG���3;n[$�*վ��d}Y���z욈u��ѾfK^�x���}G5/Io�����}9!͚7➾���fc�5G�}ϛ�U&��%B	t\9R2�)��I�
�H�㴈�~0��rD'�Hd�e����Z�,�j��ImU��/f
uLz���	cX}	\����h���b'�x�Ό e�ְ���UYG�04A��v��4&�?de���D�����:��7��6~:CB`|T��+,��J�_i�A�j�g�U��"��T*V̱��h����&��'ΗΪ�W2�16�]��3��	�'�(�O�z���T���s��1w�6���=3Ӧ�?i���L�i&�Q�N�><p�K\O{R�N�0�]�vuUPD���	����~8h�.�G���3�rʕS
�Yfawa9�⳸�
�bSF�F�d����'iP���$�¶%`���I���B첸��]H)PJ�
G���0w�pʵ�웯njN8~��0�a5)�'s&߬�6�!�puL+F�{b��%�K-$�˳e{���$�h�hL>

_Ip���a�#	Ĭ�Ɍ�e{Z��"O�L(M�@�%;!�|,!ߖ�Ր��"%JN�> x��~�=۲�)��Y98���ׯ�4�x速�$�J4���if�8/��%�dQ���:UT+{Dߑ]V��@D���ai��U}B_-��"	�
�He'*t��Zb2�T�W�Ro-2���V.;m���U�Y�S*1\��*ˆ�u��!z�P:og'3ƋcP��rYl���V�I$J�.�D�����X�Z�\Sj��ajW�2���!�԰�CD��L�����}��i) "?�A�mza\��>�r��0��	��%�7����
�����9F
?he� �n����b��hK;3�k��q�O�>~q���ƒi�t���4�O"}D|D��u�UPNT*Q����������G��CZ��z�4¦L&@�� %�����T4j����v8�1HA̘n�?,��CpÆ��6�X��~��1)]L�+��w��0�q��V�Tn���0LR	�<0�@����e��5-X��Y*�.�ʷ�[��������5�*�eUT����ҩ��t�D���l`J���2Ri�������6�rm��c+ٔ�������O��F���x�A��4��QZEMN�M�O�'L'HOP����?��#Bƒ��H�$��xx><t�p���'�'���x�<t�8O�0�Y�i�z>$�I��sO��xi�i��	D�GC��x���	F�A��,�;�S	��z>�'�$<C�'�$<Hx���[�x|z/��Œ�x=�d���V�<~9��~?	_��i:�M'HM$�:h�a��i	�1��h�p�4����fl�]��'�G3c����l��_��p|�'e���|K'��C�𧢞4K>'���x��a:Y�a��o!4�N���di�o�ob��~�v=����]����_��1�os4��+��%Cud��y�����n�y�wqv���~x��G׷˯l�a�.���������\9�~�[�jli���*�ՙ���g�/;~�|ܦ}��ɘ�2���<�s�k`̶L;�Ų=\�/կ_�E��CBs�1Q$��-�L��gӾ�෎��.d8�K�{���G�B/A✷��i�<��7�9A`L�.O]^���'� ����ӛ-�=�.�N��ê� ӏN��g9^wǱq���̮l��ple�\"���[�7&�8[�ǭc-���f������o�i�޼݋�i�1��	0��p���R7�mż�}�y�N��x�Zh/%"��BS�?$�\[�Tq�q!+#M��Y�ec��6��TGKa��O��Id�MF0�@e����8�%UA�[�x�C"�ڛ�\�+R���	S�l�-rbc�G	O����k��dZU^MU�LX�\�t���^8rU�y��<��*>��mg$�͕Xӕ���ё��5 ��h�w���'�����e������*���fff骪��fff�ª�������	�<"`�:`&�I��iGD���㇍��l���.�%Y/*�u�X�Qn&ڒ}+��$m�Sev�cE
�2W+�CU�4�(��h�Z�#(�ڒ�[(��I%�"�Ț5!�X���PЍ%��H��PrY���r[��vd����'d,D���+���'ѡ���%V;r�k�|66���N@`�V�F�70T2:� �!b"�V!�$�K"aS����`����Hg3��;���vK疿"/j��sφDs������@������=�\UC,���>&	���lke�H	 
=O[�5
ka�(���tg4I��~�OJ]��)k�u��Q��P��*
�yE��H҇�gԈ���O�1/��م��P49���.�ت�؇��ç�&Ƌ4r���J��ڪ�4���Ir�V���fQ�0�fx�i֏�UU�k�4�g5\,��n��o� ����ʨ��20������&[���ܾ�0iշ�ֶ�2�׏_?8��ׯĚi�J:"xM,��yg("c�g��l�����V��J�ϸ{��N��5?LU��x�1ί���ܵMo*nnjg`Y�oya��µ�ӓ�q������2پ�7�MV��Gh�� `��P�	�X�^N(����A����U�I[��kq:�7F�NO�e���1��P+��ޏWD5TY��NA�.}N�(�3��%���c�r�����Лm׎:���=z~$�NQ��if�6_N�dDz�)`��X��E���*��:s�8�����E���S�-��_qpM8��Ʉer��#����L�����{F�|r����O�]c��0ш��~��6h��,�%�u-����?L��Ɖ�s�L�}-UY�.|��c�#}%}�1[��!���&W��Ɛ����\��uv�_�����V���92�2��7������>z�����48-&R]U���ǧ�af���j���֗-|��w�a�q����0 �i�(���4�O]�?Q���u3*�Z]�Ui	MJ�^ڤ,����	��M��h�R�0���=�Y�n%�-1nf0�`��Ļ�����/�_��?R��·oyg��4�x��m?=n8��;��j���5GIӛ�À�t]U��H���r���z�a��o�t{߆�w%˻�NQ.���!��l4��ˏ�e�Ӭ̴p�#L���4��/��'M�`?yxa�M!*`�4p�&����4ӆ�pD�Y���ܼ���o6�R��Î��kƜwןZ���
}�Tw�CN�)���r�9�Ȝ\͋)9$3g.b�ͻ���9�ȟ�JŊ�KS�R�[�c��O��6[$����1��<���	�U�5��lw�ڋ��x�B�n'�2~z��gN�;�\��k풳��Y���O�"�k!kr�i�~�Tz�C9F�a�(�x�~e=��1�m3���.1�;2�}r�F�2�a��rz���\g�ط����?����������뉸�j�~����1m�Y���Y�h�%��Mk5˒]otћ?|m���bB�T7XDl��2�W��d�ƛ�w �lY?+F���WQ��w�p���z����9f��a�q��]�צXeǏ��?=q�4ӆ�'D�Y�w�E�v�SZԖ�B0��K��\UZC�?pw�?Qc��gNѯY��9��d!��n�s�G9z$�6Z�%��F���*�,����򳷌?V�>� �J{��z�l�?I,�C���"@Ѩ)fue$�kThC^7?]DO��d��FJ�60U$�q<m=G޹^�;���a��bo~G�GN���gh�!�A,�D}/˲�)�Ku��㓮ǳƗ�̲˯\~~~z��4ӆ�'D�Y�����8�H&iUiVQ=���/F��~�˿�0D�t��>�W�e~��a�u��\�ss.󸖱�X�q��}�4o�O���F�9QI��>�ɐ����M�=_6BgVv�ڣ�p!Xk8j�X����G�C��>��x/�9D��ߏ��+��=;���@���{���Tj�~iu��&<z��X��1�I�	{��E��gݟ}<<t��~�LH4�NP�>6|x��R{�n�����y-0r},��}��EQ�M���v1�ˎG�c�ꙍ��1���gp������DI.嶌.�Ha�W=Gh������~�r�E����vAǛ{��2y�����ڼ,q��#a��4D���]����?W�n�;�^)����Z����Jr1��~����#8~��ÆS��m���ADӅ0�~�:`"A��pҍ:'���=u�ӅSRw�{����T��mtj�O3sj�W��Ʀ�X�c-��@F\�9���MKG[�B6�Q��J�i*}r��&,7r� B_�������y4��Jt_s���T�)�n�wž�틓�!����";ɇ��0�j����߻8�$Z�2j�W������&�Dc�皍�y�.1׭0�=�a朊�L~���\�b?+o1�2�^ˣ{����֎WGk��O\W9ۅW�������O
��Q꺅��>���|��`�:Yၿ����h;��������#��L�Z���}��*�rV�,�!��H���å4�<t�D�4ӆ�4�K4�g��Ș�&�R�bĦ2U��-c���*�UQQ�����o��F�tY��~נ��<p�h�Y�ˣ�@�~!���ާ��O
J�y��z���i�Ǐ�i�ϗ����e�72�C��o�����,dq�9$��v���7����٧LL�Og�b�>录��U8�/�lq�����0�7q�������%lp��	��~6L4C����"x�!<p���t�$����i��	�	�$iF�$B24��I�'��JG�	�Y'�ě	g�'���=/�_���|l�x��ţ��<H��xx�=�<><l�'���F�D�<C��d�!�'�l@�SD��C'�O�'�!������tl�&��	��A�a<'��c�#�G���~0�|O���<~=o�����G�:x���d���:J��ţӇ�������'�G������������~_����dN-�,���ؐ� ���i�hI4��iÝ4�0Ҭ�p�tM)4Ҵ�R0�#K�'�z=��^�n�N?o�_^i9:���a����Wy�7�wM�MF�RO�p�۷o���ϗ�Р���gf����Y�����*os�����U9O�^���n
r{S���Fy�����^>ԯ3/��.�K1��7+o!`��~����z�*��\�s�_}��T���eA�z�w0� �����ۙ����aU\�����ݕU�������U\�������%Y�i��:`"@�<a�>6|x��yR*�!{:H�Gգ��å�Щ�!�h�y�NGt���,������l����V�?,<w�K ~�&���s.�&d���$�g��5e2������,�l�װ�+�R��¸��,�uq��}��|U:je���d�/���o���5TQg4�4�O, M4�:'���(�x�
$�L��ս�G�+�*��j�L6���A�͞���Y(��+�d�=2�'��d�0�f/���̑20�d:ph�̣(��՞�(�c"Y������@:��$��Ӂ�re����r�!��r��������t~&�����|���?T�Ѹ8ec�?Qo�߁L!�6]K9|�L͙Ƕ��e��Ҿp��,L?:X"@�i�NtO_��w�"����3
���yd|6QB�5>ۙ%X�o�!��]�G/�ƈU��NW�˯+����X�>5zjBr�����hʅ�*~�%���#L��YR�k��Th�6󓞚�Okwxq��v[g:�o��>�f"s9V�<.�L}$�3����V�O�y��8��Jv7�0�mR����A/="FN�>>;Y�7S�����yV���T�0��vw��a��r�4{7.[r8�d�m=�n,���/�|��>4~�G5�H�����ع�SĒ�ۥ����	��ϵ�{��
k���hƓ����a���4�O, M4�:'����7k���*�!�4C��^d��j�F��﯉$��_vW����a�ŕ����q�b�JM4@����?���:}��}6ڕU,��[���8���1�y1|[KB!JY]ER�F�o�oߗ����yo<�VOѶgx���KV��,���h�q�i�V��v�F&dۮ����^<|�n��W��pӆ��if�]��	��(�Wf~�0��UD=Bl�h��z��Ԍ1}��کZ����n2W�0vbL4�:\Og1|��G�z�ْ��.�]TE�[�̑ɔ�e3le��mܛ��y���ߕ�~�F�y�l�����L<CG�8:�"'�\axp2�k�,�(��GuF�h9��������њ�F�A��*��C��ߪ����<~q�O^�4ӆ�4OK4õ�W�ELO�4�E䨖�Y���!�!�Ҟ4ۮI����)YY8�&=�o"̭�Ѭ����1����RL���IB��w�F�� 'M�%J��5A����\��$W�z����.3�bJ¸��i_��G��eOЕ�+D�f�U]7�O�}.�ܖ��M�8�M��YSS��9�ve��x��v7)�0|�1���؉8Q��x�i�	gKHǌ<a��fϏ<[�v���e�2�H䂲���"d�f�&l�<����깜���\�W��U�l���Xԉ�ܪb�r-u���X�V��� !(�t^7����r_q0���kՃ霛' �����8�yͲbݳE�f��g������yP�v��:�����jw�Xpj��u�3GZa��qq���Y�R�����_x�C���˕>=FG�f��#�O�%�2�G�g?���߇�0;�D��O�܍W
���L09D!�;k,!�d,.�%3=h�~K��Ȧ��BÜ��--�R�k���=,e�#�O�^��k��j������d-8~4C��	���Y���Np�<x�������]2��m1�,����a�ٗ1�Y1IV� $/�O�>^P���L)7�����-r�D%^0s���̦����u��Yb)g��.��W橣�5��$6y!����]6V��F��Q��a��V^�#	+-�W$������>�8��|-K�:��2��r�H׾�p����ϰ�xј�1���~q�^�x���H4�����1٢'�8F���j�������1���~��2�~�Ҭ�bŵO��6���{4�+/L�ߵj6���{W���W��;����a��������X̲Y��������'��uX|j���*}2�_�s�߻��q�=��Y��OD�`5�}���G��U~�$m=5*��+�۪��Y�:�q���}���O�~>8���wta�|+��>d��4�Ǐ�Ǐ���<~u�O^��4�t�Y�LܔE��9Q1!2�A�UUO�uX�Ѱ8x�a�!�,��a�@��oq܈���b�2\>̻��.�+��wGc�X8m��ҿyo���Y�y?F=�q����0����E�ɸ&�H��t�,z�Ѡ��>LO	0��]|X`!�%k�tF��fN1<���G��+���3���CGM�~6M&%��g�#�<D�6C����h���~8O����yS
H4�(�I&���1��p�8O$6M�`���?�~/��8~:g����:�0�0��O�'�����g��8{˟��4D����vY�p��ĭ���C�����W�<O�,�./'�'�'����6l�~&�G�����x��v�zI��Ѳ�o����|O��|z?���?��ö��8v>!��~6N/�����Z�|v����'c��z>'����tx��:%��<>������t����a	����OEO��GK�־4O"Y���0�JM%4JЄ�0� ���#��[�j���h��^��yn9Ҹ�~��h]>�)nY���'����7�{%�`S�xf8�d�k|k�L[�NEqrK�/}{�ýY��p���nTӒ51�sJUf7=���&e��[X��b���=px��t|�Dۯx�0M��y:�84����9�]�:�һ��S�/W7�[qe}���E�����N�<e5i�Y���͹uw�~���b��S+]��'N]7,0}r9'^Gq�;�V��Q���Ӱ�\�y�E+�7!<�
�[�c��+��l��$�ex�;�ǫb��/ݼ\��w+B�;=�f]��^�i�����v���Ч�ź�ٹ�wu��pW�1]N�t}uq��5�ڍ�?��ܜ��>��)!�
!��h�&�n�Yjt�6��C
�4ܷ�1f�©U!�q�Z�A�jd�o$@Y+ev'h�,dM�`R����Zm[>z�<�O�˒�&Ռ�a�>�"0m��c-�m�i�r�\�FZ�E��,C��eUp����	km��/�.{=�����ffg�ݕU̽������W2�337wv�\�����ސi㆖"`�t�D�Np�:xM,�~ٹ9GyU܎X�_����K]�+��	]�q��,���V����a�v�O��U`|�m�j�M��vB4�!BF�F�e��d�*Ȅ҄���v��K��+�qmEdl��F1?���B�#yB;d�:!�VȜ���l�V؉����@���8�O�lD�����26򨤠��n�*W"�4�;ad�hn��ybcg�52<� ����7�pof^��/٠�<~3��>�-���d����t��0��7���������9>�ɷ��1x�ekfS9>w��']�t�Y$�10�����׻G��o��bz��y���]e�S�J��(~�a� &����tex��=n�\������66�)��Ʌ,�%mr��C�2>�a���A\Ww���k�T퉑
�}�fK[�ƾ����|���'�c��-ag㱈�f=�h���q��_�V_��?�?t�D���N'�8x�.�3&$oj��t�Q�Z��m�+&�4Z\,�EjU1Dmf��^���+^�gWtJ> ���8�g��Y��Wz��lᱟ�c!�L��h�F�!����%���%������Ц4'\'ֻﺾӞ\�^NM(����'dþ�+NG���r�~!��3�7��鮷�[���^:ۏ_�?:۠�&�4�xK4�L<EIs�)>�˳Z�UU���V��x��OkRO�ٰkTl�0<x�	�e��O,��n�Dw��]�m�GNUA؄?�����:1dW/���Lo)�K� X�)����2CY����T0�������{>|�o�i�^��c�Z�v=��Z瑳��+�E�UO�Qܕ�[9*�抮tt|9UҡN+�R���4�֟�z�����gKH(�N'����b��4����Ň���%�Ϛl��k�M'�a�a�����kԞ��-"�-���xժo��_P���:��~Y��{�4����X��F�T��3&c��N�%�?g���am�/*�~7Rp���U��]K>4Y���I6hר���%?N2�~�q4�Y)ɑ��i�W����0�a��ʲ��,Yx��D�?t�D��4�xOZ��ں�K�#LM���g$��TC���,��XA6�NY��2-$iٕt������V�"�����mRԎU�2�f� BY���?{,��l���4�u~G���f3�G�{�w�~�p�lQʱ�;8�rU��}��>���~$��f]ۖ?r��J�(L��D��Z8l�'�����-��F��_0�V/���OV�BV�H�� ���k��]2���<a��z�#���bg&�ˑ�ѓ�N5ƣq�fo����� �.�q���nV1#!U}BpD?WZR�8��DU*�h|�jV��w
���&��YGO�<Y�����Ζ�"Q��4M�<p�=ꑵ��m�u�UDO�(W�Z����3��A�7��+��<W��w-u�7����/ƵF���ե\0�4~��b��6�����Q��,�^�������-JhJl�����(��dc��}����A��.�v�[(��,�M���ɣF�H�ч��~�n)꼖4}Xm�-U�3�m��~??�ŝ, D�M8h�>6x���V7�30����V�H�V�d�UUk�z��W���ʝ����^,���g8@C?U�8x����{s�9[��`v���_���Af�3]����fCF�]S�c\�e���WSՎ��`�0�,F�̲�c�;o#��NF_b!��iQ��7BTO����!e�ZR̪�K�߲�����bx�e,���:X"@�Bi�D�4�M�4I�õ�f{]�����TA����3{�C�����RW�My5�b����N����ex�hGNe�ut�NQ���,D%<a^��w/t'�����C���F;BpC�hNw�d�J?%}ճuǱ�MI<nZ����.,�f-����}��d٨������X���l�F�&�-��c&�0�����\�:��L\N2�Ǯ>~x���=$�&�4O	�K4�V��+���W&&�)P�,�B�n�!L����겾U���մ��^f׫D&X�Y�~��`D�mW UTD����$���M�0�� �}���W���I˒X�w�ì��x�vj�ǆ��;w���o5��z-��G��(�0�>��c��snF�q��
�V\��ی�G��y^4t=T��K7F9�MȾ˨�j�؟V�r�+�d�h�X�3>|�|�ƙ6S�r�g�0S�f#1�m�4�}�����]���пJؘ]7E�_O�}~�ވ��ܶS&m�D[������Kӑr��F�����a��?��"d�(��l9�>���	Ӈ��0��, D�4�xN�Y���� 1m�Q��|���E�c9(�j@v�-ꪢh��5�}G	��,<B�1�>�ʺ;D v�ƍHB�����6&u�S�a0��Q�0�ݹ��Ѯe�M�&'��bǻi�Ȫy���99p2�.���D��-z��>�v�ex��X,q��j���M�J�V����:m����c�0�U�b�8Xa�Κ0�ΐ�����&	Б<"X�&`�&
,N�b`�:`�:ID""%�,M4�ΚiD�Q����"Qb'DJ�0��'^���*���f�Uh�HD���"H���<"%	�A,�8'N��4�M4�M0���b`�tK�����x�ӂ��'�ZE�"ag�a$H�p� �<I�8"xN��	b&�`�	g��wʝ����*:e7��>�5ϡ�+=K���z�_rN�ɘOX���ٜ�Ϧr>����rb.�Ӽܣ��G���Yy��|j8�,�s�5�z\M�ϙ��E�Yt>��=�$�y�͂�5y�}�v����粒��7�'3���1�z9D�ϹҚ.se�|���\ ���k�œ����1���B����~N�b�n�Kɋ�|㙹�������f�ff��ҫ��������U��������8if��Y��JN'��㇏�;M�UQWP=��b'(�:�VUA�&����9H�FQ��=<���ڶM�γ�3��cOc���8$Vp��ea�=]�`v��ڐ���f[x6}G��7U����C��3ˡ�3����]�W�Y��4a�U!��i++(a�����.���9A\��V���"��q����񑈞y{f1�ZvV���G�ǝ��!���<&4����JN'�饚'��r���}$}\�s.ȗu�UD�O$t	}�2B�O��a
� �N��*�O�G�V�@n[X�,��~�X�5�2|�䵚��1�Ǌ���7+1T�s����l{o0����3`��e���>��[baLn-�ګ�����^�kV�"�0z����Q���Vժ��1�cЮEd���,6I9iQ�艆�:x D�4�xM<Y��뙞Au\���vԮ����n,[Ѽ�s�f�ӶGeUbo7s-ٛT2�@+w1��IlWb찶6Y>�M�q�΀ ���u蜳I�m�R�U���ܜӫ4WV0���|g0�qf��W31��Y��s�8#�8�5�[��֮s���M��,h�U,�8��z���]x��Ȕ�j����~q狨����6��ku�ʅ`��
�V]B�����,O�N���U�#l�׌6v��r~ǆ|t�4)�d����������X�_��UVF�֡�S�*�y���p4Y����`4b|JH�'�����񆉇�Ξ D�4�xM<Y�߮�f`����NvTA��}�vK�V�ʕ(�c'M�$b��r���.�Qɱ�t�R5��Ėxw_Kp�H��k�T���eT�Xy}V�]8��b'<s!=8j�ц����I�#U���LŘ,w%�o9���n*�Z�y516���0�'��,��U��ҦJkߖ��+gу^է������G�+N�uǯ��,��! D�?4O	��4x�TW�J26��
A�+�,�ͪ�!���I�:$/|�r2�l�5��.��5F�D�>!�|�.�r��Ά�f��E���P�ec��̟����kJ|X��t�]MG	�h�����d���5�$cmsttH��7F����z�9Z9��l���<+!4h����3|ߍc��]U?=�Ǒ����/�u�^�~a��<"@�BQ���,�n�-���[.�MmUQ����ĕ�֍�\���r/�j�O���5H�>��٠�O	��L̲�0�3*�]ʼ�R�	����	�r�~�(���}�ٿ��õ�a�Uaʄ00�~���|����5u~��Xg�a<s�~��}mO�1���^5����$0��&iҎ'��ŝđ��M,��N;�A3}�(�0�s`n*!*AL������Ҋ��f�܄�m��9��9��y3S���o#b�(�JF�
�պԨn5%RV0���T��?  ������W|y��W��D�������/{ُ��N"G㏛������������mkA�8��;�l7G�VQ�o;U��d!�o�	"�0��::CA�:7��d�,w[���+����%�T�G5�2��4C\,6{�Z�p��gO�w�-��]��VH6[-Ktn�U�*���� �$����pi��ab~ŝđ���%�Y�J���l�)�l�MmUQ�ח�Y�,m��|�{<f��?o6�z��X�$ϫ1�j�l�#�Zx�1������~r�2{�<q��?<ǼiAF�	��W��7�R���i�b�0����-|�m���5s�n�Y�{����%��p֏�;_	�,�M0K:%�"%	Bh���:^�?Zͩsچ⪢D0i�.��tM�'�5_fv۲�4F�|�>�O�>|��˹�x��O_���3��ӹ��RO��074E�d���n qGV��FH�}������O�ߣ����=[myf��O����T��7���Յ�@J+�a�wXq��0Y����c�<��~�ed���\�:iӧ�L?tKDJ���,�ǼWd����9ɢf9�rBL�zUTA�r>Y=�;E�Q�f��a񔔖��ֱ��yt�b���Ǆ�L�V�8�g�{���x�u2u����mˆX`�<�Ѩ��������e�<YZm����'8��<j�ߏ���Y���Bտ����$�>��>U5�Q�J:z��O|ӭ+/�+�����z%���%��&$	��(�(K���#�t���"""%�"Q�I"�I��8i�M4D�ŉ�PpHHN'C�ӄp8 �It�$I�X�"t�DI,N	ӂ'�M0�DM4�L4��,�0L8%�bX�&X�Yç
:'�L8Bag�&I"I�DH���D%	�xO�X��0C��O
�I����V�E�>�vr�������Ø<6G�K�j7N�׮�w���I=������l��(�9yG�ւ��Q�'w�1���os��)�r4��U̧�Û��r>���-,^�Lkx4ݞo2(#�{qu�F�L��p��mN��rb�b#^�W:v^'�ݼ�b���N�#5��ѧ^�����Y��^�\R����K���3��s��<fI�"Hf�E��:�����=^ڵ���j<��/���X��q�f7���"x���;�p:�!�b���2�6�/g�L�ϖ�ng#�6�b�wݢ�S�4lF��M���kt�S�ս�]��	�Ͳ�;�Y^�J�njc��V�UX��+�q6HX/nlܢkZ�+��WJ���j�OAb*e��ƊYZ�YI#�r�E#R���Uزѩ��T��k#ݑ3�/�XI$��(��N�+{���oiy����X�dQV'~Q�Ӷ$(�Z��-��2;5f���D�L����{���wwwx���������U��������*�f^�f���&�i�4�K:%�"%	Bh�f�i����rH�"J��ev5d��Z�%eU����[ͥkM�:Կ��CLѤ�mX�I~�QZ9�v�V|���婫\PQ���$�i�FQHڈ@�!����"��&Ԋ�H�l숌!�Q%UQAD��I\d�+aXYP��K>m�O�H,fB*���"N7(؛v�1�Ӳ����:�*>R��FT)Zh URV�U�j�+n�DӬ��D�+�cJ�Up�G-nh H�ox���1��<m��?��3�
,���ǵTr�'L㺟
�^�	W8߸ZN�ZЊx�	ʺ��>o�8e1������p���c�=�6tk��79.�����thH�Qg�������j��zb���a�g�j��FY��<Y_ih_�l?a���r*;�X�d˒b�1�ƙQEϽ��[=��X0��a&v�cN�O6���tKDJ���,��t�� ����_��nFȞ  �J�e�Jh.����ZIzs�~�����vD�\�~=n\\<���8r��?b��2e��l>���_���n��J6��{z��=в����5�h�6[z۫1��+rZJ��	-�DU��qa?ʅ�Y$��U�>,���?pN?W�a��u5$ؚ���gҷZh�=�Q�	��""R?�Y<"x��L?tKDJ���,�>�Dzb(�rw�Q�*� �^��9_Q�ë��qc��]ʩ����m���1�l�&~�S(���|h�����^�d��F�:&�'�D��h�ɕ�S�t�B�,g�E�c���9m^�`�K0�v+ܯ���%���ؒWO�H������:s�@�(�<X���%��t��<t���%�~����R�b�74K���ĵ�Z���UQ���BOq��ލ�%��(��&������XV��r*AV�~Q�i�bRj�����a��7G�[���\����	ev>�MM����1��X�̲�Ӄ���]G�^�o�;'�،�+jb>�>�;�s��u��G��>�՟~Ĵ���U�ƞ,��4�K�%Q�4�K4�L_�N���oٓlܳT���O5@R��6���	��f&�!e�F5�v���/�Gb��6��&��WYe��`k��՘��4�:�� �6>o�ߪ��jW1�>b��k��Y�y��Gd������O�� }��?F�q}�L�i+i�xhܔ����>�wZ��6^8|�؜$�e֨ퟙ%o�M����?4d,C����s';~�~:p���a(���1{�j�/;��(��*ܪ��"���S�-i[�Q��t<$OpzXt�0񆟌4�<"Q�p��4�N/��z�eay�L�Pp���UD>�h���?W:3ㆳq����l<G���z�nX��3/���n?n�W�[���q���+�+�������A����b	]/}n���z����y�,�a�J7��0h�T�9�2�~�4���9a�?&����?����ѭ����<�ȍ.ß�&��D��?ibxD�
0�8x��+������#�H��UD>�߲�����ؚ�>�t|﮼z�'��ُ�[�,EuM?F��$g��N��+\���V�P�!�w]��N;,ќ*�ê,B	�'T�0Ї��/�;;rY�����k��}6�U��K?V��g�O�}�?}D�"~:~?	��?'�J:Y��<x�㇎�2���mj��mS��-�oȭ%���7�a�f�~�还�
[wYw��k�̹4{�����u�2�|XYT%�#4�7�6�ŝU3�#4��T|�'ŗ\����|p>:�E�I�t��,Ѿ��A�ڲ����P�4m;��C�<�;l��2���RHri�.l�M2���=|��޽e�Θt���<��zR9�c�X-ao6(&��Epdn ؜M�j��î�]�&��>�}���9��9J�!�%��mn��\E�=N�ٱ�  ��AcA��������z���O�`.T�T����5`f'��U���x�ā��Ǐ��yiQ��͈t�ź���^�J����!�v2��B􈋮4ˋl�{�&kg���~��S����%���~e��0xx��Oj�ԟ���a���э�8���i��i&j^kWÕ���,�Te���;E�_i�,��D��:"Q�Θt���<s�KK�#�-rK7yr�����>?l��,�o�@���UU'�$��tHg��G�$~�~�-2��h�}]ź<�].�	G��Xa������L�:�r>i�|�.�g��������@�J��3ɭG�Ã�t4wʇ��7D0��=]�v���4ɔ���Ǿ�Wra[q��L,㌒���cW�>���40���4< �"P����%��"`�&%�̈�,K�<tN�$ DDDL0Hy"Q�xJ8pDO�o[w���ƍ>W�+���f͸A��$	$	��$DDD�0H� �%	B'H<"X�h���h�Yf�X�`�P�%�bX�X�,�'N��pD�0D��Y'�D�I$I N�H�$	℡�	����`�&	db:P�'��>���Dq�Nk���Ϊ��t���5�nN�{���!�6��q�m���_q�Sd���O�'"�唗���G�w���9���ﵨ�zL�|�/E�c�����i������s������K��n����2�^{82t�K8Ǹ|M��}��d[���������G�;6BF��}�_���+֍3v�x�2/n�zL��󙙛������s33s3wM�ޫ���������s33s3w��4�L4�D��4||Y�Θt���<J*� �tJ?n���Y��Gՙ�g����D�6{�����2��k�<�W��Qp�.���,�&�#;Z��Y`��+�q[����q�_��;*L˹}�a�*�W�:ѪC��$��Q��V�sthD��C"HB�+Q�~}�[V��a��qב�e��ێ<%�h�Y�DJ0�Y��i��~�W|�>�c��Ʀ4���ڦb>{��<{aN'$��I��?*�.��K�w��Nzsȁ�l�Y�+�g^O��AH��>߿�`�c[�x�l�+�3���ڂ�*]2�������3��]a���)H0�Å�������S��mxp�V;�~m�MG�=���4��}�kG'�~����Oq�_�&'��:"Q�p��4�K4�m��@��e��-�J����إ�򮢙�鑡U"o`186�1�~����c"��h"�r���WaU�� BO?�����5��󘢸�(�ן���]�f2�^�,���c���1�V݊�j�Xr��(��^�}��s�~4�$�(��1g����y�'�^s���K_O^�S���LG>������sFո��⪽�{��m}���V�t"����@⌣R���q�&�#w>����ߖ�Qg�kN���:x�����K4�Fa�4��<rk����E�(�u�Y�f����,�ϕV�;C^��a�h��!�4ْG��6J0M��4ɿů�˗]a��c*�a���f_��g������U�&#�ٸ������W	>p9��B7dV,�]�Ip���C�hO�ͩ��Oۖ��wj�Oц����NZ���!�2��o�U�!�؛,�O��:xD��:"Q�p��4�K4�4b<�,��ZӾ��"e`��n�l�:�&�0�85�,���ؘe\+��U�k�i<x�m=���܆�y2���et[���D��и�J�e^�ۍ���Y'����㳻_�o[U<�l�=V��x�n�L��	^�&t��ז#�D��ߊ:t��if�Y�DJΘt���<96i�f^2�qV�U����=��>�ݴ���]e����\B~��l���J�
���Ր�#�G)�Tv��hD�_QluU��Ϯ3�Bp�z3u�pL�P�Wk^�]�z�~;�-������J5M"Y�(���%��	����5'���q�ѣA��	�O'D�DK,�D��:"P�a�4Ӌ�������i���XY)��������k>"�S5�kͶ+�[��˩϶��K���UET�RʔOYr�|ڑ�/�kz�dȳ: M�9�d��x\9-��g@5s�����\���w���o&�L����s��c�6��M�]ѱ>�Н�U�>?f~|�P��Met������ؖ�B���X�:�eX�e>v6e[����Z����$���e/�e8z�B}���瞷��r4�x�������euS�[�Y���I��a���4Y��7��
���_������f<50N�a�&�i�D�(Æi�=]�'��h��-�UiN�.���o��Ѣl�]��eZ04&R{�~����y�n��T�G��qǱ����̪�V&�x�PҬ�<Xk>��9e�	�;}l,�K�U�,��3.X�ᣆ���Q�tM	>��ar�Չ�8M�ְ�%+(��(��Mq�ww��4x� ��"if�4J�8ag�<p���|!�s\�{�^�Lq$���ʫH�=G�+1��%X����*�޺�e�V�М��7Dڲ�Z*�,0�'N�吹h��l�ڔ~�z�D��eT!I�}�m�Y�2��'���U��{�1_��bj���UZ0�}C���>���+���c�8�ȳsד/�z���?	��?i�D�(Æi��Y��]j���i�*�"pM��MW��\V�]r����ja�{��;��ْ�2�	ch��{��J��phׇ����T�6pI[�����h��˳�]`�F�j��2�jM��ƇB$��>����sg+ ��SF�i�+��<BhL��C-���d��8X����2���|&a�	$`hX��"P�=��<'�0DD��ı0K,�,K,��:Q �$������H% �H�$�"Y��A!"IN&���A��馐A��DJ0L�D���8�|����M4�4��,�0�0�0K0�,L,�9(D����"aG��$A � BD��Q$	℡�xO�&	�a"Y��9����ro�8��)/9��O�k�k3�ΙƵ�@�9����e���ڳ֘f�eX"��Y�	�=�_d2C,���S��*��[�����.��wC3w,Y��k��1f��QL7$�c����->�8��ad\���+�bk�!�l=`c��;�**��N�&���1w���+㷷;T�ܼW��N�ۘݦ��^Y$��͏Uǆ�}��u��模���)P�-��1KM-<�.u6�j����N�q�Cy����9���f�6nG�Y��sxyn�n��N���3ve�;�\2����q=��sb��	�o(�1�$�sqK�s	�kr#�7���י9Wd�[�����N8r���P[�:�U��9Uv}]���Eĥ�9w�%$R���K,I�'P�埱�eb��%���*�t��jԢr��"��m$�2<pp`H�Q��Ė�wu�?7�d�<��"�'�w\xIkV�hш�UY�`|�P8G
��O�-�P������%�D �b���>nǒ�u=&�V���EW��mܻ���������ww{n�����������www���4��4�4D��8h�%p����,��"����5ZM�~>��J�դ����de���D*e��oִ4T����6�c�H���j��hlE��l�iR&VIb-����CA�!A2)\s��
��"7�G��"��Ǉȟ
K%UYEA��I�m�P�+����P���v9Y>LNQW]qX��S���`�#�5YUU5Ed�����O��L��q������V�$A~%��+uW�R�&�d�87Bb&414s����W���sc�;��n�Ѽ��)�"8��M���7�~��X�ry�rݣB{rw�C���ڢ����%���P����닇�ı��?I0�a�vx¢QօW��4WiѮ�pK�K�ᇫ¸&�����vz����Q�����wEˀh�|Z>S!��QҽD���gM~^�Ҳ�\2�v͙G�Zv�K�d�B��q��|��)�j�4|Y�W7�ܑ�W���4M,ӆ�BQ�,M,��<�ȧ�%"GmT���&蚥8z�E��>���9�>0�aޣk.M�GJ����>��VI�q��Zr��7�n>����a�x�2Һ�Oe�=vi��*�I�lr�:Ո�ƔU����VOh����fVQ�ݲW(�7�$���XV��f[ic^�fs+�<��&���I<i�Śi���p׬�e�Oz��ξa�U�:�3�ڪ�'��%||^
4a�����ozY��a̢�H^n�C� pN��BR?�F��5����n�l��H�[1�2c�7�n���?	e��'h�K!�T�	��O��,D��~���DP�q���BW���Bs��(ѳ�L>8QӦ�h��p�(J0ᅉ�O<t�~���8 `��m�K�^d�}UZD�	x�p0؞���_#���]�}Dcq9Xd�[3L�Q��5�}��%C�`��n�[�ld6a�%LV�Ԧ���8���p�F�'��8�&.��ά񭈈W�QtX�>?,"�yW�gֳÌM�O׍<u�DM0ӆ�BQ�,Oif����kJ!�8���6±n�)qb����d���-�G��@w�U�Q;>Ox:��<�**��P�[P��J�'�̠�7e��`��VH� �Χ����>��g������ |�d޾A֥�ް\|o�\N��.oDh�/q~<�&��5F$�<�YG*f��F�Xe�4t�J�;F�,h��T�����_�iƞ��}�����ef�m��m�e��p؞�x�ôh�r�Ҹl�;F��}�=V`�u�#'�p����8`�F�K�,�?Q�4]���N�x���DO�p�(J0å��ǎ9���wC�X�r��S\UZD�v6lف���0١��ۑ�����ڃ+��k��?�5���?x�5H��8�F��7͐H5��M8���볕��^�j6�0�\��D���(؟WV��5�����qq�1�J²Ӎ��n*�*"M#~X�>�ᅝ,�p�L4�5��=e�/6��>u��K�jʍZ��Ui��_�.�wcl�X�Xܵ��>��ӃﳇM��ʲچO�#w�Zn��(�镳	���6�!�"c?&�!�L�i�V8C0!��.��v�$���ʶ�ʮ�Ҳ�|ՏcQ���W����RR���B�P�.������lLL$�M0���L<Y��a�&�p�(J0æ	�M,�D}���n�-$��!$��6�����t���<�yҫf^ϧ\ӌ�~e�q����CVW)~�G�S������l�'\�]��ߏ��W�����򴳙�,��?-�J�퓫=�ܶr*�ܪ�n�S�{o����Wg��3�M+	����{�+o_��<�W>e�]q�����_�8i�	Ft�<i��M�&����\��]��5�Ĵ�e�����z���.��V�X���.c撵�n]��*�R2c���1;!�rf!��'�a��������ڸ�w����e���}j#�?d��Ư���������������-�q�͹�;x�|W�^�|r��u����k]˖�,����~�UV{��d���!�4x�||a����Յ�MQg�.C?`قw^Tt�)�`�e��n�Գtw�'Ｍ�v�8��Uުמ���0�|�J�S!O;�n�yrfd�C�օ���^�ѣ�{C��w��h��!
��A�?i�Ξ���~4��şt飧��8x�i�WXk��l��|����q�*����<�����8����PhK1U��6��{RF��,��ǎ�Շ�1�ͮ/�x�\�u^��a��9&�n�'�'�R���*$#�[r&G����Ē]�e}��xM��フ����a�5��/�ڄd��$5[�,D�d�����Q�;P��C�>,�I���"$�H�BX��	�,L�L L,K�3�%��<'N	�5����DI$J$�H(� �"`�e �@�A$� �?�A�������D��DDL(� D�(N�'�Dâh�i��h�if�a�aB`�abX�Y�<t�%�"x������ �A:@�@�@�(D�8P��:X� K0L�����9��t�ޗSY`̎�p��'��^�9/�Ks1�̪���.n^�!�L���司�����HZ���,Q�D�%'Z!�js8�֨	����x��^��9������]�.���۫���_o�.�2�������?w������]�rl�^�����#�|}�+|UV�aUگ��*�z���Yyqt�Ӗrk����k��V{�����O�ÿ[=��#/��痙www{�����wwww������www{�����wwww���M,�DK4ӆ�P�a�L>6x�����L4�����Tb̪�YjѢ��~{�H]�G��<YI���a�2��k��\��G�,8$������'����B�?��>rFU��T��k\�z���Nƞo��c9������'����X�q��; �'��}��dl8��
�C誈�`�a�{�������4���M(�J�0�x�K4��i�j��V�.��E�7���_���y�L��˭{>�2���D�"��AZ�cE��~�����BtB�X�Q���3�/��O��[�`���L+�]s�&.:�n���j�5S��,���g�C�^M0�*���1�?2Ԫ�H�}a�Nt4����^��t�gD��O�W�IÅ�0馚a��iF�P�a�LƚY� �D�UL�{�������߶�0D�=iY�nbŉŕB��/*i��51,�ZԒ��DQ1��T����Z�R<�jU��������ތ�ϗIUq~���-�{�~8�Q�|3;֮h�'���M��{�Q(ݶ�~BD����ÊɆ��Q_m���&`���j��4��M��*.�i������`���*B�����3{�I0M�������>%ՆU��I0Ѣ�v��	� ������/���cX��d��Z"����6��Ʉ�_,|���vd�Op���%�iF�P�a�Lƞ8x��eU<0�1%�Ż��v�����|05H��+�?
pL������$0S(Cu�N�T�S�f��YK{c'�6��`�W�q���0�V����a�_�|��rL���&�T�a�L
��ƞ������IU��r˗瑨���{�qYW�bO���L~u��_:��i�iF�a�LƚY�	�r�Lڪ�'L�8F��e��i�6z�����U	���}��p�5{����UvXxCbY�3 ������������L�%�r�,h�"���?�7�8�I��{��o��麫�@���&�h����0�g$�+j���-�v2uY8d�Y8�ЙF�5�Ѫ9+�ڲ1�ڼN���0q������i�Bx�L�4�M(Ҍ0�x�K4>�&���n�w(�o{���H�M��t���0�v2ˢ��GXbɕnf�/Ś��:��Ŗ��J5[<r�u=R[eY'[rW�\4�&��u��C�X5�w����C��wPO���蕂pо,3�CF��?�I��8tM��J=F���qS�_,s�̵n��kj�-�9:�֚z��>u�Q��iFt�<i��N_��ب�}���We�n�>�$J�m�I._�L���h�1F��㣂�Q�����> �`�M֣g|���8��nHw �����}Zp�7�\��F>�w�v�[9��um��:ua}�\c�ڬ�����9~�{��qGm��]�L�!r�Z��>�.�i���ƫG;��a�ߖ֍��Y��{��?xl8]�RA��&Wiܧ���[f1�ᓑ_5b���^���֠Y!G���RVI����˘ �����Ǖ���n���w�L(�L4�K4�M(�J4��:x����G�eF�EB�$Is��D��,���>a%��4H��8r��Y�*Q�Onmq���W���m�`��q�;��=�<}F��(ѣgh3W=~c%��̆$Ĺbeh/*ý2�G����>�0y��&�V0�^F�o��x*`��M(�"Y��iF�Q�:h��g�<nU-)hF����jBHR�cln�7K$�--\�%F�%$7��*�ǎ�ƿ���K3:u�Q��~�o���i��-�/,�ghO�2�������Z�q˼y�L��仚F�PU���5�ޘCG�*�4W̟N���U�S�4��?4�(�Q�!�~����"��k}�'>4�"�#�4��4�M(҄æxM,ӆ���">��"dV���O95.�x�3�!�	��*Q��2��yP�05�>�-�OJ��\MC2\�œ%���J�L���t��t���Ѫ;��0u��1;��d����F�����0=�?Tb��Е�ˣ7����ּ���N���|�;���$������M)ez�Z���A�l�8����3��g<���[�z>�rrN�;��BF�$&"X�]���滨̩�3.w&,[��Y��0)b"-�"E��#YE�"�Qۃ�D��D�"E�"�Q�$Y
$H�FZ$Y�2,�F�H�MD�dM�h։��"Ȉ�D�mh�"�dD[E����DYE��-�h�4E��Z",E����dr���h�!�mD"Ȉ��-�h�E��D"���2-�h�&�h�-�MD�mDȈ����4[DE�2-�"�&�mD�-�Ki%��ɒY$�"[Ki%�L�D��,�Y-�KL�Y$�D��d�ɒY&I,�,�Z8A�ZD�D�IdkK�%�K$�I2�,�,�$�F�[K"�im"X�2�ImY"ZB[L��D��i	bD��%���[$��Ki4�$I�E�i�Ȗ%�4�M-!-��-���d��Im"YM�id�m"Y&��,�m-,Ki%�Kiɒ[$�H���D��d�$�I"Y"Y"e�4��$I,K$K&X��id�Y&��Ki�,H�H��im"Y2Ĳ"Id��L�"K$�Y"[L�&��KibD�[$��m�$��4���im!#L�[Kd�i	m-�%��K�M,Kid�Ki�KibBY&KibD�2�M,Ki4���HI�!-!-���D��$�,�K$��im&�I�[H�K%��	i�-��I"Y&�$&L�Kd�����2[G	�>[8B[I���[%��K&BX�$%��d���L�X�H��%�Ķ��&�I��bM,H��m2%�Q2)�����H���I��A�g�8BLY3Dmi�&,��mdš!�����h�&k#iY3I��b&-3D�F�d�&�KCH���6�i�F֙�b�L�3���L�6�i���bĪYM�;��Up�$[D�""�hֈ�"E�dZ$H�h�d,�"�t���"ȑh�-�"�&���m,��"�!!��"ȑm""�DY�p9m,��h��g8�H�DE�DX����,DE�b"&D���mD�h��$[D�k.8n9pr�",��""�m,���h��E�H�$X�!��8$[DE�"E�H�rC�YE�h���"h�4�mE�E�"Ȳ-h�&E��-E��kh��D�2&�m5���dD[D�b5��,�s[pDZ$[DF�$Z$,��D�tC��D�"E��F�h��$H�&�#D[D�b&�4B&F�&E��b&�h���a,E�H�,�4[F�,��h��mE��DE�"�-�"ȑ#YE��&�h�-�#[DE�DL���b$[F�m�dDYY�E��$Y,��X�DE�!dDE�dH��E���$Y(��5�[DE��!b
"B�h�h��DE�dD[DE���D�"D"E�#Y-�8,��"E����""ȶ�DBкpnZ$,�h�Z$Z-�E�[DE�iȄ[D�m���mDȈ��D���""Ț-��Y�"�d[DE�M�b$Y�h��E�[DE�b-�E����ȶ��h��"�4E�D[E������De�����",E�X�"h��b&�"h���4YhY,�E�k"ȑdH���D�di�dH�"-�ȑh��H�"-ȑh�d[E�B���mȚ-�h���YE����"Ѣ-��"�"�kBȑ$Y-�Y�dD[DE�h�E�h���DE��Y��"�"��-�dH�H�$YE�dH�,�h,��E�E�"�#Z$[D��"ȑh��G.6�DY-�#Yȑh�,���#$MD�DE� �E�Mh��m��m�4["4X�2-�m"�E�[DD�Ћ��4Y��M��4Z&E��,D25��-�b$,��b4�""ȑdDL��#DYh�m-�E��,�D�"E�dXxd��'�YL=�?K�̣s鈘G'�?��v�m�+3lְ�IXt�����//���ۯ�v��x~o���#���?�z������=o�����'N��w3sh�bsOw��8mG�=~�nu�^����:/��j�?������{����c��������7��������lٿ�<~�C���oo�g�����>�f�����6l߆q2D%�������o���������N��l㌛8��L�������w�/�]i��<S�f|]Ͽ6l٣�o��'�|Q$ug��mɾn�3;�������g,��9k>ٟ����b?���A��c���^C������=X�Ǐ��rۦs�4�%�����;���8�N0.$@&�\�a$���L��Lc@�%H$f�@f�D�]l���a��M��;�q��r9�������x�1�_����ŬzY��7#aD���(�����3mF�9=o�w;{�����[vߡ��ާ���8-�ݻ>&����#��݇3G�}��?���u��vB�lٸσpi��<���}n��;��ۧ��|�r���n��x�c��w�޷��o��>��g�Χ�gV��m��"y�Y��q��Ѿ���~Ws�=��f͛7�l�w���v��C���|���s��AG�{�l�g�y��cf���͛6o�{[�f[o���>��\.\�{܎��}��������N%�!�:l}��x3`�7L�y���^�W-���or��cl�lF�C��<ۖ��>=FRΧ��)qK�C	?���Q�w��¦Vf�d�����eY�J����m��f�c����U�}/�ٶ��͛6o����:���mNz��������?g�;��n��y�rɜ�x^y�p_���m�?{|���������'��}���og�o�f���N��l����/�6�6lٳw��|���v����6��Vx�G����l�����*vg�`�ӹ��Oo�����E��9�8c�^-�nG���sɟ�������dr;����ќ�C�u�3�rt76����:��͛4ߝy��m������S��M�o��s���z�7�����m�=9��c������87N��㝍�}9�a0o�kg�ܷ�rl�v�g���wswg���͘7��7<px���q�Wï[����q�����7�+Oǜ�#F�K  �/��H�
ȁ� 