BZh91AY&SY�g����_�pyc����߰����  a� �               0   iJ (@  ( P �!^�U ٖm�YCp�@�pP�   �  >�	����9n7o\���zv�Ǯ+g��w8�=�'��r�����轏�����B�����B���;��ȠU�G�B��0oH��o��	E+�R�=y�r׬;;��=�n�y�m��owg�7�q΍�^��Ch1�݋����+�Wl�q�3���VZ.�w��ڹr��^��H���)VWx^�wn�^��^�nox�yں�)���7<��w��GP��7v���{·z�k��:�:���wzS��2Ƕ��^��e��J�7�ڻ;��]7m�\z]ޝ׻�����j�*��=�5�dZ����k>���=����Zx�k�t9�#�5�׷S��������T	@�`�뷺��y{ѻ]7Sw��z����ط9���#�=29s�A�ǽ�[�uw��]��{z/`͝����{׽��7�stwn��,D �     aT 
��� $�0  h    %ODcJR��dd� �L�1  i���D��T6�#L##�!���O"��T��i�0  �M0i�J2d�`�L�����$�4��4��ѦS)�4��o&��x�*�A1J�LLa	� 	���6���A	ADY d@�F-'Bu�%C��-���:
����1�=�
*8�&�
��>a*PJ�p�sDmo�U[�=�ij �4@��hV!	 _�ApAQ�Y�mV�"I$��������� �3��I$�I$��|�( 9�/�������÷�)\�;HL4�~��C�5�y��>��LX�ё�PΌ����]C<<L�L ig|���c:�U128Ί��ESK0<�0|�K���R&3��BGN�g�y�Bc0�<A<��"�� ������g��ť�D�����2H��JLgH��P�X���$L���p�x�L�Le���B�,�V{�Ib:Ap��Le��ȅ�d&:Ta'�JEĬ`�r�{�@��L�TxgR��2P2�D�S�u0�W�@���yP�J�YC���1ï��"�c&Ԓ1�D�HΎ<1�<4�\+(�F�c���'��H��� xt���B<�I�L���ס3��g�4�Zh�0��xD��:"���t���&�$:1��<3����t|��LD3�p�d|�!�#���1�w0�0�Ϥt��2GΧS	�2�Йm¢}P�f\B���G�Q/!t,�-"K;��z�{��W<L�a%����c�B�ǒGhb-&]�Y㴙3:[7dx�	<CXA|�0�����YP�P�N�aS�'ӧ�t\� �q����$z�1��Bs�a%�bRx�u2 ��+p���Q��``��8^'�C�q
�aY#(t$��L������W�,,e��B��ftI�ﰙі�0�å��<�Le;i�H�K��S	�1�¢N�j�1Е�:�&`�aiQ�ɗ�::�P2F<�L�EH�I�39�/��p�3�԰fAir��}�LfY���=���p�G�u8\�FBL��wdP���R^)��D��bԑ}���2�bI�+�(�p�����Н.0��e��ʶC,�,`���,m+I�*P�g�#�	�<V7�X�gG��@��*!����.��R��=�b�2�u'�]��G)��2�k�f�;L�X�2�#(��>$P���\?.I��&Ag_aAc^��Bc�2V%�;ސ��ɐ�>aE��,fC
:3�e���tD��aGo�dI���X�/&��:����:WDx��]>K!�2"�1Iz2!/+�.X�%�F(\�� c��C�(��n<>�,(�p�Ɩ0��P�1�f�.Q2���!B��r��X�c��,ir�Y��<1�!1��ĈJ���c��d��	��J�!�@�K���1�O��	LcT&2��c��3ǚ�2b!x��Bc�Q��)1��VH�8T#���@�z����8�t��:X#ǉ�G�ey1��]:\cB���5d<�YeB��!ґc],ã-�3?$�21!�����c<c�adڑ��5A#�g�2�(a�=��ÙQ��0�>&A�%���xe9P�,f9Q�0��xC�j(�FH�A� d�g�(c:3�у:�bx��x����2F8L�ã�.0`�1�|c,��2F;Lf��1�׆1u���p�c1چQ�B}]$vT1�}V1����#��\v��������0�>&2FKI?v#:�C1�F;�D�qGg:�@�(c<���xe6���E�G6��QD�3�yʉ(c/��i�C<H����ҋ7�Fh�`2��#�I,����;Lfy6t��j0d�D�:t��g�y�C,g�(c:7Ń,���(e����C��ITD�t��Dx����3�;�L~��a6A��U	��	�i���
�2�:��t����gVg,�)Jc�2ZE�ġ��(�3�7ּQژ�%/��:�GO3�����)�3Ŏ9Ta$�y	�y�>t�@�%cjI ���B��TZ��i�I�Q��1�2FI/":2F8�d#��:tgi2�xgF?'!AюWN��1��Cy*(c�Q���gEmG��t��C^ O��t��i�IcI1� |��Ȅ�'�c�\,����1:L��j�JFu�gY#���2�C$d(�@�mDd��t�c1��g�)/x|~P�v��3��:`�n#:;IQ-*IA���C!�D��p����1¡��%�F1��G��>��@�C�~L�ڲZ\|XEB�H���g�Q֒�ZD�I�v��:SH��71���"0gF1���aC<8L�I�1�$k�&�w�2�@�����d2��?qq��1�>Qc,d��Ң�#���у<�aC-�0e��e(�]#�2J �_�3��AӤ�0�� ������z<2�8�Lg�7
����W�*D��AbgIL�t���8Ȧ�Q�H�	�օ#��dAE9"
|LǊ*���*����(�u��T'Q)LCk��ӳ�I�K��Gj�2J���"FԞ p�Y$�b�=)tc�F�Z�$a�d9���%�"F:] ��^;"R,��b:2i1�:K5�.�+��:2!2FD��1��fC^N."8�~����E(E&1�,H�"b��abLc:q1�DX�X˥dęC0���:H�	�xeuI�0c���*(�����������J��֒C"���<P0�]�1�ƒc)����c��Y�Q>/e!����H<��e�S<3�A�0�*�(C��1��*���e>�f��2�f*D�C)�<t�A ΢��چ@ȶ��<y�3�=~P�X�mF鏉�E����(}IH�qs�����jH=�:1�cVA�0p�1���1�	���&3��e�����p��<�#�=)3J��kHgY�
tJ-U ��NT��S��,҆�eC��N6�b�Pt��f��#���D��s�=���EO��F�۳�@��$Vny�]�	�)�^���#���;�����'�&O�I<�vQ��>�������w���;&���]�i3'|�y-��}���'�9�_fgW�;�-��t�gm���})��Ǉ�����\�&�ֳ\�*�ӷG$��;��f�!��tfߦN�N�E���._Ư{|���,�FL�� 7r{s%ɛ�gL�l��;���n鶑g�폽�2�wdʫ�{!�k�������<�R�b���s�������K��H�:Z�d�FKț��ڱf};;ݟ��y�K�y%���?<ف��밞��Z���Yf�[�v��C|�0z�{gL#������t�'g�w�v�`��s2�'��Eu�٣/q7�����s<��3Ӵ$5ﯺe��+�p}���u��혝S {7����[��ۧ��d}��\����Yt��Q����{�����͛#3����w>�$���Z�ܘ3.��	M��e��̐�>�u�{�;b}�?wL�4����o����_V��
�7d��a�v�f��3����I���>� ޿��~!��>���2��S��?w�jo��;�]��=}�)z���4�;I<)�ό���k�;&_3<���t�2�t��t�D�哫�_d�}�wT�U۝��3��~ioR�R�~��*�o&�t}޵�̙.�M�s��q�vt�Ɂ�=�-��N�DK��o�����g"��z{Z�>�S����R�����Է��þH��M[�@��ab����m��)�MW-���l��rn(�ua}���KF�~y�ʜj)ʺ�k�M��y]��{�7�g]���2��Yr�3����7�4���:t2�r佒}iL?v�H`�N�+�Jx�{�Vv�lY��&�3ɭ�(љ&/��� 9}K����wVzn}���MȤ�zcϏw'����n3:L��7w�w|컄옱�>nnV���nn�u>;�d�u��GZ��Y����������;�~j}�9�0Ž�{&��[�'�e��ɍ���g����$�p�/�u�g@��+O1o��^K�vK]WU}<�r��VǕ>�J����E]F��+w'�V>䒽�龞_G?OC���p�|6��i)���w8gwfٻ����q`s_���+W���e%o���-p^����y�;��t�
N��aۙ�����<�u�Μ[�y�p��|���ðk��}��:���~�L���I1+J�|�f�HC���.��Q�se�5�Wci�K ��HW�?��M�l
Y>T��z��3p����n�29N�չ��a;z�g!�;��ϼye�S�w��UU�L��{
:�>��n��~�f=�I��{�ﮓ�5�0p�\�Ǫ��H��V34Kf�>��/�ny����z�99� ���npl�lx;�����Oñ޼yg�*�~��e)�����F?d�fG�(�;7Om����)M�Ys�¶�l�CH2�!����O�/�d)���<�'-�;������ub�o��þE�}�wa��g����yܶ�����w/s��;�� ��&�Z"zzuf����o�}�>�fd;n�LY���w�}�Ť��ǮJ�c�{wX��+��'�v�8%�>۾�[������vy?w��tX]zǳ%�>݌��>����}?Od&��4��~�d3<���ޏ�;�ɒ{~o~�ޗBx[`�t��c.�LZk��~y�����c5��O���0>�;�y���q���m��$0�Ӿ�v2I$�߼_hY�ӧ^;�����*S��`d|��� ���ޏ�a��o�&O���̙$�Hn����yT�a�n���Ѫ��zP��yִ��1��fL:w�=��O7�ѝ��y�O�����؞����<��]��څ��G�̞����O�3X�eLϐ�&�{ض���;�������������M��fy��y!�F���4�!=_;�{d=�!��㿏�~N�c�]!|�vWC���������c{�:�����h���.N�����Ù�}�����o�'��M򛲫se��P���n'ާ��ܙ<�Ӥ�.b�������~܃�C�{������q�9{+��϶q�����=�5���yl��͚�3�ə�~�e�����Y��%�n���g��ޚ�T���!�;ٗe{'G�ݑ�=<~�M�/.~~�DGʗ��>��+��OBլ˞��(~�1�2`�l���^������K>}����;b����!���R@�CLyd��^c�o2��W�F��nl���[s0�l)v�?��糲v].[3��t6�l�d٘�o�'�gO�m3ft�)������E�c�y3�� 3CI�*y�e18 ��vn��t����a�L:�Y/�^�A���ݏhq_/�+45?-����$�n/.��$��z�������̲��h���O����P�Xi�O������a�o�s2l�����
y�wŋ�p���L)�����gG���c�:x�hc�߇���v�xԝ1b�Ɪ�i��W�D��g��yy��0�}���&��Q��&I�����?'�I�d�� h~�`S���NW���}�'s��(Ȝ���I��nH����T�Jr��T�K���l}5����˓�voxNӷ�����4<g�IBn��\^��Y4;�n�d�3q'�r�.`������O�ܞ����,��æe�ۓ�/���w&}�؜���3�5y؜f�ûV2��l�:�,��d>�=�M�q{m�m��K�Ʌ���ɝ��a���w�� �6^�v��f�}�d��-����rO��|�3��w����3-v̛7����!����7�7�?g��/K�g��W��z���.|�j/%o�Z�O�r�˫WV%�2��?�v}$��<O>���ut�T��;$�&������Ҝ�获�
g�_	����;��fI!�s�b����v�N�s�:�O7���鯯!dc�}���u�g�v}�a�z��$O����U];������U�N�:UV}߷zm+c�ow#����B��{�/�!�Y���~팿���ل=��$�,�d�aѝ=��Au��Nl���%ޝ��	�7�����]�+�_92ffjkB���A��ޝz}݉������_�^��xk�Y�}��7�t����i���+g-'�B�<|%@��	�%�4��R��`��{`s����GXsn�K;F1bpj�3���n��&&P�Z���2�ɥ6f�A5.M���K%^� �ͱ#�ܝ�H�`ƛ˴�e��XٴM����#sr���f��n& �[��mةX"�˥�5k+���:�&��̽k*�Ζ^�5s,��%q6૿�.<�RL�<.�5��(�Wt����tK���x��"v��UTp9k���I͵�Y���,�G
���@'k^U�"�4���Dɍ+�B��Й%�����nv�t��~z�{��{�|6�M�έ.˰KX��Ou�z%r:cf]�`i��gkZ۪-9��U%��Y�y���o��$_w������K�u��Jj�v��y÷�o4?���'�S�o�n�ڱ&k.�X͵��7:�օ����Jji�V�v���=hEm�@c�Q�v^�%�E{�g<�����|=+!kt�4��Զ�$5�M�R����2v.繱S��N)	F�R��)^�8�8�S�>o{��G��(�VX��������:8��'%T�Lq8�)l�K�Qz���~�� 	~�~��>�R��N���.�+t�;6_�����b�[h�&Y�#X��z�@%�����3@`C:Κ�{l�uմ��鴥��\�a$c���"0*��xSn���7���a2(�qU��V}���'��.�(,�e3�����w�SǶl�Fn �� �`�$D�d8����S�̲Jt���Nt�cn��!�J�l��=8��ѝ�����ɼ/C2�9W����p�5��^e�Ĭ���IRO%;�l�k�.��nl�I��$��i�/#s�HcpM�8�aP���Qzrr�"s���ĥm�;�J_j]�Χ������ZJ$�q[G�h���F�v^��á�
^��c��`���lϩv�!P�d�SS1Y)��ۿN);�H$�G��
pp^�&�.��<�qآ�,����|bg�{<ʲNT�k�u��؎d��ےs>�����IF�j�1L[޾�G$pb����(��]n��sr��k14����h�&H��4�f�9�fx��m|@��[�
�=UtPU�kIo�o���k/Y30���?�$z:dOO�@�ߐ��_M��$0��� 	�{�;���( y?'F����=�ϥÀd	A	 H�IdU�FDBD6����Վ9p�n����W/{��6�~lo��m�ݱ��m�6�m�p�o����m���6�~����m�i��o�m�m�m�m�Lm��6���m��������.��p8(���"�$� "��� K�8q��Sm���ۆ�m�m�M�m���~m�m���m��m�6�[n[m�m�m�W��6�[n[m�cm��lm���}m�m��!��m�y{��� cP�E��Bas��pH8	�pr�O6�nۆ�}m���m��i��tۖ�oͷ�ۖ�n��m�m�m6�6�m����nۆ�oͷ��6�n�M�����ۦ6�m��m�G8�8%�8���;��Kw[m��m�M�m�m�鍶�om�۶���m���۶6�m�i��tUUU6�m��m���}m�m��&�oͷ��6�w����{�(�	IEdY$FAT	��`��J�� 8E� n7i�x��(�����BB{�������#w~�t���!E%�1:$�-֙u�]i֜GO�3`����xg�'�@Βx��"0c��$c�1�3C,��3X�(e���x�Ė0���1���@�"@�!��������t��Qպ�GN��&Zi:0ac�2F1�c0f�0`�!���Yьe��a#�1���X�&3	�0��Yc%�@�c�3�:ӭ��:㏛u�Js��k�y�
�� %?��lZMg-��J-)���|�χt�R��f���u�O޶$��_L�6��v���)��zzY���ڦ֮�{2�$"��ڱrv�m�0
iD�5]v]�����aiv�f�s�Zkwb��\��(ٵ����]km���:)kHX��u�3B1��/��6놸�b���a�����ѩ}(K
�g;SG����IH�9�C[j[�؟�)��XԀӓ`�$H��hi���6�niq��a�Z�hp��E���~�g�jP�)4Z8��l�`
TѸƔ�m��Mf(ؙ�}�%=*;]��"�,�f��m�@�V٭�,��L�{ �!�í	QE(�ŏ6��M�%�͔�n�)�5 �C��%�̯iJ�5���Xov!�imɬ�۵���[n�f�[{,m��	�X�Fe���]���V���e��+U%�:]HE`�4���8�a5W�s�4�$%�m�&�V���t�hͦ�a�&)�J����vpr�,�7M��x��%�%l�-����e�Km6�-<���I�M{�;mԱc�7.Ui�#32�,)�8H4TZm�P��4v�I��Lخ������y��������Av�;2��iI��Rm����
SV�s��h.Ҥ�,s��e>gA���j��mu��s�j]�f�W��VWkZݐR6�e��W�ҷ��m����I��u�Z������g���YC�j�mC��H��h\&�ۍҙ�5$�ݴ+�sr�,��ͩ�]�H)�E��b�پXԾ��"ғu&.�3K5!�	u�k�LVbcM�ٹ+�9��.��2�feu4������YC�hV iL�\m���:��\�A3��)k���7�j\ݨ���K썕��f�]�l��\@��-�c���R%���m���X;L�(��噌/T��F@����+�׬��t���@������$���u�WB�m��~��)
G��s�t�:���JL�8s�����n����x �n���m���h�pz�wwv���s�����������9��9�B�4�Fif1�YC(c$d�a��{�}Y�y�6�i�pEnV���
�̴�&)-� �]��Zb�L��XÒ�%�m�Ƭ�mTv��b�%�)E\��P�]���3���q��l�Ĭ-��֑���M���I���wfZ��Dus�wf�k��x���	�p��f���3G�U#7V0�n�Z����憫����+���_zY}e�!��%��!qpJ{�O彩��z�=�*mV�|q$E�Z������&V�̎V��a߃��������C��;�s�&}�.e2����/A��a4z6��(��uT�a���S��=���=)�sq����
��7P/��A���#��ZV��ag�4�Ɵ<��,��3(ed��<a�U�a%ǂC���ɺh�y��w�P��4�ڝ�D����;۴����SMG��2M,6l��Ӡ��Ԛ*�lae�_�YVl퍻�k^����ٵ>�u͛g�b�����.�m��)�:�&�u��f1�YC(c$d�a�ʑ�(`WEu)�n.�Y"����H�#v֋�RwKB��#��l�?�\��g]"A�	eJ�.t0`��S���_i�c\<�,�����dd�!�p���N�>��۸ma�d��OO!�SҸ�/�;M�}Y][���-��HYҋ0c,��3(ed��8xi��D�b�0D�2���
%�#lP����o�F���3.�f�]k��΍!Jv!C�S�OI+m��].���8�g��Y+��"1O���n���r���c�)�!gQ��M%�rEe���I)�&�:��Tx���F�|��1�Y�1�2L0�U�L��[�s���W��yb�9-%��FM�m������h�nU�'d�&,T�9��n����ɮW�)�]C��lM6�4`S)��*f�J�u'�����I-��f�]��P��6�H�	s	�j���mX|�ٮ�6�uR�t�aOO�F��1���)�Ⱥ�S睧ڦ�y&*ZJ`�2�0�NԺ�}Lײ���JE����>=��K��r�<�XN&A��ڱ�p����0�	ã����[�m�ɶ[q�θ�:����H�0��f#�%3��� �ag�U�;��z^��S	�y�rrw�32�ԡ�|v�;��I�9:�t���T�;�����">���,��֦�j�$ZS7u1S��x'ofV�i�{7�K����2�b�yE�գ�Tw)}��_Uu�i�[8��u�u�\|ӭ:���8��:�k2���������NA0:�by�#��i�]VXF��8�Ho�r'��\I<H�{]jf�EڷMͬ��ճ��FXzi��Q��%&v)�����b�F
�|�Ú�1V���S�3�_|��9��Q�ӈh��1�P�m�~�lK��P9��Z�U�%����}����Ð����v>�VU�|��,��]y�q�q���&x��q��Om%Q-]�i+���Hh�MP��d���Ț,L5�h�fdt�N�N�ؓ��{�����V�����;�P��z�L'�];K3H�)�'��/�	><��2�딱׹O;�K�rb�L��ɦ+NS�m֏�i��u��,�Όd��<`�vwR���#.cױ���ql����f��8-�81A��I�5W�ץ��)��_����5�g+j�)�wɕ�X��R8��E&���Pҩ0$l���UTf^[�RY�n����	��=ҽ��8���3˥ͬV_*i��foIW�Qk�M~E���N�0�๻�g����ʸxR���eQ>qĚ���y���&d��>���9�������a�tXpO�vs(ܹm\�� td=;�i>'���&0�S�.��PL�`����0�61���i�"��R�)��� 4�,�L0c��u�]a�q���8��F�����Rҭ�(i�rRA�ϧȳ��)�?yx��==׼̹fhQ��n/�Rv%zO��d��C��7jբ*Ֆ��+Uv��=M5�U�*����q�>;!���z�]۽�m��w�즋�{^J�+�z�Z�a~L"�]��'�'�ȶM&��H��iF���Y���#D�!�F�L#L�P��J�~����/�#���_1���YY?���o0�/����F��h�Z2$L����DC�F�F��0�4����/�/��+�/by~yo'�q�p�L0�2�-�O-yy~i~y�O>�����y8�x��"�O-v�Ɩ��(�4h�|T~�zKF���/�o///��y~OI���X��(�����'���{t��߅�g��*4dɤ�4Zi�pZ24��Eѐ�!�F��F@��4�4ax�"�LDh��ei4�,�.���G*�e��b���?f[_ɵӒ�!�B^�c�_Eȳ��M[���W�`v z��\23��ß�\ӿǿe�����t������̻��n�����333/8n���������gOi�3L�3:i��y�^e�[u�ꝴ�H��3L�h�t�� m�ѐ��\� ލ�d�	CF@0D@ф���O�1��Q�9��A	�d��'ܼ��5�K�֝���:�٪���W;�+�zj%#t,rK�J�V�%0��M��� q�ߞѷ�'���~d'~y[G�,D�j��qJ���)O�)]*����<I:�&~_�@�"FB��J��&���3a�C��`~ZN٢v"2C�J�6�����.��G�yղ��_�y��1�Y��4�M<tfa�5Gʪ���A!�3��Q�o:^�~@XO � !;�!!�	��|���K�)���&��
ŏ��RE���X��0���6���P��(��DR�C��ED�r���pA6�l�8yݵ.$��o�!D'w�V�8�t��d;I�0Ao-MI0d됤��~?4>&kS3TB�!�ā76>������u�ۂ��tw�'�z����ZH<����ł�&FjSkdۏ<���:㮸���x�I4�ь���$u.Jk�u�{H8�0R;�	ƛ����l�.�ET�n����p�>��sa#�Y,⇄-����	�����\S��������:�r��T�3Z����� �!c���ql��$l�J�����ƹ�RZ$I�F^�����UA�ܦ��&[�^�)�9��{�u h0����r�zM����qRRъ��Z��V�îBz$�Da���C��=�)`d�N��!DF��Λ�p8r2L��=�'4�n ����4���<�qD��hM_"#le9���5NU�J.ԓ���I�d4�շ$�@$���'t�!�9d7�1$����N?�e��.�'4�35yss�of�!S0���>d�,?	<#�&C
#	�a*�LU�%Usɜ+iLS�8mƜx��a�0�4�i�C#���ʪ�",�&�&��"%IԶCE�a��iC��"c�c%M�b)��;�ѷd�"u�!�;a��p�E}��>���ʑ�P�ޭ�O,)�:�qD�Pq���B��*�~�rw����O��	��Dad��t2o��ہ�m#��]B���Sr��%8�N���i����j�xǢZ�\�3.��$�?2	紑)a�e!�Ʌ9?}�u��L�;g�	�L	"[gp@�҈���5��`��pJ���\i�����8덺���/<��2뭺����1rI$D�!4`gͽ�v"%@��х&2��AO h����B�.I��Aa���҇2�f�"DaD
��"CFHs�ÌbB�:�3���u��7*���B�;����Ԍ��'YTcs�n�L��O'r�>�	�KD��?�Iaa�"��Ԫ�Z"5���Eu���Jsd�������P��z0�|Xq��d�{l�N���8�8$=��i?A�����p@;I�!$E	Z���]%?��__����q�1�A�M4�O�.�{�b<��TDa>5��'�� p:�i<�&�'����pHbQ�Y!DD��]�z�]t�o9j^���k-mP�:@M)OŁQAd�2~��Mɐ
�D�>f�٥,��~���Gj�� �S��کa��~�|vY&���@�B�`��I}~���r���E��PB6f��N��J�rɐO�5pHVH�JP�e�M'���h���}Y��NA<��0B��2��S��a؅LAF�|i��2�4Ӧ�I�*�^�^�����������g��+s��D�1��z��$8����*�t�ɐS�8��z��#_^�騭��M"B��;+���nKHⲉ� ;�~� K������~�ゕ�����۱��ls`�'x=ɃAy�^�,��GZ���Ċ(*X~��*p�N�.�S]�ݤ���'�[IbQ�)��RON�@�ED��	�0��!D�!XB�����vw��!�	�(�,�����ᜈ|m�å�(9+��.�!�>��w�]�p��8�!rj�L�?J}]�&�;��;�y&M��W��=��w��ϗ?D��,N~���~-�O"t �=���\��9^gDu�
9�8rMF0��!����Cx��T�6U]C�r�?<���n???8덺���/<��2뭺fL���9vZQ�9ϵUQ!����Q���B�#!�pd=�l�L�DB��bԢ'�%C�������IT�Q�bd�Uz�� }|�d0Hd;I?2v�]H��	�<��C�g:4e$�����(��dAHCP3K$��@Å�a�q������C��W.��7r���N�E,aJO`��R}�pjt��7���-�Uq(�DV�J�&�O`�=,��`�w��k�b.��U��䤍EÔ�6��0g��P�4�M4�OΏO�N��UF@D22DD�Ȑ���ꓵ_��2���8��+2 ���Y`u�[!��(���OO�3v��uy�C��==� �&��ɻ���LpLHY	�	�g��j,�i�������s�sDי��Ln+�G�;d,���8rv TORA4CKIY,h�阂�����Y����V�WUƖf~K~Eq}L���!jN�g�'x4���w���'_-;�(?����%a��7<�;�lB�D�1a��~���B�h���dD��qe�JZ*�JE�y�矟��u�3M �I4�ь���I$!>����@�&9Ć� �g��4LdX�����o'W��uc;g�l)� �z����������M�^ckT�[��O���e����J��Hn��QĦ�)�0$����z3�77�VN��l'�D��`e,I��@�d� 2xz������$�!�H}��{vC��g�H\,���&��ղ}��mg�,-��G`�������D�at�Y`"��<���bh~d�(�,��dP��=9*�)I�!���hɴ����X�ML.��ii��\z������i�����H��'$�����Ѥ&a��6�M��-���//)����y0�����1�y������h�����C��A��J4��K#L#Eb���L&�B��2,�$��>>&�������>4�dZt�6&Q~'��o1�_gɴ�K�y��q��/Ǘ��/�.���&V��M������ϊ'�O�����h��4�l-#E��Vi���++��_����y�>M<����a�?�FJ>!�)i0�C�g�N%�8K#a�a��E�
�<iZ-6�N��idif��}_K�e�{?����pݧܺ�?5+�v�	��=��dR�	���r�rsxK�F�8r�
�Q�"���"6�4�L�̘<�al����m��]�-�!1����^�Y�m��٘���ۥB��3���1@S��%L*��ݫ�=~���Yl
�R�1&��h,|����̷Q�9=��\�x,X��Z~�S�Ν�^��ӻ�wj�����D��m�f�����ן�r+|#���y��>K�#d��'-k%Ƈ�ߪ���N���:�y���z������
,0�&2���GYK5�������Zz�頯�5#|��	R��W~7����U�N�*���1֢�͝aUuN�A$#)Z��U�����<L0��ݴ��D��u,�Aj�v�
�\�B��ǔ�]n7T�hS>چ���Ħ���6�Fi�Ս�]j�v[MPsI[�����t1�l��d	�QF���y˒��ljR㠌��]����GR"f;�. #�`Fa����}{�����n�����fff魶۽�����[m�{����xУM0њ`�(���F�i�N��k�.v`�Q�x����}f6�Yn5،յ���)S���Sݦ�����"��T�X�u�1��֢�1�mK���N��$n��FYS]��Yk)%��-��!����:(��C\�Nwi�gx��)v�+i&��j����VX&��o-�f"f�b�6�)qLRH4X)(�'*4ɚ���Ci����,؛d��[OB�%���S�~�  ��~͢�$U��ns����=��l"�A���M=�8�U�q�2i۫Z��M,�;�A�p�K��M�h�b�K�s�-�M��a!��a8�$"
@т!�2	G�kL|�y�{5#��nRR��.�J0��d�;��L��C޺�l!c	��"!�'PL�Xa�F2Ox?�vLM��8<�Vg�s�hKŞlcbh�d�Ru�o�>�g��D��1�����[��Wqݶ�!���uؿL��o�D)���A��GyN��QF�i�0��1i�M:tc(g�}T$V���x�����ɽ���A.N�q6D���ȫ��)a���{�:
|ak{��t0§ku���8bR:��n��3+[���F"F��_������|�%g�|�tٚj�1O��~��S�F�O�����
��$��LNy����sl���w���GL�.�<x0�Ϗ�|`�(���F�i�N������򪨆���Uާ�}Y���t�=�|�.`�E�k�r��a�:V��	�B��LN ��?goL_D�qycX��N� ���ʅ��7(���y��B��w�0��Z�$FR��=LjM��fi�mV�Q��ԬGZ�r�!���m+Hە�u��C���Jpv��H��͹�b5�jKn�Ti�����`���4����Q��4Ӧ�tc(��(��UTB�s�W��S�FE��S�9�P�����2���VnmE��3N�GUH�ŪR�z�a�����Mv��V*��Skt�R�:���ԍv���WR�L
L)�J|wG	d�3!B�3�V
�&C��G���N������O��G�b4�N�Iь��%g����ǺA1k��{�H��^f&L�L �7k1'dMS����NͰ�C��*�x�O$���Gl�{�.\�̆�'z�0�d�cM�F�o���ٲ�
l��qݨ�  ��/�m!�+��.n�2��1ʤNbmb�Vnb�k�A�7���y�[5����a�i��8s�*�y���=����0F��0i�$�3����)�-��gY�I�;�d���D�g���5Y���2�劷���˺qa��M\�k?.����\5�'��'�98�­��j�{���|`�Ƌ������1��yPb��>���O��F�}��)�ߙ�~]���<��Q��a�G�b4�N�Iь�s,�˧v���앐d���Vz/��y����X_*�!�W�$�p�Á�B�*��z(�})��v��r�~ߗ�>�~^�e�!�k
�W~�1+�)������~v�:���~��烓���ﲆ�S^3����J9����WBF��1�����+���u��ޓM�����+�s�����S�Ӈ�Gӂ��Cf���)Ќ<x&>�����DGo4A���(�F�a�1�x`�#M4餝���`���UTB�C�=\4�1�IIC�fO�s�Bt,�?raϧ��e��w��NV��Z\䥄mH[$�Uj��o�%��K�ӎ2�7�Q���ֻ��zK�)�x}0Ã ����io�7w��o {���5�磲��@e�eEx�omRA�r%�	 ��!+���6���|�k�V�Ͷ�H�굛�Ԏ�����l���^�4�r�e�a�6����u��t1���N�Iь����� R��I!s�}��}��X|?�ۅ� �GW��U�Z��jO��w2�ˣ�R��cJ�$O�u6��j��ޓ�/�FJ!�<���Q?~c��U�����䬙=L6{Y���I��u�ի�N0�z��O�M!�d����?9OԌ�~��˕�J��W�Vd��t�/.i+)��4�6�����u��:�:��/2�������I@��
�[�KQ�4'�f>���w��}�g�QD�ob�I�٦x�kZ��*��+MI[K��щu�m�� !%�+�n*u�����:�%��ޭCƴ�M.s����\���&F!�/|��Pa�E�&O|?%J��[�:?S��y�`&�"0Rv-�y1���z~ώL(~(?�\��>}[r���[h�k�%2�6q�r~�_���H�ʞ���a�:���̵U�m~��X���HMB�GP��_��t����f��8��.���4�7WO%I����i��[yu��q�[iӮ��<�̲뭾0�"��UTA�?l?I�Ȝ�:��Ж��ռ,����o�����@��$G\:-�q:�g�y_aO�E���3ϗSo6����ZζѭSH}N'�K=��4C���8�:�s#�T�5��o%#(���ϨzYx���obOO�6��y�i�}Xi�U������V��
�F	�$��u��|G����0���yv�O�" �A�QDx�I�h��	�H�H�FQ���t�4L���iP��oKyk���m��ˍ/Ǘ^�I:+�Q����dh��4L�L�#��Ţb�ѤF"�Y�-0�,�,�lT)4�T-6RF�Ӥ�%�<�y�|��G�W��X��O��s��&^_�m̵�����a�J�<�-�0����+ˬ�)Z&H�F�yq�Ǘ�5%�%���<�4�'��痄�����<�<ǓE"Ӥi��҈���O�G���4��~:i,Z,*��0��L�KL'FGE��B�H�Hp��h^ �\Zl-"M!�Ƒ��U�I�iVx���O�0ē�B�O��B",�Z��LA��C���Sq�fT�(�	�Huh6Ȱ���ē��a��I��	U�0H�!�Y��yi�t�� /̇I5��:a���@P�����Q��U�ޑQ�ygl�&���s��oi����fff�m���333wV��y{�����[m����̤i�J��i��1�x`�G^y��e�[s2I$Cշ��L����8�!ק׹🶥k��o��}L��Cz�ُ?1U�G�||��V~��B͞���Z�ؘ`DL���+�I��O(�/ny8��MV�:�$un�U�~�q�S�Uqg�z�U`��o<��1he�ϙ1N<��6��H�=Ye���矜q�G�b��4駆P�|�"8���M�z����_�}��4|w0<4��>
kS*1;�6�s*��-�ȒK0��/�>Ny�6��ڏ�'㳅�Ga�2�d�D�[m<�fV���]��.O������}�+��KQ��
,>�=�.w����|Oge��p�m�����ٟ��Y�e�ζ�o�2��θ��:���i�M:i�}��PE�OE2��O�g�P(ԱI��Ю�E*NZ}۵���Y׋/�&t��D���Chk��� '�ԕ����v��Ś�)����˱~��g�� qlX�|Z�݃�����8r�8%Ӎ��t������G�&�n�3K����Ze1�������m������Tb����C��V)�5]�����ahj��8����ܦ����ß:q5Z\[nS�|��Y���R�E��I��Q4DHF����3#��y��g�}�Τ��S�?z���./�UGi��|��~q�[iӮ��<�̼ӭ�I*�wE�,�RA�e�2�ϒF��1�B1�(DEQ@X��@U3)fZLBVI�b�T"��a*� @7�$��X(,��9�K��ם��!������ã�!�q:��F;*醇,��u;��?#�Q�!$�3��_��Og�~Ǿ��5i�`rV1Kg�n��җ,��ZJJ�.��*�~�S�����/$�`���Xծ��m�wվm���%ӀN�-�o1�Բ���w�OM�\�D���{�����9lc��9!���<M���R&�d�韛��F���>2�-FRz�ik֗ll�Ue���R7�k%�JZ�;fc� �6�JX$T� uǁRZ���jA��+NbT���C���ʖ^y应��j�J�bŊF*�X�Y�KZ%�:��5��f�+R���ç�MN��~<�{|"İ�9�ڪ������3�D֪)Ʊ��̳k"��,�
�k����Z˵�]j'�����7�Z����"����g��m�-a�x*��Xt�e�P�a��3G�b�M:iᛤD$�ޤ�HA8�̵MS�u��2hu�N�_�|���ۿ�i񄥾���#e�yz$�U%V?S46l��g��-3Kc��Iq�%�M�|�ǟQᳯ��<`_-87��.3'�tP��|����Q��#�
JU�o:˔��a{z>m�Ͷ���y�\p�<0c�4�M<3*!v6Q^RI"�ô��3��.�:���}
{1�B���ʏ�tf�CU�!L�J�
k�T���V��<-�`��N�d��L5%�����D��/�7>0�G�x��hBHJ�2�5��d��=MST��~�O��ˍ�E�*0�����sߩ��ܹ�9\B�Ur�r�i�_<�:�뎸`�<0c�4�MG||�oV�|a��WͶ[k�
4�ٲ+YcV6��;�y�Ͳ�n,7�o;M�j���rp�U�"�P��[zR�`�j>�������  �\�֭���z�I��,i�<�+P)��)���� 53Ua�3a1t�ộ�.sk�y�T+�I��U5�3��o-���W�����d�2|U\�����$c��<����JN}��+v��4�[~so<����橦�Y�n��w˸���k������0�����8��#.���"�u�^�<���i�F�Y4�7eۈl�����O۫����3O#��_>yo8��8�m8t�1�tӦ���MB�W=@�$�B��JR~2|Vʢ�_��S�7��y%�<H�y�Q��'�A�NÐOчg;��y�̇��;&�/|�3�~�kR���Eƈ�J1�ݜ�Z�bq��婯�~[Ŋ�K!β1�;򊏕xw�|0Cކg��LTY.���m��~~~q�u��:�:�̼�δä�k{UU����)�����~NPo���W2&I����&`����:���C��};M��T�f�<��N1�H[Uu���n�M����V��}��҉��&&g�Q�q�;d�Y���V�'���~���'��DV���TG��Z1*s	��arq�g7�ZC5nkW/U��O�m��G����a����0��x�c�~4�<bI$��9gy�v31���=]u��m�?�u�gM��V��13i
�N�h��ݏ׿"����k��N5X~m�u�W�ʳLb�q�q+�3m|J��c�\�޺E:4�vK'�?~>,`�GfK��0�6Y���b�T=*�G����0����v��r#����^[i�|���<��^N<�i�����oV-(�L(�K^�[-�	o.4�\y~[�|��t�TL�"�#M"��#Rd1tZ&-�04��#�V�Y�>M&�Ɨ����i�����6�lZy���<y~Z���4���ߘ�O�����r��.<�-�0i�S��5bh�ZQ�O�>;2�ZzK�-_��0�'����<���4�4��D�B4�KH�t�]#ON�l�>'���GƑ��������Ţf�i����H�!iR�r���DxZ�����`�i���p�4Z&"�Gv��M��mV1�2n��b�e��NHU��+ݞWw;m�a������[{K2��)T*-u���(袨N�Dꤷي,��>D�	e��U���n@��*p��,唼��2���c�ѕ�[.,�;��&-0Մ��-k��=i�T+.��ٜ��Kcx��¸�qͳM��Ǌ�2ٖa�K��YȈ��Uv-�
�J����gH�܁s���k�NI"t��	H��ʰ��~MM��M>V��J��jnǲ������v�H��E�X�nb���H���m���yVZǎyl2)en:�i���t�cǙ
�/��x��ל���w��&�5���l&�ܙYSo�!��_�z�J�Ky�ݥͳ3Ãj@Bۑ`�Mx�W-,�r�{@��Pv"��6�T��m�֍���h�*���4�~�']!7Q��8�kFƩe0�OBU�@��\�Ķ�^�\Y��Y̜jY+A�*U6�u��d:+�+���dhK�r�V�{��fffn���o.�337un��˽����[����s33�4�A�`�0e0�1�tӦ���܁L�t�D�OWb �l`��+3�,�i�.aa�� B�u&�%�&�h�m,�e4��[�Z�0�]K��ۖ��F�ŋaT)L��6ֵ�*�HoO�1��ɸ.x�KX�#�.�ʆ)��mc[1��E�#�&�4��0��k��W6୷��X�M�����z� İ��lF�V�T�� !)B�5����8�<>��6�̐��k*�L̂�C#��4�1��Q/��>}Ma�9K�>��+.{k���6��a�;�g&C�Pٟ��R��vv!��S������w�v�z<;��a�giC�6�ŝ��;:����ND�M��Z�_prn#���m0�~:��eyL�j��ߙ��#�8�~q���`�<`1�c4�M��ID�G�b���=F���Q��d��u��[���	�\O3�K��%ݧ\B�{���^�U������R�֔�kN���08{���]L�8hc��~��s�y�T�{����e��p�V�͇�{E�p�RS�?M�}&��iA������G��M9�}O6㏟�[�8����3N�tџ}�6e���� ���E�}e����!c���=�����#I�����]�h ��ؔ�!�fwO���p�fT^�SCC~����׎�����0�A�A4I驾�||�ح���~q�MS�1]�w�v�IO�1I�_���Nt�t&�e,z�����}���Uq^��2��u��|����q�(��!��M:h���I�l�	Ka�C=N�LS��0X�������%���A�cB�cN���\��F���Q����hw:��۞|�ە?.��i_e��_R6GO?Q[����l���xh{���s�F��R�}��"*����UUAs��i|�H�|��� 4�$�
$�>> gƌ�G�1����O�N�\��Ϙ���r��~��=��l���-�=N�R��oji��P<N��	.g�=rj��`�m���;�	�-`�$ /� BMLl��i�N�5����s;vm�.u�̗^7(\��pΏ� ��F�Y�Aŵ�����+6�����ۘI�~��Ze̘�B�5����M1ڬ>e�ںYo�o�f����e����9MW�I{0��l0;z��K�4�a��#_���R��Z������"��*fn�S���O��g�w���{3��3$�åx�F`��2�b�4Ӧ���t��I$������~��j��r�)�i��J�]/:�����)�yd<�T��̐��{Z+��$�m�1M� ��~2c*�q�W+�����+t������b��x�8�';�L#>9'r'f*S �^��w�/i���_��#���w�%�2m�v�h��㍸�_��y�m������2�e%H�-$F�H�q�Xf�M��Q#���#�1O��X
��0�'��V=�u:���zibXxa�����1�Ja׉�m�6�fk��̺ �`t��f��f��i������e�Ju�I֞�N��]p'��^;����0S�Mv'��8��a��(�,yS<^9g���Z�ov8H��fSs�W�O}�ob�mӾ$ÿR�1��6�1�Ϙm�+|�y��0��>�2�b�4�O�N�b�Ҫ��>�����*~��C���~�(��C�����+0̛�I�������z=-7Xi���eU�k��k�*~�>Z+��0b�],�\��T�Di�v��kCt�<��oG����S��hu,�A����'\>�m0y;,à�n';ٟ=��	>t����xf1�3L0e0�1�i�M^�/�Q���;��5i,ܳ����S�b�*����xLk�<�nL3u�(E*���B [�\�,q���9�N9eX{� Kq	o���" d�N۔y2,#�UK5�.͔4o^�i�{�e��[�Z�ҩ�;(%l��M��"��v�"�#̷˹v���a������6�N�>|��I޶þƘ�!�]>�`r~�,�M,���0�/f}M��4�ɚz}�Ҧ�C���DC?~G�f���Ǚs^�����cJ�>�~�p{�4d��?7�r">#�p��e�x��4њa�(��!���tљ��*�O�}?i�'6R��P�ϵF�?wܲ������m�ChH,�a��Ov�S�gYq���&���<�5�ꌛ�~�==�!�����Y�J�G�[���>�v�N�&k�']g����8�ؤC����\�wv��e�ko�Uӵ�f��-����u�|�$��ጲ�c�<1�1����mi�e�e�Z:tӠ�!�$c:`ΐP�tf�	�`�tf3�,e��GN�:1�Cє1����Ab�Όc� ����Q�Ǐ0a�Fmգ��2!�21���3!�!�c,����<1��4c4f�a�xd�3ac0e�t��X�<t`�3����e���YK߸w��NM������q8�2���bi��Mm�3��a���=n�����a=���9O>��Y"��:�s�wo=&�14pX<����&c�z]����=���>������o2�337wc[m�^�ff��km�˽��7wcu��.�3:a�J4�H4f��G�1d�Ӧ����I$��"���1&�>?SoS�4�n���fK�Y��o�)O$�O���`"!�bR�s�?�Q���-�hMN,S�ux�Y�S����H������)��	����<���Hq;6�������$�o�X�FKa��C��vS������%E,ﮗÆ���J�Yc ���a�(��!���tў�2f`�N�I$ �!eF�R�)/I����<A����T4>����w����e�&e�,�_{=�p�D;�t��~]����n7M��<�!�j9O�]Iz���U��r��$�$�=���W�p�5O��U�3�?;$~���E�ue��a���e�i�'ƌ�G�1d�Ӧ�^�f��*%Llԕ�|�knlh)I����:�&��m�woy��k���<���Ak�W{,�iU��H�#�l���Ee�14V@t}�*���VVfDu�� ���3�̰�f�ʶV)'�G�^5�i��.A��l��3�!ky2��5T�+o��N-^g�~��~�|iW�𸐽�
-�a�jI�����$n}#�t�H�w��+���"=Qp43��oǚ�e��U�r�w�����ٺ��o3�l4��8�Y}/��=ٳn&�����=����;����{��dGB��
$�|Y�0���G��1�3N�3&9E⪢HrL����a����EWo���4���Nb�D�}W.�=�S!ɐ�_S�Z�s��ɍOyc��4�9�Bd��W�A)J�녇�ٹۍ`(T�=������$����`}4�(����+j,p�Y��:���8xtb]������r�Ul%����W�T�z�Ȉ����O�[[k~mƩ�e�WZG)�4��G�[H��i+�#�x�@�ψ,��3I>>�2�1�c$f�4|u0J�7����a�d�x ��E✗�x�DG$��$Eߟ�nx4�<鬭za��2%:!����B�U��'�1N\k�8N(�L�-��D�G��?CC�%:TK�[	80P��~EY58W�#4�;~��~n�<�>�֑�W�v)�����p���,,��"�x���M4�L0e,c�H�:h˺�r�I.!v/�Y��E�^�q�m��#��8ukb<,��F��R6�Xt�^�$;��f�ΚG�Z�oI��M?S�|�C�����)���L~;0��V�m�q{��]G�ۘ�Zi���ru��4�4N�)y�gu��l�3P���.4�0���8�<3@�H�:h��]��S"��Q{j&���Z��b���q�¨���1)\oK0�}��zgW��-a*m�!1��(P�-��8S�� ��s��\̈�+�
����9%+�
O{g/��2���{w���Ȃ�Ƈ{��F>"ݣ�|��c�N�|z=J&	<(S~\�M���yX�Ay�6���R�/��|H�ԓd��Uu��S+u���֚W�-O�&\v���N6Db���f��#�������^4��`���Y�t�p�Ѻ[�u�6��G4;��p^��Dᢦ�Äl��B�
!�i��E�3�M0��xf����tі..#<�Iq`����p�~����D�G�&��y#�D�Sk�-1�o�"0�֏�c�)��F*?l�v-�f-^j���Ekym���2��єo�u�柤	%���x�5��¡m0��짐�0D�هK����O��-�Z1YG?S嶌U���q	jR�<���Ζx�1�t�M0�K<3@�H�:h�<HY�~o�cڪ�(����Cg~�z|2�\��0\C��~Ąc$��kF�~����_k󯟢�������C�uÕ�ƿM�ã�Q����Fr�R��׫.a�FT򬭑j�S�����`�a�}!�")�7�{���O!�(������D���$|�i����d�Q��a���X<x��i�M4�,��#$����2]UX�����u:e��OE�H0�GD.oӲ�e��_�������^���CWT� $8'�u�>i��֎S��~D����?b=��:�}O�ʜ1>����$���g�&_ Q{��ߒ�D�?p�[go�/�m��ö���v��&i��&kG��o�>��F�$�>���+(e�f��`�I%�BC%�Z2��:iӮ���묺0��0f3����f���2�b���#$C�2FxfgI(d�0`�!���g�3��˭��:�uh�ӯ2e�FO<�<y�un��]u�����1���tg���0�F3M4�,����`�<3Y�Fa%��c,�Č�2G�(e��e1���ӳ~B�Ģϝ�˒-�י�x�	KB;��P/��oL�f2�H��C*ʪ�R��4/��N$6>��a�6�ۙq1�1>�r%ʲ��6��Sx��.����Y�Q�<M�����cƙ�ۘ��ȑ��j|Y_>]��k&��(D8Ikm�Wm�L0���5�-1
�d����ui��K.�U��Q�q֌���V8�,1;#�+-r�UuY+�"y�jjd!ܙQ�ВJ&���sWc�vo*p��>պ�N4�	▊��A9׺<��F�٥��K4ޓ������~�1
�i,mZ���;dL�WYR�k���5�]It�R�R�������v�v%,K���F�`}r,�İ{\h�1���nf��G*`��Gj�4h�])�cVf��M�}Z����r������Ȥ��;[^҄�cn�}�K��~��Y�ٽ�ǯ3/s37wvu��2�33wwg[o3/s37wvu��2�30�if�3��i�Y�22FI��|������*���٭ՙf��!h�s���`�iK�]^%�0�����9�\���ER�:�ٌf�B�;%��6�j�nԍ�Im��VkIn��Ua�֖����腊h����KK�\+]t���e,ȶ�c+q,�Ͳ�Ha��]l���	j� 7Zk�dz͍[t�ir�Q�%x�����m����ew@��`��@�c �n�d �eM{g1d$[��̛�ۼ��8�#��5��`��%��R��W�8�L�B��/�s�P`�����iD䥼0b��3���(�I�q3N%0���߽��ͳ_-�$6�.�������h����7=.�~�v�3WN�yh��s�j������Q�]��
)H)J'UDQ����V�4T���	�8l0�n%㤒x��L��M��3C�0�:���I$��մ�e�-d���s�����;�����&��:�x�Pn.�)w~��ɦ�a�xaM�)���:ɢti���N�a�rG�<i�y�5w�����,JvOn�~~a�Ҫ7IO��������6�*"[<�MWJ��ˬ�����O�4fX�0�	4f^�q
t���qv��T���&e>���q���4�Զ*.W����S�kZq��'��鳔��"$[��+��ܙ]D�v PE�)���/�@�7/��B6��ԟ�>�Z5K��|�z�ӷ�H�F�Nx�n�&�>�'	�3����k�d����
S�����i�:|i�0��`���I��Vr�&Aۈ^��I.!>{��)o�L��4�mĔ�2�7�er�D�N!fH�[g��V�aG�.��DҒD�Cq~�$ߠH��F)���U�%Zۧ�q�Q����imr�JWK��~)�l:�:O'�č�����(C��BGyT-��e�y�5V[�;_3�-����ZX�(,fx��Fa������Ux�^/kY��@�"c��5e�ǐw�OڠG�#�8�M�F6#�uEV�Z�(8R8��<��Л���H����nq�clm�SH�.J� 2�aj�1�� ���1-,n�&��U
Yej�J�HX	x5��tn��C盧�`��#t����w�5����$B��A">v��J�Y�I��	ܧS�M?�m�e��"7x�B]7�V������}��w�t��3���f$��ϊӢ,����	���[�e��R�E�31Q�A����F�uČ匢�2���4јic0c$�L:a�j�;Փi$����������m�#o�|��Y����LSXq���p�2I�����J�Y���=�-��1WN���M֘��V�S�z�iw�$�:Z�j�	b��� ��A"4�
��D�B����j�'B0��M4B�ԩ�=7�:��>$ь��Oh�4��1�a&x|xu�*�D���,�*����(�bj�Oբ?/WR-�D~w��܇e���l܋쿏��i쏑oQ����_�~
�ID�Q��ۖ�NN�������ñ��ߟK�:���Qm��0�F)u����U%��*p���}cQj��V(,E�R8$���U�6�B1X�����!�C�ch���sJ�B���ʄ��8%�V�qb҄#��^=�3�����)��Y$�7������Rz꒨*�A�K15,�0��A�jchM,�g>�T�ǁZ���&J�k�y�țZc)��5Q���VVTR�-'.�s�J�v���W�S�_k��B8���O��\ze>L�+�՘�`+���mu[IU���f{��XXʪ�U�vQ�K2Co�j4ŇOL��k�>b$�jE�|�{�8�Lj��hN)Y%�!��|݈Ɍ��9α�7 yc����v���ޖ1m��.�5��G�M`U�Qb�+T��y��w�xkLf?/R{[�YX�\�S0pK��{�����\3r�yZ[�G�V����3M�_7���0�����t���S�[O�6�θ�O<�<��u�q�q�8�%H��b�*B��Rz�d�H�$� Y���t��RF�H�Y@���E�J�m!���d�3�H)kFAI�Rc!Y`(dX(E��AVAH�I�ȫ&�犫:��]����v��S��O�s'���h�×csE�R�n�~����xh������e�j�֓㲌��)����D��]B��em�vu<����R��,������Z���F]~�N�M�a3^�:��Թo�W#:�)#��;i�<�Oh�4��1�a&0�ֽj/��F� ��/+R�uܓ�uz(]Q.����<ɢ���d�#*���FS��BP������p_UV"9�e-����^f[J��I���+x�H��Q�5��U�q>Q�&
:��K&�Dm9��h�.ܛNqp�;N��z|w���8S��]�0�~�DُC������}:2�h��raL5?C�9[H�#絺f��ۉS�b��ٕ'�����#]���0�)kbHħ��з��}����<-X�hcXIS_+�D|��0�������q�Ǎ4јic0c$�L:af�J2�+qUb'�Xzt``�4��L�ӳO��C�O�,F,�Da�!�������I&����QW�����=Ha��mU��a�}�Ӳ�[�����F���n��=0N	O߻-���C!�D�U���L�|R�����_CO��̓�4��8�2��G�N�պ��tf1�t����3a�0�Kǆ�:Ӭ8�F_0��ӧ[un�Β1��R� ftc0��3Yє2���Qђ2X�1����:2I0c�K�c,e@��:dc�Xye�ǞG�+�#�t��cC���1���3�2�2�i���M4f�XiE���xe����K��YG���tc<`ΖH��(��
J�EM�K@�He0ևX�� jCRx�z�v�x�pq����SXLa�d�*HVE`N5Ra�A@R)1�!Z��2L'��Hv��XI�"���j@���-�@άXfJq����1�b@P�(G).Z��ԕ'l1��MI�T:H)S�*H(y�A��\a%Hv��&���xGO��9s�){���D⿊�����7��{�������fe�d�����y��������m�f^�a�J4��4g�4јic0c$�L:af�̄�K�G���]6ˈ�%qΦ�u�Df���y�;;�{9""g޼ΔN�9�?�3	6ɤ-hCm|�_�ūx�ϗP������w�K�^m�G!hܥH,���'���[Eh�ӡ�;($E_}� ��J�|�"�D��.�G)o٩�*���q�~y��uƖ32L$æi|BI$$$��|�U���}cj~�b&�"ף�9�K��?��4O|������4��.4�;�t��/S�G�|���\]n���{״�����i�G���m�H�ڧԕ^i�ߵ�}*i��#��̲�-�iȓ�X?7�)m`����?2�|x�M��32L$æiz~}�����!D	�5f�fk�'n'L�`H��9�_����O�ETع�g��kGƋ6�*�ZQ��ãf��n��ze�y(��L�m�� Bb���ul����)i�+��A��y���o���"�������/S�>�)��"ts��O�i�C���"-��Yy�TۺZ>SئX�TL~�{���d����;4N��G!��'Ӹa���2�L4���=��P��놈������6�]�������XM�ڥ���:�>].�a"-�4�m��ϝy��y�X��0��Y�+�%$�����4�Mèp�>��5*���!���ͭ�a��G<�摭�ߴ�����dL"=�āX5�an:��e���H¡�5��טr���~*��v��Y�1���~�^�Ki.��t�U���$#�8²�-�;��%#��d��T��V[ɩ�(R7m��a[I�����3����|6/�Y�L�̾.�����֗(��i�>�i�0��X�I��t��+��&*�D�L���8u[}6�|_'�=�Jz{;�",�1�>�Z?~7wW��f�g/��Lw��1ÙmM��=N���?#>�z������'.r��瞧��W���*�~��x"?oŴ?v��v��?~n����SJM��2�8��#(�şi��3Fa������a�4�i.�����Sȿ%�L��V�z��ʫ�R�F�C�Sȣ�)�#,�֚"1�$s�ؗaJSiD�[V�C.�,�~���̢9\Z߶ղ��Z�0�b�ah�>�l��oԑ�N5]|���-�7K�]�0�|��|���S����KGy��8m�|�~��"Te�ki�"ΔagJ(e��҆h�4��1�2L:af�w�1��Rx�u=���R�99�T�$8�*�SV+��/��}{*,"�զ�鮹a�V���kڶ-�_}�x����|�60ڿ<���X��$o= VAfhD̵K���M�X��a3��m�O3�<pF<��;��ҩ(~UEթ���`�a�ågtpFt|`~?�w-��lm"5'��Tۈ��������~��|�%#KZ!�[f�Ͼ����Db���j�WH��9o�kS�Y�SUy���m�e��r���Q-S���L��/��]rS�6��4������3,e�d���_<!�Df��\B+�xE>g(����&�#g�wq�|�9[��rKm�~��Ɯ3g�m���<����'H,���Z>[�"�����l��F_�}}�ΰk�a[c���mk6�]6�m�\۸�۞ư�}'g��l�$��J ��Z)ᅈE�A�p��ӳuY�'pO��mo���9�8I�ϊ<Q�|P���2�2FI�L,�I$��3��=h��w����5�h�X]ar�W����u�R#�[5���j]#M�N2��7=���J���GL$��ۓ[�hp<;Tf�0N�{���)�ؔD���c��=�'���u�8�tĥ�ם��m���O�\�<�0���'���f���q���Q�3Fa������a�"�Gr�S>UX���Q��'��Cñ`�*��Q=���=��rF�u���22ƉR!8&�L�k���%d�x�ӂy?y��w���w=�F��=��Nd�H�֤��FkL9��M����Կ�L�6����k1�m�Q�jݬ��5����a�L-�����3��8y�el?0����n���:a�Zq�,��3`����<2� g�HΌGK:t�1�@��F1�&P�XtfgF3�0��3X�2�e���b(��c���	 d�0c�3���X�ac@�@!�Hy�Q<z�%y�yh��[��錱�c��1�2Ftc����3M4њaa�3a�2�u��,gK(e c�3�ጱ��YC#�&R�nH�O���#�,��mWbl�+	6DL�J�c3�,�Z5:�fXpv[KP|u�K�n�*s�C�y"��"}�����ke�zE��&�gC�ɼ��\���֪ӵ�V�X��Q��Zt�W��Xڥ�����a��<yv)�G��Z�Z��e�mx+;20m�yo+ rܲ7K;c۳��� �)Y��Z�Qlf6'Td&�!�ʤW�(���Y�oe�]����Y�s�/�x�fM�kt�:z��)q̘���c��m�e����AU��X�ڑ	����Һ����e�Yr�lK����LuX��ZBb�����5�7#�m�mm�:�h[6��2�
�t����ś\�r�v-Wuc7�}���kp��Z2�f(���ae�k��m�%I�z{�POWys���_�����ޛ�������n�www|������������m� ҍ<Y��҆h�4��1�2W��W��z;�j[�lI�7GAJ�rV�ԮԤW���P�)^e��i�}l�Gi�F��]6�B1us��¹�UiuWY��],	s�ͦ����Q�b�om���]����n�j�4*�u C6�MLr���Y���.��fؖXh�&o��"��̸e�5���JMu�5�Q;Fkqԭp[��R�����M�M-ԛKs�JD�]V��:X�:Ӗ�� 8!;�I��ɼ��y��V9��1�jR�Q�&Y�4�'�Eo3�)���ۖ�xe�r�7]FJ�Oa��0�L�~�Ȥ��#::?�I�DL����s����Da���Sgs��"��Te5M?}_��壏V)�8�g����	��O�`�;>Ta�D���,�x�1b2������-�Y��1�uţnT�Ǻ�mڳk(��||i�ь��X�H�0��ܽ�~UX��C������:�Ԕ(@$i��b�X�^���>��"^vүE�I�UO�S��L�����̜�}�xy'BR��(���0���eYK,iS8ݗ�Ǭ�r�2:���usP�#����JO.�{	>ea������#^���{
<}�|Qe�Yf�|P��,��2FI�L,�8�$��@@�G�|�?��/��m�d��1���s���ںr3�����{8`�����ڜ�[�ģD����WF�
E5�nÆO"y�#������SDN�{�V���(���7�?[s�
a��ӳ���yL5����:�5���UXi��i�_i�ь��,c$d�t�Ɍ�z�kX�<�Ng�*�D�㇧�BHtX��s|a"�0�L�˳����W۳F𰙀�3�eR@��:,G�+�,�����#�2w�����}ñ4��Q"��~��=�����{��w�.�S��N}=��Ȟ�,��l���e�	ܖ�ꨏSt�գv9	ѹ��۽ON������i��XZ�4}]e��R0�5&��|�O8��^mםu�X�H�0�ŝ~��S&uGb'&=�m�����Fz������Ah�|�1�����=3(�xvbς�kLd6�f���I���&Л��qX������ 8!m}>W�ǚ��[F��4�t��n�>U7nI1�E+��]�U[۪<�m�v�qmj,��+��I��k���N����moF���8d�0O<F'�Ku��*�V�a�y*�-��L�{0��>�)��9�}(��y�N,�*�/���^�c�G��k������,.e���[�׺�2�#�֕�m�nrM��M,���(f�f�ic#$�]@l^��k���> �=N�qEDJ~�L�I�H�L0�5�1L�L�϶�ב�<4�ó͋���W�DB.���-F�/��zPA�rD,�
uh`�N�{�p���-i�(rC1V�Q�)Zj/T��4�=Ka�1��x�-�W�Ȟ���3R��a�v�.I�2�Z8��0���(f�f�if���a�����U>UX��`�2\�����-6�EDq����5�isȯ3O��D_ݸ�y���-Id�r
���}ū�Qf�xp�X3Nu=S��S��Lө�iGÇr`�"��t,�q��ɶ��i���8�+7�b��p7�7g&&����V�FU�C�%33w�[(�{��W9%��%x��#yӥ�{�
1!, ���1t���ic>(f�f�if�����7D��U����r|p�N�вQ
va�y������G�m�Ά&��u�����}r�>�Ͻ.^^��%�Q����
�D%���@�!����R!$*-��a��Rߖ�`�n������S��s��9Q?E�k�L2��a��<��^mםu��,ђ2L0�eg�p�30�.g�=u�r�jlu�n6�13��k�g.U<Hвև������l�q2A����#��֚xǣY�|۽� 8!_kI���LM���H�(��f��ǉ��,�uf`�5�><���w02	;�x���&�"�ݪ $6�I�ϦB�Q�i�ώ	N�������GyЁ�H�K��BQ����X�&���i�,�PN�幗��B_�7K4i�'Ѿ�ɪג���̾�D�r���U(���~���E�q�8VƋlt�8zd<0��:~cz�Y%�3�,�K4҆h�if�h�&x�-,�IP�RI.!E���X4�a����,:�g,�Ӆ!�M4�
y"�w�)g�K;7����fC���h�" <G:��J!_}~��߽�(�M���qH�N�1>�Sl+��B��l����D�g�����-��`�1;=F��Ԍ#T������R�SU�\���v�8����8����i e1� g�`�����3`�adE3�$gFt�N�$Cb0d��F1�Cc0�I�����@��,e2�b��Q�xr��1�X�H� d�C�&@�3�0c,c,gD�Ӯ��":t�'�e�ǃCA�!@�bc�3`� ��1d���c(����xњi���4E3a�2�Yᅌ��G��1���xe�0��!���j�d��=GU{���������l���9h�mv�̋�E-S�7wwu������www[{�����wwu[�����ۻ���<A�Y��3J���Y�$d�aøTFw��O���a��7�w���>�;��̅F���4���ӡ)K<(Q7��S�0Si���nv�`%`�XN��}�E�Ku�Z%>�gR"�m��G�9ץ�4�7�/يb�8Q��������Jq���(�uڻr�m�q�.8û�/�i��J�<�3Si�I�T��0gO`�,�e�1�i�2N��8��$���=\���1��v?Od����yѣ�\��+Ԁ����s#V�P��^��˦f�ӬӐO��J0ﱙ>)�
p8%�NC$����TVi���z��ii�s|�r��=���{��O�F��xy0J(�"���M��V���-��O0˭:��h�4c,�J4d��<`�I����=(�X�;,nA�,N��Cި��`���)�˳8�v=�!?���l4��d�QT]�fX���P�C�$�U+���u���]���� �Bk�
"�H�CĠ.�.�&�30�/�lo[Ez�Bf ��s$|�6-ȡ�N�(a��n0,R�M�n����v����ts!�}:01���I换�1U�j��%I'Y0�0�fD�!���4�4���M4�]aW%z�6�i�G���H	�w<�2j�w顐Ғ��9|�f%q6�\���"3�z|먄"��0w���)�+y�<`�4e�1�i�2FI�0|��*�$gp���Q'q>�b&�F�'�?{2y>3C�imV�Ѧ.��;@���GS��J����8<��v��	>1~]�{#JX��dEb/�d����&2�����b,&V)��5��\��t���2�j�m��i$�����9s&"xQ:�&	B�|�%�n.7\ݫ�f�ɸSZ�X^�xi��R2���vuڧyœ�]��>8Q�p쓧�f���0���%;*j�0˯4�if��F2�4�FH�0��~UX&P�Þ�n��aO�b� "zt{�`l�y(�
��T)����ӭ/���D�8-�w�q�7[|;<�{4�C ��~ȥ��m��D�#�ι���>��mSN\��۩5_g�>m�"[�,��.�%eQ�^b�il6ۯ�4�FY�0�M(ђ2L0�J��_�E�	�0��^�����4�C�X0���S)��}u�3[��L/),���m�@}���y�6�ާ*�+.��F��M��r橺~�b��ղ�_�n�-�"*�3��Cɉ�-���o��OA=QDF�}����_'��K&��p�B�^D���|Di���v�`��~i���4��h�,�J4�FI�3�q(	Mg${-y�pe�~�6DJ,�+�Ƌ���]��$,Tq�0�s^Z4�dU
�)*5�@�h��tؤ�G�� B��A�t+�FZ�,���[W���!�a�n‷Ua�]���ʆ��F8����چ��]�9��3>��KG�p��#űXcˬF��f��a�FwN���]]8��EE�~<:g	�PB^�J�.|�dH��}'K̄��mD�*2'4���%��X�:�v9��}�_,�!pr����~� ���?|||`�4n>y��y�XqƜf���I!+nA:�4�G����S�8&�#2C�&��q��������d�P��L��J �,�#�K�E�,�
x��~�v�w0v���YZ�յ|:�X3�z���Oaɚ�`��8}���C�K>�CC���'m��&��|�8`�0��4f�2���i��a�q�rW�U]z�ɣU�+q�[�0�4����,ן����/��:�����xO�<7��֙�&��_6��C��kԤ��U|�z���z �L6%���i��e;:�U�z&w��K�	�.�z,�`rxd>2h�C�M�;�v|�a��QӚ@�,���0e�3�y��a�q��xJq�Z��6O�铴����~�z�#}�j,a��ƶg�B�XL�O��>9O�mV�N����e��j�g==N�a�`�~��*�����r~�xp?`i�u�0�a��<O~1̖��*�lX��0�)��������DQ"�ҬR*��{�<���tp_�B>�a��b�n�Mge1b��Va_@�i���{2f�$�Hxr�b�JB �B�	H"��rHD	HB�RP��!�P�BR� � ��" �A��b!�1A,eFD�D%B��BR)BR��D"���TB!(�BT"��"�Q	H!	P��A*B�P�%!�J�B JB ��R��	H"��%TA*	H"	P�B ��T"�B	H�J����b2 �ADF"D"#DA!"0DA ��`�#�(�R#D"0DB1F�A�"$H1"0D�2"��H"2"DdDH"D`��$��D��2"2"Dd"D`"D`��$"0D"0D��ȉD"0"0`��$��4D"*%"�QB)(���"Ȁ�
�QȃD`�$" �`�D�2 Ȍ��D`���D�"" ��2#Db �"AQ""0B""1� �""0H�""A�EH"�\DEBR��J�DH��"0FD��#b �����"1DD�#DdD� �A ��A"D`�$FDH�DB"�$"DD`�#H���H�DA"0FA$#DA"2"ȅI7	D��D� #" �" �`��F" �`�`��FDH�`� �D�$F� �FDH��$F�	D�$FDA�Ă�F�0D�`��D`� Ă�"0D�"A���A���C�""$DFDF"H� �F�������"0DA�`�D`�1F�""##Dd`��""A�F���D� $""#`�#"	�"2"#DdDFD*I`�#A"Ȃ$ ��D"2$#A#D`�"�H �������� �"0DDF���DH2""#DDb" ��DF"2"#� ����� ��"�H���Ab2"��A
$��0DD��ȉ�"A`����D�����D`�"#"$F""ȐDDD`�"�B0DFDb" ��DA���ȄDDDb0ADD#" �"0b$FD��H�H#" ��#DH���0D"0Cr�`"D`��#A	�F"0D��@H�aDdD�F�"A�" ����"DdH" �" �" ��H����" "F`�EBH��I˸w2RƫHs IA��B�	B�J��*�)e�Y�1HBud ���%!�������!)��"	X�`����"T��!JB�A�b�B�0AA0*Ib�"��JBBЫ�B�J�B���]B��!*��-����BRP��/.���*RBUB�HB�%T%B!)B�]U�P�P�D%T"��B*���B!*�A@��A)
���!
�%!%!�JB��EBRBR��J�B���D%T"	U��*!J�D%!�J�!*!��BH� �1����� �D"��D%!!Q	HB�B!)�BT*!��!J�B�B�D"	HJB��B�	���!)�J�!J�A	HBH"*���!(�B*�" Ȃ2 �D �!R�	HBP�P���"	HTT%B��D!	HD%!�n�J�Ud�"��"	P��R�D��T��"	P�HD��JA�T�D!	HD"�)$A��DA"D"�)�B �!*�!)�JB!P���B*��"��B�!*�	HB��"��TB!JA	HD"�da��2 �A""
�JAD%B�%T!
��!��!�B��!Q	HB�B!*�B�!�JB!��B!)
��BR�RP�����"	HB�D% D��P�� ��D"�B	U
��A)���JAh�Z�АB	HEB!*�*�J�B!B�!�D%A ��)
�B	HRB	HD!�B!*P�J� ��T	HB	P�D%!)
JB ��A*����!)!�
�J��B	P���!K�"��"@A1��E�B!*�B�	HD%!(�� ��TBUB*���BU!JB!R�EBUB!(�!!	P��J�!��!)BR ȄD"D���*��P�%!�%!��B�	HD ��bDD`�DD!*�����BJB��JB��!)�JB2FD ȃ" ȂD �"H�"	dA��2! ��0A�B1�A"A�D �2 �FB��BR��JB!R�J�T%AD%!���"�� �)�A	���HD��v2mr����@��~k���Q#QT$$EE$��(k�f�ҿ��{�3߯�����G���-`�r
:�?�Z�;������1�������h``�%8��ߛ(I@�W�w!�Y��ڍ�abI�m[ �б��C�b�!�/��l���)ws�����*(��G��v5�ӧ�G�������D���QG��B$B4/���ҾY��O���P��$3�F/|P���l�Av�;���?�@�/`nc� ��~"�09��~�?�bFr��h�e�ʐ9��gpnf!H������A���7�� Ji�۫<�n�N�9lJqRe���d1#�B0�u~z�ͧyD�e
@R�c�� R#�E�X)@D��DA�@EAE G�_0,I��x�X)�a�|G� k۪���Â�]PD� dSA B��
���PD B
�I*+P!PVY�z0�.pb�B��̹���PbG��7�� �6����b,
(�.b��	�����1�=�	Ehzƅ�6��W���������ǈL�۷�r�l�K���&�:��9���Л��$�A�{��~���_8p
އ�y�^S�3~��{�Ew��"��{���pl+����5utu_p@<�Di���" ��9>4E�:Gڃ:B�#�)��=M�5= Pn\ /��Q�!��z9�Pk�$dHI��$�w�]A�j EF� �l'�@p[ �vd�9����X���/@d d	tqC<�� �6��a~�1qK0Ɍ�����4��7�I;�UBr�W�E!oA����w��6�Np����O�n������<�j	���'&���ת�yE�1 �2Y!�P�/��+�nQ�QGqH@"0"���������(�/,ñ�s��~�\9��;����;A��zh�AiKN��`G���ӭq2r$!��0Y���=�j����/��X���|A���s�������Rff�(��N"�22�0���op��-�0���e���6�:�A�P$i�# qE�q�#��<�ʹxR���������n� �A�f����\D@�L��0��'�,�m#�t�w�a��򞴑��h(����7����ܑN$2Y�� 