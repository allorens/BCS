BZh91AY&SYM�=�ߔpy����߰����  `���   �� �  h� G��hU%���UTP�TE(�[`��Fڀd>��P� [�>>A$��UUQ@�}}�=5�n����w��7�ܽu�_{���s�k �-TU}V��p.��}�O���d�x��^��O"�wa ��bTx�٭����Vέ�����]��8��5� N���z=��\��m��R��J�d���/N�k���� }���.���j��n��'�޷;����\�\���u� �=ޚ�������w��:��i�Z�s�P }���`����>��˼q�����z��������;�������}}��y�׮�j���qݽ��EX�D|� y�j�v�������w�Z��K�{������w�s�͟m�雟��sݶ�w4p         )*���@iJ��cA�3P�	� C�&@�Б	R�a�	�`h4Jm���M        ���	U �`h00 # D�� �!��4d4�jzjz�FzM1@TI44�J��2z�6���M4`!��H~�Ȃ�$��$�H$��H6��KaI�KO�f�@$m#�l��B���"A#d���H�!����	�6��7�?ҕ��S����V��M�I$E�T�����c2ڸZ�t ��#�dO&��m����I$���������'��U�?��W㲿M�f`�#h�̺�Q6t#k˜(]^RYE��l���dD��Q�E/
c=M��ʱz��lPph:���ZL+(?�`2F�p&A�C$�-�P�B�OŌi,h�5�L�]��LE]x�kRi��"�"�"<� �H ��xX�ّ��� �4�h�$d�5�[$�xAxItl��aRZ\2��!���JB��P���(e�v�������&�G�U��$�xA�$șID��:��QQ!�$¢��~̃�'��,CiIDԲ��	���4�����m'Uz�K�ZM2�!�>f<�A2�Aه�1	�ҁ���i)l�$�d�42Xd�xA�	6ZN�-.^`7�ta ��	����b^%O
c�����J�E�v��d�����MX��*F�I��,ȑ$?3��K�&�t�;)���%�%N��yi[��[Ҙ���"�'i&*��&�E���9%2N�$,C4�	���'Bpt1��ePsi8��b����I�W�d���iyY �JabCfu��-�X1���e��p�~h�Aa`W �����6CC�%:�|�@T�RY;z�z�z:½0uac��f�L���/����J�c,N�t[k$�;��v��c\�bhk��U���m(<!������dְe��/A�f�b��M�!�֤�2��#C#=���*��"�f���8I�'b
c7��X���Ҙ���EPu):��e�8R���/��W�a'd�,CiT2��	�����\�!�a��A�$�A�%ό�&�^�Ϥ2#ɤ)�(xS�T5��,��N[�Ŀi�`�4Ha`W ����9%�C�!�Aׄ��e!�駫�������XpvY��`�^b��T�~�H�!��)��?`�`�hL"�p���2Id������,���M� ��V�#�Ċb�@"Y%���Ɩ
0 ?0��&����`�R E�Ė�r�ci��X�[���1�	��bE@b�Ʊؐ�?1l1��!��!���D1��=����ŵmN���X��7Bz���wl��Nh�d�-�8^�[�[+dֆ�#A�ZUI�5���.�LgMilִ�M�*�>�6�V�?T$�Ե�JN�F�e�# L�r��'1�9oA�.c�$�cr.(�9B郺��{,f�Ѻ�o|3��d��1VHB����q��K�`�	��d��E��
ak0�%�����6HvHbYhk�]XL�%�q���7b�$��a%�'jp�2ɺ�Me	L���M�y�tKwd�$Y2M�I�L��,�p�0�a�ᙌiZn�Q��Ji�V��Rg��/�I8�Đz	�����:ͳM�l�enV���H�f��v^ZN˹*�4Ҽ�]cJf�+��JJ�t	tZ��D��Ru����%�������.�xq�L��$�KFIt�z��]"�K�Pe�'D�E���A�$]F�20�I�I��zxm:q;ז��y��"�h���tj�D�d�IM%ueM�P���,�DY&KM�K"�i8�-��X�%d�"�,��4�Wd�V2�ٻ:�g^D�m�$R�
T]�G%�[)����"Z(�!��يe[5l��@�*�˲�xSd�⤖N�D�D�rn�9BJp�q�8���f��Meuך�ʛD�&Q6�v�x���X��;���vw1+x�=K^���-JWpN�Jbq,+F�!�C�	H�M�Z)�zLI-��yI6�֊h�Ej66���'ZI�I��h���'\�����ru�M�O �%�&��SRU��xCҵ�ܲq�E�8�)���#��2e[$絒�{�ʽ�}�@��A5�	V�ж��!�#XdF��A�3���0&�QN
tv�Y��&#�^$��M��ZsKf�H�ٶ��:�)ɔ�I&h�f�ͤ𼒩�Z��i9���J(���@�E�)ix�u��3H�w	d�
ZaaJ��o
rS'Y%���I=Eb.�S��+r��pIȬ*���]�e�M�DRӊ�RZ���e�!�!��SEB'QX�Z*і�x^d�$�&�Ji'VT�qe
,Q��M��f����\BW�S'%�	-���l��P%�C���j��YX���n���e;:�$��Ae-0��e�tsI-�$�R��d�"�,��Ɋe[7l��nʻ2짆��I�4�L��4]�c=�xSd�KRq�8ԜaKK�VD����X�F�	�FE�E|ɛ-zS�l��tc9���6��K��6uJZ"�ً3g�N�N�^�^�r�ji\��gv���٫/�KZKZ)���PY9H�e�ѡ��Xh����V��J�%��딛��RV�TfiS޻�v��!i�Q?���=�����h��)� � ��y�	�%(Ҹ��C ��Ѣ��kR
G����d��e�q��q/�:%�׳k������ڹ���ךS��1P����i�����fh^Mx{�����a�s�I�ó�i�d�����qU�������\��F��	��q8DДa$�$|w躤]}D|���	�`�n�M?�;���4i�/+:\I&�fYҍe&���t�gJ:�eU�7�����IUU����l�F�6x�I0A&Ll����I݌2j����dL�G�x�q�Ҹ�.K��.�Ӭ�r,��g0�%]��&����YV�KC�����zQW×�o�$S�Ny���n�>	���-�i��N�-�{d<x��I��[{��8����O�\3�=�����94U�F��n�M�؏G���р z�0�,�������#r�Y�N�Q�����M�{�_�T^Jw��А�O{�@�uyd͉�����~(y��;�;Nw�QK�|k��T�n���	D��6j͸ʃfϬ�&�����xY��<n�
뽉���9�i�[�Jӷ�/�o����N4Y�=_sy���lQ��:r����f��WQ&�`˝�f�Q�x�n'�*{�������hܔ�C3W�Y�7�f�.+f��(�7{bt�ѡ�=w�t��S���d�^�#b���.+9�UPY�m��G����y���5���zu_���o;�C{ P=:C����>[�Hx���
Q0b��"ٯ�(�wU�慐�pс�{n�5��{ޫ�rC�=i�3��8m���n��I'�rS�vcJ7{M��-7�1T���N�.�E<ܳ|�ʫ�$��c���Gg<�~9?N��g��&�$�M^�o_�/�I���Sύ�U�{��Itg�j�-��uFxxi�83���.��q����c>�7�q�{�^P��W�rn*� ��[�2���w�K���	�QSuK�b�_D��7�����,�]}.,�}u�$)�����1n��!M1������ˁ6H�(���7ye#�.�Ҧd��y.���&���f�X\h����Y/����'��|�e�����͓�p��E]�m^n@꞊�'��Q%h���B,���C�$�ԙ�*���6d�0��_}�c̰Ҹ8`��AD��0ea��Z�]up��QG�86�h�bb����n��U���O��e����^�����n��ٳ�eU���~({�ˣΨ�7y�I1��څ��x�%����o�����0�~ɿ.T�*��6I6� �L��1��i?Y�{:y�W�;�+�a�0�3��2�'bM�;��"ī��6L�,�vGu�\�~M�/;%w���
p�$�l�eA�e�0on$�TK�n������H�I'�d�P����g�-�g=�p��; @	�����l���o9�f���o��ZM/?Fh��ꋎ2h�erI�j�Ov��K�?}	�[�M�6���I�]g9�k6Hi��LP���9��'�����yM��y�l�9�7��5�G�
��N�C)��W��9�����B|xh�'^U��K�T�N��S$������z��j����fՒ�"wxсi���Qe�N�N�ۼ�f�:�'(ݳit�ˆ�J�(��|��*e��Nl�
����C>�]�:x禞��'G���;�5���)����7��!�2C�K���@׫� �ц�y�4MD�O����L���5F�,����>�{ z3���a�	���Hd�H(J\��<t骘��h�[I�ՕFMGvQ5�PA����9:�:�G��4QfՕQ&6�8��G
,vM=4���6����r��	���|�s2@p��N���?>����y$1��@ �x[�Ҝ{��Fͣv:���Y�ŒIq�R�fI����=<rzw˦CN �87��  �3�M�^���6e)HY�����',ɲ�`�/�I�*N���𧧁�D
9�l:0�M�oy��Ç �=��zEӲ��:3F���'t�:1}�-�z�)�ۼri����;���M��Ēʚ��q�<}N;��P��f�ge�j��Fp�<����O 
���G�8����4�ӡur��5z�|���W�9����OO^�,��
]8�3��~�<��I$���c!��y5u�lvj릟���O�"��d?k�O���O`ɇ��O+�8�̢�2�P�'�Bۧ�����m�y�K֙jս�n�J(�z3��gI(�%�#N�<N
"˜�">BvN�gN���'�H�D�Ի��Rz1��xQ����PjOXZE,����[�!<�c(a�sW4ސ�@K0�:�(\$A6WT��X��u�5f�W�1xhdS�SS���EZ#�O8SQi"c "U#��協��&���MTFF,�|h�������@���m���_?A"-Y�M�l ,�<Lؤ �������~�Ѭ�]ݚ��K���P�F��I�>�u�~:lH~�)�hO��r~��~D���C�w��O�'�o��7�?��jh���H	���N��T��Z,�S;n*Q�'��6���L��,�C�c5��qG�,¹G�k�"���SP	i��u�CYm�B���P���Y}�;}.^�*� ���V�Di�ʳ���-8Â���y��_w�7Ü���96h�HGL�#-�*��D�.Fr�8�Uhs�y�ɘKoEĆ/�Zvb���M�i�
��f$�����Ǎ�a&w�^���K��Ӣ��u�Ӊ��� ��m���@�/�$�Y�uEM��w���ۺ<����s�١��[;v�'�R�����w#bQV� TG5�:v�VV&�3r�ǩ��a퓩��o��cnYי�����hi�'9RŽj�'��[\/�=�1f��v3��rd����H����\�(�:�}�)��S��6�Q�Uih�^���N�kD�i�qn��)l�ID(��r����Ey�N�&���n���*_^x4un�+K�q�13Õ��뙫o )R�u��>��
��4.$�'7OA�SkF��He�m�����Z\2Y%x	H�z=g�)vgb���&\��Z����l�h�=V�Pj<K�FL�^���,k�(��T�b5���\z��%�)1���-�ΰe�f��xw:�;w3���e�%oz�̈�:u�Z�li�&�u=!XD�q(�;ihi��cU@j��q����3V؁ �5�a�:���Y��1�� ~���*�Q�dT�q��!��j���h8C��~2����?������~�}?2@?��u�ۭ���tۀ�M���m�m�m�/wen�Ʒ��m6�m�UT�e��oXm��z�m����6ܶ�t�r�p�m�p�m�a��m�m�޲�m�m��{��XA�A	I}��l�6�m��n[m���x�m��wcww]6ܶ�rۧUUT�p�m�e��oXm��z�m��6�m�m�m��嶔�m�l��m���m��m����mǽ�<x ���������v�[m��m�M�-��m�a����[�����m�M�2ꪦ�ne��6�6�v�m��l6�m�e��oM�۶�6�R�n�i��x�m����m�ް�m� (�7� O�=��{�����v��m�m�m6�om��sN���a��vۉ�uI��vۆ�[m�m6�om��m��m��m����d�M�-���6�6�v�M�����{�ڢ\IK�{�t�w���]?6ۖ�6�m�m�l�������m��m�n��]��m�m6�t�r�p�m�4�m���m��6�m��d����6ܶۖ�t�p�m�m6�����������n�nXe��m��m�z̶�6�kt��޶[m�۪��a��m�-��x�m����۶ۆ�6ᶛm��6Km�e��oM�۶�6�t�r�n[��|�@rDJ����1THUTZ����_����~��W��G�!�O�~C'�?!�+�o^8���n�q�;x�\z��n=q���q��i�+�N8q]�i��xۍ��N1\8p���q�q�����Ҟ������ÇW��t㎛qƜq��n4�4�Î+�����۵q�8�nx�=q�W8�|������Vǝ��%�&�Ť>�C�U�)�Ae�u�1�b]q�5d��:�b�*"��aY�텋�XԚ5)B�]� &4��wvȿ
F��$8-֩���D�nY�$��J蕉>v1�UKrY�Q�ee��k ���yc6��m���JR���\0���,HR�Bū���!h��FIK�h�b��F���J]I��e�*�5��5�!}v���U��hB������D�%!���.q/��	����u�$�vEףkt��-r�ſ���5T�e��Ճ �ڠ�MT;S�
���8@��6�L�k��s�Q<����� �CV��R�'M�-6
�QH��ϭZ��gh�V���VTL\�u�Ff��Q��s4�4.��nj�*�7�R6�nK��5ls���a��5�b�I+9n�7QF�y�n6��1cR�Xl�5��s�-�o;Ѵm�eQ}Z�f�WO�\0�aE_bcR��\��]�K3)-%�Ɲ�l�Q���4ҷ�hCOok�O%��(ʪi���"dTj���b�[��݉mt���]s�ؚ�f��5��)��b�]K���`��i���l�&�aB1F�m��ΐ��b8]I1,LjU�K�Qn��$�XnE*��]G5-��fJR+�f��4�u���,\��R��t�~T�ֱ����!Paj��Ai�0��`崥r�KD$��\��Bϫ�ojf�[`��![�b=��&�j�إ�i�x�E.-��9d�Nm�;$F5��$D`L�ͬ��جL���Be�Ō����Lg��`dB�l�SQ�-�J�h�&.�Mma��%$�[u�̊,�6�63�����M�VB�kqt�eLh�l#2B�@�
L��7.��(JQ�蝴`��[e���`��FjU[r]%]�#�IW�H[(�,��5�ñ�N�Me��	�G:ކ��n����k
c5�f2�we���'Dm�m��vмĘ�	50���$��H/�}�M��D��TEq�C�� �V�������p ������Ī��<��2Q�N{��1�yEG�=�(����g�<�*��%�����ǑA��Jܻ��f{�����q*w.��ؠ���.������ؠ�&�MK	���?g�jR��ų-�,�d�q�Lm��Wm>��m,v3]Xm	�qaI�m�l��c3�.��:\JjK�Y-��J�]1�At|�JE}�٥�IH�IMt�\R���Q�d�\� �۬���ƚκb5��72]b8�W��͖�Xd��r�1�L���(���\��["Ȧ���5�̕��(YiYD�,&��v�L�������,�me�V	$���"6'F�Z[R�+`������[i�����'ᤴ�֪I�:�pfvJ�!UO����Ӡ��#��u3��W���8�(�Om��#�7 �j\YěM\�,pém���,��d!��x� C=��kˌa>�c��ǵ=m�Xͭ������UU�c��]v�0�)˔�k�B�X�b�[����l�w/�&-^,W���+���jwmn-��V�4�1�f�`׾�>Y!F��c��qs-�4�H�MQ�˪������)i}I��S8�f�>|;��Y�����T�ԑ�D�`ؠ�����Y�ઘ�<���$�D-qVj�o��;:&wS�*W��1�W�4�1ٳl0��u��S�<�O���qq<U~G�I5VRѝ)Ѕ�gH�n�n��o����7�ZiZ��VE��Vb��!!UHM�MU&m�MrI3���O��'k����*�q��m-7N���P��� ���n��H]l��9�&�4���.s]P6�k�啶�9v�Hk�!��^�����r��U�2ѩQ�h^��ι�����a-��&�����j)h�I&�3fY;�ք�S���צS&da���y�He�L�Lwra�ra�WwÏ��;BI�(ҹ��/{�E�*�Oc�ٶc��j�X.Kl�
�]�XҨ��DDjm8;��]0��� ����[i��Y��-�v�U�u��r���q���.�����m%W3R��̙O&^<r��^!,��8 �L�:tu���zqÄ�dks� I!$�i����'���pDG�s��"-)	
x�lz��U!Φ���d��vfl�Ti��<bc�x���}ڔYuS�e�����أ��}>༮nT04P W7:b�J/Qi��lٶcQ�h�m�w:���=�8>1�.sX1�� ��F"�Hi6K�䫎��LZL6�i({D�L�[�)����:H]]$z�xi<��Hki�0h��,���i<`Eמ�x���t�jt�	��;F�r&���V�o�۫FSNr�ʉX�x�\ٮ06�-���)a��j�$U��,
ШBEY��4k!kՆ6.��ylauMm� ��ZknlA��F���2�������ӧF��s�PJ�&�&����̒HJ2�:�C�ˁ�#<u��=<fN{
�g�FLb��L�Ū/���t�X�44]@M�,��,�f��%E<���0�
�@=F+4w��{$%J0�d�n�"i��5���ZrTɅn{�������|9$�"q2*�H�C�):h� �{tbod�6b�w.J3��&�j����BY�uxME��<:�gMǤ9����M�&���,����=>'���O|����x�|N�if˂,�|�	�G�6�c�d=�$��h}��G<Y �
>���~OÐ��*��NE<(���#��c�C�G�#�g��|>ta���O	�d�>	�<�l~2B�����|$�5�G�4��M�GC�'�+����O'�O��<'Gã�6>2J��G��|(��Ezsu�#�c1f#,11fĩ$�o)�H�O�8sw���C뉈��I!����fB+n�R��G%y�Fa���^+���E����-&z�)����،c����w3*���}U39�p����˻��g=ß"��]�U388s�T�]�=�U3c�>EI���9�*OwtWu��פ
(@��,�l7ZXX�ag�x��QE$$D��ll$���f|Z�P�i��.����I�!]T�'S���I��^=3d��۫�H�S}"�SLQ�W�ݚKAᆟ	#��) �2��۞���䧉7�&]��e)5�BJ�8m1/	a��,��2V��"Y��ՙ�(��*�;),�!%��/�%�J�>�%��	h�)��AYaıd'���'8P��Q���	�9��}F���~��m�~�U��"]��D�4e�h�x�UwfSO���z��'�#ȱ�~�BHR�3�������)A�㥖Ye��U��e�����G�������s������*��nd@5�E��[Z�eu��Uk2�8��@��u��*F�:k�T���{\1�K�4�n�m�MVnͲ��`J6�$iŴ(N�nc[mU����돞�����'��Ԅ����Z?���ç��U	
�P�]we�dNĲ�)��1)���Ə�$�G t�R�֗,:��M�S��0i����:�(J���U�S/��������-"p��atgM�L�2�M�/A�p���_[�V���FIV6�����W)�0@�b�&>���J>��z��M4�N���1U�=>������]EQE��բӮ��$~JV���KXL�(z�q"p�%�rJJ�ZC,L<:��&ǳ�*��_����Fq�U��j�i���Q3:Q#��dR�'}�b
#�$���ĕTJ�>2���K��5�iP��	bt�J��>���7;b����%�������|��cBy"<���q6JHa"h��ҌC���&H���Q�Nf�*1g��z�M4ӣgnԁd�}��WHբ�(��q6Ӯ%-p>7	6p�&R���b9�RS	�	Iƚ�I�$"��h�J�h��J��R��Ex��چ9f.VX8eʊ��#$���*UU�6�Ì0��'ZW4�͑):��1}�(�͗L���3H��0�d�'�CN%]�6Zh�.��RZ������w���:x��M4�g��Ն�%������,/B8EZ+�ѿ���m��Ar��-�&�n+��UwS�2*�#�s\,�hh�4�_6��r&�2L�{�If~)�y��;,t�d�K�r�n��1��"�WFL�����j����FȚ �`��&�l���M��D��p�$<īm��i�͞;VcLb��sκ�}�����V����)NG{�jݭH2�d����V��H�;ͅ$}!d'}5zC
E�*��6���Ӥ�En6��Y�1�K��6.m�uY^�h:�)e��ʢ]J�SX"RE�ѠK�y��$|�JL<�h�R�6��#�&0:�JSl��Za�N��q!%��%o'̓����c�������6H���Q�S+�A@c���p��Y0agF�_7�KX�h�j�l�cm�F�qdL�`�^�,N���R�O�'��&����x��M4�N���VQd(������c�c6]�]�뤤���ilG��o2�n̖�`��=�H��É�Sq[ђ�ap�)>b3�i����F�[`��"2���"�&�3�3��M'R�F��0m���N��R��	䆎�`�#��:�����(D���>!
Q��I2�Յ�B��L��|ӄz��L(Pލ&�Ț�m(��iJb��.�l�cTYtVC��;dGG��!�]�º���ب�:b�4n��)4�/R���Ha��`:��) �9%�|zHlܒL�Xh&��cD�D��i��=##Fb��*�];Fh��giyg���ctxqڰ�4����K�uu����vRd�ʤn8�^D�4�_�&L�T�V.���b��}��I"'^�'�}u�(�d�QzU��(�	Dh��I!�l�e�$ã
�2k�'�eD���$(!I�'�i�{�6��a(���� ������H�YV�]��t�8��%%N5]��'����d��xw���I��<=&Eْhtx�O������|=<C���#&�Cdn����Œ��(�����&M��FM�&���<YH>��'�������2>�����MŤ|"&����x� ��G�'���O	�2>����|&��d�	��d �Q�5�Gâ�^��:(�Dz1Xp���|`��|9��xO	����G��4<<d�	�G��|(�S�r~���WtG��I��4^=8,L���D�'+:�D*�����O�$��.�ݽ4܍x�9GiD-1��D$�JfQ� �!T������6�e-��"Qt,�+&x�R��'(Z���¥D/f'�.�g�t��޽/�z&��7��6oe�\��m�z�d�e�|)��_ �O[\3f�*���&��Q�n�v�:j<�M�|�k��#��W�E���r�;7��]����Fw*��;Nŵߢ��/bu�LQ�*�;t��
^ˬf��d.F�d��EP�cn�BI��aTV��q�3�a[�����O���Lq������s�S=��ݗwUC�>EI��컺��w$��wGv]�Up�䔞��˻����&{��{.�ꀐ(P���>C�� �)D~�}}�3gZ�.D��J������ܹomn�5֥���jj2l��ҥ��e5\�s�L�F5.�����!�L��6�4�a���m���ik#	�#"Խ#^$ΒSSM��i�n�m[*󌱐M�2�1"�j)*l @NBֳ�t��J�j7RLD�z�Sw���n�B�%��^�I6ʸ�zl�bRf˴�ZU�h�۶�.��7�,���<ip�e�r1V]i&$�w��|��O��H%�O�1?	Ɇ��N�#�<�M��bj=�	Mr���HT���;@��ɇ	��'�;�#~�bM�KF�QI�e��%/R,�U���|L�T���߭�WlGTYi}��L���R�k�Y}ۛ��&�)$�RL��wl�V
)8�a�	�%�����57��e�Gq��C�M�cӣ�ѡ %�C�s؍�9J1��qG|���^�>K[H��@2c鄴���+��)8VXB:H}�H��C�v����R�*�_i���M`5B�Hy(�h�ܐ�:�IQ*�^�T��m��8��pخ�nkG����am�IjI$��j�m! ��$HCES�!&���Ի(�8���6���^&>�%/��b�0�I��Y�d�1�:=;v�+M1�ʶU^��8��DgZM]�w$f1Lh��H�SE��RQӉV��P��	o��Rמ)�]@j��T�0@��o��d�Z�GV|��/+M�i�$���K�1���Vq)��k7X����y/6�Q`F�]]]&�D1�*�d	|kܕf]|�Jva�fϊ(���ƈ@K,��S��-��F�F�x��{.x24@2�Jl��*�ƺ��9�%����#�o�CX��1��T�����<zf��H^	��O����E+P6Ze�"Fm�� �R�4E+�NN4�s��5$���l�e�*e��q�I�@50��0jM-�'�c�f��X����1�:6x�X
(�������t^�?�{��Vݨ���*��Q��ҝ�@W,�$R�޺�9��r��]z�9�\��S�U��Kk��}�O��E��T���cn<���Ypq<,S��ߙX�;J&#�J�,�oJ�
�S��(��p��1*m�JN�࣬�cFn/{� S%�_y��r����L`=ӼNy'�UHu�3����F��V2G��l7�!)B�M]X�2J2�x�*`R�3)I�E)��˘{	HCf e90�u6�=ڑ$�0�F0�zC�DǍ� Dg�Иyd��� �%5�I���ݽ�<:qU��G��Յi�;�7նDy�\�)�>�k�Qy�U��#�`����a0�{آBoZ��U�����)���6������ZUda��<�~t�|�-7JH��\:J�$~����2ꬩ$�SI���ɸ�Ii�%?$F�쯒ZM4��|�}զS�v�0�Ki��� �#��������۵aX�6��O����=�D$�B��K�2��28!-������%5�%�y����v�l�4����6������w��7��1����6�J�@,J�������'x`m��'R��l��8L7ײ6��+0���E ���>���W�$67݋{���E�s�������ު��&�����&L2Ѻ��<�e���L#�ϓ��k�էʮ�txx�XV+O�?d�TT�O�ou|*�����u�^܅�5ש���}H��FB@ۄ�¶��@�m��-:�ĒB���a�i�KE���|p��I ǸMK�M����#�HF�Fb�K(��lG1�E/-)�	I��,o�p~Ux����V�}��_�o�i����U|[b�c۶l���ط���9�GƵF�5ܞ%���54�)�I
FN�K�������%!�7�1�F{��
�i#��XT���4�R n8�)(�+o�H�7F�>h˲>cpG��aM萘A<JM����x�� ��{����K	up��Huƞ���& ���'N/q��*A�H~?��c��:�ٺ{t�l���7���CτN�`84$�g�,\{	%�W�7�i9�J�Jz@���QѪN���`;I&df"D�JX��o1 ����mD���&?18G�^(�͒��~�%����֓&t��|��G��� �D�UGp��2�H�jJ�K#k3ն���?,n6�P��N����|��Η��t�;�I�:>:N���h|l�8C��/�����:>8Cgc���&�%��,����<��,�'ǎa�pM����l~������$<C����O>/�A�A��9�"dQ�%#�D�`��� ��O�������r>��xO�'���x5���T|(��#�G�l|5�D�z*�=�c���>���O��tO	���G���48=��`�|(�q����8+�zy9�v�jm11/��
l�fV��*U)�5�<J��)�m�R�Zr��G36�it�J��G$��W`� ff�)��q�����-3�vȱ�lPX��- ���%ݻ���{�%۾t��K!��?C���~�~˻����&{��z���w$��wt�e�����-=��=Ywuø�:{��z���q�t�wwUe���A�U�N�ݫ
�y����=��u �İ6@.'4�E1RI@w��.R���=�R��*�&�A��̸���AF�!�������ڻ�&��ɺm"E* ||����t�Za#ö��Pĩc��Rm2��#ն��K��1jy<�n*��;r��0lD�f��B!�ǿ>�&~�3����=|��wI���UUV��ZG�/)<D.�=���]�w.��dHKSTmHļ8�I�i�H:2�|Ԓ�����m%�r���ƒњi1��H�H<`�JLM$o�$�L>� ��|��ZP�'�I�n���J�X�|B8B,�l6hH	�?C����K˘�,i�o-\{}{�a4�����Q���;�C��Lٴ %Eڕ�0_3�/�a�!aY����X�F���M.��f����q�6�P��fܙh��6��N?H���)��l���q�h�_i��,�p�@i"h�B��@�GPud��솸I!�����zXѧ��7ާ�$L��hi%'�L�=iIď�&S�[N$n��(�
�Z���VJ.�G�b�Y5����Z��� ��Ǌ�Ν;V��#�j$�ɖC�P����&���O$�2�Jdv�P��d$!n� VH�T�H�ъ��袀@߾���r�zb�G���2ZQ�����Wz���Q�KbB�$�VT��i	��L�������R��66�HX/0�5�4�d*Z[жAp"�d��L��$ O�z�`��.�LB���P��%�d�����������&�v�6�TbDT���7�j&�c2e�EfND��(�.����2�}x4��܋��G�/zp�Ӿ=�����X���O�K�Lܤ�~W��vlYǏ?F���Y��œV(Z4��V|���Ӱ(.�i���C�Q(��' ���r�d�=$Y>��-j��x�DM�A>vr�i�sw��ɡ�}	$v��Mt�x)2���t}�;F=G2(���{r�08p�ԸJ*HF�� RY�&�H4�2�I�<�-2�ywH��*��NL�]�x�~=[��:Uq�U����V��j���=���c�Ӊ�q��8�f�`}T�.��LbY!/K�%�cf����Z�5�hEǶ""Vkev����T�He2��(o��R��X���Ha�4e����ө�&HCf�OA;/W�e����ssH'�ij'j�f�5C�oD��o�
�ꌲ���uI���UA�}��K�+.�r&0����Q�k��Yea��g�)�AF���W+©� dJL����IN���$0aa�ϝ&F[�Sj�pw2�I��OpTL�"�ױ���|�V(�^;G��%x5�]�ˡ����FH� Zt뷯GI��<�xh�>8B,xvڰ�sϺ���K=���6����)8�7��� κ�ϒ6�ɏI8�:;t���5ڔa�:(}��������`QE��>~�O'1�Zdm�����\4.��g͸�^1����ӶՅb�����xW���Q�=D�������q54B0���'G�h�K%�,Z�1��$`��7?I,R�%!�;�y��/]�Z���q����M�Y��ڏh�v^��i��W���-Jϡ$�'1�#O�M;=�c��ӶՅc�~�Ӳ<q��:�J��5������If���<<W�f�~�*����Q*�ܒ�&ObB	��--6�y=���Ē|Β���o�{�7z�O��̵[Fp~a�V�0�����5�@H��*f�^��p||M��#��N�Gm�x�<�W�قe|M���	�<t�^�'���t|t�.��hpx���a���|	�|�flrl�=G�48<L��Œ�x	>>$>'�|?�tr0N��< �DD舙z"t�!���|*�.��OE<Bt�+c���r�!�q�+�x�k�:&�EȐ�T|Y �����׍��\>$^�G�'b�HN�G���?��W�Ǆ<'���:5��rp�z*=<DsJ�(�Q���L�����ޖ�K�j~G-~P�L/��9�6����A�D�j#x(JȽV�0�1�N�rri�A�֯v �ȸ�'��5��P�R��֊���gW1�u���k'5��{�ܹ�.��$�Єz�~�q�W:�ǧy���$�훺pm����5�o���;�u�v%�"ּ�yCZ�xI��ʊ��E��R*0��`��A���S��ơ��ӯ(��'0�)�ش޻]%�[�u葛��'�v'�G:W���s!5����߱ũ�Mu�P@���ws�h���@uC?
�S��8N'+�zseJ�K��\H�B�ւ.�o9������8��.��]�(����.��wGOwwuUe���<����˻��y=���U�wø�{����.�q<0�wwUV]А$P���C�>B	�o�>/�.2��]wI�!,�(�E��s��c�V:ke�K4��ʷ2D���e|ݶp����!º�o%�˥"z	��OG�m��F�kksjF�1���2łk&�u�.4��].	rH��i�.Mz�+e����M�˱lB��$��t�bƽv��q$2�ƺ�6Hy�1=%4�
3F6��Z
���V
n�����I-*��l�R�����X�+��Ǳ8�L,x"��&��MuG$D�ִ¢ķe=�\a�+؅*�,��!��(�h�qGƱY��{Q�wT@>�Ǹ�t�q�*�r9M�:��w+ys�}�dMy�gm7 ah��ꌛ�{l��!�>c��X�r؃��R��ڦ}�W�"p\0ۇ|��I��FQFK��V��e��FO7?����YJHL4m��@�+~��D1�6�#Á�*e>mѣ y7�|��r΢���Ke�$$YۺIe�u��M��+�$�dt�[X8L�O�Z�WsG�:V1��ö�c�}��T
��-4��13��&L'(�ոl������V�~[�e���v�h�ꘒ�]��i	��
[�0���L�/� g�~KK�hfyi��Q$��O�C�f���p�v�--�]�X�_d��j��!��at���l1�N��y�UW������;.�f�h�����]���+$��*��[h�y�T�1j��rDJ��}WF~��*$����}�v��QfJ�n�d�r�BI%�J�*1�OQ��ҹΕa�+T�!g2����n~{,���ڞ�tc�x�?Ѿ~�$|�Mg��s�F�F|���6�� H�q�-��u�bh������p��5�0�&���WY��Fv�r�^H/LSE����md�Ѝ�"�w���L&[��ޒ��Y"51�ی:��6՟�?N�Yw�ϔ��Y+���;�yV�����±�v�n����&�[,�;B9 �_fj�r�Hb��C�**�ĒHp��>UcoX�=SӶ�c�_�a�&%�f�޼O�&Cf��t�N����	a��O����_h�7�����i�i��/��]��x����{��}ƍ����$4&Bf]G=��5�*�۶1�)��$nd��f��0��7[�|���B��锾S��!䉸���TK�Q�ރ��U��S��Č%L�X��O���d#����U�}�� nz�CX�A�qx�h�$r�P�
�ǸsWUR��JUC��#<R|4CO�Kx��w�:z�g>��g95yWN�X��Ǫ82@���ր;\<������Nǻ�_τ����z��_�$�CY�ku�Rx4�DW�+�##��k����a	��h��C+>L������L�u�$��ç{�:�����6�j�v�c�;;m�Nx�?[���𕼉hkL�:��QF�&���LAgb+'$m��@STP�$�-�Cii֜��Z:�YL�Y�	$���͛U ��Dx��ؿ\[�#�cᣡ�nj֍k���P�F��Mm�a���Md�L���-���DǞ�h�bQu��-u����uْmpuܔ�R���3�dK����l���=�mҫW�W�xX��B��;����11U W�|�����A�iI�rHH�nL�0d6r}�ܺH>8���������HE-a�bbb?/�s�/[�8<�!!�ؐ3���a��1�p���5Pk�f��1�4z=�ӄ����!��=\�,ْh|n/������:C����x�'�D<j.�����#�tx����&��l�tN������l|Y!�d���G��xa�x|'��|"d�N�DD�Xz"t�p�t�'��"?��|0~�Bdl|&O���xzx�D�d����D|(�S��D��آlE~'����O�FI��&��|'��!�6'�#EG")���B���b/r-�Aw=$�<�Mwe�gY}+(�B
�L�=#��Ӑ����6�TQ2��3���N�:A�;)%`�n���6��P�I�5<I1�1��
��.����}�U�wø�{����.�q<0�wwUUe��xY��˾�����ꪬ���OY��ˑB�!@��Ǉm������\ǁɎ�͏�=���:N'���I��	$w�מ�\^����bਜ��t�2*��e]��	��'ɣI<�ޙ��&A���|A��&S�Ci��b��6���]�����`�Rd;$-,<�0h�M:	���h�"��0@�Ѓi�cx�kN���0���-˪9�A�[�ǸM'�h-��%�{�񗩵��M:L��K�JL���GM�!�� �h�W�>I�m��ZۡlL�r�]ݷF�Fͣd�Ǽ�J�u�Z%\�#*�i���[K��IZ����1sl3���L8n��[^ŷ	[�ҷ�-.�V#�$�<~��W7�TN��7�M(�tn�!
NXr�B�r�$8�,���M�'q�U���X�L�:��h��O-�S���n��<,�v�N�*��W����a��v���G��ts�}+g��B0�%'B�q�]a<���W�S�}d�L��c��qO��"����W��RV^ʬ�Ϡ>�,�Ϗ�,�>�TW�wIO����q'�.�-�"�'�J=��ꓵ��Xm�e7F���T�M�Ò�*�ګ�Ӷ�c�׬��l�`h�i�a�̆�o�/�ƨ��ЩUE��Q��i>6��y4�����������M�Ijƴ�;�>v��gFP�N���x�6����Zd�o���½��9���a�ʬiU�ӵ+o6�Lˋ������}G�o&���9���+$gUF�j&�ь�)�6�����y�7���8���4�6��q�iJ/��5$$6ZG	���~JO�#㧈B�!�A���>_A�{���a,������zҳ�����Ż{2��L:�R�F} W�=I. � ��n�6v5�*�s%Mv#ue�,�F�����3ąĒBI2��j���}Y��"#�a�F�B�7CF^����h���R?k��c��$�#8d�0ϥ����B$�J�t�j��b�2h�gp�e��r�w%3'�Cç�ɓm;Uc�������(� s���t��4`�U��I	'�t��6xӓ���.��m�L-�Mi�w]�֯����.ɺoi�<�I!��`ZSaQ�e�ܶnwiMwW�&:mU�ʯ�G������ɝC&�.�J3Y�֔�`�,k�W�p���uM�Ƌ�c�1/'�1
E���MܱQ�*�C�j�ΕЕS
�_4�\�
&�=$*�1� ۠����㥆�ܞ	�ï6]��oXҫ���ڕ�Ӡ��7�i#I��a�������H�e8�0�ݜl6��a�H�i�r�{�&_;�I���N$He�:a8vI'G�򪉿V�A�
"nV��p���9������-�?I�V�0�	bY�t�~&�E鳶���O'�c����]����x�<>:O	��:x�}'�C�QL&����'���<(���c�ɱ��p�tC����0>Hx��Г�#��<3C<>�>z"n.�F�	�D,��E�5c�'«�WĤ|'��o�X�|(�L�!����t����r|H0�*'O����&�Tثㅈ�N?��	�>!���+�xzx�D��r$<A
>
*���e�.W���͛�I'v�ق�U]�m@La���2B�ٞ;��zyԟ���]��_6x�8jl����e�׺�s�����	�9�溶^�|�pp>��5��9W���O�ث1���L9�El�Ŋ�%�Tv�~�ԃP�ٔνZ�bSÕ�4����D���D	�Ȼ$��WcJ�F����W�$̑�F���!E��'^y�syy#��tqq�]�������<�X$-�i�+W��[A�G.��5�Z�Si"�[J�W*	��ͽ�j֤�P�Y6��f݊�d�W�JC޵��]�E���05�Q7b���=��Ƿ�uUV]��'��wwUUe��z�wwuUV]��'��wt�������������B�!@�(P�� B����F�����6����]�=�1�Im���:]GmI���'lI3^c�2��Y���u��ʛ�L�����IKI�t�8Ʒm�b�Yp�6lqzGXMq��&Ó)�L�4]Q+�+f$�4-$Ik&�[#J[k��#.�uŘnd�m�ǜjK'�^M��H٦-+gXi:R�R۲h���GW���5n*L,���Gb�&aH[
b��^��9��сX[l���Tq�d�U��,���a��$-��λjM��T�I{��p�>?>�O����ipѳ����)�c���m:��l+�)mD�<���:x>����_���Z�R��[\卨IB8��&4 A�����ޙ�G:��qfN#��X�U��l4@�>͖Ɋ�dI�[��d:�d��XB�ӏ]"d5Hv;����Nm'�it��&�.Y���\[���~�(PdqQX�yZx(�Rm�����BJ�O3/^��r��I�a��I4a<a6�6Q�NA�ƫՎ]ܻ�� ���g��AIЛ��t�y�':l�b����[lUbDX]�BԖ�wwr��;��h������'�hИ2]�1Ã!$'}�����*�����ڕ�_>a�L�ad �(5���gIU�#rI+�i����B�.��e;7w4�Fc�AhL��T�=֕��U�4W��R�N=M���}鱨|t�i�F�fH�L�)zi)5�C��� �hA>��c{����c�R4	��6�ʤ����m����\.n�fx����;�����F��n�W&]���y!$˺a+
�6ݫU���c�'J:��f&8��=�g��q8��ɴ�p~H�4�)�ӖY�f�i)2���i�ITl�vx��<p��!�OW�GhMd��|C�!A�ԼG4Ur��b`�oeUT%i÷4vBB[ަN=��d��s��Q!�	7���1��b|7����'�P���IV�m�8�����軕~�U�x�|�27����8�1ӱ�ڂe1���N&�\gEVJ�	�4Y�X�+��+VJ��Gqc�9��jWǺ#I�_V���d�ILP>N}�$����a���hČ& l�O����>f�H�H��c�2H����p�s�x+9��G]7����}��'<�ʽ^�PnmL�Cj�EM���vJ�����O6�7ި�;ݶ��8���M{�"�&n(,ۜ���	I�����x�5�h�nIF���}�fH�r:�M�d�α�ڡ��K^6x���Z��C!�)��D��QX��=z L���I"q�N�+LW�1sq�I�b�[E��D���mo���o�^�e��@Ok(͒�*�[5�%A�(��hJZ��tKr�-ֈ��-ݶKB��6�C�$D7�g�y*���s��kY�jMnl���u'I�B*�|�?D�:��S0�='�&�i}�<�#צ1����ԭD�I���5dT�G**�PTu� �*6E/�оhyHV���r�_Y��wŷK�,�iR�RVߓf�%��-�M��ov��}�[�Q��`��e�>>~Mlγ��"zYf҈F߮H�9�F��a4�cI����x��6lΡ�HB��1��G`�-�D*5]�*zSm"w݋a�z��R:얢R�j#�0�J���]D�غ\�ͭ�aqj-b�tK���h�CYɲ��lB�"F��$c���FZ�p�c@Zy����:�"S�L�8�L�&-�/6�'SI����d���|��b�zŶu��Y}���z�2~y�=c��O�WjW�>�Ice�R\�P]`�dUF�}�3F̥�H�g���ߓ>~�&�6a��98�>zO`t��uE��K���q���߮��>:}�}�H2F������=Y6��e�AVԼx��6����z���z���m��z�Ǯ=q�\x��m��q��8p�[m���x��n�iƜb�p�q�q���W��*����4��8��ӎ+�w��8���Ep�Ç;|��c��>|��b���/��Ҹp�p�=���Wq��f���F��i�@�A/R	��d��j#���L��*+��GpM��^D$^�� ��إ$�^ f*,YҊ�ݘ��i%�Y��e�t���dwD����W��E���+�C�dO�VC���l,�>�j���,W#ٸ0~�vL���t�����������������������������$ �,z�!�I$�m:�v�4��I���~3�p���U raH�8Y����"|����l�!$�<��~�'qӮ��q)��i<�pr�fn~Y�ڪ���6�<Uv�y9���BaD��=?d%��2�s���8�ݾQ�F0W�\V�J�J��S�G��h�wįHd"a%�0h�R�����+�Q�_��:��ɑ���c�1��'��А���a'�Q�E[�^ҁ�ɤ�<=l�aj�B�V�e�QA�S .%�m���u:�[&���i��|�i<�%��bY�`�	�8�r�0c1�	��p�N��p�'�[N<�#��+�f�FB����ݰ�)M�-&ܿ�:/�C����rI2��!��cv���R���f-*�MFڙl��^�x<MrBa�#��z��f�|�ExB��yy�"�_�����ŝ�BI79{8yٓi�;M�|w�I�����zm�m��#v\�ŸK�d�6�G��A����D� �cm�����q���W�������1r^	{
k��AI�v�Fk�M�kĒM|���$N�$Hu�Ѐ�ؐ��Q��W_I!��Z�g�\N>8�-�ʘ��Ui�SI��d!�1�v�vWl+[�+�o��;%5��p�j'+tz�/;m���˹qӵ,e��I"Q'��w^���6��u:�w����G��uÔ��Υq����UUUD;bu>m:�(D��4d4"&�	��Ϙ����&Y	8�ܻ9'��ms��Gx�*\l+v7�7CwbL��V?��e<R�c�l2ى�A�=lӭ�UZ�d���V[$��u1�$�#���<w�������	N?&���.���6�M&Q;���c-/�=X����j�z��;���׿O��c>UR�&ں�LƱ�:��ck825=b��:ch�hD�}��bH���D��+�w2��;�뉄���cu�_Q�ǓL�6�>u�����j�#*z�ݗuuE��wi�����He븑0��u��ݪ�4h؉d<B��Љ��
3����#�&���]����[�)��uó�'���q�����!7Q�a=E�M��_X���ᶍe�ٴÇ�s%>�2�Me��$,D���2h6"h�k^"*�`�!]������8J�^��\;���#)��t���a cB��=_;"l����LKɧ)O{*BUT�Ґ���Q�dK�"_u$d����'��gF��Y�f�pك�Ov������N�q�8����Ǯ=q�q��4�ÇV�i��q�j�N4�Ç�8�i�q�ǧg�������q\vk��Ӎ8��q���iUÇq^<<<<;x��>u��6����Ϝq�n4���0����2%T���&�Ů��>{�d��DN�{E��3e$��U�y�wZt�����=njes�3r�A�	!�vMR�2�)(E��*�f�S3$,�n����Uu{9�ɵ�"n��L�J�:V�D��A�Ȣ����o����OvNyg:���"��q��М�{6�I��.ͼ����κ�=o4�����|{�ȯJ�R!�U(�ț
wU"{5��w����q�x�2dl[��y$mXj#�s�EJ�X�2M{V�TQ
l����uL`���y����;��ff{8w;��ff{8w;��ff{8w;��ff{8w;��ff{8w;��fflH�A��P��!�O��=>��Z�xvY�l��ԒbYv�v1�u����sf1keT���5t0���c���޺�,��aep��و�p� ��dy�ʹ��X�V�n5��czJ"�HtS\Q�Hb(�
�AEK��Q���&�9��D��\�I�JR��^��S/]IQM��<&�5,�τ1%1��L��Rf����h��Ya!�A�d�(��6Mu�7D�t�M-�}�OxĞ�\�2�X��6���$M���E�]-�)5��t���\�.U�t�N��������&LY���O���:�Mizc���z�qq��}�w�++x}#h��E�E-R�(��)@����3�wy-Sb"B!d�pD�E<T&��V(�@�N�L'���o*��(�i��I�T��H�ך�D��y���GČ��y�|���^���q;�Ge@lE@������"a6��&SFC�BhH�:�e��^B��qY����S"�v�ր�r���Q�x�{������~U�/��Z���J�:�v{�S�&GI�S�c�	��6�W#���]Ǔ�����1|l4	� C����p5)%���<�Q�Q��ؑ�� ��OHƤ�	���;�FN��[P�q4�	��x�q�Oz��R��xl�bS�����v;�OѓK��ƕ[clc6 Ak�����d��m6��ӂ|�y����U%ǳ29G0pj�d�2���`0H�G'�C{�A�<fYOR��8���b�I��VUp��*�6�5�v�k�d����R�U�"b_g���1<��ع�CiN��Rh��}	���w��>p�Y����4�r�(O��s6��>=�їw>��qGh�4K(�'���O�N�^��1����k���X��8����Ԧ�MF@�&�6ƈ�*����s�MI��se��c(;��b��\"#������E��Q�����'�n>���HC�i��9JN&R��M��8c�1������h��9;� B8��$3	ϩ�����-�%�zסu'�1�W���J%��l�����x�'`ȶm�K���1&�t�Φn�BjW�m� �3�1X ���Ց�kX���"��ᾠ�|�yF��㎕^1�ǭ�cz2Y*���Nx�-+�Q��82A��K��%EU��9R`��L�S5��<�}��I椄�BB�1�����0n���6U���3r����ѹBb�P�&Hl�'��A� �_��!�[�-�tn��tu���-����#�ڛ�ת̌ȭ�RT)[]KmI��J��XB��TcA�m)�l�k�`���kL��i�k�ڵZ��E#0໊b3���K�z:��l����j��T$KOY��~�K���'{��N�S�0��ɶg�LS;�����Є2g��3�;n����.��8}Mt�D���m�Ӷb�V�����X��*���O��bm �P�!'R�I�ƓŜ(�Ox�d�j��)-&��R	F
����.��Xn�S[�J�!(�ܪ�:;CCf�>x���z���z�m;v�q�׎8�ƞ��Ǯ=v�iƜb��\8p�m��v��n6Ӎb�p�Î+��q�ǧg�釧�W��O�8��.8��;q�<mƕ�8p���������|����_/ϟ=|�8h��@`1��Cf��
 G�n2�V�IC��PQ¦��Gv�n�OT��/E^"�$��Ff�Ⱥ�Dn�N6��zn��ꁚ�f��!�M%�Lڍ�Ϻff{9<;��ff{9=ǻ��f{9=ǻ��f{�.=ǻ��f{��ǻ��f`H �HA`�h4PPQ��J&�t���I�%m�
��6h�g5�O7wukm�i��:z�f�v���a���u��Cp'S:�ݾ$���2p�V��ǭ�������b�wFe$�h��\�CwZō��:FFj�R��T�����ݎ|�	�E�RRi޶B��$v�5~���i"s��OnY�z�<x�[:UW�t�1�ó�c��g՘��HRS����0j����%F��`Jg6���[����=�&�']�53�tK�,��.rM%�$�se�K4����|ƓI���m=�IUUTM�K�I��ӭ�N�z�t�l8u0�'<��)�z.��d�oD�2�@��2P��E�T0�b�w�˯xCE] ��!x�h4@�판���ԇ�2�ry�)�TJ��Ig�4c:3�_c&�Gyk��<~����x	p��U�T�]3gWغ�7=ͣ�!ވ��h�2�[���n��n貥��b���2�)��I�յ��EQ	O@��D���Z�~v�퍱�~6m���e�ՑGK�at��q�|�؊j�0���4Cd&�a0����,�kټl�����d�(��s��(�&@�y:a#��8�.�HwUD��"ўk�Z��������z�6W����W�x�1��c]W�K�$�SGktp���>�d�.]���d��+J���Wa�m*'X��6ӛ~�lN�N�8M��@�:�ˮ�s�z�2�jBG��-_'�'�>��q�J���Ǧ�M&�F���B��N��c[�p[�5j��q��/����D��[nr�:�L�)o�t��=�V�Q��+.��*k�aI��%���K)k
)$��&���ɛ�۹b.Jc�����TyI�3F�N�M��޹--)�/�'��M�L�ģQ�$eɪ��w��1sׇ�A�M��[Z�J�ve1JLK����������>�d��t��VV�lЉ�!p4a�;�&FNN�fWl���l��K�0��e)�d��m2m�e-O<	�<��(��2�7!F9,M��1/�b�c]C�1�6V���wGۣ(�J���x&�U�Ո��Ј�a���	Y>��τ���v.�oRY1!
�e6��O�6`����6r��X�G����榬!�m�H,��l����`<S��u�q���p�0����$�2L���L|�1��l0ÞM�ˍ���[
�j������X��{3Z�e�m�����0~w��x����*8~z�KH�Hn�B0�Ǔ�N��]&KJŏ
�K�e����V�o&��������)h_ª������Q�����?�?�8`��	?���ke��fih���G3�}�xKa���Q�!B��� �X{p��a��%"�E%"bT�PY%IIRT���RR)(�RjY&
%�%)%B�%D��E�(�Qd�X�X�kXF�E�(�Qd(�%J*E"�%�*F$QR(��T�,�E���(�(�(������QR(�QD��Y
(�Q(�Q�a���E�(�QH���$QP��E�,2�bED��QD��QD�ĔY
,T5�T�(���QH��QD��E�	a�#(�Q����E���EH���F�u��\*�u�K��i
,XJ)T�(�X�*ED��XeH��!EIEI(�E"�$Qb(�QIF)�E��Y%QP��R�%��J)(���QRQR(�EB�E"�P��Qd�,��IE���J*J,)%�E%�Y"�B�E��!ED��(�K��E%B�
*J)(�)%�Qd��E���Qd�X�,J,Y
IB�E���)Q(�Y
(�P��J*E"�T�,EJ,E"�X�Ċ,��,�B�%B�%%"�RQd�Y"��E���Qd(�E��I*%%B��
(QI(�QB�)%�QRQbQS
�r��(\�FE(X�e!b�h��Ab��,RZ��B�%�,�i"�D�B�D�D�b�2��%���,�YRZ�PX���PYIeIb�(�D�K(�Ih�I-%�,��,���(�E������QeR�,RK(�E�X��b�Ȣ�b��$�E�X��K��,RZK�),�,��YE�K)%�,��-Qb�e%�,��,RKYIb�)%�X���Ie(,��YE�,�,RYEYE�Ie(��(�I,QeK*�K(�)e,Rʉb����YV*%��K�K(�)e,U���T�*X���KK��U���X��dQh*E"�R,�"�R*E"�T,�I`�,E"�H�aJE�H�H���!H���H�R:�0�!DT��d)
EB�R)%"Ĕ�D��E1C�5�j9�_�.�4%	���ޟ�~� �� ��� F!�RW����_�s_�s������?G������3���������/��?���!��?bC�������g��&��!�?��!?~��E���S����O�~
O��?��?*�������������?��

�0���LUD�)�����������?�C�~��Hh��)K�x'���� �~��'��?���~D?������w����h����$�ih�iC�-��p��؟�4?��\JJO�M�~"�4~�k|tn�'�����?F��b�����\���oE?���Bt�$�$�C"D�T*""
��F�[�B��k�]�U���l�`>�����p?�
 ����T�-@���'t$�*�$KET��2�Y�������|&�����'����G�ҩO��&��R��z����?����Z�����QUD����%���Z�N��;�g��������	���\A������������!�����G��O���M~�������?��c�*���|:����C����1ޛ:��_�L@�?i�DUQ?7���9�9�C�諰?m�P�?i������lh�D���1����SR�?��ϑ����#��ӣ��d\�C062���)�?=hN]������۵�\#�'��z ��6N9V��_�������"����e�I�D�O� ���?X��o������O��C`����]O�?П�)?P����3����?�Q����H��?�'������?�~@��0 ������TM��L��?n����?�;�@��ҟ����'������w�n����T�Х��^�4д3����@�E�����~ <�!�w"Y�t��.�8�0Ȋ�&��$�A�G��gQY����G�'�O�14~�G����6�>�H�������eR��x�����'��s�O� ���?�~��?P���:O���A@?@~��T=��5.�ݽM���������į�C�R��=�M���?��ܑN$x�@