BZh91AY&SY�����_�`q���"� ����b)                                            *AH� J� }M����<�   ��  0�   �  ��J �      P @     � n��"���UT�� ��TQJ����E�P�(�)	J"�((�B(��B����N�!PJU*@*�T��� k��w��)�w�����۪�<�C�=(�ý�b���a�[�<��n�j���B.t�;����z�   }+�#gEj���6o��{��ej�j|�}�U�����w���7"���� z���9�TU���M� <����Oc�` �   u�_m��$
QOEU$�P�� 7��c�� ���C�����q: )��JRpz݇�����_@{� ��}� �=誥�v:yh>���   �u>^�k4�AY�w0�� ���(< c��O�}`s�����=� y����c���9�p>����� > @ Sq}f�0��QT
H�T)5R��k��z�}���� �}瘝�����ǟm�9��{� ���� ��|�UW�>�����   +�}&P ҭ�r ���� ��P��:�� w��}}�X���]g��� Ǟ�=����`���p� *� <}/mi%(|H�)*UD	Hڪ*� >��������py w�����O 1� d�wX��w�<�� x�S�	Pv�  Xy[1�T8l��������@�@9 ���`t��AE�{�<@ʇ� r70 �� 
����� �RUTD�J�B��*� m�ҁ���9W{� yw�$�k b@�`C�� z���� m�y ;�  P��>�kZ�%x7��2 �I}��z �`������=�Hx ݇�)�4�`���A�   �    O )TɦL  F�S�"RUP 2� 44d��O�*�LiT�10&i�i�FCL4�*A5IJ140C ��a10��F���H�@ � �5�R()�EOh2M�Pi�2oT�䟷��~�u��ģ��ꂚU:�˶�^��9�7����*���`�)Ï}�DTWЊ�
���*+�����`'�����ҧ�TQX?�ʢ?� ����T�)AE��~߿��Q�2��`���
8�.0��2 c(&2#2(c*�0�c*�2#2#�"��������Dq�^2�� �������1��
®0+���
������
��2��*���.2+�"8ȁ��Ȯ2�c�2"c+0� &0+�*��0�1�8Ɍ�Ì�ˌ�Ì����0�0�2c.3�a�.0�2���0c2Ì8Ì8�qǃ�a�e�q�\a�\`1�q�q�3��a�Le�Le�q���q�d�d�d�x��q��a�a�fcq��a1��Y�dq��e�Le�\`���d�q�q�q�1��q�1�q�q�q��0�a�a�La�a�\e�q�q�q�q�q�q��1�e�i�`1�a1�ƙ1��Cq��a�1��S`1��/xÌ8���Ɍ�ÌLɌÌÌɌ���2c&2c2c&0c2c31�8Ɍ8Ɍ8���Ì80���2c2c.2c'x�a�La�La�a�a��fLd�Ld�a�q��<N0�0Ɍ�Ɍ��3�ˌ�ˌ8�c!�&0�q�1�q��1�1�q�1�1�1�Ɍ�d�La�La�1��a�Ld�L`�d�gd�`�`�`�Lg0e�Le�d�a�q�1��d�L`�Ld�L`�`ƙ�L`�La�Ld�L`�LdǏ8������Ɍ�ˍ�q��N0�2c2c&2c3���Ɍ���8��Ɍ���2c&0c&0c2�38Ɍ8��8Ì�Ɍ���2c0�0���Ì��0LÌ�Ì(L��8ʦ2�2��.0��� 2���� 2"c8�	0��(� ���2��8�Lc"8Ȏ2���� 82��� 8ȤɌ �
��.2#� �8Ȏ0#��$��2��*c
8�2� ���&2� �!�@1�0�
c(8��2�� �
��&2��eW��c
���0	��� 8�&0��� �Q8ʦ0��c��2)���8�<eq�2)��c 8�0)���(8�&0/� ��0�
c 8�2��"�
ee���(�����(8�0���*q�q�N0��*c
��0� �"�¦2�dT� 8��0��
c"�ʦ2���(a\a���8��2�*�"�0�$Ȧ0� � 8�0����&����M~��?_�>���k�"��ON*�I��Z���+�O%�T�A�ݕ�4�̺V��ݚ8E��D������  �E�w L�r^�Ѯ+F��M��qUz��U��{�@>n��ܻ!�V�&�74	wnv�Q�]�V=��2�Z����X?�݂C�����E��1�gEK���n��<�'���q��f�h��u����E��n�K���g^���Bъ�հ8p%JuaY����q
�b\8,�;[ˇ	�j�_sd��D������^��j��I�9P�^�K�K���ڛ'|e��/l���7���9˚��OM�U`����گzov�(��j��d�ű�h������蝋d\�pWb��7��t��8u=��קo�GH�^�To��� �b�Q��s��+=��]�wu,f̍�p��\��E1k5��ҵS���ߺr�ZLc���rnqɊ�m����5t����׻���V^�eG����v�ގm�j"�-�#�n��Z�sWR�ƈQǻ��4��왷�LVgB@Lv*��w8�}�F!(����L6)]�([��`�o:��M��si�i�8�u��n����Vǫ�=�3���;S7����t�"��ݥz>ޝ+眻[�+;���pl�U{hAcmx��0�����i�扂:��v�x�7^���]u%~ް;���ؕD`Q7כ���Y�x�wu�#,�_v�y�L�9���)��oh��>�:C� ɿ6{S{�]�Ŝ�o{�o= Vp3f�\�EM��O�o�I'%�ӷ��;��;�b'fQ5ηE�Щyf�x�f88Fj�7*����N;�%�E�`sM����PmQF,3y����P��1�%�כ���[��Om�{j��~k���싧z�ܭ�b�� ^3y�Ɉ���.�a]�ˣ�i���2����Z��N�/D�9����d0�J�Ѩ�w/�u9as�cOtz���L�UIF�V�gN�[]��6�z�郤B�� �T�u3�!�A\8��Շ���v{ �48��֥xM��q淢�� as�K��l�}:�v�mY��I����k�)bFsEXwRE]^�a]��#���?P;��[F����݃AӉ����}��N̚z����;&n�\�q�;G/��${[Y�Tr�0��j8����kё*n;zs����l����R��u24��<�G5�En	�^8z��%��T�pDh��7z^h��fK��1�waȗ���^>��,ӻ��44����I,�:p��I��r��u]D�z�qszv�0Rn��^\�kwU ��t�f�=f��`�V�=U�I0�6� ����ROy�0a�Ȗ3�*�|DAjH�5���M�w�A�q3wIשP��j�T����+����C����ޚ��q��v�<�oVq���25��6YJ웸{��WA�:+QX�o:���k|
���X�b�I�\;S}Ϲf��N�|�Ի�݉
��(Kf�v�)�0�6�+K�fq47.��H��Aӽ���+f����:Vm��=����g	���(QwW�>Û��gvo�>��*�É�����1DƧ�+:� sw�H��o!���S;4;M.v)�ɸOc�Z� �}�5hi�@��rwx(_ڌ;�y�y;ܬ�VLDɛ9�0�[v�R�u{���9f�n��������Ճ��~���q�h�0�9���䜻�͔5�Ju����u�����ߎ]�!Q�k�7u5 +f�@j ����3b�.v/��V�};���F�m�;�8�%ɂt��p�=��t��cA�+�.���Ť���{Y�6��cFN����8�{�ݲ	j�y�]�
�1v���A��`�L����9�m"�O�X2[�\vv�C_�Uy��.��TS���L�C8Ov���K�Q�7c�j��M���N�7}1ku+�n�Q��lr�1w��Y�Wa\�����9N�wkz�^��Ձ7½iŸ�8�^Ggd\��6^�6a���1p�K,s�&�b��2�8	if�����16=�+�^���
H�2uwٸW��b��-�����(��z��FM��m�v���ğl����pj�x���7b�h�X����	ۭkÅ��;˂�f�{���Ք�ɼ�14.\źP�)�ؓ�s ���s�H�4�`��`Xe���9).�cJ�(�.c�n�Ȩ�����ۇzq�Q�oxы����=_�6�Þئk�M�or܃�&D:���-)̽֝=����@]��#�PQ���v
@����'q^%���5f��!�@������v=*U����v�'ϑ�;:�f����z؂�7&M����d#�ǻ�&�3����޻���!�Z���n��l,Vrc�l���k�{h��4�wF3���5݂ŝe)t�<;{������!G�r&q��N���(�\7r��u�VwWF��@�O���o�=y�A`j��'tjfb�1����:����M:,����4|�F1�w8��Q2gYe3t7o<k�9
i�7Dlw�зa�Ex�3J�W5���WwM��e��.���P�}N4.h��o�%�M�^lН�O%�ld� m�sn<�iB$�n��h� �q�E䮹;Rɴ�Ɖ����zWnq7�c�ꐫ�f
�`Ӣ��Op7�!�[���O(ű���vR�2t.�ƙڗd(%��j�be��\u����Ó!35�+�(
��%�:�-z��oZɿh%Y����`H}r�#��Δ�q[fL�7`��qe��i��H~x���Y�ݺ��蜹�`B�n3Rم��4�q��3@�uȊg,�oj��gx�*D����9�(�pvL�v>��Xr���}@3�V�"<N��a(MߛԺ�#���mS��F苹j�X	�d�Bܯd�
#�lG������okf��u�%+7��(�����.<ov�s^vM�]�*��ۚ�@T� =�;Y��;OGX�����$��uA�w��ά��ɳ�&ו��Y#�ogJ�.��%.�t�w�,�(��aD��l��F�y֧�t=�㝝�^�"�q�Ggo$@X>C�K�)ܵU@� ��C�ˊj+'\ъv���I�}qn�#�#��X�nv�����^3���9��(����ҵ�I�"�eؐ}���;h;9�8u�N')�3z��˳5��Y���u����pW��ʁOв��:��k�f�Pj�`���{P�8�v���w	�;�T�pu��I����\�)k��rY�P������r��}�evܖrj�.�]�DTf~l���<� <R爌��N�n����s��;�M�Y� ʗ���q-�L�nohK��;2��擼�U�Wmz;��ҹ��yP�&��Ӷ��8��d1�.a�P����	�ëGaC� OsUÜ7vg-540�d�ٻ�|���.:�ZY*�2�	]@��a<��d�ø-��U	t�x2��T�2
�i��9q���G�������u�n���*j�WN�4%yl|�p��{��a��G�L���XN��l�5ҧW�6��?�1���&.w�Ġ&�8f�z���ֻWZ;��}8���A�,ۼ	�Dh�� Zt��;6��rh�˚�/1�:S�9wP�=*W�wg� 7u�;ܖ)�G�+�SZ�3� sn��_�{�V�^� 77%wgi���r`�1����s�#��c��tu+7\�3J��;q�lO��#�h�Tw$y�k:@��˕,,�/�]�ZJ�0���^>�6�J�p���([�-�3�t�άîܐ^�nܣ.ʞ�ͻ�5�ݯ�%��|L��7%�#��ˎ8��9w8���t�`�lU�۠@�%�E�S���Pg��9���Q6�;q\�mq6��ٮ�&�2�J�4�;$n8�;�L�<���Q��6D����b�78����׷x��0� 
o7f*!��d�c�nGtn��̏A�81ظ	y� �ċ ���v����)���_��:x��.v����:��dk*F �������'��0���ۑlI�C�s'�*����ѝ��ι�q�Ko�z�ܸ7dc�Q�S�v�	+;]Y��	*�V�#�x���Z��L�Hڢv��Pw6쐀l�ٯ��5r`���)�|5����a�[9��i-.(��o�D�\c�T������u�b/~���.���/jtt�靨��	Y;acY�oj�^��^t!AeLv�g3�G��V��p�v%��t.{�wp�iZ̹9Yn�# �(�a�{y*H��0��zG��]�6���Lu�Z�������"�Y�w��)��mX���뼀(�XV=s���9^��q��\�c�4cW�bb��7X���+㻡��[>%�;L�Vsr����%�C����I��s���o�=$�{:��Б�b���G�hXN^q�78ڐ�����u���۹Cј���i�"�聳3%-�..ι�>y��
[�%�K9���nM��c���o-/�P᳴��V��ӂj��3Yk��xlM��ܩ+�r�f��/hxs�k��[�t�JL���9\4��$��j8dx�'v^�b:v�x�Z�]{u^�IHͽE���3r���poSpR��[�]Kz�#�j�ے��9�7^���8V@Y�{�Ұ����j�C� {�k�	-(�V;d����A�ڹ��)��p	�vf��k��]��1Uwa���rgj['����NבW���+��(G�h�CsD�^UR��p��u.�o`]-'gL�N�;�.�n�\��\�1t�:���Ow,���וlD�ΙN;�+5��7n�����Ҿ��EF�j�*�h� w�Y���E�A��}����M}�K\����@lX�⑈�WRH濔�pΙ2��ΔB!E*z�S;��W��I�m����.u�i	F2�C^�8��=���	a���ȸ�O���;��8��s�NZzk���ES�\���T�����m8k��^�����9�l�+_�Lޡr!�p�,@r��ߎ�ɢ�����]f<o&�'v��U���軻�=;�r��wk�2����ס���������詳Or��7P�hz��l���6�9'1��3^U�$XÛ*/��}zpfv��P�!����mո��h��
����{z�*|�<�h0�f��҄)�PN%�4�.�8�9$}�qO���[k,]��"�$�=�^��f��+4M�'�d���_���#д��n�px�^�(�\RÞ�ӘQ��! �7��ܮ�7��#�
V����yX���.�2�>�TWo<��Ʈ�0*`L�	�t��'^�(�p�(�i�=xv���s�ή.���ކ�-�J�����z <�u���F�����tl�sA��03�&�FX����8��5c�8չ&����	��٣�1�٦�������|��p�����y�u����S�{ľ=�c��g.��g|Nl������D�on�Z���F��^w-S���.y��ޏu��1l+�N2i�i��֎�o=���n��Gk-K�8�.-�;m�OHf��f�LM��EV�j���yf�oq���,#X���7�=�1^�;<�#TE������
��l'��)��ݗ(� �e$o�y�Әp˵��"�]t��h�´��Ǉ�I��҄�v%c��z!�D�-�J;''���Q^{v����k��#,PgB��ǃN�Xg�n]��{A�w��G��E�{z�_j�"��e�u`c��bݺBq�V�����od�P��3�����w�A�ܑ�Y�0�{Z��`u\����Ν�c�ڶ���ѭ�LѨ��N�`%�V9��um�� 	҄�`[�7�b���V�Ӹ貯���:�ɺ�@��;��D:K'�Z�S�0�%k�yf"�Nl�2�Z�ݘ�O�p��ж|ϴ���y�h�j��u֧R�T�R�MK5E����V�-e�t�\'�FTR\�ӂ̢����i���n��<O�sq�a`Ix���K�<�f1�nH[��g\�~׿�u��ם>��ol}�e�_w��O��q�5�PӰ������ID�[��-��^�3Q�Ǜ�x�Zb��m�O�S��PϊPn����P��F�!1�����ꨞ�B���絇썾��~8�Oq;n1פ�K�UG��1�uכo5Q��*z���]VóLnΖ�N1�7.��_wg!�n����kkX�"��ձ��X�A�Z�Ӵ���b6�����hw����C̝������j���g��=�4���d��s��uC�� h���핖�u-�����g�y�ܶ���%�8��O5�e����ETSj�P��i����^�1΍3t�nk�%t7����{:c�@�G�  ���w�#r�O�>��;'d����N����A�a헡��؈�q��&��#��^�{y1��k�b�8»�����\YS�M�Inȿ������1=�1!����O���d�[���γ�]��:z�}&A����N�<�ћ�}��wE|g�[��=Ej�Oݙ1�TӪ{�ɫWڵ�/K��/2�$���{��lk���̦�z��/��� �f{���t�����
�x�ZpUhe���7�<��4]����1�ڏ䱌����m�(�����i����a�J{�mP�#"]�[���cŌK���9K�&�%��r������	q��"�>})�*KRt��J�Jk[VcAt�;�ض��KR�2y6R#�7B��/��&r��^;�Ă��3�#E􁟡:����V�t�����=��ݒB?��~����^��D��P�A?XU9R �BҢ�ҁ@�@H"P*"�R(R��"!P9 P(Ҋ�$S��B*�$U�-(� ��H�Ң��@<�9�BrDC�r@�@�@��4��/ Dy
�B��"�W�+@�P��*�B)B�R"P���Р
���9
!�Ey R��N@�С��4������
%( R-(*�(�*� �(4R- ��@)EJ/$Q�(DZ�
U-Q_�W����,h�3#���Ȧe�;�>nz6�ܒYq��9���[7O�W.����*��5v[���!�]n��Y�ht��؄���X0ñ���X����N��E���M���'R����Dz1�����3�ff.��:|�I+���S��	�,�j�̮d�Y�G7����r�j���Ie���L�Ւ��"P��7��՚���KO�ƍ�Mܭ�z�o[���FO.;BjP7+r�|�ڴ�Jj�i�ދ���@������1b�����%%��֡�B&8{(��±5Rx�kxB����ZA.J��n��G�.�G�[�}� ��s��)Nb�#n���&���{���� �1ñC׏�X�a�!7��/_��e⁼�QӿK�'z��;����l���7��t�K��S�ղ�rTKh�J�W˅חZM4�P.&���j���\�
ƍ�i�E��Y��(*���~���:���o�;�{�����_�������s�?>�˟����:��[u
��]1o�[@��ע�劓�;�����-�N�2UZ�,�;������;���{y��FS��ٖ����CV޷�"��&�g�rcer�4��/{u���ErɁ>��	og��&>�2������`[�>~��䞺��s�4nY�^�v>�:/e�(�{Vs�<�:��j�w��/n �΂k�*ڢ��;�>:G�����g��O�#�1ܡ��w�L#�7�fn�iλ�<Y���݆7��1��N�Aa6ļst�}l�//+�]38̘Nn��f�6��}�wM[_��]�}���v���gzxދA��޺��۪kq���ң���g\��{�����J
�����x�Y�.�W���:>k{��x���/e!zOxO+���Lq���d��xg�^���9'�\�s��ſ����9�a�$�{�9�V�b�X[�U�Պ9�9���K�!�� ���=��=\�@�L7).V��0�{���P�)KȎ�f{�nL��{�-�/��^�Q�r��9˼��&�L*۬w������L;}{ȏq7&��;��<P���s�~��D�C/L/�}��C�{	�0ӓׂ����׷g��㮺뮺î��N�뮽�:뮺뮾�u㮺뮽�>>8������ۮ��Ӯ��u׷^�u׷^������u�\u�]u�Ӯ���뮺�㣮�뮺믎���뮺���^:뮺믧]u�]u�]{u�]zu�^<zq�]u�Ӯ���뮺�㣮�뮺뮺:뮺뮺��:뮺믬��﮼�t`��lf�O2�<��k3�{}�ڳ=�ϸ�0�"�{���������`����d�ޙ������K/���O�ݹ�����QL[6h��3���2����
f�>v6\��F_3��֢�It���8��<4VL��ݶ)RSy�v�����2c�IW������1�L�i���Q�4�b�e��y�ist�s_}�
�[a^�Ԇ��^�q0Ӿ�z�[SM�>܏5�b�\���B���{�@�M6d�ϑ3K�]�~����Kܚ�sM��M�=��l=��'�]��'D���p���mw���I���yw��l*	��=�%�#��=3���֬�&E\���"_��t{;����4̬4��e6蝒��s��a'�Q[2�^�ݘ|�o�f�g�NxN���_�w5�����u}�����r������,^����;`��� �i^�"���$�p��i]������8+ꌃ�Nm�.{��P��C�yS�KD9I�z��+x����3'�0�o�,�Om{�YS�i�����}�d�3���|�og"�
�7fOU���������.��ݲ���g�PC`X��n����و��{�����~9/+��1΁y�Ώe��}�Y��b���L��Ra��{w����]��Ӯc�����O��뮺믧P�]u�]}:�:�u�]u�ۣ��뮾>>�������]u�G]u�]u�뮸�������]u�]u�뮸뮺:�뮺�ۮ���]u�]}�:뮺뮺룮�뮺뮺:뮺뮾�u㮳:�ۮ��Ӯ��N�뮽�뮸뮺믧]u㮺뮺�u�u�]u��i���Mk� �������j��7(�-�rY��2UTb�X��ar��|��5o{�g��3���-};���
E�7=:rk��ҹ��Q�ӷ��fƁk��;�!��w��bݿ:JY�K�}��������St��{���9�|n���g���1���������r���%�[�&�cb�7�~n�y^;������b�/�y�4}��������g���N��@u�cp��v����}QA^��v����	�׀%"~��RNe�"emԮ�����eE͋ӧ+곦q�7ǯ���O��8O��}��&š�G`_V�����2y����3w���r�
͇�� gg��oo��G'����]�Fw=�I�8����C��� .�Md��u���L$Q�ǌ76/`������/ac���<u^՞�x���Q#� ���v�.���/_>�Ր[۝pޫ�G��7;,�r��0��
�z	�}ۺ��-^���w��{ٸy�R��?w�{�na]9��<��Fy�۪{�Ϩ��ô�W3Й͓"g3��>���n�b�	>�����$��8�:bc��<�4�=��JY�I�9�&��p�5��<:y�W}����k=�e��{�^>�q�>�o���ۮ��ӣ�뮺뮺�뮺�n���=:뮸뮾>=�>3���㮺�㮳��뮺뮳�����ۣ��뮺믎���뮺���^:뮺�ۮ��Ӯ�뎺뮺�u�]q�]q�]q�]x뮺뮾�u��]u��Y�]u�]u��u�]u�Ӯ�㮺뮽�뮽:뮺�뾷�LF=��:w�Vl��E�Z�*T�;WI� |<%z$d\^��v[�-n��!7z�zS��|���"�]^���+z���/v��E8�ۗ��<>�fx��qJ�����O9r��MLp�{x�->������0���]s��:C�?y���}tX*Q���l 4�o��Go=�f�m��C�3w�+	�9���=�� �
���Ź���9Ѥ�dv�{���x��|�[��"}�giϾ:���K��s�;���Y7�`Y�_w���ʭ~�u�����}|�\��q�̮��Ư���p�~��|���B�
y�ݙw�\�i�:)>3	��o��ץVHx1=����v��1f{r���+������z�3tk��B#�-��rxK��-�0�z�x�.{�{]Z��y�������w��B-bU{s��x2txJ�c�7=�;pc��z�y6;�t}�M:�;�]���F��I�����Lf�ٽ�0
(�zt��K�����5��F�L�6b"c��1���u��}�,ٜ2cŞ�C�{�@�(�Yv�|n��gn �˸������ ���f�B��s}ޜ���j��=G�<Ϥ��9ng��"�hݚ<��[Ԗ|���*E�Z�E�q�z�ϥѸGò-�&d�U��}�E�ݩq����"�4b3�a<�����&_u�~�C�cN}�]��9�܃��1�r���Բw���<��%��p�]�^{���5c�*�D�JdyVK�c�,�䜣Y 3��l��S;��^��˺��_`�_�q�{�R�Ԇ}��~�^?_a��F�|�y�Q�cw_��6wް�3'���{~�w�K��5���Y�M}�!�v{�ki7�M����k�+��2�!�>!d�rlY�ϵ����;�{�囋��*Ț���}�y��#0c�b���=��n��gG�\�S�Ogv��Di�y�=|�d+�@}�7Z�8H�dJ�MXV*���ja6A�Q
׽��l[t}�CvHh.��G9��)��Q��;��(�>j�� �a�ug]���>�ͣg�yd;�6\p/e�+���g﷗��䈏Y���v�}v�|�������W�0#��o<���+>z��3+#��sn{��AŪzg��I�~'
7)z��!���jC���ѝ=����ֲ�eL��ϸ���O�9_f����9�Yٝ�ㅽ����Ce�w��c���ɾx�Y$��L�1{Qk2a}N{ˇd:y�y9�-�e�f��ßVB��F��S�ܩ�y�%��+��5o�����3�,��*7�RV��r�oޝ�L�y�@rv(XMks���稿+�ݾ��1��䡦iR��1�q����
Z���"�n�k�Z�V�Xǒ��p����j޻��h��ٌ,kV�f`��｝����(l�ÔaI��D��_n�s%���G�Fu����nY��lR6�SN������������޳�;f�[gl����N��;�!�3�����ˌwVn�T7.�pɞ;�n�q�3�y�����w�^h�}���G`��}<��]�VzT|L��z\<�����hX���ߌ�,�E������鞷:ϳ���{��϶�҆���nx�rl�]�?��,+"�2�B�NU�T�j�<E���δ=U�����s�6\�'�lv{4��r�*��=���Y��@������YC;��1׈��V�����;�=4/�3~�m�I�����n�}{�k�-�dP��>Ʒ�o���m��#S�;�s9�}띱9ˡ||�׍�n�z��ʻ��/CH�M�����~^왎�y��7���h���4�f�,NҚ.����֕���>���7�z?&�(1���^��~�3����/V��қm���3}Ӣ��g��kX����J��}��q��뗞�MY�i{�2,�f］��{;įL9�����4�	Y0{�x{s��ܻ��<�{׍�z��VH�׼�3��bЯ�u�f��pOh<}���Z��X�=�G�s�[�������f�7�����>͌O�\������"ݤ�ӻ ���x4{4?��!7;��_���،�6�}��������j]=6Y��s�y�BOء�BK�+���ox�O#{�ys}��/�w�Nz�T�w��r�bQ;(��%�%��Е�����vo��=�!ϫg�3V��K����h�!�1xm�>�Q�:�c���Dk�[ط���r�~���pkֶ��+��PP����=���r��c���riԌ���z_,��1���5�^iγ8_b}����z�V4�Bf�1�n��рT��1r�3�zz{�&-b���^]�j�=*�u��7�{�����~�	���w.���{fm�o���N�t��e{7���^�bW)��꼸��b鷐V����}�>�l��3��{.�sS�Ȱb��37<t��9��E��y����4�(?1n^��{r{F�派��ȿ}��r���F�3�V�=���k�czr�8�g7ӱb.�"~�o���v��<�h�rf^��#�H�j�r�8���K9H_J���W��'lp��]��J����$����L�񹷽�ˬ�~���x}�V���R��;���gG��g�ы��p�&��jm�w�@BW��Xn��Zأ6T�%��6xL�nf����3�>�]<:L ��C��h\�[�����.ɛ/�.Vg�����R�w+�d��`@l�4��o=\q��g��[�Y��F��\5u��^�DW=�(���=:H(��/s�^#��{˞#�����]my�Rb�7�}�턀����� M�oy��A�6�v��{Wg}�w���qz�q�;�8�v�=
Ei-x�c��G����ۦ�7���/b�|0&��T��x�,Ԃ��,s�P}��̍=�����}�:g�Μ^��7o�n�~�]lc�3���7o�=>s����6��F�_��nX��כ���n�ޓ��g�{���Iz�0�ޕ�p�����V٪E��ސ�+gb{��m+���|�	�Qj^p����]:z���6�^���D��ެ�e�/��p��C��;ʲs����汾�~�_�s��z16ok���o�WQ����_/�W7�Q�io��Ky�>�7��T[xd��ܸ���G<��>ř�d�S����Fm�k2����]<4�<�>�rrP̣/��ݶ�~�'��1�-��2}Hž9rY8�|_�u^�3��8�f��D���8�#s_dHt���z���H�u�vt
d��n�W�M�!xCѧݖ�~̙�j_d(�]��<>~�z+�b4M�1FW��g���nN0�3٢�s+CߚC�3yY$�AuR�@- �����]��t4�A���Űꗱx�MB�yTn-�(I8��Vk^���(7�S�y�.�%��- �ɖ��_��{쒤����2�t��4:�%�wN��w(����a���n?<�bc��/A�GRU@=o��sݽ~�g�PI�{�]�}��0 A�`��4L�7�=�ڐK�pPwn��}7N�o�[�=n�|�@.ź�]�i�������������o_I3[�ػ��Y�����i�#����"�$��w�|�x�Ni�>��ؼ�랞\�ؼ�NI���7�yA|��V�g{��>�ӎ{r^jlݛOR߽���A��Ov����fͷ�.����Q/Sxf���z2��}�z�k����qp�)�o�yߓ���7g���,:�ٛ�Q�Gy�O�Cl��B=2���ٺ�]�K�B��I���7Pzt̙�T��k��}]�����<(Nq���wypV��v������9_9͗tvI�/f���f{���q�t���{!ѽ׽��Ѹ�����x�0�]�<��b�������ˑ���%y�Tγ7N}��xC���>3(�e��vY��yr\,�{��:U2����v��o��MΝC$�_f��%>��/�� ѓ��th�Vb�rb�W����:o��[�����{<̮���PϽ����1��rI�8upٸG�C*�"�ޚB�p{�� ;����53V�'eE����w�o���_��Q�=��.�'%��Ǳ���r���=Z�;�M��îo��yƆ�G�4D`��u�üv�{�ɤ�y.%�{G)=�:.r�E��ϮV���( b;�E�e���������y�r�9���=����Ǧ���B��r�[�Z��;�$|����h�g�<T	.��U�}�4�x��8�κ��-�j���ؽ��CX3[�A�o"
;�VA��7/=:no�p�^G�D}����oQ]г�S|�{U��Ě/wnnw/h�o�8G琛�ެ�%ŗw�̻��{7#Ry��{#����g��]�b1c6+�pVUZX͊�E!s8�3/�7�H��o��{6K��-;���>�{�=ހ����Pkҏ�v��}�"���:$��o/]kw�xw$���SA���l9n blb��w�Z�S�;N�[��/)��pq�z�է�Y��u�a2�f{�ǣ]�%��fÇ����;��eP��>��ۭ��p��'��9� p�4$�`'|Fwo�q1r�3��8�c�}��<��Og�����{L��ن���a�w�_t��r%�۳��sxp��F�|�9�c��g�Gs���-`;���ok>腦��8X�[��^(_{��;ï�ܭ�e�����}��B:._������������������;����W�������7���r-�MmY����$�ZV)Vw[<E�{qe�9�>8wǻ�!��v�^S��������ϣ�hp����#�y�],�u!�y���᫰a�k��B6j�j�ik��������7��o95��&�2���k��+yc����~q���u��#&ӔՒ�۱����H�ƍ�<�[װg����)�V�.��71mc�M]+����t�7yC��o3*�⁠Y��r37kX��Bd�9L�z���F��Ig\�|۱����l�m�s ��'nچe�ɚ+�՘֢E��GM�j\9]h��e�ޥ�7m�	J��-��-�9�x�
ګu�/p�n�-�Y�{nwm�Eu�<gA�Tk��K��vx�
��	ɻ���az��J�\rx����unF��3�-dS��rsl�f��������ö�T��<�l�Wv��-���R�cV��T��:�����+;���#Lq�5�0i�#�����&�x���P�m���C� �dª��8Ii�i�w����M"�^Ս�v����푸�t������+��/n�mq��+��C�c�,Jڞ�kG -�k���vή	�tb9�n�m^��V܍\A�˞�l�'���O[�b�Vɼ��us�3�U�8�Mƞ�{���=.���nh���j�ݞ���S�|[��'�@D��)�(} �1��+��N;�8 ���޶�Օ�1�t�X������hV۫�rѶa�HXku�b�٘�&V�akmZ�a7,5-��GkO��N<=i��6�.�sg�s�n8ٗU�#ؖ.�d:�B�]b�JJX�2�Ջ��Ԛnݲ3F��D=N�ݩ�%o/8).�f]2l��]�+����݌��J�p�m�0[�Ƙ�,ь������5/-�B��uɛ�`��*�ծ�F��a�����Z���!��͍F�*N�t:�����e�J֬�%x�.j`�5�n,�"QXM2
�%��D�6�f��Ȇ�l��5-뺶+�ǭ��R�y�A��*´ŕ1B�aL
���v��n^��n���s��;<��+מ�.�n�p�3(>ۧ�z˞.��v�cs[6���5�ہ�];]�&L�M����&lf�n�C��KG�����V�`͒�L�z9mQ��pu�)�ւ�gm�3�؃��9u9��Q\
��{g�[M�ݷ�;��`'�k=�'�׭k<v0��|�^*_e�ns.L7�jݎMƌr,�<�����'��HG[+�J��XR"PV<y��#��f����m�ϲ�q�����w���Nx汣�3�)��6N`Г0t4�r4�h�6��,\�����FH�<M,�u+�c�tQe��!ֵ�WFD���vS6�-q�G��u����n����pB�E�-V9�h�+�:���ɺ�G�@ڊ\F]5���W@a(���!�|�e�zj�θݍ�]�ݢb@�|�v�\=�Wp�v����v����gr��L�D�4��Z�-�T�{bn��q�bZ\EwW�����Nw<����<�K��: -]�V�:��=sZ���ٍm ,]���\Z�^�r�[���֌�{�={<u����'�-����J��{Vl�]�%(�=���{uY�ZpO9�ܜ���tm�]Ų,�̩.�D�YUћd%��9@"�Z=�{\�E��d};=��Ԗ�������wK�e����q]�*�\F�e.3f�1���F8ڠ��oi��J�q��l؛�Nm�� �E=�r=�G0cc�G)��WY��ђ(;g�`Ŭ�`}�R��9��y}ob��6�:x�%�f�[3x����'�ֶ[��-�cl�X�.q*#t�#CLF�6����Z��E�(8��H��K����b�5�]�؄.��2up ��űIn�����6�5��Ƹm�ݸ�s`�f�-�Uݝ�6;Y]�6Sͨ�:��Wy�s�u�rW>,2�ɬ��$u�a��vIZ-�@Kh��Im�̉f-�v�j�jC�Yx"n�9�Cdbx[��)F��Z�kqè�l7:x��j�>����.K��JZ��*���;��lA���a��v÷];�+�up�\G>�m��^n�s�,�^Ўsu��n;/B�sKuԊ)MGdI����N"׊xz/чg�8u�r���G��u��<�ʫNk���YE��f#��\+�F�WkF��B�R.�R�]�I�s	�٬��Z�N��O����ŵǰd��7Wg2v�'m���S����a(3�a��Cdbsc�ƺM�p\��x�wd ���l�۬��0���c�s6�׎���cP�>���Nn�g�Q�݆`�qڵ�%��R;JŮ�M6S��Q&2�H��3iaK�*���=�r��j�^��=Y�P狗G3n�p��;j�k('�Y��b�.Ϫ��v�.}u�/;�5�����ˇ�P��=�m�:nc�O;O�ո�ݺ��9�5Jd{D�X]FKSCv&�F3i����:��|-�Ȓvr�8��/.=�V����]A<����X5Ҽ(���gYZ��˒*�f��pg�x��zOM����upK�ib磕�^��#v���V���;e��N[���g�7)���w\M�k�wn�g>�+6�p���uB�є&��Қ&;&�V.u���@�J!�Iwty�:��Eck��yq�Æ�V�v�q���!��W���vY";5�8�¶������KS��n:�u�`�����>�ie�s��J��O:�9:���֮���]Z�O^ۤ۲�XpE����s5<�;<F�\��}n֨�=�v#3�<k�G7�6�-���5Yu7QX�1c��mKj�g�;�sy�^}��w/*�nK0T��<{n��ٖa:�
@LU�� +��@�ܛ�0�J@]��"WD]��[^��c������Fڠ\�j�c��^�S�G��&�<��9���])�g��%�sb�l��)�0�9�o-�7�k��t�&���k�|����v�]v;g&cG�s�Π�d�4���#���t�;]��X���OAj`痗�w!ڴ������H�2sv-��W���ˈ��g�=h����6�mv���ה��-\Kp8���]U3&¸�C����O��<n��f��Z@[�v�c3T��5T%�Q,tXb�j��W�iۏAìќ'ۥM���v�7q�Fx#Ɯ�[<�ޏ1�-��0l�I�ۭb�[d�5�lŊ�u�Ű�b���[���-�v�l�s�]t� (ݎ���vG��e���s�0�Dl�#݃q4��f��F��h�9e��2k�b�dOKբB�a�S�n��t'q�:.Ҵ���tC��mۚ��qC�,�5X�h��e�q�"+.�㫧\�i�����A� �&G�\]t�y�.ۺ�1��E�:�<�wbk�v�����ρ�L>ĕ·Y9,����=����D#�Ŧ�sr�t,�����G��ue��Z9k�nE1<��A]nsg.��I�s�L���Ƕ,UN(�+b��C-���JG��m��������QY�Q�E����Q�3t^{vv,����{le�:�{]��[�ۣ\���·��nœD��B�g:m,�<R0���:���.�n��D[js����չ��Wnjp�����N�펑
n�LV;�����;�����v�֋<�ņ��$�ƶQMx�4���iX)2З�Iff4r�W5�!v3F��l����2�k��������s(NŅ����ֻ��*�M	��l�/
�L��Ų6Va���7�;q���ʻ�nm������ ��v:x��{m�t-�qN �OY��p�mh\U\h����}��r�V=<�6�Hr�\�J��]��/5�����FQ�YBa��Utѭ&iL��l9)���W��Fjnvq�y�kV��SH"���A�hzыjxi�Κ:�%�|��Z�C[GM��a��ғɞr*hsq��lM�l�.����GMtb[V/�k-�H7�gۘy-f՚��gY��:ݙ�M�����gF�p��L$=���K'�r݂�Pn��j��u��t�3���*[.Kpƺ��<-�����m���ֶ`�v��Pf� ��
9p��ϖ�C���K�Bq*h�^�ƹ��x]v�i�vt�1�:*��^0=i�ژ�gcntkG5%��o^�&�2W��%�֋�)�05��U��۳���]�G3�e���-m�[���q�(r��\d;0�"RP��5�sL)�t�mØ�G��J�V�:�ۥ���f�,�î7]��]�u�w*�����VC���q��sݳ�������gUg6Mn�xz.��jrl�a�M���;1�\��n�l�k��v��h)]ln�����X����U�з]��]3íp�<��밗l�$V^:뎳�O\�ӛ���
��Q��9A���\9�b凮-�J9v=�,�Lםڮ^���0�@�M2kK�·l��Y�.��W�H�VѪp����u[Y9�w���hǬ ��ڄCq�����˝o�" �d"gn��
����vG�i�Ry1O�Ixb��j�*P���Ϗ� ��ƻY�h��ƶf��J��Y�s,��m��U��lz���s�|-����Ѹ.C7T<v�-�O|��A�
�o<��;�Olu�]�Yj2%fՋ��{5�	��3� e�p1�>8�4�ô\-�%�A���2ěM�l�Ly�!n:�@�n��v��:Y�@�4�i Xh:�X<3u�P��Z�5��qj����+���V\hX�"$���QMI���D����Y�������������U\���4GWd[H����!w�I�3��9PQG'���RDh���3����x�|u������:&j*&����i��q���F"�B�cU�R����?3�3���x�Ƿ����:)�l����$�X����-l^�� �%�<,�`�-�$�H�"�	�e�z���")�0���E9�D�t,㊪3��ֳ�q�k�u��I��H��
4I܍P�#�I�@��t�	؜��Yu�lh9%�*���D�
(��cH��*%DD�%T@�`��IMZ@UF�Ʃb�A@bB��`'|��� )$B,>^�x�T�hi��%���.�UY�Ȑ$'҆�jLI���B�g! ����kxQ@�׫dR����[e蜄yH)я3�N@�AQ�V�@F�y�1�R�2� �>�.=+M���JjM�EP�DeM�"!%�-����E�"��r�@��!�X��h&�sd�chmUhSi��X6�X�Z�P��Iihi3, @�s q4�#�m]0-�[B�m�;a�@w��Gܓ�����OM���eڹ36�s&l�g�vy{������Gĵ��r���k�ȏY3˫���fGf�b{���.Zݭ��lCe��u�xVʺb#�����	]���17��֋wFv�{v�½��ͫ�������.Ycq���WU�!�n�ձ,1���k�S
v/c8:8�.�2/\ٴCxx��홄�q\����rt68��֮�.�m��ۋ�9��jl�Xi`콕�7f/�f���w�1��59u$�V8����Aƃ,i��Kn�4��fb��ڜ̄�ө�e!�׉Z�0c�D�]���U��ʼ��.��5s�n��*����9��[�����>2b����jw+sh�v��lvc����4����ڞ��2��!��� E�\�zݪʧ^�11ٚ5�h�]$/]����w[s���^��v��F��:�z����{��k �)^�!3rM(̺u��w!�yݮ�w2؁L���v�n�#ْ܄&����F�mw\+���J�v2���YЧ�lϷ<,���J�gA��Q�g[L��8�h���jN�PwH������� ��k�Ю����=r�\���m��q��8M�E:���Qn�cD��l0���ѻP�#l" ƍ�Z����Ŗ���u���[G9��xCN9��^�g�zٔ-ֶ��	���Z�
�1k���&i̶�,Ͱu��F�F7]40iE�e�5�C�!�w6��-+�g�n׍8ꑆ[��sn��b@�$
)-�aqc\`�����hۛI�Żhug8�p�A���'kY��Y�v�J
)C�ĸ�[s�v�^��Ei��Xą,u���c6�[��jd-Ce��i�����J
.��ԳMz⣠ݔ�6c��M�ɂ�\��E�$��d��$T�Dk�7f��]`I[�^:�=�| 7��պ�h
��]:I�h���X���m�+K)zRаJZ��͵��e�*B�-+JBV�/),�/6���Ie�U�ZQ�m�Ō����ԨU�[Ye����XIe`�%��d�6T�c�6"�:�j+
R�!V�U�P�a����z� �,[a�m���KE*&^W��c���QQN�{��ĕ+XR�m�jZ������8g$2�iI �EDM���rS<MN��߈{�a��E\TAo&�(0e�&��Q�N���_�o�ǃ��ך���Hu��x�X��	7���b�m��&�&�L��3���l� ������R�e��>��P�H$�E�?�$�Ƽxv�	����.Y�3�}q� VB�&���D����I$�kk�-�H����M��S��bצ�D2N�tc�+|� ���`�K�k[ 9;�q�|-R{x�����g�&��}b��k-�^�k�tF�K�u��<�l��ʒ�M2��s��%�v�㑽Qν�kU�\�6�g�^7��k�N��#D�
�@��S�wXk�g��żR�w��02�r�#}r�]2�ji�[΃D�zTIw�^W[�ޝ���_�C�Cw�+�ؑ��닗�4'mڲ�,��L�3h��~ӏą����|�I'*������p䃰����e���\A[��!#d�.����'sz�-;�lʒ
 D�f��u���}z�A� א5�9!�[k:d���/[&�jъD�O�g��o ���9'[n&t�f�y�0Pw��w�x�r�1q�&�\#"��^:�QAck�@�鮚�}Mn0�$׸f6��'"�d�/����s��)I����y��j�� z�&sm����<_j��2Fb�c��S�v��'�6�|u��mvjl֬9X�I�^8E�)�d�`豁T_k A#&b��7����/�#.9 ��O~3^X�Y�D��,�W}�x�70���g=��T�� 2�v�}�iW��z�^q�C�͡���YW�3��wϏ���8��{t�=�ꟇN�/���y���jc
�3BLxf��Ã�L������y���#3\*w"��e�Rd�:d좨��1v̴��17C>�rA ��.#Ē[cYE�Z�e�m��H̷�9 ���t��:;���ȁ��(�l�Mm3ȍ/K���u-�$���<�	c�A�|��U�iO��,�(L��W\i]f��70�\D�ͭN^)q�6��Ny�>lQ��n�����[f.7��s0�@� ��W��X��5��Ɛѓo�//�0 _O��O=��$wdD��.��c�-��-��
[�`p��/t��Sx(�Kf͓���$XfA�59��F�!ρ$�D��b���ǻ�	[��#F���ȟ'E�A�V0��yS.Q$��D�{h ��[�O�7���z!����Ư�����Z�[|����8�<D�t�)tC��[�[wLJ����d���#�(U�C$k����=}��~�%K(�bΖ�e��v�?�2�cjս�F�TCJ��	ͷ�Y[�q��mDg��a�����u���/::�F+��r��sD��8��q	�N$���E����?l����?�^2w]����� ��8�/5`1u�-\�x�fXcxM����*2�tO}��Yz�Iҷ�N�pH6ũzC6���ֵ��	ʾL�A�S���րH;X�9�,�Ll�xɣq� �|���	�3K�b]���r��H�[/1u	"�\9>+���C��݆-
��g��	4�A*�&�����b���W������s�J铧��F���0m��$KN�E�Hm7���]y1N(ݩ���Wnl��S��W:'� ��A�[��-��Q۾ܵx��Y[��|������<��sl�4��m�gwR�W�:VՌ�K���m,�&�`�@U�(ݩnL�krь��=]p���4m���9����]b4�?7�<���4v��s�4	�FP	�W:\��r�#�h�;Z6����r�V�#��BAL��(���G�LPt�;6�&�Ic�3iwG3�^�6x��׫�
��Ӷ*����U�Ѱ����i��;t�#��"q�5ڣ*�8e`�>wl���Ɋ��_����M$��$�m��/op�j��
^GԮe��������}��)��<�/�'��э��M;/�{z��s-T�^u�$2����q ǓL5�9�(M��u/m�<���&�3G��^Y�S]�A��$a����lQ[p��	$M�$Vm�O����PcEӔt`*�>����Uߚ�W����<�5�iC���������������p�~�-��$�`�EP,�� �N�{��F�M�c0�9z�pB�؅�Ï��m-�>>}��k�ո����-ѣ]zjʵN��'X8�tC�.p��.�瞝����]���k��h|V�7��"�F�x��T�c��ȸkp�O��Ȃ.��"�3���$�k�A��O:�L3^�-�.%�V��uu�Mz�[ඨ|��_ +1nn��,Fg���C�d��ǜ�����L���r���o��|��Z�L���a�Iׇ�"<��]��y"D��a�%&}�!n���[�zٛ�ʹS�2s`�z�iPerv�����L�s��.�\Zef��b�ւw2����w*g���cE�������B����M�O�u���j���4�K	i����I|Ш3�d$Ȣ��̮��2�r���u��5S�@$��{"������
Y��� {F��9P3N����ˋ��3�9��ת7�;�>xL�H4�����$C'DG����3�����p�m	�eS�³]ψ�q�d�t'�这�fլ(��ˍ��}�x$9Z�Ω��C�����lz�יVE3�uU�E� >y�J�8o$�����cE�z�꬇4`�;�]Y�����as=stZZ��z2������޳�Guq������pև��sݮ��"/��_�8���}��}����y��U�{�(n�ܼ��#w�Rr�W�|��z��A&L�ÒA��g� �v�m����u�������p����r�@���8I���L̊Ѱ@h�^�^1��q����F���E�_�ϰ	��� ��FR�1���:�K�!�.��<���tܙ�K���]� ���?ԟ��1r�l��f���O��_6 �����3����D�Ⴕ�<�7�I�S[����'�X��5��	$^[���_�-� �`0>6���y�ūT��ƚF�U6�R-А��&�o�c0����p ���Zvy{���g�{ȃ9m�Kv��mlPD��S����Pk�k��MJ���}��H<��᭷ac�c�M)5L�����!�*�� }7�����{��%g[�z띳����;�{˽���u�?~6�8�����zr�U����o1���T����vQE� <��F��eU�^5KH�>I6s^�y�����y9��&"��Y����0�\�"�k��(�le��۪
��۩���y��0��a�4y�j�k���3T�����V;ͧt�!ןT�$�m�;��3Bk�����D���{�׮]A�H[N�G�����tj�Ħ�ۻ�G� N�D�H�Z��z=����7�y(��3n�� ߐ���4���;4�ݞ8�*]]��\��ȍ|BD�$w|H'i���s[An�+"���굞������a�/F�:�%@$�.�;�fm��%4�z�ϨA�XC,o3�u;sc2M��E�!=�D��y	���Q	8�,;����{�������eO>�oM�c:cO�d���&[�yi�dH$al�޴���켷q��[h�l�t�����RS5���.������n:��5��H-	j^ۛh����@90P�m�;,��3�����IiIX��!ff�g;�-���=�8�V�8.l�E�ۮ�J�6���c�Y.�S�����Yq1�jL�M�h9�י�R[dGZ�U����h�C4�j��	���a����曀������uCnp'b�OgC�9� �S���糲X(@�@�Xjو0��������� 	J�<�H�l/�>}�5�q����e�1��@$*j�'Ł.��Kx1�2�	��f�/�mx�����i�5�x��N�.@>*.��:��w-���Q�
)ؘZ|��kS��$&.j����4r�Z��w/�K��pd�)�8F���YǶ�[nK�Q,AK��@�F3��126)�^r����w<-�ȗW��]�[�&^u����ۊ��E�m! �M�`ʿ~�B�ٺ�������\�^e�P̻h�f��h��F�Ζ�{seշkP/�^���C,W2�o���jn��Y��Bn��h�
ke��t�5kh�`��u@'�����_ _z�ci�G@��_������پ��1�Ί���z��4|���w\L�ۄ\[�[u�[��^�W~L��6a��*�R���a���K��dk�oə)p(�����Ү������ �YH>a������P	��i�Rw9h뽪p�$-5hH��\�HN��3���Z	.�9>Kn���
d�d���JmQ�'������&*�=$�Hx�)���XӪ^����ٗ+p��UG��Ca�A:A����^��#��!��
-�Im�ʚ��֝P!}N]�����a�D/� ���K�µ�����k�����s���R���E����&%��&���8$�����i��
m���"��U������	ܐ\�u8u�� �azc��� �mT�H�$7Y���C����������ո�����fU�y�F�H<��C+U(����<>�m�;����t�;�S ���:n\�}�6��d]��B�k�Y�Լ&������!˃����(�a*����w���w�a+<����{�b�z�z��}�M���<���W5�� �' ��\=W����tI>,QKE��M-�JGN���P��/f1gy0p��7�<[e�;��ҏ��7��v���]���q����Z�f�8�Ҏ��;�H��9\>?n�=�1�gYâZ���yC��x�X�����=N<��ae��W��yur�GO��Y�y&/���ph�����j��]fn_�HA�=�F�q���c��j�����;&�n��C��ﺴ>�h���t�.�x���Q����\uŃvm׭k���|�{Н�1$Y{ ��l
�uē�Ǌ\�iFG�+���*n$�g��A���yĢX�Z�����x����>ߖw��̗�}k�w	.9fk��I�������ұ@@nw���n.���w%�ɾ �-.��r���>��شw.��2'e�\��	����XN��۾������w��z7�w��w���93�u\�﷼W������۽{���r��Z��^�X�S���^Lp��}���{ܴ��&�[�4Y�>{�.����x�v����,�gv���e�[��Ş��z�y����`;��8S{��gdt%�܋���c<=���g{���G���H����|l!�����]X*Dz��1�� T,��`�ѽK�*��(���q}�w)��x�D��<�V��I�PJ�+ҽ~:�q����x��~=��===W�wZ4r�iF�ּ�u�Eܞ3p"-sR��Ui[KjҚ�)7'�Z��?����<~3�O�^�~=���YYF#�hH(�lK4�5$zx#^��=2Yג�h�4�P�Ao�����x�gۺ�yWZ��ku��eeee*)$��2
G-�!�.��t��2G.K�]���i���(b�Q˻Tw���dnTz�T��e�t���-�%Š�J
0�N�J>2D�
���9��19P�����2���� !��-z t�R��V���$���^��l`[jH	�,&2㪧p/��S��}z��	�/J3ǥ���P�C�qUg�&Ա&
�4�����C�֩)H�:��P���fJė+���C���|��"��9��%F��KR��+!*�(hZ�N��a)���S���U�"�p$x	@��O<s|݊�c+ JX��xD
Jg9Y��^ߏ��fYG3=�Q�ƍ�E��i
�����(�n}Lj��>���PZm
�+��&Im�rC��DP>}�����4��{�}��A�����
4�ƪ4JJ����*��*4D��_�>O'�>~o\���@i�SVաQ"k7���Q#f3��Hc��'fQT
�#� (�O5����Z�d���#��3�v_<���{���dr��y��;�z =6UBէ�f��V�JSB�J���E;$��>��<��5����������\k��tN��mb����upO;09{N���$o#9��ߜ!2L[zW�_SG#}���=�x�73�R|�<��S�T-%���Q=���Yo����lm<�Υ�='��T�	��JQMW�g�h�M�A}_yZ�xD����\������dkBj���~�Yg��|�����}K�K�8C�8y�^}z���C��/Ϯ���&�rO�p�>�/�61�` !���D��;/�s8��|J9ږ�2��Q��R�(���#T-P�B�n��w�z�f;}wo/Ҋ޹�q6���WH7M��u��U���!������X�i*4o�wG���$�xLѲ�A�"oϹ��>��uپ�{��rLc �=w��bV5B�A"Q~�ZR�J ƼH5w8�= z7eLF����5\Q{5���Irz�8߻��+�,����3�x����h��dƿY�����Mx����w�o+֘]���`��fR ��~J#;��*�hTIG~���Le˗��|��x�����P�2�3�t���>o�7瞭����9�=��QM5�=�&���+�ָs���ќ��y�d�`��\j�n�<��-5�&7=�gU���6K[�b�O�ߣ���/.��U���5���Q�ƨ�)��`���:����h�^}}v��B|�o�b�P�sh����m�`y���&�񨅥y�oM�*�/6��x�	�vKvW�4D߻�(��T�m�n�}�� m5�f<^�����\�q�>s�"4H�S�;�J5LJ ƨ��s�N�)J���9��>g��^f�מ���h"B��i�0p���Ģ���TR�Br:��z�=K�JN�˴��}vy��=�9���*Ҷ��j��|���hB%T��A"g;����D<�w��qs&��r���_w�9_w�ζ����6ITI
/��j��Q4!����6ѿe�bjR}�ϴU��[�nw����r��CCU�_o���P�F�1G�}�V���K�&p�+ƈ����h�U�TB y���*�76���ݣ�g�|wS��P�����{�n�*��6޺<>�"�O5ˬ4�)D-Ӗ��`T!;O)s0�i�|���U����~;y��z�q�f'� >�o�����E�v�Ȟ�0#�E�j��d,Ģo�x�q��w�dѬlO��xf���	v�mpA������v�s&q�����#0��j�����[q����v�Ҹ����a�N�ݮg��]v�n	�4q����۷g�(��+���k*�xn�w`�,���:�k��Q��$ځ���ؓ����+ɹ_sA#�wm�HDL�K���:�	v��c:rWv�y��;�f�^=]||.\��y�wk�3�n�\k͉�T�B&-�Gl�F�5֗ �-l�K�e�m������-.�K�q�|'O�κ������-o��>��%䠟���(y��x�}�Q�)���g��m���b�j�"��A)"g>� ؛Zh'J�;�r��[̻� �xYG�����As�}ᵊ.�Fpɫ��@R�k���Q�Q �D��w���G�C�����^���A��@]���`�߼'�#��o������]�+���o�(�T-V�#�C�g��lk4F�	��c%���Q�׼�F��A�Q$<ןe��(�6%���tU�頉��+�S	p�Pz�������)�v�]�������Q�l����^Fw��p��'�ϝn���'%(NOϝ}uɯ�×��g
� �j�5�9�lM�=���R��Sɾ4W)���uF�k�%�Cx�:�x#�Us��˛�_��q���w�Bw$9)O����5Ahn���
+���4��������9���W�CLS4�hK�
=�8[�:�rD8���!��//��r�*������
�l��4?D��~��t�r��'��^�tL�h"F�$J'{�j4V��s�M�z�3�8Px������B�J#)�����6�D�}�޷=V˼��͈W��T^�y�kH�y}���[l�\*�U\�!U/Q���ƔD�C8�-I���l6�&��|�U��O9����iQg�H7w���Qܻ�+=y�u�p���Ji���i�
���o�����N<�����rR��=0/	�󯮹/d����|띝���s��	����i�,๓.�������7N5D����.s��F�]4=��>�ܼ��O��&���Bl�>0�G��ם�K藑�%�U��>uZ��>��{�.��,�����Oz�O�np�� А�)��Qr'�y�G �{(�SوIy$�s�;c��X��b\ ����{�fzN�'�7��$�p '� $�/��&lA�o��O���/�-) ���l���	$�w�H��'V��x�R�/��|�՗��[�,�sf�E�JcF���M���ļl]1z�kYH���}��qT��f�d� O�w�^K���$�a�zD�4Zb�\�n��$��aΖ`:�cfI�	3��)PK.&��䏣͝{��{ ���K��	 ��}0%y<�H�E ����(sWt0����Kg�)�M��\ $�3CWCx�@3i�`r�=�}7b�h��7��L�]�s��c|X�U��ר�t�eB�!�%<L�׹�(����c/M5%�=�I�w�����||O����i��@5Z����&U��	��ε5�g~�7��|&�L�<�� ��LΚ�	������fG|�K��Ǡ�@$��t��>Ewsd �q�Nq���V$�c�!��wF"���!�����mt�,̀Ux���n%��Vl�b�lf��y%��y"��s̭��s����B�6Ȱs��C/3 �Ȼo]A���.��<#�i�)b\-� ���7�G���	��q�@���9s���H2�I+���T�S���Y�/�=�~0!�O��$�JXz�	�d�eUAsƼ�	��k���{i�����+�_��3$Qy�$�@$3z�L��T/u�ƵL�9����Y�p�L�'�VWLI�`�M�c�2$���u;��1��FRAC�șE$�z�L���F�ɓ?�f�x�&�bҵl�KW�(�3�o�A-,�wuē��) �yo3���X���M�r�`�:�5d�!!����t����e�y{�Zgyپ��nM`ye�E�4����k)�T����7�~z���έ�e�o>��f�X�pd���2�
I�""�		�i��AH$�U��#<���UF���kI4�ș	$��_\ɔ����8�V�<q�։��S�4;%�gN;'vAY�2����s��ҥ���k��Ք�ٵU��>�O䲷,`�pJz6ҥyO��-����@$�]���}�m=�(z��͛�>��37�u�I&}�y�s<Hp���I��� @	y'�D��^g���($�P9�$�d-��	e�Ӎ��>�@�*:������N�U���I3�1Ø$n�2����8���efc�|ǒ�	 O��CYZn�<���nلYx3E+�W�Q��z{���	 ���LDǙ�d��@�	 �M��8��K�Q:�e��
}����,�3?�f�4CɁ	$|�iΉ�ً�aԆ��I.�y�!#�%3-���H�o@�J7Vm�{T�aYu���B:#�b�cT�x
'YҔɍ��	���s&[=����z`3 ��{$�H(�{� �?hd�x���4bH�-��Г����O�i�fR�+
͑�l&F�=�j������U�Dw�Ļ�������ol��=n]���ۮ�:�a�J���M9�p�����Y��n�OD!�=b��3K5�itͭ�Fl�$�;p#��)�����za���oR��bh�=К6�Ѹ�헦px�u���̈́Չ�s�f�E��<�Z����	��+vH�x��+��E��,�6g����֛aCk��K�(!t��e���tc�K���?���ˑb�;���q�d2IX�c��fH�_��D���(dm�]�ۍ0� ��]�·.`lv(&��U^@)|�e$�Z�W��!�F�=�/S���($�I�@&��I.�o[�lv޷��Q���S-n���^w]vjI �vdIs�2B�ͪ�[���@$��Iy7gH���;���GP.\�|�7.�+�ZT?Ĝ�*��%��/	�I$�o�D��@-�n�<;N��ӝA{��:5<�}�.لx3���6b,�{|C0Ȧ��7w;D��\O&��$��b�2,���O� PJ��O�w	�8L]�]H��R�+�"�"Vf�Z�]u���͆��.u��Wf,�(�ū���7�$���%?H9�l=%$շ	��l�@	�!�r���UV��i���H]d�;�ڌQa!�"�Ӿ����R �zgM�#��;>�(ˮ�������OP�^�J��=.'��3kD����j�A��Iz9�f�T�L�R���U�.e3����q�� '���e Ƴބ�I ��z,̄�>E�~�! �@_b��B;��e���$&	�1ft�������R|�K�VKdHd�%b������k��D�eF�IgKt)���'��o(i	���ޮ�t>@��~1!%�d�ʔ�@$������6��gR8�8�P]�%��3���ѭ3,�Iv6Pm��w�OnJJ���	 �H_4��"io<F�&��i�W����a�`�V���b��9Zۜ���!�;��vbZ�x`���W�Wٜ�1g�
�NSLpiA"�S�.�@ �ݵ�e "�d�l��
F�7TM��W�Wm=,@3�o�y�I'��w|y:d&��O�;���8-�sP�Io)�bk��uv��%�Z�v�famӦ�Ud���F!0��"�z���}I�ڠI$�?z��n���;��vرt�/�f�Y�>�����£!�pV\�k�5uH��E����,N�P(g|���o)y>�dx&����A%j3���I-n��A7b�3&gH8c���h�~�v���s�;�G=VѳA�G��!͘�I$��=����O�=��2��W�ֆ��͜�Ф$�g�R|�9"�:���'�ʖ��H���zI ���8�ϛcF��a�������x��|�m�FW�uFܯ6�:�q��v��%s���5H��jݭ/�=��IE�r�D�}�;���@{˛u9���X�@��S�����B���� ��T�3�cW$�Y�	3�O�zJk��I�*�i�����md�G'ؐ��3$��TB@/,fl�� H�W��կ��5*~��B31�b��Ş���i�	��f 67�s��I)�P�Jg��� iI$���W��dL�dH@�~�hY�3"C�������ݤ��$f����,nu"	$��ƙ�*�0�}��7�,���;ԡ���<7���P��|�鳦�|����@x{Zz�$_����O;V����nm��V��>�5�>
A)�`F�ܒv��hԝ��u��1t*�-��($�_̉>�����y�A$�|�3 ��d�7�L��+�\�|c�ѓ,.�$����+�>_6�u��vWH����6<=E�^<oSW*���F�t7?����_;��:ШˊO��I,U�/!#�S��\�\���DJ_�D����	�r�Uh\zf\�@4�p�!1�Uka/"��H[�H�d%����=��v�˚n-��Lh�t��m��dY�	3�RԀQ}0"BI+5��D��F��OX��HgyXN��>��A6�z��}��������?��߅�V�*�:̆�8L�����2�&RV�v^RI5v����F���L͹{"})x.�)�ݑ!�|�PcvdBI$��ڢK��ڢ˂�o�^y�����@$)Vd��$=ͦ!7������a�iNn<�f­N�7C��ߞ��w�q�]�]����q�fާ�4����ي����yx��pK*g�Ƿ{8�1�x�z�pO*��{���2�ĩ)8Ҟ{=����n_j�׵�b!j���_e0���Y��Ƿ=�����-/��}i���L��w��{SX��� �ڻ</,�>�`�r�'i�_{.tB��'f���w�Ps\�p�Qԟ�d�Ō8{G-�����؎7����6�y�������w�:��{�"�{��$�.�\u�ƫ�.e{����v����س���_
����[yv�o�C���M��Y���[�s~��n���L&�L��O;�w�;8�=���%�g<ˣ:�j�8�X�?h� {���n̝؃Π�Z��G1�ڷ}�y�������v�p���?z=����6�M��N��댘����]����=ׅ}->ȵ�����z������q��E�;Gf����݀O4o��-H�8ͬ�{7W
 �α�O�9C��d��0�7����������3o��R�ܩ�+�Ã����}�鞼߸���g��'.�FB�ΰE>����ǰ��77���$]ʲ��s��)�u5ۼ��Nq�:.��{�%)��Sl���1���{��]�2����cm�oj������7�l�Eƾq������s��]`��;+���)�OǻO^3$��~ލ#;����Zs�X^2���8�()�L0"b���ˣto�@l�������-�����t�B�H��_�[�G��
�=ר�'��5G����B�{�W��~�TCq�l*�����|7���-DV0�D��Ïԃʉ��O��i�S��l�5�&d��UX�	X�s�A<�x8�Nm�R��,Z�d��m#@�һ]�jSR�Mi��u�_��������uz���Y��K^�9:c���+ُu�*Eq�E�$�b^Ἡ����oA���~>?<x�gӮ�����}>�Ooo]uÎ�:��Wm[�,ADj$dRQ�f���#H|z'�pws��"����||x����O������n�[�֪�p�me�I�� �5k�Ș�������6{;_Ƅ��6�Ѭ���'X$o��Lrp�� Xꛗj�u��K$0KbD��-Մ��R�gsW[�LKLbK閡k1bO�a�����6���Ҥ"�[m���=�d8�l^�|z[ͭ�N�v�H��D	�,$�	%j���KR��:$8�����ù��S4	�%"i��I 2�@Z�P�K*������yVC�<pxU��^U+#'�{�<&�	6�)o9�5����SN��^�ܔ)��Jr��͔�V��8��V% t	�	��Y�k@������|�H�3X�+���bsD=7�r�U �nTkr(�ND�׊�	�|P
�6��F��A ��)�a��|���F��Cz��&�g/p�Q��S���67M��״=��֧�/I�͎M�Zl����������ٸT�J�=r ���vs皨��M�f��3��D��t�k�\�W�t㍗���-�U��u�䬻6�2�=��V��huv�<��v<֎^��R��;���z����x��-�E�
@��Զa�tƗ����f�5E>��#�9���wR��Z�r����n:�7g�����en.�=�	�V���8k15��]�Ӗ��ݞ��v�Ut�v�dC�4"#
�3;�k�u�V��8����5�e� �
1�ZdMwT$��(&<{7�ܛ
�su[��e�j7�F�m�q�:g�8�A��4��؀��vH�v�O���r7\�{c��9ܦ��ɢ�3R[f�@M�u��#���js\7'K=���j���t�%71&���"���k���س�>�"ws��幗���v����lnr��]-cr܌J�6,����ؖiQX�Wgc/��V|80�;]6��	�W�'&�i��:�;�c:�k\kkQ��r�<<]��ă�#�QR]���لm	�)��6L�m/`�u�޹�/�G/-=�ݵF7W�&WGO1��/:�P�f��l�W���\�r6��ݞ��9kz9]�gȻ��v�6���+x�n�5�=��-,I.v�g����܍�U֔��-\U^�����5c�GiiyݠW{�8�u�q[w)ۂו=��#t�l֭�Cݱ9v&{k��r�.��؝��3<��j�mxi:ʏ��t���RJ���A�@q[��Uc�'M�^�c��؜P��b;'A�k�	�������Hjk �I�u�!b�dcE ;a���Xi�B%�fJvKI]jKj=o��p��I�BHt=y閊�ծ��%�rZ�ّ���4�ks��X���F9��e�#	���rN�ۏ[�#-�9��G-���i�yσ��q'~�����^�v���^6��K��X2�2҃ZV��kF�KP��S*����eS�oL=��Ōbr�űm�٥�yn�c��gy�ݲ���Y��ş0g�q᮱;s�hp����us�,j�p9��lsE7���n����7I��[PmvCp:�]�v�4Gcy�aI!}����e�v�0�?(>^���t�~dx��9|�+�ϧ�3~v�B���N�ìĵ�dO� g�0����@uz�
c�pC�KO�s�_��o`��ʹڸ�>@�Vt���fb��cЈ�ꀺ�6v�ڟ�g�&��h�!݌�-v���K�|��7 �@/%��U���4m�H���&��z�����v��ȳ�;�h��T��4@���3�K�̒�]�.�Ho/�$$JM���m���lh�{'�R�符�$�,�!3��{�n��шI �U�1>3q7��wt�"�@i	$��}1��	vtȟJ�x��/g����?|��q
��n�aF�����j�=�7h��6{=9�l��������}aKm��훊u9$�&�\@�I.Ι�
�Ǫ9��kH������%�� ��K�U�/�JځA�"�:03�x��d ��G��ȯ4�~/� �����{nG��ܒq{t=�0�J����)�(�i/o�+2y�Lz��9����|��<� hD�>�s�]��k�oH��C��I%?lȟJ(>��,���wkJH���b�rB�������Iu\ǄHH�G+'ǈO����O� m�%�=�0.Tfp�!݌
��MNV'�+��N����x��F��uS�K����	��CvK6 ����skRAe���Ё�K8A;�37��%��)/���I�� ^���}��fyg��\TxA�)d�T�2&W��H�.�bz1��s6��A �����$b���D�vr�2[!��I͔��ɳ���sX3R۹�?|��cm����>� ����&�7�t.�b�xV�
_;T�]�'��
�fD$Vtn$,����$��
)uL��(��F��{[nM��ّ2���d������@'�Pؚ{�Ù۝YnJ�AсwiGvD�0fA*uy��($��y<�[	�KUt*�1ؖ���؆�d�/']�K������'���e�X�|�����'!ŕ4m�)���A��{��x|����!)��<���$xtۈ��	 ��dH�7�a�S��Ғ���%�bܠ��OKb ^'j��4�@�H�x��$�$�ai�e���K� {����]-��\�5C����ۦ�iqk{ξo{�jHI�ٙ#���kn�ԁ>`�{�"I&uOd���K{ D#�6V�!�6�6��D-Ms��V��m�GZ�>���acuu�Q�آ.�-�/������m��?�o[.
K�?�5�w�}�PH�q~����/`�K.]�¾�>�W�^�[��Kl�!��p勽
-���}b6k��Rב�Q&II,jޗ��y�6�3s>�PJ��嶍ޞ���
��H/32����9���32Iv4�H��qm;󽋠�@ ��wK�I �[φ%�WNK�E�w&���ܬ�\�D�~	 �Rj�&'���f�K���	&�L�6Ŷ3i|�A��s��|����{����ݧِ�ջE1E��M��4'��[������,k�T�L�V<�8yJ�a������ >�A��(\ �$��R��	+Q�/!%��_�d�C3�T�Y�7	 ��$�>�ܲ�7)��z����k�L��	 ��B$�ޘ�Rۀ�.a���a��f���,���!3Vb�GG]��%�R1�!�]3�7RmmO����&&�����3"Ho��I$�3�2��\�)��*�t��� H�/��b-e��d�%Up�?�_��,I{�����]1P�^	 �Ϧ!%��	_tȂd$�/������Z�����X�ԂhQ�E�Iod���$��4Z�W�� �N>y(`̗k�B�%$���	�I�+'��%��v�7bl�*|� !�LHg���/n�O��)q��z,K�4��a����{.g��:�u�.�8�.�#옷�$�$�卑"���Sk�F�I^>����Ń [�R�X�\�z^R٫#{B����Qy����rU)z����*z
7���W��ߡ�ծ������-I�I���M�&x�`��=?�L�T6L�V�i�ؔ��p���x{�x�dN��Y���>�{ƪ̑�E�=���qڲ����̈́ ��CM)b�
��r+�I�>�ˇR�fmE!*�IEV�&L�"18�rbַ��Ix�V��Wh�|!ϪwG��Lv����@��c��T�+��7Z��Ӷ�<Wt]���7U5ɐ�v_]��)��s�����YZ�e)Y�v�`�kn�̬xs�S�k�����r�볂�S���ۊ�qe�*66����2�-�F��Ƨmkny]k������?���)-�7�V�e�0A)˘�_�7��f	!�o���N��W��� h	���"�H�v���;��('E�wcUAqər�i�Ժ�3���SE�s9��RH��-�f�G؟zBH$�ԓ[l��磂��ze#�S 6�*f���g��zd�����(��H��׾�"$I�V$�I]�H�D���gއ&|c	'���� �K�.�,��C���X�I%$$@*���ϓ�2K[�?�����bh��]fH�O���"C3%d��d��
mL��~wb@������YK(�өެ��fs`A$>����I]��+�2+�GTuՂ�c���Ӹ3�rG-�K.&*��)ܑ���홶N��>P���xX���~��ј�!È�~?%�s�'��`�#�O�"<���-n��Dw!�,���Os2&QAc6(Χ�$��P�b�g �S�9;�������iT�|z�L�>��5�=xV��3{|�=��?Bzg�)���>�%���=��n·���S�rƠ�%9��Wh�4h �s,��@�FG� y�ДR-,�o����O*��־�>I���NL ���(xq/sU2J��%!>kڶCK�:�c�k��̟A@$M��	$���N�r��]ҕV�$������>E]�$*���%;�Y��h�ݕې�f�g���_��eFz�DS{Ȱ@.[��$� �F�x��+܂2C�b��y�2C����a���&:��|��$�ퟥe���gwsɵ�t��7r�D����Ј�~��i��c��2�%�)�$'�^�k=n1���X�\v�f�l�
�A;g޿|�"�2�|�$��8(5�.d)f�^�@	$�Hk�H�@/iǁ0�ej��r{��@8��f�ۄ�0NK��K�v$'ޟ)�z��#.��s/Q�BJ��#o����� ]�!y"k��;��8��hf�n��<�38AM %����>^*_.%���p���Y��b���������i�=�ϧ`A>9��D4��zD���^�$���a~��<�c��_wWB�K[������xz@!��a�d�*P�(G��	_t6$��	W|�1��>�D�R�S0��:.C;(`1��;�oY/��k�-0�I$��d�L��C��4tR����e{���h��gv)��_La�IY�xu��r�?-�U�r����Q	O�3 �ng�DǙ2Kt4_������O��Q�H�ϰNn��=�^h�HXD��s�r8����|�2�b���ͅ��Y5� �	 �\w��$Ż�は<�Z��R�z1���5�mxA���^�I�kQhv��� d�]Vne��� ����
|ʅ�D^�����K�݌I��"�r[���v�_R�`�0fr��ݓS�@������y�y���2p=�78��yy�%�u}"D��	{�d10;�=�J��8A���N�:�f9��*���'o�$�H��Π$}>`�O��8�yh�%�L��qΤE;&�əB�`LX6twV6�<VY8= �=������Y�?/-(]��i�����?�'p���y��s�o7����*���� �JA*Ј�����>f?^Y�}"D�&r�ن	�r�L��/�S�Y@ex�'ͦvY��m(�.�>�G���K|��Ϯ�*�3$k��O�kV���S��p���bں֛b��]�uxu����knĸ������>�|Oߡ\�'w%<�'�ؓ)$�Z���	!\�`��ڞ�Я�*��&� ��ss�	/g���!�w%�f|�s�}0!t=��_���5zY�3O���x�
%+����
$�w2yŸ�ܸ��2���hH��5�(�H���D$���[ͅ�$����_�6b�����	������PH Y��!!��x�8`��K����.�
]z���w����,u�� ��}0I0�mt����y�%�=�{�� ���g�fp�
X���6	y)���Vu)y�^�?���mp���35�$	 �mt�V����%�8���!s��w��dU�4�f�ݫV6۞���1{�w���NR�Y�X����'癠0,R0�}����2�C���	�d$�Ac��׮�GY��am/<�uXI�n�*=����v�Fg��Q���ܮ�G��_���k�rO�ӽq��<��8w�{B�զ}��k�z����Ʋ���m�v�R���fP�-۩�u��훳ٜ�!q��U��f���Wu ͎f�ū��'��-���{-�6���K]��1��&�X��%�l�qNڮ�nc[�Zn�j��gs=�;�W��	ffUr�teG	�4�Ō�ծ���k7��.�vS�|{%�g�$�W���$�HGuș	tS+茺9uy�-�_Ё0��$��?��gy�&i�Y�Kגg��Ha�է�w�h\�N�^�~1$���;�"��6���
~��D�a�4C't����*��#L�^@$�u�I��'ׂo�l���O�	$�[�@*|�2JwzD�\�0$RL$;$Y�	M�cT+�#Y���m&!����A%���S�Spj����� Sf!-ۥz�ذgv%��3�YSd��b��%��[^�{�� �o! I(��L�^�Р$��Yzjk\���;"�̴2�ҸLX�rL��s
9��U������K����~�}{��.���b+�D�@���H%����\�yf6�L ���xB) ���"R+)����C;*���Q�y��������i9sFmwvЅ�tgf�%OƋ�z4����M��l;����ֆ�WsMe&�olh.�X8-��9���c"2(C!� P P�ЊK -�{�}�ĀD�H��Q�a��B�K12h�l����k���'��m��N.�Wl>��W˝#�$�"9����,CD⌣�y�o2*z�(��j�P�J=|0U����d��ڗ~#�+�l�eϬI ף9�N�R-䕻l(�G���gN�
A&M�Ɨ�2�ɏ�S�̑E[����3$oFs�L���r����Z״2����S�	+��(�0d�[�BK��sوM�������@f���Ļ��M�Ȭ�a��Ţ���i`�+�i]�܉5r`��,�̋;�)���]S� �H�ŏ ��	�~00�V���#�����]��	Gk�Y� ������
W�ev߽v�L��ۡ@I W��!䀕�6�e���4����e!S���`K�!��y�UKiT �$L����k�e�|UQVQTsG�h糲I�C�o��;sU˩D������LIZx�}���T��}�0?z˾��z�����+f��/?r���6ǳ�69�x;S|=��zf�\[�;v�=�<}�`Kc��ɗ}s���t;�����gw��M�����A����O�۫\ה�t����w�|��ý뗌���H�����
L�ث�Y��WwtL��]9୵�Y+�U����9�9n]=�;jT�����m}����K���IDӡ �t^d<2��g�ڷݭox�9��+ Ӿ�����\SZ�]��_������z<8�����4�X����ކn�]1��4C�l�MML�)���7�*���T^��b�d���1��l~� ѹ�Nkq������=Ig�?w��>}=��}�&�j�NM�xM=�>��@ŊT�-�L~���7��3M�o���t���y�R^���b�!5�����'�xv���`����k�f�j��װ*N�ʣ�/��ŭ���Y����1F>��-]�$�U�{�P٢k6��Q��^n�Q6��,=.�7ϻOzu���:z容��q	����=��G���aa�s��]끽�svvP�n$шSu�v�CY��5�5��o6�9F�d���q��lL��¦�S������_�����������঺��6�47��bv�om�o����n���d�8/����O����~��3�����U�NN��xM��dľ7��<{i��C�2�>���˧�B��9%�m$����� *zR�ϖԒ0��Fa�9&4u�c#�2�<���Ǐ��}>�u����}>�Onvz�����4w4�Zt�ƒRKX_�Ub�*�.E�^e]�ƪ�]+�������>�o����o�����3���LM���'�!r���LRP�
R�D=��ZZ��Bd��.x�o�u�?�_~?��o��n��IF,�#JA�1�Ԥ��b�H*'�'��*�"A
<p�Ŕ���M9q�%2s�h��NO9�I��	��ӆ0��a�<��'��wb9�I)'�o��&��CC����i伲���E�:X��é9"AND��a&&�<�L�K�ؤ�0��&$@���%m��"TQ��ĨА��FO��ͪ��&��������+99Fseb^���:Q�ed�"0� @H� k	�(�"������U �Z@����!ҨD�@�@ʴX�2
D������Eb�,Ye`u9}�"�������"�Q��T!�W�H�B�*�u�{�z�>�f@,��$�@ 3���$/�Y��;�;��ޠ�w�q���[�@-H����I 	�m/I$Q�� &A�| Ŧ}�ݙ�� P�[�E�,��ɐf|�%/f�~.O��z��
���@�*�d�>��kt"a$k��@H�����f�|�A��M�����x�i�Cle���e�3�k��4�5Ĵ&�F�qv����hALᝑ,�ɭtG� �	-��I ~�2���H���76@�`$��{1 $U*�r�ŝؔ�a���|o�i��]c�Q�kZ��2$||_��j!"R|�	�K�>�A�������H5�%�x2g�V�W:��k����2ݸ�d��M��k�<7Ob�H��3�D�	�D�Ck-����C;*�]
 b�7S�G�o�z��) M�����%��@$#���ZR�͢E=8R���|/���˼��- ��<�u��w����;S�G����y����ܾkd�H�6"vp�D��3�����i	80�C �JF�T�+��y߾v�8t�t|�ə���ܖx����D��e����A/C]�zĐ��Q 	 -���W�R�s�	-�uWK��i1�VD��jS��Kś�=�q�n�1�}���:���z�B݋&�Y�]���b�� ��X�	��5Vį)d��.��P�[e���	u�?�^	$��"3z(hAZL�ݑ-]�xh �H���]�����C���-���I ���&BY��c�Kࣅ���e_s@��d��r����,•Z;�A g���?�� �m>R��[4�~| ��F����y��K�獊3��8dJ�n}~+:[�Ζ�,�I$}U��e$�J��	�xBb[�V�Fc��3�Η����f��%Ð��{0@4KD$��3y�̖c@�j�b� u4e�	.ݹ>@$���`$���hֶmk��:&�V���ֹF�k�P��{f��u���5��d�w�8�1Q��q]6�mh��� ����&��3K�̀��Oy�z.��r�w����?c"$2*C>�Pa;�z�{0�eԅ���<$u��u��L>������C]���-�i�V�h
qR]�����	cM����Ǘ�.���,Қ�kd�We�:��Mz��l�m��v��
v�6�k���A��f@�5�c����S�]�R�K]#�����D��^��X���=!V�۷�U�.1�;�M�ge�Tf��B��-�Zlݔ�S��Z�o`N�ra�&�݇��@�3�';�o�fvwvw,��@1�0#��$���@�^U��	5y{�vz" A;䐼׀$��m�aݜ;�)���%Q�
�S5.�pI��[,�ф	A"ku��AI,�3_sD"���k�ۭ�v�^ț�v�Ƅ��;��d�� BI$��ƈJ<ވ$� @�3kf�a� ��?m`�Iy �_<[��d�_4z׹cݙ�ܖN 7�������ⅷH�J_Y��$�^H�[<�H���F6��v�h9~�S��%���L�*dއ|n9��#�V�����`]\A�%�=/��Q"[_�
򶧫��E�G�T$*BNK��y���nwD�{<ʹ��Lh�!��f�n�ړ׿��'��p�'e�w�ߢ<H�-����~#"���i�C�%y#m�����$��ݝ2/l�������<�9��c 1O�����*v'�=q�r�F��bU�����k)���"
���[
d�"%�:%��l'V�'��{�T/�+�~�Bpd�^H�
��)H�K >����ڀ@o�I!�����U}��K�cU���_v~��o��t��?l�/����*3Ս�{�X i�c�$66���V�p���It�{�׭���>�q��+���/��]L���!������dY�T��fޜ=ܷ��ũ��m[�hJ��뛘��qXd�D>SY�V���X �S8>�̌���,������$�<���C)��;��,�@�3��}!��!Ͱ�	�s��2�,>$C��r�Q�7{^�)���?kO�<�K���۫�26�ݡz'qIâى�x�'7v��v[k������l?��m��/�;=/6+��}�� ��&��M��yp��9���e�:i���p�'eo��2H+���e��i��S=< ��p����"7�b'wEc-�ݻަ�~��ƴ�9wp]�xe�!k�^<I�0�+�����5D�S�Yy�`VU�޿���w����%�?v�p���}�;gu˝�ɚ3|���_K�þ\9'0�DO��B}\C�%(�(-"�(�*�η�t	���$�����7�+
N�ᜲL�TA*�|�j��<u�E��pu��l��w�`G�י�_��Ė=�s�7/�NՒ������h�u���9�^w^KgX��>;7O�x����A{�n}�o�>o��� �G�v�T׬�㵸�&up)^X�4���^�z͇����|��z��}~�my�2��S�����~���PS쾈.�ӱVǸm��ߕ�A�~x���a���;�Z����$#6&��j'.ݟ@D�{k�$�F�ɵ��0�.q����t����bA'��2�/�.�n�"<A�� K���4��q۸F�Eu�A>$��ަ��9wp]�x����og��n'����6�w�x��}H;��v����WSI�(p�v��M��ċ���6U�޻�GC��Na8����4�x�b�ڞonû�uT_��`%S ��� <8x�xHeT�Q�Y
��u����l�I��0v)�d�b�@�����']��-�q ��AdvG��Ty-�~0^�/F�3����0vv)��kzE��tv��:�x�,n�܎�3�j�]0�0\��R8����
�A׬��A=S�$��/�<L�wk[��m�\o�����H$�،����wwd];�H=�o �3� ��-�Z�fD�߉$@=�� #z�=>7�0j��O:{�"�w"b��-2l��M�?��&��a\uĻ��E���7�����:�\vG}\����FS`B���	 ���	/��ơܮ����+��RL��L̗n���V������73� Ef\�$�!�ٽ@ۇL��Z\�R��{Ym,0Ӭƅ�q`�ll
�i�
�}��%����w����v�]D�pd��������9��H�f��]f\��:��}��@�c(�0��80�@�F��	^����:�ݡ������zY�E]���X@�mhh�W1veb뛪Z��KV�q:�,%���l{BQ��]� a9�	Y��͙��H/�Hq����9�X�b�a�-�4�A�h9�"9����������[�k�	M���n�A������1g�����69Z[d�n�$����-�ݥR+b`��5�N-�4B�ۮ�N����K��	�!�K��P%!�!w�Ͼ)3��2g����[o�����{[5VBt
�C����/6���ݭ%#� 这L������@�/I�MqN,'z�A ����qd޶�4�=�i[���X:v3>1�O'Ğ�ǀ'��r���w&�H#�v{:�Œwۜ��L�����;�Z�'ۇ�^�/�.�x�F����� �EqeIflm=`�z�Cy)�l����;�5[�=t���D H��n�9c�z�;F��A۰�r�u��釾v;�4��h_'�.��&��ur�vs:n�;/�.�A�/;sM4&��	�����}߭���J`^�9;. ��� �v/�� �]���Ʃ���Y��f�e�L���&{�p�T�J�fx���m�D���ô����1G���/�>ӳ��w2M��OwU���G>1�X�-��f�M=u�]�������z���$~�Ea�B��J�J"s�ߛ����ϯ�	$���.9��h�|�QĤi$:!�
�����no�A�n;ǝӸg����{�� ��]����.�僺eޚ2��s+Vsm��A��x �I"�6 �}� �Bƨ�k��oB�Y�x�ugy��;�X��i�<{"�\Y��N���l��I��Omt 5\wT���a,A �ir�����q�ɡ���/�c���\�z_v��{���5����<� ��{�n& 	5p���I9�� 79k�s��꫋���c�#sz�[$�;��'� �;�&}ܭ�h^Զ����y�w���A3�����c>7ͺ$��|OXɒ�;�%L�$�l@B���LA~���ζaj��/��q�oʩ����W�k�'=�׼xGl��ogP�s�;�\̰�=�K�y���&���!�0�UcT���A��H�(�ձ�7�/�L���n��!H���M4�A���;%�X�/��8�=��X0 N_t'{A�Юq�{ė�؍����k���X9v1 嚜��|I��x7�Mn)R �;�Dx�E�t�"H�ވ��������|��5���,j˕ڐ���݁�cha�ɩWmp[�95�b���o��].tK@���=8�I��_�*^�ޘ�hm�3�+����� ν�H���������>tC�L*��M��5	=׉�YW(o_;�$�k���\H/�q���#Ā^����5>�Um��H'wt�'�4�Dj���↮ǛC�4�Q����q��@�V�dA"xl�E����y7Ls�#(kt3��x�c���n<�@��B�d$�u���_3�>
])y��C�ؑ6�r�5��ӓ�>x�6�[^cD�ݳ��
X���e^"����/2�<�nn����qި^��G燀�"�0���P�����c~�'/`��\�2�T}���@�װ"9�4�t�=��%�3u"|I>]�$	H�v�m^��[
;̉p�Iw2�v^�X�3a�=�7n��ѫە�;��a��G"M\�&����2au�o���١ii�}�ǂH!�� �U:�4+ʆތwH'6��#��]�o �3�wD��9��9U"9#a�t]2�k�s\���@��[��3�H0\@��^-قY�6������:2x�o����	�[I%�!��#Ʀ�{8�xڪ��ʼ˱�#Ē��{�>P��6����������4�+��NP7���w^o$H�}���3|�b��Dx�`�6QgwD�鞤F�vp(�k����xi��-=Q� �՝�H��� �U4��v[�1qτ�e���/e�Uz����sj�wL��C��S���x�GR74e�����g�c%��,�Of���^����/��Ϻ��A�r9�\W��J+F{=���^�rJ2��PT��e��y3�n��c}���=d%�\;<�{u�wx��R�(�w��6p�k��bzc;����ݎ<���'w{ܽ�~�����N���H����Ƽ�^t�մ��=��o^����I=�@�ǚ�aӽ�>~8��:Nm���`��Ż3��n s/r�ޅ#����+�t:�Z9r��G���*�>��"�37�qb�?6U[y��uo��}�zΥ/����D�a�ܧ�^0�i9�N�W���0�
��d%~� Y�_x`qcLf�f�|)��	�lf��Hu~�v�<&��;Ow}��q�
c}g��6|W��^�����q0��'���^Ʊ"v������N�}/�k�w��ݣ;_h��}�G9���.�����xO�߬z2�U�r���6O��}#.�|�S��0w��=�r�B�/�y_[��b����j�(Y	�.��w��l�B�^������}F��vq񸸵��t�����.�#W�f���e������u��w����=��=|��{ޛ�	�����U����f��H�j��8w��9�I�V�{sc��dk4ԏ1}��K�C�4s&�q�4��S�,ƂeEٵ�a��7M+9���o{=&w��U{n���������8�v�:4�^cD0�7��Z>��7r������܅��,���5�v�ރ/�l��珐8��ba�b	�I<�F%/�(�-���x���_R2èf�d6��HH�)X���.\�<	��}��3��~�����~WkU��r�[��1�$�+���8�H���N^W�*��)�^ aҬ�)&�Db�X1>>���x��}�>?�Ƿ����������@䐀1A���gb�$�&$��!R!�b��!�,
�	�a����e�=����~3�����ooo����T0j�Ķ��X�1�(��Z$Y�X��(Z��Z�U;�r'D�����@;�+j ��؜]���	�S�p@���Nı���+�Mnip� �H#��O�:Xt����R���Z-�7m'�R��"^pqFj�	�RA�*�mH�}'hmU2@�(��V� ��cX�ֳrdPݖ^�,%b��Ay��(/�H�(, �99�� G��':1:�&�u"��P����C�>�i7�RE���Is�����l|�=���MP��ԑ���^u�[m-��iƅ��%��	�w����5��oPn$m�F�����3�n�5IC:2⛁�MF����Y��gvL��v�ӕ�g���������7/��u���q��kd��7E�eݬٍuI�=��^�81��Q��7�����W����7ZEV�U�Rf�$f��!q,�'��� Mc,�.2�t�U�d�Q��bC��n��xv/d+�^�Z\�&.T�,f��tΛ�+<>N{y-+v����ȉu�p��g9zX��C�Gg��w�l!-� �u���{QV�[g%G���Ŷ^ݳ[��9�@R�2�-�am6�i�ն�U�]�عB��w!�k���# �'��)rLᨥ!��0i�43ӹ�b��d�P�n1�<�)q�ms��8D�٭��^ztrvՉp�mk���38Dn�^Z�k�8�v�^R��6��v��-%�"�ZX����U�4p��mÆ��=s���lmo^K��j��4�g�>g���[3naݹ{N.kdV9՟�i\hڢ�fw����Ҟz�m�c�q��kD��rո���-D�uY�U�i4�����ty(�ܝi]�&�e��_��X�+W\���{s�¡c� ��VQ��P�"�ӝx��ѣ�iU��L�=s�8����u{j^#s��=�f��Su�]�2]�[��_�3פ�^�;3�e�+��볻%�J-��\�lD���'X�s�iQ�m��;��u�Ѓ�柞�i"�T�٣�[vՙ.�M�6���S`��Z��W@��AIV��\[����Oi.��Zz프�-�l��%Tb[Pźy�N�z���.�6-9�������/`
�$��]�sn9�uqō(X�]�m۱�n�BSk��*��SDf0׌K۱�+�J�:뫝�W��/c#�62c�`d7�Z�uNu���i��2PC3/�M�Ry�b.�o*C��.L��ؒ�2�S��'I����#��a���$��+����zK�|�iD-F�	�b��eeж��2��bB���^�h(D�m�3��Ϭ,�p������#v܂��#<����ޮ����c��Miye\%��s)��[N��Z=6�^�l�<��:y���ڙ�q����'k�O"�9�Wh�l���SL���٦��]s�ni+mHV���v��wm�ޒF���^����fb6ؽv����ӭݖ�L�X˳�S1�К�i���,۴HE�\YxK����/��f`�~��>\̷�!M�$�G6��;t�_n@����$��v�ɫJ���8o;��Tb5���zwe������F�L�M��	pc�r�
n'�V`$FB�$���>.ݰx�c�y�;6�*wȺ�[-�H$���z'__�$�6Cky�b��U����ML4�Y|��lO�(��D���趬�0�m��ּQn�x�ؒ���d^d�h��� ����pmT�Tk�{�w�H'�ٱ����x/|��4��7��*;�
���δ#^0plј�r ���ABd��u��������K�aA�?=� �e��|g���g<����lB�Tv��D�l&6�A!Q%��0e�l�����3����DSw�ҦJ1��^o|[�gh��ImmWB5Pj���UD�N����eC!n9�g+vC�R",z8�D��j$���F�S�`R�RN<�V��ח�r��>�ϠA�����22�jb7��^d��bT��;�������|W�{�$�SD��r���Y�H�́$:��J�>I3�v	�	�^o��_g�ܼ��|��fl"_�i_A8�,�H�� 1���o;� �	���	���Ǣx���gt�TϬ`���<��̈$��������i�z����M��f�T���,P��u�pݞ�t9wn��(;8tK2=V����3��t�ǉ$����H���
a]�3!�C���lx5�:#�v�	���,Y��('g���x�-��g;��+'Yݼp�@�̈�@<�p��y��T����}��\˶칽���ʐk���K���­�1ȶ+k���6,v���bq��7/U�r�ȩSޮ����|?x�^��_�?gT�}Ӗ�����E��j�,xʪN�8�(���x|<@���aHeNJ#P@)���ߛȃy�A��>�j]�p�vc2]���A�4��({�%�ĂOdcǆy"�����+�gi&ꧽ3�U����LᝂcZ���o3Q��ȯod��G��{�#(�S���s|��u��	��a]]�>��77�t�qV�Q�ۃ\p\���|�Ι���=���r�ˠ�ᱱ'n-�|<H�ށi�5�FO\H�'���D���ooX8gwv,��n�f��ݐz-9`�6���}��~�-����?D7�>0��{ʓ~�;4M�,��$��̂�؂Es�Š�Du�Ƶ���c7<H-�K.= �Fs�'�y �LK:b�2��zD��{��=Q��A�$	����|7�#|�]�t>�̻���F
5Uu5VjbM�Ub��ș��l9^�Mw=���999ps_���zL;����5݁L2�S��s#��jc"C��tG=c��~�N೹!���4#������x-_d��hn���UDz<�Q��-�[� �Rr�#6��H��P�����q��c��4�t�5�;d��m�/d5�e��	�����ߛP)p����\^; A^Iyn�x�9/͝[b�ٷւ�d[ƭ�����C<Z�ނ�]� ���X��N��NAv ��������ƫ��_�	$��ϐ ����|y�Kb�EkF��v����&��;�.�P;�A��q�t'vA9�7�dk�{-�@��B6: x�b(�����gwI�=�7�(j�U�@5�O�wkǛ�9�kjE�%�:=��'��݃`�R�ؿ H/�;c�э��1�/�ў2	 �<�hI�툹.�>�t�w�W���N��i���h�������f��R2���`�xj�p��x�c����zܸ_x����՟~�/�2���32�����H�eB�� ���׮ι�i��?�s犛�l����.��.x㎅��=k�W�5�9�m�īnB��cl�r���ȶ	�#�m˪��1n�z�,�B���e!:ݖn2�������v��h��G]
�nWK-�)���!�����*&IɎ/d��:�=#˴�q6�
��nm�`
�S�C��y�0#�z��k�ZUs/�;���رy瓱enwD�Z�t�T����<+��{�Bo�￿�����Ki�����׀H>���O��x�2�
}�]3�;����� ��0&�x؈'�#�ǩ�;��ȏ�O=�A$�k�}鎇j�]-S�ޯq�l�����km�ִ(+�s�+�[�/ُ���ۇ��*��켢l1(�����u���!�緡1�^$���	�e�<I9���%e�x:�ϛɼ��:d���4 �d�K.џ���>��;c�1K�����D��<�8�� Fk�-Q+�x�����f<�� ���d,޼�L�o[�w\tg���hXʹ��.�ѭ4�uy�>Z���#v\�Y(�g�I��~1㭒�q��lHΙ�[��q�=�ȣt��'gL���1�� "lS��]���/a��b�s!��M����q~������~ͨ�w���.:Ɯ�=0(V����X;��]s��p��>��@paH`.���D��y"y�">?|��Д��JJz�H�ހK꼰	�Z��3��0���q�A&�L+�\�kf*�� ��������"	׳Z��仠]���؍��8م=0�\y�e�xA$�;Y�A��_3H��e55VĞ�ȃ~��C��ÆOT=��Bz��cDv* ���;]���_FzBʓ�:�y�Ӥ�o�nmR�5�n:3!�8�/Bg��n�q��fܚ�(˘��N��32�#�>>~���J�5?C	=�� `i
ER�����w #��#� %�;"�(�O<U>�Ҹ^	s�3f��9 ���6�#ă���
o^nOw?
z���Y�����f�%�}J�49A��x����f���(�ܸ�7&XG]�٫уK�o%:;���X'��^�,As�vO������.�l������K�+f��ge�C�y�o����C�u��=gڇ�݄���J����ח�^T����(�����Ġ#�Zؐ��d1�T��Z^�j}�.�j�$�������_��-�ٴs(�k=��`xp����Ue��%��"H  O�\[���[oУej�&�\�Ə [�^<��{�bl�X����B�wbJp\!�,�I��!��M9×�ޞ]��m��k1�;V�����e�K�p��������Q��x�	ѱ ���só60���B������^��p1wwdN^�e6�&�����d��{���m�'Ă}Wy�g�x��N�#�TUv�xD���w��T�s2XL�@$K;��(�哱 o�_N���y L�vc��wY��'���@�E�-��^鳔Y�����f2�v�뱨�!:�H4�/��>����$<���g`�x��;�Μ�g9���fhYf)ޝ��)7��bsCغ�4O�jҙ�v �	��[�4:��un��@��������9Ϡ~�P�R�*}��wc�EM�6�!E����*�����;󁯪���ZZ�)�<�u�̺� eSűN^IK�3����z:D$�^�m]m/n����<c�uq�.�Dݿ8/�3�仠]��In. ��$c�r��N��5ݿ<x�|o��>�vh�%�N�;��������I�%�u�]23�)�I����u��@��e*"�܆���*X�vw(���ح�	&�w('��ڡ�j	�z�ldI�x�$O��z���H�wf$31S>];�8CkFG^0$�w@�A>�׳��}�fѷ3`����\i�)��˻�f;�b9�$7�{���\<�^�������W�z�>ݞx�v�3|�M4�r��ǳ�2�'ӵ9�8i9s61j`T'��@�*詸˖��W�O���dn��AJH�M���/�M���	��̍�L��.gs]p�g�c�˖:�����C;!ɜçw����S�.e�`�J�%�Vm������� �]��zڪ�xwM��4��aS��m*K`֪8IR�c��M�"8�:K0���n/�o5��5��N��n�s� `�:8������N*�eܹ��Fj.�F��Q�s�XH�fcAk�]�&6��^�j7J9��tm��b���!dk��bjH�R�Z���i�G���az�v�jV�Hon<|�,�������:2뭍G*�p]��kGC;:���<�,���yP����A���?�_[��?Dz�<�0 @����u����vϮ�EٚF�a�G���z� �%��ǉ'���|�q����/�2��{��°����M�r^癈 �z�c������OG��0��
ڲ-wgg�|J�,\�;�]�����{�����NY�|Kl�A#�"}W�ߛ�N�Ds���D���g��d�w> eM�"������ '���ے2�,�y�:[q�%o $�o^@�AލA��q���A���Y��ˢ�v���۬�2�V�f3�]�P�"ͺ�i�Q#�l�ߣm��Ki�����:��q|q��I^э
��:�Td1�^c�"};��Ȅ]:.R�^/��Df7s1��s[�"��$�.�ܼ����uwx9xZ�e���U�y��C6�>͏���ܛ�{���p��ׯW>��Xaa�{dE�	��:�LiO}���(�߼ރJ��F�����0G���㚓�`]�.��K��$A˹�A'��=�^�[slF�9��؀H$��_3D�.�;���g�ɝ���!+�^�$�v�}�@ ����_�B��qJ=dT�xɎ���w�[.��:f/B��DA���S�O'&*_����]0h��@&k2]�(9��AR��2{���C�qT���1scOG���7c\��Y8g���^�����G��D�v�F�w(�Lr�؀	"v6�|@ox�O8�7�z�圅��/���G�$���w]�3�vr��Q��x$���Ӷ��Z��]�3��> ��6 I�� ϗ�ܭs��x�D�۱(�gb�!2<[�c��U�<6@D����[˓��俒�{,.ܴ�������:���g{r�K�^:���x�|v����:��8y����ۀ����N�E?%���-&�юI�6�Y2Y�d��[�X�|0��Q�z�uWZ��[��RY�^���"�l��)d��9ᱷ;��x/M.��t/]���y�������|w����{В���3w`'��P�f�o=��"�{xF.�^ݛ�"����ꗙ�mQ�Y�/jB}�ľ�F�˔\�9���bÇ�v��hл�橞�$� ��4���pJ�Lv�	؇��6��
���c��N�w=���٩�ػ@���+w�{�J_���zj�����Ru���w)u�yç��a{�bg�u���|�j�spcĂ9$qR�
�"4=��睢-��|B��O��{�ع{�RQ�@��!�>�F������scg���f͢1������~^�y�_^]��.�=��-���]w�q�W�gp}"�3wN������{),�ׂ�����vy��:��gϫy�=m�k˞�W�!�f��oѫ8޳� Rż<����&sP��Z>�<���Zw�r�n��:u8�F��j��ܩ��8y�!
����g�'�.�͐s�����;f��H`��� Uz�^KgM=�{�F���:��j�<4m?7����j� ��_�>q�]H��o�z~�mB��3�0��+����j�"�c��cgú�G�$��m� �B��'�z+������<k���1��	 w+�99!����K���K����J#T� �s�9s��>��σ�Ϗ���~=�֫���f:d��8ƳD�ԅF��"�Z�eD �F!#)HRN��,�\3�Fg.q�������ϧ�����{{{{}��t�A������H�$�Ā��x�;��'+'�'ODI�+"�Ex�Ź>?��3�~3����~?����o����[g��$NcrN�+;�-J�8H��C��k'Οf��,�UB+�錼 �)e�$Hł=J�kH �=u��H��Q�X������	�����ADx�yE"rI�IN�# 0�`�+�Y @9&5z<#���mT� �"���dk��C���*�/ t`(Q��ȵ �$��	b��I�8�-����DhF�b��QJ$����DC����R��G�dşu�D����ᬵ�k8Vrj���Q��qZ�1�D�T���u!��}ԡ�[bA���A�n)&�r��{�e���e!� yχcD|I�t@ �[�G�MTY�IӰ.�azݦ�}X��ؼ�I�x� �w]��9��m�� L�n��K��bF:6kNN��)�A��h�sAO�&ym��J��t�dkK��H�݈�'��H�Fu�An��E;���C5�Z��v��Y�vu�а�0�^�E3�[K\�/g��0�0,���xg1wN�&b�;�b/$[���(�Om�C����ҍ�f�uw�s��}�:Iݐd�4�踀|͝�}�;lT�d���	�����G�s�&�E�t\�����]��)�3�窀1� ��q����0PL�E O���E�{��<��c�	�gb�!h�;��]��.�+O�y]�%������'�c��}���zd���dW�;L�G�~o��鎼�,��y�vǜp~�;7�Ӟ�C����V�O&ȗ-d���P�x��|V]Z88�C�{��'80�{�{��G����+ԝقr�	����I?\\Cdq�"�Q�J�9��{�q�y�Ex��{��~֛�v�r�/2v�9(�E�S68��ѷeW�%�]2��9?�����3F��f���!��'o^��ȿ�1�s�(�ng��x�{�E��D�'ggt�Y�^<� �����F��.�u{:���!u��H�F@��^+��7���g�pAڝ$��̘(�F� IQ�{wk|�9@�+oE�H�܈�H=ё�(�6.��ۖb�ݙ���:a�_6�e֝�#ّ�$��ׁ>H����z��9V�h+��@���p��w.R*�螈$��><3�����yznn@��H��M��@�/��R\gU��e�Vɇ�iJM����ܘ��7[V2U��v�p�7��(���yix3�2�Z�`5��3'}{#5�kr�B԰�:{;��I	Đ�rt�"t�o�ZOK�B��E�K]f���6ۥ.�f6XM���t�,�f��s��מÔ�Kmv�Sk{ n����#�bM�9gq�J�Gl�8ܶ� ��K[/5%�z�bΦ��e�g���� ��qs)�������Caԃ�U�3e-�J���.'�6��%{/mq��榥����+���#5@j�띴���e^�9�6��{fYE�lj
�H	��`3l��Ҫ���نc��}������)˒� �uL@$	7��H}~���3I]x�����C
����I$��<h��Maᓻ�� ?��-q/"Y͡	w�m�=	$���ͽ�q��خf�ږ��t٥�;�h�I���spty>~�p}�Gi�Uѽ�wF؏���&:��"���3&
PhK(�}H|S�DO��{�� �n�w˶�.Vc��AΡ`����٘̂�� �x�~퍉2�W�<gn� '��Kv��H[� ��/߿Y����tv�f�lm�47��nGK˩U7':Z�
gu�d�� �������fw,R��żJ�ǀI'+y�t�K$fLu�z^G�\A �f�L��9r]��븳,���\�%=��ؕv\E�K�X�Xw�/�KK�������c#�k]'b<4ºZ������2���Lp? ����d��7�_^�#�y��O����E�>�AܐY�i��;S{��D��tS`D��Ļ@�s������!Q��FٟU�Ok�<Hi�>��"��3�HkX������y�A渤YH}	�m� �~���@(�������׾�� �Y�����x�������u�{<�{���/�� 䅾�h� �	5��"��7'�F<#؉�w� �_�;�`|	=�QKG���<.��9Cv%��%ctf���eD�!�Z�S��Ӏ��S5-"9�����32���Q���G�n�<x�G��D�m����X��)��n�;��m���3�E!ANň ��禗e�s�2 �~؏|H;�Q<�ܵ�'�$A���TO]�b�;�t]�I7a�� W��&�� ��{��ټ��3DK�1��T-w��;P6�_|T����r�+ޡ-CA�`�z�d+ņ�bS�
ө`�������W�L{��|�/��`�D�'�}n�򟯭�������[%8fvEڨ�'��
7".���M�I� O^�ǈ�d�rt��qD1��Y�b	��і'b���'��U���W��]i�bz"�O]y��ɝ��y�ި�(��~PZfT4��~���<�����k��C],\��<iY<c�U��K�n�lRR�p2�h�ϟ~�?��9!����D�LP�m�dd����±�N�Y��=�jD��wfc2�ކ ���'�p���ٴ�	$�vd�z��Y�u��IU�;q$��4�猉�7��y3�E!ު1}Q����}K
f�$}���� �w�I�%���ote x��3��M����deR�Fk-��H�m�~��'ݹ�!�g��xd�Vv��df�]�?����Zqq�>��ݬwbﳎ׻����<�Y9�����b��a�_��A�"SUB`��0 ��4KXA8fN��
��3�����	�2��"��=@�jq@ ��Cx��㠳��nĒ\:�b�7AΫ����O�-a�]��J��F��t�}�?o����S�I�A�� �ӑ������ݾx���l�[�g�ǫm��톻VH�k�"Ey�9!U��x�? ���o|�,��u�@$��;�̡�����a,d�p���b��wn��N��� -|�����ʙ�œ0��#��vDxW���=|j����8t�E��x����9�Mf��A����t��K_=���-;��p]��7~UH�:�\������f�͇�)w��S����u�N�D��h���BM�|��݆і�LP�l|�~����mm�~�oH�DP2��@�cv��7�)��~-Z[Yk�y2�OfnqU4�[��F��7�������[7o"���8�*Jq\k@׀��!�pi]m"�#��А&��cH٠ƃvQ״*)���vH�7%Ф"�qx��x�\��5�5�z����TJ��n�Eٛh�+�&�ݺ��JjB%�-`x�Pv� ��:�pY����<G9'���k���<�'���	�b�sn���,��6�1�E���O\�\L�\ݷY�>��k��'H�ds�Xˬ�m��1�����;^�.��,�C9An�1��E؄�;w���x0D��� �N�B�@o-��������M�/w��Dgכf���wwt�ח6>x�Qڅ����NyF�D@$�D@'��4�fEv��������TI5�~z����?D��w�n�1-;d�I9�� �3_��qd��çfcY��T��M�3&W4�~|���ܻ�$�g�"3z�e���	�e<�� >�1z�E��)
��[ƹ� A��IzWFD
��[��07d�T��K�t ����lH�iwgg4�{!��$\e�p�ם-t�l�C�t�!��P��;�8p]�l58�T���"5��o�����T�x�@+2מgk�E8E�v��!��C�2���y���wr��?�+p�υ�J���	���wG?f�]r�CwE�������*N�w��f����_�)Jj�y�K�>�$K_��H�@�A�^�A\ǀ���	��>L䳻�I�X4� �^w��ļv�ؒJ���@ �F�@�H��wR8Hr�� ��s��ܙ�ξ�G������ �Dfl�">�����,Ψ��O�ظd�@� �l<xI�x7��e7f����yY� Gol@3{�V�����۰`���-��d(f:-��q�MuK4ı4Ĺ!����~ϟ~�tHwt�C@�j:^����	'��v�x�Fe�b<��K� 2�w��9H����Â�&z_b	���G���F �|�r�'��Љۓg���ce�l^@�p��$]�.��
�
؇�H$�ǀAn걱��B��nೳW.�7M���٪L�Rd��\ST0���^�.�90&����Oyk��������v�<�<�]�;�?�R	MQ�k��Ѿ$�M��� �G��DxΪ�pY�ܤ��������I��d`��@9]��w�ZΚ6�t͂�$tc��R�N�$9gd)���� ��^]��1�Cz�%��Lג�|� H$u�DN��@;@�:5��$)Lt2`�����J,q�{R�+�V4����]a
��0x,�G9p�����mpb	��9� ��؃��̨)�D�r�Gws�7��R���"���燸���v�[R�wC	&�� x�	y�!x�{���O�n#9Ԓި�H���8.��w����0)���䁵k�0�3绾P_��3���=�;�)��d�����)��2��,V����O�7�	��]kax-=�!m�O3\⧵R�\�c����9aBӑU{���LL&ʭ�}@�^����%�5�t��s��v@�<�uߏ�o{���;�9/�~)��JT)�7�1 ��ꠊw���M"Jۈ|E2���)���D�ԝ���}I ݽ�_�lf�;t(�}�n���:&i��k,�K4YV;�u�\�� Jű��z۞G5��ͫ�#��B�}�����ZE���9��J�^> s.�d.�{7#j4S�鮛�/䉫����dK�	Lb�<�ty��,�l:v;;�3.]��^H�]��x�']����`j\fc�BQ��Ӹ��1$3�E!C'ۀA�Ui�w	%v��}��.���Y�$��؈(�F;wG���5������@�Ϻ�g8l��,�;& �	�Y���$�Cwd��[���O��Έ7��7�1����!;@�ܞ9�$�v�ɢV�{�߉���@�n�ބA�=� no�Cc�AB�S�Hv���=
ǖ�;��]�.�|��ߍƱ��������2q����]
���p���JY�w(9���V'��=�5����q޹Jr��N=��[Ѭߐ%S��.=��}���{�1����c��?)QN���~/=AG'��I��1���f^���<2>�s�����t^J�=b/ydI	l�ٽ
y�x����'���!���{w�h�b-�^�Or6w`�_v	'=��ѝ;������{I��7|L3�]��ʂ�9���1��Fвݞ�]�=���zWs�a��//���LN�Vuh��]ؾڻĔE�+g�>�2�����5��ݷ��G��}R��s��8{��o!�f8��	zP䫛x���q�0[�fՔ�&�-s����9��.o&=�3��%d�@ɻ�`Nnָ'T�ȝ�hŦƬI���^�~޻��Y�{ov�(�p^(��xv��Ǔ87�Xۢv�����}�c������'�軱-K
�Qw"����e�t��( 7��sN��	��*��ts����j�� '{�0���;$��Bj�hQ'!|�}ȩ�R���<�h���58w�/\�k]�f4���c�vvk��erT7HN�6��n%�D<��z�}z7<����tv�����}-�)3�4����$z�,`M~��!!{�`�hQ��nzIq��-xC��\1���{�M �����<b�ۇ�d�!��{����|;) w����;8����m�&��&4'=ط/°�$,"c�[��E����<y��$��OҰL�2��G&��Ĩ�(�
I	~b��[�Ƕш}�����@�u �+ N�	�U`B^�����o���3��Ϸ�����{{{{}����!�"F/�I��:KE`'>Ƅ9
�$���G��r���~?����|u�eeeeen�SU��d�"�QbA��0�C����傐��.p�u%s����}�>?�������n�뼞a��# ,�8(R4�
��$�������!��'�(y���!�ч)�!�Ӥ�D8��E")z!�1 ��� � �U��F�Վ�dc$�#B������Z	 ��� ��,���tFLFS�J�!�H(A"AP�"�2+!�(/�R� �՜�
�R@��A���we!�U�U��25�B�R$G�FAg�"BQܕ�y�	 ��Vz C�HA$�����8z�Ń�'��5����2w�R��5��k���;>˺˸��6;S�r�N�����^}[����M�֊��:�W)�&�Vs���lu�7\$g���Uy��4&�v�v.Ů�.���L�ڝ�tt�9��hY+�λ=Pa����NvY�����=�K���ΜI�֓\��;7L��E�FU��I���K���+�8�t�aoL��I̼�,���C�\���͕%�DCc���ѹ�+ͩ	���t+�Hf�l��3y7�m&�*8m�[�����۩ThG>6�tvg��kRN�Q��Χ�*���k�B@��#^\�G�Y����K��1�ق�%і��Q�M,e���'�,�#��y�ݸ��.�h��lU̦t�;v{&7D��"�u�n)��)k+y�͒쒸���kT����ۓldzcZ�Q��.�6��}9�mlm(��^f�`j���z�a��]��kc-�e,n��B�l�8����a��	3+\k���\E�+4��<����ŕ��gd��>y�᧥��Mo]�t��W]t�".�5��0Ь�+u�I��bn�w��lhf��Y���ۺ�̇gX]d3Z7��7�}��lU2�e�"�k[	�vī�m�HB��K+5�:X��6lb#��r��)`�|��y6,�l.�s5�.��������lq�Н�k�ox���5ۋ���~S�|��=����e����sK��u#�Ơq��y��ݜ\-�]F �p��ݗ4�ݧ���y���>3sh�U\d�Tu�m(���l;Y���)����ъ�H���7u��;X"��\��k�٭�D�qz��QT^��[������PйE�<��l\e�I%�X�4Y�8ؔ�nc�^�ù ���,�����]OJ�E.���u�3�z�� �:K�Ɲ�c<9��u�2�hY��<uٮZ��p<	������v�[FC�)�s�kNW��z'�-�y?�~)�J@��sQd���%1�MJQ�y�3"��2�Ka��v��ƊH�$]"�@e��Ǔq�j&�kI��]�^M�	B��D����l��_�X�h��X������;Q>Q<�NВl�EH�M�ի����af�u��k�a��]�g6F$F����H8�������]�u����m�6م+�,��5U���[R��{�ض��x(n���vׂ��#a�f�HF�ݔ2�]�Υ��������U�;\-�'�?]�yW�ۺCH�� �tU\�ک泼k&�@^K��U��tA8��!݈D�A��#Ğ��U|H���a��|��D��Q�Ioc�����ꌼ��z��v�H�.
,��N�PX]w��G���C=י��u��Ē���;Ւ���H@�.�<�� .��s�u�y"У!�$��H=�v���|�44򂽓:RJ�vp������	z�b"�{��T�"��^�h�$�W��#����_lX�Oa��� m.(�n����Z��� �ԙ��c��[�X����>�vb���=�{UUz^<��� 	���@'�'0k�ff�ҏG]�HM{�;02N�3��Mr'��["c�E�'�ν�ډ��&��f�ܼ�S��9NX:�G*ih=YŽ�}ڽ��M��^�Ǉ'
R���M[zwck�O�q�X��s�R��鬿3�_>FF{��=����5C����!�/"�6#ă�<�t��V`�m��Ԅm>�:��̃�U3t��L�l+�x�LB����ڽ��6�	y� u�#�D�$�!�$Y1����,]������<~�3x��{�~`��'�Jkn�|�b9��P�߉�Hw����$�kk�#�ݞ؞�5� �E�lz$F�G�a���%*^�z��-�
����hT�v��e���^$�f�Ѽq�0u�a����V0!��Ϣ���MQq�)ߢ$�j���������'3ļGl4{g�r"%y?��2`�gc��2,�'k��}����f[�cs��>$9�"	�9�y	 �da��4��=���sz�2vrY݃&�s�>�qMЈ'�y���7`��4S?L0į2�ǈtiNӋ�
oj��;����Ax�L,%� odE���r�����5&MrZ��6|�mu�a���O	>�{�}��
����]�ܾu��d;�O>.���%Qއ���N��8��b<�$�ͭ�<I#;�#�2I��/���b�.��	�I�9����繏Y��לn��f �vi�ǈ��x�&�I��G���H<��݆dl@ѕ�jV�qƓ`"DwaRVlbj�����`f�Y�����$�g�;� zq�ǉ'v� �_4�2n�YT�;*��m��ǎ��I-E;�H���؈ kcm�ׁ�_wj�= ��������	-�1"݊"�T��9?Fn���e�cA�0L�'i�s!�$���I�ݍ�
���<�`{s�	�����g`��$�9��u[��q͆	$Ov�O�^�aS��b^m����N*����L-�r�^1\1{�.2���u7�3E��m5�mԊp*����FY�$mhl��}�c�G8�v�wY�����m";�h7� ߊ.~�ތ��Ul�� �CqNWdA>$/��5�z�=pwuE����� �b]ݶY8=�[\�ӣ#]���X]Y�4�����6�����`O�t��G7G�m�8���9�~ި�޳8em�6�9����c�<j*�+�A!;�� ݝ���G�� �A��0�y#]�	�}�ŲdIm�k�nbfl���N�Q,+�C#f $/���
���i�M:[�7�_��kq�D�L3��X�r�&r�
�[ݲ���Y�0su� �f���X�|�y-�~5ш��!��	������g`��|��H7:�]�����b��j�o�"
N�7/F�O(k����h�Ҽ�?��F�?K�#5����P}�{�a�m��l�}u��j�D��M�B����/�oD�|�ؐ�	Ù�3����a�T���\�gCSImk����P�[���a^ɥ����5����e}x=�7-%���ű�S�qmA���4#\G%���ݙ�=Sg6{�Kd݊��ͤ�N�u����c�F��d9gɐ�i��;p�'��y�����^��*j��M��Yx�&ZdceƎ�XKa�u�����m��ak�;�yaU9�0��-�[jË�iCk%;:�a���1zɻ���t���0��:,���O�
A y����� �}�XL	 F�@�|{2��*}~0w%2c3���Є����yq���|�K�݈��@����>$���Ζ�����o+R�(��)Tع�M��XQk̀���A ��@�@'�_�}�6V�1,��LLϗ�a�r,�W��OU�b��<�����X��cĀ�H��zl�j`�c��[��=�!�9	�g!;L�s!�6D��<O����mo&�^��N�	�=�`NWt7�dL� ��߻�L�������#����t�6�-�b�#۷Q��VF��@�:I�c~��,�ٓ����j�$��n�"	���x ���z�ؔ�C�T��|H���ǻ t�L�bZ�'�OL�A>��f,��~�~���A{��af��$j���^)w^)k�x��O���yA�Jo~�[�Y�6פ�XYƳ�����r���4]�*��{��>#�����/��o�$k�`�H�ߠ@*8t���g��������bōU"��&��Q��f<7�x��ȼܵ\�F�u�8�X0���7�w�	�Z��%�9,��ͼ��4̶\�� 4�A��U♻�	$����1\*�s��ͯ�	��W��v&&ؾ��7�=[�U��-���Y͆	$w^�xϐD�V�ev�fݷ%�;�۳NIg.ᜤ���B��y�b,��iڹ�vN�+�yyE���y��_5
2�1m�d��'n� �o<Aޝx1]�RΊރS�-��$�n������&v	�D�k��N��i�u4�^=w���=ϱ ��q�����(���{\Ҋ%ܳ1-2��#�<�&��O Y���c{R���0�����>f35�˵Sm�\�*�s/6n�U��4�ְ���קn�C�J���5�[]x�����D�~�<@#����}4J�W�t/� �ӯ=�^�R(�v,X�~k�$>59�1`A�~x ���A���7�_]6i�3<w��I������Dd��?H ˹�,���v�O�v�D{�ڇ���_?���j������s	����w;�)벐r��]��W�RȚRaa�k}~��}�u��`w{Z" ڛ�y"F6�=��e�T��0�w�ۭ����H��W?�ąD�ۂ��y$���5ߏdC�& b��2�٬�AV���٪V�[C�{��Ιq~�=�a�?���fb�nI�Ԉr��Mƫ	�\�0�Szރ7�X�(�7Ă��;ܿC^f���W�䤐�30N���L�
\�W�Ve�1(�f��*�s��tG��|�1���\ ��}yvLmt5ύ��p �?s�$2zF$c(c���/������(��-o4r�AðdK@��;�I��r�2�hg�� 1�A$�}�H���M�`f�utѩQT�a���F��jɒ���#�zE���йv���6��݊]�.�B'�xy�"~���y*"�	@d�c�����m�W>�Ԋ,��k|l�~���	�Q��V	諈"_�L���ugU�V�) 0J�`�;;3:f#CfV+�p�k�w-\�[b�5��b�$���߿��,��D@�����<nu�� �Ge�@1�#v��Rg�j�|S�D�|5�����[v3�� ��d`Uh�;ʭQ��j���O䀦�� �Ǐa���qj��!�_�L��f��ˆ�Ay)����kw�k�ѫ�L�?��&�ވ�7������"O3�]f$�~��`�y� �;3"$wm]R~�Ei����`��F$o� TR.�"Z�=t��z����	\�`���̈́o��|{݊�᫤5����,7�����Ol}���0ɯM,�ׂݘq��ե�z3ׯ�aOo��GGwu[�����~�-��M@RH6�#�t�����y�4��5��[��7S�u[4�e�� �)g�+�mq��y��L6g���{;\:�[I^�h��`����w)�Aف� ��n���!s���q'����^�u�y��!g�8p/�99J���9�vʩ�fp�G��vv<���l]a�Z[�dZ�aqol6˒��m����۬gH��mc�L]��u�m�Wfe\��d͗2�uf���6aZW@�u(Ds���~���S'L���э�&w1����'��"��f5��%t�@�|�����zo��dC9.��8a�`A;��XV]43\�K�5�N5�@$gTz=&6�p�t������8X�Y��,�z���1�d�A!�zS�bK=��F�tzy�xPf�E�;�w�@��|�Qon�0����x$jD��D�D������1*��F[z :^�~���������7;+_Z��5h�mU	'ֻ�$@ �1��)���A�`��@-�����*SJ�BV�)ʵZ]��Ѯ�GrΉ��yiN�;1H�r�����y�{1I�>��^%r���[Nn�H3�'��~��:L��E��� *��O߿��Xg�ckvBi�f�(8B8\fB�0�2�����[-܆`�s�~�����`�!�����Oކbs��!�Y�	�������v!�?\'�[�mݐ!�����:r��m���"(c�.u�t:��$�g�|D�����}��-�E��"�@��11�On���kh���I7t�Dx�g;٧��~ٻp���ɧ�x뽒Y�ő'[c�|P+���j��$���k��� ���� ��R����
3F��(�I�r��,�=��� Y܎��i]�=IZ�ݔʬ-��űv��߻��p\;�S��k�|k%���ۜ��M��U��4��<g\O���`7��ݠuNt�E�A���!��I�О�6lN�� �A���`^s�^B<�M��Ή�y)�/J�W<��)�&a.�ގpo��ڈ���{�UP�{���MP��?]Se���Q	�D#&N��BH�q���]zG!����{���}�������
��n�wzgb5Q<��yT��x����H�@���{PLŎif�acZ�ȜďF5����Ӑ�a���4L�����i����>�X��Y�'�Ǥ�縼������A��:ͮl-=��F�p�qI4>K+B�����d�=��-��LX��4�y&�1s�4�9>����	p\M���!>����.��v����y�شa��l�׷ӽ���O��x{�2��cfI��fˉ{�ն���.t{�	��[܌�}u�{:��|f�u?wbl�C�X�_Y��/zv�{�!��z��spǔHn2DX��o}���	�	�ٯ��Rx�w�|�9;� ){ ����V��#Cp���_��+�_{��M�{ݷF�g�7|ݾγ_i����y�"���߮]�\�9��㟷���w�K.�^Еw��x��ڐ��e5��eҠ;\���4^��ot�q���������>㥯�|����V/o�~�%o}������k��vu}��	�b�o�8�[&�uh�7��L��ɬ��nq���ɽ��}�w���r�3�O�>�y��?i�}���s>�B�{݉"�s�����]&[x�	�*r�e�>M^8E� >kxG�j�k[�K��^s�U+�Ͷ�~m�����JQsR�pZzJ�ŹƽM��Ƽj���m.�1[�K� ߜ�+o�V�)O��Z�3���ҽJP<�v���"R�R�$d��(�BIH5iQTR4Dc�!��~��3���}�?�OOOOOM�*Ǖ}���$�c<#�rI���#5�@(����⨚�8Ug���~>3=?��]�v�۷k�H�NH�!"Gǣp ��"��7��Z{8ڭ#GqA*!'ӯ���fq�>�o���������U)�<f"jK����#�)�xĆU����D �wEg@��pRVڧ 
rD~��b �4"�$���0VH���yH3���b�a'�G���LD9� �p�����@���E��%HB��XN���$JZ�D�dQ��r��ңKB6�^8!QB��=��NJZZbDQDEQ#Qx��8�"�@�
Ƒ B*��'@A� g*qF�"% T�2�XD��=��Ҵ%���ʇٞ�bU������}��Fl���wg� �:r�ӻ�%�3��!�������'Ɵ9�I&�6+�H�:{bku��[����k�������	&wp���� �@�Ǯ���b��mx�͌���{A ��;�n�y�X��I�h�De�uͶ�
#���H[Xؖ+�L(5͍�YSb��"H��%�|Y�.�h����x$�;�x�*�O��:j @$��� u��"��w.AMRxk���z=�j:���I5����V����s�A��$4im�Q�D�Ed�Rp��R-3\�M2	$����Ȧ����X�4��� o��5����^S����/��N�&(� ��vm"��lS�l�MK�o$A�|�Fw=���y,Z\4Ū��� ���MY��N{I����)]�=2L~{n]<����3|��{��kӷ3׺=��G�݆u��~�!�Z�h)��_|����[���+F�Ǧ~�!�e����k@�U�g�jD�?DA�q9�ԣ������c�q"��3,�p�W#f�����n��%�jɷc��u��5=tw2�j���	&wtCݭ��k�r��(D�K��փ1��4�����Ay79�6�Q,��[��c�>�V���xB�&^	��^3Qν�s�҂�S����i=��x�A9S}H�vvd�j�h��M�$_<`)]F��5����uР����'H��W?:۔*�^���Ȃ	��Y
'k��D�*��3�OD�E���x�N�
rHZ�����l���hڬ��ى}�z��G����P	��x�`�a��E���5����3��!����Q�����+;�!���yD�$#�JC��e!K��ᧂ�II��@�/�Da��`W��0�,�rh���ǜ�e�# ���JH��!��<a�O	�i	z�"�R���7MƆa�۰��<�=6��P�z3���uu���������9�zzZn#I��mu)k���`Q�hS�U��in��r�Ap�l�����G��{Z2��/TM��x��yUѷW.rk\����-���W#K4bh;9Rh��5b$u·M���&� ii�X�W��6�ʈ�	�q�M+]�ߗh��~}��&tt�����~�� 0/#���P�j$�U��|Osd(%��BgwE�U��������q"㶣�I$^5I=[����^q�-۷w��y@�g�pΝ�@��!C=�b�/*��Iy0��+n�3`	��\(�o��0�~�i�X��߆��ᚔ�dV�'� 1� �_=z����p�3��L�z�����R;�!N�"�$�d3�D	3Ӱ"=qlҨ��e�1q�fsc\�C�E�dG�wM�_cJ��F"u�i��v�[lt�[��MPB��\��>�[uw�v`��`����y'p�	�A��]���ǂ��1 �~y��KN(�9䈾ވ��u��bg@�N��U�a��	ܪf���69�I��˶cJ�Nv���)����Y=˪=��	f@	{��;�c���W]�CO�
�V�(`�V�|<�/�u�】�oD�A����$�3#YRs/��b^]>C�L��*{��� Aȫ�M�q��ko<X��D($�w�2�!��F��fk�.�34�=)��u�[x�T��9��q¬���2	�g��х�W�3���3��30vv,�h\D"�����Lm��}Ɩ8%� �NDH�����B���S6�N��������K4���e�5]���rn&��;b�l�Cu�č�౮�C�ߐ�e��#_ߥݱ�|f;`A��;[�@7�zn(���)Y���$�f.��NM$��@�
�ںa�f��Lztd�Vm-���@o����W�'��TB��2`,�-*��%����iN�')���.���OZ�P	 �_c��36&�̲w.�t�$m��
7E3�=g��#���Y��Y�T0�k���,_�fM�AN��*)��0DתM�F�2LR�x{��H�ˏ2�]*A,�;^@�L��*$��٨1��M7VI=�� ������A;}�~](¶�N|(a|�x���́�N:fhE{�) f��<gD�Y|Ǹ�4Dd��W�E-�h� ���Y`���1���᎒(�.S3��5s֎&;q�u��ᕝ���0g>��r���}����RV	ۤY�v�����D�T�-VZ� �rކ;���+��e�<tDOv��j�E�A�R��, �}�.R�1}v#:4L�rY�%�J�Ҽ#Ƿ1��ϒ ��N�d���f|�D�>�5���$���Kt�5�t�p�����x�ǘq ��Q�y#�v�"	lW?���U.����o��Ez��^��ɣ�b��+�F�_����|]�y.YYY��{��e�w�X��ͩ����`E�쪬��=H�r{8�]Y�H����s�����n�-�@�͉�� ����5n��\�۬H�s�� �Z�I �ODc��*���1(�g�/�L�4�;9	��6af���Q��9u'�sŜvR��y�wg١�@t��&f���ӭ ��ׁ>H�u��
���+U\k��	9}� ��;,C��wA;H><����(k�Y�5�W(�|	�%��Ajz ��0*��j��w\�$D���bU��E2�]���	񮋈-�++��]�ʅ�����+�{���4s��Q�x��[�+��۬X���/6� ����>^�n�B�����	�M�ă�yn�������� ��j���Pl�x�o~�>��㽰���h001�j�s�S- �2ɓ�XE\94�͍�/O.�Db]����M�?o{��/��g�N.����A։P�a���-�7�;��OYN��@1�1?��`8��w͋/Lr�1׶��+";є�	I1x���"��=\i�ӹ����sO\۲ey��U�,;K��a�V����va�%puk��rG�\���=�ն�O[W��a��Qw���{`�=D�㧂�Zۓ��U�s˸��K��#��Ƿ4��Au75r�&�ã\�r���	U�u�j+��]��<p���˺��{se���[V���4nBC�;<ѳ�^j���Εςjv����߾��k�����}��C|Ù�n`�j0lb�0�GL }h;��A��>I�����t��&f�&�w��i��7Bml��骴�`�H�˨	����H�b���[��绅m"݋�	�E��$k��<|�6�Ns�z�Mݽ@�[�m�Tzs���3� �`l1!�N�U;GF;_�cH����Y�� A��y0޾|�bvV���v�O2�7�$�3��-2
�i;��o�/��Ǣ�gP����5�q>� �ט>�!:�z��^���b���P��D�8��[F5u��Ȭݳ=�{t���r���}���6I�(��ӛ�}���^	$������� 6����I�'�I��'QfNK"�UȘ�o��|:8�6��f��cɅ�����fX)(���7�Y^����E�X���x�e�Ʌ*�4�Ⱥ�b��VyY�ʷ�o����m�$�f� C�!K�k�#�@�	LV��cn��8���ڗ.�t��feK��$�5��H�%�i�L����������<O��N�!��;���A�ѳ��h��D�_��	�n�D�A�y5���C.
YE�6�	�w�!y!�-�^d�� ��؊����0���rZ*\@$��ȃ�H��o-���w����K���.���4.�i�¬1�nG�3^��6�.���"9��￿!	���@/��
���A�q�A �踏�������� @$��n2�1D�Hp���%������\V�x��"�v�\�{n�<���E�ͭ��8�2rYz����I �E�RDzV�Cٷ$GmDM����/[���*�j4����>yg��vŌo&ȅ���7���^��^}��2�C ����rÇ��i� |2��� ���������Y	#tm��sS���������	���#5��a��m������w#�EYA��;���A����H�����s*���w� �Ol�r��� ���w�6�0��&�ؒ<7�t�烘��^�\�m˛e�#	��T���������`K��̃�o� 	3S���� ��Y]�.4�u=OU��Y8$�
��~�q h�ܡ�y�UμwG8�A�R5\��-�٠�]��.Q.�$Oz���  ?��-�ĀW���h��3�d٢/����:::��"I�̜�I@��ﵪ�M�E���$�俠��dl����]��X�3a���QM��96f�ɒ�*=L΃�����^԰��n���ͣ|�t�hރUNu�����w�wY��YO����DNwzd�k�r����fS ����@���_g���L����6���!��!��7Q��o��T���w�O�~�=�W�5�)��l�v�,�v�-�j��3�xys���:M��T�u��}_�zgV�7P�	�I�H��q��>�����9#m+PS���o躁 �v�c��܃�0�X��3�a�:��v�:�E[Tt+�>^�l�A��x _�s�ͥ���v={:��e&r��%��z��A=ۯ�H���B�������� ?����A-�Xo\�8N�M�K��Zf�1�:tp�O�	7��`U���;�v;K�����7�%�c��AN��I)�f�Dx��zm+�mB*�F6 IY� 	��"=������Z	��:�=�T��B��%�ۛ������0nx����1�.xC�e+�}���[��[�!Kw9xi|�Ź콺��VN���ș���n2��
��9��>�}�5M9VB�#�{M��v�}ٯyz�;x��_D\ن��m� ��y>P$���T��l�|^�wފ=��Aܫj�U�~����P<����.;Z��W�e�5�r���f~�����"E��3�Ga�>]����w��Kp�&l�ޕ|`	f�%���C���3���ׯ�i�{�i\G mj<�j�S`�Rr�Ig�cf>L��Y����w�O���u�K=���/�"����4{.� ����a�e����V��3�CY�.D������%�q�����7�Q�I�S�&������5}�K|�X ��.Fq�`; 5��^Fh��]��Q�{ר`��n�%\3�|��Vw��h��}�9r���[��������w�F�ۜr꽓�J�S��9�k��Dρ9�����z]��݈@����7=��5�=n�{{���}��ὍBY�Zxw��7���y�-�zy�=<7nh�R�g���ݻ��y<��.�����s��c�}��y��Ǔ���t�����ކd{1B��8�W���S����jO=�����^�rҭ��G#Тs�X=9�Y����O>���q@Q�G�����G�M�e�o{���������=�,˩璂�kJ�m�:�_cȆND3�*.PG�U@L`u�Y	�Ԧ�>�f	3��գ���-B���ҷ'&��T�Z�gǼ�#2"��r8�\���?N�8��}�?{�nݻv�4&�$"�,@H�T0�� /��&�;<đ9�rZ)��
�����~38�+u���VVVVV��E9v�&IPQF�\�1'|xE\��IÉ�(�ɹ˜b���~>38��+���YYYYYW�� �(�*��p|Y
1bpB*"K*C��AZV�Mj�f�;���Q�H���ט@�� qX8Hd�'Aq%�,NAB<�<�B��@qm�RF�^B"�䕤�qY�� t�T��@�BE`$xA���m$�)��u�p� �D�F+	匤"�H�/2��HBB	ѐ�a!�E� ���H� 8%cABp@�+m�#�[)a ��'�$�  H�
��/JDO��Eg)ޣ�C��x���EiGp���F2��r�K7'��vz���m�[n��;M�N�c�����*�J�MW9��I��˞�rM�.u�u�l�\�O<`�q�M�=s����vxK���ӽ.޶���q��Zn�=1�qvť�E�Hi �)&�	a�-\�����r\^W[��\�2�L�c�+r����B��l��v��aa�3���8�p�ˮ����svv$G��/]���p��qf�,�,	M4r�6�e��&%��`��B�[��v�NNdH�z�(�p��m��W�ܛS�Z��Mt^��N�D�۶��N���^:�б�=
���j��X��j�j���;��2��Q��y�nzz��#ܓk-�v����(�G�e��q�x:D5q�8z�>lM�[
J��^l5�n���-�m���BG���;]�<5#�VŇ7w#7t�c�tQ��ݎ��u���s����aCiua�+���su��@�1���ь��d&���u�L�e��6��%�z���v��nP1T<b�۫�Ǘ+�$��u�Sj�"���*	�1�Xʥ]�������\�`�`9�Յݡ��t�^#����`��3Dm�9Ğ��t�Xkt��D���� ܋�9�7)�p
�(g���6]�LŪk2�^ր�kx��7���cD��}�E�]mC�El#����T"BhKZV9!��=�6p\Ӷ^n)h�)����W���˸��)�RؽVV�X�*FŅ�UÚ�h���H'�<Τzr�[-�יXZ˦)e���q��cRi�^����J��pnv���-�^Sq����c���ۛ�NíU�������S(e礑N�Օ���|�n.+��.w`Ńc3@�Mcb�{�� ��GY�����V��D�m���a�����W���v�WM�u�Af+���g#z�d��,��K.��Hk���K��-V�]��s���ʀ+��e��+aKaֽ��p��i��I�����V����!�\qj�A�ⳮN3h��y�7m^�Q�*^s�6��j��6�`�hl0+kã�c�[�!3�=K�=�k����m��Iz61
�u�bM�U�kð����8ͱs�q����{s�r.Y8�qrr��n�Bo%c�]WA�2ʼME��i�E�VE�\ݵ��֛p�,�PƁ,���ś+�eгGd��CP���,Ȃ��e�Ͷ���]��$}���htw@���>O/F%5���Q1�h�wvN�'i�h�DDK��V�9�V4�%���͈$�}�	O)�mq�K��PaH��'�T���D���!��F:��T�;͐�G��ވ �M�LA��d�L��)��k�N9�<'�$h�qK�{���2�3�ME�웼9�\�'H�'sN���W����s�_k���O[�<k�"oe�~����]h����tS�o;"�I3:2=���ڹw,�e�q�]�5���iI.��={�>�Ѯ_^��1�=�1���bvy�ǈ���yy9��I���xw�m�LBwpS2�5����vԺ���=��l.fڊ�b��Bv�XÑB�ո`l�|�T7fŝ�ꗖ{�A�4�g��2d�}������0c�G��3�O�|U�%gj"<�`�T�`PюF�o'h�&=�����v�l�k�@�>�� m_Џ���g<.P���s�bALN�>���0�\_��*��D��5=U4Q�x���?���{0I>ξ�L����{|�;�^�:�i"�;��- 7�33i��׸�
h���A��ީ����-dO�n�<x���f�Y��q���8wK۞�������XI�8�K�շl�Y��ɻҝ$�t滯 �rD�j�b	 �KY�I;x-�-V�_"�e{�	������@#g`�JdslDKp�ۯqѭ�k7�A�_B�]��|_�
=���5p�C=��~t�gd���;8�Iz��A��!�>B�)��&�?^Pck]�É�_��y��l��)�n5�<���ʆ?��Fg�eAM���m��9"��j��=:��C0>$h�o�$�u��@'ٷ���u�N�Ӻ	�d�"��[I�K�sBM�	���D	�݁^#WD�J�w���`;60��pA:�T�DA �Θ)p��.�����$M����C��x�Θ���=�=GfK[�N�$���L��I��9�tf�v^�V-�L��d����3���^���8�k��I��x ������G0��Wosż��ȀN���wo �rD�QZ������N{�E��Ty��WDI�彔�� -g���8_��<O ����J$ktD깈>$G����2gq�>���"|@ NgDI��ɏEV����Y��fS ��֕�O���Lu�.�K�[���x���������	^x�-3P]m�٦w���'8�ӏ�Зٞ�
�\���*B�8�����q�>^x����Nq1`K38< �x�����f�mc)��߇��'cy(W�$v�@�D�����q����5+ӧ�� ~>�s�F�q z.����-�%q��v3����ܹk�義g����%w��tA 
ޗ�A͇��:��x�ר�ӑ��A� ˮ�˟X4��� �������5rh튫y ��Uy|��ݗ��TnK�9ï�I�:���:.�2V��z#�������,k��TtI��z6hgWD�����Gw`̊�X���}D��Y	&M�O�A��:����X�v��!�dg����ڟd3�L�d�k��I�ھx�:��+�Dg'$�׀���ѭ ��u����X_)gP��SF�MU"�{Ӡ�{f�'�cb�{zc�׎K~ZL	����>����r�}�9\\CD��󵚚�q
kA��J D�v�������|�y?t�|�,��
�[�;��q���˶ɼ��yg`nu/���fK�2[����v}&9��v8�[�!;�;<�v56�u�]2]�D�md�9����#p.�F��Ws;������sco#m<6��rBۭ���-��ñ�:ݽb���vA��v_��a��eG�l�FJ�:f)]8̫6��[?�<�U�%�U��x���֝�5��7m㋮#5"l�ňa�������зu��A���4Ih�a�~���N����f�@_x�� �=8�	�*�w�p���J��H�_� Cz���L��	�$0��')[�'~�!�4���v��"�"yd�@'�א�n��:Iř�����D�z������(�t�ٻ��A���u��a6��r�ƀk�#��O����������� �vU�)��+�˘�� �w��@t7�P'L�b�$r��7\lĻ�,ȨA��b=��*�����-x�6����n����#������L;v�n����-L4��k\�+�����t�M�3�2��0JM�`�������U��~��Yٸ�D��A>=�n;p�ts��ia7n�� /_�<g`p)ݝ9t��H-�-�a�&|m�FT�jk�I�S<���9�$߈ �u�WEw�{H�;!�mg,�]��"���I�Ӻ�ѧ�� �xQ�qJ�y�ގ� ����
��)]���	���CY)ܱ(;]�>DuF��F��sL��x�z��k���`���E�T3��`K@%���Ȯ̰g� ޞ�+�x�7��#�i���B�h�4)��2�p#���^��$L���q��5����[�����z ���� H��� ���������ޚ�S/gj�Z��K�0�Wh�贆�T;c��7M��о�~?�?Gk�ĨL���ٸ�?�8z9�w���f-E>�-9�}~^�T=a �w^]�d�Ɍ�p��y���w7z��5�I ��}	'�G_�A���Ϲ��E�m:�)ݝ9t��A�]��#�x������l�:_fQ�@�z���Ŷ̄��d`�n����{t.(���{���T:U>����ui�n��H��g[Yu������y#���9��������-�#z�	�pĠ�M�<tc��I��DWeǠ�
V��@$o_G;J0��^�z���q]��J�r�L	h@�h�rI={� ��*���$K�DA>��-��}V>K	9����<��Z�-�R�\-�n�v.�VۓV��T!VkΏS[a�{�����3W@=����)-9����	!щ�2;�6V"����G��0���1�p'vvf@��1 �u��P�j&lͽA$�Y��I��� HRzv��]�63z����]��L����9$��Aoq���خ��jΦ�~Pٹ� �{1��ݝ$�-䎳���7����@1 9�$���A ���y��OU� )�b�ʘ-���S\õ'�قʰr�Xx]v��sߤ���r6a4cf~�^�< ��/e��K๘��J\��3���BR�(�h&�dNJgJ�|�s��3�06�U9s|经�J���M�I ���,ϗ9H*�J9)�'\�-��Du���lk����Z�l�Xs���+=�$�Ž#�w'����-(�����4*�N��qN�z�kX���w��g(c�A�d䉟Θ�7O<�5l���N,M��5Y� ��=�M���,��Q�̷d�[ۭ~&��r�׉�����K]�l���v�$���-M� �����$_L 6�Ȱ]��L�&P*��1��j�k�2[IM ��s����z�h�[K�jkbC�t}5W\X�8,�]��Dl>�$���������n8�竑 ����:���{��(�y�.U���#8�5�SГ��ܱ3�Zr�"�$Ҧ��|��9&U���e�^�~L.�yj�d	�y|�����# ��:���T�C-܂���u0b-,�
0�8r�u�u��m�k��ՍUP=��ٜ�]f����O��CC�v�q�a�Wv��9�zm���횸\��iF^�Of9	�a��77;v�[ύȎM�@Ѭ
�ɵ�k��@��b+��݌Ke�,)w0�ȶ%>n��#���\���n��;g.�:�4LeP�t�kc���i���ֵc��-ˮ�k�x��	8wnU4c�[��xɲ)�Mc�~gx����Aۖ5?ԃ��n�A�=]1��6�n�t�Dx�r�]�2�Y)���`K@>�!wT@����ٲV;8���NG��r�y/=��H3E�u��lꛀh�(;NH�"w�=�d��@$���Cő"�*[_���>5�'�OJ`x��@/��@��Y�;�7<��j�����$ؗ@�{1�_� ��H"3�m�kI���_d��f���]��	��U�c��7��]��q��O��"  �e4������8�݋Z1Dk4�,�r�$p�\l۫�cv-�n�j�Ԭ%�nWB��#�kev̦����r��㯷�#u��sU��^��zB��<�^D�d�$⻦6�|h;2p�e5��'-m���ؙ�4��{�}���+x
�R�:����2[���uׅ�;��ފ�ф�����tcvl�b��uv��:*��jV�m�7V0ý��w���-�a>27��ݺ������;�{ۙ@$�X)0%@��b��3������d!��:}O�.Z�g��x�U<��H$n�Dx�U����; Lz��:��7�j8a�D�#e��<x�{��'<�7K��	�w}�0W���h�=:d5�;2�L���  �ܻOR���M�H�m ϐY�� �m:̡����TN���^��?�geextЍ�u$Κk�����n��HV�i�u��������ى`��F7���>$�^�x�N�L7�&7!��ȋ�]�$��Dx����qwfp��-� ��OʆP�a9�~p�5���قI;�0q���v�%���j͟̜8,@�ȍ��>Ă�fTA�'@�8AS^�֙m��zv��z$�쏁����UᢕN�z�7<z�Ct�f����jݱz���O�qG(�}��gӮë���zE]Ѝ�v=�e����׶�傅�n@��Cc?��yw�4�&~"?nض���,��3��4���^�#����vhɜ�B&L�H��"R��^���W������ރ�2X���@��Q�b��֯��w'���{k��{�B����\���W����E��Xў��cU��Gom��l�;�x�g�������}�Y%�`�Ll���ݜ\���t5n�~���C(��[�'2^��p��y��G��#�ڇ��Z��W<zNGS�o����L��~�	���S75�����`#oY{�"�b��aW�}}�sچ#�>�r����j	��S�-��5�!o��]��7�H~�(�ݘ�)�':����I�͊��5OXw�+�఼��L��.��sK�:��c��ɊQ�!���𗳷���绦L}ݐ�4���.ܩvݾ��.��Q��;8��c�#�S"�Q)�+Wu�L�6�jVM��u�e廹"���5�@�ra��8:g�U�4W��>����bc��ޞ���};����{�_oU�����:��e����w'���\g�UU���$�Woggc��[4"����L�bP��M�Ф�gm���L��,ofD.���3����9���l��.V�v�H�i�2
�$TQ��r%_�JW#J"�-[Pj���UE��~<g��z~���ǧ����0@
O���+��#��H�B1�$%*�Q#"up(��\�������~ǧ��>>:��VVVVV`��8�0��䑌b@ #�P@�&�M(�1�I$�4����5�J�뎾����������̛�+��5Ĩ�Q-#Pc)5h � ���I�Ocr�X$AXr$��8�"�����Ē��UJEE�Qh�j�4�@0�,N���1NN'�=����`��Q��@(��� M�Ʈ�+l�X��H���D[�d"�ҭ ��$�yK`B�c"N+ʧ�[16��JQ�0E+!AQEjB5lPE*%��i%DE�������("[�5.R���5p�53��8�F@���8$`��������.�Pۮ����_nDs�.Χ���(1�ኈ���9��9;Y�9����*�bvy�.�����|�����'<�S&L��U�/�$x������,T�Z^�@���[\���|{ן��Z�~��
K1L�#i��)��X[��8n��A6�&|�����טp5�;2�g��^�$Ud�{��:z�=]� ζx�q�뗏?�oN��0`��F ��o2��]42�,�xc���F��& ��3 �t7����W'��qy�M��dk�g3E��[3�*��G; 8^I颵�B�]5s�I�/fI���:��h:d�â�dw�l�1SW>H�@�O����a$f�A������'s�t��T���_�:3�?ñz��s�ߐ�a�{�Պ欃��ް6wC�Wj�Yu������mP�����L�5�kL;�z	9������)��ኆ��<��ۏ �<�X�޼'ɻ�G���~h�#;9��*%�nh�\��$�RE�.���J����u�6�q�wk[�6qp�A��d݇��'�����/���xq���$�gD NUʧ�ݾ�q�x� ����G�׷��:];�0t�M.,�~���Y�>`��is�y俔��l�A
�-0G-B�o;+�ד��fĦ�4��$u�<I�������Z�$⫆�vtE�;�w�9�3�����!yY�x�B�O"&�h�eU$�|\�s@$��؂L�-�y�;
�]ڙ��O��u�l;2p��c@k5=��L�lCE�
욀G[��>5�����՚q���h4�	�!�.T�Ю���Ӊ�vI�~>�sԍ���*4E�/�F��w�����C�pj��om(��Ƿ��G����n�����-�[�t���眥���2�m�M4�*�L%ͰۊWv]�\����;�b�k[��nhյ�W�9�n5�s��!���!��t��tsZ��hP�9�y��`�u^���p��*kDV�ŧ:$����m�&�h��i9ֹ���i��q���M&B�f9�tt��logM�e�5�pO:LT��Pv�6�c�L�kq�G��	4���n�*Ÿ�nvu�aC�C�3l�]�[��{ڹ.VK��q�����L��� 	ё�j�Ի�����Ǌ��WwD�Oe���L���$إ�ǚ�ut�c̾�� �n���'�� yQ���[*��g6ă�:t���xM�P �r���r8-0�Y��o�� ��ȃ~H��={�s�f�����[F���- �J���/G� ��<�5���� �D�����:-|q�"+ʼ����2�s�|���k����$��ȇ�y1 �<8��E��Y ��	�����Zqk��g�r��;4Ϝ/f:�g7	�'Gu��:J'��ٝ��	�sc�@$��
I��v�<��j�����/�" W�'.<ə�A��z"{�eS�旦i�IlSiv�Ol,�u�Bmu�
�xj�7o$eP��%I�Bd�wp�[	��8����}�ӤA���^F��ˇ���
��x��|��c���$wu��	�b�Y]�M��=d;d���c�c �8�\8^J����e��mz} �yw`�%���@��A�z�l���&t���1�&�g�HH�/G�B��BS���E7l5�1*f��x�\D��E��ft���ţ`9-�v��5@��(uAoJ�	Uw	�e���: 1�,@@�}�4�i5GL�vɋm�ei�/��������s���w%̃�.p�7�7-��9����>[�_��u�ެ4E��ꀀI�e���(wm���3�p�@�{��e�v�� ���+�/bͶbޅ^�\�	5{m��5Uّ�}�W-��ɐ�̓w^�lP~�=�UߕY�V�8m�Kv{/%VcK˫MNQ��RM[�G��1E&��S�CN����T���.�#�~�7��oKx�[���R��˹h�x|�H�wl#č��H��',�d�0w@�OL��y���w���g�iy�p|O��b�?� ���l����%�d0�W�7�8wp���.��^/��3�H�e���DC��`X�^�W�Ăsw�oG�0��y��I5��5����Ld��k	��8��.��Dm��mjPq1u�é�c�ԝ��}�@//l�.��r����/=(!��;�^kg�h�0��I�[ɶn;'��L��=��.����/F�Y�Hܾ� � ����Ay���O4���"a�������읋�b�؋���$=����f�7O�D��G ��oF�H�5ٞd�69�L���
����cY6�@1/o H�-旿<�����r ��z�!��N��29y�b���P��p�Sp÷�{cJm?k
�O�a�+����{y�J��ή��=�T^�<N��\�f�z�<n�ޏ	��,{rI�x��=�^� ���XT<mS��>��G��M��#t�;�v�8�Ꞹ���#�.� �q��xf�0�=�OG�ay�d3���sZ �|v�`A�t�M�h*�<�^=m\}	�ٻVIf	2.�Ёvx�CAS���/2���O��>틈 �[����fB��>���;�i5��Os�r��������>��4\�[��N��E;'b�8a�7>�����o`��(�Y���H��茞��}��V���|���1LB�!����	�Ǟ[A���v7�,��5�=�;�o�Z��	����u�F�M�M���	҄�Axz�^xorz�;��������H��B�{�)����[UՌ�R=����[��ZL�����y=y[��TR��-��qHcFy,w2v]�g��H��Om���efZ�Y�H�:W��,���mjƻ;t�V��ת�니^�nu�o��q�1�m�;U�VR�A�EQ�F�B�] e�*.��)��&�0h��<�;��kn�x���v�RjU���u�5��wbk��^‭";��z�&�3v倣�vN��F+����&*q�x��Uh��Kvn�kv̝\g8���熧%�sr�W2�0q&�%��G���vce�s$���f�#NdG�/ ���A�OYl4�r&	��Ifݏ@!y!��?�hP8��w:7͵	.8ص�X����Ɖ���}�}H)E�۫�l����Gyv͐Y�f�: �w��k�W?8�x�[��+S�e}�	�W��gL���\��tK�{����VA2�c���_�x�|��f$��E�~=p�p���@��U�H�]�Iٝ�8NT��s�yO��3�#���b�Q8���M��O�_�D�T���ۻ{�i�F�p�
`��!�Mu�+�%��z�m�]TZ�#c�m;c!
���I���2S����n�A���|xߐ�y,�st���"�h�;H7��i� [�{l´�0,�!��F�o��a�:�К����G�i��7d�J%1�A������"l��W =D�&Cĉ�=���\�B�ka�+���2�q�t��u2�ϒ"�" �N��z�/�;&v1�vDc{��\;��[��a��;y �l��m���������	��6 �u�z�ز��A�3��"�[�Y��N����*�%�C�DA �ޖ�~��}e[{���VMG�4&@j�]'�|�42�sܥ}�����#n|@��9��֣v�&x�g��3[ 5c��B;K[(�V�Lhl��n�j0ڨ���,�>~��;�p��n�+��: ��@� ?8��op+��@=�� ���aT�;((^,w�<��SB�����6��dtA �bHD�R`P}%t:���&�ڢ�	�/` ��1I��C�H9�!J��1��ީ�A�D#�>i�3G�NW.�[�4#���@ԨA��p�ʍ��	���hu5��K���8E5�w�����ף������z;�/�ē��A�G����b�3V��Z;�f<�����o�v�K��l�W-��	+��$^ux�,��a���Y�}����aH-�Wo��H�̏q�v����{;:$�����y������DQU$sQ�L0��
ʳ0�p�vrR��%��ˡ��%r2���!�V�C�pΉv�����I �͈rO��3Ӻ���%�������)[��UȤ���ӆN���A Ʊ����K��{]��'�-Y҃A ��ȂN٪ʫ�yǋ��:��!��()��tǜ���_3�j=�Yu�����$�ˆ��^$w?D��nY�1ً8c�Ǫzn�4��i������ �w/�@$�3�o���{���e�X�8*����6��)��a@�z�t?�#�w���S��N���c�)�;�[���.���J4�b��J�Z#�{3եᜐ�4��4�� g���5�{��N�>�y��H�݈PD�M����l?>������ݴ�llGM�����̓s��׬�z�-�n,&�f��[n�����e�vY��f^	3]��$;� <��7"����@��H
�F2��\3�SǗc؅���h�ު3��rH;w���;ϑ��3�H��v��ɍ���H�u��׃�e��^� ���I ��� �$o	vxf��S�����Aw�� �N��4�d���
A:���l�QZOm��jc�	�ɷ	��lq�_@�F6�+�b8��{����	�h6^�	<q�<��2�_D��Y<��o'b=�ι���?��s���8��*�����Q�|�����H (�?�z  ����:83� y
�41 !(H CCC(�C"�0C� @�ȫ2��0��� CL�2L �L��C"��Ax!*�$!���=`� ��(qEL������`�*���z�!���"$! 	J*B
��
�! �H�B����8�pBR�T�$� �G!� U�!�!�$�!U�Qa	aEa	a	aEaEaa�x!�H+B�J+B+J+@�J+B+@ B�����40��*�*��0*�
� 42
���������*�40*�*������+0��B B*��
�������� 4 !"�1(C C�4��!(�! @ CCC"�!���!*H� J��;���pp�~��DfT��?��Ϗ������� ���T������������������o����O��'�����������(�������O�Q��QEb�/��D����������?��
����������'>��4������o@s�� ���\+���DEX$��Ve!�TY!��YIQe�VXdd��@�VREYdU�Eed�!��VAY%��VVXIQ`	da�%�TXYe ���� B � $	XB��!	P%$I%d$	!	� ��BXY�!�"���
"D���h� A
���EhR��EiEbDV� ��EbV U�QZX�V�V$�AV!�Ea�VHe�Va��V!U�`�V�VdU�d�V!�AXrpx�+ �H��?xp�?����O�UDiU�
���@�������AA����@����9�*�������O��g�?����8� ���?��'G�������؟�㟄� ���*�+��~�?��PAE��~Þ�@E}���I��^��p/x�!���>����`�*�+~H�����*�+����=~�[���O�:���>�O�������UE��?�?���(���a��AI�_�p�p=���q��M� ��x{��EQE{OA>���q�@~��������&�_�AE�L���^_�����o�?xq�?�1AY&SY'ѵ��DY�`P��3'� b_= 
)C���4@V�m��ٶ��J[E(�(6�� ��HF� 
5��6� ��P  ;�(<�TH""T����
UB�T"�
�TH�TIQ**T������EU*A)$�J�¢�HUP%U!*K�                                     >        � �6���ͧ6[U�;WH5u�j�E��J"� ���r�6�n���uݪ��M!p ;]��u�56��n���Z����  �y�����V۝�v�M�s�7]�K�{N�����
x��`+�h��� �  `粏B��4��a�@�� �=
����  }@        >( ̓�h���g@^�@y��`��� �EcW� �s��s@<��A��4th�o �w������S��v5("U4��� >租c�����
�e� �:Cu�׶vͼ�v��Լ��ɫg6Uvթ� .\�&�o]Ս�Թ����w\�T�wy�B�4�D� B�|��    >�    �J��ݻcY�e�wݸ޲魏v�;����z W��9ڸm�m�s�ܧ�^�V����-. r����ܨ����1$�*T
�/�  .C��U:�sn�%� �.�5�nϹӫy�v�۹�ZN�km��f���V��;v��m�家�Un��0����F�R�H���  =�      ( =K�knf�4�\�t_v��f�����[i�t .�3Zsep���5+���[�[Ykn���Fp���[n��jf���6j*G�  {����Եl�:�jÀ��m��i�V���U��Uv[UӮT�f� ��f�7v�[R�;��Mm�]٭�c��Z��R*J�RU�  �        p��-�Y[��J���v��7r��n
�s��li��Q%w3��6sn�� ݭ��7$�9"J�*��� ^�С9ع�[�j���n��[��DKt��[mٹ��N wUJ��ʻS���#W7R�b�`\� 5O�JR�  E?#)J� h�ʩSƩ%  !��?h����   ��JJ�i�14`��ML�)!@G�w��?��������UZ��?�G���L���$�	/ Z�� I[HB!#�@�$����%�P$�	&��BG���������&��ۭ�[_^����/�bef�ěYJCdwa<���%Y�'���P�ۖ7"��+jwtQĆ]�9�J�qS�����j�[r���o�2I��n�J���ձԍ�V݇2�A�ӗ2��w�Y6kjF#[um�f�s	ݷZ�[��4��F�b��Z����ݨ)�ׯr+voẒ�lx-��XU�b�`�zFS��P��M��#p�%�ݟ �%<ޚ:��C�+s:&]�ԤMFҨ1����]��K�Я��Zwv�+�{.��C6�����v�3�P��9h癄͛�u�̄�	�oWG���X�e��␝A�j���"��eJÁͰ�F�J�%D�.���eKj��2G��
hȅ�jZ\h�y���⦴�����ia%wY�#W1�g1�F��ɛ��G��"�tHg2��t�U�P������X�[�+"�@oE	K+d�����0�i�b�U��:��5��'o*�ss\� �J	c�mZ�fP՚&�o��w]�N�M�Kf
#���j�+	ݢ)\N�N㫥"�ӏ��1��Y˕�����jn�ѐ�'7*g�P�8B��q��@�`6;�����wu��un�<c2��:F!wr���^�L�P�[+f�эd��ڛ�Št�z�՚��Q;aa�"��)���ְ�U��M��{�F"�wq�wB92�&��x�e"���zf݌$cL�Lp-r�d��{���R'f��]Y��L���8lش\nȳ4�;��`�k��+5�32��f;ɢ�b�b�[2���̺¤�(	��K�DV��j�ft�g�D����4�w�&hQU���,�.Q6�V�oDy(-�Or�E��kK�kn�ˋ�LѺ�z,ǈ�9K�-�ڲ�n��.]v��
�=Xw�ں&n@Y��7͒f�����6�m��N�%IC3m�E7�&��{�4��@ҝ��q�3t�lAt�r�#"��lk����RYY2�F�[�UYYwX�mvY�8��ePM���E�%��Qhݠ-^fj�ٱvd#�d��cź��Ѹ��Ձvf��Ʀ���[�kA�I�ɶ��ާv��5���h`-��۩/�(GN-�&�fq�n��yu�Hh̲c��9��7�������c�Nrҭ���L�)�شHRշn�%ɀ�c9:u���^Y�Y�Kٱfl�y)���̭�"պ�nn�B�/h5Ge4V^�Z�,˼8+vu`��Y�����1�e%W�B��� ��8b��+��V������J4��n�"�̦r�a�5i�L���4mEO)����nj��eqz�f��l�[WcBǣ^�k;B�]Yzcɴ�]�.��ѐ֥k5��F٥��,���U�)�FQbޕ4t!���+ȍٺ(i����t]KL��e�ۻϲ�Y��1�U�Ǵ��ue�[q�b
�W�F��ƀѷB�ʖRP�l��]�w	�0���,�mZ7�6�i'Yz�G�)���0��f`�S�r��*�Cw2�.�7t�60c�[N��ʺ�Me]�[�!��hƦ'���u�WQ��v�k�˓j�\okCy����tt�6L�Gp��� ��R�]f���]��f�I۰u��;rr�(Cn@��2�;+G~�L��
� b�{�[Ci��m'>&bg%Չ�����eU�R�y�r�3��a�6D*�4�B���D����6���v�$�o#��UJ�V��vF�Z�����Օ��^��2,o2�Ĭ�I`�j��j^�{-�>i��fft�2�}��N�kD���i����lXhV�;ۋ"ɭ��9n��eݬYu�}K��}���b��P���Y��qe\԰m�)�����޸���Fi�'9w��i�QEvA��z�?�0;����o"���v�FEP���x��NZ�shn^+����b��V]M�6�n��a�����n�'�xr6��̋C���Ŋyb8�h�dn�� ��!�X��Iu0��0��?:r�]*F���8sɹ{|��1n��	��!6�ݓ@[6m`�ڎ'Swo0��n��.���V�iO��v�5�XMoϫ�!F�"�-fMmƑi@��xPV@�5�YhK�ġ�J�3qI$����L	���n���GN�W*%5��.�`E��$T�%1��4�U�t�:��n����I�y�͚���[�f;�q���ӎ���h�k���*��0 +5��4m��A�R�l	��qҲ�/��h�:O�qܲհ�]�[lw��v�ЦEq;4heŒ8����V�i�����c�
���u	�c�J�&����&��vԇn:u��U��O�È�n�u(�E�MAZ�*���/aY-K��c8[w-&�^�̘M�C ܅��V�2��.���1,�0��I�l����7r2�׷��ٮ�R���`����d��V)��ޜ�#b�4�5My�&1�^7&����g��>T�UYUF�!�,�W��0V3��~t7fڛ��x�I��K���f�4 ����Ź(�]DE���cyeVd�7q��U��R6n��òJyx����x\F���1��Ths�oV����yGŃ\�8��H-ʺgv'r��#�e,ϠЅ�,�˴r���r��3rcp]���N���'B��Ocǎ�j�y�����p;�C�*��lڙ���v�`�p�ʡ�㜫*�m]�sS8�r����o
��]�wKl۬�ڷHZu�3�wS�wb�f�z4!�1=��S7�8�˼7�jI��zYƞ��F��tY:5l��xFӣ�3"��F������{!Y�v��" �����M0�ܺ����(���r�is��V]���A��0��V���N̠��7�h�%��S��[�[� Eʲ�l<0�on*4p�+(�< ͂���(�a-���Em# �o��m3Z�X3�T;�w�R�
&��	�5���6�M=��wE�G�f�в���vl�M*���Y[����ʺ:ܲ����<��yL�yJ���ݖ��	�u�ƣ��F�tfѫ"��{�U�gukñP9L{�E�ʱx��
6���lh��i��}�Xwup�sm@��lz�ŅH�Dc!��Uެ�6�ke�����a8�"�kvٌl 
ƞ�̙5g[�K'o�YŦn�pcmk����lJ����u�
ėS,�#�U��	�޳���S�tL;�1QW���0,�1A��"�!�	q3�� �i�����k�������]���ݭ�1����`�[{���eM%=ϥ��4-�pة�C��RY1�Wv$���Ӽ����Ѷ��|C?H�^͂VLof�A��[��-!�óyH��%Y�+r�u�����9,ّ�7���b��[7*��9�@x^4�]����L�ɸ�ԙSq� ��v�2[(�з�WR`�`��a�� 2�!�'E*˳|#�4I4��9l��*���	es\"�{�������wJɌ�1̓.���cZN�8U�U�;�e����o1�\	h�c���*����'Sќ/0Ro�"ݝ$[������x*����#k�,�Ņ�I�yww{N�L��k	;�K��7�ڒ�E!��mb��� t�</^�uW��2֦䰕J�E �ަ/&���?(��3�X���Um]���)봞e:�y0��9�0����j��yW�D)�8Y�/1�h�cI�Y�X`9AИ�s��z	.�A^)�Y�XnS�u�]�����K>���v�9n:��o*����T�A^���N�5�f����M�5.�I���9+�q�F��� Dw�2k��a�c|j��9��UT��][0�[���0=�80�cObUd������F�ܳlZ�nhe]��L5��u;e��y�sU*�����#���ǎ�:�ܶJ�Z����ɩ���ʶv�nj��1ݠ,R��������E�kO7�uVpCVCsV��b��㓆�x���X�٧D���Hg&Pж�x,6��Y@e�HTF���0mH�a:*ֈ���1���۽�gu��63E�7qῥ8�,Fe����eR�^�b��A�z��.��ȼ���j��(�9/]��`Q[ w�n(.��*݇{ӫ'ë�m][���Ԕ��<�Mۼ�xb9r�C�f�a�p��Z����� Wz��NY�0m�ӛ�/re�5EiT�5j�Q�1E�GĲ�ә���`�S)еLf��ģ�i�n�0if�X�Ϭ��l��7�nP� ��+��>������r��L�(V�A�n&�4��r� F:�Mܓ����ɫm)�&b�w�9�\����Ĳ�N\t+%[?����7�5A�E^бt�e��ԭ;�at��>�p��-ۼ4N�R��a٫"g=+lݜ�r����kc��ᠥ`9l]�V���V7�i���9Y�{�e�T�ЀV�]��S�݂M*�VNI܀;���%��ťV��i��$ERy���Jí�c����w�:v��[X		��z�dv(�u�Y�W�6Ea�1ʁɖb�]*�]m�[g%j#o�Y�qY6"�)|U]î�����Jr�#�C��-֦�E��VN.9�S������b�J�ʶ5�ˉH�,'z�oiͳ�n���iȎmYe��r_�I�ɻ��7��Ϯ�1א<�]^�R0�.���:�f���[flWd��j�uwZi5f�ph�A;upA,9DK�J$�J�t���q�F��;ݭ�C4-��?-��=i,�*��:+^��fM��B�;���0�����hڙ�!�w����P�Mm�ր�)�9,21K�(���^krS ��&�*5�/4^����]�K�p;�F��X���7*�$��UFh�*�T�x3fiU`��o{%�Iiͬ��S7�fܼ�e��nm�̓i�Nm�2!OF����{�ƉLa���t��^d�L(�&�f�/�Ĥ��
��4�e���wϯy6��a��&��v�t���!1�o2dCԮ�5�6�
GFaݬ��`̔0݁����l�y��So^V�u>]���RK�ޔ-ǗF�o4R�`�I��LQ�d�ךhۗ�Z�����3i��E�����o.���@n��A{4��H�܊�e�t�̴�1�jG#˥��""Ȯ�S%+Y`FPwg2�<oٺ��ղ{V�iEH($-T�6�QR��kwux�pAo8̴�n�}&i[�5I�J	�SZ�a��b久�c�jJ�qb�����in�Ë]���7Z[�r �0��TT���WG]nYE��婪l�����8�Ȥ�b���5m?�[���Ua�XVD\D|
z�]٥�Ʋ�ՈMi[D]Fں���[Zf����.����M�E]���$˕�$ϚÙ�]��N�!\oZ���1f�u
��5S4n�"��^YD�t���t�[�8{/_mԎ�4�F�.�4b����,%kQ�k:m��A��
��qP3f�5����R�e��f7JIH��K*��1p�7.���Lɳy���wI�h]�H�+/)�̴-�~ƅnok�wT٪b�\4Xx�h�5�d7j��[ӸoNܽF�79YvayKBkspAt�2��!n4aPEЫ���M�b��u�p�r�2ݻ&���Qf�֊�7�o33{h����M�m6��7];v2h[�m�qb��q�u{�VsA6��}N�4lU:}ʬ&H�����)n�J��oM�wj:�_^�|�Z��Ǹo*�ݿ�[�F�[��ě�)��јY��Fl	\�u��ܥ��Vp[��J��bMfG��\��.=Y�ۧm�6�U^
����,�h;v�Z��ӑ|��#X��R��(��sM��Qwle;ɹ�sQT�<M�ҫ>M�o��V�d��i�8m��E�@�"�fL����ym�e��_Č����J	��ݍ�0n����l̿��41c��V7hj���e��r��^�i��YN�Ւ4�30�\HU��\T�uz0�
wa\mi:�h�SNI-�o7+, ��85'�蜭0Z)�u��L�V��nS�
�Lh�D�ܗy����9{x�z�%�N�ّ-/1yn,�ŗnX6�,���Kc
��i�O��.�"����lk�( ^�^ˣ��U#���8�)�[-�5e��`�*ʎ�ԫ�U��sŘ�J$RF���3l��IT�A3v�������d�G�\5yr�b΋ 	�c���RkB5��^�B��Z����x�X;��0��{xK%�̵n�-�t�5Tn�6�J��n<��7�`���	�s|E��2�tj(s��`=O6��$��X܈��q˖hZ-��zO�N�r��7�نԊ�����KI�w�V]��8�Zܔ�&ԅ���"E����{������	�Z�n�M�pS�VBEe��*;����e��#�$��7�2�J,�𬺴ƣ�$���*� �KYOh��`�)X����̰�z�̚LpD���+C�$�e=E\�g1[� r P�T>R�B�m�@��x1��e����� t&�p��N�V�e�h���`J���K��I�!t��Yl
�1�V^!&��"�cE�n�ԥA|�\U���,����3h8�lN��q�yYOi�PMe��s^�����5���J��2��K��-]��n�%���3\3��.�	�yG��YO\��q^�L�/(��k8P;yN9����.du�/3��Y��Ǝb&^�[�e�B�{j�o,��Ql�f�mCJ�������4����j�B��b�-����g�Xf���Io4fL�U�Snƺ��C/S���T�m9����7-֫P��ɣ�=n�7�!�$]�_�gw]��qWgU�WSi	BI��M�HIi	weWu��u�Օ��g]�$��I�	6���H�6�;���������:�.���⺨�㪨��*���뻋������;�����ꋮ+���컻���+�.������������:����몎����⪸��;��:�$bB@��I m!!����躮��*�뮲뻨�����芨���*�������躺���;�����⻺㻺���*�������.�+�������룪��;��:�*���㻺賻��ΐ��	�����%�ע��=��;���͗!��I���U��N)肺t�*��\Ջ�l�r�N����V15��	Z]mA���ô��Э.K��9S�.�����Vmk�[��s�����{�1���r�b��[ӸJDDr���#�i�;X��N}Z)w�ۘ*�,ް�e�,^������+�Rq�M�7�k�K�w���⹂V�Q����Ỷ(7����:���w;.X���1q����g�� =Cw�5�vq��nJ�K��p�w����x|��7�˖�V%��vr���Ŧ�Tټ�*'��n��R1k܍��י��<×q9�{��m,8.��r�V[몡�e71l�+
��;�/V�^�ZpB5�P6&i��-�U61���*:y&�ACmE[/qm���oyʕ�Ӥ�e-+`
�m�+v�u�a���ՖJukP�@J�gv��37��gT��M��o������a�om�2�Sn4&����|8�IJ�R	l]�M�v%�)e�v�K������(���p�ծAm�o*6���N� T�嘾ni��ϥ�33���ۺ/���ͽ�70��څ��rZѸ��gr�f5|>۷��=����c�:s��碆d����E�)TA�VQW>݀��=P�``��.�^PW��n\0�]h��\����B���$U��]��R���)����y$�L�B��\t��r�Vw�_J��O���͊-�
�h�T~9��	�	�X"a�[���ٸ�e�s�}�>�2��om_i 8�
��ƈ��v�!0��NW�Ɯ{��H^�N��ҞbU�sgU�2�&��{v�a��*˭��:��#(��j�<q�:uM���&��˔t`�nS�7S��dL5Uw��n�5Wϥ���S<�7U��#*��,�
+B�Yts��)a�kH2�3�-�aT ��Rd�Ga��^u9��]��QWF�j�|��W4��*�Ⱥ�k��!:������	�}�]��	�F��͡�P'� {5D)�٪��.q�u����F��	�@��iL�Y��Ӷԃ�c�1�%Y��������׳4�Z��Z�z��W�v�N��f	�Y���ڴ4P��b��B�m]ޱ]iI1ޅv��\$9g�;iTn�r�6�F�/N^V������>RD����f1�HJ/5��{{}�gB`�z���\�U�#�-�7-mwm�du�
�N�Hm�����1�
��/>�X������{��!8��ޫ��3nз���}}R�V���	ҙ��HP�f*�{v�^#agd��qz��'

�j�na�t:���CV�9�LX[I�F�g��I�v\ހv���9�T��7��4-�[)Q�c�d�
/�s�xz	f�_3��cv�_4�uk�1�ڬ	Zf�����~Gi�8y��U�7����Br��9��1�1�/Jd��9`��6.o9I�VֹKpNn��g0�km�Bf�p�Թ��6�����Mw.GkNU�Q�}vU噪󶂺+��\��Zq+��$u�hV��6ܻ��<�Q�UgIH�u��rӈ����lLÙKdP'�:�Ks��r����K�����{�FGi�#x嗚�>�߻m�[{7&���&dLc�[l\�.�2������R���"�Z�
>��ׄ�ov^�\������V|�pi��k�/�A��k�]��U4&r�q"bx۠an����a�j�@�aT�>l����]f���Cv����t�Q��M1�^�R��u�/��M������ˇ";l�ٲ�e��^�8U���ǼE�2;���^ʘ�mI���l\�Tj���֎��w2����SFkBw-�#,%�ي�]�h���mI[w\��	�6�#	�vZ�@]���X�Nޞy�� �b�=x�Ǥ˒�ج�S�7�w�+h���꾾w�Mhq��	�1����@��?k;Lޕy"|��(���e�2��o�[5ْݠk1v��Y�+Wa�teM��z�',e�A��.�2�>�n;(H�볗��ElUI�-=�N�����Ǭu��ѳ��[{W�����%�̇��a1��Vt0P��W�bnK�m2�,[Ǻ/����#��9����|��P��n��G�����Ok�ܶ��^u�Ԙ�T�U���.��͘.�ŋY"�/FlQZ��W�)n�y�P+"��1����N�F�]���H��9}��M-ɳ>�A�u��犲t��Nc��W��)t-f��f^��31
u���1l�o���XJխ���n�)�ʃ�p�u��Alw��^;l
�|�i�n�v��qal*��u�2������"[x]�/�WS�p��ɉ���:��K�F�ZZ�0�4I�!n���;�w%���kp>n�Ec�2mhZ�X�i�Z�V^�=�;�;l��[?���6]�n��u�L��i����na�f�����e.
+��1��3*��͢�+�n�z��2�aEe&蛒G�Q�K����*�x��]�V�D���}�&�W�5;��G���?��띪?N��]Ƕ��"c���t�����-��C"T`B�X�5B��n�eʻ����f�]�|��QT��	�P�9��a�dE��ou
���َ���*��⮖�p�����Q�PY���<�������5u�\2:��D��s�F��}}�W-q��qn˗X\����x�VD�m�r�:��\C�Ktm�LZv�Szm�44���ٴ�9:��q���"����;��	��X�;�Kd�'$��E��k���t�k1!�+�J"�k�R�2�s6��W�U"�r�]��%�/�tP��s���7:gN�Ȋ��Y�c%�p�0oK�ڮ�������S�n�>���ɹj�u3�du��n�Q<���9Y�t�0��ne
��W,�ca+�}�<�;�#Gt���"���a*�r�'���}H��b�̃��[�r�ܸ�o�溵l�hŉ�݇v�e�\n�9y2KmquHLZ5��`�!�;[���":�GL�j�q�8��"�hӾt��d���n(:汁Ģy��j�,����Z�o`�u׹��j]�njp��i觝��R9�rƫ�7(�ōE%�޵�:����Q4��C�7�7J��Jfdog�^Y-7j<��d)u�m�R �W��p��wcY�rGSf�oh��j��-]���,�Ձ��{�� V��g3j]mEz��@U�|)������u�Y]�Gz���8f��c��jMղ��dn�u�VTZqm���~�l^�ӑba�j=�s3"�S�H��jݮ=u��ذ��op��#�o:�z��+OT;�oi��JBӶԫ��=��\@�f��P�u완�CV��Em�̕�X��o�h�0�+d��i�w��t��ju�>|��Ljy��Aƍ�Ko{���"�w׺.�h�9#��˨K�sof���xCW�ݩ������K!��Egzн9O7�\鑒�[�|���B]�zrR�Ϟeg��^u�sFA�P�fNp�bRg]�T.���Iv�WQe����d�Ι��mK�0$1�e�T1�.�+(�r��EL�T��v�8�U,f�;aѓ�_9$��bd����,%B�\�/�e����՘���\9L�T���sP��v�:�e��oL뢪;Yc�T���0�9r��\�*�4���y�0�:L2�ˑ�vo3!�dٹ�j���,+�t�V3�n��qm�V��2�3�V����o��eV[���=yۿ6�h�MwJ�[Ј�q���a͠��;GU���w[v�bG��NB!kA}G�X���
o��6��n�#���Q��j?K촒9WobZӃ��L��]�e��̘�r��B����GQ��&�%����/n���՟��v�r��t9*�Բ�f�W�j�R	Ge��h&Y��B���6`����#��5gc��W�v�ۘJ��9}c�N�YpL�.�5@'�wqI�b�b�\�z�+�ƭ�]ૂ+꠹r�b�r�n�.��4���V�5n����`�I�3�X�?V��P�2��;Ԃu�ً,�r�f��1m�s���v�K��%��6�H+���M��U�����i�c��?���t�'�dL=ݮ���C]ޡ��N��2�=��h����ˊ�ر�(��tfu�0�B�ܫ�2�B���ww��gCe��9Y����Z)�qT�yE@<�����u1d!q�Aoj���1KfpưC��㗇!#��K#ou��s� �uo�.�6�_`�]��e��FBV�A.����o�����vLk���S�4�>:���AU��˓\��ێ��]��*\Y�_�nwI8�\��mpï���Ŋ��U�Q.d��#t���d/.1R���H�n��'6���a�y������t�%_;���٘#�|�F���N�:P�K:�IC�z�����'��B�ټ��Ү��&俱oU�/ⶠ�:���!+Q1�N���}�-���W�B�Ϩ�4�Va�;{���S���寋W3.����-k.�/-3�{��\J��ܢ����&7]=#A�b�U���9�v�Pܮ���U��"�]-"۪�tW}�p���j��!�AG���>���Z;m��,�5�cY��^����+1�Y#5I���|Zf!\��}:�K�I�*U�`it��JN����Ъ�a�ѦzԵ}v;m�b�@��Î�T�W���by�1�7q��бdq�	�G����뮹��X�C[V��.�};h䂲��c7FJ��-)��Z��:آ÷�t���Z������vUuZN���k��z�7s)e7EW'Э���,��5k��[)�	��l�n�}ջ&+.<�Wa���j�L/Z��S\xv+�fa���G;��ntNU�m��x`�آpU�{�KndX���E�P}��a�ui��FuvG������U�X�]��y����%F��q�ݗn���]�Ô�v��Q$a՚	*+��B����ȳ����qM�r��̧�U
��j������IA�76z�e�%V�d%��$n���Pʹ�/(�����h��'S�Gy�v=�k-bD�q:�]3h�ew,��quwK��j�)��E�s��6��b��6��j����Ӑ�#���Լi�ڎw)O�t�C�U�3ljk6`\�]�ݦ�y��]�]eu�&Q>���vr�4��sv0��z�o����-���{�[*�9�U⮦+���һw:���R�:�ѝ����b��6тz����R�ǲ�w������Y�@�J����X$�Ī��A���c+:�Yy;��E�L=�H澾L�,���NT�23tF��U&�j�8�9Ck,eҽ7ב��ӷz��s�sh��1�̉N�:�z�P#p��sX��cɲed�����	N���2Z�7Y#6�$��i�n�(�u�h��KK�ྻӖ)b2�wu;��UCtS_
��l^t�%�9�DY�+ML�*ͼ�Vaͫ]C��� ǥ�m*���A��%�SJѳ�<�2�Cb,0cWIf_lu{�2�C%���=�x_�<n�KU��r��/1f�[�N�y��t�+�ܡw�i�紣�{�*�г�%f�ʛ����=V��BQYB-wy/f��Z̉l�|��U��3��e�ل�:T]�pY���^�c�S���������M����	�ٴE�bb��ꌅ�w)Mʔ��R�EO����M��T���_!q�ï��v�-;QB�`wJ��h,$Z���Y��t�{��j�lڂ��.]N��+6ss�ܱ
���ZOe����`W���ë�e!|:����S�4&gk�R���
+--m���!똞&�>k�)�2�S{�J��R��0�I�۝W1;U�*gqـ�3(퇥���[�+H �Y:_cz1��\���g��y�[��Y�e]^�A�Sȶ���[0��]c��M�kl�U�8g������g1�uŲ��r����LF�7���`y�uL콭��X��j�ϖ���Î��c�xmK�!��x��n��h����\�Y�<�C�7����iA�v�k���^*�32�VcVd]�`�Aء�`��~�0o"�R��1�%�#���\yE��ˡb8�1r�U[�#Y#v�Oj��
�徒
{�1�7q]d��B铧gR�6b3 �S6X��Rm2�u��Je��ٽs��P��O�j���'OAP#q/�.��N!���8>K���P�s^	c�ּ�;�o{�)D���n
��u�=;2��B���똧K������j�;��\y�n@4ꋧۜ���B�B�qv����K����f�������R�,9Y���
]/C��0fwk��v
�cU�:æ@�b�u���%�%5O��eu�9fiYۯ��t����J2�_�l#��R��9C��EA�i���쫤J���x��J.�5vm�aRy�ܸ
�y,���>�]f��bI\� ��<�z{�*�-�{I��)�F�Pۭ���$��X.Dl ���nWU��)UI,��κ��W�o��j�IT쒳]�#��fB��soEհz�
�u}LQ�w�5�i,�}kM�R�v��b�-�/���ͫ��sz�����Tu ��cڝ��w���͙K����V���c�m�sx(�w�Q�u.af�pW?�v	�*���Mj՗���b��s.���x�i]��ژ��St�zMMv$��1�m��Ǡ�*n+��w�dܵ�e.�y�}t)?�k�x1=��6���`�V��C.w=ű6F
]�M���LB^_[/py�.Aw��*d9IR?=�^͖��զ4�����W:r�����N�
���ǁ�4�Df]�B��j�[�9K?U�5Ou�y$�eM����e#�7x�9mђ�l-�zvI��5].˝�t1��������IT/{���_�O�i�[]��n[�wnSlb�(ޓ� �'�se�
lp�;ng�7-�%��fW��8dS;B�q�zwL:�g��;*h��K�6��j�GZݮ/Kے=s �I �k\mSfM�4�ݯC˜<<u�u�GF�e���ݮ|�7qn��nמ�!t�w�B�:�V�;'��
��G@>N�㐃��K��v^˅9���u��Y�]���{k�t6}�^�uƭ;������E볶��|cI�Ų�ĻlF%�{=�y����챠v��:�5���[�m�b�y�M��s��6���2/Y|������;k���m���f��.}��d;7`0�3��^N��0qR�}�Kv�� ��;�]� \�1����ۗɩ��=�C>�����>4��Q���rPnnv���V�PvÍ���]�����p.xnV��y�>����a�x�`�s�:Gu��n�5duN@/X�;;ָ;U���Z۶�y���9;A� ������ z�:���-��.݂v�sm�mv�*�b����ػt�u=���c:�B<Ǜ]��wa�=���є�/l��C�Csn\�1� Ք�]�z���6�6%ܛ�z6u!��n�.	o�\���q�����ƶ�s1IɷnP�n�jvMn8[@h�U��@֫�eݹ���n�ⶶ�۞ۅ����M�-vf�/<���v����������m�v<A�ϱ��1����9A�\����[��=���!����]�t�cF�ȗc���v 5���5�jh��sm�\;`"�p{m��n㎵��wXN#��qi�{m�n�:x�t���ǭt8��M�\l�9�OFu�cu��)�um������u�=c�=�y��]��wG��2jwb��q�kn#�n�k3li�m�i'n �X��7n�5p�:�Sv|s۞�v�)�0v�9#��sӮb�j�F{k�ݷ��]�����F�s�L�ƻ�o��ng��<7Prg�{uy��uMp���Ԛ�#��ņN��n(�v]%�KNn^����D\��#���7\��v�[F�����1��!psqr<���g�{N;FGw�z-�ț�0��֦ի��E�έr�u����cn��6vۭ��>/9-:Mm�έۻ:�N9.q�^�����������[]����#�	p�V'�у�l�n!�)Zܼr.f��M�v7�\Z��Ѳ{Y6��<�8���g�81��G%�M<u����Ʉy�ܼup�{X�r#�m(4���s���P�ۑ��{s�c��OR���]�c��-[+���p��;��X��A볊|1v 8w���Gs�/8i�,]�-�qF&8-����Y�u��S���I���5�u���1s�<��nx��Ͳ���c�=F���+������{ h�ku�+ϑ;Peu����ͻS�]V�{	�{�Þ�9ݶʇW+ر�7Lq�@�7/!�w9x�1�8��`�-ǰݕk�u�`��<US쮌]�k��tz�|Y��&�-�y{����ۧfNo q��K�xk������ۮ�����{v�Ƹ��"�6�0mͺ�<���{unxl�q��o���熞�ŶMd�i��9�&��瓞�p�(Wvwnv�;s��������u��M��&�9�!{=gn�A�'h*W�n�o$/l��PpLq����c#ͣ��vU:wz�9v��n�r�o;K�L�uv���t��sѱ:�O6����Qۓ�xom�β�Z:����۫two[�y�5m�3lA�j��v-�v\��e�+�f�
��uɸ���c��\&�mƢһ�Q�����!۞��<�Ƶ��zۭ�v��z3q��.���U�姜�.�:ՋGm���Y�T���:��ӫvp���`)���J6�ɼ�dZ���wn|q�q�Ln��Ul���g�ب�2�$ط^e��P;�d���q�Рe��vR�B=D������wc@�s�9�yG���od6�c.��yq!��KB]���:kcgl��9�Y�v�wcr<Z����&�o{s��K��mW��h�㰾_v�Ϙ�[qd�dq����AQ=�.�{O��x:ҡ�4\K�D�۹��ҍ6�g�q�.M�hŷ�&���N�/A�۶�[�jz��8�nW��g�n9�v�p�9���79��*�bv��kvp���;n��se�e��c�A��ݺ�#�n�6x㒓���Lm�gZ{W8�[o�г�렱�zL�B���\�1��,Z�ۀ3ݍ��m��n|qqkc="R�Lqz�K�U�[���N���3���N^n�xɪ�Z�\�����.�Iu^v��Y�4s67g����/"�iq�kV��m령1�1�l�f\[l�R�p�Hv�� ra!�նm��Ć��\[�g]-���m7	)���;v֨-瓓�v�q�Gc.;��ukͮ9M�bݗ��۳���l��]�d<�&:��,gͣ�����r�]nm�ڗ�j�����k���ױ;��������X�A�����v�.tr�RK���L�ew3�\��v�s��f;��Z���  X���0�n�b�66�,�k��q��Z���j��;C�s���7&֭χq��,V:r�W(#��y�v��8�1���u^��spv7N�[O]���C���9��Í.���m��	�sr �ͼ��s�P H�v,;pgf��Z㦫v:�y��9�xx����n�m���g��r��u�Iև�[��Vx�ڧ��'�k΢�hWts�/w	���cu��%����q�;��������odۄ��s�����J;K�K�ggGk	qqb�v�#�s�v�Ǳ�q`%zZ��M�;T#�]���޺4�:�<��q��Z{u�`��4Hp\���������,���\�z�c���.���C�d��;�r�lm{���:;g��:�jn2�ۛH����팠*]v`
[��8�H�.�n���v�r�Ż����;�%�G	>۱�O;�9�ù��<�'*�ѧ��\�j�uŖ��k�t�솵[�s�5���L����wl���N�[unN�wK;S����G6]ă�CЕ�ǎ6�w0��4��� oWY����mm����jNp[�nS.5���d�۰ܔ�<�ۋG<�u���[t[n�k����'7�kF�f��rnˋ������e쥎5�lF��v�DF�����f�sX���vE3���\�W -�9+��;`qvM2�1��B7d�����vS��l�솻&�ѯ\n�
��Z�fy��[ul���<x�D�u��}y�F�^�^Ǝ�Owt���]��&&�1�u�w-q��v�<��J=���
1x����<�/i�K'mD�VNz�ۃt�WW#Orvrv�v�&[/��Uͻ�s�v���i��t0[������s���N����]�\�QY9���fdӕs�66a�.nv�L�h6ݎ���	�[��˱u^�#֑�LcG�NR뵦��D�w�y�Y���Xc����h�Zi��s[���H �磔��F���dA9���k<'	�%g��'b{�!�y���t.������v�*+ç%�mE8�e�N�']�	i�Q�n=��ln���&^NtziVrli��k�#�z3�^ݳ��{4O`��Pݮۣ�϶:����æ�c��86���{�7rA��r�p�Dqn�	Kۏ���%�uv��cmp�l�sٛ�ӛ�v�Ir�3k��滷�
��'�}���ލ[n��|yw0���q�Wn'�ͺ��7Z�r���9�pz�Y�t����n6�;�5�'�[�݃m���Ҍ֘�j�sv�E�+s����-�;G���9ݤl��\B/���\�L��j:v�d�Vz��z�:�
r�	�Zl��O]Ol�qM�s8�.,�W�ZR����#�5���)ʍ��n^��RmnJ��Pv�	���'�'d6\��)ɝ٣����=����]��-�-����Q��Z�c���Yz�k�Z���rv�J5n@C��Xi�۷�Ns�\���-��m��ҫλ�m�[L�ۛ9�pW>͹�x�x�n�-�;`�ӰEmy���p��gn��G$El��{:����8��f��<۫�&�Ŷ�=iܧ,['kZr7�^�Lgd��7[kF�y{V�6�l�3�{r��S�X֒���m�VL�.�=���KsϨ�^�3^v�����ΰ �����'\9�c�+��,*�2q�v�e�s6,��uu<r�;a��C��ͫZ��<�$����y�(�[���q۟\u���ć��ɒx�}u؂��h��]sn8���".l�͹�;]-�nE�9-��tt9]��LL"Z�r���A/#Rݶ3�u��ޱ�K����C�[���V����@pj�k; q�vTG���`��b4����yJ�F����m�2y���lQ�����b"������7/�����۷1���rݫ�wF���7=�Sn�n�&�nu��ܱuGj��nD�{vq��[k՘��g�h�D���:��kq(<�paM��s;G&v�n�]�:��9Ms�G�B����nv�um�]�ݎ3����\ur�6�omI��*��\\�n��j�䗖"ݸ��N��]������f2/Y�o<=W�8�n�u��:&Ơ�mW"�ۺvnS�ݺ�x��nP���j��CqE���+���6����]ۯj��v�����m���
��]�O*>����z6N7E��N�8�:����t�v�Ƅ�=������=l�Q�,�`�.���u#�K���L7<x�ʄCٻ�y�a�n5[�+�Ӛ^(��z��uI���7\4q�.�V�掑c#XzMQPUL�Z�\�G]qm]
ڳj�Sp�%�qyHZ7l%��k&�Ɓn]��࣫=��M�����ǽ���n.��e�_�i�fu�FY�Q���N���3:��*H��C.��eͮ���iǟ<��J��<���.(�β�;���:)<�˲�.3��:��,��|�<:�ڽ/&��w�����:�8�+�n�;+��Q^���˴肳�����:/+.(�^ՑqO��':�l�{w��kYGVdw9ϵ_;˳
�j��ʼ�����)O�۲>ZZYE���;��.���{u�fwG{k��2�6�]�vpM���{ء;��:<�
({vE���;,���$��,���[O{�y�y����w%Y�b��|�^Tr\|����n��4��<�����Y�gchHλN�f�lu9�� ���{�{|�:��nl��V��=n4�$nc�C�w8��r+ζ!��:���`μ㫖v����h30�s�P\�GE��b�r�+��E���8��
�ۉT���W;�e]����v;[��%e�D�-�=@��>L�v"ܵ���I��,���ջvx[d7\�&]�qn<[�-�����s��UM狱���v[u�v�s��`NT�4��$�>�?��-�{��;�ult�9�r�<v��7\��t�7m�X����Z��72k�x��̽�v;��X�:�O�n���̙�7����םc�v���&�۱���q�����]\����5ml��7]���x�{v�2#���ra�nۣv�<l!Q�ɻk1��m�đj��[���,Z7B|݌'�&��:�:n�Asƛ�X��0�v�"Z�be�:��o)���W��s�@޹�o �p��fLH8�Cc\b�<ո�۶���Y�����'���m�ׁ&�=\�8�{[����s!��˻q�|z�1F����L�(o�+'��7:�<[����k�ݭўW=;��'�b�������]���ʻi��yoV�;��bF�9�u�F�N��mv��ݸ�t[;�ۆ�M�Og������6�u��ݎ�vc������G[���h��tļ�V$��.㮷n;@������O���]ވ��;m�3� \àݍ.��rgr�Y%؈͑���^x�<�����]�!���-ͪʮ�9����녮�a�������D���,���Q��x�m�br�5�b5j槸7D���1��*��	ʛZ�u�^p�O\^gb_[F��'�YM��W��m�]��7](m��x�'^n��Q�u��L�n�����w6yM˙�/e�g��̳ó�x��Gn����]q۷v��2u�V�=C�Q=�Q�B�v��RF�6���>3�<�.y��v��oD�Vt�]5����EQ��@R2B!������{*a�=��U�Q�DF�#M�D0�J8EN��r{r����Da���^�L㷍��۝��d2=�m�S�e�����V6��({ǧ�4�y�v�m 1Pj9��CNj@���w&���^�B�l��!�	����L��»���e;r)��\�#�y7�: �i�H�?~}�� VQ�c�~g{��l��~$HVr�p~��F��'o���h���*�%e`�,�|�B�w!��8�_����(����Q]l>�̞�~IԶ�������R��\P�W��f6��l�M�����g	}&�$�坔~��
��,]�y���k̎<͹Z�ƴA�?r�P{mB��*����X]��5;����o31��ԇ>������ʬU�=������~���|+�TWB�rw��v9M�^�*%������lo��lq؇m�z�c���v��G���`ن����I-���/�ӽv��X�-a��߳ ����U
9;ίa(xܽ}�
ǩJ��5a��V��bŶw����G�����qi��f����No�Ԃ^=�W��'H!�F]F���m��bft�����=����	mhw}�ʳ\�®'������i/P?λP�w�����Zӧ�.O*��6���vX9TCӾ3��o������N��]�_���6�� 	�5t ���ى�E�?8��N���g3 ��2����Я���LP��ӹ�_�K�Z�E��x��w�+���� ��I�Y�ϴ�I��3Myu���B�>�{�~�Z� ��6P���3/�&b�^y���a�v�g�\��.^tay%�֝n��a��ۥ7��Bk�;���SB���gOl@P�~�`�͇S�˦�Vh�������sW��M��*�Xk�;�t�3dS��5(
�y�^�ܙ&:�:���V�ݧ�k�D1]��F��bŶw�����T�Ao����j�ر �lR�m�r��m�(9J��6�n�߯��}�Z�����͈0֍/Y�C���(fu�T��i�|H'�=~��}����n"j�)�Aص�����V���~ ��ɺA3˷�ͥ/�o��`�{ӷk��ʹy�R�Pt�W��bϛO�;p
��FWs(��������<�M=���4lyɲ�˒�Wk��U�.�i��qGi����`M�^�?�	UP�X���R��[ݮ���aP�tE��}��{�����$�g��`=�gK��B�~��	97~$y��,X�y����/����N��� �sj��I$��M߉���gݴ3�vׅU�<���\X�qf�*�*�Xirg���$�>��$��:�����A>���I�����U�S��\�YXԙ��~����0�;���(w��� 
6:�I���?y׷>5���]���̃�u�����&gm���𙃝2o\ޒ�cH^�����;B�`8r��g]���"u��������ޛe���no�I�!�q*�*�F�PDQ���Āy����i�MX�̲�Ogy�0tw��N�7������O	������y.+0����r����7]�6�2�s���m�q�Ua�rs�|c}��\��������'��$��?n�
e�vѸ��Uu�� �G���7�
�X��=�06ƍO$��c��� ���Z ���� �~�'ms���ŻZ)�v�ł���h>56� zy�~�	����rO0+K�����"���o�6�V��yB«)yM�r����q����4��\T�%��p��,��J�]�
芭Ӿ�z4�	�I�
���U& q��TOf��w6:i��4n��2��L��Uޯ7nh���g��#,M�/���B\pBj�����������J�I�]j�X�O��ΣK�2��a~n��2I$-�,�v����R���E�����k�>M�x^(N��؟d���t���[S]����Fӱ�{n�s�O3t�lvǝٷ�����u�9I�����շ:����<s�nh��yr��ͣ��#�n�1)���I��x{O<��ƹ�+NΤM��ac�8{Gnw1n���Z���竛WK������c�x�s�ݶ52ۧ�g��rg]���=	�,k��e��1�������cT�/8���K�,�C��e���I��=:M�uH�;��ns�������7踸ѹH�ԡ���� �����9pRg<3Ͼ�@�C�I�	���:M�I��ۤ�wA����}|�
��_R��U`>�ٺH��0h$_���]���+��{t�H�I4o�4���ʪr�&g��sGw��m�v�5ʒo�OĒ;=&����D6-��o�||��i����17u�V�#�V�Xk�{'7��G�Y~ե-~=���&�t�ӛ W8�3��z��=���ԡ��u�<=��ǔ�l�rgл�c[�6�G[Fi�Y�PeIS��x���;`���y�{���7ӓ�>8��T7�g!2����W�r-����9�߮��Uٳa]Z��>�X���·]r�����?�ެ�@��ӧ�/�pC��.�]K�e�gC�u�J�q�OK��U<�z%���ӫ���׋1��CW�j��|4�Ho��A �a�����n5~d�,ޜ�}��6�q��^e��3?>f�^��~k���V�����'�~0�{,��7�
�5XU�����5/�db-�1��x떀�����ɶ;������=M�*�-M�,�1?9�M&������w�z��?_��n��8�� ';͇~�s���s{��Y]�U�(�d�[�1�\{n�=��2�W��\M
U��x�u������Ԋ/3(�L�|�B���(|��61�x����B_�G���?���R�f�劻ll�k�(!}���n��ږ��  ({�� ��6 ����{�v��}���W������Qm"�I����!�~ߴ�AS��{쾤��m���Z��m\xĭ��Sj}J]PSB�N֎*�����%�Q�`����+5�;C�����\+֘K��:����R��ٟ?N7�)�Z����3��x]����
��	{�����o��W{�m�Z�H{������Q��
�����M�4�&S�$DI~��{[����g{��pݡ���mY
IZv��\'�����ø��R[����	�:�C���ՈjUm����n���w���
w�����{�V��h��s���������;:M�~���+c��j	Xk�gu�ϛMo"������a�ĂFߤ� �}�M�еʺ\5�Μ�M�s!lT���3>O7�<�I�~���I<�f�x��6㛤�}��w�e������a]ڡG{i�(!�B��S3�u�o�H ��zo��5=[�d����.�0+�������P�P��t��J��EDbE�������ÜF
��vܨ*�z��wa,�f�����s�-�������F�P�T���~����<��$�kδ���e��3@'_w�h$L����?/է6����ߥj�{��U6�/ԲP�������]�su�W)ڊk�>r���8�a'��~w������"¿�w���Ay$�?K^Հ�U�!k�g/:c�w&���7���8���yŖC�Y;5n�0^�zn�	���`)�b}5Uf��o0H���+c��j	Xk��w1��)�4�i�Eyx��ɒ��#�ɣI2׷�j*Wt-PJ���:睬�3y�F�u�z���=�����e�+�(
��y�Pº.��f{��8%�uT,+�t(�Q�C����ffA�˱���� +��U����bݵÃ�:�X�xt�b�08�Vi�!q@{�{!�c���:�2�Qx��к6����I+��	St�ӖJ��������:�ie�2d�QQ��5�J��g>��[���wYT���0=\۶���9�<�\.3�w����/k��t�N�e�r;[g6Nr�d
��ۚ��Vw=�p<��d��X|kA�(�\n�
ۗ�]l��Qq��t-�3�I�-��ֽ�uݑ`k��'�S��q��..|>#�:�O�-�=sr���8�x�S/�G�U�)�{e�b�ͮ�q�V�	���\�S�O<��.��=`m(��mk�%=��*�JԒ�߼����DQ�e}��޿&��i�
?H��{tsq�ϧ_}�rf&�m=ә����[��-c����鏂��`1��n��: �~g�����*?�k��dw��[���]�Ev����O�;�b��m;4����%� a�i|��OSU�b욻�Z8=�&�[o�߇9��qL�D�F�t�>��=o}�;����D�"����]]Y�4��ӯ�{��c���
�D��^��H�~�7�G��j�w��ե哼�JM�(����T�5kn��]!�]���ڲ-�lq �cQ�4�P��W�'��Y5vn��t�Hkst��'��7~7��aKϨf�L߉^bPP*�j�;f^_o\M�qm8���Qxӽ�֐՗ژ�F.��f���dQ�|��S+@w>����Y{�Ď����%)�q�pX�2���$z_��H����+�}͊�o|.�a!�VA��}t(ګ�R�3w&����f�H$߽^{W��ꙧ޻��	{���	>���~�9��V�v�gޜ���Ŕ�O� ���c� ���l
{��+�������._(������w]Y��c��R+G>�2n�H�G�n��?Z:A!l����s ½����z��s<����ڬ�7+�U7=r�5��:ۮ3֭t]M�b�zV�(�
Z��=��Ĳ��p�I�\�w�P-�&>=���^W}w�kΝ�L$�e�vM]��G>"�� �/��S�;���)�>�{��B�&���x�.��fA��Є�$l�h�7����T�<55���o����a��X���h�ͯ܇u3xS����6:*mlnd�]N032P�� �Ӄc�ތ[P�':�I�������G1cC��Zkg5Z�=#�83e��WɈ6�VΆȊ��)7�v����}�Wj��]:Ge%ln.�^�e��A��\\^'�o*.���Wf�j���bP�L�r��R�Y]2�YĲ�4.d̊r63�aAv+v#Z�]Ki<_eV^�E�v���ڜ��l]v[३}
cD���N��uٲ�����xyJ
��f��A�����}��,_Z6a�B�ѽ=xm�n��KG;1A�I��n�j��wa�A�v�9��+l�i=vx
�9֔��
ח��r[OpM�eT��b�wW{{���Ҋn�.娮�#4�[�1f���M�MLMN���(�nk5�еrH�[�;yiH�*�px�k`M=�e����Ĉ�ią�N�Ԯ�R����S\�w}Wm�P5��}Lk�pl\��ح��Nu�gvQ��$���^A��ԍ����UX4��Z�����˅�+7z���.���^	i�Ӽ7{pȂ�(�CXy�#Q��Dd���͠y�}/ݽu΅��@��-kh?�z�e�U0�g]ͩ;Y���s�sK�x�28�z%7β�����E
87.��n�b޼�wbP{|��Y�o2�Alc@������˵�kz�����f��$�d^���Cot��m��Ĳ9��]�\6�,쭮ÆV��ڕ���Iǒ�u���4/��GetG���n��U����=�z̎�W�Ï��O�HG�~�����b�[6���à�z��(���)�^��;μ�yGtsk
���QX��㹭�/�Ŷ���{{x�:m�a��.��|�}��;�÷��ї������8������wE=�嶯Fלf��˃���.ʾ������_.���Q�eon�C�:R��u�6��;=.���t]^^s�zĄ���:��U�q�w�y��Vu�^�WY���;���ｺ9���Ygt���޳<�N�&Օ����/;��+�8����z��vu�n��]���:��ܝO�v^v��ok��i�ݞ��ޕ��n��2���^v����:����^|�JmW�����Y�wǵ{oH�N��<n��zۯ,�{��(�ݙy����l�m�˱���on��op{�4k�W\�ck�������z��W��g]�3 &�m{3�9�ٓ�غ�~��5N��
�x��������w=5E*ء��V�M�d���,.͛�k4я0YnO{u\��k�;8?s�m�@| ��e ���{�;�����y ��WTjH�P���U����Ѳ�z��h��z�ze�R[b-h������P�*EG��޼������
�A��n��+��z�ȖV�j�o��
�����li�yy�YF��U�u�=N̎^UW��BI<��I;�=�L���Bܸ�j{зc���5vU]��G�q�K���h&>�C�
e^���A���ֳ�T�w�:>������2��o��zs<�iܡ�t��Y~��$�n�L�qQ��_Zc�<%>)��K�y�n���qﰺ˼�I�������k.����E��cΔ�w���ʺ�I��=�=�i>��4��s�J���V[[	����hI>��h;��_��^VC�o7@�BMA���T�*7��Ux%5Z�K���n\Z����d��b��v�ܽ`���8{�5Sj�]���u�ښMe����$7�t�{%�ƪ�+^@��W�_OjϮ����rK+"���{��M��L]<:��j�?	��M��$�����D�#���\��wq�bξ�e*���&cs��LM����.��X��9A� �c��$�6��$	,,F��j��Т��Zs7��L9��{Ɲ��L|PF�ߴ���-��Y;*��7ۺ	A�4����,��f�n�H$���F7goM�� Şm� {۾l
�~����=3� ܫ����fe7\6L�V�t�m]�L}�95�m/yޙ^d��T�yL�w�<*����Ʃ\b���[d�N,�r��QQѩ ������q��(p+��[vv�����u{[�����!�zݻ����'�n�3á�r��Ҕ�.�ƽ����u�*K���{{>$�m�z<�t��7-v��zD�v�s��ܶƚ���j���~FCq�Z��˽^@݇�]��j�c���x�'kCj8��ٵ����ǋn���n(��s�`��Le�w)�]i�b������������7�>�@�R��[ή/�բ*䵸E���؟��nf�I$yW��C�r��g2Y�v��4�m��O���6I"�ٺ
�@6{�`�x;/H#�9L| ���� �~�J��������*� ]��u�wtm��
�얨��	�%�=.G��6����W���>��Ջ�j�5�vO7�dΧx��w���	�8OĎ����\����o�|t������pV#V-UѺp{O�����_	�{�%9�H<��w���5���ȼk�����%b�A�R�v;>��Ԛ�6C�2uu<s�e�ha~���ro|\s�A�, �^��Θ_\TE L��t�㢤���mIۤz�v"'6�W]�&�P֗��L"�[���0������f�b�{sʄg�B��NU�Tf�a�<,WT��*���8B"vI[ax�Ha5����Y˾�*��܁@}"���
���&[���/]MR��t ���.�����	f{ۿJ�Y�����I �:�0�����{)�4Ý�(�v=kZ��ѽqg����<�[y��w���Ɣb�+|��-0�bD�y�q�i�1�3;���b��4sse�mp-�hj4��y���K��-t��{{��7��������~�v�Ƃ�b H{���N����u�_��h#����A����~�}H�V(�6�w���alQ�[���S���v�!$����ˊ���6�.�Nmsq�Olmc����/��G�<9S���?|����C���A�h�أ��yܢڶ�j0 ���;�}�؆�W�u��]^��o5\�4q�w���>ADw9��[��=gLz���68m�q��s�G��6������s[��-=�n������1F��s=�[E��4F(���QlV�4��is��7߾ʏ��2w�]��__���j4����7��o�� �V��24o�̠��Ab=���YH�������g
�W����<�_8뿰z��c��k�r���or�z�8\cGVX��sWa��̘�P�E��i����]f<ܢ��Ͳ���u?|#1����H��4�Q�F$� p#�~��PY��fʲ�~QcDu�o�����w�:�b�a��4Vw�R8�6�0"���l8�AǛ��H;�����5�^�w]؇q����v�GynlӸަ���ǽR�1{���`��F�b��QƖ�e\�z��t.0��4Oz�E�X� �{��8�c҉�҃Q���R\f�j��Mo�3yy�}�g/7�l�w�N��ϵ��[h�н���i��)�,��y��Gk�� ��?.��o���Pc��8�I ���Q˂$PDq4řU|A��L��[z���f�U���ko��ԋj���(�&}�z�im&�����`�ݔr)�!���n`�(�����Y�I��[����xj؆��#}�����F�'����p��+_{5�}���s������G�Cvkǲ=vBM�c�����c��v�e��iF�iG�swG��F(�Q����{�h��_|�h�4F���f}���i�iD5Q��9�������{�֍��:(�4�\���y����ZoJh6�b"����"H"8�G�*��3��6�Ͼ��E�7��e~u=�{��w�p�"V�l��i��Ah̢R�S�����D��ON�}t�����vL�Sp]:��9���J0�>��(��"﫺�l�7��6渋b�ٺ��4�F(�4{�fQi�ikgף39k�S##��}�؆�Zq������ �!��D}�=��bf���Ժ���c��D�1	7S���G�)k��m]k]���=si.�'��[����>��[,e��Hi.��f�iF�iG��|��(�6�}��8�bG��|�ϵ����-���ޢجa�҂j<�n�`qk�ML��RMm=p����=���"�~��jmk�s�Ϸ����� ��4׻����`F�����"؆Ս(���v���N�=�{K�/�|?���fG1t�9ϐ�X�=��A�Ѧ(�1���}E�lA B ���̓�]\� B?�q�{wH8�8AD}�gԋb���㚞��������i�|ϲ�fO����2�%M�5i��J?}��H#Q�b��{�G,#DM�ϳޢدX�ǅiSQ��z����$-�\O��kQJ�b�%����Y��h 8�I Ͻ�Q˂&�������F����}���20#Q���ԋbVҌ"a�w=�����/~�؍�s����s�ǲ\�ǅ�fn�Zx�E�Y]��,��N�[=stp�mv���+��.��A��9�3(��>�6�l��Qp%�L�x�*-Q��"q��UH�m��<V�[������e9c[������V�9z8g��X^8�[���x���7[S��v'���veS��IȽ�+���<�M��]���>�xp�n��T��2'զ�:�{r=:��OX���|3��r�]�x��;�P�ۡ��k�'5O:d8����ACqp=�8z�プ���Y�Lqj4l�)���m�ؔ]�1t�ѭ��ERn|�$��'B1M5t�5"Ұm�r��djU-��vz�ڕosM��G�h�y��b��b�#E�3�,��j0##,���`[#A9������h1Ǜ���sPCb���}H�cA9�r�;��ַ��7� ��{���e�5Q�Ww��{s�������4��a�DW���E��lV3;�z�b���)�\��=��r��_=�7�Ki����j`�oz�olz��L����-;h#�D$��z�1�"8�G��s��-�Mi�9� ����Cj3=��"ڶ�j4��;�z�alQ�w��p�$���٭�#G�����O�n��E1m�bG���5m(�������{��-���Ƃ8�׿�k�k��f�m��}��vD�G�wt�v4�_u�5=	4�ܛ����c�=�-�lCb�����8{�߉[�ۇ9�xT�6���y�E�X� ��>���l#J5��׿�.4��rs;�y?sz]i�$U*���M�X댣Z�Y�����y���c�T�����8�a'���ϼtV�4�����������������"1Ƃ8g=_qg3���=�w�Z߀m�{�G�׆�`{����b�����V�٭�޴9�[E�G��|��F��F/�E��}zת�f����7�nº�mѽ�`�+?d}��̴��G(���$Ҩ��O/��xY�o��{˄���.N�Ю���h���Q�VҍF���p���q���9��H8�9Os;�׼��ñ�g�ş�E_����IU��k\A�,�_��[5�b�{Q��������YY>��yz���:4F�4F(��}}�ح�bJ'��g��|��Y���y:��e����F������V�sy���|8�I �������s7� ����������R-�W�}��������b^kQ��f}GZb��:ܳ\�Y*�����?o/t�'�|$���4o�w(����~���N���r���#A�y���A�PC�D��w)��WU�Rw��_�n�y����O��/upX�ܷV������S�ܨ����ӏ��1�6W����bL[�{�-���@iF!����H#Q��D��s���h���nM:�����q��g�G�#JF!�go5���i/uLOj��q��4�Ib!����? �#�>���>�������� � ��7����#؆ѫ�r�ƼҌCa��:�߾����E�ޖ4������s�UR�Q|��ƈ��o�4�6(0��̢ڶ�j0"d`?t�2?P����^�RΡ�
�9��y�׵v�61'����fۯ ��'��*���n"&6�zno+��9���(?h��f�va��F�8�@q����59F�߻��;�_IKJǩ��G5� ��+�q��n�~��\�Ս(�Q���q����"�}��-��#Dh�Q��{�[3��ܫ��o�m-5Q�ﹿ�.&i�5�ߦ�G�=�Sz�o|-�l�}��#��1@;�gh��g���z�;��y�A�o)b)���~��-�Q�4����v�alQ�|}�例�Fr�`��K�y�t��ӯ]d�w7=���#��'%u��+;���������g�%�K'�C_&�g��1c�F����ձ�;��`X��oG7����W=������AF�� �"7�ܤ[���k�O�]��{sZ֍�����}E���'��Gn��6?����ƃ��@DQ�b�|��m�"#��v�1X�4�Q���gܧ�������W|��5~��5H_�+��W](���CIc#G2��N�8�B@3��h�"B�}��j��2}����A��j3}�}H��4�Q�F�3�[b��t�V�7��=nR8�7�������3|e��Cb�a=w��q�i������=���F��_~� �?/i���fog�Vp�*�T.�X/�-A���}˽�˻���x�Y�4�����`4�=��b��u᡽��ܪ^�w��P^�� ����>_�3�E��w&֗���Q�j�F�r�G��J5Q����M-0�o>�Z�W4w��xM�m����-��#Dh��3�q��҃Q�o3_m*f���Ň���$�k����vR�P*9�l���C�Wɞ�]��Mѹ �����C�����Cޞ���oOs``��ｗAi�A� �3�r�"EGA��Ԃ2�e���&�X5�g��e"؆�6���v�ach�xw�(s[�混&����<��h&�ܭ��g��2�ty�iF�&F����ldh#�Cy�oh(�Cb����r����f���y��G��ɓ��ɩ��`ke��u����g��M(�1F�4?o=͙�s���_u4|� ��;�gh�+C҈j5���ܷ���_��'�]t�n�4�������eW�r�!�I~�v�[�D��9��"B�Cp��T���������R-���sU�i|�ZQ�����0��!�Շv͚oOzz�$�-��#߫{
h�Q0�PF�Vg�iWټ��g#櫔���L�w���0,dh#�C}���
Rp�$"9Yܤ[��6�����j�>������m�u,���6�6q(��v���N������+lka�x0��]���l�O2�Kl�{����B�V��h���/�of�] Gv`���ܓ� ��ӖTl��u���h�󊇽v~�ėpc
ʲ2��̥]��eK�3V�ݽ+*�>i*���w�;I3d gʂ�B@sRHۤ'��f�h�O��M�(�̐-y2i�'j�.�S����ٙJ�]�d�o�qU��#���4/&�z��I!%衹��:�rɛn�r�/+_*�%���9�X��{B���밡��6�s���5I�9o3�m\�r���5��Ru�}aT��2�X�c�����df��O)��{:�]dv#��;���?r��5�/H$��=t��_z���*���wN�֠L�N�R��(%&�Q���u)�����tN��ڃ��ԡw��e�����a�� ��|h�ɑn�_bf���-��f�J�x���tAWn�ݹc�if۝[����ݻ��`��&�/7����3����W�gֶn�6eW
��~�>uR�?;�^��є�g	I)��7r^���tm��c��0�NU�yk�Y��[@�v;��#����X�ˏfS��֨Wu�xTI�y�l���ط#�8lT5�48����z�_[BTOuڬ�|��lmt'��^�.���].k�|���{�`磳{m��Rc���z��3�hv��w#������^[i����FVήpK|	�%E|�ί;K�W�yu�&Z*�ա�^Zoj�w�s�(���|�z�^yԙ������;ú;���/k���mwd|���y^}�㹍q|��EeDgY�t|���$���/�iGEy�j;K�uޜ�Q����\�8�m�o>Y|�u��j8˯�}k��y�%'f\۫"�}������گ#˼�#���;��<{VyE|���f�ׁu�#˾E^yב^w��%y�׾j�+�n���\tS�u�Oh����}��Vw���{ڎ�*}��ފ��z���1��n��۳�Y��y�w�)��/R(�v���/X��mo�h|�^ayZ��9;�qe�>}Z�����"$�	g�Ȉ�<Y���v=u��1���j�@!��Y-J�]�+#�sqے�Y�����l�Kvk7��� B�� �Kݸ�i����wL����[�]s��Ӹ!Lj�_<�����\g�Ru��+7秧nu�]k���ݦۙ٫6���!�;���8�{q��������C	(��)v��x��؋jq���k��a��z˧f�\q�1&�Ý��-λ�e�����k K�@n�������v�7XH������㣄��H��#*v�I�]1�ok2pW�ӹ�n5ɭxM�n�&֯rn,�tk���h�Y,�q�z�i:y^�ˎGV9��]	��3�)�.9ݡ�f�Mݼ��p{g��ۛ�K�a�'h9;'[�3�P-��u�m=�%��n3��F�FNη+�^��]�:��8�O;I��=bӞ�>�:l;&ݘ���V��8��f*͹ϣ��+����U����j��x���m�^�w/��ո8ǵ�����i{$�{fО�=v@�b��R�yK��xD��7=^	�Zi$.w�ncm��;[92��W�Q�fg�����g^X�w9�sR�lsշ������gWFٮv��!ϯC�;,����>��Y�哆J�Qڂؕ��L�PE���W��K�q����v�n�b0�9+c��[�un��74�1\�����a��9r�c:���{�Ѹ���z���v8�Xq�c�(k�Z�M�(�{\
puƖK�pv|hӺ@�^���<����7�v���=������t�G)'.���	�)�"����ts�mڞ��̽�g)���
���^3ٻfn�w' <ϛ�m��;`z�m�"���[y��7>s��qۊGL���ɑ)�s[���9N�.�%���&������:��z��i����^@r��;nf9�n:1SU���&	�4x��;��A�׃c/���3d�u�`�����f�\���	�M?���w�9�d��k{f��t�Źr�5�;\ޚ	��'g`L��X����Mk ���e���/N�X�l�. ��i�pp���g\�x��A�0ウC�p�Yl��ў�:�{q��i;vs��ɶ��ϟ1���j���.y6Ǵaz6;�9�c��vݘ�][[�qvyt��M�[�r�\�n���v�k�Ӻ���6r����=;q6$۶H�X��s�k�;*��c&�N��g���p�N[�林�,lַ�G5�����^����Q�ҏ=��RiFb�Ch��;�E�[Dh�n�\�ϛ+�W��1[3>��ح�iA�҉�����T��ۓ�RZ嵚X�[M����%���C�G+���s�u��^�(�"B�4���H؆�3���"؆զ�`�ߩ��W='���h��X�D3}OjdnIk��3�5�o��q����F��>�GV5��˻�ת��~��{�g�0:��h ������AA(��w)�k�L��&�Ԛ{�e�[��(�:��Ǿ�W�b�g���iF!��h��g��h�����=�}�[�TT��w�{���&�J5�oh��|u����5��0824k.�Ac�!�@3���r�����������~Myﷴ�0##5�y�R-�iF�Ҍ#�>�-��Q���W��^����6��	����z�5h](�����,�h�h���8�GTp&�ή֬i�c�A�����ڭ�&�1D�1A�h��ޤq�l����؆�r��z��O�ky��Ai��׶��A>�w)v�G�ɽ3A�ַ�G5�A�,���X��Ck*�ˇl��n��k�g��$��֕,s
���\ J�X�!�԰E�r}�)�2Z8�1o'��9k,��8g;��U����������V��Y�Za��%���m4F�4Fw�~��CiZj4����c��9ts��%�}֣Ie|ܜ���U%��Ƃ�#G~�}An��	 ���(�"EG�d����S�h#�����}��5cJ5Q�L3��(�k����i���rK\�dϐ�X�C����q���o&?��/0�Q�h�|��cV�6�����,dh"q��<���	;�>������W0C��$".�=H�!�Z�X��c�ܚ�O|Al��u���6�iF�J?�_l�����_k�jS�,_1�s;�m���=�^QlV�4�j4��y��iP�0;��E�[�k.ާǵ����f��;��g���C>��d#��-��S���Ғ�q�~�ϋ	O�i/ɡ���}�,v�A�"H{��9aHA��G37� ������{{�}���}�x��{�R8�(�6����-��F���t�ٽ1��OOnN"�,h�y��PѦ(�1J��_~��Շ���(��iA�����/�q�c#�<�}�jlC�W;>���u�Q�{�H��A��3Ajkz��k�#=�r�3��M(�Q���Zb��CIg_�}���<�t]/���I;R�Lv��WPO_b�$�A�Ow/m]��,_l�
�//;Ϋ��";��>�����pܯ������������4F��fs���+F��(��ܟ}�֚H�}����d*	SŶ��F����}ɽ}���ϸw��q��߽���!ڂ#�G��P��Cj2���"�i-g�^��_u�4ķ��).4��m���54ިE1z��li�4r��q�uϾ�����b�c#wݻ�lCh,q�o=��QPC���w)b����������#3��6P��+V��+�2�(�A�;On������Ż];���n�"lm�y��� G|��[��Ql���(�Q��SJ�A�0�h�y��m�#D����{י�sq�����g��-�m+����'�i�4���o�X5cP��08������h#�D'r��8��ts�H���h#�ﶂ�L�6�/9ܤ[VҍA�s�������6����z�G���}�m�lޘ����n>"�-�+AM�F(�����5m(5d`vv�?��]㙭ex�����@q��?w� �PC�D��w)�h#�roOCv75�H�H#8Ş�]�뻕���}���y�iF�J<�i�Rb�#h��fq�i�4F����w(�.�M׳eJɷ�߯;,����S������Ǥ�x��&z�ܭA�`ݲ�K��Y�x�^e7bG;<���Z�-\-Y�) �}��$��_�Q���������wzަ浭�kc������w���1@>�;��Z�'��i�F��g=7�1�zʤe�6���;�E�i��J0��;�[b�j�*�s}��]�O�m�LmKCv�|��t�duf,���yػ5��MQR������`�(����1�+�6��0��}�X5m(5��3��p��F�Y^q�7{�s���߶���ADv��R-�h#���c�}=$ܚ�O|Al�-�ה[,`F�J5�߹�C#��o'ٴa�(�6��~�-�m��=��QlCiX�i]��kG��;_.�J�h4���q��[z[�Ӛ��dh����!� ���D��&�9����{�p�auw�g�2�w��#�Cj�Q�a����6����WcN:��X�]O�:{U-*���~x�"1F�m�w��4���6z��8��F�'��ﶃ�w�ѯ���#Y�}H�cA��7i�or9�qg����lCbV�Q���(im��o�o���9��ch�Vg�E�X� ��=��(�+�lCy=�Ҡf�����̽�j���\�i�W����Ե0EP��j�Ho��v9��eb�8�$��H���Δ�=]�mz컂�#O;o2�}������}��غ$5���2N��n���+l��ڎ��l���g�}��+t���;N��[h�}%ƨ���>{v0�.n{v.u�8�.B��O�-x�]K��\��`��[n��'=pώ^ѵ�#��M��9ۍ:���ә���q���`�q\=E�e�=��Jw^�g9��n�7Nv��S��L�q˝���7kwm�L]�{���ݶ�vz�\�������;E��΋���<�o��.̶[���}��֛+q����ᑣ�w>��mN1��e���#�O}�e����|�k���t�+��)k�(�60�_�E��(�����rji���MCy+�A�/����{���ӷ�>�x4Ѯ�eմ��`A�����G��AO}�np�%{׾�N��e箑�᠎o#r��Mɧ57��b�v�e�#Q�����h4�1F�,枼^s�����>������l#JF�j?ǹ~�MV�?N�}%�RH�LCIcCF�w���C��q�ӌD$+���1�"8�G;���i�����=}��[W���磻�3<��C`j��Q�/&�˼�>���T�����7��捱D�1F�//Ԏ4��o���~ר���ᑁ5\�x[�q����mT�!���"ݴ��֋����)�ko��ct��ϝ]p�,�ŭ��2��cM�'�#]u���������[ޣ�� ��/e�(�[1�m��m؆(�9��q�6�5�.�}��u�i�L��gh�+aQ�ě����kM$}�����r�UYQ�m�F�f{��8�z��{�k�?l�ϳ}��oDM3$H���mbe�/��P�y���72u=�T���R����T�v�r���R�#�G���`��>�� 7���G?("1��G&{�A�P����g?v�R-�mZiFe�������������-�1F�w�n���54���������h����P�LCb�#Go��-�iF�20>���\�g�X&F�4q���AAPC��#���"ݴϷ�܃�Mɧ57���]Ϩ�x���3w��&�_mRiF�ҍ��즕0�Q�b�������h��1A���Ql_*׺{���/�{��:Ҥ�iD�o+�J�i���;��Kb����Ϛ˷7����1��;�9d9�+�t��V�����F�8L�R���`F�w�v�ƭ���A�����ƾ�?~?n{~�3S�.��\�W��T������[b۲���Η�vЛ�����Ź���������n=�&#�M�}[
M��0��=�G��������s��-������޽�o�m�o�������9u�e"ݍp�[�ZR�ַ�G5� ��{�]�C5�k��罿}��w��V��vbiS���9Y��-��#Dh�Q3;��-��F��*��#�<�ϸ��/�,�'߬�����F��d�lL�_��v�A�"H���\" ��A{�K����9{ҥ��;�;�iX��YL�J.�賖�ˋ}�����Y�+|f�&'ѩ��r]���_����++��k���v������5]���mXҍ@iFa���Ql,b���z�B9U�[�!�����g�i.�{\_��|�WȦ!�y0���h��iA��6�~�p��4Ƃ<���}�����3�< ���gԋv4��H��m�9��A�Xžs��l��j(����}Z��k����OZ�F�D;~���m�4F(���E�ZaQ5Q5L�ԃl	�/ә�����޶i�jl��ޤ�f��mxW��f�u�:�OLq�Nγ�|]�$��������=hss�6��|�#�1@;���r��"8�G3Y︃l���z<v�{{�����<��k�w�E�m(�M(�0�޿Ql-�4g��c�ִ������#�4G�y�4Sa��r_��y�j��1��ﮋ�!��3�_�[�F�8�7����m�|PD���:��GSG���UH�݆��&��jk[ޣ��Fq�;yt[,`F�J5�Lˣ�J�A�0�Q�n��}G�ʯ���|� ������-�m+CQ��'}t�Lwo����{qк��q w�#������|XE���zo���D	 ���bݍp�g��6�Ȇj3��}H��>�>}Am�E~���7J��[W���-���9�C��Z���CKݢ�^r�v>sb�Jov<�n�n2�yKα��^u�]˽�f����$��k��A�~���[LQ�w�;��޵�=o{�[���~�h:4S؆��ߩi}��}��d�_08������`[#Ab����m�|�$Q�{�E�h#�;z�Z������Y�[>�>��iEH�X�h�q�Ր��8z��Z��u�"�k��������z&��� �1�|���6�iF�4��w�G�L"b�Ch�s����!�Ho��=�>sr�������E�ZaPj4�j<��Iq�������捷�[�#���/�;h ��w��wU������}\�(���n4��r��l���Cj&w9�մ�Q�o�u������j{2��y�4C>�x;Tp�Jٟ-�����k�_c��y���M[JF�����P��^��:����Ch<48�{.�p�!�"@��s�R-�n���U_u����U� ��>�;݃�|�l�yZ�{��ƶ4�Q4�ɗt�l8�D�"�s�q�cDh�D`g��Q�+���|~�t8���iF���=Iq�i#u���"-Uȭ�Ŷ��C�g���;h"q���}�=�r��]�ů��;ͺ���Ѡ���x�l�2�g���H����J0=��(�A#��x�՟�K�;��r�N:3I�lf�z�3�%�}�i?~g��g�Ot�N���VcH��[���]%�|����S{>*�N�;�	$��V�����d��9�+F�;<�ь�ю�p�����.����D��m���4{]�;��Crdָ1��NSt�\�ni�n��m§q��vŇ[���C��Nmn����Ck��qöK�8vv���$|Uک�.z�ٺ,�Uq�y�u�ۮT��]�k�g�-���.���kvy���a�Bsƚ�c��;�wnh�]�v��ے{�7<n&��j�ӱ��qfD�X;;�N��0dw�Psw=s`�:U���	y�'�󅄄��Y�>C_&�o=�b�0�Q�h�ݿ������6//��؆�L��������;��R*� ���z��q��G|7�މ�57��b�s�E�;n�5�����Pt�:��o�Ay՞�������Y\��WwD*�j�T:��L
~�Ɂ@P�n�ύ�2:��{Ҙ �~�Ѥ����~'��
�#J���%�>N�6�9��T3�s�> ��:n��'��]Qͫ�����V	����2+���ࣗ�d���m� 
����D���;u���~��n�O�s�\�{Ͼ�m��s�͵;]��5Hm���r��`քz�]=W)͠�Ԗ'��������Y��,��z6( �O& ����<;԰w�}Ͷ� 9�́[|NZܱ�&���ӻ���]޴��r��2]�}��һ�_��e��'���"R�
v�5����QY�ʜjfĪ��OR��uO*�h�-�R���MO�_{��$ �}�p�c9�~�l����4ϳA�{�Xͭ۽d�`�	X��6�o��@Tޘ�
=5�'�R	/N߈��L�I#�v>V�uUwDUP�� |�3��2�(�� �~��N���L@�t�q���gb�<�'�U���o�g9�Z�
�,���=�|��m�~�׵z~����@��=�����ﮊ߽��15�g}%ͼ�i�	�Z�a>uƲ؏8,���/mN;Bq恋q�g.�i�9o����W�z'/.�7c����� {ދ�> {�"t��� �6,�<Z���{�X�g�B���+G��&�����������H$'^~'ޝ۠���WȫW�x�ry�j		-nX��}�֟ɴ���l|�W��^u����m����m╁�=��%\�T�qʾδ�k�ݒo37��[)�N���sgAOK������Q��]ySS�m�f�4.��+n�(vr2:�|�r[۲�޵a�gz��)W��+�y�([�
�}�;��j��]���a��G�.�WwL��3+��3ۇpw�do!�+a�b=�s�{UJ�`�oXU���/����ō�T����ʕ��fsf�U+v�u������Z���\;Q��M�ޫ��饢o��[�zP��l�:�,�YF8T3u�wW0��B_&j��|�t�t��k�۫���u�IV,�BY�2Vv@;�Ѳ)V�Ùc0��(m���:,�ՙ���eq�q��9	����:ˉ�H)�5��u��`x�RBNT)�����b��Va�w
��9{b����;h�������n:��P��͕G����5�9� ˢ�Ac�����t�鵘X��6d�fǩ\�����F=��;o���ӼL��D#��󩊷s�a�Xwg1�5��ݛ�ƞ��͋J�e�E"Y��7ƶmK��5��P�\WP0��6賙>+r�4F���>�7�ڏR�0o�<��on�U�²��cpޅ��X���1k�3:��1��n)�2��VfP���U��=��]X��$0��sA�[Y2�5^��2jꭖ.pK3�&:S���`g�ս3
��t��6��k�`�Y�ykb(s{�	��L��Yo~7n�N��ҁ9f�2�a�j�����5�΃FdK'L��]��q|@Se� P�������+��8⭾�e�m8�'o5o�yw��ue�+�nｭ�'ͱ���������v�Ӻ��ȭ�{������5���_;��|ץ�qf����.mEc7e�v6�{l��gcݍ�ϣ�ܝm�ܝ��avv]y�iݝ��h�3-�}�{����>o�Cl���(��q�۳J��g_}�}3���(�;<�˳��ڶ�i5��>��=��9�v���󤓣�,�.��N��Y�GE�ڳ�:���M�����ۆ�]�y��9;�+*��%�m�l�
5�/{s�u��uy7l���]��<�,���Z��w����e��W�����X>�+����r-,����6�I�<�<m���zfe�swf�f�;,�.����tg$���z_2::���y�Ew������󵂌olM��-�?	$��|�?��{�����S���~��Q5�b������c��i�Bv�e :zF�)v�4����+��~�I��z�U�J�A���@|�r�>ó<�R� #o���7B��~n�>��������d�rcu�66c5؜�{k$��y�B&�f�n���('9�uIAªK*�}�E�T����b��>]���Ӛ�ӧ���ʔ+�R_yll
�YWw���g�n©�Ǜ�3��R��`PWF�$�{��C��v+'E�ǟu�:/h�hR�"�����g�@#:{�~ �&��s%��~Zk^$wsD��o�`V� � a�n�,|+��������5W�%�ɺ~$����h$ޝ�K�
�#1D��7U�,�:��n�]`D�eK���of�O1��������S-�T��J�X�Y.2L�]�ݷw7��ַO���W�� @��&��{|��'�rL5�OO[�"���}�n�]Z#8��٭�/k�L�M�T���N���{�*�[%E�F&�Gh��k��J�Ϣ������ƶ�OQ��h�˛��������9�d�����3H?[�X��[���,�-q�V�����.Ly�ڼB�V9�v�P��� ����Ns��ܹ�([�P�~���+��e������ /,a��U7ѷ@����P�"B�V-:����BA9�&���},r��v��8m�z�5w�-^�
4�y������	���
�ԃRA}�s��~��
7H[[�]���ͼ�c��<��	��O��h�H�۟` ��ٺy�l�Y�)�[����j�g�}ĮQ�I-��nǺu��f�=��ʸ�Z�JhвN����:���{��j�����EOQ�?��}��mVi���ޫP��xi��rb�7&tY�v�Ӵ�/����m���l���Í=`�lT����s��ő�Y����<v��ӵ�֬��v�j��%§��Н^�=l�5뎡�<^.s�63{wO9�'mF�X��{���g/m���燞������-�>8�ݹ�7r�l���-��8����)�q���C�<�q��ގ2F�0r�rL���V*ő��Ӯ8ԨV�]!װZ6]�S��V��������.�}u��bm�G9�0�K�lђ9��<�����Ѥ�:{s�?y[��7b�&�'������d�`3պ*d��$	��6�A ?f�C��F�qW���vo���T������]�����~t�W�����j��פ����>#��7A"VXHm�iX�A*G=�n���{B.z�?'������'�N��旞��ޮ^> �$�b��g�.X�vʼ9v�+u�J��D�j�y:dfvkS�ۏ����i�~$�9�! �W7ͳy��_-���}�{n�EGiT�0����Z�+�^2��v��;��v��\1v�i�U���{��n�rR�<[��$�}�s�BI5D�7�2{C.��y9ٵ��|jk�ku�I	����$҂,#��y��X7��d���~�H�O,~����@�z��-���7N�=7{.�jR��&1���l���
Y�ϭ�Yx�ؤM�u��Pa?��Ԅ�7U��!$$��^]ڑ����9�B��r�y3�;���uc�ƅذA�B�l�'l�	$�5s�6@4O7�j��D�=���]�t�BM��n�5��F�T��ɘ�L�����|�t����$�I3H�l{��K���PY�og`׃(���ݒ|I�c�/.Ŝ���e�[ͶM{ޏ��b�� � ����w���> S9�Ń^���V ۮ��߽K�;2i�dmB�+.�ۜ��&���A˒b�ɣ�xm�ټ���n��M���~��r1�)d����wx��@�w�d�I?oF�8�g���E������L�s*��� �R<	�LȖC~�x�<��g%�I$m��tI�I�wF�ye�T��m�.��w߀J��|px���3��f,�@���3 k�ɓܜn��X���;V�n�YY�)���[|�_8���YGT��-J��wJ�*C�^�*�j��1��w�.z��Ù�H�GY�U?�}�}�%��|�7���{����w���<u��U4�o1"{|������{Ǣ����� ?�����d� 5�@2M{��ڵ��\u� 3=�������8Ud�×m�W�`}��ʇ;��Ƭy
rO�?��d�+y�l�I�G� ����9�b�[x�,�g�2��ߛPu���a�\v��Y��sc����#��������:�M�>4�Ͷ@4Mw?6�4I������-���W3W7� �"����:��e�GT�I�=�g�������,5���z�I��35%�Hzv���D��(iv�5e�G4j_;��#y�,Ye�^[�٢@����O�I'v\��{5�b >���X1 ������ןuq��8 �e1��^��"b^mk&�Ě&��t��Ol�$$�&�c�9�/������T�̩t��G�67��u���6��ΕcFt�G��챙�[Eg#z�ez!�
3n��x�T�5�#�k����|���!�w�g��~_��WSL�[�~��s`�@�}��#u��R����s��#s[N��w�� ��{��T0��ս�:������V�y�x5�ϱ`'�q���m��և���M���*�_����H�Ud�����ŘI?۽�Bh�Ǿh�Klv�=����뺣V�n��?Ool����ne�-v2G����i�ǿW�|G�-�6� {���D�$�k��@+�\���j��z��jI��I��s���P�@�}��I��;i!^�޻
OmļD�oϻ�I$E��hԀv:�B�j�A���w9�k��@	�{���4I��?{�h�[�-��k����w3`)�Ƣ�	+��g��?6ɢO��oGM��}�1�&s��|�$\雨��H��sO��Ւ�a��1�R���*�Ά���~�ׁ��LS��}62�F�V鷻��T���5N��w�V�:�%�4�.��}���K[ٵ��]�*��ܬd�ӈ�e*�����x_&u��zS��GV���v덀2S�; m����n�3�����ϓ����y��#�᱌�y���^��'kv,g�d��Mqdm�eG7�g;#n���c��G/����\=�S����[p�:����؛�����h�����\&����U�k���c������P�j��f7�Q�������۵��e�>v��){M�zSF�6r�O�4�%#�}���B���p����c��$�Μ��h{�ZtN�j6e���I�&�&��4�U�N -r�`)��%�)��?6���>0u��Ӟ�Ȕ@߻ۚ�(=#��PJ�d$��K�Vt���v��*N�c$y0Z�s3� >���� [��&��ox�	 ����W�/��[;�]	X.��e��v���o����xn�"	��\y�RI$�2G��/���=��4�L�+�������T.Ŝ9F��&����$�3ӵʨ}�}Bk��Q&��2I&���kl�I�Ol��r�C��gw�������O�k�M@��vO^�JQ��Ng�L<���k�v��_���9�.��)�!sY��o-��Ř {���>%l��RZl��5x��S �MN����ގ�)]L%3���66��~�}���]ݤ7dֿb2_c�Яk΂��A��֒IlgmG���c]kn��!�T�
�7�eǘ�F�rdg5?!$�V�o�y#g�視��L���$�N��K�V��^��)��sj���Vǘ�/]�%��~����*�j�o	ВI;p�Izz=�a�dB壈���-L��ȽG��x�(��"�=�$J��rK�C����yf��Q"�w�d�� ���Yxp]�=�ͰI�����oV��5��O�M}�v�(�D�I��
���t��ߞm>�`����!*���[T��5��U�R�R ��;%�	��˝�Z�cuN@�y��0@|�{����|s}77䮇�-���a��F��IN����
qo�S�����b3���$&?X2Z{Ew��Ԓ	/zG��$��g�n�5*<�(>�Ʌ��B��u��%�L�g3����k0 ����/:���u�7(8DLٻq�yKV"1��n�h:��qϛ�%��x���F��w����ͦ{kg��		}�{��$�$�g~��H�"�����{5���U�G,y��w��K=���6�C�I<��h�]�I�I�A�=n��]���ݸ7��s����Elpv�@�.!k��b�I������^�K�;bzH���o��I5���A$�k}��6���yT]���n*\t�ݱ�>�g�q�Z�g�����gV�+�����&��BH�k�Low����I ��盩�A�L�H�����z��o������`sK/H�U",n�d
�{�uQ.��H����禷*TI$��Mi�~$V��6A����}n�ݠ�߆�֙	GL�_wy��?h���t� y��yqp����/ٹ;���D���=�E|�?I��M��@��k����o�t���=E=��ѩ|�HG险 ���<��\R��*�o;�߱���2��,��Xu�њ����{z�<��o�#^J�t�@�UJ�ĩ���,�j�s_^v<j��ߟ5�}��Wdx$���E
����=��]
B�$
�)�{Ř*$�ۭ��#�"�w{���&Ni�II|���5_{Ѿ�	S�[Y=C�����6s�)�qb�,aN7%���Ɓ��[����������	}��v+c���
�|�{;p�H��陠$�Kލ�pH�IW���"��!MѨ��C��w�HK9v�ddjJ����s;��s��7�_ׯ&�g}��@��J��}��H$�~Bt�(�����e�J����F��$z�'ۤ�ލ�I7hv�n�{�y�$J7��W�{�=�S��rET�P��w;��y����H^�߷W�/�]$}�_$��绞NM�h�:� W��ņ��y���Ddv��$�!4I&�v��#D�w��[����Ny�E����d�$�v��I�$�S}��7T)�����KTb��pX$ՎSeNJfk�z(PO��!����^°.�3��  "�������޸Yy�Z�Ѽ�Q��)�T-m��;��'�����w�R������B�I��i���XE�3T������l�q���'ۆ�X��0�r]Pu�������;]�TMc�n�� U�E����Ħty��6�Tˊ�-���;"�Zvm���T�����I��Qk��ڪql��Q�<n��Wϱ�RN���pm˪e������[n��/5�_<v�����6��P`,�Ƶ��R�T�,=�:�rUb��0�#��2�����-K�P�*�����b4����Sr�ڷC+-��s�uf�Jp��ZU��g۫:�6�PHuK'��ս���'�dm�i�N�f3�8mL��fK�A+ڛ��v�2ĔE��]��:��Z�T|�&�[�l�[�\N�n�F�}��k��oKwgL�
�q軝�S�	��,X.�X*S9�i�B���͗E�`	���f�}oWw��d�ξ��&T��nRw&��b�\�u���O�jmq9����uk:�"��J�͋;A���� k+o�2��n�4���b�᷵r�gTnڙ٭�����u��;5��`��ʥ��ÕZښ�[����uܙq;nj�WQm��5�zӥ��=*�3!��"��ۯ�M��p�(,j�̼���J5���,�Ѳ�5�6�Cw�vdf�Ҧ��+[v%X�2�� k���M�u�/�O�>F�a�6i����m�g��q��}��2�׵o5�m�3kt�����|��i���=h�����=�eY��Q!�n��㭭ݨ6�Y坕6�y�u��+:�Gk����w��o���p�a�'v<��N}ø/*��3�6��������=m�Y���̗˾{���m$����:���.�g�y�8�̻���ޓl�ȳ�#Z�Iok���Y��wz�ﾵ��]gy|�kwEe�g޴f���^��tMj�^��&ם��|�/m/�yps�;-8Ĺ,����󬽚��m�y�e�s6lוxxE���<ݗY�׭�O m���l�y9o�W���޽�����Ӄ�,\�h�ÓmJn��i�n�Ƕ�K,���[ݒo�o>���oQ�y�9��[#k�e����6���)��e�÷gFy��P�gs������.�v���C�Z'vj	ݶ�zһͻqus��i2��V:yN3c�̥�N��{��&I�&;:8�d���:�[8#�v�5ɍpݽ^7+����t�����)�m@�c�s�ۚ���v.��&x�Ui�}v�X�.[�M�IӬ�oY֎x�x۠�=[n�H�4����걺�<e-k������ݯkj��� YR҄bS��:�O����v����A�,G�t��`���ǌ�8ܥ�<m��v�����ݹ�y(:��th�:�=��mz�k7<����s�����v���ێ����b��^�Ł$�O`�v����"�;g���ќ����: x+�E�7�\�ku�]��0N�;%�#�i���s:�WUq������n�qA=�7��.�!�qٹ��^v3jϣ�v��v���#�yNӮx�{)�K휆q�kr�Z덺ܳ�ŷb�cO/N��e郧����p�z��5q��6��S��ô��o0��]�Q.'�G^���ԝ�s㳒;<̹���=�<����v��9�q��S�{BP��A��(!G!l���4�����u�(fyn��2r�q�9�p����v�.d�+�9Lw
��U�]=2�����Y� =���'8�Br�*/C�qbyUlI�X�"���+�o7sCP�x��G���>=yh"�y��v���Lۉ�Û��Z��n^R�Ge�:��
Fqx�9)p��K�N̅=A��ιȏ����`�A�B��vcy�֩�rX3m
���T��'\����0�tq��l��h�O;Wf�9�q8�ŀ������]�%9��1��g��{���X6۵v��Yk����s94[���#��Q]���s�q��\�k[���d"�q������ǰ{.���n�]�p�{k��ރ=�x��0/c{��ˊ㗇�*''
�l��۴�n����㊱Y���k���_����#���ݣGDǨ�`�����,f*�t�N"��n	�����{=��7^-��\�qc�5�Hc�< �y�ϸ�#�&�� ;��˹����a�]&�����=]��	��(���Z!�7N�n�%��5�28��fꗇ�wf
];q]-��~>� ���n��c��#��gn�s�pF�҇lyh4�g�����	���Ѯx�u�hz6�i���ڊ�fڮx��\0W7��h�E׮x/8Ri3������m�it����h���Ѫ$	�9ϡ4HM��ɩ�yŒ��)��8�"jo>�h�r+c���
���������)�$<[M I?T�>�|I�MQ��րd ='һ�n�g�t��	�F]�%T&<;{���� Y�sX�l�4o�1^AH�y |�I5D���� �k9�f}��-W�,���U�>
��(�i˒�$�t�� J��:$tzM��c��M'�I;������Z!TE�@C3�tjI�s�z��U���j�ΐI���k2N�Nlb���&fج�C�6:F�4*��U�η���7Re�b�wQc&M�F� �ρ*�;]�E���ߏ���%F��wH�Ht�7H h�北�n�cwe�V/d��$���{��{7�P�Gd$
����p�qK�v�x�;�h������;%-�	�uu���|�2���_q�ܪ�Ļ�S�\S�hUV)�>��o@�����N;�m�����}��Kc�P��A${����I/�?�n�$�&�9x$�{^owٽ*���B�:��=��`؃���}�;b~�z�*�ۙ�M��$���<�a�I�F`�qF��!���<�O���$�M�l�)����z%	�;�V��M�7<뽸 �Sz�i�]�T\����GU�>A_�ͣ� {{��Cpj� �I�����`��t�$��t��2�]���sK�[�\�l��QJ�m����_n��箞5th��d7[�
��v�����x���H(ꆼi-�l��$����h��tn��C}ޘ�t5�����͢~��<ρ�"�Xlߤ�!?Q*9��&�//]vjM�I��P�玉4I���O�n
LJ�����r���ż޻\��;d%����,d�'�������xg����Ⳗ,�;|�ͫ���:����cZ�(i�;;� �b�,�r��-��g����G��xaa��F��-`!
k=ϫ	"��9�Q��{w{��U��H�uj��o;�����������^��J{ӻ�$JC_��'�t�a�vk w�&�"b	��M�������t�(�}�M�Z�bqf�h/=i�~'�>$�iﵡ��-��h��t��ZH�J�Q�V]��vv_B�X�oV�@.c��Ӯ�}�O��u�Yb�VϨ�[�t� OwG!$�i�&O4��{}�~���ᨗ6� �ot�Q'�f�[�HF��`��w1`߮��������A$���I|�k������[���٥��g��N�9SE�Gc�|Oo�����,�y�X |�xU�c���jߨ�I�s� ���=����z텿
2+g����۳�z�y3�F�+y��"I@��ВH����4=W�D\Cՙ�o@n�<=�PX*(�*A��7Y�1b=�Չ|���˹�;���A)��j[8��z��~)����K�Oox���m�3��]��'szU����ˈ\������<��=��1H$��k�36t��$�$!��tD��{��]�����'��#\"v{���;Qێ�$Jkyvz��p����J�Ռ���}�!K%�p����$�)��6I$�'�4��Z�\�]��o��I�Cd��R������.�*������x�|��o-z6	�Hl�3BD��{��ڊ	h�.�^��V��{=�5��q12��P�!k^��RB>��JJ�A��:��N�]�?�_'I�N��C����7�Y 励����b�y�J��xw�&���$�I���:$�L��o�c���������`o{�l-�(Q�X�^R6�j��~�Źׄ^��KV衑2H�Q�h������L��*�����e���70��ο1M]�--dv~����r����ˬ.�-�z&�KcA��wU*�ꨲ��p�y�]�`���މ�6���q�d�"ʽ���gm�\�<\X���q���U#%B�UH(��*�x��K�%uôk�J��}=�n�;�|
xKg�ۚ�J*���Ŏzn�n�[�1�tk��l��[�&L3��9�ާs=\h厺�Ҧ	�lX�n66�ܹ-�]�;)��p�a�O'�Ϲ�ڣb��5b��$m�;Z�Ě5e�l3<u��y�E�)u<zx�8s�n���8��7��ad�������\���?!{��f  ��wZ� K��wrZK6d�-���4j)$��n�׬�EB��[���w���޸+m	��T/3s@ԂH$��M��"WM�I	5D�u<�)?r�2f!����	e�U0�Z���1����sl����������$�#��n��K��d��ܬ�d�vF��X�n�|��W��k$�1ə�"d��{��/��1�ɯ_�� ���m�oVp���X��_��bI����]ǜ��0f��.IĒ��$�'���I5��h{<�^:�����×����E�����Ƚ콱�rGǓ�����\<��t�k���M��߿gm���+�$
�{���3�����I��3M�#=܇3I�m�~$����{��z�5%-���#]�޹�G�G1|�e����l�=�*{3sa-�t�]��/�9�4`˰郑��n�:i��o��yY�:��u[�:#�n�����F;��>��6�����$���}��I�7u���i�f����V����BH�Ke�a����� [���4I�qф�ZC�q6�+���J?s���	 �������e	f�UYj�L0<��߹�л'6 {��{�I��7	ВC�=���W���i�ohs]���5wڬp
�(ao�^O��'�jwk��/gIt�>㶢I\���K�'���QI ��{�G��v������V���ЎG$Q>�k�۬�΍�k��j���EnÀ������d�"�^Fs^���� �s��` �֝�P&��QF<�צ� �^����O�]�3>���,7�5�"L�߰����
�w-���J	 _��'RHyɻ��`�㳒��I^o=�%���F�j�V���ow�m����w3 ?�
U��dy��N@�y
����o9������͞��-.pa�C|�<O"��[l��{,�hZxP��7i&��}Wï�6�$�7�W�m����F|�w��n�o�P�J�[n��=���>�X����ۿ$H��5�_rno� �o��n�L��t��g���zYC���l�Z��/g��0��~���w��x��H��愗�$<���	7��{䠣���0R�cHlgC��su������FA�����hrk��<�� ������뱸�:'N��_wy�	$��&���%7�����3z�ŏ�ټ�g�����woKĄ��")Lχ�:H@���e`�*������#�&愉A�7��$�ɵ�W�9�Zc��sO�v�\�J�(VQ����,��@���BI?Q7eK�ˎ��kjQ ^����s��7������YmVG�2�:5����&zr�� V/D�ğ�?7���	$��v�����V�<�o���y	�J�:�l~�Z�e�z��O�3�)[�������o]]޶N�S6MJ�����(�"�����-�׹=�I	d|D����Ò۫N��PVl����_��}ÒH��I�EW��ݒ;�s<@$�q��I$�~�t`��\W�����D�V	�@M�&Z>�M���6���=���V-آ���߿�������b�=�.�=�0@ ��f�� $���i�4����hW�Z2ę�ݛ�@r�κ���%S0W��b����E}�}�=\��$�8���A��tL��_��D��e�!7`U�vo+`䲘���-��]�{��@�B��}[�{^0�+���w�/�H?I���e$U��#"����w�K�)�ض�K����H$�/�n�$���۴�X��%t�}��m��*���U�����s����/{�����=�����X�^���rD�q��E|��&�˂��;�Y%MBn��\����r�,�rÇqnk١�^	[xv�U�n��b����^j��H�)��p��8]gH�aS��꯾>̭M;��ǭ�X�A��c==�;Tn�V.j'\w�^�������qFGy�i�yv�Âx�]V�]d�hͮ�z�S��H�l�m�ۂ-�f^���Y�6�\=���!m��<��ݷ�׎��<��=t�7!^�r�ng���^��E�S��vK2���r�"��'�[�㣷 qa;�9�\�&�線V���#�:.xSF�׮8���aь��K�=�`�FMd���=!=IŘ7P���~��~!+r�3_�׾����D��3u �(�&� �/\���J3|�I����$��{�n�N�hR�P�������uf=�\[�qӽ����_��ssRA$~�p�J�9���v��:�.˹�8�(IA�5�~h2@���٢I-<��~o��� �^����>���Y��� J�&���f��t��60v�ΰ��!�� �$�'���4�?=ݭ����}�p���>���ܡ��؜Ty���I� o����_Y/ޕ���:8�BH$�$��I����H�P�g�ƽ�/��[$m��V`X�Ya ��:�g8'�h��vp����xY���������5I���!����$9黤��ý$�$�5ף��f���L�D�S����-X��]��i�w˶O�$�z�b�"���{d��iED�����p�݂�ysj�Zq�Uo����N��&fΣ���HXL����I�*�2X�Ǜu+��_���z���PIOM�I��I��%��RS���7cչ�jC�V��B����0�W��|� o��s{	 ��:�zFy����"D��$�'@^�{�� �.N��qKF�cS��z�+f	�ɹ���~���Cޏ@�A$��;�$���z��3ҷ�)��T'�~�f,��=y�%N����{7�!$��k�u v%�����l�D���:^��q=�H&|��-������_O�����\l�Be��+p��x�6pYz����n��?UIKmr�o��q��8����ۺ�_$��9 �I�7��Z�����G�zk1��I57�d�~�z����W+��.w���� �ցN�������IO7��$�I3��~�RC���P�����d��]g;�WF��}v3-'��wt`N�n�H�Iu��ۊ�^���1�����ʛ�����St�Rm�P�ġ�W�M]ӭĠjUg��I�T�e��[��m[�s�H��z��9Ɔi;�m�ekU`Y��&�[6�f����c�´!t���v^���	��-�6��H�U"c�*��9��a�!
'34)+��#���)U[b�>�2X�3]vk/$�7�w:��nf�P$�Ie�UۮաoGG^t��;yC�VR�5�ٛm�uzi����h��]B�n���s�,�2e�}�t�Yqg�A탻���m=�$�+\^��e�c�Ct����]Tq��)��: ���<={V֦Gv��"�J�m�p��6��2ɽ��a�Ls�zs-J�C�|q藹C�J�]��k*]S��P\lgn��A�b����Ik�Vr.���ϦC�Cr�V�u>o&�7{v/d�g&�ܽ�M"$��莳 ��VQ�8U��6��I�����諸(+�7����Aa�Gco:��c�9�[y�������y�}�y���]b#-:O�� j�!z�A�ce>��r�%�\S�)mke�9Cl�+(==���<��;Vڥ��@۱�����+�*��k��3e�M��*��A$C���䫺մ(#V��3�'jE��q��zV%հ�TS&�iuMƔn����00Q�t4c)��M��:��DQ㵚`]+a�pM���X�\���^^��lW��{o}r��8Qڸ0jaK��yv&=	��O�$��I��?#���c����<�{i�������I�fk;��wg6��8�8�;8�y��qY�m�-9:�(�Z��2m���m�[����Vv�id^���wY��:2�&lnl��k4���"98:sۖ,�΍�����nu������*�Ţ�7�{�dƻY�ÊrK�� �i�h���^I�l��̴$����Dt&�`�-�G
ZV:GG�G�hr%#���8�,�3!m�q�ͭ����mو���9	�a<�G/jÙ��m����Y�3.ŷd�E�ۛF�[5��i%6��NrP��4L���-�� 9fqA8�f	N2���
�I�7s��m��@����"�}� -��?$���7�O�g�{��S�B��mb�g���{SK��]�t�=��o`�@|�w�ˀ k��qk�[��"N�o#�䔫ج��ث����V};tb% ��&�7jeݳ��^lMs�$�y���$�Iow�D������w��L�{��5j�ARv��mO i�4v��7\�E�-���u��o�z�n3�߿����R��Z^2�9��`����-�I4=��2|+k���g��$$�~<=��Z]�>eh�ҧ6�u��0{�����'������a4H�X�I�׻��8���1N��}����k|�ϩU��UM\G]�r����s�� {4/{��[ײ���OĚ5��m��{��f�7�Ij�H����ݚ"�~r��߉4M\�H?�����h ��Ȩ��y�͐�r9F�w�n��{*v����]��6�US�6�s�FNHD��x�-߽4sά~���Z�/(��.�c�A�]���$����y�Ki�XR[-�W���Y�9����˻9�jt6��l���D���O�MQ$׻�� �'}�dț�~|ek���cm�Ρ�t����z�u[�n;]�jz��(l�l��	��Z�qrQ�[5��z7L�I57��d�I�t�'��d˳A���G�&a=�Dy���s�U�n�U�n����>��<�}���XiOD� ��i�@{��7���g���M��A��ꗳ*Ȫ��`дs~H^N�'R��}Ȕ�3���Q{�i �Bz=�D�=#}��Hz��E�J�Ջ[z��^�ҭ��x�II!��	zF�x$�I ��=M�u��k�5��4����]�V}v3-�G���D�I ��0��u7l$�9�7	Ԑ~��pI$�~黫��p�M�}���@�Ǹ񓵚�7r]n��i�/@�ۻ�E,W� 3�!��6�9T���Æ/3���> Sԧ�uApKU\w&C���{mv�n�m��q7k�Mvݣ1p�r;v�sLMس���pF;�ںԦQx0\&�u���n�nx���mi��.������\ǟnqj�;y��ή�K����y�p�n�n�Gnݘsi��t	��nu�;f�h�6V�v�p��j��=���R�t�^���۱�9=��sK��{��3BF�yw3Y�R�Ŷ�t�7��m����=�&ѻ	g�7s�:�l�#gF��"U{ή��`��X���]��%���_$��M�y���Raʮ��ow�E�n7��&��P�AVO��P�N���[#�N�>Ą� �%$�~��rI"�f�E%+�K�Q}��������4X\~���5�96@4J:����z0a�h�H��}��H ��w�H_M�"�]�+,6Mb�޾}���.g<t�L�c�P��?ho�Zd�M�o?x��u��V��������szpj�Y%%Tˋ�v�3�����Y��l��Y� מ�w�H���F��Dz9�����z�ߍ^	��nJӭ0�υ"qEu�Ƈ�.�$�l�V�\�U��ƻMu�|�~x����s. vNlz�$���6I$�Cӹ����r�C��V�� �?��h8r�}U�e���pā{��}�߃1w��lN�(Wg�Τ������F4����u����@P��&]r��q�_�vHw_+ɞ�Wqת�2���j�
��� �����W!$RG��ܮ)$�}�9���+�׸w;���\k�6 ��Kn`����6���Y� �	���c��=���	$�G����H{�s�4��8Z��B��=s��ִvf��OD�絋 {�{��l�w�I~������5���i'��^S��p�֝V<ρ\��X��{{ͨq�D)�k�H�H���I�קsl�S~�����lwb���D���n����B��=!6ǵ�t]�ج�ݳ�u�.�:��d�����
ʭ���v�^���w~�}���$�5P�����_�kT�t�4H���l���>�/2��a̶����b|M+�9�W�ލ:d�'�M	=�&�M����&�Rl���v���~Լ�I1W��l����;�a���{�� ���(������V�)��/8dX*6f�D;j𼚹�����سn�U����ʲ���ޥ��� v��q���2��[ЫK� �nL��c�1���lw�=Ϲ�a$$g�=\F��컻o|��]�������_g��S����N%P$H�ݣu�K�����$��h�i�pu�Ű��,��L��///3'	��>jl�B~$�5�ܐ�W���x�D\@9��5� �]�{�� s��i�F��{뮑Kk�ȝR��v�5��M��o���|Վ mt�����L�A�M�����nIcN��$
�o3 >���D��?�sL����y+��A�Q�g�1}�>@s���{A�f�2�Z�T������K �/y�c���y���$���(�k}�� �����O8���\�0���30Xs-&o{�AȔ������B��n�X���7}�2I&��� |k}��2t� u`���-�w_�}�{L�O>9&�6�����$I �{�%!�shS��Z�����c��ЁE���zZnz�T�_A.u�՜r�kb���a��T�.U*;ȐX�+(e���>������i�W�`��|Kn`���t����5&�le�JŹ�4����w�H$��n�($G���@��������ԫ���Q��S��]VŽv熽��Z���}Ch��5T�;3�|���`�B����{��	 ��L�H$�H{��ߒ��}xC�ޚ��J$�'�[�懖��8�+�غ8�H^l�Б0��~=CE�S��w��  ����k �{��b��T�q{���^r]w���ޛ	U�ʜ�f�H�I�w*HK�����]�����I���	 �stS�ƬU�ZB��fhT�')��g�!^�%;�ͤ	$�����ĒH�����D���n�G�٦I�������xI�����VU�А��n��%�^s^���Z��~���H��	ВH��5��z>�䘉�x��U,��):�`��{�݅+�Z��*Yrf$-��i�luE��X�r�ֻ�K ����7�,Vp�n+6�Z�ۛ//2;�u~�(�잎�?��V��&����cp�l۬'�]��݋��\2����Å����7�`�=ku{[�R����c7�s�.
T=.m��kn�g1���	ٲM��C=�+n��<5%��R���PT�J�V-�������m��۴g�LHv힞9�ۤ:�z�f�s��$ێ��7n��"NȈv�L��1�ˋ�ӎ�{��e�Cvm�m�րvdn�=�$�`�ss���Aomp�V&�\��=�5�������!��-�jk���`�-�Ř�I|'���Hb�;��o���uW�6������Uwv
��uz�>�K�&f����	��rH���f  ��y&I�{ݱ�I�I���}�:�D�&�x��rR��Ǚ�+��,���v9	$�7sӥ�=�^����z��I��Ѩ��Bz>�'��/�
�U��Y�v�����0�� t (����I��$}�O$C�y���G�;�x$�A����zy�ݮ���Kf���y����v��%����X�P�F�&�?O{���H|��恩ۨvh=�Ǯ[���%Ӹݱ�9�#��u��+�5wV�R��N�[+hݲ2�}��UqKi\��=�.�vf��K�wo��I5���)�C�^�&���d ~��I �j����Ы-�R�1#��ϴ)��}{�k���Rj��Hˠ�ƶ���7!ޓݮ_�q�[�~��k,[��e
��`�3u�~v��orC�Y<%���tyʅ
?Ϫ���|������B@?v�� �\h�{/j�Z����K����KIm�(��z�>�Ȓa���_$���j��杼H	D���d� 4{b�>]��nJQX�>u���^�`�́�s}�n�I �/��hI�C��]�C�ţ l 6��d���%
˼8N`̫���]��4M{���s�S�.���Е�7�wI�H'���I@!������{�mw�3��t\ke��"�Tr��Ȉ��7b99Υ^���"�g7����?���o��-LT�f��9�{x��=�k0I������I�6�1�=�qi�C��7�� �{�f`n��)-u���&��F�$�5s3Sa���_Bj��w�� ��y�Ńz��vh�K�~�}�^�!�.��+Wk5wM�Oğ����S`'�ǻs������z����S�A�N-�a�{�f�S��o&i}��Ku�ҥ���!�V�I+un�Z��nY���L��"�����S~�I$��{�QI ���p�xUx��7yx,�8��>���ԽWSN�I!���H$�K���sBH�~���}��y�cmsl���&�P��d+Gt$36f�%ޓ��%�:��#��O�Mh׽9�A$�o����p/Ofmso�ױ�����@�VY6�h���bs��om�nۡ�&�UAV�Lr: �^�k���*�Z�Rr�S~�f���k ��I �6?L򣦓�h ����lF��X6.��3�z9����2F�V=��}��I }_$����[�ި����/L��^�c}VK]r�������0@ �;��=�?
[��'�V9��I%��w�ۺ�/�v�$��!�%".������ޛ�.��p�Mω?M��$�Mn�I% �oj����<�~�|���M� �ҍd���QKS�Ε���{�A%��ϓ�t��1��:;ns]Sm�7"1gl�(+d�޽̕lc9_�Q���_������='�� [$�\���s{؀H��<Ѫ kjU�z���{sR'����$�A�{�J&�\���ZU�������qG<�.a��\0�+Y৞���^}'nZ�I\r{9��2�-$EV>�����H{��B Ov����#�$��F��=D�9����Kۂ�uV���YWo�΍�~'Uɭ^Tj�ӛf� ��t�I&��Z���"�ai]yۈo����c�����u��B�j{�l�~�f/3�r7m��I=��$�� -����ݚG[�r�W.�wь�x�<�/�����rA%�H���H�o�>rc=x�C�;�Ѥ���{��Z�kl�X�v��|-g���l&�g:��/T���0�Mc�� ��z< [��_*/c@ד��0`�.ԺV5
ƙ�Ɯ��T�4#��.��n�Et�e󺻆Gw.��#
tqݎŤHq^�xxl���)���n���%���%����D���^d�;��Ί{�D�Dnm��f6#-h������b��u�ώ*ZMc��(���Hv�fGrz��\HJ��+�ٸ���MLǚ�CH��1�ի���a�K]U�%ݵvp����$��,��)Wm��-Vc�7&`�&�#���n޻�2
E���lPg-�͔���2A��j��:k��,Ty0�nI�j��n��}m��[I�y$�e���2�������7c&m ݓ��`���mͲiP�x9<2�U�Ă�r��홛N�� �)��:]�i̖j���7P*꼘�X�+���2+Fi#�5Eʑ��X;(��n�u�[ۺ��8�r�2�[W��7C�V�k�*�׼#u}M��ޜ�|�T2�~�f�pU����=���"�,�.�F}�oٝ�N|n����ȯX��[�EU/��u��uЋ�{G��T�Q󾽍�'4�Y���t@	�M�Jٲ��#�r���Pj��Z�T�9�үF�H-6Pio�hƁ퉹�-]8�N"ƽL��eɕ�Q�,L͔L��>Ý�S"�B�h<��;���Z�:����C��Z���>�ΰs^��z6�=˖������S��j�/��ŗb�7*Q�3�8�X���l�V+K���֌���>��P�:�^f���`����bm��o��ѣ:�c����\�}�6�6��cm=B&�ue��'6ɖ�kjУn�i�nkgX���Xd�`p�l�af�V3S�e����miD�l٭�l��,��9�:Ps�p̄B���v�
3skQ�pա�h������"DS��2,��m�A93r3M�w	�'��:D�	9���LЖZ
�"DM�Ӆڳm^�I�i�˂����:�Gm�m� �;k�Y9n�4Kk,���������Lƛ����we��gy�����qN�d	[Z-3�v֑9�8�m,�5��{��)Yݶ��譵�����N�f�kdC��'I�7���"fe3�E���`m���0������E�zTд0b����7� ���v,s���g0\�+=j۶�����؃�Իs�m��8�o)lv�pu��8UCZ�9��N�(����m0�05�hw����'\Ns��ۈꇶź�r���q�#ۍ#�����k�����c����S�j��J��Ч:��n�y�Ae��ۢ�ky'W@A׬\q�Z���j;�^ݰ�'j��v����v08/hx����y�(&i˗)�g���9�ۚ)^2��*�m��k�]�'31�s����M�Ft��P�#�`�u��g9N����P�{��f=���춪<�s��wS��[��k�۷c�/��Wĩ�H�".�vu�o[]��nֵv�O�iN��]l�s��l[�Ҏ��:����l� 3�۵]���7;��^:y����ټZ�����.�X�^��Y�(ɼ�����נ��m��p�n������Fن뇦�x䆧�5��zݙ�*3���/;;�R�����n[:��j��ri�^�����'�-W���{]�6�8�玻�4��+���v:@�t�a�M��W<:vKKgHl��d�GaLY��.��W|}��u��<��
T�l<G{l��ĝ���P��gs�Џ`�q��W���m�cxh�1���Ϝ��<�ӽ�w>V�:�n��v|�x�c
��u�%h^�&���7�nU��WG/R;�b���ewY�'�K�ʝQ�gyMR�ub��ΧO<Q�|���-�4.�ϧ��.,�qx6<��iz�E�lSv�GOklRNخ2h[a�]���f,MwW<�g,�&���n��[�t6:V��E���=me�=��
��ƣ`� :ۊ�k�;k�1���dy{jzCX��n�g��v;0�}u��d�vqGb�2��DZ��#��۝���<��9����\DWK�D۷79LT�ݺ�v9�����t���(��{s����}u]5��3+s������ϛ�R��ɬח��׳q�nÝ��q=<YH3�g�')���^����^:zY؍��n[^���=oO;�ٮ,�kc���)���5&�j����뎻l�F;X�׃�e�u�A0>�� qo0z7��o`��G��6�v���<��r�:�^�]��ײ��U@� �4�=�\m����r���[s=����F6�̧:}��&��I�	�����Qdx��^���}���D����șK����?����/?��/y��a�7���@�����:�A
�Ӝ��������Y��o�ZC*r�DUc� Z�wZ���-V9�$������;�� �����q���5��eQ&�!�p����T�_�k� mw��Y�@ۻٙute�o��%��wF"�H?ln�<���e�9�e�3~����
�X	֠�Iν�:��$�M�H�<���3�M q滙��.jb�T��Mڡj�o�	��7�^of���W��tc��~���$�k�\���yN� 楔oѹ�u��ro����j ��N�n�/��v��n�������Ӹ�q�s\۶����o�����r�/7��ȟ���m�M~�)�BxkTx�[_QC}��Zg��5�Ł���>�ڠ:;����p�Fo<wP��W�U3��hFQ?� ��n�u��{��(�G՝]j�������SA+d=��e�s��������}4ZCfʅ����c���R'�I&�w/4�$�I��)�'Ě%j�함k7ϰ>�9�v7+�r�`+�ܦ�Ēg��$��t� OL�O{|Ԫ$j��2 ?w�������.��%�,ˈ\�fq=��}��<� W�c��?Q$�r|ܪ$jr�N�n^�s㼯h��k��,7��uZJ�N�y�'�n�1	4MM^HaAx�:�pOͧD�$�9>�h�S��;ӥ�s�{+���d�J�(�[U���e�g�كv�H�0
�\=���s������]R�g�Mw{[`�O��I$N^i���(�{$�S�6� �<�I(��co�FJ�)^�3~����p����ǚMS� �&�|�I(��$���� G��;�t-�g\��>@݃WTN}x���{	$
�\�����D��E����̡�{Ӗ�\7�w[���ȏc�����2�n]����Q/tW��1u���e��*�z��cq�t+w+��������z��"��sՊI&e}��m��_��s�ZR�)]$*��ֳ�f�uc��.�A&ۛ�rA"Q�g4�$j{��"��r�$ �I {57���Y����f�x��y��ϝ:��y�����ʏ�X	$�Byst�$�����W�~��x��+���:3ۏ9�<v�sֱ�D�]m�L[�L�v�炂��P���>�IaQS�������I$���$�K��怕�ta[=sޒ�y�O�4jj����r���˺Ì���zs��Ļ�4��oG�BI4I�M^i�I��N��~@�^T��Ͼ幜�z��:���VՅy�Y��4� �o��,��)��k.���&�d�������:AH�u/A�A�ݢ��\��}��漎^� .��}����3M�A�o~��y��[�O&��.���Gj�+�'\i�`o�ݶ�at��6{5���Pݱ�f�b킬ps�!������t���V?z{�����}�i1�v�Կy��lf�R���k?8�l�I���O9P������_��>&��I�~$�k��n��I�9����E���QQK�!"����uS�9x��zv���vjxu�.λU�̙⧶������nQ���w��{� {��}�"@=羒Q/]�Fu�&��̃� ��s3�����!JXܪ�"�����'h �!1q���i�L�$
���Ԑ	)�~���#�}~�uFķx��滚u��Um�R�}�b��k�lB@�#n	�zuГ.{S$�h����� ﳞ���|z�M�IU�^�B���U0�c��$HowF�I���I	4H���&CʳJ�"���O�i��<���uZ�R_����s�x�6t��i�]7	4&��$�'|���I�M�^m����D�R�Mj���g��~N׻�U�	�^9�7ݔ=;�b�E߱U�&�b���t�|�%mlY��bX��8�4�!b�9�����5o�[;c�8����K 'f�@r*;'ҿ懣ZL\eU� )�^48Νt�5�Eg����\�i�N@�t�s����y��%�V):Ń�gn�spv��<�c���ls;oo�䰗.8�;�<x���m�;�[�v�881ě��K�Ƒƹ��E�]����Q\�k^��� m�ʈ�y��v��v;n7\�2�ϛ
U$�^f�4l�x*���/Z���o���gn7n�BƔه�s�v�l������QZ�B�=�>��o۩$�orA$E��愆�XB_��&��4$�=�%j��X�*��h�J�oBf�D��J�6@�o1����{3` 7�f`���vh|��ƭD�f��sy4�k�UQJ�k}�wr�?Q&����� �)l�a}�<�/���Q$���t��Ζe�,]�P�z���C��e���b�}�����#`I7�:$�$��FJT�I�߹돈��}���������GUqЙ���$
��齻^�;K���ߤh��y�*{�uL���~b����x���������6�`z	���g�+������r*ؘڣmX����Q�:�U�k���w'�H@4M\�H �4'�4�&�ۣ��:/�{=$$�h����l���JꐅTz�Y��3��߸���%�R����x���y��F�5��ʗ���L�IG�ҙϲ����WaE�uH#0:&h��=A�5m/���)��M�|�ŎW{u�Ȕ���p��$󝻨��-���\��H=ˢ+�*�AfV��u��/{�ϳ z���n'y��I5~�m�~$���h:�9�9U
��UsX_s��_as���z�l$$���J� ���	�{{��&
*=\���j�&��m�Ӷ�e��fe�a�]Q5�Nm����>�9�Z��[���M�m ����m�j�5<���/�z���� 	�e��F�rT���-�;{[��r{f�N0j�)qJ7Z/1�=�(ӲU���sy�` |�kX ~��!,E`d�Z�K���d$ѭ�m����G��w��.a��{� ޷-K��|���~���d�$���.x�g��p�D����Q6~ːV��uIYT��Q�q�]�h����������0�/�N��N&��f�FJ<�h.��j}9�hP�Ÿ���w$���gm�r󕚿�}�l����{uݙ��9ə�S;a�� ē�f}���k~���Y�:�W�S,�՜�{^v�9�b`�ݢI6�T�$�=�7x$�	/������SWJyxC�*�c�6���$��'2���cN�n��4M{7���OgrWuʉ,���H<���H�c��jg7�yk�9�^�"���D�4ڟK
4�SWN�\=m��x�����[	�k�Ev��K��zʂ9U����q��y�{Ò	 ��f�2� TswCOn�D$Bw(m�V��%Q�Mg����ϰ��;P.�� ��a$U'�`:�I�ݍ���g{����b�-�]3òU�n��$�!$�����  �r]�j�<����$��;��I$C��ߵy��*-ERUG��+�u���\2h�����>��A$~���$�x��W��=�S۳L�����	?�N��h�G�5�̳���g��v�ؾoI���;.��*��ٛ'X²b��ȍ�U��;�͠;�f��
��L��#�7��Kǽ�Pw�Q<�����$�D�~5�to�A�O��o6���^ky�k~y�/5���ݬE,�Hڮ�'l�r�ݷ&�;X<f��G
��d����I9��uUd����"��������5���x�玉7����������i��7��R��f,9{�-��v�eш=��ǀV�g��)l��ztluI#��Ӫ �s�ĨĂM�k�$�ۇL��s���)�o_���
�}�Kσ{9�� 홆��U1{�����o���w��3�~���(%�*��)j���½нz�vgz���=3�H�V�a�$�z^�D�k}�I��嚃/�?�k�����J�QT����>��ŔD�g��*���E�x8�xM?F��MN��6H ����:���g�u˵u��H�m�Zɂ�$Բo�ݙ-Ey���Ϊ�P����ׯ�����X��ZO>{y��L\�RVn�Z\�����v�I���k�1%ι-���PƓ�m��tCa2�#�[:��ѕ���d�j��V��;qkR��"�{pN��m�ձ�<��gs���q�3ú�&�t]�����l��WKG�0H�"�S������+�0U��=����=��n�W����2r��+���Eük�A���M��9'� �5bl���Mat�獧���3���Pxu�;m>��h�U�ЎC��^wݞC�m2�_�[��D�'ӽ��I&�;�rHN���E~�ف
�{tE��t�����k>��GQiK�ċ����&�l�{4�>~M� 5���d�N���Q$�Qn��{dyg>|��`v��j��;Z��I޽�JK�ooH$�K����1��$J^�/u"�A�owrI�k�5$�G)���o����]��̢�f��I)wb�4I���B@?�v�Os�����H�T��e�[-E�����$�H9n��������3�E�4I�6��4I���$$F�����z\{Z�Ĩ��겱Z�I�h6C�5�5ַ<0Ѵ�N}>*!e��*{��T��HJ�)O ���é 瓷�"PHzN� ��<<��W���ǹ�l�I?o����Y���ZPY��)��i��8��GY�D{ԛ�ӭ��n-{�)l��Dc����4e�f�yp~C�$=sY,�-�#2ve*��N5muվf�\�F5W�/�I <�ww$�K�=6k��I�1 ��w�<WHZ���eÇg:wI� &�ϓd {HÇOP؉ȥ探I;�Ѱ'Ċ��N�5m��tM�E�`�e��~���ε��)���	u�f� ���w5� =�K՘��we���� �ۡ,��������(�� �v:�v'��x�;$�9$�I�I�/s@ =�غ��;Ϝ˻�_)N�o�{�qF��42@y�2��'7k�Vy&W[�E#R����A�bp��B^mmx�VK-E�9{�o{@��wX���I�=��'ڪ�*�n���{��p��{]�}���n��D�����j��jA'��o`��%�^����JF�˒�h��cd�;ӓ���2��,����ovĔܾ���l��������uϰ �=������{4����4�]���@���x�ZlEl1¶&T4o�4�v;�r��&>9�e�od�Jk_Ǵ���w����gV�k2�Wv\���s!T�xs
X�ƛ�i�*�w�m�ԥ�☔6�Ht�O�r���£+bξJ�̇5���57R�f�����tM���Xڵ���Uv�J9d�������nu�]HLK�ݵ7Vn`U}IVd�ڍ�U�e�Y���7w��u�4�E�p�&r��c�p:cXp�k�WW->�M�QW{��y� �7y}60���ϫ���\ҭ:C���Z��&�Yz��Kgf�G�s7*�sY�*6�N0��*r�e�*�t���N(�e}�6�a���,���f��"	�&�����Q�H�a\Λ���K�wE�13��t���e��rXg&��We���sH�QΙV�ɺ�:4��ft��uv���v
}�r�@�dA۷�R�����w�R>w����Nr������kUS��<cwD�C��2�2�b
o���3�襤��n�``��vG1�����糊�I��:�㜁*V��pt�=��<Yc0T�f>#����sHB	!�z+���Ȳ��ȾO=��������%�jd��Z��\%o<[���vX�כB��S������R�^���i��r�N<�+t����r�+�O�]u��r�qb���l��j��,ݪ�;ˈ`��Ί��/J1�T뛢l���a3؄�.V`m銻�/7)ѹ�p�͠�K0^P�;-��{��_������s-9�c�.�,�[k#���9v6��B��s���V�e6��t9��ܗ��Cn��iYnu��kf J*::�Y����=n]�J�nW�`w�1��gig5��n�,F�g':#Mmc�֎m��qPr�3[[��IIIn�'Du�iNFZm�4��'�G:mXI�brC�m��mgN��9����{vY�ڬ�A�okNyc-6�ݤq�"t�ge�:�S��fvu�g�e����=���'-�%�J�BGm��y�rr����!%r���'�G�P��̳Kl�E�r�ZH�q�q��8�����9:�rCi���mI�
NRJ Nm�:�l�FC�� ���`;�*�� �{�����s�1��ޒ����WWW��_��L.�[��/\=�t���u� �{X��>�{]���{�YqP���i篹4Z ����@�y�U2'ں9�#=y�QY�Y��'�L��_v6H4I�.�J$n���;�
�H�;-PEl`�#c��^:�����,��k[v����@�Ԟ�ￛ����2�"��<�2h�L{��4I$��I%$`���ڙ����uL���w�1c���o2�7F�&�� YzTjԭ���HBI'�?y0�I�.�B@ux3g���5=��>��~��*%P$���]�J$�O�>r o݃c�y0lھ�[@�=��� ������N*
��
��U���w:l{�y�� 3y�l�$�>���$F��]/_�PW�|��|ſT^,�=�ץ?<���M��:핵 ��%��]�	1�\&P�̀��i6{����w_�N�t�^���#���g�/of��-���sOד�B&��Sgr�X�����M$�a�I�MMS�|H�r��f������o��~��n9al��^<���.�fݎ͌v�@ۋ:a�pFn��}����vSl������:dD�)�}	���5��I�⎯n��d�3_!(̓$$��z@&�2�_������{TZɢw�w��ܕU�~���H�����A$����4Mw��)&��$$��xE�ˣ`���uz�>��H;�0��z���^bӰ}~�	D��;�z@ �����'��]b��p$��0.wuy^���.g�����ٽ�� �{��$s�G�u֒��*jz��>I
}w��]�
�b��dh� �=�n���Cw^I 	/������C�&� �&���7�7��p-�<͛V�2���(noi+ˤ�u�sw2�9aM�1�Ȗ-W5��'E�]A��
�6c=�i�ʘ�To(}b���2���uY���v��wQ{r[n����7t��&�##�7W;G��1p�٣C+��Wj֩�2�Ύ�O@za˷q�t�q�!�םS���p��{L(�x�d���7�W:^퍰�^0׵si�Kv�<��6���`a��ݝ��=pF�K=@�������/!�.-&�hWlӈ�l�X[��k�#���h{y���X��Y��d.;t>(�(�3��?��h�NKe������� ^��� ���F_��������uS�� �ks����gNj��'%�\0=�ő�w7vO�8��J�5�A$@��sBD���q�3<�VL�J��9��$�ñz9�d���f|/s9�� �voF .���,�����v��� {������f�R�*	Gs�o���Z�&j#�@�=��D���u�Z 7��3#�Ǵ ���b��.�Z�J8Rǘ��f�썷�gy��g.|�����l��{�sBK�	�]�)��}�BV�T��Ê#�f��4lj�<svn]��� ؝�1�vb������祋�g7��X)Ti��d��Mwى` >��;?h�������W���;����@#���yrT��R0�._+��H��s=!r�JTꅃP�N��5�i�F�؄�h���0U�m�Ʌ�h�f�b�l��0pA���=����c�8��K=��������z���gy���yTn�x�i?ige�W��5Jԍ��.�w�<�$k��P�=�:�Gq�G"R� {���@�7��7��>�ΐ�6[D9�/s9�}�oQ��o�t�>�M�Q'�I�>����dCt�,:$�k[��{���!K�%����}��H{&h�े�x�������:$�ޛ$�$kϹ�����M�wn����,���n�f
�U�N�Yw�\����7]���^
�V�l���~V�R�����\��MI��\��I�H��i�Ml^���.Y�;� Q'���	�.VY��b���hB�Mѩ%�@���Z�gf����'�L�rITH����A&��*Ű��b����Ę�U��j�ݜo�=�шH�ܛ$����~�ٖx 2��^r�-��}�����V�7Y����%��Q�`����s8�k+}0%�����b���~o�l�i�]WR�u��o	�.{V[X��� �y� ��5'�5hUD���jߒ��Xx9��Nn|A���7�� �N���`�H�r�?eSTѿ6}�K�����a���YD܆g�޽�� oy��X5 ���վ�q-|Y�;��	 ���2ē罍�Mj���-gq�mX9��LF��=��c������ob��0lY�)�lX�`��-��!B�PJ;�|s[߷��Mgw&��My�&>�>��JB}ϙ��i�	
���X��լ��A�K`]gn`�-�ME�{=��[P��4� y�bd�L������
����|]ɛV�qUI0jz�\X0h�?{  �97n�J����~�5}��0`�s�3��or�eu� +U�k��eh~�
�k�9�H�{���&�����&��S��A�*P�|$������لt�9�E�'ar߸�$���9����֠�̷#��Dؓ77/���K�>��ת��w^��+u�)r�-ӹ�w��j��h�ݍ�'�LӴPN��a�{������5���6�8W�u�]��5�bd�I���6������f��]Vm��6���R�Y�T�m���m���/����J+dnV�|�P_{��D�,�p��B��ŀ�9ۋ  �g����˿S��B���=���I�~�σ�S���BQ�a�o|����ݻ�N.���η6&ɢ@>}ɇD�g�����TIo�y�Z���*F����5wk�I��=b�ۦ���qʄ�~&iZB�o\G��h��\HΝ�������h왵a(�NWB5;{��f��b�����;�0�o��$�$�Mg�������i*�ݣh�]e����%mu� +&L/9��� �	���V�yw��,�K��4�I|����O/�n�K���H^ݔ�\��۱��y{�:����u�^�`���z���|����Q�̒�Cq�h��J��6��9o-t���W�I�߹���'�sK4��4�S�
|9�������;F�������뛸���@';�5g���=O8{5�^s�9�"�Y��zǑ�&�ض9C]Mۀ�Ne@(��n|�Qn�3�=^�8�^܌
Xw\u�볺��������nG�n����`�X����[�Bv9tm��{q�;�Wm���d&�j�Pr���(�2oQ�\���^PC���l�@�2�Nޛ;p�;
a��h��*��#Ƴ��T!��}Ee(,�!.�ӽj�	�-jN�=t� �3���l��֝Q/ưיZ�0酮x���y�����ޒD�d�:W���g3��zWG��]�C-vs MN~�! 
�I���H�����Z�#β��$:Ye��F^U�X�򓤄�~&�w��$��ǛC��]�Y�8BI3ϵ�D�
�����{�����$��Kb���p1�Ƽ�;��s��` >s�njH$��zN�J=���|���;{���IGr���υo;���/{�x^F���˼	�	/>��� �T~�'R@/9�����ɠ���o�}5�î)�o/H:��ge6^�s�䣓��
.�:4m�A�����K)$�lﾬ�Wdc�ds|��P�$�5~�H2M~��L2SW~u�����<}��$�I
���Ԁq��[ �Y,Ra�����>|�w�y��z��*�Q�����l<���b׵�&�����	�sv}n�Ŀq𝾢�p��kR5�u�j��Ha�E��m���M~�I }���4}���E%Ո*�Xv`��y��$�T���'��߹�Ńb�s�o��n{�O��K�I$���hI>�r���[��eT�����o�����zԷޏ�MQȐd��5��L2M~�s�w�n����9��5ڵ��>���Q�#v;c�x	 �~��Ϫ>��K�阺牾��A{ͦI(�Gy�@w���M^n��5��kA����r�ݴ����i�GA��G�m/F�׷j��m�l���z����R���x[ֽ��	?�{��L�@?O9� uT���d������Z���{�\ϐY~rG�qb��t��R	z���T|�ל����~$��&~$�O9�'Ě�S�^��j#ތJ��3a7tEU�]إ��y{9�D��s�B��������KnS�yHP/GSB��閮О�����/�5U��Ҩ��7ю�&��+��4-�&g7=��՟z�y�O1v^���� =����07�߳6���ޗw@�ˣ�f�{Z���>QzA���H��{�$L{�t�H�~���rv��*
�3��1�V�w����ec���&��D�grt˞�b�-J&�n ��<�Mn{�d�=�ߟ�}?���g�m2�h.��t
���R��ke��$��S��8�������߭�u����ħ�S$�D�s���'�$�/}��7jWU	�g/�+��N�	!�5��?���G�$.滙�Mo��>3&�@?f��%h�ks��̃D������V�ibWy�D�AB���v�WKkU��i�� ��0��R�j��!�Ѥ�$�O)� 5��n�<�ͭ7lh��j��}�SW�{H[�i��ozor%|�_�愉K|�>������;�/!9��P	��fM�<�E-D�e�8;�̞֡������n�J��4�n�հRT���z�i7b%��I����]�dL,�"��w�f�$ f�ۘ{��kG���{3`�/���{�����k�O$�vG�c����l���v���\:��\u�\np��˞r+~�~g�Z�j�ڳbߔΏ���$B\������d���K���m^���� /^�4�{��;U	��b�۔ɢh��c{n�=Լ؄�M�sO�@%�v7D�Jc%���(n�u�f�>y���5T�R=.滚x��3��ϵ�y�x�|�s���	/��&�@$f�ۘ���]��ŭ��&+�~��XR��:�H�Z�7�����y0�4I�)�"g|C�b$W��N�7�1i;F�U��0��}��`؃�S��E=��^��/�d���M��tH����� =�= ���R���rċ���^m��&��Up�.�+-�vn�B��6�ʹ��Z�
^s�*�\�yN�>2�,�ۣ}��F�*��G[�e[����+Y]b�.{w;�5��<�Ɓ��bO���`T�V1H��M2�_G��q"1�0�'��Ǧ�b�����T�#z�ˡQ
�x�7�[a��۟I�m}Y��d�baHB�@�y�V5�c6�����j�����{n�ΫS�q���r�E�����r���/whά�x^���|�e�.�e2�#i�Ϡ�.��������QiS���)��c]<�S��ѳ;���r��ԗ����3	�Q�ېo��ۧ)ˉa��(��RN	�t2&uo���=�ŀ�ֽ���O�wgA�[�T]os={�ub��lu�ӑЃ%x�3w �K4VXݠ�Lf����'���H=꼙��{��2p˖:v�*]�0�Wfw��J��di�����*�i[�'6��i�7[���<Z�K����9	ws3K{2���r���B�vFWsm��
ޡ��oWU��v�	.֚��2��Y{8;��� �+�x��m��Q�� /����S�{sL�
j���e��m������62U\�f�X�&�hG�����\�}��-{��;�gRB�ETۥ�� �j��a��u�u𬥝Yʖ�嫐�H^�F#}{{�N�X�V-�[7_����o&q%����Y�3'^cX���Xނ�������.���;q�W)%ʗ�_f�ū�հ֫q���ׁ��e���)9����F��9PX-gd�
(�yÔ���A#1#;"�m6��6��̵e$�4�J���G�"L���twE!p�8��`��v�;,���8I6�kv�t�i�\̶��r�kaja���q��."{vpwy�vefq���n����f�^[��W���.$#��՝�c����݅'BQ9�:γf�荷'ֶ���tڎ2��8v[c��'��m���-��4�-�V֞�y�yq%�E��j�9mZgm�Nv�n#�f�8�Y��f��vu��m�f�����I;δ�m�q�Gvub۲�Y�n�F�@Dr�D�&^^q�\RU��&u		6�����"N$ t����7���>�綨�t/n*�{��sj��wY��Uϛ�;6�v8ݷ��Y��º�H�>�G[z�;\�ڇn�&^��l�ڴ����> ��gkʮθ�xΐ��C���0��3n��������V7Ez��a�Pv��]��X�k�{��$�qe�tk�4� 7`����:7���]�H6@W�cx��c���y��x�������[pb��Cӂ�ף���uݺi�7W]�y8�9��˭�{�,/8G���/Y�򃓜��ĉs�6c��q����u@sq�ХѷT����9�Ϟٮ՗��;n��k+\..���8��m
vލtt��ze{���3����n[]�7E��v�#�̈́�&�_�y��Zr�n���,���̬��ۓQƞ-��vxg�s�\4M�6�����OG�I֑����ݵ�0v��H� �Cϱ���Yg��5�'h��������ol]8��x���ɋEڽ���y����9��;e������b�q�W$õ��d3��et�x9���K�ͩ{e�"�ݙ�@nr竘�`�sU���;m�k�\v�m�;;��<���7�n�ƭ�[�{/M��/l��`�k&ll��۞vk��(ú�!�[ō�]���c	qp���q�-���Z,;'"<wm�nۣg���a:���#�vf�!�ˉxg1j3���ٜ�.6ۈj��	��$=�;�>���8w.�Yd#������B=�7��TɑxL\s*�"����4�G����8y�<��v{>�z�n�ɧv@��^,�n���:��7'/�h�D�ajV�L���۩�0��pp`��Z��tn�nz��Æ��+��)Ɏ��x��]��nm�����Dh�Q�>Bۗ�,gF��6x�c�{\;�{��]a�mt<��v7^nހ:��.."�S�ݺ��5�7[Sp5�:B����1��&��݇l[; ���qn��5�6���I�\[Z�q=-�Y�ڃ���g[F���5�c��
7)�ή�q���3��q� m����y:0g]j�=��F����%���)8���]G({g�'A�ݍ�I��Q������ێ�[<4�\ά�{q�ZY�y݅K3θ;;��<F3�NJ.3���,��+�cEW�gr�.a�vշ>n2���B{>@Ъ�����{9�Ջ#�3p+�]4;��q�qI�s���Şݯ\��=:B7� On %�P����g:Y,���zjk�ז�D���|I�$�yOI	������N��Q�d �buD�v 9��w��Õ��)�$'�r�w~����֥I$�9�L2OĚ�)�% �����y�32=�Ξ�I����ZUDݛ��|3�>�@ ߵ�f=��|�w-�xž�g!��&�}؀ w���������vU�V�{��{��DOGf���n6I'�g���~$Ѯ�7�B����]x���v�w]م[nN
Xdϋ�s�Ǵ��{5�}��u�{փ�I���&��O��D�~5�绨�@���&�4yO^u*<6HU{���.��Nx[�p��^�`��T�n
PF���j��w�S�jʩ+�;���@��|�$�Ml�I�+w��׺-��ġ�;�ܓF5u@�UZ��Y�+<�D��dz*8���ͦ\Y�fhjѝ�c(�|z�F��}aP�M�4)�^��l���y{�PfZ�r��/��U�b��S8s�&�b��ǀ����Y�}�r#Lչ�OĚ�M{����$���̂M��=�-#����n/j{e��+v�\�_o���	 �{}�b�����M��l����+�9�I=��ff��ȱH�Hܪ��f��G��ܿtf�OĒs'G!5�$��=���&�4u����G�>��@sm��)j�ʣV'JG�|q�[�K@�A���3H��o�{!%���Q'�MQc���"I{Ꙣ�=�q�A�u]=�OY<
���=��yT�����엔Y,a�ոu�Q�y��ES�����ܭB����߻��1�٪��>s={�u�ia蘮,�} �?7��uS�t�Pc+/.�Q1����lO:g�_��<�zo����ω'�sF�v�׽AH����o��l9wC.�2������
�{����|;���I���^c��IA��mV��u�^u]vs�	G\2��N�m�pd�P����9�UnTq�uT�G�1��A �����g�5��B�?��e^���zG��1���w, �y0({W9�������X��ڒ�U�a��/+2�5�b�>o&o�}���V<�^��Bb�u��<� �������=|;֚��>�wtp�e�uϜ�]�� �79$۷]Eۚ7&h��r�9Y봒{9�(�:ⰲ>�??]�V����6> {ڹWr6�����z/��MOs`W8r� ]e���U�s��(y�j�9����� �y����͊q��a�7ؾξ*����3�]���s��$��ɚ	#�G~��[���BI׽�bm��s]�o�Q�ab,�XJW��}ޱs�p?:���h�]�f��={tI���)r]~$$���`f�<(<4�Ne��W;�@���i���𫨩b��qfؒ�D~VO��c$S;ʶ%����a���1���څ?�-R�m�3��ox�5��jC��H����ص�@{W'@A�X�[�����εq��N��À-�i5����Ϗo�&���bN����I 
����u~�_�T�Un��f>ߴ|�L�	��H������[/rIxw��P�{u�1�H��yW����]�ƎȰkK�zL�S��䩀L�}�A�e�O]PW�.��c�~��� ʼ�W��?�O%�
�vډ7� �������� ��*�N��uB�[�����w0���\�;u���A�j��'��� {�m����_���Q�����]��Y�C=-��V`����������9o�P�۩��>�xH�9�DڛQ=z���c�T�j�M�j�8��|�|zcK�>�T�N��������������ݮ��U#����>��+dy�s�u�����;��Q�������.a3�@��]<��[�RP��b��7nn�k�v���!g�!�1�z]�΄y6�x��Q��/���0��)�=��+s�k���hz�ðt�ma��/#��Ap��R��!.�£�5����{	r"Bnԏ�-²vPp{v^zS�w�Ӟ���͌��:��knx��g&�Y��<�θ���Q�RhmA4ө�����4��9�0�%ͪ�@PC�Z�	�lm��/�,pU{;F�~#$��<�u���R�b��������b#6o�C]��g|H$�e�$���h%�����5��i�~� ��LY�J���T7A_f�g�4 ����7�`Gכ�4���>Qv���8n���*�Y�[ȯ.|t�x���%�ϰ�I��Ѥ�y���,�=ޛ�y��d��/�Z�+���1��|��o*��Ƀ�Po�L���n�r�ر�0�J\h��uMj�us�&����0�t�3�G���ѻ]��]���ˋ�]�[T�Z���jk��Oy�y�� }�l��W)Ƒ�Ç{Ue
/gy�ğ�[}�֖�l%��\I����f;���]�dh��ge�ؤL�՜��33VX��J�;(T*C���l�:}���s�d�Vc8�kؤz�Ք>_����l�� G�����g~��ũ,#�*��g5����7�4Auv���u����f�I��}7A#�1iX6��7Ct}�3�:�]u�M�ӷH"6��&�{ʚɶ|�w��`��rP�0+XMѵK>�k��?q�f��z���E�+󛤀H����$�3��?o���^���};�1R	�b�a�Cd�8��-vc1�5�w6�5�����aF����~��`�l��"�����ۼ�`W�hp,ӥ@q;W+}3�}���Wt*��ҫ6s��h?Oe�oE�e==�d�(P���t>���ټٞY���p��$��Z���f�}���+��U�{jZZWsɛ�2��Ru�p����h����ln�㗫�A�I�y�����,*�\�э1��&Xq�*�ē<��$D�facz��7TJ�b�f��)��iֿ.���t~X�$���Ҧ0�e�/b��y��X6��*����3�'{�:3�t�NǮ����t��-唾G�:��o��o}���q��B�h�r�6cnq�G=r�/"I#\5,��vf��~~o����2�0��� �R���#�7C=���лr�0)劝��,]gטM�%�nO���O����n�R�;�`���5j��#���j�:�����
�!���a7���t�_	�|��m���r�X�g� ���,�@T�����o׀��\�������C={�����O�������L����¯�,�5w#�
-��n=�I���g������~�[M���[�9�ǖ�&�9���V;!��%7hv���Շ�3�j^��u4`!o��}�W�Y��p�)D�����4�~m�߉4g�f,�瀈�m`����� �y��i}P{����z����Ω	��'e<�Y�v�cF{g[E������k��n��V˾y���N�;�s����m��O{t}��t�uo��2c/�,���Or`}��s� �a��oy��-6���\]^^�~�� ����^��n��c���w����J�߈��ǝvF}y��l{_��>���L��{����yvo��$�I�#�}7A"#�F�Ѫ�n��z�F9��{�Vry�L|�Ol�Lޖ�;i��m'��Kٍ�q>��VUK]�����^�J�O�����!���f�H$���}}�0��隓��WMث�/OF���J��,�2�]xd�'�)צW��2��N��)��+�\��O��D@ܺ#��Gt}�.T,Rb���%s��eI;��G\]ٮ�W*�޳�q�3�x63��=�세2n�;�]k��W����o1�R0(ty�!���ʇQuc��:�9�=�Y�ݻɛ���lZ��]�=lx�:�`��v��[�gqڹ�OK����$M�Q��-9��ݵg]4{b�ke���n%{]�<Lrg���ne�Ob�&x�'i���3rn����Վ��Knh�U�m��iu�S�\��6�\����o���+�B«^-��?Ko�i$�LAP}���	>��<��u��F��������������RՋ�f���L9��Ck�ݸ7�|�{F�D�Vg�'v����&�l�wm��eX�aR���j������=-"( ������y뵛��A?w��� �{�1��d�P��r�= c;�?�׭0*�zb�
���� e�ee���+�-��%N�ƻ,�ƛO|�{{zƶ��_�k!"]����As�1Ov�n�>���h�5�n�����d�GԨ"ӵہ�X���]uې�v��%;F�������۝�L~��n�$^���$�l��/�#n��l��=-"=�]".���a���~L<�^�.�'G��ۿ�E
FG�� �]0�f������`�(�R�mt6�;�v�^bIl޺�v�Ŋ�R��v^빞'�I���3�GoOn�H7X,�ߘws�S}��S�JҠs)1��j��>��1@=�l�7h^{��� �z[G��s��P�� r���*��dיq���~�.�f ~���n�O���>�$�ta��|�E%wG>��Ã��=�'��:zJ�˖\�,��P�=�����{{�Ý˞&���$+��0���֭��[sF7n�ˆ�uţzA��&�-MPN��x�:�rV첏�c�b��9�ďyɻ�˞]V�!T�b��M�OަO����5In׽�F�Iw>����I��٠��97@$���Y��r>��`�l*j�t.^L��4?$»�S]-��J�9\���t��k�ftt�s%@�������c8�	������qC�IK�o��׃!�ʭ�r���6����X�C�<�nX\�J�Mf�{`��u��U�6�4p�x޺v��8�v�ƶs������7'Em�¹�r���J��I�qhCx@��¯�`�3r�/wz]YE�!Qi��k��e=�wwu\uYcz�ZҒ���m�!���*hqY������˻I햬��-�O���N�u�iV>#����Ա�Vsr��N�Q;WV[6�N\5�P�雬�&�,w`������~Y�y"5Яv��=�؆u����Kin%�Eݙ)��p���u�FSX�ve���
��fE�.�|��,m*��]J�h%+H|ٙ���n��-���i��<���lGI\7�f�(����\%+�K)�N�m.(^W��Wv���32�ˢ�٠��P�V�)���ũ҃�cq��)�i�ڕ�ك��j�����j��uW�ժfּ�:��: |�p�`�f�%�v`����qi�r�]'rE����������is�̡Zw8�a&༥�uw[[�&*<nY�[�Vu�Wd�w*]����P��ù3m�\W.���,tBvVe�d&Td�n�]�W,W,ɵ��5��N�t&vms�hV��<v�����7�{�0[���']�M�ޡ�ve��0T�[���+���p),�,օp*)��L2u�ӗ��l*B��;.bMH�(�,��"j����[�Қ�=�r^�9s�o�9��?yMZqq~K�N��2�$���,��(�::ɚm�Y�^��)�yY՗dwHNt��m���,�:g��;��˭mgqDt��(�@)lۂ���;$���:smsn����FYfrw��A���tPN ���m����Ҽ�8��/;:8�:+˴<�;���V^j��۬�˯�M�ȣ�rw$�9���їeEA��gIvwhq��p���ptw�VgݎpE�'6��Ӈ'rO�Y���9NNG)#���N�gE��E9w���_l�mqdQ������k�[��:��� ��g\q�v[j
+�DEvwYq׳vZ�ٛ���Κ7�}�&h'�Z��4.��A]�*�Y�ڷ~���yǛ�$�rh�Iƽ��z�L�@���������G]�cu2�k�I5ɞ�bm6��ٯ���\�kf��$��n���� �F5�&%�w���Ӎ�QH�Q�F&Ƞ�g�uv�r�9�e��["l��+UjITRs�9�݈�AWf����{�h ����	$u�C�李��²�wI'�ܚ����VN^4,>�������¯�{B;{� _��4�1�n
���d�5�+=o�����]0b�Q�j�����^���'"{�Q$1{�kˠ�*�{��`���zn�H8׵`���_U�&�݇��t�0���=���ɀ ���T��c2�z�풬���s([�.7�ד-�հx�"�~�q�3+���b��~Π�eڎF�Y�A�b7p�'!8��q��^�sk�z_���7t��M�iPY���Ƭ|�O?�ޏ;���/&>^>j� �����Pg�h���6�ݗ��@7���r�k�.,gD�-q�f5��|8��AR�ʤ���s5�=�(�m7NN�tf�	�o����7���J�=�΀ˣ�]����{��	K�ߌ^�|*�OZ]@T�w�����`P��.��M���g6��wpb��(�zNh����[���b�pѿOK��k�����	��{w�~�2aQ4.���������U�Ĥ���8VaZ��B�.��t ���n�ٝ��1�:�e���^X+3(�/O�����s��ޭ;��z������;���y�n����)p>܂ޝ���{N��I��$
�x���ͫ���,:�`����n���Yc6�w�m�#�6a(�����ⷺo�zd�܎2�bupUq����tը��GHf;%F���ܻ9Jn�SZ��&ݟCn㞶�lۤwļ���e�n[l���ZM��O����y�g���E�`.��]��-.+;Yy9^nN5�Z�[q�����5m\��7i���L8n;'g�
pm۲�'q;X*�ǜ�n��u@t�<u��u�{3�]�N1�`�n�z<Ʋ�Z赞�56�ѕ5��2-m�V6��`NPi��6!B���켇d�]�ͯ�Ee�j���뚭�s��}�������Xm�lOP���X ����������*V�U&���w3��~��vQ���3�Y��rG�߈?{��t�o�_{\�yow���e�w��&�E�Gk���o��0(OI��AQ`A�|}��π]ｘ�m{��qgMwvG��겱�g�o3B�=���o�[�9�(W��9HX�W�
{�$/5�(PV,��-^���$����9���'r�*+ �?y��{�s����� ���7S3��L�H�Uj�Q
����Z5Tql��J�b�[�-����]٥%���xUHԱ5k��N�3������ʩ����u'd�e���Ș{vy�$y�X���U�I+�������V_��l�50�֠JKX�F��Ҽս{��6��f$�ޙb0�[����&�9��ĺ��Z���S�xAܔ����P�I�Լ��Θ����T(7&�}_O!�]�{XE���t�R{m�6 �_�B������.fk���77I�7٘uڛ�Vj�4.��3��מ��[�Py�T3di� ���劀N�]��򽓆5���B�V]]e�yY�D|s�R�l�6F=�Wv��V��o��4$=y���t�����m��}���AZ��#V	���ʁ7"�ZC����Jb��9����M�Ur���{���7~��kמ�n� (W=I (I=��T_T���e�{1��ky�ii��7�Xॉ�]�O1�H>�qoMs޷o��$KZ�������uٗ��	��]@{�[B�բ�WcG��X&l��I'�c8|O�{kˍ���˯m[L���)m�Ⲡ�2�єk	��d���WT�S`e4��.�\ K��:ڼ79@�I�#mz� h~K��9�L
�p�:�U��wyF�z��?>E'�ئ;bH;��tI��M�JX���k^j�=���,Q7f�n�d~��~��f���e�t �2@y�s`P{�9��z&�s��t�sS�r��#Vȥ��^�X�ꣵ��v�f��#Z��IW��q8�T�.����*�!���i�9�f6�~�7������J�%��\_`��{t��d��h+���-�{�?I��u|}z��q����۠�G��h�+s����t�޴�B��b�]�=��}3�9^�R��,c|��=�~�o����l��1��բ�Wct�+ӱ(;��]r�&���4�Co�� �^��N�Gqx�����s���K��i�fx��,u����x�sVf*�|q�
�N'�e��s��U��瑃K��Y3�����ŉw6U���;FJ�]�η� �|���-����%M�L�z��"y��'�&�f
허9�F��hQB�؅
6�N�P�"V�;�<gE�{N�5�jՙ���֟�)Z�7f�1�����8�I�	�^՟^λX��`���0l[�$-VVK]�=8��iV����O_k���L|�{}̀ ���P�3�l�'����:=��,t3�̲S�=筏����O�p�{֙�y�d$����Ly���n����m[������y3��j�<	�~L
 �_;�@T��߫9�j`����[�4�����J��n`����U0P�Qsgچd����4(h~k(	'����J��s��j�A����5<�n�d�A��V����~�$fs��)K5c�v'h:<B�M�7�vL,���%���2PZ�t,�/9�l%mz�n�۳��[nR'���;<��-�-���Jmu�wgu+���O�1JW��9,Pv�c��N�=�r���;v�����m���J[Kmƫ�چuoWh{��B:P���]'�]�'q!��q�̀�ѳ,���\%q[�h��O'M��u��[uV��|WI:tڹ�[;�n��~&�d���%�W��;j���ki:w����������iq��8�xm�K����v���N�*��b���3��M4��Ҡ)��l�����.�_g�=��$vnY]�o�",_��ѭ'�h-_��[��w/| P����rw� z�nN�r����	n���iF��Մ,/m�5ﺝ �:�p��U��<y�Y�m'����W���D�&���%߼��7
�}7�ԁu�;��~�� �y�(
����i}���G��׳,����M�5F�b�S̜4�<����u?9�!�h���N���&����L�oa ���q��O���ŝ6@p��k���c<�s-\s��멿~���}��`IUZ~<}{�Ay�F����1��O�޺�4#O]�	�n�/��WB«	`��t���p������^�"�{B��)wu-��]��E��F��0�.�dx4��m�E�D�q�R�5�/*��m+X�enC��X?��yɣK��UHQ�jֳ=γۇ_����,Zc���>�ܘ �L1���ܮ�֒w��i?G&o��ݧ
V:9TzN?g=��M�����B��Z
7}̀ ���_�$����79�{1�y�ˎ���(���=o�(�����&
Eϭb�
�~~lP��ﹰ>�Ѭ�L���fθ��{��Y���>�&�؎u��^n$�y.���m'ͺ��,�����S���U�I�f�F�nL߉'�Z�m`>����6G��I��n��i`��Y)*�[���K����$���m� ��}$� ��7t��]j�X�³����Z�QT,U����{�ƟϏٚU��=���d~�Kк{"��W����g>�$Qߝ��pXn�_�>�<��A�p��;��GWs��b�z�b�>ɛ)S���ok'�$���n�A }�����l$��� ݚ5�g{�3=��P�������E;ha wG��;׹���w~�I�����B
=|��sJ���߷r��������f���������bb���n��8��琔��A����;�]=Eh�T�܎S�ܫ������E(�
��T�ɯw�A _maOo����y��޹�y: �c_X��
6Q�HX��=�O�ն���������;�B���?�S��٢yNL
��U���� ��lz�5V> ���A �#ʵ}��z���̀�$[�}M�~�o�fi:�p�TJ�ڒe]�h�{c=��Zٕ��|߷@'�G�I�:͵pfy�m�cM���r�������`�s�o��=�����s��n�W{_���F�|�E+�vq���k�!��>������+�� ��4�8E����u�.��φ`�m�:{���{{� ��L_+}]�a#�~�'�}�����w37���Z#b������Of�b�F���k�ƔR�"i���B�;�(�)SU��xo��Dѹ�I>�L�g�ЏU��g�n
�s4��O4(!DX�@��~���I}w��T��)yO!	��� �7&�$ݾ.�3\n�����v��Tn�.��͛�|�L�I?+í�ʎ*���tPI����A?�Ӹ�{�ԇ>����b}��d�2�}��·<��*z{��>�{�p�F�ĕ���Q��&^��Yˬ�yD�^��!�g`�=C=�9]��o��	�s���ʺ� I_�@�$��$�	/� IQH@��hB����$�	/� I_�H@������%�B��$�	/�$ Ib��%$�	.$	!K��I_�H@��(B��@�$����%��$�	+@�$��b��L���{���=� � ���{ϻ �����>               �T���(�  �H 
�  ��P 
�@PRT�����QJ QV)x���>��[�x�/c�F��Q]{Ƀ�Z��}�xV���A����z=hhi�N��íA�]Ǫ4b�P%.��6ǣN�41�4@P78��]g3(���z/��}l��f�4(u���AN�)[e0�>�@�z�+�i�@�0
^}*���PR"���h(l���F���[0 ^���}�4��(��֍��s`��
)�ԯ|
����� 
�PQ�E�VѦ��=��y��}�}:�:2)���P
�_�@���Ѡ2�`�C{@Pv�/oC�� �G���Η�z��zi1�@�(zm��     �� ����      )��e)UF��     ?L��S�<��� �   ��RaRJ �A� M 2 �S� IT�       ���S	��F�22h�h53Q���x��w�m��յ�"��9k��M�����������
�� 
��6?���*�g����7�?���9����3 �0� (�v��@l�4&Ҩ��x�8�붽�?_��B�*����ӫNxL��d�o���rӎEu���_�kk[m������sߐ
�zq;՜o7j�+�6�)����{�t��)��/*4�/�P������o�@OU�g�d'���Z��(Pl��<��N7��zhw�Ǚ��Pr�wuި��V��#�'w�=ƭM9N=fp�#�J�h�Q6� 6���J..n�z{s�@��X��{�A�5������:���r`�WGg5��G��zR�,�A��;��հ�6X��M���ݽ�e�*���tx8�g/v�ͤ�c V#8�����1���󦑕�+���o��Z�s໹
���^�;h�2M�ۺ �3tu��o"`&e��oU4���k��㨳CK�)���&Gu�÷.�WC(Q-�3���7;��Z�$��f�;��!9�4h �4�
��uj��B��Sz��=�W>�B��8��a�)�ɧTF�����!�}��8t��4��r���]6�ٲ���w��f�   �ћ�p,<�(�2i��ɶ8����h�D0��4��q��v$���Ѹ���|L�ĆD�[�kU��L��I��ې���l�V�JIBn񄛪���oqݤ��&�5(�[��.��t�&�E[��g�G<���::�x^�#�Mok���@=\�x:��ɣ����M�>���5�Z�:�%%Y�T�x6fY2^�h�@�3��I�iCl��{�z֎�[/F����û�p��sBj'�涬����4=[�+�)��k)�v륹�����i�&C�gYŦ9I���o���' ��-帢�܁�d�Y�8��9�(��d��d�Vi��n8��SB��,}�vp�؆�IE;��m�tcZQ�o��:`��В�Om�����E�p��5��ص亹p*�Hn��:�륊����N��;�=X[E�0d��T/^�G���;NU��s�Ś���p�Wn%�Խ�Dj��o7��^-\���L�է<`��Q�����^*;�_K�s��xK{����!K⊦��8�!�4U{*�Z8�9���������{�n{ts��J�bq)O4�m��k5��{;{4�+<~⽝]G��y�15]��\`��B{���q=�s�ü:-ɏ�X�!]��(ݜx�-�yl:=�� 6�Vi�բ(���*��b4��[���{b�N��֏H��Ȓ�!w�38[)*�6D*T�.wEOw�8/c+aس�����
ЕEt��ζ,��z0�N_�yF��*��n�fUB2G�b��u�Gڸ.ؗu��r�W6л`Գ{���;;CS4��ӄ��Δ=6�	B�|5*!S�ǱqJ�y�vΏlKtzW�c�e�m�X�x&:E�'d;P!�X�rk�]�oJ�r���ŏ�׫6ͣ8���
�;P��Vr�-��20�X�P�� {�8���]̈́m�{���b�u����� �c�V��i&d)sj�:��|��897x
��޷��۳i�a����v���;�>�;�k��9L](�WZAwpی۫���nW�̘�!�4� ����0&�ou=�8e��ok��+L"a3�Y{VQu�װ�
\br�C�24��6�`À"yG�E4�vI�:�򜺕�e�ȕ�yP�Tb1ݸD�0-�ӛQ�(�\����*��^�L��)Wv����/ �U�y����&y�֗)Ŋ���ո'ggt��v)Ey݌�Q�S���|���5����^����q�WS�b�ݽ��G$h�'�ŀkX���:n=�T8��{a�E< ��7{���b����.2�GN�X���q�Ą��+����5^\��Ӆ0�6z�5#/͇�f�XST���F�2p�a��FƊ#���q�:;S37v=s깳_,��wd!�}ϷX�.�p��2�4DO&;&8��f��"�h�r&�g���b���Z��{MՆln�&�Y��2d�(0p{�]�/�t�K݆��0�7u
�z3��ܺ��uL�ǵ���Z�U�og|P��f�G���!kH��]ta�-��ǩzìv�k�D�i��)�F�x#B�4a�&mE�6!�t�ԣܺ}�V��\��4��H2%���,b�z�0b׆�,쩵�ۤl��e�i؟4S�Gk�&��^=��4�B;��c6ʎ�{@R��E����H�[�((Y�r�5�5�h"����CF�(�1G�7����iJ��;���	��m�v�V�vB\��;�ҢG���0c���U��zsw��M�U�S�e�w�Ƙ�.�`�:9�I�M��0eHP��N�Ҳr����+SZ.�m�:G������
�`�}N�Ƨ:I�;x�)GI�#qE��%^x���ۧO�N��R�GE��h}�-�T����7S̈́����V.�����x7%Q>�=ɡ�V�<�LFـ\Rt��Hœ*ۚ�s��o\���X ���|ul:D���T�;!F��LC�9n�6���WBZ�f��Vn��a�a$�W=+E�7�gg7�]�*%���M�;���}Y*Ɨron,�#�oo ֭����c?�G�{y�V�q�aҺr�m�Q�sFǁ�
yJ@"}�@�H�d�*!J�� P� B"
(�H  M(-
�@"P(!B!H�R�䢹"�
�B���  d����- "H�@	� � 
�!����x{���nק���fk�*��#���n���߃�NA�- �}GȞG�|?����TjJ�����;`��m��Z&N�����a�6���K(��wD��L^>�J��S���[W����=��K�:��Y���d�����'�9��z�Fg���^��|n�;iP�p�<�Zi��j8�����a�����^��nh�<|22r���w�Δ�fy������-xG�����K�D���\:H{���ݫ�w��j��Vs�l�D	ػ��[��{Oy���w�҄�m�Hz�K;a�3`��ꁌAճ�S�{����@~��c�����9�d��K�W�b:�z��z��SC;ӱf�8d:2|�n�/���_X�+�5�Cվ�*��h����ΎI���Ηvp�����]��U�k�&&tF���B�xM�-β{�V�8c���Ǘ`q �q�Q*�T�E۝Tu�74(��R��3Z\FF�^�;�'ϵ�7~��T�߮?\7\�<�4F�f��?'�e�vv(ԙ�4�ͳf���Z�]@Z	�-[�a�ݷ�XX��5���ˋ������{U����~��Ii��<ᷡ��{=W@͌b��}�*Ov��;��;��]�C��N�M��E�/o,�Aٞ��S�'w�+�v�n:R�E�(�����r�T#�!��#j�u�O��յ�(�eWw�أKyl+Y �޷�G��MX�yu����sw��f�v����a�=�m��><v	���	��5ή���s,�]�<��������qj���a�	���"�f�C�rig��.yV=�H�7���{w��Z��	��'{�����C�k^)�v61助f*1 U�m)ۊn�ho�wp�}�'a�49�F�������0�2(-T����xWk"��YB���nh��cTb��8Rݴs5��@���Yn�u�%ݫ͛%��'��f� »i��>�7)�D��$�}���X�Ӎ����`߽1��V�P�)�h@�y�I�SkvR�W��#��T�8B5[�q�JX\�	�Zo���FS��&s��d�jORw��u��\�L�����G�qv/u�Ӎ5�!��^W~�>�;��0�l7�]�Ǝ���uV��Û��^y�ø��U �Ĥ��u!뻨E���{�y�}�^�\yt}�`����%S`���/���{z�C6��;��[컷i��ܗ.�"��}�����W��]w�CiǬw7��|��+�w����5�e��͹�������b��X������{�G)��s�r��W��/7�S~α�(���z��;`�|��zŸ��ou7rG�������hv]��9$;�f������=��t6��Sz�A�ON�Nw�59QT=�X��yUm{���×�p���O^����y�^�z@�G٭��Q��<�����%ٱ�{�{�|qw��{��*������$�ӤbO\7~c���.G�O��^�ӄ �ǵa'\ro��׾19g�>ɛ�w�՛�z��<�RyT0ZskX��m
=	}ǂ�\[
�~�|�={����)��^����fC���\����p�qa��e�0�#Y�F�����M�LIS쳐�b�~�x�L���#j�.�J��Uz3p�\k�0*np�e��F�����<bm�e���ܷU�BvS�w=7wkE�;s�:65/�g%�G��~e����)�m���ɨ�B��	A�ٻ�� �˧���:t���ʓj2ug�����0u�t�ny<�Q����`�hY0E�iѣR�d\�c׍NA��%7#vjV��mΛZ��]f-&u�Ԝ�#q�������o�&NM�V�5�l#&댴Rg�㯽�σ�%�5��&zc{�^���xpwֹ]�����N?sr 7�yki�Nx�i����\�j�����z�vM�\o$�^��-�w�o����uqP�\�h	7/o,�^k�}鳝��H��摳�,�6��=����{tto>�m��0�{��G�;(�}[���|�����7}���}�J��a/r�K�dO�S��o����������2\k�W��-��j�-㛆d��1��5Z������{$v{�b�m�ߺ�<=s�W��nz�8�C�sK�	ѝ���T�{9�=䅈۫���H��e�"�sK����8S�Ջ�F�_ڃ�x�S�B�SU^Ң�H�
)���Vh*S���t�qQ�#E-�۹�M}�j�=�W̛��wo�x��>
��"<[;Ѹ{Q*hܩmж��D� G�� ]�C��F���SG�|;�KTߊVl$����ٷ
��=������}Sd����9�����ǄC�\>��Ʀ��-��{<�Y������Ӷf���Ϩ�NѴ�;��������>�`�Hm��F�������� |}��:��^��7-[��Dq��HhT/�-x,ݻ�z-[�d��5�cwϨ�x���۸0�-{�)|'ۓ�y�F�7���D�F-Rx�U��|v���N6��#�rg�h�Q�b����a�"��co{�Ob�d�N�"��ogl��އڽ��Ւ賔�t�^;�.��.��gIxƳ�F���=��s�yl���T���F^0zf��j�8�L��t��ʳ\D��zc�N����gKv�<��Eݘ�1�ޗE��B���տw>��z��f(�	�ܝ��a)"�V������PU �J�(sv��ә���M3xYy'����U��F]-k6д��i$�r�������붒��`;g������Y,'��-zNu�;c�k)E�^R囖::ZhME�CڃHqr涣��T�s��2�Ϛs��J۳���xțG���m!���d9��77cp����I�#/!y����ɶ:��k���i'��ͬ���xo0��9;r���t�������N�Ym>�t5ưu�t�����Շ�u���[��8��m3ǧ�1c�O)�۶`��P��L�v2��b�xwV�b��^:Q���h]��m\l�-ۍd:"�c���݌Ǭnv�����y�Z�F0f�A�'�"���=�6�T�� �,�������=�=AzC����8ͦ�ε�j\�Ig3��' q�j���h�xZ[WK7i�0]L;[��rn��ϥ����h9w6�OC����\�n�a��x����{L�1�Ԇ"�4>N{�oT�B�l,u��lgR8U
�k%�S�tF�`�]�.�[���N8:ѝO��:�s7=��ݩ�'��F1��V��t��8nP��+&VL����ˑ�듃ȆT�8�͎������	�Ll��	mkb�֔v��]`�/g��%^�]��7&�O&Ń�ϊ�qqҝxT^�<��ӽwk7����k��Ĵ+��F���w'#^���5э����v-��5\���4v�1ʻ9��Ԋf�]/k��m�s��b��Y1H�0Z�bL�ZR+<�+�1�<�=v8_7c'l@�kr^&kv��J��ίT;u�vI�^�8���@(�.G�\v�����>�^1=�k�3�y���p� �:�����Ġ���v]]����v8��qb�Ӻ�y���ۘ(���&4.�!hao��6�%��"˲e��cWknW#���ת�������,��YM���Q� -��Nm!�`�\����k1ōc�L��c�v;�2�H�#��V�VP
 k�88ܯt�<k��s��:y滃���:�8k)�6�1a�a|sщ���ɗ����	ED3SZ�.Iw"��[sf�3rg���8�̆1�f+��,�2����Se�,�,��j����ui�;[�as��,=T)�Ks�6�ۧ'g�UCVP�6��4�0*�tM�v�rx��Ҽ��1�*r[ư����2�jf�J�h��b��pݲ�9�jg�d0H�D�WX�<+jlʮ	����d{���R ��[[%�s����x�s�ڌ��k��]p���Hɵj��(m�4�,�lW4/k���֍ʑ�-vWsH�M<=\b�;�Ks�al�qo<�!�/F�ݎzǮR���x����݁����q�d�Jl����דsh��ϝ��3ݕń�l� ��r�<�$��tb�8�/c���s�3�5��s���0�J&"J�My�l�v��tXF�]Bš�uآ���=gn�ޖ;Z鎷ic���b���=�u�,!�v�b��a���h�;�ηd�ۂw�u��[���v���ןa�*,)��](.l��R;P&F��]o,������8R9�����n-���I���a��ٰ;�nI����2M�x�m�'nU��!'x^�$6�������1��%���W��>�.�G<��6;q�.,�fw1�;u��u�<vx�yI�r�:.��1�f�d;�ǲ��+'	���]����ܭ�ڶT碭=c��x�٪�j����kf��m���̗3��[k��j������؉9�蹹����n���d��h�M��X�w;-鮻L���k�4�Иf�KM�Ժ;�N��)�=�]XZӷa���nj�㭸��GW[m�'K�X�=p�f�D�r��@q���ڔôf�N`qs�o��mI����Dmuٙ4#��O߭l￿Y?��8&F3D&NfUT.Z���F�716��FC�ı�o�6ؙ���Ym!Z�5�Vc��f���-c�K�)$*!���MB�%[T��TAZUBƠ���m
����(�Wr:j\����b"�X���94�22r��5&�cY��.e�0P�D:�3m�Z1"
+��u��[/2�I��ɸZ�]�����(j94��L�b�n�i��Eة��=;a��`�ut�3ډ�g�6˦m��R�n��6�[2��x��6�l�}���^N:���X0��s��[8��W��I���F	�Se�/W4��U��G=�L�ۢ�uMti�s�fiS��^�דj��>u7"t�l��?��$1���.����u��尔.����.e�bj)f˂.5a���F�SC0�^&��m�bh��3�n-D6MD�P�v3%�v1e[��N4��U`,�ӝA�5[�����YteC�u�����0�&BG3*-�*����&�۩j�Z*�HPRh�q�Z���Ā�ʗ
Wn�E�}�v����.a�%B�`5)-�ţd���� ��cV0��(ʫ`��Kl��x���x�Ĉ��
����2��j0_ݿ��?������yo1�S?9�mL/9�0q8oĞ��*t��j��Ȋ�v��*IN�(`�F�[�
}��N$O�8�W2y�m�{��[b��'t^_�-��<kޞ'�bn�F�/W��,��;[�Úă�3�c���}�{�w��N��2[w�me�{8K1J�>"������7��1�$�N*�+��d��}��������rxqZ@�^�����O�y�������YB�p���@��rl�'���g��SlL�͞t-+�Yt���������(᭺�R.ŋ1��{���8l��kdN���EwUS���2B(h�q������yv^��"7��A�@��"-�B�����tZ� ��;�A�˵~s.\ћN!� Hws�Ê�Q����4�b�TnE���		�hL庄�l3F��`I���XL:����ؖ��&�����<�"�W��hQy�����˷J:���ጕ�5���ˉW�f �$��Xp����2����d���P�%@e�]Ω=a�]Юɼp����mk�yDUnԜ�Ҩ�����S8�6I'iKK�/aS�����w�dd��ᩌ��qKv�6��>�A���� *����,�P=�k�q#�y4p�4�T��xK�^�R�8{��A't�p�D�!��gvE�qT�s58F�|Ťk�v�F��5y�[�����t.���Y��<�� h��4�-���Õ�[���RRw��Go����bit�0�n3B�����6,\�����<%��<�xN���u�&��)o�;�tvܚU��-�����f�	����q]������m�����[e��svP>�a���!8rp�v��FA�/<^DT<��nLO�\M��4Q$2�D���r���f*��D���$��m#q+�)d\����ْ�i@�uʁ#u����F�T�kp�Ba@JjJFָv�VS!�w���_�n�W�E�j�f�i����f��v�mE�r	���j9]�8�7��O��TF�Nl:�x�&����s;�4*��m	Ód!�Jr��Q�B��S����ONy��A����b�GɘKp������_W��"O�;��,`����;c(���Gl�����7��H#HD_&�G�H����,����3=�Q�I�ll>/D��&"+M��`?]z��ݨi�&�����m���ߙ�Kl��;���<Q�K�Ybp�ƍ
ȏYqz����h��V�*�4Q�wN8�H~�{�yg�.���O;�;A�`�1�5�6٫��n�����~���o�z�wZ�^��;�9�y�۩:�{�kJnT�f�魫�ѫs������l'�;��5�n@d�����dU*�	[/V͛����0�q������e�v�a>/�]H��1�kؐ�%m:��&}�o���av�5�0�������8�r�"�D�5���t�1��W�[���g��.k���&PF����',u�HD��=�V�ښ�>�ƭ�G�j���	�W��,�"���q\��J�΋fP�i��Gjzsڨ/ה�o�En\��T�MGe�TfnZ����9�4�!�s�O�;{��Mvd�Ó5s@�i�4%�İ1bY�Kl[�8�6ӌ�ޅn��I�y��ˮrK3�F��u֬��`�1�+���8(�DU����I��WU��M��6IW��oҐD#ة+pْH�L�Q��PE6����8�驦q�w�AD���p�8&�H���,�q{�+�����1�"vI<䞄S�@5�R��6��%6��=��o>�-�Λ$^�-�/#�MЀ�1f�'^q��r�{����7y���S��;[�f̨��	���L�uV�q#%zNA'c��^��߰�o%n�6���jBqn}��˙4���F<:���WfY�A�i ���ש��E!���43w�6Q�~��jme����,�jz��3H?+�9��\EV�=I�<^D�D���
v���>8@��i����]E��~��5w&"o Anq��1گe��pD(50""�5�[����1���^�Uћ�����z�wF��s��0G�-���qO���چ�J�lG X}Ȉ};�i��lk;�b�o�U�4�b5�ٞf��h�,�M�o�w}�]��<j��e�d�e����p��ydU^@zwW�O�����t��J�`��v��a���U;�{��s�j{��j�>��cً_����F�V<�"�p#v�Y�a���t\�|�ݺ���}��"5�Ȳ���Kbw�n�c���]���;S�C ,J��V��jt��ٴ�����F>�e���r�E5Z����$�o U��RB��)jqi�C�!b�",�+$�Q�Z��&��e�2����K1��3�.��і4E�b&AU�م`YFNVٍ�����e�[FU���dPSQ��l�E"FFHƒ�˫�0$� "*�	QP��p�5�Lq���DZ�e�e�ؙe���j����h�jXC,���*�'l3 ȭa�efm���1%*�4"X��M3$H�ZKl��2KfpB�r\!!�b܍;�;��?�"~C��֋q#&U�Y��ϧb|�yz�褵�dQ&5dN����(��^�wz����Kcan���1�B#+�|`��;��6� �	%�	=}%��SAXBQ�5M���lz�T��&�";+�k�Xp�#7BBp�o`��%?.8��N��'�SC�K�1Y���°��zh�{�p7G�z��p��@�^� �Gt����WD��1��}�� �ߨ&5�A�쁏iANR|��FJ#�`�2�0A�=t��w2Z�2U�H6|�ޜ� �sgD�ݢ\EW�)���du8��}�M܈	ðp�	�\.��a� Y���u���!�3�M�m?�5Oz1=�p0�w����A�k�������dO��P��^2�n����[+���0��x�ݘ ��u�.����̏d��Y�ܺ�bFh��&���M)��c�Pv������Oz��_Բ�5˜��8}��.p��Q,��	AMT{�݇�pq"�4�D�Q�+���Q�~��nf#ϲ�a�ҏ�5��3��ã���V�t@V���w(�#1ȅ�ld�O���[��+�qK�Dw^����>��Kn������ڌ$���z&��ʳ����d�дM�Pè����#�)�}�{'�$YDi'��زyez��i��H�1�Tf����	5��]�8�tNq�A(��8�=�{�̟D�4��I��c�3�kBo�(�����#5����6�v.VN��b�M�����Ph�<}�����T �0II���(�R���ur�d��"W2&�MwZ-��g�2��� ~[�ǀC��<ҍ���*�B��m6	���͸s
�F�r�&��6��7 ��O1�M�%N�%���zS'��Y�����#IcZ��L2��{��!����O�#$J�=O�ן\p."kW��h����P|l��v��BӔf!�	���۠A��t���	��9e�WveaGٟ��o��/��'��������V���[1[!8��:��� ��HE9��DH�iv��1q
5��f��v�q��V9���Ͼ��k>�(��	�V�N�#	4G�{�ʈ �΍~�dQQ$�����y���`7{��&�y��$f~/���d�s����>6sh����X��L���Л�JȢ�۽��*�2�$d�9A���G7c�����Ş�j�On���v��Q�G�"��Q`���k\��,����%/8G
qÆܽ�O÷:њ���QM�4,	u���:8��ΐ_u׌�\/���[r�dG���D8�Q1���g�?�%��<�&9�$�	y��t��p�N���'��H�4nF[-׫.QTI�0.Тm�K��%�V�����J�Ȳ�9�I��;̡,�Cx�
�2�f�"m�Yg��'��U5ҳp�Drp��������Mċ���EA�!Y��~"�^;����$UY&���u4���e5Ł���OϘ�<K���Y���C��}�c��Y��xtƾb�3`�^D�@���TA�Tv�@��A�nk��^S����u� Y�&�/����/}�{��xl1����l�1s���g�q=�Km��~�fd�5v�M莬I����Ʀ"�>҉] ���x���iØ^F1�G�ݎ�y�ҡ��*a��%�3�8�tɢ�[|��}z�H����i�Yc��d��܏~�31��8DeG]2.��I �/Q��T�գ�����XFm6(�ۿ=�{��+l��&�Fh�C�Ϫ[=�BYp��DgLt�(���'PD������rMč���!�xf�͋�*�t�HΨD�5j�l`�I3O+�sIS2�U��9F�ꫧM�uu��˹&j8�|8����.&��#҃�9s&!?ayv��϶��"��
P:���(���������y}�u� ���GLݕl0A:�.�5���YJ�I8�"m2A�6Sw,�e	e�@x��]HljB�d���C�I������ f!$U<�WUŠ������`N+�]���A�2����ay�EG|�z��ʤ�(O��m^���{��<Z�=���u<��u7�'g��S3ӐGݽ)� M�[H#fOY�wh׎��3�뇬�U��_<;��;���L���_u���%�C��xѓ'ŭ�{]���5��SXJ=D��w�j~}�+�'�����ZK��φ�Is��b}������)���X��A�:ѶO{Ţ���GJ:�b�br�	L���Ná�!�FE�P�d���:n�ّ�އ���UT�=�4���Mh�)�b�o��͜2gd|��gg<�6�r�����)���lS-7�|_�w�'�
*�Ђ��hk&d��v82�#Q!-�V0�5HZX��V�VkFϬ�oAl	b! �Yyc���&��aku�`n]Ŝh�v��q���YmB�lp��Ke�/��n�üX��]��n��JDY���, ��i�
��!,����B��$l�4�����)YM�[��-K�E�DZ�%7q$muiZ�ae�!��2������r��R�A5�,�ނ�ɱ#�����6�]5�������tX�������َĊ���ڹ�&Z��:�N*m����mn�J�z�4Eʼ�	�f�B�UK�B�V+c�ϐ�-cJ&��/Uo5� �*�rY�4%�"�9�=���޶�8ض��xC��l�c
�gջZ�*l��ϫeM��v¹5��n-��]\��λ]��ȳ �ا�6��a8���3G��ѫ7]'H��Y��L��q��<����v�L��Bl�A���=���6���1���� �Jֺq���gn	w9��.*�9��r����a��nu8ݻ7Mu�Y62'M�ؼ7]bWwQ`.�!Wg�n�#��ۍ����2����ä��5[W]���̹�5�n=/��[u�N7FKmV9-ƴO��n�iBǂZk�q@��r͋,B�A����<Z��4m^�e#�p6\�0��2���U�.����-[�h�`&v������%Hd�,��/Z��M���}������ )��(���8@y�|r�� 屈9��۵W]�һ�,op�?o��5�&J�J]L�{��iWT�e�j�����V��>G3������e��P�^����Xr��^���W;��w�x�fڜ8E�I�n����]���$�I8�NүI�l��\U!�b��i��͖����.�Mte�ǡ��������n�~ }����/��pd��D\=5���?ՂC��I*���#$ !���m�]e��k�����u�"jE��߷5;��Q}喺ݩLf�4L����y�M�q�LEM�gm����q{��x�(l�D�M�I8� �6��kN[��X�M>F50I&�F���x�rfp.������=���I�p�a��������TX��'>A�?�YpF#�:|���M����u��2|�W�!�:��Ҫ�aA�^~;�4ue�祤�� j�(<TŘ������5����nP�NOd13�7`Φq�bZ2I')3����o�t���-��ܱ^;�tM	��������e�d�b"	3�0EbdY"��E����8#1�V��X!�H�?{�����	�l��Ypdh3�9�k?�l���<��G~��{(p��\Y�%v	[��Ã��� ���מd��7Q̓���*D2�"����M*��X��"os��♭�s6gaf�D��
\�{0�Or��;�÷��ױ���5HS9	Ē]��<�8��"1\��� @�H�����!���(��bHT�NN�И9�1�)ɷw��999"_7��*AD��Z�a�q���`d�q�tt�VE)�6�Ӄ�s��	c`ک���r��ص[J�-Κ1��	�X��`�����4�.[����9�^��LI�J�"�y���D��� �s�گ�Q�?�ty���-��C�Z���.���ۗ{U�"���L���P�6z+w Y�"eFi앪��C$Od�"b�`��ܧ+�8:a,q�_ݟ��Ԭ��;annĖ�QG^���D2��c���� �u�uV
E��V!�/�zS����y"�9�v7X�V�3��������X Ϙ��^P�U4(8���g%�H�U��=�h�l�M�f�J.�1-@�,@^/M!�5�hNc�U��l�&�:�5S"�g`�Ⱥ��v�gϺ,h�76S:�l+�����r��fן/8�J���&e�5�#�*�D���HńAA�8r*�9o�2����'
$�Q�LVK���qbp!��6��:�v�s�[�3��L�}�<<���o� ���Pq�_�~܁G��A��˻�T6����"��Lz���k�} �&���sO�M�Y��&�Ggm������E��En/O)7��G��x�!D�Z���"&׌Ww��N-[�뉳���#�}�$�AI�c/��e���%����,�I��k+��W�`��H����(C!�&��*V��gf$/��x�d|Ogh��+R�A�A��C"��*��H{�TBl�Zh@��q1+�����\Ol�����P��� ,��L
��H�B�3g	$� .��	ŎD��k��b���6I97��$e�I')��s���C�^�@F�p��+�"���Yph�l��t�B�@ί0b���p�j��d��iU\L�c�+baZ��K�H��gꪪ(�֯X��۴��l����	�yЎy��]nf�g�v����Aѣ���M0&���Uԇ	���]�\gM8�ҍ�cR����0\��lQ)�~�
#>���r[ �>�s]��Q�UW&F�O�UvB�ƻ����9�-(R�������I�1)Թ	A�߻�C���pߋ��6�)����%D"P�rJ�@��?}����ġJ�rz�
�h�J頉��2�^h@�B�ǟڟ�� �%=��یPlC�d�'LĤ���)Q>�1��y��t�[j5Q���+'��G��8�- q�D$(� �/!D4(R���ġD�瘔�K��>xm	If�nw���雷�:���4�l���ӱ�V��	Fu��A�%.NI�1�Ƣ C�ƃ)�����[J���=���B�)���ADH���}��G�h����M;��*~'����*�Y۝�j��nx�N��:��5	BRw�%&�2�!�����r��ms���7� �w{5��-��(�!B��B�D�J�^{�׳�q8� E9�%	BPj���M�2L;�ߙs7G8�܁��J؄J���(R�ޅ�cA�)��:A�(R���P�
o���~���J��ġk�%
o������l�h�Dh�]Х
U��o�cU�D�J��@����1�q�����r��U6��{��}=���K�щBh�������2�}�J�}���G�P�
P�}�-�M�s:r����>��U�����NىBPF@t톤6,���>�iC��?�߻��8d�q����x�34�=p��k�U�5�%bP�F�����}�{�����p�N�����9�pu� �v]�1��7�Ğ�����fO3���?B��Nӷ�JR�t�ozf�D�^�*�I�p�e�v��x�ʟC/`b�N;�V�2-{۔z�\�E>���;C�b�~����!�]��y�S�s�8}�<����kл=��1���pTb~�-���xBk"�kո����U�a��Z%Q
'�ԥt���[[���S� P��&�4/����w}^�$�	�f'��Ľ�����</r�Y��/��g�778xtڀ��s�7wwhjN��ۍ��aBZI�M��x��y9��x�o�3�z�v���h-��r���K"��`���G$Lb��B�I!	iL���]2��ڤ˳.Z-\���Z](���eȺK��%1�[���bL�"�B�KE���"I�i�h�N�D�bj+3љ�2��ʔ��F�r�Qo4ۗ,��,-��DE!e�[�Nc�Uc��w��|
���Gn�m	K�9H�� �럍"�>�>��?{�3[J���w�-(\h#��J��Nܡj��U�4�5�[F4F��G�\�Q��4Dߠb��Tj4rJ�\�n��uġ@��҅��ġN} ���F���J������/-qsB-ۍ�&739��ן��Z~@�Err\���A�9&I�g]i)5&C�[P���%.Ӓ��o����c��J���(�!Eپ���ZP�Ƃ$�,J��O\�J-* ��M�=�q�����9nn�4m�'� ��J�Hi��F�P�k��=�z�y��1(��� ��J��B�)���fh�z�i�� ��J�����r��bRjL�������/���?�E��Z���2���!f=�K�jr.c��_G�  ��{��"<
}��g}����e�G�(R�HQ$_�iB����GcA���������(|��%'s�����}喙3�ͪMa�e���;���Q��M}��)B��(Z��P�}�[A�h3�����)~�ZP�F��z�D���?^hM�k�1(R���鼪�{PC�Q(��5��ԙ	C��<6��)z�_��Z{�@��o����4cF�bP�@>�-(\h#������J��B�)B������~����Q��O\w\�lMM�	BRt�9NBP�qƍ�)bQ$=����}�|(R��$�|�D����fh�~�ZP�֪5��� �'U�Gd�J�@�amWZ�Tj5Q���+7��w�_u����9�?j���գq��t�d^�Bރ��¨��Mw,�ؖfH^lc{X�wr�^�P�i]�cXu<�uv7���u�n�V�I��g�ڣ��i�S�k�5����zmc!ٱ�<gItX|�X�����-��҅���bP��v�.J����B��65i�(R�(P9�[F�#D���\��ġOni]B5Xk_����(Z�D�@��ZP�ġOv���J�;r��������y�1>��\j�P���Z����s�{S���۪RnI��˦�i�rrOr�bٿ��捥FH�w���s�B�r@/P��q��h"Mn����2N��M�w�mn����סm�!���-�Ѧ��D�@�1*!���(Z��g��� M}f%A�J$�� ���Q��P�
pֿo�vϟE����ە����9�w.�3����3?����#Q���r:q�j�r�9�IBP��������V5��JߡX��?sgv��-(Z>��(�!CT~;��c��Q2��Kﶴ�L>Ŷ]N����Ӟk����9wW�p7熡(J���h�(Jv��j���ڸ���C�#Dߴ{���J�pJ�(Z8�[U�B�ｾ�l�P�
P�� �B�(X�Z-����=̏�4&ҵ�b5G���쪮���)H��b&�o��u��G�ilj%
_�X������y�iBѤ86�BB� n�/��~�g??�=����	F���BP����J��-(Zs�SȾ3$�]����b0�~��3�'����v���	I�5:��(;a���>?~�i(S�2)B��DJ�s�d��@��i�%O�R��!����x��Rd8A�Q7�bP�X�j�p���L�V�?sg4��-(Z<��HQ$^��	��$x�;�FttC1��Ј*�blfzv-ܥ���TҘ��xx���|~���lG+-uؼ4|����A�j��( w�h��
"q�q�$�Ȝ������?y� *c1��5�eq
Gvi��D ���6�ZE�M��L�����C��R� ��Z��k#�s��(����'�5=�o�Hv�#q���Ct�3	�I�o�(��W�_*���Q
���0M��֋z�̬ʱu1����$}Rí��Z��v�(����5�����
Q�iE�K>ej�t��}���뎸|*[�i�	��]0ߏ��[��Ĉ>u�{�/I1��0�m8�p�b��6Im�E���يC���L�n�ҵ?� A�n�͊�d���2��,���7�כk_�ZdHXߍ�ơ9��l*�Uv�hQ��-�? �j}�VX7ve�[r7!��>k���Q�s��n�\qֈ�������N:�D��s�#�A�a��Z �-7Y��u�-7j2�+���Y�B3E":G]��2�{���wS���B$ޡU�6;e��&����l���[*�&���EU�q��2Q �c ����d��&����L�+1��~�d�y���b}�˻��'�t��yz��#��#��������l-�Qв�gb-��s���<��4��9y�x�j`Bl���p]H`�ow�U��`k���ɻ�.b`+g7�{��u� ֶH$���w~��x����gS$�k�3��$\���o6�cq"�$:A��r�d��Cp��L�ׂ����C�\���5���^���&1�DC-%U.M���6�Ͻ=��}ڶْ��F)��QJA�Sg�x�N�(�,"�Q$l�a,N���`�bF����3����!<�M�r^C@���AYR���ŋ�����8�X@���p�I5MJ�%=������9(9Af0ɴi�}/��٨���Jd2C8��M�w�{��]���A ���0�%�,���=!Ú\�me*p�($�@)��jU�sS�p�D�����m�H��08[1#]w^�p�I�A�/aV<��aV��g8�wC��x"�M�Q��w1u�����#�oB?8yQ��J,��Q:�n��~/_�}O�m�F�ɘ�6�5�mDG]���8�D���^,"�#1�w_	�*.�hP"m���A3�v��T��H�lF���s�q��1����2	;͂I����rH`������Rڽ2uf/fdsU	E�f�"��ݨɽ�Ws|���GTM�9�.��n�j-��j�p��oh���S��xOX�s��){�\ޯ%H�{�3������:��ma?�_2�~�7��CU�=>q8�y�=�m��:;�_t.ܚM�t��/g��4v�'iC|�`uK�{ מ�������sڔ�tE=�4	�o'�]d�ՃSV=�)���>�{���{����]���6���Zl�5����Cha�nn˂�֥���ڶ6u�K$�e��&o��	�\�׵��2�
��:���5e'Kfg)�Z�'t���%�+]~�G0�(�m�r-F"4�j"4*�DnJXj]�Ԅ!�#J�Jd�22
�3)�3��10f���c)��KKDhQQ[K�AF��]Z*���+�i�ʳ2,���r�� �l1FIde�X��%Ȫbs������*�0�*����d1n�KZDk�Ȉ�I(/32��B
�p��i��Ѕ�mD%$,ׅ����\f�q�lݮ�,N,���?2��K
�,*2��Y[7v�E�}��ǈ�w����h'���-,s�%�%y��� �Zn8l#�\�OBn}�k�L��vw�-�=lG�ts�a�v�<�8�Rs���pݭ\�X�ũu�f�qu��ъ�MH�.)G��Via�k�|�LX)�[ym�kg�Vm��t[<��S*�a�q����v�g��dwV�[H�x����9xՆ���;�Йm��l��+lr���f��;x�ۥ:�u�Oc/57��݋��jo&v�;:X�L[����a��j� c�����֔Xı"���bK�d
��ջ����/T:s��m1�{�f���F�UUVZ�ڒe�o[qqqԜ�{l����kOg��͏��rN^�u��eF����D:�pq��!7p<Vu蚞@�i�6,�C��%�q����l��Jrd"�Q��&��^wZnԨգZ��3h�[�aX�ٍ\�?����q�U�����pN�U�n&5{Q�\4S������n{��c�jOm���N���7����S���cu;�8�1훯�~?f����}��f��u�4��(e��kG�5:��wS�B�ӈ��K����b�L)�'Q����9�"2^RT�M8n�������^��1�}]3m��G���Ҕ0r!cK�U��Yq@��=]��.@�Oh�Ml&�>U�E@��ZLS)`����]��b�6��~���o�gҜ���z�xֲa���NCck�q]�H�;]�=[������vm��71��76��	2��ʄm�2�ۭπ�;S���|��p�����	�#P�Mk�3��L�]	.6"�{1e���qK��].1�m�lܹ�}������d!X�va���f8�N6(^�J}��n�Nm˲U�q��o7����;�)�n+*%�^T�=��^�2\���a�&.�^gQ,؝�sC6�YD�MK�����g��Ύ7��U;���j�[w����~��k��#
�9�2ۖ�7�����!�VL��i����;mQ�Y��׈����i��dVJ7���Lq*�bg���٨]଼�tɊ�]qŸ٨�"�R#�m�����/��T�pz�N�;�b_����T漿����9�~>@*�-ctŠibb���D�͡�,y�������Cb�<q��ݛ�񕑆1��{n���y��p�qvn�z��vl�]�Z�6,�[Wcyߟ_�}���}b̞�ˊ�'��K�I��^���1���6�M$�TnP��Dq��de��Zu�v���r
��5:�x��̂ƭ���0�f D3��P�!(p�4�:�9�T���Ŏ������G���˚����i��5��.�%�RȒi"af��� �W�(nT���D^�˯���u�4E�s�e)ǘrC�3j��8O!��+ng��"c���vWJ;��L�
5^m�!n�@j�;��͈
��L��h+���B�R�ʜ^�C��Zq�^��n"���S�s�M�ů�Q�p��C6r��6/�L*r��`l�l@w'k���6.�j�~�S��72���@n�ꐍ�����xX׻��/P7�_��gU��]����5+�[��ǂq�ގW�)9�2�T��%`�W���D�3���qZ�f�#Zq>�Q��nP*�z����}%U-���%CG�~����P�ݼ�z+�J�18Ӽ"�o�x|�_m"�I�{��0-�R���ݓ)D��E, ��Q�M6)�m�������'x��@��F��]gBq�U������^����V�@F��W�N!��N�q����ڻ�4�s��ćj1I���S�]�C�f���{u�L�7���Ol9v��� w5OA)��%����\s��4v.�h��:�͋W������b��-c Y���ر���t�.�(xx���^��ܰ�[K1�4�N1�*9!��6���q�w|�q���@u����ߞ�ò����۴�����۽����+dg+"���C�8b1!}����������u^Ems}�(��˧->(�rz��BiZ$�m��k���wߩs��#k��QWY�Ҋq �AS4��8�{�N��b�t���"�'u��	��Z����MI��H�Dv���	�G�x9�>C23+9bH=B�,B'�W5��]޽#���ۙ�e#6�v�!k��L�q���8����	��Un���v��vQ�{��p6��"���5��d,}sj������E�� ���{�_�֦Fﰟp�ꯉ[��X�J�M�4�-'��Ӱw�u�A�~��ǹ�c�t������Ji�3�xn#f����YR]{�v�f�
�H�xd�<�K�����˃�ӛ�]�Χ֟��nhVy��(�0��60�����)W��{}�I��������=���'����K;�{��`�L��wfM��ӉwQc�S�����t�aӝ}�{�<�@]���/�0`��1�# Wg���uzۚA�{�k��Y���Ǝ���|y.�و{�2�2��5����	 -&Y�XI\��RƕS���w�9���q�<��n�q0Q+.�U�Q�F�3.a��(�1�7 ��+��"R�i�`q@%���9Ix�[-�T�e1F:��X�X�k0�DMD1S9QT���҈�S���ERB(-FI��̌��^�|����];\�5��ܶ�`�9<]
�v�NV�y�G�_�?y���w�W�_\K-�tخQ�mC%�U�J��z1{,��['s�+�=���ir��8��ot���s�]����y����o��+X�o)8����wz�ř]3�v��L������ޞ3�5�m���R�p�A�]>��ә8�����U�U��i%ZǠ6cЋ)D}y܊q1���8��*�z	Z#��/V*��,K���r���B5;���oۋmv�#�mUޠ6a�͗���$��������ʲ���IIeZ��Rƈg;V�4��	�1#���5����EV��$�,���I@,:��ks��Wt�#c]ҍ�ݼ�.����%��b�$!�Z��v���z��㬇V,#���r⦠t۴\R�����6��s��{{���=����ǻ���S��@����٨nN�q؛�P��4#�w���*�y�N(NdDr�Cr�v*��uĻ[5��.qf��e#�v��~&a�-����q�e�-����}h���~��E;J�y����%�u�fe�SMW-9vfh�<h�ȼ�ʘ���	����^��q+���S���A�
����KՊ��
����׎�fo�Z�Y�;���;kV�'}�{���{�\�:&�TB�]�G8��l�֯�/1ddu�)��
�z�؊��˓�;5ᐆ]:UD�I��js��\�d�!)������s^Ma��]Ҧh�:���>��hl��)�G]Kb�ջ0pf%a�c�U��Q�PV6<6P�@fAꝮ1�&bpT$�M�
(M8���I�ME�Z����^}XY��g#4<�姽�������n�]�Ew/J�읋S�C���b�]^>.�ӣ�C�ـ�%������fn��;��9W����^|���Bk'�N'e�1���5����Euv���$��g��u����O���hE�6�j'9-S�f��q>���U�C|m?����Y�{�p	JЈ���v�I-��E��г�˨ˡ�8B�FPp���u�S�b�y��E�֮��Y��@�`:�
V��BU��(�5P�	��_g�QT*Y��[*2�c���bn��)�<����s�w5.�5Ӯ{�u�8+\�e��Bx�{mz��l�7��7ge�xe�j�Q+k4�G8e#�]�~}�Ҏ�&��yYh��.X�[
;L)���b�5;;URqb5>q5;�&Z�`c��.Q�eY��u㰝�Ԓ�י(+^uU�N�l��a2L�-�ḁ!������J�V�D�k�H��8ȓ����ǂSfs�7Zt���\2�p?{�S��n 3�d}�`��~�dn�X��'~�%o^&�����9�=���!��ܫL����Y���Ro[�:׿����k����(���%����#*20E͠��Bv��܋�+Wf	��,���%8����m፛�3פ�C�蓷U�PQw@�M=�8Tl�Na�3�>��6c�U��a�B�mf�;�&�5'Ԅr�;[��I�9�n������X��n
��;����xF/u���1eL`-Ĝ]�Q����3=��1#h8rq{4����̐���k�e���՘)��vu�Y�6�XJ���vh[�37֔jd��p�s���>��΂V��hF��~���A_w�ȏ]����m����t��a^Ws-s��瞉��7�/��x�����y4e���'T�J�އ����8v��C1�2�� ��/O1��bR��&�'"�N*���Â^ɦw�|1?����/�w�Z�3������ye.��#a�,�;�	�ѝCm�/��.��ܸF�� ںC�پ���/M���G��'i�tq{y�M�n�Fm��vۻ��;{xE�{�gpؤ���<�]���g�PYa����n��=˰r��NL8�n�ڤ��I���'bwsYcu=�@�����q�k��L6HR=�pAy��Z�@�So�=�^�!���.܌��2�;��if�C�Xu�ny;'vDi�e
�t�ט.��1uݚ��q��<��6,��pT+�w���Y*�Qӑ����p��~��U%=#*h(6�f��Ș���4�4��L��*�U�%]3%Ҋ\%E�T0�-��&ue�"��(CF]�TKq�����iH��.��mI���"ҋ$326�
�"r��,��ʬ��j�Da�ZT\}O9��K��Kl́��K*���u��t��tm���c�u�ь���ݞ��Fآ�����sݧ:�OGe��OW��8i����vu��70�n0�Z�n�bkM(�\����;��X�tnz4��4�)t,�@�@�����pq��чˠ�^�0����P
ͨ��k�L���b�Bĺ䔆�JCp�����Ƚ�6؎puw�fh�n�.]a��#MIC[�5�6�X�E4A�ΰ(�V펊n;.�s���Kn�ڥ7!�d��p'�ysrq��D�4j�[[�gv� ڳ�%�6��`z���j���l�Ϗ0��낚 �m�ja��՚WlV��n�ێ���NB���۶�5U4i�E�e�M�k�!��K��,ń�c�n��./1��ؿ�!:�[մ�LԖk���\������xz��j��1�bk&�饛be�:�ƺ�tO��Υ�GX6�6؄�y�`3n�r=񛳚�eݫ5�ۀ�K�I�$]3�b7����o���M����-D����3lL���֍�]`s���]FMd�z�c�noM�ﻗt�h\'�6��6�'�.vjn�(fN@ή���Tk.�v�K���)�}�����D�^��H|�.#��b3�X9�ё5�\b�*���R��Z\4r�]�wCj����}�Y0)�F�j+*r-fE������#UM��n!���b�re�-��aN��33"yU ��D"�D ��P�*!�j�������吅f^'Q����,'ҽ��y�옝����(�����ޗ��8����7��"����'�+f�
�����}����-��ZQ��R�y�N<��~Z�}�8����	���V�R�ښ�;G�I��N�A2�%��p�1	��q׻��{!{��~�B�>�t1��}����N+��G2;2���V�yV��ӕ��͈���:[#ըe���Ʊ����Ԓ�[�`�m���b������T��_����s*')W}t��B-��n��ܞ��)����Tt�pM�m�������'^
����OV���I��B2��S6f�FPp���Bw��z�����Y"�q�،.��L�����W8���뱼�����U�^��]�Fq���I��MNA�2������T`Y	5cur
��"�f��;�Z�zyܝ��^�rѭx�����6M��6�=��+��K�=3vs<�crʍY�0�����\F�w4�ꪸ�+�9�=B�vQ��%��*�CeM!�Hy�2�4�n��G ��.P�O�eN;�6��Yi�sa8ء����&�~��:���U��*�3u�a���S5�g�k��
ִ���^����(����{24����A���Y!�;w�
Y3������N����Wگ���.���R2�qz��l��I���yU".7��p��	cWWA�-W�����K��`�Y�]�(⋢+;G�c�J��QT�}�Y�����ο_!z����uʋ��b�=�1�3��#;ϻ�J�������q�1��Ι?x?�v���01ļ����'�h�����^�A3�SJ�������)�p�6��ۯ��}|j�+P�U)���07�"�-/tU%H����Y��N!���:�P�]5��r�������sdV���"6h����wm�]V�X����_x{��yF�[Ce+�̶3�^j/��U3z��l�1�i���m7Ci���47q���,�<7S��j����s��-��?wn\Kmg/Z|S�C��?f�3i��o��?oz,pof��կb;�x㧻^�~�q�:p�HDS�y�;��	�Z�^�*e�o�$��{��M��7<���c�\���vt]���7&�g��V��˨t��4C[6�#��1��fL�3{5�b^k綹�P�̏iG.~���>���Z�Z�ϗ�#\����[�]��و��P�v������l!�X1�O�КCc�Xn2N/<�!V9����	�N���h�`f�f!������jAA̷KM�B��f�M���}����ǧ��ls�~[{�B���tȇ
#�?R�d��zw/�rz/<Bla�sX���?�׻��{��`N$�C�^��
1f'�	��=�����嚜���~�B�$Xn:(u!K�Y��j�^�6r>'��^�J��͆���m��[�m��w5�X{'X�C���f���9��Hr��0!�`��9!�W~oߏ�;�S�hl��+f�� r����-D{��+Ă�7!�:͑��Xbt����7'���a��>�'�/5�t�Kj�\]T��Q�(��`���u�]�p3�Ͳ`/�7o�@��D�'w٬�84fo�۩�e�����b7#ַ/U��wr�ñtD�v^끲o}��q/!�%Rycz�,w���q��|V�7T�a��ӊv\8r.����w{w}"���r���u��)"lu9�o���vW�7�z�TX!��w�"Kٯ��gD����>�8{x�C�9޼��u�Yk`��w�C�}�� "��^�F��v]��H[U[�,�W-afd�Y�f�P�"�[�,��"�T�NDPq��EQi�-��r�1DĻ�6E��T���"�b�6��A��A�(���mR�H%�(B��$*E ��.6�j��FEh��4�xxz�O�����p3>�_Dp�@n��\n��፿l'b��Y��ǽ�٣����%m4����a4TGoh��LpK���XmF5���C��<��r3P�HDь�|��S�wL7z"�v��*��0rV^[B1]���:�2�]k�T������D�M[Ge]�� }�Bp:�FY��_d��w���O];�� ��n�t�l쐜76��Co��R�d\/\������ý�E� 2��zO�tHx"F�#P���^�
Ε\�����s�О^�����Z.�;B5Q�XF��Vdd�oF���B��.��<"�`�q��0]ջk-�YC���#Dh��I6 "��T���3�-����CHY�i�jk��ib�PC)#RK۵�7%��P�뗊KM���=���7���4#���-���la�L�n���pQ~݊�f!����Y�;�����4gW��	k�{iV��cu����nk��B{y5jp_7�k���zu�^���C��������vS9�K�)��Ep�c�!���H��}B��qP{A�
��.�Ŕ��;<c���"��k~�5��ud
7����@��*�vs�5de�-�ED��4��L�{wf�H�1��*!eD
�j�8���祉��k���lH�o�g�g���:.�Z�P� �^��c���7��T*f6����{�h�����}�z�p~��n]�BFx~�J.�r��d��MnVDE��[hV٨ޝ��Wm�OJ�RN��>�Y���OS�nU�.yWB��������/��j�J��.��ۉ��U���8#;ws�# ��#g-%7h]�\ `�X��.�E��#{˝u�M��[}>���,�������Q���w�&�	�q����g܆�ߖ-�ԉ�Q���\8�����t��/�jл��r�Vh;z�6��CtUf^�v)�����u��wufc��ݝ9�t�Ӓ!���4v-����Ƿjo+K���9�m
t��g�D)1W��I��~HC"-��"iVaD�t5œa�Ѓ�R���p�u���;������Ŵj�rk�J�劑Ѳ��joKq@����)Y�V;M���6��<��@�����;:5{u\t�-�E9ojD��Cw:�2�D:ΣA��kщ�n��R�B���rr����V���ɢ��w.��������!����H�nn��fmU]3����ϣ���<�'bwy^!���Qj"N.���e���L�J5���q�]�	�k[�������;�^fWOO�dP�W�B�vÕ�Ν��[L�E2�� ���>��"[7|���$�^x]�11�p�7q�DA.Bn+��=�z-���c��G;��������$����8#��Ű����^�q�G���A�܎Ȭ�����]�y1�yP罚��FE��dl����օ�H<�eb��4ˍU8o�N�E�F��H1��0l6R�"!��7;O7'۸��8�'rب���w���i�uGF1|��p���B\�X2=��Dɥ�xV+�������;]�h�{/Т�O�-U������[�������Ϫ�b�:y���z!��d(�6 ����Q�ښq��e_"�+Ө{v���b����j����x-��j�b:�du�b�M ����ʘ����M��bq\L�j e{b4Gr�)��b�z��É�]�����%D�mR�R5�ec�ǝ~��n]�ٶ?/��o�}Ə�㼽Ց��Wf�`�B)IN��}Q\a�!f�Ho����vC}ި��[��{�=�x_n��|h��
W�7T��H�͖���p��o?n��@q��V�,�ID"��DC:UF8��`������Z��x�k�`������%���^�ŏ�\=d��z&�9�t�W�_i��탄�X��|��'��"ӟ����	�^�B�{TOxf�'2}I�_�o�9�MɊ�d��# ���.�$/�^�����zA|B����Q��̭æN�9��h�A$�J�$Ȣ� ��&���& � ��wq^5�k��D�[J����QT���F�"h�hCVHf��QM-fe���
�Y�P�e�TQY4EM3�����21�3��b��-��]�5���T�fUTڇ+3M-F䨑%!��F!η�E���H���Ib��נy��I�wnzz�_.[H���q�lNշ��"]�u���+��6�<8�ᓋx��N�t�xqQ���i��V����vu%%�h�e��坝ǉY:�Fǩ�3�fx�tm�&�ԋK1V
@!�hU��v�f�Pd8�̠L�̰%�;Gr�A9,m��Kt�A;��nw��t�7-��nc>�7N�n8�o^ѣ��m�{K3�4n�c�ƹm�;��V&��2`��,�L�Î������˞������O�l�Vj����F*N]��m�v��	�����wA��0'���Ϋ%��+c���T�iS��gPHФ�u�҃t)�.��=[n��f�]"�N�'9n��4��ĸ+	��,�rkO<���X���6���=�7�ܢ3�U���غx�-�,1�ȓ����x��B��s��s��ckIS]��r=��ĭ�06�k%6��~���z�z�z�Տ(Vt�Ji�k^ʧ�0�_��%==|��{O%����3�{��2о ��8.�5zm{wqq0c1��p��Eޚ���x�#8_@�g�&�2��gU˵×;��{�M��� '##6)��S��'�n$d��fsf6w�&:/�DH��,�՜�qAи�;��8w�}��q��r�	*�	���i�k�����������z���jЍQ�r�*��lvq�/�7��Jh$�aDL�nF֎���6;�U���)cЧ}��ȂH�o����Pn'6�jI�SЉ�׸0�E�Ms�,o_eUm�ANdC�R#-��/W���WE2�8aʻ���d�I�~b��ɖ���c�![q#ea&���u �m�vq���w߷6ѻI�CQu��6o���rzI�������_D��gթ���ê�I�p�'om��V�4z��,0v��QJ��'HP�z�ʲ	�A�k��Xn*�S�<���� ��=}�IS���Jߘe7w�B�lg����L�q�	�B�*����6�CR]�`�fb����L��n����;�ޓ���}փ��<A��#=-���daÛW����`�j��Aӗf�#8�uE}м�]y�Da���=�i��'�ȩ$��ϲ��g_��r#�n&�p$�k�
1�	P��*�u���k��]rͅ��nѣ��	�Vt�1]��}%�����u�v�bK�r��p�ɜh���uc����:��8\�u]��w<s�b[�D�
N���Ϋ%��:�f�3���S��1�_{�����a�ƭz�!w9N@���9�KBq4v�&gr���&	 �6H"q�A����c�i��<`N�"	���ҰI ��3�6
=��K̑�GG^ȱ��1zi��%cd�t��
��Q�A��=��=��}�5�2�T�k�Ҩ��q]y�Ê�@]s$����O�İ��E2�8Q&����ib�n�,����������OL3{v�o+2(@V�$!⣯�U��š8�i2(�C24��Tf7�!s�YbN�,�kI���!�A�a���ê(�H�L�wq�5/e �A�c���o�R$�P��;M�i�ٿ���s��G��W]���z̾X��/�p�qT6�$�\���ݦO�/yE9�ȩؠۂ,���	ku^�NIN�j��c���D��\�4��������e��"����d)�N}�
է�TJt6�dh8B��V×��A��k�$��D��>;�mmw�w��0��]�tH�t��]ô�{��� � ;��+"&�2+��1J��%kzB"�y�ݷ�u;j}DÉ��ô)�������wX`��u�Bn$�ݪ����"�}�6�*+'���]j/���:��7�v���+b���J�$�9ڐ���MK�g�� #u[�!A���4�6֎���
}���α28�s��uW��[1p/K�EYq���u6�9{��QTG2�1QqA3H?>}�dÉ�V�G-2N L��QqndY�l�TPM��d"Lj��>�$G?qH'y�C�����r����lA�%�}QI�Mg~�ν�^<�����~ɧ����V�lX0�5k�xq%Y�Ր�������I�4�Nx��m�2sm�\���9�Wb;�������Q97։�j��%�a�h�n����mv�-M��5pn/�t�$Im��x�Hy�#��E\5��>���':X �Ak_�s̷u���Q	�J�k��$��9�י)��Eg��w4� >PI��-0/��(�q5��$��PH��s>�qc�y{����v�-m����ˬ���s3�{���|�r���8�{��إ�8��l�Q.���fuٝCs.gU�Ӿr�if��~�j�R[G��ն}<�c�O���`,��Q$N�0Nm#���I�:�q"�S��D���j���Sg)A&�)5F�DaG3����hg�7-�t�t4�)����U��0�X�)��w���y��݊���ޤ<Nri�rk�^/�����g���l_A� �E?ӫɞ��a����+�SP��{��hPẘ�+߻���x�>��%�@�����O�}��Ć<P>��Þ�^e�Z�w�뺳���2�� g��ph�Sv�U5�.SfX�^�+鹧}��ɦ��l>�x79�E�J��.q��"�^6u��f�;pn#C��c���xZ����m1ժ�zv���ɡ4�OuoyNθ.OY�v<��YNɎ�ʥHw%�MD��x�]:,�̣7��;�C=庽tԲy%�m�����{n���0'��Y.�a���
i����\~�ysp�b�j�+n�dE�)��-#�
"ж����\Q�阐T��ʩc�%&�(�"
��¨2h6���2�"�mA	"���B �X�E�\�-"-R��D��NTd��d��TN�Ȥ�0Ɗ\�6�Tj���' ��,����5%�ruh"�M��-$�7��Ay%������lu���`�U�/K�lH;F΍2�m2I��M�eIn��뼠�dGhJ�t�˝��{��q'D8ٙD�VYR�2|��l�qY(X �������V�C͡N+�n��p88�#P�^�"@�M��`j*��ٹ�� ����d���ME�Qz���l�e�(د=
)D(P�(A�O\K��ĵ�,.��z�R����RqZ�B���I��;���.�6�n��g��~��K-�	$�|�q�;"�ܿWd���l�i���U ���1 �6L8��`�+u�[ cB�nye��D1��A�2��[�ņ:Xj$l�`�1�,-�A3k�|�UO�nL4xw��ܻ��F�z��o��&����#�����u����\\��a�9k�<�&z����u)��Ćfv��ye4�D;q��Yw^�8L:��F�.��X�d�u�k�IK��-5�ŗb����{���I3͂H�6��i2H�n6pq4d���=HX"9	����nY�E��%Z�>u���ug�-�	�}�dÉ�W�"�N ��G�0�7i�;�r�:�Q������Y�QC|�O>è���Ãl;��n����v��W�"J>>�bA�RjP`��Ra\5��Z�M�sL��^�'X#nwnG�T��P�2m&R~���=�!��dƈt\��7��tt/0o�X�"���%w�i���}���۬MR��`�r��]�R�IH�٢a�\�`��zT�>@� ��n+�W�Jpa��B����B�2D)����a��!LZ�IT�u8"��L�5���=I��Qq	]�Ίiv�ذbu0��^$:�dO�.�U�ݲ5Ꙙ�b4��
��UA������0}Vَ�|U= ����wS#}e&-{2䵺0C� 筱���s?.8@Z��[��ࡺ�e���7ϯ���q]���r�#E�9�u���u�M���p��/��u�錁�J$\�`�>Dˎr�NZ>WԠ,�/�=��.��I<@B���s!j�5���u̴w춽��֢��m/�n���K���w^�#�e1�M�(d&ne���� *�3�d6�(4L#*7;GV��_}�6��s����!�@7k�ד�&V�Sy��O�Pkˣamk��kv(&�ɲ� �&}r�cc�H"I�l��a(���}��ă�"6S ���[��$���@WjD��̭B$�A���[����i��1{�*����n4�Z��ʷ-~��@�Jz�	n����
��;y!����5��t�5p��3������f���v7����/m^����e0��V!����u��0��]�cA�&Λl�������f��_q���+��Ѡ�hG�VQ�A�F:0��YH2&�����E����������b�K�"7W��Ok"�N�Ի6���y�j���0�ϴg:EGi��(��K��y�����G'����zŕ�l�kNgf��]���y�v�g���v�����>�N*�qTd�N��i�]�!Ы�lK���Tc���
#:��i�F�+u�F��7nȎY �v����d�����^���
���wp(�P&�F��6,��k���+:|�j�C�������7ޏҺ�u\[H�D�D&����k�����et(.����l��:!�ka�FS���`�-:�q�/��d�|I�L��+;
�Wsm�W8;�CmZ��]� crF6fj�TG��$�ɵZ*A�q�����o[$��k:E��fgQ��	;L1L&N/#v�"鹉���~N��6��R�r�l����}�
p��D���RN��h"M�f�EXJ$d�d�V��#%���69���	5٧�*!�VHEV�t��xޡ����5�l��3ptB=n~��7o��l��k}x׋���-l�m^�ޠ��"Y�2
��'H�kP��D���>/.J}Y��l �5(��mc������m��>�Ύwf����b HS��V�(�s{��'#�AZ���i��zN�jr��E~���O�&m�'ݔٷ�YfC-�Jm���O�Ngً.�^ ��,X�^�m��Qq��}Ǭ���*=0�*��時�*����!TO���AT�����3͌s�w�a�����v7�۬���o��vD]��T 06�;���7�q�;o�x�\����Ԋ�����{�/�}8�q��N���ۣ����شz,�ly윿�s09q���8�ڹ�/ ŷ4������ˠ�
��'_�}:w���o� ���TU?�C ����4��=�o��������� ��������?��{?#�n�<����*����������MC�q��so�tA��p���M�蟠��������'3�����;�o��q������Ъ
��{�t�x�~��G��AEϺ� ���U)�q�Foᜥ�k���9��xv�c��AT�����<���3n��~�vL��ǚl��m���W�z�}������|�r��;�pUS�Ǯ6��?��ڟ��xz�����q���4�\@��v|}����}�n�K���>�a�xk�����?��|PU=O��n~�?X��}�}ӟ7w��?�0��|��`� (�n�}�*����c���߆X�Z��]��r7�n?�p��DU8V����:/�������`�r!|�@�7����K�e��u�Cw�i8���3�#}͹�0?i��
�GA�����_4�EAT���?&�>�P�~g��?������:�a�>��M|=�a�lo�z���__os��I���!��)�����~��b*
��|_-�O+��i�b���4��TL_�p��nn�����t��c��:��;�@�����8�9��L>��iu{s���1�|�t��П��y���~���ON��o������{����Opr��K^���9���G����W�{����y�7���q~���	(����A���=O/Og�����|�jx���_��}ۇ�!�-|t�5��������ۺ=��O���"�(H>h�5 