BZh91AY&SY��{��߀`qc����� ?���b?~| �Е���Ғ�Q�h��D��k��d��F�V�U$T��`b���Q6i�R���b $�P�)B�R͒�ٺ�TMwgYF�IY�f���E6b[VZ�Vd��֖�i%h�5�,��͵�HeZЦ)���)��mIKV�1J�"�@7�sԞV�ZՃZ�6�QV�Ʃk-	m�4%�ZڭlԂ��d�ֶ����[l�+i�ѵm���e�h�,U�6���e��-c3k,���N٢�%�x   ,�n���Cu�u�k
=��mj���z׫�ӏz�N�/^컚�zm�j�\w�k��^��{ݙ��sl��T���{{��Ύ�����RjԱf��f�kEc6�Z�   �}�T�J�w��{��EJ��q����J�����*��'z���T�RU�^��
t2�y��R��Y��zU��!�P	n��=)T�y�M[h�m���XHfڶ�   �{�T�ȝ�ü�)B����z��T(y��J��=<=�R�*[�ׇ��
9��J�79T�T�ޝ�R�����J	T���j�[D�[h4�mZ�5���  �U֕�ҩ�)���J������h/y��"�hR�Wxv���l���ҤJ���7A*��z�o�TV;��*J���V�U��U.�V�L��J�U�2��lk�  ��UR��ʷ�k��eQ[b���{װ5R�.�%!AR����w�s�m!B3��ڙ�<7�Х]�������pwU��S�Z�i6�5�E�cm�֥
�  ����_Z�q���=t�]��^�J�8:�T%RC:;�Y*��l:�J{aj��/<�^�`���x���T����KM
Jއ=�m�W�{M�ei��jf��M���+�  ���
��.����.�T-�Ͱ
^��z�ʔ���{\==4�
����SM	)y��BJ��a�u�V�W���e�TU����^�U׳���U���l�P�,��  ��D=��� �q�^��� ���@���^� ���yA@��=
Cw��װ�Ѯ���=+�&�Rzy�(����V��Y��PP��  Ϗ��E����]ޱ�T����=*��W� �[һ���48�B�����Q�T:�yq�B
�y����k+Z�b�Fl$|  ��� ���T �w��������@{ך��B�o#t��gGp
QW����
)w����Y[����C� � T�&�R�Q�р�1i�L��{M�(����F  �����U?T       �~%*T       56�ARR��I��  &���CH�#j��54�='�������I�}�������sG����H*ʻ�j�U����l�q�!�*3p�,�����=�g�yEp"

��DU�����eTW�g���+����C������?��0TTV�U_�����g�?�Q_��}?oPO�%���$"�Q"��H� �(?�J!�?y �*��(�"� �� �"B>HA>H>I< T�!�%D�!D� Q� �!A�%@�%� ���*�ԅ�H	�!Ċ?r� ��H"�('܄H�UO�  ?r>I�$C�PO�P>I@T�!T~�"�|� ��J(��!�J�'� �|���H��(�$�$��O�P���! �% �%���}�{�O'�}Ͻ�M�k�]�s�.]��iۊ�J�$U�&�YF��,����Uv�)�*PX!����ä%�V�Ӄ�<YF�3I�S�[�o6�p�p��b����q��,�ݖ0b�҈��8k%�	\�è2S����Y�[5	tmZ�@��BR�GL��P%�Qg��:�Y�Lz�6v��oDj:�&Еv���I[*�$u�P1ǅn�C��XR�mX�0�Ԏ�Kۑ�%�[1�����.�^��Mn����ɷ�(���05�!�d5r��E���gVz4c�E�ݩ�"lhX����r�bڙ@@��:� �3
5(Ón|��^eEXVҘ��@�n$��HZ��2����*Ql4�S%V�u��8Ca���tT� n�4�n^Bee�G6^-��V�E���,J4E�ׄ�r��x�E{��FC�*�&���m��r��3`X�sN��(۠�j�,d��6j�˓s*?��WF5M���Ǳ%-�G6	7N@2��em�����ڤ.�C76�Y��Mȭ�������1�тrX_-j������T���gQ}K�;�1qe��ܦz�%W[���f�yW��}��E�
�#�2�c�l�N�+7�������+yͥm*O2�4��e^�ڂ�3[v�˅Vޖ��#,�!n�R�;t�;�^���8d�V���-�L庺� :6��ژ �E�jʺ2:[ʹ���� ��C01�B�v�E��F0j]n����F�Nbx2<f�^�f��#L��i�����,|5m��	� ���v���ov�L�ŧ�<*�����7S}�^#���ö�
ze�{)RVA�F�U�����4��$��"�؆�6�	��Q^Y!i:m�
�c[l2�`A���Ź�Ԅn�r[��@У��	�.e��iLِ
vgۈ�k#�d#�*�Jg������{g,�����L��t�$�"��Q�<��fT�{L���Ƒu3�����ڴo�)��Ґ[�"�l�Sb�/e�]�"{T]bl����o U�*�(�`�l�f�[�f%�A�M�C�v�#�������6������缪�:m5c4P;�(�E�4�Ek懹��٬�k���+@���9�ޙ�#�)q��+X֍�mݖ�iI�DT�;���Z��!b��n��kK��z��.��8�+G�)������#�8�ܨS�����A��$���ț�Ա���7H]��jn�O鈋�A�"�N�̉J+�57F�ݝ̡��u&��J�˸�bF\�cQ�
��� R����tC%nkf�=�)�؉d��lob��(��V��OE�{���R�HQ˟	�f�P����vY�f�6��H.�4�d�%R�[�R�&i��_cnE1Mt�Zu)݁�/R4�F�p���D]��]^��r��2�a�4�e)Bc�bc��5�Yw_]wp��Y�
ka+C�b��&M�N@����ث����ě�c*���CD�0����ۻN�{q�e�=����څf�z!KM���H!�����������Q�t&Qhz��N���i��U,%��]�) +��
s�����5a���,��tk��ˉ�y�Ph�����S���4�p<�fb��&fe���y&3t�3$-K�R:/f>�/!r�4�t��ױV�B��Fm�\r0�i�s�(�cvoi=ߠh�&�va�$NV�"1�I��]m�U�B�8�룋��/_WS
�}�6)<.n�]z���jJ�0ʂ��Ì-�!��	z�j�.iձ�%��ݤ�4�Y@sh�
Q=��{ZZ�4���m������v@����i5�& �2±���ZL�yH�&�QT,u.;V�eRU��䨑|1��!����f�V�V��)���t�V���#`Ks$[�2��r�e;��h�śz��n��9��p��i�s6��@��O	���)]'�wnm�h�:4�
ϐ��d���,�B��eX�sx��e�s�V�1d�R�+��l|p1���p^m�e�$
��eQ�+*����l.dYd�H1P���
:�:��Iև�;�@�Sb�f"T�Q���4��v����wn[�d���Ŭj̃U��ʵr͌����c��U��Ù.�Q/D�p�ƯRf��D��bMM�0�����3hY[{��
�1�LM*��lb܂��m#8&a�k�o�!OB���k[��[;��$�hm$�-�G��-��ֱ�yb���`����0U�Yb��-n=ǘì!n�F�>[K��U��<ץ�1���ĺ�i�ӬM�R���
����so��j;R�6���P�Yb�j6��:��I�
��d�n[@Z��pK"P5��PMs��������
�wj$���Y�Mn�n�շ���C �YcZں�Pҭ��W{4mʘ�3l�OjG�Q�x����{P�v���HX��f�9W 7sJ� ���f�(�*d-���Tv��pM #��ܭWi���*����ֆA,�[o��d����`�����\W�-U�j��SE�kw;��Ǖ���㥷le[m��r�6�nlYxY��ȶ�t����X�C�ɴ��VTEL�@�eލ��O�4�&��u�[!TwR.E�����46у1Iwu���5"�EG];����!,��7�6R7��'���� ,I`�@�n3 ݩ��RG`�K]+zV�,�l�n)�8�����Y���]�J������2vݔJV�mP�Tȍm쬰)CP�J9�*-+�[������ej��L��CQdjVQ���B��e*Q��H�u�Z�v���e�)�)a�e]XX5*���Ȇ�t���Qg"CR�7yY�Q�f�S��/�_hb�(����0мnh���ݛP�=9n�ܣ��o  Fg�����#z�͉+wY:Ɨcw	Gc�W��tֽ$ۅ�O��*�!z��fȮ��k5]��IL%�ٸ]��|�ͭ[e6Z����yOd�vd��j��X�f�E*U���Oce�ݕ0��%Cj�O�t��[��e7]*i���j�����K*��զ�Z07wJ�ݚ+5je���h��{(ڏ&�J4jU� T�]�� �i�[�-,�x-QD9�V��)�/qԦ3.���˪#;01��6��,f��pS��^VL��U���3N�OBY�J�iP,��K̭�w�ij���}$y�a�*�<kH;�ye������Đ�Ņ|��N���`�T�ʳ&u��ʫU������jFG�wO"Y�cϛ�v3 ���\$e(ȼ���f�Ǌ�N�S�ۛq]ғ�Joa��]kM
ɡ�ը|]զ�����h�i-Ƀ0B� DU lNS>�u���>&%��e�y)��ZG%1[��J�L��Xp�:el��*���1wI��L�VO�s;�AtA��iu�l�.k.��n,���j�����ю�b٘&�R���AՂՕ"���ɫ,޻��Ou�͢c���Vn��"��m)*���kD�v&�4lʇ/�QiԚ(��W5�F:����)B�&=U�i���B�����V4�q�U(Ǜ��v�Ѹtd�0Z�Me葱W$��N7�� �km&��R0E���d����JBnB�V�-�Z��e�-fIf���n�46��>K.f��Ksٴ�n�%+v�4sej�h܂ƃ1=u�q;��*K���kw!�6�v�f�h�O(^��d�I�D�!�[ջ���Ҥ�id�����-�Q�`����-dph���RA�!�L�T葇\�u���@i�R����(�wX`�-T�;�d������*�w��鋭�&����¶&�ժ�c��eB���v�AQw��� ��0i$n�#,���c,�@�-U����A�e%n���F�	YXO��4�eљD�f�e[�6�8Jy}��P���s�3u@�C����K;vuM�6�V�.3��Vv��R�)�䉽�Z�QEF�<�hc&��A�����ZA�{x½Mn-�}��5˩���"�Ok2hp�A!�,��j�V�f�q���Ǵ�f=6(%��YN�T3Q[�N�fV�4�����/M�H\E���YX�_L�*jJ�ȇ��c�i�	���١&j֒�M5�W�])��F昆ꅼ
[ܫ��0L��j��[�!dɡ*tżÎ0����I��Dj�aC���!�#�u��+Kk!��MO�r�ަE]���4FR�.�w�V�����hn[,fm���&�k1�*T?���U�,�2jn�e�t]g�^��10b�M�Xy�C�%͚�j5�fk7Pf�Gn��m���M�f ����hE�M�)�lX2Jw"�_ۧ��n�NG�9�Z$�6�6�цd�*�:�!���V����[������F-۽�)�w�07�꺘�!15aI2U��I`;�Y�@JK�sro��ih�zHL�xɿ,{� ��|�$ՎoJ�؞�|�:B���/������ݺ*�y)�͉NC�9��	@̀�L]M��V�h�n� ʒ\�v�hE����6i�s7,9�y�i�3v=*ʺ	�Nk�A\����xjen�ɷZ޼�%� �Z�p��f��X�N.7f�#��3(���"��
Yt~jR5r�$ʡ��'��+s�U�kջ7p1mY��y�n�1j��ֳLbմ>�����y�(uXh�-ಊ5ڨ[a-|3$���lr駨�JQΆc�@�C���/J�2U�� A*�767L�KM3Mae��u�0�4��j��Q��5CV7PDъ�屮������-��y�g�J�,��J_&������Y��n%�K82J��:�vdˬ;�]���6��`J�@�Z����tZg(��̐F�-��A��b@욎���&k��ucKŴtV�,co"{�P��W���M��fm�eB*+��]	.G��Qk�P�H��r+:	�m��>�7v%��ՙ�+E8���nAi ��v��(��s����f%�%��3u5�bl]X��sU��Ei���U�C�Z⧈dm��K^m����:��h5�2�ֆ���٫7.�
ƀ+*c�-�n�壯2�\۬��W�`����RB�`yK
6ұ��e�朽�r=%�kf�U������%e��2�c�o-�RbC�+�v@+-�F;�t�����Pf0�GQ���\�--O���/
x�S�^ݬ͵��u.ViH�n�w{[��ƭ��^d�d��t7$�i�b:E[Ĕjf�9t���j�!f���x����n��.<ʘEX5��YZv�q�j	XvΖeR�҄�4�Dؖ��i@m�s+)��V��YS3C���[n�	�f����{
������V�\p�*�#�8�f��<��gI�d�S��]�gNY����r#w������2j�X\���<�z1�^ ːb�
�Sv���f�ե�,熦s5�����!��4M1��bM���X�Y�YX���;��Ֆ�C��&�p��YL�n�"x��!,B�ǳ76����]0�˨���p��ziF�g�n�\#`�yh�e�Z�	�+N���Ƅ���&fX��O4��h�%�c�,��V�
db�o0f���y��Z��j��u�Zb�S���-���.��'(��Oh�����p�F��e�V�m^�,���ś[�>Đ�#��O�t���[�gMsS��f�*�h�ĳ(����,��I���j���m�;l[z����\I��tp�fͲ��7Z�=��7 [�+J̱�F�[Q�	�[2�%��5m��ݏ%�2�v$�f�{u�� XӇ30Vey�c`9�h&�YY ����\ørP�� �Y��-]��j�JyZ���H�o�>h*�@B�����ͱ�t��&�m��n�c�l������O%�Y�E�W��[Q&�W�����֨
�j7����w�s4���t���t=9$u�&ۭ'.�%
�
���ͦ�h���bQõJ�F�	RǷyX*"0��������I" V���6ݒ��h��/r�z��Z(�ہ��8L�k͡����.R�6�Q��([!bجl�y�=z�ce�T�]����-�TL��cV����e�[P7Vv�#��ȥ�D�P�О6��ԮJ9xmŀ3�6؂Q;�X�35�m�Nn����!ћ��d���r�XߦP���Ղ��qBV:%32�� ��H.nVI��&�տk���5%q���5�7�w��Ȋ{�� �ߞ�[5Iz�/0�eJ�� Cffi����(݃[�rܙA��!�֝���r�-1�r$G%&������IR�:���d/(*��f�����jd5�6l):l*��D٥4᦭��U�>Qe�Ǥ4D�AbY#V]*w ���xe��x*��ݍ[�%�{��0�Reڤ�z�,#���2�X�:�ю]��
`\!�P������P�ͻ*�	l��r&�B�5�����B�7���o~�V�a���:���\Wg��;�5}��m�1��	��݄��'��=�-^`HH(��M
�"�������i�Rhߓ�hS��Z���2,M�-����`33U��I�G6�DI�ۃ$v���D�S+h	V�3�R2��E%�wl
'�%�ofŷ\5�4�Ͷ�`j�@����!v�T[���Ư����z1Vepc7I���m�u����v�-Ņj�������WB|[;�u�xF��&��P���Vh�@�Y1���%��CpZ�m��k����^�Ӯ�b��
��I�Ό;-i�4v��E�ţ5��h�R�t­bZR2�L-#v�����oA](�.q�t�waXd�|��
��H����ĭE�U5���s+�@,���.-�a��?�>��Ʉ�yz�܀��c�_7��r�*�fAr3�Ǜ�Ct�R��%��U��6c��nr[�}5�Ð\DK�,O6m�)�+G�1*�u�O�̣��Z�`"�-��+"crʛJ�,��3e�.���Q��Z�����;��}ԍi��%g,s�+&ͭ�7kU�B��gi�q
�.����S�պ}{��H�d�i��� f���8� v��2oG�1H���?{�A&�I��~�>��bĝ�zRu�g+e���c}F��=	Ыna����k53��N�k7+�<ɖ���`l��U�VR?H�r�3ܮ�5�U�8�ċ�ڦWC�rcQ�,c;��eۏZ�������\��g��+{6+�V��&��+�ЖY�$�IU�!�M�|j�N�tcP���Ș[Y���Y#x�
��4���<9vD��,�L�a-�T��8A�4*dcՠ��k7�L�:�����B�G)����D�w:%n��;�ǘa��5�4���Ūc�[8�'x%��l�"cw�K���7��t;#S�a͙9v�:�}	�����u�:h��qd��,�vT��g.�w!]���t@�{�jue^<G�l+�BP/����ͽ'� ��Z�T8�i���G	B�*�Im�j�Zn�<LR�髦��j��n�~ו��G��`[��^֋"�	�,"��vYiK��/ \�LC��7G���N�S�#X��1��m 4P�����՘q�K��E'Onp��a���LT�M��Z:wt��B<G��ν��]�`^N�]���R���Э�b����Ďӗ��@(:��s��WwVZ���s,�M>1�{��t��ˈ�S�2*u�|��R�:b��6-�u������a��1r�%V$;Gn���`�������N=�K�Ñ�\�}�U��B\2,�IN��=w�mIK�`U�:P˧w�i�����Ooxc�N��@�m<F ���>�f�^N7�Lc[sWr�Sf4�E���r1h��Mhָ��*�pLƳ�]����E�똜(8ˡ�Kj�UK�͉�0)D/S��g9�v��(=���8�RS�')[{�`Q���z��ft��v�×f���8G�0�wQ� �J]�} ph����d�gSR��;o���˘r��闦����ٙ��	Lf�#:%��<����l�T��[�^�u��F��%LJ��R�r�y�!��`�{�������E]�#۬��]v�v���}o
dd7�+�m�BIMuܹ����Z:�1S�5�N,��@ 8p��e�m��y�X��p��W¹^��X��ªn�t��}d�*rqb�kV�[!�Q�z��|�ƅn'�P�6��Ac:��B�b���Β�N�C�/��[M��F���1Xk���f4�ל�W[贁�%�9(T���^�`廘�ǟ�%he�WX�9L#�Z�g`t�:V��6��8��J!��w����h����U�Ƕ�ֆ�r[���2w�v�A��tRR���ޓM�s U�V�}��Z��T.��h���4�]��x2�V���"�*�x)��<ɬ��)�#�휒�d�d���-����WF��̫L;�[��܂���J9>�����TtnS�|�	�ڟβX`�%� $5V�+���xhxU��O6��^�&i��GZK��p��,:�3�cֵ�Bw+5'[n�l��\�k���y��E��D��ъ��]��35���E:s1۝*�*�s]��5�Ke�E�nq/_4 ��`�3��7ЫF�Ź�nތ���u).��zwR:pq�mI[�#�CʦX�(�dJ�U�>��]��y�Xe̷ݤi�7�l�ͅ��՜}�|�=� 6�i�%@-�K���p��j����Z��d��r�� L��=6B�N��R��(�5�(��$��R��`P�z�ʔ۽aX���Bnł��*Z�Q	���Ԯ�v7�8�5z�[����.��̕�Lj�,2Ҧ�Z�U:w9��lf���ӛjFm��際��V�()���Ѿ�Ww 0g<B�t��Lٓk��іn������O{�Һ_d��x�W\���3RrE�2wtΓWf[��
��:ܔ_�̀#�5S�(��v�՛��oQN�����Xj]���*��;kU��� /s������:�[v�\�-���v�b���@V�9���|Xb
ۙTŸ�Y�o�7��!X�bKT�:a�e��ˠo�=%Pq��I|r`�e<��$��B�:6M:i!�n���1c�ܤ���,Wb{;�V�24 -'
�*g�7k
�Ε:�:._3]j%`ա���ljǠEkv�����%�I6Nr�����dj�z<�R��6�r�����M74 u=�b�!�3���wHbt�!��]���:�[fl�/��O����$��`�]`V.�`��u����ܢU�I5��P+��$L䳃�ucU.=uu��R�]rV��[
ɪ}�����e��3/:��mA�qe���9\n.w1�Aj�J�Vd�y�1� ְ��Y5��0�5�+)�	��P��jLT��{ ��+&�5�<��X��i��V�w)�Ďl�$vG���-ɵ�C ���1\�U|8��ǽ�t��~����gfWCQ,y;�FD����%��66uͥ�V�J�˾a����X��j�	�[��xg>���q��#`eۮ�����]�@��-�ͥe��"Y/f�5�%e��#5�����V:ɫsh���	\�c�A�մ1���$EkQw+c���\�n�s"�����1Qg>�'Ec� O(P�;���H�՛Z32l�j
.�1 ��x 1��P��\��Rn������<�+���xlD8�\z���o�q+K�o3��I]�u���Rz��z5/�[�����C]~*�����i�J���jN���]S*&!��3(R}U.��)J;Yw��%�}YB�t�����X+^�`7�P�ۜv>�W&ˈ�J�îXu�ެ���w&PwS����9�<��0T���{i���q\��<��C)��kLFq�j��;�,̆f�d���f<U.��q���*��\`���ћ5�7Y�!R�n�ƶ�ԧ[���d;��rB'�B�.$D����JL:���k��+>w�3�i�'�ts�����ræI��Yz� �W4�c2��Zi7����bb��
y��Rڔ7l��Ls���&�_iu��R�%�9X��!f�|�u��`�o�����]v,����Ѹ�n��:dՑV
�}�f�cChf��j%{c���$�{Y�i}��,�y��,�E��kt[���9.t�)��զ^S[�[�\ݰ��Uh�9��&����pv1Hr��5���c�no]��p�l`�v�n�J�f��sz�q���{a��M���Z�m���[�kœV���œ#��Z�Eu��<�\i!�[Fվ�y�lch�`�X�Fd�Cw����F0��2�B��+�C��j����j��2��q�(�l�5¸�vj<��wM�7M<���Qu��fr��НM�Y�z��e���k�H6�k����LU��O��h ����]g^$nf�,-�7�X�7���wQ���\�|v�`foϯYN1���W���TAN��C{k�y����m��m���6�� Z쭭':���β�\��Dw�=yx�%[\�0Z�nf:�C&��D��˳��O���������	��+&T�{�ݵkm�ۛH;�Q�o��hh��Y��b�m�Y]A�ε�<ػ�7��ͷD�t�̉Wf�q,pг'k:�d�c���gs}�F#�	�Ft�}��r�j[��p�Y�9�[V�c��m��aE��ŭ��_s�3i]g)�DN���(�iT��c�B��G&>�����L�1>{Y|֣�����<��TW�R�'|���⹎�M��x�;�LggTG��T2#��[e�n^T��+h�ӧ����t;2���
��y�O�W$FT�aԕK��L�|y�\�|�'n���n�X)<"�I�*:��8A�ˬ=v�m=s��v�M�O��� ���W��.���G"[IM���@�MX�v��H�HoC[+�'�N�6%9��\Iz7��V�7�EW�Q���S����mC+��� h�Y��M�::X�*;Y��{��@͛��7 ����iH(�e(�4������iaV"������L�B���E��1������Kq�[Mf��L:_j��vv���sy��"����ꎅ;�"�7
Z�V������S�5�h���w:�e5
��@&mu���|�p�pR�n�ؑ�H��ff.q�6�W�8֙W\ȝp���ٮ�'�!���;5i�W9�7���0ŵ1��D����؇RzyC#����q�Rֻbt�WpOr�i�W��8rZ������J�dɇs�}������\�X/��N�gn�e�L)��df�e��Cj}��w��k��	ue%�^����,�Ъ��Z%h��Q��AD�,������
�3�S�i]o}��}��K�)� SV4ZV����u�v�K�g����x5��K:9!��-�O�<١V�[ڒ<�,��;x8�qH쎖�TN�q*��-end����\&^ۉ^f��ؗ�T�yh΅P��3%��$�s���}�7U�<Y�}�ڬԶ�^VV�ҦE�;���f4��9�9�ڈ�lu*jN�؏<� +��Be%C{�(f桁�x�L��{Է�ƃ��-�'Vc͡^D)��V�)�x��^@v�+��[k$vx�X��h�R�Z�Q6�;�=�mE!ݭ\0��hc3�V�͜U�[�l�ZA�;R���l43u�S�w<� �!;��k}�[Aؠ�C��_8��BAɜ����Ppr����:���jO:�j�Ӹ,KU�.K&�c�_,6�����{m��ne�(Ú�y<J=�R�%�i{L%��$&rAe��K��.6�
�j5�ѹ���AU���@թǊ�U�l4��Y3n	��vM�XL�n��U������H��Ӽ}X�f'�kh�-��7[�������6��@�ŰU����Tq=�y�VY��kf���B+4E��6#�h�P�نJ�S��Z�Yv8��P7lFmkŜ���ő�Ƶ���)C,"'t�1����_GA�Hy�1n]���8*f:.e\Q|�GKB�īw3E�ٝs��� ��F!�V�.�u��v�q�1Gž��׺e
�Rr���<�nH*3�"���g3vH���-�`9�������>ŷ�L��ii"ڒ.�6�:�K6RX����v� ��B��ih����&���vWN�P�d��6x�ST��Ӏ㦕����VEe��n��Z,M�R�|VhX��ӷY`5���jbɌ�x)6�8���OAw�j���u)������ă��ѷ�����$D���(�Ll��z��p�Rv�:Ԭ��id�UՂ�G��X�ֳ �ܕ�n�ʵ.5���>�N�k}s����φ*1�K���,�5�,�cM7i�bVh-�3t���;O���6L|�j>ʶ!�$EoqS'oW2�m+�Z��F�#qr�mK32a&��B6~�.�ᦦ�}P��9�L�O�W|��N�
�v���6�Ht�#3o��`�]Pq��:��AP{uM�:O�g'�Zr���Vk�oFD�O�5�T�7�e8ld�{�����}C ����,�il�m[��.T%�	=Y�^�Lޠ��[t@'+Yb�:�eĕt�/B��o��hn-����{"F�勯%���|ST�nu�㼬?bK`�C�YОݥ�-�qW&��B�B0�ʻwm�A)�Ȝ/�Փ��X�Mq�o<T3]]�`����f�Vk"L˶
e�.:�ZC�ejb�ub֩ZG/�Z��Y�����ka�eѹ��<A�����ZX��S�{�3Oqf%����ّ
���ӵ��^�Y�#3��	������1VM�NmJ���:�/�����g*�a�ګ2�4��ђ� ��ה�P�;Y=��j�{_G>S:-R��{��x8;9��ЪQ���J����2sݭ5�+�TΨ�ɔ�.�ל���ћ�k`���%�;�v�IgP�5�5BR��;���!�о�A��Ho{�r׀kk뚕KUa��`��i�K�޻����5�sz�*mX!^!�>q��RΦ,���������k��N�j��%,�� ���=͟��'v�K�3��I:u�y�e܂���`��H=%^�@_(�+H��Z�2�у�8h󏸼u�)@C�XF�E��Iշ��1��]xgv�};�\���fFFmZ�%u�B�����ƕ"�7gu[�ZG,��f�c�Km�wp���0����Nh�Oh��=DP�r��S���N0�s/p��1�#v����v������y%�+�$d���bY��c�LB�s
����\c�8��5˺�����W�fa8q�����"_b��hUb���tGIZ�o+����Y|�~C;IVW:���
��]��k���IJ�Ǒһr�p���]M�%�9�M��G�s�v�]2t#��z�����T�c��ٱ
�tJ{5�<�f��FYߙB�>h/E�1��c��������u:�5��t�>���鷐n��m%�DWp\��
Q10����w����Y}��ѴIa�L�QК�������wJ%�W"+[ή�-�;���o*��nP���4�R8��T�ԩ�&H�TEI3�{2�jT��$ɤM���Ȣ���L�#�;�RM�u�$�$����rI$��$�I$�I�I$�I#�rRG.N����'s�I$��$�"rMrC�H`�_HeJ)Y%n`9۠����2�zl�]�3��r��C�+����8naI��Mn(�o�#a��q���4M�
$%_b�w����_c�/O*�&�+���s�c�m�n���w=��� ""�����"
���~�Ϫ���?">�����������>}����}�����M~�T�+�i�Υ$9Y�B�ެ��
ط��õ|������ۀ�9+�y�w9fsl�;RMZU��nv
��"Ю��B��)���Z��޾�L�L�C;-���q���(���_Y�7���q�D76�S�5i��c۬�tgv��MN���5���f�T�t� �ۛ�N��Ǡ����V5Օ�r98�ڬ{>�@�,-,�njCN���F$*�C�Mqp'��$�+��%�)n�ǫ	�8Jx�:�3o�YC0�Y�ă�����1�oYG,𛃌���tN�J�dJd����G�]il,ru�r��n�܁d�`M��+3Ews�9Q�iS�ΛiVg�q�을�w��vX\���@蒳��y�c��":�u-Y�7U�L���R^_H�W!�K�P�+so�u��5�9��c
`ض��C�m���=ZA�ƶ���*_t�!O[O9U�7��w�(Pw���ڳ�ڢ���J�`��T� ;غL4.�cz��s�j���f�x�Xtp�Z6�>���&.�62Z�֣��`�V+��^s�(\J�����U��TwU�����e0H�A��las��a�i_*��#ȃ���-h�s���
�'�8�2o��XS#�$]�7�D���N�r�{�]�I���]�n�t3:��h��w��!��`��>a.
�S�b��5µ�TT�S�0�ۓ@ᐹ�tk�p���G21�ۧ��3Z$�t��Zj����ɸ۝xԮ�%$i�f�sM�o�
d�t��q�EK(��"v���÷�͵4��T���4��b�V�\o�]�]��C�λX�<xn8�@��r����
�ڟu����n���\�������{�&Q��ۜ�	y�sn�ǁ[U!��mS��{p�ת�K癒��*}�m��*;Ӥ!��N�34pxI�nK}��\�a�݀VU�	�ou{s�r����d��e[aR �I뻘�I�}3D�(�mu���*�y��w���.��VYH��h��f2�]̓�9Ϯ��5v[Et��m�0]e`}SF�CY�=��/O+v��� C�d�{��똣�]8�ӝ3/hp'+kaK��Xef�1�]k"d>.]��>���L"M)o{�0m拠t%�2��X��k�/&j�hV�W��L����9�n��IHLˡ�����uę�w��n/5_pA�GWM�d5��LfZ�ʇ'��{]�,���c����鹡��F P�30�����+|*��D�	��0���-�.Q/^����nh��{�Z͸�Q(���g�&��ճ F��lv�8������:�ܯg"tX��uj,��n����Gt6���:�NT�\[WN�M9��nf�X;Vȥ����c]��l��x���I���,e�r㤤��an\4ˏ��y.ښ�`�%��"�����|����0u��y�JV@(v[邶m���p�b�Z��]�Y;w��4�I��7��F'Z[��]��)ǫKs6���/���ct�p$Sqm�j����s�8��m,��ƚ��:��䕗E�q�2�+7��+s+:�v�7C1.Tfc��Z�����ᗎbX�*;8QƬ�3I'��ݕ72�nF.��[��å�l��B�}v�bO,�f�Ȼ�M��t>{[���+�*�A5�61s�,P;z^A#�����آn��/�[��E�Aؽ�q�y�_w��=��u�ȋp��U+c&��k6�d���f�&�%��$���+�Ϋ�_J�F�9�92 ȯ�%+& 4�mY�6�᱃)�k)�!��G��jKZ�NmXB�X�IJ��I
l�>�:���T���Ao.\�]i_af�ueeK"�I6��6�,�Y�MZ�f��(Q{H׀���.�v�m�7d���㧅���wY@eFɲuc��� ��u���M�a�b�-�MY�awċv��n�)�ڨY��S�����|�%b��v5!4�����GI�R�r]��o^�F�]k1�L]�7�U��$�8t�/**�a�b�ene���qJyK��ji�b�I]�SXj�
���r\���}B�������la/�h.����/#�N`�/��ǙZn�;���(�OH�rp�5s����F��,o�
-�N��>�DJ��`pN���8�k]d�+U��Kv.H���,Oc�2���S���x�F��^JY{���U,�(tU��52�{H�Z�e"�
�#(��k�j�P#�qy-�xMu��u ފX�c�J�8�����}��.X���1�N�x[���Oj����[�0�a�ّ��p,�Y�{�mɿ�)�I%�v���o痮��Mm�y4�6$L��cl^�,U�ޤ(A��V��F�B�AeY�Y�u���N�8 1���tC�õ��<ƣ���!�\o���n�շ-��l*���ZV1�͔/���*hmKS.J���t�$�l��eK��� _P�k��Q�35;�+P�ӛ� �Ż���$f��:���n�I�7Uu7u4]�3$Ŏ�z����ڎ���<�_nNWٔnV�/�E�%�{̛Q��G��e�����Cx�Z�qΤQ��z⇪��e�&�h��.�-uJ�-��.w$��5��A���Wo2��֤�R�m�\��{z˛H��9�ycp�O���5=��aYh:�7^J���]�%o_fޑs2]��h�(*�٥YB �2��]���qR9\����P�3x���X�mTܮ�y�������ӄDIeY�K�YB�l7���;�9�1$༺"'����K5Jt���`��3�\�7:f��ޣbm]Z7S�[���f��ۙW/�m�@�w`����OVq�Κ�
7k�<5��D^V'7��*wop�ٲyr<L�4+[Si6���ܨ�-���|Xk�
��e�ki�e^+���1N�RI�Y���"E�*�GI���y}园�g�˙���]
V�����j��f�d�+��(⒔h��8�����i��m��o�,żw(����;w5h��K��j���T ��r΂���V*��,�+] ��E�uԂ�.V���ۤ����픝\�m1��f�<���'VڭY��\���\!ѳ��z��i���x���EF�[-�9��i�}u��_D�R��-��*�Z��]���c(_n��}s&���.u��L
��zM])�.���O�܄Sn�E]�R�쓘$e[�x-To��	\w쥓�eo������zus��㸹���l2���`p��r�*8�g�8S�vs�i`�������rŃ6%�e�p���o���$��o��7�����a�n���oj����%�7�.Ң �@	�,{%1��3fc�\��nu&4����3��Zřz3��ፓ����:!ک|��wy�T�i��`�g��#W^j�]���KA���j\u"�u��tD5e�5��B�T���yn�ގ=]�#�A4���-��R�g3rM�!��F��:�1��Ur[�P�2��W�����5�p�kk��;�m��Sݮu��K�u&��n��1��opr^uh�qjÛ4�";� dD&�R[G^ڝd��N�FV�xBBE[m�v��������4�����w��P�Q�ݩ���)T�h����gj��J�;�A3����N��:�h}6�f9�d�W����:OpF�WQ9!n��U�@�+̫�:QI\.w^��4�w�\�	ڹR��aSt�gN�$�ǹbD��J+���{��b�3N��7����)f�3b����;��N:[����y�)�^C&P͌�k�Yu��oMq{u�>WN�Lg��W�f�kDS�䬂p��5���Rj��*�r�'5,�ZXq�F�B�ш��s���e�3Y��m`K��sz'Zq&Nh�]l�(k=,�q���ɵI5�Ō�\S�CZ�T9�[��KR�1�<a��!�1w=��p
Z���!wVt������af�],��A��;��sm��(�elu+1���oz�zq*u�-�4�w��L;i��es-E՛Og V�vо*. *wT�<E�l;�&Ѯ���a#l�`nȗQ�ړutۡX9��lv0]��J��ZD�R�D�G��ۑX�@ΒZ�}�PIl�9Vd���wuH���׉��I��k��^��_VI��C��t�
E,�ÏB
�uKWG{:H˃R�0������܈+rC�+8N/&�3�`�U٢��f��eͨr\�ܢ&ݝ�3��%��4�QR�VRy��2g贾H劳4f^2�oE�T���q�_.�6h:��=�Jo �d�i?����sr=��숈G�+���LSܺę��[)R���e��%�v����+S��3m�|�nq/d��q�Z�s{��{�pYIu:f��2%��X!����J��Ҧ�=]z�fG��#� ���&mA�ju�ɝʴ����]���i���-����^⨰���ͼT�Kf�
���>2�����,�۝\�+|e-��r��g�rf�vܷ7^�5(���{���4�8jn�<���;/m�k���Գ�!���;��������H�21��.9wM���Z��Qt4^>�L�mC���-|��jm��Nç�˗ØѸ�G\汙 ȔIZB��}#�z��C�Ei[�|�E���z��m;��b�.�����f<�`9��)��DB�;wo3��A"��S�m@V��7�!YF4n�/	p�L�����ݼ��������z�N�3E���ZY��֥k�Kk�Z�R�V��@.�Z�;1`}gV�j��i�kX��ϕIÙfa�0@,Q|k���"!�03k ���qDF�V��3�zZ-��Vhմ�D��h�����X��9��Jo9A]L+���[������d�v�L��
����9���eH�)*�p�F��Y%�G�r��nQp��x��B����H^Rů�(w'JT��4�U���Ң�ĩ�<E�;�z5ə��,�&�4l:�����:�Jn�;�2�`Ԅm����f�u��s뙁nE�J���t�L����t�$�W��٥��_M�����Pk�x���a��}}�7��S��SGA�k�]��剈< u-ܷ�å��8�����0�..j�K�5Z�'#�}9�6�_d-q
��h3ClکIN��p�ck/:��@��YWSH����@�V�aS��N�غ�3eK���:�u&*RܶQ�����ٕ�h���*K�nr�̗ь��5���Y����]k4���)��;�kN�ރ{�`����oC׼Ms|�+/����+����Wik�r����J�9�q���A�x^>;��ղUl �
�
g ��1�GV�}ۋ0u+ԡb���Zd�2ޥFdn>�W�hN����r�����T������٘s��i���*Yw]w��q��p��p��U]Zȑz�`.�8�j�X��ଡ଼��D�;м�cK�ԅ��&��rh͂����+���� f�rmл���Y�4zL��y\;�Eu,��렞8�n����X�^r�r�n�	"�ml�Ƥg��\�\v��6w`f�l�	��@�յ��:� ���04����>q�V��U���N���1(�FP�{C�pں�ΕP�h��n�q]�ݧ$��#��Tub�J�]�u�Z��G_o\-�:�Vӆ(\j��w��t	:��=�iU����imb�X�EX�s�m�O
Ab������!�[N�W��˦��6%b�Ves�kDqnMuX� ʫ���̙��+�!댠��U�쏒�q�{�H{�)��6豝$�fQڽP�#��#!�3s�drfΈr��`G��m�5M��˟S�z��\|&1�T��v��=�GO��pJ]9���3[5JB��(n���$��iҭ��}�Z�d�
9xj�v���7�n8���1�ΒkÀrٔ�o�=E���ظ �E��m*�Τ�����)Oݒ�x���s�G��:���!S�/#�jH;��ȹK02���e�ט̨巛M���0�V^�\���p�gl�r*�Ք��w�����Gpl>��WPjC�YKs��H�j����Eӳǈpe�V1�ga+�B1Ӣ�ec�Â���R ��Z X�_طA�}ҭt��vk�#��-�/C��`�}�5SL��ܣ<s�̹ƟM��ż珵�,܊K�t�<ܡ�J�:9�a�C�Im�Mp�t��،�.e��r9��d���k X�v��J5���uFВ�v[��f<�uɘl�i�n�� �K�n�:�q����v�I�ؓZ��L�Չ�8:����z�6��:���5�HоۏDf�ǋ$��I:�T�>8��sw�^l�-�7�i빲�yr�yA�m�t���c��VH���X��4/�v���{W��D*�v���:�>���a6�O��o�e��y	��W�F<r�7$����u�V!�*��5�k|Ѳ.��[�SI�q)�4���J�ci�~�QFY��R�����X��x��6S.nꮎ�� �oV+�E(���3������ڭ���u�}�G�f�idi�P�YU�4�R��k�9+2��ӊX�AN\��z�1�u�=q�J��,1 |���R{mv[�Ux�Hi�]N��w:�n�A�O��b�ӭ�1.�F �.IWE��6(J�W�n�kݬ�����}�m�,U��>�gg �F�����}os]K�����1�}�]�����Y["��Wk�1R�.�A��Bi�����)�V!��%��5��>�H��c��!K�r�v)V�-+R�o9yvr6w]�EZ��#�*k�gXy-�9����ҷ"7,bz��4��-FG`	�|�*��.�sW�K��z9�!�ύ����#W�îz���oC����)5������?�=��x{��@����������~����}��x���>��? ���h����9'��nT���-�^JL�kKUo�d6��K���u��jbM�	��[hPY��36N��.Y��Y���~���C&���u�nJI�º.U�ܼ�)�|�K	���w}�Ǐ*⎙�
���;��ڡ��಑5��;�
�@֘��2rp���V�fd�t�k����E���]���s���F�F �9f��J�B��;RkqVcf� ��*������	�_Y�j���]
Π7�RbKj�v�%��T����;��u;��Z�,�rK���.����H�P��JK���y.������uz�6e��U#��o�[�S�`x���{�j�7�j}���]w[�ìvʖ	�;M�5ǖ�] ���tQ���؄�F9��_	Y75��s��XclӔ�uh����-�M�/z��;#�Oaӡ�3Y��${$�~���q/��|�����G�6�c�wt��o�����o^'��d*TX�QԻ�TV��������s�� ���e-6�������֬5���
o9�S��L�� ��9��R� �F�����`�v�=E�Eh�6��5����hLZ{���������V���mq��|�$zk����^��%�V'eM	��I�Wi�ނ,W�N	������Ύ�r�G���{��i�|�,ܮ'D{%RY�«�a�#6�JR�$�I3��E�{�f��A*4x�C��*�ݏ-��Wy�?J����QMDQZw[�88jO�ϛQ1mZ���kY�����Z1E�*h����Vڊ�(��h���v�WG�l[A>A��j���EE�(�=گ1�m���3%ETEV�����Eth��OZ)"�o8�Cևo8�v��7����ᦚv�DIU�G�SGNjb�m��UEEQM�4MISW�b�(���+݊���LEf&������RE$LLh��Um����\yb�*�ֈ�';&�Ѷ4A;j65D41V��Q1[j�iذj���#��8��X�j���&�cF���UE�MS����D�DAIA��c�Ay�j/,�PZv�m:i������5If�m2SUETZ1PA44PhuLTkTQ��ti�l��CtTFؠ}ت��.�4j��f6U5ZUUF�Q�ZM2Qh�y�TLMl���PC��*�d���i1ݒ���:,pw�|"��WT��o2> ��CV��c]M����2�U�D��媎el����	��n�|x����7V�t�J�ܻ�X󊓋�P����"��n#sO����Q�zyR�ye��U�i�z��rs�V#k.��{ޱ���2�b�i`�V���n�;�H�S�g��^�	��E$��V{�x�]�Y��Ufe�/��+66��P�D+�8YƽԒ�f�CL�>[ї7�kU�m�6���ކ��7�!�R�+�{��̨zVx���cxS�rS��~k�G��X�ָ��f�$��Bkuq��J�{��ma�3���?5,�w�o���zB�-�]5|��b���ג���xO�#�4�W�������%�]Ʃwp���M�Vb��|bV;�|�1>ឮ2�?�@a��D-�=��ڏ^^����}!�vӶ����l�K���cb�j���4$yV���єy}�Ī�pg^��!Sm:�]����&\z���YݼZ�&yt�M�z/D�5p�7N��my���9�*�۳'U�WLT���"�^vgt��sA��%�L��֨,��>�7\�J3��7�"��T��9����;�����8�r��i*c"fR�w2����m#Oj�T�R�W�WaJu3^��Vi���yŝt��~�w���=�Q��|��Y�� �Šg�;4��Wo$i. ��d0F�4�V�B��������{l��e�\��D�RFZ�=G�������G9L}�u��̦�Xg{������վ?<Ѕ�׹8�v�Д�L���ow{2��}Y~)a�
�-6=g�yM�fOf�^<��<�Y~u��V��|�W����₼J��\(iFm*���������7��N�m�JC{}�:��P'T�%}��=�k&YJtO�[��S����h맷���'� �XDm�%c8��B��"xg[�����U�nuA�������տQ,�V�5���ի�L,z�3d�/
��肇����O�}5�u��R)}~U=����e�rW��jיCǽ��b��;6����^�מr��s���i������Y��:��}�b~�V%Βr�h��u�s5��O�_!�@T�r�(��45l�G�5���8�&_f0[��hüoeڑ}���[E%{��|���2s{����Q'�D�3B�U�N5�y�����N����~�I��^�D�` �Ч�{ԯ�{�t��U�+�6�b]�m��{����@x���V��e^)�)�T�YYsk=T���r����W�,��2/�Mݥ�5q��qXj��7'�>�__S\0���>�^0[����N��}�+�]
�ݞ��u�ﭷ�N2���5�ռ]*v%zgbP)bf��[PV_�9\�~_o���!EGjQ��N��!���fB6�%N�C�b��3�*�W�o�x����Ӽ�X��
�󼨫cM�O���#F{�=S���7D%�H����}ʷڅ_$AX����t&�W�J�����9�8�7?hUA���t����m�$��L��ٗ�h�<�C�U��@�MU��p�2�P�E(��d:z���N�6��
ح����a6��e�d�FQV�7Z�ZҞ�����"T!_�C�9�l����4��TP_vZ�����j�MJ[�-�u$={�D���c�R�=��1��~}��<aB��䠱�����V���MFl��m�Uέ�B�F��vF\�5mr����cv��{6��M���-�W`��KwS�����&���iޡ%虾$-�IJ�+7`.;���
��E��ƻlǲko�h��9��N��~g�),3H�K}H����nJ�;뫹'Է����--��| P��:{c�u�_{����R��a.&���)q�U=��]��)��K�
#F
s�n7'F�Z�V�S_����쨺E�H����6������>e��;yuҼ��)���߫'�<L�~�4i��F?Iw�w<���Hk� k�6�8`���m��E�ף&٭
Z�+Rc���~y;w���7��Y7i�A})3t�2M�_����3��?N�����J,
�v| �� �s"l.��4ԽJ�j*a_��ǗB �>�X�C�"�u��4����s�]zw��T��k����Pg[yT4��U�~�aHeѤU0fۓ�bg;�):Q�x�]��}��k���v��; ��6�>-y֡�u�<P���Wv�h}:N��L#^(�Y�y�`q۔�>�sl��2-;�EwZ�cv��xVVt�}BtP	|uZ�Y����{-\�w2N�'^a�b��47ۖ�ŀ���^���,����hX�0�M�
�+ln��l�uKu�r�z�,��W���v�l�Ԍ�1�k-b���2�mD��]�;ʝ[��Du�*��NT�߽m̛��kٝy�j�U��ED��@�¬AXKP�Ȋ�W�VJ��H��+:4�T1oWnG5�RXY~ŜT���^��q�U=�{p�Q�����x{�%��Q�
Z�Q6��J}<9�rJ��me.��e����%��EN�cẸ�1�����RB󈯻WX�A,i,I#q'U��֔[�sEu�9�V�>NW].��\~���Z�V�������/�q߼S�����b�ܬ�
ͤU��b3%X��7%.��A�"�e@�]�}�^X��EwQ�s-����[>5��2��/�>�z�Q���1w�����G������YP��E�q�߶
ꁅ^�/,R�:Rb�	r?@M���X�,ޜ]\��|�;wsU����ś;ܜV��ֽq��}$�,h��8<��r��4�̮�*���	��4n
#�t���e����O�4�j���]��YH
� ��_k7S;�G����uӂ�ܭg��."�C�#X�w �7�c��P$w���ڣ-r6��)ס��z���W�|O��N��Nݓ����G͚�k3n���»�s�ra���C��e����:���ob��������h�������@r1�g2��L��Z�/0�lt^0["�*�*�����<�dî]5�s7h(P��Q���3j�J��K*���)G��)*XLi^������b���u�GR�;���EF�q�5��]8g�V��G�ȋ��G��=�N2B�����$,P�S��V�g]b�ˆ�'��m�k�J���jA���q*v�^�kC��������ET��I�.��$��j���н�|��7�>���R����M�v	�n�/@�1V���0�DT��[����D���$>�ҍz�€@����69L�F#�#�O�*���IoW��]:C�	rZ�H�3�T",�W�\x]��r͙4q47.)�lu�������(��V��\1B�tI��6�D&��<������YnX܉kL`�o5��d���t�u��7�,�ϤŇX�q���U�^b�v��ܫ���!����Hoo��3��-�b�X8��ɴ����m��mrH�?++#�4vB�y(�#n)/F���C4���
R��T�Ux,���#��Մ�̟o_ѹ*�@�FP��oF,9�3�qβvpvV�!���֒��Elu����#c�=���������Լk�U��(�g�oO\�:�勖�!y��m.圪�Vj$q$���ʺ�g�^w)�<�c�-�Jr��h�^3#�MB����G���������9�t�
���Y52n�pGL�!����x�o����ӕW��������~�.����j����^�8��ޕ���P���{��B�]G�j�}�Z�r�7Y6�������]$��Z�ݨ�pґ̔qh*�%F�F�i0&�����Q��{(���~�U앒��_R�*}0�]�cZ�\ϊ�+.��;��9sY�E]0�����6j}2�aQ�$� �Wzۛ��|�	��+�5���j�x�\�l�w��d�6(2�'�G:��"���6�Z�RrM�F��0��v��X�S��6�GRe�Ɩ���o�����9��T��Q[�.�\�g��s����nh^����(!��^��à{�o�
��~�#o��e���s�e^W{�=�t��'S�+E;L�/DL\�OP5n�;W�*��wzVj:�_{FY�	�c}��!R2�(jt�N��<-�Ms�5:9N�^(���z12�K�ʊ/W�{��ǽ�D7WޯnV�O*<�*^RE����#M`_w��=��K5+J�yvoU�Ĳ��pU{t-g�:���p`)����X��,zOCp����;��t-�V}���פ��c|���vJϩd��E�5���Ze��D{bi]/d]y]� �ȣY�'H۟�#k�!u��t����S_����Ot�t6����:���y0�e��0��W��M��>�]��}�0�.���Gɪ �΁Q�TT%�U��$�z�omu��!��]ܳ9�e�Q��9,7XT�^.{Ob�:yӹ�+wK���#"B����c/7AS��������6��]]����Ш�\n6Y�8R!b�Ŋ���� t��tr�\�Ҥ�Kż��2�RY��U�H~�A��A�YWI�מ|<�6���-��l���r�f��k�i_I�~�7�߽�&�b�(�|:�T��ț~�ߥy1���e|$i6��oX�od] �p�D��`��{D������~�A>[���W�?#PR<�*zu~g�T��g�h�n5Y6�s�
���$;��C��^�b��.��@��V�YY�3cC��;:'��kŶ_K:�N_P��m��ю�TÇݫ5zu7Vvz�3�J�dpp��Y��=Vw/�q!��N�WՒlxF�T�s���Jv��
Լ/�X���n�r����gPV�,r"�{�d�Z��]�3�6j���:�_�
��bz�:��X���{�j/W�ۑ}=������:b�]����{4n �2���D,�%����-Ϲ%b6��]�ލ�S��=��j�J�^��Gu��*U��ƼR�-���MZ�z,��ph[�C�ڧ-i9��t�Q��cm�g��;Y�y
ҕ 2M��@]mWN�@�)�l�&��ga�Z7�R�cv�Ω.��� �q�]��`�B�iV������̂���Mr:;�����=��6�RB�ں�J	���Y�;��'g���&��qK�;ו:���W��uԬ�@�Wk�o�t�G�ޗ{�{��'��a���U�f�G�T�۷B�BٳRP�m�љ���=(핀r�V��W���8l�����hU�aJ�'A�&��d�8���WY/��T]����b�H����Z�z=`r�F���}�*�����h��,���'
���þnf�7�.�]&<N`~����}I�^�}��Qe�'dڀ��ߧ���s�f�^��w�d��_��e�����:%4$yl�n���PR���јp�[�&���w�Щ��׉��"8�G ڿx�a��QghI���l��}��1�q�>lt��-0�+/�X!��
#�;%tgU(����b{��Jǆ<��J�$�;gJT���ﻭ�Υ
F�#�&���%�e�e�b��-�\XI]N�Z�3�cB���Ε��V�[}���fh��t�.��Z���|]�Kj=����p�]���]vdX`P�턆�ő�V�>�1с݇��R�E�ۦ��Va��}[�2$���XX���q���oYs%�Si�@=v�Z�	��${�uͷñ���,�).��bK:��6]k�oM_!�7�(�f�U�Q�okMbI���.�Z�Wc�C]�kaےr�:��cƂ�hdZS�F�+��
^e�f�%�$΂��r[}z�����_���Cw�����qe��w��3��f>��0.�P��i
b��.�Zɧ���A�T����5^�xsl�x����ƌZW-��2.�q��M>��Ke�����(D=��Yk�R�j�Q�1�-��`Ӓ�7��U����Ʌ��E]zT�\�DeF4����!qAW��Vѐ�09�Ө�u�K�u �t�n��dC[z��J����3Qt�Xr�mU�@�$օ�Hm��z�7���|XvT�s*m�A��]b�+m7)��&��V�

렺�3lҋ��>���po_H��@�a�1���qѡCu��KXi��`�ӴCCN�{D�e�+4�-��[�w��3�Y�N�����H�a�ۮ��wS���;�8��܍vC���s#�ɕ/k�Y���ϣ�T��9�)M�}�d��>� �˫���3���J:R��8�l����B�uZ��!J������r��"�:�4�n�Կ�vS�ޓ�����W�{){r׋��m7{��%�LB
}�r��B˙jW:�XL;)�`uva�.��&gv��ǩ���O�U�s3�p�AF��֔��̶3)p�G@6�k�l�o/v��.n�!;t�ѡ�N�Ƀ����4�vW#2�]�P� ��h���/��U�[�,��+c�:��AYZ��C���N�uN����.�VlQ�ԟ,QV�a�U��5�ڄnգ���s!
J��Cf�ͺkD����hm�h�b˃DKj<�%ޫ�|q�i�ǲU�B+�P\�������G:�^w^r�8�U7�}��	I٠��΂
U+0��Z����-<��R�XƱL��7�]g؄���ی�n�N8��u�����Z�lp�!�]Y�]-l���#y��Y�#�|�\�׎i��u���c���R8�О�4�}Σ궑]�yR�g1�\U���me�$ �*����6�@P+��$��z	�s}mn��/&d4��J� ������m�3�v�{�S����B^�1�г�v��:�������ͽ��$��.�,�����+�j�j�r5.N!.5|.��FU+�J
I&I$�3�>��>�_�>�qvl`�*&�֐���v�:�AIL��4�Q�EM]�AARSu�=��DL�U1LQM^Z*�.-���uQ��I1=�S%D��	@LD��%�sj1U嫶Jf&�jb&��$�"�
/w]T17��M4�Y�H����+�Ӌ`�U%SV�Km������U���f")�(�M=�$��bb�*�-`��QQGF;���TQ���SLTF����ڍd�&"��(4b
��٧mS�V�1�55M�P��F����Ɔ&h�d��b(���S���LVê��"��d�A�*� �Z���*��/6���ګX(�i�h���������
����-�Z��b�j��ƨ"��1P�L�[gX���d�� �*))�Ͱm�UTK�D�B��`����;Ϧ���������W�Lž�IJʍ-,��B۴j��aH��g(�{[���.XYR��v�$��/Y)�	��d{磌�P_"V����z���j�e?|�^��s���F�8���-lQ�w�9>Orwt@I�^�HׁXΤ�A�l=
�2�`�ߎV���8��q��z� �7�av�D�׮_$��,w�ٵ۝��:�Eۤ�A�CG}h�ʅGzDǭI]w���Ȏк؇�����~v�$��N<w��&���Ze��>�J)���0�G�)�Gaܢ�
������=W�I���yk^6/�?j�~K�jn]�<kѹ	��q�3�3E��O!R9Hh���-�R��h{\xxe�Ԥ�_��9TA�T�7$6�!׺vy��w�)�a���M�5��@w�,Ȧ�=��:��N�+�[i�Y��w��`��U�9&��sભ��v2�6��������ծ'�{{a�[�	>�9�Q��6qZ�� >��E�N<nT͹M����3��j��py^�sң�0Qer�9���+�P�b���
1��dA�S�|�Lb�p�r�#<�2#l=-�����X)����W��w�\
&��Ӱ�zJE���fw���AgM�i�/� ��}su.�iw���tt9�OR���k&S<���.߰\CoG�]��h���e�^!��.�q�r�\<3y`̸Eq^�=jB+3����Z6�b6��^�)�v8�@�kF�e<N�Sv�p��Si)Y֜��K��=�b�]�l�	�z(�spY���.�B���@�R�:(�Jl�k�,���8c��0Ö�`�.���fO`gw*�H����"䟸{���q�W}���^���[sP���)z��h�>��]�`����C�8���8����j�.�����R5��ڬ0������=0 �
1��k`�:J��|Q���F�ͪ���m�vi�[��[r�� 4��:�������dIM����]p��P�-�d�'�yi��t��t�W67��g���a;�-;�[�s�0�t����a=�!ު�:�|xa�.��	~;=��D��O?8���GW���)WK4^���+Sc.�_��gA�ǈ��F,C��X��i�g��n �q���A���7Q��o��}s��.�Fi��q�K]S|��!��D8oil�įu�z�Ĺ1s9�PH�nR2îLTW���>�@�iSY�C7X�?��z9J}.����.f7&��9�!��qW�\�:�.�wy9)i����+� ��"�^�b��i�b�AU�^����(�#Gڗv��u��mAظg���/���j>Ke.&�ɱ�T�LVM�¬�`oM�Q�p�eJ��Ttn��7hr=�����3`�=���+�O:{|e�W&��8��U�m:u���Ԕn�f��)����k%�j��FΫ��^�kNqS��Ȭދz���d��Z���b�̫��GY�� #�+��9��U9xpu�N�
�ܭM��Nӑ���qf�5A�X��e��̶`=�ا�ߣ갅z&4�B}���*�<8�Ϝ5&���%�{����U�L�cr_�m`r�t߼J�� XN�Ms��d8Ѧָ�k��-B�^b�Ae_�	��F��cn�l����*_��@Ň�lvo�U�,7���l�>�y�I�9��s�'V�]�QR{�Y�0?[3q�)���P��+�8���=S�H��`@��r��^:���5��?�Tx���'E�`աU�Hԝ�Y���tS�'�>�D�1��4�V�����n��4�7Pt��,��X5�uo��6��O�>�}n���h��Ӷ���л�s����;@��p��ĝq�e�l\Ǚ���8������G�Li$uV��\$����a�q�����Y��������~aE���.a���^Al��w�D�r��>��+w�uOkܘm\���m����z}\���ЏR�ԕ7���U��E�i%uF��GEM%��9�m��,e��kxO�7"/����/�tc*��F��"U�C�e��l{����P���l��0�#� ڶ���_4N���ͽ�z�k=պ �������ɻqֹ�sX\�#:�+H�чE��יB3%+�UK����Z�;-�&��h��E��^�����,�<��j���|������Gz-{�����ei���t纛p�,9!�XcY�X���Գ7��=��^l{�Ga� <T���f�=�f5��\z9:�WS�k�[�x�D���0��%Z�fc��s�1����&��?i��C�i����.a�-Ǵ�o�mOk�?쾈�Ȯ	k�{�<�v�d�LPA�Ň"Пg�t��>t`�ͫuXY��d�+v�%ԍ,}a����*��#mt_��(�9s�
��n�pi�?{�W�#Q��Ga0z�^SWK��M�q"�kL�U�lgC0�fP�0�,����q��U$�wD4���E�b��}X���3�;O&ǖ�]�[4��X2,Y*L���A��z�A��:�N9����[��9������Z�ƷJv�Lc�r&+l�v�����bNC=��p���[K�{n�x����L5��uH�ލ���s�������WmT�J�)߭8�1~�^��kvHf��SG����xR���
���16��<�gq̫��jl�*^r��,[���V38Q؝��ՉZ)����*sC�$��q����9�E(V�}E��i�aW,���w�J�2�cux�����#�2������0� "I߻/#��8�a���zm���\�6�C��5�Wz��Mt���Vc��[U�"~ �LQS,�y���ёW�M��I��g뷆dN{�G����O>Μ�'v���V�-�5�1������C͛�=t�4>>��W�6d�yFO>��ZRv}hN���Y��²a�S
�5s4Ĩ^�Tr\kj�ζ����t��p���u�?�B�vz�.[Cb�����x@���n���~9/a�iA�bpOEC����]l&�:q��0q��/[���qv�D��1�]:gV��6������Oxi�.�f�<��8k�G�T{e>�w>�8��c&�#�u��O���)A:���V=�i��ܻ�� +��Q�/Ӑ$�@�gi�(Q��Q�l;���϶F��,y��81��WFa�ز/p?G0�����9�lߠg�׽9��4��D�p�r����j���>+qs羖Dn�1\qDA��U\7:;�%��vy���i�tǌ�(�����'�x�K����68�q�ֹu옅	{��xw<yb�W����4���Y�Y[AQc��mk��SC�?�R��&�g���͖S�X�����$��,5B��fT�ϰ�돓��_Jr�靼lj���������Cv�M1���TS���4]��3	�ז#²;a~=�I~8��6�5�6'��F�T�=;W�2��O}�������F��E\B��"}�q���E�q�s઱�`и�����~y����Q$�}�Fb^�&������J�vYpxߣ��N�/U858]k��o�j�j�o��e_�'m�9��a�E��^@�Fě�^��@tb�P2:�����^A���U�ӵ���2�c^#n�_S�lsõ���%6O����1�p$��SJØ0�Uٹ�(V���w�.`�6g67K��F��[7�=Y�� 5�\$�(~�²�Q�41�Ŗ�S�?uEO���Pd��^�v����u#gR�?G):'�8*`٨d��b#�w61��<{�N��/z_���9�5*N|<�
9��A���gɼ�Hわ4�`�0�CK�!e�b���H� �A�?�s�B����ѐ1��pA�^9�Н����89��Ԩq�+���J�;=��:�0zF}�$���ع���h�����~�����{�������*r��,Meҁ!%:n���d�wH�!�*�c�w�n�\�W%d���4���4s�u��Ef�7lh��X����氌zo]E�Q�����a`4�9\��rS���n^�}�wlܧn�����<��a�$��f��s�ڭ;ͫ�<:��E��JF�|D�1��ݻ\osx������1�7�B1�s	��b�싁$�C\D{��i�K���`{�D�PR�<
Q'y�4�#��ni�44�l&2�)�BqLx�%�(k�  �Ż�;[�2hmR3�s���N��XZ�g�8�z7��Ü�Hy��=Ǚ�"��~�@g�$�[���7�.�׮=���5�R�lea��}}2�L�T�?N�X���x1��P21��D/oٶ���I����:�]bK��M+���.��Ϸ� ��n�ʙ�%��i��Wtj�m��qe^H�)ߠY�lS�~��XB�]6$�!ꨂ#��s�x���Z�!����?fZw"�<)�pn�:dv�����-3�Ua�	���Mtq�Ɂ�L��!�$�b���_���L��\a.�z�5�'~�)~]��f�`F���1'H�C�� ��M����M��'MG#˟0/���,P3�����m��څ����$q�͖M� �f�Ը�mT��1uNIP{�LU���ە�װjЪפjN5���n��T��T��}v�^����W���[�vݭ��kW�f�a��d������f��ǲ��Œ$��/�87b��S�y�������v�j=�Yoǅ�QZ�'05R���+�vS,v��vn�sڮr|��J�K�q��:���]\3�d�lPjcp
Qœ��'ps�U����-���D�#����.HRa��c�X5�} �i���)��t���}�yr{ӆ��e�<������	�C��f�gC��Vˈ}�x�c<����zUl�O�ˣ;�x9��4A�1|�u���T`��6�����S�Z8�a����;S��*+�0Y�	ɳ�6C�9��;-��ވv���p�c�Y�xi"í)��
��?Ǐ[�������c���V�4/		ϛ�DX,�Ņ�[>5{5:�D�*�Lx5���yU�r����
簩�����;e+~�a�S����W�d�%�@�ʗ�����g;/1p��|�&���"wv�1�f5W]FG���>���<{b�OH�(v�A؟��LfU~P? n����Ț����_�;(b��7��u��L[�h�pǹ@���c"w�D_Z��`�"��3E� �LY��^� �#A������S�F1ʢ���0��>�
y��]��"G&\4�a���9�o@����T_�QD�9Gp*|��G?l��s��>m���^H�ܭx��V��5 (w�L:�?F���i����Bѱ��뜭\h�9�����մ>IW4�n< �J1U����2�c���32FJ��ڽ��e�!=��ʈ��ڕ���[*|��t�[��6��.�+r�+v�^�$fEMݗ ���_P�:rU�8?x����9~SWK��YX�`���Cv��6����}+����������`�� ��h�#T���ǘW��;O&ǖ�]�['_d�����:��z�Q�ۯ�h}���HS��,(X<���cb�n��79��ɍ�P�ҙ�<��W�`�u+����\<p��X�_:���'��չtk`@P�#t$�\��Q2�=��ʌ�A�%��X��xu1y,yP�&2lEh=BE1F�
���K�8;/#��gl=v��/hL�b�ֳ�*�g��Ze���ntj�?eD
��
��pA�6�3eƏ]Dw��z$��TC*���R�2��Y�����N��IN����*�	H��Bp�~�iv���y��-BL2�%]�]���*aĨ@,����;�}������.����W�������a ?�	��f�����ұ	{����8�YɅ8m|}�58�����VR�-O��u<1p,=�4=N,e��s��oN�q����"/��=�G8b�S)hN�nb�w��m�����n��(��$?�]Mx�����y�NɘklTB�ꔯ;�g�ʞ�p��|��թ���6��һ��#�Z���\����vb���>xU]i;�d=��b�yM�Ҝ�bt:b�H+_	Ֆ�L�BfV��n��Bh��S�~*-.��+�/�#>c)ū�����[�]�g&�#��%D!y�B��N��U���>�5ߠ(ƵH2��[�/�6�a�4�=�:F
W����(�J��a)U�)MO�����,ǴlC��^9��ߠ#9����"�%�p� �Ó�>D7�����ɝ���YX��r��W��Tm�#AUp���6�!�x���Q��}�v%�zM]�D{)�sS��m��p��|-�F�4�_�mϤչn|U�Z/�Kt��g���ڌgy+#����(�	s�S������}5b�le3q��dC��/[�۶�����~�c�P����G��z�Iȳad�ʹN}>���
�b��B�v}�dA��b�Ϊک���o�F+;��V�er�8�g<�;NsQ`�W�*�Fě�^��@tb��@��.݅F(��O�O��g��ݝ�u�h���oR7e�O@M�gۯ�g�%6i�[�a~�6<��[�j�v�nK�KMl�>��Y�ƒ4�{>�P��f��nTy�Y6�z��v�; 5�1�5$0a����(h0Et�"��"�[ጶ3Bώ�cp�vD�\��ћ���v��lA8ف�8����͊^�oe��e|̛QE� W�.�ĥ���ڏ0���WPQ 掵4Ji��$]�̖�U���J�'e` �G:�Z�ھ�ި� ��Ӊl`_Mc�	sWn#Q�BN�W�{����BZ'N=C�R�1�q;��HÛ�}�gt�w�g	6�R$����7z"r�N=+��]�{t�mI۽�Hq�s���Q�L��n��Վ�;��w�Х�.:U�8��R�TDU��f�'���( #y���Yśōt�E���	T�p�j��N�i==�17�>=+X륜��v�'}3�6�����{�X|�j��r��{��V͙��N�G�É��A7b��lD�S���6vj78|Q�\�Z6���1���f��^R1�[�W���ވ(_��ծ�ӝ&\
=Wk�N�)����Sw�N����°hT�<y�=�9L�+heA�V�V���M١��	���\�B^��%��!)ooTV�2�-6it�E�-`6�d��B;MYY�R��uXXB�"��֎�-U�����,�A�XA���3e�$���rͧ)��s'M���%A\���ce9wPu&��F
wە/7�艍����،z���Z�
���z���W,�՝ ���GT#���W5��V��˲���.�U4�u9k�wF��G��ݙ�-������k�fo��=]ز�����J�QfD���B��x�w,��Am�tJ�9����ߣ��㱱�@1��-{���k�!�yslr[Sh��h��I��)b�^G��s�T�un�Ĩ�t+e*�)���x�μ�2������@q�R��sUѬ�V��='�4�S��'�(�f�M'�!s�j����<��?�˩�͆�5�o\�$Ia���.⸫���1=iu]q��͙u-
��~}�R1(�MG/u^ �F���6��_M윎S��B*��e��v40���]�K�n��<�,;2�5����H���bn�<$xS������q]b/n���I�� �@�qƌ�e�*YC�˵@�=cO��hu^6�k3㊳����:'N9�<s�l��c���v�z���/*�I=̀f������:����Հ�S��j�Z|�F�ӫ�/(oWR� ��1>�u���������{�T3zZ�G��b�`FR��*6��r�K���z.x^ܱ���i�he��������M�����k���47>��dM'�wiu2�*��<��6�9µ��ЎSx����\����	ع��Cʚ�S� ,�N�V:�o����J>`�K�Mf8J:��0�r�A��c���=Au����R4/�S��f����S�Z�'u���77��($���q���M�����XF�y��p��QZ	糷eD2�p��i�*dN�^B��s���-�]wM,�����N�.�$�I*��__���Y��}�;�r��u�)���6�PD�2EEv�����U&�D1{�DU@Utb*�"���l�QE�5Q-TD��ɡ�TE�����Ѷ����탱���4��&m�5AQPm���N����b(���<�`�����4h'mTEUT�WmT���4��Vآ"���F�	h��t���:�m�M�5LM4��^N������Q��lm�L�MQT[i����1ET�TUv�h5U2kMP�h41Φ*��4t:
*�#(��.�B*B�X��B�
;��j��%����0SD�R�3!E5Z���/�R���.&*/#Iyd�(��h���5�)�b��}>�|{���o�:�]��K:��/{7w&� D����[�����|�}f R>��G�X�9X�՝-�,T\�{cu��%���ŹRwU���If�8~\��<�k�v����t���Jl�|�蟬੃왉{W�P2�����q���^��[@P�׆����ݐ��;�HCW�qAy9�������6bo_-�z��m��h<���\p}bΆ����Ҩ��m�N3c��bu�az%��\�ѫA�/{v�s�����a�L�/�p �vqb�=11�yFBl���҅-���ڵ5�d����<�ox[��&��3�DS�~3�(�ȸJC��郈z�n�/j���ᮐn6�K��3y�y�Yч�1#�11�Z>��LU��Qǎa�^��O�e�z_��vO�7�M{ ��Lu�Tu�O�G�=ƘsкXr��\,L�D�ʎϣ�����};,��M4���m���ށ�2��u��^x��Qm�it��q߃r5�U�_��m<�"v���U���n��G������a��[R��DбF>��;��R�ǆ��zm��5N�UV�h�fާ4��k����T+���«�t�T�	�#,��z�����Dx\>���͡�Ӽ���S��[��������h'K�w3��"u������V:�(�t����F�5��Z������t�1lS���:�mꬨ��T��[6����N��v8t��������*��sX���P.���i�"c�>�wlL�5�A賤��1ɖ1ۢ�Fٲ6�}��IT]���
a��X�A��r�
R䯜�r�ǖ0g�l�rj;�Tsx�\�^�Ns~�7i�����0.F�N'�@����]L�����A.����R�rim�\�8�L���^�SzݨX�v8�,։E��V>��ˋ�(ih�c���Õ�]-����k�7Rx�f�f�����=�A�qw]Pm�.�l�n`E㨃���ct���ր�c����A��<V{.ߤ�Ҝ�9�evUݞ��U�5�*:^)�=��OF�`}���x[�ˎ�;7*�����W����������<vg�k}>m\�v'�
03C\�*Ջ�!H���8�wޓ]S��,@��T�	�CT"�=�`�I��S
���®�,.�����0O!�zí294��ƪ���M$�Ӛyo�&�����>����	`f���8�"�,�ů
�x^�B�p̓�5�I��5ڧ��N�\(>� 	��x���4Ֆ�fU�p0ө�q�,gl����G�ǃT>�r��bYߍ�4�Ň��2�hN���7'4��n]���:d8�c��)R�y��Ju7���/��f�������'c�;w}����(� �{��5��3�]�X�AiEv��d���sy�9h���r�f L �^>��N7�Z��D��^��Jc�"k�t
�h��X�{٪_}�f5o��.63���}:S�Z�;��:�|�9��:2�5�#�iV@m�T�M���S"z3�R��jc�mꋘll<����e���7��M���~���T�_˷N2�X"�`��W=4"0��]G�6q��T���40o�Ҫ/���º�r���q-8~p��Y�_�2%r%��]D��f:(��@��.���p,�!
Ì�Z��nۗম���j�&���5P�g��{�Ovm�\�ua������|����(S��u'�n\,�oyvIl���u��w]?d��Ez��h��x���FK�>�DtX�(�Ö,��1y[�W���Z�Ɔ�B|V�o=[���YFN��r���r&�4'���}Tt]];/������^��;W0"X�h�Ofi;��FGj5p/���S�&���h�_@��w��9�(�|���N��w��3q��@a%hΧIN��ƭF?m�9W��'�	bJ�������_�ry�аwV���ٴh9I�=6�5�5������D�1{:p�����[��892���h�k��Dp�Tˤ��,�,�m�@��Gx:���#;��HΙ2��24�3#�tݩt�Llf���2+�ht��8�f�WiWN��*��x����W�g����ѱw�wZW3U�Z����@�G'��ղUWB�v�Bϕh��aP���T'��}��*����9�-�nj��U/n��9W0� ;�Dv�jI���g5�b�1����� ���j�5��{�8t�ح�*q��4���#�'��hΙl�wװ���lN6(1e��N�����p�M�q���MO8���;��q4�8��ǩE���s�+zuxq��y�E��/[��N��Խ�׻�6�]�5M��8�b�+�Qv�v3��G?4�
����a��"�j�cq�ʫu��	k�oۮ#�fЇ���5��T�*�q��/�2��@�g)�����w5P�75NlX�x����]7����U�3[�r����k}9Fh������(��l�Ū'������U�9��'U�94ÐT�7%�yڷj�mz+�gb\�E��G�o��=!������;/�O��F�I�����
��amϤչn|U�[�;X�b��.��s+��̿-�'�j^_MQ);��"y\@v�ԋ �x��Uc��T�Vu�|�����}9��jyy�q�N�Ɗ\��j*h��f+�uNM�w�ok���[��iy�)tn�,��ЭF�TT�6��4���'ugM�&6qSo�8l�N�Z��ֱ�Z[���q����61d�u7��x�7Ҧd��}��_<���z��޾?O0��ZY�	�+�B\v��"�lZ�\�P����Z�U^v��������'�=%1�S�E~j�#BO�
�p�@�ޚ�d���
��Dp��S������D��,qYѯ���t=
����>���VL��D	&j�@��E{�l�S������~�d�c!b��ƛ��1�Q��fR=oD�\v
��Mq�z���(s���:��a�3��A�<�c2��8!WC��F���U��Mww�W}	�9�˹���Eޤqh��� m�)��]�E��'>�X(����-���������
:)�\t�J��ݗ�nzu���m8h�]���Y:֢c�W���pA�^8�1�=)V��$ӣiE�ɵ�%��kv�$/���p��p��v�G�11�yFBl������M��u���Q:_��{"/>�l�`n��Fv�h�����_g�ICHy���B=�Q�{qO�/+��q�Y��m��]Yк[
�11�Z���Nu���qLx�'�:P�������Ls7?,V�ĳWqk���|�*z���&6�y{�.���R@�WN���q�g
�V��>;��{��U�ワ;�����?�{��uw	����ٜ�<�8��wM�p���7�s ��9�����kC�d;k�_W�W�V}*��I���EM������7���ߏ��=��s�?P�X9���Tv}�OJ���m{�F�Q=�5�J2"#�n��*8\ژ?_C��S2fX�����/�ؾh���۝�%n{#
y<�� ������	��/Nv�b������!���U�6>��ύS��{�h���}�k�x��x�2��k��H��;�U=�a����鼄��p"��n��f���78��#�=QZ��;�`�0���61L�f��}��IT]�z�p�8:hs��g���e�b�9s�3\͘'4HG���;��ۜߋ����TX|f�b7�o�Q*rD�Wt��M��9~u�h�ũ������^�^����+���k�jl�j5�PL�A8�T������1G!NK$���%�]PP\�9Xe���R���(5�0�^�@�h��݉��sE�YM��f9�nh���,OC�:h���7@�p�X5�o��6�v�{|�Y�{��O�ƒ���vi�f1N���@�+�:Lg�'�S�ր��9�!������3$2�*��I�Ou��K�.�R�VV.r��Kq���ڗVn�9�_��>�W�u�6ZKACry��\$F8��v�
�%CV/�J���մ�����0��
<�TE����2yH[��ɬ�dҶ�I��kw�+����T�ipK&�����M��;��	�B���8�v��_�/���"��kd���h8�f�UG����i�<�d�u������]�Ga��mm=Ơ>=W��k���`�����Gg�.�j�k�����gK�����9+}Z��q�����E�nb�^�����/n!w�E�q��Zx狫������q����JoJ���N��^�=�؛�^��~���}X^fv:}n��,���N�ۣ*W[R�c�A�����"%5��_u�;K,��}(B��<6����z���*��� ϯ"�G�C˞�o,xdԄ>���fc;�o~�˃N��j�PE��D^�^�`%aC��[�l��7�8��v�I�-�M70}���'<�j�����jJ��"3�F��Zչz�5�1��a�3f�~3E��^l����}�ڳ�>�qV	�Cç4�iW��ݷ-D�5-�����p ����K�q�´r���-�C��Bve`U(ɹB}�,[�����>�r�iymK�k!�g&���N�o��]T@�VnQ�4î�S6`�:�cTX�_ߑ�}�ew���^;�u!p��
Il�gz�3��7(o^��|�������yG�;)���q���]u�����\=��ʰ�k+�^F#ʚ��д��S��ީy�8G�q���Ϟ Ქ�/ot��|�4� $2.2�#�C2i|̤��!j�;Kg����k�ra(��e�Û����G:�[]2��"OH���\t]]�N��F�a�>[�Ep�R�f�����}��F�8�r�{�ݫ���3� �[���1��9�ɹ�k�֫ͣ�7o-9��{�%�l:�zf�IN����j�L?m�U�%*#4&���n[�kf&2�0�N�ʓr���r��TGt�{~���M��.��N|Uم�Q	N�IP���Onnln)���Z�
�7X���*�����P��Bp��}�V}k�d(�Ss��ىӹ��)��G�^	X8���@
'ei|�2ݓ���=ܗ��%�!oܜ��]�Z^�c^icqť�I�w�; *��%�C�2�a����ޝ^�}�"3C/s�R�۾��z�����!�??4�^��s�.�K].?��~b�+����+z|	����e������4�Ȏ���<��`�`��_��ޜ��# I.��@��a�ע�Q�.ݪ��L�AZ�h�.5���\�ύ��۳�E�kM�b"ܯxx�_��=!�U��W-Yw{K�amW)c+j0�U,rڝi�ּWgC�	ϝj��뫮�h��<���*XY��&'S^�v.VxQ�hjK{ܙ�J��O:7��]���	˪�燀�ӷ�qn�X�|�����_V}|��*���n�Pxo�7і�/��Kt��Hh�������3���
&F��&�b.�"pu�0W�Ϥ�F����j���n�Th��q�׎�N��P�J���4�Ox@5��Ufb<*\�XB��h�I�r���UnW:���J�ګ!緕wV=B9���MM��1�s��������D?*���ԋ�������ET���Y]�l�z2�7@�����7]i�S�ߍ0�Ã��k����BȦ�.��%5��!
|I�/	u���O�<��L��ͫ�hؓbz�ы����ZPb��T:�R�'���B���<s�t>�����u$7DˏL�VL�|k�`P`�X�=�P �S�c�9����J_�1���1��V2RY��i��_.��1]Q�3�E��p*sK�F��^��eU'	��,��Ò�T���2�pU��?o��;mV�v$�r�+yt�5��^[�'�=���@�!D�b�(�]tr��R��K+nBP��r�=]�V!�S5wN�U�7���hmc��<�^��S�n3���''Jk�C�@�-��mՆFf�tbm<��D�]��X��s���)i�
	��A�};�>Ek� !.+Y���ŹB�yb����?������+�Ћ���7(8�<�^�7f#s�:��n�ո(��|��*��&z�9�}�x�m#�
:��	�ؿ�a�:���o�x�a�'����s>�^�?)���96M���S;�qa�5"��Z���,b�i�8m����#HAM��A�>��N���;��y|���	�6v�k����<��.����Z�ܿV�ހu���*�Y���������=Yр.�Č^�!��hF6��>��	�1�E����|���#]�2&R4�s/�o�36:�v��`oE�g�����B�a�}�(\,�99�7�鎧�ֽ\�ܥfr}��'6�D�hm��U�q��eb��}}3��9��!��V9~��ֆ�,N��dEu��Wf�ܽ7���h�(�����f��C��U�6���1�]�<��Z�3�\������K
�̴݌j�'#g�`x��+��yz�L[�B��7(�j��O�y��_�h�\G��#��nb��?C�����6��-2	T]�	Î3<x����1Hq��2nz7�)�c�qp��}���{m9�B�������7¨ę��8hѼ{�+���$��M�����J�Y���!6l�.�fo���i�wQ.��m���Y�
�4�}h��"���'�һ��끽�]g�Y��Gy�k�M�pG��K<�E"�8�U��=I��)�tWf���X����J����)!Ro���f�*�*�v�P��
��Wt�d�bl��E�4��BԡV�P�ɷ j�k��n�����r3-�2-�����a3��:�
���b�O-f��[H	��7��ê�F|̕w�����W!Hul�g��5s��ċ�`�K�8,�nŕ*⦷�/nn�(��2�Th��.� ,_b�9A���$�<�rj�n��_=�ak�,�fX2gp�F��DEj��j+V(!h4SRec�j��[yU��(���xd�wW=�q�]��V�r6��Ջlb�%�O� �MɍX�W�v6�lŸ�M��m4����Z_;ȗ��#��N���;�lS58�n����1��7V���mt��rc
��R��1��a��1�`	�2ڦm�v��#��l�}t�i�|v�p��ynk��������FYi���Ss0jYm�S�%���|��ft3f�cC��h�WHm\n��r�Ǩ5�3�;XUt�s�f�'^�~�m�K�ځL�;-�����iE3����N�nU�o��X�hu���M?�v��s�n�B�e�Ż�Ʒ�|���xT
�l��C'd���j�9��R�!W��.J}�����IZ%�x^BL�)e����MR�T��%U��Y���UM�Հ�(���K|8멐�5]�xFol���|�+�_�tf�}i7F�c�b���b�������X�7pj �P�ub���_*��O��]k]�d��+���b(;��d\,IM�Gd*��2�^A���J��\�ٝNnk� �^�;�;�p%���D'�+�V�6I}CM���║B�ّn��jrF��ړ�=�pu@���=p��vc�;2�^-o�u�_V�]��̫�t&fi�h�sV�l��L�yb��%���]+���1�	���z�7��k,��p:5�Q8���+S&^�&c'qX�`x\��k)����6�5i�G���oa$VǢ���F�S�;��5�Q_���5yu�p�ǥ`\9�2���E�j�e7��S��Oc��WG�;���/\Qw� Ŷ�d���E0�=�^�,�u�.G�*��a@j��D�S#Ю,Ҫ��{Y���D�Ԅo'nt85����V�����c�Y|�V�]J�\S諐�)��Q��NJ����PZmf��u^H��45D6�� 3�s�6�TG&n���2��@�b�e�e�e����3���)�<$�����)=ذ/���`��*�=��MsW�WT3�Ж��Q�R,UԹ<���)�Ì����-g	��q_C�櫅�d��å_@Ec�[�g=�9���5Y-�� ���aySC���P��u�7!��e9���!���/��I$�4h��.�� } �0)&
����!��뾙�R�@]�l���>�hz�>J�GC�l}6j&64����H{�􎆐�(�v*����:�:MyN�2�S�o8O<1>`TLy�P�	EQZ�
j��<��ȪJ����JC݆�����%n�X�cPDR�IT��PIG��J#�AF�,m�w��5��i��N����"�*�~ �2�OEj&d�&%�&=�.�+X�"��Rt{�'�m�JP���<�1�Ӫ"�U4�UMDQ��妒��N�(e�1y�IKT-U:��j���o 4'y��_t=�{�斅�E4Dy&�F�J{b�����QF�P6���J���h*����X��Rj{��3=\��j,��M�Gu�a�-���~�{GpjN̔������	���`�3e"�9��`>�ZvtY�ױ��� >%~�N��G�7��R�7&�Ԯװb�,p3>^�f�5�7�7j�*�����.e[��z�Ւ��V9F�0<��[4�����5o�U�H�	<P0k�p��z�2�c�:���f�v�9@�kI�d0c�b(�τ	0����p����`ײ��k�z�� _�7��݆����ֿL,5ENƋt��gE��:&U��@�+����\u\�7\`\��b,"sn���;ơ�l;�c������'S������:"U�3@�Bk��S��k&��b�Z��?L,�řӆ�;6a����6<��V�0��>�*���[Ȁ��I.+]�=�u��u�s��T�W��1�0B�۵fK0zOZM��-�b�:'!�h�(gv���{��KK�t"캜3�#��a)�*e��5{-���[�>��8��P8'�������Tɞˍ1�n(���{.1]k��P:��@�RQ:{=Uյ0��>��>�6�I�WB��f"����m)�3�p�7�L T<�ٷ�/��� �Y9���-���Lv�#�¦D5h�nV.�k5g�:�z����6�įƕ蓘�snLI��E�J�"Z�]9h�C�T
ԶZK�ho���8�8;j)�^��ձ�b�LgJQ�v�kd]�h�e�WY�&7a͝��9�[�3#��y�'-M6�[���O�R�@�*W�< ���&�Js3\���io�5�F7�a�����:-�`�F�s�y5��1L*ط"Пlm�&�������x씦4�~wg�B�%�p�5n^�j�~ޑU��	m�"�&�����L;�#�$�D�VK�(J�@�9�PcJ����j&��lA��ڷ ɭ20/B�'��z6�T^7�篻��K��QBè��U��r�.�-��:�XV9p�j[�d;u��9�̚u}��r�k�'�:�Hk.A�~�Ɏ͋&6�^��G�9����ɜ��Dն�	1�<n�~���Fv�Lc�r$��_�.:,
"��x����o����=�u5��(B��1�rX�u�2�r3�N+�4Ap2����0nG6�mD�t�������Diw��l-v��0�lΧIN��5j��*��X��`�t�nZ%e۫n�-9ԵIܪ�.�=*,�Dw�7��=�=p�!�����{�_p~؀���(��i�0�5�=��ŷ�8�C.���O��u�xώT)^��m�;�*�В�A� �φa�J��z��ƸӢF��4�&��~�I�#�#���:9�˸�}ꆟݱ���{�`���^;-+{��)�H�ɿt���J�|Om�J�z��!J�r�>xZiѧ���2q��S(򵏆T��;u��^^&;���wgK.�<<=��m��[��U��@����A�dxk�/�X8�S�OJңa�[�U�a�l��Qu3���8���-��`x�L8���VT��\M)Eű�Qc.��9[ӫ�#�V�H�^�������}��-�fol1�%�Ă��b��xY�.(>44���ԝ�݊-C���zxUw��Ȋi��w�,�@m��Иkwm@6��(��Ip�՛-������j�,m���X����Q��Z����,S�!� 5��:�g6}��4��}Q��⽱*zzٶ�=�� `xa�;��V.��
����a�ª����7j�b�r���rմ^{���ߟ?Ua��*��3c�G{�s싧��,!zm�&��s�U�V�`�|�N��Ӻam�B:�����jj�ڌi)��ϱ�C�vjh~�h�"�� �n�zk���)���o���oޖVo�lcϟa�cU�8'�����)�+�B\v�Yy�k�F��un�#*���Y�⮢ƺpjp�\��v�k�l��Z6$�W�+9� ²�Y.乓'�jw�̤j]FYh-� 4�TC�����C�V{U�k5N�շ	�~4�pw�����������t�ǥ3m���N�����<�<��I�d�
�G��FhBr-�UnVp{3H�z��(k3�[8�"���˳QՇ۝���| +�Մ$��c�?}�W�Gj��;�a�36���u8s��M��$�b�g5�,�%��ޒ;c��#�(�m;|2dN�F��٤�cw�6ܘ��lއ���q��MWk���Av������1ǪH��jtT�KS��3�<Vp��&t?N���l�`�pL;��<8�E�Qۣ��H���@�u/�ƫ8�>Ɠ��>�Ĥ+v���降�g�Yy̝�쵰5�|Tن���>S�dP3Q61i���Lu�Y01�����z|y�E��GO%1�ę`���jw�a:�q�5F�X\+T�3{4��\�1"��m���߁����
��ת/_-�Ǟ���ж_����q�r�f��#�W1���V��7Im�]�XCꌰ�e�N:�&�!�'�T�d7y_&꽌/SbF�b7��pm_�s�u��z��&b���5[zM��O2K��p�,A�u�t����ދ��F4Þ��Ô�Bl-a(� �|�����e�>D�c��C��^�t���U��`v�D��́���;�nG������H�r_�Ի4�z��g���wM����+�X����Ϭ��w��M��U�cT�7�"��nZv$��5f�.�k�����������fH��6�XCf<u��vX�Ѭ��]g9�Gc��ZolwYbo,��qʛ�6�:t�}U��W�r�<�\��)u#_={�'�#XC_eBl�.yR�]�ߗ�t�~!j��o|�_�Ҧ�"��]2����j��S�U[�۱�z:w��|��=�韧�	��4:hs��؛��z�h�ۯfNNc1	�<��D_ڕ�L��8j$8M���q��-�~FIT]�XN$����!�
݆zA�$>ku�a���tS�yP�k��8e�9�{K�Ш����ՙ�ׇ�i��S����g���O
g�:� �8r�J߭{-�����:�ڛߛ�
���c��7O��
ɂN�_S��K7+r�
n�l��5�L���=Q�Ekk�7�Ӭ�mF�	��B�,>��23�T\Ű֙74A{!�hm>tpj��J����J��IDd�qL+�A�oxq�EH/�J�Jr��S�d0΋0���T H"��c�Ĉ󔯪� ����Z��Җ�g����O0֐�x�7����c;>O.g���F��!H�K��][}���g�-��j����s�^�
b��o�������E��V��hlJ���일�����>�Z��\�4?[U+^������-�s���J���� սrv���g�M��HT�:@��˴�̻�.��x�MM6Z}�%�r�1c�[���\f�e3}\j36F$�n�Af�?׳���ZxcȩMx־�]I(0�fU	�ѵ�L^ձ���  	ԼR�.�i?HK�@�0��0����љ,��'�&�q����b,nc�Ўg����rw$3	����gP����]�+T�	OqS/Vi��#�[�>��8����o�4ۉ��z���BƥC�k�La��;8���$P=�G������F5m���8�/B�D�lZܚ�YU�Y���C~����%}����YR��"X��J,z�Y��u;�7�sC�'ľ1Hn������Q�IB�{J��浃�}��ۑvg��hM1ni�w^t�Kj2 `uv&��\pt�C��}�}��Y��Ib�-SV��v�8�i���ݞ�l�ir��42���e�-���Q`T�'�@�9��(!cJϬ7m��SWKnf���nx��S�w�̷�!�=�Np�诬*�����Ô�)��:uO9�c�0�gLw��⤟jI��Y;]��+m��9�c|�a�t�Td��_��,�9ٓC�~l���g�|�Nז9���T��Q$�e�1�U����N�ۗ�5�*5�P�}��Ɍr.D��=�+��涏>��1:y�Y�n��6��~E~�dd[�i�MAP�h�ő�| ��j)�Wnk��32���U��m9���b� 0�@�;�����c<��g*��<eũ:���3/��EMeU�	��� SZ��������O��.���تK��X�SH��l�b N����^�����q�u���l1��O�4�W��8�i�"t�$S`+�k�2<�,S���u[턼��^����y跎6�o=
6�w��)۝ƭG)vl�,��n0� ��UH�*u�ƴA�Zc��qƀ;5�"�b���ㅰ���K��Ӆ]���n!md�M���us̼���j�艋`e�����S����K��+�Z�Ց�r�k�4��̀��.l1[[(��{v�G{�C�&���<����HO�#a�^��@�
�0�9	&A�6��R�;��ܛ]R
�F��-lQ�[���O_�(����(���a��r��Q��2��2wFꨧތ\bO��CI���z���`��H2�x����_�CG�~l���5ˣ���_N���wC2���WBa�>�� �W��4]�62fz��5��iG���d=T�޿_��о���-ǴlC���<z1��=#�E+���\�W��sԋ��8K��P��R w b�g��3�&�r
"���^C�Q��7�u���F�T;3�z�7x,upG[��r���6�ޫ&U�}8�3�K$ϻ���۲�O���3}A�	l��(c�e3X�:�;2���;4up����4P\ɦ��@�І�z��H5�@7�vA�K�2gr]J��{hDT"TRk�Ϟ����z��4�6 ��j��Y�8�>/��X��_�����'���<�H���g��-�aP�\��r��Y���.���66��c'յ/}4DlX��#��ȇ�W���JT`��|9cQG���3���8T�Uc�����8�w]id|mL������>ܹV�TU�jwo�k��k�u�"���S�S���%��v���j�x#`�t�Oi���<C�L���NG'�l��b���n���gאtyѫ���tk��s��M�5䖋,1^��&Y�O���^w�q�L��m��lT��2�Z����K67�7=��a��]������J�������˞���f �����0)�*lT�KS��A��V1���������7��ڦ���%���0��88'�0L���&&��
,z룔љrO�K�$�	3y�LNp/&����	���8���X��6\b��b���-A}hQ1�w�]�S\C��j}���L��=�rl^�5*�,�L8�ԋ�j�������.f�*>���8gs㜩I�'��w�S4�L���;��6��`�X�k@�W�sE�u��ƓU�/T��eL��X�'pR*����%�#��]v��^f�Ş�8N7�@�f�xW^s.�����&:�χl�|
(+�V�ʅ��x�+��� E���U�n��Y�n6���
���Ќ��G��������T��n�F�b�ϣ\��/��{3[�7<Z�)�����������8ϳ6�à�g�>}M��LC��Zڭ��]����	g���~+cnYm#�1�d�8�H>�\=٦�p9���GaϠ���{uc#�g5��V�I�]p���ٶ3�|��|���M8f>��+D��<�M/:Z@��ni����h��˖M�O���P��$^=�f̭JŦ�P203��79R��蚱I��]����ٙD�#zcaD?=<�5��:�!� �7�5J�UV��o���ӼES�&�韧�	�AMp�)���=���g����']h���xG`�qF�S�?|����A��p6V���s�l���OtA��V��y���,<:htq�04i���7H�����u�̦*,�lu획�~��q���qٗh�۪1=7"}���JL���*�ص�X�b�37k�joN��ХՉUz.j0v�_;G
�a��=�(�d�A���G6i^�y���V�;����~�yp�&^��G�)զ
ꝰ��ۂ����`���08	�*__���bo�v�I�����FMc���ٮ��r���;�Vr��eڨA�wN�S;God��[��7�l�%�{��K�p�Ax���u`���:�Ƶb����a��|< 𗠞u���4U���6a^��:����쉯�D����=,PT��c��aq�+8���Q�k��˦=,j�Wl�p;�	�S�NR�C:,�)�2��B�+�c�n��#]����iXK�(tc��f�� ��ɼ`3y�^N�3������M;�O'-GTf�SuE�E�,`�@����^츂�QVـ��~"w�G���͠��JǿS���K����ޒ�*���2�ɹ��h]�^s�6��<:���9+}Z��		-�b#j��-��q��j��LOc�cP���<Qv���f(s��ZD	����L�Y��<� ����K�2,ג�z��pQ�yr��{v|�=��d=9������V�nEט��9��1��ҋ��UK�C�38{��y�t4��ӡu1��bN�H�8���6�*Vug�4���Q�˻�i�w�	�O-z5:�d���Qf��n+��GB�x��[��v����f|�.��4Ŷ�a~�ٕl���Q���E�(T�A����u��(/�5n^�ݨ%�c;�����},W]�uކyz��U
70��d����$�c;d�̠WtW=׋E��K� ��N/k�bK�>[�ro+�F�t�l�ѵ��in�[�e�c��/X�F�}�HqR�Sz�d�:<{k@ı��'C�P��72c+��C��d�
+�M^����&��W���8�-Wb jv�kt[����W;+Cpyi$*�kN��)�,7[<����F�C�zW[��VI]��N�ů-QL\�Gc���e$��}%v��[�̉��b���m)��k�rF,"�³a����ۧ� ���\z�R���O����_Q���2�yr�i�p�1����3�����-���k{���4�ŅK�q9�� q1��RJ��ȵä�O�׌��Wx�陻S�R��, �A�����%� ��KLKF����������҈v��uN�aK����2��sk�U]���<�`V��!o�q?�]�N��GEԽˋ,
p&:,�J���1�d����A-;o�8���VN��wZ馟R�ŭ2�������������sPw��R�7*!}4�d���B��E�����o`���=�xJ�דpSB.(��.a����]&�	}��fX�����zn�rh�W��]7Qr/��h@$�W"##o:K�F���G�U�
�)�5g��Y�l��S8�mf�(Z�Qu9���9W:(^1S
o-��ud�8Sы�*j��G
��mAB.��-AQ�KU�x�����4��83d9��6��LJihh�y��xf�L���Q��6
7vN�Q:��i
���u�[�\�	�X'*/e�����1�Vw"r��y]J�G�J2
)�0w��PR�k{[J���+�C�p���H�9p��r+p�Y��5}��Vkֆ��b��=�L�ّ�C
���&2��1iycV&f��儌r�]lt���S#Z����JXz���$�WFV%S\�FW����+x$gh=�{�I�^ֳ"���M������V��Y���2��Љ�M����{��֬�&��_=wrgI��$8)�ѱ��kJ��v\�)|�q�`���V6�W#N!%b)Ҧބo��r�t�����o8��@tb��qM���	�Ȋf�=�7�������P�6� �kI)��*�O;^�k��JҷUp���+8*��.��cƮ�9IEX�WA3��3t]��ʑ	�1Ҳ�K��Z�OT�LL$���'7[�؄�!�'��s�>��)��9����v�4m�cFU�٣:�oeJN���pQ�w�CV� \��wE�b�� u�Pe�.	�0
9�Y{�{��)�/�e����e��+�#B�Hl=tj΂�6�KYΦ�j�ڽ%m�EKi�}�2���=�CQֹI$�ou�$�������X6�f�5��c�ƾ��\�j�w���q@,O�[�mN�f�Y�����4�NjR�N;��*�R]�I$��`�7d��7jë�k�sM4�F���u���E�ԕ10{bi�����f""���o5��0y�M14%'��x`:uBSAO���lkTS]>G{�y�L{�����6((6۱]Tlh���]&�+˧��M�y�S���K4�TQ���'�k����f�"��q�;��y�I�=�E��~M!O�E:
+E���G�y�T��lۻ*)����ǐ{����)�g1�-*
6,_�4TM@P�S4�:"��"����Z�)��5�4�I�X�+�iu�M��F#N�#]b���1�<��8�V1m��C�����8��5����sSHV��5U�*��Z}������Tl`�1ڌV�V�C����;d�T���uTh��4��kQiĚ��z
��>��_���Ѯ��D�:*p9�)L{��7�<�y%�+)t��e��ɮq�xP�)*knÝ�/���ɣ����u��������
q�M�f��{0�6�K�g�*J�Rs�"���q�nY
j���-��dO�ə�!t:�o2���bUi��N}�z,���8�|r����@��S�!�bz��D8�i�iz�'=��|f�ܟ8u�����d���^ �?vd�����#&6��"uV�M��q�.vn�v�pE�jdc����7^��wm\�M��r�
�����mEtS���=��1���g��Ϙ��@Q�K�7Rx�s]*�g�V�D��8a����ņ-���	��_?�O��/ �6�!�o=
6̧)N\��Z��q U�%Ҙ̜rg GR�-���pB�A��q��#�9�oaJv�(tr}����8Uٍ����d�T�<���c�������>�ڮ�`c�nA�a�L(y�zVK��p]c�$)���P��:xP������&:��r�a�ϟ	�0pL�&�e�P0p��B��ZTc�=�n�mXd�֒ذҪ�[�^͖`m�&��6(1e�����E�˜E�������SM�}0럵�6g��?w��~X��cZ�[q��]">W�넬�fN�>��a��0_"=�#�e]�j�>��qq]c��(U��N�Yf+�)MP-Nc�1�^��[z������,O�<�����ύ��mUͶ.r����������2m���_6N�Q���<ɜ^������ڙo^�3����,t�1;0�'�u��P�l�%��r`��F�1��8�)�s�Y����WBa�#�T�!\.2�/ͬ���	��h��� �rl�Q��߭�@n�o�,S�lC�[�s�<7����+D�/x��L�NQ|2(�\p�	0G(h���'Ξτ�a��
����{�:l�W���17I�C=�&�;<�NI�C1�jf��N;>��1Ⱥp}�XBƛFcrw�^q"9˜PI��u��K
�̽�c!�klOm�>��fA�
�=On"��07�J���E�I�h	��W��s0����G7*fܦ��Ǐ��1�*�0����R��~��?ܟ�	���{ҡ�&��A���M:hm�;V�lsyϮK���%<]@j�XFĖϺc:��ә�zq���S4>�l@����������	�~�^�f���t:��>�M���3�+�w�7*��n�0���TL��P����*aIX`�.���RY���ۓ���p'�:�_V���fX~T7i%N�	2��[�\&��@���-z���^�{9���\�@��D���	��֪Yc����~f�r��̩��S��GJ�}Y�aLu��L�P���i�أ���_g(����D�*L�sKGw#���}�i*y��{����#v �7Y��z�a�t�,څ��$��$��S-N�{ �X5���(D��nf�"��.�,��������8O�?>����!@�z����S��K�V�A"R�铻Q��9q���	�(��ar�^@z���NqC�2\(�2	���&&0J#��TvU���ݙ~<Oxg_e�	�f����hN��bw0�ڣR	�>��Y�.f^g*̿X2�+��d�4��ִ�=�댄�GP��<�[L�B�7H�Aj�;gѮ}b��>�t�ه���y�.��I.,[��������+�5��7��>�Č�z��߭��Q�;��-������c��e�:nI�1��↸Q��ۛ�,9�@�ط�������(�zqRVj|h�KP��?����=��ƾQM!Kӝ��p�4�]6V)��}xE�<��^��؎�|x�����Q};�U�^���<�#��H�zs��t�������cF��b����L��9)�.�0��B�(1��8nuU[�p���E�NF���}[�z>x��nl��4�*��3��w�jʏS�s���ٵ��0L*�2���	�uݙi���5�t��bf�"��_e^��)���ĵ���'S���O9��3ĸG��<m��绝��#�ڴ�,�<8V�,$ӕ!�*9P�(&̫g���N*6�q,�xxh�&'Tq���ꒄ�
�84�CzU�_Î<p�j�8O�lb����-��o�q���\�.��Ғ�6����B�b�*XRp����y�E�e�f�������5�	ݲ�Z�5
߳f]�\ױ:`���\S?;:0���+~�������l���6�r5a���jU��뼆�;Rak�gۗa\�g�������4ϲ^p��@�����{�T�=U,��B�_�%�}�مo/�r��=gdMt��t'���T�V>��Cκ���܆�6;�V0����~�m��t��m�JF|΋1� �Z���4!��GgOk:˻Po*���B|��Yq�x�c�x�7����c9;�Q���F��ixܮ�gK:,���"X���ߤ��Cr�&����P0��S
���*��/AR+�6�"���h�}��]�Hf9����q,:�jb��슌l�fD
��&��HO]k��A'���#�=\�p���h��0��n^��qiL%=�xLІ�MYo�k�0~٭k75ӛ�`z�{�u;�7�lyd�c��D>S�X��㙩S�^�����׵�LY�
�������2�3��*N9~ڇʽC�8��d��k�i�Q-���]r`ضY�mDsrՒi�Z����jbR�Ҹ��S*��n�1�+����
wm�B��w����-�7�-��q��mK3�5�*�nGW���-�O0�׍G	�-J����;9q��P~�S���1hO�9���d,긚�1N:Gz���V����xז%�1�B��7�^�e��K��Ppޛ��g�n���O��j;)Y�=�q��F�^Y1尡�4`��'ދ�X���"��%�p�)�r��Pe4�k�L�}����Ӥ��f[;;�mhh�����h5!��3�#��Ǻ�)J&���ט/�T�Wն��oi��c5��e�
��k�(�0�22_Cl��t��yɶ�9�Y�E�����w�Q��w���Du\,Wd�ϕ,�&Dt���:��X�)�Ö/f���.[��ߚ���ŗ��S#1���5ֹ1�҅��L��"�M�=p+�P%�FYY���N����>;A������t&ҷT�	x�N��\��b�T��Ȋ�cMr�#�C�����8���s���H����8�a�n��F�Ir���ƭF��v��s�:��V����M�;N��/t�Bi?�&.U��m��PWAf\��O��䖼������
|B���Z���K�ntuu�'V�����B�*��]>�]6���b�&2���c���\��m�\3`:"�@��/黲�d{.��}��W�ٜ�3���x���02A�{JZ�2r�h�W�M���ͣ�A���Fh>M?��9�:��y��vZ"aXT"p_���7����d+�Z�
��9f�Wo���[ĥ�nnw� ��YƩ�>�m������ro��`�"�߹��3�E"�,�|�k����#��L������pM���/��L@�b��]�H	��}hn��u�Ƿ(sI��/W����s��3�gyx���0jdM���8f�j"�1<i�8��D卞���㥩��>�`&*<��z8ϱDSN�t�^��n�WBa�ݵ ڸ\w��V^�GY�.J�W��{U���K�"���`(Q���Ú՟X�Ÿ�T�8C[�sso�SX�dqøp�ɬ�ȈɎL+L��Fh��Q:8�H<0�>h���$:�Ɠ�È;�#dP6�M]b�R�eEf�6�����E4�<bM����d��d�����,!^��8����3Y}�{�̑�k%�*��S�UnV��6����z�`�ږg�DlX��#�O$�c��/u��fOz�S$�������y�2�l޶a����/�Dy�ٲ*{���_K�ӯ��1�ss-�B���7��ݷ*�N 4�Pʏ��g]If��8��u
;����wY��g63�|����nvȺVq��P�!��Yu2�!,7��������w���١gHeIم��\����V�����zz�cN�2S��L6�s��iZ�6�庍/�������Ys���s����pjp��%���`��^@��o��ֹ��(��8�����z��tX� Ⱦ��Fvϯ ������t+G�{�ߗqRX�\Q�z���ߺ)��B0KpOlX8ю;͘h9n9�2da�J���),���m�19����cf�aQ8��mO��FFrF;*<�3�m薎��$I�A	*n�:Z�s{��X5�v/�n��������h��З?���j�z���R#� A?mUz�����[��<^��ƪ_��;���'��<�������'bu�09#e�|�EU\(����K������r��%�1���/�,OGf����jw�c N�	q���k�j�of�|F3��s�'�n֟�;PS/�EEx:q��eѭ������VD^r�f07~�#j�/���d�\A����v�i��l�l�^��IC�y��QM�Vd���=Y��[��8��g�E/�A׏jMɑ�Wn
R���D*c)RǂQ�� o]�/v�S	��q�R�I�ᵻ�:D���w�R�ϭ���޲�).&��k>�f�B��)}��"��m�.wc6m�3�t�˕���U�qqx�}�Q"��u�WۂM�}��|h��oS��jUL~ �d���Ƃf��P~��{�L9z&�wT[�h�n�bЧX��������������'۽��ߵ�e\�B!�#sEZ����19jf�_Ll8=���d�Q�ᩮ��A�B�K�r�݋n���a��A�ʗ�6�V)G۴a�=���UO�su�������8�9 E�[��p��ʪܶ݌h[��l��g"��7�]�s�Kټ���|�
�_�%	�]��B4���x��M	��>l�7ɝ���:�^qf��#������ٸhtŴq��4�T.����u8]d5-�Nn����G�{�ڴ��.��y�7�ndę�BC30�> �c�KlZ�,p1�\�:��qO�+���ݛ���7�������8�,��NQ�S\0<���+�=ȯR�%sgt��u�&פn��(�مz�@����=gdK��� ��Za�F�+>��縝��X0q���~�o��?Js�e��ϺD���#Mv=�0H-�^ݨ��wJ�^�/U�q��J�e��좹ک|ݭ�7QY��u�������b���ʘK���f��qۚ�yT��_�P� ��}���8��շ'P��T�=o�L��
�4�Y�*����X�2,]y�vU��r%q<�^�f�<���xF��5�'r��� W�_W�_���@�2<?}��ҋ��/;. �|<|5�1����C7������!F��C\�C!y��	��;5Z�D��3^Z"�)���o���Cr�7l/b�������. ����fDR�������5�pjDK=�0O!���x��^�CD�@;��&��2]̨��c�Ćc���T{�Ɔ�܂ځ���x��n�k��ZDza)�*e��;6oMGd=�/��
�^��ᨨ���I��n��Ü��ZϢ��e�u�/>5�]�@�5k��f��/e
UOf��o��t��v�j�}����>���x����/i���
�U�i@���q���d�}E҅R+�4r�����1�Ib�{J���~X1��=�t#}�5��	.�e����=�c��b�؏q���w�S�F4�s�smixr�7j�GՌ\�L9�=����f��s�$d{��dQD�a�Ӟ�T���pi�+>��ݷ/��Ҫ�FeO�s9��0u�{g��u��V�5��'v���z(XU�N2m
����r6�p>Zi�T��O �%�p����P��������ſ�{�`��A��\��|wL�u����!��C�g���(��z��G�2�}��c�� ���)��R߸���k���+���mQ�C�,��)�,W>�n�q��E�-��_���n�f`�i����ǜ9 ������C�3�,�2#��NE1�̚<������Ċ�7�e���?w�b��df/<7:��!�P�p��q�qA� ���n �����nu���
�C<yx�h�~��<��n��\��Dʽp8�x� �dI�Y��.�QvY*��1!讁�}K�;/#��8�a���z|Q�ө�S�;�5j!-�s9_j̝��ݲCKg.o��`m8`��������d��B�E7���n|��73(9��V�J�x/̃,P��]U����Z"a)���4����Y.�u[��#i݈���#��Y~d�3�����'���<�lme��Ǳ���$X+H��zV�V���;in�k�=��ҷ�X!߻=��M���YɋS�g�U�'=WLR���Ӥ3��>��f��uv�+��ۮ�Ӡ�����3�<���po���L����\�3{5E���*��_�r��X4��U��(�V���fǾe�����5��F6��g,P!שV~u��ug�|�L'�!j�4ˊLvڊ�ѻK;Z��6-o-	RόpDEZs�7t�+lt"����NZ�����K��v]�§���]���xp���y:���1*���}�'��gR��c��1`	�
�Wa���7\~���@0r�u��17$��B��ܕn�*-�y�����S�}�#�Y�ɕ��B�g�p������lJ	���{�s��7����ʖ�PA͕9�ٽ�4�[z�g#��@P�ʮ��걘�YI%Y��)��@)�gY��/�t%�5;Nڧ\�Sy㳣�C,1݁�'1.�mM:�i�;a��(\�[/���_6ֳ�K��m��K�ظ[��n�xdѴo�m�e���a�S��m��qp��t���X����j�h�����[R����̅�M v"����=��:�s])>�4��)}+	}�t�7�����F3*j�&*c8)]�a�W4�˨�Ԋ؄s:������� Wg7��|�,�QM�J��Ԛl�v��P�Q�;����HI/�����e�Y�z�OJ�QY|0�lp���@p5/V����{�\WJ�՗dfQ4�	�N�+����Lq,X��Q��4��7���rs+(�H8"<#�����˶�*<���CK,�ɴ��8m����gѝn��/Uȧ�x�ut>lӺ�x'=�W��`Ju�.WF����{os�J����(m�������1] (�"D�;
j���!lË1�떦*�}=�F���T3��m�[F�{e>��N쩫�u]9h��(�g*����d�	�ҭJ3�ŗ�gpd�&iQV�z�N�u*oA�s!�+7��WP3d�BoV��|*?�E�`DX��q��oy�ol|f+�2^��8���ިۮ������/~n�y������kU(D��(�6zΩ}��7c��.��9W(m�Mf��hL��*F�7)�n.j�u�f��iT��U�|���@J�AY��Yڍ�Q�wk2����:d�̀,�x�F�zq;��n��݅LZʁKO�i<ԗ]�8$�"�}�������"���\��p&���g%l�����q�l�r!��l���5Ś��$dV�ٕ�x:]CB�Du-Ĩ�X�n�D�(�{����#�;V��B�68g���}�ҫn���K�������/Ea��3r;�`�1;2u,eg^ 9�Pt1��=�_i�Gd�xA�0��9O�7��vT0Α���n����L+�5Vm&���-A!f���Y�wR��t6��Yź�SNl��n�r��V�֮mp��t�|��*�RA�ٹμ������e��վRk�ϵ�ZƧ2�פ�9�g���7���X�e�%�'�l��ܝ^q��N��.fӳ�9��{uƸj�G�|QI6�F(��]�i-ޘG{L�:�pw�&-W�}�䢪T�e�$�IR�$�1���_m�ܺ�3V��lQAlQDMQV3Fںz�R��֣`�����lb4�1�b�_7�;{�N��M:3Q�(����RO�gZlju����yWZ+�UZt���[��v:�IX���A���{eѡ�i���=���X-��
"%�V����5F����n�F��C�4��ݩ��N�h���&�y�-Hj��N�6Ѡ�Γ�+�4�u���:-j��t�eփZ����Ê�"��b�uED��A�[V>-v7���)k��Q���y�t�0��5�=�qQ�n١���
)=�f������<��� �Pm�ىj�V�=:�Z(hѶf��`�w�tW�5��5].������m%���T��:'��h�::�9�4���wp�PP&7�[q�-jCb��t���A0�u�F�A���������t�����YBQږh_\�3�i�ae-����wnv�e˻��Q�X'���2#��lb5������P3������N4I|��@�_�L��sJt��
:m�sُ+�̨��vk��:���oWַe���{��xQ�/�EK��
9KD�}�"����[\4b�k�����zA��,6�!�Ŏ6d����u��9aS�ʫS��.�n��f��m�$K�p$��p~��8$թn|U�[�[�wl�S�ƿ���ƻ52HqD�mC��u##kA{��+�����u"�ǍϕV9O�lcϟa�c�i��7v0���մ�'�GUU�7U��<+��8Y�dA��~�s���X�q�p�\���Jp2���1��ퟻW�ef�c��فLx؞��W�;�����f|,���y�F��jo]�Sw�z����":�8��j�f�x=�(�ܦ�c~5�0(0h+�$͊�rV|sv��J^��{���O��g�_��Q�6ziZٽ���O2�D�:�f#�s�b�l�i,�{J�v�w�4.�ľ�]~���P�K��0u��Z��'���9@� �[0�k�tmo?5�>셴��
�K��c>z6�(�P�t}�Ќ.,Q�3�P��*�n�l.E/뮟�yg�z��6yEO�nf�ޕ�����&b��t�e�]�[!�+I��S]H%է^m�S��v�&h��4��RL�\�Y:(�1q�B�	j���  K�ٷ�	f寐�'�[�9!r�G�ې��l���9�U�0$i�4	�ػ�m��b�ToKd�0��ձ�t�W�a�lA����8�;�1�'s,5F�Z�Z��Z
\t�m�k��ZJت�{5�m����EE1�����Q��(꼏8�[,�7��Z}�	�1���ą�T���x���sl��8��K��"LC�Sv�3Q�̳��&�U�Zq�&*z|�Wi}����\�Cv��
�7HN)��$��k���+�vi�/D܎�}�]�ڧ-�V����	Twy�$�5�Ü~�p���tNGgў�ڕ�hD0�n}��K��٘�<jh_��w9zx���'6�~</�K��z����~��9~nŵ��P202q�]��}k��H��y�m�~�G�)\B�]�7�!�>�3.���/[x5��9�o�+�+���*�X�kq���3�\[y�pt���-Έ~M�!��s�s��p�:h8L���=/���V�F�ބ�E�9�J��������C�rr`hҴ�n��������-�'9��6v/�u��5f��kL�}�=����)2���Y2'�.��@������.(���s%��XZ7��\#f�V��Ӓֵ�r����^!�&��)�D��Bܹ�����.rr͒_L�5�n�u��""}���kgAB����|Q�=Q�<�~�ܟ~�AE�3c�#xf�ę��Hfn�&s㕎V�k�1�!�b��}5��+3�B��c�34��v����>ι,#������ ���0<�H��7�Pwlr�2����4��^ϫ�c;#O͘V������+��:(P~���2�v�ӥ>�k~����:��Cԡ`Y`�g�+��o��F�Jr��+t���
0L��<�FE�G�E�%�b¾��
�.������`�� Ǔv��{��c;>O.+��J�؟/w'Yyr��}��c��pI�Ü����<E�����fTA>^� *�L.ĕ)��^1��Ds��]�X|+agƆĹ��s,)�i�L<�L*�۵fK0���*�R�I<3�l�h�]C���t��@�����E�l�jk��ZD�P���.��d/�j�C�Gs���/�e[�>��8��P8NvϚ���YNz@ǖ/�XL��HE��x�9�Vs*�b�����秞�ע�.60rvN���<���;]"}Ր�eJ��`���������{a���Jf�X�o������(!�v��W�l|^5J�Ɇ�5�U�FX�#�t������M̽�Rm*����Ȟ.Ѧ�rk3;�iᶨ�rds6�����E��`z �I��lԏP�ƪB=���D�%^e(�E��\N�y�<�_Ͼ��zJӅ�y�O�`��迾�з1�s�����1�Ib�{J���~X1�3��;a��<E�]���9�Qy;Y���G���)���]�p�m�5nX��\��W����|�O<��鷃v�6�E��Q. ��s�
���GE/JϷ��q��N+s�D]K�O�SW���Y	5n�XdF�S��B¨�L�ώR��O��5��j�)��b�/ݪ��Պ\/-�~k!����:�'ZA!���2�Ý�19\���C�Sއ;�R웇��Ll[P#ml�#0/<79���&5�P�s�2c��'���1��&br�]°�7��C��<A�e�J��K�7~I�ϵ�2�^��3���ѩ��v�TTu�x� �V��A�@a���l��\ĵ�FN�Ö�`qF�Jr��ʝOA�3�ʦ�x���ڍYQ	N@��V D�4&������
�џZȦ���:5�7@�3y�$�颻ݱ�G9���Pͺd1mZᘌཇ�0����Y.�u�t�%Ʉ�g��M�uT���LLF)�gB$��L�{ޜ���/x�(��[�����]7½�(�u��Ne�4/7t$���F�_<`.q��;t'��X�� �?�O���_;�G���쭵2���M1k�ۢ�+��)�.����{u,���]W�kO��W�վf�5_�8���.��^�#�}hN|
��U�X�-�#(9m�x%�`��ZB"bL3+=��O�iܭ<��vX��S��,�{���|]6'��90��O��R������w�U����)g)Ԧ�_~�h<��v˭��A�ޝ^�����Y�uG0���R8Nti �\W�,v���쾂�377[�:�Eۄ�b�L�>ᔢ�_��*'j�e������=w��1�u ��z�pi&�NkZ����/��$�@�j�S��0_���7�_V}|X�y<�9~�h����wi\����ƀ��L'q��4_L�(��!��*�o�.�bp�� spK�g[)E�޹0����#�^��k�7f�c���0;�#`Lm�N:f��PMl/�ye��9�w,� ծ��]<n���X�h�	5n[�|������C��8؞�1��ڗ��C߼�q0;yHN�J]b\`���Q�Z�+�׭ԋ����Uc���<}��J��W{T��
�������N��x1_Bc�vYp�b��s���q�pZ�}��ox0q˲8��6�R0�������7ɺ��t��0~jԭ������kfK9�7V˷{%<�F�yoXɰI:��i��'g�=(J���ŜK	ޡL���pj��핅WQ�"��^�`�j㩢����ӐIY[Y�J'�8N�Q�����R�ҹ�\��-(c��_{�_��,�Ω�;M\
���7��F.��n£Ke��mU��/yՙQ�Ze*A�v���\����M��$��]��a`�$��Ôp�2�P�UK����[���������F0��*)v�ъQ�veV�K5�`�4`�A�7S-JC��>wgϲ=�mg҆���1�x59� �U��t�gh�XaGe��udr��@��~�HM$0������Hv�vv�T=���NO���X܅����8����{��H�q�t@��D7|pWΫ���b����
�X�宒n���u�:M(�^��\3�.�@�3=�Y�Bt�v^N�zm�K�v�G�11�y�M�v������q
��fά#�𗽻Ԧ�ƀ�]�Z(��2��7Ip���/Z��������o����PLl_d2�-�/�Cj6[�(�������n��S00�/C\(?q�\=٦�j��o9��.:"����yM~ӣ�lt�Z�f���v�VԬ�9�j\��n���oI��9CnU�Ӯ�DS<�����=)e�<�NxE�=[|���x@7r��I��O�$b�X��{�ch�fM(�Ƴ�EkYs�Q��2��S��kϵ��Y]`�����q,���:�k��8��2�K�-�9u7.�?=�n����u;�����iy��Y������7#C9�Ro=��C;[+j]����~�(����T�������D������	@�8nuU[���{o��ɇE�1��.�{̀I1�o��{�Ы�(׫��LH�!�M�!4���8����h8N6,����TG&�~�|�y�:�����v��󑰴�)a��?���4i��!�@���"�޹ظ���E�n_�"��zq�{K�Ш��͎F���Q�3bD�)���R�8r��.J��Bt�gn�NU�x��=�Yg�@��fn�����P��Ɂ9B�,��~�.
z�8�&�f�М�u��$��OyK���V׎Ƣ*����}]������}�Ț��!da��Vm[����r�;��_ѐa�AӃ��c���^˷�D#o�S��cm�R1�c�T�1�щR�ݴK�P%�\0  �f��tb��>R��!�x�c�x�f��rТy�<_����q��դJ=�a��`l%�k������Oh⹆n����f�T� ��X�9�\��`�6�lG�{z��h�'m8A��w��<�z	�?mH{Zl���zk���o�s]�w���:��s�^qy�Զ��'9^%L>hV�/���+5�n8���^JO��d5����i���;��u��R|wWփK�$m6p���q?��}�[�o�J�����50v�wQ.��c�c�=f	q�\Dzí10��0���n�U�\ϵ�V6�j�I��6��v[�$q�М��E�,��|�V���{5P��R)��"�V�3�]�c�]u-1i^RɎ�<&^��P�}�>V���N���C~���轮�q��u�/dI/+�n������#ӧ�� <T���f�9�cz�2'a��]LCϟ����Ʊ�������r�[{�n'����<�{��~N/օ�S��n��b�kXpߝ�r��[�7����S��"2+�Z�Fh�D�b�4s�oߚ�k��|�X��Ab�)���q�`�LR��t�[H�������mꊳh��xr%��H48��k�뢚��@�Q��Ga1�vL�PԷ�|����#&��[�'����#�U8f0z�T��U���Nug�G��G���b�*�Վ\�,�dy��8,�2#��NEq�[���<������	q
�v|����1h��23��s�]k��34�L�F���R��Y�w@�V�f�.�\�����������;���'��O���Y1u	Â4�(m�9wZ�
�o9����*�eۦP;�Ti��nQV�V_'�k�`:�cӒ[��$$+kZ��ti>W}�e�ES���[H�|v�P��[������"��C�O��(��DWC�;/�����K�7BO�|,̫׸	�6A2򵈦�s��8����p{�M8w�8��ã�1����.bZ��#'[a��zm�����}UP|���ٵ�(��x�Mt���0�1��n �U�%_�#8/��L9k<�;5�"�E7c:�v[c.��\pOW\3`ʾ��l|������Wf1v�B��DL%"#
��
����u����V��U���ۑ�yF�q�0�i���?R�E����Y
0Ɗ�Vj�h1*�JH�oc^�5�R�w"�tIQ*{����n�d��g�;��$�71৆��UeI�c���Ps!�l�xs�Ŀ�Q��������s������t{��"����,��2'�4O�rxM*"�Ixu:��5�O1E�,��%��5���{%]��d�]�2��x��!��|�\E���J��mXD�ޢ�3����=�>W�4_�d	%����P�Ӂ�-�v�-��	AΌ=�4�R��m�����
�x�C�~����sg6iN}��p�
xa�|��Q�Sy=���/�pV֟��vm8��n�.��/!�II�^E3�R�;r��dQ��?�8�8y�~_{��JȐ�N��-����(rxf)��U}�`�d�H�Y����jg
�-�ݭ��˵-P��+��Ξ��it�B�V��Yu��=ՇA�������=��$�B7k�#�q��H9B4*�2e�j��j1��pN6��6J�ח�l��`\W)n:���O<�ii��
�#��FN<q�:K���%���\ɨ=�Ɵ��ᾬ�0
Z,�c*an�����tU�,�D<�����u"�Ǎʙ�)��<}�����j��w#d:/�/E�&�2흗=_OX�[�W���N;>� ��1N���E��8]k�ύ!Vg��bD{;��'m�9��z��x��
F��}�\F.�"�뫆gl���yѹ�v��O�ڌw��d�^�ٶ͎�R���Jl�k�,��Ń��`09��$?���e��]=��3�ō��7���NTh�V�o^��.�=�ul�k����0}4��Ε�ms�H���:e�T9����C�pB��ӿo���b��?Y�S�@�mq����/cz'��K+Т�ӎs��J��y,|��	CW�����N�F9�G��F+�hy��]����	�.�ǅtLR�X�宔�0���>^V�p�-;�[�<P�C���$f@~��{f�j؃$�FF�R����V�Uy�$:'�IZ��3(���JqS�X�}�o(��f� �	��ܬ�R���&ƉK-�AW��T��ܔ���R���ŧZ�C`M"���F,�B@�������&�g&��,P��$���V�[�j<��ŔkZ��C,�I��ީ�d`��g�uq��2��B�V�s��tPO[7L�냮�(��oU���%n^}�9
�m}`�.l�.�1�O��M2�ϝ��&�@�w3Щ�+Rț�Mĳ��Lxg�}�xn��z�����R+{��i�l��3W%]��W��O����4eG���7�<����xW7͇�9Klխ�_N̕�W:ac�qs��m��Μz���]���J�n�r�LLbR�/w���-���u�n��\K}b�Lr����3;E0�P���Z��{
�Y͹��`R��덚.��O�����9#�ӝx�-�y�Ic:+bh��'Q�0Qi��V�Zmn�����y���
�2�Wק��E��&�c��� VP�z��5��m�t����g^Vk��>���)�:*;#��awz̢�u���9�v��0=}�@��A�;������6�� A���d4�&�*Is��Utv�F�;[ubԸ8�mL�:��stZ.��1�#:K8��VZ_VB��4�!N�5q,�x�_D�ᚪL�P��RU�h`�����74X 7���q�Ieo,�oT��|_S�d�3N�s7�f���Hǉ�x1 �ε�*�3Q��r&��z4�Nq�/wKՕ!7��%qk�]����2l�N
����ո�4;;K��D6��<��x�b�[@^�L�^+/sh�N�r\r`n�"k(�.�GYH7�;@X�n1���o\����S��S>s�m�Ld��^�/��V�; ^��Zژ���ѹb���@T�5� Gop�1ܦ�C�Y�z�w#��k�moY��d���{5z^�B�0-�œ4`�z\��̌ZV����Q�{�qf���vM����+�d��v��m����V�޼�Z.����t�.+�ͣ�S\8��NG����uu��� �:�;�Ǌ��� |��:/&t���m�Cd��^E�rlL��x'^��Q����tshR����������^����b�E
��.� 	���͔����%��c�;$��f*����@|�8%�;}å�X�$gS�eK�������wav�DR�h�u+ %B��7}��Є`����]L��LiO~U�R.Kc�. �pa�t�����6���ċ���4Lr���䛘���0�C�V��VVbHgl��V����j��+v5t# ǝ��,B��cc8���qn+���G��j���]����w��^��7h-颕��;Xx�!�ђ�E����ɜ�#�.��WK�s�.�ڷ�72U*K�rI$�\��f��w�:��V�/~0�5u�F��*�tit=��Et�|��j�U��=���o'O5ѪJ:MV&!�F5�c��l4���{d��Gv��]����]{>L��h��gLA���y�[f�����V�yn��1Ӽ�A�cgF+��ml��ئ�q��=|G�M=M�oHzt%�OmAT6���|wyy֭���@�'V�u������vرwj�Tm��iӊ->��`�y�C�7�骡�<�{��:-�uT:��u�;Rt:qov�j5��u�OOE=$vɈ���w� ���6�b|��`�jاO�A֨��:�7�=wI��GCճA|m��N���Ѩ64�N�ƭ�F�e5�ccGZ:
m�ѧl4:*j�4���z=؋���f��;���:�N�~<�ܶ΋d��{:5��;�J򤢒�ZN�64i(���D�h�"�;%(5������ڏ r1�0�r�;mYP����jA�}�Z�bV�q߸S�(�a޼k9��
��7e����e�Y���ۜm�r�v��2}����=��Tw��o���}V��q�K�rlp!��S�X��n]�9)}���j���G8Q�dT��:��f�0�ŮT[m�7v��QM\da�/��	�5�G�:`��ݥ	��N*%�\A�)�v���xUL���_[w�_p��no`�Q���鍅p��8�<q���p��?q�fq9	��Sfo�z�d�?��_Vz04Þ���/�)�z�1�|��T�9٧�Vo.8q�!�t�xL�!�&��.2��f��q��fp�!�K�rכ��E�P21�_�t��}�[xrߧFT����_f>���WD�(��+�܋��0o\A�����s�U[����k9����}��{�\Yq$W�L#����Ӑ��C��=���<�qE�W1|q��ki�QJ�T]qz�Yx[+E4��'L��6F��-3�Ua�p�8:htq�04i��!��W���8�=Qz��q����L��a�~���͎�o�TbLؑ>�Hfn�&U�~�_W��a�ǽ0��w��}��yb�����{mM�J?\�9rY�Ӕ`���_wk�1e�::1��~u�'�Gy�*���RW�l��wP��&F��<Y\ќ���qЮE�V�K������SnX劺�&�pg ��ʱ���:���{&ޒ����p,�apn%뮸���J|��v@�V�-���B�%]����4�l��ّ���q_]��B�U����+E�`ՠJ���<P3�م{�{����vD����u"�c��A�^Ƥ�#Dz5��Ŋ
�<9`�c��{4K��a|k�Ϻi�9�HH(���e��5LJ�稙6:��NY$p3���qۇh}��������h{_dΙ�f�Z#���4A�1|�e�C21O)��
�!H���wޓ�ˈn^�n ���o��{]z0!��ɳ� 2j��u0h滻b[,�c�E�%�qa֙s׻� ����^���EKNX���;���@��ky��Bp7A����X^�����.���P�뭟����MQ:Mvt��Dp�W=�ze��5{-�̅o�6�a���Xck>�]���ԿC��7*���t�;/a�l9�AID�쭳���#ܝ�ҺX������#"{юĮX�{,M�&?W����˿�ana������� �Y9���M�ދ������*́����¾Fû�2��x5�p�/��OvE�M]�M1m��."d!��1���g��}��W0EMQ�氿�zw�wX�8��,�m�W�jMSA�x5x�"�p�aٷ�BA���h��p�)PQ����3Z�������b�8>���+�[���I�]��3Q7�����i���6�s��F�N9�n�W��T2�v�lNߚշ��Cu<���x!�dv��<H�L���ߡ�Ø��	��	�h���@#�-�
A��k"�}D��;�"z�������s�F�9~SWK��Z6Zj�*�Hϧv׌�h�T��3�y,�Fz��[�K��uq�\��R�%h� j�s����j_��y�r`�ʖJ��9V=��U����z{�ODк=Q/�B�<9aB�/`žX�Fb��s�]k��t�`�jdǤ�ϯ
�=��ئ��uݱ�%�4'�
��:2������^ڿ@Q�K�7Rx�u�2�r[��e��z�vf�	��*��P�N)�G�HbL�@5�}'Ge�s�j2�oz}k2��'.���#�ޙa�Jv�ڥ?m�U������0��d�ы�)�m�bc��鹽�B��/a:��97;�_��®�.ʈ\�U*�T"$�Mp���Rdڡ��z�ω���=�d��>9P�`�X��M�'D*��"�TP+4ǖ�ymi�[c��Mc����J���nED`Ӟ�HF����"��ŞSFt�l%��vz�.[~lPb�g&-b�����7�E�4	nӬ�̖��ǁ:lt����!������%�M�|���W�Bn%x!qT�<��]_��v�`cD����X�Ya+������H��NZV�aw��/�u9I:���q�����K$O��ܻy����+���jՋ�]wk��W�:Z������S�����7�)ዋm�e�0���~9[ӫܱ��y�E�^�`o���-�����s��uV�q�1E|g�t�u���<���ˎ�cw�y��r�:�|���}=�N�VF_XeT���uH2�Fh�c�&�"��v�����$���hݙ��5�_0��1�*؇�x�@xm0�Ǥi�K�B�%�Ü(<0��f�\�׼�+�]�r4�z%�yXC+�`�M0�`*��m^Cߞ,q�Tv}�1&�^ʗ���rj�8��v�c���M�,Eрpi�6���V��+~�c!��q��޳�~�ψ��UO
T��^��o��������ss�m�`/[�۶�Lے�P��譸�#�U��pD�QW��)�'�����(0�}BP�RDw�޳�W;���S�Rs�s}t��C�wh�Gwq�8�g<�;N2�����
F���X��Ŋ������.��?΍9�^ So���u-���9ZSy��
��&K�L�Y3k�`P`�V I3u0����էbƼ�8m���3���cyO��b_Y�G`�R���5�*J��<3�z�~[�ٴ=�� ��ʱA�_-Ng1B:ٺy�0#���֋S<{��zb�ʯ����yZ�\r���_t�M�W���D�Ӧi�.�}�y�<�P�Gw������f��^�CJ���62Y��	��F��l������]�{>�٘��:�D�$���e��a��qܞ^���S��T��X5�un�
����M��ƿi�� ��j�(cF�U�-��A�𛉡��tX�ӎ3�jiQ�V(�,nB�j�������/>���֋���m�]q����&���bh)D�J/ז�Q�d��7��3Bw�ae�B�q�p��,�B���\v2���O�GX3�a�/�p �vqb�#*�}����M}w�_��7B:φ[���㈷�6T����gū�����&K�K��"8:`�����$B���lڔ�;���7y�y�Y��Ԙ��z�ni�Q��wl&2�t���a�^���7^+n�m'�wb���N�r;��^���Fq��h]L9~�P�3���ϣ���jXk�]���k!���bf�"�C,*�Tv���1��7У+���b�K�r���ǿx�dx�?e�F��b�٘"f"�Z�˝�t��=��m;��R��uDO���5N�3N\
{=)�툡�Pۀ��WE�&�wcD��u��Ƴ�� ����/7���/b�y���%��#��޹O#m%��.k�/d)�1�g��%;v�!��ώh������+�ۃj�j����YbMGG8�Z;�뒎�Օ�r�������n}uW:A�?� h���)���w���"�ϐ�F'�}�d&��@���p".y���U�-�d�cLM�s����y�̛^�547��S�6V���NL����a8����:8���ѥ�5Ni���0Lz����w������E�����u����-��y!��,�Ȝ1>wLp�d�����q��F�@�ۮ�KO>)gc��ۛ���gM�����`׶���ݨX'����.����pS��b�\'��K
oC�� N�_¨8fp��]-���Z�Iڀ��͘W�=Ϻ��ѫ#v�0��7�0�x� ��������Öv}�k�%���������)\�o�j嬵�1��t��<����:&]����"~���Q�'�V_E�>���&�#]=m�Unf�h�7;ᗩ�ΒT�R+q�B͇ln�q\gM;	���=<E��\�7q{����зՕ���eLw8��֠0�Z�ϊ���ρWu
�X�S��5�X+Ods����ّ�\��w+W/qg$�j��&M����	�l$'��Yf�-xV��W�P�u�|./���t
��%N�Q��L[D��\ֳ��H1޹Y�����"�_��¤ȟO��ѤD��3���-g����/<�a��µ,C�u��Vr�]���z�B-19�ɏ7���n,̸��N��W`��@o�sAH%�(�-*_o6�R��4�u�g$͵����zW8_��*~
�A��Jw�/Vi��#�߸i��8�r��;c�t�G�ʔ��G��K����]��r��[�����@��S[/�ݳ���#Ó��WK��7eԛ�;���OG���GR ��E0�P���[��4 �>�(qZ}}��蹆Ƒ��G�5�׶�ӹ���sD�&�[4��r+q�7�f���1j�zh�-O���>ϐ�B�����\�2��9S���,�ޚ�/~n�M<�Б�Y�_��(��9s�
� ן��g΄[�y�M�p�� E��#CO��{/�)����d<5�	5�FN�l����{y(K���=VU�nf�z��ܑD�@;j��M�P3�Z2���^��0a�/�"=K�^h�8�a�S8���lpl�q���1,�$O��s�]k��(W�=��&c�ѷ�r޷������A�>��C��J⧷�]*�
5-��$�\�����&5;�{ѯ5A�X�F�5�#4�'�4AL�(�W�_@��z��qFÁ��F�8�‰�R�+�wr��������aX�u%�U�]lJn�4� ��c\�z'}��?"~�9Ī>�^#�4l���tM��g/�
���2 ��/���!��I�����{9��h��E�k��س�-cn��K&�Z�� {G�)��U�w�IZ�NR��Xըϟ�� �`J���?hM �7�Ͳ�.4�r�A�by4�	\�Vx]��R�;p�:9=�_���Uٌ�v�Bϒ�yו z����Y��`���yX�
U�R�"�D
h���e\��ԝ�_Z�E����Y
3㢦��u��MTT���{��]v�@��@�� (����X{��d6��à��s�-�X,��1u���pe~Ĳw�>DÙ����憎	���M�k%��W��`��"/ ^�tt��c�㌮ܽ�����G[��(�@�^��ǫ��2�ǖ}�#����/z�~I߰�n�wy#�7ۮ#�Q�V�0�}�AV�ǆ[�/3�$��S=@g�)���qn�5,�A��J�	�L-tcϯ���]�3[�r�����o��l�2K��T����ƹ���F��
����`�����	4ÐT�7$6��~~�'����wj3�۶uRX[j'��{k�;Ɩe-�:}X h�H�&��s�UnV�v26���׊'XF���Q`�����S��l^I�42J8��NU��Lh��{0�h.�aŮ=�]v%[0u>:0f�.M�{=YW=堓1����6o����>:�i���ŵe��S���Iv�o�E���$7P�wY|�,��lΧk�e�����2�B���QN�k���!`�7���Q�h���4����06We���k��E�	ǍϕV9O����fǻ�]+��km��9������|�{L���������C�z�][�F���B�{��]��H�����6��[ҟ�;	K*h��
F���`.���ԠduMC3].�Cb��U.��H���w�oь>�����U'�����)�F���1��8�6ah4Jg��SGLs�:���0a���d,
�ln�c��.��1�혆efIf�,�GtT��jL֣$#��0N��SY�*�}�kߝ[�rt>���;~��a��Oh����<�F�.{���;5[�L[L���:6�mz_	㘷d>-��f�*(y!�DeZ~��h�#77���xQ����!����C����}+��a��L��^X�&��r�ϧk��\�������Q`�5"�
�8f�i`�3LH���h����ܿY�A�XX���39�c{V���ZU�ב�Z}�	�6v�kSWg�����k��������^�~��n��z�p3��4n� �b�h_��S0�cW�`�'��Y���^����CS_���K�:�U�Yki�u,�BmYU�1��\����5O�T��Mcj�`H�A�$z��3*��;��^�:�p]3(a����**�(��[㟲O�Ϳ��.��N��'�S�ni�Q���a1�p��8��6g&f����vX�<9��`�2�=٦�nGuE��,/�j����>�\,	��Tv}
Uú�M
k*�5�1���O^>��D�hh���v�w�5�l�K���j�ܼoinz�����$�՛z����U��p|����3��k�)�1�h6mFP���v�wDn���e�+2{]��gޯ�!����A����_J~�ͥ.�rpL3���]�q�?���-����rN���\=�0ǪPsO����|��`�Jn�r�J�^�s���im�y�<eh�;3�6j���pU��4,v@�J��5B�V�r9�<�wie-��io1y��mW���|�s���3��S��1G#� vTꖋ�v^
[�%���k%V<�w�����⡎���orL�A��X
�1��9!�ԏiV�,�������琞#��/��d0E��Ծ>=
�tP��ecӑ������ctZ�ڒ����Y��(ݲ�0��DH0�&EE_�Qr���e���6�.�%l��a�nq�a��m�F�gm"��\n�n���ݔ��qc�.�Xd�b^�����f�=xU�kD�]�c}(J5f�(��:�E{+ V�ýҀT�����S-W`�9M�M����\={%�AO�_�E�(K�!hO�q����r�6��`N�b۟Dh=�7�ű�6t���3���$�%#��ˣ}z6�Z�2!��5�oX�1�n�͍�**��h�]Z�O7�y���\�"��H�҃eL��1����fU�v����$�|M����1��؍�X�N5�r��]���������c6 Ì�fލ�eGġ�;�&:�e|S2�\��'K�_
�1F3�׳`�+ҳ�ǘ�+`�7Ft�ب.D�K.�)�lu�U̒ƳY'#������Yx�Wr)W]�wىQy�p��I ���k(B+L���)D��G�r�[��!�+�-+T�Y�5�����4l��@*���Q�F`a�S*<ZJ�R�.0��L\�}���ik@pޕ93��8iT�Dn5��4e��qI��u�mx>�-�*�6���+$ü�E=t�Y���-�:����k����&8�dx!tgˋ��h�S/��k�@3(2��A�F��w,�x��z��vlW`Q�ؕ��F���jiVȩ7�ǸbG+k�:��ޙՂDZ��j�o[���$��J�J�[�l�κ]�ݜ�EĘ�C
��p��VP4P��0�E�tNU�U��t��d��>�f�����r�:A	�X�­��z��u<f� �3zyIZ�X���ؚwR��sUה�/nc1�ٙ]��B��r�i�zx7�ήWW	Ҹ@��s�,h��Y�u�lB*/1��`�2Θ-J�����S��'�]�����g�:N��W}wQ\�-�l���K��qZ�77@����T�_uu��/��kE��ۢ�*�r(�K�3��fU�K(�����V9-yخM,F�ٯGa��c�k���.Z�r��P��#(3Qv ����;7�ռI��.�ں9�3�:��t p�ʝV�J��:v�4�f�R.��7�(��^M o�]$.b՜nA2nL׺K��lܫz�$�赛ܗS5�+�s���y�U+�+(5�����Z��q9]�Z�=�������ʵ��e�U�\;��(]�K"��eCJ�=N�����o�j��%Kh�N�n�g��ܲL�Ǆ�A�5�cDR�n��W��K��]���m��|�@jsD��R�rl���:Kƺ.=2j�/��ͬϺ�.���1���9���n�3ת��X�>j^�)�a�r;��$�7�L������m*�P�V�����u�f-ۀ���
�&F-���qU۝N�ݱ7s:��_9rI$��n�y��Ϸ����������u��+��d�i+N���)��wI���=^G�N���آk�ט�[6�y�����o��J���F�Ph��wGkh����t{ݷ�����M�����֨|��ǖ�γm�_�������z]j�h��<G��AQQ��"��t�m���\M���uF�r]�����ǘ<��ݨ7`�d�{tv�!��h�e���TEӯc��X��ΣF�ƫW��WY�bu��â�(6�Z릞f�������>;WT%9���!�8�t�ړAN�)��:h�h���ES֊�O���h�7TZ��ZsEV���獂�u[n�#�;c;j;�N��661���`��7sG���*��%cTi�!)�6ՋUV��5jl�m�1W�����"��A�[j�b�Ef#&��:MP[D7c�(x͆�4lgF����������G�qV]uC�����y�-f�7�-��iX ����:��9Û3$�H���w��`N<������rf�[q>�;��N�6��a��JO��,�l�6�B���8(c�5�z������E�d�lWdxm?k����w^�E��TWt���ۥ��C��O��;��n�L�"��1V��
4$-�+;5�_�[**� �a咽�U���\�D�{�0Tu�z=�tV�!����ґ ���V8�,6ز�/zk%q���>�Yڼ^A�ރ5����/E�{�Ϭ{�kXV��c�qX�b������םws֨7�`�� P�qCy�IN���ߊ�sFn�Vz�c}�^�ݹ�oS@W=z�ì(F�O����]>[t��F)�ʓ-��h�"��f�.��?b�iS��M�jyF�p/˥k�d��3Ot�#u����(4bZ�-�4�����v1�M�~��lzLaC=�9|}ޖrlZ����+9;&�z��zu�(�τnK��Qb��۷c���l�P�b�5�Z0�6m���A#���,wvM���Kw��jG�j�� �E�+����E�0Vl4�37��s��=�8g5�ٕ�pQ閝'bu%A�F����+q.��Z=QJ�/s���L�����=EOo�-�X��hI���-B_�Z����=���;&`y0�@��li�:�Uٗ}�z���C�$��:�^[K�8�Z��.g�qb�v��f߁q�V�^0���W��uh@}RG���:��ۻ�N^T�=~�O��#{yH�ư,��4�	�,���]�جVz ӯ����3�r�v�,���YT��Y�*��'�
��^�ӧv����|��:�����Œ�8!u�[�F��
������)�ȥۦ7��P'��k�^[�	�9�,�m*����M�:�+�φT�=>+b�pA_]D�tǝU�-��� ��v��� w���QZ�ͼYz��K���`��xt�¶��s�y`V�=3�`��-Jk�b6b�r�:�U˅��4�3��ud���$�����Z�}��o�g�����g��"R���k�l���\���|��u�6�������wʍ��|j���}0'A)�~E�s�W4&v�aL3`�>ýNs�Vf�r�X���L����4�_f�e�$Y[��iŒ�y\��(��6ܥ��d���35\���M�w��z�`{ScwAʁk��6-����k�{���K��-�a�BU����:�\�6�(�](u��ϝ=�p걝Ó������̉�'�|B~��/ы��\.FF�)��h�;�X��t�� U���o���h����1=팞QF���މ�_�H݊i搅}�����g����.�^��k�,��O37|%oX�+��Cj[u��HMyϸ�n��/8S��㢐�\�N^�
�����K���zz�5�7%�:�7�m�>�ܭܡ�Q��Q���P��3�}�`�e�2m�m�����P�(r�����'/ա;:E�0�j���pi>����|��_l�/���z:�+��;��L��Ŀ!Gw�3��$�IU#�/��K|������=c���6�l������N|��:�f��]����ǒ�!s���JJ�u��+�3:X%P�����w�ҡ���S��J����j:O
�����kcn"���4j|�ǻ}]�(Қc��F]uT0v7��GD��ap��}��Z��24��v}�Ja΁kV-����/�3���ө=|Q�L����W��ލ�٧L���`�� _�(����)0������������K״=ݜ�A�z胑K}��{lNG�p�K㱱�B�O��p�{�
ǩ�`{n�f�m{�96z���؅�	�h���Y*��D���ᦾ����fk���"%(��J(��_bη��rH7�!��~ן[*��Щ碮^&�
�<���e����=�^�]DJ��z�k��m�����C^ˍ���_z�r��v]��D�+��;����}][x����%���FKY/��]��O����WZ���q���4R~�"��5:�a�|]���LW�5^���6��	�*�]y��H����\���A�qM��Wk�c����v��}�
H�{�54^�9E_Ok�}��z��lgu���8�c>�~�l�k���e�3���mXl��I�b7%_�=!�=�o[Lӗ���xX���JʂM��6�U�@j�v,z�=]n"W 5m��i�v�%�Fm�K��Ν�<� `����.Yw����̛	>MI|�|�;����_q�(b��#8`�2�8���a̦�f��y�%�f�(]�p6pmJy�v�~�~��E,졾m�u�����y����猠\����z���|Pg~N}9K��<���nPn��X)m��Kx����ّz��I(09�%Iw���}6�_@�_@]��x)n,�pn�Ľx5��ܼ3��7���{�b:S���p;��?@�RW֏g��s-�\�G*�9���٬眄H��'4�������o�p�rl(�j�b/���	��y
@�k�ȸf��U�sׁh�ATO�(�jߎ
$H�Ɍ*	�>'�o�X%{���:^���U4�岬u@�� �9���3�ek!��m]_k��k�r�?16S`�m�,�ጹ�==���S�q�Jc+k%z1��5�]n���=�~<���6)o�͙���+�;���]���n(�X��9CvE�IF�B�4b��V�j8����,wbq=و�hZq�������HL�����<�<B�d�k�׈�#fݍV�Y[1�TG��޻�Y��y��U��쫲�z�k �q�Q�٪��������LL�Kw�Đ㱩�Si��2���u}���2�w�W�xR��R�+CŪӵ>����Ȩ�V:�~a�F�W�l���<6�r6n*+ە��\�T�u�x{��~t�ϱv���$�	�<6��hY�1}�4��I>�ƚн�B�< ��}F��H�����{u�ٯ��
3=�Z�	�W3�"MX䠮(��1} ��6���M=�:ՔS�''k0�ȧ����jz��A�MW�h��y�|v�2��۬���#����[o%�]�������$�И��Yk<�k58�Z�7~���1C��S�����./��5r(��M��#���yGR7Ѵ��h�Ȫ����:{�$�����,�Z��[~=X+�Y!�>��m��ʥ��I/NU���})k�Q}�����6�X8�Z�1ꙺ��zO^rU'r�8w�Eg@�	@����Jh�.���xF�]�_��>����T[�g�'{�/<��{oX��aT:���	&{}�^6\���2����-
/"�v�-�7S�����-2��|��\�%R�"튬��)'�K��A��0U��,8�#�Φ���@�OF	{��u$س���'pxOVǫ�>� �#��k�~��h��4>٧���7�(����F��T&��z��ղi�����TkB��e�h�X���w��H5���þ�ٛ�yQ�6��\v.�XV�(��VK��|��cU}t��7��G���}F�����9�_n�>�,�ŀZ��[�Ւ��ц��S���ش��6���)�a�Z��ӏ�I�0�-kk�{��\��&�нљ4!P�/w^��qAv,�>C+^o���{�Z�a��լ_k�����PÕ��w�z�3�TB��V;�p���e�;�_ӯ�t��T���o����PX��G#��Rm�~�����[�i�����}��mQ�GT���ɹ��U���P���?k��y�N��*�)����!ސ����t+�f����ZX�ɽފ�+��6����yX�MǘQ8S���.0f���U(M��fZ�lj��{}���w��A\EK���k��y�c�%��m�q�ۥ��0H��ur�?AY�'�ѹ�s�u�u$�Q�=ϗcFc�Weo✪��vk��j�b�Nڵ1Ğlձ-[x�w+��;�(��)��a�l}��� �����*��k���3X�Y~o����?z\�]{�����'�S�3MIQAu�ܸ��TE��|^��21v<�r��d�>�WA��U����+u�]Vj�!��E(��B]c��`��b�����}�����e�H��K�͈�F{�ٕ��zj����tj�sV���X��I�m�R3�&�q8vf�`��^L�1/���;*?@�a�m.墌3z���h��Jud��7�vg�x�>*K|1�����bǃ[([��k��s�p�3��(�]D/G�����R�_N�h���k%zc aU_�C2���=���>����|�S�f����V8�Ia�$[�>['�7S�zVT>5����=��C:��O~��cߏW�6^a�z����ﵰw˯�z!�V�嚫�Onk��Gxr�*�@��{���WV�����
�Z�]��P���0ʃ�:Z&��j}fi� *�Q����՛����>�����x)C�J.�2��)3�M>����e�fу{������H��ګ]�Ƥ�L+�hn�${�E���H���P��I/��З˗�� ���&��l 5f�\�qĠ��R~�hX��Y^f�2��m�7R4�uaY�f���Zϩ�Ͻ�y���Hm�7G]]J�5����Fo.�+��%ϪJ�Um�o|)�'��d�z����	lm|��
�V�WK���������i#���j�l��t�ѹ*���.7ܺ�_C\`�d��!w�x�9u����D.�^rv��}�[�|g�#f��U���b��
׼�YȋP6@��_�A7�JVQ�[�^f��U͓��D%X��+�����������Π��5E�KqL���Y|�9]hR2��O��HdeK�[ê��K�L�^x^0���k��BDI�&��w�Gn3�y$� (�{�����X!W��1�$y�}u��2"3��!�2��Rٍ(B�K{dy���f�h./�Us�C�	LY~�ef\I����NA^�Y[���iv�"����r��F��I<kz�!ϪV�#DS��sF��e��Y�OQ�yAD��=]�E�*Ъ}r��()�L�GJ- �hX�ݺ�A��1ӆ�b��DH ���w�L� i�.�m���wYpb��V�f]q���Gڤ����wD�6���aRr=�էK�U�`�;y�q���ӿ>��m�5*K���P�Q�C��.�hJ�խ}Y�wC}�U��!m�,b��<�)^�M�߆W��8�Ըqx����G��~�!껝�F^_\sb��-��ʕ���^�O�.�3;�/�w�]dy;��Cu�C��Jw��Δ`�VZ����Ȗ�*���&r�����E�}��{y*�\Khh�[F�ޝ�5���������O��Is�o��7^���L�8W���%O/Ahͼ�����rz�x`�����>f�1-w��y�On��l������rd�vg�����P{�IC�C��qVM���4�'�V
)����Ǌ����}���̿`�5p�mIl�8��B��s]��/�i�1GA��;���]�#}[hq�쳦
ٿ��}���$>�-p�����B��8D��S�4ғK����L�(���N�L�G�C�;���hiڌ��ʉGV��A�ڄ�����v��Y�b_;�Mu��5���9�J�*P�����9��ov^KF��R(e��ִ�!��Zr5:���*�����>U���jw�-XN()c#]���-�T�Z��ͱ����l*�F�Y'keNW���e���UcC2�D�i��Ԧ<�;؁�w���^���ݒ��ǲ|Tt���`U7�s�3gwjKoP��ۡ�dt�u+bHƼ�Y�inl�3�s+����up-�`���3WD�&�J�T��uŜ�-�[�v��'��+��ݻ!}Y{b�}A�:7N��-�6AK�\�f5f�*R�0 Svm(U�+��K,�=�5�Ю����i6�I���ψ�T�GA+t�\�6��[X�ܦ��{�W�:ofT�O�Y�^�+����P�54�k-�Iãb��%]�:[[�;N��r��`Y7�]��$¹�>�d��V^�%��d���Ʌ齿��(��Z#�U�
:kX�KѼ1P8)o#[ ��� 6�un�y󽊭��V�{�N97��_fѭ�v�N6�uԨ�wLu�7�cK����2���y�C���p����,��F<[�
�C���r�dJF4�y���];[M'��Ѡ�3D�ͻ�"�th�i�,� �\3S1e�e+���T��(�q�]�@�+��OW)6��9^w)ٮ�l����eȵ)r�-c���ҵ."ʴ3���%�db��BM���D��O|���)���τGf�q����vWmv.A�"�ee;or��!�[W�݅*4��5}���lf��K�H��A�����-Xip#,&.�&��Y �݋��c� �(b�$R0�M0��Z:WA-k6��rDp#˭-l�[��A7H������Wԑ�ǁW��ج�]:	�wM}(�WQM��9e�Ӧ���"[��Ҋ�$��- FΙFWN���;�ɩ�.;b*L}2��E&dxm�Ɇ�[�r�[c�D�N|V򼕒MW�]��N�2X�9y����ec+��+�.9*u��rnW1�Zm��w���gf&��Y�^>�
��h��]i�.éi����{�D�q���k�,Yt�h+����Z�'5f⬏�;$�H�T�5qu[�hӂQLC����S��H�������G��>RT�i�8�<�@��ʽWؕj�$��N�m	�&�Xڼ�;/�����.��$�d�F&Rp��%�W]��a��·L��T�η��y�������-Wb��mک��)���E�g�/
�c������w��=�_C}"\�	XE���޹;Ei�՟_*t֠��{3)^�/�0gr�24�m��I�r��*�`�`\�%f�<��rHVm���P���6����mʄ:Vo���r�VF>ccsݵ/V��1I�9�T�c�����V��c�'7c��W\i�4N�9L!$�I$���=�ف���6]`ݱE_����U�Qh6��i�E����4���۵�l4P��5���AF�j�>'L�f�(�|�Ѭl�ŃI��E۶��X������m�T֬`*ص�8�֌[[T�t���7m�qyn�5Z�O���l�W��I��ы��F�U�U�t��"H����$��;j��KThkOs��e���#���v��"�6tZp[h"
-�Q�X⼷��h�Tkα���"N"�$ky���5Q��כE��=�t�m`"�:;Z�j4m����PSUi�{��>ƺ
��k��Z�8�FƘ�mDE&ڒ��4TT:-�{��j��X��V67X�`��Ӭ���DA���A����"&i��t��o �q&֭�hj�h�#SUT�cy��V-PU�ӊ٢ε���*���ETu��(��8�Ql�u���щ��1QA�["��w��V<�}[>��s0e��N��U��7fuN�Z��j�z�MYZ�	;6�>����,l�|��f�k�J�Ė�S� b�d���O�Q/�+�p�PB �ϲ���q���|��F���j�#��:�>����s�u�zM������g�	^�ڣ�>�X��=��6XP�`@��0���#w��گr�����[w݂�Œ����iee�mn��U���s�(��6s���8��,a�������c�M�׼]iSު���~m~�'����E��n��ǇE����-�߼���H�m��Sc��1+3���u=v�`j���a(�f���L�k}���Z�m�&Ǔ]��nM���h����3��d���S��kz�b���m�^�蛠k9E��=�xU�Mc~� �3��ud���j���Tt����C<a��<�ia�#��ڞ�KgpS��ōpmz=��6�_TQ��Q��ۃ��`�]��oT���
��+��Ň���j�}�;�gMy�ڲ*�����<�π�-̙h~hWi�l��1�a����u*\pR�e�V�f��¨4KgnK}k�����|��-N�:�\]��o���Q�F�3��u�VmN��ؙQf=���qSq�4_L0��PpfJ{�ig2�	��*����cWzA��'�6J�#���E5�l_�y���a<*ݸ�w�A�+�"��r�wIWrr���|�U�͊��~���ۊi搅(���7���뫱��)�wW�Dv����i�}=����v9M7��d{"�@��i��g9ԩ3՟0�3�����Q�W��������@�a����5�n�gޝ�aQ	65o���5��X[�/a�o��4��5�*����*������nש(=�Lh-UQ�9��0������ϧJv�[����|����ϒ���Wx�_Us�b�����5�����q�;�H�ؖ�z�8�~n	Y9s¶�y����Z$sF��r��p���h��0ϰ�+�X��s�=��r/ 6W�y�A��iw)0�#>�Sِ�؈����	��
ɾ�];���8]iҰ�c��\`�>+h�-��.(�\�C�n��,�;+���t����k*f_��~�L��S I^�͔�Ըs쵣J��%wFlm�6( �G%��FD�L3X���0�D�FQ�75 �c��˹r]ynӂ�]��BvFx�i�K��>�/�l��E╗�E;Au�aw�".!t��=�s
BK�W�{�;���N��	����b�Y*����s
9�`�g9FORi��������ε�47څX䐰ޡc����5����qM(��%LF���[`'���q[�E�{��_ϛ�m��G�{�u2f3orD�3ȭ����Vn'�kBu�N��(��8r��F��ŵ��;�H�Ozo�{�SG�d�z�OD�p�z��4F��]���\m����K�Cd�I��I��*V֋��񫗠e��� �������O�&`�jR�8/��o���{�ooR+#���dI�hX���n&y�Yn<Rɳ�FGK��A�=��0�n��rN�RtܣL�Ga�5�jY=�[j��HC�(7`@ޕo���n�x���{�`���N�a��{���ؼtbrlؔ	���YKl�x����c��3��:��_����F�-c��u��,��ZE[S��IV��D���mĩ�=�gZo\��r<­��̳�\Q�퉞�ي�Kpm+�γ��D%]�JBmf�x�ዐ�9���/t�xwy:)�D�\�8���y;e��^A�B�/*?�β��S2'��}�Q14sa��@�G�����ύ�x-��������`�*"���*�[:��ށ(q��q��&��o�gZB�Jn�����nim�q�J���NS�����X!���8ґ�ʩs1�؛��gD�e��\Ǔk3z���'�s׊4J�Q�HZ���7^�
7����Bƺ��ߖ���tu:^|
>�=s��Ҏ�V�3�v�U�����*ǲ��Q?�w4�{�y��[�B���!���	�Pw2X~��3sDyB*bz�#�k%X�8�T�u��U���e}͊�"d��]5r}if]���.� �j� ,�h𫮌y=h%����Fgb�s�K�坱�ދ�Ã��Lv���K]��w�=�����cǃ�.�T�}�z	'�5�U��6�$��C�S�>�����kv���mT}y��������t�\���xOQ���i�1�7a�l�٨Sk � +(b��O���/��=����é`�I��T�K�_u{i���^G�V�F�%��u�ri��Vܫ�
�ɑ�F��lN';HZe�0��(�Z����1NF��u,�Lʕ����X�\3!�R��F7�rN������`��,�|��a�i�	�y3i��Ki|�O�v�l��:��<Z���!
�X&�z��{j*�dL��]ue�H��n^��w��(6��s�+�;\�m���*��{�ݯM��<��^�VoWG_�ٿ��T������^��{���<(��,�C{��a��[J�5ڹz:�i��	#��YQ7ֵ��0�l�2ǒ�`I��}ư,�>[O@��㜍3�4�4а���gm�P=�!n��?QYn>���E�&�Vd��n6�3:�i�`��iE�$j|�z$�*��c�}�>���]{���*�`}8r�/�Z�)V^_�p�`�\�Xq<���.���--�!��}Rs_���"�GR"��S��V���a.]궶��_uf�Q逘O�
��O���R�Y��q��rN����jYh۴��>��i�P�(�3�_Nif)�9��R�aW3O�Q��e**Q�9>v/֭W[���ն-=k;\�K{D{RWp�����ֆ���n�2$ΞERh2~�X��Ϣ��;�$�ި�Pn�>�v��ɉ4�(L���+�ʭ�y����U���o�_Ũ��=��VJ�:�F�U7j�C��8_�E���}]�0IY[���v��>��[���ְ6�=���=V�惐d]Q	K��!�s�@�Av���a�7;>C��[�������$&tu�|�R�q�n=4�Gmh���m���!N����
���JT�xG�f���;�/ޡz���y�:�ײ�f��A?X�Cn)��HB��W[o2��Ԕv��(��o�4�rh9��=����y��lܗ|�
mKc���]'ݵ�'��i��=���4>�i�m�:��5_d�հ#p8SNɘO$�H�	�O&��C|�߇Xv��5��g��,2Oό���V�����
Qu�ss����`�:؁�R����'��J�3G�X�,�t���qs��ٯFXK��W(����޷�-u���9i��j���7�tE���WH�)�X��b��f�1}�u��o�٦N�`M�uh/%��6��o�_J#�S��f6����;�Ne:�Z;z>�g&����`r��2�F�]I��#�%/E���T~��}��U���%Z�n����{��TMU�'�\_p@��lj�md_w��@���X���,y)3�)Ÿ��hNwD��MDv^jG�v�tmv�pA��'����rߨâ�\g�\�]]-�`��C���#m�p��t�>���F�G=�d�;�u�O7�/���7ؽm'�,?;e�
��4f�Vk%_�<�(��Mnp��<���ں�/~���{�|7څ_ܒޡc�����{�:m���fqjc����2�G����s�����ϛ���Guh�Ֆ�F�P��Gj
���c�M�V�y$�w�B�������7=9�Ň�x�l���%�t�gr�.��3�˶G7j�oء��4R��"���J��r�֌�q���jf�����q��jV��y���=LC����Aޠ�F8��jY�n~��~J�E՘�_,yw����멗=~le>���H����#Ѭ�0��vQ@5t:����)F]�.+\W*�u�/3�Qt&�&�����C�ᮮ�g�yʠ�NV9����6��S����)G�˨˥Iŧ���'w,r��F>�b�-\#��gV�*�N�}-��)b����j{]�l��~�����|㳢_��hH��²��1XTW��[������G�9�1o$��7RP�x����-�2C�,#}hU��<�w��2�+���f��".��9x���7�?yi�V$�W�6B�@�Ȏ���FVwFj�s,��d�)�j��<x���Cˏ/Cs�`{�@}_Ie���[�׋CWG��%UOg�a;����/5����pxv� �	@���k�"�}6��������?sł[�ϡs��Ǣ�V�a`�X��8�~��n�L
�I��I;�fqf�z��,��mk��`�6=x�B�m^=���{E�r�`�CBu�o�~���GV�,�C�*��T�m���q<7�lZ΃j�2q椋Z/��-<5�X���ZnWmؽ�Z={��������x9k-K/�׻ �찈w�'q9k��~���n	��=��E���]��|P���i�#�N���lKS��kZ�2Z��he�%MŤ��v�/�������M�n�t�7EG�!-i8�Ͱ�K�U�$�����*��Ѯ��#.��x�S��f�_�h�ULj�u���w�ç�N𨾓�_C�\�3do�����G��Z�"����]�!�7^�s�RS�F�x�k����ĝ��҆��Uug�o�.a��^l���/TI�xu5]	�.��Q����}����>�u��ǋ���a�m�Z�Gs�z��W.�J�ɎO*8)�kD݅����dQb��>f��|�X�o���A����&��њ���[�S��r��� �agM6�J+:���N�z+��N�&{-�^'����ږ��qz�5�k�mn(Jua��n���44I�츽��l��Wtu�M���P��c�$��E��'h�oks[��U����]�=W�<�$J����ԮѶ*u���~�9�͒���ô4�TyZ�x��v.�Xw*�͖��p,�T�˔���9{f~w�{��[Y)0G�I����2 +1X������Խ�c(V~rN�|��2���4
u��h؋1tk^-kq�3;�������;�$�������;���w%$��9�uڈ��ouF�Dv�$��}A�nei��͌����Gj9���R��x>������_�M,�ɰ�G�������R\������KP��z�G{a�	�au^�s��Vj���<^�\3ۡY!vHeC��A
$pj������}��ihՑ����v�m۬k����iB��DvU�a,��C�o�h�7�`���EP�Y�&д�(�� w}l��}Y&Ǫ'�S�ѷ������Q�W����x�>f�����ǻ�U�M`o��=��}Y+���őY3��X�\`��`�W[�������E���+���m7��"$W9�(CQ�k3/e��f�sH�v�c���	Ҝ�}����S�����5*3e�eo�$o"2&���PD��4��Gz��Gp��z �\z��ٮ�Z�c�)��Z�kvIJjP�V�YY�Of���f�a׬M!�����G{�8��
[	::�]<�V�{]�b��KsV�+�"O׺�oE��,�r⫶{,�Ft��lɁ͛�G��c�*���2/�=�^8�{��w,��Z�Tlo_s�����QM��ϥ�Jg<�C
f-Ǝ��ɡ��Μ.��B~m�����;"�R}�V���Y@�%u ��8) ҩ�S���]u��4��ަ��hٳ�\|�mò��oQ˫�]�+���ȯ�t����ڸ�[B�P���'{8������[� -�UŔ�2��.��t��y����4�SXcr�U�β�t��VS�M�%q�r0�r�����e;DdU��c�v�ؕ�
��[���+ap��gk���Yx�5��X�9k��M:�XAd�m�m]Kf�79����gv
1���ҝs/�-����oc���o:=�4^z�����ʴ �%��R5�����$�Z;�ʄ�ʯ⨩�$��+���:ŕ�m�,��cwE6E�`5����+#�(q�e��Yp%ʍGFs�V������ �º|����;N�2�>P�ʖi�.}2wWp e���t.E�Bp����:x����a<2�ߧkܸV��u�@��.����U��˦$��'9�;Zh�ޑvd�H�֌��F�������!����8ڎ^m���'>u{���Շ�{fKR���@QP�J̒.����R��B�K�"z� �]�y!98n�ݮ$
],��-���ﶚ'+�ɔ��C�w� �)�tdO"q�I�-�:�,��׍�����)6���~�V�ᛕ����8L|Cb��7l�m�x�-4�5u���s1���8�N����$�Y�Fhe=���/{pZ6���0Ƃh6�n��*��Ł��=��ड़��:9pɽ�zTI�G.���A��w9�yQ+��D۵%�by/\m�n]�Z̫� E��iskR�]��U�����l�EB�ZCT`���ٳ�41]����+��M�BS� ��7Vf%)7L�0fX.��ʘgdMX��Eȱ�� &���/esY�ַ�T�A��\G1����e�8ŉw�7Ah�:*�Wj�Yg!u{�7|��g*)ʝ�t���{_;w�R�Z�� ��i����.�n,�Pfby8Uܝ9�l�w��w.;P����H�*K���
����yΆL�_^)�B{��[��n��uw�]9������ ���CR>���@�aS_�d�z�a�ӳ-J�bї��:D�3����3�?$��NW��tox*��!�oB�ci�Y���l��Rem��gq�i��%SF��&r�v,��YR��i'�X���,.�KNa$��lɁ4G��a����/&so��-؛��-�Ow���hfi�Y�y�)�q1C��-߬'}����B�^,}%�y**�A�M���O��r#.�ׅQὤ�T�t4^v���Y�2h�j�m@D��(!�g��>h�PN�n���(��j���56ѹQܠ�I$�8Ba�'SW��W�X�4E7��m�͢��(�5�ш����(��'�ED�j�>Z*4ૣTF�kUSLh֝Qvq�5TZ3c;�:j
��jj�i��QTM��U�b�j�����j���.�����CZ��QD�M�5��lQT4QA|[�j�4i(�v5�v3^ڊ��I�q���(m�]��U�b�≛X�*��-���]h�*�lt����M�k�4t{ɂ)��L�PW��5嘙�h���]h*�&�'mDEA�qN�'QG����m��cDI{��Mwc�tti3QWmkOZ�1M��b����#�^m36�tt�EQMLQRA.���LǞc��툻a�*���4mm�E[b��*�cTWX�`�m�Pm��@
�O�y ���ݓ]�vU�gP�uqL�B���L�m������zNL�v�J�r��\c�{+��i��η˹��'��sO4�����A�Σ4�y~��vg���{�~��Զ;M���c˭�9��q65}���/)���zf�6��#U�H�[d���)lu�]k�)�'�+���p:²��x|�f�������n�1��̨Q}{��)5�b�DZ����x^��k=���_����*ϛ%HǷrDmH�ժmlVn�'+-����@�G���8�WUs������y�����v���´R�w��gr����h���@#� U}#��`���5����}6$m{}ÍǷ�0 ���D�R��.��pA��p1? �m.�T�>ϳLy�^������4�!�"�������|1�`�_��b�udꋡU��&�kx����Z�;ϋ�
��4ep�f�j�B��l񠮷��C��,x7B��z(�b���+�!�!�1���ݪ�I��B��>�����Y�.]�m�Y�2��(�:�(QϮ�,�D��*�u��$S<e����V�>�U��5�#��z���}}\{^Be09���.�si:y�E�p��̅w۱u�R�5`Q^��Me�U���:�e���oQ�vq��tS5�뎸�4:���]n��y�:>=^|�Ey�n,�#yĽ��bf�Ɗݦ�Up+��{!����P�t�I~�ϫ�k�'wb�^�||��N��<�VW��	ލ��M�/T�N4R~HxU1��ͥ��&��Ufכ�X����X5Y�"���w�A��Ǒ���ْɓ�8-�o�+�wCm�����<��Y�{]��<�+�Lk��iǜ�!{q��a1����!�*=��0�N���f�kW��s5R}���_�G�]����(3}hҭ�9��m�s�Uw-�Wu�o��r��w6�ÌG;cZ��𞎯�l�7(`ݵ���-��h��
��TO	txV����_r�c��̀/SwR`��a�䲰ݗ�J�&#�@�F�g��0{w��;�E��h����Y�ށ?!Ơw.�8jg������{�-�}����rh����u�E�FĶշv�[ŉ=~Yg������PT���T$�>�/��r�b5ݨP�F���&��6�:+�s��6La�Iwj��L���R��M�\4��J� ;���	��;$��I^����7N�S�c�����
'4�83a��y�(�Nn��lB��n�ZÎm��^ͬ��[��6��ل:^�.'s�+o�vj�R�ƏA	�P�W�u&HM�t�64G�[+b�A�Sր�A�k*h�O�]O]�����]��jޭ��h$�T���:��V���fN��{p��.�ݸ��B_�`�1,*cUM�ï=��7��v�5�E�ID��D�`J�Z��ȸ��fns��	��!����Fi��}�,��՗���s/|�ؽ����W�1�e��va��D�FE ,q�i����½T<X{ŷAkx����L]�2b�N[RY�3G�포e8����e$�B�SY�E�����
��w���\�.7rr�ҳo�Țz��n����U�M���5o+}f
�q�U�4��u�2��Km�J\�К\V���Q!u4���-	o�z`���#��[�@gu��S-m�6��ژ��N��n���p�u����l�{�V��\X�tq�	7���Y��,wh�Fb�I{�0p��Z99���������W쓆�nK�����;�܉ؚ�*����v��*��+z����=�n��X'�,0�	 ��
c���,\A��-�&�Wj6@ԡk��,\�6��Pm�����2�:ʹ���J��]�I����v����&����wXZ�p-��-���.�\�n�]�"jD!��P�$.w�|��6��'qo�&�Vl���=:3o�&#�مD�x���
C���|��
�$y���Y��Cb�g/"�Z:임�f)!�������`4#�q�k�]�a��(����t;�#	���}���I���ʣFՃ�'	�<�����L��xj�U���?���o�[���m��8u�>���d��D�*�w-��F9]W&{��C)��Y���t�X��OX�Q_f�Ւ���魍͸���o������b��ƆHbW��_N�{z�%��Z�\���X�]W�Oj5����>}�ZJ41�繙W8gZ���qa`RW&,k�x^�/�>,���6���m̳C�p�ZqR?v�/[x@��:��~�/QJ��n��w޳�<�R5k���/�y����#�����}9��bΰ�䵬�@�h˝���ތd����9�,`{Z
��ּsx+�����^��>�{F�N{Mr������o%��`���гW��]~p���v j�M�l��cDL���6^|۷���]�|�]���N�J%����?IAb�x/z*nU�S�w8~b%��#�<M�f{Nܽ�"��j�5��;Ԫ�{L���������m�a��u�K�ļ�=��^Y;�Z}��g��{��ƇR�}D}���sYͺ�������ߓ�G�x�h�����;.�1�P=,3R�+v�Q�:]p5�����y���N��M���5v3Yu���
�H�G�8�a��w����p�yw�x�hu,���{y�=��K,z�d	��G�{��Bj͟mm�A���T|�vgH��:�/p�V�|#2K�07�E}�|�w�r����v���q�6�pmd9a��� uՈ4�2g'C���*G�V�qU���K�.<��ɺ��[/�����\k���0cۀu`��Υ�sPt����[W��A�����ϡ�����.��Z��3����UpmV�/��d�y�w����;�w}�����N�	�}o���@�^O��M�tˀ��zJ��#�GN�[-�e�
��34�b�������vz�Q[Y��uP��/��׼��jqH_͠B�zk5�7��SIJ��o�;��߽[.����T.�Z�w���/>l'-�K��F�:Nɯg���｣�"�D��\�_�ƅ��}�����Ok!�=��mH������yI���v�Ϣ�9C쫕~Q?0�D�qo���D�]J9�㓦�g���#pX{����#V��<�ĤO�h��k�Y��!3F�N�w�G������s;`.���ߔ�Y�m��QY�O����UM�J����z�Zy��]�ԹH�G�(ȱ�`����߷k�[LO۽��	��d{2N�΍��P�iT|*�.�#렺�U��Vx���/�Yv�C�QAT'�zXFż/D�ۍY��^��]�"p7N���}�+�c���Wl��[�*!]2�z�stX�f[hVST6�hS�$��*k�k�ozܼ��ZXq	�5�J��D%&�%��1���'��G
��o�z
��y� v��n��}w�
���0rr�RԾ3֍��#� d��_�C6�j�"��]	��xV��/��~$��ư6M�#èޏP�� ?T���7�"#�t\�M���Cf�^�zN�(���T��nu��'��8���Q;[�6^-�����&��Nx�y���˟��q�H��k!��5���j�D��f����16���S���%g˛A���ߊ�G�����
�$����{ٷ�5�x��˖y����aǸ4����%7��3cG+��VN����Ϧ�ȯ �T�,����HaOT6�����A��))�Ƿ^���rA�}��A.�tV�Y�X)�e����Ec�8V��<�U��)�-R�����������Eu��akV��c�q~���c�{v23;;,��]a^�X9h������n�f�5�����n�Wg�12�0hCiؽ3���^a�n�|A��Wh3����a,1I���[|��R��&  ���CU�7�R͑��,ϋ7�3wn>������F⮘�[�t���|�>����О�k��N�٦���yjj�t��iS���Ǫ�;7��o%:���ڝ��)�C�=P�ztw�]1��7��^,<��w?��gBj���j��uif�����m�͉c����Sb��!g���ʚ!a�$�Z�iV%-�$Eu�`;O#�7�ȠW��hz��n��+8�p��	q<#T�=�LD���3\�R�pl�F���2���������^vyy�(��rS��7���)�x��޾���B�o�pɘ�}b�0���v�
��P▊��>���N9k�9b��HsPo�����q�n��՘��*�LB���7�K�U�>��s�{>ļ���lr�Cmu�!�n��z��K�ƅ﷤�o��ɧ��ՠ���4����}�U9�n=�#�t�l �~���
�#�G���y���N��^o�D��
h۱u��%7�{'i�FOf^�nxH�@�Ո���g*�ԙ��V�3����n���H�;�̚�0��2e\����#�ʏT-�Y���[��`.`ީ�S�͛�θC뵽Ԛ;�I��̕o�<$K��fg�����^��k.����c��5Cj�yoX{���������j�0O�_����~6��>�UI��U�pD�L0Nx5�I��+��p���q<z��x��CN�xl_�áϢ��>0r���w��f��a�㌱i[f8���B��rs���o����5�?1`���{�L빿�p+�y;������J����Kn͜�V�e�aXKZ�N�	�	�o�F_s�ɦ�[YP�^�c#��C��t�k���Ξ�z�'����]���:��{F-Tlr�x����U����(�d[B�;ϭc��U��;�(+��S7���[m�n��]�|�^lm�%��Y�.��[�Mh]�p�*cM?1�Wڑ��[X�D�h��`��;���+}�_,�~���_����q��T#Fpn��m���+ ��a.g>Z����n2xTZ���h{VԄUͳ��&Zy�Dv�4d��^#7[�T�r�,mk���;osE�%�-��������ɪ��u���ƄQ%g�
�5��E�ݩ�ŧ5e�^��+��v��@ڽ�0J�{H�+e��uk
�M��E����`��q]3�����U�QQf��t{P��P=}di_�\�sm󣳇'�+�M]S�6h����2�nT�:a(5��5(r��g(�]��ԟC�6S��ձ:�d6GT����EB�ޏSj5,�F쾥طcn&刄�x�I���7�@q'r�M���=�!�8А��N2�9L���{��g��a��2?p,��H��;���G�ﯬ\�m���N��&VS���aԺ����!u�����y�hx�]�O�|��o�q�agt�2��D��}�i����O>tE}�9�FJ�i�4�1�2�a�H���Bv#G;�Y�ެ�]����*�␙�N�v���@Vr:�.B��B�b�����˿�hR�-�u���f�����N+���i_ge�i�U_�4�$��.{jǖʺ�E���������?�o���밟�
����E�����Ƞ���?��������rH �@" �����q  D� J   D�����������W��
����*� D��t�bUV%bEV!UbQV UbEV$UbW��bV UbEV$UbUV Ub  �EX�U�X��X�U�X�U�UX�U�X�U�X�U�w �EV$UbV$UbV%UbV UbV ��q(�,J((�_�o`�/����B�R*�3��;���������~O����������#�����w��������}�@'߯��>��>~�ox{�������W����EE~���Q_��`@?�>�p��?�?������QQ_��O�~S��N	>����W������_����d��� K � ��Ċ �!T �
 �( H��)" yߣ������*��)@�"7�a�������s����1���������φ�a��;���O�����|`��_⊊��a��k��������UEE~ਨ��̃�W�
�����#� *��9���3��'��g������x~	�����|EEE���/��_�**+�}~�6����O��߷���������;���`TTW���������~c��1���������}��O���>���**+�_F����$������~_O�}~�������|#<�Ǡ�������'�����������)�㒋�sH��8(���1$7�{꾳�"�P��b���#�;��� ֩;;�WZ��P$u�U��H��R�]�
�6�!V��̪��Wm"k*��T��GL���iv�ee��ZT-�v�ZWZ���l۰j3i�l�cr�V����]��k!]�3cS�ً�T ;v�CD�E����MM�&ڶ��,@c���,mY��4U.m�Vm�.�*�B�Ym�F�����LEP��ݶ-Ref�f�����d&��6uw:[n���m��mf�w]bt�t�����6�M�Z���  ��y_e�v���a[]κm/Sw��M��{v6�i��u�9-�N��
��ݶ���-v�y=7s�v��7k�����vm����`�M���Ûu-�������yz����wkY�Q��W��v�|   ��B�
=����C�W�>��B��(w��B>��{clm��bFE�л�p�(P�>�(P����}�m qת{ޝ:zҵ�+j�ݴ�����צ��֞oY�ZT���woN׺^����y��&��G�v�C{��2��   y}��MU���i۹��k̯oy�w����]�=��]:{��p�C�H���)�B�u�uݽ��u0=5����5��Ӡ�o^�u����oR��z�hdTk
��pηN���_    ���C_-�M���[M�[u7���P���ݵ�q�oo2ڹonj3Wo@o{��n�����mi��zhe�ۻ^v�o{������o{����){�\�A�:��d^n��۵��ة Vi��   s�֨ =����֪Y�qYV��\(�˃�*����5�	ӹ��k����eWl�*�i��hS��m��)�Lh҆&֤�m�  ��K�B��8���9�Ttⵢ�wUs���l�q KA;�u*��� �i��UG�ח� �j��lմ���4u�t�6��   O��>�!@igi��S���
������
���H�=��EWk:�4���]�K�]j��z� ���h3j�m�Vl��|   |  }pp ��*�� 㮻@V�0  6t����@7q�Ӡ um�� g.��4����.��m!���r��  u�  b`��;�  И� A��� L���[u����W���:  z�2F����x �.���!�m����*V�ٍ���  ��� ��Gz���#�z ���h �[���  r�� ��g� �V hPv��@�Oh�*Q� )�)IR�h0�Odɤ�*   "��Д�@  S���" � �J�ª@���?���?����K�7�.?��̟�Q�':3�����Q�N��h�/^�"��}���z������6�o�c��0l��`�1��C����0m������z��?���WE�m�fQQl��
8޳)�q�rh[%�Լ�nee<�aܺ9�جB�T��z�m��<� \;4��1ܱSR��b4f}��V�CL��YU��hY�Fr3l��+�̣p�2m��5L\�IY�_a+���l�̼��@y{A�n��U㒆S`HB�$�K/i�7$֞��DU�*Gt�v�4���[g�Uj��Ѯ��VQ��B�ƧF��ġk@�
�d��7�S}��FԶi��� \Sj6���M�M�v�6���u@F�1u��	����fj�	Ȳ�\%���h�&��{u �4��*f�V�Y�՗�/Lڱ/kR0��aV�S%�"6P�q���n P�w�N���E[.�Y�e�NfD�y*LL@*m^�`��PeVk�F�9OsY�n�(�K:�ð�F����n7m�m�%�l6.��[������ԍj�rݼy�'�����-�� e$I��Ui���U��^%�N8��Cv�`�ù�&PX�N-�JQ9�m�["܋p:�yY��!
,&�j��K����#!m��P2���KhTy�*5�̫k�x��17}���[;�bMʠ���b�+wm�麱VV�5�"mޘ*�{y���5(��.^�F��@R��*c{�WV� %(ѽ#4ܲڢ���e�5wp�#��eœ gp��f��T���J�,;�@S�1���Q��ې�x�2(�6��4�m�`���U���XT��xwF9A��FQde���ʺ62(^]��lS�r��[wx�^X�b#E]�\!B�!lKܬ*�V�X� �]�)H*��wD<c:�sD/F�	Z-R�.��)ZXk.����mdaQ��ZǰfLW�1���kNh
áT7F�l��b��d�PF�^;��$x�c�f�f�|�u�[���٭�������cYZ�nf�Ԭ��؛{��9�jyڼU!Ӊ�V�[.��Վė�;��~�7��Hn`�ԫB̋27YR�}��.�H�m�
���tf��c��vHӒ,Ucqe�*��(۬�R&n�<�&@�[��Y�]�N�F7�7��v�&�+wFe���kV�V'�-oZ�� �G������l�p+�Sː�l�Gv�f���*��9&`���GXi ��x[����`&�z��C\͆�S4�nͽ�nB�� $ඪY�+�V��8s�*mbi1ґ\�K)�w������GE���K�I��#VT�5{ ˇ/%��a�te�[�ac0��mX�k����`FĻK(�Gw"9C^hY$;R�QVjt�b ��kʶFI�����aL�ky�!kUH椷��-�0�^����A�A۴�� �2J�*����uf���Hm<ؕ�U#���pհ	���e��6ӛ�g1Uv:Kh�% ��ԛ��`����U�E�������D�GP�'4�QF�8[y�B�i����
�<��6���.�i�6��VQ6:�� hn�`��5G7�6UE,���7V��������Hf�z�sB�U�Ål����X�h�7��6� +զ:��ӳPY���e�&AN-ef憋��qj��1���4�"X���k��vʱ��#K+U<6� �7	��o2`U0F,���Q&�r��f'�F�`;l�=���Զc�t�pV����wt�C�;��ҡ�U�wt+vTKXX��A�q
��L�-�5m�V�jL8K�U%k6�هkTJ���$�3a`խ��q��Zxta�f<��ِ|�wZ��S�,1FnK�,��m�FXllz�#㐨D4���c����$yKQ:�^��U��Hv���U�̍�;��o&N�Jׇn�;XEX��b��tF��,kb��N���H;�1^d���"�{D	1�T�6
f�	ϣ�ߔ��:y6�Qvڎ%enJ(���[PR[b&.Q��K;Vh�B2T&�;x)����� ���M����)\� ��A�b�Fh��t�6��+2��V)-��hKcY�JRn�ʴi�QB>��#$�@P;y��{j^��Z�F��A���8^�{����$Tu�FF]m�E�MCRxZ��b� 7]��x	5��J�ð�,X{����S{�`��a�v����ٴ7m�Q�V�E���ˉ��n|U�W�e�N��kr����2��y`�vn��t�k�it�F����M:V0��*�Y(��×>ٱ�t�C�[ܺj���q���W���Fؖj#f-�jl20�K�Բ�**�aejɃ ��m�K�ͣۚ�:��l�j�1�ɹ�EZ��ǖ3&�����5ŵ���5�E�wab]�q(mաd�H����Z��,����R���M}M��>ӕ�(M���gaP�^^M�Y2��+H�v�$b�IZy|�k:-�Q�Xk��:�4���WZ��{�ҩ��X.6��aL8�=P-щ������[�@��4ҥ*e�"S�͡��A)���w{Jֹf� ʽ+f�[X�{Oo^�`m
��3Mn�Lʵ��2�ū����*�JWlC�VU��b��!�e���Wbb$өH6�n�h��%����r�ВDk�*X�h��K���W�W�nèݙ�2J�D�Y-	^e�i�l�{B[�J��`Z�r�ѷ�'�z֢��;���N5h�
1wU��ʔ
@l�L�.��vo��j���Ƶ��)��&EL�jn��l|���u��U1�K��^���-@�[�)�V�M�W{t+�3Ӕ�2��C�2SJ�����	,��R���]hd�h�ɹl���Lɫ1�a�N�pQz�j��X-�m����Z��I#�.1��ڦӓ/Yy���TI2�2�e��S9BRxlн�zE�N���TnAYPIQ�)�cyl^���/%�a��!swD[�u1mZ2���"�۴����:�Ħ-,�vm]�,�4k.^�`:�= ����v�FE
tO���Vډ�����d0��JKO4���ef�AA
Z]*Z��FV*�J�a�s
f�v�N���n��XŢL��#%��
�F)�DH�0�{rn�$B���N��Lo��ʄ�-��J[f\���(U�7�m����%��3r�6�-5�&�)��!��[�)��$�JIc�҃r�XI{�M�0�4��n�n��S\iG{2�����k�h^
�-m�D�5��E�n�ӳZڻMe#�7`�ER��fi��F���<��0j܏>�sfm����t3$�-�R$d��jX� �/2��D���ci:�g�n��3�:�	0e��M
��bҷL�Z�QC�,��Y*����T2�4�D�R��f<�t��n��nҭ�B)	���+)@�rJ�m�El&���ۼu��E��� ,�Q�c�jA`ˊ�F����Io*ʭ���"��yn����]�r�ʒ��YM�y[&d�Rf*��T)E+Rd]E�*��߭!E���S�&<�T�RJt�̭�ɸ��t�9���;z�=�"c��F�z	U�t�+
��U�#��c�n�[#`ڶ�J�JL�U4ѳ-�a����[Z X�e������	������W�YU�[�p���V�]*vr�ܴ�V¦���lwЈe���˱1ѽ��"D�o�I��N�-��d2b���g`6Ӷ��� ��`�e ��{�hVm1,���0�n��}ek�����Ԛ�z� �l)oVR�hBa{�j�O�9�l:X��ǩ�`���@��G��e"����Q}�5�kH�a���w ��u{Kp��oP���gW0Eg �󱉁k�;i�z�]'[�aK6M�p�!Ed�W�bc��	Z�l$�EڂlmfKv򵣙q�H���I���LL���$�퍺��j�����j�#6�E�&Qe;M]�l��^���R��MK�۫O��cu��嗯)�C,E8�n���R�N�݂5���F�뺔�Q�SYr�_"?�����ձB��Y��գ-��+mc��~'F�5Pe�ط�"B	�w������a�Ұ�j�D�ۂ:��]l
UWY�cr�9�	��kI�����BP8H7M���պLY�6��SU��,�ܛ��y�e�UdR7`|4jrR�w*�9b+
�����p�I7�xfv��Y���b)��ө�G٩�Q����6a[���YF֩���h�;����h�[�����^��)T%`�h�B��ݝx������X���TS��[��V��C.�j}�w��̈́���ޭ�ʻ����l7�M+ 9�%v(� ŵ �t㙂��K5e�����m�܆�5K���:*���,�1SC ��^�4'��˧�J��.�;�n����6�P�lm�8+f}�d��2��:ǸS�e@na��R�dVT1��z*��P=t $�Ck-ݚ��&���K!dV�v����*�v1U�̊=�A6f�r�25e)��� �Mh�aٹ��l�ߝ��dʶ&�2(�jѫ����R�b�2;����-+ņ��w��ܢ���P2*łFӭ��rm��$�R��h���X 9ĭ��)�Ȓ�S��9�[�T,�뫗�^jQP��`��N��ed@Х���\�x�~7�p|XoGRKt�+2��2�{A�&��Qb��!�rG��P5ZM��%n
e�i��s]eYH��Ct�P�{@��(RB���I)�u (Pk.���#�=N�TU
�<�� 
�e?�uCr�ҡ�R�,k��}e'�3M`;Fk�����ἫE#b�[�&J��j��͎�Ղ�F�yksr�*���Pӏ[�%n�b��2\n�YD�v��;��ء�7m��B�VvR��m�[Ba̸�a�9y��h;SFF�su�2hn��y��CmPُk"ŗ�j�8�@�ٻ��&�-���D6��� ]a��j^dU�%�^�%l׉f�i� �5R�@��D.�GVR�R�팭��J��ܫ��̬��Z��T�]����ɑ�rf�)�)P��s
9�Z�C >+�j��y֕�x��lf<dc�������W&Q{�b��1Z^���1�LgׁiE�LjmiC��b����ݳ+5�0�]醆jҼ�s犈�V�n�j��@*۠��{���3t�jn��H�i�[N��X�&�E�|En�hSj�k�r��k)3��4�U�h���52bP&w
�{�6a���q�l�H�S������5��[�.��*S�/.�ϷN/�7��nKQ9{7������g3d�sI��K�I��&��]���gkr�1�H)���3��+E�n*tT�ka�.Z�lc],��J�[��c�kZ���G&���R�eǫ!�^j8RM�n�7S@4^��j&�������ӕ�sQ���SU����K5����!��;�ooL���wm�ul��@fE���"
�kǷ��(kZ�'i�E�ܡoB�J�ʌ�b]��ZW7Z2�3���EZ&�GU��q#r�� ��,���-82���R�[;X)�B�U�0���35���^ʍ��uQ���#&I��Y�)F��B���l�2դk2���h�n���"�첯ic�����YBkD-�׸�
I	B�uV-'Nd�0�iZ�/p֨�[ݭ�ֻZ�T�V����A�2-y4�2���ش��Z��I]K�cr�ܕ{j����܆�9W�Qik3*5M�1sT��˨"�w���sj0� dن� [(g��T��H��{������@��5D�o�Y`�N�ȴ��>�U�;ヅ�{GE�q�V��mÚe��9+���,X�F:pI�aW�����Y�D¦�귻�ѡHE��+q�W�n���34�At[���h��9�YOT4�sJ�{W�JQY4�0�kf+�.��{�<��Y�m*:��ʨ���lк����r�ȝ9�0jǉ,T�;ʑ̫��"
�Va�GDn��|M�9d=z�e�A��7B�*:ܣ�KA<�%-C�v����1l�,LO��e�oP{"��f�i�2Z�"y��[���I]� h�S �@�+"XV^����#j��#��
Y�݄�C��߂�V��y��Iyp,�v2�F�K�x�*�4�C*{�����	�c�O�P�iXF�u5\9l�k,�rSX[�s ��tB��f�v-Z&[�{�Fg�F�E!@�c�ћ"	�u5����B7�EN�f5S7�`aU�eA���J��H���ݕ�-`�2�V���L�0D�gUM�K���w2���׭��a����8����6�����K2�7�aхP�EB5�5�c��sc���K�Em{4f�D@bkU�Y��UìfZN�e����Z�ID��D�V�ո�zjlyu ���T:&F�Y6`�5����ܬm��d�n�q�hSm���P��I�u��[��:�HPkK�(��k7�
M��ԑ-h�7�`�/I��'��h�z5��Q��J��N�I�p�*jtMmd�Ƌ�D�V��f&����+�6F�\ ���UH�6�y��U�v�ū%&-0��i]�gv����md���Cy�{�C�O�Zġ4�mjD�fUMCZZ�&R�6i��� �c�4�3��7d��#W D8����0n-����kr 싃i��˽�Zsd��n�T��'Γ�JV���a��/�-�;u5�N����v&��(I.$w.��ղ��R��%_�Tzr�� �Dh��`��ݵK�k+ۦ�bn�]V`�%Q2g�����l$��dP[E�q�05�ٸ���tՇ���n^�2�I S�����v/ +)h��^L��s/��Ee��Ԗ�înL���,�ׂ���[{m�D��	g��m�)�Ҿ1��coa�c�$�ܭ�b���^t�.�fD�Z����{�q�sG�C�}9�8�u��K��Vܧ�s�s�q��-d� �wXL5>�7F�`OtDRl�)�r�vul����9qA��e���u32�D����%L�xvn�W+��r�j��\T�r��ؑ9E1�@y0�5`<�	�yN�o�U��h�`d���v�.�V�U��֒�ܾ�0�[b�esH+�W`����XoM�hU�DX�}ܠTn�M�.�$���Jw%��Iњ4V��ӺE�n8Tː�$�V���Г8��GP�iLs)^��oRC�$�̡�|oY���34���BغF���_X�2���@���:x�m�3J�h<̕aYC�b>�� bś�:�$�f�Šj�Y������x�5��	���8ۛ0�t{x�m����0IQ�!�jw�\��Di���$��%L�,��x�t�!�g#�)�2
����.y��Y9k���L]2�Fͺ�5iw��Ox�f��MW[]ݵΤl�$�V��9���kk$��0XBdcݦ�WIд��c����\�����O�Gi'��ۭ�i��J����ׄ��{h��LKYjᤧ��*�v�B[�ǒ���3%��&��]��P:РȺ
�uAWy�Z�d�-Hob��|�e��Sb�֛=(�dkT�fM�]ogP#t?���Rn��y�k�U�������J�z��ǖ]'�m,�r��i4�j�0-z3dPQ,t� ޺k�l�٦'Ӥ�Ԛ/�T��-�wEڶ�iJ �{���ՊPCl݅��.W%=H�f�v�-Tu4U����;�E1��m`R̖��J;������N;���dǙ3�ӓ[��u+��/me�
��-Auv���骆�z�^[����`U��`�O�R\��ES�O`�ڢz��BL��EXW���ec����iڙ�ܸ�����,�u'�r�]&e8 7%���Q]��~8P���%��fڐ}���W:��E�U�޳VN	f�� ��OIR��J�;L{�]�C�����u��0�*Lש�cw(�u�#{%JRIh�K�t�+�yR���wyb�G]ZQ��&���fs.�*�0��J��ɳ(Ҋ
{�F��E�[K0�۫yUԁZt0vV����Q��t��`>n�v���,[�Ű���In����;�n�*7S�j�����z�X�D�W<d�zU䀽���J�;���[�CBU�I�]=oS���1WwFh�DSW����g])��	�ț�_Dq��Z�R��w�5И����\P���
�UN�����t�Յ����R�eշ{�T/z��Gg=�|ΑswV>u�d�I������w}�MQ��Ew.{ԝ�����q5;�O:.��|7��7(E����2='P�Η*��Yu�H�p^�]l*F��N�c	�2��ՃT�sWj����w�|������7x��5�����LR��0�o�2���o���y]�e�*�v��q��4�[yRc��9��t3��������siX������p#q��9$���9�6w%��h:̎�WU��G�;��>X\��gKS������JsnS��yx2u%O��}�%���)�C��G .P��e-}�}����bޕ�*ۑF����蕅u�'x����ũ�mG����soXr��w��6$0U��ӓ� �݉ÿ���ݕsr�����{	E�V�YD�+�I���;�϶v`C�K���&���Ω���'R��&����N�K�"��{����hJ�L> �(�Ǌ$8w�����ba��}���ѵ�\A��)�Π[�]����֩���J%k�h��M`8�7�[J�jUs�u)-*��COZ.��86�eܓ�h�Ffu�;:+�9�����\��,G�C���a�L��IĪ�tE.%�9�J���p3W��gA<[vN)�H�4uB�ŗZ���J�v�]C�P�Z+sh�5X��C� ȅ�c��������^7@��t��^���{�d���m��v��3�\�Om\\����H"%VHx�n�kz��p��Y/�E�_'����xh�wlL�4ɒ�hd���ɦ>t ��괤�&�:����gkuΠ���<�n���`i
��V�Ky�B��^g�L�Cg �+�M��x��ֻ[*��ҕt�s(3K%ֻ�n!7�U�x��Ryb�� zjݵwKfI%t��.��0;n�`� J���qZ-��g��v�Zb�(p����8��vǐ?������xڻN�ڋ���a!���ӧA�xh�|�K��<��u,�%�.ĥ��y��0Pz���!6�j�c�{U��]'+Kz��(<������IV0�I�Q_`�
Y-٨]A'Z�j�^c�7m�G;[ٺ�{4����N�Cv������Phb��Nm
o)^Օ�5]x��vG&D�u�Ȓ_NH��P� c+u��^��u�η0�;P=z&껨�)��N�Ñe��.ob�M�u-��\�/�D�6����ۨh0V�&�̊���3������laY.��)J��2�]�M ��z��P%|Ⱦ�����G�$�E���q�eh�]�������U�vf�����*­�I61_p���i�X�����%���BgR妋D'�1e���x�ܜ�t$��J73W
�[b�J�}%)K-h��ݹ�b��5i�2f}ֳp��*p$'e��qv�^t=}yOi'�hy�[Y����3�l�j����R��p]_[���d/H�w��+{t�/D�]MR�t��:�77��Ur8
�t�[�T�g����ȸ[��ώPˡ
Yde"��X���t�Mn��p�H�V�� ����6�s	����	�M�vFh�Ho̅�]�r��]
�&+��}��3-��\�n���U֩��άR�CS���N�d:�����i��m����@�EE�0*6�a����;�FM�A�(�8�ň&>��e�Ũ:cqO/��Y4�>�0�|�닰aѥ�Z�6�DՙB�6��݆�#n���\�n�9���X�
N�k��=���{�ѐ�k��i0d���W/��[9 Ѿ��^��4���nE�v;�ilo[�N���G�:� ����v��hS�뾈�n��|�&��^*���*붳9\�zT*]77>
+�gWu:.�!3v@D����r��\2�m��M�%�Zڕar���N3�f��_tu}��hG,��Yߴ�V��e臣���w����S�kÏQ`�u���7��|7��J�	^��]։H��Vj�B�/rCV޼DanX��0SYK��^�v�Q������O��u.�[˩i��Һ�k��c�x��ɣ~�q¹�:k���Eۆ�	�E�΋O]�|Mg�e�B[XfU�D:�v��2��$9��VT�K����Ϸ5� 	�y"�wف&R��K�T���w�tzn�}j�(Р�����D�m;�ɝ&F����ܰ,��d��c�@���<Xb��A�a9�������N>G+�ϑ�w%�*�u���}���B��}uE�],A��'�i�W���:�SO��B'R��l_wJ��}��^hw2��ܺ�Z�Y�'+o�iT�O���r����⸍�T�X�:�;�8 ܶ'[2���<g;�q�U(8�
F}}bYi����!���y�C|���.�Y]IU�vͻ�)��u���g#m��]�s26�*f[����ŊNz��T�/�vc���)��)4W���+����]OR��r�q��*��\a{Z[�)}e�Rw��YJm�o���VP'��/�v��GMڳ�.p��8r=y">�CJ�]d.[�q�	�ot���	�&evgHu�^�j�ؘ�Ӓ"<�N�N���G����{�`�������'@�ٲ���4�]�I�ǲ���8q'ⶱ�����\�v�qt �r��ؽ�8��T˩�=)��pa�I� �G��������j��.���Z Va�,aB��+��;z`��VbL}W���5.��@�;�c	�Z�*"�Qu�X��e
ŝ�����[�/��-�|���Ǳ�T�2Y2^��ynl@�nΩg�ͫ�oB.޼П	�ܻ/����Qc#�N]�4;�|*��+���H�Bf-��muG�9����lܫjSb��U�����]!�+Uѿ
Ÿ(e�k�}F����iv8�Y���\� �nR>�xT�������=t�d9�I!����m�B>}�"��l��_l®]D���"1<��R�xY;)\U�6.۝��-ϔ3�]Kuo'�jI�:fZ�yy�4�׊�@�n�e�reX�N�K�,�՚�W( �6]B��Frd���"_QsZ�mS�g�Y��릞z~Y�[Y4S 7W�l�"퓝�Ht��-�$�7�Oy�2�gR���;|"�o��]á��w��Z75u�j�t$�țX"�`�)d�U�'Q�o`)�i4�7f��Wa���[�A���YT7��b	^'S�.6�=��e����j�,c�fQ!gh��)F���b��V���5�#�4&����uiK��wn
h�J�j9��X�E�X�,�q�-��PJL�-a5 ��d�북��è�R��ɽ�􊓮.y�hb{tݎ�m�ys�?�*��Q}���%:���gNG\�T9B�Q����9f����K��ᶁʄޓ:�T9vC6W+��\v�(��=J��Q����Q(�>�7�9L�ԺD3��Dof�T�t`\��S�18V�W&�!��j�̓A]��2[3�������R�m*����;�	Iӣ�ҵ��JG��P�IG�X�;y����W΋����M�Љ��An�[j�_+Z�Wڠm�d�]���ⷷ�X���S�{ZAGl����%E� 9�N{sO|�+������ʼ�}�B�r�\�b�
�{F�m��/t�b�se(5��J�[w��\��y����-Eu{m��t�c�U��SHײ���6�|��'�6�#���(��剃�n��u���h_B"�qow=YS���?e�ܧlQMd����7�&��]9��y��FM�x3ݹ��Jm�NVK=�4v�r=�P�!��XZ��x%�
Wn4�R��ξ�\q*w2ou�S���t�8��:�?j8r��KWStf�˰з�VJ���;�DzQܺNT60�Q�*��R�f�������\��׼*�A�WڐJ0�i:h"kD��+��Q��s#�5�ρ�V�S�W$xur��WF��j� h�G%/���2�m��1-v����n�[w��L!�kj�*�����u�n�:EH,�ge@��関��,��/�4'�
��񋒫[V�VV��}����:���1pPO+%.�8���'���7�[��v�7JG�	5���M�^Aqc27�x܏��k�$Yh֪�ٙ������n�n��Rc)�UJ#c����O5@�!�F���ߦe<���v�C���o/,�r�
r�1�[��ǆ�`���*����?j'�,�(����)�T��8���"�0�;w}AC��5|�gV��B�Y����AGS3'u��^��+C���� �5e�'Q:�Mp�0U�[��ݧ���P�6gr��H 9�z6V-s�k�T��N)�p��K6�μ�+��L��j+"��.ͽ�*��2���}v;�W$n(iP"gs�Tu��w���� ��z(2�Á�T�%�@͛�_�MB_K�Mn��.,��,����u]\����J�7՗"��y�؆-ǔ8�UV��ER��@�у��#�����=�-_8�>�f�� GB�V՜��pRWl9ݒ�l�cz_��"̬M���N�[��p�ǉ���eCe,�n��˽�zg1FN=R/U�f�k}�����}ط_1&�ۋl�1�Bҳ�ޜ�+
,=�U�{|\�!�5�"Ǥ�NL]���ۧ�z�Z����.��Z/����v�\�ޒ�cHs���V�����#m \�t��ڝ6lԴ�n�e��{ >o8�i����t�E���8�&Joeoיv,.Uj��fpj����V�^�����S)�����q#*��K�N۫�l�������T��e�ݜ��P,%�q���r;;��E����N�ں!_�[�l��Χ6U�`5}"�N��d�Cz'*���C�k�B�x� �{�l.Ⱥ�MpƆ,����XVe"���r�hM�P[�nfc��Y����r�f�»�`�mLʓ���"���#4H[���@7�԰4tui��\�ե@�׹�����D��V��%4�o��ݏfu_RVnq��g�b�v����=Boģӹ�Mܸ�����-z�W'�&ռ��(�+�	խ��m��Ҧ��E��"�#ε��v!-B���9Hs���	�}�'e��ݚ���M�T�CCN��w�EL�Z���U�L6Uݚ�\�Π��WR!����"eb걢t�cL�d�w�k��߰�t��Ny�U��4W-�z��*/��d=��A`}e/��Mo��W�2�r���&�I��:������,=��@tf�hm�:0Dǜ�2θd�5��
�i-��r�9�*���lM�ۺ�h����l6�����Y
��� kk7��ɋ{�j�1��`�u�ڄw)�NSZ�9��Ď�F�&݇ ��B�ol<[撻�f�����c�J�G,�fMQ\ظa+*��j�E^�9ZO��+
ٕ���'o�d�0������Qے��:q��ܞ��2��z��6�E'�v��6?�`�1���Ǔ���������xy��q��f��\�ڶ�����閞��f�aAIR�8����
�
����.!�r��u���{�vj��"����jP����JT���ʺ�-(����Lq�Z�Χv�L B�i���NK�ח�s8��m�r�S�2ޮas�4�ѱ����������uv�X0����'0S�����̮#�1N�yQ����������H�`I�7��d�F��7f��"�|x_m��K8� :j���=���d�h�Y�Z�Lv����w���
�
�tWS.��p�)s�QVQ���?i��-.���p�M�6���*�|�W�HP	1�d�n���f%�7��RA����w��}��gR�p�,|U̢۩w�K\�3��r�j{V]r��ܥ��Y+%���
I��G.�Y(�T���u�d�t��SgU�G/�������n��a@l���Հ��Y�X�̮�|%�ϵ��%�#��,	��)��;j�;EX�b}�Ѥ �B�s)�d�*���l�mdE�����5d"#g*X��m�)��j���N%`ʬK���Y�N[X�w=ı�xw)��-��Zѷږ��y�)�Wb�hH
ܗ���Hŭ���Joڙm���w�[�@j����K��nٓM[��P�2,�:tWv-S�)���{,�h�ݰzc������"z�mm��Y�r��/��ȡ?_�9�@4�v,���K�Qi4�����`�Է�Z�n�q�ҫ˫ꎗ�9�ֻ�Y%g0����"�Zi�S6B�������{Q�Q��J���y�,t:h8T�l��(�O�[�ÁY�M���w���z9g������X�4����+W��--��cV^u��W��X8֩r��>��!�%�}�>��)�꽈9��U����V��E�0g��JԶƹ�z�|�*��2��/�PI��,��[VB�NVm���
��x��P��7id�T�\�ڏ�ܗ�!D��M���wzc�;J�{�h&,� ��z44��]Dx���4fU�U�0򫭦%ċy}J�Q�6�U�@�%N~���Q�'4�;�ů��o=F�AԝD���ffX�C�x�>���w���,bp���T��xY���Q��h���鉎�p��Ln��ȱ�l�P���t�nX9q����)��[�Z�l����1ԅ�^Z|����ґمEPS��}O�����7��b��:%C0"v�9y1��S��S���ծYMG��}��9�F�FL+�רBB'E
³8<�0�uf˒ف���4�SW���A��/��Yr9j�ZBx+Z�;�����1�&5`(͟$(bU�L�*�_��Ԟ�F	$�:��n��qù30�@]��HQ#6�5��)�)�\VSP��Z¢���rW,ݻ��B��N��v�k����N%V��ʲŕ��^�7)��1�]������X<���I2��V��
<,�7�*w[jM�\�����:X�`y�ut���Q�ӂ��̸����e��ƏLIx4e�g��lЖ6_�.�,)��d7u�+�*��ܥ�����J�t�Wa9����('���kXɃP��r���\X�6}��������ܤ���۫�A2�[k�������G|�.�^��<�J�6:���D���v���3ĳ���g����=�D����i�J�.i�i����_;���>��[�6���M��b�+%n ����b�P�S-�tęOʸ�V�R�w)���`6�T�v��GwUi����I���	�Y 4�dQ������1�X�7�Ҝ{ D��&KI1W�".�8[ޛ� 2ow��Zn�����t[����EQ�)���o����ںyZ.@tn��\���5I[0�"��Uv��xl�2@|a�s��k����*�'g-V�G���d1�c�+��ź(G3���A)�uB��ݢ�pǹR�ug��OT�wS�A�`�ݛA��-m* �gwӳu��M�%fJI�&�ƴ��L���E��M�{w��+���,W<A�n��<�+;��̵W��;����X�ͦ��4�a��O6Ľ���J�rX��o�5���N ���k2�w�\�6MՖm�b2[�fڒ5�
���J�M*��e㕰��v)Bu`=��pV�ЈP��Л�!�197&�F���$J
�V-�7[�
�mځ�Z���R��l�p��\�q�(��ݓ1�)����-��_^-6��]ܖ���ˣM&�L|orJmi6��0,G��ƻ1�G�p��|�W9�E��E�_Xy��F���%A3��u��͉����!#��ޘVh���{^�/�;
���J6�5�;�7�!|��,M���{�kH���jl7r�r�����P�m;z�S׷��Gm�PJ�	8�Z�RU��sSݫ}�H[]c"g\+ܗ&O�Z�^<V�)�ܔw���]l'-Xgz���)hM��(͎��`3+4jQv�x#��]�r��x��=c�qC��.����b��|~�)���M%7���˃'J�5V3@a�M��
�ɵf�;2��T2]r� ��@*Q���S��5��s�C:�k��z\9���c�g>#���+�T7 �MΧ�S0�E��й�h7�Y®��Μ�ص,�l���pw�uHn-�5�h��1����_֍�F�9;]em�N����{2�Zx>e^�38��w@w�����3Nh�u��RV2i�);ڰCb�gݑ���7�Y�D�'���E���G[,v�P�=�e¸P�r����.��"��a��`�LZG]a��_=��C���|�C3u]w$�a�!�y�
�������o@���g�@j�l;Ϋuݝ��P�u2!��
�=�V��b�$�W"!�{�3
�Y������t����s.��{A'MuC�i7��9�'dn��m��d%Pۂ��!^�r�[�R<�^��,*�q�8�qKq��S��Γ-5K6v��Nh�%LNv�Z�6�+6����m!{9�%[�s$��S����ݪcʏ�)�0i�[��JKR����Km��sY[j��N��h[+�S������R{��wʚ�ӧm��^�g*�Ŗ���oS�%��.N6��ŭQc&�Yv����Us��&�E%a=�w�W;6��u��L[�/i��a�[o�����7N'��[���i���ػ �*A�.��-Z�CP	cto�t����m�-���眢�Z�h���6�NUh@6.�����`��7�X�oU��p&����j�/�J�r"����)��n-�π����k�V��<��kU;����0�ONE��}����a'�>����q�7ٗ,�@̊�vr�O=|�)�x�����B�</	���V�J!�Pv����\�m�ٴ��B�R��m���s�Vn�d*9�뾧r$�� ���i�W5E�X�����������)����U+��Z0�ڄ|M�Lu�,��i�!�tx�O���^�3�_G׆Z��Sw��e^���<�}w$U�G���hc�+��[+7�L���bU+�Iۢ<
�C�6VS�S���m���V�Wr� y�NQ6v���S��;�Y%<J�l	u�8P
˒uwW:��+���;p��V.�-�Q��έ�IKx͜6�zm	�չ!��α�F�:!SN��u�q� ��@��1��6��.3���)-��2����`mj�$�4ӝwo.qLڱ��E8�f�M�ج�}m�FK�gP�]\$0�;���.��h�a�ޝz�6�,���T��u�6i���
�#��l���4����\]�8�U���=Cs�9��(j(Õ����ΐ���N�(��7dХ��=Lt2��u��\��Ī[����묬罔)F�S�R�]��/�ܷw�`򛛷��æwbT��)Lp����vQ�ڂJ��I�VG6�*��K��{jYV��2�e��d��m�札mr���J@ᬜ�솫�b�[ԦRw�n
* B�*�l�Ǐ�n�WTipі;�����,.�S"����y��qTS+���F��Am��zo1v�f�1�6m&Q޷�g\���_)����Ά�kM��9�����9:�W�����
����T"�:yzh)��O�d�A��ҭޣ���S�9�m7���[OP�/E0�v���Tf�+O�̕�:����Z��̅8��m������-��澡.��2kxn��zM�����c�t�̣*+�t��ɕ��M�8)�,��oFt��;�/�P���˩/s���4��C��90@�x�m:"��H.Sb�ʺ�}�|�RIJn�(�}�t���+w(3�j�����Op��cy����F��vZ�6�w=�1a\�n���x���YWs��m�c�١]���{�3�5�Sd�#����d��Q����,�DK�Y0��j�:G�Y����Z�oV��,�\̙��n�����Q.WZM�
�j;�2�!�5�=6�W0�*Cvլ#����+�Vy�ɽ��u"�dza�ɔ�gbⴸg%}اc�FI��V���4�hG�J���u����	���Y֠t�]ؓCc���;E�KUedץ���:���mv�X�F#ZuT�K�%�}�kXy�
X-�w����Tʹ���id�*������[���R�~Cz��R�2��ٰ���n>+E��i0y��q�R؀����V$�a����P�i�鷜��Ll�F N�Ь�0km͍�$by����{��P@̊I����� �j��Brp���e�˗w���}�E@�:�Rd��qc�\�|r�`�WV�MɽQ�|���s��n�Zws��=}�`���B�g)j��fk�M(��A�<��f2��r�r��32�B�D�%\�ұ���da��VX�f�8V���dS��m���$[\��.��I��k�]�w�>[qک�����r���Hk�J�֪5Ҋr5No��l�&�)�u��)ؕ�귊;jv�5���Ck��ʊ�F9fq˃9�=��Щx����1ST.�b����+�l��ҫw�� �Js6�.��F�|�R�m��X�x�ې�b�ҝ�&�ȸ�ьۼp��bז=��w������9��>�S1`��~�E�^%i��M"�R"�s��v��Pb��D��}��pue�/*�5ϸ��m�G>]&�*�N�ַٹ`�ZŻ��cmd�v9�� �[��˷5��j���ĕd��wإ�Gt�e�����Z��;�1��T�r=ѽ���Ģr�-���U�}u4�|G{)����,b�6{������􎵁�F;�ʼV�,�n����ry,�E��e���dJ�+b�-�#����=4D߶6/+!��j�d��ʃR]2��\�n%�V"^���N�r�p�	(�.���{�O�'��+���Tu���h<jJ0b�����у�',�k��Jp�V2K�x�0[�-z�x��=;G.�خ^T��y4�EJ�����7�B59P60�\ѲM9q/�
-�C%m�rd��"�5��eL�4����Ǥ�炱_<[fq�J�59��O�w��$7A"�UX��Rf��)���i�#ÈE�;{g}j:ո����<���9�Ou�wq_MNu�w���J�@
��W��#q�����@�]se0��[��8ri@�gD+ue��N����vj���[{�$RR�tɨ^&Q���y�Km����7������RwW9T��ta�GTmJ�v�'��EV$tK��*�S	O�eEV�2!I>�iVo� �8�Af��	]��cT����X�5x[�'QS+���v���*�3��/��0������tg2d�N�4���e������I���dbvuf+�&�N���N��4�R4���q���VuN5S.���@E ��'b�!�p�WR%�Rn��BQ)	Y�ms�����t�x0�C�����gr�ҕ�D`�t�pJx�Wf��G#�@�t��\qQ����M�a%Kt,��W[�u>��X1[��j]k-�;�t^˨����w��(�������-	0�(���2�+&ml`�sn�p�)Z��a��PT@�*.�����6��[�o��R�#z���������K�i��Rc�z�]�l��C�HP�k���%�%�t�ݑ�O9��n�_2�n�u���+ZM%�n�)ץν� �y[+�v�/CW,�߹՝��
8��w%V��2�S%۫������1�Y�P�9{HID��YW�� S�".l1XJ��n� ��*u�6
��
u��;�z�c-��S*3����&C���>�)^*V'iܧy�>�{~��\-�Y�b�n��V{:���C;�����ךf(�"����}���־�}��q��+AH'75>V%)A��3i�gweQޭw(f^��0+:1Æ�,*�NfP��qp���E�"����WNl(�k�6�� X+c�!HΗSڟ
�,�л�D	s�1jgE,\�>�3i�G0��,J�'w]������I��JC)�)p,���g��' :��`�o%Jɹ�� L{',aK��*Y|���ˉ,��I�����r�#%!j�w���\�3F���v.�|똚��h�nR�5�aŦN���B�5�}quq���1cH�-6�|3:e�p�kۑ��v�'�2t�EF�;��`C����J�T��΃d��4�H$�Ƴ�ỽ�)k�B�|�q�կ7Ю&N5�akv��qW�E鬩���A+�諭�����ﱼL�����&bz���%j��i�O�J%9�:��f��Doc;9�Ѕ��n�j�9�ܺ=dv��u˫��8�I_q���(��cU��5�k��|'+����&YMT�vhS�,�p��+��kȮҒ��vZ�=�:]�K}R�N�iu3ו٘ST�\�@�
�W7zz	D]i��Q�8��@]�I.�с�>�^F+�:��U�K�I��]��l��^^����K��XUk�p��y�v�7�_R�j;N�[6Y�2���8�˕a���n���R[
7B}�u4�v��$X��@�zAxI��>Թ����"
,�2m��)�Z�!��[u'��ʌ�*lw�����h��X���1qbv�j��M� ��ԕ.��y��}.�Y�[���{�N�+���t_v^Ԍ�Sč�[Ե5�U�ҕ�Y���1H�$!���r���w�愦qm,oKa����d���f��٘.�6�ܒ����u�ZYoU�1.�&n���)n���YRB�^�I��L;�[���7
�J�z8%�×S7�:
�Kop}�Tj�9�M�o��?'W��C�,%,2�rښa�{�i��R�꼮l�)}`�uM,;&��ή�2�S�yrF�$�n��×�� ������k<^���v�y�̧�;�:����\����nꢧ�����1m ���޽=��"|��)��E%M$=waD^�䰪�Z��%4�$T�D^��E.n�����qdwtvk��ۦPU�]3��q��
]���;�'C��멮�\���q���3
�^��/Y�hy���VK���ݹI �,�{�;3�99�d�d��0�wws	wq+�9�<�L�!;��C���u#-��z,%r��<��s��i˖�Q�������Y�GQ�����y^'��軸�nNk�DN�^�y&xn吇��NE纓�n�n����Ve�-�Z�Ұ�]��5ܓ�L�T���뇁�{�.��wq<\�z�nY9+���)/RU�!w=�	�9:���;�䚮{����y�C��\tf@�s��^f�z�{������Ng�kr\�Ku«,�����X��^�i��F;��]���꺇��Q�h�SY�Zb��=ʈ�@��3�}v�)v836���;cMj�r���/��Ɣ,"���c;��f]�s���Y
],��>.��c���G�ۢ��cq:q�m��i��,��?��V`�r��WQ�&#6�����n�/s)�zZ��:���q�V�������L��h����yHD{��mW
vj�*�V��N�&�y0�R>�z���Om߶a���{�o~�̖�W]z�G�Sv�����:��.1�u��i�A'�ևq��dK��V��X�T���WX�@(�~�8nd�{gʔ�m	nl�!k�&�Yމ��������fv!۸s���\��8+�uv�X+ש+�X�\G���$t�ھ-�ʜ�氻,T�����v���e��1et����Eɽ��0�W�Z`�ȁ_d�0���о�s)ws�K`K�T�������p�`�v��$�{n�B�ڷ��SVuO@�a��`}?Ld��:�\4'��`�o����h8u��ؕ�z{�|'z�ct�z�_���e�Ӑ-�M{eL��Squ@`��������kp�U��ӌ=��.��F��O_��B��O
Q�����KM��]u�S^� �����U��vGQ�H�2�Xt�Z�2oG�E��&��1z�2���r�OjK&��m.;�C�_s���pI���:ٱ�	L�˅Gw�����U��G����3�k	�)Z�z��+�e�8��M��������u��>�Ը�35���`�����}k�ćS��?c�Pr�2L�B�v�wsd
w�]���ĉ�`KUD��#�.vd�m_�^u9��2!������Y�}���
e����f�$����@�B<Z<�)ߑ��iNS�Z�=6\�7hȗ9(
P�rQJ8�]�Ǎ�]��z_� �ׅj��_�{���@��'}���6��^�[u���'�;`l��޵��c;�| ��Įk�N��|л����O��M���IQ���KflC;��)�]�x�g;3�����T��`��d���d�� d�\�1q>����Z[��ǳ��8:%��r�vL5+�v���y�~I�!�5��۪�6yZ3�=
����]�3�5��T���&"��NK�c�dwS��W;.r>*��=]����ö�������բ������&�F��M�Q_z���&��l�M| ܞu��֠Ω�^��iQ��~8��~�^�lM�?yܾ�0�ȿL�뎰YK�ODG�
���3^�3}aZ.���8�u�P�d�U�k�f0;$��E����<£l����˧]ڃ�,��w@�Qn�i�︄�'J��9��7�Q�yj� �J��
b$v�YӔ�>�ޗX*s6�rvY��ۮY�.F�
QY��������I�W�w�����ϵ��giz�B���Eįfs�S�n�y�c0z�F�<O�TO1��EQy,
#U�O����W�Q�S�z�&�*�X:����������N+2�}�s�Oɼ]�Ta���ho)j������#��"\��鰵�ϻ#��E��aX�k-竵�a��i5ސߵ5b�K��u�m����#��?s�Jq2�Zk!���srɺ��p"�;ʚ�w #�_�5�ȃU�]����59J����Ѝ�S��@��\�RVa>y�WV�G��^�.�(%|L�)��V�r+")��8[#����	�<��Zu�V��B&q�9��[5�!._y}0wN"�}���4�����׎Ė����\�c������o��>�~� u\�QU��tZ�6M �x����pa�L�% 7� �����r�m��À���8�& �9A�0=+�r|�(a��~��r��kl��w��`i7�����B��3�.�Լ�Fn�Yi్�G<W�5O �%�����oM��Ѻ�3$#��*{�^#���o�b�a�@�O5Y��'�����[gGt����t�4/hҭй,�ʆ�JJ�E�.����<&���-�$;0��Iq ���!�6cޙM�sQ��u��+-�ԥ"�CA<���7����W�Vjqn�#���¶j}J�-��4�~��Y�)�I�\�s*�����M�?6s����{bt�Q��4p�g)�	��N�F��0���zr"v���T�
�nl�;`����^�ʱ�wX��c&�i
���1�c|o�뮓��2�U���i��}݇�P�U}�W	6WId�ʛMS���|�\V�}�Λ>��i�b����;�q����?���Q��m�%�3d��V�2��7:�d'��Z>�
v�a�z�}d�aɯM݋�D��
B� w�m�4��w�s����#�"�q�$h���3r�P�D���s��zQ�3q ���:ciQ��;�[�3q�����u�g`V���m�o�Q�ԍ֤Ͼ�@W/�ۥQZ�.����M��9�؅�Cyӱ�*�}��W�9�;@��i�Q��i�Z�� �T2���#��b!Ȧ"�W����ɖ]B\�{#D���T�R�w�<fg���� ��T� 8ׅ`���U*�G�SiW��p�dK�7;�'� b��EɮYFXY����W־Y6���.��i�{�|u�&5�\�I%o���c��X���s��ɗ��v\mbHX���"��M���r	�cܝ{���Z���n�#���^}ب����`R�Q��Z�����'c���ıN�	��st&ؤ(��D2v)ؚ���H��9�qC��٤�FL?��#Y�<b���L���:��~�F���4��XZ��uLZWwm�n��P�C��<W{P�/>���nT�F� �@,�w�J�g�wqV.���8Y��b�@?Y4��αX�]�r�Y�Ծj�\�ꯜ���%ә�Q��jT���"��M����&g�$h]Ջ���ǝ�b5�Ҟ�)�O-�m^Xa.�`�zu�j�OZ�,U��]��{�8���G݄�[W7=�D�#�=�k���d�T��xZӒE�ֱ��,���Q�#Yw2�V�`������JY��,�ڳ�aV|'7W�ɼ�n;�4�XFqʛ{}�
�:��aw�fE��
b�Xϸ #o�
ZŝW7N5������2m�]�dM0@��jf��k\��;wa��7���v�q�n�u���GGD�h�7d��o�����������
�ʬ.�:�<�s�wm��Yw&�  X�������_��&a�"���h,��4��ȵұ��f=�ɻ4��yVb��߷n^���1�"s,[��<,2��N��(q����ք�㝺��|p�iD&c��:��v��܃�o�Nͭkr�t�m�W�-��9���Nv/Do�_������'�b��ɳc�\�F]�����1Rn���A��|�y��H4����r��;~Ϛ��u����~��gV�h�~��Z[�Jn���҉��]���9[��=�+�OO�_Χ�(#W 2����N��Sf��W�Ļ���������sV[�F�u,26#��{�S3H����@�D��0r��������f��$>g0�6g�r}i���?e�j/��y�(��K4�.)߀y��{�.�n��w��yX) /Vc�Īw��fL�Sk>ϥ�S���2�V)d��L��k"�|�D�W&I��*(�60�A��j5j������2�@+q(|����˴������0y8��އ�<�)�u4��<��!wc��=�N�ֽQ�B�,��é���9~��V%Z>��������69E^����A���>��)��rr=�>����v����Ԕ$v��F�m��W+A`X0����]� �P��Jb��\�X*V;�~���� �b��Z���1�^n���ک*7R�,���S���4s��
d�W���%��e/z�D��U�����,���-փ���AF+�ҧNE/k8Q)_4 3��u�ڒ5|ܼN�u�H����ި�q���Dbq�=]��D�3z�A����w�P��MW>�%އ��2Ϊ�<��,*�2㥵�Wx\gD�X��6GG"y��7�*��t0^�=&��]bb�~���o�t���:��1��;�+#��f�O�u�Ɉ�A� �|3�VH��n	�=#;�8�f�]Ü�s�V'|�/)P{ ���G"e=�L���h�g�{m��dʢ��t}��Z�TR��˙��/jF��4���Q=y���><ç���}3׽�E]m��ѩ�<O�TO1��TU���5^�{��7���1ke�h�ӹS:��@��0�|�>rr#�TfTzcS��L�Q\���)�]day��)�OB��¸�u�K;wS���>��ȗ2���H��݂/�� ��BGsE,Z.�RH�_fTː�2M�:m�
�T��'�~����2�_ɬ�tV1�ꌉʚ�Q�`+Q]
��P)\xx�F�Z�uˇ�}>��B�/.����O��C�4dB�Oe��q���9��U�����U�
�%|D�,-�/�7������V�ՠ�e^���@Њ�bŅ�X�Z���+�nl�q��� T�8�N":��(k�eI�Zk��~^����� ��Ѡv��J��t�*M�w��V�{��]1��;,j�v��Ƹ==�"{tV�+��;)���0��O97k�S�1�qqOzCŠ�H��5���	S���'1���\�ח��8���>�@A�5�wr�YX�����쬎��y�|e(+�2����{��+P=io����PBDI�5G�tU����4���.*n�@l��2xw�0)9��;�b�^�������mW�cp\�{m�/wT.����H�)pm�t��Z#P:'u/"�Zv,n�9⼙������U�/����c�i|�D}=a�;R�T���4��֮����w����9,��a#Y�3uVtK���F>U�?f]T�i�nv������w�4�)�t�sӓ���
�su�ssи|����F������mAYyK�ЧP�1�c|Fb��N_�ϋU���ĘNo������KG�MQ��sT�n�hcYq[��Λ��9pi����~.�QƖ��zEJ��-\&_?z���-7�j�*13�ga]�S�=�r�/�Z2���S��O�z�`�z�2�ld-���\g��v�)�f���e.b�*�F��lDwb�".��a�8\"r����ۜ���]y`耠Y�v0s�k@lD����\��;艅�+�����&��yL�^��CUե�tu���݌��r�t~��U6T;V_�g�WI��Z22;-R��ׁg��vr���V�%md@Vu��v���r�v����7)��d�{fep���*ŰW���>|;������n1C�1��6��,ˎ�Xd��2���nY��=B��#0D�t���F��ݗf�lD��µ�0���s��Ai�v�m�Z�ʙ�zs��>����9@�!��*>d)�촂ߑ̊c&���ܹ,(�)߳�v�8��K8�oq
8ԡ��ep�f��|��Q4�S2�����C�z�+Ewd�ZKz�H�W����UNhqd��ȪrH�
������?7bq�B�T��d���I9}y��[�:Q�8L��_����c��jRx؍8$7��6b᪁��B����^�]���ӰKiBh��_k�]	��6���?�#8�L��0��:��P�u��dٶG�Zu���i{�~LBn=��{d[1y����!�gZ���T��f��-[�M�;{�*��}ر�U^����p(q��!��=sL�ɢDkץ=U�Y��`�����V�]�k��k�]��@�����N����0��p���zݞa��ؾ�8&��1M�凾�"�r�nL���"q·;]���}'���-��o��/◊�^���î����2&!�Y����tT�+��v�j�k���L��+��W$���J��uAl��k{�F�}E��t�;���4�DǗ�1�{ut�Х~Z]֩�%���ϔg�z���JY����tG�_4t{��e�2i�b�rbl��$	��A�Y�B���N�vXNn�)�҆��8j
;��W���|[l�Q�-.��sԧ���@��Έ�ng��s2�v��C��;S��v ޑUi�}֪o$��# �q1Wd���T+���Å���W�{���_Ӑ��uP�$T��I{�J�-�{�����F�����~cI�]��#2��� ��?g�p��W�љ�p+����#�ڳ����κ�&_�³�5a��G��~f����1.<��q].ܯ��h-0�5��T����p���w�N��dV�mMh�I��^��`���^�Ļ��T���W��m��؎K԰�߸|���g!N@��"	Ww��ݧZ����I����p߾���B�.���U������!�����*��.�ns��C��R��,���S�fd$���
:�{�s���3��3�Sk>ȗ�N{S�@����Ӟ�k���(�v�9�q�;Ko��v����f%o��(T������T��-�n^сV+���*ao]��q3P[8J_�� =���u3i�j�ͺb�ͽ}���[ۡ�Y�q�p[� �����|���A�*%qb�����	�g5P������f������HI�}�W�����4=8��N����;&�S%��\a����gQ�O�-C�t3���R��˪2S��b�`W�*��
��B����q*!Ov���k:k�܉X����������P�9�*��"������79Sk��7�N�,���ĜHi�'��ҫ�h������,��0�p���MΤ��7ϵ�F����.� Λ��H�	���kF�T�.-msN�A"ȫK2�krE[h`{�v���If�NPP}�Ӭ�Vu�o,&�ޓ�c2��W����5yKVL�ki�`�
�'�
��V�`F��뇃8e-��7Mb]���]�̂���\� ���"��:`�-jװ"#���x���n�e�9�ֺ�(N�V�`���Y��Q]�ޓvi�^�����9V7���1��rua��Q����.�-n �eh�iEpw���0>D�D]��f;���
��td�fg�-OX�e���_}�gk�ip�4�,��6u�6j����e�hQ3*������򛝡�a�\c\U.�Z��3Q���VJ���}��(J�K�6΢G0I�j����&�q�����V�1le�w�##Җ�3��nZfM�[��*�N�'K)��\s�u�$v�zT{������,����?��m#|�hn�7:�iY5�ţ�`'�9,�,gnӕ�B]t35]&VP�C���
�:��^�,���w���N��&�'�{D*���+���lܩ�rܴVl;�]sZ�dr��9	��&��r�D�,��4�ˑ��l:v%e���y��Z��f�/�.Z�A�4�m����*���QrA9��;ݨ(Hm��df.ȹ}�uH��ը�@���h꽈p�R�}w�Qt�Ø�F�Z0�V�̕����N�CkZ�[C�YlىE���}�K�l��ϔ�V�N�48�:���ț��2B�ɋ8I��F'V_k�=�Z[X�*�]15Sk9�D'�qH�!<Kk^^��*V"μ�ni�n������:ؾr�u����LAo��Đe:b�I�@%B ���5�Yb�t��<��Tԛ�_��:�X��î�]h`�N�(�
;�;��N+���(���E�COkr����w�ʥ�I�p6���*ڷ�������GPԯ�6^P�a_1LT���K--��twUl2|����D�ҁB��թ�km��X�s�n<���Y�n�Z.��r���ЧL�$�wQ2��%��E�@�÷ \
�s�rW7�����eX��E���m�s@��y]Å�.��<��%G˅��YB{��J�焒�r=K�'=�ZQ�h���Z�Wws����u�+q�!����[L�[��r�F�$NUʹz�Ѩ+��!�jhV[�����G�{�gp��!ʓ¼N绡��G]J\uC�\����i
��C͸z��.f\���#��.��(V�C���!��A<�r'M=t���g���I��,�'+D�r�#,�Gu9���ᚑو�QN�PS��wK/�=���n�D��kN+�h���j���j�:������q�S�U�.�Y����<��H"r]��e$*���ȸy��.����犇��:T�E�y:B�j'Q+����l�NbaW,)=Т�.x��C��R�f��S��w4"(��MK��qL��G-]�\�u�<*@5��P�]yyW:u�X2k�sw��D�����4 X�t����j}"�'`��,�|�p�ɚ�G�ǲ�.��A18"��ۯ��쿫�;���raT�|�ȡ'�9���Q��_�y���ۓ��<G���~F�!�|��������ۃ�a�]�{����v�=��C���6��w�i#8������Y]z{�������1S3z/��ސ��ܝ���<;�ڭ����zC�i�y7XS}g.����7߰s�۷��N{��xOɼ�&��=pxw����]���zL*�ɧ��K��x�	���m�/S�wٝ#&>������e�������xw�k��7��yM�	ӵ�_`97�'>����7�9��|���<�p�s���~Nt�r��׎�����^`=51h�'*Ty��>���O�1
~����9���`��|w;������
�����������o�rs�۟_vߓˉğ���)��;|t�m�97;�|�&�;|O	?�܁�!Ǐ����0�維��n�#�����g�}h}�����=��o���M�Ϳ���l��oo8����'���>��Ǘ_�ra~���6QC�xC���ݷ������1�1H}U�P��~�3_`�B�v��ʳG^ �\�4��Gz�30'��!�0���=Q�]�� |O><|v�y���|��<?�9P���c�o�O�o}��bw�k���;~~'��N���yM���뿃��*�Sw�~���=}��Ws�̽�WgSU������	�3�<�����z���9�'�=��	�]�����90���x�'�nC����'{v���z����o�N��!����.7�$���o��7�9�׏~z����I��.� ��!U\8!��￾���]����w��r�{�o��<��5�7��xw�9܇�=��<&}C������yL*�;�?���oGx���7�99���@���Ğ�����Vu^^�>f�j��c�1��!�{���m��&��YL>������|��}v��!=,zw�{v�y�{C����r�y����ߐ��G��}M���<�|w������z|�Έ���B��<z{�M;JϺf~�f&b�������<щ�Z����';{����}�mߣ|w���ޓ
��k�z���a����U��oO������;_Ǯ7�<<��ʞ7[ro�O�-��=�h�Ȍ�����0�a�q)v�V�3�.��g�%�t4X�RcV3]x�N�w"�b+AVU�i���j�yф�(E1��U�:���Տ��{� QS45Y��N���!P����0�|�
�So%���zł���ip/�Mg��t�#�KsT^�.��;�~cǋo��������xv��9w�￼m�0������ߝ��|;�N��O����G�݃ÿ'��S���?!�0��޷Y|���8<.��y>?|�/���.���\��j����>��iޓ����n�� �C�x�^M������s�7��r|�����P8���S�o��;���o������=�ls⮼.2���^lx�x�d��󘊓
~(<�&����׸܇'?��:�?$�q��>?~|&�����8�o��=}��<��o^~�;㴁�/G���oΝ��;�|���?����>��j�D�����{خ�n�*c�?�7��|���7�ϟ�yw��]��PzO9��&�P(
(~O��ׇ낣O��o�nNC��4��o���v�]�������|C�a�w�Z�}����ǵ�(��}�L��?|'��*�S�}v�����S|B~;rw�ĚB|���ǔ��1;þ!�m�����=�s�i7�r���P���%}��G�}�����f�?:��]�^���?A_PX�>�+�n��*�W��߿x7�돨s���ݼA&_��ۿ���?�˿�����o	�!:O�;�bM���xpM�7�9�÷ }~��i����+�ަ&��-}���~�8��>��='8��p{�roi�9�����݃þ��܇�}��rraw�>}��˿;������Г}BO�~�<z��N'�}���'}w'��o��G�$O�����Նa�\\Y�n�F���_�wTn����W���]+��uUԺmy�:w�i��ݏ�_m��������o���o[���ψ��ɿwΜxw��������?'��C��~����������>��� �E*�Wl���	;�{Ӽ>�s�ۓ��=@s�u�~�濐�]�5��oHra�y�����]��w�=��}O)������{�I�!>ݽ��ǔ��}���ޓט��G���j|��.bǅ��]U����<T�o�U�<;㴛�'����L/��?z�˼;]�nw���\/�����������&��ɼ��?��<��I��{q�|�Ǥ�;۵����;x���'���Q;޿{G�US��tM�sn�ݧ��e���ݺ7�����c)<A�sa�g.U����
 
r��l�^�-_dј;�$�[|���}����]K�ڇ�,ѧ�9ft��!.�$ƞo!����}�m9Sn�U�`���/�&�A�$%��C�xէ.s�|�	�"f>�$�#'�#|��~���N�>�!8]���q�='�J�����rr�<��Q����I=��<&}~o{;ӿ?xU!���� }Z*���Uo�`�ި�<Q̙�#��}A����r�����D~I���ǌr~}���M�>��	�[|N���	���?='�;I����۝;ˏ[�xM������&��A
��k�xk�#�����n�_����_��;���O���1S�G�+*��?C���C��{��xWe<z����O�[}��˾��s�ۓ���N��m�����P��U>'��7�9ޡ��� �>��*��)�C�!�-���|6��Ç����~D��c�1v~����������|��۷��q��G�o���xC��˧i7���x˿;J�������9ߝ�����˿'����{|NL.������S��ra���������)v��uu�j�c��}X*����_/�����x@���8�Gx��nM�	�y�÷~��'�=��������~���.�����˅���|���S�y~���>��ʾb��+�*�}��m��_[�^�s��_v�Y醙}~Ɉ�E���=�&��?����q�ՎWol�0�����x~;y@�����<'��oχ/]�L+�������>وD����1��O�	����ļ�"�٪w<��D�w}1Q?|g�?l���Q�B�m�?~���M���?<���bw�q��������\rs�~����aWe���~�*ǝ����}��_!���U�����ȫ�ҧ�,��mo�Ւ_��*��� (�_|���Qɾ����������q�I>�{y������Sr��P�����0s�ۓ�X<�/�����<'��>���}�N��>�������*��r���-x�{�����g���}~3r~��o��0��z����r|C���w�<+�&��=���x1�L����ݷ�Iޝ�?A�;�ro	�����p/�
��|���W��{����b��G��'���7s�!T��}��c�Å��7����s��%}�M�>'!�?���o?#�!�v��?'&ۮސ��w�}C��;��\!8������ѽ'���<�]��_��|��}���X���,o먯�:C4^X-����Y]J>6��g�ӱ1����e����\��EM���v�f�$N�([]Ʊ��8�.XEչB��y��#z2�W����A>��cIW�ij�e�J����tۀl�׎�r�٭ӛ�;]��祐�
C�>�u���0��qG�𛐐<o߯��ü�O�6�S���ӿ���q�&�����~��r�������I�!}�I~�&��q�����waw�S����g����S�L��n�-�ژU�G��	�/�[��m�ߞMϴ<���}��#!Ʌ���{v�F��;�ͷ}��ܮ����(RO�޽���Ӽ;I�!>���yO?DL�#ϣ�=C�vG%[h��Q��>�!������ߋ�o��V�����(zM:v��������*7���A���������~M��S���~�>8����8���c»�i���{�,}�@��e_c}�<����
���e�����;���|m�ռ�roE���s�k� }�ro�N��|�c�.��!�P~}<�p�C��xM�99��<��p)�����t&��1;�z=�����B��1S��܏e�y��"����'�e�����1��~3��"�C�q�\��b���_`��_P�w�:�*|�Ug��<��I�����/}�Hra_v��I�7�$�}��o�o	��ɽ(R�~_
%���T}�q��Uf��_��;����-iK�	�fg艘�'��]G��>��1���ύ�7ǜs�''������?'8�|����=&v��Ǐ����?\�}��ɏ.��M����}�zOI��>[�=F�� }IS˵Ѽ�ϟǟ���}�ͥq^�#�;�)�����T��L��}B2��$����χ;I�;׏=��v���=k��9�����z?�q���[y������C�iӵ�~��ߟ.]��W���}���>����bw����/��v����Z�B��ߢ���1SD���c�ǔ���9޾�r�M?�?�90��C�P��� }I�z���ϫ{v�?��P����N=�������z��ǟ��!���'�������p�O��N�N��cw����Z�'�FL}�b��ٯձ}`����V�Sʪ
�鯨���Zj"��P���q���r�R�=T�Ż�������ɓ]�[`KΤ�{n`�y�Z�n[B]�$�h�+���j���;���������},Ц�������"��v��|攸�&�-4�:)�	sQZ͆�e�L}VZ莔��Ѹ�p9g"��N�^��հ��`����6u�n�[�
Jh"8nv�.�K�u]�X�1�� �{�dɰ+&��bY��6�L��)a9���o�����y��v��o�fܫ�)T`�z�nWzT��q�wǀ�3�]1��T.%�sW�c#~.��GO�t�9
r �M�"i�>Q;�&�-fx�Mr1S7,3�p����]��}F`��A\�!���8��a�s6qL�rl���u��1nn���Vr�*���
~����#��&#�ӫU�{�ʯ�O�i7�X�Rf׈�����uh{���d�|}��|�����}���K���}7�ے��zp�~>��v�Y�ޞ��Œ�lȗ9(j�)����0G(�/����>��*6�q���D�S��Tge�m#�J=���ˈ����t-7fC؉v�g��T
!�H���5�l�z0aG0�M������7���椑���#>)�|ڪ���Bn�K�{�6D`�B��<��IjNUO�7)]m.�6��Õ���I�!�5�r]�vC��������,-�ZV���\F��U9PNMFʺ�z6s���ԥ�U�˜��g\�5{.�-&VG�i燺��]ȇˊΛ-�u�t���`vJ�=���Wo�7�"�3��ǹl��`T��V�y�\��H��[8�ԩ��|�X%�5ڮ���˝-̴0&-�@ۢ]f��L�S7�|A�f�J�V9:�[���]0y�^�*��Q�I�x�>Pŏ�KG|7��a�F�������2��{�-X=�}.�~G�^�I�g�I���:$�D�켶�zMLWzf�@�H���̽�|����t�;78�o�l�r)�aFP�8���#d��̿�����yP�
�~}�UOvK�Q��O�j��,W\!�on��Ҵ襼,�g* ����0�a���O8�Fc�=����WL P3��n(�d���Y�� �5�f�έ���N�[.���s,-�6�y�g�/�pF��c.��ں��nT|�@�(Z����.��,������?g8v�w�e�h<׽<����{��ť�c\M˚! ��/���B�*�7�n����BK����c�y���n�XD2�tv7��zzc�3���{\�N���-an�ʼ���Oh�u{�1��wЊ4wv�)��s��;��$���ʏL�z��B\���~;��KsVg��B}%#Ij�F��������v���
��>�~� r�Ej|Yk����u�U��Vl��q��W+6g���SA����"�� &��[�L������#�����0�
�6(R������A�nk���}]i���,�Cjd��*b�N]2�Ɩ^]-8:Z�w;� }�7W{Y7co�+@�-��w�[ia�Q�qĦ)����Q�ϝ�c����p G\q�LA�3�	ꩦ�&l��E�]A�/^�O���в	�����C!��5u��w���Fn�Yi౟7Q��Qu��v�m/a�����E,�^'_�"�(y�����ӽj��.z�f|�'wsG!�P��iI�����5ڻ�qi6o��_ϰ�p�l�EVwG����=u�&z��[M6��&ItSX�i�&�s��Ç��ʯ:�p�C<�C��@����<�ރƬ꼽լn���E�~��}J̸�i��݇�D�Ϋa;���e�n[�g�o2z�׌��O=e����IN�۫y�l��Cc��0�nd»L06&�P�Mgċ��l�D�;"FT�γ��;'�����j�wvpt�*��GS���G
�1eRa��ym�4Dn�'���\L��f3�dЇ�$q�vG�R��*�K<�>]�F�]q���o�P�LX����/y����EJ�Z��}��T��*�MP��3�巯ʛ?vs�\��A��r�ө�� ��VuZ��a�)7)��3�'��C+�@s�E�yB�5%�]<S�Sx��vk�@�����L>� gg�?4�M�彁fJAh�ܖ�A�P�y9�|,���[���8EL��4J��O�4�`�=Bd�[�tc�so�o��Z��z���>۸�z������S4�Ӏ��A�����T��@38:[t�,�	RY�b�?�qXnނı����͉��]��E����������r���[=�a&�3�p��x���Y!�A
��᩠+=�C����U�)=���V�~�J(7��r�G�nm�+_Q��n8RaLl!EƣfN�x؍8$6��h@����u#�}�aU�������7>{j��P,��W{a
r���qʝ����X�6���ڟ>�A��Z�ؾ�Urրz��a*�X[?�X<��\�W*R�5�.I�m4��-�N�{��K_z�c�}>^=X ��Z8����G�U�טv��xbލ�s<���U'	��3OnMU�_N�2�ӧ=>�����-<p��	��KPC�����=��	e�q6E.SA��Tt�t�����ޙ���)C,���m���K��n��)��3Ǘiٷ����°�t���c>=�>ϕT>
S��'}�J�Ҵ/`|4R,XߥY^���]X�[�Os�<�|�Z"�Î���n� �N�q�:4�k}N�S��Xz���T]s"\�h�x�J��pgَv"w
%�R�Ӂ%���y�urKD�΃�Wuw,�^�����W�`���V�yE�@��n���� ����t�?|A6��T�l�J3��->&M\��O %y�ׅ_��4#�.�Tʽ�狽ɘ�#����c�S�Xo�#*�/�{Oq<9E��F�s_avX�۫�ѫ���<6�s��V7�rW���o�`s#Xn��+��8��/�>@wK
�E巾;P	'��(�ӹ�~z97�7G������-�.�q'G|Y\��k3�nM�.��&m�GP�QR�O2�OB�8|�nF���:T�Me���FB�N4�^4]�x<�u�I�7��;��9ja�B���b毒�AbX|���>�|�΀����ܥOw6	C=�%�%��y��>�ɜ�����A���\�!�]Os�A;R�����k�gO���/�MQ�R�6[�zD��7�E���
3�����[���LWn�w�����[)�d�����M1�zs���UK|���mV�d��9���Ԥg��.�B���$��h{�ʗǹ�S]M%�������d ��xѮ�J�W��zΚa|�JY�e.'YOge^��)h�����ҵ5�%�ée��w�`۠~eZ�����/�JxP3��|z��,�ce6������;U�q`e��Ӻ^�i4������$�� �40Q�޷�lOLlT���h��#��HV�~������떜�ک��s�7sB�+�"��y�>�<� �|l/��E?�q?/����H��3ֻ.Y�oK
F����� \�:�}�# ���j�V`Xi��/a�d�  <��6��8�q�"��8���N~3rw���쎶q����U��P��B5���/���`1�����zׇ2<B#�*��
��u�!��'�#;�KȎ���9[:�z&
Y���5��f|��z�߂ӽ{z�u�Q�e�8�]���c�T,E�^Ի���ة���GxVc����0W���^�m����ya���7U\�+����N�1ԉ`�}ɩĥei��8L�̿�/jw�����ՐZ�0�;yKK"��j��vs��۾�]Tr��ͮ3��;e�b!�z�̬��T�g�{�99�1ݐ��gVP�s�(��Ŭ���L����p˹�S�uN�I[wS��˥Ӑ~e����>�w���"��C@Ixʞm�K��B���ԩQ���7._N%9��?g8v�_�F��e֠-T�-��)�[E�#@Z����5�Z���W����O���.���-�_8/�f�3�]XeX���s��ؗ}�0K��8��R�Gr4^[Je8��i9�n���]�|���y�/�;K1	L8�����?v+.�ݬ��'�tD���E��dU�d�ڥwY�V��!l���x�\7J�Y�G B�̼����/T��d��m��ݪЦ2�1�RG0Be�Ȝ�b���hEB/���^b��D�*�9�X�.�R0�7�6��0�۟hO�7&*�K��{-�o��ն����#���OR8U�`��D��d��Vx���iVv8+`�qnw�]tD��s����$Y.j���1pd��u7)�V���[�M�.깢�eX�vu֪�j-̅�K����Q��)��i�����P�fc�F�ĵ�;�·X�v�!���8p�Qf!���6(�+�~��T�*�n��?um�:4��u���7C;��Z�So�n(H"��^��b���u���N�NU(w�b�J�z���LR��׸���58�1����\h�� {�����U]N}���(J���u�I�C�����b(�ʱ7�:�j�e�J][=�v�z	��e<��m!;d �F�w�75d=̊���@�)\�J����V5�^��PCo\:�*WBڃ��iU�]�L7�>����d�SIG�̐�f�pȭX� �H�v�/���q������51i1ĵW��,+�{�;f�:��V�r�]�yP�VRլ�c+��/����U�XwX�b:��:s}�ɷ{,p�CMm�Ak��;/nQ�k:
�:ro<J��G[�z�vf�I��W[-����`Hp�������i |�=y3�Vd����M����R�]'P�Qf�*�"uތpn�Ҧ���j�����H��>�dOm�jc5u93ZeQ�
>����M��^Û��ru1/&�|�aP��Ԣ�f�����LJ6�Q�ˆ-��J�g�V�Z�$�W���-3~����hiR���ڇ��k��rj�j�6�ӖpgZN�+^S�O��� 5��9C�Q�e�K�[u{*nG�YIζ	�_I���OY��\C'q�aZ��s��m�_)���4"���v�@fu�Y��� %��]q4N#�Z�&m��r�����0Λ
��ض����/2[cf�ĝq���Eܬ�@�d��Ss�5v��c���a�=��ѧH�໩3Jb�ˀa�ɭ��"8:{l�>Ckp'��] 1�j�x]�J�j��P��˒3�m�5�/�h�j;Kn�@:.N��Z���V�̠A�'�o�܌�"v�,�RY��g���'<+95�=�WzV$����+���f�*���J�i����xt|���vU1E�i�����[,�BV3�yN<�;��I'��OGn�DQ藒id���8��wO*A҄�=]���s�c��;�rr��.;�IY�8�TI��]��\��\�((� ���nC���E�䊺V��竸�QF��fJ�I�ʩB���BH�22V�"��R���\��9�z�DP�f &�Z�b�V�R+0#1U\'$�t$�QU�ͩi���Р�4r�<!$���YI뺁l�P�O�M��u�t��Ry���RuNEZ�I,D̋�d�qå<�wp���tr=�;���(�T��xb�y�������N���z���TJ=���A���W\/=t�*�M%R��K���#�$�!V�t�u��wt�R�f�EJҌ��s�Ԣ�OT1$Swr �r]+k"��^Q�԰4附��3*Z�10�(�-�"����&r%D��$�aU ���eEʲ�C�+3]��Q�sT)2�E�/I6DZ��gJ�4C��V_���؝�*A�d^`�nGO.��AJ�×���ȧp�XC8a�ֆ�cH�k�����0`/{[��ƅ�NI6�����}�|�}����Grg�~���
�"*`ɖ '�Jf��K��5P���qO-�7�3Z��]���''�eJ(�m�����Q~��Qd���T*g��=�|�pw_%���y$l�ܬ������T�{{d���A��$,�Grvd��&o|���]�����}FG�iߦs���>wL�rǪLD��c~1��i�lCC��lo��솫&P��~52X�&-�}Op�l�:v*��$\C�U���w]F�!�܅&:H�Q�c�3s��VLģVκ�<��k!fUT�,H��p8����xv��]��;�_���Yi఍Ps�����g0�"]K��ÛUo���^��i�:�_c��i�G#�zվ�uC��w�K5n�O��9��pG�@ĳ��6zl}9�a|��k���>���Dz��c�6�1u���䠓ݕS��z���'v�2!sc���ά/Ɛ_g��N&P��8s(�Q��K�[r�\����p.��l�.��Gvs/]Q�N�hg��\V���x��Q�W���������3*<�L���)�Y#v�r�>��K3>i%���P|3�ͥ��X��l�]3�G�u#A���W¦M
:��Dޠ9n���;�/��RT��E�N̽�K�W١�y��H�z����r�����Pu�n򎐛S�'�2_JB��W�}r�t�5��vX�JNDU�gE��х�s:�����;>Mg� �p�9c���+���2
�R�@��+�D�|o����Z��R�bʤÑ����z�i����Ϟ��GoDw>������]��wT
���G��n~C��!�����$t��³͞�5t7n�!����*
����_!W1��ăJr;.ͺ��/�چ��j�L&Mgna��������s+����D9x�$4���:`A�rZ��Ζ{��O,+�Q\}dw��Ȥ2Ǹ}p��b�b;5���͉�W(� ���iæ˘��[��]"{��p6�&�!�ד�m��+ S�B�	��ԨM�uhW1]f�2��却�Ue�F�L>�,+�bj)��zBaLB8��l�	�b�g��F�f�;4j��3{�cL��h��۶*nPJ��_+�z���\�W{a
r�2>⍹Sr���S�V�|������]W��~�� �q8�U���u��nZ�4��_�QC5�1���\
����M�	n���e�is�M��͠P��r��]׃��B��N��2ݣ�g�/)�G�ܗ���gx6�]��8ԥ���4����$�XQ^�ᶝ�d����pe��)O7%f����RD���#��5�}}����ҍyٝU=?�����0�Ng��q�2��1q@�ˈ_�(���Y�ao�t�.�Mt�+V,�;]�0��rګ����)�?%������>N#_�ev�г-<~�݂�fϘe�|�-z�?.ʈ���L:�b��o]��s��O�E\��b"N�7�"o`���]��~�����r�C��Y�T��M\�\M{��깂��WY�&/����-�j��}dR(����9s�n�TC��>������k�d�O '��xR��l�5\���R��!�޶8��K���Z|u_Twv�*�*�<5������ꡯ ~c�.�K�׋��
�l�ݪ9�*\v%�~��k�WZ��dk��}�E}`OL,�st-ݹ)�)���}N�v��s�s'�И�&��m��ve����T�FR pX���uJ��.��L�� ���5���K2�;|:~r�Ԃ�<�}���X�+��<9Xf�dc�"�@��k�3�A�squ@b��[9�N��/�Y���躝�X�����`J��Qnr�I =]F{h�׽c��P�{Bߙ�C��'h;6���9M\�-����>�by�m�}U��G^�Mڭ>׋���yr��$?����^�=�y��BJ�S�-)`�fll1��Pͽ�*�Y�K��}��0rz-�V3��a��e.��ﾪƧ�!>�ƷP��2B&d΀�jM+#�$>��|��������+�$8u�ae��On��͞�
~�u`� B��$�bj�.n:��]�Q���N̙�t�� �\�j���[�;����'�nwC�pQ�������%�?'��wC�N�y_Jվ��w����q��+{�{ OKmZ��@|���V̫WS;é$/��%����:�N��x�JX�9���?�WoRϜ�sB��J�иMޣֽ>Ib�).o��_�'�}����t�뉞/��P�>��{6��rX��"0���j��`�������L�i5�F;\5w�F��� 8��a���w[V�o˵��|�>�饕�6�S�T)<�!���`܋� Q.���G;����
�X�.���9U�tA�*����8���J^u\�-b�^h�=Ց"kƂ��r�,ᖕژ[�3�)��7F}�e@��E�Nf=�@r����]���t�g���Lˍ=p�>b��+b��cUs�7������⇀�@�1~��Ks�>E�Y�a��0M�.��I�:�4�5��$��tUE�P@F<]�o�nod��u }x��#���|/��lM���+��k�2��\�a�:��N��;,W^d��p(�u==���Ֆ��ڥI�3r_gH���CH�oS����_�����3�>�)9�w��>D�������ʕb��WV��d���:��]�����ˁ:����JV�p]��*!!�u;�S,0;�0�=Ϝ��Fc���sq:�T��M�Jr5}�:^: E|� t���t�-���N�F#��#>e����Zܖ�F���pvqIU�j.�~�A����1<�b9*�Q�c'"���W#Yg7��N��>!j�)�E��{��;���_N?��#�Y�>>ϔ�����l��&��6�#�ߣ�.)���`��O�3�цQ��۹�u�gg"�hG184ã#B�P�r��2����1�q ��b�2��-S|3���Ee7�fU�#S����M�}��x�"��ܺ3%'~�5J��2N��xO�c���"��1�\j"�)�q�G��n�� 땊,o�Oy�Stq�
�i�@]k13�c�C����I7����bÕ�0|�(]�����~Λ �D�����	�u�p:��x!����gy�����4k�`}/2;2��fc}{��X9��&�7��t�Pѽw3%��~6�_�%S�{���c_�s���=�K�����&�G����P �gN=B�ՠ���ӧJNûiK��ݚ�̕�^=�VڽRՋ=\�(967��b���_�k!ml��F\��ꯪ���n���:{g�ŏi��x�&j:�
������C�h�t�*z-GT9�R�î4_ӛ��9�|~3���_�9�Tr�zl|�u����Wm��~ey�}��fr�=S�?S����~s�j��/�+{<ǋ��V^4����)�D ��:߅^�������bu$�%�uo9�u1����Gvs/]Q���D5���s��>��u��^K�n�NN���KW� ��p߆�� ����,��Wi�T�ɬ�䋧��D������+���h�Ln2�3j�;t�^7�8!|ǹJ��^^��x�¤�������7e֭٬�_�UZE)E
9G�Gʧ�<9R�yF>k�b8;�Y��|�
U}�S&��m�2�Y�l69|�̳�@�"ʤ;L�OɌmNDv]�uv��K�L`S���L%Ig�۹���c�qP�r5��ʈ�W��f-�T�5p��^q��_R�5-m�Ě K���^���ëG��⧀�,F��s+��Bt»�_�,�sU�n�T�)M�L��X�k�گ�.��f��!�@�����r�P��dP�{;��z���=*����By��J�C�9�fm�5۰�?LŃ��b=��0��6��=���J�M���+3S�a��͋���S!5��Um�vf�Q���#��IJe�\��͵�� U��a����v3L����Hς�rxl'S1�؜��[�ՠ�����zȻB��H��x+�bBU��P�q��fN�Rx؉����V���}�iik�`��n�.�c�B��
���TP,��W{a
r������P���k�<8��8;�vX%`cA�����}--83!7��ȶb�� ���&k̝���Ɖ��z�}�'"Y���V�{���ی���	���X7����u�@X�E{|���ɚ�H7�z���1��?6�,dN�2��:s<����x>��Lm�7-�&t&��v%��
VKǋ	)��\jȠ����]����)��?g�B	�5H���ސ2����SC)�����@�t�"��p{}����R�W0C��4�(V{5�cޱ�o���.8Ճe��j
��B(:�7,�ai�2�ڙ�k���aؚ�4�ޓ�����`�}�L9+�v7ek�i��k�ƀ��uB���ێ��/�)VD���М:�=��,ɻ��a��dS���qw"� �o�(ѻ�8����zk՘Ҙ�y���h3}2�ge<�4�{�C����6�`�{v	>�rN-�X��_m����(ٔx���h���vDu��^V��I:�::�S�v�|V�7|�q�9^��>������S&��dϯ�:�<�qݶ9]}�:WM�m���k}�@t�rA뙫}�5m�KH�A�ι����?g�o&輧1��wf\��_���w2���.�v:�L�{������h8����4A��^��Hv�o���p؄�[�ج��I��Y��m&�vm+�k��Y�$�7_����rT!�S[�c �,>��zxvUUk�Wb���N�{��E�����F#��K�\�B׾F���;&s�����R�3��93���/��-'�޾�=[g�|�O���Q�L��E�$��̄�v%�������V�s��U��F�!;��v]���^u)���LJ~>�N�%�1	�C��d�e*��2�1��m��$2S��yEy{ OM�Mb���2%�Jڭ��X��f��$�I���/
/�RV�$o��J��<���K>ssB��tw��W��p`w7ȥPo�Ɩ�׷d��{��COƩշ�m��#H��
}�cj��[E�c!7s3�C�ڑӛ2�fV\	�6/e�@��o�R����I �XY����Xo���\sTԒ�6�4#Ɔ���`=G��,���b��7_�ή%�7P��M�GT��h*P읋!�����QK&�s�%�P�6 ����Ǡ���v�9����#�E�97X�VV��"� �@��9.��}siv�>�[z�z5^\��B5�\lmK��=7��ԔY;,_؋�Ml,�q���Ca�<���t�z5��kk1p�	xk�\kI�m.�f��NK�h�j�L-���v�MTo�]��eD�8E�7�_��=��sݱ�h�'��L��k�s�!Lr���#����_Tc˫�y K�T"p̺���[8a�ғd����ws�T�b(K���/jvT6b��Vf������ok*�cL�n���:��b��Ë2����GS���0���0�|�>rr��b�itͭ��j�|���K�1VP3�� �ʸ	`��o�p�Ѵ*w�ݵ������N�+�1��66،a�}INZ[k��sk�"pՊ.'�F#�����2gj|2w ��[y~V��[�_���%��'����e��C:+��鹃%x��N���Dkq�\��u���K�Ľ�5�]ǹ1(�d���>>�j�yϸ���;��:�3��ڎI^�Vu<���2��p���n����ŋ@@��Y��g_
ݤ�r������=DR���\�v�J��ř
�_E���	&3��2*C)>ΟB��"Ĭy�ZR�y�>릕չå�j]�'o͹tj<pM�y�s�J�-�޺Ӭ�7�����>�"��NGr�|��H�B�5���r+>�o ̫�F���$�"g+�v���J2�Z�B��N��qͤz�T��\�>��g�)��LƐcQ��S�������Ϛ��9-�)�QZV�n�ܿh�A���L�3���;ƨ�7I��
LdGu�q�Ȅ�Ö,�6�}L�-$/�ȭ.`w�����$q��U�}t5��>u��:��<M� �sJ��E9���V�	�΢J��Fz�i'�C	�N�V�����>۬�?aif�����k3ݸ�����yٟt�ż˜A̪�N�ԙc�m�.'�E]�a�i�Xܒ_ �ƻ�gq8E�e9�t�sӟN�Ӓ����R��w#�����b� 5��r��8��+�&�-�5Wz�9�	�1��i1�݇�|����e�o쾟w�Ż�Mݤ��a!t	<6E�Q?�u|��L���V�g��v�`lMΡٗ���ak-^��mL�!z}�P=�0�K�a/��~��E����r�
�0>��%�9��/����]����u�E+yDL-�����eeʂvrRoi*�=����{c���-��ijcV��]j�R��£7���C�VsZ�C>[NE^Q]7}~.�f�N�9`�77/�t$ͤ)8���_U��N��~�"e����v�2��灊ښ�����M�S�DN���g��G��%k�/b��T��t!���gh��0A%KW]]��[� �FjX�"��b˖�'O2��3���{�%��N�CѾ��%�](M�u��<���+�ƨZL��(�vs7�iO�v�h��Ц�1�l��QP-Qew�{r�I�_,��:�����۸��ޢ�L�`��v�uܬ��`�׉��:���Wb�ڨ���5sb7�}��L :�l٘���Z��nH�S]v�*uw��0K�����$;Mu�Woc�_v��pJ�̍��N�;r���E�I�R&�A"��[�7r��9�Ȑܑ��d����UX6p��2�c���B�)�9h��v�\S(+J
"��WD�ء��ն��
��J=�� �4�Yc4L5�9%xb��A����Z�.��&�mN��.��J7o��.<u)9(�+p���gW^aպ����R�)�70Sh�9&�����C��SEq�f���;:��q���t��ӽ�G,���9�|�M�+����a� �܆ �c׷{Ff|j�E��?.ϓ�3��֛��#�+���R�a�_s�ldԂ�SPs�Y��N�Xٕv,��&P��&���х��\�Sw��9�kF������Y�2�r]ڥ:�b)�Wl|�m��pc.�eM�#�m�z �����	ւ�u
�LGlWb��m��N؅�@n�.���+w&���';v�5l���q[�.�q��)-���!�볩,>\dž��U�bg�춟-M�@�ͭ�5��so�q�ֻ.���_t�أ	�%��D��K�V(��A��Ʋ�
y���kX�
��˒�t�Եb	܃[�v��8�,fB�G]�vL��T�Z�e�#r1�$@�4r,���)��q��I�;A�h��v���R�C���P��CIޭC�R^|��Q,�%G��N��.��Т(�:iz���/+�eVm���t�5o=�j�Α�[��h"�[��������u��ɬ���|��+���\(6���F��\��2�+6����?�R���D�'K�U�q^rĈ�{�D^�pU����b.�Mw��Mf���WP� ��.�\��V+@Ώm�q�guZ}j��aYy��}BM��%u�1	�8��/H�@N<�����X�&r�Yؼs#̟�z����^�i%.�J�L`4�r�{XS�Oj}���@�$�>\���\�*�����L���Mm��3�� ��HiP���a��������7Vp��ZMK��2�S	S���5H[��z��r]��\�vK��J���Q(�]A��w�MB��0J3��'P{HxU^g�3�(��du�Nyt�4C(NXi&�$�H�6�XR��Fp�2%CL�Gw
�D�s	͒a��"t�@�M�N��2�b�f��H��\���KS%0��<"�-H���)�!�VE��H������E�+V��	�+ݹzj��U�-��y��{HU
���v��`n�z
^l�V�⮕yEI��5$�F�Ґ�W/v�P�2.�a��Vh�����H�.��
�qG=��	t��g��Y�Z������^�IQ�UZ���Y��&�]dT����kC�q(����ETZV�E�������iJ2��#QGwpĲĤ�B6���h����4RZ�"J�a	�+ft�gJG]�VF��t4U2(�4fk,*-�)Y̐�%��f����ej�,�h&�UH�ez�t�#wWC�#Z�GPU+	�*�EB���9jHt���ŪD�":��BĹf�sWWV�Ϊ���[OpʋA9{{��fZ���5> ������3Zz��G2�YAJ\�	N���oDޜ�����=e'�興��Z]l�䬱�?|r�`Y#3�ie"ϹG��g.R�(��zn	`b�#m?��ۍ��'o�R~�����Bt�:�̳"Ȏ��C0D�,�}<0c�h��&�y�g9�F	���\E��E���'�0�o:y��8�������*���NP"�� ]\TWRh�ȵ�[��q�z�!�{O�A�ug�X|>�	[ѥԱ��V�͉�W'��ꗽQ ����'��U�O�f���B�p���ד�m��+>�# *�'��u3.IbL��X����֭wa"�E���!ElM<�w?���j��!E��ٓ�Rx؉X�ɱ��sg����M�,�}GUA]Ƌ���A�G|�����"�jbV�:��U�xx]?f����Ǩ�}���q��e��m`c`\Q����Ҙ����n7����l��D��1#I*01� �p��ϴ���eg5�.r%����l�K�3�b���@��r*WL�_[B�Q�;\�us��#*�����9P��z�L�����jx��k��O�;��?��]�F�O�h.?����Ҡxr^a����v��ʛc^z��d^|����|�%��e٧S��m��̜A�Ҙ�ԗ�a[PY�}C�۶aZ��*^0���r�s�s �pE,�ܾ/��+si�]"�[�f=����G������J�MOOe�3�>LX9֖�h7��=�)^����{������Q����x�Ӛ��7=���cY-P�]K�=qճ�XC֦�4J�)1�{|���L�dKrT�R��Z��&�H
����-(mA]c���������)Fj��{5�X��ai�E���Q�Rٵ.�ۆ=�i:zX��z5���:*�*�<�q��1�G��d]@�s��*�û3���g��[�=�_W�}��ӷ�N�{E�;���I�y9���'�a+�`�L�ƿ���X�e��d���c&���m���z<2}J��r����~=Z*J���guw^Y P)���K�3�\4q?_,�F]=��V漆�c�n{7�d��9�,����sJ�W
B=� 05*��p�ҘrWT!�S[�2���!�y0�<�`w�����#M����%o�`�����?�%�m�����0��$�����n_�^��F��5y}7��r��,�c�KvOH�* /~Y�� }�3}\���E,ahCXp-ރ>
CBV'oR��x�$U���Y�P�t����+��Hp�,X���W��oJ�z�}h��j�Q�&����(.��i�\!�赆@� ޕ��y$7�1]��� ��so�r���e�Pk����2Ռ���_}�Cg�I�[�����&v"�Y�KΤ��;�^��d�~>zBӡ%�i�|lkZ|�z_�l�٣ϲ����0͡{(��L�HR�%qV��őV!L2P�a���F{/G?B<=���<z0�$�9Q��ϒ�t-7fCؗnfzs�2g���^���i��1O�g(S�`}R$�$}���:oE�c�d#H���g������X;��x&[Orb��K��/,N]��#�{p)�x<ڠr]o���q��[z��� ��ԝ�����'c���ꂽ�~�"�ne�^ǃ+G0XU���jѮ��;�k�;_E� ����w<���|�*I=ٵ:��vT�o�*v���q�a�P��d�h���T��ܸ��Kn�6P��ھ���X�f��9�)�B�;,F5W=�~�~+��8���m�Z�936��wc�Ϩ�?�8��R������!T6:�WV��g�+���o]L�-�����L�6��^&1��T���Q��u;�Y 0���0�=Ϝ��!ҝ�/��u��+Y~��܆lh�aB�+bc���bc�VR�3>��W�mo�pPW��1�Wp�w�k�iu�x��vתѐGؙݍ�
���=\c`J�n�V#,1�W M)��ރ"G/R�*�,3��/�I�
�bE�P�_�������;�L,�nuԟ�����D�G�%��-�5Z�e���o�_���ly�N�d쓜0�$���}�\z�_e8?��������(xW��~3푮&���3�s�6MfvA�x{��s�jw`9�:��Q�׏�����?@�&��6��^��+�=L�A�G{.9�����t�R�ψ���=J�7o8�!���Z"j'�]3�\�3h���ǻ�fX�s7"Qj�L�VSyr�dwBw. �®ѯfu��V7���MI������s�h��,_�q��=����o���i	c&�GMMl:��-�\?q��u��J �. ���H���3n�=�Rc#�8�n»�V�
�*,�os�=̃*�1���J�8��$q��U�}p:��x!CðFB4�FqZ�d��qН�x]8՝��K(����I�y�g��W�BSpl��-������[s�'I/�����)J�,�j���3�8�̹�ʪ}����c�:��\O���m��s�^?��a���{��!��b*�nGo^��px�\��w�Z��,�⋼�D:�o��
�qSA�X�ƍLg$W�0QE=ï�� ��Ki_c�
5�۔�v9���rPn;��bt@�L]��;?*�iͪĜ�+��O興�>���Xx�V0}�otk�3��zck)�UNa������yՃ���=m
�b���|���~َ�2����ZT~��
����7�{~�G��N���}�R��N:�6-�W�xQ�w���r�"��|6WU�g�t|�QY�2a]��,��.;Q�XV��g�[�$����=W��B�f�o��]%�?�_k��g6�Z�����С���w���]��YL�-,�)útk��/Mf_9��`�!G(���O�xr�R�(�=G�+{g��:*��xv�U��U���;S'M��Y/��*
ΏHU�iw�VM����Fios����v��9�;��&��t�s��;��erw��(l�D�m�yFɌ��G��W�>�C�n;,����aE���	[ѿR�v��Z�͉�3Wr�FJG2^��/;Y�_[�`�S3΄��!�tp��ϗ^O�i���L%rtQ�7B;�:�@����۲�+��F��|9�m
@�ه����bxK�PR`ǎՍ�7O�졜�$��{��u�37_e���Ɛ;�{I9�`��qT��B�Af������zdng�cNQ	ZP�"oJODv�qRJ^b�Hv�8Z�t�橝�]����71.�K�V�j,M��S�Oy]��]�ԦFT*�g#Cpݺ��bn8Y��_W�W����
�%��Q�+��g�Z��s��:g����%}�ህH�1��xOZ�����f^y�=��ӳ�>Ժԙ�6 �@,�y�p�n�rɩ����F;L�V\��w��U�_�o�u�BB��w{��ĳu��j�eә�d� LYgnq��S ��)<WvtՇm��m��GAʇ=Y���.9=�;�j��E	�U�^�Ga�y��.Ѝf��}���s��B�.G����I�vx9I�D%Q��2aqO0�]L�5jv�+��qbXY:5��>��w7=���B��?z�~�zӨ��9x*����B����j�$Ɲ�u9A�j����t���LwPWJA֛�~��c��y�ּ$-}
��Y��i���n��/�n��c��;S��v�z��<(�UpT+�x������+�o�X�w��&��L�q��b�Zw����ӷ�Эw�� ����� �aZ��G��. S�MP��w2��2~��7�7E�9�N�˞������{��U�!��{����:'ɧkl�Yxr������(�g7���d:�N�]� os�Y{{��$HEӝ��iҶ�=HU�*ܙ��3y:�g6�;w|uqeK!��D8��g�7cxv�B�t}@֔��BU�Y]� ����'ʛ�W�=��G�&��9�-g�~��=�G��2<���L_uT-����+s^Cb+���{����������ֽU���W�W1, ����D�p�Z�s�.�[nj�䱑��x)b����n����#�=��)0�T"����%��9'^�x������T�*&i�%tk�T��k�v��;A����x���xs��S��j�6���	wt�F-�+����%���f/�N̙�mdC��:S�@n�pW�;�b�]��c{c��ы�Y�J�HN^��:&�w���S�S�Z���*v���\�.���X�*�8y��v��^����骘�����tb!T��v��Y�K>sq�4.;!+�B�vA�~ `�;��w�����9��=�L��u�>!w��>��7��v���S��W9�L	�9��d�a%�t�F�4��OW�=�� �@��K�T<,s���~���}���>�?c����v_���B6���C빮���2��Шo�4��v��iW��=������	��z�δ�'2iU�Gl��������ɼ�xC�"8�t��w����־�JK�[��k�6�m
�@t�ifB�ɼM-���.�n�ra��^�)t�D��f�λ΅+ius����
���3�7oT5|:�V#��q~��#ﾄ��a49gg#�ʜ���rU>�\����ܫ���gp�� 	X��>��{W#6׮"�?k��CqXx<�Q��)�/�U�����{�^��>���S��	]E{�Y8�䎫=�P8�y�Ʋ�g�S`-������ʓ*!�ں�Vf:\c�s�{o�^�Țԕ��8+t@%��>cܨ���`_Dj��V�e� <<�U& aK&�Y��9�Ԋ�F}��Q`�ˮu�U�`~$�G�%��-�Ҩ��>�}�I�7�aߨ����8�=U�r@���`��>�飥��q��P�����c5�q~;g����	QY��؊�e<s�}���e���C:+��n`���)��i>1\�w&����w˥U<o�QIŷ�jr�9�����N0��ЩT.����n$,׹��'k����G�b�����7�XZ��3���?���9e�;��$�"g>ݒ�)�E��펭�����1�xK����ӈ�i��1�j"��)�C`:ن���w�h�wZ��s����#E:��>�2�Q⯴Օ�����RP*�T���OoǭLf��U�� [��|Gm�X��=��>.����s]��V��ZkbR耐[�B5%�9���+��}�7*Xݱ�����P���V�x(I�7�m���G��}�����}Il�Y��.�T�ҁ�a�TA/���"$���6\�ZPd��A�K�xr���?��VϪb��g��O�s�/���uƆMo�U�:�B���i�ڣYG��ܓ���7(�ޓ��#u+�AI���"/��I<~��Ɯ}��j����q́|c�N�g)Im=����bN�ָUp�pr�X��/6<ke��3)���K'EF���r>6�:K��ׅS9���D>���Q������q�\�HU�Wޫ�:'ʆw�dVv�J}�Y�U>Ca2����ʃ|�C���ܯi��/��2�Nf��>�#+vh�NhQXYp�3B0���n�ra��[#y�ۛ������&�݌?;��Y_H�u��
����00s��L�����2B��ϖ�~�~{T'eX��7�ʽ�hm"�%�u3f
���dhnqCXbl���Ϡ_Q��-L����r[�Z)���(E,�eV8cF�kFn���u0�
#0%��U�ge��i7�F0o��t� uL�ᓬOL�&�X�A�=Fݮ��]���<�FfǺԵq���*)YՅc��:��U|R<.������s����sQ�}����\�/�K�5��pn�3v}IZ��p�/���M>������1N[��[��7��˵��.3�7����Ap�k��8��vdBY�\��(�:��N�����e\��$b_��ȷL���M�ح�r7��xWn���N �޶�)�D���w��'��^�eʲ!��MK����8���󒇙=N �A]�%s�f��놗��od��u#��J�YZ�̵K�+!�T�QS�%���ܱ/1j�)��܉��H�u7՟F�}Y�;�h;�l�\����Z���`�ܞ_*f7���//8��\�y�{���7�\rz�uq\*��s�2�-�;����O��yO��6y��)l~e�-�tΧ=�<�g�.�K�����_R���_�};2���_�b��(gx��c��OJ��2�y�b��`�����iR+vJ�mc�%YwE����i ����ut������;v�	��j�n��̤Ћ������"�Y,�&��:���ϖ���Ҥj�;���5�c�
V�Ԑ�R�b�6�M{p��/�락8�y����N�'f�n���]
YmD��:6�<��ұ�2��m�l�b,mv��M�i+<��UҜ�!�����;'��ı�uK�.�����1Qux���V슠u뮬cNu��8��@B��`h�g�/�T1�mP�CfSt&Ve�v�oiӔ��w�$�S����-yٵ��{\�Ι�t�EV�(w�i4�[dA]J��+Cd_d�؅.�x �b�����H�;y�u隊�UB�+T�עGc嚞�܂/���[���}1�ϔ�4�+aF��q�����j䈁�j�Nwb�z�
��u�Iu��Յ1#�Gݩ�ǃE�AT�.��7��Y�ٽ7v$���@#��
F���7���P��e��ªT��Vo�U��y���60�Vۍ�x�l�m���D�O��os�Ô��j]+�o;�Rn��blʒ�E�X��Tc��`�e]�0��2�+���qL�%�}�!(�F�)U����5���Te]q�Z�5�w�)5wB�kZډ�9���u�l���鍛�Vۺ��cvI�!�Ľ�J��J�5Ɉ���u�f��ܒ�^�O�&�� #
�Q�ֲޛr]�-�� \i�n� �9����k�u�,Xk�bm)�x�y��6U�4�t���]P2�p�{!�({K�&M�Դ^�^�����EH�j;��^Rv�&������AM]��~����Cj��ĬesÉ3It4`�5��ǚyq2t�تW1w�]��JSUp�v�R�]j�a�Uv���rl���f�QB�ۅ�ڧ�Spu.��6�U�K��^ +p�G����0�S����^���۬��2jr��5�G�]�mh�ܩX��y��&��޻x�ikKǖ�١���=�h��f�{����Ru�*�s�[�X��{��̺p�r��c���ӫ�vZM�$�[O^��mrv�X:��Еcne�"�,�͹2^�j=��s��>��w�u^j���e���.���d�GTKR.�u���v�z械���D�L1L��c�u��v+s"�6�;;�j*m�¨���IW�]R��	�2��I�._kܜ�㸊�8��Z�㭖�p�([�ި"�+�<'���pQۂ� �
lu�,���0��3W��{#[�x���R�պc�W+�m�9���quˬ�Ҟ����yt'Σ.��:0��V+�y]���|Ф��i�����"FW�s;��,���-�Uz=b*����e��% %�Ԩ�1���9�]�R�c��y%f�u��՝J#v�
�©����\CJ��j �W���^\v� �w[�(ܔ�XԢ�,�X���_R��0��B���*2�J-�E	�eȬ�w;�i��s���Vb�OZ�P�8(;����p��3uݹQ�Ze������Ъ ��r�������sB��.���U��uP��9��iJ�����RUR���f$E��I�wqZ$밢�
L�0�B"4=\�V�rw[D�S��F(����� �aGJ����&J�RE�P0҈HP�Α'�NF'J�J�,�*�+�	d��l2�Dz�z���%	f��J�Bf�mT*ڈrY�bX$��,�M��E��E�*s$��	L�:uI+P��*�H���\��D��բ�Bè��!��"E2;IP��F�Pʪ͖���*�(�SQ:�����+(��CB�����ZT�D2"�D��M��g(����U�GN�\��M7��	f������Ī�!b%`����ɤ������j�y�sm�2��d_,�I��Y��n�a��7}K�O�U$I����G�B+�"S=Zj���ڥ�[���`�i�����w���xNg�����J�m��I�a���ϡRnq���SڗU.Y��v��tN�2�R���]�����94a����,*MϲCꩭ.�������E���z۳��wX̩	�u����	dpv�477bM��l�/n+��^Y�U�(]����,��g�5_H*㮝,���H�os\5��L�l�[6��;{�������ܚ��z��,��I������r��șK��L�4�6Y&���ӈ�vDk�����ZQRp��@_�pIn7,�d\S7�R�a*G4V?���_����Z��q�78�;7%|N�93��[9ݏ3jF��j\B��8�g�m,���a>��c"����+�,x�WG4��X�%Ȁ����]�!���G�Q-�p�O5�C(姳P��6�L9�����+�y8K
E��.ͽ���&��*5�h�V��7��q493|�;U�Vn̮&�e��$orZlJl����	�+:X]��T��;��3:\4y�Ba���|�3g��$ti����}U���Q��Vy1�=�]HF:r��6�VB)�Cz.�6�˷�Y�¶�i*{�ёZu���*�02���X���]�,��#������;�����]鬝�q��j�q�]ls�n[7�W��%��/��]�7j@T$wpc�ν���g8trP뇕_F��_D�7;�s	�Ot5m�ƿ��x��>򴧲#�z�;oYA�̴�?m��.�p�3�����v-���]�}����v+d�����y
��	��Թr/S����ɸM���W��D��ݰ�QVoo�"i9[.,�a�MˬZ�A�/�[��ioyǥ�����]3�[��dO�wW֡���r����ƐL��w�����+��G��iw���A;.����=�K`� nFk�$$H��=��\c��"l�Of������b=����Rvd��B���W�S�d���}��<�0��Ü 2�3Q��[֙-�h�<U<�4M���ē�j�B��2�<"�-�A��!X���
N︚]��{�Bgtv� �{f��5ּߨ�`����E:��ǎr��b֦9s4)>�ﾪ��.O4��eq]���o�n����g���p��O��q7$���c"Rλ怠I�ڨ��!ľ�d"�Xw�U�{�^�_��{�zZ?q醐�v�4�y7+Ǟ��.#�j���s�ku7�&��<��@@��3oy����dY��1oI^�+�#�5{F0�����-�u��V�ޞ���rwf�,��ZD�q4�t�]&k�ݿ �����P�ξ]�N��я;�[l��x嫍T����Awr��:
ip�s�e�rR��Vv�$��&�n�Ni��,�t&ʕ��$<�����a������$�q�WVF��W�>I�\-p��c��_���P��:87ѥ�}�3�d��Gw �,�����ׅS9�.p������oe�F���=
~�4Wzٴ��������ҝ�m��*��e[�%�{}���{EP��_ى_4;c&���_Ɔ%ג�
aǱ4�h������t.��+8d��ҕC��u��"�y�gj���]�۱�!��]�o^D���cK��(�<:�`cMŵ��p"�����Z��n)Ust�f!M8T����������zd0�&����~ͨ>C,�ݗy>�b�����G#G\��4���Ϊ9���IN;��	�ruc���f�Yǩ��%�7��O��7ʕ�gc�g�JR�M�;o��e)�r�r_��:�v=�&
򹔥Y�ǌ�Djq�F�(h�v�478��0�g!�}�����M	yR$��g/4�Z��ri8�z���ώ`A*\C{���p����잹��x樤*wPJ'���7&�tʯ��,��I��S|,$�>.邮�A*к�.��-܎�zv�%' ��"%'7�$���L��Ƌ�4�4���o(��q�{\7���:@̜�_A��%�ҚũʞJ����R=rӽ��r7��)�����.:�P]�`������Au����4�6��w��޲:�-dKf^O�\�ѩ�V|�_,�YV���ӭ���2"�r�Q�}�aФ1$S����Ŵ������{��yL��}�(��>��J��a�Ω�ٕ���1�XW&�m���4�����r"�u�8�*� �F>�M$y�.gs����@:�R�HJ���tYɤ5����>��x�\_w�����R[K�|�e�uAi��n5�ţm|����b+�gӋ���Dؗ�ԃ�r�)�wQ{Y�W'�WK\*�����8w���þ�}Xc-�]Ax%#���'p�u�쥱�������z��=�$��вgl��P���o*��.5K��cup�g��v���<vn�
v����mcq��q� �S��1�Zx��z��t,ã�%�u�7!�n��N�E�4L�q���79�ru�ݝX�iS�U��V͍�Ut%��!�L�J��i)���	dhq���ö�!Y�ϖr%>�Is?)nx��S���i�M�N�
lu���:�%����nN$�l<l��E�1m�����s6����7l���Jμ�N��	�d�=���p��	
Q�L��3W4�D;O����S=*/�g�>�v#�x��F���Nβbm�Ru�S�o"�+����f�`�oy���l�v�0�m�oŭc�W_9A������@E�5;����XF�T��#�G��p7���]7L�'j��l��h)�\�7w��Iu�Mӟfu5��Km���g{�r�
q�J���ﾪ��\q0�5��k�yv}���\.��WdJ�nI���(K ���.dSᏧ�����q��"�V;�kG�f��*!�7ri|K�ETWu�;� ��,cɴ	{�!�������/9v��-��0K�*�Q	��+5Ru�1�������E���+�GYM(l�R�L�O�M��I��Jj��j��n�U���D�+�����Y񴺑MsC�.����p�o�r"��M.�o}m����L�e9j�{��p�b:���������TL�#��8]��ĽF��sE7����4T�����lu��H�4\���Ar�aõ��Uap����ã��u��V/5K��jїn��_vF+���OJs
;����������\�[���r��m���T�-�1��cDN�X�}�O�r#J��e�|��Zj�L��۰���P���޾�1�V���NM��	na�����h��3K���wd+N��;u���*�÷���٩N��Mm6�n�� M�����.�dרn�y�Wh��jR�e4��� �Z�#g{�(턹�1�����ԼЖ�EuD�����G�|�i�ŴM���#9�T����g�I��q�Yc>V���e���ж�z����0�oy$����̏����Z�s^?4�W����hy�W��p�8��[z[fl��֗W��v�S=Q ��˨:�E��ؐ(�����]-��n&�ϝ��/�`5�z�U��^n#�g����[�w�٠r�ծ`w
���o��p�녦O�[[W��B��m�i)�Z!��E�U8�\pMb�ݾ�	=ϋ֎�8޸fnB��5	�o����|�A���g���M�-n�n#S"�d¶w)q�`���Im�[�}.
��LW�I�	T����G�~�=1���.�ǚ�=<|�1�o�2�}>�:�uҪ��@�J���I��6�u<oi3�����i��ڜ��{����l�M�j^9x�*@T�����})�ڼ��l�H�g�l�R�.� �(��1����r�ݝ��WWR۷u���V��z�5v��c�f+�[�֔��C�$�$ii����� 2���Fu�f^mg5����
i�Tu7�	�o:���Ⱦ�[�n�]wo��N_`�9�F:��w��諭�\��L&�1WQ��}ɇpٺ�����s�Y��*{`����N��6�&�8�띕14�R��Eym)�:O]\-p��6:���=�wp�>V�<��x���޹��o�Kڡ�'���i�%����r8tn���ǽǃ��g6�yX}۸�}M5�[�<��������.y~���+�'�̋�W#e�^�!�R�j�����/`�ݸ*}�FV��G�i�!U:�d�����3d�þ֡�ܧz�D�άx4���"x��18ZP�(��L��.k���L}��)7)�|���B�Y�6�Գ�;^��VUu�zoJ:i�Y+�W��,��gѡ���n&��e��F�uv'kt�����Jd��D�ﮍ<���%�߽����=��D��#���<7r�j�kS�&��2eE�K*.:�K�3�S|,$��8>��Nf/�_r�Qm���V�:0/��,Uq�2R�dsT�]T4�4z�܊�X�FB��«ŋ�l�wC>ɂ�:���aJ3��&S�M��vh�y(�]7/L&��37�]>�1�����o��f��d٥`�ãk��y#����}��TZ'���n���Z`��gPK�����Rz��I:-Ll�Qj����qT~x�8�Z^K�{S���@̞__ %�{j
�{Wպg�4��s�=d��&�D��%���S���p��)s�����\�	cU´_)m}����Pٖ�^)N�~T�9Qj��WRu٤;Ǧ�qȷq;�G�dm���=d&ٺ�-9y-ƺ��n�6^�c�9o�维^)k*�5�W��*��,*=��y���r�^#�F�RV���GS���!����Irv'F�޷�ԋ���"����QJ������@���_ڍ����Cr���Ae>�R����y�Y"��6y��J@�8d���w�^|��-N���д�ϟ�v�d��krɯl]*)7T��1��Jn��}�L��Pwh&�;��	�vGgV<�D���dI�s�Tm��ʋ/�0�;h�i͸%!���	yئ#h��]�g�ǿ7�Z���9���*p�?l
�i�w$�"�F�bD��U��l����ԥYg��u�)�ak�hsš�A��쬾*r��=�]t�@	V�Pe���nkv#Ջ2�W]T{��>�����d�)��S���oo�iCYae�
�s���g�E�ú�ycB��$R'��M���(���O,��uqj�t����&��w{�}r�$��L ����?5�����
��t���5+Ae��L��E=�,�=U֞�ks�m��i��q7&�������:�i@A]���!�f�J��u�Ֆ�g8k��p���W`����?��J�i��Q����ߥ�Z������W�l�|V�w�o[s���4s��
k�g�v�͍$r8gy����K"^r���ۜ5�A�Ǚl��Z�V`�_#��%�g�h��C�Ƣ8���̳��P�[;bf��g$ӮK�l����H,�!(�Ⱥ\֮�����qȔ�&5L�zl���Y;��{��n1�Y * ��	���]՛e�?���&(<u2�&��qH�m�N\�5�/�;0�o;�,��e��eJ��R����N+f
}l����WeZٯ��E�t�l$�8y{�{�qw|�n4���諡t��J]��@֧#��h�4H���eu�*�;͋Sb#MT��v{�
�)��Wt����{�i�	vs2�,��E�R����=Vr#Ԩ+�h8��ʥ�fJK�m1o����c�V:$�H�^��f@g�DF6�%ӭڜ,;�1�������;ڵc*ɺ؂�@��3��;�4�c�B����9�(Z7yl�Yn��f
v,X%����RB���*�����Ĳ�O{��޸f�,u���1h�����+�J�6B�a]p�l�V�kU/��m0�n�h�I���7N�$�%�����vy.��0EFn���h�N�cmͅ����j�]�tAfN�:������0�2�%̊�bGouIͤ�ح�9�_w�=Yh[�*����ݶ�ĔMdh]��� �5�2��X�+���2�5d��-h�V�T.ݍ�g.q��{}+,.T��e���򾇍&�5���9M`v�u�O�<�ŗ�]\���*��RԒ�m!���Րp���a#W9G��&��C�u���6�oV��Q)p�S6��F�Z[lC�۬y�gJ�	��q+���B�n�i^�Oo���`TU�]w�m����N�V]�by�L�����4s
�H.��&�Vm+L��N�h�4]�+���򕪹�]K�8����ܤٖ�>�d	 �j9���XYc����*.Z��O�n���P��B1� �,���V�S)�͂4`"���m���hp��&IF�{�Y1aޘ�<��)a	�ӗ#!�ڸ(�U�A|�TU��fҤ���wf�_{�j4�Q*m�WԮ�C:U�f��ow];/]��Ib_[��f���rX׊hmVv��k1�R���%�zJ���Uu��H��+s[Yy�;[��v�+�ǚԽ��5�Yt��t-���J���ڶ�tX��b��;2�d�r�Ҡv5����cS�Z�c��1H�6�3�Mۭ	��.5�1q�"z!���#%�G�C43,\`u�Jڙ��=���V
K���$��x*��e��G��mZe0���*D�^7{�KToWt�	���`���(����������GL���qɃ�ӣ�[��R����i��K3�g�Zf�u�\��g%�)�Ni�⣼>R���^�Ig:rK�W�9Ze0I�ZO�^�H3���ܜj���Wq#W��|бK*Eۋj[aN���S f�o��r�j��\�#��Y��θU�|8��<��^�������-]��r�Źv��)����
���,8E	��C�g���LT̴�+f:*�֫|�j���ٮ�Z+�D.�r�R��iJ����ܦ�ݪU4����r<�݄�
#� �t$%I2!YP�b�D�Hȓ��Y�����)2-*�4Zr��TVR�U�T�4�5S(�KaIBjjb"�Qj�AVs4�����T¨��EFW,���VV&�l�Jdhb�X:���DR��B�2NX�D�0�i�H�&�����C�F�̹U������q.T���Hif��$�VU���-�QQuY�&�r����*���%C:��QN�v�YE��T�:�TDU�+:T2.\���L�t�AW��EW(�MEJP�B�B$6�����8�is2�	��W*�!"�5�2�j2��i�JКtM+L�՚D\%T���Qa�1��D���E0�͂��r�1Yq����\k���p�<ݨk���[��8+)�Cq�C{6���M���#��-�~�VIY�X8f���r��r&8���UUU}/�z�gJ?Ţ�������q�!e�s�5�Rj'\Kť��� �,����N���+i�}����z�vr!s�G!���U}�_ڥ����N�e�vt(�Q:)��r��]RSڎ�u9�}Qy��з�ٍZT��ó�a	go/K���읡�Y�#@[9��n2�U>A>g��vjn�[��v.����-~�\�_T����K*������,\�=�[M-�I���~ZR���|�g.%����ߖ����P��z�E9�:@Z\�ޔɭ;���f�M����;=���Y�6�L�|��������)�L��qN:�7�jv�877�c��!6�;O�_Wǰ��jRR�V׬þ*,N.�.�{�=�0+�j�zy�[��u�i��A\�� Li��]�y"��?�@�X������}R�΂����7���릕����v��}�n���C���y�5�׸�^��1��7�,��&H��h��ƢМm� �G���������y�*Ϸ�U&���q�79y$�%��r(^Nb��Ĝ 6�FsU�éRW�^^㙐�҂܌�Qڞ����G�D�I�V��'�=�})t�p-n�!��S"�d��T�4r���������⻦�nr�t��8�,�������O�'%�ږ����1����ю3���^s{��ٶ�)Z[�	)Z���U���qtn�ߚ4�v�s U�#����f^D�r�@T����Ap���iY��Yh�v��i>���l��Eu�a�͛��
Nj��dv$��3wUB�E�Kt�N?�S���m#ݱ��Vo>�W�!'uq\*M�ŲOKV�2�hZ��ʳs,K��yW�o�K����~f��ߑ��s<�j��&oH�����F��o�/��:��eꝩ����V+��s���f��=�7Ѫ�a�֚�����-cV6�f�A�u�3�T?Ne[����{s����1A�D�KN��+.1Rn]b�M�i^A������+�R�7���@�/�;��X�mu�b�����5�La��_t��8�Eq��ۃ�y������Cұb����\���g1ae׫��^O{"���q���ޔ;���&9,˕�la
k���^JZ)��ua� K�\�nCG��������:�2�q��}��g�F�g%�e&�>v�d+=���_g`�F��z�f��G{���_]:��	t�Y-��5��g>v_v�n�e.�Գ�ë������U�ѧ�s�Jі��Cu����mk�&���sb=K9|/�T��I��D���:�Y�;�����M\�˪���rx�oJ�ݜ�CҎ��fv�%q7$���B%'=),7��M�4+X�0-m�0ҳ�/w!p铒���N7������i|L��f�uF��u���j\!�wa�7���4�^r[/vZ��T�%�o�+=����tc�K���"&��l��A��YQi}-�y/�Wq�Q1N���Ybc��}=�����[E�#��u��	��َЯ��;�t񌼷ؼ���U�����vD�Z���L�M��B�@c9c&=8���Z��'��Gq,曹8݀�����N�6�u��Bd���S�'O�ڸ�7L��;�,�.�C����}g��ˆ������0�y�h]x	�2����dljҨK�pݽ���Q]fK9Y�kV����nG	g�꯫���P����;u�c��ێy.��	���Q��l�=��Z,�J��ͩj��o>N��On����n�B��|�\<��/T���:&l�Hd����iHǱ7�E�%���;��/!U>Z���{�]��S��L�}֜n)�e���޻�Ƽ'c*��Ms�ϴ���e����v'}���Bh��ǞB��� �Փ�CݟZ*���M(k>�ⰲ¤ܨv�H�J�K,�/طW������w�F�ʉ��V��K���ncz,(,��W�33'cL�d���}#�k�E�j�]�Ԃ���,9Aq������(|H���y����ks�m�v�d�' ����C2F���sԲ�&m�ƻ�u���o$�>�vk���2� ZWrh�̱$��b�N��RZh���������;f�6w �h�s�돛���F��R³t��}ΨmbԺ�SVr�����5P\;�B��Ǘ�LzA6�j��-:���\v��X�6�R|���$�h)���%�5�1�i��e����!p�x��M-y���B��!]�gkф���u0��X9#}���n�l(���筆�zٯ�U}ʋ��hI��T�}9[����L��6�;�>�Ǽ"{boNk���Y�ݞ�u&Z�A�f����
���4���3M,���=ӹ8�N��*�_.�BW�.�:ύ�Ԋg鴱nF��k��8�}��\gq�m�y��G���S 嬱=Oz�"Y�-�����Ջ���ܞ2ںZ\��7�����&��qR\TQ8�F��FVm�d��z~�W�!'g>\����:��&� ���rr"��������{��0��d̓h�dw'�X�⩜\�[���/��}����G�
t)��Ad';���W��D��܈Ң�q���������%&fC	���f��.�
u��*��1�=��Ǫ�,�rf�3���mQ�6�S��qk�������䫉�c���nY}כ�-����_l�rjԢuw;��P.�4���c�tj{�3���B�ŢZO� ř�STQ|�juF	���4�@�}��&�6���@���Np�bh>��eC�c�Sp�g��u��\+��PՅ}Y�Fm.�o-ϐ��S[�Ν��Jҳ���W�)7�8��;=�6�L��u'�	��6��.����F���5;Y����[�	�q�}���`9�:��S�k��a�]s8�
N.��t� �q�uqɾ��n�Z�[��ۛځ=����O�_�r�L���I,\pId.���갓܈/Z*4̡�Ŝ������8�n�v8=9N��������s�kv!:��[4_����qnyx�S���ѣ	��K���1�Z鼫�(6�~A�K���<�f�^=�������&�P�%�����V��aw:��[��>6�K��y��[rƓ������R�>�.�!6e�K�-\j�AS�y����s���+���n^`�k����仓��Ai�_͸琲�򸼁�����Ue(�w�%ۗS���9Q��wR{Ky��+ő��t�r�5�X�=k�,�YzM��$����ߍ]�.�G��\�I�����v�B���5��Y~��=��Ы�C/q9�uY�{S��=�����	�����nksۊ�5�&oa7�paF>�`ϑ{dl�s\������]]mk�/�]Xu��(�%��#������~h���Y�����nU[s*��jl~f���t����v��[��#���Yd�T_Xއ�������'uX�fW�%j�3/8c�����=��(#�SV7׻�e�s�a�O�mgv�J�v���;��\hqQ�\ ���)蓪|�����O�{t�:��D�DO[��__dӄ�C;-�|Rnq�}�MiwӞ�
TL�S��S�9ǚA�����ʈ���:����K>��l�'5�	�WA�Fd!�I�c.��Q�����`W�����H*��O`WIZ�!��R<rc�����Y�����dp���Mɢ�M|�T_�i,��Ϯ2�N*�ͽ�9��&�v�P@�;��]��u�3�%�7$�΅	9����"�j�%��������w_�L�'�Z�'���t�AWĎ�++{T:�e
�P@k��T�ɛ����^�]������;;�gKB�=����&;pN���5jK�Mܙ�i��V��W�[�F��١��R�3+��,�I�Ku���Ѳ�f����*K�j�u����K�Z#3Wb%�y���\��#�B�	h_�w���#�0'�s��Y���^��59_*C?��A����J�Y���k��4�҃w��(�t�/����71�E���R�2������u�\���]X�w�~��ܭ��{�#���ٌ�m�[T}���-�F�U��Ȓ4��g���.���x�Jy��T���%�7O\*0��y.��	�.MN.�����\Ҳ�ȭ����=�W�zyj�A~����S��.p��ϰu��9`��T��E����Gi��%��RҔ��U3:~���;l��a:-k6:��͢�e����e[
�%�3ݓ=�j3��sMN���R����d&eW-���%
|M��X�g1�Y�7��4���ⰲ�+M���G��뮲Ot���0������gVv��K7�YR9\u���P�pv�3�J�ψs�"����
Y�Vl�2�n����{�(.�`�zzl1Y�����ۮ]n��]��p9G����eݫ���V�Yu"���u'v�{��)��[ziWk�)vT�:Y":,=Y(𾬱���B*"�e��e+u��6����y�rJN�cQ�<J&�*������x��e��l���zKȉuJW]��O�5)RY�5�a6���k��>��t����4T�W�F`Wk"�T�5��e_=�'>]a������>Ϲ�]��u�2�>�����}gD��q�6�y"���U꾈j	�����W��c]�3[s�[�rb`=������l����~�,P�^��И߾3��zJ��xA*�|��}�����_�NS�(�+䣧�}]H�R\1���96Bw�"�;�Ƃз}V���/�q��
��u!(頹уiuq`������^���x�Nl�\h�Gš��W�2�[�j�*z%<��D�9w�0��E��==�6s���rz�UF�5i�殶9��*H���̼�ي_(|Q8)�J�n�vu��;�\r�I:�s��:�T]Iy9����L��k����7u�u�JXr��-e2k-]���U���#��G�tt�m�/]��^mս��cⱮγM*��j�l��c���X^G�pe��u�yn�ƅ��N!�Fx�Zl��f�+�K�bM���D��N�j!|������d��r�=���v޼���\�B��{zh^aL��u��;l[�����uh�}�M.��Ң�d؉�����W�K|K��ǤruW���K�}����NН�ʿ����lɌ�Q��.���#d����Z�r��{�����j^�YQ#�R�T� ��	��oN��pp�[��Z�x�ϝ��g�����zr���hoK�zY�NB�@�S	F�k#�sx�ϓl����}���.Q�g4���u����T�\��:��Øµu|���9�[�k��05+i�����E��ˊ��Tɠ�D����.���ꔞ}Ui����D�tR=�z��8��zٜ�T���rj��_%Ӝ[���0��#�j�*�2�ݠ�iy�������t��8�*��"]/��̃4�)�|�Vo`���㥊̎�lO��^���X����(v�kM�};$���s5[��K����J�FV��&u&���Z[��8BNl�:s�L���nՍ|	��%g�M��U��" �ک����D��N�d:��teu:wI*:�4�״�-W��L��L�C���Y@��9b}�KFoJ[g���H�k�a4�*:���j�3��;l��Yŧ����p*D7}i���;ťP����lq�;/F��-E�39^W�\ՋVV��U�37��<�P;H��͢�@3��]hx����6���|*l��%�p��hP�"��`�<+��OT�k.�mgd�R�T�'^�6e z�i��&[Ƕ��Eσޱ#���<n�N9r{X����L����.�YNM^����Dn�C���c���o6*Ovه��.�>j�bqu�kr�G�n�8!��6���P���<�R	��I1��DF��Π�J��[fQ�ׄ]X44��b�M�u,vJ���vz�jJ19�����;��]�ȣC/`;N!�t�UǄ65���x��9�J�v�aE�Z"{l�rU���}6�����f����6��|��W��N�h��VE��2�-Ȩ��]��x��1n�:K��ҲXڸj&�����$�+-��!��Võ�X�Ζ��ނ.��z#.����S�S%��N)�뽡WI��%�.��)Z���e�����#��и�1���ҲL`V&\���
[9����Ĉ�!j�b��d�.q���d@oe�re��Ԝ"�%l3r���Ӛ�e���$��O;�31��bf�� �̓R֐�W���zN�5�-�{K6�2��9[Z�/!��b��r�t��3�ŗ��������4�	���e�ݭ�[����;���􇬎]%�Jb=�p���ȳ��T�I(�p�7�튘=�,�y�O�ޅS	�u��bݕyܸ0#�tsYkS+V�U�|��+��/.�K�9������
u}��@Y3c'zR�첬���k!��Om�Ȭdsj�T����۩�m�1񅊏���eIa�YL�F��D�[W��㠘Y��RP����;LR��\k�o�q�rd�Bl�ybr�f�����9[R惂hޏ 3]�w�٤wH�d_�U�a��^>�w ����tߐ�Y��$�lv�ջ9�zG�ч�Ύ�U͖{R�6��V���Q�u��.W���`��Ҷ�l���3d�'`d$���i*�
ˍ`2����1�7jk���o��Y)�򵝨T�A�!B}c�W@F�h�sQ�em ,�޷J���R��o)�պz]n��\ѱ7��=w�P�_8��,�yif�T�n�b|BnU��%,��m�ͬ���Gtu�,��WB(������9ˏ"�T��7��+��C��M%�2]�eh����C��Ur����7.W�P��o(��R���)Zl����8U4:�e\�5iQHt�SCU�U�DT�r ���ұ4$V%dV �R�Z���2�EG-J(�ep�.is��bQ�J�bdl�$�q3�\�X���"Q�XfQtE"CaEUtQ$E�iEh,�1CU:�V�E&@r�X)#RV!Eə	d&d�L�I�):uP�"3L��(��
#X���T˔PU!���B�DQ2L.�\�.Y��S�DU"*�Y��3�%EK0*���t���B*8G.Z��
&�M��af5L8��UR���I�AsZ*�*2*�a�U�d$r��"V!EDQ���*��Ua,�B����IT�jr�J �AȢ� �Z�5H#�R$�,-�A�$D�r�]ZZ��QQ]fV��*�T%��):�T�8��#��t;�+N_H�ǌ�ا;�Pk���:���̍ݮ��f[)�9n�`G�5v����h�؇��-�*}�	{��>�ԏ$2>��ߏ�Z�ꗜ�Ľ�j�aZD�M$۹f��B�^����n��Nr�;k�a���s��2�%㗐�ʐ�U�F���[���h�x���?�E����<�i���u�ra�f��Ni���j����:"~������������v�#Kc������bN�[0�rCF�|�*�h�R�|ZgfQ�/(��U_ED�T3���c�?S~J�e�����?rO"S�ΈȽ�����چ�y[�S�g�.7W
�wV��9g뜶��-0RaΒ���m~UO��L��Xۏf�!��컜W��W��\sv���)�g�L��
+.2&����8s����P��ȂU seSk�+'�N�3"SϺ�����rQjU%��V{��/+�Kj��L�Gz�=Xř&�ȞY�]:�P�����hno5��t.�<j/�_K��51�b�LI!4^;R3_,�R�V��p��+�(��̸4�GmL��m��_��ᳲ`�z��(l��nC�ҡݧU/D�~�Z�SE�D��M�	��jG|�K)5g��܎�g7V�5V�PB'6Kn����=�RHˮq�%�4�
�+��}P{�3���q�F�������=yw�@I]<a��K1l�u�z��)����e��r���*��,�:�@�s��x\5Ef��+�������k�\.�fu�&����j (;��/�e��ґ�xڗ������L�&V�ڜo\79P�2fDU\-�Cr�����}w.�W��И�}BzN�r�����jrs4]Ѝ�L�����׬����:��nzd�Ym�7q����-d�e�B�k���J�ޠ��z�ێ������$y���m�Ո�q��ƥ���v��gq��Y;����/>��^|�'bJ�ؐ���FR���/���'��"�7EBGo{^�Ӊ����\'��_[Y�#|6�b^�<D�K���cp��sJ���5m3�K��E:��.p���p���.b�F����]=QڄWuiTݮ)�k��j5��87R,���$t#\"��[������F���K���Q�ɂ�O��>�"�E����ov����a畹I-YԾ:�����2A]�C��4�� uc�a�â�ҙ�֨�])
|A҉��e=C9��{�����u��U>Z����sm�t��Y`�k���A�'�����6�`+�=m9�Z��|�7.�o �Sٮ�O4��(�gk��Vq�텐�ߍ��M(keŗ�����sty�M����ɝ��~�lk��]x��,��{G;���uX�Ӭ}]�������ևd�s��g��Q
^�ޞ�׍�v_d��6���T�J�ځR������:D�+�����H��5�[����;O�񸛓PT�Fj��P�q2�s3y.W`��. �O>]a�u[���v}�c+L@���h����\��aZ�FH��1��JI|����횖�w�kGc�od\�:��&��j�.t'꽷�?���Ez��&���Nik��v���Q���x����]�78�d��Q�>�\GZ/�S
���Ub��5�[ ��u�#y����x�)=#FS��i���݁�ڟ�5�:� �~������.Ur:,��G�{�6��R��r�Kr¼o�u�Y�a5�G�4h���%4��20iJ�3�l5�X�¥�N�Q˭\���u`��"V��i�䟺��~귊nȥhQR�RȞ����Yb��]�j��,ڑ�k�憥Μ&̼��^|�*@=�y��Xb�`�&��t�<)Z����]q��m]\B��q����	7;�������}�cZ_e���S�V��o�����4Ω=���ã����*�� �Ɩ���1��f�xv�[Ϫ�=�&X���;]IOo���QT�L^�c�m�tn�Q:��ݜ'4��MU<��}m��5m����=��9��I�g2{��G��꣘�ڥ�7̯MK�r��r��myION�����))��n�p�]�zy��`´������EQi��<���χ!s�C��%�D�Qe�J��q��Y����q����}�8��g�Fv�t�X�虉�j�2��\�8�B����u �5;Y���aM����|�b����R��n���6+��¥�мt�o2H�,��
��:Ty�.	*�^�!a�e��g�Y��7�j����fG������'[���df�����z�sb�0���Z��:Ov��'vFXl��V����\m���g�U��T%��>9�\+WWɾ�eݥ�P�dVs6�v�ugj�-+��P\ɨ��}$�q�%�.������6�eƘV��科�ꫴ�V�v9���3�����fW�l����	i�d
�manR�����l��X�'�&��HQ�T�~�"k�<�� S/e�����q���SK"^s{��ٿ����hW�I`#�?�_Gb��a�Wv��/��k>6�v���#�⋤ٖ���^,�p{B�ؼ�����Ȼ�R�yO�g�iudr]|�vٺ��Nh�nA{�Y��S��'u.�1�� bj���]q/*6��޴����-&�>w����_r.w��5�uj~��:�m)�B���_e���p�,���҉ڙ4�<N��Ony׫�qs�G`뇕���j��S��U�neo�D�dY�	6��V�n-L�<�1�N9cVgn���2�,�8p���1��0�V��J���譱�̣��˺�vXޘw�G�S�]�!�2���9J���!�k
07�FB�SG.�WQ�����������j�l��쮳��Y�J�13�"�h���Rw�e�*��je��g{6��ˈ.w\��{aqαY��-.�q<��V^��99��Dae�|�78�Wd�o��+U�w�iX��j�S7�΢2�8=;�D���w�4���LhnJM���}�_f,�v򲃄7�����l�t��ϖ�k}q蝖�[���l��#�=�8�p�5&U�f�����>907���e���ڙꀝ}
��4��7�[����xap�5��y�幮��5������srh��A|���ᕍ{�b]��;k�=G�%��~�����p�k���q|�+�&����Z�E��+�/9�t���y&Qeu�	�]2r%k=�'���|���\k���b0�-�w�X2}7[���Q'"id���N�鞎}17��B�u�1QI7IGN�E�A�do|Qj~�3�S13NH�UՒ���D��x�jC��=�-�٠��i3����J��ks\�~r�{R�PbV��fɎ�Y������ۻ<�
fd��J\�4�q�;o;�VfN��M9������K.�wZ���]45�x�d-���؋��ť7�kH���U�2��y!�S����\�>���:9�*���ʧ3��+M;�r�Ӗ��ן,	ؚ*z����^Wє��8Y��1Yj�O��)�nV�Xv�z�+�H�_�T:�M�<��Q�Irv"�)�5ҕ+�[{f����c\��t���z��g8tq��yU�x��Q��'�����g�{�JC;Ǟ�k;���*��a:-l3c�%��;�X߼���W�4z�uC��}���3�˔�y��d��}U��x�1/����Ҩ9���Q+���o8��[x"?U��{}�JJ��m����z��,�ݪ;��>v�b�ݐ��;�Z�l,������yt=��x�y�ߗ�s�Yρ����-kx�ϝ��/����Z��ֽ���q��5D��`�#��놱F��;O��%ĺ�x���J�y���u)@�n*����[�n�f���]�����Gj��.g�ӌ��g���Mu�[\u?_N�{)���5՗Ն�u3x/�%��rTW��ҏo*��¦��@�<B��Vm�j������y��Z�1���(ng��]q֛�]a�u[���v�Zc]X�6_ vF]���<F,q7*��ξ�X�������R��+Z"�<�C���G�-܎�T�:f������9��s��؄8�g����j��;����#���ܜG���nq�2�7�2�Պ�7��}ykwƢ��jQ콼{�:�iCfZ��nȥhe9~�m�ַ��{nB����)�{i�)���넋�ٖ�%�א�*@e9j�L�b�:#�����C=�[ʌ���l��V��=m��K��M�<�����lʆ8gg(�w�%Źq�����Z����t���'���z�����7&g�ү*�$�i�Y�o��d��.e_G�Lў'��v�)�GO����D)���ZP}�N\�J)k6:�jy�����o�/n��S*R������f ����T�[w��`����^���;��f`#tF
\S� VNׁ��}�o��X�ol]q)r�W��X,��\��_b�s�[U��톘Lwc�{�P��+����\�ep��ʱ;���T�*ѝ�|��=ԓӜ7�i6�m=5������~��Y��u�}�YS�aeK(T���fgA�5�����;��_�Tae�V��X��ܾ9��6���'a��%��e��3dmmZ>�j��[ꓪ88W���}�8��d<:s��u�ޣ��r5z6��p���㮝_Z
�5;Y�p��7-��_k�<�����z��|���3�|�Ϻ��ώ`J�a�S�X�wU�Y����̴����"�O��蛒\�؀�D���Id.���w��E�6�j]�[咽��q��PE���h�s��fr�R7rW��P"R鍘'ɷ��D�Jh�/��g��1����9���O�[��t�&��	=���0x��Nk��.�m��M@��¸)��/9���7dTB�&.�tp"�8���{zs̶}yޥ}�#Ϊ{"F�5��Qui�/>��] v���ÞØ�.����tՑ��%�KM�
Ș��U͹�������q�]�5���^Y֕uB��gt�H�/LF*{Y��3�[ȣ��Sm+ٓ���۽r�|�*��qI
;�;������b�U�C��.Ov�G2��}��+��`�dȡ�� ��֪�:"NVR�Y��VDr]qɇ6n�NA���E�m���=�N#OG<y�����ϯ��i���,�+ɻܴ�~T$���4_at���'�=�^X��z�]�?g����y��/�^'�i���?טvb�v{:�A�+�s�9'^#gg�S����}f�G��Q���͟V������ciO�"=�cgϷ}�)O�s�~�C`]x��b9W�0�,�k���t?R�{�����?1Z3ٕ��ʒoӗWY����v/��v8t�����Ӱ/�­��s7��}3.���{/�/�������g�/WP��)�\����Ƕ����NĂ��=xF�w3�/ҳ��H��߳�8��v��v��q�6Ujݗ�g��$����NUp�����NL������[�#ٓ�g+kB��8͊�qԉ��[lO��$;~�����S�;Yfm�B���B�{*ՏtwE>�/j�{F<�,���'2�ǯ�7��O���L��zyEe�Y# ����N��_k�v��?Z��ʔ%^5���݋�J?v@��؎
���4/Z����E���}�q�-��P9g��:0wFCCqs��aЯ�j��@=}�:�JB_	m�)M@�_T���q��s��T=�����L�������$�폠]`��@���ۛ��D�*�~7)K)��C���u(T�r]8�]έ��'2�ED�X��y�B�K��y�u�й<�Oc{N����� 7��H�UEu��Y#�S<�;2GP$oR��|���
U��|�yi�]k@/�Ʋ_r��)h+�'�Ż��)WǾKC]7�-�_�4��ፃ�2�3�w˷A��A@����2�e�ĲpSB�t{3�e�ɱ�A!NZ��M��]�����ע��M9cLckfػ�ȶ��[|�6�Ǝ�$�=�iC���.��
j�����	fT��r���[�Fm���ӧ��-�wk�a��0���r��mm�1
�1�X��Y[��;9�ΊE{Ī�q��`�MH��Z��x�o�Fk���P��f��\"]q�}y֮�4���+#��#�*{q����`�i��e*��L��=�����������G�06�җ���^&M:ת��5y�Yi����f]���jU��٩�`B�!��5J���Ѐ=Y���O5A7o�+��[�F8���D�۹Q}��7��;BP9��e
�(	��+���nHb�.���`a�{E���TT�ZFݱw݋���g5����ۺ@�v ��8���*�˴�pc�}-B�Y�.�Ko�r��v�ʾ��`o��d�����y(b&۵Md-��`�R����5����ޡH>�K{�ھB�d]��q�Y��ٶ����lu������(J3*	A|�˃����g���	�.h�&;/�u��]���Vs�p��U��ЗW½z!��4_'۾�ҭ�|��������4	Krbįt#麓���6�a�
85��ut���o[�ģ�b���Ż�;�T�{Ӥ0H�Q����3lMR�R�0��Lå*�Z�P����H��!����\m�Z�aU<����j����zog#��Ƶ���{3�k\��#�gS�sKU6��gUܠ���j�$*:�M����lQ}5�=+,^�H�z�;�2[.Ǽ�N�o���r�}�S�
��� J��n(+�)��5X6,+jV_pC�e�wJ��/f0;"�v-T�B�9˲�Ky6�����U|��<Y�W�+[�һ���PԦ�W5�xQ��L5�u�F�vg�mT:])T*��x1�EqU�N���}G����o�㽉$�Њ�@7�
�b���"��U�]שN��T+K]P��j�Z�D���Tp��`"#�]ld��͘��h���$&i��rI������hgpc(3ʬr�G�׹���6�j"yN���X�P�r�)Y��cL�1bn�(K�0�f�:dMQ2-I$�������Ĩ��кe!HEE�UHF�eI`�A��r
�L����EP��) ̹WUg
#kN��t�+6���Q(���&����!4,�9A2�Sd\�(NEh���Qʪ�L�C�V
�� ��u6H�L�"f���N�5
*"�ND�X�dR��f!Td�G*�EE"���( JjR�)$�Њ��5�C�e4��Q�$W9\"�V˅֬�ɦPB�"8W(���*�D�*�J��DEtVP�*W.d��FTEs�1
�9�+�*�2A"�EG"4J*�"r�E#�$�9\�R"�
(�T��R �E�DT�4LP-���A� ��S)JB*��*Y�2DL�IJ��U��RH��*ԨK2K�\��S"I?X�WwutZ�m�
�b{���s�0`{������][d1'[�i��Q=&�Q�o&�\�d�V
4$����}����TG�u�������)�r��"��Y�{��T�2;�X��{["FHB��ڞldۆ�#��ƒ�c�9�� � �^T3�P�~�5�z������~��s�z�o���&�z}Yu8��V�5�b��T8_�L�.��lО���%��b�;�?<s��q��{j�|δ{y+k}�B���q�wp�M�7 �K֬b�hx�1~�gyeI�+�{��tO{�}���pv{f{� �>��lxl�;yS6��bD�n/m�������MX��ׯ�ޔ{o\xQ�{���&��=�O��3��w�O�u"�S ��*�ճ��Y�z6W����7��lzW����L����߽�cz�]���\����ɲ=�B�U�{g$�ml�=��������T߾�[>�e���<��t%^# �vC����k>�����r={b�.�snkƩ߹(z^��h�=��w;^��=]>ȫ����X� v	�>=k#ҝߎ�������^_*�cȟkv1.�٬�G^��[u�>�9�׿ePY���8����%g_���~��TO��P��O�6��իUM�K�[�1V70̘q�ԡ҈W`pe�}���g8��Z�\�:�+� =Nă@{es9�K���������E{H��v��T���n��:K�9�nq��jm�W[ô:m�u1��@q���g}��)�ɰ��j�ڶc/�nِn��{޼�F��3{�� ���P�\+��;0��g��	\��G�/\��\u���y�O�?z��_��l<Vd��3i���@�A�j]��W������m+J�[����bSkِ�8z�}�������Ǳg��VY���9�: �z�V����p��>�ϯK9�7�h�nB˵u�շt�sw�������|�W��G����v�s�g��'���#~�=��!�@�3_HHzp�y��g.�3��ɼ����;��doz������%�E���~��w/Q�N/�+�E���R�J^���M��>؏g�M�E{�:E�@��\+Q4}���՞��'s��{�G��.�����K�x�~�T�tCۘ~>�ZV{/����,����Ͼ�Vzt{l�{��2@���#���s͜�P���`�'�Nɻ|�������i-^hn����w��9	��R��Ƕ܌�;ٛ��1W
��M��3!mѿ{�Ʃwfn�����G[y�{�xS�>b��6��1����a������W��HR����ܫ���^�t��Sҡ�r��:-�%�����
O�ذҨpA�v4����xR,^ե��+�<�S�h���(��y��h��d�Z�p�i��]:r9���+5�2Uʻ�'*lW�r�9{Y9C��1�X*A�t.�~���N}�&�om�"�{=l�j�_�#��̱��X_?W�O��>�{�X#���k*{�gpPA���چrk��G�t�-�7�9�t�ߛ�-��xU~�?+���_k��S�����y��7���t"�u��k֟��3�> �n}>��9䧷D�ͿQh�*ӔO�}n�>����W�Dgm\���N�`n�¡x\뇕{� u��q^�P�q�i���n�{|�ҡ�ߋ��y�t�et�Pĩ���OA�/��7f��n��*�Sދ�ݞ�CEטoUz&�W�z�Ņ��Ǖ��<��^�q���Jy�H��<�^�.��'�xp>��ۚ�>7J;�:؃^���p��FBv�<G}�x-�,�uS�][��'��l�_�ՕD{	�z]Ċ!��������9��^���ȍ�z���kc�Ȧ2�k�w��W�G���݇!�Dr;t�πC���,�ڿV�ۊy����9T1�F@������[~s�q^c���̳����o՞�y��/�< R!��U�a�k0FQ9�X�KSo�O���y=��ۡ8x�Ӯ�w���ҔR��[)�5�����PGZ?f_G/���r����tܦܸj�X��:�
;a��������[��Q/i7�����\����N!��_�\��C3(Y��]�qq/��2N#�a�|�E���g�l/u���\��yP��v�dg���,������^=�֯S�rl��R;���)������?+�Q�bC`:�G?23ޱ;q�*��U!����ۭ�����I�=�5͙Ey<�rȨ�i������n�b<�fk��=ܹ�5��E�C�>���"�%�I�5�[�!s��� �1N}��YRq5���X<,z����Ǹ0�.�v�����j�� �75P�`��o�6�.�.ܒ�u>�>�#�sr����Z�t��z�K�1qk�߿/�o�^� U���P`�����j�r���sc�7W�)ν�^�$v��;>�Nn��^X�}�w���1m\�s۩�l�'��y�%�	���N}�lv�q8G����<�BU�0�vzv����}j�<v���ê��#/�^�o�f�/Ho���cϏ>�lߢM9�E^�C~L��Q��{G�!�_����^b<�"�?^�y�%���.�g~��?v<Ȥ=�48vUzcX=i�g/���}�x;�O�/~�8�_0{�=�ϧ�F�nȅ�H٠'��,�\���D2�t��ON�ˠ���:ޱ˕�
�w$8��z��&�r�8Z��d�f�\LB���Ç_`�o*%�8��Js-��Ye�*������rLܧ���s�ɈtQvbEKyw����[E�U�I�6r�W5#-����S_��
��� J�n$Q
p��n�|���Vp��D��ϣ�'7]�u�w&��#����e�$k�qq�n�f�@�z,Q�&�c�;�m�o����w|vs4�D֝Ʀ��x'}�j�~�O��1O��Ee��Gn�� E�A�HU0&����:�6���|wr)���{��p��T�>؎�L��zyVY�`-T�A��S2����q]��},����lzv˯���EdSy��S����K7��C�a���������%�H�ȡ�ϔ�8�H2T3�P�~�5��bB7��؈���a���Ϝ�0b�f�,�}�lT�:����K��ME�	�N��9)sX�N���9���#ʎ�!<��n�O�w]�cwE�wqPC�7P�}4@���V���1~�\�<�}��Ԫ���o�7�;>�Vzv�hl��Xu��5�Tͪ`�+�>n/�s���^�����G�W�JNR�^hu��La���y^Xϓw�؉��f{��f��.�_ʘdF'= K;�޹7�.��D��ؔ�@BVq���Gb�8w���I����6�t��� ������r��5���^k���Zsh��ѨӼ�.m�,ѽ�*o�0Fs�缺2��_ds-���!��c^��Ħ.�5��,�Bsn�6�[���q.5��qF�����r���(/ݑ�y��_>�̻��>yw&}�B3�L�모��be��BϷNz�h�
_�z�NA�Dߎyg���a�쇰�����E����܊;��)�0*��Hd�^�lK*Ώ�����1`�J~0s� r�mϲb����v9=�`z:��C��5���GV���.�h�g^ʬ�v
�뉮��"�o8M*�1�̔�E�3�TH����;�{g�m��c��גHӴf�}�\2`wd
��Ǖ�W�dZ͍���y�7ii�L��Ffq2��)��6=����/(��Mm��`y��n��,˝Bm߷=j��\g����{��|���fC�����x��܏x-�b�Iج�6�m��E�G7<��y�8wL�ĘK��\�om��xJ��Ϲ��{z��{�>��ޯx-�<���}���{���$�lo���d	�)��G�rm���g.�=~���-����z�~Z����,��o�W�q���r<tV1'( �f|�9�!/UI�K�r��}��7>�
pK�>�f+l�`�l�w�A:eT�/��>�ܞ�*��w�ʬ]:�w2 d�7���^����H�������z��������qt���\�lм�_p�W�Z����B��i�u�8w\�sz�w@[(�˝Jg2�6ku�;V��Ջ������V{�ome�Ϲ����\�>�@�޷p���9���W����쁐j���q1�u�S��ֵy�W����ﴗ�v��t{l�y�̐2=�����j�*y"e�`Г�z}�U��ou�P�:m�Y\B=��9�ps������H�p=��dyހ���S��u���l�t����,��%ݭ��촱M��-�ll5O� ����6��2����\�{]���8��mU{O/E�G�*�}���b�Jȕ[;^�EɎ�~"��A~�/��b/X�쇕�����zyԽ�}]����B�@_�xq��״9È�n���&�'��s�-N �?v�5�7��}���y���[+L�j'����afy�_��o��jΣ��#�m�xw��{��;>�4�c�~��ϭx?*����/m��u0;�T/��pݘ�-���]HX�7+�*�w��@�4z9��o��=:����s���<�'`홽�m�NG�z%��v����7\c�b]��M�w�d�t��Lj��P߬/C��~^y	o�􊏟��¥Ϗ�����ԧ��O=��n�/h�20��+)�z�^�7xfi�P�Wx�:/�Q��FA��>�{\c�鸶���|B�:���'�����\g�e��z�ELz�G�'	85�J2����N�O�gf\���������0:�L�㓔��R�����Jv 2���.�>8�|�bz�^p��Bt�=�Ƕ�����(��%����,~�?L|+xt*\E��@���QM�z�wLds�佂=~�=�޸�ù]�՛��'�$��#�Ea#�ug�k�� G�?is���t��N���hۥ�;�ɬ��)��j/��W���L�O���lVz��Ӕ���H�)W�m��z�����vn�γ%��Gz	̊C>y�a������A���@NtC�r�"FWLϕ_�����2~3�8}K�p�Ϡo�dg�SC��\2;����bCC��Dw��̌��N�z���{`[��w��t�ņ�r�c�Б�FF����1E���6#~Ӟ����������3D~�ߴ���8-
� p�
��Ȟ�5���S�ծ��z�T��؇��Y�lzcY�J��{�{<0z�@{}q�.�U,f��"ih��o�c�E�nN�Eס��5^n^�Yٜ�L�I̹����]d{���������HA�LN�20{n:���ۺ
le�����ɬ=S[2���B.�h/$3�gE��5�f��^����(���2�i�Lɸ�����}�:.+ĕ[C	{��Σ�z��3i�E���m�5[�cP�>p��(	˗�@-�|�W]���m�{���D[� ��][\���r���nz}ٸ�[�匇޹�x���#"Շ�z4��P��A�yS:�Ek,������굇��$<C���d��Ju^!C>��Z���>ܹ����F�^��G�Ո�_�G	ђ�F�z�s�M@и?|{G��_���|��Vǭ$�]�/_��jZ�3
?�"?h�+F}�C� �6"WKϪ�pt�*�he���L˧�����.�'ϲM�A�M��M,V�Ѭ<?&|W�`�</o�2��0?zUp�JT��~�U^X�$�5�T}�'�io��_���$�z�/N�p�,E����9w�~Z�ۀQ��{7g�8��VU���>�d����J�q^c�!��>^�S��Yfm�C00A��r���Vn��,L���~�V��ȯ
n��C��ީ�}�w�e����ʲ̬���L)�Ǜ��fZ#5%��$�}�k�3�-x9�r�½�qG�o=�az������X�����7�E�x�;��~�3�2B�'�+�A��)��~g,��o֦���HF�{��q�s]��x�2j^�����
���'aYR�R��������]ߨW�������c��Y/@��v����`��#5}�/���+�i %z2)��u�K�$�
���E�,V<���Ү9��|�}(аLv���֎: �1���d�u����?���߿m�Tڪ[�2��X���C�1��s��K�����������7ϟ�%���>�-x�;���<��v�)H{�&��@���V3���k�>�n��m���u�7(�^��{�G*L缽�v�hO������ ��h���P����u�X��W�%WW���,o��;��P7�p�;�S��]�D&��=������d�C�nXڙ�����7����za�8�z�J>�ㄎ9K���4�����y�X�޹�c!��2|��ux{\\[+�;&��>��r��2BFLp�]/��8�yJ�FA�솟�ȅ�>�����:�[��: �h�=����z+6�������>b/���7?�>'eV�s�ֲ=:K���7�>]�*r�S������h�u��^ۭX�*�w"��GW��٥�>Ȟ������J�Y<s�39��Ϣ=o����8�^I#Nћ�m��t�x4y\:��&,�1���Ӥ�4=�̧�/�3q���S��C~�e�|F�Vd�=�7����L�2��rY�D���8�tfV[d	����9pƵ�5.�N�� 9�ri;:[̂�r�ؙ6����3Oj+���S��WP@�uO�U4gu�U�^r�|\7I�P�%T��6�]�[�r>d�m������|H�*���hD8Y�N2o��E���G�ق����h��U�;��n:Y2Վ�q5r�!�e��A�\�̘8�ݏ�r�V�q>�Ӷ�]n�Y��K.��u����M\4ij�M+Jz/�l�*��(���t�����9�ס�t�&DdVc��E��Vћ�a��|x*�T0F���Y|�	���ɛD�}t:�kQC��B�\h���e4��O���|�L*�hd���ul
6�tCNu�[��&�է�
��|r,��v+�ή��5�ߡo~ʊ�&�p�k�cf�Oh�g|vj���'Z�A�{j���;Mf.�k��1�� �ھ��F���)Dث�,�Ǖl^��(�/�5|󖽍�%�e^t�r�8���ԩq�(M���u���7\�m��g��_uIU�} ��x�<�Z�&��nJ��}+E���fv����V�Jػ\9�[�e�'���kҬ�vF��铳��>�����O�����EG�7��&VdvR������޾/��C�mv����I����s�Lz�ȶ2��wXD���!-e�}B+35�7T���)XZ�s�0w�9Ժ�
}�������՞�x��`vY�Ki���0֦��@
t�.�U��2�.��UE�ӑj[�ur���d4^3�B'0�t㷕)ʷW���TY����p�7����uS��+�!�j_,tN������mu�Z�t����k�E�ĺ;�'d�A�x�Xq�ʷH�e��gS��Zҡ+'t� ڂ�Ml�/VZ��Q�9����_b���ěV1+��jn�F�t)��Q�r=�z�& ���#'��}��΍�zp��.I۹>�e��y��ܺ!{e��L��:U�\����P��WX.ʤ�K7K�qM�u��˙�'�|V�mow��c7%�7d�d[j[�림51*����V�ۺ�ǝ#�@�k]���e�1ѵ��P��~fv�Һ�}���]�_+����u��oB�gEG2���*�q���NT����ո�5�0Cs{;�_7�P�ee�ک���NӘ�K|�X��Ԃy��,HiIV���ip��.ż���X8�ܼ@-�o�Ke�ل����yZM�R<����f�wNз2TSGY�H�T�](Kj��B��3�Z9��nk���ܮ���STD<�ũ�F���3:F��d��iiU�-��銎��QLL���v��K�J�VN��λ�Ib[._%U��b��&{LX�&��4�۹զ�T�dX��u�嵪ր�4<J��	&�g�Ȳ��mH^�1,��c�Ls}��+�_o�f�!����{4�X�Q��䦅}+����,o��BI/�"�P*�J2˖i�Q�E�u��q��N����Nt*�Q2:
��Ь�KUQgS3�-n됊����ER�yG!�ҕ��'.V"fHEn���Գ���R�ݚ$鉇]wJw]��ddP�z��*�H*���{��dҊ�+�T΢�4���˜"$����$��YDxu�4�C9w2���tqҋMV��v��jm��h��6�f*�$�W\�8�uJTL�A��t�KUZ�eӎr�"7R����Ƚ�(jE�ea��G��+.J���JV	Y��."��y�$����S������V�p��e��yȮY' �)M�̐��j^��ZY�:98J\��¤%=��L�Us"nl̢$Z�2""՚�(+,�MD�QB�J>J/�(`�֞�멌��B��NkuWt����Z'U��ne�d��΍�뜵�xYJ�h�@)��z�ǝ)
pt;�
(�+��CÙc>9^�llA�fC���k����܏x-��,����7Q����YY���ǳ���P��Fz�ꜻ��q���߮������佂=~�ީ�|7�^�^�5��t��ׯY*�;Y�^����FH��H6)���;�N��^�U����go�D�"�tc}�(����c�԰w����CȜ�������jB^��5M��r��T��1n6F�Z�W�k�w�5>��:v=�0��������[�Y9A3�@�M�b�ѹ����!����ޒ�)j���.
���������`��� d{�'o�_�*�PT�D�cמ�u�$���XՇ؇����}����)��棘�EG4�����Z��>�r������J�� <�z���xϾYშMFZ9齅��66���\��z�|�^@xO�S;�"J��k2�۠N��vͮ[��������5p*���[7n�;��E�v�/�q����,G�~�X:���=��ŏ}ʌI����`���چr&���|q3��؂o�w������FDW10I��z��WԠq���W	繶�`���_a�&���P9���QŇa�C�V����tne�8���w}QT�xowjMJ0���Ck�)��z��ʽ�9J`t��*_.?(�_'ع�rU�ma�Ӵv_5*u9��Ϯ��7sG>�׳ssۭ,��k&��1^��-�D����L�%��y!�;<�.V��m�*���gּ}�y4FGm\�eT��S�"B�
J�C���̔�a5e)�Fz*�����A�N�o��=;��]WD?\/:���2NQ���鐞f�����OU��nA�]�y�{�Yلo�{�1�U�^w���`{�esay�%�;��=�CB�Q��J�����2��F:p�ؚ�+_��3��η�^�����	�����S��W��G���v�w�9Ɯ����w>+��
��/��m���W/=cӗ~�N��:Q4z�}�'�aڞ���Ǳ�x�°��Gn�ϰ0��g��×j�V�N׼-FX� b�&<�����;�s���gO���lw�e���ψج��ϧ(!p��
�C�rʥ� �y�ӻ��Қ�<�B�D&n�=~��7�᰽��\��T'o�v�d�
���Q�p����s��\��g2��S��=FA���.
��"���Hl[����fFD{�'M�΁)�F�cݒG�_��,	]u{��JK﹑t���J�sУ�ܑ�R�;�*�(\�M�����kJ�&�ik�&�W]u>��E�LdJ�[�	���G��C�U��T&n�C�Uˢ>q�\�6�y�tm���^����;c�|+�mT��z����SvdN�C�h\O�؍��9�
�ތ󡙍��-�� ������UA:��}&���n��ʷO�9
}��ʓ[3�G���hrŇ<�Md���{�x<7����q�4��P���ih��g=c{�,�w��>�]1����rwwu�r�n�����>�yf\�/;��z�2}�C͙��캐� �N�23��R��]yN��g�&�W�y^�7�s�g��:߯,>�L�_?g��X*w��H�������e��{K�[�;�h�O�j��b��|������a��������}s>�^9Q\}�r�����ﮕr��O���Ɣ�kҲ'��¶���t�6��z�ǔ;��������e��/�����D�XԷ�g���c��1Z1~�ò*�;q?���Sr�_?��+��ߺ~ Z�ս���{�zV�����e��w�zDo������S���Q
p���ǧ37~��'��5Ǟ�{GZ�/����lw�Z�C��U��0<dB�������vB�2��m��!����΢#xq��u�V+NՌӕ���wr�e0���֨.���\�K���M��3�F�;���1.<�q#�bK$�G$C���Gǥ×�bwk��*��0j�F8Õ�J�+{�VA��0�,NM���\8�M���qo+�ټ9%�~V?B�s)��{2a�{��������b�Iج�6��M�����y�1�4�uig<�xQ��YV�ye@c[���C���w�|lw����v�̡lĬE�Vm�=w��V$m��Hg�n"I�L�vZA���]xe��ෞ᰽S����K�������sy�ܵ�-8�GV1쑒<-@�j�9�=#8RAJ7]����G�ئ ���1�֕BG;�c�:�t�m������9������L�Hz���	�5^CT���~&�tU��������dws�ӎu����:���(!����*)z̓m>�p7|3Gn�H�Z�Cw�\+�|r�� �{��O�_��~)'=M-8?d!��\���sz�|h�G�6��M�X��xu���||�Ŷo�17~��_�g��'�Аt��#r.c̞>C{N{ ِ�kf���=C�m��22�d{}�c>}^�a��3ޮ��얱aR�\�_O�v�3�\�=z��|��?A-�^��܇�睐��bh�9*�I��3�~ݻ(;m)G�)�ӵ�h���QW�\�yGF[&��9��u�M^H�#�Qc0���h�b]A9�K�7�r�wEWݽGa� �z��e(f��Q���jb���iT��ܡʲQ�ZV�\��F�]-0c.R�v��:�]}_���YΎ����B����1kA�/ߎʷDD۟^o�Ś��r�Q���T}>�l���׃��׳��X3�.��?m^$+Fv�Ac���-,(��	$
ӌ�\�LϾ���Nÿ[��Z�?U�p�/}�R����
��YP"p�o�WA�	wGy�J{�{n��>{��37���S�)��6=���0���i����lR�~QU݀��M����������=��2�A�Q-�5뇜=~"����܏x/Z��w7=N�ș�_F�����ީ���
l����C����])9UH���f}^����z%���&Yn׷����߸���ވ�Z!�^� �
s5<��8�Һ�0��M���B�Xt��(���M�Uk�s���9��c��C:+��ϕ�s1)z�vSn�'&���Vf����CT�h�o��SR=�^��>�0��tr��D௝�����u��g��OGC�����|�R7�l!k��#���3��,S������d���	���
�T'KeH��Y��:߲�Q��e�^��~�(�y�m���/l�b1��"�oZ�f���gD嚼Y˯*���N�N^8%���l��w2��KH��,4Uu�5T�w����B�{!�K��&�BIT��.�Mx0��J�{k႟C:�JI�����_S6gא|棐\и9	�������ۑ�w�7w.������^�Q�]��f
�2�©�:��e�g���c�5O�";�\�Y��?W��ޤ<��WXO��ֺ{�w6�d�5U>A�R{$�M����W�/K�F|_�<(F��þ�Gq���N�,G��^�z$�a��A�@)`�v���k�#���������aWQ���#���}���%w��u~��y���ͅ���ì�h:�����C95�!vL�V���1C��߂e,C���)K;�8�������Bw~CY��V��Mp�m\�B��N�u0;7�T�^�j���|U�r�k�c�wϪ�A4U����K��s�P�p��c�.;#��}W�͑{���%�{���A�4o����:�pos8h�!��N&�W�zw�t�<��`�ط7�s��s���5�c�R~��1�����TO��Y2�_�F|m������Y=~��ӾZ����Nd�_+'�ܟe�����}�9�B.4���>2�dQs�~���J?�+U��S�?b8�s+2�g���3��w����~P�F��u,=}-7!ՀbCl�c��Uu��ȷ����MJZV-��C��٭��(�4T� �o�"$���m��E�7u+��ivX(n}��ф�¤����2h����w}��a%R6
=�Y�p6�NDo������u��A�#0 ��V洲�'�g�Wbhvyj�Ͳ��5ٕ|�ۓ_��;ފ��lw�e�~�> X��7@�!�5�����Z=��\Wo��}oeXly��W���x�^Sy���z�_�Bv�ە������v/���~_�i��������	n�#~"���n
��"���Ho���";���8�P�܌��Sc�y����g�s��sh�zL����N"�}���>b��5pS��"��)���W�;�޻�<7=�=Wp��۬b��UAz�]Cy&��S�V�1N|&�(;�]7�������3}S��qLg���G�X|�P^~h:��u���]��^�����uq�'ںx�K�3���I�������yW�l9�~y�3P��R.!S �H�GT�a ���k�����G��؈�9I�|n6O/n9��yc>}�w���3���n9�ԋ<��)�Ʀ���(�g����0uB�k;���<CJ�FA��+��7�����:Z�b�x�"j��Awa����O����h��0 �2��n�lT)t�geu\5v�;B�ޤї��&�g1�+���z�2�*���
�C�x�i�\ĕ,`inf�g5d���c��Tflg�g4��!��R�����<��C�)����͂���xn������M=��k]�H�R�gb�"0����Io��,x�Nn�*�~��Q��{G��_����x:�L/X6�����o�jݟ$3U�V�?^�?1Z1	�:K��gɹg���	���T�v|'�7|I�uoU{3>�o��e�a���W�:7�u� �v
��!I�U�Yޙ| S��r��S���I�A����"S~�H~����yjIj3��F���ァhJ+�+���c�5�^���3ލ�FǾ���|���a���`��u�;a��>^�S��Yfo�Gn���*/ؽ#o3r��-i�`G��x\
WU��YP���4=~�ީ�}��C�O/%u7�=��;W_�"x����F �2 ��D�ڙ�촇�~g.�+ި[�p�^��d:��7�<���/W�v��礍�#����H�\(>R�U�
Q��~�7ݾ��-�u����F���Lz5s�G�'G(�����ߖPA�̥�=bj(6hN�!�\���U�$	�.T�����-��d�J��y�ӎv���:��(!��l}�a�Vdx�6�[J�x� ��jp�N�j�C���mk�����,�ZnY�1��Zl�{�%�-z��e �J���&p|��Z�[�e+zg��E�e�)vo=��b��@ b���&+/6�WR�m�����z�Z��vp�;�!Z�#)r:��������Q!��k9SӐW��w���=,�4�eL٨�k��\��ȳi^����?�~W8z�+좱XՔ�!���1qpٿXȄ��G����f{��d�=�aMR���"z(����a��@<=V���ᝎ�^ca�da~�l5wᏫ��{���ų~?�Ol�}���-�v���+����3�\�=z���(���^��܇��Z��5���}׫��b�IŻƠw��(��V�������Ѳ����ӿ,v�6n��	Ι�:/���A=��wѧ2������j��u��/e������T/\���}������91��4<-Z���=37�Y�ߡ߭����6W�;�lZ��������O��շ���j9��ފ�=��n�zץ��陸���ה��ˇ�yWO��q�R�Q���]/օ�mwXH�meM��,�f�S^K�e_�o�v|ǳ�/���kˆ���G�����~�%��:�U����:�Jf,�`hr�i��6�K�lmq����zV����cѣ@<�'�\�ݥ��G�Qk�
1A��%�^����=Y"*�����K����j���={)�<�����n��oH9{F��J�mk�cR����n�ΩK�:���Yt��:&͹i��s�6�M	�>ڎ����+�� *�2���T]�욫�V��Gs����G���ߣ��<tVqd�A��LH�r �N.˦�5����U���Wl�h�gg�߾�qɝ������K��!��X�<����>R�J^���Ϣd�3T�h�ޞ�����;^'.}O�f�)�gN�}~aq���caڸ9�S1>Yoɢ}�r(N^�o�:\{�S��1�4=�\3��F|=�t=�0{��2@������ܾ;Sb%:6�<����]�;�$	��9��sQ�(��O��Q�xo��nA��O�^[��p��/�ܴ~ٟ�Y�HL��U�Bk-~�M�,�����}�.&��.+D�{�m���y%~�=�><��yp���*���$N�U���a�����~"��@o(NmL#���[�х�ٝ�8z��{�^�c��'��n_�\<�f�Y��enM[mZ�r��
��F�W���rÞ\/�9�ft��oّ��r]�����=�����9P��Wz�mn��>��=���7�k;��(ώ���I�������ϯҶ<qY��n���o~��s��Է�mV�>Ĵ��pb��ݖe��]�$a����Uj�[V~�S����(���pܘ|��Ǧo6F>��g�l��9���\D+��W��H��뺵�o�ֶT�1M��{�\o.�A[|��f9Xsq�E�]�#�<[:�M��1�,�Z͝�,���(�=x���qX�\x�Hq�,K9�9w�qT؀�y���\L��%.#*v��]��!0ky�u��G,�!X�G��;xp��Z�૚�9��T��@���ͮ޽B�8�J6ُcx_}�m����9Dd�z��Akf�;��m<TY���[��Ϯ�N�r�u��^v6�gn�k|��jS�����](�Ǔ�'�R�>oh�i�Ǜ���7ȍ��ɾ�(L���J�
���G�k�Ð�Tq�3У9Խб�k �N��Y".���#s���ۀf��0�����+UEe��-�--o ��'6e�&�P��(��j���W4Xv ���C���7�r�-`��JѾm�(��vu���G8A�V�at5�a�ćY��U�o�q"m��mly����kL�/k�&���t�[��ב�=@�5Ùͅ8eݦs����4�tle��X��A�34ݣ��&���bX� �.�[��x�ȗP����Ʀ�M4�1�����)�(�U�k�ക�Y������|tN���v�.hT���$�N��Y�
�z"x��5��k(+n�k������d��v�,f�H.xt+a7y$�KK�Y�앏�Ӗ�����K�]���}I�FdS�9 7�/Nov�n.l�f�eݖ�����;�x��������
�Z��L(�Գ9�!\U�T�̦'"�lEL����ۄUE��tso����#E�v�)�:�Ps��A �sfqj�&%1�WfjK��۱��|�C{�1sx��xG����źJ,�[����d���|�̬�f^�s-u7!����,9j�%�S(�]��0��]5]\�UG��qY���`��1d��/Qi�A�3�e���(e����q!�c���r�νȨ�`���d�O�R�}��O�
��h�'c��gy>�wYx77�r�pfe$����[:
T�qf��}���Q\�p�Vv������w�bUƥcTwil���<�,#m�`=#%��)�wS��\��zJ�'i������zZ*��K&��9Y��������b� ��o�'-[�O�$��I�$�~�O����8Qc#�ٝ�Ǖ�����;������.�狁����d���@*��J�p͗�I��ӫV�^��ҽpr����U��@�i{����r�÷�z�˼�%t�5��+�\jF�
T��t9U��s��x�6�����ފ��]��c�lR"�J�\�b�ru���v��J�
J�E�c�Q1�l�k�V�Vp!���N�}�|D���iK�f9j��� ]�4�D�.\KA�.���ĝĉ2u��'"#�l=s�Y��Ҋ�L��eDd���V!,��:ΖK*�V�k�AW*�jW$�YZ��YH��E&D��u���w]�t�J��ι��\��"2����3	Ԍ��D�]s��w7#�'3���=O7&z��S�֨a�f[��(���+�T^��	c�aGs<³���D��''(�-�<�T;�ȯ2���s�A�'��:�S��P���.�̪�i"���Naf$��@W �<�L�����r��©4Ē�rt��n��^�G�z�{�:��kH�vdEz$Nc�z��*ʤ�&��(�(,�
�wv����r�H��E�W��b�Z	SN��ҍH�����|��O�'p�\���]C�z�h^�v�ƘΉc�V�y@g�_ps��G#G���c��^U�R�@���*0���FV�`��w�d�%Y��0j��7�z{|�ҝ����~�^u�yq�9�/=�sVk,�o�O��m�t�p�X6����4]/ ��U8��W�zv���q���{�=��^{�˽[��l�RB�~a �'��5|O��/��g�*�_���1~`v����'�+�N�׫��4MnUw�G�M�ﲽ�]����B.#N�p�>7���Qr]��^�T{�Ǟ����e�X����TVwxΓW+�=~�:���S���l{.=��������G����{ΦG{پ�'��<���˵f���{!�ܘ����؎�W�;{�2����b
��h�A�]y^��U%�� �P�g]ߠ�?�3��{<r,7~�~^�0v;�2��s�"���x��RR�}����o<�=# ���]:����E/��9�\R���Ho���"6��2z�9�>��R��J۲�1��Bv+��c�G��?1?�t�*#ߏOsP��-ו57��������]���^/�z�����-�� ^�.���6&���T��k��oMM��s^������Kw����v"��@��Ƈo��H#!�FAp>1՜w�nu�C�-β�R�r���~��I5vح��|k��aT7�K :�oQC�6�W5�ܵ�G�2���rZ[�͖d���WBm\5�7O:x@ɬ�]Ζ��=5v'���5��\ܸ�^��{�ʓ�{�=1��X<'�z�bk�O��^����푐lM�И��g�L��I���lv��Gz���T�}�wray߀���w��fW��G�0'\C����xi�~��z@yp덞R�7�r:n9{q��߯,>�L�~�=>�G.N���MkN����M��g����č�F|:�_����ae4<�%^#gd��	�\ϭWj�p�5R�\s�X7˺�z+=�s!�f�!�m)�D�t����N+�@Ἡ��q�ر=�Ɏq��t�N{R�(/G�dWg߯x]q�x�x7��:Ń��nY�(��g�30�f���O����}������[�zG���/����_���0;�TeH�
r���������C��̧�^���_�N&�������ז���j+;.�f�nx9��Ϫw���^�{Ьz;��}j��̷��ɇ�=����v�_��cي}'k,˹���gM�v�1{�n������q�9V�{am�b���!�!����S��{���EJ��?�f~5�B��#V��(�@���k͹V�����J㸆�'aJ�Q<�QW��<F�հ��_:'�c$Ѧ2d�)�<e�fV��L��NL��6f�D�)P��V�l��v�e���̴S�%6�+��N5)-�T'.��83�}�,�YT�
=�n���[��tyi���,ϲ$`��9 L���3�����3�^�^Mao<F��QD��{���u�{t�zl=԰s|���<�!�g�C�
���*�>�e�f��R�F���\߾7ا���[#�'Gz=끷�bD�L�\=bD�hK���{�^��#�xϋ4��i��!FV}�إN�{��i�%���Q�\~�;��q�%�W귤�>�fy9�gx��r[�:�yM5�s[Rg>O������l�2<�f]����>����Ӟ��+Ŧ���ENx`�Q��z���lֲ��a������R=�>�L�{�*���:��?՞��=��ۯP��^ ̀�Ыgi�3g��^�A���~��e��^r7�����;�X{���=���X�܍̟o�2o�=�B�U*�����O�e��A���g����}�����_S��`����^�k1�E����9��/`�����N�5����*��:lhn.��)�V�7Ly V�r�/ǳ:};	ߖ�{��x>�9{77�u�80;�T/C�~�]ػq7o��ϻe. ��{2�Ol����o�:�H��)��%޺l�I����*�&(�7�W�ۯ��Ӓ�e<a��k�y�7�ԧ�����3 !�ćb�ml�s����3��%:�-Ǫ�6���ëL�tUh��r�x��䊎e��=�����g�/�dv�,s3q�Y�u��)C���W=��h���up�+�(�K�V>--v{���F���q셝�F��x���37���R�?z���WW�yڕ�{������b�=}�C(/e0�U{E�7߮�q�q>cMz�_O��&��Ξ�ok؈=�:e�ţѤ�x�3�z_STG��I��%��	h��W����t�G?^Kq��rb��-j�4z�}�3�P:��c��drE!�c� �
s5<��j��)���o}���
�ۻeJ���}W7����'��s����>~y;������� ��3���z`���/Mv��Ӫ�*�U3u����f�7��0���D\�>
Fv�}9A3��wB��s��̐�g� a�^��r��Ee{�T�{~@��� {�N{��̼^�M��A���+�k�mP5쏤L��:QMّ����s��?[a�V��ttE��qt�%Ӷԏ|�{3~�b��S)����hM}���o~Ym�%�~����~"���5=�/ۗ������"�Ǘ[t�X&��u�@eH�p�w���S{uA�>��dJ!0�Bnɚ�P�β��G���3z��B�^�T�1'o7v*�������<��2Ҩy�q�rwS���)vmu�g.�1cr8K=��g�<��:?Rx��G�?�Uy��O� 돎�R��c��v|.v;�-�s�kM�#Kҗn�=U'��2�g���,{��=�Y2�װP0��C9�״G���T�e����+�\M���>���{�7�9�t����s���.�?UMqW�s�*�o�Ln�{�mB�5;�̔N�*�4X�
w�9ey$����gg�a;�!�ϯ�k~�͚#�*{���я;.F{ZR�ޕΥz!R�$l��Ȋ��!��@Ἡ�a�Y�uU�uI��y֦�wf��T�o��k{z+=�塔0�HѦ ==]/*�0��]/ ��S���~��&%�z6��(���h���n^` zW}�pI��z%��#�/�#�	h뭷�Ή�~c�����I;�͂�5ǳ�=�u��o��7�e���<Y�B/N�p�,�Nv��D9>���^�v�xf2�!ԓXW�`٣+�G�%�p��D����矫��-O���"�ۤ200�</!�e�j���<���M�������}m���H�{"=ɇ�{�ӽ�xv�z�Yȇ�s�7��wD�ߎ�E�_~ouM�V輢�:�2�[B�R��-"����4�J�sh�W�涎��3hm;s_#\����i�*�-��@�:�R�S\������u�I�n�t5�L'�7���aB����SG���5����ҕ�zP�g5fdL�ܽ�7�)&�aV"o<(d��15�J�3�-�ٻ��_{<r/)���>uϽs,�נ��W��N7Ie�V�$����&��2�(�S5��)�٫�A[�ȡ�ZA�?��F�[=y繧��cНO�����[p��!8
U�z��7fFO��9�ڛ���HsK8�����������6�q��G���wlT�ʨ/V�o$ؚ����*�vy�Ψ~�8Z�l��K�F�
W�����k=.g�V<�լꌉ�v�mS ��B�)�gz��s6�.��ґv�u7}c�����ϙ�ʟND{�2���o����{^l��?eԁy�������괈·Nz��H�~�_�l�#�9^`���!��_�=;���,>�L�P���>[�mԺ���׃�X�ʷ�>�۩� �F�#"V��9�$�J�F��z���>���+��7ۚ��:�'ɼ�9Q]����Cڭ��xNVD�t��������� �&���٥J�ʐ*�sgkMQ�F�:��
{޻^��+�~��l~b�b\��}=],UFpr�>������A:�6�S�t"6��E�y�PЛ[�W�<�D/��}�՚<z��e��R����:u��=�d�������ļv�/f�5�Q�7#U���[�i0%���0�G�Y;��@���v6%V����Hbo�ȫs�0���-��i�����.��o�zfT;~�H߽��~��t�����k&QU�͟�<��8l�磟�%�Eϻ=x���s>{/�z�k§a��zF�{/��)�������8;]�V�[�Na����_�_�Q#E;�dY�0㹖� �fL=��`��Oޣ�O��f)��� ]FQ'�o�r��{�z����VFQ '�h�p�U���[w4�G7�`�_�w��=�$c��y�_��v磎W�����*&�[
� uNf�����ǧ~g.�2/޼�ٱflC�T|7#�Ir<���xǾ�S��7�R�ȍ��fE���2B
ϕ�)�K�×֒����}�nVsG�G�Sy�{ا�S�cC������tz�Y9A���J�z��d/�����y���,t'�:��wxQ�������9�a�O'�$����_�*�
2���Sp�˹����^H�{��_W��+�3�\��ԙ�����z���l�3ζU?�-�k<ё����l>������R�ȀhMF_�zƬ������A�"Y����H�w�n��기�N���f��pns9f���\���cB��7tc��
������/
�\�K�����
t�L�cR=c��;	�f����gq�\�f8'�b;.Ph��
a��dGj�%˽��YW�x��8��:��tL`�o`G���-�݃?p_�p/��E>^'C�){�ln�8f��xu��2��{s�n��.2�w;;����M��Ǣ8�`X�{�2|�Ҽ��$g�kÍ����(������M�nF�P,���~u�	��h��샱������E�������џp`z�'jȞ��W�w�}I�s���
��>��T��A6����ΟN�~[��>	�^M�ٹ����Fp`wEv�a;ŷ9Yg-B[�]����\�{>��Dh�fGr�L����N���)�����F�v��E���;������av�z�yQ�D{��j��.��{��37���:�Cc�q���g5yI�3�R?�n~*���ߦ�����s�<Q�Xsٖ���\������Ӿz����s��nK�}r֮;��eF��6� �U)� e���ӝ��tŌS^�F\���~p�#{s�O���#7�>���{�l{G��#�@�3	�9�� ��~�6�ڳMEq�Dx��!�=y7��=&t�=n{{�,��㢳�NPB�C�㋋q�]� lzd�.������ګT$ז��=�φ�Ӗ�h�x�kF�Fm�V)�������O�J�mR�
?��6�?�ݖH,���s �A�;j�Iȅ� �Jp���+)I2ń���cھ��jF���ՕfɮC�Ŝ�	���}rR�[j�˷�3�*�Ъ��3u������߳�{k��N��z���B?V:V��Vo�b�x�=LO��S3>�4�/�j9��+"+�Z�~�����~�$��������pi��|�xO{�sV����H�l\P��)�22����G ����O�؝�#2A5����^������.������:�*�T��t����?Z��[`��[��6��j]>úh�7ٚ=ﴜV3ޯ <6�|�y�<W�B���e*��9������bdt��哓��{ޕ�Vx�h�/�S�y]؅��=�{���{3_�
�`�چ}�h�>�i$;���G�������8��{�7�9�y�.v�e�>�˺[��6�s�����6��q_{7O��{����=P��B5k;����I_�����>N��k>�M��͚"�̸1����;�`fwDa�}>�{n�r!׀눑��0w\<���!�.���*~�g��W��8�<�gwV����y���KV��G���u}�m��YUC�5P��m��.��-w�x�K�7���߀�~����6`��O�T�:.�eG|���4ĺ�싥��w�}�ՉH0"=�by-Eַ�Q�S��#%B�j9�Ĳy��Y�լdZ�,=��Rxhv�yx�u��c��7��7h+���+Rb̭[.�x��x&�M�䄕q3%v<����=��]�LzƱ��B[��ȝ����h��>��L�U~BZοW�mM�ב�ý>]���g}$׍+�y�_�'O�����]���XDgeV�``yHs��UMʼ�y�hyu��#����.Շn�/��r�p��D�k�[�����߽���E���!y�߻�Uvc��yj�`|*1��J������[��=ɇ�{�ӽ�xv��e��s�.h:C�N�z�<Fz�}9A$ ��&�y[�Ö�d.y�G��"�)����|����|�A:-4u?~�|�t��6�vН�]�Y� �:��*�u3A��"�b���ſ,�>ސ�W��žռ�xo�Ǡ*�	�T�9�X��U�W򪐃�R��bCtdo�S�s����Z�sk��/J[������J�����6�c��G��ۇv�J /TІԛ5�v�VE��ٝ{���'|��ϖ(�O�����k=.w��,=Z�~�Ȟv�n!S�_D_��*'�����`�-�A�4�E�66�]VJ�|�Թ0��M����'�}_�;�*���`���[����������h��cm�6��`�1����6��ݰ�����cm������6�o�0l���`�����cm6m��o�0l������6m����cm�6��0l�6m��b��L��q�qd/� � ��� � fO� ē3�z@�@ R�D(Rj�(+A�l����BT� 6�J@E[iE%J�h�VU@ P��@ԍ)F�Z֕V3B���z�;��6ɶ�Rһ���ʛb�LDkX��ԛm�6��5�;whĵ�mi���W��Q�V٢�k*(E5mQt�����d�l�[ZEhŶ�Y�#���6Օ���5kd���ͪ�m��-5m��Z�jBX��Ii�R�6�f�LkTB��6�m��%���![j�eH   mS���A��0�fk�ۻ 뮭ض��nӾ��=;��ν����=ƶ�t��Ӈ��%U��7r����;�����Z�ݽ
�X�[a��/:�M�SMBKX�kFf�F��  ��W�5�ǳ�F���N�o{Q�y[��j_4oz��4  �(�D�th   :(Ѡ( ���xF�  �q��   @�>��=4P zԳS
�
�}9J��՘�  ��� 4�{>��+���S�����\��[�8�[wk���q���qb�f�޷���ՠ��s�wA-��k��]GU�Lke�FU�V��^��|  �>}5�m���5֔���{������E�ꢽҋj�ʷ���^�Svov����i�U�w�\���h[]'n��N�oJSl������lYݻm�ơ|  z���M�ۦ�u:�5��6��e:��^�j��{4q�9ݱv�.s�����{�-j�i������kn��٫��ql]���ݲ<v�R��8��ݭ���[[64�ec[K�  ;��Ѷۭ�]�)�i���t{������WuS�u�f�[*p���]�aqʎ�n��Gwk��ӻ��U�[�[��;��ޯp;�m��m��{�w6����5�v�ն�Z��m��IMz⫬7�  q��Mtmv��-w\��Z�-B��ݗ;�_1�����l�����v݀6�����+^���yo]�����w+c�!���q���mӎ۷oN���[�����ٳ2-�
m�mVV>    ���v�jڪO]�cۻ��:)pk�������x��:��:��m�]k��h/<��{���!h���(��mwlݺV�����wz�m��syO]eK�'z�H6�-�V�5[cU�c�    a����.:wvgm���۶�+�:m�+�w�w=ӷn�j�u+�۷h껵ezk���n���^���e���^׻��T�\�ݺz��l����cmK�{Z�S%h�jB���̆�   ���mU�jUo��oI�n�=7��)׺�^=�\md�-�vНJ��=��{�9���==v�ƍV�l{��RQW2�Ni=b^���a��v��C��T��&ʤ��4���
RT��  ��4�T�S�MM��0�~%R@   �?$�*�    I���*���F�2������?��v-/W�V[�߮����`�\:�-���b��ټ������_����$�!�����$ I$�	'�� IJB@
 �?������i��柠cB���i�h]�)6ݒw5��!e���w^��R۔w4Az�Io��1T�=,�'o7F�W��+�h[��.�;��Rf)boM �S�,Ō�����j����{E?��[�`ך-�V���p�)��`ڠ�B�9"�h���x�A����Y�&*W�DG6���[��Uj���p'z153�:�R�w�����C*�B�Ԩ.�A�v��7f f�W�r�k�!�oc��Z�{���*�Ȗ��q��Z���n�u�>͘!"RV��)*f��7�ڃT�5�5��oqnGx �5�]M��©.Gn�&�F4l�vl7l�̼t,�7@�B��%��.��[���BF��٤�GY�K� Y�-B�t�(t�^Y-�;%:A�RTئ=J�k���Ff�7-��/~8�iM#l�{&n;:�Q�-��O!�B�V��G�!7[L��#� ���Q�T����X�o�Lm�v���-��8Qz��O��כh$�!�ܕ���{(����ɦ[rôwR�P�oh����l2��0e%|I��0��@���xƢ���-�yb�V	��2�&miv�˄��$j��f��B��ulQ�n^P���-ʻzG�Tz������v.�醚�ڕw�.^`.�<n�w����JE<�ՇW���.������.�[�$Y�Z4�ZC)+8�[���ȱԌ"�RX@e�7d��xt��m����\�?�4QW����LX�s'R�F%�\)��Sؑ��jkJ��;�uj�KBKk�2QiM�*���&
���ĲQ�xh�ԑ$�ȋyN��3YX���A�5���h�D�&?��mdWk/gpۤ���,�y}|뮲*�B�b-mF;ۻ)D y@�as2�ѳ.��{�SKI�|Iݤ����A�L���OQ���lUQ�/A�h�k%��-c������.e1��mn���3-Z�ֆ�w!�k�:�ш�.B"�(ˆ�C���j]ܬ��:��Yt���1}Z�꠆�g���b�sGL-=���2}mZ�c*�ų[�	��!�� )V��8���σ{N�.%j�wt��6�Ve��ݰL܎V%m첎����)ݝ�ab�q6k��l�a>6Z�]k9f�{�Y�x��=\9�me�����gκ�t6���;��ѩ.�����B�ׇ/.$/�����e[v�R��[���M�u.�[�E��4�ڷ�en�����q;�/4�R���[��^�v�Z��	����!z�#rX���)��t�/M�-P�9ѷ�EK�pD*R
\�3�CAW���nĉw7f��Pae	f�KE�x���^�QE5��x��Lm����Y�8H�.����+$�5j�Q���`aZ��'ϭ�*��=�#�l�X��Z\�F`�e�=�fe�SSd�յd�&柋�t&M�X�2Gzs�.�LaJ��}w���p�U���T+��ʙ=D ��|q��èo=4��\���!�ۧ���.ō�m��i�Y�՚���ei]�(������i�6ŵ��.N�&
�W��!�����3omAux�J�wR�(�����A�����[�#,�|�"�ܨ�ޘ�Tm�u�+V�6��[Wx�ཬ/��Z��8�tƫ��,�[�%�ɒ�j�� 7��A,ݧ�@��m����Sj6wC�Vi�1FHc�2cg*��0Mժ�k3)*��e�r��3L�w�h�*��m[Y�����f�i9 �E�Gi��L�%�0ӱK�1]�n�.�N�|n˒^�͙�m��h�n�غ'SFj�'x�-������q7j,�/3(���j�����րq˥�Vmǂ٣W��0�.wo_+#YI3L].�6F�!Gn-l"�o�,$�ȕf�շn��ǖA��&l�Ю|�F��ق�tj(N0�ș�^#���A3�D;�(�Y�eb�CT9vr;�\�t Էf^�^0f|S�U���drh𥇕@=#s(UqH�oE۽KL���ɻ�䩤i֍^����XЂ,���-�Ѫc���ۇc��Rɡʣz�8e,j�,`�xv�8���٠V�죗B�/LO^歚~l����#�%���/n�֐��:��6[����7ӥ��5ޙKr�d��z��k6�M��p5s��ѥZ��ӵŰ/�^��$j�j�E�˧�H�<�+R41Kw4�(�4>t�&�Hu�DB�/0벝i���Tq!Y�k����;R��{�ū��Y��X	���Xu�M�e1���X��]��!�z��zq�OqmVnZN��Q"�͓ �sB�ڇ��7B�xR4j�b�D�[��k^���4tq��Y���)��B��O0�|i0Msr�M�v��g��6���T�V���w�v�0�Y�ST��T�7%�X��]�Jm��s$�In�o ��յ��2�Z[�}4buq-Oe
�&�2d�F��:7�^�(��ˎ�J�+h�;>r7�M�B�V��h��3.���]8�D����d���M�I��ihOF� ��ф�.�ҥ���ԸA8h��]��̻�T
`ӻ)��9v�칰)We���l�FkX�4]����2�#B�b�w uY���|�i�|��)_,th���z�����H^�$=ZM=�x�i�|J���[���*����c˱b=�(M���B�n���]�u�n�u����(2�eF�Ѫ��6�&L5y��-���v�����	Z�my�D3��h�Z����
��W0ۭe��b��^�\Az����k���DsU�U�e��x��ẘ����[h��wu�Q�4Y��7Nmݳ*�P�l;��$<��s
����5t�����-�?�0�&���Q*�pe��I��Gb��1V6� ����K&��۽M�`��F>X��G^��k�zq"���p<�WX�(�ek������w5'��D�K;�`3`����x��n��"��M���%6�b�v7\h�w[eg"�@��m�eL�s���)�A4h4>VA:��;T��ijw��f�0@�8w[J�c�ң���াw:k0x;�٨-�v`���cܲ
v��;6c�q�V��qeH(3cak1j�$vaPk�2���N�,;Y�K��(�+kdF�,�ki��I�kL�[/>��0������jj�@@�"����څ�[����h*�w�$(5��f��¥]���j�§M��J�8�?��DY�]���9�kL�lu�����1������ulWXtC�(U��l��*勅��Ff�sr۩��w���,f̹@�zц��Z��2;�����5-�7��M�F�����̬n�t�@ +l9Y��*��N��SJ����V�h�@=�+�em$�5�bz��c
�%`i������w[���ʱ*��im(�ր��l2��gv����3f��QD��-��Ce�4�!��ax�@$�˵� �N-�6aد*�a���b�m]]7H��A���e*��ޚ�R�n@w[�Y�JV��棘[�3��I0��k<��̲��r�pV7��᯳z�,�m���,�p�@�-FkxK�
�SM�L�:��Ǎ��E,úSx��&$΁R%Ql9WMPW�+P��t�\�-�5Q�0 I����Ÿ�L����fX�g.�I����\��i�	��0=��.����v�ۚ�8f������d�b��6,�jI�e������ު�6)Y�l� E*���\�������IgynXI�41^獐Gv�/��X�e��`�-|^���F^�6���ff�tj�|s�&���[!uwz��gU�F�s���rC�Ae���c��r|�:. y+4��LἼ:k�*f���c�$�� 0},����b��XZ%XQ�[�)���5�BݹY�r���֫u��k!5zqVk�F�'A�4FK�Ҹi�����^���/={5����ذ�Z���oc=���Ք`07��kn�P�`ۣz1�ѵ
��ȪdSh�%�JZ/[&��D�V��)�6Ly&M����ۤJ�=�+\8
���Lf�g�ChG�]��2�^�Vf�jb[�ęzH©����:D36�m��]�y�t�����f<T��������vc{/V6�#*�v�r�`��2�	ѩ�LyG\��R��7��>}l�j��l<���w�io2��h)#��oX�4��r�3	�
�7f��M�
-�Ӽyi_
뢋d��O5��x+)=K-F�!i���-RH�����6����]1E��P�ى&�D%&�Y���H��6��&ݥ��h�7��W����Y�(��vc� �׹M���u�l�J�koҙ|��@n�`p�U֨��IF�i� �]���:�ʫ}��0��էs�ífZ�2P�p��h���b�Fhm�W�8������wu�A��H��� w3u��FM��[X�[U�yA��n-��ٛgH���ԧi�w��c�L�ӵ���	\�R�'p�X�u�勴R�eY�6*�n�f�����[�
��u����Sa�&�y�w��e�(�4m^� ��Q�6��<�v!���6{Y5� i/�-����sM�6CX�p��q7�af�k7m�3��.�mY =�D��JX����mw�r����m��7�k�hQu�پ#R�:Քm��:�W���m���J`s)�Jl������J��y��wXH��-��m,{��?p�^���h�PP�djz��`c�ncۦ�V5���f�!K'n�p�1[�������e�Y�vMn�T�֑��pWu�:�q]�:�˶BI`m�O�z7�����DQU����/���St�:t,=�k5�- �R�3��/=����NX���]��Ve�̰�Bih�p�	MDB�֙o1ڭ�+^]]_v��k]��v�4�29i�R�5���0�+-��PGY{�Z]%r�Lt�Ue*4M�.�Ј/J�):[�]�M̀n�e���^�Z,�6��^V�^�I��y4�(����1J���J���ϏV��Ul<w��J��GQݼ6W[ך�^�i���v9N9�^�6�!t���N&��Ô����v!
,>��7/T���h���=�mkYI����V�L{��
�W��U�\�gКՙ�&�Qj�.\���M.�ˬ1�Xc
���Z�˾��xHeRq�᷻n����?�lv�謵N��]$�"�2��R��ŧ�  v�۪����LCUk��]�m�Ko��|��G;%��X[ǹ�Z��zm�H:/,��
 a<S�)�afc�E�m=�G"7�b(FX����S%֫{�f���kYc鶶�&3�%�t��snK����j���6���8vf�mm*������ը����I�7���ݥp�d2M���k�䘂;�ź�>3�)���޵�Ӽ��*S�(oٚ!��չ��Nd�.�mn�O�a]ݪ�GԫE6��4�YH��y��Z��f0��J΅��9`^��ܠNWu=����ĥ�y&<1�45��Q%{����h7kl����д��-����(`��.��������5��/K�-JQˠ����E���GW-K�-�ad6�xU-d8�D�6���ovnY;���/1�V[X����L(GZ60���%aV���VLr,1cԕ�%�.�,�YcAm��2�"`��*�h�i�Cr� � �K����լf�<V�:ZrV]�tJ�E�n�K�"'mǵk�&��ߞZî����f��ۄ�;�VM���_͂���Ŏ�۲]��IÉ�&M�x�y���n���l�X(mU���L��� ����e��t�TBe��.]d�cx(��1�X:�g6�A�hѴ�|��G�o�t�_����{�ТZ.�o4m&�#r��S%��h'{���z�f��,�f�.��򅼒^�+7x���+��8֠q&�*�m�T�:��#5�t���/` ��T�ңR�,@��0��[��ї3n]#ݖ7if«B���!Ͱ�Z�m��d��ˀݗ�IJa�'�G�ٽ��0���+�u�6�i�ƺ�oE���7L5ËVy
"Ŕ�+��Wh��A�����-Cf��v�䷃`����Ӽ.�1���0ǣd����I��>J�t\B#�V���h��2�/E�A2G��:( ���v��p�ɴ�~�Ɓ�ӗ��A��
v�,�nK�,)�m�hU��Y�+n�IV��;+'�0�����Q�Gw���d֠�y���n�r^�m@��!�8�G��-E%v=u{g�OwOY6U�Nu���M+{��6{E������$ivS��# ͦ�՛�	Vm�N�2���U��~�tc�ۛ:.ڂ�'U�FeI��i
�la�r�%���V���֜<����M�ƌ/r����U��Z�)��	c^��{��$Kn�Z;�6�,҆࿭O�\G@՗hWQ�z9�4�az��xŏ[���/v�`LV˭J�{{***?j�s+rLK�IaA�X@���hl���ܸ/3Y#wWP�UWK�l�pUL6����.�&Y�F@֚��	�4�!���0j:Y��%ۦsP����J��1��v^�EHF���U衰U��kP�x��[�C�rA�3�;:p�u{tB+c�E���>�ޣ�-��R��aׄ��q]�_f���c���~WY����dT�+(#a�4q�Z�xc��W�Y��^q܉J�2�0˛(9�p-O�Sn�f��cN�uB�G)��Y�f7��SU���BYYh�
��d�P���)�=z#Сq�x���ۺ��ma�)�6�(�@ո����o�L�Y�5�G��/�ݺmS4���{�&���bד.��l�P�9���|T �+lV퉳�q=Sm����/�	4Z�VW<�	�
]��wg)E��JF*N� p(�V:�ޙN��\0e_n+�N��l8�M[	��U3�t�)���Ge�+\�9K[M��9[Z�-M���ز��R���p�µ�2�V���m�s���Y+���4dko
��C�a��9]�[Kf���Vl��^<��������!����E��Ν���N���s	���h�͛ZК��.r*��|r��f���~"f33(��@�\ͭ��&
Է��w3�R��9�Y6��gZ����^�5=F�K���0b`��:⪵��������l�6��W�|��u,�D-����on����ѷT����$4��MD{j���^�@�*6m�t��vY�ї�\��0m�'U�]5g5���t]�W;��k�豻��7]��Ԅuw��o_�6�`;�(o\�4�V+�c/d(qʻ��;(#�5�3Pn�nl�K��wpY�f_N��59L]w[=;n��{���q���1�._8Om�!���S��ܭq���2���u���:��ԝ;�Ҵ9ٽL�׳Mk�s��P��+H�z�2�ݡ19d=�ܴi�v�SX�0s��+�^�y2Ƈ8� �uxd�%�Oe^X簻���c	��ż�v�A���R��l|�	.�� ��1!�����Ht�!w4��e��U��B�nhX�q��LCw+��4i�{�*㨮�7��{Q���Θ�#�<�h�����F��][��D	_a���7n�%�*
��]9وe[���X7�W��=�mJ�Z^�߻+�2ɦ�Ž�V�#�=L��:e�:3�w0�V��PՑ}���f`�Z��v>�0�Ԕo_�9�{N������Z��4���E�e��-�/=c!�ֺW[�������9	��AM	�Y�Q ���avI���c�65�T�͔ίb#O<69"E�����yҲߗM��ݎAc%�g}�R�ZtK�1��:���*u��yǤĕf��`�4��Af��,mr�8`J�k]�)έ�ܮȖL���;���H2]ƻY��>Ƌb�&��D֠�+������50��ޢ3$m� ��f�QE�_�5i�t1�.���'űT]����J0t�R�-��IC1��̼��/	f;��Tؠ� Q�Qw/��<��Qp�B�)��8��9�S&�6_uA�'�+�FS�J�������+N�걅 ��Gj5�u:o�*�^���b��.Wy	��2�L]�-��4���(��=�I��S�h}�y-��u=�p���	����f@��F� �����987���S]m����3J�����h�rH�����4������2<��rn�6�7ٯV��S_d`�c_�Ņʹ�%��Aa�$��͖y�LF�u�5S�ȆB�-��xkn�[e�-I��4�xNt9;#5 �`F�̀��� ���hip�X��5{gB	
}יɀ�[��ˆ+��VYذ�X:�҃"�ŵY�2��'|���Fi�fv�DuUȔ�0�2`]K/m�1�`�m>ܔw��(�8�G/!���}��+�`�sG�}t0t̓t�i��֝��z��̋�R�.ʤ�,"r�n�<̧l�躆�q�����䯄��#�2��C��%�Pv��ϊu̎��ٶ3Vv�4ˊb��[vB헳s|{$����	���rPPg.�� Ի�R�B-[c��&n�L���5Nl�y�51�&��y)�ȯ�c�<�_�7�t8{��Zu��ܺZ�������oa�|��bՓX��oEV���Kn+b�z�VxjB_��b4�: �%m�6l�+Ϭ�GXG��<��P9��;����j���H�<'=���8	���ٚ.��ڕ������W��f@lcV�tէ�]���i�SyӶ-�N"2��$�.��JUu�WVʻ4�=J�ԥ@��tRpev%-!{91���/r���{F�gU��K�i]A����]c��V����=8J+�o�Z��h���௢b��b�+y4��Q�s�Bj�i@xmݻֱp,���N iޒA�WJpWXG��T��'R���K�Кa��H��&�[���iޕâ4!�6ڴ��0	zfR��e�.�w��8�4E)�����t��et�:o�Ey��0���s;�;g���
�Hv�Y��wK�H��w'��Yǲ�n���A'R�O��&߅�h���X�Ekv�]�>��ls����.��}y�hS�9�+t{Mo���' �l0�Ѳަۛn�S/J�Bm��|����W�&�Z��OIz��c�nl<,ԝ�ᬍ<Y'WV�[v�k,�J�u��h5=C!c�z�=G׽$8c"�ܾ�ѵs�K鐌マ톺�1��Y�Q��Q��WJ�X���jK��P�w.��b���o6z��lŤ���SroRW$,/��}�gl[X�:�b�N���P��� ��"q�e��H]��83p�2�6H�"sDP\���^$\P'e���9i�gZ����[���6.Ņ�ZX\(�pY�Q^�V��a4p����ZF1k*�
�ki%i��I
S7���#�(]��Հ���*x�:�=&���mC���+��ˮGzɗ�r�j�ic��T��3	����ײ�F�=��s*�<�ɢ�٥o���nP\�9*4�M��8�2�K��89�{�x1�9���װ�}�c�v��L~7pn+X�]�)9�%�ۏtPR��4��S�����jk7��J�An.ך��Wd���ge
cO:�7��!�,�:E�}t2�cG6p�v���0��=�.�w����:)��89��X�DY��l�n�Nț�i��2�d�s�Q��n� �"g9�j�H�7�No[w:���������_t���ۡM�ٴM��C���h��`+Ϸn����`��I�وw+E���� N�I��Ŕ-wfu
3�7L�Q�a� ���j�5z~}�n�p�Y�Q��ڗګ�x�����]hl�d����e�k���^8�[��A�6Z\7o�	�;�z�jL6�x��9�Uٛ ��lIu��idNzj�*\�R�]�Pޑka��>���ZF�;O�Q�0�P��lG��Ɓ��k��U3��^�_$�b[�[���u[vr"�7�.�H������}a�fS���h�_M�9����8����I:���k��T�8�A�b�NOsFR]N�]E���<Ͱ��ӂ�=��Q�uUz��.�2�-��=D�;*��NT�]�+8�ڮT���jhc�"m�w^�!����VB��]����f�E%�Ʈ��)�-���GuA4P|2�݇���ǩ\��=�U��ZE�2���b���{�'+�J��h�=[0���X��G<�����!ҭS*T�!��f�a_�~��/��=�+��-�!s���x�	Y�ұ 7��!<���>��ۦ��{��&ىe��|M�-=z��*g`��V���;����&��(�����[���l��J�m��k3� ����Z��;�ټw���BV�"D1Ъ(�J������j<��b�}ĝ��[%��O8���0�n�su�V�	�fK�6a}5���X��	��-D�K����P�k��b%Ƕte<�E;o[�(`�����ޕ��i@��ۈt�5m[Y��K+��1�����s�o;�g%������E�;��l_<W�Q�Q�yƮ�5ϲ���16]�=�!F��L�����8!�
�I���V��0%��dhΚ�'h��KF�p�#p��f���2P�&e�F'+�V���o�Ҟ�	��˚� ���T5����T_�cl"Oev���,Z�^�f�l�&W7��+8^�,����e����ѷ�;_v�o��70V�0pXy���*,�SE^­Y��V�b_Q`f� y�C�*�r��ĝ�t0ۻ�έ2���o¹wd2��jw�5o��<Ȓ�����F^�e����[\]+2�>�K9;na��8����޻����	+Vx4��� �Iiu��]oAHK޾,%��Vجyx�<�(��ܯM㚫�`؋��BEȐ��}���YE�{�1d.��IW��+�������{6�7���c�;�i�)0]ʵrr�"�Su��8�ɧ�8}����Ixr����,�8zk����oJ|�æ�N�ĵ�,\9����\z�lu�#U��f2�Yrj�S'Gǥ����}����|V_M<����,���Gr�]�Bp��w隴N2S���:oSYW�K|m��5Q�-�8̚�w6�ܾn��jԑ��]��B��5����x6�9T%^a�kX|GS37ys	&�d-\}A��:�F�n�x�m\��cL�k�$E�eb�0�nd��Ì�oZ��I�6��DFIww{�s�Q�=��n�����p��*�{_���[��HX�G�k�8!Ke<M�:Ӫ��@��Y��!�{l���{B݃�C��u�wF#��n�K��k��Ep��m
ʽ����Hv��R��v<e�#.���X���Ok�����:����(�F4T1�d���X�f!o���\��A�n�����o۝�7�貎VX�e��I)Ecxو��+��ow��]p�.Q���I��EZ�
���\x�9g{��]."��z���V�*�v��1rl_b����!�u������:;�8�4[ܾ�:	��b�(�z�cb��q�XC%o��+8՝���Q����{g�jǊa*�DH�Ebޜ�������f��L�êg\���*�	y�q	D��L�Q@k�J�E�mty��rUAv�a�,]�]�M�@��\�ӣ����}Ėn�|wZX����h*?xk|uu�9���xj��|�Ȫ��C�;�
ۣ|G;�C�xe[a�9m�Tw/	r�ʭc�r����O`k]k�j�Ee�
t1Vq�۲��{=gs*�E��{V��c=6u�:���h�Ү�RqD��X���r����|k������%.�m^�l���[f��(ѭ�p�^�`(��@�r�o��J��Y��c<��aU�cU/��v҅�{2�1wq��s._}�h�ŵ��YȪ͡�-�D�a{V�����^�O)q+�'�e�ү53{%I�}�s�X�� K��t�
��Z8��N��WM=�Z�A�}Y�f>x���5/��{2�::�Z؆�Kbr}���;�Li�h���%����k��G7���E.͕�iLwG@�\N�#y��Y�e�ү2��t�mcB@6�e���	튮��������tHJ�����U�]�u$+I��ͽ��C���e���V��uX>���7$���+��9���Ղ/�%c���9���[�]�낱�r��e���	b�"y����M����8�=~E�+.��8�-�x�ǂ=[Ywy5�Ʋ��yq�ydX��7�ұ����^N�PiR�0;��]���]KTa��3v���"���6�գ���J��|�ՙ��+::s'��N��:�ʩM���l���2�J��ɫ+pn�L�GD؟N�K�tV��˴�d��&^څ�c�pʾ*��Nv[�/må��P�Wqx�[�#-nm�����2�ALs����`�����c^�Nd�T���lrYy��u��U�����܁�����5+��Ohέ[�6�Y����5
��z�����=�N�{�H��fr��V���	Q�9G�v�S�2���^�.eD�d��f�m���ĲC�v-��0��V�
���n6�9'6�i�$3�xS;�J���tS��-��c���h������u�Y�n����"=npX]�*��0+�$�ahw-���1ӧ{݊�]n���#����:��.:]f|�lfw��� ҋ�PƄD�yID4�K���X�6�[vi��;�V��܍��9"�(`�R�J�+�R�zb�7lJ�$��]����������;�<w���%�S���r�Λ�q�䩗�U�r��b�,ÙwFD2���scN�b^kqJ��i/��%u�ǘ$�{֬���E��Yv�o�۬�d\`���������ߕ#��=�h��Iڶ��C�A�����F�S;w&sd�y��d"�AʉC�+U�pܧ��t��S�y�Xk./\�ɒ;��Sս�Z-vc�
%=
F���f���Ϧ�W� �^ԝV��븃j�C)�+�r4#$e��a���1N`f9�]ݾNl���	�ܼg�p�;7�Qy�܋O�H/�繋XG�i	{%��WoG1��A"rZ�s�:�i���9�&���(jb�i�]ވ�2�ۇ"l!��YI�:\��r_G���燅�ҎE܄[ ʲ�[�u��$K�H��v��]�2�Yˤ@���
PN���V=Y�� :l���BVk���r�o��L�*jt��'����;��[��|-���<��,f�}&�8�r��#�a�:J�ƲQ�N;��*s�.�%9�r�J���y$��\0�Nm��PN|{��4$2H�B�!���e1�*R}�M���B��6Ҩ�o���rXC2��;v"͓�3��Ny
5ON�;w��I$�I$�9�I$rI$�F�m��m��m��m��m��m�䛰����r@�tu�,�2n�n	u��1c�O�:A��x���d:3���˕��"h;r������4�-����N���x6��\�hRV΄kv�2n2�w���,&9w��N&ܷf�p�>����܇]�޾{N�t�l���?��<< ���?	!I��w�����sY���O5�/�ƽ]ia���Uz���h�bu��ഷ�+ᇩ:�{9��;e��9734��]�K�
f����m$��o3��yX�&��f��w8�Yp)����tu�ɣM\�}�m-|l��8ǒ>���q=Zt]U渌[�Xj%E�V���\�>�v��7բ��/�L���*�
%a�>w�"n�Ă��O���4�:U��q��������ܮ�v������c]ǫun"X+�Z1�ktM,�����3,�ƴκU�*v�|�����jy�,	&\����D�V&��t��o<Y�K,���MY�=l�H���Ԥz!�ҝC:�S�}zMj�f�N�&��r�KF�l��
���L��w6��>�=x��� �@����X1�M�-��Zі9^��k�
M�hU���6�������<ܩ��X����RY��0�ü7�T]��.��xyFr��KjXv.Ŗ�[�\�\�9b�;w����ʳ}r�=�	b�Hݍ�ݏm6+����h��ã���$�Ɔ�����:�W�SZ�.�f�;īD�.������  ���MrMu�
���n�7T���Fi���˘�W�N� G*�,���%sl#�L�ȡY㓓�C��x�t��r�DBfͷ��F����3n�=�eMo(D�� f�v�Y�C���N���On�q��a�V��G6K�A4��އ�Pm�YR�[Klz�rYݩ�eL��M�km��oe�I��)��ل��ÜV��ZoI�%(����2`��m��*�[B��іi���vGu��S�#X^���sw6�m�7qR�iŻ;M�!���2���5r.��5X�-�[v/���Y짃�$B�7 tht~��l��V�*�K�o��8��N8�Y��55��o%,�lκ�"T���CF���]�3��8��i	����Z�[oo hn�;�,�¥l_3)�;��H��ғ��[V��-�0p3Db�:�}4��wV��N.�fj�(��ꆁ�N��tu��F�鐦��U��ٖ!����qVh��9"�
ua��������1TO�X.����L�v������wj��[ĵ'��F
�	��e�GI��0�&=MR�֢��O��`���f�n�Z�KW+�4��(�gVh��P�\X�&μ�9YA=�wo�j���kiJ�4�;�� 0��_J��ٗVIh+�4oSN�:TE��3'v�Ndk<��nmN��-p̦�Rq�?jS���lw�ع|�lC��$�)�B;�+��˳W@v��Y.��@��ʹ�^�0a�Tznr�Zi���Ay��f�	�%@ŗ]�3b��X�W��'�FX��d5�ʢG�f�K�z��$Ul���xgue��!㰄�c�������v���������Ng�R����<��._��1
�n\��u�턨����V�y��+�;����#��]w�t�|�|�jۻd��+�Q��Jw��C��LUۭ���g.��f�FVQ$ѧic�r����2�wQ'�5�Zm$��x�N�T���wG&�	y�aw7(㘹J\\��L���+�!#o@��c,�zsI��>��{�0�g�ӫwr��L^d>���dp����*|כEmBq��Y���}�19�Uq3�:��y���dU��q~��g�2�h��&�7[c,��(��n,�9ҫ�i�Y��JlL!�iB4ڡ��J׌�Y��w�LN���dQ��켅�Z"�p�x�z8�]�f��B��Ig7;-��
h.z�aŠ�ye���Ț�;؎.⺆���$Ӵ��Aj��V������-J"���]���{zШ(g�a�i�gu�����I�n��N��Ú˜�n����n�n����.�k;-�B��Mj����[FetZ�EwyM=��;����2�<�����ì]���ʵ}���o
� �^-�5�R�36�H�Ԥ//`V�]�r����&���;���̍��	g�#AW[�0�xt�Y���\	%����3$��4�n此��J*��{R�5->Ә��jkp+��ƌi]� }a޴Q���sKk:O�tv�K�=S�GM<�7@g4t�0��k+y0h��l[<���՛�F�;��!ī���)�ː�^�J��:��u$N,l�|h�M�M�{c�+pc�]I�;��;Tz�3�ue���ͥ���{V`<@uz���R�zhFw.�,��l+_֝<+^]K.���P-�;nv-J�#)JqVc�~+t�I��W�^k�������r#|�K�	�8�(k���s�.�� j�`��$�ޞ̾��'��rQtX�e�٘d�)cfe�\F2K:e��#�xg�ﯵ��[�%�H�ӤB��������bh[��� ��r������H9.fּ��q������v���J�9�u��� �馕w>�m\�ڱ�"`�N�U�zH/#&�h� �s��1�t2��d�����W�180���+8H��N'���SMswD��5	���C�����e��VtحΦ��O����g��^�Ϸ�ޗ풻���t�}e��8��.�m����8�nc���;��*JNB���W�V�uz�-�Z���t�1�A�9�.��oe{3.vZgp��C1�8VN�j<��e	�{A�v��%4}�90ɲ��n�/9� m`�Fc��=�dov�V��q<�Vej3��4aX�H��w/����}q�F�n.�vD�wk#6�I�����Ԧ���Q�Y��ec]���}���,�B��|Rf�Կ�g�V��w�˶(��s�VI��C�H���͐���]�H�#;6���ǅcN�IG-��M��+��5ݻ㸭j�N�֛�G"S��"7˖�6�q�նE��޼�D� ˮ��e���eŏMXr�o��Y^l>ts�ȹf����\��}�F�~���6��F�ՑT�d�%��D�ˁ�=х�Y4��:�/J�(E;�%^D��IPcCu�d�ߎST�Ȃ_N��f�ᒎ�R�d��ӂ�*�8lPŁ,�)��ܬ�3�)j�q�}[˔!��/h#�ː2�!�U!�KQ;d.;^���F�LX/;��R�t{d6ǖ��_�n��j5g� Y���4 �������<T���,dv*�5��T�jA}�04
3�-s�n�C}N;�7٠*Gep]Q��壻pHv;\@�7p�I����1L���6��k�w��f�@=��ɧ:�5I�ՖV*�@[!�uڐ�<vvց5d����:ry#n�e�%m�hE�9kf=����тqJٱ}�'c ��t4��_�VR�Ƌ�+P�=��̙��_+1�
9�I��Њ�[��GH�I{���*��[�(��J�)D�`�Xh`��-Jb��r,����tt�7�&�D���P��z\<M{<P����E�� ���*� ��/y��XN��зa�xM�+bWQ�1Q����Tzq���|]i�˺ɍu�����p�]�ԭ9��-Q���t쒰�1O(�ܫ�d�鵽�L��Q�9����C7y������� 9K9;΢U�1<�ν4�M�wڸ2��%��d3���j_D�3Ҙ��T��K��@-��W�!�c%c�t��V�5-�᷏����ާە�	�up�E�d����6�P��L�G7C���7�~[�-;G+��7�b!,��F�e��j��XPH���eq�@��Z6$��VfS��^�	Xf��w�^h+ (�Vl]
��r-j9�}$wǦ�z�cPW_J�E��3З�W��'�P汴#j�`��zڋ̤�x�7���Z�9'vV^j��̶p�tWK��zN7��[����,Q�un���6�����8C�U5褮�Lү<�����V1ƪX�����z�����l��	�Vs5��w�1b���f�+��� ;�K{�U��t�=�[cE���2^	a�3睶�f� �#�}˸�����;��%Vnqb�.��ZH`weY6�6.��˦�b����sn���U[�[�x�T��(���!m]�a�J�ϙ�<���Dꦞ�8�����b�j��/QÌp��fi\��|��z��N�ĻցF�nCp��rH��:�&���tb囹�{�x�ʽ�Os,󢯚�O��V�]��]yLE�}[g��=�*�%y��3]gut��%^:��3��I9���M�+�^u2![۔�Υ��v�=A�=GٝL��l`J�E�H_`n�fQV	�����|�s���osO凘�P�}&���q!7�:<��/�g���@����DO��/e8w%v`9�A,��d�1�� ����eNKp�_]�LSU��+,}}e"�H��˩Jsٯ6��'tn˥��1LמǊނ�K��r���T���/�6 =4N޹���^�p����Z�3��1q�a{��V�+���o���(m�뾅M]��NS�x]�`>Tx�I��g
�
�呐�Z�(m����irҵ	y̑ƽy�v+Ђ��c0X�u Ծ�A�M� Ĉ��N���W==�E��/&Л�S���w�
GKח��IW[���h{}�7"�Ed�9�����M����@�Jw��0f���z��9�E��<��o)��;�q�W2։1l�|�ED,Hrv��j�?�pvsh�V�S�n���n�<�u��P��=�
2ܡ����ëg�[H�}���^躺��)�{�z����3h��9�EttM���]MO�)�[�x�����R�!�G+��c^��]��x��M��v�]���lq%b�����s����S�Z��.�lm��@����]r�2Qc+#���3��3���R
�&*^i�9�eXƧ\<[��b��I[��q%�cͫ�Hu1��p�Tr	;#��*r�g�ՠ=7�]d����N��-G��8�l��01��N���U/�(H� "v8;���i뙏���n��Ћ wQ2J��yO�3Z��YhF+	�������s�p����F�-�����+�ՍlȩOEݚ��pG�X�k��I����ê[�ojͤ�p�GعmCTHJ��t�v8މ�3-�/
W4��ŵZ��Y"-�}h�!۬�e�fۋ3�`訩EǞQ�����\-���+�&��7uvح�:�R��T��=��-[���{�d;�+��.�K5Pj9�k��ĝ��;5T�0�%Bz��q�U�:�}�P�kn�����Y��d��gr��ye̊���:��&6�8����<�s�u��Pw�K�a��p����;˸m�i�>�`O\��wT����䨃��JpR��X���.��tv|��4��t5`�WJ��OA�m
e�[	d�
��v��Ƶn�i융*$�
��gfwQ�D^���N���]7&>����8�d\m��U�����B�]iwʀP��R��dru��7ݙ�[�`s*'w���s���Ս�q��c�<��/y�7 A�a�vM�cj�7��[��-d|��g�GV���(��*r^>�.�`��,�wVpWEt�(�6�Ȣ�=V��ُC{$�x�ʲy�����2�t�W,,���"-R^�!m�v3[��{N��d"�q�4L�����N'�6p�<-�,�:l���X�	���ʺ;;����5x�d��$T�����/�WJ|�G;%cNQE|�XcFg�4_�VD��fM/�zqY��m���֥����5Jխs3sR�KNU����hs6ɍ��[W|�4�5Yy�-,S��%�}����������M�z�t��9�\�L	5�C����[Ȯ}���o E���R��{�W9�9��ܸw^"�p�C��U�S3Kز޼r�h5�OZ�<�I@�PZI�X��)9<��(];����lò��M:�u��M�YB}W%O��0v]N��Zc�Ќzrݞ�N����}�
���`6+�D�M�)FZ�ys�gڊ�� \)pZ'f�9f��Λ$���>m�ŪW�Ï�ޫ7!9GX�D)��u-���H>��#�5�Ŏ��_fj(˼������L�ܬ��-l�����ڧϰ$ʜ9a�g�z�nVjdK5�oCo��Lͨ���+�b/ec��@��s�;�gm�^w>tQq͙�4�WZ6�<$[7�-O�j�a1�P�SFRZ ��e8+D��Q��z&��Z�n�ٱ��%#��р'MZp�ɹ�x����٬�y�D�#r�� �c ��܎[��߬
P��+������9u%�=��H��)o��kM�]7رwTD:ksucy�BbXJ��uHpҗ�#����vT4xݭ��e!Vp�΄�-L��	l�x���U��Z�G�i<���౪��f��{B�膦�K�>'t�:�/s��_nj��Y12S����ʆJod���(�1��-;�M�/;��S���e�s'�.b,�u�QU*��V��p���V�:{K:�T��ݶ	�z�;�W�9dv.��n�]�($և��Zk:kV�J�.���R�]����uF~��#@��31������y��
f͠6�	h�����b,Y/z�I�D^h9��s~r�X�rt���(��9��{��)�t]d��Yމ�
�)�S�yb�9�Z��6�S:�`����ΞJ���;1Ӓ��/t�o�<��C��70��:��s�4��u��`�7/��X��No7:�!Z��cQ�����o��Iu���	r�C&�Ηy��Q7˲�g� �Yy�#ih�e��S�˕y�Hr�G�������/��s��o� {��|϶�rfv̯*�Z
ΊZ��E�����N�xe*�S4rs�x�醞r�U�]��:�s��9�A0ћ�t'quh�p�iΰ3�:2��aڔ�s�d�_*N�����c����o���r}{��|박n	5��o%�8R�=�[&��C���(S��r�P�[7���C�9���WY{s�
Õө�Y-�5�P=�Pr��8��ΣڂY\��+|0������Ri��𿞎Eiݳ�������4ve:��־��ٓHݝWdSVZg]��N&�׽Z�ov�q �����[�0��t�V+SN[N˺�렰��A��	˪>'�V�%�@�s���ژ3�C�����4U7�n2��bj����%�2�0Ȥ���� 	K�f��N�j��9om��C�x�I�#'[���ƚ�������z�W<Vy'KE�< �2���E�&�7�t��� G��qG4[���G{o�[z;sl��+�]"�N�z
������[c2e�	}K"�6]����9���]��Ό�^|t�.�S�^존��o��-މj�q�f�.�ǎfݩW�s�c�uCifw]�t<S��3�{���OD���7qp��c��_!��ʕ�z9>W�Ҽk�o�(
��n���[h�}!�"ݚ��3�sɓ�R��#:ܒGy�fd�2ɐí$消��v-���m���e*��G�l�V�j+VŢ�����b�V|�1-k[l�!X5�5(�Kf�G*��[iQ�KD�h�eJ�h�j�h�X-h�Ҏ	YUPQmF�j�*F�J��Z�Uiw�LEV�j�[jҖ�ێ"�4Z\k�iZ���cj	R��c�e�5�j2����.�� �łV���l�V�ҢڴEU@�e�h5�Y�\km�*��iF�Z]Z�Ƣ�X��SnDF(��)*1DQT���F��#���b��
�
���e+(���j���V��Z�+U�Z�-�m��������E-Uh�(�Ԕm,b#Z��SZ¢�Q�*V��ѵmT�����q*���m��F�UA�ӓ���c".!Q"5%2�Es-�E*o(&%E�&�V.!ED[�cQe�k*�F�m��F�F�
ªT1%E1SlӧPUT	|h�I$MC~�]���w�V�0w\T��Ӱ�KF����tt�-A��ûC����yJ���\�8�1e������Y��.i��:^���@��g��i���J�Z4%V� 6�K�y&he��w,���X��^>w�h.|�2=Ǿ��Sډ:��,D|+2�����x�"۫�ܶ魷���	[��,w������!m�y��2�R�.̯4M�i�7YR��7n�������K��8w����e����8G������f}�,��#TlE��󂞥f �gE�)��9������D5αu��ׅ�<7�y��-S�7�I�*Sy���8S�$�0&���X1�<u_��tﶡ�l�����T7�ϋ,^m�3Gg��y�P︛�9��̂K^��D���o��m,��ԥ�,m�+թ~̪�u����L��^E��e%�zk�C`����s��d�Df��e��N;-�g�~1�,4C`B��[�l��*��^g�Z���!:��@�̯lh?�_��[}S �BU��(��c�^v�qOi�n�gȄ�ʿS,�(+5��yQ4�[����\:�a3̠���h+[N)��a�#�:R�ѕsŇ��V���yy��ݟn��d�2��C5�}V3[�u����&f��}�G���r��Wӎطu�B\�j�x�k�r�{$|N�*���߃�d�Qԥ�1��N��hK�m'DJ�hF�#(��3�5N}x�mW�ʄ��Y����
���%k��ٕR���.FzQ˞��α�����V�[�N�9�뫀���@��4��Hp]�Tϗ%@�|����d3ƾ54V�I�U��w�{��-�o��f3���A�QU�&��G��Q�p�N�s���ŝ{֤:G���Z��5��Q(�m�y�>�>ɞ�� GR��!�~��rP�˒��w����jღ�.nj�@�)�]e�\����[\\[\H�+�2%���[E}HPv���fjx�	��g,�_�JO.���fO���b�r�N�C�K!�7Q,����p]}����Ÿq�e�Z����c����^  � �NGAh��\h:�����r��:LI��Cډ?���]�!�[!)=f����c���	8V����_ۋ����n���w�Uɴ�WJ��*����0�y��K���kE��>�_����_�D���e�<���7q���{�K�{}FAg�wr�S��$A�R^3�z��ĥ`l���c|B�ͩ�U��=i��2^ݴ��ч�v�٧!��.-��,ވ��a��#R��{��$�"��˼O�0Cj$K�|��Փ��{��7�t�u�N\}��[�n�q*S�K���#����V@����֦���;]��Kt�&�t�M�c��Y\5.��В\,9���$�A����C��2��<�ϥ�^�	#�9~zVY�}�"�[c=���fD��5���$��
��Yv�ய"��kYPob�Jp�m���s��Ԗz���`�~��`!�����T�U��w��q�����L�E���`?zZӁ�^���\ʻTS����[��x��v�X�����~F`���P�8Xb�κf���ס��{/�C�
�����<ת�x��2� �yZ�)}޲����$�z|��:��
�.i1m{q�R�ofm<�\��Ps�ׁs�K.�O�Ԅg)2"�pt��T�λ�J�I��%�;�xv�;��W8���P��d�hy��>��F��+�p�hw���K�`���P_+F�ѷn�߼T���v(����<f�Cw�a�2c�,]z���~\����Hx����Ṟ����"������c3,X�E��LM��̡d9:��2y�(w�C���c���l���k�.�If��P�|���Y�(<;^�hF�Y�P�` {�~ì#,��y��4��]�����W�5�(:��O%���uϑ������[�z��m=��J�Os&]�egY��Ի��]��OG�[Jﱧ�S�ޘ�8�#��/r�u	���8��vZa2ٮ�˻Nr4ΣZ�9�6W�{ ~����b��)Ri$��Y�!�=�{Kn�*�L����K�o����aV�_c��SHmd�Qс�~)�MNIf�����H���<�.l����E�ufK���V���P�`�T��b�&�
u0��$}ډ.�4�o�Ʊ�;kHx�#��E���lU��&)�P:Q�C�<�ޞ����3%��'yC�-	X&��Ӵ�mݽ͍>G<p�����ho���l#7܆3��~�4�z��G~G���Ԏz��WzP�dך��f�d|�p2�V�!wΒ�� 6-�������<�l=R�墒��ݏx1�5���^J7��ݿPæ�bP�fR�]V괙Զ�=�}w��L�&�5�|��C��cO���-�6��N`R?u2ҹ*���|C/�X�N�Vi5��} ݜ����nE�'��ORp�{�S�����L���M�~;�"Wi��'��0�B�BΣ���w�p����I|���>#§�x\d�}�\���( �u���X^�5?&v}W��-�/�r�Fnׅc�Ҧ� ^��sojv����k G����oI�p�򎽼�/]Q���C{V���W��0�g���R�����'>��R�l�eJ+��Z��4b'�ks#;	���#����w�97��[I0`��]����)-�d`+"����4/�]{q�ۛS��� �K�J�ʞ�L��"fV�9>;�{&	�ڜeȹ�fjYo�{����M0I�$sU�����1��3vz$=7�(��4"1��vzq���Z���W�J�ё�ט@-�|CG�4kG3��2�x{]�ޫ���hE��5�p{��e>� �o5nPőE�n�VEXn�%]���]^��/Ҟfb�^s9�;k�=�OU�8s�DۘB��`���EX٦K\�9��c�O��T�۽��;�G�A�N�]˅;�/��;��a�|�B��L�8-/��߹�s1��>X�k�狫�zk��!�J��hz|e�]�ey�o�=F���Ԅv�o݊{�:y<o������ʵ������G�5뼋GJd^����5F��x�jݬu�]X���l�����hUiA��}E�8:�!�a�9���>���^g���-��c�ޝ�ϯ&䭏'�n�/���JFKݟ^;���N��P_�^�}f^I��v1{sr�Z��� E���4\TҩӾ�(��5��e�w�o�8A���.�*Ѓk����&!������k3sF�46hL�4�m�}An�S�ZM���Squ����[;ר5�$�����E����N��fgb;��3f]Mɬ�H�c��c�J(\�wI�s��7fJ�y��=��2se�<N���^�+���|~�V��{R�������.n~��9f���ԡ�qu?ƹ^����w�9����yw��P��9��w��X.�4�w��(��S�z���������a�W�=¡�����f���C�zB�����3N�������R\"��X�P���iN2�q���������3�a���3����#C��R��#3�6:��0�@u������a̖L=��=�|i=>1�x�Q��q��K�xث5��M+�����2��P(_&��	3�1{�&�~ָ��/Lr��&�S��N���#_�#�R/��Ŵ3{nq�~.Wl�}[o����H�ئ��ϫk)L�q�.�Y��!���5%��h�70w��DU��wc
��JX��C�f	�(y�<��>�/M�#�:pL�|o ���|b�)��]�u"���ƥ
�BZ>��H[�C9K=��e��D�36�3��e/��z�V����hv���%�V��Z�.+
mR�v�KU�w*����L���OI=R�t��������Xާ��LD[��I��v�����"�oF]t���>mA�7lYrSuj�v��E�i�Ի�99Y��f%o��udg�*D	-����6<G]��*��=Ee���:�����i���(��\A�����{�7����T��z�x&2�/~����c�l-E�.��0��[�x���E�"t�f��%c�u��$��2)�y��RkE��O��u�g�P0����ᖕz���hi���r�|YY��#�z��Ed����H����������)X���ؼ?R�%�ltͽ�z���Jz�C�f�M2�=jc�z��UZԪ��s`7���(W����J��}���hg,���2|�ևQ'ƴb>񹩈 ���i�����y3�uz���LY[���u���#��hp�ԯ��(���A�Y�&+ut0g���;���2صS
�c��.l��5$�27=�Ç�>��Lt���JK�	�Ԫ�m*�u���%v���3'��՞do(�fz��OǼ�y�H? UK��V��u^�~aK��{ϩk���X[PA,bt�8S��~��4�*�b��C���~����w,A��y!h=�Z��n3�Vl�)5�e�J¬$��U�F6����f�f���a����,�bLZ�z��(b'We�u�˭���##�c(bw4U��734:�u.�EW�Q�d�Μ��Nu�g�Q�Q:,X�L�b�k��g\8���p�!&�E9z�{�>�r(GK�bM�=���mƜ�o��je����V� W��[w�0}D�u�=ৎn�J�=���K�[/�mgW�-�]o{��=����9��'��5雽Rg��.��d`��m=G����X�;����J�ϗ�9C�ɼۜn<�C}�3��vMO&8�x��6���Wr�r�t�D�T[�v��"��R�{�{}�Aa��m=��(�����Cy���Tu� -{O���+B~���wHd .݈�$�72I�LHzƹ����t��޽��''�;h����p%T~?#C��y����)�}����Z�m��;G���;`=@�����l�|@���^�z^�N�T��o|�<_:�:�������R�Aq�-��Ѩj<9)���n<�e���G��S}�t�4�o�J�#I��NhMb��x�k7��Q<���uA��m	�0��BSef�!3$Qn^!\/-Kg-g>��7���X�	��V���kp�X��Γ��3jv��D'�`n����6a�F�����+|ڗ��U.9:��{��{�߻}85҄��!�@	�Md��	+���{F�d���n��y�m� ^�^tR��펹f�i'�	��;��N'qL��v�rv��U;��.�g���GL��Zo6��Յ ����$�O|�*cTW�6'�u��0�ݯD}=�j�
�����O��AV7K�bM̓�]�)�~q�Z�wQ����"�U���V��8`�v?���yysg�����O�eo+h��h�ҝV��w�^���tBŊ:��@{{��rb�ӳ0�Y!�y�r.�h�A���5Nú�V|����_v��ۛ{EN�1.Ə��n<�ňts=�"��.��Tu��:�T��G�t�=���UJ������[�.�@��r{D��x@���5�kf��� E�U�Ԗތ93�wf�=�0�#؞�ҧ
�"����{I�߰�Q�7���蠩�>8C� Ӗ��� gk���Qe�ﳻ��!��c�gmң�ƾh�!�¢�ϵ���:�jw԰����h�%iH�sJ)����]���[����6��o)�e1!�^_)�f%c9�����}z}�m�[X�"�l�.��Qe�iG��^ў��e���ŵ����71nίGM_8v�l�b���q ��	��G�Rf��K��]�G��f�t������.��<9�����%_5sNhq"��>�� {�t���}�q��=�ڨ�㓨���w�|�9Wf�ox��5�}�Q����[q{5�Hds��ڡ�H���pf}�'m�3=\.���ʁ_E�-���V'w����{�V�	q��Y�דZ��
�cv����3�������������ӧ�ȋ���F9[����e��W���Gm�}��*���IT--O���w.�g��S|xwv��T��:���>@��Վ�3���k<Ͼ�#���y���CV��u��e�X���C]b��FW�$αH�jv�j]A�+�A��z��*S.(oa������� Г�o�u�J�,ؼ9�S���:���ÒVl��ٝ���� !q����X�
��Teh����ѯCr�����Yq��Qُ�]�Z�?]�\��o*��Y�kH���1�!Y�����9lwc|JZr�v�D�4i��'���k���f�C!v���BHO���gs��U���eh0�*����9bgnc	x-kq�5�U㻤T۠8�rdj���_;�Q��r�A�Z.#�û؎.U{g�=#N�����sZ"�]o��X��'Uޣ�{�fE��i��R�Efdxc�c����8�6*�7��
-(��f:t�*�wKM��3YW��tY�+�Rk)N�����](ԋ�CD�]��g4%k�t�83[:By��5�t��[v3]�P��1���ufj�N�d]��dU�gp^u�H�7C+5�ݔp��A��^��V�KK���'��[�H�؜*Lt�}���* ��.Y��%&h���
l�>�aٍ���gwx���&��C[B���8���Lr7{�����nS�R����.������IsP'�����ԅun�,+�W}Q�p�Ki9z���۹�zC�xD!�"ڱoNn@�_4՚���[N)ku)��m���۵u��f2yR�D&<b	w��}H�-�7qTg%LXf�kOPe�qoy��.1���M��v.�ӢcHf	�N�&m=�W�����5`��!W΍E��У���uv��lov���Ѻh� �/�6v]O���C��*W|	��))8"Se&�+�g7t�%!
��h���GT��Á��:�GO�tT���,�srq�E�4�j�2��E���b�=@�;u�v��N��)��A2�L�R���e��%��:��;�3��̪��Ĵ�Rx�訽�^�Mᮈ��fM�]���5o��I(�t.����k�o��3@�l�V���{yBl���L�B1o�6�1���Z�I�z��zK'�s�W���)�8�W�la�Wvk�#X�΄Ҿ=Fm�*Y�`	�A`�
,j����-MV@��l���n��g��΋���}��Ǯ���WZ�y�WiCX����/]<b�!`SWM�
n�>�k���uܳ�A�A�E��e<�h`����e�5,ݻ��ɼzN����ԭ^j�Ur�i��r�41�\%�:��լ�� e��fٳr�-���y��0���3�'�����0��˥n.�O�,�����;�#[��J�D�(�)��]�)`3�#u��G�Kz%�-q\v����v�0B�d�|&\�ї��8D�Y�lb����v��ެ5��M@���s�s^L��b����;�Vˮ�>����};���(��,TDU��
1TX��m�V�F�)Z�lKT���hb���)�K�X��3%���.i+�e�e��,F��D�iV#Z"LpR�Vҵ+���X�--�((�SPB�k�S�R���R�,V �eb�
UnS",UUĪ#[u��Tը�m�Xi��ʱ2�E��m�2�r�k*�ʫV��Q��
�ˉ1bV�R�b ����TE��\J�����#���\�c�Qr�E!���Z�X(��AbbQ���AK�8[h4���d,�(��+9L�A#��1�.�4�[-�4����2�v�q��+-E���b�X�
�ʕ*c1�efh�����̦R�F�DX��X32��q�2!�**+B��
(6�AmE�",7��v�8ٍ\h���V6�Q�ӊ�m���)2�1b�YXV�TD$Qf0�`�h���}g�A�Zsu�-�Eĵ�����Ac�q�\n��i{ �/n��m�Tڛ#X.����夠�]�D'v>��8�sQ<yJ=�d�~Pz%+!g�z;��6�;�)�Їp��*]f��m�C��w��ܧ�0o��W�g�>�Sf��xn���	��{�K�T���|�#��^��z瞃=����9z)z��׷D���E���d�@�����ϐ!��^��>�]�#x�.{�c��/{��v����7=~+��=޾B;�_7]V�e��t��u��j(xެrİ���:����lބ޻/;*���b�}�gg��S��h�mѪ���V��>�{�nJr�1%=����xL�kwk�hK��z��L�����˧�)?@lGC�[�T{|���`^]�Du4�R��VN]rٝ�f���ۃ�=@|9Ծrޛx�ST/ݽY]�j
{>е���T��Zk��)4cPg��^����}���0y�:���*��;��m����as�k��դ�k�Y���*Gq^��w%p7�#�k���A�A�o�͊�Ǉ+ ��i!�j�aÕ�H�^��q�C�U�Y��@�\���޲;�m�[�zx��ۅ�1tǏU��&�+��Nq1$��KVh������Q�9���W��wH6�`��5ֶ�F���kk=ɏ<�1�ݿ-�A2U���h�ի��L�"�:����n6]��F��w;7��e?ac�����\�'<I�E��S��E�F�yį����K89K ��I�)�nꜾi��U뭩�����{2���EO޸	�@\�������z�������k�Y=����f3E��+zϪ�h��h�_�z=υ<sw�IV���}���q���&w���2��[_e��`��u����rٗ{�f���Jk��f^(��4A��$*=��6���'�w�9^�O�7"G/|�ۮ�FM�g_�g[Y�Y�\ֹ/T�����Kwo�O�`d��u�+D��o=��'u5��3xK��%^��{mc�W��6���h�@��-�����,t�)3G:Q;p��3']����̢8����|@���N�:ݼ���ޗ:e�SR�| ﷐�-���([�V���^=e��:�INSv�P,�`�.��<`�^���D��PAs,r�Ew�cv�{��F\��:S�$+m�Ԯ�{{�a�۰��>2��оso���XLc�dyK���Բ��΀}�_�%iG����꽯OJ離+]}7����F��������=��"��D��=@���P]�����G��خ=�t~��5����䚩����lj؀���t�ﳱ��)<��߮�����G3�L9�G�c=9��y�C&w��}~ZZݩ;��j㊢�+{����yE���E�ǭ�e�:��uė�{,�F�z׋�r���7����=~�N�%?'��
����u�D
�E�;|�u刽�{5��z�!�����-pr��ĕ��w:g��m��i��O�=6ﹼ�x�m8�lio~=m��
���ě�`���V���0i��������|�����|�zú��[L_��Ϋ���En��^9�t�"��z�:�LܛF�5�5	[�07{Yy�g!�z|�<z�
�wJ�=�*�A��u5|����GAڼeX�qn���L�LYŚ+��Von�h3{h򮠝�V��v%o��[�����Y��E8�c�Cz_a��o=ͷ*�9ȩ��7o:+���s@��)�av%�O����C��}��-o��v�O{E{�ڒb���3����o~���r�B�G��ќ�3tR|���|�)�{�_罀���g�����b ��/�n���*�vx��>�7�~f�=�Spֺc=���z��=�4�����0Y��#\��gto��l�6W�|/oc����yO ��"op��ђ�fwn�陻f�A��R�L]���VA���Yb(�ғ�W���K�3}Il�jeG��>�&��W��gl�b�����"p'�p\`��w')�1�oYn��S�7�9�9�Ճ��V��Y�����7e�j�Z���^�{�8|��v3�g���?�_|�:��}�PXO�l��u��P�<�O|��*r���Ou}I�@����5�߫��i�'��7^�'���+�	���N�a�����XI�ϩ��d�5d��Y:�����:��y���I��{�:�ĨO;x��O��|PϪ���cU�_s��ߗ�z�1�+E��1Ng2�E)�t�������c�DO�_���TG��+1w%V�ڮǅ�es�Y߳����1�x�HcVL�;r�~n���Wm�"�F��1�]2�Z�17Ob�Afۺ��s�˙0�ʱ�eԜ�m���2�QR5�Q���ڃ?/���{����f��:����2i=2�2OR�[�Ru	��ء�N �y���8�Ԭ��x�:��k'Sl��y;�d�����{��oϿF-�O/P���쯴g�����%d�GԞ�&�q����'SygO�T��� �Mo���Ad��0�N��*{��:Ûǻ֟7��5������������,���a�'R~d���q�����י'O�Ւ���y-YY:Èo,���N&�)���L�C�,%Og�`q��X/���g��t���~���|���IĜeN��H,�0�)��@�^�<d���6I�����$�	�l��'䆭YY8�&�l�u����2O�q7������}��}�g����|�1�~����X=��2w�ݲ
�\���O�4���:�&�9;�g̛;��d��\�IR~Hjϐ��Aa�����e?w���~��s�?!��I�,��&����m�c~��N>2(m$��y�>d�$�ׯ̛d�'{���'�6�r�|�~�	��5��Wï��w�MW���_����*
�~B�m�m�8�����Mo�C�N3|���$�s��O_��9������s�<a�������W�z�^��x?$��@���<:u�ޒx�2w��,��4{�%ABq�J�Ԭ�@�'|��a8��5����������7�p�$��<3�����_��z�U~�(�w�Ms��T�I�O��q�d�ŞC�'P���PY'���J���S�+'�Y4I��}�oV�7�C�u��y>���]˯��W�oB�����S��{�0��=Ϻm��|ó��'S8��ӽ�T4��6r�qY4sxi�q&��$�RN�aY>v��N$��jeS����}������.�OĔ�.��+���Oi�	o��eXD8��!�3�'�V�d��י��8I����1�j�j*Š7A�\�b��+�Sn�y%�Ͳ/;#f�Ra�h�;��{�5�ap�7/pܗ�\r�ӗ�v���hj���'������z�N\Ԭ��F=�����Lv��'��Ax�l?~�d�+�w��	��;�i8���{��q��|��O{9��I8�g�d��'Ұ#꯾�[C���w���P�A8������vN0��:{�!�'̇�����l:��X��N���gY&%a���$���'Rq!�ٴ�d�+�RI��܆���}���7ԅ'�p~⯞��_�SN�%v����	��'ɹ�2OSg�d<d�!���d�N����@�Ͳu����$��Xns�:��14s�|���hm�=J�<;������+����<�����{��z@�'C���'���.�|��V�Ěg���:��Y��	�>��m��:���d�Cl�A���z�Xo�é�I���mw���Mf��;~����N2m+!��6��'��;���I���8���'�d�'��=I�ze�d��MoY��	�>2I��>�>C��A��>��|�[��;�7���7�܄���:sX|ͤ�����'=��=�d�'���܁�	볞d���$���ÈVC�c'S��8�=J�W�P���������3�a����/?g���uCi<A@��
N2q+7y�8��s)�i����:���O̜��	��'5�I�I��3y%d��?%dĜg�d=f�8���p��\T��ϳ�����^뿙'�=gM~��$��b�Y8���)d�V}�p���>���:��́��OY9��N��}��a8���IX~d=<ֳ1��l�k���߾������p?%d�'���C�i���SN!�g�M2L}ϲd�V��a�N����� ��d紟2i���u�&�9ߜ�|�������˳����w�����Ϯ{�VI�vy����Դ�
��,4ZC�d�T�'�8��~���I1ٟd:��l����N2u�w�*A����N2i'���{�}���{���y�X�r��%t��x���<[�\o�g��-����y�巷�����v�U�G��� ui��\9g-sɩg��(J�X����:������t�3&�ʎ�*�:)M�f�eDt�up.Iy�W�O@��a,�y�۾mt�<˜�:���,_�T�2x�i������o!Y'���d�	��|�I��'�8���$�'F�`|Ͱ�g��2u�'���z�_+�� '���Җ���cV��7?T��VI���<d�I<�'S��$��l'��&���$�Ւ��79g�VN�dє�q�����q���e�q��!���9�<�|�s�V�������2N�C��d���^a�M�����M�~I��НCL�;�$�Ւ�I6�IY>Jɣ(0�'Ο=��Q����� ���{��^P}���{O�ܤ�'w����hl�̜d�=Cɝ�i:�9��4��X�
�x��!8���9���MO����'<��aRh���'�����|�}U��+�|�O�&�P���^}������C�s/6�g��Ԓ������:�9��2q!��!P�'�,�r��OY9�j�S�B$�|�.~��W�|�}�Gƾ5	���d��'���N��>�~{��N2��_̞2qO��'Y<a����I��k�d�IS]�d�
C�w��cv�O��s�]~��|׽���<J�}��z��T����/�Iݟ���ĝLa�I����p<d�!��~gY<aĞ��2��'Xy����*����;E׊���>��pJտ��P����v9��P��I�OR��}Hu����y�$�&Ϭ��?2q�	���I�d�=M�>��'O=���'Xu&y�y��;�k����~�����&�q'^��z��79�:��~g���8��|yܞ$����'��z���S��Ԙ��&�����d�T'���OfY�I�*o�Ͻ���~�}�\5��z׼��٭~���l=a;>�ɶN��xOw�|�u���	ĝa�k��'��,�N2�<�d�'����	���d���C�OZɦN#�xyCL���K��4.hĿD���k�f��ʶ��W+9'4ҷW:���i���:9;+���ıs��3,�mn�tPF�r���z��?mHA뼥�����_������Hn=�'E��/t�0A���8EL��u�ȳ:���o�_���]�������!�{�#ކT�����I��08��M��`!�N�O'��'u��k��N��d�'��O9�:�|��7d��u�y������_�k��{�����]%d�}��VM0�
�z���ze�a>B���!��8�ԩǜ�):�ԩ�l'u�2�2N0�3 }�'��w��g{���)������j������}�Z6�I�!�a�VN0��`|�I8͙q�~C�M��C�,%u7�C�8����
N�w�v�,�a���ϻ�y��u�m�j�û���t����h?O�9�ԓ�����B�O���d��䆥��+'XjZC�I�lˌ'�8��é�I���C�8���>{�Y���?����_�J��S������_������;����N2i����|���O9ܬ'�M������k$�XL��
�����8�����>a�{�}����z��9�k?o�ӌ'��ϲd�C����$�����a�O�&�ïxɦO;���'�6���&�59�%a8����*
9O���J��8��u�����s}�߷��'��N�d��~f����8�<�ﴟ0�9�'^0���OM�w=I�O�ݓ��OXm:�u�$�w��N!��o�}���F���̼�������^�7�*
�i*M���e�>d�	�O�ן�:�O�Oyd+�'P��ru$���6ì��=ɦO�z���:�d����{�_�z��<�}��ٿ�	�$��x	�&�w�T�&�IR|�ɩ��d���N0����o��d�Ns/6������7���N��|��s=�;��S/}������۝8ɶ)����|��6P�C�M�d�a��̒�a8�E��,e'Oya�N2}C��M�q��P?3��C|w���?a�Y�ӤUS��wܩ呁��H��2{�WiW�
�f���\1pmu��e�W���j������s��r���i�W��l�(���7�<�,w[)V��f'E�A^0�\5���F2K����Z��==�,�)��� ��ړ����m�Tه|����B?���2>���a�0�'X��AC������!Ԟ�h���$���d��ss�w�O��������~��y5Un��׏?g��g��C��'�9́�m��~����¡���$��y�:��a��x��?2���!ԟ�5��ԓ��n�]������OY:����0���_ޚ�=�}��ֿga�I���~�����<���'�:���SL�A}�$���ϰ�	���:�ĨO;f�|��T?r���M{��& q5�߹�~��;��}�~��ώC�d����XO��6�����?ki:����~f�8����!�N�������6w�:�d����0�'�7<�q��~����/|�}�7��yy��ֳi1��生5&�?&�,��|ɴ�Y�I�Vkz��N�7<�4��O>�|�:��?oq'P��u6�=f���~�}��矛�8�|��&�0��?$����י'̓��y%d�S�OZ�I8ʄ�1���Y��5��Ad�����'PY7�0�N��*k|�����i����o���}��	�O�t9�>�|��fd��O̞ÿa���'�^d�I?;�䕇�CE��+'Xq
�z����2��?!���� ��>ѯw�~�{���ֻ�}�}�����'�X��):�����d����s�$�X{/p�2|��ߜ�|���Y8�|��y%I�!�hz���)5-���q�������/�_�7z�A���u��_����ﭿ�u��X�y��Y;����ܐP��a��'̚I��d�I�'~l'����!Y'��sY%I�!�g���y��o��u�s��Y6�ö���~M�Y'�Mo�C��$�y�Y8��x^`x�w��2~I7�3�<d�&�[`0�iG~��B0�����ٚ~)Q&�5����qR#`{"C�J�wT��Z�3Y#8K�Fd���][��_������h��O��]uK2,��n��L=aͣ��L�O����n:�3�p���;6|�����צ.I�w� �.Kn�Jp釻
����5��sZ�>w��
�x���XJ����ΡY? �ՠ|��>f�)'�:��a�Y'��d��'{����z���d7�|��_���N��
��_V��;���}��=f�<a��ԓ��Mod�C\���2r�%d�VJ��N$���XN2~Mo�C�$���{�B�2u�?�?W�}*P����&K�87�'�0�}��'�'����i=@���N�l������~d���,��h��J���S�+'�Y5��@�'ڦ0�`xo�����߯�uV?r+�`_�&��b���d�0���u��q���<a�I��N$���!P�'�,��!�=d�7��'}�%J�y;x²|���Y��C�Y�]�S��r{����/�*�q	���<~d�{>�$�6�s���$�Xh>�a�I����N �7��*d��>�:�Ԛ9��I8����ﾕ��ƃ����l�L��='�}����,�>��vj��	��6{��'=���&�u'��d��N��ﳬ���?a�I���'Rq!����'?%a�ԇRz�6k�;��a�ֹ��~������\�a<d�d��'��&P�>�q6e�'���ϲ2q��<���Ou������N�v�z�X|s�:��14y�:��VA���+�?�|���}�[��{�{��d�+�@��M��I>d��ȻI�'s,'�ԛf̡��:��k!�a6y��l�IԞ��$�d����z�X}�{����/�W�=�v��=���q�m�|�Ԭ��;���~$�ē��^h��������d�o,'�Rm��g'�S[�C�8�y�a�8���O�}�\9�<�<Ze/͕������z���U����d�9�:ͤ���i�N{a<�8��Oϩ5��	�Ӟd����ֲi��YY�N��Y�I�T�w4��}�1oL�*��f�X��Yo�r����[��d趛 S{ӂ��1n����)H�ݭ�jS1������ʺ��*�"��}%7d�KÏCu�&��!ٝPk�m^jE\�O�t�h�� )����JU�v��VK�]��k�M������������;gSQ�m9�Խ=��kĲ���6���y�1�_̰���k��[��Q)ۥ�:�et�tm�n�nάw	/�C��%elٕR=&�"�u�LX+�EU	ç�=�i�r�jusb��.�i�oN	'R���ѡ�������J�A
Y.r�3]��h����n��؎7�ʜ�K�+���0ukb�z��(ˍI[�I�Ũ &Ұ�X߻��-PTXŲ*3��0����(	H��]������[���XQ�=J�o�ͲS��2�!z�A��k�R�G�<�i�n&������J�ĺ���+�⍦�PBftX�AX���k����`Ǧ��,�ZMd�!�Ǯ�i���.����y��Ձ�����i���p�'x�jQ�!���d���o`�v[�T���8����3�C.�������%\5Ĳ�M-ѹsAD�7Ѽǹ�lI;�.�tGZ��W0�i���õ"�����
���E�]�$*�kApe��뭉uۭ��'v����ƚ<�ɊEx�������g`En@q��4�P|k$h��7(Y���0�滆$1rR���U�����-Z-���:�����3J��_9�w`���۟bu�I�Gk;�aQ���cJ�i��>������.vD����(m�m4��YCY瓌A�JRVӣ�ཤ�X�ٯe�_h+��C�ְd
�e�w��b���Un�5�':�;	��^&��-dc{LŒ�O�u̕fM���/4��E����mhW��}Wӑ�V�������i�D@�kG��}fb���&_|�)��%���e�؄;&1.w ���0�&#d�j4��D�R���w6wJ�Ge���)��M���k\X�N�1J��X��я�p[:�����yݛ����q2��5���U�UU�wz�B�P��B�sr1� f^�;^����q���2]���1î�m9�m����psrf���C@�=t�ʺkUގN�WwC]��66��io-�wE��	+�p�"{�wؒ�yd��Ti��ho5	�����w�;4�_���-�k�*�;�z��@-�]��R9���1m�9�wukm�n�u��&�a���H�
r�0��bvelʓ:k���;^�3c�iYy��8K��w��^(�����k<87��Nػ
�dZ�v���j����q���'���v7���P�^𫹄koBu��I\�l=*m;�\�O�&]�����b��)�H���G'Y��6K��X%<�u��l]��A�.gw�As^C�4)��	��;�=5��#�矷�=���Օ����EEƣ�THQVڨ���1�
,Lk��EJ�-�b �F4�����l-��hi�����
����"��e
��E`���57����J�ֱEPT]fb�YEq�DX"�,U��a�EdQ�"��G(��
�e�d����RҳT\�³Z�X�r�:�HT҈��V֢V��0(�m%Lq�e�c�j�X��*%Eӂ\�Ur�(b��+0�Z¸�݅&!X,�֒�E���\���TE�6��d�+).����uT�m*i�
[��b"�,��]ې��AE�$D�m�l�Q�+Dc����� ��)T�Q�J�
(�������b\��eIiH����Y�iDGj��Y��Ս%MڱAe*���(((��@j�����\Je*(�%���H$ �H�@�-��l>�Kxu�G���0�j�3��v�:�WP'�&�n��6f݂��aތ�Ij��n��u̎�e�?��8��m�wk�������~��uϬ�d�V}=��N��k�l'Xx_��'ϩ?2zs����O5�I�I���䕓�|��}�����}p�o�za�;�_y߹�.vC�zɤ�'�~f滁��A��C��J��<�a�N�f��P:�����Y'Xyy�>|I�'����u�&�o$�	�:���ם�����?w�߼�=���d�<d8��i?3�)�i��R����=&�`u6�1�ϲd�V��a�N���l��~��N{I�&�<9��<d�F�y�w��w��X�.�_\�����j������}��}�V�Z|¤�ZC�d�ne1��'f�`|ͤ��>�u���/0<d�'_P��p��7����=���;Ϲ~����O4��� ��Om<���3L����z�e���7�>B��
M['�8��م�|����>f�N3��:���zw���o��߾c�~��<���y���C�	���0�'�&�9�x��&�wvN�6�o�l'��'5b�8����	�,�
�Ԭ��@��>J0�@�o�}��o�o��~ۋ�{��i.O��,���_~�|?W�}(�s����gp�'�'π^a�M��Ý�:�d��o�hN��M��q/�RS�lzU����]f��S�=��b�+������#�K�7ҥ�!�GGol4�r��WvΥ�7-�r,K*�RP�j��gg���H{ҫ���-����ĮN�K�ۛ<��Y�ɪ��*檀���};�Jҏ�'�3�sB�px���=fT���X��"}��M �;��Zu��,m��ܼ�3�<�_��d�R�^�{�ľr
.���ɼ�ݧq\�a�q�%�;�g]x�w��o��ݧ��3�a�o�g^���^Y�gXoY�m�Ǘ��T�ҋ��V���-A޳ػGntgoL�  b_s7�{ԷgST��8f�_B;�`<�@�iޖ�y��6X˚�Z�oǴ��[����Ok�e�p^h�R���1ܨ����kO�s�^�Ұ-��C\t�ɝ�k�_����H����֧��s���Q����uG��<�_;�pGd���wWe1���o����/v�l��{N�`>�@��W����!��V'��WN����y+�+�37���p��;=Y�
����;�(��9H}�IK#������v�����Pnv��ʮ��������%��
���ěޙl�C�	�`�\�=zxt�<3�X�{���֎�8X�^�y�K4��n��*~���>[[��g3����8{g��h:!}�X��9^����1�ލN��S���Ǥ�3ٚߖ8��)�ڧ`;���M3��ț�8-��w�_�~����n8d���/�#K�Y|P����GP����]ytlt�Vn�:���-�|j�C�s .7Pή�W5��%�,7�G���%:�'*�y[8�n��_�6�K�r̐�k��A��@��}�e�##����,y����[w��������gqn<1g7���h������X �)
���Cî���y�'�/b�c��;�����#}��ĈK�lN����|��)�W��M��>�Y6�+�{�W��:T�yS��p��� ��V��v=L\�іX���u{{��BzTw�M�_A�Ư�q��a|�{Ht�e�ݕ�{��`;���B��[YH�<�>]=�f~Q��'�}�~�ΕO�?-<|�+<�N�Ժ���+'.|^y}�����(.�
^^��K�����Տ�*��ɧfep����rȂ�[+�$l�n	�Ӂ�]C��
\gI�@�Keܭ9��Q���-]�{���|���!��\��-�w9Y�珃�+�[ţ��g\����F�	�j>��s��芩�E�۔��y�\$I����:���l)��� �B^ XA;���]�&��8��^=�b`��B�.*�#|.�e���ٵ.�fWI�c�y:�܌���+�B��a���Üc�gv�w��䵔f AӉ���m�]]Ԭ��1�iN	��[�3&�e6ӑhr���N4\�������y��g�=�%���~u:[Q��y�U�4v���YL���X)��d��;��ҾƅO�t�7���	s��S�d��_D�^�[L>�f��F.��������bg�{̿�7Zԛ�z~޿�̝O�U�,4��4sp؃}\=�EoY�b�V\ﲜ���;�����=���1��������i�-���W�2j��A>�.��#���ny��n�6�^�b��)3Gz3�x�g����4�@��J�ϗ�?/C��맪L��B9K��<�g[[��^�W5��xI��a���u�eεog֫�h��=;�Z�h�o�\�f9���yr���I��τg���q��,X/�*���}&b�ŭ����E�J��������M���Qͽ��z.w��]������J��,��G�ޓ�jY�/G_�,�^��Yx[�fng%5���hX��dFJrp=D^���S[�>tE�3v�V������|{����.�������c�{��ډf�Gt�=O3��6In鹑�Χi.s��`2��U���U�PRUv�np�qR1��ꯩ�A�k<���v���ug����f�d�ۃ�=Ϡ'�ק���D���j���Vͽ[�>ԋ�Yi������j�q�
�x5:�[r�.�ǫ��@�{lg6}r��eZk:���S��q��+!�sk��Zȹq�������|<�A�[�t�ٲN���ufU��ڤ&nG�:8���I}�$�u�XZ'�$�����
���rzgE{~Xp��yn�E�'�����kX����bC���:N�_^=3FZ���﮶�J{���,Z~7��W����t��&��`?[{� x�ٙ.�z3��8ά�\�s���x�@�y�u�=�<sG5�_FM+��y�2;��\w��>�#ٶ^]��9��׹1�7�����P�5hg���f맙й����L���ڠ_W�knb��X�ls�U��e��K�7W�\��pܙ�D�s�S��r��n�`+�G��L}�D�2Y�5�7��Ļ��\�9{Y�]��{-�,�>�q�F3l�ܕ�
�^o�+��!y�9׮-|����+�	��Z���]
\,�}U��|�j�9?j�@����}����1ge8�>r/,�K�����Bm��MO����7s��N��~�WZϞ뗛��Q�K�`�o7��N��;��Ѳ�J����
l�}Z���Ll?n�t�;S���)jo�t���U�k��<�+���z���J�(�'�W]���5���Y�_��VQu�*+�㳷ϯ�D{���@��\]B�s�=0p�����wq����D����3�8Vň�dʞs��垢VQH2��������B��P�q�S��q��=̕
ZrRh��e=�{�b�9u�P+��w�} y8�w��:C$�������1���vunvy�
�*=�H��,`^�w9X���St��~�[�����g��d��w��uE�[�s6�ϴ*y�k����)ds7=��yoi�z�%Z�]��[w�/�� p��a-+��.紁�gZ��qqG:�s�ƭ�v]��C�&(�OSY�Hd��ǜ���*+��/@��Ts��;�:�{P���a�YΞMT�t������8�4OY/������ﾪF�ΈT��Y��L�����ī:��Vo��='��
��ѭ
��\Kޢ�s�����0����k�g>���	����Ń�������@�z���=�>v����-�s��d�zo:���8_J;���,M��~�s�=�&U��Cމ�0�4E��qp��G����m�i�)ؗ6=�4�CE�W�q�VS��y;�|X��OAY���G�ܺ��|����PbT�#ڇ^���N�oמ��uӤm�;�s׷�-b������f�)=5�z��K����u��j���g�ߛSx�Z�٫������gc�6$[�<��7n���K�]�PێP�ھ��}F{��.,����=��될�a8�6�j���zg��W�!}�p�S���;��UP'��-���H>��9�9�Ճ���z�=J�������^ o�`��Q�N�lL�����z\�VQ�F�|��1!�1?�]��E=J��=���a{����J(�͹�	��%s�ب6������Ou�M�� ᰐ��|��'R4��*��F��][;��]e��E�Ո��������%g�������V�!��wޟ ��)y{��.3�ǹ��#7r*4i��ؗCv=C�&��'��f��Zk;Ɍ��^H���5|+��<A�x��5]��m�z궁�H��d\3��w�߰���^�+�Y��<����"���"4?w���f�w�n"��/1�޿.q���;�[�L{��ns���Q������飣�ó��Qӊ+����l*G�R^�N���ֱ%vA/����'Wr�'Ȫ�~M�����ss���^���U���>̞B��G��jM6��mƘ�O��fJ۩C���O:��q�a��ѺvO9�܊���fk~X��u���m�:�^�֮�����Ps���НP1\����^75����Nt�sٝ޸m﯊�{O���{^E哮�h;P!��`|�?Z�>w%]��f�Ґ��M�*��]��5ή^��ļf��S��(�q�<˥Z���O0���\��j�ն���M�v'�o{��嚣��i�-��JD��p�_e
��j����˶;��ج�2ikX���ۏ�b�o�����_�����W���������I�,��烑x`��n�n�������EM���b�)���'1��kjx9qٔ�B�o�㪝��l[���u�kS�J��u���~����w	��OH�|瘐��+����â|�j~o��"��L,��>����y��i�}c"�չ䯬��<����Evh�v�=���|0ud�x1:�^(.�/f�jp��#�ޤ"~�v:�Ԭ�&��+0v�k}b=�d^�[�N�@��3D.!ޞV�}�4$�Q���$~��:2w��m���A�*������y�g���Y�����w�^�;י�T�W;�7}�x$���{��;�R�=C�U �����28ԩ��f�]ս�z��o�Ϣ]����M¨Ͼ�W��>h_�����$� ��I�>Y���L���ޛ�p(�X�u󤯣̴�u&�OW����$�$XιsW�9�}�6ii�KMR��^�^��T�X�]VM�bG�,�X����y�v��O�p�2^1}$�ATBzU�5oi�A�&z������Q�̏f!�$�/��}UUK����<��l�����gZӆO.�N���^\���$̃�면�kxl�ɻ���y�}UM��n����޿�k,���@�1�s_���Լ^E!�Oz��������Q��!���b��q9���{s��{�z����O+���y͕3;�2k���rPN�h5\����h�~} �'�כ=Q���	���l��`Ŝ�r^�%���7�,q��n���z��
����]OC�>�\��}0�T��U�9�5ڢ��K��Χ^v���UQ+��g�/�dl:{��${����¶�,�mɞ6О��s�j��v<&j��>�	BQ�^�8+j�ֻ�yh=�n{��S��*��6���6ڸ�ed�G����m�K��=��+V��漀���)�q��|'��{�+?�ŋ
��֣�j�^���n���+F+-h�NL�͠i,��\m���3k�ug-����̸1a�`<Hŏ[A�nM�"��4���Kr��&��`�졜�ӽǹ�d���K�0�&������sI���9��r���Y5i�:X��g�m_:��Dp!��)�K$��R���uU�����ѻm���d����Om�(Z1f����l�0�w�y�]*�'���2�GT}�V����I`�؝]p���+x�`L
DƽH=����;�g&�������sQ�3]�ͥ�P��/�H.�PK�s�k}���)�85/@��+WoW>	Ϧ2�)�7j��z(��Vnvr����VQݳv�=�`�]"�%�@�q{�w�&�<�wG�qk��j���l��g��eZLnN(�	���}���ʁ�m�*�3Yî��f��Ȟt�%�f�B�Si���q�;�އ�Z��VR�Eo�
�[�Y'���V��5��w����0��֣	ݮGm'���3T@��d���s��6���&��-�wIT�*���Q�uK��w}0��ڻ�2�ۗ��k:�(��q�����̸"�w�W5v��`�u|���`����8�K�E��!޻ߚ���k#7����x�V��k"�4w5�{p-����Q��s��f�v˩lܨ7��ާ������xR�'^�+ww��7-���u��A;��n�jk���tpwN,��׵ '�r�1ޠ����$�a�@s����Ú�VB��(�/Y4��{�Ǆr'�
|�=�q�f�d��]k{.˥�c�u�~9I<�Y�7�zl��9�6��Z"��ZMT���
�-$��Hv�fs�uW8������D�S%̏��p�\ze����^�����r���&a[s[�b�H�e^e�-�&T3��A�e��ޤ�=��p�ܨ��G�>���Q��:�V��	gA6ݛBT�j���g9�T�O���q�{�j�Y\� �pZX��Ceq/������D����E
�ue\y/�JW��uyE�w�t�خ�}�T4Ko&��L�zU6������#�n՞�;���J����w�����+L��y��Y�$iUҝ�٣��`_+���W�#Nج�آ2i\�Z4P�h�0Wg���C��\]�#��w)r:9S�_�k�i�#��X5����sr(L
h+��E
��5����h��U8k�1�����0.U��JS4�SvV��:��z���G-��' ��}�:�9����KJt�4���{T�Z̈��B�5�X|b��k�8Et�wmY�y�;��.>��tvҾ�u4���ѻvm�va��vֳ���'i�M�w+
%Z��.+ڍ:ni��"���0v4t�,�MwK�]k~���՜Do�qE�i�Z����9���t�S��:��ef�fɱ�#d�H�oL�7�t��٘�t���HμϮ�'� ���Q�qV�L���X�&���!]*���Da6��,��J��qamSMdAUE��f3%�)�bZض�TUUA�Q�i(�2-֮d����.�JʁV�#ur1�(�"��R�c������V��*���c��֚AV���)m���T#4�CT�uLC�J"�VJ&��$��J$R���E��-1�0QQdR�*�mXUFڄĪ��LB�B�d�+Q�k
��4�40��1DGl��ZP4������m�UB�X�"ʎ�1�Q���-n�$�v�-Z�j6)Ea�ɬ8Ē��U�\����H�ZjP��g�0����X�C:N��8�s�<����q�N��ͫ�fX���\d?�}_}_U*G��%��;��Hx�Ґ������R3�����Z��Lu�j�γ�5��^a��=�6�+���c ���y8�w��:�'�g��o�T���v�˶�bp]�W���L4���]�*y8���b�>gv�w�^���\�N�r>��y��_u[�3A�V���zįz���� *��-]x�t�6	վA���U��V�h���>��v��g
�>~O>��S�?a�l�bW���q��;N�����=���k�SϦ��ݐ_�����s�=!�����]��GpDS��u�[�-U�R�=;"^�� ��@�K�{���s�_��"��h��<��7W�CH:�[�<��3zoȈä��C�{x���=MxX����f���F�W=	v�^+V)��������׶�`/c��~~���`� `�k���k��\�nw�m��ݙu��:{�t�_:��h!V���`Vھ��ᓹ�&(G��Y���X��+k��'�	0�
�L7��fY�*��VK]��i
�l���o�i�v��k0\j���C�7����z������ >�ox�zfך������/����Kj��x�G�བO���-Ho}qF�n�~�������R�RWho7��pr��Eq4q{j�j��7����}�&��3=���5�S��i�a�hvV2}Y�y�G,��̻�.g,�k��y<�q�t�O�61�9�՟���n�ݛ֝�������X,}���gcY�Ro��(3���{\uRj/�-$d������*���Wcy�oR�����lv��`��R�~<o�����u�NmK���G�AT�K���D3�����qє-9�M�i���/4Ź��l���^�UN��~þ���\�j����Owlh�g)lq;�03�~�����W�V�y�RVfn�������6���η1!�.	�s��9��=�ϵ���X�G��4bt^�/HE�<�M��g�)���,�;E�Wj�^Π.q�\ձ<r\���D�G#�q1�Z��R� �]��sR�#+��0�����t^ܫ�V���H-��r�(�����ɾv�ڂ1�)H������G��<�ޱR��O՘�V�v[�у�G���؋�'�Lf��{C^�r?4�ĩ|e��x�G\#���ȯ�G��3�'[/�L���v�����8p�~�O���6h!:������������EPqz�w��{d�>޷��[��q碗��[��5@��J�q�TB���.lu�~��w>���rz�F��vS�qȼ2OX�;U�uw �
�µ1�&����R|��ˋ����`�kjw�\b'{!��?S�J���Ul����Ĳ�{+2����3����D���U��Ӊ�$�����t\���ջ��cА�ǵ��X��l���(L�ޗ����Иs/~��@�/IO���:��j�
�o�����@C��d�g�6�����Lk��[���g�>�s�A�~��z���F���^��%A�L��W�ʲ{):�g[F���aځ�1Q4)��r�z(ߍ��X��X�
c�"X�I򷀙YR{����t�;	��9f!����Ss��޵kN��Bl㶋��s��7H��唵�/v�c���wv��S*=hf��i��U�Yy�{!��{���  x{�/���#���~91�[#���/�g�=/+�was3�B�հ�r�Gy�<��a�Z��;���2�GH��Ok[��ʌf�AlW���/i֨v�OkB��1�����)�ӷ���߾v�=Q.e�K�~��z�-�,r����V��U;��~c���$8�G>�b��yg���+zY]}����/�p�ນ:��G_ė�{wٛZ�*E��]s�~�?InsL	�܄GhGh,W�d��s[Ծ=]x��j�^�u��l�n�y��j{��ܓ���98���_�4̌=�=5�����rxzM{�Rg�r<��,��n�\��׭��u���%�U =�@�-{�O}�n<1g/��Il]"�g�9��@�f�����x=�([�����B߯��<�k�K���yR�h�<�h��;�v.�S������4e\��޷��vUƈ�{V�d�%rx�l��C]\u�J�"��o&��-�\��ʱ�{
¨��u7wW�ۋΰ�aᵳO]ք���}�1V4��M�`��'�u�Zz6�F�c`�S1"�[ju��\�������^�ߥo�JB�W��ڃ��y%�q{pƹ?��K����Y�U\��h�s���ᧄn�BͰյ�T���3W��P͍P%	d�39��`9�>с���j��Gw�pU�a8��hj��~�Y�V��%o!�����Ѩ!��'�-�8�Kzl�Y�f���;C�i�gT�zxv����A��
����~[� ��!�;����m���5�Ǡ�'t�_c������W�;����q�����] �'��#���vYs������-]�{�+���X}ݐ��l���p���btV����3�%��7�OQo`��q�ۂ� ���^����V����9Z�w྾�Qf�{]ۚz�l�gGS��nN9��Mc����^�
�(��FZt����4*}��K���^A+�I�	�\���<v���%�T�eq� /A֯Җ?)����:-y�o<��'Q��"�X�L!�l4�6��x�i�θ��f_Qͩ��4��(Ծ�Goc�tnv����u�!p���';F�����;A���W�N����;�bO'&�4f�4�Ωٛ�t5&�1�1ai�}_}��W���nb����~"+���׎{~��)�z*��돽ֶ��;��H��z�	�+y�9��'�ɸ*g�[��-�����-��y.��Wz������4B��d��t��{��5�Rc2��jWW��U������s>6�l�yc�(;�/�<ON���{<g�V\w�e�����'����<��w��'�!,����~�q�݁@O=k4���;{��k�+rp�o����,zJ�	���Oì�y��E��n�Ω�ƌ�}ݽ���3��!��&p=��M��ǘ6�꩒_l>Y[��:g��'�tC�`��@�T}���/V{�<맧`���$	�;F���Y��g}������)4{<���Ϡ�e1~㾁�ƚ��rMTo;Ճ�lj�۵;�d>�;��J:��%S����j�T:�9�cزN[�B�W��)fLw����C�g|��⒩D�
.�ӶR��qWim���7�2�]��(�}Y�YW/�:��]E���U?���
�GOYZ���񻭜㙹�++N͕��
ȯ���f�r��>�)��9���}��W�7ܞ~�-�1��!E�}����Z:��u[G�S�ЮI��ִЕ���,,w��N �-�_�$�jר��;j�;s���/_�TZOϚ�䶧{����$����t�c�h�8��vu����+�{.ϼ�\�:&b{kN\W[��V�hu�q�\���9�:���b×����[v�tv�|�la�`�d�����6|1ܛ�`T��~+���q��5Ob�8y���u��Gh,Q����^�tyeۘ�j��7'�c���j���L/�m�5�K�]��ۺN�.�������ҧz�M��=l5��~��1g���Y=��#�E/T�ma�7R���63ٺ4o+�_�<�Թp{|c�]H����[�E�&�D����ү4�T=��)�o�{V'YP�Z[�<�9!���r����x7��:^��p���z%#Sʼظ(��Uْ�������q��vAv�����̾ϱ"$�esf��*�C���cX��E�.75�fv�Է0�ue!��1'�ͤ�m&�f:��d���:M��Xu��v^�*F?}�W�}�Ȥ��;��������-�����j��蛨��*�t��q0�0���`��n��$�z+�gj�o���~�`=@����ԃz"������d5۱�z�0�jWT�+�Oo���`�}s����xyR�B�=�/:~� �%z����7�u/���χfޭz.?�H�KT�M�+5=�E���tX�9l�Q�;�o$��!_�|<<��KNBM��>�R�-�y�Wg.���C8[gt���;�C����Z ��u���-�<��J�ܫ����V���.TA�S*������p5���#���i����:���[Gm�}�1apr�1%,�fn6-(r��|xO�TO�dZ����2Cc ��?��:�Y�]�bJ�v}��G3�f�}�%H���'ޯ;o��^ӣ����|vO|�1�wP7+&'�v��tI���J� ��jf;�i���r�o��QX�J�Ј�iSF,3�!0����I��<�S��9ol�����C�|%'/qӥ��B��3�dl��YX�m���Sj<lV�MX!i��s��Bm�������Ӷ��)�˚�������_2���"k���'2��s3d4=7�_�������:�Bu1\�!�0`����&U�������׿��d�#W�#ŀN�h=�ftO065��&_�7�udO���Q��q}����@b��qn|�^
����ިy��w���՜��b�o�$�E���SX��[�/�k�����s똥<�{��̝(U�byܗ�����,ܥ`����#��t[���%Я����I��Y�RΛ�x�/��QP.�˿�u批=F��|�g�u�A�EL[c��m�܈R�e吣�6R{���M{w�"�oK���0�,8)�W�T:h�����<8o$L���,�"�=[[��f�i��/"�>Dl�<L�B����,r��@{<�V��.��n	+7V����N˼����Y���^I�틙�lX)�N��3����''�X�nSϼ�no�^N�2Ǫ嵆V&����.V���i�&k����؝L�$�n�MCװ�f��l1��N�ݡz.>p�����[�T7�;��e��#��-���RL��w�7%��o.�{|jZ�q�/=���yg�,�-�+ӫ+��֠}G���/v8�z�Sw����B���=�d�d�B��0յ���f��5
]Lo5�mJ�Xs������U�\]{��7�5ݚ��b����Vp��)�PӪ��x\�+4�8MJ��>��9 ���<�����׾���P�{��[}S/�H7V��>D e�'���3U(�-�$��^zTz�rcՉM�r���:��S��e��Ӫ�����e�5ԏ��L�h���h��^��͹Y����h��ؚ^�F)��ɇ֦�|�sB��C���:|�k�g]t��&ϊ#�Nݞo��bKG��(��ɺ8)�3<w�H�d�/�Y]�1�B]m0Wo(�`:���,�{��h�Q����wfeO	���[�mi�����U_.ğq��	c�3\�,)!B.$�o�@�\�K�WS.�
f_S�;��(y�%�7����L������0��0<�|o%O/�C�@��i/�w�Z\7/_��f웲��l�26��B��LR�"���b-3��~&�HC��qH�S�;1��ˣ�Q:�Ͻ�9���D.�$˙�4.����Q&+�n�2\�!1*��=����_$r��*�4?)����t��U�`�R���qt�T�]�fnЏ�]�Vn�B7O�b��Vm�@�8��Q�݁���4�u�&�)�.�2]�
��TI������a���y�,BY[�g^�J�	:�NT�I��y�{G���M�n��W�'ѝ�Ƈ
W�����6��ƈK]*�r���G3=��B�9J;
�]bC�ץ0�++����NΆ�ͫOD�棇N�]�`���j�⦰4֜���$����g��*���e�v y>��!���'jWv�u׮��¾˒���.Q{�8Vu�n�:)鵂P8F���&���4�NSZ�]Q��c���|E��U5�SW��X�,�M�I�Ԯ]�K��bŪAnv�k]3�ć&K��x{�����[x�son��e7��Ӯ���ٍң�DV,�k6MdC��
c�`O���CrR�Ň�	���E��]l�%Y��{(�[AX�&gu��}���k�\e�5G1���dH��N�Z�3\���{�.X''k�����9��d�IU������YlX��Et*S;�h��Dmܲ�L
���3^ڽ�7�j�h{��!�/H*ĪuB�f�υ��܇A7C[ܘ�6��qXr�;٭ޙ�!j��c��ƣ���+��ʜ��n�-��#�7�Ԫ!�W����nq������42�Vj�m����R8���nL��6���5)����u����OY��ʩ�+'�[S�S�^�Xkq���[�0Z�n�V�*��jj}%q�#'�!	�7�D�r��}��C�h�iL��Y�`]bQ��*Şg��r=�b?4��$���D�;X|� ���La�ݎ��S���ݦ�*'D�s/ih<�E��}؜os^��Qp^��0�S�v��%�����:�G�/p�W;[1�D;�'�Sa�ُ�����Y7�]Zv�;W�R��JKB�ZFnS;�Z����5�Gln���X��\R�,��E-���+�:���J�����I���y��6�T�����ҁ�i�O��fz�Kڻ�UB�3ZN�	�D9j���2�XJ,S9Yj��Ut�NRj����	�j�$^ ]=��b��Utu	�;<3q9��!���Ί:��۾٪�Q��$&�x�|�s��b*5���E�u���;���/�.���v�͕44ɮt��˪ѕ�L�g+�g^�}B�.V2��y0�� ����`�ffk�#q,m6h�wl������)���� �.�_����_�ן0qӪ)��7V�Y�*SI�X`򩙹4^��W��-P��O�>�l���U��>0g2ͳl�>C�N�F,�}f��x����S��S�e��%�;F�/nū�lD���X`೩�Cz.� ��&GR��]�8˛touiH�l�Ed����H8��u=I�P��˥��:`켓��[Mź�ޝ�.t�XLjl��{\�I&���ԝӶ�3������Q�|j�S*(�����	����m��U��-pE-��\Lp�b�X�Ь+(�bcb�TAX1Or��2Q�B�J��(�E�L����(�UJ�Z���LB��UH�e�QQE5l��f��B�@�W)��Ԡ��V�1F�eTY�1̹��j�.Z�$��**�%P�TQ���%���sx�W�(�E���:q���m���1V,r�UQ�C,��QEAƙh�(��c�6ԥ���qF�mxY�U�m[k
Tm�F:��\��E�n	��9��iK(��
Q��)F(�km
	�b$B��T��V)�\��D�YS,lY(��������EKX��*�cF�3)*� �D�mዶ]F���˳�*f7����rv`,�˗w;�ŻK��X�P#�Nm�1Z[��\��SẤ\��,�V�+'�}\�u��v�}�������}_Q�������9��mnu��޾]����>�r������>.���[����:�?d�ߛ��;����D�t!±,�o�0X쯊}�ud���t}���M�W��p,�y!�ז%>�ܷ�L�yKB���yu֝��{=j�e��Y�����MC��Ũ��*	�_��~�H���ݥg�f��+��a�y��I��P��j����S�e+�">�eʝ�׾���	W��D���[�ف}��'ס1���O��a�s,T�̶y�v��ӝY���@l�梱�l�~���9B�d�(kZ�me�\�z�S����2�}YUW��UiԮAC@�(@m�]P���WqO�<��bA�������:{os��
#ge%���tv=� ���I�:&B��b�2u30������mЄ׺�VJ��s�_�unլЖ%�[P�W]=�N��H�l�iI舺�E��]��H�:����А�=�v���U��X���9��R�Φ���^�����9sv��yR]{l��a�=��.�v7ƵF���ْ+�r��7}^���x);�;y7�-<����N�9o�z��j5��poV�Ih7M�,���H�<Ů.�	CtjT�ۜsD#��reN��gF<����������/���}��&Ȓ)�x��ˢ�����9�|\���ΗH�T�����\� �G�{���q�hk���+���,��!J_��Ҟ�%'���}�/��讀&��IE��r�s�ٛ�틠M�n)�����W� �1f��"��˘|4K�Ծ�B�W��F�)�f��h��GI_]�ePtV�R��j����(9��Q!��]#�e��1�YDLY����Sv�ϫ#z'�h���Ȏ���GP�u��P�g��S2�\�D�3��W[�x��>�Y�������ă�i����ǧ�m���^VnS:_/CV	}��ƥ߅<׋����tg�`h� e}޷�	����O�ٳ���f����y�����wwx�n��?\���Q�m�3�Ι�zG��lg����/�ۮL�v�[�!���\�t���>�%Ps�V���`W�vD`�ca���\�K5J�#+kk	u�͎<e`F��us�r;GN��.�x�15+X���k�B�A��$6�;g��~�p$㷙I�:�U�ˑ(p�r��9�ɩ6�-�,~>�k�� ���+]���Ulb�Eڋr�"�:s�;���Uwu/in��c�rʶ&'��:��,̘�t2��R��f��e�**�`�B�A9�^JIf=�A뽎�Wi�����8iR1������y8��aͩ��R��=M,4ҋ
��}|*Dlc�0���N�
�*��<VY��4�7��D����|�:ȣ>/�X)qh�=*�X=z����������X�\�Ç_�ا�+i�"7��auش�*r	k��Ft��k��j<�U�OB�aOM�������s���O��`�^�&x�����`��j��H��G�&j
@��Y����]+��t�|�C���b�[�O�2��9أb]wef��K�ש5WU-+C��o7�z\����F�O�i�z�4ߦ.����ɩ�99b2m��!ȅ{�4)˧Sg��kͳz;L�.�42R�f5�PR��qA�״̶�FLW������^�u��9��5WAɼ���!V׬��,E��I�ݚd�w)�JW-��Ѯ�e��_B�����0t�4�����]U���օ���D�`GW�r��E�.�k��%Xa]
�GT��s��p��}x{�s~Ex'.į4O����!X�dC��6& ����\:��}c�|���
���r�pn�t��;��ɧ[X�{��ߝ�
�O%|n�;���"���p����M�o;e��b���w���[�P�J�,�G�������
�5J�n+������`u����Y�Z�;J_yN��z\,��ꪪ*�ڞ>[�)��L�~�t�b�?@Q�,|৩X�|�}ư�Ny���HЌ>�&��Ҡ���|Q�e9�؆.�2m,ƥmhs�P�L�އL�ـ�|��}^7�re�����zg���%�*��Yf�|�Gڞ+�����c&�q���N�P���GQ��3�k�av�V�+��?]��+�~�'�p>"\z=�/c��r;\�F{�)c~���{�](�d���;[
O�P��}A"�i���_|o�U�]Iג<1��y��}�^Sd��z��eM�c��r.�շ�3��jRn�C�>D#,q[�K�v?ws������t�;Ó'7�����uS�<�xf��N5�l|����W�x�i�et�=z\%��z�{���*���)P���<�I�tb��,�}jjqb����yM?��o��8Q�a�7�V��옘���p�T�$��=lQt�͕`�mM[%#���>6{��W��Vҁ�9]{�.i��c�o�	����a
=N�]D3�eM���0��v�>����YH໇C�Zg��b/ByL��ң�Xg��pR�֋O�X�f	�����귇�阪"��X]��`��&v��v��E����}[L�h��#�l���푮e/��*�x�;i�PM��LK�թۗ��딝h��
Ҽa�ڕ��/�W��}K&'V�s���,���l���j�wdS�&﫩�t)���:R��B5��N���~ݭ��kؼ���-���lU�{E���r��\ER�C�Ě�y]���y׶UO�q�|��:�/_Z���ȃ�A�R����Za����%��EG�n��W�<��>��en�}o�)<8�	z�-�������x.��^B��1X���J�|%����T5M��R��a�^v���g|~`�40�qpC,���8�[�(��|V����4�ދTT[���x��cЂ�~C�ؤw@��Ϋ��=�$KR�7S�}���'�y��b�t�2
~g�9ᗁ�����B��x�0q|W���)�8zQ�w�*�u�R����s�[����*��&������Y;�L�8\�g,k5{�ɍ�X��xʤs����$��]�u`T��Fe>s���xHn���SإL �Uz�\xk �������oU�yw��)�\D�m��5h:�w��u�-g�	Ag�\(ut0�]R|S��S��ȥj��h�2�%H7�u�i���z,2���˕டa�+���/8S�6�(���(�\_n���ݵb
���9􃭋�nE��V3u*�/��ov�ُ��0�Z#�7��h�p�PJy��5:���gpM���'^�.�'�{$%fa�־�jG���,FF?}U_UQ+ښk��7.+?�uq��T%g@�0D�1�C�+��c�f����s);�~�15�TP�;����Ra�ꍣǥRXI-�} ^��I��D�U��b�2u3-+��^8�����ߥx��9�>�?2-����W��t�*�S�}O�W�ڐ�Ͻ5	���n���Η�c6����g�׋�>W,��*#M�&	:�Aq~��n��<�ˠ�����k�-��Mv[���z���
����6�D���f�"+�`'��+�v�//`�^m�A���7Ҧ��m�fP�5��4��'�L����z0<�@E���k6�u^f�oK����'�9��(M^���3P<�����KXC��r��+�Jb�^�跳6߲q���H���4�*�K�2�M�~橜Ϻã
l����� �H��ц�}�W)}����Φ;�'Z$�y�b��I�|�r��X�n��S�%��➱�6�7�������b�7f���t<H<��.����<��d�^qp|�z�M��,B����� r���z.����M�k���� Ȭ"�|E�c�{��eȯ_q�G�ɬ�P�o�{�N�����8m���Eyz�ȉ��=ݬݘ�ƪ��Z\X�֨�t��kӥ��{��Yj˗�4�,\�3�*]��q�I9�.r�������דSۆA3#�;�ΎY4Y��g�&�C��.�%�yb��U�o��oU��9"��A�"ezG���[jP����4q��xi�W�VC=���u��(����n�7��U���UB�*�Cq�؇�;Pf߆�b)���4�]C��0�cY�'��g�=&�y;}l&M��6Y9�O��x�1E+>����v�A���`��d1f�Y�W��6y%˷�L��.�0Xf������Qh�ZU��>�E�~&}�Jf1�کK���=�w�4��hg҄:�y��~Q{�4�i���Ѫ�紻čzV��޹�v{69��ܮLy����E7:��]v-8��3�8^#� }V%*e�fǟ����:�T<����wz�ϩq�{8S3s�L��Q�'y���6��t�JDh�<�q�j�Y�V�s~����	��R�0Y枞�:��zd$,��!=�W-�FF��O޽���u#lw�2���0s���8�g��VmM-����tY�BG����(go?a�ρ�=�Nz�}�����=%�]�g�'�[E7�p����/å>���;���h�u��^����G�3GUu��wY̜V�kJΥ�)ڹJx��
��������8��鎟Y<N��{r/��0KJfɵ���E\GG�~���}_UU4���*y�R�����$V��P�u�P��(<״���e�����Y�n3������w���KL���X�EL��$�n�2U����r�@�z��#q+�u���k�O�[Gx��N��I״ʫ:) ˡa�a��$X����}Qb]���k^i�K�ns�te�{~)/r+�H�qSD솞�D7���x�}��-�~[�;βK�����w�x��5sz�B�n��Z:S"�zX���|:���.�gڼ1��rI>K[`/x��v즰^��e`��z���[�]hl�5'�P��[HO&q3�\�v��M|�W+f�Ͻu�d^��Ar|W��ʳR�Oem���/b�=�P�n�`���bq9�W�ZQ�;���ݘ׌Äׇ�iZ�`��ӆi�&kU�Hke{�wS#T�sTi�ֵ���T7�m��c��o��
ӄ�H��
����(R��nzX�s;<�{ō��N����}N53*h�c��E�:���^#R�uj��G�u͠��OM��V��`�ǒ��zW=c������K8q�L��԰j�)Ҫ8��9)^9T��QCR�J�Τ;[8mպIf��=�����^q�ΚN���a�Vl�)i�>�`a��84r��Cp�j0�u�5������|�n��]����pKY2��꤬��7/������W
�"d��.T9�:�ߴ�q�gj��X��t|6(��]�J5$�om��7kOi�*���J�#�V���4Ҷ�S&�&SS���	�ձ���Hi�^��Y��*<j����3�����T�����D��(p��zDk'5�FA���.{��}"է<����tP�T��H��+���&e���R�� 
_��tc�SV3͎�x_,3[w����,��u&I���6�a+��t�X�Qg'fzo�^l�׼��>^�Q�^qj7FfI���$�:rd��y*yx�C��Bl�%�G�����[���f�ˮ��.�!�K,�:D�̔���}[�>���`x:[\�3��ƙ���7.��§Էz��0�gg\�D�b�������6$4΋���{��4/�Tp"K"x�u��7�o�>c7s��lL��/�[�O��P�s�`�����gY�*�Х�_a�.v���̆*�_1�HN�Qի![�b2�5�	�礻5�O�L�
�y&f��� Kޅ��;<�z�X�4s��]z>}y!��FU�2�;AS�XvAx͜����\����3���Wn���9�,���"���횭�A�\Ȭ��t~b�&=R�����i/�石�O[�Aن��s�r0��/� �Sۼ�&#�a��܃��3�z����M�=4��P���t�mC*�6�$�4�xlOs���6�M�dmz ����� ���{��s����,'�"��7�J��m�ƫ.廭_��h������`���������W�\h����[���hp�^��=�.��|(\�y������K]x��p����`ѬÀ{1�Ɣ����S��.Pֵ:����E!{�ݑz��.�z�K�V钾΁1b
�jx�)��+@w��~�xie���f����Go����G�JK�*�Z=)���J�Z�J9��J
�FR��Q�����'ug`.�Og��4;¨D�Ljt���t�4�H�������{�w�������>r���W���F�؜i�f�xDi��&�ZԺ��S>x�po���g�-�Eo[�]��d�:�휞�[��y��-���f�"+�\�{�q�:���1��>*X�ܱK���ř�k��NG��-x��EuR���<K���NL1�9�*�%kBme���f���
�o�� ��[ĝ��n�:.;{yR�Jйfbp�b�Z%����)�jwjKr�k�!�x�{v�ј	8�#��,Yn��<D�5���=\Ü�UY���������֢WK���U�����"��j�&�3��qۦq�d�u"F�ᳰ�ͼ�k#���2�n�o ֆԭ��L�%���=ݖq�dhZ��@�vl����ý��fwp�$�N@Ȏ'�m%�jXq�bq�V��w�����d��6�00ẛ7Ye#�/uw35ᗢ�*Bb��KQ��wkM���W>��[F��:gw$� ���g*r"��R������w&����f܈�w�1Lbw�����Fdၾ>PѫoR��̹��
��Fi9�=�j;]6<}mn�uj�3+=�����!=��%.W_\ϣQ�/]�j�;� ��t���U�/5�k&���t'&�����!��Х�[�b{�s�vo���7�`�\���&=���s$�X�*U��@s6s�t�x�=m\k}Lt!��j�Tu�^���%"m>]�\���	��YR�呰J����L�
����u�_^��ؠ9�>�G��*� �n��Hu0eMkP82[MZBѱV�-�n��ut�4˳oD�n��7�r+{m���B��Cz^��ǚ�M�K`�laʜ*惵�2nE�d�Z%��j#�	�ޱM���&��o�Y�k�*:21Hnj�hѵ1�2۴�J1�����vh[�1�*-�RhYSU�c��d�!�D�Eȴ;�浳��}�M딝!��$�����a՘�:`#T0d:�_O��wF��2iTȍQ�������$�zƫ5�r�ouf�5r�i����j��6~r`V���]�<{p,t���eܲ����\}�p���u���!�7Jw8N�l�r�͂�%m��vT+
[(7���nu�S��8��S�F]��A��z���>9�,(V��>�RLkx���kEk��D��t�l>��ס���}/UI�r�*�Y�t,��-���(sT*��9�:����6]��;2�n#$Hɣ�卋�Q����@��X~���k�����]ş;R�WԌ&��0��$�Ѳbe��0y���]��%v���M�u�đ��'��^oP8��"���!�MH�Hj��Y��WiL��8z�6�
+�[���"��Z���SΘmߵM=�ʙ��^�<����;��lknp]�^{j���V�bhٞ��-��+"�c�M�y�"�q��D��x:V�� +Sy!�.cVv�{%�5����$���I`ݵ�x�|�߳S�L���(sS!���Wn�!���]��M�o����}Yt�b�	�͹�BZ6_I}6V��'3k�I&n�b�#
Gķ�S���-��F��1-[�6�W�QV��iP�*#T�[d�m��R�T�bV�+�Z2�����1`��J���M4�2�#DU�QPc�F�kドX,���¡��+R�%dKE
8�DAL�*]d�\�*�dۼ��*�f8�s.fLm�6�"���"�j�i�e�2��8��ZT���
�++���0��ej�k%EU�XV�H��Q�k*i�b����!��Q�U��JF�ȭi�b咢�F٦����J¥J�F�e\�m�Z
]���YYPFJ��6�l��Z�)U+���E��6�V��\B���U1�f�ݢ��
�%���%���Z�ʃh�����J�FЩm-�I�6��aPm���+��������\;�@�
!P�Q� �J�J�AKiP[F�!�kN=�����t��uDj�a��s+��ݧ�[��pd��.�/��1�lwǮU�Z\2������a9���#��W��}��~[��x��숀��4��Y�WS��1t��b�!�KN �K[��OZ�����|��μ8`��ʉ���,��ܡ�P�腺T���3��S�0<�ܳ+g����}�獴6��GF�<W��N��I�,�Ӕ��Rk6��P�bf>1���z5^<���v����P7v��)���Ҟ$e�.�T����`����ע���n��-=�b���_�$�o�4Y��9�d�0挺���Kʬ��c�+	{�ٖ��j�k�+G����=u��0�zG��l�O	��U�U�wz�a%{�����y��˲��iP]�t�j�}�%y�{�9��pO�����^�zv�W�5d�)�y���u�8=v�;)+�'�p�e˕�a(+�t �䃇����l����SY(3pq�+r�L�''O�ݱ�F
�UP�k�%a��8\�ٴ��%λ�ݺ����z鹭Q𳳜���Ț�����K��,hx�0�P�W�u���� �1PvYY��k�YX�WT��S�6U�D�u�����*-Wgz%�9�M�u�c#5�����Rt|�Z�t����I��p����fp����$O
����]]5���t�J��DU��	�8�r�KX���˨*S�5~���m�{��rcoR?����+<H���L.����˨e��.@�B#�5�y��USM���n���Cr���Ey(1��o���dC��I��[g>�f�D�u's�=6f����$����n����d�K�hz�^��g�zx��Sw�L���к�ݷ��'6[|�b�ݠ�ۗ<�6o-0g�Y)r>)�|�Yު6��.�����G#�G�x��(z��j��������}�4W`�M+>ل��3�P^�aӭ���2@�j�+O�z\�������RӀs��*�E0Xh<D�n�2K2��JW!�����[�R��d��7�_����#��.)\�)訓�h2�Ίt�hhXk�Dt{�n��C�UВ�g���y��^S���� i���ȯ).̯4M�=F�B��g�J�P�V]�������egn�+�&�U?l�?X���tE��OR��u���$�z�k<s�۩@��!�x��Jk�἖��t͇ݷ�FH��>�_k�ɚ�?`ׇx�u�3�^�ѯ���hVԬ�z�P9��_�Z�M�C�w�F�"P�,�/d~a��'L.VmY{=+A%�=��d^)�xΗ8W���6mޝC1�Gl00�֕qXJ��,��̨_#��|SmE��y'8���o���Avf��Ǖ��c�(ASD��(��,���/$���j�u�z@snNtZ�},�N���!86^��f�W}��p珉|~�VY�*�u�O�3CB45���;��k�c�{�٦���D���tF�c��o��
��T&�B���i�"��I���r�G��;�]nR����8Nbu0�eM�c��r.�շ�2�dx>������ �:ϣ��y�BYX҅ʂ����N�eB�Q��+]�7�gU�{��>�z��t6A�8.l�os+�F�P�K�M�C��l�L��:1M͖L>��)\�ܐ�bK��>�\��W�ϐ~�}z��0ң�!�wn�.J�@_&��X�������j��i-��̴/Dr[��v�+*3�� �/��@4���Y��z�9���/�s̩��Ho�1���ꮅS�{bݙ��v!ܰ�n;��="�XGR��$:�@��D���h&eŦ��3�=�3}��o,��������gKr���2]����C��P���8���뱂{R̫/E7z��A�#٫�s�V�����t7J�� :��7|�o����yP�\�\ՙw�Hk{횺��9>j����m�i\�ܵe$���b80X-k�T��ҧM����xG�3+��B�Vt��ˊ��sf�y��F\���Iȼ=]�p���W-jYp�ޖYt�7�fJ{���P�Q��C��_�����N���{I�r5���9Eg���%�t���C!�T�<I��Cډ1X��ek�<m�Oh�S3�H`�	>�e�YeKt��S�ܺ��J�P�~��oH���V�����`n�Z�𱞍�N�l�V�*at8An]��̙��:�#+$"pr�Q�W���ڵ�G��Ș9���½%�>'~�<W��yKL�*���u�f���t�ҋ]I<_�;�ť�׹:���K'���
T�{��r�cC�b�}��VmZ��-��;�������Yĩ�t����A���0�Uz��<5�"�yY�ʢ����Y����ڦ^�O+�����x�\C�e�(/��LP��a~�fX~���9B�_�'�U��kt�=vx=	����_5m��@�?�c��{��Y� �1b
@c���
��d�%��KuQ�(�u�}�ϡl�v7\+
�6��D�>2�%�ҩ�|1�UK]�IG�d�w�v�e��]D�һjR�nƾ�$�z�Q̂r�3,��e��1j�{6��b�:;tB(u�c�ܚ-�z���jr��Xu�0e�i��A|v��Tk���۾*�jv�I �D6c�7mx�GA����-��b�ܨ"��/�U}KӛSqf�i���^\ӌ�|�>hw�J�,��/����|�Z��D	��O=��fZ�i�/.�����>^/J�PK4;�Qk��$���kQ���Lө���~=��;�>�6Ƹ���5J������Z&�ͬ�-����$hT��+B�]Z}�۳���1.Ŷ(P�t9&v�����c^ ���A��}^b�9��#�}����xL�:��Ϭ��&X#_" B�v�5a����u=�\gH�liEKr�[5�guBi�f��+cy�}N�C讀FD�IB:��b�^�~-_ ʈb��=���i���_�pڡgyV9��y���$�IH�V+�WK�1��1������j��-q�ow�L�k�lR#�ܦ�$�t��S\���:��	û�g�/O �|�������s��C�eQ@���/�sS��eynZj:}Oy���E�}��+7xQv3g�ٍޡ��m�1C�y��4q��x�O	�j�O��{/�x�<���5���1ԘgA�}j�Ko��Ϲ�=&ۆmJ&JzM����l�|����1�(F�8't���ʊ����J��ɒX��n�-v�{�gX��7�L���59n�]]iګE_q�3F�x38��TT�~���R^ٰž��J�*��[�O���KNxԾ�+��}]��xϼ|�	}�Ľ�v\�|�g��fb�؝�X������,�|��ȗ%���5����n��1158}Kۖ{^Ojbi�|,���d����{�|D9j�])+���Z�ͥ��{��X��5���o��UF���M���	bW��4=��¨z����E�o�5����{�h��_cS�}���xS�^O+��u����Z_99u���/��Ĭ��v��h��v�m�#t��ʬ.}
K�����|��9ւH��2���r�e(_��۽Jy�z"��,z�����\ ��=�)E���Ƀ�������{zR��nڈ1Т�-wnL�2q��9��Y�|h�҈��+��h�V[y<_���^gl�#g.�E�/�ݗ�I��>7�uۡ� hr-�C�"�7f��u�P��Ǫ
���z�K�Oo��x��Ji����8��[]������*�,�`��&۳L�-ܦ��u�&�Nŝ��!�����t�0���Q�z����4��fe��OV�j��Gr��}�Z�;����3i����OL\�sN�x��NMܕ�/-��c�8�SZ��.��,�EX�r��<u����ne��Z�&/��\�{�G�K��e����w�p���h9�Y�G����r�)OED�{L����̺B�C�E���L���R��ו�vۣ�w��|�Eﳫ9s曺ݔ��P�W�&Ǽaׅ�HW}�9˹oi$k��������i8�l��'���>���2.�ޖ)c���<Kw»�."��IL��:�{:�՛�ʆ���Wo��Q�b���}��c(R���`�/l�ݾ�>�=���I�9>�|0<��%*a�IAr|W�`g��n�;<�@Va�ZS�۾�\�YX�t'��!��/e�=��z��z�8My���k���
<+�4mfe{?u4�S�x����{�̕TEϣ�e�.�����Q�>%C�}ACՍ^�x2P��g���lS>��t�6���!9��'S��#��E�:�Tˌ� �\�+��q�Ow3�����d/�����LP��5	�b�C�j�w�z�M�QXk���U,<�����x����*p^#[U�eB]�śA_�@���K����0��\Ӽ�.���/��а^>GhX��}O����U��K�W�,�n�w��4�~�-�~�K��]`^�:a�X�X���fD�{QΡR��vȇP\O]�<�����U1�9v[���,[�+.#����ɷ��;�ݑ�Ht��/9�R��.r�_}�/.����߭��2�����1P�o�Z�x��:?2�\=�(����e�<��ql�{I��dΊ�ܿS���U�W9H:EV<�iV��?���Ŋ��]?Udb,E�x>��SCt��x�N��}X�YK����e�Px>iV�	W���Tj�;ڢ���|��Pw�Yx���t\�i蹙�e�Vt��%��*yx��\���{����9帝&Y~<�%+���qg�)4=�I��.�xey�0�X�	P�3�(-~ٗ{�]����||I
�.)�{}�,����o�Q��yأ�j��*ޟ#㴲sn��6�HZb���V��	]a���a#�FVypcNx�=�]�$��;�WW
+���y�r20����@P�fS�/���UP��˺��=@�,|R�7:�j^U�E[��-�o,�����7���U��`�5xm�v���򡚂2�m�Z
m�}E�d�y���v��W;�޸�}�4�>�N޿BH���iX8���	��{��]Y�'�J�:;��Z�3�-ˬ!��X-�<ql�׷��sE�X탈uB�vR5�[Ygr�M�Xyk��t(�D��ou
�a4坚���Ӫ��W�;z��+f�������\=Ѫ׷�.r�딅NӃ	����(��+��������_G1]�¿�u!�k�㴘7�`�u�L.*8tc���(n�`��w����=7����Ƿu0]�9�\C�e�(/��LVWW3{1�oޖ��ܡz�/G�l�D�/M��f[� ��;x,�	���3藃%��b���C\����u�Nü$Һ����bع��T�I��Y>=�`|e$�z|���? :w�7�}]#��k��rtKeA΋^.u30��|#>�Mߪ��IbL|}r�Y��9pH�ew0�WzǣR7��߽����D���1p�D��ݾ>ϝՙ�=\%�QI�#�t'�槎1<��=�=Y���-�?B���~�(g�3�>���U3���%�T�&WU���P�X�O]�y�W���1��X��bK�n�w=��~1����%Z���?)^��Y��H*q�˱v�-���" B�v�4����+����\b����KXC����*��s��8�m���x|7�r���r�ʳW%�Jr�YT�T���gꉍ>܉r׌�`˻xQ=��V�3]�2t�ڤ�xN�����[�z5�[�Vq��eh��޷Z����N��Ջ�����o�}P$;+�D$7���ط�m��P��s�ݲl��-�-��$[9#����Mǥ�_���6a���|�W^<�M�*��uO �ԮU�_F�N�I^�#��^Z):X�y]�y�\�+��;��5Œ���{�3���]J�n%£&�
�f�� �3�rXu�8��g��Ŝ�L=�OW��]����ehr���v��3|�.��W�1�|�y�o�;�T Ž�yۘ�GZ�ۧ���N��b��Ҳ
��P�.�!f��žY����4wv���'�p�j�'��O'��	�,Ub]E�I�/��J��J��+��.�����ZU��_e����7�9��K���w[ѻ��`U�����z|�Ä��>�����]�zb�Rk�N�=���-m'���
F�̋�����1�Cx*�l��+���r>�8{d�|�s�ڹ�6q�i�N�X �]NE�-��į3i��Va�C�K��m�^����wՅj���<�`3�h��7�1R%c'�I�&5]�M���2����3��`L������k�~�S��!fØ���Yt�CX�S��QdC��g�rzw���7���r�����M��]]G7
�ZZ�53y��6D��-e��F�ZsSV]��e�E�7���h��gc��|`�&�ŷbgb��7�pW]�:7/]��!�3��yDՒ��ى��G3YJ�V^�)�����gLF�l��Ѣ;{0J�K).������q��Z\ra���oq>�ff�]���#:�0%8H�h���l��+����Y�J�Q&��z��SkYޓ��o�ѹ-� ���`=�����i�т��kf��7�e�S��a��`̇3��Z�3�[(�F��J���+�d����whǻ���ԁ��]����ek|gubM���v[�";y���� Cpd�l��{��+�\��e�	5j���lw��_wv��G\X]���o���; ;:G��z�gl��vڿTL�xh��w�i��oq�\!����CMP�����(��ri �Ź֍���F7�����r�L��E�c�ky�ئ𩳫
�b��R<� 6aKn�,��|�iȍ�=h���T�5�n��ܷ%=8�㔵�Z��x�$
�ʙJ���t�U��M�Ե�An�����ٝ��5SfbY�|Ykb�ޖ�(�^)}���b�dR8Qɂ�,��gyĥuU������o
C�Gx��k@Z��
���9P�����@١��<�zί�w]�]p�	Ӝ5�����	O����T$��4�Q���e�SrM�{^�,�[�o:��VİKsK�1q��ʾ������w8��K7���um�-��u�Dd�X.�b�YS��n�yu.��YJ�(M|���6̽Y�Sp�p9�8v�눲��N�惗عJt6G�Y��s6�[Ӑb>;����C�NTA�}���!L��+�o �j�-^�h��:/$���$�hr����u�2�Ҡ$#o��<5��:u�V�(�LÔ�eb�໥�s��&�iD2�;GtV�cDZ0Ѹ��;����,�ء��t��d�ވ���&2��R4���v��1�x����eb�1��-�S�y��֡�� Z�d���ʛы��Vs���sa�#ӳ7��IY��k�V��b�� +YY��]�ٗ[R8һ���Pdem�
������D�l[�����0�q;�eC�=���c��	9�D���Ug�㼻6����4�[�;��ʙ�I�,5������6;WG��i�`5��.�]�]��wL��䨻�v�������}�f��-1���H��祈�x����IWN���3g:�op����M>`-��Qv:�w��5���L̦��U�B���A[$N��dn�W��\k0�Iv�%��S�,�.�C�g9�eTw&�>yH��f�[n�r� �%�1�JGe�<�yeWL̛0��l�pd;Z��M�Ӱ��LK�ՈU��D��3֗��۵�'i��j�Q�S��X��d����:	�6Pئ9&s�H�nB�#!����r]"C ��#�l��h��W����J��),cƋ1嶥(��ŰZ%J�VO[�R�-�5P���˪Tm�1iR8�aR�!EBT���QKi�.o!uMe%`����҉�Z�QEl[EP[��a
��&61%�a��6�fm��2e+Q��F[J�h��M��T3)���r("[M��ʵ"ʹJ�[-���`&�V�R���j��Xc�f�*"i�raF�9���D�Z�Q�Sl�+j�h�VM[1�c��j�1�$մkk]j�Z˪���-iU�D̵�H���J�q�f\r�(��+KE��[�+eZ9�pV"\���&%�aZ�3Nۦ��.f*e��v�*�Lqr���Ue�³��&b��(�
�[m���B��1%�L�R��.R����k{��l(Ҵą�ZT�
��Us0����1%D�,�f,̮k1�V4�7YX�C\F���m�%j]8∢���2�*"�mŦ\r��* ��63:j�7��M��Т
���+;ڳ��M��4��S�O��f�ǍƮ �1,f���,wG�<�V���QW4�wD	e�����DѥH��U����e���/��*�	� Mf��=��9N��z$=7�(�ˤ!���}7J��j׷���RO�RU�X��4�R� ���Wg˺{+��m��|5��ǂ�t��S�"y�����CD9��n��"�7f�ۨ�(h^�5���[���_|֝��ꞆE�/�X2��"O�����$�M2z��k��b���S��������%Ր�ѮÂ�=�r�TI�o�UY�I�B��v"H�6�o���VF���l��u��8���K�Z�x�M�j���4L�"�D��4�B;딄
.�r�SÜO�~"�i�*�q�YB��>�޼�~�L�ޞ�c�
0��zT�YR��l�==�_{3QP�Z������|��W���%���=,QO����a��}���f�.������������3��V�&? ���P\��Ȭb������<�h��/YS/��s�����e����7�s9�����81�^=�	�3��Mr�f+��/|Hw�cB�ձ�J���
�Q<�y�R�	���+��zf���vugN�nu�:�fg(���K�.>̷��W��r%Q�%����I'1�b
��d�pE�����c&��V��o4v�ivDY���v�\w.i�_Z����of�c��F�o�����W�`nF��3d���������0����
��o9��@�Y��m)b��
���	S*�����Lm��?K�0C�Ov��]�Q�b�#���Y�d��痦���;H`	������%�c85Q��2��3J�y����o�{������J��ؽ]���Q���mh�#+`�^�e���:1M��ɄI����clU/1X2H�S�z�&Г��h���8���������E����{�å��׼�ST���s�{��{�DtVWq�*á�*��DU��L/��`��~���1�I�=}�N.�hM#x��i��X�ͥ�T�p���+�6h*���"ߦ��#5��6<c.������K3'���t�m=�IbP����&�~^e�B����l�A��vxM����+�B�ʼ%fq�u��,�X���]"�JSb��|<<���k�b�lyf���4X��.��U@�,�e�ş%�t���Hd5
���]/���?eT�ɵjH�K�u���!���ޝ}R�Q�/GI�+�=�.��״=�3���Yh�D��TR�$D�Yj��m[ �Z�L�R��~�C
�����K];x��Y.g^�R�cSX�ꬋ`m0����ʜ��[f�\�2_o8 �
����9WNr���T|�<bx,��_�R�Z�7ֺ�;��>�"<��
�xDsǆY�`��{�o�/p�}�j��8V�xځ���'��zK����X~�O���C��ND�jۖ,�$K��u����\ד8^��ȺϽ�q8�Z�b)}%�>'~�<P�yJxN�lo�#h�؟��}�I��S��5��j�o<�ϙ|=�i�+�G�v��뻯�o}1,\�n4�єk&�܎�̞�����2�Cg��0s�P��~�����c$��mZ:���]R��7��5�t�]��g2�+-	A�b�WW3��w�+%���zw%H>�S�,o�š��{��V[���P/�n�D���]�d�3�Ab���0�y�*�2w�nT��S��=~k����x�#݉W
�I��Ѵ|x��U$�z=� �ݱ��Ly^ujI�}϶�ryd������F/'S0E�t�C�@|��
�u���Ub�\��8?��-��W��|�������Bk=5	��j��Ra،�gӂ�3�*�P��X�]o$����z�w�*u�lmf&�[��a��bl[ƃψ�+����=����X��wS%B��,;�B�̉��T�]�:�ǭ�����|�X��@�Y+ ���`W8���L�[y�4�jS���m9�U�qV	���������~��L/�=ܴ�`��g������qOj�7}&u`9=*��7�mf�-�r��ez�qK|���J7����\�_�(t��:-�NO~��5��O#�G��w1��:R��U�^+�u3�~&	f����I�GS���Vz����1�~��V��G*E4�N�ׯ���WXZy����+�L)L�5Ie�����:[��3)��e�f��(�����p鷍eK�PI���YqV���T�|�U�n\87�4���h�%5]$~S�W����\�T�Wt�OeJ�b�%�)q�Z�Gj:]_k��|G�(��B����K�t���q�{~�+�\�W�f4O��2M��(u��[�|ϑ�#��U��ڎ�Wo�{�2���c��^ox\Y�[j���4|1�hĞG���'����=
�4f^��։u�����o���Y���^Y���=G��W����Hi�w��,�:�[3=���[khڵg2Y's���.K���U�7�}�I�8U�����n����O��5ߖ����0�0�9�4�����qC~۰�:ӥ��QW�uݺu��o7���~/Z���>%W��X\���6�\[�dÁǷ���92^��v�9X�
i�mlZ��f��t&l�Q���e���e���.S��jc�oh0����jfi�=Y%Cژ���dCV�z�Xj-�ZP���!�Yřc	y6�G'��	����8�����O�S2������X�!֥9β|�>/�X)q�Wf��9({^�mi��(���
��	�}�\���DWI�&��i�Ƨ+�v��\懲v���D�*�R����,����r���-/cݞ&1s�Z�rw�.ͬ�O�M.������7/�O�-�QupR���49��0Y螞�:��.$<��W���
��:��{˶)���D`�a �����Z9|}��ϭ��/17Ex�]�ܔ�gd�{�ޛ���e��7�{�6�Y�S�n��,����Iu��(nR���Y�/Q잏�������n�/똶��2��D*�b(L%�i���
W�K��P���{�:v1j�RQ'\���Z5�Cg����J�:� ʫ:)]`�h�{�
L�t����qbYđ>��8˩��C��+�wO/��+�).̯4M�=F��lΙ��˴��һ�:���^���N���]f�;�#׋���s*ZB��\�$\�ز���v��^V���c�3��ZI�qGN������$�v��7E���]��&MU�Y�	�ڸ R�١6
N˚�G��mI��H���%=���C�c�ۥ}�{S�VÈW����H��7z�-)�w�,R������|&#��ǹ��sطe�[U��y��,!��H���+��Mp�2���	~����=2��%w:�7�{��DϺ0�������^9�W�g���N��GR��~�6��;�G�}K7���\^gz�MO����{ �-��[[�b�����HN_fz��+[������$���z���[��>���quHkGbu2$�n�tF�x�8q���!<D̛��o�aM,ĎE������mu8N��m*r���09x��~9�-n͘���T��4��F���"2�����k�P�`ʅ��iN2��;;��������1��\�����n������3�h+`�\�in:1Mg�=���{��՗-��m��'�lQ�R��N4;�����G���1%���zآ{6{�������}Ӫ6��
�����sȯ�sȎ�Y]���EV<�DW��c~+���|6k�b��8�+�[��m�i+�bf�-�&�xk�$�wt���[:��n���9��%h�G[�:�A*�ЛW�7^�*Lb��NWn����C7�ط;qTBN���C�
�h�rV�Vza�6��v�����Xr��Db�k6�%t+���p�!��R��>Rx���,~�~ɵ���{N�l���U~��;�E	f�5A�H�FwmN��oz���j%��N-߫��q��t����kY�:��)��e�Vt��.��J�W���^��~��h"�СC'�g�ۮ��\:=,�H�����j��1_���-kD�~A��p�dz�hǱ��� ��r:G�����{�=�`��p��+�x{;ǆ�_�h1�\gDP����"<>�b<"/<�;01���0(Kӷ1���[w�Ӝ݄���]�m�-ju��Ca�,R���ś8���K�o$��0	􅰃��R�,SX6��uWAA�a��K]N�@3j�m��k���3�x�/���QY�p��{b��ͯ5���P�<K'3������9�Ц)��/!}�vw5����C=Z���#0�^u�ğCG�b��R�����W�5ǆ�f�*3��O!�Z��L�`��\{nX��T˾����}�b�W3{1���R3�f��~ټ��8��X���8�c)�@3ی3۵�^4��w�������:�E�}�6�܀=�^;K��#ޞ�J��y���>pq�)�����3 �V�hc_ua,Z��RX��B�#�v�b�6�1�8���h7z��6`%�_��G����J�\�W��T���)C����k/*�/��j�>�=w)��t/��T�����ۗ��f��y*�iӲ�K��Q�uÍy���W��u±��a�f����|���k��.�wͭ����� {:�p�(��'S0E�s�3����hY�l�����Bh�H�wٳ�,������ymHMg��<tK����g΄j�➮�hr�=�������ݸ�6�Fu+��Aqz/��Q���MX�B3>�/�N�k��3��d!�֣�I�z��h�s�n\�ݕu��1U\�m��8�K፩��\�=!�1L�9��ژh����<~�&Ŝ�%3����},�2$I���Pz��^��i<��U&�v�_Y�7q����׆���d^GD�+�L)}2���e�����B�bٹ�]����k��{Y>�L���ف訐��.���z}�ĝ<$���=4�2�"�Z�Bp��k�}V�!���O��)�R�9��d�hh��iA�U��O�H�<���.�r)J��g׉���	x�Qg۰�Y�P����ms�J8n����w3�*�n�x��m�T��w�'غ���A��M`��]WOd]��1X cn�S5�q�ZJ�MC|�Q�e^%�2�/4���kV%#��U�sO�7�s���u��:�P�_���<�`Oݷ���&cD�9�d��}}�3�ȟ�n�o��c�F�!H�Wn��o����7�.,u�����<�@h���D���gE�A���rMq�+���ν�z��P���WU3�z!�]�pm��C��ů|���o���'�Ǣ���3����~�Ị�`Xl��Y��%���^%QJya��t����54���T;�`�AÀ53��]!rzբ�|4��s�X�^�+2*���n?p�z\��k���{ s){��ΥU!��LE�o��~=�,Jtm�Ҭ�:���>,-��Xِ���+�3է�}w���U���&��!9/�7��i�h�����js�ӗ(����i/!�C��m.Eu����K��C76Y3�\�ֆ^�<꫚���}xZ���gVg^.�).��T�A@hpW2Ef�O=%#�|7=z�o	���nm���=P��yĉͼX�����=�����~4LiDp!��COڪ|k��4�G{IN�G������b�{!��~�wg�-���gET�[�����{�$Y��O��]7Ξ�7��e<�^�ηN�w@�*�9�ɘ�4��).T�P���Ը&���ּ�B�8lERo7#�L��Jۥ4��
��O�T�.r��.ժ�~��1�/�N��3HNG���6�Y�C�A�3��-�I�Ց-�Ve���Q�e�|��G5_!~|Pu��3��_�1^W����b!W}F Cߞ#A�G���R�x$���sݎ��D'Թ`֗��y�gY�3���p�J{Q']�ʺ�|�!�UX�K�ӷ���g_�>;��f_�B�3\}u[��Y�3�7E�Xݢg��B�^h����~x�R�K��~.^n������"���*b�L��y����^E�)�v��K���(��s�;1��Q���y��-P_i�G-��b�[�}���Z�ͩ�Os��/�f�ŷ�����5):
��� �<0�~d��>T��'�����!`S��}�4�=˟.�~m)�v�PVz_�!�=�&K�e�=S׽��>$4��vwޛ\�)wE9�V�1",[\�z��J��{�]lu��y�2�~���Ov�{ZQ8�{N�=������z���(=���/4��Y��1Z��g��b�OS��:��̬��#���;Z����U�u�.�\&�'�S����i8)ܙ���h�k�qB�"�X3K�'^��85u�V�
�u�j��Y��)���\܈�8g^� � ̎A�Id�1�팋�y�%�e
m��geF���:����!JW-��*I�����	Mґ�l���Y����`4E3z�vk(.38��Ċ�{P��h�F�B\չL�Ow�#�*�(la��EKB=չ�z���1��qξ\VE@�V&���Lp�d,}
_WV�[���̺�*�<�c�Ǜm�y�NnC��R�sd�F����fJw���[��eq����v�iXpŧ���7]^99��Np����J+���隍�JI����N�{d�����-wj�l�yX7lM��@�h.ޘ,��%��"Z�C��#�L�Rc���>[��VZ�G0�/H�V�.Ռeӡ/.��J[��+0M��NP#�20|�_#�U2��R����W��@u�Nu����P���%�Y���b��\(f�i��ʆT��N���0*QF~���YW��cTRô�cC��wd��e��b��>�sN�ܪ�f�D1Y�^qX������132�=ڄhHr�V��͊x���5U�:��8�5X����X�-��_X�\�v0�੪=6��z�D�ǘ��4ƴ�.��I��eI��SEv�Y�f���f�;�`�/'��n(N���YIT]��sU�U�=� ����3@�eT�N�A��F-���r?Q�QZ�K9���@�	`ٗ�?y�S����^m�����4VMh�#,�՘�����S�";cwn�)9�a�mf��N�E�(a�s���H���F7uxsI<�Ѵ;:�H��\�N�Ά5V౩�v��E���v�B�e�^^�n�ͩx�d��t�Y�B�a�6��Lg�h�#O�|�ה7sn�
;��u"_7n$�ԩ;����Ɲ�}}���U���2��}�"d��oWp�"'m��ޓ��t �Ty������M.��mm�kY���Ub̂e��5��hR[�	=����y��;-V���*'n����ܲ��]{�;��KN�%�-�O��V�$W<{���=w��q�j�2���vx���Ĳn(ٯDcG/��lr�ц�������#f��!/�rj���LG�VPZ-�喛���#U�7C�i5qk<]']K�mÏed@��{"��x�g,�O7������MU��q�Y`��;Azw�I�����R�]IкX�5��n��4��7ԀE��׻�d<e<H�UX.S[fE��21
�27z/�a������J�Gj�Z����\�N�K��CK*�A<�=b�u���X:��95����ِ<���c��u�`��#xM#�(�:�_Q��9��z���6d��;rC�-�$�̽��"(99EѰ~��~j)���Lk�ֆ��p�0eոY�3�#�u�®k&*
Tm�iS���"bSz���Kw��c��v�Q2Ÿ�(V��p�*$�%�Q�3+��,��ʍnTLk�fD�EQ��X�Z�˘�l�LG,�+YR�L�9��hi)��+0�).�ZV�J�Y+m�neq��N�cTimƸ4H�T�nfq�Ӊ�a�1.P��e���q�.ZZ�M[&Z���V��(�t�cE�PVТګi�.Z%��Qՙ��*��Q�
T�c�M��L���mSmb�"��k�D�SZ.R�X���r��e��)X�*"Ya`��%�3.j㢖Dj��U��P��,]$��сV"*���Si(�ULTFUUK�mmK1�)un��c3+��t�qƭ�ն��+��-id��[Lʪ�L��L�����9f7-F�,E]ە�Emj�-E�\�1V�
�KZ�C�,��xVG)R�h�3"�i���U�̹s1Qrժ�QQ)i��UK2��``ъ�c)0�1��PE4��L�n�t��Hf5ժ��U���GEl�[�4���D-һpv��W+�˓2m�j�U+��iSI���뺝��ev[�VP�d�ݖ��("5�YQ�=ک��w`ױZ�Ij�e��C��s9ĺ�'��zq���������{���^]������Ԥ��Mm��c��p�ap�Vb�C��:�4Z��yu��mgp1�R�Ŧ:~��U����l�Q��=*�C�X+���Ŏ��Vt8W��ct5��֏��E�>��Y�SS� R��s���]�/�hg���2�U���"<�,�]��k�n����� <m����P�Բ%w��A�QU�&���Y�5_'�G��).ssg�G3�GF���+�����SN�gԆ8�iL�I��+H��YW�=��)K~���Qu+%�.
����)6�ҋ�e9yX)�y^�fgVd
�����m̂NY��#g�@�p�KԺ.I������},�:K�H{_?y�r�r�k�lOK��W��3�>�m�;=D��!}�g�P��ŉz�-�R�2��4�Q�ۘ�����Q�wU�uL��:"�'��,������Kbg��S�/w�����.,���ܝfwL��n%�]3��z�ĥ`{gL�:�x엟�����K��ZDɤQa�شK��:��b��_%y����~�u��X�=�*�9B�,y!%1ڷYj��LPݽ��(&�gp��@��Ǔ�+����u��[b���mN��4�.��U���J��re�\scۛF��NfC��Ǌ{�m]����g��LڜG��{��O�B�!���q�>FU��ۨ_5r������ ���X�<�гS�W�{���4�>�N5	#d�v�\��E�/b���x3��K.��[�������=5��ۚ�=W���=��Y���K�Q����kw�}J���Ƽ]��|�Y�׃"�Up;���K�����f�(;��dX�o�;��l��<�Ѝ���٨|;Mx���ڨM��mA/:�����=�lO%u��<e��Wo�v�����B��ayw�L��kޗ��g��:sc���kNOoY7�v�!V2Q��N�f)����`���
�uOv��W$������&,)��羐+��H�BZ������r���kJ����a�����5ZhtTE�bLKb�qz/��Q���MX�B3�b��4�?'�7j�_��[�r�ؘutD'T�t� ��(P��~Y��bn��֏l��܈z�6��S��G�x���n��H�t{0�1�@y�o���t��P�-��q]��sɭ�2�/;7��k��}��Ȳ��HP�E��l�ܰ��7H��*����#���9'_G�V#��.��k4S�}*����|����d�qѺ�JHM?Jz��g��L>�@DI(��ʶ��/f��q=P5���F���6�h7�4����������]Q+Gށ����Z_a<+�Ѻ�lz٨�e왋���n��늝aԧA��Q�A�X��Ep���OR�ޱ��ܝ�t"��j�I�,t�3|z�u�'tD�̩N]�^Y���3J'ֵ'���bs��'���{.[���W{��3l3�yY�Cj�oJ���r�^LƉ���}���^�w��~H�w~��+<�u�������\��~5/5��y�ʕ�=v����]��.l$����]{���D�t=��_��*/����o��}v!ߴ��G���]/����2��9�2�K�q2p��wxX��a�i}">=�).I�k��yW�G%��ڝ�AY��3�$8���!t�H�w�ݱ�9AՌ:U��}�Ԡx�{��H�l��.���K�N:�qq���s�WD!⫨Z�`{7*@	y�f��<Tm���k+�����|��'"���O�d+2������)�;��WE�=^�F�.�/����R��<r�����m92ݕ��mo!P����6�.����x���Di���"Z��W*Wi�l�Rs	4;-C1Q��EH��E�߲*Xl��(_gQ�����k��I�b�J�{�'X��Ŧ�6�������9�Ž9�w�O��O��-@�A�#iw�*,{n|�Z^�*�6Y3��ó��\�q�o�wln9�8��նre��"F��
�������>��-�~A9q"t8TԼEr����4緥!=��]WFFU� �i
"U��v	<rR�� ����=�}�;�_<�3���:ϸ�!|�y��۔1Kg�<�M)�a%��>;���"��׼����݌e�X��~6�C��a�m:���[N�^.a
�C���q�n����ʙ�e��Q�v�8������o x��f�}M��>���To��%Ү�S�����Op�S]�����$�r���,KЭ��!ֆ軫ݢa�B���.׈��i^nf�y�=����֤+C��*�UԽg"�^_f��~��|:[��ryAS/����6���|�!f}ݝF���A�}�ʭ^"��m�C�k�ᗖ�n���H$�.����@ʍ�x+MծF�߷�哤�%�n����`���M�&�Q��S���Ve��M����v�'�n�R��&����Σ�Y�{4SM##�޳�-��8ʤɱCq��xorn%����
����ءC����Ϋ]Q�̓;zI�K��E�_�O��}s��|Z[��|��<�N>�C{ӄ�������%*ad�<������k�%��oF��P��g��7��+H�� ��s�'���8&V��UCv��r��������[2F��r�g*,]���V�b�T��b�����'�W�0gZ�4e�]����e�v,�0	��%锎
n��*�~(�u��įo����]�܃�Vه2l87r:;�2 ��x���x�5)0ng<����i�F{��61P�{|�76��n��U��s�j�Fߧs�;��skڬgE�v�dhg��IkE}L�=��IK�=K����j���u�h�Y��MJ慉Ƈt������M�ȴٹ�����(���ng��Ǖ�e�G+�!�;����gJ�9�RS��*�͑+F,���秛�0�^�x{��4��a��x���ϩc�6����#������=��9��q�z�d��	�h=n�b�D3��'�P�]���3h7-V�Dg�/�����N���c�y�>����mr(�c�e��l[�z�S���bYD�-̓�I�'[���(�(���j!��:,����Ŋ>�*Q
ƃ��LW)0�&��VsM��X�m�7b`����t$���~���|���Ǿ��{��H�F��P ��V)t\�=��җC���!}� ߍ�v�eB=���Q�{^z8j�Xx�X���Q"��!}�KJ����
�W,���?RВȍ9�g6R�1�ڣ˦��G�U��3bCL迢������	C�e|��#��:��e��~ޞo79Zu�^*��}J递��B��f1Y�L���!1)O	�'N��*{����~��ꬑ���x�\�su���=fT�ET�@��c�HW'�4��rk��b��^���g`^��+)c7/��5He{��CZ:Ǫ �eR�����MhY��(��7�B��o������ w��7f*��D��ш�m�R��ؽShC�V�ު6������=��7s��\<����^��JK��^ue���e7� {lS�/�{	��=7�&��2ڽ��4�V�)��ȥj�2�yW+�F���#	�T���дxQ�n��J�44N�b
�4�=r������z}�c#����C�O�0���
�������*��.�&s`s�������g�&��'��,���%�e<�����=�?#*U�Gx=��������2�Q�;M�	'(��Z�;Џ=ux��)נ��F ŃRI�6�5#���.>���,�:�ِ�NA�_}���%�O{����I+;�zK'��BO��&B�d����"�q��V�!՜�c�+n���LN� q0{�6�z|��Ҟ�@���"F�P��d�k����|�F��8Ӣ��]��7�e�0z��^tP� a,u�«�����)ʘ�L�#3�_�eG[��G�i��+@�8�w~�Ҫ�^�O�y#T���'yL(t��:�!����7��G��r�\��ٽ������z��A��F��>9�[�����h�I'��4���D�Kl�QZn��$i.M��]J���ރiEKK�#�%��S�BeY���'A��F_�T��9�ť��(u'���EL��W �Lj$6�ˤt2�<�G+;;�*��	�ӛ��I�v٭Ӗ�г�^Ga}�P�}�S2�'`ȑG<7	�^�{��>���Pn$��J�0��o��:�{�L�'��Υ<.�ߐ<n���$��/ާ�q���_qu�����t��>����O�L(j쯶��~6���T���U�1�.����c_E)[�/n�AԲķ5��k�F��]������B{�Mlu[�s�M�����m=J�\���,m��\��tx��A��Ƹ��ի��*�M9wV �I�!�Y�l�V��?[��Z��諭��\1�]��F����
�Cy�5�C��L�_Cp�g÷�'��'�C*�y�@���3o\E�/3G�}2�V6a�1�4�&y��Mją}wJ'uY��+O�	;��D�� z���^ʛ�1X5ۡy �Ϛ���d.�K��]���m�!�2���mE2���R��tNԹaP_����R#c����������?c^����/ǫ�C5�2ī�GO�V
\]#l�K�U��]7��K%}�o�������bpe�'�����j���e�@�>!�a�m.�Ceo�GE�Z^�*����ڳ^��Iu�Ga�����s�:��#�l�,�(���0U��|MqK��R/C�1�:`�����ݕ�`�U�wY���3_ι��+NldX��F��zm����#{�͒�]ძ!��Ϣp�/k��i�#�Gfܡ�"�Eּ�+�I��7�ͦ��j�K�j@���q���~f4���ԫ�ܹ�*ϡ��6�+>��z�}P۵c�*�M�Â�s��"�S�%���R�fBʨ��:V���vt�{��X乻�q��Y��"�V�,�c�AI�⟬-mk������������7�}�mB���mʘQhA6�,���=v#��ﾤ};�2,�[����F��i���r����Cy�gY�B=b��TI���x�n�u�w�t[���F���������f��:�=U�hά����쟚�[�ZՇ2|~�}����扰٧������%�*b��-w�{�B�Lf{w
�c��֜�R��n�t݂�ג�(e1H��������k]�Y�k��,�,�p]�P��zL�r��R8����=%�K�A�^�`i�V;�����Cf����ɦG:�W\��&+����[���g���۶f����#� ��崬��q�2���˦��oz��rf����8My���H����8K8>���5�v!���#Q��۹���C��$|6D���f{�_|��Ρ�3����M��VW�?2��P�tw�Ƹ{=��'�m��.���?3}�����BI��V���FU�,���+O({��0���f�1+o3����cj|�4�|������ua�y�yz��t�bH��*Fk�;��O��dDM�L~���ɸ�r��L����xt}�׼��?�&������81��]+7�q�����Z�{N��m���h���dzi��P��ŁSz�,z�����8#��bﵺۊ�s
�÷L�W�6p�:�������ʲ���_cC��z��+z陃b���3�æ_23�hU�+�V�@�3���y����V/�"��&U�W"IĨ~]�p}]Y��H�,�K"Wq\� �K�=�i[�����웛^h�t��t��
	�|үa��x����c�e.ju����u���w��h��t��U�CĺG�� ���N���(y�
��nf�y�vF}�֜?.�ݾ��Z�άჱ������E��Q/R��S<�����ޖY�������o?'���Ƹ�5��(}��ҡ�	~$Q����>����ş�N���8���{�f.-w��9�C���] ��!�E�d)�*��o熑�~�*~#�V��K��/o��84f�3n�������Z��ÔZ�u�K��_;]�Ӟ�u&X���}1�K;� �~�Qgd��zf���c���UϠBБ!L�:��'����<n�V�Lش<�ÝeU��*�>[/�����s�_ګ�ݾ�z��,�����6�ˎϷ���]��7��Cv
ݬdg]�
R��k5�9���P����z�f΅���Q,[��o,ڃ��(p��/>/�G��D�ml��If/�O�"&�LG���m�M'P�0fb��816Y�v������.�x����%�5cx��5^itY��y��+kn�+��Fyb�hR�0��e����Β�����e�ɨ��K��Y�m�A���)�]h����sN�m`�snQp�=�]̈́>9�.�\�-�ڶFD:��J�o�Hp��yc��j�ų�8�	62(l{p��7�5���1��/�-]CN�l3�s0&�@Tf�����5>k�Ü�%>���<b]/lEX��洣�>{�k6���yʠ��1��=,���sWL��ЯP����2����y͡�k,%�V'�YU�,�v%��a��g#\�M�8�W�}g����v6��D����[V�\'6t�Hd�	}opW��N<�m�\N�ڵ��D����[���u�q�Z]<{f���8��Z������(�-��-j�x��r��9���M���4<8~|�^�f�s�Q�{oL$��Yݙ"�.wk����U�᝚�9|�������o׺ @}�Ϡ\�o��DSb� �9P��5-z���廛�k&f�(�yg��f�d˧K.vJY�a�}uFl�u��S#0�1��Q��v"��D_gu��׎�G���ʆ��SM����q���Y!dZ�a ����}�M�=����LNTY��7FBw����`3/{��)J�j!z��v쳉X�:�)ո�o�}��.��Ec#4�Ը2*��廕�=|8�U��[j������+1�}i�30�N���V������K���T^L�99��5g�u��G��m�c�>��K+sA��[�$��u�I���%��P����s�o��_��ѓ6Kˢ6w3��@%��Hٶc�u�wX�dy�5�@�˚��)����|-��:��K�<]3�����5�g6p�J�M��v��ѭge����B'�맙��M��ģ*�炡���
��WRl���f�f��v�i�$�G��;X�r��]q�"m[�br�.%ff�����{�0�\�;���S�����]����[ө��x$3H�h&���5�ۛʉ?��#��c5i^���#�d]�b�n�n굋�2�=&m({tG͙��Re�#K��6��3�\��z���T�D=���f�$
�1E�g�`I�Z#2��a5ܲ�p`�
'eٚܜ���c��j�!IIÎV�s���z��t��EV/��}ǢVz�3�Z�e:�s%�y��%u�\�@�Ioc+eu�ht�jq���]B^YN<�]u�
em<Gp'�s��Y��ƙOu���H�i������kS����P�;}�%jT��(���V�͛���n�o�s����H
(�R|���r��V�&����i�ꚴ��q����Q�P��1��[�EV�2�rֳ�Վ�3T�]9��n�T`"c
P֩�̸�R�1��10q��3Y��\��3M3W-�K�f"���9���hi���n�e�9�Ri�+LWA�8��-���\�3-����XV��\��jQҡ��̫�޳SQ��Pա�aQ�Z�)��dղe�+k6��Ve�F3vQpAB��r��n�p�X���s3颮���J��kVhADKh����k�<ޱ��+*�G0̥B�r�\���#j�+Q��&2�z�-��Z��L(�8�`�e��-�S2���-Q0b�4�񪚥WYc�T3*�����ͥqe��A�W
Z�6Q�顪ڎ���7p�Țe1����m�3n��V�i�*����e�\VfX�o��3t4�.Ze�R�n��)��4eue�WLusM�ֵ����R�h��)Qnf"Z�����ʫE�uqb:i��X�����*�V-B���.U��V���Y�2�
V�A��TW+V)ijTi]S2�je��Sm:���Y���V����Q��nZ�j����Qk]b\՚p�sS1�4�,�QՅk�I�`��8)<=�g�|�ו�F� u��f�ք�v�3&�#�)��٥���$��e�(t�ę��m�x)�b����.�?U�i�_ԫ#t�秩�l���������Y�.��[c�-�"���Z1���=[���f�wB���(n{޷p�m�#εb��t"_�e�U��v��*�Bc�^�!��sU�]����r�3ń���;��2�~������*�������Lt�,gҝ�[�P��ݿwH�y<���!�p�ơ��(��]-��2<�á�T��%ةʫ�,��7����|v]�.$�S��*�:��[�d+"1	6����X�|;���`˰�ysZ��׏gpX�i4���g��)�
R��&yW�ʿ >�y[�5hcټ�,�n��=[�`u�*�P� a;B�|N�z�����(ach_g�XC%�.;�⟩�8ӅV��Y��(L�L�(*�	o)b��C�2YcS��W���û�kl�=�^���9��sϕ�ҙ����|%�&�$���6Z��=�����!@ـ{|T�^���I��1f��"�b;%��Sʊ�:�5���]]����������MgK�X9��L�����kƲ�+6�^��k\�]R��r�h�4"�k;Ff.m�r_e��]]_ޯ�Vw��l%0󫶳OE�R����re���NV�G�AG��$�l�۴^�20)BR-#�`�����ߪ������w\S�� �Lj$6�ˤt`v�Puz9�������/��� ˤ�_":��yh��X�Uf�z�X�n��S2� �LWjf�%�_m�ٲ������+����]�����@p?��C}�o�3x�n��j�oJ����P�*��r/{�x����L�L��C�ʄ,�Wn��o��/���O�L<��e^� ы�; �Ƕ˯Vפ�]-q�7�V^��캿o�P��W�U3=/�؍S9#�M#�NÁez�`T�6�ڃ߆�qC���d�3ݢ�4��/��0�N�_^�1�&��wץAw�d��'Y�҂��B�[Hl
D��P�.��y�h��O!v�R��vE�b����D��eRՀ���}�o�BL�L�~��3�瞮�Uu��
�=�y��w2���I�WgK���[e�ߪ!����MkB_�ԯ׹f�E�B�T��͎�����bӏ���^���Z8i�l*��V#��[��i}�L�T���ݾ靴�+%���;���l��U�}��5�Î�K7��j�-a���t o��fg:�$'�����(Z{Ą�M��t�>��y���t�kedd-�I����� �/�|�;�z�6���u�nfa5�er��MH�)x^l�Nr)h�ͮ�uɍe�Y3�<5�`I�|���6�K�{��G��(����Z��+���
�ۣ��}
~�"k��}��X��36\Hx\�b��.����=����|�{������-��=�KK����f��>A;���u�槵=����k�ܡ�"��w�_/O���/G=�x���Β�ܧ�/|P��gm:���+�3)i�.a
�]B��������K�3�Em>C�[�i������r�(�5�pSg�Ϣ�)�y��m�T���1Ι����(�:YA�RHA�>	����g��K2m��4V��{�a�g}.v�ã|9> Ox.�!�HV�Y C��1m��go*D�O%
��t�Q�ɯn��"���.�����R�&j��E�+ F�ϡ��l��Pf~�r{o�Ř7�`�^y���Gl���}
�1�f̴Ϋ�t�o}ݼ���Z����T���bd���}�)�o���]�
�}C�@��k����f<����z��x�5jŧ%p:�o{��O�s/)�S��(dg;x��iWj�}�&掩��+a������r��[q�0����+�)[�ڸ�h��yI��8��c��1�����x0f�z�٪��ݶA73��J�E��R��H�޲�7yc�r��0�5����G�Ǣo��g�3��DX���%QOB�^�q��\wC���A��v�/kO�w������PH�iF�:�LV�S��#�W9�5ń���t�s�,��j9��n#R����C�|�@�O������罜��w�=��3�A�@4�L�R��y��v�l���=�|n4uj��>[OIҽ鯗!J�ڝugR���:1E������ŊW4';{�$�(��`�2�h)߳ӛń�=Te{�]۩�rT
�M��N�㾑B��Bצ�C���W.��\��{�2:ͤ:H�@�5�|(�HpX.��2�>���0�SN�gԆ8�ik��]��5�»|p�\7�ȭ W��������]L�3E��)bo��T�cm4�jx�=���Ɵ?X����8�]��S���!�t!|٨��.g�X�\���І8f!��lU��$�፵|�6O	0|����Zӂ(}�O/~�0w���:�> �F��;�෷b��`k.�v㯵�È:)wm`*�jf����J����q�v��횃����,��;3������[]�`Tcj�hS�.ǫu�*�5�Sގ���1��l���6�t9�ڬ}O�{�[.k
H� �˯��&G��O���r�ĻzzJ�^%���LJ�cڳA^�׭.Uٙ���+t7�>������Nx�=�U`�	(9r���~r�Z/��&i:��+zW�����o����������Ş��
L~c���������1SV�O�����ӽ�1�f����#|%u�x�sh���\O��K�Wx�S/����FI]������q����i$Nw��i�/&:�U�C��;�E�ZD�+��H���_n�	.c�2]��e��ç���c�ѱ�<�rش�eQ��TgUdWb����8�X�]�m�s~����OB���WW3bu�G��z�d��ng��vT:i�[�]�e)�өw{�ۻ�*]��(b�|(@}}E���8�Ozһ���k�.�݊�*�I�wc����B3�C�~E��`~$����Լ s��X�F/:���ŧkk\~P�^���7�.�:�>�y�C
�&���Z��qw��]�N�H�KS�N�^�&��m��/7��{��e�"��p�vִܲXׯt6�OΌgp�靴�r~�N�꼛�z�/J~1��OA��z� U���Ow�n��s���h�ͧC�4W`���[K����{�h���w,�}�3Z2u�Y-4MX�,�eQs���V�*L���}�t$Vo�ƻ��,���`%�0|��㸫�A�cg��<;�D�io��i�^�/��o6�O�ys*�Mo6�D���f�	�@����Ҿ�:q�L�Vx�P��o{����|���zCh9b��ӛ-�@LUR�ʺ��;5U�W�[���L[^���db�.,w��
>;^�0[x#�k}R�ӎ\����J`�Y��^S�Ŧ0חp�'���PB=Y��-/
�/�\��^����'�a�Bb�>���p՜�˷�y��F露��ḳ�i�n�N$]��\E-�GydS��/;��L��(M9T�Y}���\�S��S�oR#���:����d����;�E�/�J:�?��J�ގ�L75k�5Ǻ{�뢣�Q��'~pS$�r�<�%�yb�*�����J>���!���T�/0o�y~���z��򂮐�ϫ��t�VU[�^�����]�+��GC藻���U$��L
���)ڃ}C"�:}�y�c&y��Pæ�Ù/�V7ʷ%j����#_1K�f���뫋��H�R��Si��rV$i#�'��Nte�h�c�7je��B>Yqv��_J�!o�-:��s�m��ZX��2s�,��Ȃ0��Yق�;k�٧p����i�r���>�jG�2��FF #g�|�y�gN�w�sܯ�&�g��2�tȃj������J���rz�/�k�#"��V^�>�dzt�p���å-����/,�G�	�}�7����	U��GrЊ�=G5^���mAm�6t�n3#���Y�<��P��-������+,1Vp��b�'8m���{���
��[����N^1��G{�]C�_� t��Ԛ(l��
%�ʞ�ᥨ�X����}���Pl��]�.P֡3k�>+�It�xOy6�=Wv�7Ư��]oO�����:����b��4�j����eą�~<�d[Cw���g��/���f�o�sx�0��4k��j�R�I����>��'9b/����2c�+$msQ&�g������O���g,B�^��]M=��u�s�2�E���&{��=��zao!�=Zy;�ՑXݚd�n�5w+�7�<]����W�2&�����xT��������_b��׏@j��By@l�<(F��07Wīw�|��[׼C�]���R�̱ ��$^�Ͻ�Bxh�Ƒ���8u�#r�m�mP��2�dV�}�z��Gh����#-�������~�wyjn��]}6�剳0�R�{aԐ�Y�5KɆ��RُT:\�/.94u�B
"K׆8�-��%8�s��(�zm��I������2��6$4�3��uD3�:ɠ�\0��,���}X;��l�M�R�>[���E�)�v7��^ƨ�E��~'>���*��.5�?>����crt��;rXY﨣��J�O�t��x>�Z�1B"�O\���wh���`�K9`������P����%g%��5^+,�^m�3����W�
��3�fVZ���KSˇ�GQ�Ù��Xdƴ�Ä��ҵ�ǥ�8K8F���Ds��e)/M\�}��$ԸM�΂���Flsaڰ֫�4�T9g�$����t�1�vm��_�7��n��Sd�1z�|�̯oѠ�Fl��w�kG�Dx_`O�#�ӣʴ�h�c�oW��蕼t�	�����C�yQ4�����^o+�;|6|�#C8�����U�=&/�>�i��*Y�� @�����u9�̪���\:�dg�q��b]��K�ޭ�fa��E��;��.#�P��9�KG���K_p0ud3�~���	���FW�^���=Jp؁�Z��T�]Z�l�\3#ܴB�Mһ�ZN��`pZr�ɗm��|��T��,�Bu��� ���igaa��|q�2�rU�����ՙ�>��N4�Ъ�S]a��������TB8Z��:L��cd�n���"���h8��[��V(���wp��������5b���,'~���}@�N:<�v��}f��)@�Fw��.��Ƒb&
G���b�DrvfO)C�ΈCo�����>}�o�k��� g��g~ؗ���V"\�A!�fe��ml���{��E����EMF8���Y�=Ĳ<ݎ�iexqh�:uzL���%�>$���<��W��p"�]���?H�I�� H:��+�p�+ѡu���%���J�^�^S�X�>M��`Kپ�q�,�b�>GC����Zs�)��U`�%|���t���xk��(��X����B
͞�W�Ñ��r���z������c���{��S腜�wٍE������B��w�|N�~+ؔ�����3H��^.�go7�;�^���e<Pt=aT��[�#:�v ��U[��u��c��b��]U�����������l�Ȍ�]f�M���/T�6�y�<7V��eQg3�x���"�1x�͛�6|59��X�`jg2���_R=�5:��x�fkLhP�7���t\5ҴЙ���Q�LV�3Ǿ&�DO���6�n�u�M��p'�7"�LG�N�TӛV�R��&�њlƄi�n���'w;�Z�ꛓM҂Z��� �L���0�Z���VWWC{��)�ա�O� ���Z���Q��O�OnmT͂�����}Jm:~�����]��+/���)g]3\��A��+A蟏x�iM��N�����X���d&w*۩��U�,�8�Ih�{��K�9
��l��}Ru�<s��5��_d�o����l��X�
L���x��?�����f�S��U�mHMg��4�mk����K�{��=�g��-�`t#VgڸK5Z���z�'<}>Eh�O_B�YpG��PL���[�f(�z�5�G�5s*�ky��-���5��"��V����:�e/
��^rb�A�9E����/�=��~1���uV͉���[��с���܃���P.󳟛� ����9���/	,;�]7b<S׈<2�ӟ9s�\��PM��j�+�޷�c͹�|sF�e�F�:M/
�GR����OÚ�s:î�.d��THm���L���=��&#�X~<���;���k*WKi����L�������2��ݲ	C��oE�U�mM�Pa���D��L�z҆:]��MR��,���1c�� �]�H�\2����y��Ɛ�>��꾸֗�a#6���R�z����q�ƣN�y������Ga܏p���6^��f�'���I�of��ɰe	���!�c��,v%�̝k�jp6y3t%��ei���{���K�x��Δ�ul��a;�s7}ڞsϕ�K=�7���-�Ԏ�o:��N:�����9V#���\�<�=Z��2��^���h�X�w9j����8�sfU�����c�7���{��A��ArMTV�"l������OE�Y�5׎��ᗏ.v��g��e�Xܖps)4w[-1�j�Sc�v����Y�A�N]k~H��9�^���o����ǵ�+IC��KV=[�~�so��}�.����2���f;1�ʒ��J�7,YD�������dWI:�0�#˷��ven!ٳ�΃��G!ͺ;.}��υ���/��N�h�e�o+��U�vl�|oz�/��X� ���`zE>���E���;:�H�`��eXLe-�xv���mvA� �꺵��u,k%EI�5O&�I}�q�f�����]<wd�HL�h���Wn�5%)�^�"���X�ټ*��.�MP2����d�c�kdS���� ��;kE��f�I!�+�$�>�W+)˭��#Ϯ{[e� ��i[癔�t��CD�f�寍��5ݹ�%VEu͋B�Z(�P�Ĭ��M���"���bɇ �Z�%���2;4���Ƞ!П-��2�pp|(v���t�ȉ�a���P�68E	1�yʰ�M(yS篹 z���z.������a%oK��)�#��%���ʗ���n��cy����+l�¥���R�֍]Fm��S�X�Ul��@P����#0���<Fí��baG��*8Oe݉ ��ю7Y���������H{HD��p�"�naWth�L��Z ��Qj"c�͇�e�vo�x�pk8�ïC9���������mge"�]�j�Gar?���t�S،�ٻ[�R5k��F�R�̝D��ok3#�LKPPJRj�ݚ/W"��Zqu�4�T�*�˫ʹL�ћ�t^��M*L[��3y��صF��L�D{�@�ag+BK-�K�rKj�m�A��Ws�l!;%�a��ᄙ%�|"x:��֊�9[k�QV��Br��+�8!�����Ng5����o��ovq3����N.ě��A���dv�34��䅑R��θMg�k���;����*��
���q=q�͕ռ^��Tl4u-�s��FTɹB�N�̝��S�˨��}�� ٺua�:�t}��'.A�hp�Qe��КS4�2�� ���b�ռn�ˎ�=Ft�{2u�R�G55���wP)�.\�}�zl�9�FI�"��O�47-
ʫ.Y\j�E��i�(**�V�CV���\���꘺J�PҷT����*�4�[�����N�u�����&1�q�Ն
�-��!��h�f\�F�Zj�2�*��f:�3.%TF�Ub�-�㕴Rk(�R�ԥ[f��U��cK]8ceҫ[��b��L5��k`��ְ�7v��Դ���S���;����4�Ъ%|˚��*��
�8[u�]6:aYZ,j4sY7����nar�nbTƌ��[���Y(��mj�ŵtܺ��s)�q�V�bD�����"����-fb]k2�i�.m*ꥪ[_)��2ھ5T\�m.�f�7�je.�q�����%we2�R�un4�m��R��m�Y-�
�Ջj��e-Ʈ��8��6����u����s-�5YQma[J�m�l�.�+Z�<i��*���i-B�A+��5�2�kV��W�ҫD��
2�\E���m�h��(����R���ե��[�p���J��m�ea�B�QR��iDDD�JUj�kJ��H���k/�}k�_=Ţ.�7�@�k�R��kK:󸂅
��-��x���	�ŉ��Ҭ�F�y�	�.r7p��w:n��W~�I�ϛ�CE&f�� ���Iv��1o���\J;/Dы�������|���o�'�ww��r�E��:�UK�2��boj:C��3��o�3x�+ib���`��o����D��L*�mLR.+�>��8����J��YbWv���ɺ�:�n�����P�Y�;ƅ�3z�C�mӵm�lV"��@k���f�]ޱ���v����nߑ��vmA斘;ij�n�o�L�WR��}yyB䃇S0{D�L�wǹE���nEݙ�bqwj��`�YK�IX�1r�\} si{�K���G��}�zG�+[��w��ލ��MY��C�p,�!Vaߨud�ٚ..��Xb��)Ďs���.�����Rb�c͓5�w;����S�3ŉ�+�^#� }V*e�6=)�ɘ�,[u�{\�W[�:ZS8S3s�L��C�r|v:��	�k���@��
�^�"-�7z��"�Do/zK�K��]��3�=2���L��`�rx�z�l����MԴ�G#ɬK�rN^@W)(��e�!Ι��9)`9�廰j��9�r��#Υ-�b+�T��U�%��V�9f�;�S�^�X���g��J�2����@�2�:��i�홒��0f��	ʨ�����{�J���+R�s�+<@J��Z6��h��s7*�9��|V�H#�Ž��˚��/k������q棿M�C��%��%�v�s��b�f����@ƔK*��_�#�ʃ,�Z���PT�a�</;-t^��*�/Z�ȹߍ�sL�*��E	��_<DU�ݚd�n�5�)\��<Y˵���%�c4�W�F�����s��SI�o�X��Ve<D��'E��^�N]qa���f�]�C;���'�hY��e�������]�^h�z���PuD3��M�ؠ��~Z��&�t����f��	��w�oå2/zxR��ʌ�/�<K�8׍d�K���r�,���_e?='���˕��L�|:[�3��p>�Z�0l-3��ji�̛���O�6~	n2�!:�]����:ciqkK����v+z_PA�x%��"������d����J|�c\�<�>�o}Qiԃ������՘�4��5�quHjt��W/��|�yF��kW]�wC`ɺ#69����_�j�p,�}g�$]6�HiUoϥL	��~����CQ.P{�#�a�mq{V����ҧ���a����[Ș���^̹E����ַ�3Ɓk���i�+'=����5ՙ�QY���Ɨ�����V�zt�qǛq���v���������	L=�A�n=��@�qՙ��,u�wo7.��N$\Ԋ�D��!y(�5~�+�0|�K��+��zCd]�m�L����Z�׮���w�F�/~��['���u�W
�"b�X�P��A�@4�Z�W������n���O�j�f��Z2G��m�=� ��.�J�!k&bW��տ���ŊW4,N4;�RY�	(����Ro/\����:��i�,�z�8.�`��U�n�t��xl�k϶ߒ!a��Ԫ�M��]�jӞY;�A5V<�ώ��L*=N)�\ҫb�H��4�p����z#�?0e�3���-9����V%%�3(�0R=n�� 3��:�t�B�>��ok�=(��tfd:-��x+�x��2]����@�l�KՎc�{��1rJ��ǹu=���s�"ؓA��x7�K�=�����C�F�C��K>>$�o��W���}��{1��[�� ��y�!ߜ�g0���J��TpIP�ׯ;���5V��nd�9��W��3"�2��;i�Ӟ9OGr�s;�J�9r��3��9�F#S2���Py�1���wA��&݀$;�<�t%��ᵥl<,\�������Ȇ!�Vz�D.�E��mB������]VV6u]-��`�B���em�%ll�,��&+(qJ�^��-6
�X��6�E�ǒs��r��@�%}���ھ�;����g�P0����ᷙ��i�G���f��5J�KG�y��K2����V�s:Lg��%+�:}4���v3O"�پSL�3F%���x���o�E��Sf��=\�}2��֥U�'�;�|P�y>�!��Gp�T��F��{V�Jtw��'a�������#8_�5��«'����t"}~�Y��l+v��*�&;����k̑$�]�1]�Ҡ�!@�:��(+ut0g�:�Ja�hfS��/¯��=f0(hqI��1��3�S��P�RXϧ�p�\~�Nm*�jaϮPp��J�Ǣ~<i�\����q�=�71��J���a�{��Ғ���Uq���Y6�4L�O�Q�o�G��mH����$i;���x�;��j��A�J�M���1���=�J\��B�^��%߄]�7a�k�,0���T]=�}��j͉ƻ��C�QI�6��/s]ˮ]�Q]�yU�Ӑg<������^�Cw�a��˙U�[ͬ�m&"1�f�*+���w,̖�O�"]���ԩ�/A/�k�m��"m.k�V}�8cPxi��뛕�/բ��J�eot���`}u���|5G8P��t�6�Ŷ�}8�Rn��v�ʽ'�2ޫ�yϻ�_ۍ�����F�=�Ӝ+���-�yn9:���k#NCƎ��sǕ}~*X�ܱ����-��:�2���I�=9��$&*�P���)�佶ڧÞ�\���(���"M!s�a³�Pu��3���1f��T����T����+V��xM�Z�̽�ug^0m��)ip�du/@{"�����gXu�๓�j�h�ѷ��S�ú�+�M^v)�䒑"�p�N�>�珷��0ن06c�\!w�����w�3�=N�SI��%�)f�$�It��f�g�!��������1g/Mz�����B�~�o�ޞ���Y(�'\�>��9�u�3�r�z�{#еqK�6��v��/7�<D�r�/�f�QO�u�4k��)���/V�)W����rS���v}�Y�n��n�>��QL
�o��x`���
�!�&Nl��g���%�t����S6�M�%f�-ZN�S�^%}�)Z�()�-Ѓ<�p���A�<�F�t��bh�bT��Q�wcѺrf:�`�YK����R债��m/x�����Zuovk��q�K��2?�5j�AVۺ�u���6�!�+8�6p�p&��I��v�U���ͼF�)IbYV�3\�[�a3��E���J��+Q�5�<�|�B��u��T���0�y����7��wc�1[�WnThs�F.L����5�����D�Ӏ,�&}x�>#���)g�R���p)�^xɯ9yߖ�j}ɍ�H��Pd�#���������g���T�:i�p*��j=���/W;��/S�S��|���r�/�(ZXg�L��<5�p)�|�}��	�k���F�w�Nz���5��~�����UC��4��5��*ꛭ2D7�!+�E�j��p�o����绸�S��.���
�������4kG:���;�.j�+bϵ=C���F��i�핪ǲk��۹����S�h��W) ՑVݘJn�8,B׸��SO`��Fo�`�Kx�^/��R�m>��[9���!Vb(LVEg�٦J�r�ĥryř}V/w<���>�kl�V�-�b��}Q']�X��VC(X�X��$���%�����^���{�2�Y~�s�ݞkK���6��K{��R�.��扐���Ͱ�g�I�r��[�~���9G7��,���7.D/�z�"ߺS"�oK��5G�^�W=Yc�Y=�:�e��N�n^G(�jѹ�E��&�	��N�[�e�+�Q|�(���x�AV⻉�2f^$�ǲ�r�$CWm[5v����V#��C��#�m�ӻ��5QǅsYx�bqޛ�����]�=��q�=�$ʜXN����#��QR0A'&#y�����X�}��q�e`��N����l>���#>�D8�}�&+K�n
�n
�������ͱ���ծţ(AS�%�	�*�K�<=�y)���3kA���Es��nN����ǧ��Ĳ+kR�&V�m�+թ�?]��+���*��Mn�����fu�>���ɘ�=�lԘ�O�P�j:#c��Xõmj�v�7Y�	CJ�t/�G���o���2�χp�PU���[�fs��;�1�{�U�3��F� �V��x���<y�)'�ŷu�D��Ɠ*
�����ʇ<���S����Nk�ڵ:��s�폽$�)�ٗ���z����,g��W��S���BV��a͙U)gC̅���'�C{|���
���`�,	�(�Hp]�T��P(_&����!�;�t^(�>�d��v��V�|��vnyB̊��:�tU�&��@��a}G�Ö�uPpѳ��d��]o�{��x��ǹؠ-�>���}3��Z�GRd��4���&
G���,[�C�R�2}�{��;��[ehm��.���{V�[yF�
��������dk�"�nWf[O��yֹ��e�՞>ʱ�Hn��Zꡍ�o2OMv�ٜZIU��@�Xӻ����W$rr�����6�4�b���ś�G�K��e�H���'sƦˣ3վ\m���}r:���w��S��>:�� �٨�*�Lwj�l�7g��zp�,_W/��g�ؓA���R���C�F�C�1U:����V�Cո��n+ʪ�m������$g�nC�˦sI��9wy�3�z�C^:�SzzWhMhj2�o.2���NM�x�#FֽI�e��_i���u
c�`$���z��L�[5�1����I=���ctZ�n�����zyK��H�A��y.�޼/��P�B
�&��b�=�Ƕ�Ͻd�l!k�R�K�|N�+ؔ�{g�P�C�:��u�M��u؎�j�����8�.//4���X�oX�E��'W��
w�����Luҫ��1��O�g�/U����z=X�bO��|�-�^0o�<�3v���Ղ,43��,�n��4�<ٜ��M��[�E�X\N�)�6��h�T���Ɣ���e?������Q���72�u�V��밸:�	���3Ғ��r౿gRκf�A�����s ���i��O_!�uN⋾:����nV��BJ��f?I���[���%�s#|{�=�YQ��˿=h�*(S�pCp:y�E**���Αp�@;��6�l�W%�Fbb��y!u�I[�$gp�݄`B<Ɖ2�Y}�$Ziu<�k5�r�S��kQ���8[����T��;�Rn�O��*���t�m�	:-�2� �:��Esk6��P��_��b���jϚ�@ꤴ�_Z�h�? �fU�NmU�W��#}���&��O�R0t+c�k����:�7��]�ĳC�#I<�Rآ���Η�}Z�7$�|�rxn�K�je� ��i�˙U�[ͬ�و��&e&�U��'�oNS1�#'�vX��E�n�f��N�P�9�L�x�&i�*Oop����:���8`�4ND�?q}�
+�T�qK݈�)��({dw
�u^	�ɼ���;��N� �X$��_]�ePtB�W��e��Xu�����F��>���;ӯ�8mP���}ʻ���>�����f/-������G4\��a����S��aַ֏.0{�S2�<��LV}%�)�ï;Q%��f�g�!���w�QP�������3>}X���K[Ҩ��\�W�1�\�W����yhL��!��v�+�neo��9��mS�8��V��
��ı�7Ä��yY5ɃX+1)g']�n�X�U�g^ꇲm��q4m[�**��Y;uH��Bb����6e��件 �W�;:��+g0����RȘ�8�F�`����T=!�����6���L=�K{i>�d`R3���v惝��E��o����Pȴ����q�0��Kz�:&�gQd��y�LS��4]iv*�Q0�k��o]�sn��3qC�Cz��d�����\ʮ7=��kbw�Uc�d�wh��9������(�`�ِV�e�z�8b���-y���d����{����{�m�	u!YpU��%c���G���^�	T��m���/I�c7.�ӵ\��M���D�ӟ,�&�aT:����>�/=�&5�w;�3�#�i���Q�lg
q+�jo�߹WbӀN59Cw��.C�,4ө���f֞����T7UJT/���(��L���T3se���2����[g&Y�a�,��o�ձZ��{^�p����i�$G5ｲ�U��m+��76\H\��G��vU"O��$�{����oa��ߑ����D�J"y8����9sp���l�YQ�����vݥ�qp��}�J�vϪ���?��2���F����߮�/��^�~?n��B��`IO� IG��IO��,�$ I?�B����$��H@�P$�	'��IO���$���H@��B���$ I,	!I�H@��B���$ I?���$ I?�	!I��$����$�H@�}��(+$�k1|(�  h��
B,��������S����מ.� Hͅy��Ρ��
VfP �`LM&L�LM2100 4R�dё�	���2�F��%P   2    $҈�d�?T<���h4    D�#S�S5<��4�4@RDS�jd��e'����F���ʨ��{dI����R�VH�$��a��V���1HeP���K��n��QO��%$����O�&a
�*����),����[x�I8)#(T�iPcH�!eI�R2���������*�@(�~?��O��/�Q��T�d�h���M���� �}����,I$�$�'jϲ� ��wL ����z4��t*C�ќU-�01j´�:b�j**���Q2��)�7�&b*�:�F
�eNI)�$�vzɊ�b�
���N�eY�N�3U*nncZ�%cR$T 	��pH�A�P��Ó����7�����l�{���2���1;�ϝ���ƴ�R��Y�ih�צZ0�ǇX�h��Y�d�쩧���U\�T�׆���;�YiTFdf�ek��B+O�bTj����1�Da�-m�9&H��Մ�Ǔ��q�^M��\�46O�B)y7W]tۡUz���V����0$�`죽�@�;� �^;�jT��D)l�pӨ�XZ�#�P��b�6�Z�"�-qq0�l4UEQ|��QX`�b#ʎ�$1�]��[��t�����]Jz+M��P%��6�:`���4�j1�Dצ��v�D�>3~!g�)Z)a x�~�&��އ��No��+ U���=Nb$��E����V&"�ɰ��CFu˔��}T.�!TD��U@B!
 ���� ��N1�.ТZ��c�0�s�����
�V6�)���ާ�A�Q @����_��G	`(!Մ�.���l���\/�0R9�+�s.V�2�@xl��5oB��BI̘���T��m*��p���K�%+t��n�b%v�j��������X���I]�C�੟#�}�F�lL����:���=���g!�� ��v�w���\��CP�T"
TD#�3��d�o/h\����͌�^ӊ Bʞ�^�N����:�5Lԃ�)�� ���r��۫���Ğ��v�����7�)��eIU������t Maꇓ�u;�5���ډ���y�,�<��'f_2 G ��֫9޸�ʻ��zfg܆e��k[�d���{ک�qP44� �z}霎��h�v!c۬���Um)� �I� �I���1���\���݇��Mԫk
;��y�>S;N��A6�w�Տ=OG�>��WgFX�����n�3���q�cw�-ٴT�+��`iv�m���n�\q����n��37ya��/k>Hi�"���a78f޲�=���1���3�3ɉ�"K麬xV���{.upM{ճr��/qZoZ���F�������.��C
2"�M�ً�7!5��9���r(>�L4Z����fW9�M��h2�����n�"�T��u�%�f1�A��Q٬o������"l.�������\F�
��m�M;�Ef�Wut@[ԤH�3�tڛ3���=2NI���ٹ�W�0���f"(l�ח,�6g	�7B�J<=2:���Y|x��˽v:����y3h�%�7l��u�t�!�'Upb�"#5x�<���F��xS*�bb��t�T��'ߑj6lv���j�|�\�WP�{���)���BN����U[�8�N�@�ŧ�� ��G*v��.iA#vuFٶ[&�o͊�w�q��ر��%�GnS��{7Gt>""/Un3�u��6�I��\|ln��eie�Vg�eK�[;�h�a����P�ө�:[�3Pf�t�b���ֹ��e�"��4z���`�O{����Z�U�hH�{,�z�=�H�sAcG�TR�F��.�����׋�Y��EF[�i��s�ji���vsd�
Kl��3��8��l��o�ͳ�(�]rgT�[E������vq�(�1����,��]1
�a,����!zP4=�e"L�(���Y���"S��N)V!P+T�����k����׷Myp���:�$��-�]JZe&,N)iĔc��"���O�K� � ��`̨<���T��L��L��4tƼ��AG�%�#���͆�/��Ⱥ8PP��-��(B�B���n&ŇA�����#f�X?B��tMߖ�hjʱ'*�:��
sR�����)R��.T�R�g��3vL�1R5K�����k$�B�
�˿ִ~���_�*�X����vpQ�;��s�*J3�����vQL���������h ����Fn`��D��΢f� i��:b.�R�"��b�1b���4�6d.�4<g����G;(m֟����е*FKY
�![l �b�Y�x�t�w��8���&���#Z��{|{����!0rR��5)���Z/�1.,�:��y�4���_�#*(�q�����􉵓�Bu��s�]�ύ7&\�\sC]�\��#�ֳ������{%V���d�R>����f���w��G���j���I5��M��)*�n�>IEgS~#F�&��S�%��qթ*Z�*��` �lTG���		�bӚ襥U��q����K�X����bč�`�&M�!&P޽(�����(�L�Xs@b�Y�UeaIf)�p��]����/��5£%�Ki��	��g^�"C0Y�x�2a%y��2Sh���22�(�I�a�8�т5֨��1�8��
�of�"�v2��o��Zjs���9�u&���>�0�F��i�&��uҋ����J'Ki��u��7�-��s@�jz�yzXs�bU�r;��pq�0JQJ��֖A���F�S�H�h����Қ��#��hpM����oF������9�#<���f�K�}�%䫤����XnP�8cC����R�H�5;di��s���*���9k��4K��8J�݁�n�H�w*r'A1�UaT�qqnQcu�&f%CE��R���{��تM�6K��ѫ�%�Z1Fl���Q٘��5���D�H~��>�y�.<���Ď�=g���s9�N���'��v�1I�bn3���&F8�Ȱ�%�����+�r9�S�Ţ9E�ɉ��۟���)�ŗ�0