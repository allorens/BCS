BZh91AY&SYժ)���_�`q���"� ����bG׃� *�  ���ѭ*��d��J�XRB�V�"[5J��%%P�mi[hP���Qj�j��$%L�5"�X�-iUI	IT6�H![6�X�|�欍kSMF��iV��m��J(ْ�m6Um��R�(�mV��hAIV�&Z͚�1�Z�YKjͲ��ڒJ�Ҳ�[KZ� �ԥ���E���ݖ�3Vf�6ۀN
t�(��j�lh���-�l֍�6 IET��2JՅVѴ�D���֥��e�e�Vd����e�m�yw)��mH���   ;��R֍�r���n�[��r��ݵ�]�u6��2�[��9 �m��Xi��k��j��͵�r�*�����F��Tv�a���l�V�е�b
��   � �U ,�PR��Z�p
Uֹ�  h6�q҉P�h��8 ���`� ��;.p9P���h��)����=�N��J�Y���m��kU�x   'w�ITP\� �7v׼��oS� ���;��8@��{Ƃ�w��oa@��e�x�@�=��ix��3R�bٖ�R- b��   ͼ4�x^�OA�=i�;��  ==�=	����@R�Bݳ�z���q�� ���N� +l.�/o�(
�G�轆�3�Z�(��Z�P͋dj��   ��n�
Vooy�t�T�wP��
)�`�PP��g� �R�=�
 �=�E]� =ú���F:�C@à�ISq�l��m��խcmf�45W�  x�������gR¨ )n�: P�.]�@( v����n�Y��+��� ;.v�B � �
j\���m�����EJ Y�  �  ���tƴYӇCA몯xw:�t�k�sJ t']�  w��]wS��v�4Z�^�:
�� ���m�ƴmiQ�kZ�m�7� ��(�'v8tУ�ӷ h�� j` �ÀC��ա@3:� rۀ�4`��1�5��Ս)��
b�Y��Z�  ���ޮ� �� N�����p ��\�Z� [vۀ �s� $�;�A�W�Z٬����[m��<   nx  �1� ���к2�]�e0�T���v��֍hwS� +�p� n�*���        S eJT�F 4�0&	���1JT�� L` E=��S� �     �?��CL C 0�M0RR����6��#S�hڛPѓɨ��RJ� 2  �� 7����,��C��������r0�C��N;v�۞=s�w����^�^�*�]�2�U�*��āU�~O��*�_��{�������S�%T�ߛm��z
�U���>�B���|��	�G���',֮Y9h壖L�f2������NX�d壖W,\�֜�3+�L��S29��3+��f0���&e3,�a&�&e3	�L�fS2��p�)��f2���&d3	�&�fS2���&a3	�L�3��f29��&e3!�L�)0��̦e3)��f2�fC2��e3)��fC09�2L�a3	��fG2����s)�\��.X�er�,5��-',L˙�fBl�f0����r��',9d�,3!��g9fC2�̆d3���f2�2��`3��fI�h壖�哖�-#Z�刹b.Z���d.XF��Y*唜�W-*r�.X���dW-*։�D�eK�%r��d.X��P�j��P�eYSX+����.X��*��K���d�,#��։rȮX��B�jU�%\�,KZ��rȮZR吹a.ZE�$�jS��9h�i,�Qr�.Y*��Ur�ZYUkH����W-J�j��
�jZ&���媗,A�UZ�rȮX��X+�(r�W-Erʗ,Urҗ,��5��eU�T�!�r�����k@�9j��Q��rҫ��\�r�Zҗ,��W-
��9g,�h哖�Y9a3	�L�f4�fC0��̆a3	��f2f	�̆d3�L�f2��g2̆d3	��3��fP��fS0��̆a3!��˙L�fC2��&d3	�Y���G09�̎as)�L�)�L��S09�̦e3�-5��-.Z9d喾��~���/��
�����￷R�z��cdZ�CJb��b�Pl�.�3w#!kjJۭ�m虻�������{k/�Kr+�GW�h����ǀ-
�j�G��4����$)^f�A��q �撛kMEO�%��*aܐ���5ї,��X�3
��:�L�h��sh!��rLXUʹj\�*k��䱰jl�[l���5�X̄FҸ闳mP����5����Ѧ�ZD%�y��H��S[1�M����S��c�j���h�g'W�1MJ��[+��4m�JfӲ��2Y�!I�6���H�5�� ��=aZ\�՜��є����{����;bi4�i-���L��-Wr��o[6++(P 1Q3ge�����.��f�)�Ѣ1c�LǢE��`<�M5�t��3aH-�\86�iH^���z!85^i6m�Tˌ�Ș`5Oj�,�6�FMac�&9H�����JŸ�8�I���ol��0��Լ�kp�Q���Qƴ�¥E&M�h��bm95���̲[�ˁ\(�8hn�嶭�^�o8���mǸ)�X"��]����u�b�	�#:�d��!�z�����bQ�1���X���'�n�O�1*�0[R����э� Z�ݙb�
T�]Xtq�y�V�55��*�9�.��9����)�,�z�8˘��`�yפR+��THw[*i�Q!f�l�SJ���%�p�+h�0鹀Î��$yb�+K1��4D�֮]�h<��� B��*�r��*Qv(ڙ�ÆP�2�]��LV�\6���k�_�m��7D�zD�f�Y�%L���M��[��G������ul�.�Q�Tq���Q�z�X����TIռ�syY)�٘�i�YEݒJ�R(-F.��S�9�D�B 8,������r��x���@�H�pk*�\�gal�W��1ǰ��`�X�̥z��60��kQ��3e�����xҝ"Β^-ܘ��*�.]�ƙ��	���=���"劖t��И�.ڨ�eL_*Xv���Q�2�wl�6F��K�r�h�1-{�Nh������[����-��T�JʡbΛ��.8U���b�ʂ��B���̬��2J��,�'hQ���#N�ɀRr��:�&Ya7������s%5C.2���x[/��Ɯ�Dͼ�)�O7U,Í���YWn���-��[5�
�(�zV��Dխ�b�.�i��le�4J�[f���EM+[�w]*E>�-��IQ�Ii.��"ɛ��)L����`ۭ�*:~�\���-�pX�n��Ն�m��S���Eb(mJ���A��O�*ԩ��5`�3#�n���G��o"�6�n2�U��hI�#)$��B�4�8�"�TܬFaW�o,b�8�W��t�g�օ��j�ɚ!��N�Y�Ղ��e�/��w�7�0�U��0���Ptt����W��q�An3I��	R��ۅ妙P�jH��X�x��ө���%?�^�l���X�d���V�j��۔i��c���Z��b����1���j�m-ٻ$��Di� ��j2f�v��b�N������A,f��Xq�;�x��5h����t7���b���_G�	�ܷ�m^^)(�Ct�E���Q
qeF5%�mL��E�m�K^����.)2����K5�cD��l��5
��M������2�nCR��U��x��7Q�N,��z���e�Z�ƫp��Һ]��^_a �{[�
���5*�!peڬ0���k��o[8 Ũƚ�9R������O+���ic:�9���`3I�r��r�M�{4�Db��*�9���u�S~�Pn)�3wC�C2=�n��k$.��#emlZ�AS���˂UVf<DEw���R�'.���o1���S'Xҭ�)�W�19sA�^a���	UB�s"��P�:�B����\ȶa����Ѡ�I4�U�6��mL�&;ט���|�dXÙ�|�����PM�@鸝E�uZ��H'D�őI��Q��VC*��Z�3x�d��wN�L`�˻�"��u��[(�o(���nf�{�	���)�I�g%�����(c#Mb,��u{xh�,�f����^�i�7V1[�t�JJ8������Ն��A�ks J�:����<;���^�hy�vf���rQ��At��4�1����l��+�64�YOh�Ǭ�yq��M�l�#uїA���l��.�(K��Y�OM�Pe6%��.�^�ܚ�I;$וc6Ω����.�&a�[�J�B!J���Cb�rጢ˳V�'�l}-�y$H�����kf��-f��ܯ��A.�����d��<y�(!d��.F���۔�*⤵^+�܀i�n4n�y2�W�^��HA-�ME�e� ���n]�Ln�C`�C��hk�25i�Í�QP�m
KMe]�h����2tX��I��I��Fo�,f����u�r��ԭX�1T���K�D&)X#sY�&E�w���7��6���dJ�7^�a���V̫���^)�рa �lnCX��TNc��ù�ط�VC;�oF�yn�W.�$��mi�e`Ctc"�衙&^V\�f�$d��%��ݘ�*ҫ�%K�w{��A�ju�l����ڂk��B����t���+j�"�ɫ�a�Oq�r�7当P.�;UZV+
�;Fӱ[���z��4-���U�e=dN\�&]�\Ce!Z���C2�������i�T>ThMɎQ��cX&�Ò����=r��1�o�����{���;�M�N��++K����cV�,Y*��a��1�34�9��{v�Ŕ��m��TG e�4�͍�d��B�X]�NQL{���p�(QqEr@�f���Ȯ�f�e���4U���N���
��L��<�o�Q:5���oNe��bGI�.� �ni���@��f��(�|L1-��F��ͪ�53c7.�iCv×	�d��V�`�hw+b���t�c�b5p^�b�wQ�q��ˆ^�C��I�������c�è�B�����ʴ-b-�M��ݖ�HգʷhŌ	�4n�O�����IV��Y�#&���V��sv��;�D�Iu>�7��nШ�.�x�r���e:��SF�)���\��7V�=��nΗ2��0M�້n�K5�M�7m�ʒc�
elݷ6�ݦ/-]VrM4r��j�NKB���YcſnU���Jy�8rʓ1iƥ���Ł�ks��v��ue�5	�����&̴L����;��ܳ��L��5IL�sA,O v0����Ȭ�����dը��!����mq��{a��=�S���H�Pr-��p<Xdj���Xt��w���+B�i���2r�a֚
�M�elA7�;��P�ÓZ�]��0���[�Õ��4n�
��]Ga�.�j����Z��)ӭ�TZ��Bj�0�͙d�5c��jU^�Ks��Z� �2(u�ș{72[B#1^�u4AsvI��4^���Yā�������׆:���%+��
-����R����hy�{s^!�ICi�m�Շ fD��`�Y�Gꐒ�V�$�ꊠr�0cWm��I��y�Z@���R����Z���ʢ�>A�2΋טM���g[L�4��XYp2��j��D�3PC0��[�r�"�mFJ�AA�;&=��7�+A �:�0,Rk˻f�V�<�`5Y��{7I�s%�Z0V�S64;��f�ѻԭ|q�OQ��V]�r��[On][��-��1��!oFԱ�d���ZYx2e�&C6�+���l��-!Ф�l
,�0m`��̶7I�F-���#�[D�ڀ��n$½fd�oke3[Q�#��)m�J�<&np�8('����vAf�f}��#��po��Uq�uU]���Y�҉�Y�h�3za�i7~��SiP��jRY���;�-SvP;F4�YF�S�����&�4:8PAkZNG���+#�p�44�r��l�e�b�^[�v��=ܫ��i�����ˑ�M13oh�5j�	�TF�n��M�� Z�a:Y�,���ڎ�m��,�����Z��B0"wlҢ��u��fob�yub���%�u�KVk�z�Q�R5*��a��í�u��Q`d^��fe�4͢��u���kZ�����Øe�o&.�,�#��1J:�5���eY3wN<�X�9wb��4�#41(P�ٕ)9�������d�:�����0�V1�&m��]lIc�&=����4�H����gQ��m�b����*T��q�.�1P���-��K�� [��04�H�������m#�@��.J�n����ڂ.l���b���1-��a�8j���u��4,,���a��fG����V�-�ʷDMA�KPJ��b \F�@���u�5�`ۼ !XP�e<%,�53Lp��o6�[���P�B��ۅ�j��jm#�R�T �dg��^�u$�Y��W��Lؼpb.��UQH/+4Y2��j���Na�A;/�T�ݤoN�߅�bl���S\��:uQ�b��Z*8�{H̼hl��x6F��Ź�Q[/E�5�I��oH֘3.�8�C@�t�M\��8�e�4�%���TEm:�l4ʉ�F��r�/�H�IP!�tB�h��ٴ�y)<:�^�W�W�싳��[�\Zo3r�k�����9�c��S��>D�u�P�2e�f�%-[�r������t�v�Y�$��;NgfF�&�܀E��8U:W���R���7b���������M�7ћ������|���	��ʴ\�����ˊU����(�L[2�9n��+b��@5���hUYwnDma�/i��/1�r�,ͤ�B�)fjz	��?�����\�ˍ꽥��Z�l�Zo��[D^�1�OL�ܙfH���3�!�+���r�m�0^��@ʂ�������{'.��%GJ�v5��eR�L+1����HSf��m-fE�G�#�ʅ�V]R,=l�	U�	�����0nY٧+)��uƯ͓�Gj�ɘ,�)��]��mx�c17y.^G�{ȾZ�哅��hdV�P-��U��`-էF�h�M)��mѴ����V����CQ|��D��E�u�HL�U���4�ͥ*�m�PkBe���&�M���oV��YS]Ǻ��zF��rV��h��BYFV/�c��E)�!ob�qa�tD+h�� ��뭛2�ȑb� ��2K�`��H���e=�Se�11��F�a���u�V�uEn���ZgƑ[��7R�^嗇vP�)��ZPQ8�,m e��m�J��S�X&����zwDd��ӆ�cں�)	�u+��nfR�����V�nE��픰,�4�[*���T:�N�,Y:�<��;gE���\y+�(H���*�ۢ��ͅ�i9��Z���ȯ4<�ڻ5H�E��t�
ׄ�UY�40�j ��m,��!�*�a��X�Ӽ��ʰ�
A۩{!�z��v1Sb�)��N�$��yei�r�n`�*�y���ҹAJ�gk0��^,lM��K3K嫤�2��Ѣ[�]Ќ�8�ƦP͑�(��c�([jv��ڡ�F6����#qjyxUI�X"�T�w�2:�av,R�<9��Ӛ����P���Swe��!�x�:D�\� �kx����/��(�V�"����02U��4%��6V�f�B�VT��ܙxm��-O�ej��V*f=�8bt�Y��Uz^,	��˷6�E���fchfne�i��wkD�.8	�5j�����qT��6U� U��VY�m�$:�wm�̜bMMk0�k#��^��3u]��x��V��6[z�a���M�0!zE�� �Ap匁ݺXv/h�u����O�#
4��LH��Rj{��3x27I\x�e]�w 3C�̼x�vb/n�d��t���r$��{v�߮m4��dDXƄ�X6PH����6:D+���V����IZM��M�����r�Le��N��[3��k�T{��V2ȴ:7,�n^e�mm�&�)c�ie뭵�2���z1�?�պ��Ù�S#:���(�4�n}��#�3l��$�Wn:�mr�Zɻ���;�}�؝m"��f5�q, �H�=7���^^���\��K�\����2k��ܫv�hUl�z�M�E�ۣl���4���ǧ`"1���Eu��8�Qr�Q��6��k �Z�eS3nA�Yn��j���b�N��)�7����y[�N�X�tL�SpH�����ss��cK�lU��aL�m�:�^2�T�.��[4e����zw~yU�-KƬ[:F�v+S�p�5�T�;����w4ÒJ��J��(Bb�M֌j�CT7qT[�7E=�gA�2e港sEb��^���vm��-Q�j��i�6p4&|� l`��{���f�f�����B�M�I���V[�-(3	̀���IT7�.��ΑD���A���Y��f�dk�5+M��6�W0���N���
l(����-F��]�/SA͢���u���XLbM��Z�����L�����yYF�n�X��NU�΃|��+ ���	H0u���t��Z�fL�"���+��{P;(�a�`X��X��`o��d pW]a�ܵ(W�䧼hE䢄$�/��<��G�?�$�0z�����F�p��{^ ��_�0p�p��C���$(�	�sH�_U��!.�p��͖�0��H��D��6^F��C�B��1n�r�	������fE���䳮+v����:�N�3Ʋ�bR�v��ֈ
7ŧ���w[mncod�f�����4�"�ەC�Ɂ��8�1��7'p+<`��80v���54��B�isDk?l˩�Ѹ�������#fb\�T��T��[������j��������z�'�0u��;�̿����}�}��kʁ�T��iz/������v�{���i��;C|r<�U�6��Ī��i�E�;uπۙ8ڥ4츻���ѻ�.�S��U-q�׊�b
|�)I�{�+t�2����5�b�D5�urKyں��-]��&�\�NQv�\iHL����#Ot�;��B%`��k(J����D�&�I�3i��hb%G�������R�:��K�Ʋ+x�J3h�c���BN\#�5`���V��lUH����/��{;Z� V^���8o-*����nC���>Z3���I٨	�S.��_] �Z�[���SrnG�/_Z�Y���Zm��M�B6W�U')���1P�)��=2�������,;o�t�z{�%��t�2�a�ʭ��,v�j�r�]�#Ӯ�T���Ei�0����9�-��ڏ��W ��n��7�e1�6S�Aҫ&��7�x�����7�4��ٛyٗ�dYn����u��[)�gn�hܢil]�{�w��A���P��*7]�Τ�^��F[<2���;[V�/Z���=װ���|�\�zGH�Wl�V1����tM���wgK�
���Â���$��j��î�;�>jL�n���gX����sJ���s��7�
�+W����{���[�aZ HCE������:PX`w�ikN���/��﯑	u�,�/0��f�t3OX1㾚Ĕ��:]�xl	��+���wzI���.>ͱ)�}�ֈ��j��sB|���"ʛZ�:J���-�f�ᵡ�U�;%,�ߗ2f�ȃ5k	(n@�M�i�&w4%��,s��&�*�۶�pL��D�Q�EH��k�vE>ޫn�T'D5|����(Ww^u�#���vK�dV���Jk{�r��(�îV��C��h&��"Xy���������U�7u�Δ��2yF*�7\9s��sd�����u�>��}�o[�Lո6l�;*lmq.@��qi��Y�M��d���;�L�w��:{�?����0i�_!���j�.�)��[��'�ެ�$�S-ج��''*�eB.2��r5Śx}����wv���ڪ��&��k9�G{_i�˧Q(:n\�(�|`א���j�l�\�S}��%J9[�������r�T���|$9���ʾ|;�%0{�0��/g;l�P����F-f���,�77Q���8_6+��)ꕻ�c�6���D���	9mF�R�7+��n�����%c*�3N�(�[+R��vq��$��Mg��U�y��9L��Sv1'l��;̍�oP�}̱%�7X�a���8]k;b�0u�f��:G�F�u�O�J�������j-0ƂO�T��OZ�h�59�vY�$z�j��v�	�{b�͕-�\|KK(mY�n=¬	��hV4�k.L��JacWn-7�ek�R��Ѷ��F��ձo"nq{�&��M�.��Fr�%˻�I=�*�!q��U�]��-������q2�»{s�I�0j�%����F��U�J���7�Ŗ�ݤzIB�<����˾C>%�e��ԭ�-�8�nj��2y�۰��w�;�g7��r	w(.ՇJ�t�vwW�f]\67�KJ�!�4)��Z�&徫�������A�K�gLra.������]��\��D��y�ܓ��s�[i'���p�f���0I���e�&dA`���S
wmJ�P�l��CÚ�UP�.rx��+E��h����jIHP� �1���E=�Jp�h�=�"��N�̧X�G�3x��%��ˍ؇a��*��;��򬒉�������W2��#��w�eӁ�	+0^B�����ך���F6l�1`X�+5F*Bh5�m���^`n����v`�}\�`�[ѩ�ܻjk$�kK;����ݹ�Ԃ� �<�c@U��[I,ڶ�e:�������5�+e�m��M�xۖJ:)C���k�2Juj[����,�+��'�	����Oq�k��݇SK�Ή*�z�.ʔ{	���7W��5u�GkFX����8��%F��V���)���n���x\#�}X�K�R��)�U�N.�<V�Bw�cJg{E:��-����n^]�q�݃��49�w\Ƨ1 %�{�e��t9.	k{�P���"Xw�^��R ׽��x�ل֗"7���v�\\+;��7���X��B�=�^D���{}�b�`�m2N@6����0z��x!-��守/hei�f�$l���ڍ5�|�de��XW4�g���RL���垊IۣM�=����r@����;6{7���Mt�ì�k0��,SΗ���w���©��VT�PNN�hKqA��̣ť�VX1}����6��bE:��R8`�(�Y������5r�U[Z�Js�����d��e�I"���(NpҴ�)��R�t[�/�$�2:ha���YKB��վ��#.��x��ޣ��dSǉő�=݁�&�*�/�oC�9�6�]L�8�^�����X'.��C&FgbX�q��б{���`�#:�2Y����qq��n`�	�^dU��كj���C�u�.��{�Ď�`�7��8�uL�\w(��rw����G*:RY�5n�]�l0�m.1�t���N��Vk5Z�*ρ��4�������i���d�:#]\�U��2�!Ë����\���}U�X��%Z�(��^����_҄6���"�D���y��8��5��v*`���d@e4��7}�g#!��#�I!�����:R]ˏٽՁ&�a��UWaC(�J�f
ǧ,�EZ=c����޳�M=�H��Gh!W̚�1qǍ;p�OAz;�	3d��:�m"%ش��w�'9�Z,���.P �׎h�z5��4*f:�&�݌<�rd���@���ob�-���
܈v;����SN���&s�Ʒ�sk��i���Lh����L.��.��
��� �x�7�����[�`ի�WԳx�g#�Q�:X�$j ��(ެQ�\/p�Yh�F��30�l���7ĩ%��&`����1�d�4��|�!���N^��ﶜ��3���r�z�R�VnM��R=�ş��t�ef�`W�B6��v(/��A�LQ)�Y;2�	��� {�R���S�(�ohS�Eht%l*����P�E�-Ry���Mԫ�ge��@�7�/���Y��zM�F��ڥ˻H����<Xr��9h��L-�*g��X��^�bډ��ڛ�n���zC&��P�'��/w��+��yN�[t���X�Ś.B��X�]U)����8(p�VNP�uUC���ؗW4��V"�����4q�(3K2�g2g���%�F!�&*ʝ�>�fZ_D^��j.U��y5���C��W���t����Ԣ�JgpN��\Y��p������4��1�KZ�z��n򫠄q!��V��x�qј6��ޙYC���4�.k���"q6�L+l���w,Ώ*Ўm�8��@ks����{j��3%��n-�bv*V�V�2�:�5���N�9r-��E��B�TJJ�K���&Q}J�w��-�W�n&.�b�0�Sh7yj�3y��2��vꞽѭՙ�³]�-!�j��s�9��q�]��l��u�[ԛ	N�i��pٝ)V.n�ԫ(fn.��&_3��k3&�v��Etv�'f,���S5�W[j�t%žN�t鰝�X�5滧;%�ĩ4�S��� �v9aj�/{kz����eĎ�&�B�%�-S�Q�T���6�r���ʵVW�_�XUmwF�@:�6�8r��w��&r'��_V�獚�K;�9�.�+e�o�5�ۃt^�ai���P@lK�|�
N�+M��o*k�zx+�Z�E]ղ��˭:}��7)va�18b���[��x^X-�V�J��;�Vᯝ�P��ٍ�;�Bw�u"�ֆ��^a�r�������f��X��\VF7OR-����)Ӗj���B辄u��/�.+��O�k��y��nl#��O���J�a����PFQ�m��&2��i�3k:[��{����tOo�S�u��6�=��]��>)��!N�M1	�]���OJT��c��A�R����r8q�����V>������n�b�5n��2��T�5�
�Rɲ��䡷	�SX�[I�Hug\��"H��)[�`���³��44��!(D�Tg���p9��f�rsK����f��y�tS%���/M�6ݻ�[��9m*L]�f�"1^��F��v�k(JYJ�Xǀ���S�����c�}а�̝��m�aʀj73kk�����5,Z��7~��eW>��u��v��R�!�4sC&�Z�mD٬�.�����<���6��J_�zr�61�w�)>Zn�����g�*�Zu�-l���W�y;�B�kOr�-��;�-u=��D=���������N��q�z�;��`��)t�]���޻�+E��^Qm8���i6pA�3�i/r�cލ|b�ܗl(�mnT�خ�=��H��V�gk��V��Z�����$1fkġt�b̆�Վ˧�iC���+�pD%Z�� �l҇^���*������T�+n�n�k�N<+1�<�z�"֭�8h��̀�)ݚ�z��wuÔ��,:M�׭ڜ_j=ȘF����`���0;[��^��+;�8-]F��u.׭�y�4<�]�@�s;,�oS�u^�H� \��W(���xɶe�.;�gp�l�;q�0��M��G��M����anc��s�/U�oC��7����ǩ+��4�}ӴK{+x�nq�/m�Ŭ�S
t/h���cm�oj�C�/]/��UN�o]%N3�Yh��*� ��V����^<L�;j�]�Ƙ�T;Y%]_e��v�i2n\tv�gi��\����zB�݉����V��i�FsS��趙�^˻�*b�D̽��ӫ��f-��Y]M�7�/Za�Ĝr�(�Vq��sm#NM�Zˣ�4Ui��Sy��w5ί�y�8lj���㎎S���6��F*�CWs����u<�V�Lֲ�`q8
6i�b��#�".�[�fɂN���](u��Q!����Vm��/�o5��gJ���:���)�Vfʚm���:����uu��[F�|���i�wVu�]tO:�]=t���N�۳�$V�f,��ݚ��ak/V�Rh������O��@��j���+�k���,���P�3���G�S�=N�CE��J7yzj�s�J�ܤ�U��8.��yڣKD�1�As�9�����Z��
�EL�����܂��<���*�	N��3��B��Y�8S�Y�.ǯ0����\S�,�oH�vH�N�N�.i9�xc���g���t�ǎ<w���:�c�2��������:�e�/r� �f��	���5�t���+v����qd( V'�,Ē/)�unt"��4_H�<��쬺��n:�x-�={KY��ηFH!X��^��x^����+�n �q�.c�tl�W@E�	��f���k�������s���N����.�s�]����-����\IL���㛘����	�V*�^��\�T�%�."�)�_I�]jŴ&?��=�9"��U��Wuذ�RT�t�ۦj.t��^1ݶ]�[�:�M����:b�rv��L��e=���w1r�g
ˆ�W�Ν���ˡ�3Y����]���'X%3͛��S3`��/-����ż�)�s���*�pC5)�U&d�I��S�E@����i�+���ٵf��6/E�6fKSH	�
�����{�-&�:y�J��d:hN�1@�)}��a��C��t��4s��yx�J���1GvĪ'E�Kd]�'��0�8L�+{/*z�S����q:��Ǚ:���l��|H?^���,uˇM,:{��G.ŋ��[���e2Ou+3tj�e�߉L��y�{���̓;�]��l�<�p�7j9���ڭb�����1Յ����1��db�N{m��`ƻ�/���)����n�r{xj%4���@�Κ-EQZ�U�s���?Y��Q��xKὝZ
��v��Ʋ/���f�՜��i���˷�_]c��oj�wMd=��*=|&gs_.�%\��������Rn�pe>�h�����ޠM�U�#�b��kY����_Ǥ�XɯE���,P��ʙ���0�n�X����'}m�El?N����t�|�����d��o*�x�%��Z�o��zT
K�m��A�mZ��F�
E��"m��-"�N��-��
�9Y�Bۄb@N�j�V��ܺX�k�k�5/`��ғ4d��E�G�V'@),i�J�V�}6K��
�W�bu�Vތɤ�@pZ[;}mISW���]9�a~ɟl�p���G#op��]?��_d�oA:Ĩ��9ǩj��#i$���d�S�͍d�FZ�/nEY%4��yI��%��Vff#dt݁���˸*Z�"��4BLl������!$�(��e��C��+1ULuae6��|R)�̖�p�.��'���/����쒙f�R$J!�("r9D�LD�6�ڢ�eMIM�H�@!]�ZZ~�ҙ�a}�!F�դ3\4�oXՖf� -"��\�5aK4]B춑ŏB�T��@� ��:EeBG����R&��p�9J
	��`q"��Ț�նYB�	� ti֨�&��_H{$U��50�c0��'*ۖA�E<\GV<M5��l�&�b�%*��3U5���h������Xq�$�qQ���I�1.[xv���+���_'R*������z�]���'�I"�����������ϕ��ν=����ӝv�*�5c��*����vtu��Z����T��7uh�H�����Y�`-PŜi��Ɔ��ru���;��Ȧ�p����j
��[�$�p���p����b�j���x�����uor�=�-�4���VV^ؗNfN��td͓E��X5Z��6�]���g4�*����w�a��V�cϞIt�%oi92��}qebv@�Bn`�DG��y��=ab�Fe��e�n2�j6(��۩�r��:��X.�EV�|0�Ė����؝WK��rdVt'��md���b�o���+t2���#S6�!��v�򥝙���Ja%}�˳%5���Ȉ\�F�ñ�W7�*S���)��}�w�(��F�+b �}�f��vaʴk��gᏆ6ﭻ�-q���5e�A����3�Zr�r��f�/4Su�9�F�]m̏7���km:|E]V���a*���< ݾ��K�FrMn�DLR��N�7�
�4(������ش��ټ~x*L�ֱpV#8�Jw,�~�sFoh�(u\�͒~wah���C�@� �R�R��g�Rڄ�Ӹ�_L�P4�!�t���u\��:syaʺki��u�.G��*�����1&���ƗGe�w�'��"�t��٧1a�7W���i�Ђ��]Kwp0�9lI#�X���y�Rh9\oE����8����~?�|~?^�x��ׯ^�ޏ^�z��ׯ^��z��ׯ_�^��ׯ^�z�z��ǯ^�x��ׯ^�޽z�^=z������ׯ�z�}��O��ׯ��^�z��ׯ�^�z�����=z��ׯ_�G�^�z����ׯ�z��ׯ^�z�z���z��ׯ_�G�^��ׯ^�z��z��ׯ��^�z������=}�f�Fhz0YyW�i�.�
3�A�Yue4�3q��pW�,�d�-O�r��[C5�v�<%n٥���t3{`=�h���C���J���A$���h<�sq�sP���Z�}Ǩ��`�"S��������x��n�:��a��m�)"s�>�ζ^��)�ǝr��΄�4��]1i����V�0��O�]�N�w6���6�	��ɜ�,�}3O_a�e�ψ�������4�2�'�h��Z���j�z�mXq�ܬ�L=�{�z�٨���s������Q�rZ�Iy8�&4떭']D�u�i:�[#j�����0+��e�gj��o7ޒ�Pȭw���&y��v�L��=���*M����d��Q��[>�y�,�[���n=�z �#��㷐�V#�[�vu���,jB�[��v�D��x��,'Í̉<�2s����n��{�WTq���L�����_#&�"e��<��4��*c];�Wzp����7Xɱϕ^�%�zkm-�f^�; �,�7#є�+K.*�F�]p�mn��֪�9���������ǐ�e[��
T�f�t�_c1'1fCz툣K3�� Y��gMt!���t*���/A0d�Й<�����IR��R�y�sHD�v)��:�r��aJ�e��K���}���C_3�����}��ׯ^�z�z��ǯ�^�z�z�z����ׯ^=z��ׯ��Y�ׯ^�z���z��ׯ^�~=z�^�z����׮z��ׯ^��o�۟o��ׯ^��^�z��ׯ_�Y�ׯ^�z�z��ǯ^�x��ׯ^�ޏ^�z����ׯ^=z��ׯ��^�|z��ׯ_O^�z���ׯ�z������ׯ����}�v�`�Xs8����2���4d�����{y�*�zdp�.�"oh4�k�1d,|��,��rQ�vQ�E������mѧ�d��)L���e�x�
���^2f�x뎈ɔ훌$�Z�!��ʹ�z���A�B��VWD$�/l��c��(�jUet�MTg�n�T�ʞ�q9��w$�f������_e�>XjK�m��hj囝"	�Ю��۔L��u��u�7/lĭi���h�
�� �aQ$���MĪ��92��Al�[O��Y=���lp`�e.lS��{݇r���Lŭ3:��n�Z�Ž���p��6t�7����ZMTw��D���A�x�^�����z�몽�V�ǜ�P�+�i�s@'N�/H�x�m��(��/���u��_�>�_sd�Shk�<ȫ�f����}8i�ۚ+I��	����V2�b�o0�`��!7�#tFn�B�\��+�Fe�j��v�����b��I�R�ô�U*-�	e�1���!k-J�D�U�[vT��ۦ��X��j[�Հ�� i�zu<�΀-F�^�j�I�/]aɹ]��+mɃW�v����0n��#&����̧�z�JN<��ͣ�������Pܩv����g^��������2�[����z_3�4S,̮�=X{����a��r6_i��#��\[��m��Av���fnFR4�f�s�=��N���A��������EQ��-�����ue���$}��:��W���j�ƻD����:Yhr��i7�j&����uU؋ ��\��P�u/�op����5��ˊ:�T�|@vf�m_هkW4c1�z۩٩�	SI'���3Y�pݺ�m������t'*�<Ք�ԷGu<�V8������F2'�s��I^_|��'��l��7�:�D^9���Z�lvSʁ��i�$]�&Yΐ�}�#���]s;�����	Ψ
DK�Z�_3�mU��wa�, 7U�����4C�b��Cm��Fpɟ0�B�ɨ"Sz9%}yWq���F�ZkM��V�����1����M��+=J��Å�r����ˉ�M1L��e�&�Źp*�X�φ\��,�2]�v�t��c�^���� +�����}*�aŚ�1�1vCœ!P��[;-��H�]��ƀ8M���R�0���%��U�wV���
�34�9��(F�X]�jD"rXcM�ei�UX7���*1'kJl-+��6��^ԛ6�k���PA�o.�|��|��a��.�>�]�:�������i�gu�u9é$M�ӕEҝ6,D��uv@�볳�U����V���ɏI[l�%��6�1�g'���fP�nr�A�������\�Y��`k�s���K���(�;�c[[V�wg�P{��;A9t�.�K�Z��1�e}G��p��%���2�
Z�G�:릾0�_S=֤G��Iej+0+&\Q��[�!3z�ñI������n���y}��d��=�q��j��(�*%��.�N�l>�}�Jri��oM�b���tH��\�a�.�Ra�Oq	8�n,���/q�	�0'u�vˑ��ɚ�$*�G6�iVU����͠&a�y9S�扻x&.��J��/��ٛ���q���x�����P����J�v��bh�glo>��t�9�K�X[y˻h� �vC�.CY�]4�X�
�lsEǸ��{7�[���+���J`9�6q�9����/8����Y\�C��鶰bY(�N�Bܮ[��K�&g=BH���g_sCOr�De�pv,�ٴhɍ�5��W���ݡ�Sۣ�cbuw.f
=�sՎQ�U��q�ׂ@E�L���F��;�SF��*m2	���RN��Ff�%B�_�#}n�)�D y�>�H��w�v�9���c�Ks�U�dZ\L�xK�f]14���(P�l�l`Wb� Z��(��ՙ��e�]��l$9�%�G��o]�T�9ɶv/��s�P6Wu�r3�eeQ;ؕt�3���C�Aݛ�i��i�AV��qiJm�F���`�㩷}v�Ƀ	.8��5�YLRL+CQ�V��(�շ�6̭f�)�9	��E;�BIa��6r�@�7H춱�@�[N�4eX[�u-<Z'v��&.����%�b&�F�WAԃO$Tk�#�7y�R�uk�]�S�F�W(b�a���guK�y{G�|y�Ҙ��n=\�n'��%�������#n���vկ����^1MPLuKYp����OjK��m��M�/4Nիq�mazh�L�����`��e��m����ț}PGS��es��D{�8�un��;ir�,b�G���7\J�]�n���8~��:ֻ-o9@<��lY���V2�׌չ�T�}��W�mܭEg%38I�drT�*wՏ��rn�f]F8'�ctwx js8���c_Dqu��M��'
�=]�-F}��3t6�dpv�4��٫_�y�(R��f��J��Oy��f���#�����J}lډ⤦sz�H�/�D��b12�G��\|���l����Ϋ�F!����!	Zl����\!/~�"8Zx�X��*�fYQ�
	��fP?j�l��Z��YW����J�q�[̮�$'Ks(J8qQf�$b�6l�xv�ĵص�z�{è+�.�I+��<c��o�I��L�$���0֪YBk�������C��O��3o���F�ݨ�-5y������mX����Z�\q`@�ꞑ7��lpT��`�Z���]�Vm���K�'O;V񥡺�r��D�J���Y��h�F,�VΛ2��T�Ė&���:��#r�/�8+`�flrLr���̵3i������H위봎x%Q��z�;oI��X�ƓsR�����7Ie������A%E4*I\�o�lț&S���x�������{[+���n�+O
�"r�K����!�%���z�PI��6�c��ֳo�Ѿ�i&����u))im8`oIL�)�/T;�y{N��@�P����Om9�
v�b�F�q�2�N�ң��6=�m�j��b.��E�yn�gS��aj���3���I!n��r����{:!��ن��̖�����j��c'q��R-<6ո�ݾ�=Ï��	�"�E6d��_sO{':Maj�;1���@$��U�cN�U�{n���o���W3Xa��u�Pyso�r�z�j�ԡ�Q�?��0l�k�;�nޚ��=1�U��]G-�(L���ˣ��-UÐ5QU����qu/��VbƭMЙ5r��L2��0��*a!��4���q�׵(�nn��&v�[��2	}2�[t���]������zo�׆˷�)��3��U�3�5���Y���?2{k�3A�1�BNe�z�7/�A���rnm�� WSqP}����u�e��bc�6|r�`�Xj�.^��Nc���rN��!���'o���y@��@�v���|h���HT�A..������U�Ӗ�E���;(XW���Y�:�o؍�dM�.��� ���N�Au��|PQ`�%�0[1=�]� 7�Ա}�v"��n��L�e��ƾv��;.)q+U��a��Tz�u�|X�
��}�iu�lRi���Iʨȗw�S7VRܓ�[SG��n�<�*�bIה�W}{*K���E��lX�����7]J�f�o։3�$ot�v�}B;|�lL[�P!̠��=u�N/�D�3�7q���F�+�c�dtI;����d_r��s��Os:�&��sSe7�]���m�%�ԲA[��d��eL���HV���[���.v;@4���A��뮔h��p5�)Zo;�a�ot�\�99n�
��NB�Zѷ�v]�l�mE΅J�ڜGu3ݔ�[0�T��pm8XU9}TRW��_�;�	n����$=�5�G�2u�X蚸K�M�c��T�<����t�]�B�z2f�,D��hk-R6�u�}����;nq�ʳ
Д �%Ѕ�xue�{�/z��	����_J�þ�3�賂��Pd�ڑL��A��/�mb)�,g�׳L����i��QN=s�dɕ�<���5�3XU���3�˯G�l�!�>�,٢��%�з����Ȑ���Dn�����Z���P���KNbR�6�VR'�Bpk���J=��M� �@�$��0�����[����n�`��@�
��Aw�81w-Ψ�w�3fu'X8�/�&�L5b��ӵ���]K4��t�"�rO��k�.����[;hA��-*�y��+���\�S]�%��9�sU��xwjs"����̻UMʐ���f	6���9�$E��`�VVD�T0o�Š��9���JK_;/d��v�c:������2܉��mf;/�]�L3���������בWT��_S���G �.f��qѠ�R#���˓U(00�
�s�j�9�-;ᐥmU�/0�C�%�n��x!�JcuU`ܪV�
����h�KW[�-�M^�Yŭ'd;���s��el�{�*�ꑈ�εtK5�i�߉WӲ��]��j�	Bi�]�%Vˎ���ܜ$�U�=",�*Δe�E��#,顯��ۂ}��0_M�G�NU*�͝��n��{��J�+��.�ku$��H_8��x�(7?ī�D��z��ĝj�Z˸��WM�:/�R��m��1V�X���E�zr�=���F���鶕0�w;��::7���6-�� ˩�މP�ls�wӸ��ļ�����[�}�� qIXU[��7a�T��nKeة�Su j�F��p�:�<vu�r�T�K����TgN�d��1қ"�'���7kUo��J��%��]�v���+Q��λ�,N�ʓsr�Wvu�|�]�O�i]}�c�;�}�Z�l3c�c��O6�]yZ�X�#�ZrA�gS�1o��X�
,�q�H�»>�f�Hҥ�Eɰ<̖�
3sU\�v�yYcB:�����жÝ^�D�<�If>�T�`�e(,��
.��e?�B�j������nv7�AS��T;]�kO��PN(�f1S���"�Քm�׻G��EY��b�[���wK{h�=��Y��AN��`g\!��/!l�"m�����]�%A��r��Ѩ^3_$٫?sZ;A�L�WIKc��Σ�{���\��ׅK��Ě�=����-��,���z+�Qs&]��'�[V�=);Wj�`;F@`��T�R<�siW�:�P��P�C�H�J�uc�Ѫp�:�
�s�ַ�򔙗��ܫظ+�.t����������ܛ���*�s�Y�ԡ��;����hh���Ka� 7�r��xҥ�Wbۣ{F��.M�B�̳��W��y�j��<�w��;�����'����U*�}?o_���?��ݧ��������s���Ot���Y,��lY�1e���i�G됞�������n��v�b~�J��ff}ڋ���0g^��P�V/��I�3P)r�B�M�rMqSȑ�팸n���J��9�Ыc��@����eQ��
8�f�B��]���
�M��b����#��@M��3A���4P/��㰺�*:���p�s'�n�z�V3����Y-s :�;#eZ�����/�ud��a�$lJG������Bw)����ō�1m;��P|��W3�m�XVw�]oT�����u��{N���N�Y���uc\Ȭw&��ay��n�^��t�X4܁b+�&ԫQ+M^��,�v*#�	d������o�����̜:�6�)���|��^��47k*�bp;vy,��7�BR��L/6R��軣�?#��Ō3-���}�D*)�+��s{7$nt��Z����%�N`�[�T#�wa}$ ���6j�M��R�u ���@��+����X���f>�������@�4��"s�ԚcI��YY3��x��f]�"�}o�jۘ��ʗa[�.�'i:�˹�e�*�f��Э9x���O��>����Ь����;�%cJ���w�7�Χ��jU'�W�(�?�i0-�4���$�/X4��;\n���w�jK{,,�� q�Z(��m���	�Ղ{r`��ACA��[� H�4K$GT�Y�R(��n���K�ni�"����� R���*����f�l\�:4h4h�|�Clb�CA�#Irs�O�������~?o^����X��}��m�!�gAK�j�sY�m�ݱ��nZ9X��sX��֋c�s���������~?����~���m�T��TcllkUk)��Q��DHTƫ|�8e�+lgb���sUp��ƍ�'O�1�*�5m�FgN�F��Q[V�1zۑM%����涃ki֢��4nnp��=^y����ѵ��k�M�-b�F��kv�r�QZ�b��Umeӈ�Z��h�"���bӶ�DgU�i��մ���m��\�Ѧ�"-m[�^�1Ѩ�v���F-4��z���k��ض3�Å�9��ÃT�p���s��y���Tsr��TQO(��9F�Le�>#�=�7�a�z�/��rS�n\�69���KmM��9�\�1�+�p����j�(�F-F��FqR���k�Ü�XKj���Am[��V�ks��y�r776bZ��Z4X|��G����p�b�\���آm9�cr5ˁ��qu5�Er��w�~^����/Ke�}�X!�*�N���������V�9j��y5�5OO���[�,6��b�t
K�Mk�{z�f3x,	�)����B��лyW���?�lw���P������}��E��}'�i�_�׻�u��C(? ��Sj��X�y?x�̚�]��sN��{�cDtI%��r_{�ߍy�,�~��ϵ��.C�&��I%��Æ|,�L�T���iPon��ۙ�`-�Wq�G�p�m��$��{����=$K˩K���1�<�5K�f1��{ڸm�߃���ۓ7M��[6�'sc+=��＋>�a�&��xw�m�ȡm��;n�&���3O�y�$�"߷�S�v<������p7^�Ei�_�R��>����O��~�xWOVg��r�Nݓ����i�g�s�H[u�4�[M༻�;ݵ��ҧ�%�E?�Ɉ�"0ѧ��Ӕ8�TQ�����C���!�(�@���7��U�W=uw�Vx��j���7����Tu�1���w���)P|rs�4T��X���]sZb�U�1����i)���z�9�bN�ˬ�̫�sc�FҀf�]��[��F��K鸱WV��.�������$�@��q�ܫ�o���%v$qԬ��\!�w=k��� ��ȣ��G��ڷ��/�����;��{��;����n|���h�J�j��R��M�Wٰ�G>���d�e�;q�$P�#a��c�ޯ4���A�8=� 1�)�Ql�������k��ϓ���C
TOW�[��y�ȋ�u��Y���dH��Ue��ݚ�o:��#x0���;��|����������$e�:@7p׽��^��n�=����M���ե��)�_�;�d茈�״�g�����W.�m�����A�x^ͭpR�GݠD����p���������7dr��)�=GӢR�W�o'���y�w�ʭ��������M��c�à}lV��_���@�n8^�����~��7�&G4�;���θ�H�FQ�li�{*o����C��������ϓ3������k���M���U���G|lM���Sz��%��)g�m��#�{�����oU��h^�|xۖ�ˇ��Րp�i��Գ&HC�Y�af*��/W��c�fy���M؝�T�W=�X&��Hh�Ӎ�C}2�κ�ܗ��쳛S]��+�����P���n�Ix0n����t������SGWY?}]���#7��W��C^�3���'�uTN�(�>�Ǯ�˯,�|G/y����7��	��7e1�vfK6�ؗ�M��a�K��!}�WÆs#t�oXe�}�#�wd���;����#w��i�><���R�s��J����r|)��)�~=��re����u�rJ���O^UZs���/T.��@뿏�4�8{��7:��6�o�Z
�y ==�����=6�!��*��T롩�a����B��#�>�i�<�{Sw�6��b����/o�R��ߊset���yl/4@5��~�s�\��O��>�L<f������]Dh��h�y�2��,��r�����2�|9�� �P�b8[���P�����8��=��5�ݲ�����؛�j�*��W|,bǼ��"�g��M>5��z���eºp��"Cz*��ݴ�����U��.^s�o�y+�X2��m )ʆ?�+���������;��Qͥ	�s�˫�e���Z{����*�Z�v	m�����ur	�(��cȍ��v6�rú.��]�_Dŝ��͜�u>����6�"_��j��Ί2$6�1�|Z�2g�54$~�<���������}�IW�E��NO��]�@ib��G�W��|�MGI+�ߝ�b�pu�dk�hs���5�P�o\{n���˞��*v���%x/p|�y���)��{�{�:?��A�>�#D�ͫ��Jq8��������mp���k��|���c�����Z�W�3sKU�Z68|���g�v��D�,�Jl右��t�5�7ƭ���Ʒ�����x���q�|��훠��j������U��9���1�:�'4&�\zS�վnf��Ϧ���뫩I�]&6y�}�!��i����T.�/g�k�˓[������c^[H��x�<4�]�U��ϼ=�5|(�|+އ*Ӻ��?F�$�{}+����/���Ȼ�&�K�?UeS�Sa�X{�=8���^���Ȼ�Pw�K��.�Uwnb��:L�a� �\�>�g����� ��u���&f�0�MeuA�Y9
[*�:���G���BWa�l��u[��"z6o\'y9
��]'��4j*��El���F�%�Oɤ��H��w��.���S:8��Ȭ���{�fw���ӨT��=t�{/2;���v<�=���fP��"k�k=��U�0b	�inMZ#w�œ^RT�N����������O�	���q��ګ#T�}���.��E�Q�ή^��-�Qq�ic�U��{��5�����8���|l��XV��^s�b�x׻��z=���"��ժn���e
�G}�^���d�>n����f�&�����6�g�xE��`��ާ,et5�D߈���Ǥk�&���x��/=w�����3�׊���-g�P��Mp�z��z���#�}6	36k�9C���۬��B j�p���,g$�d6賓5S��R���%7�k���
B1s]C3�2�Ѐ���g99��Ul�^L3Rn��+��ط������:�ifz'[Sΰ�Z.�MT�VH�h�-�Ʃs�v�Nׯ>�<�X��P��Kǂ�7��<T�#cVd��i��E�u�R���0"b�-_���> ;�:7ۧ�37�v� XF8"�y��;|�&�<�zgV˽}�D�{OnW�gSp	��Ɋb�9gg�o��zI�y�ϲ�V�s�Me��c{�V�OfF~��zNݩ=0�:���>��*d�}w�L�<��z��z���[������]y���VW�������'�F�W��n��q�{F�I������ŷ���.<Z���hס��N�K9^�@��k�d���-KZ��|߳{7�@n�lm`�����}� h�>�oV\���`��#S��˹��+��v�z:=yo�\;���k��V]u����[�W��=����t�(�k�;5}�k����ۤ簇<�4���y�n{�D�y>~�}��M�T'��6��l���$ez��GH���6Z��PՕ�e���^����_��
k�qb�����&�"=���{K�w�� ��B���|���4�1������m���łi�v��,��d�W]�Cǈ��/eyxW����=��.��P},&�:�����9�Ep��6�G�mM�g��<tn6A��n���|�J*Ǣ*�D8}��#BM�u*�h1���m��Cv{vEM1�*���(�;��j~ر՛[��i.�9�C��P��#<���rd�����=�a�S��*������sp�^Ԕ�]}/X���wF��gxK�;����<5@-f�G��;���b�S��Rw�c=O+e<}�&g����[3��e��>�=၂�N�����u��S+�b/gѣ+6_�Wy��:A��w�E��r/���?U���V��u�Ey�=�ծ��m�}7��N��)�}�eū͝=�Ɏ]9/4�4���g�.�_�5t�
�/uc,�ow�^,�.�D�}I��}�c���&��|s�m��S�)�Ng��]�C�4+wr�W�H9��P�����8O���e3Wv|��Nį{��W�tBj*���tG��z����~�s���BjJhɌ�]�j�y�z�W��P�m�78���a3�KY'^���'�(o����kG&Ȭ���ΰ벮��̝I�
�e�@�����`�,�y��U�2kLvn��f�0m�+��-c:�X2��&�+����jvu�	�Ǹ�^p��zm�XU��c�o���R���D�ISjm�?o.�y��/�W����BU�e��s�d��|FS����dIok�NJ��U�_D${Yt��^X��pU}����ŏa���>��D�N�ks{=�V���W��i~�D,Vy�����q�*��}��tu+�#�r�����K��8�Z����{|�-���^솟��}͹�d��n��W�m��t�ӿ4z����;�ՙ�^��g䈧e�G+L�G�L����)���[�y��z����w���{c�����}�j$�<�I�B��q!���m��5���}e�z6��Oyg�|�F���z+P�C��2�>��Oo�0}WU�ʰ��ü��5��^��Y]�e����������d{o�+g�M
%ߛp��b���=}���7ꉄj�,�PCW\+�y��۱�vcO�h� �<�M�9���y.kE�+k(l�d����5���(�b9}+e����&�%+�3�n˲qb�\x���wya�
',p�@F�q�Z���Շה�̬x�2��rWowi��I�q���Z�OH7�_"/i	3�Ǝ	#�W��r��̦�K쎜�1Pڴ+#$���Cͽ�s�"g�-���S�����>{"���;�����cC���u��ؽ�h9�['���s4�eM(���R��&>�/�C���2���:��q��j{��IΣ�O6f)ƻ�j�~��\�ە��\���<��`�XC{6�$�Y�7���g��J�rB�zJn�h}�`z��3Z6#O��v�̀ߙ�s`df���2���y�=�%���΂�9��U�62�y�|�j�\U���hӳ�Y3��W����z�J��ю� ���o"�b�q�N�Oyxte��b��K�p�V����f@��"v�t�dO����3��}���uN�^Fl�J.�周2�	�"!��}2�r��=����g����n���UY��i���>eѝ��;��:X�H=��g�l�ɍ��ox� ߏ�<�����]c/x�^ּY�+��)t��^�N��[2:<��ø�;2f<2�m!\��>�j���D�kG1�R�;�]�;�����|����y�̅�ȗH��k \.cdt��ǘ�}��O"z���Su�:����<����12wY)s�+�U��F���(�u.OU4���mk5^>��"��z��r	���y�lԚ}��>�+�M��;���U�ؒ,��:\�j�đ#��V���3]F� �͸p�����?z�7==Tm�oty.��]���f�S�w!�H�#�=ȁ���]=U9��{_����f���f�CG��E�z�F��wd�[��8�>�!�=x�g�5��9�'��,Ei��[��m�y�7`��U����9�"4�9I۲zf�������}�ھQ��{b�O�r�Yi��7��S���g�|��ٱ�k��r;��q��\X���I�꧞���@��`o�k@h +����3+���b}����؏H��<���ٛ��|_��G����W3�N���}B�-Q�k��J��Y�i�:}�6�3�h���������~���!�������s��=o/~X��	�܂�uB���캑g���&���y[���Rr�h�r���*�i�D�9j�؍)I ��':&���0�
��v�Y�N�*Z��6��&6r���̬�C���tW����;in"���s��u����x�35�,�tZ��̬��Y-ů1�����k��.u���[�i&'i=��8�J5�jZ�!{�S&��}������;;�i�3�v�ӎ:��ȫsj�(�.s��m��#6�d�:(vOr�ɠ�صe�z5��e���DY����Nb��Ǔ(r68�Fu�9����=6�K7C[�/�)�$t77GeIfgf�/p�ń-63s�M>��Uz�����[:�*����Ҥ9Kݩ�٦I��D��k��=�o~3������Ƿ��R��1	G���9["}�1rگ��E�� �r�qub^��T�ոi��8��5Æ����jͤFv>�q4��\7��^��C���~���]KQ��N2)�a)s5�F��2�8��ϯkJx*�b��Ή�n�#��kqX=u9	�6�����3��ޒ��/��1G�R~�9��w:�{Ka�e��H��s��:���^�O1��Ȝ�m�.�s����k��5���5BXEI��e�ΞC-B	�&�92��Yb�(�rZ�gU٩зFK�#s����n�[<�CjF	WӞ�a[u���wbӪ7|�;#��hfe��=�
8�!s�SI�q-}Z�:Go]����uc��s�W��՟Nmzw�0�x`��h���	�2���A#�4N������DtY��C��}�	e��8xqГ�ԥe#�N�:��c����)��΋�Z�\~�{p�`�����zt���ތ�C��tj˝:&D�l�r�ak��/4i�1���!g4�r�n�k��g�E�e��;/D�3-�ib+b�3�U[R��q��)�[ʳdJ�OI�����rTG5[�U��3j ^m�u��hq��5��4^�9fr���x
��ݤ�nĈ��DG���ar��z�8N�2�f�-6��V@��ڂ��M\ך�e���]�S�g1k�F�:�PΩ�Xw�C��Έo@;a���u��C�]J��9�^9�}F� -<���c��N�={D�Iy7:�X��af�\�;{7"�v�bhum,K �� �u7�"���O�e�ݹ���M�:Bo.ܥYx�Ril�Ŏ�d��,&rH�$U0�sD�ѝJ��Kl)sV4�n��F����xPR����(S\��E*��)�kТhl���k�$^ />�O]�Z���������5����Q���po�	�ҫH�RF76���)��jhގ�r�f�r��(���.u���_K�|Ɲy@�ྶ��/+����sv��7���U��Lge�w$��4�fJ�����y�~��������ͣ&9k�nb核1f��9q�d�[��T9�ٍ����nm��V��[�8���79�g��y������������~?�������߽�cA����m�2h�m;\��2\���m�5��s�h�� �9nns�ƞ���<?�o�����~?�����=�v��G�sq�sr��9��j�Ʃ�W���r5��͵�njLt[�nnZ6ۜ�5�s�W9p�kU�m�k��LZKT֮s�q��lns��5��v��fւ��9G+lm��6"uQEm���ccQF��؍��*i�crל��E�9ͳ��gF�+͙��QSm5mh3�cF�W��9���F�EZ�m�H��������4TSL[j1�����5�ͩ�����5��y�rrE��7�����8k`����3���-��(�h�F�[b�ъ��-�lj��f�m�Qlӵ�ެ\؃���9�\��mm���5�;f�q��sVu�i'Z�
*m����v��Eh�u1V���*\o7�1���d�Z��Z�5�ѶX���ѩ�3���V_"���`eAj�ZF��"���t������V�x�2l	��}���UZ�}Ie�=���Y���1�˛�I��}~o7�<*7[��s��5D]?�^Ӂ��u��ͬa;�H�E�Dx �S���1��:"��l,�+��2�O�r��N�������P�Ƙ{b�
Qx�Y�oP���,ӽ�[è%�d9Aw��i�a�B�\%�]Fhk��{���B�Y�>�5x a4�F7���������[J䩛l쀃'3�fg(�EP�f��]���������e'�ğ7����n�a^�+�`��دN�l']e�W�����y�Oe�|>7�;wD۩=:������o����~�k{4*##c��`�BQ��-��u�viOGS?!�������%�p,��B��՞�e~PR�A�2��"q'^���h�0�H��0�p�����z~�.��D�65H�7��2��#ny��.W�G�Hf�@4:	γ�j�gs�H���B-K6И!�E��>���4�߰�NV1�J��7�5 LY}�%[j�&g�;s�oj+��.�xM����a����9���ê���c�A��b��A.�z�ð��P5�oe[?O=��M7����0�o!��i�9�aᖽ;�M�3�ɵ��"�@.�`�k#2��|�ٕ1����UoOT���x(u-��+B�ׯi��/�'���8�Ą�����k*�s�#mʺ�Yf1y�A��o���Kd6�̹3�����m{��u�|ԭWݱˮ��v�vMd����g�n���n��o7�M�7���s�j�@�$����:LK��� C`t���'��g�>W� N�^֙a�͚��hԇ�z9�5�����_�����A_Ho�/y �����D�x�eG5׶��6�M���9�2vg~^�4/�?Ia�^5�{�˦�����W<�����G��AZ�ZGE��d��������z���ޑ�gRN�F@�H��D�sP/���-~/��6q8u՚�Ẩ��С���Bi�L,s጗{v�y�3�Ȝ��v�q�`H����@ƏU:�6Fs���U�it��>/�m�08�'P���ަX��YF��5��I�o.�l�3m�]�1}�A��C�^ZC ��˴��|�����D�����$��xC[����@���X�ms�y���:e';��QC��d8Atpd�� ������3gW����zw�a�Xd�$�>c�-/$M��et7U]�Fo=�#���=�{zO�`� ��k��_���W���:��o�y�]���ꓴ�F�ܩb�CU�'�y��x}�W!_����x�Ƀ�;��yE'V�P�r���5+�h;���m�8�"�������T������d�Ő1�}E�huX�IZ�^Uq���eL���2��:=�Y�W.~{\���0���8���ǣ%	}9�����4��^*�&(X�۩S��*�%����a5ՓM�nq�'���}��:����H��i��+�
_�c��vr�݋8߭��>g
����zz�X���Y�H������L��xNy%B����ne�yv�Mjݏ_E�����|a4��WN7��9A���u����nt� wR���L@X�&�P���cu����w�#�^����O/ry�؄���sȾ�,�� ��Wl[>�ZҎ3���<��m�:�n\H����zk�%��yD�??��ׁ�U��s�A��H�7-���q06�ΰ��:��Z�\�T����P�	��»�Aö_����~2�ˡ`����t��a��K�~�Ol9���d�,)k���~��/+���h&5
�//���%u��n?lWJ�������6KR�hLl��p�b��N���`�%픿0ն$>��^��H�S0k:zi����{^�4?���(-��P����2پ�a�C9*�6��>�2�]�L���.&�.mf{�o��c�C!�/LY.���������p����}9�%��>��5'[�͝��[�#Ys\�����X皧���;_�̟b���h������T]�A�E{Dap$C�|a^Ql�J�]�2VV"���T?=ǥ&*R��V髐3��*�f}.s�95.�x��T׏voKЍC�̂=���1u��ҳ5zc��c�����a�Bv�wZwkZ�G/�}ڰu7L�C/�l YLj��"��/$f����q�;=�������U�r	#ݎ�'���wO�!�p�o�醓�-����:����!\6� ��i�<������5���lF���
-C�/^K'�
�y�F��`��
����l�Գ�"�k�n�ݫP��1`�=�sI��Q��R�eT�5�!s�>��Y�)�m)<��zq�q,�Ѳ���6�$��ޡʸ�[�z@�鱰C�vϞ��Xک`9���M�`&G�
OH2f#�b�W��v�׉�J�y>���zǫxjkgb���K�L��W�k���A�'���ofU�u�����s�{IO0L�����P��z���/��[PN���!�	�_�.��nE��ȡܞ���83�{2y��/�:�Ǌ4�����a�&��� �6H�0\�v�+\���l~v({i�7V�s��_@]0�ʥy~���lGO�{��$A�Ң��<e�}��nt^թ�=݀ne!0S���УfS��eWC׭@��ʂƂ�0�ԜK��x�iryQ96k1��.��0�t0t��F�
���p[	�J�ޖB�w �n��|�/3����~\��+���"�����kJ<8�U�S�iu���YA�vC؃�t�T�٧��SA�ͱb`��X�z��7d<�b��V�v�;aY�����[B�EYS�>ozB�*������h���>����դG���ÚM��q�ql�8��ـ����Aíp:�1-�6KS-�>-�(Ӿ]��+M��S9���q�ؓG����T_��|`�N�`�� ����;k�v�m�՝6�s(����a��G���5�^�@�[�Lq�ۄ���}9�W����C��>��k��:����+��T��[�g~@u�ff�y?���	;(��I� [��s�]�,&��&�+��
�ވ����R!�_�:����w������ma���x +�<;���K�J5�Zv�9��T���ԟ�{�uu��kgT�!�??����]N�_���ei�^���J��Iw)��R��m�[���m��y���p%��M-((L����uuS�Od�⩛o�v�c��Tw2�X�k��������3����r��U���AI?�!e���-}/�ο7�_�E���7mb��Vڙ:h�H�oր[<5��Ԟ�+�[<���V�Ts~��&���=����9@�S�ѹi�ő���&-!��C�N�Cy0�Q,��J��`�i5����q�gO^��B��j��2�{1�!�!˸o3�Y܂��<j	Pk�y�y�?y?e��I�^��\���t[S��U��������P%���d��,�J���q�^%��}�DЎtS�݀/+��ټ�D.�GS�rl���ӹgem�϶�p).ׯ֝K3e��y����N�I;�Cţ�����/��/��<'I��"S��S&�����s�O�p�˔j��y�̛YU=�<��[:0���7�]�#��0�w��O��Sy1X�"�U�9��mTH]&U�͑��u�S���ѱ���F0� �C��nm�=�`� ^�5��K�]7C�zO�.�f�4<�WN63N�!Q\����p����&i����!�[xa>S�Gi�4���ȾzLx�1�0�ֺ�Zgm����2Al�����nC��G�1���5�w����Oy���w}�q�;����`q��:�T�oc.�ڱ[a�z{y�1Q{V�� �]��ɷ�Q�
�|2��H���(x.!����y��֔���U�m�:P�3C����T0ۙ ��;�Y���UC��P������!ۤ\0`,��B�v�U孹�C�YСŧ�鰽K���z�F�u$��df�D��LW1n�VY�z�g�xѕs�y]T�!�o6qL�����v�
9��F�3�{���`s7�n�m};'ń�f��q�b֑�U�qP($��J��p�w��� }_�ug!/4g�L���ߙ��u�b�)͍����7�~�@���ĳ\[�.�!lg�>�H���0P��U�6�����������K��C�+��6�Goni���0�VEFWY�TMs#�Zk(�7�=�bG]r�\kf�,RD�r�s�Wǯk$l�]��f́����Z����z�<ʴFYDi@�xu�oDn�}�/q@�_>S�g�����֛���@?`�)'�}�$�qmF,]������ou��'��c��4�$1(y��F2b�8�r�y,�j	�z͜eY��ɤzw�o�h��PF5)F�eK�y��G���/L���V˜��ln��A:��B]Z�9~����/m��8����lY�}zĸ����p@]:ɫ&=tB��r�):���(RXKjܐ1����zgu9��#��a���5�$F��(2.��'j͐�^�	���$�0ˉ�� V��U�7�Q�.�nVn�{�=���)FN0�;"��-�bc����%��>�9�U�����w��R�VSt�Ef���W�(����AF�T�0H�+��k��nF4Ð��` G<���!'kLjf����.��1�Y9�6�E�.���#h��<ע9���cPA¿tC�N�Y����a����2����?�����L�3��?��W�âZ�Œ���Ƒچ���#�3�TAd�oNj�~B�#M�R�~�3s�xz�;q�K�y��ʏ���N8�T�Z��3*u���O�\���DWw5В�*�������Y��}hTS#R�;K_H��b�gJ�sQw9Y���kR͛{�ZJ�iV�2㡕��Z�*�`Tԡ�¯[���7(һ��ʌ�Ejd��O��JIה�E`��M}��[�u� 廱�&�ȹ�/7�� *�k�T�b,7�X�`鵜'�P�Z��еnd㎿1��ђ����Q�/��j/T�Y�-dƉ�C�R"�c�w3�½B�j���9���:��XcW�����߂~����N�5V�L�cl�0k]w;4jj[�����V
?zy�����'��!���4O���n�v�磤x��G��*���U~��xư@�7�AN���	��CW�ƺ�@�(�����<�j~XE����=N�4���݉���ܛ�/e�Ҹ���`1N$��i��ʽ�6�ƶ3����~9�E�q��*B�v ���nf�kߦ���v5�^A!�vA�%��gͷn��L\:�=�Y��^�ȭ�W��{���B#XG\�DX4\�ƞܪ�ƣ�]�9�A����V���/�.x=�TY=���3?{a�mLÝyg��scN	���q���1�����tiM��Be-s��1�7�D��?E����_���w�7VI������q%�B{+�4��O4^�ל�	ndLD'�̶�D�r�"%��%�PX& EP��d�=}Ǆ���[G��!���уo��A�SM4?T�c
ڻ�]��q'���ހ򀝣sL�Ϟ3N���ʏU�\i�d�7���⣙��ݗ盖['ѥ}*ߖ� �mݘ-��R��r��^�dj̭�/{�S/��e'U��k���|�K���雦�Ηz�^�����ޭ��M��*{�8#�.��S�/ K"���I�߮��ι
Wq�U�K���9oP���$m������H�ha��]�D�u{��>s�t�G*�]`n�cKz���s/P���c��j�,�yx�Y��h��nh���Є&50t��/��H;��S�����"����a���\�AS
妱�������������(�s>a�`鵜��~����d�`��#�.�Te�֣������R���z��EI�fC�K�6��x�ׁ�޸oo��1�o�׹�����l��D&���nJ_n��Ӗ��f+��u�μ�&.�Uϧ��ܱ�TB�	�>��j�h�f�z��]�vٰ%bU1�}�C����d�A�u>X�>�z&9��f4b�>y�8f�H0�E��^3u������.��j��u�vO�3$3e���c�\�}���_{B��a���$��f�[3�W �f:����=����ݸ��&����/x�߻�7Hͬa��$8�}�d0n�}��������*:ǩv:gO��]y�j��z9�FK�x��^t1�l>2OB^��ov�����f��X	e7]݅�?/ֽ|�e�$Ԡs �2GX��JLX��q�q��m����c�wlW8WW15�7�iG��tfj����p4�ۺ�L�kO&�(��;yX�k+Y�wL:RŪ�s�z7�)��j�B���4�) �z��7yL�C���9��׿o[��Y�rg9_�;�����{/�~{U$�_�yKLϵB�aq��
tlm>X��Iz��i��m��9N�ܭ獣�8�(�߫�*�y�R܈���s?,2���o�B�c�ax�Q��w�0�����xY�CDjŰ�wC2�1�8#\eR�)��(ΰ�;�1�ޭ�[�y'�"XY�P绐�;kD�w=�*�+6G
��殈!8�Q,��)W��_����]�#q���ΞE=�Ⲩ�>�}�v�����!Z������_e��z�)�|1�ީʁF�[\m�6�O&�vu�(D:��Ó��J<���z�)�	K7TƆ2/��)�]č�4��yР��(�p)�D%��P�7���Ї�_�%���_��� ���A�N�g׳�E�v���H�z]���P�����U���1	��~b\�<A�����[7��`�ZC^�3�U	�(�̰�P?�O+�
!�/o-���j��C՘�zu#$��<��0~�|{��.��惶y�QЦg%������|x٦��%?o�5�y�*�b��z��ͺ��� i��}U�U�S��I�v���[�ft]�	��X7����T�F��k���ٌAiK7����e��[�K!rl:�i�\��E�x�or*�ڡ�۶(����Fֽ�u��������:+T�P=����6Y=��*�v��b������-��Lڅd:�`��f`�6��5k�54��w;��87;q�Fl�(��Rv�p��f��F�#+z̑t��k&;����*C#P{e��fY��d�W��a@��8z�@,+�ņ��@R��O��p`�E}�4C����:��wJ+9P�zu���R&��r�����J��8=�H���AVɮ�;�KZ�:�-�7xϠ%.��r�$�[N�%eR��E��/����˽��jH	�un�TQ�G.s�fG&�R�#�-�v�K��([��:�41$>����V�S&�N��î�:�1;ʺ�N�8vr{)�hV�x�͂XX�zZۘa����n���8� �b�q��l��8�9r'}���w����ܩ��M
7�b���^Ɩ�H���h�Ku� ���aX�Ȏ]�2Z[�^�}�{'Ay�)�6�Z�*�y.�E�۶Fm;�/d��\8Z���zU�:Rv�,ԯ���ԟR��N�U�c�"`�R�37��-Q�')T=�*�6b��p����A6�],���<��\
�]�wu{M�Ц�2��S�E�傭=�$0b9��gL�߶��aB�2��s�G;�D=�h���ؖiB]d]��NjR��61��2!K�tl�!�2�t/�vkT��y���v�U�//�����Nt�@D�8���lwV�j�����De��Y�����o,4^R�1+��>.jU���l���)R� ��J��T�,YM�"�p�;�����Xj�r���u�.q���)
�9Ev��YӔ�8wq���^�ŀ�Wbˏ�3�2�����W��X&��%F�0Gm�Hs�0h]�� �ҙ"׃�Ѡ�@�<؄�cW��I�����/\�lܨ�m�DiC�]�P��z���:�	n��A1툮N\�^�[���s�K��ͳ�G��?J��3d�5����u��7*��z0��}�5�4����84���sw(���pW��d]Mк��2�Hvt��\V^)G-���	�pAd�O���P���ѡ��Bh][��P���&��6���tި�''�����u����@\�I��L��C)����S�P��]+�r���K��O���5J�8��YӨ�2�Y�؎���ٗWiu�Oh��E�Ǵ�VR:]`w�����i륔Wl�dG*n=nK�ϣ�(vϬۋ����>}J�	[X������廽]}�#CM	G6�=��+X�W���zw�t�.1��>R�g��'u9��0��Z�\	�|�&�|w��,����N������
�xa-���N���T.�
b��w n�)'i�	�N���R4D����:��G�=�y�|��p�?�>KU�����Z���L�*�"��Sƫ�8p�N�kQ&g<~�_������~�_�����?N�'F�U��Z�EJq5�h5L[cF�;̜�kh
b�f1m���*�sǯ^�~?�������~������*��>X涎�\6�1D�3�:7#�I�(�bh$��1QDIU�6����CkZ�UDLUUU�m��c�lh�����'guz�Us�rb��Q[`��Ew�mMMc��"*�]�F�ΌT�֨����ٙ�ъ����+8�6�љ��:#�SMDU�6)��j���"$��Xu5Sl�+d�l"�g��<���X*��Έ�$��mj*�5�{MEyh<�6)�M[��5Q\�<��m�kF�O7h�����k��j#�Lm��b�mZX労��ZqVh*�mU��EUU�8�Vđ������4h*�(�$�l@�� ���7"헚�7��I4WH�W�v3#4���i�F�e�wX��癄��&������l΄����Zbfv�)�ρ�t������T>^p=��?� ejw�E����Зn|����a��e�|�}]f��|_l/�A�ݕ�Z=��nW��� �(^=�kL8����>M�Y��% �~�DP�Hc��S���yԸ�~�����?PkN�	ؙO��E�������s�Y]n�my��Bk��vyj<����"�ڨ��c�ϼ�������4E��y��@l'� ��o�k���vr��nϲ�Z҅��HF��n�Mބ&�N�d�q�5߽����\����)&0y�� 0�J�w73�.˞n���7_l�G�{`���Ź,��3���8ʆGy��Т�{w�(�t���y�<s��TE	,3׮��e�!?ˎ�hk� KK�Y��c�Pʋ�1��Ȱ���v��� ̽!@��3�bS���>��O<��2׿r�N�j�JĪ,)�x2�oa�抎��8��.[�>H�oQa
F`�I��CW���=�)��tBd��b%9x�a�=�qy�A9��ٳ;��!*��[�l0ȶ�э�cH�H ���g�Лntdٱ
�~Q/X�����^E��g/�g�$�F:�k T;B��c�5b=�����۵Km9MЉ�]Z��U��;��Wt�Г.oN�d�{�2��],�.K77;N�m_tu҂��r��r��ȵd�un�H��/��א��gm֭������� <�8 {�f�i0a�m�*k�'�̕�H����.b��]<0����0�'��a ��MK�TL��9z�Ǌ|;.��j>r�3�>�5�'��6Ⱥ�09�������ߙ����h8Z�h��.P;���fg:�\ԓB��&B̮xj�r�͂��X�K� a��� �~e�#6���OlUR����M�DǞ5�	�B͹���l�J�aV���*u���O���؉�5zKDe��i�b���}mj��s?��L�Ll��B̀�N8�z?��j�׍yp�Ա?U<�����5~�tO��]�3HB��@���k�a�d��a�Y�P2*�r�d�T�N�*��mr�tT3N�&����1�^ϕ���\,y��?�? ��G& fZꈧ��Ƙ��AY���n���o�KLIr]����L˴��c]��ϵ��ϴFK^�d��dӄ����l����z-�S��ܖ`�y�h���� Ș�8�pok��>g4^�q�[�������^8�̒����۱�7�Hyn� �W �="<΀���꩞��ei�L�6Ch~���]��j-Lۣ$����]��G�e�h����%�k��'���mk�\xh�ԼYەa�(@�c<�L�}�뜵��V�i'ѩ�i��]�R�kw��AN�)M��vk|�cw.�|���e1�������F�Qs�"z������Z�#��m�C��9N''2��MF�vL�[.P�;W�XS�(�r��M�O�u��=�1î^��𬘸w��,��#�F	��!�zz+�tk%cj��s�	���V�5=*�6���Gd��ۑ^�麦*(���Ŏvg������n}��+��j2��KɆ��L�[�Y�>7"�)���`��"�]���z��	z/]��c�����Ou<ae�7;��b9�C�B��ӽ2S��x�E��<Q�������n�N�@թ�^�����v)��P��^�/�|�C$H�^�a�_E0�~�E����z���r�9Ux���f-���מ\�;ۼ����AX��-��D�2���)�u�Qg�`U��g�7w���U����՚���q.�z���yG�:mi���&$��'��-�܊%OK�0˥<�Dm�W7���
�	9��^�?c��aß�k�����d�2�綗Q4t`Q�ڳysn�k�J	{���9�������]�~(#	�<y"u~;���/5�U�x�.�ھ�g��5j*P��Et3�miZ�w�m�'h���eew��>�� ���bNٷx�y[nU��͍Y
-�u���:s�6��Zt��n��V�U�Yp5��M=Y�ݔ�\��r��z�fQ����o�����@�r(���_�~��_��}G������u�8�ca�u>_�)���1� ��1����}�����}���e��b�1�t%ؾ�d�l�{)?Xc���D��zA�ź=B!�Hݶl�|_��_w�S�|���6�V,�0�����Ҿ�ٳ�!�z	D�@"�cъL�.'3��1UجS���}��g�!c��!��,��[�Xݡ�>�Φi�;%0+0�vÛ��Ӌ#���,��@~��~H){/�r����LX�ii(M"22��ǣ��[f�#��7�qTn�t�voAf��x2���X��,����r���?��RO`�X_��<N�D�N�B��|��7�q��'��;�Jl��Pd�Jx[��ј��O�ѫ]�3�S�N-⋂�T-ǖ�[��t�P�P�Dy���wl��Klt���'�T�jSL�J4�Ϙ&;_Z�Ƕt�n�#��·���������.1xlIv`2�9��� ��y۞����d��H�T
4��0�>D�P��f��5�-��Oqp���i�,�@Lpc}�
�.��I��"��u�Zq�K7d�3E��3��(i�H:ܝj�ݘ^bU0Z5��%�ʗ��з�6a��X�>�\��.� �Y�]+.��(�n�ӄ�kQ�׽�7�.I����[�X�*f���_U�BPq1��b�����u޴jN�ѱf̾H�[Ư�f����i���!%��2?��9A3�
�s�}���������s���#ZØ����}M��! �� B��86���Q{�.�E��	��p��L��Qi�Al_:X�A/K������a>=�m�4�>`T�P�@���^����[��CL
���Y�-��خF����/-H�0�Tw='�q��/.�ό�����9(��w���˙��o�ӥ���̉/K��)���������،y*�ʦXطvm�`�Z�x>S�W97]�_z)N�#Ƀ�y�d랽.��>���0Xw1���tzq�Ix�V��{��u9iMwq;���䪧��	��C��΃�M�[Իw��6�vP���I����0$8��ب�����c���s`�����A�e=�z�~^:��/�#+��F�[�Y��R�_,���t��v@�� ��q�:"���x5�%��4\sH0���ŶS�Y��r����t�p�k;�C3m�_fH���vA)����˶6�'-���e�,��d;������uUs���ݬb��'4
99��%�����g���U����}�����W3+߻1�(���(�m��>��wp�*.��+>��|��$�W��,Y��t�Ɣ���N=��淄Y�;�EY���F��6���%C��wht.�˝���L183OM27���}жc�dUj#���q��F�+6�#���CTRt�kR��������q�<�� xxx>�quV��!t��!�3�l.�$%`NE[W���t�q�.�g���f�	ݑ�-���c *��fo0Nޑ���LIv�ӬZ�L.z�-~O)�Z�RmflÍW����&��Z�]z���]ŲQp��3��	�A�p�<y�^�7	�t���t�?=3e�k�����}6�s��6��][��*i8���a=�m
�}Pށ �4�t��k���V�x���:�γe��|}E���P�Ss�ȼ��)�Ɓ�l�|��a[�!#ZD8'����h�Uu�)-�}�΀��-�7:���
�Eh�8�>��敼�4�O>��?<�lg���Vwf?�gsoSIܢ3�)�!<��E�^S�q�8p�a4�Ts�Z�@�*Kva�gw���v�K��~ep���yt����t��&���ΪNг`9��.�%QaB��s�R�ap��?Q�q��{si�h�{e�n�`�6��v�� (t��4*�Ni�jÙ8��X�'��i&�άݓc3W[�/��>�4�+	t�@p�|g�>'5�e��XkB�k�q���4�VՋ��vڔqt��+�0ݛ��f�ͯ%k�xs��B��h�7������4��mss���uv�W�������u�顎	 �ҷ�u�zx�h̸�T��[n�sˁ?�mYS�s˗b���.���J��,9ݪ�J�2���|>��9ª'�}��]��s�����>��k�C4�R��z-A�����r3X4�����[_l�gRk��f����������A�)0�1%�f�rb��g��b���Q&?b\>^��;D�iX[��pXS����<����3з�@aZ^��$���O�3t=2�tM�˚��!GW-��&/[k�PfR6�I��F���E[�n�kH��C�S��\��W#^m�Q�E]��::b�ܿ����E<��,/~B�+�ħ���쪖Ơ�H\�ve\����c�,��;a���p�oN0�.b��lS<!
��Ղ���~z���کnh�M��&�ӓ�5Wf�2�r1K
� 8�j�&Ǻn�2�6)YE|���f�	� $2�9��+m��Ŝ��w�Yz�I���s�I`��B�FNc־��z��x����EL:��.�@�(���C^�8�\g���qT����d]`n�c@�I�;��y�)�M���,h��W=������BE�6Ϣ^��%vI������U]!>�ii,.X�K;;�/�ׂBZ(�']2ve��m�owoE����M$�壂;��H��܈^�B�Muڹ.�K�}��8�Km�݋Z��f`�6y�;g�lG=9ɴ�Wȃ�
6Y'Y�BfM�.�,�d�$=ͧpNI�6�Z�'v��˔)��翼������83�(���~w��
�^<�0lp>w�@�65�"���n��B�N�xYU��j-?6𾁐Ϙ��]�Y��}.Q͒y�~�3�]`�6��������y~���x�k�'(_*��拇�"��=-�ٞ�6�T�#y�ߩP�z sIzp�; 8�#Xw���\\�%����7cf^��'|��B����ƶ/�6�{�Jײ���uS��{2��u�H��@A\1��y,�զݹ��-}:Zٚ�ºS`7\r��s�N�m���[�J9���1/A�v8:5�`�,��]�����Yy�<����N��|7$3d��R~�1�'�nD�^}�D[�����I&ꧫd'n@TK�pr��qq*l���:W�A����~��xne˧ž��{��5���v�v@�O�EC��!4��2o���=	zǬ��CZ}��L�5�\:au�s��buK	CNP#�����}�ZgK*����}��8��/X��O<.'�1���q��άe�9�ͷ�$1oR���$v��ŧ��x\:E;�amVg����Ŏ;�Y;�/}��NC���*�S�E^h��{�z>�͊%�h�7Ja<rg�t]�Ғ��T|E�}L�����Y���?.��)��Xuo}��5cw�n�,r�ڜ�B3�7�����4y��Jاe_j�sM'ER��Q����tnrxb߼�V�z�p���9¨�����r�DG�p;���~=I�V'b�#y	��� ɏ�)��%t�
=�V�o��k{]q�����[m���8��U�����v�B��U�]�qC�K$��)U2�J�M�X�Z���om��f�h�uc>:�� ���.͕��O���$,.)��Ӥ���P%��]lZ����eǸc�fZ��˞j|��5�8�`[:P͹1���K0S}%�O���OX�Hϼ��7=;4`�;c+�.��z��5b�Ǫ2|�� ��b6��a6�|g���~������J�.��.Տm���b���R	z\^GP�0����S>`�Za���r4�X:��D�����m�f�k]��Qx�N$k~�PK�>;�����ь�C\v1PlF+NK�k����;s�S"y���n��mw�%?5��o6�}
�Fkӻ!��������[�l"�Ƙ�f0f�����5�G�%�9OB]���H��d��c���ܺ}Zfy�j��a���N���9��!ݻ]�$��P��|�/���K�}����I86��Jޘ��ec�ü*Ө�q�2���N�Uu�����}�/��?!~�)X�����ޙ�:=��.��Y �I4C�2�VT���Z��شc��m'R�hJ�)��]saZ�T�^J�ݻ�x�֦�|���>�<����N��ϗ�s�/"����Ñ=���Ǉ���-�s�\���F�1\������$/� -�5�����E���u#Y.��rΰ��
��c�/OG7�	^&i;P��T1j��$e�y���!��4\sH���)��ʭL�l����c<e��l��CzQv���aښړ��x47=B��	�� �ó��|��P� �~ǰ.�}F�k�iȿ �%���#:�C6q��l��v�'�,�OW�B���R�loH��D>c�
��؜����O�u�N@YX�]Z��<��"��/�����(��A/�k0�u]�W�I@�V`��v��u�W�aG�+�eo|���ɻd�V.�"��o�͟n�C�*�c^y���@�\:�.2|�0#[�`Ⱥ�I�|��S�0ͷ6L����E͆���3��n����Zi�Q]ZJ��U�ߢ�gd?��_�q��z@�1�0��2��q��jnb���~|����
��|�7�[�j��h/5������\h�6U%��n0���<1�۱
y�,��/���򁏨L9�=���ت}}RS�(�K�`sHy�i�}w�~}�l���ѥ#�Q
��FU w�tu_U���:���J�O/z�{���h��ԙ��X���e>w��'Sϝk���\A[Rv�eqe.��T��2��S�{�a������tS9��C�	�U^9t��qTj⎐�ll<�7��x����r��ǃ)�Z�vӳ� �˅h�3v�Wd�O�%B*Ȟ��C*Z��\C�>�o�2�šS\��Q�ջ�#1�I�T6��m�� �9m����,{�Y�z�mDz��E�&�l�sۥ�#t>��Md$�Y(�����Uetײ��c.�k7�?	��!U���Z��7ܖ����:<uv�u��v�8�ə���;�9��gvRM�
�$nB�l��a*�uEW��>��x롂��-�V27wE�k>�u7�ԙ{��NiK�s�ޕ��u�޹+]`�:+LN����e��񾖎�#rD��K�p�7�m;�xF���Zlo[Ɏ��$�s���PN���B�:G��9+\ˬ�Q�4�K�	�N��_���}O��.�c3��p��T�M���1�#/����kD�\>��k��Z��k6�5�}s$��|�nSmT�r�YSo�'b�/1a��m��ܻ��2Vn*0�r��l14�e�4�2�[hTL��;���c@�:')���ئ^��k��ވ��:9�x�]Jw!�Y���Ȁ�U��hW��%aU�;�*՜�u�v}��[���4Q�d���Sj�$׳0+�-�}��c��)�fč�do������I��\i-�vHR�ٙ�L�܏,�qob�1͏�m�����^-p�����N[F>�����}i��R�<�NYk�#�]�mXp���ۧ��RyPQ���.|�¯n�{�lxvY�\�-�[����v޻�<׶�+y�t���4C��:��ۜy)5�u��;HMw5]`̽�am[V��W��ͻ�$松Wv�6r��X�ɧ;U(��Cta�\�6ɬ�8����x�H�k&��6��)Ǵ�{&���]�j���;��u��.w^go;��Jc������{�`z˫|4q�m�o#u�v�z�����Y6C:���-$"r膒?m
����.�ٮob�]l�9\�Ļ�����;�=y����u��mm�X��݇d�܏��Z��i�6�r:T�I�O7q�%�����U�����a���|��2�l܍�{u�÷$���76���ے��x�-g��R{Ǵ�q=���٨��7rnM�8����}��i��"���	-o-ƛ��!:6g]̾Y-2��KqU����	�MwqM̰2��\+)n�ɛ����0��}��łwL�^nV:f�'tGz���� ��Vd�[�w�7s\]��Ar�vZ�%�a�xcZ�du+5��eY��מ����=X��8\�l��cE�8Q1Sy�Eƨ�klQES��*�c���<}���ǯǯ�����~�_���ڪ�n��ADƵPSV��[ji"��J�g�IED�E?s��j��9����ׯ�����~�_�����⊦�lAAMQUETSELULbqTW͂��uEUN-h�%��-�EV�m[$h�j�"*j�
�}٢*h�Ws�譍RD�T�A4�kPDA3SQ5,�RDQ�[���j
Ӎm����^Z�������*��Aj�m��ML���UN��ƨ)$�J)6��O4m�F��'�6LEF�ت���&��(����[5U�j"�3MU���Q��M1%SkUPD�E�hѢ����ffh�s��(�ɵ�4E�M$Q�55AMSh�RSk�QPRAm��*�����ō�m�X�&�D��#��ן>�=o~�{��.)*u��wo��hܛM�ߗM��y�d��P��Ӽ7��{�6	��V���6����"�W���{���3��R���������~z��v����"��y/�<g��i0���\���W(��*K�C��ُ���KC&�c�^���`���`�D@-����xгnd�%I`mt�-�I�vq9r���5;��F�������� �_��r>�4�@0cB`ke�K\��`v򭷋���Q7IS�5��]%�����|�ğs�|�|`0!�� h�� >'5>�e��r�CPfL.Z:F�B�_�_z�f�V����]5�h�4�j[��@��^�9�"]�Z!0�Uf!�y��(������6nڈ��xdm�!$�p{e����`����p/W�K���ګ��g�~b���(���n�0�Ⱦy�H~�PiD�0��Nm��+��\c��ڪ���2��Z����:����_��,@��Y!���K�%�z�{�]۽��^d:2ܵ��4:)�`r��$��K�j��oT�5.R�	�&��tJ���t�m�l���ӪR��o�p��8�欨�sC������X�9־2Ttx��.2���'ao�,��2N�IW��I�-��Ӣd�ch�VI���[��q~�[{,(��h*���KW��2�c{�_��l�e�5]c���E�*�X���_�ļ=c_�`��Y9�켅��6DR�G��9�9�s����p���T{��?�~��)�X���	��d&T�P��%v�����Z���XQ����,e5��$�:ځwyLv$/m׸4�_t���D&<^%9�)Ė	�B*�ߣg1�s��:�0	�:��E_��3���q�~�G2�,?pG>z�@BE�oD$�^%�u��Lh�&��1i��Գ����G���]|�a!C6H�L<1�|$J����zΊ.�Y�]`n�b�W��y8�`d�'�5���^�+��|�:�J���N��� y���_o'qT�]�ge�j6��9^�{�9�m����9ja�c��XG�̛��DkuL&��zzKх���7q��#��2�7��uz��f�P�z sO��ך$v@qB-�O��c>`ѯڹ��M�I����CG '���?�OJײ���k���9��o�8:�H�]X�2�:�{c���Aߜ�M����@�f�z͊d�)Mɔu-�ߧ��k��|`ۄ�ʁG�7L�к�W ̽"b�� p�Na�˾s��>�d�l�^�/��=%�:����x'W��`�(gl[׋�`J���}�ud=�k2s�v7`ȫsS#�n��������=��L!����}�\*���!!�ӱPv�6K�7�9����vh�k��TP�t���\ѡY�N���{�Ք˧H�!h�4V�א��fF�f��B�H!c��*��9Ȋ��W~{��}���^�� ��Ӵ;���4���~G!��T�W*�-|�{�(s3?LK{/����x�Ӵ����EC�� �--!����<4��ћCZM:�M� �w����D���LҼ�y�*�!������O��xiז{�A	�ё��;�ݝ�nvbm�6r{�^8�LcO��*����y6�u�d��Ўޝǯcռ*���vC�Z�mV��݈��c�FG�hOV0�bv+��Bk���A�MW�i=�]:¼z3��[�|��ʤ�d�ڵFo[9��+w�\n��@�B�E{%W5�A8�r�d^�J[���M{��J6o���b!�:�f>g�{�ȷ�x��2LJvl���O���/��<'Eш�䓻����ݸ��m~���J�;\��{���ȸu]x��nLpe7���IwO3�(�%ri�����\�q����t�˨���j�sj�1e�>G�e��@A�"mLpm�#uZ�=s{��^Nj�K�].�,�n��Qi�c)�./#�������鿀̗��^������I8Q�·u�y��
u�)��i�����~�ͥ��Tb�7�T\9�/E>4�s���H���v;#4��l��x�hU�eh�s9�ΜB6�݅��Hl�������-��_M�.+��ן�P��r�g8E ��ߝ;�������}���'�i�9N5vE�jF��)��5��>1.���DH�f���Q���5G�0{ǝ�wf^�w'Ȟu^�����M[�S�Y���E �}
�F�2��X"��2Qկ�No;�Z�`ϡ����K����r��a̖Y����O��W���	�z�����T�z��9m�����Ax��?04�7ʼŪ=Y�#(f�o��<)��->%YY��yK
�yB��;Z�?r����xg^�Y�E9g�V�@��u�L2u�9Z0]�`���ٔ��Fh�W�3�]������O��K`h���3�w[�o6�梿AD��E���T��g�x���7��YڂS��r0����<����)ܫswL�A�����}44�V#C�[�Us�Cvm�:AƬ�JZ¬��3���8!;N�A�x�̹���ʛN�L�ս;��2pAO>��za@L܄nr*ڼ�O����z	e��V��U�����(.8����1aȩ���J���Ϭ9�2�s���Y6C�}�-y~}����CD۰@��E�;u��or��wK�j;:*��e �Ջ+9��,�rp=�[��x�ξn�E��@W1&[��g��cK�ҹ���f�ѹ�'A�ބ�m���n�9�rn�Ʌ�d4���#�SŐ����+������� ���x{����b���+���>}�]B��*�
j�q�^��\cg�E	-�����u}��O�����Ӟf\dgRx��p�k!��^���ߒT-X�E8���a#�-�P8ށ �4� ��4w��Ef:R�ؠ7*�f��7:a�wQ��K�����)=��7l�;�K��)ؿ��̴�잵�rp�O���08s��	e�fo�Jy��m�t�ny�mx��?n�c�e��\Y�����w�E�e�!��x�QO?T�F��aT*�xj�[�ĩN4�>Z+����Q�|��WQ�eC�xwo��"Yǒ�yg�M_�w��o��2u��*��Q:+�T�Z�v��o7Y�����D�t������Ѕ��`��=05�oMS:��8k��-�٤�����	{k�����P��9��+�^P �Ao��?���7-��uqf~@WQa�C8��6˦����4�3͠�/E�3�2%� �`>��M
ƛ
��/�X/<ħW0�u�n�6�d�8ė�a��Ɉvâ-��#
���5{��`W����S[�2������������9'���1K1����/��6"��'#˜�3,�j����+����nJcv���d�;�;�Cj�|ծG����j���S�i2Q�V�uwjW�-2i�wn�@3���.�����z�Pr�Ȗ��#��*W���(T	���<��T[#~ݦax��=����H���'Iy�Q{V��YA[r�D��u�́8�B,��H��0�A��|�;�=���g�Nk�LS4r;�����p��M��d]�5q�NK�1L�7�<0h0���m%�3��7-�ú����~ȿ/ޛ��s\r��FTe
6�����	�����E1�?�/�X)�σA�{ן�$�-46�57Dt�Z�V�KsWA�o��ʖ*��vл�ջ����m�����>�}�H1�G�����2��9��<�cҘ��W�4�����6^%9�
��5B*�،�ǭ}Ǆ�a��6Qz�)�j����cF:!�pO\��קze'E�C^[�F�Y�P"÷Kn����
��K��c2�9n�8((f��Ba|�:�o��6Б(�}��0�r�E��n�{ß2�)Eg-/h��b�K��p��L�vll�uL�"�Уc'qV����=J{�kZ�cF�5�� �/]���PX��0�PN%�;`>�C�,��鏃�����>�bW��?cӱV�3���mY��2�w�c����y�/�q��O�p���	��ٵ�n٬Qڀ���4�_4�l"p%>+N���h��B.�f�����6�ܒ�u��Y��l�@2+E=k#!��r���ܰ��H�5�cՍ�ss��8\�9�� ���&s�B����|�����:}����s/�.�4e�Z��3t�w=2�C�?�{�#��3�m%�8̭��gB�}��=%��A5�(���~*>�dz=K\N5�,�Y���0j��녵x���صX��΄;'M0��o>�Sl�9Rca�u>X�>�z��g��\�b��(k��ǻ��j����ᚆ�t�$�:�^Ļ'���w�{(�[��$8��L3]�:]A�����v���쳢^����y���q5�Qf������
�9�yt{��9v�
zc}o�{#��T���H�=N����F/�F���W��O��?g��5e'�Kսn�EuS�5qO[��G5�c+9��5�%�QYAW�0��eM���Zfj�;�3����*�����E;�]���aE�)���ׯc@\U3m����`Y.�Fl�z�o
�E;쪲�4�,�ջ��N��`fp���w�c,������؝���x�M��PdԱM'�]:Fc��s=��M%Y�Ooվ�ϸ(!�;�C��&���6���\#�:�JSL�i[��S��-e;u�(�E��璸o=�ujgp�%�(R޺��)��/M:�ݱ(P�c�+���p4{(��dp�M7Rձ7Q{3���t��7�¬e[�*�ʾ�nֽ�]��%�n��D/참��h��t+�g+m�T�^�_πO�� >|�q�<����cWi��K�m�|�������On�$>Q%ٲ��L�� ��y�?D�I�ɘ��X�Q����z�F�ג�L�pm66Gd�lz���G��m"
Y����Τ_S0]�]�L�=c;{��[fNj.�WS�+K�yNRc"�U�9����#ϲ-� �z�M��V�4XU��wk^U��Q{�]��&�z����R	z���H�0���-��jm}�M^FBi}a�`3#���ѡ!�3���xn׍1-۝�V�w�S��ׅ����砟�H1.��2w��0��HF�j�vP�CE���L��U="��Gu[]�JO�c�o6�|�j��8ֳ�mls��;a8©^�i�s �?�1�-�:_�*���/�6�`��cY_z#��^CUK��%��ƛ���L�������]X�Ѕ=�~Lp7�}L�[�s~1�yHGAz1{I���f6p�������i�{���D�sQ~�Pw�xg����0(->���b�������U��2<���e�8���6�b�W�3EڏK�i��$�ߕr����$���'rf���~�OHi�m�d?��Ѻb,��!㷇D�@q7n�Yu9��*�b�ofk�2Vʗ����?��~]Z.�Yu�y�|>ӯ0���5p.լ���U�Ldn�Y��"��n�ݚ9�㘛w�T�[�*s2=���q��:6�=_�S?�*��D߯}=�s��z7���w�O���zn����f�u�9�����c ��˴�|kO\�o�5��]gc��ˤ�=z���P�<!0�=Ŷ�ت����X��A��@� Œ�����:f3�>[���O������_~��Rǆ���d�$���¦nA1�4�� �G6.�	�L�omE��}��F��i5�W>Ň"��e�J�?1v���G�=dۓ������"��t�RsQ6�Qu~�
P�0���8�:���x\c<�-��C��>��L��{W+16tLY�L�!]%���Y'�b%9��V%QO�v�a�������(G��U�C�)O�	�1�ô����f��n)���T�p���"���A"�vl��,�T�n�)�
z'3����O��b5�:	��
�/�K*����
y�Sl��\sw��(FcT6���XwSA�����Ϯ�=���t��?`�4(�x�aT,�熫W(��]���Nyn閈��Vִ�2'�M!؀X��`!~=�y2�~�<i��o�d��P+꾹�
�����M}uz�3Vتw�
[�����:���_���v�5m5�R�5gJ�+��̃-گ���g���������}�&�X�����u�	.MkPh�9���a�5NN0 �6�$��P=s5�ɍ"��Qn^;��ͱ�N�wxm����
�9{��޿���}w���yv�2����_0-���n�|\0g!����Z`l&0�[3{ �e�5P��н�0���pl=+\�%銨��lM<h%�9�8/�~��w�MN�V�W5Y��~
t(ǘvc���j�����"��4� MI�G@���g2dK�9f�1�鸺�Vԩ��:�� M���#$��A��;���t��?J�O��w�{ċ�m~m�׫G�(2>m���U�j��΅<���`L��yS��Tc#�wS0�y�5� ��T�.$㞥�oo�Yy��PˬE��,&�喸fМG"ˉ�)=�j/��cL�~�P�7��s���h����E�lp���!q����tS>,*ä�c����h���Ʈ�ek4U8���T�C�L�-��l���veK2�	Q�C@��skb��M�8&Z�%��Ȕ�Yr�]�DA�(���n��کnnr!6o�ow�&W8�R{��B���{�ᦞ���&`�`U�.�w�����6@��� ����<�:���ħ7�)�j�U|��^�z2Y���`Y�׹Y&�6;�t�c�۠)Ŷ�ru3���̮�sc(e�����-�%do8�mL�t�m�$k]�ⱪ}(�M���ا�1�hkn�+H�\2��]�q��[1��U�ܜ�L��x&�6/��ZR�jňk���.ɜCrm�F��N�@��ru7oN0jF�4p��k%���
��b���5�׹/o$y�me�VR%��oCRtώ$v�i��Ơ�-P�F^)�6��9�B��7�[��x�N8�u�K�8��y���a�n�I�c�mkp �mb�0qK��kp�X�$�l��]f��z��O��yQ�v��<d*��ڈ�V�P�]P��w�n�^�K9t9�r�.���̱J�s/(8'��˛�0rf��cC8�����u��i�C��U��^�!����!!�*�2ָ1�.�i7k \B���7.��,�-��Z��5��vvKm�g�<��]a�-���Kt^�k����gn��l(*oNw�6��FuqH�p��f�mQ,n@:�����̈́�f��Qu>�s	��T�0��]��b`�L���&�P�4i��GD��0v����v�h|��A�Jӵ5�'5;`��GB�f�z���/��דZ����q�;�\��qcқ}L�l��]��[��X���7S�h��0����صݷ����5h&ts�2�h�v}.nD����y�w\�xʆ�&�튑�c\�l�$ ��ۮ t�|��G� �$��$
������Om�6)kr��<o_`�U0Z���B�xbY|�[M�S.���x���rA8��e�\�{HK�&̘�JVM^oee��9X`�pt=�ͤ(�k��luo���f��gf�LS�y��[Pʸ3&��i��,�8᣸�u��8�ֽ�+��wh��E�v�#���ǂq�-�]`�ٽ����aɨ��+M[i���.Y�h[�[W��$؂� �� �.�!�Lg�p��ߵ]\�W[3[�A܍�r[8]��Y3lM��!-%���K;���Jъ���D�|@����=#{U#Pݸm�%\��'%a�}sY�b�++O��K�
CX�����u���(.�������<����8v�K|8��e4�0Y�#�$:-�ۡK�' �J	N��{�HZ��8�蜅���:yqg3$�<h�9̋b�����k2�{��_m�A%&l�(Cy��n���Xƺ�v@N쥦�.N��*k�{��T��7�]��ןn�\=��I[�hf��.��h��=K�HeJ�ֱ+���8���|z���N�|d�!LS���YmHv�[�M���OX8Ē��G�-y���m��ڗZ��Lf�uh�}b˘��Ӓ�rj�X���@��yqT�ݍ!Ù��:t�{��2�!�\&J�t�7�K�9�Vqu.�M754����}�	P��!)�UT[ʒD�h1d��AF��MJxn�!$mz��<�y�+�����}�h�*9�jζ5s:�m�i6�IAm�j*����(���
}���������������~�����ሊ&�*
����HڍDVƢ����+�5M�4��LO�<|}=z���?_������??�I���4
�e���b4j�i��������-�UQQ�����b�*
������cN��((b&h�4���CU4ź�1RTT4�I�7""�lTM0UkU5IHA5CE�IM%5rQO1�$������]8��cXw9����gDEQAU��UIE3��`������b���r5DDIRǌj����9�p��
�*+�t��DST�UDr���
� (������A��UE1UUy�F���-���8�Æ��Z.N
�X)���ӭTEPAD��j�(��*���/���m�����2�q�[=|�T���Z��D���"��tӖu�����қ(`��Knu ���o�i;�>�9����ss��ׯ����\�(���}oܭ��)�V�Ŀ�;�amI���!<�M�oD$�x�E��)>83؍j}B+c!���c�fZ�ϑ\��v}��~��P�f��Bk�.{���C(H��&G������;`���K���Wo��S �T7Q�NY�6���L�y�5�M�0&A�Y^X��`z�������`�->��߿t�\k�'���C�������S%���V��f3��<>�
����{J�~EQ��Z��3t��;�k�m �8x�d�#Xq�a����6�ֺ��WE�^NS�xm���l�	�`K��c��PK��g�~Q��/rʹ	�`�Yj�EC@jLn�,�1��2������L�v�{Ίb��7�/zc�n��l:�oI�f�Y�j ��Lڮ,3���́p�4B/"u�˲}��!�&�Q~�1�/�w"۟����	�3 ݳTz��p��|o���E����Pl��q&10h,&C����;�U��_5�_u滢��K��1���)���x����$o��g��_Ln���)���d�{d���X�A��A��ק� )u����39�5�qcq�RPj��B&��ʙ�e	)?��.����Rk&�?B g��V�����s�uc��n���h��>
�s�<ִ>��#Gk�r0�XCM���[;#���~�9��\��s���$�8C9ʉC�<��sk���\_�(�TtgH��f�S4�d���e(r���)>xsͼ4�yd����w�{�+��ғ$�>���p^��^К�Iz��cJY�� �� -�`���������z��i�LZ������c[=p9
wBÎh}`й��гҫ%~����x�M�� Ɉ�{�Ӭ��~�?F�#	�}�?1�2���W�d�,.b!�.�VJ�nwA8�Q,��!���6���:�ga���O�'�|r�{�=򿼰���!�S�cg�?&l��`��H"o��ɮ&u�c<Y,�}��M\z �/V�(��V5H�EMMލ�����ฦ�$��Sk:e�����3���}��\|H���k��)?I���ksb_m��_ˠ/~��;&�eQy�U�=�»]O8Xܽ0Ct�-e��۪]��&�z���2�K׷���f�H=��j�U�&�K70���B��i�B��W�ẞ7�[�9V�]�"�BԎn������=�"q�e�I�ɺ�͏��l��X���3���@�X?��̟�	��N���-��mw�)?5�2m��m�p�`r��6��c,�QvN�^q�
<��d�4;����l�z���ٱ�n���]ѰY�8��5�ښ��̮�s`6�[t(�T�j��h9��ꣃ9*Z!b����z�]�������.���L(ҳW��4����?j������z���k?��}����q����e��ʡ����A����D����|���ʢ:���y���:sis��w[r���+�j-e��~5��
�ض�_U3	��vz��tɮ[׽.��s[L̡�%���u�{HAZk��l��
�������k�G�����O�>(������� 鬬���E�C���n�my��A>�~��_�w�J��g������Kf[_jq��s�f�sT���d�i�Laubb�)́�>�����pJq�j�#.��Ԟ�\���ʻ�0=�6����)&8s��+vyXW>���XV4���q@���a-�^2��2�!��-�����3���5�-��� [��P6tF�v�yas7 ��TU���I	�ݖn�&�"�WE��:����>�H0�}ke;k���J�??���`��v]ɭ�X����sD��8����_��
W*�5�����b��.1�="z�"�^����n�s�k�S��.G���_N<y/ߗ�Nl$�Z�*�qvt�	�m
�ӏ��VrU:(�K��8�|w�ı�-%򄝻^�C_��6�����M���0̟J�ծ��.�aKev������@҃B�$���¶b�PR���GW��5�����(��iޡ����E�:��x��7�s`�}�j�w{ZfN1�i]K��z�χ���� ?����T��M)��7��q>�!����=��13R��`7H��3�恱l�U]L��2nL�r����U�����A9�0/"�	n�v��Ⱦ�)�S"�s�kmL����;6�߳���/m~��*K��A�@ �k��ϒ�xׅ�L*��熷�K9f��i��9o(���a��C�,D;���D}_6?~L�\��Q�����<͹,�sQ�w_����K�դA�t���h'�P�Zz����*�.gtD/Y.�� �ʸоn�n;���S���ʣ�H[bu�����0��<ͰgwwO�����1a�2�u^�f9"����Ͱ��@e�X�0�9@���io@��^�9�uAv<����y~}�bPD�?�4߭u�JN��v�κ,(q�/D�7c�&e�n�(��K�ok�j��h*n��΋˼ygDawhO�,EE�67i�^=����$�T9�ս5ĵj�Ξu];�0/r�wB�o��}_`���O�Yp�p��Ƕ��֯ ��r�ֲ��3S���,�֮�Y�b]y��xFuoF�ѽ-��i��4v�5*�2L��jF��Ie@K0���(r8��5S�.Q��30C����4`Uvy����#ߒ�.�u�b��԰�YNU�+�.�wl�X�mJ:�,=������79����9� f�k=:��-Je�0w�������+d!@�^k|�M������a�s�̖�J��O<A�OK�]���^��1ݙ����]��*Y�(�Ty�׷�M�SؖxBmf{�	rW�]�:���ū:�O=c[��T�jJm��BeK
U��"��c�ǫxjGwBշf7iu�����Y�LYPQ�#\I|���H��|���B��x��ʔ�5B*��n��B�kWw����V�2����)s�w���·�ٱ��nb��7Ͷ7�v�k�\�"ґ���<᪢�c���3d�!0\��,�1��"_ʽ�f��6:�˚a�b#�U���ߛb[�چE̹mwSJ�}���L8��}B1��(�yOuE��x~Y��ͥU��YTa�Y�O�iAcAt�~j�q.���C�CM�u���*Hj?�x]���Na�$D@��LIsRg��'(]�T��=�*;�̩��di���d�Ck�3j1�]��N��.}���hR��D'`�����ked�0'�c�A/rꟛM�x�.����eo��nh�u�b]i�H�ǝwb5+3�����Jp	~J\��gd/�z��cϤ>;xd�y�S�dpV�}�մ�U��
ko9?�5˫��U�;kq��5���
�ێw<�Y�%��y9)1J]}��$�� ��{��L�O�� �_ >'�%S�<]M:�� ����x!vmt��٬.4ޜe~���:ƈ�|��}8�J� ��s��f[�x��́�n*�G�s�a=����+�=�*�a�l��E�S�1�~���q�IV�����CH���1^��-�WX�c>�x�Xhl./\R�/�����R�&jK�X�dv�cFm�2&@� �=.�_E��(�_��_��f��Į�ߙ5:���3�`/K�z7�CZFn*f���I�Y[A�;���O��o>ז|�j��k�T��ż_E͌�_�KP���W�����E�{�*f�ݔ
�ʖ�����i��X��ȃ{��@�{Xn������VH�x����)���5��y�{x�M��Pd�J}�-�h6m�
v�WX��;Q];�x�o�[�!�2pD��e�4�p�l�(d���'�uy!�=Ų�ż�z���Qj�'bX�F�]���Ơ9�<������^� ��ʄp�D��]��B���f�4"6㽚����N���)��L�#I��n9��.W�<�i��n���i�E���bϺ]v$]���Lf����U�n<v�c��-�JT�ޖ`�������A&1���zp��ᗹ=�r+�W
�7ͻ��:�����4�,'��#{�8KW�mKz��&8:�	�;��u6���n���M�O:���=}���s��;��߽߷�~���l��{<�|��I��NV7H�Y���5�;�\H�v���k[�<���W��@p��߰Jh�1��od���_���n�����e ���#���0�B�m%_f�:�=Χ��8G��~z`xr��������Zn��/jF��)���g ��+8����!_��/^�G���.�G��_E��a��$;z�~����؃�hϗ6�tę�{�c��@�[�ͳ��!����;k���g|�"��zpZkgJf�6&�����Nj,)���V?{�շ�3�-����4y�ZBb����X��"<�%���|�i�u�@��������)��23L	:���j �r�^ø���;<��D�z�l�{�IsA����MF�V���g��y�^���C��v�Z]�H��$� ��9���jLi^�Y��ە�Ŷ���!���吉�Ρ�T.��ͳBt�EۂS��W#.��q���R�1�"c�[_:�o�%���B5�c�$�5��v���A��A��.0�	O�z~���q��Z�����޳�RL�d��N�Z�Q��]���'ee�4���Z�9�jd���l�7�����OTY�Y���i����-p�֬���9�St�[�+4�|�C�&�l�Ǭ��Dg
�{p�a�W�Տ�?>K����7��ol�.n�R�&u��g�ג0��T�<�@0?ܧ���D7l{ۛ�ה��v�w9�1~K����?z���>���Cr�]Z�@�c�W��������sb$�x��;R�l�u\���<lu��o-b�l�/^12�L��W�QoS�l2򫙄k�,�}N��J�ʳK�&�=�J`����-�]�'.��IPT!IN.�gN�[B7��y�gLYxS���Uܭ��>4c�H�H��n��3�U&E�&Hl	.��B\n��	���h�f ���K��v��w# �JF���5�d�qY�jo�J{��H�`֪��ٻap���"�;�����Fx!�5���>~=�F��aCp=U��|�>gcN�x2�Z���.���9bB�P�|���|y�B�v6?����-e�g{�T"��e�C{��W��\�㋱�QaV�y�� &���GO��8<��߿e�n@l�3��?�[����Lf�P�nd��ҵ�r^���a+lN�sۿs�
1�JQ�Յ��:��^�L\7��ϡ�����;f[ga=Sl;6�'!�ʜ�5t�rm���2�}M�3^h�X�Q��`�d���0A���_^��헗��v�˗�ʤ�}�9��PH�)��˲s�cJ%�"5V���\��Ay����m N�,�B�C�?������wq�Y�������P�M0�3m�e&	���B؛t�8L�si�_���n/�섎v�Կ^��0�����#-���1O9�͓z���1%�vn���qO3;�d���R�k� Au������Fz"���ݣ��d\c��f/"���Г<��WWf���E�!vi�CH�\-ffYm�DG�'I����1 ��#���ʧ;Ƕ�-�ZF<�D�C&�f�Z����9�?cy�=��F��2n��b�=�zg��Aϓ8ڪ�b t��uv��l:�t&�N^�5��B����2����E���TE������r�!6��Z�<�Y�S*��c���Hl�0�"b�!2��P���]�+ǣ1�"�邸����nX��
�F44�-�k�DD�Ux����nj�	M��9�T��ݤT2�;�׀����]��p�6�{��\��^E=��am^.�|�	>_H�5�ޙIӫ��a��T{e_]n���9C]���+�L+��+�S��'� f�	�ס/���	:�����"i��R��ƻ�U]�&`>�Kiz�݊�J�^�7}]i��� ��^~���oS~�H^���w���Z�c�m�{�w��X�o�`_��[ �J��#���j��u��ʂ�ŚS:��!����ȍ#��*ۧ�K:" �}Ӑ��F�f4� 3����ws���n���V>����o��Lb�f�/����6�;�B
��1n�|��!��Tі/7b!�%������,��~OI��J�g�Ʉ1���,#�А�}�$a"5�[������~��z��A���Xg���.�F^�F��P�z�l�b���5J~�Fi�p.���̅,.X(�;��k����Bv�2~�ܥk�PKܺ����:��Z���u�m]�	��ȶg�!�>���-0h��1~(���Vt�?X���W�Ͽ,�',yi�d��._��DW\�m7h�^�u�9�j��|c;0�����_�S�^��>Ⱦ�헣k8���;�Â�9����������|;�}>����4t���\D`t\H�Se룡�iD.��}��ّ�?��c�����C|7����l/���[���8S�e\���_[�-�I�����P_��kOb��U���#~��D�ޒÊ�h�%�H�i���X�ЅR&T�i'���z�t��B�Pza���G��~�&���B�1�˒�j97%�����w��6��q�E\&qwBs��E�vc�@��YX[����J��L�욷|�XW�!mR�!�	����pI|�-Y��h���x4i��`Y��N8�D�t��df���X��.��h��9�VPHRl���z���uƵ^J��wū����ݎ�=]��-��%t;�fe���x`4m��ש.R5���xJ=؇R�º��g�8t����A{ )���]]�D��+yFc-{�Kg9\��{��?�(s�}�*s�-��O	ZF�[t�#����MQ�|�H���,�To��|M�8�gq9	�6�-v����3�d�<Kc�r�+w�𓶰��c�� ��4�6������Ӻ���G�4 n�cp�v��U���j]^��l�˧��v�Xc:j����E�b���&T��̺0K�I����	\�F͗2��Thł9"�*y)�z1#���]45��+5E-�+Ö�&a߯W���@�}�Z�R˸��NR�9=�t�Q�A����TlͻA�NGI ����E�ʾjC��:G��ws�L,�q�mi����z�Z��G���E���3FZֱ��Zu�qS��wu4bt+ۘj$o�n��]�����ͷz�ѡ��h�W;o��$tq]�mݳ���N�G�H�=.�%�j:r�y/;H��M��3A��V�$-W:!/�حB���}ܳ�t,5ǟZ;�ٖkr�;ou��=$$�B��1֧WH�'�~�SZܤ:�H�,�Y7ǀ����r�O�
z�"v�����e���Z;K��{����O\�[А!���['G��Y�� Ý����ۃ�����K����;u�� �㳊}0]��=���nf�o�3�����;�=Y��5,,�1^SPBvf�h^1֦9��]�ד~14F�g�V��8�ڭ��ϰ�S���z�W�Fފ��Z$#|(��b�vm)9s0�w�[yYtK��1Hsۥv	���c$����E�T�-�%��sV챻��m��)��6b4�J9%�Lcܜh��'7͙Su��ݷ���#�e���k%�K��6-�#�S4��'5��f��C3 �c^�f���=s�@��C��D��.����f+���
j�Z y'K��8�s��O�.���*���{H�d7@�$gzl9J��6Zo�A\8��zo!��\��,w�{��Z�p;�u�Js�1e�h���G�]���4��ļ�D�]�n�EW���Ն�V͸�S�*�B�Y�ɋ(�\<#���9N��@7J���/KrGf��װS*�Y���ѓ��B��f5�c�_gT�wX��r�k:ѱ
U\��Q�.]g�hV���~�����74��9���P�c�)Rӗz�w
=�9��`��d��QN�I �g�iV�Y�zL/��:�
0\��pv"�h���?k�w��uUQQAQ�AESM͚�
��&���fJ(g������z�~��_�������h�"h���������A�E�TT�U�Q1Q����*g�ǯ��^�_������~�_����
���f�~mP~����EQ����(�4\���(&*"����j���@EZ���kESUUUUM4�AT^s�&��	�m�f|�5������fb��bJ*�J&"�$�(����"
ii)������(�T�UU�(*&���ԕPUMI͟$�y6ڦ�bkX���&��!�E0U%LLskm����)�*����(���E��PSA$DE�LMG�J�cC�3'�ii����&*�Fb(Z�����ET�D1s��k�s���
m;�{MD�DT�QG��8f������;��,Cc �Na��9ʟc9;�\l����ĸ�n������ɶ%+�z�gYǩ��uf<��� c�[�C��7���s;"��Xqm�����X�ןO�+�la�6c�g��huۋu����q3�+�3�i�>[�8A@�-�� #�\�Q"���k2c&�Α/5.�7�bX�F�P��w����=�Ǥ�L�ٮ�s�wY���:�����ЁQ���r�9w���R)�$i5�;��a�~q��\���W1����t� xo1��4Zf^�A�����w7�RO�!1Vt�4Usj& ���y,�����"Cr������
E��:��Lpm�/dJz�R�>�34&t��-?,e#�qsH׭g��O4���mW��:�����l!��s���^�;�M��Dх��j�cTF4*��7�^������]/�Z�`o�FxQ�0<5������A�]H&��'AG�$�6u�1'y4�T��3&upw^�I���b�v�/���o$O�/�{>r儰��]������{HY^s<����ߖǤ�3�>/�Ӵ!�dk ���?Ǐ���iO8=Υ�cq��.7-�5rx�2��D�����Y�c�;F�L8�:ds��dȢ�����،Ċ:ws��N
v�����V;B�T��q5�b9Zв\6k@%�\����v?��P�)�!�Y��4`j��0˛o7R{�^�����s��e�q��u.��j�X��Δ��5�8�
C��^u���c��^ýsӼ��9���➖�e�]S�ak;*<�
߮`k#Y�^Fv8ėj�.��	�w�冉��������ӣ�Y�
�$���/�t"��+Y�^�������A.ܔ����MB�3Z�m�u�Jv\��^�ͼ-��x	A�S�"�Us�ɶ��Hx��1�l��Ţ_�Kڅ��{�����ŕ�*I�Xt�D=��
���F�D��a4�ӿ@ke�L�-d-F��:�PO`*�,h%��^1��E�V��@fp��sb%8�mi�UJt���"#��vU���Y1��D�^фʖ*�Ia,r��n~`�A\����؛s�^�M��3��+���;]�^�BE�瓁��~"S�IPT!IN.���ape�7%�2Htw�j�N����<�$T9�V�7�Α=ҩ2��%a�E'z�q�󨼘WOk8�ۗ�'Ȯz����A�#��?T�#�o�K.�0�/�J}��xt�u�����W��϶����e����Ы���w�W�iN!3GEY��;Vܙv��}�*�=P��8�����9��v[9\����Z�x.�����pC,�:)Awm�"�Mj��n	��:S{cʍ��hr�`�#�Ub�Z�Ko��Z�~�������vf���M��)��� ��y^nF(�;��=6��2dCpeOS�¨R���U�啊)��j,6�3^��Ϻ8�7$UC	/�s�נB�����w���E�Ǿ/��SE��$�xp:0����qH�E�]<�n�i6t�ܩ�}���ҿ�x�l@w�0��<�b�2��={�-X�8��Z�
�^�KϹ�n	� ����/\ϪZ��g�Ȝ�T�s��8^�fp�Ƙu�C�+�Y\����D��&�	�f�D�F⻅=|OlM��F���DO�C3�����)���~��d�k1Ļ<ު,(q�.R$',���l���\�5�4k�3"F�e^�Ο��4>� Ol,EE�7�L�D\�t�MoeU>-T�Ih^d�h)�G��.���x��K��Ϡ����Ӥ���>���J � 5��u�g�8Yom����
-]���%�?
�z�6����5B����-s��+�.-x�ࣜ(��ǱU}G:����{��A�r�a�):��f�0�\������xLA%5h�_���NLX�ݓ�,t�4��U�ܚ��$�Sr�75} ����W��4g'����,Q1�|r}�ӈĖ�h���I�D��Uђ��M�w��zM���&�ٓ�Ҽ�ԋ��gb�N�Y�I�£�-G0�?�;����y�O�y��{�_t�޸9�3�q��(֘q	־2]�R�x�M��BeK
U�R꡹�[�mTU�sEGV_�?a�-U�e+(����cc� ��5�m�BSrxNJچ���Ʃ��LF��+a,��b2s��l��)���Н�B`$��� ��5�ز�?fTJ���݈x��&��x���E1�
4�7<󆪈O��� �5ȈL�K�e�Х�ˠ�p�Fٗx�=Qp��<���(��ǖ�_��:�p���zd9ف�u����2ks�����ɞ�Q�N�|,��z�(���9b�:Y'����B�NYSV��ffxڬ<�W��	ZA���!Y���cOW��l�j�(]���е�
����kX�~�.!˷dGF���n=��#)`��:���Ķ*�)��M3��w)Z�?�w{cW���k(�m�y�������*!nl?a��.򁣫�4NZ�������}8���Z�Y-�nk�k�L��	O���s�f��A��F�fq��9�ߡ���xK�|�Vʲ�ϑ5l�:v���[�M��.ǵ���^f��qv�E:���U�ez�5�a�|�ȿ>�-j�;�C�s{lWZ:(�a�H\��bY����u��d��-�3/'Q�n�=����e�o5.�Է���=���j��:��, ����o�˜��A�|1N�������΅�k��5v/SI��."0:.��w��^g��-��өt�kv��������=<C�4 =.ŰS�F�T?PȖy=��Ӹ��t�ۯW��z�!l�B��رO�^���|��Φi��,:��r��6�-<e[Rf"��7x�|E�]<2��}�H�Nbc�ϗ��>\�3Q�A��Js|�uvmh�\�N�E�s��}n�*�t;gK�=��`XC�,�[����=���w���-�C[�1[SQ�Y�N�6��w� c���?=��M<�fЂ�v]���l׏pk6�ݪ��ֳ�փ;Ȳ�\P��t\��e�K�zUn<Ϟ��D�'�{w�H0:vk��̥�ME��O�"Na�
�%��2K�1�=�)�P%��&��F�싇\�˒�2`���7���t�r5�Z�i�6��0Y{<�j�ic�LU�H�C���l,$��f���)N�(�/|i��b�LS/4�=Ўm�LG�>���%��K��2O�����H�oz-B0gPe�%�^g����w����QЈ��o-��d̹�����9c�Tw(6�N�����Z��D�sJ����:�۟V�\�P�O<Q����ħ���*n>������5�k��/�F� �2�.���,U�x��L��Pˬ��s5�8� �o7�{�7W�*����~Y4���"�B�`�Z��!�;�.x�ݾʅU�\�$a��ygB��{��3���h��ӯ��=F1�G�ûF�w�Hl�E�Lss"y�Sve�~g���;��DƬ�\�66|`!��͊S�U22�-ݙ��4�����{�b���4���$]'~�����W����^�د�v�_]��=_=A}�$vƲ
4&-̇u��k��
}d��ۼchgXe'�4��D�^y��r��`��e�<8Ӊ�
"_3�c?� p��y���[b1���,��%���[��=���&�}���}9p��(z�_��߃��gE�c�Ї���v=�1�>��W�$�(}I��a��`����1�VU����v�`Pv5�0%��Ƚ��W�v)��6��nT�oٹ�rF�Wf�!�̑����IA#!��m��l����B�^�>������xG���2j�z��.��m�)���a?����.�g�c�ās��7�gA@��6����Ȩ�?8ɛ|Q퉅V�X�R�4c��Y91��k1�nvYkG���Ib��˺����WO�!���JZ�g	��t����ЫTW�pUC��f�����rY�.-U�䃙�Ջ�a����g+$e�$z9l��D�ŋ���9�WY�d����^����~���)e\����\�����O���a�C#�=�A���	�,T)_�QaM@�N5����O��WBŋ�Tc�WR|-f����P�ތ�"����^��>������`�2N]�:����⍌�gۇ��y�xC�VQ�z�[B�:q���H�!���7���'�U&X^d�X(�L8�n�h�cqy�W��G��s�>{\;	́  DcH�I����!�_1�gC�H������k�SNq崹A�i[��9Ȑqo�*/�C�)�B�����t��3J&_gnkFU�>�9�����s
�Y��j���Ɨ�	��O�~�N��Vw�r��u�a�P�	�B5Լ��Ɓ��N>y�	Ul(	�O1�S���/�� �8~`��V��T�Y�nviM�
Soc�cl8��[��BՏ:��(ҵ��A/m~�n$������XZ�kz,��2id)�7����|W���d�p؟!ٕ�es՜�D��0'!�g[8��S�Fs�M�����[瀯F	��}��!�вj�\�fX�3"��3��2x�N���=�1�n��d
�\ٓ�-;v^%��t5�j6_F���W}�[c���]�lJw��x�\�xH���ɔ��V{Z{l�}wgH��J��OsnG�3NE7����z�ps/1���Q�S̓�zm��-�mE{s��{+u7ל&�e[��g�|y��d�]%�L���7�w�����1eyNQ'�y�г�|ԧ�r�ڟ 'vGP�}��Vpt7�m�`�f1�}� �~Nm$�4�tE��x���p�ag�E�T��2�̍�����͜O����y�����XKd!@�^i��v��T�
ygW�����7Y̪�("�
e��.�ߪ�H
�a��w���A�z�̰R�����-,u�/tk����eS, �L�8@��XP��^��c%~کa�D&��&K�Oռ�7�
������LԴo^ �Fcս[����!Qm)ĵȈ��x���<�Є�r�o������4��A{����8S�cX^�U|���{gO"���0�c�N�}�0#آ�=y���(�~,Z!x�F;"s�~�Lc���/k���(�aO�\ᮢ�� f��B`�汤�1��Z�!@���e�Cr�:{��y�a��J.�7E1��C��={@U� ;H��zϩH�NuO9��L��9k�دz�+�I�O���z�Z~d��>]&7��i�7o;ҍ�A�O,o�n��?w��Yᬹؽ=���]uv�w,�W���tmJ�g8�����,xG�㏄�y���c�����H�dj����[\V��E������w�h��ӎ�+%t�:˽�����I7�X��t����*���d�n�ȹ�����o7�S�6�LUs����2�|�|��D��^���"�r(�=.��f1EP�s;�+�c�{��V������|��Dk!�G�8u��&%�T�
eQ�Vr���a�+�0�V�v�FĘ����.��کf�ضf�AC�0��y@����NZ�Y���jh��יlG�CV2v=��Rn����"b�y��p�ʁG��	_o����譠4�����sDO�C�FQ��O�W/�	~1O��#�Ͽ.����x1�C�u����=A#z�O��.#�'�sD<FVB	n���
-��N�O~���[�s�Cg����gDqq�[E��d��D�l�+7iβ��V�!ò�4æ��/M�j63kח��8��@���r��;I��-xpE*ެ��	�R�t9��}����	�� `5��95>�z��i�䩚��A�Sgn���FlUr��ݪO�S,G�=oN�c�9��BËk��?��n��kf	`���l��l焦m,.�G7����x2jY^�]:��ݾ[ռ�vg��w��;�C�KI���{*�̃���y�j��OPɣս����������6t��PBuJw��'N��u�W���]�f�fu͋�q��P"��v���|�a�L���\�R��ǹ��R����np�{.�=��T��oy�����6����HK��7_i�͉Y����g|�s1Gw*��5xtA�=���ĢY(Ъ
7���Ǆ�o��$dV)���ƦAnc��
�.�yF;5)�æ�H�>���ºe2N]�?qR)�y#	���oP��1[7zn�:�O�*��s�C kLa�gn��Y�M��D�R����`c"���a�����.���f�6G^��u���ض��!���߃l�؀�*�r�i�'�Qi���b��o)���OGy
dkH��	���@!�x~zc^�3�UM�G���+~"�?2m�����t�2�H�P�
�礱 ��E번~��B��5���A5*� ��c/�G�3��j�Aڰ���S������)�x*�^طvh�`Γ�a!��;oMR��fˤ;[8������t��B͹��A�ly�=��O����g,���A��du��97�d�ח�e�-V������C�I�]��ުgJN]�Q;	y���,��=�C2�k�GT�S��A�C;>�v\��/6�s �T ݠ���do�������^*��%��v���1s�|�,ʸ��d��.f��e�P�IV�`��c�����������䦔,�K��^X�Nw�W3$z5�qoGrh�x򾚶�#z��7v�䚘�c�kV����޶'e���*�W�zi�IzQ�s�-���h<�9�ڂ�\�;[AYqѲWR�X�:�t�i'\̧�Z�IN�H���i�bc������e���.R��)В7#�De�sVػ�N�4����>O����Ғ�e�J�>���#�Ot�;�Q�V����6�u}eC��X��N:��ЄOE:�וKlN��`q������\n���6rB��Xw�&��[x������F�
ڄ;�b���Gv����k\W,:^}��}�8�׻B>�����]����Sj�45�0$ӛܲ�X�)-L�W"ka�ZA^-Ż�][gql�7Q:O��w�$�oF2#%���Cr^�q����rm7t�j�����8�3NH|m�����k�:J��	o|%e�s0�f�!�h�CKT͂�k��H�u`���tf>噅��±��ʻ�rjq��aM���M�ms�X*����|r
��;�)4ɻP�a��䨹�죃r�S�0W3�#C�����Bi��[7ha�v�ӵ3��x����h�'��̭Ll
LD���,�u�X�Ȗ�$��l���Y�g�ܼ�*!��=��$� $�W�k �W.����Z�x�v��-�B�EFTVӥNX�[nN��#�f;��;GbF;���$����S�6f��+�-�������.���N�3�����p��s��#.��1�6�&LO��ٸ��ۉ�=y�vA�����<����`���t;��#�!�ȳ�#S8tv���_Aw�`���#M���ˍù��h��&*N��e����٫%N�kz88.W�q��9�p�K��u"k,�xyc��}Hl7��cJ�\�J�f)S9)[(3��.�Y�5-��ɕ��i=bg5u�ot͒����j�o�+�Q���L΅�̗�/?��8I;�V�TA48�� �oV�i>n�y�t1��N�[��y�z�X��ǹ�Q�:�n��,�XJX�t=��P��Q����r,<c
�ӱ%G�X��]����P��쵂�y���r.��O�����L�g
�;�0��ᶝtW�b��<v`y�y���em<c!ƚr�"�Z������})�s�����(�q�����ir����o��`�2)T��� *h�GS�����N��3*5�m�k�+\SE����2�S����W�]kv���]`�W/;7�{��؁��"�0���W�(��Q�zoX�eNfE]n�(��J\v��͕,In�Z�^H�&�����
�qI��h3�݆�BV�cR�F��g~j���AF �6c8��D�m':E|B��" r[�l�F�UF���!�L��o���A��b��UDQTS1�PDKAEq��UUݪ�&d��o�����~�����~�_����	"�&��:)��
b�("��b��Z�oL�O^�~�_������~���h��{:*�Z"�����\�I��UEQTU�mU4�`����扨�������-�4W'DmA��͋�9��

���%�Z*���MRLH�LA�1��PUTQW6O��)��*����ISQ5D��T�PU�IMz�T�UTEVڦ�h�����"�����AU�IEQ�6rt�EE�EUU���/Cb��*
��������5EQ>�J��)�"��+�b
����@h��**"((��Q�PEE��f9�����~}}�ۮ��vQ$��/dǋA�W��jz�	�gT��'Zv�t���u�%w�+	C`�`���t��҈3ľm�&\C�^`����G���S��e�~u��z�=�����C`�氥�K��zkNlnϬe��vMwyl^,F��k�UN�i����Ci~c�Q~O8�u����3�"�@{�d^�Uϫۓi��g}��(#��v�2c4=3�!�%pCo�2�)��l���ެ�C�EC�yu�4�����a�;T��"r|7r^m�t���	�8�)l�9��0��4�\iS�j��} �B�N?y�KλH]:ɲ���C-{ϥ2�*�Ia-�rq�g()[/%eο��7�=����-����N�/dp�_JnjЙ'�b%9�����o&���ݼ1��,��
^��a#�-��cz<�<] �D9�a��m�ҩ2���/��L�����uY�KV Ȣ�O�<����	2y#a�y7W��}YX����{������c�%݇�$������뢢�X� �P\^�P���oP����;�\��tr�l���k_F����R�W*םE�P�+��\��/p���������֨�?T-.�����d��*O��,�u��N%C��$���;@ވ)M}fd��Y�kf�G	�/T\#j�Ց�5w]�M_>^xPҐ��
(>̕��+�v��Y$	YgwG�YjT���t��[6l����fo.s.^���^`������������y��+��I㰬e�c,"e�R���k�qvJ���s���~�"}�gL�� ���.���>.���!�!!��������1�zhZ�9��(���eA ����a:��譆j����MvLl��ܷ��0A���i���!ٕ�O0M�g%@�e�X�j���;�NTLƣ{;M��N�5�/~���,T����&����Y�Y;r���[˴�����j�����#N�]��X#�)�f�rb��c]���C�y=����{aX��Q�
�������Cv/v�0�{h��!pz^C��TFhp!V�i��`���(mgdD���/Y�V�H�F#��ݘX�څ~�܌���Za[��{z=x%���3槹t�:b����4�B���:+:M�t(F7��ās\�*�OP��ke���veK2����,�5���6+�a�B����|��sY��c���#�G��l�0��%6�f���2��p�{�.g�r�g:���6����	(�z]��X�����<����6T@HO��x����E����r�o��x�U\�z��d`�nǖ_N���Z�-].�7��?:�����`NWW/�j����C%����G�ZY���(��c;Zmnn�:H@QIF�{��ft��]	}��z*'ws�ؕWЋq�S�0<׹+u��lv���������c���%�f�2�ydIw�U&	�B*��d�>�3���|4��c&�2`$�;�٧��B|�;����2�N�@�(���7D��.tE1(ʗ��.?ʵ<�����f�~4?�K�<��k� Cmp��pa׷����9T��tS[�:���Y�6�Tj���a=\��Uխz��\�-ك����P9���J�4�ċ*z�E�气4�L<���cY7֭~ޏ�[��i^�?լ�d��y@`鱤B�0�P��a�^�YB����}c=0��¥�xb���l���r�3S�8,�^�<���Pp�_�b[NЦO�4��:����-����v:�V�)�A%�^¸W�wϻ�o�>�E���'������^�o_̟c-;UVZ��^Ѷ+�z��Ƨ��O�*��=�	�G�X%h����Fu�4�ohk��X��.�r��xf*�_@�A{=��|��w6���hvx׺�;k;�>�柮DOj�eFh-.��!�3��þ݀�s�f}���>f�ǩz71�Q�%�M��pc���7�H�7O������~x�=	2��o0�۫��^á*77���/j%wt�0z�#>T�-��L�EWA���~�^�;;�/�h�,��J�)�j7�b�|w�]:gI��nC���٦^L��������'eY�N��욇�ˉg��4.9��O6����輾�i��,:�Y^������.c�?j�g�g����g���o�X�ii#�|�No�S�/|�ظ�b���͙��Q��ə�."o�3��-\N�|ش�1�O�E;Ň�a�yp�a3�Sl	Ue"[�l�Ͻ��ʖ	��0�Z`��b�זt�
���z��x/V�΂�r,D����.ue&l�'��I�6Gdt��頜_(�E�(������u���~�j��\���T�6��V�D!,�ٵLs�z$!>��Ͼo_�L&V���*E1H�jn�"a�%�<m�/:�_Dov���p;�B��<�+%�D?��f}�;'z�$�&\/S1X�"�6^���c�v�����X��[^�==^x�F0C�y�xm36Ƚ�<���.��YC�4����&�W�����ǼA����<�4�K�����`8�v���T ��o'}�)�t�"��#Vo����] �C��A>;��Kûs�;���݋q6�F3i١�Z\�ڝ}U)��RZĳ9��4¦q�p��!#��+c�+�=ؐ��W���f��c��F���El�E�*��(����,�V&��Q�U�\�jư]�	����S�mg[O$�s�mp��l�����y"v�tZ.D��_�����ҋ��7ܖ��'����_�6|�;�\��߅9��x)O�����X��.����}a�0�}xCb�me�z,(�@C��/B_[$z��Z�2Xu1�e�ˣ��zM0,���A�����c�y�Z61�L#���Ƀ)���v-��%�>^��Δ�e�L)��b��kj��'I�ȻW�}��W�g�֝4��.xG3���
߮`&KvC���hP�]�	�ZV��{R�\���0]���l�`C�C`���a'�f��7�Ӭ�.�m��[�M�Fm��s5R��]棱��Ri��O��Zz�x5��v�
�"�@{�d^�y<��l�U�|y̷�E����;6ӹ�1jK$��$d5�S.qL������:�&�[�-�ouq]�������L�xw&,�Y���mAЗkH=qQ/��y������7��7Y�uܗ�m��?2�U���J�F�Q�s�e�(ρ�&��Co'UQ�,=]<�s�*:���"���9�Rad�
�+V�iIp��H��X1Lݭ/�켧n�WUP�:�ְ������7�,�j�S_mU���!6ۦw�(2�Hk�Mۙ]�]�T��w/+7���`p��8�=�%=�ԉ�xv�U�%]fқ$rP�=O���P�uچ�{�q��ݏ���׳�5�߯��g�L��If˳W'Q�[��s�|��n[���+�`$�L�W �؝Q��i�fw��t��L��m�Ms-$i��q�������p���7V�;&&��7_xs�ac/��/��7�V�uFJ�5J�51a�y�ONe0�
��/'�-b��1��0w.g�al/H��=^�*�+�iR4
���\��·�U�����*��1�
�t�TG)K�υ���ܸ�c�2�d֦��Adb�{���YL&����@pTϣ�H�4�97'�e��Ǧ�!�A8P�[�r�n�y�Fs�^�L��Bg��q���UU�*�HVSk��kE7"w�6�"�ӽ��A���a����y����_P��t�S�"�?@[[������}ePFI#�0} �g�v睩ގk�7�+j�O8�x;�Lz)!�������xq$O�tTk������\k\L�b���*U��٦�Ȓ*�,i�Z�Y��8!��r��fˈ�
p�/�wO[���NxA�A��:j)��s��D��p���&��d_��8(j�Z�4!G�Q�ؾ�pwj��4V9�z��p���4��&�O*S�$x�}�_������o30��܅ͫ	p��cj�^n��"'�ge"t�i��u���&���Moܺ�׮ƍ�
�=ܚ1�Y+Q]gPJ��F�������D��k�wm[�SsOӲ�T��0����'�*�y�ݥC�C�����Gv��SH�ɠ �I۹��2[ o}kn�Y�$]X���B3��Y�e�@nkk����I�S���F�(i�@�.Dg\��(ssX�"��Co@��+F����)tyl���?WK]:����WL����c�l��к��q:{k�F�Zh��:fF1����m�z�1G�3��&,x���iٽ�5�)��ם4u$OD�h�?�G��2JM{�B+����~9U�6�
��,�y�H���g,�$䃋�~�^<F�Jgk>�n�=]�����PXS��B���z�1H3�)*η��6d��(Z�$&}�ؼ4������:�ɰ&a��{]�!�21|�b�t��;�t��U�ζn�9r@�^uj�P���I��P0����{4��^���r�nt�oQ�ܺ�b�5)��nS{�I[	���Xu�v6�<�]�;���s�⊂J!>�������˟��}���>|�'�c�S�ȹI�w�X7$�8�T)�>F��t۱����'z��{Ga�*,��Џt���c���Y�_7��C��ߖ`�m�a�}�C�f�R������e>ϵ~�9�o��L��Ɏ��t3Ct�4yÓ�e�iV�@��$ά�bs�iR��t*��z�ޕ����Lh�������������>��8"�E����{5<#sQ�;��6�D۫�˞�S��ވ_sG��m�t[��g�a�2�D��_dwZ:6_��mgv��6Z�o@>;��&Ѥ��m,޷]B��XF�nCS�c0�6s�u��
w�YC�
U���̟\ә��AQ��H�=�Eʞ�gq<�u������y�5�;V
��)N�0��j�MՑ0��Ö�jܖ�}M��I�J}z8@�=:����Q��T��9ig�t�r��iQ�:���C�a����u�w�zߖ�}�IVxk;�F'Of�yY�,V�΢�}�\}�%*n��m%W'�="H�6@N]a��������6��(cܺSwC5��b�n�|"0���aٛҢcs��a:V3To^�{���]�\A��E�?��W�љ��@^�>_=����������ȡ��������|P��tZ�nsǷ�%|�hz2�&�+����� �.��-��6� �Ð�c����"�7)귙3�C+e���v��Fa����Zgl,�n��Ak�`d����[2�>@�N�͛��i����H�{�wJ�~/u�Z��Neԟ7���oT��ֺ�������y04�����%"��EzJ�S� [{Y��o{��2�V>�WN�HH��]>����J���<�}�}�v�;#;"���P�M��~�A���o�X=u�נ,�ӗ�0\BH���-TTV���$�~�9����y�W�����@�\3��@%Ctlz��ǒĘő�6�GB5�y��
ڰEkr�� �=Q�3�΁��|Ε<�&����ٳ�T0v��v�o"@�$aDl��[j�a9>�ްa
9D]ۊz��K���MѺ�8J���:+�F'�hʎ��	Ђ�z����e�M��:���j�s>��C�g|����J�k�	��{�c`��#�ٙv�.+�0���#�Gs� ���5�]�*�o�
��-�������ׯ�>��o�&rEDAR5��Z4�P�	Ƴ��&iU^�,(wa�+"B\ Uґ��O�[���=������qcW�C��\�P�D�T2b縭�vg��R�b�ڃN�qM§����g#N4�Je�\X� ;����d���B�� ْ�=3�)��ܻ<�&��@̓4�4���2��
ո�R[Z���ai5W�d������ 9�U��S��u>�ȑn� A
=Z8t�Y�]�j��X������c�$�B+z}>���z�����uF�F嘾hf�9s�á���BM�ް�t�Z�q�ڟޟ~�[=��bIBB�f��=_�����0-���=B�*�+�}J�������fڬkD�#!��Y�g���y��O�J�q2,��w.Uk��J��UaD�24[f�殷y��&��,ؘ?��a��.�T�+�+C�rr�
�7������_�tކ�Y)� ��^���jUS�hbʳn�s�a�ψ�z�t	��5�3�|���9G�R>G݅�:Y�W�D&m�D�1��R|b��Q�t�֙:9O��:
Wѐ��.�wXN�VtS�}���:���v�.(=��O�J���N����ҳ/1XG�N�X�����s�c���A�0nB� ������;��F�Ꝺ���	j��e=���b��R&�?�/��tޓtm.�mGƜ���H~�.��e�=y�\�b螛� b�WQ"�;�Q �ʚ�>��&�e%5����uWuq0�8Dع
�D����h��1[�.g͝u�qgy��{W���u	��6�H�Ũ�.��e�Y6P�z-Gj<�����V_%���C�n[_ct�iP5*��3N]�+��RL)�^ո�k�Ys��n\�2�u��'2��H cG�ݠ!GT�/�=AN�Y1��8b�|w��B|�!�S��/�Q�q��0(Jz8(�����S�R��+;tb�Z��ź��N+yʛ}�\��N��__s��A̼$˽&ؖVN�� K��{j�'\u�GgK#�u�W�U�����YQ��*S�ںKF�l����Lۿ:�j��"+B���V�ǘNaY0���4��@��h�{Zݣ�q�#_E_Kr�S�"�.����R.�S�D�@u��&�Z�%�ٖ�Ѧ���x�6���e�'1�a����}�A6���m,�s0�E�UD*W���r�����Gx�$x-���A�d=V��uI��N���B/�V:�힌j#)*��\6�'��m�5k˫F�����oj�atF�jʝ����Qdtgrv��ޒ��ɲ�$;���×���16��ħ��t^mvov�\�����0�D���vs����@�9;�i�wP��cc�ok��P�&��.ZǴAy)\x�S�f�:f�g��ت[��fm�,�d�9���`�����ŭ�+-ċ+�b���/n��V��n5��X �B�Y��.��2��6a������#lWR�r�V����rA��cV���`�h�ۢ��F�M�c����5��.��j�|q���&\�@lU���]u�k�|9	c��� �'I�.hx�����[]�r}�|;��2k�X1��/��fK���GW+�a�3��f��˽�����}��)S5�.�^��T4�C�Mjӛ�k��n�N���"v2p��b]���a�v��Ƀ�с�飯��j�V�}�1P�k<z�b�TŚ�'�l��cA����b��9m^�yp�ܺR�X����#��<]C����s���\�69rocU9�k�	��[�}����d�/� V�grF')���y��q�;'�Z\�T۴��W8��c�U�Y����Bn�/+��IIB�;� ��)��(� ��gQ{�Q@U-~g><~��o_��������~�_�S�EU�4]���1_,T�MC�lꃐws����}>>�o^�_������~�_�S�EI@U#��Q�J�*������*����)���%�`�jj"�� �����F�*�J�4j�NA�)�A���j�J"#�5�Z���*�*�JNlL5T�se��������R$�@i��_�1E% �2Q\�T4QP��b���*���r"���(����AQK�u�7��S�R�4��:i) ��y���%𖆨�����)(�����;�� t�vf*���0�̅��D�Q ��/��w{��u�!u�8�kY��J�*[���U#g�*�#��l9�@8y9��*��@z-���|!�G<m���o7�<���^gj�aD��ݪ?�]�6z������d7�8�p�&����t�gs3����B��ۓu�.}�=�	�� !�|�4?���P�� �c]cjm}����F���J�A#����+�5��5�΁5��[��-�w=A�=x����f��yo{��"F��h��{dv��+�T��i�{Y�_��թ�68$ӧcj�so4OY�F�N�M�.���yY����Y�r�Hا���!PA(w&����ȩQ\v<���<f�ص�{�(9Q�~��5g�~<t~p��)�#��,��d��.2���cT��Zf�ùLD�ѭ�+��r�
��.õP �.�i�5ؘme$Dd$���i�,�ؘ���^�=#��	ƨ]^�R�ESeU�2q,�ăF��c��s#s�ۧ�đ�Z4@��	.�xF��zx�~�b�����۽�߽� S{��.>���K[+FS�?O(=�xoY�G�W�f9L�:��TΠ���f	�*尊������7���{�@�`�[��G��I�i��jq'��B.�3t7W�WR@#r�:��[��w���&p9-�-�,)K,��\�'+D���������-T��8�P���5s��T'��<��*�X�F|���m+�L�n�����l�����/�=�|B����/zM)��V�����WT�,n�b������xS�D����W;�v�`��!�g�aʘ�MaYR)��⪶�O6��ЦoC��^G�k�a�҆�����p���\\R�ߪ���H|9���-U�V�D�r��#);{wԇ!��m��͉ȓ�Sv��i@[Z����g�خ���{A��ҙ����Oʠ<h��Nrbnzpc$WC��wX�}�zMׯК��T��:�}�OA�9��g��5��>����G�²��ؽ���H�$I �T�%����f�cz������R�X���"��%�*����d9'kT���/�w6)�go�k���#�l����s9,��D �E#g����NRw?1)#'�k�Z�:���,��KK|w K�@R�-��u��q9��9���O���n��{]ݍ�d�B�X��o����҃��7��:[�W/knn!�Z��O�A���Z�h[ ���;Y.sb��mf���2a���g��R#3�^o7��_nK1���3nNލ��6����ڛ�Q�@�XG&0����n�e:���
�]7��##d"BCo�HJ߰��@�d�sNdPYd,�:��g�l�1f(D�B0ۡ��>U�;��-�*F�R�P�g�w3lT\ƴ��Ɠ;��DqՏ�^3�.���*E���t�t�s��Q���>O:�SFo*Z�q|7���G�n��jx�:B���i��������]���^��'��y`��?z�Gv���Fc���N0�B���p+`��n�Mr!�&H�isټ�ՈءƗ+e�-kd��*{����` �ov5�W�b�otu&}�'�qgh^�z��Ǐ��i��R�x��6Z�P��4oN����E��0~/��E��n��qSKw������a����O����_s��gx�� ���r�ہXiS�����9�uӌ�jA�,��ޚʖۏ5p�a�Ѿ�A^�sf��E���UfL5ԋ�jmGSD�4���U�ܝ�X�	���)+&�����x�9�6�v�����^��}�RS'k�n��Lڶ�&�00��R�x�;2>�n���y��k�����_.�>�"(�ڐVPk��B<��@~�k�V��亼��滪|U7fTuk������gM�PK�����\3���-�ȕ�k�5آ�6'�3�޷��O4g�Lc!��l3����*�ߡ��@�f�M���dn7�^Y���AK�HG����t\�{CH0�ƾ��ܸ��b��hVY�)�&�kj�}q�ć?�݄t�+"|��UҝV����B�h���3譔lI3װ�H�(=T����u{*/S%���A6��]�7�[l�S[>�q���:�W�<<�L��qb~���d���B�Eg�9w���3ѧ�}ٗ����Y&;UW�gٔ:���i����؄�[�i��h�!�;��oTp��C��Fi�U���S�ܷSِ$[���
j坆^�m���V�t<�Z��C���].b�Lg��#cl5S��t̭���yvwPJ���TM�z�9F��$�wskb�r���(T�p�]�#�]p��iv�����N�{�l'�癵�
]�c�{�K�W|��r�Z<0���V_Rk6�M�5�եY���ogt�.�uR�dص������5��)ínN�q9y�2'�����:1,g��A�z�ǫ����\m�km�{}]A��T�]�]w��k�L�.�3��竬DVr[����#Ew_��[����V]\������"5��`����G�,�0��ܭU��0����jl�̬���W�e�{�����~2����Ͱ�]�D	��oM*�`>!P-�5����w5+�f�bP�)Vzz�������������G��b�8U���4m�m���Arb��Zy*�n}^]9�ٺl�s��g���Gd?lP�'���Pu��KԜ�^.����U�2d��>&#ðWN�x-���F�@�_V�ꮫd�u*����ѱyo��}đ<K4x�5�d��z��a]�;^�l���:=�&%X����3v/	=gd#dh����=���=Vgn���/uِb�]��tx���Fe*���mG��+Dn�n5ћ�y����"Nբ�ɵ)�R�~�(,��\M���$�4�bVK���43���2ΥmMe�JFJ���$f-O*�դ[=�Gc�����u-�&�y�b5��ھ9�Í�:p_�Hp�p].CpG�T����Fr6�A����ٻ[�p���vfV������pht��)���Rd.�O2,�ޙl����Xj�b�IљCy%^X�:�÷�4�}V��,���O!����!���ogKLsC�|>�mp���!Xj�hq��U���ql<��X�&�/Z�u�ڪ,�W�!j�C�A�Eoޔ�ޱ���)E�t�;�S�tN4�����։��;ݶ�}L�Q�)mKp5�WYx�͞K���n���S���=\�d��X1�����M�Ԃ���-�ޓ^�����m��;9�����n��ۺHiJW��3��`0��ycp�o;�1��L�9�.��ʼ~P�ݎG�Q�w�	�ߟ��5�����m ���LĎf������X�w�8���ޕ���!0&�M���R}��q�.����A�w��1aܸ¤@ۊ�^��X�\���jh�;"�Cj���;B^c��Z�2Q�&SH)jR��Q�[=����8�ˡBϷj:���4�7���f�S�����*�k$��IȽ2Ԩ,�����':���op�ҧh,�v�'�΀��$�n|0�1o��{�z4���lS��^t�yY����~i"�a4?O���>S�}�9�OQ�gh��x�^'Vd@7��oQ�z3�m����t6|�_��|�݋�=1�~@��?�j���
�E�#0d^�D�H�����[!�W~yrl�(z����o�7���B��J�rh^�1��8e���0�4����J���-��lS�-c�	'�U#U;q��7q{�G3���P�ֆ�6� �֜�W,���^篔κ׋��4��c?A��E���^�0w ����\t�wx�dzn��ƴ4�#sd��ik��`��}��vz:��CW'��Q(�^�3ё{�Av��~���*:����Ԋ�Sp��������xD�qf�{��Q�w�_�g�\�����]:���o`�Sϸ)�T�k�c[%�f�[Wd�5��G���מ㫻Ǭ�fD3c�@lAY�c�P���dg�D3+�G��c�H7�'�]�u�dTQ�5�uvx<=��:��)�W�6��g��~Q��������]f�]�9Kl�K�Jlە���ܖ����+0�H��o�58\�R��r�m��Θ����Ѷޣ@���w��9>����6$������Ym��	;U���nEE^���c�,�d��=��Xa�j�h���'ti�gٷ��O��z�/�υrע���R�x.�mx��*"%e�آ��s����F�U��;��R��(�c�魾��4�D��ct���0~����C����a���z�Y˺NI�n�	����v��=U��vP����a�;��;Qp�q_丳�	�/b��Z���Y�x�;Б(>I1��^F�,���gU��䕾�q�gh�eUZ����&���:�H퍜�(�c�O{��d3������gn��B��=t�Uߠ����������҄�}(��,?cz���.;�3�Eձd�lVq�W���L.�ɚ�̬�$uvM�D��Y����d��Z�\N�V#���ӕm.���lP)���D��&-rY���mG�����O�GGo��z>����b+����戋H�O����{�7�f���|�uDd�N^��}30Ѯ�M�t~^�f�{�쓼��B�+���cA	�I��LB��+hE�.ۀR�-�x6�Q��tH��t*������^'Ye���Ru�x���m�%>���uZ|�w��ڹ���TK��g!]�4�в�+��Wz.��t�tE��w-�����s�Gݹ<��t�d�҆V�� �yA�K<ռ)���⵮T�|�Z�d���^d���|�;��{2$[��-�+k|c�/�M�],�i�D{/c68�t�[t�+���2�<u�Ƴ���i*6o3�{}�2���}�m�P���z�J�R��7.���d��!��e���1�隆�pb\pKg�Gt�=\O��®�Y\�J��Wu��홧"EQ�<zm�6�k��kdy�p�-��[��`�+���sULM'�8�m���7��Pg
�o0�xa������
��X/M)-8�m����fڥ�\���i5�������l�=�~�ݾ��F�8�E�J8׼���,V�l-�����@vqD-2��~����`�6�p-��5I7c!��{�h�V�����r�WN�!n�ogɉ�<ifZڭ:�/�3�Uj8K�ֹ���Uެ;�`��wYss��J�<b-�a�Ɯ�	f�+�3�,gRG+A�����ٻ��FwqI��^�p>�9S�q�.��g�7�'O߾���"�E_ib��ƥB۱v-��$x��#���;t��M���(���[���h܍f2'A,�R�7�wF����p�D�KnI�fV&Bj���QǗɴ�#�1Cղ�ں�/7b�f��~Q������?o�� �2�����]#���8���2R���f���*bk+e�#U'(�-]��SH.����]�"���ә�gS��0����|K4Й���O�f���!�o��%K��'�"��c�\���Y_�&ʨ������#��Js�;����:
uB���ESeU��Pa�M���u�����1��p"+x�t�H��6����)��.�"�����{y��:�����:���%<z�.�,#��9R*�l�>�ѵZ15���Qy����6��A�pX�����o�`�����5�5g�^Z��m�V���+����$���k�dnng#��y|Փ�5���"vaKH�$�̜��Z�;��X_j��b�%9.H�땹y)l���j��`^��k��w2�w�T��*�����+���a�SL�O�����h�|�a�hJk*֚�]or|:E�_��)�,��Ҵ�W��)H����l΁���!Nlũ�Y	0����T�]<J���q��H�8Wj�Qu�8�Dc%��r��e��[�9����+��X�y0�t������NyB�2��%^bwe�:)���c�A�
�rwǫ��'%[6��d�X�c��[F���04H�Q_=���۩�.���z��<�36�2�t����p�Ĳ,Oes=+$ӹ��eݠŬ�Z71�(�u��V���ܒ����3U�'�C�C�
�ʾ����5�2�ݽ�N�ݵ׭ٷ�Y�����mT,��p�13\I3e ��[o�2e�x�lG(������|�Z�<7fs.���Y���u������Me��S�B�l=b9�%�tc�k���']�E\T*�/X�+(
�Z���:�P�
\�͞u��C|d5�[�q�a���m�{9�����ɤӐ��C�s��e�����J�Ǽ1�곝�)�gw�/���PK�]^������a��U��,`E'Q�>�Np1:oSi�r'r]n��sڻ0�:�^�����
#xm��*1.���9�M��u��Z�R���D�u��^i���w��`va������]:��:��i���i�t�rj��3���'7Wk|t�{b�Ww���^֝$r�yl;�+���@.ۃ{.� *L_^^'nSF�-3u���2��:�����;-�C��s>*%��E�vh�B�k�R��s�`wtK����bw	W+z뱙���9}���u�����U�l�*�mPyJV�� t�h�j�u��l���.$c��Yz	c��0!����lD\�Lz�u���X f=�1���p�f��y��2��J�ֲA6ȱs��@'{V����i㿇'IY���VD۰[�Y�%��4C��%rkl�Ю�A��k;A��[MP)�U~{��:�9WE���sZ��\Q�y�^�Va�h��U�����=R���Ox�יҮWL}-��ys���}X9������߮�.G.��V/ �);a��t���Y*�N�-�Wh�\VpW�ca�̆kI�������S�n���@�h�Q����
��zb��iʜ�x�6���/m]�;b��'f#};���`�܉i�Ww%�AW���)�x[�+��yg=�O�+���7:�a`��5���he�ݞ�����+i�:u�N��+e>9�%��^oQ����Y��聶w�C����ǝqW+N��6&3N�%N�銫_]�v��n8]�r�v���5�p.�Q5���D�����m�_ n�ε�0��>�V�uu�or��:6/�����l�]B͐�[uf�0�3V.�t�?4ۦCL�#@� �CD�;u�u��������s�Ĭ����*��o2bI"�h+lQIO�ئ"��J��C��=g?O��������}���~?��=N�KHT�MW툪��"H��A�ET��b���$*�q�����������~?��ǯ��N�HD_��R�͐�����2D}�G�i���b�kI�
*��ʍ�'T��%�Ym�m�Ӫ����Pj��%T�5MM�b�
))9�-Py��AM��klf��(C����ѡ妈��|�y�������Ӣ�X�Y��Չ�bA\��*S��*(��<�O���5O�r8Z�U�Mihז�ZZ��8N����i�Z
5H�����,()��F���*�农'!�B�TEZL�S��8@d�����z$�)��yS;q:z�kv�iWp�CK!W|�p��o�� bg�Շj��8HB�o��A��t�5�]t�a�K�P����O���=�4ם�����vf��ե_"d./n���m��0X�6��SuT[3��L#st6l�C����䒋�0��&�JL-�g������;�x����A~:�k "O�g[v_�rW^(��
��n@�aj#|�Sri��Q�z�b�xhs�g��,�P�q��[���֕9D�x�
웶va�ެQt��}=T��CT&Z9y����3U����#-�v.���p�;�>NmuV��i�΅�+�Pg�g��gTtE��*Y�>�<��K�y�+��$�x���p��v��JO0��[��]^�'��͹��O�Y)2�8֐'��syqV�.n"��<����{�>S%D��¦�۫;<s��3*r�{p��>�Cd�F�:ӛjE�(��u��2ݽr֧;�:��@T�^ǃ����^���<B�PR�H�*=��K���[�b����ˌ�&��ݒ�t�­����c���Xx���L6����Gy�����.N��\�"5>�ݴ+W
3�ɢ��{A�vi�0<6��u�L�9�2�<v���<��©�f;��v�]���k[�9��i��y��h��?q��W��SBȅ���u���U�T��'�qӑ�!�*�xY��T����s5l�cT!z8`�]:������~ڋ�?\����{NA*���}��u�`��H@0����:�1��"����q\ʚ	��3�{��xּ���Ǩ��Ѷ�A�Z!�5+Ƨ9,�C�쁦r6�[j*(r�+�-�Z֌new7g�|��YԞ�̵�֓�]������g���h�}R0Wwyv<x�S.��-^x"��h�ݽú��)����)�4�S�]WrR-�: �)�y'���V�gm�k��d�!t��y��7�$n#�r#*�xW7��8(��z���LuF��5nP�h6�|�t7d��U�*�=}�$<m�[5�c�{,�ܕU��v�0sh�Pc��<h�s����`f_ߗ�oc�K$�y]`S}ث��A��2o"��m?���",�⽁����Csxҽ��̧"����xn�lX�̊�V����������K�Z���T��pԗc��폒#K4�bV$Y��s��qU�lM^U��4;yy����q��c_�ڃ�辵:c�o6��@:Z�L�a���$��L�1���̇ho�bd�%��LO����ܶ�t[�j3J�֤{6���D�X{��5u^̸X��� �J�K��sn�LL�Y:"�0��*ܟP�g��ꧤxD�x��+R��g�׸��f��ơ{X�^���~�Rݮ#�=���vn=M�"aH�΂� �w����&���/0-DK�I�j����j���(��M�;UP�ٓ�OL-�%:�����S`�-�lؘ�q����N�9����xR��Lx�y�ԍ�u٘���Q<f'�k��!��a!l
�ـ3a#̒I�L�W�l�so�c��MR�#�(d9=1�`
�;�o�렬�+���@��}Nk<��X��ϝ]�
�Z6�g�ƻS�B[.�t�B��q��Jz��T��p�z�����#�sAf�w�Ε�:���<�[���$�%�U����R��~Rw��u[v�ᭃ�$���+�}to�E�X�ݑ���P!��X��Ij��O�;T��gR���̋z7����2ѱEu��
���C�W�[ߏ����{���1G�+7�a�vO�=��T ����߲�{ƻӷ`���qo~����$ͮ��]������K��`�#/�,5�\�ܣ�&�mL��+�B�����g`��fry�}�s�t�:���MѾa�,z�k�Y�3�
}���OW���QgD��U��ѓ9�6GA�h1��7��*�m�����aD���ۓ61��R����b���$�:���v
��捻���xj:uS��.vo���*5�F�F��עw\�Z1�W��r�y��.����E�A<�f��W]y�y�G�����M%��c��9�o�v��@q4�yj@�E>�P���	���hL��D���f�f���ʝ�=k���A�+�)v4�Z��66YЪ�;!�ܙ�t�ɮj���5c+�&�Ɍ��o�T�J��A۹4�i�@�<���b٥T\;�������$��
�M]K�dyV6;���?_�1\���*��M��j�&�������}1[P���9��[۸@���1��^Լ�E�#��;A��l��ۻ�T��,^N��Sf�6��뾖)�v��[��Ȥ��e%�>�+T�Jp�������bd5
���|��	�]̂�P��ĥP��7���qq]�)N�5p��*��+��"�W =gO��+x*��L���旆���"��4��_1��U5���x�gL�&����d#iQ(�����4��(�-{�}�5cL��w�Q��ɶ� ���Zj�ނkT�=�-3CpK�f�/V^<�Q�a"W��z;[a��'`͑�^#��fl¡��
�g�����0���r�qE�sϸ�ɵ�i�����nNk�N�Y�Uf_+�,:�H�f#u��ݮ�o�1�T�pf.r�鬑a@g��\#��s�D~ T�qY���.��[�^����m�eR�9�-��i�ꨎ�0*I���9�E��z��/����=W�^��+)�ˬ�Q0�2?Ma��g��.���3볏q`�΄�<e�if�8�Da���z�t�9V����ض�v_��x�o��WJ9�WgS�5Ȍ����U���nε�/K�HDL����
���u�Ge��%�I�8:�2�3ySmgQ��.ݻ�h�ŴDf:MS%]�/���ֹPt�Z�ʪ�̋�i���{.�K�sS��⥼
N��
22)���;�+��A4q��{����v�{z?��`�\���I���nc�YK^\�KX��кiZ��]=	ވ3��Vu���Q�܀J�>�>@�Yf�H�Nm��d^c�f�˰�n��5�oa��.��l��l�����,����<N�-��B�_��\�D�mU�O�(p��`г #�"�l�k�Ur�w�8SS�9긻�W٦#6{k$���[ۗs���[@3��ԈEH��7xH�D��g��[O��{a���M�M_�TB⪟n:�ԍ. ��!�,��SU:�2��Z�e�P��n23Is.8Ѥq��@�21�m�A���Gp7z�"���~<�᧞ͧ�1�~����_*\�2���Gl��n�`�{W۷v:����r�`�|š��9����[�zz���rך)�U�������.�<�����
��XԽ�0��f� {��]c����ΛN�[�(�f�A�E��IhC���6�RVTIv��̸oi-�]X���.�QFc�֬�!k��&.P�ٝ��:��͗�z6/#=�^o7�?+t�d$��}g��7�|Y��F����]Wr�Էz:�u����%�Oj]����z|�C6��pQ�۬2�?q�,���uY���+���zux�SL��2}�`o�����F�3,��U.����}Mu����q�d�}�H��&8��`s�4s`NTV�˧X:*�{��K�7��0��>��׷F���#Lt���i��g���q!#{O��M�nz�
Ջ���2�H�gE��H�$IDA�x嶮���e�;Y�ٗ�(^��-cݥBf��f\v:������4�|�Q1ۯ���ݔ�t�
�ϺYŃ��f	5�[ţ�1u'���f9ob{�^��|�W��E%����z' TK�{56HW X�ߣ�w�y4�-���M[����\��w'$ِ�:��w3�^��8�(7��h�+��L�La��@����p�	f�H��rr�B�Z�M˗��o$��u��@�A���|�b��-..^T�u�w]������$(r�Hs+M�]zn䱳n���f�W8_)=���	���N�8U�i$g߾?��������^� V���E+�R� 51�$�o��p K�ۏ=��nue��!G^m��W�# 3D &������$��L��Cl��Z�n�EuS����h�v}�x��HU�2<��#k_�;u������M��l��S#�Z�wꭧ������	d���t��_%UesӴ<γ�ӣF�j��ۺ=���Iۻ 0�,������TG��V�c�HOUq++kCi�}���ww�Rq�d���&�����Fl0����Ϳk�*h3�X3��5����lG,G����AWA�#������S�R�;��VEg?v˨��@q���zo�3������#�ڠ���Pe��n������O�AP:��#b� hd�#�|LT�VMkU	���}��Z��E�eO��C� �G�dG�¢�h��}a-��z�8#޹�u|��_:���{��&c���=�������n�3[G��;�%܇-&g��{90$>P+t�B5,/32�|.���st��i�:U@�����i�ЮW�δ����8]35������y3��E\�0�J�u���짜�����{f���)�a�߾?��1��x�t�>a��!{�4{tT�EA�3��y�Z��{�;��������󱬞�:�w�}:�/d?��i��=�6�wG�J�H��,J眿�m�^�Iƌנ3y-�!����2G	�oY��s�ԅ��5p�b�@Z=-�9�={�<Y>.��^Ɉ�,)6dЃض���[�YeM{-�z�5�5��h�b������M��� �oB�����Q��$`�|�]�=G_]��S�h
�B��W+x�t���j��6���G\�N���7O`k�S���t�rx(�
:�ژ��ضbvZ�����KҶ璀��^��t�y�lx3Sv��n�m���/nD�0�Ĳ���o�A�N��WT�-W��0\��kޓ��������_�N�>x��9w3n,��Ȍ�ت7��oQ���vM��L��KR�v�B���J����t��M��djR��!n9�[7e�Y�sd����~^�pۇ}�G^��ӯ�
um��5WQ�:Zĵv���K���%mEA�xr}F@z�fbGť��no]Áw�Xu�z��#K�v�+��n���6���n��O��������
�~��cO�2!�͟Db}�a�k�y-�Q5�1y�}�`�����3No%=��h����R����P~[>n�u�Nt����F�;�*[���O;Om���L�9��[l؀�+�2�QÀSh0���5��T/a���v�����~�XF��^� �k��Y$Y���,^ͨ�ȉ$:�b\�ٗ������]�ٶ�g�tc�6;5����<���童3Q���r-7+_�P���{{k�7GU�`���c��VhL�T7��B|:���6�y#�9��(/h�P�Ί��ݪ�~��JJ��	m�\b�︠�+��2�SNo�Ov]�w>fk�ouZ^9�>��`���*�B:�谻T�p�(l Usm�n�̪{9�MK87\�M�vMA���N���	�H�T������!�����y��P�t��U�т�}��m�#hS��������Zky���r[p����xn��<E�;���h�P�N�44R�7�.�5�N�kW�}w��9��{ytA��V`���z��X	���=��D����cx�QΣ�;��k9OE+�.j`�ۡ��a���E�T��C����y�����4`{�7��yf�7��S#�Ɠ��-]�ظ�7��R�kb-�r���f�ܳt]
��qĎ�e�$[oR�dl��ln����op�o�ծ��i_L�$�݇Y&���;����N�h^4���T���/�:U�w2�ћ���~����.����P��ߘ��M�]����%���;'s+��ٲ�/iI�D���+�u��:]��j�_�1$�hl�Y�B���{4�.��ee<���FLK'0�����2���E�8-����c��k6��v;�L�3�d����f�.��qT�7JwHu��2�h(�cRd�
�dԃ��jmm��~����˽���"Y�B˳>n���1��BG3A�F��X���ιK���}�_��^����6��(��D�+��/Mq����N�>pGP`3R7GFL\���̩�.=L!#�I;"�q�[���6ay��lMKF���{�e�"�A-�ܺ�K0ȝ�4T�mrI�9v+�V�-_, h����!�d�*� /"}�B�H�t;��3mc�ܬ��ރT�Mojr _==j]Ÿ���ŽZ�R҅�d�՘��K`�[�h�W�����D:{g�5���\��ז�s��	�ɱ����J[X�UîaZ�hf�p��Ax�l���H�����3*鸴�#9��pU�qw�����]2v �W��ˤn�p�'ga
晏������%�W�X�WMΖ�0g_V��]y	9����0w����������^�����p��z�5mZ
�S�x5��,��Y�ln�9�6�̰�)QX53�ikL��Xr��K.4�����Ҁ��o��3+]��T�|�Μ��eJ��^M�Sy��p�	�Õ�n<���Xk;$x���f�p��h�t9A����Vt����h��]��7�U)ΐ.2;�ͻ�禃�rKIu6�А�����L[���,^��#��i�;��U'�J[^�O��g��F�F����E��°��S�j��x��%�%��#�u^� �h��C�2�ʼP��H�	#��̝Xn���޼�k�s��oo�$c�ۍ����Wu�7� ��4������r�$�,V�8����'�3��E��4͡��
5x�C��r�ڬԺt:���Pev㝮�P��X�l��oӥXh�ꃦ)P�8x��W�4B6�\�/COn��`��:κX��3I�7By��{�"�����˧�sјZ�嫱��J�n�����χ��o=^��硪}IE4:�AU�k��@P4QDDIN�8b�l�>ߏ�������~?o����z�)*�����P=ى�%�Z<$-D��g?�O�������~?o�����?A�"5ZM��G6q-��lj�M%D[8��~�"�ݎU�Mkh4~��p�bJ�mVCF�[�E�Dқf�:t�����v���h6ז����4:M�fƶ΂��F-4��l�l��4'�d�E�%�8��ľl��4i��{ۙu�N�[�i9W65���Ωy��"��r=�s���Q�gF�Ui4�����m�����z��"�-�V�b�A���5�bד˔ع�\���y��"\Tm�s\���5�4Z�ĻZ�4�l��m�Ɗ1^G�TW�1cX(����Pj�F֍kcF�TF�F�ۘ��j�UcT�.m�*4V��p���,F�PQ��I�2���Vm:|�C��\O��$J �j�,W~�賰�4 ��\N��XŅ[P��=Q)����&`����<��oF���������:�<��EU>�{���W(
�>���Y�]������_C�q�aj��7��c�q�y�㫨����c���V��?	�O>�t;L�n�`$�ȍ��^�3(�L���ʗ+e�kZ}���!h�g<��c���.vs��xn� ������rבE#Wq�Q鬫�{��o*����U��w�e��;�5אΆ��x>��1���sNw%�9�j��{��j$���T�S�,(g��8�oC����
�K-�m��=�S|,f#�o*A�7+�#����;9C'h6�������gFr\FQ[:Ѵt.�l,k�lf���_wԯ�R;d ���:���O�r��ݎH����,@l�0���֧Lv�i�y�,8\���2�S;�Lu�0���ɷ�n�{LbB���:։F�ח�>�$H{_��94�şm�W3��/�}ױv��
b,FGCň16�ё��9j;t��{���Vk���zm[Y���j��t;�ǯqǰ]g���5�>�v"d�G�[;�P�w5�ct0���Aʘ����X�|:��o��rZ<i�oq��Zټ���vv�/7�ۻ7�	Pp���E�p�aDy
1�F�3WU�ˀ��݄�M�����&��wY�7l@@_p�W[��q����ԯߏ�E=�C�.Y��>x����K����i@���2�%.�c��xrt����<���OS�����Dl��K'�G9(rFA̗:�N�H駋�7�Vҁ�H�ي3Q�����D�>��[��{g��%e�IBg<j��i�>ܷUEY����jk#x��Q�JFb"�G�8H���69�J۷�k�'�O��3��q�����`*�n E�r�>�腝��m�3�c�t�����ʇ�-;y�0�z9�^�x���������B�3����
��7��}ka��x":�����C�G7���`�������ƽ[�A^S=��vC����������o�k��,�����#X[���d[�/���|�R���5����2�h�1Y�Q*7���
�wuhR7��;�HRyݔ��4��mo8�g��.ׯI����zxL+j��EuΠ.�Y����/�8��p��ŕf�eih��I�p} .�&�f}�xы�����k]�Q��w^)+3i�F�J�O�?~��~[kx{��3�Df�IM��^se�Q�[^;�J�t��:��|�U��u�_V��,�p�8ډ���e�T5Eϻ��N͛GF�%����vMK�솨��S>__��\V"k��$t3u��W�s+zf�[e����Ьm`�t2G1�F�����ïm�Ֆ��MC������1[R(^�q- �������B�RWW\ا����"�`ѽ[s�b'��g��v����)�a��;�K{)��OI�w6��=Z1r+*�[is�g����t�%�l�����z���[|6��{Λ1BL���Ÿ�^TN��qyjD,R�?D|��KT�r?��a?]����?\�}o[�+[��glއD@G�|�G:
}�P��	SJ/���r�WZ�N�o+d���F�tM3�
�2}�I�|��=ВƷarѢ�������VT�������e��'uWxI�t���{n�\�r�ʜg.�ѺؔfJ�r�ҏ�N_G�K�;'7\��,���Ӧt�u ��y	��Z������]�I8sy��5�c���H�r+�z��o���!�ͼN[4@y�ޗ��3|Az�꯸�'���]!��i�Eg	�W�Y��t<��U��xxG����n}����P�*ۤ�֠n�U`b�jA{���Q����9��QB��Dp�2Uj�B��QZ󦎫	>\_�#1��+��o[�cb"w�qmt���`b�&3�P�Y\Tx�zs���mt�`�ҫnZ��&�P��x	�f"t0*��GK	�,*z��u�,Ț�7bqζ[Y͞&��{&(��O��o�?��a���.gW��0/ܫ��6fwe'Og��2�m�Ȫ�j8��m~�_�
��	��h�SjD���!Ċ���O�ۣD��oe�P������h����,��	���f��^a��3ݨ˴�;���v!�:/�葽�����#!÷���9Fd���A�L�mE\���]tf�ܬ��m<�׍L�˛E��~5v�.���t���bS/�����~c5�&�q�sb��K��S�_?5���,=D�����A��Ҵ��{��Y��WQw񽽫�Z^ ��k���'W�n�
!673P�J�#����J���7|c�3o�=������Z�&��#"��U�Be�
z=�fQ�:���4�֬j�pj��Vݶ�!ӕZv����x��	�=�ȅdע�%q
q��|�Y�� ﷗���jj
Tkާ#~��.i��AT�B:�<!v�u��>�o��OI�/'7�$ITR�P�@��s�V�E[8�_��H����B
K6;I"��3�k����G'�'_��x=D�)<�}r�����=:�1e����p��Oo�r6=<H�災)+�ȫ�1Q ����g͘�L��v�5�Z������As�ۭ�#m<ZJ��*\���l�m�:��k*+{GKGVͥE�k0�h�}ۍ���d4�W-z)(ұ�^_���6�YR�M�������R�2�q�5����ʬ��=ҭ�4D�鰓��y��ߨ��{J4��+��#6���Qv����lM�#�[�rJ����h҅���%��V�Z�]�[�1���/9��ICD��R���ЧN={��yO"���V��5�F�}BQU��vųO���B����҉ԧe�Q^볘jR�&,�ꌘ:�� =L�;i��4iͫw����;�\Č��o7��vh����>?=F����.��9C$�����o��ġ�e�s^�5FJG�V_%�_eR#���l�7�!�q�h�Q��;�v�N�; �p([���]ǽ�Fǯ�Θ�ͦI�tWx��I�c�r�.�e���i�g@B��R�H׳:��0o$�)���۩��u�M�C�Wf�1n��������5Qy{����W)�O��88Me����+=�|>�\��^Q�j�S����P�z�l�54Х��`�t�n��N�G;hvdړIv����\�u�+��Ĝ�/4�2h��â"OE^%����,��L|lɨ:���H4�4�R��V�5#ii��	z�� 0�BkV���k�$ǌ��2uߚ�#ˮ�wtG-��Y�-�B�U�����Y�<���'!�����)Ծ[��?-�_�4ʤh��:[�/�h��[t]����N^HvA�q��ۺ#~���H��Yd<~%�#��j�r^�ڬ�9�-�y�mnf�0�x��lp;1V�S&�\B{H���?���V���=[ww]�T(+y/M�I?��"0������G��tcّ����;>j�S���2.�#`S����t>�>��
���RJG~G���!�y�|O;����TH~�?����d�zݿ�k+r*��t/L~9��g/q��Vh�>;ΥCv6S0Y}[�C7�Ox
��7��q�O���u�yk��f���&�{[������	�nC����Tvf�̈}3�z�u���J��,oPG�(qޥj�<v���F'x�����W3<g6��w��ǈ����T�q�K��t���=gv����q���u'�y2}0�;�%_�u0@��F�_W�%b�Ո��ƋνTR���cdX�@��tc�V���?�g@��0�І���^���q��]K���6<g9���3k��u���{�hEkC�_3�b B����h�:ϡ�lk��n��Haؼ(D����$<���ܢ�lP��E��`���EA���8
y�qs�A02����]�լ�&���b�\�T��)�s���@������vq6Z�\�d�j�<j���n�x{ Z���� A9����I�G����"�g���	\IWk+z���nVG��=��g�����'s���g��[7Bf:�o������Wf@K��)e�9��f�C�֎�ps����&�1��B�(���g�J\��*�vA��qh��x4հN��3'.��]*[��g&�9"�"o�H�AO��]��X�y�7Q���⚞�lɿ���'�Aw3s������K��[�Z�Y�U��z�؇��=4Kƚ;&}Ǌ�u���u#X85�[Bx"���De�]���Q]�١���x��N9R|�h�>Ż=������@g��B�T>��p��X��&��~~��g#a��L����.��꣨"eq~�f;[A��j�j�ɜw3�q3]�:a[��wO���9eP���}�&�S6
$f�-/�ֻY��V[��}|U �oLF)��/�]�����WC�))�&z_���<��?�s|�B`�Ԩ@܏V��~�-��A9|�i����`��cw2��fHo���Z�ù�nT�+~��N�i�5��|�$�Ġ&iϫwnV�|U��k=�g^����������h��'�Ō�;;;U=�כ.kb�GC�N����͠䗭�s�"^3��R�.��k݇�Y���z9e���7�/�jG�����}�Sfi��>�'��~���}F_��K �s��`J�17E�A�n�4��ӝ��ʋ����tl��_H���3���e�{����y���+�o�<�K��f�s�0��{O4v
:��y+�b�6&��;��]�>�5>tJ��hvU�Fi<J�9�Y@&aufH꧇ӷ���9ٜs�Jĳ���˕Bd���|�δ:|M�������:�̷�V��;�vU�]i�n����
�XF�	�B�hE�.!\s5;d�ћ����v������=w�4�}AR(G\�ox�uڱ�r���ʷ�]�o<��O�ޔJP�l����H�g
cP�*�vi�9���^tp��u�գ�_wO��49��*O���'h��AQ�7�m��x�`��I���3��2�[����)_:�Z���WW�Y^�����X+���;e����m<p�r������.��M��JY����eEx[kv.poHA��Qluҷ~* �{�[@k-3OJV��d��:�`�Q�;2Vbr��*�,s;ݗ+��*�H�mC���>�_S͐l��i��_f�N�4�Oiu����-�1Cj+�>
�TP�K��u�5��=üSMv�w3xw��[��-�B�F��-Do�?[?0��Eⱕ{�<ׄ��v�+�Ө�<��Z���`�<댈�O�zxE����4����
���=^o���p�����0p�����7�8(��n�'h>k������6�;���}^-����Tg`���������?]0��ʻ����a��֥W,�V�H��\[aj#�I��v���W���8��T�����
H�G�t�W�Y�������*�`_Y-��g���-��z���m�'�j���i��pO��<�E#�����>�$w�/2ò~������8#��-��t[����>��-5�����e��Bè�5;=6�nkߙv�����u]����<]^�F�ק�������_'9.IU*��H���/���"���N��qǆ��֕�ZW��e��P�!���!���!�ZZ�VY���eYejh2�X���2�e���e��!�U�Q��Ł��-C-U�C-U�Q�U����Ő�!���,�Z�,�-Y��X�����jd2�2�e��!�(�A���C,FZ�Z����-K,�,�XYk�K-Z,�Yh��e�ũe��E��-+-XYd�Ҳ�Ţ�%�+-Z,�,���Z�]�v]K���@e׈-P2���� �2���%�,��j��e����@e�X���d:t.�Z��(d���-@e��,�e�r��kR��� �$��C,�kZ���Pe��� �Ӣ�5��Z�e�C[X���TZ�d�ma5�Y�Z�[Z+��5�ȵ��e���2�e�2�k5��!�)ӧB�C,�Y�2׆C�(�Ue��Ue����VXj��j���VZ�VYG�gݏ�����(+j��ZR5���9迧�����Oi�򽝟����o���'������x�o�q�Ns���}}]����IU*��Q�~���bP���Ī�f������h}3���O�����������o��/�zN�l�|���x��|O���m�j�IZU
l�&����ah�^���d��c c 1�2���@jh�d�-UVL�Ť����ѤM ��,-CSUjZ�P�i����dj2d4h1��Q���d��UkB�7�������H���؃b�-�^C�������_?�Լ����꒪U��������C�׺}>���p�����N�m�%T��y��=����;誥^�UJ���e����*��.��T��×��?��}.˩�<1��>�	�]��N���J�V�G����d��|�y������>�7�׿��?p��~���$��v�O���D��{����M���|����}|>���z����N�~��xN�w���C�:�>��~���zg���i(U����:ġW7��ח��v��r=���PVI��Z�g�@��v` ����������}
J��
�UJ�*��U$T��
�%%�1$U
�R�P����P��R%JBP�ERU*B�U
�%BW����V�T*"ATUD�)DRITU�PPIHAEU*DT�UT��PB�d��R*RR*�J��+l�)���T�"�B!R%$��BJ����T��T�

�
EURT��J�T��H��QUDUEt�B��T��V�DR�$T�  ���2}���n�݊��]*��3]�s:�]��v�V���eL+i�5ݮ͝j���鵝�6M+m���s�A�jT��
�����M;��M��
E$���D�UD��Q�  z=
(P�����P���hP�8����(hP����+����yՕ�p*��h�.��wk��E;�]���B�˧��h��@�j��껮���q7GT��P(�QE*�
��   �h��n�#-�r���K���sm]�c�[��NJ�'�WcM���b;���v�.S7w���8����띥i,4��V�iII�l��B)*�HQEWL���   �Kmm�v����wMn�i��Ķr��Ll���ۭZK*���\����90�\��KXl:s��IsK+�k�����R���� ^   rU@k=:�:VU����]8Rڍ-�XZ���[@��XU)#���k�ku���:$s���T�B٪H���  �U
�54E�Հ��N�j�J��M��4�ڣQ�tmP��)TګR��sKt�	WjjV��Ӹ*P �TU!��T*)�  }�}��PE̦�]Shj��t9��jAV�m�5��P  � �X, +�������� �T�T$�*T�K� �� mT� �;�e@t�� Ԭ  ܣ
i�ܖ :�[�΀v�Υ�@P�� �uI)PR$@(U*�I  �  w� :�5� 7P� E��� ��@� V��+�t���A��ۣp  U
�BR�JQJUT��  ��=s��܆  �X  E�C�C��p` �uSt�T ;�VA���+ Am��� � �~Bc*�H��4i���$��@h  �����*��d  O��*   �@eJT   !)6UQ  ���]��W(ntC����l���NF�=@��<��l����;S�g� {ݹv���E�U�h�"+�� DW�YPQN����������ß�Z�kSo���7Y����Cu]��C���o�L�Ӭ��dBi�o*:�l�u�Jt�-J��h��
j��̹���F��Ӆ�aG{�,E)D�D^�V�i� �#Kp*�Mhs"Xv$J8w)f��C�dH���� �9�Fԓ^�v�Ҏ���`���[$B�M^�6��PyHϵ*,顏jފ²�֤2w8��7%�;O鵇[�p���M��!�c6�<�hW*֧-X-�-,@ܩv�8>�ȶ�eK�N� oqe�L+�$�3uJv�aX�n�KA�,+�7[�wX� �p��6��xѠ��^a[@�?3�C���h�����k�%�N�e4a�[��*�#*4�CLp1X��y�uC*f&��u�N|��{����̺VEl(e��wXފ�w0�`�sm�֜viS�U
n��5���E�v�+���I��	�jf�ǎ�D�V��qϞ��p��*z�Z�f�  zlw>ywSZ��ߎ�j�պx�*M�@�B�-q��Id�a_Cw��#��Cj� �'(h��P�B�@L#�<ϲ�m��kHɅLWm֩�*'H�!�R,f���:TF,4�Z�����ttV5��VrjьA����bC�2�W�6\d�%mˏ��k���f��[I]�d���Y���@�&�Vةw����խRE�5��N�t�.�K��HNq�!�33�n�Ty��H�K\�.aʽX�e�AY�z�YI���)E���]k���̑�J6N�W���
���qU��!�$n �m�z�"&ۻ�h�K+Uh[F��Գ�ӀmKق�fL�ݢ. �@	��B��1��q!�;�Æ����)v��d���2�"�`t��KBYVPt<vLIŎ!1ܹXq�)��Z�tRd`Iٙx�U�k�,�7���*��3Z��lS�3az�:C�,ۣ���XM�Cl#tܳ�S�=��MS��LI�.e�[���f9��V���4�M�h�F�b��P�zX�s)[���3mڻ	�'Vk	&�N�m�mB2�k�!ލQ������O2��QR�ㆵ<n�'�$���� 0�x�i˱��d�ׁ*7S���Fc&=��<.��n�WW�m=���5:��.�������@-Q��@�Ӊ���qR6��P�s/*ݽGsb�$8�Pى�l5��j[(P�	�l�,c�@`�l{m6#A�e�07�5�%mi����k)	)�B�Pf�[�Hn�U%ῆc�u���b+ci�;�q ��Kr�;�F��'�V�:`��(�ɀQf�=U��R�0��	��Ϝ��Yh�����t�����5栢��ܡ/!���S�Dx7 �:_�ゆ�B,��هl5vv�"7i'(}��ٱ$N��M�G�^L���Z)%���� �B�� ��7W$l�ջV��)��b�L`����{O �a�R�ɧp7X�m�a;A^Jz��mM&�<#j�(i�d�=��m���
���&U���n�v6k�AXWKh �%`���B3^�������s,�7ؙp����u���h��N�d�lE�'(FZ��-�ؽX@u�aɚ�´6�ɨٻp��\E��A��P�¢[��*�l�v�5!��V+n�;�H�����^��YW@�0�".����hKa��c�Q����@A�upj
iܒfi��>f�U�˫e2�	��'6=KV��W��ڳv�͗.�pਓrV���F҆bC��-� IE�־6���ݍ[�[�+ V-,� u�H��>϶��1�E�!���=Hԏ\�!5�bR�ټ�j�U,�v���:r�X"Dκ"�VF�X�:KP�7]�����[ 6��]�.;�Xeb�dF̻׻K	�:�,L�mk[bf��{w:d�o����֤,Su����귋D��k*����v�ἅ:�e(H1L܅�!R��v�
*m��f��eJ61*-f�
'���ћ�����t�2��!��7eel@-�n����(ɉ��@j�--[�,X×��n-ԄB�ܑ��3�X$L��lT�GE��@�Zc]XȖ�m0�Q�����U�l�CK4��嵖�nS-P�����L�����J�7����n��PQ��b��hl+�0�K$~Z�MCt,e%�Z�u�����hɐ���z��ň�.^ض�4+!CJ�n?�2�5�W.�v @3sk(�btw.6���7bcǢ��''uz�e�l6(f[#��V-Ki��wf��(5�5��ҭ����-��1a�XE-:Ul��DF�,1Hس�I�8�&�T�G������{��X�q\�T�F��H�k&sW-�V/4j�ى^;­ [Ƣd�s0
t%e]�J���fc�8ʡn���2PM��~'dӴXui`��^5y�n��5;�tL͚uD�"���81h��I�΋�5@ �ԏ$���֐+�B�ml{bdLܫڹ]���7Z4mdN�=�*�u���%֌��lR���)�q�,N���NV`�T*Q���(:
L�W&���{��σ��u�،�I鱺���6�RG�����I�d�Y(H��-逜�,H�A���[�u�4p�PEy�j����R	z�ʗ2��tA���N�l^�吆����Z�ۘ�>T��4��Ћ(��E�ܑYU<�"�V)�y�a���̸i�bҩr֋�]���KV2��LJD�0����Ae����7��2��-���͢�q�'QSI��h�F�1�v��t�?Ef0�X'E�Y=��-��w�B�j�WL��)�a]�J�n�#���e#�*ؼ�p;%`�4�(�ґ�z&��t���=�M`�Ɲ�h�ᙂM�c�/[˖�-�2��� lŎ\�s,:0\�[�-ke�m���H"����nfD�k��!(I���KM�Z,Ђ���[3k���7�*�ujٳ��_ӺNC�-6��//j�M�-۹������Vl���X�C�#�e`�F��Z*^�@Gy&͵��4#.����X%f���6n���nF����b��m�Ղ��������	ݒ�K`M�>�l)c��nb�hXb�pE�;�!���,fê�b���L)Yn��Q�MV����Q��G�iʶ(㥀|�� ���;���=e^Fo[�Vb�+buY�ct.e�YXm������Ӻ0�M�sn�SS�.TpP);��u���T�(�+B���t�z�J��ݧ��T9�KlA\�r���w[yi	Sq�ȐN'{��h⭂L�M��Z$%�B��nV�F��ܻyW��v������sM�6��&��r,�
V����;�a��o@wp��N�x�J�{�M�O7,�U��6�4[����^Ѳ���d�����$�c����@���xP*J��&!�F>xuln���[$�L�a�3[l(ζ��E�k�7���`���"Y��Э eۼ8�%eʵ(�I��P˷�*X��,��-��ΰ"�����l��T��0?���)lvnxN1aZn�aP#>6GRZl�ɺ�5��@v,��ʌ���Z�ߎé[�e���a[�� �4�_�� ���b����+r�j]F��­��1�T����u.�r�[k\m]�����CE�P��,'W�u�CTr�{kA8���V>92Ѡ�j�I������l�r�qZ;RE�n�N�ٓv�#r�S%V^J�A�tf�cr|��hX�)
2��.a�G+M�B��a�5Ki�0aL��ݻ�n���X��p�ڗ�DV�W�{��R;*���[�}�����oe�%tLeP��T�C�%(L���+�׷v�(b[p7Oe捓L7+-@�&Ir���X�D�䂵ܼ�v~fCX�Z���ۖ�:�m��[5a'tE/�F�f�R���kHG�xt��1�7�	K��Y�YBU����p��ڬe��4�J��%��P�мv��KƉ�\+\{{���"�Ƥf��uz���d;#4�xY ?�9�-�V�^��r<�tɢͨ�	7@\O�NS/n�O����`{6�ww�q��M��V��!ISoFa��pe��ךt=ȭ=Ү��8`$�Ɋcӄ�����؋6��Q��[���f;[2���g�ۺ�P�3C!����V-��3j�`8�I�6㭫��o��U�JKbrn��7m[9Y�U�Cr�%��)G+#�^`4Fl�K�c�4mm`L�0Osj1���i*24���1�&�j��˃w�ʬ�q��U(�1+M^Ɇ�,���.e*nնA��U�R�#��NLw�1��V/2�� �ے�0��u��#O���N
p�[�vb(Y��-�A�"[eV�ŔmL�����X�~X��
�L�A%�
ܻژ��1^sw�[NEf�XX�L�f]�vΖ�Ћ-��K(�&������4i��5��QI���ڴV�)P���V'���ڼX]�JE(n���xܸn�߲fn�͆�D�xe$��0ہꦈ�maL�{p ܱ�LN9c/r�j�K3c4�Jŵ)仢��,�*�q��K^�A= ����$�!�Z�y�Z��%`ܺz6�����,�kA+��;/ѥ���������3Q7-�dK�Cu�.��%)6LF�9/����q�z�[U���������]�A�{s�X9+&聁�!��"�7xt�#��((�]c���s
4�g�):��c"Ĺ�YX����9f�g\V(�'#�.���b�^ �uh�p�zюÚ�f���+�t�,7Yˊ�қ+3Z/V2��Y��K.*��-K�pkwK+)��B�.�n`�	L1��!�&�n����[MR`�	�d��k��Y��]��j0ۼJ�:�m�VVۭr��[����2��wZ�Ы`��@A���NlG�;��,�	f��P���9��H���DR��$Ve��N�O6�Lx�1�9��h��\�q�+RrXӡ[��J�A#�v�r��F�Ot	sbD&��T8�6+�3)����F��p�E�%l׈���� K�f�6��sn�7���b�PT{XA��nҘ�q4�ԑ��M'cDK+ "������qT-e'v��j��a�D�1/NA��Fch谰Q��:(F�]$�8�՚_b�r�F
�e��(�zZƧn�#OuzJ�e�uk膐�����a���lm��G,���k��b%[E���(��o�Հ�h0��s^̻��/]��Ehi`�1,l,�p��K��嚴�D�,Zo��4V�ȷ74�يn�bڼ���)K�j�����j��C
��&�4����kCCe%ռ�t�D�9t�t���+���\Mʽ��,,�z
c�J��W��H �tkm�r��he�К{��(ͥ3p�ue�(������v���Y�.�EF����B���^\�BoFC���MT �Kp�ԩ��c�sC��J� ��Ֆ�����Z�rZǖ�]�Z�iGr�̚�=a���A&�
��Y��m26�5�'z�(�ɲ3�x�
��1XV@S���R��V����b�3T5���l�^Ǧ[��Z�(֦&+l3�%��譹c�L���3o��`�F��А���[�.cI��#FG�-NVh�2	�wa�i�t��a�l�R�X�1�]L�A�̭h�"����Ee�oMܻ�itI�r�Ƅr�/m]�� Ejvфhײa��)rk�Oj��f
�P��Aw��f���^��ǿ�e����h�u%+��
�+oB�LɁ����s�����ݫ� :7�i�GJ�j<H�K+/ 9u>�K]�O4X����l���d���
*|��v�Ջ�1Y.�3*[�m�-ǉ ��C(l��[3��K��E�n�[��,֖@v����*��WbkwmVZ�R����g.�h�"�)�w&K#[�F3�ÄR#q86n�����$�Y�5��){��XЩ^w���r�0Խr��� YN�|�N S)���uHu�[Y;H���-�v��ו�iP<���7��W[O(V�"�4�'�uSݶ�����Z��f�k���j�K10���쿐�zƼvu�b[^��D��������j��5�Z�5n��U���cZ�*��� %&1�*$D�ۺ�_�q�W"5���ꆕi��*?���H�e��JJg[�ȥA��"�(���%^�3&b��%�IE�'�R�[hGS-���n�,���n4��G�%m(I��j��dXf�����"[IQWz[$�P�YJHbջōcĵ�j�Y9���l�i{j�K4[pd&��� (ZN�D©�"VkF���f��Ɗ�mKŢ�M�v�Hh 	x1�K�) 
HS�t4��Kf��Ór�m��IH%��8�4%]�.���FV$���B�w���t#(MG��ֱP+��U�@aZ���e�
!U�3P��F�V��Y�XMd9yM�V  U��M"5���b��)�V���g(#-虲�u�
����ɠ���J������ ��ulM!d�PX~�XF�t���o���Wr��30�#���U{�c�Y�����Ɣ��Ĭ�&h5��3�QۭHJq�RD2�����\��ufմ-��Y`��\��cpŐ�q��H��ʻ�h0�Jz�`/���Z�Z���U�^ڎټ[6ʣ�Q�,@�MN��ᵯR�ZI4�+���i<w����a�YwC.f+�ȅh��Z����Z�!����4�����1���V/2��ByI�+3��6p�on�¢����jD;�5�Áƶ��ާ�|s��ަ��z����u̝�W�ڽcv(v��^ȡY�CDN�9�5�1��j:��C�S��Wh�x���t�A�+J��E��i���K�-�� ;isOQ�WH��_��py���J�e���6���RڙI;�[v��ݪԝ)V���)p�T۩�WK�aIͳ�e����}���+y�d����F�(�t�eW7�,�.{�k�C�K�ˈ۫�7P��}u���J�ք��,�Rouu�G��/�3+��R�IG��7�뙼���Aր�"�|������6d��4����m�'�Cur�o�L��]ݗ Y ���n�I��K��h�<���\���Inf^�$/R:v9���y@��O�n���Y��m�'V�ii(�h�e�7W �i[��E.:TՉ�t�{�] �Y��\��ôb�\b�f�r`Kw	�-��9�k�b�׈����{%U��U;ul�c��I���ra��z�I��ݩ�\����gR����wRՉS���
b $�M����}Z�C�6/U��^�	��Uͨ�4����kq�;��a����)]]��qk�ePG�T��ڹ��1�/����,\�Yʴ��2i�m:fwy;tr���|���Q�=��1�Kxr�n]�K�n�w9[ֺ�xOǺ�a|��E�WZ����f8�n>4�H�,��Ն�%�]����b��Ok)�R������O
�vv�˜����� .�[o6�����>�Z �V\X��ve�f�mR^�!�9��!]���Q��Ն��/^����+R]W#oXFR�ugZ���ՏZ8s@ʫ�U���z���"��S)4 �8v�'ǲU�݄���ﷅ�w��>H%����
Q�2���ư����opq�dփ�W,�gV��m�]���j:랅3�H��M��(d���۱Q�5���N�+3���]-��u�Z339��I.����=��f��2���6[�3256C)f!]y�Npvn�u���������n���#9��$*��^|:�h��sQl+�CVDE�[����Dva�J���@�#�dns�Y�:z+��f���� �
�b^�ٽ�4��ʷj��Z����w�a�)�;mm٨�����X�;��J�}�+Y�s��C��ዓv:���4�*��n�4�
R]YYۙ���"�q�V.�u���!_;R�9N�2Z�w��;)�^����z�-�D㾥pƲ�u�:KТ�9�� ��a���`�`�r�h؄rNӭj�N%j�kmW'gu<��ʌm�뷊���l�)wwi;�`��'��E�����y�1q���.��i�ya��2u`�_^Q�]㭁S쏛�]�D'�V#�F_uc:�X�j����RH�I���n�ow��M�ՠm��	=�ؕ���yK�PMޫ0�xC\�{]e�g�/d�,����]�uw`�pv���]Ar���lq�TIԭ�d$��\��'&�y�����7bs��*�`�:����ܱʲ^B�+�]�aE��v�M���\	�fS�w�2ݼ4Hw�%t��k�p)����_r�Z�����|�rw�7o�U�|�ɰ�G3]�c!�$
��[�Vh�Y��gn�p�RLPwbP;�5����#,9+:d�5�Wp�����q���nq�F����S����f����*Z5�ceg�EWu��mwt���w-��;�0�u�5a��:��\�i�.J��{z����L�n�G�l��5�睤Zf��WG�c��9tK���϶��n����\�0O|�/8��X�:qi:�Ě곮�YҰ��r�V�h����C
 �����pk�PM]^�Txc>��	�֜y��3�Yʜ '������w�?�FCX�
z�!�
r��:�sZ�yٱc���I��1:x�(<��u;�1�.�3�tU4Q�{E!� S��WKQ��X�.��m�t���C��ӼW�Z�;ɪ���#w�j��#n95ȗ��E�Oz�;LX��/�;�o:8n�-��n�m�L2�J��;N�s6%r�<�i�R�T�ie���Y�rt)ioqaSn�3GKL�6����ŎT���i"M��z�u�靠 [�c�y8h[�j��(a
v�^]
6v?�����G)o��X_dPUK�{��j��@I�*�mC���#8]��RبYq�J��%���B�I��i㰅7z�[׼�`�zj���j��(릨���uҍ\E�[ه����"�
�ʟ�Ú�L��|���n�ԩݮΠ6�4&��$܈@F�ؗ^�sX}ݶ�2�c*n��H`;t1��
�eՕ�tM:Y�݁R�\����D����o���W_/�n�e��wR�
	���}�}�p� �u}!n��V���c��~�⦫�݋j|��C�f�M-�܁����ܔhR�!<��������m>1F7W���7T�d����ύ4����*&�MG2,�'2X�셪����`�!F��5"�*<����<�T�j�9�W8�4�eE�u���o ��[_g�k�v
����rT;L���rw�Ki.�����.T������[�_:��!g�>�л{��u'{Q���N�J��@���n��M,h;,CV���FuP��\H1�/9�쌲�n�i�V���-�p�[:�C�lF��4���m�α��e-��I]Gbw��#n��o#R�/x��{b��>U����AcH�� ��SM��sźL�Q�+C�a�H�B]>ce'`+��#��f��M�:�6��*��o�ӭ�C����)l8�,swF*Ym�v�K\�/�G�XC�fr�At�L.��}s��jGyxW�n�NQ�C&�����i��f3�^J���.ek�*itT/�k��er�Mָw���X]4̾���T���4�uc��e"��lK�nA�q>����,�T�cX[OSV �u.�Pbi��AM ��=��-�t���;jg^M:KB�Ĺ�����\�����O1�� �^n)��V]De�a���m^ΓP�2����ۥ3��"c[>���cC����+�t[���W���-�@G�-8(���Ag�d�����{{�scj�I5��ɠX�����d��N�d5ܺEݚ�X�0�2�^�2�u�BI��iծ���l��qH����67+wW_�����Q�����S���2s�8��_qox
�1�}��DȤSU��yw Z����"��j���:]�YwF�e�uz����_W�E�����e\���#�(4�:���%7�k+��ۡ���%G[���>�]ɘ���p��*9�f�e ����u|�8����mд%\�ټ�:s뎗>	֪St��ޫq��kӻ�(
4���e�L	j��vJ�Y��7T���9�9/ۚFl����+�C��o��Ֆ7����5�d�$�-,7M����r���뚇�D����޳��yS��--k�	���i���o)�[n2�muW�JP�|2�^�Es�θ함4.�a53��ǉ�ohv��Zv۩�c�1+���|q_���R�E"���5LZ�\��ֈ�	r�B��x9k������m��D��>����(�J�Y���c�ׁ־ZV�h�'rK!e� :�chefZ��-nLɔ�w��_)ÏE[y��Ǻ�id��)أ6�1h	����Tk��;�K��\ے]f���}�:]�d�]Y1g��I֨��W#j�k+V2S8���o��#]�)P�\��L�D���W��q�wt�.���Y7H;�i�켚�"gm�3��� 0,Ь�5q�\)_,�a�$��=Ȍ�}\8��;i]��;Aw��z9fγ�N��Æ�F�Ǘ�㘎��M�>����&�����
1�lAv�������rܡF�ر�i��(�K��]��V-%w`�<\j37��|��W\tsab�A}6�ԝYx��+�|������r��#�Ö��]�HS�N]�mU�ɓ�ͻ"��7�b���y�IZ�:#�s�����أ\��{�}i�34����#�蹻Fã�+2�hޏ��o�r*7}�e�Ůku�u�3(�Hu����:xu��YoI���\H�q2I�z����f��cX�/�$R}�F����ܢW�·F��t�NA/�P=媣ܖ�M��f_�W����i�@ຏ7��x�^��hEŹ�>�ub��@�vx�f��,����v�`�[��)��S)>�ZV�O%\ɰ;]�L�}�19�7�m�d¹�l�� 6��9!kvu���=�T�OxL��?J�^o1 @��ieD*]�B�����|�{6�õaS /��$(6�[���³V�B���-�+n����+�}���A������yP�5�dcрP����ʵdʉ��y�"�x܄��s���N�Σ+V�os��!l��<�4�}3'ks{�;���9�K��U�ū����h͍���;���G�f����y��逹 ��J��������c������WҰ35����ۼo�#��N���nT����k��`M�[����oLƯ��u&�쪴��ӭ�,�E�Uf���E�˩�{��f�q�v�]F؈t,-X�F��#9�����c���p�FS�A��`p���ԕ��1��3C����=�=��!Zu�=/�]�{_(����*�Iu�2����(�L|��|���J|��x9&�V�"���ݭk�-�c����u���l6�*u$�c3�yS"��`�;g%B�����p�,�9ˑQ�Q��Fs�[!��.�ީ���7������w�3�0��DD�"���9I�Y3�=���n�}�7RC4ժ��+���a�����nwd<v�������妭Ѳ�vm��;0H%f�/O2��	�껼Y���lIk�;��j�X�������R3��jc}���M�J�7�4<�׈�*0fuMs�m�<��.X��[!ݼW�����{�,sIV��}˰𩄁/7����Rn?���L شEL��M�пz'��^ �Ա��S��ݷ�	A�]��QM1���9N��U]�oe"R���k���ۘ;��)b+�n��PM�^�X�����s�o'�5���3�"���we�葅���ҳ)�+vQ��������\�*,�`�����;)VG�*��qEt�A9�9l�U�t����v��Ƭ_���}w�g)T�F�_d�d�K5�ll����%罍_���q�3�M\;��D�QU��#h�<뤻���>��ɵ7��!9,�;Q�� ����[n���Prni��ݿ�I�nW6��Qu-�gL�/5�5�X�|ũK�N�	�mV���u0�ѵsU�)1|;݃�:6@8ixQmgi�7yr��ʗ���cx���Z��A[!�؇�k���ߞ���AG��`:�r�0Dl;U��j��JQI�*uj;��A��^-+��Y��mo�1��k���ʖ�5�d|�B��i�>���n��9�Z:��N*^���k;��y��B���w9��6��B5�J�p=��u�)>�Mh���5K�y�֨��<v.Pr��3gz�#]:7�Rq<��7W�3z$]vY�4�8e=���3��q��MǮ�ֆ.�ɡvqx��L;gǊ�}ٔ;*��o zj!��z���^�b
MՅun�t.$�j�!���mZ��Jx	�;b���4=�����'v��arv�El�qjǷ�����i��;�0�����v�V��:,;�Ww�aM҅^�[ A�V��mk���2�����g*��S�	�٫���E�\���m�. ό4��*�k\9nl��A�O7�Ʌt�</NDW���bu��.�l���/���3�>0ou�l=��f�{�vBWRs4CZ�]�:_=��BP�b����¦���V�&�ov�>�vAoy�z�K�裆�v��9ýʾ|^;�ֹÏ0"XE��.�V�Wh���3U�|UN)�<�����U:����ۤ%����wR@i�t�wМ�ZE�<'NG,��I u��%�6^J�S��U�-`���eN�?����k�<�
K�L�q����
/2��+{v�^*�f'��]F�d�r��n�J�L���Z�a�oB���(�{��V�1���8�㹍�"��S�B�%H1���Uܼ}�M����FL��<R��V[�v)_|'gmj��6�^ƫ���Z����.`�$<u�+^V7�jAE�=�pΨ���ͥ�+�n�ոw�ɹ.-0�K���^���H`�'.|*2<ݨ��;yBz�2|�l<B������L�5w��q7czv���+��Ṋ6�=Y�˹�`�(������}��X��[ �*5d�ѕ�]LUOuh(N񿷌D�z�(flJ�w^1\M.�VX�q��J':�]�i��G�뛽PJ-�@�"�Р�N�Y���N��r�]3���Y̋�vH{Bծ^�6�V�ث���-���\v��T[���G���L��`gB;�v#�"�ض�e'�e�7�Պ}w��U����n0�d�̅\���\F �B�VR5V���VX�.���	l��|9����<����@�򝫕����-�i��ە���3-����c��3"_;�@�c,V�Vy0��*n<����"�(�~c6���iԯ���^frd$��J�ܕ��s��gu��ީ&R���nr	�R�E�8i���q�\x45�%ϯ,��w3I��ˮ9x�dH,M�B.�7���㺞�Z�R.*�;�:wt@1�z��`�f'��+�we��!��\�}o&řD�}��D�I��ú�:P���N���w��+e^es�Ǝ��<���}c���j�ǗtѴ!jun�(*V"�WM�Z��Gh��y�6j=M��7;{��(��,޾7�ҏt�w�.l����Q>������ ��)�� DW���=ן߾����������1]��f�0��[/@�/�=�h��YرF�Ō7��u�N�F�j�L�Dme�hAE	)_7�+Ty�)ذ����3 �!r9��f��'�K�Nv1ܯ�@9R�g ��S��I�M��5�E�NSUtm�2=��;vmA�[��s>��8H�tB���ô짥�7[��� �x�e* ��B�q�݋y/���+��#\.\s���t�r��M�GL7�7�ܭ�� N��)��g�b�ɨ���᷏�>�{���������;����p�ܮk��Cgp�D�y�5}z���v�Yue+��M�����M�V
Dfj�;V�oI���ܥ�E'N�����j�ǝ��r�\����X)f�����aΠC#�y;����#o�ۭU2���}�q:A�PZ_KZz��6��u�e��#�{���ճ&̮���=�A{.�D���[���Uʸ��uǺ�dCd�$�����eҩx*F�a�DN]:�E��n��@�.�k�	k�v�t�r]Xӭ�P�.[���cY�w]!X�ik��݊c��s��Z���h"؝&��B.�< ��&;��ʓ)+�l��o>%J��dfb��ux�c�}��;�z��:�u4I�5��f�}u�%q���,;��{RґN�țN���*@]A��1딍��E�6�Y��I�r]X�v3�L����c#�M8A)
��z��㪉ru���oU�;�]m�����w�9�u94�.��N;7&��F�>�7�%�t\�tvۃsCU�Bހ7Pu�VfU��}��ܨ+����l�7�5U�-�'H��v�Ү3(:�_!V񵢚JC��)����� ���[�ӷFgi4찲�<(.����P��A�@��;����Q��HD9c4u�ʊ�Ym�)Y�U�.��	;w�� T����|p<i�dol��c'ҴUc��e"X��f�� �X��ݗ�dY0t��h����Z�1�	���9wsdwi���ݘ�}\��9��{h=���M̕fc=&١���v75d�X�4k��|���uE��H����9��tm�/#<���:��k]��6�U��v�e��\��ml/(v_U�'�p�t�Zf;�#�:�|��ފ��T����T'"�y3����S�	sjZ��{���=��h�Wz����0�\'(��|�!7U� P<gO�K�Nu	VN�����+^�T5�o�G���/Z�u��ъ�W��z�-�q�Y���ln�:A��9�U�%�B���u��LԬ$|�x��X�%�u���ս*Vֶ����qCE�Z��@�ufJ:~�ֹ�>�"��� �D�І��jn��A��V�Նe����v�.��X�v@�[���=��,�Y�����{�2�;=�y���J��wog_Z����CgZ�ͨ3��!x,�w�6计����v�<,�2X9����N���r�n-]|�F�����(�W��K=�]�}L�VoB�,ˁ+��#!�����!�:���p�R���	a@�us1��ަ���bS��=u̺7R͡,e
6Z_ έ�N�%дi�h�����/�o`
E&l�Y�,�\���h�ݤ��b�o9 ��:�ܮ������:��RO/�y��PшV���f*��C�&��梭�Բ��B:�omm�eob�0�@��Ҙ�/^�2�t��.�ͺЕ^B�̖E'Oz�)̻텮�ݺ����b���æ�]YL*� ^�1��/4,�xm�����`@�c3;k�oot�F��_,���<�t4��E��P�.Z�L̙׳�a�E�� ^�4)��5ӛ�� ���ol��p��ĭ.��g�;��	����t��u%m�WY͌��_d��s#]�뇗Ļ];�1��w{S��tڳ�(ގ���;#"΅���ʴ�����*����K3:���$8��kq��[�;�飗�iJ����C��>�6�u�I�Đ�S��S9uK�#���+Eŝ�H��Hn���	u���m�hK����Ĺ|��H�])�P@Ef))�;�`�/hN��'C"��]��#s�oٶ3wB��E)wڌ�];��!<z�B^Ǣ���J�,���);t�u����7�PO��ȁ��ZN�픺"��Zp���k��Hm�
Q���q�qDZ�q�իp�(�$$���4^��Uoktok�K���Pď�Z�Ęy��Y�S��s@��x`k��nvȫ%2�#L�Ů.ͽ�)U�ͼ� �-�+;��}R�vP�T+���a8{fS�ʹs
���rZ�v3Y����	�PRT2��Y��y��@V�<�^��C���õ�'[��>'&�+lR��K�,=�fT�<�Y��\��]5ۉPӰ�������"� 0�L<?>A������:��x���N�[��kU�O�@r��*,y�X}؞]%��:��ꇣ2��kF��:h4�⛑6�(:����anS=�蝥a�&�hM����6�h&o����Q�2��\*�+�j�f��)At8�=�
i�*<H>��E�S�9]w%L�~ב޽��n!�g_+Ϟ>�Xq��7�
N�k��v+��W�aU�:�bݫvC��\j�F����en��mZP�Tzҽ�E�m�).Cz�f��	�5wq��R��u�k)N�Z����sc�:��o:�����;	���s�:`K.
u��ȧ���];ֻ��u��͢+27��}��"9�LHP�ջ1tׯ�g�i"�ܹ�/�ol�z�3�͵@M���&����q*FWs��<���!��ܵ�݆雗�Py�& [ø�K�@������*��]f�5���-Ui�U-,9OlȄ<��ovS��]���Й�OY����[z�髮���fȫ�:Yulv�X-��!]|���)���Xw���"3r�:�,W����z؍�f����,���S��*�pV�� �J�n��ڕ����W�۩���%���v����rk��Qޮk�v�	d7X헵�s�Mb�O��d��w4L�Ѥ���}Ra��;2��>�t
5�ѫІw!����y�pP�'�V�%*N��.�1�vaWl�aݹU�T| f��{J	p���L�b;���&�b����ފ���s2�h{]���1FR��V����@r�G�n۷M`;�B}9�e3]��r�q^�!�^��Ġ��-T�q�N.�:ס����<}¦�}��p�Y\��Vk\ ��wO�<�j������;�]����RgOs72W�1D-.{��ϊ��L|�t���tloJ�n��Q};L|:, ut��4�2���]O����\ZŽw��4-
�a6~�4V��{�u����_f�B��B�4����`�߲��9���"|y]ց�o��o3KkhX��[�>f���0��;r�[Jf|��^��������*g��h�Ub�Z�����X�t�{���`Xm��$މiiĭ��#��R u�����ko��wŻʰYwB>���+s�9[r_"w�����Ů������u����B�}qN]��w�M���������W��t5�94�R�w�]nF.�{6m�}:�:ӭ<�g=U!�	������BՋ=���*��06w��{a�ޤ]�����U��\�����3�,H:��C���v�8�����&dbۙG��`�8'D�A�2�ς��N�c��-�ŕ|�0}B�!��^G�f��zX=Һ���=�̲��_U�����͝���C:3V�u�:�D�ۻ��}�%v1�g,U(ڭ}��A��C�72�e@U^ƬS�ۗ��nj�)k�:m�Q�̡�E�vrv7���4�b���k�Q�U>�XO���8d�jѳ(Q_9W�ݳ*��5'���Qh��y���f�n��97�
[j��S�����%_"�Wѭ&5��:�-b �3�^]Gq��n�R�k7fd��[һ��T�g��}�*b��>�B�����7w(T�qu��3��f��i���ev�S"G����	�k�u���8&v����mj�b�tH��Fdk1�:�
|F�M�L)u���Z�X7˗mY�)�V4������T��q�F���Xp�ˬ=K�VΕ���Vf�#s�Ź���B-�]���/[�Z�A�:��@bC�/fu^�Z�_.\�f��Cz������" �H�e��$�֜�s@Ȗ�;��C�-:6�_U�é����ӵ���Ϲ	�Y��,]S�k��99]���]�t|�i%�
`NV�m)����E��桊�+|fK�|��q��R%����x���#��V%7Ž8+
�����!�}�����r��pu	u`�%0s�WB��uj���С�^Mfխ�N-!P�k�c�OwXQ�¶�;���]6���r�݌u�5�N�u��Q�yoVQ'�cX��" 6Ne�8. ��8�3��'sP��{�D'c�:W/������J��vZ�q�t�F)N����x��af��D��y�^��t��KtH�`�	�:w�>f�.W��\OֻC���$��%�2�f�Xs5�dH�nH!9�Ok;M����#��.��Z�ع4lodӻ�`#�-��}�_E���

=9�l4K�b�.JTS_|�n�ٕ1ԥ����u��[w}FZV0��ۓ�$��/#�R(�M;�g04�+vn�@��G*��s���:�"�w���5�w�D���i���\o�vb����J9�G��ICY}h�[���i���{��k�c�M�Wڜ'3��i:)@������2�]kK�V�{i��k>h�j�ً�cRW-&���E���ԯ9���Uu�:�ԥ[��^���^�*f
Y#��R9V�/W1�DE>QO��{�s�CM��L��8��
�b</�]�wO�u�=g^C��K1J ��ˤ����%��<7�p��t�CѦ~��,NFR}X�0�!h�]�u�gS���O�7GV�L��vv������Fgu�:�"y���e����˩B&�7��p_�G09�\�e�c�C,ڼI�
���	ړ)��9YK|����ԙ-v
���Jmmw �r�(��1 �*F{+�vc�Y�p�X*��&ݾx*\�R1#tGez�»�����X���؟gv���t�mGQ�����	7[�t/(N����Ә�w7��}�[�],%;�-a��t�!�ޝY���U�OuK���#v6�k�|uP�3"|w���3��	:7�1�*{���P/rok���ru�0�I�h��	�%��{�(�ĝju�9w\e�h�֗_���k+y���	�8�X;�+�A����C1tū���]�l����PF�F2^JG+�C\l�5}���;�m<c^��U��N�!�\8<�%n�]��="뎥��P4xbgB,k����B7� ��x]��i�U��X�;��\X�������:ެ�l�ŧr��h��"S�bpV���d*���s\�*U��E��IK�m݃XFl\MK�[��X�
a'JW9椝3u;�M_n��}MJW��-Զ��lƑ��f�_fd�+�v)�ИҮ��@�f�R,jHQ��N��V�BR��wfK]��n��B���p����buK]`��YYN�����%��wC�j�_,<�
%�v�kS�o�B���4Iص��7��`�@SK�5̢u�t��e@�/�A��f-�Z���L��9��g��K��x��V��߷��w,��GOd|*k��و���8�g{�^s�R�c������ҦG ��n�5�E���{�����e��[���Ė�3/3�o��W�R5����d�E�V ���zL*�Ѿ�W�1ʚ�f�3c�^��7z��O+��W� sZ��،���;��v2�D����W%FH��E-�P����JV1�T��˔��V�:Ȫ�ܻ��,����@9�������R���}R�R�	���%4�u[z6<�a���w�b��L͊վ�X\O(������n��r#8+�ѫ���ob�.�x��R������S��6��V�ꨍ��Vs=���]M/�V�,�'����2�1Ogh�^�wM���n�.fva/K����A���"Y٪�R�ze�۫MvgMEe+�Y�1�q3�:˕�����D�lTbe�T�L@�#y9Ӏ_n�ԘN��0-.ݘ6������̷mi�M���O"ju��ڝ�Y�/U�_$Z��[#��G]u��tN�������Z�XgX�y��7��Pt�ut5���͋	��T�cM���ḶQ�YY��iC4�Y,vV����X������bSs~�=���siV\0���nK̝����2gf�Ruګ���1�t�=�V�Jyv{��a��W�k'U�����V*�Q`Ր�J�a)ڬ;'&���Y�1�g	��s��� �[��k�(��;���!;@�cF�Dp��
��ʝ���<�[c��n��T�C�9�p�2Pa��
!S�vtĸqXՍ
� �2J�����yW� j��S�:H���(�;�jdd�wK�;C�i*=��Ҙ�e��ccie!j���k���ːS��{+Msw[\BfL�.:��Ĥ燸vv����u�Ρ���C D2Nz�(�GI�ϜN�¶#�՚V������;�x�U�����y�;W�n���"� �V#}���Y'Sm8�2Y[Y���ՌS$�a�u-��)^D��3���#�)�5���b[�f* ����W*�zk�9��'k)�Kkl���F3��n�ܔ���mq S�����Uر��$���n�xب{8Wr7i �����-U��&�*p�L��v�1X��Ad����P=D4�b0�w��nG��:�](�[��u�8O����GQ�]sU6���� �����։���p��i;��{1�d���s2J�A�\�5����xk.�6�;��P��U��0f���j 8:7�����Z>�f��ټr8�e�JR�D�hv*N�p�[&a#�b�$��W�L�Jl�rs�(Ϋ�ٽ|��vq����N�f�d���V�G}z�#.?�U�}��K��}HIٷ��2�oXP��������㧵�Fs�Ev&T���1����,P���gi@>ea�~@�ggrV*Q���I�Z���-0��[CpP&�
�����WYY][���	���FV�.��QWns�m'r�����h����p�â�C^Ҿ�\l�m�h�INO)[�mų�*�����W�s���
��I
n��.�B���(S��(
C�^�n(��W��8;@��L��B�5o���9���q����wb��2ԋ��P���n\%�K��Z�٪�iEn�9tq]N=�K�i_әU�0Lv\<���V�;ͩ�o���u�NV�7��3���u:s�C'+�������a���c�o2��OD�B��γ\NWV�Pu$/u���J��ՅZ�㬽#��,��Y��������u�ΥA�ѹ@s����J�n�'�tiZ�<u��gٶA0'��&��s��]m��Z�1�.��@�h��%G�z��J+xot�k�b4՚0N�c+P�B����e� �w����ބ@@Y����M� �F��Jtc[ʹ�+Z�h�Zm��$�����V�mf1�*ڵcQ���86�AU��DmK�m� 4QUD�h	��X���l��j6(��-�V�EUV�[	�	��(���"���h�Pj�kآ�ք�&�*��*��A��16�mII��i��Q��m5�F؃lE���&�RS���I�ѪJ���ֱ:6ٚ&�kl�A��;��5��t��EA�՚-��Ɯ���J�b�Ś��փA��ыEm�cF��*�N-�6�lXΫEDm���-�Hm���Z4kE�b�����[l�m�J-�h�A���Z������j�PX�
i����J�4h�h�Q%D߇�h�Υp���9�+�Y"�i��l	����]v��on�s;��+g؞!vv���غk��b��r���bj��K�\�Oj���8�h���n��S5���\��z�J��C�4\W~dW�d��nbd��}��m�<G�j�u��atmA���q���=Ƭ+�
��'�ޜ{��$W��y����`:7��.��Q��f�DYq�d�Pþ�~�z�����E&�ԶqCӌ�[�H�LWG`\�O\�f���f��H�
��]!`�]s�^�o469]1���ݥB�,ʠ;�g����zg�����A^�[�<�~C'�f>\T��Y���vB�"o�����z0:��c�����*z�(�+F�w�89k�s'K��?Xp@��Π;���!���6<���yo����n���v���f�8�R�kԶ�ηm���,$�h��ѯixBbE�+s����߹o�����#Om��z�o�,~}c��S�����&���$�K�T=��SK�؍;i����Q���ދ�l�����o!��>���[q��*m�|� h�x�,�6[!��ۜ�ȅ	����,S��p̆sK}X$v���j��&�L��}+�L.�����n�zZ�L�pK.��g:�9ѹ�"��	@3�c�Q���C�����V7��]�E�����ͷ�of5M�S��Y�D�t�ذ�VɆd�vT�Ԇ�ϧfw�V��E�ё|��Gy�i��q�~n�WJ/�jUeޔ�YϽ(���͜Q�@��B'�O��xG�N���[*3��w~��7F��R,�m�B�w9�S��P�_x
$\�]F�����Iu���ը�[�H�X�v���ID�D��x�t๪��V&�<D�>��;&
���
+�Ձ�~w�ӯiwe{����n�����)���A�
���Up:k�~�@#��:�T{��gt�Y���Z��m�3nW��@��̚<u�:��5	*�WN���y�5�~}n�����s�=kq/{{����:��4��!���x�W����0y@�Ws,�t�n�v1;dNR)��LOpضF��C�֒/6\;٨�qiS��Ɛ��|r��ȸ1-�hy��E׹�+g�po��_���R���9�J":��qh�*�����Sٷ ���\ݣ���o����Nw�V���Ҋ�:Iw��!DD�_%f,u:���2����8h���nߠ�U+�n��QZ��W����zشk�9�����,�m<5�j�)d\��2l����gV>��ʹ����iĎ���[�����}4���G�d�y%iE�-�M�"�t��n���o0���+��Y�|��S�K��<��%�8��ǵ%̣�rF��bɍɠîܵr�nK�}9��V�q9��`<�8�z����pO�"M"ty��ti{UlŲlj�S�:v����m���Ȓ��ףp6x;�iO#�V�����x�Ւ,;w��9ߚ5�b��������K��霮�w]NrԊ�^��Ǭ{Xt�3��9uB��h��#�=�9�Y��9U�Z}�X,|q!��^�6GK��^�3��[���pxh0��X��g�1�+������t��|d!R�&�<���OhKݎ�]>/r��iQ�_T;�p};*�m	��(��8�B#�ҭ�!iw�LƂފ���0$��U���d����K�z��]j>��^�%xSbOړ�6L a3�-7����l�k�dу�=LOnv��-F��&�Lh�4�[��WK�G3G��}�����w`��c����b���4Ш�p㰊ݕ��ʦ=$o$�Ѱ�5�"��fI�D�#u��e(\.�V���<�b�ic���������f�%or�� k˚E\>���W��
V��Y�k�6��Fo��y��z��-K�z鸯5_m�����ﳫ�I�����r�]�خ��M-���y�K;�^����`����ӥz�ĥ��X���6O�J�Wr/��k�R��K�!)'DUlz@�J�B�;$��)�����V��5x�����̭��{o6x`�\>y�
���<5�݇Py�1x�M\Y4���b��T�NPn6wh+�e4bH��;�����t�{N�i׶B�:W٢h;Ҡw�w@��/���.�O�p���X�N������eo�)��@d}�^u�g,�����k�d芍g�U��t��4R��2�:��g�R�+5C=�;�"3���Fxz��;U�\J�L�:����|6
o���O�Vۯ]I�G@��;��J��,y|��I���X4�CY�.�^�(���)�ET2��fS7L�r���W;��sO����T~�(�~��c,xW.��v�kw�����Qe�k �*��g)����yQ~��Q���,�G�*��C��Wqݍ���g���s���%�x�/�U���{K6��C�cQ�����0�r f�� �r�T+t�k���L[腋"����no��D����en,�]ц�>]y��"u�?��������'���=C;����Ew%�3V[z�vO��+b��{��V'��$K^dh���
�B��=�,Wt{M �Z`>d���{�M⺝ۭǃ���\�����q��q�Q�t�9��
d8�8���mٌ�4��HKh�:�������7���s�v��aRÐ!�AoWGd�m����цE���	˧v���L�T���n+i��7� \7ꑋ��m��N2�µ=��]n`-�,��W�\yR۷��W(�Fh��o"��Gh�x�V@I�rj��&�iC�5+�qp���9*d��c�4nT�r��
��S)���[U���X�����Κ�U�8ɡya@�wN95W$#F�@��𝤴��W�咀���G��?	��N����ڃ���8�i���U����|��C������S1���|�!�`FQ�{� �}�\�^�|b��-}Δ~���m%����|
G1l��׉ G����J��L��_&+�Z��=;����$^x���0)���A����:b��j���^<M���9����x������i���SӘ���KlTW<�2��
m]�b���A�߫NjohX��'�޽^��RG|���38�̄3���x�jf�!�3�t�5���뻰{�y����)��YJ� ��&�{R�j�]++N�Wn� ��%�H�,v�G������*u�2J��M��cXZ:u������jG4Y���+#�r�>8sEr�N$P_v�3��3@���[��o��c���	vT�vx��3�������9��z[�ȋ��yf�b򟕥RK�o��:�I�[���r?oE�n��t��Q�^0BQ��]�Q"��nE�ER26��*�f���h&B�8�򬾅��%�N�ʈ�C�
�e3WWk{�-��f�`6X��Dׂ�o�s�e��>Q����Ͳ�\9]D� u�(�f�F�����V��0_��t�ze3��l�ds�K��vU���W
��,{�؛���e��k0tE�b.@�;I�'�Ng�ʁC��������w��S��{�݃����Q��E�T^�'��h��"0�"m	�`ꝣ"0+�5�� `��֣n�"����x�_s0�Q|�na��%�:؋b�4AdO$h옙[M��i�>͟xv�U4�`�-�{5\�\G���V-�z� �c��1�\�S���#�F��b���w�3�z=~�W�^�b�*�U�{~MH0��&�m�G<�o�Y&}��*qp���n]%Ivڙ���{l)�11#������Gd�l��h��]8��=���}B����i�W�Vn~��p�G:<n�]��f���"�);}~˹w#����m�a]��^ֳ�c�O%e�\�]L������k��-x����uu�q˾YS+�4��vIz��Z����򦯢�l�����N��}>rh<�"v�w�o��8zG@R��U���7#��{��l��6 BÑԧIl�w�Qp�){c��Q�_���ŕqP�&`�KCbsm�S��1J/Ȣwl�9�+�=4J�����Q^�t_�2�A�T�ȧѵd<�̤�>�^�L��Mސ�ϼ�ܲjg�l����S�D\g�̦ODu��f]&�����Mڶ��,�	��WM���J�[�/V#M���]e���S�|u����˾%�Q\N͈��C&�S̾�����z톬(���;��I�N�:	`�w�(�����#���!ە�v�$��t��F*Pl��{exN�����`�C��x,=�Ƨ.GI����^��c�(`�K^	�>|��)��ۏ^��FC�G8&�>�6ϝbf����8O�*_�i�t.^�'�;��wI�9wQ*��$\OJ�W^B�����\�+J����z=��s+hk�Y��ނ�)V�~'�Y�״;�l��+E���s5�d�+��:Ե��&5ʇ�i�I��u�g\��a#=�)��伹�L@�ffU��%J왰�Ρܧ���YVi���/��\b9b��[��Ҋ�ͬD�����͝z2K��(�`�Y�v��K��}�[�O۹��Ð�N���N(�Z4�# XRxO}�'��H�H������+މ";O�U���N�t��EͭB�b��l�.rgyY7Y���
d��+��" &z�7+�M�-+�,�a��p�B�q�C�f�oA\��9ŗ6�aM�#<H���e*�vőm��)�����pc���#c������u0�9�"��;4[ c�B�b��vd�Ǒ���N����+�Z��Q)�϶��슕�2,K�����(��(�rwsq
f��&ޮ��qZٍ��T��ک�^��j�ez�����κ�UN[���띙��4��A�u٫��:��+/��}�����Чg��w��U�N߸������;���M�6��#�`���y[�&K�m�p<�A��΋y ���`�W�2��W�V���u�<.��T�⾺@��ł�	�}a⩮e��*5�MW�\ޕ����'\ʌ�t�{b�G�X��<��:��%��هB�Ǘ�䨄6@��<���W\�`5�n�w���"�D^ �O�)���ȍ�V��[0v�V)Һ�!�����Ud��<Ռb�j����O(����j`��N��t��Z�����:�'n���,�P��ՠj��y��SH5��oe[��x��L�� D+�gY�2���.����t{$Y�.����e��*�n�Ի1K���k.��vj��lˁ[J��f�u臈:P,���-g��� )%��ͪ���# х�mi���������q�<+�Ϻ@��`ą]q�ᔓ��<D����r��:�W��uа�(�<ITdy�
`�{n�K*��sUh�Ѻ6q�5H�ܭ,s�dm������cm;����� �MU���z��?UD�ˍ����9e�iX��q�Y!����k�{Ћ��qS�HK�0�H����-κ��M��U��n�{�����>+6v5Jv�	�-.F@��	˧�<P��+�%�A�l���l��l�?I]�B���(w^�R.���d��^�����"�{�4��u3�n
��!&"{�'aɡEq�*.��T���S%��.�3��s0�n%��սz�"�q�t�d�xA��/�)gMl*�^��Q��ړ���i���J��pb�/sN�*�$��#��׀����}�j�:���ꍨ:Su�l�\Z<;��]i��QBΉ�o����.�ʞ��B�ܕ�o%*)IV��m���Ê��R�
� �@�S���c�6_5�Ջ(u�ݿ���1QꜦ��x����ͮ�GB�6,�P롳iw	p�B�e?����'��q��X�Qo��9ڕ]=���!��`�0��qR��7;u��.�G�Qp6�۸�/fr�p:$r�2|�FD���m��tħ���1�13~����2�|��eo���'c4�"�١�0\�;����$4�t�Ub�1A��g��Xt��^~����R�-L�;��� �z�2�J��G��ݎih�����"3(�q>W5�OHg�À��z�{K��UI���/pKO�J�]����	�4~�[�.cZeC���W�"pW���0;�Kc�,F7&��b㈹���y����a�(�zg	Y~��*cl�$�$�,�4k�^���s�Zᇭe�eՎ՘Um�P�#U=84��Ǵ!:T��;�:�����N�A�u�v�y�>��Wqw���v|�H(�k5I+|s��/�i�[�
,��y�9�@]�W�of�����㊜�Yԣ���K�:��;3��S����un��F�J�eT�.e���u��v�+Ȭ(�@�����'VϽg�{����J\j��:Ԯ����}kG��J+l����ZQL�tRʩ[�{��޵t�$�σ��.��L�aOV�C&�/]REJJ��a�O:׷�0���[.���'���(]	�2zN�G.�\Gd'�\ _S��D���ڣ銔��;9bi'{(D�ާuļp��jT7�������f�;�K��[���(�ŕ�zb7_YB�;8凕-�],��S�op��1Jn�X��e�����8��{@"��o�@�C��M�	�:OQ�0��Lu���a�or����d��ߎ`Ms�3u� T�-�|3���al���F�#r�H-�����.�*�ב���Y�KAe9�wܶ���]�A���Qv,�Q�5p%Vf�Sʊ�
:��;�,��y��w�k�5��1d~o�R�݇oZ��R�S�N���[��gY�y�oI����&`mӈsR���k6��.AR 5p��3pW��J��b خ��>3a����]��c��԰K���M�q�Ys���zhr=Ɔunq�������+9U�MVG������a%fҖ(���)ц��)p��WSR���i�N�v��#��N$���	�3����1}��7�l�j.s�@�F6.�v�e{���hC���m����� �J�]*6n&���=U�vg78�.�Vuv;�}�;;�N��mҭo�f���'q0��F�:��,b�B�"�U�*٫_B���p������R8�V/�>��u�/���n��^��k*ZEb=z�[���!U�B�ޮ�v��ެ����S��Z�U��ƍ�be���[����D�@v�.�W��J�Y���l�X���V�t�p;��¯8]rv̧g��"޷A���/;{/j��I+��p��Ӆ%�e�����b�榼���h��m�Kq��[y.f���`'#}�|WE�"՞rf8Ջ}G�	2�Z%-��_j刍OI �� �#b,�zf4�o�պft��y�3s'�)�B��FZ�|qm����঺��p�E��u���kkn�8Q-Ŋ]��4�r�w������������ƺ�^��A���[�M�-�iffܩ��M�u��s'c:�5݋�������Rv�6�=&���,�����-A�`�� �r5n��[�.��ŏv�DKq�{l,�{*unt��݆K�H��q�W4��b3�Ŝ\c���9�y=�����nD���q�<�mX����}W�É
\�G�$�C���r^W ��g]Z���]�QA��� ��[�ϳyJ��
B���X���8 �M㋦��zy�T=2��+0���5�7rY�s4'Ь4�J:	��D��T�7Qt8l)�na�0��)��bъ�ḫ�[�ժJ�a�g���9��>������bR��,#��T���1�o;�mڦj�DEY �֛tE�����R�U0�N���x��Z�ֆ�wyD�/�f�<�Ż:�7�v1�ΩT_�hւ-ZGHi�5l�DA�Ѥѭ�h���h�э�
-�[�حQ�d�h�M:J�UPkcQ�*�1�DZ4EQEA�u�A��[j'm��i��m��QIm�:5X����I�)�j����A��"�&�Ѣ"��mF̓TUUl��bZ4�)� )u���mUh(��8��EllCEhh�mb�P�KF��kF�"	�d֋F��)��V�5F"$�����֝�Mm�'C����UV�ڶ	�ق]�L��L[cmDU�Ӣص��6ɬTF�f�5�0TE��h5�����D;i*5���1���
��Zժ���F"��QE��������5��"�lf�Elj
֦)��QNH�m������EP[�C���`�F΍����"�"����cAII4����&������*`���M����t�.�Di\�[�5�o"�	T�^�Ý�xjS�p���ܹ��.���O�:Z�x�d/*t�Cz�A4*�ŧ��5�׼��w�tF�������Ӹ���'w�r���'"�G�r�m��>ߠ�����BW��?{���{��|{�ʏ�w�~��u	y�%�y��T�t�h�?y�K��|�@��n>������|��[��2{�b��{�C�{/#����:���`�{�S�i-�ۓ@z~�*B��0r����a4��I�{q�~����~���s���ϐ�O���~y$n�[�s��~�Z����`��@�R=^GR�_C�y�w?��ϰ�7��`ӥ��_7�C�z<��ߘM<���;�˫�)/��K��=�Oo1�N�B����?��>û�y�����<k&�˼����>���",D�O<�O�~�O��{���J���8C�4��7?��#�r���x��ri4~���x=�����=W̼�C�����r_��v�}��#_>������Ӫ
�3��Uu��Ǽ`z⧟r�O*B���C�?��}�w���\Z|��䝟�|��!)�O�����/ �%}��]-�Pr{���rӧ��>>{��K�9!���̼��9�qx#�dy�w]�W�3�]8����Lu!/1�Ov:��.��;8c��nO�tv~�����y�>�d�>A�e��뾍�	��w��;�}�G�J~�~���a�rh~{���(y�����f����kf��Ut\X���1��<���'q�?c�|����rNG��p:��|��ۗ�>��K�u����y��p<�?e���>�����4�wg��{�B��4||�]/�>�4�G�p���Qǽ�{��d������#����O|���.��~�}<��~�������Pu��9>���`���J|����sϐw	T��>A�?`��9�`�r����i����wx��Vs�}��k-���C�4�w�C�{���<���Ƅ������>{���~�G���>�s�]'���_�z�T����<��7��S�?nO|�S��S�~x�;���#艊^K~�����7{.O��>���~���^e�O���C�e�r_�g��y���߼�	T{.����p?A�/�O��8*|�K�����r�����\��ʎ�����_�}_3�.�X^���ߝB3�j�	x{8���82���`G-�JT��Ү�77����nK[�i黣'L-�]Q�r�.��?j�(�fp���@�T�Z�2���R0pR���ns)��k��.%���=��hp�fL�כi�-\��4HWʭ�ú��.��+��i��׼u�_/c�J���%�a�����8�BP��/�tϒ�d>s�i�䜏���_=��u>G�r<���8{�J����:�'�9!ߛ��hk�{�=��*;>��̺��g~�����4��Ù����� A�s���G�]q��~�����??y�� w��%C����	A�_���~��"0CM��i[�:y����g�����z� �%��4?��t����y#��vs=@{M'[�?_��<�G|ǰ�y/��?|��;�������:>��tQ�u�:_gO�t����[?|��#�#sqxQ��[s�5�
�m���>C���=ǧ<�a4��.�{��>��J}����N^��h(
(?������-::9�����^G �s'��y���9ǸJK��{c� �Du�I5%�w���aU��yS�]'�����=�˓�'�������y�ބ���|���s�&���0u�^^GP�N�l>\��(J���0w?��a���#�NG���Μkޞeo�����,�IOM[�@��䜏￸�(=��z�$�K��z��C^ǲ���z�w?e����y�!��N��^�;����<�G%��0����r�������S�¾�����_J�
��=V)�M!�C�>� ����O�O ��ߺ������O��{��{��4>���{�:���9�������h�y^K�y�p����$|{ި�*eL^{��]���%�@w	y������~ˠ;z���/��Ժ��=�~��y=���/P�?�!�߽�;�	��~{��Q�J���$�>I˸9��x=@QA��y��}��~�R&��t4�6�aj�d}��.��r=?��y��d���BS�;�=��K�׽���~u���=����>�����������%�k��=�~Gΰ�~>sޗl�]U�_CŊq~����x��=�?Ue�/������r���{��w0}���rNG���}��)���n�A�!(�����O�rO��q:�����~�pƟ��>��~K�}�M�>ߙ�*
�>G�o�x�R2�X+��lq{Q��{^گ�{7+�rz�ғ���Cv�tB�Ӵ����7�R�QW�2{���u�C��,v'Jm�{z� ���طe;RkoT��:�d0���ɝ�[74��]q�<��p��dҦ��T�oM^�F\]�9}�������>����w_.w���\)�]C��u|��RSܺ���>Gru&�;>��>G#�}��n|�i�g���?����)���~�s��ǽ�n}Q���ڷ�Ȕ'uΟ�������x,#� LW=���1��뮓���/!�|?yø=�W�|�}��C��.o��O���K��<��藓���c�}�s/��l�����"L1Xc�#�>k�Q�eW�f�]������׻�N��䇯;�S�G$��G�p�Z(?}��;�����{�װ��^G?��&��r��<��w	TG���;�������ʟ��鈆"�H��>��f�n�y���۞/���_�zluT������G>�5�ǒ���GP~?���>˶/�������s�y��付������$�~�����%?��=��: p����b������}j{�W�?a�$�����}�����vs'PF��Q���y�k��:��v�����Q�����u=ˣ�|��s޾IIN�]�����w'�j����z�{�@�G�_U�9�S�&U����w��;���O�>ǧ:��?G!(���A�{���9'rj�A����4%�`�\���^�<�?�ԝG������pra��^��p����`��>��u�1%W����)�~��Q�/�������tܿ���y�(}��μ�|���M>_M��Ԝ�#���y?��rN^Og7P�KE��?A�K̝����y/��r�@���|}�=�Cg�&��5[^~�����~�pr�߿qz��9����c�yS�'����4h�_��q�^���?�=�|��!C��/��9�C��u:]��_������\L@����� #�Pp�n
�]�SYI��7�D^&=q�}��ǁ�(<&��|��)�<�zM�� >>�ê�a��?���=�N�~�ߞ�����i�?��w�>K�z����z�si 8} D}����hә]^���}����t�?����~����h��rOd���(|���;���C��&��}��z~A��!/��~A�<�g�9�*O�i=�{P�X~q�<#���� �@ͳ;v��u'�Y��x���^�8'F\Jubi���K;-��&^�DG���w.��3�R��1j:*���h&�A��sr�:*VtK{F������Q�ִ��ru<��1��i�Ӊ�xŽv��H�V�w|
�m�ܮ�KfK��thʵÕ�����`L8��=�����:���c��A�:z�<�K�:���Ǽ�GD�Ο��!��_�u��T��������o0�>������NO��>����y�����n�U��!Ǫn%�{�ue��� �~�u��%�A����_�;=GP���O��_�������8K������c����~���pF�e���|�������/q�HP~��	���~�u�*�Kn���G�0'�w�z�e�/��u�J{�l}��sBU_�r9���n�:�i�>�χ8{������;��?��{�ʟa��:��}�����|?���1QMW�0.�����T{�  ǚs��Լ���ރ����ﻐ��/۞���u=ˣ�>���䔔�?O!�9��M�R>G�r;�;��
�����(�xQ�^z~�~��\_�i��S3�1�ܮ���QC�P���d�G�(+°i��jE+z�e�C�w�M����`u��x��پ�W�S!���g����;���U�{����gl�irpl�*]+~���b�(��K(��޽k��V��E��nIy�`��]�5y�E��2
�t����@]����^�����_0< ��*��A�ޟ�������j���۝���;�`�r�f�{���Ɔ|mUUΏ���s���<(��Y �Y��������G���q/R�
�Bt��϶�*,$�#|n����<�~Wzwcُ-\Ő�Qқ]I���B۞�����7��͋��S���u7b����JB��z��o=��&6�G��
��ۧ���5�f�[V�?cr����Sv�wU��E":ip��U
o�<f������;;����;5�9]9��(��l�N���y�QU�o��>p���L��8앗ЄY!FA'7ٝv.�!�	��~��o}Nf�� �I��5^I[��|sO�m}c��a��
�j�w���u�G0N2��� �D����h�?]mW#)O�JGE���N��0���ש��Vd'�j��j:�|tF�r|iA u���'�N`�*bu�рKj�p�eF����Ƌ�q˰��Β�����F��D"���చ;����\�.��l�0f�59輓��s�ncj�v�T�!��&�u�;���b�+iѿQ\v�;L���C͌	b4U:���_x(\�G�uB��N��*@8X3��M��TL�����ґdMC�\�,K�5���h����=�Zj�W�Ox�e{�`o�y��i�oUq�"|_Z�;ԫX�^�o���
�y��~v����d-:��-��#O���y,D�z@H����?�Ӈs����]]�U�[��*�½f�g<&�^.�bb�>���GJbo:��"F�ܘ�9bJ��F�sm����� 
եL���G�������*̃�� �Q2U��V��y=|�/)��
��� ��l�x�vķع_&d�v�27�}S��x�/xn�~�3�v�i�њV�;��Ȥ�[�`|�3�EO�/"?���sOܵ��W�?R����[���6F}찐�?nW���V
�� *>�UO�lI"Ez�}&V��[kЦ���T�H�f7O ���2�.�K!����4{��8�s3��N6�=V�Ʋ���b��C[�f����k�M,��z%^�F����>K�����V6[�x���-+)��-܀��2�+��^�2�^_�u�=v�Յ���;$�46�c*���9<|Z��A/���U>���������NC�;�z�{*/���|�b�΄{'lp\�E}󈃮�����Z�J����R*bv��Õ�.!��x�S��۷�v�|� �0���	:��;��|��͑����z��xX^�V_$O��-�o�mfZ�Nc�*:��|d�G���B$�ZM�̬�k� �9"���u7z��ۮ�,���3��i2��G��H�� �W�4�`�S�S36ޙ<'�Z��arÚ��l�ފ���G����������$�ړ�9+˸���9�;��O6Hz.���2�Ʈ�nc��8&�\m|ut��+�u.Ǻ*3Pw���+��z���"�׈9��H��;X��3e"����B0k��@)[[��6�gk�Q|�\At����ɥ$�Շ��f��X�p�U]��S��=��;�ƛ�c�D}N�#xظ�z���To��1� �"V��`>O����-�������K���Ӟ�5ʼt<6�?�a��A�=$rN�n@���#�4Ļ�ԊhJ�ah�=m����<EmVt�Vj��x���ᕛw��U"8z�\g���Έ�5ˈ�IH5�L,��5%�Ϋ=�	������Q����D_'�1�Rz��f�9)0���B&��f7d.���iw��[m.7-_K�2*]-�ݾ� ����h�8<��D��pp��*���}��׫�*D�0_��n�x=�q�v@����<�%�F��W�s��n��W�"/���Q�y3G�3��o�KE���t�3bQ|ǵ]V%�t곏"��W\�a�#u����c�v�Y�r%>a'.l��A�@@��e�נΕ旅:�|��P�X��	��Ek��Y�N�o�n��]�}���!��54Ӯ�k��hT~�upD��6|+�S�WoDG^f�Kbk���`:]!]�&����� ؇��W��8���z�����3W��>;�!�۫FK���:yR�Ӑ��8�,Ӽ4��\e�:*�Gu�t0U��øy�5!+��a�N\��%6ֺ7C4J��װ�%�qhH��㜷/鯏m���N��Ym*�b]&$8�s���W]Y(��J���
��G�ɤ�u�Ц�{sS��p�E#��<���s�dm㨅����	��؃d�
b#zjJ�����dl�����lq�~���	U��ڱD��<�;Jf on�e�uhթ�0$̵o�V�͒��޻�!^� %v���{�EJ�]��kѹ�N�#	�-d\6�M�me�N;x��W������,�g���b!W��j,R����{(r�p�j�1U:x�1~^2��91����`/\ߪ	�o��:	�� �C���"k��;��s*������mnK�E�1�Y>~�ԉy�r�5����Jt�(��3��	魅��k-� �nY8�1��unˎ�Iz�{�Uɱ�@B����xt����H�d��-8ɸK���X{�uo2P-�m���+�q|�lnT��;�8��C�~���m�����ٜ�C��A�o6�SY�H��)�$��}s>�Qy��K��ޔ�m*�2�|��c�۵�+(o���\��K0�Z���ԙy�%���v��r��eì�Ѳ�KQ|�	ʵ7�h����T�Yt��B<S��1�K��t���(�5h^[Ƈi���|}��}��a\ޛC^T�`�l���i����d�����MNb�~§u�s�v�`��*�=������\�3B��p��x���^!�lu�l��->&�ۏ�u3�u�~o�T��j�V� z�/zwj{�-�zy��^���ƀ�tUp_
�����/��W�l�2Ų�jWf�sݬ5���=��Ae�^�W#��[���ɝ<,�{����Ɏ9] v���ڞ㾄��*��C9I�Jw!z���UZ�|��λm���'U#�/��KX��Rkݛ�-��'dh��s��s��c���"åN;%e�,����;�A^��h?7w�������+�\{P�U2ϫjADw��V���|s�|���5�h{��FVp1�^^�#��m2Z#"I���D4��+��8)��GG��*�=�F�U�}����`Z����=��/U���P��u�@�H1�HV��i��S�Kk����p$�ݯz=Jd���l��4>�L��"�0!p:H<��F��h$�ÍK�o�%�j6m��".��n3źD�����Av�J�� q��0�c�.����]%�o��R���z�����N�L,5�S*ts5 ��˹J۾M����87��2qK_{���I��X� �^�dT�L��u�e��`s��J����+��!����jٖ�>����}[�j��T����
����X&�ЂvE4�X�:�����?}�� ��ʞ'p����w�(��Hrv9*�W�
���uW[7�?P!3�\�|����K�v�c�����*�N��7��7�/�]$u�D���9T2V�����a(X�|;�o��Ӥqz�^�k����~���v�.W]jwh���My��C���Q�Fy��]��Nrʝ/���~DDp�`#!W�xr:��#@͕�٨�qiS��g#�. \�3�Ɏ�W���芳f%����g�v}a!\~ܯ1�@u��g��v�7��̛�N����~�2�Aj^��棸����u1w��ݰd,4U����1sg�ON�r�m�K�q����#�!�5f/�N�d��{<���?O-��X)���E������s���̆����j��u�ٖ!\�E2��yF��nߚ���t䝈|7Q�>�����]�y����H~'�;$����UES�F*PaD#�y�L������Z=~[�r8:0Q¬�| �#�;:=�t���ă��V���z��_���@Ň�E��Z���t������n�ۥɃ����LYw#=�vU�U���v��9'��t.�j��m\���ڣ�Kqo�7�%���:�Pr;fS�����(��|u�	L.)�qW�lԦs����r��(N[˅���>Na��."iX�;s{sN��Duќ�9G[A;o[FU�wv���[˹Q5L��+V���� �iz�9eϔլ]��K�T�'�L�*V�<���X8)��'9�ܮ\r�����J��x�䪽:FG.��㘚�S�z��n�]�v��jNc��,�X���V�Ђ�W(��gT��J^Ҙ�Vm�Xw�r������ϰ[ъ*����&��K!6x�5�H����ԫKj�A+�2n]mdqm���[��"�5}��QgmHE7q�v~T>�}��t�O0+פ�RN{�|��8_4UkZpD]]��.�0]���ls� �ݘr7t��b��Φ鸉Z��}�=�h�S��j���i��2�d���o�nS�3�@��5m�_v��Z���sxX�/9,�}l^|��]��N�4��iZ�P7.�YĽ�a�Ch�ܺ��@���u�l�XN�Wc��H��D�����7][y��NF��y�֦�ػa�Y�C�6��=�� ���l�Qa��٫qÖH7�.	�b�dY����vqxF���t�>}PUĳ�S�Y�-h�H!��䱦`=d����l�Ws���x9��w8��1naT�zm��U<���LG{z���7}Zt)ch�XZ��j�]/�f�2�����k�x�/����W�Lͽ�&E��&g8���u��Z�XĮ��s^S#��r���嶭q�k�
�e���
x�=�n���̓j����Z2-��qp�i�<�L�o,�u�B�j𥗪l.�e�3��K��zc�Va����e��:YK��Q��)b�
�M���c7P��\Sã���ʂHV�c9�ɨ�>�[��j,����w_)Q�*fҕ�ݭtd5��^Z�S�ntlz��Eӳ�H�Y��#A�y������.q�Cړ���(���|�W}]V����6��J���rA���;���u�]��E��	}��=��&�SH^teq�B�p�S�L-IL��!6�M�)�!� T��3��sr{�3k.$�H%�k������A���Z"�o
�+�Z�1�t�kv[»�U�j{�x,��no<��{��E ���:��F޻O����SԾ�٤0c�H���r��d�֫�(Ż�)��펧��NH��.���9sμ�����+���#����v�/v��X�}i/�:��O����)=�î�X��Df��$�qmŮ"$�+�z��J��%Kzr
��>[MjJ�v���Q��4��1���L��U�!WF����+�J�5�4!$�8R1��������ѝ���������
qT�ƴE!A4�TEUSF�����֨����:"(�USAMP�UUT�4��PZ�؈����)�i����֦*(�b�����l��v5SF�ӭU45V��EM3I�UlgZ��j �ґV���X�D�E�6���+C��ű���8��������
�
���( �Ѫ���A$�M��Sh�$�UD�LEiuF�EQED��[h��vӳ�h�g1CRLE�Z�N��U5%1Z5EU����*�Z��ө�&h������
Ӫf(b4fjjh�������EMS55UF�� �&(��*�b*I#m�SSM� �a�QEE1�UT�DSEE�KULUUUU�!����&��l�(��� �1TUUm�������5Z0Q-TTV���;�>���uSF�ͅ�o��SQ���/)q���S{Q���$`�I���K�����3>�e��^v�L�%0M%?����uy�v0�"8����;�X�B�$��Ep
��C��]�V��z>�Ї���焼tT!����H�Q�����c�q�p�N݆,�G��!��I�̬����a��{�fO����M�v:/��>:��i(c��䨜�*k�D"$@�E�l ��@�,���x�d��-�W�'I.rg<^;}���'��
<I<�r����cܔ�YV��" �ǠW��9����<H���NG@q`��K�
�!Tf�L:ע������JWH��.�U�Z�>5�����4�a��hzUyhh�ԝ�9k�7��-�+k%7;��N0!P��ђpqd�FO���"����r��r�����8>�]�r��pgM�'��O�4��$�1�UR�'v2Gu�����0��ŵ�=4�Gu���wV4#{n2�՗:��y�>�<�OyS�q�N�t �k+����E*{o�ܹ��'S�#�=F�t��ݞf�o����\��uA�5,�e;S?XB�)�9(�����MP6�,ם%������)XBtg��U�$��'xrJ�Vy*�A��d�E��^k�(@����Da��!;��Z,�9�]IS'WT���V������ʬ�\���}AWkoZ���F��s��w�YS��0��E�� � GY[I7t�{t�NF�eV���(��������k���m�C���5=����];�nȲ�����F��KE�	}���6'�����:�eDf����]o�z,@6S�����)g���e�F��a���]n�����<#K���=xS�>���;ч&�`�)�g7F�j��ӞG����\BۙEYd&d=\;�g»�_!�S��;���۵�w�9���c5�
3�<����W]=%�%Q�!�h��HAs}���8.�vs|�v%����BS��f�_H�}�G�+���d�GH6B��l�ϻ��5ԛ��Zʬ��tʅǂ��Q.;�2v��@���f2�գCv�fRt��,U�:��o2����D����@<���1�k�kF�'��FoKG��-ID��jIg6i�z�{��/(�=��	U�D���_R<�j/Ԥ8�:\+q�W.�
E�&�a�\:sG3V���n�����v*�.\�h<�e�}�4�E�=��׽~UTɫX�v����Ă���^�OYMЏ���"q��F+*P��Wju��e��v�.l����^��<7r1�OG4�&Bw��L|��<Yz��x'��d��[�kd��w��Ӽ��o]�$w�Z�If�G�9�*��?@�����Oqc�st�ߢu"W�
P���'�U:x��f�C�kk:j�~�$%�zkA�g�W�r���@���55%z1������5~.ϢzY=B�� �{��zj�|�z�6r�����skoH۩����@s=A}��=i_����{�5�[����
���>�ƣ�sc�'��L߻m_�)����ekWbx�bS��bD����E�=\(�#`�n�p�-X�ճ�O��[��s=�^��5^;�c+��{��x1r⎰�f���zk�-��@7tUp��x[�ٔ_0�^|D^%G�o���F]ׁ
2�Vz3��6y��0�o+���ڞ6,�R�?Xu�Bt�V�&��Q�j���	,#� ^�5C�X�RE}�Jw�ۅU�=�]���p�G|\]��n��O�y��ܮ��7��G3���Y��ONǜ+yC�ҧ�V_B�8H��B�p_9u/*��Sk`���Ȁ�����}_=�m�6�}�}��g�>��=�o Tqq+cr{�i.�]4Y��C�8�H���=g �*=yI��J��^H;�5���֠�6��L��Cm&덊�.�P�	��,�]��k�N��/*� �[[����Ȱn
G�U�x-�:�K��aY96�GQ�c�ȃ,2Rţ{�<<<�kMwbrlw�����  +�:�����3-ό6v.��7ո�}��,�n��N�<��2��:�>��^��Ug�nA��v ճy�xE}�U��g��w��n�$�U}�p��F�u�M��t�gԈ�g�`B�'I'�u���T��ۛ�|Tė�٬����ܺ�������&�%X�+��l�ȑ�ˍ�`%�1�=m��X��wEmј�9Oz��(���%6�u? 0J�� ��ꜗ��+�[��W��hُ��� "�������w�Ѿ�\o�����2h�n�9�:�څ���W�6�s�J��J�p�K#Ǔ���O��Gl�uo�x;�U�^t�{��Dc��"dL�`��x���c�A?Wl�tzʇ4��E]��*�½f�g<&����(1��y��T�!�����0UmX~��8�{>8��*3ݙS�V'2|W�B��#^��D�l [A��N�own�x�D0��8�e��c�>r9����}���]����d��
�x�^ղV�.��d�{�]��b椯����	����슘u�M�l����Bb�ܻz��b���==٧�[8����%6�����pB�%��������[o���W�S\�]�����iǔ�y�R�2T�@&;Ý�[�gv[X+�F
���� W��+����!G�g��(��غ�_S��8���m5��x�Jc�[��KG�=XW��ױ�#;�X2�mҪ�}rF��,B��&��S/����3�3���It���sǷ���d�
�I0�8�L��`u��"��}��A���6�ʮC�*��	��+U:�+�_w�<+Nx�x�8��>��Z.�G���*`��v�noͤ.�����pT�_�q�j���U���\
4���*"}����.6]ЗF᩽�d�sA��Z���$<,(]�\cъG�4<�Tr��,Џ�B �ZLÌ;����1�nV�^QX�X�ݎ�u/�ru����-��<�'�Ɔ�:�<����Q��S�J��5�~���#��vh�������#�l�^ T�ʞ��i�(������*T�ٰH� CG�PV���)��$^��[�~	��,6�w*�>Nz��t.�ڻ$6�yB��S�Q0��4�J�udC����W�ei�o:�l�L��2_p�Rw�cO�va���۽�� [�[}q C����9��f#{kq�*4��T��Wi�}���=�ˎ�^8�Y��G�w,�f]u�h�r�fZ+��f����>��è�L��d=��IJ%Yɚ�U�8��w>%	L��K�1on{�p���S��{�	�6��Tc{w�Ə�\���*+eْhqD����.ȩ]C"ĩxj�rn2�յkK�iڊ���QѹS�ͪ��@t�G)@I��*��m�x�t-V�0��y]����>�}7�����2�VOWt��a3�J��������T9ٰ�Q�S0/�[`�x!Li�[ɟ2>7:�}O���lԌ��c�[;���z=&�S���wPr������.S��5�&�<��v9�+�"�W�U�u����*�'�S\�$Lc:�W�]T4�a���zs����M��b*�p��d���P�	����lJ/���ĸ�1�*�[ǁ|0ema
�ZL�V��wmq�i��`r�ƥa�p��[��������>�E`�56*��ӋDT<ok�C7ވ�
z�g��t>�d_AvT�P"珓2�(���3�}���kpRP�铘n?RWp8ku���$(��:�{a;��r��FIF�<IU�>bE��h�S��L4�t^�#�+�geؖf�iJ�f�:�Zq���N��E�L���&�&��Y^�cǝ�^P]��M�O1(�g.�kn��؅���Sa�pR�2�.M�kQT;wU��g�͏ ���G�%5�o���4��q�;^u�f3�k�����ⲷ�\H�Dw\q�N�a�w�)��PԎ�Ԭ#+������ ���Ul��A;̈���I����&3�U�㞤Չ�L��6�C��}�l��V���t#�5s�y�蕥���2�PFS twO��GD^��5�l����}�HǸl6�حxf������s�d�����J���(�U&Tl��<�j,R���+��9�-�B�6���nc*�c!���8	�V!ׄ�J�=I�29��F	;MQ\iV�yݺ�/\|Zݝ7�z�_�{��T��%L�qע�q�Љ�fw!э}�
0O�+��,.�4һ3b���]�-�&��f!�7.#K�Ɍg�z�N�����oGA"����9��qA�O�a��{Oq��U��+��V��@*6=E˄��s}º��J1fK�u/����{p�w�<szS6;m_�!�91\ʻ�R���5EqI�r���/Œ�f�:�����kJ$dY�RnH�&�m(��k���SX�О��^,�8g���P��wi�Ӌ�E����WiX��u�:ۉم��]6/EP����e��s��^���܈�i�iVj읚�w*1,1�}j1=��T��]��*�6g�3��Gxt�I�AgY����X��Wt�����)/���s9d쬱n4�8 ;�uv� pa�F�M�\���!�0ow�W]����� {�84ùظ��ySO=�<�}�t7��{�S�ŖJP}Q`��C�p�lˊ�ش�\N��(��MPB.��=ǒ��^�#mUhCG�v�C'�p��W����V���j�3��7MiAF�%vz9�ӃO�,{A2����[���r�p1\*,�Īu7�p�^�`	����L�-�Gյ ��bq�o�s�;Q�����Y��GHw�������c���O#gA�Wt�V�r2��t�tx}���7m�|�	�Ļc���K=-��p����@�tPTv �j��p�h��w�����c1��ܸ,y{�>�M���q6=��:l
4ϫȈFx���0(����zvF�ö�:5g�#��r�3A��DlW&�F�"E�\"h�lE�ǂo�GG���p!�+e�zLu���I�����A���7��(.QC/�M ����C�#�W7�ܺ������� �Y���f�|���@��=���T�v��J�|�߭5@�yd�&���#��5n_��u��ː�"��nۓ^�gN���z���/�����<6leP�k��r�q1��"Ʈ�����\j��+{mQE���T�罍�r�빵��N�b���`8LN5x�x^3Ё\}Jz�n�B�r�t�r)��'vX��;'ko�ʕm�W�nS�V"uUW�_UW���������%j�:�\>�c�UMm��9�P�AM;S�x��j�*��70E�un)�L�`��z��Y1����P�m��׬���	��\<��( �����쨘�|��|�8����y"�٪�n � ���v}a!\w+�f�c�q�{'F:[��Ԯł��l���X�9�ʟ9�sQ�py�W��wSc���`�XQI���� �GVZ:&�1�p{��sr2 ���B����a��6N9����j����gN���T۸7�!I���$�s��a�gh9S(�\�ѽ�b���)������@��v%��f�Ż���Lz���LD�D�s��X9�U���F��ۂ��3��q�5-I�f��%@�5~�]&w�x��ӕ�E-� �<�
��ף^}��em�]c�^;�Y�Ӥ�u�ݷԱb�>aӌ���MX}�V3�.�Iۢ��!�*�+r���{���hVg[vj��b��*\d_��4F�s�����v�<�d�hG��!��:n�N��)\��s �\�E��ﻋ���wa\h��:�T.v�MT�O��|��n���j(�[���Wl����k�gՐ֬��{s��3��Ӝ~�u�[��/Ue�%��sW��N� T]��{iZq���M��\�8fatql� c��W���}����˖���{�tp�X���u/M���i2�ʀ�|���+id;/(l����ێ^fDB!� ��WA��Y��q����C���� 6p��oɻ����.��I̭�Ar!G�ia�4{��" �L�
���fz6S7���S��9�mg�K�%��ռ]�>�Z�i9�;�|Hu],�[���U��f�Y��4<IY[4J��,����f2�2H�ޣG���]�&��:�Z��i��ub.^��_n���t�N�"���l/5��z��"��S@'."M�	]T���Nף$wX��>�nLWj��-co.�W.v�CǍYB㺩��AF$)��S+j�����Vw�͵o/zth��>��PWYI�2�aL��}n3�a�5�T�j����g�W���x^�b=3~���s���(�����}G��+KG|N�8��߶W��{��p1�:A������cX�^˼���0�#~�VFErp剞D���K�����ĸ�1�� �7��iZ�)	���[��mj��_to���(Ӝ:�?jX��=�U�ʔV�Tc%;�1]���u��M.��_lޭ1��{L�ݥt���-�u�h<X����Ȧ���Gu�����rX�ufi�j�^1N�����kqoۓ��L�)el�E]6g]3�7�r�Vs�`�5#��H���k�X����_w�:y��֩:��i��Hl��p���:9�v*�P���F��e4�����K S�6�D�˧�L���A�|�of88O�]�8��fp֝#���#� ����j�
�:j�:��kP�BѺ�9���ܫ\��e=��T��lUӔ�YY}.�mD�U�W[
2�,�
s �C�HkX�Ͼ��dZ��ۏ�\�n�뒁���=�9�Z��f�.\��E��N�t�o��q��׻��cl�I\��c�s��;=ϵm.��g=�*�,�}; �m�b�<��G@�om�JL7�Œ�-�0�V2mq�z��zt�e�u��%B�γp�c�.���7-ly���|8sg��Q$"��G�����ed�q'2��a�Ƃ���T�k��3s�gPI�:*=V�ب��F�Lnr��&L�n��$��vs��S��\��6tpsp��c6��Nc�]su���y�|^p��R�Y�AQ�Ea	�Ϟa�{��(�w ��c�)�^�Ň�~R<�1;Q���/V�Y}N���a���C�����l2��t�t�4������MJ��R��<Wu,΅�G�v�\��\�R`�k`�Å��Q�t6���gWgF^�[;� '�����sY9Zۋ3�CB�d�(l�Wp���m.�Y���<��:0��9S!unl@Y��V����gܠ��_`�-$	IQ�X�ҝؽմ�7kxS�r�{h��(��2�� )����u�+E�^)Orq9U��:�]m���Q���J�^uhv�gbGn	�8J�Vk��@"���V��5�,��ʂ'eure$��b����\�z�̃e�@���Ԟu�ZN�|��A˥��:Ş���/\xiWq��]W�ؤ�M�˩'{��tee�&�����8u�S���(��oGN[�ܱ٠��!ro1䧇%���r%�ݤ-f�.����Q�Z�O��[(��Ԯ�Grh��%Z�]�V_ۇ���n�3mkO>���tt2	AtԶC�6�|ﾶ�E�h;f��A��p��_x;�ՠ���i��{�����,yAu�˜���u�����N�a��uZʙÏ\uó��{f7έ�[��!�9�[�(8b�kR��%��>��;5y�f^�d�v����G�˹^�.��ɑX��b�ȯ
g\���<����y]IS��Y\	y���U��T�B�Q��ҔK����b�C���"��N�**�=z*wk��+B�$��QVa�c�,���/-�UN��_��}?��6�UMM��*Zu�(Ѧ�%����*"j(������m��UT�L�TM1EPV�Y��*�b�bI�"J
b�*�$��gTTDI%1RMCUUMcm[�]5DUS4S5�QD��SDV��j&������f�����TMSUQUDDU��b ��cDDUMEQTUI��3li�"*��(����!�j֨����
��"�"��
"�(���&J�
*њ��CQC�����ZL�UEUUD�3A54��SE4�3Q�EE豊""�""	��f���������j6�1MD�T��QT�bb!�����h�b(��Ѫ�
��D�S�UULE���"h��&b�6��4�q�橀������ϸ;	�Ѝ��W��V��զ�@=��j�:�09�˕���Qv��]|P��ʹdu��)l���.����=���[[���)"��u��Qzk2w�q�Xl,W�n��G@�<#�p(�P�=�q�ɱ��������iljc��DW�Je�����xȾ4���*���U�����|�թb2��z���C�ǯt;�;<M�--��ke����w��]t,�d�_$�� �lP���2�;�b_�������^{��K3O��Os�dm�u�����Oޝ���;�I/$�rogm��^�@��G@C�R�[�=��һ�B\ˎ�nd8�8��şf�K�M��A����i��Y���E^�uҐ�;��@�:#Dv��ͭyRF=22��C+�-���:=JǇ��׻�Fg��x�9#��DV��"�jaq�	.g����Lur�<����3�������`�-�,�"�*�ׄ�*���*N�L�v"{�;N2�1#��b��\1Ҵ�a�t;��8��}^䩒�C�/@��Szx���dw�Q��دf�m�.�U0�q�ľ��ѓW���^�=��M�� !IJ
�æ����IP����qR����謕�6C�]�ʦ�w�֬XsU�ˤ�R�MX��h�8��*^dѦVq���\we�7��|�;�������W�t�8�9���r���h���=���}���wM�u�X���F��KUVfة���J.$v��������Y�����冏��]mf�˕ţ�����p���\�!�%����ʼ��z�~#��N�d~����j�xV����������Wx��x��W��<���J>���L��'�x���
6�8
[�e�W��M���#�3P[t^E^o1'�����j����܊�+q��EW���Ӊ٘\�W���Ҫ֛�>��0h
�^�/ir��ʩ#������omO��JV��r�[0�����9��ٵ��l���;�����q����1Jn{@yN_��n	Y~��*ctKLm�Kb��ӕ�i�8��O��FUz���`!��Y���i���dXt��Q���$���Ww~����&���ih{h+�L��R��Q4V��9�_&P�H�R�9B
�E��An{b_�������T�GAD�O?���?\WU&r��Yt����=��'HJ�*6��;��cO_�\{)�_������Tv��y�ګ�f���;�ܴ�{D�Ws�6�*���P��@��QTB�c��{2F�!yٱ,�e�UWUm��c2�s�sPؘ3�L��ɠpi"�K���A�}��x�IEoq.��y�*&�쇦��e։�
��J{`(�}�Y�-[�\ҿUUP���7Ю�'�W�P>ԩGAMP�z1�]��݃���>P!���t�<��yB�RԬ��=~�9�.����n �Q���x�\L\@B�P�� �v'H,��q��i�rȨ���I��=G(�;V7��)r�|�2kɺ�/!� `���z��ڹ�Kl�\��������`��~�}�Ô�x�3uv��[�>�c��&��p����abǈ��;����UBJ�Ux�f���;�R�qY���ya@�§�j1����m��QV��9�O%����l����2���U���z͍|���Cɲ'���G�h�ݝJ�A~���약=��ςڮEY��@� l�ϻ*a=�Ç:BӶ/�Hv	E�������n*r)z�09�Gq����컩���N�q˒��A�e����7�J��3 �W�܌���OdHq#�u����6N>��~MW@��+�k���a�2{����F��lOR[d��N�rGIb���S/����`��)Ⱥ�rC�T�VٝSs6\1_o!f�.���}89�1c]⳻}��Ĉ��B�}�Cq�)c�\��׶�sZ;�3"�xZ�K��O�!�Z�NX���dNT��[�Tq��l�������]��]�y8�<��ә�j5{<Q�ɻ߇�=�x5��JB˹��ΰ~��Z8M_���������#Y|��B��+�~����=��\����/��X�����������(xW	T��������1��3�7ed�۱�X�����E�\B;A5a�����Q(�'�* Gq1 !�&'[��|3u�TX��Yס	H���}����.�ztY1���glp[L�O
jv�BUg�!�}QKE����O�M�v:,���3��Ѥʿ*��<��z/r3r��5�we��/q Y��]��iy�LƗu{���.rg��7vmR�+8��a����ٮ��X�Q�$��K��& 09Ga�~�����t��wC� mʂ�\�Mz$~�a��u.��6�X*Ȅe�A�@̎w��Ƞ�W�xm��=e����Ԋ�w�Os7�ΘO�EIN�	��Ш`���.���Ϟߍ�Eߦd;Z��^���c{2s�fͦ9:5�)��h58��׭�1���~IzX���
�6u�`pĄ���R�x=���G�v���ũc�F.��[����z���es��2�k�K�]��Cn��n��D�zR�K�w��S�=7.�m��Pr�K�6���©�|Ư�9�q��I���]��u|�iN�A^����,]j��������S��w_�uf�k��h^մ��ZÚyNv���M1Om^u��^����^��Vj�W�M��kc�n�s��^�'���Q����u�;�
[��#���W�k���8��ʰ����u�! v>w�3��l(N����\�P,�n��e<w��Ʒ�|��eY�������sJ��PLn�]�4u��t_W,^�/Y�&�,��9��cf�˶�A�!�G�AΨ��߬_��ff�\9-�9C9��������5��}n��|����v�w����%{0�7�Љ1{�mWK�IR�n�ce�i4��W��Y��ѩ):*�~��7S�<U�^W����'�_����)<�sm�j�Fdjr�Q��}�ӊ���q����/wn���)�[�qO����`������m�M=C��Ky�P�4�.���}���И:s����~Q�]1p�y�����E�G*�o�~�~�G=��%�x�-�h���e��W����y���vK�'ep��Ce��=Sk��3^v[��9]8]��@(��XP�#k�	���#Uv����kUzn���Hgq�=�������eT��)\E�� �;AN��ɂ��>�;|�C��$/%R5Gi����['�X5�L��TI��˅nv,�}_.��-
��A���Q����޸�fN���IN=�����X�tUK�ܚ��Z�m���N���	Б�7��3��bOa��8���U[6�+;�4�{N{�5F�0�����<�Ψ��ƺ;�S"ڷ�-�֌��[��~�r��w�����`C�g������.$��O�%<�t{�<�ߩ��}g�m.�>[Sy�5I�����Z��:��Kc��jI�|vk��9'�s��וٺ�2�S�&�(�q�GeO�3�2_,[hY�wk�3ޣ]��v$�󚴅��-��*�9�w!�}�S�f_R)��L�n1	�]_7R��m���v�N;�Vŧ�$��U:f���<w6�J��Z��Pě���î{`|��V�^C�-Y�̳�fG3��t�]�gaV��W���-���#���ʯo  ���z�f���!��_?(8GV�3B�U��Ə\/�z���|P�������+z��w9�:��]���'���ꔦ��V�����wrRe7u��yj�aeq�߀��</U�����}��%p�w%��h�%J�[��Yc}ko:�t��-�EU�cW;��ZV���p��P�ʤ��O�=��6w�΂�37�ҥ�+~�е�lmߢ�J��/wFCK��Ԟq�Բp��ږ�m�nS�kZ�b�m�S�HT,��1��}���j�J����_TO�bv�'���ޭ��b����qS�]i٬����]���9�;�'._�y���ѕ������|+䗢��D��{(xٖ���ݙ�4z�+j务��^��5�μ�Fr�y7��CcF��٧�T�:!��Ԏn�ˎ�;����k՝��t痻݁!����4B�'�<�ޯr���.�=}�_���s,�����D��������$��%vC5^�;�S�u��9x���V�6�r����s�Hk8o��6����b��Y:��6�{]�f�ޅ��0g��{ _t��,9�N]wmΆU���nJHTb����fk	po��IVmݎ�;IL�)��;��I��N�oS�	�`Jn�;t5����d���8f�n���\P(�o������7,^�Ev���[����-c]�유�+��XΌ�嵗Wtba�3$qN��w+��鵵�2�ڄ�v�^�'�������D��-{N��:�6G�c�<���̉n:��غ(t�n0:��kw9H�Pd/t���Vԩ6wrΪ��B7�K��A��¡�W$�۲��w��8�8H�k�I�<�k]۟b5X����*�)������[�U.��gC�����=�U��+ElC������߽����t���;�����P���;*9r�Ԗ��݀o��X��t����"i�}��uMp_��M��R�E'�9�]�Xͫ}@'Mߢ��LW��c�J����,;�+�9��r��E����pOv+�ی��1Vs�v�S�eZ1�˰@���U�{k�FT}���V%�;èT�K�3m�fb��`VɓʽK�K�������u�n��	��'�v�]��v�]�i�贱w�G��^���V�e�p�/Գٙh?5赥"`��rf�F�xj��s���	R���ku��t l��4���ZY�y�Ig�L��}_W�x�
|;�\8�Ư��Dw����M	[�b5:����s�J�������յ�Em�z�¸
�V:�zxl����ܞ�5+};J�p\�b=��-��Q\�����M�8���аN�1<�E���\(M�f������Ln��sK^��>3��k�
h&������N8ڞ�BNV��Wn%�s冎ձ�����z�y⽫v���9���[�2N߭Y���Ӝm��Y��1m��i�	YC�:��s�2�,r|�E�`�,��gs3ݚ�wX�流��|�֖���.�Ê��q�k�/OK;���7����t�|uο:��]�9�VU���3(sz��P�A���XyNe����+���,�+�(��g3�=児�����r�<�Ow��ّ�g�o�P��{et,g�_�e>�o���U�˰ϧ"2��z%R5ܖJR���Ձ�&|�9�ַ�u��u��%��r;�Zb����vd�ȅ\�k�⯴k�����a��2ۻ�oy���G}8Ϋa�oV��5{�m�8p���������ֈ�V�4��t�xv�Z<��>��꯫��ʚj���Iݯm"�)]�-�a�Ƴ�i�*�j�!��×�7\��c��R{�����%(��<�sm����A:2��W�c���%����w�`^�"7r���r�o��`��~��.:�1bJ9��G��)�����o�9u��w�~z�9�	��CR��� ��Qʫ`��u��̄�^˦iR8.�#b�E��p�)�̮p���T�_����n�yt%�t|+����<r��3J8d���t
c1�T�pc�,�=�/u��Ԍ����5�aP�!�R��`�N�e�N'D�1�W>/r�-\׻��x�ɪ5�M6ƽ����֩���������8i�R����YK^>2�i�]�ػ Ѿ�^,�2LK�Mm_�H��C^�k����[������mU�-.j;slQ�x�;m��[Y���^޺/`�˔n�:��ģ������ѷ-" ��@�ń佾�]d�b���u)�������ɞb�]�S�g�ax�ߺo[$Yˮ�;��ea�X��bc�b�sl����̠��Fw2�S�].���,�V�9!���.5{���~Uۉ<Yn�ëM$��X��̫.(��7+uL��K]��	�d<�`�����8nƏ([E��jmotv���Y�qX�b�Ȏ�=��rW;�@KE�
�pE蚉�=ٮ<�u��\�'K5<�ٕ�Gq����V�-�{Ql��vmCdԖ���7:�L/j[A������Ԩ�qj�ْ�lˉ����-m��T���!;.jka�9J>�`t���Kǻ���렺i��(SW�)�fK҂�P���*ɜ�T�`V�t#c�7Z	,+D`Ԏ�+���'7 ���E�Z3��ޫG��=�Ԋ���GBs)j�G
�M��{��晨��7"�%��L��=���]_R����('��׵}�;��<�־�2�a{�%,OE^���>�x�n�iANTz���]Pr�������<瘗H����6y��B�h�Tx���f�!�\uw8a鳲��y��K5��̲)�עM�@��]qL극J�IX���)��3����#fȄ���Y�����e($*N�;�-֊=/o6t�ն�nYMb�5D�7/�`o�YTz���ѵѦ5W0N:��f".������Wf���gIE:�*��mF�z�hԲ�:�a��c�K&Νz��ٗ�����:�[L	�܊�jR�唒��s��s�2����i�������S%˓�P�}�x
�Eh�Zѻ��K����9�7f'�\� ��J:0����7�A��jM�Fc `ø�w7���rktpAy�`���76Rc:ݛ]V�!�CO@�R6'_@�N��+��F�j����j��o)֮�c�4���V�tw��%	y´
�!v@rzw�;̤ot�ײW3�QU���� n�m8�#3��	�8�vu<hA�wݧv��-2`i�ʻ�u�S���J�2K5ԃ��;�F�x�d!����VU��t=�wh��)�[���m�5\�����]����*���r�f���W'!�wU������r�a@�cX�\�����5'haE۝|�:����Bft���J����ݭy�?\*��̈́t[�c��v�v�$CYa�*f��\��#�=���{M�����������8ܧ�`�"
�	��հ�(��ߖ��=/��z�C,^k����vM��6j������AU� Xv��&�l�R4Nm�75�a��T�assr5��@F�#֖���T`(��f�+����v��� �C;���ǔ�>P]�Ѝ�*�jv`OOX�F����f���e��γz�sM[ܳ��z�
�� �5E�TUE�*&b#böԛj��v�[h*5�A�(-b*
���L�AA	��3�TTDZ�E,�je����"���(�������т��������*�"$����H����h"��
�*�&��� ���14EATb�������Tla*��*��`���������H���RUZ�F�"f��AkECEETU��S�d������d�RRL�AUZ4�@EU6؊(""��&��h��̑�0P��A�D��[b$�b����������j$�((�)�"�"Zj�X�QUQRU5$UMEAD�P�j�f�d�*�Jb��&��j*&�*��E4QEL�E��i�� �������")��LĔL�T��QTC���(��ADTO?����9��!���Z,ou7��Vf����\%߆�U22�o.��8���x�]�竵w�A�h+qp�5߃� {�p\��1�]��^�LsO��y�HUF�fP��FdSˊ�zu�7G�s(8w�$oc�����ٞ����bM���3��N��pF��!;����>�ٜ������|�8�n����u��Db��9��{mE��Yk�V����N׶�%cKT#�I�@;O���΄�d''j}W�ldLWk�=�c���Y(v�g:V#[�l5|�k�h�n7�����J�]�~.���#a
 C�Rz}�'kӻE��;��]��̦��f2mk�ul,�'�a�|\)Cz|W����ҵv�q�f��;N�e��w:[����k�l\�IX�����k�z�u����V���w.�b۰��O��
���#���+��'�c��u�*��d������>�Y�Z��꾅ܷ�kÓJ���؇j(6�ح^8��FF[[7�E�	gԆ��5 x��.jn@/����y7�LV��E��z�^����Wեh�.+Bn��E�k�%d����F(4nR}Ԟ�;#�
��ݜPͷJ����Ǩv�YR)Dw�����AZ�H���{����E���g��dX)��[���t��(%��o��ٌ�"�*�5�S�׌B�;=(�ArmGc����ڳF�dZ!���.�X�NV�\�i65�íUg�xb�N�T=Q�{�/�o^/7���x����9Vu�t��<�h7�@kî8J���N Q3~{O��r�6�.�g=���U}��W�+{.Y&�ܲ���t\&�T�a��7���n�s����Odfs����7����+؏c��|����J$Or����%j�O8��$v>���q�־�:�oϗ���a�AVzܼP⎜،�6��vP*�Aީs��0�������C��.���L,I0oj����gYݡ���u}�H)�*wJD��͒;YSֻצWD}��>�-^�hM�v���۞O��+�F�����FW"̲���N�����[f�=\�a%M�:룬����]�Cybg�y<O%��w��֯'[=i���	*����T�]}���)��s&�Ƭ�3�`ɵtv�9=�݂�e-q]��,S
콻�Un�7똨o�r��着�Ѹ�M�X���l��;���a��amy4��*И��#N�W0�Z"y�.{[�O]E�b;$�N��E���)<�mn0��Š�6�ځD�e�/'Ŷ�dT0�}><��}��v'ǁo���5�O����s�Q&ߣ��=ͼ�V��
G{Lݑq�����[�ɥYBf���fS΃��k3�\<�i�9e#�P�c��)m��P���<��ഢ;+1�5٨nI���C�.�bT�H�z:��+\�E�#3Jt����p�e;uo2����I�l[�rb�(م���a����ft�T�ł�a޹���T���KS^M�h��F:����&e9ڗT���v4R�|�]��z����t;������9�j5��v\a�9?b���ֽ���j��VUMN��\�/\���cvlD\𑰦�� ���5c���8s-�r�uhi���$��e�w4��!ȭ��]��V�Z�����W�zA���{jE����{u�z1 q�8]�����g:w}�^���.>�(�uĒ z���2�f�
O����z1of����b��=1�]_Ww�j�k��6�v�{R*�ߕ������{}In�^�$�J{��.0K�\��o~~/iii�tY�k�Σ���N[��:{�,����	�H��O,S����9B�7�!�����5L��X���<�,���5�Z�an+ؚ�	��s�UڻGv��n+�ڀg T��*�{�UYJ������ĥw����5��kkɧ�rwoD���٣�5��c&; ��4�s޺,��<�a�uzd�������]�-����W;n�	{{<P1���S��r�kB�uMv'.aM����lgU�^uJ���o`!�K`=��ژ�}#!Mu7Croy5�4�R�)�b�'���.Y�#
G�#a�"&#r��B
y�Qܲ�����ӕ�����v;QA;�#�;��I���zA+o35	���o�W��p��+�nm�-/d�F\��&�N�*.+�.O��]�kN^������jV��&��)�������윶� �w)c�g�8���&r�5�b`�0��iRm%z� -ȍ�Z�	�ۢ�w��U}�ׯ����*}Dgt��87y�Ԍ����5�w�V;%+Q}&�꭪�z{�s��C�8�q�u��P��b��x�5EcS�v�*�8��U!���.�Op�b'���m_��$������]��9y}��W(�wѝ��JQVSւ�x��o+]���{1w�%��:�����j���g�D�^oS{�]؜�\��4=油�����������G��f���oWT�sb��������f��vƭ�*���<%)9z�X9�܇+>���*��5鳙�X�bo�Et�n0:[A>ݶ�`�frka$�V��W�aK];�]dl�T�9��s�<�|��rM�[��&��7�����D﹙!ֻ�q� �����s�B1���D(k �E��Q�����o_>r�p*���#r�P����2�f�S7uoe9MC�+1�@7�ԫ��ci��v�mѮ�k�t�5a�M&�ˍ�w2u�w<��Vm�;~��^�]-��2im�܏]vL�ڼ�E>a�S�)2�u�x�n7����Eb4�IP�2wh ��t���t+�A��>+�'�:";7�<+t��Ż�;���I�����|�6*Cz��*���d�k��f��<Uඹ���~����R�_=k���ml\�I
����+->Md��լZ�WU�cpV�?CN�Zz�7�~�mjy��ی�.��9���*Ò;>s1��ҝh�[���[@�w|W-���V ,Jp�7p`�q����s��a��F����w���z��������Fks�
��vƌ���z,%|�X�)Q=H�A�<���;�6>e�L��ޯtD����c6�|�ך�A�5�z��r������'�S��`�2�q�0u�9=�U������M���Uk�:�����{���^����
��1ݶ�:���=�o.i�����i���[A,�?e[���	�݊�_���I�N��]��3�[��
e�_��k��;��F�K�3�"�3u_`���}��(�A�����u��Aǐ��[��1�1R;��v�h�g7;m��^Y����;v�B�^v�|�<�\���nh������*e<=Z��s�i����x�#n�������඗Fͫ�w�*�WR'��_Uߚ�������Ǹ.����E��O8ќ7��C��bB�}��l]ݳ,¼�3!��m#k'�-j�9�ʬ�XP���f.�%t%8�1[}{Zr�)���@ga�7d�A�BK�[�!���S����z�h����]���:y@�mv���%��t4qB�r��yn�����':�ڮ�t�V&�j��\���T"��Rwķ׸]�b�ȉ~��@�>��,��@)<�mm�m�]��5[�aebͶܣ����!�;�Ts�˨O� [���G��nhy�����^{�=k~ɬ�0�w�����(�������A��;�g�^TNu����}��x!�E&�{��|�e��dy�����8s�x�1ap[�Or��m�|�}:Q���Ҏ_���F:5pt�:���-�����H��WP\���M�'��1�Rn�����4�:�,��AZ��;r,�t�w&���0���
�ŃV�y�z���KU��[�6d\�&c��r"�fm��[i-ܷ���Ʈ'�n2�ߜ���G���+Q�,L��x]��)�ƚ��v��s��]7�49'��аHN�O(��f&o6[�]Xa��|�$�0#*M�e�O&�/2s]������M�w
k2-�[�����>�}�S"��-�Fmg�ռ��sڽ�Vu���:!�v*E=�ԱwuZ�Jy�����5�ܪ�鶗�3���}���J\u밅Ю�����wZ�S][�os�����3h;F�q�@��Fb��ʉ��1G��I6�Lݱ�}�^�}D#^�������k��u������r��*��"ES��{��H�&���:�1�m�
������g�s�:��k}rz��q;#�\��L�+�c�@��Wqc<�-�$� ���\�ʾ�*
;�o���f����<�����I}[HC�c�[�����b�-��6�o&���˾�Y7�b��<z@[�'�^�BR�Z��ޢ){N]nű"{!�:{(�Y%}��Y�}Cp(�/Rƽ!��z���3�#��qz�ַ�뤄�8x�>�I�B�+<�)��X����Tڏ[U.i^V�LX��k;��Q1�뾬&���ݷ�G7�����-Q�(Pp�Þ��>��(���3�������	�,��a�\�˶�B���+��B;��R~8�vv9(��#��n����x�k��n2�꒿E���^���3L��Y��ww��_���yR��e���y���m�P�L�����x�w�w�u��/�Ot������R�������5�v��x�J �*��CP\��5N o�4=�j{rhn�K���}���>���G� ���2�v�	�+�=y��q�psX'�(������~��r����bq^ ����D��3�t��Y�6E�PV����y��и��ڻ�ֵV�%�+�M�����4��yZ��k���f,���V�����=z��i��>��a���4��/�k�>���*�ٺ�2����O�۲�:=H�'�+ŵ���j��Ѩ���^�5]��s�5ؗ>sii��Ϛ�������;h�yz��V��������0�g��j�Ɩ_�\�.��~Ȓ�Ƽ��&��`<�*��c�@*���RҞ���͕�3(��U�����a��N�QvlK��oc�8�@fW\���o}�|��Y��]]S�\�\��N�{5Z��R��t�Υʴ�v)���Ԟ
����]XgK�t�n0:��������QSUp�_�:��*����.�Aީsմ�W��@F79&�d#�{}/+]T�ar�ܕ=��|�W���
؍��}UzK�H^��GvX���Z��t�T s:���i���=���vU�%y�1��НJg(V=r�h�bR�K�����0��i���lT%��	�)���vo9�z6sHP3�.�����<y�����5�ڷє��C����L��ޙ���7��/Ɓ�wlTs��]i�e��o�<Ȧ��f3o��Â��;�7}Y>��(��/��C���p;����ѕ˺¼K���սb�8v�^�r�x(�F��=+�F��O��ne��tތ��lt�yft�������p�øV$)Q=H�c�9R�%��K�/(���v'�qp����Ģ�;����4��"��� �0�z�L��l�/u�0RN��o�)ۇ]�vڭ���KOy51e��9+��t"r<��J�����Ֆ���^��>{���˛�`$���6%/������6�OiQ�fW��Z]AW[�ҕ�kE�aE7�0�u�=�a�M���D3t������p1Yw�>�g'\wnoG�y�ʆ��S��65љ}�V�~��R�Y-s��qꦛ$]��c��2�+�4 i*+�s�r�Uݎ���ըP�����ƛ[/]9'f#M�f�.5�tgۘ��vg\ŝ�z���8ZTn���꘵�Jm.Ifr�?2'L��6�ֽ����~b��H�-��VR�����C���~R�0s���-�ݻV���U��{:�b/�>�]��k�wC��y�w���A��T1��Y�۝��V�q�5�n_X�4R�N� �K��Z�c�xĻjoNX�e���=�a�cR�o�Ѩ��η�����20�Z�˰s)v
�;hԉ�@eM�A��Є��{���[�G\�}h(.�ɤ{�:4���xvC�N)�F��k��U��WvT��;��ʗyȷ�k]8��7��vm�ާ���{QcޱC|��î=��;u�;�n�S���n���N�}ٝR��Y}��5�*���Q^͇I}$��2*�P˻��������p��r��;Pq��ao��Q����V%}��*ª[׋�Y��[��q�r�"��u��Qٽ��II���m�V�[�x����\e��;��&fU�V��S���l�N\Sr�H�x�7��S��u�㵌>�k�W�v,.[�QZ6\�ra�t�1{��fs|;:��)�=f�pU�]�7f�1�E]����g�f7v�4�YF�x��y@/�y�����ṟ�Fuj���]�m	�����*"^wo[�IA��w+���r�:�B3�G��.�[�a]Mrk����f�aYqi픩�9h�c/l ����nPѡT��J�\�Sr�k���J�]��@
J�6�os��RI>̮�����5}wC����w
�7u��EEM���W��:$ZX�H�A(R�u]5H�lԝcP��%�݅뒳y����w5u���x!�>�7�	q��2���M�;�t�`����b|!]f��0iˢ������B�c�7�,������h濰mj�gq�L�K0Ⱥ2�������)N�#Retz�W.�������Ju5�">Oh���V��/�Ǝeۚ�	t�q��i�}]:6qC�b����}�nF�]R[�-�J�H�Q�K��j+�ٔ�	E�aꑥ�y�bѽ���x��sl��%rΦ��͔��<��eu����;�l���WP�C�`^d�s�OY�9p�ή�)��j��pc�<�u(o�=�2o[V�"��3םyM��5]Hg�7������]Xoz�摠"�0^Pʝ.'9Ay$�����>˻���뺺��Jb��`�-D�SLU2QM11P1MU�ى)*���h�uEL�3U$�QT�M�1DQE:4��P�1L�TMQD�AMD1�ဠi��
J
�" ��
&&��
6�h�M�T�T�L���TA�TRiht�-TEF�E1UPU	AAPQMPD�[h
(���JJ��� �*i�����H�������������
���и��j(���EU&تJB������&�B&-$**h�(h���)��"�HbZ
J�* �(*���h(���*"�����.��$MMm���""���6uTDE3˿�9ϧ��_����a\4�:��vfxc���+t����*Z��b���:���R�2l�M��1vAא�<B�*�����*��6�PO���M��p�N�1>�>�[B��.VѾVޝ�xƚ��]����V.NO,aM&��k*��o�.�+�L2�Ĥ��O��GS���+&�J^�a�(�r�����W�'y��Ғ�>��mZ]�}6�e���'�)��~���p.�w)J۰D�Rjk�į|�v�$��KG�����O8�C����O��<�u�����]�9�d��qw�\�ޯK����j����JtsB͊aVՎq��y��[��Ofjx�;Ч�
��������6ts@�o�P����]1�l�^є�-���s��Wˬ���ф�tY�0��J&��7����R{kj���%JƖ�j�0��Oo�_)�U��rMU�44�����sqpX�S�w���]î��)i��_0�߱���nC�;�2�%ڳ�V�jT�xF+����\R���ϊ�V���nl��	�]J�dA2�N|��.�i���':U\Y�67|k�it�ƫ̭C�ҥ)�����<B�!T�'<ٵ��ӯ8#V�j�NM4�i�.ڕW�!��o�1�{Z@��M�<�R�6���Ιv���w�=M앰�{zA@�N(B]B��X���o���T�Aw�Ƈٚ�'FR�΢�G�kj��4�)�� ��ilP������I��zs��ٮ�+&�$�޴�hM�t��x�C��}��Qn<�vtz���#w�7��׌C�X��y.h7��;p��R��Gj9��W��[&y;���J籼�--�~�;e�w�B�)ц�:bU����]aU�ԝ!c�rV�\��W�ho<vTh,aM&Ƹ�5�����-��[ν�S�q��1#�l���+�ޗ�YK_`�[B��X	:ނ����aޱ��S:��L��~�c3��O u��Y��K��>[Sy�4�{����14�D�����%ci�k��^|��O�1T����
���x7mWHˊk��|��g��u�������ZB�d�h%xW��>��K�6.� _k������M���1R�~Ҥ�,#�cRa��lhZ�Y�x/J�TsZsk5X�ޒՇǡSq�4��Zj�xu��FR��*.��dA�k��S�tT)v�дQ����#�w�Gyɘa�k4^���3v�4V٢C�B��MJ��%=�[x�җT<�>�5�9ߕv�w���;\�CS1�h6�*91��؍w*z���W�2Ռ-�{opy�}~u�Gc��ۈf�w)&��Mv;�Z���@��+[��0�nRλBr�b�
:�]�S���f�tT)�؍��I�뢪R�9����њ["U5��&ֱ�5�1��o��.۸�]�u
�/>�� ����}޽)�q��oҒ4S�j��b��m�P�+�����CqQ9�;�mF����p��ܷ we4_PZ��Ҹw�S̎�e	t�}�u�U�gG�"��K8����SR�e��U������4;QA7���N��a|b�f�?{Os(3�Ǩydl�hJܝ�|�F�K�ד}vS��:�p��Q��o+���c�cOE��u}�{|�:��Q��<�z��z�-:�_=knJBj�On��v�wV�4f�Xo-�k�h�R���ƣ�%A�y�R�ON�N�SE��k�r��cV)V�g.�X����2��R�����tb�`����ٷRt��s�L[�w6���].�T�㮢�2��[��yDJ�,k�A65�o�1<���o�&R�~�-
�����!ԙ+�;ُܪ��N�k]�8�ʭxo\vP��w��(��_:(.7({՝Ց/s΍��{�O�z��9�}Gh=ʠ���δ��Δ���5V����?v��%�f���Ѩ�YZ�<{3�����>��(�'5Wna��v����6y���.�z*s��-ˣ���:��)����^@��W�~���9���{iD��Gw�	�z��jƖ������rZ�Ey�{$���ӟ��gC���O�A�<�9�#�u���>��{a�,W���ʭ��~�N-���}a�{`��Qߵݼ�u�ӫ�0�&�F_H�M���m�0ꊡ:��c��kɦ�Ï�l�s����;ڛ�^����T�'ѭ;��)i��<�z�`�3h_������OB�&g���Y�&���<�jˉ�oΎ:Ny[�ey)�����J�� ~�\�^�yS�R}���:������j�3t��e�|ro'WsvE[� �мŗ�Qί��ӸN�d�
���O���xc���Y��eMYˍN�.�]�̽AT�K�r��ݤ�"�|��@߼�:.�{��>����8��6��w1ϊԸ��br�֘S�\QI��?UNr��I�;oa�v�2q8��^wk�<Ƞ9����0��+����L�9��K��V�e"��AW�fX��Q���p��\q�mq��G\��s19`���l��d1��=��y�A>��8������F�1 r����7T9�*SQ.��u����Yy[�7�պ���th,aM�;A����m�ok}���@���v�V|��.܉P�z�7���=J^�a�yG���V��mV$�e�]���2bҡ���TJ�r�����W%��zF�����$o��k����u�y͗�z=|�En��b1�.��9�\��6�i�{{�N��k�	���^ʳ��q�^\�(�=���\��i`��e���^��h�jEN2��!��P_oS��7�����_X����H"�k�Rקa���Ӊ��=�ɩq���&Ws"�*�s��&���6W;�Qd���L/&���)*��t{��c�hm#�(=��9]9u�[�[%�����G!��r��I���'�:����M�1Q��7K�N�Wv?I�[\��z����-���<�U�.�͍�����0"�ƶ;��j����JT�+�����5���	��4�M(�Κ�+;�4�Ƶ=�t��ʤ���Eԥ��O/��[�;\���0[�u���z�2��b�/gq@�q@B]B��X���;֬8.�L��/}|{��+7���l?��}#����X3��מ8�nd��v�SJ�޵���"�n2��4�.�}n��:�Y���^�����hr]�\r��C}:p����>��[���%Y]������@�_��Mwd׻S��A���Iÿ2�;������۬�G%�l5\:�1���
���<�h^-���U40���{�*+�����	��B�Gu߬����nH��t����u:Ğ�����9l�Uatm�I0���r.{�.��K��e]�Czޞ=�	�c1|+2����k�$��5���K�d���MŘ�lܬ=Q��ՔXKk|k�c��Y�k�ѤŹļ��gy��9l�+��1�E��yf:[y-[�݃ymڴ&n2���Ue=l)�<�:�N�xn���}Q�������Cd�Y7��K3
Ivޱs�oz��s/l{��u��t�!�3(��30y,��e^R#NXW:�1�)�'�3u��'��k�	���Ρ�g+�fk@�V��E�$B��~^*_��(��]]�_�>����1�Y����ݱ�]�4ٗ��ʗ����V��+#U�F����H%~�-X�n(bM�y�}|�mc�ǉ���y�8�L>͑����������Pĩn�9ӽ9�V(%v�j��,z���I�W�Kb7
C�BGw����Ϲ��f�Ľc�]vDQx���[~���]�*/oB#��K��i�҈~c�']I:�;�6q���-�[X�k��[uI\\)��{:�q�����g��!�l�;1�|yn��{&�[�&���G�K�NJ]�+�g�;ޡE�Z�鋻�ù'C\�C:�5 �������x 3���i9���;��=�t��b�e�뾶�D�|�4�њ������V��#YW��+���+m��C�t�f+��񐻀Z�����;ש�G[q��6���<�1���Y�;�P��^H���R����U�\v�4�o��;QYWܕN{[�$or�Z��ʲ��(�G���C �s~��5��t�F�\���b�<�T�w��vU�_��c�&:xN�ɀyP˒�$��մ�#zC���IH�x�!�r��F��Klc�S���r���:Gn�qb[�tVY�V����\_�d�番�ZN�ְ� v��Uk�u�:}�<(���O�#��X�AC�v�~��Z]�ֵ�k�;A�U+�b�*5��O&MX�ƙ����;�3rm�D����'W��u9�/����\la�����D���'�� �v�ͯN�aŵy޸Db�讗����Fc�2��o���3�z��O�!������ţ�}aͬ��m Ս,.}��=15��֙��f�>]��囵��.�R�֠\�2b�PT��\;{��	D�˭k�Sκ;K��Y�:��omui��|��N�+r`9�����R����r��@�`�ұ�SNA��o]��ʵ�g%�xuK��Kk���>���t�=�/e�7m������?jֵ�z���j�{;Э��<�Ω+E��n��7�X���Cw����jU����l5�O�Γ�Uڻ
�؍��K��է�|�`�[:��c𓝳%���4�{~��[I��⭻���n�꾒�pNs"��j���@��u)i��X�v�y��2���.��[xLg��q�=Vme{���s�W]�+�b|h���ٍ��o�T����v��Q���v��#�7��� ~=�(s�0t�-&�cyn}�珇�-�*\�<�m��]�@#���lB}%mۊ���&:QĘ���8���M�;�n��
Tt�� �JK�<�\�=Ð�[j���~�w�|�Q�9/^o{��\i?h��nj�)��Nss���`z}_[6�';���yc
i6�YSP�6q�-{��w���.]��2�T�f�n���/�	^˧��ض��j��F���+V�{;���d�D��=�nsܢ��c-��v1�1;���Jr�Ú�(w�Mc�Oy��yh��וpާ��ӠX���7->quDo�״.�_R6%w;����N����2/���-�}iM��[��o�y���H�akz+�&5�*c��]��M���d����w�H:��3������VFg&��s���f�C�s����B��'�g�:�{{���{\fP*�˷�8�O\*�1="j����}���FXaok��y��Z��k�����h���]�t�$Z.#7��V����bQ��{�7�=Sٛ��Vv�W��͖�}[�>g(w�������a.�=p�h�v_�m��\��U�������ɕ�kx7�����W�Q�@�1ݞڧ*�%Ka��1��񅳍�̞,q7��]�����d�b���p���]����KM�<B��ˉ�"Žzt���.�Ac����黋�+ٳ���B�v�}{]�Dh�e2(���Oes�ۢ�Mߡ[����^ˤh#
@�oI�؜���su�u,������fUՐ�-�c_>n����ah&��Dƒ���S���n��N�SPL�ޱ�H��A��v+u��%>(�/H��-�� �K��#�:V7�v���0`Xw�j�Iٍ�6�ۺ��iX������|�ԙ Ȁ�S��LV�̧��ll�d���{��:��Z�LZ���<����n�6��,���$�!�J�m좓�z �n��:�c�r�8�`�d�xq�-�w]�w�c�u>:��7�^KRʴ���������n��J�~�,�����u���
P_���P���s+N�b	X�e
�w�y6_JaKJך�C�܌|��&.�Xطx*}�uZ�5ppl�Y�!�ː匹���N�t �f��4;�T�p!�{l�3j�u���d����Wm8�T�*U��=�y�/�*���J�d,���d)0{+,�Jv3�^����X�ͥ���l>�����V4r���AiB$�8�$�|p6z�ٳv�%W�T,�盲M�mp�K;l�V��88�Z�p��چ�?ZFfM̹@�z��%��	�w&�[-���r��n���\��͍U�ϭe ]k�lU�*���%���۬�=,L�ҷ�oP�}�v~�[�z	h�&��q����w
��:.���/�=��J��a�΍��P��n�^�+K~/���b��w�Ⱦ��R�7��/m@�%ud��9��Z���c�յu��X�vyҮ�.��:z�|������E���)�n��bs�O����G��⺻-�D�j�Z��aFib�EWQ�)��\��z�Yl(�y])���oK۲��f��:��hd�U�m�	�՛o#���wN$n�����}���B�<�)&�{:��ʎ4���v�0��V�]���-����hǡ���a��v���G��+�N��pJ͗���f�E��h��m��Nȱl��֬���+t<�ծ��B�A��1��Q�@V�l;R���x�D9Dq�7�OPV{�z��;�]6��IQ�sQ�Q쭷]f�V%�љ�SW˷��ส�]f��z����Ok���2������B���V��	��P��>=�,Xv(G��/�z9oӳ��Ь�q���pF6Fmo.;�B��vUl�	���unssM��cܪ�OAgu���N�o�`S�kr�-���m?��#,N7gm��{��hD��hS�Y�b�qu �V�)��}ݢ�ܪZ�S���R���_i$�W�I٩1�V3+W�/ @�߆��n����唒�Z��E˾)oo�"��P쏆J�,b`�1�X]��w�X#8���̘��si���h���MN���wS�;���kNai�e�4��:� ƹ��Z�U�hx&U��N���qP_gq�K�ӗ�V�w:7O��S���G�&iwE=N;�Q��l.�ӯ/�_?��}���*���:�

(ѯ�I�����*�f��h(f)�խuKF�A�Z��E��k�TS�N�l�*b�����i�b��(-d)���)i�t��TD�F�9�UE�ErM�0Q��m���*��1�r��9�@PL<ښ4�FM:gACE-M-4�MG0餈
Fjӭ!�)�i���i71�*�UT�b4QCU@�!TS6���A3��:�4�"&J(bJ9��@rMV�sh���!)�����*��*�9bZh������i
	!)(�!��EV�4SM���ER�AD�lh��Q�p���@?^���)OxV������9����B�a@������4K�v�p�w%0M��0k�7�xMa䝌��(���y����ri}����]}�6�v�u{��^�䇪%R<i���J
)�*N�}`������5,�s��sݸ�����C�C�
�;�}rq�lv���w|K��xn�����k���-��-���A\"���w���2f��)�����֋�n�}V9�_�|9�ryM�����O(�Y�lF�w��� s�^p�z���&5�!�Q���y�2��'9���J:���_��N��r�����N��]ʜm�W��q��f-m�5�]-VD�/u�i���,VfE5��O>
e����k��f�Ѻ�8̠_�`d�?=��,��Hý�`M�P�j2�P�����k�	���^u����\��\E1��,�x'���9���BUW�^��ud]/jc��9��۾�!�z	y��u{2&;o������V�	^�j���{SY=�D�خ�\t7���H�Ǝۣ�*)J���t�v �n#�a�s�hZB�,�Gsz���\7ς����f���0Zj٩{��e4�p���u5o�ޛ������}��H��#��tXE��gX���������(3
W��-�f��J�ut��羌�3z �]�Ϗ1�K�
�J����9y��ouí��P���c�o,cO�����X��#�lFϊ*���ίq���]�;��m���g�Ks{~���ڷ�o��v"�H��P���(��̅=��;�v�wRw-����k�Xζ���%b.�|�P����]��	fz� �>��+�oGoyf"�u�x���6-!�>�6+�\,�t����f�����0[:%k��b�94���C63�z�V�d	��[c�0����qz��B6 ����~�綫�[��q�]�����ER1�Y9�М61؅bT��r��+ΆEG���E;Y|`r;�ǻӮ�\���+	�+9Ķ�'�S���O���������ֽ��F�F�]un1�R�5�y�hUj�u�Xr� v�yT5�q�*q�F,��F戥;*8�jN���}��%�T���ܔj�4���@����	���	K�+�m3�����L����xA#�r�*��n=$}�P���ۣ�_C�&��R��2���1�&��]����UweX�l&���Wa�P������N�=.7]	Y�Զ6�S��V��K�ZƵ���rV@��Wۗ�l�k��Sb{�--���m�D���C�X�ڙy�W]��W����.�S���o��դ�����`�����F!7ˢ��\�of�cgT�N�r�YZ�0�W6�xsίgaگ�G�ؼ����>O���n��z��>E�*ڱ�18��{���=��bu{g<�;Ѵ t�����t�ǫM��&:��C9ұ�P������v��T�F�a�;&:me-�ob^5&�ۚ���^ڣ�=�k�7��5���4��V���ݹͼ�YO���R�
��g�F��n�����Q�e��5�5��ܼ٘&d����*a7��ڥ��wX��!{zJ�[�W+�b|h��HF�5��D�Wl�r1�v�gv��b��\��S�\P)lP���3֡��yd����U���<���s{�VԖܶ������}�zYT�;���ᔪ
v��ln�\jaS��
�q��as�-����B/����FV��\3b`��a\���w��ZL��ycO,ԀY�Q��'�D+���ܢ��P���1�ímC̆ݍ.ٯ#
zWW�`����FZ��z/i��9m�Z�6/�Qi��b�w
ą*'��(p���f�tʤ�,�����y�̺�}F�'��	]�a�u4�#5������cD�b�ve���lյ��X��aO&�;`�R�L�T��d�_g���"�z:}��fu/2�R��7���[�%/ao;�����&�T�S̙O`>��[��uKYfv�]�}�҇+)N��71�@�eܺ������e�[O��u^{�A]��q�@��C�^��ܒ(����v��;[+�˸�����)�n��Mw_^ϭ���8̠U�_\�[Yz��k�q�Vf�99Q:_������ä��sf�˷�q �M�7��p�Y��9z�$��A.�=p�W��m�x�ļb���m��a�C1*��θ������2,�r�gU+5��@��!e*b�0�i����Nl�]n�ç8�C��0S�S[s&�Z��'�iM�]���"j�w���e�.��Auq=HD�[l�X(Ӊu��t���C��]OL���s�����:����Z�<�OumS�b��z[����j�u�.=�#X�w�%w=힮��z{�
��X�����Bޯ��m��U=�y`ZeF� mGNb��@����5��-�}A:n��/og�Г��LI�#��i,١w=�a�̫j��>����c6ۋ.Q��f�)�M��f���w-�q��л��V!޵�����=�w�:��Ħ�^r鋺��X�������P[є\Ոo��Hv�p=)-���>�iV�j������<��=sһ&�Sԋ����' �"�tB�]��N�p�b~���]�O���� ~�%�n�����a�r�o�I���/�j�N9�܇{��;�t��8�@�m�K�4+�wRGK'j��6r|:\�F\�/����J}Sv���~����._�;������@:/*X����/��ϯ��`��c�d�K���%!]'W�['�Ty8��ҹ%��A���3R�YQ)l��S��쫠w2L��]�O���6��B�ަ���e
�*���R�Q��׭�CG���q�8�c���/��c��c��{�s*�XV��ՈM��(�a{¡1��}x۝�)�#:����N�X�����0�W��t�6y�ܾ�~U4�ǹ8�ek�����3L�o�Y�q�qfXx�y��#�(��J�̼�l�m�T���[\Nv���}�cʫ��9�;�g��ucw�k�����*����V�low�M��㎓�fa���(]zk� >�J��_.:�Z�+�Gpk�n|���J=*��~e��)�ʝ7e��faxѝ�W��ڠ��������b7P��l���3�ѝ:��S���.�;�o�z�.��ݹ�N�9�zalE|v��(�h8cMh�-�G.���.���:W���{�1�'��j��B�_��T�A'k���
_$��2��A^&�;��d,_�?fd�wS(��_���}�_�>�rZq��w�\-�u�\P@���/J��3��3���x�t�5 �X��I�DSu�o�n�`kΖ��F�u���\�Q=���N�f�k�
e
��
{$Ϧ�7�֍%�h{Lbs�Osh)�DG��a_�q�9F�.���ޙ,��	�b~�u�n(�/=j��ޑ��V�����~�-nR�y�L'c�����Nh{R�W2��1�t�{1F�͗��+Q��֧l �����F�:�3���:l�Yu��z�mi�g)��h���E���S�Pi�el�5մ��ޘ��X^V�zy���ū�$p=0u��NF�Ag\`.���p������u�_���ҙs=p����"em:2�VF��3��=�:�N�++�]����q~[J���p/�� c�U�*R�:Q:* ̦F�l�Vmރ�[%��,�r���a�Ӹq\�r�=��h�Cn��l�L��zj>>�5k���
y�z�{�eu���"��O��2���m-7��p�	;�1�)ѿ�J����l����t%y��7Wu��u������S�p\u��wٴ��˿=�T��宆�X��N��OZS�+�o7s��:�f���̸3	W�s+�S�f�`9�� ���ǾUN��D��YN�X3L��~��+��=S6�	qiܹ|��U�_���;o-xl�{4O��ƛv���x���x���#'�I;����Uù��tgNI�,�ș^5��U�˽�:4��Rg��7^\�;��t��c�M�)L�wP��[Q���!|}�E��'I��{=�S*��N�3+�d���yL\}��%��uaz k���ea�')��p��U{���e]�=R�B�?��aO�}�TM�V�,�ѱ0�쉛�*Ap]Z�����-Ym(�H}}�^�[���$=SԨT^�L�=p!�tr�s�r��@�i�R #�g8Ϛ3��+���F�p�������rq���Cy�9�S�t̰���7z�
ʗ��S�����߾*�Tx�\.6�uX�����Ѯ!��v�W~�q>#Tc{۞�&�9F�ơ�$�2��{��]5�0\�x$�^#�SG�s)o���b��8��{����OUp8o�����,�" oE��\M��+0#A�`k�X��3�u
�����Z^Ҕ����~���u�I�rG���p�J�� �E�)V�iv'���-�V���0&��k1�a}�Tm��#�.}���^Vpۼ�[��J�D�r>�D)2ͬ���Q���:����S��824�=xTe����'/�g�\���W��4��*v[�׊3����R$(^��''�и�=��ea؍�R�}w&/�I٢�p1�U������ƺ泞���}�$�D��ݸ�+�*%�^}���n�z��!��H厂��簆֚^�7Y��k��%hO�X�s �F�'����'0�\E:�=Ei{��Ƌ��~���3�*�h22��ۡ�z��Ĥq��N�bVݴ.}���T�����;�ϋ^�p�������x `��Q�75��:��Fi�Y��
�4:wj-7�B1C��L�k:]Ij�w��fn�Q'�Ո�At�1g��|a�Ҕ�lGu���g�M�SMo[X���p,������JN��+�n�a��¨��Y9�-e0L�y��y�U��u�̭�Yݹ�轗~.5^�uT��G:c��u0s��\/O��K��2�j�
�FK��=a\��i�"N�8\�ܺ��*��Y8�u�ɫ��u{Mx�L��O��R�f����z7իNV�V1��2�z��Ҡ�|rXp1[�W2��;���_\n�;�c���P3�yxv���:�k�s���y��:Xڙ|v��Wi��/�N�(n�<��us75�j��?����}�R��gI;Pf5g��*g�����iz�(����c���G�b�Y��	#��t�n�z}�yJFIf��Ux�b$��;��VGz�%�L�1=��dd%[,�]8��K��R��c���>�2�;���� 鯤�&T�L�H���7��ӥ�y�6�3��#�o�*�[���.|�i�NF�7deӫFQ ��i�k�j�<�����`ml���{K��\;�)�F������&�w.)ݳ#��S�E�C��R(�ڒ=��TD�K�����8��oY�S/�}e�ͲRѣ4Ȝkh[���αoa/gਜ��:|tM���f�w�w�;�<�ǘ��G��ۤh���C�<ˠ������
��Ƥ���[|��y�<VF�3�fw^����y>SJ�'2���KK1����^w^���v�h&)v�X:���yR���ő�ʿԫ�Hʓ��ߢ{�/��3dօԃ�ԮC�]�u�LlL%(��C���w���fX��W|�܃](������s���}G�ʿe��P��ݒ�0w?.��W��{jZ5��7 ��;`i~���F���Y;_��l�W�kaP&,�����:{����A��R��U�-�I��Z�EC˦+|����~���x����j�q#4��Vx�[��/^�u��^�='O�e�q�}p�
����ܜW2��A����6ϑ���L�����i�����#��ry�Ύ�8EO�������:W?0q�k=��YU�~>���t��<c�B�T�h�9�f�K����ҠFJ{�#�U b�B�ɀ7�uW��y��u���Q�&x�~%+C�@�Ps��;ᶨ�L��FJ`l���<5X���/YT�S�ԃ�|��1��W����GI:H�z�B�2��3�3����
��sb��ol����+��t��1�eg��'��j��D*��^�T�A'j'=w���S�����o�(�L���7�NX{;�3(��BV��/"�f'�9S�c4-��ܳu���x6��/7�n�s`m��(��Ú�X�!�}{�EK�2��-ly�H\�Z�h�W�8���\�6�f���A���n�a��VCMR��w��_W_��	/��̄'�j���r]J�6GV�۽4�7Ʌ����	���
�$h�,f9���:�ܽ��,-O�1]̌ed���c\�,M�.޺��u{Ar�Ơ���؉M����|��:�-�%b�����&@/��]f�����u���r���˳���3�y)��.��nc(MU�ku��gS���\��pF9�N�Z��H^P|]b�L�Nt��un���n�9|�M���5,��鷂k�^��j���>�-�'���T���D��e`��+;OZ��S8��Z-Y�D8}�&IͪOb�e�8f&�7
-\z1�ð��L(����,��]4,}z
1�<'f�N��.�o�:�k0o�Bu�<��(ɴD�����3��B,S���e9�t��¯IL#��9��T�lY�t�Z+���8��,}G8f��7�Xue*WɞY���1@�Y�먿�֠��HPS��3�[0̥�V���n��ޒ��Ēu�[2���x�%۸�,O����V��R�ϴ���T�n���oI�Ȟ���� u�F����6�I!q!xH��v���]9��`Hm/�O���q_E�Yi]�eZ�2GAĢ�N�����3�6c�-���w�oOZ�R�x����y��E�][I�yВ�8�q��1���y���ؽ�,�d!K��vv哕Ϛ��̘��m��j��V�(m�-�:߆�ލ�\K��A�XWkR�pb��Q�V$�(`� ���ݕf^�C����Kٚ#�g>��^2M����d�()�� ٝ/)<��{�@QU�\��w�ɬ0�j���dG��;�D_X��=��r<�F#yG�s����yI
�,�_>��z1a)Rf�g]�R렅-H���;SY#�K�N��۸��F����C���թ��t��t�v7cG�+,*
�V���	od콅J�v���]����s��u.��ˮn���Nh�l;�\�=(QԂ'%O�)J� �}�U��lo,2�a
�p,��@l�]9s`�WzK�Mڙw�]\��}S6]^�g�z�*c�U�Y�(�5x:_4Y�ӌ[]jwIY�^3���˛���wo.V!Ìej�uғ{����	b����op�O�r�
V]nӁ���oX����lע��G�˦�fb�� ���d�:�X�ޖ���(�U�	t�I�{��rڋf����G�Ԭz�-��9P� ��i[K�\,��j����쮲*.k���7�]v'�
A�V.�V]��k#;�֡+�S�2MC��H��z{�p|��Cb�Հ��[�3\\�}�J}٨��W��� (| � U ¡ӣ�LMS��*
g4�V�''CTh�	DA5EQS��[a�*�������b"�ij�hyi����4\�����T�s��A4�EPMC� "5�*�.cM4sa��h(
����)�n`4�P���4�TKEC͚((NN����UAC���i�9iiKcMb��#jP���:J-�QAE:T���[:����"*y::m�6�$��J�t�M8�l`.XJ9	��$䆊V*h�NI�#N��Q�����(�Ӥ9:i����Bk�4)t��޼7Ů+b�w�<�$�ھ�ם��ݘ�},dT-s�j}BPȶ<K;�EX���<���Ks [��/,e�rr{��S�:d���w?�Ubu*x{\�V�d#�}p��^e�����Tq��ǲr�c����F���y���3�W-�k�9��z���ʻG:)�����������5�� )-�.	���GC��ᣥ�hx�m���oڏ�����1�|v�Β�7���q]j�P%�"�:LL�qEiy�a.�]�=�΢��Y转��T�^[)Hʽx}L��|6���۸�S.g����;$���(�9]�rڱ2�Óu�iH�p��I�������-L��^�R�������W;�#�&r�Gz'�:�0ӱN*_�n��{�.�Wrn!d�&���~���_�/�&�a�7u%gF(w���x��c�l�;����[�B����گ�	'U�;�)ѿ�J�;7yf�?t9�-��ͩ��]�{�a��|x�P=1�c+���gZ�'}��ܪ�ƥO��Z�k�Ud>n��+דЗœ�y����6b[�c�l�2���+���ƕ`9�m *������ÏI�~gv��W�@��n����ء�&�/&8�z�,��`�n�+�a�ˬ�����;GyB{�O�(������ƪ��.6�)��B4�1p0�2ڡ�ǔ{�IL!Зְ��D���(EM�m_QY���3r�9�"����ᓭ�u��F��Wٳ��uȬ�:��8>���1��wo�C���\W��٩L��N��w��C���Q��{�s���l��N��9�]>MW�<��t䝢���^5v����p=g����)�ɚ���{�mW�>>�f\c2y���p��]Q��g��>��b�I;<�{<�-�wqW�-4�2	C_�S;���J����5���2��9L��ڸ{��O���X�4*�FF�[�l��I��;����q�u<n+��KN��Ѯ!��t�d9��FuM�9���|��v��8�qk�c����i$�D@H=Ċ.R鮩�����'^^s�JΘ��x����������n<��:�K)z��!��뉰J�������B��b|fӑ�M�Ӊ+���S��'���qN�	D�9@���&%*�U{˹�#���yp̯,��j	��F�rv��>���/+���ͳ(�\ �KRÏ��1ی�Ͼ�4��̇��T�G�������p�[�i��Y�%|�� G����O��P� ?�4�ހ�#����Oq���܎a��+zw�;\�OR�ژx�����*9�gH�05r��U�mV�Z��4�n�D»v��� d��1 [��j�P�+݌Z\s/"�@��׹c��믳1��qv������qRw]>��� h~ܙ���^f�S��W�KM�:��!>��rN���p5��Ⲡn�P�Q~���)�� v���ez��V����{-S�^ݤ6�U�=�܎ݽ$���&��<�}�+��T���v�/`�k�H5���酶'0�K���+������1�{W1���q�|˪��|��f�U�[)����z�z�Q9�2=酿W��~A����gg�u��7����>y��z��{�����s�9���um�)g��Ł��0�ٞC3�i�½�z�[~��P��q^��$�O���W��� �(��W-MTn�;�7o�83�c��h���K�f�[�s��q3��&p9*N�J���L�:�b����C�L�W��Y�{G�'C.N�zI�6a�ܩ�vx��,z�҅��㴤"�L�k�]�E��!�=����L����zG/]��6�i��Y�ze����>3ԅ�L���bW����Nc5��$z�^�_�3��wh8>�=9Ķsю�z� ��D�W��(�:I�3
��
��G���΅W��|K����ø-mӟZ�z�߱\^��X�t�|���t�1X��#�&��Z�В����ڰ�>���v��ۢ���}�B�}|"Գ^y�()�1+Y4�9�Wmum.���9Zd7��㨗��˕���ϝ���ݛ�R��t"���[�[o���q>.�WD���CS��@-7��Qiݰ��U���I@^ԅ�ϻ�*��ؽ�{ѧ{V�H���VO�+���>���=�!9v�<ݑ��ٛf1J;:��ole���Fq2�t�>3�����7���z"S��z��G ��&�w)��S���]�z�cZ�����2d�U$.��D���B��9���[�G��c�-��J�����ù��~�y�tץ������Q�T����s���TJ�tn(�ɫ��jW!��Ů��?>b�_�)y�D���?�u"_��?q�T'w ��(��B�p_�*%mfQ�r��j�uG�x�%㾯j��p���m��mUѵ��up��4�@SC���\�],���|���নF��{�r8���WE��Z=�x�*7/��;�>Z�F�]1[��X�/�>����뗗>T��g=Cn�v�ǣ\@����He�u��t�3e3�]P�T���⹕����?ך}�E�1��9�g��۰�L�����2¨���I��k����^>�1�U��wZ�O@�rt`��.�2)d��<l�����r?J�YƷ���B��*���9Z�\#��s9Rܽ}PG"�$M�;�F��3*���3(��@���Mw���:q��kyNW5���nV9Ү�'���,`Li�����9������\��58�{�4���5=��w���~q��7œ�+�����7� ��2��b�Oi����f���c���hS�u����y\3�3�l�{���f�)�q��@%���%vתθ�{6z��Ƨdb)��s�j�І9^�ژ��<L/�*�����mh�7�7��n��s�%��w�]<>�rY�w	���c|���z�R:	;�t=��z����	��^ޡo q����Z�=޺�n��q�[��rZ}�9�T,����.g淬
G&6rv���V�%������Ҟ�)��p��[�=��㬏B��F��o�[ӹSJ?�������� �� 9-�,�}>�C��ᣥ�hkg�l�)g��}�`y-�����	��7N�ḧn�m(�qP�&'��[FB���j���dª\�+'��r�Xq�;c��~|)���;w_)�3����vH��[N��Ǹ/Ul=�ꮋ��5c�Z��q�9�\�F����&�p�<�M��R�mL��Q�#!C���xLy,��TW^�zX�
�����-&�'�7��0լ��4l�/�nU��H�-�A�վ5fV􆃀�ip�!U�*�:�<խl_a��V�k���>mK,͚P6������E����g�}-�ޭ�R�|�Vfr鈦�B�V-e�\��� }�¤�Qq���?T4��K�d�&���_�
�e���ɕ���ц#_�o��g�aD��nX��9�������{LW}�KM���p��N�yk�tm�����Pl�>U����X�Xq�*̮?���O�ᕁ_�/��V��ͤ�U�5*}��o��QӇ�Ul�������+g����C^�ٳ�4ǀl����^6+س�:iV���@�4xvk:G_3�W����{�N�D5O���uc��^��/*c-O��ِ���PveV�0ΩwO2=~ٶ�O��O1Ԁ��F�:�����5t�5\;���gI݋�O%YJsʋQ�'�=�mV���=��g�<^����f\���+��g���w�g����$�����fd���~�_�'��<2�::�e��ґ*w�N�/|5���2����3އj����w8"�϶�hN9���<o�� �<���u=\/n�ҟE�V&�;cG�ä3�\[��O��+��;|ƚs��D^f���Q�'�@\�H�ӷ�P]��{E
u��1��$��VP��`���iG��Ld�GOjƕje7׸yj��el�v�+���^��P���V	P˥�3F�|�Z6~��l�v��1����e7`����_g��p.S.w�p��@^�q�U��j�w�P��sz'f�hq�)���a���n����,�"�}a@�)V�3��q5��My-���׍_�U��������|s�N�i7���2��)����t�$_�J}��W=uPkG���S��F�y�.>x������ێN�>���[!�|�n��u�f��(L��c�#��b�wO�xPed��D�up��Zpg�l�V����[��|K*�2\)��It�;���;ֳ���6Hz��M���V:�*%γB����Zoyԇ'�rc�th�|�|�j.�M���������Y1p�]�&��v����_��^���F�!�����F����;7/2S �y�z�Sm�v���� ��,���[bsuӬ��V��~JEF��<�u�n�-=�~�x8޿[L�+�i��
�}'�b�ީ��NT����P�]K���@5(^����|�'4��<��u1Ъ��>�T�5<�`�}�5,�b��L�a�n�E7;������箔��/��^��$��~9*Gc뇒g�,�����v���4=��#�#n����@/Y��U^]]g�d�O���qhb����]��S�l�"��G����W7��=q���pk*�uʊ��8�TY��UʜW���Bq�.���D�O���ֹ#҂X�ᙝ��oDT\2��o;�t��g�t�
�u$d|��ī���uμ�����p������tp	RN�L�:�b���2��L�[S�0��b�Ww�{�{�lU�^�5d����@ˌx��e�A�3A�av�xM�p���%�z��ގ|<�N��:��)��]�(ݝA�Ͼ3ԅ��q���bU�d�Z>x��=�~���X#����D�s�������W�����QCI=�f �a=c�<#<�����7�����^��]TOՕ�R���G9N�{$y'v�����_) oK���9�K_)�A-��wqz;�ϔy����h��uX\}Ojķ}��\��Ӊ�þn��ӫFv�l�fzBg՚�M{��(�au )փp
g��eq�[�ý)�xR��?�����ʋ	���'�h?�r���=��	Z�R#��"/�w���(uDvm���H!t,��z�m���u��M��{�����ωaȱ:Arv	�x'|`��G(�ɫ��A��eZ5����k�w3}����oUH4���̰1��0
N�A��Q;@�Zn�A[9f���ͮG�������Q�k�̅ ���V����/���p�Y�5$���0�ǩgTJ�(Cx����qm��me����.Ns���V'sx���k{m��VI����ܼ[��^��g�+���e�i�`�R����w!��a]�B��u�>�3���jL;;}�ǣa�p�����-����c�\'l/�Mk��s�OP>N�e��M,Rv���jgzʍ�"�ev���/�oJ�n_��w|}] 輩b�S�X���3�������;u��V���~��o�Z������l7
�����u�Z���'�yu�JM��\VU�k}�]u���B�͟��99s,8ÁdEO��]_��Gm *����B���L�������g��~u�_�����{�w�~����d����u�6iP�2���݅ޗf��fr=���"��F����L�ј_��p���qe��fc�hɵ㿷x\����o�AY��:�R��nO�����T�@�싌R��ȇ�A���7ҽ|.eH۹�N�����3 �LpD�&�=��,�ˏ8�;���K7�%w�5�Ì�W�����;TƩ���Vu���X�ڜ6��z�O9�G*���NX�z�Q����ޥoN�XTc���y���y]���cR��������69�p��N�`GiOD_]&}�p���Ds�k��Z1�ER#^^��j��uU3P���j�3h�ں����ޭQ`km׼m{,G�3���
Xx���!���0���IrFFu��\G01�R�u��Gi��k��'é|Z#�ó��dK��5�A��C��mQ��egڔ���0p��]7��{Z��'bV�.���cTjw/��^�zJ5�@ޯ��AKd���}>�P����5�o��	-ǧ1xf�=W� V�F6�t���w�;wh�F�� .���11<�h�E��hΕ~�+����W�Ec��x��V��uĿ@s���M�n����e���26vH�L&�����G�4�tS�.(本ڎeo	�wm:/��p/�L����5�M���ca�VZ l>��Բ�H����a�9����3�o��Zo��К����&�|۠5� *��>s[V�'�eN��հ��%��*G�����]Oa�ykm�͕�]G(I��|��:>���N$C����w��ݫ۷�&���:>�6tqd���Ո��vO�v,+u��6�w�~O�{8t,�^��9��Z:���p�:�d>����X���S�xQ9��<�a\W��J��aeGK3��������qg_�wm��T��G*|�g���q����^_�G�:Y9�f�A}P�v{��\�Q�'v��N�pjW������E�S�nN|�WO�Uý�<��9'n��*"3=�Tȩ��u[˛�Y3d�d:��zK�#���Z
4RҘ�@c�4"��{}�;nb�!�Yj��5�w�X�7t]Ez(�]8T�uvͦ��P�]�k���(�*���;��5���w�	�uݣ�>�	_*������8�eF�J��놖���6u�3�D�6��E<��#��pv����W���eӷ	��Яuz�Ҁ	�vn�9m0>�Et���8\�7xwo[<�4q�׳�G�NL��s�bbWQU��n�t���c	��J2����ջ�'����Y ����7M���F���CSO����Kk ��(�j�w��i�u}��oU�c� #lĸ; R1��hu��:v�VrS�8ȇ���)�XL�
;���b�kg����>4�đH�gJ��Gtq�]<凶lG���b-726��uw�o��{ݎN�jN«�������A.5�幢ڢt�����^ ])�5�)^����P��.�&�	�n�][Ѡ�y�(�g��X�،�޲���ZCf�Y�/�xW �[C�� �y^{&3��Kk+B�mO�D����Z�n���O�`Fm[Ѯ���i.�`�fs�NƠo~�K�Wv�����
��4��)��3z�<�j�7{���������`�܎��ȷAX�=&�D��M�1�wJŎ�B\z��pZ��4��hiQ�����4��
jسrn�
d���|`����Se�b8)�U32�t����V�5[����b���B�"��/�r�ՙAJ��0��⨮ty.��冓�2�im�m���>����n�v��3k:��^SʋW1�R���3<O@װ.� 2q
}�s���l�+Z׹FW�̃��zUѭ*v2��]�����G��чhRж�v����s�ڍ�
�҃o3������a�)�c�r �n��T�I�;��Nw�;������v.��e���#� �Tĺ��?`��:\vg1du3n����۳�R��*�������nh�9or-���J�J�*T�٦v��R��9�mMOL�		{G��d\��y�X��I;�t�[D�i$u7��?v�H���ԇhf�&�wr%�j�Tڇ�&�:���&P��r�y��%��jO�`۴��t�NP���Y����3Vu�\�h��vc�؛�y2��S�;�5�Vv�Z `�^�tva�E�ev���`����z�Ph�u���Q��u_c�a�׹��CՇʵ:ְ��uL��̲��/~\ٔwI��b��ۮCw�9w����]k����vR�t�l؊n���+���.+1	��v�q�9R��$x��V��sf�#���9g��ZHL�lꭋ��v������WK����U�n�\+-�`�};������Oz�@�_^�_f�� ���3L�����8rY܁;�;*�c�Q���4`���Z�F��h�� ^+�!խQ� �`C�a���uu�V-]:܎���A=$��	���5��h���cCE44S���AA�T:5��h(��M.��8@r)�h4��4�� SA���N���E!HQ��I�8�&��&��m`ւ�:^J�ѠӘ)t)
Z�A������l�)T6
��6��h�ZMPSV΅ց���N-*���u�jbZ���@q�O*�Cs:�h�r9#T���P4��SPh��IHF���b)9s��:3S�CEh4�`6ɣA��j��A�(54��@�Cl��К6�imh�P��[P�*��V�h��j&"��)Ӡ���m�Cl�*t5������>#�|
;c+;u>�2�{���]:`Yw��({b��*�����QN�7C�.ݳr�ؕ�\�m�"�;*�ʶ;���.�f��ɏ៶��݇h�	�f\p1�'�L�wQ��w��z��&_���@�s5f�\��ǒx?�����C��3��/�6��R�:��5��<�2��9L�L{��-͝yyr�����v����,��v�2����	=<2#n�ҟE�V&��cG��f}
-���������:ڨy�Uy�qd��#���(	��K���%γ���Ī�K����-u�r�e4{>�Cߝp8n�p�=%��3
�R�$�ّ��0����:٪�ݍQ��o�4�r7b}q7-��{�O��'Z4��tF_�S�BmL�5� �\h%5��p��q�naQ��q7���;���ơq��*6�;H����[!�|�n��]y��WU��cc_���:%�'�6T�Z�芕�F��-�Q�u9<��%�|\���$�����qT�1���Q�x���$W\��ٙ����GY������KN���0�R��ȸ;��lW��^k4\F9p5x*�El�2MGOTd��O�E	kobY�fK��탨E����j�����Ⱦ�:�z­W)<��d���:0V���ǯ���~�n;��6$yr�烢6M�KyYC��æYr�Q�43�ὓ�iѧ�^�#f�$.��Դ�SI@j_ea:Ƞo�l��}�X���d�ټw[]�v��<r�P!��p��F���uGN��p��U6��'m�`�z�RF�'���	�1��S��&�r��U�]���K�Ǻw��4_������T��k��[ʰ�g��X���G��}� �&gԇ�=���\U��w��
�c��-6j^���Tn_[
f^�ʘ槝L����>��V��eƾ�X�s�����,��w�z��b�@�j��e���Y�&�;��v�^ffW�o��v߲�x�Sţ~�B�t�9L��'GIr|2*��2���b�����!����͜���	��5���Fc�W���eN��,��(z��(\T��q��"��h4�sMe@��ӕr�|d��!�(t�y�l�������F��'j�f��RS=�o��םE��ۊ�v����;����~����8��{ ��N�zs��<���3ĕ@G7�A��n���gF�iq�(���]ĳ)mD�o��!��c���Ϩ��N��|J]�l�|�ժ�+Eo�� �˓`Gt�>�y���uX\}
�\U�w�}�s�{N'#�y�#�(��j�{�1ޝ�꺋���S��V@ђ	�vn�K�G�O;�e�vk�xY6�@��kI��v�{�%/��S��R�䚵����l*|p�:_@�;�u!s��{kz���Ev1,6����
�����M� :�]m]��9���e�	㓉U�;���<g�)�pӂ4�@W�J�	���+�[�ý)�F<_��5���\���S�شwF{l��^�9t�ёjd�]RB끴DĞ}4/�S��K
�[�F_�ܲ/K쭚{�yP�����vY�%C��=1+�2���f9��j׵�fS>�O�������'쐵��^�
Ԇo*����r.9*d�3,a�ȍ빃AK'�A�|l���gf����ǡ���4�ˢ��_��i���jj�|�����M�~����Os��u�f'��Cvs�{�K�~,��;��f˗�q��Zw*�N�K�Z�F�]1[��X�dǲb}ԧ���݇ޙ����_Kp2p;�S}t��>͔��_\?B���=�'̣T��^w�3w�nn^y�����׈�f�qg'.e��2p)>�� �W�s�v��z�P#`���7�O{î�Z���7V7}���1y~����a�^�/�^��A�@>qw�/;(շkc�qx��A���>wI�u<3~�;*t�Yd�\��_ڄ����)�%�7^�R�����3�b|(S����iڼ���% 3,�x(ݽ�wd��-��5�R�&<�N��	���yS�"��b�z�;����k�s�Á=o=��]Ҽ�����+H�ĕ�9��2z���&Ă�77�;�6��9�C�}�'������&C�7d^)M��� ��pc;�^�%{�����N�5%�l�7r*����[��~��k�;�h���Wp�5����ef:��T;T��W���fF��垎��ҼM>����;��e)c��Qߩ*�7��>��!���zq��u�
�����7{�C��5p�aX��P@�x�ZS���I�|��
���჋��sz�T��h�5���g�ϴ�NF��w/�wh����k���_��� s齈�(t�uF��s��U�C�7�=Jǃ����/�hn'[�ߛ�8o�v�&�FJ5�@]P'I���[FL�Ƈ�`]M{2�����k�f���d`���?�uĿ>����n�Q.g� 	`��v�b���ީ�u��^�ѐ��g�f�6mrp�[�p�����1�*�
��N��.hL�w�O��	�)���3/M�S�^�
ȩl���V��y���ɫ�+2h�Cn��J��6D罾No,����L��=5҆�s����-m�Y�������BN�d�W4*���8h���Ȩ�"�R��o�`'��;�ޙ.�����b`�׳qd�t&e���QEC�M��n��p"�"��
���QH�λ�ɍ^�ޕ9�cy���B��-�'�X���� r�au�g�y�����g
{�M��9��g�o�p'yW�旆|t2{~�]c+��xpu)�s~ͤ,�#c��S�6}���}N�ʟz<���+U�����p��Y;����"wHv++�7��Ȁ7.��ۧ�~��@
�����T��r��Vs�����^_�G����+$�!��'�l)r��C���q�s>.KD��e {�Y�뛓��WJjtoG<��9'n)?]_s�A��*�:'?�{ƾ3��Uq��P>ٗ_�2n9Je�������Rh�=����/���G7;;��8U����(]�v��aP�Ф����J��N�(�,�΃+Xv�K(����ўTv�H�WTn2��n�2���t�/�zxdm�:S�J�J��cA۵�]y���W���hhs�Lg��A�MT<�*��?@��i$�(��P\�ң<Xݘ��\e>�u�]��Y���O��א�s��}�)�ٮ��:�p�v����H����(�ja��\=�y��k�Y)���|o�O�&���|w>N�i7�茸�v��)���ML
Wq�'ۂL�?o�#b{�J���.b�ikĂ7ι5���4���#[Y����\��l�6��L<	���iQ]�_��Y�\5�#%�� ˾�Z��˱Wuٗ�ӆW��%�Prb9�l%�`WB��6{nr��Xyo��E�$�қ+Ht��j��{�`�4���l�{�j�&3�������D����ۼ"XМ��co�����;�z���ɒp)%t�A�"e:�WR���@�L��1�K�ɿ��Ĳ�:�e1�{tf��S�����q#����8ٱҧY�q����KM�o:��*Ac�U<�O̻�=T�=\��l����V˳$�N���o�/�%����?i��'A�DO�v�{9���]���;�Si�v���d,��0��cxm�H��������\n�5���tz���z��G��l{�Sҵ�f�ʰ�e<���H��J'7���^3{Y�����#}1νK���XNGl�or���*�zO�S���������ry6�}�S�y�����ǲ{���~!�+�Xl�d�>������S\�'>w:�U����p��Y����(��Z}�_�`��}����::���f�ӄ�;���R^�wU�{(IN���WGy�P/�u�wЯ�7S�#��:o�,�����t�$�9��"�|[�1.����b�������U����N�H)��η��/XO���X8���e��؏��v�o�ߝ,�Bm7���V�eo��2�W���;���\՘�X}jsScX�v�G��E��$hN�Pr�g�͝x���
�s�}��+rs�w���g�-��q�[\b�Hg���{�u�ﾂ�8��.ʔhi'p�&h�R����NJ��<7��j��wZ%W;��kw����������%z�/|=%4�ϟ���̭Gg70mnuQ��cd�>��K2��N�)[���!��}��Zn#Ϩ��N�S[M?��>�Y��ޯd��<���#����������ϙ�8��=ՠ�¯���7�dӻ���O�5i�XH<_�i��d1*�l�{��7��|�ߏ�('�����
���V���{_i9��7q9.���J5�$.�����}4.��9����ۥ �^a�8��(��E��l1��Yg�ϙ+�G�R�Q5q�'o�3��WҶ��	���Y��:5-��}\�W!��>���K%���8U!;��Q;_!i���锄Q��^�ꭅ�×԰�(���\==���Bj�M�t��n�_��z�r	y��}��M��S/I���pr|�Va�˗��Ϸ�i������;�>���tn!����eG<�g�x'"mU��"OՔ{�bHc�{^f�T����ꩨj�7v�dξ>^G�^���ֳVۏ���BܨCTvG�^�(���{�r�{M�1�*�8����}}��v%tW��֠�XiO!���G_),��â��a󭫻��8���|{��Z9�X��������]z�ˎ�ZN�Fl�or���T����BP`[�*��ktO��ý<������^i�|���rr�&X�_@Ńѫg/�������sd${�^�=���xノ���C��y9�����"��T�P�̂�?"��+&��ι��喞㌕Y�X�ޫ�`g1Ԁ��w���|��ϝ�g���|�W�ʝ7��Ou��^7��c#�qm�.���[+'�\k�ڤgz@k�MPaxcvE���A�І9^���i��ƭ�t+2��f�m�'��̪� �9�*�q�]��t��1�eg��}>�ڦ4�n��=���jw����a.�8�څ:	=@L�����T�s�`Yu,�7WT���'���̏<	W0"��6E���4�����.����Q�P@ި�(	����iO
�ˇn�U�d�W�+���q=6���9��#\�;���U#���}�@ޣ 9�R�"������/��d��VC��%ޚ�:��Қ�<_����:�&���2��N|��x�"x�����Lة��w��sf7*-�umv��y#h�,�1�'r�C�:��J*:��BWb�A�w�
�`{j�t2ܡ\��kNh�����{�#���{~���=/��ܸa�y�9�#��N;�s����+|T&��(І��rV��B�>X]�<r��N_�G��w���$�����=�n���|6����n�iL��1�bpmV����ױO�xS!ag�����7EM{.9�HL{R�tnu��L��W�7�el��M���sY�/&��3:��z|*^�
���Q��Zn7�\?B�Vdѵ�mq�Yǖ�����O�c���e�L�0�H��l>�*{�[lW�ii��_�����˫�p��fa\M<��'����N�w�oK�>7Y=C��V�ߍn~a���@u9�_�/Zm�M��^��v<����s�ޏ|���/F^)�]�<�������PLW��5�t�=���	Fۤ\��s۶����cʩ��T���47O}�k��_�G�:Y9���w3��3�׍��Hˌ�κ����U��y�LQ�JȾ�\ܜ��j��j�w���q֏��k3�y;���_�G=Q���*��ޜg�xnU�|�3��L�w<k��R�xr���ɢV�h��O���� #���΅$���R%J�4:��5���E�� ��1����:��=	I[�����Ӂ�ƙ�ï�-)T�*b��j��8v��T�@؎r��WZ�H5�dm'2Q�fsx�qp흈ʹ�B*mG��f�7����y݋=/4kz�gZ"�js�E°��v���kkG^�oWn�C�\�'��2K��]�^.#\�<�T<��n>G��7{$`�(_�=\.#n�ҝ�;�!��nkѓ�7����t���-j�4j�(yc���j�3�=%�GI=FPq ��ҹ	��Vt����~Z���ޗ먕��E�I�}�)���a���v��zK4�����(H����cܪϔc�����	�%���5�'��K}��+���'Z4��tF\S�BT/Ͱ����ò�� d�Ā�����z8�.+xLf�'iAs�-�/+[������s�E���Nי���%���O�;$L�\*�i���3�xTe�	u�"|z6hK��gs�I��ʵ�O���̕_)�H��;6fc���
�:��)�a��ܪ{�߄M�/m�1;��q��kWtb�i;4n�\)���eْx"w zam���+��e�~r�y#;n�˼��њ�gJ���1�N�E�tM���'n�P��u ��,���x�H�{}.���٫�/��j�1��m,7s�_do[/�~�9L�+�i�<�
�}�{V/��숋#f���o�dX	�n��rԇN�^�D��±�y�sB7|�� ����Ѽ��q�9���x���v�w5 �ųF��q�]�u�:D��P �c�WQ���/��0rV:��Q]o��������V�������; =���~�ri1�����PZ��ެ:��7�e���j���R��rI�[�	���gm&emݍTk��'�4�&¼�)��@�E���ԺN�̮�V�5� RoN���ӊ���j�r7���V���U��"@l[)VA�<�5t-��]+���V8�����X�:�d��P��8��4V�TH�`b�,�����K��w3�/%�7gx(a�\�7�x�@fr� X{M6D�%���V���WܪU�6*9Ȩ�S��z��w�b��n�Cs:��hf�#8<K�E�kl���k4�-5,��B\�:�ntsX���X|�vT�9N����Y����]K펺�RI���D"��VUo0��tLc�U��u�b�{',Y2�1���7#TɣNZ�K�-Vm�(��\%*�]F�)<]���d2=�D��n�P'�5,�r3��Ŋ�n���Z2��e����ā��.ڼ	�b�
V�
����f�K���l�'V�Xe^*�.��b���]@���0Ι�9�:s��w���\y)�9 \{�l��kuW{;E.��0lQ�QP���|]KĒ��K-k�5��1�{�����RVuO�&VX٧5���M]ˀ�TT�yH)Y5�ɤ`�2�\sC�J��_u�
�+��9ۨ9=Ņ�ݧ]�"a ��y㬶,e=�|�!uwy..��Y��8�Z�T��tiJ�v;w�tɮ)V�y]�(�ջ}��V�[㎯79�m�o�V�������C�Ԏ��,t����g�����H���c���3y1:��> 8.h���ʑu��K2�ԍJ�K�]�����p]�iR����,F�����k����}�X��T�3��}���tN@T� ���f,uҒ�R9Sep�oq��L�x���Ka��.i�P�@����{q�ʶ&[vS-���t���XŘ����$/x^�D��������&� �az��i��|��k���}9��6��v�05��=�������uU��8*=	���O���ս"{:��&���V�4�߮ z��ĸ��n@��Y76'�m��cM5�^�K�`_[�����2�s]�R�O��kܹ�
�0[��ľF�r��7!���Da�{Rf6>��I��m�����o��aVӮ�4��W])�n�cͼ���w.XB�z�5.\P��{�/�eT_
�Y�Jn-����X[�|�n�Y��\��M�R��!Q�7�����ǋGY�-r����Pl��ԏR����\C�Ev�<�C�p�ި��݂�p�#c�(j/��GZ�1���Ut�$(Z���)��
���u;�+��	�4�6;g#\��V_R�}��L�T}0�w_U�|o�0袝i]CLM�E:t��bZJ�:2��ֱP��:�̛f��:t�h��k�:M�m���HR��`)��M��Pk[�j�B��m�[m�Ei�N�
��ڳ��jZJ&�]�c��&$�F��M6�Z��mT�Ͷ6rD4�uMRd��K�l;�PE�(��Q�)����5h��S����m�ѡӫb�h�Am�V�`�N*�i֘��]mm��6�i(4���-hյ8�-�i��Ѫh�E��mӫf�cF��H���E+��Mj�j"�:��*�mTm��H�(31$����(�hJZZ�i��ɭ%kF�t&1�Oƅ ?PbP;M١�Y���=�ۄنm���z�5P��|n�km� �V,���rn�W<��N�m%V7u*�7[Q��F̜���U�kM�̨ۊ�.7�a8}�)����aL��w�T�59����}<Ǽ�N���(��~��F�-J=eU����O2x�*�c��S\�&W{kݪK�3+Լ�����[���ܯ8�a�L�rp䤼-�KG#�E��ܯ�K�p�c�G���*�e�������?�6���+�GUuFf�x�_��S��'�`��gJ2����> ��|]dU���>�0��4{��P�D'M��<tZ���Գb�z��񜘏�5uc�]��v,ǰ=Q��/��/�ۮ�+�
1��c�h� ��;A�*炋%�m�E�s�®�x3��L�X���2�+<��O�[��[����N�1�M���닐�}��V���vx��̀5�}X*�@�}4V��[���s>g��l�qS����S\v�F�1���2���fmL��t��d0��L�����6����Qù����L��Y|5|
��i��"˜�nw��ّjd�Q�$.��0I_)��S���c�ru�_�p20\ݡ����U�ݺ!`��~�tM��X��i��L�gܨI�Ʈ5�j��9�]�R/k�} ���S�h�E�y����7�KU�q�0Vv9�:T��Λ�Y���6N�WR>���#IZ,D��;@�s¡֖�B�>\n���t�ϮiMl�spv�V�CZ�dg>�P[�,� ��%{��=�*��T��1�ق�Q��HT��A��KFwFG��O����5+���}wB�*d�C2���
� �N�t�u	�n�VK�y�����\��2���a��U�.������\��c�7L.��ᾼf�k��7��'�-��{nAq:OT�l��uӬ�q�+K�Ҵ�n_�N�O-t��z���������Z����V�]��q��W*�~�6��1`��^Ut~�t�jL�n_\>׈h����eȓ���=c��Y��W"�]��ךn�3�|Y�˙c�a��*}G�������u���V�-��+Qg� �ܸAê��
g�����Q��:l"�ݳ!�xD�������*����ћu��m:E�� �2Pح.:�?0q�&{��n�Cy\.3��MOw!쿻�k����U[\iǰ�2�2����qZ��j���1����A���7ҽ|e���׃쭿r�;�՞r9��%��ў�r�r�J7�]���]<>��Vc�OgMxu7�ۂ��\��wݧ��"��Y��w;�DQvJ�SB+ՠʾ��B0HS[ܝ��8s�ye]=�ӗׄ�Gu���n�$��Nܦ�z���x'_Z}����6b���y̐tIe�Al̥6���]"�}���5�����nwf���H��ǺHqʾ�����j>��D�ps~�@H}P��R��۪�7��b�!�oI�z\�z�s²b�Q������{��9����|]y���(� od@Oç���<+�S3��h���+�ӏ����=��S���k�9�a�7P}���Qd���@ި2��Kd�2�q��)�8گꪽ���\����3�\bwÁmR�Wi��>n������M���x�_A���ayA�z7��ѫ��{YF���^p�If�rj���s��Mπߝ����7�V��c��ڒS5je��#��[N��QZr��͸�mrq	u�6���� ��3݀QQ��_c�ʌ��jG����L齙�	h���[X*�3�o�V���ɫ�3իS.��__x]��w>��[�&���5{આ^�����(f�s��*{���w�f��Yّ'��s7�.3׸��v����Za����<�v���q_���d����끕�\T�8/=���#'���u�O����	���a�n]�1����]s�{4'W�������̸3��Rd�8�����ySVt=\&X��I)�x�t$-��ɜ!PVK��_b1a۩ܒ�Mӥ1e�g���vk�w�nf.;����e蓱%����(#n�c=l�^&ʈ���f�*�r�k*Gv{�%:�=[iʖ���h��!�e��iCr������o�#k��C�߯[�T���ʟ9Y�:��u����R=��PN4:��xt׻۷Yල٪s]�������w�z��L�OzR W�+"��srr�j��&��m)���L[��Q=[�I�6_��=GI��/Ơ��u�:�7r�4|v\q2ye�קl�	�ə�';ު����w.6�m�n����gNI�w�I�x8'Bߪe���ڡ*o�틧>]�4�X�Uݴy�;���r��;W}U{���e�� �@O��(I���,���Z��#�����Y.ҫy�������rΈM\=
m�qd���OT@`�:)���kލ�]$�vWl��ĵJ�PR����SG�5�÷�\���8�YYx�l`3����]�{քK�1p&ui6O3��q�\q>���o��+��;��F�q��bkj��J�y[�e��'�� .��@)*�nZ_�L.<��F�'iAs�-�[+Ұ����֢������ �U�eJ�T��gd��N�Uԭ83�e3-�Q�ꞃ1�J�,^��D�K�	\ �v����m�4e�@-�L#&%2�f\ڗ�q9�O0��hP��VdVG����v9CM�{�Kx1Һ�e6�+V��脧�J�z���l]\*l��۾u�l%���앆�����!��;};~���+ԲK�s̖|\���M���Guʝ��3�W�J�f��9�4��p����w����am����]ы䝚6ܸ��Q��vd��8�v�$>���T8ṇv;w�lO�v1���S��W�ep��z�������U<��'m�E
�u �K'|�"�S�w��o�h���a�R��}r��ȍ�cE�{o��)��c��?�U�[>Ojǖ�m�l����O[�j��ǳ��~CW.'�ٸ9�
}/���O�v�f�/��*�zO)c_M�~����L��ݹʽ����΁���^��,X���0�!��;�[���d���P*;\5)B���>9+��{î��D�s���W��y���~��q��˙C�N��T�8.*�j�ÅqdUYˍx)GVR��+�P��
�L��c� ^�,jڞ6,�JV<e�T:P龛֌���\O���6�an��=��4��]�F(r��!:l����v�Q[R͋<I����S�^�q�J4��O4x�պ|W>�in��P��iz�(��ñĴs���	�O�W����f\���������р�׷��w���Vp�������{?�'�{��~T���!�$hgc;��%i"�R{W�n�r��.t�Ǥ6*�\��gDg1��k�O��興�%�A;I�T�ޭ;��ɓ#��ܮz�jQu�Αd�%ӗ8��0~���3OuC�2��v)-������CS� ��5g,`�_T������+r���7n�w��)��I@HJ�P=�m�X\|���\�}�u徯U{<�L�̿<��Zr0���=.iJdj:��2��h6
g���W*�Vuд3�׏t��ދ��KVُA~�h�9���'�N�
d�_uI�d�9����!�QO/۶o>���qz�ˈK��<[�,� ��%z��
�J�j#��;�9��V��y����X�v�:5��q/kh�QK&�;i��T�9���rT�~�e���q�T'w�s���#�v.�M�+��NC�y�!�/���E�U�{.��yly5W&�:��v���#����b��x�ʫ,��u ��Y=P��g'�K�������Zo���o�<�u`6�7V;�y8�۬oj���qT�X����͖>�:�d�W^�2㮖�����>��5��v�9�#3���X��<���V8�
���i��<���N���;�>F|n8���2��Á#���/M�������)�Ψ��!'4$�_}zO�t3�@��qź�}ګLl�u(V"�+O���Ֆ7:�٢g�m�:����#C���w1&�y�=�]��he�9a�/�s��k�[X��������8�s�kr��^��f�`�t��F�ڬ�	�z�_�6�u */z���
g���ʬn�U�"��T鰋'v���=��r,J���lc���v���צ�٭�xe *=��q�����;��{�u�t����vT��Qރy%�z���Jy��_�,S"�����W��P	{MPaF7Dy�jq�R�W1UO�_��ηy�=u�p��.�o�G?\�'�I��2�;g�o�X�fƷvt���rX�#�|(ͭ�h�G�[�����u�Q��e�x%�s�I�(	���L�1q�U<o���f>��%'N�\N��>��mi|�2��#�v���hsl�
+��2�����-)�~������]<f�<�j�z���µHU�)����r0>�wh���=%� oT��F!,p7����(�vI wdۄe���;���Kj���7!:�&���2��NB2Q=+��yd'����� O�T}��g��P��-���5h�k���m��1�rb-��ίv��ȧ�=2�j�ѳ�DĽ�F����f�s+xLy%�ٞ���?���~^�Ķ�2Y[W����#%*���-<w�uv�|,P���ݹY����-j,L��zV:Č��YPl�x)�b�a��%c7��q�at�BV�ڻ�q��n��խ�,����BKg-����y�b�M��ޣ}���rٕ��۪ʅ�Y2?� ��������KD���G���[X*�S9F�ei��yp�c��ϽC����ߴ�')����M�M��P�.�Nt�=5����σ���82��k�jĩf�o9����wD޼���~��V�X�U�T	�N�����ύ������e`L�ڭ�t���я�h5y\N�3k��˿�����>{4'/嗖l�r[�c�l����ü>ˬ�R�z^��q���u׫�ٮ�=�lx���UN�r��W9��zmp��
��VVU>U���olU��N�pf�A]P��U��e2{�2�ܕ��뛓��WMߏ�5�E�b�]����������>�X���'��^��+]t��͋�?x��pc�NTU$z��;������x���4Z��찙Y�X��|�^��=��$�<�΅u2�b�mP�<�l����V'w#v㧧n7��e��b�Ǻ�=��7)�t�t^�h�F��w �A|P�>��ǘ~�mdn(˧����iO��X���4z5ä3ю�;i������0��G�OrHT��j}�y�Ӭ���X�[��r��3-��y��oV��}��笫�g����J�g]c��m�c�u�[��9�#�r޲���o��2��s;���N��Y`���a���K91�8<�����-0���۽߭#�s�#3�7�=�<�i ii�]LK_+^�B�'x=�=��a���nᙿD��]��~�y�{��L��1��`�ZM�<�{���؟\M�K}�\�9Нh�|�<���#��v���r���.�N�T� -��@-*�`-.�8�.6��F�t�ɞS�X7��Wm��y��{K���n9��.]y����(t��F�6S�q+N��L���+H�*���dm<Ώe���-�Ĳ���%�*��D���g>31�:lzT�4��!"�/��T�{;ã5�8���n7�Hv�]ы��vh�7.�S4���4,��FH|:����s��]�iX���aľW�ճ�k2P�޻���;���U7	�v�E
�u ���1t��S���/I�=0���W՘n:��}��Ƌ�߭�}ʩ�Z�3I�XU�O�'+��w4o�{����K��^�H��?��9�v��VW��5/IӞ]/�j3�������/�~�9Q����j������U��.����=��z}'ײ�ö^?NñYU��J��p�#�Ck�ߪ���	o!�[��d�����s;ۣ�n։<�|��Á���w,�W.��K��
�,�6�w7Y��)�\+������GK��j]�"�=�z>\LzI����Vl��8\v3�vv�ucOSs&���%֒��:`ӡ]{7�;gh�	�f����3�Qn�Y�&�;��8�����rp�(_�Ύ��GU?z��ގ��VTV������Η�.!_�~��2��=�;V;�?�Yޙ�A���P��Jn8�}~8�ud��8T�#{}A���4��]�E�Hg���z)�����0��(��15>�.(��������O?��a�2������	^�K�!z�x=�8��{ ��N�z{g�G�Z��9��qF��c���(i%a�P$��We�U̥�{�������]�{��_��yָ�[��`mϨ��wl?�U) oMD��� �}4�[�������]6Z��= ��
g�����a��vF\S�FmL��@{"d?�A�S<=(��4E�T�����y՝Ξ���#/�m�.s	�����S�fE��J5RB�DOMQ�oz~���dd�	ֳ�A�V�i����#-.��o���.|�^�������e��ڃY.E��+�W_��i�׬��i�v���Xn�c��KpTF0�dG��  =�( *��@������@� ���PE�@�Ȁ"+�_�("��E�����"+��"+�_��"+�� ���PE�@�U DW�("��PE~�"��1AY&SY8`"lJ^_�rY��=�ݐ?���aJ��R=Ҁ��+m!��ZjB�$��$U*�%#65m�ā�0ge�I3m�٦b$�Ije*�6�LkL�+6ij�Kh�m^�G@
��w=��im��1���m�Jk�!,l��L�KVkVT6ik�Vʡfm���{�Ƥo 7�+1�+��Q��u�D s�cfP�����5ToW��M���Q� v𑧜�e5�i��� ��zPP S�{�z��0t ��Ƶ���wp(m�XM��˵��� �Q�m��5�70:�� �`���BI��;��֫���u�R�(�� v�V�F��c�l��a�l���.拰-��v�v��5�q�4�]�[�mCj��b�����[�:�NΝS��J�lP�ӹ�t��m�uv���Uu3+�ѶT�;f��)�-�X�=x����hS��J��u�)&��Ф���
�ntwm�JuˡTk���K;U.�چe�-�� �z���sV��q�A�ܻc[`�n�a&�UT�u����W`�ܻ7n�AGvU�,��B�o �z�c�u�TUn�t,4���26`-�N��)��l��ulb͕[m���g�=m��*��S���Q�Ѫ�֮�&��6[���m�2
��$�Vx�ȅ�P�N��cEle*���GN�p�m�����B�    �*C&&�22 4�&����R�M�0 L &  �{LM%IRz�� �4�M  T�A��*j4 h`��4�C@4���26� �4F#F�43D� �I �UJ       ]|�����զ�gٖ�j�4�X_<ej�y�H�H�?���q"I��RYPI$BuA���O��K�$�0�Yl�������_������JH�TTH�	$
�(k#]�ڈ�T%UU$I$��9��`dS����!$��I5�i|�r��iFOM-d��J�ENv��`�e�������W���W짪 JC0��
�Tr���5�ٖ7f#y2�@U�3�0a,#I:�H�;Ql�t����|����R�
����L4*�S�m�c季��uj��@��!����d�AN��h�kq��̘H:��3
⭔�V�Q���.�M	��;�������ZncYtH�����F��$�9x�uVy�����4��kcYY3h8~�d�vZ�7������=��`L�غ�Fn��cǷm��)�(�����n޺F�3KΓ��ޛ���U�G���3b���b�q�wr���Kf�n�hҼ������P�U��+ZG1ԕ0�F�nA�c&5(��u8�ɍGwYb�Q��`a�3(n�ō4L�0,ݚ�2�ܫu��&�E���*�"�ą2*�����)�Y-�L�Pp��a;9g ��׮�R(��]��h=�R]'V�zt��V��֯m�$��Q�R�N\8�P�_)g/M�������K `ZB ��*�
�L��0��%3*My;�(��&G[p�z��Yګ�]��MF���"�밭bh��e+A1��˯�Yx�#b��)nm�%���Q�h,P&�&��U[���Uo�"av�YT+Y$��20�G�����/�i���A��lG�J)�/6�:6�X��o1)��ˁ\���;�c��9�֪U��AM�+F�\l��I�E�ջZ��'\�����h�v��bU�WO^��a��%���v��.�����Q���^9i��R�bJ�iVT��n�����պ�ʙ��F�l��V-��˴���Ab��ܰn��Z�Э3
h���MnţP� �bͷ��ch���7�PU�i�Ԉ2�q�z���f��5����Q5D����9�����2`�N���Y�!�� á]�6o�0�I�G6]�ZJH��nMVڼ������t$��NQ��s���(�(��Xr:פ2�1�v�,9V�[�+�x.�+�\2��V��0� ��fM�.��w�JHʚU�HJU)�[@�t+T*6�?�۪�TU�v�-���z�%J�n�WiA� ޝ��^�zr�R�5v	���-Ռ5��66�����YB�ߝD-��^�H3t���V��JY��&�*�s�(ލ�Q�pl6	G^�[W�����ZqfYKkL͒�e���We*>Y�<�T�,�q��t(}���Aybի�Af����.i#WyH9Ae��mHɌ��f���o^�̢�Q�ѪڈV�3%Ƣ�"&^C5��Z�^jt���bv��4%���!d@u����,vD�n���u3!�����XG6�#���R���
�&�~G\'�r�e+�j��*��n�t�wMފ�5^�B���� ХI�+��S@�B� �A-��4�6MqT��
g*^��0�sE�F�5{�+�J��\�H�Ne(��m�)��� ��M��t�]�p٣���7�k~�mϞwr�˔��p�v��sQ���PֆA,�J�`)ɋ�qM�F��M�J����n�0K���)�W�n��eڙ�1s�WfPa]��ަ��,���A�Ց�mJE�j�ƫJ;c3eB^�qQV�t���S��fU+����Z�Z٬���ZZ��ΫAua��Y\���8(��-�O��U���Ԃ��t��ShSdZh偐�YGS0�3�6�i�%+�&5���J��C�SQًhZ�lc�&R�-�w{�wi%B6�=��mn����Q��`�V�z�Qr�U7�����+):���NܵFe,&�n����-��U^��Jee ��i�̱cԵ�5j�a3+K.�c����F��D*�v�X�����L]�V�S�%R�£ؼ����Hl�,�L;�P����c ,����M���-�:7�yoSnf�!Ǜ�bݷy2�b�Q����� �6ʶe�-y��4ph#T�6�`���fK�B�6�	��i�^�2��p�Iw{sw-�br�Ϭ+�
���7���2�k��c:� N��ټ����%�Җ+5�+��W&Y��o>��ػ��6�C��д̫����O���-���; �ygV��C�UG{�D����b�V��[�JR��BB��w
X�@L_i:Y+��h,k���6���M� .����Tm���i����)��#-�ʻ/sp��[/0љ�5lp��S*���Ǉ5�VJ�3sL�d��q/骃�2��gK@��XU�4�e���gLB�+9/c٪��Iͬq:����p��[�j��mݱ��t�\z÷� �����p2U�Y�n\�E��>�ԽWdBHA-�P����n+rRQ���4�,�Y�!R7M��1j�@{�EL����u�e��1:���r'��F�[l�b�\f,�P��֨����U��Aʸ�v��9�1��2Mb{�f�F������P#{Cu����V�3t�ʷP�����S���.�:�3� �
	�V�XzdyXm%G-%�B����M�M#��K-�V��Pj�I
��&e뎴f�����df^�r�1Q(m0AkYu��F�o]�
�m�h� �Q�5�����t�P٥%z"�Lf�4f�˻+��D9��,���9�u�3e5���A�
tQ�!��W�`��Am�(-�E;T�]+��L#X��l�VfmؼtU�1���M����b{v�ӌ��3�`+o4�n�8��ʫ�4m���b��&�R���Q�Ut�c1S�,E��f�6��XǲޫgY״��o�5��&�F�ɅF���֜���aS+\-V0k{U��nX���1՜� ��F�Q�n4�fF)w0�w�$�@#W��H��V�bVԇTƐ&#�q\�B�h���Ln���e:.�Q�n6V�[� ��,3���Z�#�l�UXlm�W��͉�*��B���b6���[1k���ҽ�4�Kn�$�v�����kaf�p���hf�m���v�XBͼӦ��5U���cu���ͼ�V�ll�u���A�Jh8���:5Ֆq��� �Lg�dGl���ۛ�	��h�3�@���!�v�ǲ���*���Sd���Q��Ӷ���f�����P�X3~�eҹA�9����n��a�:,��9�3F��À!�����52rK�V�� k�ɽQ�ӈѲ�9B`�V3��u��	�䯺��X�;@�Y[�4�I�J�Დc9c�{d��zV�u[a貂�	w�<]�f|��
�A���2�!%�����b�ں)�{ab�V�D�/.<���C5��hеa�A"U�[�U�X)��6�����j3eՠ~N���XNl
[g�V�A�#.w���H\�j�J�w6�jKmf���5���|Ay��:4�p���0P��b�֔�"[M������f��WI.���oo,��
7t�CPf���nI4n�ԨIw��ݖ� ��6��ӂ���xeK2Udy�kY�+��)�[��AFIYD�F(�&լ_^���On��5�6��w�h�fU��B_�a�=Kol�0������f��m7
d,�/ �{JJ�nS�Vǈ�պkYzʳV�T�j���jU��h��l<��YAD07i���sH�B�f:�V�I��Z�a��/��њ����6��t���-f���j��a�ܛx���;[&ֲh�{���Q�I.b�l�35
.���ݨP�SpB2:�W��U�Y�'V ����Ҝ9y�$�n��'�ڲ��șZ�Z6�dY�
�v6�4�؛��6N�h �,��cH�������晊�ö��T�۩q�p�~���TﵧO5��Uv_U�E%K��8�9^��U(SKZ8-fVZ����ɵ����j�x�zi�=yJ���T��k��)7:^�֭V�:f3Y@��c��� 8��,ά5������`��&��{�m �Һ��D:�����+T���x�4	�:7&V�r]���^���h�)>n]9�i9Cz���)�K�̇z�Js��e鐛��/6nAJΎ�	yZ��!<|v�+�r����n:ܙK�g������P�^i�p��({Ju�5L����y+����n��6��S��EXb[7]E1�̭"�o9ǂ�Bg7�YB�-���H��!g��uc��ī^a���r.�WLp�F-#V��h�/���=N�t��[W�n�}qfw�}s8�K�/'b�[U�
���#C-+ʻ�,q9��zt�	XǕ�?Ӝ��w�C�{Rg�'�ڙA��h]u�0���;y[��X���D�2"6�Iv^ފY�ͱb�ժ���
ۄN0��1���6j�g���#��U�8���ϰ��R�I�.���v�^��@+dt��Z��[�Z�
�f�Z�h��r�[6q1u)ݣ�U��J�.9n���W�&N�z��yثWs;ݱuIi�&]p6H���qn����agֶ��Qe
{F� �%����a�U���ݬ�tZ����g������a��ջxaB���x]l�w �����-�Џ9����9����&L��.M�/9���������1[v�Z8���Ѻ�X�:ӪN˖Ʈ�����Z0e���v�B�!�Xj�2U3wt�t�1������[�P��-1Ib��^\٦
�dZG�ʣm��sv!�y>�E�	���l�D�0��:f��A����kf��}��ҳ������6�라�ؼ"��Fm$���ɢ�O^���<̥څ^��҄NDR��M�A�U����
��R��h�W��0ш�9rl�g2��79ʲ���q�M�R���۬�|NZ��,�g]��Lj��7�2�#"�d	,���"��5ϳu�bo��Ǖ^��1��V�y>�,9م&��]�8U�E��Y�->�O"�7��w�p�@��K)�wx�RJ��5i�6ސyk�n�K���Wc9�yr:�am�mX���,K2�<�:&+C[e���,�*�*T�u��[�u	I�ՃE�ϬL��K���h��܈����N�r�����QfF��j��m�����d�3k�N������E��d-�o%����җ�ww�7 �\Jt�3Q�9+T23�'z�������h�&nGݱ��y���a8T�����c�����ixl��ݜ{��cky0U�M��F7Ei�R�3�F�/���z��8O��}������b��޳y�e�3a\xF��ɩκ!� ���ͱ�z��$�Η�CVѤ�P�$�J��cM�8ySW�5�6�n��W�.ԏ ��P)ŻI�.g#��%1Z��ɦ����Q��\ÄG��<V�m*�9�d��/�a�6���T������t��`���M=�e�9��YD�>VZSov4�9�� }Ű^9�fv(�|����4�u�fk;Wt"
�e�g�ݐR71��8q�c"�r�H�V�ې�j��١w��Çv7���}FU��nZͮ�I ȹy[�3Nh�ri�,���[Cv��T�վ��W��%4F,���k%��7)8�V�Uf�����xi�Hl���N��vf�_k���SU��kW�0#���4�'��v�R���S��Δ)��{�:)�{j�����ε�s�:��%�ʎ���9��w���J��_j�b,鏈�|Q�~':�0��NH�����n���ӰVTv7�ii��S:[3\��\vh�]�x��&$s���k�=�4I����KFYF����)�A�ϝE��3{�y�,+��*9,�H�M�;��;K�f���K��)�Wr��e�A���h�VDnmt)�BZ�z�TnP�J^kR-�9��d��]z����V��7^��
;�9mH�-�p�1E�*��2�t�V Q͌��9^U�,:
|vo\�:���r�mR�����+���%���'���\q�Y'y�`0�We�3�Y\�q2�NH���b%���)ɣn�kE_��R��&vl�	ܠ����}V����r���Y.���Fqbؓ��/1�)m�0^i������ĩ�T�+Bs5YyΘY'%��)Q���}�v,WW��;2�n�6�[T^To缓�x��+v�M�|͢�ۍgtn�S�_�5��W�u��g�;�3�HHFb�n���l�e��Ԛ8��I�Q�.�eY�4<��#aϫ7[�*p�w�+e�nA�s�� �b���AX�u��2��:��{Iۂ������fѭYM�]�{��oKȰ2���v���a��W��l������I3�kI�@��ɗ�^m�Ӌ�-���S3���б5�r2�K��&p��s�:�W�b�����l�n�̴�����o}�1PՈҶ.�Q����.V]e1]8��^� Z�`Q˻�<YK�)UF�-涋
ୢDcQ�0��k��*���Z���(F���r����O1������QP���{���Mnr;�hk��e�y��Β���a*Z�2��;]�w/,�r��jCw\X��]�R�K{H��%	�U��u�t����p�6A	��ZIN�q��Y��7t��jݰ��Z[���YrJX�|����s��]t+B�&�Ư4�u�zy�j���A��4λ��0����ss���K��cڜS��X#F�٭��q;G��hކmmq��'�@M��ʑ�pn6"�wQM�j.��"q�%PK:9�d�z�*ȓҝ��rU�O;�2��#At�&u��m��%�.�1Qby���\+T����j��HbE_w�"����t-˓��^���˦r��R�*v��)>�12Xin����.���v��ЭY1K�z�Rp���:�D���+�Z;Zu�����}���TR1�#X]"{��J��;%Maك�M��yu��15�������GLO�Ae˲�HΫOY��sAd���#}�����M.�.���S�]l:B�f�,3�zq�gt�l��0�6{Wb	���]B�;ʅ0�p��}�D5�s��}n$�hL�:1�{��6�j0/�F����[g��đ�Z��35��KF![���vXJJ��i����gI���2�5`��]�QY�XTs�bd�Wt8�����%e*�{9�=�7���-�I47��F��*���]z�!�컕٫��n��8r�J������V}+d�`\�8m�;8�&�%+Zl]�nY�B⁬�἖[o#��o�;{���::Q�a�d�(d|���LԻ�|�:�h�J+J� �]�s:�T���F��L�#�92���%*i9V3����Q��Eٖ���@����[�T�9$�I$�I$�I$�L�ގH�5뗎e�3�2�u����X�3Ym���D���:�fI}�p�锐�>��a�=]3E��u
� ӣ+�?��v�yI��f��iR��E�j�	��.��)T��IL-��L
��U��sv��Kȋ[��p�7|r=# ��As$�Įf�z:��:��Զ�<��cߤ����ѸvmF-s�)k�5��]i�ٗI-y�R|%m_,���'ǧ�<�f8T��k�9{���y�ȅ�7$��M*X~���2e��X75n0-u���Q��SY2��h��i�D�:|0�D��j>��Q�&�.�m��v34*�����<��/��{�8ڮ<:.�J��U�y] \o���&�𙏃e	�iܭ,9�*6p��PT�o`ҡb��׆��:f7�g\˸#/
���w�0�4�!=˿��������ߦ?V߿{>o�o��H��/�	 ߞ���؍��UU�x�$D�[�S[����_��d�A���ՠ��P�Jb��u)I�1\W3[�Ht�\�ޏ7{:���b�st��4��%G�KV-ے�KC��f-9+"���cB���$^�4����ݢ���ԺH�8Aq����V��G��ˤm������va�VF� r�:�v���Ʃ9zE]��:��7S�\�	����33@��I�2����Vy]��V����+�Ղ��'F��#L5K��׉�O	Π����&�nV^ެ+c*Q����@���f�'@z�\�ѝۀ,�⫴mKhm�X__*vf+y����� 5�z�Vv�f]�@��wGc�f�ԩa@��ѣ�^���F�#����
`�������ͮ�S�.'���xn#�w��)�B������?8���\��;NS9��)&��
>2���fڕ���gqq��{�v�	Yv>7׵�X�i��&��"[Ź(e�ץQWk/H�T9��}]*�94�^��:4�p�'�:U���<�ݚ�<Z:1����@����Uy0M���p]�M������b>�L{KD�Z��YIK��e;�h܍��s	w�QJr��N��M�ΜVT$��x���ތCz�t]��αmB�2��i�at
��9%�P�w��e�J�:�&I,�b �e�1�������s�ry*�`HYd'�}񱑉f�����*�&�s4��Y�@D������50!VG��R}�L������6w�V̓��)�s$��9�'y+nź$Eo,=��7)��S*�;&(7���*�mflEثe�AU7�Ke@�����&B`��,�s�wUT$n���v��KC^�C1@-�"I^m,�}����'���z
ux�ꭌ�㸋�W@��n��k%i]4�ۀ�e���6C�歅���t�p����W{�]3��,��
�����u��͊vvL�7x�|�������a[V�G��V"��s+q����kGvd��n����gܲ���S\��]*JL�j����6wX�e왹�Ʈ:.�5B�.n���QZn��aS�I�³5f�4�mY�-K&��D#%^J�[D���j+���$ Ӭ7=L�u���޳]�`u%e���^Q�e�&������GGF-7�J�ֺa�-Dh��vF�y��R�`��)���wm'.n��Y�/{��u��{@��cOD,y֊��Su=ke��s<��I���%����L�Û�h�ϵC.��C	�n��Dg�)[�Lf�]d�{&lP.��d�����wf^�},*��u'��;L��@��se��;(�y6.%o��ws�F7�so���y�SW7�{���f'�g�H[dj�o1�g�`���Sjq@�o���Э�h��CD�kl\�5�G�۽�������,>v��G��j�;s� `�̑�\�8��}!��Ƃ����,���u4�e]��
NW "+˗)���ȵmEs�����<�Mځ�fr��-WF�C��o�pX��&f�N�U��8��.�JŲᭊE����	Q�y}܉G�jf\XnvX(�wQ���Ԋ_+�d��PMy��nQ�Ë��&�8��ܮ����D#����s�U���Ӕ��YtH1���E[�o�ڬð�.�i�Zt_q
�gUn��B���2��]�
Q�Զ�7���oI��Ü��۳83�n	�x˕	��\a[��/��꬏e�i����'~��C$F�lm38pv� �m�X�+0�q9� ����9��wB���3e�SOI̥Ҥ.)ݟdp��q��i�;4�D�y�,a��4�(xr'�\��v;�c�Y�i�j�8z���-@��wCo�.)��V�R�����a��l2�����]뮔��xd�w�W��;|9����ۤR���4��kmD��U�zc&8��*���v^����֬��S�(�&����B��FGm�#����&�K���$Xx�k�.�DAY�-q9xHۏN��tuRt]��6���#t;:�<"(J��Pn�HJ���Y���d�N�Vy���E#ސJ�+���sSo�k:vuP�c�ШK���$�՝(�4^�9fr���8�Z��_�8$�W���z�Ҧ��4��	�{����]�&^���9�%;�{�7Ius^5�j+���/m8.
��"X�Y��0<Q`P��E����`7]UYUHI�W	$���S�=��,�I:z���H.�(uv��kh��X�?S����?ix�:ih�6�n�2JC>���+9ʌ`(�w�WcOE�N��KIy�g\R(�1���V�����]Ӯ�v'�-aD��a���k�A��SL�sz:�RD!.���&y�w��;�C�ݔorּǸcq�a\�횞�ȣ����4���4p�݊�E��F�-w�@���ưHފ�@��K�h�5�1�.�V��{����
c:ܜ��E�yBGT!�T��W�j�g]:r�Gs�GGH5����)��" �:bvhG�S�7�w����U�wfT��|�U���$�V"6�w]�%Sx��TX��hfc9U�Cde��bnhڗv�KjΗ2�Jw;��t�˞�ޕ�ҽ��u�#�+y�=�[�N�dp�x��n�͋���m!e���>WB���1�*XI�ARr����l'��ۛ�l��SL�lY�6���Q��52SC�}0<�I=���nGr�Tš���Y!�[���^u��9���x�{@I$������#��]GB�,3���7X�Zt�Q�p�Q#[�g0���t� �#"�BaJ�|�a��(��I4��[�1�&f�ސ՚O��
[M�����u��m�%��ǵ�0/:R����\�/S��*7Ep�q���tƻ��
%[�Pw�U
&�e��^K#�ƫF1�*�o��g����ou;M8�C��;d���ۢ��IZ��(n�4K�Q]z;���֌����R����(u���MKM��-N�XU�S����9��[���n]�QqKN�DU�#��j�.�U�"���:L�!RʔV�J5� K0�i��oB�lf�x��׊Uv�C���+m,�HC���b�j��]�ff[�N�1�a��v���v��{�ҐȚTyPݜM�]r]��FP�΃6Y�7���i�`T�h��G9i�UT�5^�QW:J���m���YE(3�5l*�������
�}Xj=�w�B������Y��'c�7�,/.Y�ծ�r�֤��o�����Vp�8�ꕪ�*�ku%m��og%Q�H"��3��D�����N}���T�n�
z,{+(m嫛���T(�$�3(L���)�۷v����d&��W:�"�ڔcJ�g[�\��9V��4��mt��Y`µ��VwYX����nJ���Aw@�$Cz�&��+�W��$J�,��5E]\ݮٸ-��5����m��E�L�vZ6kEbR�H��	Y�w�)y�.d�b�ձ��y{��Ջ�w��)����6�f�v*�/��cz���lj�"�fC����ς�
x��з:�Y�˱hʂ��o�D�S�ǽ��4�����	��f�V�cq3�ޣ{�2�h-�̫����J�v捃`�_1E����2!cM����ho��.��S�l���K�����ZyH-�\t*���Y�U�@gsJ���^0�LPv�U�˯����k��ұ؎���lV��]Ȗ��G}q⩒�7P��y�pg�ҵ\ŗ���![��#ʻV;K�p*�hqB��pL���Y��VQ��'zҘ��r�*}�t�wzԧ/���]�oQγ�� ��`��k\�,��*	ū��Xs��C�_<E~�ߴ$�XE��!�����׀��="<@�n>��U�E~#/zi���\�#��w���%���n�\ed�ݙI�%]�����-�%&�_Ƥ�֘�%d;�y�yId�^ˀ��F��=ɋ�s�C�mCN#̓vWWm�]�4V#Xw@�6��.^�z�Aʉ���%tk�v�PL�ϱ��Y���8)V���*����Û+��0��+5��Ca=;���Y��iܕŠ/fX����'oiM$t
��&"�qk�.�Wa �1V�8�0��;p�π��y�Bo�g���i���2��<̾��6��O<�Y�ww���P,��ǉ��6s��b�U�����L��\8ə�]It��Y�;$�5�G77{Zrn''C��*J�̗h�J첖�˶`��.M뽴�e��Y�h�I��d���  �j+*���ond+�SGM�G�L�Qh��(���!f��e���pjڥ��%B��V��Q�������hؖ��q�[W�Z-Ab�m��AB�j��\����Ij!YQn��b����6���;�r���(�!U��e2�Q`��ީ��M3&SpM\��,TJk&eYX�Y-�U �
UkEbF��Sb�G,����B�I�*f�{忦}��_m��=6��"۾-{���X�jfen��UЮLF�C�G}\�N���}_���pR�V�﮹L}������ɻ|������c��3l������)tM�E-���w8�!���"S�C)m:���h>jrM��J�=w��KG��<�!��o�]*G�YӚ���%��}��B��C�84�t؊j��Ǌ2��G{F��s�r9ۑF�2\���k8i#�hq�������'�/���֮�#`ֿ$��Bz��4�i�ON���T6$�����0�V\���/�Sed��9��-uo7U��m��������&m�f+��wƷ��JF�[�%;�7D�֦㔞e�]��9�s��З"�ޕ���&�U��rnJ�m�^�ȳ��5לŤ��T=
�W+�s��Mk�f�Y�=C�}c;����c��H�>�0�]�fes���,�u�u
�&�D��/m�rQ�U3>&��3�m��{��:c�YB{	��Ru�9Y��ܪ'�[�y�&���x�#9Tm�Y'��0��"�$f�V+f�:d�
p,W2��
���tVTf�>�fl��yn�>��p��Jz�\�=����s+��B��H��'�s��kF;9�w���EP�ʰ��������K���ţ�>�7v�����mR-T6�p޹,�&9��i9=SVM��}�E�:�(Ur�͸ҵ��_����+=y���U ����� �[)�
y��QYj��q6�$��v�,H�q���R#n�KE�Xloe��a��gV�6jE��ڹMi%��;����8�y����ZOgGL�.��_��e^��6mZ��@yv'�\�y�� �=)���H�׊�9����-w:7PB��F��;��&ۘ³l�3��r�{����+�=SO�ɫO�&�Zh��S��3�i���n��^gY�
�N�X7W{�f(�N�z��gH_]�)��D�m2���:&g\Uhm�TM��I�'��a�lT�Kw�f�o��(o���&׮7{E<��q���5]�b%���g"���-�����$X�pݽ����)^�1O]��+�r����xl�fI�wC''T�.]�CL^)dMꜸ��\حCS��c��C���o�B��Q�*��C��v��FG>}�IB@�to���c�7�
�7Uש5��t0�@s�dT�v�M-�ZΏ{��8�*I�&���ԓ]��,ܚ��۪�"��IJ+���ĳVT �0�����F�����`ܡ��u�x�Ւ*
�Y3�'�i��	ا;"!w��E�=ĩ��X�4D��B�l����ʕg�8K\.�B���~h�v�B@�Q.�崇kú&4X�3\t�U5�V�x�9n�9�4��1}�<ז,֞})�ͩ� �vڌ}0C'����˹���t9v��������4�ŌF��	�l�y�QJ��oL�"��Z!��M�o�W-��U�9�v��;��9���t�D��'�1��N�V��<\�/4���|ĎGa�����A�Q��qO��B�@��Q�p��Q
ڊ��@���X��e���Yv�N�q����V�
��}�J��Lt��#)ʽ{�9��NO�씤h�G6��7�1ڽ��~���7�7~¨�>Xq1���rO��~}5&���ӳU�/R\��Q'�6bO��2�<�B�ý$����W(7�Һ�����ۡ�4�V�B%�É��[VNvvtda��w+k���w-}$��=�v�tE��g�_���	'D��<42�-V����b��8pmٌ���ͮ~��\�W����ʦh��C��H��B.�&:q묯OH�_J'a:�Wq�0q.���a���͒x�Lx�e��m˱'��:U	}ݝ�tF'�-�)�-1��	R�Ǜ�lޘӀk�Iś˷�T�t	�Q�B.y�CtDu2�so�Rir�{�UN�����x�^��?09�����?}�`��s���:ۼ|f�D�g���Ȉz�91��
4�z�YKX;EẫZb�K�+�����%=l���t������.ӱ�$uk�_+���WQ%����Ժ1Pި�h�t��
��յ�G^�r<Ze.����ϩ���)��p�T�6�q��S�Ԕ��+5"��MÐz�u!YE1z�V��3^�����j�����o4R��Wg$�:�����&�p�R�X8�iFu�欚��L&f��0T���խ>:��&Y!݀�CN����za�:����%˺u'�I9�<}��bk^CX2J^��\����F:���I�MzگҲK�����.2��� ��Վ��W|�)��f�֞���q{���+V�Ǟ�>S�'"�e��}���p6.�r�.�Z���Ɇ�o0FlV�"6���D\n��jwoh[�����Mq��8v=Y�h�I��u퉘�Ol�;D�x����̗�a;������*u�CLX��D1'\��R���Mh���D��$?vy�jz�_*��l7y�*�ҪK}6:�#ȯ$�&�����W#��'��9��s�q���íU�}(�.�R�;�QNw��=�99Nʅe�R�Xq�/�={l���o����Mq��d쇹{[��Z�Z�]}x���R�s�:���כ�[K�Xf�M�������F��zѥ�ml��"�e���˛�U�Ҕ�����#�	ٮ	��D�Ȏ�z˶����F�Ui�
�bmnI�_w�͗�z�j8�����04��7��IeYñ�z`1�=h�<x��Wv�o%�c��ӷY�:����#�X�����#X�Ӎ��D�f1�Q�8�����n�N��X�$e���"7v28�j��VTō=�
�B��2�6�o\℈��I,�gI�fꉞ�F��6�AiU�^��E�%]Y˖mf^��/EP��-]͚hlF���Lm��JT�]����r*U��)AS\����d�B������0n��k�*P�R��{f�P9��9���N5������*��<zv��{ڱW�
��-XΨ�ks�f��z�}�5'{I<��sV�4(�Y�V�u�S��Z���VrL5yz:v�MiX��f�+s�g�kMg�om�D�c���o}��~4������3�~~vw�k��A�����.�<�����[��Ϗ��=��DB���}��y>	9&NۧpġL܋{�wP)\�ʼ��\Sx�ۓP���Y,�V�m�.k�7���9v���$n�*8k�as��,�Q\�M���T��yd���)n�<��:��;}6���le�{��D��),��R��c�����������{G@������j�E��2Q�s$�Ɇfw^�n��j�Y��h\���S3�)�0��D��s��:u�L��7�+3XB`���'_S�����Q�I>�T�4v��ˌ���8WEx^-��Id�,�kU�:	iN�}T���xW8B8/�!Wm&�yh[A��U��.�j��dSwa�j�_]nL1�Q�oy_u�������4䙿�����=����*���~8hq:���,�CM���"H��eu���9R̋��zt��R剙`��Y�B��
����_=�o���(�9�)�mm]�b�kI�����j]\������c�ա��hЙ{��9��42�a��ou(h�{b�h�5h�w��	_K�
��p�f��ԡ���7D�/�4vl�[޾a6D�ɝ�6凞2���t�� ��W�%ϫ[{g�L�*ō�/�뿑�ZM��j��Pv���.�i`�ۖu�g؁M`�]t�ծ�\.Y��r&�
ѭ�h�z�}��)���%�[=uv��ti����,�}$����
E՜�|��Rt�9I���RB���:l�xWs�7ZI���)��@4��|��f^g�ￎN�Ƒ{E��7,�Z*ZE�0���\�\CI���aQ���1���9UJ���,�u�e��kGb"�b"ZXi%f�*�"*��UAMe� �--��QLeV��
�+
"1dUQJ�Xuk�6�Q�HQU:B�XTcY%Ƣ��������CZ��ł�`�(

�Պ�%h�UU�X��4���kU�
�c,X
"����4� �]2�k��ʀ��,[QAAJʋs���}_��W����TӔj��T3Sg�m���C�%����ɐ�������f��a�,i���K�Z,t�[y�Ei��@���� C����xwR��c}��'����z�6���HU��f�G^>��#��xu�͵��Y&9J>���H-v/X�������kV�8���}�bs)���'4��[7�����(G
a,�A�"7��5��u��F�<�I�WA�>�����"G�+;j���/�7�O|���!��W�l��o���m��X4��M���K��;O�Y/e:xj�ڧ��^�u0s����}��G4v�λ5�=��Y��'�sE\U�~�.����l��\�r�\�N���u�2�d�0��T8�~L.k'_{
�{c�[�>]+������j܇���}joNW���s�~�o(�7��#566jv,�zn��ݵ�V����X���w^��j	ƹ�-���=��]6�U�V���V���B��]U�L�+	5���sR�����h���teA�ͣ2 �ڷ3�j��jI<��<�����b1��;tg8W��㇚�$?i�]��W��V��k �<V�NmN�;� f�)8$�j ��� ������`�^�����)%���볲��ፂ����Br�9&�I+	�Xp�� ��utٖT=�8�qH7y��l~�'r�V�e����}��ow�;
{�����!l.n�i?.I�T��f�hV13ٲ�������b~�ҥ�WH�(�Y6�V���4�� ���;����*�/��%V0KV1J��57��e���+�5�i�ޮ�³R5c�K6���S��RR��
i�������c�:����B��1ƒ�'V�Rf�^:���u#[��Z./P�k�z4�|k.���pNB٢]��(�����V�=Kjɼ֙9��n7� �AޚQ�A����ev�ʌ=��!�W�������:
*�\�/B,��e'!������P5���\{�|��Ә�i6Q��y�O��#���%z�'�{�as�"�#�@�#qƣ0�<��D&�i{/��:a޼U�k�O�T�� $�}�>�}�ϻ�����d�7zIX&r�m�2�x��h�2j�^�՞�N0��'��s�z{�5�q�y�|�]y缁�����8�<a��p�Ƞ�O;d�!֨c�	��d<�)�y���7�t������'>�205킇L��|�Y'�4{d���H�sva<d�;2����T4� yvW��k�|�>��c!��@P�)��������{H)6�OY;v�=�Ȳq���I���u�͚�޾�~󄇬1	�N�:M!:I4��O����q����^��>I6��OPw�u�3���\�����1���z�;f�Hz��S�i h��|�z��i!�(C�x��'����1��L����u�lڏ��Z�����
�����u�ʙV���'m�Y�=;Đ��<�3���ڞ7�f��w�qf��#�v�VS���)7�R󺯾�7�|n���|�R�l�!����C�M}d� z�G�0G�ǽ�^HQ���Z����ƙ4���>� �'�&04$��$�P�'���}d���6�m��Q�"d�����۹�����$9�:@��{N�>d�&�6�i��(OP���t�`,�8��@�$�$��ϵ��=u�κ��&�cNԁ�>�i'�<g�6�yݒi�G�O&Ol'��;e@3�	�S ǽ� (��l�5�1�} c`m	�!����0�6��0:{a>�� �&����Ol�!�����]}�<������a�7d�I�P��>Cl�d�(v�=a���I�M{@�����'��'l6�3����|������|�p��՚B�`��`u)I;I�kvHb m������N!�t��L���52��	�z�O�5������w��$�v����;Ci���(��x��T��7H���L;I�'=!R��z�+��s]��������a5�l��'�f�!�x°M}I>`al'�����Dǀs���x�	���oÚ��&1 퇉!�a=@��Y�����I4n�RK��@;d�l������4�z���?!{WK�w0�/�O)���i�1���Ḁ�C�3�i�ܑ�{�TW��_�+.yẜ�	���[�)V��&�ޕ*ԣ�������{���������A}d8u@��ɶI�*׶
d6�{@6�T�Ę{d�IP5���-���Ϲ�:d���P���4��5�	�!���%J�=���ͤ=Hu9`|�g���lkݎ����|�@ē�gvE'��!���O�Cl'�=���d:Haߔ�d�;O���
<G���JT���V�S ���{��'�'�&���@6�9d�'I�i;��c!�T�H|þY!w�zu�g���o�>`,������4��''9������N����;N'�7>�W��d ��	X.�������Ͼ䁴9��$�Ci����$���OY6�i�&���$�	�t{��G��ZoXR���Ĕ~��4���!�&P�$�ya�;��6�|���O�=�$4��$���i����;6^y�����g�I9��$�xÌ�R�gԁ�;���;a8�4��ɻ'��!�3���ν�5z�<��bV�v�V-;I=C�bHV�s�O|��Ր��4r�r�5=��=I5��I��yݎ�:��#~�i?	����{­�d�$8���O�Ԭ�$�6�8�|��4�x���O�M���w�ϻ��W��Z��U�(eKd����k�=
r ��8p�[~�}��0|�'��-*n�|ɔش���<�X�y+�2 �RR"���㩧��ToI'�� �3��N�Yd�l�
��"�m�ݲN�x���m ���>a��}��\��y��$9���I�N�`q�ۣv�i�_RB��P�<�hT;�x���a��w��X�����K�{��@� }��&N��!�Y<N0�q ��C��>d�l�d��0>���ϵu�u�7��&2t����!�'L�L�i��$;�&�r��<�=Cl���v�o�y��Ov>���<���i*��	�
��������I�:H/hM$!��'BV�킆�g��0:�/~^����p�}�a6Ƞz��Rqğ3���2�:I=C��!3�������C����C�u�}��~}ߞ�a6�,>d���6���H�|���(COI�C�Cq x}`i8����(v���P���8�����0����R2t�m��O7@<H�t�Xz�1�{���v�Bz���λ�>����>��C�$���`,��ĜI:��'̘��6ɞY=I6��4��XC��=��yO�ּ��}���=LH��6���t���4��ͰC��I� z�l��=Qp=�B�+"]�����I;�H�ɺ/:I��t;�O|��;�
޺�.PK-���W�Y�|VY��Q�'�,2���%����FR�}r���y,��E,��$;���~�~�0?�4�m�>d�S(z�m�P���d5݄�=B�ٴ!�)�'��?$�t�����͜�k�y��}	��YO�<`
sv�&k��]YX
f�'l6�NG����=���ב�~����?��^�����}�t}�`�MQ+U�[�Ƴ�x���l�9z����2�<�F*��ۆ�7$�=oK��)Tي<�U��Z|6�W]Ģ�R;5����φ�C8�:6�D#7Gsl���r[�sqP�F�Y����gO�
�~�@��V<^���@=����?=9�|c�Zֵ���ZՉ�YJ�.�0f�ڛ���O��W�ͱt��2��[��j˫��ȷ�؞��*��P�d��e�_�s�Ce��+->��a�Z�97rmeΕ2$g)eM��K�� <���I����]pR8����cr:pj��I�˼~�4-�d���d=���	ȵ����2^��H��.��Rی��VWC/�r\rg+*�u��s�8����{��^�Vj2��C�t��loǏB.3�jK�����lhТp��!)�s/x?Kr>Q7��Y��Y�F���[Ȗ�����o*Y۞�1�9A��|ߓqs�!�����q��wN���ݔy����=��=(���kOZ8�Ѝq��ef�[�q{�� �%=��u��p������v�^�⌘��~��.���2��{������m��rM���]79WY��feo���=ƻ{��.,<��p$�ڴa��b�N�63䥰r��F}�3{Ď���u�E�-�.�/���8'�&A���מ�=���m�j�-ʡ�[���K�s]N��Rݭb��V��O�܆8w�Z,#����R�ֽ9S%ڇ�x��h�Uyu>�uBޘ�5�賖�Kh"�Fi�����Jm���]�q�%]2�]A�=�ǽ�z�F=�;q���������c�z�����ۇ�QL�-`���~H�h��f�J�Ԭ}��買y��ه_�[z;*[چ�29Dʳ�p/��Of:��Ζk(Q��%#P�C��퀇ֲ#���l{6�oX7-�hT��3��U'Y�^^)0@.�+,����iXp�j������ڍm��Y:�Ł7�Q1�6����ب��y/�X�5vm��[p�����9��9"Z���^孊��÷M���R��袴rm`ؕ9���S�,�	 �
�3���
SB�j�8X���1k�ǂ�Wn	,܂L:Q]qY��]y��S@�4@{���;0P�Y
��:�v���?!�xgE��*|.�m��]�ml��7s�L�m.�c��5YyG�
����)նH���Xt�������*�s��w725)+���W�V��a2�]DM�rTv�����ۅ/�P�?;����\H���z}���-��\w�]>8<�+��g��ֲkq�9wuq��7��z	;�cwK\�ҨL��:3ba�H��nu�^;4�(D'=�û,��&-���㌒+��w7:����kY`����G6励��ro�@�О�$���-�r�r�H��t�9߇e�oM��Yv[��Y�aX�9�m���]-�%�jd-ع�7Oy2�L�(U��!���ώ�=Y�X�Y�iT95�W�kH���X�ob0-ӤX̷g-�YEM]���e��npJ�7��uul��0�h�����Z�V)�յ�X =s9�is�u�F���5���Ǒ[��T���H��O�Ss����ϸC�;K;��'Q���A��ٳ8�*ȗ0�{�|������,���d�aU�dU�R�|�`�cZ��(�@PX�T���Щ�@�(
1Y�����Ȧ����,����F�ʑH��2�U�ʂ���V�ibµ#��c$U�V,b��AH��R
cm
���T�����"Ȳ(�X,"ŋ QT!��r��
Ȳ��[(i�_}����w������ފ�7"��y`a_t'm�Z6O6(�L��_j�^�Ի�q_|n�?�{��ϋ�U\֎9�J_�.v�w�/U���ay�Vo�����j���ؔ�����B�)�-��	U��ۮ<n�9���%���2$h_rɭ��2�XX�%g0L��Fo��a.8v��l�����cy�$�z4]�J��æt�I�Y�nV�����-�n?5�]��ˢ��b�3���B./x���~��iu
��{(�V2ݵ�(��7��qn�jH忀�=�e������n�$g�m(z)1��p�!w���<]��bXc���(?µ�K姼_C�@�`޴��͹�$Nn1 U�c+��)�$���>���;xR)� �P "6���M��zd0o��w��ȤT�."�1�kF�kXX`5Q$�6z�|��*U��5׈=���SZu��f7�UN>�h�&zX�kYx�cL�{3�Sa����g15��).y8͈o{F�q�n�Ӵ5���o�w;����diFWV��_�ni$�`�����Iv^��+{M�V�H�y�bV����%.�V�	R���y�=��?z:69ak�����9����z���֮P�Os��S�Y���`7puC:Fo���)�Z���x��l�b�x��qZJ
�r�)v�z	K'	�W������D�����d�t���'qT�Fn�)3�;�ޗ�١��̃i�0�C�x%�i��j&�����7-)�s\�0���r&I<�|>>X�ϝm�����B&�Cq�2�6T2-ɔ�zc'�a��>��ٔoy<�~Uh穎-�%<���^�Z�,�0D�:�+�l�)tG�Y��U=<հ��Sn��]��1�m�[��3�����n�j�iH��tۍy���g'�d�O����AM�yy+ڣŻZŗ^�U��:��它"�K���G&e[Ύ�~�����'�>̗Ʀ���.�&��Q�w�,��:a��%~ � {�ksQN;s�����`�˪�,��iof��JۺDS׹���l�܀�&3�-��ރ�.tO9�t��<pg;2��4��#�#���5y��Z&���v��%��E�]���;!�]�NCYŔq��H�o����:y�i�v�=���bI6`g�f�ѭ���'��pѴ�m�cEY�Zu����;�"�z�ßY��8��b26kY}�Ѱ�zI�[�W�M�=/�9~�(�ϝe�{�
胠p_RJ$T6b�YO#�����n�54�v��w,nT�$�i�+��z�rA�1�:�hy7}�����;�x�D���*�k����i����.o���CIy_��R���e@yt��'��aIז<,Re5�����3p�Sӊ�W�t�=Y�|�v9��/5�j�����V�4�U�Y��n���m���Mi��4e��F���:��[)�l�3��<���ޑ.�@�O5>d���@[0+U��Z&6���*G����n�z�*pXU�� ��fOz$֜�����h�Է�;���Í!�%�U[WO�<qm�vݡ��
��T$8`��㶸PX�'��>�k�ܠVu�X͌�&�M�0�i�r�L����}U�\fD����.�}8��7S,�%���YE'�7UC�1>�U���#ngxںwk�'��ĉ�/�r�9_wr���[�q':����fko�͇�z��a֊j�����'ݶE�sN(N*�Eܛ!��۝��{��nV�:�~5�Ϫ��\�\��%eݒ[�b.^�]P+�ۜ��ө�cnK����we/V��N��Z��YZzOS�ЋXӌ؆��ˁ�`���Ӵ�ؒ�a��є����b�	��i���0�r�f�ݮ�NQ��(r1�on�q5�Aƶf�Y�2�a�6�*'3O$�� .�I)���H�K4�^�y{�:���z(��r[U�m���%3͖���@�����f���}�W�8��C�k�q���W��C�O��^}7!˜n�KIg���=^ְn}�tFj�
H����fy]n�E�<eɟ8���F�'Bʲ�#Z��S��B�+��E���h�d�)��R+1�>���L�"���myrn�[����}��XtU]M�h����ชPVOi�oK�J�㢧�m��y�η��Lu���2e�����Ő;x�D}؛>�E:Ia�w:\[qcۓ�)��8�# ���������1S�`��MPs�jr��3������z�<C��Mߡr�6��Rg[0WIx�H0���wj��s�*Ȉ��Kь�E����.�2�k���{uΜ^s&%��҉�����k�[u�{AA���g+�����Ư�]��7t��#�Q<������Q�/O8�0���5FA-5y��j���:�֔Q�\�]�����z�yV��32�gO�Q�ɛ�ZD�mo�^To�L/ے���3-�k-�،����}L�M̆��Q_�:�M������`�0�5��B��c�C��Ԡ��g3����"J#�l�GJ_xx =��u��m	�v��I�cO�+H}M����5w�<�D2���8v"tn�ȕ�l������Զ���M�
�N���J T�d֨�{U�3T]tE�g���8��ֵ!����Gr��ӷ����'[)�c��{nk&�T�j'��t���
1+O��j-̃����E�3�ݠb�X�ǏS�q���c��O^;�������e{�Q���g���P�Ria����+�]�f��zZ� ,e�z��C��=+:W���F�����9:�%��:�g_`����b��Ķ�b�8Լc,Y8�YP��p����|[���着�)���UH��,���T!�,�]3el.~����d2��̴��A��Ҝo^�{y��dX��"�u��+����?vj��y�FGa�3զ;F���e���~���l��s���܉�C�Nw�?]kꇥ�]���;������G���,|e�{���=[}%%����	*	H�(�+����X�<z�7'�o�ĸi��v��4�M�79yz;c�ձ��	��=�Ձ�?#>��~�_u��]�_�{�K�\9%�jn����i��Z��#�e�M��hd�V��[\;��;I���\��o섬&��F�&G�\��jfH�p�p�K8��1X��e�R��Ԏ��ۺoi���P�}��ktS�T��W� ��l�l��<zX���P�����y��;�L9��xiRA3]�]K�XךfrP]&��t��"�Ml�o_E�Q}Y}V�\� �0�Jn-X��qQ34�x��mA��n�9�ܨɫ3�1�Y��q����-��h�����Zn�3	UVP��y|B*}3��f�ێ�܇N2��Q�޵�N���#�DԾ7�͝2|�73��A�Xp�`ධ�y�$�0�v	�U��u1pWJ^����ZF%s5i`ݕw��s��ӱ����`�j�,y�Al��큻DӸ�7+l��ĩ��d���%�_�t;�xs;̟y,/f�vR�/�@T�a��N8� �v8]�tZ�~�#5�tZ;��pD��6�
��J�剗 ����3R8�,r�tԧ�ltJ�Z�y����.��RVkN뾷ҵN�����yXu�3/B�jY0e`N����Y�^���ۃ�}n�I��p�8"�����aw��0cZV�.�+��]@��38��z6jr�������V���.#»����͈Б4���9{��r��Y䲰iad0����� Ք��	R°�e�lY�&��U�l�=K%IG�8�=Gu�dvۄ�9�creC�u�$:���W�Z�@�3`}㮅����7�k��t�r��ΝS!�2�G�|T�;k����kT������]Ȫ(,��y`T��I�IPLa�*b�,`E&0�b�H,"�*C�Q�
(E ��0
�� )+$�"�B(J�X�`��	4��AEY4����,@QH��YTX,P��QU@QT"�����X)��A�5l�PA$}�$?��U�����r���Kc3�)��s�m�����l�w|�}nE�(�c��y$�v�L���J��aҡ��u�3����C7$F�xr�����dewsG�k�b���<��#w��4Rė7�ؕ~�`Nu��m��;+Q��Sh��z:vf4��vӞ��}���A4Tѩ.��C�X[����$1�}[�
����Ƴ$�����{4�3�9]�N�o�E=��\��3D�D��G8�oٶIj�^�t�C��}蘒��D(����Ht5��b%�9X��7�=}�=�������i=�l���Yt�vh�P�k^��n�Euԝ�˕�c+�u�,�V[W9
���{������[D�S�_-���w�%�a��7�{oI��j�6�{��E����K���{jxpT��W��~��z�j)��
ܚ�iϨ����g�Ɋ�Wa&��W��TK�7Um��f�'����^͜���ͻ����e4r�w������U�9^��kWv��S�yt���rMlL�z�YT�U薻�Y<y7�G�޺��i�+54U5��<�{ݾ�"�2���y�<�ʹ���k�SJ�j��2�5��YX��W7�����j�b�D����{w�,�3["�@�.9q����J=]7�m"0�-I����F�u+���X?9��M�����B��Ͳ���M��j��r�c������4����X"�TI17�ڽ�}Ϣ~����nP�����F�U�f6��+�M�Ѭ�R0�Z�L�d����n�	���e�7K��ţA`F���77V#AE��ͷ���5pCjF�U�ݕ�?i�(D$�i&��=%{�c�\�>��4�6";l`�#/!3Mb�ٝi����+��q4;MnLsYU ���������޷PZ2|gټ&Ku����G�u�/�z��䇖V=�6���0��%GvI��R
A[���<W�xc��Rsh�©iN��=�b��2h�7���#�)Ήa�`�0Sfv特��yF�%&j4@�=�ʯv�k}�Į�Ҭc�u5�gkV��ח�y�����u�"DoP1<',����7�/����ځ��q�;Z�S�c�o�-~�h[��x_d`��ɉ'�=z֦�`�ÝZ�!^t��4�p��Tu"����k�MX�B�\��\YD3�e��{��9I'����	MY��$F_1'��v��z;��t������B�;�9�9}�kwf�H	��񬚒���u[�q���Q�J
��Rn�.����J�;{ȯ�<����n�|�t}7��0���y��H�b������^���:
"���CJ �!�q{�7UЄ�Ѧ�g��ȋT��BTW�A$�~�L�Z"�s+kD��'���[_+�0N�h_�0F��2t�F���B�s�*^���i9⡫^#cڑJ�~�1�ǋ��Q3��^t݇�Z@T�$<���V��x�ls���G_#x-'��5�>G�Fۿ�_��(_^�!��cMp+�{=Ӓ8@�S9�D0�^��r���*��/m����H�G�(G��<|a���}���Hi�<�a�gZ�\
��2C��Ǝ4��E�~�����YI��yh+����T�F�[W�o%�i�<I�5����:��et65ջ3��K
0��vo�M�Ne1�1�ẓmIȞi/��{-i)'cc�T2d,�����ݕ��*���ޢ�(���]̰ύ$;�4v��03�ln(DǗ=۞�l^��Ha�
�����9�x�7靇�cj�`2qjmd�ӡ�Tt�X#����Ɇ�q�]a�^�������a}FQ�HZ��@�P���Ě���$�_yLW��j���1Ǐg�Q�3���zSK.]T
�eC*���q̬b�WN�b��(�0�Z$x���x�T�^^!�Q��[_��0����\8�r��L,$S�����(S�v�����͒r�=�z0�c�*�Ak�!Z��5x����#�刉ר t0�ŷ�}j�H�n�3O��U�k��d7KsY��@vXjA(D��O�*�Ȩ����J��*�\��� *���g?#�r&��
3c���_��c���D��'����C^�h�C9q��:+X����V�����l$�|�4��/������r��T��������w{��XY$v.>��Xt�����C^B�&�u�{��?��,(�˦��?Xj�W��ۡY�)[�#�ߌ#2=-"B��RC|��a�ˀ��j�Qy�������ŭv/�M(XH"�0�+s��ÃrSK����>Q�����a� ����s�>�U�o�`��J�!ާ��yg*����ٳ/��ӡ'��Dq��h:Vl���!���⍍Br�>����v�Yh�&Ay�*V'x|x6��{rP���}^
��]��w!?2�9͌[�-a�ҡ�lB��l�m�P�M�����򾯾!E�~x]�Z!��O�ő�L���<��l[�'�G<���ȑg�x�F.X:htz}m�U!Dx�H����}y4p�j�YAE��^6�u]ZC����Dvư=1����5~a�Bb���r1��	��M���������aMEz�[�0������f�ѵl&�i�&�'���z�x�i}��ڶ<X����7����Lۚ��s�\� �İ
����Xf�/9�0����뽝�~��~'��-6+\"�BX��^�^����d�!�S�Z~��.���$���׬�����ک��9�!��k�qW."CKAKH`��1i��hY�Y�+P���W+{�ݭ��`S��f��E�3���b�.z�6Z�b�g!�q��CM�ٙq���6�שL���6J0�%|=��o5�t:8�Zt��4�/��8i��v;�B��흃Ak��0��P�ו����l9n�c��*�ܪ�e����ȟ"6����HY���F<w��|L��r%��D-��,D����I	&����3OCe��G��VX,�@Q�04��V��s���g=k������8�)���P�#iP � �����W�׫ ≿w'ӱ7~��E9_#� \t�a"�3�dw7Y��ŦZ�v,��:mN);��Ĭd�df�)1��Wd|�D�*��%H'�.FE�fF)ͩ��P�V��=KK�ş�#�K�bf�!�*ݞ��/m��г����~T{�
���>� k��SKf�u{�Qk�����2c�܅VWc��;k�ZSl�,�
E�ާ�:QiH2Ls���W=�ȧ@&G�͙��
��1}#��/��e��r[2nye�ě~4���T	��(�*������	[�z�)�ݣ�oL��r}kO���}�G��*��,��������<�#_[_s�S�f��t�W��~�q'�88_]#���5�p�Y���!�R�' �U�nz �i$��Zx�6���a�M�9C�j{{����B��:djC%f�ZH8g�G��>Q���9ߤ��L_y���򗈘�!Y�V��L+������������F�0`�ѽR!{y�&���H����b��^��~�>pד=HC��"&�4"NVb>/ۣ=�|�^�˾�y���{�`h�E9��u=φ���Mep0��D�"�7�*5�Z��/.����nI�*�Ο!�3v��Ҕ�\� SU'a�����BXq�����+lJ��r���F\�nn��S9�X�� Ӑ�������(�@̩>v�ӥ�]����6kTk���3O^eXT���v�3y.)���hyQwS=�>V,����U��;�Mw���5�Y�ܺ�rƍ�5NQ@�9�eM���s��J�H��y�JX���f���\Z KI�"__����f�>FT;��Uq�t�J��2��Z�6K�;f9�wb�^O��=�Bn���V`����%���dH�������5HXY��sdʾnw]��ȱ,G��]�>�rWAV�aȳ�Ci�f�5��4��	�Q�����ߕ�M��	'��7#4��{�j陮�^w
�|t�{s	��e�-G+
;��m�U.��2fk���y�\�X��_^쥵�Yj]�����V���*���wf�Û�R�Tgg��e`G2\���E�T��[����t���0,(Y�͌a�y�dC_=$��OL�U��.7�#<�O�U��cޓc�Εݖ���R�/��e�l���4^�Kә�n��."��W4�Tː�FZÚQ(�e�NDj3x��;%�]B.d�YD��>8pҨ�j5}�;m�OmҬ���ԭq�a��l+�#ZN�Q���ʏ4l���{_&k�P`�c]�ۛR{����nT.�\�N�8ӏV���>��e5�FŠb\sY�q�
�ਓ����9[���F(��d�
�
�V



 �`�d�P�! ��Yf2����+!R, �UE@�B�12�LI-�+ ,`cs )Q`)XVi�C�EP�J�����kl�d����W`b��Щ%S*�)*�,����Aq�L�.j��Vm�EX��Hc1I��ݗ���������[��	�4Cܱؐ�9P;�$i��eH�ׇ�v��O�߭���Yr/$vuC���2B��QK/V���r'�"|p��lX��*$��6��~
�W�HQ9"C��>8�uA�,�龷F���]l5��ӷ
����k�Y�y�x�_q�C�0�ߤ�-h6�|��y�p�?+��'��z�Bp�m���ֈԀx���1��ƹ
��^
r*�/b���V��Ry�%�J�1Ǐ��,HP�p׵����쮱�'Y�j�D��y!�G�|l�� e^WD[[4�{��Aj�;�`��҇
'V�hF�'�}b�B��1ßw"�j���:tT�R9I���E��yb�M�?1_<������8N�u�����ϵv��H�-���V��7��f]��<C.g''��C�T&\�.�7���[�8���]%���_�ꪡ4���E����-��Rކn�H�IBH�*����}$��T᥏O�}�n)q���9�F���Ky˚�*w���Ƚ��c���F⇮�Em|B3���PQ$�����;�)Y��",r���>T�jf�}�B\G�D��Di���)2��.׋�ˎ:UZ����;��F�a�#5,7#����J��4�)��ON��W�
.>5�ň��C��b��S��h�Gҝi.J��h�p#6�F�a;�d��r1x��ݔ���rF�_���ҋ!���f�k���G<Vg���͘����H�ΗM�l��!����%\a�w~�U���>]�鲥�"իu*��c;��cZw��:փ�R�ѻړ�P��=�y��pA��8iE�pN���:�X���s�*�$�χ�\�vz\>#�R��&,*�0�n�^�A�4�/Ǚ�X���.�g'ʖ0b��B6�$���s9�P��St9�G�yW�bz2�@�~V�^�qz��-#�d���/�8�3��F
W}b����҃��q��~�2�'���Mr��z!ָ�Dv���\]V�YY���6a�$BQ�1�p�(V&e�>)@p$�[�+g����H�!��H~B4;�t������5枤ҽ��)x������$��Q��
��B�a��^�ǃkw}�4����6��{HS\D"�
&�+[Ӗ��L)�{9��f&Zt6�٨,��!�F`Ab�^�+�yN�����fm#�;n�ފ�E{�>2F�ڨ÷��`o 2��_�Ƙ8Z�k(�R�ƯJ��Qɵ�w>%v���4]�ІՓ��YT�Q_�Wo"�{�Wyۑ
�����5I�G��H������#z�вǔ4�9_���s��BW�ɄS^[�n绨x�7ѓ�V��|�����2rhV�F��������D���./�~t��=���b3��Ѯ���Uт�Ơ�{�ڿ���}د�FZ��Y7婮⧄��_�5V�]���re�b��b����2"���� �ݨ�&#'����	�x�Fl�8H=��Uu�҅��F辄`k5Ǐ�C�!�xE��yKj��ҋ>Z.!����pEz�>�ݖ����u��˵�� {�s�M�Xx�C\l�6E���}>�Z�E��F	#a���kb"ޣ����$�VK(ڐ[P�2=�Э5q��7�7+�+�fd��ђB�w+����Δy�,kEI?}���j��A_��@`��$@:�y�m�MJ����.������߾m����B3W��H����ZB�j �3�o��w�ѓ�԰���<x�(�!Ӧ}�H�{�-���P�6��ia�F�)�)�T*0�ah�aT��),12��E�$a���Hf#�E�yqh-F(Ůɹ�=�,Q䴽B�"�7����1Q����uX��:�l�}�Bb����1���4����փ/�k6I�����tM*p(�(�2����C���삄���b[^|�>(�.2/�"`��c_l�����C�O�e8Ml.�r�(u*�G9<Gj��/o,�[B�����3)�<�]	6o�6;�b�j���zLO4�Z�R�U9cz��H�F��W�`lSe�e�&'f�{,�(��q��+�s97"�W�%��u�r����D��5�p�H��+����}�E�"|�;4i!��+_��g��n�V�y{��DH�h��zeg���c.�m���%��G�@S�
�	�s�|wޛ`aW����p��
��K��ێ�VL�7�5d����yNK�6�#������d�w�7�����w��OJd0����ؾ�^T6)q�Z^ iU��C��xuZ>��3�<kP�r��e|�!�_/,�/�a��;�0׫���VaI>Z~�c�4+,Z�|�����r���Md�;���7�ěԈ��(ӄx������,Ι��������z�^�~�D����Z|�E5
��r-7�E(�s�J��+���Y���5�KU�^,�����b.*���Ԅ�<o�Y�e�Q�me�ijR����S-�FH�s�_oC��	֑Q�P����1�az$C�^j��De�n���/�'��rrb(�@� ���خo�m�e�v|���?���J2��!�f�|�"�Kn�i.�����n �^�!�˱aN���
)Ⱥ��ա�g{R�a��t�JbqG�P�^2�����;5.9�zN�c)|������+��`�����߇�����M�R'V�b��8`#Or���D"�]򙌩m����-I����pb�Ӌ��C��l��r����va�H���>�놖K��SИ>�\�^ڽ6x״ý��Q'x�<�ؑ�c���ZF��//��i���zS�%��@i�S�OK��w[�C��[�����_��馦S�Q�[HZ]��ۺ�g�66�B't�JYu]2�O0����2�ܓ���2M��1~�?�㼑�!���K/�\�Ȭ��c�y��j�R�OQ�C�CcQ$����;�&h���[��A�{����~�H&z�p�0(�7�}��f+5�~0/A�\����*�<D6Qx�Zg!��%K�]��}�z���gO��AT��D��!'NY�f���|��G9��e����
W�|�0�����K�}/�����Bl�F!㕌�exի�� ���M9���֤F�{YKCSfb,@1>RcN�V���
�G��{�|�׵�NN�H�iH1]<Uz�LoH��/�7�G]߷���;���	�B���v>�����J���z��҂~����݌B3�f!�w�)�v��a��]SW�&�w��zU�I��7+x0^��c13j��˦ħ&��C3D��A��3*�S�����G�I� |$�1��.vϱH0�z
�e��uJy[�N��ƍōy!{��Y��s��ظ���=�ro����G؇��cnH���MN춨LGE��.o�X=@ab<,$M�Vi!�y��^���7���K|�s墵�z�P(�(�J���p� �[��;��#	����|����y��;Y�j�;{�;�/����y�xT6|x���hF0�5V��:����ӻ���#�{x�Dڨ��/��p��؄==e�Y�׾ )�����mȼ���k$C^�����>�i���-\C��Z_ �!p�([�4r�Ti!���Y�KI�J�¼Y��I�b�I�����%;�J�1s_I9���J�J��,�w4t.��77t�e��X#X�|���}ߡ�sf���9�:|E�Gȑ����a �(�黐��%�w�����c�k����ط��W����7u?]����JZaG��?��툝�������%7ײ�}��%�z��l2+�U��H�C9�<Gdva�^�m^nv暴��i.��4�������ў���Q�}��Zg	3)٢H�P�|j�Ay*�L�ɫZ�b|W���ӀȽU#�qZZhbd��2�MBN�d�Ⲹ�>aNF�k�Eu*)�)֧*\��V�Ҩ��o�8�T�:D��o�6��t����t�+2d=m�I�d<�u:Td��X6��h�B�Ut]φ�~hv��u�S����9Q81в�J㖛�Dok��Au�v�I���٬��s.H��P�\���.<�ʲ�;�o�TqBzfM6���=�9C>���e�r�Z�m�J���
�̥��s���0����B��*мz�\�0hэ��[!]O�mt�ؠG��}�Y��Ea��3��k�ӡw6�t�홓��:Wbgh��`��eu��;�o\9��Nٚ�,�T����n��(��Yu��|�.�U�,o��0�3���`���[v^5�2GuhEV�v��D.��Y$dcd����b ���S�E��,	�p^�C!i� �Q��ޗ����ҷ+�E�e��>��egVwu�F�UT�@�E��G;/iμ!Ʈ䳶,��`��r�ޫ��T�ˮt���I.έ[b���o��X?]	h+Ҭ�7y�^���#����K٫�Rg��Ci*�U(�^V3 B<�^2��WGv���X:����f��L�DA{-D�4�ᕉ�@����U)�}78��+�uY�}������3�����bE������zb�b������V��0��q��N9B�8�CWNV�c$q�y:a}��2��&qÉ��'��^����}x-�zmN	�I�;T�q�%��gH�u�2�\�]ỳͳ�r���+5��󎾬9�k�D����ǡ��q�b�f[�W��ux˫�"du�K}17n�ub@y���1�2��3u��r^�IÜ��%�6�}s�l8����5d$����TND�j8Rr־�l��}�iY���PA�s��Lm�G�7�L��2n&{w�>�W��k�����E�z�1��
J��d1X�Vbc �J0*T��0���
�4�c�-�QR�@P��X*$m-�d�$��E���Y`�2(�XJ��*
"A�P1�E�1�+"��
ʕ��IR-`,aKAF�V�J��-�l�YQn�.Xز-V�m�eB�54�"�Z��E�+m�D�C�O�����I���ў����z�:�em;�[�{�7�q�"'.I�T+�\�s����C�@���9{mNL�ۚ06=�0>f��sɧ;�n�H��1_ԏ\�B��0�"���b��n�k�a����f�C���zp��͠�f����Y*���GL:�X�٨��j������x������ z1g�7�	=`��_m��L�muv��P��0)}�y ��a�(LD�"K~cٗSsk�0�P�_����(�!\��x��O�㷺�W�
��w��E:x�Uk�!����#v�P�T&.�91��҈�eFŜ��It�!�xUa|׌����\�	B�����3ܘbs��<�!o@)?*.=8��*�Q7Z���)uz�e�j%6FZ˻��87��()<J��z���w:ɂu�b�L\�խwYM�U��\��'��9�<��)�F^9�b�����s�0�?���]>����V�"�����n��frK�g=A{�C�9���q�x�1�'�-��4�/D:�J�u��[]'_|Є��!(�S�`�w��¼a�W���|�P'��E������u~�Ю�q�[]zx�0NИ�&�ψ���%f�4���&���z�v�{��,�]���1�紅 �!�_!xY8aF)΅�o{��������8�d?.=Z��B��P�r��i�:�db��.�s�ю}p!�P6�����E��n��ۻ���?\G��e�Z]W�P�~U|�0�W��wV��_,��H44��i�z�<N �{ץ8�/��R��	b3�(��X�6�5�
�e��gw�����0�s.,kv�Vr�5�d�ʎ~��i�����.��>�d��Z�1��ZVG�L)�8�/$��m�G�b���^�U�t���^����n�y��HLc5���b�Q��*}W&6����fw|[�t��Z���H�`!�}��rg��8�,�V�Ӣ�@{\o�&�CޯN�
-�jT\��a�z��<�9�wJ�Hx�ц�Mf�hq�s�b��<��$�&8('��Y��.Q��g�S�8#�g13Y�zY:Y��Wb�\���n<-"l0�79���.��+�Ԍ��5��¦��;Pr�Dȑ��r":2D�ֻSI�A�6F��O�q��|�	b<��!�O*4 �m���kE(�xD���������o.@�Y��jN>=!��kbco@!a�l��鵑jǏ�E�&v(wvjN���
o:�>K�+3Q+��������c��bp�\x���hF0���C�/n�|=q�^�����Xt�������<���a[����`g<�I~v��N� ��cu,�!�r�E��ZfA���(��ddDF�=��N��� �)[wYs��(A�8�xj14��e�d�$*CJ/ء[SO&����sP�H}.'6�
wHA�Y:�:sgL2�G2���|̉/W�bg���=\�[/�O�,��_OO���{g�u���!�����R�=O��Q���V#�||dP;w����V
\ZZm."�1�ǎ|~ȱ!�z�{�v��u3�������3X��VY${�3���Pەz
�=�x�Y�w�1^IN����e�N�=^5�c��m����o�Y�S0���p�v�O�A!�Qݜ��� �ū3��&��[����������^�B�P��+KMbe�}.���s��(�*�4��C��	n��;�r��k�H�fr�nw�'��c��O^��8TC�W���-��B�#����w��j���פ�ud�$��h�(ᠣ����ㅞ=9顙���ǐ	�F����	(9��9�B��F,߽�ɻ����c]渚^/�,D�9��i�<hQ�F��o=׫�dN-�E{�'*)���S�@������z,�Z��Ƞ�F�68�!��1k$X:}��=��.�d��ST|F�䊡��jň�U{�V�e�M�<Ь�b�^[��/�'�@�(�!�	�H_��в�=�ڙ��J�{w���7
�t��>�۶#��i�$8�M�\���4�vJ��-dĺ����Bm-{9�g�%�'�x�p�(���=p+�k���|��k$[��w�*���Tz!��<X�EX�6at�����8��NM������6x��X}Eҕ�x��±|e*Sٲ��7�l��z&3�_�^.�b!o@?$�� E�\r��Z�Y��2EN@�#ki�A�G�U�؞��Cm5xw,d)�Fv^�EV>5hs���_^(~�VD��r��-a��HfŴ6��|�ʷ4/�cU�
�u��o��r���$���wD%�1{����=�7��?{���FKK��x�$"��an���@�Z��-`�aK�Ά��r��O��Zp�L��#���f_�ړ��GvRθ)�ڡ"&��\�տSԭM��z-wL��s��Gs�U�k�����u��^�:�iG$��Դ�����u��8���H� ��ԡ���xY><:&����w7�:�^n��V�sHq�Q<{T=�C�i�a�~�n�
�B��Y?�mA�"��z��Q�ǁ�U�ԥn��
�H����vв�iuR�r�*�`�"f����[������ɇ�x�"x]	t<)�)���^�=t���+�.����@S!�Ta�yiZ�%��}�x��=�V���U�r�҇.�O��\]�0�>Ե^ص|�z���f�~���9!�U���W�vo!f����T6(M�=���c�c��[=E��EU{<Y�y��!ڭ�F�����&�Q�c��	�T.�_<�7�2!7�6�Q��r���b��d�m�7�D���N��o"����d�My���;t�#���ũ �{�W���]�<Y7��b2f;d(�&H� �P2��Hbͻ�ӵ��h{�5U��w&�Xa$o�;��j��xO$�~f�u#�S�ѦP�@����N�C�^��;�㾌/��O->������R��#B+��y��\�96$d_K�!׺�U�8p+vj<x�:Ym���}r�j��LH��H��x�Dڻ��������n�ʹ�ѝ�4����J���l��ckY��['qyӦ�y`�ѱ��H�pȂ�H�i��n��ٷ�y�'��-�� m<x��bi�X��V�%^��/3�,aM�E�����c�z�B.,�c�B��|%��`�g/����FVW��ҷae�Uzbw;� ��Ʀq�󇭣E^up�E���^>�W�M#�\2��'t<����<����>��U�q�>�?��ɍ}_b��>�%3��������}F��
�jM�(s�f�rǣ���-�=���lQ�N�K�׌i���"�*���rV��K��������8I֨�i>p���X�d���w�8�}��x�ˈ����s;���D����rm��w��)a�}����-S��5�C��d�_v��6\�~��Q&F)pۆP���f�8���`��M�v{���Ȅ�$���<���_����)q�t���-���l9��:�ȑ�� T�t�N���wB���-MzoޮS�4���"O-?2x�+9gqxJ8��5l�p��%��'E����.�w[ɷ���S��ܝ���xt��,9aW[��`F�"���9�m,�$�)o`q�ЮL8�&qQ��|+�7�����hp��c�:D圇^kDi�Zlm�*�=�o���k��Bύ�P�HTD�^�~�D�O�]/^�M�԰�	�K����O����"y�S6���>����Ag.
���/��OʏW��E���$߳�۾��%�8�+��P��Kƥ��A�TT
R�ebqұ$ZQ�(��(8釠��RC�⅊��^XF��]�η&�X��
k�(b��Rޚ�t�|1�c�,�:g�;�V_�8|k�
�
�ܴ���d_�^��l_U���"��}Y-R���*r�#k�I*::B�^sa�����g4�/���#z�������;�x��^7b�]Sq"���B��%�cYrk��-K{о���v:fW0�7Y�]���b!u�XZ�v�e��Lpd�'v\M��x.DjeWۋ{a� y�Of����|��_XVNu�Tt�b����,����޵��#3,���k7�Z|��*���
]�b�;:j���,�i3	|f����{|��;|�P�Vg[�Lf����Y������|(�j�u�I��tK̮��7ź\xf,z��:2��XYl�<��Q����p����w��suڌ!��H�|B4��-3��+f�����aޭ�Ə'yz�W��m<�vMC���&r�A������#�{(�h<{j��Sz�@�L�cr�S�+��T��%MZ��j���Nm({u\��a��Ux���d媱��8:f�H;��G>G9d�yT�)n�:����U'P3pL$�Q��7�� o�)��vUr��b.�3�
�N�"^���l]�Y���JY�T�Ewt8����\6��MK�{u��YN��U�5P�̻�$��AW�U��/��t;I�j:��d82NJ-a�qG�j}��{����>A=9+��$9vJZ�6��M��&�6��cS�GE��3Ɇ�H@pU�L�L���{	�D�����麴F�Q��� )ݗ��+��KF;�YwPSa@�]7}LdR�ܡ@^�d,�|�T�})Zt1^��Ш*���/�hN<{C-Q{�U�l�'�;i�&t.Nی��[�f˂�p�7j��1H�(�+/-V�<�EX��R��K��7z��%Q��;�u�Xg���fh����w��b��G�!��o]o<�^�ZD�X�-B���E��ڰU��V��ƈ����Z�ђ���OiMj��Г���P�`��X�B���XW�UACVb�KIQQbV���%n7�k��XcP�,1�Ģ˂�1V,��e�Fb,QJ֢�bc1��p���c���q�ֲ�%q�Z�L�QL�q��EˉrX���U���8T�[lf.Xt�5ciU��J�-Em"�J:bֶ�E��
֥���	g�IE�q�w���J��|V����RoeM�s�9.����'~���L�=c���'
|F�B�ʭ��*wy���(��=A߶�q��CQ6�����!��p^隑��JLἿ�HW1��e�}t���<F�~��9���9c$Y�f���[�Ŕ|Grӄ�fk�tV�R����U�N����0�*h/���紅�肋�vi�)}��=��~9Z��)U�!�L��ǫ�p�cy"�U��|��غ����i��R���2�(�XO{)˯M� �f=�����g#���1i��,r�*��I%z�Ӻ��ei���'��"���0�W�'���:Ru�!�9���C�S�\�x���C�ʣ2��G��y)���-�YVll��%���]G.[=g7e����pN�n�'5�Ɯf��^^0���`N�Ҳ�Cn���&'>
�j��|	��A�c+!��D� f�l��aE�P�˞'[/|�})�ե�f�~5�MH�@z�w8D�yt�svƚ�:��R�+ꇌ'm��}�eKKM"�u%�<�om��%�uhC��T��G��j9lq2�5�k���u�%��+K�tXW��u.�w�C�H�&��J�I���,���W-��M��	�o��r�3��˞�ʦB��8R!�I���wF�*:�w���u�A�^��MiiG��q�x�a���)x������2g��xXC��s�&X�|C�N<x�:Y�n�*��������x��C"@ח�HLS���.?���q����
����<O9#���u�����,R5�C��}���.��nEI�j3<2l�$�m+=�<6�=�M*�ڸ�;�*���LYZJ_�x��H�p��j��O����O)
�7Q�#*#���9k�s64��!���*�"t��7	�{E�����P�+�$�^R��]b�Al��_�,��1�`��0���n�Z����\����U���޷�W0�3�
G��M3����۱�ħ������&�a���Z�}�I��CH�R<٢����Wn͞�a���C��Z��Zm.!btr�J6�\���w�/sa�|hMp�����8Iۧf�#��(�/�����Z��a�Cc$�G�sm�p/�����豳Q.�ǘ�)j�N�MJ����F���6t�:�r��D\�\:�~�Z4ݓ�ZJ�U����A�	��u�oNJ�i��Y�L�uq>��Jh0
c��hN�հ�)�q�=�s��fb���ͨ���fFܞwtm1�c���N1��:�2��=3h=��Oqc$�޸��8p2"D��I�e\��q�kĺ�^�RM�_��˪Vo՜�da߈���u��D�����*�������ˮ�fa����`�4�@�_Q���<��b�C�sP*mH�1�0:	���˲���Y�Fл\||slBH��C�j$yw���p�)+DK W����������ő*(�JmNo{���くc���������Q�
�(� ����uf_��̘�O�d�C�^����8aE��.��S�E]I���G�['�C����C�V"G���WT �'a[��j/;V�:y���-5�$W6]Y6��I�L�8��@sYLt�#_+X��H`���]����δ�p����j�řX��.�츗q����efI�(���0���Mb���0:*���*MlK�nݳ���*�>���C�Z}Q1�@V.�>�^&h>Ю�d�Fb�Ct��T�S�89(�+��Ҹ��Bt鯗�/�Xw,LD�;P,�F_R���΃�e��ۛ�:u8�<�-YbΟ��:�h�ˌ�-��z�gS�-�%�p�����V�a�H1�W�9~���U�ÐN���Qv�ӱ#�C�-#ZL���<�
gS���R��<�EDÀ�����x��hl��qUfȾ@�k�ڍ|į=��X�M���=��V�H�Դ�P��m:�z�MX��	rߞy b���̌��8Pn*��Ծw�,R��˭.4۸�Q���jP��ù���Q��թh�Au5��5�ɝ� {��?UUU;&�z��A�f)M��=;���A��j�[|�$�֚1PЕ�Bf8���l��e��꺅r�*�Y��=���{�t����!+Y0���Z"L^N)�n���N���eȼ���B�0�*�O�xÿb��Γ����z����F*��/d8w��܋��D�`��T�1�--�I��x�9�u��;%Gl��1Y c�IT�j��^Z�v���(�#����(K�ޞ�*����6hT!�JJ2����e�̎����MN�Ø�o����7#a�������%i--cE�CŅ=b�ޏ"7ʶ�rM!�	�}7��1�=���q�i`��2��uw�/��g����K^�V�P��� ͊�V�ݷ�\"ZuY
����(��u-�V]X2��x����}����� �zy/���Ȥ�|ƪ:d�M�������
�
��}D�OG�� o�(H:}q��8ҏO�q�oː�yKH})>{{��YЅ��h!"&�||C¡�\x�X��/]zwBϚ8|x�5�x��<P�F���m�b>���$?g�>0��!辄�p��a~�ˮ�K�uI�#i
3�K�U��B�6���t�(�4�6}�������jlp�\�_X�0��u4j�_+���I�'�A�1��>7��ա����\<M��=e���C�W�CV����EyCX����y��U��v�;^fn��z��!>�}m�\�cp�*��F��;�蜡�}�йh4A\�k��Vi��rW���~G��lv�������@V"U�� m�k�7f������U�}(�⦳t�K��<<��$�S�(t���9�˫a��ii����i�]�޻�.����Z�l0/�ƽ��U�p��Qd��מ��F����e�{<x��e3�*�ɟS��J>=��Iݧ�y�˦ZI����a����׮r����h>�O�������h;U)Ч.�����E��c���6�0���!���́�Y��$�˔�1Cj=����H�s��6r�;�~U�p�*��6��v�
zs���w�q&z!4�#���9K��E�O,?0Y���d�6!��-q�$F\g�:D圇X�h�h��ws=��B�|n���L�a���BF���hK�d.��W��;��[�_2��ǥr	���Bi���w{���|���5D¦�����u᛽s���gR�R���x.�\�l@�;%��UU(~ィE?0�q��o�����O"_�A_]����T"��9?!���@J�父�(؎���tOk�{.��<��>��-A��)>K���h�^H���q�8�ǎ�{w���b�+�3oi����D�����$���zk�.��c�`1�޻c��zN~NFv��޼7�6��2��\D���Ѯ��+��V����V� }�Z�jK�k���ñ�J��Nv���]��B$����TD�k�V�?0�â���v�$�f���8�J��P�ZC:D(��[D��B���Y^���gg=�{��T�{(�$�8xvn�[�eu����s���.(��!�<��i�A�Y����g��wV+�_ԓ�K,v�֮s9�:1\��=��n�����s��C�˼�-#C��Y����'NĎ}�C�d��|[b��\�M\���1��5=ˍ�g�u��˹W����N�$�f>4���	���<k"���紅5�(ݝ�٥���9����*�6�2#i�Q��G�̻�r�o�7#O�����Ÿ�V*��oM���>��h{����N����|4/#�#��}�,��K^�3�ߓݺK}ٽ�mK@�A��q�zɇ�C�����N��F볋h0��)���9����S��1i-�quwt��X����ӕ���R��!]��U��G՜}���������a�|�<>��C��B=lՠ�b*�����}Y ø����yz8����d�9�D`o]g��wI3����IUq�ܪ�8J�����zGZR�;��(��v�05N�WƂ	����e�>'�Y��%���IPȷ��xDH�7�S�γ�2*��N�N�����R�Z��ki�L�j��#�a�Ԟ�΄A4Z�1����cRV���q9�0\_��f�O-9�+\�]R&w&^s�R�K��R�+�4��­��f�w1[n�4��H�K�AGY�]��{�S"���w�xRv+��<@��k<3�Z�� �ջ��.���t��^�����\�q���Wc�.�ȷ�G��d5���)V�V���4�ʺ�y�z��X�:�)�f��&��F��$�r���ʬ�N�tr﬜�ٮ��Ow)�����^��".���s䲩�r"R�u��0b{��M>P��*����:Aǃ��"��%5F�SU���5]uه��u���,��W�Cb�=���Ǖ�W�ٽY���ژiZ�ʦ��d�[�gQ�0�B=����*�V�j[=/H��.XF
N��0�v��U����/j��z���CI��ͣ�(�1^^��=�Ԕ-ie�s��vܹ�'u�r�CY��)��u�O%��U7t2��m{�V�Q�8��Z9f�Tf�S�퉈�85��Q��c����Ĳ��Κ�YԮ��A)nEA+�a��']#�J��nA{cLB���X/0�`�m�q�]a�Ӳ��� �3�Ȓ���#Q-��nI��LP���Jͥ��)s@��C*4�"�N<����ɴ;)�\O�*AVڈ=�1R�c��5��K�r�ؙ��. �����1q�E|��
����SM���D��D"�G#^�^�T�Tam�%TY1���V�CIXf��i)�Y�*Ƙ��j*ȍn�8�4Q�$�34�����L�fSB���h���\*"�k)�ێ+���U��DAeJ�1�ɓJ�et�V5�E��:��*�ikfaq+���.�j�Hc�Q��:qs.&!�Ę��\%�Ylr�����#���QLe�j2�Z����L�L���ޞ�3{�v����cX�ˀS���;��\�Fs3"�LnN�U}U�[6l�N��?X�/�0�+�Ak��ʆԘ���R���r�l�Z�%�r6;N�|o����	#�����������G[Xj`��iQ�2��Ƚ�o������xڎ>�Ѯww��=�`���Y��N�Qf��Ȼ�	|�E�a/����+8|�����]��+ck�!�W�R^�䗷��e���qh,=Q�x�6����oː��z
��d���!�!hAY��C���]c�!XT/���T:�)7���n><YDJ^<a��h9qi	���NNX�E!hI|�Js���FL(;�o�����h�j܅/{�L���|��6!<�#I�B!d��H�Da��ؖMn`�:m˸wE�4��X^�Z�]9�ޜ>�hQ��ՔxB���$�o��9�rZめtqd�e:�L�܋qI����£��Q����,U]
���%q���ǈ�F&
��`�U�����2aiHq���E�����u���B� �]0���6x�Z��V��|�� ��(k�L�X��{>ָ���������s��>�|���T��k�4�|�ѱc��o��H�g�sa��0r���t�I�jqH���h;+5�*(b=�5�B��X��Zf��S�F�]��mB�'�9f�ڥ���X�Q^�l��2�^��BT�K�׻�m-6Q��>�a|�$��󥇨{ް0�z�-|���ǹ=�/y��$+]ʗ1+���A�>#�(��p�aBj����yZrc.��x�$�I��2P���V�~��2��³�qY���R��N��#�6+^;ħ�������,ַ5�6QWJ�F�RR��޻�"��wb�_aV�z*�X�^�Rr>X�Nw�7������K��da��C�"�<j��Ǿ���ǀ�Z1]a3�,�b�|<e�=�i2�2ኻ��p#nw� ��Da����=y4)�a63-��#�<r�1#XU��G7�"'�B�D�GR2�<*��BHa���ꚳ��*v�T����3v�)��k��du5�Mh�z��V'�ąO�H�*��n܌��[��[��g	�簉��F���ꝺy��^;�a<��(���dov��7�96ct.�T/ѱAW/��56�L6�N�j��W+D�-��]�	�{�WYJ�B*=r0Q�A;�[R�����qyD�W��i{�JU�3UuVs����p^�R^RC��z��S*AX�}��7� C��t◽����'f��|jv@�
%����YQ�������4�f�b9���,��LOݚ�lM�I����0����m����KX�Heªu��22'L��n��i_�S���|fB�?녩��3�y�K�FX�ܢ�]�:kfhtVK�9����I'KF�n*����kGf�=������|�rc�)uGx���+�=ˬ�[���5�BQ���57�J��x�7HB�W;�;JZ���8�����K���k�g%GvsZM>ޒ��7���&ܦ5���8�Q�I��4k�r輋q���*j��-��.�"^c�H[�vz*V/��s��Caw4���n��l�yc����f�
�x��f� ��n��t�k\�ȗ�VƋ
'	�D�S.��E�$�H�&�ͨ��iI+�������2�P�4Tѫ�"/�w�M�1P§�/زV�''�.9|k0ꕌE��缊C�Yx��s��Swbij����)�QN�^xIh|5Of�N�2+�.�,Dh��yy�OC����j�ʻ�a:�az-�������x����"�<FZ|��hJ��GՃ�\a�����:�R��Q��oW�#�:Ƈ:�M洛-k}0��Y���qY��`�֤Z�Մ[��i��]�F.U������l&�d�k��̃�UW�*�&R,gF,bL�Zrb8Q�P�F�ػ�U�n&�`�ʦ����0c2^4��3y�V�(�gc���z�M2�L/ioe�}�(V�����s�i�}gx�%N|��c7�gJw2w�����O=�'����z��+�=�2� ���2�g��]J�̳AT=��j��q���q��\Y��૩آ�HF�3�F���5�㘦�}ǘ�>�mIȞrM��&�U�Yƽ�"���%�7�Vy��o�j�K�~��
���So��ٜ���Uo�"ےڐ��|�A��d��dro��zm4�YȬ��lFj�On=�q.�MgC��IFh�x�Q'ei���� �,�˪O[E�zo�Y
�ƦI43�}%ȸg-��t���hإ�F�������#���=P�蛘�G�U�����-n׺=F�lH�g���m����x���W��M��SJ�	b;j���՞�����L'��ڶJ<F�m^RͬI���7R����Uj�IŎ.]*���!�ѹ
���:�/x4XJ��8���a*�N��q�m:�_�'ASx��­g����ރ����03=��V�\�G�5�r��r ��Mk]"����F7�S��Q�ѵ=��s�:�S��T���2^��`��6�|'�d�к�i��5�������ѪZ�<7c��q���ԗCz��]Ĵ���:�{aB�������l���_<�̆�ծ�jF�.;�;S,iӖ��։)&d:խf��κ2;3":eD���Kwi��r�Q�laT'Q�z��t�u\�(4�:jw��U%�r8qum��%��6�n˥cN��*K�=�J��u���Zц5����Ml����m�����Y���x�:`b)�"����k��Ӻ�׼+o������[��*�C����O�f㩘���t�-�
<�z�\F�X|f�c���3Re�V��8[:��p3���ĕ�nj��P�Wn�ڛn�:���#�|�\�)��s��}T�{��+�k�RA��+5u/}����k��0GS�ˎg$v��䮚yN��&�_Y{'O"�?�1�e���+���sq��3��@��Pk�N��f�2�(;�lšF�r��EUӬ��g�^�qS5�]h�P�7���C�qn��3���F�:A�sTi�}̔���b"�{��Vv�h��xN+k2�9'���6��7�s+İ�j�K�S�;�Jm�L��{�L.c�'a<��挻�wQ� b�Z�<�T�NC�Re���eWx`��:m@�p���Ǔ;	����7RQӘmX]r�~���]� �8�E�AOIj7�D��e�&�E[�l�8�Dk�N��z�a�v9T�W.j���c����p�m���}p&�nƢ���sy������;ږk�!o�3s$B�}e���Ybn�Z�)6�dO*�!f��b�������Y��v�QM�2뢛0��.��$A�f�G8�aܴ�};AŘ���M����n*T^���Y�,B�QѼJ	N���R�k�:��h��� U$K,<�˲qܕ�f�k㤗2��D�"���fme�KyG�Q��&-�H.4ޗ�N/<艠��Gͭ�Ø�&|�^qu3���,�-��fqf,�^v�,*	M���WpG��W4���b���6�\��B�M*�>�R��Ҟ�Q�8ᓨ� �̇��3n�Ih5:�LO%���P#�t���:R_PUu��^5b}��!6�"�]I�[�	�m��ޜއ]��bP.S�G3A4�M�EN���W"�t5U���8���uD�8�P�M��Y�M�Vt� e)e��R�����\=υLa��`º�ƻp���>�=�o�ѫJ�����6t��W.b�8�[i��w�vu�wk2��JGE,Z�Krqᖷ�5᝚�&�p��j�N���Ψ̓���ή}��/�8ѝ]SR�*�Z�q��L�����5Y�^^��ދl0��8�W�&��vۆ_-��I�;�Lv��������K�fO�a-�tk�#ū�՜�ZN�Ln��	kڇ�pe���𧻓����\��e�ec�V=+&q��I��˵.:Uh��-�0���ﺌMX��v��2�j��]�v�vs]:t�'Vͻ͓sQS��V�2���ݑ91��aLqL�i�];犮$)}�D|J7p�w� ��:��L��dA��*�G�~I|A���h���het�Y��\�X֒��dJآ�4�e&�b�J4�a�l�U��B�[�\�DIZ����"�Z�\��Y�3iS2�Lu��5���c\k;�f��H�R��+��Lj��L�(�8�\�-�YsWn�3U���.faZ�̦%Z#eC���MR�s�i���� �#-���Z�cYm��f"�ܗ�̦eYm�Z�5��!����P\u�i11��_��H'��y��wީ;;p����/��pon���2��(�d!19��-9?{caq�ͥ��zB|���%Mk-���cl��:Uǽ��.�t��Sӊ�W�̮�Hi�ɣ4Ug���*�f��5�^ޚ3��{��Mӊ�ldu'��5�ڨ:�N��^^"�:�Kq=�R��`�X���'������θ�FV"�JP�����U�g`�i�3�3��R-���Q���ʹI����KI�=ݵ�|�J����3զ3z�1.o��-ziwlV`C��_�U7ԫ���^L]#�q,�Qn Q���ö�1�X���.�����P�yzo�sE�t؏������fH��n�k���'v2�g��W��@��j��;�w����ȫ�t�8�l�d����k�2m�YB%[����Zq��<en�o�^-��Y�{G],M&��>p��n�z�EK2�䷊y-`��H�ȱ�Ɏӹ���U��}�a��H��kY��mot�r�R�qO WvUcZK�qof��qv?Όo.X�f&�����}}�)��X��L_Z�ޏs����lc� �֚���YV�L�m�R�qq��#�z�j�C^����X�|��jq �^��ZW7҅\�l3ۦ35M.(s��Z%l�CG��o%:�s���rY���S$���t�E�r.��ernS�'�Bz=NgM;R���e����̢��4�_u<����~Q2Z���
ڑԎ��`M�_�ϻ2r���z����;5R4����F���6kJE�~7<w٨.*^��{ ��x��^2�K�6���NhY(m+�Q�[eM�,D�C��t3qԝ�o�q�gQu��Ň%d)�����ڐZ�H��}�!=�y��
�Y4ȞG@�)�l�ʍnpj�J�۪f��n��0�A��o��}�.�l�R��&��n�-:��_Z�n��_.�d��{ï��l ^�U"#(^��Y(90yоs@z�r֔J���ڏ���Gv{��z/����Dɶ毵`�y�S��Qq�k�E��*wx�p���F�M�s<ur]�Pb��p���������3�N���k[��O���;�(�����3sƮ�z�����mpJs5�ٵ��vw�0׬7B��,��9���J��ټ��)v:�1E������繇�S=��"����d���@@$u�
��X��g�JY���gTOf�jC�DY����&�ԩ����S+}oze^��f}Oâg��lZS�h����břuŖ;T5��I�b�xo\���r5هx�̸�U�[�9U�*��wt-���f,�*����ڸ�{z�1�vO2��!�z�I�UZyF#�Y�#j�q�L�� ą�8��g��cX�s}j�sK!��:���i���G:�6��c[=i���W��
�[G8͝/#���n�������X�.kjJ�ª�⧣��2���^;�t9I�Z^���B{�6Kx�E�W�f�-k©V�w�t<�-y�M��]tKi�a�������0�;h���KS@��[ƅT�-�\%;�lo�y�"�7��a�W�+�S�Y��]\�쾒��*�E�:�(�X֒�u��No8~�E��)� ��J��'�S+}�*}g(LgFT�e���m���=ȶ�����eGj���
�P��P����֛��Z��D�m���L���ƣD�]<8����k3|B���sA.#��L�Qz��m��2ݵ�n�z��o�q�i�U{H4f�x���{)�b��5��,��9:�#��.��=�󩙪k�j�y���Gf;N���jwyj�~���P߳&H
���e()���}[3�7�R� +U��!i�Z�|�Xws�`��7xhMoގś��	}g�9�7�����9���PC��mt������'�&d��e\�nN��K�"�w���ӽ��a�u�C�/ ���X��9Q2�Ĥ~���f����F�="�о
_Qv��\����=*CD�WIɘ8���5���/5#����g_b�gأ�AܝRw��ߜ��#o)�ñ,�D��ġ���sΙ���7��5�X]b�d^��^�]�Rle¨����Iӏ�f���>]��;�9z�j��3����>��گIT`�l1bw+���t�כ4	��[��` �=9XZ'7r�j�=z|���`��{�,�-�_g�P�8�����Ii cP���s-�׹�J�<ov&Ck��F��B*��f���ڞ��N��őIu�V�sp�L�3��7Tk��"xE�L�Czm���*.}Ȯ�W�A�C۔�a3<̻�o#�R�~(ܵ�gfWyn@�����y�-� u<���erJ��zެI%2�b���Z��2���*�5#oE%�G�V'��ǥ�W�:���u�ȶ��̦hح�m��哝���l����޺q�X-�N�	H�9��U^f�1y2�i�����:�C�qO!�	�*z��`x��&��,Qr�X�;J����WB��h ��n�u����-�\R*"�["�jcvJ)���fBӭ�������acZl��6�g+Z{%Z��N{�蟼z���) �h"�X"I��O%�RaCm�L�Iy���	����;)�4�aW[�d��z�t��]l����8�Gn���7J:}�,q�:nMM�&#�wYy�6���A�mX�
}���h�O��˞��2�6�
\Wf�S/��{7�l����n���T3��0���g�ǜ����(Ѵ�+��1(^ض{�\�)�G��7�"���ud�0狗A�v7��L��	�
���p��D��T�'p��d-�Ǔi�l��{R�:"�&ɍ�=���}�ͳ��� �5���{��X=��[�ꖂ�U��]"���8�c��4�־&�i��B܎���3bx=E�Ìp�֤�Z��kɬ�{�a�j�m`aɛ�m��sVѼ�T�9Sѕ����G��еګ�<N� ��-�ϒi���j�8����e�7Sp��7԰��ߗ����@�f�	����̼9�L�o��FlN�3ۃ�o����X�����T���P�[�piZ��	�U�ǉ�H�I�
�wqK%ve_lˊW4���00�d�������k*�
*�Kw�t߬Z�WCm7yl���\æ�v���i������R�M]g'dx�]_~�4�D�攇�R��U,�N�{%-;}uo����!�>8+�x��a�:b�cc��-��ͩ�L7��7����c�/���8���9.�9��u�jJ*�p"C���W:�:6!���{��N&�ٛ[��3�C@k� JZ�R*�SѶ�<�B9���z;;*ڗB���ꒅ�1W �GM�|d99v^�=Z�Ա���r�]�(������������,QF���y;PV�6&jx���0����t�0Qſ-��(�T8��k7:��Еy�x\��1���a$E�2z=����byإ���bgיJ"��pU���w'uz䓱���*v��(0�֫�(q'�e�`�7PQ�]�m�4��me��U��\gQ�3��ҭ�ܫ���4
`�lo�v3��Ȏ�xb��z���ɽ}wb��-��R:�V�`��LK-����}Z7���MHW��6����QL��"���XR����Uk��z\k��ڷ.��)�/-��1�n�V�D�=��9;;�1ʺf\���˭U��hC��[�նL���gSe�#y���r�cP�[��+i�f�;l���_i�J̑�����S7x���GX�lY:;P��SS.��͝rQ� #�F��d-�vxv#������91'�aO��\�n^LF;=�,�N_L�h�8h�U�Z�l-)����y���ʳ^��lf�[�b�V��V�5�WT��Z�Ui5���]Z�h���E�XdS.���b�0rY*��q��C2�4��Ӭ�e�i����-YPR����m�\jQj6f��t��e-[i�f:���6�tk�R�S�]%4��\(Ыu�d��nJ��q��h�-m�bŬ�1��b��.�f�i:!:D�-���U7J����i[�SZ��[S��\���@� ��+�<���9��y�W|viZ8u�"z�p'��Uc�
�of��H�RN�*��.L��Qw����P��w��[<�3q
��Ag";l>�5wڅ�}��j�R�cTc�D�2{IrH����x�(`٦�s����t��W'W(FJwv�7����ΟU�,]x�:�"�f-U��\�M��5�0�ȼ�]K{7�D�0�s�N6�b�79S�WN�n�Fe����m�e�˩fF���4N�z�o"հ�M#of��U��-1��3�5�:ؕ\5�֤iY�3�_f��#G��z/�7j-ʹ�gLn��!lyk[�Ǡ�*Ŗ�iVh� w<Ů�ŬX����&�"+e�6�L�7��jD��\��h��8Yq���H�[}�y&m銹�-�u�LXΘ��I��Xl�UI�ŵ����B��^����_�����%��[��	�|n�� �˨�jOw�1�ؙ�N�8�wT��"��kj��Qn��6Y��f4�"r��o��`�2\�O,��ɠϨe��׬�k؞ބ��}�5E����뻋M7\(�G{f�9R3YX��i�k�/��,N��1��g���sy�F��P5�J�Ɓ�C�c˽<=dd>����`kmc�0��I�����UzgX����JQ�/���9pT}|���{͔����'HFb��3���g6�l	(�/V�H�.�W���{�y�G�z��S&�U��*�8h��ene��M�O̍�8 �[5�BS[�Vw*�.N��i���d��1�k��Ie7�θ�u�泳�ua0ō��K���I��낍�2;67,�g�f�pݥ���R�Yc��RI3�jũMj-@|�P�.����C�ә�	�&��C�h��_m�"��8A������n<���\������޲�[��Eլ$���g;(oT�<מ����;�[K��k�� sgT�Ţm�dΕ��QR�zxY�a�����V�Q����[m�������ǯTS��3*�f���Kbqxܑ|d�i�����Y�hcf�~L}f~�w�}�z�m�=e�y�:��)zO}�0	�|�cc2M|����k{
M,��Yq��L���9K4�O��S��4,j��&���h���!����x�Q�=S�xO�z���I���Jm�1���0��ze&�^�MD.�T�k7;!G�G�/<�����Ʀ�EgF[V��5�s{I��
��d��ѱ*K�Z�R-'�f�﵍�un�&�^�Q��]N(P�M���ڔt��@s��7\�奙&>�qz����r��긭9&Ty�_d�E{V��F�~LͲ����ᗨ�c*pd`��֏s�{��~�T
���0ی�X*��͵�����zT�m��2;E'=͞���9*�8S*�i��U�r�W{sĞn�2���F�S�Ϣ;l>�{�6��mkh�R�Bt�&G��(�m�m��:M���Tk�H�C��4�e���7�~{�s���%��9�^w&�a-�e��b�GdP���-�@�&�z�o��c�R,Vh<V4:G�/:�d�����@�2-��wW2��U��ɞ�d�4�cv>�N"����ܠ	j�%]���42��f��-L�=�^y;bi�h=��Q5����sLH���- �R7J�u��|!Z��>�ִ*1�S�4�u{GX��[�vHՓ�\$h_u��zi���ɹs ���n2 �:�lM�@�-?�=��9=�bУ,rE�Oxբ���s��gx��+�Z�S!����5�*��3Smz@�w�_zg�`M��t�x��^�й�M���J�] ��̺��Y��h]����iȰ嬃~���$W7e��A�e^�,��O����άf�F�=�]�odʡ��͗bJ�V��Kq��|ģ2���Q7)��޴S����ғ���j�r��U5O�<,�	gp���E���/������YÓgc��\T��Q��+�;۵t#�3s���5�Yݜ�qlmc�pޭx� �X�#^��/o/ϓp̳��D��z�K���&�-ů[%.b,O�Nr�D޽đ���+���#�s�O1a+�΄f�o�-uo(Ҋ��x�?%-I2*��1iM�+	0�����Z�ۼac�j��v� X�b6T�	&K�.E��ou����,v#�B�ԳMU��7֡u�Bw%Q+�Ά뺛ܳ��ఔ	��X4z�sm9te�es���q�&p���]s��|k_.����Wz��ډ9zQny�u��գ�jQ9,���5Y�У��o'%��CgՈ�GY$>�� ��r74�)�����	�";��s|�d#NP��\hg^.U�DQ#8��[>���iğn��cn7IzA���M�f�c3r����XF8���=�
T�&��
���껁qZ�.������Dq�a8�}������u�T�wŏa=��hzu��*��R��>�������#�T1N��F��EVm�x�d�b��ڌs]�4���a;�=hi���^	��s��:
U`��du5Ս/{b]W�C��v\�"�>�6v|� /\v�ۖ��oY��%��Ko�QiH-%I��&����{���sF�kp�ҩnN��KYe��6��cۑ���v���c��M$Czm��z��Z���Z�G[Ou�#����4-���*l�	|)hۧl��1���C�D;^�w��Iٱ�ct-�U�u���P�s�k�EeOO��Et��\�4�s[���Ƌ�ܳN��H�̲��q���GH����WmgY5�m�%�f�,�<sE!��u�U�������s!H�D��3a���G�-�m��1��0S��K�J�T�u�!YZ$�՜��l�H[/���*���yKavI�Nt�jb�+�Z������r�xf�����Zc�'��wI{8����P��mN>�--�;κ\=�ki��UyP��.��X������乜��َc�+%�rP�Fo5͹�;t�7��*�c<m�-yW�[�;������7��+u#kv:��me������.��Z�܆ٱ��+�Ȉ��yT0J�[y�͊g����G�j[k��7��:�YI��cE�W�f`�:��MP��c��\fA�$*�W�]rh9?�_ׯ��Q���S�)Z�UP��6$��g��!$���E�Y	$�V����L�8�"�ݝ����P�eY��pd�d�͖�6S],Q"DR�H�VY		 �B@�	#?�3���F�Lg)��h��Z����n�=ƨ��T�9j�iF"�[m��/D$�<T�[�J&���-y��i�F�r.hm5�5���ra��%�$��,jd����)C��&p�Х's|[�~<(m�4Ɠ#M��$荟����d�o���h��$Щ4"I ~P鈪�Iwtt��˚7,t�쟞d�#煟�뚿�����9���xU�������#�o�Σ�IJPۉ4=��t��k�L��%�f�t�+Z=�0�$[��(����IF:99���(���z�.z3)����I�abH�ᅦ�I�w�إ�ٖjS) 	�Q$I���I�����ׄ����4�Z��s|�h�Y�~���7=1	$�g#5J��,����c��-���|�Z��_O}������r��cjtO��X{�o�,�}�֞�?����R�$�1�������󑽛��;�Ç���}T�g�˦�ZE���-���ϫ��XN2`�q�p�=������~Gw��4t<I p�������J(����&����S�=Gf�YR֑��AE.z"Hq�'�E5���D�J�#��-orXݒM^e51$o`<ћ}ȒH���Ҋ���`���,���Ro�Z-&�	���N�902��ٕl�Fw�Z��Z"l̔��3�Zz�IzKY�d�.U|�d}��H%�C���mH��BI�+�ޓ��Q�xp�I�}���76qnGޛ(��⋒9�Rned���J.�.�u�;��u���_�:$e����/��X��S�㎇��֋Yd?R5EzHI ZOn���.�Ϝ>cY��}'?n���ӈ�oG��M��1�F�T�S��̕)E�z��ޡ�/Xs���Ff�r6(�}�U[��W�[aō�w��!$�~��t�8˺4�銹�ݹ�Q�OV���k7�'�Q�Qe�iٝ�jaAcژH��J�I �'���\���U�<|�f��wD�t�N����F�8��fc�,�T�cK��M�r7�T�GtS�Y#���M�f����"�(H\U��