BZh91AY&SY�w�  �iߔpyc����������  `�����Q     � B�� �%@�A@  QE;�� @��  aG��J�J�}^�Ksf��l�2����m��AW���8��f���Jv�a�N�q� "��;��2�%��1�hh�a��S�_z=(8�uB�Jy���fT��}4� ^-Q�ϳR�J1�D�(�[M�!.��oq�[M�K��x >�!��}_]�6}�q5����::��\��*��MQ���u����� � ����Z)p�l�ѥ��l���p��,��(���UR�� �i6P TQT@I������ ��T�&R�RF�=	�   4�ё�OЈ���d� ��h �d0�d�Di�d� �   	4���T@� L4` bb0"DT�T�L�dm#C���   TR)�z��� �"�Pi�j����G���j����.�'�R��	�����W��d�!�I<�Al���I$4�!�����Ҷ�7~K���0� ��I ����V��4$��U@�:1Ga�I%��m�~b�'V��z���c���}���/�ÿ�w�O���%B|6;��=q����5٣�]���Ä޶�������ُT��5f�	f��v�2"я��\vȘ�}�e�z ^�t�l���h�6�6��m���pc5�z�c���D8!��xݐ�r��[�11�" " !�J�d�F"�?a�}��zv!��oݣ�0־b���>��g��k�~o�|:sS 7r���N��Y�
n�F7����o얝
�K���X����[k~dF6ڶն�5P�W��
�V#"�8$3Q�<n����w~��w��{��������B-7{��q�]�0���6�q�}�!�����7�Z?�3>&|��>o�<޶޶�Dϩ���}�o�w���<�/���~�^��>�x���pC��d1\9l�p��vŭj���8��S�Nn�pQ��ȗ�CmS-�������nHq��!�òzY���ψ�����
��4[E8���#]��g�uo�-�����m��M�=��6�`�yc���1ݿ7v�����Z����c-�y�6k�rvߛ�ڦ���d9��V8��3�8��ݘ�צ8-�llo\F7L�HȌ��ڍ~��)�(�E8�e��xp�!���o""=Q81ɮ�0m�e�c�fd@dF�n��n2k�|���e�dB6#�h"�Co[P�Ë���`�b���.l0�Hp69�����7{Ì���@D@C�lXٍ2�t6�y:�uW.cf8��\h3tp���F�fθ�O"�ڼ���nQl�Ƹ)�:���U���1�B"�\
Ȉ��<␮X��!M1z�#�$�����47l^���G+<����p-2 -�"��"K�B��?y؁@�O��v��蘏�[M�c�J
�q�jъ�����m�F�[�7�cL�ݡU��qH�� q���D!��.!T��Dx�����jb<�
�",���،�Rߑ�����=qc���R����x��G��Z��(��"�Z\@c�VlE��W�E����{U��)�k��[�|4��bxӋm��NPةR>��)K���F2)�"�{??y4z"�Z׾��P8��M��>b�b*���`��H�g�P6�5���=Ay=Ob�o�*��=��+��RS��䢒�+1�cx��^Zߖ�+�ӑ4*�W�	�Xݫ��b���,U�@��i��M�)9Q^hHX�CM�6��ks*$LY#ybt�)�%8X�}�Ƙ�H�@�+�׆أ愽��K^KD�G�؅J5RX��`��Bb��J��)bb�	�(N=i�����[H@��W��ؘ�^E�G��Q�B�O�R<�M_º� ߧ��殕Ҋ�,�6�s�տ-k�D��F}�|�(ޯ��p��q����z=��1����.�יs6W�uη(���ݎ/��<�""�;3b</D֋w�Y#yJ�o0���Ng���瓌P�e�n~�QBy��ϳ�Y���Z!��ϯ�m���*�����[b`�Th�խƞx^���D(߳��3�P+����l�V6R�Zϲ�wJ�7HT[z"1������Ս��Z6��۽Fy��L�_ԭ���څPۚ���Ư�cZ)h��\�P۪u.f�"h��K�6��i���fDB57��5�k�`�",v7��NL�d|����-�q����F)� ��������lU�L�q��dz � �[��Dk����nKq��z�����q1"��+Y��!��Ǫ�y�6S�����v�o^jk�ݱ\/Sx�,hZ�?��6�d?\8�r�f;�l�[n�舉�����&�a��}���_�~1�������m��ۀpC�麨p�h�0�`�P�,ۻuOKp[�AIܷ��7N[t�e�y�����n�&��1�\����<��cwn/K��7�t |
FԹz�@'�Mʉ����\N�vc��̕��(����C1pxh���4G=g���[�4M�oٙ"z'�M��d��E�)��C�����W��ff�L�y_��겋M�2�b׷���&��۵���#�t�ٽ[F? �ș�=���2	��t&���߳�
{Jk��sv7:㴩��At[ŉ���ߔ�s���d���G�z�}\��{���,N�ִY����=�'g��>О������{}>�t��jmn�˻=�cƳ�Z��vv-�������o'޽���]��Y:���ú��sw4�鵸�)f���ώ�f��1n��"v�e+�W����M_�~�1�컯e��[ gc���w��|fc��v]������0���T��潈���͞�򨙤R[ӟG��3Gf��O�w�=ݪ����O������S-�������^��K,��My2"��+Y2z��|�JɯtS��){_~}��s�b����w1mM䜇9-çpd�Y�뙿d(�JtɣU��4�{���}8f��g{&����s�e�n�=����|{95���.��l��c:��}M��@������/��%�����~�l��)}2�'ƨ{sp�Tm�l���ë	w���EzbT�{���s
˦?L�G�u�����3�{<�_L�/�"�|�l���f���E���L�#�O���q����Z�������̧g�:6����:�IG�sn���g�$>)�5���;g����e7�_n}����������H}r{�b�Soǯ�ݲ�am��>*�v_b��V�&���or��Yh� �d�|	������S˳u�xe�`eOj�G�ܪ2e�1~w�~�VdW���fj��b�^��ȯr�OY�g�Җ�yI�:�h}��ku��ə,�O������f�3��ڲ��G�gw��I��Wט��˹���쓠5٠`��4�{$�/8��]j��r��Y.貔,T��:�_�|}���8���)���3������^��p�ӬٲW���n�7��ng{����O���:�͔�+;{S���Ŧz2&��b�BtR�G��������Ӧ��[
����>��7o�rߪfo+�:~��;�����FL��yn�O׳b���ެ�c��z�ގ��{4ѝ����ʵb<%���I�酛=����dk��Nf�^]}P���<S��) ��i܉nY�0EȂ?�4���iF{��4����Й-����R��:a�0Nʷ^˶�3�d�s]F�l��SO���a�O4g�FB�E�w�۞��$^>����ï$#����6���̳�~�Eu���u?N�fJx��=5k~��x��|���2���c��==�}s|Q`n��s%3vbs��ƴF����n�=�Ξ�����V5^�I:mɆ��t>w~�(oI�񤾐���f�����=�@����۳�\���Bm7ϳ���S�c��?vN���]�7�̳O���cd�`K`G���W��{2X�gg�[0f�ޞ�ֈl�N�����|����w&aO`�}����1��M;�2���_9�:�������U�=���re$�4�3�9��:��V�����s>7���T]j�C��x��g^�jn��b;(�_��N��a��~��}���i�(�tTs/4y��������l�w̪w�=~ǻt�ϏO��2�%{=��׮e�'��G:�;�,+���3��4�����ke���^~i��g�~�Ԡz��kL6M����s&ک����l]�Pz�v��s��N���!�����A�}����V��-�;�����+�'O[���l����fjl-x<~�zrI{[q�VT��5���6��p�&!����e
j6��5Z��l���L��aE��3f�c@��Z�^��nY�"�ǭ_ظ�z������A�Rm\��蹾}�R�ֽ������=8������K����;=�v��.wm;٫���N�vG�.������es`��fM�Ǐ�c�;��z5�L���9�ʐ��;�)�z�*o�'��Sm��g���t����n"|fͭ��~v��-J��-�+w���������E��'0��;Jڥ�"Ʈ�ۑ��28��ӈ��Xj3����Q�$����� ��4�P�bR֐�!��ز4��q �
G������U���.d��u	@a��A��J�"qPN�{��i�u(rT��6������q��9���n�*p����H�Mi"#%PB�փ��+�eJG ���D8�Ӯ��	lw�w���w���񺨆q�%~��Y��Zj�P#��D�[ݐJGjaqb�
�a-8:&C�K��;ˍW ?�b��SS���a�9~��jF�����ƅ@Ğ>\l�7�3En�8̶&�_�'��k�PkBGs�+r7"��+�(Z��0H,R�뫜��"5�$JX�Ԛݨ�M$���d��� kM���!�(Ci��&�c�R����~���ن^E���oʭ�#jH��L��+�¬i�W1�����q��9R		Br�9Z�O��QQ�ʪ�$E"� Q�yK	h�}YED��b���I�Z����Eg�9�'2*�EJ�;�>��Q�(ٵ� X:����
UlDo��[#x�"��n�Q|c������C�ر~����^�=�!}f=���6�$BDg[�ʭyy����.����Oq����#������+?J_��������O�������U3% H��� h�  @  0 B <  ��R       �;����:�"�
� �.�w��u���<U2�	 (�`@   �  �	 (A33!� �`  D  `%��}�  4`�UR `x ��<   k  5�x ,@@ ���$ � �  `0  ���}��r%��}�����	S3     ��  x ,@  P� �ɟL�P� H��� 0 ƥ�4�KZI7��}�o�!�� &f&@     �< HB $ �  H0 4""f$  �� P� P j�� S3� ,     �� , (D ��  XL̩  ��h� �<  �s�:�E[d�J�ط���O�	$��mG�����������I����^�0��8=OW��������9v�a�[�˖L�e�l�t��ɓ�&YV�R�HB�*B�kV!T�j�
�^Yp��,0�edɓ&YWf[2�,�;9;;;;a]�vdɓ&\�&Yn�.V]2˶\�l��G���ޛ�r�d�m˼ͺ��J�B�M(�_�W?�����a��������*��!�Vj�pk�4��nƘ���@���L�;hr�Q���u�����ao�NFˈ��V�mW��^5h�T�e�����L�TDj���L�Ck3�I�n�qLQ	.�l%,�uY�5�N�I�vFI-lj�J`�#�J�2s�m�02�!��up��XX�$Y!���-��W
ψY ��Y�0%���#c����.��4J�ڥ�Q�AJ��\���d��&2���	��|�F҅Y.0ΓI��o2Kl>��SMF2��N�!k��RX�)��h,�gi����u��v&�^��"�+Z*	:��ԭ��7�m�~��U�f|��s��mN-�Ҫ����H��u�h���pa)�nI+d�YU�\�T�-99)y
�r�ӵ��W�t�JmCj�N�s�Ƙ�X!0���))c�3M���S,�D,0�&�8�L@h�k��r�cv�r�*�hc!T����Y�@�Vؖ	6а�!=bS�$Xڶ�B��2U�C��䮙)dBM�PEv�(�8��*m
W]R�:���)���_8_DS�ߡ�>_(�]�8w4|"�{>ֵ�{��;���(>ϵ�g�|�$�_%��wS�s@�K�뻺���x����W�ֵ���理���":W&N
pN���w��-�3Y�6ԑʩ�l�-+q�^dA)-�1��V�q���bK-�ju�BERS�q��T8 ��78��Ui[U�񰅕^1"��J%�8�sh�	u4��9�kdd��m���U),nZ��l���p�����K�����Hk#��#&F%�����x�'�t�E�<��� �K����2����20��9��6h(S�l���fW�s7�I���5�;q����.]�e��m5IO�7/v��d�!��<>�q.S�K-U��TT2头��qk�����Ɠ�/�M���(SBp��c6ϲ�}K�-��{tx�d����,�3�������p�������7���UU���#��|�����H���Ҝ5�$a�	��!aAF�l�fCf���edSd�}�U�d���R8��E󔶧dV�uZ�1E\���3�I�)���N�jv�:�w|�gc߮*�0�{8&���9�a�aȔ(S���Źks=��[�u����̹����4�q��:�&*#mc�	��s��Q�
(�P��%���@ZI$��*KS���ż�^�^@��P���֜�@�g�-��Ji�OSZ�*�B��g����2X;�U7�4)�><0�lNp���}���I�A��+mZ��M�HM�Ci|m�h�������u�F���}C�dۙͅ
��2�m�����!bs�ѩ,;]�{9>d>�Mvz&4'���ٶ��+V��%5!�"��X�Cq�[�t��[��a8�Bd�[v���D����j�^�m3����>0�bRq�a5�%�6�f��QTm1���]&M�x���N�ن�g�^�T��|0{�̟O�<�q%^��������ٓ6�>�y�P��!g�y:}55=�E���S�E�Ro͟
Q0���,Nl�ͫ�����7�.eu9�f��:�v���u���H>r�W%P��j(�,�*htB���ˆA0O$��������驚s#�����ѽ3�,;5����|�\�r�J��Kf9ߨ���}m2Y���7?Lh�8�ō>֜d��ӹd�k���Ʉ�;"�g$�QD<Q�e��h�B��� ��"g�ٸnr����_q|��Z�U�#qI!"���ԩUi�t�qt�N�0�oR��G���/N�azZ��Er�{Z�hi
'�D��G�#���Ylƕ��xV��X�a���:3���&�Kݍ�v+�G��FtM/G�ø�8^��K��K��z=:zg�t�}7^W����t=\)���z(���zS�:R�M�?�
=U�'�Q2�M���U���tV�j���DG��/F���c�i�Vc�Ҵ����<Dݜ덼g�ƿ{'Սz���#fF'������M�Q�����{��-�~��}���bƏ'�7����3�]XёZ2���׾�����g����G�U������Ȉ����}��Ww������K���ϻ��u��Wqϟwwue���w!�wR�]��wrwuw_��ﻹ���Je�0L)��:a��ph��(��X�1�d�-�R#�+ƒ�?"e�I=��1�#�&�3�+#�PC�1Wg�����b�Uw�ݐ� i��6�<���.�����r*}��A��|C󔿜!ȼH� EŤ�q;g��<L&j��)����$:��(��,�x�Q�d��RK�9�f�lu���p��70���Di�b�¢USwW�{2�3�	h_�Nʄ�eh-�o큔����0m:�>J1jRV��|o9w�q�a�$�_��Დř�N�K!e����a����y�h����.����@�Tw�@ʫ��QC �>X���%�X�n���)c� @�$1T3M��X@�ǭ�x�sQ��Hj�[T5d���!�rW���k�����Jl�o���8���z)����3�n,v�Oa۠�<���P�������\�L�_'%��u�JTF�O<���?$w�C��U�T�և��D����iE��h�(��sV���!u�����6�*�����	�	 ���Wo�֩hI*,�8�,��;(��~��a`����vk���m�Z6�C�=:{�ȁ�w^�)�x!Ͻ�C�NL)�M��l8?hH|�JǴ�ӈ��$$W�Kh�ǁO-6���=�$��&��;w+�Fb�NG[����`y����\�f1R����i̺,	��9!a��C@t˷��>,
KJdx�
���㚖5:�#�����t×M���
��$��Q������(��'�*��}m1�rz`
7d'e]U�R�۩S��5VT��8N!���<��#I���S;�8:~!	!n��u,���)��8�L'\X�m�zƀ�T���>^��4p4S
Sf?l8)�oJf�������5%���^N�y͍m̸�*%vDH�`��TU�*��31A<���F�@��E���c�uV��2y4�]�:%� n:�a@�2}9�s�Q\ �|��m6�h;��]�C��� ���﷌_q�]�94���7�rn�9����fZs
����ǸU�]�ӝ�0�%)�,�}(�YL��?0�p8k�S�m����v,.�'��a|�8~�!���':���ZZW�%����54~���f�vC��(�l�
Ѯ�8Ni2�h	P2�'S.�$��3�6��Ġ%S���O�E'R�0�%lن6e�s��2qa�|P���J�dٚ�a}�?C����+�0�F[~�^;��#`N�σo�"rԚ���h"c�E)�Kb���BA����J��Գ�0[I��l �������
i�G���A�f��T��x�;8XB�(��Μ,�h4e���J�=��}���v��8p� �l�ˋkY��Z]�-Y��n�� {��۝�a/)�nB�^ �)�+�6}'�'�4��%L�UE|�	��9�6znh+@F5�FD�e���/f_����x(�?8(�(�!ѧ�|(χ�N�G�'Jb�^��t���i�.XiZe�m+*���E>/E��
�*=�:]/�qzx^�����Sލ��=�����Oו�L����z8'L-���G���Ҝ3����z<��'j�щ�QƉ�D���tQ6?�Z?�G����җ�t�N����z'L/D�������x~>�Z[k������y��]�痵�Z�8�C��#������p�1T�mN����ݓZ�����%���<�����t]��?�ǅ�9���*����i��D���^�c�z��/(���RS3=���VX��Fbr♺��]�p�y�d1�����=����F,��[y]]���`���Grs�B�]�+Tk�}�~;�ޫj%<�>�A�	��}~˽ק�QK��Q���o����Ny~�֛��_r�v=��Ey�������C���b7�ȼ��`�&����ƅ�\*�UUm���4�@�|MBv�y��U���o�UO���F�ň�V��IJ�
Ь�U�Gb�b��QmM�J�U��[��P�/�$�=F]�w��C������>���˻���C������>�����寻���.��������I5��
(�~QT�-[=�#xی�L�T0K�	�Ű�Q��f��'+C8A	ƪ�Ո��!ګTGV��v7K.�4�l9(����ե��҉����I�ae����Z �#R�1z�e��m{�ñ���@��[�EM��K�b0X��AJ�RQ�7K�D&,"�7�:�[m�-��Oa�@,~:"�~]"f�)"X�u5}t��?�i�/TEPK6{J�M���b5F�u�{W��袬��y��7%ݭʺl���G1�
�i<p����Ѕ�QF�6x����ꪃ�W��=.�р@u���5��X�+�1�%`�3�5!�� Y�,>�V���6��V$�ˀS��J�F��NCp�vG�L)�|�p፦�`<Ln�j�GхrV͘a�f^7	�Z��R���*J��,Ɉ	ď�mӇ���-���t���v�%U�3�����ĭfa�k[�v!�����`}�!� k� Q�SHag�����<uJO���0��5%t����w���Q��%pن6i�s�����P%�R��r0��0����c�7�^�vܻ���d�HIi�b�4��(D��`c<-J�3	$��ߌ����eoG�@"q��� e*�e��'�@g���l�����J&�������jZ���y�/�K}1\	������C]9�7[�q�L8��1�s4���b���Z	G@QB�l���`���qeU7[y
�!�ڥV2;$j����R�5�����0��/:�nx�d�)F:v�Q	9��H�II�ahe�ڇ�v�b�!�0'�'���<���Hjzv=�G�Zթj�G��x�;L�0=B9m<�p�铡
0Q�>6Y��h��o:O`�F���3Uw'��g����v���`�M����m�t�Hi �y?~���+d��K2�e��$�� ô��š�}�:��WR�\�d˘<�c������d����'�Q�:h��у3&D.4q���CF�>�-�t�ʪ�������Ick���Dq�VF�v3��(mB��F��&~�z�2�H|׈JH�� Δ7b�=�Fy#��%��&0�,��f�ß�-�MLj�6d?B�"O�,��O��J�J����e�l���[JD��o�8���D�Ґ���ƪ�Q]r�2?i�ht�>8:�|n��9t|e!��
&��4P�G�c�����7+
�Zh?U<�A�;\UEA�gm��6�"�eBd��O	`e	TnE�y�n8\Ŋ��Pc�x�ʜj��li��W����ֆ�e�a
v��}�,x�i�ZRޥ>�|���2��RcqJ��P����6p��R��!���}jI�)M6���țs����r�˲̥�8���V�~>���M
�!E��UKR��<��8ԐH�O���o[C�N;2�=�f�#%����!�$��'N�c�Ku����M���X�⭱���X�@�)��S��D;�F���KI>hz��S�4|a�d4{U�?6t��(�3�l~O���z4z"t��)������W/<+�l4�.Za�,:V��G��Vt�
%zUzYѝ6]/N��zgG����x^���=�����|�ӕ�S���pN��=���G�KM����gOǆ|8=z":��D����Q:(�����c��?�O�c�x]���^¹]0ƕ�h(�աG&��o㻜�C������n�v哗$�k�.�R�'ê9�u�O����2�f��n�y3Q3[沱�������͐��J��o��M븽��+r���E��_�w����_wwuV]��w-}���Yww�ܵ�wwUe��wr���]�sww�ܵ�wwUV]�wr����RjT�5�K��Eɺ��v�2K\������ҟ|���g��|�s�I:UT�0U2�S"�ʶڔ�~�𚜉f���	�a��i�O��Aₐ�|�5�d�
���<�0��xzh�p8o�6��>��Zd2�H:9	���Jv�ڸb��uT�b�V���D�C�B���I#��y�)�v޹r�C|J/�!�'9�'u�����HKR�'�ɇ��F�t��ɒ�:l�a�я{��c����*�ֈ�e�խeM؞ሹ}���_/"U�ܰQG���	�9$j��8����WN���z�C@z㄁$d��ɔ�41�N�R�.r��sq������~���~}#;-&�:t��&T�r��)��SJP,J!6u�S��.�K���k�*�a�|��.`�	M<}�a����e>0Xh4a33��M���JD�6�t��[� �)�6�pD:E4�X�4qʚ���TĢ�e12p�ܪ��"�}��,���bl�i�&�%���x�;<h!D0ه��p�s�0}n1�6���F�m�'��0�,m����n�f?Z�*��y���ҹ;�np�=-kU�fyMÒ�Y�.�t��z=�d̀i)�%��N\�<�۳�
!��x���������}��sz} j���p�H3�ClOuy����������Ë�Գ�_�E][Ww4�Nm�n�𪪕*��L�DM���M'*�Gλ�m$�����a��JCGo��қB�.]�rݳ�)��:ޯ��:���"e��4�Œ�
�mNVI�LRlx��F+ ����C<���-�ņ��p�U<�f
c���I\���(հ�Ay��\��B��t.ː��A���'�i�"o�2�L��I�T)4I!1�$b|�\$6G)̥L�˷)I����?'R�������闐,����$�kDM�n�p�P�?K;b��U�aZr��)����f�n���]���(�@|��0a��4),|���J	�'L���9sqNN�P�5��/�]��mɓ--�E�C�P���p�r�����>���Y�pH�/Q��NQ?~)��?Y�G�kUZ �U��F�0i,#��m4&D���f��ϋ�IҊ��Օ0�K�M)��h�P�?L��Y�2�\�h)�&��-�>��B� �N%�:3����vu�7}3�O��~)��p8w��0+��nb�����.��ζI�b�t�<h��PQP�x��|����&��fO:8HvL%��8O'5�\pz�;�d�>�p��+��ȇ%'�3�C���x8{U"��/�Gោ��(ρ>>�~-zQ;T�Kџ�C�����ۖ&���L2��K��.����*4EzUzYѝ:^�/�k�'�Tr�/y>B�m��b�|�G�k9WA��z8'qm��N��z?.^�G�џ�N�WҪ�eV�U���VX�r�^��-{\-���t�6'GC���OǵS�O�~;_�>��{�� �E����&�V�~.d�mƤ��c��h�����4+0v�ɚNA�&[����93ɽ�+1D�BV�=n's�ߖ��6�ަN�l���|�}y�]3"2�%��oo{c}p:̷�/�;ݗf4c}��[�vd�V�w7��w;9�i�x~L�gw�'�����-䉐6]�tdr.ˋg&ڼX��Q�1�������Yۉ�M�����{ �֖��b1�ՑHUs���+�&����氛
�I<XS[[��Vv&�7!�� pEEM4�+��5����7��G��P��,��'#����~��Y�҃g]̸��3��ٜ|�j��&*�b�����ǯ.]�;Ӝ]�wc]���U�w�ݍwwwUV]�wv5���UYw}���wwuUe��wc]���U�w�ݍwwB򔚄ԨR�rk�J�N�x/�����a!]`�퐐Uyڨh�-��Sf3� �WQR6����k!H�%��b"b�)f��B7��`p�n7Jq0V8�,�UZXT�$�'�e�+*j�eb��*�!
�E���B! p�[��AԾ�r|��	!��u����-�=�a��H�	��e���B�#���#�����|���w����^�5��9����W1�0�3�;�a��a�be�%a]0�õNN^*�+ Y$���M8o��UF��%�S/��M��!��y��ܐ�"���C��x�v��ϡ��(/#�9/�?C(��$x��I�Q?���'����\mx�(��8M4�V�>?M��0�0��AjG�\�*�Q�t��<��-dL$��8�T��p������i�%S��RF|�>!���G��Na�tB����t�(�������O���`�a��d��NtQ>�h�I���h�����e���0�نf�1[@���)�T�B|�u,)���f���x�F���Q�̒H|�4���>։��Z{�B^k�D��|Q(���.jZ�_����~�xV2�,9U�1ۍ�[P�̖�!��T���,��aR�j�\�8�Y̙1�r�c�cX��e�\Xa<�|��lX����Ī#��FR���1	>p��Q���i��RUW�Avs��al��ˀ�檥�C�����S!�p�n̔�x����4��h�(�٠4b����t\�����fHQW�Dt���FX��[>r���O�I���Y?'CX��r�U-�[�s%/�EZ�3p�DU��;=��UN�L}���/�rI%�2(��:p�;e�@лHZi�����I��i���~!���B�nU�Y��Mގw���aTUa�MbF��FYԂg�%m�w��q>ѣ��g�&���F�A�'��J2/'��$l�M<�ç۱E��%��O~5�Gǁ����[i��I�r�v����I�N�K�vx:�xa8e��)��Z|p:Q�d��>!���ܪ�&���k��+yKL��
��ZY��W��\z"C^Q5L�3����S˜l�nKb�7k�0��)S�XR�����u#���\�XQK�!��UT�h�a������H���Poͮ�ɧ����)��J̸5S�~E��:ܝj"��].~�V��?/$�A��=:�w±C�b����c&(,��r�r�n�a��RG�GL�� nS�S����=�ý�-���L�adתrնZ�s薫Z?s>�;��3�/�bv��%��@ӽ���<��i2�|�;�S��)����G�G�D�Q��C��̕�U���.*��ᇅn���yxa�{�p��.t�e\������������Ό�����z>��:z]�ץN��>��K��������zZh�qiN���G���Jt���z'VxU\��aW+���-VV�UYaU���^���F4��S�.�tt=���:>,���~:��O$�
~�L�|j�8=�v[ib{��=�˅�i�&����zMf�	�2<��.���b�/���+s�c���ſ}WU��}����)l}�����G�����d�y�[]���UYw��mwwwUUe�wu����UU�}���wwuUV]�ur��˾�Zֵ���+v��rr��Xż��~(?�`u?���t��J��u��迤��GP�vUg� HqjC�'g��캻$Hs��C�BO���]�I`��vWU���D���6xne�tæ\�N[��sU$C"��K�d�Ue"E�m'�Ҏ214Ɔ!�q�?z[�ڢ{��汍J35F�e���KM�8�E�P÷�S	����8�*�d�;;t�h�/�L�6(�
8t�KR��Oڿ��y��7�I�U�!QSG$�ט�we#U��[B�#����
ӕK-���%k��o3ԕ�ULQ@��jn��/$Ut��R��u6�a�4�`X�R|좞v��D�;	$,�����(�v��O���R�tC��Q#!�QR���wmє�s��dɖ�l|��l���p�.܎N[1c�FimDr��&���v:��V�������3����D���l����ˣ,N|*�����7��p,)'���k�9UY%iХ�����K��=���5j�S��N�{D%N&�d]�f��GNA���Θ�3Y��0�CX$�M&	��a��Q+R�E:sG���cdm8ku�#����X/�R����I�R�J���v�L�	��UO��=�tc4m�G�ü��l��0p�5�z�B˖{a�I3�Zd<&�Jd�kB���S|�qo9�+�)#`��r��G��v�
H�;y),�"�Hq��0��E�x�a>J6e(�nUJ
��zb��+���G��A�D�3z�~�)�����N���*2͜�*��V���9N
ʬ�v�Lu�
󹒼��Gd䊎4ڂrQ�<��J�0M�����-��n
�kTcR�X3�N�Ֆ�.N`�����d���m&�g��>d_�]&�<��R��OKԆ���p�	��hZ����[PiE6dL��F8q�-(��l�46/#�=H\
�+B��i�ƍ+����	!�۳�ܔBI	�dti�tu0�S��	��9g'g��Ѿ�M��C�L�|�ӌ���K�A@�r��?MC��8i��n&��<m[ZSP�h)��)��c�Ѽ�͋�|����k���	�7)�&������B�M�蕄�����y����[�4�!��ن�1>��y0��B�r�a8t��>:ht���h�]�VZ`Z{���V/�!S��s�EX|���s�O�<a+S�4�34SWXK�Z2�����_���i�?dp�Ѵ�́�������͙�1��\H�r�����;��i�QE��/���[|1��Y+J�ZU\��ħ���8~)�t��~g�����3�ӵ~������Q��Q�i�'D�t�6^������������G&���
1j�O��iz].���(�A���~ѧG��e���#���T~�E�D�Q�Q�Dg�O«��}=0�L.	�4=���:>)ѝ4_���O
�s�������պ���nͱ�r��%�Cz�������oM�O�c�O��?�%@��Wuh��:79Cu�,v�娹.&��3�ȿ�}&�骪ؼq�͖mOQ�+�f_Wk��X���PC�+�w�o��4�T�Vd"u�5��y�i���!�ͅ�f������jZ��c�ry���պ��S$@�4T啧+�5"�٠n=�{o+�[#~̈n������p^�w1����V"b�{V��Ec�9Y��D��Ow��W�����׺jd�tUu�:�dq�e����4%e- n��E��C��X���Dl���o"���BT�PC�ZB�o���+|�-k$����WP����dSșDI�5W�<����~���e�������ꪲ��{�ww]UV_wOs�������]UN_wOs�������JT��B��jZ�!j��bꔠ�%@�n�R�r��(G93��׺�O-���UcN�9d��
�
�#�	�%���q�a�|Q;[�Hմ���]C�1�T�6��%�R�Bƣv�>0	-r!Ș�+�[�j�(�9$�Y!h:�J�X��I��C�󫜜fcm��0M����MI	&Z��|��V���[ż��H]U.��}��0Obd�j̩M"�x<0c����7�2��ߥ���jKs�٭I�~_(��\(���qD5��T�����M�D���`�˽Z�Sd��7g܆@4}O`��T��٦�L�XMKG)��ޤ�?/���$9�z�S԰��������e\�kSP��Xa�}΅/^�N&,3�#��0��i�-99UW-�^I*J���Y���J4��S����|B_���U躟�-��k*©T�e�K\Ó��)�0؟��k|>���NR�D�҃i�2.�KJㄴې�(�A����j����̨�Cf����aO6δc[mm�m[j�����2���4��j��-����$v�j��㔪*&p�N�\�|Pa+�8�v����I$<���4:Ji���l2�4(Z�ZV�V���z^�{�Ε?{֖ڭ������$����͘�$���i�$�Kh����8\���v�Ɠ���p$Ô�g���Eu����Q�,x\�N�C�xCT��>6�P���㬤��xt۸�+2J��񭶨�p����=4)������Jj	���<)����'&�|ɂ���[F��'l�}��0�x�xO*d�R�V�6��筆[h�I$>t!�IǍ�M��jCtv�a�v���`�M�;Ę��v�s'H���6b�>�v��>?&���ۭ-8Ia�F��M&K�ɔ�y]�J%I!$�o����tuШ��!'��ʦ,��YLz�v�5�$�&"}��ܓ�ɣM�6O8!�kWV��s+^!��f��L��?p�^Xd��L����+��1)��>׍�̙\�q�;�6�?qyg;ȿs��kܪ7 4�r�\�z�]$9gHe �lM6V��Q*��O��{���UD��.��ujZ��W��?����dNH��0����l��HB?�z0���Ej�Y�	E�Q��B���[Nș#m�
��S���܁c�4��&��==l:�6a�9�[�aM��|�B�nb��D�p��Ü,a�I	]H�)�7��=�V��9r�O}�u2u�6�Fm��c�A��0Q�f�A�c$%�����8t�8ģe�o�X�[	�UC.x�v���|p�Bq��Y�Bp�5����R}�Q���i��By�)�I!	f��t�\�89r�n�̲d��۵i�M8iƗM4Ӷ]8e��dɕVYa�Yn�-�p�.Y,B�j-B�-X�R/!y
�2dɓ&]2�,�ˆ�Ύ�ӳ���F��:e�V[2�vYr&!h��K��d�~�^�WU
��U�.���ꨄ�ȱXIq_�AE��'��Mχ��V��&�˒��kXU��x��������E�eUN�\��hbd�d{��J~T�	��5_ވ��ԭُD�����U���Os�������S37��=��U37��=��U37��=��U3=�����T��
�d�'���1P��G.C���"R}���9i�S6���3��U���~z�3��'R�&p��S}��9g0)�)����˾�Z�8Ŵ���NO�s��m�����@�1�/�t���c�O�--���8��1�95~.���Zѷ�y7��\�r�d�u��g�0�9��I�v@�SBxSgN�h���=ˡ����ݶ	IҎe���{ �raͮ"�GG0^K�+X��!�6(H���B1�$�UTn[d����c��6X�l&�]�R�C�ZS�Ñ��3~/�p����!2�dӳ;�А�S�	��	�ro7*�B^d�l���G�ޕ�=�.�U7��h)��)�Á�}��b�����n <����ʽ'm޸�hk^ܜ!��Gji���'��>׷p�n�h�A[M�6��%����J~� Q$�u7�޺�&{N^u�����6Q�F�A��$¾�$&�	��f����d�g6��a�BvO��fL�6�[\�mm,�C����n�n��L��|C��ª�����?9�I�����.�
4Ce:p8ͥ���o�ͭ�B΁���O6���$		IQ-�N�ˤ��He-�I�� t�z�EH�M�ǚN�:r��&���m��:�t������իRԿfO���89��I+j�*,cM���>WPZࠣ�Ԧ2�[��c�D")9Td1�I�ù�t!̆s&�S�Ξ84�A-u�����R\L�q�W$��v��a�p18�0�F}�|�f5�:nrp��i8l�ð��_=L&�fV�r�.�,��&��	׍��dIe�����N�C��:�&���0����'�=o	��e�&]�5��>m�w{�̟]_H�r�k(�� |��CM���g�D����:lO
l��p9�G�r(i1�s#m�M��0d�NS�H4��󣒊���|m>�ͦ΂aӬ`�ɬ�]��ݒ���Ii�Z{���Q����֜'���ۧ��m������4Qӆ�A���Ƣqե�㥖b}3e���X��z��ө@& ٙ�8t�ît�hi�0��I��q����� ӗɳ\�\�i�y���eX�;�a˵nh����*����&L�;V�iۆ�r�N�a�m:r�ed�ْ�ʶe���*B�K��Z��Z�V/*B��[2²e²dɗ��,�ӕvtvn�����4dɗl��*�6/!X�!U+�
����"s0���p�s�����޽X�i��x&�U�t�r�3{ޘ�{O��}o��N�71>�����}ƽ�Y�R�����:���o�w�:G�R�f\U�l�k�/�fI�Ti߾j�5S���p��7�y�m��uUE\mk���ٛ2, ��}��[��f�W��pi�ds����ɽd��mG���}�L^�RK+*��j��>&s0C-���eǻ���]F�-�oTZ	�#�&�V��zC^�ˬ�ˑ������~�d�.�V(?�U�ˍMMv'�tN���J��aTuYibm
�>JI#q�H{��X���mDqQ�H�ef5>7+���2RyV+yf�Y�96���Yo��F�����qE*�˙�8�9��7�?]WN����������wGwUL�gw{�����g������ꪙ���ww{���{;�����T���I�P�r��/�o���!6�nVr�� jAG]R�X�Pu��MWB֚�sI$*�Nu��ⷖ3#���C%`%T�P�'! +dU�6��,w��)f9+ɂ����U\M���b�k��٘�EdX��L�l|m�QD[��1���9X�U�`1�)F��D]�C}���8�L�r��Gǋ�sz�y�w�jT�Eu���
1��s/�=$����l��������-�~�f7�N�90ʸa÷''�'�l$�10zHA��I���a�m&��M�y<�&�)<�n�J�[Im)j�<�vbӉ�i8�m2t������˽;�-w��qٹ�Åp�M993�T���[o�6���1����v}�̉���uu��bU2؈��������	��I6{�>N9�e�#L���؃���)�g4ky���d(��
8p�h=�ʟ[�_*�5�)ó���-L°F��6�/^y�N���AiC��Ou���&�g��ҧM�M��|<�*_~���M
lOJ|zp8i:��\m�sN~U����#F8�#����]Q�R>C�� �R��ȩ�Y-�|%�:�L��\n�#�[]%v����7`� �4��9��wA��!$��	�:t�)�*��ۨ{U�{ĺ���7��5�t�_s�{��g;D�xd6�Zp��$$���a)���!!8��i:�x)�)�Á�n����l���4�CR����̦��O�碪�#'�Z$f;�&[K�}M�<�<�N��Z�G�:��$�!F�i��y8�\�������e6x���D<Q���F��X�YC�4�a0x���2�y>�����_��H��zg�S��*�۽6�Ԥ�l�&'^%�I �����׏�����u(((�l���~����dc�#>��[�%������3��O����|�p�Mx�aW�G�oC�zNm)�q�N��́��r!*e5�7RTч�u5=4`P��t��N>w0QLk�#]���9��M�ӌ���h��f<��3qDU[M�n�@���S���ǌQ��Yx�`�Z�#�2�rj&�iJ��[ �De��c+i�%E��GQ���|�6^��3��:�~a��<�m�ױ��]\�u��d$6�U�I��B�ێw0�i4n�L�sR���5t�R�f�4�O\�l�O���<{��[�=���
�8SF��u�y6�O��Đ1Ɂ;�����S��r����x�+���J
�kJ�eO�i�ƓDmc���=���~:�W��֪-�m
�ԉg��2����i�u6��{���L��2ó���U�'N�K���Ӗ�i�M6e�nZl�:2B�(^B�
P�V�b!j���.�9e�<[��̰��2d˶Xa�̲�-�:;0vv»;9.HHHZ�	�xLR'���B�,W��g~��/�yu�{�����iKs0W���AfkZ�V��1K���g�ձ��my�=���GԾ_M��Sq}ߴ�>��l��h��x*��9�-]��̝�����uUL�ww����US=�����sꪩ���wwt�UT�ww���z��{����{�
К)ӧ��E�^��i��aܸu�\���eI�Y�j� ���oy�:���]��be8�<��o_%����[|�fKL�g����
pO�p������{t;�zS�5��h�������3�˩U\�b�ߡL�~��7�p��fcK�_<��=!�*�XnCP�9=����9Q�7��nI��J�>���'sNOg��\�%
�<)��o-�jk�7zqD�-�֓̋���eshs�N9�Z�w8�6h�0��q�S��ǂ%��b+�N�˘�r,p��"�[B
�`�]&�5�ER�eV��&����!m3�Q���u0�8I.��1m�:�M��I'�B%�j[0�X3 �����Սxk��M�GT�F��ȳω�26P�FHl����xB����JÅ�8���N|�����sD�Bi4�p���z��3W0�p1季K�P�m�Gx�봉�O��1��R@���K���M�'ǥ
К)�ٜ�~s�M�#�X�ty��j0��wG-��ra�`o5�h=M�kB��e��'(�o�ӱ�i)�ɳ��C�'�ui���eC%2.f���.�L4��3�z�fY�R��m--�����P�;�"W�!3��a8���KO�oR�%�^�m��'X��q-��0� �&�B��$8���r��aAFHx��Rř�{�,��,����I�2ϖ2��o2L�=���wN�ێ��`��dL`�l�\Ĩ�)�`�����.E�r[]�3��(�L),��ٯm�R�c&���u�nf.��a�gp�MMz�4�O��2�R�N��x�����l�v2�(FS�fSU�s+r��n~��d���Q�h�
П��l����h͓!��<3�DD2��HI$�q֜	�(�(�:M�ɓGU����C�<j�� �Ҙ\��X�3�1W-����I#mǉ�)�eɹQ��`)8R�
pO�t�l�䆐'�m�Ec�<�-)/��$$�&�љ��q̸����5�p�ٮe����a0�0xp��ҭ0�y� s��;�C���(S�xS�a�3e�1��a�m�04�(]v�Wur��A�۞�f���eL����3��Ow�n�v��4�Jy���P��I1�����Hۮ%<���A�A�g�R"��ꪪ�F�H+�g�}�؟����K���f�U�	ٚEh����{�[�^R��Uj����D�"���,`�U��,BJ�����%N�Y�&�#m�b*K*J),��Qh�F�(�E�R�YEX��QF�`���E�-(��Z,QKT�EP�X��R�(�E�aH�(�X��QEQb�(�l�QR�EEQeQe(��#���YEJ,QeQ�ԍ��E��YE�*QE,1R1C��0-P� 1�2��}4#@Pލ�EQb�QE(��(�E�T�
,QEQb�(�E�T��R0Qb�(�EYE�*QQE�0�bQb�(�E�X��*QeRKYEE*T�b�,�eJ*%�,T��,S1 ��0H#1 �%K,�EK*T�ED�RʖT���**T�eJ*X�c�c)$��A�0F#$��0`��F$A"Fi
�E#�F�*X�QR�J*%��T�RʔT�K**X�eD�#$1"F	$EK*%��%K,�EK,T�R��J�b�,�eK*X�J�*X�ED�Rʖ*QR�J)e,R�,Q*R�*)e,R�,R�TR�%���YK)e(���%��)KK)b����ZZK)T���F"�R�R�R�e,�U,���*�R�b�(�K��K�K%,R���b�)b�V*�UX���R,�dU��U�����S�D`�����#"1UR,�EY*��X�d��$#"0FȌ ��$#"��"#P"��#"���U%QKUb�U���RA ��#"�dI��2#dF#$�`�"0D�Ȍ�)�b�U���Ub�A�#`���#"�"�TUU��U��U��$"��DF#`�A�1"#H��R�I2#H#`�����V*ʱV*�V*�TUT�IV*�Y*��X�EH�V*�T�*�K%QV*EU��VJY*��T�"�X�%R�*�XUU��R,U*���
���Ub�*E��V*�UV*�0F#"H$A�0DF�#`��F#�" �KR,����)�H�"�d�H��E�T,"�"�`)��"���"�XA`��"�X�AcpT�`	 �b)�,
�X��`�
0X��b��*z�n�@�5�b��BP�)������BAE#0L��J��?/��痿=~ǫ�}������t��Ojo�=����}�����=}���'i�g�+z��ˈ�K����G>V���~^|o�k�����^���}Q�������<��O\�?���	$��'��ߏ�}�����C�$����>�P�H?(bT�������u��g�/ʇ��?���I�j?�m�jM����_��د�>wo܄�A}������մ�1̘O��HzCi��y��}�b~�h���))?Zo�8�4�5�9��.��G�z>�v�l�6��޸��Q�?�������L�EZ*�"�l� �0�CID	����(.6d?P�-i��V��t�����69-I��k�7O&�(��I%��Z*�-HNhI�*��U E�������ʚG);��Ϝ�~�>y�O�8T���G�R�˶��~�Y������=��d$�G��7D������Q��?����?_���a�k�;��l����r>c���G	�����+�|����>/ѯ���O��O�	$�ڟ5"��O��Ik��c��|���/�\'�'�{j !����$�|�Y'���~�O�m����_$�9nv�^b���S�t
9r��IHO�$��X�K��D`))��r�M��'062���)�o@���z����7����.	ȼ�C�TbC�g�m���yD���s�BI ����ő~���ԏ=����o���I��{#�b=b5�=6��S鏔�z'���i/�'�#�a_;�O�?z{���o$�{���i�)R~o�JID�p|�^���g�g�'��7�=�jy#�;����'1jWU|x�MۊY��n��l�	t�L�M>-���|�I��w�<��6}\�>Ro6����׼�	$���K����[Ř�{���؟K	�o�'�d�N��{��N����E��oF"�z���ԜE����}��H��d~q^�ґ����'�~8
�?�~I����O��������{޳����>
�ьA�RX�yG�����]��BB%ބ 