BZh91AY&SY� �_ߔRyg����߰����  ``>u��     �=�x P(C;� ���:}�\x={�U@� �� �@�
	2��0 � �J(  X�$�2 � d� � ��� 	 	 l��` ��h�>��	(�     f�Q!D�&���5?R2?UR�d4р���Ѧ� ��S�i���       �!4F&��z*?D��A���i��@�ВJ�12` L���#%$�F�d	����&�M��hh!�F�DiJE4ښ44� �h h�z}�U�N��D���p��TQ�~̹*�J��@�GQv�������$�H�o;��|�_ ����I2���;���������Z�Ļ�^5 "F���TA�p����+α^m7��wf�m��e?N/6u�yh�^l�|�g���#����.a�8��)�,܍�����
���t��s�l��5�����S~�[-tg�}���|3өr��:j� �R_�K���W�z�iO'�筪�KÖ{����;+X�	i��m<������JE4č���vÅ���
ZbgZ����<��-�;����
�[7���L�hg��ӒTHG�)�p������2ʃ�1�������=wV��ShGU��̊�''hc���z1��N���V�1K��OL�Ī����;��tV�Dt�7VS��'e�%t�cE˛B:�b�6T���eGF�Tl��F\S�i�iɘq2RvTzvR��=Q[�x{�.V.\pfi�q�ٶ(ʏ�J�!˳|j�u��9.w%�U���З���.����{�O	Z�zy=9�����t`�_vU��GQ�)�h�[�v��u�L��bF�	K3�TL!��e�j����mj�0e-UX���d�roJ�窙h̛�S㒞�t|[�;���Y��=#⧅6���s�9��$=�$3[�!��),+�����5M��� �����j�Cg�Þ/Y��}13�a�����s�[����;��̸ٍ̙�L�:0e�|�;Ī=*�<Ǒ���N����rws%���Q���7��	vW�;"l�T�h��F�3wC���PЇcG�B2�=а�HFl�B��}E'�-��e#9���r�\z>3��iiiܨt�s��:C�H���b#�VŞ��zs]��s���1�U8`:�#��=��=s`;���5Q.$����z_�p�����x.p*40h�m�\��c=я�SJד�.o�n�u�W6�] fp��1��c=���^�x�3�u�ʴ���UKtt��ׅ�J}9ԯt�Ҳ����Kڒ�Ԯj^�K��=	�d��R\ѥ��7��=��:ϙ�bO��'�ʞ��gNC�9����>���O��L�*�;<�R��\�Xʰ������U>�S���3�Uz;<h'm��|���A��R	�a�@2�1<�Iie��Q�8���-��UC���=���&����Mow~&�]�ǽz陸
�WzɂĂ8�����f���z�f�ݘ�P�c�R��&v?N��r�m�H��f2�U�BJ�Q]+	7[}ɫ�ua4��	��Ś�c��rPI��H@a}�^��]�8X�ȟ���i6.��!�~�D�n�M��iq�3p�OH�Ò7��@<+I+�aA�(���xIi��4�[�6���5��F��%��[�U��8���
���u��dʊ��.P��1Lb@B���p���:ˍ�9�f]T��)�L(t����4�z�͕K��\����~A����lc�
�?X��ݛ����,e�>�\��f3���uK�wۂI�����7k�Ϋ�d�X�|=�s;�@X<�0�֤U���9���If]��]M��j�*{k©-�$��A��at�D�p��}�a<��5�(%��1�~~��${�)a-/N�i��bz��L���\��ӷ��:I�M�QD�������H��tEYG�A�پ<����|V����B!T|iF��P>�鋝�Q���k��]'�������xkD��,z�vWg"�A���u�,R�{4�aGM,�P
a#0"�	���A����b[L�n�tn3����ٷw\ѕn���������AG���
]D0�/�ی�d=/���W�r��L��	74FV"���U���|��[I��aƠh��Y�Y�,��zJ���fa	un!�����&�Nۘp38�R����Ǎ}] C4�W3q�\�^�*$jOf��2��}�C5�K�Ŝы�6����J޹ފ��p),c��\����ww�^2������t��CYTgq����ٺf��4�ZE8t�u��1���3�t�U��"]Gt0�#j�E�l#�:����Y�N���y��n+@�r�,���4;\ե��ӱn��Ǔ�d&�c Ŧǋ/]�--mS��9���Y��p�t��Cdn_�n���f���\��e��!��6��1��2�u7><*��3&C\(r�郦-MyUjD�k5����[�ų2�T���O"e���(G~�{�~��6Q�>�Bf����=��L��6���"�����GC����j-EF�\�C,u���+]d!bth������ʭUIu�iש�dl(�C��@�@�`�S�6륲�q��W���@�����"����hb�s��Ԓn�X��I�5u+�8���`c�K\n�	efJ�� E�Q�
Kls �
㛺G��U!Y�ʁӕ�	��G�RF��r�Ȥ�[-3Z �"rZ��o����a�j|���G�H`�m�F>��2�ε�j�q�c��8Q�֪`v-���"c-B��i�v�C��w��`��mpU����$X^��=q��A��$D[.�ԫ%N֋�?����N�饂��	�d����m��H���'���	�h��0��h$!$���_{T}\H`��\ϡ4~�/�O�j�y�5$�,ʭ��|&rf<�7|dHђpJ��7�w����?ʪ��U^�+UKUU��VՊ���rQ3�uS���L7��U|�UWȭU**�����������J����UT�h� ֧����y���ҬW�*����R�*��U|��	�$��tѶ�յsNj�W~�m&�IP֬�T$ӵ��qU�jұW�V��]��*�Uq\�L�)�;��c��h��V�d�J���Z��J�5��SA�l�o/ݵU�^*�UqEy��UmW��{}�t6�	��M���҆���!�UCAD�R��Ǌ��Ux�ڋ�{�Uq]����[�@�`�bB1a����@���#���5�SN���Ҫ�V�V�x�;۱UW�J��W5�5�����A�I��$�RN5�JW�x�UWȪ�+�]�{b���UU|���I^�\1�4�Cc��&�"m��	1�1�2r6�r%�B�e�Ͷ�O��z����#�&:��������Ђ���������˛��T��g&���˕.\�s��Ó#��Fz1�eON̏!q�Q�Q�֘jU�����jx��q�¡���V��Բ�6YZ�[UD�9mn�-d��X��:��Q�
ZHX)Uݵ�M���v�bM9 �%+e%jF�jp���*�j�t���RcMrDD�m��1���"�ޡ���&h�8�Q[�,Q��jN�&�ш���W%��Dӥ�u�J�v�#��W��2��IPK��5q|�������� ����88 ������kZֵBZֵ�j�"��kZ�!%Z�{��!� ��	4M�������$Q6�%���q8X��
Ԍ�t�h�i�\��B5JAD��D!��G�V�c2�_�	:J�1�FM��߈&)�C~�2�c�ž#sf�k�aE�p(����,�$���80ta�3�n1q	y�����(�G���mQ�꣚S%�}h��n��Y�N�:�*-���b����i�6�&����Ih�
����u�4���8Q�J
7���!��J$�NK�
��eLL�V�Ih��(��X���\m�J�6�B���$��ݾZ"�cm�ͪ)�Gk2>1����q�P6�RS*2i��9Q8p8�C�����B2it���is[,�4�([S�s�T1��#���(R���!��%a&��q�敖���6�#�mqZ'j��ZG�*�q$�s*%�ԍ�	�����A��Q&�,)H����fQ!)��KjMrC�߂���"& 1t��'�҈~��\dbբ���'L:IAF��mB��p�;"!��,!�)7ތl��k[ZK����ݨF�W��l6ie�b��IU�n?Jc��C[R*��{�j��R�Mk[�j�n�T�d�VZ� �j�u;eU*+���>�u3538���˔�@uY��F6�/Q��(gLR��Y�%C��������e ��n-55ҋRB�$jFJ6�1;ѥ�Jͭ&�o�{D�х���T��=�<>��!��������xQ���a�	���h�
0'�!�FD�8Ig���<G����C�$z���x��g���0xt��8��F�p�d��hxIF��0r<�/�h<N��;�e�ߪ�������{]��{���LCg��� �cq����xis��9��Gxta�o=z�$���{��)�ۃ���kරk���pk��r�� B�� # 7���ӹ�x��s�K��j�d1�����5h��m9`�|m�&���p�>�!m1���LjRiH1LW'� ���&�ơ16��^�D��(&���P�4+�a����-#��iqP�ii�R�к��g�5tI�H(���o��D��KO==�hV�59$N�Ox�ޙ�E KU�ĲjR��D&"ᛏK���M(��{�"cAG!
ΜMHtj�P�/B ZilM(�H��466���14���KB�J]4x�2�.FV�AI�����J$���%L8��"ZhkJi4���	�4��A�r7qT�	�E�Ac$��L<i�43��qJ�$��D
,��?U���m@����A��mY	hk��}z�9��fF�ibibh(��6�:�@�L� l��J$�f�_��F�p(�]��q���h�A%��`�'|'IJ�EN� Գ<0:�Ucm@pem�J]M44+i[�)�g�0h��	Jh4�-�m4�g�Y�Iq0f�<A����Z���<��G���1A�4�%�-u��e�UM�),V�K8�6ӈ��:�,h�Q��6�7���6�k��ML�����4������
QI�lcM�*�#DA9h�l��1�(E�,�g:XV���lHF�!l��Z =�B�ץ�.�!@�wжĸ{�68'����Țw7={A&/xf��Lh0��0�	J1�G�8Y�z;PL�RH��m�Ѿ�yB!
[M[:��������AH�ư��!�ގB�8��,P%�D���p��4�m�����P��4a�]M�D����0R���@msp��)i��î�T����F��i9P���4�i���m���a�ĞW;CG��b�i��0��8<��a�	�xp�4D� �0�0�(�ȡ��o"���Dh~6l��g�^�~	��?#t�1��n<ON��lrx�o�$~��$�.�e�=�>W�1�uȯ�1�&�"�-�ô�ׯ{�����g�e/3��=S[5��������#lGq��Λ�b�ꎡ�M�	3A|-�p��4�h�BC /b��h\��M��s�c~� ꛾͡���sV����nuX����s Ķ.�dȑ[7�\��p�����oǢ�n�TcC�Y�.'p8�PuB��i�յk��*w^��I��6J K`cs'	�
�*�{"�ق�Ԗ�(����-jWK	N�G� ?  >����m��-�Z�-�Z�-�Z�-�Z�m���m��8�P��W�+�&��r��ٶ���:�D�\,�ӱG]�U8��K6Tć2�)E*	&F��m��4XqH-Z�1�A�{��-��ɥgf6mm.���7��o���-�8�d�TZ������!J �dl�'B�Z+�!�������0��6�p�j��cM�ᆊ��qjd�0��O+E,�	,,���Ijb[g'!�׍����TDD"B��06?)�� �����yB=*�Py�w�gZH��cl�<�I,��$�YGx5 �D�(;L��3!�5�i��Z�j" �V��A�)[��\���HkBj$^o ���	���P�A1@���I`�0���N��I!���DR���I�AFH����CkђYs�՞|K���ި%_U�Xj%��9�Q�T(R�*�%�C�V���I
�%R�'���<1���42�8<5C�բԅ(Ӆi�h�h�F(
�:i��i\������2M���A6�c	�U*	ZT����M�Y�$��o��]b3� in(���Ãm�Cy��,[H��#h�Rh�
��"� � �\Z���:A&�͹o�*H���CRmQ"�cccm��aTu@S:���qQ�T��ţ��^X�U��ah����l�I0�� �z�%�
p@S��������k$��yT�AZr8I8q�$-��);K%��M�K�,��>�	%x�	V��!IJ�^\RJ8Nyt�л*Ԇ�[�G������N)��GM.���KH�8ID�XYh�MF�I��5�1.� i��P:"�������.�&�@I>��ʥ��6J�6mL0R�6��1��f�EI�${<C����lxz����ل����ي`�a�p�0�(�
cqFaP�
#���h�#g�<p����x��!�#a�8l��F������	��ro��K���ЇͰυ�Y;���[��2kPN�Y���1܌�;��|�z��Zֵ��[m�m��<�r�m���nR-�W�A�MAad!s^�F�KB����'aӉ��M16Զ��"H�����|�y�4hh�kiuqP04�X�P�-�0�𣄜$�Ae7褕'�M�Zڰ�l�E�T�q#˒H��/A���yXupđJ���f��UI�
��Å�ÐPb,�5!��>,��$����;U�T�>/��j��!U-"P%�b�8b
IoګISN(���dD����ThUC���=��)qV�R�փz�!�����ll�p���a�a���)��S*�*
WŶ7�k2�$���t�m%ĘZ��6�	GU($-Z�M 40��T�%��0���`s*f1�G	R��T��Aҍ)A�v� �ՇM4IB�㭶�V
�(\4�X�G!y7�`�qs1T����@��',�Iu8�څ�j����L���QF��4�:a�AagT��̫�q�Y߮ ;�4dmι�Y׀ 8[(��@��Z�Hu�$c�T7�4�#�tfΉ�G����ţ�߃�N�0�����qΩDD5ET��BH�j�F��Н�-��Ņ�E�9�bl�ѥ��N#k˦�.,T�K<�����i{K�Q�g�$�J�U�1�72�̐m�<�/So�-m_��U�<t�F�ag=�2Ƅe�x^JV-��F�2f�RI⃩�5��<���ĞRY���h��oKGpo��#t�ACJ͝,��XX��m��@�(6�"�sm�<t�f/)hpt���!��^=��DH�1n�#I�F�jUARG�c{�6J$��&J&ΔPͅ���s"&�P�MC����b���&��6i-�R$��V`ݑ]�b�iqm�3�6�uqZ�y]�k�R�ml�6�G����6=��G�`�Ǌ��sß��(�G��!�A�N�VE��P��(�0�l��aDɢ4=����a+���'�0~<A������oc��c¡�����=�K7'(�]����j�=�/58��	W�1!���M��&��& �!p={����c�Ly�s�:vl��Q�e�":��Ǧ��D�w8r)�ѩ�z[�Sw{��i�ٳ	��4H�$����d2��,��7{~>���Ԇ^�0��s0��$4�Q��1�,��̝ݲ@��,���RD�h�N�q��lN�*�+�75�k�P%2��R��*���;D��"p<otjG� 7��φ�m��m��E��m��m��m��`�� �{|��,�!i�m PUG#���."ˣp��*��Y[VՈ����00hn-�*�yp�RU|<��Fl��(�5%��tT��KJ�m�����Kdɦ{0��>�@�20G���Q�J�$�$�Ph,�\�PhGE�D�uJYթ7�H�����I$�}�&aKll�^��>�WQ�k��y��m�F�OX�Ǣ�:��k�6I������1�J�Ѧ�����]�y�cmѝ7Ҏp�3��� ��R�ŋ� �b6oA*���)Dp��Yݒ47�E4h�Y'	4P!��)��:�cO=�k�W���g� ��.:��%-�-e�./V��m�]�e�ml��4mb�g$�l,}~�Lil���,NՓ� 8��#sqh1ra�3
59Y�qT CÂCB	a.\�-��2 �("�-"ղIj��"#nf5�,��(<�:)ZB7�a�Q�D�0�" !��i���d�g�5(g��I8v��Zg	!��GPJgxQ�*��9ߣ���E+N:	�KW]���γU�[9�V�W�g�<I��Y��Y�X2����È����2L[4h�,��nX�eÇ��6i-�,�����(F�i�"��I�h,,�e���:>�/cpyF��x�p�P{k�1���J��ps���_D�N,�92F<�[C� 6�[8y��Aӈ�d�$�����D�W��w.�vn�i�z��"� {�0+���պ�QY�i��Gq�؉�U�Ú��F�mL��3f��K�j�yzW6�	R��م�l����6A���ԙ� ;�-�f��c���5�1��$�M�YB ��LIJ
U	քx�a�Rup��{C⡭���6�貗��h��VAX����R�]I��ǳ��S<�Zm���g
]���<�6>��<0�px;0�t��GF`ل3����m��EKv;<E#�C~�dP���f���1��I�H��xx���xx�O'c��I>����{�m��_'��o_�z!^y�y�~��C��v�m��m��m��m��m��Zֵ�&h�M���H�G��|�=��Y�g�&�I��"σ{]Tlܜ(�������e���t��$��X��!�L�h����ʈPia��:@2Q}GW��-0軃�͐k��''b�:�P0ߪ�d#��u�%�bୋ�4xk�T�-��B ��&�����!��X��ٱ�h�@Z��+!�Z�Q��j�ih��2QjW��P� ��!��VDT����s3J\��g-��I(�񳇉4+q��H�
�F��L��֔���'�9:af�ѪLg���9؆�Ԓ�daD�J��f���Oa%���tjdj�buW�.[oD����2�ֈL��(�Ryk����#��xp��Q:G�H���0��Ie)!6�KKR�W�x��I86��d�E�3D|�q��VA�-0�=�P�F�+m�3KN�5�xDX]��+%����Z�Z\J�[��3͸l�N.�tmؙ:'�b�ɥ�TC	�0MKN�-�;�pȻ�n�G\"����Z�J��D�&�G����a�%XfB����dd�˗�"L-zͩ,�hᄖ
3܅b8kJ	K6J-pe,)#g��3�9v����Fյ&׺�~�ME:���6�PA��<Te�6���&��6p6�|d4��[����  ʴ�/|]dS���H��D1��d��$B�6Z�A�G�1yB�R4x擑a�G�o�p�S������*�6Y�<Y��5
J)�ȂG��.����P��܎���̸����H{��Lߏ��~h~ѿ7���ф��'f�с6a�0����1�[�ɄQ�aP�a���=�c�dh���$��0f���<<F����~,�â�0tQ��&�Jtix��"�`��ݭS��ƫ�b��<ցJ��+�[�,�m���i�yd��vtu�t����c�:�+�����N4O��� L�+�6�ˍ�i����DD���0q�T$ 957�;�o��խ�a[�Y.�Gm�F�v���M�1L�UDH&��,u�N�
J����˰i늸Jؤ��D����%��{��U��m�Z��Z��Z���m��m��(��A��!��M��V�(��6��;e�N��iJ�̑1IҨ6���jْ;MC�P��ǢZ=g�E��4j�f���F���R��xX���w��l��c�4m�(0�e�����+����imp�ll�2��X���ڣk��fM8a�%��N�ǟ@k4���S#�#j�6Xh(�-��o@5�KI����^ًB��q�F���.$��B9�����iqZX3x�8�5G�4l4Q~Qi<���&�� jQ�m�Vu�N�ll�D�4�G
� ���J-#��^%g��0�a�;n��1�@�
ȷn��QI�97^0C�[��8�̱��J�u�����%��G����L��jm����
Âg�+)��""6�+���%ӈƊTN���d�8�b�ս�<gN�� ���^���Y�Y�`�{]<l����X//#��s2Hɉc:��~Q�6q���,��n�<�E2
:t�2�>=��ݦ��������B[F�|�݃D�C����h����O���h�[:��L�A�qIC0�a��u�#v���v���F��mCcwM�Ě8�7�`^�����ң׍�\]R��i<ADb������f��FTܲ9v;a����<���8�4A�`�*�[��e�:�[T�RVZ�R�=��ťh�mvh��|�dLȴm�ZV�m6֖�0���AY�LB��:��mh��=�p�!�D��Mq>�V���Migy�,�-�����֊���!5�g�$�KX���qT-�S�zl�2c6��8�x?���g(���	����0�aa2����,qc��¡��H�d�ǣdx�og��}#���x����`�p�;��<ܑC���tQ��gώ�o�A��n*��;j�N���6���^�٨�{��b��ښ�jFw��t[m��m���m��m��m��yEQ�`��Q���3R���W��~㈍�!	���Q�>D�ԣ�*>Z�ж�]C8�T_NY�C�7�#^�8�7�����!�ŷ��m4m�n <]&�-�܇�q�������8�L�(��S"*e!�E���p�l+�����dF��r����7����&v�\����H��Y8b�z��"K���4j��Ia�&q"�1�a��h�'K �a����� [��F�;�a�/"��ViG ��]��R�K�����/�8����͕����8���8XXv����N�!HgNCm�qk���N�C\E�y�lf�Ƭ�ՠ2VA��-f5 �m�#��hѵ�f� �ah�o+�Zmy��[[\`K)q5�>Hť���R�KWfm4b=�h��0�XZ�MB�����%o5���fV�Q�k��e�I����R��Ђa����<�m�m��r����7ͮ�Kh�(�Od�X������oƑ�>�p�IT.��ߗH6AF�Uv��x������ܸzZ^F�+�//+�眝��ۇ`ծ��X�x�f�V���h�'H<h6���."֑�y�e٤^�����L�s6��12��Tח,��om1uj���x�߶� �"�:h�����D5�ѭ]�)x�Tu��m�*I��&��J�m��(}DPxk��!h�6�Cz^�x��Y�!w�C��$c�m��6CG�N�f���hr`F�C0�0�xE�AaaT;#�vh�#C4x�#���<>��0�0f#���`�p�7-��B��0taxz��:~�yroɳ���1d���Փpm�����%ϯl�̎��^P�� y��3 ��ADN�u�mwv�"�:�Cv�������$va�ţ�B�`����o��q7,Z��H�3qj�A���-]��]��}�%#""U{r���DÂ8����"Ǐ�&t�[���U1£�܂��~S&���ޭB��!wqN��cj�H�Ej2H��D���G~y����Q���>W�Ɖ���nZ�ISht�eȂ�0�Lr5N�b7@2(��H�p��+�\)HЮW4�Ghj[�����}|���m��m��m��m�[l��m�EQ �>����|R K.9�j����cL�U2J�"N�ؔ�� tts�j�8�ɂ��D��Ɂ�c:ܣ���!�R����掯� ���F#�H�,�"j6��Gy�n`!�Ta��6X`roJ�8�[$��-i����V2�b8aª�c����k�83e��y4�+l�a�PrT%H�Y�toDDDh1l�m����#�J��y��4�6R^Rl��В�6���Bf����h�:zFY�TZ�����H��o��P䪛�P��/'���!ywH�
�� �B*�#JB��&�-�a$:�����`�>�vFI�P7Pv*v� ��f�5�S[�E��V�i�F�U�	��8�du��{��<X��q�فj�J���Gh�6oO��4�p���ލ��q9��b�:��$�Q�=4��h�J��<�10[�q͍k��K@f�Ä����(����Ȃ�#C^���q�XG���9��J����'jވ<zW3�!]�ѳ��:p,�i��Rk�:'�V��B�	������5H�ՍmR�M�����
�a�x��&'��kv�]����浺��$7u�+E�kjAWl�ƤU�GS��J�68�l��Wx�zmGX6v��f���.��U�)�Da�l{(���C48h��#g)�t)���5�0���'�%�fiH�n�'�X���b�kˆ֎���W�*�t��3�5'���m���G��]Di��ӧ�DL��$���3#�2���FFF'H8I҉:J��IGH,��,��xl�t�ӧL:a�f�6h�L �<>I�:J�p�[��n���]�\{�Qz����ٷ�.�0�ۥ{�nI��W��~�V��;�K�$^��D����;|q��d���S�����B*	���K��O����3g��纷k��~��36�m��m��m��m��m��m��o�� gr�sW��<���m��mC�CmI�b��(��Gz�
5ᤱFZ��IaFz �׵|h��7�Vyp�,�~TC.y�*�qJ�#����ޗ3QN�c�h�'���}6��m�a����U�����CKY`�e�!�l�ʩK\qHڰ��E��PC�K�kkF�ծ����<���%�#����r���CK����뙘�l�qN�2�&i3�I$�Q�H�yiw�cz\\4ON�4uC:����b|*a�L��Yn�w˃�H��^�`����0�M���08I ߸����h���F�|�D��a��Cx�Q�h�iu ١ͷ08�h��e�IaKW����Ed�.!ÈpS�H��"ф�ՊU#^&�׍�f�(�[�g��6�,:Id�{E������^@�q9X�U1�V2i�.�h�Y��'A#q>��0�✆ۈ��>Z�muH֒���!��!O��Y���&���cxDD5����� ƪ�E�W$��E\^k��zŤiuZ��F�Ȇ�n80n,��@��q<Fp�F�:���8I��4���p3#r�mJڱb�6ܮ�wj;$�I�!�.G�=�um6��6��*N�G��%e�[��l<�� ��6D��pL��\8�O\C�D�s��o~�	pӒV#�l�D&l���6�mz᭷j�%6_o�87-�)�f)?8�<;y�H�Mz
��38���m����l��.Qt�~O��_���흻y�U�5��>���;�8맃�Z�Z�IT��Bw�Q�D�+�)����[+e6��ڶx��.��:��`Ɩ5LicU��#1���1�5ь��.F5XэLicSc,j��c��F4X�ƫ��ƫ�i1�\�5�cC�hcQ�dƖ9��E�I�F4��cU�F41�cS1q1�XŌ��5X��s&1�����Ʀ0c#�.K���ь��cKƌ�����F5chƦ4ƝN����t�t�sM��kka��wc�-b��X�b�a���5��\'S��X4ÌNLM1u�	Նcc1a�28��a����X�L1��a������LY�[6�f�muìc1e�a�9��fbq���8���f5�14����k`�31i���Z�Yi�Y�Z��LM3����VcL�����ns��ý���4Ƙ��5�L��bi��i��Ʊ5�f�Yk-`��3e�F�k3-0k3-2�4��Ze�������f��[5�����e��F��Z�ek5���)����5��k��k-2�ư�V��6�f�V-,Xb�ţ��ab�b�aj4��4��Ƙ�Ɩ11����.�wp�1��1�1�1�k�\1e�+��X�Ʀ4���V4����D��0>0���A��4��ݭBE�5�q;�7]�?[�ӯ��PZeBBc�m�k|"$^���n��.�Z�}�"�`QGh�A� �(̽4E���]3��41�Ml?4T��� e���h C���6�(��*���@?2ؔ�
.]d�� S4�7�=d�̇��{$�"��b$�Y5S�āA���:��;[;�J�t}4R���2|cU
5�%��`��t~��ֿ.�|R}����C��'ܚr���}Y=_��6�0��H �xΟQ����5�5�c:DO����������O{��|�fc���Z;c�jx;.�r����ؽ���l],�:��S��_�NNO�/&�����RԆWl�9���cg����&�)@1������$"�����TJgN����$:��4	;]D�<�E�F��l'�ԧM.��qi(̧1T�h]�N��0�t�c��xd��B�MsN�B�,ҡ�:�A`��;X�x0��flf"����UNb��D9�`�O}�����;��/q;��������B,	�/5V��U�<�^�5�U@�a@I�2A�ʝ��F�O�~7s���'��\�(�|��L�$�%�,-4j�a�ۈ͂,������t�����=��>C�o�;����#/ja�������.��"Y$t+z�_;�.<C7�I �`+��3M`���r�:����A�eCY�x<��}���sS3�{����JQ������_l��`������̤}�B�a�G�TP���?x�I��9�0�<(����*Wr�ci���՜�u�q^��{�sUR�:W��7��y^2x�-^o�ˮe�N-�9Oaϗ�B:"�9J�4�jXK(��Ų��L�6m�n�Nǒ}甑G�����f�3��;�C�C|�J���U
=���w��eX��~���~7���,]����U�t����&z#�&)	О�|�υۋ|��|�N}|G�y/���h;>O�;O��q+�~����ܟ����T(�;'Z�z��I͙o�8���������Q������7�O�~B�ph#���;��M��F *���xyvO{�3Z��Mf}ƻ��2�wm�ݝ�t�-����zX���E�p��X#a�lb)��-���pF�>è��*�B,_X��_O�a���(Q���������ɸ��:���[HJ@b"1��pX0g�y�^jF� �#��K�l������QN=x���1�k�N<ҽ��>��z�š��v,�����Ga�O'���O�o���W���u梕�>׭���c�X��Vkc�Z+��46����qCi�h����3����H��u��H�
�@�`