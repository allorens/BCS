BZh91AY&SY��6P�_�py����߰����  a8�����F���
����H,Ԫ���ɶ@ 3MM��B���   �* U@�R�� J�T� �g�UBQҁ�=G����D� ;�  (�%E    ���)@�xtm�g�N�h�z�P
>�@=�����[� h�t8|�G��>����p�����(���R��rJr΋3��s5)J�7n��@ Q\ ޖ��x  ^��d4�QOwـ�`ғ;����zi�֥ݸ�ìlV-5;��)�C�PP �|�^A��)�!b�h� �����w�E�(]�z��  n��||�(���J�F� �c��7aAE(��p7��I��4> U���mE�a�Cwv�B�z���=]�v&v�J�	� z7�p��Ô�� h�[i��ý��J4[$���0:kv�����{P��)���4R��0�4�uZ(����� >y�=�  ���T���^���ӡv2PU-�r4�_ �0�z�����:z4��4�iB��;U8                       *��47��URM0�`&L�  ����h)*�OSM0	��i�� ` ��%)$�z��b   �   z!*�`  ���`  )#Dj��52cTƚ56��'����*~��"�)R�&F�	�� h�O�?_������͋S�j��{��iV4}I��~��"���q��u��� T�"�G�F >ϸ�P����Q�ރo��
���@�@T �P�Q�a�`Rr�����D�2'�y��'��X"����G��_��~o����~���9ðr�#�~�_�wOa�=�f��p0�������F���N��/�C��OˣnVrI+��!�}�8kd�g���t'��/�	�|8s�P�p�x]�/��N
�,G�<9�H���`󌬧7O�u>��D�5����˩ֹwk��c�.Mb^��iI-��7-��5�'x�ZzW�3��9�^�g�ĕ�Ru���?I<�K�5����.�]f�'1j��&�'�f�z��.��4��I�3_���kr��^7�H�kˢ)�^0��a��xņz�I0�wj��-��$�-Y<���Mf�鲸h���ù��vW�݅p��
�3Il�/-��~���It�4��f���������N'��q����2SV�a��8��xa�.,�]3�+���`xʃ�u�Åw��>+��N0�s�0÷�<Ix��s��������&ĞD���4m�HOp�Iv�[���j88,�(uQHW�u�:j\,`�80;�Bh%ĂhQ8d:'���m��c��tl�ف���+80y� ,.)7ǇCC�vø���Xt{��ҴM/׸--	G�Y�����ф��`�}i`�
���%���;YX8vpN$w�N�9!<9�����I���̶�.ӳ=c��1Y�l�c���ZH�p�$w��0�Y����N<<0�Ө�8�8�ffg,�
& �D
�	��tI�I�I���w���I����WG����aX�INԟbO�(hX�V�\���:'aOv�}�[▓��lr<�Ø{Oi�a5F�|��9�V��tm2�$@;�z�+��J��r[��_%tM��)�!����+��Ҹ'�7� �H�I.�4�����}�pā���L���{Y���G,�s�3��/9../-�b
�'��}`�'P6���N�t,r漳w����V�b���z�Ş�cΎh�0��ݗ�t�����r1�:Õ��0���t�kǗ�~ö]`���}\�9XB���{�y"m�
����$p�u|3p�᣷I;��^a�H�I�gs��&��h]q-��&�L�vƾ'H,e�/	����,o�Xc�k��mC&p+�;��`{���یn����73���t�:ǋ�ߌ#V`���
���ŗ�\��K�r�ٚ����KW<�=�{.��?%����a�/�Z���g�axU��c�8zL���|0y��a�,��b�,e�:�ݟ�kR]\K���O,���^�P�Lt81N;�{:88�F��+��g��X�gea��3�,K��������],Kν�K�|��u��k/-O�K��v���X�:���.����;X�|Y��_���ޖ%�9�,]Xݛ�/�˻�����;���Iyv�]�-~���Kē�v�弤��,^�|�S��ug�w%���,]�g�ū������y,Ir��b:YXFT��`�x����:�0�:>�tWpxw�2�yP補8a]���mيɩo�gҠ���7��Z<@��޷v�my=�O,Y��g��^�#��^,�
:��G�郃���³�c��p�hÈ��lh�9�;=��cc<�O�a��%�¬0ǐtFp].p�7�,`0p�hv��x��	�&SO��u�'d�1��2חC�����k�2!Ҙ�xdp�Eb��8f�B��a*�8+��Gk鋄���ԝ!���C���]����pp�X��G�C������2.|Û�|'�ڇ�ze��FVC�Bx;�`pػ�p=��p�h�hr���׈����p�� @��<�0����=i0�9�<.��v}ח]bO,Č�^[g�Ӽ��测�l˹3�b�)�˯3�I��$�zČ�w��?'Z�$�bL�厚�l��䎵��{ĞsX�.���u�ԝg$嘼�̓5�]�g�k٬ԼƳvN��Y��k=��x��~��3�svb��9fu.�g.�u�<�X��r�٬Խ������4P��#Ç=D.'��P��1']k=�jL�/6�wd�?f�"��TG��G�
c9���$�bG���f�R��Ƴ�'3��x�C���)�(��9���5&sX��k;�y�����՝]]�f'x���CX�{�/.������Ӗ��k�!��T�ܑN
�:����#���3�����r\Ze�ή2��������:1�X/�Č�y�Y�c�-G�{�<��g��'#@�����8b��<��$�<G]��c]mPgZ��i�Ƥ#fS�90���u=�X���y����k�bk9&��5�����c�6P�/��7��bv�b{��:��O!��Y氮��V0���2�Q-x�3�gZ�4��ƪڞ�Cg�Ϙ�H�4r�\�=����m5D��h
�G�����v����N��#}��t�qȏu��"��H��U�����4�H�3u�y���h@n��F�q�h��F�F"���
����ǨpͰ��"���O
�Ti�g�fvg���g��/�YTsW"4�<.�,��:�SFq=���zl�K'�#�{n#�#�#g����Օ|���}�N$U��SG�#�H���G���6OF�gġ#VU�#i���u"��YDв_�B����#�X��m<�G:%���$+�F�4�#"�"��$u$pt�}ѣ0��6�qɨ�(Dh��;�B<p`�xpβ�p����ܷ7�����i�h���gr��iru����Y��X���I��ݓ��ξ��gx��;8d˅�[�	����$������^u�I�%���~~޳[�Sx���H�5�խ�X�4��+�<8viP]�8q=�b�s:I�-O?g�~k4�M���?$u��;+�=�p��
gG�W��/u�Ä�+���: �,�$�s%�a�N0�	L���%�y��~Ď�\��y.��J�,����s�0²�aҧ(YN0�s�p�{�`c{�D��a�iዊb�?`3�-�&�%�5�%�l֭O��k���3O��(Y4(p�$W�u�:iPp��X��X���h2xpT�	����1čx:��ف�3y�<ȅ��lc���:0��3�]��N�7��a�M�a#���6A��xw�� �xX���pމX��
C�h'��ė��č�h�H�`���lBH��ppy�+�1zH���ヱ%����xJ�q��˶�<��ٞ��9d�zV�Ǉ�~�xW�G�#�����GyjAbAZA2�pp��m�V��d�jWq%)%Ԓ�Iu�v%�o�)\��<i+I.I.�>���K����KI�h��a�=�:z��B�tה�E"�"�U��u���=�Y\0��z�#�a�0�.���F	LQz,���i�O�]М�"4���^�
�l�Ѽ7�Ч�Op��Q�#�Ý�D{���)D��#����������>r|;���|�!�F,U����qj�g4� 9�t�d;I�+]FCy�:p�i�#�U����e��z�\�M��ay8������\b����G��ӵ�<��q���^?mæ�>��CVW?
4wq⧴�Xa̷��"-�ڨp����Z��e;|���6M B�ОE�M���$�p�
$����+0�L��ʪym�),?�P�q���$��nυa�Uј��K��m�����o9����
]t��f��f��l�D���5N�vI�>W �~`�5r�3������<(�cCL!�G��4�2[Wk��J$�f�t�^�- �ݢ�8)
��ސ 9��aWT-�)�*����UՇ*�>4oi�e���T�:�����m��HʱU$�:I��v����H�yjU�<h�"S(����9�n� [N�l�f�xq*���ͭ�n���J����Mi����c��T���_N�q��ݘY�d3����$�a�J͹2d�pçH���>y�Mqg~�ɤ
�V�үHr�l�E>N*)�L7S23�ΐ��IZk++铤����9B�XZ���2}��ajY6�b?8Q�\w�i��z���n���M}un��Nn�q&�M��ZF�6^+#O�����XSi󷹯*>q��8h�em�XG�Bh�	�c�
.o�'� S���TM�X{o.i�w����bg��~k�n>eP�QqG
���6̾�}�U7��i�Ш��Z|ɃU����O�i�������%G�ԱMX�s骫��\aMQr�U9-�s�>M5z�XS���h�4o8x������Ȓx���0���|@QQe$�eD�E-Y�{<�@߬��(P�����~��ʢ���I"��Ό�N���y��K��P#%�B��Iy��.�(��>�,9t��rLLр�8e��W�.ΐßk���7��_Ggh�:;�媵��Fi����gm�L�����u�ja҉<Ql.�x|0��έ7Vx�n��^p�F��h^�W�-y�	:p5�u�O�ܬ�����gR�k��Ξ8@Ԟ���ӇK>��D}�1,��H��F���Q� �L����Q����d���lRTt��#W�@�]͑��r��gk�V8|o>����E��:%�+p��!��a'��?P������P@]8��@cJf��z��$�:x$�ѻ�fQ>�~l�c��n���	L�������Kqq�px�8p�@�SG���]�fG��,�y�&V��e��qY�ʯ;�fe�Q��HjWM�gM �@����a��{i�����1(B?)��-B��5��,�J��^��)��8b��!�E 2�8h� ��j�K�r���������^p@W��*� ��{8�⯞�"���+l�A�4||����ӠDf�c�i[R�f�|�d��˕��?*��ʋ�|�H�؅�e�O���c4|����Vmf��tT>��"�,zQ���E��@p�%�����\p��6|*�J����@�]�.x� %W��!��./J@3����Iޝ<�J�=:Yf7�ˑ+ <]eB �y����jH�Q�� ]�m����Mo��_L���k�헶CM�=5̧�+��%d{�:h骧W��D�Ҍpl�4gI}��{:
�kQVI��8�_k��(�eҲ �<h���*��ǧ��$�m�=��hQ���6=��d�$�p�gK F����N�w	��,��c|~������[��Ə>�6x����%����o�,|h�
�`v�\$��ی ��l��vy|�Kti�t��W���,��'*�}�x�7��u	6M���B]�Ӛ��ޝ	٤:��b�U��g��ܒΒ��s�$���\p��3�2 ;������ge<�th�[�n&�������a� Iuc��晱��oK���kr�im5�㣥�J�/{sr�������f6l���i�Fe��ɣ�
JkF�3��(|�����ǆ�7b����j�0飇�v��4�
E���(j���զɂ&�ͧ�YEi���&7�4��֗�M\|��v�h�*a��,�ſ�U<6( N��۶���7��L�޳}�]�R2�]�i�|9T�*���H���d�v��nSv��ч
>��9X��ݝWFV�)�V�[#z�K|N���{Z𣹏�2Q�m�<tԲ�a�+t֕�����5�}��j�̹-�3�Ʃ�I'r:Z�k��D����<T�:a�\/|:i
1� �8bU��&��/��A$l�W#�a�=�xi��EU[�ֹ��[��|I���=�צ�Jr�2��Cf�>P�
	_�<8S�F>'M:t��3��Ft��~�}��Ӏ�FB�GL6h�D�:^���}���ׇ�J8�)�|>���N�^�������Za#J2�f�*3�L�3d�<UӅ#�3���N� ��0<=8ϝw6r����,ҧ]�8IGTtj������
#�XޖT�j;�tY�iҔ��FxbZz3�) ӄ)�盍�g|$�K(�e�+�#�t��&�����sa�x����k�6U�g�x�Q��|tѲ�4ag��$���m`��|��h��<\־�Oa��+X����C���G
6m�Y�s�(�؃��c�g��6=�m�e��(������ӒaF��cċ��*;vګ5G&�Y�+�|5u�HS���g��Fb�r��_�|Q��}+^�>>�t	��gl�:��症��6II������b&�GK(���r�l�)���E�+O�+iu�&���+�$��=��vl�	'I]fx$��Fm�x�%Z/���іpu�/�4p�$�Μ��2���$���9iZ�'N�p鷬�9V�Ex���ϒzuގ=�(�?s����4js�G�Q�K؋�1�2��kn�Q�d�0ڄ��<�~�;�[9�'Wʍ�ʅk���֥B9{_�_���x�����w1�+\�U(���eM�nTu��j�<eg��0�c{v���wG+�_0�rK	*9��}3M!�������><\�V @��{T���J��� |å&�x@��F�_d��6c�bH�&H]|��)6�/��[�7uYyu)U%���u�@7/k���7[���(��w�̹Ǐ��Q�~;g���w�"p�Δĺ:m<v��ʦe�q��]�,RU�0�t��eS��CH���+E�7�xr�ڌ����7��_<��W�d�� ��a3gV�Qä�j�����Yӯ��T�i�d��iS�tn�}x�ʄ�R��z�Ț�.��rP<�M�8B����s��.F}��ݟ�^MeQ.�$�w�>�Zuz�0�ǲ�p�������d�릞/^�`[�YVm�}e�4@�]T��d4�����;[ݏ���6�T��!��G3�iJ����P�2���KY\n���[R�Q��,��r�ˈ��A�7��4����A��y������Б�N�ytj�?��+��_��>g�F�'�����g�Q�$l���v�\P-�	Y��miJ[�w�M}Za��;tM�UV9P��<U
�=�ĸS��F��UfǨ���륹f��[v5�nHܓ�v����GEKhT9Q���֖�CT�X�@.z��2k�vg�F�"j<+h�����n
D"e�T�be�Y�[6=0B�1؀�VT9�b�7X_Q����5�\�h�-����4l.�`���J��8�S~Y�'_��8��'r#SV462�,�P��X(��կ9��:�4f�ϋ���=����{_z������4PI�m�}�\�.# �dj�����[��]�|�x�-��F�i3���rcQ��0�@�Bi� e���(>��"�ؔ.u�mP&1ƋTT3u�l��ZS'�v�P�%@^߈6��Z �č�L~6��.$����Y��j�A+��H�	rAH��R�!0�I<��T�0���7qF
/,G�*ǈ1�\����P���u�-N�> k5�=�5��&E$O1!÷2T֊Q@Ǒ3c�*���;�L�m���'|Nn+�ۯe�uok�������P�P��e�;K����g�5�β�\ńlA�򦨄�*�!�	~c�%�<*�'��X�*�&bvf��$���6���I+Q$�,ғcf-�^�K�n%����淜g	do!1Wbe���̤
�K�^���tz%�ה}�B5���������:`%��w���3%p�K9�"�j��Ie2�4bJ֣k�x��Yx���z�_%/�1�@p��KI(��#G,��<�4/�ĳ v��֒^d����8&RE�
~�]@�}�H.\G�;>�X�4.�0F1�ƅֹQ�4�-%�š��x�8�h�:�w!�j}o<δg``7�#��əJ�����9�x�R����r{��q�z�i��̽A�Oq�/2�'4P�8��Hs��
C�B�>���>>5�_3��v'����"��*�����y��S������~�O������?��>��-(}2a/̑�!'CI���O����_������3333/ ��� ��6� � �z�@����PDA 8����z�` ��y�;����`� ���yV�)$�w2�H����J�
1
��B��LR)���%)�(������_�?~�~�k���@  ��64Ѡ��l�a�����z` �8� �=4������}��<t �  �  �׵V`��D���U)@1'R�!�@�*R4!�n��T�B�^�Z���zx��C�<���4��;�zh�@v��� �6����<��h� q�@�;��t<���� 84���z<�����ZK� �+D0M����H�H�94,AM�k,���η��y�΀x:�����64��   zh�a� M zh����6a�l���8�@��y�c 8��;��l`v߫���������� 
9 �(�T2@=H��H��@�+@�H���p�JErQ���

Z
))R�,�r2�w49P4��>_�~�P�X�����}���T�}3�>��>�v��]۹ue��r�E�I/$�wY).�Ԓ��^�rK���]۵)JR���%���Բ�Kr�K�/%何�.^�r\�%�$�,���vI-K��\��Id����$��%�/�.��ܻ�wWwVJK$��I.K�WR�Z���I\��컖�n�RԵ-Y.�fwd�){Y^L�InK�{{%��ݒIr��wd����ܗ�\�佻�v�JR��+�����Y-__�y�_ۘ�K�h������2��ć3ΰ�;[q�Z�f����M�!Y�n�07::���Ԗ�M�	0�)a��l���X&E�P�K�tHk6]� �I������#�(h�[2=����Ngߛg���L�B��CJ�"�Վ��&������Z��UVSWٴ��Q��@��]�HF�Ye�1�%������$�,	GE���3@��2Z��͡�C��|>QR�h3Y`���M2��X4v�,�ͭ�cpb���m�vVWV�@���:;�w�XH9]Z��2��Ŗ�Q�h�@�4'TǮ��ׯ�|�Dڥ6��R������Mee�+M���K�v�m����fZ�`5,n����\�G^^k��*Y���f̸!uF(�����׶�҉��c�]4���Gb�B:S[�&�SUɠ!X��)6�t��]YcB8��y&CWR�)���K�P�DB']c����4ͯ6�@�Ў�F��h�l�6��榗mq�c.I.�se���Y�����^�v�Ի3L�Xm��m��Kc|{��VZ�	H�ems^�<�ϢO{��v���m5Ԋ\)�3H�q.�n��,Y����PxѴպ��aČA����� ˝���m�c�	�M#.���ؗWX��陠�P,�	��tي�୴B��[v�eM��î.�eP��q�"f�#u�}�6vsA��㋳M5��Њb`��\��ˮ�ծ�����8���@��1�9���S:ց��
u�H�r	��fK����iO]En�#�Vn��j��nPN�eJ��4٪3p�#/`��4uo��`Lr�G�]�T����:���ĔGk]p�u]6W. ��3j��CA�ѣK-���դb�2YsM��uܻC���֘[mIbF�JZԚ�4����L�vU�-������xS*|s�8�ZƜ�WP�D7j ��72�Qͽ���������.�b���&���j�q��GBYX��XKV�N�nSJ����Xl�B��P����.J�Fm�Xie��#�)nG],��i�2;l�4��,rGA���[qpۛ2SL�;l�k))P�JӅ]S�{�/z�>�۾"��5J�o���B��2�pK���\�p����AP0j�D8I��M�-��fL۸�C�eTb�RJ��k��mb�X��=����0/��liE
�G7+v2�;��%�n��6ۊ;^	��)���@[8��q�A`�7*F�V4V�K�Ўu���2��]�����y�t-��:�����醌����˰�iHK�mE��ۏ���f�˔�-�{e&�Ge��l�3y�vW1���j[���MEҮ%�A\e�B�`ml;V��I�%�c���]���kX��ch�IM��qY���7�f]I5�B` $2촎+&֩�-.4�A�@�Q9&a�6�!��š�	lݬ{p�43d�JLJ��z��# {�eS*C�eYK�\���`D�n�����3Ƌk���Ε$%Tm[%������,�hٕ���v�J1�",������m`�B��tX���0�L3�Q��N�a�IK	�=[ۂ[|�b[.6Z�Vnp\�H�ɮ8��e��e�MB�Kh1�8t,�Q��L�9�-cj8�Y{ٲ����crhe�2���ects���n��%�� d��1�m�4��6�Z^�͝LAld&Pڽ�t+t �Yn�̷!0¸�K�Km2�&�[M΅�5�.q4��iLk���Bꯋ�1	���6!��4ej�Zf�z�V[[0���e��kD���V;p��L ����ϿW�߯߆���@=@�����W���lx4��{۟_���lx4���{s�~����~�j�њi&�iF�a�0�0��<^!uqE�^� �g$L���R�L`��]&�`Im��V��lr!%�K/x��5���n�٥��q��YiEɕ��
�a����]��j�Zq�r�jjh�YLI�\f�#3��wz��c<�Me!�sF�5�Ų�3*�V/�zh_U}sij�pX$�m�x��,v��\�r٩X���UKYiHG�%i���	�-�n�)C_�6�-z�4�э)�X�!Ts��,��_�%�8��uѷ@,ifq.�J*Z�3T�D�[cf��7YlM.� KK]�+��*]u��GbTR���˱�0�z'�kk�*mlԶ�6[Y��!`�Z�]]q�[��c�0p��nM)[P����*] fbC�����&ҫ�f6��Ql�gl��9(��ss��c��%��S.�`�y�P�t�Uq]fa�`t�w�!
�����X�j������/��X�x����K��]���h��,����T���8y8Z�o�"I�DD(�Xq�8qj�z�����n��L~:p��a�5s�cy�O���!@�:v�\�M��J$�S�Ã���D{�Z�u�w���U h�u[4UknN#�*Ո��h�㉵�U.�tj;��:��"�E�3ƒ|I�0�0��0��㤑ۢ�q3V������᧗��y{p�0LG������N���ڶ�%�߄&87���&u�E��ⱒ�OK"8�G�23����\(�>"_q���\��I~������[hOy�I�:����!��!{D��j���Ƽ���}:�x1�g}ٔˁ�q�b<Y�x�."���Vj��˩uyn��y$�.K��j�c<t�����M�aU�)S��Dc�@V�֫i�^JU
 ���lx�T0�[��è���]�ȉ:J�U�qP��4��$þ��/�"4����+�Lv�A)��&۫]G��l��Pw�� �kW��0nZ:�����p�<�����w���%�%�q�:Cl�G���D����t��-Ip�}c�N( d�$�N�if�0�0��0��㤗uyK��uC*��d�����Q��Aі�F��1&xx4K$#%u�915T����m�mpڪ��-k���/��r-��At�P�AE"K�x��@pF�͌&3�&�
�x��i����m�J,Y��P��A,��<uaj��)$�8�{�q�2;۞"��:���t�82Ot��,��a��Y�OAe���JeKqQO������oC��'����g+��ֈ�Qf�r8j�"6�qPHnA��mR[�`��֭�I$X��{RUA��j*�_8�1��1��:rܲ�%f�V���k�ՂU�[D-���*�$c�vw
@В�)�k�w{kpv�իcʺ�2gMSÕ�f�2�����,u���o����Ǉ ��W��*���ڎ��r�=�ؚ�u�z[y�Pzb�ȡ:1���kg�p���G�3欤Rh��8%��U����[��Q?�ײJWd�_3�ӓn&�5�pTY�%l�e%�T���%t���E����n	�p���(���j܇�y�����ն"���""ӹM�Ԕ��I�	G�
l�����%��Ӡ�Id�$4æafa����x�%ߒ�326&�~�*Q@,^� �)F�O��S$ O0��p�%�t�{n"8��Q��5h��W:u!����|d�9S���;M�Ԟi�^q6��*�m���q��o��$jKlfR]�ʔf��:���yq�X��m��t�w��Q�c�$'Ҕ�3��x�
4�N�a��Y��,,��:H6�	r�M9c�CTbdb=` ."�&�����U�)��h�M����Z5�񂆶�0D0@�x�c,�5�M�������L�����B8���.r`�	�4�Kw���6���pg#��ruuR��Ecl�Ս�ʆ�ah�֠-��`�GC�o���5�b�Ѫ���)C���Ĝ$i�0�0񅅖3�I,���"(�e1�F�/� +�"�ֵ�z�w[Ґ٧OD,-��VTd�jiPuR7�%�#���kޕ▢�D�@�2�1�4�-�&V�+��$g����=k��#��͙��ʚ�D�Q\�$�Z`�����3�Q�A��HW��D�t�G	M4p�j!MV��p �J���FID�$�Fa�0�0񅅖3�I#�YȢ9WfD����،#p'b�i��%аl���W��Ug7.��q�Il�9�u���,>;� F)�{V�Mq<��[7fi1ٚI7G��-�C3�V��ʽ�U�h�or���f	!� �G�r���D����BF.#)&B������L-��K{���Tz��A�v�^���W�qK]J׬|D��ۨ1�I��mq�9�k��P�$�Ax;]��{A��/"c�c���|;�s�t�U��u*��XCh.�Ø2��G���8�D��Y7%k�i��ߖ�A��Xaґ��	|3>�����"#��ov�y����j^��~�~�L�#$�.���oe�B�餜$0Ӧ8hᣆ�`��@fb-T䅑��-� !r�j'�P�uON����_.����3��dp�z��G�Q����*��4�S3���nWEGOh�	�{�8�pۈ��� ��<m�JP��q��׬�!s�����V�Ź�D�)N��O�ߧ��I�~���X�q6�˧8vt��ٺN+�����л2�i�����gG�!��2�I�G�����xi"��#Fi$i���|i8,�oG���-.�tg-��m�ѳa�3Fƴ�H��i�� z3���(�F�#ќ��5�n����4��h� �L �/GK ����Fa�h��0v?p��F�Fi&����4z=��� z3H#F�%I���z=o�h�kL#Fh�iI#����Z>��(d�z<Kq�����h�za>���i||M��x����<#�����|�O��z��_��=`����(zL6@�i�~$���rܷ�È�|(#uc��r^��t��,vi���7��$h�zd?N�G���!���F�H�h��oO���.��:3���{ɏe��=�G��e��D{0��0�h���	��y�<���G��AF�?S)s��a��"4�Ը1��]:�*�$��6UL��I1�LuJ��!h
�D�j_*��az�����N�;n$��u�|[ﰯ�����3��Θ�r�Z��e#���B!+;t'Kwv9����'��N:�m��F��ڠ���y��SrV5�]��7�FG#���f���#��Fd�PP��M����>9�5� _}{�^��s2337wou��L���$
��w��̌�����{�S3�l ������32s33;�������"��w��à<0��������+�,�r����w/��$�%�{.W/���W�V��[��fa���xۏ'��kN�4F���L��l6ri) i(g��f��y�K �h�&A��'y��)No#ˎs'��{ն��,�aec{�9!:y04KԆ�N`�=tz���Md��&���_��Jٗ���f~���M�PJiZI)qa�����I�C�xI'$i��%�N[�Cx�z���U��'䈂 ᇎ1m��Aþ��œ1
���&o�xj�Xk�i�i=�2zc��óx�l����Y\u��}^:��"bhCC	CJ��J�	,��4��e�,�gK0,�H,�"�r�_�u�{x�@ 	{���d�)�z�R\�����5���G�;���2Jv����$� �@~���Sa�i;Ǔ�U���Ywb���'d-�rw�/3<B�. �gq��-1kX��K5A%���!���x�t��(ps������ �I�$x �\��+���XpL@IyX&�5�pa�C�06�r�>�j����"���G�9� �N�7���!�D&��!�xÒ�zy6�?6�$������P�a�b���Ř��l5)�$�a�P��+d�v�$5��`�xeI��Q���L0��,��Y�x�Q~�
�����d�k��7n'ƷW$n�b�r�W��1:L��F�%�E`����:z�m6�oB_w뱾?�����:�����T�%���u��a"���U^-�wcɝC��s�������Yy�S[ا`ژ�g`�}5��ձfwt�0���m�eX��t����sy��P���=���҆�TkҪ�p/�����M	hª1c���0<YN��v����3�@���K���.`k����8A�����)B�8�v��{I|���2�N��=1�HvA�L6`��#�E�(��N�9�#d��Xpi3���t��Hz�b�M��G��`�$��\��Yge��xD�����âNX$8$;!ԏ'O)�tb<��xGF�%�֝�'I.��<���q�iN�<H䗔��`�^]�:TوXbLY�%o��6��Y<�}���D8I�� S�H42&��ه'�ѧA�D �3���Ie|t�,��<aae���)*�K�?&�Wz{HЖN�:��8%���-&/,��dJ��<�̈�t��H��f�Ry���2èb�rI���U�$��P���'�N��.qAh�t���c;�DZ0�O/���U��Ⱥ�c��8zp0�d4C�\!��xxZ)�(��: }���m�<��'n�&�3<B_��X8~NҴZ�j#�vR�q^�p��a�ҡ��%'{8"���C�\p�pƞ0�ʨ�OD<2�K�QN�H��z������S	�\k8�!��MK�(\R0]����2C�K��L�!P�i{ÒG��<t��K4��L0��0��X��P��{�8��/m�t��[����dDA��!����Dg
9M.I��oÕ�l�<0h�}��_d���#�&N1��a��Ȉ�d���7Q�rK����K�A��ף�MYj�(��W��!W	�D
��vpb��K�$�<4'hI4%ϑއ�2:C��4�b��V=��|o��*��1���g��1	���̊4f&>�aa'D|:��0���#7�ļ0�b��
�'����v,݇U$��r�R=8A���$�k����<���"5�B��G7���é�"�B
9Q ơ�E}��:Ṙ���PW���|�P9PRa�����X=����fӥ)E!���]$�[3�6��׃��<I��?æafa�,k���%�>���,n�D����U<��� �KӾ���^��L4G�+�v�7�`�0�����z:(� �N�4���-��{��	4Ū�@�P�EՇ�Gg�L�51X������HRHa$%iF��K�#$�t�s���]��"�8���ۇ|��Gd9��}$����3K�1#�iѠ�Hx!9$���5���hԝ+�d���!�NX"	a�=WZ��ֵ��c�AM��%�o�%�Շlu�a�H�H0��8a�f&�Ѭ]$gn!ٮM.�Cd'2�sMC�)(�,_4>E���iK9^�,��a�A���}'U�41<�$( �Ο|I��4��Y�x����O;;�b����I�+�X�xф�唬K̵<�H2����%L*�:�H�Zo߷�;�͂�ە�,��մM�]f!�	 ��@�^�ec��TR������oUΑ_������Ϗ�-V�t0ڸ1�f$铏��iy;+/���8H��m��}U�P�v�Y���>�w�xz"�n���� � �u|JL] 8�<V�(a�HC"��!@���C8G�}��C!SM'}'$9�A&'�i ��i�;P�o'���S�~<H?��l�"P�<A��E�2}M�%�#!�i��F�ź0���{5&Fr`pJ���Ӊ��90�G��ٻ��ى�FP0����+T��8B@�o��H�l�yU�$'K�N�#�Lbd�Dx��,0��0�k�tm}�$З���jD"�����nZ�����b��W�����b�F��t��L�<HN�8!9��zN�Jp�Pw[�D>uL��J,�+�
82ω4���|t�,�<aae����G�Ph9�8�
�D"��(\\�݂"�!�&�Gɔp�O�H�Xu$nIF��K�r��,i��D�#ȑ������ʚ��R����_����i7+�I��]�C�'��0�q�gO8M@z0���i��EZ4�qORʘ���<��K�PPi{�5z�Q�[�();�t���Ī�#�����x�_E�YX�����kG<zyOw��z� ��D���X�pkI�}�Į.i$��h'�IRj�|���h���(8@1�M\7��}86��z�D�B����PB���Fp�K$�N4�0�XY`��]B\��τ� m0�XġRd�1�I�%��~��"�VB�.�׿U6��xGGI�: �x����V�#g+�X1�I<Q�2��xܗ$H���3�z�����SG����&�i�&%���-y�2%W���aч3!��Q3n�g�\l�J���e��O�KaA��'F��f&��6c�!���X�k����D.I�]�j�Q��5↟T�����R�a�<굤��	9<��<r�̄�:!��+[�p�����0��t�2��ב�u)!hѾ����z0��|tg�#f�,ӆ�4�0�XYc<i��y�!O'�%n�8r��B�ʴQ�]�e�YdBYby�&�'�Ȉ���|Ę�� mZ��i�����C"Q��K�"�
�B�iY=��-ǂM	~���Sʂ��������8����G*���q�x��D�!|=T��($a��h�1���&I�l�La�p�pT#�B�0t_�j�Pa�}>�&9��]�٪LMs�!���I
T�+�dS�$�Ѷ�dWF�4�pA��{.H�pF�6A�Hh���=�k��	8���E��|I	�:���p��GQH~��Vʈ�6�oz=����䒃�$����l���ǷK��y��A�8:�(pl5�|=&���z=,��9.ѳH��&��M#A�<�L0�K!x�:3������m�M�Fƴ�gHѱ�5� z3���QF�h�FQ�Y�p;x����,�M0�L ��Z;�A�����4fF�F�ǣ��ҍ$���4z=�����=FI�
+Fk�q�њY3G���}4���zE7�>�Gg���>��٤xf�i:=�Ƒ���Ӥ@���h�I���4�4x=�HZa�#�Ӥi
���J&��(zL6i$kq���m��f�1��> Ú��x<1�^�ч��.�4x��#��A��=#K#��<4�#F�#G��/H4}4��A��h�� �tk��������O�����Q>��G�	��p�|A�>.�O���o��{7�<m]�P�qȰe�9[A�R��eU>�J�н��fP��YYG��}��ht��UGY��h�
�؎�BJ�%��
^L��T��W/�)]���U��~��vj����_)���S��awA��U8q��3��ƛ�h�O�i�g�FUS�K�ڴ4�u�][/z�T
�d��>��E)z([�g�i�@��4���:��D�Y�7Y�H����"�5[�5c�-�5i����41�kġK�&��r(��y��FIL=�����O�x�]�DUN鏕�ے��������� �B��n�9�����h����ݛ���uc��;f5~���䂚��8�Yb��2~�Vl	I�z��&�YV�K�WZ�K��sE�.�؇Q|46�Rl�Z�.�h��Rlݐ�Ú��/�W�0��.��(ѱ`2��=��+OV�U���1��j2�iŭ��U�k%R���>��P�������ӻ�����}�w̹�s�s�}�����{��e�s����@x4}�{���+��9�9����ѿ����2�er�dY%�Yg4�Y�x���B��u	q�9�N@�����R�-��+@�H�g3Xݩ�Jmm6����=_y� L$a����L�R�Ζ�	S1���h֘��kJu�f�������4�M(��gg��M[pk���k��s����@K.�����.�a��v��f�
֫���,Ȇ(�G��V�γdm7^�eԺ�ȍ`�.��ܑ��!Zk,A��%�ZU�L�s6ٴs�~om�vγC\����ږR�R�b�+�X@O�����Rx��BV�(D��m���˵\6:b����������ڠ�
m��o�ۦ�@�@}��l��Х���ٛR�Ŧ�:c!���6����16ƀ�Z���ts�l3�R��2hOy����3���*l�dc����Ƭ ����̧��1�4%�/��t�'׺�8��˿S_�v���I�0�w*܆�b���E}��<o4w��Af"�-�:[��:���G	���3�R�'��$�/���72/�S����;j�J��w=F&��"<�S�Wf68\My�$�����\PP��D)>��C���ӫLzg�F�tӤ���I(�O!�&��1�aC�0�"�����8�p������7�

#�������-�Y5.f�D�\� 2�i�J%4q8�@���$�D�:����$�ӳ;83yq0�O��$>��\�HR��/��s��Q�U��	ӀD�������p�9����ӄ��%uB�Y��cC���K}��.}�Y�yS�6�6�c/ؼ_�\MX�_�<�x�m�
<B(d���O�J�
F0�`��hiE��d(i61��$��J0�8||t�,�<aae���R�c�6�1���ݖYe�A�'I��DK�N�(�(��(<�J�(�PC/G��G��%1RM��q1 鸆���&�z������$K�����	HD�tF�11!��%Xa�y���X��'��p��H�La�\�Ӄrp�m�F�0��0x �`����� �}�%і�aDR!��)�������e�"
#4v02G�wi;X2X��OI	d3ھ8[8���L��iA
&�a;R���cLE$b����1O�(���pq5��[臢XbH<���E�`��{�BNA���% >IQ��|p�㦘afa�,g��;��K����H��,���H V��1�I�%�
 lk�z#8LL�N's����N���W�!Ӹ��O$h�}8�	�H��v.y���9I��,$�r�b���q�Tr��!��1̔R�J��a���T�f�y�K�k��t���s~}p9�o'<s�l��G�c%�)8���8�䒈Ӊ�aJz4�8@�$#�mv����X0�������:b�}�ב��CPR<L�6���-p�<A��A��K8H���%��%��uL(�43��B�&#�䪟7PQ�q�%,%�>$%R�AB($ђtҏi�>:i�a�0���x��g���� ��ST���c�1&��CG��(�G	9:Ӳ�Ӥ�҃���e c!@Q0�����8qI!�<J��AGQ���pa��:$R�A�c�+-N �� �L,#�r2qѧF��M2����5$�	�;9���h��A�q�3$��F<�k��5<���&f���ւ�>����}���ĄAȐvk��/p���IS�2aB��69P�0�=�!�ʨ��a���D�:������L#	��n�F����;HW�!�qu��p�3��<q�l��m�p��f��
�ه1G��rTW\)q0�֌�QєQ�(����M4��0��X�4[WG;��ꫬU ��ͪ��i�y!�j����]�8	��7y$��<��j���ܙ�,��Yl����~#EQE@@��w��]^ҍ��c�gQ�i���Ǖ1W���;1���d��^�zK�8t��9;�U�Sje>Ȥ��q�ɻ��:,*��uT;z�o�^��g�d䊈��5V/�_������p�\SrKj pI*��� vP�ە�C)87y�D�8��( è����S
>y!�"V4�ƚ��!���N�M'DU!��Gri0��Np���I��&Py�R������0�r�b8;���������z�C�qNA��yc�Ƚ�dѫ��A�@�a��S�Ii'�trkG�xbGi�A��5�A�bjD0�	5�T&�-D笄p��Y�7e|$�YDHJF��Se����n�5/�-i�t�L�(��."P��#ʑ���!1�F*c $ep�@4����\��ۖ&~]Aѫ <`Μ0�
,Ç��M4��0��X�4W�Đ��D�㋫,��,�O$�ď�t�to�c9���"�$��G)������0�S4�Oy���!Bx�y�	~X%�����p��%>=��A-b1YA(%4b����	�i�F"	-J(dڅD���t�8� Ω
�ʽjQ,(vêp,�J+�1v�'����ã9vsᷓim9#i���P��7�DUO�>�`��G*i�Օf��A�/?%0A�A9
Fti@���t�U��d�t`��r�h:e�A�=80��ɒ4P�����t ��t����6����^��Y[�x6ɶC�=�vF<�d����(�E�||p��馘Y�x������T8|�8�� �mUF�n��1�4$����7��Ihg�%R�S��9�+����'	5�vFI��XQ�����z۽-8jp��h�4a���9!䃮�qp$6��x�G��])A'H!���"�(a�"E)�
��! ��-H�I��#�
�h$�1Z���41�0A��d1 �\N�Sf/��l�2pFI�A��u�,�l���%��I�Ę�04�1t��L��H��1�m�q��hnd�W��LJ!+�q�M�̡��&�^�y$�IC0a���@��#�%����C
ch��i���!I�!��x��Qf4�馘Y�x����B���c����0c-�����o'Yj�,�� ��C�M$GF<bd&0<I!Ӥ��ɮۤ9 �=��	=��K[�:�gE��-��9����}��8ra�I�g��������$�����@Ό�Ө�R�!VP�g,���M��t��:B�t�Gm�-0�w����<�:N�(箊�hh�V�q	#����ms����ҹi%��!Ϛ�ɦLtC�@A���';LL�{/i��-&&J����Z(���UD��ἤV#g����0� ����z:�	�m%)�`�(�E�a�>:i�a�0���x��������YH�h�/
��a�2���	�quj��NfK��8�"��&͎�R�*��>�1�I��=�3Oά�J�0V��L��),g����N�[�")c���5�9�}���$V�aPC�x�D�Uwbt�%hӫx\gr��>�Y������� q4
��#�E#�%4Je�8H9 ���'��՜=��ͱ;�z�+��up�8
R����� ��J'��FI������8����N-�'�gZ{#i�p���4x7�lT��*���#��Ѣ� %�(CG:@KE�G���q�G�'.yMN�=Ϸ+,��{�_D�A��b�G}��Æ��q�r��ba΃	d�Y�]q�cI&����0�b�~�Y�����t������s�ñ��c�҈D2Ƶ0��L�5�dpА���/:]5A�0�$�D/"ϾM���K�E����Q⎔Y�>:i�a�0���x�r��(`;8͐U���e�W;/�8�"!0���t�:�aE!J���qB�u
���j���M}��W�STO9~KL�>\��#�D����?">�C��������e&�G'/	�=��l��<N�zM��h��<�<�QhgZ{m��胢���$�tGr y�~n&
��L���C#㨤��jQ=8R�	`5��j��5H��f�N���L!���)��:!/#��Ԡ��2N� c�R��a�I�M<�D�s��,��.p������Hg�h��zl�#G���4�zp���F�M'G��h�2�-��za�pt�:3���׼�����e�'�Cѱ�YFH�e�iD*4��8=Z84f��4g��,����0�L:I����<�h��4�a%�ãL&��H�H�zt�����{���F@�f�p�"h�f�E�[xi���kG��Npz=G��PݎG��n(�(�4f�G��N����i=&���ΚN�G���zp�2<ޑ���)� ���[�GC�HZL6�[�� Ѷ��f��tlf��Sl���f�h�>�G�χc�k[���G�g���L?���`ύ0����8L��>>�&�����4f�F��z=0�Ot�(���oHc4��}�{(��G�}��E�I,$I��G�}�>���O��+����b~�f�����R����34f��P��m�(S��Sy�Jd���N�ݿL�Ҹ�ȷg�VQ�9C�_cJQs�q4�8�O$#�N�w�(��o�k�fq�b:�Ȥ)��Z���C���8ٮts_�{-*�b�+K��1�I�1[}*-]x/6�b����P���c����%�Q�;6~���^���ffeffg323+�Um[�9�y�}���v7�}����9�9��`�:ow���9�s�s����ʭ�l�adAe�QeY�M:i�a�0���x�T�D����\���q�)����G��u9�����q�WX3�E�W �b�w
DsϬj���5��(����B;K8��i�O
�" �(��)p`����F@�e���T#���>#���х�>5�|dHS����r�d��U&�4�0?߳�2�VJM�upw�B>:�%"��WF\h�Ӈ��d���u��vba ��=��&I��r��U�$��b�c�=�%t�ê�0�-�=ڙ���� �%s����uin_�e��(�R&0�v�T�ux�����V�P2	 ��(��M:|i�M4�0񅅖3Ƅ�r��J��2�T�� �K=�4�:/V}s'��ER�qvQ	H�����h��G�i41��[�ח�m�@{m\�O-��u*G�R�h�b��'C���N�9q<�99tt�w�,�+�:�ixf.��2YD�P�����7���tp"<&qֵu���4=l�Ӄ:�����dg��7��������������4��",������#���%&#��]���Ѳ��d��c�I`���2�N'�1;G�CT�����$Rݢ	$���iG���i�M4�0񅅖3ƇV�U��Ҩ�4���?6"�&c8֤�t�XT�����uT�y'_d���vV�!���	W!������8О(��6�m6�4.^蜰���,���&H�%�rM��34���8�9�>�ڹ���cL�»;*�5Q��;/�z��C�j�Q�"����e^�a�u���(��D��r�'��N+9�r��!֌_e�"ǉ�\@�2Q|HP��j�Fz�w�uQ��F���:2��<r�Đy4{�R���P�4W�#4n�H��1~���J ���.�^[��n�
��"JOo08�z�dDScg�t�����UV;&ӓI�b�8#��h�h����/'p�m��1r�C\�i2�i�#E��F( -��p������|ػ$ ��#�l~G
DW"^j�_A���X�B#Åk�,P����((�H(���0�L><i��i�0���W˝Eo0�4`����K��xfa���c&�q|�;d�XPl� ��c��a�B:R��\ϗ�"�nK�8���K�D�Tp�q|���%P����H�h�E	1���<�s܁�Y�Y���`xe��K~���X��|t�蹑ĕE8�!���C�A�|m����"�����b9�I,�=/J�^7�8�Aj��N�|����:h׋!<�a$t��4��O��i�i��`�|�ىQ�*�8�	 �	B g;�=�bd�wP�KZ8$�3��P�qyj9��d����d��ֆAJ����OF�騄@tgQ�)��)	O�ќ��9N&H�}��!�7ӈ5A����:4P@����=S����k�]@�I]!i>#na>&����^o2;��r"x����G��a�P1��T|�u�߻�uTn�,����%	������Oi��<_�'�e)��pܒƼ�o��ќ	4�:Q��i�ƞ4�L4�XYc<i�b�.���.#[q��}��#i�:�A0�N�Dp�nwQ��-���u(�����&�`�4�Qu�m���+ƖlA�<*P�i+��,�8����P̶6�x�<�x�k`�%A�D�-�������������4�L��7�@!	��h����c(�@龢�0�������<L��oQ�a���C><�y4�p�0h�J	>$��t�M8x���a��x�����=\[��<�8���L�. M��M�)WV�����1GȐFHF�-�#��ո��X}�@��~9A��U{Ԧ}3-��݃����i��qn/V�Z�j��'��r�X:v�y3h:�ꚺ ��5E�j
�uy��U����v����M�uN�Q�B:�$�S���P��c��T�4��n�"W��+���%G
��S�&t<3D�k!�/#�Q����97$�KM���>��Rt:3�g}*��!�"TQ �g��H�$P3E�ȴQҫ�q\)"TZ^\Q� �I@�W��`#�W.�P�R���Ua�Vź%�I)�<ח�(`�A��:Hט4p����{F�n�<PA�8Qe(��i�M4�M4񅅖3Ɩ^r;�S����9�`�)
"[t�sؒ	 �	/��|�˛��O��B�-T:�������:��G%���I*���UDC��s�9ȨL�W����g��eoȥ'N��"��_ʹ6r��3�j�2/��*>K�J0%.�`�By��(��"EP)J���$�DY��|�@becx3<�E�z�j�w�|b<rO�|�82�զXI����0��t�
0�ώ><i��i��4���`�8F��8g׮]�}�;��:���,�}?Z4�h��z})���\#�7�>�3�)8	��=<d�13�<��ζ��h�[Xz��G�x굫�����T̓ݗQUY��[��핛�Bu�G'��*D���)3h�����:�t�pd����f6�ѽFk�� ��|�_,�4���+.8i�5^!z\0�fh��A�c$O����qDya�T��pV�R����/��:HQ��(�(�(����x�<i��i��<<3��z��Nffpg͙�f� m�޴�M����u@�?����� �GJa��"T����u��$I\H	�����$�>������t���}AэM!8>��#�B�2�y���g�0�ŽGBFuE?������C��`X#'�e|Ci�&�r&f�p����I���0@x�
]D�|Q~Pp gȕt_�s?d���yX�e�|�&��n-|1u#�|iB��3��CeF�f���v\i:=�F�ȡ���zA��8F�G����xiM��������;�f�56֍��f��ѱ�3�����o�*���83Fi����g� ,����a
� �����<4���`�zaa?�h=4���#I$��A���z6=�h�t>F���z5�cјi3��>��i����B�������H����4�N��#G��n4�o����h�4�,�ǡ���(�
<A&�#ќ(�(�a��!2�Ѷ����h��m����֏���a���֚i+����P������G�����c�zA��?�����x�[�x|B�a�,�|�u�#�89�Z���M�F�h5�cѱ��
#Dh���FD�\g~���!Z{�QK�n�k�⪶��@��Ws���]����G�v���e�d��jbͻ���J�nN��sf�"�i�ʉ�U*�9�WՐR�)�����������-b��}xti�/~�m�KlL�4��r��[Z$V�N����,��%ʧJś�ݭ��阍:�4WP�����nȔ��Z�e��Z�����ܺݹ˨i�z�Rt� ���Ĳ+��mK�&I2�m���[o�u8>N	)ֶ���#��@�p�5u�8��"���2�+�\��2��ꫭ�����<���x���մ���795��#e����
�+%�v�We�B�Q�"8�0`��Y�*z@�v5n�a5��{���ó�\���m�kft([\T����im��x�K��@��	֢�nЃ�-sz:���u�q��rX�η���}���k����a�{����9�s��}�����w����9�{Ͼ��`�����\�9�s�}�@vffUUo6-�,��QeQe�4�4�4�ǃǆt�$�Q�%I.���� $��k�ՙX�A/M�7U���*���(�fոٔ�Ĝ���:��+.�f�٩-�y`Ђ1vnִ�i�)uړQ΂��X�f��ܮ��l�5l6���[v՘�ãFʹaB�qH�,��R:��X�-1^�fJ�,�me�u:�ψom�-�׭X�R;HZh]�^R4�Fˊ��GKq��bH�*�T��D�Z�����kbMCkHQ5�ͪ�S���m��v�`��c�z�(b�Ƭ�ĥ�|���7��/�W7:��ݶ���J��7m���\9Z׭��f�W���3�lU(һR�1΍�h�m]�[�v���p�cy�Kf#kk�gX5����VMV���L3cXܰ���j���V�i��x�����[}�LÒ/��1�H5/C��{�m��ݓ�gKr+�fu7��zl�A��Ƭ7t��v������zt�찍���*�Ƨ���B�7�ങ�ޣJ��H��#�v����J"~n$��[a������g��q8�h$f�Qqz�(�������]���:��613&#���؎��0l�>0 a2����{��cc���_)�7Ҽ�)@P�Gp��qB�"�3}u1�C֡�g�C��3Q-����!}��ʈ`C�"�\5Y�F�P�J� �g�0�
>,ᇏ�i�i��WP��_{Ϡ�R8�J� ��5�cm�I�V��I��1�?�/vO"� $e*]:����N��pR����c� l�Y��;�s�B�
h�O�H����۴��i��[����eu=%u.����$!:|��/,"��BN�^͒m�r�9�kgT� ^� ]G2�k�YF�!�0$�5�|D��I�3�d g�|oM Gt�Y�βBҏaE�p��4�>X�{2<"�-�)�B�����M�I���ID!$�L\�9���/����*[���)�,�Ҹp�F�
�FRZ������>��_3��%�
�O�X 9%3Aʂ(��j��*�u4���Tu{j2۵��vӐ��|V��<�I�����ѐ�#�]�W�
�4b-��#E���D.~�6G
(�殮��)�y�s�(��4�z^��s��Č�'
$�����FYF�p��Ǎ4�4�ǃǆt�X�34K ���"�"!3i����N�;�㈃�Ǝ��82>���XΥ�nj��q_�u}֗����@�%�e���LfT._G�9-G5D�8Z�c>���I�FZ(��O#���jGHժ�2D�3_̈� (��F:�F=����	8O.�r;�p�Y�&3O�+�Ʊ֩�]LϑB�Ym�<up#8>�t�>P}�`�X�g��Ď�xeaGJ>>8|x��a��x�x�"��?/ce(X�WA.�DT�RʐʷH#B������*CMK�5]X��;cSjȳ���.��b�A$^�Ԉ������_gtsy���V�:��Һkλ�N�a�c�wp�5o��T��Uh������<��� �e�e�Ӡ�}����;��y���]�y�Z�yZ�t%K�J�9s��Uݶ�~�3��>>�C<���PYl�Rb���#�<������% gK\����֡a&���9Ͼ��yN6�dr]�}`f���rd<^�h���AJҠ�B� gJ_j��}��L�tdD#��JIT�	����\��a����(G�-�8���(<����r�D�<�cM�����Dq͹;����&!"y�%](��`�D#��LagaG
4���x��a��x�0`"���CE��A��p�� �M���m6�oB�(�x��w*������z!�E��[n�ɜ��q�)Cή��<w��6�����{�$���y��X�xf�Q�"
����:��s�HZ��I�~�g�|U�"|ڤ�:���w�VY���G��B ���ɬӇF1���5.N��84�PpgnQ���q�J�['Q���0��,Ӧ�><i��i��<<3�wД6�r�l�ι��A@��m��m�h_��b@�UQ��Q�}W�})y�!:����~���E&3&�'�?���&x���.�tLgQ�*V����p�p^!I�^ڮ["*9� m�Me�aґZ�ʂFb^GQ��*�x�*�g�T� ��#��>
�>E�װm����qw�UI���LM��� �"�"��ќ�����P�{,���+�Ĝ0���t}><i��i�<<3�U\��fj�"I�o�@ ��BOt��O���1�8<�������ه�.T|�J���ب<4{V�	�n�-/15��=^�V�_�� Bh6DGBNȧ�Og{; �-M�}���#��1����~]S>=����@1��[>D{�����W�1��2�{N�<3�B�σ���!��Dt�32q���ac%��3�^UC�\J��p��>0���ƚi��a����:X����gҙCUDh������6蒹p1u۵b�˩kŨ[M�[�]����Iq����_� �	/y+�!������+)�+�{��{:��)x���{��r���4�vp������q��[������%��K�:__d>�F�T/�f�*ljT�FӬ�襮����Q[��u��]t%�D�;(ei�oV8;r�p�l�(���b��1�"`A�k�TI�<՞����G�p2�D��v
��������	:��#�J�d#���ߨ�Q9T�j�lv+m/3������Z�A�Ppf#�IF���!�_30�#���"y���t��E��OyK(�3�/W�D#�>q����h����{�;%���'˫��^!"FT�#�c���ڎxM=�P9�����I�J>4�ƞ<i��i�<xg�:*���6���9�=�'�Q�2	 .S�}��"�"!3�%��JR�$�p6B�Z���KP�_	~1�����4���_���-��؈�2���f��f2�|��*C�С�XϞO|�<���â��Fda�Q��9�*b�&*"b*E-��g�M��X1�J���e4�������@B��:qt83��O�5�Aϐ���>,�g�$���0����K۩Id�ܒ�K�K�{/o%ݻW��u)JR��%��Y�r�[��K�y/e�.K��K��.Ir\�����]I/?,]��r�vIu.�ܖ����]�n]Kr�Ԯ��%�R[�K�/n�%�KrK�.K˒\��������vj]KV�Ռ��\�W��)IjKr�^�r^\�-�u!��0�K(��Fi��i�0�L>����}yw}wn��)[��)\0Ђi������&����{�MJn�W�����`�(��Zi�9�7�][�� 4��q�l��d�5ልTуWo1�5���Ă�z���
��i!��QL�}D�lj��{ol���vJݱŎEMꡮ�gh7�1������X�tj��a��U[~D݌�S��(�oz�E������C�^J����pU�r��C�R#j����]��ӻ����w���s��=�� �t�{��g9�s��}����{���9�s�����7��}���\�嫗.��[��Ox�a��x�� �����y�AD��V"V#���u,9X�!j0T2�\�.�T���4~��&CFd3`�1�k�BF|�'΅"O��]8��}�5�)��
�i��������.b��@�]GnN�W���ʁ��Լf�BT��#�T2a��A�ϔ�k�IK���`�4�3�,��8yYz��B�lա��!I��4I(�p$��Q�&�(����Oi�i������B�S�S�!�D�CM>o|����3�i �@:���*%~MCb���0�g���f"WiZ9��pg>�L�25�~�)b+�1q|�.)E��Z�F�J)pZ�����gC�%�#�{���8x d�wj�y^,
�ۘ�Ǧ�X���n��x�\�b<�Z����]��ּ2)��g:��F'ȳ�4|t��q}�]#ˀ�Dt��J<a����4�L4�0���خh��G#�'.���5��V�9�x�#C�\�#Bi��ܕt�t�!*Kkc$Sp���Zm��m�h[��}(_�]����q]J�(��7zl�u^aӥ���G�V'.���!on�moZ��ڛ3uEqZ�O��G�|M]�.q���CԊ�ֹ&w+[|���W8���� n����g��?��T�>'��l�N�߽�$�I�ײ,۩$,1Y��|�@Xȑ���G�b����.!��!(8��{�&I����J4f��
��F3���qOiI\���>#F�G�L(�Q�޻���p�n�A	a�B(��!}D�ܧs�U/�AR��۾���tw���I��am0��\�hͬr2�(�&�(�>:x�M0�L<yu��.�q#� g�Ɉ,yaQ�pDAD"��Pe��!�>k��E�VqAa��&B0��8�)G8����&a��Gj��U'Q��L��`�J�F�$�>�tL���"%x��f�E��(E��p�'~l3}�2�Dz�dÏ��RƇ��w�P�A8�������0]X��F��1�_��""�w(c�j�@�D"� �G|=.�bh�f�mVJ4���iYҋ0����ƚi��a�ǆx������1SH(cB�|�E�q�xM�%��� �t&��_���ǹU�Oqk���a9���[�A�G�G���V�W!���((���~Xn�H_���L:Jj�UUS.�j�|buj��!������	�dB9��~\!)<q.�G��BgLIa�N|�m�.����m�� �(����:W����C�/~VB;r���j>D��p��4��M4�M0���<A�Ɲ.Ix;��l�N���>��Џ����$���u�yiJ�Z�Q�9h�䁱��:b��z�,�*��
��%���c���qGxO~����\ۥz��ݙ�]�sۊ�CGH5K>EZ�f��:��0^/־8���X��GB
=�r�D/�'�����"G�F-�=0�1�$�F���c4���H�o4 ���/a���K�A$��I�N�0��Ǎ<i�i��xg��ܺ˵^P�H��-�ʰ̡m��GqT�)5oe��4r�Jb�uGl����,M��4KKe"����v�	 �	/,U����u��P�O��T£j��Q0�f�ڝ˪d�E��n�eQ20F����Vs�D��P�)2-�ZJ�"�4�UIŢ�+#x0�V6MҬ��l�3��#��H1Q���%����q_1� 83 ����D�PKc(�H�<�u|�|B0� �ьgS=T%q��³2v{NM�v�4ۻ��LG!�ppA��D�We��ȵH�v�{��v�N�F�Fc�pթj�}�rG�#u�/q�ц8Yj�B5z�qCG�a$��SgY������Q���iC4��t���0�<i�i��xg�:{-=��|�ӵ�~~� �t$��&�	<81�:�|=�����J>n�l�T�Q������Q�6�ĝ8�ϱ�"GѨ|�CQk㈤����%43&̈#��1��/��'Q�$pR-�J3�ߗ�G˹��T��. o �����AEi�����I
d�l�B8�6��$��
^�p8�8���(Y�x��e�tJ���队���Q>�H�����I�'O�0���M,Ӈ���F�`B¨�uiʕD��[0MĂH$�K��
]�0�m� ������1j-�83��t��R8�iG�<�R�ad%�p��g���j�J�߾B��)r�~���:Qڵ~F(�3?|�\��#Ikǀh���f�����۴���hO*ooxӤ���p�G�+����Efa�;O|��2s�ʸ=����9j�*< ei�N�t��4��0�L,��x��v&7��U�d�a�@���'��"�W>�i��i���>���cc�w'��o�d�b(�0;�,M��=3!�G��Q����%��bl#`Z*�fƶ�y�wa����Uqw�Z��R����aGQ�m���p$���ņ�<���m�Y�����.���ð}%��|�Q.�����5���%���b8y)>C�zqOTL�%���x�â���j5uA�4���4��	��I�Ir^ڔ�I-�/$�$���;�wR��R��JR�rթKr�[��K�y/e�{/d�.K/e�$�r�^�ڒ�%�$�����)ud�R[��\��$�w%�u-�wR��31u�%ܒ\�/n�%�KrK�.I/$���[��n�]KR�ݦg�.Y+�ꔒԖ�佒^ܮ�r�0�a�4њi�i�M0�0�ƛ��Ӥ�hhhQ������@#�G���6�u*��b�4���A��+6��Z%!�⿌`�:H�r��qQ�ղe�UY5A�zڛ�����W�.��
�s�*]ʤ8�u���\擙������Qu���i���=��2�&�j�\�5ײ�օ���Ǝh2��*V�41N0�ڵB�4s��[;�@��jC�CfU"��/W]ܾr�R=�2�UW�tN�<�N���`����T����^ɔ�c졲gvT������ӄ)Qa��
w�u1�(R��}LJ�UM�=��U�wYՖ��	�Z��٫+�ѓ�Bov��4A�X$�0i�*�uS�n��/1v�
��D$���\啤�
��*��y=V:�7pd�����M4@Q>��=�7�Y���_���ცJ�5Z�j@`}$ea7��0L��ua�ң�����7���6���њX�Лv���[i*�X��+`�I�i��Rb�Ikd��eҷ*
��.KF�ܼ������t�{��g9�s���� =4�{���9�s�}�������s��9�>�M{����U�,�j�ˢ�,�f�4�4�M0����3��5z�-L���s��[�{G-�R�kB��X��	M� �.me�k-����*��e����Ui+�1��`�VJ��tir�5��ͦe��7-�MɊ	ZK�:�]2�xƵ-�	�`��ݣsj�n��@���tPpU�U�(�!m�ۖ��M�V���ZT"�!),���ȸ�܎N�W]-���R�Y��\��.�Vj݆-Hm4`UƍT3�l�l[Z�l��]B�`��E��i�[k^
ӄ�kA���Yl�Ӷ!n�,n	���1��

+CY`�e�K���;M��;�Cfk`X��e�f4�kic��̳�~� �t'Ԉ����)!�ye}��xjl�̓r�V8^��<�E��.<]�n�b3m���z�*ǻK�ʾ��@���wVgzoq�4�
M0�t|����!�i�� V~a���,'��D%HAaN&���ɘ}n(�|*%���n�;�n�×RU�K^g�I ������E�Q$�9��JE�����m/#G5����ג��E/�}��Gެj��y�v���k+j��Z��4]�TG&���&��IF�b�&>Kˡ�Y=G����
���0��$�%�4���ޞ4�M0�e��B�|�|���E���$Z� XJj����6�m6�4#?5�˛�\:rN1��>�W����#��?�x�X�)��4q�4|�����PB:B8�+�m7����Gy�2�Y�\`�&����"Ŝ���B:�<Pt�ϲ`MU=��&e*T�r�_QGOK�o����"P����6�a�C�!�҂W����ޏUy���%Q��p��AFaǉ,�a��K4�i��,g�3-�}��$�H$��������$���\M�G��e.��q�%a�N�N3Q���;ci���6���,>_Uu*�*nWFEB���~KUߏ��&7_W�� 9s�������D���TCi D���񐼼 8R��Q	�A'

(�Z�<y!�l��b1w[�ŨË�"):J-Ye�,��A�I<Ig�4��x�4�Ŗ3�Q-S���_]�u���Bb�f��m�����	 ��CA�q���q�,�#�^�H2L��yB�Æ���҃���vK�鬱E]q��~z���E��^~N:U�Q�@���eCF�m�| 5�&�.��h��(��Defd��6`�>l�<<yOOFӔ�J����cl�s�Z*NH��S�%`3��ʂ9T��Q�eqA�Ə:��4����D8�p�Z����:b�B㕶P�x�O�<af>4�M<a��x��YC q�����r@|��ۧ�� ��*�.ս�r\���Ȥ�n�l�A
'�-"K\�,i����|���}�I���ef���^�Kw6V��g�!|o��4��fvu*g�uww_�;��1��/PfQC�2d��q�����Yl�de���o�=�������������B�� �r�t{�9�ӷ�hl����)����c�u
>G�����w%�f�
��,򰡍�]9c� �az9^Xp^>X�::���s��1�'�}F���)p���q�1s�����I�6�/��쉷Bj�PD}ѶˈӤ:1�>J�Z�p#:A�I0��,�ƚY��0�L<Y���-mI�!��AL���DA�Q(��H��":A�gi�XXI��t���Bh�*��<���+N�#����s;����y���D	�����_>����� �5�S���A���4ub>�l�>XR:��$�Ө�ux҅go"�\�S'_���6�v��mʣ#�X����}#;J��v	�D�P݋�!���#M�<�-1�@�!B$lsӄqt$��x����af>4�M<a��`Ѡ�X������7�)[���U�����M����z��"h�W��yAA'W������:yW^��|t��j�t��K�ׁ�C(��ڎg��.x./8����Z�j�oSw�b���@jxv���	��ç�H��:>�szDATak������a��/��faJa�Sgz"P�\]Fd^d}��Ż]u��7&�WKm�q|�y�>��\C_Y��U���QaD���t�Ɩ|x�K4�4�X� ���%��-����M��M�MTby�����������3�,$��e�����/N'UK��߁�&FI���c���Z�^U\��&�p�ǔ��C	< ���"""���Q'[��(�Ȓh(�S�'z���:�>w�7·�T1��ݙ��u5��6IDp��Ç*4 �"�(!.4|���l�AK��
:8���q+G�	�I�O�,��Ɩi�i�,��AӚ�r27�(�n��4�E�vNT1u�c�P�%t��S_�]W��ic��iQ@����A$^w����R]��U<C�u;�~W�N�1��o.�cU�K�DY��{j��8�aA�cbT��*)Wy��Q�N��fe�s��}�8!;�ٮ�Ll�S�Ҟtȃ�U12UM8Y��$�O�m����">�DȎ"U"��8�x$��x���#�p�|X�%[��A3�����Æ"`x�A}��5�}�>��N*G��uq��oB�V*�gW�6�H�Q��X��º��Z<>6�}D�Lԛ�	ǑG�Q*g�K���9�::{��tQ�A�8L��Zl����D�0�Ėif�>4�M0�M0�e������d�HK�O��2�u��o{�i��i�����EDJXA��ÉXt����� \g�_Ba�c����Iӊ�%�<U����OGG!�R4P����E=G��<h��XYO�fd�Ϫ���w��Jg�'ߝ�B2D�M�Gܧ~&F��Fx���E��}A����@�#�	Ҧ�`q�����@R�����'����x�|�G(l~FI�Y(Å���vI-�$�/mJK$�䗒\�K۹w.�JVJR��.�Z�.���eԗr^��g��\�%�r\�%��rIyr�^�ڒ�%�$���꽔�-K�.�.Z��]K�n[�廩ud�I-�w.K:�^ڔ�I-�/$�.3<�r�-�3:Y�uKVK����J�JIjKr�^^�-�pd�aE�Y�a�4њi�i�M4�0��8a�M$���ӣ44448h3Fi�[��=u]w_,}����(�������dix'tq�D�O�]�mu4>nۉ����<J�c�0�X���h9��t��<+���Ma��G���w�@j�����q��9������o�Y��Õ���9�Um"K#�:�U��N���-�������bP��#�q��$geBІ�˥����]g�}��������s��9���{����9�s��� ���{}r�9�s�|�`7��o�ܹe�\��%�Ye�x�K4�4�X�#�� o�q��m��)���0������6Z:5G�;�8i�XR��5�&�F?���"x�x�m�ꅅ��\�術�B�淰�D��K��`n���l*t�Wȕ��G�g>�[m��١ߛO��s�xq�|�<��خՑ����(~TB.�!�?WH���ID�E��x�5a�^VF`��q�.���S�o�<]4��>/������2�Q�	<I��a��K4�,�X�#��ΰ���n:ޟw�;�Td	䎀Ejh+���Zm��m�1{�y�(F����HVp�6z�驛�v6sy���"=�v��kN�E��:6�-�u�yIá]^3�8�#��G~��� ��Ahƾ���SP1h�Ρ�:p�[n�|��v��n"	�B ��cG]oQ�PH���(Fa�ԫ>�ξ3�%ӥ"��B�!D��o��If�a��K4�,�X�#͙�l�=L؟�yXu���h��\5�y�@><���R`[e�e�5XEР��-�I���֑�l�uq���^�>����=~g�0�cW�����̈����I�2�v�"�� c�ͣq��䋎���*���&�����qmVr��.�����j�Z�j>J5��G����m�5Z�x #���"�dt�C$�9��U!�$�߇�<8A���rbg����Ѳ>�T�e��i�B(�ew�)p��q�����.�VY�Œy���;�;�PLIu��U,6�rP��G��|8g�xha������k�3�k~$�O��0��i��i��,e���q���<p'HK���:��Z��b5}�̈�"�C��"&*`x�Eu�R,���cd�/R�󸈈��q:�\�IQC$>G��`x�lrR �uQW�+��I�v��R>�{ȵE�W3{�\YQ�R�c�֤�(�C�B����������S����B��1���D�\EP��#˄��qb�U�c>�*06M�i��т�T�Q,�7��I�0�K4�<i��,e������&8�Co;��m6�o�^{ 7+����LW�����+��}6\^���6�����m���!��&�(��|B!b�
��=>���7F9t��T����H��$��^����^��\�߉8��s�.3F,~P}���zV�����&	��Q�_6�х�ƶ���$�8��
%�c^cB�/����Ǐ#���8G�M$�M:a��i�x�X�#���bbxɩ�M�6�����m��#*��qnL>�`�[5IB�l�-K]G�����N�^MG9���8�S&�J��_�g�����éy�j����XW�E��{���� t�s�2��eV�G�(�8�2�S4�D�m�×�MW��l4��>m�yZ>e�����#S(Z�y|HYM��Q��#��y�*��\:@Α����O|t��K4�<i��,e����i��A�f���� �mRQ��&p��tti�3)t���c���rp"�A�lc�-��(U[�H˒�l�����H$�K�ǝh��J��y4|�n��RBs}�r=��	8I����pР����ݲ��"��a/u�d��l���'\C�uK���}�n=������5ϼ��_0�Q%��re����RG��>����q��uv��>�H��4�)�7�8�a:~ֻ�ܫ/��pρ�G4:��ě�y��G�����.�(�hsQg.s��q����+)In#14��.��GY��PX3��y;�'W���n�0��t�M,�L4�-x��}}[m�}�84��4�N ��Z!ղ��Qi��T�ӡ�=�}Tz;�Q��\=:��3��(�U�ÁB*��"����0;M�壘��N����߷��x�`b5o��g����#�DSI7ژ�ğ�/�C�q���0�Ka��4x�R�O��mJ�gO��N��%W,�G�C��7d�$���Y��i�L<Yc,�7V4���ٗ��۴��Jޒ���{�DAD#��DB�A�Q��>D8�!p�����h�6��XuB,�K��I���x)I�;�t+��ɺ�����"���ėqQ�4HR.S8��UdD2�x8`�R��S����uE-�'���j�O]>�x{�����9<�#�5_L̸���,�Q�.%�&�@�lf�T�./�H�"Ǥ�(��N�i��i��4�Ŗ2��ṍq4뼭��S6�:N��H$�K�?��$�2jϩt���"��a�`8�fc�#D�� ��
BE��}q�:<M|�u���x�F��0t����4(!r�kmAеս
VW��HGύL�ܽ��6�6��/0l@3וډr�bY1-�|��)r�C����(z�����k�0�,i�y$�:��ÅP�> fA�2I.^Z��I-�%�$��r�]�Z��jR��e-^ڗWR[�R]�y{/e�w��{%�r\������콻�$�%�$�^���]X�]I.佒��K�y-�r��wV�%�I�b^IZ���%�KrK�.K��]�vKv��j]KV3;�i��JK/kU�$�%�/oe�d�we�%�ː��:A���A��Q��i�K0�:pÆ$����CCBO G���z{N6�}Ύ:bړ>�o%漂�6�f]��Ur�9��t�-	�)v�`���R�Jk`��⹹H�F�K�ڻ��/khB�g^�&Z���x�n�w]N���Hv�_C�,:f�%�LpT0��)DanePxOt�%9�Ð[i���A@��́كn��Q��%U��:�o��X�릗8�y���[��"��;�y�ޛԯ/�I���WXi#�B(Kpv2�Â�,>�-�^��B��֕̇3����e-N:Y�9�`�R�A��-U�u�X��PH3�����B�EH������]nnlH6���hu�
Y��1Am�����d[��1��Yt�
�Պ:�4�����.�DMK[X�=����诩X{�z��jN�$�YK�*r:B&�%����4��r��Th��e/&�+�����޽�����;�����sןs������+��s��>�� @�����s��9Ͼ� 7��o���9�sﾀ�{���.Yr��˫��\����K4�:i��,e�$��?q����e�.�
h�E��M��ky����R���i�Ү@M�L���Zˈ�6�j�Y�&�F�0��. �ǶГm#U�b<���/�����3
�Ċ�x���K����{f�kT����+;J�X�!v��Չ�����B�5 ����C�`�kbkz�i�RXS\�b��+���l/\D��k"˲3�ݘ���m�,Ռ�j.̆&����BTfwR���Y�u�h��ڥٯS��.,��r-j
B�!�*�Q�P����L�nx��mD�	F����سF�h�ek�к�͈T�wfq��v�:�xV�nJ��3�6�/@*\4�ZFjLQK5���m[��m�F]����Tq���֛i��x���埽��{-��\��m�	��ι}L�������}���5�����N�ݪ{�C�xC�vZ9�Ω]�N'�l��Yryq���k]�����]U���e4�3:�F�
��M�{�vA�؅L6�d�E�󮡌c��ɯ��#�,�Eh٨�`q�^��R�ר����a�g���#�����ysuʘ�["n�׈�Q����qv5A`�Vp:������q�AgZ���P9a���j���CdB�s$n}UT�B�b�� �l�-<^P�y�I��L$ҏt�M,�L4�,��x����9��u�.*�-֠���qoi��bi��\��%��Yi*\G��=��5K��$�࣑�M3��-�v):�W �<@�ß5Д�{���ˠl�m7�B$][��Q�f�V��%Y�m�h�e�wa ��,��K�v&,�1ꙜBlm)!��WB2Nm6�:O��:q���ul9Z``�8b3��b,8HΞ$�&x�ӧƚY��i�L<Yc,�%��]jچ��(h�*`��F�E���1��ؠ�È��w������h|4�Ë�(ޜLz�9�	���5C�&B�xJzX{���2�*tL���v�OV{��q�6�E#HG������yZ�JA�'F�j��U��|�9<�sJ:��w0Ȳ³i�=�z��CpI�ֽ�R�����E��|���8Q'Ğ(�L:|i��i��4�Ŗ2�6q�l��ݥ�Q ���-Z�(Ǩ���=^T)]^UЮ�VUeP�xL����4�v�}����	�w�iP��Q�K\�X��H�h����$��4�Z�ۑ�W{�q��LD*||�q�*fL)�_[g����mچ�8jM
�>�a�"!�5ӽX��4>,iїz8:<�"!�Zc���|J=��ZRP�<Id�(�4�K4�:i��,e�$���Wµ}l�*�^T�K�b���J�pY �v]��D��J:��@R38�S�P�1�2b�$UUCD��z���њQe�F�ςS�	5�k�����'�&*�P�t���J�<�Ӻ�_n�ZY���s[�m�܎+�F�ZC�d�����������+YX�e���[��!�+}W�P��%��@�����O!�\��'���$���V�σ�ƯD���FXuA��*Q�:���ƍ�qa��`yx�B��o��8h��:�$�=�QE�~zq ��NQh��t��ᔆ���D.�'�V���Ѐ�������U9��W�֗�US.��b���� ��xvW�E��e(E�!R!H��#8x��:Q���ƚY��i�L<Yc,�s�{��oE��!�E7�_z @�	G�Әx���'��53m�G�*՚�G����ÊE(DE]M�oaa���n>���L1܈�:��>��Ry�N��uY��;7[yc�ZX2Wg�|�����sZ��_k��5�3��F'):)��,�l��ط��͸H����	Z�4��f5�J�5���hE���p�J4�N�a��i��4�Ŗ2�.y�Y�3�l�B�.�7b��?� @��&=ˆ(���I�ˆ�GC����#�\6V&�ѽ����P_e�>���#�+�B1�����V�C]>���;N]�V�:�1� ���c�����N����������a"�j�_�M��JXCefR�E���ȊD#����D�tm��J«������<Iҋ4��Y��i�L<Yc^.���|)�V�ҭ<Lv��	�p]<�<����T���4Ϋn%{�G\�8��'UjZ1�Bb��>>J��"��y�φ�a�8X���V�m���K˧�'!��E�O�x���.�qJuV�o�\�p��8��H��=/t�%zG�;�Lle

hpy.px/)P�ģ�Ä�X�W�yx(��t���(��:i��i�p�X�<I0v��i#	wi�i��i5l5R��1�$18q;A���F&XB�"��J�[T �����E(He�7�)��b�0]�.�/��/�4J�"���z�t�ұ��ٕ���FB�e��Y=YCh�����{;>7�����7���Ҳ#�_v�wz6e�9X�d!�j�xJ�B��T�*�'��G��E��1��c�yh�r����E�x�8��i���B������"-Z�v5�(�ag]�z;-��1I'C+��b\���"0�b9}J���)a��~s���ȣ����WA������6�i�-�l:}k���E�dD(:y�G[g�7ia�Y'	<Q��t���i��i��,e�$���9{�訩�QT��666���iH��G�!��ᶝ"iIh�d��7��٩q]�qӎ��	��I�{��jX��R)8G�Q0ݰӊ1	uޭ3��Rض�E���7,�����8��j4+�R-\�J!_�)���Ӳ�N��e�ɵ�ps�e�V�HB��[��5[)GK�Ӗ�[�r���V_�Ie�Iw$�%��R�Z�]�{%�.K۹w.�JR�)JRKV^�K��bܺ��K�x�\��\�%�r\�%�rK�˗���ԒԖ�\��JK�-Iu$��%�%�.��ܻ�w]�ud��I.��yu+$��K��%�f.K�w.�n�L�KRՒ��gvJRY{Z�)$�1;�^��r��d�]ܹ%��`a�|i��4��4�L,��8a�H00004�񡡤��A���/���dXdkH���$}[yl˫p����,}����앗�A�U����偪>4�.�S%��Dʥ�̥�p��J�eދ�"E�]E����Tm՞\��1SG1Cs���-�����3�6�.�5�{h����
���Ӆ�
�`�L�t��T�Y�3�l*�R��ǺlS;K���ǜ�	aP�|]�4Ȫ�M��}BL5�1����_*��1s���w��Jg/{�{i]��٬w��-�Za��n��|� o{��s��9�s�� 8���{}�k��9Ͼ�� ������s\�9�}��`7��o�\�e��,��,�N�a�4�H4�Ŗ2�s�ccch�*���D8a�#�~5�r�������.����Gg}ș-p�DGڬ�,��ݒ1�D0�Ϙ����U(�R��p;X|�p�-�x�0q��% 4R�4����f��F4�8=k��|�hоz!}1C������R$,�08���K1QG���Ox��0�0�L4�L<Yc,�&�C��.�p��\_� #G��=�����r4m�k�)����_+V0���}�%�ʯ��PQ����ãyET���N��å�����i�xj,<5'���)�ç�-��6��|���ŋ�m<GID�QkP�$)Eu.�9d�8��䰅�5H�AТ�a�N�x�0�0�L4�
<Yc,�#��[���U�p�^�l
>�������l:��5���Npff������QS?B��)��u��rL�jF�r@��EZ��  $g��|�mU^Л�dO*���F����f�t����^%YJk���v��aM�J���Ј�Y[�9��.	�O�mPFt�
	z	d��Y��d�C��*���LC�GF�]���a-$5B�t�IӀ����b��p� ���F�U��y^a�v�b\�� ��}(_.�`�<�|ڤy��h�qx:���3,�Z�l���N��rt��U')��`��yI*5^ꊿR�J]�����}�p���h��9Ո�!x��*�t��:I�K(�ώ�a�4�M0�Ŗ2�bփ�662�X�G)Ժ�4�W9��p�m�h��գȴb>
Qэ���E�8�`�4GBŠ ��Mk��`��5/�{���O�B%R�P���!���l�n�;qR<��Ϛ����Ǆ���{--T%���eG��z��	!�į}P0�8��#�O�M("a)���F����]�tђQ%�t��4��i��aG�,k����:5r�� ���ܒ6L�FL�5�j�k=)�d2�r��#��O�ξ��O.{�>�-�����qD�o���#!g/Ø�DӒ/v�t{ve�7Wqn�������O�9yo�r'�A*���G��Z�(�7�c<���޽�&bd�&"~^�:�#�����RTH�4���(�L:|a�4�M0�Ŗ2�L8�Hа�>�_a�` /��9�SΫ��{?�;�y�/OYD202ʢ�-g6��LL*t������+Q��������ͩG���J��Ě�^Yz?�0#�y���~�/qN#����
����눠4�Kc�5a�(�㉟Rr�"U���q���i��Z x�/��i�8#�܉Bc�q%F�e��&�iG�4�0�L4�n�<3�I,���
��%�p4+��	�=�_M�&`.q�r�ܮ�U6Y�1"ַQ�
�JB,2�ti>�wI$l9��h�)g�y*}T]N݂A��'�e�X_vͰ�=.��=y}���L��Q9�"��F���qf��y�u��t��Y�1^9�w������;y�ֻ���oA�
�c����ϑ�F)�ۉ���<Q�'o��s-[��yB�Fj��#Z����a�m|�:9�+���F�*���B�
�W��Y�($�>��PI�΄b0�L\ʖ��钼��i��8B1�F��6�e��'	>$���0�0��4�H,�.�)��V�4��6� �ϲMR�yk�ZXݱ�qu�E���qfB�7V`�D�VB�����$�Q+�Hh�&�q��q}�P�,/�قX�&"��"Y�#ؤ�Щ��/Wq��x���ޟD6�Zyi�q�F����ƣ�"�؏���a*K9���"���5��h�0J�m��$�f�I�Oaf�>0�a��Ag�x�'	v���Q��h9����q�݆�^k�i4	!*9=� oX�O��7!mEu����\�>x�y�#�yR�$f�8x��ۄ#����#2�(���=�ks�T�ND�m�j�R�(��o����7������X���;ZL��e���^�h}���<0�_öٝ<�j�����5���iن�%��LB,(Ѣ^UM�'��y^!yx$��Y'ĚQ��:i�[xY��i�3�T\���6�j�jn7ހ ���qui�Q|Z0���E���È�y3D�0qLB�.b�͹ո�M�8.���i�WҔ����Z0�Zz�KE^/<�yz�%�2��>���]�J���p%�ⲖJ8�T�(�ŤgxuG��`�Y-�e,>�h�CO���)7��}����ZP�W�UUU#

�a���'�_�;8?���+�χ�E�0��E zR9No�M1��6�QL% $H��L`�&	�b��&&	��� ��a��H�X���� �$� 	"�"$�b"H"`�"(����Y"`�"&����
"$�"H$�&"&"&"$����%�bX��@�"&"$�" "!d����"�
�(& ��& �&� �"��"& ��"$����%�"XX��"�""$��!`�""X����$������"��$���� �"""H�� ��b"$����"H��Y���H�$�"H�X�� ��"X�$���$�"X� �"�"H�%�"�$�"H�X�"%��b� �ab%��b"X�%�"YbX�� �""X�%���%��b�!"��"$"H�%��bX�S%��"���&$��"&"$��bb��"&"$�H&��	��b!f �""H$�b��"&%�"b"b!f"&"&"$��"!d�B$��"H$�af �bb�"& �!b& �""`�k40PDLDL,D�A1D,�D�ID�IID�I LI�D��A$B��$DI ADĐ�D�D���0�̆@8�$3B��$2C$BA$2Dđ�C$C$D,�I��0��K I���$I I�IA$$A$0�B��$2A$!0�3L�0��0LLL2A0��1$��D�10LB�A0I�B��$3@��@kX	�XBT�� e ��``RC!L�� aR��``XRT��u�j���*`0 �Ȅ2��qk����"RCP���2,�@�00@Ȱ0�"�`�4
@
@Ȅ�a�HA��F$5
`*2� ��00��*��&"���(��00(���0,�@a`(@°2$��@�%��`aXQ�� ��H eRE eB�@��D��A��A��Q�`F `eXD������`dBA XD�� %HP��H@��` ��BF@��`!	F@��`$X	FCPd4
@J��@J!(@@�	,0$00���ʐ����!�		�)�
H����b`���9�
KC2C2C30�
IC$1����2��C0���2��C�1����1��3
A����2C�3
A��1��0�1��C$0C$0C$1��),0C$0C$1����
I�C$0C,1��)$0C!C,2�2��
A�0C,1��00���),1��C,0C,1��0�0�������
K���������C,1����2C�
L1��C1���!I!�`�H`�Hb!�d�d��Ba��$�a�f!��`�&�	 �	`�%�`�&�&�`�&�"	� I �$�&X"	`��"	 �	 �	 �& I`� ��`�	 �`f� �� �"	� �&
��u���DA0DAIA�A�A�A�A�$A0DA0D@�@L�A�	$�D��2AI@AL�1�L�I$�I040L�3 ��$@�@I$�,�@K@I �$�D@2A0@�0�2@I$$�AI�$$�A�2@2@I$�� �@I0���	@300�L0300� �0��00D�1�LA0,�C04 �@L�D �00L���!k0� �����&	��`�&`(`&��	��Y���"H(& �&	���`�f"& �&	��`�Bf�&
	�l��6~�;�9σ.�N)�l�=O���p�AZ�	��O13���\����g}|��G��I����f���}'?q���>�������s�}��G��})Gǯ�+����}i��|?k�><�|G3�����pw���?�����>&������fAP���������A�|�C�EG�B��* �����>#��?���`��H�ڲ`��_�����w��#�������T@��O��8�㊃�ϙ��x��~��?�p2F�>���I��������n��nξ�3���]n�q�iyN#�TD�{6���&?F �����!̪�&����
�@ �@C%Q	��ThD
T]?�Bt���=Bf�����6�y�9�_��#�?��(#@D"��  u� �P"��@���g�u�C���}���'?'�+����G��=� �� �?�}���HG����5m�~�� 1>� �-/�����������~G�����/����;���}o�6���?�N�	'� �'���Y�~��y���t~��P >c���wܴo�~���g�GG��c���|G����~%P�����+�߫���l5�>��=�~�_!�;?����h~��Dyy\�j#��~|�&�p*��0i?FϤt��?�`h`��fr8�&��ٴN6'���?#:�A��g�q����b~�����?W�����o�k��@��9�����} 6q������߿��>����$��_�}:���s�����_c~�~ԅ>��O���x�_!=�R���><?L��+��O�_ʠ* v���?��w�~I����_ �����4�>��(c�J">��`�r09���]g��t��/���@>i�~	��m7�^r�^���@T �Ⱦc���1>���?!��@?,����|>���N�K�#:��g*����C�&�>?��(
?��~�~@4|ע����yO��t���>I�g���1v}��щ��[ר�?��3�#�&`����N�����rE8P���6P