BZh91AY&SY�HBxݑߔ`q���b� ����  b@��           u�-�!*����D��dU)4`
����U%IED��"�(DH5�%ER�TlhE�EPP;D��S��P�����!ЛQ�HJ�
قJ�J�E�E
**ѐ$
�����%UA� :n�R���A�b�a%m�p��fDE�ݚ*B�*�"�J�IIPkRB�ZҊlʬت��HIV�2�TP��)V�5��r�jU��  �JP 
w�>0m��HaN���+��*z�q��AZM's�U�S*�6��m�ХZ�˚֨鰽8 Dv��{hT骪T�F��¯�%$ �w�G���@��t4�R�:�]�y��J��^�E�M�����zVD)[�{��^��K{'�=W��i����RUH�W��p�IR<���P�.��E"��$�3EAQ�$� �����T�D�_:=�=J�oO����6�J�y��EUJJ{��w����*��8�R��{��RWmR���<�R�ۭ�7��)Mz+�{�J�:�T���J�JB��>|�  ���j��l��ץZ���8��
�n�����IUN�<�v�%==罵T�R=����%*�lzn�WM[�{�
�N���T�R�=lن�c�TɅP��R@ c�:��@�)�/{ҥ@��{ޥ*��G��J�:��Oxz� I�{�"��U��D��݉��]5�㧧=J%%.���"��U"���Z��UI�䤀sϪ�JP����*u��wn`R��g	T�Jw�ڥR*�Ig*&�����zP�R�wPU*P�K�WcJ��p{�  ��IJT��L���R����y��| <t�[��
 gOq�E�[lU*3��B�wC������ uE�\�(�  o^�UUTA	$�(�|�@׾h;cp� B���5��h�X� �t�@ �X` v�P�� �p�@rTQUJR�֠��F] 1�X�4
7U�N�8 �a�	Χ���� cs�G� J� 4n�p��I*��R�� Ҁ��JR �| 1��ց�:�)@3�  YX �� ������@��\

8  �>  
��B�M	 �S �J�A0CFF`�0D�i�IQT?Q� ��MF@5<�%JP�0    T�"dT�A�	�F�d0�&LA�$�J$��I��d�d`��4� $SI$��&�j��&�#���G������?����a#�������g�����.GAgvC|�n�� yR��܈ *�D@EO�@@U��舠��~F�!�����?����z��dPV�
�I9��"�
��G�`z?�@�H/󊨢/�����`���Ŷ-��6Ħ��-0m�l��`���m�l[b���m�L-�L�6Ŷ-�m�lB؅�m��0b�؅�m�lB���m�lض��-�m�l[`�
`[�6�-�l[b[��m�l-�6Ŷ�b���#b[ �-�b�ض�-��1m�[ضĶ-�`�)�lJ`�b��6���-�l�-�i�l[`��6�-�l�[`���b���)��i�l[b���m�l[cL`��6�-�[ش�؅1-�l[b[ �-�m�l
clZ`Ŷ�-�lK`�ض��e�m�lb[ؖ��-�m�b[ضĶ�-�lK`�ضŶ6�1m�L-�LK`��6Ķ-�m�`[ؖ��%�m�l[b[��Ŷ�m�l`��6Ķ,m���m�l[b��6��$e�b��6���-�l`�
clZ`�ض��-�m�l#ض��%�m�l[`���1-�l[`�ؖ���m���[b[ؖ��%�m�l[`�0�%�m�lb[ؖŶ�m�m���li��i�l[`�ؖŶ%�m�0-�L`��6���m�l[e�#؅�-�lKb��6���m�l�`�ض��%�m�lK`���%�m�l[`�ؖ��2ؔ���m�l[`��6����`�ض���m�l[e�c��b��l��b� �!l#ض��-�[�lض�-�[M!l��ŶlB��)�[�#lBضŶF-�m�[ض�-�[0-���6Ķ�-�lK`���6��lU#[`�lAm�Lm��1@-�-��*6�@�
��؂�e�P#�
�� � � ���(�[`�[b�lP`lm�lTm��`�� -�lUm��lTb[[`�lEm��6�F���
�ت���ر���E���V�*�[`#lEm�-��"����(� [b�lEm�-�����(�i��� ���"�b�lm���Q�
6Ŷ*����@-�-�E���؊�[b+lB؈� ��ب�[`�lQm�-�E� ��K`) �F�(�[b�[ ؂�[bLE�*4�V؊�blm�-�U�(��V��X�؊�`[آ�`�l��� �F؊�[b�lEm�lX�F�S-��0����*�[b�[[b���E� ��E� �-��Ŷ-�m�l�%�i�lb�ض���#-�l`��6�-�l[`�#ضĶ-�m�l[b[�lŶ�`���m�l
e�i�l`���-�lb�-��m�lB��-�l#ؖ��-�-�lKb��6Ŷ-��l
`�ض���m�lKcLb��6��-�m�[��m�lb[ؖ���ؑ�lb[�6��%�m�l`�clb[ؖ���m�laLm�LK`��6��-�m�lal��%�m�l`��6����m�l[b��6Ķ�m�lX�Ilb[ضŶ%�m�l[e0-�LK`�� ��s��75��W�fX����J5���:�9W���l6V-�ݕkIԊ$�H���Z��E[��P�����:��*��ڕǹPCpZ��B��6��aooa��t�I���i̫*�֘�ɐ�6P�E��͈]z�U�U��J��c]�AM�K/} ��XmǒXx%�6�K&�|��R?��w[�^���h5^U^%��Rd����k��%e�LkwA, ѡ���r-r�(�)Ƕ!�n4wK�@1�)M[�-�-dJ� �Op��+R�ـ�YQ����D*�0ȆR�I���X�{�7����J
F�ܛ���w4��bh������H�gJ̖T�%$ff��Veiu�eahk���!�1��mk�i�[36�k��!�X�x��,Afg1!1��h��L�A�=��ǔ3b�9yx؋,�:yJ���9lZ��y�hnh���)S#`v��a,%�lDQ7�v�0��N�\`���]�Pn�qZQ۷���NLtV�6�ۘ�f$�[�j��m@ϰGvGh��f��l�櫱��w%7)kС)�P'I!R���v�S9�-����Q��6^Q���m)��%�N��*�8$sE�nh
����q��U��P��ܶ�`�X�a2������[�X�cV�
�7L.��RbAX��Rb4£�2bͪ��pLY��3%Rw9iR,y�(��U��Kn��[�t�HZ�n��-݆)miLT*�nm�-�/DåF������
trP�*^��j8I5z�&jV�a$)L�%�KK�Sf��Zͥv,Z�;n+��&`j�� 1cŧ.�^<�rQ�VިTr��%n�[�[,���,�טsj�m"���8�Vj��9�yV��ah����n(��R�A��yuqU˚����
K#*Ģt������Zj	4B�G�0eۂZ��̃}Hbi�y�j:�i�֘`�-���m��/tT�m�!�&4�f�L�9UP5��e�3i,]�mK5iJ���D�a�t�ME�B�����R	�w������ҫgO	Y�1�F�H���	��L�<X��.���$2j	5��ʨ�ѥ p����Ö�H0�UV�1h�����ѺIJd�8���*�N��KCr�@�6��%�;�*U�	�sFԖ�ܕ�I'zQ�����l��RU�t)���ݻ�,]8C��lX��B��ݴ�'������aS�����F��D����Ef���h]��!�5�QUd�٪�NJջQH�ɒ��m�(&ݔ�D��̏e�(��b����U��B�eA�ho)X���
$�Y�)�k_�0�T�:�B�
�(fl"�;�In���U���S�diͤD:�lܧNX/a���#B)6��2m��L�C.��I�60�2 £V���qF�
�B�Z�[���^��b�]ͩ�U�nIYusNAwt�ٺ%J�kf-�I��;x�J�L�Xd��˼(�ȕ�Mʶi���r�,�1�D��q%�� U5�v�U�PO`Rka� �hͼՄ��v����7a���Ge�������zk�e�F���d�ۻt��0�g!׭�0�̰���+.R.����wӲ�ӳ�ʱ�"��5i+G��Z0�
&��T9k��я/m+�݈�4��p+�4K�$G�ᆦ��[.ءdx���L��z���Y���1��j�
��6�d�̥t*f�N���C&h��'�Z�D�/!b���3 �M�g���E��Zk	�qR	ܚWQX�0�T�9-��D�;y��N�C!��l��@�'
O�!ҵ�r�:�9�V�2�T`R��Z��G=�^��U��1�F�r<�з�s8�0䊂�(��tq�7q�t��@@ ��3CW����G،,��y��3pZ�ܦc�a��d���kU4�f骽@��e�E�чH�n�%]��'t6Qs�kBbAPf���n`p�4��s�;A\�Y����l�o6,W�!�Eâb�r�	o��{NU�u�(RX��Z�b�1+h
Y��Sl��*CD�y�Z�i1R9��h�+%��6ֳ�iI��̼�%�lܵ�0d�ۉF��n�b:�ݺAmX
 ��h�aʲ�JS)�u$Y��uR�]���b3X���|ͅ����,�v�(AV�[���Nnԫ�T��Y��,��Q��xn���p�,(�u���j��\��%35�b�Hh���I˺q��$KgPM��T
��uU.�fe��*����@��b��	����àUX�����Ѭ��yb7��o��up[�����2�V����u�F�P�#i1�B����;VY���
W��pc1�0�+p����	��wm�-aZ��&�P�h���v����.�͢��*��0&��Q�����Õ��M�L�,L�1ASb�AIJHI�i8�F�q5-*a�R�w2� ����xD.�
W3$�X��td�mE��qS��qJov#iXV\���3�%y���Ĝ�
f�ؗ	����CL5�V<�n*�jMP�`�U�7A�$�4ݼ��f�Խ(S�CC�:ݢD��K�(�U܆&��؞���2�^I+-�+ZqlWp�e�z�L�&��UU���/ڗ*��-\��nj,̓CY ׶��o�V՚�]�bu0�m�I�Pn��U�҇/cUPF-gIm^@��ZcO}��K>ܖ�`�pAS&,�d�R�)Z����R� ݝ%�(�y��b.j��M�����V���� s�j�`�ܰ�7w6i
טmjɛ���aSqmْ��w.���Z�nVl�S،43iM�ek��%�e%8]��.��.Q�tw�;6^[�̷/-ly���R����P�{lJ��h���i���Oע�j=��j���*�C�S.�0��٘��B�����a���&�gv�a��N�H�"(�����e��MtX�Isc]�Սy�V�1$A�H���*�B�jZ���-ȴ+ڤ��=j��u�Ѥv�
�0h��+fk�I��9C*^��fe'�@�7�R�)F���v�ʙWK+Q��Ǭ���Ҕ(3��,���:�$GW&�b'[���k�Z�Z̲�fR4��SL\D�EDb��۠�������#� f0�2dj���&�`(�T�%j��u/Z�j�����q�D�;�캊��]阦�^�6�X	(Q.�bklScu2�ͷՈ�S�q�fL���bܺ��6���`+:�R������e�r��m�5m,��A!~�H��.� �36b�KQse�&Qo(P�t���6��tJ��0��Ae20$��4��N�W*�#n�"靫��k��b�6��c�2���3��Z�c*R��ۤ�36�ȽW�	cP�A��-�+F6"�ͭ�Y ���K�wʶ��e��FVU�Q�vj465�6K1�kr�^ؐ�xw���E�Y����"ֲ���$֓8i]�k/6�lK�5W2��^0��a-,�B�X3ne�a� Y�4�	���{H��x�\4Ŋ�)���L�.�!zX09���)i���;[	Ѝ �S����3�����Z%��`8��
U�p�y�(e�a�`�{���"'($��l�r��@q��0d��xa��5K۸Z�Y�QN���8v��hVe�=ep��G�J�2`���R*��DeI(�5[r�;�[i�&9�E�;�KC�(,Ԧ��ĠփL��)��&�"a�C$\T�m���3f^���zhqB�ާ�VE���F׭�d���B�$'u7F+e��&k��Bj��Yv)E&�C�V�n�V-x$I�Y�c%���f�y�U����	W���eE�^�Ce�C�F�<�̶�ꔢeܦ�������utΩ�<m���/'�/FM�õ�ͳm�M��&J[�eh��Z�Йv4Z,Zʻ%�V�`��]k���I����$ص[t�I-��+��ٙ���ə"�W�k�%�V�JJTW�LŮ�	6�UUZۻx������vM�ƘlT��u+�4��#1���(
˫�8-�kP��3H�;�o���c*�#��������Sd�FX ���q%m=I^��/0a�aJlʓ�ޛIŒ��y{�������kt�eh�cota�n0Ė�FUli9&A�X-�%m]^�.�!��ZN���^�u�/i��aL�3qJ+]
�e]3���^�Z
�Ēblyw2���Wc@&1q�֨�p�B�jf�J��mZ'��͸)=�~r�^-&�Kn�e�mXւ��5�E6�n�F�2��.��E�$r�nVY��6M��ВŊ�F��z7,Yʺ�Y$��ҌX�Z-����A��X~.줩m�)els^��2˱�q�$ކS�����5{�JV&�ԉR��%:ЖP�3!�%CJmI��]�a��h�H
�q�~m6m�lm�z���PA���M�,�մ:rZ����S��^ߐt���d�pbm:g�W�U�s)^!��cc\�W�ԹW���n�j��Z�*\�3{���4V9h�.�sN!f'c2,����2�1���P�:�{�T��N&�1��mV�KĊ�-����EU]�*%J<0�W�I�KR90^���|v�e��֭l�ha�f�o7|ō����*MGj�CR95�I�c&: V���D����3$�Q����f`���Kx�lnk�U����:H[� �Jf���uD�Ѻ1a�b���dj�%��sR�@G3)�r�0�zM��7GZ��\�*+F`�f���OC���R�=4��w��j�$��'-�/r�ۻ@�f��b�x.���[u�)Dp���+yLf0����T{W�yj������ql�Zl<���i"j�i$����^�ZN���yq�dX/)C��b�X�ba��������z�M:�s.6�H�J*�e[�qn���§�nCV�s�b�*Mz�%��(�p�ͳ���k5
qc(�F�X��j�8M�d���v޴�Q��"sp�5�tZ��Z�Fae�y����-�K9��xr�t����x�]ZQDōX�hۀ�mh�R�T]�[Bb�W4�"ͼ�e�pI�����-K�Y��(��#�o`T�z貶�&^���t%�
��@ՠ�͛�ctYC�����#U���$$�ubtHf������{�I�3X�{-�q�΀�y5�����sw*�J�1�W�j�1�aC�1#�FR�Qj�2�tQ��c9���Ak]\x�+a2@�~�9F�^U���[�e�j���VT&lۗ�k!F�$ ��FLE��+��Z��2AB裞�(�:X�x�R�[F���t�a�@U<ֶ֨�Ncc(��N���cp�-�ݤ��Y�5R�Df��Y�B3Yn�l˭5UU*<%hp�R�wY��0ݚ�w�}��&i4K�h����̙4՜��b{��Y�G�r�T���H'<��YM'"��o`ddӻ��J-֦Kd��ۗ�����ۣ(����4���{w��L�K�-3swf+1�nK!���Kq�F쬤�dݥc��+���(ݻK��:��2���Kn<�t�9����)���4i;�ӔD~��9�J�����v��y����-�QҢvn[T@F�jωgh4����44��(����e�aX�k6��RV�[�仹�$��5e-���K�35+��7K�`k7,A��,C���r�Xb�J]m��ޫ��-�%`Wa5%n\Q�pJ��Ƨ�eݫ�{�JaQ̑27(���;�B5q����x�)Cs	�r%K��^iH�#B�X�GXE����QD¨HΊ�����s��U�j���<��w��#5=U�Q\Q,�-_&��˳u-Z)$�V��-l�C�]��ru�rr����MT����E(�j�-��X��K"=�J��KQsj*�.�@��&��m��C��(��m���ɺ�Q�MP'Q��rYi�T���Z�W��[T���8�KU��AD%�⺮��沑irv�F�iĩZKRKylFԼ<�T	�n+�`���J��Vj�>��k�-Wɴ��iō8�*h�x�&ִu\T��ֳ�r��Ե�&����u)�iE|�G�ĩ@V���z�^�f�< �U*r[DKR �)�j�OU�{Irx�.�]����.$�H�'D���4ⴜJ%���(��qW_\T�i�R1U.��g+�ԩ�ՠ�n�q�ռ�JN����}��]�Q$����T�j�\Wb�T-d�)�I��DZz��w�F�RX�h,��W��6�\���K�(�W%1n.jr�J"
���{UR��7�cĞ�i5�dR�V�wKY��ٙɋ���#�����mKE-E��
U��-��Y�Z�N��cK��/��O+Ž�v�8�KWr�t����5JR�5���Y�<���I$�*JRMF�X���0n�⦕��D�qH�,���{ٙ1�TR�J%�%�RԴAx���*�-�ifެG�e�u��G+OSi��f.Ԣ�]�4�ĵ*�z���҉[I���D�-j��VR�Y�ZX�Q���Đ;��F��H��-P����bv���ڷ�A6�����ԒR��v���#T	��YIZx�KRj��j�4>4�Z[�j�I%�RIP7���p������-=�`�n�y0g�5����>H�%Z��ĭKR�҉V)�R\�Y�$�,I��IjqRN%�h�Sjz�Om����qg'�Qj�^�`���Ir榥żQ'�V�J&����+86M[j5|���V�T�DڍLW��QsM�ֵ5rRՂb:��kq=J�jZ��Q.�5x�'V�\�ԩ.I��Z�Ҁ���I8�y��,j�o�Ѭ'6�][ p��of)a�:e�MnȐ;j�Z�4h5q.f�K�*��[я��wV�G+�A�E-��-J��@�Z��Ʃd.R��&$�H�֞-���VDȜS��
r�u���~C�[��D�0?�ķG��>������=$�x��3����)tܾe����׋9O�1wY�����/F�M��D�l�[I%�.��*�eݩ��n
ڻf�5pXY�*!.� hǽ{�:s�]sD��=�"��D��8�b�*Z0��g#���K��V�૕�¨������%σS~�]��Ϸ�Q�e�1|i�N�/wWdR��g��V
'(.�S]-P�A����$�ݭn�v��h�o4	���wn�y�L��z�fd�����S�u%a�{�WT�hͦDRJUs4Z����[mGWD_EO��X�SO2�<�|� T����(�g�k�o��(v`���՜z�H�zXjNe&��� Jxt_[}�n+��9��)tV���T�7�y�gG%{[��3�{�����p{8b)�0S�;�&��olt�4�Qr�.�Z�l3-��e"z�n� �s�-����`ڼd���f�K��4��Wo�)$�i[ֺ[Y��Z�b]x9gM��^�ޗ�>�qޔ�>���Sua��Q��P��t7T�N����f��ݙ&^ꊜX���/���;�eVt�ུ;:-X�V��ݖv5�xż�r-�Ѹ�圖n
/4�4[}A��ݹ���\u�1(�H��r��h������zX�89��׽�f?_)�Ls��f�cxk7�"te�	Ne��{��F��tsreF���d��oY�yv�J7��IWcu"���k��ɣQK܋:s�,�R��Yj�;HTĹ(�Jf��51�Sjj����74CWV8 ���8dN�٢��v�v�����/���i$�����V�<�p�SDΥ�Ӄo�t���"�=ǹ�z�F.�<��]LPI]&wa��,�l�Ke_gt�T�j��Q�����z��nU+JyEykʆ�\8��Aƣpv�&�V��wS;kx�<�{���wt=�i}��^�+\�N�K��>6���v�B�n���*�/]�4��Z���c��)���vsftY�9f��(q9�U�2�]�͋UR��dC
��h���*��*摘t>�oAu�������ޣ�s��\,�[��������j������m��pRԸ��T+�6⺜���	gX�뭀��p�NdW�M��Ģ�UD�3��9���ϱ�eѣ�F�_RЪ������Ar���Ʈ�g�g";�s\j]���`���斌g+����`����Ϩ��nؑ�[��0!6�#l̕ԑ���ACX�ꦐk�gMuV�nq��\�ya�`]��c};�6"��r�arŝ���
3�F\���F�.^����`�
����uk�d��hf��T��t5;xE��1M�7��3$�;L���B6�9��<�>�(�'9�wnF��_){N�u
�v���T�׺��q�F�N^ԙ�F���AӖ�'��ܱ.x���y �]��l��[Ak�S���u�Ϣ�3�قgK�R�h��n�:���"7�*�o����W;,`�az�fV���l*�Х,�ӻQ1}ɇo�����VШ�A���X��v^�]�B�(٩Ӓ[���R�:�Lr�J����CZy=°�.V����;�\&̵��ɗ3YL3k�2i�1����r�������M���+wx�)�:�Zr�rPۢ���ܭ��钊��p�[ebV����]5k{�X��lG�N��H�Ry�T(r�@V֪�V�|�K]|���Ob�A��>N���=�7�K�ֲ˛�d6u��h	�;����٧70��!d��ÔGb���C��;��|wf��F ��
�{8Zsr	�']c�T����������xzɡ�5�tw�"��L��Ⱥ���|�\�tŉ��_%�wz��h<(>������xk�P;��-��2$S̀��5����l`CO��_�]���������q�oUң�\���I�*=�jA��y��ګ8��p���a��c+vʊd��-�G����$g�z��Shև]:�)�����7XS��8l�n.i�s}EɫU!�s�)����ܱ�9���л,;��6$���R���o��	47pTIғCZKҪgNQ�g��fu1ru�h�֍غ���{Or�*,��fis�;��fu��u�lJ�VPQf�4B��P��2��ǳ��yT�JZ�C78f��#�Y9B����f���;���wT':�m��=ʍ��Nk�����+�,����tW��a��-+�B��jT�ES�m�MŹ�m'�<s�cd����W��lGp��6f����T�K-3����Ȳ҃��Ǭ^˧��)�G�L��Đ��'Ccb�7`����x�۔��D˔��ȅ쪡b_J�z��r�7�(gX���U�Rz���2�<,A��<��ǽS�����d|�"�ƻ�1��a��͓3�1�ݻN�mJ�#u��On��9JN/"U݂��N�Qd�2%Y�`kwr*|N��_k��p�͕*#t�S����Ź�:>6Z�]��<J�҂�9�Gou��O)����t�[��G�eFH53y�׷�V�W3{{o��� �h����'�3Be�����ꦢn�o��K��q��$���ՉVS�g4�e���n�*��u>(a���m,#���U�ѹ�t��\�ԃ�Ŝ�`�)ζ�qe[�4�p�țDP����A���z$���9N��7<���o4}���YN)N��8.��eY+k����ˇϓ���	��U�,��F.��Y��*��bz�
tr���C�����)g�G��Z�4����l�YU��k8�)|J�,
�g-��&ī�s�[���;�8`m�(�9��X���ݔ���
:�ك�f�`�:\�Z�˙��է`yٛ���)��q��R��������� l�+Y��})��l�1mH����b`/B�<��� �C�'?�Z:�u.�L��<���'Q�kK�ي�9�D�|��5�{7��Ǫ�rR�w^#����с�sv�	B����#ʺ�U8�+C\/FW��d�۽.��f��4@e�/%e�Ai������$��9��n����"�^6�����g9V� �A���ޝ&�jM������N=8$Ofw���C��4p�r��
����١7v��MLu��+�u|�Ņ��F>[��v�v*6H�_M7k}�em�.]=��nE1]J�+�3�����5����c1W;��9i֜��� _V&-�x[��^+�8u�e��2�j1��S�5��A�%qL���Y}�)AۻBorͼ夦6��W�S�Y|L6�G*o=
C����g^o;��]p�����-�NH�u6%5q��ヮ��r�N�g"/am�V�X�V=V�$�Z�UH��x��g��]�:J/�okwE�\�3�9�Ðx�h��w��Y6��\�U�J*�Q�9T�TUx�vv��8�1-2y�N�CYg,m�H\eu��cMs����\��쏖gt�
�r/]��kg)5'�v�y�:ܭ��ص9rܮʨ5�f��h�d������+hPJr])wWO��告��*ܫ�q�PWx{R;]�6�T��͐l�'d�ʦ��XYy�ӴR���x��F�X��1�eK�Q=�z��ʼ(v��K|�����H�*�D�X8kk�oj�F��!M�|�yuw��eޢ�7R��z*��4u۞��U�v0���O��QdL�#����e���[�r�������$����Vf�'+u��p�oK���m䧣v�����&��JB��պ�+T���$�(��TI��i>�:�A��@�;��fǕ|�,,,��d����O5�Z{k*�Z钩h;��9�ig%�ճ\�V�K��Ne��n]mC:�mJR�(�6(���M�!:���1����3l�$���JGe�6��Yop�ʵ���s	�G��')`{�eܝOs:�P`��r��1�&Q���)��GQ.�虁�S��{���*��u�{4�l{EVX$ߵ�U�6V���5��KU;�s�c�y��ַwJ`k�4ks�)��c�����4����Z�+B�V
�e�2�ɩ����[�KZ��9��ugHYq���R:�J�l:��7��:?$��Xb�Tw�6U��8+�;F`�3�;���u�@յA8�J��O����o��S��h��T���y(�^���P����f���6��v���}�%�GSݎf�u�T��T��R�;�eb����4�L�	p��$R�%�ҫ�c��x6��_-<��ws�n5�΋/�����=ڪ|�X�����L�e�T!.Q����|�qn�:u�� ���2�q�w��9hǿ:i�m̤�:ߨF�+Z V*ˤ� rȌ���;fҭ�o�44B�i��r���H�V�ު������3/N	ؙ����rs��J���_,�ks��(w`Ô�9e<��^Z��>��G���Wa�Qzj�EY��W�O��ǹwIj]��{+d��nV��q1e^�\�ؓ�K��y�ֵ�;�����j*�nGѩ����El�黯����YJ<���^�p�5�j�E�������8�茶�nN�һ:���-&�]��H�ʮ�l�JV��Lۨs�B�97�L�+�rWuY�z�vVKٝ=��"��qI��H03��u�7��=;����w;��tE4b����+��S$���;q
�H�w��0 ���Qf���L���wV!��	od.~Uy�t{�6����1nZt�t�(���Τ��%�hp��b>A����q�0�{�7J��
IΝ�������a�wL���J�1�b��r��H�15�XwZ�|	�حp�I����ͬ��Շ��k�t�C���a}�A��3�r��u����G9o����4�4�cL��e�w���ژ6��R��3������ևۡ��*V�&�ri]���w-���ބ��M��|�t����;���%�]��vvÔw3�B5V�����x�+\3t��@��Lj�e�z��XO-�������\�Մ5�Ju�ӛ�fn%e�7�gv�Y�ɼns6��J�BZ��B�w�0eލ�y���dK=մ%+t����{�v	h}�[������m4Fд�΄�}/a�t��!9��`�Xk�'�B�6JX�h`:RV�f�f6��]�ϱ��ÏMN�rq�[��+pS=[��b���v�Knj��Xɍ��y�u�+��C����G:�,s*���p�ĵ��̻��&����rm��j2���p2�Ι���Y�b��ة)Gw��L���ee	�ß$��uxLɥ4�ٰ3�7z=�u8��O;Nɶ�i7�wue�moh��o��
��V�켋���b�X2�t{RY����n�K�^kxz r�^��[�;+������ �o*J�u�,w����h�yz�v��%��Tb��sn=�]��7���5j��s&Z���.�n�=W����b�Gm�9v��1��w+6�t��cZ��q���m
V����=��Z����F�m1�&)r��;�}Iͅ杠�^Kw�ݗ5cT]�Lw$be]�Yo�����f��!VhWsIT;'@�,] ]Y�,���mj͓LC{Z���ﾟM���	l;�rlb����1��[�:�޶1�X1�C� ����
��QQ d���O����oױ��}���B뷍'u3��5�+�(ݼ�Nu�97Ƶ�3::��/A�J�F������1
|=�0q�o�g��+%$��2�9{Aٷ�a:�|ml���97$�د1U�%9�k\ŷ���J����݌#7x�H����y�w��������H�p�+��h-���M�*��<���9�v�U%�3oYݝN��<��s����<�+�������&v�^OXq����ݶ��X�~x�Q�:���lM��+iw�]2��b�i���\���^f�8�u�DZ���#�+c�Y�i=�f�m�n���A��\�ӵ��7�i$dR�	UG�NCZ��E�n �t�Lʽ����"����_f��.��q޷��y�W�@=�o���R�+ˮk�X�%��� �*_h�GP�_.���#�r]^��u<綏�Fk���|�ެd�����=���;�sz7�T��5"�*��<�yj�p�¼�IPة�� ��y�<�sV�V��T�p��ȂO9�97[��ECSz���Z�ӱR�n k|�*�bw�.�ٸ�R�n!ʧ��){+t��/�Y=��ʔ!�{	#H��
 ���_,#�_Rk�y�Q�R��s��������|A���ɕ�O������(��/�����p}~���C������Ui��C���FR$��7CA������K�ȳWA����:X�j���N�Ƈ*�WbHk��t��ԻN��O��N��'G����MM��UyYQn)�eu��
��h��ɯ���ظ��Z�^��=��)�R���Kj("�N�L�N�G&�қ�L��m�n��=@��l��[���l�&۹�3�K̼��+6t���M�cR����M�e��dѡS��e7Է{x
�0������Z�f뇯��*ÜT��w˔1=kiu��3�f�V8��q���.,��5�K]R��9�[�W�v�-������;d�ҙ�y�ӵUd���łʔ4#���T<;�j�X�2r�z��u�w1��hj�P�V���ݚ�Y�o��Wa�{XPv,gSh^�[��%pm��-$�)N���s�移)ᗲ.unk��zM
]k�w[�oēD����jaj����V�4�ɉ�HKX;�B�ޮ13�y�޺�Qa��z��%�B������S��o�(%�&�yt������s��� ��|����
�P" ����go�rs1gn���I�g**�3�rԖ��쨪:z����np׭Exܙ�`�,�ën�Q�E�;�	��<�b�pr���Evc�v��1�n�8���q��q��q�8�8�1�x��=q�q�q�q�q�q�q�x�8�8�<qƜq�qӎ8��8�8��m�q�v�6�8㎜q�q�q���=c�1�8�1�q�q냎8�8�88�8�8��ӧN�t�86�8��qƜq�qǎ8�8�8��8�8��q�q�x�8�8�<q���N�I=ï(r\�6�[ū!��eQ�yJ���KWZK�뮙Ԩ�[�l;K.q�d�tk��*XZRŨK�Ʃ�4�hѹ��Q
�JX���i��BThb{����0ip>94=��j�f}�<�J���P�����l��ƯV�S<���&��vJ�ܰX�2 �2�wh;�X�ۚM����=o"7��&�3-q�������(<@�C�ǲ��ԫ\� {maX*�K�	6���j���91s^�tʬ�x���eٺ��:R�g^�O��]�=y�#�gn+��oKbY˂���xd�O��+��Rw��&�7���$��S6�E�M�47��{Y*�Pnobnо�l�E�c�����\S���2�"
	�xGF�4�{�׶n��֝)��!T1qhJ�j���/T�61I�ç�����FU�ͧ��rr�hCyi�{�Sb�d]O��:Wt�бO�.,�ي^#t9���f�xuw)a�QՌ^�jTbm�"�^U:��o%�f_VA�
�GDum��zr��%rR��чV$��WG۔��9��q��i)����ñv����Fo,�p��b��������9+��l���ҧT���r�\��]�w�1����ǎ8����8�8��q�q�N8㏎8㍸�8�c�8�8��c��8�8���8�8���q�q�q�q�q��q�q�q�q�z�q�|q�qӎ1ƞ4㍸�8�q��q�q�t�8ێ8�>>>>8��N8�8�q�q�q�t�8ێ8�;pqƜq�qǎ8�q�qǮ8�{���{��u �$�Ã�����OokJ��{��v���*el֌O&m;Ņ�WE�ΑUR��<H7Y"���L]����E�<so��5$2���(K��Yz*��M(�b��*q��*}�>�u�
��W�V'��k��u���������ۖ��N�q�SH��2����&kRWC����7ġ�5�pۇ�4�n�m�χ�ܮF�n���u:�-�-�"����N��惩mI����w*n�X�=�`y��[g��/a���L��8aZ��IӶs�;|L�pe����/�=1�D�"�K����0�<����f!�.��qfi.fM�9v5`yPY�A��FA��X/J������i.��4n��y�+4�/.H���S7u��S]�<����ŝ�;ǬU���,�5X����ﯲs7o���6&��rtx�QU���X�X9��M]��]��ft���T���'���"[���,U���(v���[�vv����]֖��O��(�h��9@�mH����#�>:E��+���r�-�&j�X7/���F�G%Bs�US�U���S�j`�H65�7e���h>s���b8��i0�v�<F�Xg�H�������~�?Ow��;q�8�8�=pq�q�q�q�q��㍸�8�q��q�t�8��8��8㎜q�q�q�n8�N>8�8��8�n8�8��i�q�x��8�;q�q�i�pq�q�q�q�q�x�8�8��q�N�88�8�8ノ8�8��i�q�v�6�8㎜q�q�|q�qӎ8㏎8�^�n��r���*����̺Hs�r��3zEWڅl5o�uV�HA��(�numK��x�4�ɝ��5L=�˳g&�T5�ɲ�4��p��!���U����1[Z#uGb����E{r��An���e����<w�b�^�+�F�]�r#�T�pA��P��v�va5Ԩ��mʌ���F����{�\���u��."��(9�Ru�o�h��T��>��{�L4R�V��z��)_.[Q��k�k\��ª��"��_hv_`ѳ�������%���ْ:�sPY�$έ	e�n �X6�WWC�eahgj���ZHmɶ�+Wc��+Z*�T���N�0v��Z��;.�I]�D^vĂV˦)�Re�L��]yt%�v[�����`Ѫ��Vvo=�g�ge�\s����Z���x�dA*2S�Q��˾��c�^�$����`֜���1�B�SNMg��t�WїY�x�gSi�n��Gr4�٬������R��ta�o)<K�qNӦ7jeYh�mV�["�mӍ���B�*��T@s��9%�IR~>J�ԭ�z�k�i��p��Reٲ�n��K-CF��K���������y�w�r�TR�J�g�V�j�],�����������{�l�k�q��rm�Ζ��*��{l����6���gF��b)Է(s0��&�����'Z5�nz�<���+G��k7���фWM܎����D��������[ܳrj)�2m���Q66�u�^�ٚk�{�˓i�iQ���d�y��K++o��][��c�����[S�Z͔o@Qн�g���喵乎k
���ջ�8dG:���Isf��鎖Cb���V�gX�};G1�&�������'�sWV�Mwk�������֛�3W@ɯ��* k{����Ҟ>'���hM�K8ԫx�%o��۔*�k�zNQ�j��U�^��Xy��ר<.�]��%lB܂Zg>̹T\�j�c��W6Be�w\�=���j&L���A�v\� 5[U1������ͨ[�e��>]���WCo���W��b��(<D@v=C����{�\���c�c.�T��<�}��[� jFjâ�b)eh��qwȷ5����Ee�kEU�T;��XU1v��:8�w��iZ�
��Bq=���Wm%7wg����Q�].��Kj��p�����÷ݙ,K�zj�w������hn����'%�ʶ���(GW{z�*y�e��2�$[�`�Hoz��"XǙ�=��0^��>@n������W�x^�0���}�!5�m��'b�����Ür�YT���2�<�� j+���@Y۝��;#[���Ň�	CH5�q��VWj:��@kW9}��4P��\L�i~��xq�٢=�05~R�q��,�A�rse���t�F�̽�Y��݈y;ʠ�k�T������3�+��ma����
ʡQ�5zl��"���6���X�N�X�i�R�
�/zCq��$/�1B�u���r'��I�k9�Q����t�,�����PVh|��T��n8hSFC+�V.;˿�p^����ly<���W�rf��rL��ڇY���]J�AT��o�x�oU;/x��ݎ����������uwFAEK&<0c��Xff/&�]*E�C�+�}�[�U�*���[\լ����98AYJw7*�u�ڀ���>���(C��Z�1bb ���mL�=gi^U{�L�n��)����q��9[PZ��*��ۃ�0�w_�M����;y�n�@z��X� ӭ�Y�m�i�+��8�H�K��D���E�ǭ��w�o���M���x���<$Uή�� �'3���ڜ\0��Y6��k���:���P�I�B���ht�D�����;P9�Q��b�[��wr�f��w5�t��e�>΁ӵ1�NX��5US;��V�ɷp���rCp%J�gX��VD0�1���e_���o^�-�̥WڍC�"��l��Z7 �^|u8ܨu�A8��oL2[���i�l���Κ,`�p�
���寣��m�J�7OXn]�*���(�AwZ��p�Z`cS��ˏT�N�U�Z2�d�Wb��i$bõ�^�͚�<�n�W�ݥw�	#�w�`���HU��GR���*/M�6o-�Yb��,ͺ&�H��b�+-���z5�^����݂�����Ac=�h�Y�7�uʖ"�Q����xO>�{��z�����R�P1([]��UC6!�Z��츬>�ϑǶ&#����%�xr�$߲`�4.I�}#Ŗ���)�6���� j�čJ�]@ۻs�<�y9�����E��k<BËrT�YZwL���R��{�FhU飏xֵ;�ݯ@��%rB���)s$愲vH��Ux�x�f��p�V�l���c2]�y��vW*ܡ[��1B����5�]��{��B�X�SWn�O����WNꫂU��ٙ'��yr��o&r;P��K�L\w��n���|�r�a����ŚH�aÚ�!m_�M�7����$V���c��Ќ�oz�WT���1����s�K���^\y����9\X»�۹Ҹ�R���n��IN�T�HIb�WP�}[�wjU���qT~�t�����ս7���'-�.b�q���i-�Sqb�}��.���϶̓�xp�O�\ꢶ;��
"R�Y���}ˆ���j7���5��d�<g����r��GOVIiX�.T��Ǯ���]^cc`�����6^�������4p�tL�qe�C��9�ӕ-�T3�j�/'�� }1��b�E�$��#7fu��O2U�$%�6���_'R��ޭA*|>�}1nh!�{-z��]�=����RrjQw\��<�"vR����t�,�peCft���[ږ��7���f�[--�C�W�
b�J_b��v��7�����'d�:�� nFl�x���0d��h3�0n�c+GpAн/nIw�e�*]7G��Nu�	
���U�m]Dk%C��U�^��ᠲ���ÒB+6-y�nV,rٽG���6+2�)��ۧڬB��2��MAw{�;��t�
��E]�s�GN|�6Uօ�-���eYS%������U,�fu�:(x-�P�X,u���)�K��ٶ$���{<���Xĸ�����O_D(���k��#���"�fK�1�U4�2h�J���\�����cn�؆�J�6�:V:��S4o����0��ں�hkT]�ɲ^���j�r�������J�%�窱�)���@��n�ݓ��]c�Ø�H������Ƴ":�딫�*�uB����p.�c�[��R���Xf4�f��Ы9)ќKT�;q+.��ET�ܫ_ort�){GVLLgZq���ۚn��B;���[yɻk��5���f�����T�웈)��A�:	��"�������S�n;�����R�f���6��YW�xT�VSTp�(�]��7pm-�N��Z5����Bc�ķn�WNK�����+cͮ��m��"�y���VgX�����X�|h�(NY��М7vp.1u{�SC����i�Z7�>�o3�u�e���±�,��������*X�r!�Yua��Ҩm-�M#5��E�
�}"��H���L�#l�-:'c*��z�F;.D}�^�f����V�!xF�EW�5'��b:�4l�Z�nՅ퓎��g_%v�:�������T�X_jX���xM�b��)D����Va�nR����*��eb��;�j&�39�h%����.gU��J�P��qkF�WP7!&���6�j��\�mШ���қg:�-����=ϕ�wS�E��9�Ū��R���i���&gLk	qه�ț[��܀P��(<�����lm�aزV_5��=�#�7p:쏞��:��1ұ������t*V�����&��O�w���"�*4r���R����D�2�
�\�Rؕ�ΰ��Bt`��[��<&l����̺,!cYU�׶����j�J��s3���L�G�wm�f�##>Qk-WLa��_V���UZ60�y��Acr���=�V�%tK!�O]�SR�}�b�س�Ws��.4ư/b�2�S��tؑtZ�3��8���4������ݱ��l���m��a��m�Zt�8��,7b�@a!��G��B�p9Bkxj��l<���.�b�8eM^�ս�l��`�B��ι
˔[=���u��۳6��q��0���M)X^fnb��q�h��II�*]B��۠B[���˙���%�6�>s��6C��s�F���b�<-;�.Rx�����!�
Yg�4B%�$:�V��g6�Y��Ř�,�l1afh�z�^��+~n��K��ku�˾{�}ߙ���
��#�_�~_�����/����R�I'�R���%�&6$}H�h��*~J%L�Q$�P'p�`�bA�m����C��qF�)�`DB�����@d���h��F�h0DI$�) h�CH�23#)�B�H�L$)���j��PhטhN��%�qJ
4|�T���!h6Sm2J�ZNAa�&&��6?#$1�#��M��|b,�D�$"�h��D T)9 A�@�DHd��I"~H(�n|B)31�߲Yj�E��D�E6"
CM�P�0�J8�i����c%�W�Ώ���C�F?���dyLx--�o�(
��=3N�i.�r���v֚-��l^f$�D]p�CŇ
�����J����OaIt�I�]�Eu��X���ܾ�)N��A6�3��:.���.K��5zn��Q�ۧ�[4鍜�tf����ni��;ʕj��K����QY�ǘ�I�����r������#�4Z%v`��ہ�8�C���h�u�ΠUCGr�y`·6�xɼ�o^��\���1ס�{[�
�A�Yte�q��x򲺵[Y��X7�>n�L�����K՛���+d}]w�/RV7	�2Q�y���]��M%�v�(����C�r�$⁵ogiC+��Ov�)d��PU}�V�,'T5K����k���۩۷p.Y�P����lb6��v^U�	z�ܢ;��V�X69�bd�>qa�(�F1WN��M\�)�s]�.��Y؋-n��:�m<���97�kk&̂�T�M�ee�XNVqu�O��j�u}���n6���R7Zd����m��K3�����\I�Ň���ۊ�O"c���8E7�uA���'�s�N�C�;9=�#{�3��]=�n�	��/�`Lb4��$�M�J"�"�3R6�B!�"��F"Dd."�h�D!@�^�jEXb����"�@�@��H���	�"	��&Q�0K��Ќ�[m���"9F#�!��!A$#c,�4E9p�̂2��M�Y�َ4�S,�L����P��Q�L�*PJ@�M��BM�b.چ2XD�hH�RO���MB���*��4D!-� pōB�AQf�h&E0�4�q�`e̅O�	��E&�m��I��E��h2!N$$��E&��3�#n6�B6�E�T��ƂF�Sp�4M!I"�B.�D�B		�
1�&
	!1�$�E�$&�$��1��4�� ��r ��2��(2��e%$� ��� H�	�~AHPi!��I�`�lB)D\�B#?HD,6�!�"!)��@�
0����@�[0��2LNi�H(�,,��%���M�#��¡O���(^'F�EJ����;�M~��{ۃ�`�c�F��~�bG��a5U#��6�ӷC�n=}q�z����4�ӧn�5*Ho�O��1��r1{��&��X�{W?7��O���Ǯ8�8����4�ӧ�[��6$�������˒Q�J$�3/���7��i��z�8�^�|q�N�:q��#X����D[0��mˇ�$�&b1��76�GW�^�k���/.���!��o�w��ܼ�^<��y˓m�m��뢶9���ܙ]�۹�%��;�睫D�'.;������5�].I��Q�Fq��Z�ɖN]ζ��n��;��m�7�pݭ�8L��+u�u���V���N�\�5��t��f�"��ܜ�;��so�L�HAu���);;�p�ή�|y�˪���ڗ;��nx>���5�w>m�:y�u��c��e�מW�IEJ�$
�*2ݶL��K�^d.nRhLvs���v���뮎w5�;�dvr3�5�wni��h"�h�ϯ/2XY4L#|W!y����DI��F�4��@�T �}�}|����@�$��a0���؟T��@ʑ%r&A87*B���u=HV�u7t`>�Y��u��;Yi����
�����]��f0E;\g�ى���0�J�!��Ԃ(�l�i�f4��&$_#��!�b��g�L���SP$���P�
�m8؊91&�H��-&L)� %(�-��a�_��8w(���i0�jE�Fd#%Q~�̖*��=��諕�^��ע_lF��z�7�XS�-������Z
�Sa�0���N��	�I)y�-������Q�[o���˶gn1�R��A�*|�U>�4v}��kA����*���^'*0�sV�ǫd����Cc:O�͐�PjmHIVcl�W��E>�iy�+��)x�c����ȍ�!�9��c��jܳ�`��_]	�7�[��䗮n�U���|Ru�1)l��[4�$������=]%SV�0�.����fE��'�^�I�H0�NbI^ס3���/�u���ܚ����NC:D)u$�E�+UNm�v��}�|)�k�n����/C������-���5t���TQ��;iԥ�������0˨O�$q�м�O�4�jN��# =�Ȳ��ticl��8_L�����_Ay.J¦��ޏ�wd]��]cu�Z�!~���vZ/yu=�jֱY��u�/���l �(� ����m�{��X�#&�io��i����5_*�u���Z�j�g��O��{Z���w���f����¨xU+p����G��C{��j���|k"��W �U��
��,� «�4�C,��Ȓ�����5�dk�h�W�ϭ'�KCN��m��X�+�A�35����S�;�d��^��^q�4:,�h�,u�Ě6�j�CBQql"���>���m��C�'�������x���9�/s���ٷx��I\�+T�B3V�h&�dazB2�s6�6��Ѕ��{��
� r12�|zB���z%F���o�������Kd���Y�򻣠}�>q���O�����zא5lr5�Y�Urn�A!L�f�-���d?P�Ot�l|����\��\����W�IN�2m=�����@��Y������`1MK���ĭbm�(��[TUL�b��>���Y+�R�^YY4�k5'��}��%�lO���n��N]֪��i٬U��!v�R���Bj��+JEHЙ}֌8T��ς��=�	+>�&Kwg�9w>�
>�g©{�YT�3j�M=.,lkʗ4r�.���(����j�2E���dW6ojv	2�qֲnr�t��4a��Glc��U��y���J�����z+FH��-�QJYJ̲��9��2Ɍ%>h�mY����5�>з��!�uwZ+Sn���#�iy��F�rEd��wC��P��P}gy- ���Z�����En��}²yŸ<C�iq߾۲���_���7
?]-�~��=S9��L�|��ز�r���EL��C�%����J;����j�Շ������p-��Fo�����ɓ�U�	��s����5�wL-�5��Ub�h�P�'u�N��N$�G���ҹˡw݊eѬ����B���5@�g��F�C�+�%���{(@F
F@������^5�J����@�h��ѽ�� [i��7��o�+_���i�w��2�U��w�\6��"��]`E�@B��ֵ�FqX�3�+�>#T��]NdN��Nw
���v��Ɇ��P�'0<�E�[M�C��	f.���jK�չ��-�+G;�7�RJ����ξ�jSF����/%L���
��E�z���p��3f�����]G�íf�&S��K�����T�o{�wFV6�P'�`��P����v�QP�7�c��徾���CmetS9�L�j�
3����y�¤d�oM������`{Cw(O�O���'��>C����k@�Qq�f@�M�+e*��UTZ�h�lYU�ᵰ���1ӧp�R1C�	l�����>Wd��r�Uշ�fDK�(vl�/y֏�~���F+޳�s�C�h�8�+uC�kQ��kbn����-�-f�ul�\�T�s->�_Rz%��R�SL�&�*]$�����Ơ�:�V줯=P��'ϵ��c����r��_Byf�a1�X��E1@JԳOjϽ�<cp�?Z��R�q#��J�9�Jj�ol:}+cQ��BБ7H�|Ʊ�R�ʷX���b��/Ic�QH55Hܫ���{زV{E��G��3�
a�E����[��Yi�aT-!*��cl�2�4�cc�ϊH9Sg}����5Y9sV�\X�����#���L�rM]Y���k�1�^ʴ�y��87�^Kp1$��c�gv�P���Ƀܰ����������`�Q�:F�l�/��1��Dw8;i=SiАfJ[�т�p,ƸHѤpH9��},�0�+%N��z�Ѧ���G���9��$�)rk-�	Ӏ����m�{�h�a���|��\��~W���el�Q��#S�/��F����-��g.�י�L�-�eH�s��r.�ঠ��N�jܡL���6�"h%B�ˢ�}��<�`=�F�m�֠rI\�}�8e��{��Rf��q��~mCK:m�����5DcY�a.�w�f���(�A�.b��AN,��I�i	,��N}4]�o��ņ�r}�����#� ׵^�N��ڌ�,�rq�t0�3��&i��>��Η
�L?*�p�1X���KLۘ�:V�B�ǺH��|[J`n��oO�����7s�⭧����F�lה�՟9�/�o�c�l�Cm �rF�[�Nh�XMTY�7��;癯����o���i;�29k����1���_��E��
�?(&�C.�!:3��#"Z2�fw�J2꣫+���'��>���u�Z���g�G���`s��Je:yy\k(L�(�R���
gh�&�57t
��.��of��)dޫ����bX���f#|:Q�xy��o6=�;�6��I4gd6� ²�
J��&;LVșFwB�����cZ�
�D�֒�J�@2մ�0��Z�\�w�>�"�65͝ ��_xwƬr�y!�D��i�[�����I�U�Kf=�O�)��B����zD(.����1��_���xE}�!�%7�k1����/�T�ry=��������?g�p��r�S�ȝK$�ul	CǗ�́��~K�� =����Eܶ�5�ߏ�)�Wi(|*��P�}��}���|{�y����e��w)�����4G$3�c9�]���1���\�(�Dkg^\�n,�M��X��"�3���>i������Zd"@�T�X�X�;D�x�v�\����aϴf���@+��'Q��+נ�yS�j�6�ҽ˩33W-��k
Fj�w�.�W�o��y)�x�h�_Q�������>�F�wd�'��,j���DD���/��hbŢ�����V�=ԕL�P��Ŝ-w9ڶX�R�]1v�Gt-��[�xU� ��8*�w&�h����i�i&1��
#�7�Y�<�Ͼ����X��U+��( 5nXY��K��Cb����1P+�`{�g�3#;פ�w>b�"I�P��ϖpe�Lޢ���VQ���
��c�l�7��b�z֍��]�e�!���¸���r�
<��U���f��a�2}����>3ZBo�KL��(a��m�(��>��[� �.�[Q�#5�X����L��mI^r���wXz�}�L�)-�o�ɠ�i}E��Y%,ې���Z��x���d�G��#A:���k��6;1"	JI)`v
�*s�}x��*e�"5mN�=��a��Bx2�d��E겞kk3���Vߢ{�������Ձ���uc H�56K��u+dӝ� ��RѬ� 39_�E� ���N��2�9���Zʓ�_o���{��iʇMov
4�(]�[X�2���Sp��Mq�>x}ǈ�T��k��;�s���{y��\��slgi�������X��ͻ�(6�â���{��1m_��F��F�u�����rglݓ����@!��6���77��˟-?k�ʫ��[�[���桝"g\h����lxj^��7Os� c�M�YN�-Y!�n O���Z��!l������Ro�X!��O�*q���,.��Lӂ��
4Џi�S���O��=��ʐ}U>�	Zr�-����b��f�3��ǅ�F��m��x�k6�J|��bo�A��eG��Ͼ�X���[����D'��dskn0Z�|��6�Y����:�#�O���H> �G/�����9^��)Z�/
����^dmKm�Y��ؽ����)��&�bp�q�}�����+J��;�*�YB�H�H�A�V%�Z�����5}�+�z�7�#Rwr�(�V٤i� ���v��o7o>r�ST¸|%'�߁ؑC��l�YL�ܔ��Ӥu�C�p�wrE(�����ۘ�^՝�N$yn%q	�X�������솮��4�����Vm��H9�=j�E�v�qXM䃷E�ִ���\J�:��}���q�����x�[֧=֗t����b;��_Z�޼5z��]�ֺ3_E76u��X����A�$1��wy,�J:0�ZFӏi���AU�Aen��KV�@m �<���^l����WUE��8q,�{�K�v���M+'wwĶϒ����_���8����z��*�63^w��j��^��wM�	n�$`,j�3f�r��a��x1:2,�H@A����Q�;Q{a0+,�f�/ȭ�+e���,0�cjg���j�햰$��a�V��5�a��2|�u��K�j�#\�X�4<!�:}"��%��:��t+n���1
�d��Le�j�L����>l@&�h^�k-t��ea��f'�є���b�Q4Sۜ��p޾}���5���
�4�K���<������f�����}𿐌��"{u�·��lF��X�����S�Rڔ�Ov���'�^UlZ��)I77Kq�y�f-X��qo��]aQ�za��Y��B�[�K7e��V�.+Lܬ�u��l|�Ɋз�]�ܛڋuU�>��j�)2��W��'�%J���/�7ujg��a�%Kf����ή;�����U���K�s�W���|]��cIyW�e��9)lTו/t�k��gԁ��J�ڇ�Y��{]��)=��\��U7h�@��T��SK�5,�d[P�r���]�5�5N��a��0Y휏%JS����R͆i�ج�+qqSk2�e!��$aO����⋒��J����L�U4�:͜Q$�f�	쩢Zh��3��7���9U�|��O����ُ��	�gAخ����gω�9�X�v�p���H�e>�O���[v�c6Uw/��>}mer��s��o�č��O��%�d��m�*2��5�Wm�A���3�2<+=S;s茏>d�>���b��Z�e�^Ka{)6>{b̦�){Jj���n�ϵ�ܬE��e���F� ڙ��a&�b�����[[�tqa�����^;��c�Pk�a�qf��TnP�`�qڭ���.��U�"��UΠ�\�U���JM���f�َ�.�}�cy�֬A�p�r�򮐻�ځ��~=1��1N�N�ǩ�J�Esܾ��;i�h��v��襳[���`	s�ޖ��$�Ť^�5�i>�^G������[��0��!��{.�jԠ�hN�%m=��m\US4ڬe�c��^�T����gm��e)��Φy���D��U�Ts[,�ݚA_��h��m���Q����r��7��]fǁ�;Q�]�M�b!��㭾<�2�ɏ3�p'��!���smu�}�-bغR������,�\�x��\R�F$�kT%�7"ͬ���cz���e����{p���-�y�R�L]\���7�8[�W��x��6-�$Y$���N��-�:fM*D.�Ի.�\�lA��d����cvvҌң*>��|)|�
ʢC}y3���ۮ���\k1��mv�h%כ�K��;tR��+}!YZ]b�9kT�kjq�{-���c��J���V��E+�T���s��R>°����"P���e�oZ{�{�3�Ֆks���޼!��V���z�����S���Ֆ��Ev��>��7�erNܔk7z^݃iWR��ʠ��6��-����)���kPB��we�����Hqq�Nͦ�O:ii\}n��ųks����׃x9ť之����9��sr:�6�r�H;f\�)y��U;����8�ɉ�����p��-;k�e���^1]m�nUZ��0p��k0��+rǑ�O�������]��F�y}Tf�LD	E�Q����#���s�b�`κ<�v�q���"s&rX�_
�z�.���}���oc&�7{��z�*�\$t���B��z"An��Z:��o/PG�i_U�,нR��c�I���YӷR�\��8vI��9M�M�8;0���E�ݎ��.���M��l��.kOWdXR�tD�Uz�ڹ��'Tx�q3r���-gl�ǘ�=ԕL�"�N�a/��<��bYU�����#��[�F�΃pv'�����C,����7j)H*�K���;�D��d��d�|��з���^�݉�1j��Y���y�%Xܬ\�y��;e��Yy�E�y{�Q��"L�>�w݊]����!����]�{�Uܳ��%�Ս��o4��{�sW)s���tv¯kK�pt�K.�Pum��p�mW�Zk��Cevtw��:=����4�Kü�ͭ��u^,x8��VKYW0\��]7U�ӆPq*�����h��A���챑L2Pbi���F&dd		�9S�:vǏ���8��Ǐ��}v۷n�_o��BIE�Ҙ�64Fc�up��F�\"~���������o���q��x�����n��}y�$	$�ID�_n"��<PіH�"��@��$	$��#�����N�4���8��Ǐ���ݶ����j!#	$$!	�� 3M�v��ۂQe�w1�]�&��J2b��,�h�S"(�%��F&Tk	!�tC���$24b(3ޮO��"�Fd�B&|WDXl�h,`K�ۺW�s ȘC����&0F7�]0W��)�;����s�#}��'��$�)�7ӳ�]/\؍	�"&���[ė�e��b�4gήb�B�LM���/�qx�!$� �!�;��w�P)uܪ�&e�e��`��j_R�yR锘�ȻSv*�rrwإ��
O%��ܮT]T��44��M�kgy��l�kz���6�m�����)�# 7�kЮ|g��D1��QϠ
��uK��|��l<=�����.tP�i|ou��b�5��2`0����޿����t��K),����e�a�x ��$�� tqL����}|�ib����R�}�7�َS��Ч�eݡo��s���_�!�\�DN�
�>��b��R����SH)�=���S�Ć)��f;�t��B ��Y�����/� D@3��s�?#}TՓ�9�'�ޡ����7�M���y�n_�@�F�5�=á�����1i[�2n��!�s��=8~e� �_>J��۟	�[U�V�ڊg:�7�<<`8���G}��L�7�I��dS��o��v����v�y���v��AH�]PL�������xu�c�Ft����s� ��/h_U�֣�.��v������*�vh�o� =a)[4��d=��w������~5�{��|}�y߳�.`f�j�-C\QN�
����8�{_]D�!_r�l�*�{��Y#;�YA�	*�� a<�\��d5xni���	�d<�<]/ o��!�tέi�h[6�n��XnSN��X?���y�cO��_@��\�H?e�{b�lwTi�`?����[���cW9;dsd_89Ѓcm���\E;���$t�@��
kDoD7�4Q[��>{���<�����<�����IZ:��C-��S��8n�|1&�0�ldLjg�{l2����,|�|��۫��ͦ���<�m��:��Q�%�um�C `��0hp��!Ia�z���`���wL�[�&��p��� 3�7SS�TIf�������5���>,}��1�Z����hndzj�}�.����I=�{�v6��.-t�)�z͕�Ḍ�e}�"wD�������A�	��{3���p�������fjEݻ�{>ۜ�����[T�k6����+p(�-�
S
&^m�]���G�j� �G��.陏
��5Z�����4xv���E�^ׄ���~�z�:5w��������t	�x��t_��H���aг�7L���X9D>b�>��<;��Ѫ��CBͻ�⣇���G�t���W�0{�@�\?3�k��/o|k�O���#�䲈�����U+���cuC�פ����>�}�׶Ɣ=7$�oc*��F��.7�2�e��{ɰ�xCw�G��+``C*{�r��]���XSW�q���~��p`�~��۳�ֲ�۫�ζ���m��oTm�����8��I��!M��1S��������[P��P���w������Y �.	����r��7�p��N��ov��F��2��#����I8�j�}}jK�v��a��[�{��x�.����e����� ���(wopG߆��/��}�n���Y������]ή�	�AhT���߽� �����z���ԝc� ��Jkkne�4`
�����t�8����z|y�oW��>K������.�����q̙��/l�F�����)�����-�n���� n�9l��<�xL8���yI3漽��r�� �|�b������M�.z�4wB���z�]=CV�k�5���;��2ފm�9˫ʽj��T�czEE�e�>���mx��_O��ŁS;mGM��J�٤�v�u�a .��<�a8��a���5}�+������Hf�i�!x������[��>�}��|t�p&ґ"�Ⓓ�1a}�Swg[���_{�:u.5�j/g�SZ;V�vvk��%fM}1�D?��:�T{b�W�X=H
qK َp(wA9�c�S	�=��,�b�N�?eS�E���.4�|	%��P��"	�h^�|�k����gr�i)1qAdxTu=}ֵ��2��W��o��
�I%r�6p�@�JNu��q�� c�=<��Q����������Yj�,���� 
c$��I.קX������vŰNu@��}���z��~}o
��66%ڽ�4!��u�����G{i?�"G�4{C|W� =��2L4fZ��S]����#;V��v�I M^�����kG�����ٙ:Q�#�X��ҳ�ƒ��˚�5�{9w&9���o)N9y��t���`��0<��_/����/���Ht����ޫ�6O�����uS��Q�nR"D��
���u.h���Ȏ����8����H�\��kǂ�D�� φ�Qz�lh��$�ˏ��nq?/��f�������P-���櫶�+��q?�����X瞂�H��u�3VC�����3Z��X�w��F��=�����ܠhq�T r���B9�}�W�7X�ʏ5c�nQ�S��W\������V��������+,��[Xu�ՍbK\���t��&�6��c2}z�ډ�qXz����i������=���\~̊��;��L5v�Vk��P�E�@��?�!K(mɧ�4W�FX��Z��f�&g2p1�o��2os^tSouͰ�љ1�B����+��9��"sY[�o2�	^��b���� i������6��ulh_M�w�ڲ:��>*�}G�����ꓩ/1���k`{��s�,��<º�� \��_=���;d�-`O@v�Nry�d�M��˼C���w���c��=�ֶv��-�cܜE%�y���}���f �Яy_)�OB֎f.���5w62ҷ�ۤ#����r�:�MK��N(5-�omȟ߮�MŖ�Ws++9I3��A�_�7_{i���eu��fB���E��v��[�7_+�����;����k��6���r%��\�ߗ�?F1��`��y�y�L��~Xa�Z�P��G��OO�6�sn�9/�B{��1�櫫ۚ���kn���=���a��4φW�6���X]a��S,��ǑC�>l��u��oQ�ne��Hw�hu^u�9�i��%ׇ�<,~��,�ߑ�����Z^)Í��~���4��� CW<����.���t�Vwxk��
<H��<����^�5ֿp�l�Q���⎭�"�a:a�8¸��3�%�k/,���ZPm�S���`_x���W^������,���@w��0=�#:�(��kF�ȅ�V��҇�4��#$G���������J�e�B�-�i�"�M��P�_����Ӿ���`O��֙�L���W<�~^6_Cg�|�ib]��������G�e�k���I��!��~$H�����+UƊ��(��v��k|�Jc�_J�G �`���*�ԟy��ݹNT?x�[L��V��_s�I�{�
<�ܬ"ySl�I_U Ր��H(�F3�N�ó�r96�"ej�.�E0���I���Id�'��e{�w�[L�7�ay�;���R��s˶�&;6��koY���������*V�͸��(��c�V�9ǻ����9�}9eV�od�.��*�/�5�q��U�^Q~��r�S�W��q�[�饎kqk@��}���`b����Ir3Sy�Ť��7�o�&�1�1��I$�1���ey��x4���	�����#^M8>�cﳢ�����M��]�k�����6(�_J˷���gp���>�m�0��K�5��͓q�3�<LxDtv?wC{�+��{W�l5��`�o�N+�ݎWx	U4�.�n�ӏ��~�o
I�Н��ېf��A/3�1�Y�|����q�Ë��eD_�����O���ڮ�3r��K����~�`a���d�h������zE����n���(�x�I��ח�:9}�,AK�RG�<��5��5���s T��'=$�{58��J7p��~��5���\�`)��w#@&���~��j{5bA>~K���|�
�1�U��ۉ���[��	8qw���|*�Ia�ru����JKJ�{q�C�>Ȉ�f�M:g~�2�*Ҡk��6�7y�-�\&�'��|�S�mws�һ�Ƶ��O�lt�`]�&��|[]�����s{���D��ϕ�������q����7_A�T(����Jq���^����ƶ��$=Z�/��&�+��6b���¯����+��x�Tg�D�ø/��uY���ھ�x��ѣɛ"��g�vN����(y:G��Nu�.'�}�H�nu�u�]�v�&�8���2u��]�����{�Y72>���C�l��'���	-�!Ah\xm�k���n���.��o{��k2N}I��1���h��T �/��n����~n����^�rw�;�s9Ƚ���=ܣ]�k�aPV�;� �9qq/��cA���+���j�D���oᅮv��G���#����]9�m�9(��!���,ǣ½���@7��z����S^���s�^*
��p*�u��<&ˎ�}ڽk�K�;U8��o����F��}(���@�k�u�K}�;>� ���U졄�G�l�޷�9��"���ц�D��z�Ra�E��覝|o3t<�q>�Id�Nv�0����p9���Pw��;�Wx�V�M؊����^8��ǩ��>� ~��x�m���1\��s��Osq�q��{��}�1�=���_��@�?<�����P�X�� t�=�~�<�Og�yR�)9���~����5c���������Vq(A>dfw�R��u<xc��&�gLq�k��!���su�tM����5���mT��XT���^<04�QE�� .��w��#�C�`\4�a�R�>����W��#L�b�t}u����4;������\6����Yi��m�F���[ z`So3װ�+�
��B�()�%]�k�7v��@,;���v�M^�a8����|��6���2�Y��})�Z3.n�ֲ����+훤�uZ��A}[�]�u1֙��Z!U��)�Q������tξ� �gKҺ�GyZ*tC'y�s�wkU�pZօ�aw2�Z�r�P��{0�I:�%���ǖn�ݛ���u�Z�5�ߙ�<�*=��o��x�0^��q1��p��_u�� �U��=��[ņX���7��-WU��,&�� �� Kp�'���h?@dמuP�yW�峮v�o�zE�	N�@Z��q�+�����==�\����O���Đ �:>5β
?l`��a0q������:خ�i��j����J���d�;��Z��yzSN����*C1�͝Q���gޯ�kά,#�Vq�(�O�+�^�Tba����҆��f�]�x�걻TI40����N��Z��8@mv�<��}^���k�.ȯ �q�K�W�2�& �RS�þ@p��Є��9�l���|�?a��{���эST��Зx	�l�����zj-\^G��M�f�S�v9�e����F��p�{�W=�cG3)"Gx�Á�� whq��<��g�yH���聳�>�"9��H��7N�n�i����%�aˣߟ ]1�_�:�ƾ�M5z������⯖�p�A�O1�Ap}���(�3�m�U����پ�&_�mp7TKj�}z~����s(^e��@�Qw��*�G�<r"�6T�n�.���c6TSZ��w���m�եe���@/��^��ޘ`����vn�Y7/�s���<�֎m��<��e��Q6��U��xm��4�,C�l�(��"�[}|)K�dX;EH( ���һ�f�/gJ���<�'+5�eO<�5���@>�cBi�*�4*��AO�_�3��������;9��p�گ���Nip����ڣ��E� '}��$�Y�/ ���}U4ٓ<Dӛz�mxa--�=K'�x��S��(v��2[����E��3���Rq6�j�q�
��mv<�:��ם���G�Ϣm^O�l3�����*��/�۹�,dwJ��}GB�h����xCt(�ǌ;��h�� [�����7�y]��;v�;s��U�<�� �4��K�d���0�!D��έ?'����s�O�?��#o�6��EG(Nx�h_�Y�mcc�F�ML�T��� Å
;ݱ������+��x�}��O�z�)���(p�]�c�yW*s��ys|=�	7ϱ��P[;#[z��vj��z���>\�}cQY�G�����.룍�<�a����Ħ�}���{P��p�}�4ǩ�DI^�� ���M!������<��y*M�g=��۞��.O�"�1茶>��x����6|2�Yᯆ6������R��"�y��Q�X�F&�I��C�c�F���c���L�qO�ӌ͋.G�e)M���A"I�I����k4���F�~VTm��_A3X@:�;��?%;�@>}+���4[���M:��)wk�_j�q!��Z�OH��7bW� �of�}��=)a}O����1sf���������޻�k�,�~�~�ƒ�� F��Jhh��� # ����{�{3�w�<��o�/qD�ę����f�c��S>�� �\��]ðVUx[�Q�� �1�)a-�؆�̖a�Q��qyn�	�A�bb�XQ�ߺ��O�=QL	���:ak=t��'L������P��$�fNS�Y��a'��"|^�_U��]���ii�s�,o{���6��<�_÷��m�74�q�Kr󵥵M���^���7(�{��:�*��x����P�M7��a����k��Sx�p�غ)=g�UkK*�jk�0�9��W��{����W4x/4yw�m���7"؆�5Ӎ�\专=<��d�vׅ��y*�WC�ͳ�w���x%�0��׭Oj��@l�������?��z��٠�5˨���g���{��Vș^��:�3�&�n�pU{b���.O���>�oA�L�>U�숑�t}T��D�i�+�^3�|�����$�u�or�#f1�-L��s�z'wb�Z����o�J#�s��;UT�XW�"-�=�bO&j��������u{��ߜ�k�NwV��r�+�\��_䚳�lȎS�ho�77lיʡ�0u�^u:��k���F��0B��8���κ����lX8
�J��UI	�h��c3:��{w;-.����c,m.�K�T���^_R��0��3���3v^�N�U�X-�'WA����VN�������1ǽ���6�§p�ٛ�A�4q�vQ���,�[C��^!FW)R��{K�'V�/h9Z�7��{��xqt܉���k��J)��S��qa�7�=�n�#����8�kLQYC��s����nbڍ�B�v��i�fp4������zs5��{��@�*�" �)ɺ�\�+U2�7�c��b���&k#M��!��o*7�l0<Ld����ن�����\�L��.y��8�ac��յ�r�J���+�3�����w��g7��g]�ٝR��C.��Rɕt�A�v��1����B��xi�r�(
1*{�I�3#����i^�]��d��N[�o8sQ����{�L;�غ����'7F=4�*�� t�e+=��7l�v��C�>��,�Msŕ4�h��-��T�nU����N����̨P�ʭ=�(�:���܊^<W\�ƺ�݅�*\��me�:���ƕe�w��&G*w���"���rLDcY�v�r�c��9�.ڢu�Z'�,�en��4b;I��-XXo 0+�oW:�b;�D
�/� +��;[��Bi����B�UT��J�"���\t�+K*p��-�dD3T82�,��j"@@�$~��	d�*c�H�(��E�m��qH�^�7��3�5�]>���T�t���W�l�r��@77
wީWõt��H� ��7�l���ʒ\�Y�7��za�s�j�Z{	'/X�X{q��ٜ�A/�zu�ܬ	��v�5o5r7Kv�>���2�x;]莗w���,%�H!f�Y��;��S�%a%WRB�R�j苛�'b'mM�$;2�)*CW�hJ�ѵs��y��/[����/j]rO��!�y>�D_��q�B��Iv�aq�B;�PWKRbm�<zM=/.�!x^t5B�.pp��m�L���ۄ�3���KܒgJlqA�襼rc�o+��9}WH�ۏF�Wg�)Yڸ��Ә�f����eb�d�yE��0�#���rY٧{+ �Yp���{���xɵ�u}�ƻ��_/�2��z�y�]6�e��1�vWq�w�=��h��^7�L��J�s:���Oi%�tNE�1v���ܦyj��G�k���\�μ�LC� �^�fwi�{V8d�@�ִȣ;�����f<��4����M��o��`˝����_A���j�%�4���U�,�e��De*�v�{�鳴�wg�V3fm��	A:��
��Cr��	<��,�<�^���;���tN��4�hV���i���Z��3�ī�]�s��"p�ȯ�����MG�������*wy!x�����@P�M�!DEB �$!�I촒$������N޴㏯���^�x�����nݾ�6č���E���\�	R�_K�LiݺQ���$z���ӧ����___\z�㏯�ݻ|v�����FE��	�RKO�[�+��N똫��K������J����=�����N޸ۏ�����8�ׯ��ݻ|v���F�s�J�œ�_θ\��ۑi(���̌cRF�Q�31P`4�(ň�Y1g�k|xM����+r�^H�J�\#22~���,�LE��o�R�>�pھ��;���dϷQ�ѱ�[���d����ƼU⻷X�5\�B(���u�盚5$ZM�&b���6�X��7wj1�E��* �ӕƠ$�\���\��M�r�N5 �����7�ѥQ�$�##���AH�E$�?�&��D+����uε�α�f��=��.�M��{��u��׍�AN�3/Uqd%��#�~yղ�$V0�f�S��M'&2�i�S��1#	B~���F7�16�? JQ�P��Q�e���\n#�2�L��I��"�L�D#	P��T-��#O�C?O����+r�M����n�kV�d�"�"H����d���~|���.��o'Xѩbų�����;��ٍ��j��ig��������SqX�X�����^o&�w�>�JKHŮ&1ǪC�>�>�cb�G-���a>X �,7�z~���tG��c� �a3�2���DeJ�5��KrN1�jI̋���� �~vz}KV�Ey7;�
z�4.<���̋�c�`�
�e\^)g�e`-}��xw��H"���O+�Ny}����>>j�!�t�\3[�G��w:L�3��qꖙFg�e�w��Oh��j~�������鯺������v�'��:�"����<�����k�Gw������:�cP�O�'����0{�@���Q{WƼ��`
��cuu������@3:�]�����ҋ�Vt��+0!�Q���T�8�0㪥������_t%w�%����
����ި��Taύ���s�2j������uƱ�2��ٵ���:�un�#��A��E"GA�x�������ϾVF���MV��^�f+��V�F{S
�x���Q�j�Eۊ�ݧa7��M>���ռxc\�>&�gN-a��<&_w�uM�/��S�ݗ�A��K��r5_+}[%m�\�Z��:7%hU��%[�L|7�UWe�ނ�^�B��W�"CЏw�ã|���rRھ�˘����	�x<\�ʍ�`���sX:V��=���d�pP+7C�s��^7��44�4�� @���0 z�N�g*{���|�q�W�b�~��o�;�<w��!WB��<0�C6Ϯ;"��*�W��h��lN���0x0伲���ƹU�s���iYg����e�>�?X�7{��{��~O���ƩL$R���U<�{����#��3��{x)�"���j}W�v:�	�xS�Tb��R-9N��a��Sw'�ñ屒�R�m4	�I�{�ؗ�hY/�O��
��F�t�_o��+z
�v�����Bo&ƽo���b%Ih�?<���G��s���5���	�u�UH���[��������`��2j��v��AhL)�!�3�J�\+�a����|H[҇��ׄ p��K.|���bcܼ�~���;Y��qܯ�6YSm�%G��N�\ߦ6b��;��~�_S���8Kweؓ���n�<ix����/ӆ��q_I&��>y�4�WX��-ޘ��}�G\Ƿ1��uz���ůbЅ5=�(NG?FC�8�Pծ����_�t���L�� ~�t�����4:��
�)�>S��%��Yc)�s�A<�1t(tY1�����ߎ��G$S>�i�4`I�|A���ߗ�a���s5��}�L*Y�[�&n�>��[����whm��D>y�F�Uŧ�;Z/u�i;�o1Ŧn�Ѿ���w �'s�aR��J���ii��)��iX(,��l�����&�TUHQ�F�G���="5���߮s��!ݶ!uq��>�!��"_�[�7���C:;n��y�o�+h.�FG�4y�3�+Ɗ��}������l�_"5��sW���L�Ϊ���V`��t����11[�Ac����tx���k�S�X>����>���nL�Gzφ#��>�gk����W=��ԴO�D��*6P:�|��	Y~�v�5�L�) |����,��X��h����Xz��Ռpv�f���d��a�۩�_�>B=Ɵ�uh����9�KcSӗ��~�����/�����;%���_�)�R�c/�[K���0[ޭ#����3������nhɐ�<\�9����9`5�:So�+q{�0<78/��Ň�Ma��-�	��Q��/�g�{`W�K��,�P�K�'O߶l�ٟ4�<qqG	��qɱw����8�1jOf"c`l��X�D8ߎmԇ �!˵�,k�U�u�t���̃ocr�
zo�,�3�0#��9X�8��c��ޠ�x��gV|�O�t��H���'��v����T�%l����dgZ������.�V�'R�K�H��"�\��Zҕ�CYD�m��\T6����v�eҜ�6�+�ч����`����B;9vߓ3y�f_��ʝ�'L��>�W���"�CH+M �QQP�>{�Ϝ���v47Юi��ru��e{=s����D�<; ��	af��ܱX���Ժ2�>��r�/̹�c�;�f�)���Ϭ��a[��f�Zà�,�t��?X&��gt���f/�;&:'���ѭ�fA��66��|�o�kҥ7�䒺�y�&��0�n��ú!�e�l�Ř'�i����C�����3+瞸9X�����ɸ[ݽ��B���
Y�	}7�+]F~�@j�a%QW��<�g�;;�-���bm�҈�c]�n�����}�BE�=�P.����g˞��b<B�<�5��,�8GO.��.�h�z�K�^�g�������8O���u���܄O+m�
J����k��xn.1��9!����}耹��P4��Z�:g�n���ʣ�=�$�m3�󃶡�>;8�Wx�����F�rWP�`�g� �/���ߢߢ���ߨ[j�z�Ʀ�][1t$7k�ݷ<_�:��^��J|3��-�3g��y?24_n�{�)@M1v!f�54�[��{v����)�䓅��G�h���+��Asn<͑M�ҁ�$��^8�(�*�\�n��]�Eھ�|rޮ�ze���iԗ�LxN�\x����9��ԧX�%SD=�]K��=���������	P�"����}�/���=��wS|���OT��a(�»zZ�t2e��k2�M���g�o���������g��c]>�:���r�RXN����t��Ŋ�"Wt/8�n	ky.����_�k�r	��(#��o�O<1��g��{����<�^oFf��{v��ot�[R��e{�v6<9C��,"1+k�Y6�_�������FƝk�&~�2]�,w=�����7�%��=03���w)��w)M��~�`�vo뼑 �\[�9M"=��II���ׂ�ЅKڽ������t�Pޒ�+�'Z9�,���R[�����{Ɵ�ź�Vm3x��umÔ����+��2�nh`{b�y�j�����FE4��g]�'K�����Y�$�5=��>��~$9䉺+~G���:�l.��Jo:�6���9�58k��a���Ó�^�}#���d�p��Z�q��]�<Ϛ��\����� ��i����KU7�f�-�jp�߼֙>���C�c����y��--,��;�	�C���Ժ�6.�iT�O���*��=�I_u����{�@�\k�ܟ;�N�E��#����-��+j��=�U��Nا�N�TcYk��o*�j:�5��;�u���5�j�5�ra_���DeCٔxK������,�]M�"���:��ve�!��]G3]�ޛ���[�k��@-�QB�T�E5��w�u_=���_9Z+[�f�������Qy��{Y�C�붖��A^g�,�����ú\뵞o�̟
���د�[J
TC�}j�����m�K}�/a��-�&_��LY�p 0{�]�׻�눹�;+��}��~}�Ƙa<���ݮa��ｽ�Q����9�۔7�.��&݄�ñ�x��0�-�8>��f�WF2b��/�>�66�L���n>^�>a�ٷb��2���z��qM>���M��/xZiM�t)����5&��8f�L ���B�q6�^p.��WcnT�dn�ʺU��f������bI��M�$q���^��_�=eH}Q�3į]; S�uS�loI;^���砷�k]-����I���/6�4/g�B�A��C�5KS���9z�8�����P��X���5�ǵ��
>��H�}�h|u��}�';�v?����H�.q�b���z;c]�l��~��;��,�+ϒ��(�E�^:G�J|u�BG�U>��O���/o��~�T'�]R�k��GT|!�L�;����F��u��FکN�ӏf���&e#t�SY���*�J'��J�c3�f7/�WI��}{p[u�"�Ά���e=1M�����tś��\��o����.v�w7U�!>�}�$~��J�EJhiF��"�Ƭ7�_��;`��<�N(1��},���D�C	"�iD�!�������¾��Ȥ[���kK�a��>6����i�U:��#;@k�4q��H���T�P�ӥ�۾X_��^�O�+;x�xn&3V��Y<��OTe�(�]u-`i�;�3�W=��1z����B1��٭���vg�>�Λ w��"���%G;��.lH�=�U��C73J}ib%?�-#�o�Ê��>�����şBhi�� �q���7�l�K�;l��ؗ��|'���O{}�Ȟ�F���L����+�G֪��ϭ���>�XxL��4�zf��g�rk9 ���(V=�qA��jT����'|����5~`�y���M��8��S�nQ�M^F��p��}X~�z��s�~�6������Wj%FɓX���u�2���K�gg~�p{��
0���	�Y�\�9�G+�{�xE�	�Ls
�Qo�~;*h�O_e�p�u�HT"�4��j���\�}~a=1�t�:���S�y��_ZH�ʿɃ�g��8<�P�ݮY�[�cT��C�������sE�bU;ﳑ%uF�}yֱ�D��i��$�\M6�e��C-��[F�����;Lb���˱*�se2�����N�k�/	yc]Ӟ��[�wkyP.����=���w*OUGO�����B��"��y�9������j��Qɨ
�`M���^9υ����A��j���U�^X`~6��+eV�j��]M�7�q�\���D?��L�v��xe>��-��+�1:�wK1a��-�^���<f4�@o��o��P���g��e'�p���<��o�;b�9�v�o��Y=�u7���S��e����
=��i�q�ч��dV0N0A`���G����"-̷�4���T}�Pѧ�4`c��QoN4u��j��[�ޥ͐s�"
�˸1�mV�[�9W���NS��Q9�A�ru�0���+���r�Y���q#/��l������^:��[�M����䎦����y󫇇��4�A�1�6�y�}	$`YN��c��{��;�^�I���m���^���87_�����L��4|��4�9��N&���;0��@�,>kT�p^b9�ip�L��S�;�8��L=�|�bs����<o*�0�|���jD����@�,�jw���^Z�O��s�MAa
.��>edy_7������5n������c7G��������w�<}��]W0�3�n�d�N��V2���`�V�r-P��*4qܱ�n;��;�r*�E���j�p�2�.���u�D\��]vnkXg��J�W�^�����4�TD�4�ҕ@ ��¼=^��]ҕ�>�%������=]�y�l��o����w"��h�0��|b�a�0��nx�S���
�k��S#|��cU%}T��q�w��ܢ�Ք)m�_�td�k������M"�,m�-Kj�o��ػ���8��Vٳםyw|}u�7fi x���KT�ƀ;N.�s]d�z��|d��=��q���Z��,Eu!�6F�&��0כ��&v�����+#��{�V�Ok�J~K�1WvR���&n�j꩙���>lY�a�AnNK���l+O�;uƳ��ƀ_�����Lr��q�!��ɸ�:a���Α�b�q�f��,{�}�O�Õx�J��/���E�)˖f�� J��w*97SCpE��)�_�v�������+¡�kþ0���K1�⼼����^�m���\Cu���<���y�w�g��Ɗl���s�x�Y��J�f�$z��Z�D~�&'�/4���`қT��z���mN,���R[j9 �&�_tC���ē��x#Չp�=`����uإSR'ې��X(��Ak3��i06����J��C���g|k�⾘�ũcȷ
����J/Y����̼��.��@a Y�#�|�&T<RꬾY�F���s!���*���9�2�7v��q�1*6�s����Mis��|����(��4PT�(�������ᕫ��Nts;��fn_J�f�1�>�YI��+:����0�kj��?)�t�k���q�]kun޿P�xV>����H�>Α:��U��v^�����u�G�|oo&��c���7��s�4p�>U�35��PJ�3�\Su(_��Q%�z������;b�i���3�k;-�����υ�7��P�jq\�<��&n��D���>h�B�G�U]�Yⵂ��B;�_q�^����#Y-O靠�B�/T�m�%9��SV7F@��#
f�;��pf�)��Qm()Q�h=jm���י�9\�e��t�ha�Q �__�^va���ڛM����r�޿����F�y��_;>(;Vo��2:-�'�7&�|;]pۑ�M�(��ۑX�vsl�?ew���i<�Oy��=0g�:�|�ut�m0������9��˕�X�~˹z�%����)��2��z%��?�Dm����{߱������0L��}�'��Sv����"�]��m*ݘrY�s�{��&]�J�U���7W�َb��,X�U�d���NWZ��y\��)w��Icpj5�����j/:�թ�Z���WYX������\�h�3Ov]��+%-�u4Re*�|[;��l��S���cݻ�0�h�T�%e��M����������i��5(��"���q,*\n�J|�R�콣���S����՝X0)z�R��k+�m7���)�P��ݚ{oxd�C)&�[�vk]t�3�j���Z�+�n���" \�u�r
Ü�6��K^�I\��q����KZ{I�o��Rle[�����ٶ��A�1t��.�5����vt֫�$���`�ޑl�ɂ���^�v�p:,�9��ْA��+
��^rCDˏ���[�E��]Rn�q�}�~��{O���V�o�/Q����*�	��˧��)uc�b�c�$�۶z�6�}C�WW#�&�f�&�ٲ��b���ΗN�(仝�X3J�G�K7�eҠ2�
����RI*��D�ۺmֺ��|.�i��-J�׾
�XgR1�YD
�0mE�.�������'E�s�2�r�\�͇����э�
�����UN�.���.��:��B֜:��kp�<��S�p��c��`k����r���91z�.�]��m3_�x�!�k�r��"fVa̹��bqI�6��I��2A������X!��H^`:��ğm�E�&P��ζ�CZ"��pe�z*�	{���갡
�����Ï(��n� ��N��^+b��<�,��=\��7}t���/^�2��HN!b'g��K��P��p���5"=�{P��o]�{����W	[��< �a����R�>�x��{�U��6���lT
{`yB�C�9�P��M�2���^)ت�;/f`Ѣ���QqQqKT��tu��I���3zQ��9ۖ��#�ړʰ�	��F��9p���Ϝ�ƫ,d�՞gym�B�4��oz��2.Ă[w�{�u�Y��0����k�U���|�zr��M&Z����&n��W�K�*�Ҹ]K�T���5V���u�f�����'�`���\�x9�e�t�.�تQl�CkNRO��-��|��m�ۂ���t��etQʋ��qe��yc�ӕh���]7qKuR2�[Ӏ�[�.ê�,��4����R�=�1;�@s՚�-�fD�tOo��&����zZ�0�衄����p�c�֦��͉��}��o{�ԍ���}֙=nekQ,VyݦE;��[����D����w	w|ӫ�/,�]�{z��+vl�M�u��꿊���F�6�NDh�m�]�6�5��6!		 �n;t�㍸�?O�8��O��ݻ|v�Pd�ID��&�W#FƂ�ȏ����];x�n8�>��__]�v��攐Y$$�5���9�ő���߯���v�>8�>��>>��v�ۧF���%UURB�P$�R�L�����dE%A�$��$!+����ж�e��W������k:��v"�Ab���|sX,X"�6��-E�\�2��KF����scb�r+�6���[�~7aD��1��ܐ���/>]�������KAE�6�E�҈�4Q_J�+x�=�6�F"���
H*���0n�畋����s�=�`ۮ���N3�M@��;Vg^7P)���8q�-��;M(�(ѓ���n�2�@~����4
SCJ44�!�2{�"ޛ)����с��}�Z�lt���<����;)�lѽ%��\�"�_��63�Ƽ7I�K_/.�ZT���'�Ӛ�����H��5�b��aC���9�1
����^�u�s��{���(s���K��C����e����P��RS�zwvZ:fN^��O�z���vl]���=�Q:������󪄏<�������ݯy�-gM�/3{��>�or���j1�d�*�������|��U bA�<�@xBo�Lֳ�K�?A���x<u�W)��t��!s��	�����z�G��0Ɓ�͉ݛ^W-���m=�r;�d��{��tfx0 v��#�3K�a³�䉘`HYo��A�f��{-�=JbZ{>�.Ř)�ᩏ��X��,q��u	���*�<B�#V��Q�nc�J�3
�Ud�<����(/{��!�U�
^�c��u�����\�ˠP��Y�z�C�t�ʸ?oB���yJ7������8���2|�;h(;��C�G~�*gY_��U{_w�z�fJt{�7��VJ7un�Aw? B���!;�N��p�8�7��L��-l�� ܑI�>\\<)������UJ`�!��bO�o�^��
�8�w��c꾂�݊�p��|�����_L�Zr�6�N���&��հ�ܚzv�����	M(� ��"�P����R�~��
"-�ov�2��|&ߎ�����RV`J͘}�S���B��_���~�$L^�b�y%�1����4�}�EỗM���]
Yr���vn.�v�.z��[W}u�Y�z����+��t������G2��,���gE��lwmk
\�;��r�6��cT7eO<'�*8;�%P,���֜r+�D�0��yO�+��<���2�S'�(L�衫K�7[_yl�Ƨ!f2����<B�/��4��0�ޞ.+�AOph�I�1S�|���n��x��}=kN�<�,w���L}��ơ&��xe>�oIoRˡxW\����h���I���+f��^z}���χ}L(Н!�P<b�\#g=��	/��Z\Jz��]�dj~���%��&Ӑ�y��y�/�|=� �`��0�{ ���dyW�n��K���}O������$��'�O�3��������F�X����bv�	��-T�l�!��d<��%T]<�*�Ƈ��&�[͟2m���&��w`ꌳ�n2��2��驋����($jN�\����kʰGy��C+G�j��.86Ҧ��,�%��]��|��#�W�X����W.qSss2��ԗ���V]R��SY��T��Zu@�ё��m�͞�=g���z���M
��ЁM  W��w�My��5��,����|�f��
�p�6d��uBL9�9���-%�4�L�i��S��X�<��������8Ş��;@N˚�o��Xq�,҅p���D�8�7҉���>��WM�>>��4�������B�؟��X��ڜW����b�^�Z�d�K	3�U�f:�`q��r�!��Syns�;��yB�s�(j�>�{	0z�
v�yV�s�11@��+��w˫����y|�λ�ɎI
C����g�W�'�}��|d�C���d�9@�^��}�yzv�׮'��"�gr�#��S�p��9璈���ˊ���`��Q,�Y;T�}�B�e��k9*�7i_<����<�{��'��[/�	�{ݒ�2P��O1Y���>��O��g�D�z���R;�8c|*K�����v���������&?Ɗ��y��A.��1�I�fwT�[��D;��{i�d&���/O�m��(�\�}�1�I�=/}��*y�<�>�q�?c�l�������F7'�΢y�H�U��e�ֆXd
���俜!�=�("*�~�^ŃV^����ۅ�C�W݋���hh����F�����*낌qpwA�n���F��*�[v��/g���-�=Xm���z]�sr�.�h��z1��n��Az*�J��;��Ԗ޼���Ѷ&�U_����Jhi�UJ ����\�&��u���}������i�D�޺r� e�Pa���zVXv�p�����1��d<�Y��B�;^�/�V@�����_K�˞nk�Swc����L������5 �.Z����$��>T��Auy<��Z�'zK��h祚��ؼ�/Uί_3���8կ�	�&�@���C�0Z�Ő�d�0�/SO 94��5�3��7.��8�TSR����p��1�A@z�����+|^z�rmM����cw���r9��r�0ٌ��栦����36�p�����2-:�]�.z�;�\�S���? ~]�^�O� �O�睞PʲI���P�8=�=ߕ�Geҭ8��8�v�W�i�����Ff�/5����RȎ;>��J�<��zOU�vO��5�5Ώ2\x��=�@ᰑ���~ju@���r*�,�� ���K��B�f�)�X�&U:��}!�p�9�iv�4<7x	7S�s�Jn��g>�|�d?y�FZ�>h��/P��ȳ��gj�Vud�a�,���B�P�h$�H�7������Q�SEoC��h|*�j���
�J��Z4N����u�<�EJ]�9k�w=��Ɏ�nZ� �Җ��*�8+��/i �m�Yd���S�w�k����\>�z�Q���i��Dt_�=�������y�h�Zi���ϫ׷���῍~�ڃ)�P;�Xc��x2*�<�r�Zф��xȜ����C���L����F���л�ٔ��Ə����N�;�;��\O*���ٵjx&�t3
q���dN�.|��?�r���׏]��'�eE=z�ĴV��yc=�~�y[���o�t:�5�.E�7s�|�<������;�jP�%L���������A�p�~w-���ۃ-|�MҐ�y��R���T�ސ�n���䃫�RC����ׅ�u�"G�D�u��Y�<��"��*�+�6��f�]��'\"��s{;��t�=���'��GX�hYϔ��a��B�|��	5���
T��W�օ��mk�f;�Kb��!����,.^���r�H�k�jٌ X���	/<�y*uD�o�����D��
�����#��٨�O�U�AD
�*��O,��3꧁��@x��з;:�us�qoY�}L4��p���E�v�)ϛLBkoRPZ�"�J T��T Eu^���ϥI�R�]��~g��l�_r$־�ŬZ����=u4�(_�c�a�D��q����Z���@o^���Feyq�9��;��V��Nᛠ���5Nfʔ�2C�pTzLĥKu܋1�׶� ꜷ�;��T���T��hV����ם��d�s�\����> �E���P���k�x^b��P5�����b��UM0����3�����Ֆ>o�g�=��zg�#���b8�z��7�]�d���^b�B����x�a�:��V0j�6�o@�F�P�ZB>�qWm��p#ܜ���UX�l��d�ۖF5ℌ�f��ϊ�dcH�	���ѣ�\�+�!����,ӵ��岯����X�=>�H�Д=��P�W��_Ƈ=�ڟo������{Z-��؋Cd��f��M��.�o0McaM5�d�^9�|��0kf�'�,]�9I�h��U謾�^fQ��-�������1�u]c����>�i����.�nǰ3��{����[��T��j��{w���ۥ�>5҇���Z
ݑ#�z�?0��bvk���9�Y�����ｲϫ}8��f@U����K��W��2!�cz;uUs�id�Uڠn[�vc�_��V�s�9m>��-6'�G���Z�ș��C�#��g��_����,�:�05�]�t�V���k��un�jPDC�4b[���<�|W�_�C�Z(�16���΂%�0,��lZ�I+�W�Kz0j��۵+�1y��ٰ��Wՠ��cx���C��s��X9C��ø���+����q�+M)M-{�N��=����W�y�3k�s��P�����Խ^b��W�o(� ���7��*w�ӹ��q�tu^�.�d���`�S�|`�9`�Km��x9�����¤	n�}"Z��m9GC����쌎��Oc\���	�1�w6�3��s������y�7����UE5x�P�L�F�οWy1|�{��iJ5�5@�k����{�B[�5��ز�?�PU����}3�:�b�g΀��>�A7�+����3o �w�9�k������г���j*Q��m���e�|:��3d�������щ���[�֑�\[cdt�a�/WY�6�ֈ�bS���n�hm���&�n��Y�F�ݦ��>��CH��-B\%�^�f�S���}��]U�Gw6r���Ֆhh�	�8����w�W����.��A�v��&d��k��)�����N�k����h�O��Z��:��|g���}[�H�=��Pw�Kʁp���N��u�*a@�)�va6��+Y�)/Ïެ��@�z9P����������}:O�}޸yY�R"��t��{�D�;�ñ*�泿u�]���
7_���4���6�˼Θ����`21��)3�鿋e�6�k3:�h�2��֠�؜�fXA��9GJ5ʻ��S�M%L�Z�5}����\Ȧу�[���+(@�^Vi|F�Ұ��ةF�\K���H�9�[��x:(X�\iWrǽ��\���wGws�K��<�����ǟ�?�y��=ۉ3-�ny�W�휇�P>�Y���H>�
�,�b��1��d k���c�W�5���������,�-���q[��f��a�B~"#�L2Y��Z�{~xF#f�;/.�����șx���lFV9N2=�+)M0���9/Kc�!��@�a�]~d�΄�8�+��5�7;2ސ� v�֡�;�S��|���H�WCl*�v����K��"u*��ꊉ�h�v�ɸk�&��{�cS
��c���i���F}l���� �C��X���eqL���٤���.Oڙ�_os�&�=�������O75��7v:���裵���^������A��z��������4z�M�����c?;^*��u��'rR~ڻ��_�C;��*�`��� ,lv��5	q�������&�N�f�\&<�s2{B�\.¨cW��*������A���64��F�z����_3ʐ��O9tr(��<v�Ǟ�Z� i�J���9O��u0ޫ�8�]�^"z�7�7�/�1G��H��]�F�	X���;��m�ǓP���s�H��E����������e�}�[C� r��s+�lN'�T�n��Z��ip�+&uN����Vm�gv�!���*�{J]Ӻ��ڗ��J��K���������M��{ӥ���k� �{5~@�ԹB�<�����g�<O@��J��s̞}�π���[:6�٩]T�
�GB=W�7�&����@����*��	����*����,��|9ƴ'9��]��x4xz%�}���%><�>��*��B�v��y_S3�.�cz�>�i��Y
F"`�qD7��gN4��KhkK��}|=�M�m�(E��*a�L�qS깧�-��_L3���{�7K��Ӕ;�P�X��F��6��G�w�
��W:����JuE�����
ؖ൝4��\b�o�3�l�*�fS��^C�h�����ά�|��E�k��L=8�Lç�Z�8	��Uͺ�|�vЬ~�20���)��q��^og��Q��Xw;$�ʸM�/�[jrA7P�wB��sϡj�g��h��05�t7u�;*���3�ޞ�nw[�bs�Gr�O�TJ�:xQ�}����}�
gg�ݍ1N]T�zB�mM��^�,<ٺu�-�U�2������Z��1ZC\O�*w�<w��O(�K�ޡ�Jo�z�Knx�yyuv�S+[Y�YV�~'����	��U�s�M:�b-���[�;ۯ�g��λW�&�巁�n�v�+���G�����Fڼ1dʝY��5��W����p���:y�1�4�/N��R�%��ͫS�j��梂���h����7]��8�#M-44��3������c&&Swb�,'�)��;�g|�Kχk�1�|� ��6���Α��&�[�Y��޼�)��xɇ������P��ja�D�ZA/��\f���r�s�Y[������鋝oN�2�Rc"�Y�AT5�yd�bv��p�*b��� ��ٓf���yкi��
k5ŴGC����QQ�tIhǯOXc{g{��*���q{�4t1"m{��@����겾9aY�+ӆ��67�iz��h���ޮ�Z�&��0T�<�<3�e�Ǥd��������G�H�^��|�������Ұ-��H�e�|�1�oe������t5S(������l�$���b���Y�{��ù��pf�|gh��z82�"��l��
��_!1�y�	��|d�W���F<].�r ��Rl��C�8�5ϻg�����	�5���[B��ι�Pj�����+�����'�@��x���-�Tl9�7{�@~�k�d���n������_���]��ˈ�Gx���q|.����h��x�v����bA��}�&f���қky�l?��xL��'�؝i��m�X@`�j�%C�dD��Y�(tTHۻ5���т��O+&68���:e������6���8[Z�YE�*\$�C)�y���mc��Vf�Ėv�&��4�q�����p2C)c��f��;*�(]%��wv!U[^K+�f�Ɠn�ɖ�ȳCñjōq�m�������JNP͠���Of�;J�a���b%+wv�Q�9\e��(���QCD�g����f�Yw���3q�w�[�3�0�7�!X#o#�U�����MD&��I��At��z��ٵ�a�M���P������B��Ŕ�恒��v�S;Y�ִ����j��<w"����]�Y_\W2P�:���7t�1��o#�"��,j����5��ѐe�xIj:����}P��w�:��%|�U�V�mZ��tW���cm �r�gP�u���7�E���Q���.ٮ1:�� ��beو��a���-B3X�WMw(RHሌ׀@�H@z�u^�!��"4�k`c2�2Ɲ����sr�:H��U|�I�f����0�ەû���\ȫ�l��z�Ř�+!Ͷd��S��ڸ��d]�UΙ�R,�	�j����X�9T�Kq&
L�D��>�Sg-��9��6�uz�D�P��ߤ�燗�ĹtY;��/��^ĖW����V�i38-=gk�md��=es��Kc%wcB}/F�N�g]2͎���8Y�,1��<˾�D�*)J�75LN�`ɉ�z��U�2�,qd8��뺾
�(�mJ�]WY��I����'[�nN��h�Rǹ��9�h͙t��-7/o1�>oR/W^fQ��x��r���)n^��wE���^ӫ���ݺA���]�:@���nfqq������	M'YWِZ֣˕f��S����՚v�Ŭ�q�c���=���ٽ2l9�׸����v��E������o�qA˾L�^T"0��Nm��a�̶�&���Zs�ފ�Xr�С�붽5�V�w�^�*j{�dh�yD��a��k����Ć�L]a�̱>ݼ�ev�o`8��M�7x�K���fj��81������l����
=���� R���/��n��bR.�T�X�W�JM��^���eЭ�.b�Y6��un���c!x7�̹{ �����g����Ǧ*�E���A�Y�;݄�uR@��R�� Wqw}�]ڡ.�j�Vvu�ĺ+ޝ����&�
��V����N���Uh���}N���V,�l�bS�RpЧ.%��5��㽥n)-�q�]�*<~ϙ� �������֐��`�6�d	I*!Q���o�:v����qǯ�8�o��ݻv��j &/��x��M�ch���\wW(��~��|߻�N�8��8���q���nݻ|�'�]C�nQ�b���j��w��+�΢*(�����Q�	���Ǎ�v��t�=}q�}q۷n��;�#"0� I$cL�W�\ŌW6�Do���7�c�n�ѧ�����mȷƹ%b�Ź����1&���b�K�]�1��m�������nW��m+�(�E��EnW4IQ&��Fư�M��cF�WJ+�WK���Y(�lk��,��Q�2@fQ��F���/�
�F�ȍ�[����܊,��b�U2�x��hьi�[�Dl%F+�lIS$1���\F}p@[�UR#E���J`��)�"I(
-�8�)Bچ��H�@���NBb� ��D�q0gG8�0㧊��u5&�m��F9��-�L]�]4n�|�T,��D�S�S�\��k��k����"��0d�	P� ��`Q�@��r6ȊH	?EL,��[m\�)W���AE��@�DH��n0�
c(�B��D#h���2�BT�
������L�$�D	�[@=yR�%����4�CAM z|�S�u�hx�J��R�	,��(mj��l�1��_��D�/�	Ce�[򾞡��#�2!g�=��S.|����a5�ȇ�'����j�a��fL
����aq%E	�Dli��]�>}� �~Q�O��:�h���S�Ƞ�[7��5jl�}��a�V��*P)�?�����H�z]�����G"�B�S�m��?Es�_�AcAt�9k��엔
A�8&#�Z�&��T/�N��0��f\�M�b���HЃ�O=y�5��1����l[|�;�߶_E5y�ĞQ{)�:Ξ����dp\�)�KH�)��;�������	ͮ�8W�VA�ܬ��|��G��@2��y8`|�F�����y5��eyڤ%:��q�����y�͜;��������w<�1lJZ�%�8lǾW���Q�\�h|I���y�x��l%_	=;_g��?�r��メM"x�פF�\��)�k��{�y�MIٷ�7��6 ��FF�}����@Y6�;I��|E�0D;�<֎��8R�s��k�#}�ʜ����aQ�V�6y'lλ�_4�T2�#��M%�:i��WC�NUE�dWf� ����$s���J�%]p��Dnˑ��wTwU�����ng�sp �tB�r����l�S���;�3�X���40�}�󜯞޽�Ԡ�h��W�V��^�!5x��Sz⁊�������<���}~#�|�;����D�?�No���ې�H�q�A�<����o!�%t��]�zz�<�ۓݡm����;W��!GϏ��JH*)�=�0�צ���{��s�aʗo	ޞ�HR���n�x�����IsU��sX��F�1�PX����L��+M�K&D7kx��~�e5oH����Ӵ*�祴��u��ځv��lB�1�� n��yݙV&8V4٭]X�L*h��oËz)�[�gH��un�6vC�
�v��������m�4�.���ɵ��3�0�z98��X���vȬ��a�Od�-�PkaCHo3?R������5V�����]3w��3b�)��py@�����a5����r-�������-�v�ۄ+�X!�y�]֞xni����@�j{\��=�A���\����8����p`�Խ�k�Y�.1��'�T"�*�D����F4�z�Ȟnk�R��OAԳ���TՆ�=��ܖ��ۡ�������I��FY\l@�Uth��e�]�r��Q��a�5�ec�U�z�!��G����Τ�Ò�e�[��g�Z�����¹N��D0snrR]�*Pub\l�����He=�:v�.����C4�C@�3��e}����}�'����@*�Y�%�_����Sך���V
Z]�U{�Xnd���av�u���)�7-�w��fO��}4��5k�,����\顁��\�R��"�uZ��˹}!��R������j�5�D7��N�����A��H��H�y�*�]�p��s;��a�_ܬ�����]S���סJ`�A}fkZ�_2�f����T�����\(��C�|L��T{��Ӫ1��bQuqA��;�SQ����w�����h�p� ���1��,slK�Gӈ��Xw�yz��K�	�I�uz2r��hAބo
y����#
��r�Z��W����/���SW� !s�]E�j�M�6ɄSG��[,�Ή]ёNj�P-/^D0Ӳ%�(�w�T�8��1�T��e�2�.�
�2���fK�"�g_�y=�(��'�����~=��P��'�X[_��bO���؆�����b��_�N���3�U�y����ʢw<�����^E\\���f�M㋸�"�[Rc��,{���)�kF�>�V��ﲓ�{�p�!ZS�zͶs�����KZ��'6��n�b��#R������Ǔ�A������|,��=[iֲ�዆6��OF䦭��\Z�]�]���`���e��.��;��䓅��}����=�W�?�y���=���1���gm�ś�3�ͮ``��a-��.��x�3$H=re��>�1*����znpt;�e��	��v�ܸ5�k]�Cf=% Sqs�t��'���{$=�+y(b�D����y���5$l��|����h/~k;�"0S�+�M�b�I�q̺����`�\���O1������C>�S����J�b1�U�<���Ԗi�q�֕k�����k���N�w`Q$�=��Չ6����|;@����zZ�D;	��U��7y�P����f<�{�up�|�G�Ǉ��׬`ei���<�����{��}�Zm^���|�k�
�]Clc�3�t�G��R5�ӈ�,@N���3-���zxh}�������WP_�w��%&o�����k,��|���M{�S��%@���:Z���f��}hY�}�	��G^���UD|�D�.���pą�1��|�~K�=��ařúOD$����'���W����ǳ|�H����8�~/�� ]ó��Yq�YX] .�e`+�|���Π��+�$j�L�m(�������t!*�!.��ɏw5L˦�fQҋ,��c��C�sڒ|4�����W�f���iv�'-�wk��_9F���Y��3�l+;�u&���Y��w����>jnVj�%T�}~���
hh\�}�{�(x�}R������j��3,�+��>IZ�w�ƫgP��?צW��˯�
��7��36Q}�����|�<��{���)�x��3��u�XN�w��Cy�����f��V�"��m7�L����L���k��^-W��=��*�&�6�.9�*��O��.�P�����yl_���j���}ΰ`ȠF��2�t�7nE�����@�q�`[�����8�n�Ӎ���yb׀����,����vv0P����@�'K�*�B� ��͏��>hcO���%��v��v��z6L��؆�UE";;�r��x�dd
��
��w�ߢ�#�ύX���	�.^�2'ڢ;;����>��-���M6ڊnԧ%�'�,��%t�C��W�uh=�k�ѫ{՛v�V���~�=:\P�;#�Zg��=Ŧ瞖`�X��ŏ|r|)���7U��c�v�/s�J��4$x���iO0��%B+��y��h�����ũ9w��+vw.Ӈ��5^���_�
��H�v�T� �A�hw���n�<9�|�{�g�e�������\�͘I��DͻZko��Tkc�㛐Y��eTN�� N�1����R�@�X�Ǆ��'��<� ��N.Yʕ×|�4�ҳT�n��_H�r�'d�����^������p�c�vR�"T�������}'_��
hhD�;��}:B� �b�7�+����QM^4PᏛ(�;����ޠ��Y��JC�Tuζړw4l�g��4�x}��;���ʣ���U�W�w�_Aǵ�y~=;�FUt�p�����͞�;>|%W����-d;;�k��L������w](����SEI&M?e�����Żb=)��_�e��,�8�7�	���E��sNC&��˱D��A�}5w�7Ɏٻ�e��z�d�Hf�x,H�6\W���J�4�+����21YT������W!�o��|��,]�]�������E��=�TЪ;��ػn28�nG��d��GM&
�2u15@���j�O��z=��<zy����KfQf�E�١����{	�u�G�n��G�۶�+$��K-�7#�g�G���Mzys%z̨,Q�s'�,�8v�g��W�����x3��F����OP�c��||��ܷ�~	3�ֵ��m���^��?�"�W}9�w�}0�,4}��|��hك�SK��_w��꿦7���xC�_�VUю��ڰ����ۥ~�g^Y-��&��I�&cĞm�럺�4����Vf�⋬������K�\pn��Fh�KxV��P,��P�)gk���9��Ίg,�Rw������������ 'n�lt��v���w�G����=�Ouн�}V�Z�d�:I�4y7���7�l+ٕ�@�A���ɉ��=Cs�~f��v�gt�k�uϻ�s
�������э$ŝ{����r���8�zl�/��w�M�1���;ǻ�Y��te�+��>���g6K�9Ä8.��cK��O<���1U�%����1����74�Txc�mz�������^��ǩ�~Q����޷(�)oT�$�;�������5N��Cc�_Q�b �w�vs��]i�V$=������!�\�F3}�=y�sSP��]n�]���o1�Suþ�A�e԰�ɩU�>*)�PN�������wf�8E`V��v2G6������-�b��ڭ�#|4§����P�`Q"`�k�b܌ydvTC�X����ad&I/�%��6�~}�BC�t�C��X���6�l�<� ��L�I�Z��+�Sm;h��)v�*ig�«�x}�'�e:��}⽷mkz��>�����k\SGEp�hB�X���m�SX�굴�>���e�x9�x1�Þv	C����lOgZ6�-Z�Ʉ�l����vY�{K;����vҺ��v�G�L���GK�eD#�C97���uw}�*�e��T���v�V�Ɇ�Qޡ8�K�Z�[�5̮r�m�c0}�ޫk��d�!h��<Vk��W�<���+�|���Q=\i���j]�^k<�ܙI����w~L�ò01�"[��|*nH3���xA���Jn�lW�m'�r���5�g����˸k;pa���#þ|;�6�6��7ʂYB�����똇�Qb�4/�_�{>���C\�#��^���޸�{^s�|�����l=����r3|�o_nK��wl�f�]�D���Lh�+����zc^�@�3������̉��Ku�1���6ٯ^���7li��}�W�B$^bSA���LC�3�<05Ӗ��`V��^��*�#���w�ϵb�>��n����KWog�P!�.�q����;V�<��M�x�ư����_{AW`a\�m�kf�"�_�����'iڒ���y��Wq�4Y�*��~<��۞1�)�XӒ�.䊧�W��Y���)�UӬ4rR�� Q^�l[[�w"���χj7�{��(�'^��7=���,z��z�{�U��`O	�YΓ��f��L'ݻ纆�v��`p�5N~�oA��ь��z��VWeqŜY	��7qbt�hVw<��f�Abw4�QKW���<Ik�\�]��"����ałe�-Ř�]|��,:.�vɲe�v�l��u�(���hn������&�I���Ls���Kw��9'F0c�|��_;;!(��l��S���hY���8�;X�9��|,�`����FIہ���Ξ�MY��Y1dĦa�w��v�C�|����M��P�	I����J�mg*)�S�ɳ��˲�� ��Ɋ-_��G��O�@�@\�kLs��wΔ�K���%E�^^w�D����H��?,s�m����+Vw�7��:-��8�>VED��������I+��%Ck�l�kjiBK�8�bk烈���&Wi����_�yդ���U��j�����Y����-�h)/C�Wդ���t1B}����A�tWT�� lD�M�, K�y�Ơ�h�5��q��*��Xgz�C�	�L�#:e@�#�we�~*��L����s������e�Ne�u�s��o[Cp��8�.5��^��S�#|ڃ�FR��թ8��ɽ�y�[�۲G��r�%Y��D��%�L�e�"?�N���3�7�z��S=P+�n�ӏ��V�x�7V\,���Lۘ=�BD�j�7�۔ڲO���DѲ��W^c����;Z�H�c~>�mn8�ӱ�}������~���`����|�E���se�g�������q���
H����`��p���9�y:F 썞�Ls��e�7y;��$y\J�6��ζ���+���Ul�>��!��/p��'Z�������G��>�/��{4�r�j�աV�s��<+�W)�/��ڮ�4۹>�!��7�yD�2;jYE?{^K�
:����t��l�g%�8��g����r m��۾����%�7i�g0Xuapy��Bx��ֵ�X׻����O@v��(��y.:�]���x]�y��V�9c��vO���F{,�B).��o���u#u�.�bԜ��]9[���uz�]3��ϫ���	i�����b�9/�KM�F�la�ѝ�X��G@�J�f�N�?V&�͜%G�;Yq���H�GAO�Yg
���s�O�:/�����|��g��rm��K�#^�N��KT+�����'z��c���Y�uWy@���1�ϓ����Ƥ���\cdDC��Ru�=[���5机��xޙgt�vǯO�k����	��P s�tR~���5��&�:w"��y���5HR�0�a�`9�j�ݟS��n�q�o���G/�
��{�c
�ݴ*�e�J�*f���y�~��q{�c3a��^�^+���h$@"}򗪎����((�uӗ��kx�z���p_ޢ�W68W�o�I-4\5�}���-$��`�����O���� ��;>�!*�k;WY�]�p�
����?�<��z`��B��6ǖ���i�������Y.ʕ���<��t��T��1d�Y�f���%����Sۃ4L�Y�s[.�7�ji��ޛ����V�ï����5x�Ww��*[ə�]ͩp���(r��\�Tuz���������I��.�Jr��gp�ܞ��A�1*���U8�!wy)N�,����P�IX��E�g��$b��:�X�*`]ʡc�d��9�ؚRa�#n���Y��An^��E!������hE����ӣܴ>���RM�Gv2+]yp1:�ʗO�������:f�[�#��D{���Y�!,�Gz�v��A���>if�۾c�;�/'0aݾ�50{5ɵ�»Υ�A�+���=Ӳj�ξ���WYӦ�xew50g�-q��Tgk�Eō78��r�q��k�"��S�|�"���h5h���_�}>o#�ڜWg�Kل���
hf�*���!κr������3�PG�H��2c��Wg�Å��]փ�����@yv�4���!�W���Z�=�7ۧ�J���Y�J�Q��9:����V�����oNo��ޖ��UP����s~l�Gę������z����" {3G��}�$���rʄ\X������������Dh&�L��3j���M�b]P�D�V�,����"/�uQ1-WHK��k�(�ʰ�N|�K�}�'4kنZ!�8Ab꾒�ϙ�u��O�
���~羟x	#*�����ؗ8��Ѧ�)�I�ͮ�o[;m-��u��M2�s�����ݳ�=�R*+�'��W	z��3����J���']p�4\�J��l��>w!i�B���V��jX���&�V�Aŋms˄�a���Ÿ���̽�n%�#�;��<쬕tVwCw����8ԝ�;r۔��ʽ�̇iC4j���,�W��L��c�ӱ�ei���i�%���믗Lec̕e�m;�Ͱ�є8n>z�Ff�]�VMq3P�p�:Ħ�u�r���3)�[�Wm�S�[V�X�9���7y�X��n���{CI��fs�7TÏh����Z�b��H,�)#1�aO�q1z�w��q����Ȗ�m�7�QXH���.��sq�U�U��Z�� �{�gM�٬��Q=`�� �+��Y���A�V�N��I���Cet!r���
��V�)�����<����Em��WO>l�]��V�5[�y�����1s�6���tn��Kr�鲡����׊I`\���x����i>s��5��3�B�شջu��rv�it�n��d;#9�Er{��\��w�R���n�N0�37)I����@��=W��ϜN:����z�W���r��+�nk#�!q��II"�|x��n�<q�8�^�N8��ݻv�@�M���� �lZ*+���nh��5��W��ow��n���:q��}qƟ\v�۷����>+������cx�r�nm�cX�幢�c x����N��q�v�^���O�]�v��Ȭ��j�P�qj HŌW��Z��j��5��u�m����c��k�J�)~Y׽k���o��r���E;���.+����6�����cFh�/;�ccdط�ίsw.�G0��_�̢��W,b��W*��5�6�^+��ΣlS�ֹn��\��\�<��N�\�v��{�[�rg;�F�N���y#=�k���{��� �}���]��X�.��7��u&�Yjp!�UԞ��/�f���6^D��5��xxW��{�;�-��v�-%X�~�~"o�&���V���-����-�>�O�5��7���MawŶ��
�o&A�5���v��q%�߽�Pj��w�U;���c:�ܸ9�g�F^�~�"�D�3TݰL�׸���k���gl��y�dN}����-�&͎�_7�ԅs�evW�6n��w�U��~N[�׭E'��ޡlo˶�n3�ѓ疛������Ѳ{k<�j�x�o�RH/c�h���{\T(���Ǭvж�ׯ���C}��VR������c���<|���n��v�O���и,�fC?� �]Z�1!=s�.�Z�T������CUY�|��}��l�5��r ��xW�][�74���k��4�T�~���?��o\k��j���{OŐ[�سn�;'f������X�c ;��UR�����z�4_K��'y�AY�9Q��91���ɻ��n�����M�����^#?=�N�
^�w�{�-��tTSW&����_QvgὝ%�P9:��K6}t���C��F�n,\`k>_Ɏ��Ӝ��#�q{�Ѱ����hjn���\��y;�;{���.oo��>U�V��c�Lk�ʵƲ�f��� ��-TB�,�dװ�cp�;{d7�h�L-=Y�2�1�%�k@�&E�'��p�)ܗY�N�Z�o�-y����x��7:��^��~2.U(�(&�ӮqzQ��Aa��K��g���r�_{F���Y��\/�;�˘�O��С�?�,��VP���y(,2��)���0^�.�l[|��z��_7��f ��% ��|�<GB�W��/g˾���79���r��c��OI@�Ƶ�ح{1a��A5W�}��)��gJl.z��?�ߪp�+�_U$h桽���-�M��Y�3_O3<�'lxn-�J��x*j��I��~t���`���T"�B�]���i�f�/'b�9K?3u9gh�f竃,��#��;��L}s����KwH����T��_��:5�����H��=��]�.{xO� �kn��l�S=%��o�p�!�SmdH�~%Y��]���e�ʞ�5%�$t[��y򚧗��u��)�����=��9���a=7�/���0�Wz�'r�ۛ�q�;&��g��}�y��O�!�q�\����dհfC7�#��+��q^ޱeѮ�+޼K��7rd���u�q.4�<�Q��lh/��	��qpd{劂�9K�o�<�[�0�M� �%<��pǭj�2�wEF�'���=��u�
���J�]_�԰�����8w/w���d�:]�A��gt�-�ZÑu[��x1�p�X��ưojBZ��z�ib\�4�`X���
�Va�;Q[5��� k�7�y���:��Pi�$��v�����ۼ�gl� �<����s��K9%���_�C����L�uO�w��j��cn;����$ḼpƸqP��JC��Fg���y�e��R�P�0�5%�|~�];ޒǺ:�)�M^�^�w
=/�S������������`j.�>�LZN)���ߊ���2�%}E���2=�B��{�4>�M�k���va�����0GpK%�_L�ַ��AM8�DEs�,��B�^���cy��\d���GkT�P.�z+9�����:;��
�	aS��	}޸Y�N���w�9~H�c���y �����6;Qk�l����;��'�w�v?Toj�.�:1��8��us>�q�dK�Ն9Qt�:�u�ϵo�8���<|��G˄O�$��
{��Ķ��y~}��j-����̕P��b���;>:��@��7�@W�-Q�qwȎ�]�p�ؤXKhq���c�_��@� #ݖA�����cX�G�m��v�:0�lT�v����~�ѐ:n32,e@髑M,YD��p?@7����;���!�ʇ�Ѕ���Ѫ5�jI����n�F�ȃ�Y�Kr�t��r�'5����c���8m�t�{��ԔAw���&�O�m�!ۓ�ֻ�/��5��ᦚ��뙌Ld78L7IԂ'|�QQ�%�;��LW2�lu~��<+���{���L��-l�Ǧ���z\���O�������{����dnYr&�qןX���R��X>�[^T�lٵ��І���﫞��_/9r����z��p�����LK�v�:��hI������e�Ůz�$o�jP
�f��s��1�X��^!��_&/e+i|��N�Iaɷ8q�c�`g)�7�������y���7����r�8e���<nWv��;��0]�����P��%q�c}��p�>>�Vݖ=��$^�q
�z������=�4ZRTqq�AN��[W_3��z;2���n���8��ѮUڻ��nFF5i�U�率|@t���'�xc5|z��~Ybo� �K����(���E�b�ob%_'�my6}�./XF�|E��sO�Q�K�ױ��rGEwAc�&�(��|���$��$������� y�[�@^�TJk��x�� �5�痍�%��w���&E�����َM+��3L.�d[�LX� ��lp�ﷴw�ˀ!��X���{�[T��������N�>WBW�مY�U��38o%� ģ�\��n��O~X+m�����`�Gj
�����=٪bt,��s���x��49$#{w�[F�w(���1,���i��^�����䷝��M��v$�6{���<�`�y����p�a��������0�����pu ����:`휠Eaݕ�8�X,��#�a]�y?7ӟHѮ-����^H�ʅ)����sĿ��X�'�;��P�/���U<R:��/��>y��+�9ۃ�P��$@��(��0�n2�ֶ_DK4�.�q�HQΗ���*�zc����'�_�m�=iH��3�?B�aM��IޙuӔ�Qp�gF�v�_?�z�/��R⮢sbbb�[g���8��)�g=�"Q=ߜ��j��0}�x�u�$��Y��<[�Y(����nj�����W�}B�"�ߏ�8����Z1��_v�X�h3��u7����3���� �>�����N4͊@�\J��ۂ���1^,Q�O{N�J�n�%���RM�ہ�%�m�2׫��~ΑM��s�FC����@�ĚǙ�z&s�����]>+9�T����ߟ�	k��:�D�^�6zz�4=�=Ζ�B��}V�Z�d亅�Ӛ��⃳K��;��Y�P��>�y�����^�K;�[XP|���ׯ��[0��f^��ܴ��O�?�9�J�v���]�U��w�uu[�3���kR`�wJ)qs�\�[݅���1P�@G�w�ALMޱ��`^�fd{@.�5*Qs��R\��eh|k�%�/oH3t.�F�jU�&\X�v�K���>#�½} q	c}�S��X����+?^��r�=�[�h�v�r�sf8�^$�mۚ-�g�}��v�{���qϑ �x�}�g��hjH�4�����k��oX�MR��-�3�a[.:}�z�p�����_�\�&��q
��]O����+cx^|" ��S�:��Uzz���)�_v=�l�gTD�	��X`1���^�fD��RZVLe�=`;k��Af�5�aم�5��k�����ZQQ�Ǯ{���6��t��e�B���"6�V����ύ�k@�����6��]�q��N�������1�|Z�U���}��1�H���E[�䧻+H�s����e~Y����vf ڍ��O�V�p�{����-�ު�������ۿO�+<·��XF{�d3�5э	�0�,˧�A��P����t����u>��A�D�@���|��N�f�f�5�Ӿ�4�����3�Y��\"٧��4�����y���|�ϘX���Դ,�|sx/��Z������;��D^�(���y�t���v�Ο�'sm�˹���U�7�m��^��	�3��tS�WU�e�[{Ӵ��E�7ܦ��1�*`�D�����is��(��t�qK���x)��0�Ǔ�$�Orڮ�|��R��e�}�79{�+�92c��ښ��g�o�`�K ���`�l��
��Аb��֊G�2���yny`n�����C6�6;I����5�5"�/��E����2���e�5�)�:�kbX���N��1߽�܏�o�����Դ�/��c�׎jj��2ׯY���ۑ����<Ӳ��]rs^E���f�v�٣�Y�]��ˤ�\��>��w>\K)ҳ&����g�i����k��̡G�c+�ކ��%��p,aS���i��3�P�gh��c1F��֍�#a�����1�8t����m�S���].�@�$gد~Zmx������w9�Wl��v��4oG0��o��>�.���n{ӧ|������eqMV��sod���6NU�cɣ��_�<�ϯ�D�AN���z��йఎȦ��.��d�r�_M���/s�^��4�|<:XL�~���x�Q��R�Zٞy�\e�Ҙv�Ƴ\��v�0��k�N�^�)��F���c� ���.H�ʄP�ɭ����I��Y�s]�q<�^E��}��xCpY���Sx��Sa�!��� 4�m��Y7>{�'��g)��uKU�U�A@�/�8����y|��t����V��@��~ll����H��Gs�/��o�Ȭ���5ؖL�����S j���������3	צ��]E\�z+w2�,��3xe�W*�z��Q�r�����;\^�<|������������,~;)�^�*�T)�����#�"qy���TGˇ�P��e�x`$���u����r�՚��'�����[���������7��`oϝAuޏe'�I���^��Su�+������{�����i�P�]�#���[Mb�$����
��aۆ��Ǘ�x� �f1S�\����.�E�~gl�!�"F#�*�[�	�7J����4�u��l����UM��oMK�Xb��Û�,�X�[D��`���\Z3ݹ_H��[VI�f��Y��h�X��>�ǟ��z�l�����<+m�FPM����v����_,_=q�D�yhj�F}j�]��.||���oS�;��=M[Wcz�J��d=�g����tSm�>p'�k�j`f%̸�Agj�Ǐ6o}$�J}�ʏ�����o��^y��.�'��]V�Z�m����Ơ�[L��Z�h�V�T��J';��s��VH�GTizϦo�����L�OHZ���͒[��m���`?d��8�=�Hq��,^�ӽI��K������N�wե٤��̂�oZ�j�X�k��E�s�n��}�`�&���/���rRq�"��㳩�e�)kld:sYǺذ�.=�z�Vk�����<��&{o�(<'?��d��t�����z}S�o��<�D�Wռ�c%�mD��4n��FTR�$K֖�ݭ-��.���
��OH��x�����%��'.�*#n����Ey߭��y�����9^@NA���ʺ���OY-�~��ly~��k_���e�u�1��\��m)֟� ���qm��|hE2���.[��z�X؞��ō\�3��w�05�>��g���kƆT)�셮��
)p���Oí��j*��ԮUk�N�o`t���CN)5Ŷ6�)�0/aJiQND;X%A�4����8�t��x�,�d�d{�x8��w��S��iO�E��u��fu3�1q���Vg�����KLn �z��] Do�q�fǧɮ��w�dH�7DS�
���ݭ�=ҊH2(�_��Sv�j�N��Pz�
�B��'���W��!��}E�XR�
&���;�΢dq�f��8yY�w�dw��|꤯ʀ~����*Ж��u1�����P�j����f�Chk���������s+s*��kx����vֳF�9�n�Z挢�=�dv7{"���P{�8z�y;1���|�V�3bQ�a�\��T �]35����y���Q9χm�/���u̭ku�p�L�G��SC4yߟ	k��5/E0�C&�+�nn��n����Κgq>|<�֫���[�4���S��c��ˋ.w�6��Ĳr��gO���v�ر��5��j�m��vl)��=[�:mn*�.��ݹ]!�G�	6l�K�^xgw%~ɸ�]��}�."&�2'����9ީ�v�Hh���3d=�ݒ1T��׆Ȼ��Zr^!�#��swF03>��:��t�deX�7���x����"���|Hd>0$��]֣v{���l`}�O�h`ۻ��Dv������ibN�
dlƥ9����v����<�4�jqr�Gv�V�so��v���d<������/:l��*�b��e��
�n�U❧7׺kCG?;54˷oV�1a��V� ��d�y��Vy�Ֆ���-�-�ZY�e�
�P����Ÿj-����Y�(\�9�\=)�3$�^�z�n:*:r:TMf�C��D�v�Z�)�����KTEU��	��)�x��j�lؔQx�/U�b�4���5YY��t���s�aQ�:�[Ъ���wwWec�Md±�Y6�'v]4�����k��� ��l�ȱ_3��[ �^}����˾�Vp��֠��,�˫9�Ȣ�"���pʙ,ǀ��u3�j�t�٨=Q�Lm�
��'���^��/�v!+P�uvWS� 4��\\���f��S�i���9���j���+P̭ctf˩*�6�s�J����J�pʽ
�2�n�;�v�dǯQ ݈�7N���\Z�Q�y�B�l2-X4VB�|/%���7��[�-���x����D�+1qSɦ��̼�MK�}�8(z�C7in�*a��d���{z�i�[Qn�x�Cz�muk��"ڝ5)�<�b��v�b�
�c�I�� �9�U&�ggp��<өm3��T�q�����zj�3t^����]s�"������U��"
��[�7[���塬45��f��H�&3@+�>��gX�i1���)��ķ$Sn�Y�v{� m	h�����\ƺ=t���7�n	�Vu��S
�:�K�t�ii�hK[4{F漪��a-�@�]�jn��b���8�
�Ol�5c��y
Q��gg��j)@9�Ȣ��v�-4���`�{������t�p�6V��^�Y+���!m*�~�Ѐ���=����Yeu����Y_^?�Y�[�A��9w�9��[C|:g��bט9"d<�	ٴ:�۬+�������^�"����(PH�.դ��	\H�A�sh�b�t��57�\ba�O�6�t�]�w'��	4��q�Μ+e)��4T�i�����.�l���Ԝ�S1��R� zV���ة���_
���CPdڇ�c&ˤ��JNrt���/g>yEC۳o���G�H����g?���A7N=�J7�w�N�vݾ|]YWZ�� ��n������1�zԧ�/&�zH=��*�R�J%w[1��M[��F#�����F�p�1�(�����N��"���y��P�;{��M�E_U��t��:�1l��tu�Z�xy�(E{��"�����(�g+�wW*�+�}�2+�����4A�xF�)�oe�/�7lq
�x�:Z���X�k/8RZs�p�WkL2W%X�^n�'l�t�l��p�S��0;��]Y�4��w�Op���\eӥ��E`�c��u���Z�V!��1��Mҳ���kSa�w9,WV�u9M�QI}�+�z�mc�T�/�%oR��S�+���^e��N� �:���IJ�koeך�|ٚ�����"��wD�T	$�I#���Zt����;qǯ^���:t��q�HI*���D��-s�W+�s��/�����N�8�;qǯ^���:t�ߵ/�~W�}79ȫ�����_�
"��>�ӷ�\q�8�����ۧN�[� �� ��"��J#��ۻ��6��Q�~5�<n�K���z�6)*M��[v��|��Ȩ��:��������o�r��P�����ʍjx�;m^u����Ѹc}[��J�5�E��y�W7�S��^7M�EG���}�$^�����:[�ͷ�EF�t�.m^7-�ۏ��{|��:�IDcm�
I�Lr��0�EU8IjC (�i�
0TB$�$�=E�j�����5����5-ܰNYU� �^���&^v�1}W�-=�E���|��~��pF(����cH�	,p�\a��EH��hZ�RB>:$���.4�?D� ��&?�ND#~%��a��F.$LE(�N@�e�ТS�1�@�p9E(XK��rE��.�]x�uR�Ο�E44SCC^��s/S�X��
[6��,^樘��_R�y	��)��4�s(������ĸ�x��>�ݾ�c����7Z�O�����u3F�X@�%�c��z|��j!�u��zha�6{��X![��w2Qt�S���(H�>5K��9�x1�ˇ��:�dQO���Y�e�	��==�^X-x���@樼G���Y��!�����Õt����&v"�f���Nb��E{���a	��W=��� �S����t;k�XF���^i��-B���s5)uY�\�^߫��ۚ�G�pKq�x�y��n���>k��lz��5�\��.۬}&��	�ѵS�Z����;@��we�ԵS�����!�`Q:YՍ��M+n���O;T��&�hC)�dow��.ZEr��Wq>51���Ec�y�ܧ���90y�Z�D�ҙOb������س�;�ͧ�9#���e��G�]]��'��*��d�J\µ߰���g9���EY�k`^����,�5�e�n��^�O&�{�,���l7�7��֋j>�B�>�WM��})��C���5h��k׸S:����2��;4v)*/��A�o17=�W��{��<�þ����\k�q����R�L�o?r]�*I�������0�m5wm=yH�81�-Ϝ�w~���٪d�3�x�^Kc���=�����<=�< �TWL�{t�ȪIR������������3��:舨z&FB`�/�[��5P���͏�y�]�UeǷs�|�Q~���q�v�C���SFa�F`5�gT�� �N�<�-X!>��/Sj�f.p�9a��3�ղ%dY-��d�ʓ��v<�V3I9@�I�<k��q���L�$cf71��p)b��zqEa���{K���"=ƓH�)��6��jK7����_-�,���/^x�w�غ|#t�M��3~l�<{7�5�olr��%�;��dѿu�o��k O��3Oi=��9����K��C��,�Y�_��}�/��=����`���1\��*��z��Қ��]K�����:�7iP���
G"���d���V�f�Kj}+
�n�Avq:��ɴî����ְU&�����8�Ϭ��������s��%�u��"cPjb�CqoT�+sv֩�1�U9^<�߃�C���w�9�^�Jq�Z6Oѳ씧�˳nư�=���憪��~�W=��m��S;�܋���
ӧj5�J��H�꾜���P\��x���3��(��%麛o3$�W�҅�N���?����������o��={�ڱ�3O��\B�:'N�G�<���u�j�}^8�
5Onߗ=�e�߆n�WI,�j��	���x��V)�׏ٶO��B\P��&������b�E�Ej]r�3���&}.��tWo�n�4Ʀz~~�6�eZ�&I��rPs4�?u�?��s�7��cJ��/��`�Ξ�<4A�k�n[�;������R�Ԅ��Y5�,9�m9�]�~��=ٻ��l��ٝ��X�N@{�1��!�Ti�.A��-��2����,����gMQ����r{�e��@Xf��7c��Wm�ɖ�Z�=%����'C]U�C>cZ�?���1ҹ�#����l�k0���ǻ����ׇ�{Y�u�	C��K&��R�T����*��TuWǩ�۷]�������ߒtZ�A_@����!�wi��䃨M�	�����*{�?b�o�9����75���r�5����lU�nU�;R	���^����נ᫞O/e�;�G���@x��ו�j��/��ƮC��<Y���H:�c���o���3�}�O����o�ޏ4�@��9/���]�\J��z_&�<n&���Qx���:ۀ��� �}�*@��|�]Va��"t�{��M���B mF)�������L���y��B��K��8�k��ŊZ��2_)��k��|�Et��ipg�[F�f�j������a�Ǘ�ӣ������3����=gw�Ɏ�v?wK�05�� @"c.K2åڻ��fCػ�ɭڏ}}�8O-wgm�j�����j�,ѽ�i���b����7�>��8Ӎ��a��%�^�8g�}�Q�o��c�j��A�[;�l������k�u�ݪC �{���3�T�u��e���������!P��G0�b�A��t㷝�{m�z��(m0<����ω���~%i8y�1hW�*�|�PGem�����W��Ǧ��E3Уxfu�Mi��qF�5i���JR�$F{���<|}��c�a%��b�_-��k�gd�@�H�U9��Yt]c���M�n\�k��l߆_L�# �wWq%�7��4`�m׼Z���������r���db��5�B�۠����'�����ث�l��w��^�@L͙�".z<�����dz�؅� P[ս��B��ʵ/k���[��&&JK����aUp񗝯��i���ǽ�OOB�	0��̃���/g���1P�H��>9u6����C*���Ѝ6���G� 뭃W��Q�b����9{�ʕ d[ͫ���K�����Wb��
P��q�@��zg�z|�I,�o�|���O{o������z�Do��@U_uo�b�s��9Av*^�a�t,����c��Y;�{��h�N/�~����ǭ�&:�cO���U+8����"D��p�A�r[9���U\��� _�}K�׬�wbl�j�[q�3Y'�oGA.p�ㆩ��7}.J�Y���7�B��T��@Iy}��ٕvy���iOؽ�>��^�J�r7��l�F�ŷ��jI_�&]���)B������%����zW��Rq
SFZ3z�e8�����=}�E[>"���\��ؾ�xp�~رwW����oʁuf:wA���z���~&��-��;�l�^�2�Z��^6Ԁ��Wd�YG������ͷ��������ec����z~���e�@��\��lOfD��0���A�^�s�1�`�<�(y{ޚ�L.�y�
�&�AGf����%}����ka�n��Wڡ�b���D\�N�⺽��]�V��o���9ܯ�����3������s��w$���sT^��肪���y}�-�톋r�������F9��L�N7z�4F�DoLw���Hˬ���9v�PCf�.u3]��4/%>��{Ob�W�rX���e�+�=a��)l�]<�w%�<Ğ�pL:��O��!�F��.4w6ڽʜt��Un��vl>!�����w�*��a�I���!���]�~�_!�d�8~4q�5Va����qĜˣ���)j���m�,	E��Yv�^��ʺ�jP�L�7���"W��kkupr3�d:�|G+���zk����9\
[��N���L�l���$�i�gP�?E�������TRL����_mB.��w\;�`��]����Dq�_5���&!�P3h-�ll��Ր ��LM��,�SV����E5��vo�5j�g�2�7���c����7ic	~mtB�+�wP��4Y��h�	lx�)��P/ƻ��v�W��j�|���A���=�H���'����*
��s�9�wf��F#Q�+���\���w��芓�6�vם�v�IՎ�yB����U�N�����Һ�-*�^]�������A���y�P+�f�RC��#}��I�n��TQ�&�f��7HӚ,� ����&s���7���-4{�x�ƨ�[{�j} �g`\Lx�oVl���6�|�cd�	���;��Wɶo�/f�]:�ӖyW��\y¼�Y$lK��ܙ�9lh���S?���e�>��GA�1�+�ӿr�;t��r����z�dV�Pk�8hK��E/��'g«��[U[U,���ϟ��w&�ʄ�&���U� a�� +?��%^}ֆi�^n*]�hǬ��^����9R�H\9�NJW�z���{u9`�LVK�
����w0j�y��o7����I3 ]�|���]��:�"����۵��}�)�m��c.�ˆ�jv�ڷ��k����4�-��ױ�9 6���oLb�5�V�V����3fXљ��d�u�s(佹�d9�}�zZ�5\�Y�1�0�ך���d��>�����6���6��C��E��������ٴ�d���ިm�q�����1iu`^ֻ����f��\:�?�Φh���"���n�����S�s�獆�x�Q�xzţ����ٙ�t`�m����ͥmh�A�r�����/��
�Pw�H��;v��N�=R-�q!=�ä%�M�9�қ�*@�bǧ����R�o��;p�ޜ�]�LHjCI������-�23�����%�eqb�6�bhm�����1�͍uV��t��k�x�]�y���=����
�$(mĳ,���T���[�0VGʞ ��]�D���9\��Q���Բ�۴����Xͧ,s3M1��	²|yP�6�t�e����v�a�s:���������dC���v�� �Xq�&�7g�����ap�P�3\3���y��o0���؅)�,����m��ֹ��P��.��^�3�Қ+��{�؆1b�Ou�w��0f�f��˛���nqҝ�^陘�GN���;��ޘ~�=�HF�]d]n6�������t'�K+�K��<�fZ�u�B��[���wcΈv�Sӕ��T�f�F��#����s�8㭈�����y���3�����0���j��7��7g˕�u�؟>Ϗ�����߲�u��[7��']o0P���
z�uSR���w���v4e�{�(�zx��L<�c�;����p��"#{�S�t�?oa���.�Pՙ�0�o5�K��c ��޹@=������")��GS���'l30YkI�~�׏)5�˶{<Q�u�9Y8���ݴ�l��q{�k�v�U�lZ	�U�LM����_\7����Two��<VǚԸ�}�^���"�\��^<�S�F޹ݔvu��c8�y]O��{�8��:�TS��-]{�l����8zj��^վk��}�5^�_d��@���21�0�����0_%)�� &.[;�����+��'b�/*�Х�়��\���\眬J�2�E��Y���O_^�t�7y8�c�_���Wk���j�k�c��L�U�j
J���R��o6�0��W=�͖_����vm�ɀ&�����k�Ώ ��bÎ�K�M�,��z��ow���0z�5�s�6��Dm{��^��h�L��r������S���C�lOi�wF[�����s5<����<�y��xn�r�e�Ym��wP�h�ʺ�����˚ZU�������p\J�O0B=}(b�[3.E��-��||ϗt/7�vl��2z�*�H���/ثV3Vs� �F�SF�h�!ÿ���<��U��Yt�r5ʷ}
�����֬�\>?n�5uf�C���uʟG�c�F�F�AGf�n�䯫���E(�3�O.�4:�Ro��t�F2�O(�Z��*�U�J�PN���XQV_6B�gu~ݝ0�l;��Կ�ϯ��>ڕ����뷼W�/�H[�������!��4]���@���_O���/n�5ǜw���aiH.��,`ٗ��J������4���FV�S�o����!{�>��|7T�ʂ�$�$�%�LK�0�8v���X4��VD�
�3���d��<U�Wr;Z��6�J��z��r����s+�J(����U��[�7�z��W%��1R��E�Le9���je���V��Uͼ�g�;��g@#n!��2���(t�A���k{��-ѩ�L�����p#��e�-���p;=R�&�9:�d.��H63k6�X��l�hZ�;8�Vem��6N5���_@�҃E��P�j�Q���Z��t0νOJn��=�����gӼ[(�bޑ��_P]��SS�8l�ފ�#�z��xU��"�U�,4�y�c����kc��g��hVU���[�P��4��Vr��,77�Wl����8o�h�3�he�b�"{mD.�Bx��,��h"���p1K.��[h*���iupVJ$����f�B�E�^%z�;Gum:��{ ��4���ܽ{l�μ�щDG*���TE��#Q}�t(4��AG"���2�Εy&*]:��7�m��ʲ���%�R�C���=h��2��9�Wb��캼�;�Jϲ9�j���
`���j�έ�4�d\"�M�s'Un�F�f��>1^U5�Q)^�J5\��g<�y�5�,�xю��b>I�@!����u].5,�m�+�=�2�۷xVӀ �t��Y8c�Au���݉��wݹv����Y�%��RM��^y���i	,i�Z],W��lr�\�����H�������N��}2V?h�̝�w_\g��S����7��*�n븖�(��-�",^��5w+�^e2�Nj:	�����q5�N��b�K�w�ޝg���;nn�:��/���Lغ&ԫyL|�Up�x#�U�xDz)ڄP\̈́�,�;����t�1ǎ���Pۮ��{�Wgd1).��S�eYx)əضWf�[I��;�{��'Z�E}�"�0�՜�o�S�S�7eCo�e�o���t�A�s��;L<[�V�8�¦��*�\N��1)DT��g7��sQ�{1d��=�٢=Z񱭝=WW�Q5E��H�/7uj���<���t6��n�ȸ�X��蛹��B
��hZ���a�=��=o4����� ݳSbڛ}$�P" ���9�S���x��^�7���|�tcZ�㸜#�K*-����-�aV"�.�f��붯7mfc�㙔YRm<���\�&����]b�*��+��
os��;���S��2�:�z]����,.&���hR�e�݉[jo����,�@�v̘����f�sq@Q���w,=��"��1*×�wD;�9��5~5�����W-�sX�B�P$	�@�q㏎1ӷ�8�<q�ׯ���ӧO��FD�(*U�[ss{9o;�v�ѵ�PI
�D�=}v��;q�qǎ=z��}v�ӧ���J��*��ү���%�ܵ�5˜߻�|�X�ێ8�<q�ׯ��N�>�j?;�	F��6��Y-�����;��v߾vKθ�wU�s�q9�_��F�7���4b�(�ؤ��w{�Rl���^5�mӛr�~����wmҘ2F���^q�یdӗD^v�+ţr����t����c���%IN�E�0�bd�ْĒr�]ݙI���殇�Q�������%\������y�;��RM!���$�%rc�\WdH<�4�������y{�2sǻI��%*��&���0̀h������ݩ�y߱�&�J���}�M�=��Y{:��j��܃m04�H�֫��@|�G�&���ӛвs;&��2�T,�6�T1MHz>�8z����ĈO����6��q�x`����60�	�=����b����i�	��ǥH�i4x=v�+��h���C�f�I�8[l��r�|�+��W&��{�@s�=�H�4��#��&᪲l�O^hr�c�Q9A������t-y@�g��x�q:3<�����*� ��U*z��m�H�lL}~eP�L%R)G�Wј6�Q}��0�(w>�C5q�닞6�=g���9�ߣV����)^32G_]��s�6�d2�IM��� }��0{֟��ū�2������U�7X�7�[�,̺�k:����O��c��l�Һ�\rz䣳&��y��02�q�o6�i��1A�u�ݏF�.��� ������1qzH��=m���{����U���C��A;*�VW{��r�+8[ ����;4��-�OT%����3;/�1�S�}Ь�������y�]��7�����qe<o;vm�Od{�\��Ǹ�W���z��ۨ��'n�L����d&u�������#�}[�d�mwL1����n���[�m[�nc5[{}{�/W��i��v�R���A�n����*IO����v#����r�㓩�N�S~ݵֳY��Y�Ϧb;L>��7�ө�0Nr���R��9���c��
�^ �}�ӛ�H���y�=��捜�ɓ�V�J�[Ô���Oz��>�5��V����|�=%�
j�H٬�8O3�&�����p��C�r�Vg�&;�m;u�z�>�Xf�S臓�2*��7Ž`w�S�4���>>�)d�b���9A���5V*��$��ȘM�=�vXf/�;Y��5�����˰b�wj�ރ3��F�CքC)��]J�����ذ<dy����TI��P�%=���\G�������ð�D�	���omu���ri}���fW�O�������U�6����e"���v�k���U�-.�%�]��U�<|9w�`uu�����eao�at���ٽ��lam@v�<�P��&Sx;�d�W�H���x�����v����*X9�}�;�_x��В[�D!P��hD��I�C1M��r� �f�w�}y�:�������T�{�3��_�VFx�nu�;��PX��z8l��}�u�p�J.Fu�I�w^�Kϵ^{*���n��.i>(��`�S�B3�jp�O�M!��T�NP��4�;�ތ�ЦN����ؗ�]�y��}J��_�]c�2=t>罕ǽ���l��v|�f��c/�T�4�xVYhl����:�C�Y�3����T���:b#3�6l�oh]pU��jZ��C�ȱF|ê3k����4�w�&X�ҷ��ȫ�꽋\�ޞ5�f�ɣ��vHr0xڮeS�妪��4r!����Q1�+M�=Ǭݕ��6�l�.靵�f�G�.��/J�iC��5jkf�EoL����rt��Ԭ�v���w�x�G�ݝ|um|'��b�"#�P���da���럊|C�vo��s����Sn� v��Wj����B�C���8M���%J��tO|��s�kHMk;�7��s�2������ۙ���`	�
��k�uè�ub�m��yJ1�f�]��c�K��m9.r��}��Mu��W����y��8� ���w�a�;�nH���򬞇���tN�5w�$�zj�z��W����K۲�g0�����a�d�s���1�x�A���j�;���ΰ�]���I�s�l!�0ry����8*���q�79�Nx�F�������'d��	�H/�_k9�}Q�P�[%z�b��z&��W�!��@	\��>� ���	;�~����nwXȞ���=6s4҈�T�Z�=���W�ѻ�^����;�r�8��w�ň�̅UfM�u{���S�D�3�D�\��H=8�&�Րx�ݖ|�ե ����V�X��ڷ��[�I�Uv�Q|~�����`���ҧy�-����y���]7`��Z���UϹ�ɨ8�v���m�m����٨�se�^Y���g��}@��?z���7,b<����
�ȼ<u�4E��^=���e_�}���"�EX�F����Y�`��=|Q���v���)�����ي8kH7�����"�����4:|.�>�����r�S��'6���{M4
,�S����g#|�Z�nJ�q�o7��z�����2���q��z�z��ٳ�R1ۅv��W���s�Qm|���P������tVv)B�	=$�0�I4���{s����̹js�hk�b�[oS73^s6ʹ�g9q~K�ϗz��+�{�%���dpܪ���y&��6&vR�R�͞�����w]����zNǯ���N"�>N:�Q��@/�ڰ0h�Z��Ne��v���||ih�m\C��FL�������"u��	˝�����典�hBN�$iV���0�
a���<�&bչy��ޗ�6d��1r��*��#��([̗/���s���=�gZ-���@���]�-@�ʼe��|���}�ƚx���KĴ���|(w�TA$�6�_��ț�;��;U��|]��춵�'��C	�����2��+=�3�x��s��8�V+��]"&�и�P�Z��	ٴ�gY.���+3Q�j�'l���TL��D �+�ꓻq�;��̋���'>k���]���16��"P��9uPn�h��Պ'�P�_JA��䯹?>bt��E]W���N���aJ�e�+!��*d�t�H��W����:�8�u�(���.4�_�e�3�3E�r��P�Ko��-�0�vA�����^��UB�8���*s�_�,��F�&�Nt��DUBɌ�0��`so�"%�p�ss����Qܕ�ovePηx��T��>K����b��-�4�}�q�^9��Gݕղ;�����ؖ!�S�k�����g��yA����ɽ���φ����l.��u7Rpd�, x��0��7�wb��p���
��^�{�W���J��^`l{|e�c�*'7&ˈ�gc]���5ҙ��ډ~ܡ$D
u��P�g�48��믩;���͠p�1�)7Y��;��$5��]�Tl3?T+������V5��ގ��i�=�^����h��û��t-:��Oy��)$m˼�w�z���u@�߯q=jF-Q��4g�鬤���cdƱgV�PE��2�#��;���\�wzإ,� S��Ɗ˨l���%f�r\�xR� ��(�5�H���X��ٯH8�"g��4�Y���/"�ݴg_d�>k2,���j�ӂ��asDa�|s�;�3D-�5�������Qu��+��>-����c�ٲ�d�0IB�q��� 0e��-̹H׳y�[^�@4ns{'Nԛ��4�͎��R��1tFE̽6�Г4�Լ]��p.}��㳪��w���ٞ�b��l�~�r�%��qf�NL�+��y,�F�&��H����b��2���d���Zf_M&=�
� �����/k/��(���M
�@ĕ�×o6#�/e.:��k�M�3td����d�z4�涷��Y+�]R*�݊/N{�bQy�݇��DI�ŋ��;�e�q^���r���Дw�=kE=@�dܥId�����L�8�z�uسc�\ٳOo:���1�����B~������u�],�׶kx�zYTu��j���"9.�����*۶[�`�*/���Z"��W���D.Hff�.�Js���F���fa^։��ِ�g��#����v�u{�Zl�������q�dئSu�cH��q^�vP���0��ٝ��^#�m��.w��@��1���s��4�����Uu��7|n����]Gl�\s5�b��-ЫD�z��ZU���]��3Bs�.�_,*+w}�F�:�ݴX7y��o7��3�ʴ�݇bY ��L��۸$ŀbu�+C���3ܦ���h�n�4����d�8)v�v��+�O�o}wϺ�$�y�����o��땭��Ws�/L�m.�tɺ%&�4u���}A������/�@��!r�%����Ú�U�޵ee3�uH4�TWjގ�c���>{k�!�)�{k&=��`�d.�=
�,���`�k��w>ϣ��6}��xK��D�mL7��R���,t{/��0��eYeиo �)Jss�������Za���9e{�*��Qƣ]6'F��pmx��k'\��;Z�aV�bm�ϓ��|�6QlW8�3�����4�k=v3w�*R+� �P�lü��Si F�!$�ל ��f��3Ě����Zi�@樽/Q߾��X�ZȧϞ�y��h�#Za�k�=�ʹ�2j��ɝ�ڬ�8��o��R ��"���T��S��3gE��������1�N�3��M�Z6�e������,]Jٛو[yϣ�)*�'3Gd���wnWZݨs�yj��y���������-����-�f<k2��5KکǦv;��N����2ff�_c7�n��Q�eV��sk�U�g�����fṟ9�[�y�*�4�)ٶ����3�]���S~Ym�/���{U���)��K(�3�5{
c�0�6�� ����.�V��]�-�E[ &Z�b;Wgdl�x픬j�sOv��qh>\z�q+y�n��V��P�1*<o-J݆}���;iq�[wx�a6�u��ہs���Ο��H0f���2Ku*��A��`�;�ax����W��b�M{!@��@-[�9�m�Q4�u�|�'+��]=����a=�ל�w�U�;�R��b�m�p11'�3�G�_�TᔓA���t�;�z���Ѷ�<k�!���R"7�����ct퓏d�:��ǯ�R/J���sJ����!2"����53�M6��Q�9��C�fUܪ��n��&���H��cc�s��v���oo���n'�f<��"�bo����������r7���� �y:�U|{��Q耮�{���=�&f⫙��AlWs�#��Υ+o��o7���HY!Ԥ��]��nz����\��۪՞����M�����a߲N��x׮�O�5d�ZV*tس�5�7=MC\�vV<<��Kd��w��A6��n��l���������|�T���j=v�,��W!�b��Na�V��}$1�]_xϳ�l���?�|��������딖�^i�!l�Yr~W`�B��i�4Ǫz��ޗ�k�DI�����z+{j�4n7Ax��u����9�|;��RC��{�z��Ό�]Swb -�`�U�v�߬��.*=jS��36_�n{����U�����
#X���b������"n��á���e$�����BYCR��O�m+=�P�n�/Z�c���[Ect�������ec�-���:뉈nlu��1����H	[܀z�]]Gd��Y-�{�"�\�hU��_d���G%V�����h��.ZX��`��j�ME�:_��1ޏ�C�q���T�zѡ������ܚ=8�8j����Y�r���ʓ*+�Z�Y���o��]�'puK+P�p`�Ǯ̤vą�s�N˚Q�on,�K��yY�;~:ᵽF�SC�:��]���μ��j,
ޖ�WsW���اpm}۩4�(f�҃g;�s����3V��c�N�C�d8h^:����ϝ�^,�BN6-T�-�Bq��igS���g5
�����g�i�����]�W�0f͙��f҆o�=8�������J$�\�zN�-��pu��*��4K3�S{6�R��X�R�H+�<g�T�Vm��^-�3_r���]��CD1�옮�\]��ʃ�x.����{8i�s��&
�k��{lT�.WG�tz@�k�j�Z{�R�ժ�8�Y���΍��������ճ�L�<y���O1�s��ʗ�H�ER�"�ѼJ�S��s!�녥ha<l�s�='�^����.L��3�;�[�,v�|w�;\��h�����L�)G���}��*�|�m�5ƻ0�GۦK��ܛu��9�Z;U����.��疵��p�v�f�U�}�y]a5�s�[x��IN,��S�w(�:L�=W�M�S.@�@�8���5�ث�HP5,i߶��ٳ&��洳bL_MlL��88���w[Z��q�GnW�N�_��RDm�@��۴V��T�>�xgb"�Yũ�IQ��>|���FGM8$
!ꉫ��6��7�b�D'9��z�� 
�<ϭ}CX�������Ȍ�W����eۤG;L2_e�e<����E��,�v̧�oM��tt�(c�KS"� 7%'�:X裗�nҾW������k)Ļ4����
�*Q���%7��=���Z{f���L�|��1����ۋ��n�A*K��eԎ��;r�m-�ױ�}�n>��v�"�35F7|�O�W�6X=�I%���=��l���Z��N�G{N3*�;�V��e$[���[�v:�]ܰ8x��\np&�!�cZA�(��U��ZV��:�d���ȇ
�d����*W�%	�����e�sr��U���C�h����=��l��|�C7-m��c/m�G�&�D�{w��ҝN%ck+�3f�T`j:]w{f;�-%\�gH���qJ{��.V�h[Od����ݭ;8.��[�&�튓l�ܷ��t�/��\x�2W�=C3�ܫ{�kTH[	��GoWH	˶vZU+2�%��y'r����E��q�k�F�	8Oo~YV��N���36�'̜|`��:ࡗ��^�飦ҙX����<�)��Z�#{��ҹ=O�,�ӌ���8�0�vnW��� H<+��s󮾜�z޶��\�r+�BT*IA҉
�UϏǎ�Nߏ_�8���z�]�t���P&�������μ�.m��{�0!�U �I�(��n�;|;q�q��z��}t�ӧ�����I%J���ׅ"s�;�xع	$$=}|}|;q�q��z������o�����E����������r`^�L�ߝ��stE�Wyܞu�<q
�Mr�7uqz�D�.����Ҝ�K�m׎~N�Ԧ�û�,����;����|;t�)�p�Ef�����_;�wu���.��.�1QI�qB�\�up���d1�z�A�y۽]����v�9�S�9RD! ܻ�P�	���
�Hdq�n�nB~���pI_$��FI@[����¢-��3#6����q�06RG�,Oe�lW_Fs�R���ݛ�glYo��7]��}�0��d�^��s�4s/��,�����+:a�M/���cP�Q&L!4"B#�@�Db\�D�2�p&
r7NO�	|KN3@"(mA@ڐ��h$�qA��Be@�22�l8A��J'��fH�
B�����	��i�?"ch& DG,���~������)ҕ�|�.�
�̃7%lW����JB�m'��q��'^2E4���6ߨ�Y�d.�5zF΀ڪ�?�	"�c�����"�8��}�����=A�
���Ҝv+����^	©�V�54��ѫ��j
�Ԝ�q�S���E�����f������qKֵ�T�f¨���|=���l1���l~6�p$�Қ#��N��־g�n�4`�n�̣��NO�W:��w�g{pmM�6,ʏ�Ƕ���!1�ב.�x������Y!�T��G�]z<���#0;��b�����m\rb�q�[-��5��ٟ�bL8��lL3[��uFb�R�
2�w����!�lި4������(p�[>���l6)��@k.�X^��u�������i4�I�w<�.̔yO�r�8�w[�wSq�30eV�2���V�Zӳ��q�z믳�fh�ݮ�C�*|3��s��F��Kö�KÌ�Ƀ���T�Y�Z���ٖ�����ʴ��8�UXF����qت<�x���:�ϳr�ԓ��mԮ�p�$r�N���8�F{h�ځ.�q�+�bΔpܵ-��y��o0J�^𒙽/X��l��T_^A�Q�Hi�{�ʽݓ��<#��ֻ�&l�6�!��z�v[���Z�uS�Up�ךpS�-�,b[f�]Ga�k-�@g%�V��*�;s)�Boi��Q=g0F+a�F��Ζ"7�s4�EedҮ��q^�)���[�]^��:�Cn���d�t�iڗ%�+A�J܏_��ܥ�{v��<k(���4�{XH�-n OvF!�H:�D�~��h�ݞ�~c>]ȿ"�u��^<�Y�Λkz��vp����5���j���xrz^���)\���'_�wf�Ӭv��b3d �5��h����:�>�U���Y@���.���m�g��ߗ����͍fy̶<*T ����T&7�>��2�L<5�q۴`�(.�P�=���֐G�C�6�XKխ���\��4��H��8筵Æ\��wS������s�����4q�EP�6�wM��귢��6G������}`���:���YŎ܂��p^��n�,4r�H']9�MTa�����{͇���&��y��o������y���*��f'��P�����
9z��Վ�gN�Q���:��!�o�j7��&H�!$�X�u
^�=�=�&�P[��E)/�]���Qbj�&�|�!�Yx�ޘ�K7ͳ��g�&�HJdX�x� �ىgq*sf7�����3�����H����ˡo�mL��9��\>h�q�����z�뉃�o�����sY�@����>Wڏc�L���egi�oV[J�>����[}'����l6��X�e��Fw�G;=��MXÎa�(���յf{��=yC��O���KX{Vڬ�qt���ͷ��=�<M��l��c����y���ݞ�����f�;�Rmfv,n"�-�w�Dy)��օ�M1��n�¹^�޺�Q�uV.v���0�H�������&�� �>I��OjZ4��xU���8u#�N�����<�K��D7]\�5n]ǘ�M-���(�W25�{H�;V.ë�a΁c��v��MÚ�z��l�on�]W����O�6tLY� s�>�9-볏8~�|||||6�wN������]i�p�ge���d�7��W�z�G�֧��;X��z��۶ι4a���O_�	���Y���.�̸�Z:r�U��	ǉ�p�9ޟR��x�|�oe��.�%�ߎ����,g}[Ed�.ٽ��x|I���s� +�"��V�r�]���̀.>�㆚�Љ�W�[Y^��k��Y�r[��g�iՔ-q�N5@^�]�u"u����F[�%&��ͼ�0�H��f���1���`r4L=��7K�+�^��,����j�cQ�ݗ�=�>��j�NgW�����]��B�3OV��#�RF��4���H� ֣-ж]�μEz���"&�݌��ˌ���َ5�Z`v��H��v�i�����g�����C��kl��Ϋ-�Kr�^��T�%�^K'+�<�E�d<���)���;:[!����q}盰]lK뒄m�M���^ZuU����3�,���!��9y��̮��Y��El]_G{�5��F!ϱ.Y�����9CQ�q��R�N�a��7E!���Ү�RQ�Ν۽X���_�^>>>> 9M�U+�:I��>�oTz;�gQ͝�9��iKi�uц�K=VlӍ��c�N� lw��NgU���H�
Guj[Ǫ����Ѩ�ꍬg�E�ES�W���@�17U�|7#�l��r�e�Һ�'#�ݙ�+nY�02�j��s2$\c�HƎ�p.Wlz�y�yl�扔_{1�Dd]�d�A�ϵ��U�g0wMʌ��v]oE�^p�ok��c��MD� ��+s ׍_�p�Vg/���q2u��M~F���<���*���ǌ��ugz}i'�����@�d�����#�g��j��c*���Po��	�W��D�������7u4V�3��f��ڥ�4��c��b�CX�LT5�]"g@��9�Z�qĦ��YĖ�ͥ�"�v�:�Z��م�g����{�}��:mz�_g�ӷ;.v����{Cc��0�^T_@FC��p½pg��'����v�����~�֧q	X�M(���o/�/{>�˲��ʀ�X�Z*���R��/�{8_vn${"r�����ˍo:.��T�n�&cw��1��mm�G6D��d��8a���ޡ][:V�:�e6cI 2�9���oZ]ܱ����|||@
p�r�f �4�1�/�!�0����>�T#)t���e�Ӳ�yQŃD�l����|H�� $�R6��KCY~uk�afH�=gr�]δE����U��f��c��u�u�G��� ���c�uz_:koA-@Rk��z�}���Y2*��e�	��Ï9��n62��KL;�0r��<�W�6[U͙��U��*_�b�� ܥ�s&Ս�v���ն�rf���'y���D�v
́��&KG@`��賏�eO�Y���k�ive�m��n�e������.E����A�Ī���;5s;{���=��䎕��J�h�d_��n�6���l��:K5,ސ���[恄m,��qJڧ�mv�ƣ�@���5�{�J�Xf�
�V�V�QYf�<]X�Z�Hݮ�
�(���\��b<2`3�ؙiWJ��gN�ݦ��Ļ;l���r���=�[9:�\��mָ��y������_=#�W�2 �|~ #�b�Γ����]�:�U�U<��h�5�l5ݰk#qg�O�Ȝ+�%�c�}��d41�=kEY�LU�Y����y��a��s�Ȫ	�l�1��~.�ES��B�t������(��4��y���S5Ms�mCa}^��;O2`�(_�k6������b�z�T��	��q\�����6s'iZ��n��\V4��w�����p#�m�ș���f�n�l��s���$jF���������}�[�����%c��LtvxZ���;Ž�v��<�t�RN:X�z����f��� %��m:ۅ��"��t)Er���F�R���}G��w��ػ*��Q#Ske ��x��=]^���3Ty虱�B���!����ȅ;b���{�27D���89�/׻ڒ����}��yq0~2s�;ͳ�ގJf�۶%N]�[疅�ް�91^3S��eZT�9�� �s�WY�6�HJ��v�U�g�e�%��11=oh[�E5h�W���M�f�i��7�9�1�:P[�̦�+��%m)6�MJS¬�a.ӢRm�.	�f�ͤP]�"���ZŻW޳}��w��d�'7��4[ckPARw���{�n�����[=�-86ރ/O����y�>J:�m~��2+���wv^Ou]R�n���-v�����3-|���鹹�(���/�;�:�1������[5�r]û7mQ�}E�eͥL�mfgw{~��oÖ*�Eik���ҏz�v�J䷓aװZ�tQm��^*��Uč��wc�#Gl�����t�*ҭ�B˅ة��+)���8�Q��B�m٠���{Mc��v�[�>�3=�����𕼳��� ���Jf��{�����q7wO��9�Ts�4gww�utvg��*���-��\���d��l{< 6�W����!M<De�����)6ܨ�(���ۜ�)#~��4�@z�xy3T��:�PS�I����J�ؿ	�ky���Qay�Y�s�P��wo'��P
ok'[(���>�|C@}As-��Y�9�nO�m�Ř���x�w��s�N-���� �x���a5\�W��b���ξ�߸m]�)S�m��0�ܼ�;he�W�Sx��@�G�� <,Ù��������P�4�t����w7�sf�I�ݢ��)]��<�:h�=���ƯZ����?{�P����⠂f��i��ܼT� �N�;ۙ�ԥ��o2v�{]*2�D�9MQ�]�)�hY�}��'��o&��b��V����'�%�o)G?��ڟY7g���%�Dy��	�K��8��k2��U��A�=.�|P�m�z�)�-l���l��y�3�H1�2��UG�d�����]�V�=��^��\*�zR�~������|��ݘ�ķ��g��x���47T��*���UԖ_�{�+�����3�\�_q���UA�����M���#7Җ���vh���$Vi֙UZ	"3؟*��c�����!��â��G��~ҋ6��C-2�K��[�l��{Q�Q'�N��YF�qT�j����Ϸ���Aj�IR����ۋ0�TA-�ݼ�پ�����	�#Z3�+ ��<&�)��ܩ����\�O��u.Og�G�Ev(�������kS5�5����IQD1���ӭ����8�f���Ȭ�_p�H����w������4 �F1�d3�H�s�_>�۟3O�,ک�����6sG���}������݂wiUܸ�¶�>��=��@�Vt޵�'���* ~������\�zn���	ޛgǽ3�-��_���������]M'cuk���i�ѥ���pk�=���ꙸs��~���E�u]F[d6��E(��"���m{�]�>��t�R*ȯ�X<�^��W$9�fx��:�{������!��`�p0��f3�ʤv���f�oZb��y<�h��M�I�}� ��ǔ���kX�pw�Q��d�6>�����yZK�X����o}W 6j$H�@Q-�l6)xƫ"�:2�#+[�����iB/ ��%�n�����8����u�@S�ɉ�l�n�TE�B��i�<g�C�k�"�v�da	�Ǹt�� ��W8��N� ��mYv�ik7��i�Pw@L�9�J��l�L/\*O�o�2�rt1�o-�t�e!��ͽ =�U^g3>��y�cIS�[ߟl�ܷٓL�e[��d`Wa���k�tc��Q�Bc��wǻ--��r�����M5%���r�ü�8��vrwZ�����0��n�$-�26�oe�1�
�)u�N$�b�;��Y֊�����J���ن�(��5Wm*KG+�����l���)��o�Lm���X����X�I�����eQ�aEx틜�PQճ���p4B�.e��2��r�o,ܝ���T��>
� v�cQwp:-Ú�\��vp4� �)�jY�����a4E�X:kW]��wZT�jeI��J��gGv�7��ʾ�c�{����R��m��q�1�w�%�%fg9������j���d^\'4UVCj�Z�˛��%ݢ/��"�8}���x�d*���n�q��|c����C���S��w�Y��� ���97{8j�mP���b9��L��+�X�f댾����Ԓ*�n����1W����8�J���V��/P�Jz2���M�[蓣 Ֆ̓ӎތ�B�Ft��Z��AS6�37�ʴ�Cmg}��M�HK���&�h��ۻ*yf	|�;uiTwJ(�&�ʠ�iӗ�Z�Y��񐖕��VS�ٖ���0'!}]��[-��kB�
8�mZ��4�gy<z/4t�L�$�TI��H�Q^J��u�8�0�7<śhX�7A]J�׉�9�Ny ��S�%�B�U�ć��)+F�4��C��:AyW�c�qY���C������P̖A��\�.̚;��iҦ1�ʗ��*i��9X�Vv���!��;N�[���������nYtbNª�����K(���K��@:1lwZ��r�ݤ^������{�+R/sM������1�G�\z��Ӎ�,jn�&8�.ʸd��c��x�^9��W`�/k��Tht�҂�6�����e.�k�+���p��;�I�Y�@-ZŬ���w2��Ei涑�,$�R���!���鹿1�,[O��@����1m;��w�������v�J�jmeu��_e��͔�M3��=������9�J��1l����|���9Ut�wr�ð�fv��	"�v�����b֞X6'R�n�o.
��ʷl�,�otf��,��:���Sc�zj�W��Yym>ܝغl�RK�d*��wSS26fgs}v�q@U��ME�k��:�c7�U�]���ZD��ӷ�o5�5\TRi�f)zi�T��eL�/�XX�ꮭY��l	�/�UM�}���r�[�rco,�B���x�gi��w3��4�LYW�c[R�s�ȤEf��Z�h�S�/���Nj�]㌒$;%T�dd���Ӡ�\^w.�*1���N�q����׮8�=z�����N�:}|�e@�#%B�!�]ˋ�<yܹˤ���wq$# 2=�K�G���]����qǯ^�}}c�N�>�/�jU�L����錥��eh�BFB]4z����t��q�z�����:t�����2~�n����D�1E�+�$g��wA!)�q


]�bB��s�%%�\��!,v颛e�s;�!�,cF�×Li#D���u	�t ���d6.\?����K�� I${���,0Y�L�"�M��戓5���(�RQ���1��\����
�wb"9ȁ��)$S3C�]+�-�9���,��d�m���p��[b�G5�ӵ�N�7je��OX�7��S]w��!�l@Iܫ�z��'t$a���}¾��xxx��
m�+�V�(�]���x����_��$.�:�WcE[v�'��uo]�t���aS�0K0(mq��`Z�F{�w-=���U�� �>h���ٞ�9x_g\�;Ԣr;���&��1E����=>-�f���$L>8s����:C�ǋ�r1H���SZnN���L���wa�ۛ�;?o��͝��o�����e�#��*n6+�g�tɺ�dz���ܘT��]J��Q�[Xӛ�a�����Q��ړX����%Z{6ﵓy��ܸ�2������V������';��I�X�b�s��;ُH�:�=�U�;�K���R��PX���-h�z[ʋ��10�Y��
*���ű�}�-*7�n��a��@��֚��kQ����]��X�К��;ׯ0ܦ����ݽ��{Y�g�oX���0��ى�hF2r�a���2����ᗯ�|��:�*�6n%���56��M��U�Gx8��:�'����:h>y[J���/�n�{�!ڣ��N{��<ՎQ<�����)�L{�����FSP�������y� S�l(҃)���>}p֝է�=b����������v���%��
Y�)P��}�7�z|6<֡ϱuz*��͞�9T��A�3d"׺��jB�I>e�gs�������7�[��o�A����������e�6Ow5j�
)Q>��T8���,��4�	�$2�=���R����7f�4Z%Ee�i�g�����=/>�.@���/������E7&u�G���;���d��.+�Hpe���q�9=밾C{1h{�Wy�]T�J-�_mZ�n��|��ף4a魁��X�$}]�Ucbh�l�0�O,pك,Ͼⲏq���-O 9�j���/�t��.����%���4�I�|�LǼ����ˉ�$q9�-�,�}��ܷS�D�
UEm�\�/��O%-��ڟ1.�:��~��!r?��c��V�uV�as􎄵%M�=c�)Sj��7.K�,���<֮�-=���B/1ݪ�-��2�F��W�J&��c�A�#ڑ(@��)��з�_$�2��5j���(�`��p͋G!�݊G%f�yƣ��] �B��&��hE�PB����+��������o:����:��t��R*��bOS��$����0}N��������P8�������fy��e�03Pż�5\�t��Y�Q�R\�
�ؖq���>��� �Z��ȨS<5�0X���zN��6�
�~�|��Iى��Nz3n���WW�b���¸��85K�Sjn��*�u�}�E�{E�P�Ykd��Y�	R����s����7���-��^�jqu�R�g�.,	+���PU#�M�U?H0� 3أ�!s�P��h�eq;����*퐪j�C8�:E�.�M2����wi��!6ξ>�d���+ic���3
�,�a�%�_rO{��x=S���
�S���r��N����.۳/SR��V�����Q�^K;n�x�|��n�7�kd�=�A�T�ç��<�y�u8��rwk�G�UW0m��*���ܜ��tVN�F�rd�����r��֪����u�j=������2r�-ؙJ-��"�DpYc}'b;܄Wy�o@����&%j-wYO��X��u�y6��욲�ع����D��f����<<<<=k�6�d6m��Z��݋����ئ)��_�X���}MD���qAa�.i^�W!u�]Y;�`D�0���G��������!N�\��������|�${N��οw7�*�
KG���H��^/��=�6�p���u;�vSڤ2��a]K�F�+��U|��I2�}�b�,�'7�R��.oӾ��2��ww ��emރ$<�TS>ZI36Js,d�2"tl��6��+��U�Z����+3LM�UDK���
&3Z���>���ܧѼ�}~�g@$�;l�6�W8��9*�:ε`�q�2�l�}��d��[��_\�ut]dueQڔY�^꜋�T$�%e�:��D`%��!�y�l6��ɇ�x�xx]U��!o&5�#��{"�z<�Ე��>F�kY@�ʈJ��Z33�A�wwf*���1�kK:�֓弭�ǈ�ۏ����l��n�+�R�������U����ζ*�D��Z����a�ݎ��ĽФ��B�bs��e�R�0�}����B�gO��/iI/���x�� |@��UQ��05����7'��=�0&��Ni
@��{�vs�#!��Ϊ0A��������9>k�|JDMT����C��R�=Úi������7������Ie�O�[��~�2��H�Q�3^��EMK�����Q�dh��q�+����.)��S,�]�.��&I�W#j�R�μK���s�CKw��:���J;��l��u�m���r|`P�Kp�R�w5ZB����g�/b!_NoF�뤗���*���|s+s��JӶ��ŒVU�i�C�1�Gݵ�zR�ݵ�x�-X�O-4^�V�j�K#��U��{�,�G��jlޱ{�Ƭ1\kp&۴�8��/%�ż�ts�&Ze�3y����y,f��Gi��\ë�,ѿ��}��\##:D�V�=��f���;''�ǟ}b��R� l�>��6�4S~��٤k���e�:�ū�����F�sx^��HD��=z:��h�ܵ,��sD�!�4�i�rھWm��y�N/Y��X��s5R���f蓪��)�����;�.w6/gj�_q7ƣ�c�A�1�w�L�+*@����<���J[��Ŏ��O��>�C��,���0zNv��tƹ�L��eu�ë)d��@+@�T��X�mED��%9��W���Qؖ�xvwY4\
���X9~l=8UI:��r��\�u�t^�2X50�ai��͗�?���02�>�&�&�^%�"�;��a�m�B5O�_�ҡ�K���<GY�2p�`Ǫ���ݹ[O��.V��aKق}B}��2��nu�>�>z�D���m�n�ޣ�t���l��4%��R�����?y�.����,1�z���`j؁�{9i�Rb�l�b���yH��v�H�x	l��������øb���x��1]̢E.T_�ݫ�{���-��5�I
����� �����93O��4���&G�`׍�s�\	����~��\r�S�Dѽ�sj���x�K�h�3yݬ7E�u1��x欧ڀ�W۫���i>�P���,�T�u��s2�"�>�<*[��#�����:�C�KG]�CG�e�)������-��{�������٠@ieu������׽���������.�7���'�.�b�ݗ	��kxЊ�!��M�%���$3rGs^���Ŵ�D�Uz����u�uqZQ���=�ذ��u�f����3��,\i*���A���� ��l�~�Yu�3�9�0�dM�f�i�tE����xn��>o+���H����}� ��f�9�wڲ�����S`7a[�;�|���O�Vψ�� 7a�mfd�E���/6]�H�ll�\��������/@N�{����\y�$V���nٯ*���|d ǣ��hD%"e��=�Gu@G��y�\�b�F�����Q��L�7my{_���>d�Mú`ڸ�zMyH�Pո�f7WYY8���a�
Y�^_Q��V�<vt�󓎵����=1S�s9�enڤv�჻�`�=�������,�x�7o�<#��G.��h�Wb�z�����ƭ�Y8��h�#�)�N��{v�Y����>k0�N�����.�*R����x��/�wd��V�)�y�u�MO뎹\�,D��<�cu",b��v����:��'q����;8�y��c2s��sQAs
�>�e���iջ��%D�ѷ�^`�y���^�B*�|g6���]�ps��P��v��5¡�Vc��qoD�d�N���$GES	'=����.�9E�|M��Ai��ҵ�H�M6�w��a�J}��jj�d��O@� �MA~詋�dfN'R�w��L�]hv���)�=��5T1�m�齡�ҵJo�ˑ��:�Z6�S����*��˫�ޚ�i�ϛ�Bz�ѹ}T�!��w;fu�\'��SZżW�&���9ޠ6$Y`�]b�yx��ؘ�ڶj�u�P��-��7���)��ogk�5~�����թ�&�%�^�䜃]�tf'�����y�ڨ[��#~|����m�i�}�k���� ��g� ����F��ܺ�����"����rQD윖�yk[���G%-gKPɔ�����ܗ:@���Nz�����x�~߳Z��+o��Q��k�f����ٗRe����-
8o���	�I�ή[�#�}���V�N�=5����H�ۙm��_�҈�KM��������ƹ�3�eV|�g8n��J�o�7A�����y�'U+�o1ud����|�$��W�mp�������@�1sGgy�M��e-Z]����:5&�W�f˝��������W3VP7�[��>��7�՝��d;�#L��}���$f2=����+c�WS��L)����l���.$k�ސ�C��������eL�=Sx��Y�'|��͋Q\��^6��69I���X�A��6���j,�e��2�Y3��*61���uϷ�Ȫ��;HS�!YJ��4M5�Ve���٫	\��#6<��a\�S����d^$�Q��62���/�d�vg��^1�4�t����y�5�.�z������������we>�iU��v�JW7]�3}N� j�þf9V){���srb��6�h�g˟�S��wd���Z�к���ɰ��#A�ǼE���n�K�Ye{�7)���5h�P�����w��ɸ����̎�gﳮ����}�Sm/��ؤĮ��-�R��Y��a�Ɍq��޽����KOU�
u��|<���1KLO�&����S׼�a=��˧�yINd��}z�M��;�^M��KB���i�^w��y�o0�U��������l����'����]>���l�@�yRX�k�m˸�~5���e�t5=����-"�A�ͱ"l5��̉�W+S�%d�<W��!����:W~�VO�q��m��1����Oqڞ�������Әg^�T�d�+ui: ��kz�^������yIߋ�5���B�M�z<Ŏv�.(ˤL,j��m���*ұ�f�kA�&N�+n_����H|Q\��	�k'�kڪRd�)�-~튷���{������9��5�zD�E���Fc6C
���4�b{�i�zx.ј�$6 �Tc�$��~C�� ��	<OP�m{%�-��H��^�w ��:�Z�eu~[���Fϡ�0wuk��.����3��Z�B���h{\��(@J�l2���0xw����k���}?��C�Z^�#���
������������(*����(W�Ȩ���J���pB���mSSmKZ�&j��ڦ,�S2͵�,��R�KQ�e�5-Zd�U����cU����2�MMm56�2YV�љ�TԫMMk56Ա�����[i��LY[LYV�YmK3-SSV�����MJ��ڦ�jj[SR�6��5<U�ԫMKjjkSR�56���SSkMJ��ʴԶ��ZjU���5*�SV����֦�Zmf�5+SRښ�i�Z����զ�ZjV���6�V��jjU���5*�R�55���MMZjkSk6��զ��56��֦��5+SRښ��ԭM��MM�jZ���5-SR֚���j"�E�6*X����5-��j����V��	���i#`,`�DR� ��!  �GU-J�R�ժ��Z�`� B�U�!`�B �lJ��B �A��Z�j�j[j���U$ �� H� �A��Z��RԵ���mT�6�R���KRڪZ��� vX(�����KR�T�6�R��j��Z�jmj���U-MUwkWm�j[RԫKSZ���-MZjkSR�4AB! K�Q�B!20M5*��j��[SSmMMm3,�MMZV����2�5*�SV�,��T�EB0�H� n�F�i�kf,��J��ͳ5����X��c�fL�E### C�&����
7>��((� (��*"bs��_�~9��������0���G�����?��߯������C���~���������@_�~������Eu�"�
����@�����t��}��!�`����e��������l�"��3�����p��
��p~a��$�Y������
�B$Q"�P D*�[-SU*Ҧ�6�mR�JԳmKm5���Kk-�[MjT�J�[SMZkf�Y�Kl֦[R��F�5��6�ԛjZmP* �B
H  ~	@�"�H�� 2 �kQ�I�L֢�)Z�j+i���ImL�M5�f֥֔�ZY�I�M*ҥZZkSTե*Ҧ�-�ZZ���U��jmh�AX
j��J��}���� ����2
�H��G���/�?���p>�z��9���@Z�A�����������މ������-���X�?���Ƞ���ޟ��>��@@~�@_P�H=>���p��x�"����� ���R�����=�((?�W�g��Q��l � U�G�?�C�5���
��'�@w��#y�����y�0�=��������
�
�;�D?�� U��x|�z�D�+��>���x�ʃ���������� *�?I�F=?��R��"}���a����/�g���D_�|����M�"��>�c������'��W��PVI��K��$��A�` �������/��<DT����"��������T�)%"�J�IITB)H*���B��Q%P�(D�"B�HR(�	P��T�`"�$��A�J��!Q)*�)$�A$�Q) J�U*E"Q)Q
AA%�D��)UT��!$) �BD*��4RH��AAB��RUJQHR*��"UX�P�!!JQ$�Q�RP�T�  auIE)P��P��E�ClkMj���жj4����#m��eUk+
����-UV�j�T�mV�R��S���ЅEB�P�m��)RD�   maСB�
bF�qќI	�!H�c!wS�Б#l(P�H���H)M����е�YV�mmd����C%���P�چ-�@R�b�M`�UbT�)*��U$p  �j��
)0�*�
�
���2)ha[(ձ���JŔ��l�f�4�5��LiJ
�ڪ��6�-����X�4����Vڤ���$**U$n  �JF�acUT��d�VڅD�$�UI�HյE*���` &�a���L5 ��k5� )�"�d$APQR*��p  ��e��kJJ�R`�4եX�
)de)%)hf���mEL�CZ�6�@	�� (J� 	T��T�J����  Z����fS �i��hlZ2��Z`�Re
�2X`�6֍@
@*�[cL  "�(P�d!!*UQBp  � �mM@  ج h�  l
 6F  �X A
�  �L  ԰  ���-�TD)J�  ��4X�@   �0�  4ح@  Z0  �d�  fS4  l� ����E@�P��*��   ,p� �3Z@  �  ԖB�f,  jX  ���,+  6�5�  ��TH�Rj�UT*�!�   �P ;[  ��  ��(  Z,  �� �  �� B  (Ֆ  �"��JT� 4��a%%H�� ��LM0�b`&����R�� Њy2i�2h  z�"ʪM C5#`�d%�L�ij,&��p4�I��x��
�,A9�Cҁv�P���������K���[Z���Z����:������mk[o�յ�m��U[k�W���%����������N�&�Z5*��B��z�1��j�\��ib8�x2�P5��&k5r��c�V
W#ZcO2P�,�G��&��ɶ��3v&�J�W����a?��V�1��òÔf�ճ0��'Tɔ7)}D��hU��.�U�G�zT.�h�y4�{L���S�2��c��Ve[�ma�E��2����̺��ʔ5f�iPc�Z�u��M��i�<��
�.�]�6�t$��Q���4����j��X����
29W�b�Wh�x�<;P���^�N7a��#bOX��^��]"b$k��x�bj6t�Sh�:6���ݭB�	�94s�q�PU�Q96m6Fݓ��/@�*x�5��������K7cMۘ�� �R�Y0�u�kܭXRw��b��P-դU�Y>�
GM�U�t��YB���:xK��I����!�C� �e��	��*Gq̻�X�\�b���0*˽�_���6fs��4�U�T�3}�#����]l%��mM�� Z�%�*��1B�p<a1D�v)��D���,�4��Pn��M Z�̶2�,�Э�P��
t�v2�	2uE>�5���ε'CM`h�®�)u�M�V��"�r��\xɨ�J�.QFB���MMd(���l�!�R�������Vq��y��M01e��m<ʒΡ(��2�,V�ی:.�!�m8��ՙXU�
���h��dS*��Yvс����6(՝�4�1fR���i4�Ua"jFe��8����^����V��Ql�����A�DP�<B�4���5���3t9�Q��a�v��z���ɕ�������[�g-�n��Y���񳻰�H׊iv]��Q�3i�{0�Sc�n��=���H3X6E'���e�Z��S�����,�72���oT:	7�����l1D�*�A���W@*�h`l���b���)�6P�ܭB>:��y�}�v%�acE�/d�Cm}a�Uk�����8�_mX33�%���?n5�NM�#�r�c%md�RӻeH0�Ԓ�b��]�#���7&�����-	��T�z ��T /N��Mb�Q��	�6e]�g`�ƁǤ��E���֞S�S;����I���XUԈVf�XYe^�[{d-�*u��[.���)QI�u�8�sFЫ�(%��J���Xj�;��K�O)}��а vܥ�h�e�����`����%;�AJq�D�8�$�b�8n��r��Ct7�CJؙ���m���Q�B*㗷�ѮM�a�[���*헵!2S�堲^LԳV�I�BlCY�@Fҧm"�p]�4V]�5��T�n�ֺ[W�1�铀�:+�;	�q��5v��<F"�rMPA�q^X�)�Ǜw�oMq�0`lܪc�aٺs+!_	��a�Bɴ���"
��I�]���iِ������h`L��k���;Xw;B�n\���QM̧B�n̔Ek�������˨m3���ۨ^,���!������f5'E�e�u���
{X��$�b�v[���	6�Sfň!q�{�q�FI�D�� ٲܬ�e���é:��Q%U^����V�\^e�ɡJ�#NƂ^�kLK$8��9yb]������q�M�6[tS��N��6��h��e�r��w�s!/��6틫h��K���#��R�7��2�f��r�ee�Ǆ��kUfS�Qe�T��`hR���b,s,�.�V��.�ɤ䣪 ��{wB���6��Z$�.�F.�emk6s(�X�1D��b�zْItrV��0kT���֕�ߠ@�%���](V�ݲ2�i ��Qm��T^*y�$02^\��L(fX�p\�*����6]V&���
<�i"r��Ypv�-K]{>l�{tr$�e2�mEI
��7+3 vL�d�WC4�t��>�����J��v���+)\u�Aв�(v+��Q٠�2�o$���ҢU��V�P��F�
�3(�aY�d������S�(�L���C�S"���][Avj}��%j�²@G�"sv, Jt��ɚ���hX:b�F�X�ԫ�R��㼲��"����yҊܕ�k�UL�4�N@���XB�I:.֬�4\;�� ,
��^��,U��d�����B̐a�H��b����t�i�n��:XM��-����g��l�ڿ�����FD�7��,����t���McXv� *#F��mf:���, �G-bRi++�T�5��Z�İ�t3V����C
�{��������'�Pܫ�f���6�S�M+3�[l1�Qq��	�L�[�!e�5�iVc�w��g.��Ū�ُDӊ�fVR�>T�IT07��N�,��O�����I�Ҭ8�Kx����1tp �4CjTB�kn7�h�" J�wC�u1�̡�n]<r�8�̂AIX9����I���XŌ�n�`[�A�$�^�a����՚Ҩ'	Ԏei7A՝��QÔ�^Ԭ���ޢ�I[�@HK54�.D�ΰ�ق^ E�)]�X;�Ll67J�(m�rd�1�w,�7YX �z�m\*��
��ۏ\p�6�'�4l���ٌ��mj�I�vEp	*�Z�jT�5��(��im����9RۡG@�:D�kM�{F�,��{[j
PTW�v��$��iE�Hu�$��L��1P�xKm!Zsq5��Bݵ�"�;��f�QDo�%�&��d��sK��C[l0���sE�0��u�9ofЂ����FG[�@���;N��/Ht(h���V��lz��%!���N���O~Qس�WI�c�r��t;�0k�t��0���1v�G��*�sR��l[1�B;	y{6�Y�z�ҥ�\V�G� ���E
�%RVYݙ�U�s)Ԇ�d�2Rp��	�F����̧��T�tԲ�r}�Z��kbM�[zX@���6�*����Ҳ`�)�,K(��(�(�x��&�U��I'F�$�f��6�� �)4�2 �f*�8�W�����w�E�y2�	�������+2��S�d�ƕc�x! {�1̎cJ�1��a(ܫ��yZ��.�Ԭ�ه�Bm3u�YSr
�>��}6�\[�Ԗ�@Წ++�Ǆ �pDhn��݊t�6�'.��L��sv�&h�c��MB�0���zD�c婩PU��1#��*TIǖU�y�n�68�% J�dlb)3h�
�ݹ6��@�E]3�F�զ�.}$Se�N�-e�kC������PD� �Rݒڴ𻔲*�L@ik�X�)����mG����]��v:T�͸Y˻KS3uǮ�K.e!��V��S�J��Iۧ�[2�tM�ň"�^v��X��/P�(Tcsik���n	�j��v16�%Cée�Ѳ� ڃ��o45b�2�Ax���j=T�
{əu�i7�eD���j`""ř D:FG/k���z��+.�0��,:�pn�X6j7���7�
��h+���V
�3Bj��wR;� t��*yO6��:�����F�W��,������P��0����Ù���Kb��4A��9F�H��B�r+S�`��$j#C��٥��ãUKOY�P���$%��(�Y[Jm�@&L�2�� ?n���*�n|wS��@Sa�e�&@%�m��i�P�"��� n�R!L�
n�-�u^�M^ӄRI��t�]�C�ܻ��QB�e
(�aU�o^=RD�b�b��-YYZ�&t�����9sP�� �<�Ma�=�T�y�&�9���"�]X,I�C.V�e��cM�U� ��ë����m��p���Z�����^22!K2b5a�_�G{O ͵Ze�m*�T�����h���Z�@0���.�w�PD�D�:�L4�!��
S���k	(������qF	�1,�Z�`�u�W��6���	@�[���ٵ�Q���)6q�Ǌ�Xv�^^,�ҷ.��6�P�R�*}LZ���ĜN'�\w����b�k��3lE'{�kv5v�J�z��� � �P�[V,�X/`�oH�1���Q)�(\���d�X�6sI��c���;/*���]	���A.�X'ئ����9Y�R��Q��2�1V!Y-�⬚��[�e㩐FLx�7svf��k��u��FT��PJ�������+q��׹x�P�u. �۱C�FY(���by���7�b��Zuc�m��IRz���Z�)ҭ��,�����)j'�D��=���{���n�5G0#P��q�;^K[�J
�B��H�S
�
V�[v+��"��^�btb5��[�<"V9q������K*�taE�tlK{u5��Ѧe�u�Σ��
��6��֝���g@,�K&Il��z�tt4�tH�a��)�+36�K����-/�ԣe��� ֳA-�cv3C�1W
��"q\w� ���*]Ib��ݵ�:(�u(ս�On��f��9�u�+REi�N���.b��@�Q�C�~���o]�04��"���h]/�V�3!�����0�5��1޵��F��;�<�ݷ����7#n��l���sfmX'\�-�YW��+A�4Q�6n,��4rѥG[%�U2���Ome٪�%�����7P7��0���*N���u�-���W3cڀ��)���mR��WVj�;��:њ�2g��t�i��$��ht���U��%݅{�ml�:7S��wfޤ��o붎S�]n�s%@�
��,�l`�m�Sh���&�[�@!����F�֧��a�l��9��ȃ�V�ٕ�fMYt��f�̿���ǉ��[��M�:)-/-�t�/RW��:Z�ۡX�0<�Q�r��������l*�ʶ�p1lr��a������aʼ(j�LݥA����{u1�Kx�x�k�a�X`RA2�m�*�Q6���b��9{,��u�	�ⲷ�0nal˴T�Y�2Ďm���-�U��`+��Z�Ă[�_�M�v�Sv<�����)��$��V���cT�����jS0\���4*��sV-E"Ս؁ݎ����Eͻ^��)�ө�[�j6����j�z���XOЩ�E�e:�u�Vh$�KɆ��Ƅ� ��Z��Pdz�|��P�[7Z[��,�J�,���DLgF4�c�dc�X�L�%��u �&�z��U�P�u����3A%Pv�v���)K�+�Oek��Wn�vX.�n�o	Jdr��T���pERںͻ�\i��-�
�e�Kh�����uCL�k1n�6�WH�
i�80�`tRQ����T~�q���R�n�ZS�M��ct�Ӊ(V�Ŋ�I���$m�ܘ����kf�ܛ�2�cBb�VSj��L̬��Ƶ���O~i��5��\��xv��'��cRr�&���>����(H*�h<�]�b��$2���n���J9Bk�P�dw��հ�����~��V�(��ַ��3,;���!$C+J�%�J���d�q�-��:��;@�ko�{�h[��(3kS�q�Y�|��/ ��9��9 feO��̷��^�B�� p�QW��z��F- �������`V[Ko6"6�c��I���1#Nk&3h���h�]��"M*�Y�i34�ª�ݲ�<�1Pĕ*n^ȶ�\t�k�0cF4�!�#ϵfkܽQ�V�U,��8�A���?���:2�t#��ݥ.�9�"�JD�L3);Ec������"���m%����
�䳗mH�e��cm��6�֭�GD��)`
��ۤ�a�p;b�!�w��y�{�k(�{��H�bY���BF��n��w-nB�%��b�.��[j�[4%�%��k6��@�
�^�0�sh2X"��N�T[�+rmc�5��"�Ða��S6\�3`��;�#"�ZX�ƩM�W'�K�b�FvT���G.�b�u�ґj�8��J����:���[oIt%]eTń�%5�E�����+��%�XUJ��9`�b����&ԫ����{�AK6B�(�#�)�RV��MCN�t��$:�EU�I�a�2��pi\�H����F7sn-9A]�����},\��Bj��I�dj�T�#��wbELLp㡰�$uV@�x޸Nɐ�4�V-[7L����A���[��E}��5�:��ZZf�`�[��[�˺_���%:A��zqࡡ#)(D\��v�a����
X��v���m��&�$�Y�XMu��z���Pr��RP��B�,�ys$V��o
�Ce����i�]a��ʍV�x1J�Y^��d\�3Y�WC\ݻ*�z(
щ-�i^�jn'w��,u1�s	�zR�@}8���v�V[)QŸ4c� ��\�`L"R2nʼ+��l)�MRb�S�/�i6�f�О�ú�l�W`	nP����-���Z���B��V���#`�72�_rC�z$[�����8r�o�h���f���*����-}gb��BY�4�PA�� x�����[���0V�R@L(+K/hӫ�q��СV*3�mKO^�!qZv(f��nԼvhY��İ`��Jf��+�x��J֫�YbjM���^�ҙ�M��OU�+��X�/f`���l܉��h�Ql������J,8�0��z��MܽI*n����W#���{xsM�� 5�*�����]i���^��Ie�fE{)ϱ�e�ĢZmj"[��3�/
����)���:��BV�m`����^����Gh��1 %�;�
��'��k0�j<�d7.l�V!��0�@�Ӧot�#��-oj��vE�rT��.�ʹ2�޲��b�(�
W��|��t[*���h����r�DU�Agv^���J�W����8�̮7��{&�L�׻���h4��5��>��;5)�������.�� }bAx{��ݷoT�x���杏���X��@��a�$w����7�[CZN3ٍ���gd��91�:b3����!�[�B����r�4�f�hi�ٺ�K�y�����p��E[S�.F	����o<���V��H���w}]ܲm�k;5�m5.B"r���һF�˅}/�a+l�uCbV�e�|���+\^�qQ��e՜�����8p�.�xuQmȸ&tQ�l��pJq{WN��U�}5�1]�Y�Ԭ뇒�Yi`��bHR�IGL]�'�AG� �@�+���OU�z�N���� ���3��#���۵�9��6����{��vh�)�����}�Ùut���A��E�C�������\���:�`�-�FD��ywq�h���󢦥{V�U��V6Wtʗ�L�k,R�ǫ�9s�V@�[Yܠ��h�՝+�U�l]Lۗ����*��Z�7:���F�w��VV�L��ۉ�:fb��9^�C�vś��9J��l=�*䃿�X��N��.�8Ef���\������D�1���.��B�� ��'3>�Ml\1f6�pۋn�\4�:u|���v��U���'�ʱӹ�W��^b���l�Y���π���k�u�E���d�le;~��I������^uH�G`]���^�÷�8�������[]gf��u7�a�s���t�r�C�._��Ö����E�e+p��W�ΔoGno$��Gl�Si����u��$��"��
P��8^ܜu�[���ZDe m:	�ɂ�9.����\�5���Bn�8�N},���f�l����#��NwU���й��׹ E�n�[*�K�e9]�>l�v�o0����;4��.$X���Jqw2�����T�WJ�y�0�ԹJ��RάU����)p=�ϲT
n��[��V-�I�xr��K����V|�q���O��GL�V� ���T�0��}��\��ѕ��&֛��-�\�{O@ʣ�,�Y������5Z��e�cq"���ʽj���8♼*�9�h�g�R�D��� ��d�+Tټ�Ч\e���!�g�wsm�Sw҉����rH@d#�� �/y�5���ڼ$�b��[f�v�}�b�3��}t��������dm�<y���v�Π;A��G`\�_.���{]��
9�� -��4Z��Pe�Ɨn�9��o��X3,��(�%� ^�W�����*�i7��AU���S��ӛX� 5{Y��!��2.�Y6
v��%l~��k��h7*���%�[y�z�O�Qa*	pRּ�Ѧ������3��A6�m���IU�+/���7��49�'Zޣ��Wkg+@�U��Ӵ@rʹ�K"�%W����J@�(.]]�iM�j��+\1�mi}�d�Zx��(����<���#�o�k,E��:�%�Q">���i��U`]"�B�<�v��7��b��ųѴ�muZ7��QR<�4c�|!t�i<�:qp�]y��v�^�f�j�=ǣ>��ZŜ!��%���P�U��_M���P���2�+��;�5�z�]���:��6ض�#J�"\�ܪd|wwu�ѩ.ɃEu�sj��4dgu%ZV�,��x��d�uau(�gZ씝_�N<�|�g�-�M�1���eP�n��ð��Φ�6J�{n�q
9�T�W���侷��c�����@l���b�(���m���m�{tV�ݙ����J�ި�	�����.���c�g�"i�m��a͙5�oa��PB${��W\���G��,]$�nWn�#9�Ҿ����cʏ<}�+�r��սF��vͭ����@2��v�<�=���+pk�/M��mE\�3��-���ޛ����*[�q�`]�[{W\���T��TivB��nF���Y0�u��ؤi�}�����R�G�{���:7�N��Z�"ƾuJ��Nis�O���sT�_U�è��q�5⺵W$��7�/�_2|'X5k�j�$�o8��,L��/���	{J��و�}��-|z5B�*,��k.�>9�,�`��37�Z�,V�&���R�|X��nN�.�^�}ݍ��c��ߖ@���K$X�Eܷ��	�������JTA�G3z]<����Pg��u�kS-���X����w�+͍��gGb����	�A�X��գ��4�f�KD7��[��8*v�������"�����%:K!��,	���*d���L��^�e���q�F�RwI�{&�9Lh��x򻲑�yH�Q�U���r��Nߓ�qͺ��*���3(@�V�Ji44�T{�!�fwcy8
�+/�:[��w���7-��u�ہ�E�����v�S9�iO�Y�d%����dA(g���y|�l��2�wj�n�j�h���l�E���ݧ���1�nvs5Xޮ��ueV���W�B:��j�5j*i�j�>�7V�ty�:��ꆙF���fZ�����>�a�D)�N��uR�$��`yf��v�I�|\.j�v�]�{A�#��i|�Tm���j$^_(v��uϰN�|���N����������V���nvK�˔I���]�1����� $�o\�1��c�3�E�F�E����T��uڄ���F+�.����M�������k�̛��kSxM��e�qPΰwu��w�mD�->��^�����kT99�����|BG?���8<��\Ԧ��eȝ�wU�zm\�z�;�g�
���bԴ�Xo��Jc�N�d�z9ϱ�̾Q�qҳ��nmflj��6��a�9�R���!p��[��p�f�M��U�7�A�Vv��0��=ű�$k�X�}ۜ.��ʈ��}��Wj��>:C�DCY���P��<�S�&�nk�;4��_r���H!�ΨaJ��Wb:(<�ʾ�X��ۢW&VG��1�ڷ6����b�s{u�]ʷ3�ʛ՗˨���1zPY����Ѣ��ς��/�Z�JA%A�ڐ�ٹ�ش���A`�[�J�JƜ�\��Kb�G�"���o�9.׻"�%��)PWw����E���:v&7�Ze��D�E�W���6����'Sk'�=��+�#�k*oW#���,�
x&te��.�c��!�Z�j
eu��x饱�s7��7�U�V�\�2����uJ�\�+x�,��o8�����b�6�j�6�ѠD�oјzi�`¥!�j������v_n�X���k@�E�z����t�=Lu��#	�֬h�7O$��Y�6lV	"'��7�j�v����VK4����n�Օ̘�
v2.ޘ!���X�l�u;.�ܲ1*���2f��vyc56��X������i��^�Y'H��ThN-�YKP�|�pD�eǵϮw.��ާ�"Q�+6�X��^)�R]�{����"JV�R��ځ����A&뼭���O�v��[�k�>�n[�jm��3�ɭ���Z/OɷEIXc$5���D?������2v<���T <���w�Xtu9�H�����
����� ���PS)Z�x�D�3���b�{�tu�i�5�d앏%J��%e��[�z��΋��I(�'��v^X�k`y3R�:�6RΥW��ق+#6�{�8w\^�����uX�4�-D�;C��[ꂲW$�58��ԋV1�p̷�ͱua�3��rɂ�p-���t4���W�g�n 8�Llۮ*lGPY����5N�����b.�uj��.'�0t��B��_M��킷_]u�ʹM���
cL]��{X���eg!�EhP�����g5�6l��,tb� �$���Zc����@�zbH�r�����Eȩ�4�SY��y�}����Z�ᄝ�b:�=�|�g:�&u�l<��J�xSP��2���%�K]�{A��w���2h��(V�V8�6�&��e5��_uK��,��	iR�Hl��|s����tb�yJ]��F�AM�%0`�g���R��;�h�;w�w5ɨ�^7����P�5b��m�=��E�z����V�!F�t����r����	thW<؞*f���ы{�ϱmJ9�><l����C���h�A��Gؒ6��\�]9Z6�[�����On��&}���a5�+���=խ�*<�+*��I���4�F��@'C�zs��N8⮤�8�Ԁ+���yt]�	�3�F[`T�}f�.�z�8�O{7���z��a�d��O�M��c��E{vz�w��w:�S�/*����`����[�;e*�P�r �;Q��PϷ$��z�ٰ�!:�s�])NC7�G��r�x.Q�=.V��JE���[�:�AO��ծ��l�V�p`��ܨ)�Q�i�>�7Z3rd���R��Z�LCap]�hK����K:�U�8fic1�}u����v��aЩJ�{Lmu�xp�N�ݡ�VjjѓCT�p�H�S���[�l�E�s"��F೙��PEd=�[t@��7.w(z�� !]�(ՖM��o
}�V���E҇��'(J�0��f�%�VW+4N�KL5�[z5y�jYˊm���^�#!�<���(>�0���-�͍�����ZjS��Z�ao������[:�ʤ�S� �̻F�əG�a
��2�]�Q�V��"��Ѽ`��Ǒ���ﴯ�qWk�E��)�Ϟmۏ�[4���^P;'p�)˻<ͽ�I��J�o�ݗB�@���� �֜��ԭ�����,ys��S�;t�uv27*1BWvR���5v����)pS�l}�>�k$���1TN_�����E9rT�m��r���
;�
����:�j���^}�`�vn^:��d�Y1��`�;�`��צ*ִn*u���U���;�|�:{P#h��q�髦s������bD�PlP�>y���΋U1۱
�Κ��+��N�'3�Ai��[�h\� ��o�Z�d��kF}���y����;�9Qʾv��=D4f:�ûA�T�`��K]
��r�iG�y|��I�U���=u��;l��u�*��+e��4�.@7�7k��.�d���R��+�P�Ǎ'�D��`� 4�sz�����8d�{l���E&���#qJ\��S={D��A���ŧ%m�Uan9�o���ʲx9�IJ�Y�p.����b���:�%w�ܰ���N��tδ�h���.��'U�܃��r�y�vJ3��ݺ�V�<tF%qɷ��s��K�smS��V,"4
{�%�ٓ0A[��y�夆(S� �R�gC7�4�v��6��%f��0"��Y�\pt4:�<�x�1ݙ@a����G�6�$�t����h-��u����uwR"�p�̵Y��9 ��|�`d�Z2�Վ8����"qȄ1;�)��[�Yc�h:�6��/fX�p���;�#�2�ڲ�6'v�ԓ�2�y�ǭ4v�uZ���cr�]"W+Y�5r2���_ypo(�wI8f��^�:�s�AEc�wM�Y;���X�z�g�r�7�9T�sn���oW\EMּ���9��[y4�3�I���
]�l�0�f'��c-��KWf���,��5J���@�t!����"�!)�=�&���hݜɘO��n�Db�V�2*���xUN�F+�Z�v��齕��-\�0*��6�cS ���w/_h1����>��t�^���,ɖ7"��vZ��4f^�v�Z��B�Tt�F�]��w̞��)4�#��V^'K5x����ͳc��[$ ��2Q�����Yڴ,�ؗ��SB���ϔ�B��p�K���F'��XU�o�SvA����y�Z�X��k��4�}T�l��!��ܐ{O9dS+�#�mɅ��2���e��82�t��"�m��	�d�n�7�����!��-g
8��r��ua�����:�w[�x���@Y<xHu�/��{�Y oli�ݤ�|H�(��"7�����鏟V����;w.�iby*R�U�o��;�7����<�C8v�Wϵ��9�*��a�}cob����\��]�ݘ�� z�f��*(�m�|���8�PӱѽݩZ�P)�NG��;l��p�wbݗ�'a��1%]�5�K�u�v��f)4ѣf�[�um�ږ�c�)R�!����jmZHoJ�{���r�Ht� ��zn�Sf�x��Bӊ4�&��Zh�v���A|q#���x:ݥWd��uBX����]f����[�s����F�W*���Nm�`s\s`�xQt�+�h���HZ 	��	�wa�|讕�[�v��	̝�Í͙��@qYx��8�^���~��)@��';���7u��AK �� w��<���ǿJm�4�h�.}�r�˕�ۖ�K)�p)* &ޡ�f�������S�f���:��(�V>��إ����t^�b,�e>����-���.bPcSXMs0R�kN��\�t)��5����e�%��4����
�`܊���ӆ؅P�k�@]�"���oN���'h:%��Lc*���I�c+_��E澥�<aCq���w�cd�L��A㚡ygK�n��p:���)L��J��❔���oq�X���Χm��fW1p��-�\y�t�ө]3\(^�*�eGL�y0Qc)���޳�uB����9�Wl�z~�FN$�Mͻ�㎮�{�±�������ӛ_@�2��"���۩�` 67���d/� �����b��Z��nq�F��4Md����#��b{���Ժ��y�b0r<�����HL	oM��kM�V�k���ڝ�G݊ͥ���Wp0O ���ʡ�o8q{��]8�R��ݨ��u�i��Le��,A!��!����U}UUU_}�_U}�}_W�|���~�B�e�WR�ZSNǸ%��)�[u�8;oYwZ�u��k`��okn��0tXww���Y��'�M�˥:��{*�G�p�ll���C�te'�����/j�9r��o,��7D�gr������)��Q����{[�{GC��f�Y�r�Myl�J�y���.Yv��{���!���d�'0a��'+F���p�:��崨9aE2Cu���z�g���*�.8�=�S�����w62$�_|ECO��}x(��Zt��U�g�T�V�m�f|͗��z������櫠X��h6��xK"�y����Sa_mՉO��*Y�=Չl�r���-�G:AV7Hk{'^th[�:��j�A��UF멺BQu �=[Wsi���"����A#wT� �$��]��v�-�8 ��_lclT�ua�Q��u���WDJ�I3�_^ᰚ�:�Kl�jL�
嗧�Nh�\��N4a+ D�<I`WǌLg8�f�M.��Hқԭ�'��1�X��w����T��j�Jv)��Y����8y�wD�}��W]�hS��YpP.�v43a�A�w��}cH�]a��(�Қ�V���tE��l��*������>R,b�*�]ʴnQ�4Y����2�ț�R=��L���ϵ�)K���rݜ���L�.�D�z��t	�A'����l�tmA��L_<���vi��ъeF��⥶�jZ:Ge���AV���G�j��hͻ#:���7�o�35�b�mO�һ�Z{�gʭ��1>��wJ;�P�G*u��q=���/u�(�a�R��A��|J:]�CjN�.(t7n�)p+�����0�i!�7��{����S+V��w��Y��e�`oCId�:�,G�W*¶�S���mXi�u�
Z���7ͷ��-T�L�a�n�O3�Y>ʙ�0Ǹ�	�&�*z�
���f�2K��!�,�;s�;8����߳[�kl&鉝�5�{�<N��0\¯wgݺRr6��⻖�U�/��ꎶl�ح3�gP!��<�,pл�ufI�0�U�J���pa}�D�Q<�tC����r��Cfc3��¸(�j�C��VgX�uΏn�C�q12�'2|K����+�P�-9�]�|R�ky�ľ�N�����-�5w���˃��I�"b�eY���bSJq�G`̜߰qʊ]JV5���/R��2�)֬�=���n5�ja�Y�E#:��Jb�]�G��0��X�F�Nk� �\n�P��K����2.v�*Շ���z-h'��H�WLwu��%�Yt��;еqS����g��9��(�w�b��x2�Q��(�S%�,��VU��^]I�'v��U�y,�+s�/h��[�ʦ�+��U�c�fJwp�]QVj�B�#2Q�K�]r���q=&�U�:Zt���ժ�պ�<@�����X;i����)T[N��/��묺u�tE��_X����W<������>H���̺�(S*(�:t��U��RWۊ�=;z�lfgR�S�A�H����ֲ�xtSCqaJ�We[z���mtR<�6����%`�̵ԃ��{�s�s�@[�����Kj<@a/����*Ti�}Kh���O����z�n��v�l���{�.�˫���f�O�0W[-�9b�j��{��+���w��/��ܽ䱽²'�s�q�ĐS�W";��ݵ���uv�u�ɕM�G�I{�8�R�����C�k�VR�{>v�7R���U�}3.uc�۬ۢ3�v'GҚ�
�t�L"٬e���Y'�q���-�����`˓��.���:|�Y�̤���`��fj�!X�u�1*���p$=��"֣Z����ΝV�#ֲ��)ӝ��̺R�
��e�L��vΤ.�Yo��Vɽ��R��Sh��o�t�v�CwI���[Z+m�4�|�b�m]�0���8�]����l^VՋ���[��N'%��x+y��>z0��y��\�Q=>��Tw�	�õ���n��_7XB���e��u�E�Fi��Ұ��8)po��B���hb��7ܢo5�\J}���n��.��(��2b�IH{-Q�}��9Z6�b�{F�|����A1h��X��2Z�Q{�'�o�4�K0MZtVؤ��K]�#�r��*�;Pq��8�.�E��
�(h�k/u}�rx:�qf��q�ǅ��6�_4Wb�LX�:��D�����Nȴfn�Kh�Y;Mb�ZͰk���Ϳ�t�[�Y�X V�F��<�;�(��EQ�1��uX�gKf_����mw�=�T�GV�Zh��U��u�j�j���8�KWְ][��s��J�՗t
�7��e��e2��Q<�o��s`�<Dc<�N�3�m���i���e�u�X���ڔ�c�y�Yi���q�A������W�Q��k �M��C�G�oh�uy������)#��*5k�#pV���!OcR�ᷦ��.�ب�� �yc{F]aX�V]���t��c��[%��$aЍ��uTJɥӻ$�\z<x7�ךlz��)�WT.�B��Ƭ�wxj�WV���e5�G��(�%�D�R]��s^j��c��b��S'��̮5u�EL��.ޙc�_l�RYF��X�^]c��RJ���k�5p�\��)mB�yۨh w_C� �]#�sZRb�v�]�t.b�9��p��m<�^c�VLa]񜥽�sh�����ฟglY�*r�h�W�FW�\�=5K;��ٚs5u�(r.s �RN]�7����ac�v�V��Չ��C�!�,4Q�� ]Y�^g#|��vl2�&wK��ǂ���
Γ�[�촳vIG���Z;�ֽj����[O�! ����rV]�З��1�kze�q�J���"ziô�
{G��b�bl���6�M�Az)��۔�RW���4!Jt�����(��Wt��To>u�����0W�F��Y���"J���{�ZY5s�眕NSëU���>%<Uݵ������R7��H�o��B0��[�-M��֎`Ϋ�-�HϰY=�i��d��k�5AL
�y��X5:�4m%�p�ѣ�։��p�`%3
u�
���rA]�7Ye�gX���hmݱ�\��Rp��ކ.%��s����hNK�2Nűg`���W"����� ��uK��f��oz�S�l��ƻd`�����0�Nd�ݑn)K�-��^��V�����@�/f�wSa��g.&��v$��	����*�ڐ{�	,jB�DZ��˙5R��Sn�lT	u��7QV��Sj#Lq���wf�{˓�d�%����Q0+P�K�u��F�E�A[L�cvif쭻x���7z�W��������e��*t��ܫk32�`ߵ5B���ըs	�3����oLl>��4E�;��7b�L�J�li]���	����l�$�M��{�g
�Gn�u@o���mK���Oxg:�Ɍ�>���ekHں�a6�3��F?�����[�j�ʹ�vo�⺼ZH��n�Anb\�<@��B���؜�m[�wZ�z�v7�V� <z+���rΟh��A�Q e�8�,�-�$�#J�蠷��ũ}�9�X��]Ύ��	��g�<:��"vp�9�Wi.cNb�v��YB����A_3��ֲ��7
�q�Í��;xVf.��
�B����u틳W�0�[ή��ŒSVb�C_t�K�A� *�ϒ�xA��+rk]N�vnv-= �⮕�JS"�}�]e�\��/��g9	�-��B塁SQ�u9/0�b�Xn��24�ʋ���OW]u`6�9���Ȱ�q�x��0R�!יw�f��(���C!��mH�QZ���)��Q�-"��z�2\�4��Yt����ֲ*��2�%&"�1$vuшӉR��P�
�L`����]���Y0u�<�P[ĭ�|r_R�X�W!2�U���2r��ʜ;�b"�+G/u���N{b�ĳuI���7I.��q�]�)�b�T}]Ck�X�;�l�M�tP��J�\=����� ~i�A������z�šW�
�'�x��pz]�O_?�:�sin9F�޼x%���΢VWZ���q=xx�eo�c8Y��(�$��B�{0�H�a�¸�b��Z�m�ԏ!�K�;;�e`M2�S|k�ѻ��IG�0ΜՎ����*�΃�ktؐ����Ĭ�SsESs�0V�9�^�}|F��B�ĺV�MN����}@�h�1#�f�T{�O�f�����>v2������w�h��d_CP9Ġ�f�P�p�$�Ws9]J���jK��=�)`"b��P(�ae��C`�+6r¶�d�,�+zFf�­a��2�Yȱ�-�8�M��Jc�p1M�C��N��|���pw�Y�;��Ɂ@�I󦭮��2����%��˞�˓r�N�᧭��1��:`�q�x��Y[��ێ��C����y�-��X�t�b�<)[�b'�ٜs��h�Ez�OmT��6��Si�2�������&�)+:V�����trΖ���X�y|��|��D�Y�/{~:�/]NnC���֮�$�ԍYY��W| 8���i���l�]�leH�����z�����D�o�u��s}����c����Cxha;��+DG�+q�U�fң��bXe<�+�P���W4v��=�d범��,S��]���]��t��Քž�ރ���1�C
���y�;�㳴u�Z�wU�{��c;�5�[��-���e�]t���8z޹�UZGT�kQ4&�P4b���A*f�i٥w��	�mk�ﻖ�l�l�vwp�b��N�
�w��~��fc���yړs-1�E��ov���}����7��'e1��P�4�-����T5�u�`K���ip+*�e�}A7O(�V��A��x>}s�3��I��J[�^�B�x:6vU���(���]���6.��<��[;�K�̹M�e��j�u�y"�q``�}���
x�b�݀��H�n���������q�(]�J�d=��6�! }]k�*�|�������2軙���V\��U3����lwB�VQ�y"z���S�`fw������!�
Y�@U���0f��R����ݡWNQ�5��"�� �X,^WN���k5oY��q�"�[�ɫbVS���kM�/�]��co�=Wbbc��������@���+�Zˡ��Q�۲�%Z�+T�y��Ki�b����m�ܻ��2z,��c��^�3{ruAU܋.qo����O`�32���^���ӳ����Ѐj��]V��KcwvT���z�iZz7A��զ`����ȻjG'���Fs.�l �*:tW����p`�N�nwt��4��c�n�������u����*Ԉ����'��ML��3%[�e��N�"�<�ռ�rSW�cg�E<�YU�f��e�Գ�V�'n˕zBȫ;�O$�:�U�RYa:��9��nS쾌K�@�K]\#��	J�՚�S>��}�+�h�B�_@�(�bV���j�pt*�s<j���5_3��V�5j8��,�6���Z`3�m�Z�P���Z����u��\E���k�nV�N�֖�ä�g�Y�L�r�kXT0� 3Mv"R�v�Dj�{�/]dL��=���ٚS�����_ʴ+EY�+�*A��t��{�v������`���L��6i=�X����˥�'%��z=����d ��N��[9mқO��,���ݵ���_J9�"��g>T��Ug`�7S�]>؛���1r����X�_uįf���7�k"C2�.�b!n�NnwL��5����ֶ���L�Ķ�Vl�hml��������Kb
��C�>ʊ(/�c;v�-�R�[E,�Kr��+��CK�	Ɇ�yh݌��.6sOH\z%�f��l������u	��rڮ�ᅓ&��'���{$j�K��"�L!���q���w`7��E�wh�k���{"m�ÎwةM�(»sLm�z��Ԉr��2��X�Rk��9��r�4�mM���4넵;n�sc��1D�Ŷd�(h�5M{CS�p����|Ѥ+7�2�{Qn����u-.gh'�"�u�xv��#|�i�ZwF��Q��w&�D�������.��v)H���E��%}��]i��h��Cy�tlA�������\"�n��u)on�G	��l��N;�H-���ղ▕t�g��ձf�Z��O6,IS��kU�bSU<��9w5N��� ��+�
��i\��s'#n��}�i�Jk�[�ND�wi��Ǘ�F���r�5�i4�s��[6K�[���ep�E�k���C	��dIZ�Kb�y�g@���t�w�
3,��f%�/�Ws�Zm>��Ӯ���V�Yar����>Գ�GS�x���\㱅mnI.�}��4�P��R5f�g��w�]���L]�w5�:Ah[l(�n��F�U��P��ͼ���p\A�S,����WY�����$s��;�%vU�ۮ��܆�N ���Ԁ�;�Y��T���ᐜ�%���현)�o�x���Ә���ݘ�x\�N�{�Es%!��4��oj��w�=G������[;"WO���8�/�G	��72	�c�5QS��k�N�}��м�|p�v���\�3U�D��i[���e��F�^�bu���3%��
��)���aL`��Z^�#Y�����FQ=���,q� 	��Q⛳���P�����g6u��D��n&F��Y�zҠz�0R�����s��ц��<��}8d g�d7*&M�n-�3��E�����{w��+��*Wjt�}ݲ�3Rf��G7�7�GDj�r�v\�YW)s�9��(�^�h�.�:3�T�:�򌬓�c�D}�}G�}?}�R��(���üR��K�U���-źx��w}X2u`�,U�:+�[�mW��xI��K[!�;V��{��y-.ALvѫ�}Vt�>9�l�>\�d��:l�!�d�&�`]��>m��Fos���2:�硊�Z�(q苖�/�����Q<�'ML�]C�V�3(�ŕ0-��p�iwmdU��U�&)}���VL��[�m��[}vsD@��:O���vn��;/"O�p�oq���	n�r��,n��s��Z��,v�⣛st���4�=Y8S���IZY�a�@<�W���+�)�%)6�t�<�V��t�Q�]2Ō���]Ai���q>|ͅfq7ʤ�����N9�y�'o������Yw�Wm����؎�⎚�*�љ�A��F��Oh��q^�L]�m�F(����5/z����w)��3^���A�ɼwZ��DM���汍؁�|�Z7�X�Z*Vy�w_K�o��4���I�e:��r�/�T,���;�`ӱ���Y��ŵ�9� ��E=kPЄ�L�\H]�$:��\3pU����ыn�h�Xˆ�a�o�v�os�"VkG��K��Z#6��j��q���y��ę�Ω�
��o����2`ˠ0Cqr�݈��)�ҊS�O�n�9��8��V��e���@np����啎;�%  )�����P�������.�"�(���!��G2"�v0#\��A΁����wn;���wss��R4�T�+� ����mѓ!�$���t��MG9�(�B�$"!�������2���u�S-��E��D���&	��S!���M�˦�%wtr�Th�hĚ�d�FlFL�# 	w]�C0I��΂b�9��r�]�Г�d����s��# �3�(s���vawuw]&��Hw\D6����
s��nC24�:SI�D�a�0�%��H� ̤��6Xe��E���s�%.�1���\����u�D�H�2r�(3wp��"��� P�
�|FA�h�Ĥ�������⶷re�������UԷ:؎��Ȥ�Ļ�W���\ޡ+���I6;� Ҷv����ܹN"wPf]V���A�����
�H�T��/����0v.k"�&@k3)����~�sGV��!R͙��w[�����-��S^"��i��v��o�Z��o�8�7���p��\b�����q`s^G^W�?
�-Է�?����)k�'Y�`N{}�������jq8*9�|/>��-O�,7���*g)���Et�E|\�c���]GkF\l�z�Ҽ3�UYؼ�Oy1�}qC�Oa#���P�^NoO�j�+;�88Gb�	�Q�X�[(	��D
����~��Y��������Ȭ�"{��y��u�cك����g���8lW8�� �[L�j�8!L��n�B�ՙL��R�]��n���`��;���z�Ö��a�l�X�����Y���@	y:Kʰ�k{��G��#��r�ޓ�oO��z��P��������9��~��NU���=��2d�
��7)��ٌ���9���[�D�9�7�+/nh9�����`�}B���JJ
�;���^ �[�H�
&��ٸ� �YX�})^x��<t��r��J|2WV����E���wo%c(YF���sDp`�qvl�=�;a�Zl�aN�B8��ǝd�؁�n�9=]])
Ãt��w$ӧ�f�D=G��1v������3)ߍNW��l�p_��g��r��4��k*����]@r�{LJ�|��d�n8I��V U�ս��b�J�����l�U�/i�����c"aW�#w=ޒkg�}�g�����M��o0CX=�n�j�4 ��$]�9��ԍ�&���m�[)."uL�ݦ���v�1b#VM}FFԧ}� �����Nd�R�"	�31v����5u[$��)*;���
J�+�P�:&ۃc��Y��aY��q�"�����P��2�Cu�2� w&�E}n�� .:]��rD��?t��{(5/�馢j1��T���)�<2�
�IS�0��(���������ە-���%MsI���8�#�(Yj,sS�I�b1ZX�2J:C���b�꯱�����.�_1�LoM��;ޞ��b{��~EbB����j5΃50��6�ٜD_�a���uB����Vfo!=�:f�߷`�4�Ё���^aSo~ڢ���R���]ۼ���J��r����*���LsPWP:w�VX��x��]��a�����)��o���Q���:�Ѵ%��SM�xk@-!z>��+6�pϻ�-�J��%������}]#�G����;�ԅ�ӷ�ś� F��v
��B���j�r-tf���̗���Jx4c�d9��s�9�S�S3�c��>,	����a�Q�*9D�1_ v�Or�Z�D=��U/c�����:�)�r��;��t��\B��O�/Ҝ>�X�m�t�J���vz��LT���ΐ�>eJ��,�G��Wz�s�Gb��_7�^���X��D���*������j��q+�Y�2�L!��7�/�Ι��޶�ڠ�6�,(6�M�}�r����yEս0A���[��ً��Y��U�\!<5�F���0\c�h�;���U�+s�b�ʙ��|���jc�
sq.b�D�Pҕ_[�G	�F�7p�
�(���1M���تzwqɈf�T!A�,��@Jj�0G�pR0&���;�]���XƎ?�[�B�����Yi���8i#����c��V�Z^THQ���#�S"$��1b�lkt����ع�[���Ə[��:�|�p�,�{]�b��%���a`��P�_M�"��/�[�]�V����mhw��S�8�nbOIE�S�� j���L�Pj���8�1{,X4��+�0s�@���Pw�R+Ps�g:�*�{C�]|�����rWԨ��1g5��N�'���0��.w+�_ǚ1ѥi���f��N}.�;�OH�Ժ�<�V���9#~�
l����Q"���%��1O�w^#�]	Sp#��������ED.�Sz�*��FL�Q{�xOʟ����'�>��:�Lwy]���X����%�հ�-!�E�Br��K��M`zs�ݨY����cɄ�}�t��J���\�r��$,�E�J@��`���l�y�*�|�����4E�V��C�f6����l,��3f���[�\�W�s����/��5�4���:{�r	��p8c��3~��
��dO�U�q�e�����ӣ,�푮n8��EDwK�0Kޒ�2₳�a��rwN�ŧ��'�浽&O�Nτ��L?�P�U�d�_ tP{{%��F\_T�9¹M�^����z{�sGt�xň�aQ�����f���fBz],8��;�T���3r{5��j�5����l�:/�iҾ���u�9��c��阌��ݼ70p>�����������|0O9��cB�}�`>�y�����c����xn�솕�J�"Ռ�צzj�ٌ���fmE~f���n�G���m�]��ɻ��
��u��oy����;��\=�i�v9n�MЯ�o���Ws�i��0uY�b���}��I���G�8=(n=�̛
Ut�{�K��K>ͰJa�.����;�8��캽�QɎa�zs�<!ņ#�S��s(��������.�e��3ʜ�*��\ܪ�ȡ4cB	�C��v���
�����]:(g�1)��@F���Z�]�T�U��
&�t'����!�B�2P����H��á��*t0t]+�߻��ې����$��|gh�_t#�Cu�H�'B�q�1�
�jB��b*������
���S4{��'f�̢��
��G�J6��j�v>Ֆ@�.��:ı\���r�>i���}�����D m7�,�t������ᒮ�u5�/�=��l���5ۑ��mFcT���V4���h�����z�� %w��:�^c*���ʻs���Q�j]�
{s�b�2��l%"~���1_$�M�U������:����9,d$1f���J����ˎ����Q�:�Rwm�1�u�\BE��3���5�Q�꼈S�̑1~�?{��/��k�\%�âP������pS�Gs�`cUu=��B�TOq�W�'9�FnV5Ϲ���r��z�	��]��-מDL���E��l��
U^em�\l���k7������4���W�0Q����*.5�5:�AӐ6����j�W��/t'6k*��	�Sc�&����n�pu�)X/l�b� j��g�K�H����ZR����y�2� /���9 ����u7����U�F�ruv^!�{���%�_/w�.��:������v0�����Z�?-GLO.
��ggs&�zb�'�:�t���.5�O�Dp`��Sp	�u�V����'(��ݫƂ�Ȭ�q�4\N��XT>ڎ�1���Z��%�����n�j1����UwJ!G��;:~�6S81��i���U���Y�#n!��d��V#��;���KLt����7 MW ��x�|)?+%��� m��r�2�c�c�kɞ�k95Y��޽�YN ��}g�f���=���08��
���]_]F���=Ġ��O�f��xmN�� ��=C��;��B�Q�ܲv���N����������ج%^D3NJ�����t�>V�LNΤ���K��,C��<n��ݙ[�U���-k��c���!�������>F׭�����E�����\K�b2�kTI;��5�YK�O	g��I�sW�6-CK6���u��7$��m�p��<CtkU� \	3��U�{&�����/g�ߵe;e�8�N�Y������XΪ�a��6�vF�^M���3��X�6a�%-�ud#�p�n��z�j\��bH*	q�/~0����	��t\U݊��n����;�pQ�*R��qs��sʲ�R�䀡åGmd�N�t2[2��0jf3\mF��d�01��Κ%
�t�1Q	:��S*��md���K�M�k(���{��r}vd5�^�곖��K�%P�*��;�x��m��)Y�<�IYHF�4g�	�R�d�q�=P��ۻ_^���3���Yc#�wn
j�I���XΔ�f� �xN��a�_7 `�@1W�vȕ��-,{R,��wT|%�>n�t�)�m���T+Ɂ:�+��\��׾t���`{�hf^�c�xG����z�.��r�ڎN5s�+�ylV�E����;�����ck�P�j����R�����bF]����;2����W�']�9��(!Q3��d�q\H��]M��ꦎ�{g���P�\�֓9����-"�D`�=/誰(�,nL�2�<�W����}/�:(bͨe���x{q>�Vmh�b���a�R�U�΁]�<�������u��}�/�պ���e¼K��\�*���y�u����t�"�7����z��cE�h�Փ�*.��]��+pP�x��Ek��}R�)��|��S�;O�\�z7U_Z�*Z�[�N��9bKT�g��'��WɊ��q�%�s9�˫�{��m�3�fؘh8��-����t|8��&'p�j��p����4��$����Ƣ?5G��g{˞���񲪚�����K����.�9��p�:��<,��!�Z#��ho�!K��T�Lj�y�fË�=۲���v>��T+�3��nc�!q�Fx�ȵ2���&��x-���c6�:���5��a���D���.��.0��nC�SJa�T�3�����r@f�gG&ݹ��
�2���
�A�#A���0��D�����Pʂ��L%�h�N�RDP���%m�<��"���L�@u����ڲ�9+�V;'�T��g�y<|,WP�*�{$>H��ofl@���ѳ��� o���VZ�ܶ�ߘ_6�������K+�7��Y}��m�s\-�%�B���?��Qf5�#�U����M��=�C���꩏���8��y�A����zJ��3=UA������gY��g��ꯩ��G>�J��r���ϭ�ay(�~a�m{CId�d��B1���a��#zn#�~UQ�/����N5�qW���+�rF�{!U�?d�z���Z���
��j S6w]�'�������U�ܓ��ʕ�O)�ΧG�S���h�V3�3��wBN83�� �o�]����wZ�<w�W(%����H�}}�sxvt݅bn�ɪK��B\��6jj�E��_�0ꯐ��Z_ b�ٌ�t*��s��f�Ɋ���_q�@�5��+��R5k������B��w�� B��d!��a�Z���`[9ZiP^�2��V�J#�O��;P�D���L�
>�u��E̱��t�΢�j7�lT�k�,�E�]A�}Lp��^	���+�@=������`UTg���py�ug�ӝ4ik=7)+��<���i�����b*Ӷ(��w��ߩ�&7{Bv�����x�ҳ��b�E���i�p�q��?h�y,C�.J��/]M����X��/;�T# Vy$#K4��<����:����)�ǅ���N�0�J���Bk�F�;O1%W*Llp=���<eT���t> .1pj7������T��ú��J�{�n=Of�I�8o2���)��PZ"���Ղbiun��a��0�f�,�0�E&�]v�Hgs9T,�E�{HA�ŀ:���Yn�2!�����~���c�n���L/�i�5���^�hɘ�B���,�2���mH��v��X�o2�V����ەw+j�c"��wk�\��{���(.{��=�	ȹ+#x<]�Y��H޻� �O-�,��J����{ٳO^�|��R������Q�Ӳ�[�Xdѵ���:����N����C�U���#en�VN@h���F�Z�Of|^Y��XC*�P�P��z%=�MT��2��fkJ
�P��#:`3	8��p�V��P>��Υ��vV��u]�5c�P���[�3�j�Q�t�@dFӸb�P���^x��U���tVk�A�]8ɛ+;�`�Q��=X>���Y��\�x���(��D
�{lj���j*�z\`�����S�Ȇ�7>��8��3���k�����Cb�yk9C���
��H����ܸ�����nh[ٯ}��S���41u����k+u!�u[g�t��[�锡�fwL-:�g��.#y�c�w�Zi�CEƼ5����FŃ�V޻������y�(\��Ü~h�'7��\	aٴ�2��ɍ�5�19����h
F��YHA�QGr3$)���j�2���J�*.y/&c��U��)��3�rzk�W����#N����ܪw��YC"j�;�� f� �V�����p��J���9 ,}U�Z�K��U��_v��=�ea5�^��x�1��+���/�[�a7�e�
�wH�v_ʙ�@a��M�u��m?��4��X!WLʷ���7x�3��[�+���E ���t�pd��ޘ���0Ӡ��{���lt�r�ٙ�C� �fv}s�oma8序Z8o�ӗ[��1`�AB��1W�}K*V�b�H�.��
��'2H;��*�ޝ�̨���(��W��ȈG�R��<�ܨ��XffKx� ���գ7�u$��=�7�.�,���n_ͮ�23t��Vշ�A��6:�=��>��#���t�.��Ҍ�/��yVPo /���ޖ���oVͽ�w�\���c�v��'��_;�":���4�DlD]��]�e!G;�c��uh_u=Ȃ�"]F�|� /Sv���])DPx���q^��DK}�%�yV�
��]Y�.�������gbh���Xp��#��ʃ�9GT�i��b�p���[�{ԣn���z��ci>M�&��4�j�����P�mj�3�uӶ�V2c�kz��bL�!�ef2�bIիm�K�u�v$��f��E�ؕ���l��F<C�@�p9�/�����\/��}�"NV�:�BX�j��h�����S�{[SG����S���kB5�u��n�<���o&�$ʖ�N�F���Ev�
�>�줯v�BL9���@�Rj�ŽV���n���e	��)(�G~Uq\���u�o��y�kOn�P�.KYq8!Һ�<�5�nwۙ��U�9t��5L$��
�U>ͥ��m�JK���=yE� 0L�h�(i�7fem'�E�A����T@B'�\�ͽͨ`�em�j���ry؏kY�k��˥�0#�lR�!!*�WTO.�@T([�C��Hs��ݝg8fd�39���Y�&��N��ֆ�S�r�� �(P��.J�mm�9�VHܦn ����>�ӥ�:{�t�*]wE9i�q�Rc^䰩���ݗ�	f��A�,R�GL{�%Bf�wTB�v[$��A�Y+��K�I����E�d�Jطa$y�w8
ƩV��!��fX��AI�1�Nb���H5��^U�5Zr�fĊ��KlȘņ�.jMX �	�1\�z8������|���
\��ąv�O��t���#{��os�X˒��	ϖ=� w�7�2n\J��5���;��5�WX;�6e�ה�V�Vm��LO�@����k&M���p�޾eX�e��կ���H,bf;&itp��e�����S��@�m�I���˝(S|/^�&},����3o�ýND����{�Q��6��ٵ�L6۔MnjF�����i�rŴ�.�;�݉ʺ�����#�
���f��*�R�w/��5 }�;Uq�溵d:7��p�+��5r[��6l�1,c�׶��T�6A}W�B�>h܋���r��1��!{�2Q�-�Xc'_L���ڙ������+��1��GW!�i̮\�������G�����>���n�33&���c��!i#	J�DiC)��H���9]Hň$Zf�ݹ;�RP�.t.\�H��! �v�)
Q�*�*	1$���a ���J�a�4L�(���24�d$DȒ�݈b�vb��u��4lBR&)$	��#067wĀ#l�fA���0�st�PB�
6(�7.\ES(�e0���D�D��ɘ�,$�D�I�� S A#�1$���Jaݝ\N�iB�s�d��FA#HI$���&X������u�����������5�`f[3��&�A�Y��LP뚵�����ۣ���N����;{���}�V
���G���|��>/kA{߾y�[��x��>�^��G+��_�������=׮�7�{U˕��
�k��}�_�W�����_�C-ʾ._�=��}[��|m"!�߁�o�����6���!�"�/�;rߊ��m�o��}j�ޛs{��߭}z~-�����z^-����G����zW����W?�]�_W�_��^-��W��_�+��������0�� r�3}![Ý�'����Oί���/j7�ռm�{����x�-�����\���p���������s^��Z���j�\����ڼW���W~k��[�zQ_v��Ƹj>�DO���F�ʏt�l����^��W�_��_����j������}^/kA�z������sW����׿ޫ��_�Mx�}�W����>�����~�m�}���7�r�ޯ��+����m���|p}����� �b뤭�Xo2�g�Q����~~}����6�w{\�[<��|��>5����wm⾭����u�h����������zZ?|��֤����o�_<���Q���.��꽪��_������"$DADgN�ޑU��p���S��ڿE~�����j��_�����߫r����WŹ��6�]���_�w��5�}W?~����}�W�����oMx���o�|��徼������@>�E��J�B�K��u��p^��z�zZ9W�~��}b�{k�~��z�x��|o��/~����[��7�zW��W�G�����F���x�w�W��o�r��^�v*����w���ǵDW߅Q>�_A�@�~�B����.��i��u���#�@DH�>�8��}�(�������o��ow��1^���-���_|�j���_�����h�V�x���/��h7�ί��o�r��ީ}"8P��6"!�#����Pp&�ϤW����izĈ�DD!D{����~�n[��߾ok}W=/�����+�o~�^�߿}���7�nk�{^/<_�_}^��s�o�������+�n*��4Պ�����Xj����h�>��i�E�짞����
����}���5���G+����⽪�ͽn����~7�x�����ւ����|���_U��{W}��^��6��}��{W�����y�z����ջ��xۖ��ok�W���Fd~�_��l�&Ѷ]#0!'"�;N7Ϫ�V���7/Afj.���bL��MW.[���s�Jf�����m��R�[�瀽��o_2�XA���[&_ y��C���-3Wئ|�S�ƴ���ރ^��7 f�&)��J�I����k��R�w[�����5x��}�:����=-��_[z\�����r��������~-��Y6�������A�_DH��>��{�QF� ��S���D��-Ϩ�>�" ���>�菺@{�~���f��<����|��ks�x��m���������[�kſ?�[�~w�_���~_�W���]P��1}=���>��}��~��8}������|{���py͏x�k���}��5�x�}����r���r���-�����z_��{U���7�߯7���*��~W�k�zWŹ���^����ֿ�����[�^�|��^6���mϯ���E����$G�"ȭMj��1O��]m�#�h��Cy��}DX��}��޾��h���}�/M�>/����i-�|_��-���u�|W�\�^��k����m�_��zZ5��o�ُ��� �[��}�r∩��u�vM?�}��Bg�"DG��_�}�������������^���o̺��G�_R^�*�>#���b������6��|x?=v��m����h�*�E!���(}}bv|�Ƽ=}�׻D5�g��#��>�	���E}�}��}o�}_U�o��o�r��|[��������{�����o�_7��^���k�\���~���k�>v��v-⿕�x�^�x�6�����������%C���\���~���>��|H�����|o���j����+��_��^֍�_��^_����Ư���-�\�|b"A}�$D0��m}""D�׎��1B>�A>��#�G�|�S��*_y׺�"й��D`��Db�Y�/LD��E^��^���7�n~W�����~�o��|W>�������j����|�����ν-��z��w�����_�z�* ��������""�{�Q�������l�ǽOn��*�SHUQEk?|B~��k���7/KF�W��o_�o������5�oKs{��|^��n/��wkү����w�>��[����/��^>���Ĺ���|G�����E�HT�;�{b�����P. �}�D|Ǿ��=�G���Z�/K�h���{�\����/�/�׿?�Ѿ+��o�~W�^-�����^��_��k�ƹG����{U�rߪ�{���ͽ*����
��_�N|�\��;�sQ�>�ag?ܚ1+~��%�\g�2X�l������6��R�5�o��+݅X�ܒ�j�D�6w��
���X��4���OS��7k����E��f�]5gL���]��Wn��C�����[�ߟ�U�k�ݷ��^��~�����皽76����}]���|��b��*���YQ�0}TEW��hB����/kF���{_�k}^�����o�� ��DGu!Ͷ�wbV�l+���}�{W���|��~��������o�żT����nn�n���zW��ϋ��?}k��_�rߗދ�m�s~5���/j��_<~���֢�U������E�D�]ߞo��M�ث��ג�����>�t��=�#��(��B8DGI_�����{Z>����������^*��>y���zo�_;��z^*�\+����{^+�^*����/]��^
4G�Ǧ" �"�����/ʯ{h鬑~y�+;�����b<�Eq#��[޿;�~��}��������wU�������r濭�����{߿�=>����KG?o���+����}�z�ʱ_PAUk��HU`�+�ͽ�ן��#G�Tmr�yl��}#�"4B>�?6��nQ�_��]�����^�ν/o��*���_�_Z�=����{|W���~��~k��ڽ-��������W76篟�oJ�]�����|��-�W�}޵�����{׸�VS�{25���w�9z��?�_�}����_�z_W�D��Ź����>��~.[�������U�����=�⯋��~u�M����~W�o��nn���-�\��s�#z��ﱟ�}􏅥��G:��^�r����no��|��{U�r�6��~y�j-��{�߿���{5r�߷��V�񷿝zm���1�w�����뽭�������֏����+��+�^�=y>��#�>������>����ޱ���_������w�ּ_�������}k����}������-����W�������|��^/cQo����꽷6�}�W�<���ss_��W7�܂#b,�!`� >�������y]o���ϻ�����zZNj��|W��}ߟ�o�������_��o���[����Ͼ�"]߭��x��:(Qn�ZD��囝<�U��Q9��8���*�8$b���~i�F9Ҿ�?`��C���N�oT,\��yB��±{��s��##�sxD����쌮,N�f�75v�&�î�ǂm�o$�O�/�k��:����Փ/�*s����n@*g1`!=�N��.�����*P)T�4��L�/�v�B����� p;-��
�`=SG2[H��j���y6���d�=d#R��:����\(_����03��^�ʱ�`}�w�*�~�v=R����6�䈂���g����@��t�j����!�ݩ�U.�F��H���`d�(�T+�S��#�R��7گ�aR}�0�^tk�b����=da�U�s�@�+�v��S�����.��*І�3�W�C���f���tc�*K
}[s}&��&,O�9��sf��� �ϥ�� �rz���-�p�1Olp�܇o-�W��ۯv�aI��Ϙ*�T<i�_z��i�h�j�hЂ���m�w����:Tls��n''F����"�΃5����^Y�:���k=��<�z� ���SeN�q��7~����'b� �@dt� W������ڨw����N����BϜ��5�L�U�-�>^B�O�?�r�k�{ �<~ @�w�ʗ�`���L9ܲ0ŋӵ�������C�b9eN�.pa�袂X��E/�U�W��K7Q7�(5��,=ܹ]gg5��.��ĹLCx?h��z:�/�/��-�x6S.�vs+�!uD�sU4�Ycs��7������f�xݩZg}���ǜB�.��v�Wv
�餃���N�����2�u��w�u�H�vMqU��CPʠ9A�|���Pܡ�]���7b.���M�.���{�)U�U����>S����,;)��iO&4TB5�19���=�)ށZ[t�S��ʮuBh*����S�EE����1�ު�W�e3�!�.We�R�|��q��y�Np�~�r�0Xt��n�(�0;n��&��
����u��'�w�hN�⺳�1~f��3q�s��jwH	�{��Nx� �י2�����F���쿛B��ꜫG���]����p���a������f�M�H��PB�:E��lWН9�Y���T@��-��2,�]gIH�9N�	���c3���������8�f��t�f�.����q��ą[�|xC�W���E��鯎o�Nᩞb{���!��~����<�����z�;�s��֪q܉z�OjQ���n�|�95�!¹"~������*�N�b៛�����˳�c��a�OӜt�wu<$.�T&ۈ���Q��cd�Q������B�Hs�N�0A�1؉�4声��mњ��r��V�}�[��4���22�Ө�l-d�T^μ;z�����E��@��4
E���<*���Ӯ�f��@r�IO�
[G5z����oF��gd�.���Ş�o5��y�6�G(�J4��U�����q_]q�W���{���EU
ﯼ� �z���m�>�2���{�倪�A��:l0W�C�j�=E��b!�y�;*���\�:�R<d��4���^aU6�⁳}ಭ�nؕ�n:���@O}��@�xb��au1<X�21�8'Lira�[R2�2��ԙJ���WN�çNK�<=TīS�v�`�&FD�b4[y�q��S:po��ph��Z�R���,[l�Zd'5��&u���a���o:P_l}�^g(A�_�{>4�� �<nw�Y��6ޮ�T����gԶ݃�M�[��1�|r�����������:[9��\P{ܪ�5u	9��$�wLݸ�Ki��|>�:y}n���������0���>�������mC����=p��ź:���j��~�G&U��a�K�Wd_:w0UO.G	B8[V���艪E��K�ds�=w�cs�!��f\!���w�[���'풑��tO�[�Le��NUm��ʛ��H��'I� G#x�pU�V�w1!X .+�`r;��{qpz����RmRq
x�l�`r�ՔUǋ)��i�6�M���T��7��]l���y�R�sP����&�c$3���}7�zC��dפ�w�e�Uq�Q���M�X����{���L�Q�eJ�^s�����A�N�ݩ׍&��5���DD}T�y˹�b<nsC��_����gK�m���ٛ±�4�ۢ��fL�jˈŷ�����QVT8�ԡ7T����G�٨+�c��v�@+�j���Hwd;2f�0j�y����2@�t%#q��M�bF�)cw���!�����M�P��Tb�|���g�r�0q����_�B�m��U�'�T��g�yd�c-!�5WXi٧��_C����r1B��@>ª�3�d	�rģO�'[���&����`��y��d[]�V��6-R@��Ŭ��Ėxc B�V��M�N&��e��d���	01� ����)+-NB�7��35� 캇gMj g�:�o�pECyFU�@��-&qa�˥ޕE\���ʄ���lV��Xvg��g��<�n"c���
_)|���ȍS-:��/dM�xÅ�B�r��0�Q�<2���W��d�| _tP{Ɖ�՛��yǮW4� 6|�=qT�9���^UcbUк��~@W:ɐ�l��<�e��w���:J��E.����'gE�ad>�-�3�Iw{��9-�5�ޭ��0���:���y�ψ�l�>SY�e��u�v���%�ݪ��w�uh�Ak��Ld�Wh��˔g!68��[������3�$(zꐋdr���}�Fb�oRg*�D�>��Un|��ŕ��|g���4����l��k]B�$r3��%u��l��Q�T�N���k.����c��.M��2+_���r�;�0�V�:����z�J����#!�:�ahS�W�~ct�X��N�m��5PA��VpMn>����^�\����Ѝy�
�����WK�v���t�7����a>�92/*��yԜ�ޔ���ʖ���^RHF���Ƽծ1|�!L><���+�v��
��ع=�l���T��.F��g���m�a����'��Ϩs^#�È��W
��NS��ul��yJS��B��>�>�>6��j�v'���5�v�����bV\�&z�Py1b���յh���(X�� ��r�eÚ����!���c�s�n�o�9X�KG8�9ŉ�����ug�>F )n Wz?-N�G�X*�,)좕u:μ���$꘳C�|�G9��Y�L��(:�P��3�1I8��mUhy�v�;���"E0��ռ���ʱ������;�ͻ�)I��Az��z�-{w���X��!���v��u޴�ʈk���ZtX$��H����0z��7t��ٕ6uٶF�s�rm��Xjw�]j��YzvIi�gY����9^�{���M!m���`z">���OZ��X�tDr}=)���C2 ����Q�A���@fӸc~�ڈK���{�GC�Nłﺧ]�%F��������� p}-m{Y�YA1�j�V]U���pS�g��ږ_���sϦ��5�s'1 �T�r��P��*��^�^B�_1u-V��� �^��<���ڽZ� ��,+�b.����_�~�����3�M�EV�|#l�9�v�J��hۛᆃ�'�=s[%�93`�2�]֦s�:�t�7(h���O��E���B��x�2����f� >��'O�e�F��!+ói��;�S+��2�S�,���yo>V��Z���h�۞\�5:Ȳ��ѓ1��j�����C=����2��6�-,6�oy�1ϐ�b�����@vkpk�������B)�[_q����5z��%V0��<�P��C������>��6�܀��*��*�v�7��
�p�r	b�w�}�n�!a�*\q�����(:S"�N��,�l�b�`�{�e�zm��ѻ~d8ׅͪC��ά�%�S�(xfKQ�����Χl�v8l����y���Hn�W�*�S޷�gH���]�����9����p2�'�^uin2C��q�O���/��\4�D��()��fmB��fts[b��B1��T9k#[�}�}]�Ov�Z�ٺ5��_!=}�&a�PZ���4Cʙ:�D\B����0��+,GF��{��8��>}S�r��z ����W����F�rz^Pi�ȫuP@ge�]�R,�Ǩ�t�����F\�0�?V9zw ���¯��x�7�~|J=��;�7��͝~�������@uœZ.Rn�r�Վqxb,p�����������p0Sgw23��:�T5������I@o�+Yʯ5�:�K��ٮ�0��:��YL�y7'�D���tY�UC�'Y"p��}Z�O��C��:뇧7v���mhW���6H۟-��*Xp�����P������bx�vdg��+�I�\��mV�Z�\����s�^r]:�L���r�& S6ȴ���pfTS���df�+[����)"�lgs*T�`�G����K5T�C:�^��{|�F(v�u���5�M�j.Ը��ےnͨ}Zj�o���n��j����_2�������?=R��DA:c Q�@ЮJ�'WvA�f�vؼ�ݽ���8u'.�P;g2͙����T�&��Qn���W*w1:��
��Y���;ln�+��'5�np��i�NQ鱕xkEDOsf���v��0��K��{è��hj�r7c%��X)S�9��Z5�oF�ӕMޝ`|	�dw��x�ͻk��]��wWmJ���ro9p���k]�eKU��$f�[�m�p���r���Jx��bZ��Ӣ��:�1D�h�g[Jwq���{�O�]Aݵ|� "1�묾)]��xoE�bl������n�=���WK�O����`��o+U��n�j��n�����1XZȢp.qI�|�8;t��k����9X��幢���(f��@x��g,�FP4'?��zk����h-8��Skp܅�8��o�����CǷ.f�n�F���a�x�FtWsξ����U�ȺM�/���F��+:��v�<T��Ӽb-R���[{�|�wwB_&�f	ۏ��0�54�k�m,B�r��)�s^!0V-h+ *5�f5ج���3�|F�_g'�+s`]]����:�wܺ��\���A�t8Fk��F��
�Qs�˙��dg�*��p�IU�f�+u OM@iԾ�Ҥ�b3V]g|h�֨١��d�zE5�3>[�/�"��C2�̑M�Q�k�P�|�i͈(>�b�>1t�9f�����K,��+o�\��C�CN�O���ye�uϭu��ó2jWS��.���y�Q;�e-�����13cBw���|�ݥ�`[+��g:�m��C-s�*f
�0�j:v�+��0�C�3��b�Lٗ�T�����֪�Y�9M�s��7U�������ZoK]C4���ѐ�ǟ7��FRU���<�Gm9��_Y��W��ob��r7}�R�y ��X�U�n��]:zl�?��έ�w��	QϮ��c$)t=�R��t���>��2�]_	�����Wס�\G|%`׀���-�[(����Tp�uK1T7������,��;\):$�t��W@D�jM�,w+�%���ՒSM�3u����C�e
�F�Gn�[#L�ӖN[�9+Ue&&����C�,���pV�WgK"iM�R���4s@t�.�(��݁��k#N�'�_Bl5v���^�_P��u����Ἤ���[�5H3q�o�v�{hÖ�o�N�[�A�w��J�Y1U��)-{uq4��6\�1�6�e8�Bzٸ�u�A鵴Y����Z�\��ޜ�H��v�b�6sVRSZş+��g3��FcxiVs
\�*���8h�M��ef�[
���J�{�]H��t�ut�]�&e*fP�a4��2jj�n���b��yG.�v�VȤ�gME��[ZC���,4����]�t��V9E��@j�|7����V"���qB�V�M+��٨r�."'N`�U^�.��ŵ�.s#xᵝq:F2v��i��\�;.IqA�(
��Sws(C"�'.&�4�0�n�30"3�� ��d�QHc���,Q$&%�r���(�$�+���`�f�$w\�3AM��D�I�Lll�4�Ja0�h��w"a,��	� ��d�C2R��))�1w\M���;�%"��Đ�';9\��$Fw]�»��10ɛ#%),�l�h��`�w)9є"`�D �&2�ݻHDL6R���.\(L�f��Q�Cdwve�¦wt��$�"�75��M�Q
DA�v�Q�e��D��R� $�t�1!o�
 T> �
���:b쎡�ӝ�)�L�/C<�b�*Y����Gr�2��c���Y���A8Z�h�3E�oݽ0 ���g?����ӱ��'j���kf2����0�!\zR`u5�<,��.�}g�h�}.ٶ�'7�4�VJ6�Xu
��h�&U���)K�Wd��~]�S�ȌuD�D[�
[��F����tj��j�]�����17=EpH��|�5*�����e��_s��.iB�`=�|Ug�P��������G~N@���멋/*$+���Ɋr��+��߹w.'(Z;�i
G�xԁs7y/�_uB�:_�p�9U��"1�:�������㒹A�ɥ'�<pG���>U�bQ�j
��R�0��ʜ��1t(�8�e��ԟT���dBxj����|�KD0X�ߢfɉ�[Q"��/N��Q�!�P�uk#i6�/����ZGt���LX_?O�}��J���[tܕ�x🟍�vxC�`(̼�N�Y�vp��݊�p9���-ݍ���a�*Q��%��3A��ɅS0h�f�.�*M �r�BZ��5#���fl��Vkg�|< ���x�Tٸ��C.}^O�"�w���q��bT�J��8��vyU�8� �o���v�������i�;��Z�r���·��^r�3ݞB���4��Lՙ����e(�f�g4�ϟ-���D\���o���WJ�s��B�4�RqPQkp�]d]�kGlu�!����$�磌���7+ӽ�>����Pw���zy�&�LA�u�;*�5
5�<"�m��!�#�v����ޚ��b��A�.s��\f�΢.pV�#\�@l*����x�.��kkV��n	�\���޲�S�j�l��y�eR�^�U�*���~4�_ /�4=����28�n����EL��0�����{hu�3���+�u���]��5�%~2����Q\^\�m	՗&Ċs��q\�k�׎�f��G�f���qU>ѽ��G�O�4�ι�-C������N�::M�E��(EF�vS)���cE�x�����Z@+�����O^-���W�q6�y{,/TD�Qo�b
)���eB��iȍ?1�o�別4��2�������4�z���`T����H�k�����TAc�i<l���R⩏��Y4̯]Sȉ�3w��X���=G��K�t���Ha;㰎5��Ѫ"��U���ca���}t��:��n���n@�2�FD'.L+�`���x-�"�J�`��"�P�Yq�ȔS�
Ƅl�����"�Y��(	i]`����RQC�k�]t��`�8��wX�`���c�Y�T �+��\/F�2��/ :����e��K�\w�6��6�F��y�öᜋN���xu�❜�.�]�*�9M~���>�b�[�j\u(���L}��J`
���"�̣\�6rH�LU�����wt�im��}���0R�!�$%�Kj�ϊ�bB�ݰ;�z0!B�nO'��z��,��Z��f��u]*% ��y�5
hC�ee�uVsa�����`S� k�q9^�Ʌ��_x�~����p�nh�	�*����
Z��ϳ�:�SƟw��6�V�����/�efy���
����.\����3 �aVp1�=V��Ҽ&s�+�P�~ҧ�ל�/�{�Y鄥�/w&1��(k7��?h�璼%Y�<%
��𣕋������\&��I	���@i=�tƅOr����Yv7�V��^B�B����k�{�\���җ��� ��� ���([.��_5u<3��,�ӹ.�11h�Ol�7������<��$���������@�x�Tn���9����0V<��-�!��y�Ϩ�KZ���9 ���W|��L���>S�e`���')��0W�ƴ�#���9J>!H�b�X�k����?�'��ڿ!w,���9��HZ�c��R�]6�]�>�Fv���C6�9W��om��Ed�f��{�ZS�W�um���~��sy���Xu-Q��,������X��ƫ+}�M���	�l�unW1��9gMo�!DD����������<�s4�<���@S%ܡbf����"�._0�����+�͋�9�g����o;%`������e�z�(~5lC�اds����L �O55�l��: �\�ɧ��/��p�ˤ�p�Oq�����`u�_ta�#Eʁ�Ё����G��u�ࢸ�纲�oTU8�p��$q���[ X�oZ�~R�hƐ���Q�"󽚽a��Z�ӆ�%��I����N*{�\��B�U��tn���ԈD�#9�eh-��{�"&���I�݌�͏�NN���@Vy����C!L�5&ޠ5�y\c:s���e�S��zGs�p�D{]�v�G�O鈅T8m��)zw>�	)t�?-= ����&s��n��º�;�D �؃4c�U��΢��_Å�����D�=.���u9nwC�b�l��ϒ��c��']��U��s6���M���Z�5�k�?�c����쨝z���Z\}+��1!���O�2q��56k�q'�9��l5�Y��!�N��6����ɡ�5�o��{@�n�Ҿ�O��<�Ano��=�zQ/�h�qXn.�іf4Ĝmm�\+���fғ�駎yHV��:���R���}e���j�sYQѾ�syi,cI�.j�����uN3��Z"x�t���#�;ִa��������i��G��=*A�'�� $J,W�UC�S�ڝ�B�Ѣ�\�1_t�iL^T�B{�yB��A5]p�2]l舶v4�\�	�L�k�}u/Н�uC�S�9�jizN�*���M�Q�bƅ���V0O��'g��K<�VrkޗC:Pz�|�͈/�W�P�{�%�����*����|�8��j�xnU�c����i{O^�+;W�~��[���k��n����:��>7�	���Onx�bW�EL�k<xO�*��\7ۧ��d��܂�n�-V��҃.X���WL�5���M�1��
RQ�Y��@��M���Y�[9Ʊ�<;u�:=َ��s���9։WԼ7/���}^qׄ;�)�.PƁ��:��텰��Qq9��f����VF�$j/����t�ϣ\���qZ.2�!e�D�lL�v���6E<�M�֕�C�X��3[�u�	��9���|j/xT+�:������F^����O^mB�ѭ�Q���ui<'��W�v]SvJ����l�p�X��1���!�n��TcLǪ�@]W���l\>;V���yN61�6.<s3uS���+-S�w�i����1��
�}c�W�؊��m]�v�cLGl�|O\}��KM��9�z4�hʍvk��������>1p�;���Z��s��Ӝ��]��	ǆ���K(�J��^�>���>����iܝ"�>����w��Ӓ�P��`�W�%	�� e�\/��Ɨ�����4�RPܨS���jKnCsrb��^���t~R��[>շM�]��	�?+EnגTz�c�;�������M{^
��CQ���2-��l�̱(����EM`z]����ح�F��ky8���k��l�g��-��f�`��a�s4z!w1�k�[u�;��k,�н=�왮����RZ��=x~c����v]C�Κ�@ĝJ7d���EՑs+r4�Q�(��ҐL`��p�,~�b�]��!�R��
�����n`I��ނ˖=���2Ӌ5��>��^#^��b��gʸHU�~TŢ���_^EMV|��N�]�VIX q�cQ���[Y|;#�ܣ��i>n��̮#nh�Ә�=�Y'F�����D�S!���n֜�0�_����w�#>�c��Z�����e'�Fo��e�u�=��8�����:V��4�z�Re���)��jwLh�U}z3䶤G\}�{���_d�=��o3$���Zi�f��K���4�?�p6�#�s�s�5fZ	S	���U71.��zx}@Xvh薊&�x��-��XA{������,h�)�U�u�ul
�Vw[��z������.��IΕ7͓9��j�����/*(��(��12��'��}�}C}�����N]?���qE�$��VT+�2�Ӌ��9�����Ε�>�нzxi�p�=�Њ�qd��*�s1aC�����#�*\v�)�ʙ2���g5C��ӂ�|=3���X��YB:K|v��Wd��{_$X̹�;B�����5rn
(8M���~=86̣)�:1��A��w]6��H��3�'������WG'禯&��GKʱZ��%u1�vt��@W� �e��rZ���{=X&+Zb���<�����;œ3.�:����"K_Ǒ�������*І�����>�G;���G+��k#Ӟ"����5� W/�}3��tG>��PT@�5��Ɋ�M��;�Sy����1l�c�:.]�������P�3Q�V�_����N*Qg�t���ԥe��.��i,
�9�)7%�rX�etE�#Y�f����.cY[��x�s�4E���ONͷ46����pY�?p�;P���(\x��롆������q���[��Z��>�P'��۰��(�G�N	��5��2��s��2�f���[-���v!�Ԟ���ѳ[&]uf����!:���%P0��юrY�doRq����#-����KUC��k.�c+9�i���)~�����-q�z�K�j@�d
����9���7�]�5Y�cd<,���oHWQ�� 쉍���9٬��,`F� #Q�ˬ�����
�M}Q�������W�j�I��gXo{O���c�����Y�f��F��k�2:�Br��V�^<0?��֕�+���&13�I��q����$Xpzp`;�V�[�:~�0�M�i����2���&6�V0�L�7��9��7E+P���K��J|�i轧��Z=�g?�����&�C��E屼*�r���q�j��}sF�b���)P�)��W ��絏�zǔ����~����Fk^\�
�w��/�\n���������@{2E��a�[�r��T�e ��<+��EK�����B�]Ÿ(pQ�@�P)�Q�t��d@x8Vڿ�<��?~�֔��V�7�Ä�w3����P�T6m�V��!�Dû�����:�~����nܻ�m��<x?�6���˝G2|wN���ϫ�a �2三y@s�;���r����/O�D�Ǭ�F`���	��3*m�n"&�b�Ř���<��
�ݔZ%g M.�,�)�{v�L�ڠ&i�� ��s��'_+��>�*9���А���n��b��Jb�P��p�;n]&��t��Y߾�꯾��eb-��r��=�P �S w����J��T8m��_/a����s���J������݁;��Ҥޫ��>�=U��@�co�� NaV��v��8�18X�x|/k���KvtC�W^Wwζ���Ӡ�_�TŇ
� �vu�\������ٮ�^�u;�<8�9 �j��.
��0�����"�C'�̈`:��}�%�q�Ny�F)N�e�^	㖐ij�L�Y%f?�'*3^����Jq��w��d�b��9���y}m�i����=���P�)u/mS�Y�ά�v�;\�n������<ʕ�,�I�w���:*�;W�iں�o�y>���ss
��iP/�KEۈ�o��䯸�%p���D.7�Ҙ�u�]���*f�3��$�i(Ks[��u	��YI\����u���V42ꔩ��
}Ў��ͧ�w�5��ϵ;{JkyC��׽K�mu�Ru�U�5���_&T*�7U`A��T�;��D�rT��V�iU�a[j��o�{=j�^���{^TY�g�κ�M�xVdt��@+'DM���ΧC�5{MuX��{��1}����u{s�1L��tUL�z��en��
-+9��_	O���y�ޭ�E�ͅ�ﾏ���=�Ojp�Q�!rUe���گ������9�����	W�Xo���1p�e��[��=+"y��)D�mM�.���U�J��r�q��:K	�}����)r�O{��2{�>WS��<��.wc���Vu�o��@��_>���-���X�ҥw��c���<�U�H�{>��:�����y��8�Ȳ��Y����V�M)f8���6g5���7Ep��L'ӨL���s���8{�tu7p��Te�����P�Ig��W��׻�������T��;Y���>����p���;r�K�mMU�ؖ%��v�I�IھGfm^#8�����TgHu���n�5t�	�κ�vT����3+�7�:��1�E��b�3��Yӊ.3���Zj\A-��:#���Vw��[W�W��\fj������PzTw�fSm4oTn�C�A�٤q�ai�=!�c�j���6�+�N�@Q�9���:�S\�f�d�m��E�]�H��6�xt5��n���d�x�� H������ݵ8�u@�ǝ߃�-i̮I߅*�M�Yz��\�5V\�RQ+s) �
�̎���$9�;���8�1v0wLݼ�"�#9S���f��z��b�{��nR��R�Sn����v;����C����m]���a�dG����Q�kǅ�'��F/vѻ:�DNL�82�(�����u��v�8! ��-��鐒�3�Y�k]�A�lǷx����)y3�q��X&eQ��3%��۫�����	&��]�hʎ�Q���%_ʇ���s��n��3Յ��iar���e�^��x�o��md�{�2�<������o&GU}lW�FZ���ze�ꗗ���"��b�f��j��ӣ&�p�9�[<{� qV���2�r�DhPB�[V����NN�x����t�m�8<6��G�,��a�D� �V�R��ڴ�2�	B�c�P��l�m�
��4����P��d��$ثH��t�Z�i����1��;(f$}Z6���y��ĜVVӰ�[��sTTl.�ہ�*Z�s�V������y����=�l��t�֮�,�u32�&Sk�{g7H���5�ef��b0��K�0��2��p�`��@ӭ�"�
��os�cUԎ��9v��kOZ�3��q�4��H.�.�g��� -�qL�Lr�r>oM.���r+�/4 �6��v"xޭ]�ۮ#�c�e����;2=P�P�}��O�oi呆D����ꬾ�x�VbX�L��U�*��
)r��2�l\�]�;���������8���s����	��zfX�Jr���\�4���$�B�H����y��]���ޭ�w�5����"�ut1��j�>�ll�f:_\�ʕ�
*I���Yp\މ	�٣���n6���+s3�졧]]�+����̈́^%�Sv����1[����[)�{Ϻ���i��X���a壦�7�%S�G��T��C-�+-@�\!Uʳ��V��m ��Ҏ�5}Ӯ�W�o�1*��bӖ���S���+kz�ۭ�NC�=�0�S^6�O,j�ޣ�M"��qن�5\.�Pa�Τ��Jءc$��=�
u�(J�th|z0�=�v�)eӷ�^�;Sd[[�03[����{�1w��Re��Y�[���ٝ��E:�L\��̓.�٬�*`Л/+Gm� �ǝ�k�9��ZRj�MR�֟�{:����ޮZ�RJmqz>���¶����q����w�س��U�yơ5�*�KV�)c�k��N�R���˴2b����m`�³z"�� �" � �&$�"B�ș���0�ɡ�DI�1 ������C A3% �2H���P�3�2@QJTiI$C�H��$4c)�d�f,�(��f�bA�1$���l�U�b"C#�R5i,Q(`0BPY�QJR9ؐ�PX��RM**LS'w2PBM)��"�,��Ɗ#��"�F3&S)�Ph�P��&B�����LP���!Id�$���ɤ� J���I,�-˰�i(2Q3)�]�b�ot&��X�g�������*bl�U�K��MKU0��F�m�%a璲hkg�U+G�����,^�Qu�"e�_�>�������H��sJ?CKz�	�i3ܭ�C�T9�(���T��{�j��`��䶔v�ˍ�J���5�WfƼ=K0-�vī��QJ��ْ�fOW$}�n}ʻ��S��S���t�����!�V]m^'�s��p{���:�󨲹�iJ���ֿ��SZ�Y[s�RTUf�֭���	��w�m�����>Ue'q�օ׸���6�d=6GT�=XL�soy�;�%�P��w��ܚ�)D�]�N.觎�|�ݴo�fz���Nx;�л��0nS��i�u:����P3�mɩ�Ϯ:�]�Y�yeq�+ �H���})sy�[�qN����*��U���nM�AZ���^�0�]�w�_);�9ޫS1���B/4,��uf����U����uv�ܞ;��j+�S��Z��{�҄���1�4�V���*㩻�WN~u@��}7q^^*f�~;:��RX�U����֜�o�iZ3q�bU��R��.L�-��ws��OSK����;nQ�J���Mv��-��+�}��8�bK�W7�k	��x6��c�T�x't!�9|��u+�T/�aܮ��������6w���'�}��}�D�H�nY���[y��+��ǐ��B�f\Bp��bۋ�.8썽���/��0g���;���5���*�����I�ksy¬�}���Jq�q:����Fk1��mQ^z��e.��k���/�WA��ŝp��Qp�=_2���P�;C�\�~:S�+9�:��d�Ů��vw���Gr���{�5�h-�A�T=Eo݌�޻7�ݵ�zr�_oK�q��\f���V��y�m�ѻ͹�<;���J��]�`��&��q{h�6�T�~)��ޝ�^-�V�,9�1�2�Ry3���vL���s�v�5�dY�_E���T����i����<M۱g�c��c�}&��T��ί��=��'K6�?o:���:u[^i������.ꙧ��Ỏ{_)�Q�Vl&BP�f�ĥ���8ݲ�PUSFY�����n��&H�p5*?���O9R�KʣߖŽ�N��O�%k������7�,VzV��,��!������LېۚF�fgqS��z��;� s�o#ӊ�Z�3�#Nh�9�����vuLH)�b� ω޼@MFVd�ynQ✛C�U}��Wվ�2���˜��}�$���}�������K��{_I���H���Lͥ����С�vj���[��R���Ծ�NQ��ʸ̪�I��J󕔆H��nNk���1:�[�Zݎy�c�U,�d��Fp��3= S�B#�+��;j��3��1+^_��e�W:����+l�p�2�t+m3=Yy��o�Wg3�~Zi��{Y�x��lVtY��پ92��:Ŝ��M��ǁ�dsHeP����\y����ٗ��f�4��>c)r�w���)P>f�_l��.ֱ�*��H�o�'����Wy�ꨈ-��ͼ˵�t���O[�:��&��nc�z��O�T�Q�Y����h٪�����\\��Y$ծ�oӨZjz%�V-������)M���N5�繓P�;��V�h���9�8��U��P���!F}�u7Բ�u
�����o�N�1m���&s�!h�ˢ���}gr� 2�{Ϗ�d��)mO�7;��[���nH���[��+��{+�,�miǜ���(���ݎ��:�r�X�R��}+�^X��]�\5f9��&��<�y�����7t�_}U_Uf�C��y�f�~���y��g*�1�b�U^f��{�,��;2��J������]MvV<:��]�y���s}J�,�/��mj�auq��q{����0*_�_e�MnC����/���\b��H��Pbu��c�0�:���ݙ6���2����wN�T�Lիo{�&Н\�V]��Q����v{��nuz�Y�u���ڍ]݊m�Z̷�:�T���;kg,}.f�1�ޅ�jJq?W&��L�c�����u.������zݻ�q���;��큫e�[*�5b1vɹ<��t�+�[����}��e=v����?��U����)G���Q��l�2��ٖ�&�)�MR{�D��!O+hc	D5
h��a�-o�ʉ�+rqj�6��}	��.V�Rc.a �䶔'�=+_�)WG�O�Cے�'אV�=e��ZV1�5	v��h�¸�ʨ���f��Q�f�'���3�}������z��Ts��5����$垮X�pF"��}{C�a0�1�N��'���ov̔��P�^�|D=�G�N���w�L����X���X�\'~��˶��P�e�`R³;F9�ۙx`��Y����}�#�o���e��Z��gMk�!_k5P�8k�5`�vs�@j�;L�T���5=U��$���8��Nc��gHt��ڏ��yE`�E>�3V�����������ng}����Ļ��K�S�{~SVU�g8�̔�N5o�{�s��X��ׇܚ0�[\�]��磙������_���5��IQ6ܞU1��)ͱFo<�|�y�d�/�c2Q�K���+�U=���\4"EPz���˕Yqr�ʄTO+nm=U�W�k���r�T���j�o�n&ᕚV4{�-�-
�Z�Y��;ݮv��5��BPg7��	�9�8I[��MA���,��ޔ��������;$Q*��R��u���ҝ��W3�mc�wӴ��Ƕ����aZ,mk�<+2�E��
�d���Y����CP��	B��jo�]4��|�P�������8	SzeK�vLQWV�+H���+i�1w,捪�B+��bH���s�˳��m�h�ِ���� �N�~�c���������)ΤY���|e��9:�5 �%�]���{�.lMH#���Jޚ��B������W�}_}t�o2�5rl��7r�Fz�C���ҭJ�/������|�R�TǇ������ ��/y�˻�o4+�q�N���8�zQ��՜3�vS�N�?nzh^��p;�.S�n���n�;���*�v)c9���SAuWg�]^,i28��q`�Y�̰�~��]%ke�j{�K�<���'� �z�jŕ�n3mnX{�f1c�
�)�f�'���dԳ\i�z�UG8
�a���%r�KOo�����w����r�G�!���*ƨ�hꑧSz�uC)�W��Cތ�c�).Ҽ�����o��-IBszQ�.�d���RR�u�s��v�a�^C�yy��wLm�P��Ine�ot֨?t���::_rye讎|[?QHX���#?A:;S��{�F����Q�}�3T_R����^A��ݱGw}Y�^ui�����n�B]�m�oS���J���اۗ՛�#�y�*�Cڽ@�����B~E��ޔ9�Yq5�ˡȝ��,��a�����-�К�7xR��ݎ����0�@��3��I;:����g?������Ѵet����������۾����=a��"Wx�^ڢ�T�Ǔ~��;�k��S8"�{=�S��a��f�ٮ��	�v���Z�8�,�WR���u7q�q�����Nv�v���N�אy�V�����|�.{3(f�ۭ�+$�o�6�L=oq�5��J���;ic.���b�(�ߜ�%r��Y/���Ԫ�ʚ���ԱG.�P�F8���n:�V!r�P����Y��D(S35���k"k[Sx�kuR��Cl$��W�QNe��9��n�ڧΊț�xE2�]��x�V�[p�b�q�J7;u"�f��3�D�0�`՛`ĭypfXW�^���0=�5e�kr;P/8��p�e|�10��A����2�&�ݸ
�ٔe�X�]F]�l.�
��s�a�}e\:��'��*�O3yIv�G�q@N���]��+(ʠ�o���XB� f'�2��3_r���R��M�30����K�Lt葪�nKߧ6�OfӔ��j� �:��y��o��W�$���_o$�]Ǩ��-$\����z� S��DG�DSd;�7+��|�&����Ể��*�N����+�|Ω�bpe퇼��%-Zo��h;�7=T�:B�Z����;F�Tk��a�7�s^j����S�(�vNG��+�y���	���^���y�<��"k�.�����9�ү���W;gQ�6��j�^�}Ju�>�6�i�ݲ�V�ޞ�y��"�Ӓ�^A�NA�=EAڎ.��Q�Ly>�f�=���}���܈q�wN;]΢t��J����\��������d"�I�7Ret��m��{P�<���t�vlX{�"��g�Y�A莰����]~�1�/���>�j�QS���v|��%V���n���hs[�<R���I��B�5y��>Ue.��Q���=��}^O��h+'�s)w��{��k_ޯ�P����J&�57�.��U	5�����3(*K��p{M]Lv�M�h�5�+&M��}���J��ȱ��뎥�5�ڇ.R���y�O�:ښv��=Ԉ��RZ�.ں2���s��}͸0 &,�����|b�ۅ�
5�2#����Ϙ[6e^v�7՜�C�:V�����.�i5��1^��:õ(�]�HT�/H���O�uݥw�Z�Uy�o$,͖��*'JOᙣ�%.����W�-���k뀻0����w�mt�w7{�NO8����V�D�Rb&:B�k�BkwvS13��x�f�K�-ݸ�r��6��W�'Ц\����B�*$�*���P[q9[����9�Y=!Oݬ�$���Sm
�S�ʛ�}j�s}y�ZX٩�f��7��%�+�+��'�ӧ�0���|�c��Ļ��;k1�u�|�A~�9��?$�P'�X=H{�|Mij�t=[��f�6��{95�p6Í�^��j�}�b�Լh�/e)a^-8�Y�=N+���WПn��b�hI{����(v�2�s���׫�/;��I�}�]�=�~Bo%|�P�W3�]�^Hof(�z���x"Gr��vi	�����͘�udf�jg#X���1��w=/GPB�R�mj�"aow"��sw�b�}R�l�q�usQI.-r�+�J�;���z_kG���c,��AV�t�y��^�x�#��Y�]�.4�b#��[�6H�U}_+o�z����R�8}�f�����k�iec[<��9l�:����:�y	0�(���nj+Z�<���q�*���jv�&�s7����X���͉��3Uf��|��󂴮��5��>Vx����
���s׸72ݘY���(���o����q�ж��û����hJ7��jn1vm154bcBW�z5U��w�;�[r�nU�J3�fĚ�έU���:�.�+�T��9S]Fq�7����P��d�:E9�K���,rY�y\š�1� ��185�v̿�s���n�;���B�C>�(ģ�Qs�'5�v�i5|�wH�c��4/�{�p̰�Xy	wZ�����:��k��յ��m�<�
3��Neȯ8���V�/'U|s��x`yoL|���%�����pUà�%�d�O>�3K//�;��M��*)��S�c�1gƲ�uv,�Ån5!�dn��!�o��ٱY�xH,��G#��3<�H�R�Qu�ʼ�A��43=9�z�q��P�c�ԱGx�����ݢ�Ϸ�X��ٚ-���EbJfg	�]QXIN��e(�d��y5�v���N.��Fݫ�\�)���<��e딭hT+�A�gmu����w�%��
���58�\#�4P��K�����e][��h�G�7r���4�츨Mc�n����l�.�)o�37koz4x����u�8-�ؾ�(ު��S��m�u(��̈���*1#�4z�@�;1�)PjNO:�g5Ġ�C�s>_>�e��`}�.�1f��p�Yz>�	��Z�14�:�Z�ޒ0Q��xV2�nМ�IEn+/�l���tN�T���#pZ�ф>}�Tw���³���5�([U�ZUɘ�ʛ��*�F��z�G[h�+ڝ��¼�҈�m̔Z�]N�}%�<�N9ͼY����̺+�V#[�#�R��ۙ��KT�q���]���V�in��c-1]����v��5�X�8ʮ��ԣ]y���.���.�]q��[�:\���+�h^���`v�T�xü�̏���#�*ÍK:�T]�,3vm&k+�vw.�i�� �\&TS,���1�&�\�t�����xo�;�s&H�S .%[�7���1ݩW7���Gj�7dU���K�9H�g�V��o���
�;���E������F�� |���Ϥ�\�V	�[�Y�iԦF \����YwE�/�8�2�	9��׳��Yt����&����
m�ϳ7c�|��It�)n ���gKs�L۫����̇d����U����s�H
[Z}�^�_Rt�����p�x��s�&C�X7�g�p{�y� PX����:�"���X\ ���72��lPNG�jej�
���E/�&��j�'�}�ֲ�ZÂ��=	�`���^:yq���+4WqkV`��l��Z���b��ҳ��fM��r,�w]u���E�d��X+����M�%ԫ�zWR���p���P���NB��ّ���P
�z��|j	2_RQ�v�4��� }�.����+�삲u^㩭>ܽ��9�-�g4�Q,�4�0m�hŀ�N���Y�;�'auk>�ޭ��1ݪ�I���S_w*��֧L�q�8�Zwc�N���T�`Ýgn�T3FR�Ӝ�)��u�<��I�K��Ď�/D�9��jƱ��b,L��!�uf��2+'��q^��P�n8�I���`��غAؖE�<��M�e<���1pz,QdL��ے�����ⲳ�'[H`��<�(��;2q��h��&]M��x�Т����{�>�}�(�����ӭ����{.2�Ct�5�7��Z��E�d�Q�sy��eˬ��9�kq ��7o��oEY�E�o5��`�d�_U���w}��@v�QT�t�;����Q�V��1��uђ�X�q{�L������w�y8��U
F�F�����ƒcE�,BJr�k�4�e��v���t�A3
@lP0�"ɢ4��r��M24SI�M�Y�8&!ˈ�ۑC4� ���&@fRr��.sLP��!Le)�"���D
2Z2$��A	���d
	�ݺ ���,�LIB&��,4$ɦE)	SP`�-&�]�C
ȥ��L�ۮq���Δa$���I6c@�RQ0f���&2w\��nn�w��It�C2 Hcr�Q"a��2e��L��
.��$� P�wE$I`d��fY�_ՀW��[�VZ%��>巧.&+�r��P-�:2�ç�p:�>Y�]�֩�,���S�8�VvE��VG+��D}6���� o�7��6���@��o��w�����;1v%��Z�
t8S�Q�!�B�v��ɨ��\�.;)μǱ�Z�q�^�V�dɽ�龪�S��ꃫjO/Q��7����R��;u����=���AZPC|q=�&�/R��RO�V���f��7��ݹ�PP�o;2X��y3��S!�P�Wg������:1��կ������J�nr��q�{�^6d�T�3T�	��t��\9��܈\oӕ�(����j�}jhޓ{+\C���70��Zx_[ؕPU�n&���M>T6�i5Y�Xj��k�tW3�Pk��oש���>ۆ��)�Spx-�L:����dIպ��՛uk�V��ܑ�����+�m�ݨr�|:���Gr�a�@��LָN٘Gg"x����=�.��T��_��r��e9Fz$�9��Ы�jU�6��	�1.]��)ИЦֻ�B�g,�ہ��H��m��fZQ�,3��nb��-�Np�;7b�=���a�zX�ض��˷4N�L\6���{�c��R�Ac;�@�ݨ��s��Ҍ�0;b��}I��[b�T��7� `�nJ}wv^'�e�T���U��`x�{���޸�=�)髦Y�H5CZh\�y���^�J3b���u�J�I�i����������U�v����.�m�W��C�JS��A�v��*P��_'�o Ө��J�[Y�̤��r�x�*��ך��j�sY�k���{d�I��*m�W΁鯋}���,�6�K8T���}=S�=ert���]��n�T::�ܘ�S�^M���n�9����-uȺq
T-������W��1=5�j��Ku��^�]<#�/؟�
J�E&����#��{:��ꇂ�8��*�u/k�YQA�;�c�c�5����s4��K�>~K5;y=�d��*�Go�����f��b\	���6�MҚy�b�f���R���cu��^��`J����t��I���h���^c���k�u�8<�]k�u	;��Z��l/���9���W,��.�
��Q._ve봥�;�ץ���G��3��Z���`+���Y�@��~����[��X�ԑ�q�/Iʽ�FM��Z���0��;Ͷ�e�I�1��?}_Ue�o�{�=5����n����y��;z�����Գ��*J�`��O�6D�H�[�㖪��E����~��>k���5��YZRcWA�
m�V+�[v�!��r��-�����>Ue.��j7�J6�m�5�{ �iWi�D9 1�K�r��ڇ[w�mD��)D�W&������iG^ͫ��E�'�cWP���5�&79�q�髀���	ta�ZE\}ws��|���7	B�w�원��K��ޠ��w��LR�z�T��Z�{ �ảd>�e�[u]�n�vV�X�_��s��S��O��T<7��nS�.�p�:[��aF�6r����o�y�)m+��>��![�?B�so�_�Q�Y]�����ԊW��.^ͧ�)M�����i� F2�.�2�v������Y�46F�_$�J�\�����Je�=<�^y��ּ�Ҫ,Y���O��K/5���L��Z�x��6��C�F�)%S%���8�e��]�*j��Y@<��7h��t��d���M(���Lɿ^����F �� A�;���{�\�I)ٜD3s]�G��heU�����)r�Q���7�mz����K���&w�y���/�v�7t6��ډ|ʊ�Y�k�=�qz�=79��?U�����I����L�<'}���|����DM8����[�\��fMF<9M`�*�b%Z�B��m=�E����u8��q�����Q5�ۜ�ڨ��Q���s�t)jt��p���� 8d�r�mS����rﴬ����׼�;��K.�4�k��#�M�'w��L�Ήu�q5�dY�Qe�Дbt�M�YYd擷a]�;ya�і*���|�^U�D��shc�����Gw���VM	���c��v�VJ���o;�SM��+o�P��P����Mw59�o�{���B�ˬ���-+q�*z�׳��2{!��EWGU�d����n�0:M�UhZ��W�b+uW�_u���8�r�Br�\a��>w*�u�i�:.Z\��j����oo��8��1:q�[�B��ҁ�ح+ھtu,v#�-�>*�f�ys�T}�I�Px$yz�:�s0dZ(q��h��3���w}� _fH�S�Vl����
=��vU�)Բ��<u]���rj��?���)��ݖ�H��D������.̸	�v���/G6�M9��w��g����ac��^�ϻ�V9�̰�Xy�[J�,l��1&$H�n������6�%�t�GH}��cٱ�r�7�&_Q�s���V�U=�Kv�)��4��[杂j9����x�ޜXGƄl_=�A����=]+�d�)�'P+�.��j��\���e��bp�J+=��Ci{�v2�J<�o�`QKYڌn�[�����PS��mEO��3!�j�j����r��5��=*&#���k���4�{�'%��Z�Mѹ1i��ny����*/)Λ��m�Tb�u���Ңc��P�v��L�ݩ�3(4�=̜���|�ڮ�<�P&��L8���]S��^88c:����oB�׃�S"fs�Uf?�����|�W��:�jkUqU�N�[�������T���ɹ����(]u:��V-(��i�t	��yO�%���HYY��`Ѫ�͎�|"@���W
��Be ��!�4K����]݉s�,���3yЎ�t�mEY���Y�C�`9���m���*6�p�ʊ�!!|�j��}�c�y�]�tW�j�P��{1
{�����Ī*w�t�i�T�k}����[����4��;��j����>ۆ���k������P�d�g&bWmN��ܹT�]�ױ1[��_l�6�r���9�s����RZ���Z�՗���0�i����Ԟq?Er�7��2��O���]�8ŹS����@h����:�8K������V���w�5}4��Z�oc�����5�jB�Ć�m��Ul�xn3��e��R�W0�@��o�bV����ˀ��)<��e�� �;я)J��GJ&u�����AwI٤Y���.���°bWd��f�Rw��c�/�q�p6���+	��������1]!��L��{r�=�BF���J�sK��5�'��
�vq�rpz�N�+�rI�W�.f���M��Xq����4ļ��M�m)�ռ�ל�i�3ơ�7�;q�Tu+�TL�Q���Wl�y�����o�:�5hs2w6Ⱦ�c5c�.�l��%u�|(�x�f{M1�����]C�n�����Q3�9��]�&:�j�hZ�M�aemRe]jR��ԍ�[3�t\7��+�ژUvA���'�_W�
^���z�?�EW�hz���?#I.�*r�=5��-��Z���8e=����<�v��W��wN�Khz�mWcN(|
�Խ��i�fo�LƆ#����Rx�{���j�j��l�=EC�q�8�~!{�-S�����q����h��Ģisr���������X�v�4ӍS�.\b����+=�.ҵsw��5���)��Ou��;��z�mJ��	��r��jN��l�w��H���ro���Sw�	�7�u�`�V�uv���E�6�E0�f�ĥ�B;�~=��B���q؆�O��y�۩B��'-��u�e��%P��&��VV��a]3Z�;*Ƿ�)^h/(�9#W&�O�M��}�2��P:[9O�cR��ry��\�9˽�yu@)�JNw(+*urA�]7�8��(V�TmZ���YD�/\�-��������(����3D��]���J�ۥ��!-z�^�6���ue	Y4��FR;�,]���V��ҷX���+�}o��[#݌�ÑH�"�ߧiOMʷ1r$Iy�R��Q8y��x��k6:=v���Y�z7n����Jv�+c�{�B,��:-5�/n� v��j��X�a��N�:�kݰ�~���ҿ�p��*㩻���w�	�{��)=A�ŕ����lE+�Uo����jɮ����BN���/j9`���c�h�P��h�Jk��/��i��b��g�X'�T�7Wa�YJf&�6�̋!.�8��q�W�B]p}�3�ˌ���Z�}�~J�{�FG�װ,پ@�;0Ԭ��]b�ƻ;-X��n"�f�㥾 �wh>¶5[�FO:�?T��4�j�/��_oA�Q=�\.{�����A^�m�����)w/���~E��P%�8��Qkj����Z^V�?GR��"��w�Ѩ��P��f�I�@����V�qʣ7��^>�юOءs���y��Egm�5{��T�MNK��T=�AW؉�1Z�Y�Qe󿴥�:�53h]#�EJ���wM��K>��㺬7�GH���wwgc�g�R�[��gt��>������,�����7x����8�/z�3�"�QU�c8�n���5��6I�`V`u��f�a�v�a�t� �����>�ڟ;�Q�W�=�i�]<�u����6��;�Ue&6Z�mN��ۅiE�rf����-�K'���x�u�6�������qB�BۓS(����`̓w��m&��s���N)c��W�qŷ-FҞq���LJ�:�8�K���[{�ML$���.�Ҷ4�<Ю)r��9R��h}�+Wj-/ kү���qS�����z���.s�����P�B��ӑ��{��6�aȩ���<�Q�^+s,'�a\��9Iu�\;�
��e��}��;;W���US���son3��3� i@�.�>G�[�n53Tۇ�T=��&9ӓ_O>ۃ4���U�0�ڇҦ3{�}���D��F�q�_���)�N��8��nISž�u�C��fU�;@�Tj�����mF��8�Kw�t�����&����p4�e��d�dCB:�}�����J�r)��I��'���L�����YϮX��S7OV^��!���m�o?���߱�-qT�{H
ˬ�ESBrGa:�:���R������uMت<L��Y�}|��n�������a.���]=��]R�vwZ��}]��I͢�/y��Υ<}\��{ݻ0�����[�c�D��;Z����v0t�}7~]K�OԲ��	�|(߻W[[�_��W�n��ey7����=K�=���dy+���iں�k@��<�'uI;o�~��9t��O=�zM���b3��^XJ�X:����kU��STL�((e�ۍ�[���E���~M5��r��L>{l|��MB�5d�u�&*��4U�C\���W��@����}��Lj���B��c.윪��(䩘3��-�Ҳ'�NA��i�7�-�������d��7d�TЀù�p��a���ǅ���9��^g�u��=�t�{����kP!h�u\�E�k�l[� �8J��НR�����>�]u���պ��B�+q��.+9�wr,�����O,�)F+�j�9m�M�+^_��c������Fe��O]�DqY9/#8C�ن'ʂ����v��K�q|D�p+�Nw��mp�|�]�UX��s���)���k�%�XU6�˫��XwuF�ܹdu�}��
���N����*����5o��y�5�\д��!6R:��f!�H�
;�qؙ'lΠ/�x$�d=��-ܖ�0U)�`�`�RC�78��$!]W�������6���]�[C*`�j�͙�H��j�X�{a�.�SЊ/��ų�����(�|n�ȵ ���ǐ�H�R���>l�m�XOd��.�8�||ec���]��;G\o�Y���oBŘp��j[�e�ђ�΃��f]NG��e�c�+��Ҧ��g_p����1�Y�5xm��;���P1��4h�*&��"b��q�[a�e���o �S`F���+Y�w܅���������a
�n�2�g=���h-mĥۚ6��;��f��ޤr�"���ݙ;�8��o;*#r���fT�ۨ�����W$-�a%�6�<�/js2�7f�>o,��qn�,iX�+�R�@(�����G�P�2�@][�.���	!c����<C<���=�GH6r�n�C+�v8@���6�m����b/�*��2h�K9ˬ�K�6�=GK9
�$V�T��ۙ�}�t�yr�3������G%+I�Rv�q�t��R�����9�O)dV4�yvU�q����`��)k�%���p�����D�(����SRC������dG�u��v� ��{,ӥwUɻ�S+D��Wfm�kJ�䬼�pd���L��T�,��S�]D�݇�jno��R�AB���F�8�M}|8�x�5ݼ�*���"b���!ק���p!.��Di+�5�hv�O�C)�����)�T���D�'έ8�+�:\\�Ic�<��h�S//p�R>���4���"��Ԧ�&m])&�GK�����s�-CY��S�s���˦���[دFufwS���|�W����[R�G�ݞ7*ġ {s����J�1��TY[Z�-R�[ܵ�����1��ȫ�[᩺��n��i.�SgdfR�7�n�̙x(��;���CN���]�M�SG��+>7}M��(|���K�C;B���4�3)E�Ok�b�{��.�z���V�D��W�MIn��G[�iv���y��ڙ�Eٽ�EuJe��$�Km%̎�1=��-��UXך%a��0��$��*+�)�eE����D���.֎o	ݽ��]��G>U�w�Ѝt��ap�:]��b��H+j�bλ�x;�e	l�1]������z�*T��4Z�38��:%nl�z�)t"Km�Z�C�9�o}l���k�:ֺ<�gB�ރJ��NU�]����YZ9%���4C��5���A^��M�j<����T uh�|�=� �,v<{����$�*�oC��xz��+��(��b��͞���\4�&�H[Z%w�˙�*��%�@{q��vC
���~�����B2wv$LQM·v�0RD�`ђ�Fis�f��%i��s��,fYk��Rns"X"�'u���@R��Hb6ws2ۡ�fbB����3LdIHZ4M&P���w]H�P*7wA�Be$*%�%��;��AJ ƝۆɊ0�&�δ�DhE,b��	�4l]�!�I$b(��E�u�R	�@�;ǔ	�"y�<I�����0Pbv�) ���$<�L���(1!�b���HW.Hx;�M2�Q�nQ�)�
	�-tDD�SCP�P�|,9dǵ��������3�I�v�e���ٕ �M��W�T��Oq�O%]%7�"wH��s5�ߞ��1�Ҍ�p�9r?�$�X-�E�u'f&)1�T�.�D���չ#Y�l����y�6�Õ2�$t�'�
�u�5��q���E�u5�MG��-���Y����'���^^ʈד��l�K��	�_���)ݍ�'�����`�r�k�f�>��ٜNc��gHQKY�ݽPl�J�7��*�fry%\R�p����u�q�λ��U���'�tt�,��a��[-˹&��t����^�6��ڿT+����6��+c�}�yƢzֽPsB�_�rk=�+{emw{���,^!��A�=EAڨ��^�'���-�G$�a<�IK�{+�p~�\��ڈn�u��/0w�9��w���o�oN�8�,�W�mB�o3�i�ϩ�gV|��
�9�����}Ocl&#"��v���?N�_Y�Qes�����>}��oL�%&��/�t�'~{����*'i �W?bn���3ދ����o�_�5��S�%��-��]lv�-�.�޽����r]!��B�jK;%`�ט���Å�|+Q]�O2����h4n�� "a�Up�ΐ�F����*���)��Ѝ}$��xR�m���ξ�Xf6%(����]�k�Wq�P��/�ܰL��Z�<�u�r�Bۉ4�����.sv,�������K�[�ۿ��r��4�+�ܫ�	`�Y�ls�z�)�z�s-s���Y���zUB����]	�:�WÊ�(�P�s�R�x���o\5{k�\�]B��p1��.�bb��SӸn%WÍ��S}#��v��^��c{��#��]'a8n�y	FC�S�s�;�<�-E�@k�aG+ɚ{y�M<8�˧�*e�G�P���^�'	�:�R��ð���k*x�;�`o��������9ۚ�=�(��V3Z�Y�	]q���S��^]����|^��^[߯':��lUB�<�ŪB�q	A�OuFt㋅��|�rk��^�{�q�_<~^�}]���m��/}@�ԃ��-"�ʒ�?]h*�PBa�.��X�7��.��ݷ"�u��
j(`�c��u��S��[�l�c�[�vnmko�V��%+����e�f�v��ʵ�oN����Y�էh��j=UФ�۾I^N �n�s���c���R��j�^N�9�0|�JoϪ��;�8��S��Op��i��ݙ��K��6�p��/��x���<�c�_T��{��7�c���Ϻ}�ܣ1����8�	w�厐g�tU5���y��Z�c�y�%�P�FL��蓛����ڠO��j���UN�_N��k_�nt�=Ɣ���J�u���*����������Mv\B�+��*�P���;�1O�M�
���.�/Ty��[﫼f�1;��m��6��SM͞q0�6(�;&Θad����N��*С�rNq��o�W�;���Kt��:ܫ�0�4���9L�u~{�5��o�j�kc��/�S��]/���7y1N�#���4�w6
��\����nM���.̄�1"����G%p��Ԋjv-
�R�WS3	�bb���T0sۉ�~���̅Y�6s��Sv(���R|��k)V��3$��du��9���e������"8��;Hp�|�.n��6�1�Xk�r��r�k7W+�ڋ!ˏ_%9��u�Y�/A�D�,ыJ�ޱ��	�w��q�`c�f�}So�g#�"�L,�n<�p�J�b�B�7�j��g�ʥ��Phޭ�D�cIi t��O�6�7���>
��P'�-��nB�\��_�����5]����j��/��q���q!'j!��
�#]�_�z��F����5����}�A�Q;-���6ns�'���}��I���q���R�.����?RO���K����T�>�_t��X(�\3w'n��.=�U>��N��Q[��!G��7j�R��_'�=��� ���t��y�V<���x���A���Wq!r�!{iuN{��]��ʬĞі�T�9�{��ۍxz�f�C��~����ˍbGv�w�LԦ�q;��kui�Z��Ʉ�D���	]U4�;��'[����$���q��@��އ��΅5��Y[IN����z�P⧩�
�x��2M��nF;����lv4��d��V"����۩F+a��Ys/F�s���~�ҦX�~e=;�g��w(-��-G�)��L�����r�Ǧ�T��uᫀ��+Jc��l�_oVq����{��RW5���;�;[L�8_,�V��-38��f��g��Wu�}����huB�תѼָ��[.e_5!�RR��\��t��R���f&]�B�Ǐ;��ٓ|�ɧL�r�_�U-"���pe�F&��X�\���!V��N�
��S󹹨��%K-X���+]�ѧp�}:�P�	wAR�r�.�%���V�l�����H�!t9w��&�!Y�ԣ5����͚�[�����:Wk���#S�0-4t<�������M���3���y���b�5�b:B���:��>�*m�L_��T����s�:�����J�<�<�=�󱋽�w�Je�y� �C��s��@}O�_��d�p��\-�b�^NW؞��d�B2�����TKƣu�T��4�_ϑꇶf!���q�ЧM��uD[�?Ae�ӣ�P��{`�Q�ym�32�A/�ɡ@G�gQ1��Cβד�bμ��ݜ�9�͜�B�Cp-ȌI[��R̴��I�#�`=m�bޫ��돎tv{&��8R��guhȬq�|�{�V�v�Rg�F���vL�b`kk�h�A��.��N���h�}}�;=K��>5^�f��j{�$@�k�,6rr�g>	�h�&��Vj�����*��GR����7}��R�	E�5G|�����y��kw=���o�.�=9�ͅ����nC{*{�xlټ�����րVM���H��֪,򯬮{=�9�|�e��
��ܑV�k��ҳ{D�>�޿�+/[���L�ĥ�o�R�v���U 8X��o:*��ܾ��:��YݕVА�S:TB�D���S�d���p�7��u�Bٗ�Ӹ�Ҭq���'�t��l��	VդU��]����{&�t.ᎦJ���1�n�+__���-;��zu@a�զ⹔�}�Y�N�ml�U��7�#}�rs����;���n�5���uv&��/]��{t���/=���Ƞ+�Ӿ�d��ØKiXN*B���'�;�'�s�̼�3<W{u8���Xz������_;>��駱i:"fc]u�AR��Jw\��ì�/7�qoc�sl���Cc]H��k���U g]^���z�J�O*6��2�WŌ=kR����n+���>�k���6�i�l��#�gw2h��f�3;w�؝w��*�|�mv�RO�]�O�Tb�5�':�.f)N�u��u�X�f�%�[)�#q1�ܩ�O��m�]���ŀ�pŕ��\�l���%���uF)P������#u_{Зy�}3�ˊIydZ�����P��OT���]��t��)^��!�z^��ZW��o\�{m[�nz��z�w��[T����
�Ւyz�y9�o��(:�P�v&�u��(O�O���8�O��.��ǒ}��qɴ��6�.��'��2r�����Q�Z=�U�r���!{O�s�*���N3�zc�꜉����v��[z��_�bUhu�5�e�U_4��t�d���X[wE8���֚�Mʺ�Y
��y���*������׉[6f���
�UY�/�8����}�v^({����'�Jd���l{��r'��V�)���a�a}�r�WQ��\	3�{��fl\L^%��E��Li2�̾�i��.�j��5����	��;4��2�[g��?� ;v�s�+�콹L��]�V����޵;���
�F��؁�����9U�}3��޵΍NF��8��m#h�����~���\�ºeS�M4�[	vC�ڈr�@=n��1G6��ս3Ѧ��o�*�I�^��'n�?;���n�R������q���QjOٺ\��Ny�"u%�T	W���71k���/������l�{9��C>�N�d���,�q��c�/��â�ne��/�/*�����@���T�R ��;!Tsu��8���y���v�:"f^Qwz�f���\�ܥN1Pu�L�N
��Q?rvd���A��-��q]yz�
=�Yj��.Fs��9�
c:C���h�Ю&5�=90�5��ģ19��fj�8}I.�+�����Pb6[�κ*.-ʞC����"��f6��Q8�v]p�k��R�ſ.����ړ��"�0�8ih�	�=��:�� >��,��~��w�ҫ��B��j�>t�I�e�[1��P]�M{���hg���dz���JG��_y�7�]��z����s�=��3O�1���U�GN��i�X}���?~���e��q�K{������m�؝W�Z�(���"���߻�q��s}}�u�<X?{�g����� ��y+������W���f�Ӓy�vK��뎗��CPz�'8�v����R�	_�f��lE������%r8�YVg��Gz���iJ��w	���΄���;���1+�N\N�=�4����N�LS�Qes�哥;�p�*{�L��B:������#�l�c���A([sPbR�����݊mP��uK������*v�9s����(��ٮ���0�T��j~)D�r�7��/J{��I8�������jf36�{�����<ʖ��>9m�&��@]�h=S �Υ��\�m:������Z�b���5P0jۉ�\b�[�OrJ˭�턑�ռ�f�\z��K�ެl�w
�����BVj�O@����ih#�[��byd�7�q_�#�Ҹ	�ઽ���v��N֙&U�m/�OT�4fV��F���I�4�ӕ�p�]t0.�I�(T\L���[s4D��_Ka�l	Sx1u/w�q����u�&o\�G;�:��{��X[�V�1j<�-�C��:7��i��_u�duT�y6��_V�K,��ج�$�g2��L�Y�����1��W,�������3C6"���0�{��6�X>���ɞJЊ�}Y��&������L=����%׆����;�P�6���8�&j6������R���ϯ#3r7YwDYe���'��{�Z=��Tٸ�D�r�}@-7���ݭ�N=�8�{�]9>�q1w���Z�%C�LS�p�9�d�O2���{�E�{�d�e�s�"�2kJ���n3�#��g����h�>{#}7���	S���_7^�9�q[���gt��:�o���ɚ�A�i���S\P�wǾ� k����`�_1~��Ay��j�e#UKZ�vS��s�2څn�mJ��{>��a�WLa:�dςy�!��k��9�^g��^n�;��/"��-7�^���NDרm}İ�}F��K�	�}5�w��L�d��:�|5W�^S_3~�js#*r��MK����={dp�ڦ��{}@RFX�������'7�Cjsf��rb����w9�F��}�i��(n[>�r<W�K��W�W2�q�@l�9�DUH�偱�p��y�#�TKS���L������>FH�aڽ�>���z���&xδz�5��t������vslˊ��&r��S/���dv�G&�u��Op�-�+�<2�G��[鹄X�)wG�o3�dt�Ou+LZe���U����e�]�WV�G�l�1ӫc.�J@�`�{���U�*dCu^�ƀ�fr���o�� p�����u��.V�.ꅑ��1�hE�r%e��%�h��9C+���D��h�{;[�*:�qj������Њ޻dj5����-�It��u²�3t���1�p�$�,^�;� �mpv)W(��,y�C|{`�j��b�\WI�o��\��rJ,8nV�Q�|�v��}�N�]e�*�{��-N�ʕm=�느�`�pAl�]`[�v� ��3*�Z�|9���f|�֥��=g�K�o:��FYK+wSV�7��五�p!j.D-��Z۩�k����_=�qq�km���%��z7f���&�w�7���29���t0<��Xu}i��b��,j�Bh]�G�
���vq!Lg0*��a��U�WNj<��Y"�i3|��FCv��'t�}�ݻ٠[ �儫.�|�v�YdF��JN+�=��嗒h��W�M�֙\%��|�P�G9PCCR�uP�Xj����pk�݇)@lGp�cQ��ZR���V�͕!���s$��OV^?����a�f�����ϝ�_vq��V`Nۮ���)��zּ|�{�76�یvs�iC�o"��CC_`ǜ�ӟI��h��3nGs6��׎Վac�{�mr���ʡ]L��(=��=.�^
G����9𼷊�5�nAԔ�x1��Y�bu���S=�1�!a��Է���9�;;
ɫ�u(ySXI�ݔB�}��K���I˻�}��}��먣�K�V
�>(�f���x�0Օ`��zF���֥�g�u��u���n�D����Rn�h\*�#�SQ�cެU������1	�-�����P߂�:#�._q,L��Vp5��i�T7k�����������U�9{9��VE�i��7Qb�,ӷ�9,��2�&Z��mU���U<'��W8q��We2�:�}���O���,J���	"Yu��K[6�yr��ń�o�7��S�|���d���s�Vk�V@��t�����d<v�ˮ�Zo���9���7{�螻zJ_Cqu���u���q�A��Q{��.�fe�i�1:�':x)�w�k�]Y5�7PB��
�їl�u�CN�Z��G�Ԟ��s�>�b�(Rd���	c�����Ó�x`޴k�����wJ��EN�:�Ku��3�d�77z�hX��%6ʅ(@[X��'��{����7l�O#�f��x�a����@gw0؍e��ݢC�ve>��Dkr�\CTFL�{��X�+l��i� Ԩ��r���p�N�N7��u�/���9��JY6���uR�Eg*m��a��p�S�]eQ���Ib[g70Dr'�Eh6�D�����4�:�|���y�H�>����,���!���Ix.o;�"I;�.�I.��I��Ji�Q�xᄄL�y�f\�3��x�HB�sx�0�w\H;�����l�$R!��u��s�8�+�Y#2D���v���dQ%�;1�]ܓw�b��LQ&�r:r����71��Nk�3;�<�.�˰cA�QNWD�7Q�㝎\Fr��t@��.��N��뻝������t�wt��pl��\I㹻wn1����nK��wW$Qwk���"��s^yћ��ܹ;����a4�t�y��h�	'���.��:뻮t���y����w\�\ws��.rn�˜�m�;�;�����˿�������O�t�r�P\!�*I��>�^�:��.��t���AX�ھ���т=�h^�F�������,�_�xz�b���l�����3��o��	�_���f�bx7o�n}k�ς�������s���9�>
�/��.{��m"�7���ndHy.jjى��ݹ��~����*괏.>���ݑ@D�����wr����á�W���g�������)�N�٘s}co�@�b�.���ā�ٺ�14�������'���d���l����'ы#R�ꁌ����)����x��j��n��ղkK��7�鷜�x,�ht?^���E(ў��7�z��;36<�H��W���u��VW��nև�|f]���=�魨Ui�gv�x�3>��;��q���b�z*x�{�Z=�3�c��C/�����-���!��g��9og��֐�
s������k�O�^���8�CU�Sp��������#�����1=M?��<0�*뇹��X�٭:���d� �|�?-�/�=��*��_^d.�7�Y�6A>CܴS�>��VUCÓ�s��u�1����@J�Y���j�=�*��:�`��um���H��̻4i��K���y�}�|9з�5�`,�8n�bt\��v���M��篒�yp��S��^�v���xk��RM��S}��0H������8b�hK(Oi+"�V�'�X�v~R���gA�4;,@o�딹�+ן�o�Ylp���B��i�8�paS!�Q�����o�>����5��V�̿9{��f���X��H�m�k5�����mJ+!�N�.�0VEU�1}�q2���c�^�Y�O��糮|̏+�޿aϟ���v>�O�۫WXՖU��
f�Z�eU����=	�Fu�x*�K!E%����5M��.9�q��:�_�eK0�\S�/(�/�{��ۏҒ*s�Z�ET���l�__�2�>�aW�~���lg�蔏f���z�Q��"fV5[�Ud�,t��ޞ�B�29͝�ݕR,T�U�����ͨkr�Kґ���m�/6'���v��K���]S��,z�oFG�����7��!���#*%���݃ǢuC�t�y#��{b�-�+��'������@�=�r-̹!zO����=���f@�����Owq�x���v}��*:�w%���+�{l���?X$TB�;��]����w1��5p�̇Y�H�{����'Y��B��r�M�7��R� zú���2��q�B�zG�^�3�x�~#JX��q�Z�K貊[sq���5܂�ƺcΩ�t�x/=�ii���^oG9�TwV�p���D�f���lz)ϯic�[��p��m�S�\vᇛ�`�%�$V���:��gc�S2k��γO^K&�\�3Q�ǩM�F���O�
�fY�?e@��Lα~^��u�г�cU�>�>���ו�cٳ�=ޞj6�c���d�Ϥ�vsY�W�q�_�%yd��^c(��X.�O~��|�����ͯ'���=�L?M�ؘT�~����s����d�>�G��ؤr�nE�	�_/y�"��xvuH��ۅd�\�i`o�h4c�i�x*�j��^�W��=�b2���}~����|/���w�mh+*�ʌ����9�/b�9�u�P�H��{{f<�C��q����\	WM9��Oq��{Gj��3��	l�Ku��6���ߤ��-�T�����Х�b�&w��e"�:d7>�������+�nZ�����CȕT�V�=�ZY#�G�98���"*{�
���o�a{9�,�~�g�uG�^T�b���ޱ3���������:��W��'>% �棠M7@U�^3y0��_�P�9H�uv�<l7ۛ�ҷ8q�Y��7��4W����2
ʖ^F���`{g�Ⱥ������mCE���RMG����Sc��l��zکs��!T������ܱH�m#.���^S�J�ZL�7V+e��8nT��U��Uz�q=�6p��S-�.�Y��H�q�<M��E�ބꎇEf���3����)]�)��q��:��R�N8��Q�\+��r!7VB]�j�q�*�G��,����__�܇�Qhl��
gz�FT��9�C7������f}�ϊ���T{�)�j��î�x�N�(���H��=�r-̹ j�3��nA(��a��͏v\ﶱto(�%�}�9�FAr��@,eDw�����1��{�8�ՠ<��q���H��c���i�|��iS�u��וm����,eb�%��zi��/�=�Q�e�����нb�ɘ�wY�uE�܉����F�i�g��֗��}^)P�+�UG�x6TJ~:(�o�n���̮����x���@T/X�F���o}SX=�>�ڇq�^���3�mC��+8��}t6��ྭms2���#����{ʛ7蒎\��Z}=>ѻZ��[��P�ȫ������]�.�},.��75� g�z��vTM{�e<Oa��(m��FB�A�f�~+��Y�h眡Zw�b����N�o׵������s�G<���}�<b״�q��ɕ��� *��"�Ky�*�ʈɭ>�L�7��]��#�}L0����l{+�{�Hn�W���� f�*..�u�3���-�4!h�{f������W���<i+�Ɩݼ�ʥ7GJ_o*�/6leܪJ�$�#p��n�ݵ����R�Ċ�9&q�\��PSgL̊��L���"��]��J'���]{�Мc���McT���L��8Y%͘��<��};�������]1y3��>	��u������w��(��$�s�r�����/�֎��ք�D�����Q`Wz���e3y2���0��÷m��G�bw��Iv;)��{/ÅëV�AYR�g�@S�.��"��1M�>NJ-�>���3-,�~ް��<�~v�����q].�*+N?O��k�B�J���f�>�����މ��B�fx�����`yJҙ�,%}Z��l�z�9�0�"�n��ez�1-�gey	{w=��G����Q=�Jd���g�r�x�����^,lm"�<C.�=��3�I�/����r{����xR5��,{o� ���8KGw��S�|/�]V���Pz'r.m��iT�P�y�A�F�l*�l�H^���11O�h�ѥ��`�xW��:[r3����ʑg͟D݁�=8 k�*c�̛�/�#��)���f2<�~x���?��~^@��ٰ�̵����C�U���1���se�H��`�C9@J��K�7^��φn�hq��c���� !J$)�+e]	����zY#�\m��عee̐^�iK��Rڭ���W����)��0ф6:���u����ι����5ΰ�X����U��jF��-�uM5�夝�%[)�r�)�B�4�u l�͈i�c��V_s�.�g��F�F��Tu��zX�3ZPU
������.z*x�o�w���V/�S9��S��,{~ۄ�F�A%
u=������,��W�<5N;���zT���5~������^�	(g�F����E�3��ϧ�3������/�Q�@�\GScU[ Z�W�����/s�+���$�3�X*.}���m��'0�Ȋ�xk+j�z���5�uH���� �=x��e5���S>��MO��Z;�e�jY��}Z4�Ϩ�������n0�gL�L��sE����;j�܊��Xy���z���������Ac���u���*�	����<���ާw_��ѧ7���u�ǡL����w�/���>���!ի�k*Y����n�}�o��WP�ί]�:��1G���
}�Yl��-���:�tf��w�?Q�C�TzL�<�h���oIi�ښ�kg#ۇǕ �"�E����J�u��W������D����W�Ԙ2�]UﮣZ����j�u}-�zdy�����*�X�^��/���mCU]�׷��_SQ"_�iW���A��N���S������=sV�1db�5(-�j����b��9
�84��q$����hѱq��o7d�\��� 4J7�����X�;+����V^:�y7%�0�ъ��G�gX�(����$�γ��紲��Ęy֮����]��t�jAv��������n�[�zn@�>sqd��r������9�wr��Yc�&*go09N��z�P��G{����n<�^�`�{r�[�rF��,���YDS=�'�<�����w�����l��}��RڤB/��T�����$Z�!����/åvq~�ޣ���8Jb��癑Q�u��{��ø]^���BT�2ǡԀ�S�2'X�;5�J�/��9>�(��fd��d��j7Ӡ�F����,V��o�'g������, ���~�X�Oh\*��	��	vo�)Ȫ�ٵ�a�ϴ�zx��`	��x\jWr�1�	�,�sr�q76{�1V�vm��|hOڢN�����n����q�U��4����]�r�ye�b؜�F�HMR�>�$�Q�LJ7�ݺ�q[��r��ݦ�nZ+Y�4�����/fe�7�\��L�
Ug���ЋQ��no�Zu��U��s�o�xH�=�:
����I׌wG�{н�������z�s�	����U�N}Gb=��}�u��۔m��-��7Y38_�<����K�����t"$t�z�_GV��3�_s���A>���i�����U�.I+tm���y��$��]���y�lY�S��0��q�6E,"ԩyZ�ѥFYA�c#�(Eh+7q\tLn�_�	���}ܥa�]��T|�F�6��T�KOIT�A$o��~�L�_�3��dϑy2��+�����x������\yf)��y�����5������$�ߎI�7U�Q�@���n2e��e����ё��zb��S�6�|j��T^�$.�����*������½f�`>Ț��?StZ��8aq���h��}7���UN�.�*��-��~��+������V\�����}(zs�2.���\���B�9��ѻ����{�6Vz*��y�z�S��{�L��������Z$6l�g�*df��+(��_^Tf���*���h�7���5}���_�p�w�G"<�C��4�`d� oʼk���o��Қ�쩔�Z�)��W���f�W��>��rc*>�W\��s�{�9>����.&��"�������לt�̟\�:A�!���C�&)��8φ��Tj�%�^�f�/�=�'�@�t�HN��Ww�!z�^�n�
]�3p-D������F�i�g���z}]^+�BXq�o��s��6'w#�к�gşG��<���g�Ay@R���h�|�EM`���wj�=����c����1� `ͭ(J�h�-��b���]k�^��~�j ������s[]nc6���p�K��B���(K���AW"|fq�K�5ܷ��f���A��c���q(�W�����ͷ��}��B��ȗlM���	E� + q�+;J��gd��z�~���wZ.5�ܢ�:z=�=���w�J9:������e�uho�ϲ +����k/�]F;ݻ>�|;�o�(.���o�תQ�\��{�eGǧA�1�]u�ħ�qy7S�ӝ7��ސ��Mq��O�i�Fz{�k���*�z`cw~�;ܨ��u�������@�˯R]糧؏��ë"*�2�&��\d��޹]�H����j��[���u�P:\�]Q��r�=��~�����m�1~��ϧӺJϪ��k��:��ςyR�k��>���>�]ή�ݬ�cஷ���c����{6�Y�ӛ�8�1@dWz���e3���f��ѻ�UPxW�;k9�bao��!S��|��}���কxt�,�{�;���s�6�7p(8Z6�)G6���V���ud������aƹ�.5��\r7��ߪ�~eK/#L�ٸ>t��z���+og�[�:o�?}7Z}��x����aV�_��������F�:���N��������v�/ޤP�w��1(weT����Å�����W���;����H��1�?R���v��Y�4��*����{�v�j[�#��\���6L�b�_��֊�z�e��Ԗ��wU�G]�k4÷h8���0�%")!j���t]o�vk��ywۦV�y����gI��p��Wv۪���Jnj�}��,GZ�}����s��;F�&n���
G�tO��P~�}^G ���	c�
{����������|�D�ȿ]��+��3���`�PD��	U�x���Ղb�N��/Ǻ;7������/���܍�͏)P���������vX W���<�]q*���3A��ݢE��I�,=uI˿Hȵmpu+}�n��<{N��u�o���H���=�>�Iu��Uexl��]�T��e]�ls�v��*bj6P�3_i��D+��z���.z*x߽U���9V.?��h��I�?�x3Ўjh)��iS=Hg�gt��'Ei����f�i�]^���U� g�>�7��Q�܋�9��̍�����Gw��qȓ�;z��۳�XQ�5��\���`l)�@����	P�וw�J�2�|��,�?o�5���]�'�0�ʨxk+j�z����}$xe�/7=���%�p7��;�G��%޽EWC���:CE�M��K9��CJ���b����;���&r Jd�NxN �s*z����φ�G�X����޺�����dGz�*�}@S��dUX�Cм�үQ���-rE}�:��u�͋�t��Uv^���ĎK�E�l殳t�$|�RrĆ�$Ԯr�V���b�s��Z��r�7X��i�{�Y�<��Y�#Ȼ1�����J��G��*��<yiV���=T�X�:�<�#C�;�ƮX�K3��Sj�1B�;�C՗�f�Oag^�m�u*�����Ct�nőY��6N�W�2�E�n�إ2	�RIn���kd��u۰���#g%���6Д������CV�����♍��G	U>�u�&T��9i����W��%�䩠&��Q=F��]�i^���͢�%o��a�HM��0"���+�A�O�f�i+c�®P2�W��t���Qˋ�GNWv�s�;c��ͼw�:ӭ3z�(BV�m_ۛO��=��+���%�>B�|0̊�} ��^`�rC�ޮ���48�i��s3�ko�.�
��:q��'ʑYBIׇMf�24Fq�g#+4�s9T�&֮��-Cp��C;B���<5֯*�2��wM��;j�sK�ؖ�"!Z��wB���Ԅu��ם�2��ke���{n�F�'��,9�z�ձtz˚�.<���Ũ�jz� 䂵&,�i:�xdɉ�\�[�4k�̻N�k[2��X����ج�tccc���n�!X�N ��̫��)���*���:%�z�������cE���7�GSFܫ�J�',�t��ݐn`CX}��D�?Z�wˤ[θ�<歡hM�\+v30w�\l�7\	MJ5*w�t�Y����5��e����U��v�$d���WN���z����a�y�㊞i���b��)�빑��LK���x��Gh}]R������t��l�$��'"�t���H� G\�qdy�Fvrdφ�݀�cϖB�SkE���N5AVl��ӛ�������:ҋ �B���\��?m�SI$!��4�oog׬�h��έ]3��x��@��u�����`���<,�p�ݠ�<�2��WˑO�P��7��w� ����;�^i��|�Gd����ڋ�˜�a��6�fQzd�g^ˬ�JU�
���O��|9�+&���9]+�v�-�i�EmG�n<���T���j�jlZ�r,���á�6�U{l��g__-Ii�y�d�o,	��M�Wut���vZ�H�Ka����
��Z�+.�g���rU1o݈�4�V�o���w�6�4����ݑ�&��}�j�r�v��L��r�wVV��v	+�%퓩h�������ά���.�SZ�V�T3��ə�����>���N��qڷ���J�)�Ǌ���r�:��װ�3�������n���qw��kq�w��X@�oZ 2����.3(�{;��;�Y2���x��O-u�"�O.��^ƅ���r�v=�����s/V��� [*7��w��z[���q�č�����wv��L^�ۋ�$�����\�y�-�ns�������G]�f����q�ry�������ss�Yݻ����k�<�yss/:��ne˵u%�wWs��n;�e.�v��\�;�S���َ�[��n��+��k��s]ܻ�q�ı�r ��ܮ�.m�v������s�u�]ܜ]��Gg�3\��әs��7H.b��'wk�t:trN�HS�Wws���dT�sGs���wd�w	���Ӝk�tn�];�wu��띹����q�$����G"�ۨ'u��ɜ�H�9��K����:gw+�aD˻v�uۺ��tv�.��鹐���6ww:�u���s�lw;~_��������d|�|;�6�,�:7BczB��|���RLL�:['6����45廡�Vtx�0��[�.������2o(E^��5�c�dϓ��!��^��?K�h�{�G���q�Ig��DWUZ8�R����W���9qW�)z����DT\�/&[>��X��Z:25ǫ��{��6��u�2w=�X�~��_��.�᮰����r�Vnt슩Q2��ԯY�¯�z�xc�.7�=�����2�`c='��Ύ@w����v��z�|rzy�UH�Q+�b����ن�E�qctlW�jd�۰��|�\�>l�!����������E�W����>spvHO�(����g`����x�����UO=�z^z.��y�z�%��NO�=�`{r�
�L����G�=d{*8h:gz���y̚�h�tb�|�^�w���w���|�]�����Iw .��*-�zH��TCG�/r�V��Z�U��]]�~w?G����^ׇd�WʅC��^�����<�~�p=_�/�a�5�:��ƛ�>�2:�GL�Gg�/G�2|:N����Lz�SD��G�6�	����w�9�[F��2+j�_�݅u y���F���ʮ��dmn�w�^�}��f�����ݗs�b�-�vP�;�	���LLf\Xtn2}�ܵ��1��u\�s�v~��TTd;���"I�Ï;30z���u����P���=��]X�H����:�Nu��`H��30���-uftHs2�0i��x5n��<�V��*Ȭ�kb�AuU��=��t�>,�c�'�7޻G=�X/�x����;q��i�醣6�N��̦��r�c�(���x�� =��v�d[��>�ʡ�{�kE�߱�;t�0/��&W��Wb9��@��q���,{�>g@�M�q�� *s~2���7g�+}�<y=���'�Z
�)���9{ghf-+ѵ������ɝ�Ƣ��G����-������}P��F�ﱋdb�;4�w�#��rϢVփ�U`M�x�dγdϑy2��x���^g�=��%P�r��F�Brw�����&�ѵ���}�Lܹ�\�U�G�"�)�ɖ�#��b�S�h)Q����<|n)N�7�S��ˍ�=��� ���p�G�6\�g�Qp&)��^3ѓ��x��t{�3P��9�^��^��õo��z�;ⲥ����x�=��2.�[�3��`[{泌5��������S��G�ks�G��~���}�y���'E}����2���d�ٿ��l�Fր��_�#�v�E��P��}��&�x���9�>��nz���x�}�0���.ED[�r@~c0J�?.�m[6�;��}R>ܘ�I�4?���s	�*{o!E�N��V@��.L�i޻������Gٵ)Q���$&�Z�4��B��ZՀ<��u@�'#��3��գ�;a�r��u6+�N�Vԭk��l٢�+�����T��Q�T��nu�+�G�D%���kǙ��JӰ����!�J�bڟzf�_�@c�}�=q�~*Ua�7�r�==ްH��4]�{�V��g�u	c*�,R^�f��I];�xwI�o(ME�@����� ���w W���
��OdD��=���0���t��/O���4l^��n=z�f}�>�T��m]�8��S��9����Q�u됻����ڇq��=>�x+�:M�䅪L�2�1;�CT����x߽U���Tپ�IG��c����yP~3�N�E�sVܵ%]�h�|�V��<=�7X������O��\����5�����;�z�=`��퍝����O�/B�r2�kOabp�������U���n}�+�v�FC�F���,�G&k��z�}���,�]7�n���>���@g�������^񩮉2OT՛+��s��3�/�+����dF����>�����a��]1q3��dςy�T�:��{����@}Ѻ��r���<))Hｕ��j����i���9��8����&����F�FEg���=~���T�Ia�嶡��&���`=�����c-�s�"�JՅ=��PԱb�5��]��w�vϹ5p���4P>U�A�6�yd�"�I�X�Ɍ0w^��0�n�T��V�=���M�OJY�:�vP������"E;'vI��v�Q�;r��1 �:�;���|�c�4���x��e�x\:�lVDJ��_���2�}7x���Pz*<$��Bu^�Q(+�Е4n0����w����Idx������^�+*Yy�@l����M��7B�����x��T�*X>��5�l��"��;��[f2;�ߎ��7�uw���o�u�Շʏ`�F�J�/&W�Å�����W���;����H�38��:+�g;��U^��`���S]wʚ��b|͝����#�����;�ý�ǽi��a��c|�NO���P=����n���
��6}$/t�`����m��{��͍�����Q�]=~����+��M3p_�v|U`_��`y�*U�5a���!����5;An{ܖ��(vG�qZiP�t��6o��@y�uX=��P���sF��i�w�P4&��U�z���:N��������N�5���d֖=Qk3!�|�T�b��:���U;���bTZ�,�ߊ!�ԕ�߿����}��=�]~��Z=�D�؍s���`LGW�</Uk�O��H�ǵ�]�&>�:��m��jgNx]:��ӷc4#�8��5/$u�/r�0Ӄ,�UӅ~�S��w�4���QR@z6�T�M>�H����uem��Ky�M����'�8����G�f7:L-t{{{*�o"#�i����;��J��J�7���W%lW���{�?@1	���3�톿5O\��k�.��S}bVղ�;mGM\�fE��t���~`z=�~/9���Z/�Ew��Hë"���{���q�@��&�u�DU���ӳ����c��+���v��?WQ疇�B�L��ӃO������ޯUه�E�[�@�g��|��~7�>}�P�k���/�	��]�r%Oh
WV
�M=�e]qԻ��П\;��~���]/�!��^����Z>��.k�1��ܲ�AH�%��ܫ��#�(�"yP�*�	��W>E�%�䓽}T�ю=+O��� ��N��P���^��k�ګ^��E;�c�I��ʩQ2��J�u�L*�V����M�=w�����dǻ�΀����g���i�����UH�W��|K��f�4�%��.:�O�s۬-[7^,��*�m����� ��{�졐嚏_�r���{7�R������x��ۖMf?���F��ƣO������\
���@�ۗ"��uNH�^����tJ��C�T|4*
=�/ �(���C1�"�E�k#xi��{z�7h��V��3j�p��X����^I�`��J��k�΢�:��p1{�嚨J5� ���j�y�v��I-�qt�M �IemlN���N���z�ؖD�]ɪ]���lp�u}��[Φ���5X���Yn�]H������y\�;��=�5�1�����/��}'b}��*~��$z/JQzmc�ǝ�Ʌ=��u��nI�V����|�P�L:��znb�o�<��p=a�Į>*.��M�$���X�[ ���&â��7Q�[Y��O�I�t�c��4K�z���ޗ^�펇�s�ʬw�<�uTu��Q��ތ���ͯq���3[L {�f/L���Lq�8=ڃ���>���D{�NO_�T6��/i����#���i�醳j�䇹�q�#��՜���9>�L:���爷��,���ۡp���_���V���.zd[[<���;y��1Rӝ		Xqs��T�ޟ�xzo:a[���7O|�z��Sǡ=��ǚx�E�1W��{nF�A�g=��U!��Z}����HNo�3��z�J��\�����j#�n���,�N����֮Ϧ��Jt��D�kAYV��cc&u��&|��Cq����יqa�9�-��d��n�s������3��r��T�f�s3@tT� T_�3q�,/gS��o��>1@NB�sG9�`j�7x�P��sev� ����P��C�/��"o���ي[6>`�0�X��7��2��,�X6�'1gή�_]4�3	ECemG��b�<%h�}%��L��H꺵(+��`=y�Y
����n��)e*�4L�*��AG���j�]����+�=�%����#�JtA\]�c�\����DME�����J�ݛ&lP��]���w�t��B���������@`�~�_�dJ�˽2���@{�"����Ч}��s��i��U�]f�4j�����sސ�g7�:+�����3�.0�ѝ{[��\Z!�詑�N��̈��3e��ĮKW�7���oޑ��{r�,=;�C��Wa��8=�>r@HG�D��ϫ,�������>��p2�����S���铻�uK��e���]�jU��<� �_���/�B|��L{5�MVѽs�=�X��`F���z��<w��4�ʡ�͟G�P��e �<n�
�����T|��j���i�q������(��ꌃi����C�]��t'E}���m�����x�9�j��7q>��SX=�#wj�cR��`9�;ԵG��������}���w^�ܲ1*��_�pW5F�Gz$��>��8��:�ǺP�tn��B����֏\d�lޖ�I��,	�^���5� gz|����k��(��t9�<��y��ڥ8�8�`�{��?Wh����mJ��,	���Y,@�)e�H�}��ʣ,���vb�T�� �z1C�=cv%3Dd��s����A��I H�8�dV=��62�ɜ!��J�N�E}}]7 ޳�^�kG#�4�Ӄ#�{�2�Le�l���X���J��>�>�TKq�둗5�^O�i�Fzz#�j#S�s�������L����W�N�Z���CKN�����³�h��O�aK>�c*2kK�;㬁���G���6$z˞��
�w|�gԈ����^�W�{-��ܣ�E6r}:��a��t���dς~��ڭ�6j��N��D�˗�E�],>��x�'��C��
�\ڒ,7=5�w���޳��Sr���^|������мs��=��W�[���:�ld�,�{�;.���ދ��㋮jfǻ�	Eֶ�m�����e�޹���$n5�>-�O��J�x�����&T�o7`�5��5J+<��A�@5�R.�׀��S>f�e�Wա��l���
�9��@ߢ�6�1����M�� ޑ[ޅNRG�b���yT��-�q�<3�hU*��
oH��|�XH�?w�2�i�p����n��9f�\
�k̈<�D��3�KGw>Ƕ�����Lz��Ѫ\utyӫ��>��+>��@w�̂*-׍�S%���!{�"�LO����B���2��w�[zi;m#��r�I�+K�'8��hoMT�iE��!zS�]��t`Ok�0�}��EK��HM��kiM�F��306H�iw@K���X8���<�eٜd�˭���u�"Uu�90Uݵ��Bk9>'6��r���
������cp�b|9��!�@��X W�����5@j��L�c�*��[6�^��nU�n@p�d�/�WI��JҨ���T&.�͛���r%�`�|�P���.�{��~7�O�*(�A�롃���uo[M�Ɩ>�?[35���Ю�Ƭ��Ld?D�5�U1�c� ������Jr��}���>��>:�z�����댝����ge��^��Uk���VQ�73��b}>SG\V���s�W����8�n'����ƿ5����I�_���3}w���.�����W���Q�� =�v������EF{�h��=�r'�0ꙇgc+j竬���u����7���uoOl�2<_�����������������(/��K=�>�T�b�X�3�*��<�X��/Fh;��}x��2��w�������q�mW����:��}@S�z+�!Pr���>��AW�h+�U`M�q�%9�'���2�>�~Ӟ/���d��«WuͿX�����t�j��𹳞�@W�ϝ �*�	���|�2��9���h�����/�
��V��Xl����̻].3���p�,܋_s�M�Jʠﷳ][]��|�c��[1�S�6�1$�c��L��)�2����>�ݏE��_N��Z3l�����m�j�N�\����T.6f�+�_e�C�[ �Z�2m^v�u����{����wN��@�C��*��Y�O�v��E||��U"�l�H�9��«�_C;6�o�A���k3�7z|��N��<}��{a�/��[��(�!����>ʩ*%z�Y/��z���:ܣk��M�(+Us��S�}�u ^}��4W��w \C��ø'�n��d{���х��+�UG]ypeWr�#��w`Ǚ[��k='<��/<k@��&)�9"ר��"��E���,�첻���e�����zw�;� ����&<�U3����ND����� :�`�W���(��[�<��t\�~�lvn���V�����XʌV.>ʘ��B�}���'#o�^��u�1��#�[~��]^��2*�E�����ix|:N3��K�%��<�_E�!N�Z�M��B�{�5Bzn=顾����*��~��n�_����+Ɠ����X�אK0n�2�{rڐ}
� 	T����E�ϴ�?U��ب�xT�ܙ�v���Ӕ����sU��gO/PI�]��k�c�}��=7Ԁ
�_B^���xJ7�ݺ���Z��������g��{�rH�i���,���R"�+(��`JAy���:���ŕ���ðY�:k=eH���A:�Ž�f�����[�ڻ-�SVw��9����Vb@����ŝ`D����S
����p��/�(3	�c�vˬގ)J�dc-�L�hq���k;�����K�.	���sҳ�vu��p�+��]���o��;����״�����
4�岇nVSyu�:����{6�;ĉɏ�b&�ٗ��"CCY���e��mbͳ�;:]�"wQ�F�9F���x^*9�ϯ��-w}0;[����m\�x>:��z���6��3��v��db%��:"���@����'�`����\�}�8�����p�X�8�4��.YK��|��ɵ�ȥA�0�9�-�i��C�@�!{��rW.��z�}����aG��-ĻN��+�ϱ��2m����_pGt�&4�8P6j,�t6�R�|�k���i]������k0�H�`
��w���v�՛�(���lVG;��J�1fn�ϓ/����S�f�|�}��h��i�!�MR=���#�K���K��� 
.���g�
�M�&h�3X�6����Ү7g!׽�j�=S���f�;ZD��*J�C�v�QG^n��C
�+��GB̳WM� ��DfRn�qɱ�t[�� ����V4��T�6ع�ud��ܯf�D�������LE�g=
:�m�Sr�p2Ž�;eN�s&�=қ]�s�(��a��r����p�h�f�'�I�N͡�i�cl|�i��ѫYG�tI�TY�'L�2�)%�s�N2�B�)���x;���4#glef�f;�u����7�/l�-�̽܆��*<�Xgi����?#��+��F��ubtٹ@S���H��f�h�j=�*�r�>�+ ,���R����xQR���y�,��Xw8��q����������Q��:�b�k����@�jՒ�aP��g=�,�W�)�42P�sUm@a��p����u ��IS�]7��7km@uRv)��f�4�����;�>����,<5���pONW׽�%w]ײ��)�yZ��E[j�AL����uWr�k��.���K�/3cɾ�@M���ƧJ�2��k..�ն��;n�
oNӶ�+��h� ��ֱ$u��[�v�W;�#@��Y��I�T��r;R���r%&��-��@���O�
�\�v�����M�����
60�E�tc!�$_e�Y�hD�\�v�Xu2Bt�8�#¶Ō!(�U�����8�{x*��Z�u���øX\��t�(�;@���P�Q�%�N;\�R���&�]N;���J;�ӝdm���Ҟou1i�zۏ���q�)���X�-J����
&��G� A���J�X9t9��wQgv�]��\�L%�)9r+�B������]��K�]Ɖ��\�8]ݤ���r��Www.�;��\�뻣�&Ww�v�t�w\�r�ú�w]��:���s��r�8�\���s�����Muݻ�q2�㛷+�i&!�����ԗ.��K���B�q�	�.]�s����uӸێ��2��;�N\`t�sw:��뫘�uƈ7;�w�nD�q��+���"��W;�D�v�NdQ�\r�\D���sww��w;����"'n��t����ArI���u�v줗wwur�wWM;�d�w\�;��v�#wt0�.nȐs\�]qݢ��MԝwdI%�S��b�AK��.L��$��&��DI�	w\�1DH�7:!�@
��%Ж�@�sU�����.ܨ�se�{�3��n.+A�p�O�R���������i�ݸm_D�$�b���FHo+]�SC�~��o�~��.����t��{�;�$o��6�ϲ��(�{ܝ�p�ofP��ൻ�5�p�W�TFMi����cY	����m�z�L+�����'��y���\���/�~ae�zOꑭ�A�?Vy��t�1s�,^L�73�_P:��O^��~�#5�X������[����
��n��8˛��(� e�S8Kو�U��L���+f�x���z�f���g�^�n��c
��;!���n�욋�4���r����ܨ��s*�q����v7qW	�F���.��X+޿_�L��e�@!�(zo��3���y���ھ}�C_)�s���9�����mCF������sސ�g#}����E�Uz��~ȹ4e����T�D�����/"}^G3�XZs6_�E�T;�%���'x�o�zC.!/cq`zB��i!Z�%\H
|e� hx�*���s�:2�i����W\��s9Ϻ��o�����tx�3ݳ>�s�u�ِk�5� \B�->��n|�	���h�>�%��F�*��;���k�Йwk�@1胅Zޘ:� �\�V�\�:��,�rց-,��lH{�r����Qu�]����S�L��U��JA���8�@mv��ݥݓ5ӚS��N��o��J��ܷL n�\���[T2�71�pӄu�خ�X��OU�j���h�Q�*[W���u7Б�<���Υ	�ty��r��<�bN��z�5UQ�ɫ�{�Y��W�
���ږ�Y���^���|�_���*Ѣ�	b�UO��~�<�����߬5�ϩ~�m�N��:��6�H�i�����^�^��u.7�q3���w^���O���w��{E�Y��IG'T��c|�
z|#�J��ݭ
�'kf��{�a����c3� _ϽS���Q;�o�_�mc�Z�
s��|x����O�P�u�#.#&��>�u��Ojwb�{=0&a)��C���qX�L��}	�kM?���C#?e��V�m,�=f�g|n5��G��{�D�=^�ʮ�\��\�&�#^��B����<���(���Q>��VUG��+�0�gsN�;걊�\Ձ[�⺫u���r��ު~=����uv��~_k�No�s�9ɨ�l))���I�[��9y��9����&�Q��6���c�G��{������ʖV{�<j<�
��g{ǲ +ΝnJ�`�E�n�Uϓ�6�Dw���t��G�iQ�|}5��B*}�L^�e�����x��-��̬��J[_�.�Z��L�*��VE�rrM�^Fc�
w�Ϧ�oI����Ds���ަ����m�Зx�:{�)�<^2xR����3��j�d�SZ�ws��M[��ΘD6N�J�\ɾ�&s�O#;���4�_qW��tޟM��@�>�� �"�E��.�S>f��s��~��z�:���Tm�&�r5{�E����a�����.K�����R2��^++�3�Q}\�Dtz�B��W���˖XO'��d^�ۙ)�9�Y�|���(>�2%�y%��{�6Ń )�1��k{��{�:C����7�S�U�x������?@��75�GyNDV	�{�t�m��	kV�{c�5���P�;��1�4���i���@{����{,
y~��U��n|�!U�=������'=c�Y$m)�>���>�G��	���ue?H��e�[>�z���9"h�>s�ؽ�������Cg"rXی��댝��cL�ic�
��ު�鋇ފ�;#,�cM(T�/�X��Q�״Z4=��ţ��x�EW_ṳ�}q����k���m0&:�q����s��M�!��*F�mz���җ�#'�<�ي�x�9q���G�'4��͚�z��'����躲�ҁ+���
k�
��@g�W����oE���碻�O�aՕP���î��b�S��"u�Z��[S�RF�t	�o��':W(:�]_K�-[�t�N_KKi�oc�'�.��'W�/O�e$��36oϻ�4V���iMA6̲x�m��mt�:�s9�ty��Ãv��ʋ��Jvk3ݧ��@�_T�6��
�g��b�s瘇��lgۢX۟RT��y	�^6�a^�>qS{����^L��
����co�V)d�>��.;���Ѿɞ=X�"N�q�	��K�"��p�ٱ�窱	��\;ɔ�.2g�����O=�b<_������5���d���x+L�gr�7���G�z#ܬ�d�ު�'�DUϑc	l�G:��t�tf�ƪ8i�跱9���\�����r��z��ςʖc�ĺ#�@Z�Y-�)����c7ǥ�}�-Z�H��{�_�{�Z<�����W�<:
�M���!�T�U"�^�lC�|���V�j�7���n���,[�RG=��P+��C~�MÍ'�W�d��U�:*�NP����$���m�8O�w`Ǽz!wT;����(��g =�86�S�7�y�MCUs���
�xz
���tD�zu�ρ�������G�U2�I.����L���*f����|q�T��O��ć2BG6e�v}�DM�"�O�{ 2��B��*�����S�C�,Җޟ�'��V���t���.�]��x�ei�O�T�ARZ�4:�;�{�]�W���߯[��T[Y-� R7����\${�5i���"��g�k]B�r��rnN���u�v���ܗ� ���:�3v;g�`�Ñ.�yu|� �����jz�F�/	��@�nVsU�֍zpG����Q�?��� zǮ�^��ߕO�숚ˇ���]�d�t�Ӄ�[Ly6��4�t�L��Ӟ���zIC��}q{��9�>�* ��z��F��>G�*�=���a�ϴ���r�(�5�+�rBա�}�%Ҥ.#UQ���'�鑃W�Ջ�D�p�B9�ڏa�G�n�������Wkў��Xn0�M� �+���
�Y�2�	F���f�~c]�� F�L�k��b���s�EJ���R����.��v4�\�	�~����;���\V�Ik�{�k.�#ی�&���rڐ���pj�b��ѓ;鋍r�2=���OnZ^�Q�>����o����a=���9erx��,�r9/kAYQss�,_�3��FL��2�p��J���,�.�ͬ���g�m�g�#�^�p�����܈�be�T�*fh�����i���Z�����˝�h��k�h�}Oף�������Y��튣q�~�y�g�@K>�������Eߵ_�}!:{���y)l�|k�~�p��W��|�f��EG�~�+*Yznk�cT�s��Yv}�F�TD����]r�r�7ĩ�w�0���5�u���5!c%�ہ�C��v�vm����.��m]�����jsg6��η>��k9�9]K�S���k^N..��H����0p�L��K�����vҞSҥ��L���n�Y�����4j�a��m�}8�gb=�{��}Ϭ\)K;�N�vlyI^���G>����L�����P���T_uCs���{ӼJ!�+�v��a�7�ϧnz��0�}�ˑW�&/�LO��:%�U����td�r�C����9}B�:��5�9�Z��M_�����9�����?U� (���c�n���}[F��s���R�N�Y�5���9k��_�|���֦���C�r\��p$���5L�)͚�����y�q�J��#Ό���9#[��>������CE*����o��wc|v����IF\��%��d��̧^�掾�+�&�}����mG_ٴƇ���C��cT�����<}���X�oޏx��;�h�TyA�5�Q�o�]Hn}�Z��l�ic����d{�d�}�\�����55�f���d�uQ��Mђ��(f�댼�ү�
Ӭ���q`'0,�A����$�����sT������L��
}���7����ۦ�[���ӟ�~7�@��y|ȯM�Q��$&�̱x3�죈;U�.��A�~���j4:s��v��U������˙��ٵ�ś�+�#�w����=թ#���X0wFGMz��\�ts�ř�Q�˪���K��R��&蔳�7���Ƌ��0����f�k�Į�UY͕��P�TOvT��2�P��*����������v�w��P�E1gӘOeT<5�t�Gz�뀀�EM��y3=�xp��������z���ǲ�k��4d?i�}�U2Y��oE!<@v�;�2�W������^7�>�8��9�+ŭ���p�TS]R�|���b�����x��#�+�z��"(��Gܧp�Kӑ��p��x����iF��)�z����q{E'����o��@>Ȫ�u.�(y��:�:~��k���4��9sQGm��SY2c^���z�p�{+�X͘������FT��Xr �^9�1���Y�B{����-�.[(z=�E��zF��]D�������>fΉA�}U���[|�Vr��L����Uo��(8��q��Nי�/k���޽����"�Ш�-��!{��l�T�8po��g�9G^!��/O3��a�����[,�	�� �~��z��S� ��z+3�y�=>#{�����F��l��/O��xiP�u�sf�PG>�8<ߎA
�{�r$0>�^��*�otT!�gD�<� �V������E�����{�3Q��Oܶ@����jbt��=�O��ί ��d�c޶(]JkE���iw�32�Oj�cui�;��'H��f��:�X��w��J�/2��D�TfT�V_���X�3��l*�u���ak옗陜�
�9�Q��쮏^�G�U��<�?~!��bO�{"���܍��Vp~�q�5L	�9{� j>�	.**�,�8y�w����������g_z��B9q�ۏnmo3L�A�2�Dު�>59悕]�^�T�{4�	����^WV0{ٵ�`;��>��������4�t���z7��;7�]�Txms�%[����=�Ay�!��pO&Y�;�N���63P�>ч��|-շ_�J�K>��f��d�?�8�����u�y�^xM�ܧ���s<�D��;����g�W\�}뇄�3�s�i��w��y�_��^��Y�~�=v2S�靦�l�N�{���ۍϓ۟��)��,>Ϫ�	��DUϑc	c������V�/W�/uL��K6<�.�>G�OQc��]>TyU1R��J�u�<�����O����=�9��^�"��V�k��=��k޿dz�D����e�?���Ѓ>��'���J�&Vn� ������c���n(! +��:4�"�/�0���~i��=�����"��Z\I���W)���I1fa���Mͽ�k�� �(wy�N��w�������r��=u���Ѻ�{E��]d6�"��;��e:���gNr�Up_�����j���,9��W�('����_�F}��wG(��`����
�԰g,>5�mO���޿a�%��ɇ�_v��ܾ�x�\�)D{���ː��8���C��9��S�0���9#�N���n���N��@/�t�/Doz�����ex�Mf��;蜺^�nkn���츿<�$j�<�\z��䑱G���}���T5�#�VVa�4���3$�F=�t�����T��S�0�O��ˇ�Y��O�I�8=2�T}�^�Z Mq^�Y�.5/1vd��_YY�#�y��.5��	Vm��F�ʛ���JB}�����p��9����(��B~��x\j�,���;�L�{X���%��wo������w��q���z�f�G�W�M� ����9�;��+�{r�W��և���o���;̓�%�(��yZC�En�"�����5����{ ��=�"~Os/f�\[���jGqϧӃT�fp����L\k��i��wkoٕ��ryMA�5_DŅgk�JVE��[�+��
��5��2<Y�ﵚN�Lu��	�o$4*rѵ�عlb�ܥ�O��Is����F�8�WZ�a�qU�^͋M0�ˋr�8���1��v��]��SV�嬭&CR������:�>!/��SG�l~�����`���V~z�r��3=���L�7�>E�}��5�U���w.���{%-��)�����yU�����Э���.WǕ��S[��y��}�c�	��UY��>�L�^Χ����ף7��{>�z�:�]��V]F�	��@-�i�T�X�^�..���u�ﯥ3q���z��N�8w+û~u%��l��}��ful�M_�S(c����4��dUD�\
��N}YPѫ�P߭#��S9����w�Wg��]����v'W�}	Ғ�Ig�:'��$^L���(w�dl��}���T�li���ww�����x�zgt��%̹0�xO�l�dUa4�x�߉�9������G��=�j�T�<}��n#ޜ���˃Q�$T%�<cٱ�ɉ�մN�^��x������+w�-�L\�n�>�sL�B��ӑ�:}��P�ƠS�^Ed��=�C�"�W�=9B���ʓ�+J���
A���O����9�~=r���.*�����VL��4~�z�'`[WfՁu�*0�'�M�TZ�#��4i8��/>�B+�糽��+<�=��wA3�h��Ya�g,R�_'b���CN��c>�5��vFPδ�)��%d+�����<�"�eQrU����Җ�'���cX�tDwe1�_u�sq�>��S�J�lV�8)m�ʅ}��/�u��ն���v4=���|9
?9C{�!.��y����[\+*Q��`��.�cy^��K�����c��>��$�ն�W)�j�$���{���>�ڿ��� ������`�-�m*{���+�e��Z��TY��vх�����s�R�V^���[IJ�p�P<>�����Z����t� %�R�@�Rri=���x(n�ְz.od�x����y�f]��$��e�KxV��b����*�y�̐V�kT�n�u)��Iv��œ����\��y�om�]W^p�6�\�@�\��l%�n�>��L�[�#f���J]�>"o
%b��%�a�wٻYg:WK�$��M��Fv� ����(��(���{'A|�n�����3�ۭ�H��%X�D�O��iW,��u%�Ѵ�������TX+�;��Kt�8��s�����n��6un[1�c���́n�P�މ�v͔�+9�1�\ﵺ5�W�`+!&�T�{ً"Xk�p&�`�6�Y�����r[۷rY�uԦO+ݤ���Q�Zc��y��w�ynI�zZ,���*�薲�b��N�z���9b�ܪ�b�j]�1$(��Vo)�p��:I��+�}G;������x�iJ�I�s"�R�㯯��2tÐ�t��fAP5�y�%.n�I������.�Ĳt����u�˺JW����n�Β�����iq]hH�w�*=�0:��^�"(�r\��{��E�ĉ7�f��o��=j�M��v5қ�f��!�j[`Rt���O'U���T(K'��l�ff��N�nI�ԕ����w@J���H˼�}!���
&Y+m�L��C0L�PJ9ʄ6�@�J��Ԧ��]��@ovk�M�.���$��+;��;���Q��*Ti�:�gu��s�b	Z�U8�KM�i�8`U2����V��W�J��Y��eP�F�t8`�]W��X=(�K��J�wY9v_BjL�S-۹#G�s]m����ԝ.�M��$�ڣ��5�g3
a�3z��q�"�z1־����!6FL��}0�g��D�Qt�ʼ��K�a���i�xTƘ6�����\�r'�M�O��n>z^��v�Q�v2f�*�Vi�SS;�!Q=�N��վ���z����͈[����U�1d��Kw]�hX����J͗M�4A5��zQ�����5���Ӻ����e��l�r����(�&�æ�k�}� 1���7G���*������+�'�I�Ns-�̼5�]M�+z5�t}Ғ�x�u����$�i�ř[��h��1e\���*�7Q��ko����]j�R���[z�w�E'B�wX�v�u�$�qݱ�H�.\���M.��Fٛ��d[��7:���t�b.�
��iݝ�7v೻v�h3����� ���2���liKL����$1H��őN8��7D�l�u���] �wb�!N]0"wf09sgw(4���'71L���H(I�;.�A��u��Ĳ+���M΍�(���;�Db��B��+���r�끛�Eh�Lc��vc��%"	wk�H�wnc%r�u�I�H��$k���0�������ss�1�����2���&&IM
PE�1�b9;�$;�� �����û��˰�������7](Ww2�@��������I$)�pe�:(���V�+�IDQ{iS�hG�ko:���ʤ��m��yˈ���P��m�:�b� �� J���]U ۵���zJ[�����T��"7v�\f�=���?��e��	UO�Ɵf�^��k=
j�}�i�����U�X��GL�p�y�O���1�>��ѓ������ǉ�,�T{!)�d)��{�*z�[CF��6f�ӧ����e�rN��}�����+~Y������d�]�)�����hS�@���oL�'9�n#}����!�~�BLβ�f�Zc�9���i�LUE��?Wa-k.Ue��}
�{m� J�^��ѽ�e���۔b�{�����'��>Nj$lu �kv�q~�a�W�{�s)��w�!���</T�{�q��v�������6�+B�����(�/U��}a1I\z��7�,/����}ҼZ�׆��\r��ܭ3����fg{��%м�_����r��4�r��!/NB^ۊ��HV9=�}'}���y�^�6�1wst=�}	^,�]�x�E��Ȫ�e�>�C���JQ~��w�pxXN��]�@]�����4|ُC�*B�3�0���@�W���1-���A�UHʉ����������~�1?G-S����t��&B1���mȶ�b���)kx����)��WW]3�孝��AW}5�]��� S;�r`1�B�:4�ݧ[��K�r͛W(권�w�,�y��[������һ��+�bn�5�[h��W9%�Y��'��®��U�˰��O�=L{��̰�ҋ�����w�y��Q�3�<�W�~���PuPk/л�ړ�돣�|����
v��A{^{Հ;��JD�w��%%�\2��Ey��ψ֧Ղb����'���	����	����/��=:g 
��V �'t��љ�f���k'=@t�����C}���[&�����D��*�z��~�=�=����y���^z���)IU���&���ܭ=<'�e�35��=P�T>�=n+�պ%V5[��̋��1��QS��޻��r���L����Uu����}d��Ǽx��:Sj�Yw�A�;􀺕Ət���=7�M��{rp��z��HGn#��܍���˨��'�v���S�Y�4�ޞ7Ԁ�SL�_%��W��vV
���_�z+���>�A֑nfS��k��k��vt÷=G����W�\]K�o��}\ye��<�z���w�M1ּॳ��+��F�9G�2v��3����&o�|6��P�y{�Q�n���;�9�ݳ�¬�M)��+)�%�o�Ƈ%��
�oU���U���\}�I�Ʀ��>"����@��l�7����s�R7}חomV���ֽ[��_-�E�v��s�i�s�7�yS 2�]E��{���]_!�����fuϞ�P��n�}(;��f�^�t�������u�AYV����ι�'�΂�g�Ӟ8��aVZȨ�{��T�<�>�z|��)To��>/� J.^Ss�b���\�.#&Z>޻\lr~Go�bAl�|2���|.9�O�۫W ,�f;=�Y�� �>��'����<8���e3)D�\�Unz��yW��/]�c �H\q^����{/�
c�0Ķl�}��!��^�\'��No�1齠*"ϼS�چ�{��ԑ���PO}@`�[��^��	�E��11���߫���n��=�Ʋ}��!wL�,�Ԭ�Z;�0�W��y��M������P%�:}���z�n*�r#fβs����8'�SrFS�����%��Tz���+�����{��H�����^P�u#b�W��UD4{#՗�ٻDO��i�k�p���W�������yn��(z/�ϯ�鍇>�=,(��{�`[���*z�+"r����z��)l!�2�o�nWo�]{��j!����ߛ�)ȗ43�����;��|�eU�{VX_��M���9�n�sn5��W�v�B+���b�M��q丒�!	������[�q�'p�W1,�c+�L���,pUX�Yb1�r�-\��t�!���P�&��;�{y!M �|���V��W.��n���s7��q�"�,�.�ŉS�e���Zw��9,1�RǵUE�J�E{�#$�4&�w�*Y�8��@��$I���#�C6~�;��xטM��?'�ÿx��S J�W����o�j|'J�ݻtĆlT4"��]ޫ5�ƈ'�z;�K;s�i�u�#/+nNN�i`o���P�*�Y�9�1>O���ͯy�OO�����"�=�G����D�K*�ʌ���2g}1��s��d�o����
2�{wHu]ئ�fP��k���=��n=�W�G{nQ�{:Kg'�Z
Ȫ���%Yb�ɝe�>�~��kwm-Q����jo�:6<���{+�.iTek��a\kF휓�����-t�z�l���m����g�<���b�<�z27ʼ��φ��Wh0�Q���s�ol	��y:�}��O�
^���1M��{&aq����t����x5�Lh��/_�.�ފoY3���U�;7��g���Se���"�[�r���}���v߭��!g�-y��/mܬ���8��A�X�w��A�S��l��
gz�F>F��X^9�>F���u,��l�L�A��Ep�Wjr���rmu'bS�u,��#���u������SV�m�+9�����dmi�o�[�2j�;Z��k�1����,�:iU�c�C��D�*b�J���)k:��2���Cs]9�Z� ��j���1�\r����Ǖ�3��q>l�=��K:�#O��`��T�<�GD��"*���=� �Zt�+*��`��ۚ��A�,�)�ޅ=Nb���S���fA��^$
T%�p|&=��	�����fR�
�.����5���>����τ�e)d�W��[8_�yNDK�[�d ��5UQ���g�eUΝn:ri�%6Lo��l��O���:��Qj�0��h�?H��T3����R3�\,T{���R�YG}\k�M��͇�wv�כ^�Z^�5��UK�����<E��\���=�7_{$���x<�fߢJ9q>��*��7"2p:�/*��ic�gC;o�=WX�7�ƪ+����=�͑�����J7�1���|o��{M�O�Pۈ�u�nF��w:+M��F�f�t�.\�{oށ=� t����KT�ƫܧ�2�����鋅�5�r}#���c*2kK��OW�T����F���W��>�����Bێ� ������t{)��{mg*(�D<B��};���f;(J3��#�܊Q��)BwLa;�ؤ�:�1�ާ�ު~=��k�lp��i���7ϺW�7p
��פ�.���@vh�ÅQ��v"�e�,28�+�kr��1������Y��o����a����w��Z�"�jf���	�"�\�h�G�.wR�5w:�R�M�R4��S��bq�Պm�y���1NJЇB��5�A�/�Z|r��=8숚�o�p�0�g	�^)*����~���~/�=۞t����-P��������YUw���+�����nr(�\�E��7�C~���s���O��#��R��L��,#�u��z���VT���E:�UH�偗)3Y��	�K�'Bs;q��3������l��g����C߆K��91-����U#�^*�yo��[���8����_����>����3�P^�R.r7����y��P��D����P|�E/N�������Qw���5�� {�9���=ŋu�����~`/G���?_� N��ЮIr+h��W�����⤇�r�LLW��N�܁0����Of�p^W��>.� ��]Q����KW���04�1ԁ�uE��k�gѻDz�Vɪ��?���r��U�����-�Չ%���.t�����'�P�=t��S]��,��D䱷���FO��l�&M}��LY�*�8��h�6/9_U�;��W��O�:{�:��r���zr?T�g��뉽w��K�@�G����߲`�0��X�·,��5$B�ܯi:�!sWf-Y����X��+�V�{�Lɽ���CZ�o�5�}�5燀^n�Ck��NiTY��#q�a\�;׀Sef!�iH��s!l�h[�� ���B�9t����n+O�:s���=ݽ��gє��N�G���z\߽46������+
�8�߫�=��=�f����o\�Wᩋ�|���Zn#zX龯 ����{o�5>��ݷ������q碻�Ї��=�����^Uᇽ��BÓ�
���@�\ux�΀�W�������#��� #pq�L
�lY�](��]�}�jQ��}Z4�Ȋ,eDemÿ�g}7��L�>��a\�>�����Tw��s��hͪ>���K��{R���h��%֍L�޸w�:�.2}I��2=�j�R���^�w%�|�R+O���<mڨ�~W>+#�@S7�s�U`O�<���|�}�;w�������=�;��7I��/��G������U��,�_��7��EU��1+e�b�R�ڠ5[���"�%���~�_�5hk��:��P�W�<;���i���w��*���݇U{T�<T�`R�"�������g�P�B�H���M��A��q��4_�T���t]Η�Oy�ג�м�sqd�#+�~��	h�f�?���ľ�x��W�d:���6n�Խ[�#VZ��% �ۻ�c�~~����]���o7�g�o�݌���������d��i��}�c�tџp������I��*�W'��8_)��-]��ҕ>���ɦ;z�]G^���.釲�����[M�S*���n$�U�π����"�2��:>,\A�)���"b�����wN|KÝ�1���#����p��y�r�a�g�zgQ�7�R����[����H|uO��;nHߩ��B��>��ue��t+�;y�K��1l�)�����s�=c�@^�II�8f�v�i~O�czVz�`	KvU;�'��t:�C5M�Z��dgϽC�r=SCiu@��`ңq�#��I�wG���xfp��t��F/|�t�\Fm><�=Lx>��9��%{_�v~������ˁ��4��|}M��ʯE��-�Lx�}*�;p��̘}�Zt?��� �^�M��ڿ
F��{���m�����fU׬y=���O.@X\�Ⱦ�+n窴ޖ�o���	�>�i��9�/gtdϽ����e_���z�������ʞ=�R;�O�pjϪ��ɭ.�ɝ�Ʋ1�1!�y\]�eW>Q��͟U��z�TF*IϨ�f�����,����������|����=F�GTX6n�\o��=5���γ쎙�j��#������q�V�7!�nQ��L��\�.P�r�l'��<r+��.�vYM��e��\��p�G/iD�ȼ��}0��Q֨+F�'S֓2�9-bŤ~��+��8�V�;�\�����\�׶WJB��t�ls������c��h�Yoé���&����?h�W{ٚ�Jm�h�Q��&w��V/{���Х�c	~=�,/t�,(<�z3|����r�,���!���9.�hgU�gf�h���fNw�j./H�Q�0�����:H渟��o������c�����s�o{Dv�5{�{�tQw�G���Ҁ}9FEԷp-K�t���Q}��[e{ܷ�;]��Xc�#�?Ep�����2 ��K�9D6D�w�2:�Uy�X^9�>G�L�x�X��n�O�:N���ʝ�}㨖s�a^��ȫuNJ|'̍�YdM9���NO�9z��m���u�(���#��=�3��.U�>��@w�̃V�Vd��4G��jw-_���rww˫a��|ɍ�����/�`,eB��_7�l������K�_��dO/�p:�2
շ*�^��k��v{�Wp�6���['C��莦4T*�.�]a���˪ǣ��(z9����z�Hנ�x	�oz��*�G/���&��*�������{��Wt�ƪ��\�-m���G=�Vs�w��x	���6o�IG��������'��������Ϣ���v(80�'nA���%]Ə��E֨_L��<µvt͈����yodGoA���u@jX�%&��;���1r�b� `���� x��xZ��}ţ����mr�Xvtʻ�A!G����ק�{��V�C��e����d��֪�
�Y��,P�$*�Y�w����y[�G=3c��(�w��O�������r7k����u�\w�U����R�m���"��N�T%O}01��)�̨��T��k��gU1����{#}5�2V�.�RVkh��R��o�wR=�L?+y~����W>y�v��F.!�|gv;V�{���5���ݤ�UC�_c���n3�wRۍ�[Ө�~���^�c��|���_n0g͡&��P�%F�7��p2���޸x
n|��j�x��;j�t��ɽCܹὢ}�Ǖ_^�����d{�
v]0N}F���Wϓ��,��{p�w8����c���UcsU�V�<>��=Ň��[�=�(�}���>t쪑u.�r��5p����^�C������+�ԇ�{�َ�)�9�0����ǫ ���4�l��P�H�����=�갰%c)$U���}���s>�aT_Wp�ߙcc�Tϧ6g�z�ďz}5������OzD@�W�x���	�R"`�Sㄤwrß�wJ
�����7zE��#�D}�}G�}�Q��m���mk[o���ֶ�Vֵ���[Z����mk[o���ֶ��kZ��Vֵ���km��[Z����mk[o�mk[n�kZ�~j�����j�ֶ��Vֵ���[Z����mk[o��kZ��Vֵ��յ�m��1AY&SYUٴ�Yـ`P��3'� bF����Ԡ"�*A"T�mkTRJ�k-�5���KC�ZТ��։"��mmbJJD��e&�b�B�b���l���^��֨ڲ�&������vѶі�T�s�u�l�l3[l�U����:հ:�ݹ�f���V]MV�λ����A"����*lwh��_s��u�̪2QM)��'G.��]wdP��]����5�QM���:�Cwp��Yjش��]�n�#X���Uݛ���ZJN�&ڪ�j�UEh���j��Rv�f�   ��(骢k�u+kX.�(�k tʐ"�V�a 	��AP�7Z���:ȨQN���҂��UM�ʊ���)#m�RR��  q��o���Xi*̮�uW��B�����<z��QEQ@z4o/^�EPó������{�hѣEQF:����F�(���}��(��(�rڞՅMim�8U�[j��t�|   �K���L���u�L�	h��i��]��(T���z=J=��8u*%E֠iM�E����Z��m��Uk-��T%$�   w�U��m[j.�n��W�ݪ[uѬ�/q\;mj�W�w��z��3Q=:W�
��˶KU4Q�^�mwB���6���P(�l��*C�����m��U6eZ��:�   {w����ۭ��zr���&�ݞ������q�ͻ�[kj�ٻY����P�=��ج���:VkZ�+XCCV��7�޼�a@kzөVh��m:�����l�	QR*�;��  ���Z%5�f��p)U���n��g��m1l֑��12�=�.�J=u����WV[iZ�v�-ov�Z𺫶^�N�̍�"���wz�Y�Zm���'MC��U_  ���W}wwn��])��.ʇ�F����� :3E�����t�j�նX���HÍ�-T�[���� �h&�ut�ZoC�ԝ�P��uuY��h�  ��0�2���=p��m)�ïyO]5@ԭ����wGMV�ק���i3w7��[/YՖ�)�jUҶ�wJ���֕뫛4�]w`4L�RleUi��¡{�u�Y�  1���(��#���0ҁI�\�PW��v�z��f:�����K�SY��w��)v�\��8]�;�כ���j���v���l��D��-�Z��iM%��  ��إ6_}�Jz�ֻ�g�e��F.5�U��/j�ً��͝#l�mr���vi@m{uT�n�7م^{.���؟ D�*QP�L��O��JR�  E7�LU*���  O��T4 5O�4J�h&F@	4��U� ����Q�L�����ys�7���F���b�2ˏ|��~��������2B�����$��		����$��B���$�$ ������y��O�3��������MKX�X�/��kj�ի7PÅ�["v7l�):��R'2�c�� 'MV�D��鑳!yn�ӎ9��b(f!���/��7]8��L�Rǲ���o&=4��h��J]��=w�oe[ MŐP��?\��X��Q0���:Gsf���- �p-4�
Ż���.��7�2*A1�i�E�fcx�ȫ[
Ȳ�di��&��E��nVҦen�yI��d^�Ho)���0lIT�X�PXUa���3j���QPED�s/�i�M"���Y�v�^�C��(#[�p컲M�`MQ��G�iπ���ܔJ̷d����u���n��f��j[_:���- kvf!LZ>��H�������h�N^l�sd[6
�[��m1n��Ф�+ۭ6��z�W�0��1�q��)#���!��;H�6�f�!�7Yd���kT��j����k^�f���6bFA��!!ލt^Y�*��Q��,���F�S�'D��V��VT�vIg0`��)���3t�3n!*9�Y���7y(f�Sb)n�o4�[�
Z��Z
5�l��ZpSj�nX�`�}i �RGor��3W�a�fi7N㳍�q��-�X� w�[��=(����V�4�J�ЦXV��ܚ�p�a��ƫX��-Ӷ�?Y���=���M��q�&��:(U�V8�4��l�i�dP�8���N��L�.[xKV�2Գq���@�����X�Ȩ'J�!m9f��S�X)}����)����2Q��>��1a;��An��2;�����^Z�i�6�ˆ�.��՗v�hߓ�Բ��/.�R0��$�/i\-�qݴ0��/���/�w�������4�U��-�[{��!C-T�a�4Y���w�4����GŲ��&d%ꤶ��l��e`����Cp0��͗%ź-;���/S� dYjV��'áQ��oop�*�P�3�h�%���B+Z��3r�A:r�w��QDͭձ�PG� �J��n��ucRJ�V+ܰ�:���TP�n����-a9�z�E-n��#wnMI�څ��qe.e��h��ᳪ���{��V���շm���p�@a�N��3�b�l���xY�eqn�����2�!�ݭ����4�ki*[2X�ks4�V��*A�jc�2��R\.�W/2ֽ҃�_ʳ�h��-�56Р�"��z�������ݑ�"���"��yE��)al�P���/��.�	��OR%����׋F�M+9��b�@#�d8T����P����+2^ NU��
�M�e��އ���r�**Fu"�Ӣ%�a̶)�	��"��oJ!
O8r�t�φ�L�4�E,Y�ʗ�E�HLoA,Az(��x��;�zh|?%L�*3����!�	��쫖L�Nܵ�=�-��y%�p��T�	��^�xm:�ܙwij42�P�%Ie��0=ť#�r�V�|��6�)I%����L�ѫ��w5��q��%��!��ʹL�n�9���7��Rk1�:�CVE�� M-k߆[��\z]��T4��'�T�Ӗ
	et8���F�Rn�eD�	�H(UV��+d����F�H��kK���Ѳ��Z�j�SZ8��Z�;̠N��f��b�����X(��pN�q"���D�ޡa*VwRt�sh�[�$Zb�� éQ�f����iġ�I��Kj���Z��s��Ȳ�NZ������]jhf�GF�J����/T��)gJF<ӫ^��Q��	�A�X�+��E՘(D��ͥD����+j,w���12���D�*�\sB��)�#&'h�s6�7��بD���6��O맇V;'�V�^#�.�s嗎I+7a��A�����V�a�vP�B�Z�J���{y�e��j�6��Х��TmX��	VQ�ό�t]�Kѕ����	��Q���evѩ�S+^�u�� ժ�V�2��ځ�cƓ�Y$+F̫ŰL�WX�!X�1���A������ �M ��u��EQJ	n����v[�Ho[�4<2�D����R�C�����K���;���38�Y���.\R9��)�,�L�Um�pn4U��P�*%)G���ŭ���U��խ����ODKq:д��~`S�G�Jw���խ���ϣ���Y��V�hQٰ����2����eJ)��v�8���-��`����̢��H�T]���;�����n�܄�e�ۗd=R?��R�XTP;�-��Hnى�J��{d����v0�p-��%m���ޚV#��v�J8�╖Q�f�t$����ܻ�8Z�����8�Ԑ��6��,L�J	���.�:x-nPa�1���YD��Zౘݚ+)�e:�4*��̒�ʨ�\;Dm�-�f�X��4#��ct�Yٸ����9G^f�b��1f@`�C�!���SEnYXa-�y�u"��Tƛ�eh���1V�<�Z!�))R�JFe$ݴ�j�+m��N�c��V#[p[��v�֑r�KJ/��Ħ�謳%�T�{����y�ӑ^�T*1���Ir�+7[��5P��1dؓ�SLyKksF��S�6�&�Vl�Z JkY�'�]µ�9��n&�;Ge-�J�sk@�<�n�BV���d�G"��z�%	�ئ�I&�M���o�Rqȍ`C`SV6�Ӣ�e��̒E�֐n�
)�e	�W��J�V���V��U���dڙ�����˺p�/C��ie��[;�&K�1u��0��Rr����`^���6�G5���E��VT�]-��)ۛ���iҸ���I���4��ű�+:�J�d�q��ņ;i�!
A�<�6HY��&�N�lSM��ڙ�bȝ��Y/a�A-��*�t�H^EL�iOZy8i��ҤM�}4q(!\��J��n������j�#t�]!Wy�s)�xQ�ֶ۬	�ϵf�m�o�l���"Vj�E,��y��I���
�#j�VքY�.�Q�b�O�ɋwV�����y
dh��v�����I��A3!j�8�KrT�Z�Ϯ-'L�����X�V�1�%%�����1%��5��Ьc�ډ��-*�2��"�:*b���Z���Z�5������eَ-�֩�Px�ɖ�/r�R��X�onb*Gu7J�3m�RJd�h�U����^�j�e�3i��7�&E�����
X�bVR1���Ŕ!�$ҺT��vAZ�J�2���#^�ʭ� �/VZ�ÍbۛZ5�W)�׎�\r��!�[���j;WGr!��K��dS�ߣBʔJ�\2UhJ[�t�[��+Ԗ��bᎠ�R%���S�l�IZr��28�!���n�Nk���bK�qB�Xe�̫�3r1��Be-F�!6����,�V���{����sM�1�ڀ��
a��b3t��,S4i嫦ue��@�KMi�b���մ���JR5"�:��+j홸�� �'y{�AX3lhz����W�ܩ4���٫^��0�&�Vf�-kڲ�^�mFP�Z���-Rh5�t�e�Y���a�N]^�Ur^2�ֶ�q���U� ��0�	Qi]����.VEun'+1�@Y�/Y���n�3m4�"�m֏�[qj��K�:��낦L4��;���k%0�[��>	!1�YB��X3]�$�X�d@��Oh]���*����S��n!�S�g&6l��l[m�I,[�ꃕ�S6k)��H��{��ȴ�򋒳b:Mb/NV�y��\�n������Rd=�-B�@.��kI Өp�����)p@C��.��e���]�^kxS�sg��aZ�Y(c�6�5µnFd�a\�cAQ�w�g$L���=,lj�eh�˒�r��O�^�dU�c�k�q�&^hi`jRܦMf��e�&��� �^+� �g^-��=���U�`�ڌRua�n)�f�t;T�e<Ӕ����f���:��rYʃD�H���t0dbJ�-æY4	w���r��m4qj������I6�V�k��Т4�n�x
�ċ-�8�VG�,8�^�uː�Wݓ�y>fn���n�F*�U�#��-C�)k*�b!#�ad8.�6*#/@����IՐ�١s粬;�7υ��ot�3"��O-���L\��<4ӕn�asi��[+^e]����T�%(�aH�I�݉,�-e,�i��^ah[ן
�Y�.��@T�r�1�xVl���	}Aj�(ʂ85��c���G��/~�[`�G������Z
o&
�Ӓ��a�hPV���c��+wY�Ѡ���C2MFQ�K0}�l�� 6��,�XU�Ȥn-�rH��� �(B�R�l��:�u��m�B����Y���aͣV�Q�Ou����+(���ӗ��
�p���N�W��Cl�v��KYu�V[SwS�4�d�.��G���d\�͍l�-�3T�pҨ[Ne����r[E�c��dۄ��pa�ڸ���&ln��V4z��:$6��q�eȹv�R�U�����\�n
eD��ֵ��-�8T̰��cp����(�5�M���l��+�\���{�����
s�w݅��ʎ����';F6i��r����o��sd�<�6+t�O
Q�eVn�x��h�)�-����w�P3H�k��B�+�Ej�*Y�Pcoe1:"����K�ܗ�Ζo�J٩�s�Kq��/��z&��[Y+0;.D�{�m���#�V��%��AZ�`)x4q�Ң��;�Q�����V���ڸ�7�V\�: ���n�؜�6�Yq�v��J�\ypfE�(�B 4���ڦ%-([6,b�8�R�h*=�.x�C5�nK�+6���5#߉Z�WJT�
����t.�6��wyH(7D�m��f|u�+�5�� ��F,�W�p�©bf-Q<HIy��Pݟ�+{���N�O�AP�6�; ֓32�Y�yv��,��y2��Ӣ�X��E��y��=��h/.��>*�rn&'X�n�UeL���"áK�o�{
xt[�eI ,�Wz��s*�#ݴ͙���t[�f�k��U2�&<�b�ױ���X�7�m<ǌٺ.�"�sY�^��^�T������*u5S�rb��1�E�J֡#�V)��#C	��f�%=av��x��E8""mXf���N"��P�f�di�s|]�y���Ǵ��%Ѥ�n-������VP�ܪ���8!:��9Qn����hJ��VS!��@���.�oh�5�X�9�]�~.�ЫA�W-�*J���[��!aSb*ܶ%m"5��lEF��r�׺���G���2����wD��4j���.�/i��n!f�����W��Pĩ����k-T����-S���Cd� LUx�%!���$`�]��++c�ܤV�X�U�.��V�M�����1fG�j���=�L�Ĵ���:�f�{�X*��$X��3M5e�ܫ�-�1e1��r��7�@��"N���
��7��3�â�]<�iE3K��ݴ*a�W+7%i���ַ��њv��135 �7�VE�/*t�[�7^�U5��5�)��	�=�����0F�cr[�p�WSi�,��1ZxqP�+X��E% �2�wK��oFT��j���)9#��B��FSa+E��s��L�CR�ͤ�v��ح�*�5�i�Rn�*%ɣ*j�ͨmioQ)�E�jR���&�gq`w4�c�^���c�ѩ˔�(ݑYtt!W�E,u3�eBu4k]��аK�����Ê���Fkq���2mo֮��T:F�E���f3R�C#��S�Hi8G��DcyDb4
�����z�ÊG�0u�>���u>��/%e%��2�\ܥ%k�d�5+6��eiJ��win&�gU��Q�[N���LѩA��LQ�m�7���FN]J�0�j[���j�5%X��s(]ٚoL�Y�5鲅n!�ޠ�9ѡb�cZ���%��lⱅ]7\��$�h���\u2f�/eL��R-(U������å��[�ɇe�8A�����ҭN�K�u�f.��ĳ\I���;G7y[�B@�]6�;( 0ɪb��J{b� �c��#9�M�)nAN&�`�%Q;5q�wC�pw*nKM����6j#�ݛp��;a3l�c�vС�SkkS��%�BeGJ��Oƈgm�f�R�5]�̷{�Qxj�ە6}��-�t���MT�ʗ�h�;��hǵ[�!���%�n�.
C^ �1����Qc�8`�����������8e'��!v�[c3k014\���3i��[{�P�ƃ�����1+x����4Y�m��[�+�.]�	���/Q!6�U�*��w*؋�r�c���g,��X��{�*��7�����(����XE�T�"��Y�*	K*�s)��k�M�l��D�ȓњZŔ��WP�by!�$�*��w��R"��R��kn�kS��[�n��ٌ���)�7
����gj�K"n�W�i&,ۀJ�J�n^�!����ѪIC樼�[X�t�x�IM͒O��[�Ǌ3�F�RV)s ق��f�;���ܭ�i5B�8.ZR^��3k`pk��.��6�&�!��/)9j��X4S����YyyJS.0��iL�sI�UR� i�����'N�Y�R��v�2�?
yV�*a�F
�F[zħ����e��(F>��ɠØ�ԬŤcO#�m�V�,�G������3��OV)ZB!�q��li�,�%��?�G�q5�ٽ:9�u��Э�܄�QLV"�w�Lr�.�N���J������w�NʚZi�z�j����M�
�Y<�]nR(�-!Q	�2`�r�������=X��!��_˔���|_qfW8�T��{k7�aew�r�؊�(@Y�a�[ٶ��a��v��W���e��o�Ѷ�٨����i�T�g0�1�ݙ�L¶�.�������L�x(:��a�����u`����y��eڽA�5��n��^�r�9<�=��qA��^�=ET��Si.�κ�f��Jp�I��cʳ[l��V)��m���9Gے��Q�l��̢��y3:�ܜR�q��9�F���5�Ki�:m"�I�s�"�7vY�
������'j�_]�|#�`��[M�&�!K���^k���;�jҊpO:f�����I��fp�YX�>�U��ꊦ�f�e�`�GTr�� Cn�Hda����T�|�VT`)��)\�N��!�;_ܶwX����Ur58������}��t>)��kǐ\��@
� ��-rn�X&�=|���ckkMo���Z��d�F�+6��p�ۧ	6�3v��^<�����0���'Z;]°
NC�M�w{mA�m����*A]\��Ԫ)f\��+�Tޙ���V�8[:ڝ�����P��}Z�w+~�}�j�E�hovb�]Y�|/0�N]é�8�6���ˡl�8Q������;Zb� 7��ћG�H^$�*��v����u��߀U��α�{<q���v1�i�¹�Ȳ��E�����:��w`T(��n�cb�j����ޱ�����S���IxR�)0��ҡ�9���p�?M��QB`y�}!)��ԙ�/Fu�����,�������	;�W=>�F�`������rЇ�Җ�mp�(�޺1l�޾ɃJ�H���VE���Hoj;��ƙ�n#̮2m�4����,M��{��Sܒ�mvJ����w��:�V�i�f��Ǌ�N�-_V����šL�k *�r���t��)n*c�x�n>X5%5)Fy	���#����%�z�Y9��I1����J����e�ߎQ��6�vF��ܔ�ϙ�j<���obXҏ��%G�4$i��N�)y���NR���8ޣ��4��n�ܳ����x#�9����B�"��4�\g��\3U'��(�M��Τӷ�b:��S=t����L +��:�z���D���kY��YR�T����h1�*��B�w-�t���^��0�E�1�c�]	�
M���2�_p�rY�ύ��vz:�ރ8�TF��sXQ�k^�ݡr��Ra�1s{ont�(��[�^':{V�����v.ʗqs+Q�ǜ�VsjnX:��hSo7,k�V���L�P�����U.����6[�;<'�_>�j�Ÿc9f��D���:�����a�yC$�j���¾}�(j�\��ܒ�w���	��FŔU�e;�[��u�G�����E��P���T@�{����j���kt&�Q��m�B���K;3D�nl���ȯ�4�]v;ZmiQ�k$�t�n�����s�g{*���+�G�q*o]�������򌼋o�s��%�k0_|#f�ò��w�:nZd:2�s�Ywo���d�Y]a�M�{���n��{����|1=L�N�[Kne:�"�{��T��X�]u1�c��z&Աӧ$�˚���A�7�#sEζ�W� HV����Fc��+�����0'B��rs��=35�ľ�q��wHT�)
�憊U�Z���	ȅkg�Y �R�2���7s�縉2�'k\��/b1ֻ�S�WO��đ�x���M��s�|XNպ�Y[�b�+0�.����h�.��+��ʰ���E9_���gs�}�0��3��!�DE��#��eSd]:�ƨ�,Q�X��7��Sћm��9���~�v�N{�h7�\�1��p�ڵn�rnr�;����ԭ��x����\3hL(��l�fTl�l[�d��f��C�nU�wvqF#p�8���3��F��"��b�g�`��c3o�z�}o�׌Թ�zZ�8���$N]�� �u�h�v@sD�hٝ�:�i]�5+*3�M3G�%,W�:���K�	�E�BJ�G�o �O���>2k��L5��Xv�S��ąu��w�*9��{0V&nS��Z�P�Th�s�h���>�.���w��1c��5�TB����k��!��V����AWF厾��}^v>[��Fb
f$�ce>t��F]����ۻ@��V���8�Q;�0fQ�*��%p�����j����.I��v)�@�X�Y�,[2rX��ݍK�)]:�Vk�Ƃ��8jk��o1GpY��N����wB^�kE�"Z��i���:6�2Ś�JA���e�� �b������Ud]E	�J�[���Eu9�ƭt���ޜ�n+���S��+���P�6�6OK�>J�OEM��1���=���x�5<|kG����d��C��C&nP��U�뱍��륇[���������Z][m;쮛p�H
��U���
�wE�|�O�l���o����XD�K���W�1>[Ҙ�z����λ[����kY.PA�}��>Ȉ�]J�ʔG�OH�W'������F`*WL��(����Z�V��g���B�5��hW^W��E�;�4�7z��Y�IE���L������/,cU{`t�%Qut�O:��A])�Ֆ��G&�B>-�	�.\��>��}�1a&�t<��չ�b㣙��1���hj�8��o���ܻbz`�+SS,-���L��	(�:�Uw+�$��k���X@�`�X��߈�ޡ�L��O���Ło��;�z�+�%Ȳ|���r������i�Փ��g^�4+����RgW)s�	b�j��˞��D��3��<Lǣ5���Rӂ���O����
�ʔI��vég^7;�]�������&��7�`�Μ�[o0:E�oJ^�L:�tНIµ���h�Z�W)����B��%}B�7ټ2�<��m��*۴1`�)��\��D[5�ѡ�K�w!�	S#7��
Wt��{׺밐�{:r{g�4��{ ��D�Vϟ^-\]q,h�[������ݷ�+-�.��(At:;!��(L�a��Ĺ�WU�\#��k��Fd�	�R�n�vX/�+xc��Ws
l����$3ub��v&��7ia��j
�}}.�I��P*�r.����T-fL2(6�³�*��R����`��)��-,�˚�_�:c�vb��9�\�Y��L��m� 憯i;]��8�m�:%����Ww���|��֠���?r��uڀ�iE�R�E���+���y�݋#��t�\�m�$]۔E�^�ί[bS��=�����ܰxc�)E=�9r���k�p��)G<}���k�X �e����Gڪ.kOT�Y܌͏��d��r`�&�*j��^f��	�D�nhTI��4�j����P�Z�Ss�S�{�'�-�_*��TH��#^t�a�5m�*�u�������jJD�V�ҽ "wV޻²��m����)fCi��n1�X*̓ݐ�͒�5I���l�G9�������c��<�-`�����Hn��QK�1_*|E2����v�79�u3�y����"څ�����;����:���;sμƎ&櫈__j�PB_:(lS�J������WWn8�q&���s�\M�X�6�o�Ał��@޳bG��>J���ܲ�*�wd*�2��*�Q�/A�*�Jn�������l.K�!Ӓ�J�<��s��C��i���R����p趰<J�D��z�j�_X8[�oŖ|��A�Z�-�z��ٯk���7VN[G���L|R�����=5�'���w��n9_b/������Tc�|̷��+x7Kν��5���YW�:���Cv��j`��vˮ8,��,�[)B:h�R�<z�ʊ�	i���9����ċ��s����;�r�-�<��N�\�d�����ɱ^S�]d7�����W��c$����
U��{�=�7�\�d��Z뜻t,�1Kɴ(�}g.C��d�7�	r��tJ�a�&�jw�k�ղ��p�)a�m[�Klj���b7��x�c�KvK@����#N	��E�X������iQ#�Wa�`��[��N��m���[;)5�:�g�N��^¬\*<'h��/K�]�YX�"�'*���]�u��jק�R��k�p�ftͺ�W`Z��<<�S��y;b��lr�c��! -���иH�~M���=A��Í9C���� ��{Y"��p�[{�����(��1	������*��;��q%�XX�B�f�=�G�I��k�Ӌ��=y��Cb�b��$��]t1*z�$��U�*"4���^��;s�ت�-������u�u���P��e��5��td�L�#�#ifV��:�3������GE�NH��z	9���x�b��w�O��(i�E����Η]~n�fkFXu�:3�(�Պf�6wx�qU�
�/�'�T��\�Rk5]k<�NEdosu|~��vnAQ�|�9a�UD..�)'�]�.G�Z�<��p{�Eg:v�m*ľꊓ�~���q���r�)x�iyG���{��L,�\�l_d'h��� �/�vQt�tU<=�i�7���Xf�FΆ�m2ݺ|�ݥ��5kx9gF֡A���{z�#��%t�hLCFHm�V����jԋ�y�*�b�w��M��}8,�&n=uy�dǺM��N���e�y�e^we��5�Y;U����WL�5	�{����-�:�����"��[%��tˬ7����zqU�m���t�쳶B�µ��{��e��K�Ii��<��wԏn8p�7Ԥ@�q�Y�'gn
w��z�
�s�LsMm�O�}g�
���Qh���A��X�ǖ���va��7ij�X���r��S����1J�uu՜8w9ڤ�ń�ih���ٖ�N�/�b��L���Q�+'is�z��Ֆ��g'z�������W
.�Cv��q�;�v< ���a؈^�ڶo@Ҹè�T��H��7�M�»�D�fLD`ޒ5b9�4	4���U�rY��EfU��D���ч������>录���k��gml�[p�[|���8�k�	��d�U�)<OpS��w6�#��ޣ"��X`�_t��G_ל��ǲl�e[I���m����͋ka�ڄn^�c#���r,x-Cڷ���[y),�����4R��[=rRt���o��in����X��[Z�Y��犬��'Y;	�Y�MW�'R��}\x���7�plrk�[q� .ˀ�7%�;�����1��^ho�瓜��lL�=��7ӊ��v�_N����e0)��eݕSNm�G8�\����Z>����n��4Ql�;KTl�2��]`��m�$���v���K����j�X)�Z���q�#��H��ۭ�WL�(u�yU�ϫ2T�7>�#�e������n�v�Fqk2j0�-���%U���7J⻫s��3�.ao���_kd��m�Nʹ��wy
nS�+T�E����w�W\�%��9E԰B�^�tCA�.�'r����i�N8��&��Q�z�GEF�u��(5T�z܂fy�3��S�>�Tχ���p�Hn;;����������i���R�гxx��	\\�b�yu|λ�7[��ekM��E�3��[�R�TS�*<M���X��ռ૶þ��+4�����]ZɣP}���r6� >�:�F/�_-�I@��d�0�p�--�o~�ɰ��I��"]�	kw]_SokF�ܚGWes �v6u��N���i�Bf4�d��z~��J�������}bm���.�Ʋn���-0�7Bˈ�q���{�@gV����s��T.���F��0�P,�ۯY]���dKC�Z��ŴՓT�=�{zk9��#���#{+�T��D43kpJ|���f�溴��\-�U��R�Xq9��T� ���߀4���� �@GӢ�����ٻ��dW�%���f����-_r
_`#W{]�v�l�oRϻw-��m�zp����a��w��u.r�`X]�]1C�0��|k*��f�e����J�#F����K��)����b��u5K�Ts���9�m3.���s��B���$�#�{��j}T ؕ�ǝ}ۓ�&+"�z2Mb�,,�OwV뮥;�P���T�`��r�t�3=�8��C�g
�g���}�I.�9 �2�b5��+��a��e%羣 ѿ�w����5�a��쒌lM�iq�D�F]	}zNK]qS�e5����]��;პ:���zK��|Ί9Q �xi�]�OƲa���o��M*6��ޔ5�Op��B�e��t�V������7y��(p�6N@Nc�|���I'F����FU�-|J�5]Xz���0٣l�k@6��K��9ddU{�,�=탶�ȸ����yrW�U�ʷ���}�,�b�R� V�X�P�͡�E���m�W>�N�$�q��9[�5Ҷ�p���eՠ�6�3HVg���B��׹1-o�sk��b�Ȯ�b�%^��!$� �	/���oC(��u�ޗ�AVq��5�+��`�nd�e�ښ�T�s�҆Gs��@�G7^��O�3�FFi
y�	�B����peU���􃯓�J�P���r��Y���ynJ�	�>m��vm�.��&�~k��v�&����&p��mw^.�'w�۷�9m��>�v��G�wNѝ�GZ��F�W�<�϶9�����		�H@�y����U�+����Iʵ��T��%��V�kn��J�k{��2�̠O2�0u*6�)>�j�o+aY��o��2�!S���X�\�3�
���nv��[O�"���ؕ3[�V��f[e$�Ugw9�.>U�:�ݕt�BJ\�V5[/U7�+k�e0��޵n�C�������'}��GD���WZa�z�C�R�X~J�L�^8�70��ru�S�x�������uUׅN��؂�8I�\�e]��l����Wm��V��5�;u��pN�[:Ao7dX��6xZ�����_&�p�F�nw�ՠk��s�w��X�ī֜�g�٬&�!k��l�'�[ξQaO�ި+K�er�l�Gƭ��ΐ�Y7�
�viˊ��� �P�鷧ǅ�Q������q�nP��rg*j1/r�q�HW���{�9l�����Y�c� Ui�[�V�=YW�(@|�Nl��Z�M� �������Z'V�:
[R�Z�RkN�5)f7oQ�C#o-���c6����n�aŶe����2����a��Jt(j�6��6��F遵z�����Ԗd*�c����6d�h䴬ʟ��]�̲5]�_:�I]�]!x:�D���1&�*R�]���1pȟ
WqN��z�e$����-#J�6h����$�٩�d���=��ً.&E޻�%f�dӡ�[�S�Y��B��M�VK�:�=�c�Y �z��J^hJꝛ5m�|�>Q��D+��V�u��Fuչ��FĀ�}��o\.X�~t�P���s)<.j;�\o*�i[�3^��e�yϴ�Xi�kR�0�Q�`�.j�o6]�y�#{�#-�yf�yՉݫ��*;�6>��N�b��'�	�e��Ol�Hh>�pK6J���&�#�>$}�H�l1�7}{�z�K����J����@iW�������� �����n�g<1�Z����Jӡs�B�e�8y�;���"�*�Z7�cy\�9�ST�	˯$æf�FŻEC�7j� 4hlc��\��k�1j�sŷ�v�6��s����M]��c7�˹�#��m4��6��A�k��%fԎ��1�v�["T�N����hV<1ءΕ�SB����}���}1s�OQ���(*�qe�B�K5��6���ۮ�!*)�v�Yt�-�*�t�k<��M���5�"����5�'��v-�j�C��&$�a�Kɏ/��8нN𷛓r���X.r��*i !0�6q	x0��Ku>˫n	{;7F��&�3Iff���1b�ݘr(��ט4�+IK.����h����v��:t��0��C�
��\e�CM>fS�(�.��s��&�a6ݑR����q�+x���]ʻ�7)y<���Ր�˻"��1���a�%C�.�6���q�U��P�ʀ���HtD ��k���̠n���u���^NA�΂�.EG��Ѯ��:�R��mʋ�������g�,���eb���|�XnPl��˷�]�r�M[���պ�E����z|�X�� v��,L.�t�M�Ej:
�������v�Lp����v�s:�l�)���K!�H8��v^	�i�muͺ)��}/ShX���]���+v{d7��z�>��yl��+�sO�ڼ��uu)�|*�f<�n�yK�1��J�.�}y����R9���K^{#Wӣj��NJ�)�B�ȺI��˵�}v�����د1��wB�1����+$5p@����n�u=�6ې�i����;L�͐X&�ȸ�IJ�+S3�}��]��|��Uv�����U�I�%��}�{n�"���=c��]�#U��^��+ǥ�]�t9c�D�u�$4��Z"KeY�g+�\I�O4l4�
P�u�2��t�Wwk���J�Ь�� ���X"�/��$�VtE��k4 ��'[oI�g��f�˗:�Ё�-�[i+��R�hfV'�C7�lr����P[�Y}��KF�+��Nx�F�^[��(��vR��c��|�Wn�9�QQv�xU��H���R�i^�Z�t!����e�{ϫ5��YWp憚�-�2��w���P���e������-�$o��i��W^�(kT������)֊��Б�g4�2:�@����S�X�k	�}!��J��Z�R��b�ݣr��,n&յE�]�U�J�L=���i3\���}��۬�`]�7
��6��Qq�E�am�'Q�G�����e��_i�>Q�{L���D�	����+g-.���o1r��^T��g�<��zn�����(ۨA�Σ�9��
�
�O
�[xJs�Kz;׼f=WHR�r��̾	���F[}r�!mԜ,��͗қ�c/�*V��s^Nđ�t�v���b��M7��l�8�Etx�Q複�\��\�x��v����P�1�&��ջ�kË��z�&��y��y���Yg]<&K�a�6�4qhkw)�����8��@�I�f�{����f���Xja�OO���Y�fu�a��[Pj��5��
�Ow'�]�!�e��>����#Z�EL��y������=FNg���.]�is-*غ{���RO,�5��rɛ1p�"[}�����%��&,���ak��v��t�6���X�=W�P��ֲ��|�n�)�,�wu.W��]�P�U7��+����NoK)m+;)�(Q�∾�Z&���:�����N�$)�q��������0�z�AYj�_r�E l&;]�K�z�3:��"���Jen�b� �o��O#�.f�@�F�a�^��Y\��tyvS���,�:+�[����L;}�R��QYF�����{N�f��P��;z�Ն�A�.C��}�����:�Sͩy#�L�^�3��HD'wh�u@�^֊3I\���@�V��;�RZFO��F���N�̔ŭ�=q��3��U:�,ށL3le&33--�澋��J���m��	���� ���8��\]u�-c�wt�U n����n�pT�m�F�P�0]E
x�'/������v�`ܻu�:ё$�B�)�gD�,D\�ެ�*c�V�`t�r����[���⚭2\��U�g�m��Y�k\�/4��X�����y�ܖ�/_Z��ޮz���&�kv�ѬK(���K��Mm�\�g,�>�d�urԚ��օ�b�J��(�bt����_[וـ�&�i�nY�R�F��.z&�to~5��´T=f�2J#9��:C6�L����l�K�Y����I�f����Ň�t���x�z�ͺB%����r
���K-��7��g �Ɵ�o�5z���"d�dj���ɨ��)�E�?�:�T�gJ�ފ��'NT��gQ��ҟ�.�rD�U�Y����-��Z�nL�`ȳ���-٫?k����FH����mVE���%�{�Ty�;���61�q�U�`�/������;Zg7;��j�T_r�鍙�T���u�}�4�e�Kv��1�aݵx
��Sɲ�ޔ��50*t;���L�})aS�I؅�Ek��eմ��E�d��z��\��I�1{|�Z�ѝW��c��H�XwT��}OJܶ5�1B3�֋C9i�`�Bt�H��&�j�nC��2��%�vަ��Ubu;r\T�T��<�B$挩:�*`��\�(�H1o(�{7s3��7H��&hД��ܷEЭw�I�u����sPky�p�rYleq�#��r:E�l�N1`k犷��{��媙��E�ε��Sژ��|p��XにvVӵ��h۱t	cZ���|E:N�S��܈��(vST��Gp�5k��NO6�D� ΘcJ���r��nW���R�N�4+/�p�1� B��+o�Un�`A��W%�b�В�CQ�{�+vVm���7�ue��Zւ�W��,=����r�Z:�{��)S�h�|�s��N˸�e���<�z�Y4W:����������-�o�*3��)8ޤ�R��e�&�f�����v��H�8��]��%:*H��[ֵ;�w@[�X�ǡ_X�3��)B ��v�N��/V��%G�#N�\ڡ���Ȃ�Gc�l�#f��K)��PW���^��ݔ�=�+�V�U�\�A.-�a�f��i�����F3�.��R��Z�'Sf�o%����nC�)� Ù�ue�\���9��/%��S< ƍ�Y�=V���7@q��A�E����ʵ��`C�v���8��GP؜+n��w��m�����:��/������Pm��rW�-�V(�ف��Ʊ�w��dVQ��1M��a;��X6�R��z�n�� �]� 8;KM��;��|�W����[a���<1��'o��Dfrϯ@�	)����;Žg�b�9��=�$U��sɧc멘�v%Xj���v���)*yi�8�T�!�4:��*��a���A�y�f�ʻ{w	N@�q��Jf�M-��C�,�����\�$ys���:���j��I��z�dʘ� �X�7v�{��>b�+�J*�ꐰ��]r����9m޲o���S:-n�R�5�R�;�)�g�JH>�! Vi�����k�me��P�A�FԨ)����	�&�H���8Ɠymxg4U�w�`��bLFu!�$D���� ���1X@85c�ŭ��0+������oa�sd�j�s�oTV![�;Q�c�h�ywQ�&��&��igYMh��:'�0v��G)ސ���;�{)�1�H���we1����K`;t�2t��ls=V�ZQ��T��I�6G�<�Hg�QQ�x���K`�]��n[���� NlԕZWQ��S$XWvvs���P�Kf��̓y�Sb0-�X77�|�}=Ś�\��wa��������2����N=���>f�����K�L�ν���%�S�o��6����,0����%�U��W�#�n]��[/��8��3�5��n��ML����O�gθ��[wؑ��r�r=�i�e'����@�
�­c0�B�ha\0�Y�.����a����
u{k(�)v"�l��j�TXg�e�����Ϧ�yu��m�_n.V�۩/�b��X�g�8�.�K���]��r���\�m:V ��4ś�Z��}��ͺ�mnF ��NK����k)��|^ecRI�6��yw�hU���_5Xf�W;�;��cv���P \x�rR�^ǚǼ�\ڜ���qzm�z����8@��F���'Or��VRp�v���e�Փ��b��F���:���5���`$[�*��<��z��q�����M+�
����Ǜ�x⻌�l:���]\�K�{V��(�R鴴�~iv*��w��4�U�"e�q6�a�*���>n�N��MSt�mNe�)���~k۠F6ps���#�'h�v�V�;H:WF���W}�%�����LU��N#��N�JD_VZ��\��
��\�Vp��Cn���8�O, `=��&��uj�B��K�����\���+b��0�x.���aR<6�`��f}`�t񺰲�; ���*PuX���D:��bł����-P>5�}�lJ����ol��9v��[�WWpf���J�͜��
����%;6�3z�emb#U>���[��
�J՗`�غ��\���ݗLҌ�Ӽ�[�eE@����`��`xNc�P��x�Jkafl{ m��l��8�+���xR��{��F2h:��-� H쮽������k��W�N��u���Y\�+�Ƀ"0���ݧs�-���7y����9A�䷔u���=���T�xa��%֗s��1#�S T�¼WK[L���L�`��-���a�,�v���0j��Kl�G;u>[���9�$�C�©c4��n�f�oj��p�-������� *���hs	;���h��h�;����W�%� ��r\v"�\�k%=�]ͱ� +,�t�G�Z��c07Z���+ҫ�\y�-|H���!��l����۬�ױAI���tC �ڋ�vk0KX3/��R[�q|*����]���a^�Ε�폸>"��ݐz�.I�ZԮ�)5m��&�}���r��օW:#Xr��咫 ٞ}!���!�\~��.�.څ
�C��u�h�F����a�.�c�x'i>�|�ٷ�:u�6�m^��v��Wk8��p�6%�h�F�!�L�vM8N[��4�q����]���a��1Ã��*�|}���e�iu��&��kg���7gA�)��uؼ��D�(~��zT[y*�*q�h_Gu�/Jt�� ����N0%�#�f'��nڋ/�Z%��z�c��7�Z�2�n�>��w��[�hiA��t-���Tt�Q����|'�ѭ�P+s&R�x�!�'1�0�ud�5	Z�k�3�]w���e.�}���mVk����8�)u��oZ��F��[]�9����91mv�O�駗�����sf�x�͛�e�;k�x��N�RYd�.�\t�_.J5\�X�˭��^��<7R�c���d��w�n�\[YA�׾v��\�Y�90��@r
c�����4Q��1]�C���#)4d&�b2��Z��kl�(WبQȎ�۲�O6�B>��Q�Ek�*nNAŋB{�o`Q�����Η9#�����x�gZ���̡oY꼻��
����ea��\S��������љJ�RǸ{����EJ��4\���8Rb�,�M��'oE7K������#O78SΑ��J;��h�]��]�	*9��]:3m��f�����-_ƆkhX��uQ���{��{�љ���ZN��ڿ}�ӡ���cA;�>X�e�a����ۢ��H}ܕ���u�B����&<�t���#��� -�[����lg&D�����qe�V��#X��+��ɇ���B�]k����M����ue��1_�w�h:�[Ed'B�춵5�!rj�*4K����pKz�8ړ#�k᧩�\�xjj������7@ꚃd�N+n��oo:���*�����]hnX�Z�n�t��"��Y �}�&�2���gge�|]!Q��ې^6!�k@���Sg(c+\m]����
@��I�t���z�-�1���)�w�0(�R"ou���,���E��a($�_iͣf6�3�N�f����+v�*vT�(���t�53�渚դ�jQ�Q�z�0v� z�`��P�z$�Gt��|f_4��oSm��J��/����^��֠���®�|9T�K���Ks�k�A���g�e�9��tzt�՛W�~-�[A�����#�zv;�9�uj��U��׌0GY�̍�qm� �s��7V6Xg3ܗ
�� �93�fꌚT9�aT�F��꼇�k�pYM��6��wY�_t���pB���\a\C��~�V���rn�n�����Wի��l.վ��h�g���}�,��I��T����d�:'�}+�rWh|�}6Yuf��k)=2�vr�t�&t	���=�懳Q�����x�R��[��b�H<-v�J� �e�L��oRu���T�s�n���PW7����^S�1��>b��X�2�U�J��0Ur�Ea�\�R�V�`e����T[20���RܵL�5��(1�QTi`�Z�fdq��V�V兌�ƃi\cJ����e�"�ci[J �bʊ&Z�\�m����J�-e��*
[hؗ)[hLb(�
�q�ZZTm�F���R��hbE��E�m�噅\d�"��a�P�AH(R�**(���*��Y��X�m(̉�Ce��R�c�9p̲�jbS-nf!QE�`���r�d���Y�I��+��m
���s	X,\T
��1�AT�
�(*�[-YY�(�ƨ��
 �*���["����Җ��rɈ���0R�+��j�*T��Q!ib�̶e�c-��KQR,��
V�V..R����o���>�~��ٳ<�D���ܓ���7W�1�����ز<r����=��v^���*��k���v��΀�����w-�Ze/�M�p�����7q���A�|9�P�:z���q�2� �7�Cy����=��:���w7��TG&g�D)�X4IZ@(ճ[I��
s�D�
Nu�s�P}1[Y�*�-{S��i8��)�s޺�"q�lhf�N\���+�,���><ڿx9��&��WU�Uz�	ξO��_\G��^w�g��8|̪wʪxc���5�p��u�n��*��o������w�dLGs�0���"�Y}�bU��F�W�ʇPݽ���k�|��o��I���PeF8�>FBp</�:�	Ҏr��oOX�����5Hd]Qg�W*�u5��Ъ�� �v�f��*�e��)�{����^�>�P�N�E���:�w*�u}-����gJ�qq3�gY�o9q��¦�˙��ʋ�x�f�9[�su����-������3|8�С+L7L�հ������]l}̅'537�u�\����lB���#�\�lR�Zh׷u%��줝q[�(����x_�z�<��}�8�^�]P�:Q�X+�]���|��Wu�eolw��.֐�ZyP����z��X$���^mh��M�N�i�>6ព�}Y�����YVWx�:y<\�
�[8�Zu��=��m,ɪ]����%VLަ�{�j�E��mT��m����6��{�8��m��ǩ��PY^-�E���qҸu8�0倪9ℐڪ���Y��)��/�^{�E����r�W�׻R�M��e{�ĥ�נ�^η�_tj�1oy\2���C��F��Suq	�[�)�U���u8��T*�^���O:�6TL$�e���ɴ3F���P�R�t�W!f5��A�ռ.������|��N^��j��c�MNY51<�.�
�*S�]3>��b�+����E辕^��/X�c��H���+)c��ϛ�Qxi��v��Z돎E�*��]������ss�_
�Ų�Օ�/p8)C�	�4�,�܂�!�O���]'�c�C7]t�>�/)5���oi륊�1r��0�K�y1we�Ϭ%y7X�N�b4���P�Q�!��v�.��G�n��I�3���@��Z�vqݴ��Ğx�;��Y���u;R�0v�m��0���un$�I4e���m܋Oh��3[�o�[��� ��8��i�j��Z,�,qWl��MdIN�.&�.�G����e+�1.�X��g�v+�"�0��zD���9�r���c:kS�]ҭ���yr��rTW��pe'��s^�x;�S����m���Y����٬�4�.[��Q^�[q�k}�r�=2���������i��9*�ӣO�~����#��j�RG�6��ivx���z�&��7ɞm�=�ki��ndNL�S}Qr�}x����n�jgr�%�obC,8����ϳ�β��n��a��e;���U�N����-��rz�b<��)�/]�K���_�[\��OE0� �=�d[�kY�����ŷ�݌����=�xubB}i[��aN�R_gBH�}�U�"��p�=�U(&�ճ&վ
�]�Jz�j�>Nᗅ��h���Z�Φ�[�y�R.�c��}bmt�x��z^�Y��Q�sjJ�H���L��*6VqSD��ĜL�a\s1XgMv��$�@V�S#�:��]��U��� `�[�*� {��n�*fl�%�i���Whޮ�'C����U�"����%��v�m�f�b��u��?#�cbCk 
�#��m4z�O9{��B�ɴVRsяF>҅���̷�6�d�.��/D9X4O�-�
�A�8��ݬHﯙz�|��o�<1J��)f����i�S3q�-��<��ۻ�캠58�ά�8�d����Ĵ���Lʑ(L��N���o�-]�kB�~9�K�u�o�q�^�/��@N�9ő�6��%���7%�����>���q�ڲ����^ʺo,��w��]3�P�dʼUu�j�~����3U�=yg�yC�Z���	ԟ���1?y�{%/#75�c~�$��P�������2�eeE�m�#r�[�u�\©�����t��I�{��nmW/&g�"��0qx�C���b�K���[����UVۋ�������T����w�s2w�i��
=����T�{�.���� �g>�H�eK�6�rW2Pީ���5CWW�K@!�:��{�vC��gff�%���DWw���Q%γG�	Ws�Ck� �y���cI+�76�DE��	ݰ��GS]���n���͉�T�RU9��W.%M�N6�#9�^��c��o����-A����sm�W'�v�-3J���9Ǯ}N6���	�Zv��8����o��%��z�+{��z����xvW�:�YNz�ep�JҖzZ8�ڿUߵ?O`x��9��Sg'��leG0�Azz(.Ȩ+k�au�D�#k#��̸܍Nv�����\9����n���ah������WU��^	��;��z���]˭ۚ��׹E.u9ҹ�ñ	B������n��[���W�ua�m����]gx�aK��Rtc{z���<��5���)�M�rq�!�S鼉YU��p�wn�)�<ڠ��n��s$��(�R�9}r��Uy��b���U�,�1��2�נ��Үʬ)���>�V�����7[c�޼��/h
����6�G���
�09����VY�?��;�1���6��Q�t>�� ^e��騯/:5���@��o��8�k�[��V<:k�媆�X弟�OW,�w�u�ŋ_tޡc4��n\�d�0���&�i�jD���Y&K�����O�VДo$o��\���\�v,��q��8��pdJ�P;�ğ�K9�NK��Y7��J��oR�S�fU��ν�.:v:��OE4.�5�1�ɞc5����'��4h�L|�8�}��s$�x^}�ʹ�Y���հ�*>�ڜ��Ksg��]1|a�~G�Jpy�x�e��8��j�xet�}=�F������ٍɤ�<���z�v�Hp��7���u��>�P���r�UfŔ�;5$UWn����{~[˺��b�����OL��l�&:� ���`�V��(�9nvb�!N+qȩ��#J�M�OS���[��=sN;[��1'*����x+Ww�\��~�S
w���edq�)�j�w�wB3�F��ȥ:f�6�����YCw����giP��*�^ctϞ�k3s#f�^���tUR�0�v`����U����mby��Pb�w7O����իG,䘳����^An9y��"и�\wVNē�랒b�C���/s�w��G&��QT����l��3¹�G0z�7�B雜��l�֣3�Gl��7R����}�Xi�՞l���냪��z�<m�`Z{ۮ�=7�E�=._\=�R�$�7%^���5p�pYTa�Q"��#���8&��O\rZ�$�ըW�����}�x��w���v�V6�� �g{��/�Lt�{»<�y�U��h{��y2j��\TgF��Jv���Voe�i*��Y;1�}}b��O=�a��8�j�I
����������!d�l����U��$��D�N���Y��y��F^�6��d�3���\d0��,����qdO6f!N�TECʚ]ܕ�rট����ҧ7���Q���\��SB�E�5�ia�;�.xzn�8/����`�p����-�����k���]��� Ah�Nx��ac�$�ԔR�<�e|ϖ����Ë�I��{�\�z��-�����v���ϔ��b̭���s�{d�o�c�a�*ȭ�i�^V�^����ޭٕf�mk��̛O�=g}E�Xt �:��v��<+�I{���@���0ox^o1������ƟJӽ}�G��\�d�ў�R��w�9�e�QE�ݪ�^�nZ��\��:!�l\u.R��jR���E:Y
�'9��J��鶌������������d#o���C�6�jឹ��4��HLZV�r�)s�u�3O���v.:td��/N�Fp�k�Ȩ�9��t�x���3�Ӽ�s�"��Wx�榮q^W~jTr�,w�+J��=0]r��x��\Xx_gQJ��Ԓ����V�M�'E�e腐�lHo�B���ki��E�*m!��ΩnM.�z�sm�r⚣	�0�L:����~
맪�D r�=�kVOε�b͢��T뒬����*FS�A�Zo'�^@�è�^92T<�֓o��Q�)u������]d'Dl*dh��3	��w��8�Q�xxa\oWeQ�~<���竷��4�uY��+V��r��]�t�|հ�n^�Y����ί�W�{j64
�$k:"�����6[����N]��7��A�F���VR��d}��1������zA����n����wf�!R�oh:B8���׽�+k�f���}�*Z�+MՙN��=}|�0&��F���ʥ3_�`X�2{c=z��{ʯ��6OZ����y_�	��p��t���B�ryUGv�\�.�5�%�J/+r��q�b�i�ֳ2o���d��O�[[�<�{��F���kݺ���}Jߑ�	���%r�g���N��*R��3��CڱI��O�����g���u��W�9!X�מ�z�5�����9/�G/bǵ�����];��r�V�V,�MRQؘ�f�-��ǖ�\�^5�Ğ�.���U��RU�hꙻ�䙼�ӑQ�b�l�LrBS����`�$vf�w٬7��=��<;* ���{
��Kǡ�T�F�҇Mi9<�7$|��u��ɱݒ���L7E��.�®��Q��;
}u��=���KL�s�N��9��웄�ܼ��B�É�ϰWE�=�ӥ�N�I��e��w�!{�_x�S��'s/��&\=�[�����D,ޥJ.�-��dᡄq����B�s�����a��Iɱ(�Iաъ���E-ʐh�uQ��\m���f��a�*u�]�ۙ�ohD{��V��^��G�U��w��r��m	�J>A��i�(��wo�٢ӯM|�x��δ�,F��Hf��]�'[8�]�^�s�J�oԝ�f�r:umsN=5�E�Q�/u\���s�}�w��^�����g8�fv��3{-.Y��k6���f|�J��/]���Ϡ��U鏥}t|��q��R�L7����yص�ف���5��yő1͙R����^�J�Z��]��Lo]�+.�r�{D�f58T�Pв'���x_ ui;ysw�*`�������TS�\v����b:��S^���+���k�c����i��;+W8��w{����b9�2��wo��V�>�l>��r�g����A��؈��I��W3Az��i�ΚřU��eF^5y������/v+C{�w9k��
ޞ��UW0r������سz�Z��LTf�X.���λ՚�^�iԱ�jN,��xky=��4���.^u,��1�A�w�_�;"�Xf�Kz�R*���5,�z�1=��_V���BG���(p��}H1M��I��f�����k��V�L�L����WY��)X�;��ɴT�J{����Sz֊�p%&U�lyRl�ʀ#��P�:s7�&t�z�n�>��Mq�|ĩur��{WkM�0ffSؔ\Y�x��QX%j��cn��PB�t�1��7y`55Y���������S���z��'W�p	og��c���{�Rr�+�555iT:�)ҭ8� M��bץ�tRkVSs$��z��n�fM�l��.\����u5������t��
�	�8��:3�n�3��6S�gE�x'i�1����Zz���sF���2-��f:1j��Ҳ�:�n��Sf��%�n��d&U��IvG�N�zV��;�
Ff�M��wCB�6zq��D�K����S��f��E���{ɸ�n��d<��!�5�SYh��@^哴�aeOཛྷP�);�/���8�X��[Ʒ[rلg}�j4OY�H	wծ�V�V<#d�ke(m�nZ��Pu)��H��g1��D���ڝ���^;���t���$:��s�q�N�x�q�L����̤5�-Z���o��t��ѳ|&��N{�%�����CP�	�8�2ήѓ\���n��t�\��"�2,����k�Zp���@N֝�ɥ���p��΃5f��4����������4�%m͌�^j��R����4D��7}�e���T�(:��\�*ģ���c3B�z9i�G�Ve�C2�󭻰�J�f�)e�w�B3�I�l,�Tzsf:���*��w��īkq��2�1e�T����-��u��f�:)��@��y������v������;;���ՇM�T��p$h;i=ld�mɠ G
�bЖ��b@U�u��cb9O/��O�+8��Rݻ�Yyΰ�6�t���Tb|�9���&���׈�e�
;7���'�\Ty��{c#�U� �=��'ɷN�/���^���:�/��l좬��"��W*��Y�NX Y�1Cc��jF�4�`�Y��]��>*����q�v�m0(�z�%�gq8�`^�Ik�V#Օ����Ңw��;��S'�Pe2�yٚŢ&�OgΣ=)�,�VY]�ܭã����G�鐆�<��݇�0��NA%�(�{s_T�yoZ��4*�,�8+��Pinv�q[������k�ؖ���Yq-�)ĝ���]%Q��f�$]��C��}�I�uO�㒮.W�!FmD=��s��	M�a�.���Աµ.�)�k���� p�mv��墵������>}4����t�BΩ�yN�e`J��x�ٮ��&�?�p������p��]]^��+�Ge�s��_[���D�T,�*�-b�#�*����ц�*"��PU��9�}�Y|�?#�$�
�b����ʊj[Q�A`)P�lQ�V�b���%E��T��*�+ �+[m�"�1b%eA��P*ҕ[�*[@TT�*Kh���E�*�%B��q��ũUX(��V�)lm��1��La�8�%h�X���%���0Dr�`�c6Хn4G-��)�S�آ�*��)m�*��V����*[T(��X�ŭE���D��J�Ah�KK���T��EAEUA�"�R�����PF
UV[J��(%d�(��5�J�V��*X�V-[@Z�c"�#F��YPKIcZ��h�AUbV�EPm"��F� ��V(����Q��QJ5��Db���X�1�T�R�6���-k,����X%)([dkDTP+Q`��
�*E�B��b�潻��/�����4�Q4s�}{�{F�X��>�6^p;�Iv;���:���3��7қ̒v�.E�^G}�ҹtȢPn%�n��׌{��(�n�;���닻�夿K�o����m�����m[��μm����m��7O�B��c�z��y��Z�n=��>�s.�F8Z�v�Z�R�yZ/�VDq�)�����!U���unwj�ƴ�v*
�k!�W>�����1,�P�c��;.�aȓz��n�1	yZ;��P{\VL���g͸��w8WwU��5[��b�+��N3=���7�8+��մ����AYl�hyʲ]#��v;U�\�+��:�&�uD�p�>LC�X�Kg.VU@j�.�9Oo��\�J�N6�Sw��(��2�� ۴�d_��1P��AW�c�R�m��x����d'ǹ=�Т�2���\(N�xB��N,��l���.���j+s�~!w��>�t\�`' 'b�\Y�/�v��A�6פ�wd��ez�
�}@�T�eS�YE�������pe'�b�	!,�����o�=)���u�Ž��E�J��
Cr�X���긲��X�΢2+�X��w�L�(��o���'w�\�;G��&�R�zo�d�}�ڹܲӽ�p,v[�{��uV�5z�Usehꗙ �r�*3_ח鵕7M�EE{հ�n�7S�\�����$�����Uz�|�˝.��_K���N�����є=L��>�|������{��v�S�i|��p/.���������C�姡�Z��[	9ׯo����ՙ5I���z���{N�������^U(���XМ�j�)So5���ٺav�M;�X���]���	�f��
�ꊷ�Wpϒ�^S��9�G���Y��t����f�L�~���â�5,�=s�=^+��v�ؕv(sy�p�[�,���-e��+��1;j�%`�#�m�7�;k&��H���,O;�Nz���1��ev����p9s�(�0�ۈN�{���
���!���W�,q�-9\5V>X����j�T&���+�E�XJ�?1)�P� %��~�x=F*<6��B�7�M��Pz�v�[�.Eoi�/H�jNg��V�;m�%��c�X�g9��L���V��4e`�|H�]�9M,�Z�P��66��Z�t[�<�>�{BQ_`�uf\����O����K���N��erĕ�i�\+Fv��+zS��f�-<10��bT)��М˝����U���Eϧ��;)�Uf1��:ۿ7<"�
��U����z�,�[r_�D���gؕf�d^J�"]y�;�
9�$�<[�z�osa�h��6^�y3����ϫmTe�w{|��������ݏV�y��c�R�;�CBȝp9�y�^ur���U??fޤ��a����G�T��{���C�e���9�����k���rx'��C<�������Y]�*ڡ:����=���Y���m����y��~EQچ׼�F[���ݨQ;���n�J����qx�^$+yRzz*�վQ�+�n�f�U��O]������^g��o��;�$���ܓ���2q����'̝d���MoY>O���=�Ѓ�Q�1D�ۦ��μ�<C��!����!����̓��<����z��3���'Ȱ�)��^s$��S�d��I��N2r��1z#����N����ع.�wD�?�����[���v)K2�{�wvK�3a�ՄV|o�
�sF޼��	�E����ei��L�j��Q�����ɋdcy.�4�c�M�;M��2G]1ƞ=�ˣ.����І�yηz�����K;m�O�zx.�����y�����>���&0=N����l��7���g�C���'bw
�Y'��g�+'Y�!�ì�$��!���y���!.c�������~Go���Qu�?�[����~�8��|��0?$��y�r�u5�a��'R{���g�M3���d&�T5���	�<3�VM����N$�O�a�P8��'y�������3����o�{�"#�s��=�#=�&�x���8�ğ3l��̀�M{�?3l�3H��'P���ߺ��4��U�q�w
ɴP����_�k]�k?s���3�}�}@��I��h�x~̄�B���u��|j��Y�����m��3i��a)�sP�'���s$�����<;�	Ԙ�~���;�|*�^����r�� ��D}�'�L{�=-l�['���Rx�]�'��C����I�<g�쳌'�O&s����i����h���Ý�Ԫ�^���٬����b��Ey���{.b<�1��k�3�$�1I��'�5�@��I�Of�8����3�	�C�t=ġy>����=OM^�O�*>���_w�5u�}�u߿{�a�:�i97CL������:�䘋<9��0��aud�a�o�+_�'}ϵi1�ɉ8���|�q���p+?2x�$y���3^������ر� ����L!�A��+$�<�X"��h(2e��o�!�La��aua:����La�~a;�d��>d�Vd6�3���s����륫yE�����=�6b���c�G���d�.�I�L�̇U�q<.���'ք�垠zɖ��܀�VL�s�N�nҰ���q?_m�g�kOnv>N�����$�fWoވ��D}GИO�y��Hu	�x�2u�I��O�4���n�)8��ú�M3�s!ԟ��y�d���4����a���o�'�ۆ��=#�T�;J���+��*"Q��,�]7��-�_~��p�k�!̰���YMٽ�^NS�\"�-�;��G��FN�d��V:�wK*v�V���������:8Y�Yq���z/���QTD֣ܛ�J�t�E�^������Ky�9��4H��D~{0Ly��	�й�>C�|��׹8�>a�Y:Ρ?}!�d���:���Bz������I�xs�X|�Br���7c�*��|�o���4z#�{�����#Dz��n�	X������x�uB|��5<�RO�x{����5=�	�N"��O�8����	�'Y�w�M�t�{5����B_���5G�z>�C�̇���~`~C�4Ý�|�b����Y
��{��d��C�Y��&�3�I�'��N"�y�';l������^�۩t�݉}""4{�L}�ݟz�eg�OP����OS�!���ԇ�?3L=�w���	�����<Hh3���'�iu`m�I5�0Y'�^s�����]�O���9kg�y��z��}��O�+	? u�����Cl3G5�רN��o2Cl��zw�ԇ�?3L=�w
�2M����Y8ϒܝI�'Ȱ�z�ƭ�'+���;�?>��]�����菽��a? _?d��I��d�$=C�$���}d:��k�y�����ZCl��L����O�V�p�u$�5���h�L�J�>�ںC~�� "=�����Xxe��O7�$�'�;�n�N3��@�:����C�m?r�Y��{����d�����1�u���>����w����}�y��q
�^R��8�O�²mAݝI�Om�� zɯ7�Bq�{I�i'�2M��?0=����O���o}�M����L�����ސ�/?}LW�Uh���M���=d�qP�B�~��
�$���VN[	{N�m'�I�h@�����q��<�����c&���3�Ѡ^E7�;���*�~��X����1&�'��CL��H�i�f�d6Ɉt�p���Iϛ����q�?2{�'$��^�'�����������Z�=i�k�pX�ʀLw�g��^�����;��:ke`���#2��K�Y�����{R���4������&V.�]�&�]�<]St�0�:�{ ����OF���We�e18f��dwq�U���\�c}�����}�[w��~�G��G�{�F�|=��X�b�C�u$�9��'����2I�&"�;�tA@�4r�,��5��_{��{�u��=#D{����f>������&�c?!8�t<�ğ����Y��G׬��+5��8�$��ì�"���C�>d�a��C��9>2}�{���(sy��7�Y1y�9϶�����'O�3�@�O�<5a�C�1�>��d4{Ou'�q���AC:�^����~��Qd��N�<�C}��x��l���~w]y3���u�z��?g�Ѧ8~��O�'S˙���Of�8��f��wRz�0���1���O���i�����O��Qa1����3��4�Z�[�ԣ�}7]{�F{���0�=(x����Y0�s�N�xs2V|��N��2�����Y�I��$�By�=a�N*��'�:��wǾ���o���};����"#e�GQ�z�G����&��r��=a�iݰC���aP�9�$�����Y�>d��ru�|���$�)#��ϻ���矩��������VGG�D1�����'�NZkvhMo�C�XO�s����	�~���SHs�O�C��~�	X=��m'�i���2z������^�
V!��z=��Q�1� ����'�N���'�`q��'�Oݳ��	�wxI��	�o�Hm�$��'̅C�\���m������<�{�s|��y�������L�Ci4ɠ��$��^o	�XM�Y8��`{�'����62`q3����	���é8͡=;������iw�}�G;�<���������Y����=r�|����a�'���)���G��a6��9�v�&��$�'-��hq!��S��!��O!�#�W��E�O3�6�/1�(�U�����Ė��5C�֓�e9�����O8@L}HԠ2��beaytR�!���]�V'YW�[�E���u<-j�)5ٺEtE�g��ί
���޵Τ�d�Qӻn�ؿ��lj\�' ݜӡv������z"#�:۞X����
/}"��~�w5	���w��gY&�ܢɴP�w��6ɵIXC��g]I6���v�q�$�O0=a��i?'���;��f�몾}z��=���=����s�u��1����O�V��+6�u�*M���]��M�}l�<I��I6��;��6�q�����޳Y�_������k�� x����~d6���{��AH|�y=`z� ~;ܓ�<d�u��u&0�aQd�g;�&$�(OŽ@�'���h@���9����_:���/�z�D�m���1菽6�=#���=��L���2ΰ:��|��a�:�79��A�'�i��'i��9�	�1�A��TXN$���VO��y����u�o�����������x��)>Hx�I�d&��~���	�<>�u����e8�~aԼ��:�>�9���R��C�>d�SÞ`N$�k���������5��_m�+pQ���=��Dq>�9Ɂ���Ɍ�`x�I��d��w�$�C�ϲé<g���|�L��!�u��{/2I�)�}�I�׻�����n��]�&�2��C�
��,��7�V'N�ϵi1���8��&3G�`N$5���d�I�J��|���*s�A�����o_�s�������o��I��a�'��?~�@�-�M�u�5�8�u���&��'N� m�3�'�̇Y��<���3�&��|��:�X{�����?����k�߷%�\�}�==� ^���h��f"�z��N�>�C���zɖ�G��@T�!���'Y5�¡�>Bq=�2��$�Va=a�u�7]��Ͼ���t�y��������<C?"���8��z�E'�`w�$�<�2d�l��y���|釧����Ϲ��2�Ѿ�P����N_w��N���u���p��|YZ�����yYO;>Ÿ��z��y��.��v���+eJ,[�h��< ��s��%c��73�����m>#3����M9�=I����=��Ң��	,uWgN�4v�vT�j��w}Lj����|�����|z��?}�{ތM����[��F���ܘ����Y'�q���ɉ8�'��q���a<@�s�����I�|ì<OY��`~I���I���>{��Ϸ�{���j�}�s���DG�DG�=���zǴA�4ɠ�y8�m'��$�)'�P���~�X~@�'-<9a=@�h�r~z�~a���u'��C{��6f�\9i��S��jC?R�A��}_�Ͼ������+'��!�w!�<d�3�VC�d��1d��h<�I�XM��$�'m�~a�-?�C�C��||�<��G�������5�UV��y����GВ��H&q����!�j���&�O��²x�RL�Chx��,=�Ci=d��0RO�<哶�6�>�q���~ۼ�����߷S/::~]
�����PW�7Bq���u���!�OCy�Rm��C�ΰ�a�y��P�$��m��z�}�ì�$��!���h�ԓhG�ﳶATi���jM��q��z�ѦO�z�`y3��:�׬���u3���6��NZCl��L�p7��'bNس�'Pѝ²m&��H�{D�Ϻ�~w?	�k��w7����$�ә�O�3�C�i'S٫'�=`x}C�3�m����!�׽��6��4����C�LC���Bm�!�> {�Dt*�ɸ�U5�j��[�an�5�
��(N�3h�>����Y5���N$/�'XN'�VI�?0<2�2C�~OC|�P+	�s'X3B"./������H�=1�wm�}Sf�}z�i&!�z�����C���'�I//?2n�>I��<|��q���a����5I�=g�&Y����s",D|=�tl����,�k�WZ�f�e�����4��>�~d�&"���8�2s��d�a���*O�a/��a����T�`|���	�C�7�Y�!�$b���"��5�����H�Su��P�gÀHd��Fu�C<���`�j��bu��y&��s%��B����xV�]/������8IQ�	�Q\�(�7��wEBȵ0J��.Ϩ���k�B�\Hi�ީ[G/o�q�\�xj����1]��w�k�;�j��a~�=�D{q�w&�Ngw�{�=G�g�3�&�����O�`zr��=I��G<�@�7�.��l<�����$��2�W�M�8��1���	��B٤�m�q��1ˠ.5���."C��|����ɴ��N$��Tћ�qY'��x���@��-M�$:Ɍ5�aua:���%a�|�s��m����Ͻy��X^y�\�w�a�2c<��!��<a���m'�X
c��9I�L?s!�d�O��{hN�1�MZ�`z��3}ϜI:�g����׷;�L�n�k��*���A�"����́�Y�'��:�|��Ri�>7g�i���O~�?2x���M$�o���4�n�`|�C���x���U���Ja�^W�C$�����>����:�>��C�~Bu���>C�|����I�r��u	���I�N"���ԝI�_7Bz����d9�P�ί��jk���9��W5[��\�}��!;?~���O]!�;�@Y1'��P�0=�0�|�̞��zj��4�י�RO�VN+$�ϰ�d�,�}I�{��������t�����zǹ?P�'�<���q������������i��;�~d1�?wR���hm��<f��j�|��5�0Y'��'O{kbר޿���*Ϣy[9�}Ǣ4����d��`u�޲|�$��ì<O����H~C�4���2O�O���&$�R�Xm2|ϐ�Հ��B<���}I����t�o�������{l�oFM��0��d�8���`q���j|�	ԋ��z�o�Τ?!��&�JβM���J��|�u�F���}\�Kw�C�6��1��`�=I!������	�O9�n�&ߙ:�ǉP��4�;���C���������3��?2i�wi&Ь�ﻊ��KRW�
9��c�WU�"�G���m\�z�QLL��G ���/�
dg���l�]�9�9
d��>GZ��-뇌�̙�S�t���ϽL��T��,Եx.�O��J�� �H��%�؟c2��A\ec�x(�iu���/xV��2�.ѽ޹=���=�K7|�{�7��2�����fz��	��ɴ�d��2k��M�o9�n�N3���M��:��08���x}� �M{�����y�]��[K�������}�/�'�6Ɍ�촓�Vo�*,��k�²uCE�N$�'���q'�y�j�3�O��Oud���ǽ�B$��Kh��&�����[��{￸Aa3^d6��4��?d�C�Lf�op'Y1N�¢�8�������3�ui>jOL����m���F��Ǭ|"=���#�z�r�\��}&�8m&��ܳ��=g�������$=f�5�$�&"͝��&���XN�紬��$��3�a����>�����;��g���1����4o_o��'��+?!:��Y8�����c�I�
˺C�'g;�C�O�!�d:��LE��!Ԙ��k%Ւq��`�{��{�g碦�`���=����Mf��i�'�:jɶ�c/�`N2n����u>�d�k��I�����:�$����z����OY2�|�=���`־�>�Fc^v|���,����c'g��䓞�@�O�<5a�C�1���	�C��u��8���AC:���	Y*`~�Qd�IT|��
�9aW\�ð~˅\�?.�W����Wڬ��=C��u�T�9�[��F��ڍDVV��9s���Yި����~�O�׽��J��h罨�S��z��{V6�F���reW���}SO��Y�7��b ���wrcm�����z�u~��C�8��w��̹��:���!�.I���b6�̙�V�+��֘���[����`���c�jI�}����V�|��2Ǫa���},�.I!�ȵ��N��T�-s�ϕW����{|�xɄB���d޾��/�YX��W�L��8܏�ݶE�\� }��ׅL���ƝS�*�Z+&����h���ڛ�bY�^q{�¦��m�S����L�;^�\��J���.�3�� Z���h�bMY�#�Q���٭�2�V}.�oA]-���[��M��P��w}�
�a_ѡ1�E-�kW�e��:-�x��v1���<�:Y��GvV>���ͱ��q����(�d ��\s"�	4J�3j�Q�bܛ}E�{bw�_i�u�����¹	b>K ���q�{Iw������TWH1�c�q_yY����*��秦�S��5�v��q��6�1��q��uh��{l�.{�m V�U�r���δ��C����j7�����$����/p�˺�z��u���U�A&��sh�^#{G��\˩`떦:��T&3^�IBu���j�V�w��`b��⡯��Wʈ��tP�s�ŴF����b�&���X�����S�Yw9����<��YCݗ�r���;�	���jȚ#5��	q��j�]h�ɑ"A�8l@H�Y-<uUőa�4���-�se����ڕ��1��0�2�n�F��RYՃ&�Ώ����wt��(�Y��cx�%8�D�e���R�&�i�]���^�t%����D�x��\�&Qd��c'�$Qu�����t���MQ�V��sq�;�+
�|�Ǔ�EJ`���,�jR��7�b��BڱV�Hbb��q�ڔ(=��B�O`�x�g.��Α�O� �Uٵ�ڐlU�]B�Pm�0� i=���3��t_*�3��-��.�����z ��a-��x�>�]�ʖ�c+],B;3�q�Y���f��m2�ի��*!P`Ʉ$j��Kw_��Z���L辶I�(nf�	s�upQ�{ ����7�Fi�|t`�ϰ͉�r���[���'Z��+�c��k�Ai#���oҨ^�Iw�c�c�:���m�F�]�6�r1�X/7;eu��.9k#[��ky�G��{)��^�>Gӣ�b�:��ψ�t��_j\́����4.hӑ7��1N���:�5�����8�[^B���fL�}3{mwz���FQn��M$�#3u\Ʋ�#�{��B�S�`L���T���Pk	5��F+�;�\���T��ʊ��ò�������xP�((�����2�*ȷ3���r/x�ktgm���[I�U��i�+�LVU�������u4�G_-��G��)�Ź�a2��n&�^rp؛Y-+�+b6�*IQhҍY��i�T�P�e;����� ��zpSK��|�`  �m��j,EQ�TEB�b�TB�U��U�Pb�6�VJն6�"��kU���U���X�E[e+l*��
�R����b6���j�Q`ڪJ,���
�����d�X�"(*��k*[V)@m�У��V-�eT�
�Ql���*���EU�X��-�PU-�%V
*!Z�TR�`����"h��X���R��
���,�-�j*�����YmR(�ŕ�PD+ڔJ0��EUdF��"B���aZ����VV*B���TPKIR��H(��YPJ�Զ�,XVA�6ŢEDEXJD����
����Z��+%��ʩmZ�jZ���KK�+���J���%V�%J�,�UJ�em�[-h��["�P�ږ��*4B���0X�#R�o�}��/�~��֦o��7|;9"Y� ���Zb�A��9fcx1�^��KE�G���	x{�LŰr;�YF�u~�Dz=�c�z�C��}Z��Op�]E�?'�͝�`���]|q旳}z�/4�\v����_lf�7�^��{p�n��Ò!neWh�@����on���x�9�-ڋ�S�٦�1!9����F�ַ��b�(.�y���jO�w�f��?VOFx��I��HLZ�v�*��.64�5�,�͜�ym�RF�Xz8t`���)��lg�{�к�ղ�����-�sM�%��Z|�x;/��<;��+��D�Ɗ7�8�OA2�"fmt��W8��9�6�FZ�rے��f!�0�lLz !�j�L\j��b�$T���{'���AN��c���b�va���CV�֢��ŭ�m�F�pH���s�ъ�-��Z|��.S�^5���n�I�v�k�_d���\��<�M6ףt/S��Q��}��m��1�;H�	,���N���"O5b�ˍ�l6�zձnd�|д:a��>E=��tA�n����w��R�G���}��[�S"��C+ve	��WN�0�@y]mc����2�뫐~{T�=�s�~��-��Q]�oxY�������n�.��ݞh����Q��U�����ږ��n�1U�+# �⹝̓�vܪ댘��qd&�)���D�g�6%��\�A�M��J�_�/�(�J��^�ޫ���T4,��p�=����^�'nv�Wnq�����f��v���\M�qв;��_��һ��pF+&����0_�U��N�e�76�|�Zs���ox:��Q��/��l�bݦ�	�98{�ɏ��6����9J�~�uR��ީ�÷�y��3�u�X�o!^�w�O4��$�V�yE�d���(٦�����QSW��W���&�>�;��?7��|�Bk=�d\��4����8�p�Tf$�r+R�w{|�5�q���i����W�sڨ�<��ys+�ъ�C̕��9�Tq��Tb�X�;�p���v�v����0�ca��Yϫ�ƕ��3,^li^�U��b�y�N�:���l��s���������4+\{��Ӗ�Ɛ��v&[gU���GX�fPK_L�h>�]yx���S�¤�#	HӶygQ�u��f�{
>���I���y��5��T���ԑg� ks�ވ�z"4�x�gk��U��st:�U=N�vu�uz�t]��wP0���)��(ƻ��5���k����ס:�P'�ܿz�����iRHT��]l�hT� ;�۝𝗮�B갖�=��z,��=E��Oe�}�׉�T�q��a��ዺ��ۿpQ������V)�q�O�m\7<1^T̩�#��w�v�Y���U�gt�-G��ʏ���4Ug��=]�x֦�H�&)�H�At���d��
�ˌ���O��.�n"{�j��N�
�PΧ
�v+�"y��ysn�e0������]���]��W����}.���[%�ܗЦ1ͤ�����c��5�u��:���}�.z/v��me��>��Q^�n:���:5*�Z�s���;	�zsg�������X�}�9՗�C�n�W<����Y'�C+����r:��.-��И��܎ۖ��r"-�JmL�a۾9��'��ۃ8/�5U۴�2p�j�Jw�y!�7e�X3gI�c�K��z!O]=�X�|V�-��֯%0ޝ�N��aޕz�K���������z#��k�Z�s��4�ԋ�N�i���\������ړQ�i>�>ͫK��|߰Sݞ һ�%o	�lW'=8�Y��n��ͤ�X}7 ���s�@ޘ�+��Z�1�ucB}�ծH�z����MS����R*Ɗ�Ԗ�=���R�4��VE���Q��v�d�W	K�\sR�_l�'��SK*�7=G���3A~��VP��9U��:���,�P�Q��!B��ys��Iv_i�������ƛ�]�S�`�U�X|��ǙHᤨҢ�g75g��WP��7st�����=�аh��`����T��[�ry��$�=��c>ڸ��ӗ����7F)R(�h0ed��1��R�7U��YwK.����6���l�s����S��L�9�p�w/_o�Z�_���ml)ީ�9�y*�XG=J������$X���e��Y:@tjM��������tMI��c��$aE$"��7�^Y)g}�p���J�݂ʑY|�Xtgu�I�#��6��v����MJ�g�n� l���N��?�5��*��K*<�/D�843����I�;wW#�Ӕ�꯽���m�ݥ�'���M���&"W�Sn��a0�
��o9dl�=5Y�+��ݐ�6�v�}r����e�y����9���8�<�y��y��}�)A��X)�w5�;/������[VX���o���W;��k5r�y��\[=���=����v��@�3]�\�I+=P�?y�M�v��]㊊���>��Q��\���m��+-��J"�T��K��3��k%ʙ��������,�P��=w�^d���c4p���j(RRk>��7�U�>��k&f�<�n:��	�v�r��6�q�7Z���T�ݻM��u�$�V���a���J:M&:�	��M	�t�����;[��U�]��w���=��c��A�sQ�_7F���
�(GS�Cf�����9O���/ѣ{G0�{�؟)h���J�hL���_X�k���pY"��:���i�e����{��5+�7�¼����[��K7��]U���8)?a�2S΁�s�����]��/c���H9��.=p��4m�ww�[��}r,�x5r���
Y׵�W3�;�z=�D*�z�tgr���V鞦�j�(ɋZ�m[v^C�
a`P��+T:��Nq�|���u���*��j����={E}{|��ss�MQ�M�����#}�0V���ǵkv�BHQ�!���B�٬.ڥ��g_����VFٕT ŧ�0t;έ\�Y���As
ƇQ7�Tn3�1��2�<�vU�&������S|s�����v	U�^��9�J�qX���1�|�k��
���Z�[�8ۂ�Fs�#�9
^��:��m�^�&��e�c��v������qu�Aq1���82��M"c\�x_���"�Y�#�|s�����D��R�]r�-���{MjO�²sj��#�M/ޮ�ty�w�;ڛ��ߚC������o�b{՝����\���{��W���~�iN,���ݭp,f�\�ϩ������:;%e���*��ͷ��P�+ �mQ6�Ws���兴Pۺ�g\�^��B�_Z�W]�VW%#{��e�Hu�j���~�z�k�2�������d��b0^�<�ވ��ީ���Wr긗	*�Ԭ��s�i�h�s�8������6�#��Y0����<r�ާ��ﾯ����t����Ž�l�������I5s����j�X�7��o�����s�\�[]ٙ]�a�1�i\Cmu�׻2�v#�iڿMTnާ6��k��Q��������&"ӷk����tCm��/��;&:�t���%μ�\�����#\yt�D�^��O[o9T�2���.z�ԮUWh�b�2.��t�Au��=N�,�P���M�辗"M�d�/	5�(�����ZV���w��TP��b���%�ݯy��Om�y����uǵ񵚟t�ӛ/��I�z#�����@�[8�����k�f'�j�Vwm�t�S�����*E0^,$��˕�9�N�u�lN�d�K�=�<�v�Mg�����a�L)��ŧps��b�U���]\����ˢ�|��m+�AS�z8X����1�D_�uߏ�x���K.x��{l��E�R����V��M,}���;&aƸ�8s�k��K��6���k~�|�-�����U��l\�Ev��v#s��y�fV���0>�/]�F��̱��*G`N�g�f�+O\�PU�zM� q{Y�����.�n3�Q�g)3�>]��U�Lo`��;D_�T:n�qJ��X����z#�Ӷ�>}�˂���=�~�֣��@Q���p�'b�# 'ZQ]��I��Y���D��ʽ�J�彲�z�u=�5U>^���W�w��XvX�@��(]O��1��eY�{t��Qz��U1���or�\nϾIC�����p�P9K�w�u'��,��yo�:�e��׼��N��#݁�s��Ȥ�q
�77�^j�̝���Hp�,���,ns�9�����ݪt�決��\�⼅��dj̚�]����b�Vf�
$�={͕9��W'L�c�c�ؐ��v�)�Sm�q}��ݘp���|r�zHa^<��<G"3����ܚ��;��{yծ��ӱ9��vS�mf�-�CQn:,jY
��zj��L�W�L�u˫�f�B�Ӌ��3y�.m.p���h��1у�`�s��T]r���G�Jvcc:+�-]qF���ۂ.y'���	*�j${	�"r��^�8�=�6���z���u�vP�M|�v���1VmL�,�����5V�]I�sɭ���}_}UU�5DO&�Uf�;�Ba'SQO����:c�u1_��?:��#�Y�!�t���O�a�JZq�
�8厽��M������9��D%�F�d�����\�ӉyT;�+�:�y�r�I��ܙ��OJ�it��q��6��=�T2�YgB<+%i�Vtܳ����<e�X��"��M�m�7m=��n��J! F�'���zV�f*�^|�J~V��*��)�"K�'Dx�i���R���5Yرd����j���r��¯
5�(��7������bu=/Ưr�(�wX�{�ε��1��j��^	�&�	��~�`!ن)H����2+kV�c�-��פLPx�>�����XF�Ӄ~ӂq�;]\U�w��Xpe�qR6�'�#4��6OU�\R�K{�+U�'v�g��	��a��� Gds}�L�s�9��� �qW���Ҙ�'HR���Mnwr�DUR}d����q�*f������ì1������gG�x��~% �e�O67A\���$�*�~~K����Ǧ�FA)�%� l��LS��f�V頦{��t&0G8�q]f��ͧx|B2{TR��F�E���o.�dC��9ć>i��E:�M�,����7ꝎJ�L�C}�W�_VƟw�^gu�y���c��W��k�V%#���+:p8j(�͖1�a��;{�n\�f�u%�u�;�F��N�_���(�qxVA�<"��0c�ة�����3][�v�1wrx �땰Ɏ��ԩ	��E�(J�^)�2���
�C�ݖ�eg��Gj�ڸJ�FWK:����y.�1�	�&}�:��K�T�6fE���f�)�|��t~�����?F�
��wk9���\�h癇F\���&*�������֚i�5[�� �:0�g�ږ'�
�Â|Y��~�ޓ���(.o�����m�yI\��~0�Ց��R��	��ğ/�MG��W��T�eM2�횭�Ju9}�7k-I��=N��U�pX|�>�p�v�bA��;HE�ͦ.4�-΋����k���݊4��m��r&lIULO'qC�P�0y��G�F�b�iaP��ٽ��k{P�a���!fi~�$�Ʃ�J��u���wBw�XE�;/�V���?{*+j���Y�2�D�el7y-y:�èe^xp��Ѷ�U�����YFL�-���<mk����M���.`�
�xk�'�)ا���f�]��Gn۹�`�ɮ�?�7�v�E,ǀp��[aS;��:����+PzOxmio+�$1��^崱L���o�ݧi���f��z��g�@`�2����w�L9ϵuNLö@�q�ƣ��K��YR��βX�^��)=r��o�Bҧ�%rN��g~�u����u�$�9� %j���Wj��9u�~m>;v���rR�5���i��p���u��v��,��P�ѭ��i�$*��a͹�k��])�4.	�X^��9��σ,��}��׭����Ӓ�޾�2W�_z4������pvp�#��!6�wN�i���Ļ�5�n���*rIi��wj�$����A=B�W�k�䳯�^�C:bWӗkj�$z�'�n֤.uՠ�� ���r�Y�_a��[-Ҳ����ؽQ�-�:�F��h��T;��`Z׻m�Y��Ӌ��N+�-u_A��{KH��YDS��M�{RO:SԎmX�;:V��`u`�M."WT6��,\���Û���jذ�؛K!4WV�{�b��c�RO��5Ƽgl���J�)�(gf05�u.��R���U���6�V�W��e(�w��'PGp�,v���x|�����jcz@�5�f7´�X�9hDk��\�!x�;Y��c���uۦ�iR�o[a��:`1�E)�l
2�nl7�y�ό���u��у�ű�K�j�t�b�Uo�L�q����*[E��Z�%1oR�1N\����|C�+<'ғ���Ɋ���h��*'�d�H�٢%�t+V[SH >�8��}�o˽�[H�^kB����6KJ��9�6�����,:թ�=v]�(��ma�jc`i�e\4U�s�4�p��3����GsN�[��.��G�Yg��.]�q�%1��1#�An��9D	��v���S95#�d�d�;	�*�Wk֪GZ�5j�"�\�NB�wէ����,Ǜ��Vi�t/�� ���N��U�е�q�j��1�a�<YC�9�3��e3����《�5����֘�J���"�W��
j�����A�V(�oN�1��䛂i�L�7�"��C�sL�귥q"�����Y�n:&��p8��B��+:,�is�7C���ŏv��}��i�iƵ�4d��Nj�p�)F�Iv�n_�t㧀p'yyz+�J�Z�-p����8�I�oU,U��!b=��tjI�d��/5TB��忐��16~W[Y�[���N��\V��e�B�Ʊ���i+Qj���ԕU#m�*
1��F�b��b6���j�E�AUKJƍm��,�Z%�F��E��������
�T��Z�QR���-�VU�PKK*�[h�Klb%kih��*Vڒ�J!D�E��ѫkX���1KV2�E�
�2�+bR�ҪE*��U`���h(���k
�TDP����*T��`��kKe�����Z,mm-�d�+Z�KJE�B����( ŵ�Z4�b������b�EZ�-��`�R`���
�ڲ�E�j�b�*��1B��X1D�
�k+X����h�1�X�(�mQUb�T��iPV0U�m��B4��-��X�[E������������Ҥ������+QEE"�V,��(�"�Ԭ��+"��,���T*�XZZ� �J�IYPQV[jV6�H

�¨ʍ�H,�1Zʂ,dQE*QX[
T(��F���B�bԱIzۿ7��'��q2e
ޅ]=K��4^q3^@c�k�򻃕N�B�>��>�e��g\>' ���w/G�2���g~{���kmk�˥"��\����U��� "�8��\��8�a�j9Đ��a9�{��VYm_k��up\.��%��\Z_�Lua��ռ���lRq	;�b᭭ړ�
*1p]-��wv���vr��<b�м^ �u�ή̆�i��n���N0������W"6��n�)��r����!�ˮ�-W��N1���DQ�5e�꺥+�p6��l?sY�y���Fzz���`�e9lI�EO�޷z��`�~�6����0�����:�P��!�>�b���Vo'2�ft�T�rS���mW9���Ig���ïɈU��v�)fpA��-r����zs���%0��
�TZ���rpJo�%��e�B*Xu��uY�1���cE�=�ׂW%��E��.\�U�ń1E��] �2_#��S2]�`j�V{�^%�)�O��+<�����7B|�hu9��5��E
��;���u�֚�b���񥻝˖t�q�k�{��s>�)|w�p%a��.'��c=Js��%ϯJ�q�
v��70��F�����ɂ�p�ʐC��6�Pʽ������`����з�������+�yJ���������E3�Q'~0��zǥ���Ⱥ�<���Y�8o�찱��6$}x6�ĶU4^�h�23����_{@���lƞex+���֥F��4��f����=C5ų��l{�����h���.�EgF��)}�U�ݍcCWN^�Y�����Q�Rŉ�R��{F�H>��n �2����@(�`��n�-t���ƀ����h�V&K+ʂ>�,$�T��5�����x�4�{�ä��,Mٻ�<��I%,B��E��n��Q&X�"�hzD�֦�[|�L檡"I�rp!\Q]��YΤ�a�s��.A�N\�����w9n�R6�yPܡd�������V�(1L�j��À�� ���2���j��Å9҅��� V��]>!j��Im�~U�c��P�-��C��s�����������S�lG%�&,MF: ��"Fs\@�i���V�xV�������V�m�����C��^�"eG�oA�?k��l`�o���"o{f_�`o���)�W��qU��C�ZT\8�څ�46)Ts4��z��#��:6��,!���}6��v�o�:ϟ����2�X��������60�HEQ
��1��Y+϶��G�ԥ���J��鹩�cvjNH�V��,-�p��W�;9Oqs�/ya�l���C�_:�|��Sw��[�3���F-���~^<�W�ԙk��m`x'JX�J�=J���]���t����{�`��h����aͥ����=*�xx����u�
b]��8�G�	��=t|�f�B��z�͉՚ӡV�3t";e�R��$Jͳ��,X�a��ut��o� *2b�ZK;/oeh��e;�/aD�����N�;ή��\"�|l����:ϯ�=��s.����{jOq�I"�:z��-�B��]h��x��oV�o�����8�9=���j�wK�p���K#]OZ�F%� ����QO�a[uC���������G�F�ud.�f��On�d�(T�%g�d�2��aB�n�E��Fb��)5	��0�wK@��R�s9bSs�R^�K��i�P�+�YK@�8UDO;b�G ])bʻ�b��s�9�>SPέ���az�	���I����2����>�������ߕ��f��f#L�����.z�h��� @�����7^����ן-Q�U����V�J9�Ia��5�V�Ź��R�Y�lt��<�ؒXb��Hb�UhX&z�]5��5+�]x:�'��Y(jы��uWh�W���w&�ޒ���o*i�<��Y�bz^5OF����Yh�s`�!�x�iRܲ"yK� �c4��\gwV�|�b5(�8f4�Z��M������C58�]�;,ʲt��Y��Ijb��
	��	������������ޮY}r���*��z5���PМW��*�baH����a�ѕ0j��/�M�9���on(]f��3��ӂTtŅ]��)k�&�#=Y�D[��Ȭ����t���^o.b��+3�jk���xz������]ܯ#��f����eI�U�LL��g��f�b�������f
�S墦�T{M{
�ux��C�peu^C9�<�+���=�f{�~�
1^��q"�OQ�
lӧ�����c L��ȳ��t%��ϸl�#�dU�8\>M��wM]�HqRY��xVA�<"��	��p6�T�.f]Y�z��I�O*�lc��өJ.J:J�T��P�*�����qt�9�!^d���	�pc���q�Q0��"�Ùb�i����ł��
u�.}��&*y�.�cٱr!X�����.�a~���<�9£//޿o�N��kGy5;w�N�F��!���\bY�^xlr���m�W/Z��XX�����W1�f����"w�Ģ�Z�� ��;3�0�6�N�@�v����i,�*N���=�l�"٘qjWy:����N���V�72�=4zjٞ��ym��K�A�E/j"��8yņ7����8��k=5�hm��7�R����着��Ⓩ�N�*F����}��1P�H�`���t��ay��W��2*|��&ӥ�k���Ǎ��3�͚�\�D�ºBkń+ι��ũ��T����~��3m-��Z�Y@FV�a~*�,am�	C�l"�O�,������Ii7^�C��:؋����>��ڬ�����tl��`�{�*�N�D<�kʡ��3�"hB�1��FkRtp�i&�e.�F�T��5�Lm�e� �) Ƨ��a�8d�pH�8|��0��-��~�S����9�C3⮼4dS�g��Q��Zq�Ø[T"i*za�������l�]���fs�}���*������S�ά��Luo��}ڇ��$)&nY�`��xۍ��7��s֯T����2���[{F�e��P"`c.�e�H�}�3.'��b�~���5t���?j~�7���uµyEX�^��Ѭ��U⣅��ɫ����zޭ=%���e:Qծ�c,./\�'�N�h����j�:cg����WJl�N��º>���+i+o��*G�] ��bЩ��;NP���jR��Yo��;�+{>W������+�DƲ�6ٝv	�!/B�x�nGJWX�F+nm��DȬ����G��	`k��@�S��-m_u+��ѤƥF��w:�'u҆�Ύ�.� l.����͔%-�ˊ�}AN���2��}��}U��>�N�%?F(��zo���6v�|!�6�;P�%���҃�۾��(I�k���ֳ�'[�8|�1tO���J^\OJɋV)V^C�!�|��3��H��G1B$���ѧb�Զ�k
%�+Η�Q��9B�r��7�|��'(X�EY��*���/s�v�;�.µ'І:�^#���{eb]���1�>�[إ����+�o���<c{�����2�54&9L0f!�-6v��X˱�>2'X����N�By�=�+P~����iTHBY�J�(�N�L:�bw�D�+��56�$e[�&O:<��{�D�R�"{n�r�/��؏�T�E:�&�K����c��)���cʴ��o�N����U�X�[Y0ᡁ	�bv��g��y8��b�t5$DNK7u�����vc���xdB}��i�9�?�T\j��y^�Dy}2�C��{�k��e(��$�\��H@���	_o����(�^���?*�>/Lg�6,!�Q��Of+\̗�`F�˫��ȬK=���Dڪ`��̪zb�n�u꧴�l��$�RfMn�kԵ�<tF��u�����^�&����!���+�����ʍq#[�ُ��4�{�W��}Gq�{1k��쫻���q�&���gZ��� �� ��g	%��_�^[u�]�6�gi��\\�C�)~�Pr�xރ���,_���z1�"c܆�a�:%���hu��ʼ{;ˣ��{�P�qVW���
�ì�j���l<s�V��f0z�R����{���1�Ȝ��ᩨ�S<$8���Q�R�Tf� ^	�U�!���z�7jt�Ԫz]q��N�����}�N���o穉�:�X�d����U�Yl1�9#�8*�ykx�U�^M"������Z�DLL`�:=�Oa��q\-J�s��(P�Y~6A��E)�K��&�ݫb{��Çk�-B2�d;bU��F@���S���Uġ*�`B�B�t�fBJv��9�F'�����A�8%8�5��.���h4=$�K��I��K3xx��1�Fw.��&Qʌ~=]5�X��s�!c3'<�Q��,H�|"P��x���T�)B߶��㧦dCGE!�C�F�ߦP�r����ċ�.��º�'[�/�h��e+���{V%}�n-�ت�^�vX�0j�~��z����^ �ּɐu�J��c
Z�L�iCy���G�4�|�4�]�=%��sk�}���w�#�/#�f��r��;�\�|]�-��"�����en.P�ɴv�}���e�ě�{ܬF�����L�����@k���V81�q�0�vŲ�dI�a
�
u��s�Q� �vp�К�q�R%��3�b�����!��62E�:�5�.��b{�0��א*,��ЪX� ��֔f*��y���X�+&*|rW�D����J��v-"���Ap�@`&�,���~�$v$|sY������|)�����0����b��8��ܪ�4\���v�����Z��F� ��1JFV��l��\f��$�K=6>��ko_��z��S�Pv溸����jGQ�k�#6�Η��s��qlny�;���r�v�� r�C�6Xq~���l:��W�^l�1�+o� ��==�U��Rq��R�胎�D!_-���-����|<M��:bVW\�ݙO;�n[�ޔ2��1�S��d�Y�K�%!�X��N���ƅ�5|��]ro���C�-~�aӪ�/�ھ��V�0���˃UY˂�z����V�}��-��r���ve�(y��٦����̮W*��v��,�q��[wXZ�\�e���� ��������L:߳���o�G�kTe��j�)\��K�`@�Gn�$)�C)��i2�М��1l�S�"rjW}�f�6-T���|���>��{޷����t�b~�e"wT��D�ĺ޴1�z5�lVT�xT�*t����9[{�	�9閴,Q�Uئ&w�C�0聆���Tj�,[��b^G�&��*C���Xy�9��o,ס�㪴i�	CZ�B���*z˳,={J��ή�C0��Y&���=��e%{�jl��8螀����ؕL_�ЄOQ����산��|��Mw� ���W{�ҝ懲��f�"a艇^YGA��]zNAS�� 9b��N�/Lf��30�cp��������8�iV
q9VͲɡ�.��t��bD&�a�N����]��B6:كQΫ�GB�yڸ��LV�Ƒ��@)���g�WlM*�E�ō���x����/��s�8��ܿ|fpLL޸ȓ�	3��\� Zr	5������[CtsK�7ɬ�����&;�b��ܱ�e����po����k�;�o�I�$֊)"�˹�����K2$��(��9�����(g�ͳq�4^�_�H|��D�7�JH�3Mk��l>=�!gÀ,�~�(���*�Oe<�b���6� Vk�Z�-c�ZY^����J�3�Q7�����4��ۻ�Z�Fĺ���ba���w]�g����R��8�#i_l�e 2N�' J{G���}܋x��z=�v��m;5]}���ۻ[�8��E�c���	�h�ƧR^�ux��泇�&&�%���x4�FOvB�[4#s,��B�s֯UOl�O3���\7L�.
��=�O��N;z�t�<��j���n`u�1��ΰD�c�.��Y7�k��CyM`g/�ȣ�����g.W��ڀ�(V��UB1�zPCc������^����t�����X��TĽ'isLt��j���e�xR F�\
�9��*��3������	#��q�k×�T���Amw���b�pe]%�é��J^\OE�,!~EQxX}�+����0�W	�Sz�5.��g3���d��R�8Wi�K��9���8��S�]gIܲ��f�O9�9��w�ޚ5'҆�	�h�\��VХTw�lIu�Z��O~�sjLR�dG,n��/�q�{]^ǎ�>�������bb�͆&��@Ba`�"Ce`6Kq�ɜ��d���L�\�A�Z��2�ΒΎfn�h�V&.��Xłt��D�:����q��I�|i�F�Z�ò������Vt�y��Λ�G�zT��������z$�������[�c+q�����v�t��kzS"42�髜#}��l̵�:w�c`u�Ӵd	��4�a�L��t�#V�g]�+P��IZV,|�iq_0� Yz�J�>Ͳ��c��v,gRٍ�T�0u)�"-�kuܱEb���qkԷh6;�up���[XK�-��oq�[�ܠ��J�DY�ؖ�:�#�j��3fZ�k��=;�	��Fm[k(m$��zb�J�q��Y
|�utW �������DǻwR��#.�ܕ�핬��,���P���[ ,�J�`=�یU���";�͝��O����VI��ˠ��ч\����Bj�J�_^�Un��s`�0����뒣>�k�woԘ.�n���ZУ���m�k;��&�3"��%�U:�z�Rn���s�wڐһ�fL����E�AˬZ�R�{w͎U=6m�	­�`�r�����
�Ͳ���}v�p�uK��n��� �V�L��M;o�+ ��{��.���V�I���4W]�&�x�b��W�[���P�&E*��U����A]���v(.��Ut�ht9���^�X2H���\o^u$;#H*n�'+f���P=��lZz�=�D�3�]~ٮ����&mjJ9o�tR���4C�^^�Zk'^��\<Es�/������A�|�k�+�"~�U�z�;���u��b�S<S�U�W!w4>�vc�8�N�Y��*xM�ݻnBT0�o��S\׿�q午��V��@�aZ��q��:����ntJ�׎Aظ;Տ�S`5e@�.9���F�����y��j=��WC�4�p�Gǳn�d��˦��@5���r��d�,�[�ͮyɉǝӈ�>�KFT���Y��zW��[E��<"`&V�w�E�X����;쏯k1�����U�Ճ+�7�.���u�ѩ�h2>P�n��j,�]:*C���Q�b��Ӧ�ܩ���1�<�]]�~�RW��]�����8�-������;�y�o8��^�L�X�����P��ۛ�i�A���"��GwO_a�Y�Ը��첳�E�6��P���{��� �x�q��{M��͜N�}���B�s�W%�d�}v�t�Z�-Њ�];=[Pn��Q��r��M�Z�^� ٧D��5U��u.�r���q��XB�U�۠��t�F�v�Y)p,�˔{�k��JS��@�Q����f$�?��8���-��<LC��-��-���u�֥I}aN�~�*��+)\��M�_Ul.[pR�J�v�QѴ�ҥ(Wj
ݮ�U���Vu]��Aut�c�k5�;���V�G1ui�{G���t;%�-âv��U��&��l��]��{N��%ps�-K�v�v)�4�=��6�z��)mJ����H��J�EZ"�J[mE�UX�J�Ȋ�PX�*�
�%�)5���DE���X��*X��V�@Z�P�E���
�jVJ�dF�Z�h-a*���(,X6�-�*,��X(����F
(VT�m"��Q�+
�Y"�m�T�U�,ejT�Kmd����E��Rj���("�Q�Ad���"�R-kU�VE+Z�i"Ȥ[mIiIU���U���*����-EE�¡D�b�T�!R��ejV[IU�)l��J��d
�jV+mb*"E����6т�0B�e�Ubʊe"��T9f ��"��,1�`�(*�X�QeJ��9s*��AQ���P`�-���U�,��f��+X��Tk-,�����*
LB�W,dĊ)�3*�Z��VJ8��=ךvT �V�8Ù���{ԫZ�-��&<O��t��&�� q=�:��,�(Y���.w��xZ��=����(���}���������u/�ƌ�^��C��}���2)�q5���s5<Խ3�tăTr���t�7�*�}�Q����Fք+(��c���� �|�T���p��#�vS���u���1�����i��e�E�0߄���뢆��~�>3��B�M-��!E)�ú�c:V�Rw����Z�@�� Uo��m�4��I�ٺs�Qh���I� 5
l�w�{^�ֳ����Om+4.c	u�
�O<�*�� ��|1����ŕ��Q�l��ݨ� 6�wt.�եE�q�T�\a�e���%Q��]o�_pr­P���2��>dD[*���g_R�3��^������ߓ��0��*�f�7S���㋺�ug����`���b��8��V#��0����9���,Xt$
҃S��n�\v��W�=����W4��4���o,�aT��fަE��p�=�k�Ŀ��@��[7!�͚
d�lM�Iʺ��Z-�i���ښaLwJ!�&�d��Qn'�Z�J�q��Dc�ܮ���4�����u�w�)�[�.�T_,l|F5�nӻb�j}��X�.�Od�HWWw�m�5���9s2��b�ky>͉f�D:Ś���{�j�xŌ9+4R���j0Ǹ�A;��-��w�o7`�V��:M�$�p�~�ꯪ��{:���]��:�
���S�[�3��)��D�7�"ʘ��<�f�*�*W,�w�2d�.��׿.��T�����]h��k��.���@�yW :9\]g��oS۫�*����;j��T��ߣT��������2M�Rt���,/DKt�=�l�X�sʪ�M/�Ê�p�'W��
�Զ��P�cc��N]��"�J�����8���
������K��<MDڮ�"�軈����:	�LA'zÒQ��%�}���0�_�Y]��#u]IW:���>
�+9T_��1p��. ��:s�ۼI�Y�ׄ��'�m@�C \2� �'!P����\|�b�~Ui̞4��{n�>Ed�F��Ω���%Tk��A�B�y�3}J�-xxR��!>�kQ;K�M	�}�m�c\�r�T��y�22f�a�*/�3�\��-b�5�Lf��1z���
��U��6���\1(������-��L��Fa�^�����眧����6-��hɡ� �X�w��e=�>����k�u���Fn��X���L�u��r��.�py5�Iq���{���Z�s��T�9�U�a���SR���,�Z���s��:�tkV�Mgv2�B/���^�9�N�^���x�����[t%�I�����{����r��m��bH�h�үӌ!��knuO<=R��*\ߣ�4��>\���;����a�V���l3�yqG+��H�3��.��F5^��2��p������̙v���⩶���ǧy�5Ro+�����W���3� ����q"�'��P#f)ӁÍ�2������s����!�bPnf�1�ھ����%�R����Y�4f���Qz�y���_G&��;�t��s\��v1J��W�r�2!��i�J���E��BT
6�*�=�UKu����SB��g�TY�!�\&xõ5����QP�Ǒb��i���j8��CºƊ��<gq�7�reps�LU��0TZo��X�ѭ�ҍxu��������v��v�N�gw�uM�c�M�QT�֏}k;���v�y��l�X�r�uJkB��:+ҥ���w�f̻�浽�,+�5zk=҅L�a���&C9S��]6HGEw��*"�N�*o��BD��ͭK�moD�sӡܺ�o�#C &pLl+�	�+�޶p��oV$8G���;wL>�ƭ�.�m�0,0�(NG�y�M��e�6���v6N\so�O1)�,�t��t�=��2�kol�Y-w�B��zݎO��nj���P��b6��2m���7�U��hGD��6��<ݳ���U�Y֦N�{}���Cz�l-�앢>�1���Γ~SfSe�U�.`�������B�d ::��:�Y�ҵyH�kk<)�ƫ��!�-���a$��T+	�@��pIS�\�"�tgF֠���j����k����o��o�ר�.����Ԫ>��a��2�w[�ty�>�Kٌ�^�~5���/��8J)�f�;f���l�a�����V���M	�	Bwn6�(+=Io1uܕ�[��B���ƅ��E+�S�9�ʃ!��d(jy�OTNt�&�_]��V���=BmOq���1ޞ�1�z�`����m���~!|��T��ui./_O@�,#��X)�gC栯]�����Y+}�ܝ�x�s=2�n��������Dnߨ����*"�;#YEO7�]�ƥ���랧|wf*��=;���}7�zoՊi�fp��R��yZ���`���h�m�t�]/7+�Bi�^�y�\Dj0�k����1o82�.O7�U/.'�*�
�R����G�LY'R��S���דӅ��������ق-]���&��:����[�m]�Ӻ����m�ښ�9�����ˬ��O1ۚ����7���(>kd�M~>�Y��ܨp�S�Pso��>+���b���Z�FV�}�;{/:���睊�Gs�yյ�lV���\x�R~�9�+�W�q� �+���^S���R�����]�Q��{�f9;~����c�w��ա>�N��
���-�a=e�o��]�Q���^�z��or��G��\����&-*c(筪�0�0\�LuX{�%����*��CU"'�}�wg5fߠJ�B������f�\��U��s7G���1n�	f,Tz1׀בvY��ӵ5��<�:AЭ*�:����M��G����6��ݪK�y\4$'3v�k둄=o��H����Z?=j�6����
�P��8�ާ;��5��w+査��mS��VA�{[�Ⱥ�𜂘|�,�S��_S���S7�!Efxu:�uw�S��� 1��ᲀQ	6k��g���;�!=>I-�WOʯ%��Z�l��e�5��^�kn�G�t2���vh\"ƓM3Q���8�,�+��������c�C�)f��k�j�j�ƈ��P��..Xs��Vh_���,`�Cc��l�/��즸�ոő�ʗu�$�͛��il�M�2�.�R���In�p�z����}j\R���A�.��3M��IiZDn$e��ݺ�����; ou�b��E���L��#����Hiwη�ʷ#�8>��r�I�[u�KC�q���ˆ�u�;�4��_{���U�ɴk7xV���,UY�CFD�����P*0�LZ�c-��Ǯ��B�@q�-z�*w��s��i�C�plVt�~��B��O
�.f� TaА7�Pu�Z�6l�啴�=�w��OCA^]�&X]�ՙηZ��cCa�e�-��ZP�GDڦJ�,2f�b��4��V�ע�#a�-M`�/����tXl��ݠ�|��V+��7�R��r�xE,#F��y��*<�{ޱ��*��p Ҹ;�k����/Q� 1�*�A�<�2���x�fR�K��W�6v5ʮ'�ʛg��1^�����R��'���`1L���>�ֿR�L)�o_��*.!jh� B��1��ꅵ=}7�a��xmcr��̮�/!W������G����HѢ�/
a�\P�|<�Ù���s�ى�n�$!�#z:s{��¥ʖW���T\/��ۤ+NA�Z*�p4�+>5�����u���:���v�ۇ6e�����xQ���N����i>
jV{��a:��:�40��6u{ɑ�}7�nf�V�$�WK��7V)L�zj��;��ư���q�wB�R�0>�I��z��v�L�eg'�(��_Z[����ͫ�ab��f���eo?ng��V�:vf%����� C��`
��W�]S�%dz����˽f	{W�5�sv[|��� �;�M�_G�ѵZ�OU2�z��Qyb~(h3ݸ�}��
�R�Ҧj�o�^�t^|�G�V���茋u��7��+��b��	[��3
��a7�'���S�!�"gB�\���s��uػ�Z]���y���~5�*���l�J����"�99�md�ʽv��dƅO���y58����q���ȭ�ռ+}��O� �z��G����餆���8��Ӕ�yg3��D-pm����1�5�k��PN�=Q�\l;������4��f�й���:�y��2��qW�U���K����*�Z)��D�����p�5oе�R�����rv8�e���p��W���.���0%�t��Re����;@uu`��'�K�9CG�λߜ�y�ngX�m_��]Ʋ��a��gzO
�#k	�&e/5�k���˜�e����Q��5�R�<}h1sʘ�3�R�%z�x>��2�1��=Y:s}���amY�ë������P��t���t�b��3��(s*�~������e��.
�_:n��
,��L��p���Sꆋ�ȳvq�娊���u����}����:�jVc�Vuu*�4�cټ�f�ܠ�.*p�$�^�h����Wg[|�lƟhW�+)�Yˤ���Wv)+i����{�rn-�)Y���q���n�­U!2H��Ij ��3o�|�V�o��Uh�����90�x�4�D�=�s�	E��
X�_M�W=�i��ٷ��3�םos�=G0�^�N�Me�B�����`�&6&�^��*p\2�q�=�x�����WV��-ݞ颊7&5�C�Ul߂�C Zq:&@���(�a�et��Vn�[�"������<IȒ6|;<+Lxl���uGKe�����	*��S&O�]��v���Y�8h�ų-�_�F���T��<oF�L�K��U�w��5=X�_o6}��\�z=�pc�0�"9ØXv�X�5�ܤ6̲��	pj�8���M�yL���P{��;U{3J�M*����xֲ�.�>�7n��(����Λ�<�9�]պ��)nm؊�l�*ݩ��d�=X�4�x�	��*�/>L��D��j8Y�ʴ���Ð�3%�T�z�����4%��ky�	ۈ�dX�^mm��=N�r�<uj�ɀ�4@m`�q��~��eݏ`t)\h= l��1t��5o��$��Ⱦ��x�o��}�5n�O����]d��hw�m�|r:�GPS�7U�f=�Q�\ݷ�`��w)9}i��wOyν���`J���F�6�E�ꐖ�9��z#б'��s�UZ"����'6\�(#J�hƳ��:�rs%(NJ�6���E���O��sĶ�N6��.�w�x_����өևU�V����+<Q�\�GV�ўe���d��3�5�9����ԋ��7��<���L�����씁�x�����Z�*�\��������IK���3c������R+���5����A��_.��9�#��5̫�I�ݬ��l�,+�g���D�T�^�+�Tx��;"T�UH\K�E�c��뀣{����6��#rwȍ�`;�|��٩.�t�ъ���u�x����dFE�K�VE�Ѿ(])�7�׼�
JX�.-��1p�2���ef��ޓA���Ou�♽"�Uw$=�*"���Ȣ��\��*m�I�����?���K1͇(T�o��o>y��V}�D�?0��e#���;��%?:�Z��]��$�N�˕���-�����R��˭+�B��� ^�rx!X�D]P��xg��G��o���w�17�����U}���(�!B��X�[�w����Q5�(ySooEYRҥGݞ�`וh������nRĴ���3�Xah�#���b�JB����g]Fk8�f6��>�Z��a��煌�v
�|��_L�r��v�rx��;�W>��Z�(��*�1S��PJ��慰g�%�58��Y\~=��D
S:�noVO$�v-��2A���
�X�d��h=,L̉��Rz���}W�J.�sԻ;�e�<�DTt��eѡ��MD4&,N�'ae��9���VP/W嶱����<��*sn7&a���p3�q�h�<�s��k����,�M������+/�w?r1�`��#��*�ݾ�4_��TTf�(�:�1��n������@��a�'<K��jBα7Ռ1�s׸�d��cA�Շ����ŜE|P|��z�q���*���c��b�}�ηZ}j��/
�_��a�OS0_�����|�u���me�'|��!��?l���0����Ƨ�Ýl\Xt<<�Д��OR�s�JWhVI1�N5Mb�M����	�^�����j��`�e�mOQpkj�m*��Z4Qbw���<w5(��UQ�g�c��q�e�Z�?[޴��^�ڍ�����#/ղ��;Z��*Ԇw\�Hv�ózN��w�q��q^D�]��ʗ��՚�b-ب�
�Y�%�dG�z77e���D9�t��#U�<絺��w9�/��l�*�2��t��?+�
�)�x���|mv�h������K�S��#n��=EW1���c��sCoY�w�O-b�ߣ�w���L�����+G��w�]ҷ ���˽%@�l%۵� ��R���n	��v�(c5$���,v�ͷ,���9j٘�ĵ
��ea� ���_V�ug:΋9�/�H�0��zj22�4�s��9�ۭ9�%J���J�H�@�g����]jt�dX�%.��ˇ��]��ǽ��0�m��J{��E"����T��J���l�땸�1�7��r�3��}���}��NR\�w�5L�Y/
�����6���9"��j� � �]�B�p],��.����h�5+($��=*������k6�KV�\{��ec���D�����T�ɄSr�#s:��8㚁W�s<���[��^rAn����N��)i�Q@sC��%
{rU����>��u�;X+w�}��Qu��%����cC���4��渳��EꫫH���aO���z����U��۸�'7]�[)K嚀_Mà�P�F��[���切����3���(���"4���4�{����<��Vҡ�����˔��1va$������+�M�zo]*�0��e�E�����qc�� ]�%����cӸ�L�;6 ���R���H91�Yu��u|(�9gJ捭�f�u��d���/%9��Y�X�;��E��M��/���*k=F��V_L��C��on�(ӷNZ�ye�ڼ�0�o��9�fB��M\������LƝ�ݮơ�7��q71Y��F����;PIJ'�.:5*�)!Ǎ�9n����WR��Y����Y����A�{ٕ�PRe��A���6;YӪ��2�ia��8��wZpeS�-F4�u���Pq�a8�ئ�<��]v��v�ª�u���e�jLL�&E�-�p�y�;�Vjsų3������[E�ň����
� �u��!�u �,�Ge���*�Emv�VZ��eZ��/���c��U��u�=����RZ�"i>��j�ueq]C�uྰ�Y���y��E���r�R�GUc����)�78����=�^۷��uw�Н��F��`�T݂g�Lb�޼���#�8�^u���,gT�P����-���OXs����ٰ����1eZZ�TF��F�Iʴ�ޮ{,�'p�PӍffF���1��X���R=�v���//n�#�>��uM��8�=���/�ͷ]]�ƻ[8�Ǭ�=�7.e��Y�XVN3U�j�k:��I��m�.7��XX^�.���.�a�ydp�O8�q�M��c��m�U��4��0s���1��B�k��,%���*C�M������ܣ�AW�ả=3�{)2e�3Ԭ�y�#��u0( |M��YP����Ńҫ��Tb"�lFE"�X�,+
��Q`���b��D�"�-�c�iT"�-
��������*�%�1*�#��E�̘��� �m�l���(��AA��XQ��1-����P���AV��(UTEH�T��Ke@QdTdc1*bIT@���l1�b��1�̰\Am�A���LEP�V8�f2Q���R�TT�*�J�kH��"�ĕ�����*Z�0PX��R�`1A��VTRT�W�A�	�U�2.Z
��R�+�aD�)X�#Y+�#lRV�*ER)�Qm��X����@D���2,���,��W(LI�(�����>͛^~��/�	j�i�`:�
�ym�w�yto^���*W�k�*�Ɣw3�\r��fab]%*ʚ[��Wg�����N��DP�}{5����
��왲�Vj�z���m�d�G�ːuro#��(���г)+����x�>��<MzJa��HP�E�u=�ICm�B8�X���<�sqUպҼ�ڛW]VN٘���Ⱦ���I�<�<6��H��b��׬�*7���{ȖvjL�L��A�R�
������ȅı^����a9���7K��`�K[ʇ 𪂆vz�
X�1`U,K��N������j�3|�o��k�e�z[���Wa<Z*+���P�y�AA�B��w��N	%�#!NT�h���pVt$�[�����ks�f�^3�U^����v#��H�͓�МC���n����[��b1��dehpOY��e1���鍳.a�P��R����}�]�݆w~�	�a�_G����
N�k1�5�Z/*T�Î�� y�3�i>xܼ��=���M4��O<�w8!VW��\2
;f�,��{`4�:�]�~H�E
�{p�T��Wd���9k���b��� 2��Y@����>��#�����X.r��FR�iA^���zFݚO)�J,r��<z��^Wt�2b1+7ȥ2��8����A���ң�0oe����-6�j�)m?�Oz���A�}?r�`���B��=�Pf�芇��[�xxd>u�k.X�;~t�t��R�u��MԔ�譹�w�ыӰQ�,���c:A��c5�|2:�ȶ%�q.�:m3��7dS]���;�W�O�ؘB�`�Tb�M{�� �c�XƓ��W	���mx�u� ���~�2�߶0fy`�}u�$+C��B��NO�<:j��U���������EG+k�f4C���J$��^va��j4�*@�T)�r K+֪�"G�S�]�aa�Vm�Bۜ���RGk3�i^Qp�f�%�/L*Z)@��!��s���+��bWaW��J�l�&��l==�ߋ��cWz+"�!s�0�=a�Q�cp�.�_bq��CP�uH��G�;�y�s|�I���P·R�ٰ�������V튳C�+��Ù�ٺ�&��G�N�z_-Þ�́a��+(�{�t�1U��	��l�e�d	�]S�r�+<a�(���Nܷhx Cql�rX�9{(Tf�V΀Ln��L�8�W�����ׅ�J�J�;��"�8łӒ���-�Ome=(�wxU�&uZھxkj���|���Ӽ��A�z�ѵC��*��N��P��!O��U��:r�m�R���9�Y1��ix$�ќo6�55%��_gu��v��-QK�l֠sx�w�Mo;��r
�C+��(�N�wS�[�M(�Ha���i���;j����,-~���X�u�[g%S^�S.p��e�q�$��c���&5scbk��]>Y%.���m��;��Ҟ	�ļkYw����68@����P�Yc-�s=~�Q����!+� ��+7����׹�m_��Y�1�*���#xh�U"Y�8�8a4��8}��HVf�ht
"� �K�[��G�Y9f��!;Έ"�OI�z��,g���3�m�M���
��Te���A�XyLk:.=B��%z���1��/3�a�����ԋ���=��w�lc��ڀ��Q��]��7����V;Caq�=���*6�z�p�/��w�N���7-U���Cz-��rud�F�3��d�>Է�����y��E��dx����Ӟe��b�Q�(R�q<���D�*.X�-�J�ً�'��y��q�������G|�Q5Yb�O@V�������y���M$�{7��mu<,EF)x{#U �Z�Cf�zν.�H�ԼF�[��(vu$�,5:�aT;[����б+oN:���{$5e�Y�湞�Wp�T~��b1P�n6��l<{���Q����L�v��oh���+�܋�aJ�hN�;�^�zJ,�S�Z��֊��ա,KOW�ח��tm�~���
+�a�0����J̡U�ix�=��t#X`�-�s�6d�f��Y�q�a�&���z-��0�ط,lS��#�PG��XXK�5�>5�l�>\6���߱/eK���
��n�6߂59˖l�Z����i��,>t*��@�}+�oB�(��Xূ�z� �a�i��Mv�&)�y8��F���F��""u�7�*�0�衢������U�!��l�M;���n[����q{B��@:0�)
X)�jtD��P�5��DL�͗/�ȵ���y���1�ŝ���$8��l�4.��a/��P'Y�U[�C�������M��e�4|3x�M�in�
͙P72��bÞ�k��l���P]����c�j��Z��Z���yƤ=�[[X����o���u�lw���a��
r�q���U8Vg%to�+�I6	���'�����cF����ܸ��t$
rc����wpX&�}n�lMTmA�g��)Vj������:�K�Gs�i*ʞu� �����¢��C�V��Iw(DoH���Q���E��;�s����g�_j���Ks������hN|��vqj �;8�*V����f����[���14����W.��wV�q�X?����u���ef5*w:[)xT�|u�ͽL?�R��&J���j�f�,�Ŏ�s���!��f��h���ݩ��G\�Q��xy��)��k/U$���������Xqjt�/ڧ�k�,_��Jv�!�
Z����K��lJ��a��zM�\1O9>�]�ʢ�2a�3��P�F��7:�N@�z�m��*�K�<����ɬJM;
�7Wt컠ƀ �0�����\7<a�[��4�+ϕT�����Z�7+�����Ӽ7��4��Uv�b���$1��xJB�	��mK⧳f䡸�S̓��P:��ܻ+����^7H:z�
�U�֢��
^�t��������X�	j���{w9��[
M�t-��9Qb���a:���>O��Ꟗ��^����nӟHy�����{Cʘ:P���0��%�S 1`	�R�׺�T;�f*��.Ǒ]y��WgcQy�N�Њ�ʋG=�Iu�%
)�|�pI�KEz L.���vT���v�sA�,j��>S3~����C]Q)�q/�d��x�S���:�A�O:�_z:t�V(2���͋�����c�n��q͙v�[��3�WTa��-o4����a���e�~��&]]uS��pOe[d�w��WB�B���]7���g�%�r�k��5�Ymׄ�Ő�a�f{\T����wz3U>:E!"��|ev.�v�g���ׂ�X�dV׫)�鋍�p*4؇1a-R�oXK�r>�za�]����[�o�]��tu�"�P�!��,�7�8�A
aa�F[�0(�[�Չ� �6��F��\���A���
�jV���.]����7\��TV�KK{B����S�{��7�X"}�i������λ�d[���@^}3+�'
USE�2f[\��嬥��!|�V��Ry�Ǻ�a%Ղ��Wq���%B`�(���~��C�s���8��fR�t��R����@L��H��)CC��u���3|����C���&ioZŧ�>/�=���).�B�:]��J(zr���2�L<�[r��G�K�I�^���pк��by�Lq2�*�q,K��0�	c��6M
�S�Z���Ϯn��$��[��b��f�q��6�C0�����A��h��P[�4��8.������&��h՞��)^r�"[�z���i'|yT�,&z�D��Ŏ���jvúy�}ԡ�̖���Vߟ�Ԃ�h{����`�\����-��(,�B�Q�;)�ћز�W]��$	ۡ��seRgB�gCVLh����x �@���׾�V���e��Ɂm~��	�רw[�)����Esz����$�׎.=p)*sx/;�]��뷽���gl�bx�=�)��7W��-�0n��T?s�tt��]zK�����2t$�˗B�9�h�(lF��(h{�ٸ��qI։�R��!�q�=335��~�Y�Oիf<;|��)������uj��hg�N@��	<�>�~n��]q��+�o3�3�N�B�`�#���h�S	��<oF�ƍ�sյ�׃�.*�=�����t=yJ�/]x����*��w�l7�xZ5{�����/#� K��j�s��WY���j� ����u�=��2M{�I�p�]�<�-/��8@���<W#�K�ݫ�Fu�빒�L�h�+�]�z<�Xy��b��ݩȎr�xnEy�řW���^fz�:��{�}�X����l�p/rXf�
�:������`�~I����)�r��bٙ4A�N�$�[���!�3�\:+b^�V/��T�|țT�2��u������)�'ݏzr�F?&
\��z�q�ߏ�j��L���Q
�!^��z3�8�t}�6�Q���՟z���P��\�`:|T,���غ�5����D���靹i���o��s���Rl���f�A��_g�mԱ|rg6p���uŷ)�o;v�SJ�}�Zj$��r�P���o��_& ]W�����cb.\W�d�H�:qt�z�H���#�Z���0�����¦G\�KI�427�(`�2�˔Jުg��]�T�U�M�]�(Xy��V{e�E�v��t�;�Q5�!�f�����	�UY�W�;�ֹ�Gv��	rXphB����P�7�]���njK�@��5��&b:M�gH]&�����jNvUn_^�Xk��H4�O��R��d�����ٹ�p*����v7���RN��}8��ǩ!�V|3��2��ru��6d�n/SƳK��lŦ����FL^�=9����
�*S��\W��׍��*w��C�R>\r��;k�f�j]�Xu��on��-�;�͝�ڥA�҄T\�@~ޗ�b��)�߄� L>�ބ)��"��S�d<m:�ӏ�S�m`f��A���ԑrBn����Dޗ�dp�7J|t��J��5�s�qj���(`�o �QN@S0�*���"��7 � �禣Ҹ��xD'�:�[��B��	��9���XpV�鳅�a�y�ogw��-2��6[��c�v�X`�����^����p��x ��i�,�\ÊO>��l^DֹQ�� ��5�]Ҵ.W�.v��O�%����=
w��1�yY-�v�6����U��x����:�n��0e%�b����]�R*6��,�k�/1�/�c�u壥��_��β}mׅ<ڥ��.Py��Vh-s�P�1Q0%I�i��fy���y auz��ǶnN��,`YN**"sj�4�7bW��:����똛�c�'����4};<
{^�v�'Qѕ<�A�����U��[T�����ϥobH��\iAR�y��zo�UGuNZډ�"�Թ�m�z��GC�'���o���~��I'����J��J��ha�Os���q���ܻ�1��B�ã�,�T:�K�]����B��}JQ</\�7�X����U��򖯨��#(@c��4�"2�徑�G���ں�P�}]5r�B�N3���{��{҇9u�\wc�&�7�f�+��k1J���������������^�������|����1y��%��*�I�nGs�"��V��?�R�u�IuX�ġ+ǥ
��XwS�u�ׇA�~&�]�h�ǻ;Kbh�∽��>�����>㵷�/��_�A�c�o���I��T��qe2�gFjdǪ���¬u�,m��xB�v.���VL*�5���_xFDO�+T���Q�� �u���ΡSUԠ��!8Y��>37.�]Y���N����q��z��Haɘ�WP�� ��t֓>��Y��D�\=��O����ۄ��xt��qp�7�s���.b���|�(�u�x'�']7��>�5��ZJ�Ef�ws�f���b�`i�Q
��1;N�����q� �"��Bj̪����-�f���mm����-S��V�L��-����}�=C@�P��0"o���u9�3���>��q!cՈ7���9mp����\�1�����*C�����6x��}�=� 0G������x*�B;�=�8k).X�2��i�/�c�Y�9wwof>��K�i���]���L��R"�pd!�W�ҩ,_�G�_!�6&�+|�N�ǵ8^��p}�¯v�����e�ѷR��*5��*4�1Xnd��q厠�M�{|��X��t;��{I燬�څg�z;���=u�SH��rY�$b����O�;}�\�&㔇��X����P�>�(���c:AӪ�5�Z��5Q��5`�4f�R��6�%��Ê�m��;Ycώb�6�E�39�^I|��������3�����ub}ফ�n��ʑ�:[���5γdi���]{J�y�7��Au�V�!k�h#�9e�x���η�N��0'x��\r:5�z6=8dz2�E���
6�j�H7�(ho��l�[�(in��L/vvۃ�=�v0v�ë��)��~�DQFY�D篢]�����V�",Ρ�F��)r98��4�u-V��Xmn��tL�+���A�B�\�DY�� \���+B�烒I*���+ƌUoS��֮y������,�Se�U�5�E�3:G���5d�J���1�`�N��F�5x���[���� %�^��F6����#})=em�2}
��فv�����f��u]�Y�E���{�2ai]��=w��rwć��l���'gXf�ʴ��� ��Y��s��p1��A�L{r٭���{w6�ꆉ�g����<3w+G*z��/�)1LюV����
�:�+Oקje��)F���h9�d���gnW����跴=6j�EF�a�pQ�D}o�n��W,r����t�o��f,�*AaWj�>|*�*�:��Y�qٝ��P�bU�mC�Ѩ��L������N�۬4([�h�m����PYW��h�l�r2�R��s7Oz��d�阖��hJ��J�K��s��>7��Gr��*ﳃiT. $�y���\3$���V�[+T��ދz�����j�i7HD1MU
ښ=�5p���ۍ��]�����ck8OKí������7�c��3�E�o��ƕ�)5KGf4��G��j���H���Z+Iܘ�>D��q��3-(�S�V��
{d�Y�U�Va�@�6�8�8���I�R�sD��ܢ�zev�JY���(��_�ז�v�tIt"	�YP
aD˚2��vWi4���N@��4�7iZ6�R|�ƹ#}7��Dm)�����r��9_Rtk(#x㉊�o*/n�"u�-��J����:�4���s$��>�(���m��t����=ڰ]LQ�����H��,U�;W�mQ��3/h�Xno,��7c���6�1��w+�9M�*��p7��.��M�������e����Ł��\�d����wsNP����%�vR�R��l_
�kN��}ޠ��9,��4��o��p�<	}&�J��ٺ����*\AȺ�Ma���f���U���������k0.s+^�˻4f)��]L��w��m]˘� ��į�Q}Q�֬h��+o���:�fjغ���7{�J�g�����'��d�Gt%b;�l��;Ǌ����`U��*�h�����]������X��Úٖ���C \�i=7s%���bи�t�t�0����y7ff
�[�.)6|���e(+M|�@j,8��t�`��wVq4�X�`�n�����|��}��u����ߘ�R)�JZRz�AFڂ��UY*�b��EX�B��H�jUB#(,Lj�J��J��011U��PE#�+�V(�2��l�AT�E��DX娱A�fU�VLj��`��
�*�2�i
��2����X��I�d,U�#k[,q�*��TX��L�d�D��c��,*V�1r�X\��+%A��5Um̪���bTR��Kl�.P�,(��娱TV��F���G���"	�ڢ�AV#Re*���Պ��(fW32
T.X��+m"�"ʔV(Q.e����Q�V���թR�6ю]�i�V^sm��N�,h�OqMrQ7�{�;�\mT��U������,L��Z�uD!Տ�]oI6B�1��c<���`��#��sĺ�����N�P�Цߕ��V���<�;g$v�-�r�80}X��G�8w�`�W�)Z%)���\��gT��tQ�����yݭ�f+9P�~�,L�,�؞�W�t��D�d��+�B�0�MF��Z�\�IXk&�z���0�tLK���
g��yƣ���R,J�E:CN,`D���C��Y.k;�۩Z�nf0n�RLZכE�Ra�z�Ѹ~0�	��cI�8,Nj�ӡ����r+r'��9AY)-����;�+�^��[�.`����&B�:2%�Nʌ+�y��:밗�ӂ��_�a𕆯�����r��1t%U'Z&.�v�)�����iۼYo�CgE_��i5Μx�Jg��C
�,w��1U��M����:��r[o��w_��3jn��C��<ql�,S�\\`ʋמPОA%۳U0��=4���L򮭤���~����~��0�]�m�^����d)���Į2�d�r�س ���~Ԣ�k�w�%�J�K|<9b^:�ȻK^!�C�G�Z:�0^˵��l�>^k��\�3�w�3B�@c.��m������nV�@L�G��,�:�A��3o�j�B�v���
k��,�E�n�bz�5X)ຉeRw#o�%e����墉J��X_�&�E�ֆa��mP��J���4���u&u��`fυe,�
y�Y��6^�yMu`��PP2��U��.�f��`�imn�:1vP�/�7(40����s��c�D�;�9Gh�B;n�����\
�͔�ס��p<sb �z��y{�$Ʃ)��}';�=�z�}�Ƒ����)��#�EO�9{�\�c
��ܾ*��Vև~q�����t��H)fR�82��}=KC��k��p"�7EZ��Z��K^%<5l�9����l+M�2�o��G_���%M��C�[�@T�;�AkZ�l���W˜#V�j��f(p�[�e�A��@����Q5�!�D�] q\r "l�\7��,��jZ��{�Rg���0���u	3U ��,4:�7%��w�DT#�g�](��GSw'��|���W�����/��O����t�3�W���T�~G"ګT��٥���O�fRW��!�����\Y�O�T��D��x�2M�-��Q5/���9���i��\���g���f
a� 8.�\���I<¬i��#@��[d�i+-�=�y���i�+��؇�<�$lCV����:�K%)Qq���Py�#�@jt%އ|c�����:�^�y>�飛/�(�fΜ��f.�~�摕ە��2�{
�*��(qƫ�.7�C������g��B��o�;��)Yw�𧣷M��1���U1~D��O	�*nMD*).���}��E��'���v��)�C�b�sRE�5�\��L�ȵ��Gҵyqں.�g7���'�N�(�o �Q^R�� ���*�R�[�[�2�Ŷ�pK廛��x���5�[x��Vd�S�ٌ�r	+� )��vh ��hLX�s+`TM�t��2�ie��[�*!�h^zgsfq�f�*���ڥ|1�89�����ee�.�
����;%�`�A"�l5���nN�ط,h�q1xa@�: ,���a��3���K�s�r��ܺ٘G���~�{>�>[�o����V����[� �$����e].{� ��x&@A��p�Ňz��zWtN���S��^[�oS>����93����W���=S��xx���
�OJ��y�G�@l���
kv�\X�]μ<�';��d%�%������ފy��s����+�t��-cK�Sݏ��Y1m�N��gه�ݫ�jv�M&�{Yewbw�^7έ��o����Y9��̼�B�m<��{R�#0+9*��q�l�ڧ]ȶyq�'w�Ae��Y9'Z�m�O.i�<[9��`�C�q^՗[�î�J�8΢�á�)}}E�#(Y�F�$�E�����s�{�g���9��b����\J�q���cW:��{քߕWf�D�0����%8f�4��*�I�\ �U���0�DU3�<z�kڦ�QA�]��f��ԓ]U���F�ni��7�Q�a�(k:OR��P�҅xm���K��o�e:NM.ޣ�&x,s��3�n�$_�˳1p��I�Bb%���;6�iȧ:/��_��Ǣ��)M,�90��Bt;���p��1<����M�`R,�T*�\{��K�m;��s��=|�g_+	����f�����Ӏ�)c \2� �&f]��
x�'����[�F�U�ks�Jzn��M�1��ʋG@%��H3
\sd����E���tݹP�9TO	/�x@�[h�U�7���9�b�y�ux�xJ�l�MT<wM5�:[|�l�t���M	��u��r�= !|=x>C+C�	�ù����S�.7&�b�K����9:SJj2�wM酃����˒�R�/(�6j
Y/��+ʱ���,5Rl��8���4��n?rt���$]4��o V�[�7���5��V��CCs������9q;�`Ql�����2�2��� �J��M<y|d]���)׾yDM���*��;�C�ضg��D[��:^:J���.������{����Pqࢲx0q��UƮ��*Oʜ�t��Q
���Q�uY�<$+_t>����g%6\^�!�z�l�ɿoK۬1�i������t��X�Ջc�*sEZ�i��b�&�8�۸�rU���N�Z���|냯*���[W�Jڋ]�hm\�׹ϗB̽�+��z)q.����tH�V��huC�k��|K��7(1�sHD������V��m�3MƦ�ʐ�
�BT�X��(e�"�*]��J5���v�+n��o'��x�w�_[/�Øs�P�SԄK�5MBЩ�bT
��!�<%�����s;<��%�ޮ�k�N�W8<=q��ڌ\�h�L0�K�P�LT+��[���}�J��W�m�[w}�,[���ib��-�ĥ��tr��}���¦�az ��{ݮ{�r`3��쫽���4YXK�.p]/�����Q��%U�q#C ]'Z'�PuY
p��r"��{�h�s�l���0"�D��d>1����#s���(J��u�G,gA�$E�u�t�K����󓁛��C�9���vS�é[�nP�!�HT��Ց����Εo�ZJ�q�9�F�wTw�9H��6��Wu�0��:��|��NPe��wW)����Y+�Xm��mi����>g�?��i�k��G����vggyFIX䩴�tݙֲ����_�'�u͖xJ��EoQ��Fa�x<� MM��,yQ��m�����*���V�"{Uެ���u�B�v_��Ҽ�l䦼-�ܤ&�%�LS0䞭{o4c�)��bjqQ5	S�Zs8h���D���]#��i�`�� ���������A�)�;fC���"յB&����׹�{�{ ��{����7���Nuv$ڭ��S4�f.M�%�xd*���5б�3�hמ����{C�^��A�J�n2��y�ý�ݮCR�V&�!�3��xV���
t/��^$�XyLk:�,]=������G�W}��0����Y+}�{����rz�p���:���o��,��%�����g,N�X����������A�����\�ʕIp��z���h����A�@�s�ڤ�V�VM�}>��5��I]��#Q��G%a��V6	B�G���.� 4��r�e�sQku���f��<�*e)�]8�k(WN��#���zH�Sfhw&�� Ǫ�v�[hv]����m>t���v�;z�3ۻ�Y��=��9kiӺ��Ǫ�K	��J��'s���)r�cy���S-�C:M�+�ǵ�p�/�<J�mTXb�E�d���UMn��%�>1
�
p�Q|wV�ov�7 ��j���sh���,EF)X{#e��a�����t��3���غ��f��o��Z�P��plG@���]��A/����X�o�m:�vyP)*c(��#�[�LS���\���L<�O�
C�=`ϒ^��j�
�l��M[Y�/K���¦>l���z-���ד�1����5಼�#����]R�����.P�_	�F�c�6����ڬ�qN�Q:鈗3P3�K�1q���Yk�WQ�}>V�!N�(�W�t�e=Tp��>kKt�C�,:��V�oT�Ɲڈ����$�=AX�܀�ѷ�I����EohC��=_��B��A�f���>�TT�̴��o.�HAe��c{�GzNޘr�O�Go񬼫u8�b3��!�Dt������X�y�F���unr����T���/2�3��*9��wN��V:��ʨb+6�@�Ì���Ks�Ey(���՜�v�U��_Nr��N�mio)�5�t諲���5�k.��K��r����t,U�m�r3;�d�\����(!�]q,�Ǳ�IW����"8!��r԰������q�t	��F܂�̫�뛆#����f�����r�L�z,W���;��8�q���"�����6k�'��ٗT�矆	o���*�s��]�w;�ĦdU�1�g�9T�q]o]&�5g�-��m�>���0:�Ր4Q�<��#35/y���vz���d  �`�"��Z�7�n!��ȶ��,��R��u�w��{=��Mf���u��^]�R�(�Q��&��XX��7,&��<0&wjn-�Q�Z���#{�sv�{K)`���,u�rVPxm�D�z���,X��t*���-V�}f,��Cg|J��|����!6�C����L\
��9��\J�m��,odr�>�l�8�<��Y�&����7]��`p\��q����0�@��p 5U\ˮY�r��f �<��tI�������=N5Ս�L�D=]�K,ӕfT9bGy��b���jK0ؔ"�U��R�|2a�[�|s�I��Ӿ��,n9�G��j�$Kr(�j�D�&"X�z%�Q6�i7n��,0�Tٮ|���G�>Pf��A^/4g�����׋�n)K`R�biP���c �L˔Bκq�yt���)�2��룁"*Ifd}wO��;tbc(�߽<���(��/�1K��=1������	�Z-�׍����,�p�xu�얅������e���M���RT�ܨ�vpֱ�(qɶ�X���7�>������Ǜ���H�#�՜�m��5�j����>,Z��
��Qp=�K�0 �ruV�$�i�eG^.���	�5�	v����j�ʭ9�׹Qh���k�A�B��X����w���9�`G��
U���A�a-�V�L�K�Mxe�g�B?��u���8�����	���ʸ�`>��
2t;�	�ùYHh�r�tw\Ә�m��[)�{Y���NqP�,:��W�֓�a��o��HʍB��Fid�o�A��Qr��}+m�u����a�:񃖨{�=CG�\ڏ��_N��������[��62.s|�S;��Ն�U�M.��.Fl�ɿoK�:��i�ȇ����>u�j�F��L��n�um.X�
�l	f�R�IHDu�C�+�??P�q�Q5��Ʋ�s4!Oy΍�1r�����*��)r;����İ���'�d��Jp�	�X�Q�P�ݕ�8�Y��8R}��2v�:FM��S1�n5*Bo����P� '(dl�Q萭v�\Kyq���i>"]Q����.���MK��vΊ�P���v4�7!�+��JV[�Ґ5�S��+�}�iLk��7Ľ�V�>L?9m��;"�`��%��9+��|e��{�u7��dD�*r@�5�ˍ
����Bn�;�	UӨl\4ߕ�bs�P��,2u���ƣ��o��|S�:��=�������ޞR �ÁCF�OYw�v�T�.y�s�ã��"��)W:�he)�i�����{Z���Ƭa?x��v:X�_M�W3�t\J���x�,T-f�Mc�*`�F�ED��-z+����\�Eu+W��g����C�/�����L*�+�\�qB
�X^ݨJM&A���T%IR7�a��h"�u��чWL�>\)����i�����sW�͊��zy�QMP���	��Q��/���< ���9>������<獻,5C����V�K��f��5(�v9�@n�)�{��E2;����|q�������eZM(�Y�T�Q�)�t�.B A�N*.�h�2J�rc#�N��f�q;��]�^���]��e��Di�{L���F��lȋ���1p�%�g�J�E�;K=槽==���^`�a�	�ƕE�A�٨͚l��+}�пb�,/���^����L_��]��p3�t�;$������m���_^[fCp-Y.��D�Vw)���u,��)X��яzu�
��3���'�6,�=�KJ��w��WN;Y�;m��s�#�Y���Md<��4]Y��Ȏ�嫇�J���3r��x�Y�U�;ke=ѫ�9�"'M�ïO|J�a��w�qy��M�S:g�C�iS�V��\R�c��щ�BUŋ���C{Y��i̭�\�o�����f����Ю���]Z��*�\
X��+�G]�o��M����nݐe��Sv�t)J5��&17��_]'
��eݧK
GX�H�p���`���d�R���񊻗Z��4��>�b �e���V��V�����s+h��C����9S^y��/��w�I�k������E�CU�N[9�f#�Uw��T�i�e�;-��1業�S��G�zU�7Jp������\���]\UL�+O5��A���ڶs8V��S7�b�i�łY����toQ��Q�f��c�*ڲ���������M7��8�^��% �+V�	�����iQ+��ni=x�7�b�a�ǔ"��*P"��]�e�=�S��z���fr؈�-�6�Y��gP� ���z}����3�+K�}Y�i�r�Ū���k2����
|;4�V��W+6��/�k�ث�T��,�J�+���ì��,1X�F���"n�k+���ثi;+�T�K�yj	2,W���J=�T�^��zk����˜'JIZ���=�́���M�e�j�Nn����U�X�]����hS6�V�J��wiи^*�4GΤ��x����x�^ʻ��VJ�t�Y�: �}�/2)3��n�<T�>������]�M#s�ΐM;�L�|(���I2kh@Wu�����d!�ϲ�d�.�$!`��([�eLE6�J�#�;r���@��<�� u�R 	;l<�}��[��ԥf�*�g
�;~���?-�,˪`b�Y��8��sgR*�#]�ƒ3���p�P�N4/o.jY��V�?9bt.��RҚj�Nm����6�E̵E�Ǽ`O+�h7D8p��$�[P*v�gwhM�Xr!ssF��Zo��:G6×g庚z��h����F)� ��׺vpx曷m�i	T�͵2���s噏+!�6�:�b�j}n;"����J-[r�� cw�jc �'t}]��h��т���&q=9�ŝ&(ي���)]��u��9XC�8;G��>Ǩ��u`��f��0���[�B��HS�Wљqoa
����}���ov[�e3�d�ۣ(����|�;���*(��	�2��ݥL!{0��˹�M��zk[�H,MS �@�Mh���ҨLʻW6�����q:ٔF�i'�g�x�mbӊ������`�d�1�h�ܱF,6*��e�YwW��i�Oi�UV�[�V+�LF�B�m��2U�ZQ�rʨ)QZQb�h$��b�cj�"4UF�X�Ţ��0��E1.([B����ps,��VZ̦f5�\E�.Q��,˘-VZ�j��*�e�S��T�֡X*�a����-����F$��+Q-r�Z�-�R�,j�cKcQqr������Qm���-m�%���AQZ�a��Ʀ!�cU���X#\LE�&FT�XV� �J.8�b�Զ�����,�1iAr�Umh��J����m+YU�5���ALbʥ�Qq�
��RQUm��f6
b-Q�jE*��e��nX�K+m�m��-�Yh��kR֖�F�U��J�+j�Ym��MeΤГ��e��x�%�rưM�v�9�Ys6uj�Kn���)��$ֈ��P����Cry��>�'[1qi�c/d�֌�̒��_I�k_y`��rk���e�Q*_�ܨ��=�X\6�.��F<����u�09H!�L"�޼�����Cf�s�.�ks��C��R��z9V��pJ��$���`�ۖ�ʉ�%���U�|�+�{&UXѱ����V7=2�pxt�e�i��!T��QT�>r�bh�ڷ�g�U6�C�
c3�:)i-M�Ƶ���#wƽ��'
-�=K��3���ʰ�F)V^�Aa����4�D׃W��2�:�ė������n+T����� [������^$rK���DZ���Yynzn8�I^�\���/�
��8�(���oD\����Z�����o@��Q�,�^e�Q^�ubo�a�/h�B�D�=��5�q։�c��)�^)�D���O���ގrw�F�SoW].����{4e?���GǁĠu����K�Cط�>�ı*)^�
a<��9�J����,Bs5���/+�$T:LZ hu7\$FJCl[�}�b��*��F,�}G����}9֬��
ٖ�U��.�j��dJ�J����P��]s�v�K��i|{]�����Y:|��͟O�7y]��j5���Θ�7����ܥ�ǀ��%u8۶�9�K�u��䗞�]�E��Nv��1or产D� ոr� �\kp��P�x�N.b�!A�\�B��ns)S��]L��T΍.|g�YLD�%�2 >0�%ी"��M�2�����EU�R]�!�K3`�8�٥���[x��V:�*|\1�x�ᐠPkݴĊ³��a�%����uŐ��I;�CMLB��[��{��͙�1�UF�dY�\+��3yϽ�v��t���7��}��h A~�.��!V�c�6�u<�0K~�I�v�F���H}jsPQ��HWW��lb~�-t�����4�=2�u�*��J�o79���qT�6v��FEp�9�z�7�m���X�7��,��H�Wx���_bfHmm��'�Z������
��Uoq�e���gv�vF,o��.�e]����il�뼯��(*�r��u,j�xx0��/�
�V�&[6���k@����˫1^R�E��X5�:�Q�1G�F@�@˪����xk6�k��`ss/'���ݞ�Co���q�'"��bn��aJkGq�A����:�l h�zqŸP��EN�]a�?`*�w�nI�K��vW|�Q�4��f6�qwY���x��]�gB��H���0����T�B�j������WA��2tۉusxanr\@�Ov��;���/J�����O�kz��%��-k�����!ܪ�j��]�.Z}�MYq�;Ƽ6���ɯ'*̬���D��Zb^:qY|E�6�*X������:�P�����o�,<s�G��n�$\S�+��ãp�X�<ĺ�V���B��n��]3bb m@���X��^��o.H|�e��7��0+Φ
�:��=��y�8����ce߁�ێ����B�f+ �U�bv�P� n7�n��5���Ŗ�{���S�_��\��<U�y�������X(�ʄIu��1n]e����|��mV�x�=5Xݣ7�/
\���*��_��a�(d��3s0���Lμ܇u;��V�����j+	����qR+�3��4'׵�Hva��mp�v�tVT`ɛ�T��^��Z�h5yV���}��>��W~<��7'Q���BH�"�n��=8*�I�N�V,<��R܃i<��;#�R���}��ߊΆ�eN3�,�HTby�%HR�J�̥Jdv�_�u�y��p��-�V������tI�X�$�b��^�%�Ud�۱����|��О�S�wl����ݺ��r�ӆ�0V��c�}���-��P�1Jۥ-�
�������-Z�Rn	�5[):����s�w�ݗ��a�����DU<ׂ[]B�6Pb�z�d،�yL,����Bs��3ʡ�t�������񽢪���	�`M4ꗶJB"�u
�T���	��MF������_m��E��[t�X�j�?>u�S��bc���gA&�����*�W���S��&imw|�<]x����#��b�K�c0ߚT��S�Pɂ���H(�L��2#�P-t�v��r�� �oJs���v�5Dç<��3�
�5Ms
��K�����.�^�xO�·�+�v�tP�-Uh��#��z���@:�I�Q�L1Gd�[b�ewZo��WW��r�̡���(��8�d�t���/Y���N�L-�0Y�.c{2�S�o���%b�:pR�.����ل�V$����j���;����;O����o2��d�&��>���bƾ)����c\PT�ۀU����|�lV�]��6����=���8�wb�/�i��x���	����$Q�c��ޣ��&;Z:��x��Y-}�A��qz4!�Y�{���kkwH����:�a�C;X��H��Ӥi��%R��K��M�xJ4:!#��:�a\����0�
��v��S���W� -ly���^��tAv�6����D���lJڮ��u�݃Q"G�u`PI-��<�pNՓ�rN�,I��U W(�U:�	����P�h�>ʊߪ��߸R���sH֩%¹����_K��D:�TRR�jN%8$g��X�p:tL�4�.wsǽ� �H��0p���7���X�0���0�]��N��h����vf�H�L�^�;$ ���PxE���+F�E�M΂:����t���U���=z�v?Yg��B�j=�oZ�U]΍�� �U���q�P�S'�TǨjy�Ԩ��eC�ݚ�p~N=�TmzO)5�^�gRxںڿv�[:*��Tp���Btz��3i^�4��3�8Lr(��A��]�a�犽�*�h��&�ߥ����0T��ya���Q��Ǫr������8��Uk���-t�����עxWq���y��q�W˜u��.����/�X�S�J�8o��,/b#aи�4ʅ2�����v��WNjK�H� �㓺vF�Ū�(>�B�W�J���T�}kO�:�!���s�����|���>�N�q�U�XJ�z��s���Z��R�W���갭/>�K��G�gX�'�gʔӀԺ�ܨ�[��+��y�#'xŸ�ϕ%1|��ٽ�WX��A��AC�l�[Br¹G���Y�sz����>Bg>�3_@-kKy���|V�j�>.������%�!V[j����e�GF�\���V���gnf�4��s4�E�tn/�X�S�`!u��{�l)�Ch���0/Ⲷ@,�U;=*1�]��K�����1p���9�n�L[�bj�#�t��N��=��qFk��5���2�����ʬ���f�r���W�?s��/y�]�|���5=��XU�6�-QB�SB�eY�]o���z�zP����{��=�na=��]���[�F[��SYCF��)���x>3�	�C�j�P�9xA�t����6�e��1 �D����˰�+�2iKg�fY��b��R[1`�@b���:�X���w��׹bB�]�j������)���z�	u�Fy��,�
7}A�_����sC�R��xͺ�S�B;��~��.{@�f�ZS��V�-��}�F߱z�Ƌ}/�Ʈ�k��\���q�0�VlWT[4����i��\&ృ�X�1k��T�c�bx�]��ХlZ�����5	��r�UsҶ
��y�X#��VJTwv��8�#���n��j���Jy�k�L��Ԝ�ݭA�wK�w	�	C�{�\�q�3\/��(���{�BA�i��]��9�+���z����K�fΗ�.:	��\��kv�#�{<*&����0$�0y��]d���u�֩z���Q�y�yx�c$b2|�U�O
�,-,2{��
�e�|����U���6�^^��SV2c���á�������X��xL~~��F��P���QUl�&{�DYy��O:����d6���1G�F@���2�o�դ��m�	�Ǧ{�m\�֛W�I"��eNp�U����U/`��c�"t�i&��t���Y/Wo�h�Ws�J����7�?V�=���ן?�@��uMCS�e�������xd�qF�877j�R{whd�2���x4rZ�#����ߍ_��!�OɃN��B�P��c\e��v�jrmV�=9y��ܢ���z0Z�%^	�V:Q�Yf�m���<���f���xU�sԋRD�>w<�J�7�Ux������~�nq���:3*Y��~ny�D�;F\�I;G2���0Xd�.�瑘����-Q�U�S'�;�O��ȒϢ)N$��P�B��Zlu���^�1-���߻��GsL�g�rJ`o]��;=�Z�:@}�~ɧ�f�9-��ռ�����GT��Y���;�{����ķJ�����m�*��*�z���l�&�jM:r���tů���HH�}��E�To�>�V��pZR�$�,�z%�rx)A�v��fڬ��)�7`۶�o}z6���'3"����iތ���Ia��9R�����Ѫ��3O����=[�s�F����7U�w�4(8F8�L�l�/φ!���X��u�S�9|3"�"�ᒷ3~�=��\<y��o�˴+���;\U�$@OgF��v��I�gG�����~s��ːV��<֥h��c4��kC X���[����m=���Yر>�j���b�ȊrhEɚj�d������,3p�O=�4������5;TVr|���Z(=՘T�/%z��N��JBR( z�]yʁ����Z������ə|�q�;/�dF�������z��mO{/��R:є��O�|��k�S�
��s�<�;L�6QѪ�j���<jl4���e��j�H�yf���'�4�g�Ƶ�7����1�Az�!y�՞�h樘u�`WF�'XR�b��n����{Qo�zٛ"��C���48)=E��Y�Π.w�X�&g���&�U]+h��h�U����ˎ�
��%g^4u�=���U|�Z�`B�"Y�<�B,dn��j���:&�8��u�\�����V�c^F`7�@ ,df�_��[��n�R�ʄ\k��9C	�As��b�Є�j���=ea�]/j��B���<<��J>�{件e��k�W�����]���8.�9b��t1�+Nʝ���Z'�ǋ��e��Gz5[=�*�!�E{���iҋ�Z�ny���u�k���k���jub�k��q&�鲅�U�/�3�j�j�(PbƇ~����b��z�]�mk[[�Z��G��R�4�ӱ�X�(�=[\G{U��pIS�T%��B���M�=A�� ���{]y-q����h�b���˸�\��N./Ȼ�l�9�I*E��q�f-&�6��[עJ���	�em�=+�T��]���J����s�͹�k��Z�f\	)�݊��G�R�4*�Q���t:E�)A�t��7��gy���vww�����b��5=�i�lX^�p�s�v�z�D�p-� v�WϲZ�#}�)��b�~��M�\�?jy��]���)�s�-'�֋u��fV�Qg�pᓡ1�9�Lj�W���የ#
���j�z�����*5[���<�S4�_H���V����c��!k0tWկ�B�.��cM䃪�qX`�Ἠ�1�Gu����R�%82�Brf6-T�]��i��oq��a��P�R��1�o���t��Ɗ�<�~�ʬ+��F媱�)VC��IQ�{�_s��˼�K��:��-Q���:c��!�2�NC,F��aTn�1%����������p�^�2��Xu9pO.'�(��F)V^�.�޸W��Gmi5�^9�{���3_.K�b�R
�Q�(
�cnX�A�l�b*1Oa�R��*+��NI�n��S��~����2e�u���[B��V@a;�ރ��|7��@}y��:JŜ���������b��54&�L0g�h��M�"�`�T6��8���^�E���f�p�+Pp;ԩ��3	����mՉ��t��C����&�ċ�h>����׃/�|��E��8ì�n2^�̧Q��D�b+НU��4�i��,�L�)E�}.tz�Ю|���@`W��
��0��8Zh�E�ٸg������S3A���$��z��KmT��3�5�3#�����e!P(1H�A����á�����h�D]@o�[j�z�	�'��mz�m3�<��oU��Z*W��X0+�KK�"\���c?X�85LB
���ڧT�a��u�nIQ����ŤBmlq%(U��������ݶ:�^�ݶ�{u�f��'�v{��T�:u�b�11�H�s4X�}�~����҇�SA���5�F�B���èe�A�Z')qݜۜ�8�|ҵ9���*b�+�<�r���Ds�SM�ն�Z�o^���yڴ[&n�7�@[%�(p�M�]�j�0���9
Y8���>�1l��"���Ӂ��������O$o9]͔�2!���/ | �]Fԣ[����Jcn���]�l9��1��z�'��}F鷥�;Th�f��ݐ����b�p�C�z�^Pm�`�ve��ե0��Ql��^��X�Θ��]{g ����Fk�5�Ρ�b��r�*���>�����u��c�}��F�'�0�aU��w8Xy[wn`r�i��y��-^e-2�i"�8�(WEA�D5u����k8	�:�Cza���u�vώRIl��f�mM�]�i*��~2R�w8�r�4�`�9Vn�PP�]�|č��lc�^UǢ�ܗ��{V4��:�L��դ񵓨SH[��wh���xb����� �)�!��*�yg,�wx�t|0���ѮJv񨴗���9�r d�N3F�MsaM��TѲ"�%�yN�Z���Y�A�2XE��N1;���	�U!_Os�A���|q��EzP�Εv�U��dR5�� �;M�+��e#��ћ��Ԙ�6��/�V^-F��J񕹶z"\�׽�z��Eޕ�Y�Y��^V��iPқ(�VH�u|��Nж]�ԅ��f����K����4�*ܺ�/[�(��+jP���t���U��)ep{vQc���vmd����Z���j1���o�޼X����`'�^l��iH�Ŕ���抍�F�i�4�R�ȳt�٨�m�+��7�h�8E�C�+��K�<sr�x�5X���*D�
�;z���G��-F)!gwB����D�''�Jl�ow�^ʫ��3��bw4�����Oo�ʑ-؎�Kz�l�l�$��?S�T��D�F��xKy�.�0]�)�Ƭrn�(��1:��EL�n�,�꺥�"�XBnڦ+����6�mV�i�&e&�6����mk���|��0?j�!�ɫk+;m4�v>��Č�|�����Y�t���I��P��c:eU���6wv�,Qx�¶�o-U.�s�&q�+(��~��ӕ6K��z��/j���5��H<���/�Hvzf��rU�e�X�ӹOo�P7��TLt^IM��J�61F�´[)^5*,�]3R]K��Q�C��a�\i�Vh�c�̴�ZZ��Ĩ��X��� إA�(-�Ѳڈ�൵1�Q��F֋Z�ҹ�ahe��X��er�d-iD�Z��UX�5�jű��̷̢Ŗ	D�m��XU,m��&7)UhT�e2���j�ŭ�Q
�iq�131µ�\j�Q�flZ1Z�"�V��p��[E�QVڅ[VW��J�0�2����4c�k)VVV��m�#F��2��PP���ؖ�4
(70���-��A(�J�V��Q���Kr�Y\nR�D)jZX�QZ�m���DL�m�\q�)�KkEdch�V"��Ub*ȕ
"��b-+-�Q�E+m���X�J�������m�j�ňV�Vµ#acT�Z���?������wE�`�,*��>�Aw��/&�1�n�I|A�<��@�rv��$�ǵ<��Xq��M�����f`���?�w��`U��^3��dxz���������,��dL�o�46��u�Ê�w(`���0�|@����
�X=��^+�~u������5��HB��sz���]J����\��AʷB����+�ň%g���U�gi��2.�~�܋�^���qza���9QlƵU�}�sM��\&ృ�X�9�
�ͨ�y�sFsqm��qT��pl�{����a��q�[7��ݩȣ5:j9���x��i�^��N�zf�&N���nXW[L2o�PU�:ue��d�u�j�o[���k�U�o#�Ʃݩ�A:ظ:��x!(�ʝK������X�
�5]dc{RL�޻����-V�\�P�:�Q�1G�F@�A>�fcON��L�܏\7X�(�Wj���v�<r�y����/8����@�uR _�B�U��7q�U�g5Fw.��*��3�;nn5��9���uMy�Ve`tĊ|"Xz	�:����8���n��4���<k����$$�U;4����v�Y]#MVK�$�L���Y���^��M�+jǃ���4ܢ���m�����)�'Z�n��N�G���,�ݴ�ߧ-��R�(U���N�z��KN�XHЕl�]CJ��z�ʾ���[�rI�q��"{�����o,^�]�C��G܃&S�"jCB���0�'�X��Cq-�+���*�{�������u��|M7r;��O�x�1ꮣ�����B�s��t5�9g�O;b�b��UTnZ׮9�)]"
�W�q,_�N�f��\j����c���6��%]�
~Ļ�J��
��ox:�� gnxf�N����^�K�&����<)�W���t0�2�_\���b�(��G����`���MKD�NT�/�"�E�����N4Or�1��ڽ|��giņ�T1q�4�r58�8My�kE_�p0�c��НLK)𑊵�3��n��R���K���{��nM87�8�t�v9���$���7�$�N7�q��[���nsc�Er�~� Z�`��*#6Xq~����������y�6��/)�8@�$���K��]zln��9�69"*M@��5-ތ���zXca��X!��.���p�[��G���.�_�追�1)�,'�`K4ꗶJB"��(��@ѱ�,��;�����ݍ�J���(>3g&QV�YT�W�+��1ܜ�����ҽ�
�!��֮�s�����}K�y��ə�n@d�`�kvޖ-󒜡�Vu��&��Z��f0�w<�
w����"��Hv�{(*N�Dh�Cj�[�]Ʋ-
���tC/�=5�H��|�{�x<�%���}�5�Z��S��M�ŽT��S�cp�4�	�tY�r��Q�!�;c~Wm�����s;y�K��BEX�N�=9xu��j���"�C��VD	�&y�\4�2�Nc��,iZ��Ъ���z0�d��DX��ֳ�Z��@;�w�\3�1:߄��y�(Y����D¨��(�Hi9�
�R��fz΋�/d����$��-�O�o/j�M;�+�߂��S��8TK]zI*lV�bb�t1�+H��Nᗽ.��Pj���y�gOmHדh�L��)�	�v�'G�
��j,V�:.A�����R��јNd�7��t��0h�z�4�����8&��^N�l�����#��?;�����(��Jy�z��!U�T���T�;��:�R��B�`� �xrR�.���ͮ]�ˁB9���;q�2M��f\�^GH�^�	9�u�8d�Ö�@s�ӛ��#E�wev#��:x}����_�j+��DB��]������̇�a��ڸ׊�Q�~n�L:�hj�u]�|z�e7�Eפ����;�n)ԥt&����q��1.��͹^���<Z��R0 +�Id��ŗ_v򁼭�i!���"?S<N�a�s�p������������q�Ht���^ �c��]�W4��dmH�X��n�j�J�Yh:�x�!J�ʜ���W���i����.U�Q�t������z~�i{��z��ڵ��lXʮ�p�j(�D��F��KN���'���A�����M�1�C�X!k��7�x׶n��y^�����h��X��-�vvg]TtXvrX��=����u�}���\�+���5d��iO�����[�F���8C�ِ!�rV��
��wQ������h_K��e��hh:� ̼�3q\�oY��bwI�4o�P�l�����1a
�b�e�F�)+OV_P4���w�[�W��Maq2ɠ�;�v{N����Qn���H<<4VQ��o� ���_��*>��]�o�(o����	�.P�3*
{eZ]^�q��|�q���֫�k����&���/z}�]��J��9�X��
�
��3C�����=�'��lE��ZTB��
SdLtn�ʾv9�u�o\X:�jC^v����.���F̫�2�U$�Q#q�6cv�.y}nX❮�]�gN0&s�	�d��tnh]�/gR�40�^�.[Q�h_|�['UiNoV>A�.�2й]ӏ��m}Y���`5r�_\�3�����+��h�h���b���+h�����ًj�(�Q4&@�`�":r�hc��%�ޞY�õ��������l����:�&�K^M���R��\+�$0Pm���������*8�0�n=S�\�,XЧ�8:�f��H)���1p#E+xӄ��j�s��3̫�e�poƾ�]��L�QPT�ƲP���F��I�v��w��{w��k2u]��)��(�u�^	��+ӊ/W�'e���X�����}�{���R�����}�:��&OC�,��hLX�r���	
6x8%^��:�gu5�5���R;t�������GeE�~���gqpb�f��-�jW��8lO2U�Ţ����^L����;��<v��l�A-���T�WPߕ��m/^�ۈ}<g[��<8{!�x0E�47v��ݫ!��hʙ�#o�!q�.Nm0hHEQϞGd�Q��z���k����M��M]�W�O�����:��S��:}��N�	z٪���`�"Nڨ��G��#��[��y[�X�x���px����6���Nz����T~�t=�6�֑�觠���ɱ�&ͧ�.��3�'�c:qλ�lF	�prT�.�8���H�����S����(��z��.p\�z�v��%��*Ň��}7z����9�>��:;e�0��ͷ�;
<@9�VQBU�n�5'u���k�oz� ��!�F�*np���R�Q�Y|��~K���UE�v���+s>����.8T������6׹�bd��lJ�"���8]31��2��Ub��Ԛ��e�}�m.KO�g8�,R�@{�� ��։q��yO���7��+�"�aȃ[�-�4?+�qS��Y��G:�#m�Eɨn]�y:��P�D��vԇ��ps7x�)F�t�X�@qC m��9>K��W	�[W�IHJ~]
��Ǌ�MݯK}�j�pQ���}T�h�o���H���훊S��Tô'��-�mM����������R�(��#;�n�W�='�U;��~V$�AB�����LJ�w��;K���@�X�B�biP��q�Vq�uK-Q�U�2xV��K��ּ2�r	�N�
/Mau�N'���AN��6+E�b)����dUpNea��B��n%w�i�s��Gf�*]kv��iTq��{S��A3��BpI�v
��ׅ�\�u�^�m���t�V`�,��3�G��r������Gs�$<�Dv�𚹃(_PO+ml�i���,�b�2�pOrcv6��麚��0�q�R�x�k��z�fm��*��)NR�i	��&w��4d*�+6i��b_L ����U�����03�+y�En��Z���Q�N
��Iߍ�?5���n{�\��� 6<�s�����%]�G/{{����~�u�ܧ��(��h�%�U(F4�ޭ7�˥�KFl��tbǚߪ�<����ǧz�L��6ǟcw����������>F�c�V*~}CFmp�4�^.�}je:g9#���,3q
�u�U�0\6���λ�S���gEĞ�b:>Ӄ�j�*�Q�e\n�!�`¬��M�,[�t�
qS	�B�ܡ5�tY�x�����\�O9�{�����[�$+���C���9X�����)�������5Pԝ�Uo��u��Z�y�Ԓ�+��r<����0T��JE�>ka����Yۮ@yT�m�"n�doj(-� �u��jJT꼊��Tn;��)@���Li$����X������bz^� =��t�6��7	�)a��������&B�:TKj�����,m�ޖ2�3,OS�&6�U�ʻ ����V�1d�����ҧo`���Iv��uA�w�'hI_����z�T�G>�&[5NU��'�&�IT%vFN�������������/�b���=��e�e2�Ƃ�s�YJJ�`��sy�-ݚ��U�Ȑ�YxBz�18��i�f��6k�IxN3�1lʩ�p*���N��b�>�0/�=YL��W���9���+��jAe������t��J��G���s7Bg©brQ���,hw{8ԁY��oV���gL�Rm�J&��X��:���"LN��&��T+��`c�aμ����-�����o���dc���+�U�6�s�e�Qkx�W�tpK�^D��a`R����Fp�&�������M/f��/�]E�����`�sh���uh��Ԁ�ʞ�N9ҿ;\֭:��Ŝ"^e--&kr+〪�Y�>4/���٩�)ά�[�<��8yv�n^Z��'���<!W�pt�ҳOf,`���ds�kbcz��E�a����#O�
�;!���j���*8��Vl��¬�ã�޺��kt�&�
�T,�j�	�]4�ˠ:�nd��d��b�@���7��5喃:�CV����qJ�h̗$Tj��}{�^���jˉΫY�(U�����T��a��O�.�x�����9Y;�p&��=����������83�5�O;êm��ي��[D�~/��7X���c�s�Q�1����;
��^{ާL�)���7�ff�#��I����/
e�˕�A=ں�ء��=v�d�t���H���-��͝]���˔75��uqI��&�Ls�l��.hd����(�"B
-J��6X[�LSږ�������pM�L���/�L�w^g
���6"T�2�ĹD��l��+�>�۰.�%�U;�{k�ێT}*� �Q���B�r�aoV�X�U�Cv2P5�x�7�9l�����c9���X�X�;Z6%g��f!�R� D��`.�j��/`��9��v�U�a�1W�팢����n�8�_����M�	�Rķ0 19���vû�Ƈ����t#�!%�%
���|�:����wMB,D�n� g�K�0��֥�v�=��=�@�*Vg w}�8�!MyDjƋ������-�����P����i[i���썀�'E�el^E�0߄���(h8W�����Qb��d}����x�sq�l�$�����U�E ]g.	���]+�Q5� �ɔ`�T�q�KD��T�'��y�U�x�{w��8���B�@y��H��,a5	�Z�1�.C�mp����{�?.�{�Փ%vJ��b�4&/�)�D��dnsZ��C��s������ۂ'�]ŗ��p���0[���?H�K��MZ��l��wɊ����m>\�xvv��tE���N�Ѓ`��V[�\u�*�C��v
�\92�Hm��=�j(�tio.����O�U"�2�������1�v/2��o�t ��@]_E?`ifYb�}'u���Z�}��6���8��f�((&7�1��p-s�ywWo�J+�����	���X���1��/Up��Uh�m�%�Y���:�~5��lN1/��9��ܷ(k�ٛһ�ʘ��G¦��/-�ٷ���xS.aa�zb�R0԰��d��%�kb��1�2��܈�M�2��Sql*�(LX�u�GYȋQ<*ԲPLu����8�C�#�l&����K̔0_l�Gg����㛦&�x����17;jP?
���	T���������,65��xV��o\�k#��O��ld9���t5�O��>�>�*vkY��S��خ�	BƓdJ��Rz��k�z��KZ��9�2�e��f�H�+hxe�8�3�m,n���B+CÄ� �9X�zP#Ia����%��b���zc�t-��̾p�r���a��"�E/�It���&��X���c�zbc,��E\M7����*��<�aY{�b�ԯB˭�D�N�����@c��U�WLQ@ ^F�U�ѪE�F��rk1�C`m隆���R�c��6;�CB�n�M�b�N�%8[l�\YA��
wh����u���m	F��lѤ5�d�5|�k�4QQW9���\F�,���mҶ�n���c"�Jܭ?�43+@w��ĝDQ�*��!F⮉�A���T�+7Y�x��@�oPan�K�xR�ij���x)��4 ���V�F!Q-���y9W�wy���(�٬5]���uhZv��D�u�� [HժD��DM�b��եaP:S�t^�z ��9�}w�o�0�4��b��:$jX�F��e�ڷ�3�����e���8�tH�ܗo˾�c�̫�ܹ�!yܝ/�Y�R�v1�	�.b2K�;_m�i���viѸj��|̗�CB��VS.]kb�
�=�T����C��fަw
��:��bT�r�=�HRx8݌��\A��P������c���.�+�&��&3�X3%$�8T�k�ۼ�W�tJNЮ�A�����[�`͇ �}qnntw�-�Ӿ�`�k\fιܧq�K[=�ه7�2�E�I+!�,KS�����Ǉ�:�B6���]at�muZ+5j���0����}ž&rq2�v,�&d�����)�@���mciu5���T�Z�U�����XfS��ێå�q+�M=�������Ėe���r��
Q>ξ���q'�����r���3�O�65��4��I�lu�Pr�1�Un�Uz�h�p��yv-LV��S#r���9oe�;Q����v�q�h�Pו���,���9u�V�t�� 9Seg]��/��d�O,�}f�j�+66��
���]��L���g��=��׫�\��i�a��x��U�͗[n��=K�"kx��piedQ�\�;w2Շ��y>��z2���9��k�w�K�v��">l����*ȏtpӆ�����8���F����g=[��Ȁk[B�1��9ěj�)N�շ�vn}u�)�O ��:�Cŭ����À^�&P�(Ѳ91z$�w���ʒْb=�kX���j���K��]���-�>w�Z��V(�4VJl�;�C��#���cf��3��j��PM���6�b�A��7:�7y�
)�h�ūRZ�1T���D�,�ï��9�\�����}�&:�����Kb��u;�/)��д�*�<�3�5�$���)i-���ʲ���H�QKsSImhS�-vP���bևu��+��R���M��u7���Τ�A�
[ָ��o>Һ�5'z���p����ާ\�]���/���5��ݡ�}�W�}/�M5��Fj�Dt+=�*��7=�)�=ݳ%m����G4��1���k0��z�,�إ��e,dp�$s����h��z�����߻ޏB�

VŊ������b��U��imiEf��ֶ��4��KF�E���Zڅ���
Ҋ[*�(�̙��E���m-��6���nPiUm�#j�AE�m
�(VҋiT�e��am����aT�
b�-�(�X�[B�J�-��
5��b��V-�eTF�f*)�[V"��Q��\�c1�2�J�����h(�\��´G32ʨ�l���QQUG3!\-���Qb�V9h��im�d̵mmF���Q�pL�Z�k����[m�[X�������Z(�TJ�DKJ12�Ƣ�,��m������neq��\J�**	��)��j����b�e����ڕF(�ڵF(�Q��Ekr�VQ�e�*,��#b��ZT��-��R�Z�%ʷ)rµ�DWmR���֔�V5��-�airю5���Q3.bWĴ��"C.Zb���*�Z�.4LJ��[Ibj�ڪ%���e`ȩ�b�0}N�g5Bӳ�v
�[����6+�cGx�c��d�ȅ�VT��mm�څ���y�'Hު�x_5x��5��s9tS��[�Vƪ3�@�|�SP��D�u��MӜqe
��P'uc}�V͸��y/V�:�@���A*R/`9��.c �Mx'�0�t��7��uK-R��Zy�|U�|<�L�;=3���(�pT�iq��%֪ ��dplI�KdXH��s��V��o��{&��Z���3�ڨc@%F��@e860&p�hNs��5�;��`�f^��Hz��j����|4�w��[����s(Ɏ�)'ZLu�Ft�u��noUnG��e����à��;��� 4�k���֔=N֏ i��˄LM�o}oyc��|W]��yR觲�e2��Oyr�X�'ؤ鋣p#$�s���,8���\�-��^$��Y^U�7�P�}O��n����zM`K4}��H�.�P�s!�q�y<�m7��b�ށA��i~��4냯uV��p���o9�5~���f�#���ۇ+�OĨ��OOo>n�.pC�T@�TF:D�)cD:A�u���3��t�ߩ�g�P���nR�o����;��\���W�..�T�u+\��"�3�t�-��v�	��� a��K 8�BIVk���k��Jk}�)���� ]
m�)�RV)�_�yZJv��G�[�[��Q�W�*���i'��=�3oK6���kH�Enq�7���Ð"��X�Ht��d��_	��,_��Ac�9�����.�ވ�}��&e��5�̡t��V�2�Ip�e�P0�62e�j������pa��U ���}o�t)�v&���n��k����p72e�s0�1J�'�r�1-���8
UBs�֫�c-���ھݚ��6k
��й<�EF�8VUya�]+�a4�M��r�aK	�OȵQ��qBy�=�T�"�:p'�ٰ���o֝X��+�$0D<�,����=Y.̿m�DX�k\�����6"�7�m��b�]F��C�S�.����2d��}#uJ�՜�^S�����v�qֲ��@g���g��y���:� 'Ě7�s�y�����Kn$�L7bZ

�G�l䦸Z.e�-z^�NP�����u�By�Jz�ntҽ&ӊ����rļkYu"��A�sh�vM�E�Sg��.���Nk ~�gtVmS{�]�Kp� 
�Y�:���R�5�V���ה�yH���)�5�q�T�k�ݧ�5�"YZ��f|��IpR�u���n�˫�� ^���o�"��W7+b�k-q��V.�+r;�Ѿ��[��u�%��!F&���dm0gW�'��y�ھ��:�P�9�w]uh�&��&'�������8*�����;�tu�Ōmn�rv���1�Wgb����h���ڵ�]QU�9���|\
�t�ʛTã���ֈ�+���1�m���[�e|��p���w3y{�,�5����C��)K]�`�E��r�y�C��*����]Y���=�Z�t�|�i���/4��~�43.��é�Z�`Vʣ�=9}õo�9�ֳ�&>���B�{���Sf�>�b����82��T�.yq*���UfӶ�)R�e[|�ݬɓEr�%'�:���$���i~�հ2%N
�uH_��%���ptwMf�=�\7�v�B�<=e�Dc��yF�`��봊Ax�5�[�֓Y[W5�p�ˎmV�Eb�ȫQ�ty.o��7�Y��F�bҦ2�D[UbTN�XO�q s�:�{��N�I8#��ЦΞ�^�^U�w��Sޓ���S��#�6I�Ly�c���|�w�
z@����!p֋e�\_�W/zs"�G^�,EBn� R����<@j,��cǨ���B��Mb����d��+v+�Js�]ÇH�S�i��9Kjk��i��pk����Σl���w����h���'d�ZN��S��q����!Q��gv��3���
=7� �1��h��ԣ��
G��}�g�Or��q�A�e�	\K�ޖF|;j�Xt���守�3�灨W���ObZ�k�*�K�R�Zva�b�M|q�Լ�2ߏe�^(�Xwԧ�b���
R;�;����Z)ƺ �l�@t�s�R2ĨU��ߛ�6��D�͛�1�1*���D)���b�ZaYc��r#����puܼ0��T	�y�V��F-�)�WU1�k���v54U<��7������]S�q�qpb��F�-u��8@��fߩ)g�_�a��BW�cr�&6ǉ�\u��R�������U~*��Z'g�i����Ƒ��k�g��c�J��|���[�h��!q�.{6X����p:�czH���aVs�����mƳ�^���Q�SJ�+�^,���6�0��:�����s�a���֛�ۤ�v.�Hd!�ٴ���c/�4P���M���p�bb��c����u-��Q.���g�99ڧA��'b��	N�9KW�#��&Hu�C<�PK}���/�9[�(R���V��yм�q4� ��Fio��0�J�K`��X!��w���vxZՌ�/������{(X>�N�E�#��G�$�1�9(3��}7����� 9^��bg Ry�{��;:��c#o�
*�p񯦑/��F���%��r��Mn�7�I�����m�t�V�,cK��։�
6�����i\���|�$�>�k���(e�4"]����o\��������&�ve�G<ە}+���oB̤�`��K�^�A.:q_��h-|k�)x�H�yL�}u+Nٿ�NOI�bFju�γ0��&^��)�Mz&�p�C6+A�3X�8�y[�JK˹'���N�I�]�|X��qJX�IBsɉ�w�Z+������(b�C�?�7��7*nΠ��0�� �6�cg�vb�O ??0�*�|��^6�b�Ի=6��U��z��������+
��aUk���P	���q8$԰�J��%9��\�FxN���ͮ\�����5���~52ۯ	�#զ�����E�VK�a��@h9��n�k������G��T��*�J	m�G�n�f\�:!�{� S��WI>�D��������֪���%㘰�-А�xjD1���Ό��E�*[7�Aò< ��[C`� �	�R����형��L�s3HoeIЊ��9w:����{Fu�_`04љ�N� ���Y޼ܞ�SQ~��ϼ)c-q��L�,;�͛R��1���:���l�Z}����}���[YIe��~s^.��1��6�W+����,�M��g��x��Ԯ<(�x2.�,�*�T��[]A��Ǔ��ޥ��7�C 8E�i�1�i��}O}��k�X����h�[�.��m^�U����fE��+�p��
^��t8L��]f�N�u
�D`�ھ���w�tu7F���y�[o��z�eA^��&�&4P�ub�Mn�cYA����L�i��!2_��|�������;��{|=X�7r��*��n�B�5�l�^��p�屮&9�X5ǜ�5�aen�f���^v#oMC&��팉��IN�(ɖ0Y�e4r:Ϯ�p�;Y.�e?�]T�6hc��N�G��'%`���p�:0����5�&&)@��!��s��s~j��1�J�]�GV���<[����^ ��X�s¦ �,c�'�<\KU��s���f�b��i�$��ۛA�*�(z��K��U�~�ɡ�S2&6�Q��I�`�Ykn���T�a����~�xK�ά�m�����6��;�,��#�������a3�S���Z-��,�+�^��4��^b��w@mvռ�Ev$��57�S`K=]][������þ7�է4,��ZN�'yh��l��G�ηX���}�T�n�$�Kg������ݝ������@�N����[\��[�Rh����-�pU�萈*vP����p��8=T,A�����k���.�M3ٲ(�3I�:��&5�n������m�`����Xo�H,Wa��9�h���:����}A��Y �.�P��j�y�cR�widt[���U��4��,rļhk.��W�k(`bQ�2�5)9�[��ozuv�Ǔ�	^�s@�y��׻����Kp�;����ƅ���5t�:����vvݣ;�sY�\.�դ+.3f���Xq�p:����ً7����r��d=��F��^�5t���,�t^��l�n0����1�c6Pf�`uʡ�ў�8"�*�4��pq�C}A��KS[�.W0`�x͵[�nѕ�B��v���j(Ҥ��w��+�s2�q3��z0�X�B̾�;�YxH������ER*-��@�،�H���6#��s�1��Ր����9Y[��l>���vc��Us���V62=2�
���*ܢU�f,!�a�s�/u�X�s��Q�҃�3��@�٤�B�}�(tH��P�~;^U���YmNw���*w�*��5gv���|ŧ�/k; �������6� ~����4X�m�Iv۫G���F��|;7뛕��\w�.�r���L�uuT~�9Gz��8���&��(�S���j��갻�|���i�_H9�}3��6{j�{9C�y�X]��ٯw���D�KE:�D8�h��w��n���~EO��ggv3�u�I;��}G�&f�Y�jDԺ;���w��<_e�267���O�l�+-�J�m��Stcq��S��FT��v�L}�U5y�VEm������;m��Ľy�UfD�V��r�-sy��i�W�W�iֿU�.{��i�K�N�F5Td9���$d��o^�afofs�XN�a;"|����7����|��l���*�؞�������T�W�ő<ٟ)���D�o/0ؤ�Cns�� t�r���;�)ݸ��5��Es��Q]�����
�L��Q��~����}�$������Q�-i��s�R^��Q{syy��$�����I��O/L駙��Z@�L'ƭ�v��TLz�e�+�n}ګ���MZ_Q�$����W�N�g],w/lRZ2i�n���@� ���x����S�@U_N��|�tt�	D�x�1Q����������2$@f� ����U��������m��y��?Q�_?t�U|�R�#���]*��)�}q�����,[��9ӎY�oOSm�=�Lr��{��f|7ކ��Ox%;���d��Ru6�3���w<\q�S�?7��Y��r�>�jRԟV?z�e������5y��w[�䍻�F��޽ٿE0��e힜�=��§�&V�r�.�w.�1�Ɩ�i����N���X��K{pJ�+��Y���inz����Ci�l���*�j���b��'̼.�7O�Gm(����yoq���lc�Y�I��[2d�Y��ݲ|���㕺�p���hk���w�W�"����
�r�V�W�����w���;��{��]�ݛ��6�n+��M�z!�,$������h�ɡ�cg�������[�o'��t�)��Jxb��sPๅa�ma����n�(�rOzw�9�/z��^�s8�I����������"W1��_v�h�ݵ��P6�ϯ�At�����WR��E%�b^���9�.���etD���;/��vv}EI��f��Wi�o��xW���r�3��V�ޕ
��C�t�)���m�:!���VHՆ�>�Զ��,���pU�=v��Ҿ�%kwA������-R���5�cw���'�Y�JT�� F�=�]$���m��Q�SjdN�ᘊ�U�-�l��86��c���ٹ;d������c�Ѝ_����M+:'��Z��ޥ�Ж�L��On�5��y���'7��K��};��5mc<��{ڞu+�<��XQ
E>�|a��fd}��⻒��y���,�L�ɚo��D�jk�2��}�5�r��﷫i'�}���Ś�$���0r�����]��Wg���^��s�퍩��2�SΎ����*.8�!�������<��xZ�	g�3��ro!���Q�9��}[�����><�m��/ͼ��i�lQ��I쾿Vn
�}s�Q�r��&��n.��ǨĸS9njy�[{9K�yl��<$���Fvt)�؞��z=�G�I�d$�	'��B���IJBH@��	!I�HIO�!$ I?�	!I��$�	'��$��BH@�RB��$�	%!$ I=�$�	'�!$ I?�	!I�IO�BH@�bB���$ I>!$ I?��d�Md���n-~�Ad����v@�����;��
 )E
$��� ��* *�J��\�qH�TT�D�J�J�+�B��u�Ƌ,*�(��U�Rk*;��2�L�U��a��֨�.��7l�m1�c+M6�ສ�a�
 ݆u�,��[(,-�͌��E����X��bխXɲfPWtWj�%m�X��6�)(h�m5��e��4��V�Ԣ��M�Ų�f��i�!�b��itڳT�%�ِ�6iD����r-�i��c3��(2��TE�g6B�d-���j��f
��     �ʒI@�4 12� )�L)JJ�CC�� �FhsLL�4a0LM0	�C`F)� ���       �12dф�14�&��HAI4	���<OD���CaO5'��e~�����kz�۳g��	7�a�CP��!�Y��� Ԅ ���		L�?��9,$h ��G��������蝇�3�@T�����P��T��	>APY&����� I�>��Ϯ�oq�?��_���:�}���  Il~�.[/�}e"Mɩ��&ߣ�w�)(hP?��t�9A�c���;�ǶsB�jQ|PZ�I`Tю#vm����w��ޢ��n�k�z�#B�7�o7S%<�y��yB�21A��y� 6��w��C#1�Mբ���W`�m�h��Ts(j@��� 
��=9SO*Z�N�Y�WYc~�W�[!�y"	��0Q渥[��+v�����#Z`Ӕ�e����aڳb��r�w,�F���p�7LY��Sb��2�K�p�˭�H-a�<�g 1�z͊v�0��X�@n�Y��3Ao�b�x�XۭQ`J㼗T�0n�%fd�1��l	ٗ]��T*GA�Y���P����)TVU!6���̇b;G[���%����d��k4�1�Pg����1ٛR�l�r�ۡf�WCa�G��'i�������lRכ�	�5�싈�ފ
�ڰqW�ֲ�O7���t�x~1͗��܋Z��!Kb�^�!h��q^�^ma�2=u���VN����Z�@Ն���,
�.�X(��m^*'7Dj�B������M1�k7,��(�oi]�����"��1�@ͷ{�$�V��K1Xoc9���:�!}�X
v�*����YVݦlrT�Y����//nb�2&��	�P�sMK`���B;ZL������AU���+
d6��Be�SҚ٘H�����S�B�[,^c"��es<��p��ѥ����VA�؁ͦ�Qݼl��C�6�ӹyO!��u�6���e��f�hrL��[��D�R��cå�0m���ڱ*7��̛��+�z�0�t�H��ԹQz�g1g������'���jJd!/wwn��Ȭ& o!�TJ�r,5�f�;���]% ���U;�3]j�1"}[D4�X��Y��ر�
�ƭC2��V�C)��p:5�%�I`��ug����jY+�c�VKD��l������b�gq>+�Ɋ���ڷ2���\I�PX���5n}���sv�VɎ[��=����: �ZMswy�M���/i�T�7��3wQ�#o@jۻ�6�їvj	7M���&z�WIw7}ZM_!p�|Z��*ۖRyt��]�ck@
f�*[�@#���j/�4�^���4�$�K��и�4o��*Q�l:�������5��
7���vM��(�4��37���^bw���) �B�ą��h���CmZF����t�:Kk:�B��YHe�.�\V���0��W[���������U�)�R�n��t�.�A;vqf<��څ��V����p!"�(����M���%��A�Pъ3�M�k*�J͎��#�̫a�5����z����5��L��*���m[#��
T��U�WHg�o($$3��$ڐ,�����VM��4�i�M���F�-\��%ڭ����wF�e	���E��ٳ@?�2q^LS]�$�a%��c�Ԫ+�&+2��H�	:NK�Y��V,�Zd�vvo�b"�+��0�կ^��j*�&�X��u�{�S���?�*��Wz	���Fv�:v2�8�i�t�ە��Y)K�;f�͵�7�iJ�9M�jX�J�4��A'��� 1c͡?�K���V�xm�޺���˷��g���ԝf��a���B:�����=��_h�����Eэ�P�أw7/W3�t쎺n��>�Gw�_8���i%wR��W0'n填)��Z���6����^����3�,����;{ub��bG�K[���X���dK-r�]�.�(�t�$�lj�\�Lc!%�V�Z�T�ˀ�[�ư��fp��!^�e��m��jt��@Ù��J�&!خR�iʉ:��m�j�������\٧)Y��w{�@e�p��Z92��m ��d��qV�+ms�ƺս �����h�C}fQI9H�u���d�u����[��W`�H׶V�q������괇�P�ʎ*�e�
ب;+���sf
�kUt�SP������=�I��w4K��ەe �`��ow��5�3.���̑j=a�B���iw��\����CI`�V�<㿒ƨ�m��(b�U���)T�ԯ�t��E]%m�fA\�K�ø�S��ю�Y�H����~�ꖌ��z���G�|+�ˎr��	�����������<y<�vƻ�坛-��l��Q��z��!��,��ȡ&���f
˲
=[#4�!G��XO_p""*H�����]�>�V�jd�936��,�y�����mD�$e�G�ߙVkD�+2�s��4�v�MQ�.ap�Η@	PLV)��EB�نW9ktt٪�f���wQ�@*�`lnV��$9i�{��r��l�_�᭞�����󥁭�.���X���r�VQ����A�r�ݱ!v�K����`F���x.���k�3vH�L:rke�ࡻ�y�욂m����';�� �]��%h8b�S�Zfm�2�V�ݍj;��6�E�=<�l�w!�qӜD�[bc���G�t��H$������L��W�OK삥X����9}��]�Ic0p`\;r�
vwG�2*&���<Xj��Ūc�mЉ����a��K�_*0nM��w�l����H7ɉ���;M���y���t�擴'
;m0�t�ڐ`�C����@7ٕ��>VJ���]��}�;b+�U��7�]�w'�A,��B�J]�Q˿��b�0^���QF��g;���v�z�c/t9��Ps�+R��ɝ*|+c����Z��]���^E��ҥy�l�́)�u���(E�� !�BH��t���\��5:Tqf�D�z^�k�0�-��M[}!u�K���:�c�8!�%�')��R9�W_VIG���}69w�:�Ύ:�,�NS���s�I$�I$�I$�I$���Ms�9	�ɾ����#r�16��S����|�4�*��Sו��%��5��T��N��r���&+6����ًmt/4��G�.P�[9���v�s��ma]w���w]FȢ���8UԬc�;}u��4���8�9�!v��Ѣ+P�ِ�{z�i�Y3�ʕ�Wd�ڛfM�
}mbԑu��b���g1\%�������a��gAff��jh�@G�ZA
Fͣ���9�uq����4 Z�G���u.��swD�#[������7��}˥=\�,gA��_d7�h�E[�ڣI}p�r�Q��������]y\Glꛍ�ս9ԛ���U��A`��L-�1�q^�R�˝+�J6g���Ϩ������G��5�p�k�֟���o��D�B|�I~<�@��D�@��?�O�����n�ސ>�ċ�J��6���pWy�}��^v�q�Hɨ��%�.o'Z!:�����ZN��, ծ��2�.9|3m�-J��fѠM��t˻�E1���9�2��C��K���lJ[��)��c���uʱ�<��+�``��f��;<h��E�.7Ce-�f��5}��۩����zMn�^�4���G����V��Vd毟2�p�nێf�.����P�O+�4�m���!��.	K$7���I�9� ��%p�or�I���
��l\��N8b��	�u���!���f��n��ߔ���o���v�ږR+2�tj�r�b��j�TJ�:}]M��/1Tz�`�Q�EI��AKWr�[�����wv�ECɗt�5�:х:�śt�s��a��
4��5���d��NU�6���hg�o��e܋�Z���c�[��	f�9��"�9�em�9�Jǒ��
�z�s�ϟR�
u&�n�m[-���F��;��@�C�Ί�oj�Ze#�v�
��Qç��Z�,�I4��V��Smty�������z�c5�5����a����}�_D��Eug��l�k-(Eg^�����aˠ4��̮��p�y��6�Z�~�2�r�@]�U�6}��-1��+w�������6�ش#�2�"Y9�	�0v��K��ݤ�-�V�z��ؠe]�z�޵M����bH ���[�hRx�G��h"q
�<��u�@�!�1�UPX[��g�p�g�N�Y�`�i8s�w�����'Rڼ�Ɯ��6F*�����X��!�Ȅ����#��٪U��eq���`���t&�u:2k١��C��i����F�i�EA�y5t�˻��	�Ũ����|1V+	
�n��b�b�F�v��[;�p��α3pe����M��ї�un-�-!]z�ݐt<�������A�S$ó�V>/�|�8�+pR������	2���%L8D���G$��zt�sɢ��:
(�vR��A���򄷷nP��W������CrVl^SuՄ`����=�;Pc�q�)>��#uްQٙʩ@9��9;̭�ycXdy�7H��Y"����x�[-#y���.\���ײ�WI�#g2LV��hc~�d�0��;)P���	�7�{Rݘ�*X������h�:�Xe��9+�:����V,T�*:�v�ʗm\F,p�q�%����ai��vf�����hv�C���Xfv_s�T��-l<�d�k�wv�>z���ѝ�r�R��0��i#�⑶�m��6��\E�{�ջ�ޫ;�(C��'AKޗ�gb9� ��X�(*���[�,�k�@��H���<��7r�=/ݡl�tO�&%�V�ε��i5pݺ��H�
�Vԍ��5��� �1tL����͋�n��Dg�4�;)��x��v˴e@Omɱ���x�uA�9�t*�%�|�n*LVꁎWmc�Zg�R)�b��|f@���t�vv#�vK�e��|,_W�ي�g$�C��/�]��&JOHW��if\H��t^e"��9�������w��L������dr^ڇM�����<󾳦��oY���ϑ>� @�b����b���.@�tD��~���;����}}��"��B1v]�S��TX�D.�J�s���b����m�[��p�u*���
^u��̤}������!T-�q�����{h��(V�om�גᴟYpٗi��K�����Ů�M�n�WL��/ȡ��wFK�sGζ�'qp� {:��N�jɱ�M@*�g��-NM���-b9Q�nj�n�m��.9tܮ+V��Tm��e��,�.e�#q�EUiq1�V(m
Ͷ7v8�
ZP3*�an`�1�"�ne�m1�-�i�nL)Q�V�23IF]H������=���:�5��.[}������H�2�J T4��|��z�S�w�_�L�LB�V��l����6r�����Nεߔ��x��������z:J�����:O�7{a�)��So��M�w�u/��9G3�M�7�3<����>8�{���s�fΐ���Т4p�>�V0C�Wj̮��a��X���x1�>�s�K�5@������f�W�������YY�t�!7�v@��R�I$q�܍be�r����c��ٴޚz����wsy��n�L���&�T�2�q��N!���1�{��7�r��N��TS��4"&q���;׺��HW�{�A�W�S�;�N3-&j�G]�����>��ݾ>'=�hqק=��=giY��0�y�ƻN�������:C�Ǧst�5cfmߦ}Z>���������cJ�d�i�G;V6�'�$N�Mk����6[*7��^�]qʮ���n��ūW~�w��Y�*��>�+��E�< Ƶ�4�wE5��4��z:�v�,��x�T�6��������g�XoW��y�6�ͥr����11�;���)�Q���N��|C�7�W]���^������1��5�@}�b�.��\����ӧ�o�i���Ys����;Y^(1�Ǆ>�U٩�<�[�]?"��UK�.�)�xf���3��(�gs��
��(!�!E����*Em��o�xW�8|�V�LAX;�;�oG
���ot��5�s�����ͦ��OO,�2j�r��4t��T�v��xt��E�I�C��
�?L14�g�[�:O�QgN�I�9���w��穦x��,�c7g��6�����E�Ω��(��C�K�=�Gt�;��J���NQ�&���Z�謊���:鑚�A)'��"�,GHO���ܳ���.���N���C�T_|���ޫ�PSL��Bb��U!���r��Wyz�:���^��Le��p�����+sh��c�+�{�/�N9��
���F2�:F:I��Y�|��t���v�M�����`�� �)�^�E���e�Sbq�t��N�N%M5ji�TF��\����^M�O�Y�~Luv��}p��t�J̎����q�GF��F�׮���묿��R�>]�V+EWC�
�3^�	B�vv���.`���C��!���/z_��b`���s�z�5���<��,���@1��
���_=�G؅h��|j�i��i�f�������n3}�Y��j�y���m�7�QM��W3|��
b	�Ҡ+F�L|�<���j��,W��X�*��S�2˺:[���n�k��x;��N�+��aQHc�����{�H|E�*,fQ��>޺�I�8�wv���t�u�5�C�q%xη�9iw��s���<I�{2�8��j��`�6>��yUX��,!�;����<�*m�v�;awKsμ�ӳ��ND�4|��Nr��/h]�"�{ƀ�,Z44� R�5b�������iC�f���?1��UJ=�}r���E�Ə�U�10ḡ�rj�x�u=������R��MZ>o�7�W$|An5&�����Ք�ev�i؆�u��5�'n�uM����}zG��Z��f����;f���c���������j�!�^�׳٣X���!��,5c�����U�������o�3�5�r�פ����J�jg]sF�{�I�W�R�R���!Co˻�y��X�<(�
��R�V���W��*�S��
�?Dh���M������w5-��H8�]�cu�#ׁ��v�#e��=��.vm������59꒠�>��xQ1Y�*ZzZ�]'"��y�4���u�5���xm��S��W���)����C��.�9K�.�wE�^��bz����ƀ5f�'�+�m����{M|��p��ީ�9�~���)_S��*e���꫻�{��K�T�!T-��vT��b�ڢ>"����[�v��RW��P���J�	�(�!��)Μ���MG�q�w�e������T���5K�����PR��\4o�tx|�m�=��S�t�gnا{�9N����z��+���L�tY�ݾ{�7�'mO�����x�gZ�I���{B�OQ	B6�0F`��V�}pB����x^�LC����ۓ�v�5��3�h�P�#�����B���t�_I��
�|���\��с�n��������[���?�]F�|)ܖ�̘x�Ok�J�ԃ{w;�[R�[Ft:O�/F�Mw������a�Ȇ��Ű�0���Pq�g�U�����g�ճ�f:P��ggi�pf��DC�թ3U�q+�D�W  �e^�5���-�m^'��u&p, 
�ks���)��O5�h�N��Ef�آ`G/~O�q���w�h��ڲ����tx���.@�
�:Cy�q��7-�6�K���m�,\�����wʟ=�u�/�9[*r�Z*��m�NN�v��k�!��N�c�@���V��R�Ĕ�*��.or�,��r�<21λu��˰�'���WD�[6�ʴ���/������~?�R�[�fZ[am��S1KsQ31�W�Q̸�-md�LR�YWIp�)na����k!��-nR�2fR�1+��l�i���I�.Z��1P���C�"ʖҥq�+mq��2�����RW���Mïg��˽"U�(c��|���DvRYv{�i�x�CO�o]����}1�4�7�EPW�T�h�֝`�(���g�����3N�ݾ���hs�c�t��6r�4j��}�����JX����j����[�vͳl16�{v�ո�h^��i3���{��|����v{EHcY�nu�!�}����s�m9lX�=��၈>�[f�� ��DA�J�y/�ɲKG���]�ݗ|Rݰso#����S�N)��I#�rtW_�r��v�3;�
o�P�^��׫߻�;{OG�;MyaN��N�Z�Y�n8�L���:�0�u͛�l��Wn�Y�st6�Y��u��8&j��~"
��\�Ҵh�)i��@檱d�`ư[�����ӧn��t�:���ַ��HT�8�{|{zy���t*T8�N0ľS=7��0ᣚ�SHW�~�֦��1�_�N�l����s�r�ogܫ�$�-�C��\Rw
�G�yj�vUu��j��U��>�E��{��V�,��S��P�Ep�,TGn*Xj�TG�����z��w��7�ɉ�oxuߛ�'�v��n��M���_u�N��l�N3��-��s�^����@|f��`���7�;w«jr�)���Z*���a��u��#|h��Z)���&>0����E6�3Ti.0L4k����S�Ǹ��N���t���gzjv�S�G�қ�F~�Pf*|�j/��yw-��g�$Ƚ�9BC��)}���ɶr�M�i�Wǒh���=	���yd�(o�=��8�+���hx��>ć�I#��F^	��%m]�m�Ҽ�c��7�uf�*�-GѬg%T�Z����%\N,K��1�~A���O�wb���ɺWS��x���\��֖묛#|[�G�nf����k�|яw��o�!���`�BK^n��w�/��F�3�w��|+�=4�c?�ױs�Ȫ��n�V�ί������������������;)���KFv1��<�,'$��[�b�4:�׭R��Z�M�7���#'*�5s	fT�sfik�2�q���齢�#9:�#��{y�����aW��uh���+⣴S���h��O�}U�{�\��m�9m������yo4���탦��X68�]��/a5|i$���l���cFȬ��v���t��\)���N���� ��r���wdް$����s!\ڪ��?*���^�ug�}�V��)��FMR�4DZ�3u�Q��y�Q*����?�,!�u]����ʎ��&���Jv���EL=
Vp��]tqʺ�q�1Νj ��������ҳ�ov�|����#J��L�Q�e�j�4Y����ٞJw�C�����d�x(�G"2Ri{�E����w�*�����]�MG��ߑ�y�	[��������L�/OvG�>�d�N��ç�e�t0��5E�m_�V�}���׾�S2����O}M���*�
���W��c�͹u:$�9#�əDnm�S��~[�T�X��E>��)�4�y��SǗwXΘ)|��#m#��w/�G��?�M{qK:C51t+}v�#�ێ���V���L|�zk���1���u�w�R&v$�B�*��soO��z�_�����	�'��� bC�N�!�@�d�d�@�)!�$7�^n��q��z�;I'� E m ��$�}e�W6�>$�2��a����Ą� _z���%�a?��z���3�З���
��z��c�{�����4��\l�xx\�;���+�	/�42�r�yX�`3aB�8���Xaۘ��em��.R=}��G�䮅	k������f���'�x�hн� ��ˌ���\�����nt�ti��_��?4��p(�!�O$�n���*���R*����{p���_9�j����U��3q�^��s�5�:U;��N����sZ�t�C��pB^�5>�7m�:'Z�r�Q�����R�l�f5C���l�W&�V�+��dZ!Ux��ל&��L���U&-ۼ�C�dc��	��Nʮ�j�����Y+���Lى�dew|�����ɘ�jʕ*K����r��l�s+�-��J��4Ҳ���J�E��X�q�T�KRܳ2�F8Zث*Ki[Ej�EU�W1��ffVҵ)D�jT�#Z9�eIYh��1r��jذ]\�E3%*T��F8յ�QQ>M.`�ߔ����קQK�;�W}����|I2C��Rm Rl
�O�$+�8��`�|����RC����XCj����'!����0'���5�Ԑ� �c$=d�$߶�q�=CI$�8�k��םBV� �&��k$�r���@�v���
�v^�Ԇ0��<@��@�!+$��_�$/ņ�`k��y֯���l���|3Ԅ�HB�!�%d����><�|vI�iR'�P�i=�!�bC�u�^��D� �� �$醐���� �&�i!a�=�� t��$:�&�v�k���q�<HC����]{ԇIt��$����O�ē�v��Hz����9������WK�@69�|\4�aWS�{f�*&^�Q8�#�O��}�W���}_+����PVO�$6�L&��B�q�k�gHC:���y��H�i8�$��@���6�l�{����D���;d��m!&�8�N�i�� �$�;��TV\��H���x}$m9&
~)ڟ�M�F�r�f��⭤+�$��;�f&a�����E,�R�Ds͞�d4ǭ�^+��/���vY�Eٹ����M���pavd�x��Ͼ��z�x=eau��
�U��V�I��q���r�ĵ��N��d��Ktq��q���n�q�~,�q�V�Ȫ]��ڌg�=���Ʈ%>��F*���Yӳ��2�]=��z�O�x��/�.��w�-Y��zxb�H���+���H�����Ν�݃����I�qԱ��-�$_	ո9m�l�M�.�zo_Z)�7��o/����;��so.���.ӯ���p7%��m ӻ`�.�~I�yn��ܵ��|I��`���|żDJ*F�P�$Y]������zҟ�Ge���57��~/�,=*(�����9躰�z��Fe\����|+#�n�a�����iq��p�`�T_I���M��'��Wme� {����_z�a�<�b�iZuk'�u��7(�_�~���PKNܻ؈�<m�W��F��K���#���Ǒ��7�䝽��;�J1���'� �0�w�4牻8����������c-{�+A<ޑ���6��X�@FO�ief.��E�vү4h�7�����Ǉ7\�+�H6np�݆�K�ws5{y���T�b��^ߴD��ȧ
=����5��E��/Z;�mJ�[�vS�����`�Ys �kD"�{���y��v25��x�)�E��fU�������&�	���C�2�=4"Y�fs�h���*�v�,V�F)�ꯪ�����D�I}��_us��w�"[��]�Lǒ��褺��耦��l�b��r�{��0/�"Ƿ3�+c,�G��Q6�K��߶��X��l��䒿vi�c��v���J��U11o�=��b�C�{����B��Ț�Q8��T�}�}��E~v3(f^~\^����w���lwo@Dp��m^żr�+7v_m��3���3��8G��E�Ro���K�8f���d�������g��,��oޚ=����r��.]����uD��5�W�����YAd[�U��n&��\��$������䧚٢=��=(Ҏ����t�׶Z�5!Z7�!���V��Lx����#��ူ]�eg-�{&��U=�=m?5ǴP�鞹�����1Rc%5s$�U�Y�OA~���o�.K��j��Z�Z��4�@!+V$����c��ѽc�m*B�2��#�Jx�9�셙-*n4&76��ډ���� ՝*��K�w� g_L���VTLp�����!wГ�'������9��m�X]u�m���U4��U���C�]�w��d�;`�)�����v���ki;����g#;=��蠒OpKU(�ڮP
f��Iֳ�����[ц5u�l��/��9Vp��kv��4�r:i2�4�D�1��P˾��	\5:��t��s���5����-����ͫ�Q�ݻ��qa�4_I��d�wsZx��S̸@��w�����s��.�vجJ�4A$��h�mD��9L�&m��ˈ�f4��hR�M5s+u�Y��-n��
Qkxkw�-��K��b9e˖���"Wnb*�TV��:�SM2��Z�Y�w���K֥kWYq��T
E	0��|A�����^���$C�m�꾪���7��V�[�? ����>۷�h��B5��A_�-�}~{��&�}c��[ub�ݶ����4�n�b[�,���\�s����גi�3������<�"A������^T@�e����悧�jv�S�Gzҋ����K�g뤻H����-f��{�"��vy�#;_vlm^�%�ҬV�.�����;�8�n�)�ƀ��6/q��� U��{f[��&�=�V�E<���{�U��1�������:n�c�+2jE�mrrc�J(?}��}T}���~Aܡ8hjl�lb�yz����y��:��7��ּ�����jM�'�$C���͝��{g{�mw�cѢT��\�y���v�z��p���]yW=O#�T/F?�p��+hȤP��2B�4���ꯪp=���0U���n���>�ty��UzO�
iŭ���U~f���g����RZ�V
�k"����[�q��"cf%��v�Fu�&�<�Խ9�\d��=��4J�V׮����b+ʡtVn�"����Ds�n�I����W�}_W������_�_<�����ȮyY����ڮ�����+.�����S��۸��,�tb�>��-1<�Ğ�a3]X�YV�Gŝ�¿��x�VጟBȨ��<|9s����ed�os*�[���m�r��W�)�����^�y�s{�~�׼,[ev`� ������� ���>5~���-o�������=ξPY�޻���Gzqe�ap��,����M�����Z�nUq}=,��w�m�a�z�:�.֐�q�zE���" 4��Z6�����p�(�tE��APӶ��Oqb�Z�v,�u˝&��\����U���s��`yb������<�W�~m�̞:B�I)�4����G�Lf��(�:H�7���4�yׯI��tʎHDE91�N~���<��ߢT�*s�Zif����s�W�,An���*�����'X�d��G7��Kl��m�Y�n����xA̮�3�t�|�W�b�h�{�K�D��W]}+x`��aǮ��Uن�)(�*����ʏ��}�����~��������v����9��Y�0�72�a���%c���*���w?L�.�P�J���k%UC���Ե&t�6'���n�X�Ǧ�J(.��*5w�=��^�Ɨm�q�rk�ޝ������6^������u|���lǮ���d27ص���rn�:Ƅ��[�;�GB5 �:Yڞ��kh�V���â����xk����"�I���i���U/;�+G���S!q��o��>��*^]��t��,�����э�L֗��+���Tё詓(R�j̖y�KF�kXt��:n�8Y�Ǣsw��t��;jg���;.��m�ݵZ�WG.��S5�(-ԅ���n��&�/m�it[�l���ȃR��ȁ��_��]X��=�9��X�c9
���a�y7�*�����;0���N⃷* ���9�-lc��7�[�����ce��>�}�d׶�N�S"��\j1�D�Լ�6��ms��"Ѕǉ=��6pF��!ow2�ӧ!r��c,�u�d����bs,[��KqYw)� +�;Tu��u�W�:�����q�:�r�:��P�w�Q��Dޙ�|�S�as�*[b�1�3�jc$����'�UEաmF)��*���2�Ԩ1XѪ�)��j5���m֛��X�̢�*��S7�-eTīVDF��Z��QA���#���w�������www^�	DK��^j��%��_}U����}����-���z�2/'+b��u�����a[�r��G�p	<،��KMK':�]xe�F?mg)c3֚̑�ݭ�7s�Y7��[��h������x��>+�۠��:*u�h]�s{eFk�W��\����8�����	�W�*@'��棖~
����v��"sY��Vwlt�-t:����gQ&�]�*$jǧ{%dYͿJ�Y��O�Vy7�s��c9�۽N�%i�3o ދ��6�Z��x���\�8�NF����U�g�k���}�m�����"CuڽF�B�O�}k_��W��j��'��wN�g}Tg3���j�p*>[���#u�֝���k;H��7#�ʋvM	��T�4��'z�R���X�Xw��q���sYJ	)�ꯪ-9���f}س��i6�?l\+���@P���7b�6sF�6�jfz�ߴ,��2AKb�ic������)t�B�
�%��ã���^�͊���6���g-�a��?*V;Z�d��t�n5�.��Ё�E<����#���\Lp�]���;G�"gȒ��9~�'��i��6nB���G䳯�������<K��K�'��e�M����A]�o{�����;@z,#z6d�S��5v�N����'*�Gch�z��ӻt-W{f���5a��RA�{��v�˾ym�Q^��h�p�����R��=��up��[+�uVr����|����k�}�-.�
$=�x�����RG��4��姒��S��ֶ,4~�<� v�R~g������guI�Fs�ȹޘ�NsdtϪ�+�to7�'�*��%���o&%X�ol�x�7[|����x��E�<����6�� �����C=vt�u��������m��d:#)X��_����������{Y���+��\`��=3���;!n(TR99?W�����]���_��} 
=�`3�_��P/�D��^�(C۵����5+����/ܖhȶ��i�Uji��2>v��̟D��0>|��,cR����@z���جi(��hԆwa��-��>����{�ھy�6_�>��� ����̘�����3�]g9#��mU�����mA��L��ߵQ�{�Zv�!�Ü+v%�n�_FVqmon⺞�<K%���7y0-r�k�I|��U���x��׌\�夰a��N��G�qH�JF~��~����:���9w��`]�T�L�nǢ�rE�P��]H���R0X>n�Bn��ݨ+���f�5w���5��7�}=f�}lQ��y<��U*�V�W����w%�s�b�¥qի�Y���$��*V납���zʙM�y����f5%
η\] ���BM����=��ol<��LSm�<��5�;���Kےʲ'm9�˧B`�շ�Ivd�T:��:�/�m��6b�:Gs�i��vңIHQc��s�����
Aʅ_2ĆI4_�ʏ�U�e俚�B��Y�X�Â:�v���Z�"��x~�f޹���8�m\�'�ǜ���X��[�
�C�[��q������8hV�a�|��Z/�P[3 ��hu���I�f�Ur�&p��rS�;9:;�#�M\'8ź�wR���Y�p����X��`R�w=[+�#;H:�a�Q���B�3t�F�2��[ڨ�jj���-�����\�ښ��X�"��SIB��Dt����uh*���SHV�J�YEY�Yq�X�"7t�;M�� �����λ��lf�Q�у��=�ھy����o�:*�˗�k�L�lO��Ew;�*͝�o�ڰ�\H�yTY�q�ΑQ���Lۛ�qXf�vB����x>�zH���5�l��R
�_�����C�����m={Z*`9��E�92z��9�w^���s����>
#��0r2g[�CK��p��^Z�5#l�}��
�*
���F�J��=-&@o��"��i)��p�x>@i?dզ�$~<X�eT�6���N67G&�(�-ЍFQ��n�RF�2��������ҳ`	�!X���9��o�%�Ǫ���0پ� ~�ƫ)R�/w�=�gҝ���rz��O�Qye��ykz|��o׎t=��
+�&saB���v:�Z���*���+�T2�S��
������9惼��猒�U���9W��xm�韚	D}�W�Z��K�2������F;�x��$�蝚8@ûa�!<�t�[j�5�^	����뢇��]�J�+��1���8�*�wY�J��-Ԇ˃d�]����3������S��cm�D^ll1<��6���әsfOBz©��]�bT� 地�� �F*���b�.�>�����n�k�?!�L��=;�|��A�Ҭ󵲱z�٢�\�pGA��
>wmܤU@i�n�q^1���9������=���g�^G^�j�K.����������zF�^f�(�<}^*��+ ^[�W�gWK��]e� S�-Q�7;56�Y��W�k{!B�9�e|:�x��n�_�����F��.���Fۉ�
�􏹲���}��� Ǉ��H�Օ����<�𮷞����\$��Ŗ|:
�j�։*s�W�}$v|�Ognаkּ+k�K���z��V<�1Y�����M���{z��Wmͼ�>1t�烤v�p�����J~����u~�eշy�~�̪*mUl��<
��l��i���_]����#�;�} �����}�}'TX���F&��v��-F9_��ܚ��͠�u��+�`ε"�I"�:�>�Ϛ�ʪ�>���?69ǽl�T��*�J�Lj�$8��;8�;�y�����������;�� na�9qS'���u��y�����\�������1�4�v�"�<���]��wҦz�4{�T
�l��.��ܺ�Vb���#Ɗ>��Cg�cf%���N�]K���R�o��w�mpLW�V��^��z���=6_��+8�ïζa�|���7}�ښqja��\���]������l{j�`7�3���^]d�N�?ai�~"���2:��h�vU��"��ԯW$��%-�]s�IhdE�Q���(������6^�#��r��
�l�y�qV�v�]};�a������"s8��쫺�Z=���:n��f�5�\oe�V�yN*�ٴ
�e�{���K!�Lnn��>�X�oƩ0#�ׯ��f����L��Z\C ���	��`77Q��]l:��s��ȁv�r�n����(]u�$�*MUp[w�����.'�)t���l��{7��}�݁*+:�� I�NΩ�d�W�]��ɨ�'V%�:��U+sη��6|����9J,*�lUV ��j���³�+7d�������Y�R�F.!U�wk�V���L7M2����Ұ��e���1jTDU��i���ҵ�*ږQ3�Qj�EE�Qr���<�^�딒C'6�/i���������M����k�P?�Py+����p+�Oi`�E3镫�u�.��y�Ej�vR���;�K g_�s-���]tw$Ҹ���a�hVp�/'���u�TM ��/KV]f�.���Iڊ-�Tz��#�Q������t���C�U��ga��5E��.���{�libwd���VZ\�\Nxn�e�Ž��������l�he[�S�$�Aɫ؁��ٕ'���s�`/[n{[�f0��'q��������Sg9�N�݆���E?}��}U��ܲ����^��� ,-=��ګ}�ŰʓQ�.�o;EO8���02gU֕m�Qp�o��6�&;.2�`��9�Cq>�ZA��;�'\��\K|��Y���c�$��^5�5�xø�Oӎ��o#����W��,��r����G/2�v��[gI��ɬ��1
W����g�W��H9O�Uk4���5S!�UcQ[�6%�|�H�yu3����ݼ^a&��=)YB�,��Ջ[{r�pԓ� 5wΉV\p�w�)��!������7%�v��������{��V��r��^����KY�֌#��>�k{2!O�7���W�\���;U}���j�|J���ɳ*P6b����ᰚ��<P�.�IA��nR�8���6���aMHT���՞�G5���4U���~תl�j�˺�:&⹶nȃ��y%��b��F�Mr�ym5����"����܇;���O��,�Y:Ҩ��ɼ���c��\.c��o�o-����/�ewO9FR��*�v�K��]�ͅ	"(��+efh��%T\��k6��{�K�pR���-^N�10q[Kۃ߭�"ƌhj�<�\F���{pp�p�>���_���X"��}�����Q�);��v��o�@�1�E#���=��ٔ�����h^�r=Ojv��/mbH���.�ȶ/5Lr���c"�k^�1'D)=���L����k�z��ۀ��_l�:&�pD���8X���`]7��#[��;뜖�LNԤ��\3[H�ć�>wn(����ܪ�OM��j��֬�1B�doaK".�1짏����!FZ���[���E���Ĥ�~���Z������ ��u�5p�W��b]�����Vy^h��v�&�Cj���|�Q��g���w��k��ա�K����:L�,���o)Բ3���W��t��z�6q;"ZK_4�m�;w�l7�iI���\O�ᔵN�o�V=ī�y�� |��� ̫Kh9����q̷�.L6/�Skd�߱����6wkýj��TR�����G;5=�WΘ�Afk*	&.n��Y�B*���&ֺ$��v����>P�F�5����p*U��ġE��ŋ�����;�VD1K�os�4ࢫUM��v�Z7�%���mk]���<�.=�9��f�ۄ�]-E�b���,Y�ؖ��y�&��m��M�a
}u,E����h�u�+�_Y���9��5�.�;����5�[[(JZ�O��a�ٮ�<4�e�O�F��U}J�D7k5B0kU���'pfT<�s0�������F�v1X{j���eM�Ě 4�!�QY5�����u��r㕱-�Yn87�1("+��E�P�8(�A5j�l�X��i���F�c���1r���11eL�01��M]j��q�j�-��"�\E���%Dr�W*I$ %J���eݎ����I)'&�Y崇��[+���5�C����2�q���cF�����R���]�ֹ�G8}l*7Lfܢ�:�����j���o�QՐ5w�=6���R��*�bT�Z���EO,�^�[L����u��ݍ��bs��I�qH�+7��g�o��}�;z�\;�_�[$�M�����GJ�-��0E�����FK�C#�hrܕ��'g�GNv;F�eJ�%!dc��ս��Le���q55�XgB��U�z��R��Ub��z�ӎ�� �������޴�1���Kea�=`zlzwM��V'o�a��&� x5�y����b���>�4pBNu^��7��dos|R�)�<�o8Uƽ��;���݅���`�_��"���[�-��f�	�^�e.��X4Ǘ��v#��q8��J�;T�y]V^�Jz��N��%{�u�X���爋y����q}�	%L%���<K�6v���]�W�����߂Ö��fO+TM�M�ŋk�2��F�I����(|C佘��
]�n�u�{��x���ڊE0�>�l�oO��ק�
l�x�呃����6R�.���ճsPO�*��ӝt��^u�ZuZ�Z�P����|gnי'rF6�ȝr/M� �u��Ӝgp��ݦ��3���Tܥ�5�M[�O��49�1I�G	m�8�C��Ay{�ރ���ՙZj&�V��65-��.I�9}�[F��Dq�ݐ�CPc�W����V;���NȌ3�x�s=!���YՉ��)�P��U�x��6�D�ص;�QػEQ5�I�u�p�����|۔��,���`�[f���&�`�b���R1�VH���$E=�mUK�`a�b��u
٦���]!���l����$5fyf�d�'��4Al���9#�u0^��'׎��GV������ֽ���}�ۿ<K�P�J�c��kPj8�>�@߬�eXV.��C
���b�#���{��{��u��Q���8?�S��OEZ'U�f���e�΂hE�z�}�����t����_Ml�^�l
�����M5%Di��u�qnP&dbR���εu�&I$0(܁�������_VԜ��A�i�.�����b�g�x2���q����p�qc����NZ����ɵ�4�'��1��y�`إ$��n���U��屙���V-W�E/Ա'�]����r8ax�jNu]H�6T{u�a��|z5w��H�����I�NN�[�a��	ẆD���zb���F�3=������6���'��_z���#@��o6S]��w[�j�BO�
9�9p���[���e_9V�[o��9t��㬮:��V��VQ�{�;�q���t�:�滫ں���f�q��Z橐����1۬ʸ�eYԍv�⺸e�oh�a��]ڧ��w��L*���ՄV�Neۣ��R�v��0����s\��J�N�ut���]�*�fV7((���Q��ggj��b���L4����2��-kvf�ηΥ�w�B�0���
�+��s}Jz�}0k���BP��-7+�F��+r�P�Jn�9��x(5ѭ`�נa�I6�E���?o�+���ڝ{y�in;iY��IXƭ����')��mE�M�2��]�룾ߊu�ݸ�ej�K�0[�K�ۍʡZ�i�QfaMk4�f\�(�Q�ċ�r��$����b1ʸ1�aP���4��A�VLk�h�)Ri��5�&:����8т5.fL���\q�����Ӊ�ߍ�b\���<����:��&�w:���`V���Gt*ظXϱ>s�j��~"��Q�x��V��t=F��z��9�L!L�v��'�M�{I>��P=#Y|;���-[Ҫ��^�q��Jy���+�<j��N�����U�qk�bC���;�k% _�S�W��>it�����D���z$�iŤ�Z3�r�o���ymy{_	���Met��28��{ސz���2*Em���Șd2�p9��m��pR�@N!{xŚ���O�{λ�2�xL�8���7���`W/�t��Oz�h��Ѱy�olDB\������4OY\��F��h駆�+�Z��7|zWk@7�{�+p��N]E˼�<�KV,�J��O����4<E�PYcr>�j�Q�J��r5"e9"��r���w"aoM应�y�R�X$��rN��=zkڇ9�}j���wt�9BqW��h��u�6�3�/
.��6����tY�xz�� �����wC5����tUM{������m��ryF��)�<�QJ���5�PH�|\rMY�.�Gn)m�"wy
#��q�7�����S��g	�l\�w�X�1X\v�t	��yNvJUL}*:=��<6��t�axa�"z��0aՅ��'�%6&�=��^W~�������wT^����T�(8np�݆���I%���vq����ra��7�d����g_��R�G���p塥��<�m��������3Lg�c��Ã@��������<���X�d8��-�����)��C�O=Łi�-mV�s��k�]�8Wi<��v2\3ZH������K�s/x�ͽ���~���j�j����x ם��D����-�j�P�yͮ��x]qИ�/�����e<E�����ߍ+Z�:#��|�q�7�� �$��tTۛ�t�8�]�-ۣD�9RJ<J��Eޘ�n�1���^�nZ���	*.�ׄ��{"�l�^ߕuZ��ٰ�B*�%l�t��Ư�ge^�R�Y0�,���KqF�>�\#���2�����W?/�
��]������7��X#�}Cs2���l�l�0�
0Bِ�褔��ln��;o��9��>�(��������]!�Dfl�j
7-e�����z(r��K}НĠk��3|T�����</d36�`���̈�7muZ��4�6�}M�9{����{�
q��k�Bs7O"�L�	�nb-9�Qj䏷�.)8xmyհ�h�Z�.�1�N�P:�!��%�5�jg!fP@���'aGM;��Mv�P�-�ee��"�\t��<9C��
�Wq�n
C��c��<����^���^�+s�3q�ԙ������`��B��C��IԺ�@
��,_a��h�맴����x�A����1�)V5}}w}j�Wj�R���j7Y$����`�js��T�9]\�@T委�W�ln��
tʀS�(ВNs�:�"0�@o>y��s�'�R�Ӏ��mp���L-v�Vr������/;��[�[ohN�i�R�'L7�vn�;2p�2�����L�(sy��ȱu�ulz�G>��뼔��b`����$�q9zp98v-b�����}���Ϧ� �wM��m]md���.�Q^+.�Z6�U��]WϤ�)]٣2⼼"n;��I�'ne�*efl=a!.�����6�]e����dz�0̕���T\s0q�-cj'v��)��Z�"�.C)r��U����Mf�Mf[����[1��)Aƙf`Q2�ܦ��hQ[q̩s1F�ƶ�@!P)�1�	��V���ݡL��W~���H�1U齰8��{�9�Q����!��R�w��~"�V��Ր����hq�E��#p�@�5s��T@�ޠ����Ti��,ۥb'�*1K�Fz��v���u,�� y2��2��nt�v�rcѐɩ�e������=
�0��eY��<��V�X�|�o�$�r�zt�i3��_a���.94���He���z�+���㐄�ɱ�L�*�"��m��g'Vx�uԜ�V�c(�� �n��tl��rMC!W��1��>RBp�B�j@xrZt/���k����kid8�:o���[��k�UyF�*a�VTi/��+`��3���WE2��`�|�g;1�A:"v�|d��`É)ޚ.��^�V�����{mu6�9�|���l�'ݸ����9:v�{�ǥ�A���2q0����ZjM�_����2
{<��v�X�<��� ��*i5}���F�����Lq�SEh�당^���nmJ�4-��[�]��u��m�㥇<*�C�Bg�)C��1��zIn#xt�Z�H`�]�� X�W��9��H'�G�\6��];��s}v��x��O����Z,�E��v5l$}��䇗�m���=h��ga�y+�<��c4�I�k���L���CQ(ᛋu�zj]Z�QEI��Vt���{�Ⱥ7����I��ެ9vB퓉B��Y�f�
[��4+��<a�Ь�:�ļ�4�-�8N��F���y�Ii[���h�z�n�'�nVO�15q��`�8X���ݝ��VVJ����9��"�B�r'8�7zwI�u�WY����9�h;a/*}�b���� 	�l�U��wJ۴!��N�1�ʊ��
�Y�f��*� �<��n����S-J�žk�/g�ϖ�{�TC��N'Ay�/Z=|v�)���Vϓ^�\aB�Gݻy۰Ƀ0����0h}A�g���q��8�.ӌ�CI�C}�ך�q��L���o�u��;��[�uM2�걠��p��י*����#?m�V�s��;ɿ�+�Ƹ��Ʋ��pol�k�t'-�t��=3}h�u��z5�*m�t��awK垻N�t�1���N�7��SO������Qgo���mh� �� ��k��^ЂJʾ������Y�i�B��N7��)�W�;aߖhc���om)՜�/��i�����q�L�Ӭ�S���pN{����_PV�e���ϫ�Ɖf���4!�Sn8x�֋S�|i�a���J`Um��1��,U!V+e������
0�|�-U��kv���V�U����:�YA+�w��oZ�*��Bf��]v���Ow}<�L�a�İ~����ix��I�M��%���'$���q�M5�y�Iחᕛ��SxUƨ�� �)ٻ<>bi�+a���1U�{��ֲ�,}8�+��AO֨
\jƾ��Ph���H}]"�W�4T[ӗf
�0S���*
�m��f��v��NҾ'��4��<�����{H)���>0�`�-o�5HP+�j��������͙_1 ���4�q�r]=mؼa�Y=Ls��7�O�}��@�_�T��R������G-?/������Y�$�&���'��3z%&e���Ϳ���}��=�Gˣ+�xHHB�PL� z �	ju�7H|�x��a?N�O��ф��R_hx})�  I��� y���S��_����>}d�g��?�Òof����5I�F�D�������9�����(Gf��a������@��d=���<�k�}��a"H}�$��@��#�� I��l��#&�������h}����<	��������o��'����8O��OȐi��@w��~���'��*�dο�d2 o�r~�g?��}��	�̻�@��֤��� $�}?\��~'�~�÷�4~�	�8D����O��,�${�xɮ���]�萐�(H���<6 <&]*�y��+�	s?/������9�����@}�8��d�����?�_��G>s���@5
}������������d��'�D����O�|�����������>_x2�M�2�h8C����y������Y8j��'ϟU��
'P��_���N}���x��!�O��'ϰ��F|�~G??���ȝL�HO�>�#����Q�����;�'x)�𧿻�Ϻ�}$ I�8O� 	?����'��� ~-%�����Q~ZО���܇��ђB$�p�qĞ�Ƀ������$	D6X:�`p:8��zn9��`���$6���?p3a�F�k����MBO$�|�������d8@:��� �R2G�?g�I� C�?)?����>@�����?��Q�����V?��C�>�O���O����C�>�g��g����M@}��>������� /�!iHO������ 	,���r~�=�?��@����}�#����>�D��a�?Hp�:�8r��`1&�ￇЄ���O݁��^~ x$���������w�S�I��~��O��p�$�>�d�=� ����>�>��C�?wp�|�'�T'��jJ$�S������h!I�`n@� }(D$��d�?@�}D��#�O�~��:�~���}�>���N�\����8M�<%��!������6p�E�}�'��?��'��:����"�(Hdı�