BZh91AY&SY:w����߀@q���b� ����bD��� $(�                                      
��QAl2���$) P (� �5�h2
�H	(PE �4UJ��*��TA	
U QBA��H	
�EUT�TA�
�B�
$$  R����P��@@���(
  UP$�(��
(u��BH�J �  �}G�E�W#l5@::W`���ThӮۧAk۬��U�4QĶ�4mҺ ���45AE"*�x   m^��V�AI�V�[i*U��L�*���㫺
���Ʈ�QJ�8\ֲ�)WY�%[jR�;�.���Us]�1E`��;jMcu*ARH)GF�PJ��  b;�[i�5��]�QF�JL뎻jWM)ӛ�*�BGqZ檒�J\��oj[j�*��s��J�)�,:B�.��+�zN�%^9{��)J�
��"�T� QJ�  ��
6�Y\��5�[V��K�[��OT�M��7�z*�{S[<�x�
R�N�����ʥR^��{�RUIC��޽�P�*�V�nvզ��`�w^�)Zji�uA@(IUQP
�(��   Z�-�����)
���7P[jض���:[Mi�N�vմ�s��j��V��Jm�2����Y-�:��Ԭ�
NpZ��3�D��Ɛ6���� �   {u��+:Ҷ��hU�;��T��i0୵),��Zڲ�kt���e�[m���*�jWp:�4�S���Ց�ZguWq6ʫj�p:�D��TPT �   ��V�ղ�qm��ԕmʷJ��k5�uK�k*�V�R�����U ���+�-e6�V蛨Gks���Uڝ��
3@PP
*�JIJ��W�  �u�����˫�5��:�5Uv�j�%TZ�QWmkV�Sp5�l\����V쫵Ѡ�'Rj��Z�R���ґ�R�I
"��  tx���(�euR��Y$��6�W@���jUS�[��v��.(Uw93�T�tuu�Up!H�UT�D����W�  1ށ��l�]u�D�5Q@�
�EmUcB�SCQ]4�v�iU�:KUU�N��cT�T����   @�  j`�J��  � L "�႒��� 04� �)4�OI����16��B)�)*� d    � 
���1      z���UD�4�� ��  ���򏑾�$|��D"�S?-���͓��9 �]ӭ}[��j�acSs�w�   ���׊
���d�Us�g�� ��m'�k���徧� ���Ӏ���U���W�M��#mV�����6�2�x�/$�Y��g���9��V��k�6����V���٭}�~���Z�*����ٵ}���+_ek�}����3U�V�ͫ춾���Z�5��+_ek�ھ��m���٭}�Wٵ}�����V��ھ�k�۶��Z�6����V�ʷ�j�*��W����L��j��Wٵ}�W�j�-_e��}���U�lͯ�U�j��W�j�-_e���`,��X�p�E��*l�%�ȋ��.o�֭�kU��Z�٭����վ�j��m]��Wٶ�_em[쭶�͵[쭶�ͪ��[V�+U���V�5L�m}���eUo��m}��o�V��U���@�b��X��\��4�k[}�����U_f���k}����Z��ͫ�ֵ��ַ٫[}�V�������[o�ڪ�5ko�[m�����Z���[}�A��C��.VIM�%NV[U3j�ekk�ֶ�6��j�*�ͫ��}�����Z��fW�Z�-_e��}��٭}�W�j�5����ٛWٵ}�Wٵ}��ٶ�ͫ�־��ٷ���f�ٵ}�����V��W�Z�6��j�6����ھͫٶ�������7��ǝ�̽��1�Pf��;v�	Eo�sbDõ��}��*=�d9�T�1�.F	�U+�Év.옞�wl�Y.�xJ;t���̠܆7���o��n�U#r�ky
˼�=��5����V��MQ���]�2[0v$�#��vί77G�}^�s޹�?x�ɝk�}�>�`C�l���ʴ8;�x�9b��PksxfB<gb�(Q��/�"e��6�.����=�(j���5�3w�xk�h�J�^�%�F)��~��D��gV��);%ǧ6غ�0l�e�V��)������\l�Y���;)��r��(	j ���ue����qt�w큮T�Ҿy8]�;ke��[c�����m}�v��7�$m���o7���Qy�d�̋:n�p�ű�=*O�xry�J�xNQݷV�7Nͯ����'�zwwHDm�l����=	�f���#q��Yې��)��6R��`�t~#��������G
�5��.��(:���y�r<Y�SrD�no]<����dԮ�5�.������k��F&1�U�qS�,`��w��Ѡ�n�����9wo<��*�o]$Pe*'v��oE����9����b}8����xa�8��0�������r�����/;�.cs�����j��7z��E��m�m�\���R�޺7�
zY�Z^�W��}�nk��=�p�$�9�(흯g*�XGg3�,��-��qp���ō�L�YݵP��1��\;���,�a�~���,}@�.vX�۠�iv��|��s{�j^|��C���+\�s`���J�n�&L�d�C[Kn�@.-����{.��+8n)�N̡Di��8`+ۥ���k�O���0ٓ����̓�ܠvU�3�{Uw�%�E0�-��G�Ap�~	,X}/��� Sی���F����qЫ줲7s���]�XJ�f*����Z�!���:�;ϰ�ʐ*��qygvn�����UX��Sbyl1���~l��ᰎEZ��<C���WE�� nk�!�Y�2��>Rvj��Gn/��3Xшީ� 2m�.,�E��6|:�m�(�:ݔ�hB=,nj�WČ���/d}.j�g�Gd⇙Q%NkӆA;���3��v�����	�B�n���Y�t�k[P+[�j�8�\gu+sG�w,Oܣ������cӳ��M /^����	�f�u��u�Eۿ���q�9����fh��8^(�ۉ(��ޑ63�����n��5Ԉ�����Q��s�!wIZu�mg{pg5��w=�j�sN�;Z�6�̥��y�Ͷ�y��6�ڦ�j���Y�ym�s9�FW�Q�I&��z2��pq<eـ�r'��z�0�'} {��Rs.���5x�5�5��!z�z=�P��3j�)����s���5v����%� ��ec��ƃ�CA��`��`��,I��pHNpuŶ!ÎE�#ͫ�l,q�2��7�U0eZ��|zMW/ȩڷ��z�|��Ժ�u ��Y�O��Q��=���vk'��O-s9��r�1E1j}r晫M��5"�%Tu�Ôg'�R�:���w%��4��P�H��{�wgkw}���º��_�\G���g7��"� J�������m�|�M�c����@��{41�8�0Vqn���w6�6<y(�Xށ�g6�y�4̹Ϧ�u���-9��Xa�m�/j�*�ι�qz���W�Wn�5ՌkK�M�EQ�ٛ��l��^����wA��c��C��@,��M��j���r�B�{�'���z;Vt]�Fo�]�,�Q �S��jr�p��(%c���@�\��.�	k����ᒺ�����.Y�:>ڄ�F�Y�^Ι�aXd���+h�Î�}��+{�c����9s/��8G� e&��]�{��B�Mӽ)�5���uj�RVpck�Y-�5� (��s^\�cO���@�F�iƎ�u��O �\vZ7x�����8,]�^����i�P9��*�Z��쒙8��3n���#����I�rc�����'�����q�w5�����:��rQ������ ��AO��^%1��ҁ���S`w�|b��.^�9�N=�x����5��WV,:3�=ݻ dK��9�a�0ݘ��N��S&� t��g{�7f1�7m��!��X�����Gu�>�oi�߶v��25��2�)f�ó�{�wqE��3WN	���j�A�;��@��䷵ji��K÷���%�m�.����4H��+2f�CZ�bZE@�pe-�b�BFú��a0��͍ɯ�;���緊��-jһ74j�Z��"�v$;�)�lMΫCg.QT���󹸵FK	�is���r�.T� 3f|�,١jvǧ���+b��&�=����ӕ�F�>����:F�>|�n�]M�f�In��j����#��a�������z>�^h�y�\g�k��D[��`��N���G�ֹi�����PN����8o(����gsy �amc���xi�����'Cz;��*�/�N&�,�D1�t���͒�a 3q��`{4���2q�+��&&�G$��{(RͲ�Z���dʵÄ�!\M��wP��9ї;K��_������	I���M�;L�!���+T��4��h���3�ޡ�H�4��OmU�1>Ғ�޻Z��qk]ls��8v�7!��#︷��8����ٺ�Ɋ�ǵ�;���ZJ����₾�����s���1}����x;S�5��e���뜡ydzNֹ&�%w[�iI��^�#�'&�X�}��G+�ض��t�`���t�ty�խ���#K�b�|��u��8�B�kr���n7��d��q���n�x�q8~��Xy��m�Ty�\�p�i�>ݽ��2�ݐ��g.i�C��	�$��󻃜��'h�	(�:�G���F��ږ#
�G&�f�z�&�ܒ��n�{	�u\��7'q��u�u�v��������.��z'Էm��I_����='f��,,=p<���	����ˁd�$)F�8[z������횳x�'#���W�[�]�J�fODsvT�p���k�Q�8��!3�w"nW^�&m[�YӁ�825u��� ����zYg�ܗC+�s*;a�kY2Ƕ��;>��m�# �-�.��YZ�:��������J��w
���Tq��Q��;�y�=���7���*��qhb�V���3�Fl�2���{W���X��gC����G8,�w�rnv�ܼz��7����oi�Ǘl�����F��\.��>�z�E���Jλ�ԷhVVuaa�����`I�Ty�@�9��,������ޛ�z��'mR)���N��b�yx|�y�l%5�N�zM��h��w5,�ľv�r��XfꄥmG\s,ç�F��d�bZN��1���Ϸ7���y0n�.�ur�"ː�dއD�ȱ�pr��r�ql��Np����y�.����3f���H��a��Ӵ���`\]�.{^�u�r��*��!V$5vШ�:$�+vv�QKS�FN���^Si
;�}V��n�'�1e�"	^��rS݆�o�밢DuݿN�n���f��P�6��f�^p���2>Z��^{�b�N�o5��2��q=y���r��˥��ݘ҈�gG���m��.�;��Gtˍ�Ѭ?�ll��԰��ڷ'V�Q����+x��Çc���� XxԖ�{�nV������'	4y�oW-?���Yf��# ד��77i������C��C�.�q��<�Ոf�i�1�܄��X9<�z�Hˮˮ[s\�3�#6w�pr���y��8-x��>Lt�:���Ń;���gZo��Q6h%Z��]���:��Ϟ�wj�lX8=����fB�}��59��Y�f�-���<<��5�+��+ �aZ�Az��4�RX��L�)�
��1�"]1^��LU�;z���c����\�<{V��z��,7P��n]\@c����.��<C}�V�(���(�J|&�^-ku,�[�,�,�Ӹ�9�O� �a=�t����}�TᯚR��wu���Y�T�x���'O�K�'���F�P��Y�7��:w�.��������e;_m�5;��k�i'����Q�Drp��:��8�M�I�krd�My2�����]����gw='���U�պk׼*|gc��6���]�P7]EX
|2�F�p�}�^z�o�nv�v���bӴ�s�p��s�99f���-��um��(^�'e��GH:'�v�oR,Zq�w+fr���	N�Q���㸖�i�ZV��a�k8���[s~�tDtM�9����FK�%�.���3x�h�y�����;'E�z��1(fW$δU��^Qp,{�.{�Z�\B�q{�|�Þ�T+ղd��p�ⷓ��$3��y�מkt��\�u	h,bzǹ����tא�8�k �3�n��N��$�1�i]���.�1�<-�qo=5>���K�v��p��Z�t�nv��]9�/J=��B�r�{�&go�r`$-��$�a�[9���,U\�������U\t�#�����X3�[�:m�6��㔝�nn���#�hk��
LL[��]���t�H>AȺ��J��H� �ؕ�������i&B2��p�w�n�Kt�7r��"�w
��#vS�J�.੸t9����sD��O	�4�뒓�k&�8���u��:x�q�x�|�`q	N�9�	��f�ԣBBGɈ�`V�4����N�?ub�Z�i��bԧE�q�O��<DI�׏`�� ;s�p���0��u�mE��/^�ċ���7vL5�eǧ���7F��䇯nR��)��V���Ԃ�KM
@1��,��ɹPcs ۜt
U`\]×Gc�2�Do��ٳ7p����fX��)�N�Fƫ�7�w�a�i0Gb���;63��Y��0��֬�b+j�iڞ��K8��<A_W�(UM�,y�y�:=��'�GRw���M�{��M��]T˨�<-w���A����pэ��B���ɡ|��D�D�����Bl�\�]������ye��e���[ot`��qn�Z��*�z�/l������P�p���~X�J�8����겑d��wA�p�2b8�]f���X�������*��kX0�Ѝ���:9�+8UH ����P�M����_`��f�A]�]�0��D�3�4�������ރ7ly�i띐�vS��`>����:��a�F�.�}��{ ��Ƽ6��p���{���i}��u�<��W��Jo@��,}���_.����N�dg��G<2��V�F�V[��ɴ7\��}��v�F��xh�zdtͽ�7���m�!��M��#��o֧�����D����̉�Eyb��}�7�ݬ�c.��� �x�j��O}��/܇lj^E�0 3{���,����i�T�s]�tˣ���@�!㺍%�8�hX饨�����a�ᮬ���ŧ�Pi���)g���ƙ9c�튳��++���\��G@�z����q�*���єާ[�S�ud�Ԧ)�:�.�ζ�P��%�}.�+�xe�^�rt]��x���������I���o0�Ѡ��=�.�z%�2�-ZX�pp-]k�.W��R�Yˠ�N��Z�I1�-�������NZ�r�ۤVa{@n�((rBwA �����Ȳ:��/�9�,=�X�-B��
ΐʹ�N���hypJ�	�0�Lf����pP�[2�t�]����Z��g��H�O>�t#C�9��	���;=n�d=���P7Z��:��7��!�W߬�r�ʌdFj{!w�Ov��Y���>����w���/�wk/�l'����v�ס��:
뢔'<b�(/4�+�dh�a�:؁�����0==�w[&��[ 
�!���ť+��Lɑ��[�;��`(��r�0�p��^8�x����GG��[q�gA8���M1�vt�i0Vp�1f��kt)*�tU�{,/m�]x��Ӧvn���F��R%ף!b�zr����Pb��yoo	�
j�06��ǔ�S�!�nǀY�G�@5�>g�݄k�yh&$:>����:I��N��WGh���X6mc{s���q�\��Z#=��:<w7y�=���4ZH���w��p˚+z��l�.t��v����TT0�~^´Ǫ���.%��jnqZ��w)�ꈖ�D��7��P��;�4S7/j9r��G�KWCb8B� �-)2�B�뷾=ӷ�Q��A������4ޫPґ�	iK� ��´f���1�)ر�Y���Ʊ!�!=Zodc����ݖ�a�U�'�DJ�V���+]�/Jp9�ݬ��y�c�H����w�#�D��!8+-��%5�M[}7���q�VnXC��������x+X����x�>e{�~Ӵ���d��i��֪�:L��d"�����Z���i�7�1�L{�7z��fo�R�`�_�d��Kݔ�ϳ�-D��B=������7;ox�;��x�|��I�K��L�l���hG�,���<oS�=�q|_��h�O:L�x�ece�ө�+�k^��lӇD��1o(��Ѕ��y���f�3iпC4�,M��n>=�T�sz�x��������0�����u������Q�͜jr	u��;F�ݥ�s͒��_#�c�o[��/����v��xg"ڳt/5<�{��n	�P�e��7.#g-����̂
T���ۆ-!u���LO�X�޻��fr崍�'i�΋�ʴ�r+�br�q���W_<r{#�yg�s��ϛo�=���W�Os=��y�6Fl������u�v{�a���4�jv���k�@]ó[�򴲾{��h���^˭�qwtG�����kL�����dg��b��r:k�v_z&�u��DO���O�����O�r[/����o���a8�ק9pX^��H#�ٳ�q�����R�.�ʺ��>�k���nG�����{s��op�)�����j��L��v����s>�7�/��}�n����8�����v[��F�7"C���U-�B��v�p�]d�������[ɫm�}�2PJ�{��;�4m��d%lkviG��([6���l�(qZ39N�h�r��I���yΓp�+��ts��Np�9p��u=Ӯf�n�S�~�k�Y�G@�g�b��$L��.#w��!Mw���"�f&�g�3�X��KR�1�bᅽy��o�y.��Q��J�{Lro�o���7�������|��%�O ��W�����_X�3@�#���n{v���&�]���M��c�r-ۙ[o�隲L��g���й��|f���ܲH��o�S�y�l.�վ��:� =�x�S�M?F{��>֫�i<䚛��rz�9��pI����Z��O������Ue,��N��<��J�<��s �g#ŎO��Gf0�2nזIN�_�!���Z��`H˜�p���ٮξѓ�u���7D�W;V@3�ޞ^���f���7`[�b
9�=9t5�[/�/�l�f���*�����x�X����U{�⠤���Xs�k�=?q|�݇�r��e��Gtkn�C1�GM-|���'��o�a�^�y�{(�1\�/L�Z��6j��ǞW[I#��vD+e{�	��ar6���2�ʢn{��6&V���F��N�;���V����u�ۆHD]#s��������<k򙽐a��*n�����=#�/|����ޥ�5�t8$,�4���k��^�}nk���0�]�I�A`���`c=��9!��Z�dǓWb���%@im�)(�{��.b�bɒ���
���M��C��'a����z��8�Kߩ[�t���CË:#Wqξ&��rI���`/G�GT�:���e����+��Tq����!68�pX�h_k_�HS8-u���Z��|ߙ|VN�2���f�읋v��(�.]aK!��b��;����V<˧�L��g�Ǻ%-K�{��=�{����hK��A�r���Oj��&�Vn����p��XM�l٬ݠ�Nte79���Ve�]C)v��L������������o��<;���l���3}_K|��������bc���{e�ٹ�P�f�}�[�|E�Q]а��B�^�^̜�*���SWg��!!=|��u=mV���TG^e�[�xr.�A��݊�����&h�-�t��@��B�|�na�x�o&��v46�l� f�i0ԗ�"f�_:�stO��Z��m1Yks�n�l�1���i�7ဝ��*p���G��{{�`|f��Ȼ`��gj�o����x��G��K��aw�)��-�������;�%�˻./= �y����Z�78_pEL���,�j��*}��àtS��O"�{~�wz��iZy�U���흾&�{�k�y�.��i���e�16���R �ºZ�|y�Df�&�A�Y-��i0��{^{�� ��7�6�!�?!܉zcd��d���S��_mNlR��n:{n��7���,7�A��p�DQlBI�~⽇<6��Fx�jް�s��gxzx�����XVq;���.�.q�+���z�䙭��.�ͣ�uu��4a�5�9�p��ihܐ<;n͐Xu*��r�I�^/	~ �=޸���x���}���5��u�z �O��6�}7��5�2���էo�7��;�<{p�Hr�;<��-��6,9���}���r!-�<t�,J\^M�<cݾ�qpw�]��hC׸l�r<o�'�Έo�zx�+��_Es���>`L�7t��Yї#�:{�r��G���l��9��qQ0߯�(V�y���Ƶ/�~aN}:�<�>P��3��[��wjT�O���#ؽ��<L�ҽ�V��Xm���K��"�^q���5����Bӵ��3���W�W��Y LVK�r�c���M������;=�9/����BƄ�}@>��Uy_�����%ּ��c�;�l���u�=te!���9���Y+������̪�]�E�+/g�"�%�D*��'�gg��������ǽ��9�A��m��X�9�a�L��(�ʈ|oT����`w\fYܣ�6L�"�s����0�#:��:d\a��s�|S�=��穤d3ؼ��z3ϻ��{v��po�}m�+r?
�n�����g�"���]��\ʭ���zzo���:ڃ�·�=��n2�y7k��du���ez#��/^�d�]��OFˬh]�<�% oьjЉ�ku�l�؟(���]�Ǽ�܈�0�^�[��N��������6C��%^��mK�u���O�6ׯ�]*K<���S( �өH�W��yQS[vm&�b�+��T+&r��Թ�� )���BgE{a�>k��}6L�8]��A֥�sP"ܨ��b��+���Oo��N���Y�2&:�cQ���.�ڊ�=��13x�I>qA7Ď��������C�&�lQ�g��,��T��bs���5�H��᎝�)ʳ{ȓ�y��P�W;r?�����y?|�h�$�(��I��ǽ�O�]ѳ�k�6����m�и�\�Fۂ�<X&�z��k}^�=��gK����:s�7��-�w����]9�����U�L�%P���Nz"D�V^�w˚����6i�L1�)V2��ILɆV/�
�:R�_f���P_]
!l"(�c�0e$�Jغ�ΣM�Ȱ <zqy��q}����	�x��R��\�����P�&�d���pg�b��*!�V��ӛD=ixzn��IG|զʳ{�[��r5�Ȉ7�db�,DERw{�NV,G2�����RK
��n�x����u�ǬC���ǉ�p��k�=3s���������H����	}��a\�+Ѐ��tj�;A�t/^{���N���o�8��fk{�o��Rz|b�\�̒��ޭ6Udt�W@����7�u�d;|E:�>��46���i9b��oὊyL�ۜZl���K�6l��>���G&;�f���ʹ��W��ͳ��z8�I����T�<'��/�u#���u���1���X޻�:��0�#o4b��u���[o�t���)��n���2N�A�'8� }'R���3�,�[}�Iڇ3t�b�Y�7Ǡ�������bC��XN��yY��Ǘ���}O,�vl�G�� |�Q轷#MK��|��7�3�w�����{�n0Mbb�E}P<�թ�����HN�R#�A����ɖ�~���g�����2a�^l�.�^�|T�˫1�%u���K[Z�_g^Z�sb�w6��X��*|h#�:Ϭ��d���Cڹy�3sG�ܘҘmq/bur�N9&_R��겵���hc}�.Ŗv����	S�4�4���2��OE��;FTW��6���|/�Y�xxf�NNn8�2�]=z�_+�W%Ҷ��jd����J�Z��Cʕ�)�(m�w��6U�8��xz�7�2��齶�uI]࣪9/����BM:� �![�GY�M�#N���d*�ꖅ�fTq�#�6����U�Jyy�1+"��KD�(���bL��9�K��.�ԗ�xj�C�ҫxbL��n�:ǳ�Ϗz-��d�ᢰ�V/���+�w����5|�X�h�8�߲�:�j;�0��KX���5�T���v�kC����b�:���3�˸�7���ٳ<���q:�c(�+��/�2�"�	\�Z���O�ZX���h¶[��غ[�Wuu��zT�.��ۂR�*c5��wt������:C�#�:�i �^���/L^9�l��͔^���3�8ĸtg$���aX��PE����E͎nV�)�X���М���)�!�n����y��C��Tr�����F�9�a
�!>�s���l�p0��^p�>~��g���O+�cy5�`h�sjVJy���m��oT͈PFo���oOc34�.3ǳ{=�E�jHoH�E�l~c�;u,cĘ�;��v}s�,����'�{�?%��>�㧷�ۛ��iXt���x��e�Ӄ�U0u����{ӵ�;Yv�<�=�H�N���]]�ص�oo�p�<���ye���P���8�]���n����ہ�i�ܻ +�St%�o���iN;3˰D����9�r���bfK�9ݻ�r��nV���C#Wa;G&��_���;�S�=�$�N^�лN� Y����M۵o������k҇�ѭq�>$��=�����9�c��������>�<�jӉ�������m�P!�x��}�&�JL܋����yRJz����R��U�i��V�޻�9e97�vmM;�����J�f��j1�n�ZF�0"0=65�V��@N#�\>��RH��1�<ܜP���*u��z���zx٩��{4{٢t�C�6�[ا�cY���g��8���j��� t����a��͞�9�=�C��塟�}���ݦ�z�sx`S&�??w��[�~�l��pXx#�'j��aF�Jfz�#+A[�|�E� 7<���<��sC�w������]W8�2�,�gs��;߻`3y�$k��|�P��r'S1��Y��L�J:n�nLy$Y�x�8_+���3w���S��N�Ž��!���j#�^��͘0g��w�U�`*�4�ɓlmEI@��I�g���q/]���E���%��
��^vp��5�5��(g�c�{C�{"�[�� �ޱ��{�񷱯N>��|�/*��W7C`�YF�l�xEZN�
��s�2Kk�����K��{��䨽/%d�ӭ�3\Sw&`y�e��Ϊ!��S�#��ta��G��_L����E�Ֆ���}�Z	W*��#N��&��yZ�?L^|�5n��h�������v�]��5�3ӽWw������zK���{�ՍJ8bo}ݹ���M��8j���ս�xdc6�7�k�^Q�Ā�y-9��۝�g?/C�Gݕuؖu٥+�0%�Z��a�I�!�;7H���h��rN��҈��[7@���Z�ެ=��Y�滷�>ע@Ah0�I�u������N<cO]Gx�?��6ݧ��p驗ovKz.�h@��^��6\���Ģ2�P���O���9\�퐇V%����L�F�/�q��]�"���ڝq���.Ma��i��8�n{�{�!�0��٪�|���T�Y���F�Θ�y�j�c��2��w�����{%A����T[�����!��,�������հ��q����,�#��1��j�ۆ���`Zub��Ke�R���	�Y!T��ɓ�99�MKEt�G�Z�.�(=x��~�l�5C}���uo��TZiW�b�����pkF-�n\��ה��j�ePu<�K��C�a"{;y}�N>i���Ǥ��z�m#�Ӧ�覰�M�_w{gr��ԑ��uwX[���=k�̀�k��{�bo�uA2�u�vo.����'C�K3�Eƻ*Z�*^�����I�F�5Y+	�y�%�ח��VIb1X��Ļ�I��t�$�]��~����i�b\�.������#�s:��e?{x��v��V�� <�%�yת4�s#��54R>}3�ϩ�l�t>�F�Kl0�vC˄K�x�u��:�3��M�B"�}:���[����Ӧi�K���ʌa���;���R{�gr���Z�)L�O{����&db�U�=�Ӣ��
�g���p�=��<�*��k>��YP.�B,�h�Qa}7x[��R�������>��5�v�p����f��V�Cu=�����x�=�c*f�0�HuD�rG���c�v%OҴ��w�Z��{_b��κ�j�P4��md�w7*�;���uM�E���XO�|�{�&��ٳ�5��w���m�vP
-�nE�����]�Ý��0}}�9�It���Y�;؈tGu�e����
�����g죗��:����jM�~k+�C	�{(�[�U�����~d,�cw=�m(ϮH5yeZt��ݪ�"���Ͻ{����r��P���7}*'[��g�̤,�i�#���s�cA���y�����%�½�<.t�t�G�;�A�l�S�ޮwb���;��g`��~��:��T��*-O����U�̭]ʱT�	8H�p�kӹ��)5�UOg��u�v#/��'�3��C�,%!<����:�P!�<f�n ���3P�F�={�Z
�2b�H�r���\�^�:���}��1.Ӟ&k_^�im�������дM!_�ۨ@���v�oI�
-�=ȟ�ޥx/��M��Lvx�<�v����"r�>�8����I/'C��R;��<��Ne�"I䲕�m���O�_"�>ė<̌��j�	ծ4g�f�!�}���̤��`��{�y�b ����Ps�31��π�#��>��pC����<>�9�~�>�5gSG�j��;����|`�q��H�aA��[�f��y0��?��R�wv>��jAog,g���}�1��_���uvgf���6k�vݺs��ӆ���ٮ�����٧e>t���=ۥN���H�ָ�"����S̏��'Qu�O��ٞG�X�h��~�d�H���8�#YJ�VcK�L����v�7�*A��w"�`a),�޴V��2:IWk�T�G��+����F�� �f�	�X����ty�s��&��o��"z�����8���9�{��ص��wN<;칋���(Jx�.��2u�;^{��X;����4�]�����x�+X	��nMYjG#�k�[�oq�ߚ�S���S�C���W���y�k��XM�=p�ZjQѺ�e���;s5H�l2�l��(ok�����X��kb!�����ԫ����hI�^�E�p.����JY�{4T���=�2�#�$�L��85�k�$�dI�j���i�
m��Lv�j��jt�N�bh�94�=�)2VU���k�+�'@P���6��+[+��X5<X�;V�~�p���4ڠt\<7����#�/P7X�:���ciypj���V^G���ǽD�����b�>����c���қ�B=0�'ug��Ⱦ<'�v1����n\��ݾ�|sB�FS(���y��Z@�/��9�/7��{[�#�v5�x����ze;��Xpz>�݆{��z;���'��xݪiܛ{QJs�D�u�H]�Q�6��*@{\�ӡ�~�(����u��)�3̓�����c�����͚*T,ɩ�(9g��ճvnj�h��BIx]<�k14^�ⵀH�ٛ���㲵��_�v�T����Kz<�24v�޸�+��x�>a�~,��D����KVI�e��,�`�Nhq>8\���x��w����T��>��y�J�o�\{V,�ǧ�ځ�/_C�t3�5����4e	�Ca���ܵ�nK}�~���3r�C�{>�0�a�(��'Ը)B.p\��\]�N�k�n���f��5a^5Y|�ތ`'a���+НP41�&�/r�.XJƄa^U�%���R�s����S�{݇dI'pw��k�
��4釽��Ãlgz�*��s5&l���#]\�r���?h�I)T�u<N�S�YV;�d\�PcHHk�}<��g���F�tn�FOF����=�9WN���������[<O]K7�F�u�i�zP)�~d�J�?o%�v��E���8f˿k8`V7��1x����(��y'A�u��ξZ�/�P��
=��LNZ���y�?�f\�����G��@��>б����J-��"X|V4�B�{�M�^~�9�6z��p_���|�hon66 f6
����RTH��n�XK���U�7&�΁xN�X$���
o�|�p���3��cx��C0�f�|�˦jc;�R�M�6MMu���ɖ/qos��t<0=��O��8t-�6�̨�V�oikDu�t���:z�G��L��__X����D���'W�b��Gm�<�G!ܗ|�75�>^5�|a_�s����lc�WyxyƎV4]i�Eg��7,s�%>e�k�������)��Z �p��%�Bp���>׌�&Jb&jk�W��Wkh��*�P@/�ܳ���6R������������}�<�&��N�����^�H�Q��e��:c���m2�jt��9Jˋ2��ME-溌il�6��n��;�g�f �k9ɳ��~��ۅ	� 2o��l��2罢�]D�`z�c����W�m��Af�c^��",��y\�60���i��2��xT�Ī�!dOZ����q�+E��tb;٫W�/>���R�"v�kxU�>&�lݓ��t�~'�i�u�5�ڜ��������]̧�ۑ�H��և-?;�/tZ[/�U��>�������8f�T�7:�u]����+��Du�X���M"[r�Ӽq$sZ{$�`��o5��[ǻ]s+j{��4,o1�$�L��)BmwՍ:Y�+o^9�SRå�l��-�ڔ�]� ����;��ݑ��4��j���u�ZG�t`O�{���{Oj�����t2V�iv�>�{/�����gC��e����!���9]t놘S�n4@��u����q-������Ӥ�g<s��%��Y���lzJ e�e���0:<����(�o.�鱄�2�8��ٴ���Ԋ����=Յ`#e����w���~��tR5h.q�gv��=�w`��}��y�D"�����^��ac���:���g`�g�+�T�s�90\��SS\�T��B�\B]��Uҷ �`���bb����_N�eo���ó�ᐓ鞘-д��]��LG�����J���b|ʴ%�嗌����\�Gt��]�x\D����F�13r��.oa�L���`�`%�ʙ�N�R��-�3]zA�ٷgM�vl�֣�혴��o�;O���B�G޼���^��|�������d~���1ܝ�1�;ȯcj2{r�>TQd˝�4���f����m�9������"s^�������������K
׉dv��0Uڡ�]�r�y{�(&�Z�
�i9n��
N3�6�p,�Hdǻ��$md~���{*�0�.�#]�n����w�u.��#ה9҆�R1(˚bCh����
��i�{.�V��n��m�y��ړg�:�j���Jɵ�=޲��zy)u,l9lY����Ʋ�N<�إrE�%���_wE�é�wq­��R�ʻ���A�R�zz��T����R�T箻M�׭���Y����;J��\��9Qˣ�낏�GG��0�î��{^mÝQ�k��5W݉p�O6�7�e�=lC*�rPz=s8v�4.�8�s�b;wv�w��oa}����h��r�g�<$՚����L��u�3���fy��d�N���{9o*B}�۸�����K˲C��73�W����l�[׌[��F/{6I�y�/���ШC�5�ِE�}�w7Ø��]�sʝ[�O��Gh�U�!����o��ٝ�����~���+v7w�M$^����F/ ��0���ix������X蹡�|Vw��\|s�S�i	7�#{}��J��wl�c����wڭ_�U�1�n ���ѧ� ��<�@�MQ��X�����9q�/n􇼴��������ﺣ�$	6����"����x�r��C���7��t��'�G�[}87@�Ӄ�zGC7BT͵��-�ʎ�2j��+x��Vr;���;F,���)����no�7X�Z}��E���-���uA�\��ͻ��-���3e�	��{T�x����*�F\�4M�����t�����D��~؝��У�#�d�)n��ƖG�u�s���vQ:h;޸c,�{CGOw�����������W��i>�-lӗc�F��7T	�+k1��oZ�;�v��z�)$s5�� -jsi|�!�	��c�K~���&k��>�|��~���x}�3GTȗ�R<�Y>ĲL�]�s^|��ib�9�h���ʸ��5���T�[�/9�5��yQ����\�=UE�؋�%˩��[�w��\������ѿI���^�Wp��}�&�C���}�<���=t`��ʃ��8�d:{���FSY���M�rs����:Έ0n�M��!츩�M���A�y}�f�\/�|����dXV�������]�5����^��jfnnl��|����q\*���a��2Wr����+ޝem�t�w�WM�U�'g3�^Xq{�������r[�Y�һF��`f���<��2R� ��W�YM{��aa*p*�J~�{%B�������'g�r�%��z�ї���b^P� ��k5�[�H{��n�-o��'`y���0��� �}ݏt=úXq�����i^���"��m�wg��/�Y#Bm�شw��!/d�iwW�jGr�׈�c=�P�ɱ�~ .ݙl~xY���/V��jm��X�0��ҹ�2KkN��e�v5�t�C^�L�Y �ص=�O��/ �Nn����#�yb史�3ؽ�;����A�lǃ]�xt�U���������=�<�Ԟ����]���_���$�w<�}m��d�luX�h�D(E���7�<H�9�=�®��Qu'(]X��q��� ��Ѯ�\��H��fͥ���y	���96�k�a�&���wg�ˣ�'���Ԝ���>�;ϼx\����l�>��oj�{�P�wχ��|�;�o<}x�)�Ҍi?gx/�S{�"4#�|�~�Mf0������7=��5���.�NjҶt�=�^$M:"mF� ]>�P1��+�&�~��F/\���+uvM��:0*�ærV�ԅ�Q�A�崷l=�tjP��
l�6��L�WI��bZ�L��᛻���v�nM�Ia�n�~����.��݋RZ��e���9L��yO4�'���t::�K,����[ ^��y'w)�-Yg�E���k������l�=e���y�n]�yb�&	������*�U7�B��p��}���C�3�����I��� �u��R������ٳm�B���1j���-k� |��1�"�� V\����eh�\��q���M���L�x:^�F��>Pk�>�s��ݴ���=�����޲��/�b�ڠ���N��RLy؁Q�_wLQ�μ�<O��r)��y[ű��d�TA_V����}�/-�v�+ߏz{�g����^S�s���}���^?�>L;��r���*  ����y�����Q�Lz���䯼w�Jq4�UN����Zh�Z�_h��&����׾��.�x[��bL��=��[Mf8��,c�֮byP^�W^Zi�6y��h�x�䵴���b��.���qZ�iQ���hضlN���z�jӂ�,�Go��9�}GO�[y�+��S�(�{����Ԋ�y\�u����=�	��C�����������L؆�m���������c'�����4e^�G��ZEhs���:�N�-��0�F��֓���FMk�sr�a��x{"O�;�"��v���hO_�d�T;3�8w�NU����")˄W}j��?�7<�����	c�G�{V��TJ��x4Ec��֨�+n�����9/m��8�ِL��.q!C��^�G���^ɷ|2���/Mj�fK�
��2P�A��+8��d�s��c+����w��m0}�.�hk���i{K튣����8�"\�"��t{Ս� �r�=vz�,i#��(!zo�8���g쾻�9Azݯ@�4�مy0Np���z�����F�\:}��Sm�7�����ќg�OI����H�7�Y�}�v����>^#�xQ��2���1�ۚ�q^k����]Ϝ�\'�C;D�W��`��(���l��M�'����$q�b���i =�[�~^j4`�<��]�:u��ۆ+�z�9�C�]�\�I���u�J�Wxd�M���}B�^����m�z�>���[���ͤ�<�}�Z<�Cs�5�8z��k]��(^��8�����?N֯OE���i
�� ��� �=�_[l{x��)�_oukZ��5 Q^Z��ZW����n�Űw�&��몮(}��	�0e��5�����%��H����.��7DBo��凸#��Ъ��r͇��d�E�)ۤ�0�z=f�����{��@���c��J��O�9_m�\�*�,gf?g���	5k��^.<|�q�=����篆Q�3�_	N_��]Lj����q#���5�Z��xë���&+ɽCW\|�Xg��e��.w]�_�\��h��� ��$�l8Pk�JY���$
�4`Izzk�j�/���C�;�a��ד�ybҽʯE3V�[�r���e��~*����L�{�b�gug�9�A�Bi6Qׇ��͝�y�S�ga�w�����zO"��۸��Ȍwnǖ�{�C�܉]�V|��	N��	�UVx��a8o����H�浭��M�G #�a�r�GF��� ^a�-�����O�9�ϼ���\`���"����f�z�z]͆��t���p4qc��;����yx���s����n�X8+^�z�򜄙� 	Kx�y(?v엦�j�fD��Vum]/9�.z�p��^g�^ys}Ƀ�=����A��mvԓ��8���j�Q���V�t�3��>�5����9�o��s�͘s��(A��.��u�Y�M��È�t�u=&�c�����7�;3�މI�q�hmch�彛hWu#7^��T��\B�M�;}�a8�>�2G�_��G>�./_\J���;��o��gl�RN���*�`���'X���V��z����|���h����"u(��;�����1w�(�p_:H��=DI=%H=��t�����0��V��n����h�Q%�]��ac5�-���,m^ͻ�6��Q�d��Wn`{Z���^Ǵ�n�ȇV"��Ȝ�!��;r�+P����Os��[@�#��}���Ѽܛ�J�,�9x!^zᷨ���b�`����͔O	�i���A�Y�tٕ��}�6{�`4�4<׬�L��������r�6��gk���}���~x���g���w���xQݹ�Y�r1���u��L�3��X�Ӿ�J�H�Oa������{c�ԟ��c�!�C��]K�(2m�e:b0���ԡ�o�����GtIrG���yl�A��٨S �M�B�a�vg�WQ���i����nv��w�����e��� {&��.W�|v>�6{�=3��x/���K&�P@�ļ+��fl��׆z>�s˦�CA�����2ZW�6t��p��v*@���5�G���}���k�d�y>�[��n%�K���bھ��)
��2wwQ���f�ǚi�fq~���{����x{��<�����]��o�]���wu�t�[���}��o�\l�߇}�� X�Y`��$P�0`��r��3��)�X�.���BJ�A'A�t�H$��o�Vſ��cEx�uO������X��7:����Wb�q�k���]|�!0��׏�S�]�:.S�=H�#�Q��5}��1+�nZ:[=4.}Gg�<C��]n�>��/�[1��ݢ���zK���^�ݎ1��2�~zÖ�r�H����2�lV��t���vCÞ��~�TZH�-��mޝ��}��G�^�8,=�dJX��'N���#Ǿ��.w`RE���A/ydէ��F�^)N�C7���@��;�B��}Z���]����ي#W(HuVA7���Z�1hዶ��J!�Û���{��|YB���lڹz�@�W}��h����''l��-��!ga��Ɖ!V��m���N\��-���4��존�Nck�v�]Ի���*m� ��蒧%կ���Xb���^�o�S��e���۾�_,5�1DBLڧvIB���`���۝��M�-B�9j�m�[�5�D!t��3�ů�v�>|�V��Bv�
r�������|��]<M�G/�˪ᨩ"W ������s<ơ�f�״��������6�Ե79�}p��ux�X��MSe��RI�e>���1=�˯A���s� [�5x���f�������=���v�������`s.��ۊ����-���M��t�}O�&{P�v�����o)�Ci�8J�������@6�e���M1�Gb�0��X�l0��0�p�ƾ�aacM`��q�h� Ǆ5��k c0FD�`j&S����~C��M�#ɝ�;���
RgvD�w�ͻ�����'p���r,�.�"����s��)p뛁�1��r4rg6�K�Y��"�ܹ��v��.��r��Τ�It�� {�{����滹wa���軎���wi:]ۛ����븻�D��s9�t2t���"d=��&���nwp�vr��9��r�����9�ܹ%�ǝW�4�{��؇\ҹ�wivu�1D�3w:-t9h�CI�뮻������vu�u��wg]I��N].���N�~���Į�sw;�+�
�N�:1W#�u��~{�9�pn��]��qĊ���@"��g]�"��뻮E�y�8w7AS(\�@�����\�Nw?Z�w�߫�~v^p�L@]gwE[�T��5E����B�
�&�:�����ֈz#�|l�zQ"�_�>Ի|Y̹�B�o��(		�p����I�m���N�cͼƏ?ꝧ����R�~r;�����˯*zK�7�V!�b�o�t�~�����k�y+�S���>�s@Teu-����v��!j��ߩ׌�.}D[c��^8�'��5�m?^C1� J�?(Z�s��m3s�N�u��hqL���o�����Xid�Ľ����Ne!��R�]�Y[R�����k�;��V5�
@Jy攩�ㅵ��O�;��b�Y����6��ֿAv��J]��I���QG�{���4N��4v��I�}�a����p��MO��O�g�ꃦ�U��"���G��
s�:���;������?�����-z��ynS�{�r����^����~��=?g����'�;�kéU������VΙ�����`$K�1Z��D'�y=�?fy�~�?�����yZE�zt�孰l�����y{� r /�!m\:�/�C�{gz]ns�1.ڑe'�"��]�"͖�ݷҳ��m3�d旬J}�]JB[ɮ���m.��g2�tv����vl�HN{n������{u���:��z�����y��r��7`�$���S�U�R�ԼU�r�R��ߧkhOG����0o4�o��W+#�&�E]Uǖ��7�Y�V���T�!��%~��y�Iӻ�f����7t>khCr�B6��ŵ^�5���ew\)y�5�&�����oJ2�������I�x�=���=�����a���E΢���'a��pZ{�ަ*/W����S�_QCмX�ej��t;8�$��������΄��
�۵I������^>�{p>	�G����H�� ������l��nÛ����n�瞯S�y�}찉O=���z��A^�7��<1���;�����@S0�n�N,�{���y�������4�׶`��*�*����B���+_��c�z��m_�o��/�<I�_�����j���6��^�2���p��??w��I�?F���?�q���/y#��y�ڕ��90�/rQ�[3��W���,LmiZ��g=��n����Z�]w�(�B
�&�9�e<0��� ޫ:�J&b5K��R��ά�"�Y5g��=���b�%���^>�T,Ta$����5;��z�~,w���<�~~~��<�>�>���c"]ޘ|��^�Omz����3���lb��b����Ρ�3�y�^��u��y���T���x��	��b4U�k�m�{AcバT���]�Gk����a^�'{��k��B_�*�����+q�V�N&�������_n�n���T�U^��R>C��}����e�ʝ�^�_��-wp���-�w��ȑ�$�߯ӯ����=�W�w�*���c�t/t�1h��܋�����o��);f�k��˛#��	��dL���i�{�ǛW�Y��u�{�E�YB��"V��U{����2W���Pn� ���^��ç��~�,���A��P�����'�����t���o�%>��?96�E%esTEͧ�*�׽����i���5Y��{��-�r�D�n�Y��f���`{�����38`��Q˷��;;��S̨rJ�a�����]��w�`�+��b ���ޥ4&�Tfjnn�v��̏"/�Ryݛ����u\�f�J,��qwu#���"�:g�ɝ�u4V?ƶ�8;�:8p��ƒu8����Χx����_~��� ����[n�:7���s|��7���=�'���|[�&�4g�NU��9��x����\�3s/@[�<��C߷=)~>��~xǸ�x=@�F�g�6͍�rѺ�fٚR�w�͊;4t!�����+�9��{�3=<*�t�� Yqu���_��G�Ow��g��T�r��k�:��u	�}�T�==�5������ ��t7`�΀a�ys�on�T�-�Y)��ރ`�?�~�>�w����[�d4�T[�Z=�;���]�3gj����3�c��e)=�O'@K�Hw�-A����nn�/��Ի�X�JO�e�[n%�w'����Q
<}Z=�>���{�ן�����)�b�UAW6~�%l����7��6��w��S��+�]�U��_��J�П�OS���w�%��� }�<�g�}���=�%v�L�`�r[uE�����Pj��(}�f��G�k׀#*n�*$3��i�ސ���o���N}������P��x�k�?z(��~����z�I�0����v�~'��9q¸+�6�ޥ3r�����9���$���hj�b0q��g�׶$�0��ӵ�d��&{�{4s����K\��s�dF?��b��`ĨH��sQ;��w�@�Z�
���K%��vx(�W����ed������hh�Fgt��2�eu;�D��ၧrV��}P~����R������5{�kP��qwz=��M�����~=���y����=OG|��U��m����+�uylD�����ݚ�7�]��� ��ux��=�X��g���ڗ�A�1OE�mk�ULg���8\�"o�;�A;�x=C�0r�]�u�^q�y_�+K�P�� {��K���;�]�E��/+��d�	��gY���G'w�~@���|g)�~�ӗ����>�`g�5�(�g���ʝ���S]O7�U�o%�f#��]�
~��ƽ�������KvAA���6����f�{���-�)'_������>���ǇJ�m�a�a��Y��{��+��F���d�*��'teGg7�r<GNI��C2_;�f,2�xr�������x+0���Ԛ�(��I����ʱJm�^2��k��%��7ݫ��#�	Lt�H;����qא(��{��� ��e�����H�m��#�<�o�:'ثϫ}��q���w�nh�7�!�Dgso��SwrI��a�`���!�>��=a�><����s��~�������ͯ3�8y�K�[���z���Nme/nD'�y=�*����]���V��Z>|�oP�7�o�)Խ�^���Z�ϊ��О
����o�Rp��뤶z��ث�1M�L}��8���h����.��ln�B��sƐ%��1���� ׁ�*=E͸��F ����}�B�;Yjr���c���m�ejN�����e�=ߞ����,��������)��u���}Ai�ޤ�/W�DU=�����T�w�1�L�33�ᓿ>��8����(�r�o�����a������B��}o����}�Ɵ�x��`��70T�R:_Iw\uc��O �L�� K�U�x�Nԗ���`�����h���FN�����}�/zk�څ���׎Y��Z��/H^9Ӹ�����ҜY��� �'�x5��wz�HRo���E�w%���M9��rǬA�	+s�����n�n����+�����b����1ߧ�=흏E��i�S�.V����;�Q���z�5|�B�7R�������ow�j�[������x�X�;>�`�'��t�'���&��h�N��'�T�{�gzx�Μ|�F'Y�t��v�ᅏ�gj�	b��h�Zk��o7�9��_��z��y�xM��刊��Ox֥�F��-����S�[�*��c�~@~3�;���;�'��\MQ��!���8�j`|.��L.׈����6c�R�'���;뤫���y^��
�qw��!@}^^҄��aJ��,�@��+k��^��,��e�<�}畟��g�����!��V�qu=�n��N��W�=o -�.z/O>G͖;�/��>������G����5c������P ��~��.7fPecL��
k$����8%�����䭣6ա�7���3��.`��nxhl����<0�{�/?W��͚�dV=>�jZ*Wr\$�E��5m��\��aY���ص��m5*��Y�l��p^���m-p�칺{��L�J����1��"�~�L���5)� [�]T�͐~{ӨL��]������ތX�ɵsf��c@�h�Ef�V��)�ex������xz�Y�fW��s��=���=��zh�y�u����wz�Y
��Z����"y�/�]���~�x�ѱC�\�VWy~"����T;�׽�Oxo{́	�n�Ҹ$�뷼�'7ߋ��;^8A�q�v�;j�\���oi�'��`�K��8�+���W��1���W��{�^�{^���/{<A������d�\1�7���P>t=S=S�sҺ��Pr'������=�����cS���l#���Ym�WV��*�e�g�c��B���K����K>�ý����Ukx�{�y�eMi���LBH��z]`�p�q{����;����Z�n�9�=���&�~�6'��.}Un���W���)�k�A�`��e���'��N��i�5!=1�˼@e��|����4�s���=�]𳏒GےM��%���!��������|wy���8���/��(I�������ₘ�1cl�����	q�̨�m~�]Ԧ�cy��ķu����ud���0�4�"�Z�br��NIf �X�E^�p<=4OI�{.������ۯ=�8FzŰ�b�L�4��UWGU�cu[Ǩ�6WyJ��j���Ԥy��g"�c���>=�}���������OHo��1O�
�I�2;�PWh^�"S���O��x]y�W���3ނ�0��������0x�lyx�`FHOz��Z���b(j�.���V֧'�`Z�td�T�]冁��Z�^a���	��T1~Y}꛿����؁�)��>%�e�y�	����RJ�/G]^��k���4=��d�uf�/Q�����T�]����K�&soD��eOV���;���?޹\7���u>��5/���k�����8�cΌ�g�A�z
=��y:����=�}����|��S=4�5Fs/m�d1�6k�� �h�������̚3�M���'5E�c>+�JU/Z@���n,���[	����
��y_��ױv0���1K�W4�w0@�/�x�������5��e��1�z0����6MEQ��2�6 q���l�6�Z��.��d�EM>B�,v��5��~�%�.'_n�u7��j(����\w���m"�A"o�;:�C�v@���x�U
~Ė=�!�������^;��ޣ߷%x:��6I���pupd���n�5W��z�==ֹ���K6��y��S&���Y�Z�^>����/��-�$״��c���k���O�fU�g��feܞS�h^��QBO0`�gG���3׬O<�9���1�{n�+C=c��^j�J3gͯ���W]��=^]Z�A�N1����=3���swͺ��r�U�0_[��M�;W^��J��Cu�\�5���=����OH7�+۝�7�X'�I����W����:w��Nn~���h�PLx~��w�!;�Ǒ��O9�^}�D�C�4���ꏪܕt�^R�M�FW�X�z%{a�ҙ�yL��nK��y�W���m��G`���ݮ�G>���{�w��������^�W����{G��T�o\]<')S�ĳ�X�H��׶�lE�����W��Vv�U{�f>(37^��)�(Vzc���ފ}�dN]�!���v�fv"����1zR3��电�a�
}���������FL�L״K#·5@Ģ���bON�N����2MG{��?����1�JK�~�\�#1 Ǹwk�mT{�z4yC�9a쀅<iG�lt{Ӓ������� ��~x���axn�ňԛ�c6S�����q��w�d��]{�-\�|7�������X����^���������=y��}fr^�{:���	q"�<ۻ��B����z�K�i���\^�{��vz穧Cev�	^�}�nW���s}�,����,�1����!�=��?]���q-`d�_��K��)��g��y�uъG���u�v{61~j���[Y�t�j�LQ�|M���mS�.Λ���&;�����_i�K�s���F�\4��$��+�l8=�.f��h��>ۃ����xf�V�����R�>��wj�Ռ��d��*G�����n�y^~W�|�{�[M� x��ތsS�� �q>y��O���r��qu~�7����1h�/r�Wz�Se;���Qʺخ������uo&}��
3&vh�Z@�z$�G_3b�'�<�i����Þ�VKڗ��xjގ��d��5+��Iӭٱ�K�	x�t�m���wf=1��? ������|K��^��dN!��#�˫�E��j"�N�n�/�t�
�ȧ���9n����K���[�~�~�j��P��TEV�~��\�5"��ȢqG{w��6��C��y6<sL���us�)�|{��i�U�^��ŉ۾�Wr���g�p2�����qw[e��E�R�D�+�3F9cf���"ח�1�P,��Z�ߌҨT �]��
�٦n����'C5�N��D�:T������vh��S��z곻�p��{w�{<�I����s{v��u>���
/7Ot�`�j�۔N��n�>ug��iPY���V���#�!۞�4C������~|+��,�jD�c�ľ�U�B[r�(:�e���F��7��Ki�-7�q.{�0c�;ilI�U�n]f�z"��J�l����̳~��~�Y��焤�:�<hw�%w���U��Ďw+�w*~�oPm�6Й����pu���+�d��QT$��K��
���n���U�DT��i��}�r�m�@ϕ7y�>��r#���O�^�� �k�ڝ,ڐ����P��6vn�����udWc�}�^{@>��[��0�l��^?%��}ft�I��ӱ�@nP~җ��<Yg����.�1D��=�T��Q+�n�4�ԁ�E�y�Q8e�ݣ}�i��'�Q�����1�ӷ4S�c��]�羘=�<�]��v�j�V�yht���!�=���M��x�Iט�x+0���9�MEh��;�����������}�q�����W;���n�B9�ۦ"�uEr�\�����s�G.�p��v�t\�ۻ�;����]w�]��N�w]�d��IΜ��� ��Di��wL@�H��t�)	)(M�wwr�.��zӮW+���\ۈNn�q�"S	.깑�����wI�wB7w���(�Cs�D]�6C�.3	E-��rH����!(����S��]����.�	�{r���w�ޢs^^]�����.����`owCw�k��u���^���w:�����s�u{���]ۤ]��u�p{���t�z�e$�rn�.�\�;�_�޼�㻸�l:�]�;��ݻ��{�ݻ�wa9״�����vm�^���2������zN���v�=��[��D�7wwN�nnÎ�݈�w\��E��KÇ���	���^�B9ă=ݺ�e���<�=�wnfȫ�~{{��u�z萅���@�`"�f� ��8�j���~�^˔u���mnR�.���zg�f0F��U{�W��$|���Ś�|x���Q�롃������+�����ۻ��9o��bts�h9�f�0R��Cy����	��A�JȤ�[�����Hdr��sIw쬁��D֘{d�����gul�2�;} ��Pɇ6���J��NJ�9��G��Ϳ�.�HT�����ʕA��ǟ	�zj\�3u���*��q�`9����sFK�o�w/2���6��D�<Վ �@�[E�E��>����[/>��%6��t�����J�q1��6�ʬ_�{����u���іx+M	4J��U�u$;��N[��RM�-Y�]�Vg��:ۅ$�q\�	d�-i)�V��kw�{l�t� �)ơN9>�jof�\h�z�l���R��p�&Ԓ�:"S��b%9�.�LJ2���u�5>Eê��E�N�~�4ff��|�|[�S4��Y���Xa�-�aqJq�6���x�ZEr�ZÚ�E����&�]N$C��'KX�m/>/
�!#���Ƶke�<�i�[�ZK���='�Zs�����T��#b�գ�%�;{]�L"B2��#9c����n®��gE�ήҷ������� ��żؠ_��0�jj�3w��5�~��c������c�j�����G��d��c���׻L�`�_��{{�
;(Бl:�s3��ѓy��N�?bs6kb�����Cvv�${w�w��$=fuj{�y\g�b���)��k�ށ���ȩ�V7>O~��1Ơ�C1`��hg�0ϑn~^WFŗ�0%�����J.�]�V޾Mu�b/�_Z�GS�
2+�>7R͕�E�>
������9v<tP��pbWםn[�9�a0�cʎv/=c�hnAq�l|L�8ż���c߾H�f��u�R�yf��	0��8Ȏ�(�� ��0VU����)�q�'���4u�Zf��B̙�0�xr�rY�`�,��X��;#Y-���s�MUZv*��GC�q�d�1%�� ����?��VƸrW����{�c��\��-x������+5ټwR|m0n+=��3.Od���E�2�u�ijh�X^J��	B����
`��d^�5s���Z�%��̦���v#�qV��!���椏��5�� �l�*�����2j�qtj�0�����]�ʼ��&��r�$�Ͱ.��H�\8��lod[9Z���7��W����^X�q�M�����i��/*��(�ƻ"�X�FB��A�=�N��U
Jd����T[W0�u>JJ����h������l޽a�8{:���u\�$�����W������f��X@N����V�Ve��K�"����Ӭ����5;�y2��`Y�G|�CUx,}�����Q�vk���ou{*���[�m���EZ<�m��U~��g�Ǭ����p����G��ҷ���f�g����o�ŨtBd�1�ߒT-XUE8���-��O=/ye^<��d�0�,��7�q���Ύ�!��heB�Y�k��eJc@Ą�?��I�,zj�r�Fq�b�8�Ce�W���+�eٲ�]xhɖo �kH�!9���a�	eeK�����S���k������qyZ�ؗY�0�G2�x�f�ٹ���Yp#����a�Gofq�h`�s-H��	���(aC�i0��s�Z�D�{y����7��(�e�� �[���s7�&
�V���Vetq7{�HcU�qI�*�KG����U-t��R�`�f��2A�_u�Gb�j�Σ�/=�Sj�X	��9��r�jéX㭗J�)�錨%����dr��T���Wbr]���ba���78��9��e��Xk�*�6t�=�iY�@���C���7�M�<�������0��!���rpi��y�:� b�Y'Do/T1ղ��b��GK���#bUf_\��-tcu�3������%��dO!U�ZK.4�B�zn���piT�­����x��y��{��v��w���>���G5R�ݼ�=�����8UZׄ{�ǝ{�=��_?�>�yz�]�G'f;z8�T���=$�;�5��'��Q���~�%Z
?n�6I����.��+��J#0SK�^�p����ϝ�s9���o��(q�P.�Pdq&����1<��d3P�{�F�S{{wH��G�7^�s�ME���b��Y�Pyj!�VHB���曌�M^鋇\���y��[Т���fg5ڍ`Ȱ!��z��u5շ�R�cQ�!s��A�yfP�T�p��M�1��,R
B�:,����w�CacMAiD,,�m黦�����M�Ȁ�P��Z����\�n�����������Q�)��e�!�T��C�L_�!^��	���9�7���M����e��®�G�����IP&U<сf�Ӱ�Md�a�e���9C���ho�1,q�u�MV&]R"� ܼ�̬u�^%�u��L[�Tx�`���(�\`Y�AƦjt��a�߳�)"��'���Q9�J��U�.�,�'L9L"�{�)��P�@�S�f������W��Cbi�_Ͷ��>n��f�Vz�ޕ!2�7B���*ʞ��j-?5� 4�z��k�\8��Y����,'6~A�z��Za�U;4�X�6��a9BV���إC��oN��S��������&�^�Agbr&}7akצB���ś���l��~;m�`퐫�2)�чC;/e�P�S�gC��1%vDW�n!���5�Q�܌��uwy�>�^������'��_�%q���f*j�[ۘM��7qʗO]��B�%w�7(el��s�,�$��! s,:=p�_�N�6����N��S��<�4�����{��d	�O����m�ló[z �,8��(pY�.�}f�n[X*��n����T�+���kj���vv��[Zc
�-���fy��ܻ6Ʃ[_W�1/��>�_�F�cP:mƕ�s��t�U���YQ��p�̢�a�IC�@����DS��mq��^�u�7+&��~���y�����p�"jW=ʀ3],�A��6���9w̇���q�ğY.�7�b�3�$ۧ+:qU9�M�wDAii����9����ٸe�t�,:��#;{�6G.��������ۍY˩Qp;K��N�b�-gg�˙��T����ׅ��5yty'f�;(2o'm,�Yd=����R�d�]���,%����f��cԕ�� �(	i�d)^|:"�wO�C�Z ��5	;>��6j�k�W�O-K�y5�WN�<�o���x/V��'�K�&k̓����r�.�]���\�Vw��]v�B2���bN+�;v����ϯ��I�� K. �+�^�W�?J���Qs�|�U���GGr*2�@wp;����,�G-��{{��"kՕ-vrȹwW2����$���7\Ww߀�Xθ�C�'��s ��(�����r��sP�fd[�K��'�MqX�V������%�;�H2���H̛v7F_B!p�����>�y�s�ᜰ$g�PΥo]-��>)��t�bQ���=s�^|��M���l�.��y�ͼ~�>C�����2��A�2��̧~�P�j�> b)9Y�>��K�.��,���y���`��V�Y�eD��rC�������kZ���-ky��͈��S�8���gu��'ɍ�dTA���2� �^G7�;�T7� 0��A������B�S����מ�[�Жׁ'��![�WxN8��wNa�q�F?��%�� XPC`w�����ɡE�zjj�.iXV޾����!��jK����6�~�t$�R-I,���1���467��ȫn��n���`��+���"��*9M]|��Χa���1�Υ0�_Y[�����}P4{M�>|��c�L�����m�!�f����{B��p�5Y�����R ~�(����0VSH:S�d�)�7T�xͨƄ�U���2f/�G��)���[�kN���Bۻo .�d�4]���{fs�6J���b�30�t�8]:`qy+`[�%&V%cRu�Ӎ�����f[���z&�����\��7|�p��=�s��h!'���kG��<+Q��U��=[��aۗ&sHt��M[}_�����j�F�;�K�m�	y:E�d,���[�Z����Q 3�OQ���\[���:�v��y��U�t�;bl];��_����}�y{��b!*���}�8�����-�=y���%�����D{��Ҧ�3��/���}�,��RlZ���;o5�����YАp��d�E>���Ln��!,x����*�� M�5L�`|][ٽ��g7T���4h%cj+y�O��a����WV���{j
V�4zPf �,��/#6��)~��59V#��PFs��� vE�4�u�}12׾QI��"QUE�2ڋ`&�OLt�3���W]G.iv#�ؠ�k{��k�/	;W�e����L[��$��饟!����YIn33��%��X��ϒ��oL�K+�M�8k�=��򵡺/�����.�4ҤɽORK�rlv5U-&��Vp���.+�jNnԍ8�MRS�xdAƘr�OH �a�,��:���T�B9���GW,�g7����I��)��=ZP�~�.. �x� �c��K���v!�\�.�n�Y��Z�0h��<X��W[���M]
W��
�Y��C֮Qy�Z��N�p�f�&��5������ڣ#|$�ߚu���;�`�h�>=�B͹��.��,*�O1��XHOtZ� �^"s;WK���iE(�c�2�S14�2�l�]����T�UVIkV�fxx��'7��	�,ku���Tre��z��3�=�Hi-j��و��,����xW�}�%Z�s���e�G��z��q����j���w��SeN�l��6�7�<=��;N)�N�������>`鱧�U=#�k8е~u+u��Z�⠗��PK�^Q�8��Y�\���ݹ���fA9�0���,�@�5;.�s����)P6t�8
���nZ�F�ʮ��Xv��򖊽�kd@���wPD�@�<�<R�8��=�����ni�G��{�ϬD����{- n�l� f���hBX�D���;I����ڈk7�4ZW<�\�W�����+ch�vyC�2	^J�3����'��`A�����sa�u?-C;��em�5e'���{kͅ�^͂��Q�@����y^i��t����lI/�O�	�U�%�Xj�u�!@��)��3�M5�M����,�t�<���r�>o5;v�����}�8y�O���1P�Cs�m��������e�l����t)��)	�z�U�om9��Žhn=��2���wQ�)��e�-���}�C�<�{E��˪������&.�\��%}/���{�Xkw>�	���7Eq�4JpGQ-�Pr�� /`ٍ���w�A��E*ra��~ؼ���������4��׻FX��� ��C�E�=��5��w|��*�Yn�Il-�"�ܶ�F�=��L�y}����{�{=���%w͌jT���_C�g"TGo�1�4.3���O�ꍜ�]}#�O���ٷw��
�f� ��#^��e'E�Hs�1�Q��W8��a=y���ݫ����]�=�W|�1�+���5�H�B�'yb��ʥY�Cl����5�N�R�ֽ���4�+�;Z�8*n���C�=!1�0�
7��������='��
�ƀ]&���Ի�6$d���"ɷ��9�Ƹ5���&Z׋��+l��4���冴>�*��0�j;���Ef�5��	Veͯr�����BL�Ϫ�ze/g�SVm�DpX�]�/"Y�i������{�o��+]��A){���l%��x��g�z�LL(�=0�����A�F@�4�k<Ɖk��a����������2�;]K#s ���yO��G1ʆbA��d�����L,�����rx�i=gv�k�r:���}�pcϠ�lx�ʑ��ϸ64d�[_؜�8㶬w!�MWLZ��-�ou�'i� C�8��9���Ih9�3k)z� ��ꆐ_E��ez2|�tm����t�[v#pS�����)k?�2��<'�����O���mf���è%to/H�cj{}�"�a6c4�s���܊�j^W��9G��-���^�=�:�\#hm���ǹ�Z>^�䦓�w@���S�kʎ�!�����������˚������:�t�.�n��֊�����{�U�}D>�O��q��s�y��,`�h�nx ������JŽ�a��:���E<5��<X���'M^T��^Xjmޚ ��loX��Ӂ�-�+T3��V���5�'h=ٶ�53��?$��^i2|�s���>��v�֌�;W�"$�f�����%7X]  ɖ(����XP=�@[ռ��|�
N��g{���ꞋUGtvF��:8d!Y&���N+ܢY������f9�q�ɦƆ<j�Ƌ�jA�<�K�mQ�Y�4Z��N͔%�05|�i_A/�)�|1���,x�I���K�߿{���]ꏰ}c�)΢m��b/�W�C�4���f����m�LãW3�I.�E'+�5����������M��#5���l)�-N���~2�0p^^:!6Н���6�^�v�0���5W�+��z�x����j�{��y��~����q���
�k�����i۰����2Mn�h�@�;A�����|19��߽��>�W7��0~�=�Hk�Ka�,8Q�ap�q��:-�a$ʾ��r7Z�`��� ����B~k�d���گL��6VŻ�l�0b�7�}>�g������}��o�����>1��d���?r���̲ ޺�H��GZ�[�g���8J�}�ť��-�~��G�FQ69h'������sq��Bp�&zf�Z�}V.�n������M��}�hsˎ��؀����j�]���oz�_���T
�o���݁N�xz�ݞ{r�w��=ԍ�7��EE��7�!�,��}��>K�୫�O��
��(���S��Q�2�u��ۦ�/�l#�C^W7������o��)�z�N��9����Y�̄5q��N�o���z�y٪_x�O����~���U
0�i���r�Ξ�yo����o�t�
�HF�٠7(��V�3\��un�+X|'T��d�u�L��(z��f�ӷ�W��+���s�]ԓ*u�$��-�h�M��燥�E��4��)�D����]�W����f,��V�Z=�z�Z1LS
<٣���n �uS�+�{Md9BR��7��M]i�8c=�V���krn��Ѿ�{�M��,w�v!qƞ;�V�q���w��{f���^�>w��,栒{�z�9cܗ�Jl|u�7�	3���լ��>ʷ<���L�ސy�����<�?�ޚ&� ���&���a�.y`�~�	�y��*�Z*'ݓ_]hM���qH-��;�+�޵��ٹ ���3�g����S�#]���������{n�s��:h\QkU)������亏fů,���_=�Z��/�K��	�yw��s�z��gy�t��Ҋ
˳�ou��kû�o�(|A���y�n�&�W���ͅM-b�D&�V�`�`M^X�`����+��w.���B���榶|n������܍`����v�L��Z<��޼���ݸ�:ʎ��s���pw���YQ˧�ؑ>��a���W������Хb��~�E�5gN����{�qy���`�7{�hɛMsE^���yfs2w�z�C�]�pF��ޗ{}�ޙ�Ң�ނ��ᶣ�q�K2Z�w^KO,�#.�׳�c��'��&k.�D�����VD�����2;���/k��w%~��R>В���GP�]z���qȱf*o5���m{u�>~����c��& ��ݮ���K�����J�x�/���n�� �W�
���=�|����ߦ��Qs,��y$��#���w�i�*{�t�����N�:�!.c�Ӽ�+fb����n\T�f�W�.zS�!�����󥿇������"��}9�d�`�7gc�W:��s���2���#8>�ﵒ�^�ŃLݘ�_v�V_��N��Z�W����Ý7}����]�ݺe5�*�Վ��C�ԩ�����g\'�_g5�K����M+���].�\�E�s��ֻh�7��t6G��{+�˖��u�����x��b7��F���.��P��oR��ᄡU����p	:��/��o��{����9��X K�(�o=��ݸ�^�#��r�u�绨�E���{�=t{7%�ģ'wJ��{<��]���p1������ߎ	�u�0��LwnI��]Ӻ$ߋ������%��$~wf�
&N�!2&�$O�\vSR�����v�0�h��w�Wwp�7w"g��F��oy݄��IM��`�9]�`Gup�I�1H'�t0$ ���Dd�d�0D"\�BRi	��@r�u�PRa'�q�		17���4���̙) ��\�!��;�wWC	d��!H��((FP�"f��P�ݢ6��3&m��0�g.�J���$I	���\���Mdw\0�'����~o�w��������{y��!P����*bo&�|���/��xK�m��� ��yR��R���ݡ��w��;H�XB~��D�^�z�!��˞#.�<���g�
)�|��;�`��%�=� 8Ϸ/�j�^��1#����Y�0��u��9�sow��n�#;�rTcG�܃��U����r���3��֣����k�⮯�CL:l/�Ϻ;M��I8!���؀*(��n�)��Qm�ي������n� ��ǁ�-C���]Gd=����4��nu�q�.�,����N�mN�Ue��MӪ��၅䮴3����쾭�����NV�yS�����õX�D�{����LʚuQ�k	N2@f�y4��A[B�A+�5pT�VȻ=��ʺ������v���bPJ+Z��A����Hb�c>�Ͳ��7�d������>�k�~�g;���Q�;A��ǞX5�
�y���'泰�zH;lod7��VI���(�l����Ym�q�c����(
lD󌇂�1�vL.z�-{��XZ�R�QaLƫ^_{�o�\������+]�s�W�Y���0�k�xIڽ{,�/�1nwL��	��9�eąps�f8�Qճ���'�"����僌�,�=7�q�S8G�l���ٴ3��r�G����MD�.��w���=s��ov2�[~7��g�~�w�˛�*�4���i�+��E=~�7w�����6����8,�g��Tk �O����u�f�o��T�ۗ�c���V�6��^��}*��]��<����x�'�N䇽=�k0*��U_��Rp�f３S�_��K��sȢ�W�GM�f�xa��o�B1����hҍoJ.o
SYV�"{ݨc�.�Z�I���m�tY�2�xԞΓ��X��,��GQ��1��O:&���չ}T�6S�7�ߥ/e��i0�+���=/�^F��l{��0~(�d2��[S�OaS̷d�Y�y��Vܘ=��@L��y��Mгnd㋱�����W<�lR�a>	��t����j�!�������U�y�`Ʃ�*n���k'�i��5�f������.��S���|�o���uݪ�&�1����S.�؞jOa��08�ft69�d�ht��-��,9�
T����a�k}	vq������}��,���n!:u�1�Ac�P����J��[����`�(����7S����^�.�a۱��fa��c�%������XU���*+te9����y�k�񂌹L�z]�[�'Mz�!�%���HX"�t�&�X�����y+dѼn����z�3��ж�*�E�ME��X���߅�J����	��d�(My��]6����j��t��qv�ݜ������<ԎjZ=���iBv�$S5�Dk �Ձ`9����ť-��_r��v�X\e�X��2'X�u�Oy�NvdXf��t+o�ؽ�������Ʃ����y�є-���e��L;L����+��u���W�{�峊w�IWg���@�g��"Ô�D[��x�ƞ��R�ԹH\�]J�D���2-���gv�������#�p��僉u�Z�+B�qAֳ��T�ݵR���%6����f�Zm}��CD��珌���o��逄�/��C��Fȋ`i�+j�{82���Z�B.g�����	��J�w7�Zn��-D�pGQ-�ry=�#'6<#:b�\�Ngu8Bú��F�#L�N�Ĳ.�
�ceL(خq^w0_[X���-=��>�����&�,_3.	[ǩP�*�$J�)ދ�t�{�J.�s�7���+�z�m?fz�9�w�k��	������@���Za�ꞐXװ�
7��������,h���<��L��mJ�uK5�r��k`�=ځ��0<��#�zu�ǫ���QLn#�/��]�P�`}ww�uacf��ܯV�\�@�xd����pX�]�yz�8��;_(-,�O���6��-"u���o-`��:���/~��஥�ht[�!�<`���f��-����d�M�ڞ�ʟ[An�q�M�T��St�Yf��n�mJ-��鬱+�m3�,^ʐEO��e���g��eXǜ�f�}`�I�����ȭ�ƿZ͖��&��G	�+��7��V]iDl~F�n�`�|����~��~��Z��o�m��f꭪à��ί�����1��
���GS��N=�g��ܳ1a�������ϰ\���s��C⹴�u_!�~E�����n[�q�NKj��1��vP���:"����,���Q�&�s��#�A�h�ka�i���	�!�V�X8�s#6�����S8CQ�뽈,����!���s5f�V)����ñ\3����e���cl^@�z��f��,:�,�K;6��gmor�{D��Θ��S=�2PP�ϣ�1��<�w�<�ˣ'�z�����$E#Lڀ�<זN0-E��3f��M<,�	T�Riu+ς����J�
��0k:70%Q^��	M��PdԱM'���XP=�m4�^��� �d�%*Ls2�1Kfmn�Xm��е������!�D�/i*�3+�I��G[�WcŪ�t�j��%�5����s����S�O���a��'t�ğ�q�JS��%��&�޹�Hܢ�l�>��u�A�.s��f��K6���eXe�)�)�N�T�ሤ�W��S*x�DNnN��nA��85���w���}�z��Q��4���"N�i�;������ksO=�j��ygk	�C���Ƶ����le_�`D��}�GJT�`P�V�;�Ȏ�2{)[��1��� 3�'�V�529I�w][kzK�Zz�(ͼ��g(p��>����xxx{�^���f\�7>2Mq�Tw�	�����ؗ^������~2�=Â� �\�o��c�F��E�=�I�����Q��˦lv̛�֔{_?O �����]�0��a��XŴa,��75Q��=�O�o���S���3���U�P�#X��*;�������*b�p�1���Ƴ�[��e+��ު-�X�7B����ʂiJ�r}m�_d��?�f�0K5�`��cI̶p��]]f�/�6w���E���|Gk9P�~�0�c��.�Vߤ�s8/���[<�;��p�+�R��	�P�`��W��跬�ߔ�H�ps+b}��\�e4���w��U(x�ݓW�s���	8��A!)���ZZ���쇷��y �q�Y!�H�%�Z�ʃ՝�i��.��	��tE׊�1Elz�9(p!2Ĭb�q��|zk�9�8�N�D�f��:����v����<�@%8�5 ��i�ƴ��6�h�D��{��n��4�H�C���D��F,������&�ӷ�8�-���91j+$����=ٶU�l��sӹ�z�,�}�|+�c�T��N9Z.!�uxd[�ݹ�.Pϙ�R�'%����&��.�ዥ����� ����<���
�a1]�Pg��qS�)6̏�W�Y�a!Eb���`le�r��q	���vU㙜0p!<x�Y��rp��yO��߿���~?�kj��֢�&��@����G��[z9�G'�|Ǧ�5�8��`ނ�Xa�C�]Z�@�8��~�^��}��z6�~�q�!��R��|,�q��c"e�c�Ru~Z�R�p�T�MR�MW��U�+�`[�\�4t)G"U1^p���#,��;`��n��LZ�D&I���7���!���}x���y�{�P�~UE8�c�)K.��L�>!ƃM>G��R�_�λ�_�B�X�^ZO�{{N}���]J�,�x	��%�Íb:p�|�L� �pTŴqʺh��fĮ����������,�v�5)<߇)�E�(c8x\\^��0	Ư,PA�J�O��>:"|-z��:��ϫq���~yN�ԉ$a�¨Y��^�r��PX�-�L9�,�Wvs���U�&���|�3��p� �S��$9��y�F�ف;$��c��­t��R�`�WL#)u�c7{2��x!��[d�D	�OH���q�j�J�~eҵ��[�QqFrW7�66�gE�n{W�G�$>4i�N� ��p���\vۖ�z�_�_�ˍ��a�0�-��˻+#�{Y�*�WSslwL�o\ɝ��͍복z���i/{�J8/_o�:VËP�w'��r��"���Λ�~.D䆺4Fm��ȷ'��H������[LM�ٽ�����cۗ�sZe��z����&X|����<<<���<77N�M�K3����b���v��Z���ۈN���uƸrP5�asRg"#>��>�Wo��%�1�X�	7/xWTkҴ���-�sRGƶ�����z@��mû�]:au�7���!�]0�W8˷��u�Y44�$=��p1ۮ�悖���Sj�~&Pgu��w��N]�f�����5Kp�1&����̈́��tŸ���"k�W)E@�9L@�Y���>ccy:��uH�P�
�)}܄x*��2�\��v���B���]����2D��[r�.o3���� ���
YB=e��<��!�t8�v�������沺����v�Y��kꪳ��sm�RX�R{U�B�q��z�IL��e�T��!���w��r1�2���$���غu��	��)͂�0L���5l��k�<'�[�	<s:�M�Hn�5S���Gef��x�2��D�eW�T�N��K"z��m��c怭F�	q�a���t�[o��K.�>	�OSЃ��J�U��^S�ʥQ��cAoT7g�Ч�����q�y����[Fݭ죸mv"��\�,1�m�w'�]y����g��tyߞj {�!J�+��[�������ە�lHZ����檐j�+u��W�;j�/��vl�|�X�
{�����W�7\��w��e�����֖������xxy�{��f���0 xY����g.��p������C���n�'qUeWCը���	����,W��M.�X֕�����B���0^�`-�,[�ӳE�����WJ�UI��U�k]�˛Ѭ9l�a3`R�����׋�e�B0�1yx��r��5^=����S���*3+]���΀)�n.���t˗�~�f��8��`��B�/����{�mUeG5n
d^�E1�Rcl����O��G6���6��!�k��=ƪsM��!��ofD�|�|
���~5fC�y6��*����_�1�I\Ze1^:X��i�MM����L�
���L]-}�NJ�u���bL�{���K=ƃ����'H?����S���Y�}9���a���'�9(G Rv+֏A���#M�`>���8*_&�.�I��nu����U����Y^�]����qC�_Q�����S=�g����P���\���y����덓���=��㬳��n���*Y8��v�Ǫ�xǅ��1��,��>oK�^�O9��;\N�ʠ�{[�b������0�:*Z�y��i�J�'u3Yg洦�6��_��@�>{:���G��]5��']pZuM쟞ؖ�<S�sLy�)�<ߐ�f�s����8�oVV9���^rW��%��~������Z��U�Z�6ՙ�����ox 7��U�r{S����=+�G�TX%{Q^��D��P�&+�{�{a�bL3�ZlI�v��W.*%��K>���h���D�DKjd"o�BJ�nwA8�r�d^�SL�ʍ&�~����1E�A.�5��]�Qۚ�b��(8�)�>j�+�t�CDb�;�?�CV���_N�~�|�s3�6��a�g��R��=Mj�I�o�/93K��j��Y��2���I>��}����D뾭���7l��
����1�K��0V�G�Ȅ�S�����ڋ�^�A)l�y-UwL���o'd+a2��r�O�4\�/9��
f�D�^���q6���އ@��(�s��_t�ev��b�%[O:���1�&��"�mH�0�?s�|wo7iD�b�-��C1�".�����օ��͎vz��$Ȧ4 ���e(-���8���>���l��wf�����2�Im�U�=qd�ǜ7h2�P=��E����Ḭ��y��G�U�Q��V�y�d��B�e����z�<�������6�q�sk8Fڴ�{G�����I8!�
<���ޛ���������v��<� }�q��V_�{����yck�{���H^�H�=7ܚ��*�j|�Yy~���g�����Q"��	�D λ�c�.�[���6�=�T��FV�':���b\9�V�W���"�?U����O���=��x����I��O��6��5mj������V���c1mo25�:߉�[���	
b���Yz�-b�Q��ۋn��2aMMT.w��gD�x���~�� �s~:ڎ"+l)ӌ���[�%p!4�"a'\�Ò���ɹ��WѻjZ��&}��L�CL�v���"f�8װ���n ����:R�%T.���7V�v�ˍ��sȽ�j�նlVӰ[�rb�\�Q�g��6ʱ	c�Y6t�jh�x�ͧ9W�Oh��"�ُ,zk(%��m�zO�`���Ɗ����?^�>�*�U��پz0�6��(3����E"�����ɫ&=�A���N�],�U:�Pz�a�f���9�~����b�g��4�xLS����Z��r��M眱'�[:���a���n�iٛYȶ�@dD�┊DU�����к1��A�" �Dl��kn53�5����ҙ�l&�uL���_<�/^+�b:oLjJ`�� �
����U���&sbcY��f�ڕ���e�1VU;H�O�_9Cv��4�������1�q��7�����x��=��o�����x��4^Aי.iQa\L�S�U��)>�"��Љ�Q�wLk/<�!�)�+>�u�֪����`���:X1�ǯ����k���ac^�}�f�{V��<��e�q��e�j��{��vy��jUK�{{��Y��(A9�챟���f-�����Ŭ���Q�G��Wt_�=.ڳh>��%F��t#��(�V�9\]�!��Q�<�-n����O����t}�_Dzn�vv�x�
������������K�Di���$^�EP�����E�I��"[�"z�L�5���<�ڝw
��-�������N��}�����8+��Լ���(��j�"$�ˎ�0d�1�2i9q<���x����v˖J��������2����6�k�NkfއOM��k�^"�N�m�t�Nݥ��$�w��=��<��c���oS�=��vМ���m��5#�e��K�8�i���Y"��$�%�G��ϒ��{�[�4��֎�=�o�������Κ�=�W�ْ��ꣲq"�˦�*A�(��L������%��k�R��B�c3��ׇygn�Jپs\�ާ�)x�Bⅷ 㻟�-���f�o=��[0,������݋;=�S!ۀ$��(����Ʒd��;=�_V,�8���P9[?��Z��x��u���g����Wˇ�5J;���b�x���ƍhu��e��Y��F��w�-��\S��+�����%��r��F��ٿvs�k׏e%�\�?�u�q���t���n����kk&�o{��!����W{Gy]6��o�H����/�Y�oys���k]λ<�c֯���7�5�^��X�a�ZQ���_U�������I�����Ni�����E�{��[�N�y{F�T�g����;F�T�%�o��#|��z�D�?U��k��Z����\}�]��Q�\X�N���jw���4�������F`%֏:�N[�z�P���K����Mka���A�e�jd��D��a]��~���P��G�6${�����w�`�]>F=p�Os�8
���}{�2�L�M���v��;&�*\���fd��#��|�:�ۂ��➻�f0K�ߒ��<Yz�,��]�����
yop
Um�q��.Bh��~urwu���X���J��s�qL���L妀@	,�圮��!Í���ۋ�gˇ�����#X����1E�Ay7؋f����m{f��/ZT�����{��kA��2�+++�.����1�`��Y���G�dͣ{X��#����������9��=}�.]��L��V��fQ�(�.���T[��/\�qB����^=��]ս��2�����=}���O�>��������E�sc�*c��A޳�\8�����^�ҷ.)=w��G�q�_e�KG]��,�ɛ�����*���h�
��}���� ���L�d4����f4b��Nn�$�H�e'wi�/w#aH�!�a��W<`�"yؐ1��bI�d��(X��&��&\� �%*E�{�$�92�� M��Q�f����4��dD�K	�)7�`D�%{�PI32Ȧ"���HW8a�fDBdIݓbF
\� ��H@0(Ȧ�ȒS�Ec@Ȣi���\(D�F��(E#4�PLb1�ĒA��yq��d�+�	�$����єPR2BFc@`31���Q%%I
��c&
5ݷ ���o�-�o0�O�
QVF@��/n�kfʳ���:{H]o������nǮ�y���T#7"���.�'��r����,lG+�w�7燼�o���xoxxx0oxx�_q�j��pT߄8�y�A�x��d�Ŝ��L*�Os�Z�E�T狛U�3oB�|�T�v��m�5a,�	��Y���76ג��Taհ��2q��E�]<�cw���f�[}mw�g�<��/��'� k��������@P��@���4-[�X�u䚥�nfnC��[N��E�R�#�Ʊ�A;�0�|�<-c��k�r�5��)��2��ja�j�T=���+���]5�|��r�ƥ���/@��dȗx1
C�z`M�'����0��p��SW�d���r쿾ϋ��:���ОO��ٮ[(椚��R��%�������K/�vVލ#PHJׯC�>0�ۜnY�N��쇝1>c��	@A�����E����Ӆ�D
Oum�٫rug<?!H3X��B�!�S�
h�O��a�<��p9*�!8��;F��l�UY����q�]�se�]J=1B��
A�#���\5X�����}���T��kdO͹��w��Q���OL�q���76�b��sS8��X�8Z=�����{�;.���G���r�s�����+� o�j\�R���6-�=;h:M�:�~�����Vb)��\��(Ki[�R����vem��G��qa.\鈩Y���4F��F���G]��^�^ѭ�\��ǜp�37ٝ��'I5�������ڤ���5�[bڊ�J�V��ѽ�o �<DB�ݟ"�ߓIl��Bd�O���*�g����ᩭ����q��p6���4�; �SY�xp���r;'�5�d:���ħ%B`����G���Y�`8�1���<!��i�wL�K��:�q��_�+�ƽ#�e'E�J:M1��&�%���m~Ow�c�eI��ȫ����'���\�p��ƽ�H�B�'{/)��R��g�3�Xf����Z���ߪk��ʻ(a�L�ΰ.l���ka����h
���^��Ɩ������/��6e��sl��q��C�P�@ۆؘmi���'f���6�����]v�bCJp@�8~�_�n}T~�3��uI��p�����@pX�\��=g����z�1%�{#���>��	fՈ*��{�J�)�z�>��Գm{��q����@�77i7�hi� �lc�\T厘<�Q�uȷQ�M��!n����eO��}8��g��@��1/A��Kg����̝�wv���,RA�2��2�Ӑ.�3[���9>m^}k!��Q���xi����M�VPc�a��(�.��A���Jj�f�+E�A~��x�/�	���k[�*��j���U���'+tW"�]E�J=Jl��/��7���$���S��m^'�"M�nY���9�J��7OFu�����-ܝs�ټ�[���`��x|����f��=�UF+آ��ʴW��<��u�������s�����%僅M�b�xwA�����}����f�Yƃ�ͬ`��r���K^Lt���['T�\^7:r�3�6$��(G�ԝ�е��Å-g�2��ѝ�^Cy��3�3��'%���׹�Y�ɚU�,:�YA
����i�2���1���\�����9��f��q�-�s�+���^%�S8ˊ�m��R�����|ؤ�1��>:�b��ek'��y��?�hx;���P��b��oc��^}��Jm�2ef$�꺏Ϩ�9���E������,����#K� ����E���
�D �P�Y���e*�&��CLsqRA�ܚ|�|����mt��%�s�����(X���^p�D�̒�:"S�>�b����&�ƞ����?p���g}��>�c�^c�6v�?bӹ��o�����JY����eXe�)�)�.�,&���I�#VP��G-.��fӣ�/"���cG��K��0R�p༎��q羕qO��|3��>��o}u�g�ZT�H�	��E��<�^��ˢXF zC�����=~$Nʙ��0� n��$|[Ty��ɮ.��}����4�A���#[ѧ}��}�%��ڷ�v�v&�L�)�x�{w�c����ه�]-�ܴS��Kw�3�Ku���Pdu�˖��0�W���0���+\�z�>��=�7����l��m�lcd�X��cjeTF�5�*ƶ5���mh֌Z�`�����{ϽZ�q��T�[��TK"�*�X�U�v0�/-H�0�
��'�q�Q-���~]�=��2iz�ڧ�e�Ƀݻ�']�z�s���Ơ�����I����o6)O�D3fT���Fx<*�Q88�t�0�.�f�v�����<it[Q��p�Vl	�������nk��C�'�a�I�dZ��aKϖӻ���c`��[���:��� >�u��f���i�l;j�K��v�,'�k8��/�c�w��h� ���(XXŰ'-q0�́;#Y.����Jq���=U[�5��n���ǨIQ%�x˱bN"6��80���n�?�J�Z��iL(_�Ц�e��y>�\��U�Σ��e�f�@����e�ԉ�kljO���,���3,�=�O={�9�S�r�XOql�ؚ���^Y	-����Q�g�n��"�2�"u�Mʭ�����Lt����e�x�F����P;�mEco9	��� ��@�/Y�UPl�ŧ}�E}[�$_KϽ�ⰽ����e]��hK�B}"���n�m�t밷��
��e���Bp:�l�'�E7�+ӗ�"�<hȟ����5X�	�������K���4~/u�R���?u9m;������>W��{f	G�5���S����M�ǁ�|q��ʗZӅd��P=TM)2Uʲ�x�������	�#{vF=;6SX~vȾx|�y����`F6�fh��ѵ��h�Q�V5����ck*�-�6�"���o��_����b�g8�#��B��TXSW���t�#�e�[�u3JcݾGc�hM٭#�aE�S�bކ{Y��c,�L��"S�IP��J
�#��Od[B����[:AÎ�a����,٘7jD�m*Wt� ֌;`�J�,/1V<�/Eq�lF<�RS�HtN�v�kkzl������3���� ����UeSמ����oئ�Y��9�o<��vk�D�.���싫z�;m�;*<A�R�/��7sк��=&�V߰�aUfW<5aj�/XS�te�ݰ�<v7'b$>&᪺�0�(�e؍k0<��	l/�ζMгnd㋾*��9��Ջ%�{�k�~�����Ú\��D�!���S�6�Ά�m���Y�#�naTR�՚�sk9qI���a(%���t����Ԙ������4ǃ�~��8H�[�z��A\k�&��*�t�=�i����<��{��ٛR���Mg��ZwMfy���/'_c����ߪ'Y��v�ÔXW��5�eԓ[aKnt���.�?~A*fa�l��	Ϊ�vqS��D)�d�tJ�oVF���;R걑غބ&vr������ή[��'g�[���~��pF��oF�:�evdw?f�޶�4v��XY�2�:�<YF�l]�V�R$~Q5�v⎛�sv�4�6lۚ��u�`33m��kmm�Vص����ǳa��'��<$.��E��W/M��;�d<�� ���|�Q!�U������
X�9��*b�&��P���;�
t�T���)�->�]�Z�X�^z9��J��['���fo<n+-��iζ#�c��Rq��x��֣�j���$7A�2�
�6n볹�Cpc@,�l�󇡽6�m�#�]��\��Aֳ����+D������X����BUKsPP����&T�@�2:2�L�ǫ1� Ĕ� �\5K`����L<���yXl���j�CH�S�]Je~/�����1�t.�d穌7Eqٶm�=�x��1&ck�]r'�Kv�U�(`�p!�kK��fRu��8�d]m�Lhi0���� �}��Y�|��vW�R�����h�˥�BzcC�*��w�1I��Qu����	@�Lf�?G>v~�66��;<�Hk(a��rf�u�sd>8���p�~�I�U�'�j�NL_^i�m��{���j�8�ܵ��j8�8� ����#�5��
�#�DO>�w7�&��s\��F~�y{ac�[�'������s�'�T�.h,^g��XؕZ;�-�Ǩo1����-0I]�]�P���0��s�Jje1���@SY�B7*t��iU�[�۾�x����%4#���M���7���n���gYW^f*fdb�mb�ɶ�J�s��t�咃�v��o4��X[|4��3����ï����c�	�L�P�@���cp��#3T����Upl[�o&t������%bU�N��[��.dG,n�L�^�)`q��3������
=�7Cm���6]���R#��+{ʱ��Lm�u>_)����j���f.ՙi$���4hʝ#��V�v�f"��W�.��E�֙h�˴�}}(�Xc��C���8�р�-U���9]�Pi��854t�[��x6����/����q�䅽z�e�.��VDVU$����`�d,>�Bg�bO�҄r);�`���Z��e����ws*��BY)n���3����[�����4�' ���YA
��Q@��O^�)�Yv22h�.h�k4i�t�|Y�-�Vg7ae?!5>�{5�l��"�;�[$2Y�����6)>�ռ*"��R��M�YJ�k]b��g�|�ȇ�y��N
����W�x�M��Pd��4���s��fo��=
�s��$�x�_w<I�߁q���`v�BA���B�I�nwA8�Q,�ߒSL���-w��P��k�|��Q@]o�Qw���޷�1['���{����ӜN��a�������%wӊ��|X1o���^��P�,�ޣ�<r���=���&���{^ _�Z_i��5/���CPMJ��^Š�7`i	E��jb���U��l��Qh�ƭ̪�����罫����g1�V~�y0Y�ѤM{��f�W0����ŸtbOǸ�޹��SV��(�<u��y�v��i4������JQ����i�~wf�{|�0�0[�M{v��2������;3Qw_R�|1���F�*��z,���`����yx�\��y�!�U�ri�'J-w���1@�����˵�M���-?,O ����u �i�O�H~�ь�q��R�6�����=����O����7g)Ʈe�ԍc@�@'�q����]�|�٤���`��t�8|����1a��hS���E��,p�z��\Cj����)?5�2m��J|�|�<�������_��Ժ��m�}�wfR��8�>0�i"�{L�p�
́= ��m�Nٝ:�2oLy]��;;ҽ5�̇?��>�>Hr�>�i�6��m��g>ϱ��+#%��ܼ��>0�>�v��8��M0�Ze{�W5�nX�q|S,,b�8�H	�Q���V�^]L��uۺʧ�icH��F,�^�4]�ö��Ո�aK{Z1y<����rW_�����p�R����ޙ��B��%��ǪcC��^�]�ۏ~=�7�,�1�3m~�\6�������pyf�n�P���"*S{Z���k��y�����x�x��'����%�y�}�8�#�?{��ko�ز��<���)�#%��(^1�ST������� f��f��7�����QKmh���Ljsr�m�<7�זe�sL�v��� ԉ�i�֞^��<C~�WCd���˛##~�̔�(X4k�����j-�m��Dm.�U���:�T�jC7vK���!cNi��m�BX�}0L�^B��0]�7fP	�y��.��t��kȘ�]ѓVe�#Nz��ߔa��l8�~CN���R
͈��+��ˣY6��\��L3h]N+�O jf��D1�[qE��"QUE�7\)j�R�@�LS������f�r��L���1�S���ԕٺ��Z��X�z$����r�H���]���Ы��$�3t�iE�N�]��ղs�r(1�R�����]�M*L���_��Qz�\h�t�zw�xat��w<[�&�V�>�l �"�cO��W5!�0Ǆ��eN�,Ԥ�|��]��-灱��~�r!�m�����sL� M�A��Q�A�\�.��0iհ���+a0��+����^K1�0�Un����q���ӵN�wK2�F��i��͒	��s�:�7B͇2q�����!�W&{��h�����h���JדIU��toe�Ң�zo*i��c}��[�Ğlٳ�nv ��\3 m��j����;��[����y3]�����p_	�c���{3��u�k�ܫ�0����	V��9�.�,y[��8�t�_��?��ߟ����Ѩ��EV����|]��W��X_��8��'��^緬�yWW�p~��r�_�N�m��\�˛�����v���$���1�Z�R�2������{hd��A���b4^��n���!{gs���I|�,ʼ�<v˲�&�0�@��6�9C��5-� n!:u�1�A#p["VY���C���lK���{B���iR-�wE�ǣ�XW��\e۱��4��0��1X���|eN�>V����ll�%xP��*�Yi��^��� �BiN���n��F�3�f)�L+�g��:^�w0�b�]�-�9<��Z�X����S��6i=vV{՝i)(��k~�v=%{l����<*�ň���I�<Վ��P�
XHn�$)��24d�8�қ�fu4J��[Z��:��aTe
6Up`^<�yu�Z�(p\��Aֳ[�ewN�9u�r�s�Nn��x�F���nj��"Se�R*b�I��H��5�;�k:�W�ԶG׳g�v��P1��_���PsS>�� �/��WB�X/��	�b��q�x�4{=>�_����������_����{}P�iM�0"�E��#1	���O�"kX���Po�Χ�S��]��m�>���Z'���k[�M���^Ӷ�"Y�s[='��7M�P8�ë���)صlݷ�(�b��.��%Z�ňxry�Fg�<�.��Ѿ5��2�޴�N�X�F*���r=V=�����n����MC�w��\�y5�źx��=n%�Ý�����y#��!�b0=��>�����W����G��?�Ea�ۑ]��V��,)>C���{6�>Y�� 1b�l��~�v1)\\d�E�s�b�e���j�/V�8�:�ќ��z�o�,������y����j�1R{�^!�?D4�
��W�0y�0*��}��x|p�w9-��%7��� >��od=}w����̓��z���~T�ڢ
{s�ӈ�^�v������Q��<��y3���U������e�x�C�v9��sI��|����I�x'K
���"���dr��GMw�5o�û�.o4vy7���CE�r�JԳ�w�
��8�Ҿ:1c��x������y�b��r��{ӹ��y|�_{�v�x��u���I��Oj'Jozq,�%�+U�򣇪u����it��F.{vv��@�����d�W�J���M!p����|3AG`#����	P��l:��uJ�g�����#���U�[������L�XwCQ�=~�7����&Y��m�����;%����I��{s
F�v�=�Y��
� �{(��N�\�q^3hpUq��Zϳ�L��ۼɵ��;]��P+���R�K�7<��f�؉��M���ζ��ga�QI����X��2d"���ںޮ�ۈ�"���% �%F�K%w�u4��о� X5�jC�����~gL������=]aUE���r�0h�{/U˦��ta}瓀՝m	j&�G��)�f�f�|<x���S���$��M�����5wS0 ��:}���#���n��q�xG��؆��g���v3�8�Ƽi�8;��_���C�^h_w!����[&�x���Ȧ}��m1�������g.p��xp+ٲ�V��O+)�N�i�ęb����fݨ�<�ޣל\w��)��\�ک����3��%��f��7����o,`^��[�����=��;�����g��V�Vӝ�~��5��w���z��Ol|�`o9]g���R՘H��zw>�f�?Y�]�8vD�����t2�@�ҷ�4�cz�Ӽ�q�aȊs��^'^R��9��{�v4��rݬi�ë�8XRd鲝 �&ɴ?6��z�|M��l��� $�^s�+���r�i�f��X���=�������/`�L!X��-�}ӨDS�-��g����<�Z�n����,EOQ�ȷ�����%vgn9�]:��H�}�=�ڔuv��F��ϱ��yԳ�:̫��f�#�����������wu��׿��
̒R�]LŌ�D�2�(`������ێus�d�rcB���& �э32҈BQ&>�1]���#"I0�X�Jh��is�"3D�"Ј"(�3)(Dw]�@A!��0I�iF,��d�I���Jŀ�\�fJJ��]�B�1�	�$(	�"j)�Lf��
�d�&D�P�i ц��m2��F`�S4mbd��M�vJ@e&$L�fF�aJ*I�(HAD�"����bI"�#F�9���Q1�H4�,bM	@�MD�T	�B�KHE#,Q�@2L�b�f"��IHķ�����_���~uߟ�y�W����}��rh=��t˰��s����k8�lݯ����;�)�>t��3^��zv��F�ʽTi����a"�F6��	8@A�,A�ZD:7���0oxxET�Þ��<�d�#�
��6���E2z��T�
8���3��2���YY�ǇV�=M�-�g䲠���K��/�՜�eX�1�����.|����$J�4���b�����G����~����������������#VA֏� �G0nLɎ��=!1�a�Jh��eֵ^[��{:&2��]š�����Ӊ�|�rQ�GZ=d9{mn/b`y���[bG�ݬ�xs59�k)�*L�Յe	�ލF=<����@�1Ԇ6��c�H�+a���If�`�g��j����\؝��J�dc��2t��i�8�%�\�l��m�SM�H�;{{�K���7����g9w��v@���-�Y�U�t�f��2 B4��(�|��}8�b9��5��}�}��-�5�	���R�W��m]�W�.�轚�/h���ۆkq8��$6�>�Z�+zr�A�l��Y��.o�~�<�{�klZhbrW��ZW�S��ګ=՛ �To���n����uMf��j�=��h}܄ϦğY.�^D��ZYr���9�z]���e�ƭ�<�Lrs��V�{zR���ų�� D�<ω�[�8#�y�'g��^�h*�U�e���%��Gm�y�8��̦"WV0ɠJ�*+́f7��X�ҫ���0�5�Qz7$�	�s͖���qr�i>��	^2��C� {s'���~����7g�����n}V�>&�4��4�4;$���YA
ɇ>��OX^Jg]�B�v~i=��&����7�Z�F"�B�No�S�/^��Ơ�*f�eT�q�b�H}�i�������b���t���7Mprxk! �
��E*�`��j+�7���c��ɩb����}<��9Bb�gqj�k����ĕ�'<�EH����7A��q��>5�K�9;v�-ŘL2��}VT_0̝��z}h�%�i������$���XS�U���r�s�X�N>�"��t���Y�%�{3��������z���F���,��j0�W�/53K?�s�\=�Z.�78��}}r�h�h1�}u3�JS���*I��fa9X9�Q�<Û���#ϲE�����Tz�N�����q�M�kئړ�.��M���-?,O ��7��]�@~���w��+�z�f��V���*g��Zv�2%��3�k]�^*ԍcEGsׂ|wڢ���clҿ"���6�g}���,� ��<�!دAV(Т�rdSM[]�i�^Q͒��y�?���'U1|Xn���5��?����{;yҪ���u[#�=kY��ky����K��G����,UW:�1~���N �PԈ�ґ�X[iw6y��OQ���Y��"�v�*�]6Ý&.Qvt�c����P�L�Ӿ�c�u\�Js��_J[��[c�3�v����z��閫9gw���fY�)I,���10\ip�Y�0����hZ�R�wJ�K��̤�/k�/7ח��G�y�/�1�i��2-��|A��1�sS:6եY<le��+J��Q��Jʫ:ľ�7��b.{5F48$�G��$,)�1ju�h]a�a���-֞c'^]�O\���swH��p��\f��2�X��q�DYz�o�Wf}�\�>�P�6���4�ˁ�F��6��,�ru�r_���f?������%�(�A�0Ә��=p�ۍ-P9�um�I�맾�*�\A+�-�i��RݯsW>��حja ��Ÿ���os��M}���r/������[F���36��M�qp�Q�ˍ��E4v-q��{�t�1To97��}"ُ3�p͘�05d�h�R�ǥb8r��v���;������8߃%��u�aO㮲!:�9E'KT�D*��������*��8Z�C��4�R�ֈ��D�Z���ͥ%۶�V��j�)�9w��J��UE?��E0�zh]Ӎ��x�k����zN�.�H�������G'���RQ�/��_�Y��w����|.sŰ�ua�3{epuR�잔�UMf���^��2���4X�+����wz;��?[q�؃ӌ�R�m�\���'_������՞S]#�����`��`��o�>��D(A�_K2 _v�4�2�^b��E�)��*��/fg��;��=���q7~	��׆p�|gd�OH �zpȦV0�v�5)<�d] ^3վ�G.��֪j��}yG�]'��'X�r��Gk�9��'���n� Ja<,���5m�"�`:�5�ߣ�3p��)�v��fʯ$L�5�`y��Hsf�|Bgƻ�Q���m�y��Q�9'�D�?�8�Qa^���f�V�Mrc��NF�`�5�y�����ڵ�2 K-�[v�B���B����-Xr�M�8.���A/m~~Xí¶�2	���y���@�k��1��U{YgE*d >'�0�s�0�)P6˦��ܡ�r���02޼^�>�5(�b���]��k/���W�.`�R�;!��w�E�+j5���KG�_.,���ƿi�y�)Wݤ���?Hk��Ԅ���K��HQ�
��\i�������vy�ӄ=X� �����d<�,�j�./4 ���t�@�m����1��;�S�8UO�e�Mi�V����|%Z#�K6_O��_�|�2���f�~Cw�����${U��ov��a�fl��{��0�����^�_R������9l�mBl�拋��\��X�s�Sz�<\4Uҭ����&�/%�gYGgg$ ���v���>�޳�
�� (�qӝ�sVs���ƫ���/��p��#g����5ԣq�P�PZ��$��K�f�4�u{����qc�T�5x.R=��J�Ne
6
����.�� ��xkk�w�Jw�~�y^�XSo�t����+_��=���s���Bk�1K
N��Ei��z�ot�#�H�ޅG�vMe�c�� B�Ӯ%� �}>!���y��	L�<'<T�	��J�h,����Q�Mt�J���͞�;&��ɜA�Sc�g4��bH�[���$�,���g
A͟UT-~���P������1w���z&P�'��kH.͗�.z����$J�,�w���}7}���^����^�tgk��<޼���� j�:���� �p��M>X/��	�3��ۜ��:�N�����/c�{��1�x�f��m�� �k��{<���S���{JY�И9����H�a�kj��O��SlV�.�ǣQ���uߜf�'�wL�W��"cu2V�����ז��/�	^D��'f�Lt��\�a>�ҵ�9/R�Xæj^>۱fi�lj�hbԳ�RmT=��k<G�_����R���)�q��a�|s�cn��I�?I�s{���.v~٪.��v�@t:��3��W4\��bB��^E@���T5��->��xpN�1p�k�%\��^��ܽ��Ȏ`�}��C2�CWz��y���������8`�P�
i3�l�W���F�<����������FE9ȧ0��Z�{�{aKu�3r
,3��`3�B��K�^�i��x�����r�Z�0�0z�g�]<�e���b*s���P��2B-���C�������}����}j��<CK���|����9Cz�b��Y����� ��^�R-�N�xd�8R�T�S��FQ�ٛ���^)�daqCY�������j�A�Q�1��Jkd�D�K#*ڛ����N�[Y&���sbj})��g�%L�vd�-�2(���6��Y�M(I7Zs5O< R)�48��a�<����j��[/>��D���(2jX������=�hF��qV���]���ئ�ǌ�ГD��=�%�Hn��hh�S�c@ĸq8t.	�Ұ���Q莮�%��xSLl*4���o�C���A�S�B���f�r��N4&ln���CN��g9���lD�I˼'%t�cC{c�ZVK�G�)G�b�jf�.�f��?{.����<��?�����L�W���g�|�y����j#�+��5������v=`-���h[����򽡞5Ӧ�/���ㄕR��q�]d���nˎ�κܺ���{=�ᜀ�XYT�������&2N$��j����Yt�ؾ���O�?7���m}A��3��.�}��$�b)9Y��6+�cG�ϵH)xߌ����_#��u,z����ezT�Ɔt�R{��
a�Y��C�Z~X�A/^�R:�M0��칐�B�ܾ巳�>��-�Ϙ(֑�8�Fı��n�S�]�Q*=<��Q�o/g���kV�
��Rz����b����$_JrYj�,�hc�~�vOƧ�W:�I�Lk�M[]锟�E�h�i'(T_3��r������^�wf��$�[��#A��ipk=�ٙ1�<(��{v;����@�����XH�-�����/<Ų����!ۤt0c�����ZQ��8��|C��&;:���7\�u'�;�!�$��df�q��g���t2\�Y��/<�e�K��<����s�۬��k����r�k%{��@ÝBhq�.�8˱i�C�DN��Z.���R5�٥�^C���d��9p�,gN����Mrv�c�/,�4֙'�iN���3�[ͭ��V֮��6��;:Z4������q�����$>F5����WX�Z��A�������ɦݒ���q���� ���0_{�Rs`����3�3rǽ���nyۚ����A�2���ú߂��u�ٜU,�&NU�hnV�@��4�C)I)f�ہkW��b`���ư�����ٮ&Ϟ��.1wo�V)N5�{$����J;-���=;��6���k��{cV��H�:sՌ���5��ȇ�zaB&�#c*+KL�M�v�k�+��7u�Ď}d1G�@�'����4��P��A��1�	�O�گG3��*�w�Ѭ��Zŗ���N�2���-T))��YeE���:��s"zU#!�K�NG�޼���Lք�"�BԳp�})���~ �Jsi+
d��:m��E�*���m��^r�s����8P�i�l���m�]�i�I��m�(���"*��/�p�wHf=��f�"(���`f�}����Z�3�Q�������ZTC8���/9�-�zښ)8>8alL���7/4CwU u�af�8h�,��!�`C�n�'����t(�L*����:���["%�V�6Bs{���!������;n�K2�R4\i��lu�7�|Ͼ{b疚Ko�����T���+]�U-t��:�|��>��H(Y��06��S�����Eʺ��J�;(Z���Y"�V#Bպ��:۱�̍�e��cp�0�'b'�ݘ�-��ߝ۞��.\c�xR�y����m�n����.�BWӉQ,h� ��n=��P�N֮Dh��J�K��`���D�A8���>��rS�Z�Lf	��Y�c�a��,�f��tF�=fQ��u�\��l�c)�(�c�R�na��Ε�C_Â�B�ucq1������ya���[�| =���v��gRa�C
T��{��s��s?M�춢���M�#��z�%����ɡ�ใrrCӖ�=x�d�0�ͪ�~�츰Q*���s�k�)�1=Vf?&�T���%�:^˓�HP,*��E��#���h^Aa4gE�D�<)>=���5����ϓ�u~�ݵ�Zo�by)���}CP~t�U?q��4m��w���M��.����n��C:	-@�^�Y!L���)�t=C�yg�X)��{�8^wrD񩛦�竵=��PZ��T�5.2=�veK2� �<��zm��skDS89\��N%5if��ʱ�ɰ#�������ݐ���M{�BeAb�I�Wm�zs^�4A����M0�&v�0wp�E�k;X��l�A�逐��q~!�g)-@�̬�JseJ`�U��%�R%r���l���qU�M���n��h��%���C�O|�ƽ#L�N���/ش�wE>��'/5���g"�y���q6�~L(>(� �ZbͲ53S���;�c�g�V?//]L���]d�n2D�8�2C6x�V���:U���܂/���b��\��A(p��~���CTE�>��7 ��ed{s9LéM�"�!Y7�ƙoN�([��º�M�w��6����M���:k�-�B�o.�Sڌ���5�zVM[�$ ���vf��N�r�Eֳ�rz���u>���L���sdkT�C3%�����frj�ʹ(��x��J���������<q���[c��hC�V���S�Ժ����a���œ�kC(�	���4�X�6��xa9B��Uz���
��j_/]i��K[����L��9o��Э�8a�ȃ�z=фD�vzM&���c
�ҵ����{�ܚ�C��g�[��_m�f�2-����!��f�E��:�Z���<�����r��п�C��s��A4|�Ͽog�wz�}r�ڽ����c�P+�.�٭2�}�S}Wl�~�aU�dz�%�,o�S��j��1��ef��m��!�*pr�Cap�����f�}N혶�n����Qu%]揀��Z�@�C���h}܄�� �E��Rv.���W|*gf)�\�+I�+�ΉZ��Ǟսjޡ�#73M�,:��PFL8y�㌠�;�,�9�~����;w�Ǵ,gk	�������Q��ٜj<�3u��,�`X�������^�w������}��o���������s�j�+�֪VN-�zA(E����b�4�ph��S��WcI��%`�c���8d��+/J����E��dcn���=�[Jւ� �7q��oo����/��1>�[x��P�>����C�˽���)���u-��dֲ���\���p��n��i�l��M�K�X��nn�r^���NX#���p"'�|6�nn{�iOUg�'�O�o����#�7�a��VfҵǽWb�k���f3���.νK;2e�I3&{�3���)ڊ���{AU�=�/O 2Ny�'�ѝco���t�.]��8f��v_.W��C��qs�6L+}�v�nɿv1�BК����+�������wo���"���$�,pc�/z������!�ᤞgם^��q�V=�\���ui���hQN�n�T/gu��%��b.W�-����ۦ��U�4�\�*���v!��k�3�7He�4�5�ֺ�K9׵i�I	+�2��re�!�_:Ƅ���^5�;gv��Qqs�:����m��9=�ӹQ��D�C��ƈ�݈�.��#Z����������g���Q��X��Y���I���-^���.d�b;|^���:ANi��Q�wHZ�Y�o�vC���f���?O��^���z�Ix�ܕc��[��1�	*����@���b�x�8^���*�x�*�N�������_�7������r<��:�U���pY��*5�y�QX�7���;lc�;	���8]��ي7q��-r�3��I��՗�+X�z��ĺ͂��9��s���jo\= �}��,a�֚s�м�7fr�<P#:�W��|3����9|�����GdW�N�<w�9�7Ӕ�!�8�4,���{R���_f���Ž�_P�y6���˂���K8@��.�E�{ �i�Į��n��m�����9�_f�ř(��bٝ�{y����;D����s�M�pc���g`���iڠ*-XYg-�ɜ��������N��+����<��Ԝ��іT4���6f���F���|]uf"��މC��E$艹qo�nxU�rKj��`�:�%��%�ճ�dȆ�j�]=X�u��^n�_&�v��
�=���a'j�%��d�5�q���'d�S��uPB̚�8��n[���r��⧏�n,��݇¯,���;���r>>B�T��t{n��ۤR���G��������9��w)_���b�Nt���%�p
�1�"�>���a<Oi���+j�إ�4�r���NH)����Y��J�d��l����rY;�=�P�"�ů�	 _���4���������z����;巟K�v{}\�4�͂Y�뻇�7�5_cX�_A���mW^tw�o˝-1*�as�!k�s��ru����������}�>�*�Y��g-�ӛ�Z�Ы$QIfX��IR��@ȀB������a��2��%�n2ai����a#4FfL`�1�h�"�@0�DDd�IH"ɨ�����J1��jK������b26L����F���b���ȄP�-	`S(�i��*"0�I��"H��
��I0F@�`�wF	�D�5IL��t�c�ѹr #&���!�X̍y�VL�(�F 2� `��Q�)�F4^눣/+�F4�u�*#d��ˢP	F4�$a��F��cE봦�!$�@�f)F��7����0i�����g#ه�����n���z���q�
�����T�H��P��s�L�5�x����n[jU���l��W��2������?q�*�A*����2|�s����p��7����d͸�d�;V�ԫ��W���'�-�v)�LI\`I�xq"��" Wl�2�D�-�t������l����S6sQ�Q,y�%4�£I�BW&�0�/�2J57��r},Ԙ�����:P��}�"����z�_V��z"S���b%9]X��F�[X��ƃJQ��/��il��c+�gE;�Tuv�S�͑q>���K02,�w��$��S���Q����5�/A�<���	�.�s=\\���9�S�:YP���:m���R�l�S�(���<�^��ZG&�%
��1�m���ʪ��ts�۸À}@�
Xs��lkǆAbv�2���Z׆x����,��
��t���
Qѷ��'Z[ņw'%���4\�w=�C�~5=B��ɟ
ba�f��kZ�&a�k��!�j8Z:M^�:���R�eߗ����Ԓ�oi���4��E�����]�j]�#yW�GGnY��v:S�
�c��G�:LW5�a��d[0�h�q�B�֯7���=R�!ϔp��o�m�OS:�W��� j����h�KzaR�ksWup�D�Bv���B��{�3k삫p���s�?���^�&��*:[&�'�2�mӺ�(W��sR�k����(zNۼ�7S
�m^F���v��p4j�3���w*G���������q��>�6酌6��İ�-���+��/�ζ�D�)�=y=��\Oc�x��Yx���=	�X�s�5���A���s�Mz�՗n0퍠��q �/��)(۲m��,�����i��U���M��p������X��m�9�>��,Ӛd�j�S��d�xA����ż#;�Ғ/m�1YX*��%dq��
�4�n�O���.�k-t���ݎq��eV���C>�o偩��Xn��ƭCu�ǋ��j�J�ﳷ�t?o�z�t_]���[�S��[��YgB	���['���+����M���9٤�9	�VQWyl���P�P�w��+�㥻�O���nĀ!���QIխT)XUE�5ym�5uEáGU��w�߼�[(} i��x�ｪY�3��^�2�X���L��xNy%B��U�ߢ�Dѹ���5��-�wX�m-h��o@��cL:9��2�fY�4��.Ӧ�&Y��l9��.Ճ[iϟ��?K�I�"?S�����sn����Ɛ!�O�= �����*���$�>����S����K+#���������r_7="Y�Xh��Wb�w,��Ծ~�ӽ�*x��/C3:G�!|�u�e��L�ْ�V�|ڨT����Ts�ǝU˒�ݦ�y�J˅[�=�ZF�d������,Њ�nM�.�b�zs	�⺅?-2[�d*�m^n�?�l����j_W�Φ<�LY��g��GY#���v@}�������3�\V���7�����E���X�͕&���a�<;�w�`�ݡ���p[��Ӟ��)�#U���7�]9��S�X��qTXP���f�V����>ܱ���ʺ��c��'ݰ��}�eyhX���2mJ��hg�B����s7y�c��цA9�η)xf�u��l��!���4��������,9�aJ��t�X���+�KsU����ٙ����ZN���e���p��P(`\����N[���-�[Ti�q�.ɭ�X�SF�l���SϹ�o{�'<']�?XRلC4,�(p҃�
��/Ƙ�M�V傺9	�v�W���D���A��� ��8�`�xm�A����� ̮�N��8�B����Bg>��n�+=P���+}+:�[���Y!
^i��S������������K�5��5�mm����ƣc*���.29�A�Y�(�'\?oM����s'㶪�r��1�C՚4o���ٓ���dGߎv�����&]�����^g�Ez���z!��Ξf]_�R���Qe/.Ѝ �3�zg�X���0wӹ)mvz�^� Gv���,�u�PM:X͖�>C�w9�&$�/u����ӗm����3�},�	�N	�iAv�����ږ澂%6w�HL��
Oj�h_l�lt4�<���ܻ��j�[Զ�Zmᥩ��C��Aq(>T�HM�x��/��WB�G�ģ��#�	��:�Q�7�v0��{�mD����Ě% ��d4�P�g,Nl{��I,���pd�f���U�m�aNۧ�*w��� mF ̺��X��58K�v����0�)��"������ՠ���Іʓ�ڊN�_���OW��z��f�s����Q��c��-�W.��i'�5����H��'qUeWC�zM��)�{���sA�����d0���=[Ok���Z�D!	��f���6��r+x��c�yfw���:�Ŗ`j�`�1�M���V���{�����;^D���M����W	V57.��eA/r�'f�a��Q���g�397�vl�r�\c�F@��f�>&�5+E��;�l�AT����k��pl�=�e��;Q/��q�)�jnY����@�!��j��3�_iVO���NX�wce?6���e��r^��\��t��{����������d{b��~���`�ܟ�!��(��}C��/y�Eo�5g�oN��l�R픷,�H6�����-�N2hm�$�B�;;]����-�q��ش��/�ww���n��7�Q�!������IС���!����u�im��f�Ut� ��՝�{�-ק#��C���	�`;��hp7rkX������X;Bcs�w�Xms���he�+�ۆ��
�a���˺�R�~뾕�����PB�2a�ȼy��M��Ji�MvN�¾ۧ��)��]�����i栩TS�z؋`�,ځ�A�,�`[�D^+Ex��4�������H�Հ�?����Et
q�@�e ��'���)�t��G���W}o��c�Q�V��r33��|��w�5��*a{�}V�Q�*�I�WB�`�ar"!�.�u��;�w:\mn.��כ�Z����K"���+Q�i&��W��/�2J�B��,�3yjБ��U�����`�T��H����:"S��D�6H�%MM��<�&3���o�1|r׼�{��oY��(̬�ɚ�7,�BT�e���2���I>I��yhb�a�F�Ӆ�6u�.�����E\w�x���yլ�3�ڋ�.��tڟ��~D'�K���s��b�ow�j��#"��w�f�U|h��8�;�͓�l�1��'�M�����O]��GB�7��w�ep���H�j��nQ��vcY7H�z�nx髕^$-y�נ�4�W�nLn�4�v�E}].��\��<<9#5�G729�L=��܉a�F��-��6���x���2%�EgE��k���Ŧ�:�T���G+����e�$��/#6j$e�rYb�,C09��qͧȡ3��#��g���}�5�W>�Z���B;_d��?�f�0K5��10Zip�Y�8������!��B���M�\�]:���*�����ﳣkT��@E���Ǣ9��o2z<ϩ�w6��-hV��sГ�{T��i'���-���sQ~������}��Ύ��K�U7U���1hq�'�,������c�c��s���e���eAb��zyeL�lS��tA�/%iO��S�B��yj��=�f>y�~M|.�T]�e�>�[�}�M#���O�N\^v����v�4�4i�PW`�J��w~��]Y�{7����؎(;��RU���k���D�
����!�oլ������<_'�Q\qp��]bX.�|����.Y䣐)�W���7�� ����!�nc^+�Y��[�Pʋ��C4��!;��΅3��q�+p�͗N�2�s�Fa�HA�u��Z��ۯ)�S�G��ʮ"�]ONh��DX֍��f����ҍ�r����f �U7P΍ž>VBO�ˊ���8�fZ�ԞU�w��Q��t�&�b�(m��[�Wc#����v 㝎u�$��������<)y����o7%}��~���>�:��2as����RukU
V��
j�nq�^�Ы6��3k�4�\��ܛ�۞Lx`\�BV�4�r�K@��n��,Z�D&I��Js~IP�`*��\�5��2�r-U�n4���k�Qm
��zGƱPq>��P��b�öi�I�x��Wt�h[a�;���OF+����V�@���lRS�Apੋh����װ��T,�vhL�4�r.��:�d6�Ѭ0�z���P/�V���;5���e�0�2�نq����fN�����'��_v�P�I�P�s�D��i}孻�ۄ���f�&��A���M�-�3*0�g:�����U�V�M�'P�E-d߲qSl)lkt�J��k��ja��yWW������w+��M�]h�B��`e��w��6�|p�ڬ���V8��	Z�9/L}*9���'[���5��{��v�qoW�rb��a�A�����@�4���zv]��Ia��l�k��E�^���4cgo\e\���T��]!8c��:���C�la)\���,���v�Q`|�x,�2]W!�m���NL�L��{��|��o#��Ġ�Y+�mo\R�v�q��lꊽ��'G�����tv�c���eu�w�Iӹ#�{K����6@�&e$��VFᛁ� 
1s`kz�-��^���+W��fk��z���X�)m�p>3���El�?\W�����@��ox(��2��S�]�wM�6��NYrWA��^J�����u�i���'rc���/��w������p<�Ht�Ƕ!���u6p��A�pS�Y���<��Q�q4�ߏ�m���������]��՝c�/A,��&|�.2�7C�:�|+��Ա�婫�+B,�~N&.��_N�*����y���2��(Q�G�=oM�́�԰#X�MΙ�6M���r^Yֈ�Ɯ�z���v�zu�X��nj�"Sg(	���B��ƲB0�������3{2�Dv�՘�S8�,Y{�g�A�t���jJe��ڝ��!�`z"������y�2����~�y�n���I#�K!Ǹ�(h���^���l��fv�B����2��S�i�lP����qFe��l�K6_��6��9ѱ��iD�m{D(Z��"�RtÔ�.��cKz���th ��Q�<���y6�U�5��v�,��F�M�*BeXn��I�U�=�,h���PX��0���p���o]I���~�G��d#������/X���Ԃz���/�f���N��R�#�}���rbh��f��q��D[���$��[~�[�v���y�7]�� ������H�$�T1�1��O5��ƨsrq��+���w��z��p�t���,ݭ_ߪ8ߓ���=��U]o�:mi�eS�I����0-�܊��Q��Z��3b����\C)[wX�v�us�ۄ� ���m�K^@��z���j��-l�)��]+_#�Y���-���>ħ����=�߼G]�SM�I�a�`�
�K�"�y�*E��Mo[��ǗS�}i
��R�蔟?_������&k�4{n]�t�b�CP>$��
!/(�z��l�l|g(N4j�GX��u'�;���(�[���Y�^�1^�t(mh�HE�
& �u������c
������ʱՄk�ʬ�P̀u��&p/V�9�F���L��bO�ZP�_tz.8��;�o�y+%��F��}S�F2���{;�5�ٸi�kݒXu%�Z�yMͫ���P�f" �d�6"�r:4������ةY����1�Nv����z��Ư.J�f�;(2����fp��?�1�>��YIug�񘯆o�N����[E�E�.=<)Uc���bn�ׯ<hZY9|��f�\ڽ�x1jX���UӬ n)�bJ�-D���S��v�!���U=��i�	K%�d����)H��6<s�T�5�飭�--��8��@�ۭ����¦9[������g�Tv��8���G�b�t�'�c��'�.�j���+Or�ż�$�܅��d������딫<�H��8Nו�F����kK�3/�~( _�x-���GA�o��A8��%�{)M2Re5tF��cC4 �(8�*�!�݀�z���]N[�Qf��XdhB�N?i�W㚓���� ��斟H|U�jQ��t���K�2̠#9���X��yp�f��B2̣a[�Y��	�`�J�|1���F��.��|�ޯz!�/|���/�g�W���)a�A� w�sZ����c�F���i�M��Z~Y:A���R~Λ�l�˾k�y���P]4�A���-��i��+N݆_%�EgE����ܢye��v;/׺N�,29��Q�Л�@�������ap�q̀ F:|�N͛{}�Idh��؄1B9U������k엟G?�f���%��h0�s�dyE����{���L2"�Z��Fg���hZ�R�p/����O�`��i}����+r�˫��]���_}����wʾ���YC��z��/��C�a������B�K�G={O_������u�2�ܢ�{����bǀ���!Ö���q����J�ޠ��0�P��4v�Ż����x�=^�/o����{}��o���s��o/E��Ó%�M[��	WX��r�����K�R�`��̥�/&�����c�T<�S�Ae�xC.�%�x$�X:$�=��O\�/^��vxl\>��?%����Վ{��|5�۾�Vx{�c>8��!3�SΈ��}���[W@)7�Gn"�k�s��P��q�&-�Z_px��}�g�=Z7�930vV���T�z6�����ҕf��n��N�$�v�p5z���k`��p��[�n<¿eo#��a�.��&5=|۴�Oo��x���	þ�u ���u�C�D��w}o����΀����i�����>��Ȏ�N���l';؆�{�'�ٱ�q�/RD���39]��y�e����P4��P��j���ފ�?H��ܱH�;Xe��[�ɕ�����Z}&�]���Y�x��g	c:q �|V��,��o�z{�c�=7��p�a樲OH@��l���2or3(�����6Ĳ0ˍ�?o�%E�A���٣m��.�bt�SFc��՞T��' ]ξ���ԟ���g�ZƱ��:�^K5k��.�w�nB���9MV`��s�9^�c2�oT��Ri~��m,�i����������ȅ�sf21�f�7�M�x��t�j����c���*��bH#��Cj�B��u����Oq�Nv�(�'Fq�9X�?`WZ���{;���go[���Tf��喃�=k��,�44nV�϶g�_3E�s���yA��
i�m��x9}���ܿq�*c�w8Cq�d|��x�u��)���z��k�k8K���/eӦ��w/�R�ټ�]x�{�H����v�G.�,�m�"�Ƴh�[�s\Ly`��sbC���d�5�t�Y��o��l��>^��<�g�'�S�;�p�Hxc���u�}�Z�t�>����Y!��u3!���.�Ǣb�C�=���>,ɽ�,�.����wdK:դ��^��q.�v��1�z��+���t��L���}�ީ�{4*�v�~Yw��j&�����1x�Nu�Y���-x�g�r�]��%�w��VU�}���������<}�JNl��}�ؠqxn�y{],%��MF��u"����/�>�X�^'�9^�:z��ǁG��E��������LO � s�!�}5M�8]o����_O]�²���M]ݳb��ĉ]�j��pLp�{j���*Z���ͺ�:��c��z/x��Q��nD'.�>ҥ��<����Ѯݾ�h�^�K���g���;�E����Ն6�'����ӎ�%�z�:5���9Vz
�ho{ބ��+ŀ��ҧ��<��}��s��$:���%��:��,�f�X�nr��ո��k?��r����^�~wi۬ҥ�)v��i��`	����w��#�$ƇBi7�����Ә쨠��8@{��k�����2��1Ez��2V(5`� ���}2p��t M�o�um?זA?_������LS�&߶�`j*1H˻��Q���\��PFH
�D��"3$�0b�&�D(@B"أPF,E��,���*L�Q(�y�3���$JAD�H�+\D�RW.�HB�Ff�D�9\�1��B�W1��s�cc~�5�f̆N�$B0Q_��y�H��PC�BEH�(�&�dB�cdFc0��!��R�*D����!�HT�7��(�M&��\�F�Er� �4�H4�Y�ņbW."s�"d,�߯w�l��Y�����$"�T�iݹF����翏^�u꽹��N�{�07���;Ҍ�r�N�@�2��0��5����/-A���WPjvV=�/���)�T��ּG��nx# ��u&��A���	��㙄��̍�6��I�c��ra�^J�A��j�+�u�yb��;�����3DX)���)W}�,ݐ(�#/�O����y4��A[h97CPw੃I��b�{�5O9�v&M蓼=�n},������M^+$���4���6ʲ���3M{ir���ϡE>��*Ղ��ֽ���:��z'�`eEc.r�q�A<{�m�Ǧ:n�P��A�s8�7�v�zx~�O�y}����	^B%8U1��^�dՓ��!Z��):��P�~UE�5�8��$�˦QJ��!m��F0�p���-vi��w��f���Z�D&I��"S�	*��q�y6�g���9��z9�YC�|n���M����0��j�2�fY�k�٦�}Q��W� h��}�R}+8����w�)��(RG�s`l�y��GЋ	�A4���BzA�a�,��X�8T�w��&�t���
|׀ܥ��*V<�d]w��������0N1�� �.u�	�n�a�m�O6���)�����R�sR$ْ�k���/Z�E�ʒƑچû2|�4`�k����m�t�3/�&��{c���o;A�k\�2�^�}�l��*N��fT�3�)y�[�-&CZ��x������K�����j�>��]R���(��g�4�^.�OX�]w�������s���J�6<I#��u?6�.�h|E�mz���6��Q�*�=2� %��%0�̾4���{����~i���?"��&):�7B͹��.��,*�O1��X&�������u6���I�ܞ�w��0dC�r:liU=#�hg�Ԭq�t,~A/m~���M���A����^��Y�8]�5���a���y���� k��E��X[h^��^����K��|mcߋ
>s�{�rkn�N���u�Ò�@�<�<R�9/N[�׈�(��SW&^*��,��-Fo=�ʘ!�'���˷c׸��Lpb�M�'����Y��1�c�0��*7���y�QK��o�v�[DӰ�yC�{L�C�J�za���eF&��ڃ1��>���'�tSteaܨ��VGyn�q�𦌴ݤ,����e-{�4"k�"�)�P鋇P�$��T]���z��c�B�P=�8
e��*h�wM-��-tvd��IҨ��z�P֨�kb�Z����;�u}�<���b���-�>�0Z}#��l�%~��nnr!5����;Lטv���������k>a�'�M�����,Yh�-��T�����}|��y�x-O�(c�A�=�]�C��M�u��w,2��Wօ�J_Os}��o���&,Xt ��.�{l�'��Ft`���hGϡ�g��D�JOe$�CW�79���%�˧���:����?+/{w7���(ɝ��V7G;3Mv��[���O�w~ȯ�_��<ʦl�p���cė��*S�
�[�o4`Y�+�	4K���=��(h�{.��<Jh��&e���+8��I�qkkҺe'XĲ.�7E1�Q��W8�ezYq�f�e���٬��;\�;��{�G��m����71� B�)�يN�g:�=�¡�+�dYZ!���sa7W�ѫ+:��pT�9`�,��!,���n�i;��eWCе���[��{rZ����T���$�:2ʬa��<���w�Z��4ف��O-P���'(]�Ta�Z��3k8뵲�x�wofu�Y�=�e�; �ip�; 8!��Xa��z�@{xk�|�in����S����*�?��~�s�1{=0vw�߇m��a�#��`�
i"�y�׎�\�������^�v��/fy�eO�9O��G1ʆb@1a��p�C���X^}�;�g�+��W|������?)��r�n�f�ҋ��1�!����/> �P�ѓ��k�r^r#�L&��Uݪ.N�U�/��*)Ns���s'�h9�f�0��y���- �'�|_E����7��p�F�q#�H?�	��*�����
��M*��&g!VT��f��Σ� �Z(ޮL���Ե״���F$�h!��@��֎ծ�9L:��^+�c[,S�?�_��� w�g�>�u��䯲`[zL���{-�ZS�	W�ҿ�߽'�Ӟ/Y�����N���M��e���4go]�༳L�^;:é,����n�Ň,�p��{��ʹA�2^h�ߔQv�ةY��×1�Nv�φm ��vwC6<RZ��/��oo}�?R|������>?�G�I]�	��Đ�
�u+ς��	mT�lni��BqH:��zDD�f��[ؼT�ɖ(����XW�E��M<Rh�EH����[B���[aVv��[�����By��N(r�d^�Ja�GF�4�pf��4ǋɢy>�N�u�����݋ʵ���Jvc���!�%��)�|����ƁF�[X���{[O��F��ݬ�:�C�<�3[L.�m���ư�0SfT��J�r��� ^E*i{ve�,��]Urh|ýܵ���:`������<t.k�X��g�N�q�Y����v��z��ɂ(Όl6z�5n���}E�<��t�	����-��a���ф:���e�^+dɭ-0���i(��|���}��A��߷=�I�4H���b�C09��n9����z����fQ��Q^=��iKv��?�|3��~sgM�UңP�C�;��n䅒�x|��\z#��.��¨��	N�tԧ���4�ձS\�^s�L0\}�Ȱ�������p�A�˞� 3ƃlW����x.�^yՙ���*V%��O�"综j���5����NȦO�h��)����#&�lG?��wf���k["�@u����5>��;��΅t��펱�T:}��B�(L;��X���ձ&+��}����ݳkg(�����Μ �a�����254�j�h��^�9��F���8����j�H��u��M�]��ޛ��$c<1i�-g�N���ۋn�
ɝ�j
�S�=��-�>@�|t�:�*�����U"u�8c�]��\L��X����������EEz���a��ۙ}��Nfwrf�5L��%8�7n������A[��	^��?L$ʖ�|9����f�W���ku׉���A���&��Hj(γ��2�Ο��� �`d��h2�~���3v����ס�zaQ7 ���e�B}e�	�� K ��j�o�yQp�4úP�-���$ٖ�TÁlF�*H�V�T��N�{ �_��tB�B��UO�v�MwFP�>�e$>��|Le�/��i���Uղ�i�,�R��f� _Jb��'�)�x��R\О�CoDCF	�K���.�y��nو�s���˨T��7�h��S^��B�|i��m�:v����>���L��}v����ݏ7��?*
/�x�[��:�JW�>ݘ�]��M���ۦ��}.�vnލ��;؅C�w��T��,����B�����ǖ����Ǧ��@G��Z���
���g�-'��~k�E[��Qc9�*��"��+�pf�Ӿ[�	H!Â�-��,CF������u��꼋��Z:��v��w��!}R��(�E��(c8����m�61�����g7K@���eV�ڵT�6S��Q~�R$��a+ӯ�SD��i}孻�p��Q,�)%�0znk%nY�z\� ��D@L��y��Mгnd㋱�Qa^�y�إZ���kl��/�X�Z3�빺�֭p�\0g�����Y�tǧ�smg�B���JװT��`_�.����y��ì������v��]bKV=�s#�0q�<��lsL���-��,9�
T�E�K*]�_"�#�1K�������;�Z���lm�#M��\k�%�P(X\��95n_�gŋ�S���p}ĩ�9&���Us
*$�P�.ݏC��1��ǜS9~\��Pwil׹�2�Q�.����{_=T:��;Ǵp2	��{��8�
[�by)� ������{%�V>&:.:%��fW/X2��G�.���8�=�@���W7o��E2�Lps����vRϵ��.�3�;��5�{�'���v���~�%<�wg
��2�����CR]�3V9jsٴ�^� ����#�����|�~$z�!�����5u�OП?M�0�O�~�q��@����{k��kM�[��/�d�)�pk�o��]�p��I0�Z5u�FB�ʞ�����z��H;�8S/��&���[�)���A��B�R�j��VV�d�y�&�{�o8tzm�%G��й��#� "p:ޛ�C��*z��O�Y��.�ч�H�ɻ�}V�³`Fg�&F�Ř�SCK�ҜI|������x/3���&�ֈ{�����C!	,��Nm)LR��]�o4b��\e��CW��E�(�����PX۝�(H.��'187�fU���,��n�bQ�ß���]D'��o]�<����^�_Z�K�{�n�ϻ��0!��K�/�XG��>����V���7��j�5ת�j���5��c�=�z��mi�su	��{У�S����]i�?7���=�L��[���F�g��%w q�/o��m����ޓ6��a9BaWt�I�U٦6�&�^��E��1Ԇ6�A�$`C�k�`�_�vi�X���ʼ��̆���7��u�;i�ܐ�pJ��ڗrMG�=��cq��=����)j�A厭�]iT�^L�۩��E$w�� ���z�:��\��\?E�wQ0'9n;O�a�Oݹޔ����K���]{�IV��.^\����[:D�osÀ����ݽ���鰾��QH�۱W�յ}��c��:���/~��]3]{�8�0c�+B�%��5>Ĺg}3�n���=��]����l��LK%�k9yI��|h�ܻ6�Ŷ�lA�Zڸ��o�9YXՉ �nQ�}3�_���8�Ncj��03Y��j�8�
[ ��Q�nC�^�1&�?n�wD>��ȸ�D���;�!(Q{j���4�L+� �}]�[��>���UuNu��OP��)̘d�Y�9���
Q?�V�3ӀVE���ݨ�������n�!e��[�zF$4w fw�oN���~�xή?T�zx5���9�p��#��>m-4�}��:��0�s�JYW��Vtn_qaH\���R�4��@��ɷ����+�63>N`�3͇0�a���.
�&�l�]�r�h�W��|��j�U����"��a}�����r���h�߄>�W���&u�#c�Q�D���:�U'�T�����	�o�e�>0��`:v�wVV�|f�ȜV���N��d�$j%3��Z�b���R�Z�[�3���[�+Q��͇p8��ق:t!C[�z��bW)�N�
�qf��n�1���� ~'=zn=bF5��Ǿ�o�#ΦS��ȣ�{n���}�p��!��΀�'s����@���<
�q<+��_<�#u�z/2vE;t�/ݽ�o�|��w��n�>�5�ՎB��KC��g����}��%�d�.�\�u�0�qM��6��R7C1�a�9ߵ��`�Zr�/{揺iE�|������VO<�+L��v?I�K�ƚ9�������k�ַ�h�DjP�x��RMxAT���)b�uD���a��X�Z�b�k3���;/'D���E��3ת�y�\��]շ&:N��&�^��Kd�����h3�9�&�n�e�|_f�=@c��`�vAw��3�W�F�tԬ���S�F�nX���4;P(��Tk��9kh��$���eN�[�.o��y ���I<��<�]�X//�<$���yF�7�ow������Oʶx�	Q�x�����vY�B�y���6�Q]~�UH�Wԋ�,q�u��'�Ѩ{3��{*�[�3��A�No�K%b�&���ݎ��7}7y�c��3�iZ��p]���ߵ%�ծ^ݒ����c��VE�M����f�%}<=7����`�Q�m)�m�o�95����̒���F�f`��s�o�>z��ҁ��)Y
�i��Z�Q�F���ޱ�é����
�����!mvdړEv���bXDmwD�"��՛��{�AM���B��:J��Aer�hᓦ�5��emM<]�޳^a��b��y>SO�)�o��[�CEh����\���b����2a]���w���]C�x�d���{2<$���!���+���y�u�b{o|�r�E����t���%q����Ndn8!��.�׌ё5�-��F'3jG�*�h�
2�P�q�κG��������C�ْ���v݌9�ݡm�kХ*�S�|�Y\�tq�� %��Z�׽j/Q�̓��v[Ha���K��r"Q�9��\��{}]�}����^_V�}�������>�C��r`��y��	���q��V�e� {=��W����{���o������|�������:� ����0׋c�T�r�:��>��yt\��_>5y�vw��KBn���#��[i��"�z:�k����MG���"���f��<�p�>��7.G3�6��w��I�0��|Pۻ��E{=��9=�v���]�n�}-�a}�q𶨽u-�%S�'�ǃ���.K}��绻�'���^�xy�W+qɝ8�6��T�_=�{�F�G�*P�Y��j��-)�{��%�\��"<Oj�Z�����;{�皠{sL�6.�IG�/��>���a9y���S�^�/x��<z����~<�������ʪ��p}%�M�/	�ӻ�贡�wm�LJ���<_�NQV���;���(���k%���C����.�n=����p�>����e~ƉĺW��oNx�O5ޞJF<�滖�$]�WD��G�'�O�~٦l[ry�2�p���'��:�X���9 ����ݙ����xe���Z}�맶��OL���`��s���t�k�Ν�ݠ�x,+@��Al�Ě�y��:^�ս͒���/a]�@��&�o��A8O#;k{]�b�=����J{�׌��Z<s}�q�]�V-={�|n?*���[8ðH�O< {�%/Q7#V�v�/f�d��:��EGt�#՛�l� �ڜ(�k�'�%,���0
�Ykp�ٻ�0���}Y����Q�۷Svd��C�2�QMY�W��=�g^��E��qM��x���{̯�.<�zd��{�&;;U���>�Q�-Ӟ }x� `8��_=�׳ۗ^ۭב�;] o�]��E����Y�%#37��Ѡ�ЎVpfq�j�1aT{J�,mҹ��]{K?�`�ޓ`m��s�q�1C����9���F���߶��`��o��K9�y�!��c�%y�)�]�����>������f��Ȧ�	�$�&�7WM�u��D������NE��=���u�4�*Wy<�y �����~!�t۳5eIf�� �Į�s���*W�\
c\kEE7:����%}i;���V�j>���z�ԡ�*�5�t��H�7����`'�|;�.5��,�f�t[(79�3��=y�+;�3�}�tr�چ�;}����D�þj'���0\�S��]�G,����
̜�c���+X8��b�vi����g�F`��"��iX���vT�o"юQ陇�5V��q��5+��f���ܝ0��Wr�u��G����\X�Lizg�ʟ�U�B���g����%>��o����������~���x��2����Z}0�ے��n���<��K��r��k��^M�b�c�q�(A��"i�>V�۽�t�/cB���i������Ft�[�%�%o#�ߺ���kkS��.�T��o9*�%C��&�y眯ȸ,.v� ��/65��%͋��\�Ɇ��j���=�C��۷��ǽÔB���g�| !�$�I�Aci4$�&$h�� $���4�2$I�I��M7w�M�ݮEG㦙iKFƀ�,��q\�].b�X̋����rI4�41(1��RR\�$#�4C1cs]�r�"lE�9U�I�E���N���S&�i�6LlIA���%H�Q�dח4RDX*6{�C'u����,FCF�K��X�+��r72.�Ac�8��ܹ��,U�(��5��X�-9�ܱ�ۦ ���%s\4�7]�*
4A����;�"w\��r�
(��p;����o�oY���l�0={)���ܕf�I&��	P`Ɏ��Ղ�Lj�;O?`�r)x�W�g�q��)��=[:��|�y�u�{�����}PU������1�e�zO	;w��$Y�_j�D|��}W=�Uz^��澪���ڵ1��hv��q_�n�؞�F��������[� }=ީ�{2EC/`�L}�Sv��"����]�O^��h�/S�X�{y��4�'�$'�4��7E9u=s�뼞ޓ�o��S/�Cݞx���n��DH�#����MW�B�����k�E�edotJ�1O�K8�v����עnz��\�Eu��&e�5����簾���$�&���L|w��ݸtǤ-@X���K&����Ԣ��S�19Mx�����~�����S�pA�Y$eBB���
.�h��/�F��wDy�0�K��	W<.�JT���SG>���� q~�L_�?t!1�>sv(��#��F��iS�RV�*�l��Ñ�`���2��+c���M��%� k��Q4y̼wx	˾:k���畨_֭Dr�?{�^�] t��V����Kc^�]b��2��K+=����y�{H��P��Z�Q��{b����#��v>�{Ӥ�7/�q�\�)�����:���E={ed$h�p��yd:�)�����"���󷹦�Ǹ��9���Q^"(�����T��������f�ܛ)�h�yh���Â�Q�B
�̿�CLb�]���!�փ	��h����,�حڎr����e�3�{�Ÿ��zM���x�$��ޠ�y�ޱ:�M*��YJ�\���Ɏ/��#�hz�D�\���;\q��0���6#��5�nX&w*s���B)��Z�4��1ٰ4���c���{�WT��Ł��,����{��EN�*~R�ɭw��}��Ͻ+�w�����������Gƾc2n`�{H���j�{���(C<=z�Xǯ-F�F�b n��m�i�MD��}�{�ϲ�)QO�� `ԸN���Y5"����E?E�>gs�-n�6>_O{/A��Fq���a���l'8��^�j18�q�xe&"�k{z��j�R�T��D�r�o�C��^+�ך>71�%՜Ns�O6��I���0���)��R���X�P��39��5�vK������Ȃ�\����i�<��I��{^G�t�Zc|H�-[��56��E�h#�z���d�6�oP��n��_G~%�8��C��,�F�:ӛJE�:��{�XGP�$��Lk�+Z�ӛ����	����!mr� �)2h�{�_��/{=���O�t�� d������oӫ}��BnκP�*K ��Sƫϵrۉ��R��Uڰ�?{�de}3��;ͯ\-�\�|L��F���Tqq���t}���_Bgrԟ�������]�p��6Do|
Ӊ�L��)���;�� J�d��A{��f?��>����q�W���^NC�:�|��1g��,��ĔP�K=� NL�/�ɟn6&��Z:/ɻZjҚ���~��S�J����	z���U{�;��d�m�TV��s�U�^{ᙟbқ��tI0��I5��F���Җе�QRR�{L5�4�[��|u}��N�7�-!Ad��n��+C���Y˺s�$�G��þ7���wN��'�%�W)�9w��w�7;�y��wxq<\�`c��弒����܈��K�x=��wI�����g�L�/���_��|��O�ֱ�-��{tJpN�ϥ�������|�ҾI�j�����}D��x�j�r���{L�΅��g �b�YA�� Y�B0��e��}�e��N���ķ�6ڤE��^o�VF�����q����uf�u+\�w�j�|6w��$T���9WIs��ltS�v@�h�gIKƹ0�:�꾍ۊ�#�^Y��t�!!��/�M9=s�(���)o��b�ĸ�~U�tZA�#B&�����ҁ�AO��&A]7��պ���^�.0�i��\���QvD��)�5鵄�٧�t�O~�z�q/W��~��1}�tW�-c⫊v��޹=4�"���&�����F�J��|������\�\u�R70�{4(�DE�Ko$tә�g@
�d����Z�CE��λ{~\�����c��O�<o;I%j��)ܟ\*Y!���t�Lis���3p�ś��Wfi/a1�v8��?��`�&J�-���̌�@����gϷ坨��D�Ӊ�gơ�ccO(X)M9��9=�V��o6糬��iǋ��9#;�@/."��h�5;9�����
�٬�vBR�J��#��ʔ�\<��9}{�F�;��%�C69e�g���N�b����k*oh������ڿZ=�4ﶦ�Q YR�YMF�h�|�g��c����t�b��w������8I\��J}�aqS۔�W��y�H���y�������p�\�+s��sdݒ��P���ɣ�=��U��)�s�E�#)����0�"��޶3��j��oC	t�v��q�U	^�<X�:�м����������ϩ��.?=�c��x���-�O��5Z�ְI����{���E��.����ѳ��f����ҽj�񓛯��7�� z��>G͒���ؙ�l�V�T"}Ÿ�� v	��N�#)b9:Yw�GJ}��ϗ6-x���9��W������h$�$���1�ﻬO��+���=<.~�k/��lO�0����־���"'��z��6��<��|{{��E��P��у�S��^�8w f_�:�Jv�z��؞FU�L�(yU����nqa�_+d2�A�2q�G[�(��ss�^�re3WQ��i6���,|���Zq>�������xcLR�������7'�Js{��R!2C�G��9ʢG��K�?�r�|y�um^>ָ�e4�R�ݽb;�^���o�Yq^������N�1C��E|=5��u�؎D����s�N�q0��{��r�kV���a������y%ab�JN���9V�7%a]�d,
�DN�Z-ϛ���bB@�zG9
uB���:�W m2��cz�rgZ-�E5��i��΍`���|�Ur�+x��)+���8�U�.��}U�҄�(���`��❗��5z����羌Us�d!@��:	Z*E_<�����a��v&oQ57y�S��a�\75�}���d�����듅6�+\�U]/{��o.�X��^f�P	���/���u�_G�-k���*���0kd��\��a��$�� |�((���d�o*�~����*KS.���#��L�G+N�LGJý�]U\cd��ZR�=�ҟ�`^J}���/����й�y;��Ί��ʑ	�H�4�9Z;iQg�t���c������cH凊u�0/p��E�w3lߊ�m�����k�߻�H�Hw�q�֙We�L%t���w`�q���Ͽ# �t��{IH��	u����b����� ��1�O'��0�u�[�Ź��C�ϼ�]=͒7���ˤ�)Cyr�1c�N�Z��]��ܡ�Վp�&���(^ zy�7S����=�zMq�?eq��<���\d.�b+��#.;��I��g�v~�`E�Y�����0�z���B_o�|�A��˛�:#$����qI��O�wtl(x��8�ҭ����ǠD#�%'�^�k��E�Uұ�Nr}x:PBf�[{Y�U����u�[�����	�B9��4Q�͕��l�����ҔF�F�͙})�����g*U*²w�X���Ա�{u�7&�^�N�鰙Eڗ*�8�?e���!\��N����U�w���w��ja��m��B��f4�9��*��V�:At*@�EU��|���}�3}%�r������1d�*E��i���9n�d.Plழr������w}�;�ߢMC�<�T��
��F}bO���W�4x�<l=��,����c��=�
�Y�Q�sC�9�!x��r���ڍ�i���y/)��_eC�Q��t���3Y�?>�*��-s��<�G}1�A���`�\G�{	����TU#�/&�����s^Lh.U5���r����+7�k4��d�yqMsu��:�;o���G�TW��4=������M����տ:��;K��'Oy�X�U�HEJ5
�_(�\�l?��b��q�E,�i1��kdv-H�ˆ⮷Mlk����q������G*4��PR�Kw��%G�H�U�����������tkq��z�)C�ݓziS������T�@/V��9Ǚ��X��Z��'$���A�;���C�"��|P��l���g�Dw���2�uݽ�Yn�J:Nѐ:����h�q�8궽�'��c�ޡP�7�/ә�^~}�4Ɖ�T�q烢��1����`�CӰ�w���e��
n�Cu�
�J>��q��Ҷ;��<��N���#�j���s������:�9Cݢ�77�f-�u k�S��J~��l<�aZ���KX��X�9w��wUB&��\�1r�-�vdړ��F���'��YA�y��C����e&�;D����߀[aW���V:�����⥑g��V�8�[��a�����I�`g ��$��ۻ;Q�Z�fm���f�ʒ�T������Uz�_�]5r>�]����n�c�}��G\K�˻}��x���ed���$N������W�j*�vg�~ex~]�鞯��ߏ���~O�ɻ�?�9=;^��T�O�M<4΁�PD[BB(9]�����3����\8��1'�}�V^).�1ƚ�mӮ��p$,��.~ff�/MS��g��c�y��mMSI7ΑV�$�:gg�T�2��~*(�i��P�l�����nc��U5�=,�T��65ѕ��v8�`�n���I�rn��록_|�>�;g��á�OY\��T��R�ͭ6�ݢ�pX�1!�f�;���6CvV��)�xz�N}>+�b��/��r@��~	�kB�=o8��a�`G�\��W�5���-O��O�'�v���+�e�J�+����n����o@q�|y��}݄W-�*� ��q��^��#^eӔ5E�>��ɠ�O��&K����V��y�j���o0�,��2�#!�3x��X5+b��[��U�^
PV$��%%��NЫߎM`��턔�g7/l��g��=�U��3<n����1}�+�:�����Ӻ=T�����Q��3�iOެ�K��j�~en�0@�N�׋�%�յ�V�48�Y�����OH�no���٘O�"�r6���W���Q^�%^Y�I"|Hr��R��!���uMe��{�J��<��
#�YjJ�j�����V�>�p}�:�+�S���<�Q�"&��p��M2=�{�=TF�v@Oz��<"��m����FJ�$�s�����vg�v4�R��7�)�A~�f���ąj_7Ork:73��1 ��JJ��*������ʷ�������xsm2M�a�r[�����ܵ�DE,"E��dP��c�x��%U>���"�ټ�˟��=�;��r�t'^�2}�Ep"+x��)"Ί���<S�ά;���躚;3��k|�\b0B9�kӼ��TSXΒW)ED��پ��z��i�6�����͐v�&�M��(����V�������{�}��g����{=��g����w�s]�d⤑��fZb�eX�0_���R�������7{i�t9�/jw*\�Wb{,@��:c�=ܒ�����	��+}8��i���V!�_Orɝ�-���r������}���2+b�kw����fӾΊ�'�}����w3�n矷���u�^���S��w��aǡ�`��մ�܋K����l|)�ʭ�z1˹����F����}���x�-Bk��4��X�^Go>���10�;��r6��P쟍b ~�7�\زɾWc&o	/�h��Կ>��Qؔ�R�ln���)��{��f�H��;268���;i�\^�s}��у���=>Z3JS�P{��9I��J~�hYK� >�t���k��ݳ�+���Զ��x�ݗ�u	��!��]z��&3p{$����'xo-re���v[�2},=����U	L���n:Aq)�:�<���fS��7'ZT���\[�c}�O��<�~���wn����V�A�J�:|rE5�7fh�B��8��<���������)�T�s[ZZ~���7�.�Ӓ�>:��[��:��WڸV��8΢e];^'=�|�߼T���<���Pzǻ�o�j���.�ϣ{ђȏu�jz��m�ژ���w��y��f�>�vg�n�bW-Ş��a��q���=M� �8e�S��H�£d��f���;�[�����t{�L�y����6���}��������qyF#X��{ï=��V����Yχ?��o���a�A�G B�P�5jZ��ʾ�&Ep�ZM��wb�%���Ѣ媍�2���z'�ķ&��
�j�C0ݧf���"��U���o�O�;�n�/,Y��u�,r�hf
���&��-]��ޔ�z2{e��j>�:
Dè���t��6��l�\����v�Ӵ�h��9��9��nWJX|q��M^de��)�g�[޼�Q	&����T
 �B�v�ݯ�?s�F���>x�v�W��A���c�Ml��Aӹ��l9��ߝ�L~�A���x/oojWu��8*�F���Cά]�v���}w�=ڽ�"�xa�Z�v�òc��ˏ��rd�t,d�;SҺtzq�p$祧	�P���U��C��w��D�#�2WN�(�So7��/cB��N���>W��`˝j8��M��V4*���c�ZT�;� Lv�Z ���͌p�C'��q/�>�h��� ��g��BU�b�=��X�'Ł{��T!>"���#y��t�H'%�;:7�0?e(�,�Y���^�^;�!�'_��ǖ�|���{E�f����7Ȍg�M���,/��]Y!-5a\��c�Jяy��;�1@s^�,��6�[���6�
�s{ρ�y@)����r�;OSc��}�;�^"D�ר�
�J��S^а`T�������㬪�W峹A�7;R�[�1�y�V����e*>c�hf
��U���h�t��G�����`��W�n���w.�ɷ7-��wwv�9�#��d%��Er
f���4_��<�� @\�g��w[�Mc�������u�v+���v�4������P�9r���2d:nQsNn9����sD%���]uι��r�vwq���+��"���4�vu�a78�\�]w#r�li�����b(�QpɺN�n�5��3�]����,]3���ۛ;��t������8\�cwt��t�wqTS�
�M���]�bNιӄ\��]Λ����t���\����n��tM;�.�.��nj-�ҧ9w\�I �����%�$�Ʋ�&���	��
(�_޻�g�cݾ�Y<���b���tp����ek��s�� ��BJ���5�3s��Ǐf�]��E�S�}� t���� �pX�XR	����,`�v�ǽF{y�O�][��pI�3�^��_S���|��T��Y�<�'c;:t>Q�kM�'�z�s���q��^Cz~�2�f�x��[�z��ͨ�&��n�Y�-�Q5�Nfϱz��}G*����jp��!,��/+ ���<���ە�I���7ZT�q��v�Q)���ݙꆙ;���p1i4�	��M�o�1�H�/���z����z����$hD���T�!��T��C0W)Z��;�#o
�F�U���ae�;�O�ý��Fz�EZ��#ȫ�>ا��3������d���j��W3sF��6ߊ����A������͠p|}j�hF%Å�1lb*bGA���՚ͬᢣLJ��1��Bz��mi�ȋ���e}�U�h��o�B����xik��
�����-�H%o��;��^�Ľ�W��\�g:��-�<�)��AѺ"{�m�XWGޝ}�Щ� yam]6����J����������ʏ8 �c�wb{=���[���k��3�7�
ٚ`s(rj��5���9`!�,K����>xǋ�v/���}�$��B�u��4N�X��y:]_ʡ�"ȄDwj��κr���)Q�](�<3�'~S-%"����e}ߕ��j���Iȩ������$rj�i~���ףZ\�u��8�:�*|)����H^t�>pU��-ٽ�vzT����sw�r;��5�1�\z��ُ���!p���H���\O��O���ꞓ}�Ѣ�%�rM�,���T����Yɘ�"F�MC�l��Wû6��e�S����&��_)��E#Wt�����]�a��n�w��헳������<����I�4��V��Էz(IW���w��36�>��C>L�ϯ�7��ȿvd^��&0��f���L�]�R5�ҥ�� ��:�txv���� �<��ףYl���گ���ɸRR�����_���)�j�ۍd��LE�b,yFO�ٽ��PZ!�OԟӵP4,��eb;w�:\�I~��	+O���w���,�:ygf�p��0�On�<l]��h&�
��ё���s4H��>	��f!$��WB��[X�,�U��3LL�򦺚�ݶ����ẁt�Wm�����v�T�P��]��DǏ���5�i����#�<��������&��_����Y7ş:՚�~��W��VDO����kǹe�踂�b�<�QY�DZ����zSݮ�}dǛÕQQ�H�@�Da\:�Z.���rct���A�ń�����D�쇫\��^�_�)�+E���yu.���(��ꊉu# ��Af�!e����!K��z��b� ?')�Q�����s�;�4�4΁��]�B@��m�{��S��w�ù s��gG�I�8�#r�O_��B�v	�)�G<����5�[��n�^h��P��c�"��L��|�;>j�.���E�u�gfn�������ǍƑ���Me*���ポ)��ز:eך��g���³n�v��a.B8�.��٠'��*�?Lw�������-P���7S�;����珗*7�+���}�ۙr�rǻ~<����BQ�s��U��wK~2�q�=]��[�t�[����N�e���?)��=�w��(�-5���)�7ݵ�=Y���c�Z����6{��P�:���5p��>��t簰Ot")Gz	#߼�}���dV�k���n[[�%T3g��قGs�����m2��{�[��u�����#zk�s���̚��s#�B����qg햠��z?)�;�w�~}O����������\�����z5n�Sٙ�B��ǧ�^�˦�ڢ�z}:�gV�Ma�y
ӂ-0wv�G���tT�ҏ�Y�5Z�<);{������T���OlU�� W}�ъ3�d�A+V���|,Ш�f�]�67��,�{I"BI��a`���5V��s;{���W W1�K����>��{�TW�Z��ٜZ�9��%��tM��Rt Y��O��PP���c��̾�N�:�u�]Ɲ���^�i��/�}>W��g�mq&�_��:�;f�\��v�UWY��g7T���W�$|�J��+m�D<q���(����1�!r]���6a�8Y�28u��8�<����_�^��gCzg~�<��-�ah��ò�i��Ax�r�W��4��h�?bEG�[�r��R˝�L����X9��,ۯp*��߃��_93�G)��{@��N��;����K=�����o���{.��ŀ$OR�F�]�e���AN�]@��)*�f����na��c��5���l�R	p�d�W"��锕��ij�����FMʣӚ�23	�H�B����2�V��"�Pѝ$�Ʃ�����)fg��ߞs��N�����Wߥ|��O��J7<����=�G��=�?{'��uIN	]/�x:�a} 0[�j`���"���&l�1f��={�sϲ�ʡ��Y��wM�2»��Y�Щ�nw.��n�ދH8ų
Q��M�'���D�P�F�e�t�w��͐��
�ه[��fA���"5�&��ל�����r�2vo�G�G�	��C��ϵ2�B0�e�g��}��z����"��7˱Uu���k���,���� `F��n%����u�!�[i�o���ړ~	���C{qR;���z�4]s�m�=C�g������c��݋��xa@���LӑsNs�/�*^��+G��%�9�KX�0LNŸ�]:iX����H���Y����N�|$�m��'V���Q�ӏnsL���:P`�$�
s ��>߿R�u �<{^;ا�v� �WW��W����z� �$kkDI��[�O���؄�%��X��sU,��Gv���<a��v����3��i*M������ׇ��L}�_�-Ps���L��'��g������MX�d�Ϸ�[CܐJ߳�����׹���}ͳg�����|*��Ю���������'���]�7t�������˻��/��k�h.���C��ף�_#��4����{�Od�8���8�4QT�6:�ԍ/�%��q1׆2�'�73B�FU�E`\�B�)X�\hy�:��=f|ُ���!z��k%������D��;Sb���f�^�0�W*\�>��|��S�r��m��}k�9���R��+���tl��S�/��rך)�Wt���P���Q����U5dQ/q��Nvt�B��V�N���\r�If��n�� ���o�<��pt[:���-��O���=6�Pu��ꋙ��Ne�2T�b�s�����	 <��;��#9Q���s��*��Y=��`5o��{�ur�c75�	��76T�<���e�m:_�u�y��}�]h׃�u�.��Ck��Mq��C�}�|����.�߾K��}N0H�u��^rWZޘhG���U��n�{h�U�A� u����]����o{}B�K����u&�����P��G���=!��3�G3��0�5?|~��a���G`�=���ӗ6��=����z��؍q�ڽI��Z��	mi.��z.p�ھW����"F��BDA�x喎�nD+����hW�-��r`m���6 �M>�Gbo*�Nςԁ�G�4
�+NP��jr�V�bw�`Ɋ<�Ԏ���%�U<�g�&.|�&�e�=���o��-��z&(z�������!Nu�ZǇJB�W����i�p�c���g�Vo�N#r����{�}�ۚ����r�;��I�������tpM��9�3&.����1����$��E�U\2�h }��B���{T�C~�Y���7ၯ�z/
��U�����z s0�d�r���k��er#p':�5����#��|�G�{��x{ڀy5���E�!�&�����iuX��@�<��w+���������
P^)"��^�HܷSْ��>�w1GfV-�p��~�Eq�tN��"�A�Wm�m掊~��ΚF<m�
	yWO~���:t��}�������a,��\o]���7}��uoc�\qa�K�K$?�#��1��UB���U�Nwk6��qmU���}����G4��T0q����`��"5T��g�~��h�]���?X	���NF�35��^����+w}K/����0NmU�˯}���xg����i���N�[[���:M*u�#V���(��6�����p-�vH�y3Q��ᬳCE�0�cvaF��]�3����ɠ�H7`�	=̅֝���t��<+�ƟpנV�5�2D���ߧ� ns�&v��{���Hhw�պ���`<*5gX%�X�ڍK�����wh�,*;6�F,��7E�(:�\og��r�{�Q�pE<r3S�"��� �ӷHL�|2����ĒV-zk&��îw]A�"G���qY]��:�7o_������Ԕ�΃����8��G%�}*.ۏ�}�`�{����rA� [N;�7����o����bY1{m�§��<Ys�8ǆ��c���}- ]ݥg�8��Ҕ�]ٗ����ۄdI�M"��O�g;���'���9;������#֤�����\u���E�)�3���*�dÁ3P躷�;���8�PD���ё��!^�F|lɣ=��s�sW����0e=�YSk��[}��P��v�ˤs��T)�$�����U�_�F=U�i����B��M3�W��t���8���~�wђ}^��2<3�|d����O�������. tWP� ��}yt,.Η���Iy�<�P���{��������@b�)�@�n7���d����_�YZd���x.^�s�|?OI�2?{�|���?)�]�K�PKR��W��V)�=Pi*�s>�\�G���=���`FS7���ԝ�)��7��S����Ck�F��x�T����5�[�������:����5��������Oj��{uoڗD��}�b����*�r�+�^�jU� \={�J�$�H=�e�ӝN�o$g�SF�o��}+��e���+h��N�l�v��
�%����B:L�u�����᣾��뮺6V��^�˚7��ķe���������G�&j��m��J���݆�J��JU9ݹFT��w����q3�@܆�����h>ٟF2������3�400n��}��ޏ�>����E�ծ���xVs�;�gvS��)�Ya�
5�y�I��O�oW�����nC���zLx�1�}p�k'Ӊ�~��6�E�ZO��_e>��R{�,BQ/��;�!��Ob����j����{+Ga����z%J�{\�]hI�����L}��t!0kDo?�B�����b|�D��w*���}���䂚��l�g�g���	n���?��uC���s�.�/kdk�UX��|��h��6�ɻ��55��ӻ��ϐ�x�NE�+U�����O�������{?/����{�����N('�խ����/���v{7���/t'�Dzn1
c�)P�h��lYi�Z�����֟�����e�5y��z��(W�gn"޵���w�?<����)zi�e�X1-���y$_�����<�rY7�J/��ՍfM����T�q���<u�K.!]�{�T��Nj��97��&��<$��]���O�J����m%�V���кo�;��
%���I�0�_.y�\�5e�{��7�L՛�=�=� j�R7���[�[:�N�H�T7;���jҗ�]�lI�7u0$Ŧ�e9�����%:�w�E<����}=���郳�y���u;��ތ��CN�����p�{OAm'�\���J�
W��q�s�<��!�ZQ�
�ڤ�㦬17��A��Kwѵ\��5i��AX��,�r���{/���>��+�s{�\=�y�+�}Խ;;	��	\�]�&<A�0����bM�s���wB~�~۩�<��Oњ:�o������΃�Q�nN��？��{d�6���+V1�Pf/�@w#w'�:���)�.�EY@�I���`r��v��v��r^QP��VNc��A�/ޚ1�H�,�)^\D���f���V��%�CU�����7�77}�p��'i1����a~�@�e�	b�L���35�=�N�֛�E�S�9�����xN�X�q]$VY"u�t/^$�c%cF�̈�GtaR����7�e긇`JM���UX��8�b�k�C/�p�H�����T�?�F�>��ܗ���;�����pS�x���L%%+7Xӟ���=����Ǝ��2	>�ig�T^�E�B�7��>�'*k��u�y��o�#Ǧ��/�I�H�潋��=ϚUo�����*\b�q%v�M��J߀���5cW�������������)�'#ސ���7[=�Hep�/�g��_�y�lw��Z�B�7r���y��9Q�v7"�yA����>C|td�E['>e�]��8���������ȥ����.W���q��`ss3��<bK�B~'�LNݩ�f��!�ap�rmyyC��ء�wW����	!�YFZ�r�u�f�}�}�r޲�U�s���Βx`��H>����L�3oym2[�+��J�U�>��޵�7�[�0��(Ǡ��[,���!w���A��m��������@a��7tQ�Z�ڶ/�7����P��jol	��n��������]��t���������[���%�2��Ȓ/5ɨc%C3���F�{����Y����c�W�����t
H�C�L`}O���)���~bN�J�������Q[����GA=v�:���޺��kc�����œ��K��Ak�����f$B�=���Y���f����GYX/xƶF�~�0l煻��C(k�J��l�]J7c0��0��ݻ�+������s�w8���˘�;;�ۜR�EȨ����m˕��7.��ݻ�wn�r鐫��˧���\��ȝ�t���s�r��c��wd�W
wr+��Er��������Gw<���"�ۄF5Ø܇v�7.�4[���]����v��n�K�M˘��W79���ķNE��N��nw]wus���wrw].�wt��7w[�p��N��m�\��sr�˻������7u�gwr�ˉ���M$�ˤA ���˹��wm�u��.���äp������H��"�솽�=܈��A��\K��vt.l�듺�����F�۔�]�r�7Cu.sn]Ӱ�w7n��'9t�Gu�;��.srk�n�{���$��� �s��Α0� ��Do.i=ι�#%�ԅ9�4���]K��r��ھ��(���6�4��c�`����P۰�ٙ�c�k�P'�5�US�@��zB%���xr���uf'��q�n��a}0��[�^{��;\.��R+P�v<��$hK��d�@��)�M\���rM���n�M0�V��[��ŷ�'6=&��r5>�쎩��g��^h�b�]���Կd�-���mã;V:�`u������l�hל�����o~�r�'q�l�D���~��~�b���Cy�F��>�4��榡���^�����l�O������T�='�R����,8.�?b/L���)�/mG���&}�3ނ���S�~���zw�\ٷ��K?{�Q!�o�~B��J'G׈��Io7@o��c��6�y��E���&���O�h#k7JA�c��Sw�
"��xJC�Y7��ydF'��" �^�,�����y�չi��X1v����^��K.�78�)A��@��y�(��9\o�j_Z�t���b���9�7�R��������!_Vlq�C%�o~S��{> \"��_jm��_�����\��נ�{�s�fWi����Ƿ��������}D'���E�jj��j@�@�fM�=OY�n�hL�����_QJ��_�=Ә�� w/�§rQ��v�LΗ*-���")�������x׾���#{=�Yt,A^w""�=�P�TQ�rk#�s�Aԝ��6d�3�=e��{��i�={SdV{��)me�~�Ei�f�IqxF�EH1Ʃ��r�uVܛ�O;m9x�q�c�8Tz�B"�H8/���:<�69��U�B#3P����g��LP����uSY_W�o��ӿk�N0ħ��=FR��;�Y�7s�9��#:�Ě��5�M�ݼ���+g���\���.���5=B�*�.��gz-����z���[�=F�{�w�ϻ�ۨ�
�����[��
���!�D�f���h�i�(>WvONuI�'�]�!n��Lq����kz�z��-OCd�j�]�AV㓣_o��\���fdSQe/פ5{N��q��|6'��u�[���h�l#�AY ��:p��O{��x�����f/wo�,�w'��-��g�{<�s��8چ8��v�]�kߘ^W�Г�m�rNET�E��v��֫��%®+��ݦ_����<>����.zA�����As_��	�B��<;"c�&C��	@{cu��)e�a����}�/5����g3�#Wo��7{���c��AQ��K_Tc"�OUOl�O\;�o��v�G�|����r^�HbzJ�3����`<*4e�7����i}l
Sf�Ŧ"��x���ڐ@�Z8�`8*=�/��h��IH����p���Ϗ��מA��n������q�M"��S��=�A(c=<��3õ��w���Vg7b�H���z��\uUْ�o)Ne[��K;)�	�k�mU{���m�:��'!�VF��Z�XRrV��DYm�tF�fY����H�8�� ,��	��$_.�Ag�B���<�k�7�}ņTɑZO�J=X���m�M3�V���H�@��ޑ�M���������l,e�->�Z�ٵ��7uw�½J`�4=~5�or�ܸ�>'�v�.⡛7��*i]�y2�A�9��;J�A���K�с�-11�Z�=�tHL���'Y}�3��Z��k�J�\{3�-�g0q�T�5��P�������=^�Ç�Y�<��f�3�i{w=[^�o�~�����)�ɖ�쯏��Ng��˺qe'��$��>��<�|�mn�N���8A�e`�fp]VE�T�=7U}Ů�6�Mʡh���h�L���O���u�<�����Z3��{��b7Hz�W�=����}��x�E��g=q͐mt�a���̵e�tk�=�7�S���;�H���"�<Z�����QҤ?u����&��*�İ�WE��η�i���C�~��`�#��������|�����?d����:=��o(�/ ���u��^����`?Y��H�O�&}r}�-/;\��"����'_)�%�8�`:(���Їt{,�Δ��춽��su��;��Q,�Y���IX��x���S��xA�ML��'��_�9����ϝr���߷��Q���ǫ�b�xt���<��sw�ϻ��/�ˁ�Pˇ^pt���r1��(Q��#�e_c�m'�,Խ�
�(��:g41��ѥ�^���;8=�A�j�r�j�.������gw$iJ��Y�ݠ����<�zUOY�m����:�[�kl���w9�h׭7o{��y��@�� Ѽ���ݰ�p؊�j�ډ�z�/c$�Bz���F�G[6�Rz�զ����z��Z��W`����U�d>��!mH-x�����ywOԎ��}�-��-/�Ю<H�*��nxj�R��l5M�u�ʣ|�S6sxj^�N(�y%)GFx��V�j���S�*�]r�	������9&���*OxUP~�t�F�4��~D�������O�����}�Oܒ�\q�O����e�v���~���R6�w2���f�C��t
}C�_A�W&�+�QC�.W��5�soay����r﬉κ��ԅ�an[�ޑ+�ꞡ|��k袑��(H=
��ё&�{��X��}�����\l�Փ��Y���E񯴽����-��=:*J�R2@�`��f�G���
/ٓ���z�P.��Z��VnX�0,�o��Ё���mṲ䛗PdT�"�Wxz���f8��jD�S�(�7�͏KI4%t��u�mɹ�z2�䷜t׋����X���t�l�)���`��6��x���K�` �r�i�\�U�b��r��'c-�2-���������.wH;Cg�A��;�.Į������o�|�l��M��U����p;�m��:A�2:�J1k�	������z��X��5t"�~�n�f��^�:�N�9�<,�̷I��8�Q��Z����f����9����4���"$i<%"K�[晶��ƞ�<��Y�GE�MG)o{4�p�^3=���uW�g�Rc�9C*a�}���*��o��*�Ϋu#����@��]���F��V51[�Onoa�'h �6��+���@��3��ň:�[fND��畩�7�kn�z��N���	�ސlɣ:��^t�Ǧ��Jjm�~iU�/ݹ�yVtR@�a V�Zw5�Jˮ�{��f����J��1!{�暳��6���� W������q
o�\c�Љ�t���;���,`Aý�fnW<o9�aOo����)�+%�I>�V���ڼ^w��t���l��<�v���{EC�3���V���83|3�]����p�w�����Tz<3��N�x���}0��+u3�+�K�Y擝�)"���W�=��-�3�F�q(�0���N�3�K)˰�ʹ�@� ͓*���	���^�ꞔ�qZ˞-4B�<�uy�}^}:�Q�`��9���;g]eظJ��t�Y蘬��V�Qy�H�]������˯�����_��;�G���'	��������B�q�[���z�8��z��g���U���z,�n`�s��t�S���OH>=�ߟS�.oW}�z2��y��i~��Йąl5����8o���G��G���y�=g���F�]��9�Ra�@��>_\c%61��qњ���\�.�jt�֮���ش����S�΁p4YgT_*��o7B��v����k����H¼tW��$�ZB�P9���g�bc�IU�۴��Ԯ�=͐)!3�Z'�O=�T�oT>�xz�����L�o?
�~���<59�^%J��n���ނ��m�͔{r(�ԋgB����Kܝ�f�|z�z���x[�(�Ud�1�+{ѡz�DL�;���iþ��k�_�g S�>>n%�s�9���>y{�����;vļt�M_l��A��ǋ-ʽl��O.��vƑ>�����X:��+�%v5�G�yo��ֽZO� ?s>7
���SlXw`vè"WjY��������U쿏�P�:ؿ[�70��c�˿u�Wʭ����YQ>HH��$_.�΂�P����C�؞t|NiS^��U&~��U�����e��]�ɇJ@�V�'��=�/ �+�������䢊z�l�ϻ�������y��ڝ���<����iy��5}�8�a- �%r�V�r�u�k���m� ��KU18�6�WSf-Y�P���X���QD���0�[:�*�Ua���ތ�yp�(|�hF�ug��ȥ���k��kݤ��]�p̓�t�B�"��a���<�A�ǥiK(��E�r����/����|����>���{��R���^�?H�n-�d_T�r�XRsb��_[�v�R�%ֆ�5�]/�_��^7�<�85:,t�{<����xm����>�w^k^/��Iퟧ<K^���EN�v�j,���6̚��I��������{{��I�8k�j�B�����7��y�l�v�&im��gc��O�����ju[�/Frm����ucPo����_�N�|�ᘸ��tqn��>:(Ϻ�k2�0#���vm�u|��7�-Ia =�ނ��ryU��f���+�B5Ũ/�Ć��wp�}ܵ��v�Yѵ�]Qהs�����w�%�HD�UҜ�r���篶�4�ɍ`����Y�lBU#~���׼\��~�<>����ޯ�F⍲���93X����{e�����ɠ��2c\�|�\�[���3���~/T�n#�x.i̊*�P��<-v��g�[":��r6��}{��܎T9JT
R�)�r�F�u"���
b)��Ur���p����o3iĢ�"�h���z�Th���luө���7�R��wkit+�;�D�D$�.���2��9��vq��Y^�z!����ૃT{,
���v�l���U/Sh���Ñ�}Y�jl�+�*�k�:�Q �\�`wM��������lP�3�������zy����hW������#�c��hm"�b�K����|��l�����n,�7%]{������"�5$��/V?n�Vm'CF=�p��"7�_9�\��}fR��r�'۞�1������r*Nv�=�7%O�n���[NF�+���~3����sx�x���}!o3�O�Y��.ǀ]���C7˩��l��<�ܯQ�b/jO�h�'��=8y��IQ�R3e�y{ބ8�7ˌ7Lӈ��A-_/�Y��K��'�����I���N��)�AW'���o���Yx��?�3EI�s�[��l��=A����{�:@,{�
�ek2#t���ܿ���/L�R��g������[H�}%�Fka�os���y�V�]�|�-3�P��.o鷞!F�6ͣ�f���"t��oeE��F0�W�9��	�>�^VW�k���O���Ey����������Zl#G��&�I��@���Ns��9�꧇�����X�w�Z}*��k�z�����g��664�a�-͚m�4YVel�l�ٕ�6ٕ�6ٚٛYe�f�2�eTͶe�f�f�e�el�m����̭���m����̪�[,������[3m�[2�e�f�el��f�2�f�e�el�l�lͶf�Y[2�f�3m������̶��n�Y���Y�fZ̭�[���Y��+fU�k,��Vf��Y��+fj�ՙk3VYVe��Y��-fj̫2�e�ʲ�Y�ٕ�5fj̫3k3Vfտ}����m���j�f�m���m���fkUL֪���fj�L�����]�j��WmUL��L��3[Z�kZ�m�������L�U2�U��o_���vm�ٛUS-�ٛUS6�l�US5�ٛm�e����ڪ�m���m�-�ٕUL�m�6�lͶ�2�TͶ�7�z�m�UTͶ�2�m�j�eUS5��j�f�f�7+�fm�5�6ٛlͬ�lʩ�Y���y���j�[2�f�3[2�el�ٖ����f�elͶel�lͶe�elͪ��v=�m߆����E�J�e�R&Y>����O����o^���}�7~_����4u���?\��M4�>�{7r��pW��=_/���D�o X��z׉���z��+�?���H����9��nɃN�w�7�W��S��O#��3;��֫l�mmi[-��b�T�m�ɭ��kUMMUR�USKm�m6���m��m*���֪�Km�[6�l�ڪ���f�m�J���ɤ�K]&3E����>P�J̤�b����q{|��n�0���5.#ſˮ �����]6z��o����>��S�6:�}�\f�wX��������7䀪� ��㹋�<]���l�:-�̐[�.�\��k^�婛|=�gj�ۗU��j5 Ug8�www *���0n����|^��y����fO��{��H�w��G�U�;7�253'J����5t��{t=m�gè��s��i8�n Un��\89M!�5���[��8�Ԩ�pgz�a��n�*%Zg��ܸm�9�t���d�Me�%����f�A@��̟\����yQ֩B�	"�JT�����"
��J" *�D�B�I 
P�
+fU"�(BR�))%*�P���2�5�Y��*����fȘ�b�tvmU���Y���ebh֪����bKU��a�XىfQ�P�f��nغ��jZɖ*Zٷf�ًfm+{�t֖����6�,�&Dِ�m�V��i ��l��:�:[T��
�}5�Zb��m�$�����TQ$I+lڤ���)�Җ����Ŧ�1��k0[7�  �}��҆޷N�`9٫�$V���.�w,�ʶ�c@tg<�=�֕�r�za�覴�˳S��n��vM
ڢ�e��7��J�Z����{^��T�ٯs�e���؋QT6R�  �p�(}
(hzF���4(Q��|���}���A�#v
�Ç�B���}u���v�okm������F�ws��of�ܧ���W�iT���.�l4�v�3^Z{n�ӭ��Z�35Ueh��K�l�   =��{am]�7���CEme8{t����n���w]�uv�LqݧJ��ݕ�;�ˏTU*����ݞ�A�ڜ{�^��[g[koW�{޵E��7or��y��v�x�M�m������[,6�wnV�   ���T�ݴ�+��۩����׸[������v�k�i�ݳw-����T����ʽ�U�-�ZS��{�{:�ө� �	ov��wn ���M��$ղ*I33k.�|  oj����n �5�p�TMW��ѭ ���)UE��tR�j�1ZԵգGrX(�P�vے0�=u�1[amf֫+6ʙ�  [�4;[Tfu�YIW;uP
\�K��	{�E;J��J��sA�E�N�4�K[
�*��QN�M�M��5i�J�Y"���-��  ��=l��q�L;�T���}�W�<�[al�
3ڠ��YٸP �` )�3�۠:�{��֫%f�F�m6��۶�� ��/��[�� ����w�� �8 @<������ ����  ��  ��p �Pw�+6�X[k,��lY����� 7w�i� �f��P {=�  h�w4/`C������+���s��� Pr�� =.צ WA�\�� CΊ�l�m4-��Y�hM5� n�}:� q�p�T{�8 A���C�;�\��P��  �K۴�= 5̰t�s�k��n�^�  |���*P)�IJR�`  56�T��?J� �~%)P   �� �*   z����� '���������9[݅}n�������4��*�MW�}��G]��7�����<=�jiC��[j���U�����u�j��sZ�ղ�ڵ��=��klֶխ����km�����W�zW���^����~��[����ct��4E*��A�p�H�0@`��`/E��Nâ�G��f]DkF���:h�2Hf�Y��,-��F�V�,ZѶdBE�� �c)�&���.���u��fk�vlQq)�N�2�V�<Nc!jĒ4"�4�,,�H�ovś�'�(�����Z����2�9����A.إW��!�T�Feg��='1�m��{u�.�X�]M����J�l ����޺b�p&��[
�_�T�j�a9Y�ZU�+v����ӡWxfE,AV�!�iנ�̻Z�4����(��n���&El�{���_D-j�x��/#[yR�2`չ��Ӥ��٩X�Y���0�6�P�n��#K�t��3���R�^:ύ",Y���^�`[2B�V��i(�ދNR�k�pC�r�䖀s���V��l��i�[l�L-�)�'�؋S��;o���2f�6�k�Fo�'h�u�73� ��*H��݄�-Q#n�5K[���{B�^���ݬ9�ܫ��B��4��n�k뤑R���܍�R�Mvͫ�Jԥ�ٮa���rɛ.=m\�P��inMoN��2�[T]�{�p�H��YW�\�D�Leڔ�u��6�i�P�
Ho
N�6�
��-��5�,3p�e���miXp 4<�($�s�IM�/6�l1y�=`�6`B���]���V�cSi�SL�#���1a��&b��ba%�:�ɠ�34�e�PLtȉkJ�ɶ���f=��ӆ�Z�6l,�����]�5*����Jmi���ڊb���f��0䮺ib4���Ȳ��ۑhq�e�Yy�N�h2�['/q�w��/R�r1{ON�ci1ADI�eVk9��݈],�	�mm��S�]%$�4i׻�mL��xr�M�ڭ�l��k�AJ�n�&Bj��f�J �M+���+mT�\/ۂmD0� &�N��CX�kW�E
�j���n}��YW@HVCZ��`��2;є����ڔ�`�c�ϓ��ǅX#���ȩL��F�f;	�.�d&Y�㣎�olX�P^7����
�P���+�^XX$P',�ZH'*T��ґ`�qL+)e�Uvs&�9&�<�-��G'۟EFH2©w��,����;�u�6n�If���Ϙ2�鬭�,f�e�㺋R/�6���N�vU��r�ލ�Ѵ�����^�,��(l�S+L�r� �P�-��.�e�H+�ODV�ܼ$�ҵ�.�D�x��͚Kn�P�Β*Szj�%ͧLYq?��T����Fe�e-5�&ޥ*�oUA-�ѡS�2���j��Ae(2����Z!��Ҵ��Y���,I�qdd�F#4�Y/)��W�f��ӻ���.ƥ3��v�'�BL�,���۴��q5�Z���Xɲ\Z��	mL�eSn�n�{iT4�n�љWLZ�Y"�XҨ�n�R�u��n�8��d��m�a$Ŗ�t����c��Ɓ\&�',��z\�m��X��K�b�c���#[�-�˲q-�!�
[�2���%Y��@ܱ�Q�:!9kY�P�2��AH#��F՛UyJ����0���	z�*�+.Z�)S��p��n���Li1Ÿ��lXAhjm�ް�����{D�U*V+��,��{pe�Am��Q�I�J��dn��l弘�Lj��q�"Y�D=��N31��ں�}18Ed��U�j�zc�;����,3q�7`�t5[����Q�ٙ%fX��+#�o.�&�u7k��b�G��(�$�˃2��G�1ӥ�nj1&�숝e�b�WW�����ֵotH�<�����$A"�ܽŀӒ�/����: �٦���m�j�b�hE���z�U���i�fɧ%�q(�+�/m��t���0k�v��F���%{x�6�V�Z�R��crKv�q�^,�MPPj��a��jH1��_�Yqf@�i�x�N��6-��t��6v��6��Q�@4l6�0afە7S�R��U��-	gBJ��6J�$�����&��b�U��$��:���qj���5�� �ʑ-�����������$Kӭ�A�!m�
B%T�WM�JɊ�Q��6Y'n�a�\,dz��V��ֻ0�.�kU�ZEmX*�Rc��TdJ��@[��ƑWL|���#�4X������JrA��4p]�'m���ɶ�T�'�WTRo5�Z,�Ȯ�]�.������̷E�#�7_�m�17���!��v��Yp�1�&��J��i��%ua<����#]29or���;�!�M��4����"V�P"&!nb!`�,eM��Y	P�G U�����n�ױ��.����
���C�jz��X�iꙹ T�'P]0�ϴ9��x�m�SI�֎�*�c��U�bR�Y��1]譒��DF�X1nliɶ��*��^j͢ ê�*�SIڅ0��J�BY1�1��h��͛�kQ�6�Q��ϭ�� ljd!z��+{�	t
Y������U6�H�Rx�n� ��;��:ʕg�VJkA����}���v #u�SnΝۍ �ڴ�aP����L���G���9� �Àɱ�Ċ���;��6����h�;!Z)�%M��P�F����F�tGRX��I���q룥IP؟[�v&�^��S�9JK��JC������N����VX�`��h�����MTJ,�z[Ш�1�n��S�F��&.=̭3u9X����1T[a�7q�mbx�ꩮ��S:n&R�ӊ�]<G��m��2e�AƆ0������Xzլ+40*�	nӓH�bM�@��l��*XV��Q <�7$Bٽ��zn���,��4�K>ݔ
��EF&U��7D�7)��&Q�cC�����~l)N5�a?��Zkǭ,��g!��QL�e�Zv���T��jڭq�r蜭�Ӕw*����QX4Vr��R��YFjY(f9�RU�^ �Tұf*3#l]�e�'`ã(�rͪʘv�����6TT֧�#D�^##�;�lQy.�(�(5��ۡ�[ę��!�i(�TB�ƪ�^=���͡PZv3^V�ӐnĴɳ^#J�6U(���Z7����Y�s╻4h�ZN�qRͳ�=��D.e�R��:0�yq#��.��2�%ŵ
� >zo.�J�]=<�{h%��̤D�u`�:.Z{�4�^b�+�n��X�5���P��e�SooR� ��4�O$˥��0�锭̛��P͓��p
���qP�ken�-
�Q���TM8L(++���Ze=(LR�� �X̖ib]ٺv԰��͡*[��J!z�n�Ȉ�5��i4\�Е-�7B�V%`�Ym�e2�l�y3`�����^DZa/n��p&f���� 6��ڱu�+0���1�ۼT0TK"���9.%c5 Qlڙ��[y�i��v��6�V  H�;�7�ܭZ�S��}n$�1n�L�q]��c�`�K*�R�ƽ6Ϋ�H�Ю��i�zv�g�Ʌ7��U�5�a�U{�)D�Є����m����KA3��򥁲�J�M�R&e��AZ��#q�j3/To
���0���ea�܌˚�Ә,�a�t�Y�%E��Yy3i�wSmdn)�穅.A��^\�s'Ʊ�.'�Z��W����U�q�hSJL��M�I���e�CvS�Um�`U���iEz#�dK���$V\:�f�M�����j�9 #@�Z�m:��>a�}������������`���w02�H�qeV��(��iPǗ�^mK�eV�ܭ��k�-Ez ZI�4m�{e*j�vwE"�0��4�i�jEIQ�J�3-�ƳP��v6m4�t�Z��6�&�2R�݅�c2 6��u1����F�i8S����lX�Y�݌�4ک�ό�YC.4����"u!�F�JB཭�i[FI.��rX�Եֵ�֦�^V�H���Bv�e^Rh�0k�L�u�Gx�;m䧏�DI�&�W�����X�h���)�f���R�����
wN�h+�(��^<��y�	�a��%-�9++E��bۂ�nh����qr��@�Yt��qӺM�*�ړ*I�w4� F7��rY�f���3ea�Հ�h7sjn�%���L��2�elz�qY*��U��Xˌ�Z�2�Ƨr�X°b'Ae��3%d¨�&A�N[o��cE��T]��׸�f�z1���V���;k-!Fh�ٴ(d���I	���f	fk6[����b��R���2��cage�.2V=�f�4��Q]=���iU�j8�S�ϔՐ�y ʉ�5�Mt�A��kU
P̨�YK1S^ÓQL��R�x��-a����k�RS_l"Z��L�2�5#�u��E�ӈ�ʕ����x�Qi� ��F��(�O+s�r�'X&��n�`nn�HՇiq�3D5Q��Fܥ�a�^��)h�R���=yV��pJ��:�qm�z�ٳ��nÁc�U�ǀVQƳuc��ոn;	�X�0��K*�U��Q�eV�V��,.�9j�:�G�[��дT�/C&�gP���r��e]Ld����_k �Wv�(6��6��Li�4������QMnB�䕴�cZ��"*fn�ى�����Y�d�a���H�S��H�[�%������y�Eu�c�z�P�f�C��Y�]j�C����bM-Sb�&���x��3X7E��		B�[�v�1�f�a���+����`\�aTA-PPX�G0jY�d�(�5J�7DU��ͳ�S�t ����JfL�2�E�q����˨���JM¨|D��gF)���A5��H4��`������uV���ꀰXN�ݟ�x��Z���P��p:�Y�j{�z�,�כ�ͻ�c.�,�T7�k�������Jy�t����dT���(�-:���w�n��`T7(�p�]���C%��bp��T�D'������+]�7�&��o(�7r�BK[J
`c�JK�4��z�B�&�hR��ڙ���k�F`�B'*�Z�V桂nF-I�M־�6���Z[�4��.b�˻T�di���%�7%cTq�C{Kv�d4�Ϳ����CN��V"�PӟJF�.]��V�	3"3f�K7�� �*�#���Eiv7n��yK/DV�u��і��!v�c��E"�\j�t�S�+�G6+�;b�`^�T� &;Ҧ=$����5vԶK�˿�#6��M¥jSe�����%yY��l[��3"��]��L�֗ܶڥ��(��Du]��6�a����6��qM�c�[���]���`�+[X����\�PGi�o�1�ի�x�4b�2��l�A�>�Y�S����oY)��#°iԈћ6n"�$�Nn��2�b^^�vXLo3��(�Q�U��k/,��"��*Z�A�d`;�<u�	bJIz���.P��N�R���E����$F�,O�}�cě,`�ysv�ݜ��D#��z�7m����X�,soh\��TF���9ͭx���</$����v�7VC�h��ktf�*Cj6�*�ȝ�������Ysٕ�FR�eX�5:�޵b��c���qШF\�e���l�,�2Buk۩Y���yD}%^9x��k2��l$vfإ�Y�-XBN���ac�)�oj�̗r��9�s +)
D�ӛWY�zs6OZ�tQ.����%�ˬ��۷c�㲓ƁTv�4�Z�бX���eu��ϓ�[b�ǉ� �ସ���H�8t��&�y���.e��2�[�͠+3.��{v��m^��G$n�x��"�@�O�w�N�׆E�Q�`�P#��CaѦF�EWM�ֵav�v��K5���BP����%R���D�ڭ!ڡ�1l�ڶ��"��7���:��e�WXˤ.�z��v��i�q��&M`J�Iӭ�rAn�ȦD*����Aس]4sm���`-ҕLغnZY&�gu��,d��p�k�2Tx�xɩ��-;�Z�kX4`� �+F���	������[hLn]%�=e�s.�[H:�$#�闳$�r]l����6�h�oVc8]9iP^��:,�Q�\9q(q�	��C�֠K�j�w�V��̄�+
w2�,*Y�X���ڱS\�
����r���h��)e,D���*v������7��e��kP�3�oKq��(\R�2�������
Z��j͇oN2s]�7�2�"����3Lm���eb�*; ���m@��.n�%��ǲ���w&�S�Y�T�eG�����4ݒ�[S+aZI*��$i�l�cde�X� nT�t>u��!�����w��4�Gp���Z��m�Wou�f�CV����e���v�Ż2`a�n&�AE3̺��Eɢ�0=�P{MQ7( %�=����fh��T��<Ykw�"/D3lq�kv�I�h�.�d�6!/o`´���Itè(jy�K�!��v����(^P�d��9i)��
�X7p�v�K
�ki�p�9nV�,GCq��ފ9yb���� �X�u�X����v^�;��cT���$��^^�O+sP[R˭�0ix&+�OQ_m�øPP1����F��)����ZM(��5�,�Ml���#��-�k*�bٽ�Z��LԑB���EB�ɂ�G���փ�yt�vv����3q$����V2�h�Hj}���V���	Ķ���x��I�tc�n�)��I�l�h�n�޽�J�e:\ܥ4�jѠ�ee�GӉ� �x��2[�l��F�kK�si-b���Z�h;��+��sy�Iե�J�stS**V�^�]�v-Z�IDP�w��Օ""d�p!�%���5z�s�и7h���Y�|-q��/����	EG<h����i��i��*��ޕ,=sܖ^��P�].ta����;��c%5&X�o��ʑF��,%�xEv��#�Ļ�x[ɷ�[G4��l�m�w?�WYYqԯU_:���V3��\ۛ��1T�S�{Uh�,�8�o{[3���1J��`�D�.�]�e2��l�]����=O�#1lᮇ����{.�ِ�9�2��&�X�V�#���+�G�ы��LTA�ܞ�.��/��r�1�^�2�1f-�i�c�w\��pV���`xPw\���f*��Y��q��$L8O��5����L��Aֹ�_7vn�v+7z����+����S���=]W}$��gg͋���B�7��D�5���e�;�]�x#$�ܾ�zd�ܑb�sN_e��z�`.���Y�*��gSZ��yλh���m[�W�5�8n#9j�2��I�7���5^
	<���8TH�\�W�����^3g���eS2���YL��ږv�
	Z#I�+�o��.��`�s<*NW<�{���<_!7��u�\)��s�
<u-�|r�7�fǭQ���\���E:�u�hͭ��g�$�=6|�^y�S���={Y8��qA9)��/.�fm��,�OVC�1�RI��2i�]pq�b�dh�;[���v�V��)˰���3'<��˘�ۚq�.���mw[�++)���8ƘϺ���}������7��r�&s�*V+�Y�+�qm�;$���>U}4�?nݥ��z	�t��2lg:9�^r�ȵt����14����M�C7�l��9�.�lq��5�b���j]��;�K1pi��+؅�SXxȊu.�<���'�EM�d ��u$�s��QbXa�Ǖ��\6(�*\�Ż�N�j�u��i_|E]K>%�[��֖U!w	��[�����lC+Mk���������eA1��DW+(4Mc�Q�{gV�(��g�Y��06%�7U��S�6��^�	�'B7v�؛�'p���F!
�X��nM���c7��J�0p�p�=��Y'T�֙��{�dVeh;�E��mFZq��@�)�׋u<�R�2k���$�� Z�ݭ�����1�Զ��.r�j"��H��{����\��ib�[J��Y�.e��^^�F	B��.���[���*ݼH=n֣�9e�ù�ě[�%:�N����gF���Z���#�ܡ�-�ɦX���nq�}�IP���jU��Z�F���yܲ��:C��EV�$ؼ�yO����n�UoI�%��un��.l��c���ڠ�1֡T
c��;2�Z�p�B1�d�i���.��'fY�\�f��W�90Ji��J;���\lj�EYGX1:'em��ocq��j>緭-f]�Gt3�/��s̬�)I�<M��؂�YV�.�ܥ��c!�9�XȺ��+w$������Iq����O����<pT�z.��:�Y�@RQ���4pu��mw6SXYy&����L�p�E��n*Y�2�R���{��%���q+ni�k��( �N�^��d�L]c���o& �u�D������eYT�����ٌji�jﵞئ�[������
�E+���}�ڗ�Q�=1r��J̣�l��a�ϱ��/;cZ�Lf���:#�:�o*�ݑPa�u{R�PU��]����-�!Z�X�Rfq�6E[/&�ۤ9�R�>���	��w��8�N<�v�j�v�E�J'B����].�<l��g4�:�u7���Km�<��·n)	�1�$�tM�;�yG\�܌n�|\��0Ѷ�� Ιr���N'[٨Ǹ��=�
Zl�R�����{"��c��,"�l����,�g��E�o�'�̙lQʔ\����݀��{ӭtiJ[�_-k�z��+��Η7���ք	.�Ց��1�=C����]�3z��_##�i4:}^�����]�o��B���Q��r�=�84v�)�ڹ��XԲ��̭�'T��V���(�9q�.��yk�˝��X@bt#��>��Lj�<���;2���V�网d����L�7r:�r�n�H-�s��ċf�dƄш�̔6���7*��d
_�%	�����R���Zl�yl�u��r�bC���:�:��>���f'����=��4˫����^>E��d�:ѷ[�m��qލ-�f�y5��<M���'���n�y�k����aj�lk)aVގT3�G���i���k&���.�f�*�����I5S/�F;8���h��1_�ᮘ\�ɥ�"v�vSL�͜�>BK�1�x괚��1����'���T�A�"�^�{V�З�o4B2�'K�UQ�zn�"X�gI+��QQʜ�����ѵݡpZ1^gΔ���эFaYXu�-���u�p֐<�wP�ԧN�v�fn�('E���x�v���S�P������y��H�&�rI�%�S�<��u�^[eK�V�\vr�}����o�
k��ͦ��c��|]��yY��bюm�
p'3}˽Vr�ʢT�l��Q�E�0L�xvqɍ]?��0��zff=6�r��\�5n���(�Xq���E�,�4��LJ�b��tt�H�S�Fo&z(;8\����WA��UD^�F��b��e����3�ރ.���k2�	B��̵�)�뫏��*u�.u�;{+t�W"��O�*�l�t��Bz�6)�%�+k�վ�*��uhQ�O��c�E��V��2�c��qSA��,���iO1�[��Tk-t����5���Z�fd���2���!N���1�`ׁ��t:̾���b�/C�q�����p8��n��ɴ�U�I�W79�p�GaÉ�����n��r�Q�6��v���ҳG.SǱL�Pf֛P��B�W��:�ϗ6��
ݛC�WC���k��a�
6���7w�yb�cM�pU��[�L����F��W���V""�KyBw*�Kc#4�AFԧ�(��	cۗj�m�4Ws�O�N��X�0�nU����M��L[�����}���ԓ<.�ӳ���9r����E�q�t2�#ق�u�'�fUF��Am�W7%
��J�L�ړ`����6��ռ.u���
҄��"k�8�Utz�h��״��2?0m����O�+w�u!���7�W�JE��l��+�,)�N�]�w���_WRp�/���RXewD��THmEhE;�HwJf��Y�����X*�B��b��D��!s"ȏ���Z֡ tay�D�X_b��W���S�㥝V�DX���&�԰Z7)��ߤ:$�1�WgmB�Aq�a[ٗcb�᭾7��������Xv����hH��J��1K��Uvv8���־ޖ��E�2���y�zW2�����]�'5}��ٜaz(:"U/��0I|x��Y���
0�kyӬ�[�ؽ�C�&�!�(��|�oi!ǋQ�٫l�vY��7)�e��{�Y�'n��.�#�ؠ�M�����35\��� ��������6v���ڵK��ố1u����w�V�N���I�ӂ�
����Ù^�uO-`�����(g�����֐�ӥ��՗{#ٺi���(ô%UdK/pH]��k69�K<��'m���I����m�x.��L`���z���h>�;e^�;;Q\��I.j���#C+o��9�Qn�����R�ޓK�U �#*�d5ϑ%�˼oKt=��w%T����]	��u9;�.ܱx����#
�gIx�@�Z�SR`�.c/7�y��1\�����W	)鼾/VsR�j�q�,�e��,hC��Z5�NmX����4k��jo<�z�& $Zvzޣ�N����x)��;% pl�/C��bޏ�FZrvU��3o���H��_��;�N�7��m� O�ү���1f��d����>�	�q�T�G���hx��}ʧ�i&#>�WY��M5i��ۨ�m��
	��������͡J�Z��R�����m�|���N��sz1��]@�:ʊ:G��:��l[�d3\�]�+*VoFX�D��w�.�OQ�\��\R&�:�ֶ{W,��"�t��#�W�3J�M���p����}��̐K:�v���5�af]�D�@�7��#��8�F�CPtz�|����b�]��I�r�of;��J1�����\��Wu��Y�h�Љt��N�g&�U�Vw�ưbR�Wu�ʽ!��;��Z�נ�u�'c!_nA:�s� b�'�w�QUl�.�oݵJ�D�ō��ݵ�/ji����1%�E�-ۜ�PƟ!E�hA��ն��;e3�*b��Ч=y.�aQf�UVS@iӠW���g ���#pv#x�j�\��s}0���"ͦrjd�&�a�����k�1.r�$c�q���Z����z�(t�kxl���G���+���Hû��>[�'Wd)�+�I�Pj��*'��Ÿ��"�V��q��n��K�*��|��uS=�u�h�;��#{�̲j��f��#5Ğ�������1i��i�97u�٠m8d���4"����cyͧe(���v�х*zod{%f�](79����`������^���n�Z��ܡz���ɼ�	��[�k������}�P�.��'OGzЋ���뫎�k��z�ź´�IB9�K�X���0̶���5��f�w�]��v=�v��c�j���R!�+xG�E�؜�q��_�zR�x)���rC�W�ȼ��h��T���v���3��A�����oi�r]h#DjT�znc�$��uy|���`mQŖZ�;l�#8̏�W/���粦�ײ�s�9���{.���omsh)z_N[W�l#h"�3�y���a�*�Q{6f>�2���pySH�Ye�����ȻGk��2�>���2�C&���u7�.��OI	�0���I�ÌN��j�k�ڥ�Ewr���;)��L�R<�i����#Z�8T�:� ����&��LཬX���j��� � �hz�<ާv:��r�"�MsÉ왳ab�U�D�%<toy�O6Jx����}zn���8tcPD]K���js��0���T�F���X�1�6�h#k�uڒ^nު����+�̳{J��a
u�=�s�z��%�YDB��͵�E[Kw��Y��g��V��%�-�ד�w;�x_d@�a�/w.�r)�x�oG5v�7d�u�D)5k�]�`�K	�����j�F�ŵ��7M�cV���t�+a,SaV'\�@�ޟC����S5^f^Lܭ��y��/3�(v����3��qv���m7�p�q��Ni��
G�6Y����÷GVp��EP��9���jK�oJA�Y�� 3�)է-i��ݕ�NV�ϛ���:�˫�O+�fw��`F�'ٲn��։�����=I;�NLO���]���R�.(OI�1���n��L����x2S:���3�O�Z�a\gEњ.�I{H�Ū>u�Kq��!s����	OW.(��r��+���E��]IJ\YB��X�QO�7�gc�\].\�U�QquK���.��D��!��bc�_N��g&�T�n������G�4XU���p��U���A�Ր5���Y�m��Tt��P�z��Qd�*���B`#�S�P�٧��nT�,W��<r)b���m�7�q�F�R�DsZ"ڳr:O���X]�z�L�C�!��Z�P׮�w�-�4�IWќ�n0������HP��vcW������=�����ʳ��ǝ������˕ð��	֢#E�����SB�e�����m�n�ѻ���+2��/�Lg�.�}�b�jB�sT�.��8�)�^�����ͷ2�ɸž���}�u�h�rm̢l�Ӛ3X�3�6��q��+a4wV;1���P�,V�բ䵭�HrT�mh"^��sW�;{%5�@��L*u�;��n`������>�G�t�]h�z�q��U<����'s���O&��Ɛ�Qr�ryr�	qV��)4���&,$�͆����aq�J��[Q�ō9��*�֠s�,˰�r�]�n8
�l,�8;�r�׺�
�2oҌ`�@l����f�/CK���z5��E�����ut�i�Hu���T��|e�6��Mʡ���U��mGaÙ�q���Q��F�e�*ef]툓ݢ �f�]����k�K�F�[����Ⱥ.<D}�
M޶@��_lH���%��d\s�\�R�[
2zʕ�j%<�����W��K��˶�K<6X�TK7K���v~�x����
��`^�歘�re�0�m�(�n�T���4D7+_;��B`�z��P�`�L�{���[��t�q�+a.��lWng7�o�HVe��s��*�Ᏸ���v^,Y�T �f�d�3d��"�����!}��b�/k���+^����-\�u�J������s��e�]8�C&���k8�������"31j������bn��T�f��\Ѽ�[Z��53�f9u��p�S�l�f�|ɱ3S���>l]�V�����d�m�#˄�����]��7��,&�'�hȷ���k��n0�<t��z�P���e[�R��^K��k��H��̭�t1x��V!+�o���/j�ɮ�Va��;)ikt�Eҹ�뽍��E�u��f
a�kK�E�he_+IS5I$֭��}Fof)�;5��IJ�fa}�m�^6��-8gK��=���*�걍r����4��{@,���⸕^���M���Q�G�oI�������\��u󦢍I8aY5���km���mm�[o�>~�Ͼ���w�|�ߞ]�V�6�q��ފ�y��epV �Z��܈-�k3���� w����j.�!���r�65+NK34�Yڒ������%lm_<r�hŐw�a�F[O9V+����lc�E����F��o@��WXt!k�Vu�W8f��$��
�|BEA3s <3F0�L�-�wv���D�B/�;���}l>��'��Kp_]#i����Wo�۬G+oI�aP�즢�[I�s07�5������a�+�� �=˻�>:��+�/U��,��i�����n�
Z��>�]f�����)<��z^��S�pWXI턄�;I$�\	�6��c-w����v� ̳X�Ե%u�KX�HB�3�W5p���"���[���8��VF���h����:
��zi��"k~v�9n��<�/���WL�cX��'f
�Gn@���N��7OH�l����"O�'i�هi%�7[tM�1����;>A4��m���G�4l���f���u��f��یf�:�=7Zi�g�89G�9fɊ�I2v+��hu�P|�]�eղ��5�b�:Y7T��J����l
z"�"v�ٙ���؁��oT�1gq:�W]�5�b2xMe��Ej��}��s�-e`;Xt>�3,���=�vZf���SE��#�S0-ƞ�0QgD%�b��e׷P�H`v��&wt�K��-?0���۪�˂�n����]řY�}��:�;��/�w-{�&a�o��9A��c�sha��>9���bt�H��#`��J��j�B/*<
ז'j�@��I�KV`�X��q�������N]t�A+#�\&j������v�Ӆ���%Ŭ�̛pc�P�G#b��;��D�f�н8�	4����ݑY�f�K��_Hҡ�w�v<M��MQ�qr������ef�XV:�v�v
��1r�̽�`���m�YN�^X������1M[ۻ�}�Bx�9
߲��1v��%��QQA0��h�n�vT�[�k*����y a��/�n�#,V�Bh';u�����a��	Q[x�uN&�Z�i�c�s�p���z`��&�$��Xn��e^�%jM���ŗś����,' ��U,R���#2-9�M����㺼��z& �}&��ಎ�ne�oA�& ���i�>U}�G��6��˖:1�p�Ce�h�	z���H�ܨ�m����90�^^<
JY;I3�a�Wb�i�늁��,���OCv2��徰u��|혖a�x%��� �&�;��u���ER��:V��j��	-���j�Ab��rRm
7]�.�P���+���Q��d�S&�,f�J���߹C]�D���U���]U�����n�'��s�ʄ�R=�j����X]CA��6Fz� 1��ї����Xf ��DB��+/��.Xy���	��%@�FH���!ʻÙ��C�f��r�Zw��� ���`��wg���Od�oM�f%f*n�MT���m��dJs�w�$Kg�z�ugOe,��']]���� i���a�PZ��A�U��P[�RW±�ƶ�ܙ*F{y�d׌e�i9��T\�,���5��O�i!�+9k�����WC-��z*��v�ni�ٷ�2�]����#q�6�&��DA6�^��E^��;�8u���[u��L�N���Ilo
��G��yx��X�8S]���-kܶ�Ԓ��<9WF����7.�7�l�;:���nM]�Ej-�����6���T������v�y.�.�tɹw��w�k(�'����c��t��5آ@nn'���sSz�(�*���%_!������r�{[�,fS:�k3�_��@�Z��ޛg_56t��KnY��C.󛊹mst Rĺ�U���K,��4��Xm�"~��}��s-�r���lk̳j�p����ЍN�� ٭F���]g^��D�+Uw\��1��C2�l�]
�p-�5c��:�������ݯ|�Vb#cT�˛���.0u$^vn����ܶ���7��-̵؉���;�|�0������z��P=k]�W�[�6���qf����"�	���D�݁Uޙ|�X3����Cx��q���i턩�p�$��	j�w0�H��iWpk!;Z�It�3O}�ň�=�/3C�Y��zۖ%�o��쎷���ֺi��뽣�Ӯ��"���$w��SY���`k��JG���� ��h�VqmǀS_i��{��9���ĎV4�h��5Wt��ҖA�Y�c8
�"�.�Y;6oD(�YAr/ъ!g;���ιSTmf	X�OA��4��j�����!dC$��vo��T���]�dwTW�h\�H�ӵ������5�N1b��=;�PS�;(��p��i���*�K(��g��E�A����Ɍ,7�*�u{sGf��/sn�� �`���goU6�������2[5*N�Dn/�����yS4vn�ls�̶�B��5���j�|(u�%�ػ%ٴ��	�k�1.G�����=+'k�0�f�b���V4�R%�W�՛�iO��w\AY��/�� ��(Ξ�B)�ܝ�Q�����<+���f� �w�>�WD�c�y�b�;\{4�F��q� l�Y�Cv30�G#11�Xy/��nmu��>;���g�k�{G��"�Ԭ�Ō�ĵ��\W}Dl�{Z�Gu
k.�R����,ծj�a3�Pm�[-qb���̬c��,{�P��v=�J����Rj+Z4����ծ��m`�ky��-�"j5w�������X������*Y��r��.��u<��窂]�۰֋��L�	��;'A
��)�����t�:�9䃫�{�vY��4�eoQ�;��O;����o���TZ���;J�Rgn����x�0��[��X�P$�rj�ڰ�nَ�����L	�_K�}��.��ׯ��'r�ui]�K>�����M��뤖V�MYzֻ�.����c�@1{jVt�X��O*H-mb�QL��"7Xck�,�	�Ƶ,vhcFt��Qd�T|��Gd�6>�q:[n�^�Cb�R�tͭ��ۃI:�R�G��뙽O��;���B�4���Mv\��+�7�;`�JV�F �mx�՗�%:/�z�b�t�w|H�^�L�'WN�ã�L�M���+�q�y��6��%����׼����J?u���,�L<&֌��Ok1�
�ޕ�J��]�Aoe*t�Y����m�Z)�Oz�2o7V50�ʍ�lDzI���b�����y�0�pX�F����0�KQ�V�:�j%rd=��
�D�
;K��)�����tpV���o�J��+n�3���86���Wʍf�J�1�n�����%M՞�Mœ靹�+��P����`����t6�ր���uve#?��'���LVQ�L��'CTkxZ��;gb�e
��������\��#�AY��١e-n�Q&!̙EZ�4�Cf���!�ۛ���M��y��sv�f��@`#�c�:�־q-�B�g_1�@��� ��#�2�g�NL�yn���.wm�� ��;2��׵{jޗ����'<�����>������b��N�����hf�'�򻚜c���˴��[�V���UV+vD�*, ۬�����b�̸��G�+8^��y�y-B�F��������Ӂ�������Wr��w+i�r1x�ފ;اKM.�6�
(�N� ��NML�Ub�,r+B�v�@��/��,Wr���Ne���NbqE�aQ˰\�����ۅs��1ݾ�եG7�.����2�A�
*��T��D�H�tЩ�cv��@��R��i��!�ŪځۥY�3e#(v�[ͤy�@���1��o��ݨdd*k�0�����uVlS� a��ܨ�\�
��rK֨�])Sw�/gD��m�}%�k�i��q��VUC���Rl��2v�b�"�u[e+�I`��5������H���iy���0��3�msj�K��Ί(lЌ�'l*9y�+gQON��$\f�{ǟbfCd��؃���F���Hp��.D���ù�*�Ѯ���fX���c�뫎�wAlv
�0$� �)�㋸GJN��q���cf��,k	v�U�F�(0ՒM Od��$���Й}p,\j�ʓxst�B��*�xH�w:�\��+��Z�wG�+�Uǝ�/o;�4��4ˮ�4�q�׭"�S�r���4.(s&V'�d�t͑�#���a�2�s��1e����:��g7
@Ga�E��p����ۢD�h��-�����a���N���\��;��)���'j�++iWjw|x�y�f;!	]��z�Rۼ�"do�E�+Z�|v�5��U��H�����ȁ�Z�8����+o�l*Sy���N0�3`�d�5�.��!qգZ��.ħj��`��{r��AS��`�IMF���Q�A�ܤ��r�+��,��҇��k�7��p'�5I�v�A[#Ux����phz�e�ݜ�Ԅ��*]搽���D��#GJ�X�6mu�u7v1c��rtmR��o�	r�C��E\pIA���˨���muK�]u�ٸ�dT�ػUi}�WCm|z�Y����F
�;1��0�KG�)[z:�A�;�ΥJu�D�V������v˺��-x}�	�B=�+��/�S%��=Dr����٧.V,�r��5�&;9�C31��)�Wڤ4e��G��{Pu,X�D&��R��+�8�s;�V�G.�^E.VY��X��V �_n3�R�.�`G��2�82�J������v�but��}��9�wh,ԙ��A����S i�{�stZԷ%���@��� j��ƣTVH2��ﭑ�L1u0������v��fDi�ܲ��5)9�\�.�ba��/���J��9�7�xD�nV�s4he���f�u��#�Ѥ���Mb����k�:b"��C�(E#�k҆WL7@�v�A��KcD̲�z(�1,�\4c��W��� ��b�P�{��]��P=�2��Z#���^*�iy6�C�hŀ+=a��yY�tɏ�$I"&v3�f�lǕu6�7y�����n\��ղ�̰�]����.dx	u�@�T�SF1z�ص嬎�\�a���ML.�%j��)Z����SC�+h�j&^f�S�wl Y0*�5�.F��6X�5�B3Abn,+���"�(M�.�X7O�)���x��8���&qo��՘�)�9%�s��pk������:��w�3�n�}@u���lL
��B�$���d�{Y� ���]Z�쿛��G1�O�t]���3�xs�BNf�K�7����W�o家�܏C��!g�uf�����)�G��3�]_@l�f�Й��M2]���A�3��^}5䧒q�"�L2�{2���p�oMO_EMd�۳ֳ�-5�n���p�e�4>�B��/j�Ւ���7q_9X�Vf��H�hvAk�m��x�f_T���@|/=�z&�5��W��;L������[}&�[|XgfB��Ӥ5+�
H]�b�BsՋi�P���:��V���+����)��mXX�[�O$*�6lEL��']�ۃ���wL�s�HZ��g��z�]�L��I:6@��a�u����u���/ ���J���B����Ķ�f��*��ഹ	|o��v��ř��-�.�2-z�_p�ܚ��ɯM&�\qaL�vC�������Lr�/�9Z���0�Ջ�1�;�q�u��ov��wBhH�tL1�m@y�/��h`1BVA06�U���;+���cv*N�-�%Pm���7�rma�x�r/w�e�<��"�@��Z8qށ��=�f���e:#�&�J�bd���#��ky̭PV�Ѻ�ؑ�xϹvj�P
+X�"��\�^Uh�K[���^I�TIl��"�D0�v���o�U�*��Ƿ]J�	ы���}"1���c�kFZ��U��ofԠTө�:֚�}rN�� p�:����!�`�e�� ��9ֻ���o����׫�6ü<���c�J�r�3��	�dd��s��gCƓ'xS
���pT���|/i���Z�NI��낰��AU�:]p�wY�ԩ]�o�Y��m�t@g�
�|�+�`!&��Ň2��D&�yѾ��ڮhf%{�@���T8�<;TK�
��#8d���H�:Bv����c�S� ���LF��>�`���W��qj��k�:}-ͬa�$V�:N����(�c��-�`�OJK��!��Ԓ	���
���&C�^8gU�
S��]0�W���5��SR���X��-cb*N�"�X���ܮ]6-�X�<�ڊi��E��=h�f�v��#V�ဤ��S����v.�7��ʆ��;p:�����^�r4q��ckD���B�����BY``umf�3U��P��c���:��m���8�N���d[n=�K �WW]�X�D�
�<d�c�����M�am���n���iÙ=W7aQ�	���jצ���9w��2ٮ^u�L�����ۘ�u!�p_{���9
+sJǎs�Rڣ�皨�vS��wn��Z�)mM���++�m˽+�^1/�/dy"��*�ٺ-�>�9�T�T�`��6�@�e�;�^���h�61pa�Wo ���#�:�{�6�'t������Fu�E�+����oy�z�I�Z:Ĥ���yLm���;�������.-=����]���9Y�0̷��D�{���uJ+72<��ew&
�lK��c<�y��Ž~/��0�ꖍ�fY%��u�Lq�Wk�驅�e��
]R��c�3�{r� �������<=�O{�U4�ͭ��kt�
�^�f�Y��}��*c"��P{]��Ő��C��Jp}OY��m����)0h]V�N�k�����/����w�������O	32�,������A1�A9��̏����(om$yd=�e� g;w�ˋ��(q�F��ng|M��,KG4�oz���C8y��z�vErB��9�ܽNkh��6e�����N�"�m��k��Y���u����	�Y�h{��� 3�zu�ٸ"�MT r[���wj�JC�֌D��4�.�o��g��$��צ�K�4]�oM��i���6,]�L>ɦ\���cXYQnc`���,��t�����5�"5����b��b�,Vn��j���$Z�l���d
d�p3.��Z�;q��vW��X����*$�<CQ=�,e��h�{I����dܬ�=ȟ+̪^�)�jxQ���Z�q#��+&t7�&�uX4T7�(�LbF[C�b�lMz��s�ř��&��2���5��7ǖZ��1�!t&�rr��<y�[��,ɜEP�1��!;{p���v�T��8��5c`��I�؜U[��)�ץ���`T��Q��W��*v:bꝺ�o�L��,hі��8��� ���
���Ʈp�ג��
I��d�gG#J�`�.9�*���wӶ�[�x&�Y��u��Vc+��b� ��Ÿ	!�81�ƣ3����1�9s�(�&Rq�ēb#s��
��1��Q�B2D)Ѧ�1&�8�D	�D�b�C$s�B�@�ȋ��\��P�(�2F��	�Ɖ,9�79r�$�I	��IR�cƚ ��Hd����q���.X��D	rq�W4�M!�D0I4dFLH�G��
a$f$�@�1ȉ3!BSfI& ��#q��� f�ȍ$�E�bdB&#$�{ X��7o4�h���5�Dj���nd���r>�av,��p�n���뱭�h�Bc�d��I�.��Q$E7��ί=�j.�虜�C���I�54�"�ZG��[y�:�栃�T�ƭ=C%f(s��)���N�Ύp���;KŌ|�A^�P991�v���.�z���A[|�g���:�y���U�V��~WC!����4zҙF�+B1p�-}Δ~)��'M�ת�.&
���t�<l�w`�Bv��
������d.�&�@��%J��	������Ԧ�6c��];�x��h|������=2b�,�!�0�5�stgwk4G}�h��U{ֹ�v�b��_d�<�\IXoF�e����B�|�N��7�LvAG��p��z{���jԇ2���]}\�3X��k�6a���~�Fe,�ws���t%`��U��
���Z6wd'�ٌF�����|��UfF���U�g(�{��9��ҋ�Vl��s��Om��]�4^�8����wq�Y����O�lq��;8$'���oI`���iq����k��D�6G��f�Wy���ӆ���D5A��'f���]p�8��h��*��|W7؉�ʼ�u��wv����ǥ;�����7SrN��f6�x积����T��J�'T�S���y�ؽ�Xo,�;�*��w84��ڒ�ν�k�5�j�r��C�闠豸�ƻ��ō0ڿ��Q�z��{���!�t�L����4��QY��s8�Nt�h��麸*�g�!�ӓ�\:�c����1&��L�]7vq��a��f*;��ڤ%��N�&�u
邵���e���c49�L�=w�����%�#9�S���hխOr&����H��x�":^w��.���0�V�[�(b.X L�:GV���0n�w{6��ϡb���d���[E���Yu\g�g�o�1W�������bn��{����y��~ `�q����S�����.�W��ZrM�<Ƒq�K�]a]�˶g�wUy�4с&R`���i�����)%�j�J�� �e/eM�0���Z=�vւ�Y%�s��˅����oܗR���tܬ=Iʱ��cs�3�e��r?.��*3�����{P��"�6��&\�E�FF�g�,���ƭ���[VX��v�0��^k��;�Wց�5��{���[���yׄ�c���!�S����8����V��U:�������jo�3EC�~����TUa�E.�;\ _M���o�{���0�X���);5�tE���˂�4h�An��3.oO6AL�)�3n�F�ψ��]t�˖�\#�����/����o���;����Z�%z%����,��⨱��D:Oy��$<�4�Y0�1'T�����M��c��K<��-���|ug���.�ٷM���q��(	��Ft�RK��8�9�p�k��V�.#���!�K��y9W�cvَ��hd�Z�W�t�ef�,�/�=Mۅ�-ו�<��4!���T�ps,<	�aSg���G��A�x�2�K�L�y{�%��=c�`�5-o�n��:*a>�G?\>�T�C��4�&�H,}�&c�Hu^�f/0wf�m�z4 ���߽�k���1M�}&z�97�KB2P�r*�3��)���
����\��^����݋JR�j�G���@=����X_��\9�./9�=N�/{��`�sM=\��#�֐_|=ݮ��3��u����K�ߢ��n'��~<��b��"��|�A|p��{ޘ�+UrD��TZ� P�x�U���]s�v>�����iU�ľ�a��B���:a͇V�x�ɒ��UI�(aE*�A���������׽jR/�K����̉vB$�i�F�@��x(�)Y��O���n緼�l�!�N�Ջ�_���\��3����S*��9�:M0)_	We��3�	���S�s+�PH���p���q�h=Ds�+�<1���m,���rg4EZ�c��x�W��Y�2�whR�yX�nt/
��ni�=9E�s�� 'Qs�QzmB�0���7��М|�u�^U�V>�+��tқ�X1�	`I$��C�H1��n����3틅{o6x`����K¶�/}��H���I��5d�j� ���i搫 ��np��j�p;�J�Y�;��x��&9x�nv�������c��U�Y�����f+.=���$�S�����d������!.�F����5{���CO��\�ɛcm5u�^�����p�A/�^����K ì<̯N������fS����]�:a�J��#!�L*1���1��`10�p�o���8R*J`j�=ˉ�q"�SR%�g�x�#C7+'Y�dچT��t��u��|+8B.��n���jkieX�x��U�؉�ʁ�b�W7��<]dݏ��Ll��P�1���V@5t�T��f���[��v����*�%�x@=�lz4�B븦.$���@h�~Σ�yM��|�8f�̉Z/�\D��'�~�@�S2��PS0�9��H%M��Յ�9����ί�H��v�j��_%���������չ`�z�0iԸ�.��6����<�3I	�h�q�I��ԍv���x֬]uS��1�N{.v0�^���UR
/oz�9Fܮ5�mC��UT	�3%���/Qn��<�����q	^�����N_ΊUT���:���HJ���"d�xcE쯪2����>D�s�@��==�"���hdQ��ي�d�R~UA*��Z������4��XRYZ%�j��Z0�q
r��O�~��ܣ\�er�Q�Kg�xk�d6���ɾ���ޝzL���|�Ӥpy"\"���o��CGܕ00�q<7ǡ�cbޓ�Q�F3^�zf6e��������3��K�"�U�m�r4����5F����i��S�C�k��3�x9�8���~
�W��݅�Pl���!p|r�ٹr�H���Y�70&y�̘ƚ�ѐ���]F��7d���ڬ�5�Z��υ��ҏ���&�ܼL�EB�+��� pHr���T<rgXV;fCɸ�P5	*TZ��=CPp��j�W�:�N7ǹg_`8>��c.d��Yr�Wc�c��sݜw�v��.���t�[�܇��ޱ@�xW��t�veQ~`xX��<�An��6Kc��ۡu�;6��Sw.��,PX�C�簐�ED�]ˠ�e�7S ��xGg�A\.5�����nIܝ� 8v��X��O��T�
����o�xb�}m�(+A��	+5A��Z�e%V\�*uT�* ^�Z�7�o,�.qDNNv���/���� �z�mN�גL5mى�X6��kq�TG�
�TN
�G<Z.�s���A��"�k}�Ǜ��b��'��rVjX4g�*܍�q'�G|Y\�cU�pW�+���]C�/v4�Ӥo�R���6t��{p����.{>�;=`�kGN]R\��u������wm��t�W�ԃ�^�P�r����f��o�v�˱P6F�����R�[ %b�I�@
f`������y@�[�j���=M��i8�C�~�97�-v��u::�1�P���AA���s�r;�<�/;C&�E��bF���Y�O�������j�sz�&{������ћ#]dm���g켜�u��,������i|���6*������7}�C��@A'�0���L+w࣮݅��ͱFR��'g�2!`�qo��[ێ�9t��_�Lk@����j���t��=�x���ŀ�9��,�\�쩃3��T�z��(�(�[qF$(9��(B�嫻�T�^�ч9u�����с'�y(R7�	ίr�� b�cՎ=0b\ܡ��:��hލ�DD҄w��F�u��M�u�wW�]�a����{���B�wo�"�W�����b��47e]svˣQ����b����)f�L�K��A�c���6M���$�f�dmv���5�e8�t�h� ��e�<�i���,�+�G829)d��Xn��V��ce�\l�����F}��`�Z�Y>��C+O��3M�z?���'u���:zѤ�Tn����!��=l����f��T��3<!>����"�4.���^ƌ��s.W�������5�z6B#/��̛�a� �خL��c���e�ޓړn��Ӣ���ʧHfdcԮ�&6�.��(�oy,�n��:ye����ԫ����Nw���y}=�ws�Sm`s�M�'���n��c$Ft�Yո�0DePv�͎�j+W#�Jr6x%\��g�<�u���p_LQ�&����'D�+��z��Q�h0�1�G	�C�3B
�~W������S����tz�t�ج���E^^p�Vo�Ez0���L�r�x+F%��ofB�]A�+����K*s!�KSW�[lL9��w3��,��J���`�ep
���!+R��;#��^��Nk֬���p���/��e����)v�J.vF�ŘW7C����|*�U�d��@��ak�l���5N��
�n	�Œ�W�.�x=yT���*�Q���ÈPCK� �|ɧB����˃
��x"k�2�vQ>��y犻ع6�d�=1���]�Zo\���}�특Z��6ɳ���+��"�]��lb��C�] ��뵵�^u6���*�w���NqE=awd��򅭯7�>H�z@iU���»O�+Ӂ���i�⊿w#~��38����6y�a������<�& �(��@� ��f[,f�)!�7��ZD��!I����!.�A10�|�����8�I��+�o��ey��q�AsReO`�Դ_˙��hA䝂-:�֦����b�q�t:ٚұ�W��0G����A��7���*����{�!8�$뼼&S���kY;^��|�/'��HC���%et?^6>��b@Ýu���vP�=g��
\'Z*_��7i�|ǽ~������gF�;<M�`�G1�J8Z񪌘ɾ�L[�2��9mr���;���-��
��U�&~h[Vb������TDz��t=
?����<r��βDh9�ڻr�$-��W.������\�3����>���x��(��j�NgZ�^'�P�ֳ��b�W�՞�C�J� m9�q��J��#!�L,��t���9�`�,c8��N�6��(J�N������y!^�&�3�7x��˙��R��lYy��ߊ����F#tyu��̨t?nq�t6alM
���=�{-��m.��"��U��^V�!j���ׄ��)AD8�j���_U�9WM���=�V��s����rm��ĕ���_]W~��#�U��Y��Al�2��?L�Y,��n�����e�3HJNj-b�Z�\��cXd4b�������do_��$?s��s"y���}5q�[:�a�:͎'9�Ξw�L�u�&�l���Oy����5�q���J^2��/�vb'��K{������aDr��m�"V����N�7�?�d���oÕxS���q��noH�&h����k���;���;�!���
���n���;��tP����qdЉ�v�UZ��we�VV��Yڥ���=ՄW�ŷ���Or�Um40:��0�02�,T��PJ���ԂP*�ay�w��g��P���#}����u��B��:~�K�ʖ!�"q����]�t����!��U�SJ{�u����	V�l��E��M=������ǈ����N�=�$��=��=������S"�����8�C���t�k�7�W�)W��S��\�l�P;�,����w]�L�0�9�!77/�Q���{mG�98��+/qv��8+��[��<��һ�=v���]�2�o)]�,N��4+0g ᥲVe�W;����K�\��t#a�����m�<g6
.[�RgqW�v:��k�Wv��K,Kv���ji�L]���!l7� t`R68d�V�F���<�W��A f��94I����l���l�]L���;c�-�������Լ���Y�	�)�ըʋ�V;S���ڛpY���l\g[���x�f�_-��qV�jT�֤*�q�T%1Y��R]U'�R��ӑc'Y�#�4����{�ֲ�S*��e{qxE^���T�L����[n���F��r���$�U�|+��:q;2����
f���9'M�[�3s�y�*0������۾���WNm�h2�}#�;�pW3�-�N`w_�} �P�y����Y{n���̊wc_<�W���eL+e���Q��#B�\I�F����F��ᮐ�q c�75VEF����[�w����V����nSE�dEa���
�����<ޒ;��7wx9AUq�y��7b�[�Dl���LэJ�*�k�b�l�7{$i��j�*J��@�U�ǻ�Ƒ�!J�����w���Nv�Z�q��l�D6:ro��Hls���1����0�+:����]�����ڕ�5q吊#m#"���w�����M��Χ[�L};����ભ��(�e��;��%!ѳ
�Q�`r�PKQ�����V6�."��jꕺ�c�	�� �YA/��wrj�2ܬ�D�0�h�X$̓�ۜ��3re7�w5�{����9�vx�)�x��S���Xط�*q�d9�Pj�B ��|V�'�k4�E`����d��M'�n�b}��)�Ѳ��3P��sqT���Z�E�2��[�a��fvgIgh8tdN��o�Jwx"�I�F��G���d��n"�t��Y���ťKyU������j�Y����aFn��C��l.T���u�����i��	�ym
*otԞb�3M�=����U��m��Υ}��lh��
$֞�Uܩ�/�I�ԭ��T��n���Y]�K8�w)N+x���s6�/0#��U����mj0.8�!O1�G��"�OiXGh��-�8�}��t�]Z��Z9�U�Y�o8D�MF6�F�*�WʸS��(���;�A�o�Q�eZ�eX:���ّ��d"繽ig/�%R��S��Ŕ:��o8���؏A�c�ޝ�Ѓ���bx����I�W4�b�6�r�Mw=6Fm��։��tő�i�5غZ��.���h�����e�]��pAW��wÆ�v��kj�+�As@�L���Ӄ@�'[oT�P
�
��K�˂㥽7t�7�gP���ͬǖ�5����yԳk�9�[s�I�so+�n��g_(��Ū�Y�2����@Jm���d���h�CU��h͕r�F+o����
n�N,����v��qnCILx-�V��Y��vy�E���¯���^Ԫ]R���!��;{r�v1�Y�j�����9�G���Q���M�&s���b|����܆ࡴ^���Foq��avQ�]5���f�`aӋlu������iG&nH�qjP���0�V��G��N�׆UngZ��it�{qLLM7��L�ץӿ��n̾�V�ݷ�s�u��v�Jս]gq�W�Q����lVBs;�umM[̲ьo �wz�*���k�ZE��Z
�>����`vs*����Hΰ��r j�r��yR�ȱ���WK`H��a��U�[��&R��c�7��u7�M�ש��j�P@�c��Έ��Z��p�8�hV�#�Ħ��5�M-Փl�W�X�ش�,YPd�B�PA�͙g8;�4��$]�4_lr�6�*�ڎ�es8�������Ov��ز���H�NH#�+v�ot
�E�9����.oI�,����ڰ�:�c���\��B�|"����n�ϰ`S���A�~]`����{w�ϻIN���'}�2K�~���"�20te������H[�/[YGA��D�\�X�w���,)|�clw+(��n�xu#��X�r1�Ͳi	`wj��7X�>L�yvw��niΩ�s��{Ry��I��\�(k� �5#z��n8#4Z�9�����h��d������ D�L���#"�q�1�Cs�"
)4P4���#	1���90F�$�Q%	�$�RA,�H�$�H� ��dc�(HaFJ��LdC$�K&	7g9�qrd2�8�Jl��d���0���`�F1%�8�d���"D$���ȹˈ�	DI�
0�D�Q�d)�0B�79�9\ь��"��H��J4Q��d�K2$�\A����R��M�q�cd��I�㈥F�˜�(�i""I,!De4��_� ��ɖ�h�9`��bXk���TW�5�r�KP����wZ�mN���c�q� ����x���ԝ]�L�m�gVZZ��/%��uϰ�7m.�Ú��]-��k�W�t�{�+�r���s�o��.������m��-�]+�}�ջ������s�������������U���~��{~{o���b7KKc��j����`�ݞ�\�9��t��y�X��q��K�W��z�鿛s����|x�����u�x���\���[��WO]r�m�\���w����KŽ.����U�~_��}W���~��П�1�����*ȻvX[��G=�T�\�r�߼�ݏ˦�6��μ^��nu���.yץ�W����?s���.7��������]7j��*���F��6�ߗ�����CQ�?/�ڽ��\ R��܊z��#�U�ڭ�7�������z]<��Z�o���7���|W�����~�-Ҹ���λ��x��OM�{�y��/Mq�/�7�u��k{W{��t|��.�龺Z~�M�����v��?C���9tXrB��s3�=�\�'럷���Ϳ�����]��=��\����m����M}�}������_/����׷�t�|��w��W��t޷�:ۿ9k���{�Ϋ�����W�}�M��6�[⊘�|����%�҃����}f`N�����һZ|���o�����ur��M��}��~W��n�B��?��k~W6������|���?~ｼ/kF�������[�7�����z��B-Ϣ\:���Ʈ;nߐ�9��\y�r��5�v��ҽ�yn��鮗��u]���Ο�����{޹v���mҽs����6�\����[�ߕ��nz����騷���s�}�㿜���T�f776j�K�S6ʨӱ9���N��|U���F��ή��n-���_7�Z��cQ����{^�����{���WMҿ��ﮮ֍�_���^7�zZ�v��qo]w�w���].�V��d�8�|�DvI��#s7�ɚ�v�������{�����W��[���~]-��;���������oͻU��/����ݷ�n5��?���m�t6�qo�ӥ�W=���5vߖ��]r���}o{��_�X��1T��[�2�_!�L�6~�9��?v6"�����םj��-q�{�u��q�n�M�~���ͺ��oן:�������;꾫�O�_��y��7��m���^�v�6�[�tۥп�������<<�[�V*54����m]��7&�ڷ�[��^:�2�貕�bƛt2���ի+bΜ' ��
�Wٛo+D�����)3s�Jc���!]�S��.����CgѲ��lZ�t�աD�̣3�4��7kEZ�*M9m_Nj���J �I���}���\oMyy�׮m��v�}���n��v��~��-�y�v�6�\��9���彮�sWM�~k��y羯�h���u�zk�]5w��r����ِG��w���5���ܯ���#�#�_��m�u���U�]�﫶���������{n�V��*������{~Uz�u�/�}[�~Z+�ok����/>�o�Ӣ��5�����}R�_��Ҹ��q]�9n��n����\n�x���s����x�n���}請~m�t׿��{W��|�=����K��z뽼n7��ow�:����6��-ߟ�߻���[����eMWغ�_���?d���c�_���-q�[㧭�+�x�-�K��~WK|��^/��\�i��������?�t�W������6��-��s~�<	��yOg�=�
#��
{�svr�֣�/�8G��^��3?9��?G��b����M����^���>��u�y�ݮ��\/�w���ݷ�ܮ���?.�z�˦�ns������]r�����>�hz�� �������a̋���꯼�^q�ߟ�~|���޼��ok�]//�~�W����έ��_��o�^u���qc��n�W��W��6�\���x���U���y�w󖸷K���k��:��}WOu�/M�U���{�M����:��˿~\���7��s폅τ|Bd{�t��s�<��Z�o�t�{��{�.����_�}�{o�t����v��qo��請��x��O��u�J�����/O�v�n�ϗ�t�o��yþ<���z%��TӉʾ�/�"�aa����;�n*�w������vۏ|�+�y��鿾��n���Ζ�~��u�Z�x���>��^���������^/mt������[�DW����]oKO����W�9˟s��s�MUtn��a�<�y���� g�׼�k��>+��+�9�������������q��=u�������W�}h��q����]^��~W�y��׾�k��׏� >��f��w�>ž�
�	��'�y_��9�v�y_ߺ�6����5��+�v۝r�rݷ���_Z��|]���׻��+�]-�v���t׺��w��ŏ־o�^�x��͕S��2=�(�5V��ݳ	�.;��MNKF-E���yvxG?�k��q̐�+��M+p �{d���9�8Ŏ�yay'2�-ʛ���֔�:G��y���-���kKc�H4bz�w�54����U1�%��^��V�FR�٤ZUk�=�ʹ7�R
��:��b����> ��}�����r���y���qWO�O^r�hݶ⻿�x��Mv��|�t����_9�U�t��+��hߝ���o��>����>�DW�*����am��z{˰�+Z��}�}�S~���b!�	����qx�����|��W���6�����ݽ��Ӿ|^潯M�������M��׫��k~W:����]j�o��������>��Y#�w$�3ALh���>y�;k���j�]v��t�O��|�uWcb+�����U�i�6�w��龼[���]|z��ߜۯ�^���W�{Z��}���+�D�����UDG��O�l���ߠ�B�������u���߿���ޕ�Ƽ�.�cQo�|��oK��Z���]_[z�6��v��un����-����opU�������+��:���}U�/�~o����W���W��U��HW�_#�@\���P��=������m�n:k�]1��+�����5گ�^�r�o��-�\w�]6��Q������~u����:���n*����~�4n6���k���_���w�un���]+�=_�ysϝ����W|�:���7w6ｼ��>����4�F��꽷m�~WMzk�\W��똴��x��뫷�ޕ~\ow���Mz_^���_.{�ںZ�����������yX[�{�G�}�}�Kh�񃊶RS3٭-��ݍ�Cޓ�}���`ID\�/����[��t�w�zWܵ��5��]7��o�y�o�t�k��㥠؋�s���Z~���o���<>��A_P?���n�*����亍ߞֻ��1c虙�}�~�Џ�]-���U�\�m���{�?��*�q~m�������oKv�?�����z�~�����t���^��v�m�soWk��*�6�9E����������w��]����W}��x��>��|>٩�������~wo��ѽ.u�Z�}W�t�������n>����y�v��ŏ������Wk���r�����Kv�_�vݶ�\�Q���+���]}�|����y��L_���
WVi�u�����3�"=��/ޚ4n-�u�k}^.����r���Ҿ���ݽ}�7�|�z��^+������_��xߕ������5���^+�Ӯ[��^r��<m��A��9��~�f0��;��赀��+S���]�_]p]Ö�B�4,�;i�:�9T{�9Z�{{(�Ch��:��YzF��{��4s$�Y�"|`m�YȐ���'J�=��-ƅ[N��\4�s��N�5�8v�|�X���Y�Fk�J}��	����}������5�t���m��һZ9�\���n��]�˯����zmǿ�����6��ϟ��ݭ��6��{��7�߾��o�ܵ���[��]7�ρK�Q���|��N����U���������:�-����z_������m�~t�O���ѿy�|�.���������<�WM�׾���/���{��������>���tۋx�=�=�zHd� H����䴾�J����<���/J��ۥ��m�sηm�ns�?>^��F�ۜ������������o�r�o�z�7]����k�}ux���h޻����K�_���\�Cx�F�1Dx@"<J���[�>�&-,��z������:�/��*���o�~�o^��m�Ϟu]7s�qW�<뵼W:�7���7��Q^=�hѸ����.�M(��[���_���n����(	C�� ag�ʾ���F�������߽����㟿��W��7�u��t5�\o_9�+���[�_������mү�����5����;|��ֽ�������Ϋ����qoy]y��ݮ����U����qw�=��o���W~��������֚4��4�{ퟜ��3t��������Z��}o�}t�M��_w�ު�5��wϾ��^փou�����|WKO{��=Z�����y��{^֍��ow�+��[�]*���B�۝r����ׯ>�r�U?t}Q3sw���5}�I��$�����s|v�qo�����z]E��U�]<m���+���~=W��?{�ex��LdC5�stgvU�S�f��r&j�����h�����hD�a�~|�8��E��}f�	�������Pr�b�20�qu��GX��g��p��M]C�>��v�~�¶6�P���wF2f!�2��דh�t����	�;Uc�·�y�j?�ۑ�r��N�;��#�5�qv�\�Y�qp;l�h}Y���֤y�ih���q�W-J�� ۹�R��
���!xJz���!.s������j�R���̎un��F�A*���K��K!��w�][EI�2b:؁���$� ������#�V-��=���K�����DO"�F�9v��&"◹�i��	���'\*=����kd��H�	5r��Aj�b���\��F�o�5A��'f���\)�

$؃Y��׬�n�S��J��o�*]��@3S�Ы��h}p��a�_T�6n\wg�q��vQ���lrV�ݻBz���ȼ�E����M�.�Xhm�`[�j�b��+Y��t����S��:�tKệ��gu��R]����z��u?b��XM��n�*��.��ݲ����۵����*�1�+���@l�>rg���D���\�@+۪���} $4¶�eE> �-v�m�X>�m�1�`&�5�K.fvo�"�j!�W�"S�_e�w(��t�U�v��<d�q�"����{&�O,��!�Wo�^�5 UL��y^s0���F�v=+��É���������Z0�2tC�u��sY�7{`(�R���^�V���g����c�p��DW�DMFJ0!��1֎����2�R/�253<!8άyUq�\�uQr�=X"G.���|���ٷY
�C�����a�䠚�l`����{���(c7kk���G9�Ő����6k�x�M;�*fHV�g4��^g�oV�Mu(l���#j��6J�]8�$Y���tVM��UɌ�=�uP�-y�a��ז|.$��n�:Sk�������6D0��B#/���޺�9{���@Ȇ���5��^]f
i�b.�;�>ܯ�-٩�ǩ]�	��vǔ�%-��p�L5"�akR73-�]�8UC`[��m\{��[k��S<O�ĺ�8�Ua�eH�fWCy�%�h8wQ��R�Y����uO��,"��@�6��5:�_c]w;�'#Q\�L㈚��j�f���FhA�Z���u�"��a�L&9;w��V�.BA[�Tfv닧��N�)��� |+���?۶�ϫ������o��9�:�c]S����2�i�T����f���ƍ$��W ��$%jU�gdt��額�,Sޙ+<8�S>P�^Z��ږ���u�h��>2֡��Li;�Ҡ��[Z_��F�N^(��B��҂Y:�iF��뎛�X_�ʞ�9��4~UAQ�2��~?�ȩ�Z3�1y�;R�r�Fc�1�c�~I�A@u�����p۽yX���'���q,�
rVg��fk*e�*�fwn�Ýmu&
�z�
*��N@�rq�6���
�s�l*��x�>:���[K'p�i\�1r�7u/�������L;{S
�R���Z-��8�#$��o��u��܁�b���̼�>敌[Ln�A�Z�^���6�B_��T���k}�T���V�i�y;�#LB]n��Q���U�|�ْ��UM��iah��v��]CP��=`>cK1+�Z�ig�:�v(hrL�:!:��y:���9���q��+�B�RiF�K ~�v�=�dTl{�\/���v��A��A tёz�l�>ԍp�5I���.~z�ԃ���k+��γؐ?T9�^��>�fW��"��[�/�Z�=����Z+o�����P>D��hU�&_���#1Wk�К���ttRa2򺷚˃;+��:�GNK����Ͻ�ҹ�Y�DG��� %��NOt^]�t(�c�us��W�xEDZ-f���]�:���\�������?CS{E+����W��ٖW3$��8~���ƒ�l�@(�U:�S���*����L,�5���`��VymC���q����+��6��O�ّZ�R��e�����:��+%Ҙ<dU�d=6r��5��SV�5������ݶ��4#�x�����bC�:��
�"� �m�<5�=�E�D��{@;�#df���{+��t.�'X(�e�z�Y�� َ9���k��mB��oU�ȫ4̋�]N�ef&��}�U�N�W���һy� Xz��έ��]��=�5�HݱȢ�U�Qˍ���i��L����m֬"��Tu�%q!i����5�L=�U���x\�0=��>���ӣ�E}_F�����ب-Ʋ�5ڔW'��!��cT����+E��C'7�?�N� {V#�N�w��nG�m�M�Vb�h��\-7;�![W�1�g%^���DV��Й���r@�&�S7�Pַ)35>�:9�dMV��t�դ`�/m�a���OrUo�P\���yѲ��� l��r����-҇�䏹B���b!#�����xe���N�~җ[�8�#�7K�kz��8��:�MJ[�Tx=����a!�J.�7K����o�糣�P_/�V�q�Ƚ�ON���e �%ә�S0fs��ص+��ڕ�<�"�P�c��S���J�{T��Œ��#�0��8ډjMr'�w>&�P�q&OR���e�p�X�+�n).hѳ�Me�`n�XHlr��7�a_�;����]dN��[�ƏZPW�`�K9%�ǻ�����oM6)z�9�51�ؖ*�{ʲ:=�X�@�N��OB��|e��&ff7�hPO%<����ɘ��*Yvgf�M{|n���e��xГ_�f�d�
�&��0�����	g"�����Q�h,6ѧ׫.'�ڶ�N}�y�W��+�f��^ec]\oY��(<zU�!Ѧ�䕥ӟ��>�#U<��.�T+6���0�4��T�%9�
d޵��>�UØt-�4uL�%��k\:�r�ݽ���ךi�}ma�@I\½��q;0�`xO�� �oM� �]AH��}	�
��6�f}.:�U��6,w����{�}�lW0�7��fR���ҍ�a<%L��|�������BVn�}˘W��=�g����N\] �<�
G��kjP�<0��fr�T���֫�Y<�ѓ�^=0���9N��O������S�S���ՇK��ձ)���V^�5�u�9�93GR�����;0�L[�7��!��p�����ȳf��[�q�&rh3R똨А����c�~��ӓq�-v��u:9��,��u�c2��n���Ꮘ��`$�Z�E�6�&#j���B�`��zz]4~�`�u�v)��PCƑ��6�=�Z�q\.&�����@�TK�z�ثG����;��Y2,N�.Ǆִ�"ge�mZ��\A�'���D�����ex�n�����h��r�u,e�8�U�iՙEg�����r���^��⋢����9{�d{w���%������� �Q$�t:]^�n��LAg%����E�M
���J{(T�*5�\�|/it�\���lqQ�8:��ů�.x�m(M� r��Ze�SQaR�wm�EE�c�g���}����)ڲE�w_�N�m�0�M�HjYs3�q�s4�T+���|��ّ�irysV�]�����@���hi�K�O��	k)0�ٙ�����'!���Ch���n����1`�<��?;~������Ϲ;����`yNkfJRD���B̵�je�m���a�ꃘ�w(��)J0!���@�ͥ.�h�˔����@l��Ƴ\�e��i�7O3�����pY�ڇJ}kR�����T���PV�a�3�v����gݬ�oG��R�����):�!5FwFF�}V����Rr|Uu��_Z�ō����@Ь�X��ε�r�Nj:fj��8UC`\:��մ�L_el����@9ˊ���DD�֢��BO���*D�
5=�d�0�W!�*�9`J������ʿ�t���Fū��
Ib~��O���wݝw�p�15Y/MW�.��/���eȰ�Xx.!:L,v���f �nҁ'oA�cwsh\�!jv�WI� �m��GfA4��?7�ʜ}� _@�>�}�Mj��(]��#5���31`]��,�*Y��/iV*��o=��x�x}�Y}���h/���[���Wm6��Cۢ�w�����u�l�;kZ�t�hJ�Ή�����+N���j�\�9�2��+���)��ҽ�C"ӧEN�)�3i����7R��X�i�ʌ2�Mh�Tk����%�Fe+�CH�M���L�"������݌�hMU%�#U��+���4��8�r�o!�E��-^���޽"�Lc�=qq��_ke�mы.�e�ì"imU��]�l
��VP�cM{Ǯ?�t�g�����ݧ����P��ov����Z� k��iJf���.V-�[a�V�C��EU��˦����0cS���X͸�K�v�Z�3Ƹ&7�C�ʗ8�|\�d*������f�ҝ�'d�h�9r���}W�;�2(�_Q�lZ�X�w�08މ[*k"-��tkS�s޵u��gu\�S3����zp��.V>w($+�j�4�M�4&�)uc��s..�v�i�\y(,��]8�z�i�K�P�.�x`�P�V�-H�R;��+������X��qoY�X2̪s�W�p�����3�շs���S.���=�B�Ar��/�����gR���4�ɷ0c2]ë0T��1�})D�7�mɪ�UP�x�:��E9.������yԂ=�s�V'��4���=�Wpn�ܫ�N.�ҧ2��͕��r���c�ڷSy`|`�B�;H�N��7�0g#�SɃ~��� /nD31+���WN124��Sk�[��V�oN�j����Bv	'�.��$)+ë6��A��T���ې�oX��OV�K���w����[s������7ۀ�M�a-��k�q\r�gK��ڎ�f�d�G	����z^-�s�G����IO
�A�t_����f� վ�Aͧ���gF�^q�E�F�fM�a\ۤ�hb��!����5������a�3��Sq���A�ER��.YmdЖ�/�kdS��}Vu�NM����J�r�*i�\uJ�3���B��,������k͍��>\lȏj���na���z���,��x{jRH'Gb���)Q��Ю�R�w�]���"��Q�hj�]/�܏��4
�Z,:P�k�Jv�t�>di��
��V��M�0+������PT�U���m�ќ�#I�MI��`,��00�gK	_T2��3O�є5����o�`�n���Vn}q�j��ٙԶw`)�c^� �+����g7���#fnVSr����(�w�@��)�v�4�3����ᨫm�Th��wo*YKz���[Q�+)�j��V�vN�;�	l�+�;d�cw���H[��A�*���ح�Cd�n�ы]a��L�y+Y;t���ؖ�N,���9�٫9��A	�] �
�uwFN���vR���m�S��^�J��u�Ff�Y),#	�J�dd"2i$���f��b�4TD�a.�q��9�b6��QAƄ�$��2
���I�,��j)Q	#%0�A�8یPA�!�e.8�h�j,�㒍Dɠ�#G9�h�1$���6��1H QhLf�Q%���b�&�(�Cb�s��1�ȉE2&�5%�h�Q8�"1���Q��ƍ��A���dhCThN+�X�"
��0@$��LbB60E�����L��"�1��mI�s(�8�32D��&#P��k
lR1����BB��К�i���^�믾�������\���^+����ĭ��bgQwWS�ުҕvGPS*(.r��e�/r�I+��j4�ʏ?�]Pp�9i[ˉ#?BN��|*��ɘ���:��B}�Wq�vGK��O^�+=���ݜ�ren�.+-2���F|��+�.8U(��&Z�=�P�kv-)	ೖEӧ;��AH���[d��\e�t�ʰ��6T���N�d�� U��fP���r;���aU�y�,���ݡ1�.�$u��u�$[~2�ױ]��:�Ƙ�	�����z��a�K��ܴ�k�Q��R�Ը��م(@.�ɞ1�9X[B��Y[�٩n;3��UU.�� F���J��I���E�ԴZ�D����v�S1�*�Ugua9���+1�*5�&�bԲ?\ WJ�
2*6:ֱ]jWB~��{I���`�\���W*Ҫ\0�]QN��β~�uR3i��s+�����DMu��	�CG^���KrY=-�cf�%�-u,uF4�y�*�2��|a�uӇ{ڦ�f��c���b(,}͜��̯]+?Ty�.3m[����Zg��՘���{'��@��6k��@���Q:hd�V�6.��+�c��p��(�{pH���ϒ@�m,*@�⡎�陃1�YZx.��N}e�:5ᾭw�K�2�ɝj�Sw�!��9hI��䳖���=4�j�H�W����N�C�:���ip�����]��`2��ZcU~{���jkmR���YHʣ�z*"�ku-X�����#��c9rT`�+���쿺�B��3Q��(1��)rQDE˄�ٲxK	}�K��ϋ�=��8�V*�J��#>vS	Z�ۚ�ي���W>Ig
{�w��0lخ�ep��XxFP�Q�F�nVD�?L�y
`*�����9#2a�c����[uH+3Q��@�*n6���	#�[q98����u�{u.æc�D��g!��9ˈ�I둽>�I�8!,X1jKa?{ۙ�r�mO_DO��f.����|LR�K���/@1��+E��5;p��1�3/���Z��p:��Y�r�HT˞bȋC�l�mě�[=�"|�,ũ9C��1�;�ˇE
لf���I[z�Ա�;w��^��!Ƶ�w��a]�«څ⍼�9Cc��x;�y	#(<���&lFk����窵�(:�r�����59���aΩZu����ʛ�!��W��k��}�R�<�k�D��qR����q8�U��m�t�"�r�7�qR���p�,��M�oAUU�B��O��q6r����ޢ���+QEV�E&Rch�$REQ���ޘA|���%uͅ,Ha*qw��������H���lw�ߎ��CG��)�)愧$�g6n�.�Qȯ��˕�Ias���e,���c�ݗ�7~� xt��<�q�&М������g�& 
�Έ�N]�a�}n�˵�(�ݣ�㑜����2�*r�W
`�ynSTh)�&\���3��!�����j:�~��b}�`��=5���X�zM�h���;y��u�����`s�t������Bʮ���.��l8�E�l�K6���	�k�5��_i:n�Wxʫ���<��Q��~�x��M)h{�I�L��j�bT���HT!ǟ�::�5��Y~G�w>/ܫ־�o�ԗå�1�&��R9��_ɛ�����T!7f
�
�{O
�t_0<%Y�̷K�����p䶎�/�ڿ��d�;>��]��f�]C�"V��W��VF�W��=�3×oZ<�O6�~�����ֹГ+��.��(d��슳�Dv٩ˋ\I���Q?��ĶU�Ԗ��v�k��F�P3<��L.��e�ϧf��{p�(�{��b�r�@�F��*��q^E�u�))�ܒ�΁�2b546X\�L֤^�j�7�9kLt����c/O�ZOz�����sCW]t��/R���X5�����&<2�2�9��7~��v.�x4���}pд�����gj�q��W2j�퍺���R��Yq`�bN {Js�y�u�-#�L�GV����b��V�+��l� ��åS_������R�(Wq�mdg?�K� h�?���Pb�?v%<Yu�0��ɸ��uY�x7&���K]W�mz��Ƒ�a�X	9��m�-�=غú�~�r߬��zU��S����w�V.7����u�A|���OH�చUK|��[h�o�::gv]}�/w;-�T��9�,m�'��;���+۪���
��;8pؗ���>6��c�CW�|�0u��\����E��%P��R�cy�/)�ׇӱi���(x,��b�@�CH����{_ɣL,��"�ffyW�&�YD\�&�m߈*m7���$��Y�ͯ
t< �T���վ����^\.L�����L�g�gI�o�[��ս��l��}�Y�@n��V8W�����[x�zbb�6Ǖ?f��}]IjW�6ͳ<!>���F�$gT:R-jWe{������:����[G�/n��sEo3w�2�4c��S�b��bTgtm���vjn���*=���̧oӥ��+��v���O'f���2���Z��D��r�C�p�iq�6mW�|%�_�ф�=1�C;f��-r���^�tcs{Wnv�&�ׯpp2a8��5�v��4��%��^-<�8N�Ɩh]&#q���{�����ol�����d�t��_.yS�T6�1kj�G�."�e����օ/u/eR�*����l1Hîd��먆���*�C����|���ٌ��NU:.X����s�~��ѱ異M��%��F��k�4#V���\���Xx-:L,7��}�gp��p�(�>xo~� ��ف� �q��P���㵷mq��S	������?.B�ރ��Mn^�W��p�%�M@�����x�^.Id'��Vg6q!�9m����n����e��v��f�rdg\v�C��W+�J<66ɖ�v]o�ݬn+sB��la��_����5�K����.��V�[��|���~o��O+� ����L��ɺ��\U��>�DQVVj��"�@����R�L6:Ò-�}3n�`F�\��A�1��&�j|������"dJc�@�{�������o
���w!di�α��u�;�璑cB�"���˕�w�MI\haTR��j��r�<7�����۝����%��:�H~ױ2�_`gD�v��̣�B������V�	"��E��ȆW37��!v'qdd�S���t	tU���wo;5Ū��A�'.7R�M�v*"����o�� ��ɫ��-F�͖�W�Vc�հ"���Y����_u��5��������K�x�}�����E��ҌZ�A��҄=�i��W[�uP����W���;A_+�	�p��uG����1β~?F�5 ���NT.���2��.�I6���k-Y��b��թټÔ���B�e����8|(�Y�Чg��@��3���'V��;����#��|,�FLd�v�c4����o/�OkT���0?��"�;�w/0�l2��Y�J! �`u�d��'E�I�����}p��G�`g�f���5v�s��T�uuԥ᫛�8=�&9�f��,%��������r|uu�*��2���l�[�7�ä86q+�Vd�ziـ�
�k+�`�<#5.`��Af�nV��VR�����v��p��s	�c�����P� f&cG��V����yp�I�rk���D���>N빇�O'{/�C�Q�̽M��;I�GK�Ğ��o����7l��acW-L�l,�u�S^��E�ƨ1���6�qB'�d:t��uL˫��f�l(�ƍ���W�C��1⭗�ZC<��96���:����^b�Қ컶���<s�C-��V�I!hC��3���s���}�Y��X�޾�g,���PZ�,���a��C9�6�-��C�.���f��x�����S��<�<<.)D��{`�X�gj��u	��W3�/�^7�P�p�6���u8g� 8;���c�S�<�{�^�������B���
�ZE{P�Q�9^=�QUo�	�D�kʤ�V�UN�f���0�K��D�RaU�h|�@��(s�3u�uHr�w�z_���޺���oԊ�9����t�@��9G��a�=J��Β���g��p�n�U��`��k�kq�ʩ��}bT�1�|~�H�K�3��`����-J��3��˪��h��s˕��x�U�a��s��aLr��>�Ѻ�L�-ә��>CM�����u0;��2�P��"�Q�k�����]\�:�B��.U&��a\$��b�fYu�;c�?7�r�ܪ�"5��ؓ���[�j�ƸV�bᲅ��ҏ��=}�鿳Wx�u��¨x"�3�"]���"�h���p�,�X�BJ��!P��Ɲ��5l����oqpS=�^����"c&���5�ҼY0��;!3s��|+o���Up��x&T6_0<W��I�ܞq�H��y�hi�,��ñ��*{�����?ez�cۈQ�C�t�s0�bl��+��׷�V\C�߯[��A:<`��1�N�lu�3��޻��V%��.dٻ:ʸ��:�M�9�t��rA�q�Ԓ����BsY�C�"�V�с	��� {��S��M�^��ٟ7ָT�I��l��d~�+d����H��v�	�KJ�ӡa�D>P����Ř�Z*����Y<�����IY\�ܩ��]<ޏ��n4��EĜ5�.��ʘ��dn��es\p1X~:j-+T��^9�֨�z�u��BC��\X�ܼ��=5ҍ9�/Ś!�;�e!�b�����=�6rb55�����5���-vaN�4���ݘ�Q#�mnn��y(�`�Z��<ZZH��VD�$>����dC�~�lt�ٮS��>�S�׹܊�.��K
C��e�P�^�Ƒ��j����F�Fŷ��u
錕8�˞̬��F,:��ek}���U�~lf�:�n��]�p��c�1(]i��XM*[��$jJ�e]u��'�U7y5�!�����&�N|(�BO%��ɞ���y�d���i;rE}k��N��֯_y�#Ԥx�3�t�Е��Z��� �l�˙���j�r*�G��M�������1i^�Q�P?5�bB����Ǹ�޻��4`J��sl��N�팸����L�(nc+�o�e&�]n�Fa8U�4�����De�/k��t���@��۝s�M��V�n��:]�\*
)�Ԕ�p�FvLʾ}z�Q��6�����nُ���e4I��N\���f��[˟��j=�{�� Ƶ{36=�+�{����ېs��f���Y�%%��c���0b\ܪ���
�rpl����;��YJ���m�^�!#���z �[<G��t���J�����13�7Cp!Gl!Ԩ��ش�����W���Yζ2�v�η''%�Wdgڙ����u8,�uC�"֥w)���ChCi	��;�fV��4k[W`��Z���Û��N��N��MQ�ё��[�S|�*��3k&�u^iP��5��BO��YE�$�nt��F�ܔ��N��v;��X�~��`�O#�Gے�_*�?<�Ib�Iz�:�o羑[W��WHr�0�s���:��u�t(�I%��;m�1���j�3����W��,�qU4#ak?+�eȸe��5{��`��Z�eZ���\+w�ا�V�t��"2�@�W��~7����ui@7�Э7�R��|L�Ӕ\�:�CJj����&c��0J�*�I��32��`�v����2"%wG�;�ӕ�5�M���+ݍR���RT���@���T)�n�a��6B�ǜ38X����-�:qc�E\"a��}a�łSh�6��:ہss0S����}���=~���WQ'�&�$��N�]��9��f�t`٘��fq�X�Ƭ�,��j��]�k�6��LJ��7�_E�����u7��_Y�jf��{��L��sc��B_ ��YT4�J���w6���N���@�uJk"PT�f�s*R��qkkw�3B���/E>D�g��������	�H���ɍ�zf\h[�zֵ�!w����C�D�d�FC�Vn���)7��n��R;��8���3��	=v��ם��rޮ/ |��A�q���}>�5ʼuP��5�z�g��p�F4YaR7�\d[�k���#�l�R7�����J<1jY ��ǁ�4�k�����]��4�ǉ��ܕ�m:�3���M�n��2�f����_���,m<�met7������~�̖��%Be������q��g&�s��.b�k2�Y�1r4"��]��1��^����Q��:N�%>�+��ue4:Td�OhL(͵ns���'_45f+.?e쭜�{�wLUt�Q�����=*���T��:nըy�j�*�[~�^��||M�bx࠼�b���:��i���Z&��<�`���M��ۉy��|ǹY��:|1ׅ*�E���ޞV���ӆq�4�a� �#��-���W�ĵ!y\������CQH&�7r\ �]�)+���]�rŐob��[�!hiJ\�i+��E���8Ue��$j��Q�1u�XvV��Z�5τצ�CVkMoB���)�	���yS۾68OP"�&M�5n-|c��Y���K��v�S�`N��ڂ�Uh�Q1��f�V72{T�r��d.��<�h+|��v�9M�w�l��z�]m�>�jS�o;�w4uƁ�6^�:\}s"�Y�YN�Jg
�r3��e��{���p�dÊ�]xj)��묛]�W%�(���T��'���xe9ӍJt���3@V�v&��Pw��� ����7�m�r�+�s7��I�iXh��vVM��:]7+�)�ܾ;�L��z-vu���Y���Vi�����c��v��wqf��`k©7���M�T���u��c��M&��IY87xprYh�ylL���U�H�}¶E��5�-"
T�]ov�{\ᩉ�j_J��&>T���,G�
,s\���xA�r����t��/�t�-Wn��!�dH궜��	�s2um��Wj���M�R������u��iؗ�ؑ�W���x[�{�m@�s��5⯥�u�q�z	�l*XxoE5���-�8�J�g����]�]�`�T�dCv,k�"\2�Vbeor��������Jg[�vH5�w%֭�#����7O�v��N��X���G�Mk{���z���f��v/�Z}*|��-�F#���'��������ٹ]TYO��	{T(p��E�m�1��M�o8+��:��X�QxS2�՗��DC.�vɧJ�z�V8�tvҦpЙ5�jp��#ͤ��"��'}��y��{LXҌ�N6򮠧d�\�GZ����μ�r_����o-&�lk%V��ړ~�/��j��N��A)`��0W+S�zZV6k"ǀw0�9.�sWT-��F�8Rr.��^]��q��H,��x���R)*s37-aH2��@��I��R$S=\\l�t1���J��f��;��ǳ�W���S�_hɤ*Y�ƺ	d��Lr��A���(WLʔ��/��?��CvR������������]�%��Q1�7��m�1���=F9ή����q��Χ���ի5�U&㑼|�����b����j�hsچ4h��d<����#B���,'ݙ���zwӂ��*���M��6_�Kۊ���85KOdŮJ���t��%oՂ.�r6�n��y�q���~T�|��R[7|5m;�vԝe���1�b���y2m˪�]6�>�.��-����1#�0���Aŭ�LsYڹc
!`�VB�D�\�n����)�M嵦#\b��eE��"�.v�DM��g2��u��Lw�˜�߮O��u����&&h�+�b�0,jL��$`��qqR�I�I�4`���1��ѱR�6��4Ph)�#%���J$��M�ID�C��K6(e!&�I9�f�14�DV�EI���
2F�FEs�ͣ&�IA&�7�b�r�I(��n8�RQF,DG�5ŊŸ������"��L�Ql�X���j1�&�hKb�j�AFJ�FK4PE#��M��Z6��q��M	d�M$��QIY4j1b�Fɢ�na��Ń(�1m4DZ4�l�mi1Lj0Wl�"�6�cF��d��Y61��I��8J(��U *�U�Ux
�K+\��r�&�1[��|&nZȅ�T��iۓd�O�]�F��Zn�Z��w���{�lmD9�*����֢�?<=�xx8�B��$����?;<��]1�h�8.F���+�u@�<%2��<|�d+�V��%-b���]�fy�~�0�YS�6;>�z=�EM4�m�2������\���2�(dHq���%�;O�qe]�(��J���9�u2󓿞��[=st8��
7�)N�VZyb��q'q��l,]w�ė���!�F��H������Oȭ�ɧ��n)�R]�'�mL�:4�!b�BAZ�s�2�"$'�1O���-WsDb�)\�3�i��GP��*��icf�=O�5��xő�dHJ����S�ox��B.���Z�GFEt��x�;yU�8��2`�f�7�{���C�wژ�9׆\!N]�k.��Yt�fO��V�N:{+�&y-��1�}�R�-��/);�	���s�Hxx���廢���q�v�X�7q�H�}.�μ���%���:���ҵF�.��K�Xȭu�kb�D��ё�P�j�͸s��-�j���.LCt�t59Fa��e�z4���+��fA.�Z��,f��cj�(�u!��A��܇�z	л�J�h\8l7x�Ŗ�b����>Ӻ�Lu�sdm2Y}.�"�L[:����������j(G�{�-����ǭe����^ k����=�����'I5y�GR���؜^wF��>
9Tl�ڹ�p��џ.fe�Y;c�{���ب��W)��;�ǫObW(֊о1xl������s;�M��(vW��1�u�dXMZ�;s�3��s*�oL��qV�jT�:��p�j�J������e���;qz�X��3#�zs�d�\aL8f�����uֻ�N���\h�k��W��t�vs�;�}P+�#o6w��)���tͤy�������-��(��-el���Z�ꡟ�f�o|�V���ħ�zt��6�̥���~���I�esu�l��p���J?�nF���G`<��Ƙ͘eP�۬ڻIR溔�=�c�hqH��D�/F};0���=�LE�4\�D2��V��n�uH� ��U�e ��*��J�
��B�+�aɚ:��pc��]K��i��n��wzW��_�J�����[�ou{m�僧��]@1���K9�K�8��/������tu�1��èS4�NNd.�[Cm#igk�ѓ�Y/y�O�(��c{W�Z�JH��̬I>�ďei�H�l�-�5P�j*h�ּ��˨Jɉ�n"�x�����߅��h��;�R��s�	���BosŴ�`J�T N�;�m3��u�+�F�I ×N2�3W�"87$���}��{�����S��ښ#�ϊ���Z��އ8�n�����qL}P�J&R?Mh�*�a�䥘��뙘��Up�$
$8wP�nB5\.���0�V�e�r�?6����qF @b:��5Y��4j�uֲ����$	t�D_]48�~s��F8�a�a6zC�Nfry����8����yԮX1�B�O]$=���x.����P�1�)��\��F���Eu9�w��8D��ܼ��m�{��	��J�U�S6�S�kr!���gת��czk��<�һ��T\�p��ܼۯ��͆�lO�u�Jqq�cp!Gl:��ش����8�Xp�7�<�ћ�����#S�hg[��D�1�P�YԪ�?s*��	�0˲���ƭ���P�갇�#�}3'��a� �خ��1���_[���3�n���Yrp9Ñ���%nQ�?���2������ )���-�x�|*v/w,���-M�����*c4�wv��й*4��*����閧%��^�9W!� �%I��������d���φz�ŽDU��Gn���W
̴�k���:����9��:;b�ͯA��8�����%��h�D���;*Q�n+#�SR������M��}��ͭV$A������5��n>�f�a��3�d茗MS�ԩt+<�|���mG,u;s�t���e�6��yi�������5R�s�������.F:���wV��V�[s ^�r�����i�(�h��'���l�W��a� ��ș#�D��Ҭ��]�*i��_O˥қQ�P��j��@�c�A�ЫO�:(�$|��׳��6T��"-���<�틬�O���������뭦H�P��=}>�-�~�Tp�h���69)��z1>��L�85�v+��ӉHl#|ޖ`��!�`NR�̿w�Y��@4���<�R��b(Lo���&R��62a�s�c5�w�[}�m.�
�`R�1H
ڤ$	^;��1��F�b{�|o,S��}��j�Z�Ad���
��-n����_�����ܧ$��C
)V�}C]�K�x ���۫��}W[Fg#��Yd�i�#��0Z�c0W�w��k����5@����LZ�@6�p
�B<��d���]j��9�S�9����ag����SɓSЃ�uE:s4:���[@���u�U�atNm���\�^R�[�S6{�)�I��s������'%ܧ7�]P4����!�xnݷ��V7ϨҬ�,�C�`k�N�`}o����5�f7�%F���/� s%\Ev���Vc���u�/N��/�EcŪ��t���^����Vu�vF�ޚ�}��� j��EN[��Û��s��e����15��50�d���/&��n�ZP�FOh�ڇ�p�*c&.s���}nD�v�3�B�j�V%�zn�#P�k!��k��%P��>*���ҡs����aCϒ�J����Ȥy��q[q��0�PA#�dW�d����hg5J���K�m��j�m9�8+b�fZ0�;���:�^�L?����ϝ���5���6`6]P��uEp�L��PSJ������خ]�����p�7/43��Y,��N���K��j�4������e���[��Qyǝ���[������?"��O7{9���\c3/m;��5���8 Z�=�:���SĜ�$}'��~:Z!u�SOk��4^��1p�Z-���$Xꬣ�kab6���sZF���fw�b����T9��b������֑���\a4�-��f8����"����t�S��F�� E-�4�^d��a]�¯�5�_f���ݥȇ��F��;[/ t�J���������·�9�pO����N!��ʹ2��8s�R�uz�ެzz��P����񴵷�p1
N@�UX�+	L�p,̝�u|I�ԥ��}�j��u���+6ӘvN� [�ڹYy�8Wd�����xx{�M12�)t��E�j U[�U��X�]�:7<ߊ�#܂?u�D*G}����a��݅�3�fSYEr��k3�u���Z��K�AȜ`+`�
�Ep@f�U��Am���*�ڸ�e��;֠H��W!�.�+��#�J�D�s:�P]�DR��竁͈a�&[��B���Yc�A-�����T�W[���c���-�j��L�0�9��s/$>[\���6�r�$;�:!�����c�1�Aa�j����t��J���u���C�32˨9v`kF�tA�j(r�}\���J㸕�5�Z�l��J?kf�Ngx�>?`;��2v�m���QT��y?�GX[��_�sAB,�P-jB���:;"B�5�����Ʃ�틫�L���.W/�e\9�B���i�MPR��a𫴶�W^]z�A����qb����I]�fg���3Q|���ϊN������U�`�Y['��8�������y��m���Ꮛ����0h�3-dO;����%esu�������s�V~Yx)�1�!����];�S�2���E:ۃ2�nZ���:�5�l�0�T�֖ۗ�t<�LCdR�����ލ�7e��t��S�T�D��Z��r�n��
��������O$t"�����Z�N!�|�9�˴�q�_��������rg:��bY�R���ky�����)��DO2�F�9v���b��&��>�L�U<uz{
.�8���*_Xr*��D�0��!z�0������]��<�{�NC<е���S	>���:��� �����Q<�¯��H}-'�S��(�n�Ť��7�7.�_S��M��]�9���l}o�Q�lx�Z��9��a���M0n�9�W5md�u�PS\�Nִ+���Ӏtvϧ�Z�t;�1)}!��y�E}�e"65P9zҹqIh���e�(�>:����zt�	4����p��.�㴔�9�p1'L�Ϗ���"�]K��#�3�kCO.a7�Է�6�k�ٞ��]�����1ת��2�[ʱ=�\4���ھ�<w	�:�^U�=t�̻�b]��uƦ�7��N�_wUBv:����o�}�W�qaEhg���;ǖ�i�����o	ׂ�xj���k�j��{�V\�jZ�Y�A�T��h���,ckA;��:�=Li����ִ�ieB��=�}�b��.{����l'k*���x3׃'J\h���Ph{�ұj֞�\��6a��V��c0$���y����n�-��.���g-�������C��Q�t�#��#��^���N��Gp�H=X�-��2��1Na����ֱ�n2(e�;��b�V���9��4� *x�x�4wt�Ż32��j�US��[�Vm��i8u+x���Nz��Q|����77�m�[�8�fP���&Z#7S���m�0T�!]H�1Z�1�CW?N7%$�杇�k6���:jOT�M~���q�Y:�=�X}��=�J�Zʂ�%�w����]sZ�YꔣU��On��;lq*gj (/��]Ob�>�`���:Vܥ܇8g�|����C�z�y4�*u}�g����qQ���d>�O�*�'�����+Ջ�^;}8�[&VLĭ}���	U���:L?�7�Τ�!����hc���e�� ԙ�r+r���|{��	u�t9!-�<�7�b�&���?{���)L��GZN���|I5mrx1��u�F�Ӷ��$Äw��+uMZ�8TH�:p����-�Q�H���-�-]z�/Ku�B��@�W;/��
j�LE��b���l(-l�d���W5������z�p�2�.jm���wr��:�UW��Jy/M���s.}˶
����i#� '�Ի3x&^�횹[�S�|���/;9��5*��.�ȤP�v�s?O]@Z��]�
��v��kVcU�9l�o�?$����!q���S�6�˵Y�=wʙ����v�Uտ�׵��m\�:�m��;��x&�\��Z����yHm*�G�,��Xz�\�i��a�+_g��oh����p�[�]�f�1&���P�6$�q�-�q����)d���^�v<c!=i�C���4Vn�Uǃm����Şs�C��,�����VE���Aw�������S=[�4��q�����m���sWQ7�k��Au{�SŌXޤ���;F��Y.֤wc���K���}qK�mgW׶0�R��WR5��geE��я��fsKh6z9_�Y-�,��6�֬���:���C٘��E�B�G���3[a�I]��X��5,�ּl�SY}lI��	3M��@B. h�S�����7[;w���.���G�`y�.�ӻ����rY��u�n]Ub��gN�ɗ�je���Ә�Ν���X�li��.k$p?ʪ���c��8�j��"��u�HJE\D�y=����L&������fL�܊M�.��e8ۙ�
�f+i%���a��-;֥���쭂䨠�ܜy;�ؚFtk��}*���@�Iɉԕ�ӝp��?:}³3`���"�1gzs+-�9�!c]!P��ﻨ9��oBk3�7���L�dZ6Ů=��*��J��'7�/�^䟓s����1Iٞ}[��5�p���Ж�9KUQ���zt�%�9}-1�U��P�(nD�bm�n;a��9A�q�2L�t��i���>R�'�I˸���qIؘ�MY�
��5(����Ir/a����=�՜�����q�z��v��:�|����r�}�Y�h��R�~��9��ϻ��VT��C����l�5���]g��/�Y�V��s��y��x��!�ᮕ�����vf=�[,���C�M��-Xvx�ۭ��v���ZCojy���,�h@��{U3v��D�\��%ݍWq]9��\��;0�w/dn�]��H�7��A�}�h��Q�	<���.5H-XS�N���e_V�q�J�����ԙ���[�K���:74�ʾ��9�n���ˡr�Øle]���<V��]%��vT�E�qm��b�˕}��H[������/<���{r0�p�z���jΎ{��a=yh4uw�7Ɏ�r�u�D]�-��6[�qƐ.R�Tg6
��gv�U=���|;�Y�=Gq��wk[:��^lm�Aѫ֮T��k�6�G]mQ�U���+M썌�sh&�].T̀Z�_8�X�yg��j	���g������bf�2�����XH�_I�����í��*7uq�CfԾ�i�`�*�PN����נ�-�׵j�4UM�9S3�^'X���ǭ�䈺4�ov��:�+�UwۗE��N��\uztcm�rȋ0��]�]t�/G5�ǭ�
<�����p-Z�$�1:Qu���Y��.ͫa�����:�+�}�e� A�����زfl�f�>���s/��⳶�ZFK���0 ��`�B�Gc�&Y�2i-6_9F�N1��J����	[�s�m��䩣#��z�;��#��\�Z�h�	�`Q�h]L�2q,�VS�%T�h�:a��B�c�vql̂��-��륉e���1m7N8��ov^%�X#-ְ Uc��[������9�����ӽ�,{�1�:B�L��Fq��q��˼��|��Սb���nK�5��n�ə�jf�m�Z5� ��j�[��73�`�k�*�݋c��s� w54i;�Mh�U��'�[��jgj�M���4 \,�@SAа�K��َ�l��uS̛��x'j����<�8Ǝ�]�8˻����U��ZZ/(�[�h?&�K��6����m�<����h���~|���V��S���do/yDr����U��5�r�j	u)y̖7��:����0+c3�HGF&��fk�VaR(�TB�1
c��}*#�����O���z���==6���T7(4{w[�]r#�Q��5b�4d"�Y���s�v5����r�s7���右��3�:�v��S�z�X7�5�1,G�#N���b۠��Ӷ�tt�����qʖ���N�/����7"͍n
�d_N`�F73�4��������4�v�w�!=�wGb�u#����v��݅Ŋ�[�s�:dc�W�k�pL��(։�_1�+q^;��it��L����#+��eJwV:��fS�ocBp�
����n;Sk���n��-�E���ڥ���Nq�C��"�*�5h��]�햖r��v�[0ǉn�.KRL�V�\�u*��1^Z{\r>DS��
��l2�2Ob5]�^ɢW��� 4i(��"�F1ƌ_˓����@%h�c&DL��4�IQ&�EE���j��##Q�+Ʒ�Pc,	�5J4QQhؒ1�cAEa*H5�LDTRTn5�	Nr�(�X#A����4\\UDD�,��+E�QE��6-D�ƃTPF����Ƣ$��ب���&ش��4&�	�(�2�F�j��ذm3	Eb,X��F-E�1E&�X��F��F"1d�!*Li(����I�F�,ci+a��D�E%	��X�Q��f�]j,����L��Z]
8]���CJ�˲��i���(�TGn'�J�;�u)����,�f_N�v�t�g�".��9�oN�J���Z��e�"��x�����쪴�j�➢7ƝLu�^Mqgh��V�����q'qC�{֫ڽ;ؓ�e���Z[C���b��7��k��WXbk���(�\�\Զ[�]�k6�leudP}ST�I�����_��q�,�/��W�<��7&!g7��i�\��k��<��ay�^iX�L����i�G�Ҡ#��U�N���[���f��֕b��F8f�a��X���?W׷2u۾����{I4h7N���S|g����JoNu	�{�w��m���=_wϪ���1��Ύ�kV#!_`S�\pOav���<��o����\f�b��I�*�ﻨ9S��c�b&6*n��5.u��C9k��tҸ�3^��=��4�b�BVYB�ج���F�S�ς�^ؠdǞ�S����N��Q�K���%�����PW�FV��t�3�9��. �zC`��[E�뮕��B�۵$3h�W������X=1�8<A;xk���׊g��-����r����8q�/��@��b�ˌX��^��-;Qƥ�n����7��p��6l���%J�D�Xk���ئ�G�nFӎ�Mf�!c"{�vD��q]�ܚֆ���&�X��Qu{N�K��Ѭ.�3�Ҍj�0�E�\�k�	�믂ܣy�_rҹ�藏�LIU��M����K��6�]�����)��ml2�]�F��M&Ŏ݄k�k��}��UgZf��l��p��x�io	�x,���mtf+b��y!�:�<��y����~���-�>ԩ�����)ʞ �Ժ��}�`����Z���]���U����r�TTi�@T��֮;���2LT���FF\�'a�|l����.yWY9�QQ|������;[kN�����K�S���-4Wժ�����
�F�d��j�8G���lE�%w��n�VC|��;歞ݸw��Cm���P9؏�.��:�7k�[�y��,���������M>�e=��(F�o�B���j�0.��Y��%^՜�s|(e��b�>a�]\�x/�-�n�M�fxpgF��\��LA����Xje���.��"W;ݮ�!Mpvנ¥i+�����M��s�}D�R���1�\��-�^<�V�$~��2#Y�#����(�٧���Eg���Q�Y�7ښ��C�i�˛��կ��)��FL�Ds��g7�����}}���v�UNh�mr�e��'�����o�
��Ϥ�q(�1N��i\��>����d��Y�gb|{��1���{,��3�=�[�	v�s�0��p���Y.G�-��s�Cx�ޝ0�J�^ѓ3
�)1��D�M��V�1�%'�a�
evD�G����]��pOu	9� V^��M����2u��?6�]��Y�
��x�u���p�?d�:����|�e�ݮ���KK�,���NCn1��s����敇�5�1����r�8��%��ˌ-mf��W�8t~��N��ׂf�yw.�ڑNAym��%�&�3�S��z��y�6�*z�ǲw�����O�E�H��yu�ꐂݕg�ڴ�~��VV�����������ߐ�&D���}�4Ǘ����t4I�R���7�}2�;�5 �ռ��}շ|�12��t����C+pCf���Hz�~�K�#U�g�q1��8;�j2�eL�]��c3W��=����I��:}Y7��j�&�]��Kڈe�ض4�E��8f��#�F8`�I�ۼ�6F~9�г��0<r�.�8��'��]BW�|kU��tC����t��|�>mn�fջc�sv���U�����s`X(n�I��mE����bq90�77�)����|p��/Ts5Q��[��"�����qN�:z�t�r~Y-e��}l���k�ȏ��dEW�d:/��%v}C�$r:k��G]��R�n�JV�=0�z�V)R��{8?[y�כHo�@��"_!�%�+!�{[��Ե�G�++O^�����<l[��yru�cΚ2g���@�IɝI_�Nr����W:�7�w�C��)���N^s�nsL<c:B��]�u@r[;)�xҠ�Dj0����ifco�[���֔Kܒ��a��	\~�H�ʀ��C�M\g6��p�Kq����\�����[��r�ᇒ�� $w.���vX�M�nݳ��	�91Go�$V���s�X��s�1�����w\�9��4�j���i4��%�~��݉����k��W	�Y\�-ɼ�i�D�vWf��O�:h�K׫�M��B�N�W1�.V��>Y܎ʝ"(�?��aIu�}�23�M�D���o�2�K0�y'.��!qx��=�::3���<��e�}����t�\a�q�J��D� b�;�.ƫ���}���0�K��Vl��~µ�����gx8�r�mL�:�i���J��1��`�F�ꈛ]�b����l�Gڛ����Mo��v!���];z_Nu.����Er �F��0�.��E�8C��ΥQN�/K[�:�/���$�*��!�}i��e��gZD��sn�l-����g��^���U�����E��:�n]7�nbI��Y��.����ywc�Ѕ��9���c]�J��'YQ��B�op��~�hU�V^��c%n��q�熼l�`���΢G#iшҠ"�#8�k��ჸ��[��*�r��/9r����=q�gh(/��I<�VC��
��ݓY~�@v����ih��5)�j��\պd�IweHc
�f��-33.hnb�NI��3���t��9%g����8T�4��&�[��=��3c�TQ��,Ҳf��j{w�
L+\��!N������*m���&�3���ԻS���}-b��M�[(�����:�n��~��Zػ�&XYn1'ݕ�j��/�[���vF��?<axw:�����������u��U,;�1:��C9k�a�8c5�{��mΟ�0�[)M�gD���̛y���T��=��s��F��I�r�K����R^.+��d
ܮ8�'��_�,vD�(ٰ�ю+��;�0�N���\N82`�aN�b�R���ԧ-�u���x	��X�o�k7��$��y[���rW)]�U^c�4B����k����=do���uCӚ۱��g�d>X�o5V^�Uӆ�K�k���N0����vF��\�_�u�����7رլ������p�>���5�|F�s*x���-B����QM����,�s���'/��|<c֭�������Lܖ$�<U�/V��#j��q������T��"1��[O:�GGr��_�1�<_���r�����˿��l�Y\�a�R��1d�lgGv�����4��Oy���Y���D��h��]���"i��Hl�}[9c����KCx�z�f���ݶ��s��T�}ih�ʾ�����V��Ξ��s�.��ށoc�E�O.�8mo_^�׶0�/%�F����t�j�C��6���ʰ�G	Ύ	���Ms�v�uٛ��,���U�����*�G o��R*wηyw�i?�u91n��O��d/nC���� �a���,GAG�s�_��4��:�#�$B�����e�Bi��-��FܕW�bi��wj4��3�_�ع֒����a�y|���q�o��p��:���V�Y�W�����ָ�*�>�A���L�5��q����}�O��v�c�s��NE���W�t���r %�cB�s�oN�[���û{�h���;JXv�ļֱ��?6�c��餏ӳ)�\q]��M0��ybڻ��gN&pc��t��0[}.�w�\gݼ�j���+�odH����'���E�/��%<]����ʛ�>uٺ���+|�\�X=����q�ȁ��j�ep.�)��[�+T�,9��'������E���[K�A�sO_AҮ�A�7zN�[93|�H$�<%jU��5��qd�u��B�7�0���u�����1�垩<��zY�> ���ۍv��Dk�5�D��<���ow��!2yNR��w�4�����Ҹڿ�2,p��t�<2���ͳɚQY�54��N9�����K0��k��zoM���������u+�D�tPk�,�� �G��:�k>�;j�.��=b��y�}�Im��^���Szyu%�Z�9��.m�ו�,���wS�F�V���s)��O[��s�MOg����>]aW7.��6��#�j݌1�sWV��:�B�n�J�]ϖw���8�����~����S�۷:�¥��lH�jLS���ׯ���?���z��2����j�6��<�t��M>�Ȱ�6�����|������^�u�J�(����o/=����B��ӝP\���G7X;�L�r�ꀾ|����d3���i�ˁW�n�\��w�#G^8z"�Z����<<�۔�f#ovʲ6�UȖ\�)igtj�I=�C,��Qs����.,I��I��x����a9Ω��|���)3&�]pn��ő쭶��\b���Ժ]�K���������H���r�����5Q�,�%� ��i��1�L�wϨ(��:�����^c��N�vR6�f�]��������s�a�]!HJ�ﻪ����a���P��SZ�*����{��T�sz҈��%�0æ���srb}:c��S���.�zl�j���zt��9}-D�r�!���P��%�
�E`8�xҵ:���]��j�3���c�rḶ���v�]JΣ;���<E�z�X�j�psH�-�xS���ӽ���ث|؛f8��Zٮi�n7�î����g�Y��>G�{۾qSJ�7��p�;p�åC�[�c�1�z��M�K��^�
���yR3}]�{�����zS��rq�g���Ϲس�sN鷘���VD�+X6�ZX����7�/��AƝ�U��D3�����؋v2\Q�t����l(��NɅ�;�}x���g���,��h��!{������=�j:'3/Wu�4W��5�����l�˂�sj9F�
�@�a���������Xθ�fu]�2� `�ǋ�N��	�N-�
S��E^����r�N���s%fp��4�r�7q�3�s��sk��[y��^|���I��[�1%�=!ݩ��v�yص�][��q�+��qZ�:Uw��x���k����3I�o���Ƭ�c܏k�q��=	}�v�Oe���Ҡ"��!,�d���1&t,�9����-9痍><��d�WܦvT|��i&T]ˮBzhTU�\��;	�!͞4cZ{p�Zیp��� �bL�}�9���n��!#��J�9���`����M��-�����ix�t��L�QgM���<ु����`ȁ��gRY��q������Ŏ�m��J�oGb��N�]ma޾k88B]|�J6O�9m+���ޝ?$ҹo��;�]�*��s�4�v�9-�˗�>�E���?NȀ�ш�j��0�N�̪[�{�3Zͼ�x�=����*����p��r%8Ңܣy�8�X��s�f��[���z]���C&�ޜb3ɰ�����U"�0#�mM[yP�����5P����3�R�0dμ��jL�c0�Ee�[y��ܝ"s�guan��|4f_d������i
`盡�̗u{�6:�w2�n�Y�	�z�n��ep��j
�5�PB8�K��K�J�K/$ugw�K���H�Kw����ԻB�\�ԩr�אz	�2%�K��;P
�6�b#bw�f��T1(8�W6�(�TR��f��C#��wY�sm�2B�/�����	A��9_WV�|��!R�d��?m�O2���0(�R�K���}�Do��m�I����c*�_l#�����m�y�@��� ��!��b��]��h$���(���]��rY�%np�Y���0�x�OkGP]�,]p��axE�;2�(�XD�M���2V��5|@a�����]zn�V�^f�n�(�a���a>�
�h�ź�IY;��v��Hd�r�5p��qQn��.t�+��_,n��!Z����#r�ho�qW,'WV��nt��B�������c-*��3��,ƕ�϶����m��W��c|m��fJ�QΔ�axD|J���+�a]�,P��nb�o��\·��E����$b%��E\�M�ڦ��Ȩ �.�-5,[,�ͱy�m�<�-��Oc��*Z���R�k��,%)H&+	����	�8����Z�R�T�C�gv@����g�a��j^G�	n8j/��{m�5/r����']��E����:#�sGG'�# .['9��Ww#��۶%ǐ�{�[���Bb��+z=9}����'�
���x�P�����{�Lj�m����-�gX*hƆi�գ������O�[�y2�ɢ�7�v�fåƂQ���+���=v+aiє�_I�ou�����0�>�9��s�Wd<�ں��!��n��]g
V���C9	���7;�{3�i��������*�Y�ڭ�k-)�+��F�����ݽ�r�Y��Y�Ǩͨ4��gcZ�+�h$Òb��u�:�[���*v����L,�����Ht�D�����RG��0�Q�rc��dd �Ֆm*m%:jq^��eҺ�[���}G)řj�ǳx��H�#����1M[Rv^1yԏ��8��9���� �ӴD&��O�,oK6��Wsr�G9�9T��ڸ��@�!.Y:*�Q-�֞Z+H�n��Y�����*ws�(�*A�L��k��YV��^ۑ�cJvN����9�{Jhƴ\�hp�,i���;8M<�����.Do8�,��Pqe�N��w���su��:M�J�V.������W$�B�6�"�e�<wU�_t���o\\������d]@e\��:���JjfV-z��:ѝ�Wh���Ha#y��e��x�)6Ų�6���@�CV5+�Bؔ/8K��
��ب(�6�F��&h�F6	6(�Q�Q)�%h�ch��&�2`�c��h(b� �Ɖ�� �J�HH��5�ō��lmE�"� �I�-�5����"���)6�h�cF�������-�����Z*J�EQ����6�ĚZ4Q��EPCDV���b���#b(�R[��i�V��ѱ��Tlh���Ab��,PQ��ld؈��F�X�B�&6,PZ ޾����=r��Ͽ�>���{��~��5��
���p�Gt�
�N�q��ּ{�~b��SW��a^�O2#���R
�x���ӎ湚w�	�&��bsF!���f�Q�z-nDK�qf�%�1�\��1W,�n��q���6��;k\:10�v}�d�)%%��ۍ{^׼|7���Yl<��/gn#5=�/a*}k\kO�geѬV�[qH���k.f��rkj�qә<�s��U��(Pq�qS�3����\w����V�9ɫB����Ջ<�0�Qo5��6�U7�p=���N���������y��NF�P���[[��G�5�K<ˬ}^���`�����ױ�"^����ysg�m�U�0z���[�jg���O�ѹ�NY���V��u�?[���M>t�p;]�8�TΡ=����w=��!}�5�����{!�HF!h�oo���\C�zSOnk2̽���Q���$�I\�3<���������C0��.�����ٮ3l)Uc��v-z�����Q .�o�X8J�e��flƕ�br]��]�H�CZs�f�(uͻ�IٚfE�uw9t�P��e��E��(���^�jo7�@�t�)����čU͒krf3�g6��o��CZT¹ُY3���^�oWo@��4+��	M�IE���h�&z���|�٫sܕpSy�f����%H�q�Q;���i��XƗHR�;���%�~й�!�B�U�M�d>B&y6�|����o���o̓��;b�	\bi#�쀟T)AH)I��/��e�oQ���zt��6�Z�1˸C"�5�v�s�#qV}�5S�8�4��Id�������r�->���rq����v&.�peȵb^�
�n��z����zۗI�vjҸھL��sn'rݘ���6�oݛո�~3�%꜅�WK�g��iM�<��M���|^���6���uzC�k.�^s5�bDg�X�Sy|�֗ma�߰r�j>�3xL��C����y��cVg.��h[�����v��+f��b2ㄝ2'=��N��u�Z�=��X���W79�8��]��vmE�b;֕���>�bQ�5K(dk}X}s!�]���ɬ�&2V������������U&eB�b��k=�ʍ�nu�	���*]��Q��P<N@q6\���D��&�Y*��F��3g�C���L�{j$P6���Ss�}Cj��H���s.� j,�f.�NË�J��q�'�	ssl�֏n����ܺ*����:{+�ղxݥ�9V'�+i��	\he\�r~Y-bi�y�>��x�_"��y����Z+���9�]GIx���=��O�#L�<�n-��n��}l��K;�$�W)���|���+!�^�v+�)a�y�7��u�r���Za�0�(����%'&'RWE��5=���-�ԻVj��p�_csx�p�
�%w�����d�l�}"Ņ�4�Ը��b�固�4��k"%�I����*�	��w�զ~����t*۲�z���U���=��	sP�KR�ʶ.2E�{Y���+!�$�C�B���v�-tb�������y'.kl���lC�ګ�u��J1��p��s~����2�=��J���~�1]�)��P}5Y;=C���,Ֆ�3~�M[�0e4q��A�6�0��Y��5�i�^W֐A4�(qw��ŠP�]�ڰ�����pYu2]�25mL��
�8(9ԁk���^�&*ۍT����̓����U�J�&�e�'�.n,a]ds�ݳD�J�͸�p���9�[{")�µ�4N�M�����5��D�L�m�w�\:0��)a:�Y�=�'1S��_D�l�QV�$�Apιۈ�h���p;<��ާ�~�r�Y��_ZN�!<W�Z��/_3�H���8����>��M9C���>�L���{1*n�c�J'�)Vok�<᪏+��)U@���Z��."�nno�0#b�M"_�?y���ν#2
�ҍ��b��cJ����账]3���3w]���e�W�{��ro�����k�Q�>��vg'�7`��o�ֹ}ض[��>����w�$�W)��%�� �[Ǝꚽ��O���d'N�Rx�K[q����l�D���SN4�l�uT+����{������gZKj�2�����X�dk���0�*��'�ֻ���UN�3��h�xX����9&���V>�N:!�m��y0�+խ�HR�Q�͓��C��Y�3�ؼ�Z���#pv�b���֖���,L-F����=�Odr�!/����ا�::�s�iTH�4�\�%A���:��q���f�̄������|f
�����J�)����M+�3^�����)�gIU����⋣���N��H)��ٞ{WW=�5�:Ri$�|Kk93��ƥ8bԤ�aBq�����Z��]�q���oVlN,�,+� ��������O�)��r�c�.)G)ډ	��-ʶ;wcq�A�LP�,fb��WVS����j�|�9�ۍwUk�:�s��ؑ��	����-)C�[�k>�o9�>{�M*�3�\:0����v�3͛����k ֻM^�.Ndf0�������^�i�\kY��Za��@���oe�iv&�����-�%�|�`�h�j��>
�1dĭ�W���]N��6wt��}�s�]DK�~��?M&6ꑠ8�V���@��wd�>��Wi�jwHayE�����߇���?hwN����h���T�9Y�g����hc�O�ֺp�/EDE�nj�̻jwA�M���k����A��81̹�R��K��5ְ�Puε/�?=W��Jإ�����^�A��Z����czy����v��ʏ5���Zs �$�����gɎmc�\���;�mE�c���NL$��v�����������b���D�9�[��]���֩�J��z?-e_ӭ͸n�O��S�������N��o\�[��x��ہ�>���Mu;��	R�\�7��=��	����d)w�H��5$k�I��ٞ�{�3��9��̽��ˎ��L�e�$�
gݗ��i��U��wzֺhɕ]��
��~���Z��F�Nv��2d�a��l�rC5j˝�V�oݐTߟ�e��;�$��~�!��U��Y�ķt�K/6�[i(���1�%��]�HJ�IF�ƢT(�c&@|���w4n���w!�>R�o��C婸T��N��ů����6������#Mܤ�,�ھ�s�a> ��r6�]����`J�,��opl3������v���7�}���Wf�]Eo'�yz���������r�Z�Yr'�Z,��lb�e���=N��׵�]&+U�9���:�R
�_#�%ط�j���:��Θ4ty��X��t��*z���Ι��2�'e�����*��"�E�n�d�MK���U؝ұp汻N�Xkm�r`�yQ��B��t��o�>[��[����{�ZSk<�����練Y�Ч$u�Td:S܄�=h�]
�����TF�c�D�3w�{r��zۺt�_@!�9�Z�ލ���A��r�����\�0�wS�S�1W��e�:��Tuj�(����=D�Ev.r�7+�g6�z;6���2^�h@[���oe�I�쁴��[�����D�CW8��ra.n]'�����m�(���ת�i���֞������	^�Tcs�%����WkzKº���N��uo0v�ݱ��.gh'R95�cIx�눖�nWGK+��z�m���|ۇ�4���1&z�L�@P>�Nwt��u^�!g6���=��J}݅T��]+���Z^p���g��}A@�I��squ\N�Fk}�X���2�����V�q��/����%W��r�������'��]謂��z���J��V�D��܎ゑ�L���O����U�R2e;�ŝK\hXIV_D�}��cKw�)ɚ��c���]ˬ�Z����^�����	UY��]�kv�q��iݎU��z�J���s�S�F�eh�s�/��^�=�W�{��TҸc5���%�0�`��n^=quF��]�o)��\�Ϩ�q\�Ki�N���o��v�_I4	��)��{5�z��Y���
�i�	ƛ��ы+��;�|���-`���L����K+�Jr�g)0���v%mĻ������j�5l�����.��j��h��sn5�q���B���T'c5�]�b�����	G(����w�n���-7�ե㶵ã��m�Y�8j����#��;o;w��M�-uoq��ME��(;I�.z����d���%Y�=]���RS�,�ŕu�('9}�(�N�*��"��	�ڑ�*>�1�<\�]�o�٧�HCڝilu/����J^���.�n`f�2P����#�u�O�nm�N^�V��T�̺���-�^�Jזֱ/���YJ����,���{+6%3��/o�#����ˑHGKk)P*�ȧzyprZ��f����c�}p�Z��^�;��
��"���Gܣ���c��.��i�>��V0ѵ�˃6XO��w9]˯���5�5գ/p"� G-S8lk���7#�6�w�-5�rM[<��r>�w��בc]���r�>�id�5MzABz���վ�5��z�����I���3�L����ۘ�"Uf�5���u��!��f����K[q����l��g�B�{�K�.�!��}��\	Ɓ�i-�|����[��Ԟח�ǦOa%��ﺽ�q��r�L�ϵT���o5}�!����ΚV�~c��+��q;���S��������L)�q�%S� s��\�CQ��:�gOH]�Ѹb�>([`f;N�o�D�Ҝ�:��.�R�dHH�Ȉ]+�����.�V�7gM�pc�>�-s!7��%��!p�q�v�Bg��-v��w���,Նm�k��uZ�w=0�㿓D����k�*�]���;�����WW4&�v�0�=9?U�6��,�씟=\m\G&uk�K��u6j�D�����P��Qy |8U�cW�FҎL�\`���#|;@�/��K����V����.Qiẜ}�)��A�i�]��Qljq{ڞ�5�/8�#�&�^��\��c�ۀp��JZE6�j%�x.c��&������@Y�N�%�[�sA�wr
K~���m}y�<����ی��h��*z��>�*��b:}~��T8V	�=���wW��B*��jޟ�,����ƜќWѭ�'u,�x�lUj֯`'�[Gv���-س�s�\>Yu�&��B�jNi�}{�Ͻ�T�/�~�=���wH~�^FR�y\N�l�w:�W�4�D����ƗmʎW#�Ʉ�{�C�ճ۷^��Co��`́�x���N�|<���#��N��z0��q:ܘ���i�����;�v;"��8��r�K,&ng*��m��u�Eh�.o_KV������`
���o�c�G7_��1&UG9�����c;����2��N�\,�#;��ϻ;T���t�԰��W�=-mu%*�}P��L�5��t]�C��c��i+����
�뷮�������u��}�r�~�C��G���.�cx ���f۴�"�����hm�:�ʗLΛ�T�w��V_Yo��@tf)o4��@���]�|^���m�w;�c'R�3(��
J��]}T{���k�RU��e���^$���er�¥ݥ�`�!�tꋱt���t�Wgko;��F��a>7������T��o{;A^�S���������wd�z09j�)�R��p���m��\�-�#��\����wDQ4���j�z��Gh��-�&�ge�����b��EC�5�;�'Eq$�#�h`��e;v*ȋ_��-�q�o6��_QG��f�5=���(���tKc�s.�VP��d��	�f���N��U�d�Wju�k��oF �zV���&caY�g;��-V{���Cɕb�dgn�t#w�ea4ճ<��ЂA�/��h���)n���k�,]E�K,(6��ހw�WP�U�>�/0e��q���)mͭ��aC�1��.��n��x.��+5��s�P�X+�p�z���+��=<:�%/*gB��G	�È���+�95s8L��t$����A+c�F�ν����SyӼY$�r� �`j���9r�{�1Q�p�r�+"�N��]��;`U�q���9�	ŷ��t�ю�����gi�ZV��o�L��J�Q1�0���+W-���������(�ӡW0v�N��Kt���+���N�mP��hգ��XM��wZ3��l9ƻT���Ly�<�,����>"f�A���ĴP̎+3���5��%"$�V-���fo=a�a�����4B�:x�e��Z�\��B�*nA�n,�Z�YǑV�&��-�'�����&�n�t�$�rZ�*��9�L4v�!�Z��1r���	��L��ؕݲ��s��w6V���ad���ۏ0������D<��W.��a�A���2�q'!�7�i�c5t)n;���I�L\Y�^wP%돜�/��[�j���<j��ͥf|�,,��U�]]��4�Uܺ��(�e"�e����3��A,m-��4��ɼ�a�H��:}�Wwf�����d`�v�y3�E6�蘲�M��1@��U�����,�@���/���4�yW�I�x<�^��g�����ӡ;����d��[2�,K]�HV���+E]���ݢ[�0[U�u�T�G��N�S$���-���J�M!%α��u�y�fom��ʋp�':��m�a`�<źx-�o�������D&..�N��%'Ruڬ�󎧒�}���U�}��ĺ���a�v"��2k$v�;�/\ ���yO�i�;@��.E�v��wA��Ò�%�T3��+qLɉ�31�s]t���V{q]�5�eC�B8oG����s5H���򸸜ҟ,��i��3p����wB��rAdkUc51�ܟ�웧v'!!�㖮�0�x�b�B��Ȍ<mt��ۋ���h7���-���xUP�U
���h�mHI�ɪ+�9�p�	hƣQQF�6#lkFƍEQPhьk��"��hѨ1�X�lZ�dM�6-��h�Ƭ�"�3Qh�,�F�b�h�Ţ��*(��\n+�6L�V"���cAX5�F����b��%�bbL&�2EV �E3L�h�ɨƢ�43%��((�+d�Hh�)F�#h�F6��DU���U	�uag=��B�7��0{�}���?]h�;�Cu"+�P���cS��Y#2ޑ#�ֻkf
ge
�\���s�=�ғJ����C�[{��J�4��R���qK'.����p	�1�{w>��x�bZ�m��6��!�_B*\�����7y�Z�."B�.�=Tl�ڸ�Zas�~����rCn5��&��A���u�Ӱ㝉Nw"o�Ļ��y���5j�+y2Nv̔J�\\R�	jf�A�	��)a:�MF��y����ڛ��S�nȕw�ܬ��ң���s�I�x3-�Ko�+��4����c��Z�7΅��.�vb��&�x߻��}�{�4;<��]:`/�S�6zɿj��2�&��iʘx�.�E�͝�N8�|��ns�g6�z;6��ǰ�LK6ƍ���Id�k�F�,�tN8���R���O�vdT�dw0�.�:sy��_8]cL/�WQ#Q��F�	_�W���d��U���Й٧�5�li��-����PU3C���sM;�[�M�Â*�y�g:�W�%��T3��k];zs�biSx�p�١L���-��f�YAw��it�Ssb��"���=�k��M��V;�Yx����ֆZ��T���f���m��{W������޹��'R9�]GIc�s�v����p|���Q�:��8z~M=�xę����W�@����H��q�ؚ�v��k�U�NO/�p��=��8^��#g�ފ�u<��v��N�,�1Y�x����.��ӝq�/�[��[�no9�]!_!*�jUn�ܾ��%�(a����R����cCK2�0���SJ��j\�6��Sw/�Мqn�7|����%69u��B��:b�[�t/�a�S�{��M���˕�c�؞y;t�1ev��rf)q����W
���#�*>����d>�r��������:�$-1.�-��电�9�p��o4a�Όp�b��c�E���0�x&��5	��\�P�X^^�MX���<��}�-�8��7���6�go�<#
XLj�g�S��@")1/	�̒��6�yt��I�5�.�R&��2�����Xu�b��Oc ��Wf�ۆ�ܬ�ͷ��[u��	�QV��C�ϕ�Ʋ�rX���]n�7W\P��m����F`��[����W��ԥ�VB1Yp�h,�a�xH�:m>����9��gN��Q��M�S�my��SĜc���'9mq�j�۸E�meX.;�0�U9����;Tti�U��C8���w�b�#bx�'��>��V0�)�0�����4��b��XR5���}SY�+Y��V��۪�b��*_
�u\V�iP�J��s//_+�%����R܂��d�^UFBλk�=W8�7sv�f�f'�*�lkQW:�\=���}t�w�;ۙ���Ly�b��LYMH^�)�p���I��d3�F'���ko�p��o��)a�7���cm��7d�m\��������+�����0��v��U�C���s���,��K'����2g�����D��ٍ毐�0��\:i$�;�uQ�Y^���qEb=�_����LR��'d@�cJ縆��ω��Efb�n���� X�ۖ_@9U����+-�[�d��,ePN�X��L�L��w�C�$��+�ê�] S��N��5��rk�[K
	�z�ܝ[�&����Jj܀��h�4��)n�5&Ӫ����9��>ݾ3�fD�0V���Z7�r6�s����[�巐�8Ą�쀵�+/ww���˻�e�UF�wr0�N�\��7�ḷЅ�"��S������xf�q�؛�4�ɕY�Z&��ںk+{���j�,Nh�n5��U}���1[Ŵ��ή-^t���]�ه�W��u��v�p:�+\3�u.�|��=4���iz� w�2�M��~��S9�i�����$���Řc+���O���h�W��h?N ��KD�Z\����}��ʞ�e�	��{[�d'�5�:e��gZW�^�+-�t����U��K��+��X�H�Jm[q�wM��d6�����=4�zp�v/l�e�,�ל��]	w�#��ra$��x���u�0�j�����ˎ�Ջ��L��F3k�ƗZʿ�[�Ἰ�����ݫ�4M���uv�h�;:��EĘ=�P�浦�(�ss�Z甫�
��vǙS��� 	��#��4��%+�=�52��8�(�L���&��ѝJ�����p��t9�6Lq �pz��:,)��9��]�T�2���]����'<ښ�:`etj\�y���0vge���ƚ�w�a*UX�����I�Q՘ܜ�9
�.I��y��V�A�	7�MlD��s=_�t��;����ѳ�V�+:)�E����q�~�}8U$bL����ؔ�OӼ�B�D�yQR�#и�a�U�v�%��!�Ta��1������3~t�!*�*��6	�:���S��m��aoN�I�1��C�a��]�P���)�w&��ɞ���hc��Tx���MDc�s�o���/��u��eߨ��ƫ���.m���Ul�ß�N�y"Έ\埓�
I��ٞ5�vs�M��q����(X���uҝ��Tz�{s���|��i�I�m.^��m���J]�V��P��n'O<'�x&��=�'3�E<��k��Td�Vd��{&�gZf��j��p���k�g�D�39���Lr�Z[]еXc-A�[��Pt�� )�R۰�ɝ\�xW�2\�ݸ��n*[����j֑�>w��kP�Y�Gf0D�|�I/�����M�kw���q��'%
J,-I �N3�*�X&�*���>�� ��Y�2����kn���Q�K*�n���So�#zS��r����3�/���DƷ}K��+������9�qP�j��Ƚ<Gd��{W���e\B#&�V�P���iU�p�s"%k:Q��iCW����R���O�a��������ZE?���Y�*^�����ҡ+���q���u��7�y����x��V�=�j;l3��bF�4�jx��P����NNP̵��Ǻ�i�q��l�k��������3
*"^��+s��T��3<��t�4;�G�����5��V�y�U�d�wφhLt�6b���Yg����b�k�ӎ��-��ۍ�i��c
df�-�9Z����P��1�5d���%�����P'�{�M+��֞\��8ri�2�*��kiqԅ!=Q�F���ߴ�{����8b;�S�7q �G^<���̱E}8ٱ��"��fFiʉ��#��m�m�F���I�:�U�Q�������dE���6�(���$%9�ۈ>�7S�gu(F��&3j�l�v�c�v��ْ���k�8�a����6��G�W��8�5�66JCvb5s9ّ]���ԧ�I��):P؞}:/��f�xjN�
���s�C}��gǉ�q�xI˸���̈ޜ��_�P���=����B%������"���KOڭr�؝6������$�J�O5�~����SUg3r�m���+z�V��դ��'���%g���e[Fe7���V��R\D�����q[;q���4����k#Y��Tϥe���x����R�x/T�7i)�1�n3,��9���Ɯ���Fo<#����(����^�%�)o�_<ej���녽�WXbii���Y��q�/)���7%�w;C�k��+O�v�ڽ��
�Q(Ԍ�������E��ەm��.��"[��r{�-��:�3�����U���kn�d��]�gm�k>U]G���j*5�y-�i�i����ӫ(sՎtī>�O}�Uy��N�Π�W�I�k�'!n��Nmzn��I��M�N���4#�f�V�du����i��F���sh���x1���*���k�:��t��x��;���ڱ�X-����H� ���˓���Q�|�a�V�[����P4.wmSܞ�Aj(ю���KF�<)�ؓ�ӳ\�M�1�)G5�k��gj27����b5%д���KN�9c]����lq�5�o1�#�u�)�T�ɞߗ`�il���%�6��lԚBy��GR��o��C�s��d��?:��p�����\�u}Kǧ�4=��Y=Q�諪SK�ۤ��њ=������m�������a�{��7����0*�hH5�I�x_����6��������:Z����o�W���	�s��C&L:�URPc��=�� <�C�yx�Y��O�}9W!���e�)SС���&�wɿX"���O{1��%�.Ic�s4���
�hg*=�5�k���e���9���K�O�p��>56a�I�sK�%�����w��l������
��5�!_��t\+��v�s�yח��S=�3��K�tM��!�j�ס5R�{Fk�S������"���a����h57Ҫ%�V�# �ǫ�̊�{�b�@+t��J�e_�Ld+T4Oe���a1o4��!4���m��Sj�/����\�m���V�-�u��vWη:�q�\N.�'v�T�x9us�c��`լD����)��GY�MS�5S|<�R�t�f���+y�O���9����_�w�y����;&;Ք2�S��n*���CZ߼jc+F\odi���k|�D�|a�\��ljh�s��$���y{+]-�50��0F��+���\禩ϩW�����mW�]���-2�=9�~���>g��hз%�g�sc	�]g���bg4�)ϢG9�O���X��7/"'|}"o�q�����/�T�R�;^Ϋ��dv�z����z ���qa�8��sCȹ�T���a�v���[^����"���y�>Bk�jh���&�e�����U�#�� ��Q3�Qu��Y���W��ѕ�-I��'o9P�m[xoZ�+�}*֌�^�3�������y�O�����?jh��H�E�
�O �O��p�>�w�����b��W��֐�u[�o�[+��S�q��Er�4#�A�������܎��{�W��+�vGHL9�#x8|�u�~��xg1�7 �{޸��g�I�zit]��u� ����fTЅ��5=¤����S�o���m_�/�{�ǆz�|$oW��H�U�馒ܘ���x^��գ��o�o�{aM��I��L:=�NG�m#��N�J;3 ܩ��Yӫǂn� ��"�k�{�qN�ㄥ{; ԓ5���c���i3|�$ީo'#թnvp\�GS;�8��[ �I�P�\�k��>W� ��U�[�>>"�.�E\w-�>���o�ϻ��۽��f�ao+�Y�u�X9H�`w�,��,�P�G�b@}�v�~z��N�!߬z�3��2��獛9���"������=��z�3�{(�z����y�6=�Q�\�~we~��AR�f5x���Az���Ο�:��������ϋ�u�V��̞�R<6R�z�/t�מ@]UU�v�]s�����4�h1u?��wȧG�#�a>&+;���y��,�~���vw��}�!��N�V˳XF�ӯ�-�2���Ң�^�H�Y��{�;��W�z���W�mJ��������k%U���]�L��ȜT���<�}2V��"[~>���������Ibߢ��Y��cNb����t�ҾK���GT]o��_[3-�G]�?�gO�s}���7����ç�|�K�_�ϓ�]���5ӫ��԰���@�0����z���ǗI���t���@C�������}�|'���7��~�>�]*$��ʜ�&\�DE�^��Lb]U��J��"�EX(���N�vj��3���_�3���b��dдOvg:����j�YZ볍9�$f���:��l��C��O`�gƭ�/F�,1�5�1��ID�U��]t�ڇ��:-�.�m�N���aD�2��=���Re�"�m�����b��q]s��R�Q-{z0�xR�б[��I\2�����x���]�B�j`�vCt��Xݸ��5n��K��y��R�ؔ� �b���5�Y:�F1-�����Qˡ"m�$��6b���$1���u�Զ�j��!�6y��Z)!,L�&�FuKv�Yu|�jX�^�?��m�u�aЖ���j`�Ght�Ή�Z�f�lS��p�&]p�I��"W+5�{v���3��Ƀf�u�˷�2��I�+[�ct�ӻ>:ķ��y[����a���J�Z.�c�5��Z_˭p��Y�$vI�s���1ikM@�c���Z��&�gC�q�u�+q#m씥+�O��U3�i�u���@e���,t�롨Ŋ�޶K��7�Ed�V����K��ogYrH��<1c�ltL[���-��z��l�Y��o˛��f���۱6��GX/W��vM�lh�'��Ye�ؠ3o�T�j�N�eHIn�� ����od�Z�g���e!mVV�UZ��m��FP�/%I�yh�TK��qoLա<�3VG��!�	[���A�ە�)-d�����X�pu��;�qPŒQ�t_Wx��YXG	R�=����we��@vlSK4fZZj�P��V�㘂��U�g�B�G�L�d�6���VV�w`s�A[�[,Q��C,j�Mя�ik%9�;n-�����_����71i�pj��(@�Q�{[�%el��TxX��<m��Ѽ�{��׀�U�J�Z��]�F�J/�i�>�8,��:���b�bg2�.��>��M��P�H��b�i����o�	�ݏ�:��Y�r�{	��5�22��S���0����tQy/�|s;yc�Q���4��֝��&�\UiH�!��$���nuNCh�n��KC��t9^V���3%=�0d�`��̠�Eəmc���Fp�@��J-n��q]
����]��Ne^am��a�]&��8��(4n<�7R��Wn�극P0�жW^1yTq�Hkd�Z�-���\r��&uP�����
���v;^ͨ�����ŕi`���Em�#��)�Xsz�'$�w�n��AqeX�]Ӫ�l-��	��C��	0[hWT��t���j�E���M5��I2k�r��JJ�;��2��5hU���v�+���'Jc&���� �GfFm�0���`�nJ��٠�%�-�r9`Yљ�]<x	x�H-�����(XC5noFky{�l�m�Be8���JI��^t�C��N�w<���G@Q�1�5kg2�WjR��O�ee��ûD=�V|�oF��r��\����jl���菇��z�B�xP�Q`�Ŷ+m���ţE*�54b5��VKF#cE��cZ(4F�Ti*�n8��QW���ۋqE����K!��+E�W��TDQ��7h����6�h��6�ۍ&Ƹ�\���Tk�k���5qW��UUU��9%ɛq�7��i�-:�}��4	�c%�v�oO��R7����K�k�:���>N�	�1��m�VB�U�#_o\�{��Q>�9ߞY�TV�yߴd/T�>��\{U��:��"� ��9�"c~�"�O���zgT���OR�
V���'��:+�������k��k�?~�Ϋ9e��o[C!._��_B/�wcFq��V�G�zԩu�\�V��{���
���ᵷ�緾�К��όQb�
a��k�����\u�Cݿ0a��bvd�؍@+s^�ǜ���O�{� ���d��z�d�waU:���4uE|j��y'yg�ڙ�ɕ�~�٭��=���L�>>���H�L��!��%�*#��ER𿇫&W���[0�h��9V�<���|�o�����k�q��wB��z|Eǽ�3����u�7���o��x�(�G�OD����{�NVJ��;���9�OC�fD7����.#�P4�w�8�?n��Z�ڋ��>�-�K|�V(��GF����ͫg����םw�l�r�N��C?L�<��xJ�W"��ꐽ�&����J�S��AJ�����]yu����>��'nu���[���T=�{��^p:���ڭ�;{��:,�/
T��f/����BgOgew�y:��E����.��rǗ��;�E�Я��gC�.���-L�GDIRR[�[�J��u�b�Lx��R��;eKy�k���`8��wc��8�vU��7"��A��+��H��w�c���et����2�C�~�
����O��l� zq ���Uo[9G��ʜ��{�2#�a�4z{!���CH`zfY2��N"�yFG���o#^g4�ƃ#�y�F'<X�s��?��7�z�I�ue��t ��Rf3т<D��6�cȮ\�羚�g�>5�m��\.f��������(��~ ��{�_~#��Ȏ�\g�X��^�u�#<)���<iJ�vi���7&���zr<����z��b�{z±cqX�Wګ38��3>	��`��P�O�E9���U9��Y�ǯ�_I��?^�ǘb�ۘ���nܸXq/#��=�gG;aJ������1~�?}��#�~]Jj3��~<_�(���\�r��=�5>ҽ�.�9���؇⧀���5;~& *�2�O���^=4��Șڸ��/{����c�������[b|:}��{�_���fn=Y�G�TL��3qeͿg���j�k�yX�2|'�vvM��y�J����Rc�W�����zw��ɒ��UJT/>�l�2��]i�\�-Q�$���׎�f�~J��0��,��]�.�����Dg7O����v�[�V2;�py7;�_����c\��zF�@���miy7a�#�헜u�yޔn�왱���<Y�C��w�����(2���a�.��[XΜ�ȓ�3�^�UF���rb�jo-�p8�|.�\C��o��z���N��{g��5W�\�������V%��!(��Z/���s�]�O�Ʀ���_������ʫ���{ާ3]m����{MOO��Vr��b���l8��UN_�S���ﴚ��jo��rØ�|�K���>�Fk��FW��oC;���0���	�n^S�Ճ��moyg����S���Ӕ����b�w�g���5����j�����~7���������Wf,2��?m|7��"�j�,X��;}�3�_-JF�696c�B9��'�O���ɒ�^��`��W��t��>�Y�:ͪ�˹�_�Ze�zr=t�;��wy=|r��ر�X���hG�kp�/��Ċ��㬟}l��FZ�w��&�x�w8��G2�]��{��uf�[�烽�}b�D�p��� t����.o�Q�b�1Nݼ��C�s�(�@�O�ym��r���{|f}��n}�*��M� t&4�Z�Z(o��Z�/҆2w'�z+q�KL��OV��b��cҚZ눣�s)oۤ��{@�yKB��4���B�j28�/�J�:�wu0�+z!�oG=�:�q��%�I��c|�)�m��!�����]��xr��z':��	l��U�fC���2�[Y�(2�Cc�jq\�0}���1z��o�g�Fy23�xz�' �.�x��~˗ H=�c��D���
�	�F��y\W�A:��\7���e_��S����T�P���>�4W��^�{���b="�W���\��F:�[b3�V����Wh�z��=���肧�s�K}���( �MK�<D�P|*Lu���S�o�����~�����xV;aR�#�0]�G�^o-���MFD��=08��B��n4���ˮ�W�K��b}7��qC���^U�m�Ž�.;~��/x�-��3�rb�_�Ԏ���|j����^b^����k�y���s�_��>���{�7B��ύ�����罕R5W�F$d�j>�Rt��A��9���Uvמ߫��[����^�l��^>�>��u���޳S���9{ʷ�1{��4_�W�y�F������>�8g���/��wȊt}�3��{��y]�u�9��{Y��3�3�)��\&�z�U� ���R�6}��6nG�nB��M�G�:^�H~��

{~����ݏ*�XD ���=�+��a+�Bg֡X�1�վ��]�>��L��X�ҡd�L����H��z���ٻ��7��yJn�,�w�7Qr�]S��k�r�p�0W)7z��ؔ�p��k-���wZ����齌�Z:��'N�����#�F;�Ѱ�v�C�5��+�|2fg�4L��^7��a勉sw�}���y5k=�=�����eOp�y]';h�)�`�0�z�����{0�`n����ɼ|/+9s����r�/C��\G����]���}VzL.�S�0���"��$���W�G�b���,�!��\=�w"{��7�|=��	�z���V�r,��T�O�!RR��ȫػ�^^3>��1�x�z��5^��rn;��ü'��~�uǵ\>�X�'?\o/D�2�^B6iy5�Ƕ�3�
s5�^s��s���z�T�W��������*8�y�F=&����嵲�9�\�w��ȟ!��CB't�ѐ�v4dc{�;�rxU��֥O�̹��J���VbH��=���Wo}qZ.<|b�1A���f&��^<E��C��\M����!`��a<yvc��~n��@�������x���=qFW��ȩlO9����m�~<w}�'׶ٞv�H��J�x\y91��j�B߼T�G��3�P�ɒ�aS���~�^U�>��Ok�}�$VF�ϐ^v�vZq�`���|�Uhg��Bߥ�yVڕN�.��Y�鮲����GN�x�;�[�y������|���8��%7���wC��8�qM�;�i�(em�+��������-�Nh����τsQv�O^'��L�8����O��+0�7g�q	S�װǔ?;�C�/{�g��	��ڡ���V�3�ȏ;���V���t��ѮÂ}���I��/��5yp�?]����>���ޘ�D�/{e�2��Q[��v����{��9P����vk�6Qu�oF�s�λ���gݑ��H�%U~�{z���3�zs+[�5ލ9&Jxk�2D/@��>��{]����ݺ�t�ٯ���ي�OG{���W�^�VǼ{���f�xdvWI����LہP��a��tN{����y����t�<�e��,��1��T�t���1��<�R�i�9Ք6���۪xy*h��N�w��1u��m���Q-�^�����{��\?�7+�=j�ދ�?�9O<Meឧ��ۜ�< �ߢj�]�u��GTӮ}�r�{��=�<=��&:�0��y<��<�^�P�k!�K<�1�)�����"�3Q!���ʳᐳ1nٹ6ׯ�ӟyO��nb�պ��'��ڴq͍����ݟ
�!�e�P5|�Ҹ��[�6d,}��òb+�>��)��"&��d稚����.n���(|�PB�d�(Wp��]d�#J�[�ԡEu�S�Y���<�{)f�����:U�K)'&�����s��/���n��]�ɕ�uj;K_<8��]��R颟\�O�Ђ��/2ܸ������>�m=���.������{J�[�3��=�Mh�e�w7A�3墡̷\@�^k~��+�>s�F7��z��Fh��������9���~*x���煮ֺ����̷F�MU�֢���������!Hh,�C9hTk~)V�������q�z�g��+bP�O���_e�t�G�e	t���:{a
~�Rc��~�o����_�����*��1�x��if��3�����|ƍ��9\J9!��3�e����}����&�A�'�Sae�w���Ԓ�\N�0cK���? ��9P����i�ݶ}��o=p��K��:eX����?T�w�<�O�|��������^͛��UHߺ�3����
���C������Y�l2;�:s��V�z}חӑ�O�>�O�^�sZ=�'���/i��FJ�ڇ�ޙ)��3�5���O��<?nd����n�9L�o����y�G����;/��fz�t���ǚ >m`{�t����K���h4iĕ�WϪ��������K>G8TDk�S`W�{����N#���G2�-��U��G�YbU�e/�wuR�5&�ޫ�Yz2�o)����$�oC���T9Z�[��n���=�
�<�&Z{O�Ț���M����eh�Y{҅c����K-��f��S�eLq�:�v6�9���y%^�x]VO��h����<}c� gδL�;�����~yf=;�c��:f��J�qk��9�kE��W��\�Y>"��fXy�7/>���+_|���A�=���ѫ|�\d���U�S�z!B�4��s<EC��}�J>���b��0�{#o����n�vf��^�>����F�����ϸ:W}7A, �T8��}����)Oi��)�co{�F���)������^w��S�]��3/��y;2\��`#
�gʂ�lP������p������H���C�s�g��c���Hc���cޡ�\{}u;�LP�sժO���[푃�pq�D�&zE���u��-�*VC>��dz���oު靈�������p�|{����8�*J�$�ϧH���xT��1� ���S��Jܹ%��J0&O�D�����q4��V��0cbYu��b&��k�A���^]5�q"��ٌ���ۆ��Zm��br|���ng�z<=3�_1q�%�.�L1"���0b���,"�o�F�eI$_��_�e�Ѳ�b�cD����:(&7�
Gv��ʶ��ш
t:�ZU�Gi媐�f�`�6�Y�����6�K���Ci�E�V���4=ɲ�z�t�s�z�З�d���^V_+5���kf�����Z��Q�\ཤih�����ߧ��}S>+�z�3���n{�U#Ux~���ѷ��ǧ���;��w�.�\�����Hlr���.C~�ᏼf|]g�W_��n\�ڬu���ҾU;<f���������ȱᔧnv�}g��(��oS��,ǃ��OǼǕ�W{~�#���rl�ʪ�=�y����h��
�h!���W��gke��6l��̜�\z}L�g�r�#`d^OF8�Ǚ�e�N�������h�<���xf����^�ဳ3瑠�d��Kj]Kb��Ň�����.4�#޲�4�t;7�U�����\a�_���~A���x�_un��=3��0���&������\���>�QVzJ�5:C p�������Lk�k�U�>K)q�A�,�!M1������{��3}S���~�3��=*�X<�`�v9����J�Nn��@꬙��w�Ku�זk���d�7~�ީ�|=�1�ڮq�&��}�b��o��dtI��Ѱ&y^���d�6��;���Ro���N�y���C��ߪ�%���Yd�����˽����OF$�X��;�DD�,�yQ�ɐ����6T�JvnM#�K�@��]%�a�ZhE��;M���ke�e�[LKKmIz��,�Ljek�aS�Oh8��1=5�v�
�R@�ऑ>
��X�i�l�O���U��%�wt*�S�%��:�p�t�}�R��/6���+aK�r�is�~+��o�+G���P`�-�����qi�Z� w�Op�G����z3}�<�q�yۜ���}Y>��d�{=qE�z�\����:����'|c)�ŝ�d�|��q��x_�NLu����JG�����c&LC��Q�S�rhn���r����������+$'['c,�8���𿡯mǲ��{O�q�x����cn�nr�:���P�>�ԹymP���`ezz<.]�'��.7��p��ïo}3�W���Q���Rg-�S���b]\�i{��/X߸xbr����}���]pѼ\��:�'һ-q�=�^���ld��1Z�����9����3ާ�P^S�΍��ҟZ��&7��늏�Oƙ�r�эm_Y�q�˚;��~��?'jr���{վ	��nw�X��=��`fh�x�0�n}�}�ŝ�p�I����Ǡ� ��Ҧd�&��8]/z�}�1����O%���ue���LD5>�W�I]nN���b~�뉮�|�_U��{���)��͞*[L\��J?vCe�����#�:�ҷNK��côRG����p쪭GF̺���c�P�D���3U�u0��Z��=�Q�Y5*#�#˰��29s_)�6�wi�vV����x�2@�W�A�;�l��3p�f<X7z� v���&.Qɤm$c�*�^�E��؅�ܓw���B������׷���W�IV����"-�yҊ}�__P�Pb�׫	�)ڤ��&n�l
�|����4��S�ۂ�ճjۭ�f����[��q�gޱWt��qErړ�����3�X4�ݾ�G�nsSb�}I��7i�x�U��"��e���h�.��"��cl���@M���V�-g�su��S�leg.�^̸��>��g���5ܬ/�y=aGc���3�h]�v��G6�{�d�-�n�zi)W:[�.Q(Vm[�,��Vf��+��y��H��h��b��#�<v���]G�zp�.���� �0蘫�F"��:��ھ��*��C%��Q�1L����L�يh��*���׶�KS�����s����w��#�r�&7r�fI�A�.�p���9�<E��g���ou��3b�1�u` �t�_o\c#��<8�!A��)\vi��4�u6�QG�y�˗UqjH�
2<��H,�􋑥R�;�$��Ɲ,|�`��}]/ �-�X���x�K����r��Tn���ǯ��m��W�A�W=1�SX$�=��ÿ�S,0�T��uk�DP�N��b�,_9P>Ɔ�r�]�}vm{m�;}��l]@j^�X��^ݶ.
��G2_��NQ}�2�����hB	.�Լ���PfH��wa�M�t��Ue�ȱ��9�<����]�:�q��x�-�##�>�c|A��.<]�W�|�ꊮ�p9Â���ŊfV	�#�
��s8u��Q��O3�Z̘�9v�����M�ȦT��2������M�,'�Τ��M��|]�����Ac`�͞��])�P%�N���tZF�'j����������;�u8��C�k���Ѻp����o�e�j%1X�f%���%,��I����	�t��&�zYx��7ufњ�;-Sɢ�&��ܰ3-;¸^RݡNCV%ȹl�-��M���"�۪p��l;��Vnf�|�n&��:y�p�91e�P�U�wv���صn����u{��*�_s�ۺ���KRM�z��)!\���c�c��ʖ������e<�m;l�ܱצ���� �8�S��ws�%]s�R�6uE�'�*YR�؍u-��8�������Zl��{.�!�w�f6�*#j�(*ۖJiM�x��2����t��ˊ��m
�n�<�YnR��Vͣ��FJo��)��rt־:�wc
��Ie��uћJ� �m�ɇ���I4������Ϸ6���ێ,b����5s��X���9r6��[��\\X�n.�&ŮKq��r����\�ˍq�q�ɷ6��s�+���X��9��W9ʹ�9˜����js�%�ě�.#��9ȭ�qō�q,nis��m�rӜ.4�+�\jns���p�r�h�q��.3�ے��\�5ɱI�7E9ˍ���A�"6���q\9��m��Q�.�s&����8�\n+��(���9�J�k���9�+�K���}{z��_{�|������"e�Y��h���VҺ�R��t�5-�)��{C�+�^_w^K�/��Q ��!�P�]�֜�^�&|uw���S1낽wB���0uz]��������\?�n��O�Ĳ��:Ŀ^���#����'^��zUlo���i�D>�y�>�q�#������9��`>�]e�55�ӱ/T����Rn��"��H�n#��>0�훓mz�=9>i�,���e�y^�����}���t������O�����[>&�B^����ۧƢ�[ƫ��B�3��{m�_���yu��/i�~��q�*kC�P���L���B�<ށ�f���}4/��i{H��G��b���pn<|�K^C_��@��Ƨn<K�?:��3-�>��º�X��Y�\#J�yV��bC5�6G �MF��£Re!������;"��^�߫<)T�6�6��\M��/w��������I�VZ=��?�)1�������[֣����b�6���>W���ʯ��T�բ���G$Ӯ�3���{��mx���&�M�w�@Nk�}�����^��^s'{���@b?NT>��`�Mm��u�o2~��^����d��MoP���}�phҢվ��� �;���wZ(�ԣ̼1<}0:�K�l�>H�Uv�(d<Š��v*.�"����q�Ȼ���#�U���Xŝ�sKꦎ���jR}8�Սl��д���	C����^?�n���t�ͬH��)X3�;>~wu7|gƮ��5�=�U�3�\2�%����Cf>����س�(��~�@�6�u��/Y��=9�ϧ�'�2xρy�ɮ�=�%��8��ߌ��c��3�IeՆ�{o�����A��,�-FB�~�n�9����_�w�g��f+or�Oz���.���G(��f��.�C��K�:�Vp� ? ���V��{)���3�Y�����Dmϕ��v�3�F-�_�B��&��^�%�����~c���������G)�y����:H畎�޵q��Ў��5�π������W�ߺٖD����^{�K��J���)��>��N�{��,�>*|�g0�!v�C�υ"�R>��)  ��̼c&s$�+lr�N)3�frg'��xno�Ϻ߭ϸg�uҮn� R!đQ{�/�4*�t����y\��D}�����0}^w��|�\o���y�D�\��E����w��Q�Z��Y��LΪ��2f�x��
l<����~W�}i�U���Q�����A݉��a�$,|�j����L�a�2�>.o�:���'�_̍��pS���7�9Ͻ��ۣ��4OY>���
l��X!�ܒdOiwC;��hx�9���r���k����*�z;�R1D��8��<4��kX��p��/��U�ͭ��45�&=���"���?�����ǨM�Sg�t����[�T�g�؏��7!ޚ��(����N�1����ɫ��O�IuA��j��9AyQ��l��b�>����{o����њ�x�ȼX���'�����z�|�]�U08�MT/\Mv?E>>#kh����3+F��tVgz���~V%����7^�}^��g�\d��������EK�p=���p�uyNd_U篟U����;��׶�8��и��3>>��Ώ9�2��jA�^9昽wV�g�ĳ���s�=���W�t\m���69S�q�yp�]���3>.��v��{r�o}؄{r��*�$��s��=��:r02���v�]�>����8f�?ηq�G�!?V�(��ޡ:-�.�$t8���G���`�?�����1;[.�PٚU�_..d��dzq�}M�c:,LR�;�5yv-��f����M�1AQ~[�����^s͂fg���$���TS���ՠVn����?+hT�~>��I�F�wB����5���D;
q�����H{������u�w{%�]�V��T�e3\N_O�ŝ��m�r�wj1��o(�oVh,@̩��9�N�C���m��L.��}�"��g:��(���1��1�ש��F0�
�6}����:����x��y�C��h�rh@{'#g.[�C=S<�Q3
1�'�=��Wl_��<�]���ܖ�-�f��y���s˗��A1�>+�g�a�}t|E��Ji��|���Ox�F}�����o��d3��uҪ��=���2ߺ-U�Iz�~u� �Nf<�GY-ק^Y�Q���߸dGz���/��̷��,to�VO�5(���wA��'_,���Q���č[�x>a�D>���z�T����N�<����F�b�sܸ�W�``�D=��m��!�M�`�()"j�}Bn:�y��1](�Ї���V��o{��ʟx�nsս~�������\x��(0�e��k������OOOJ��F��do����#3���;�r�=7�ۜ��@z<.|G��7�����z�_�*[A�1�b�qSd�O�*���\�J��y9�ވM_�?z��8�L���\λ.�U=��<?K����{כ�g�&�+�?-v�e���bT�5�1��������g�w%u7����^ĭs|�h��Ϣ{T:�De9�VK�KF��Iާ��	�����]�C�U
ѳ�d�̵6�h�p9�ݹQ�pa��U�͎�+�y�e/��+NpTQ��ݻ��y���O���=Cb6�q�?O�o!�{ι2�L�E�7���4AW��u-�xOI���r����ZoU)ׄ���п䗅�]��+�v�z!���Ԋ큝����z�5͜#��*�*����k�6m[<f�s�S�Y8b��v�BU�흟|�Z����'�ni\i�2W����ݱP�f�D;���.�>��{�h��䮵�w�����̛��ӑL��½���������Lg���`n�¡��Z�d���=���M�%��^8N�� �t��1��eNDKޡ�G��>��6T��i��CriW��V��V�p(�v���,_�Yek��H���^������n���~�e��y�W�6��VDE'��ҽ��RCg�n�j�� �y�O�E��4��xܸ�W�{(x< ���eT��e{��^܋7{Y֯�}���􏲂u����G$VXO�b$y7�U���i�v���(�B�'������f���,�w7�|:ߝǻ>~�n� �Nf�%ꩱ�۩��!�%�Dس7mT�ڽ��ֱI�S����>aw�pm��FJ�ALO��P�<ǓvT��ܳq~�Q� ��=��-�j��+�q��q֟!��O{|jv��.hê�����:Ee��MI� `����j�P�1��8�
��g4���\k�����J;�M�a��P�������l>׉�Μ����ga�m=ٝb;��5}PɃ\��Ow��9FU���o��ZGMw�k��́��f�'Y]���4���ʝ(�1��������w�,�"��G�8W���9ց�oŰǫx{�G�싈��{3��������#=oR��:�<�� �b�P���⤣M��B��������~�p�^@x*Ňu�����ˣv}��O>����:�UT��!z\��N����[+�ċ�רO�b�B��U��fmn�q�e��{ޯAϸ�W�Rii��4�d��!���]���fz�By���ڭ�]��W��?]����wSp��|j���3]kٳsq��Ruxbr������Љ�>�̻�*�y���V<Fx{�G+�=7ח�r'�2xρy�q�'�������C>��r�x*����{�ܾ�Q����f����u?�:��r�>�Uk�����V흚H��(��}�,��-/���V�CyJ<����v��o�j������L�����K�Kq�P�4f}v�h�<�+���8�O��gW�h۪s�J���:f�O�`�N'}~�}���wvܺ����4P��dv���d{�{�k�;#3���ʇjer_l�Ơ�����.:ٖ��S|0ڪs&'ot�s<����G�V�ұ�p���Ft�������.X���R��G��0b��Zŗ�Z��<��G|�C��qp��u��km�W�Ҭ��(6�j꾭��告���7+�}��C���g1X�[w9<����I�kЭu>�{�%�8��]���GOD�����q~��D�"ox�w=��||T�H����y%����إ��%]SZ'0�^>V��wuޏ[˘y��z�}�=��{�~�>�U�J�0�j��@���|��Pw�Wi��1>���>�x��+��~�<ϰw��>uپ3/����r���ʛ��*I���~^���g�9�^�H��y��!����� �u[�{�`��ʹ�}Q�E���G:��|��QuR*���M�6zE�
~u��>EJϡ�[b�T�X1���Og/��k�Uv�m���^:�Uq �7O5��V���b�>���w��U�~�eW+�u=��n\�ޯ+���B���rYe��IyHG�쏡V��S| ��u���'(����N��o��wSi��=�����ɋ�~�R*`q�/���M�����5¼7I���$��v}u�8����^���?3t-�ύǽ~�����sq��R7��V�F��ޟ毝��9���O����!����ˇ�߮�gϼf|]{���	�W���d�c��5Ϩ�j�!�+�jo�r��p\o�\�kFZ-�N�/���V1�<�����{N��-�EQs;5�{k���n��^�������s�:���8S����[}���^-���;2���\��Z3X��+LSz@wA����p�����l���z�{g��=���8ezTh�|p�v�/��oS�ηq�t}��̧�w��+��r6��#Z=�7���W\~9���+�ᵷ�W�񝭗�6nG���������b�ѺY�#��,��FϢ�Z�H�������#=uZ5튇�&����}�i�������Ó	$�Ò�nә��g�����}!���X��+�����`yt
����nm��q̗�X��.��}��}�۲.#����D�bn����/�Ϟz�O�eY�0�N�zV�������:�9���=��
FH�������w"{��7�|=�=�ʫν=��~˘[��^������1��ƫ�0�Cβ[�N���x_����G7~����z�)�x��n/uׁ.�1<[~;���ݑ���H�gȊs5�xU�Sa�>����RJ�sk=��U7X��^���?j�!��CG_��Hw�|�`Z�;��`5ݍT��O�ި���\|�,{;�y[�9>v�=[�����{}qZ.<|b�����B�Z�y􌯲.���!
�zy��sӸ��L<��x�h�V�+O5�/]���n�&N�o�I���ᬡ�sP���84=��D�RI��j���C�s���2���9K�m��Q���:������+�Xs]N�]�74���;
kk���u1:�UB4j�3� ?;�0�X1��,�m�ۜ����
���x�ϯ�)��r��Ӿ�pV�7�ߪkG�BG�2������?9���5~�?x�����ﱃ�&�mc|����ќ��^�u�l��U���$�{���K�H�J�k�q��'����g�[$��w��7r���}3���n��a�P*��S��G�ˡ�2p�>����4l�N��Q���`_�z2;׭V��G���P�mzk��t�X����W��;���ó�� �1��a�-�j���c��
�߲y�nv}�����~3ާ�yD���@o������c~����,l��Y�eun��ŭ�S5��5qS2����^9�^�k	�3�=��s�jr�Sv����z�\�r���鮧����@���p��^@(�s3�bk�S����x�[��U�ݕ��"�/�u�q��z�}a�ݻ���@X��\�yg�G����(��,J����aY5�P�G���U�N��i8)YٽC'�~��>15].��'Ƣ�ٚu>�y�>���������`ʣ��k��÷m�J)����ډj��M)fȽ��T���:92�!�)��wU�v��~xu���iܧ��W�%���.���O�X�f��*W[�VfN�D�G�Ȼtƒ� �Y�����ٶ��9���܎�@����I���hf�/R�X|�=�/���H�b��H�o��>�1�NG�e���{��a��~V��"<�����χ?3��88C�~�jB^��S���X�T)��s{��ӵ�+1O���g�_�g!{��[Dh��#E�,ÿ��0P��#$g"9�(�,�A��z���:���5������yZ��!�ǧ��������\�__���̫��E��g�ed����BB�t�����9ց��o������ߠ{Nȋw����GwP�>St��ݴ�)�Ы��H\_���&����7��:{P��q�Rc��~�lªt(���L�p�{���Y�DVx�0re��q:�^ȔrC�gr�\$_pĞ$cha�=�UU�9�~Wt"�~�E�W�{�9@���&�j�R�}(c�_}���z��UI��L�� ����S�Wy.q?]����~�L�\|��7=쪑�����}�t�ȗ�L�l��o]�����k����D{�����q�y~�꽡C�m���~�^A�����Y_}ߖ�:Llͼ�l�NQ�(t�����ÌF�ݔ�|(4ͩ�n�]Jm[ɫ�=|��5wW����:ף+��s�Vv�]���4����e�;h2"E;�1d����u����ŗNNq�%�2��s�^�����/��b��|��R�7�{���s�_Ch �(&q���ޝ:sM�s��k��'w�m��Rg�K���-�.L�/�����������t�u�ڰ:-��uua&��b�s���!�Ú�P��6�w�.,��&����G����9Am�����n��m�S)��AIv\{J�]�q�v3���aXpa��������d˺JWm�P;� ���V���堊��h�w$�vѡ�v&�x[P�t��|�[��j;�\����x�̽�Ƿ�*�xEj�\ջ�W.R��ZZ�����B�n;�VX;��<�A��qX��fqbS�wO��ÀrC.��1��cX��'7I�Ա׷[S��yw	����D��f���)Xt��6�v_4��r6���4ـ���ԥ3�vE3(Q՝cu�Ł�Yru��-Y�U�sm�ݼ��U�q�/�o�+��3 ��ay���`����V��r�͆�T�ӹ�)�O����3b���׳*U_*�Z	�x�4-XE;';JI�q\:̴	ޭg�5x@�.�n��V�xPs�l�6�Ȋ�[7���~l9Mr��h#(����W ����3o�F_Vt��d�7���fb����:�	E����|��;ڜ�E�F�M2����-ע��%u� �N���
]������'���:h���x�é�*��J�3��U�rpf�������g&��7-�]��o�ױj�#_��;1=��}�J��V�hvt�|�keμ�6�G�䃳�k�I�V�ὼ�BW\VI/Y�Ii�0�'\��%�7]T2*�l�rDnɺ�61s�t<v�[�x�dK4^Ec��m�h�&��2Ī���)\�ŹP�O#�.���mL���lf��4,+{��L�9��;{�� [Fv̭e�F��0���Ӆ����:�oV�	n�Q$���6�X��׍����!���9cY���M�V�=[VZLݜ��[��;��u:�q�`�v 0W\��Cs�LhU��!�ɼ�*U��F��3fy����9+R[X*K�(d��<����AN��#�cv��_	8[n��%�U�nP}�9i�c�)Ҵ[ê2��<2�;Q���me��7tr'{%��_Lk�_+�	���궲��}X:�N�C�w'p��ǆ!*b�j�e��&@��X��җ{PwP��=��8:�ʗ/�H�:��XM1J�C����9�7&t�в��8b�V��S���[�>ҍ٦%�t���Z�=+8VX�͎f̕��gA�8s��qְ��T��S�FV�q�{�")j��<��	��VG
dwц�61W*�E�觥xѠ 4*����(�s�q�F���j8�خ'9���s��99�\�\QDn7Z�7�s���AE9ˊ�9ɖs���.a���p����Z�LF1I[��s9�eecA��qq�4\[�+�2ENs�W9�1�"�Q��9ˈ8�R�ۜ�b����h�c�\\i4�cp�,�9�9�N+����P�CM���W(Đ�(ܑŸ���B��9��9�	�18����⹋E&�� �$�9(0����F�#b\nP�!)1�`ȝ]dFG{��T�ƣ#�m�1�a�3�J��[H^eޅp�n-:1�{ z諼��o$��,];X�+5qn�B�4�yv��x����5A��Ƶ� �C�y��Ӕ����~~1�u�G���Q�����H�7������J���|U��ԏ+=QQ�[�Z�+|(�W��fu��̎ε���hC��e����K!�p<��^mS�?M-������,'��q�Z(B�U�W�ZYz�Bt�9�c��;W��!/m�2���t�i~e��t*�n�;ͭ��ps����ϲu�H��q��s�x�^�>���4�� ��z�����E>>O��3�d��>Y�)�;ys�rW�k����j�~�>��]7A�p��L�b$[;���k���FD���uy��}w�~�u������>^���T�Т3ȉ�����l�7^�d�y{�_���$X�fyP�L�Kg�/�6�3�(�~W�}iu[�V�NF-���H˱��۷ჽ	�����b��P%k�Hn�FG
~wb�A�=��BGȳ9�r�����1�o_�߇��{�+;��T�T��j��"j��6����'�m��c�!�^�¸ډ4��j�Q�[9�Ҏl����7M�-���.e�z/�>8�Y�p ����K�e�r�7������xٞ���XS��30�
�r��ۭ��^l����
��|�u�T��v��:T�b��Vj5�O�C8N�$��o�{׵����C??+��5~�9�+��>�1�,���T���k�C�ǧ�w(�o;ʶH�9�����؟M�+�������zg}�1q�'�캐U0:�]�dZ��w��SQ:�Rr��?|�����9��o\>׶�9��и{�3�G�~���cM�=���ac1�-EZ��\�=R@lM��ᵒ���ݺ|<��ʟ�f7��f|]v�n��7q|��u�k�����9n\��-����@�r����u�������O��:�Ǯ'&=V8�Y
���߫��ݩ^z�Bj������W����S��n���
Ty�j��^D�$8H��E�����̧�����zG�g�/}�I̡�x�_T;R5rWr���\f�����s�2v�z�E(;���c���y����+¥|[��Fz��Y�eOpǵ�~��Z."��'x���I>�����z��x=�
f=ez�S>k��]�<��z��=��Wo����ĩ�������W���I�d�_�6�|��T� �����a��8�4�|���Ox�F�O����{�/ps�������58+��\vd�s���(�	lf�V�R��M�z��?=I�s�r�b#~���'-X�U�UmB������\� om�
-�vTֵ�|om�a�8�t�:C�j1È�©�A7��K1��Y�yt�+ټ>�ޤ��jn��q�5v��[�8D�x1
��O��;5~��o�X qT��*��D�w�Ku��yf�.=~7&�������Ww<M�j��x����л^��[�p�E��$\�
�3�E9��T�*���Ü��w���p���m�=�7�fy��W����|�����P�����m��!�M�`�)�$K}Bq���`��w�3{�v/r������=޵*}^eφis�~+������>1F!�)�n��c�n2}�����c/y��#Ю���kO�	�o̹c�(g�d���zf��z⪡�c#ٸF��=&�o���􊗢ǨME{��D44�W���F�j�A�ԤyϏ�g}�|�+t����إ��{O�}��
0���ER�$��n2���C�a��&�-�{��@�v��p�g�n�f��@!7S;ޏ�M?�#Ƽye^�cѮÂd��I��/�ɾ������g�tۇ�-�x3=���P�5��z������p��T5q:v]h�w�#w�r��>�ܜ�r�s�-�����M˟D6|�3���=�{����zrL�]U��g@�^�Pwm:�l���!��eZ���C��kC2����$
��ʃx�n[�[؆rKn����:.0�:["
�{VB��Vuo>�|jIg��0[ҵ�Dz����z�ז #]��+�P%�a�d�嶆�W,㡤��&g�Uh"��N^��֗���|p����vF�.�L���^8�z=��Ό掎��?g����εw�6���X&��� \������x~Fә��M{*r��PϽf1�g�*W���U�M]�pNf݋[���>�ue���tbGT.�޻��8�0�uz\o��st�=�M-s뻕U�'����
�{֮;��9Ք6K ߪ�� �y�Y>5�[3N�xܸ����c۶���RSMO<��2=�C��������'X�VRz�y���X}������oj>.�]!��������C��F���N�=9�>.w7�|9����W�b )g��줭�r���J��F�}
��U���W�=~Γ7�^�/q�|�ò���p�?:�0�M^�`���<+7�zbyzE�@�(�u6�5��W����>C��⧀�o�N��Panz@��d�1����Mpס	�J��M�Sg�_
h{u���*7��[c z���2�vD*YV1~%謿fr{{������zP��H~�'"��O)�������w��A��$op���'o� �+�����Y[��C��W��RmܿEp�	���m�r1���ѡ�1*���7d;�0�M�V��F��O�d��#z2�F�����x����3y�[Z�����p��Cm�1ά.ӭ3��Ψ@���{l���Ķ��Cн^`1�=Y�=�0re��T���
�^��j��d�6�>ރR?�Х��pm�d��Y���V�}ȉw�+���(���O{(��M*�,�`_Jw+���뜬^�W�����|}��W�SWy.s��wSp��|j߫�5�ٳs}�5 �W�Q���yE�싘�I�l��|�z7�5�#���t�yo+���>�l�p��3�_��֏X�z�]RsA��)�Yq'NB�Z��g%@��F��r���ZV�n>�Lg[�NS'��~1�t�NK��	�ή����+�⟾Y}'��(g#l@x(z�]�'��4���q'�W���h�k�"�7��=��Y�ɷ[��������8O��	h�O_�t\����X�ܑE��<D���}�O�y���W�'�Ԇ��zC��� �q�����5��˅9�"�9�>�)��x��B������,��T�[*��N��D������_�Ϗ��)��R
,09b�3z�z�+$P5�L��R�J}�O����b����\��^����{���3��s� ��^�:�A5��#���k*�^-�u��:�6��)N.Wp��Um��k�5nI{5\I��ik{	��M�|R���H%�~�Z��2�Gy/l��>�"��ٴx�4��*��peo}��D2�����f�Ս��%��s#���J���7�m��V�\��c�� �*M@�1�Ű����0}^w��|�}�%h����mfr*}�g$����>�q"�f!T��P�3q-�H��M����!������Hf�_Rp�����jW��#py���p��F��8��"�PЎ��?����|����rq�^���a�][�7�>r����1��z����v�~��+n<O�I�T�����AyQ����ڕs�>Z���)K��+����\��ǆG���<�a�1ES�MT/t�O�Cl����f�ΦϮ�z+0��M�H���"}*��M�l�d}>�Lﱋ��~�R0����MB����q�����H��=�R�3�~sz�𶽷���n����g��޿L���ឬ�鴯��=�'��H��h��W�����>Cc�>ח����|���V��J�^5��6v����+�ܹ�=�Yq��NU��ˬ�No��p��~w-{3�^�^�u��BZw�o�+�V���{���Wq]�h,~b�Z[u^��>���pճ�f�g����+�hnU��@�q�q�����F����<P(��h_$�ZCծ�;�慱s�5"��u�t67`u�����^��y�U���Y��>n�Dp�{cP�Y���ͷ̻w�#��]Zil�Z�%���Uӱ��^&��Y�y���c�;Y�����|�s7�\zTE2�����_�i�MpV��-�p��^EGF\t�1_^��k��S��7�i��y5��ּ*s�߯�2=e�,�ʞ�k�C��<�]����s�M5y�����
�`?@�c����__��y޻�y��bm�/z�~�>~%O��������\1�y�+'�}�wH��A��;��>"���0��}=���n��(�Ź��oydWu��j�_�gW����uһ�*��8�S���#��n�;,ׇ���L1�\���V"sǰ���9�6<>��_b���Y>��Ge�H*J�>F9��U/
��&��F�Fv9�{������{x{֋�u�Z���O}m�򡣯�o�+n<K�n�	��6�fd��2�VO��^�4'ʫ�V�)>��S���ns�V��y��@^�\V���,Pbˎ�t������ku��DMX_V"�����s�|�OM���ۜ���"��{ޭ�y�d����VG���9,�EzVUmȩHO9O���t��\?�'&:�W���{�{�}uRf��k�1a+-`	V�����w���z3]%���3��i��wy�KL\��Z����g˦�Z�S�U�C*]�PN8`̾On�lwTyN�@�N�ї}��0�N�-�˝H���r�CǙ�1P^������1f�+X��7��S}��}^�c��	��`��5���$U?�
�O��워��8������x�M������+���'������ǽt9��#���3�Ȇ2�z}�Ac�G�)�\��]�'~�}~���ۿ<��Cֺ<�N����ח#���!}�5�[�����r��Iʿb�-�Q����t5�}��Ϻ�ʯs�e�z����>�q�w��n���~3ާ�Fk�}�$�^�X/Cv��oO�ޏV⊾��\�^ҵޅ����+���vF��s2b���!׎xR��x?:3�6�����w0�׬Q3>'э>��M��LہQ�����迁��D�s2c^ʜ.��C=f1���lG�0\����w/��~���f�KWr�/��ҫ�<����S����W���0��u��=�n�˞g���f9������e�1�YCf��@5J|~���ƫƣzٚu�z�}لmn]_�o�u��z"|�������?^f=��Y���)�t$q�jG�szaS�9�c|�1��7��u׎�{0��nK^>���>.w>����q�υ_�;��< S<�o�F*�w��6cd��h��{crX��VގZ�����zg*~�DY��S-<{�:}�v�'m���*��uo���\��ʻ[re��$�'y]}3�7��ꎹ���K��뭱�q�A����9"u!�驕����9ܛ�M��#Q�tv�9|�G��u&K�������35!+R��+��K�����3l�^�|���-�"4u犑��a�r'>���׹�]v7�+���LN#�SA3�O��C5�F
�,S�:��;_������idk;��y�нS����*S3-֏P��l��Mk��C
�p߭�f��_�=��藜�=�#�i����G�<(��hMƎ�5O�I�VZ=�S���!"��l�7⽗���?;t.�����`���T� �T��(䟩�x�.n����d+~��k�tG�|/��O���wB.~�E��z'��7��(��NezcK�4v<tx�7V�珴I�&r�lG�1^�}���.zڻ�s�������O~_�[;���V�Ɓ�c�?���(d��AۃKo�w�`D�F���>;������yח�n����/�nkB;٤q�6�Ѩħ�Y�m��O��S�\�>�a�A��,�=FB�~�n�9������Z)��ށ{,c��[���l�Vz7/d�ʲ�p��@x'�e��yJ��%��V���L�&�
2a���)��;~͏e�E{*�:{yS��'��h��u8�+!���B��Om��θ��/�[\`��]Q��|�e�9���]ڣ�[�>I.�ʸ�J���7T��:$��&�T�ID��5�L��
&,`W�o�_1A�İ��nJ嗝��}^.|�G��ñ��%����?�,��8p�	t��W�t5]ۍH�ay	9v�gy��N:���Ϯ']�E�e�zF��-\odC:�g]V��)n�t0K7�{#�]�립���\u�,<������H���.w#�/�a�S�+8A��i
���F�N48�=�w� g�G����%V,������9*=�^���|f}�����
�����H6���[��q�J��t1� �Q��yu��t-w���0G��bZ��^�==��LVFZ���_��7�'n<O�܋!3>U��}���M���� ϑ���>'�Wy�F\V��x�L{�Ugp�n��~�]Nߨ�L	d(�5�$7]#8S�s���0��*���.��ZY����\�����##ս~cG��{�+=U�R�uA���u	^��P}�{o��u��k�f��֋c�!����ܬO6��σ�����?MFD�;f(�s���=bC��y�.�]��@$C�H�0���BF|�K�L�'�,��=}�����km��[j����ڵ�����km�[j���v�խ��mm�[o���V��뵶�m�����m��kmZ��kmZ���ڵ��kmZ�r�ڵ��mm�[o���V��뵶�m��kmZ���ڵ��]��km�ͭ�km�kmZ���d�Me������~�Ad����v@�������à( ��A@
 PP�� ��DEUJ��A$�*���*U����E6
��R	D�[d�D�UT(D�
��U�@'��W�2J��ʵ�i���i�6���H�ک�R�x �#)kCj�	�     sE����Y��mJ���Jw� ��ʫZI��el�I���Q[5J�-!#YJ����&$�Fڲ�(f�ƫ[��5�Yu�n�C�0�T��o ����Ka	j�s����5'@�wqJ�u��
j�n�sP������z6��يM��(�6Grֶ@s���6hu�v�J�mN�
����{fٯsRRf�#[�mUZZU��Q[0��II*������Ŷ� 6�M�[e���U �T�IjQe x�v�m6�����`�D���VMkcѵ�0 ��{�8�z��S[6�&Em��YFm�*V��      "`ɕ**C F�h14ɦ��OhaJ��� � �c�bdɣ	�bi�L#0S�0I*���M0i�F!��A)�JD�S#L�� �ɉ�L�	4ĥ#A�#"i��z�hl������������?�����+�]�:���ڒI${�����I	$���b��BI$�� 
A�6�ᒄ$�H�!�����g�������p5��|�6���"��$� `h#~�$  ������)��I$[�����������_������h�$�F��/t��=�	�@��L8kD
W���[�?ۨ��&�o�w�n�8��9����*s�`t3*\ P�wN�=�T���nZ,/]�oD`�h�ɷ�����n·F��
Q\�?տ΍Vj<6��W�bR�}��ϸG�p.cMk�Қ��42��f���N��Ƹ�����;�{/l�l�2 �|xQ�
�j@�IX8<�����D��IyT�q�fؔ�BfN�AطWq�ݢ���5ދP�W�u�rk ���Xo��rC����P`�v+��α�ō��]i���m�Ҷ�8ǽ�<Ѻ*������uX)qO���7��ڴŁV�xWm�}�W<G�%�v��ڕ�;�L��j�3�e��wa/$�me7"����S�����D���T-�&�3��m
��\+��5�����\�v��� ��|���7�:���X�E[b v�l�F��U.�����J��!�4�a�E[Oh��e㪳ק�Oa��lBbgv%���÷P�(�I�hK�,�b�:ܲ���Y@�g
.weٺ�1D��<n0x�F&kb�-�_"m�?G*�}��<�N�Ύ��8E7^]��F�=�#rr�EA�{���bʘ�L/����ԻՃ^������<�lg{7' �,�����9ܽ<<ٻG*j��m��:���(�ɝC�cU&)���
쫦sf y���єV��t�u��t����Ep��"wg\UNݺp�e���)��:�B�U�Cq��;t�{ӹ�ڂ:��J�[�j|Cd�T�������[C�-����-�6L'^uD˓ �������b\c��!͙Q,�uc	Y�Q�{m!���f�L�1ji��`.-�/����ɻ:jٹɺ�s��`�rXMlr j<���7�t;�\F�:s��L5��6qN�&<x�>l��O�{ː�ȩ �k�
�5D���p!v֯��L|��2���r�53�&�(�hI.H�do^�4kC�������ZW��9�F�YgA�y����������ܚ��;����':��4����G�i��z��,=�:�ɡ�r��?��$0��7�˗�S�e��T�:�\�١�;�y�vp���h��{N$^"��i��QG�a=���u��/B�{l�&a�Ɏ�)�3I����Ӷ�8�UEsبWP��.��i��A4i��z��n��6t�d�����PBna�ᵘ�TS��gCc�x�ӽ�ˎQPa@:���]-ռ���{.�ϣZ	�(
����%3wX���]��O��-fvLu�Y�Y!'֫�*���a���
@+ �� �Ҳ�O�W�x_u㮠�=t��b�pm}����ЗY���qt���%֘��7���ih猉q��̌Pq[ܻ{�y�p#�#{�5a�[\Λ9��u5�Ύ!��ۼH(�����T�{���嫲�ja�
��#;���2�\3G�t׺^�V�q�N��Ȯ�J�%��|r���8l,��}Fl�]��tu�8��T��&`d������������zK��q�74v������tY��p Q�I*/#B���!s{�g<[�V�*wVi�쎸x�匚�3�������s��G���6��n���P`^���>���{P~�g�,�����ըҎW�;D�mX|���*��2m�\܎�PW���"�%ܾE"^�m�T�H��֐8���=��ˍ������dJ��3c�e{������:�ے�(����5��&�b�z �^i�_>����X��5�%�ʹp�e��[��i�*C���PxH#Z����sP��|�����;��V����6v�Ϥ���M��1�����S��6���/x�v���Y�A{�����\��ǽ�K����_8��\=+$�Ů��:{�{h���zכ�wk.P̳ŵ�`�ҭtrɇ41D�����[��`u�-v8/7���pE�l9�t�����C_�P䝵1�Ui��`�ޮ�����V ����'��ء�*�㯘8�k(�s��1��� ���9+n@�9۹�=�wV��,t�F[��u.Ь�;�bĳ�sx�����:w�E�0��o�9�Rw;.:�3p���0����ׁ&{�{M�K:n����@P��LJ��<b�Tl�SM�P���u�ǈ�g"�k�'f�+*�r��r�R�4�f�2T�5���v������Wd�!��Ҧ����7�.,՝3{CS�"�Ox�ش@�����M����#�0�U��؟'r��V������dK��&+W`�yC���n�A�h)��[������\����;t����.(Z�/N7���;�34�5�L;T�7!�VA�]�F��=����#�d�A��5��$Y�4�����Plr$�ͽs�� �����C�p��
�U� ٗ�0r{��ܷEstv,��w
���O����"W~T�8'�4�f5�T44{@�v��ɗ��c�V]����U��2�cI�<�)�w\�>ex�j3t%_I!��Zo��·��7	�'��ѝF����%� 1�c;<�.W�s�)o.��[�o�C��ܡ5f�$P��v�:N����PzaqX���#�������� g1�3���15+�a�>߾g���.!g~ߴ��{��p��M�Uovy9��2��G9숝�&1N��}����C~����	r�(���}�;Y���3締�)H�x��t���x�f�e8��p���u�&Nв���rf6/�ޞ����X;���qx��dO9����l~��9�j��הeZT����:����S,�����q8����Z�v������\�x����8jeh<*�KX���RNd��%�-��fEXWhh����} ܭ�Ϋ�R�.׃L��)y.�J����|�7��}	�K�R�YI|o�>�{��̻br���u;��l���͹�Mo=�%�2��m�;�c�$/Y����wR�j�~hqN��vB#�0��&"�w��� in�|��٩��M���B#��y��x��oxG3�[p�$�
�X���w/_B���f�H�;E�	�x�{����&���N�c���1���}���u�og:=��}+�P����Ύv���n�30&�ʻ݊��*��%]���p+Wk%3�M,w�Җ���~�<��Oob��|�7<ƫ�N�sX��y5��$���t�ի�ըK�cm�DZ2�{�.�w�7p��j\���tP8۝6�K�go%_�r�o�ɷc���E����Y�;�Q˻Uso(`���O��H�~�wK�$�*�Ч��B7��of�/ J�;{�P]$���G�k�YA�ܸ<1�e�+���p|{DZ�^������7�SAOF.�T$�r��>(�=F2ށf���7���u7�t���k��n�xU�G��a�ܗƃ>�j���r�,�]m�D��4���oV�u��a����g�\�m:�����}0�d��?-n��.S�'죺,֌O�����G4x����ڰ��Kq��`�[�Sa����p敚h�w��%).*���"\t�z��WKsE&� ѬFVq�	��� ����Y�t����B)6v���Y˧���D-wp�7[q���!\z=#Z��}���d���$�1�Q���0矑Hh��o!En�"9�7�	��w�_9�'�1Fn;Z����С٥�&˫r���?57�E��� n�y��Fa#�oNY�U��7�׸����8��=���.�!�}�{�ָm� ��N[����s�;q	c4���s%l��R�+X���qNaS�zN?c����}�ŅoIUJ�2��Of���y�{ۦ��1���s�o���l�z.�q�R�!O�{XP^�[��d�;�;yvS��P�Y��>������Wi��MNZ��f�Z�s&�"�xv�f�}���k�o��T�޷v���r�C*R�0t���T�+��z�wVE��%e��wXG�6j��#:@ⲗEiY$�yh�'tΕ�X{=Уޞs�h��9�*���+���\�`�w�J������7�wM�e� c�p��rZ'83�����7D�rm�O^��Պ�.b�'(�-�c�U�j���69�8�u��J�z"NŵQZ6�mJ��9Ckl���)�F:��n�`G��Y.����Q�\ݗnU�������d�b�^b�<�&�W]#4+ѰL4�=i�Em��])��>��0PP���qP���k��/��{K$�W�<<�<7d=�f����@�߽��|��s�q�o��Ǒ՞�c0�<}��"�� �.k�����+�T�m��ެB4U�"wc��mRe>�=�R\�<��냎e�-�/ֵ��.K�w��f���9i1�@+c�r^�+{�z�k��lWT k;Ō*f�'0�z��4d>��>�����r�"��PzB�{�]o�m5ᗔ�x��{=||M`�գS�[��e��N��M��$�����wm����3�3-��)�"���]��n��=��Z^��-�ʖ}(PRn�_�p��IWi�J'����
��^|jg��rҗ.����k�������|^9[guY���$�L�^��dv���گ�b���q���{����!�Mi�BY�Y�f�΂>�5b6S�=|Qn��2�K�9Ȅ����5�����H+�ש{_ae�ْ0�|�Q;�zT;y;%�5��x��cj멼��Ȼ��}ib&�-��^�.�IR�X����]z$D�..r�ݮ���+L�Kv�y�9���a�B1��a��f���r]�T�7��I��q5��92E#D��I$�I$�I$�I$�I$�I$��GnK���T�-GMb�����9	Sl� �`Òmk����F��-���g����!0�c���(z8,׎�"g�(Y�y;u�M�(sR8�^n��\rম9ÐuV.
{/�h���f5�i�����;.l���xW%Yg9|�U,Ν.�uZ�Y��:�o!�q#�Vq��Z  u-�������p3Ǿ9��f�����{Ȓn�k�<ޒV������u���aw]ySN�v���tZ�=>!Arp�j��Q� ے
�r��kb�V�f���ZT�{�#�eW�9�.
��{�a�r�<_\P��$^��t�J�7����k%ԕu)]���R9���Д���}�����L��Iګ~p@��Z����f�44��f��)0+�s��-B�i��9
C�W��{��oK��$,�D)�H��:�tK�:IٝR�;���J��+�ڬ�Y�.�.��c�	����]��wΥ�hh��+hoTp9�q�X�At]��ӣ��ڟ������U�}L�}>ÿe��}�����I�C;S�@�w�$�����V�5�q!	$��O�5��y�>��*��wm[�7o���k���	��qCa��'��1�����͓��9���P���&;�2�o(V���ͅD�m��@hq��.[��w	��{�`r���|���te0����� �����m�4�VZ�=R��9̐�)ý*�'[7t��iB&h&�i.T�<��������yJ�l[oX0Չyu/@3!��L�/i���s>/�}�2�[���n*&e�0vA��fKGI篈�v��x�Fg��<�íi}���iq�*�]fͧ0�`�)�5]�"�W`�Z�y�Qp��q�Q~��_� 7x�0v�~�
o���^�pq9��ߓ�Z���m<��IL��G����8�A��_W|�Ǣ�{�����r���^CIi� 5N؟������p��e����yO,� ̴�/j孾|��W �x�^Q+{_[�m��6E�ƭ\]��=��g3�E�M��1�I�p'����=��\V.�j%��;���E�����G��G���Phw����n��<�Kr�G�c��d��ߺ����ox,��c��U��ўĢ��G��}Ò_���5L�jㅼ��g#�w���p�>wJ�h�ծ����K��M��V��K�.�`
��|�@y�~���g�ѣjq�Uv�+k 8q�Mw`�4���w؇P�^U�{������ڍ
,������C]�&��D�f�al��+a�A�6!��dt8����PQ;t�c�{��?�=�xp���p��y��ϲ���S��6o 2�ҙ[w��8��<^�"���x�0e����ݎ͋8���p^�Tt��p���]��q2���Y��3Y|4���HW\�e�}c��%��#�:޿�e��-r��Fd��Y���K���+�B��e����dc�$������ �n;�,!̓[.�D�C��9Ól�^a�u!�։Ntf������Vns��H >�<�G��z��]�p0	y�`Ģú˼��R��˓ᗽ`O̟eQ؋�g��
��l7�m���8U�v�s4���U}r���Lh���Iu�3�T	�<4R���0�0��}G!�[��M�SE�:�8�p�;���f�qlȃ2�tR��XJL��1���5X�pe�mu����e ���i�ȩ�vO |h�`;��AsmRG?2�S���mٔF�������$�!����8�4��L��ɔ���w �L�le�QV$�sa�N�3��ɹCS�uF37�p�e)+���� �J�!��>Iy�d�
ъb8==`��u���_\�"�bE�Et�W���Fcm��l;��^������L�@����z)�c��9�w�b�a��5�����pm;��v�ڹ�F{ɸ���X���|�qn.������;��6闔��m�R�k����1�����ո�d0�솭��I/
�&4����u�;`P혐���D>u�����(��F���3�f%{�)eb��Y��uDk�Cz1x!ۆZO��	����op�<�a�am9�Y���2�B�>.��p�Υʲ���Q�z�Kͽ�J5�C	޾��?���fE�k���vfY�������2���\\2��o�D��|[]���j�3�<�~s#�%��r-�Ƕ��}u�Zk|��EB�5��2�a�PZ9�A��j;^�;���,��Ih����{%߳��&r�5�x~�M��)݇�K�$h9-�S�y��9&pc"Fh@�:x��gj=�CL����z�y��~E��j�:N���׈tnK�(Q_���s�n�KJǝ�]���;��e��4d!̾N�����6���P3]�
tk^=�\=���a�E��.��I�yw�w6�[�=4y盃�=��/YP��Fd�<���=���ȱ��'�=��R!;J^q���H��<��J.��q���t�֙�����������f��ӻ:�Y�wU&f��&�� �k�c:y]�c�ǈ���ub��8�\�3���Xͼco����q�b�lb����D愖'������Ai����U5�WW��|��W~��nX�([��ك�d�hMD36r��ni�RW�������i���#���.+_m���Ч�fI��as���������C{ŃlHz�Pٳ�_X��q�B����I�`�!��X�o�C�*W���8'|x7��U���X��^����T�Wy�E�)���uAu���]o���m�f�h��L#�ص�cRlҽIeA]z���H78rFI>y�w�~��Q�84yG���7���t��9x��{7V���;��>6b�Rv�xa۸��mK�|m�5��A�E�Y���	�[�F�1w;�	$ؚ%�uJD��8�~��y�J��״�7�$Kײ�wH���2�5Z\�.gUmfDk��Rɽ���W��r�hm;y�u�8�mo[u`�s�pj�"�Zq�+:@��&�]C����]AC�D�]Ƴ��k����*r4������=��������^����@��;���ڃi�O�%���.�i�3�td6:ڻo-��^�BjO.�ܠ��Y�Ag��;e�����|�Ru�R�%��a��{���U�b��n�Q�<�úۜ�{LJ�=�:��2wrF[k^���2	��Ϡ��@�I����	1����|>(D�}>���vI�?=�@؎�wHv���C��S{Bn�4��ݕq�?�N�<�/lL��J*}��Z�����J��$��*�������� �����q�R錭��w����D�(�3�'I�>z�ؚ��׮p������>��t8\��Z��!ڛ�.�;�k��h"�Q��E"ot├�v�J���B��+o8�������d��v͈�ʱ�o=����qڋ�1H`%��9�{��/rB��$8��p��{# :<�5�,���_��K�N{�� ~��/�?6����eE�\��Х�D�E	�;%��qD���o:�|�B%2$�L���T�Av.t���=�׌=,�Kl,�#&g]E����2�X_����|��b��dW8mt�v��\��*6ޣ�,�N�ɼLEW�B��{�T(��1y������Q�Ks4�v�#�/�=�6v>\��������3���b�.��$T9%������m>rN��0blP��\v ���
��|u�ױa��*蕍
�H�`�{��/��K ����r��,�>~��*gߏ���snmb�}����A
7���e��9�[��u�X�G�f́r����7����m=Lht������Ss���ΥOg޳y
K�25sߠv�e��nj�o\\�>A��6����'���;�B�6̮���nV��b�7[�iIv,�[�f$G�zޓ�q�JJq�bkFl�q/2b�>�ɴ���R�vۈ�Z�#�M �v��y5���"d�u���i'���(��Z1�q;Y����J��g�g��ʐW�����k��S�����j_@�/V����UO
��O�s��Q�eb�}x�GTL����z�!a[~�������X�k,_�����h����]��^��=#�$y����c��׍I���ņ�.V���}5����ś�X�<�4R�Լ�����|8� f,�j�E�X1��ީv�'YS�I�d�:c
�9]Q�}�8�Ćg0M�1C�ue��5��z���fk*h�v�M�}����4�G�n�����pļ���B!��?]^����E��YŦ���Wx��ԍ��mY�O�}��c�u��[^���D9���+��g�6�����"o%��o��'TX吔#�>���^��QβߜA�}��s�	7���g>i�J�����U��&Ue�ÔA���r��.t�5��ijGX�o��}��\��d��l	��|���U������S�Q{eǻ۠F���m8*���Ǳ�t酔��{����ի��l법����E�XP�Ok�фI��c�v�V֑���ZHp�٘�1�{^Ƨ+�3�v3n̥��ܡh��Fb/����Q7�������1�
|�)�۹u�Z��E������t3A���l}�{���N��ѣ����ؚD޼oq\�_�[�ܶc󹵱j�$_fC��w}wF����ON�L*u����^B�����sF�F��yS T'F[9>��Y.5F*�0^|��E�08kNqΡ�;����'hn|�}^��9�z��FQ�&�ø|��<qVD78�4��_J�N��Լr��G�KJJ`��j�;`f1�S%'a���*���>���g�Y~�r�{�-b�w��p���U�R�z1��[���]ȹ�]����W�%�铉������vIOt;-�����^ũ�������j_��U2���w��	�
���WTn�f��\d/w
z"ECo�t2��H�Yo�7�hEt�࣎���v=��c�:gk������ͼآ�<��D���1ov��`5���9�$����Cjaѻ�OR5[��s5,��{�7�GFD������S����~�ֲ@��G����Xfz��Úi_l�y���r��쯗{���Ԧ0&��w�I#�x^=�zAaK�Ř��g��(�IۺB~m�*!M�(��3֗=k<Ju��������D�w�����`���I�Xw��\�/��f&��L��<�#ӕ|y��Q�\��9&��u���6�kA����J�#�b����՚�޺�κ�<ܰ�o+��>G6�v�s--��[�2xW2o�:C�S5,���0v�pv�a�)>S����%�����˟Y���_�i�X��߼TgDCO�䩔�9��>(��G(<�͘ڣK��\�<�������ߡ�6�oE�/ҎO�JNhT�9��Y{b�鋫�L{�1�<oE=��>�^�[Y�^�΍�bk0��G�q����!���������8&��������5��.���ewO,�_�����r皺���:�����ҡ��ѱ����e��ׅӥq�r������E�8}�8�e��x-%<c�F���K���;�Е���m��#��];�v�Sf{�~�*���M��~J�*�s���7�ǵmKu��A	��`?}�8�O�����@�L�� Yr�;r��]�0E)���A�3�Te�JH3Sm�~3ƽ��m���`ԍ�9o��̔�9�3�WR>�zM5��^�^n�ytq���A��z���53�������*9�%�f��Bǃ|��3��t��Z�ոp��<�c�4�3���{~K�R:B~���P��^���{f����8}Py����{�D8J���\����n�N�v�Nk&���ɚ��dGj�w���tK�H�؅u��P�>�X@�����H�pى�ᤵ�zAq��y��с�t���T��}��glI�);аm.�����JnR��Q�u}��{�v��Ag�2�	�<�]gջѝ7�;�C>��ڷC��:�ppm�`��s��#�%��%*�]Љg�L�n擂�&�u� �2���'3hښ)[v=���뷡z�K���y��O���sb�K�I��v��Gpq��
�Wr�T)]��ՠ��A��!�Mt�8�.��n�r;��4�Iߏd�|;�+��.���gh��N�w����P���t�P'E'}z�6�e������N���C���Do�Hӣ��Ľz�R�b���%CNHz�!�w��aO�[|�7����ØͮvW�̼�i��c-xC�fK��ɿlsع���� &Ѭ�����a�8����x�tK��x޷y�Bo{�a��ɏZ�oXJ7d#Y���v{�N�(v,�έn����xR�&��й�%�\ɯ���ػ�̮ޠh�nd�{An�u[��7iK�'�P���hI����n� �L̿2NE�0��Z�I�}v�-O��#qfqtQ��=�W�*�D,�ɒc�'�s�V���$AyI	ha���j�v����WB�%Д�/IL$"�7
�̱]��s�M�*�h�KD����IF@)��ѳJN�Q��W��h���d���.�����^Yabe�����XJ��(�2f�Y&F�k�NX��Z%�^�D*e�2nLܵ���Ó=��Y��V����'�Ow�9���`k-F�/J�E�=W[=���g<��H:f��9>��-����^V��C�	�Ə�}�g�*�>[=tv�(C��ì��N�p��
�K�ה%��vl�GyL�8�wp��k��eB�1��dS��<R�뛛�:m2�j(d���ޚ8�3���1�$i�֡�|i_p�T�9����v���C���^��՝:�KZs��#V����%�<U���Mjwg����P��V�y�����z���Za�5�`���8cj��xw����W�j��;�ؘ�O�K����2�N:�8��*���}��@�9W/k���z}�"c��P������,�}�u���}�����Ӗ���⮐��g����z^ohD2������"}H���;�Ko����|�b�����Y5){|Ma�ޡn?^��%m���4ɘ�3u�c!�D�o:���^���ߟ^����[:�'uM��kv�^��g,�5�'�+�Iƕ�7Ƀ�đ�+��������Cw���UΈ�d>O�`��5*v`E����PG���!g�kgNfģ����b�_s���Tnr���y;t5��g=��_{�%u�8���g�3���>-��*�f�=\aۡ�up��S;��Pk_��2h�ف[���GWy;�Yb�ס�v�K=��a�e�CҸZ�/ʭ�Ԡ��Y��T�rfi���u%�٤�n��]�
Z���}nG��üߤK��c�U�^�
�������ݝQ:AU��Q eDמ*x�瑧��=��+���2��<��+�D�f9Vrk���bru��!�Øe�Y>���E��\���iSJ�IIP�#�	�����>\�{���F���b��Ce3�H�A^�hX�6-hK�X�"�fz��7�ςG5��/�)�`�T>0�`^h�����ŭ`�iP4��%\���{x�m%ƒ��1#���A֑�#�	Sa�*�Ɓ�S��X�%>���9��s��"�����̹$u��V:&r�+�Ǟ�?|-��9}����W0���zM�e�|&�eIv5�e��W�Ў04��cUP#�!�9�J�y��@��O��\k��"6�d{k���-��,HlJ�Kϭ%�%�5� l�BH���#Z�|iP
ؼї�ds�/��:ΰ)�fA�!`.4��S	i�h%�li)a� �糑�W���-bց����<��]���KK�%֐��0�/�2�J�|g��{g������hA� ��I�H�K�F���E��4����M �.������4#Ya)i.�L4�G�ZÍ$C ���y�clA��|]s�S[��y���4��A�b]b�cI�X�;�rG�1!��[��3�ϣ~z�D��1%lE4���T�l�y�-��$�4�p�m�Ϟ�̻��Z�+kZ0iy�4���`H��Z҆%�]ic-��4���T|�WϞ���� �E�#�<б��1.��a�Ix�@�K�bKV�i#�|�l��(X��ׯ-~vه�b^���ٻeҘU	SR�)x�C?�ʻ����v���P��Ќ�T���I숸��u�QaM!�i��|iy���0F46�5�� �)hbƄ���^���DW�iK �IP��`��u�IC!���k��Gƃ�J�6-h|>w��w�;U�_��i����Hڀ�kA-y�q�>4[��2��>4�6�_���q��o+@>4�i.4���4�l���[<Э��%�O K�<��/�|�^|�ݬ�-iPh�%�m(�D4"�K��B^g��)h� Ɨy�_�x�ܟ��H%��p�q�3X"�<�������	[@@ľ0T�T�e����7~���u����p�l����D��hG�ZC-�����q�S_�XlGϞ�D���%/�)�>T$k@ړ� �� �GY�� H��0i#b~\G|W~U��y�q�1(h0�\�D�[@�b��0WP �k�Ga$Oa%o�;��~�z��$� ��IH�k
i�2��B<����aʄ�`��$|�����r5�O����p<���o��n���\��3=�`��ޫ�0aR�\z�18���u��*2�����X�*i,g�`IS�.4/�%L]d�%,�� ��A�y����#��K�P�kօ�cBV�:�y�alZ���� �kj{����6�!���>0F4��б� ��[bK�i.4[A��t��m|���e46 Ɂ"6��?�*`A��w�k^7쿜G��6PS(�~j�כ��q��=w)���ޙ��}�a9_���c��ħ�u+00ե����P�����_K^�Y��-�y@t�ZF��)�����d�^�o��E�]�;��s������,`��(t�C��w4�}���-E����?9}�u;�]�n��8�G��[��{�s1���ɢ��"o����d��,ݎ�MQ�VEC9ΌҲ,/�?O�f�||���ǧ�vZ]�"��=������MY��z�:�;� ΀�Lc{���K��F����g_��l.�3�'�%Z���GE; �wd��!\�@�b)�o��m�;�B��v%��XӉcJ���6��c;k�-�2ULv1I��̿y$�Z(t��rQ�ȟ���{g��kة�ll�݆��U%��H�_�G���Ĩ�_�_G`1�0^m�Dj��e�g�ՍHia:Q��o�����foȿ g��t�/��K�{����ϧP��5x���L߱g�z���t���2�}t',��M��%��r�?�ϧ$��^�%��m�Ｎ�q��"��pl���[�v���s�9��|���m`6��ر�a��cd�;��*����hI��!�O��}.���W�d/a�nn���',
��$�U}_}����b?�o�w܅'?��#G{��dv{[G=���9�	��py?������#�>0�z�P\>�@��n�@�)v��Aoٳ��I��ع���e���س�U*qܳr7_HEm�,M����L!��u'O�>���'���ߛɾu�>��2w��OU<�]-{����"\�K�� ��V��^��(⣫?1t�Dln����`<�S0����Ȓm�_����m�t9�[ws�`�Mj�ֵ�QǏr>� R�kT�ny16��i��6:����o♘.v�Te�/��c���Q�J)fml�6�yN�JO�Líκ�̗�`�q�ϑ��^o��e����ti莧X����nAD���31y��w+��P����1��ԦZ�i�,��@��k�4f�g��g���$f��$o�_��nw'�ۖ�nV
�=A5����2�Z������T�s˼��J�s{:�;�;���Q�j�c譞3�`�W0n����x�N�%�I�����Zq��Z��5H�̳�e[�H�L�K���3���|<���`;��o��"�pUË����]�Vژ)M\�s˳}�Oz�4GMڛs(���#|�<#�b��G%�ߢ���4	������=�P�Y܂����v���Y��\�p��=�t�%��!��N)#�����=W�.��Y�
&�ǵ�����nc��y����.���sl�(���JT������u��Ż��� ��Gk��N��~�r�B�2I!D1����O"� �\OW(RЪ�1��y��L*CR����BO/*��ҴܧH�+1��]��//O0�Ϯ˞��dI�� ���!<���5D����4��OO,�R���)3%,)#u�Mʌ����5L�<J��J�"����$Z�p���fQ�G�D&��:"��)�&s<�Ы��\�@�=u\�&ZRa�^U:�f��bfy�AV�UPb	��TT%�'�ꪻU@
w�N���?C�o��FA��AS:�NW ��� �r�{��\����A��Z��cA;ڮP�������}f+�b�a�=W��Qk�Dcy�o烟i�lk8,������%L�Y}��5�Nof�q�����j�+���S���#O��K[�
}{�R�[�v;���Xp{�����^��{.)���2!��%�څ��w[/����U�脥�[��UX�-a湌Q�㒽q�[ �P	���ڏ�ߠ>���Ṳ��� m���
�,u��㟻���꩘ϐ�O�St҉��Ht7�EAP��th4n�&�2����z�.�BZ�1����۹�=��9Qz�� c�n�^M1}�H��嫵�3[jƅR�J���Wg?��}䇷M�|�Ľ��a΃6�n��ƹ��3ZG"��%������_�\�5n/��ǰ�����œ�>y�������}׽�V�a�;��i�,ni�Ƭ,,gCr��T���G*�صǹ~=�z"'06�}��쯌\Pe��QR'J�cNLf�ĦM	�x�l�1���v��!�����ᑠ��]���u0�s&s:��6�s��Q�t���J/1�С���5^1�x�GnejoO;G����P�}�7l>���cY�Z����y��Iۗ��6��<���Y�&p�Υg�˳�fC��h�״EF��[vF��˚lJ����>�?-�Y��M^��I�BT�(��^�<��D{��e��pv����y���,D�w9����>��t�o�`>L��D�گ��l�,�=F-k��5}o�c�g5^�4�=q��A^y�c�ܛڜ���ߺS8H�3�0������]V��:���oecI>��P=f7d�d���b���o�5[F;��d�
�ß�����L�<e��=Xu}��W~y0(��8�Fz˂¬�4�#�ɣ�<|a��Q=qf�f���S�����G�=�h��.�c��*�1T�Ȳ0r/Ec�@;������3���FԡS&S�zo�4��b:�����V���Ē�d�f�o��#��A��;~���;�3�i��P~݇�K�̼�-��;5�����5�/MeQ�gz�ñmy���������?W���a?|��������,S��o��j�ֶQ��5݅�A���]*i4�v\LL���r�䎶�FV��^Oj�ޏ{���k�}��8���#R�\��w�H�%.�tNּ�����v��T���8yg,OR	ߌNN�OV�!I�Y��%�I,L�Z�ʟ�s;�|z���e����kϞ�2V�+8�ɒ�N��6sr�4��N.�O�rr��龞���%B�_(���¯|zN1?����g���q>k���Z�� ��X�,һ�Y�+h�;4��Fv����l�+13j�j�]	MH��=�F�����Ƽ'"���灷:zJ(Th�b���y��fZ��_y�7���_��������a�ɀ9��0��2�!�aE���]V�u��J9�&1l���hCB�����D����s�<�9�+�y�����I��u��y�gVd�tפ���c �/�����_A�D�c�%�׼�h$n���'+��V4��l��#jm�����T�ii��P�@PC��.]��7?*�������"�ޫ��T>��P��6��:��1J�s�$>y�Z���P"]kՑ�QuG	v;��<��:��lr{�^�z��ћ̜]�\��ھ�~����k6&x�/`zq�EI�g8ɠVt}��'v1�kGf��yI���3+�7
���\h�3����s���#)��A�Q�X�����]~�}z�K]E�m�h�[t��t�	.���i�OqV�c!�`���ei]��ӆQ侈�z<R`�dkrVok��A�����f�_����|Q��A�yԕ�I5�c�A����G��{�*���2��2�sm&v��n1�X�vU�eT�(�6d�^�<ˠ�a�P�Q����5��76��!d鼾��_�{����l���o_D�	��&o�td�7���囨�j��KF`���*����"���>���9�����쫣/��"���[�|��9�����G���=?l��4k�p�ϔ���2\��0�WЫ�I+�;�h��y4��/~*ZTV�?� ���xt�I���uy�/Wt��Ti�>��^�Pb�q�r(M�m%�qB�����I�K��y.,�)�*�q�V�֜#�4�
#B��+;TB�Τ`{�
��������#g#㽍�&�OT�:&�a3���q���w�1p�N�W����U\>��k���o�	��TF�79ұC,1ۮ�V�1�����d����q�~堰F��$����v��@C�^"��n�.�n�o3�}�Rk�vbor�<V�.�	���M�:��k�ߴ�˿n��g��f7�s���p���%s�2�n��u�z+��-��qC�Ϋ����n#N��쁞��dX�WxϚ�`�ۛt'8tD:����o���Q�r��Bn]$u@;gr.�ró�7�o���=~�<T�\Q�˘P�L�6}�bԲx�p�b��A��͛�����2��]�I�5��_ �$�[Q����î��QR���3��֖'Xp�*����7mn2�K�q#�kZ�K�Җk�"f�L�~<^��[}$�d�e��;(H�ަצ	{��@��A�ۛxO2�U�����|�S<��ra,�����}�I��fVIY�'�_I��LR���c��[�ߒV���J3�p��&�5��A�
�H���;�Ӎ��w.�c[G��m=�G��{ڧ��3�`�8��V���S�:j37��Pگ|����Ă�]w)
M ��J��Q*����L��;9�Bҡ2��/
r�JQ�*�MqLܤ���1�O*^��d��diW��@̨JԃL,��<�t�������r�H���Uz��U^^uĊ�/r'�� ����IL
�l�J+�R��ԕ#SK#�3"��\�5��J��2H�ļ��J�Ф�!�lno�u����ϏK��30�����'%�D��.~�U�W�9����{h���?��9�{y���4Jqo��J���H�]���]ƚn�y�]���ߋ�FϏ\�����.[�{"x��d��Yܓ~^�z�k�>O����3ap�z�v`��A�oL>���qt�g�����O4-�S��'P���H�STG~K���ۙ>m=]W�9MD�߃t+�ߥEt���ҥ�4a*Q�\'���y�˒�x�c���{�ϋ��*�}�kvn|#��j�D(}�>��	n��]�&�,����Lv�>�8sܧ�.;�d�jT^�詰F5�)#6�l������{ �9��a9�u�7j�{�<�q�w�j:����nIϊ���)Z�gW��)�~�����n�?r�w���z����XP�F��<��L�Oi��3]�]]m^���'����j-i-�Bsvs�o �7�)�X3�K�Dz=W�+�����G�Y���mſ>�Ǜ�;S:��l�}םҤ9kM�3p,!�t`����z�����24������J��c��{�uչ�W�S�d��%�Qz��ͥ�wy�[�� G6�1ݔ�E�w]u�'����Q�^��ԣ�[H�]��� f��W%�`�:�{0󼟆���/����z*�,:~��+u����<߶e;�WN�擊x�f�زc����(�JI8����{ގ��X3�WK�W��Bw�I=՝hUں����au"Eq�ո��4���x@�����Yx�#7+j�b(��d6*0��>�c�r�|͞?O��p�~�b�>�b�
v��Or^�P�?]pj?q ������/��=	���d�_��S��}㵞Yv�y�-��XE��r���{�Ϩ��/��/�.ߞ4�	�j�S0(y���H�u��8}f)Vt�5�V���,v�q<���{�}���_t���F|�2�^k�m��8��+6�a�ø�1m$��T��]�+M���g��^s0g�J��G�U]��:X��X���Ή�46��6�`�&G<��K�j�VS��1�(��pgf5Tll���r��My6lvb����5��[*�{@��Z#WS8fLk�nMћV�/���[�3�ڣSGj�R��eh��n>�/�����9����{;9��-MP��v- ���8Sz9SWO�e���9�)�?�-x�	e�}�|�N2<��ҙ9�?^���~��$��9�4��c���փ�-<噶g����ڣ����
5tB�M=��E��I["vTZ�n�.�7X�Dg��]y5��CE�f������t�]6�p�"���ԛ�"�su�A���C�2����ADJ*���o��D{�sx�����gv���b�nB��b+����{�b���g���1R=7.-QC���:���;��e(9���VV'<�����Say>��YB>g�όu��lRfds�y�����]���}�\(���n�[jLֹ������m��W���U���O��7&�0 ��!cc�c'&ˊuL�O��3�l!@�l�y5j����+0Q��~�2d����)��� �Ӣ�����%Y�y�Wݻ���V�͆��)*��k���s[�4ǫ"�a�7����k73~C��d�gű�K�� ����NF�<}�*d����Լ���=ʦO`�c�q�鷵���9�w�q��o�<��񘎜�ܯU7M<���s�]q3����k�Wa{0���-�q.y=j�W�;ﮝ�������jK��l�y�$�
�:��5�x�fI����V.�o]���^;�<�̧6�o	���Y橊{�=$�5��[�ۿaO��q;4+Օ�71�ߩTfbw�����gӬ��.�Y��8�8������'��+~��*6�+�$Q3'Q�-�e5˚�Ξ��Z�W(C��8d�\YN7~!$^o��f���5�E�r��+�2��sC٧�W/�>���n���G_�砼�޻��y��g}x�m�e2:��/�AF�v����|��%��
�}t8K���ؿ�X8+���{���--�7FQ���[��� i�O�&�T?3�\ՌÐC��ޙ]�S�]c�J׬����[m棽���w1q��A�|��>���my�g9�NQI2�&`��Qn�:���>��P�b�f2_X�\�ϔ��.�Ƚ�*a�eCuі鬉�\dԞν�;�����v�Z�:'�L{���g��	aP�� ��z������y<����/,8�9�!�gy��)��}��s.r^�(a�L��a�uɫ���*L�yBV;�x;R�#��d���n�:�D˒]2^lq���nW`�1���o��;�V�1�=g|L��>�"b���oe̎���h�����>�݈m�r2�C(�ν�_��L��;D?T/2��Lc�w�<�}�C���&���x�Fc�۬��0
9�c�����
ۭ�b��8�㙂ݲ�N��Q�99�î��a항Y�y��[ƭ�(�A��N������q�_q��z��Sν�����+�'��
����p�L~�3+k!.��1��[�)�݉�J@VDn#���6�$����_������B��Or�Jb�b߲�`����pى���5}|�9�¶�Pt�e:�����]�{���K�J��z��N�_v4�\Z=��7�5~�m�����AVZ������q�zy���a��H�V���+\}Ӵ�����d3�+�L12dW��5��e�/f�de]{���.�O��P~�_��I��ֻ�پ��o�ϐ�B���w�F��˂�smwX���X���,=��8v�c��#���,n�7���^,⬽+�b�(�ݳY����sb��s��n�����2�9����CV�~���W��w����d�\}�8����|m��ݹ�
)B��4����t<>A�r��]��h�����HN�n�+SE9�{�8�uJi�����xv��ܝ���<�.����X���-�qGg��MF5q-1��V��0��t���^�w�����ZR|Ʃ��꣖�[�]>���D6!��Q,��R��L����bQ����.�g�x���g�긗�/
&�y'��:���QQ(襞QyCP��x}�'g�I^�$����ByN��P��^9{���*��O/p�r���<J�46��g~_=�8͚o�8ov&
ʍ�.��,�.�8�n~��U^���������਄�u/�¡̧w!N��z4-��ھ&:�����r�3�����|w9�޳*ĳ���eA
_�s����o��/���#×�qg!G`9�k���ߪy~z����d���B2L�T��z}Q���1�`�dq��K�d�z���;q,��j���f_����͚s�[q���8G���|���g�����|e�^>�QRw������qza��V��P�wr�I��J-n�['�W׃���S>��g��-�6N*��f{�{��,s=��D���$M+�YH]h�:�xb�Rq�t&�Ȇ�V)p]G/wwc�;���y��|�\̐�S�B*aϬ��6/9�>�Q�Qs���g�ɜj�-�yegr��g-�0u���k]�C-�������Q����l0k� ���Sҗ5+�Z밶�*1W�TT n�ݠ>��~�������󾚜�\�c]�ʦu��ؖH�v뷓��[qPq���ѯ�1��1�5�G}���¢jղ72Mv�T5]�Y��V��U��쨞�>�r���ӭ���>�y���? %�ܹxK�`�\�˗P�uv��'*Q���`��9������w�4s:'w�7.�C�7[�LS&���һR]�1�����[�Q�K��� ��;�>>3)�%���yۉ-�aا�q��{�<ny���[�я���"�
��G�G^X�u�ſ$mnK!b�'&v��E����گ�-����V۬��t��
�*
�:���&c���Ĭ�ґ1�환t�:E�}�������d˚��Kb��8m�fg�b;jg��e:��h��/
�����.�2*<� ���L(L��k��ό��N{��T�g���mMT���G_��=���˺��.HX��x��̅�5o�9እ�kM���h7�)��ꄥ^���V�������/��S�.5��%P�BIF�ǻW���i=�K�>s��:`D�ف�T�2\�,�L�TC�r�GK�ꉞ5��"c��I�r뵆�¸֎\u�pU�e�k��I^�H�^���Օ���Y�F6S�d���� �ʃ���Gy�A�c�$��K8�>�91�]��v,0Β��`\�U.1�TlW�;1 I���E�p�t�j��������C��vx�;���3�G_����:f�ڣ�8F�f��:�g�\C�ղ���_w/w=z.x�!ӇOZ�_P^��_��2�����k��n��M_/Q�r��:W�A��+�p���l�������b�Q7?*�o��p�_B��13���*��맧��p�v�j��p܂�HQ�wbF6S8�|�6v}�n�<�_�-��# ј����_"�
�9׼��Lﻼ�lץA�ܬj̓��j�T)D��"}���5�G �E�]z��J���0��B���j�/�߶aҸ��^��P�M���UFJ�9��l���Q
^�o��3σ�z�	�u��y�1���q���{����^��.8t폸��R�υ]p���,=�OJ�u��͉9�I�[���fk���g��{a�P�\���)������D��<�'#I��nD�728,_�LF����y7���D�5^�N��Ӂ��������9Y&�ن�K���O�g���E[�V��V�#����}c፨e�ǜ�G�S�\�1m�=
'���]㪟WzOvE�T��TS%�B�Aד�=�*��:��$L.nH[)��2�?6As���6�TT�y
3$o�xջ}W���/��L��v`�y���z3c����;5�]�/�����K'�N�2=����rk���ۢ��믮��@}]w�y��9�eϪ��̘�:��#;ʧ*6b�\��3�0�&�1,>ӹ���,����"N�����j�/�7���Y.�<�P�	�K����\������zy��7rd��=z��A�8 �V�d�|;{����fT.��v� ��xBmW`�=���2�|~��7���&�/�VM�;v@�˜
����ʺ���\�+���z�f����ڿ>�	��汜}��%��A��A�:�wy�ܲ�LW}b��C�Ev�X+���ũ?j������C�ָ鍮z��^���S�e2�ה�]�i���wE��̕��3�9����l�AO�o
�$����_&D+m����%���&��%ޯ�:O�u	�*-����:���5�8����Y�גs�Z�H�{��# ��Js�f����W��_�^�QTϪvTP��p�@�"Z��.���m٠)!w���SM{���.��2fY7
�mW �ۈ���E�_}���g���261���!< �0�<�ͺ�v]�*~~k�y{��"���[l~�s���l5�TE�3e�)s��&bu�GJ�/�J�@�=10iϣ])�n�c����.��	�e;�^GL��B�O��f�I5x�<,kGx\^�	Q0����ѓ���7�n�2�L�E<�3��@F��#��y�MS����LD�A}�.�C[�lr�L-㓲m��	@H�U���iw9����%p�*"�~}�!$C*��e;���y
��u�|�Ʉ�z8{��%�l�޺���o�)^T
���L��Y^���:���O��L�Ltj���ߨ��gop�섦\vHt�t���d˘��˂��YU���U3�s��E�cgu�YN�������o��fL���̙h묺�� 0������R����*�v���sȸ5��>���2D��e]��WOd��L����{p/!��&/��Ln+s�
[�"�2����	��z�v��r5��n9���>�r��j�!�
�Ԁ&l���5i���&�(�"oz���}����Orx�jp��+��=�2�F�)2�ɯ	���LLl�����'�8.�2�A�r'����֮HLg٣f���-��'��o.1�+.�>M����77��/�N�0�s�2ώ _����/��J������}g�O�sb�̂8�W{�m�tƱ�3�2���� ����\����߻jyZ�a>r_?d���nE/OKߺnS�g��Y��`��{f92gf���1נ׏<�H�Qː��亐Otn�c��}��5�d��@��rg�#cߓ�M�}t�M�![԰����C�9ӗ{܆��R\>?9�ĉ&�wv�;a��*֘7/�5��*�3��w}�0�m�([p�81���]�{xz�zԡ>�{lq��pb�h�_��Z�~�:/	n�f�]3q[�$��_ R�R���A���I�l���Sg�pD���\|�g(�c)�.�"-�v�2{n�ݠVH�s��-�r�'QV:�K�^Ӽ~#Nh[����;���jǐ[:+ã7�a�b��0 ������r�&���!��gMR����~�ۓ�Srj�ߗh���(����-��]��̷)��p[ҷ�FP��y΃3T+�pV������2��i8�J��M���r�|@	&�p[t�]��iS�Wb�(�,6��%�aѡ+rY�6'o�^�����w�k�E�u���q^�p�<s��+Onp�V<�-淂L��{)AΚ�\�I_v��]�(��:��	+�KsYfj#O�<�d�7�G��Y݅�^u���D��E}��<�/G���<�)�f�y�w
��0T��s<V�]W�N!�q4�<=�~y���
�
/*���ޓ��^�YS���*��ҙ�h'�{Ӑ���$D^��UQ^�S�9�^E�k�'B��jUJ D�$xU�6���W/)���NS���3ݓ��I���A���Y�-�N���V����7����G�@�弾w�������{���u�&[��d9$T)3��yW�HQLs�3WW�fb.�B����_[�t@w�t��ƻ�e���]�:����)�l�s{�K������k�
�;22���L0����S�n�5ɐl�1��Ro�����pK�8ל\h�v�$��m�jy��_����Ag`�{#�a�s�/���s��2cvמ�trdֻ0c�A�gy��m\39ɘZ�Ǘ?;�5���9۲v�L�6��ؑ��!��7(n�颍ݫU��l�y�@���2J۽�]�ȟ��ۧZ�P�z{y\����i��}�X�\И� љ��̗��B�֥�헗���-�U�5l��=���u���Pq��L����f�ֲ�3��[�E�M��=fe��7�'����u��ǰt��AL�tl����}�}��GZ�mqd�S͈�6M��ۓ�nI����fB�.��52����<�6fc�@5S
|MEA�n׌����ǉ:�[Qza�xTMt���[Ք��WZ�U������w��|n�=!�v��=���=���^u��i��S��8}�q�(��9˓@�6Ew�=�;}~uت��{Ғ�4�،ot�k4gvH��u�&���d�Z����}����f�93��)�|~jj-��9�N�fYƽ]<��Y��K�1��I�nS^��j<�u�˪���f��ǆ^�}[f���\=qhk�����=���0-T��#���8�ee[�ll\�q���;�]���u��=������o:�%۬��ۥf�W�P���溕�СPu�/H���C�˥u��~nԂ����+o=Y�ޛ�1�P�N�w3���M�#�qr-���������<���۸/��d3�Ƣ;%z!�
g��O;pw��='V ��H�k�e����x�9�Eۺ՛��|�)!��z��w�9���A��������SI�;��N�,�tg���x�`�lqQ�]���k���ٹ� �=p�՞��\e7Uu�l+���ک�1�NK�sm�e�LNcE��am�7`�u�)ӷ,eA�=c���{�^�oK���笶�Y�!6SW9����BD�n^��'NxR�r�aO�7���2+ղ�������y���-��+%s"s�y~�Q���9:�D�K=�K�A�������VǐC��n2�*�	u\�\��C������m�^ܼ�h#�����VO����%��}K�ܮ��CY[0	!8V��b��T�¥�g3l��˩,f�����o9;,'���K>0�B��O��uȞQ�z����{������5�?0��?��k�����r�7o��sG��2n�bE�^n�O�3��)�7$�B�d��󷞏<��n��[����rd�ɬ�l�в���﮻�g^�
�iv�!�rzEFd[g5�h�=5.BU��Bb�����-��˻��Z�~�;�A�]���*
46EAt��u�.���q�f�I�t���Eux�Ͷ7�{
c%L6�q;���l�z-���TlO��k:(��Q���)v�}.��0�O�O8|��S��
=1R�Q��Crn^�9�J_zk��ꏢ|��_X�571j�ӯ�TF�κ��sۮz�?zMc��+��e;�Tߊ�� n���B��]+��r��b�uA^��
8�WxU��F7ֈ|�/Eɷ繕�����׭�rV��n��NN��B�������̊�r_cJ�=
�O�|��/w
b�:��9'/���v��Q��;��vj���v
qp@����u�;���9P>V�w5��Mi�nB�[�����j=«��^5�n��x�á������ �%�wJ_���
a6���_�ٞ�	7J�ql�K[��$)<�{��9k��R��w�Z_z#�6�����L�P7��歔\*�6͙����덾��P�������<ypcN�>�D�_+WN����v�1��k<��|6۝|�_h�lQ1�[���9���w*{���x��ѵyu]a
�Q�]0{�]����2_��;�p��
k��t��j�oK��r��=$v0e�9�E0���s3ךW*M��$ڟ:e�C��#ѹa׷s���0T9�ى���q���P��~
��D�^��]��2[vª	v�u��[��E����پ�]Eg�/H
i�Y[Di��x�]A5b�u��}L�ꗍ=�}�oJh��G�}�������dÜkΙ�&I}�>=�L��}w1�[=�e�eS)�w��b��U�
���Ӎ�Q�8P�]����^��z��OLqx=���C)��#�W�8��vj��Wo,���������e���0v��.er�8rky�����[YL�+Z��^K�ko�ֺ��.�ŵ�# ��u�^�3��A���G*��BؗN��B��nX�D߹���;p�3J�^��3=^|f73s��A�1�BV�)��׬���֮K�����<����+� �;��8��a߻��h'fC�?Iz���53ە;"��τƮ��R�:���߀$�u~���� ev	���2]xs*}�I�Ǻ���Z��u���T�K3�'dc͜����ǡk8��!�}z�ȫ�������d��y�d�kr���5�qY;�飧����9+���~#=�{���6�.���:��O_ʊr�3I���]��^�)��o^mI-r�uçs��3���g��Ԩ��O�}��xKa�G�>�ѿ��J�xQו�VZ��ּ�,|�Pm`�t�.6�Z�C+#9;�sN��\�߰%���0���.�-�zn�%:6r
�_s;�S������s�$�f�3s���݌>D�.�Xκk,��g}����]�Aܷl
5�ջ]�\gm�^nFg3��w�UG��/F��4i������}��>��[��>b�gC�2���4�wG�눹�� 7�,�b�i��{
@V`�.��>�r3dS�L�p�vI�{�^���<�b�ѳ�1rύ�nM�Si�X������F���AvM��{�{���ɦt�����f�C��١^�����zQ�sS����[��Nra:s0J]����yA��󉉚�P�S�||W���8Gi˱0%�NFZ_5i�}�h�[�z����D9�2�v�x�8�`�YI�t����<�
��D�d�+��O��0��Բ͇�G��q���h'�Z+u��2���Wj�j2&���[k�3wd�h�yA��j�KİP@��WC�|���c���3�X[E����]�c3Wf�%W�>̭"_���+o���g���>8t/f�o���=~��>.�)�s�\Pm��ݚ�y��J�މ[��t`��ڰ��^v�]"��S��&��T	I0W���o_U���W�����W�ʼ�x�VW'a�:�Q�Ojs�X@���0�b'yօi��yV��т����w#�
��܈'f��`�{�!��8��Δ�gG}�@1Ѻʃ*�ݷg�z�{!�dުy�Ձ�}�����>��֟/�����%�x����8[8�<�&q)v3��m&�j�Oln���5]��x{I��]�XLR�eĆ!ܦ�^���ʥ��>Î��� �k�'s5ó(Ĩnt����"�v��ݾ�i
ה{GY�x;�wpZ��!ݳ��r%�_�縞U	9~5�H'e{��P��'��&x'����o\O�Oz���Q���{����C����`P@����g��PY�n۹{<H)h�&�1�%�1Y�u�˝��##��(k����-JK�e9?UU��S=��y��G���`��8IqnNE�}g�҃H�EC��3�/�
��fbH�Yb�{�y��Mn��
�mաA�g[k��q�*�.��6���Anݼp���T�x�yt��_��o	��l&�l;��>�Pg�i�sܣ�SP�f��}��M��.���Ք�87�m�M+�:����׭u�6C̑��w{ގ��<�v%�lS�����#wk� �$��.#�˓>�F}&a���3.�k֯ ҽ$�s`��[E>�p�x�Y��6O�/ϑ�@����F*�Od�]�>��n�� ��dt���Ի��p�Z�Zm���������z�Lk�-��{�����u�B)�ޏ�c<�y���-�n��K��f^p�Fg/�'ܺ�c�k��6�%|}y���:�g�v� �[R��C�mI/��_1�)X��e���=����<Y(�����G����5*�� ���E|�e=t�ϧ���������ef����B��}k�j-��7�.\"��wu�(Y��9]�2��"��sީu֫cb�-� �/����[�w����ٹȸT3"
��!�땭[��+���ۢq w���o2�\Y@��4�O����s��|��O�j���}�sϲc|���r�,Q:��?_W��|7�	���|yP��4˨��YW�4��$��(Q�P\�;�z��W�]ru�ʪ�>|f�Ks� �-�Ʋ��Up\��[������'9:�Pd��Ǚ>��\&^�c��p�j��=r��aWa��]�8�&��^\�o�{��d��z%��K�}W�{�q붼3��l�S�מ���|��qrb���I�J-�>=r�蹷U��N��^S�P����A[�Z� ��r�'yF�G���:�!�oޅ�IL"���u�9�e��F�z��j�3i
��!�����u�'��}�۳(QܡkaɇQx��;����oĒI�+����ȑ�$���1��T��.�0���1��3\�9�+�왐K^�)��ﶷ{ׅ�=k����~?���8�g���ߓ���+{��0c-�)�q ƻD)�z6�w6�mڵu���)��N����`b[�zm��V,õ��7��ꍃOh�и�����J����7�W/9.�q�0���W\�o������𨁺�	n��ڼ~��J,�5������I��=�x�O��>�z2[���V�\��M@�;u䟕_}���-�i����b��G	�Ǡ�{��=|o��k'����b6�3�ؽ���%���c��\9�[oG1uՂr�w�ڶ�?j�C�y�T��,Ə�ᝑǉ͍�Z�vygi�f'�\�kf�٭C�v�� ��������Y�(�������T'P�;}�j�5�w1l��nR��K�1����dS��ܛoB��Q�;�H�^�J���	��z#*�-�/������2�����7`N
��|����e���FƮp�������S�$����ޠN.�X9in�����Y��c���_t\�n:��z^r]Z�\Β�8�Q*�;����M�˜�+�\�%���}�n_����>E��}{]�.���?�l�,d�cτ�J�dJ�sӐ�g�9M�,���x��͊�)�9��uN�����q8wv==�jr#�S�k�Q�0q/�<;�7�P��'ד[X�1��/��Z�To��3X�I�Y��7�2>�<��ɩ{z;
0��aC�T�z0q��'��j�}���J��*���M�VD�P}m6��p��Y�A�#��5����o�!�:u�\�ä`Ǻ5�|w�j�莭�5�mÝn�6���9��j�S(CGYB�}������Hgy�yR��PWP1#fb��P�v%�\����ċ˒ƅŷ/^��z��>7�ݰlH콮�[�_�w������Y���*S�w�پ���~*D��!�l~���3_I�8�w�I�zMuk���~mV����sQ}��sK���Qcp�� ���<"x�;FV5+�h�%!����uPMda�7�|�%9|�����)��
Uc6�˃ˌK�ǃJ?[�;o};/iO�I���*Q���=]-4�˶D��r��'P��B��90�L�˗m�؛�����X�t+Jݲc����$�ͮ�1���c�6�]Ϙ��#���u�p�n"�%�׵�mc�TF�7Gc�z`t��-�#����פH�t�vx��~��K����ԛ1Y���}9۹b�����z��/-��8�����b��د2jq�.����T	tcE��[����>�V�{+��w���KA����^s�k���9Qe�%�-�''98����`�ؚ�\+�!�\�((�{}\m�0n{���\b������듸ڸؼ��	j��ƛ�#�dv�hjҙ���.��ta�D� �D$�m�����ڭ�Gƕg�eD�}��Κ|פ�%�k|�C�u����T�<�(�
��U���M1�XO ]W!�0M�e�j�c�|��V����z��'���_�������~��'>��+Z���<}�u �{�Yn��9z��Ӭ�/-5�{7�ur�}�67�:�֫L��\:s�y���w��y��J|7z�7���}�Z"��X��4�ƚ�n������x.��c9]XMգ����e����3��Y;J��� ���*v%��۫
w'xG��Ƀ#1���7lC&��}�/�m�w�VM����r���H�K�P֗ctt��4��@h2�s�� $���V�75c>RW�z�.�����Ö1^�VeY�TT� J(໵G�)TI0���}&��y���/*r�Յ�����K4�����\�Wu�	8��߃\�Ro-5�:�]�Y5o�n�,���P�[�d�eV=�˙p�5�u*J+5�;� �]V�n�y�OZe��m	{Yh�������W�ohbf7���o$�nX�j$��"���=�^@ �s�u]���R۫!��'%��Kޣ#�J�ճ\z�-�*�m	88N�k��WEHr�#ږL�,ݭ�/���r4����k#��ףm�O���������t�)�:�2&x�I<�Ƭ���Ǟ���2I�^��d:I��=�(�Y�L������{�r���d	2(O"O)�%F�x̆j�N2Y<!ÒB2Sr2ܶ�Y̝�u���R�4k�Zgr��[�I�U�����ؕA�w����ǷpcE�I�>��My){���>��1��Fꕫd�8'/]��R�r��;���A	>�ٯT�ݴ�O9}Q��܅>�XW��i]�ϟ�������&e�N�S��w��_#Z=�M���^�=MO�
|�����i��mlO�k�T�|V��������+��<ve@���G_�'�V'���N]8{�<�m���HxP��N]��iI�7ʳ�}U�L�[-*N�J��sXЬUk��o�p��j�\�*�'�	��\j[c*snM�K�s�TŞƝ��� �6�B���BF�ψ�i��}=��J}�{Jk��������ߦrm��7qx�`o<�KgAڳy��#U+�2�y�<�����|_;��^�__��{[ˍ޹�/@-��
М{`�殩���(=ǳ�t	ai��n���%���r8!ԗ��z)Zb��G�"?-�`e�'�W����`	
��N����2%���T�/�4���f�f�B7����x����c��o+'kZ����43���ׂ��}J�_�0ʄ�D[�����'��h=�yU�H޹�G^���_'�c��]�Nnq����;r�C�l�嫳k���n�P��K�'Xy�Q��^؍�خ��,dȪ9}ު��e��fy�zB��6ӗ�h�ԕc�򊍕*�sz=�\2??�fgc�w�W}7=j�ػ�4�ֻ׃i���4���V�eb�q
&�K5g忟��%�"ɏ�9�/SC5�E�O��l� �;9c�N�Et`���V�6C�Ľ%%=#c�v��0��D=���|�:3xN��7!#5zˊ1�W1?(�u�}7>�H�e�|���W+z�ʻ�{��xCn��b�9[n+ov�Tʒ�ZL�",���Ԭ֤��k;ɟ�[����{��7�k���z�}%����oE��EP��������|�C~)�ڼT��7�|��|���H�>O�+� (���4߹�C�'/a�����I��w���Ko�>?Ek��*����fFۖؕ{����~{�����f-�/rv�HG��_�O��{;F<11�p	���`~�O�4����3�6�|������*RˋV^(�z����E�6�t\�����0�ajvY-\��p����6<��>cv>.)�x���2�o�����m,�1�{I���nՠ����Z&^"Ѓ*&	��٧_���
�����-������r�,����o�=/���6�N��ɳ����O:��������v�k����u?��N7=��w�;o�0c�����S��-vo�Ot�>�����l͜�j��r����}3p��KN]��8��:r�K�3�Lm�=��m�q��Ұ���W\tІ_V�N��<O��6�~�kg��C�y��d%Z�������0g(�$�J*R(黤�/{���J��qL)mv��8Y���}@Q%h~~���g6p�`���\Dg���&��*��1�j��6���������y��ԩ�Z��(殥��A��sk��{n�h.�Aҗ{�6@����lU���&�����6N��ܢ�K�n^�r��} �1��d��o{���Wj�	�Htm���̫�M�N�Ǝ����[�e�-�c2��xvo�q�6��থb��8��kGN���O1y�[���T<�a֬��]�r�ioѸ���t��� �U<�/��{^1�u|�*���Lče�%7�,����qX��\H�m���*�1N�y(F���X��;�r�TL�&�גEOQ�|6f:����5W��R�|��x��6�����U����{����� 󍎮u���m��}|����v_J_��Ƨ9f�ZӶx�4�Vy�E�%o3�S�Mi��f���\d�%�n��mɷ`�8gw4�� ��S�0h3l���|Ӎ���y�Ra�1���>��n��\��?���=O��V;ڏ��-=�񾣽$Z]k��6����_L��%�g�x��w�������K���ǡiXu��S��y�+���o(�S��Hv����T���@;�¡ϫ��a����q�'���tY��q�D��y���ծ�vA��t�n���U��)�]ԛҵ��:�>Md��Ǩl\�mZn5���'�e�&�"V^�!�V�q*c~�H3�z��xtҏ+���e�]�d�<�}}⯡���Օ{Id�9w��j[�%�3�`����Z�瘥m�8���r�G����vg�=�|�W�-o���7	�&}�e�&ְ�<�#��9���g�z����SТjd���/�=�ol����ɵr�h�/�o�v �w����!��{�H��<������aI�x��z��_lŤ�E����+��;�5y\��1²�"�6��6�䲐�J:q-�#4�b�_Q���f����*dY6(�jbf��1R�Gz����.4����i�j��nm7V��I��S\��m�Qv�X��O��~�}r���p�7�qO��~�WR����
�={����g�w�Y�t[{��۽�zM���6��+\ڜA�2@�����~5���i��}��,s޺R����(E�q��5����)٭��c�ַ-G�i���<�é�R�Ho{���(U�����p�x> ���;w�)��%�?k���$hu�c�	�Ν+�q�%���쩸1�x�w\����&m��v�>����1uk(��4�j�©[�"�`bK[�]������RE3R��G�^+�tl74�A�t&|�0�B��H�B#tޏoeR
d�Y��N�[�]LI[y��9��z�0�D�l.�mgϷG�(������N���MJ"����h}t�;nݝ�k����5��B��3��왛��68s[9��C6R���l��b0� x����[�_��VW0�"�y'�K}P?S�g��H�xN�GsK��t1��k�Kmk��+�ׇg���`d�x�r���p{��Z|����C���=8��# ��Yg�꫾�,�y�O(`�|���ꠉ����]]�}�?i�ŷ}x�(�xa!u��g1�U�Ϝ{�R^�*��o�~�>k��-ȏ=�t���潺Z�[�����}G�C^ߩ���,��r4ܬ�n:c��z�D���K��=��S(0����#�����x��{>{��7�3�p|4�B/���C}F�+\������WF>1�ׁ��O ��	VWO��I$oE������15�U͊^��^e��]�3l9��`=4i��|��W#�z���*�o@u9=ݲ��w�W�_y��r`l8+go+�w�pkI�6�TңY���f�֨T�-hu�����}�'d�R���RI&D�sň����ۮ�k�BӅ�A�'1��Տx�ɀ/hag����*�%��s�s��.�Kk����疕�r����O���n��F��B<��|>���o3��r3ܹ�Lzu�
�(>W+}�ȳ��qz���馔�އ"�t�������	]5�*tp�=�|)	�0 ��v$*�]ε�d�%�C3ӇsS��獞���57�C���&XH����s�$����H�Z�"p�_A��� �lc�<�V��8'^Ɲ��͓<�.z�<�k�z�'+;Cn��)(���f�t���"�0�,�z.�E�{˶tF����n�����.��W��ۊtNh &!�Ǧ���~���"��w9��L��#'ҩ_�x��uG#6)�S+����J��xv��%���ZT���Y#t[�T��)K�5:�'$C�Xk���v���F�wW�sb����RU�x�	7��ԑ�u����m/>w]T'Z&j�.Fq��wq��te��f��p�(0�wQPN^�]A
��ajs�=�A���{ٵcg�����ރc��,��/>X��	����q������+��Qg���-�Y%Ħouq�z�X4*�ջqV糦�,e���^�B8}czᠴ� "n��7eM�xa��J̄�|5r\��*N�����liVلH�4t[��d�&�U�˟!n�t��O\�Y��c��.!�eE�bUg\��^hӍ�'S.�������q�N{��_'<G`�P����˱�D�~\fLl❲�N��
�k��>�^B���퇮0O/�|��QT�WZ⢉[�x5�s}��{�C`"�>�R��[�C��sϵ�mX�Zʦm�Nq�D�.g�Yj.�̒ ,�ydG�r�[r�6I�nvc�����9��U<�ݗ�q/!�W��ԙbs����b=������5���|���o�
��k����kY^��g�F�,�m��s�Y��/�Z�W�I�����%�ږ��*Z/�P�4�B}}��t��F+��sB�m����	;�v	�[�o�K�������*�q�Q���Oh�{1�����w��Κ�)SI�Kb�
��m�ͼ&�Mk�k%[OS��Y9�Z���H�.N.w\R�$y���7�嵺E����Tc�ȝ�;��4�UE�1q���ާ�w�����ߓ�ϑ\����R��A]1����޳q��b����A�
P���캫�|����O��>����V��%T�a�+����`�=b��ᨹ�]�k��q_z{�������*�E��v�.�<\C#6����LM���,۰;�K�K�֓2�\��.1kWfwq��V�%9`S���q�ߨ��ς�����c@��h���M��c. 5�i��U'H�sv`C(�O��an$\���ا�I�����9 �R��<fp0�~�x�@ɵѵF;�Z�\[L��xͮ��uI�h�V�d�$���	]�$_�N�4��뻝V׌�k�w���1�s9�Y,��{�3����{�'N�f)=Iɧz���7V�Ӕ�XY�h�e����V�rY�92s����a�����7�dz�r���]�cf�b�G�=��R�>�i��壮�^�iRZ�����MϱO�m��ɠ����ܖ3��sr�u�Z�@�՞��nۖ]�s�u���u�{��x1cڞ��]���'��Xt�u���cB����IS��u��,�oz�\I�b'�R�>!�P����h
�d,>n#��A�w<1����3��e�y�by-�8d'�I��%����|ל�W��|Y���ř��^4����/��!�K��Wt���e%��u4�$�ќwV>2V��4�m�ʷ�VkR��%=�-�ؐ��;(��]��]Q�x�A� ]e#��YK�G�qéXw�����u�����3$ql�R����\�\:�èQ���|�̼Q��ݝ4�t�����}r��v�cS��(�l
���m��(��
�@ݣ�C�JPb߭�����&W�ri�\�����կ��[W�9����j�Wq�r�X{n9��gS7��=fkj���t,�u
�2(Y�ջ����Ok}�P�6��.G͵-��W3��Tz���9����M%L�z��P�m��d+�e��E�U��Aj��m��+<�ђ�of�i�Uq���/7$��{=�i�sé�)+E��}�ڠ�WBq��6��X�&r�ϗiq��g�'� x:��_GG�yePwq�r�/rO3��`=ݼ�(���<^�V]� ��wD>˜����;ȿ�6w�?g�k5��rn|s�$�A]���"��r7q.F�Dpٌ�8pj�5{�<���&��sh��-sW����TU'��m&��ڭ�om��V3�Mgk��J��S�ahd3�B���^Y=m9)�vݭ�h�YqQ�aa*ZOk^W;���
��6��!)�nL��Rq��2� 4
�,
�`�Xؽ~�o�R��vNoG��Y%��ԣ����Vn2U]o����br&'ԅ=��P�A�z�ohSO�<�gl�f�X�)<�m�VH;*���� �(�YG;iRdm�bg�0�\�x:���˦�3=��s�d��֭�4���sCKq����XFfƶ����]��}_�kՏ~�n�7�CW_�����[�D��a�	��q�g_gC)O5�۱�V.���>巄u�7�����c�s�vvN��e�ӗp�ԣ��������k�G]�h�{�ƖέR�5`���}�~�j":�
��M��k�Uy�|V������4&߲��Χ�4��W�Y�s��l]sʦ�l���hơ1qV1�0&�}f(��-Nɼ�N�i�ʛ{o/�3���э��pk^��ũ�燦�	.)���Ռf�)�j���ݗ�[���n�Y��>�֯y�q��p��0qh��SmF�/R�*r*�'7ޮ���,kꑥ��!�w�Sњg��{����,إ{��P�����l�.�k�Ȗ�˛[��}I�������x7�]������c�7�,�~���}���R�ӑϫy��N�Gn��=vI��y0�=8�io�k�c<��~r�n�׸�w�t8�:�H%��\��\N��AW�H����!��}4�i�_���m�R�hĖ%���E�7;! /tbs�6?z'`�D1ڬ3l�(z=nQ��l�Q�1�Sf��ޞ[&f:��5��GV�fXy���)������"���k37+s�X��C���+���w�E�Fs�}��&��ᰋ�j��Y7}TE?�uv�9���o}���+�O��)x�����2{����f�bx?�п�N���i�*�T&�/F�}���|q�=����=�7]`P�[�n�u%[xƆ����"ӗ`��N�v7�괽�u�sਫ਼���U���>�2��Z1!�ȓ�x�`�pr3��S��V��t�8��H���Qq��(�W��&
��ݠ��率��4���D��"����b��jށ�����E.�2w�����5L>��0�Հ	��n��őL�������}��x��]B��X����F�'q�Y����{����4����4YT��+&E�*�ET�3f�N=�M�&���{�:�c�E�v�����͎��7��yծ����ll��OYX��e^�t5a�p��x��t�S��\6hr���oP�v0p�a���x�%E2�e7^rn���"Y}�7���Mo
����>��I6}s�rs>t�Z ���6�r0��1�;�sSÙnf���C�ne�9�����(ޤ��B=�0�Z����4�/�,���M��G�bq���kҴ���c�泑^k���k}��X�%�ζ���������c�2�=�rXױ�ƽ+][�r|�;��/�q��oW[�`��� ��/��E�+z(lrY�~�����(eQ�oi�y��z0_|#�[�b�ϼF<�}=u���r���G=4�����K�/��G�؆i�Dj���[Vg���6�2B��^%��w*b�kr)-j<��
r9��6��w谝�=¸��\�&Ȟ�|����+)n�[�Ng���A�0�]�]w���j��lx���½.���|�4��QZ���8����]��L�
�I�n(��[�����u75���qMC"r�V��[���u��X��0���+��GX�z��oyurץ�L��y:f��U-���Ü������1~ި��53������.i}�l[�_�1|�ޗ�ּJqY%�t�[�|�!���kQ7e����(�ݼ1���Q�����V&�^��)lz�y1��}άн=��f�Jvr<��j��!��!^L�ś�~g�z���"z�Tm���澋�&21_���7lE�o[z�.���/��,�ʩ��Ơ\�����W��gY3ds>ys���]}�L����WnT�ع�N�b�M�6b������-�V�<`̼�}3.�Ie9v,��r��۴���1B13�naj#��α4E���'�ќ��{�Ɲט����^F��G|#�}��7����^#��6�ٳ�[�=[6S��%&�bq���d�p7��A_$6��i3��[T��ʽ�r�)�[sgx�����s�8�Ѣ�M�=�� fE�H����}���~����e{�U������K���b@�I����j$�G��#���5�����!2vT�} �q�?�>Ç�૧<3�5���M�HH0 �*iBD�! �?ϓѮ�&��6�B@B�L�Hh�a�Ms����	G��'��Z$�G����`����~�����}�!a�4?�+�QA�pa+��x@a��2��J���@���qi_܈�!�Ƞ����BI$�#��~_BO�Kc��&%`�BI#���hBI$������	I��������������Z �?���%��e���>��N����$�0?�#����~��c��I�4�E�����Z�Pw���(C��AD�"?��"#�ԓ
�~��a���`����~R��Ω��!��4B$�C0�(���[1%2_�s�� I$�#�?��q$�6؃z(R@P}-��	
���pG�u���p��HI#�R:4�iA����
���9���� E"%�?�~�Z*�?���_T��/�� �
?�~g��A���	w�������� BI$W�(I�����:~����4g��Ӂ�Y�~�$^A	���G��3����Mо����ـ`}B~�/�w�������ϴ���$�>�?�������L ���B��F3�@�=����5�ϪH 0d���H��x���G��_������1@}8%���"#�P���(BI$��@�e�C/*G����0_Tݠ@ (CJ�J�`1#�? �T?������8b���^�&"R]���1K@�VQ����II$yH~�����G����$��C�	�I0���� ~���O���������������}���H$~�>��� O����?��@�O��kߛG���D)�(�R9�_�����!I$~��_u}������@�����Db�B�H������)?���C���������}���#�����0�R�g���AK�P������4�0�Y��xa�O�~������X��}�}y��� I$��������~rX�]��~������|m��B�{~#��	��>�	�BI$�IE+� �F�H��/���o�?_�!	$�����܆.�����~�B�>�	bh*����3GR>�m1�~�3��??��B��+_���"�(H5�j��