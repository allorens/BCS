BZh91AY&SYN�uM�_�`qg���#� ����bH               =� ��Rm�(JA@$��	
(%E
*�)(  PUJT�R�ED֑�֣L�HP�@$����W�$�T���̤��!*�D%UEITJ��a�B�U()5�UV�*��R���F��/{ P{+��TB�w2�U��� �j��� ۱�EB�p�JJ��4�Z��j�������Il�(�+cI-`T*��� �Q!J0    ��U  � 6�| M�Z0�P�Ӹ��,��M����n������hi�w��4=Rsi ���(R��j��J�+[}�)H ��#�Tm�h��lԕH�ݞ�xJZ��׏;ǳ4�^�wzV�{iT��<����V��-�z�U ���=H�{j��8=*�h��<^9�Q֤�v��HW�����b� _|����^�㻾
�fQ��/:��C���K�z�J����=�IVx��7��j�=�ǽJW��T�����
�m+�͹�l����j@U=�i�
QR���b�l�� w�>�T
�;�מ�J�]�{sͼԯAݥVry�)U%T9�<��J��]�ީS��Vk����V�ڜ����{��z��Q�wnOw@=Z��$�)2�efhR'��I�<��g�UH�z{ފ�()w���RT�K�+��T�*�oj��=j�gxw�*����g��ҩE�oU�w��Wl(�w����Z����ېU(�K�J@���*���R�EL:3�QU)x��T ��O{�UP���]��r�� z^q�  wS����x 4O=jQ( �m��+Y_>�P^�n� �rà�������  �OY� 3'��ޖ� U�׼�����un �ق�P���R��� c�� zy�� u��� Z���}���d�}� ]��랊 Y�� ;��U*�F���Ԋ
}�JI xy�w��g& ��
 gL t�z{��񎂀��z�z�� ;9�� �4���HQP�ER)vQ�Ϣ�$ �����`��Tw  �� ���@��h [�ټ <��  -�� �� �}*�     t    ��d�JQ�      ��1)(��� �4  �jy2
J�F       jxBjj�T�&��14Ѧ���R�U   44   D������ #PѦFA����?3�����BVL���!uw��������=�L{�*;{ՙ�~��N��nw�K���� ����ZS�k�C��@_�?Ї`���C�����'��������?%O������ԒI>�` ����?(��AE��?w�/AL�b[��c��0q��bc��ٌJ`����.1�01��L`cٌJbc���0q�1q��H�C�\bc��&01���11�lbc���01��4��`����0q��bc��11��bc��&01��bc8����%0q��L`c��&8�F&11��L`�8��11�Lq��bc`c6���0q��\bc���11�����&11��bcĶc�8��.01��L`����.01��Lb�8��0)�11�lbc8��2�8��-�1��L`��01��L`�8��.0�q��bc���01�c�L`�8��11��c`c8��01���0q�c��&0alq�L\`c8��01��Lb���IL\`c���&11��c�b�8��.1q��cL1��Kbc0q��`c��4��&1-��L`�8��11ƒ11��L`c���&0bc���1���11��bc��S8��11��L`�#���.01��b�.01��L`����&0�bc���11��c�`c���11���`�8��.01�����&11��`c��0�0q��c�b�`�f0q�lL`c8��0)Ƈ��c���&11��bc#���11��`c�c��01��c�`�bc�8��01��L`�m&0i��`�8��&1q���bc8��0q��`c�c���11��`�c�\b[8��11��
a�\`����0q��m��0q�c0q�c�\bc8�1�c�c�#�C�0a�0\`�@F%�����0q��bc`F&0q��bc���8�0q��`������0q��`�8��&01�b�8��0q��`�#8��0q��i1�LLb����1q��1�L8��11���0q�l`����&0q�l1�L`�8��.0�&11�lLb����a�`��0q��L`�S`��8��0q��L`�1��b�8��.11��Kq��&0q��L`����&bc���0q��c��1�c8��0qƆ1q�c���c�b��1\e1Q� 0�
���4�W�cb#�q�&1A�"8�Sb�Dq�1� ��G��b+�Tq��1ؠc `��Qq�0�����\b��0P� 8���`��Dq��0A� 8�S�c\b��Q�cLb�lq��1�*8�(�`��Q1���0�*��G*cL`��Aq�&1P� ���cLb0�*��R�"cb��E1��0A�8�C� �b�1�&0A�(��S�c`)�E1���LbLU1�&0D����� L`)�Dq�&0T� 8�S�F	�1�&1T� ��S �W��b-1\b��-�1P�1E�*��S�\`10@1�.0����c` cL`�U1�6�`Lq��1E����`c1����&11��Lbc���11�1�L`�8���e�1�L`����11��db�8���`� �1q��1��[`����11��\b�i1��[bc8��.0�8Ŧ&0q���`�8��&0q��bc���&11��LcLq��bc8��1q��`c����&0q��`�c��1q��bc���&0q��q�bc8��.11��L`�8��0�bc8��.01��L`�iq�LL`c���&1q�l�%11��Lb�8���4��11��\bc8��&11��c�`c���0q��`S�1-���`c��>�&Py�������]�^<���u��o^b��(\;u4��%LX��*r�2��2�т
(nVeRyX�и)ݞ�eb�ۦ��\�-�,�R8�b�ts\����-��4Yv��$�f͒3�Z|�ӕE�4��u��V6��m��bV��[��\+{J��I�J� ��MD]�!�#UbiS��;����ˑ�E���4�@\�K�FQ�#�Zj��K
�Qpd��b ���`����Mֻ�zd��ZJ�#�	[9mQ���v�]'a�`�$L(�E��ۈ0c���� ]JG��)���Dr���p����k[CJق��A�����mk��	I�B��Q��a���lu��7rZ��*����l<�L�ܖ2�ER��/cl�K,��s�ۼ��0���-˧t��*��&�MP���]�����.Pe
8L��.�Nkp�T�r�Ա�t��6+\A���ޛK�����*�dӶ��@$�n����w�����4*�Qy��£�R�=�C�K$u���z3<FnS#�i�SLә��L*���6�&�Z�Ql������JP 3#uh��Tݩ�i� :8f[�����e\DF6r0��Z�m��p��W�1����o.ve�2b#-<�������Iˤh��mZ�Z�5͙6�^t���ȱcé&Vu���xa�W�0\�kT�d�u)����YO1h�V��i�P��]M��z&`���uJ���=w���K�,�dw����4S�U10�e6%I4����e�-a�85����ֹ�X.����f\�,�×�YB�r!M����;�������+H�L��mlY)ǯ@Xv�6-���n�Qd�^H*F�V0�Wը��|�;��y�ñY,jJ���E�t�i�<�4$;Vc�U����E7,��p��*t�l^Sԃ�q�A`g��4m�2G�ѫܠX�����u�(�u{͘��!&L>��ւ�׬Ӗ�݇��3������FɼU����)�E,qî��:��.�R'O(ZWj�+4�R^ndXqǛ��s`PUC��#�Sc6�������L�w6K�Z]3�N�w&)����P:����ĵ����m���`�e�K[n�8�e[ɻwN��5vF�TQG`���űn���l[�Kq՘��[�9A���M��2:56���:��'�_�e�+b����ђ��Œ�V�z�:�l,�ڻf�Ю�������L�-Kk&&k/iQV��:�����2�Zu\��,<:nj��yH�L�j@mRˤX�w)z���rm��+z�k�<) 6]*�	>6��6D��3B���d?<B�k�i�w�c5/lͰ��f݀�dT�jao3U͸ܼ�-�G2�(Rѷ3Mj��û(5r� ����ԡ��c$&��l���&�"�l�L���O6��1EPY$+��(�D˷@�AOTD�xVf���i�{��wqY���Ĵ3(��c(�zj݋UtF[b+��q��zKD=�Vʋ�]�+N�Uy0-s,�[�-�k6h��L��7E��QZ�kE�66o(h�hcԞ��Iw-�Đ�)�7�^����Y�բV���d�a��S�16'sGoM�fM��%)jA���J�	�ujn��5-��ﰴ�ݫ�m�.�Yt�Q8ۆȗ0���Z+!r�7&���@ݼ�-����%�p^�Yi(�Q�q�Kƭk���e7W�Jswr��'��R&/��+M!]:����0SS��N�f;���q˄�ێ��~������<��5�M�i��MV��0���P�X�"��0��|6���YQ�+N�z�͊\Ѫov�I0ٲ��3@`����[�7`X0��c4$wW0�{v��P�{GՒT�,򷲞(Sa^ңK�I�ϳ*l�I3߰'nM��N�;w,�""�f`��J���o��D�E��8�D��]5uP*��/�Y�M�R��V�nEyc0U����L+ĄXJ��)Q�+WQ=��w�M@��u�;x�.H0lf wf�p�^-ww%��wo�J�Y/-������6�L˱Ww�0�)^�B������˶��^����Չ��%,��(���T�~/n�AblNVF%ڨ�Kr��	��=���[��"��˫�(�n�E^��S��n�,n�2�K/$R����ҕ���an�0�jXb�V�y.nТxb�wUe��E-z�ҋ�H����#��=8�
".Q	e���&Х�T�2�9z�%�LD���J՗��m<v�J��V�	2Z�зY7	bѕ�P6%�%041x%[����Ս�7W���-b�1���#�7Z�t`�� �ʖ���CF9f�[4�I��*[�ѩ�ǔ(�n�6h�݆�P��1�V����N&d��V�TN[��՗q��fQ�#oX�&��K3	Uj���V�2$�z�mf�Y�Jz#�q�Ԧ˴&n��ƅm��Wm%xs5Tc��l���1MR�P���fJC��h�آΕ1��H�b#ףx�l�^��H��T���)������w*+z��t�YS(l�5VZe ���u��t�W$1��& �=��Q�dD���n�0#Oiq�b4�{���m��U�.�Id��x��"Lk(d�+��d*�U�a\umi�VbJ�<`ڨ������9UYR��=��W��MnʆZ�3w/-�z�誵U2��Vٱ�y�y�pj�����S)KRj�ojAo(Q)5ui�έ36�G�r�T��tX7fK*����q�M#���w+s�*1l�A]��S7�bon��]%��ƍ��Ez��ݤ��<b�{K�yv�]�����������1h�F�,t��OsL�I��6Q�[f�+{qF����7R����b�9M��s!�ER�atX�ȫkR���d�h�M�촆f���ױ��̲^�v�Hš�����N�N�[w�smO�����f]��Kr��CZ�}vE�tf��b�K��m��6���$�x�onL��X��wP�G.
�h)�	��ɈN�Ĩ6<H��h-��X��sl'����F/I�2엢ɚ��e(��Һ
��b���g���7�qf�xr�5y"�tN���d�F��Q\�M�oV�	3�v&ò���r��y��ۇsv��yl�w!ڹX/�ڦ[WYJ_���[��sj[��JY{����U�;����7ww�H�a�z�5_�L������D?�U{��,����Y4`�d�ݝ9`R���c�NB�J{��A��ȌR��xkr�5l�oR��
ȱ23��h������,L�$���m�{�\M���SVc�uPV�VSm���F��na��oNuo]�Y}�;a1(��u�Oirm�w�2�]�r�`z�����?J�cwB΃L4��d�Fއn�lۨmk`��� ��xUi��� �N�ݸ��tT�{p�ri;p���ˣ�M�"�vQL�ɂٹ���,C&ӿ^���J�D҃���z�CE��n�˛���2�@��$ю���Ywəzv�Q8�����6��qB7L~`��%R��ǭV�G/,�Yl��wN�
�?lJ����h
k]�L�Zm'oe�� �@����	m��ژ4�O7c��^L�A#��n˹����*�������ˣB�������u�
3J�Eh�	Uw2�TR�[�` $;K,?]^�A����5WJ�W���d{Q
0#NԆm�WX���)P��uPV���r��B�&�-��hD��J�L�n�K35�Wm9n�X��k�V������zNR̖ m�S��ʽ�`��̈GE��ɩ+hG���9&(�R®j��9N�ٞF��:q�[/-���ݽ�L��	�X�n����5m WgiR7�Z�p�ٶE�
�)
�ͥn�ȵ��,��Xn�A��QN�m�0��t�,���K4QD��`r�.��uu�Ve�7�Up����bͻ�mLJ��m2.G*����6ũ���"��x�)J�f^�����{��0�Uh�&��uQ�1j+�D���ֶ4`�Q��Yo-Z"�"���LM�5�"v����՘�����Vg^Hr��R���c��wxX�0K�,\p+%.�]�e�5n�-����b��ܿ52M�P�NAPE�un�&��o#�6c��sY��&����V� ������3
!56ZF��ڔn�[�ѡMV��Sr�$Fl����䕪�=J�D�^��\��E�.�Xc�t�; �qZ$�udn�-%/r��R
G��l�B���0��&^Y� �Zv��XR�$���x�Y�kD ��7�v�j�������BZ�,=�
���M�͑���ɺ�S�<$$�U�"��MG�Z[R.řU��KJ��n�W��1amX�+��dBe���^�)�O%e<�b�kW�-S��c���� h���)�se���Y���T�E�-9YV&��	WHJe�����bR�s!�g��"�no����L��yc[���WUӸ��q�Cg
��gsE
�^D��.P*�Sn�ٻE,ciZ��bU$x7P��kU�8剉�w��jv1[R�����U��(�l�̽,5��tk˞f�n0E7��Q��AJҮJ���l6H�C�:�^���v�9��l�1�u�t6�+�6�S���
�ّۗae�Y�To1ˠL��e�@�v˭1�T峩�-�@�auCp�'�x�UT-�e�Y�a�s�S��a��lf�x%7N�U�t��t�D��{syW���w�ʍ�C��L��)4�Z�*��D�&�-��MR����VZ��{�u��۶��Q�j�d��#&�Zث7��Rvi�r�r��e]Rt�x��f�b��j�8�SY��D������&D�E4Cᤞ�.7w�ӓY�%f传�T�S4K�wL^�ʄI�h�Ҋ���
Yh�v��i�O$���V6,�f��2L4t�+���iabAyYd�ܑC�r@4�UجԞ��&��Z�全�eӦ�i�L�9J��J���2�v��<]fVX�((*��,1v�驲�p��[�Q,d!x��Iyzj�PW/nk�ݭ�r�L�
Q�49�٧{�¤�L��2��7MV��F�R�歬L�v/v1�*����Yy�;�j���
���v�cR��j�4%��;�+q�ʩv���//Iy1Q�u.�^�v1��IV�r7hDi<�a���c�/vX-xۼ��T(�^R��j���x�`�9�Q�l=7�.�[�HL�a>��D^nf� U�\��H�׹�=�x�U�/H�ر��'
.TɅ�� ����{�U*ƪ�V������)PI�	n�S	��yR�n��ɬ�,9.�$�H����]�R�cb���5)P�V��wr5���:�f�\�.�d��mw����p�[�*�D'rb�c�Cl;O:1<S�����PvjM�71���<�h�q\:k�*�ݝ'�kF2*�pB�9�3l�Vd�0�9�vJ�p�;�x�Z8��P�=��q�Di��S�hC	�KXŘ�#K8��k1`3��I�K�l�č�zxV��DoL��GQ���Y��a��ofC�fV��<�3m�R��YxxQd�zv�#0�T8�6 c���[�n��t����qu��[�m��&+�K�`��U�!0���lR��Q��ռ�B�b3��al뙺!�<�;��	��?(�W�t�C�Euww#���1���sg�3�K&���2��m�e4Xx�ъg���XB�(�=��J��h^�3Z{�T��Q0�n�ϑ�p���G0�d:�D"�cQW�C�N�-6w	��ma�+�U��b1�X,�u�v̆E��zO&�,�fq�Z7���7����q.	�i�=�q߈f��S�T"#�#4�<L�I8C8�����6-ټ#N#xL'K�(U�"z��4✮҉%�D8��1W.��@�O5\�>ԭ6�.�֤I�i�@�G<YD��h�^�&��E��f��;	g�Ⱎ(��(4�.J�Ί����\�Z�D3�>�m�s^[9�)M�"`��)�)�uZD�Wʚz��ț�U��`�Uʡ����M�$ye�R%�{��|��7:��*���Da�+5�V~�#��VAJR`纪Z4�jRQ`;��Z�d.Zm>M-�ZJ$ѣ�����\Q;��x�F��7ĲI.��o:^�km�%I�z�-r���n�ZKRJ�V�sؚ\�E�������%"q6�&���M�u�һFg�VE�=p���Bw�\E#�s�fD��:�Ӝw�it,���r��Z��R֝��ir������Jb�V���L�˒M$�$�I�����[�1�ի��Q*��SM,k&m3�Yal'��}�+$7���e	�,�R;������R#�8�$�x�d�Z�ٻ'�e��뾋�7���K;BP�\ш�ڙ$�U7p��(�D�8�"���CФ�ə@B���H�0����7@q�r�t"���4�=��dCL#���%�K;��Ե�Ֆ�R%!Q�U(��Q*G�ɚG�᳋��.�w!,��aL�2��ࠈ�|f?cޠ����Ã�bZ�-|��LR*��]��4�H�;��iY	����z\��j��<֎�U�ET�'�Ա_,��Ԓ�D�i��ZB��yK풁w���}g!�7�wy1ڦ���8�d,k���M���4�V���U�����Z�l��_H�D�i�Ӂ�,�dY�)*��5W'IR�rT�Z�����]j�����è�ѯf)T��Z�5"N�9�:i���W)���SR��,S���0�ⰾ(��0�+Oat,���8�Sw0�g1��fb&�D�:��՛���	�p�L��D�.M`�V��v���h;ʹ-R%�"��6�[-=2��<���[�P�u�ޭ�?�d~=�'����@?C���;�xK0���Y�~����N�nF�ں#�q'�˗���w��BC�x��&h}A�,�B�gm��������inc)�k1���fv�|e e�G-20�
z�Z�Cn�'+��X�q��ɴ�WZ�y҃��=�XX����"��p�#���2�F����`�r�Y�XP)�V���anfm­�\"W�wKT%%�*�0/*����@���;��}ϙبͣ��^D��vEzX[�בv�a`�oT�d������<t��lȃ|�]�.�77�F_:=*⠖��+,+۬�X鳓�EU�vk�gY{3]^8�ݶ�:�9n�Yk6��ԡ[�.j�.V��88��.�tX�m�U��x�Sw�\E�B��I\�y����a}�����H���o�:k� 2�*��s�f&Ƚl�^*��FN��<5��!+E���,>B����h��eϺ����yv��X-����75Ⱥ1Tl�5}��r<�,�K�gXΒ�>����ƅCce�"��G�<��˛ܺ>��l���໰:�O�"gv���Y%�{�[��C��!n��v��:�٩,��,t���ChWi�ڙe��}Ci.��!��VoS�!K7x)s�{J��*f,�e����:���i�� ��/J��Zk�#9d�W*�H�ZW�[��>F��UJ>�)�xR�ڹ}gT����6t7���i�Uٺ�"K�u9ኚ��	a!����0n���7k�6�w�W�H��֞�h�&Vh�W�a���f�jU6�:pIR�:����/��&��Z�6%�o�WLQ9BX*a2����z�������f�,�����s�B�RCxܙ�<���%��	�������;�:�oi/�Q�1I��p���(eo"	�������ś	G0b�ƭ�[��ށ�湁�}�V���E�L�x޼��ϸ*_0n���7[���q±t��6Lp+�J;��5��$
�/t�:��T��`��2镋����ʛ-d[���N��'(�]��z	lfS�̓�uT�Tͤe��/�L�:��=c��	��s}�#�Iyl���IF��Ӂ��^�\�ۻ����.��esR^�n�h�s`���}��rՊڷVu.�}���Ӡ����"k�vx��+�2#�$bR��G�c|GL�ڪ��2�e�+��q�:�dB��9�]�Ǎ��Ηt2��]j��92�8�G��]��d���Dk���Rխ�C8���t�縛Z�4\��/q�[7gt��g#����S�@��ˆw*7��Ҥ�IG$y;d�u�1mP��b�,�|��e�����¬vf=�5ە�}�wD��@��{F`���
�Cd�`�Q����Gq�"���=;ʇN�VzRűses������S��c;+s4U�kBQ����˖��BwR�}W�>��´7��� KiA�#{V�b%��O>d|.[Y;`WXY����-��GaG��fH��P�~G �����a�y��3WzE�qU�iu�v��k�r�M�+v�:�왲�Ѡ�6C}Jq���!�@�������J�VՔ�+�z�%
.���&|��[��x)b����4�r/<�'Tkb"��KGc���櫨�8�����E���9O�sOs�ɰ�(�S/3�/�Y9�����!�;�P]��ʽ��U)M�3sD(i���JT�hgS����ӓ���i�NѬ�j�l�YP�ȫQ[��v�;K��p�T�,N������=2.�td��eKA})�z����ʃ��GS�{ss�<T:ˍ>+�M�(w7��m�b�n�KrN&��ǙYsg�<��%�b�Eؾ=K#�9^�bz�Л���j%Y��W��`/�i������%q�f�-'6y[2p��c��zq�Q�<�Crw�4keQ�2�StN�ɰҵ�w�\ɥ���SP��=�>4��{o_��x���#�[d�3F�����Խ���Z��L���L�N�G�֝�	���}D����ـ��A/L���A,�v/z�ځ����R�I�!�2N�B�w��W_:�6��ۗ[s ��ӯ#/�<��7u{y��;����q��z��s٣#�O�V�w������:9w�XmW6krs�ӄ�{��˾{Zl��fG�:�s+%*�`��D�����:�Y�@k�L
�Ø%�33��m��h�ӱ���(ұ%m�:Z���z�J�J{,j��}��r����X�fS9t�31�A�f�SQ���ML̐uc�X�:M��ҪX�*������6���w�j^��z�vd4��f��+C�����,Z�������zr|���!��p4�J��v�̍�3��w!��o�<̾g�h��ۆ��*^�����Y�eH����Jj+����˺��)ի(qc�5t*+��l1��	Y.���舽+����Qi�ܴ�مf=xUWE(&�m���}x%Eh9Ձ�qʇ�.͂j�P̉�Q�λ�B�����z�4:Qz,���ƌ1dn�#��zʏ���W2�}��P!�&�Jǀ:wKV�Y&�� ���E��`�k(���&s��\�P��K��l�%姳+6���\I�⤥�7�α;(�rx�cB勊��2��kk&Ὓ���h��	����:��眃�-���Wz���	*���˹V�\V;�κ�iκ�ÔX&�'�p_-�z�(s���Ƿr砂��Un*t�P&���4vg\����KM��9�{���+R�|uf�}cT�F��W�z��7���=�Wt%�&�����',N[�'Wx#����������T��=�t\�W۹O�sJ!��"y-̏p�ۂ��Us,T�_6c�'ha�A`��+�2Io��gPE�1Y�T:������'�����=��8fɥ���<n�	A�K���m6�3u�:�LU���+O}�	<'p�
�j�b����]܍��Lt�1��W�z��m[��S���[���-��8ɮ�#N-���IckU=+$��j�O:c�mX{���q8��8��w��
ӛ[���ڷ����K�DB�y;�ݺxZ���9������+*��%�J�#vo�(�А�ke�.;
!IN��iֻ���./2�R�fR�ܬ�l��[��G/*�z���]�Z�}����RJ�;�22���7z�6���k�Ө��#�tfуzZ�c:���J
�C�����{ŕ5��z��ŏg>��n^ج}�{��3^c7ƨ�a}j���s�h��R;�%���Ԃ�z����w+���O�3�n��I��	R���R���*"���F*�Pѵt(�2��s��c��:��Rs�Y3��F���b�b]X�Um���p��=�!"��;���B������B�F���6����,x�Qkq:�W8�'�*ۤ���=+r'�!�S�a��"0��R˾k�V�8&��X�,!�[��W-}&�7]�䦈�׳�gs��!E)&�ɭW`j�Z.�d�є���#Bݾ���mUW`Ա:͓������D^h�03RʲFp����� �;ԻoP);�]��rl������D'�}�[��#��)m�*�4L�d,ӺͰ;3XhC�]��Bͥ�:����Pu!�yї.{�s�ޡ]KRܹW�Y}X� n�nۧ�!��C1_-��./U��Rz���C!�����K�";M֏; ����	�5&��H�W�W"QΓ#���N���aV-��fD{�M��'��WY�.hQQF�ޗ�6g*|����Wv-�:�oe0q��b�31à��zh7�^]]��x] E����JqX\�녍Es'V���9\9мz�U'KW-��h���$`;v3[����A��6�S݇2�\�a6�'9ʹ�mK�P������4�WC�5'����'n����h�%���J�[�V��ni���:���P�ؔS�[{P�]l7H�㨦���<�����y���˜�K�_Z����9r��C��'�-�6�+i��p��5�x��Ƨ=�C%ج��+��܁q��Ӽ72L���ujp㐣Y�멊�TP�pS#x��:�e��[iW�������p�XkN�]�K5��OU��7{�;���$S��z�TKe��̊�v�5:.�yB�����2-��W����+^�6��K�t��.�u�|�.�"�4�l@��i\1��gE��{���C%�Wo�JR���ވx���ѓ*.�xo(K�� �s
��q�Xп�|�}g���˾jT�`�W�D����������X{��+���Țљ�JN7���Lʍ��0S3�7L�u�H�̭�r��2�:��.!]� �D����m�OD�Xs�XW*�����P��ݭ/H�F[�Toj��F
�� �i�XO�A��N�Inˮ5�}U�o.U�Vd�V��ű+r��wr��vl�ʒݝH��A����j��b �|oa���f%�1t�]R}aԦ!Kgi�;�}�M �� �[�o�BlM���cp���v����p^P�Yw\Bq��׊Pטdq��f��e�KK1����x�W49��®��_u�Yw��Vح�3�\w��_��q]������t�UJ;�W)gv:n��&fe$�>E�Ʋ�#�c^�>7�ܤ6T�3���5̽W�U>;jUIYwk��m�[ݛ�٦l�/I8v*�!���RT�M^���mQ��1�س�>J�)��4n�,t<:��K����_#[u�=���Fu��!0
�	�4��g;�J�n��zd&g[IR��k�h[���t��կGS*��]�eg����M��𔦞��W�q���ya��u�1mfn6N��q�=�	��:-��F(�pΣ�N�]}�e�T�S/x+���l^˼��d�\Y}�@�;
gV�u��&ž�WW	�Jkv�*r�LL�)����3�����N�9]W��1��ݖ�V���<R��v�7U�'P���dˬ2�ӬA��μ���F�_qIآ��k:�ű�j�!>j\��u�c�q�L��Pnęq�x���}��D5��Z���\<z�Y��	��H��Ǻ�j�J���~n1�.�����mՊ���T�yf�{�k��Jޥ3�vL��G2ej�4�����P��v�q��k�'f����30.������P+��N��Ȟ�cw[�.`ޱn��u��g^ofvZ�8�H�/b�z����K�d]9^�lPθD����|d㜸���cVfy��7kq:�����XΩ�-.�ԴV���C+�����!K����!xX��>�N��5���\�6�9�!'f_tJ�Z�&��y��)]^:��ۣ�n�o� ��\۱z�A*]�=�@�;���ޣ�*ކ�hfn�f=�:X`ͷ���໭?!��
5�j�����]+��5�n�Be	���㙬��q[GD�rl����ѻ��j��>c���T�8���f�304�0C�A6r4�WS��Ͳy�WQY�v�IN�[s��x�N�,��������x���ٽ����o�ZRs�w}7�upo"��1W��I$�I$�I$�I$�I;������2
TF�5��i�h�הd�JW�I]L���E��
��)�.p@�9u�({����m ��Y�,̿{�#� w7���껊$���l�(G �/)�B=�t��ت��ZNF�	K���TG���DV����ް=�'~�O7������n~R�í���� 	�H�!{)O:��@���{��#[ߘ��Z%F��A<�Pj�J��"dV����G'p�{���CH+P�<�Ρ<�����7�w�ڬ��=̊�̗R�{�W�=ꞻ�۸DB�U8M��]�|�!�*��y��d��7ܫn=EC�����W�P�"�}�R����'j�n�p}@ :��Bܥ^�TR�&o/g��z�rTΨC��Q�y�ju���=�;�vQ=�z�p";��������H����_�(�'�~B{���'�?�����L? QP����N������??ֿOӼ��λ�N��I�f��iw���gF�C��YN,�R�q�s�H[ʫ6�Vf�Y	r�wTB�a����v�5Y�P@��%����6JJ�SZ�}��,�z%f	m��O6��tǝC���c��՘�����I�n�3!�ה�:��#qСU�W$�#/�����Pj�Ԉ�����=j��4=07��u�\ww�֤�?h���<��'��S�I�B���~ŝ���"�(o��k�+�F�_mK��ݩ��tv%=����ZkeԬ�*$��������Xm�m����.k�r,\F�C�,�j�n���9UVB(1Den�l����U���}���6+�4����V#Y�P��$h����s��u^��p���m��)��`�]���X��8m:�������Uٽy�ܲ�R��+r��*EAec��^��5�ueoj��w\\�Z}�N�Z2��"b����+��f�\�Z]-��Tܥ�2���}�F3@ \o�m/rf3��AT-����G��;�K�ɖ{w;�
���.U��橣��qK���0)���1��2�|�~�?/z�뎺뮽:뮺�Ӯ�뎺뮸뮺�Ӯ��n�뮺��u�]u�]}tu�]u�]u�]c��뮺�룮�뮺�㮴뮎��n��n�뮺�뮺㮺�n�뮺��u�]u�_u�]u�\u�]u��]i�]u�]|tu�Zi�_]c��뮺믮��]u�]u�]u��뮺믮��뮺뮺�뮺�u�]u�Z}u�]u��]u��u�]u��]u�]zfi;�tn��P��L�cFn���T|j����^��_t͎��__Ll�/$�c�]��0hЌ3��,9;]f����9��wI(���O����T+�&l`sn�rXP�H S8Py�����[)�|=�]�ǲ�	����w}�W}y�����<�V����O4�<�a��i˼�UiZR��x�9/�^>�ͪ<f5�F�ٺ)20��x��U��#]rv�[����Fa��Iʳ;a���+�1d�Ji�D���s2��4,���
T1�3���ԨP����ab���P�1;��͝���f�l�q5����#ч��h\�c��wHV�d�م�L��6�U��o�ம�iFZ2)�w9��}���%m�O���V���ȭ��nX!n'�͞�5��a��؇&�T�p�}'hu�<3�kl��眭L�䇲��`R�o��dR�FR� Z�Z9��J��i�=h
S��<=.#x��vb�7^S�wb�t�"�RT�fOa�4���ɲa9��[9z)8uج�+�[�*�݃2����l����+m�uJH�m�V�ԯȯqn�q I��M_�E���X��q����7@oU��3�\���S����A3f��l��������뮺�n��n�뮺믎�Ӯ�뮺�뮶뮺�N��:�:뮺믎��N�뮺�㮺�n�뮺��u�]u�]}tu�]u�]u��:뮺뮾:�N�뮸�:뭺:뮺뮺��u�]u׷]u�]u�\u�]u��]i��i�]u�]u�]u�]i�]u�]|u�]m�]u�^�u�[u�]u׷]u��u�]u��]u�u�]zu�]uק]u�u�Zt:���}.v�8���rn��۽�p�Bs9ne�c�\�S�&��Ǹ�qƲ�{��L�"*o]Lv�rp��]Ԭ�pLך��\ۀ˅�7�O2���͘�"o�@��Vu.���訞��)Xa޾�.��Q�g)�@��Q�O_�Gebs�9Evf#J�pŵ�n�U���-WS�ν�R'�)&��s���1����c���>x�N+Bޕ��z�چ�I�m�Aۚ�ή��Dwdܬ�Ǎ8�l��R�t��z��F�-�DH͏s��:�F�ž�~�U\��@ޜ�ɬ��\uaP�uX�Ӿ����0�\��|���M���0�;��Z�v2vL[�#q�W�C���#݋�,��m#ӆT�ݱ����V3^<@���Jw]\�k�	��5�a�A�7�.�x�l�o�З��v�cÜ.m�v
6�)�g^u��x��Ü�I�
�I-v L�Ka:���ħ�,pN�U��qJ�.�uv���\���đ��١�`���R��^i
�t��v/p��}�.9e:!\p�͕�3�5c[�2]dn"czR�J�M�
�+7[�|&Ǵ%K�ms�zi��^���뮺뮾��]u�]u�]tu�]u�]u���:뮺뮾:�N�뮸뮺�Ӯ�뮽:뮸뮺�N��:뮶뮺�n��]u�]u��G]u�]u�]tu�]uק]u�u֝u�]u��G]u�]u�_]m�]u�]|{u�[u�]m��u�]u��u�]u��]u�^�u�\u�]uק]u�u�]u��]u�]u�]u��]m�]u�]u��Zu�]u�]|u֝�{�����,���v�K~��E�U�@�������h'�7Zf�
�Ǝ�r�fmk�K2���y&\o�L$&Uu}~�� ԝGr;�5+�/�<��]�u�eS�C���+e�}�=}��4u�̓69[�s*Ku�6m��a�fi4�mK�ѫLU{a�8�W3��5��1/D�Мɩs\[�B ��|ԣC)@��=�]���IE�ҕG�@��S��{F��қ�n���rI%VC��Wk�ͻj�Bu��llWp5;a�0l���`�ؠ��t�龗J@�;fݚ���{�<<���`�6�Δ.��,9�Bԕ
'�C:��]�8d�p��ٜ�j���v��|jZ��Z8��݈�Ժ�YRdC(!ThV�I���;�T�}D�g^�Wi��.��l�����t+��c ���6�L�;	�p����[ Ve:���X�ez��O�*�7i�y��+}\�և��ѱ�������5R�]�wN�Fm��.����T�ը85J��m����J��Ӣ�eT�3&>'p�_;�j�]���<k]��^�ZE�4��f^��7��t�0��	�g��Cj��~��9��h;��E[zEC����oq�I�����b��z�N^^*�UOw�������뮺믮��N�뮺�㮺Ӯ�뮺��u�]u�]}tu�]u�]|u֝u�_]c��:�N�뮺믎�Ӯ�뮽:뮸뮺뎺뮽:뮶뮺�n��]u�]|u�[u�]u�]u�^�u֝u�]u��G]u�]u�_]c���o�8�:뮺�n��n�뮺믎�Ӯ�뮺믮��]u�]u��Zu�]u�]u�G]u�]u�]u�:뮺뮾��u�Z3�s���ᚩ��^P�"���Cg�#�z�����Ɩp���9hu�t�n���w("\���:Xt۸^x �,��k�5�R�fخ�q9y8ںuӻ�2>�:�s:��G_Y.��msn��	�KM��+ms�]��R'b�|\�c&���·v0*u1^:w2�`��{�W�}ttE�D�J`��k^$L���R�V��5ӰFF��-�{z�-
�"JT��
�zc/B�klu� ��}����:�����B^��-�DVVb�K�/��X�S���K�{�య
9v̧��BE%�=�87G��Չ�o;�ٺB��_>�-
݀+q�!�m[�{މ�sdD�Fk�wn9r���}���IM�z����E-d���F�Ԯ�^�(��U��`�%��oZ��;�nԠƲ�y��uٔj.�=�Zgf�7x��hÎ�0V�CC =.X8F*��l���]��,��b��J#J�MH����.��)���R��Ƿ:Om��q��J���k��ܐӋ��oE�8Y6C���ZV���9�ѽx&G,7s�-&�޺�}oY4�{����AR���D�	o]V�R���ڻ����z�#��S��*��f+��x�U-b���ʸ�1
�N�x�f�d%���X[]��k�p Κ#Gm��@��zX��Pӹ���g��D��1tU�օ���]��[&>ECuݲ��"�������(�%in�0Rc���͋�X���(�w�C+e����/ӝ�l�*���\���/��=��aJ�Ǝg{F�z�RR��	3vQ��c{E�z�={a��l�v�z��%��z��UU�Z1e+�3�rꛣo,�s���rK�F\5Y+�p.4|&����j��{�1I`�|����̼��Nc)�РX�B��Ĝ��ݡ�P7KٌǬ���r���:-����A�4�@�A�g����N������po=Aʿ�^�_ɑ\H*���({;�W���%m�q���YMYw�sm�A����٩���0oV` Ĭ���gV�R���t��KNoj58-�aZ�g���*v������S�Qї��K���˝�-�BZ�,v�j���y{f� І����u�ڞR8����4��
��'gޜ�;qvu�t�����7�
j4���zX�Iz��;+ZN;{��]ݼ�HA�E��h,uw�����cDj���j�a�n�fyUZ��v�<vCK+&2��2&�Y݉M̹���v�Rk_e�CA*�5v�n���(�)�r�����m.�T`P�0$�3Q��WEZ�9ezb�z��O=�-�}��*�nwS9��̓�����zn8�D@js{�����ǋ�9�o!tһ{�+��Y��2�;��A��cW���j�(�}\0��T��(��yu-�ݬ+��%��zU�:��{�S��EX���M��z�Mۺ{l����v.��&���F��X��2�	yJN�u����v�B��2J���ޙوmiVڱX�!@
�Q�Md9hoK�)i
Ԑč˃�KUV{�}�X�q�^���rei����F�4����<�i�ѱöQX�k�;�쮺�T�6N�eiAc&�����v��&��p��{UJ�;ަu�G&�$>U�Qm������BE5���<��
<�U��Z�^+��N���ܺ5؅�tI�O�!���$�yg&>�[�l�u�m]X��#��SX�m׽�\�Lz�(?m���[,�9Wt����M��»��i;�}��GY1�)�n���
W7�6X�d5~�j']�fB=�Z�Gj�9����2�p*�e�yӮ��+�h�i��u�a���B����Ϻu7��z��C"{��vV�*�{B:J�5W)�f)�ok�������3�	�d�WZ�C�pU�ڝÎ(�q^ܘ�T�O��ja˴��4%{%ZVk*9�ria�ə.�M5R�	~�[W����ǹ�\l$JZ:U�T����\�K|�ԙ�XM1��_[PF����{h�T����o�ӯ3;Z�֜Y0[,nG 9{�c�Ԯ�xHξ�^�V1��'
�YR"U�S�������h;�-���xb�U˗�F�ݍ� 	v��޵[�R�DKY�fJ��wN-�&L�Tb5��50�3�mn֑�T�]���+p�u�6�{���V^�nVκ�qK����H�|�t�J2��N�
�X�ȷz�1 �&N�ZYV���0.���-��i9���V亗��ܝI�(�C86��:ѐĶ����R��-B9����ov�<�	�n��;݈J//2MՕ���!	��_e��]�o���{ˎ��;:V�ԉ�/�'�������NM�ũ�� ����}�a�3�p�1;CV��"�y��ٔ��D��yd,��WC��d,V�6�(!�l\.�unU��w2���F'fEp�6d4w��W�\0���JgT����P�/|MFF�	s"����P�Mk�.�f�>�NK�
½7�{õ��R`�#{I��������Wώ�Ѣ��b�0_2jF�6e*����6v8�fޙ�А���y٬��+5���F����PL�V��b���i�pe�G*��.�p]N���	���ۗB[�����O���H�sq��f��j�Zu1l^�cZ��1˰�<p��f�`���!�p�DN���껨�vn�U���^�Z�:�ַ0r����t��'5}fv�Ro&Y��p�G��qV�^�׍c��>H��zp�M\uֺ��h4�����0u͝���<̧eBW1s��Թ/�с�8R�+�}��t�EU�<��|)\/�cܤ($�n��+32pb`���TmU,jiL5����bZfib�y*̂VEJƚ���u�;u,��Rwz�6�Ufi�0uUJW�I]} 7���"[��л��NU�:e]=���l����,�W��t��\2��z﷭�It�i r�֜^T���]9����װ���F*�"8�]a�ܬY	��V�c���QBOsCE$3���'$��X�)�حU�<�oW]q#M�C}�nN��T-���2�&�ldIDx��&����Q�YҲ�h�J��`�'����6�^�S9J-�.����&%`��j��R�-�O�Ex�5������ʮF���i��/u��`�tl9�-�5X#�|�,Mi�Uz��
�LX���ՌU3,��.I�8ۢ���=W��/�B�{t�o2�YrQ��ޕN�wY'g�Iz�S#*�JZogX�p���j�ս�\U;��U��.�>VK6�N��6�PR��<[W���)��U>��+nc�X4>%3f�+W=�T`޻���~£�(��4���Y���i:k�|
c3�C�.S��;���Z�7:�%�a�ؓ5�	�D;��{��s���q�KWR���6�e^�{ ҴV�Q�+�N�2���ӫ��r�ӡi�G}VJ�Csy�X�-��R��gQ����SU-Z�)r��S���Pr�����yz�sA��r��M	����w�z��}қ�Vvި�v�/��n��vDV�ݝ����N�cڮ�[�,�V'[�v��YZ��hK ��LXFIe���0���r��L�J������h����@{����W�~���o�Z�������+�?t��:�W�&� ��M9�\,��m�2/ߩ) �e��D�q'4 �	jFI��3QB�j'19�)<D$Z(8��DdEBN2�mE#l��!A���&2�H&��$�,�Bt\f��DB������.\-���Q�)�7�j�
1�q��t�Hi�iBY�#��R�j0Y	��u<FF�('&I_ܧ	��Z��!9���D8����4�mD8�1��1(HL��(� ��D4�C"9�"KE��i6D6�-�eBl��ё��F���$H���D�N�	�4#B�TYU"�C��q���t��$U��Y�W# ��R�"H*H�)�'i�<۴YaQIƉ�q�m	��"��I5"�tV���h������w39�V����]���6n�x�a��k`r5��[��oKcW�%�32���6���V��O�� ���@ͻ�T�"#�A7vȝ�H�)J�8�T-�l�
DEC�WMo2��ܬ�X�,�[v�f�IL���\m�q\�<}t�7�Wڮ�z���n
%�{�S�0�����/��X��������2=�f��+�37N�`�"����;h���������nr�!���xej�5��݇����ٲ�Ө#c�R�\�F�n�	bF�T�!L�,�iK۱��]wQ�Ѹ!�f�:Wq���A�27��KVb7c�5�e�XmC�O� 2��ͩB�nә�ة;|u+�f��ZB���_
�X�Y"W�;L�o5�Yi�n�k���D�/��|%T��(#W5v���&��;$�N7YA�:u�--��dʺN�C{ӳ4H����׷w��u����SghM	+���9�],���N&�_qX�Iy-S뛒�Iƈe������*��䋎��efU��VX{9=��ocʝ(a(#$��wnq���z�v�tXL#�DG!�8��RlH�4In!N����	�B5b�G��@-����q��BM�aȄ\l�|�Ri��H�E�i`Q��'��bPd��% �9
�N2��J-@�F8����q���4�Ap�I� ��*E@O
m0C�4X7U����2T���Q�J>��]�� !7!���I��26AP�
P�""I���A@�l��T<��M
!#E:q���i�?]�-�8LF�(� Q�ȍ2j> ��%��2\*4�b2TQ�Hm��$��BE
�hQ%#H��t�H�#rTLF�)!�D@Jp8�b����. �d�A(�pA"a�
��`�T0�7A4G[f�H(�
�jA���(�`����LD ��D��$��7�9�2HH�AQ�tU@1*(Ѐ�a(����l0DM�$-�p�� Q�Bh�P20�e�-E'�4��o�Cȁ|.�CJ�pD D�,.�a��9&��\I2�J��Kn�Q��F>6
��Q�۶�R�ʑEL�I����R��FK��БƜH Љ��e8�FrcD�.��d��)6�S�H�H�I�,���"4��aȄ\l����0�P!(&��%&H�F'k�'	�(X`�(�#FD�Q��Su!"I<0���,1��C�4�4�H$�PI b���	Sp�#��$��.IΛg�ϥ��5�ݪH�����ooo����뮺�OOOOON��蛲�@�FI�'�oj�N�:ON���w@W�v���]��뮎�뮺������뮺zM�Y]ds���v�����BVa�jm�ڏ�v�w��u�]u��]u�^������u�D����v�DSm�mgggr-eV�r�v5d���uV�d�k�������M���;��Ǐ>�:뮺������Ӯ������S�^QGwI{c����8�.�;��y�U����N��rD���wQvP��J;���9�t��5ۏ�^󪳺�4�՝�M�ֺ�'C-�Vm��Y�Vsn��	A�Yl��iu�P�m�V~o�Wwǧg`�wb�6[F��V��*�ٞ[��Y�J�\_[�������S��ۮkv�`F͛R�e��o��ڶ��ǽ�^�Y��ny��6dV�'ͻյ�j�(��{6���7���d��׵��v����ny6�KKE�A����rW�[洪K}�{�m�w'G^�+/�_[�8KƗT���fD8q_N;<� �������G|V�e�)$$:��IQd*T}�e�2B6AM�I,8㌢�� P��
B܂7%�Z��<$��!�%EDh�"Z&&bq��m��2ё��x/�އ�WC.�.m@x��55r]�ɽ�ø�ƅ���=y'9�N�(���<-��q�)�g{;ނ�Rd�E$L7�-��#0�(I�!I��`�!`�f�"IH%4@A
P��Q6%i��D��!|��I�I'	L"cA8@A�Fq@�e�$j2��(�!���P�ےq�!�b��6�E��dʙ���Ve̻��m�c��ꭧ�����ܺ{��<V��qu���(s �%GR]�K)ڥ�F��(QH���6�`K�Pq�cwp�f]zS[��OAY�Z��.����w���J�e��FZ��y�cԬJV�[Qu4�T��}p|�6a��f#k^Tו�"*��1���QL���f�"f�Nf�7a-�%��B��&�T���� V�[�Qws�)!-S(���jF5��a��/� ����?eS�\���Jo��EZ^����&g��ڳ�Sy��zR���>�.^.C����gc3"��ᤷTߩ���)�n��Tsԝ>����|������Z�D�M�±l`��t�r�T��ؐoJQ��� ����q��3��:"���Qݬ�����z�a	Y1J�W��>��I"fiS�VPƻ�`�m�T��9��Ǜ�A�q���Q;&]\{Ѣc>��!�g
0�#*E\=����2�"^�9��vp!��U�V;h�6\܆R"e��'k�?v����h������w��#�>�Q����'�m�����'^1�.�4{ND��L�8B↡-�#��2zr<MS^�D4z#��}D���������"kd��*��wo����+H�q�N�yp�_��t�-�kT&2�%��UM��J[^�0m�L��S�!k:�^�r��ө��6���S,�fxB�xXo;<̫�p�F������9�[U�Q���oչhD��o\��F፹"F7�E8��qp�Q�T��I.&�5�]���'��	��&I�k�%-�6�C�j�wN0CnCB��G�O�O�" �Y"�`Ɂz6r�J0qnl�F�w�����5P��KoU�8*�P�V��ףa����6�ה�Фk6qJKyҕ�[�)���vpƽ��%�i�\j���C�Z��uZ��N�3ԩ,,��c�]����t�5�c��YL���:��F���XPV��4eH	7��4e��(
�_}]G��p�>���霌�3'$r�p��ah��ȝ�E��:8
�7�&�Q�2��T�.�a2u+;�>�.���S��\eΝ�˽�t�+�-9��sMuv���Vԋz��WE����ʳې=��?�U"�� �yx�����|@8��vvI�*E#�߼�+��Ғ��*f��Fsij	���{چ�vZic1��j���.�_����BC`;�{�F��F�-�MeB[���/6��[0�C�,gֱ���DE��y��fs2���-�����^}�ݪ�x�]����/?��q>(�_�����QD��6�UO�4�(&�	���f}n<:�g�?
~%��zќ��8t�[T������
~^��3��_s�w�( A��;��Spv���v`SE�Z��-�T���`������ԡ���f�m��E-������B�c_,��|�zK�hE��NP$���I��gg�r�-�P�8��
->��L���a���T��%BQ[��«�����P3A(z����*��f\8MQ�ܧa4u�B9��^�StW�8�Ő���yVc�(�j�kl�æ*&���=)]�+�܆U��Z҈M8��)p7�ٗ8�ЦL�um�<�cXH9Z���'P���7n8\;{O��M��l�����+����������Ω��j V����]a&�N�=zO��E�m,���������H�f��h���v
�f|v��m[�m>@��v��7Z~�No��� �I�/ɣ�a�5@W�=��^�)�R�>eçBnlR����%Z1��[�����12X/��*BD�2X��ˉ��Z�pMԦ�x=pه8|��#a=����ջL�S�:w0m=HMd�,�e���>;;,1����Z2�O�PFүK�$j`��kM�k�G]��AMa�D����ޥ<�Q���iw��q���{J-%���Wm)���4�f�W�_�G1�=���'>s�-��X�wo\��IW�"n�ǲ|v�v�=���0��5�T��DǐC}�ϙ�y�TN�>K(k����;H�8�J��CT]]8��Ӛ���5�(A
t�iw�1n`��=�W7�Տ�'�Cs��G�����Y��'���m�A8�#x�L߳^W|�:�6�'S����*�14;������ؙ���|�v�����-oc��Fx�|||||}�M����6J�;1�:�&ܼ����M�ҫ�n���*奼�/����j��]�-fNF�UUX�|  `¬|�W1��A���'2�z��/�1��x�cum��R*��p�&0^�"�'^�u�g�խ�����ie�S�E�MP[`�/m��y|�,*��V�����z����Yw�g. �$�HJxv�C�����Qca�X.���ڮ+��L�����&��׎ ,<z�v�b�>��k=�[����(Z���8r(�{���=W�c1�s}B�d���U&#j���Q�5�
��z��e�@^�zё��(�L�H����*
/u���YƘm�U�x���r}�_\'[�5]B�ʋ�LTF��̸wv��=ɕ�Hl�6A^���C���}��ñ��rA�N�o5&��(M��JN�4%q��w��H(џ�З����[�jdZ�t�2l��aߠh+��F_�C�޽e_���d�y.���r�wGp�[^�CJ�!Rꞥ��]�J�t'!r'S�T���@s��F�SV����O]`�譎�N�ތ�M�nD�#�<<<<<<=[��5�p���뿲�LR�$��	!jw����c���j�/u�RGU���l;��W���F@:�4��0fSA"@����&�a��f���*�N�DC�̩���8�,�DBk�	7�Ū���׻����T�lLL�#�:����Q��6\�Iew�h˶�"��Eٜ��BJ��a�;Y���A%48�'��>��a��Ln�&��-,L^I�t�m���G����y���}�no,t.i�k��?���,P$S���ۿ}�5����X�7Ic�(�0���ɶ�I�(���z�,��짫i�xf �^��j���ڤrf�K$�&i�@�
}N���>Ǧ]%9�v	'@Ƣ�d4Ĝe�z��٤&��c�Y�A���a�!G���"#�z6-�Ҽ�v��.Y	��N�M�͖������`�?�yu���N���t���|�������SoN���3������Y��eׯ���m�����\U�g���Ib���ق�r�W3D�vP�*ջ�b���9� ��ufv߻�������^@G)������-T���~��t�_9�3�}r�].��Ͼ�K�]��>��]ju�%f��5`�/`y� )JP�w&��5@.�ӣt��mF�Xe�V��b���N�v[#Uy)RJ�>\�N��p�+�yJ�5��ejċe��$���@P��v:h6ߩPJ�A6e��^�*M��KrG�D;�����u��+`V��&��ɽ��ע���U��w�J�I��sM朿9MdW�8��ɍ��J#)dm� �gk��0�d�8A�5lY���^W�c���⸀2.� N��D��Z��rd�M��@�f�eNEײ�� ���>fFc,6w6�4�J}�dQ ��o��W_���7�9��ܖ1��0��������L��u��f�F��\8:�<ncN:�3�H$����g��)T1~+��`����Ճq����n>��@�v�Y!x��(���n�9��g"����͛���X��k��:�L�N�8o\�]���c�`<�#�]gp���՗�.�r����*��rcͫ�;���O������o):t�T4�/�l�E��m��sv'$�,��ʌ�c�Q�c�`Ѕ�<i^�E\��Lk哚����
���uE�v�}�o7�|1�x*��v�K.*"O�G_F����d��r�I����������F�1햠h$�1�Ggb|���;[10�x��9JÞ5*��[A&�|v��Pk> ���ȍH�*;:�y���L
����_L��{���^͹��l�kE�z��]�Ei�{`��;R	�dB0)O��#�a�I)%U�cY�ݒ%�5o�<��:�Z�Ǟ��"�R,D���Ӿ��u:3Q
r���R��x��i#1����g�J*k�~^�}�0|��i�
|L��ܣ��_-Nƪ����M�r<cF�q�5?�S�r1�������xVؗ
r�]��ð����im�_}����&]�J���=D���a�&��������R���@
 ��/;��U�_n�Rl�&����p�S,]�=�	��]���&�]Tӻ�{��]g�׻�E��1��%�;Ԧ,:v��TonRl�hC���f��e�w|Gj�B�{3��uE�k
em[����8�V�����H�I�/שe�����ϦS	}��b�3V�����Hڥ����S�n����{�~y=�{��|t+=,K�r]Q� ���Km��W�B��������S��v�q�mݰ��Z���sJp�W�X�^q^X��>�
S���W�ihk���F�+ɭ�'l��Q4�a A��c��4�4,�a���T�f���zq��1j�]s��@ܥ���Q��=p΁1�f�Z�撫TN�Q��mք"U�EA�:ªV���+hMzE�>`�!�E��5�l:��YPSejU��Jڌ3~"���:�q�_,h"�>K�P��{�E�D3�9-;�w�.t[�xV߷v�7�Ħ�f�Qm�2�^r�e#2�
}�|�Ԧd�U��7_W��9�H���D会�T+xn�>.����_S���k��%��f)[f]�'FYڸ|���ڧ(;�I�QR��n���.tVb+2��8�A	�ո�ƭp�uZ\2�-� ��|�������K)xxxU  ��f�u�[!W�Y���R�q��p��sz67 �t\�KT�.�GK�ލ��o�Yv�C^�T"��s���S;��j�d.�������7�f	���S�BI
���u8������j��`��j[/�
-��4	��c^T��d6�y�SS�=�ի��W���k1F6�z�����^9�-�T���^Z�eF�f�B�
fq"��-E�g��d_��dElRS#ul�	f�����c���/�Pl��M'�pa��9�Jb=�faf�@���Gb)�qF���v�ޒV����7�l^�}Hg�\���*b`�j�kz�(�xJn�P͌�G`E� ���1����ǟ2}/V35FM���������נn���u�uw���>u��v~�� ��:�|��F��}��E���J����ud)|f椺��ړ:C\+z�L�l����'�B�7\� :�6h����`�z��3��uWT�&��rw
vz�iSt���j���T}��X�^����V��#����s� �㩮,�_:���˔@q�ݷ���3�=V�M�땥���o6%�p����"�ػ��+��Qv�����V�8���C)�J=h�����FrÄ��7j�� �n�Hֽ�[��[NJw��h�D��q�b��C��׹�I΄��Pa×srrZZ�*�;�љ*�Z��.nS��:�GR]@;���D��k޾�c�E�{F)3;m����lr��I#��"r�;��*�_ET���Ɔ]h[;�Oq�%W2.铎�v�rk((re�{X�=3���4"�Y��0\�p�L�e˻�vݽfn��\���6ȅ��4��)V�)r��۽�]�du����t`=XH7#E��%�\s��\��t�=��`�^.�ɮ��tf�ȸ���Fr�&�zsk{�洊�6�4����T��v���P�;>;�����o�@�g�I�`��뭂�ܱB�,rx8V4�\G[��؂�������AeX�U�b�ouI�4�+gGO2����b3��i����m�yZɲ�;U�ձ�˵�y�H,�+TӖ�����n�s�j�S���&;ͼ8҆�k�V������>�$Y������q亽���"��C�]0��յ3{S�v���
%�^�O2��w_]I�r��`aT�K���X��#��e�O��ږ�9���Ug_H
ڢ�ʧp/�^J-w��6ؽڿ�5����I�mi�&�8e^�n=&�bV\{;�`l�=�/oULve��j� 7�c֥��n�gE0	�9��������vڥ�&�%H:�}#�;'^e���q�Xu���N��C#EN���9�:2�r�g�{Y|m�$�=2:��eL)�b^a�:����x�ɶ��Wζi����se	��1����/`��G'T����|�,��X��+���^�e��6�|�Bu��Ľ�Nb��\�4E�4�ظu��I5�we�q�a�4^�!۷'AC��2$�q|�j�T�	�d�h�T.�-yI�k�w}�����;:f�VPn�ͧ�98�dް��wSf�=�;(��d}V�/	l�Zܶ&1T�V�(Z[��n��%��<��v���Ȋ�䔇;�wS���L���nC6M� ��-�i�[������p�킧n����ˠ
�N�ʡ�cFC�d.0o�(�#�d㣎�wv{�p4�	Eq �	�I)��3��.��'VZ=��j��Hӏ�>�x��뮺�8㎼x��6'�	ʐ�BF:�~�@����(?��!p*�*��H�M�=�}x����]u�q�u�^<�FH@��ݤ�n��y݉Yƕ$!!�P�:iǧ��<x����]u�q�]u�M��(�$��)����:ˠ�����։�g�Q$K��@��6���ǎ�}x�<x��8뮺��ª{0�BI�i�������{|���S�5��pH�:�nve�a}+H��8����]>K\K03�ghJrDAA'rs�ND~�};⒠����kp�	{s��ے_��;������{n����'�c�E�~sI||w�8����p������J:D㿎����N���?�"�k�$xq_,.f��E�%ƧP����7��+)-*����Mw6�ifv'mA(#F����<}M4�M4�N��s�g��9�'$���/Ȭ��W2��sڰwK���W�!蓥��+���+;~�L@�3��}X�4� �4�7����kЗ��^O�`��	܄�o�|����-:Q�v�8`�Oy�������\�����0,�
�,�x��w���qꔨ����tȭr<�ӱlm�Na�Ij�C{h���<=�M�σ��'������֕aH�x���,>��\O=�J���� ��Z��V��Yuw�~�P� 9�[.J�eU`>�p���:�b�V�)r��P�+�b�,8x.rW(}������{#�6����� �1;v���!{�f��p耟Ó�~�\�n����O0�j�򔀴�0Ǔ� xo/�a��Le�O��nt���ia��X!5@~Z}\�{8ί y��w�gl{��d1됀���2 Ǻ�6�j�K�f�wz� 8O�����pj�ä
���eO'������Ro�$��o�q����&��Ͻ^�u�����ԉ��Q��\9�`t�����`o�W;�����ނ�-��ϓ7���^n�^y3�z��'�kN��x�$
`���Z@�<K�!*���p��k8/�8@�������V���`o*�a�>x�Z��Z�C]EҡRY.�u��\��o�$��C�Y�	;C$�
`)��i��AX�ٝ��i��8�b0M��'r��b��A�.��c%��ep�c2�i
u`��]G;l���{�������{���Q0�0��İ/�z8�6:���ig����bc���x��#���`7��x%�_����v;e���� |7y�B�����\���C�~��9���!�W��F�����v�iw/�t�]����D30z�C�8ȥ�>�U���c�$������m����;t�� h ܇|�>2��3﻽�Ü�Bq|`5�:���4��/�2	W\��K�������',�		�$)��TL�(������o�8� >�;�����պ��vO�cǮ��ݟK�`i�L0	��3
��3˘Cq�ӻ�����z�v^
��ze�����q{� a���;Sg��>�Nu�^��wSf��������vf��kRz姽<|�X������*>�v.Y�-7�[ha�Э������H<yP_}����լY_(6��������� 
N[�1l��[epq?���*\=�	oCJ �ᮚ���@�ف-^�	+���� U�[z���m����Ѳ�"�")���]��:�{��'M׼���XŠѝ��j��+�Ro
j\[>��k��e)痩�b�m�B� ʛ�V����*>|,�ٓ��n�/h�9�۬-U}Yv���u�6���3c��ĵleK&���n"x���x��8E����}������m�ټ���s#����zν'2�|󻳎<
i���i����߽��|���m �ӎZ��EIy��8������tUお��"���TYe��y�;� 9ϳw{P�R���Vx-|�#��9hh|��e���Q��p{WE~�����J6��7v�M)�N��x
Ƕj-�����y�Pxd˟���|`44��tt����nWWնml�p�c���t��]�{-�O�>輸��ĩ+<�ȃ�<�����5[ŭ:|{�Ϫ>�>uC`�����n\<��>k�-u�O�Ø
r<���$S	Q�4<������_����߷=C���6�W�㱧�����:�����{�^�<��z�����NصZ^D!�'7�L���2�k�[�����)�L)��0��H��_�u��/��>�gO�!��se�e)Yy	"Xp���h`�X0N��c��@��dF����	��p;�'�^�ff�	�u�T-W*'ifw�������k>]�(�	gS�nl��;�0wW�,P��>`3�~O~����xI�\�j9��vU�map��yg%ݢ!nJ����>0��	�j(��мx1.3�[q�|��ۯO��_�;ѥCz�L��o���v��^ߐ���]����
A�Y�}hw��G��<��6~��º�1����<���Ws���B�n���Ktǹ��8�w{���#���-��o+c���x���=c۽�g����j� �8�5W�D����qI)oQ|;]�Ήu��Vi�8�]��Z�9��j����ɶ�ۖ�M�m��HNy���wϟ9�!*Md�����7����p�ʓ�|,W�S�����G�H�$����B�u[g**�{/���������z/���0i���xj����X)P�M�ۖ��Á#^Y�c���[��^ `�� �dN��a��y����FL4;�������61��˭~�y5����W*Jsc�W���������ڛ? k���|�?u��*A���hR|u��h�y��=�=����c�Y�Ui�(ٮ5��.n6>�� ՞|>}�����͊�ƌ��]|) � ��{zx��`.z���03���±NWx�A ?/ueǍt�I[k��3A�ˀ֢]���ި�2߭�%�=�� ���`��V�/w1�议 ��Cy��+:'M�����9��z���{��yO�)�2.��⛻O�x(}�,����;�f�6��nhy����V,�x8N=��@�p���R%\rqI���(�r�Χ��7� SU�ki��F��Q-�=���Kv��,~|/ٗW�t{f=�
�OQ���5�hwW�.N�g���#u�n��e	k/P�}�q����崈�ki�sf�F�J��6�	��ὲ�@�3�h�>�,!u��Q��,�:�8�e<�8�Yb)��s�9�Wd��Gz��Z�W%�$���h�����&�����N6����i����Aq�@<�h�³;x 2-�5ȶ���9�����5���6��(�s��p<�|$n��8%�5��ӯ��<�x]����G�
�<2��a6�k������ƏW�jp��B�ݯ�wW�x��w'#w����3�|�R=:��ҍτ���D��iVp���b����<���>ۧ':�/?� z��[k��_��	��=���S�w��en���Ʊ��;[;��<�CxVwE2���qG��+=� &��GnUD<�ߐY\@o�l���e}��^>��C���"*i[kd�8����I 	ig��(f��g�x��UZ��qT���nJa7;�A ��1�Ĕ#)�����7�ޜ���y�y��֖���\Rx�q�=R� X��ޮ��=v�� 7�(ނ���9����\?n�Մ
+ٰR)���xH�?}�g���L�kW�m��$R�l�~'_��I�6	�M� �Z�.��oK�w^�=b`b�h�<<ŞX,����SU�~8�5E�����\ />`4�n	�o&ؚ��>���Su��^�w���x�8*���$ �b9�{��"��}Vm�B�w��z�(2�����ɽ����Йי7#	U��=�����N|䆎諏:Zt�z�a��aɮ���Sf�.J�;)`� J�.4;-�=Y�Ѻ�;���˾Z��j��_����m��m��-��D�"�2) "X��;���>{�j{��Ϩ�)G��y���t��ׂ�Gt�noP�����r|$�\?B�f����zΛF�z�{�tgY!�4	|a��ml��u���m
m��O�u��6l�Je�c��=%T4D3<_���2y�Y~n�c�����|��R�@	ޘt&��Y'IE�]]�%t5�a,���������"�ߡ04�$��[�>;��|>B4Ϗ4��������e��������8��<9�n'��b��V�˩p|RS�x=��x{�&@����u�_���v�O+�g,���`��T�\���osU����g��Ć^�-�]��o�MG�[�g�Ü
wz[��T�~�8YJ�5�2u��@i i��/�d	����^cW�#5Vg�i����]�~�f���x�3��x��
Y5Ô���a��
��ZT�M��Յ1~O����ybb�����;���3��6���0o�|�"`���0>o���Ǹ�)��Aròj�{�?^�1�E�Lg���n���Aٜ�Qz�$�A\�Қ��cW9C y�I�㋜1i�ӻ:��c�E�y:��{FU��y[�j���]�@��׮�i�ٸd0��b�C�޶�0,�|��jZV2�ɂ��6;��;��Q�c^�3��Kx�/��e�B7�Mu�$�Y��C���P���������l[m��K��`ȠH���)�y;�s{u2�R�#RHl�QO�8�A�����o�ݲV��\-��Lӷ%�A�.�u���A�@~	L|��4@ϗM�P�㤙�k�Aσ�6�ܞ)ǣ��ܱp�L������Q�<�7s�?�ҍ8���#!��m�Ζ����`^��E및^��o�=M����
� [@�MM>��Ū�	d��`>ۊ�a�{��ο�ս���gz�J7�x@��p�'��
���}��<��vy^���H܂���|%B��Y#���1;��ե�W�~�����R�Kԫ�����N�=�uY��|����=<�,�,jz;b�-ė��:��յ;ǀ�k�C<I�\��V�9��9A����˂�qt�4y�/������K3��O)�u�9�L���xKG�9��㤔��ު�y�\��H|���T92ƍp$s�[�����^����<��uq @u{�����S��W�� �]�Iv3�a���|�ϟlf�����=S.Ꮶ���D�z��[��t�T.s� &T����� nC�ϝ�6g���˥wn�#�=�t�� ����+�*z|0�ɔ��-�B����u�`*����p7�1l��8��U�Q8>��ZD��k���L�����lNUj��'�6b���J���s����=��_I��%Ty�[�F5�y�o$�YC��{	ޑ^j�O��Of),t�8��\�hݧ.����-c�ë�|���O���@���h���j\���m�ڢ\I:��=k�Wz�0o�{`6X9g���ŽR�YM��xS�v;���z`;���a��T�={����)��old�y��+ïLk���$@>��:Gƀ�_�"�4��sP��&��~y'��a������X8��o����x�����t��,�!	�����Z'� :-z�vvn�!�1V�&�=V�8�OC�z���x@Z &����<��o&��݀�{a�3�棌��,�o�����`�o�����B��pv���
�7�s�oC�N��%C(xk�!wfvm��q�0�|uo�������{h���CH��O55>V�^f��Ӧ���V���]#o=�l��|X��[-����{�O�|�<�_ �����
��X�Zx��>�:}�ӹ�iF�S~//4��Jp)�Á0���L�8�rƿ��<���אY:�w$&$�'�#�ɾl4{��U��պ�w��]��S�����,|���7�C&\34?�{���&�q9��MESޗ�������6���Ƽ���7��yo�1W:�����k�r�����k*>6�r�ػ�=]f�CYڃ*��܌f�fv:\gQ�M ��5������){��=(�R^�P�6q4k����(�S4�W�l9Y.0��.(+X���r��t�w)_*�s�(e�)�i����`4)w�o���m�	9,���z�?_m��m��m��n+"��� ,�,�� �+��r��X���	�6���ɼ]�:�C�j�n�ssbˆo]<s渀�|[���p�+�j(;kgoo��0|Ʈ ��x�p9�(#R���,v_f�A`�c�����5+vQ%��r}�I`C�A�Ɨ(�9��!����R|.��[{��s�K��8��aK:��9�����b{������u-��P��!���>�+����.�i�4���"��m ��dkt�U3Q7��5=o��t��xc�6I
pf��>>@R]������<�A~���O��[�ђ[Ý����5Y�n2Pi�/>�������}"z�|6��M�4,��'{|��0��W�H��X;�j10�&�$��%�L�@)���Y�J�E�Z��O��^�=��5 !�	�a�U�W7|��9yи��hck`��/���M�}�es����nn��{QJ�P�"<�����^����ŕ��{xB��;ĻxHcs�w��`g-qߠ�n��_r��񠤪���
	�c���� ��f��(K�;���s+� P��E�����x"�V.��z>~�_�G����Mo�s��ڕy_e�뽍�|�B�R0���\%�j�>�p��VU��)�LM�1޸+�Q�]�R*o_U�c^�ݫ��RS
��!����7qJ��9�P�ú���NT:�K���-�,��ɼ�#s5ێ�;�_ǽ��#����"	m���l@m���
H����	"���	 ����H'\����ߞ_�*�"���>R����=9�@Sz=@��,<�\z�BA�#+�`g���=�!��bINk���^��[�ӵ��ᝀg�U�VW�lघ���0/y �z1��{m�4ù=f�®\���4Kyk�ln��o&IE�Ќf8�z���h	ğ���.�	6��|`�l�*��9�����'��<��K4c���'�%ẟB�4�b{p0n��Z��^�����{�ށn���֮��N�pt�.<:5�����G�����h�@{�V�.��;�Swv��kedNA��m>�fYO�7�k#�rk�%�Q~��1���h=/���*7\OOO'ØLU��\�+2�t�VW��^��P�KjF�A�F�M{�q{��<"(��9���@ކ��k���nd���F&�{�`��;�����9�_�i���6���W+v���a�|�]/�F�duP��n��~��P�٦���<��׏��y����R�����Ɣ�ë�bd-` s�*���!�v�*�~�#Od���z(|�1�N��Rkԧ�Ǉj��_:��κ���g�	ȹ0w�[0�L����#:�f'
FnvrQ瑎����Qw�ߞ�ʁ!��R��^ܙo��}7y��D\]��5T���A�n�8�Z5�BѠ��z$�1�����%�m��g���r\n�+u����n0uk�2�u;˜�1�ڌ!�@yҦ�^�{���HK ��BZ�ˑXy;wK�@������]usT��u�$9)���',j���tqM޲n����K�e�9�<[��@�vc#����QZŇ�l�ԧ`^К�K6���K;�\=y����b��9���>���!��k]�Vj۫��T@0Q�֝s�"��@���܋��ڌA~b�㾩���ǘ�6���dېlը��m��}�z��-١���H��5�ڹ"��"�v�-�Fi��.�3��Yͼ;z�9��xI{�T9լ/.����8��em���;�9��7���ْr���7��G&����6��ѴD��rS�9�:�u.��n����*�J�̔+�`w
��s}t��:X�n��:��z����W@���)FM)�.�w����a�-�Xi��37<��]
��;i�%eZ]�7��{˘^!��9�M9-C "��������m}: �+��V *�Z�I*�
���&m;DA�2"�eW�ʙ���	g�n�u�`�C9�S~B��9�e#mk�*VJ�L;�=ue
�2�[޴�JB�MKS�ݠ%ԉ���X�V�	��}�!��W��s6�Ω�=x���ٌ�4��&��\��o=��Vui<�:��F�y�n��N�,�i�1)��*���VE�9�}τE���}�3���P�[�N췢[B�=.��O��ꖃ�:�ZH��,��֚�"\�ƨn���V˦��2�M��/6�IG��X���x��rZ��L���7�9�'�x�-!�U{:"F�Ǉ�u��iuu���&y'��>�o]2�A�X�8�8�u���zv�+�s.Scntə���mgN��J��(!Չum���:�L�إu7f��g�*p��͵��@�m���o��|ƫR�+��,fN۴��Ιt���-fb��+,@�z����PJT��`�.-��e���dw�F��I�p>�n�x[)�P)����3:�YU������H���.i��qn��5� 7�xgnѶ�y^"�o�M�����/z�����/#��b^�&�+pmC��A]zӭ�x`Nvu�̂�Q2��Π}ڦW�og^�7֚��4��/�9��)���o=�'c��r�T�z�wr�}&�-<S�Jw��S����>>'ǒ>�@F������D!�	����*$x��ǎ�u��ǌx��ǧqǏ:��$�B0�]�"��rvv����#����eaN�������u��]cǏ<{q�x��ǎ�CU�GvY��TI�Gzw_��|�&u��M�9�裏�]u׷]c�������ӏ<x��fq��Q�@ۻ��trw#)��u�]u׷]c���Ƿ�����<x�D�$		��9~4Bw[c���2�5�t[X������]��s۷�s���(����������g6������;�)���J��dۭ���-������XW�ѹ���}��v����Ym���2�#����udrDIF��P>�aNq�iR=���&՗�����]'����:ʈ�(�����e���_0p$���B&�F��l��5�x��BB�BH��1��ep��L8��a�J�6�6��1"r�3i���|b����*gwȧu}:)qUc�e=O�#ް���T���]r�e�85Ey�����Qe��!�D"S1��$��3	���HYl����2F
����bc
�	�xHm���R���A�mD"%�	-�X���"�I�bI�HT!�\0¢|I�`�"��0@d���[*
m���BcP�|J�\� �$A����[��m��")m�F�	m� � ����
g�ߝ��/<���ua��H��qe��NQu�"�Wŀi][�W�-����s����WNдl�(]���pͮ�䌹U/�GU�i���heH���[�t�kw=���i���!�5D���[�x�Fr�U��`����	�֘~m�.��j<3��w8�/�M�GDW��
���YX���U.�i�=-M���)�W�3�AM����/�1�ŗ���2���\� �\�#����әu����v�����= B���"^#}3�0>�������u���qq��ꓰ���U]��i����0>>|�	���7�B,5喥����	��9σ������݉�yM��0SYN�=^�=C���F�}�P��'�H#�ד��W0-�<��{��W��Rmj�ۄ�p~�{�f�"����,�4evr�S.!��� g�O�`
D#��E:��Z�#�zX3 �Q�������yhCP;�X�7��%W�Q�8��ĥ�9˟����W�ߡ�l]��hc�-�R�bs���>Au���q�h��Ɓ���^�%��;�_D���|���T�7�f|��sf|�f{^| @Y����=  ��pZ�M��ڵ���?C�wi��~���e�v�2�Ń����5n�\��0�;n�[δ��0k�=�JkakU;����|�@ʂ�4Q�%
��Yp�	|��bFK�y�qkaǝ\�ʖ�5f�����j���of����w��pm�������b7X�m�\ cm�+p #m��7�ӝl�Re��n)��1��x�}�P�^S���^�#�zo�8�
�'w�cwGw�w;)i��=L0���-X��Lir\	�������ė�p�� f�����,Q�����#���c���E_��ԡ�����=o�qv.:ez۹�wB`qou<y�$^��v���P�IJÕ���?����3�S��͜��yO�*|4��)�%�[û���Z�S�m��#�b2/����=xSS� ��x��p����K�
os����#?|}>�%��l���8Ck>W��s��ª���l��������Mb���"�nEIo�}Ӟm��[]Jp�<�@z�\k<ȇ���S���ͳ�9]�{i%������.�s+�aٓ{�z�r-�.��:u�pL͆cw������fZ���Q&A�L��я.���{4>�bo�E�WpI���\���nd�%�=<�y�8�����A��'p({��$�s8�8��v}N��^#����	p5���n8�##�������V@�ɜ߾$��\�{+������mx�� �)A4#�v�b�ᝧ�Jݜ�飥�Z�(�{Ln�7UO�M�Sd��27�P=��xI��2IK���X}@xxP � ��,W� J�@�_oѴ�������ھ�4�>}%�W4ԛ�Y�s�ke1��I�vd��﮲c�s�I{}�[�_�AT� ���ڂ[m��R6�h�m��
�	 �P	A@�����k���>_�b�~P�����$ڧ��A��Fh��Q�Wjܭ��}�϶�N{w�xKY����0�.�R��;\��σ@���T��Y���`'��NIQv�Ŭ����=V�施ڞ/�}��+�"�]�@e�(��-�'��
 CK�q���֘����G�SSu�� ZQ�/�G60�~��v#g1���~yjw�8����>-��{�J׬#�-��P��v:osl�c��x���^@�����)��G�O�=m6����ZY"����G���'	�Xcp����4�`t���Z�F�]y��φ�tۛ�8'lk=��/K��߀� �� =��64��>��R�8	(�r�;�G�F��k�3�����&m-�=�T9n��BO�v�>��=��Ɵ��i�zpg���=F\�`��nn�O$��"�g%}ڽ��#LT��s �y�r`^�֙�`��t{��3T>cNTe{3R��M�'�uҟAo[]��������`������#������e#�����n��4�kgV�Ѭz��a���lt���4݁��]�ݾ���ՌY�!����\[�{;�o�J�����M��H����8�G��'���Ng��|uwp�v��fm��R�[f��=�� �7���}\?�{��~���(�m� \ �m���m�U�Q�I�|�x��g�;��������������9��R����	�02=�!�C�F3;h���㊈�<d:oS;M����,>m���y�W����n���H4 h�����s&;irGG��{ύ�*1R�ͯx >=��[��@3�*�^��y�n�E���Pt�����(M������<s���0�	����(U�����tƼ}�q��� ��'���g;����5�S�!r���n���վ$~�*eO���E�eG�F��9ŀ���������ֻ1M�Ј�����޹q�c�H=�M��5$r��l�y0�ά��\9��sR��ر��<2Kap|.�u��{���|H����p.	���5zx��_}��>���:�O�B� /<��²�5�>g^a��y�&�����t��l�׎C�,�ɗ�~��)ͽ�i����힝��������\V��k �ʒaE�v^���i=L����u�kj��|��绶�5��s�Grw�v�5U��c_����j�g�>�� 𜞞Ona0��EvN3 �\�����2.��af殺c��+����ޜ顒�����^���_|Ы�ʝ)�2����(�-{�G���y��E��W�K�<���0J��֤�yۧy9��Ƕ��GW�
���.z3�JJ#P��9�m�{?�{��D�<~�\T�m���b7�I�m��T��VD@<�缓����r��2{'�%�¾K�.ڴ��=��Wp:1ߣ8[�b���]��.���{�ɮ�H��SS��|�N��p\
aß��A���k��>i/	� ��6�1�5a�����p�֖��{L_9�n�Z}�P�hf�Hrg��y�fZ¸9`)�0��&��g�Dvi�F͓��z�� c�\����c������UGޛ��<��}f�@LU\L��c����[d�{��iv����;;�x����H�F���[+'��c����a��W�#����Ż��0g��4�c�dor<�-ݚ%���s����{�+�zp]�O�dꜘ}�������aI	$$�c |�Oy�3y�{ʔ8����n��Y��t���|;��[�ZhE�9���<�"�ʆ�Gs����N1�UO]�g�{����՜/�(㥕^>���h|}�|��}�]��=��S���u�l;k r�K��p=3����'��8-t�C�����6u0����gR��X+���m��a0�B#��U������ͮO�{�1�g�f��*3�jv���	�B�
ȱ���y!f_=V�ou��rۯӞ��UŴs���i�g��A�Po&��0-�Т�ۺ�q*�)�'F'x��%�7�{Z�;��r��Fϴ>��8�Į�p�Ջ�P��㺃>
����e�[���H$q�$�����'�Gr�
����k>���9CZc�9�[�6E���f�����pr�dr�
v�j͕u4�w߾K﫻���pP#�����m���H(H�F�l଀$m��� (� w���9ϛ��-p~
���O��\�y��-U�CH��YPIV3�6�
/	�Q�g�rR�o��W5�=Շ>B4�O��69m�jCCN�e��4)j7eGC=e�n����I�U4���nĥ=�vԥew�|#<~Nq�,�4J���N�u�l�dq�SP�<U�\�\��{{�*��Ws�s�NE�u8ސ�ɻ�l:-����vt2�9��%�7�\�}P�/k�y�b��<��ܕx1z/�]�D��`�K���ݙڋp��v����p�9�7Mm�������k��:���(�}�i;0m{w�Z&���{���Gw����q�ßCkL>6ρR��Ձ<�dT�1j9s��^�wL�oT0�wq+q�l�ri��_��wr��^m�J1ǩyOР����@bzK��n�u�Ak��SmJ��ż������ޠAC��="�W����.}��+�u����v;�s����6q�'�\�������'�s����������F�� >��;7\Ԗ	��?+͗֙�4����b]��m�;����R��ZW��5��}ډ����^U��#*a��4+���e_я�}�!���QZ_r�S�X���r�h�:Ջ$[�Y�#á�V�q'���[VF���R7u�r"~�$�G��6�m���m�pd$�m�	qD�I �$$UCߝ�>gϜ���|���e�����3E�8�Ԩ�>2POa�8fЛ�}�9���M��k��o�3+5 <�5[�f���S�����f�}J-�Ξ}�.��@˚lĬ�nv�p� �<�|B��{�	
�)���W|����2w<[}{oW��c��k�v�$����1'�$C�����Uj�Z��I��VBi�!
�>7�I��hu�J�zݼ�m�]���}�G�c֠�X^3����:��|� �AG�B����$V��f�o�����*8������p�U-
u���1�Ei��o�] �_�Q�����L�b�i�?pV�R9���]�xJ�hF3��[�Slᯂ�i��>��2M���
���=�z����}hE4������Sj����l�U��򂕥^]����+�gj<��5D@o3��1�E�@ƁyD��_I��L��������up���ۡ�ܭ���aZ���^n:�Aa��l�PN�(uz?0�U<���Swj�{SԮ詖Cr�]e�7^fW��6�>v�P�/�.'ʝ����x!J� dY}El:�=
�o
6l��,x�a=����+�b���Ğp��N��O-9���zX���;�{������U���[iݐ��UV=�[Dm��K��	m���j�dAA�$Y�Y��x��X�~'���G��ᓳShO�13b<l�)�k��UyF'A\_9lR_ؑ���l��7�[���׳���i��������B|�\�.Ο��-�i��N�+�M���B�3q�ʁ�z�k�6�[𵁛�b��~�K��^����4���L��Z�3����	�������c�*m����s��=S��S/b�l���9]���9<��-�|�X����k�p�f��)E6נ��׌N�)����j9BK�az�!�b��v���W�I����Q��2uf`�˕=��S�=�@�j��N�������[����G��N��&��]!��\	q�/�Y��d-�� >գ�X����=�L�'K}�����Z%R��b����ǃ�XY����?5 �&�^~��<_��be��n���VW��v+��,�=X�ʹ���U�&|A(X@[�:�5^�xR�s9J&���r\����$R�<b�sW�;A�6q={gU�����]�}Hz���n�t,�\v�rV/��L��>DN���[�g���F�v@��r����F��t'j��R���,rKZO�R� ��V�f�k��2�Hr��(�v�����n����Z���q����1���7E$D#m�q��� [m� \@�E��,�aLa&B�q�2q�l��}9mm���TG���m	�7�N�k���N�ct5�⹖�ӻ��ǇV�(yU���7��A���1 �MM�>���Xs�W>�����ևUA��7��o۞�����dl{�sq�N[���C�Y'��M7X��5�A��e0����{��?2�`�xA����.�v�D���� �x|zwV.�%j��boݤz~w��k'�ڼQ���^���J�+�u�1���۹�Ð���H�%�����^vEoS��l܊��t�5�K\MK�4�	�9���h�`X��u@q��b�G�lz�&/ӡ��:rr������N^��ɩ�]'�������O#i&�H&�M�q��9�./֞������eNq��������S�ɑ3�Ż��>>���W��N6'>M'�q�dNv�8ٯeV�N�j�:�3�O	H�u!�\��ݞ���h��Tz�
���X���dU�u�߶�ΰ�������}��Tg�ԪWNV}z��0Ix��>��z�S%����:��eajŻ[ߵ����>d�^�LA4���?��Fs��꾡����=��e�km�(��Sܷ�����g-h��L<�V�͋���3<j^��e��ղ$p8�Ҙإ���Vsw�x��{,��7iCQ�7f, k�;8�CwM�3h������%����͇3����>��m�49�?� sy��Ÿ�H�m�.(���m��� "
H���>u������p��E����A�E47�B�E���
kت�z�2�}G�{�w��"��p�q�oC2iJ���^�l�� ظ�F������^_`S�s��_�c�޽���"�m���w䁮]��h+iz/ˣ���f��i	��ކ�����l	�l����Q[��w�����[�?��QM����!�5(2Fm��"���mឮ��w�C7�us��u���(�����o,� \�5��������6	���,��<v�m,M5 �����qi���u^��0.|�+W�����ѝǧm��[NP���sZs)�!j�K3pÓ�eW�	d</�x��_�]r}�䠴4:b�+''�����[�ے\����^�r�+�3?Gs�}�`|r-��c{�����$C��Z���9$��>+c�b�ؿ4����m�%~c"�z�P�9�/O���3 @���[)���-�b[(��/��{���cb��h��Io&%�/Cq���O#h#5^1n�� ��q�����ђ�L�8����ڂ���CrS�kƪk��i��B�S��w�4�GuϡO�{�_	:�6t�O�������|(iT.��8�]�8����z1��'cwp��*�0�<2�q��wB&gG�%�f,)��ͻ]�o��C�X����]]�7�h���,�T�*4DW��^8&�q��va�Xr�a箧��M+W�z�Xoo��]8��
��Y��;b�V��t���6|8�a���vT�Dd��5�����}��5������[[�sj�2�L�
�	Q��wn�w�����gp[�q}ctv��sD��U2�[@���+�*�3���m�r^���-3�^�b�-G��>�ap�����䣧6�!{�U��N�ї�9�����J�M5��e>l��l��\d󥱆�_n�vY��9�nö	(����M}��x�r��}0�gS�閣:g�
��u>s<X�	�wx__W���uΧ�/F�0��ƪj*�p���YCU�7���{%����{Z�ד��
�R�Vc˺�f�ql��t���ox(�4J��lT�Y���d��ξ�ͻ�+z�0�[��7��0JzYX��̜��-{����ܴwia�Guth�Z]f9e#��ZPۆ�Z6�E(I���v�T�5�	�.&IP��5v.���`�#Y"22�$��E[L��D��VeM�D�J�����n�.}�̫΢^��T�$͹J������u}2��N��їь��Dʇ�Q_SO�9�ܴ5�Wk�6��}�%��:��-��k���~A���;)k+V��ƣ���&juy����\���{�w��Pb1s˚��n��x�*����-�fJ<j4]L�OwW8�Y�Om�����z�eB[y Ƅ��oe�y�X�	*-�z��vTv��\A3+m7�m�<�U�����j}o&�[O����"��bn�=����{=S^�/i��;������r�uɍh�3N��N�K8����J�E��N=G������9S/jÍf��>k���,\�eW�r��E^�R����j'Qh�}�CV��y޶��!Y�������\[��Q�4"�`d*������w<՛��Dxa��v�z]$�N�zsl��85nA���&v��R�_kKfX�z΋��\n_�⭕%�2~�/I�������\�ԱRT���ᵹ�y�w�,�ݡf٫�V�F����j��*�ű����kN2�T��`����Rs��n��%H�ܫ�C)�4�d��L�����v���Zt���Uu��*^wu�E�]�_bMd9�5֗���C��vDI_��;��p};�.#�����������褍���ۯ��u���ޞ���<x��FHIB@�6���E�Q������Ky��ªQP�Qa��HD�6��뮺�뮴뮽<{zzzx��ǀÎ�ڵ�98��~l<��������y�I��u�]{u�Zu�^�=�==<x������
��]��Yt���(��[k�,�K�Ӯ=:뮽:�:�Oޞ��<x��![d,*��W�L�.����n�����:��+����v�'͇��W�(��(�|�qIm���r��6n�+2+n�G9�r�Qw�o�������tr_m����Ye�\TU��8��ࠂ����AK�\��u�幗Y�k�ŝ�vۭI��ʊB�:��J:
.:�|}���㯧a  ޠ:���r�N�`���0|���=�֞i^M�̓3\z��Q��w���ۼ�����ڍ����WTx�ln����l@��mV�(  �;�������W�UUK�E����CK��=1�=��=�\���[N\�?uz.�0�	\��s�uv�����uT/C;o��
b��	`!�{}+:��X˸<�#E����O��-��.���{��
#֯x�i�K� �|�������j1�ӗ��	��ϴ�T3��w�oɛ�t�� ��Ti}�:h^���E�|%�^���(8�u��Sꙑ,�˫'�Y���XW�3���s��3|�34�`O�ד�e#`'x&�~`�)���&�ɫ�<n���C���3W
3��6!�&(�^���D�h����t�O��ߍ���L=�sxh�f�ff�y�v��%�E;>��BB�
�cug|����Ƨ3�h+lZog��u���짆\/=!�����?s"���f�ڙ�X�3�ꐄ��3�\F���E�g	܎���vJ�
U�=�v��1���A�^�Fd�x����M#�l�F�)_+����֪FW8��b�g�b��lS<{�k�C�/<����]�E�]����|�ٖ��WJ�^}��~3[P{ҩw#Y����|���`��.�h��m�6S�=.�&)5[��f}wZVQ�Nj%�\�
�[�*7'Z�{��cC}�W���s"+P�}�K╋ԋ��h7�c���xx���R��m��-@���m�m�B��H ��������ι���?�����;��ٽ�b�F��jFb�j�3)YE�IL>!��҆{����F�ZNp�ç��k}�v�{(Ik��O?O=#�}��W�fb��+�JҸ�/u���~�~�V���2�}Ƴ�!�5��'���99��Ǟƨ����7����_+�,��������5�5�K�Y�������nj�/��j"��7C#o��B8�*h��<=ۖ���*/��á�����l��q"�j~�&��ph�dj�US�����\�Ö<�Z : >ߨ<���G�}�Ai�{�T���^E��u�aA�5��hᚶL�{�5�hwP%�p[Sӽ�u0�<{�Cp��ھ�M���Ǘ�3���4\@��cvi��n���:�~����Z2]
��~�*ny��~S{�(���8��!#�,n��9�Pγ�:ԧ��gI�Ѕ32�8`c��[����JOrY<�%���E���m�B#�`�b���Q\f�zܠ7k�����N*�{�^ۖ�ZD�,�b.�Ŝ�L5���_��o�����'�*�w2�UPz��Ǜ9j��W}!L/���
>�{��-WF
h�|��'�w�G3�̎޸xU�똩/4;�������>�cO��m��m��-����H ��N��~B����٤�0]�W�I�v��ݕ���c�i����,��c�j�T{���U�������m��:<���~M.��3	u
㯦b��'����`M0v��Eԩ|:�>*n<������ｫL��@�m}�8W��z�!����b^��_�}y���E�;Ob�E"��e?�j�a#�H�CT���].�61B����!j��}Ck�_��s9��ȼ(�8f�~��(���X�d��{�g�J�y������4���מg�����<�n�X�Uĳ̆��J#�*=Sql0��+�k�$U�Z��:F-�׻u�z������*f;1��ڷ����@փ��3^{"��Y^y�9#v-{\�zߢzD��]w_��S���L?Ƞa�(�ʗW_/^y��Us���A���;>>�/�uH��Y-NB�� 
�[�L��XrSQ�s�Cb�������0?z	�օŜ��\C�o�C;�����x�����U�A�/�]��j�1�澹�LPVC3*xz1��!���w�}�D��� w��b��
�N��;�L;�ֽ56�O�(�s���=ߔ��Q��d.x,3� ο���쮶���qR��E��Q��X��,�&�Xj��\�K��_o<V���߈��;��4��> �4�(���zo�q�quy��y�|ЬE�I��tG��ktٮ�:����ʹ㾨�B���5b<����ඟ��pV6�e�X�m��m�!p+�P7�w���ߞ��  H+������NO�m��>��-գ��IⲈ��������Oj-L��. n�wlȒ怘������8��O=uW�Ҽ���I����io{��ӻ��&����>�A\�o���f����r�6��՞뉖:���5��}�S� FY� ��7��}���jj��x�/t?�Lh}��r�1��:��ޗ��}��y�5��L;��WRc�����E�B���h�0�~��������)����Ɠ���Q�#��Y={L"�}�$=����W���/�-����!짵�~���d���ڼ�������� �k=м��AL3G��W=kͼ!�̾k�d:]ٶ�H��}!�v~�t�b� 05}��ք �ܔ�2}c&�>���C�:��ֹ��e��^8���[��ڢ)ۇ�`L�`��M;|�X6�0ui����/���۵�����Mq�d���������}���,�z���]/�E�u;,��[Y��s����oC�jc=��D3YWrh�	�}�K���Ĭf§篗T̨�Aނ���c��A��k�nE���l�����8x.�.��>]��X�4�n�іo�Z�]��wV����η�]�Gd�/r>?[B�m�.m���X�m��a$A�C�5(�K�ͼ43�SfdN|'i0���mkZ^�m<�[�<h�os�bW���n�7�;�\�C�q&���l���%�YX\�s�w8���7�;��?��E�7s��:tk����J7��r�4�@�Q�1��Es�% �1|w�� 1����Q���?ȑ��|�t���y�Y�hX?��l� ��ʉ�n;�Z���<G�u�����̅��{|IxO�8|�0����==�R%Vc
�ӓ�����C�.�2�<�������Z�)�Å<;��1����t�!��Y�7��^�OA��ZG��T����n)v��ˎ~��OSmq����L�,�@���]!�>~;\��������ׄø�}����8&�9���{q�V�/}��I��PX%O�>Vvw¸����s�}�����|ݼ��v2$C�_���[�/�F������Z��m�07��'��#`38Р8��mعiӝ�ra�뫛�A�}���'�
���sʷY�/���1h��(�"���k����M3�&�{�+��Vlr'�g����nꈃ7�	�
f2-u>��j��B�Ik��K�GQ��=��= tw+��7��y�^�
�ǩ�SY�q�}�{*U��˲�Xކ�j�kk#�H�t���{F^���yߝ��_"���څ��h�m���h��D�=�Ϲ����q��_��v]����dS�gﯙ	
�)��7W|��*�"�qɥ&�7r+8�����n�,�-C�=�@����<bK��fb� ������Y>��syq��{�ƅՑmŽ�j��U&��|<�����IyǦ���MP�a��{�+�>Y�PQ+0��Lv�cr�zǬ���85)��>�n �gf D��Mm�)���r�I�Arn�Í\vC�^Ol�-���wD
�nHLhYo�	d�S� f=�*�85��������u��
�E�dS�K�||C���pE���t�n���X̓;�^/l��\m�ʒ�q6iS
'ůx!E���,���@u���ϓ�m�c�~� _������%eiJ곚L����}tル�/��2G@Ɉ��z��o��dY~h���E�f^�qQ,�SF��?Y�g&]�[@�A�MC��:�V]>5�������}o�+2���.�p�c��Λp3^��x?s�T;g�����at{��YNg��_��Ey[�_38��#Lp�c�re�F��F㟻6���啱�7b�_��˭��fK$Wm7�9�~�C�z��z�aqX�n��.�������l4�:mv`�M����#�>��)wL������6�:���s�O�k��e�� [m��#m����j	�����ϞO��|1vwu�%�Nor�φ0���#a�m�t�kv����K-L�O!:T��(:ͥa-紆~���=�V�C��4;��� G��۹�C��^on�r����qŇhv�]1 7(o@����/z;���I�:�EVŰ��5t�;�=����.!� ۮ�ż顙����2~����:J=�_�X��<R����᪄�Ufg6��Ha=���{�9�܆�k�5TG� �' F���0kǥ�C�s�k��.�=�U;�<�T�UΕR�N{��Ƙ>����(|�'����B9�+��q��r�F�̮I��gMp�?�yC4��`o@����c�?Q"`�G�5���r*�_E��9U)蛶���̽îdDўa;�#��+�T��SS�E�(
�/�0|:T?C�<>-=�ܣԖ��㯽1�ǚzh k̪�<�>A���&В4�\c���;+IΓF����;��}�8s����J��9hw����$�IZ�������ʱ���]�ݖ���x�';���D��p�Or�@�/�<�a�耓��0�XP`ؙ4�1��)�tK\�P;<����5���lε�)��2���D��]j��3�s+��N���=*�ӗ� I�%�v�k��9Xx��dvS��R�ހ�׽�	����{������ K����=��﮳��� ǧ�h[m���m�m�أqd|��o���=���?~��&�i�VW��i1����]G�+藦�Θ��	5nqaS�S�M����ǤS����c���.h���ڣ�C���5�v�P����G��Y�S�"wn�x�)���[O1�]�)��u
3�KvC�����w|;���_9g�z�s�=�#�����$�(��à#���Fב�a$�s"-�%�_;��`��-Ví���0�}eO	�/�L�����'<��[����cb�J,[e��z*�!�tU�Y<��8.�`���75�Y"3��C�1_M5]����[̀o�Xs�������;E>ԼK4D��vE�x~'����1�G��?/|��rr�b~9��6�>���R�Y�VɆ_��߹޷��ms�!ޢt(�C���>Ւ����������)�����Q#����:�a]�m�ZS��MA���*�b��.�>�&����t�u�?�T�+F�]o&�Mg�Cc���7bS�wn?|���Ϊ -� �1�8�?��y��?%��.�$ڠVG4��uw�-Ώ��1^�ࢲ"��J�V��qY�^ �z^������Y�(�i�[b�F�S�����������+�@-� 9�՚�Q֮�y�/ kY�:��1}����L��ם���{�rb.K�覆����m���ڰ��լ���0����]kf�a���whzO�=5����S��o+�|ǁ��N�3˥�{�趲!�y���
�Ԍ�����8((?��x{7�Z�m��V-g����H�`�l�0~�y��M}qkhO\���������;c���^4l_Z�/nH��M���zR���~õ����>��c����+��]��V %��	������h"��3N���~�,ḆL�鳅�B��
S
m�j5"���:oP�R.��N�u��������h��1j݈�=�����v�Os�0d`q��3��m��ŭ�1H��;Żs}�m���5Z���h�8� �O���~U�w�:�ٍW�L�����<��^��9L'�	��D@A��<�?O��%�&9���U��yGk	�^��j��%7 a�Z��-�������	C��3����!��v���?O[�+4�~��}���{�_Z����(�Ӄ���Y�s3�ȟ&�}Ʊ@d!��siz�����S����o�S�u�2��QҺ��bx�{�D'��
ʎr����n������y���]X��0�(��.W`�S�9�6�`�ҥ���k*Tw/N�'�Ɇ�VM�*p�p>ã��V=���]UUQ���?[Km��m��������S']�r���? ��2����Η�%��k���O2I����=*<����օ��@�۳��UGy�����.z�'�C�	��P/ld��ǃ;:�\�H�YT�[ۮ�Xm�������_��ڮjS�T��+�Γ�K�J��5A��4�W����;�-/u.+���w�A����R�Z&��F36`����^�0����-�8ܤ�ih穫��4c�%�<�;�#`G��R_qD���d}��Â�)��7^�� ��lJ�eK�b�3I���E7	�9jus��$����[��2��v��_r�m��n~���{״�d��[��Nx��c�>}K)i��VDu�E1��yĄ���A�ϫ_����`C.��Mt�Tc�i�	�u���F04�4�]d��
�u�a.����E?,�c�����N�y̘����	�
O���k'τ@���E�B�ߥ,�H�c�4���{gi8��iVV�g�����[]z/������4rњ#Zwby�t&o73�S>j��k��| �;��}���Q]����ݝ3':w��I���V�Ź
�sj�Ly��u\	TY݀���.�]�Jӧ��m�y���j�D���[N�Z�������ݼj��:��D���/�V�����U���a_W6�wc}b���m�:�:�͑���h�y�M.uʥ_;xi�}ݡ�kh���n���ؗ�:�f�&�����V�
��lM��7�ۤM[�f��Xw��,��a�J��7li���5b�ì܅��[��qA1R50 U�Im�e�[!D:��;����لm^7�&�B�
���K�7e3(�f��U���Sf�WLC��5�%wbgSq��=����E��Yr۵WB��?�-�s{Ŋ?l't����Vņ��'��k��
�ۡe�T�f�#vh�>�J���g2ìuЕ�zy�X�T�l�x�b�b��o+n��v��m�pn�����k���le��<�u�e���'I��W?`��]bEwO�-Sv�RO/�[�8 ���Q��FhEm1��vI�����;E��wq�fX?_�+RY��\u�4§Uq�[6���=KFWt	r��{t���]�p3�b���𻃨����n`�vKq����G�"K���vu� d�[��W���eu7p˪�Ɯ��镞7��Rr���ZUY�K�T	^R�rZOB�v��M���
�ڭ,Y��eӰ{�Y��vF
! ��I�|g��:wl�k��Ϥ���g\Igא��@��W֦*�YX�w��&��̝�gu'2������.�_`-�#Ȼ+���s�;N��}�5��Z�����;�E�0�c��[u[ڋ{z ˽��o]kΡt��*��V+����vU�}N�L�d��ΏK�ghS�&ĥ����	+��G�Śe<ʛ�ٶS9LcaA��-Zo��ˊ�a]�҉�n��\I�!�eP�㭛K�4$���[�����G�|�S/��]�	���<�+S�Lv�lWc�6#3qwK�у�]���vc���<�Aٶ����M����@Ѱu�A�y0Tfp���]Z;�k��[�m���dK��Q����DWh֩�u0
iX�VN�V�q˳�9�O9�X�_,�/��gY��er��ۉ���*�m�%a��56F��	�����C���͕h�$;㌝�3Iۏ�UU\}l/�o(zfqړ�d�9��J�>Sc�ք�0a�̔y�K�Hs�ޒP��]�)��YQ�Q�Wo�
��T-hQ�)qnƼ�����\��Eެ��i�9.v���&�<��r%P�=.`����1WvS=s1g[�!�s�٤�sYz�w �:��u�[�^���o�y��׷�K�$jUEI�DZ�$
�I�q��F�{z|{}}u��]i�]z~��==<x���Ӕ��n�q�wyG��qt��}@�B�$`��1�\{u�]zu�Zu�^��===<x���x��R���滼�⋎�����������ۯ��:뮶�OOޞ�w�~��~�+�t�&QYV]ǝ�GQ�U罻��.���c���N�뭺���Ƿ���<t��t�TI	�E�}����w�wvu�g�GRw��;�ee]fq6�s�����e}�ϧ_q��K��Y�eSj������Ӯ�*��(��=���>2H�#.��p$)P�RG#YBH{׶����H5���,��{[��w�,���w��\s�������O
�e�ĳ��$Z�B�QD�bA	)2Am5	��TpE�����n��$0�<E�P��`��D1�9-��#$�w�݅��]o����4�]�d3nq�Pm��!��0�ȟ.��P+)m���'I�S�]��� R'	;Ģ�2%Q��a�	r4���)+�q68[jH�r�

SI��d�	�A�H&%��P��'�1l)NEN:��0g$&D\]Q5T	2�)�qX-I��"�q �B�� q���dq�6�m�m��[m��	$���]���8�5���8e�prҴ_r�bb�\�/C�H�v{�Ďnn=���:E���d��RN�/R@���_(1��	������z`s@��D�y�G'^X�2�z)���c���vk�|�����+��t��H5��7�,ƺ�\2z��->����T!B��ͱ��e՝�=U=Z����m�*B�nYy�6�Q|����!������>�zw%è+�ԳM.%����������.ú9��&yǥ!�����X!�)��Nϫ8��_GQ4Lޜv�J_�w��[HL���e�dkt�H%��ZBg�x܀�:5�4խ����Ռ;�8=�T&_�g��kBs;������V+��A�Nצ"��Q��{v�=���opp��� О��^z_'�Z�7�>�k��y���w��؞����ȉs�u,�����'Q��OA���38A@~��[�B#��&�?|�
O�����S7 4���/�`�YD�AC�����s���s�s� �[��t��
�x���E��/�>��>�V��/ZO:���5Gc��y�t�,�
�hia��v�9JA���C_E��{���:�^�̬��UZ�ֵyIЗ�u�bѕ[��dի��t���K��\j]�����:=��"r8;Y5x�5��1�j:�iK\U0��kxmN	����go)�����"��y֤"�S[���z{~��m��m�m�cy��������'��=Nȉ��;�cჿBB㬓�C�Zfc��X}0h�Yc��]��%�L�y�3�,Lz�8���Z�C��ɝ#�X�Z����5!��%�L��9�Q��p�8;p�|��J����!��y��w+A�½���R�`T�Ms��E�����W�IګH�h���#9�#�I��#k�юC܂�<�?b���C��
Ms��S*�w�W��ڃ���'�yy�+I��y?���C�;2�{�GX� ���]go=�ǜ���o�l�����s�:��ay�z4����X�@��4������}ܬR�I��C�5�|�)��C��"��U��I�j	F*�y�H�k�8qã�o��Q�R��5�0��8[��*f����-Ml���ϫ���3a���S�10�"�S�{3��}�z�������^�3s�LKm���i��1���{���!ف}Kg]����
,L�N�z_�v�:�/Ai���Kul�/p�o��w#��<�;�j�j�d�mz�Е��3�w�l��(4�r���U�i��W���I�֩�s=�1�uu7Fx�����Oy�˴�I�;3#7biŽӬ�7���R.��&(mY��VR{*���ud�����v�;���w��q�@<||A��m���m����d��Ϟ|�}���6O��-���wP� � ��q�oR'�<絁���^A^+�e�/��:oy��Vg:�7��O���)�δ����}� l�Wx:��k��
^Y����sO�r�p��g,^?��9�i�D�
\���7�� �P!�B�|H�z<����bz]v�զy��Wu�Ľ��c�C��ǫ�V�Is�ׇd�;0�pw�5x��N�A��cߙ4_������WM����}��d�b�z��T��I�� �`�떰���ܧ_!���)�^��͡>�O�`�bx+"ջ)=�[�U�h�8���Ì��c�v��9T�](��pn��i�)��=��z�p�>��R[�4f��J겴ӷ�ܽ�j��p����o�0�֐���b���n	��xN0C�y���t:E�k��ƞ،̣9Z�"&��뤃�|��_��W�_��}s���yi��ɀ��4�jR<��� �boO���l}�UW���M�O�N��)���Y���Vx�j롵���������Pه�]�TG�>M<?4�_�d3�,�,�"�U&�,
�y{+`�e.���ܸoz)ʺ�@�e��oF.��Av���7ԅPr�c��*����
��,޿��V�N�h�s�#s�3�\�u�*{��҂��dlxY�,�z�J��Fk�+�{}��ת�m���lm��R␉9�w���:�H������@xO�vO5�<v��3r�2+��w7�P�n�;���kb!�$JU٥LtH2�p�c�6��0�����s���1M���z<9��;���3���o/o��1S���I~0�Kd2X�H�C�|/��D�9�*c��$���U�Gu蚢�;�)���I�ĳ���{}L��;�8ʀ$:�q��sl�yy�/���J�`��j�+y��0��\oj4�v-Ժ޵��>1k��O ���Π����_���A��$2 �Y�3�ڻ�Ek9.0����I�TW��Q96�{b\0�fh�h��'v;{��߯:��Q��}��0��4N��O�-7�#h��'���'i*�� C_�I4˺rc��E�٩���������AKր������M׳��1��T7Y0�!(7Ǚ�G=�-mY�z�9��E1EZ��$���B�P���N����%�=G�Z$e�%뛬޲Vڐ�۹�?n����s�O��0���Ջ�"�6�
�����~S�KP�O֠��}�����E�����Q�xYv��^�Z&J�dW�S�6:���y��Ru5[V��<%*]�pWk����B<!��z�hc��"B��l�D���T]�"���vuU��E^����}l���v���=�w�ފ�����i[cm�[m��#m�`H$�)�9S_���W?{&FЩ͌%��h�zr����
um�%�wN���rn�X$��5Q�+=�~B|�ӛ����Uq��S�,!x;���t�����|�Ⱥ�
����*���y�S ��_�/nGY�n���g�eF2�g����������vd���X��Fs�=ڪ<}����Tx��ё*}
���c1���D�����Χ��oS&���k�DS� ���,#ZwbS��0������K^�UC�]s��n6X_Yt5񝤾;�%ȅ��ueG�,|���肘L���m�ɑ�P��6ߞB�=uW�\f���[\=���2#�����H3����=̊�X�~4$_|�fL7n�"(?]2�nZ6}͏l4�&�g�F����Ǹ�����Y`o�HAGCH.Z�ɵ�4��sj�{zg��IO,֞7����<���OW��<֚��Fsc��k`�غ����eb��٦ط����������c��0'3��]z�#[��A.G��0|T��u0�  �W���� �,�7�74v�H�;�`�~���Qf�H!���;�OyX������!�t.�����`���%�={�p�G���)J�LR��3)0�cb���(��y~+8wow���:︭A�d��"���������ſ|����_�{˫n�7;.D	���@m��m�t91�B����9�ݨm.����}�~�m��m��m��p$a=�)զz�O�T�@A������!ٲވ,�:a�Y�ZS��Ov��5GwάUz㵻3$O�T�i�+P��9����^�싇gk��O�T��.]�ȥ���
ǯp��=�y�߳�\���3`jqYiW��,�k�X�%�[�(�ܙ�T3x���D�v��I����,�r�o]T[��ؖ|�8\&��7��#��JWY�Lu�"�*�#����F��P?�$���_*�T���
���]E�f}2��owX�}��V���.|��~���+�ɠ�ي`��$M���q9��L[<s�l�>?o>�>��J�8���y������Xg'{E(�	UϜr|�GO��;Y�D�WN�㝁�b�c�3�F�wɆb�s�j�Zz��M�|���-�>���Ց����1������o�%Y�����(���P�^{ks}ǅ�F�adhN.�1�#Ր4nn�!���P��0~�owE2�����].�	�?r�kk��%d\�t c�����R*��3��j��i�A��șTc�����!��~Z�ﾕ�e9�폨�!hilɺ�ҭR4��X	�����`����UF�{�����*@�hZ�J(B������Ws���{$ތ�a�wMM��(��j�S�Ag�7+ �_���]��e��e��m�E<��������^�UT&r����,�.>9�I>:�b�1�]]Ԙ�%�����m��]�i��mnv0+�a����0!=s��[��O	=���ct��z��a8�����KE�k��^~����Iw�C�e�R\=�0�Ŵ��5�G�W������O�{)b��w�f�LY�W�@�Z<�����
x�t����-;���w�N�u
ϷbUJ�cϜ���a���N��>{�3�\�-�Ϲ8�2���Q����ƹ>��ٕ{h�B��z�~ot|���y�Z���}D/�x	,��k��6";Ŭ?s����C�ٳ8��L5ӝ�z��^j��/}�#m�8�/�L	��4����O��a��X$��?+�'��3^Wfiì蘝/�01�����@>=y��Nn��ྖ])WT'M�d��vf諙���$��;�wI����4	m�8"b	򙗶�������ȃ���8��Cg���`��${�0�+���vߴկZ��yq�l1���|+�Ykϙ!r�����<���+����i�:��čw�X�%d�6<��ԖsL|�τ���v��ܷ3w�r����}Z��2�h��x�u��@��ILc��	�!��W\��S��Ι�}n�1���f�Q�/��w�r��Ht�Ia���r{{��w���f�������[m���m��DiOV�eB���ղ%��yȸ���~㶦
b����v� ��>�ⷹ��x�/��܏^y�t(�Ԝ��(Pq�\�C�qN�����4		�ŗ�|�}��	���vn�:A$D6[�~hO���nE��(ʤ�98hm;jR���x�_z}�H�'����=��V���^�w�nCTkb�c��a�beB\��<t�?��6�0�Ȇ�kO�I-��m�=k��|}��!�\|xz�����|bܥ�����+�̶wM��)�wWJ�qD�uK����ү�"HQ�"1w70[�2w�{*=y(����zK�e&{�{z+
 ��H%��{�k�U�(�`ha�����88֋L �o;�:m��g��9��'0h��&���OL����7<���>����|Bs�$�|e�h��!�C��Y�{�w�y�su���G���1�P�TXPY�����`��>�:n�4(�=lO�A�L =<���ӝt�{Z��5���,��O��'g��wBOm~���l��w��kC�+����,�w�\�����~����J�^m�]�K�UU�m d���`�n�pf��e0��#ޠ,Vw�� u}_N!��^���b�������I�U���3�}�>�ˏʆ\����rZ7�J7W�T��i�r6�v�M4�dϒoc+�z�����F[Fj���{�o���	4�Qi��C�Xt��-��cK*�n]��3��K�
�!I��G�O���L=C�uϪS���[b�ؽJ�ՋG��3W����%��t1lj��K{7Ez�⤁>�kഊ�M宴O��.qp ����
]sUn�~�;F����S�����7��b�
3�F4����V-k�O+"�;>��BEU���F/i��񠩮�e��U�v�pDZ��2hc	$3�����ޠ�{�"�zk�4b]�T6��k[��3��ɸC�:�������#�S�7n�����YT/I�DA�K�c�s0}��}y+Q���~�2EH���Z�#CMmH4L�4u�b��UY�/AW�e^W��.<����$xC�x.a���gޙ\�_�9*F�m�dJs)�����{t���ljFy�"�iSR�����GE��q-r")��}o��9k݉N�غ���(cL5"_{�b9�[3,�>z�_b�x[|�"��`!e�|}���꣢���;<����Һ)|���d���k������aO�E�]Ds��n��e#s��q%��� ������=��S��ZQr���U�����:z�+?:�d�g~���ڟmoh�Dϕ�K�%/C��Q��/Z]0o��x��H��{�|PC�H���=�/�,o����,����J�3}Gd�c�04�k���B�ܮ�r�������/=am��m��\H�m��$����=��ê4[���Qu��Suvו��ڃ���1{��93>��D0��(bx8��U���"�Gb��Wd���>F��%�Z��ˊ��S�g�Z<v솏3�jRR*�����(꽱�?n�%3��<)�`Z�绨]��2�[����/C���'�v�}}�q��\�9�m��ϝ��.��V�y@%>"A�A.	��~��u�g�mvhv�Ӊm�-�#�+�E��P0�D	��y^1�rԯ����P��k}�yZ��v|jnԼǂ{�~�E�]>��l���5�J�F���~�#Ӛ�#��)_��~���=h�ʱ���X��	(�
�/���|�!��c���o;ü�3h4l���� `~.:-9E�VQ�VgQ��58��!��˺P��~��X*�%�9S"�j&��� 5��{�US.�Ҿ,��!��m�=���Cva=p�����x_+|���X��]����k�9s�Q�;#�!4���@����p�q|��^�Au=�Q��ǽ��K��[#�#��������.jI�i��,��"-�tE'��OX���:�4$`��X�<� �侨�ѷ+}�o�s:�6N�t"�oLX0����\�ǖ��md��A��w�����! �gbEw�L{�眆�KV^�@���8do{b��Y���E�����m#�&���r�Xvj�]68rgz���1�bb/.��O[�����I��Xf֛]���B��Ԙ��@/;gLt�����+74W]7����Ϊ|AN���V�ʈ�Pt�E3D�Q���fJ}��uf��:$ed�-�zZB_>��f��F�Vk�%I�2���}���1����S�3t��`�����CT������_nޫ���w��È�Z4�Tw2��Y�.�ɛ����ꁾ� M���K�!N.�ɔ�ky��ƻ����\��b�6ׅ��b�݊��V�x�#���ƞf���#����Ö��7v����w�y�*1d��n)tk��a2�ֺ=�U�
ktm�Ya4#A�Sr�ܙ�T�5��+6��j�GL�\x�Uvy���nble�\��]Z5�u�Y�tƸ2���G�C[�J��f����v��Po-��y3����كn�v>��!.6S��wɚ���:�S_7C��'�T�3j��~���>n-j$P�]q�}�@�Z����c�s�n�n�# g�Z�c�Z���I��r6�״����i�c�\�V�^�����캽�ֹ@��p��b����%�q�Nc�W�2ťhuv��)�x�N��Q����&q��|1�ICa�d7����v�t+�X��n�a���+g�"���I��w9�CU����Y�1�{�rec�z�����n�
���J��o�&���{C�6����)L���Y�g�*����}d���ܺ�Z�l!����4V�yj��S�eN�r�u��Ypt;��\��V�U}�y/9��b���v�tm�wp@�5�/y^��sh6+�WlNt�������]��]Z=���)WV#-��6�Lڷ8z�bJ�М؏Q��;�����wy�Wsn^�����VG:V��`Θ���=�l#�9G9VZ�Wb�GBy-j�es���P�UI���Rķ��!$@Q������Q���P�a��s}F��|!}��;ʦ�-*�VH�1��6���Q�Ǖ��O"���&���f�S�q^t����0J���2�3N�%�VӂP���ݶ�,���4��OSǒ�U��gdP�������:�!��i����r�̝�j�n��;������Ժ�����X����W�V�fӬ����D����Y �Ixi�BD�j.�J\q^|r\�ƛzzu׎�뮺ۮ�==<zzx���x�$%yvH,�ʏ!r�;.�uY�; ˹�ݏޞ�u�u�[uק���OO<o����zZGGgg\]~�)2#��J���-�����뮺㮺�n��������Ǐ��$R�r7UYbE�u`gVڱ��wtA�Li���:뮸뮺뎽==<{zx���H�$���/�d�;.��dw��O�|߯��n#β���;�ʏ��'�>+Om������Ys�/�K���_;���9;���u������k�n���f/�{l�Ӵ�^{n���璘�;���g���m�>|����3��|�u�f�)�Xs}{>|��/���I�t��d�����k#�Yu'm��1�vGb"�$�QH� YBz7tf���M�<�>��-d�e�+y�e�h���ׅ"��@�����P�"=�}���v��i����n�m��{�y���qZ�����F3���w��Ŵ�I=�DxC�v����8���I� Ƨ�(2h0|]�DI�ۃ?&Ĥ��=5^c�7����|�x�+����bа� D^}�9�1�9�nx<(l�k�.w�0�|e��U?utט
��rcX����=��.+ݞ�N2�9��e�$q�N*�.�(���η�]��$�Y]B�k���eo0�d�q;��h�P|����pl-WՅj9S0������K��'
9(w0��dWWu&�2�O/�@^h����g,�b����g��8t?�G���G

Bd\Ǯr�-�rt��������k�;��4F,���&����µ�9���������R��\��lg�������<}2��fz�E=�����Z�k����dC���!t����$����<��U�*��hY7���fn 0�vˎ)O��ʦX봃xC@��}�'�ߔh�_�+�Y}s<ɷ
̺�x"D�xT��1�HǤ����m�=��� � ߸W���5��dA~F�:k�I�A!��&�'���ʵ5���r�cu��;<��!uj�~@|��B��j�z�����>�u�ëq��W��Y�;��B���Z��<�^<c{��&�ز�S�;�i��-��
i�m�˕9ɵ����<��G���Y�?!�"�Tz~uj��p�>�0� v�%�k&A=�צv���:��ח7�V��㝝����\���C$6<]��
ډ/Za�4��<pAn��q<4��\Q��U�.�+�W�I�Bd��o�_#������u"����e��K�E�OD7�����\��z�*��M�� z���uny��	��b?���g�}�-rR���B���4�ޱ,��:/;	����dH���/&ϫg ��T4�m���,y#T��M3j�O��-��ě����,��CRx�&�	�z
?���C�p�`p�>��!�Ǫ�]t�ǽ�#%�b˻�&O�5���r+��#r9���ǘ	DR�E�n�f�ƥ���'�}����S�z{�wV0���F�y��Q��Å�h��m�m�CM�\�/W0��Ss��8�ܳ0`�C��<��ޘu-�4_�7'�D�'Ӽް��OB�{������T��R��e����[4�|��~{��f�xa�
�A���ex��c�|F�]l�.=�/G|nòz��G]��:���gn�1`[w�5�wL	Q��G0ec��^�������m���Yr�d��ށB#td�9J�5޾]�a�W*+b>"�T��U)q��Yk������<�޻ҳz�$�oo֚i��m��n�"7�_���z�k�����P̉��q����Z��f��g����W��rcb�� ��]\��'2��#$��#�q}���~t=>S��u�D.�E�,��Ҙ��|��=_5K�}�f�Ǔs����k���~�L�S#g�Hk�[��P�B�~CL7[�/�L��!��|o�����`���\N����{�k���a!=��<^���ހO�b�j�O��&����v׹0a5Ǧ�5g�����V��S��s޲	3�ߩ�	���4�gz_���|[wVF�J��ݛ�
 q"�ZD3?k�;����9��H�����EC���Y��c*q=kQ��t��RzC�a1A���Z�D��\{Ʋ�z]�C:�6�����zXT�'m���hq�`QE��M/C������*+>��4i��9��a`��~*Gm�/M�W�6s�ߴ:0jt����tD�:��߼�z�����WU����k��m� ����w8��Ȗ�bh��#ES��t��5��g��Hhwkݛ�v_���w7H���W�ؙ�|������X��We���8��f�0�oN�x5BYSo�*�d�~�u�;>a�o��q5�����t���ok��E��t,�o:���K��&����)�,�@�^�G�F�fm��PI��P�[@_��c�ˁ�j��@n���s��,�fa���r.m��/�;����}~��4�m��M6߽y����z���tyt�hNE<���s�g9�9��{�H����L�0	]%r1�߃�!�_�;��Δ�-��@��6b�0���@F}��h��[͑�s�<���(S����H؇�xf�`k�P+�Nb��e���'������u��нQ�ۍ�~J8�Y�>s�Z�[���G�]�6�{���y��P����x���z.�5�M���1g{e�<4�k�y�L�j�0��bފn��P4�㦧p��{�l��kE�L�<��3���|_\��p9��H�B�S�O���/��tz#�T=�Ʉ5�v��Q�h�+�um�Z<���n�5��p�[�hi�dޭ����=]���'}��Y
>N�v��*��r�1��s-sbb[:/�%�}�TXH��梠��t4��UϵV�I뷣�U#���8[ ���O����S�����Y��1��s=6}ۏ|T�[���z7\3V�	h~�\k�;�^LWT������חbY�f��\Y4©a�ݍC�԰sz��)�܊tV�u^�l�c���-�����ՊuӖo~��:��D`�`c�8�L�����PA*���(+dv����ݰ��[�u�}6�9EJl9�}��rm����w���M4���n�m���tr��嚚!����>�݅`�z�kD��0oX���h�Zi1�~I>"��������P��t�:�?K�r����We�j`n���;IX:��T��Q9��wn���q����Vȁ����5���U�o_;�"��%VG��|?
Uz���ش�GA��U���L�-�π�
�xa�yV���\F����������̙����6�6���tdM8������½�"V0.	����;��(t\8[���ɭX~dx�TN2�W��ϥ�뒜`����o	�3p݁vX3?��qɊx�U�U}�L�u3�8���a�.��^P�׮1��G�Sm|O~O`����-|�[jo��V�&�u0�ߚĊ�h�Y�ؐ9��]>��\���'r.���w+'ڮ�_��  q˻�}��G�$����mA�..��)���V������*
���\7�z.�{q�P���:�y�	�'4|��͞��格���=>�/�]�n��<�6O۽�g��ޅ(�Y��(a	��ō�7|��.�*,�u�FU��Vh�֖[0����N�z
�b���������+����}V�C7�Ugkꣻ�^vj<�GR]�.�,��W��tX�z
ҺΩޢ�ѹi-�����x���?�����C�6����kܿ_���ٶYtC�VX��b��k����~ŧ��	�l��9ڇ~��d�  a����W��`��Xl�(y�<�{\ّ)�f=�F���G!���co0���+��TZ~8OOM����������/��G�\���r6o1���)i5�}��H��@��(�W���}�6�
9�S8�n�	C�f����_F`��4	[%Z�	�}Z���]s�N��@ C��]:Wﾱv\	&���`�~]pu`�i�f&I3��#����ᥙ�E{U�Q���9�3R��/4��z�݆Y-�MӨv��Em6Qaz�s�S���U��k|�{��c�U}�g�aRX"�b�u����i� oO�qq�{#��A?檍��n1�I-'���Tf_a){ف7�';�ěi;qQ^�5��
Go�Wb��]��泆J���)j������r�13Ed�kz��#8�rL��z��9���qQ2����c����L�i��0_;c3{�.6U���kut��Ҹ������{wf�y��b>{�O���v�m�6�wT>����]e�n����@�ۛ&�'r]��9>�
���s�SǶZ�+�N4�����E|����v��}3��k�+��W��ɚpv���lDf�Z�E����G�{��&;�������T���h6IO�v̰�����]�oX	t���>��a�����^�ɫ�7\tµt���4��� �O����,�?n=
�qUZ.�5=�i�e�����u�����%w<�z����d;�g#Qt�ړ�od�i� K	�^[�D�F�c0n�;��O���/����-�.��1d��Z�lg���ǣ��6(��Pﹻ��{�o��X%�-��m��������/$��U�8��`�q����:��O:��l��v�2����0�Ɵ=�j����/K3y���Ԓ����F2�\��MbVk�!UЗ�-�·|��tP��w���X6��-���k���&�!׌��x*�h��EJ�l��۝{�����\d�b
�j�R}B�о�`�4��N6�ˁ9��<�_04��]τ;Շ0+#�2t�a.��	�^.3wt�o!�<��g,$W�q�ݶ�M4�M7��\��+9�9��d�'���&����9@xT�/�~=YޱK�v���n�J|t�?�� ;�7�P�8[�Jc.c�����ݚ�zU��vm�@E�����$�C��إ�ڊ�Z���$Q��F7S�-�Ӊ��0k���~�~��3~)W�H����^M����_A�x��].���E���Y��2o�@�����<m?1qP�!!��5�n�� ?������C���|�3�΁X���E�J�PqD�X��`40޲h��(��g6"��f<�Q�>�g�{j��/�T��+p;.�F\Xz�����w��u�ݾ�5��Ԓ]Nn{.:�q���V���Cێ�#��Φ{ǅf��V���;��6d2gW�"��`�Μ�G;0(5z�?,,�x���]�}ƽ=��?��g9���`5o��5xO䷘��Ck5�g;���t�M=����<�V�7o�����ư�+:�9���޴�J˗p� R�gr8D����Qc{R��u���Y�N��N�[��4e��Δ)��4�M4�M?os�2sy����}
=���w<���_D��o=�4�7tb�rFe�]��:t�Ŭ&za�g�����.}�"9�#�=���<�Pl�[pz$�fj�����s3y=y`�\p��� T��"�)���3U��/�j�Ô鐖�j���m�zH��;��̯�i����<w7�`����UKM�Ώ\�Ω�3�;$��2ٟ���l[(�h~�D�n���X�� 32�"�;38ΖP�q�d��˘�W}gi1������Lux�z����	�o��H@�	����VfqFȖ�J�M�U���B�p�]�n%��ǊM���*�pȱ�UFFl�N7���� $�G�:���B��9@z���f����M��g���:4�(d�ߦQ5|���T*��:�X��M/c����ޔ�JM*z������=�rj}�.(sH��c ��dQ�ע��˻jX/�v���< ,�a�o[[�V^�B��7j�r��N��K�9Ӯ��K�Y�WJ[�i&XVS}F��nV��u=���M?m��i���!���3z�>P^9��$} nq��@T��F��t�9�x����J�s3��{t>�]�?���[dr�y���ï���'���5�.��~��k~}>��N�-2��p�I���ޯY�f�:b�7ǐ1��Z�l,������y�3x�����Y�Y�� A��d�$�j\э��.�cm�����z�
�w�;= �~#o�(�O��ϯ��ڷYw�lb����fE,���'�:f�e���/�`�0���tb�a�zsZMwL DGoڙ���ޒ�����j�`�y��%ס�^	��ss��\�#���CT��zu� )"j���p���F�x$�ļ��ӹ>�>��r���\m�W]� k�h���WD�M�o^�k��Ҙ�1����#����뺵����3�� �ֶ�h�m��#&�m+�sWZ��&m�ז(�a��l^ԩda\w�&�.���[h�fʇ���03/^D-:�u��.X{9�fn��L­��R�k+k�c&�7�������3����ػV�F幽��Y�{���8+#���J�����N���G�;�j�Ɨ�Y�ة`����<x�M<w��ġv5�K	\̮ٵ%�%\�!+X���ZN�Za��c��d��Ō��e�޽�3mQ6�_%ӗ1���������eeN(wM�����֚-鼰#ف>y*�!��MY��V�	!ILwv���i����},����5��jŕuc����N�oxޮ�4��i�[P��o6����H:�z��0�۫�W�9�&.=ܧ
˃/� �����&���*�SYWo��~���t��oa	L<ٺ�u\t�{\�+�o�ݴ���y`D�!X�g��gpuC���\�޺�U�ݨ�4�L�ڌ)�NK�2�oS0���Q��S��}6u�mJXQ.c�M��2,u�����2�]��ˠ��9^Wv�{3�.,<��ٯ������5�B�xF�lm�ޞ��y�]ǖ�λ/.�8����x���kH�{yQ�lrHN=����);=�K�e�6)�����S�G��9Ǘ�K��N���i	�!2�9�)Ӷ�i�d`W%�V� �)��ĂM&[An���ʎ͌!���幀.�(�O
W�N��S#�qv�p�dheQ�7��1�#��1ֻh�ܪ#�eb�f�}y�$$@f�,x:��')9ۥ�sb��L���3�ݘq�eEB���ݭ}��vك������WRJU���pEQ땗&�8�>�݃MFR�� �<��ei���[���9!/g	�X�b�S�%8,RE]-f��="���Ä6GDt��I���Y3Z�Z5��u˲L��yEf��������l[�8�Vއj(L�{x0�f�F;�քn���d���:�6�ԣ�5�^�����P�\�����;���nn�&O`�s�at��K!cJ�=f�����
��ˬVX:���_�H��8��%㫬4�9�|�0�K�f���)��Ci޻��6n��X��0bs�wk&gʽ�(s)?.�en��nb��i�u^�p^�=3�)�i�Ι�a�׆TbKB C�S�]�zےt.��E�|��q�	_�.n�*/�0�i���-Lt�6!��]�hnI�`;���U�v���X��M���h��P�,og�w:�9�v�R��(<�2R�J����Vޕ]ީ��y;�^�e���ݞ��|)\��{�mUի��r��^$���8��;f��*������=�Vu�v���o�o���뮺뎽===?^�<x�!�~�wp�
�dYdu�w�w�9Id��*��=8����]m�]u�zzzzx������$	*Q'�\���W���o����N��^z�J��8�ӯn��ۮ��:�������ǎ�I9U T��R9*H�B�AwEU7�)��c�8�׷]u�]u�\u������Ǐ99T~�<�쳳��y9ye�|x���K;�oi���]�G��>��H���^Ӌ�ky�������VvYl�ߵyiЏuR@��bHdW!WL��tIq����l����޻�;+���}=mv[M�����͗��xtu%^���^��i���ס�h�����Γmki�����/(��M[���	 di��q����¤	e�v!���I�6Z��2�E�iFr��i��fD*&��䈔	n4qae�l��)��*&��w!�D�g{��𸺒NV#�Zw������o3A:+l�O\:��]Y2�����m%�tRi"�M��	�H����b)	@�"��"JMHO,HQ�HD�Ȍ.l0#qĉ��"H��(��26���pDP ��dKh�&$��D�P`"$HB1��r�9�p��0�c��؈�`�׏��m�m��i�Ϝ��/9�/��}�u�`.j�d(�k\�$�X]v4���Y��"���ݫa��������uv�4��OR{�5�4o ���k.����g ����1g�^ث���g\��Le0�l>��2I-<E]�Ţ���^�z���B����&�K6XOy�Y=o#(*[wN		h��R5[��8�fؠ��\��'rR:�o/�Dx�����!���"=:T�m��Ǫ%��ֱu�z�	�Ď�p�R��w��מ��1�wƭ��W��%�٢��w)���d��#�����o��T{v]�Y���T����"�Qi��A��wbE��ju�[~"h�w�.��k���ݦ�Uӽ�~��$��!�z�5����jHv���B�Ϟ������zŉ��۰�J/R���ޯuv�/2��@a�\�ʾM)<
��̬��mAl)�
�$����v�81ʽ�˱�Y����R�b���*-�����cG*=�0]���of�iukv.��c�� ��L�r�&�V �z{��	�����ueo����B:��L}K�9K�K���a�	�̕g���:�h��#6F'�߽����~>>>���=��-=�l(����"�Υ��کf�z[�u/`Ker���ӏ�u\�r�a�0��a-�~,�S랏>Ώwo�7]҅5�q���{��+oh�֧�hRE#�W��b�9̀0�}����*h*����_9u�]�/7;F�������; Ϸ�@��~/æ�a�d@]*��q����1'�����c_�6t��4�_J�ox��8��&�k+�i�Huw�����-E�+�$Tk����n��puRx��ұٗx�H���MOP�y<ŝ^�>Rחb��q�y9{��Aе�t5�T!�L����_�1.4�\��RZ'�^Y��-z��P��g���`V�� ���&2�����歸���y�'n榟��
�-�Ϫ�#��w�-	Iq8���=�rnc�vpQ�U�+aG�m�+�JD~����3�����1ν@ʽ~��ZƠ!��;��X�|�e�9M!�.q
���3������K��Ra�Nُkve>P�W���kmu������Š�[m��M��9�V�+�e^�ݒ�+����#�W��װ6���V��w#�&��	�hp�������p�O�o��x%=)%�n���
����Z�,��gp~ɲ�vGOvy�A���-����r���	Qonx�A�>ђ����<�N���=ǵ>�kf�5�/x��պ��#;;;<{����*x[��ǝ�L�/��!��$��tվƱ���O�Ie�7+j�}^�������@��gv7���0�wz&
d[s�?zk�˯�FT��̿_?��a0���c/�����3���sr���#��2g��yj�	l�#3Z���qQI�&^^e�N���\�:�q����&�p��S��[#ʆ���3�_�ߤ12�Ϣ}����9��U�*����8��x�,����g�.�1���)�	�dw�̖�VQ|L��k
�(��N[�7}4D2�Q�K���up�C�Դ.wX���jY�443����ˈ ���[i���(k+��r���p�Λ�ʾ���"y�5ە��oL}I�a��q�Vp��nyמu��߯��m��nԶ�|�o��b���m6���uu[Lk���ydݶ����}Kx���Ba4;�w>�J-�*�@1 ��C��{{��P��#2:�mD�f�w�ݷ�m�����hQ�z
�=��"|�xh��7z����FI��z �oxE+$�G8���q�[�]*I6���Z,޹�+|�[�3[Wcٸ��ξS�ۛ���Fw�p�%�����ǜ[�&D�W%[��l�5+j�;���w����ݹ�!¡z�r��t����j�I�~���zZO��>��X���5m55 3V����Tx9��x����qx�l���ӭfm4Q|��Uٰ�<�\egm�O^����Pq�Ip��w�.��=����^���so^�!h�\.x���H���m�ް^wM�4�v�lAc{L�}�A��A+S�(h������N������b�\N�ac��k�d8[���a����9��<�����ta��^�^�������챚.d�dC�Ak�@�h�-nf(�Ö�۽]��$��GSV��_+��E��i�qY}���Ь|X�ʥkZs��ə��������|||\\\|��~��zo���w:0�2��g\����X���"��:u=�x�����N4�ŻԗLɒ���Y����:1$jI��};����W�ҧ�*�,��0W�te*OnV��6���>���p�37����I��w-�JL���L�3����2t�v'����2�$�ݒ�I�sȻ
e3�і�&������LI^��y�� �g歩j�v
�������E��Ś{�t�	�Y,���aK���M�������4W,��I��n؊ʎ��립�i���.OeO��}��R��\'=F�<��
��'�ogn���l<{�->m��&�"t�^0LED�TP��ӜX�q�{0�p����N7����� TK��6��Z�m�ӊ	.Ŷ�"�i��%��^��_�qf�<���x�;]^�[�4��팪����4������KVX����8%z�<A�zn�����a]/��?B�o~�&ô�/�.����yX�_M���`<��Q}y��r	��aM�2;<4؉c�Ҫ�C	˽	���6F�?	F|�g/�/�#�Ld�c��sz���*ۉ_6�et+�KRv�f䔖�*v��2�ԡ�O���۶�i�������v�u�^�^��qSm}�4�������8��`�EC;��J��u>�[f^�98�o#C��r@s0���oӭ�X�O���ύ.K�5��X�<L�Dr�]����#\U���[����3`�Hj})L���z&�Noi1�}�޶"S��d힟k,R�wWu�y�1/������lB_&v�����x�L-���~��1�+�dn������׻�%^�hZ]uv�3,��y�������u����m#u˲E���f�w����T��w�+�Q��|������T�����T������z�\�T�Ĭ1���;�d��Z7��H��e��|WͼcbΎӣ���;�Ngt&�$�w��ݤ�"�>C�<<��yy���*�w{��_�ةg��EH+<���j̾� )|�߂�z|02�M�����5���Wc�w��BS�+�8xj�ۃ"UmuGV�%�d���Db��ڶު<���jgu �jm$3^&�z�c���(���]��]lV4ֈ�)�כ,	��/@����=�������qqq�k����ߝ]a�Rp���|;`�b&��E�qgE��{�^�(Ȓ��m���s7�tez���Y�K002�u>]�k� �:D+L�ei�N�)l#�J*񐻾��݆�Y�ؿu1}��S"CS6y�;���}Yأd��۹�M:��
}\�v���"o��3���e3Q���j����H(ƚ�(�P��sH��f�;��@2;��1=S�D��u���ϒ:D	�tr&Cl)��'����~� 3��+^�v�f��t��}0��S{R;:I�wS�rݽ��}f��u����3�3�N�iU�~��d-��c��E,Q�&�z�ܞ�.*y��'f��f�&���"�tp�d)_����/��{��(��yf_��fS��{)`���'P/��T��Y��p��w��T����5�z:�(��OZ]ۖUTj��:�Xyw�`�i�s�ٚ`l?�AY�v.M+�ˬg}S$ޝ���ϣ�ޢ�X�"�mT㸹�L�y�³�-����v0Z�0m������l�~��a���#]�d��6r#9��5��-��i��i��¾y~\�7~|��ߍEH������Wf�������p�aq}���Try�N0��W d�[$�|Y�%��E-�����};խ")[vQ�[�v�΃�����5�3�	�Lx�b������櫶���{�s�}�[����c��ѷ9cv��1�I�n�ASUuq�I%���ꦸP�932�4W,���]�N�#�}&���ӱX=�7^��
�ߺH���˷���,V����|{����M�i���0g`'6�yj��u��&֙e~�g���(U5���rl+�Jd�ḁ�F:A&�ɂCY�3#�O2X_�=ó�n��9ZX�kݪ[�Imf��{��/4l{q<ePRk�Go5S�gk���Ѫǽ�יxg�zd.]T�uKh�+�طH���;��3m���d��b�:c��0�[��V&f��� ՗Mt�o���S.��v�b�v �Ƃ�C�m�h|gɚ3�>��z;���<����p9b�ڷ7
�α��-^�R�+�3C>�p
�rGj����[�縸����������_��_lzٽY�U�vm�o��}�;�<[�J
�Ӷ�V�u�ڰ7�3w��W�L��u�I�rIT��߹s�?��{,)�t��ۭ~p;}�M����-�5�'-�j�Zko���v�u�\?d>��u5�֙\.-�h�:�X��q�0�9�@�*s+�9�q��v<)������W=�-U�����ޠצ�ϲ�U˻�#�?s����_�2�mH��.�ob�U�9�B"T�(�鑺|�^�IWB���2��7��u�n0�[{ԫ3#�FY��g��wL�7�����w9W�&��v<v���L����M]nk�3��n�����Ru�ߊ���/��"��EO(gj�o>�-4kV�g��A������`��Z���l��m��v{v��\���T	�I$����{������l�n����xŖUS����N
�|�{�����M��ڲ�<��͏3�؏!vzf1���m�s����^���tW&^�T�\�K��y�-J���L�j��
�ڝ��*+vv��a����� ��B�_.�5�W��1W0mY��_�՝�}��tU�<
���#{�������E��.�Ƿ�3��+��s󋋋��������Z��u�����W����tO�U���k���<w!�8�$�K�bj����*@r��x��aJJ�@[v���׋��[/uej�oru�&j�ۛ�g|3�^�������������g���q!5j�I�Z���]��M<�W��Y��!BO�"�����k#��`�۾}Ȝ��Z�ow�#.����M��e�U��d��uan�O;ݳG���J+]���z{��ڋL����}��
�k��&��B���X��&DVM;�3�38�B{<z�}����j!�t����G(o���V�.2��n]U����b��F�S\���k���2�?H���6+j���]Fw	2���]���3�	���2w�,ރݺf��KeiV�,ų2�[y�gC�0\n����F�O����~�O�0G����
ʠ���b��.���=j9�D�.���%���]קfW�KY�V�to:�#�6jL�6�
�,s��,@��W�rؓV;�y�oa��okY�G_T��ۉ|g3,j�%$t
Cc����\׽�h���5�(��I�V-���}�l��\��U�a��Qs��R���N��PA��{��j��6n�M2����ᗷվD��ǧ��z�rwV�^\��HE�+�Q��U�#�BI�47e�@J���_T��В�d(�^�5����T.��̚����F��&�P"�L.@_c���������(�a��h:_˸�`��
�Bt���en�*���h��uofm ��|�p��Jv�b�ۼr�Wl}�����U.�L�u-�T�T��J7a��áV��j��jm��u���P�r�r�����ڷt��7%���7u�e�lV=�X��.w
�y]]P:�D�f!dp�79�mM�AIk ݙ��$�*ҫ��z��������ڧ�rڗ��X� �ƪ?;��@�'�Nb7��G��E�F�O٧ ����{a����._N͸� ŉ�U���2(�!]0f	��xqe��*B�R�$Il�c�W��Q�����Վ�W�
��B@}��u�TM�O�mV:��JX$)zyްΡ��!�4x�����%�f�`]i�X��z]�t�U����WQ��{�o(a��^�ƺ��;.��j/3��f+K<:%�S.��E��f��˥Zιe�c}�P�1��u�=sm6{���b7z��*�کu�zrӃv�bod�0�Uf�k�.8�x�[=�H��S���r�ȱ��Z�wZ���-�:�=+�֊T
�KI_d�Ivc���c���j�zQ7T5hO��6ص���p���Q�8�����u�Z�;V�<ͬ�v�[�35�
���x2n��mYRޭ�o��v�6Csr3�[���kNݶ���7.<U6�Jx�xB�0mb�Q�C$y����#�������bN\�)�*jw.���a���o/k�8q�j�Kk�P)M�8ҙ��2����N�U��`��-Vp��\��e�ޣ%Þ�b�競kE��+;�|uFj�v���6^���>�ۂA8e`���u��}Ank����J��s�W�CL�[,�"����.��xb���g˵�Z��2(J�DusU�޾��:LJ!��]:�b���m������otҾ/�������N�J��t���=EUTUC&C��|���E��Qf]�X=�����/�O�d�-�u�ڛE�$��1�����_:Ӯ�뮽=====<x����@��I�Cj�"+;/�X����x�-O�D��p�
��9�ۏoOn�:�N�뮺��������Ǐ8��I!&��/ݨ��H<�����֪�UMF�BI.5#�1��<x�㮴뮺�OOOOOO<xﳐ�Q �e��,�\�#��Z2�	$ B$�Tӏ<u��Zu�]uק�����^<x��Hm�RڲL�����DD�qv%�hS�;1��}{p��nΎ#���ߪ¼�B��Y�g���k��k���,ɭo�z#�3_���`Q����m���3�.934�/��/A�m�2���6γ#��m3e����N�.u��%-�B�"��cKb��,[��z�ʃ�mID_�sno�Y�%p�;�x̌��}�����u]Ð��A�o&�hjixgV"���ʡ��g�x�qqqqqqqq�d��}�)���v�ߡTI,�a{lٍ�Yᦜg_��:⍥��o�"﯃N�x	ox��;$�Z�{R1��� �1��t"�ƞ$�����VT���N��h�Uhdή��;���&=�7L�� �<UH����9����p��b]�oN�xߑCgD�Dz
�.�oԟl��y��E�����:���_o���T����P3�	©-���NWe���3r��/K�]b�y
~�,�1R��ȜХT�31���؎��ДK�5��ƟV_M�t�S��N(r�ktz��n�����l�^��F��=�e�|��n��Ӭ��⹃,��;�ݢi�V]r�Z�-��3����~����r6��H� �o+��=͙�1�	���X�l�^�=�������9OJIu>������êD~������"��v���/��Ɂ�u{�'E���8fL��ef���H5���e�(�L;/n�����l��=}�N�c�'���K���]�>\���{�f�潱��^�j�ޛ��L�-���M��Y��>��i��i��~���w���6��9��o�n�on_��N�{��("��5�}ֹ��ְ��QP�áLT�neZ"��o3�<P&�ze��vm�xh6{Sj�#}������{���[�v|-��˨A���O��<s3�'_z.�;5l%���2�g�5�	�4e��˙Q�����<u��K����)����+��|�_�/�i`�v&�"�]6�pN�:�}y��PKfBZvkdd�Mo��ʵe�;���/UO2)�rmXn�
���)ƭ|��	jW���Tz3�6*���y���޶
&������V�{�wX��#2<�id��A�S�\�;*k|�]�n����V���dU���ԁ�f�_V�h�uY�)4��=�8۞Ǘ�,kǈ�j�_+����X˛�?֞!Ikd�׈��lڭ�m��_uC�=����$lU��S��6p�Υk��YN���>k�1���t��ٯP��p�un�b��Á�����n�x��eɽM��,�[f[���h�I�D�~���~�_�P�ȇߏߩ\4e�<�8���2@['���.5r>��W���N~fɸ,���D��fڕM�����`��M{v�3^Zj�P���q%����f��1�A�Fx���]���G|׫&ƈ�������N;�	d�ty��ee�w �Jkƨ��	kX�vK�S�f��:�f�k��Q^"�W��b�[�RިI�3qa��` Q�y�RQ�e���>ݶJ^���o@����>b�[�~����	���T�U7�-S�K{zQ�!��,��V�m^��jS7So&{�06sS;�׽е]��N��*�
��~����,�΍�E+����Y�v�w�{S�vq���u�آs�:�r�9ធ�2B/�~�3�ݾW�ҧ����t
mn�a��<h�k�&�4��l�6���}�R���b�P��U���::��P����Ӻ��<�f�r�<�R�� o�X�8-d�Mr�Eq�In��F�6�V5	ܵA���"���v�baj��ˉ��]p�m�ft���N1w}���ͮ���w�*�v�T����h��TP���}�����?����bŻ�׻�=1�U^`��c�n:�IP+�����=�aF1s7x������~^-��A#���9�Ϋ_h/!�WvC;���J�G/ ;�9zAh=>I�,b�8��lĮ�L�'�T�֭�[c՚�V���s��CH:����6�_��f*�nqmf��ٹ��j��ߣ�r{Ӯe 5H����n����k����Wd�MS$�C�O5G/�3z#4��4�	%�S�^-;"X�����݌EM��O}�E�6^���$���u��]ۇ�#s�-��f��/@`���v�Gg�G���-;u.6s�N����&�M�K����
��c�t.��z��8|��w�Źk�����X�7l6|US��%!��[M4�FpVP��
a��k�6��i�/ί.͞��y��:�O��e�;����/O;E�ZVh�妷�z�N�������x~K���f�>ܕ���3�b�5:3Q��h�pl�vGy�)5�]�9qE�彏;&�V�R��k��G�V�Ρ�>����������n2O����;W��޸͟`�(��j��ZSk�����EC�9�i$a���0fn�\t��QSㄙ�#x�����_�(qg5d�,MOF1��)�{��#�b�wE���oC��1�VGs�^�,ܞ�\���l,��a��t�פ�NG@|ٲ�����iþ�b~�.��@wzu����d^N_��0gC��qx�B�!G7���]��t=���;����<	�����ƃ���rۍ1%�z�}�>&�DȘ����Y��
0&��`h�-���L�C�sV���Z�H��<E�b�Z�wc�(�k���-Ozۦ��:���x�g���wy� �7�\H��15'1��ۗ:�zx"v��z�;yt�)����E>;P1��9�wʄ>�<�� {I�Z;�ޛ3j�c.���؆���KS���^��z;i��+K	fa,Ku�A�˒�fJ;��XM46�Pc�>c��׼�m�/��ocݹPf%�3v�˝���C���0��]n��Q쎸C��򕞏w��G�������FՓ������4�[{�c@��c����+��\�s1=)\mi��"��k辄���ZM:��G�G]P��L|ɝ�KV�c�`	�
�|6�w_���ګ׭��Ew�q��,R�R:��wf��<�:��Y�zBԺ�ldvlڈC7���n����1��G�za׏�gD����F��M3�ԄG5����Q:���%�u|��1�<y[�ᐸ|�_>Ok���jv`�m5���p�L�����O8���.½�a���\|�;����S{Mm���%�׵i�W�JiV�ʾ@CVױ�5�ݥ���Ǝ��{gf�q�/���	f�^� �S������i��߇�<252�j������~0����^>���^�����A"���0�O��>W�>�ǅ��̦�sY�����"�f��uڑ��gN���p��ged�ʇ'���W���RS4���!Ӥ{c��>nЄ��MT�s����'4o ��o�������-1�����P���Rl[������8)������s����qqqqq ��[��__���/!0ڥK�;;�w0le��}�a���Y�s��Wj:.I*ܱ����;���Z\+�m�f���(o��0��.jd
��哯�;��v��pGc!fGq�'l�ؓ���LJ4�?R�]�y��F=���yƞ��5W�i������sc�\��aٙ��p���H���yY�����U��h������{`�}��_�ە�t�s�׀�`��Ʈǲ@A�j��XO��s��]�B�.wI�߯�K�al�@$Dz�W��(#��[FkQ�XKW��M�Fx՜������Kc��ý=�|l;ϗ��I� ��Dsf���Ѻ7	<���l<�Λ�l�[t�9z���h���9EG�@z��nt|��}sM�D�1ZX�əwv,�ɸ��sf�����¤.�2�VoM���cse��"nR�ՑW���^Z�4�SJG�-�v�|7^��#��c�+�j\����zr��e�a�͚$�@�R2@�J,�zW[��w�٠�n��C���^��]
�DwiY=���'Z,ɤ�Xz���ܜ�Nlj�:�W�2v��7܅�f�rd�:�l��i��i��y|�|�3�>���_
;�U�cд�H�$h���mg�A��W��Ӹ�9�E����r�v�q�q9�|o�����#��ľ�d��L5µ��n;k'ƽW��;d����U���>�"�1pf��Zs���T��+�!^��˕A����=���֔q��]'�i�׊贱n��Ut�F�|�#� gHq�TWv3��3��G$���J3w w[���`�U�ɀM��#<�G36��_��"�Vu>c���v���봶�����j�\S����k�YaH���9�ce�\_�����x�<Y�\mU��F�}����Ն�x�>�^r�N{!�n�
��������v���R���o��u�G��q���2��%�])�a���Q�9X���}v�53aŦ`��_��j���͗��_J�?Q�6e�,���-h���|�d.7���[Wa��.�9��/�8�n��b4!�fLއ;f�*
��kS��FN�Z㛁��P�m���&�W�5�N�
�w��u��Yu!]=�i��i��i�Ei݋�^��!b���f�C����W���aϰ)�C�y��4ur�`0�#,t��d�����w�k��գ;Poǯ��Y�e'(����?@)������j�
i$���n���{R;���q���Ӵ� �-�g�fe����|+����r�"_�9]�1�S��R�[&�}2q{{�}S|DQ��>���cm$�|���\`N{Z��c��6ߗP⌌6tV;	��Ȕn;̅��#8��	���r�Z��Kǜ�^�|���uJñLY����p�h��#�oe�98+��ۼTs
u��;�x�,��Qo��4\,K���h�g}��L�r�7�>&-[����2��1Pka�
K�s."��M4�ć���f@�f�4�]~�p�sgo�^`�KʬHގ��o`ވ�ƻ=�$=%}�y��Ƚ�;��$AF���W�{>�3�0sU��]z�ĥ����Ӳ� 3;��6ql���}v�L۶�Y}[z�5�gi+�u���\Vk�ov��{��2�xt�8tVo��}H�)>�ړF��}D����.�Vy�f�f�3��������VsjV�l
���>>>5G���ƽx������l��lP��67f�7>%���O3�+���5�5ll�U��ö�B�0JC��0-+�ާ�3�uꇚ̬��%e_��us;���2�+	�:y]l�;�(��t���w(��R�e�5�^U�͗�7��YJF�<{!�n���{��q�&'P�@�3K�^Ϗ~���� �ߺ�'Z}�{7Lv}¨r�>�$�.�Lgވ�I�y	���B�	+��u���O�0��| ��`;{��ꇼ���8I�a��.f�����<(�������?\e[2�m$�嵤�2q]v#w���[�=�1�q��pI.�R�T�l�����0�;*v�%�x��;�D���ޖ���i�v����N���N.��ϖ�g�ve���q�K0�|Y<�<'� X����c�c��Kwd���e��tj���ׁ���^5�Q��T^��"�,1�z�H梎�O
�|&>���>�lmC��r
�n��;TDd:E�w%����`	��'�����ur�1#�Nmp83D�M�.�����X�H^9r�q����}Mh0ѩJe�ڃ{��.v[MkՏ��K�g>��k%��E��h.ط�\�҄Ӝ�6h,}Y;�]Q�JxGq;�P��84@�}L"6�R�i���v��<b��ď!+ef��_n�AN��z{dl�\�[t
�͕��Ҥ�_ i��8;QJ��&bB��zWC@�v��bkx��+*�7OZ`]�ۓv��{6��8�����v��U�6fS�UA��^j��pf_�4�V��\�j�n<�q=c\aK]Jq����l�R�j���K\o����6�5ފA2�Q:pn��jzaHɋY΂�t))2�����Һ�]�D���Ӷ(`J�ݞt9�*�U��3�9%^(sclP��U�b�Ew^�יRo&�o�^�J��}���J�n�*��}q!M��t��j^.��n�^0�$�s2ث��5���fG;������YNpde���|��*n�z�*A���,tz*Yp�KM圸���↶��V��@�X���,2�	�V�%�#�nR4�^$�@X3B��t��^[.UmV'%���U��m+I���s�c*�ç�JA�2)4�%�f^�e.�{�0Y�U�W�������3n��G�W�G��k;a'x�e*Z2�f�v]�ʘ?�	�L�7(�磲�,��մ���oS���U��to��V(�7�n�F�͹б�w��'v���ȰK{z�`��zn.[�7Y�U�:�vr���4�3E.�S���|1O]�*ڤ9@��M��i�HcΖ���3�غ�[��I�uu�F�h�^�V�5l歱koUZ�Ʀ�
�z&3m��������AUpF�3`W�ګ�DK�tWV�Ec�{R���Ǣ��N;A�g.���81]DU�s�UEr�
ј�7鹠��3�\�q�;��n��	�:�:�B�eӼ-�5MS{��Z�Χ�r�^���{�����H.N��<1�z�u�ДiU�l�0��nݨ��&xF�œ��7�q���;���9-�����n���Mr���xŉ�%I�����zy=ћת���s����H�
1�j�R�W��I�,s[ެ-e���:�2#�ȁV�Έ�'�8)ȖS�*]`۸�u����{�S�v)h�T`�LIg��j�{g=}B�T�;s��M�q����S��u�j�#rBԋ"�OnW������<(P�>؎"�h�5��%J�T�eԍ1��u��:뮺������ӯ׏�mT�r��i�%'X��@Z���B,٭��G��UMm��<u��:뮺������ӯ<t8F0�*�UVo�����'$"|Y�HĄ�ܩꤒ1�=�x���u�]u������׏<��B�!���
p�!ل�)Q�I�P�d��PSO<x����:뮺������Ӯ�x󌌐�`�F1�a$��*�Nmeĭ�	D')��8�%'mi��//+�T�|�^���q��v��]�}1Z�i>mN���`���βks�͸^��X�NQE"��{y�j�N��N[��9ĒK�P���+m�#��\��ֲ�|o+U����ͬ)E)Ȉ�����/3�� Jyd�S��)%�I98:��+�ĀH Ĉ'�#pV�KtJmЉ0XM�M&�i@�Q90�ċJD�i�
p�Cj|jI1$�	
0��6�|F� �с������-OE���}��ۛ��L�T?m*f���,�����lc0ruq�������p�E#x"��#m@���-ƋM��mC�@���-����c
78�"&A#��"�A���h1 `6)����d�i��DGP��1��1)H����<��GpĈ�(�M�!$s��QI�؎I!q06�qB� �B�E��V[��,�UVf�<i��i��W�%�2���B�G�M�]��?s������S!����������e�,z�&��z.�5���w9q>�O��fF��j�s�½����D=C\'��m��SǇoze�s33��8��șo�)g�[vmy���Ğ���mh�����,՞���#)���t��uW����v�4*�w�Y��IaF\{� ���W�U�쁯�"�RӲ���y��*���7L$L�p>���#0:��r�h�`�XHE�W>te���zlVϻ��R٠h[���l]M�u�}ݷ+1%[����<��9��}Nf��]���5ʪ[ڠ�ܤ6�b�z�{[��][�3P}�O�}�c_H�S,�\�:,����le�+��iUS����~ﳒ�����������Ѳ�#"碲bj�ެD�xwpίH��]P9�"���w8�M%�
?�[�:�v�����<��L9�`�"�]v���F�t���ǜ�I�mv9Y��<�iu^�u�E.�ݻ���gz�o�)�u��ES{ �ܢ��S��j�2�*_0o��vb�zܗ֫��
���{Kr����^>>̲����xhm
��#�8���@�r�I��	��a��K6uTU�Mg��E[p��T��V�N-η��#:��R�)�f�bi��a�.\{�C�Ƕ�wZ^?q�����/R��x�yD��}�#��X��╆3���F̵�ǲ��ߟ��aO/58**q��g��x'Syb��O��ˠv�;<��5�;��{��s'n�����Tl�DO^϶�7����؞��r�R� X{����5zg�S� �� �B�G*���uz��}��j�^r�_a+�鳇bf!����<8k�\f���y���w9�U�|��"���z��cyw��0���ő��{�vR����mⳋ�՚��*��µ��{S�CHQ�����/�@4b���ͽ�,Q��/�������j�Lť��ՠ��]�ς�ir�z�7c���k8��RM\�X�-���	�GHg��5���tQp����0�:���X��%�s}D�l�ٽ���M��py����)�r]B����d;���|s���nIs�~�7�ף�wG-	88l���>��W�t��h�R�x�;gXg���j*��K?�ѝ�4�W6��c4���͠GM���ä�H�G{�f��57l*�Gf�G)�i8x���[5^i$��n��s�(#���^�z���K�LM����w�Q��n�Eut���F��s������=lqnh��rf3��}qC�c\"�ո�N���ʽ�T ���Q���&��am���Z���Cd�\D[TW�%�"��n�u.].�������q��"�ݽ���
���[/���(�Q��^kG�ڧ����の�A�Q2�3��$�VAg��;�D�������/sD���u��*���Oj�ό��F����$��x�����ȁ����Y�ur�8_��=��3�65V4R�fͦ�%�d�N�:��u�i9�RG�HMF�
uH�:P>߾���Ǚ}F���RS.��ύ��<?�6�;9W�q]Mk��PZ��μ�6��!7��꒚٥��6�.Sܐ(��'`���6����7����y���s�e{s�[�>�����
~��:�;<�U���-��1�q���܁٫c�q�4��R϶Ϲ��c����W;U�j�[}g�N�d�][S��(<���Zi"k����O��=^�_�I�ޭ罙}��ɍB�V�^7C-<�]w��|�*N��H��^f����v�����qG4�b3�έ8ޘ�7��r� Ln��bk�üb*nZ����h�m�I~��vp0����U�b���g��;^�s���f�2݉z�Nhkj|I����O�E�z�<��H]��S^�� *$�������~9� �i���St����
��ث�H�g�p��ް"��js�]d��'3�+�Z/���	�k�9t�6YЧ��p��a�k�A�[}\�ɮ!��kǕ⎑�מ>�˚{������be�o:�>_%�����`�U�찅v1��6�XQ��l|*dp�+�щ|��\1_�fm��y>�>�z��ԑ���?�3�v�=���ꚝ������q��q�Ԏ��Ǝk�04�e�Lnj͕x!�b�*���1��w����,�
�{^]����J����s�D��1eis����[z�9wk0���>x�{Q��]FMPE�ܫ��ߗ�|��>��,v���J8�(�ګ~7�.���޵,�0�o��@H���ОsD	�lw�����>Dr�y�S+��$�T.{�r�z�r᩹S�qأ��{����;����T���U}��p��kKs;mGK0���������J������\Nc4��C������Ҿ>�0j|�҉^%��Ꮔkj�z�:�r�ݙ�7��\�=��1��&�D��*�CH�g�j�q#�I�6C�VcE^�^�w��Dv�G@{�����z����+��W�7wm=��S��ky�O�����)K�y{]�J�T���:����<�V�{���[i�M���w�ay�Y�RyH�w��ܳ[!��[7�Jnv�6���B��Y��!�ݟ������zt��3f�36�H/���w��6��;����o[k�����k�q��y��]�wC�X��\۲��uPg]kya��7x4G]��Ϸ�mn:c0��1A�$�m���)�s�gr�N�W[�z��_n�Qi�����g����y��`�}6K�K
�̡�!��#�N�ڨ;�Z�0c���f�{����O7{l�����D��3����@�X��X�`���+b��7s�n�-�K�^l�j:#�d8����q��ȋ�V�W�L���#�2Q�d��Ơ*:��O�q�0q Q�$�7��<��u՝q{y�rq-[�x^A��j(G@t`u�U���:�t��+���[���u[�#�ŗ:��H��r����þ?Uq���ub�t37Z���Gz���sC��v�A�-���{����ڗ������p瀶��aZ1泷#OlS{��;-�W�i�m�F�bG�����|��~
��1G8٪�u*��	/��[�;�\T�=��/t���x���F���9ad�IE�GC�@�v�������w�S���3���7?k��UC�Fq���Җ��EѶ�J�е��R`+N��Ȯw��.�B��)�n[M%����T��|�xI��Y�;Z���g�g-]!�Nww%�����+�+���1wb�G�!\om�aN<X��C�xz1�c����M�$��������q���l#�7�3����;���Znf*Z6�<�*-ns{�UХ�¼�W�F���G���M�
M�>�ؔ�^G�D��O�}6}�]��P��[Y��n,��b� =�����Gw*���ȼ8Ndb
����+e#~��@��0;X2i#�W�M���X깒IMG)���P�WR�v��)-���6�N�*a/-[M���ie���+\wpڏ����r�{R�d��CHoV���t�����/V���g+���4l�}�X�D�Ϫ���̊�eT;޼]�=5����`	�S^�gz5�s }v��1R�Ҫ)�	s+�;M�T���>�;k���d�^�{����t�[/4��.X�0�z�lE@S��b޶꺶v�W{��Ǹ��0\���4�4�8-��}fIP�b�MAe��#��[�3v�G�n�M���:P��f6D���0�7�WE�eBc�̻˺p�1�L޺�i�o�cs����fVuw]�rH��Fu�k!f��Y:7[ՠ�IWɖ഍�~��������r?��}�@�;>ݎ�\��S���FۡfR6Z�-����Uk4�*1��[xX���v�#�S���ᓼ�Ӗ����p�l��u�x׽�š[�98��`K�{��i����\�9@�X�5�L��|�Uvg�1�P�FcϖO�®�fzΘk�sZ꧁繌)���	�L��4����#�q���������wD�+q0���i�)Hw�Z��{����;�zܯ��� )m�Xs��|s�pp3�5{F*ߎv+ywf���}�g��7]}Kc+kk2k�ǋV�����`_�q{D�u�`�����o&�k��өG�����H�e]Nv�̐�|��0.l������>���/f=�\4z:i#ƨ0h/d@�UKU�r$'}�m>�g��Azx�U�l]KH�; �5Y�t�&���8s&���DA��|�7n��*�\��L,�22��-��I��H̤��^mt�[9�y�D^1 e�X<�@v��WV�_|̭�v�쇇�X.�K�ѽ��-�;������'JE��-U���hu��5��>>>>>#�*�Ӯ>.χ�X��Cl�c���8���2�0:YV;a�m�/A1�\1AMQyk�7��n[p��I8|�G�-������:�{�ܜ�?�xk۠�Q��V�:�J6ze)��2�n�#���R�z��l�<g1�_��^�V�	�����	���;�7�nX�����V!��-�P���8�%?w�?��j��r�}*�'%���M+��l7�gq���MNݳĈx�Et[rч�>�e�nBT{<p��-�L��0xh�n��8D욖�9�x��e�P� Nǹ��㙦P���Q�I���5��P}��o?oz�vC<��ho_:��Oٮ�5�閼��Sݤ=A����l�0Y f����>i����(�n싦3[�ɬ� YԖ{d��$��hoN{���m�t�Akx�'w{c����6zd�1*�R�n��΄����X-�ob�����{��|�IU8�pybZ�q��V�����;53v���=���]i��Ψ)3�E�ej"��b)f��f��ыs/w�oY:5fZ�c{GW��,�sTk��e�҈�1^sҤ!M�6�h��|<<<<*����;W���0��os������gw�Gw%3C��7�S`QS����gs�I3�g�ڸ9C��c.(ʗ�ƾD��������5�]�l�Ї��ot^�@��[�A��,������|�^�R=5w���n���.�����7���F����	��^[�^��>�5 k�vꑥ�$�l,oC���?�
�W����c�ҍ��7\u�n�̳K�e8F�!��ە�/���V���\o;��3D;0x{�C]��W��=/��zkDv�T�x��{ݸLS:��e�Os5�%8���eݵl���z�M�s1{+�\�0=|�J��w��Y����!��Q���{�b���u(0ѕ �5|�:lc0fQ�\9c"���z���%YS���)��J@M��;oM�����P���@�;Qf�7�;�#����Q�骨Nѥ�L�N�����ˍ��������w�#e��f�oYթ��jw/cG��~��j�͖����%P�>J�,:C��f�{��)�N��Ւh�u��R���f�Vv��7Z�f7��,](J��:
�حd�mQ�]r��K8�`3g^���� ���G	-����C�s��_v(�²��4��Zd�69t�v�L��z��ͷ�/��2g[o��'ϴt�	�8n��j0Wr��R��p�w�qS3�B����K!�r�Ѩt;ݣ�>����Ua�J��g;T��V�q�]%aa0'XUֶ{+N�Y�	�Ѡ�6�p|9��^G�G^V��\��#Z�N<)yhA�v�w�޸�Fj�����CtG��1�x;��l�[���ȧr7�u
}�M��{:J�%��-w3xw��� [��zƞ��ګ`��X�����y�f�o�A4�E]<���UDY�Sq�(7PK쑾FS��
���Yɻ�I�ˎ�c�ڔ:�ڊ�s8`�&�+v��毉}Y(�C� �r�ЬJX�CH����%xOks.�٪�x �h�wk��:P}��!C7;���w�R��%Գ]�kr�ੌͫ�\5���GJ���O]f�t/-�+�d$��T�	5u܅A�:C�j�/�l�.��C���Ln��v��j�'�8	lS���!��+,2K�[(�[�r�5<��5�L^)0.�U�h��*�Rd�@ȳ�+O
�}}�4l�T�5 5x�U��=�3�sݮ���S#`&��r��j�U
��e�K���D�����m��S�N��l��Lr�R�w��N�Z�a(j-Ȉ��2A#���M;WR�pJ��sPN��U[額'�a�]aNê_�4M�ö��i�ZIWXuH����e�-��c9����x�U�v9�ͮUuT�u:�Bd���k�4�w�Ch��Ymq[�#�®Y�΅����:v��]X:֪�)����e^or�g%ogU�� �Q�J�wz*���k#n��T�J�V�{��<�3Q�ft�7�wu�@�9��wq��5.i[���:�6tz��%pR�*�{]�To��&�}�ۼ3rP�$��b�`��f��8��P���s�j�[��s����l����-@X֜�Vvs]>�4st�n������Sa7�6b�R�Ӕ���i�jU��� ^��͂f@����2X�;��9���Gq��Eg<B�l����M`�̹n���w�)+M�#cm1LK�}�0�t��BP��V�T�Ӷc�n��f�݃T�g��#�ņ��6ʒq�� 
 x
�f��@H��X�K��(W���}hΐm���Rq���w�||}}u��뮺�������Ǐ8A/�DHS�Y�
\鵢s���j88N9 w<���[nr�l9��w�q�Ǐ���]u�^������u�ǜ�:I!��9�k����I��dE�C�)	��Q��};w���8(�zĩ�o>��뮺�OOOOON���߽��A��'��U���b�mD�q�v�C&�GG6�s��p��!�]6m��>>��뮺�OOOOON��Ǉ H�l6�ɰ*�%�>n�+��隒�yd��Q$%9)Ü�Ϧs�s�I"q�	�D�˲��9S�@Rr����o|����c�bNYv}��)��|�Y�>��補�Yh�I�%
�ꎯn�:�J:;�9˗��(f�/��r/͑(����μ��˽�J%�ZH�ȌĄq\t\^Ƹ�f���	."��C�lC��بH(�ͤpO����8�٤�X�I_ŞwiN_L�'��Ǟ�ν��j�v=����@U�x�ز�ں���0������p��%�����ʝ"Kn)I�uX�H�iP~��������f}�g�	Qpf�&i��m�N�4dn�K���ہ�O�l@��y�����U�3o�x���^���q�<Kl���G2��/�y��@3}��A�|�t2  :4�c��K�)D�.��_$��rk6�kU�P����5��5ex#5��]�A���$F�YS�b�Q��D�DoT�h�@l�o���ǔ�Й\�.�<oϻݺ�uY�&F�e��J��NO�7�{�0p��X�z�.S�Gr�T��5z�v"��Cp�!k�&�i&�mn�F���hs~��֚�(Pv��qod���S�[c�=�0�@2����2���o�߳s��l��%R@�f��w�X�%��ބ�#�����i��sk���F����㾏\策�aJϮ}�R�C�W���5�3K XM�Y�;�rC$ͪ~�y4�a`�f��[v������H�p�;�	P�^�kL}_u��Չ�MK�(k|gL;I2y�.�ը���M��MN��r4�;r�cK���1��R��՛��C�޷����C0[T�>��4(�²�LML�T���Ց�4��}Jm�N�(���૓{���V-��tK�ɯB1����m���|Ęffc�(B';�l;WQ.go��ע��vHw��L�4D̜~����ܓ�����D�����IH�1.V�8qx"��q�-�9׸{[e:P�?��W�7a*��̒�V��kzW��&)9Rn�����F+��wv{0I��Bu����b=Z����~�o��O�m�oݼw兰�Th:��;���:�Dp��G�O�v��y���;����L��jS�_mVq�Y͐�ϲ�K���CS����yP�y�\4K�Ã��8��"�ͥ�&|�<���Tm�7yCq��@w]�9踫���y�g�YZ*����7j���Wf�"Gt�)��1�~��M���<��v��q���1V}lή����@���\9-�\VЅ=s��6,^�{'B�c�u
�۳wV!b^>$�אe|O�q#��Tی�ݵ�5Y*�X�W����=��\#�uB���{���vVoZ�
�de\q,=��P���WX>R�n�i_f5F��ֺ>W�x���ͺAf'Y��a��k0r(o.���n*J�6`����~��ް�_s��&���q�+Գ}'/��Ս
��)(�8�.��T�暝����ʂ1���U蓁��D?=۬��R�03�]����T�3��4G��y�a�B�F�Nެ�L��,:�F;:	ƎK���ݽ^��B�sa�77��sS�!"�٣ ^9��d,+�z}��q�Т�?�s�A�9�[�4�*۶,�����R1J�������z'e��	���Nѓ7q��^��{�b��(�zs| �$�^Y�]1�g�Q�13�U��8�@!j��ǢC׫.=�߲�$���H��)�J%K�P��������s�W�WdmnBTx�E,͖�=�s"7K�]UR�Q4� s�W>��A�"h�f���s�Vq�v�'���V(�c��n�g�x��m��wCҐ�k�П���$Yrg���+�e;4�1V��4���>BV���0M<��l��j1K�o$�*E!|�w��sr��4y�r�J�פ��V�w\xj�������������|�v�W[9�G=[^J�P}��~�@~PC�œ)�t�dU	qUo��<sV��J3�[yc=>�; �'��L��\�o���Q2)�[�F�mML̴<u�:���-,�L��{;��}��cu�V��
��[����l(оp���*w3�w�3���Rݟ+�z\��)�%��j屻�d�#Y�t�^034����\��Ԓ���;�e�Q{��iw5���-��U\�2��8i�L�"2〈~�k�)��ڮ����n�e��n
h9=ھ�g�ːfȬ>�p��l��v_n����<*I���)�Ӆ�-�ܟ�tǍz���g�@�`��g�5.�%��Ѩ�9}GSMj[�����w�{����r@�m<�t]���;�3mS����k:@���;�!��X����z/Y��4-�H�O�읫_�GNB)ٓ�]΍�]�a�ʈM�WD��ל�=%�s�uwU�7U�$=ˠ�կk�/OK� �Ά�c����W/��Uē��;m`+�,��WWͼ�S��������}X�:{����Mt��f4Pv��C��0^Q�
��g��F�	�I?�oGl�W�� �B7�ۑ�#rt����ULT4��
j��֍]��`{p�Y<�o_9'SU�Jf5y�Ԏ@���������[��N_�����P��vk��X�Հw� %P�fA۽T�-|�uA�r�����Ϟ��:�DnD\L�;Ä����K\wwG�};r�{l����ӝSQ��z�;w}���ZtdҿGGu<L�m�33u��$ٶo[�&�L9;���TL�=��C�^���t�}U�������:�ϱD,ډ�ڲ�-���"�i)ɨ��y��[�6����;S�={��=�=U�����Sړ�^���;�U��Н�m}�bRLB��`=]A���0��x���w+7Q�#���e����m��Mg~����mOv<w�m<����ӌ��ܻ/�i�𥽧�f��Wb$�co����П��Q�u�&�֯�eIgE~e�	N��8����C��z,,ĺ��N\��Vv
���agS����ZW9� �����y���N�����v_wb��NeA���� lǫ�/̇n5���7:��&���)����x��+U�d(�!C��ݩ��g}��WmH���K�sF����`�P7cgۢ|�x%ހ������d�O835Q�c� ��y�yʅ�KO���A�#X�e�Լ�=a9%��>����Os��xB����sSC�b=�b5&��W���ى5}��,��|k�QwӪ�3�.�sUg��S�3�fX&�2-緘c K�'�m�����8[����*�v2�a�s�k�j7%$z@�D�de��#*��)���j%����w�3$�����xMH�Kė����޸R�����[� -s�;��;]���^����W*�ל"tP�]��Q�>y͗'�w�	5:1?�R�6Uc9��YWsw�M6^��<��I)ESv�w��\vm��y=g�� ���G2�l�1c�-���;�0B�7�L\��,W0s�����坑�K�e�7�u*�<���3���`F1����J�p�H�S���ӹ��e�t��;�z�b��6Ī�/����y���iⰅV� �h���'�d�7O�c�|�� �qS���<D۳WE�T�/{�O�U3�[����նu���l�M����qt���e����f���7p���=��L�@?OE{q�hfa7���!3;4�W��j��s��gKӼ��ܼI��3���[,��'��o9Mt�qݵ��]G��!�7�M��V��a�]������=��x���ci�t[N�@3����#ϡl8�`��tzξr����~�����5���1<�鐣� ���r����t���Ϛi�m2�3����C���j����O��g�h���w�@�y"�黮q�3�]�|�G�YT�b�ҭ�s>���yx�?�GΨ�^�:�|�';�O�锫�kF��o�[�:|�l�(�w�n��l�P���3~�*�����۪�^��U�Y��y�[��W���c4�pN�22�Wc"��`��e���S����"���v�f˹���y�J��B1V��gU����(:�r�c�6+�5�q�̗|�T�����Ҽ�y2�7c���y��o0`ݢ���j�bf<ޏ#�Ҭ� 6��>�x�P�njz�wU�t�	>�o/!�#A�!V���Bۀ"7-.�IZ��w�gׇ�1�t��f �SO�(O�n{-ml�Y}��|A����"���~�����������y��3���7*�\�zi>i�~�5��n5A�~�d�m�^��,K��n_�Y¨�=>�旌 �#��WA�;��4���"��3��td&�j��{��d�359�7�\;�h����
�с�0<�g��q�O�<���m𾛰�q���;g�� k��~���V^���mtHKu_3�3�͋-���p�m2��Tw�����Cq�L� � =�#t��D��f��h�Y�ƶ�v6�6����R����g��#O� �8m��o{�9��7`Q�!�ݕ����ꛖ�_��&���v:�W�w6I�f�v��rŒm�⊭BW:�(��V^��"h˵�ʝ8�xkŏ��.0 �0c� 3��2(B���c.���:���P<�]�*k�9*s��S�K���f*|�9ǈ�3֖�r~��¨xU7�v�:uʪ�5U�yOG�)\)Y�|�"�3�zjF\��w�b9�r���d��;#��$<[����$�_���惜�\FVh�7m�Б�b�z�e��Ae	�
2[m�(��Mk�noaZ��C*<��>y�Uo���x�Gy�6�;>DDDC�瞧Y�g}�lq�Z�w����
 p.�IP����	�ގ�**�][��	��'](�
ꉖ��g:�� ��U=(�_t���ң���kү\�B�}���gRڠ�Sêp�B>s37'��K:�Թ�S��LA`;�2xʯB3>;��o���A��2n�˝Sv����c�7g�8y��X1�`=�=��F�ע�9o��][�\Q$n>.�Z����,��nz�ˮ#���#F�����MK��:�Gdv��P�%��.�
}s�%E�XHi�Q��b�mj�n��fA1���n��̞�7��\ø�X��l9��u�����XlY��}����M�ʼ���;R.+
;V���zN�����~��g��^1��`Qכ盼�X!G)�A]�����߈�	�����mAW�C�B�kK<�z9�5�_%�W=��B�xe$>{8�Ȯ����^번[(�ݎX6�36�37lp�Ş�t��[^z��0��7�]B�m���K�v���Ґh���I�R��ލ�{�g�Ѐڄ��#�f���u�fl���b����\�:ùݡ"iz�v�l�^`���Bn��7ȣ��n�`j1uwd�iv��+S��UM�T-�����D��!�z�j^��q\K*��K3P=�m��5y�|ND�(�����p�����&�Kr�e�[�x��Bwxa5ٽn��v�S�;�,��/\���x�H���H5uWv C�j��p!&���(9ﰨ)�8$�y�3����!#�>̨�������*��@Z�b��O���ց�""��6YQ���wX��3��0A��V!#HEc"E��RX�20"1� �@��4��qr����q�r����R!#� Ȅ H2Q 1#�`1��'뺜q�:�.��U# �0##�1T�Fs��\�*��qr�����R#"�#0T���qr���'*�\�r�r\��\���s���#��R!cH��U 0�V� 1��H��1P�H�R�H��HT#�EHA"� HA 0A�1��BH�1D��BH 1��BH H 0��RQ 0��RH2Q  0��RHU 0�� 1P�1��R H�P1��BH 1����0P��BP 0@��P 1P�� � 1��Q 0��BHU 0D��BHD 1��R D 0��BHD 1D��BHD 0D�0P��D 0D��B�@��0 `0�P0F`1 A��X�0`1`0`0`0 `E��Q��E����E��c��� �A� ��P ��E ��AF؂�0D@*�� 1D  1 0T@ 0 @ 0T��@ 1D@ 0D@ �0 0��HA.�� �0�� �0P��BHD*�h��D �1��BHA 1P����m��U 0�� HD 0�H�R��I�r��ʺW:�\�r���R� ���#�@�u� u�
;���PQ	P#Tc��
�������{������TG����cH�W�����?��?��p7�����O����?�
 *�@G���:�����@���?�}(���)�b��?���P��PW���~��ދH��;���?��a�1=�+�����I�X��EBQ"��D�H,Q � E ���D�H E, �H�@!�DA �H�Q ) H�P��Q �(�P�A1D�EB"��@A")��"0� HD1P��!D�D"�A"� DBP��D�D�@��E��D��D H1T$!A�A$TID�EEDAސU *
 �H* �� "�(���
 �`�Ȉ@�$b!"	"(F �`	""@�$F �H�H�E�$V 9g��?��������"�
 �H (�����?������0�t�<�?U@Z�A��^������E�'�t�� ��L:?��֝��������C�����ڞ�W�( ��~��������EAz��7�]O���A���Ca	,((?�
��a�p�����
 *ϧ�����?4?_ӼE pxq?2�_�xo�A�3������?�������DPWOxP G�
 *�@ga�����D��_�,��JS��?���ˀ�|O}�~ށ@^����ꔁ��y���W�I�_�(���̠��=��"���w��~:���!�����e5�#�Πhȅ� ?�s2}p$c��k��R��Pԍ5J*�W�Ƞ]e$GM;5ٔ���MZ���i��F��-�vҡD��kT	duԥ(QTn�#�n΄��Z�E��Mm�[v�[gswN�k+�knuֻkwvۻ��]�m����-������ڊ�������lwh�n�Ӵ�\��wc:n�&�v�ͻI�Ս��6�wj�ӫ-��:�{�k�gv��rV�uj���;Wm�w]]ݺ�[��+W'v�Z�9ڲ�t��m��k�طT��������t���cwwm�wwmp�ܵv�q˺�n�;6Uv��i���nw��v�V�k��  ���6����mp:�m���E^�޴�]5�k��]-m��u�jv�Pٛ��.��t�mhe&����շ�{9�m�i��I�z�[[V�6���JV�[Iī�z廷]�Wj�]w[w;�v��|  �c�b��
$��tС�����"E
CD��>�H��4���mLw7mV�V�qu�]�����ˮ�k��j�ٹ�T�mJ{{����]�;m׽��!m�{����[]�t�Z���[l��]ݹw9md�ۦ஝>   ���W]�쫺��UۻWM��vҞ��=�����3��7��vV�wZk֯{uv�Kn�r�T�9ֻ���mw{�Е*�fl�S,�^��km�qm�]�uٍ�e;m��=��rvk�w|  w�A*������u���u��-1H��wV��{�&��v��{�T�l^{��**��ӳ��U
��.����g[��*�kn���v��;]mں�gN�ie�n��>  �{�rj��Ow�^�kIJ��V𒊫ް�[m�*��ޞ�:���jT�ӥ���
;j��:�B�#Ӫ�k۹��Z��zЋ{׸%mE���v��M�뻵ܻ�v��   �>�����ڵ��:�Yw���4�Vz����۝�v�u�u�u:�[ t]��ݨ h�v� �� ���� �����u�c�]�jw]uc���   �}  �w�� u�L��� ���x � ��]� z�<  j0�v��{� 9�z�  ���  =��볮�����f�:���]�   ���}����o  ����  x��Pz3��@(��x  ��������x T���  �y����{����t�+�M:��Ʈ�   g��I�� �X�:�:����7��  ����  6��  )���{� ޽x页�t  ;ݴ��j�w.�U�`���Wuu3�|   #|���0  y�p�g{�  )ܺ� =v综  �  j1�:ݗ  �N� 4;o�"m���  �����4F�4Њ{&M%*���  O�JR�  �~F���TP   �)IUD  3S�_�����겟�Ѵ������آP�L��}P���yR)Iv��S�����﾿��z?�61��l m�����m�݃��lcl�m���_߿�������ziW�S��;;�2��+dp�&8Ͼ��3��w�9	"lc��{��p{Տ�e^�tr�[4�H�q�e�ј�^F!Ԯ谮j��
ڻn��T�)K�lj�S[awKp�*[V��Z�R�af),��K�ܧ��GMj%���-0�KVvKRU֓�;zC��h�hؼ�I���a��te]�ۭ߷��U7A�$봬���t�]e��iРt�/i�#��_1
�#�"m���h��m�v�F��ˎ�+�����I���x�n%�f����*��^Kǀ��@x��3y1�]=��F=쒅:Κw5�VmO���vLA�Г/�>|�Q��T޺=��'"���JͽC�
�EJ�"fFv_JzШE�N����2��і�"�踱뀵xE�-r��<TՂ0Rem�(a��0A۷�ʷu�iGG �ʦs]lcF� �1,���Eh0�K2�x�
�V�f�%6�=H�� �M!Kn�-��2��a���X��N���r=;�?lX�J����b�9��%b�逤����Ǵ���A�]�Yb��R��D4�Q���Î3r}�;�J;��˦��.�@	�����������(x�q7W(�t97E��*6�3�]�� DaJ�P-��˻n�況���{�h�;iں��Շ)* K��j�of�6K/%r�f���n�Av@AK�R�5�!(@֌���݊�QY�N�fC���Cjcf[L�%ZYv�f �c��Z�enMZnP��pކ�����E�u)�0�$TwEef�C+2�ek/.�6�ܧ�(!9Ff]m���L��V-�02u�l���Y��93,�cT�tr�֍1���ɚ6�l�I\�۩Z��L�.j��;'q���y,�e�խ��L�5��Ys�d{�;��?2L;�%���6�x�-��p�CF9�O]�LY5��F�а7���[g���#%�0�ܺPl�ׁ�&I���,��]��t7FE%�����5c�ͱ�[	���.Ȧ�	�5�݀ P��	p5YB*IY��k..�^QZ�Vnh�/;e�X3t8�u�T�b��Fr�hL��J�a��0�Z��Z�$�L��V��4c�,nݪ@��Z@�����G���N[��:��3[Wu+v�c�<4��٣1�|˻`�������d\V>A�>���kք����vu��t��
�;)���,��u��=�J�%%�d�ng.���I짱�^
8�D�h�ˏmӫ��;6�U��:{�0�4P+!Q��S̕���Pw��eH�!��R^�u�U�	G(Mr���4��W�d��N�5������*F��w�,�A��!N�-F���U�-��z�>Vx=XR̷���a^�C-�Ε[n�SWD�p�&��G����4�
 7����LCh��gƨh�7i�"(3Y1V�X�A7N[�P�@U]�Ѽ�→��]:O �[�+"�F)�a��5`�Mأ�	��@H`)\�`�{�s&�qk�dQ���vl�Tߦ��5V�gD�i�����;8c9�a*�j�YǍ�/��Y+y-Su�]X��n���	O7�u�!�ixcۻ�̭+3��N����W�P�(��%GVu��JЛlۭx���J�1kZ@#)�0��rq4H6�ؽ��2h{�^�9,���R����[���w�N�(wm��dҜśYv�'�ìK��bA]�ē���v�]�����lX$jv�:Y�����y�ɠ��K��4n�VHv�P���X�ᒞJ�PQC�9`Ū�ۧ� ӹ�,e71��hj��e�(��
��~�C.�n-2`���#DX.ї�-�bk���*M�
�a��,�v���6��$�m�ϡor2��	e�+He�7F��Ni�5� ��/2�sl20�T�0&.�ɹ[t�L�)�jw����t�����I`Lnӗf�zm�vQ���e�>����3m�H�,���,��X�5�ݝ!b�**P��nS��k����6�64�ޭˀ75�R��I(�eą�S���Xkj�#/5�i�֓|i��1X+h���1m�`Ic�X�i/E)oL�s0b����l��M�vE��8�amF �h�*�v��kI��4*�/R;r��y�u{Y�le�2�B��ܵcP�u1�����3a֭2,��32!H��}��₞� ��t�2$q�{�.MAᡏ�-��F��d���3\7v�i8�Y�����
��F�d�i���ᔪh��,����b�Cͧ��tc�5,;�Sf�/j:3�HI�ڲ�,��+���N� �T׃Pt��j����V�Y�����,j�C0d�w�Z���-�B"��K^Rd�G4�֒��ֱ�v�t����M�FѕkM���Kr�fI�|�{���V4�ԗA� ��Zdc��,�P̧��j�\��B]m	`�{Z�gX/09*\n�� ���lgD�ܭ�k���U4њ��@TY��kbV\`�y[qR��Z��[#e��Q��ڲ��]��a�Q�l�
̏3<"8����BNI��pp�sV�Nd�1�>�0�.��%x�f�R<�����*ʑJ�Yw���kDR�9�@^����O@�
R����bˇ�v�Pdki��0޴(e���"�d-��F0TCF�jZ��ݖM��КZ������*�JV����z�*E��̊��s�R��%0E�͔f�� ���[p	E��z���2*�6�=9oh�+dU.���BЅ&M����GJ�qm�	K-!����E�L}bkD{��b��K,�!.#��M�BK�/Sn2[Kf+HS�Q,�p�̡ ���^��u�����Mmˡw�iiD2Q�2�&=�+>�.Jg��[u���)�cA�Y��v��#���)�3����Ә���Vb��
6�A�
"��;�^0���܂}�v-d��H���V,�c7\��I7.��̤6��VCu7��Ǜ�4-�X5�]�!HE@QX�j,I�ա��
]ͭ��'�;R�ЉOa��3���0��wH�e�(d&�û(1��@�4f��T�A�W-��LG���7�x��RY��pnk%%��9.��6�,:8�;i�;�w%Q�ow}!�Vn�c�i��2n�F&��$��)#hmd�؝M���/ihݧ��t�����(=�'��܂=ǌ��%9��L���i6op�B���a���>z��3&��� ���{���[��Y�D�E$���/�̚VS
�wanl�Mj�m�v2*ۭ���Q(`�B��J�@ⱆ��a=Q-����ʕ�1�)j�uS�<T��z U<�(�˹�0�w�5��*4�X�7�cB���H
��
�ң#�K�4FՍ٥[����L3�m����7U��k���p���
u���O�y��)�wF�n��uf}�cd��b�S�Q-T1i��5[º���:��{�VOK�Vt��n�� ��aV��n�в�zDEI��E��KB��CCpS�5c�n��q`�qExqɔ46Ul��T/h1�-��q��֭����� �~͐�V���tv��v���GF�U��,ͩ��[�R��;n����Kl��K4�������}���3���$�'��6�ʶ��@��E%A[KrU�:���(�Ddk&KjTA�V/1P�ʧme��f�3n�[yg1;�*;V(`�-�MP6�eX����Ybҩ��ɬE��J�Cb!�M�ǎ�}��%f]�W%��:Sw��jK,�c�#հU�.$Ǫ������SOw�iу�5�f=�ގ =�M7+MV�q`	i۴]{�+�1ֶ%%�yOܤѫ�m�����c���(�ߵK��v�=�h�W[
�I@j`j�y��ԩ`A���`ay���͎�*Ƚ)�%��Y%vT�	[�Z_p� ��W^���J���;��y+ʵ �7+.� $e�!��6H�2��:������X�*��ȨC��^=��C@��I�`��(��㕅�\I)���-#	fZ�Cn^c��]�I"�l�21@�%�&����(^��7pp�ЙD�uS��pIb�38��lf���z� \����Y�cAs�Pĝ�L^� 2�Z�-8�j�D��{�K��x=���wJ�mւ"�@nnX�z�^�۴,[H!� �j}4[��O�,D�w������S �m��Ku�wSo<OS�v�j��1-�֩���P��5^�����qG�=��ׂ�P��Z�l����i����݃N4.�-�-h���g�J�� ��,��b��	R�����I��^�m�C�h�-i���!Fh�a|RH���/e
��NӦ�šSф��A�G��I�ڪ٢���{i�l�����fV��$�D�YQ��Y��c��.� ٹ-�ӬǢBu����c@�4��X���ۊ�iI���b�Qjid���w�[8~�a�����6�J"����$tɵ�GD4%n�]����W�(}�����U��Q
�A�z�r�v\�h�OYg1bW7	kp�<Z�<�]R��VK{/�\؛��g�Ã(e#��m�˴Ɠ���C�,�i�A*ti}�˨��8��SN5����ֳPV㻆�RfU��M�"YS1k����^�q�:p��Deһ�ߨ�-f�:�:h��:�d�����Ę�Z�j�t)`���VN ��gi�%W�\� ��ob�`���V�*��g#��BWf�,S��*N��E��#�����6b��JP�c?6Z��6#���튅h;�VGW�k]X�hLM�4�E��誳W��2<�NS5{�b�EIɹA��{M\53^�y�m�+K�0���BɌf�XG>-j��S)��n��@h��	�Wz��;i�lZ٪�8ڊZ��MAE�21��8�����d:�6�V���r,��[������7X�Qj�jT���v�e�*]��㕄$��I[�Yǭ[��i���f;��$6��{Wb��M"a8���
.�<��r+��)Pj��+p�iP���ܰpAwn�Wn8�:�9g<%5`Ӓv2��7�G%�K�{j(�s�{Fqf�{ɯf�S�4�;�
���e%�Ҷ0�Uu�4�ݙF櫬�)��
�5�女4m��zu�Lf��J�Ӎ�p��U��I��!��X�aʁ2�9(���24��Q)zt	K�ȍ+��F�i7jJ�T$lj|6H � x���8�I�R)��͂R�fR��y
���@���G2m��W��;T[�I�M�Y���emQm!0���]1�J'X��ꅢ��w`e�T�55R�; 	�.]���Rƍ�u��̨��E40Mŵ��7Q2�%��ֹ�f�3\���
mF�Y�E7{�X�[���<����K2��hVium��vjV�ۋ1I�
#��B�Pw�
TUs��"�DY�*�.a	=�˰��a�2��^�4U�k��Rx	nh�Q�+Z��[k)���r�F�#@j� _��z ���;R�U╒�����3M���b7Z/)'L���&c�t�Vӷ���,������ ���ef�0M�x��y��Kz��5)�����Vȯ7	B�4�$c)m���i�j0�u�m"(լ!�i݋h+C�n��?`"L�`z�+T�@��x�YCv c�&(�B�5��#�5�Y��+/q�km��Ҋ�D����Z1ܑ;p�&��Ya�݉�ê,���6�r�֛�4\�Z��нu"�m+	[Nm�&���F]��Y�A �br\<b�j��v����j�_V�`�klު�l��U<�QG����A�)�Z�U���N$�Tp'cv7wa,�
X�j*�@���͆��A4�T���:�HA�=�ȕ�zW4�X	���hm)����5�������#�鏘P���E;�B��bd����Ms@�i���ޡ�H���Q�[-e���-�N��ب��e����Z�=&x ��Lx��ڷZ�V�E���5��vf;���K�n�ح8�LkYA�m#R�v0H�dP�&�8!�i�^=����Z,TrZ�-9�m�fcЩ=mӌ^ˬ��M[y#Lނ��?'xcr��v%��W�~�Cשh4cb��#������g	�ǤO�d�dLil��Ya�����t��|۲uon�7x2��̨vu&9h�L#@�x���&�);,�j�@�g*G�6�f@�5�IY)<�W�0V:��GM駜�H�S=�i���#��sL�e��C�S���KG�[E�
pH\��ER�-�#G#�y�m�u�L����dE�ղ�!4��ٰ�.�h�uo0��Lm�"�͢>��`����U3�ŕX����f���֐��w���lr�+�V�@���=e�j�sq�.#�BƇ1Pjgot�XݲWLJ�`�'�j7)��i�tG�6$c�k]�.=�6�\L����*��xq���"�۹{H�LPe������SZ� V��-T�wq�[�rY��-�o"e���	�f���.�j8b!P�u�n�⬩)��zhJ0<;&m�q\z0j=VR����Ֆ�ٚ!��Yq*ØVm�µ�{PI�10�e��E��1d暴J]6��C6��w�ճh��Z���g�uyskA��z����:��ȧb:��e�(�巭�����U<̽���j��І�Y�0�=`�}x�]���	��EP��e�v?^��ڏ˙��%� �)��j�+��H���6$�qܧy�9��ҏQ?\��u�#���1o�g�SK����K���ڲ�~I�C�d�k2J�L}A�6^[ދ�o��<`+M�[ړi_�T��!SUZ��W��t����w'�tP����JU�n�"P�p4�y�k/Y���n�\f�#m�Ptf�xZ�	p��/�X��l���5c�3��L���F��S�u��L��%�U�{|,j�t�|�u���׆��X�>��lL8�fR�Q�7y�\�c����Y�%}�D��E���^!~+��j7��l��l���Vܥ�]��kc�Ȼ8��t#^4��$!H�k'w&S����2��"�+ڜ�_�s��z��Q���Iއ�}�n��3�Z[�sP���4���v1�Z���d�)����0J�D��׹}���CC�1���o8lM;լ�b�h�|VD5�Ѓ���3�S8�MJo�]�¸s�:�_�d;{�F&2j��o1 �(@75�w^��*j��*�M�x�`�#�%gӮ��e �o�h��CuqݨA����ū9R�%�%-���7�M�Ύ�mh-������Ă�bcM�����@�0[��P�Ԥv�b]����--ƹ�2��%�h�z�B�V8}����A�M;���k �X�S${Plk�/O,W�^����Y%��]ä��,�:�V��1iJwݱ��df����s�6`1�׋֦}���f���]���VrL���e����!��;bi�w(oE��%���+�iQ��i{]i��I�g?���Ds��o�_U�����Gw�
ɑ2o���h�ˎ���ER�	�MdaO�w��I�r`9]�n�ƍ�B\d�/2��h�y:A%��9M���.l	w�3(t�Qݎ	UJs
!}�����4�9d�k��?ʘ�PǶV#��=��6=��v��-QY0s'|r� �KJ��-(���f'��u��z�-�|*0�ժ���^�ܓӻC�[*���Vx�7�*G�V��]�0�H��d�Еɺu��&ڌ���^.�e��ME�Q���k�>8�<:� [{�yb��6�9)t��l s4�JH��;��{)a���
�����Z�[����g&0v�E�E���٣JA�k1�J7ʡ�=z2o*��}�.����|c�˔�Ӿ~��Vj�5��
`�^Y��KNa�nXeZz�o��tX��Kd��Y��T�F�n�#�(�jw�7�+r��n�3���b�-�^����z�nU��lu��9�#������<f�Z�߯y��]��l99eu%�+d��ՖE�rnh�*|�Z���原(�T��7f��<�!�}�Uq���5W�y�l�]���.�J�Es���!�V@Ѻ[7�d1A�d��r�s�(XH�C�=�kH�%�k�e����F*���k֪V�t�Sg�B�B�n�����un�z�T�k���˓h�+S�5@J���r��q֬stwZ֕ҝ���FPe�>x�'�`�X;�|Ƨ�/Kam`�+�<�[Q]��C�K�E��M�;R���U+ڢ6���Z��T��U�3���blY�#/��m�)�F�`s�pu�c����E>`��9X�LoRqE����n��]%Qv����%&��mWsxy9��n���ꫠ��w�9ZDJ*#��M,�[m鄡x��5bu����a���5"Qn�Ch�*�-Вz/)�=��3����8r�p�\�&��b+g�aIAb��1��963$��F�\L�ZR�+v��F�7��"�����}g����f���L�Ơ-hT��,6��C8�5Y�����_+o�;z�G�{t�|��q;�b����� ]ŉ6D)�.�j*�#n��u��ն=�������*
�
9�֚�����ɝӭ&�^���+	\��פ�����d���>�|�lʃ�Mc��1�B.J4I�<~њ�@mD���K��V�h�Ybc��+:w���,n$����n�֌�+�����6��j��i��I�����Tڵ��8w$�k��=Xh�*h�d?�~�P÷�d]�>}�� �*�)�΍@���m4Z���^��O-T�.T/�iډ��ұ��^�{1��wW��m�6A��?E��r��3ڃd)����w���A�u!�t㹳��-}*Se#!ubpf�m<� �N�	r�������v�E&i�s�.tNך�nF����}���.I�U�h����-���hR�qX��Z	�
�v�ޘ��k5vR�AͬU˶{^����.��1���]��즹��W���ym�g��h�`܊�Ŕv"��CEI5�N��M�t��c5��X��t9+�<h�%(�w�iǚ�UHoM�{6�CX���)OZ�M}�r�t���tc�Fn"�l�n�<[9����Fr;}�gb��칬�a��e�V�5і��㦃��1Y-5{��<L��nY���#��9�g2}�_m�� Ѷ���o~�j��3�S�;ڜ��bu�]�!U��tk3"K��|��-�[�N�j��M��m�L:H0��V��?JV�7�2ESJ�I���1t����B{g>�x� ��?.F�e�+��Oc��5�xzp��n�b�U嗋q��] �RxҬm_[��*,�Ia�Ԏ|xf��l���yf�\!�뭫���;��嫃���/[�+�f�i�y
�p��y6n��ݝk�@Tt9�ԣ+y��L�z�wHQ'k8���&Y{����T���Td�hT�s/���gw�AꙈ���/Q����ަ��i]�x�F�F���g2wI�5�f�2)ܰ����/c���x#�pQ7��۷X��Q�V�Q�GK���������(���2A�e]��~��� $tf�T�TՊ�vT�6�$a��Ifp�v��6����©���{�T[}XN,��.�k�vD��C�d�p�1��'~9O��Hf�A�@:�%3@af���E7�����8���k7'�P��B5v�8�IZ/p�T�E�A��cQ�4���͞^�GEu��,��8�=��n��=��=�>:{+-�d�$��lN1�t��v�5��gG�Ó#B�WrT�f�2^T�#!^��2��[V0]�����42����,d���Kݾ#�<%���)�}w.�\.��Bnr�\^��E[�r�X=m�S4ٕ�pv�;��7�����w\��Z�|�,I�Z�Z*8��,�����ֹ�xZ�4��n�Ά����l*�׭�ق��vn`�mݙ�i� ���!�aiê��f���=�X���
�'RPؽ�+e�Y���ڈKp$r<���^���� %�b�ώ�o3��f���f��E H~�}�,�-��#X��r�Թ��&���"�qN�����7�_�b�f�A5`�}Q��!k0�{�p'"R�pl#N^���oNI|��K;4-cOa|b���Y����j��na�Z���V6n���7����)&�
�{
�f�{��
h4��K�X��N���f<_02�j�ءOr_�ᙁ-��'�]wDv�v�H�Xw�^%�g�ŲT�S��8���dZ��6;e=U9v�ŀ
=w��$�<ט.�,���N�dH�kR����*�gR|ӧ���!����ץ�ٝ�7���oNIK�խ����9{)Yy{�͔��;U1�R�I�3�m�b]��s���v���M:&`U��iwm�*�ft�|����b�c���B)��#�2�f�Δ�����o6 ���x�}{�,1���B��#�7" �ƞ�9fr#���}��&N�R���4f���N����h͖� ul7fӉq�𡺷w���W��5��k��ϳ�s�xK�ˉ�����p���d��=� 9ն�u�pu�F��`���;]�)J:N�	�$�ܜ�p֤3D�pu�@㘘ks�ia�z� TEe��Q������q�L�}8n]�]�d��q�_�fԹZ݄�ٟn쓨�y�J۫�!��mBD݈���	!��-���zJ	�5uf�(f__o/�;:���Ҋ��И�\���-n������E�6+:F����枵8��#�A��ӈ�d�Qo`C+pF%����i)�T��L�z�u-}��.(�@t�'7�e�8�y�%k���f��Ť��_;,rk�Ops�Hm+Wt7yظ�Y�� �4`�M��Z)�m��+r�K�AD���&a����Ǵ�Hxz�����{�-w�q�K�D��^6����ލ�Ŏx"��}�P��Ոk���|�3��t��r�Rծ$�ʔ��$�]��%k�WX�J��3�؉/.�,[�*f�@�`D���ry��*q<�e�l����dhrǽ��CCNS��7R1��(J�L�˃�"�7Vl�X���y?)�2�E�)u?c�t&Iz���a��g�/ezqR�8��$b��-���rɇVpڗ���J�xS���p�RXe�e]m�8hHz�=��m"�m�ao ��8gj=�N4�%f�ÍHK^���]o1���2FN��἖8��¼jdvn6����^��g�m׍dUc"N�4�wS��|��Ƚ���]���[7���aj��k�%�ML�@߸j~�#Q�i�#��ިxt�Ņ}���ZvQ�a�gY�Q047��oD׹O��t���ɴvF����9+Z����h��E˓WJ1����*����6,��nQ�ɵ$��:���*N��_*ɵD�-m���j�4,�Э�u�nȖ0�e�S��Jl�5��4w�<�vL��}r�Jl	�$�ʹ������o.^~�ʾe�у����Kġ;.'��2�e�E�X;�uty��2�c����;�N��7R=�ڳ�F�px�nR�M=��T� �#�v���R.'0.gpx���7o�	|��Ӭ���g����4�Z��A��k�]�Tb��V���o�dwizC�b����}P_V��(���S�i�a�ʁQ��.���q��k�N�uJ�� ���)�lOLï�B��nխy���D�7��"���Tp��+��ۺ�6�:I�[���Lx�x�j�G
��+i�WyA}�z`��/�-�.	oHy�G	�ǟ�F��d�-�8��紞�$N�f՜Tie�I깪c,�W4������uG&�+�)�e�/�>�ӽa��O�-�~���#� L)�<Z�a8������;����7ݬ��r��#}�y=�N����t0�ь��1:޶�֮㶦���Ud����S����i�(�g��\�=�-h��m�;��*���7u�A��7��P�%e�N$+�bޅ�#R����P˷�-����Y܊���5�R�S,�Mut�~˘7��}*��,��M����^.�5()ݐmt��O��']jK�&嚎�.��ٯ���;J�Ywc4Iϻ�z�c�*
S���gm���]D�M��Zvd�y�
����d����h����
[S�:�c�T��xɥ�]3B����}|_E�r}�3�Y��A��}Y%�"tSq=U
yQ��^t��f�5�6D��^�HăD��n��,�SF�m{;@��}�-���-)�&��; ���7Gt�R~i�Y�+&���zf���32����ӹ��P�H�ӧкJU�0�4	��⃝�K$�*�*T��+�8b�fF�z�J�L����&��=�6v�J#N,�+S�^[1a#7�����l�#������f���	�#��fA`�-���ʝv��Amm��XF��*�ܺ�:�|V�5���	m��}ZZW�J�>搻���E13e�C̮Yy�e=������w��6�K!�� 9��يq���>q��b�ß������n�x��lCj�GoS��͘��k1�Ԋ�M�yk�~�:Fa9�PŌ٤T߶�嚝8�Nz��'jt�X�8��,��党���	SauV'�d��	6#��w��2z����Pw+��'�ح��b�t^
�:�0�(�ڱ��F��_ R;Z6��=uy������ֶ����7��Yi����b�-I�ԋ+��p$ΔD�T��Y�.c�.�\��}I�
�[�uJG+�~[�9�NPB�uM�a�]��tb,��e$��3e���6^�i�k�������.��Þ���=��p�i�Tsc�a���Xwzh�]��D<�&���ς��7"���C19���6��۷ۊ�8��仔
r{���̱:�9[�a��e��:�gR���/�ŵ�i���-.�}w���o�f�{ٯ.:	$Kv��������1�� ��zM�ԻNQQ��l��Qb��9[���u��uuF�����F;Y`�	\Zŏ����i;%A��j�SA;Z���qx+Ckkf�@�Fm�q��{�K��uM�z��f��8��#�뫤'�,����+��M�g�qw��&|�jG��3'Zb�eX���e>�#!��Vp
	u�ss�6�vD�LɄu
0�L.�|ﱪ�R��xO+�c���,`vw.�>sF�u��A��r��Ϳ���t� ���d�_94P�%`��'iN���^�/�\�$�t#}G�/�ܴ�ʴ/������/���lĬ,��c���!"���::«L��N"ˑ�NѮ��������4;UL+�tY����(f�<�e��l�:(4L�+b<����J�y09���r�ˍ�-��X6�l��jU�oN9����^�=u4�ݼ��s�$8��tG�&�/���A|&h��\sB�r��y8��n�,a��T�-E�z�v����|�D��}����������7��o7�냚�K������w)��� ˜Z7S�����4â��{������/r~�^�X� c�`���@��@��lJ�KUx��Ke�ZW&�*�1��uݥƀ^�-�=��]��X�M-�vˤ�-n])�:Bk_�v���)���p �Ȁ�cr�f�ېS�C��πj��w`�[JXjN�ա)e��ʫ���a�ѵ�}Y���
��l����ߝ��s=�;Vn�}�\F�kT[��~��M�/)8�u�i\2�t��T3�U��*�x1R���h^��yls��s��Y��+s\�3��b��Of�H�jI�����įo�+��׵��ę|5�<��� ͸/unRPwWn�r�����6��3s{������0����!fS��iF��-t��(�ryc�4���n}�M����e�������*�;E[��[6��d9x�2�ۥe�q�|�eLZ)S��*
�[�Vr�+4�|��n���ls�*$zQc'`�u��^):�4S���:���r,v��
e��w�s�^�ɖ��ʇ85���ևj=�\��5��d;�-<�ҋf�:Ȫ�b�CHf��c���[�s۠�+'L�<�ͷ�+������#�av��Z��h�:g������A�Y������-O�B�*2��9�e�U|(��㧞�lK��3wV��_hZ�.#���I��5��L�!=������3>����[�SZ n6Z	��O����3Jm�yp�:�WX2�quU����Ef>t%LW�����T��cJ�јE�Y�c˸��>'�gP�ɏk�s��U�7S�c�Y��W�nh�wݒSV��������&ڥ��!�>��oeK���ūq<&�4)�_<�3+���W|���x�Ȯ�Z�����l|���fG��u�E�=�-rO�h#(f]�]�'�I�ν9]�0F�z{���f�B�N�̗a���Wɜ�e��W&]�;a�%j��A���;�����K%�v�l�j�G.L1P���[�gh#D+Pa�N��0�}��~$��3��mTy�y�fkAf�г\T�~bJ �g�w�v���Zu���w��Bu�q�v��QU�eǇQEٮ�������>��R��Y�-/([8bհb�j���:��'f�DV^C���#Z��)_d)��ڥi,Ld��2� ���3I�w��p�ջ�F��T�eOj<zq-fռ��n�Ķ �9�!�+�U̨!Y��i����XwK�;��6�ȉ�����Ly���h?����iKu�<��za֫a<����^�[�=K3�H�:������<70s�W��|�&{�S0�7�b�� �t\���wN��9��i'�Zb=�WE��^�c!�^���ie�<"�����fz��F����3 �ҫ ��(8l�&�k�;�����Y+q�B�����skv\�T��Q�y���j��-��x�i]��.����Kr����v^�F���;ɻ���x�Yk��t�YWY��JR`��<��b*�ݭ�`�Ĳ�&Yރۜ�Mt�y�[8{a� {�V1&L��;��0L�ͣ�6\K�϶v���=Y��H.�P>��6Z���Td���]�1-�I�ykq5cT/&�p�'-0P�Dd�s�㻂	Ć�]���s~�E�ѕ5uX4v�c�;M&�W���0º�x����k���U���n�5����.H4E����S��1,�l����9�Z�Om������l���qs��l�W]m�\欫��j�z�3O�3`S>���a�{7S�F�wP�����P������͉���ר�`��?]�a��ɻ�f:	��N�/i"�>p�22����b�뚺�糖g��Rw&O�l�5�t���x*�#�B)�۝�Yt�хb�i��Z��ø��,�ev\�k+k4XQ�w����[X�u�ո��c�a�ģ�򢭳+!ËCdp/��T�f��zu-�{�����������>"�*�~�d�*�N��[�w���WV:*EY�f�R��I9É��G�ے�w2.Z�"df�)gDS6ԫ�uV�s�s�q�Ιq���/(C�ѣ��9";�s����7����I��X���7#�\��;��y-gUIe��\ۦzw��Y�ْ�@ʥ.�U����S�f�ܖI�?J3tݜ�4���K;><B[Y�"'�����_,�i��Fnmc�2
r���N� ���J�?����3�8&�-hI5�\3�=Q�ݣ!����al+�w"�]pյ`����ݎ;f�W�f7H����Y��Hh���l�Z��|,Β��\q�<J��y[L��!�{W˧6��1�[}�2�R��`v����EVSTZ��-L������y'Z�3���-<��8�坢!�!;kNvu���*r��'r�{��xu�q�fL>�,�{�~��8�3r�el���x���C�lxe�G^B�e�s
�u��2j��
�1D8����ty�Zk:�6J�ub�l;�v���0�Z�љ��Q�FT�Ï~LN�5��(T�@���еP0m�vVR�(�V�Z �ឫ	�z33�3�́�LS�s��{tI�kUU5�k@�'E��v%e������~�I�U��q���|�����d\���,�O`����OkX��{����>�Osܺ1��|z黒p`��yl�hԫ��V�J��������G���k��ޓy�-i��z��.��
���wP��?mY�ɖS�q��>�|�2+�zi7�:�NA+ȊZ�5 t6����4	���bƍ%)��n �>��b� �-ΰ�S����C��iͮ�HV3�n��Ϩ��W�)x�;�Q\��s�Jg8�^uU�L�c�Y7B�Z���ϝ[�d��:�A��8�c5�p��Mlv����wTͬ׵�}n}|h�'��p��p�A�g5Q��I����kw�����$x��_����)
��rH!����L��&���Bƍ�W��{�����:1z��.�5eJ��4��k��Fވ�o۝&]�	5y�4��NY{����$�gj�� 7����I6�ã�ށ�1U����Nv��k�:h;�!�-Q\�q�M�n��1$/�i8ddN�ڳ��Q�5���m <y`�̭a�ɚ�d-�:-W!N���㒪-��,כ�T.�F]�sn���z��!MR�)��R(�ڽ������yݖ���6hu��^,w�"��̮3*Ⱥ�x�EnŬ���#���z��g���}qX�O��
����_Ky[�7�+�l��v�춢���,7����-k�}N�j�Y �\�5��P6�S�S8\lK�.c�����0�i�HZd�����0��|�7�����YeCC��,���Vr�K��u9m���)��v��Q����YeL�X�-���J4����^*6��/9�2@�z!�2�݄�"O�u��;C��o,�����-[ <�LU����D�+yu)gN����m+�yņ��,�>��RB���t��p��D��Z�0I�b&W>o�]g:�B>9k:����b��U0 �Md�t��j3���'I$���_�Ug��CN.xiӍ�:��m�*�oE�����ݔ�L���)pSQ}�
<�8l�[��-x�a2�ɝȈW"F������"�q˨�^�j�7G�N�v�W�јo��� �
U4�%�Y�J�	��|w��D�I��d.V�K��t۸�w˪$��"J�X�����K���
�X�C�e�3�JlS����'�Xev	��� ��[¥ΠM�U�]f=�Q<c��D�jh6*>�l�s7��ղ�Lz�P�%���*wV�[U1tO4>ZE�l�F���u�ڮ���\zM�)ڎa�IW��6+��/xIl>d�38�Drו$�3p�H���k���و�yV����<�>����"�X:^��gf��%�D�����Lx�����m�|��ɯ�m=�xa�,$y��lPeȪ�&ċћJ�_hxgZsrˤQ��2�7uP�	Z so*GX����X��=geF�Z܊�F
���66Y�u!��ّ�S�2N�i�����M�[�������B������f"���R�ǅT����{P+�wX���v�E�ϧ��uu�ps�"�9������H,�&���mh!nÄZ��F�8�[�l���=x-�n3"&pP2��9\�o*�e<�<Z��S	��Ȑ����I/I~�b��gp�L�����o5}%\�N�X��NS����R�2�v���J*+"���zJ\潰�.����e�㯅K���@�0d�x4>�D�8�WG5DOb])�'R@�жr�o�t��)�OA�����wN�cPK�lб:�a�xyAQ��X��uH�r�9T(V᎚P���gk�5�/�`*�=Vn�-�&N���G H&e�kaI�ۗ�WsKx����ӌ.�-oT;�,�Ēb����t��- ���r�V��A��cz�yt��8��k��̱�L�y���/R�ŽS+��VGmF�T����W�����VP4��Q���ج.ԫ<I���}V��I��y6�]A�O(���$b�a�۶禄��"c�n�[zc�F����om=��?6O83"=W�7ۡ�,��St�Tգ��"�<�e�#i�� �Ֆ�������V�5��ɟ	���P��'�ќ��X��J�E�����S0�u�_j١�ճ���8��D��W!ŋ�iʛ�N)�j��n7���A�/aj՜�[���eԱݧ"(�kQm���<�B����V��V���j'h�x#��,�7�(e��4�#7�7c#�zmۖ}�+��Y�W�܁vv�[4�\��8��\���d��(�3"4��x{�R-(НNoL�Ku�9���f��)�+��Z�O�{D�Y�:Z=�FT-w\��R��ɱd�qx��]+�������O9��h����i�^� �n�������Ʃ�"/���K�G�Mz���Y�]5�Lٷo3y��4��.5(5i�(te+�N(᮷�0`��oة2�^(АtK1=��������#���
���#���fvr�z��z����<�a�����c1p�����sm� h�yX�o����%=�nx����9�fH���D�1�B�|� 4������?�U��Zm�ڌ���2��6�c��gv�P������� ����ER���-��8�|�N����#4�i�Y��^��B���|P���yf}���t#.|��-�]։�&�*K]�	O�I���W��zi̢�2@��OÝ��/_����5�bg+�h�m�8�Y�ْ��a��� �'�8~EXyj��L�ǝ�������`�[�杊b����S��<���p��ac2��%9���cT�0ˬ|j_=��o(^D�*�T@/��>Kmn'a�	�ΒN�x�@�L�����G-�����ot��t<{�YH\�r�e3����p��:��WbC�T�X��>�j��6��o�6&���Dkl�58�kй���@rv�����*W�wݪ��7��N9��qu�2�I��U�yb+G��G��uơ}{O��VK@�d���ź�r�ܘt]�k��<V[�'VQWocFˊ��������vL.�k98�0i3snZ�i^P�.4��Hf�lw];*K�.�N��=�����p2+G����]�Hr�>g+)�֚)�˭K
dJ�p���&o
��]�#�8��t�����z�e�J�R/��ٴe���-�b&�ӭw�g���:���[���m�[�Ө���ݴ2QÆD����he|��<�7cp�#��~���/q֧��n��+��5P���.��t��r5qn��w��W��e�%�y,�ъ7b�^��z��o�)���1(�����M�Mք=�fd�y�ԩ��A��L��y�n����Re>*%C
n2��e��B��}]s'/%���9��v�[���86쮐-)�4�1�aX�JA%��;Bڇyn����.�[������K��`|٘�4N��U�^��d�j���a�k��l:OE�Iq�ub�y���s��V���-:
���iֲ�Ğ�%�,fK�Y�ګ���hl��J|�����U�YS}�-^�ǟ�\���!�{݌��M�≋��U��h���Ph�E��:q��;u�
�`��������;΃�4��`�:Ŵlُn��<���[���5pW�eb�m�7/���{�B�=��j`�^�a9Ķ�KwUm�N���st��q�!�ъ
�_�R|`����,���w٧1��GeA�������O�DX�f쮗��A�5�`cRe�a�z����m����w���[��H�%��8/!��1�����߶7��3���I��;r�����ҁ2e�M�M٨?��5#,.s����s�J�^�s�hv��:�|2I���ڜ��ɕ�{j�4t���d6��2�	佰#�p��囗D�1��9sNd@�u��(�ƴ��r�D�R�].ߦ��N�8���)>�X��J�*��H��<vb��uj�*=��e�[Z��G�u��x �Z�/��L5fmI|v�=r�̃�dΒ���P!�@�:7�oj8�Lи��N0[�[Z�u�Nfn����9FU�4����7q@9@rz�S�sEՕD��s�u`����䞈�iw��t������N�4���@�p��eJ)�]���r�� 1Vj����vV��V_)����{�O^�%�n�cۗ�G3L'�y�3�	� ��v�|���ح���M���o�Ai]����gmb�Ռ�IN���7��o{���N�:��^[FkhI-�b���Ҙ/|��^��=�ў)����ojk��}������+�
u������I6��N���J݃��M�>�%2q�x�*�.���;wQ��R0w?�j�O�_������Y�.��a�u��*\�;-d���_M!V"v�	�6�i�(d��v�F�Ե»+U��d�llѷ��F�e�y���IQ��l%��<���K��̂�ז�^���C���E�Յu��C �	yb�-g�U6 �֢���{V�W�4��a��r]雮Ļ]oh�fWY�Ыq�����k�3�ґ
d�V0o���{�R�뱳��.��X�E�=÷ne���bFkQˈu�	m-K�����5Ӱ�=RsyR�h�3�6
/+W]q4y�Z��sG|�U����S��ulƈ����8�N�7�fΓ.�)��������'�N�U�I�W�L�y�@�Y�^�#�V���,��!:��X�y'���|�Ca�ٿ�h�U�]w�Ĝ��AP�!tS��A��1�`\E�#Y���%2�6.XR�M��V�&�P�QVo6���I��۽����y��T�s'e4IӖ��m-�b�0^C�c�sFj\:S�qԢ�눫d�o�.D�`��+���a0�p�J�0�O6�����ۧ�qՍ+�65�.;*�vv���l�>R�K-��P��'�R(�RU�TIh��H4��#Kj�f�ݺ����J�D��uʸrJ�(��g)Y�%Y%��H�K�9�6BrR+V��5�r��WS��S
 ��fE�jG(�P�0��2��Ur�J�������\(�����4�����Δ*��i�U�Z�r�0�"��M�)u�,H��\�)QW�Ug��L�����"�3dS*(�W-T4� ����
.���*�Ӧa�-�IZ���W.VIW*��r��j�-E�qG:N����QYĂ#TӥQ�ɥ��8Q�KK"�QUdRETQ��2��(DA��2#����\�"���f���"�E'D��1 ��QÜ9(�dUf˦UQE�J�*4HTH�/R�s�"���$I}��H[z���&��>��J��l��hRc���6/1e>!�z�����Cy��Lwe�4�![]'AS9f��a���vw��K������n�Q�D���Lj�oh�����Fك��M^����:���ᳮmnPGL8�|\C�`��>�e ��Yu��V�2��n��u����k�B�\v&�΃�0����M���< �{͌�!���[������`��%<\Ԗ�IA�j�(/Go톦ߦ�=U���k�7���U�@��| �Cg��^�:���]��C6g.�>�F �3.ܙ^�ī�}���Q(�i���H�=������hu��,�ޡ(��	�g�S��C��/����};(rU~2����Sڰ��'�f�sW��"ߤ�i�D����0W���o��� �����X��ƺ��j�U�������^2v��Y��be_>D�o�1|Ez� �>9 %�;b�p�������a�y)l!��/{㓯>:d�joJ����.��\�	�u�z��+�O��vOvm����U��AHL��_%#L��������\eWo4Q0-@}�H�*'��M�dO���������%Ii�L`�ΩJ�*��p�(E�[�����L{����wz��/�{�B��#��^E��ΫU�P�i�c��N}��]����!��	|h��r����5P�bkLt��]�l�%	.�ʲ���y��sx��FsU{�����ŒZ�8Jyǻ+ۙ^c����Se���Z���00f��,T�vTϗ0�1Ǉ�:�W���t���l�ز?K.��);�
��S8D4�(�/^2v�LE���䜄�{}t���/�e��3�{�n��������NF�u���`?�U�Щ�����R��;?LZ�(�R�����G.�����%߽�f�hCç�P���W���j.�^���
�Ԏ�J> �-��]�8w��~3�>�%�b�PQw�����0����9�O5����D(�e�>x��
n�s�y�H���"�=�^�(�W{�	��z��O;f&��m;��s��O_����6�Q��rjYSf��^�@K//P;u=lm�1��!T���"��*�y��֥:��T*ou���Y���p�{n���:�*�;u�]=7=�x�x۷}-�g��zQ�P6>���5�k��v����\�.X�#�����*����x�fν���������/�o8��GΆGu�ժ���e������� m�(�=~����Ԅ�ʉ"@z(�
dk�A⏙���[EE�v����n��ά�2s��Du��42E�m�y�t/��zu��屻e:�9����͚GJ��=���y�;/K6������v?H�5BF�����;S2r����a\�����#o/����e�^�bB����}G�V��1`V�{R�ǵ;N�L�z��C��W��1Ag�}��:. L��!�AvN]Hk�e��ɜ��~��RZ�'o��i��S7Ş�t�[[�I�h�ֆ�ɽ�x�.����aT�e�.�n���zʱ Yfma�Ќ�L�
�&��q���"�=4�"b�B�}jY��2�u�3��e��g�3�6��dѻۢ|�h�x��=�Wy`��]SJ�J	�bq������j��@��N�X�)�-WN~lY�K�_��oႪs����`�.��53�V���Զ�v�����WOla��}�yQ�c�u�my_j ���A���*��7��gr�'��Þ���+�����f+��}�M���hK���ܩ�����XHhv��r͘�fZ`U
�R�����,O��m"-�D6�'@R w�b�З�ۤ(��	��k6v��H�����y�9Eʕ���VH���@_���)�=AQث�K[K1R��Uʑ�nU�K�8��i�Uv�O�;��j�����|�#^���0�c���6�!�h�2��^]�E�E����<��;Z7�������6������6�v*89kSi�%�y'������k��nK�����a�V��&�R�H`�n�q�R��r��Q��gĞ�Mޜ�
U7]`�awF�b�?�l�hX�G�~���\W�
)�	&�C���[�{�Au�W��K�r�5x�|<<+�u��
(��WY<ǊJZxг3.gq*˂�x{���D�O�5ϧ��)t<�Fꮏ��5��:�3�����8�!ؽ$��m�j�3���v/V�S�[wU�ח]4=W�K������s����#f�M��室;���عfVn[*6'4;�3��2S)�f��t<��u=�iܥ�t5}�1将Ӿ^��7����aD�j�S;�%�\c�b�!�`�A@�O�l�n����Ⴛ���	��yn熬��P,O�x]<LS^C�]V&=/z�ڧ�Ǐ��},R�J;=��H���.oۣӸ����ʈ�(n���-��o��
�X��^y�T�.��_ORV�i��˅t�~d{<v[5`؃~�ɀKW]hc	��H��3Y3N�F)+Ҡ��^�"j�
>~�q���g<��XՈ��* ND@/�`���P�������}��aU�VMx��I���f��\�W�[}A��!U����'QM���Z-���
T��1�S/��Nv�߭��yԩk�.���}l�X��Ѯjy��gW=�I�ՈH�/g)��X�Ӕ�c��[/2���F.z&5�q�N�߫�2:�������SY�SD�ǇcnA�B/�k�t��I�{�U�/�k�U����ĳQ�uFM���,�Cc���-L��	zc30E���b���X����7���=@��5�
��xG���-�Z����A���*�K(�M6����ɻ�y�ϣm	3��������&�k�^tb�T�
�N����|3-�ZO=�>��4�@{���Z��7Uh��G��n��N�p��\3dv���J�2�;��+w����`��@����cG����^E�_D4����Hwբ!�
믬�x�:���پ
G����IU��wP-ӻ��%2�X��S��_�N[��M��4�h+*��vK�8n/t��:,l�}�����E]��o��o��S5��Ua�� M[��VB�<���({��ƽO%�V�C��<X3�f����T{1��Of�:���n_!�g{��Ȋ}���פ}yDgz�:U
�>�xW7�<��\b�L�̵���̌q����8���`Z���J�D��iR�� u�*P~���0f��r���A�G'u���ڕh.kw3,�Niu.�Mka��}݄6fj=R�>��tx�(Z�%[umoPKT�B�g4��n�b��̗��:����9���ڽľ]��4�,e����`ۮG�����X0�ϐ���
_g �'d�/�\�0�%%�����m��b�6{_�=�lL�|��t��/��kб]Bqb^	���+�#���wr�pP������Z��nR�:r�j?.�&�2:릐��:��[�J j��97����Xm�_h&v��չ������_%�4�����#�8f<����>PA��Sx�%2w�y�l{�(j��$C�N1�����D��00���*Y;*��� Z�ԅ���FJ�q�8w��5����U	ƶ��p�}/��|��k`y{k���r˵��y4����Cяv(`���g&��� ����X51�[� _o�K�+�������>7�*6w���>M]@8������y|�=��
>փQt:�����N,a�
t�Ţ���"�@^H�p�źJ�X��߁����U��t }�ؼ��C��R�ˋ���J����l}-g��|�ٮ�uR/x�o���x�������3Kƶ��1}�����������ef�Zg`K6���E]-����u�+>r�Ff_����e��<�E�����QB0!���Lug�1i)5vxj#z����^S�$�S'5}�6 �4kȫe D�B>ټ)��ozv�����X�^ e����}�~�V,ԣ{˕�Z��C�V5���42&[f��Vc�	�P��V���P�򩎺��������z3����UyR��
D��J��NfܳT���*{]��5(d�+�SN�1i�-v��/paFd����i �^+d@�qO�ga�y��,p�s�Z��\��G�䫀�9��@+��*�G%�]��������3*y�d�>t0���j�`uH��K�?w���&��q9܇��>���6\8]K�|=n�S�|�~zo����Wr�tn/=�tTu�����5^�t���ֹ�ؓ�1`�S9M���5�:C��G�A��w0-c�zݚ�yٹPa&^�d���x�յ���K�{{Kpײ|yk_g�e�6�!��J���J����pg��=t|{���k�6�KÎG��bx+J=���>��L�ǟ�R�t2R4�m��="QFX+l�5{��vB,Վ㈝�PC�tҮ%U���&��"��je��E�h��U�g �[��r��+l!��/*�����u��U9�U(*=����6��Z-�M��W};6��Uw��ڎ�A�b��t�Ռv�{��$�"�D�R�3+s���CN��N曺J�W#:j��^N{�ރ쮑xN�2�8�������^�z�ww�f<�\�-����[��V�p�M^�W]q{�\�7�[�"��,��wpy8�|��I�{���>�D^ד�����D���G��uCWx�t>�yk�w�m��%$4�ey2��B�F;"-FM��$�]z݊O�T�������	����}����p�s�n�xN#q��!��1;H��mvO^Q�6�N;�ShK�����c,\jU�#Ջ��ˑG��W���O|"�1�a����Ds�4�jN�͊��kb��;�Șh��_)@i�z�.��g#{�W6Э�P�[5��(V%ؽR�'�ݪ���DK2P����E��a旳���a�N���ǳՎ��fYE�;젥��-Y����7�y�^�7�릾�c��PQ�(pCV-�z��η�
R�y`0��]?i�����"ݺ�1�6�I��ʬ"��P!͊Zeݓթ���귊���6��V��\2�'F���^�Q�������R�ʋ�0���
A(��ئ�]<�kzmY1��-�]]3�7/c��/�LFǾq�Ԅ��8��^�Z{:x~���DS�|�(H+M���s���?.��GU�ǥX��9�&)
t_*dL�Á�͗�1�+����J�ڽs�w�Q]�ě;W���(4�Ir7.'3��n����X
�3��	R�fؽF����;�>��8���H�+{%�4�5gnA!q��:P�`̜�����d�3w�W~��]�𷉊k��/�[�@D�ʫ&z{"����Lp؅��k��{�F)Y������+��*�������v �Y�a��.����"{=B#�)�\�zL��o���}Y���p���/���ʰట\��=h���'}{y縦�ja�7���AG��dM7�	�������T ��# _�xw}���.oU���S�;p��Й�	#lQ0�΋���,�Rz����
u���䀄�{�U�W	���d�9'=�5ut���S�6�E��4Hk��X-(lv�jZ2�U!7�wr郷/�L�|rF���-����*�s
�]�\N�}'�,�4gz@c2J��#ȼ�[�M�TfL���w�S�F����m�Q:Ǡm�����/-����@I�X��<o��iE��+n�̻������ٖ��ƚ>�P3��7�5�p��[�u���)8�%�5q�K�G\�b�]��4�+�cl���U<�Ⱦk����z�J������/u%��e2��2� ��Գ9#ir�>բ��mke.�|]��Y�z]f�5�oӤ䅎6�m��PS}��^-C���vj�܋��/S��rFQ�yu�vM��mV`}�@~�Lݾ.��Xc��r�ݯm�����D^EP�X�GY��6�r��\��s��1��Cʺ�����܁�5.��wv���)|^	��u0����݉yk\���33�{��d~͚'��,����H�d��t2��i��X�S��k�5��`�� �w����O49��+׮�� ��[Y��a9x�Y�u��[n��/آPӪi��Km�D��{]��ﻹ����Dn�����n��o�� ���-�졟su�.�0��=�&���y��R/�7�g�ڒ.�a=�����`�tl(W=1xR����}�V�ܱNK��
���������$1�SOo��v�h������ ��D8y�`�1�R��<>瘆�C����c@�O.�Uf
�7�6�#�e��s����jߗO]% C#�*�U�ۺ��~�ag��ņ�ת�;�WC�m�7�T�
E��|�2F�=��3�c���h�5yp�n��Mg��d�V�����bP���c%���#�����h^�\�,��i��|9�i`�+!���u��*� ���ƯŎ\�_�U�<`ܪ������{O����<�A�?nG{'=wӎR�}�Ną͠�[U����ᛕ�z��=Să��^qq}gI$(��#�zk5dO�l��V�̡βh�	3F��d���"�U�^5Α��V�.)��{�[�k�Pj�'<�>{�30g�"�O��@�p.��/(Y��vl����5�&,xz4�7�}�b�V��B��Ȧ���_��fo:i�ݶ7D�M� O��W0�fͺ�uw֎����;�VޝMΓj�=��dխC�K�s�L�������:X,{��';�mD�҄����Ĕ\�j��u(m�H'�Nӵd$"�ۻ$�B��:,��7
4�ͺ�-����ևMN$��2YsD)���{N���y�Gz�G)$&�q�nF���Fd��v@.�cSɊZ4]��m�Jn�	 &��[�9���%�M������@���D	:V�RO��w���D�]�R�����%�0'����^�����+{��2�w���ď�p��V��=�c�C��J���&�p3>��T�M?�\Ww`�l;a,�,ŷ���/c��Y��bq�D�ƺ�����x�YGn�[���o-B�<�OT���i���G��˸��(nS�|��%��'��G���dW6p���q	�%�����+#��w3-�l4tf���!v*9��<���r��jΞ[BтKY����ɳtԜv!EWU�kO2r�Jb�6�sC��R]>F�����c��\U:౉V�W�s$�A}��ش��7j!-�aȉ�
�J�D��2ӵa�8Xz>��qt��}$*�W[�]���f�5R�Fek��Vd;��S���be.I�i�j�(u7HQm}��΍�64��-�fŐ��X�Yz��8�7�d(if��,��F�y{�����PQ;�u:� �4��4)���H0���Ըz����|3x�Kx9�̬����iWk�1î�hn�e�
�b�z�\3�s����Z��J�%o����4�E��&��mCn�]�9�cY��u%�iݣ��B{��
}�M=�(�<dݖ�������v���2�.�XN�&�G���t�5��nn2V,N7��]�L�
|�:�����Q�����RW�6Bi�[�6��$:0�!��7;&t��cYI���N�V}��t�ƥ�c��Y,�ӣzP�>���s)^�c�+k��1@��[l� ξ�������[�r�l��/Ğ�geɷ�����+f[f��;u��Yڲ:��k{w�� q��K&׫vw��v_6d�W4��*}|1S�˦~�����x��:��ޱz]W�\s:ԑ�s6��RUZ�-���m��1�\��Â�f���I)c*���T:#�ٙR�D%�����{�ZCT����\ ���"��Sl���ύ�˒��nIcS��-J��HS�S� J�R�AFIA\���Q�(��$��PA�"���*.X�����!QTZ�Z&g#��a$��dA�P�)�9^���*��XER�U(�R�#��7+:��faQRM
�I�eiUI	G90���*�e\,�Z\��S� �J�.�YA�U��EW9�RS/8��Q2���N�ET�t��ETjQQIЎ�j��A�2@�9����EQP���E��NI)R
�����EG",P��fA�Rfl�H�����]RH"�$#0���(�(�":��r��(��CX"��eG&sF�����<��2��)�ir˝�u�*���V�D�"�̼[C!#�ʈ�#�Z%EjJ�JL�A �O�� �	(x����mWF*��`�]v��8��=�e��Ĕ�9³�"0��f�����a��MldJ�Mp�w)�8f�%���z6H���~���3����3�#H�H{�c�P���&�|���N��C��	'on������	$=��S��Mޘ90���o_��t� {X;ot{���_�͚�g�b�è	��9�ޛ�UA^}��@
��%��Dh���{��яN�v�~}p~�S�0��~�b��~$��{�Ǌ�̛��9�:�Ճ��������&��{O�=��PW�6��+� �
��ֽ��%��c�C�A�Еm���f�o3�fFa������������{v��S}�?Rw�k���7�N������bw!���oI�����0���v�v��9߁�ܮ�
�D�Tb�𯍚�j�_��K��ɖ䒼��hi��n�/�vmvjv��!��{C���G��Ğ&q�����zM�NG�}���P���n�{o����Oo��>���HN����_��w����?_oNO�߮�v��}N}�Ԙ \��n�L_��/���Bv��߮�p?�q�;��7��~�s�&�y����&|q��������NL/����(��9w���m��eӹ�O�xkvf�`���Y����C�0v�V��t�\
R%\�����ك��?���L5�zL?#���+������?��^w봞���S����r���c�|B]�l�j��`�O�bj��r��gj����!
"����U0U~W���u������ ���魱�]��C��������??RC����zw'�9?����ē
�ۏU���90���Q�e��ݹZ��N�v�ߨz����;���s�M�	?o~y������K�~��~�¦&��\�Q&zrң���Nާ��f=��w�һw�w�߾�\����{~"��C����O�@�>�hi����O���aW~�#�~�&�y{��N}���JĜN`�9j�����6�N:h���������Hw�8�/��~���C�k����Ͽ|߮ޝ�Ǵ�=������8��{~���oN�v�>|��������_�������ɿ�w��㽧����=G�zq����mV����/}nD�͞}�vK���(���~��[.���;�@�v�~�y�;��n@��������i?/��������8?�ݧo[��|OI����{v�OϞ����'*~}���P�uB�����Q���k����R�]Zް3�����+G(�wWw}֛�m0�'�{!�\U��]7�WD�A��}v�Y�d�jn
��.�*��;"�xz���f%�݇ �_(��ONI�ΓS�z�pXd;>Uw; L`�����aԠ-��J��}H���~Fb��?��>�=G�o+i���o�np|d��~px�k��ϞN���<I����x���'���}��O��~w�����ᩗD����.���;;y��e6Hm曬��W�?��_���;�}�cӏ��� ������?�7�睃�o��o��;o�?>y�;��ߘ����o��0����<J������so?i��gO�N:������w���o��ro�Hz�����99���[�i8�4~�ݹ�I�z�x�pN=c��<C�k����~G�~;N���w篝��];��w�r�0v��C���< ȵ���ZNt&��3'oC��;{]��a��y����>�x?�?��������|NM�~�H
({O��u�a�l�I����Iη�x�-�����x����������r�_Lv=�]u��Z0�k�.����7tǱڝ���������������;���܄�'��;����}��-�~���?����V��'�`\�7G��=&7����'?�����`��g��)�&l���h�;�8�������
�~|�ޟn=��߿<���e����������t}�}v��N�O;�#o���<v�F'�����x������۝;����w�>6�1z�Rt�f���C�����>�~��x��שpN���r����O�!���ߛ��\|Np}�{BM�	>}���7�99��k ~��O�|���~�]��_�}x�z|uQ�ߛ�?T)��?gl��X�"�
׻�����w����o����5m�/v߮�z������޷�����7����8����{���S��;�r��8� (���_��zL?��Ҧ��w�ɼ���H~O����vf�������;�nq�{���zM�����7�I�����+��~�,|O������XP>$��x~���aM�	�i3�[��o0[�ހ=�yv�o\�h3��*�	�ܑ��?3k�_� {������ap~��}�?�zL4���~�����;z���S��;�|q�yǴ߉Ʌ=o#�7���9���	2�O���ĝ��>v���w�?~w|N�f�$S���]Ȟo��X+J�m��z����յ�����đ�\��mn������I�+��k�rW��KB��o+�a6��=��0ym�2�`��-R��0^:�I	��j	���^;�U�Y��=����� ��M���1ȝEX8�1����������zI���@~��ޝ����������x�Nһ�{���Ǥ®=}���q��x�������N�=�������]���o�zw���ߘ�nw6;0v�;0쮝0���MyEqn�7�������5��;3`�ki��4���n@�?����_�����>������m�ߎӿ����?S�v�ӿ~���K��]�}��w���c�N��Ll�����őXp����=���_N?�9��;���s�w�r}���vQC�=������۽�o��M�^����w��nO�cx�&��������c�o�$Z���?�]�����Ϊ����@�������:����������������?��p)�;������;�1?�����m���!����ڭ�?|��
�y��|������w���}�zI�N�O�����v.��hv�9�z��r�=uRM��{�?}��4���s����L���/v<@�Iߎ>�;�{v��?��~�y@?���L�<��]���y�kU3�,����2�<UN!���R˫ܰie�Go����Sݍ�*�Q�?8UQQ�>�}�n뱓r�~�x|�f��׻����ސ�81+�=S��<���C��� �z��.b���cU<8�k�	U*���%A7���R�zm�6_k"i���C�zX�q��)@��y������	OCC�P\В6�x�d�B��U���fU4A��د.����"��ۃgKs�|}��ww��ܖvvHy���Qn��M���,�Ccʵ-J�����ȧ�;:"��
�~|���R�*��K�P�{0l������7nX�����Ml�ǵ�-a����8��N�#x�y%_W���P�������qHВ��#B˾����V0�J򫤲w�(�-|�i�ٺ��꯾�o$���M�v��� D���[μ�^g�E��{uV���A8{@'wi� ��k/�te�7�c^֜�z��C��:_#0�~\=���C�?v3����`�~3�f�=;����Xyx}�r��n�MC�E�E��S�9�j],�}o&:w7<�?#;.I���'N ��-�/��	�3ǵK(�c�lPȧQ����8�� �8��t���T�!����͌�oK��Ma;�d�)��lR�*�'�^Y��Nq��P�uz��A�zr�5�s��i�۞@!^l		l��n�V7N!x�S��d�>K1R���o�Bglsa+�Vp����� C����T�a9����K����}��W����#5��|䳹��F���N8$��}LqéL�i_���]%����t�x��ϯ���u�R�f�/����?.�"���$����_R�����{l���C]����� +f�B����$�$�����%8DZ�H1��������v�/�"x�#|YQ�ѯBl���~"E'��=2��T������q��ۃ�B�)F�41׆4{W ��m��;=��V�w����H9\�����6j@��ow9q�dV�0�۸:g!S{u|�}su�O=���w&Ym��Q�ؘx~f�3zVn�8���3�f��c�N�
V���}���X�X��f��OJJM�O�,Z^�w��c�^��!Ӵ�@NH��4Tӓ�a"���F�=���ǂ*L���F�vS�d�K��C��8�k��}�Uu1�SH���ӣjwBd``4��z�)����k���k��H,ˣ���X���5�uOt�N��p������>�A�۪a�r����f�@{��P��|��*>.����`:1V������w.�-��D�gN.�k�Q�Pkd�IE��V�B���{���
��Z�M�{��M,�%^�ʉ�:���t�	Q����=1n��U'"�ǀpk0�K�A/~�f���g�Mzj��w��Ȃ��yU��[5��]�Q��y�=�/@q}b򟷯�5�觵���N�S���ϓW���~��X�|g��&{FV���[<�Mf<�H&qy�U/�'2ֳ���'m4���Z�.��пQ�mFo)\�H�y�kr��s4��vV�[aR����Q]��>�1�޽�ZB�n�)��ӥ�����v�.�X9��:�����Ct�0�(�u-TM%�d�0:� |ԧn����^�;�R��ܣ�����u6PX��-����ν�F-]%!���Ä�)hB"���=����Ǆ���s��S7��̧gV���G�[��*������єv����k���B�p6���չRǯ�h��MՓGs�}�3b\&d�t��v)�G�|U]����D��V��7s���D����ij@OMjp:T
G5�w�;U��N�<�e
fJ�hkճoM�W9!����~�9��=��_�5v<aZ��cl�w�˪�=Xz�tx ~��x���+�Ǚ��$á���܂�W�6�Ѻ����+��'�%᨞����+�ns��.�	=���~^����D�Pq,��~�g
X|���U��B�%M�N/��ϟ���×��_��ͯU�=|���xx�WM)�j����/j{&뢠���J�`��v'|�0��,�7�57S����^~�꩕����e	�q�S��T�;|���K�h�2�����6G�M�	�j��r���,}�y��o�j�1�������@��	�t<��0�=���׮��,��LY��DS^\�}��t_�F;"-FM��2J���M;D���ꘄa�,פk�}��BzV�KVY��i�'g��N ᓽ#ʔ6��X��7^S��n���9oκ�"J��d=s�kU�,�1���ؖ�K&�M귆�޶�.�}� ��]�8�!�޲;WG�!��JP{{qY��2��U���}������[p�3{��1��Z�VR/�����#^o��kǆ$��Ck�@R �/@u�y��y�4^��2�o6�网���@���LmC\�&u��^j#��ihԝ�|z��V����퍋>RR(����z�͆�H��v�b�}��N�Ǐ��+���n�dH߼P�
���,0hbA%^E�0`��,+��}\W�o�=�Qu=�v,��Z����˖�6$�r�\��o6�G��́N�3N��F]���2퍩����,)KX6w]r��&S�;wb����m;���f��|�lVO0+����-���t�ʞ`4��1#�6���b�˼3�[d���3��$
f��)d������!HjS)�qD۫��
7����9#>�<������=�\��CW�t������=֞}�G��)���@�O�*��1���6[S��Ң��l匂��U�7RY���@�|/�x��K��/����
������ļ��Tny��yk[őX��Y:�vۇ*�Q���TT|>�j� +�bB	�M����
�ud �%���	����X�c��1��C�55,�PE�
�Ć{�۞>����N��+/�ʸ.&v�~�o\�N��ӏw��h�Wo��n�����3�w	v����i���]&un�)�٪oE�i�b�b���q��C����7��j2��H����׎f9%��J�- �k��pD� 4#��1�i ����oL����q7�Yp�θG��=u����AG��m�'���.��V�#�h9O��N6�d63/r?f{��/_ޫV�ߴd��]��p�
�� 퉕���eSDgQ�ɰs��sα�7��Tbݑ��2�e��ut����ND�(�T�2h����JU�h����c��6]��QR���C�h���P�x +� DaA��u஁��p|a�uV����4�f&�J5fnȣ�@�'��~�w�?3F��/� m��e��/��A⌤���j�iΑ��#$hBw�r��
��ܭ���4}U��Y�k�8g������ź���ER�S
�}�f�[�N|�'|
؈��`��<j�P&��С�_����n�����ns�3��G�6�B���r��W��)ͻ��#�wK�̾+�hwY��S8�_��Zo�Vy�cۜmz�g��Zl�ny �!<]V�9{M]M�=���7�V�Cc�cW���L*ш@n��JV�r��3BYݡa�eAn6�ݶk��`�Y$8�n�5�eң�Ca��[9Y��9HI��:Q�}6�{8�m2懼����]�ui� =�����a���Jk���h������������do7�����8�V�!�C������~��ul��/��ŀ�������36��n�����d��UP6٦6��/�Ɨ�?���`'��x7i�\|���+砆#�/���}��>'�ceÅ�W�nтx}����/}���5����� �����O.�k-þ.r����&C:��Ԧ]�1��5)6Ц�/��zm�}�Q� uH�EG�D /��.��T��ە��T��/�K�^���Ƹ�Nu8��d]��Nq�^<=^���W-�����>�����[uM!��R<'�F�k*��uL �[>;�H�'�01h ��
�B0�U)��oC�<PL��8w}wi��"a�bP�H�������D�d``79)Ĭ�÷�rL��T��[ix��0
`�:���gu~ι}6>��6��m�6��,i&�~j1z)�j��)h��y��1P�	7��Q�`3h4*fp4+��$ruE6m%k�]y�Olc'Pk��`%�o�y�#�UO*#�o�D#ڐ�t���y����,\��R�O����C�]
��!�Pv\O
��vp�̴2�*��>۰��BX��;jsh�_h�
�׳��k���N���\]J����H�:�ګ�� �4�"�ګ�nh\bRN�u���`oOw��ĢJ��-Q�poq������~K'�@��[���|lW�{^d��	<[��5�Ǌ�N+�fmL5y�����!�ݙ��w����^�w���:�֟iV�/��d9x�n����x��_X��n_Q|��׽��M�ϣ�����¥���{��]�rjX橘Dy ����2���4��bZ���[��s���1��/���҅m�頮g�J�u�y����g����a���(�9̽4`E;�M�\ejU�����=0�¿�XlW*�^��ݎ'e�������4Q��(��U�&[�PqAmQ.�E��ª�^�ڧ`n��t4n��Eus��W����ͬ��ݝ�O����u�.*�7������ηG�V��h�{R=('k�&��/����������l�t.��� $�#~��+�Ǚ�������Y�t�×e>��j��ݎ�(W�qvՓ���OEV��5�s���|Pwy��k�W�Sȣpֵl�M �:���ш��AV��K�߹�z��(Wb�>mzrh���Tj>�y者�i�[�Aʼ�o��FB�Yz�f-�F^���kfJ����X=L!�nCn�|$�ʃ�7��r��[O�F�R7e'�:M]SH�6�����4�i!�)�ܳ	�b>{�U���������=�����"m+��M�#�?<ȚwY5V�6h.Є�A�XF�Ŗ��'x�ƛ�|u�T.=�\F�������C�413fΑ	ݦr=��㮕!�������(5Ųs&�*PڙO�b[>{Vk.t����/��%p��	#C	���tk%<ޘ�+%��y����t��F����ҧ�Ŋ9v�o1(��TC�N�cd�}(��������Sek���4k��P����.Q)�gI��"a�x[�˩��B��u�1��p�0��WzP��"5���:�1��4��e�;��u��{��H�FeD�����c٘���h+<s�T6�Ձ���+������Yd�L�BECM��N<�6�d�؏7D}@b��o l�1<.�����';f�
w��ʚE�Vu�k�� ��툈����b��jf�;�۪�Li��5}a����R緆*�a�G�t�BX%k��
;�*���K⮊F��v]��]��r^�/�{`�>O1�|'9,�/�V[Q��w���>z{Fl��(�S�ԝagSY[��}�)W�s<pM,��y�[�������=yln�f���d�4u����Ʃj�65���7�H�W]<��o��r��__I5s٘�U�r�b��"�U��d��׎�r
�������x7M:�����*�:\�JN#X��T쵦���a�������~��&ըf?�Z0�}E	]˳��������Tk_!b����Jɨ�4�<K�3|Z&CY�΅\�>Ku�j�&�m2��hk��6_V��`���e���q��d�$�2���<|��a3���xp/q��="�� �����p��n�o���{�j伽��Q�)`A�Ϻw�,��3�<Ρ�v����C�נ��n�b�Q9Y�wt�|;)v\z�M@�J^��/�xo
�in-į�<(�%�=�gms���S�Ո:I���#H�'�-v*��
��u���z��[wМ��2��1oz�v�)�(;|��մ������p����>�ӡJ�K��k�N6���n��6O���5����4{ia+o�k��C�s�ifDBK4�5Bb�;
+w�o�)$�tC�Aڀ��a�Ζ.�Lso�4tf��&�;�]nMh��nIp�a�yì̙F���
4!��5]x�uf(G=ojYԥ-�:�O���WTٵ�2���Z�l�=���yH|8������YR�oZ<�f�c�}p��
R�\[h	6*�C%
�/�uZV��g2m�K14d����}��0�׃����RsY�6V��S�����@srU��-�aI�.R4m���%����5i�����n�������QW"8O�B��"�UU�	K�\�����$΅�£P9r�(�
ҺI�)�uH9�\��Q*�3-B�gBJ��v�,Id����E�t#@�������.��D�ZHQr��\��Ң��O2�"edyi&DW*(�E��D�E�9�\ĸDU�*	��bu�Hr�T�D,8J�P�^;�R������œ�*y U��P\�Ҹ�U:{CB��Qh�T��q�s� ����:��䘥r��*�K��$&�:�r�W�fU�""��H�|�8L�5D%�V�EPE�r(�d:��eQPQr=G��*+�z��Ws=Ԯ\��""�XW"���GD8Ns�𪳤h$�%ʮy4T��(R���~#� ��AԲ)*�u#gJgD���`���OV�EK.vD��M4�3��}CaEN����nH$�����}����������Q0��/�)Sn�8C6Pb��A�|TP9��U���LN1>�79��/�Y����.���y'��, �Ԫ����^�5�5��t��P�>]�DjW-��~��v����<,��~�5�]h����wj�̍�~�Dc�c��$��,w/j�v\���}����!$�^b5t�`�Ŀ@��ϲd��;u��u�7�zЗ�v)>T��Y�h�9�؛�+�K�4�Y�>�'�z�Տ0q�bv�̢]��) u	�r��'��6t/�g��G\,z6�U�$������+��V;�f�9���NN�@֬��0pJW��T�4�ͅ!-m5�c{����,)V���k���`���O��5%��׎�嘵HK�n�E�}]����{�F��S�5��_�������kD��p1\X�9﷙��im��Y������v_�C׃�U׼��=X�{�)c��n������zUomeߜ��S{�C�)����&�$�38uc5C�'��-}�o��.�����8k��ҩ
�_��v���W$7���W[Z��\0�@��]{���<�����,%N_5W��w�����\F�^٤;g�	UcE�ӣ��������Ր;}�c�ҹ��Ft���v���N�<�%��=
ճ�q��,¬�P���Gc���}U_W�x��Ԧ��p�9�ž��`�4� `�l��K]u���������b\G�C}��b�|R�LRI�c���A���߆���V�|����n-#�{ƆG�� ���(��?��f�{z}=�
��V`__[��T=������X7N��3���u]ͷ��%��p�b4\�.����E��~��Qb�z.�t�P|����t��+��#���d�{��h�׷+�f�w�O�K��U��s���,�A��z��$i(l�-'_�-��z�]��ޘ�u��Q��|9���Y�ؘ��O�g����3;w&r��T�	�/דY���p|���!,�!���;�$m�&9�l���#��>��'�))��r;%��_�G�zЩt�7���:���T�O�,��D��qyA�ڂ��6���EFI��z�_�w~,D����@WP_�aA��^
��t�pAZ�z�[�R�o/!Fi�8"h��ށ-�W�TR��f3��m�݁�t�^]�������V޼=��T����÷G��Oՠ/-�)}}g]���� �]�3#y/�]ޚ����Ӈ�ؗ��t�x.z�|n:TFww)BiԒ��Z-�մ����qq�b�eA�[x�ӝQ9S;�y��������?^���0��4V��
r�gļ=e�������f�&6�ٹ��������:�!;�c"�]����o��Ti��s���=�$2�^�\�s�uw�qT��GZ)VK~"hϰ��!���i��mVx�,�O�ǂ�^f3y�2�������R՘n��Lx�
"��67609�wtr�ݽ�2�kҖ�.{�_ok�3�ȋ&�j��W�ּmv��������ڛ�{���rש��^"�-ܭ��=��ΰX�٬�X< �1;��}�|XS=vi�*�J���2�b� j*E&vk���/�w�p�=���V�µ�4-�C�W8:�؎0�8��Ϭ|�����b6�H�;e��LЎCVjn���{>�x_�����`<(�||���+����r����Z��g�>	 ��s�*�������~���֭z-��}m��fV�߫
U�� j��7t��烴���3�&��6w�g����)�p��Юu���_5+�C�k��k��F���%�VyW�"
ߑ�8�!���ྞk��`�3�:��(�,�"�ç�=�W��Θ;��ۀ�o�w��&�~�x{���]Yq��ȧ7����{���)��u��l�99����"A��ǆT�9���O�w%��p���y �,�5c0��e���ڃt�'q�:�*�������o[��]��˙���� .vk���{�������q��� @.��w*֕O�~�ˇ���v�����no�>7�z��#ã��~��u�^���{{��(V ��Ɲ_��i��ˮ���w��&��/K{��~*w@���44A�[�pѧ�}x���f*�r�y{p�N<��'�|�J�ym]�ƣ�f�-~~�
V@����Ǖ���AyQ� �/{^��#ǐ�y=�Or蛆�G��q����Iٮ�n� $�:�'�t���kw�*�81�U�J����)��7ۋ���50������t:���/|�f�!Ȼģ|���O��P���Nk��f�V�+E��{���}���7U���WCC	yn�w��&{Fn,�U��$E'��jl#/+W;�͵=�C�}^���<ƐCb�_O[Cҍh�b>Y�W�i�Ǎ����2�fn�ϰ�ݽ�PLEl�$���������f�S�S����F����XlW^a}r̓~�BN�Sy>^b8����5Z�,�>�Y<������u]��c�`I��Ց��� �Μ���[A��EܷKu���^_	1�k�Ʀ m��wL\WU�x�U����|
<L,�S����^�Nh�$������c%	�B�6���t���!%N<�굚��2�:7Ui��y���6℅.Xښ�2�gsҋ3�lѯٗ(����\�vWnT���O��}_U}Sbm=�ϸ�p!�3�ʸ}��)F뀸��x�{��������Et��+A���`�9mfv��A�]�xޛf�к��#< �F��!;'L�B|ĥ��晛�ݔJǽ�����ۆ
C��VL���CJ��`�	�Y΂��;���"��+��<�9��F`O������<;��h��F
��Q����*�y�h������eR~����諾�p"���`gf�_�0��v{�^�puI('��V��O�]��W��{�I���	�F����>Y ��P���J�l6�F��b�)�Ptjkr���ع���&�zYi�'��hZ�0Pi�6��1n�@E���F"]���=YNe]t�Z��2�Y�C%L��G%?L��fg�
4b��m�I�k�t��$i��[ncw���zNpB��š���|��%$���g!{"h �y�*/a��o�x���Z1�f��^��ܿ�4����T�;��T�i�[M�h4��Rۃ�#�q'd�[���gǈ�!����fm!Ԋ�QMb�9-�;Y��{G`Nӵi�>*t&*Yy��s�Hz��>kE�GI���o�&d�mB��C�%���%�3�KT�m7���y��3��Y�Y�fEK��kb�mb�Q���	�Λ�m|{��>p�)���zus�/Ƭ�P)y"Z�d%$ب���bkhmT�T��ϒ��2��)��;	�~R_z9��wQ�|sf������]�����]OV7��c�5��f��"�����xש�섏�G�ώ)�Ǯ[56*�e}Ջ�D��z3!�m{%n��~��7�2��z�S�����Ϩ�[��>^޸7�j?*�����ťfb��M�
My;��F*�ޫ�M�ej��R�QbW�Ju�^�(]���TMz�f2ywOEY�x{ZF������#�'l?meF�Ac�p�����)�W+��R��/L��� ���-s[�Q��i$9�Pוaͬu��T�^�O�H�e8ǻ^��� ��,+B+�i��,Qt:k�̐��60[�3�K:����jF��q� �[-u��V:��� E��b�����a@ �<4��D��el��Wa��m��L��\�q��iu�Ӆuy��ѯ���{�L�i؅Lv@��\Fv#Մ�����C$P�X}�u�mJ�F��sH�]%ɞ�Ȳ3)Y(����8���M҇ʼ������}_UW�%`珚����кOΒ�dΙ�;d�8Yk��+B��7���뜭=ΚU��$�0��=L�O]E|��{<2�j�{~��u���E+@��!Oå8����=y��S0M~���ð�;��������F���p��*%[�"+u2��-<�KTR�c�`�*��A6��#��~�rg��ʉ�e�i�	Z�	�W��*S���H�X[�c�������l�;^�;v�i5�S�ݑ-ZS��Z�"�5�j�����sbY���W^����N����|�<��W�uxb���+�-Lci�-R�j��D��[�N-3�E��]Ϡ�%��D��>�8�g>�S̮垑(?w��bǾ������
��;o��ajz�S�m%8J�9zf(˦Kp׳���L��2�{F��z��s���z��.��8.��z��8�"�V@�о���a�E�"Z��g>$<�3n�݀V���%����:���O�����cST���Yl|�r���Y���>�_��+� �Y7C"��g1�+�[-�{W$.ƞf��gi�''Iv��:�ūK��fo7��Gm0���r�|g]��*��>�{�٧�t�,y8B��ګ|o|vz�|�Z��=%NM��?b�7�)��êo���=�w�覟E����6}~ȅ֬ZV��+)>E+�ө�+��rZj�X[-e��N�V�V
�軼K�Uul)�6�#�ć�wqa���A��݁���9�hsZʩ8�1K���VN��1F��^��Y����DM���AЫ�y~�p7��&Os9{�Y����򒧢f���=��ދ�b�*g�
M�i��<��5�+��=��A��Y���Kp�����m�%�����bʀ�۲>��kU�P]e[������p�����~�k�ǬH�o,�ƕ�L@3�B,����V=<��zRO�u����zʫ�����q	o��3!i�zkf*��-8�#)ó��W�x9� #�T�����8}q5��=cj{Խva7�޳X7ԫu���d�����?�e_�N+�u#<�/�#=�[Z�Z�`���{�ȳ���N�u}�ɢ�2��Ff<TeIw_""�cb�j*�kx�Ov�]�.�s�SI�P���һې��ɽ���fA��jda�]d���o3{�g��9�ss�_�K��^�/4y�Z�'��2u���#))�n�mΖ�~3W�g�"��[Cb��T��)�m����د
�iy}����*����Y-#*�d&�����WU�\��}��3襦}�y%ҏ�11�y�y�Oh<��5b��ez�d�WZ�fSը���K��p]ګ*wi��b�}��楊D;ԡ���/H��~L�y���6�}�?ywH�����^|}^�����+ujjc�
Veӕ��,1*�֥�����(�>�D�!;V�=�%G�<�����ŕ�ЊW���}#�ƭznׂ���B�C�f��e�n����ތ��j��ԚT��D���{�9�q�JEex�Lϖ��!��k�!��o�B��a]����艝��5�{���r|�E�1R�3�&ݴϘkd���WlmJ���SԟP�*Y�v��2��uoe-�|�G!ɇ�d5;�� �w�p�����F#�-�f9ڴr7Y�u����
S:�ٕ6��I�k�N�^�͈�tޥ�m4:8y���.ٗv/S`9�����O�}���^�������$�R�nL�}�|ܟ@+"	�'v��[�=f����>���8��|�^7�����j����!/�&�����z�S�:I�Y2��&�m׺ۋ�O4�$?< ��uӨ�������my����ܱ	wB�Z���N��jʹ��tj���q>0�l����ќ���۔	61�����n6J;�H0��zKT�lT�[AMM�J'���C��TRL�K�OpVK6Q����^��թ���b�".q5�3j����f|�Y�Ak�Ⱥ@�O|RA"J�U�o��W|u2JPą�jk��n6hO�����e[F�×��uK4R�hV�-z�a�
�٩�U�C>�k^�˛����mAꞜ,7���T5m�QE��o�����x�u<��ڷ|�h��/.��owO���SQ��V�`�����Z*,[��X.����3o��IB`F��Ď|���n *;�,�㇍5�����G�"��GT��p���L�^◔zo+�"�w��Q�8d6�_ܪ�8I��v-�uvL1�7�	WmY4px=�'���E�eV�)�Z�
#��B��Cx��$)ɢjF<�٪`��h�f�Fƺ+ ���Ⱦ\˓��+�+ڏ���&��o���(�}.���FVTa{B��{��U��yV����](	��>�"�`M��kЍ7��t۷1�
�*�Lwl�t{��?y��n\oe�U�$�ee����\움 �Go��n�(S]u�e��ұ�f�50��h�θ&wd�홠K�W��t(���|�sF�R3Yx�pX�*�X���CcK6�l7�뱖��ɮ�ٱQ.��|�p�l����:7��n�����e�k\�ə��J��8MK��8q��z����9��%'����!V{��jm����]��ўм:�'傃^�P�K4��Tv$<Z;���;��k�QHS�I�
t��hKr�`�gjg-��h��r�4MS��sB���*ХP�3���ce�$��(��:����Tʭ���ww���n�"�ss��ږ1ez�D��}	��ou0�>����%6.nt^�T4�vA��F]�-=GF%=��w^��Ym#�X���F
���)�f	����Gc{ǹ�Z�O��ǫM7�xl���}yf<k��n�w��gb����.O�i�a�BzqP�%�#�h�6�d���.gnJЮ8}���It��Eʦ�ɍ��L۹Qq�w�.j��PwC)c�����;� ȷ�t�I�I�3V�LEc��q�q�w�ѽ!�!�B|�DR�z���Q�\��W�Ow�*^��9�3.�l��N�ʲ��7�1����mn\�{����e1Ϻ��CzlL�h_Xx�S��0�<lVZ���L+)�B�7Z�֌�� �GQ<q9�B�W�oS�7�_BB�w��:��t�q�t�C�+%i2�m��|�G��F[t(�%�`gI�����j�LY1���7���4ϦamUEd�}�*]<��I��c5( {7q�wb���5s�Zaj�ZR�sj�+j,�[Q2H��:<�lv.c̍�jy�n��ا�{�����-��}�4��,�&�M���c[�W!3�]LlN�| N�]2�8(IL��wxS���7�Zb�^^°�gm�շ��6=�dE����<u�[B�+�^t4����G4���j��v�V��f�.�s7��Hk#�պ}��]���V(u,�sXS��ye�A�8oܦi�1�2�2�{��VPڕyOY�ؐj>��(�Xn͖e�8"I�0�w*֋�cZf���fۜ�[�16��d��!����{ү�\��d���W[�X���/{ze�G>n��6�¦Z
;������)�Foe��yN�^v��zk�:�i-���r�p���F�zB�'ĺy�!�e��@�k0�� �F A*s�d!C��aEF�T9#�Qr��l�q��Q�gT���~�"">R�[J���e�D:hQM6�6���]�.�9�<�d���s�ܹ97®PE�1
H�ܽ3�|^��R�᥵(ԎBIf���H���C1L:����\��EDh����7Z�j�Tr��!(��C�:�J�V9�9�-���Ie�"9Q\�����(��^<���.W�<�ò�yҪ-h�^o:�Aș+^u�r����Ñ�膤ED䜽�9�t)��d�y�E5i�*�RtB���*�3aGudOQ�T�Gq9ʣ�̖��Թ%�O*�EDU�TD�������K�ݧv�!�"<2�뫧��Yޛf�jN$A;~�☹@�w����A�j��Z��8�X���=�[:�\ҋel����q���oy�\xR���qz[�Q�k�J�K+|֎F��N�Wr�T�*6}�[��%�����BO�dG����VOOCY����B���d/Xq��AS��F�F�b%�zm�}��=�
��"���|�d��K>�j"=�VdĬ��ɟ.���cH�,�KAZ��a��"���e�2��N����<�I;f�`�Z��D�4*�gL����bq�-{�P(����B���� �W�b��{~��͡N����6�Ž��������{ݎ4�ɯ>�Q���ڷ��S*'� �쏵��Þʌ�6F�{[��l�����z7���Z�='I[&QJ
4 sY��Uc=S���^�$��W7�U�)5�{]'MkH���<���h�O�b:�^�^㋥o?+��L��d�4��l4�dO�Jp�kE�Zjgb��Zf��\�\o)<=p�Խ��̋��ոt\�0iUksv��m��4��$���T�\x��9SlC҄;t)��Mm_S���R����.��#ocĆ6F�ӌn+�%�{��*�[�V��E�¥v`���Hd��*h�a�.��������)�O)��~y�*Yb's��gp���Yr�6�ޫM8f��4����9��Q�L�{s�)/:�;���/Ŝ���>��tVpj��N��}��&��o����iV�l6��m��+۟;ze�}}x��kĨ|_��Ӽ=��b8�yjpګ��+e�פH�|v�]�n�-��v�V��8���]�w�/���X�a_�����������i���u�}G������}Q�*����EhU�L��Z9a���N]e;D2˒_䚽��i�m`�~�Ni{FPm�%��t�g.�K�%�F7Q!�,�U�D9}jfz�v��ie�ʷ]�>�$Ή�����ݲ��܀�LRܦ
�l�q�އ2�}Z�虁��6vܾub��P�EU��3#��Ԇ8���R*R��
|m�L����5�U˛����K����"[�R����
���ހ��_&z�r��E.w�%n���u�#d���\�8$F�.N�9�=Kx��ԝ��X���fWU���xIhx}������^���.�m#$��Q5l2K�Hu0��wR�@$�ﾪ�����hƜ���潥-�wh�[�e���1D3�=ף���k�_�ݞ+���l��O���fy���-�"�$�O���BT[1�.-M"�5��S�p�Ne�7�v$m�v-�%�YqL�U�ݴ	+]R�SiJ�:{ч��)�ސ^�Cf{��}~^��3�a>�i5�i���e��V����s)f�4��S!m��5W�������˥���}��c�k���m^��@�E�L���>N��lMm�ls�>�K��?VC�g��W���=}��Ʌ�!+���I�W����g����?&�����m�gF�n����!��ު*[ǰ�;�;U���[�᪟�����U=�v\,����/+�E���qJ�^�^�ga߱�zew��x�u<��^T�ueX'b);��ك�'V��")4�	uN�s~�õ�����ew����鞞UW�w�W�t+��DM������u,o�M��;qK��y�Gۃ@��]�b �G!�[F�Q\z�[�_gB5�76�+�]�ժ�9O��Q��OF��R��ԍZ�/Q����r�]�G��Zwv�R;�C$�Ā��f�i�GifJ��ޭ�d3����"5�\�o3y�1*������=�m,��@�`n���u��͸[>�䵮��PЦU���e�s�=U�7��1��<��|'aƙh��L�rR[�)S�/K$�'w
����
�e��R+)��4�D��/�A��
��e�pWk�i��c�Ji]�>�b�����eGg'!��'Z"Ct�GL��;�\4{��Z#����4=%>��W�Q�;��m�O{,��ݙ#5o��No.�'ڒB3ނ��^�S�Yjxm���ǞK�`�C���s�9�L�>�zeoJYFAͳ*0��=>޾�s��j�
w��7ТJI�O'0ݞ�6��7nz�����@j{}��K��H��P��k�'Y��Z/g�2M����Y�yL��8�uL�&�LE�z�Ԩ�/��EgM��^�����w{B�\���m˽���5�S!,�lTD\�=N�O+���'�q\�ϯ+b�^<֘��H2��,�q(�a���t��2ƝSf)�B2e���U��Yod<2Y�`j ����;�B,(�܂���0�q�tȨ��V�q9Ě�2����(z?\+S\�p�L���.�}7Eiw�;��k}((�&rA��5j�ZS������|���g������2�V��T�y�S!4��J2u5�9zŮ9)`�<م�d����[��-�\�;nyף˫g�|����0����P/ޱ�D�o�g���Sjg��ͱ�&��gL��SC�+ެe�>��]u�s�b3�Vfw����i{���%<���MQ�S訹�[>�ٚ�	��8P��,�ʺ�P����]l����Ko�L<�t����������{j�S�M40+�3&��Ρ�QF�R�`m�OE�$/ژ��=^Z��P�������be�nͩ��
�e�m4"��үX��c�N��"�X|�m�yI���K4��F�8jX��u����Wg�s�k�ܐY��sC��_;ʫ���c��lg�^�%��7�o�D�P^~On�q�Y����y�`��Ԯ�t6x�;o��m�dՏ+��L5>Q�#w�L3�{Z��&�$Uho�#BU��ܘo�Z����'T�2hƶ��!'�FNq�6;��XYF&'���]%͙E$����S'r�Z�c�x�V@���ūa$���z�����9{^Y����蝦�h\��� 9&}�}�}���Ԍ��E��{̅��e���1D(��gS�2�؁��5U��b�I��I�\ǰ��b��-:J�	PLB�m��].��(�}�û�;�z�FI��U�s����A6*"����b�y�䦚����^>K���Mނh/ZW��q,�n=j��7dMiNMh���4���k����Z=$��ԟ{5f��dX���}�aÛ6�����xh��x����$��ϋ�J.}��gح��:�i�=����/��͊+d���Y���a��s�O:P�x}�{{W���C��3�yZ�1�e��{�}�м��P�7��8��BͶ�[jj$�z�55酐x-A$��.�<�������p��nό�>�{�����>�l"-0�����Nv���^�UX��=^{G��ۧP�(���8Xm���(�@Z����G+H�gM���f�잖��V�D���aB����ROt�}��k�Y��}��+�}w;eo�S�sws����DB��<�#ǒ�.�5ؕ k��z>�.���Cz�0r�r��éV �rn�=z����?}_U|�c/5YkŨ��EsJ��>���[,�)�~j���I��S�+�G�Ê�x_�3Ag�<f�Md��-�U_9��/�8g�t��U�嘚�zSr'���P�S��(��m*|�e��s,5������WFe$��=�g{q�\�N%'n�b;~Z���z.X�J��6�F�slp�LT
qp��R���4]H^|;>j4e��b-nZ[�*��`�f������χ���wN��y�UȦ��6�ݦ"�+C-��,d%F�Ƹ�5?B�Q��	<z����[���\�3U���0����uz
��7C4Ŕ�GC+����i���e\^��3�q���kBF��t�y�8�yz�7f?>��Ǫt������^9P��U{��=��4F�7��[��b����fY��"Z�dL����[F*q�C�^���c�0����f�'w���Y6iG.a�V��j��Zl*
��4����t��"Cur5����B���FϩF��x(�{C�*B����nu߽�S�t������7dP������7�Q�����y!�w�X�!��6�&�X 5�hH��\yO�UU_Q�7'����[o��U��R.۬��W�����_��R�k�o��lB�Yä`|{��jS��
���Êo��6���/g�o��s�R�@w����ڗ�si�����BE\�6X5,R60��KR��C�"d��E���j�AX��i����v�9���k%y��Sό�ߟ���4��M`�q9�=%�s&�h���LI�H}叫|D�;����=�Q��&%j,�}ƣ�nl�L�'F�$���^}T!{S�g���\Ѯ�����P���Ÿ2�N�6֓��L��HΟY�����:Ċ�5�Y����u#[i�U�o#j�UM��8)@$�Ιh%Z.��,s���\�)S僊�S�������d�]����Ud�\�p8�w�f���$��̭�O0�(El�<V"L=X�{j��~߅1������by�������෬���Ϯ��4�`cK ���j�ܹ���K��e����I"%��4h�-5�� ���k�N�r�::�JiԃS�J1�+�������0�~3�2��U�����k���Dd���fJ(\,��M����e�%l����g��UUU��>�~MZV��=�f��s����J�"v�A��u^І����wq;n������R����U$��u=.��T;|�鉺'w�bP)U�7�r�iY{����:,�&�^b-��jhmT�@q�1hec�P�	�����~��ެh�h����ѵ\�xJI�W���Mm�ƛ��M�C���{�����W���q�Jr�����j�/Ԅ�R�2��:�A��<�qH��R9El\�᰷��[ڲ`�q���~UG��]f��Zv��\խ���D�<P��udꮊ�c��oͷ�3訹�繲�x[m����UBJr�)ͽ7��(�4�G�{�2��:��7P�*s�uG���b�lڹ��Ja{�d9^�μ��i�z0R�--��r6�M�h+�g�=�D��|��'μZk�r�ר����==�Ɉ^�=>��Ord��dA����!Z��y�m�z�� �ł��Rf.U�)ˏ�m�AB�>�Z��k%����+MxbEgnǢ�ALAZ�W���3x�P�����Iׄ1��^e�u���6u<�E�I�qh�g��V�s�7h�������x����.���i��Lm�TU��)��.t�|���ٖ���K�#���/�OZ�2���'�A�L�3�1�;��"
��Ag�P���DM�n��������6��}脰�=+
��*s�3e�������d���z��P��Z~���g��+�7�<U�>�̤�u�W�Kq�Z*eD��~~��ۧP�|����9��Kp%�)�ӕ��K�t����4���!D�bܸ���H���1�t�eQ������@��� �1��R{�K(���Ea�S�V�|B�Бڬ�Me�y���4��d#j��X��O�3k��B^�L�瘍�hn�]^O�mL���k}��"v�?�̳���ٵ��w�`[P�������2ʳ�l:ϓ�Qx��ٱ[��T�%爝�!�����Bϥ��/��b��޵V��a�!ua�;�n�m�4��V�h��c��+Y+-()jZy'�}�]��G3�3x�O�0k���w�<;L��z�qU`D�
��4����r+;��*��ν��Ј�M��_%6��U���8�u�B�ځnf��;�R�;����CwF�Жΰ�ÉWjT���C�4'V�Ĵ�b6�'P_��"^�hJ�v�s��a�j-���l^�����.6��3�&�v��kD�G9>Pm,RXwb�vK�,m
T��*��@�!n���^V�#-u\�.�r����x�{m�=\YCp��-g`�����Ib[9������,�l������e>�cC���"l��Kt��&B�NB ++{� ��b�\n[����̑�R~k_�ڂ�Yc5��Q5�<��e�&��˼zd�G!�wo���g�'S�Uj}nIs$�wC��Nw{W-���LalNx�5��\�|t�|}���8����E�
�b��i�P�'��4^Wac}
���O=��A����oD<��z�k��5_Ǣ��A�L��=�5���p��5B�-1�<rsar[f�l �=�Æ�(y�̿p�[��N W����q���Ͱn�ӔhB���������1� �'iW+�b���o���[��?+�S�#�N���`���E7����:�l>�)��L�~�s��S�j�g�1���B��z C;Wv�B�gZ��ɝT�qc�� &>���n�(S�6U��$�m�O�Pm>���H�Q	�$���j�;ݡF�E�7^�$P�������V��P���Gg8&>3��V)n����������������b�1ܭ=��J�3�a�E���hj��Ǣ8��+�չQ�,�[���5�ޚ���r8���o��*���B�"�R6ì�Ӯ��aAt}��wX�3$�U�*|��i���r��tbV�|�� L?v�
n��7f�x����=��m���r1��޵�k����`_F�T��J���'�r�7�V9���c�[8�ҋB���a<!_f$��8�T��d��0z]��Aw\)�wF%�GD��F̜��t�Ԅ�/��Fd��u��
'SZ�7Wp��ի嗃��q7���*�^���0]jc� �*�e��%��>n`�'�C�'��c�zk�Ut؏M0�Y�(���ŧ_�V+}v0_�!6
�]1�NS��k
Uq��n��ϛo������a�'��Sx��5�<{r���������J2l:�K�@�]���׽��2V�I��ħ:8�5ŕ1���;���2d��-|��G�����Z+:�fr3��G0��t%�+��3�;��{��Q�;��nt����X:1�xW'5n�z;��,VK���׋B(�K�X�:t�,�y�'FH_P���O���h�Ԝ�mYS/}VY�Jr�.��w��?�����D�zaD��<y�s̍J�S!*�AWp�\��oku�˞�n<;�r.�<yr(�<t���!^u+���U2"��D�.|��Z���J��<K
:t��*�P��r]S.'�2L���>B8���g�xm#i�p��.z$�5J�Y�U�蹐�ҸZ��	�G5(��w
�:�鮥��G��gJS'q�u�/B�w8UFrۻ��L��r�T$�Ӯ��� �tйf�(�Hg��z�Q��hhD��0��S��EU-QP�,4�\pBL����#V�daNyy�z��ˢ�\
v���r�E��V����\C���L,�Ң��&��ʨnB�:.�¡�ܳCJ�%u�+��]Aɧ"r(.L�pfXW�	�"J�$�s�U��t��o�j�p���X��,�Ӄ���$A݊Zfk�xQ��}zb���Jfb����1�wf�_���W��I��y,�$W����,-���!�j2J��Ŏ.�P�Cm�^����s�T��}�u7:�:l����.W>���>���?b8��3)�j����EL5����}Kv�)ӯ�&�_g�Xy���XY��ԩf��ߨ�,|gGj�ٍb�����7��P7r���2ʹ�e�ۧP�(�p�1�%7b�;3[�.������ղ����hfi�e����Qpn]��s�7�U�����hH�`�ef�iDfQ9�#Kӯ�g�����;Zz۫Qs�{�2b&H�Uy\[^���Ҧ|�e��s#X=kǙ�+5�1"1#�����/��=�}��z/F|�9Oo�ֈ��t��u��ݻĄ�&������C�s�ztڙ����5{U���dĕ\�66R��V�5�m�7xt;m��ݴ3��.NM[��[�E�I�%mY{ݭ�׺��פ��sR��=ҁ�t>��מ��']�ʱ�l��#n��[0���|�n8�tb���x��D��̸�J�wl:(X�*n9�"�ȭC��h�HwI�6��n� ��Q�bԏ������Q�x�A�]'AS9٫8���ꪮQn�I"C��6D8�L�Hӗ�TW�M��O;�����h��y�'�f��Ǽr�h�I�R�m�Xe��(�L�ф��1_!zn���o����H2�$�pRk[�-�4��Q����9v;��ـ)Ǐ���'ܝ�5��Ŕ��5����>O�E�jk�*q�-l�6�x_C�{
+�bi'���Ǌ/̅(B�}���[� +ժ\@on�(����s�Z)l���YV0��6��Լ�<���'X�'k�zs�����c1���K����4q�~��P�/o�������-#jsR����3i���[ؕT�%�<N�s~�õ����)�I;�����S'�h��I��p�r�I����l����6��X&�ܸٖ��`��l���+6̵��~*y͍t��Хf�{>(�*�C���4��vK�}wC�����.��넵��
>�{6��d����L���<�p�D����L�w��/�
�|s��~x���iPd^}z�ݕ��dV�x�Bjg�57yZ
����l䂊"�P�W�Z�����z&��;��h=\_����eB��7�/�Vc��s�Sd��O�+(�L�`�D:ی���ܜ�W��c/>]L��-U�3��E�ŎoY^�*�Y�׸�xƑ��+2�*["�$�,5��h�v�8�w�~��>h�{�[e�����2tk��7��x��])t�\5�υӘ�te�,�e5*u��Ӗin�Sh�}H^)�b�f�C(8��~x#����Q��#�^�s�6��U��OIη����D��B������d�H�wV�b���h*.nm��nH�)�r�S1��54j� ���1��`[=[������2z�C�U��Rٻ"��̒lT�E�bkkk�ğ�Ns�"_���=Jp���ͬD�+Y^l7q&[uNS^�B�!g	�f�!��0߽ޓY���;�����u����+�s���gz��0a���~���);}=��
��S���n��42�i���em&����2����z.Ў�Ѣ��Rv��m��7����=}F�c���o�E@=��p�죓R��G�_v1wԦ�[�3S6M�Vнچ>p�;�j����]N65�sy��(ɽu;�T��h��2�d�{��K�U��;o��/�o>}S��͔����j�b�G,��AE�S6�([�|�S�gUw�n���G�s�Q~�����'�6�ww��-�1A�'��\��Qz��	T�J̶KnѸݓ`��Wto\�g[�:���}��u�}G����������d��5��;���s<�r���4��p��gJ�-�Bm6��jcͶAQh�-��U3��xҡ��-����{��~"m?Ash:_8.CX<�[��4qn5k��4�[:�V�8'4���u��r#s���&�ӛ�t>�w�~�p9��u�¬�V��_��$s4������2׽V�b�&�Յ>6�|C9��t�)f��E���<q���G3��-~y7h�Ŗ��B�L��1 �vG]�"2+_.�H��{��$�7xx2�W���q�=���B��$���E(�1
+��Z�)E�֖�)��2��[�N����������wa,E���\R�����t�]��<�+Ƀ�+��Q��ݲR�e�������u��`�<���'܆Ia*��f��̈ㄨ����T��:%�.�d���M�5Q��^FFLr�1��}UUI$�:�W������'�ޯQP׎sq%k���
�dDl:���;3c���Ow�z�+�z��t��Mw�<�Y���l���8�

����X��P+L=�iqVZ�2���H[L�*a��L$d��������~�;�8��'B�$ϓ��5E���uH�>b�D�Cf}U�ٺ�k�y�|t���XQu��f@��[7�h�`�����w2:�����,h����˧�9���s^�'Yo����:^�}��g�K)Q.��b�z��g�t}s�p''���P���/oR��W�����~��|���S{�H�$�;վ!.���۝�rW��M��2t�����AF� ��{���F`8}<��}>�����V�{�Js~�<��m�u�S�F���5R/��2����y��Vzz_�����վ�s�(����zt��h5�yۻ�u�;̊@�7�!��l���:��K4�Ed��1������*��]��
��T�0�
p����r��������2�BLK�r������\��-^�.Ūۗ�A��]���ف�L�4������X��	ܫ�O9&������y��oy�Y���)9��ڕO�F9�H��Ҧg�އ:5���(�< �[������>���cdaȍ�d��G�e�{,�E�R�>XFݜ�{^
���|��1�^�j����,��)8`����B�A���	��Z��,my��>r�O�U����]q�כ��������O4k���u�����{@�slQ�Ȁ�T�}�ΰC9p�cU�ϛ^�'�0>D��F�7nz��D[AT�ʍ a{�8�d��@XʇR����}G,�<��	�$�&��"����}���kr�BM�\�W�p|Vl�N%�"Ay���A�eM�>�L���r��Ϸ����j���֯����F6���9�Z�3������G7��Q~������_O<{��Ή�F,��;����r�%����^*�<Yق=�~��᨟O@�mYBғ���c�v�J�;s�T�$�e5z)j���t�v^[������|�Qx�]G0�ҦC@�c�'�gvSJ��}�}���w�A�����;�)Y3�۽��Z��]��f˜���r4L�s���Ii��7��"�1.�ml��*��/T鱪��^�4��y�PӲ��@*���;��c;�EY�|����O��'��ms�Gk4[>���T�v��IJӰ^���d�0J��f_�-�5#q�&��0Wr�5�>��ܸfys��$�YBz�%��fz�OOC��>��qdb��դ�v���^oOz&ϡ=�o��w��TCg�i�'�����Ͼ�ֈ�a�0楣�� ��50mn<�^z`�r��S��U�����_���f�;�ź���b��.�N�z����i�V�͎N�#��˺>�M��{vW�����g���Ӻ�7� g�'���M|b��7�p�мE��S!zh�����e2�X�;��ںb��E졦���]�.~[�j��^��,���-uL��J�تQ&!F�#V�������yU�
�:���(UOy3Y���sm��^C�>L&&�? �A��y�jP�����ڑ��̬^#�Cb��"��u�Z�� ��-���U꒻l� ���S�k�:Rզsi�j���]A78-����Sk"�S:K���#�Gc��U��~�V,ԧ��9�ߏ�(�,�U��2/��U�;�:�db�m*�T�� �{S9K���^>Mނ}x��:���p��{�!)&�DE� Ƃ��J/\,����� ���|�F��l��H���ϻ6j^����mU����~q��9�t=�$��5���[��U��"�[A���Qpm2*��æ��*Q;Qjt�Q��ka�P�Wݐ˥EV�=܎m����1��-���>���~����V�x�i8}�$׹�����G��ʑ��W�'[͟)�5�L�[��(tWk�R�����%{̟C���$[4
|���P��6�/s<�g�p�l��k,7N�PQ�9�[��~�����dd�Iy�v�vB��y`���km[m�TSV�}��_f�ރ�Ю�>����h��S�G:2����`ٟ3��������	߷mΣ�o�r���nNNgw��FpOF@�*)xnޛ,�z}�ܿ`雁f�[b`ݣ��
:Z�eO�^�b����f]/u��g�Nhj+�[����ʲ�	u�f�Vs����]�1}K}2����m'���\��Գ�s���W�_�
���58 k�&6V�uH�3�>6�_Z��^<������F[��t�RS�J��3���v�k�ʷ�*IeAa�m2�C�g�(�ov�<'��O��{�<=��j>�~a�S{E���U���dF�S�-�VM�[�r�����6�¾��Iُn����B��K	P�U�:���3⸿5����]!V��"=����[����� �L)�MUri�f���t�Uz���U�q#�Bg�]�Fq��e&�c�Г��_rV��;l&����?o�Q���EW�CK>3�8��«�j���׸Ea��VjE&D��,��I�%���Mx��۪Zًc.�5�4��Z�R\����Kklx���{{І$/=��c�dک3�����T}�P5)���`�)��7��{�{<ϰ����b�FS򧹲�"vAt 	��5�����^�������x���q��p����s�H)�.YN))���0z��B���O��!u�U�-�t���W.^va3<!��+�͋v����x���� B�6t���U�ۏJr�T��}�}��m����"v��`Z��C	����%�Z�+�oR�9���=s��v�.��L��i<�Cڧ��x������,.�7��!�ûy�q��	F��OkK{�*�KB��ՆZ���.K�k�3l�0�]0�6��F���$�zdQ'�I[m	Fz������#����"K�����˨�vp�w[U��m���{(�Pq��E.ͳ���4:ے_��oW��v�"�ۘ�i�2�J�Q��֫�X�JM�.A�y�N�5���%Z8��I��g�hrHӘԨ�wt�[���CIǢ�M�^EBJs_��ICюlP۶��ϴ��\W�-�1�7��0Lj�^�{��}��Օ~��i�{6f����1f�3�7=�ny�"��=>)�5��;I�r�Nih*���Q;�<dy�$u�����^C���S��i�{H,ԓ\���ox)�W���L�j�v���CK�g*b�o :�}�S�S�kU�Oq6?d�����wAE�{�i�5̭��)p" �0�+�\IxvKِC���n*:�-��"m�.m�jv6�1���N�����
�1����Y/p���!R�Ly��u-�%���D�hu�_g�?C�
xe"D�d	2�w��L�`�Hq]�.�n:Z�0��vq�	��
�>ɠ��V��8��i���4g>����(�xsta+K���A��2.���j�Š=��EJ̀�͗�E�F�C	܈z��̚L�^^�)7<4s��oU�H�ڥ[0��T(d7�t���sǧW�ﮰ�!_&�)M�2�o�h��*������]���]�p��ß@���H���r���s�c�(����oM��z���ܺ�e�ƀF�Y6�{S-KX읡�)og��'gc�n
��8�dAV�Y�y�+2ݷ�OB�!��Or�����P�X*�� 2 �]�qQ�[�ݖ�M_q�g\'{oI��6��j�A@:&14��*-]�<�sX�/�wp-W��%9�z�/���(Y�׻$l�@&U�-��2[� �Ł�SX���Y٤��f"��S�|E:gg�Os�2�I3fA���)�Q��i�`H�l?=���>�F�^�i�wB�$�>�n�3��	F�Ub9wԶ�:�&�E*OS��Nٜ��#>����3�#�]3�](<❌�� t鱁i�\+](%]�fG�5�-������uq�1��cKv�sl�����I��i��tgb�'Z�0g��.n��V�tAF��t�g�j	�vY��i�\Er�/��IR���gd�
9�1���p.<w!4�]�wk!K:Ƨ g!�&���S�x]w@���ܖ���Fo�r{�7zӇ��)נ�j։�6�j���Y���8e��V�ZkLW0u���*�H�ܢ���n�� �l#�lc���w�H�=�,�~��P�Sv�-��bܪ-53J�/l�R�l�5n�w5
5�	�(D0L���zp�Y.�*�����%����r|��b�����Hg�-�9������|�a'nfNkE��tF�I��@���*�`;Ǟ����ަwM�Yy�Q�uK��ּ�˶���i��Д2����ە�I�i�����Lt��b�`�c�Ι�{)m�',���v_n4s��ƧGs�N-6�\�.��R].`N��{C��,R�)LAG{�f^.�������6��,{0��ޝ���HґE�'��v�E.E� 6��;86y��U�>�:���v���8n95
�0ud�ig'��U�1<�jC@��e*1э�a�X���ZMੴ��zc�ޫ��F�.�Ą)���˜��E��m��3�S#P�2�,�c%fl-k1���,� �7�J�ʅ�pq{V�	�9���]��F�|u.Ws��`S�VBD��-���8.�bE�.��=k������G9H��NG�x:XQTk.Ӧq�8W/%N�rr�CU����G�H�4�2pH��"3(����UP�br�����=-77u�p��<��M"*��u�2������/$�Ӹ�Zȣ0�Rs�NW��!K�S��7y���&AK�W8x��*jY��u�'.����
�;���9�;�R;��$�/=���))�*F)Z�!�f����-Rѹ����f��Q'wr�SD�A�����s��Y;���q\r�i�N��G)\��	R����j[��{�IzQT����:rY���xD')p�	j��.�U$�N�Dz!���n��I�R�L9�%���=wC�$/�)Jw�L�'�.�o.y�&sX��:��U0�N�g�45u��l�RȤ�^x�t�4�:r̍�H�Y�Ҋ4S�~$ RA Vs����S��F����y��8���ot��n䣪���j���VS�9:�ٮdd�-�����4�6����U���UW�^��[+*&���ǳrD��O,�&�D[C��U=~N����C�����}�]���+܍X��2�5Э�7�D֖BY$ٕ<^o�Ѫ�V=f���޽v�E�?nӑx��G�UKA����FbW�k��KR�_{�zc��4(�/˥f����jzs��W�s-��+�r��x��̡�رY:vUQ�h�$�<H��d�T���=P�[}��g��������;z�թ]h���&\8\�W��=����Gg�n�UZٟ����X������N^�aD��d�Xz�sZ��J��f_��ӱ*�Cw��V�Z��/'\�~h���I�Jt����zz�y���ݩ��D����^���s���`��oU�qw,�7'�t͍�kS�AQ^X�Y"�P��U=S�kۯ^�K}"K'�E&K�4�� ��ހuT�Y*�G<'(�+��M.u�,��H�;~�q�Q����1�vWXn��]��ƍj�O�8IX+&���n!�w��cK�rCZ�x�/W�i�]��F�#��NN�œM��u6�TfN���0�'E��8M�nݻ����;=5IX�Ĵ���_-��Vg��f��U���۶��צηe�j�L�>3۹m���"}o��f����/j��>̆x�o��9��C[kןZf�;�"\)z��d��6�Di��#0�"�RYo>I�2�L@3�N��hfsb��8��#V��O�fNB|N��
�b��-:WY]��r^N�G�b�վ��N�J;�umUxV��\ˉkJ/^Z�:>do��>��/�W�װȞ�[<�����x�}�t�.�ǚ���Z��$��%g�Í������Q���e9�ϭo��;Y�����ؗ��kq˺@�AOw`��������k�ꋜMs��5~�Y3k��Cgh�9���g|~;!ko�&���t�Kb�P�W݋�D߷�ɿ�������%h�����4��6}��:��?/x�M�l~L��I��.\5��'���>��S�x8Zq1�c���� �.S ��[�Z:����L�3$C�<@L�������8�k��{��K''��1�/�9�(p)܆J��:��9�󭏔�,2��J-�q91��
�#/7�ȸ˺��꼤��ѥSJ}U�l/�����ڎ�1�l��ǁ�V�R�J�K*?v� 匥Y�Z>�=$vC�\K*��h��X�z�Ŗ�:�AEhUx�Uo=W����}����|�X�d6���
n=�Nize3�J��KOS��-��N�o�%cG��5���Md��-�Z��I��r���X2�<�m���h�0�	3�3#��z��.mB����B�/��$~��D=��g۳�=�L�#��{>W��I���n�dk /�r��vJ��Ml�2|��VM*2`�׈���[�2Tɂ�SME��AN�8K>�J�L��D��W<�uşq��ߞ��Zn��N��[O�f���b2�Y��/h��j��Pq��덵�,J�^�-����KJ�t{�)F��ו�x�BGEgM���F_'O�ۧ,�����)׬޺S�N�R��ߖ���<��6ܦ��װ'[�\�b�
�o��I�;�td��,���ڍ�	)j���Tͺ��^�{sz����k��Cܥ�*��S�)��5[ ��n����t]���yZ�O9�q�8�nP�|9-���n�_3ͻJ��b/G$K�)6*f"�=�����Ã�U��kh���������w����eX�M{�+S �g�"�&���N�����/m� ���z8L�{��ٺ�c?3��!�����W�w'�J���V�8@6J�M��yW�oz1rߪ�)�[,Э�l���,6�{ub�P�ժްF�����L��vb���w��@�==�uU�m��=s)�
^�`�z��M�u���ƥk�O;ڔ���]�-k�)%P�5n��%y��)�K^!��^�EÅ����{����R>��tn�;��GѮ��4ao�Uh��M�ue2w(�,2�"IEm�*[@��G!SJ!��Ӎ3���''���˝�mE��Eyc�����7���D���t�%�g��s�+ؗ�W���@JZ�M3��U��9Kd�^�*�2����5w�Ѭ�Qέ��n�Q7����N�8�J�k�[��f��$�v�ovW��+ZǗ�F�Mӂ���bIs��t�{��Y�ل8̸G dj�}��!�Mթg����;�D�|VؙgE��Lw�Y�[�ܔ���=����8��嗣�}%��`�������+ҨɃ�^��OY� �X���[��)싦�6f,0	�n�f���ox���y}����\��-��[<�A��a�~�^��@t���t*�N�-�~�n�^Z�w+$�W�J��r���B�U�-9�B�
�bKl@:�-�(��@u���xMEE���f�u�"wJuH&�^�ئ��i�� �<�I���[b��lHw��l&`M�z	��Wj�n��,�%��"�xR�-�ɿN}�"�:Ǔ�3䑗VЭf�wT�5�d&���M�5���/%I���aO՞�n�f�ۢb��߲;E�)l{��έ{֭��'=6��Yh�x��EF���Y%U�V����m�֝>��T9N%=Q�U;e���Qz���Afn*����=�uG�s���}��l֖�������	�F<5x��$j)��݊$L&M��%-,��}+��8�m=�J�C���L@VN�Cj ܻ�O8@�=T0���j:���Pŕ ��b监t�3W����|�U�3sNH�Cak0�ܹv&�����Nm�����j�E�T�Op���/i�X��'}C͟hVn����f��#�M{�3��KBe�pv�^��+�QF�R�5�Q��T��b�ɩ�h՝��0��$GO=4�"#��[�\�t���%p�n�O��z��]^��km�a�s�s\��!���&< �b�afYSH���P֨���}[�CS��U��7�Xnq�~�
Q��\�M��p��y�xg�,%��!L� ��ꡒo@˂�D*�1�dnf���]���bBw���j��M�b����z�Wj�`�2a�)i�jt3��j1Y��0LvU�6�TeQ!��f�h�Svu4m7UW	ze30�xw�L��D�HA�Y�lʥ�I�*�C����n9��HtOIr�G/�3����mg讖�e1="n�%L,בS�s�fH_�;U�24#�q?������0�th��s��ykw�'z� tATt�oM�Hy�a�n�El��D_�L4ol䊐�d�2���)�I��eG8��z�$AOW�S��wRM���5u�������þ���`�v�-��*�"^�οY���������m[���K�v��u᯻�kVEG�6�)�Í�$����N�5�U+:�yS���u�<ڌ��Wir.{����@��h��!T���	i�;�?�"_)��)�|zo�)��<q��ا�����X	l��M�-���y�b��_Yb/��q�u���f�����V�XF����P���F�5�'H�ֿyXCr-T�9i���ܚ|��7���"�?V������m��K�7}7��ُ����>�}�|�tmh�����,=E��{;����� �G{;-�+��z���D�'zi���h&]w�K��A���Ȼ�,霰��4�N
iQ�d�xf�:��7�[=����`��{�����i11<vζ^�g��u��l�`�e�. �Aߴ�'���)w�%I�*yXٻë��n���v�R��Ǘ�]����Թ��* B�Q�,��G^���9��.�q���cI��/��nЄwt����2�m�e�Zgd+������{2� &g����\ ��.1f�rO7�A�귣�1�H�gC����M�l��x�/o$��u|1p=[�:#����봉ܝ޻͎ʨhļ�=�J���ܷ��{4e.����q5cùV���&�P�-���M|c$�!�hΣ=��0Zz����->hP�>񸺦����,��|�G��%�X̥�q*Zf8͗5�Ņ�ywχV2l��Wo��'7Iݰ�3v2�brg��e��Y�
� �gn.�ċ|���rۇ�j�֘�Z���pt;������_M�ze(�{Q�E�=�'@�Φ�2����g0�P�6�Nu�ݧ���3��ܽ��w���C;�U�r�Ƌߔd����l,v�7�~�;�=yzh����F�{ff:(�TB�"l�Ϡ�ѓo�K^<2�'k�	��E-�q6�9��
�p���r�Ż�2�qL�o����1`K����<��.F`XS�y虣Vb���#�j�������;��YwK���	�yޗ�碟�g���o�O-
7?\
��r��=� �������R�VoU@j��O@��3OT�V��}� �Cv�<H
�&{]��sn��p��}�l[������"]9bg���K�E���сx��[�x�������yL���v^x@�g7,2��01�M�"��l����;)���L��^�K��ރ�.��j.�$�:��k qz��˗̞q�B��w]z��zm��O]k�_l��A���#}/�B��fMg]R'!Լ���'A�Ʊ鳮rF�S�5��:s2ʚngHL�E`L��֙��j�G�(���ZE�8�5@�u:�ʣ=���iOmG���Ad���>͞Vp>Z�]��%�)'%�N7��c�t�h��'�����2�]�C��L���q5��vE��=��*�u�Yw�Vh��^(]�����f\�n!{�E^n�:v�w�w)��L�\.:��-��/^ħd��� )���5�3LGg�8�� K�Q<��$�4sb'Fװ�<1�Q�.��T��q�
p��`���L8T"���GV�2��7��Y �
��3�_�C�Y���q\�m�#��r��d�q,n_j~�b�z�6�q������sצ!p����%��uc�'�Co�G���2�u2�C������$���9�&89E�Cx`�]�t$*b�Ud��׶1�����v3�D�\�����|�˔���O4�f:)dr�;�l�d���.�]h�˖M��"��D�:z��ȞkZD�;�0��=ѳ�;�a�}�5�i���OG�c�����R���~دִ�Ns���dg*:�YpǼV�"�Dq��Fp�-�<�o��)��"!�׉}1y6��s�]��U��Ma���/�;�i���[N�@j�+�p��g޴%��C�w�=s�&�T4J�2�ϊj.��Ǖy�xb�I��)���z�5�[���.�u����^�w޶B�psS��g�`"&`��?����p�������]+Ծ�ӔNE��~�^�x���%A�p:�˸�,E]�}Di.��N��'s�8^s�o*w5�4@Q7��E�J�´����wl!m��B�Գ���gC�Å���?�fޝ��jEZӆ�C�s?{MЁ-�s��<mU����fB{s�R��OMh���#f�/:���>���̜��p?K�lw�D��l��ޜ�S�0fK(�����ܝ��r||�P��L����T��3ʁ[�GgL���gU��.��g�� �?m��+�i�C�O�!'�(�OE��SZv�Ď�_S?6,��h1:C����t�99�V���W1�g�cF�B{�>Auv�ke�*e]�5����A?N��t�K%��oV��l�U.�9�5���j�[RE�(�	]��V_���S+�[V�E��a���#�x�1���ȗ�^�L�8�[Eʞ]��ߍ�8CIr���YޯZN���`�E��M�C �!��g��b8���d.u���N!+��l�㵭ys���l��7�dv9���);����fŞ<,�*�	
i��(_� ��Ī�F�zU,��ok�9�l �3�Hu��a��:矋>�@K ;���Y��	
�.���!�ˣ*k���M�c�;c�F�Dcq���vuC�3uM ���pՏB��s�Y��˭Ӽ�_�]~�/F�VM�YkF��<X�KV�o��ǇR|�zn!�PL���Z��a���1�2���
t�s(lzX\;" �2�������"<:���X�{D�p2J�ڛ�Vac����*S<��6��m �:w�F�ʗ�^�Pm,�vfbMT�Q��뱅�$@Pj�cem����no0�/�c�y�l2�{j�{7�)u����K����[��
�c:�J��)����olh�$=�o���4�p+';pN�t@X�8gDı��H1}W�.<|�<��Qc�Q�zd�-onzk��j��q]��-�֫(d��ބb{�y�a��?`ks�4`H�*>� 3i�{
�;������:k�O��L���{a��U�v�<�/�iox�j��e�ǅ�Fʹy�=���qZ��#�:e���T�>��8-u�Ahn#m9�T���^^�l:����=��r�ۺ5v1D E��ȸ��G������LtD���e:���![�����\�3.�as*ΥBH��ʺI�a��)�3��i+�����owmmbH�\��#���=��{J��AS�ꡎ��rɥ�E9�1SR��=:J�v���'�ޥ����&!ˣw[[�ʶv���F�Qx1dB�K9U�v7oQ=m	�t��A�,��lN��Ս�W=Ƃ�=<=WB�^�TM�XM���Xh^#}��1��)dM)�f�1�!8)�L���AV��AL����F�f��I��["tD3oz�F��v��=5R�i���c;p&�,eK�hYq��;�r3�Z<�%X�v�ݻ�4N2���Qx�-�H��:ӣͿ3k���W���w)��P��pIk	R
�H��k�ۈ�YN�y�]�`�RZ�>�N����gغ�uo��qN�1���)�ukM�����CW[ЙNQRf,�I��Q;���mj�q{�x[x
PE��ؔ��*����r5N��n;�d�����\�Nvʦ�b
�(1�$$ft�+���%�N�d۲� x�1��a��hj��lJ��Re�h�&u�Q�gw:�e�bӥ=���{L�]�h�4�8A�G%#h�.{F.���X�e-�TW(dJSЙ�n�da�S���я;��.�z�Y{+&%RF�$]esW�B�2� �3;j�b��g\���Z!`���ٵ�@�E.�:�n��[S!GU��ގx����=�x���
�5�r��%�h楎u��X�jr���v j�:��ޥ�ҽ��N�'hOF�8��4���w���R�����q��F+��b�2]������`N:4���ptG��+4��`dZ�o&���F��D�MiÑ�JW�8�뺬�.Kv����=�̰.��צ�xH=_�m$c��9��n9SZ��8����8�*�|��ХD�R�4�TDiBd�P�K"�t)E]\���D�d{�.\�"*��dDt56瞒h�y�CV*�T� >�S��F�Z'+*6��V�i�2)9D�O�(�#Ά�]ܣ���r9$��d;������YigY�y�t��eU����̪�։"d�^��L:Q�(����UL0���(E�h����d�UPj+C��dJF!j�;�R��T��J2�ܓ2�P��KKb�>E͚��y�:�Esv����x��Y�JZ4�BұѮ�)�Ӣ��EW9EA	�IÉ�G<�sD���l�"�^���J�3I"�iB9�wTH�U�s��)�J��(�MQ2��wr�r'A;��S��G�	'�Dyi����GQ��G(�l�p�%]K̩�r��N����DİΙU̎Y	$����=	�h&m*D�;��{����$T�T�h�2��-,�!���dRTRd�bNG�ܔ��ub+!޼��{1��5j�c��Zs��fVdչ����5���񃫞�bJ��)]����YX��fe,�s��P��F+֢ߩJ�C!{=��A�+���zfxK�)��(�ÿ(���ln�P\�WcUZD�;�p���E��n���ROQr��8��}�wKc>��SLUT�N]s�;j�^�����m�����#�������2<iިzK����9�z��u�L %Qjqz�ݞ���.���m�l�)�b`q�1�!l䊐�d�K,�	񴙨Sɇ|�z�7z̊T�;U}l�K��\���鄦)�>�~����H�V:`:��ϱn�qg�;ѥmb�29�3�чu��q���/���'=�8�QΛ?��͟ ôdr�ڜ��:�8��>ɩcDĭlw�w�tG<a���f��[�����}.��VVP����WZ1��y>����M=`N�}�������x[oD�'z���U�Оˍ���`.~��Sgq��01pR�l3G>M�ক��Jw�S�Z7�[=����b6�H{}@F���d��ۇ�Oͽ�RE��k�5�pa�i��*T;�ws�ewy��e	a���Ң��()���5-�h�Z���vm��Ȼ��
x�ݢ[A�=y����w吪�r�J8qY��D���zx\�D���I�{���j�p��,���Yaә�_S�p]}6�������i�O[��{-��mf���eW%�����=����N�߼��o��Ƕ��rڗ7JT �y"�l���EzBg(VDs��ܢh�vLS����)J'`�s�w)�"��=��|0���-3��t��4Awk0��b	�w1���m��������i��ޡu6V��zc��y��m{�Sv�9í�1�
Xf*a�D�;����t��ؾ����1	(��R�|��ܷ��n00n�ML���sm�pQ��)��wB�ܕVN��ۋw�q�傂�3�7o��=yJ4^ٔgQ}�WgSF��Xd�<뒟Mk��"a��O{z&8W�@gJ��ǂ�w���Ey���_{��*2w�A��iѽ	�nVv��k7��\�]����ה�c�P9w#l��Pn;5��)���8�a�������H�Fw)N:ٸN?8�d'�ˮ��7���U�m{�Q,GC����u��?U.(@SV�,{d����&���6'��ӵP)��� R�}�Bq�w��9�����{(EaN��Zl��o�~욧h�яޓ��8����lު��e4����7Ǫ_+���差D����um�V����ry���84r��/P�"�Q�r�L�����:�`jif�f�+��z+)9L�-�фK�z��m@۫�	2U�}V��Wy��	�}��	͡���9k�ma�4�h^3P�#Z�ۦ�V��F��e���;+����k$dǷ?Ru2_�"���/�����f�==���=/���\#{��2�L,	��5��֭!�q~b�D����07T��*1�d'��NZ����oDc�8r�`;^5Ф�*��P�NK�=FG7t[�x��������,�$fK*���x�)��9�c�o\<gN�9�cv��Z(?z:K��;�<oE����3=��g���7Es�[����~!�3FK�au���Fi&�g]�R�AA��g�p��̿2[e�)��d�
�-�|��y�A�lCV��Ȼ�y�Շ;0�w�Ý�f�(lR�qLp�ĺW��M������u�a�7��*���Sk���=MO^�s��0c�Lש�EE�rk:��N ��o�G�R݄)�T-9MU�b��E�tѣy�+!���c�� aݞ�繈HW� �멧()]6��qݲ8m�6V�X��6��ޭ�#���2��cl��R��]]Ak ~>��ip�9v��>��;rV��/�g�؛�f�,Cy���)gL>W����yt�tW�@w*+��Y�ϰ�E3��E�*`1*�s�u�[��	���r���\���fLI/@Ͻ�vVX�P�"�i�M�S�z^����O$Cݺ�r�@�=�:hd>�8s6�X�����oQŝ%��WQ��s(�x�Z:�Fd\;G<\zs�\��{z��;�r�𢵯t�{Y-ݓf �s���S|�9�~��z�?{11�gF�8��}�uMp�S39���;�u��kc��1�j&��fA/�v�F��E��'k�@q��Dg ���㼮��/^e3="���:36�kW���o9����W������;��ٰN����J�/���ք�4�����MdU�m�{wY�fq��fa��ĻG��V=�G`�l��>Λ~z��UVT�DWts��dI�j#��,Μ�C0���C���%�}��@�s����vs:�ٻ)���5)螚�}X���LWC������. ��꟱_]w����RS�A��P̖Qq�1�,6�j��A��Sd��XE�掙X/�T��Ι獶Ϋ}]Sr+K���.D���U73��� �T�<?Er$�f	�Q H�1��a�zN��m�=9ú#�t��<R���{c�1�oХ��u��*��U]�v�/��y��zi0��{w�Z�a1�Z�=�T�\uO>�wQ���&H��̭�k�1;�s�`�ͷ�w�N>S�О,A���"_�6*gs��4B�=�zm����2�Х����[��*�^��n��\Kڼ��޴���J�,n�W&ҵjm���A)�Ť�<�BU��r�g��i��Q#z���٘s	���SJu�R{��8g�q�[ڬ�2��w�����'���������v���I�ޣ��"�"�Ӻe�1_��Y���� ��5��{��qҡܪfɇ.i���X��N�fw+��r�wK��$�a���OW9"�K�}Ʉ #�Yᅙe^�	���][=�{V%K+������'�]�������e�S��~,�,��T�<�e��?BC���3�����Ö#HႬL�u�4��J7�#�4�uC�{�il��cÐ�w<����Mb��ٚL���Q��u����$2��t�:�6���Kҙ�AT�D��xW[6n��+7yJ�����ù�8��кu	�	̵�R�OQr�̣�������������ѻ�S9{ć���l�􊍴;�  _Ѡ�����������u;z��.�k㒪7�]��۽ͨ�4�����6;�o_[
e7]"��L"�Lk���+���V3:�=z���q�g�Oet��09���K���u��^�l�yc�}0�K�ѱO�;9���,!����n�w+�n�t��D�W3a5Z/
�~�M}��6��_7��N{zp"�u�:�}�~�M�L����x�a��]���̓����ft�H���T|w��+!��&�f'�+�K;b��5S�X��{�'�j���+Nޭ��(#��H��U�)��r�B~��v���!{�h�+QXAk4&^�N��IRvΠ�!Vp�ʾ�f���R̠�R�Ԧ=Mɼ�}� `���dL2�b{CY�i��3�m��/����s�qQC�5��[~3f�W�D�;�h�<�1hk��d'x��d�V[�ռ/��<	��/� ���Ęq$2gxg�x�צ�pSJ�pr�5��-ڭ��fVt�s��s��Nّ��Yˌ��rڒ/�� [~a�ف��QQl�w�^��w2إ�g������}��^��E枒BY=V��|���,�rZ��
hD��eM"8���P����EƉ�O[�d��X�L;��B+�K��|
�]y���
ںS�
��Y�X��o93�	�(��A�Egd�o�d�!l�#��]V���8)��׻�7k��_cXb&���[w���A�]~|�p�}��1z-�S�J����-�Dqƞ�ML���v6,[�f{\���/r����^z0��w�Aw�����ࡵ}6��J4^�Fu�n�:ۃ��m̭��d�9FA��F�i��c�,��Ƀ�{%��-��������oq�����r�K".������Zea9�9t����~��:RǞW��c����}�t��d��m�;s���`�K����C����~�[W��C��u�)@�K��F�/46�^Co&a���[-��T)��32�����!f�k��h�-��KT�m5�|���N�Ã:�."5�
��w�n��iQ
0�TA��~ȇփFM��.ޭ�F���Gj}3�ܿ4��*0)�t�������R���j�F,	}e��3�\��
���f�GL��n	f���>ӵP)���@��.���'�z^�ϏM�H�5�U�=� �f��j��6j�ݲ���С`Ƕ��p+͓Rʳz�U���)���m1��ޗ��-7='l�ۡ�	�7h�\ v��[l�:�7<p���O�.�ؙ������3�3�~=��Hݫ��S���Q�4���ʷӐ ^�\�,3-i��+ңe6J~yl����2�fW�E;���s����������+�b̽�d<�Q���u�҇�ʬ\ ��c<�Ș��.�rTN�z=���8��	����|ꋑ�̔�}ce^����^�c����Y}�;%�Y���8e�	Rx=���\L5�3%�^�� ��,�A[D[�mu�驦c�.��n���ޘ��j��:1��,�qTp��%Ҹ��n6�NL����4Hζ�y�L~�m�`�r�Y\��9EI��;_(A�Rj��sQ���G��u_m�vl��p���p��ޢv\�y �O�u���������/�a&�rvZ=il��A���2V�ۭ����ժΓ%��Ǫ��&P̜����ݶ�t�|���X�
���>��yerk:��N ��m�dp��Tݯ[YR�稙�n��H~��βa
f=
 ����,�������箦���t��'�Cz;�Hh�5}W	�t��CFs.�x�G������,��Ub�K���� ]h֪�*s9��j��[��fqy���\3�t��)�:a��T�i�L�E,��Tr-��g��\#���{�����n����Y*v;pw��*�D�Q��΍�qM���1<'L��z�9C��\u���<�6�U���jk�: ��y�p��pȜ��@��7	�y]7�^��g��_�fo˵�J�˸&�7^z�<K�g��%ぱ6���ڨ^%u���ք�0��!]eN4fM�$:z���V��:,!��{r��ң�M6B|Ί~|m&��ʗ��by�W��c����c��%�O]Ǯa�������y̽��Y�덫x�TΙܥM�f��e�b�b+��2�E_M?FųwD����j�oN�^~�pE�eb0<�Y)RA�Tu���S�k7�f�s��J��X���E�}41�R%��J��c��4�N��*K;W9.T�jJ1]f�rr��"$��Ƴ���+OU��� �y|��P�n��x:�=ֈ����uS;M��6�a�����r�I���`:t��lw����A�8/J�}�m�3�y�o��]u�.����M.D��u�����J�Fgb�ͣWև4� `�l�,�W�����=9���y�ؗ�:�-�ٍ�s�*��~������XN{�#�z�V�ki�ޝA�ü��<���Gkede�mb���In5�H}���ѐ4�8�N �z��"��C�i�%��wÈ��_�O.���۵�as�d��˫1f�Y���9�N �ymIԡ@
�!���LGM*ʯ6L9sY�O���::���ab���CG+ˤ�7��O�\,���ra
eРB�ǅ�eL�!!S�P����$�
�cV�IPM�k�=�oLv�[!Ίe�S��;+���2�2��E4�{2���~m�qon�X<����l_Uq���yR��!���00����A_��8W�<9��S���3)a����_��3��v{qݱ^��~�)THke��1����-�U\%��0���Hn�{�U7y�qnS�F)��xw,���T�	�	��D����!f��;
������T#6�؏U�hv+�Q���)�W,*�1ڵ�#�uLk�Y���^U�|��=��#�Ulk4�˔[t,E���M�Nٵ&"��SI�x_�@�Z9Q<MEMfqS���;TG_o���}����ErXl��+ �t�(	4�۝��p*ͼ�g���!hO��?W�uӺ�?3u\�C݁>�H�\M{�?Nl�O>ӽP�7S5�F��^���2)P��|\̅6;ϗ_[
Su�y��!�=e~8��u�!#�:Ծ����P�͍�P�{���M}��"����u���|��l�y�龘�1Ob�lS�N�`Ճ3Z�LQqu8�^��5��T�b7�MK,�3�p���
��K���|�oK�ޜ���J�u��bs�fdNM�Vlnԟ{ҧ)�c���O�jY#�6���y�<�ߟT��w�|-�VW�;�}5�݆NY�v_�d.�)w�g��U1|5��!;���'�4Yl4����<	�&_t��Q�޼�iSi�����s����ʛ�u��z�x���N
�84�)��k����V϶�]�����zL�ʢN4)��B�wc�Ǧ�[RE������2�i��!~:�<��K^�xU�P{:�;(�������8DB��駷�崞�9mK��* @<�l#e�8��ԣ�Ь��ݸI�n�s#@���.�B�T�[�FS���/^Zgd+����Du��<�{ǆ��oe��a�k���u��kk�QT)�	Z���Mm�ܫ4�l5�R�s7��KG�vWǷ��b3LpL!,�e��i��%C�2I�x�8��Y��&�C�.�LU���t��˺U�؇���Ҧ�;�[K`�8���y|��ڇwh�a��[׫�6M�����h\u�^����)�6�u����G[�����U�F��xE�ʃ�BI95�6�G��+S�[oٛ�x������p�e��n.}�d�xșT�����dɜ묠���Sd)�8���s�,̶�c{��(�}f>�^"�')�D����v!݊l <x�[}/�k���*E�?$��7t� ���h��3.���>��Э���{HѶ���β���4x9J�M�I�VeL���کzd@�,92��4�n�+d۽���o���(��k�>�K��rgM���+i�%�w���#��]p��
fMͲ�VV�=R]gRxnd��.�r�Bm
�:�ЊŌ.��dL/���oף�p*�<^��I� �;�qAf2:.�-u' ��dXY�NR[R�El"�U�rih�*(k�L��˞��l��T^�Y/:�x
���v��64���C#mL���9��6���0�x�%�)泔�O�T���Z��Yf�vi{��I�d6�*-�q��so�W���-*5�Mr�ʑ
-t��b�(C�gq_?H.�&b8��.E�O5��Ў Q̉3eZw������xaK��׌�g�մ��sGV�^将�,FX-%S����gg�&�/w���LZ�Z޽���&N�h*@*0�42v�5>X��fo��LV��r�v���I��ۣx�3�-����N������<-bk$�h�ir�����[�O���H��ܓC��:DOh�{c�pk�|��\��Se#0D��9V�-��o*�7�<�R���΂[�#�
��;�����62�����yju�"�F挐�|�et�L�b����ԙ\V0S��5���P��&cDW�$-s3��s`�"����1+������t1X��V�ͧ��E�!��E|��s�(���ф�3��t�xº�[p�&��X�s�/��r=��%c~zGY�k�J]SBS�iH^���Ms�?ι�X.�;/)W��g{+YGN���8R�)k+XB�ݛV9(퀟36�7��Ҧu�"����i����|iN*�k�5N��J��b��+Ŕ,rM�{f�7r�c���B���F��{��|v��9=A�VkǼ�*I�'��-��'{[G����q�$��Z�r`={6'3^���0
ưs��Q�.L��sM�͝كF
ᴝt�hPCv�45=k��r��;!;��5c������`�kc�]����)��Z��J*<�}���9��ӹ:�S�R$���%8T�����%���#���PE��
�Mm6F!ruw7"#�1u]tQh��5��Ԅ���B������m
��P��s��"R�1�t��(�C�,����U,�E3B,ÑXhH�>2<*�I����WBU�����E%[��'$Q
剡I�*��\RJ̙�r�6T��T)�C�y�wC*21Z�,��օa�B�"��̄�S��a��nQ9�QH�2��brwpvt�H����PF:���G�dea\��505��Qβrp�'q$T�H�u��10��*�fH:��9�(�^g���ė��L���E
�i�5/�t�E��39R���y���r<��3���dR)*ID��畝Z]��sg�W	��7'R��'*):��0��D�3�st�V����ey�f�!+J*�в:yᄪ�4S#h���TD���p�QeȌ�$/=�9UA��8AP]F����������������S=$}��"Q�����j<����o55���4w����w��x+��G�&�=0b�q����,z�&�sd��Ϳ7�"��zR� �M��ޙoLpR-�����-�Y���͢�y+����q�� $����m��a��v�ո��;�� ��j�R�|���z��M�i���5�˻�[�7�Ry����Lp���vua��Ϥbk�N�.����GGl��8�o	�n�l�9�m��~���SF��T�K�c�,F��X@p�ыЫ�k��Y!���{N��gD���Mo�g��;�1�[���TDB�=��ȏه��FL9�Hͽc_j���Fv�NTsU�.���W��.:ۄ��Bq�W]s�e3}0�ff�_ru��L�z��<�b3�+;^y��X	���>ӵP)���@�2�}��n���{,zm�DM�=��و�5��W=�?���߱�AY���\�B�>l��TٽU����[�9�m�t�� ��Vn�U����"��FU��׻(G���E�-�d>>��x_�a�~���,�0���]��d"p:��KFcוom�� cuC���4��ңed�眝���mbQ2�f�`��I�t�s|�԰�*k�f��d�����7�%j���<��t��&��u��׭��f��/#�z�XT�A�XS�@��Q|���9|�'*�������6d�Kv	H�Yp˯����*9V*���:���9�yދ7zjN^��=N9�����K��΋}�.��{�=;v�t�ؑ�,��s8+� Y��;u֫�v�ZĆ�6�]߱\���!��e>p���p�|ꋑ���}cA�A��{u%�V��i�f�δ!�������x'��{�)�u��[1,��)��\B	���륺�Zu������s� �==�)�OM�Y�*���W�=t�]E�1��v��r�y��0:��D��5v�8T�"�ˈ#��`�x��FЇ&�����
��۶G�Z1�7�b�ܱG���q�Y���R�P8.��,��1	
��筪i��K�-cFu@��U���������Ǥ!��$�`�]]M�Ϲ0�y�@g*�1g�%�|:�]h����z����<ʣ�~��~��p3�g.��Evt��uU'��Ѭ��PȰ�Y�9r��/^�"�E�Ўp]Myr�Lg��j#4rѳ�;�a�'��S39���;+_w��5�6�Z��%�ܱ�h�͂�n8�kǆR��q����-�3.��/d�+�燺��J�~���b��y�M��%Mb�d���v
>�^�#��k�^��٠�*�_`�ra�gm�G�9���<�	��Q�5�׋� �2U�͸w����ͅ��7oKe���K#�\���U!�{+�����}+
4D����P�s��9�8w���vDo�3����0&#��O˴��^�^�G�FѬbWP�}�����2���y�	�{���|��?oc�7\�C�`LR�鷣)�v	��O���oϤ�åu�jq��3Fn�e�9�#�|E��&�g��B��\��a��vs:�ٻ)���ܶ�WcRm\;�lĎ��rSZ-�����~��n��ol������4��n��,���c�]�E#l�]���a��"�i��$k���/PfVm=.��:#�0�U��.��~=.�SGK�Y$��9�c4m��;�������`������,�b��==���y�ޚz�51o5��Ɍy����$�(����`���==�1Ӿ5��zu}�K��|�ޔ�5I�=q(��;��C��ݽ�RE��F@JهN>S�#���H�J�@�D�lT����hh���N�����u'c9��ܗ�W-�"�B���O v�A�M�}}�(�a�q0-g3��0^�ߛ�	(M��O��?�t_ra�@��,�,�*i��j�ɡ�6Z�j,��W��=z��}y0ӽ�EE%հ���1�-v�K��g��T_+˖�s��Tv7�d̓��xiݫ�Ygc��ze����z)3O]�[���g#7�ZO��0ү6̻<���.="�lܙ�N*�۽m�hzQ6M7�S:$�a���n������=����1��C����h�~mj��E4ﱑm�g��?�FU���sf}��!�L��*Tp_�����q���t��LJ7��8up������]��U��#��� 5P�t;ʕ�ދ?��D����3����я,^��E=DT�y�x��ȗ환B�y��*fxw1�p�C�j��,���Hu>'��{�48	���:_�*4��R��OK7�@�e��R�+������m��ʠ��F��\M{�?f�t�Վ��{�]u]Ȍ�U*�"���0@]�9�zЦ�ye���EOH�3�x�.F�\2s��Ew:��͔ͭjU�l78�LLk=<�+���G[!���,���}0�K����C�<B9x����ps{3��@nA��9�j[�7��^.���]��L=���
��� �Vvn�s�UJ�['���s����4���Lv���Rʘ�����Ӽ3�9�}�K������fڛʏ��i� ��:��1��/��4��2�!;ǯ��=4Yl/�z��6��C�\l����RCH��4��W�a�o07R���V��������m�[]��#ރ;ή�w�£{�����k�\uq��ą�+T�eoh��+�RCbm͗ޢ���'sv^9�����ٱ�Y$�Ԯb\H�\9��C}���p��8u�G�lŊ%��m���˪ܾu\�eѰ7lt��!>4�NC��N�ju��t�C;�}���QEݽ7�����N(�e�o��3�Y�jH�W�-�e�s$SJ�~7����n��U�ĉ�}NK�{��\��9d�[����O^�[R��J���{^���)�߿e���1�m��Ag�)�"9�t;�SE,V��Q��p���1������Z[�&.-�ɻܘ��M�ݲᯚb�Tʒ��!n.�ze�1�H�gC����Tݶ�6�X:�=��z�edq���a,�q�5ߞถg�54��mB��T���oR#8��N��hX���m��nQ����˪�1m����ܪ]��y�S���E:}e��-��,
�=��Obo��j0���='@Y�уz�SM.�� g�Y�ܼx,�yD3�ɣ}=�T�h�s����h��W����5�l�'xv7��)��uޛ���TDB�=�����s,�H1\�uu�Β	�Cg��-x��N�@ԺK���8�㭙	�u�<�DWL133���Oޫ���ſ�ąj��*��b�
߾۴C�A���4C']�@	��� �dp��&������o�r$ye��in��A��W)2bt�>}�	����E9�l�Eܱ������A�6(�Y�>��cnGv)�t�l�`W�Sm��z%ZK�_�s���<�H\���'����N�@�&wC�qd'���<��i1Ef�UaV`u���ja�ا����q���5,��7��5��������k�n��|��(N�`��gpu�vt�y�r IW-���:�p[��6�|���O^&{m�6d8�~���U#ka���&s�GoEzZ0i�ʷ��-������ʽ7<EJ�q����(�n�N��27;z�i�/g��:Mc�m�[�m��/:-�u]K����t�ؑ�,�ng�;K�e5��X{tY2t(�2�wxk;)�����)����f<k�:�$m�;_m�:s �ޖ!I���޽�������L�HL�l	��{bzOQ��uKfZ[e���\�2�"1�l�rT�s6�:(X����b����[��U!��\uKv��׆�˵��WD�~�F`�:�L8U������L��#�o�����<�Ԑ��X�>o=(E�&���]��m�N����W�B�:�Aw�qd'����LAs�SNP��csaj����� E�U��(ݯtª4���z�y��*��'S6�5��w^�]/Օ�9F����/�5j����6F�L���0뷇M<���q�nDbZ�S��v�e����y)��Ih�0ۣN�B��7��r�K��ʉr�w���k�1�0@u8�Y���~n�ὰ�ݒ^0R��n�gܘB��9T��ǂ�w�aА��]�H�S]��x?[Չ�Ƕ{o\��#�t��+��:fS�yt�tS,��TS@r.����CO��Z�ĉ�3\����)��yrʼg�����n��q^�����4�fy:{>�u,*�6��݉�9��ې����9��㈛ǆD���G8[tFp
ٸN;�D�Aۺ��6��G녏�����hwe�c����3M��NlZvfc���)�ɑpb�v^mI�N��RxklP��ǮzE������nV=ʎ�5��-�6���&Fi�����j�;{��l9��]�~d)�{y�Y��Ё>=sņ�n����崽{���ːZ��r9yٿ�{M�bpo��~M}4���Ly���zpD�N��e�.�P�Ƙ���[*wvU�^��d�F�짨3=������xÝV�^]u�.������#K�GVU-�sG?>�a��i��pSH(�3�_l���;�l���}ӽV��-r��/����H�˵�)���y��Cncx���:�<&gJ��V�fQ;.��4`��'�ۭ���2��#�$czJ�#��i*Y47�,;��D�k��9��qb�m�j�m)��S�ݷ�c��cB���-��qf��x^���4>�F��/ٻ��}S��a��V�F����~��nz]��42��\-,�-U����Bye��������$](�	_�N>S�#���H���i�S;�P��-^M�/�r��f�h��%B���aN���jH�jP�ӆ�-�A��1D �T�X���5�b�XU'x�:⦞[q	\&�e?i�O�\,���ra�@��,�f)M�N���[�#w��U��k���W�*������襆S�vW?6���d�r���%�TnU��ݼ���.�ϙ,%�;�4��]TT�Q���B�gL=�uM ���m|��nت�X7o��-?���4����΃w�J��V��o��U�Fmv�n�.��W�(�WS�28�W��g���?}h9���_��P<w�G���O_�l,���S���w��q���mg����ӿ��?��6��Q���t�n'}	�p��y��DY��V_:&��py~�C�� r�p�w޴)��}���<���)�aj}�k�?�N���{��g�/�ك<��˱�L*-<^��N_v�暏���V5ْS������lV8�gfk�E�y Jfv�N?V}�Ͻ���=��&��х0����G�:�%��%����JZñ��4�q�9aǙ��n��$�~�<�[pN�}&&�9����u��[͔�z+�1LS��x�,����R���z_:L�
�p)�`�ɩeY�U��w���q��R��bf�(c:�uN�YJ�lݥ�X����s>ƺ���|�4��0V�}�RʼLOhk;�;��:g�6'�WTGSsul�<N2ݓ�����}��m{b��ŏ��q�1�zb���x�	��i��YlUu&
���
Iʌ�'!M�]A8��n_:�f��3�g�x���N
iQ�{%;�N��A��V���;E�'��[=��Y�}�o���s����eq�-��ق�eD�-�6��D�g9�vK�;�1���e�	RxEʞC�OU�>�r�OM�������
�D^�2���vNb��ͻ�_m6�#���y�#��)w��a���ض�e>�,���vB��|E�6sp��{qT³��O H��}-�l�RP�-��oKzc��~퀆�r���ɫ�VԆ�1SZכ����c!oq�0�P���ĸ䡩�1�K˕�T���t�Ou���jK��m�T�Ӽ�N�k��4�Tī=Z�ϴڛ ����vf��lv11��ʽ�1\��i1��p�m5��g�I����o;��|3�îH�2(+vP�Ռ�eAE.�)�s OpN��f���>��&Nqo��P�т�C;��Y��m��"���v_���]�єǪ�7[�Lp���z��P>���ߊ��2g����e�&k���n>b/7�_��'�Ѹ��h��*Zq�tLp������ܼx,�wдB[��漧㵛�TlsE�Y���#%�2�������wt�Eu4�)����� �=�����b OS՛�w��ԹHu�PU��!�����.;�-ӄ^-ܪ��L�LW��(���,��s�17{�?������M0���`�g<2�;U���@�.�w޶Bq�[�4A6�q�PCK�Wn4�(����ͿH���@��S�tn{i]8�M��dL2��Z�i��LL��/˦���-^TH~�q��wT�oC�w�޹'Ǯ[�����zcpc��5����:y���F_f*��&"�Swq�Q�xFou4�וo{�"S���02֛�"�F8¢8m$8ME�i#9iؾ/o�q��d�8�+z/��/�b�:-��^\����&Q��atw]z_��e��X�͸m��gE��U�C�E�d�w����^�3�=����s�x�z�u�Hԣ c���%w�_����8��JLcf��!Klt��5u��d�xp,59ob�j���,k�b�`:��0��8v^e��\�+������5���u3�2<D�Eۀ��垃k^efU��-J�y�� ��0��NX�=x�ɸ��t���#B&N�1|���f',�&k 6%gj�83nu-N�V�7q��$ɚ�ܴ�ڗV�*f�Z�:VԀR� Ƿ4�
nA:e��g��Ep��`�?[��^��֌R(.Ab��_)Yn����yb������Ռ�G�SZ>0�f��MK���*�����i�|�����6�a��4Q����������v:a�e�1U<矫>e��׻��}:S!�p)Nw꧷U��@��2��+#@��>���j�6�
�-�Ƌ�2V*z���w���+������#K���Լ�li��saqb����6�����0���Ȣ��Z\�jBV�pQj-;;\�#��=ղ���R/H��ǌP5>�����%����Å��Ͼ��0�wxmڸ{����:QZ�q���M$�%��󝊝u
�K<n���ϟ4� 5\�/0dſ��B@]zǑ�l
���u*�P;y���k+��):f�3h�b���9>Xmt�հ�O$��.�4l=�Z�=d�9[b��ۖ��S.fWp��(��|-n����f	T^�h�����+��#4�h�\hȵ��:ء�,&��٬�\���,�n��A��a�Υ��T�
fSR��r�e���`�z/>�UÅc.`Y���>_��8�]�[������.���2�M[�dD[�{S��0��U��஼M��y��9�e�[�/ G��&�bǇ:9i�{u�pה�1��2&�Jni�*,q�!� 7������_U�S{9��T�n.�,����W��!qހú��6�ɿf�e�_ .Q��r7��ԙ�\Z���u�U��3z��x$�T>m��gX�^m).���Q3&�l�3K�'U�O���t�A��� ��CtCJ~�:�g�]s���:e�v1�"d�!�v�r'��ф��ԑ��k8��A�����k��-p!�g`
�*K�+��;nK���3� e�%_+u!&.�v��{f�a�xq��֐hw�U^�X��9p��QH���p��$YSqێ傭�\ �2� �[q+]i�F��/s�P/7�g�n�_2�kBY��$�G}���KU~<������B3,����bcEUc��$��� F���:��+QvT;��1�3Qw�p�(F9sq��ե��im��\�Y�;B��*�G�ŷ�l��z������C'�SN��Ҹ�2!j�A�%���5�"w7�T�9H��o�/s�d�@�e^¢[w�;���=ڤ��M8ҹ�ߟ5|����/=��������,v����$P�hH�&gm�-蝡yZ_����yH�oO��G�~(�BIap�U�WB�6�E�]2T5ȼ�EK����"��8U�9�$q%��%�9�sF�I���b�r�M��؈)�$�eJ��VH�� �=H���Έ�F�nn�kB��ȃE���r�(�p��PĄ�Q��W=�qȃ�ЫP�.DVE!��R2,�*3�������\�0�$��Z��M劬�Uf��1V��s2��r�D��t��=Ye�9�%�E(D.�+,RY;�A�!I��
'KbI�̙2�������A&dh�R�+̼��Us�OT)9(��d���M"���P�˔E��QU�5,�Qr+BR�����L+���[
�璫-B#10�U�&F�-T���+�F���wc�"�,�(�k��H/wrP�X�`Y�U"�EZ��\��"e�y.�F�t,�Y�p�J��Vlʨ��B���D��\�����z�rJ�*4,J��~>��؊yW�k�v��;�i��1�p�6u���s=c�+4j�v���/G�5���my�t�>�[��rq���[��.����t��M����S`L�[���x:��<�k�Kl��p�pWlNwSuZ�8��Qw޹�]���k��LGjiP��`����U!�.�����5��]f{LZ��`g1�8��O\�*NY�	�`�z��qQ.�l�j|-���F':�t��44o%@#
2�9��!���L!L���=�f!!S\�`�O���u���]Y0�ro��GO#X�y���l�6�$�`����o�0�ydr�1g��]尜![�ul�G�|�r{������I����1��j�z�:a򙺪��.���e�ʋ׼x��lV�s��gU���G_���<��!�:�Myrʘ�Q!z9ѳ�+��i��k��:E�h�7��v�~��UL#�;����D���6㈖���"vx��8���#8x)yM�lBuuy��{��߽�6D�l̩"!��<H���?.��v��ߌ�؈������|L���)�t�����Y�S����/m˥�;����fa���kfչX�>_���ᵿ�f\uῈĳ�K�Ț��2����jm���
��:x׼#�U�&_M��EنocK �9[u��� u��BK�jj*�e<���;�����[X�3}��7�z\>[#�lP砦�}wnkg�]�s�26���:|�D;�Ž30��\���f��,ߤ����/�������SN�g�1�X��?g���a�,�//��GU
��{~l����T֌=�_M?FŷtK�l���[�8�88=�)��-r5v�7i��f�9��G`1���짦h3=������x�����Y"Νlvޘ�q��6���+���q�sB��##�ngy���3��@�������t�91֝E�L<�ѱ����j�{�|]�泥P̥���j��k�t���S`N�ֶ�KF�j�]V6�g����ʣ�!n�h�����p6rɒ5(�	[�|gs��I*M�/�uY��ޘ�J�D�/\�����.T�б��ߍ�8C.Y2A�R� *�D�2��#�~���H��}�kx���󹟽���{Ӝ��'�S��O�[B�.��&\ �b�Y�yv�K�E���7��sd��6�8+�1	�Q�%4��1��C���}�Ges���d٦�{��4@�ñp��?z���},'���)�A��AuL�Q�l�oG,i�gT>.�=M�yP\k� q�f���aWIj��v�\�\WN�R��T/t����\�(MW��ml�RՁ�2�F����!0z�H����B-���q��B>���I�sV2�}մCVs�%�^�`V��%l6�=�J�X=����V���*5x������vf��Ʌn=��q0�hgy�1�xr:�!�ǝd����h�pV�5�[�$�*3k�F`��S��}9���.TѴj���)��8w�u*�Pt���^|�f�=y�-��X��њtI��"+��@�s7Dg]�M���}M4̦'�S��E�����}�r�y��.V�X���{'*:���Ht��j�zfK����#����Sc��.���7]"������s��������Ӊ�qj����D�-�!��w��i3P+�T���}l�K�o6S<���gV���O�nZH-M+g��~�����S�N�`��^��KdԲ�ު�m�K�@���wM�R�Q�^��`�j���H~{��4W�\�}�~���|�i��`���Բ�b{C[�๹+����Y�Y�����}�K�1鿅���1a� %a����I���~�^���eCAY��iJst�ٞa�ˍj����[�Ϋ���d����s�!=4�N
���N-�p��uy�	�Իيp���{f3+:-��߉����&t&W��k������]U"�WM�L��t�+��x�Skz�{Tѯ$��],�H����!Jc9'F��*��s�;�^J�v�S�B܃�$���8�m���R����3��݋<t*Ŕkٚ�PS�Z� ���+��V˃��w�E˶a�N��nO�)v��E��)TE��0k˵:�����;߉RxD(�8�M=�sr�OY�j\ߩJ�*����c�kn�"��eDp��ʑE3H�s��qC���&*X��iFS��Qy�h3/y!vL�����]�l���]���uLA0�3�P��*l]V��zc��m��f�z�1��z�˖��Yd�¯dȾc��9��>�< ��8DAw�3���5LA=��k*WϏ�o���
�̫-��lؽW��Ǡ`+�Z���&8,p�Qaݝ!w���3�O��$�o�'��Gz.-��K��}~�F��Fu�fSvu4h��M4�&8W�@g��ܽ�,�z4�Ru'�p٭��}"�hG3�[>������h�×��+��]�+��L�(��P9��z�Ο��Q���W����s0͘yh��6���Y�I;]��Iq��'�u�8�+��s�P���ׯgdG��W���貉b1��;k��X��N�@�&�wK��-}7]35ѱSWݹ���.���?6�R(�Lp6���o��NB��0��z�uk�&��~@m~�s��tB;\�b�s�{�i���o�A�B��Q�����'��r�N��&�m9��9�Sf%,th�y�f\���>$�ԅr��/fiV�R����U���R���G���3E�v���j�uE��f�u�-�NQ���	���`��`v�,�i�T�V��y޹$��q�>οT��ǯJ��Ͱ�3J�d��>�LM�:w;,��|t`�7g)~��_Ep���6�ȁ��~�`i�02�i��/clL�ɌgIąӱ.'c�'d�4U�-��ދm��1y�o������N�ݱ��bg\OkW(w3�T��p��i�c�Gp��)��9�Π�S�f���zl뜑�ee80�[�&�=�����v�Lu�
s��웙�R9������(w�'��{�)�u��:��&�ͧ�D��+��I��t�ܗ��Ñ�5���L ��-�|���b8�W�C��'����G~�Ȏa4�I��W��:N��:2Kn��N^eдOj�0�P�s,�O �|��*%Ò�Ŏ��sy�6���pH���܁��kdp��-�X)�_�ra
]
 �a�Y	��)0�,�iYR�qw�{��z��c��TӮ�=Տ��!��B�����eϹ0�,��U�W����Vg+�㩲�Ț��]���1S��_�������r.8�+�>M�����O4�f:�=�$p�peN��Nm�Ə��=^D	��q*O>�C�8N�7�G���g�t����C�\)*u��m@I�����
��rU�{4ۊ�n�2��a�.�����u�X�T�mDY�m���w�I̖u\�#DZ��Nc_%���g6�d�d���m�9��?���d��y�;�S��E5��*3�H��9f�����}���Q�T���<��H~�'�f`'�ީ�����l�LA[���m��)'k�@q��qU�b#���$R�°������x�~mS|%��fzA��tu�_e�F�������ܠGF.���Vnv��"��n�J�n��}�fB[t={=s�DC�׉vչ6�*;�6RUKݏ�swh�o���ا��m&�����DWts�������͒�>=t K���oA���tF�블���7��!�Fgl��Ș��Z-�����~��n��c͔�[ӂ �.�z��T��D�Ѫ=��8#�#-�7=��G`1�����f{��w���x����3w��Ц�fkj8֝!�L�ͽ.�SGK�,21�\F<�t�]�ǚN��lg�8"��������j��9/=OXT�����c�D`�f�.���i���?����m0����3��(�y����n^���?{��B�Sϻ��p5g-�"٩F@I�-���Sq$T�t�R�2��8n"��W~�l�9�]��.�EK�R�+� V�#����ڭ��K�/vWoRh�ƻkOA��T��>c).sot2#���N6֫N�M�57�آ^*����r�{
|�<)�kVu	��h,Nᾒ]^V����Z�S·]���#����Wxק�af�<�tS��
p�\�d�ԡ@
�!���5P�͗Gk&"�p��Vr�����a��6tӜB	=����R~"�Iul��R�PW��h�ǿU�5�Q=x[�Y����H��S�x[5DX���2��_��s�a��c���������Z�ܮոr�j���}�!�LW�xg�,%��!L� ���U�yR���(���������	��6z���뙺���g�ǎ���T��d��3�=�lW
~0gt0e}���.��^:{y�j��ѹ�G��RΦ���.�",y�ߕ<;�p�C�j��6��5��h;h�0�7�0L���܍�QƇn��������o�����f33����^-�y�yk>�����^jW�H$u�D���f͐��w�R� u��s�����+���yM�H�108�5�W;���y�Y�5z�<�~��9"!s��݂s�S�6�5�ʞq���}hD���]V�������,{Q��S��yLfc��<-��.��g0W�v�X	�MK*lު�m�K�@��w���C�0m���[Q~��D�G�7WGo�:��D́�r
��w��h]�t�+*�םSn�潫wl��V��\�=o��8�i��.�[���(h������W��M>213.J�_S�e68��`�X�l��-�g:QmN{���f6��:��t6�G`[L�Z�������_���5�usΛF�N�>T��0S`<2&Y1=������;��\
n�>	W��T��m��/��W
}?C��C���c�i��k�J�+�	�k���t���՚r��Mnm�dUoމ�NoU�zl�ʛˣ`n��g�x��M��ıl�p�cb7/z��ɜ!�\.S��fu��F��g�����La�8��&H,�0���c��ͱ�v��R��}�i�S<#��l���qK�*֕<�(駷�f崞��Թ����n��TY�T6�7� ��+��eR!^���9��j �LT�[�(�}*���%��3��-��;��������;#��< ���Y�V�L4GAChA
���ޖ�� m4����*���n"e�h�e�Lu�/��Ǆ�����ĸ䡠z5��9I�����36���GLMq}~n���3���E����}Ɏ;�XAw�q� :1w�9��������z�rE&�]ò����c(�{fQ�E�=�'@�vu4h��TҸDpՐ�S3ù|�4E[�tD*�s�o��5�K(Dӵ�Łmk/R5>��`q
��b�?�~�� �xnT��Ӯ���Vb��]�k��qAeF�0;���>{��Q�~Y��L�|?���k킏(���eM�F>��������p�(M�޽�X���M�&�������u�얫���q���'xv3p�|��Ӯ��}m4�f`�ʺ����#rv���T��t n�<{�xe�c�X��t
�]%�[p�~q��N;�^�Ptz�%��m"C�k���0�ͳ3Ł/����51�d�uc3�O�&H����m�M�gl��/|�p�w��{>=6?3ɥ���Xt�������j��U�R�#�V��z���os��v"��n���J�L�9�m1�����y޹%�\�f}�~��-�Fp��8�Hۻ<m�NU.P�I��{�34���N�[aR�W�\#{�����{m���0����d�Л"^�r�ɼ�DF��δ9��̍r�읞z�*����������o�˯^[u]�!y�(��ߍ?{��nSۛ�,�G0ܖ573��A@l������3�=�O�-��{A�Ʊ���+��o��J�ٲ�#~�24mҏ��^V��9gO�>͙w��%�2�yYԝ���[�#�Y�|Ӆe��; ��� �4B{�x�uS��C�͂x�,��ap��羓7n�[[�&��}c����G���0��  "��個�v�2e{q�e�3��̙j���OƇ��P�V<]o����Y�T�3�m�^��_ܸ9���;���Ҵ�N�U��5ג�ow��E�9�����[y�*"K���rD����!���7枺n.��\	���a¦
�P<|1�|.�_�ȧ4�����>��d���SS��
���dp�n�M�aN��Ϲ0�.� s��l��O�����Ƽ��S��y�}T:b5��TӤ!.�}nO��l�7�ō]]M���R��&��Z�jq�����6��d;���B�#�h���2d��ٌ�F���vtC޷URy�{KRn��p�-��;ke��#����@r vK<�����Myrʘ�Q"�Fh�8d[��/r��v磟�/OurU�[@�_x����Ǫc�;��Y ��<�8�����!�e���b�FL��lv�AU ���N;���":F��F�%�����PpN�K޿l��֗��ï�r��]�U@m��8ϋ��ƕ���ǮzA��~:�.ѫr��7�+@g�3�OYӃI ��Оc�-�m��I���=/���l�4��l�y��|Ǯa��1wF$݉S8��wq���&s3H�oe><�MJzf'��^�����ض�}��Z�J����������)Э� ���$C�w�`���Vˊ��h�ݧ3���Ԧ4@m]9�X

�*6�ɺB:�6щ7��F���a����F�׉g�r��~orrw3A��~���R��۸s�((1ڦ���3���
�^g0��m@����u�y�5X(�N3۾�B�sob�=�l�^�<u)��Gi������Nn}� �Jڴ��G�B�ɼ��Y�� Ag�&�w�.�dL��e�x�~˭���eA��=���b�5S��gF=�:
���1�&�&�	�w����2'V�3�/u��fO����v������MI�(�� ���!��������Y�
�yl{�~~H�m�+m��S�3��1Ee7v~�W%gw���'�Jiȯ]�zT�o�N���p���s��,<�w(Em���� @]wѺֈ�V�j�-��JBl��5�pd�v����wid%F� �T&ǈ�ٶQ$�03��|fK�.�{vd
�[�[�[�j\_.B.�Ǻ���{d�`Ҹ�vcG�"	��6[9*7&��/�]�
N�7�[�Y-�y�nœ�m?�Tv�tӭ� [��	�JhWb�b�c��`<��)\��*N���841�홢��r�5�Xg��b@F�Ec�M�E*�q��61����O%��TM�wW�lظ�p[bˠb��8� 6�M��gs��l�6��|�=�؂��3-$��a���e6���'u�_r8��ɺ��^"��<HGWI����ۚCT����oW��V)����
^v�Y��E�Ke�u�Y���� ��f��9Pi�*]���ª���6�4,C�ͱ���U�U�+��[�=��\?5�7�֫r��WO�x�v�Y����݈+��L��n��Kp�#�x<y��{t������[��b��dE�+�LIa���V�;d�[�1���@0'|^L��D����8��c��rĽ�$9���k5������I���`���R�A����1Mea;��z֍iϳL\0�%��>�K$϶���밁���33gr.�or���&��ʵ�r�3y'��μ��`��]2k#�y�Ҋ��;�t���ʾ�(�C�/ �&���f�$�,b�/:E�YW�s�}c�`�:����Xl:ܡ��)�4L�Hf�ۏ#Ҩ��`����J��lpl�IQ	K,�ώ�]3��r��0u��s-�ǠW3$�1��w��#p!�C��~^��׼hHZ��%��T�䜹sC���)r����X5͡����p*���gL���faTz�Ў�Ym��Llܑ��t���1�z��^|�;�ûڑ�-���Ȳ^�g���w�8���^�9V�qR�pgs�t�֪û N��Zs5Bվ���5�I7D��a�a`h�Jk��9��=*���4qh�c1>�S�\�7i�޺'��ӈ��V+��˷��i9\`�gi9eDxw��H�Of���@�s�A ��CB+DV�%u\ȊN�IʎC���;*�E+(�*�!P��=D�eH븑+C�&gh4����XW��'�D�.T�X]�U��$�J�XZ���IДT��N���.BVPww'-ZA\"#$.$$I&�(��#��N�p��Z:.z$J*�!ffKup�(�U���j]%�z�t���T�W�wwp�ZD���r'j��L��!��N��`Y\JҒX���UMY���#�I"wp�*�R)3��6���3:FI�	f�U�$B��"��I�)mJ�*�*2�`�yui^aȹ�J*�SPȢ�L��+�f�u+�K���:��dADq$�34���Z&j��L��$"�reP.��r���TҰ�KR�(E5ww5.�N�4N��eU%�m**#h[2���!I������b�QAFѾ<0n5/�5�wS#.Ó�z�b3��o;i/!=�aӳ��djK�#㌙��5^R��Η�T� �|]�Ǜ�T%����F}�1n0W�d������,`<''e81c4����x�ёq\�|gnя���{k`v�w���E�qb�>�21�zngEH<
���c4�A�*�* �h�F_#��`��}�m귛�x֌�ѨfR��W]5��^#�)�;걄�٫x�UZ�Zv����(sGT���uM�����(�	?E���9�h/M�+Uv\�rs��M�2�}��L��h��tS��`�j��$[R� *���9��aW��k�޾Wt��q~���S��y�a˚Κs�B�'ݲ��t���d�V���^���V�0w����1�ۏ� Okg��n�i�W�#��mQ�6%V�@F,���E,2�rU��/l�b����g5��C�'�~��h�r��x�ٖ�А�.U�*Tp$3�ѥ:2�!�.�U�큭�ٲ�4iFa���
���¼�����@r�{]
�*Zz+���~�nd
�:�yWܯTؼE����ц����:vu4m{����)��8w�|��a��1�w���M9����"*�<�'��vw��Ӈb<ѷ�j�ݫ8�}�o
�8.��{g�$**��f;<�P�"9��m��J�sJɌ�܊�|�B���Ww��]�0vo��P��I��U5�9�`�H`��
���9Z��l���DI�R1g5�{.���u-�Qr�����7wSk=t�SMyLOH�30��<;똾������mzo8�&��_C�ˉ�N�ٲ>��ԺH|#����Sc����aL��p�Y�@v��f�g�Fu��~���k�����l�X3��5���]���:��K��Ղ��[�&�)�iͺ$��\���7�^��اU;9���,"�,욖TٽU��
�~�r��yZ��;ܶ��C�;����m�|M�8L:�6�~-;8�M0��𜚖GK�3sF�EUomE�&"��ܸ��͝3�}R��Ep���8���}.��1�zb��ң ��;���:-�+k;r'b���ܶ?A����J��~މ�N6�[�Ϋ����`n߇K=Ϟ0��X�0�L�l�t1�ۛf����p��Z�p��ڭ��̬��~&1�Ǧ�[RE�����5Nz]r��X�����ʚnd���~5���w3�]��'�[J�C�OU�>�-��ر���_bO����u}���f����hD��l�T��*Bg(SdG9�R��LT�[^V:N�u�L5؊�� �^�'4q#|쒓���Ѥ�N��=觨˦��x�w��J���	�39@wq�N�l��,pԬR���eNU�tZnG02��Ko��w�g��5���=�P�,e�����7����;�p�@��2F��/�I�:��8;�FB�h?����|t��W])�w�{2� &g��t �^l]V�&�Q�꫙sp�ބ.G.���Rݎ��.g�Ǆ)��
� �����4 OFL���Sk�ʣ1��7���Ԭ�=�ޤFq��׻4e2��Ϲ1¼��ܧ�����m�τ�l���o�v�f��Ўq��6��#%ϙFu�Svu4h��M4ˢc�,��ʪ��SV\������f�~w.�ÿ�B+��U�r���Ƌڌ����5�
���~��iP�S�yr�Uyr�j����@����k��ןK��<2�v�]�/p�~qؐ�F<�S
��'M�.��t\Slͩ��30�X�,�g�`q#�-���[N�@P��!�ka;R�=���t(˾�x�}�z|zm�E1���m�b�!�-�Һq�!`�-����elm�5#������ɣ���q�z��zþo\����ο@����0�噐u��S�bz�V�{�{&i�׉����z_�*�+�m�SN�=yV���"7T0)�tM�q5��x�dE\з�Ζz����R�c{�E ��o��rKE�yn���Kz��\�,�c�[Q�,�^fh9+�$�ں���:i���UȽ�c�`�>y
������h�i&Ƌ*O����X`"|]�#8M�O6��ү)��(ҡ�o)ܜ���/!n.�:�����ʬqd�oE�D�A��O�˯.^�	��W^瓶eM���'i�`bs�8fKuzngzB�{%;�_l��>���ú��mg8��W�X�4��aI�k G'�޹���N��ێ��L �*���L�?^����xf'��r�n=�2�r���&�8Х�GGT�e���zlJvA{��+���]@a��C��x5����wכ$��3�f4C��R����v�S�R�Z'��p��2�OSK���j�7����ox�u�p���i�� ��{ p�n�M�l���ra�@D~'�Fvn��:��.���LA� 'Kji�)uc�rx�6�d!�ݒ^0.����ܘB{SѮx�7#'��t��5���wt�]h��c,d��p�ºC���y�э\���K=.�9o�.IC������8��!�C=>����^��eLg��}����x���(n�Svw���|�z[�}�9r�}3�qL��Ǫc�;��u��1lsͳ8�%���c�%���D��v�[���+A$R�O�5v��s�#�yb�`C_��t0�Wu���0��"��*[���{��^����x!�����x����G���q\���q,R��bS��{�1�&ӖB���M8��"T
�f%o{ �c˼���z��g!�Va"v��\H�H��_�N;ϗM�3="���:7�}�Q�%�bb����{qU����*�NTuX�P%��T�'��n��}�B[t={=s�+�ff��<K�(˙h�2���oFi���~f��k�	�qM�=y���{*�;�w�̅4��l�y�����D�0�#r�vY���y����!`[m��[�5)���֋���"����b���|u�����^E�j;��Hv�c�N��~�pC�C-���R���������i�w�/�A���'���v��d$r:�3��V�z��V�q�)����tSH<
���,�vY�5�w9�1#9��������3�.��$���g��]�5>@^����Mc8�ҡ��Eu�1Jk2*���t��.��WL%�	�!���U.��<����p5{9mIԣ %c���!]�󶻻NeE�����}�t�|�"]�*gs��4k4��г��o��)��-�"PP��]+�N�<?73z�Vq�Ek�t��m�*�a˚�t��BW	���nz������0��(�������'�s�+뮺ɑK��8���#�n�oy�\�mG[]\�F3B�Q�y��Q.�l�fYb�RN$�9:�>���L��n�9�����e���}*/yדd���B����v�(]�7�;���UW�tl�1;ܷ.p3�+if���l�n�d:�j,wtl �����n��	
i��(]DU�U�2��[-��An;6\�<�r��Vɑ|_�O�ϱ�,��TS@.��e���$+� ��٪���J��i��2��z��N���"�w�@�igT>WT�
ߣ8,p� ���g�z+�
��n�g�j�;u�okd�M}7��j6u�e��;�����i���K�)��(�ÿ*xw0�`��l*S�ov��A��3:�O3��o$?O��.]28.���������Zq�LOH�30��:�aM;"�sUYG_���͘y��q4��-�!��6�ꇯ2]$�����Sc���`Kn����UWd��l��dq��E�Lk�;9"�w��K,�r����eO8�owW;��I`��6���v��5�:��5�?6��0�K�ѱO�;9��!`����KdԲ�f�V������iڮ!���_0#��j2�6�T�S{z_V��E��M�_��g)�a`)��uxF����dk�eU���XD�k�wD�}��x[gL��߾�����M��8��h�]�Y�1�zb��&�R��^���7v�M��:i� }-M������T�b��K�Ƶ�#\��q���6�O��[�ol���f��/w!�1Gb�r�j�]�R��ۊ>�4oD���%:���9�t�q�f�;i3j,/pu'�'&�x£6�58T�)�b�:(�ێ�'�c�^�1z�+-���ཽ��ޫr���ʛˣ`n��g��MmZ��v�"n��t���b_�Dক	��N�֧\<�7�[=��Y�l��o��x�zl�$/W;�9�eF�7��􁋘)l�^��Ss$SOC���w2إ��RxEʞC�3OU�>�"pV�[/Nvz�� Iݗ���[�.n��
hD��eR#��i	��Y�qC���U�lke*kq8w^�W��w"�|
�_����W])�w�{2ʽ1�Dt%�
�a��<�q����9���&.���a��{�7m����͢�W�]���~J�x�p�19��{}�{)߰�sz�:�c]|����z��00n�MK��7[�Lp���S.��aTUG�֘�Ml�Xw�H�p�m�S��(�{Q�E��N�]�M)��SM2��f\�0۳�r��u�ۼ:83��<;��̗yf
;DS�9-WA�ϵq���'xvp�|���h�����]EoC��Ol���m�	ȁ�0��ahɷ�\&�ᔓ��).��Rht��w^�
�B^�����5�����i����w(pC:�[��;!2V���I������f�>
傯*;��{�kw!���'���+�S�ˢ�pg.���Y�d=��&�1�S�Vj��Zo�!0��>K�)g/�/�f54��.c&��g�Q?c���8�-�u�)����Q��F����<��.F6�[9���l�jP�6�k��ttE��А+˺]��	�}�G~V?3K��Ea�������x�(R�Ӎ�p��MOn����U��4�
�wG3�=0���/��}�r I��l�:�'�-��i�;s�Vnɾ��Ӱtm��|ȉt���m��a�~������M:U�>{{d@���I�~�x:	�-�j���0<��n���+�ю3!?>�'e=z����oE��K���-����n(�\�q��ݪ�GK�=;u�3�{�e�s8+�� k%;�z�g����'�-ָׅ��Ƀ}���%)�Pϻ�z.��=fe{�#ϗ�A�^�xޛ�S?M�3��.�N���j�Wv7/M��A�F���Rٖ�m��ħd�p|=���/�	�Ɩx߸��3��ӗ5�*r*K�:d�m��T��n*�!��\uKv
p��`���ÅL"�ˈ!?l뱼�e_��g.�~���.�?Φ�8��y-�#�׻�7m�S�2�}Ʉ+̺�yk�sF,j�a,��N�맻���K�=��I�^���1�̼���_t�/���AJˮ~�2"��T=j��Wx��f3���lt��T3t��5Rg;��a��Pf��c�p�̩�k0���㯺p��N6B���ȵ���ն�5�q84*�SS�<�7��_���}������zڦ��	t��<rm�!��c|����6�ix*��"�(b����c���3��=�,�y	 ��2�'o^��J#qt��:�������t��m��-�2C�uU�ޙ��Yܨ���@Y,���S��E5��*3�HhT+�9�"w2wÁn�C�l���}�n��L�fs���l�LA[���Db�|-����&7�Mۦ������	�ye�|%�Dt�c30��<K캍�.5�K�d6��[{�jӷ�P$WN	њ;6�����Į�ÀL��	li]/a�X��H������ZQ�k�"'66���:�t�r'+�*	�ds��:m���MT=zʗ��w޶B�pW��%�1c\��˞�p�� si��[l�T��
��;m�S�ϲjS��85������~���ܩ2Ř�&LzQ7lsii����i�Zy���L����ʦ�T��`��xKd짯A��zZ�36÷!B����T���y�̺d�m�*���7"��K�����r#�#W��tSH<tϬ�/�;q�z������%��]9��W��1'���dH�y�|�j�;N���ɍ�epV��xUpՉoH�Kgک����7�м�f�JV��e98�;�O|�
��:�7-3�!ͥ􏛎��*����8����6���h��y�"�0�O���3�?��5\�g����'z����>x��h��B�{�>AuM1r1�^Ɨ��q��~�vK�<(�!��gi��5V�g�c*��uO>�7uY�jH�.E�N>jq�Q���d�gj��_�D��~��.�{3�y�#��lҧ�B��~��L�mI�ƹ�����oO%�Cn���@��H��z��q��w*�&��駓�J�7��O��?�
R:w��vE���tgB�$����f~Ʉ "���2ʙ�By��	 ��J��lc91���͆�'Ჷ2�v��>�)F�tvW?[�dK$;���=�`��B�~���_:�%���5�{H�:9��Db00���n����c�
e�B������0g~T���޹ykӚ�{`��#�q�b�Q�D����1����Φ������fa
c������^����Jr��1�j$�3�b�'H��s7�K�\���C���3��j�c���ß�*�S�݃8�'�$on��D�P@pGu��n'W�{5��T��bT�
��'}�2���3y���{���1���������1����������pcco����6��61���lcm�������1�������m�`��6�lcm�`��6��61�� cco���lcm����?�c�`�nlcm�����d�Mf��wh zf�A@��̟\��yD�B$J�(�Q(��I��T ��Q"
I>�
 �UET�J��E)*�	UB�H���4-dZ��i�UH��v7l���W�	JP�SMU[Y��5�U H��٦�HJ�eOX�$��֨ j�
�Q��x�J(�B-z���*%*�Z�HAZԕJ�(Ai��m��L�����	UD�J�Fƛe���kT��i����DJ.�U��K�   ۛ���t[��E{�y�{-�+�����if��ws�3��mY�z<��V����z�Zֵ���(���oTu�ev�X+֩-aKa��K1JW� ��|Џl�̡�:Yen.����(��z��(�� �7QF�QEtn(�F�(��9���(��(��(��ۼQEQEQ����E R��#qE7b�$+����:r�I"�l�� n�R�6�Xl��oX]b�ӵ�uXsn�����1v�m������-��ë<��=�ʦҺk��Ύ[���Wv��7@I�v�l�zaT*��M%��K�  ��龷UE�N��z��kӫ�{<�4�2�W�������]޶�)���^�kt����ӎj�K���\+Bݦ�+���ۭ�����=��']���-�����J���v�q|  �ھ���Q�����ҝU�n��RڻK۽���[gu���Wn�6�u��wv�^�����]J9�{�^��i��)����v�Won�{la�X��ΥD��7��'cU�U�  7\�wj��g4w^޵�w-r�S�z�F��M��3�m�v��Mn�v�v�wHgwmf�][���nݶsW�t{�sm�3wM��p�k`w��{m����t�elP�.�Z����I|   7_>E}\�eV��sJN�sw�н3��S�۶��ݮw����.���ǽ��6�oM�Q�V���f�G��A��jU�z�Ƕ�֡R����[�n�T���T�T͒����X��  ���*�n�J�of�W���l;N�v�܎4���������z��nåSM�ӽ�J�k��]��j�=ec��ݺ�w3��^��{��'U��Z��R�ѽ�����M`��  �;���GZ)9[#�s��u˝g4tt]�H�å�������50��Mgu���RDTvsK(�5��vدUwv���۴�ӳn:����f�"E���+_   g��֯���nn[��KN����=�9Sh��s��Pj�qݙ�wN^��6�m[W���Q�z=q��kZ7{���m�[�5���'�RR�@ �{FR��P �)���U2`  "��	R�  �~A=5US@22 B�	��$D~��]~���߫�RO�ѯ��,LP���:���yߟ����Z��}�؊�+�����TA^���* ������ED�D�����?���Y����_�ܑ:9�M���n�=���Y�E�t��Q%X�D�ibJ���,`�V ��V�v�����w�oQ!-f�J�]�����h�GB#m&���c�,�x��9q�9z㧨���	R�aM�Q�w��������Jj:�n�J�hk�j���-̺Z�x&i��A�:��*7X ����oSi�Y�~�c�0������q��fYa e�:�J'���/U�ҋ -j^�� $�Gi։x�C1�2g�ͼmD�Si��cn�]�ҕ)���Mim;y��k�rX�Z����h5���H6B�쀕�HZ�쑶*M�"����\yio�kw��!)�b�D*�S�֗(�Ѭ8��sY�q�xac��F7���%�a�Ve�s�M�̷V1��7�	FƐ����j��WQ&,ord�,QP�nmi��X�Id�n�	�DsA��PX�vⵋIBϲc��d*p-��)�2���K^�5�f�����:V��i�5v�k��զu]��KV��G�I�E�%��̖J�t@����P:��7>���aZ
m#b����zN �BJ{`����U7`�F��Y��jda}
����c���j�
Z�K�4R��˂�-�,6h��]̴Qy1E��Sʰ��$�[p��<�r�~Ke�CLjA�-T; j�s`�n����1"����Z�`�h�����LmZ������K �*�aDR�N�Y���!��"��T3u<	�Z�f@��S[���L�0!	7:Y�(�t���Wo-Jf5b�%�)�pJGI�P���Y@�b�]7�7+a�#k�nѠ������(mc�4x6)���Wz��)\�$!��:Zw�QFK�;)��K���n]��-�]-K��r���S���+/P��n�(� k1�^����E;���U��ъ�v2�\���0��v�j+Yt��H��uʔں1�2�(�aX6�ݫ2�
��"%�M�R��V�kn�3�|�w$���l(yue6"�V;�~�����r�^U��s
i��Z�FAd퍏YӍBË(��d���.�;i���,� 2�F���4�s#���X0A���	��kw21��jЎjYj-��rȇ26<#Xv�U����2�ckS��[����~��HH����&���.��i|�)-�@1�XpJl�4��*��U{��Pb��U�Ra�&6�QАSk*����W&�
vvG-ZWN�,-1P֢9C- f��B�֘[Gv�5���bh�XR�J��E�cJ��+��cѬ�8���Se)n
U)��fYAB7xL1�&���*L�B�W�*�e$�lzT�tmn*�c�W��AG��͛T��r��G��Ij�j^���ݳB$F������Y���:����VH��>���ϖ��Xk��n�,f�ս�âVإ�9X��o+D��<�i��1�F�A�ib6�n;�m�l�Ѐ�ꡐi]�+v�/m�9x���(VJm�ȕ�p��5D���96A���m��{X�xq�V	N��)1��p`�X��H1{F�S�6��$�.����1����R3�!iWF������sv�������X��X����1!&�3[�3EGfc�N�:��l*
���-Ț���{[����ʕ�{!7Y{HHYU���wu�@��v��m�������ճa��Vj��X�ee�jBñ�6�D�d�q�d��x*V�ՅƖ�
 4Aǡ]�v���J�O,
N�0^M�+.fB*֣t�y��%��:U��[X^Ԕfꕑ�&,L
�l��j���zpV��+/��i�"WI渜9w�ۺ��r6�%����Qm%�ز�2YE��өxd���� �X�"�u�-�b
����H�b�l��9�lK-�T��I:�u����6�Շ�j�N^��)��,��r��{��]��u��n'r+�u'	�P�L����@�U��Q�Eu�Y�:����̱�Ձ���fJ:3Q�f՛ԅ�GPKF�j���-�QS�	KE�����^\;�	�6� 4���`Mu.�� �`��Ovaac��[d̓b�Oiۦ>��0�֍��h�`:*`��)P9��t��h�kgQ�쒚�>'^b{��j�['��	��V�B���@�I6��@��d��t�Pֵ���V���=R�>���ʱ1ͬ�9�<�ڷef�4�L�^*BF�JCVd�"�b�r�]݃RH�ݡeb:]
1�&�p�x�v��J���s��1\�7����2�B����R,�j.���"��ĭ^h���9SA+i��]�Q�^�%*`��֟���@H	�JեF�HJ[N�KMųF�h(;����T�z�ݙQ51S۽�&TՎ�x�;I*�k5��{�L����Xw�)�j�!����Z�(*�-	@JaX�������.�*�ˌ����ʽ�%�,I)�A��Ȯ�����[N��1g�~F@�w���,�e��PHț��T�*�a��ڛ/o/��)
��>
������v�^�Rj�HY��n�&0� k#% �6�i�6�*�e�V�#E�%Kt�`Z ���*��܍&K{��֭���4�2��t��f��>Fh�.Z� B�P_m��!�we'CD*C�Ǹ٣Co+h]��T�һ�E�� %ޛ7fV\GuS�S�n�$U��fV�d��G�M��
����C�4�R���GdZT�6��j�� ���e�4�/*1���zZɹT�:V�X�\pܠF=�uQ���wL�2�#K�P�H:�$(l��dc��u
ڑ�5�#K:��f��Qв�X�2��tS2��c8�ژ�2$��l����A�C��+\5z4յ���ƁqV@����+*[u�(���Cj��Ԗ�8d�Q\*��^0%
�X�K�)���3!7��P�.�S:Kn��[�-���n2v�}k@hJ�V���Q�[q�{��*L�2]�N9��Q�&�n�*�x^8jM����p�8�YyYl�SZ��,�^sr)p���f�H��p��v����;WT#˵��<�#6��f�ö���(h`sB��>����5�M*�Ĵ$P'���� ��J�j���.-��鳥�cT�![�Te�ŕ�7Qn�	��]KBY��:�
�z�n�N�����äF�Z��S�hV\,��pU�\֩�tm�F��R�P[�Rz�F�D$�I��k̶M�lhM��ܷ�҅�ʶz��Ȳ5Gf��9&.�4��˚�MVǵd�"Mөmռ�ɹ$���#��/q����~���ywq���֍5B�e��l�7��P꫔�)ʳ�#,�V�ouR��%�Z�wy���3Y+YӺn9w���Z0�TXD,��,�ڦ�k�/k֦�& �E��j:7^3uvr�S�(!5�Kd�Z��T�i��x�9l��ue�&��,ͬr�V��
s//�44�7VV���O f62 �%<Km���	fJn�^�&�`���̵ X3���S%�9X�]֜��؞V��N���1�+˺q���F 6K�	|��fR�!l��Ĉ�mkJYX�Y���:��O0�12f���U`Ex",�B5&� zK_m�h��!O'�k'E���yB�ܳ~��4Q�{��/+w��Knj��X&YE�EI1�s��p����9��+�jgyY
�Ƚ�d�����IO���H��b�ܫƒn�ت^*�'#/dy�[t2��m����Q�F����B�컍[(��Z�.�Y�m���fK�y�
�̈́F��T�W��x����_�R�`2:�4ӽt��yMj0<�u�J�:�md�R�	�2�8�`Y��/#���rm-�V(�*S&;����N@nˁ\ ����h�u63e��"�)C����8�e7���A$�431j�V�ӺN��nKt�̱ob�z�a������_iXU�R(�d�PZX�o.!i[��Զdڽ��L��əWm��w@�L��ڽ�$���p�/hĆ	n�fM��t�p��3���YƱ��'v�����7�K�`ҙ�'�2�(d(EЙ X��
�l�5�EZ���t�5VXH8C���0�n��`s&�0�
iJMʙE=Bdoo����J�Y�T,�pYn�<��f**�,@����)l`KuR��\@ ʼ��bRڽeAF�	���[s�x��T�qL�>:(9x�kBb���H�!	��bU�u�hŚj`I�]2�D�&��d�6�Mj�c��)ԡ�s���R�F٠\��cm���,]*M!{�nnK8�F� 
�+�=V�
��5�5��Yb�FmCv+N8��*�hSe�Գt�1�M�v�L@����.����$�"ĵl�Б*���؅X�"�,�oK�Z�HF@tq;��U���iNwv`gFn�1��ؐ�EU�^ꑆ.`y�B�b���N�0�et�囂�A��oi��W���懱�oV���Ԣ�8ȘR�R���L� �1��\�Z��Q;��8�k�F�F����;-�9��F[[P����܎����1=T�;����1��X�6�j.�%کF��Yd�[GQ�Y"½�hZ�V�O-`��1769�J��v�aI@�	E���Y��V0�bҔ�'��&`2'�` 8J3r��`�h��M���?X�$`TN��r�Ѭ��:�z�nwT�wuu1�+��&[X�`��L�-DÐY�e���CNl��un!󚠫+��#X�ƫ�Ph�	���z2�b��Ø��m���lV�h:q?�Z�B����b�'�RWa8!�����or�wq������T���,��f����ұ
��BX%]$wib�{U�4�,2��Y�u�����B�r�O_�R�śX��)�����d��J:9Na+
�)(v���ܔ��Ws�GD{�m��^G{SuM�i�LM��oMZ��(��l�-��
��X��SV�5�Ce������Ne:����J*f^j���B��������YM'�8.�^��z�����eL�n���̢�T3Ba�i��baE��[�*]�U�h��0�h,Ȇ�O��a��2,6�e���Y�Z��`��;� �7#&
��g��wP����m�kC�#] �5�@Y�h�si��ʶ�TE��s70@�1V���& �5݄�*�І����E�@e*�n�m�udf�Xij,��v�v�m�݂�{��5�Yw���Ȭ�h�"��^SXp'ۣ��rj�ʰ�;�y*��*�W��-!Q�>Yu���5#x[����*P[K_9��p_\Q��]AcfF��*$��NUȮ���L�}(0�h��wD�����jM[����ek�E�Q�N[&=���J�CZY`Ԣ�1���%
�#p�$?i���;'��$�&
�)�mҷI+Xح��f�ީ���M��'-e,S���͎T�H��ԁ*��*ִ1XR%����V�H|��R����x�%�ޠPH:al�v[� ��ѥ-�*-��קl�
��̼��H�YPV뭒��4m&l�;w��"�i��vGͱ����,��d�v�%�)=ǔ�n�h:�u�n�@^ "��Mm�����%�,�f��h��ٔ��!f٢�� J9�B;נbw��A�V����EZXw���Ij���BM��vk�H�m�r�%*kHJ�èY�xlPHbA��nQ��մ�3{��ݱH�A�9$�'�F�sZ�c�z�VLw�(���0Q4�&�Vb�f����ye-V�!���`m�/]��YLQV�4��.�Ւ�)(+u�"Ev�m�
��P���c��r��k-v�e�Uv��S�H�SRg>�i�V�
l׺VS-4�����!j+v�e�Fn��L�e�F�N(m�;Nj��wέ�nK�a��R�N�����H�+tak-��`�^3�a)�G6�8��X-�$�r�a�q��I8��j��.<Ջ-P�=�7Q�0�U��D���T&,oT�kcu�5^�5�
�N[�r0�K�Rڴ���jR����❋�ɱLn-[NK�w�e�t�߷DW�XA�2��WolRM����ٶ��M��K6n�Kc�ꍵaS�)$��h�g]�$4�^a�#�r
v4��^�Xn���*z�]0 �MK�����C�ܚ��j!��(=e��n�н0)��*��<0�қC0��d���K�,�� k$옭C)1/j�$Ò�S� �d�u�X�ܚ\��ٸ�`�o>�l룮���XW�f�eCYl��*��+��~�Y����Y�D� ������>b�4��6�3]MF�ĕ��<����O%E;v�)�NnJlh�d\�ca$+�b��G5�M�����OMe�:���l��4�z���� ̚m�b�H���6��h�~؊��l� ]Ը/�����]ejYuӝ�h=� Jo]�4eY�Rʵl����z^F6�}��r���dJM��7�Y�F3��l��i�C������R��"UɖU9/S�����n�$���[�qP��4)��C$�F�tQ��zq��x�'�e��Pך�5�ԃtM�YY��r�K�2�0�Y���L����%���M#���u��+w(�`Rx��EV��hU�8@�jQH��W�3.��������ˡ�hj�&+�f40���dQ6����xS:B�͒hb�F`J�AZǿ���4���՝����ж͘+
��S5����辵]Le�
�,c��NC0��m/�S�ٝ�I�]k����R
�'<�����&���6\��|��5ٵԉ[�Ck)�W(��,K�\�F���]���2���w�"S.�M���|�J�:�.�I#�b�}\�h�s����q�@�]�SE���99W���m}��=��ۂYJ��s��HK�ίK��z���g�H����u�3<TU�u�'�.j�ɯ_d�]-*���8��awp��:�;e�om��jY�q���!��\�S�����e�O4���g��<�I��&�
���2�KXj�}Al�9��Y�v�t�D_nN�y;�J����3V���]K��V�ڏ3��
;=+eɰ=H�u��$TJ�1z:��ы�oZӉh��� �啪�ӏJ���v�q�O�,�P�齞����	Xݨ(c�����ʝ=�@��V8v�k���Ψ:M�Z�3t�\�8U;u���T���ur��}�[�QYN����ճ��nMwQ�6�=�wKY��|�q�c�&5�՛�5^��qݐ�e���l�Umv�1Q-���k�[��)t�Z�$^p�g:�]{���u��ڒ{`^P�q�E$�_=����Y��6&��=�v��W�64Vby3���j֗��'.Y}����|�G��C]=�cF'R�T&�[h���+B��-V9��w�1��e��A�W��ND;�Wu�C�m�I�T�.�WNgXf�M��+J��nf�эL�%�4i�R��(U��IEZ�<��{q�]}�[��M>
���2b�C�΍S`4r�36Q�鶡��3�p
�yŧQgt�7��R����ԫ����[^+�4k0�Ԇ���,�Qv쏝�x�buM-w�1-����v���:��2��E L��1=6s� "��g��g^P��8���_?���*G�Yx����dA�F���z�p��8���B�3A�:vA�ԝSA)q���1�K�KT��D �5��Vs�Q7kj鼉�k,��@�»:V,VJw�@�۵�-�����Xsw�y��A���m�]�^���}�.�1;�:f����O
Ib�%A�%��-Q_!V��ɺ��
&�WW*��_<�����2������65�l�i6�vM�z�)z��}��W�2�|����lG�ڧ}�-�]���#�Z��VLNtpٔ;�ٝ��c��B��V&�N-��{A��`X���=/�V1�}Q��	���A�y�q���_(PɃl2��3Nu�W�6�rիP�r�U�޽����������(����n&�������[R���F捂�r�5�"�5���d�M�
���Y)��ui>1���U�[֮���g��<�wW���O��A$S̗�MW�����w��b"�	�+��珷 ����� �yG7F�����:����r}5T��G'w��	�)��j�NV�`�Tk��Q�
a���!��	� ��@�9�=-{��`<�N��;m^cn�����lo����9�`��4�l�J����ֻ����E;��ުY\�6���u�.�ܓ���m]�"�+x��7h�N&ڴ3�{0����v�F�V-��.��T�$�:�<w^�BIC:��5�}�x��	�u������ur΂n:ͷ����d%n��D�ehn��	��Z��X�^�j=�C���&�p�.�j>�-P��m{Hz� B�����v���@\���jM���ˤy�����X}�t:�����w}�vDZ���]f	��MX���ح�GX"&;�`Y��>�	Ѿ��	��z,���B��hJ��\u�T�Ouj�O _+s��X3]�b���l:���ZA�xf��te���R��Q���u����K\�$s�9�s��rx�PW��ؔj=ԁf�A�+�R�f�l�ޜ��I^��&vή7����+�L���n�29���y�s��!x��`0Ԙ �dE��{v*7�9�����72%��sn�UH�gh��pLW��t�w:1��Y�x�:�介'p������=��]�$8ȭ��=8�;v��?*�=&C.�_N'b��ê봢��Q�H�V/�M�1���w�Y���iy�=�eb�mB�\��2fëq��X��֟=gj�\��:V�˃Ӫ��]����F-�xp��AE��:4l+;%�Kp��������K-T��C�)]��xGt�J7S���6��s��	 B[K��#���	b{��1o.j7\�Y�$2��S�'�'��6���E�r��D�ѳ��҆�X�,�K8m�z7��(U������+x�Or�	�5R啝���9��2����8lh�Oj�d��`�����K�4u](�ѯr���<wc�p�멽�
���1����cĦ#�#�1�=��Lu��F�k0�Љ��ʝ�	Cm@�CGuɱ�޴Gm�;)�5���]�ݺƀ����'h�	]K�=ԁ�ۜA3�d�Mܵ�ݴ���&����_6�+��<�ڻ�';�� ;5:za���
5�\s����BS�sv�7S;{^�sS`+\��<7hZ���03W'�v�н8.����$��~c}ЛH�+�s��ϫ,`oVP����[/���Ke.�i��[k�\��k���6�^����9yE�H�rF-���m��;0>Gkt�t�_ݫ���e�8i�A�H��ή���鑻jWIS4�����l|Z�\��[���7h���[;�rbi�hw.-�d4���7N��S�J��3`��h�
d:d�i�n�>d��۾=����P�o'40�@G�(�[�@��O�T�9���*V�\�ui�����6WQ�S>ҵ�=�-U<HU�on��6�>7yj�����1�Ul��V3i�<Y%��f�HL���vi7"ɵ�wi-�s�����
���J	^55�]aE������(Z�ΈV�S�[�5���۰�C���.8��)[����\��g ��	�j���p]�n:�h�Zs:oy�g�VT�l�[�J�h��[��J��l���F�s��Q5�~�K}�'u�z��,[��eb@M�0�����ŻQ���4��$��ܮz�E���a�����w: �M�s�F�;,�q�zNRXm{�1\xզ;:�d�$R7w�����K��r�A��H�ȣ�F�%y��y|zaz���K���9���;�Se=����tk����i��}�g;4�α���S�RU�jU�L��Z\@	R�K�ܵ�ݏoIS�ކ�:�0m۔�G?�ޑJ�y���עo�^�#���o$��C�m�N�2uݳ�C�ed�9&%|۰�Rw{�̝�ۄSu�ɭ�����ٝ;@�٧,�_m)�#�U�E]�c�wJ������Ou�Z�y�V�؇�)��6��������GE Y�2qm����TM���!�ufsM�*F����۾�� e"�*��ڲ��I���*c��s���
����Em���we>�i�>p���W!��c���kru��;�[ONv�����P��>έ2��e$j�
ˬm:
�(V����֓7x������� �؀˙��o�c��*��Χ�!E]�b"�n�Z�z�$��@�/z��vՌ[n�c7c���h�����k{.;������ʊ̥���Y9��aͮ�֞�����zkb��+:�}Ls��n�0w���°���]�1��u�{�7'H��r�qwGE�Y{ה��Vu&�U��-��!�w���O;k^�^p$�`JጛNJu-��iSt:�4�T�Q�Vm�\�7D�CP�>�i^�d܇"�-�fU����D���`���6d�v�Z;:��]r��q�yl�l굎ob��k��ȃ���ⶁ��YÔ��!�E�Șu2��)�<��'��v^�j�Ή�r�C���[9\��u|���1��cb�r���[WR��A�Z�j�W�gs;��oh���t�`��D�)�Ԇ,)\�a���C�j�1���t�x�v�Ӯ����&�(�\-�v����ݶ̧.��0@,F�W{�4�����wQ(�^�!n�4�gٔ����@������ٔ%ܖz���]y(��S�	�qԾ�tXT��3���w9�]��ߐ	W.l8�\��a����A����TM s��e�n�S��.ۤ�Rѝ��6�%<}ګ��`Y��vB{/��C(\���Q���"�[z��Ou��c�Г��n���FX�X��{+J�2[��:J��@������������R���Z�:M��Z�c0����o-�MR+#�	�b=��|^���3I$�K�T×i.��v%5.i،=����\颥��>k*�G%K(�R��0�Ӯ���
�F��C������t���+j��Y0]���Z���d�t�IK�o�+T�}�[��u�C�uBQgk.vI���k=�l`4�7oxE���������%��;����U�FaJ��c�<Iʩո{$G��WaA�K�u�����8�N��:�ã֑��C��"B��|�s�Ѭ���_�T�̷�Z�U����̙�.VX.Uᕍ=+dG��v�y�'��+��Oun�1�+U�g$W{.ud�"1(�i��y8^\�+���J�C�H���f�A�����/9}���*�����.��y�˰>"�`��qt�D�y�h��9"�;f�8/$r�v���u�����8��:.�[�����2�Ԩ��/l]<�Γx6�o1�=%�ޛWr�Ok����:���Rv٭��q�Q���[,\��éٗG��2��S-�\l�u�������c�\��oyʙc+�7}��HW�yf��Ǯ*ۊ�aj�b�ӧ|C����ٝz+�J�9��-��qv襝�W�e4Z������;��Q�[!�ׇΏ��黖��X��˜�U�cvK��R�om�k[n
#����	J���1fu\�(wh}�z�R�TY��c��SnI�f�|��j���	�8f:�u�S�$�2������*��6ɇ3gM��J�:c�	=J��?�↼�r�ĵ�M��J�"x��:{������;��۾T�뮺�8�Υ�S+]q�3ܽ�)��^�*�-�%�-�wv�LGI�O#�\��L�4v��;/ANd��������O�#�W�Y�z���·��L���к|W�t*��j�����:[��:����b�.�x�v����k�K1�2�}eY��\�h��6^���|쥐3��G<�Ɗ%�wGy���e��.83v=��]Fh\��u�k�ӊn��7Ar�\��z�����y��4]�}���8�Lj�M���n�:m+b�6�y���
tN<1����mĪC=v�[�{n��C|	洆�a�f�t�)��#���yf��Z���h���i��f����ɔ�a����z˾=�)*i������뭳z�2���.R���M��)Z�"[������w����Y��C �G)��|S����ò��N��m5z^^^n��iY��iU��ѱi-�{��Y9��Z=ؖA���5��r<]ε�����v��pu�����VQW;C7X�Z�Cճw
{C��J".oR�1<��(�ӭ)*k<\��g���o�1�yyU�F��"�$�3���h���7�o�T�-�%vf55��/��v��"Z�����������=��Kp4#a<䃗]F6E0%k
o)/o7��^�}������
嶞�oi*���u�s�H�p�z����WsL�Jry㣭�μ}G{^6,�}����]�V��D��U�FU>�ٚ*�s`/�
Mg�z%J=X�hS��b�2\GF7emgA.[.��X��M�+8����j6�!���Q��κr!�;Uk����l݄](g`�8<���3�I����H�)�K��GBt���o��M\���2M{��m��1�#i��&�XWc�-̦	�v�\V8�;�7RCb�Tl�����X�)��D�,cf(c�5�O�)�^��^�y^,���($�)R�#�H�I2��eNO)�ڵ�g{�`*�͸%��]J��Z��ɯ3����{l"3dQ+��._�e���J͢8��yˮG˙l�
{��WD�a)����p���oi�}+��;e��id�l�����1�m^^[�0��a$�WY���a�ܔ�Ho�� �읮�QӼ��.�����X�͝:��W񮡀뷳n�S��*?\�GpЃ6]1e_Y�q�,_^�SyfD�n@��HCz�%��D���YG�e^6�;�.�qdЙX�C�֩p��nfYH�8Yqo%�5]+�P�+Ӆu��Z6���D��3q�f��:�	9�'���iީ����%�Bh��Y$K_524�93�`<�:�퉉��U�h>�O�����U����o7�ۼ-�P��Y���-]NF�\";�-���z5]�.8ۮ�Ѳ%��e���_q�B/-[�E�Q{�����R�ٽ�S��{L�k�T��-^-B��IJk��c���X����Ue�
ǘCh𼜞h���0c�Qh���-���(z|�;g�:o�14[���uqӦS�H��7y�y����/u���PV��I��vk�J`���Q㝥�Ei��Y`tWV�q��]��KIɮ��Kw8^�=Uru�w�aE��&��i�@�ZRs���Jt6�`��W�������Ryx�omL��s:5��H��ҙ�?fP7z�g:� ғ�]���i����[���o�/{��7���T@QO�EDz�}�c*eS��d�\uċ�/�g{���3
��W/���sxA`h�lM<\�5(h��m�x�JwI�K�ݜ��q�uܨG��7�1̫0�t;��ɐ�C�5�6}sD�{ڹ�y�EK��Q�]e��m|���e@o-x���_\ז3,��%g"�@��\��$��kz���m�^Cw�0�P�E��:ĩ����y;n�u`*M����u"����tu��uq�
>�{j��[��A>W���DYםm͸��R���R����Q7�n!t5�f��0�j��uε�����"��u��O�\В`�o<���`L� �9n�do+H��k,w�U���X{�t4���α��	7@�nN�$\+o���D>�������T16�U�rJ����󆺸"��v��1�)�Kn�>�_�ug�;�.=�cT8QWZ+���3]�33���U^e�5��}�h��W������]\$d�z�`��H�s��ƍmY(��`ŭ���>[�Y�w�H\�`��(��+��2�<g]�����e|@�>�[/uk��V[0=ܯA��J]1�o�;(Һ�
b��t�`�Ǥ��;�K���+�$������¡n���Zۭ�!������Jn�w�O	7QAjl�u�ir�nՅ�o��SoRٶi�
�Gor�9-�.� �β�[����N�j�Dy��ʄ����HS��r���Km5RL��CM��ٔ�ܱ]��,wf����nɃ�q]���sܽ\ym��!���4�7�û��k8�=|���p��]��ԁKn�哺ΪI�*�;��l
:Њ�s_&�Z�p=�3$۝j-KLj^t:�$�>w�$��|�]";U���l.��r�^�}}h�K9����8w3Fɱ�L������Y��_9��E�jt��e3r"�N�̤�[2㕺om��v ��nܛR&P��s�j���ה���z�:�KD
eb��^�/��HW�T�7n�6*��L&W��s)�;����.囚য^d�4���];zGQTCX�;�pC��m�Vk6V_J��^�!�5@g�A�t��R�H�v��C9<�
��t��ܚ��O��_$�q�?mt�*�,>��+���z+[죦�$c�ƌ��ͧ��WJTI�m�P͡#<�:���/6�7h�p�'�M�n*ed�/R������@t;+pF�Q���D���g}f�ἤ�U:�-]�?/
��m�j
e�c�p����ܻ�r6M��h�Se4]�r�7E�m8���)�X~�8��Є	��#�,Wl���ia��w�̹�2�C�T��e��v/L����^k�,�l2VҒ�:�0��R�O0M�Dt���H �q�3o���I���K�q�	d��u
j���v�%��[�a7l�3��:����d:��l�F�P���j��\U�Uݺ7b�>�uc�8�E�0��]f-��r�q�1�n�1ͭ0�8�(fq�5]��4{n�B�����j`5v��
`�Wf��6^�|
ɂ�;�ɣ��M��d���ڍ��*�ȥ�ԅ�Ia��`�� �Ԝ�3=ٮ��fo �5O+�7�[�&[��+�

��8��B�wۻ7�e�m*@#�j�^��j`��2�FH���.��H�,:]�Su�=��	�g奧Xj��C���MJ�&���36U)�-JJ��yb��������!�b�K�rۙeI�<��X㩖�^ފ��8���4���#펝����:�8`�l-����L@f �唃l��S�InS��=V�l�*`<:�Z��MN7��p�z���.R�$\���eJ7H�H�������
����І��]�,��w]�G|�S$��`��9�/M��C(�`x��Rt[�*y�]�z7��Y�W�*�۱E���1܎��b�u�BԠ�u\�Heŕ��`����N/�t�GrϢ�,c�a־W�f�ۭ��C����{�R��k�Z;P̨~����o�u-���<ņ�(i=ج^9��.������N��We�O-:��Ql�{ӑ�O3R��.�W]�g b�r�(�͢�t6�t�vWR:v��giƶ��1�	��ţ{)v�a ֮���De'@�7��|��f �[�c�U��x[�\���(��xlu�r��2]����5sł�K]OcM���{0���XFn`X�e�	���������=���h�s[ �:�{�M����n�^R.Mb�����ʭ��wN�N���Ӭ�I�j-|	�}b��TQO���7�΢4F�*���2�T!�b�݊���X��J���`�՚k���a��cQ�4���-�o2\V��Y˕���Yty�r�X�wm��n1��U �*O)��p[��W�R\J�2�T�d�O��Wp�6b��sr��T�9�y�+pБE�z���(7-�8gtÚ@
��ҺY�@�eL���6��PjC����L*͘N���̺�ݬ�R�r�Vj�ݳ��Y9u=�l�,=��U�H7�n9��׊]X��N	���&5Q��j�ڈ�w���U��ּ	�Z���.�����X���E�=��WwD�%v-�ۏnWmmf�2WVd��`d����
t]XX߷1r��T޺Mt:E�P�)�L�����6���%���N�x����b�����Rz�$%�l3��鸗[�=����ҖC�i�ݭ�V%wwM�\�6�fʼ�����Y�2�ĥ���C��qYJ���K��"[	�����)�[�yD�)J�� �}A���;	Ӧ@3�gs],����c��c�8݀���՘�RɎ�����Л�m��p����x(VV��9cj������ }|#鑪�z#ڱaCZ�n:4D��u�6�� yw�v��s������~~9�ﰯuv��)d��t�y��]wq�ɠ,�3aB��L%�����8�=$5��Ʊ��(F����:V�5P�v��mWc��\��S�����$�W����a[����0̬k�Q���aZWs��2Gl̥ñS�{eizVfmoq	�(�f��&(�����	:�T��J�ڮ������ήY�j�;cd���vL��\-]f����{j#$��;�-SJ��_Tu��߮�}W���Ƀf�*K,�s  �|0�8�|˼��Z��XU%���fu!�7��Q��
ep�W#��&��6��i����y�+tc�:�,��{i1����Y�2���XF�,�:Ցe���^�-���c �m�-'e}p[��35�G<��q�:�h���w�<VT����F���E���U�u���*�v-g�n��j�V�S�Y#z�c˦�Vi�H�IW�o\�ȭ���e�y��Nl6���Dw�z: R��M	��.�7�a��ګ��Ȫ�i� {sg�b�� æ_V9gX0i�+���ar�H���]"i��]��v��[�-����U�H��|ھd�r�#]�](�^��T#=�X;$�[ڳ�z_m*=]v��ߊ)(��f+�I�8��7�X�ɻ�.�4$B�9Nӧ�#�b5�>�n��E�t����7����K��c�<��S�m�};'X��睲E�R�d��*��P�ȵ�u˻m)׺G��S)0���:�	EmJ3-gH�
��늭�рPVM�}�y5Y9f*�]�� ���P���BN�AM��V�J�f��9�qx����|����,v�ܛ�.�M�6[Z���1�d3��vi[i��O�|%�똔nhԀʘ{������E]�\��X+���E
�+{zM��^.IM�-Kq!����.%Н��XX�I	{�����ʆ]��3}�Q��!/��Xk��Zǵ35�fSH1�N4H*�x��L�u�hrG�,�x^�v�����eZR��RfӾ�\{� &�5���e:�j]޺����!%�[�൴zY��μ��CD�It����nU��#SBu���tv6N�Zq�V��>ξ/nP�]+m-�\�R�]:�H����4�����N[cE�C�
�]�Y[�f�'wh�[q���ؚw�{�����j��P�AL[%��EcIf�����y�k��X����-�����+ �Uz��W�����hMU�Y{���}�o�W@���}[j.��\��S�:�w�F��8����h؃5���zT W;���ӕ�v_qt3Bظ���],�j����0Θ��7�V<���$!] ���r�@�f+�4V��[`I5ǜos��vj�w�A0����j�C(2�2,
�
�ZE ���`�+����ҡˇ9���.�C��Rc�D
�>�MԔ}��1>X��SsP�]ً�z��'�p]�Mj�1�W�T�咴�+��Bo#{s�7���o�ݍ��ҴND웎g*�s�'����M�o'l� �dxq���u��%��k��X�w���j��J�}j^bv5���\��DU��N�S|�!:�F���')����:�gWt��W�	��5�����r6�7��mf�,N�%%�K%Ȧ�:�7�rϬe����v��V$v�8��N�L\�nŢ
��gzG��Gs�z�W�KggYL�v0�N$�wǌ�>d��ϕ*�Fr):jEV����a���Y/��_�j����5�3��p�c�1�k��,�r�w{�@�=�ŧS0�|S@:5}�S$FåK�	x�;eC�d��kMr�R��_k�ܺ���D:�v�J
��
|1�z�.;e���UK��ܭ1p�2�ٝ;��8� .��q\s�7(P�L��J[&�;�H1J#���Vm9�Y��+�lP3p̃��¶:�َi�s��]nG"a��FV+sʾM�+��l�;S�y�z�2�����5�-�(�ox�7����M�UN�fk��jڵ9������b�7���6���#�*K.�Q�jV�W���D��3�`��[(��He�{�Y@�[�tq���2��/2�r�+N���LR��)�嶘K:u��Xp�p����΅�x�['	�u���f&��8�i��'Zůuѻ�ۘ�vh�i�W,�܉j�u;���6;�R+��d�����^؆3@̥w���S�`仞�M�uvys�ࠃ/���W���4���-AIS켩WCB*���#��
�,���#i�{l�}�e�媞E�n�>���>Ӧ-��2�-�&|X譝�Չ�bR&�����\�����=wk["u�*�}����]�y.���1��[���S�7�Qsh���rʳ݊�ȱ��C����<Yշ�{��Ҩ�[UƮ�7j��nZ.�B]=��38�=j�����}����P˅ 1o��K}9%ts�C������ƭ����me�Z���9v8. �O�fX2�Mw7gC{\d�WS�5���\�Y���ܾ� ×��X�y�@!�;�L:n۴���1��1zAQ^aH�J�{K��j�1b��u����
������x��q�n�L�;5�th�n�����[��~Hv���5���ۻ�#��2��G�6T/&��W���J�8���CV�u	��2���1�z��2,U��n�;Wߙ]zA���;z�غR���v%�6��zd�@I�
da�L[foM�g�:B��rx\W�c��ބSpn[].�N�8�&�;�}�=*�XՎ��g:�S!o�c����z��\*뺯�;{i�&��p�*�}�t
U�*V9-X�Q��u��8�6�9*eh*�w7v�QF��r���K�K�^F�'Cr�eL;�̘�
*�j�A�a����*>�s�܁�Y�@�'��X�4�xđ�K$<�i�=aX�x/���YN^żx��G's���V�C}Ck�z��P�m�)�P�ʗ4(0[΅��S��eӘ�F^;�I��")U�7_ndW�w�W�����}�;�Ĺ�e�P�D�����Vn��#���GR��n���YL�;���v����]vz[�N�8�$��x��;����P����ήoIʈZ��i���u�<�2�<��� �Ӓ������OC?*L���{7[cx� �&%e��x#Z�������;L�ڄ&�4�V�#gebXއ3���w���5���M��
�S��ǇKr��+`p �4�`���+�n᧽n��e������qr�4�MV�Wt�x���y
y��uiu@�\�4;�]b9��Ob�R�I��M����<D�7���(�X���β�b����_J�>�V�G-ei��h�֙�Q�6�v�wb}N��N������_H�÷��늦��jR������wz�Ġʙ��i�)������6ԉZ��h�gQ77]�0I�Է�f���L�����s/T3Vv�@1��Z���5x���$%�u���'�Xp����z/.��Z���hRƎ���'Yʹ�웽�B>,"8sa�7�i��s7B�\�̔��/�;�}��U��2Gho1V�M�m�f�����ܖ�T�/��/j�p��q��n��jjx�GHv���J��1ܝ+zi�P�Y:�c\�}���:�5�v_1{6�K�mo7�1�|��,��A��s��i����$M��=
Hr���q�v'rp��ήέJ���K�9/g"n�w��޹8��']D��.����+�T�B���L8���|f´�bt�ֳ!�ܗ�.AT�VA&��99h��e�������6�@���S8Ƥ7���U�����G�q�U�(�R��4r���4�8^ju/K�;�_11r뛔Ӗ_n���澯�������F���oK��_U��ֱ���	G;iW2rx)	WR�]JK��,1e_		�u�o����8v����r뭨�T��0�}fn������ݷDk��}aCVfe���a`�����<��ԍ]9tIfeȋ��J[@eE��-��iQ�>�5�A�'��\Xzs�æ�PWAE�J����T��Z%�����U��#�����
��,>9���W�J�����������b�n��=F����R�'��R�u���6r]/��;�AxTom�{����ʺ�`��+�ZQ��ӂ��Jt�Z:>nv=��i��Ѯ�+1^����"&c{u2":��|�m��NM��/,R��#�B_nY!���Ղ_L�
{X=��E��D��]�� �lF���c�Ȱb�F�}i`;wV�sj=Ua-�i	�ǝ����<}�B�y�W\�������|���2�M��] ���R���n�� ׂ��z�p�0����U�sB5Ig,��;�ɞ�ՠfME��&��6��F�ڟe`ge@��5��e-��[as���ԡK�XƦ9�+���P��d�I�ދ��HZ��^\�$�6�[;y݅u CfY��dJ��f`�){@�nN{����t��	�\pK(˵y{�n�>֬��㰷�</�(��M'	]Һ@[�v��è�K�ǣ��O��EM&f5DTHEUFX�deLDQDAE1QA�QCI��N��M5TF`�daPQ�e�EM�L�ELERMNX�S2VYS��STMU0�LLNYEIEU1STFe�D�S��XSAPMT�Qe�41Y�T�fe�QVc�I,9�U$Fc�TT�MQ4��e�LAIYaU4DUVY%VYQVNADD��fe�S�RTNFFM�QD�SM1Ude�e�fM�TU�T�0UD��M-0QIQ0D�UfPTDT�EDQQC�MDS%I�dAfd�јMQQ%3�bULD�Tde3���E555A1EQ4TIT�1STET�1FYUDTf5T�L3DRULL��4PQ4�UT�4�QTSDUDDR�TWw������JK��=e��]+����`H�r�˼;�8�I��Ь�O{��=��Guw�O;s�T%�MxF�ӌ��z�%3I�M�偻3��g�U��>�{^w�x�c<*="��U�h�����m����õ���u5񗾒[�ӛ�J��GD8��jH��o[бnO[��٤2q�u���=�'b���st�3{E��lruT�sv�i�^��y��
畽�4�;R���\:��G����� Y<����%�/WF�}���&�T�~��������n������ y�3��L9�f,���P�Z�x�Yեb~~�7L_q;6^'�����y���hRv�\sͭy����1�Q�m�>2W�u�z�q��7SN1J���+�e���V���f�j}���jS��~o.��el4fdӯ�k	�T�E^7���\�[���O7n!��^	Gm��Ok.�)%���=S�2���_�Z����z3���J���	��X_FX������T�5���� e
�-_WT�z�U���ڙvK�}�jD�j���>�u��;�|��R���q*�x���yq�Y7ԯz�<��*���]֔�V�f�z�E|sri��o`��0r-��wz I�NQ�B��	Q1"���`q�H���
�zV(3����DZs>z�.�����K�[�(]u8��Y���]�	�NW��.f��ѭ%~�����AS���Ώ�/<�:�(:.��I�����=��e]R;�;�:"�~��=�J�騅Oz�>Wp�Oc�	��{}x���cJ��紳�#�C��Y�g{|�M:����T'����F>���,&�|��Ԕ�-X���ষ2�w�U�y���t�uo8��uI�U���T[Ԯ��-��Y��ϯ�l��9�P��|����S�M>r'i��c\�oCKv���B����e��%uM��cgְ�2�9uh�qܵmuY��zp�+��JwN�/��Ap�=+'�uv�m_Z�OC�Q��F�s�{Ր��3X4�Xx�pm}�-XsV�a�y��:��c�Μ�mj�M��HS�M>�&�;i=I���p�i�&�L�շ:F�P`D8�s���.f���wɩ(�!���M�ӵ��&C�V�;Zr��ǥ��)u�r]��,'����9�[[g�{m���RjY��=�pë���i+Kgm��:�����}��M�b����61ޚ�,9=�ST��S����>�.��}��轹پ��(s�lsקǛU�po-)L~Z�����)/ӓ=E��9���mz^���TU�QY�O:��͈�	ƶ���u��ǹK��,l��گEm�	�^oP�����^�}�Xbd��!U���y��5��}�)n8��I㝸͝��O�A��ca�V�<��t�X�[�uʪ�nPN{��hYɼ¯�jV�S�k%6�F�G4�in��u��o/�+z�|�!�y��g'E�@H���,�'�!�[��ʬ�nv]x��\��{�^T��И�a�)OC�R�����<��p��c��*�q����ُ�,M}W/[�"i�r7�L�X�1�%�7yg_�P���C�=��o�=�z��̕��e�		oo[l��91�.)�әU�f8*i��h�3����XD��[YLR3wu��W�L��df��-�m���̠˭�f�Wկ�Qpx�wiN��v&��X��]��e>/�6���pQ�,�JږGd��67�z��e��{Eu�D3z{��nzz���%�a�E|�&l.{K��d=V��qeͤ��v���7m�����|k�����sp�"u�¼_d�J�k��'3���'U�t�q�6���\#.)8[	��7N�!�K�7&���m[Zo����0�cY���<�\J��_��`t���.�d�	�{r�wz鶖���e���ח*��MTE�Sǃc5@���Šæt�L�b��u^�Xz�����l�Xqߠ(���y�}YM\fJ��y�.�fV�H����ޭx�7%��\��{�~05��OYn����v��K�U�z>���W:zu�7=�JR:_����lTE��r"�mByۯ:g�T+�t�Ei����kNET�ŬTFs�ʮ����cMnz��*�!<�ҩ��Y[E��qr����k�'���7|���'���\=�[��J�-�ev�F��^�[1�zj]�i�5�7=���e�H��r<��,�l�ݷ�^vPZ�������C#������(1w*L�}7r�w@���ͩ�J�_q�h5�Z%�GwV��T��|v�(Rʏ�G*̅�wS�[wpLQ �r��p��]��u��7}���m��>X�ֽZ�b�!�����O����iج�˱y��q6�|s�ei�=�{��:�%�Q\{���1��K�7��Q?-�vy���2�m��91f=�P�N�y`�S8Vw�����J_;��f׵�idz�%ó�=��r����V��E��eQ��ͷj[��u��}{1ݎ�;f�"f��4¥Z�{7w�V.���WQ��­i^wJ�A�lCr��.zĬI��醇o5^��鮞�f���P�/b��R�*�����:����S�*u;�y�a��<q`^�H��{�k�8D�$�˂�f�t��*����>�l�T��s!��fn������k��친�dd��\�pWK���s�V�1�sMk=Ϻl�u�E5kE��l��?��o������r���RtH]��aV﹬Fhq�c8_k�_-�89yX�p=5��;��K)b2��z:����:���^��Ҹ�0�`'��J�K$��1�ԃ���'�w�Lݨ�
��sM50�x�l���f<��锃}t7��o�kث�M*2[�@ȸ@^#׽XWjy��s�z��9W��λ�<����X�������a�M�n�S�fywؤ���v�~����w՗�!��g����9����T/��P淆)������O���S���6A`k��]�s{~ƚܧ��@��b�]k��)��1����T��+[����޽��+Bwy�,��a�Ӯ�5"s��,�I�ܬʄ�M�z����*N�/�����i�\ֽo�uf�34�jYp�,��5/���S�rȗ<�*��9�\�ë��/P甩3n=�ս�	��z�8�Z�z.y��v����yF��i���Ԩ����MRI^��*{�q	�}��1Љ�&��^Toi�p?v��+�z�v�����T�o�:o�ӭo/�Ryj�,Ve�Om��v�k"^���M�$�l��pt�n�^S�$��}ըf�Wr�_�y�-�hl�4GJ�V�J��R��a߈��}w���j��;h��,}�����|��Z���h�ʔ�y�a[�z�ݢ:��ޮ�xݼatmx��b���^��+2��f<��Q�d[91D��c3W	��*Ks��熦�Wy_C�^��s�Q��V�Y��~��	9>�:�^���s��l��oA�m=�7
#[;}��f�WM�+ctAV����4+���V���\W8�EPX�;����s�#</z�~�ᙯ+�~��8��zh�3<��_��f}�Nlr�����-XsV��6ޢ�>���7���ZAI+�U�Vj�+"�	��o���h��8�I�ٸX��k�{�F ��v��~E��Mf��0��W��n��go�E�쏤����n?|b�\^c��N��=ҷk�l�ƾ���j��+i���v�����K�|����ٮ�{^��=n�j��j/�J��[���Y&Z�,�����Ml��ҳ+�㝿f·�"�V�ʘ�U�n�w�ǭ�����k|�-W���Яy7�r�TjV犝�G4�w]��or�v`�ԨS���ŵ�Hu�B����&�(��(��z����䥯VL��H؏y�sc� �����;���W�;��k�ӱ�ڰz��Cv0�7�j�&��(q�j���3����@X�E�7i���]�ގ\�i��;��O5���������O���y��gRvX��6T�s��}��P��iGWS����nzj=��.�Bc��\���n���h�~3Eg��:��-�S�fv�C�ѓ[҇g�Obf9F����pu����;ws�;�Cș�\�6����1缂@��{����ΐ�?{H�'V����<�)���I�Py6��]w�d=��r��qkFNp{V[��Z��nVu�W=�Ild���N6�}�&<�;�����ޙc_��'�nk�v���������xX�=bV\�9j05�kTBT��5�f�) ����SX�-� \������7�f��0��2[�֤�Ƴ��?W��4��9��j�[�<ho��׶zZ�t%n+�'e����!�1�1^���/h>�*�+)�ŝ[H�]]`�G��Z~vx̍v���T8[ӛhI�	���]�֮'j�_�nA���wwTى�[w�M��i��L�y���s!:U���V��hr?y��k�;�/{�g;.���60��bs��,�<�a�z��=��eY,�u��t�Zj4���Sz�T��H��~��<���~0?�'�\�m��J}�������h��9�S��·+�e�sb��}��k��f����=s��U�ӳ{�y��������^N�E��Q��*�Z��cMnE7�r�+��N�R�U��=e���a=獽�HD�f�O�`�w�T_$+9Ϗ-Q��>�9ϕo��물�,FK��љ�edj�ǿ �ꊷ�y��{G�+��	�޵XY�웎�n�R�����t+˯	�R�
�6�ˌJ^\ۜͧ/�.׽��f�ꪙ���\>��2�M��g&/��>�t�(�WQ��D��S}k��O���b�J��]
>��u��Evrb���������t���Nsvt��Q��U�Y����>r��c�M�ב2���؞Zb+v�޷
�8�.�+FLcy�U�B.��;��9�S�px�����&Ӱ���#=�S�X~=y�l:�Q�ְ�2�wAK4;�Mٱ�F��/;N#��;�V�s�ܧ�X4|ǜ��y�����P�+��G#�|e� $)��_
�6�]:��w��/p>�[Y�Pf��X��ti�$���ݳ�F��Q�]�Kw���®P�v��K��r��
���������G���&��Y�^S���`�>:��{k	�v�Y�<�m�73u�YڹX���U���'�u7��VLh���7s��W�,B��l��Y��ܧb�\ f�Z�N֋�/n����q�^�֍g�2�=�e�;|:+}�i��%������|gz����fy=���Af���(^�&tm��kj���N�8���G�[�=��ڍG�^�/7�NO(�5+�!�J���l�t��}�0�K�0b�W���Ң�J*���i���gm�&�O������J7��ϲ6v��J'Z���Lg=<�@�V�F�:=Q��U��?o7����nVey,S{�vv�	�Q*'S�+@Y���L�b�u[M�:�V]��pY~zu��ܼt+,��9yǤ�����pl��y:����:wl�0��{A�����F�M���y-��R�ҡ\c�5غ�=h�#�L�Y��mn��d��[�d���Kp���ӆ��O��ZA�l�re���;�77��d�)P�a��E�&6�R����A�3-��bv�~쿤�d�|'x��VK-�Tu��{�+;�n�8p�d+#�Xt�M꥘6��=ن�8�7&o�`�h��f����f��.�	R�e��:L5�C�I_b�F\=��ͮ�[����b�f���4ފx���$���6q�V�s���\��gk�$7G�����|7�"��ѧ�2��7VU�^�� � _|`�y$�˶4J�K���)q��/+����kV�,K2�+�]�RvU�7��S��Wj	�4[�L���yע;�f�Yɑ<=�Op0dg�x���ᇨ���Yۧ���=f����Fb�]�)�Z���v/��l���L�q�m�:�m.���Q�<�i��օ�z��lK��L�]$�0��8�J`���,��Bu|�4�=fS�W)o1�B��)��s���^�ٍ��g��@f��Ƚ
3�r:Eζ�}�X�9}Ԕ�c;GuN�E̼�I є���p����U���U���zZ����9*�te�ԍ�i�u[��~�hE0�ʔ/D܏-M�\me�׵�)�Lt2��U��B�CF+~K�{7t�0s~G�j�����!X����͙͜�;�p�WÆ�(�5����Gң[��ۚ������r�)�v��B���ID�ZKOU�{����D;��y���N��;IW�[�B�A0Jv�u���!��9�aYx�ɤ�$ݙ��3��#m�*����/2�#V��r�U���rnc�E��͚ODdᴝ���nQ6w��k���`��U0X��e�p��U]L��f�N�^�w��Wf�Q7c�j﹉(��W�h�Sם����H��9��R��2��pe�D���.�S�o+�uS]�9�6jk	X�Ӳ�t*��ܷ��f_�.�+�ꔂE��]$A�ܭ�P�8"�0�JWY��+N�6a��|���mk�(g]�2Ѻ]a�=�S�Ǟ���dT����N�r5��.����;7m֕$�W�KhR�0�ݹ; vh�l��j&KTM�k�W%K����Y��W?,��ok����&1@��كX&�c��I�r���zū��=���k2�C@S{Rh���B]r��\����ސ"Z��R�Z�t#列��9{�6�$`��
'�ȭd�U��A����Z��f:�{�%�$���M�kєd�����pMc� �k���G�7Er�raE=Cb>��W��]2;	��
Ǽ�p�e�ˈCvRZE&hq�]�s��.K��*�B��
�U�����n��t����\���u%���C�aRN.X�\�ۡxd�tmP������;{��n�@���}��~���<�F��Y���b()(�(����j	�����f������j���*
�Y�R*h��j�*h�i�J�
�
�*"���"��)����� �d��"�
&J
�(�"i��*������"��*��""� ������Bj��%�����b"�*�&�&�&*���(��
$��(���*�H&Z��� ��j*���&������R��*��)��fb&����)�(�
(��b*��*
��������"*b��� ���b�b��bh"(�&�"�������*�������4��ut����^�t��6o���W��FJ-	J�k������y;�#��֘�hYO�\��R��D���������$?.ח�O�[٦�'ï^�����L���0s.ku�4��'�ro�=�z{].���vy͝dz��e�����3��?k���*�; Buu-ze��<�F$}W/�nl;ꊳ5���]�+<>��r�ݕ���Sƙ���:o��U�v���]�)�XD_|��S��ny���ܬri4�&O<���2�w;2C�K>踋���WӰl��<�v�W�� �����äl��l�Y}�^��u�p�t�7�bU}j�����.�#.+М-��N2b�v��뢶��{��=�W�g��7��حD�]����AVzA}x�3GL�nj�)pҋ�M�.���|�t� �6��Į��[�9��&+���|�CC�*o�*�n嗩����Y�Z{U|�5�r�o���uo��pf9�������cO{	���!��y���y���b^�c���]`�.Ǐ(�;�w�
ar��^�/i����^���R+{b�Jy[Ԩ{��f��VS��{���/�f���9���LL.�$����3>˨���;�����n��l��^n.d�N�zus\5&�@�Dgq���(7���6u��zP߳ݚ��J�V�ƾ>�,ox���Ln�dzF�S�Y[ӛ_lM���n�V�Oj�^)Bu(�:�E.ʳj2��J*nd5�|yұ���&�ܦ�n%fT'�v�6v������\�mߌ=9���y��n�{Qw��Ш��9j�����YɼΕ���+vp��C���i�ޥ�[��S��+k����cؔ�z�>I�y��|3���-`�-v�8��[�eC��_�=��W��T�}k�_�%{Ӫ��Ǌ�^]S����I��fR����yF&G��Ǥ>�u��,��`ޅ�?.�A��d]�*�L�X�=��}��7�D=�R�	wСS�/�����t�HL��6�_S�6���s�%��6d��;�H��D��5+{v+�T�Z�|��u�ˤ�EĊyc'щfߣ�gZ4��]�ל�K��#C�&o�_�y[;-Byʪ#Yس�V����%.}uO8�w�Q;n���*�H�o���w�Am"�Bi��%{7�i=����ˀ-��{���I}-��A�R�b�Xo9lX|h�t.���"�W�zo�ӌ����Ӽ�>�?Vré��>��������~�땗/J�&z�O3*���K�N�WEnI垺�yn�����N:��WLWw5/T����H9���C����P\7�J�8����ۙ���p<n�m�ԁ̯<�\`�9��{ش_����zj9�ƀ���}*沚��Q�/&�ңA\1��je���q���v�jy��;�==�׵�B=���}�Hv���`�?�Ǭc���>V���ٚ��!���P�������;��=�|��t�G#�_g�~��y9)�0ܼ���=o ��vo��������u�y�\���艉eÉ��������"�{�<DX�\�H�h:��R�y�{%�dv�?I�3�7J�>o��K�؏��F�仿C�w�/$>������d<��Ϝ�#����;��V��_q��(D{DF��j_g��r?A���' �u��%��}��d|>�?I�:u��ߥw'�}�r��G�~������ީYoG}~�/o�s|��V��~��z!��\:��@���Γ�Ի����?OP������#��M�H�tw��y9!��'��]�G���roxr�+�в�ϫ�#���P;w졟E���=������_9��r���hB[��j_��٘&���޳R�A�Ԝ�J�z��?NHt���y.�f�r�w��IQ(&��SIf��x�q�C��pv]l\�[��r��U	:��z�F��=2�j�彝��Yt@aNdɫ��ղ !���&7S`Pu1��ۗ7.��ӥJ����̷ʋZ;�C��.&��̧�L�H^�&�o���
��/��{�w�<���ތ0y���=K�sz9��|�����n_9��!~�{֗RnS����~���0NA���z1_���w��u*��^1~c�˃�ߟ��nH�уޖ}����^^A縇$7[�G����}���=ǆ��>�q�>���Gpv���\���ߚ7��
N�Ȉb<�����i�\����)����tq_$�x�yd����'�w�)٘��|�I��ZCr�������9�I��_�y��=C�|����b"�~����#ŏ�wyV��M����}���:���xk ���w��/����%w�������ro�x}֐܇�}�@�����;������G���Ҩ��U�N ��sW������k�+�~�ޗ#!z��nC���r�/�Wc�#������?I��!��N�q܇�j9'�a��y�3=DDw�}o鶎U�����ޮwo���P~��)���~�����Ύ�y'���K��^��5�u.��2K���_��rG^`w{#�;<���)��nS�5���[�_���9���׾w��y�ߺ�GQ�>�ܻ���9�%��=��	C�;���O�ޗW������y�d;��{��z�w!���`w]�뾿o�ts��\����w��k��O�ԾA�y�\��G���
W#����y!پh<�p����`�>������G�{��K��^y�ir/��&�>������5���h��Z뮼�����s�~��9��`yg���ԿA]��/�r��G �r<������!�?� ���C�K��{�к��~huy#�a�9���������������~����C�>�gP�@�<�K�7>��R�
�}�|�pu���;��|���K����i�{�Ƕ>s���C�a���ɜ;�}YY��s�E4��3jx����\�8Rk�컼�`���\/�g����P5��D����ĕ���䋛��E�]B�L��T�䥻ܟtp�V�vE�MAe��ǲY�&��#���s�.�ۯqv�oK1J��Q�bQ�[�vG��{zoF�CZ;�c������yu#�voK��nB��<�����!�w�j]�KܾA�yy���_i�w+��o������A�q*��W�v8�x�w�M���,{�{�py������7��Hv��z�@��qi?GR�����}����7+���K�){��w'#���~��|�4TFV|���\eĈ���G�?�n]���n^C���sp���u�z���ރs��<=�?GR�����A��:�����h7/#$������}��\�oF6�U#�z�z�z���S�w'�G/�y'��<�w�<�b����;旒��x��zG���7:�ry�b��}�����ce�߉�,�i}�k/ڗI=J�}J�_�5��FHt�`�K�p<=�7.��~h��G�{9�<��r>��C���s�&J{����K�y	�oO�"G��@�?|�k,G{���W�%\C�5/ё�=��jOcR��kr�y)ۘ��y����r|o�~���^�ގC����|�I��_}���yI���U�����Y��C�����wԻ���0��g�F�;���O���f�?K��N��ܿC���Л�䝜澷G�C���p��{��]�k�WՑc�����_���p^��|��+�'����(����5/ђ��p��ۣܼ���O����'�}����7!��`��ǡ�D`�Q7�������K����_��}�R>�y���_d��x�u/��AJ�s���#���9&��2^�`��}���w/��NY#�CЄx��c���x%l�����_��~u����:��ܜ��/%=�~���@y�i(:����S�~���AH�M�ΗQ����I�~���y/�����w/����y�}�a��s =���y+*����\��Ń+|E�^)�:}�o��x.��d~���9Tuؼ&�\v��F��,�n��M��JAY�_���l�^:̮��[3msF�*��� Q�b�
�����):���)��4��L��)lw������7��K\W�1b=�"?{�'���S�3�Od�jN����rW�y��y	�bPn_`����(}���Ξ�y���K��_fK��v�{�]��ϖ�ҏ��zDy���}�z��a~��1=���o��\���0��^~����
��IA�FI��4%��o�t�#�y����Ȣ0����=y��W�ii��G��	��;���M�}�����#��9#�;��u/ ��9#�'O�h��G^}�r�2S|��M��d�n!J�ӄ��?O	��}Wu����N/ݫ�y�4����=>�!��!A�a��=�ܧ��x{��w�����]�v�_ �o����s���t�� �^u����({� �z>�~�y&��~�ӛ���_���+�>�އ��/Q��������<���w�'$܏]����;1}���"}�E*�}�f���]&R����湣���<w�G%�d�g�ѹy/��}�zC�C���?t/�ß{��j����r��y�r��GG������	g��D˾�������#�ϱw�y=�����}�s܎����9//d|w�n���\���}��~�/���#����{���=���}�|p�l;��%U����#�=��/:�A�^FHw��n]�Oo����}��]��}�r��G���Hno���4����Ξ�G����/��q��ٷ�|��=�F��|���O��_�٬5����7#���&��2C�0~����e7.��x��Wrp���?[������=����������.-qι�<Dz�~�{�ΗRnS�7����I�`���}��a���vu����bn_�$<�r�// �Sr�M��_������;�c@w� 
4�3$���o���(A�M�a�"���tS"�h��x��OA�[z�m�vP�e�=��䀀���z���R�[�W���+ۺ�����q`��t�F;<����p�&w���e>@F���x��x�v��2TsF��{�;jHs�h��E^�#V{�m��������o�C?��=��/�~���s�|9��%~��{�K�(���~��� �_c����;��Ԏ��X���N�tD!�"����Y²˦�R/�=������/P��?��rG��w�~���w�zMH�~ﾗ �z��<�R�.@nO��=4b�C������c�^ft�%dS����G��#��c��|���HrC�;7�}r�w��9K�>^��@����^t/�w�{��O�k��_�%�Xǡ{E�a�Z��>����3�W��p���>by��磼���O��Cp�~���!=����䟤<�4<���
|�z�~���AH�w�:��k]�����K)-V~���P�=�k���ۨԏ�G��������9~����{��vo��_�w�:��P��oIA�?����z�G{th�&g��+/�~�W�R��=�p>�އS�?w���^@w��~�ۨ���C�ט�����O`�9�\����䜑�{���zp̥��T��/�d����B��q���'��s~tw+�|�ޗ^b���4�/א��7!�>^ǇX��<���������=���>�&=� ��j�޾ݨ���W5�o˿k�:�����>��(M����/��s�hJO��{�:�+�{��������{�H~�NH}���X&�<���h�����{j�w>�N�i��ϭS�F�|���|��t�������ߴ�NJw�4���'���=�����}+�{=߽�^��`�>_�?fz>����#>�J��f��F���t�-��5����upL����������9�Wa�������ܯ����y'%;�7/%����@{��ͤ=�茈ﺣ�P�z�31�"������(��ތ7�a��'�}�k#���z"R�lCh=�ɬ̳���a��QPh��+�=)�n1�ث;�o�HH)�N�h���|;]%���{:�Uo�~����pf�Y�z��H�W�t;k�`7F�p'w4Y�-�J*�����V�ڱ���#��L����)�3���GR�`w����'�7#�h:��R������߸��nN����r�O������#�ѹy.����^Dp�h��oJtq}�%}qL�cR�����y��.�A��-��_ӓ������P�:��伂���O�ܻ����~��tk��J�O<T���}M������lg}�W�tL�7���]�����z^H}���zp����7K�?A�S�����jW��w�&�~��p�rC�1>�r�#�{�z.~7�9.������Y����_$���_H���d!��_�iw!�ϝsށ�'y�&�R�
Jp~���Y�_��vu���W�g���#���k:�3�+�JP�!z���x}�}�:�>�H�/{ގC��}����������z9�}.�ܧfsF�ԿAI�`���}�Ș>���1���j�������x�r�����W���'���)���w.� ��C���~h�}#Խ���r���4��n<��}��Ԏ���w��G�b"G��@���<M|����=�ӏ�}� ���9��O����%w�~�~���{�I��9g9��p?@s�>��ܿ��>y�~�b=~���@����
�����~�ǋ�w����.A@��{��r:�>��}���%�=w��%w=�~�/e:=�p����u�7!�nǐ:"#����E�{�@G��{o�]4�Q��u�A�<�ם+���#!}~�[�P�9.C�~�˫R;��?>`{d��tw��r�S���{���#��J���S�Ug���]��~3éI��(5/�SǛ�<����z:�䞻׽.�!z_��!Ի��X<��]Z�܇�����N�S��_����c��~��7��T��R��;�J��&�C
����kBCEek=x�P	]$��=�Â^ʺ��9�n�{�z���qF�����5>���foh��Aә�����t0o�����A��(����I�0���X��ܵi(v8���z=��+���Y߻��u)��I����C�Gg7��y!����ܿ����hJe�w�:;���4�����K���!۬��>^ǝ`;��u���y����f��f�-�����X�}b4z4E�y ��ܮNA�=��)\���G%��a�h<�p���Ϲ�(K���tw#Խ�sޗW����4���k�_r5�3����]���[M@j�Υ7!�s�=��;���C��]�^B� ��������7/# o�|�p����bK쿏����uu����}ެ��i��l�{|�]=���Hc������"=���nbrC�>����	�u��Լ����/�:�pWg�/�n����ܯ��ߴr^F@��4�%��]~�<��95�.�w�l}�=��ض��p�F~������irm�w��)�Ƨ��C����:�pR�/�r^A_�?C�:��w��8}���s_r߇ӕ��
��W�`��h�{�S{��>���ie���B�!��{��j���-'��_�٬w+��tw��)]u�A�w/g�?C�y9h���~�F\=+[�?s���k�k����kz>��w%�K�����>�Kþiy�?���B�!������J{����5+�F�����o�Gy���y����ofp:���o�~���ߘ�%�sz9}�<���;���!�}����4���#Ǯ{�<����7:�r{��Cpu/��/�=���̴��ӣ����DX��#���"6_�$8`��߸{�n]ɿ0��G�szy��|9��>���|9��{Ѣ!\��#��I���f5���Ͼ�޸��R�'�<���#�w���u+�ް7/ג����^y���ܟ�_��z��}��?���X�O��1=�ݯ���jb�P����m��vнm�{�_46V�k�ؒ&�Ȯa���!c�2p�귻�������x�7j��5X2�.O���T�:�ȅ��T?\ݳ����q�`,2L�]WoK0]Z[tz�y�\8�����6c���L��&=��W�bѷ��#���F�e�QϷ-~�H���߽�����{Ӹ5.ठ9��8B��?F�w;��yy)A�~�����Л�䝼澷Ժ���]}������u�M��E��b#�>���/�ܽ�߽+���އ �z��<�R�.@n��p�ܼ���>�sܟ���S�0܇!���'q���4c�S����԰[��==p~��h܏�s�Ծ����pw/{�΂���\���>�G$ԿFK۬p�/�a��#�G^br�<�F���H�l^�}X75q꿭Y~��${��3��d}/�_m��v)7����6D�[=���rT��B�Zb��{�/*��nŬ'�>�e�'a8���C���'*���gBx�wr��RAL�J}U����0*���Bp�Ts����SǾ��DM.���p������=%��;�9����P{���6�gf�V�u�M%U�Q�1^��<94�f׃�ˉW>���#6Te<������HZ�z�Q�K��-ԃ�ZŻ��Ts�5�6V���{���Is�o����m3���S�a��9M_�6-��Գv�����;�Cz�`~�.T��#VT�����j��llL�M�ն�o]�w&OC����5��J�o��Ӛ��a��:�@�-�X}R�~=��[�릑�ڥ�;���U�Mul��YR�>#��]qN��l�ߖ�Ki���j�˘�eũ�����HֲT)G�Q;f�\	D�ju#4m������m���ޛӝ�8d��G`Wc
ְ𣹓�s��h@��C9[鼡<�,����v$,V����l�ގ�
��g�<��7q�X�mܢ�y	�,����2��<�nT<��u�h �ɔn�x'�:�R�&9�Y�Ω{z�N;�.)�c7�-����|�3Ĝ�����
CErR�5O��83�h�����Aס�L&cT\(j
&8��#u܍�'���π��Hw4=�/b���dW1]�"{,i����/���\t��X�T�ѝ2r�yh�~Ö�j^*8���U�$|���W[��`�f�m"]�����W�-޺���)3��u;�Y��Bց�r���kSo`���ٳ
L��MK�T�AN�Q��մ,#�K���R��:��9�]R��c+,9nl�j��M�U j�Z�cZ�nB�V`�;PCpL\�e�u�����$yju3j��|e�4��L�ǅ|���N�kB'^E�rPY�|��9t�bT��kn�1w�/��V�1�ܚ��hV�
}z&M/� ��!�1�w�,�!����L�λ�wideK� ,�>�Ar�0���F�`-���a��!�h���[\.�)�����U��[:�����M�(7���:�z,���WP%&>ډ>�o7N<8�k�&���O��t�c�ǯxi��aJ�-=z4��L��f��c���vTu����M0$ј�I���Uw �=��w�qt���3g��
G��F;N��'n��l^D����=��{�v�1��h��Y����Prf�AIu�+�Z�.�s�ȱć�UJsi�9d��O�	hǫ'hF��
���	����"b=w��9a1E���S�4�����m���YYh�Ȯ��z.�퍦�k�٥����ufYԮ��)\��q<n��-�O�����rܡ�t������R�(�RS�Qw����o��e✭+��>��f�K5
���ɶzf#��Ŷ�\
#x�p����K�X�7F�N��?����{6�'q�{�޻��/�lm.C��c�vֲ҈d�x5n�]�2&'+�ڸDeK��׵�%I���<���	��r����J�%�ӹ�(az�Bw/'�DPp
	�>�;6c.fN9|F��,����w���}������W�8w�)e[M�3���o��o�����Ye�NiN�Q.kz���$p7�f�d{/w4�i)�k��wԨt��<��uJ>]QZ>���d�Ӫ師��p��v%v,���B�P���&���*��"���(	"�h������)�j"
��j ��&�j��&b&"��(����a��)��j�Bj�������
��d���i�*�jZ$��i�i&�)&�(����)�)�(��"&!�

&;�20"�" (j�����
����b�"�����hj2r������
����`��b)�bJ"J
*����g0ƨ���!���)b�H��� ���$�������*��&�������b*"`)�j	��"*d��"j�j���*�����
��"�b������,�*�
*�".�������׸�׋뮦����U���;uw��*���`z�:���X��l�꘲����)e[q�5����MUW�W���\WO;�_�j.���JvU	�� kyp�ke�Ε�^��μ��:�>yi�>V���ފؿN�|���1�������Y�	���WVJ)ˤ�Qܚ3=V�������mg�f���=Ȯ�o\'�*v��=i�	�5>�-wPY����e�EF��,����\-s�Ģѫ�����>\e���E�}��G;���t&��NLX1������sa(���*U���Q��O�����N����N�<=Q�T"}��
+��s��i�^D׎d���N�[ei>��,��-���)��12\VɤP"e�&ehB��ij��v!�%��૆f7�q��r��Kc%�X�G�ٞ����r�V
S��W$���:�(Q]�R�}u�VǨ�R��c�A>Ú96��=�r�Z�U���un=���#�.�<^��O9�:�J^ߗ]�>���S;��Fܴ�=Z�x&<�p�H���t��7�m�u����I�\��Ʃ_]�
�%@P6]�z��'b�8�l��#��ᬎPU�3)�bsk�YW��m����_P��u�Κ:��%�1�Ӵ��_�����o�\�P�۔p+�S��~��=�N�����s3��:
�Q��N8�0�y.y�+����y�r=تK���BV8A�j���U�5��g��q֜�xq�"���ªVL�4-u�����~̝���1�3�1�o���k��b͙��3y�͖-����r�vk�d�������W���s�����E��s�K6���_7����m�}��������`ޚ%u��z��	��w��Ώd�;v���������>Ɩ�R)�ҧ�ht��z�V?z���ߔ�	ϭe�61W�|��:㯷	��<�K{�+*R�c�gh�u�4��_%e��5�t�
�ju.�=4���O��+zu��������*	�Q.y��X2jQ��Ĥ��rVD���ˌjU�U��de�F\�O������<��ܥ���)?-��'��j�<M/w1ҭ�V�+��UDc��֓�-T���lP�#�U�jҋJ��8Vvf�vw��
w����MU�.�:�h;1�T�Uq�����b;$&�Y�/FJ4�)�ݗf�7ˑxmi�Y�>���;���PL�-���O���3���*\�X݋��)ͻ�ld�
3���o�z=�F]?��_=K'L��+���e�����]$}�%��6c�>r6}�d+:�X�|��eE��֏��(�=���]���O93Py�2��a&D�����N�j��6���<%�nsϊ���A�p6�<���[���t�z�Eeu�wh=m���������:�Y~/�5ڣ�A<:�WE���۞���������R�S��\�'��;�p۸�:��y2!<2�X�9����ˈʵQy�����_��:_i�pz��][��Ǽ���\��=z��ʤl��[�w5�]v�9���LRv�\s͸4���bm�:�*{��r{�<R6����Fs�b�L��������#����t��_��֝|��^��Z��f��Z�ޔ6%�⢭���Ʋ*U�V�%�f��Q�s�f����o�~䟢��T��P�t��^�nЫ3�b���fxQ����ڮ�մ��W:f�vF�)����;��Ks�I�w��-�YU�]F��wic�����[��gv���]�ҋ�;9��e�!\޲��f����S_jCgX���:�ŵ�gv���d�����;1�諭�ﾯ>����,�ɑ��'�+����OVz)�ۉY��N�Fl�A:�\�[���v��`l8���MOZ|�5|�,�޻��*�6��[@uT��&֞S���55Fk�����=W:>�������zėj[k�q״�O�ֻ��BN_��mC�����������7�NwJ�)m��B�%������c�	���>����s���v̕����M�<}�$���8�Փ�/)j��]U��;��gGA]��
v쨘���������OS�N�\"��9Z�UyMæ�	��xW���w�69cP��~\�0Q�Y�7�^|�g!/5������C��H��뫴�Փ���o����{��g�
?z2�8Y	ů't���Md�J�ٞ�z�'�t��GGG�\�o*��K�:� i��� ��w��������l�[uC�@��X��(.W���k���t"����rKˤ�%�9Җl_��D��5���c)g�>��Oc�0<����M��=!,�~�lk�*�c�2h��娗%�,�[]�w
`u�ڴ"�Ϋ97tu%ۖ�-��J7L�_W�U_f���Η���P�ވ.5���_�\�cWE��uR�i�ক���d♞�ִ[Q��NrÓMFm@yy~�u���P�h�(u�3c�润R8Wu7�^�.mw�ڞPj�y����!�N��+�i�M��-t&��^�I�˅͊���nR���{�����H;8�yK4�y�q�W��T��l���������4��7�q+1Si�+<)�ڠ�Z��*�_���\&��ÿb�ɼ�"O-�Y�=�ȇ�^�b�s Cl�\��T��z�z����!��ƌ�z�P��.�,�ήJ�ިg�z�&�;����i�Fw�<���-�we���S�植V��TAHҁd�D��U��O���=�O`�[�x"�Nc9�)�!�j��7�`�<��!
ج���h�*o�g�Hq���>��o.;L	���s"�Qd��5�_e��/%�x�j�w��/%SJ
�_0���;3ަۂ���v�XtL��$��5�&N�q�Ň���8�����xk1C�{W�'�Js��QB��o����r<�r�����f�r�_*�e�)g<�3��C�I��굜@�4��4F7:� ����Ypv�cMvj[c�����_��Sj�u�~�Q5d�(vl纥��OG}A�����u���A������XW>>�w�f�)hB|�h�)����t��3}X�>z9fB�C-0reB*�ۚ�y�p9��;1���5m�B�f�7�r���SY7��04�9%�j�f�eJڋ���+u]j��!�8my�P�-NP��D����j�T�콦.3gDTb�'ӹ�u�Fޫz�1���6��2��'�G,�j�;�R0ץiGmDxm�x[�=<5W�ry2���B��+�f�ʜ)�6���]��i��`h�םr/��ѓgnc�dnz��o�V��t��'흢�������"X6V��ߢ��`zk�&v=e�3S�`dN��ח�ݧ9���~9:��J�Y:"�6p6�D^Fu6cN�J�;�V���	<�T-��m�3���J�n2�7�B����7(:���d>�za��F�K6!&wV�\֞�=G���Uo��f���q�mLT1����+i��h�{���Č��I5p�+�OY�b:�  >�Վ��N��!�H|�J��$[��y��n�IN�:��P�\G����B�F�<����+ޙ�.��z��Ӑ"��x&��u�n��uK��6��Mݝ�������y|�Y���vh��ǕF��KJ߲\<�\��s�6VB�*�������Xլ;�����^�V��a�zt�e:�q�g_�Z�z��[�d_�c��̠��rOiiO���}�2.�k�VG�v�����ydtO�Fi�#>��sn둝TX�.�;�ޭ�����=׺i�Ai����̪������^��e�+���#���a�=�,�Lv��U����#��.�(i���W%,�F�����w|f})��s3�]=�祆��<���.w����7|�P����b=�'ʗ���d�p珯x���q�z�d
3���J���j����"����5� D����7�/���B�Y�P�N��c�3�R�Ukx��r�F}���]�-|*��;*��
�!�
�nT�8)0p	�^c3�ٖ��(O�OMF9���],AJ���NB=	�7��.�N�d����:�-x��[�Z޷�T�(㈩ю��]-fE��Ȓ�=N���^���)���{.�D�U2O+8"���cxj'�w�ܯ]hQw;�n�ԋ7���3/`�����n�b�Xs������YJ������`�پ�嶻m���wk�Br�뻧{Ȭzkz�蹉Jj�`k��%:�/�]:�y�Օ��'���F2���t�^����x�r�������G���ͮM����G>�$c3������_;~%]��KV<��� ��L���fu`�� 9쳛��REQ���5k��׷:hZ f��s��g�b>�[����+���cz`��w�R]5�9'u���V�n�jtu�����|���^��,����E}n��F�@ܬ��p�^eMj�2��	*z��ᬽ7�1��X7NC]\-�F��#�v%ᄹ�U�ފݽ���o#���)����f�܌�y]��U=0�c9E�c�j��Vj����佂�]y!������]��qY@O�� *,�H	��-�J�L�q�-2/R�>*��A��+5��_�;�or�Fq�-Ld�W�)T{ªrF��՚�����^J��~u�#|!#!ùׯu����wBak��T�I\v��%I@�������yf�
#��*�B;O\�m��~>t;��G��zf E��o�Z��2ݮ9�:��J㬴}��������kO���,��=2�2��}+I,�a�^J�K#��譔;����>�u{�x�m��+:��t�F��\j쿧N��ݐ�N�'.M��5�c(��&�:ES�������������S�崱����H�IN�kw0�=R�W:!��,�4��odA��4{ݏk���v��NhP�En�Ej6��{������P��ԣ����1�dC3*!�vr_�p�s�~�	��5�ĸU�yj�C�g���Z/���i�x�ڄ0�-��rǻDY��$�k�:X�`����[RHz��J��,��[�Zč�%螖EXL�Vt�ʋ�,oW��z([�������ּ,$Q����[�H��ܞ{s�����RL�(�j�R��m�f�q�wT66R*�{	V���j���϶�$�>��d�5�	HO��[�j�{k�[fR��y7�a�1W�-LP�IBxx�~��5vf���n�;��퓜����!ﷰ�+��j��e��V�I\��O��p��y6�j�_;�v��:��|�6�İl�����C��-;��a��g5 ��\ ��R��In9��f_�{w�ջ�DF��y��b�6Ա�id����^�ʴ������o3}�鼔,���u�@O��2/'C W��U<��d@�ONz��Ӗ�p杘N��nir�ar���Ճ�6�
�*�3�k�_�u��HϪԶM���nxt���;w]s�*��;��#��;�e@-�B����g����0g,�ź�C����^P���c�'���e�<3ثn�c��<��Ĺ��.������cU���S���䦚qK��k��V(k9`Ǯ�_r���1(���8W~��������7yD�5�1oO�Fݺy�@V����+�J��T�gW%���Ǯb�G�/rri���k5�����]hc�/T皒5\:�C⑥�J��r)�G\J�'0p0��4�@�U�Y�E'H��B�gB�9]w1�S���G��P����8,}±�<yN������gޛ��d�=�7��TC�WB��1�c��zk�ƫ��c�Dݎ��Z���=�Ps�kT���+����mXJ��w\}�.r�ɔ��ó*b�/E��BU����u�cN-)���/:�"J(eo���ɀ��8( �f����*��Ò�ަ4���:��F��S��u�ڹ��&���'iyp���ja�b��S�]����� 8چ���������L������UDC��Q�1�OLG���s���`�b���z'{W)�U�&	u�ّa�P)8���:�C��#{A;2Z�g���ܽ�͵~|�x�~a��~]����[Ck�ۀń0�G;Ekι���hɳ��p�����;��;3��u���f�c}�6�=�)�_gX�霩a��H�	��,
OM��l���YQiL���EZf̫*���k(_V�ç*[�I�ms}9 �T��=�EL���<�����Ր�ȁ�]�&�7sf ,�`�]C[i;���S��2���;�2���x�b$��Uue�q�{��5�ޖ��ƶ����D�Ln����ݱҜ�V��������K/X����b�r��`��wDͶѷ)!&ib��i��9�>4i��PƯ{N�fn�.q�A��m҆�3���S����x ێ��a{pG�9V����Ʒ$�I��wu#'��ˋ8�Ue�#�uc���G|�L�im�)�qn�gx�n�w�Pt\�}��Ԇ�hoJ"S�����_(�Ng����׸���Ƹ!���WZ
ɹةm�4�
����t�CI8�9e$М6skn,�X(�9��K�S�\M�Ԛ:���
u����Y��7B�8`�;�j9��A���ɛ��n��B�hL0Z����fQB���W���pS�=S$a�uvr�+j)�F��b=�O�r[Y[n���L��m�OLnS�p�h��tչ3;Ev�u�}<��#�6�WNY��	<+�K�08�6.�}K�������1��`<�(���C[h.�0����z.2�0sZŹB[���J�����׊)�)�zi������2/�&=vi�Lc&
o�F�e��^��L�����f>��׻9epӡ'H�N�C����%r�m꽲��x��;@�o����)x���b}7t��F��������3O=��:`�����5=��u����@��n����9��
�D�B��&�n��Yr��t�h�Е�0`<���,G;���X6�Zǩ�� U�ir�Ԡs�ѧ/w�����`uXt�����G3e^(u�\0GZ{�����IR=B��W�nMN����2�̚��23��[Z����|c���q-��.� ��^��J�~�[Rw0|oeJ�(y"��wn��*&��;fU���d�ҝN�3q��̳���}���P�79�N�O�*j'}J�����F��8A��cFA�����>	�FC1�W9��jo�n����#��9���F��Lτ�����JV�fR��G0�J��+�
o���i�@�u}\���s��<!��5vv_c�Ad�5ԗ�,u�W!&,��e3�����'H8��>��j���j�4��X1��WfAWK�Un��-��8�q���.����v>��+�{1:O5]�]��4��8k��]J�#--�[��i���S�i'��.�n��PQ��ٮ�&��oWX}���]��̫V������s�˛s�*�掀�@�h3m96L�.{f���}�%�����Z[;�f�Yܜ��Wf]r�qQZ�ܰS��p���(C� �&�)�i���b"��+�Ɗ"*(���""�����*(��� ���(��0���©i��f!��H�*20��rB"��b�"k# ��#,fb""j)����� �,���h��2Ȣ�b�f(����"����&"( �*��
(�����(�������3+*hf��&��
J*��iJj*
���*(� �'*X�,�j��b���
j�
���h����p���
 �)����r��i31�3&�&�"�$�!���Zh�hj���%�0�*bi()�������1���l��"��R&����*"�����>�{���@Fc��������_9���v��3�!]�xݚɰ�\<&Q�b�+�b3�O{`�d-D�NjJhW�G�"#�'�o+��Nȕ��(��ڦF��p4X��1�}�-�"�N->7�(�g��$�V�V��=�=5F���D#�sb�	��D\GN���a�5T#3��a{v��h"��|�7w��9�a��|��v_=�X�_��N�e[������x�<=3�M�%h�~��oG��]�����dFj��.ܰ�^\`b�gF�1^*c�P�B�K���\y,�mA^���C�?+��p�Sv$���:���i[��s�!�6VB�T�<��B��]�U3�10fQo"�SP"A%��Y����X`.��lf�׀G�}�E�\9��"�ݧ{u�w�n�jN�jʓb�L���Πj6V	X��\@L�/���=5�˹E�A�)�V5i�$���X�i�Y��λ=����ͭ"�.*����m_�q�[U4����:����K���>h�W��`�f�{:١B���䥌�F�����w�d��3zs8�ɏ�)x���ٺ'b�;�{�|A3B{,E|�+i#�j���Q(o��~ϓ�%y�U�m�N��ٺ����{]��,9��M���u���ӱ��\WrI}��ο��]�*�e�wڮ�8���������AGҹh�"���l�Ԕ2�F�>���ܦ.����def���Z�!wb[�R�V��#��r���n]�\�[뻬�GC��b���t�J�p	�`
U��h2��i�[�߂@\%G0G>ɓZ-�=]���2[9�+���Ws�g
���!����Z����7�,v��;j���)=יt�n��Z���*ē�^ܗ�ew���t�|n,���3uW�,��z�wzw6�$Gfb�\z�=��T,k�L�k��P�C�P���߹��@����x*�1�Wt�YA� HѰ\���a��c��d�7�8{S�Db� �W9*��� [Z��.i����i�
՝q)�N�@�4\��%	�rZ7�VX���;V�fw`�+�s�m�H ��ݑ�&3�::���\F�鸫N��O�Ux�u�.��c!u�Ƿ����UQJy"��Y3�t3Ҩ��̱V�1	V��l*�M��\6��C��`,�z�NM
���{ڴ��c`Xc��}��N��:���Ӧ=�=���*��qV�Ɲ���rN}��٦���1�6� (pH���V�V9SӞ|%GgH����K�C-�����c{u�7Q�Ve�v/p[.�m�CI�JL�0����R�Ox��~@چ��>�vWn��%�l�ڶ�;�eڰ���!�����`��\����(�.�\�ZgK����U�v-1qtZ�3�wb��}��[̻Gy��q�G(��.��Q�<��}��UT	G �L�Y�Ń�_g�Fܙ��-����S�A,}q��>S�s�{u�aw<۳)wP�_���R���G�A�NḊ����<"��~<)���!����{g���z,L1��h�}Ղ?]�v��D<��_ԩVk������0��J��f1�7g�*�Up�7��\;�l[�B����Hnd�6׌L0����WYuW�Ms���+t�R�v)�4\71���go<�б~U�L_��bz�O0m��Xe�h���oH9��6�qu�ر�&��T�5c7q��##S�|m�E1�ھ˭��|�J��$��GT����|h�{��_ڵJ�ƪJ$x*��cyR�<���:X`׹��9z�<%r��O
�e�����U�>;$���!�[��n:sQ�<@q��ԁ�	�\\sڜ0�+�\��5#��v��{��&�c�[�z<Y��:TwG}:�����Y"�g�Q���\5#:l�nM1��v���[�ʍ[��e_Sv�aJ���Ȃk���Mӷ�`��Q��.=C��-cU�7T0�.K��1 Ʃ��]2���׏G>{v�e��r���(�딶nC}n.�� �ώDB�e����2��][���F�W��Z��`.��d�������G���;�����n�(}�F�z�-��`�Rɷ��W�4k:�śt/����cݶ�"�k;'����tW���x��]�:|G6��`���ݾ����g��
���'��N6KnznV��3G�Y�쥳=�ec��<��.t��0�ZDz&��)�|��ԙ�h-uleٸ�������i�����i�]�ϱ|sm߽֠[�n�t�>�pÔ�,z�+���%�D�Sq�< ��I��2�hؾ�MB,<�*z���m]h�Ng[�PoXf����S���5\C�1^)P,�#+�ƅK��X��޿-�=��*��=�K}<����R*��7	��V5D#b{�.)��fź�ۣ]r�t�N��yQ1���00� =.�F�a�&Ǟ/�w�l2��^��\�5��V|7o2���[;�E��I��dW	�Pc=i�Nmh�;�Z'ދ}j���L��D4��������h���E^�ۗ����"^�95���S�j�4y�d>�խ~F-
Hx$�g7�˷ O;y�k�f�
���]aJ(淼(���t�ɒ�[�s�{�#��q`�=����^4��ǳ:�Zu
e��OC�'K�:�;л����r�9����=8�V�_�o�i�ļ<Н�>��`�\�}��U_ri�ۣ��l��>W:"��TTG<�&*5�H��[Tƺ������S���̡켤b/�˕�v�癁�U|�H)�s��\�",�S��[fR=����xV�N�LC�6���[���>m�.�Q�&�
�,9D���fꥈL�Oi]=8s2?xp|D=<�k�<�;�"�YK���@����,�a>6=6Яf,6�n�7@q��5�v"J۾IoO*�<i���g=F.�S�gh����Ab����Ҷ&�ŧƫ+��ZN��F$�L���m��m*�3v�H����9'�V�3�Cd(����Uˌ��X����������vB=;�:5����"��G/f�@�-��Vz�i����f+k�gm���By��9��=�I�0���G�B��>0�D��E��d���vҲ��
/�\R����RҶ�0�"�穼slq='H1��+�T���S���X�K���~���@O����!oD��Ӵ5�=�.u,�
�AR�p�>��vp�(WZg��C�6����/�|��vT��q�ܛ���%�0�B\���[�����;	�%��a�b��K<z���{�
�טɳQ���ױ��B|;TWdg]wj����Y��T��ܫ2�Ite�Qv���ޏG����O�U�x�2�]L�d�̻Oi�we���~O��eо�l�vѐ9�M�
n_}~�A��3��`��������E�ˎV�[	ꀂS������kh*�~ޒ"y#Bo�#�'Ǘ��p󋇜Z*EOYޙA�כ�\�� �{W��ޫ��电g�<�f�<����'IuH��|�h��/����j�����mV�n�f��U�O��d֌�%�18}�d���<< ��y�R8-?��Ó�Y�5gj\~����P+�Tu�<���8U�3�C뗘!�ժѰَ�]�T �#wf�Z�j
��K�1�9Q��\�1�3��������Gc����,v�f��A�^Nk涐��/�VQ��p�n|֎I��Cw���$��qPR�p6�4�r*2��C�M����2,�ܻ�~G¯������]�L!u���ɦo�p:�����l�}����'�Po]-!��Z�e)]����xث'��Y����mo��~rg3��B�m����Ҽ�ީ��1����W��@R'��2����Лꊜ+��{����읢��u�;���{�lX��U[��r�/`�+�+��7Aqј�Ÿu���t�E�����s�hw�+Z�d�K�Q���-�!;3�+��}��|8���2Ѽ�h�
��싌{Q�S87�����ޛ�NN9b�z&���4��mj��xi,9S����g�Y���bږ"�ԫ�OgG5��\a��p�R��^���J��2��)�(U��,3S�Fbw��a�ONx4XWN��\dEY�]��-�MU��O�������+���5��g�@�&!����aW��[��>PH/`��H{�|��R�+�8�N�'�5GQLιc�*rF��v��W�����������o�l��t'����Cau"����T����3�/.���2׵�!��'�{Jr�55�8�ϦG�6 ��=�-�f E��m/�B����Ze�2,oU�(!�ʘ�E{��K����躘�|��;�l[�B��pG
ł��v:�@�;:sb{&Y[ڙz�n��Q!�X�U{OHe��SLh��4T7.��<�8z�T>iC�>8�n�ޥ����S'Ԗ
�]
��B��V4u�ms����M;?{ٶ����AΦ3�8m;�}���[Yp3�.�)Y��͌ДɾJ��Lbs᙮�]�ƇK�k����&l`Z��鏠�����&��w=�#\���×͂�o�3���Eƈ؇Ni�Yf��=���n8B��$��������ײ�T��t�|�2?}_W�E�k��gQvA��`hg��D��,X��*vl�:�����5"�]g��Oo�W���ց�JpW�.ᡓ$��D�7.xm̡&�3�H%�������d�.*'�t٘. �H�� �rRyW�{S�W���yp��o�Æ�z�Զ���y�Y����wI�X�s�������XN���u��Y��<�4}�ja�ɼΧbBel���L���".�T!`��똶k�\��L��=�; ��E{\�"��6�WFyAː���5���yL�ڐ#{%��P�^�8�D(��BW;�̅,2h��� �X�e�VW=���?rf~�+ħ9�:'�,<�������x �Ύ�O�s�<�9b;x����L���?3[�!�^�qo"�����X
��b�5n�C�H�W����ϱ;�r��57� �����]������(�_"��)������_;����Wcn�vX����O�:7Q��)�����RьKΰ��(� �$WH-�l����2-gu߹�Y�--�	��nJ2W��۪;��R<���:f$��t�4�뾾&E���f�l�{K��r�	�!5���O�o8Z@m��$�n��b������(���|�\�0�r�6�T*������}S�����c\�z��?D�"s�;�L1OH��7�`�<��!
{f���Ɩkk��V�S��f�P�F��x+(Ld��r	�z����})�m	�2�;�hX�՗��oV�@��w\����P\E[48�L�G�+i38.r��2��rm3L��y9�u=ðs����dT+Ol����"K(f�e���Q�pdl�uLf���q;�o���Oc��]U��\]��g��O}mY�����7��:�v������b�ܯ<�͡�\C
m�q��*�����l_���������=X\��W1R&g�Ϋ�l��W�3�%_<���P���qyGб�9#zV�v�ĳ�wR�k<���<����գ�����Pl�/
��c�d<u9d��M�ZG���J*��#�=�������L;6r(�н��W�@s�H������`�[C�xh���0��È��Ԣ��/�����|�]5�<O�V���Y�:�ޛ*�wyA��9;D��%B4A-B�of�l�����8NQ��J-戬,Q�붎� <��X���VB��2���N:�V:K�؛��o���6���s����p�q/�x8S�5���ܽ�T��Fd����;��V9���ۓ)oޏz);��HIo�Iv)9��{������F�]y�z��r��^��y�ٛ̈́9�3d��R�w�L�+�j�fCꇦ/��i��o.06s�t_�����SL(��h�E#��ud��׬Ι����]pÎ�E��}KOl[�dS��v��vN�Wr�1�0���iQ�wS1b��b|0"f�����\��X�!oD��Ӵ5�����kUC�e��|_&�.J�&�'B�\:U4�kK�B�6P��߶1�����3�R|�n�M�w��^��{�]�c�]�ܣe*���I=�T��Nex�C�{�eP���-Bvr���v9�w3a��ݕ�:DP�v�u[���ǅ���.u�����z�:%��9m6�Ue����Q���5����X��#C�^J�'�B����M{��,�+t��.eU�o'���؍1��'��(��3��u���<��jV�j���֭�P��M��:��6�c�ߤ�]C�=-A���
a��uw#fH�y6�^�DΩG7�����ݸ�=V����*�9�a�(i`���>'Oa6�U���K�r�C,��N`���-^�ӌ\k���v۲��"B���O�fu�sr�c�����`�����
H1�3<��{���zM�����f��ȶ�Y�O��3"�)f�`=�@�7V��Zʗۙ����p�>Cl�vz��8T-�c��}H��vmq���y�&�����h��"���/\Pe���Y8gE� �]�����H|���z6Þa�s�#g��&�T�������
碣��q2�q��#Z�zb;{X+�.�2l�Ӓ獭o�G��ֻ����S���Fv�����T�'����N�K5��z�4{(����ۆd�R�'���;c��5�)q���y�y}�xWsFS��O/��A�5��4v�mؾ�з��o_�P�#r�tm��e�v]FL�.�W�G�9��V�)�ؽ�W7rՏX����J�Y��2��*it��{j�"�b���V�vo�-C
}d¼�yYv ��5QF��ɔ0�ǆ����HEKƗ� �]=[����7K��ǲ���$g*A���u^�KL�9O�Oqؑ߸���!�m](N�ڋ�e�6G�ʵ�!����']d��ۍGo1����a�~�+(�m�����b\4]vޥa��6�s6$���oP��v�k{�c}mwd�݈J11��@4y�wϖ���B�>�ST� ̾�5<H�f�H�E���޾Z�-t,��!b4���Z�b��B��B�\���m�Wuҟ��x�(�Ss��� ���.��� FU�kY5r�
�#o(V_m�khnn_+����
�E�ޭ���P�E"��B�]�G`�Ǌ]��W�%2�l;��u��m�e���!���Fh��*��yI���^,P�V�V;*�K貉)�E9�M;��e;y��e�'�n�ځ�Kn�=�}�`dR���u�.�u{=<_b�([֦�+i��r�׀�F�eVGS���=I�w�3����8r@��A�N�7�� �z�c�[+.���۝A0<��bk宇+Z�L��ޥN]�O�v�����J�>�LT�%�11X���ڭXG_ECyh�F^�qο���.��U�YwS��W.ƍ�p,dtVǬ>A�Z��P�$���������̉���S�ؽ.�y�C�^�ݑ�h�ro'W+M���֦����f�n6�AKx���S����oG l�k��.,U�3WT����a���[+�mn�m�ro�\��SS.�#��Y�;��q �̘�2X���k���Y�A�}�ڥXz�|��t" T�Y��y�����-n\���O1oI1ӣ:�C���*+\�PJK&&
����G�WqE&��d�Y��,��-�-M�5j��`�l���ے�TZ���Z��-��vVK��g�������OY��zQ9��48s�6�tE2E��UUVc�F0T���-4��QNT�UAfFND�CK��Y����FF54SQSQTM5Df.MD14L�e��RD���E4Q�fDUTYYd�XMM�eX�Q��8U5Nf5T�a�����ae�dYYdDU6YEe�C�ee�Qe�Y4RQ��E4a��fd噙�fD��dfc�DAT3D46`e�d�Q�ٙ������d����3SVfU�e��Y���PY�ىDe`PQ@PfaY�a��DED�%�FDNCVa��YeQfP�K�NTS�e�aAUf	X�FY��fY�Ff�da-�w���ņN�T�jr	���C�ϻBӽz�[:���*Ct����3�*�z��0���y����#�r��g����d�sMe��͘�IA�Mэ���w�˚�1�3K��Je�؄�#�i�i7>�9P��=�ݏ�3��ߨ%��X��2�h�%:�����<�*����Uoq��JNs�K6z�SSUÉ�r_z�bWϦ�FG��E\"�e1��&��8^��/ ��2z�L�w�^%A���,N����g����:hZ f�.p@z�hё��gI��u�~v�v�:��	�m�LG6z��
ܩ����3kg{C�^�O��`��B�.�m��v ��K(1S�S���}�N�62u�7@��>��:;b��n�R�=[Q�n��k�3��:bV1�Ѐ���+��/;�uz\���a\S�=�6#�iA�Ғ�������޺���#BQn���`
��	xXAi���==�nOv������KlOj����C����I�MQ�S3��
�r�"��aa�QD5�{ZW�M��S�[���ƈ���^��BcU�]�b�T��*	�8A��R�~�(p�u���ke~v�8���gh�Z�Y2��N�P�}w�[`��!�Ȯ'rNv7t&_����=�9opU�;f�ZAR�����i�|�n����[�����}ْ� ��z�]+=�+�r��=��)�W���l���X���҃^<��sz��f�7�7�ݼ��Y3.o��8d}���G���HhS�{ƺ�'j�f���M�^j֌�Ҵ����Td;�bȁ:ᮛ�>�2�_�/�`��3{�l��$��������y�Ϩ2� ��1�{KM�,gb�cCf0kr���<�,)��!Q�"��z��Qkg8~�ڔI<"����b�b������.cf�4[sC`��Z�嬯�5(���F���"�\r��u����h��K�?�5�㊜a��5�:�j�[~%9��͛�n��j3=�3�������CC&Ia)���p�ˇ��]����3��5�,��{)Eޫ:A�U�)8� �@��j5�͘oȉXK(^mS$��BTt���[<ݮ�{���#t2%�I�P"�����'�����E�ӷ�jFL�O��$��[��{�d��c�ջR�a���S9���^�TɸǴ�,`�x�[�k-A�)+@����7�{o|��J���z�(|3�p��8X�y˱�:��X��hM�r��5�j�ޗĂ^�wn��;GQR���ukA��`��X&�z�ϯn��jhʾk�qU�Zo_f�D2*;�IW6j�
�&��B�2<�4H��;���qS[2l�1}��b��5�M�mf�:�oK2r,��nL�)=rt�k%�"Vb�%9���X��I�����x`jg��}x%:H�#Ə��o����ҫ��.8�eiǎ�t����
���+��X�`���D3z�K(��5��[>�h�N�d@���]I�#�B�]��x.ެ:GQCeW�A�EG��g���w"ki)Ι���,x�pS�C	z����1PR4�\�]f��$����\D흝�[B��|��ۉ�D�c��m0�<U!��0w�?5D!^{f�����^Α0g*���Im��F��a!�N�����O�j�uC5��bc���k,m�t����K���G�8�0)b�F����(D�4:�C�j�Cٵ�z陁s��-���s�<��Բ��׮��Vg`�����c���(m��f YS�����p��sd����뇶G��>��-0reB,J�b�sn�="�K*W\��5���?T��73�\��n�:���%.�� �'���\��!�բ����"@�����]�3��0�����m��Y^���
����3��4��x��Y���~\3�5�@�Ӡ��T��'n�m��4N�?�bcx͡u�5E�mo|o#Whp�MM=S{��H�����)ՅG������;�L��U���ή��o������Q�]������N��,�b�L�0��#�{m���Z��Tt�^�k��g�9=<%�ȪU_� ��:5����l!���#�U%�(�m�i׼{w"*3L_��J�xm�j;������Ya]e'���;|��v��h��7���n���E�����:�\kڑ4X���ة�Ze���q������3kr>�6��n;�dtw!C>%�,nw��3�t^���C>�",��F��`��
}��}�r��]�&e��wZ�zb���v��m�������mL_˨���Y�z:�7�~�H�D�����m �%Sqs6�Z{}n�]��=M�c�09���_wbi%i*��J�"�y*��Ͷa�z:�'(s�>��'hj;��(���.)*)~�	��n�̃��0 ���˩���VD/����;��=��q{D��g�)v��<�1	�j�Q��B��,-7Puj�+���0�s�=��ܼ�j��o@Ws��>i	w�J�:zR뭧�B��N
F;"
x��)�����u9Q�L���%XลM�F��ɀ��EG��NW�ɳ�����\��:���<�L��L�Vwd#&�K�+v�[�>/�N�d������5��%Ԥ2_t�����կF�
���Ն|a}��:DVK��]I��.��(u������F�s�����ܹɪe��d홂S���~�Y�M�ŀ��� "��V)?-ϨS2����?�P<�k�8�6�['��쵁�/�J�M��i����ܡ��,/��'��Q�.i���15�#%�T.5��L�Υ�zW�mB�疁8U�3�ci��1>�J��[ٕ������:d�a�іZ5i�+%Z����I:�_d��{���o��1L�x�%����X�����L?��Cr��߉f���z��� OՔ�b#�ި�x��k7�P`�:����|�˻;�I��ZQ����T��h�i����)n����rk���4�	�/y����!K����3��tۭVY'5����+Qn�n�Z��1tf��d(����{�E����U]�w������5�����^,P���萞=�V�Ǌ�.�����\,mx��Z�P�N�c2�`�8�W��a�ķ1oK^��R�u��t�	��-g?�޼
�^{����V8�s.&��A�W2�p��Й��g��-���/�	������M9u�L�:�s����/Z�p��k0X{���;5)�0/8#��l�(�N)�S�黷��n�Jk�&%|�A�g5���[�y��k3���(U��\b�_{�
��gB���r���j^i�P��W8�#���4U��u�C�����U=^ ?�����-0�����z:k�iYq�K��i`WP�Zt�/N�����c*rF�ޡڷJ|���v�	��KM|�dB>�<T�S�vT�!���E�a'�J�^]K\Ba	c������1td�23�=��f����C�\�~�v`E@lD�9�֦�Y���0��d��j.6�me=+��C�u1�眮���l^C�B��#�*悉���
���est�.�� 8��NZ1�M^R����p��a�K�u�z��'��3X�oѷ�8ȳ��T�����i$�TF�WU<s�N-<��N�VC7q�4�mv�.ў�T��u羻RϺ��ɉ�e��/EÂV�%��#Ik�E&�Xۨ�qS���{�Y��Ľoa~f��ס'��7z�ې#`T'/K�����I,"
�Yѕջ�F��ꊽ�ė
Vi�p��l�N}�gfI��4�|��oQ���y�2��<����W>�q>Xp�͌�x3���I�yoN�w�m!kgF��q�W�2��|����,�U��p��n݅���-�b7
��r��R|]��:z�3se�~�*�Ƶ�=�_�(^n���XwL���f/6؛<)�����ʸhd͘}�Xn\��Z�/�V����5>{��0A�p���G��C]�(��&��]��$V��
&��f�a0_����Zq>s���z�s�;����^�u��Z:��^Lz�^�j�M��rX�� Y��bvD.��o^N`�'6�����n-qx9�����
+&-��w��a�����P!��}�p �kg_1�>{.��V�2�����Q�u�~r~"Z���:9
�FM�CkE�z�I��ƍ�'��LWxs
�����yf���vi���ܨŲ*]�襙9��[��u�S�"�s�;@.�z��\r�1^ʻB6
�72l� Ƽȗ�wP޵��c����y���^��io(bcn%ak��;���6�J0�]���:nh`�^�u/�5�GU�	�S�EKi_����\0��yg�(�|�t�/N듻4����Q�:���$���<|`Aai�-�Ĺ��G�@�׽���SBk<<w��"�;f�U�3^���u��b������ܳ�|��h0�L����=���R�ue5е%UF����_\MVZ����ɺ��(#�2Δ�W���� �>x��Vlxn>�;Q���Y�o��j��
'�����Ee�p��R$u����p�z���r��2"�KS's�XG�ce��05c�DX,-70P���0�Ƽ��(rx���_�����oΑ얡}���es�ve<]4P���@�ʣ�0*W��xk�����cw��܀���r�Ԭ���)IfUpBv����p���,KL*bV�n��W�(��Ա���u�_r�:�����/�&���Uŧ
�#�q��%ݑ�B�[2����R�ŕ�z�篴��&߾oFUs�Ux��S���P�E��N%i�t�f��Xj6�7N������(�X%\�,vl�QA�m1��}�6 ��ټ,+̀��%��ō��;\ͷ���.���"r��)_� <6�[<-�����3� ���GY�������9^�UM(<�y4�3�EDkι�gic٦�\����l�/!O
dX���lEܗY��fR9���]��ꐡ�f�mH��rּ}6���芁B0�^�	m7D���׷I�Ȭ�P3����)݌ja�n����^-�C,�����a��l�(�BE�X�������i���lb�:�z2k�%E���z{��C²v���]ɾ�O'v�dF�*j�f�W-�[L�7 I�a�Wt�֯��\/+cY�+�s����c�s[��uuv$�?_C�<g}ny�g�J�J��GAT��hHdI/�������O;dJ��R�!S��uX=|e�\���4�N�1Q���-�T��ٙ���2�~������WZh��P/��JϚk��l�X��-9��:��r�����i��s�L���v�S�gIbp�Pk�2#�&W�eY�)���B�A=�|�[�~�m��mO3\|F��]�^O��T�|;�%���c�U�����Z�������a��Hł�}�"��>Sc/��:D=�h*R�p)\}��q�T��Wl��}�[�����])<��89;e�*���bEC�o4f��f�]<�P����1Ӛ TRz��^a�����/E8��P�_N���zi�F��l�ZiܡZ�,.�-�hE��b\���7K�4���]Tw�B��K��Ҽ|pUx+��8*>�1���d��U��ȣ7���;�Z��h��*/���Z:��,�!�2/e<��uy�+�'Uw�͍�oJ���ӵ�������}4�*8d7���,� װ�~�k��4<�6sV7h�.>�Zuvǝz�֜�ܲ�rǳ��X�Q&��m�4����Ȇ�yޚ7�-�M�&�2*�X�/VA[[1x�p�/4a��d�^3�����}�^'W�y��*�=yXZ�v�X�����n]��˺l�A���5!&㜍4�]�B�.��:�p�������-��=��[t�9�^N��5��5��);���s�ƣ^u��{s�� ^�͋)���\�є�ؤ�>�V�GF�������j7Jg�θ�����[Q�x/q9��$�9𝙡n^�}����^�@t6.6�����ZC�%�1�����=������uۊ3F����ѿZiv�ؕf+`mQ�eel��l[�,��T�3��K�Ka����/5�5�{-q{n����sN��,��m��Mu	613�V��,�,C�K;����fd�1����|%G 6tm�*�*J��*hm�I�\���A��m�g����Bk%Rbl�����&>SAy���Q.�0RT%i��A b3[8�]�7}WJC��֓Q�(F^J
��o��o�F2%/�ds�1,ȇ���Ɵ��WO{__��/O�P�yn�9R�Q���9�?X��зz�u(WC�pQ�%+���Tm��^
��g#�����D,ҷZ�M9#,.�}Cg����5�j �]�Q��q_>A�ڶ��J�L��K;*tZ�a<۹�M�@ь�x��:�iT����}�1f��M.��E���V�K(�8�9�?a*���4��BQ'n�1?nm�������<�t"��G$�b�7` ;��>�R{;nDQ�D����cع�/��{ĳ�A/~z뵆>с-lC�L�͜'Ӫڧ|�ݭ3��C�G��OL(�od�?�33�v�6�M�m��6�ĳ�����^��:2Y[
�eg|���l;u�,�#�9�e`��gn�J�qO�CqG��ʈ��a�s
�e-�y��N�@��#���^���/:�R�a�i�X��(�I;�gu��`�סf��h!��TsNγ0	�4��[\���;��^5v�-���R�`�%�#c�-�\K�"^g=�Wm�k�\q�k�W^u�(����v>6��unC��ucP����?g[k�_`�S��
��UȰ�ʕ�q�v�l�
���T��w^�]	����:5�QC��n+�؄�8�� �aX���J�]���_E����Z��R�"�}��θ�e��e,�ЕN��}���}�͛Via%�$@ڝqF�����;mB�p�&�VQU]��)�O�����7\Or�:�V>C���)cm��R�\녭�� ���(��������%�よ�X���ڛV��c)봹���Mu�a�x/�Q��?$�ҳ�5֓t��:O��!�j�
���p�#������}el�^�H�X�5/`���}Hÿ�&bT�.�!ż����^�Ao�5�X�4��n���Ы-��:i"�~;�o�+��@�{��5��J�����Q��rbur���[gq�0Ci��W��;�e�����k4��c�eq�+�9E�u� ��ťc=��9۝ǀ'1�c�6�MӏX}��>�1V�H*Wf��F��>��,��7+�#�����ؖ"g���ș������í�AUم���1ҳ3U��X�u�u����w4%��P�&r�]���R�x�:�����e����1��G�_Ss�S�۾��+ۼ�Pjh*}X,5l��%��/ML��.v^��Ǻ(�M�]p��a���vި*d�N)|Iw@B{l�A�P�D2�Ł�U��'���*b�<�E�Z�9jz:���ջ�Y�g�Z3�������+*t�\�ǁ$�s����j��U׫�P8&)D
��U����+���v�x�U�uWݩq~�mg�跇��j�+��P{�N�=;�����K�υ���1
��v���;j�4��8�X#����RD�ͪ]�5'���Pݦ�s&�r/"�̵7w���oV�f�a7Dئ��7�jv&�Eθ�g��Oc|��N���"y4LVX!qǝ�f{�6PH|RG��$���d�fa��4�R9��X6aFKAfa��`PDY�PS����P�UVYYefU8a`�eYYa�dXQfU��bd�!FQT�M��Y���Md�cQ��Y���E�M�&A�fA�f9d��d94RfYf!YPaC�NX�UUL�Pd�4e��S��VY���d�DFfVAIf&Q18I�eAQ�9�L��f&�fSA�5M5���IfS��DNa��XD��ff%ef&E�df`4D�NXfd�dVCH�XC�LI�fb�a%dY��E��5YE%e�f$Te��Y��Y�ffNLD�5XԔe�EfYFE	fMD�c�AaFD5��Q5fADQQe��cVfI�ad�YYT41ady�{����P��ͥ�L�
�.�՛�k����^!��h��8Q�t ����]8�`+'9�:�a�E[Y'�[�Ix���L�A�լ�o]Q'�|C/m
�����u5x)\u�t�:�8%�������*�*��^�5-�у&�t8c�5��¢6+�)��Zq`��յ�γ��*^g���&zr�6;E�f:�Ꝑ�%ОN^����Jڅ�ԦE]W:,X�Qx⣚-gs��jG�ý��<YWA���"���(��lt���J���'È=|��c����H�FG��~�. ��q�����0�\����P��<���Gjp�@fNF^�;D�qt��M%V�)3!c�GM��p�.Сҵ���	���&��1���D�@s�(F�t�ZKg��W���7��s�LFU��!��ܘ�kK���K'��!���j�%�k/\������`��,ۡWΎ����Ni�^�^���VQ��۴�m�[�lFׯi6���\��{,�_��~����9�<!�u�~r~"� �Z�����L�b+ܔ˵ʻ�����	��!����C��0o���U�׭u�=N*��Qݼ��xgu���uĀ����h��>V4W+s�o=����z\��h�~u5a:���F��}�� X\��{�ݼ�>tww�^�״���Z ��{W�E�k���S�<�$w�k�ڱy�X�$�C���1�gVV��w�<�(D�[p�å=��|��0�m��bhr�4����oyO`�u�M	��u#���Q+�Y�ۆIA�X]qߟ	z��9窰�ň{}�mY����: AS�H���7[=%����l��x��\71��>Ȯ���.��N��l�'?nb:`�b�q&SDYР�G��=g	\^e��ж�J�z��4��a�z���o�ͨG�.gFh>�5�@|;TxRzs5�����>�kpt���@ܝ:��H�N�g�>�pL�6��O�;==����7�0X��	W&�[�!���H�
]��z��ō�7�R��B.�ve�	��+�Ϥ�$����,+�֯�w�^r�tu�hjߓ�^�� %�f��iv:���ӯ�[G�?6�xNVC�� �����=��n�f�#|}��������?	��"�ӕ$��T|]�@�Qr��p4�j�^u���E�ӌk8u���T?p�q53�Τ��>��K�J�_S��w��-�B��N%[+7��V02���g�!آ�����t�S��i�X��K�w�s�z��9M�T��P�f��7OAԕ��v^0���y
�uN8�b�d��b��.�b�6����vXdM�*[��d����s�x^7����,��,�,�eܿ�2�E��0;�6v�
�9P��Vz=^��- ��C^Kf���oypu�1p]�Kf��z!+��Eƭ��x��|�Jֽ�]q�*�C�bp���/����w*��"���dnw!C�w�u��o���{]F���B�a�t]�]�8����w��͹V���Pu)݌ƪ��cT�NŹ����h�9�:'�]����w1���!��a��f�6N�p/���R豱�,iΝs�ܨ_�r�C��sy�==�y��ӿR�aWd��u�Օ��2lr(�{)*},_�t����*.�fn)�)2����U���S�`72�w�x<1%�Ѥ+I��o�Y�{�Y�P��q��KӲ6K��Ƿ��p5�y-���c�;�f�*���M��T�[3f��Ov$���I���Y,G@L��y�����_]O$G�����$�\��1(?(��"�n�M��I�j+ql��0���{C��gҟ!F�zM��	�ذ�v��y*��%m�ȩ&A �xk,��@��,]���]o�V����24�fj&j%b�Vc�\�=��]�[u3}v�����`��]�V78u�][��H�==��=j&;�n>b�o04�/���۱���"vVZ�u��+�MZ�t%���e��s�zv�
������wM����B�	cCe��W)��Y`0�|1��ג���<�n��w��s�H�6���~��G�<�`���l�߰�����	}���tZjb�Ry��nǎ�]��uj�Gr0�n������b������j����2�ر��9����{�����b��D�A"������h�%t�Y�V=޵�1p�.�����9�4��±�����q�i�O.�!`�{d��t�},���,���b�pg�Ýrk��9�kS�F*`���G��K>�dXX�@�>{lxt�I���62�>r���:M�A��0#$�o�h(����2����ǵ��|�dM�� 	��i�ݞ!o��t-���}�s���W�'\);o�J~=VtvR��pde�V�1�X�rG=ź��w�t�Z����X�Ew���9�84�pbx�qo��Fg�� �ܢx��-'��S���,s,-�vǶ�e����š锼�U<�OW��tw�i��'���2�����+W��U=�ʏfc���hV�PX�u�üm'8�zZ0��Ns�Y�U/=���M�\z�A�ݤ���n���S[����l�L��86wAGUޠ�����uo)�+7��]<�eL֋�_9n垕dާz�5v�)W\��Oi�~���>����qJ� ���쩡�&x;��D�2ILo�;��1!3uѦ��7t��.�xo	c놁��bމ{��1�D�0�AR���;-�M.�����[W�#�p�3�����uדC���7�_�mH�uFZp��,Yر�Y:b`8&�˘�j�u�X,�!�6�i�+ު�����[�k �&��֚~l��_p�Y�`z�?B�BW|&_S�e���;ͪ�fe=���]r�w��T��*���Y|,9��7�� *�洙Ip�G��v��Of��l|a~	\V 0ۜ��N�Fz��#��11�e�Ԭ�m�LK�TZ):K�?�7,s���9�e���׏;���iԬ �\_��J$x�r��C�����I,\yH�����U�ww�&�X�ح߻،f|.�V��7�؛�8(́k��\<�/q
��G%�|6�Lw��k�>��-gRŢ�.g�*��Z�}t|0���ra8f.�X�E��Tc:Qw�LN�	_)��n����q̗�s�����/j���53�g	z,o�	��iV@��X��C��i��D+�ϑ�s��t{th�<���++3���� Ν���3)
y��5��r����7%��q�}Yٰr�qLm�.<���Q������AIã{�՗��f���S�z�5Y��[�d�Y�������U�Uo�E�����k������>��c�ΦQ�6o�͹K]0��ցyP��*0�ut�`T�N���E�Gx�G@����p����g>3]x�tU�I�,����3��1����휛fn�m��EH� �t:�uq���㑦+Ny����\��h�d��O�e��|��/r�f-v�{9��)l��B& �ۅ��=��|����crW\�O���V_6�u�5F�>R�;ۻ��R'9P����j�]��\;�>�t'3-WP�0�L뜻_ɒu��YN=i��}��4`[���P����+��T+�J�&�Kr6�b���m�r&�[�'W�{-?����!�r���%�4l6A��� X�5T���ko�ICү [!��ϴ(��ʤ"����q�/]сP�Ԣ/�����B&�L*1�'���oI�����[��gY����z(��ɔ��ó)�Ξ:���ԄM˔4�c�B�wǪ�&�8fi�͑�?�&R�͙�4l���"�;*��u�ҳ��I�N�36�V��w~v�>s֯��`�������.$R�>��9���f��!w6�h��˩-[���en̚M�5���)J1o7��rk��zJ��Z�N���k�o7z�*�Ƀ�C�o��>{�f��i��eB.V�=�LWc4�X�S�>�;�\��ysZ��;#)�!�:O
xq������#W��W�aq��%ݑ	�K�R�6�ݶ�*Zx�/8�ӒZ=W����b�d���8&kݶّ
K��ĭ#k_��v�������ى�<v0NH�\`���*���g֭��/e 3⺶���L�<�A(ӻy�rXK�g:�ij����.�_���e��u��}��mQ~*���겨�%Y���bf{�i�5-�jqPo]"y9�`
�+w�?(r�Ϟ�hz�Lmb����۲�L8�k.�+�i���t-GV�N�#pk�
͘��,���٣l���uaQ�w�eI=nx-\�V�VP���[��l�E����a��&���?T+Ž��gO�����n�,����{��nb�!~ܫ�Hp#}:�@��A��J�e��u-5OO,��,;Z��ͻk^��vB�ܸ����7�v|���R�3��u��>�����j���%�{2��c�i�u��R��/�]�;�����Fu;|zIc�h�Uͧ�e	���ϰ����I�K>]%�,����V�!�{nd��<%��45��/9f�)���z��f:$�3s�9���C��,|hg-nu��7���*�|�ָC�B}�m��E=�,�R��L�Zn&eO�B��]���o�Y�3�{MZ�յ��<��Y%�j�\�#o������O.Y	̇ ���P{J�.�9�k��[�n4�	R�����8�_�!����v\}Xt��+>��������Vh{:�-ڹ�$f��������Ք����ԧ������!F_��:��}�ЇX�`�(����8�E�'���J���Q.$�;s�TE�%����.}{}4�vyc��,V��yH\G�,6q�x��fz���n��=���sZ�iƕv���^�#��y`��:�t�7S�n}q��S̼.7���:��t51�i��Z�4E�v��kR��깒�}k�S�*Ĕ�Mc��0�	q�<��c�ۼL�i�`�%LgF���'�ZQ��!�֏92�S���QHӦC[���7�S��9$樘8�C���<�¢˹�G��nT������3�f��i��ilƋqn�1�g��9�kS�b� �O/�V�E���V�����DZ}��XQԥc Ųwd]��;�H޶��n����β�3ۼ�z�1��G�][�Ų�ߊ�زY�<�[��Ai�g�f���6��凯� �J1�9G���ؐΚ�ܗԛ��c9)��\W8�k����nK�^���ksj#��'�ے���o4��k�8Vx�Qh�Fl�Q����[�/����o��a����\����Hz�s�S�{���^,N�R��}BU
ظ_�L�ӹ�N��8��}�j��77V�/p�5���L6����E���Z}Z�%삅t8ż�_>^5O@��-NNվ2m`g�=9��ܷl{J��������r��[�+� ��bf��U�;U�T�P���jK�
�r��	CQ��ѷ�
�QXO3QZ=�D##��3OE9���|0k%�Ƒ�C�ae��`�
��^��bQ.�1PT�*Z��y��';�/��I�)V�eӵR�+\���+E
�,��dJo϶�s�I�8s8#F*��Zhb9�`C��0�PJ5�B��N�T�ՁJ��y�?\�����O	yF�����8z.�h��{g`�(�c{��U|���B���¾��K�3��0gWY{8��5}���ٝ:�kVC��\��W����l�ZL��U���'����Ӌ�Ģ_w�%�l#eq�!`�A��*ZTw�w�;9�n���nV[���]�ze��f�WiiG����)�D+��j�^`��{��Yà�.��9
�wV��N�]v���YI�ky��YYiZ�B5sԫ�
��fPΦ޲i�}�0칭�Z�eu�![r�i�j�n�E��vXٖ#Y/EÒ��+B�J�JdU�T��Y0ic��;:���O] ��g&3�Ө^�^Wp��<��<�eؚ�Ԓ� �7�d-���0x����w�����M�P�8%P�<_"
��!�	�����$�Q;}6�@�\��l^��+��涖��F5��P�ϩ�E\�p���`*�P!���f��ID��Z�����|�kI:�ċ������gH+�,E�UB
��~YK�ߪ�И�˽P�Ο�Jǚ�JD�[Lq�C��<�śt*�Ύj��f�L�eLo�%�ո��p��Rx�I����z��n�4�P�.��=z�Oj�%:�Ξŀ痆�Yb���޼}��}��-�Y&��̺}w�\����	��<���R��p�~T�'a!抱�]&k�N5cԱP�śx��oe��n��c*|�}f�R�B��hIwTqv����ɸ��9;Q&cz�T�p�Y;�Xf��èXfty�2������o�#�Y�D�&R�8@Oyt����'�$�!]�r��N�9���hWwEI����:]���uy����{�E��ە/sN�JT�h3ñL_\C�S�7�����ݗ���~�xa��R�������t(0�j�6�<����E��$�f�3B#��S4F�et�:�����$��ӭ���dR2 ����޵��/�K(�బ���!��4�/�.|K/��^�)�X�J��{2��m]Y0ۇ$�拽��Y�D�������p��nn��F�iw#���A��IZ3i��@���X�=�R�X���s�G]���֘��.���bfg �yZ����d]GK�e|�e_p�n1�ܕ��@����n�v�qe�w\w$}w�n�W�;1!|J�F��k�P�Z8R�;,����9RԬfNY�@1�tk�Tu�P�rq���ij�9$n�v\��B�Mgg)�Y�0s>e,��/�ɢ#}ܥ/�Jx���<Ɍ-��[9�r�#�����f�7��$��	�CXU�t�J �b�3SƅW�h�P:S�V���P���f��9�1�V+�bn�(�O`�)�ף�{ڭ���5���+���u�+T�B#5�L�E��؋��Q��۰�q�M`��n��C�.�|��|�ًh�(�tM��#jΠWf݇;�L8�+7#G��[z\�ȵ;峅��Kp�huhv�7�<���\����Y4Z�n��w����'�W�G�� �'�؆*
�&��|³����meː�L�Y ��!�~��>V~��T7&.��Ooͻ68�U�k��QWr��f�T7MZw҆��T�YM�!�=.+����<bp�3қ(�	��[ D�$��U��m��j�)es�������gff,P��4�bv<)$������ik���<�i���viEm�hr�zv�x�E�zu5vk81�z�F"�7�%���G^P��U���i��J�����j�V�ѵOsw��L��L��2�ƛk��չB�vV_]�\�f��yý�<y1nW���p*֤�ѣ&��c���˻!Ӕ�\εǳ'k���[���3a���L�i�4m��ӋB¤�-�r�,����E4 v҃9N��}m�5+��P�]��q�n���z�H�:���T�#�Ԧt�{U0�O��xW=�Ol%6ӕ�ML����W�PEF<v�����f��;B���/[7;k��]����֫�t�3����և� X�� z�nҮt�%-�)k�y�T�AZ�`	3�і5h�ns\Bέ�wb�=��� �Jz��v��l;u.�-oa�*�A�9�Y�Q"�.Մ�f�E�ҭ,U3�.�t��0EG'��:ޞ�T�
�4\��� ܹiS���+��)���kx�2���M���ut�-(,±�m���YcE1w�Z.R�gsh��WpE�|�\ТZ;1<���1���a�_JT�%]RC�
�F���Q��a�1HDfaY�e��YdFLdU��6I�4�Q�E4�YFN�e�UM��Y��LQ�fD�E%QM�afa�&A�UQUdeLQ�cT9&E9�D�d�QTdd�d�VV4T�VfRY�R�TDI0Y�dd�IFY�e���Ya9ee�TTQE�fUfe4MQ�feSU6Ba���T�ba��Q�AU4PdY�Ye15Vf�dMVa�fT��E$A�e�fb�5AUSUDITDEe���Ue��N��Y&a�T�.FM.e�QUe��UD��T��bE�1QQ4�Q�aPRMPLED�PfFXYf8dQ�Y���TM3͘dMSLV`�U�c�PFXFF4@QFfD��e�5�f�eQ��IRE��QK�uy��}����ﺯڹ�� �s���h���ah�B޺�_�O�La��p����os���]ޛ����#{�a,,�؝�7B��U��(�i@�P��Dj5�uQ����R���a�x����F=:C�5u���M��-��M�Αf	�W%�4l$�o���Kz�%�MY��Ӯ�9�FЧ��w%#�#7Pn��E'<��g��t`T<u(�,;�W	�ՙ�w;nT�������1%K�:}���uϔ}L��e9�0�Ot�W�{fB�R7�r��Z6���>]њ�h�s *:N��͛�7�uc{ŇG�_���D��7�I�[���������M�|�@�m�sic�h�g�q�uB3L��t����Ŏ�[�};\��R�ڔ�hq��TRL��G���oÃ���^")}9XI�Ox�]%��K�#36�'`��P�!�@m��	�kҴ���<6�_���x� ��($��R�a릻�۾�
|�b�vp9>X���tD�0���%�o�����������[S#��5��m,���ٽ���S6Γ�+w�?(r�,�5�_ɍ����)�������r�յ����>�َ���RA���1�`I376��j
U���d��T[J<b,A��'8>��#n
��>���d[§[���j������]��tyXn��ys�i݇5:>u�-�yնj�w�j�E��yZ]u�erKdY��/�|=Zd�3~�r3f�mH��|9kN�S�٣ok4@��Y�{zt��'fZ�!�̫�|�uf�}R#�z����]�ƪ��j���[�Ɲ�*�����l���z<gڶUx��y[B+Ҹk�\=|e�똡��X�-M����)=m�f9�5��OQ���[��v}��*����h��߫�
ܢW����>�[	�#2�'�׺����9��h_g_��5��{L�YΙb��̠��+�Qq��poQ%Y�r�T�3e�جvǖp�>Xf��#5��Mʊ�R��̠�`�V�	��ٶ�jr�_s��45��u��;)d�AJ�z/����!��!�٘��ҥ.^xB�*J����(\�vF�LN�\�q3�,QS�w�Pk�y�^w��w*��m��=)��/�yF��;�X �/�I��
��CᎽ�W��3�μ�����X��D����0T@�*���F{]�8M6 ���kA��i�>n��%��Rt�k�/�X�Ϝ�����"�q<뢯�s� �:��-2\���D�w� �ط���G<6���!�yt
J�>)źqa�2ս�َ�7�S9�2�fb1��������T���g����E�6n����L���=8�f���콞�F%*���+5��/�M�sm:��U�ѰdA�ϩB�uG���v��mJ�w�5G���[�<2���B��NB=	�5��ũʒ]���(!�r�x?Ns��O�e��V-��^F�t�����$��)�'!&㜍4��k�����`����w��b܉��R
I��)�V�2̣��:jv�T��J�w��:�'js��*r�dl�[K[[=��Q��@�C8,dD�,FIh�l�Q{8�@�����j7L�VP|�u>�}��[-q��S�0֞��2Q��UK�`���ukG:Z��',�='͎wW����$0����V�U]�Ϲ�5�{D�K1[ ��d�:,�,��S�w.}n`*7Ryf�I���K���ha�ON@h��=n��ߥe�Se���͵��qV2Y9�#"�Ջ�Q���4�ř 4xk�#^����r��!�5�qJ�
*�QZvT��&����"���s^T�~��:�y+��xPT��C���z%�N5yO�g��Z�Tj�T�z4q|�N@�D߻X�IW��8v {�y�:��߻'�^�[�m���pb��WE���(�&ֹ���<��<�<f���J�k�o�B�>���{�����!�M���HU!��yX�'ei���F>{&Vͨ4\�;0*ʙ��<���ijԶr���:AaIrP^�(��9B2�PU6�P�V�d0.��P�׻�.���Iq˷-t�p����	@�	s[���N�}R�V+��w�5�Y�M��	U��X�8������'�V��`m� �2i�[���v��`�gZ���J
��<k�Ď�-��>��sS�M�p�����Q�kI�p�EЮ�x:�;s�3X��e;��2��r:�X��h�%LLo�,F�^��,�K~B�J�E���4\}��#���ٝ��?U ���X�^�����wΔH�6:T�YwڒX�U�*�F�U1y�����$T��*XڙB2,�.ac �^̆�&n"zğ9DG_^�տff���씮3Lٍ�Y(�uL`���K1�e^>�C��z[�;[�]��S�����55�"\'@D��ċ�a���0����z躢ɮ�H-Y�6/Y���n��'�4%,��\�:���x�����x^śt+�������T7����$^���۰����v�e����lYu��B���9��J�K�^�BA�\a��f�v՘����a�R���D����yL���?p��l-�͑��c���P��8�*�ݚ��;ښ���\�kl��w�l7�5�I���8MK,}�kC9}�y!b�{�O��W��J�u������&:���^u�xC��)s�<�M����m��� ��Vgy:�ʮ3!s��=�+NC�\:U�vtFUr�JR�v����I��e^S�����/.#�'����u��6>��Y�PU�'~y���.n1^;x�`�X�4Uf����9x��PŵbKË��5����ŗ�]���'FZ�K:_)c�EV��� "��S����\MF)a�m0ǀ�-3o.���۽US=A���"�G�V���p�\SF�P�` �=a:A����B���g5�{͉fh�=&z�M}�e�d_J�x�����-se�!>ð�G����\�Y�$s�rtlC=�%����C9G�̴�P���y�(�p�ԄJm�]Pۍ�t�j��(]hmH�1(u\�
���6�;�>{�)�^��2�>�P����R����LG\�� 
����u�~���ג�[�[J4!o�Uqi��Uq
j.$Ti�v[Zl�W�tӌ�&72b�o:��$WZ��Y[k����:,UupY��o We�i�o]Jos �5�[��(^L�����On W>��wp��ެ���� ���W,K�̘��:����OpG�=R��f�6b)ʝ&۵���;?r�<�/��>�S~�1�K�E(��m6dL����:��8���'�g5�G(z�iv=�gб�+�0״�g��ٳ�Eu���ۘ(���������T_�5�A�.v�1A;�v��yw"�<1��&���f�E0lXkPM:�}�n妮�����=��Nj��Q|��p��<J0c���jt�����,��]�j�:2z��hu�<u�*tMl�/�F�a��y��1~ǎ������@����]�v��5�{�;fa݌��0���751�%U�l����T/<�C��S]#�u;1=��0{9k���1���T�����F5N�*��u
4�ϨO�W���J�e��mu�D��R�c���U��P{�瓹P�u�h��'�f����)Pd.
,j,��ȣ/�N��%�Z��>��Tؐ�.�/�:Z_��N��r"���>�^9ix<2�%�ҚB�F˦K�_Al�ۣ�Z.��j�S�����|z'�2��њ��tܨ������C����=F��sI��So��q@�F��՛���/�|�g֩���@k�\J��pc�G����]���Q�62+�2��j������2��Q� k	��������u:.�e<|�Y��k֦:��-3�P�2I�r�V}8���\�)>[�,��m���t4��o�X��+������\��@.��諨�z������Z��z�L욀�rX���r����b���;��H;�9�bE;��Fl<�f���A��Ņq}=���}Mm]]eIy �O\LJ�Q,W��t�s�ێ�C;�4r|�C:��,-���|��3Kج\�	�i$W�%�)ko�c��T>��Y�E��Ö��u���kl�g�Y|։Yb!�^a0��H�2(�$1�S!캅1�����j��e~����ĵUA%UU��y��p��z.�4W��,\)ʒ]�"�z��
}�	��st�WC<��J�R�j���D�}J�۪����4�<7[ۢ�b�\���5���S�����ϯ1Y��A�,�9�j5; ױS ED't��9gkb��B��6�������R�K谱4�xGZ< �E��͚
/g�3���E3���L�֒����=]�w�ʲߔ��]�oPf�V|�p�N��U��;Z:/I]s�)��u2�����廆��:�xYjn������j�+���]����]�^qG�b>gV��Z�݂�6i'�ђ��v^b9O�^wWNl82T�B�Aە<q9-%l,��֜��N��}Fo����s/�O3D�ͼ�ז�������c[��m3x�YZ��p��]�7�������]�LFʛ�S��=��S�#��RV0�Sԩ=U�'�u�3���ok%����m�}K��K}':����[�=��Yx.!=wC�6x=1yp:�%:^e�^�`;0�x4��k�V�V9SӐ�J�6pgE*��TV��S��o�-<�fG92��WP�D��S�AR��>S�D���hLj�ZT�m�^�:��<bC99%@�_�3�]K���\�k�Q�XMμ�?7�zM����\��nY�u��E�ޙ�fD8y��B��]Eʳ��������UG.��
y���VL�X�VN��y�j������e�&���Р��P�c��V#&w{k1�cy���J��5�E��8[�sS�M�p���Q5��t�ʮ#d��×�3Tr�vfN����Qq!E�l�ٯia�N*u����m˳ю�X*��&P����U
�=o]�m-�Mȉq2�W�^�Gf*#���B��:Q#��ST���=o�+K��C�7���
��j�B�NC3+=��C��g�g��(���#�ǆ�j�f�]���V�Q�|Ob�Ŷ��ר�x���4�{�
}u�DLMp��A���('����Y5.�]�u��TV��L�n�M��R[=����S�˷�� 7嗜��;%�7 Vx]���UK��S���^N% +Lb���i��f��z���@c�jʸ�gjp�@g�.P�ʦ0U��y9e�cA͕ ���pR;i��ᵱU=&�w��:�6g�QsV،�����U��%p�m��Y��K����'�2�Q�\qp0n�d�=�8䱃�<����0�V���	���8�&Dκ�h�9:�sMi�ʪ��
+&.+�3�z��X��j�k�L�i��40�:�����h�{�k�3�Ncջ~7�J��mx�M�L�}V3y̍h�	��!������0ᶄ��Rm,����5di�������u"'yH�F�1��,)���/Tʽ���MX�Y�'��q�0B���E��sq� F��k�U(-N����0����ꃘb�|�%�f���U��F�q�e�zQ���W���f���+�vW[&�Kl.�][]����,���o.�8$��`����'Z<lOb�q.)�`�Y����H6ԅ{��5^n��"�@���Q��	��V�i�X+��Z���N���(�,&���a�F�i����$dȬU(���x����oۛ�,-�DL!�O�jtRfBbybU�<�T��XM�F0P��g@��סP��*�ݯ�Zy����+&�E-8�W|;��)"�Q~'x�9�Xyʨt;��~N�,/����
x�QXd+��T:�}j�}�G����X��1�&�	�vl纥e��y�Ō��)�L.������U��՚[�Oy%-O�.-�T�a����+n���)�^���ϦT#���+GU�[[���L�Q��D�~��il��up�^K�un�m(Ѕ�ʮ-9{�w޳���'u�Y]5�C���:���d:u��}���q��?	W��T{�(���[�5���z��M+ ��%g��w�σ�O�)��9�K��'�����Q���X��_�b��X�|�7�U�����,+nd>�,r�=B�A��J0�xm�ӥuf��P�s����a������Tӂ'ٮ*E�M�8����:�^���U#�l���s��������.N���Bb�i��xS"����2"����1��n��s����B�J2P�z;"����5,��:����N��
2j"��W�A@��l��A��硪���Qd���IVRa��}W���#!�� !B����*]ee0�WP�,�@�M����yʆ��Zﱂ�C,���v�M�J�h;�.>|M�t�oNYM��^;�Gy�#Wݶܦ�:3M�-V��Ʋ����al��2@�&����u٥Bg*Բ�#�eIF�ų��W��T7x#�0p'c��#�O�V�0�{�$�������Z�2{���Z@ד�6�;���4*)<,>�� �at0f����X=S`ީk��W����LW��󬬙n��][ʎ[��E�`�֑nɤ��M�3�զ�#Q�<]L�ڞ�h���Y7f}%5C1[|+�t�3Xs���۶l�hF6�G`���C�>�~��xΔG!��Me�^�����H1,��Z�Y!U�6���Pv�I����+z$<cѝ�c�����@�ӲPZ��%��"�Yǔ���g��V��I@�Ք҉m-)2��%U�c�
sG�I����:��b���z�
i�
�#RT!���gu�K4Qt̬	���;[[7x�<���s�sYZN1���!����U��{���lW�h�0���\<>+�#����@,�Ξ~�d�`�����=���.��l+^4�Q�۵�&+����ܫov�t��ך�)�u�-�xo1ďm_%V�e�Ӧ�)�ю�
�G��SW�V]�$��QF)�= C�O>"ݪ�����n�s.�f$�5��Pׇ��;�w�y:r������BT�Ń��A� ��M�I��N��,�xmv��'��ޚ>śI����TW�x��<�yF�sF���L��z�s2�YK��i�wZ���نBE�GR��M��I�2��+y��ݧNK��>p�7N��F����{I��򸌡I�h�Q��n�޷K��LǊh�)-[\��:��K^ڙ6Ry)݊��,�"�ɩ��SU̳�O�u�.�aw:�:����r"����1>�9�Ax�U��¤]aAX=�N:���SDM���s��w��>쒮j[���S�e�ÛZ�B�Y��k�$�P��)B{`���e�v����9ݞРWB����HR���ҭ�Y�ꖬ�f���%��p��`��e�������=���V�d���*�I�ג�ƨ�%H�A؝�`�ۣM��ہ�m�J����lg�S�!F�����,�㺂$�dW����4�ܨ���m�ft�l�X�z;�Ý���r��ɮ��Q�h�NqW�v�����뮥�YgB(���,.�;̚�1P���y�x毂HF;���h]Q�'y+��;����I��l�Ss	}]�7��i'��̗�ܷH���j\d��^U'y��1��TP�%�u��(�;Q0�_����S���9h�y�ă�>n�������7�m�Q��(l������e�|�H=I�|�p3q�Ⱦ��N��
����/ᒟ$+����
����0�2L���2"�(�����rZ�̓2�bH���h������&�X�d�(�02�)ʲ"����2"��ƫ0
\�j31��0ʦ�(&�̱"�j��"�,J�h(,�3(�1�
)�����
�Ʃ
(',*�32���H���0�(h�(�
��,������2�#2�"s&h�*���r$��i�#3��0ʨ�p��)�Ĭrq��,0̌�*�J�*��+3 ����31 ��2h���j��2ʪ��ƪ*�1��Ȭ̱̊���,���ɢ�(�(�,�+	̓
�")�Ji�Ȝ3
)��!��ʊ*!�h��3*���H�,
,�3,̢�(���lpl�,���2*j���(�2,���
��)̳**����'3�3
22��b��0��3(�ʫ3"r2�+̈�0Ċ��,�Ȫbb�����̘�2�32 ��-k����˿9�(�ٽ��7Bˌ�k���ڞ�ܮ�2D�R�o!�P�k���4O;��u'B󕲳p�>r���Y�9[�sZz<�{Ƚ�Y�L�g�-�U���C�
�/�ϵ��_�ג�{[�@�������vp�}*��j��߲\<�n2l���T�<�A�b�W��	�S�P��.�`m�Gj�Z�	������g\'lk9�{L\�Y܉�+I%1�q�4�j�f5ܣ"�F��eX"E5f��}����O�Fi��p�i��7:��ew0�����Z�Ǻ�M5 ��>�wf`��������f�9��yAt<7���El&��{�I41�`?^ʒ�\(m�JR�L�6��/hw|dO��/gf�ۨNT�N�$��+��s��=qP������Em$y�Aq��P�u�,
W��7�Gю��z��k�3g���q�V�j�6����a�"�Hy*�^��^z��%��'N��Zy�(����u&�i��G���OlYq��U�0J���uj�lȃՔ�~��\]e������A%�.�6��R��t��b�ٙ�]0��r���(�cK'��Yj�ۤ�j��to�5�dI${t���Ȁg��>�|uɦ�f��oX�E;|z·�r�}�Z��xJeZOi�a\��1�jv�;tRw�M{۲�����R����_�+|z诊A7��>��C7���;�����mGAnG�p�:Q��|�χ-�(���6����|�h�"�fXཹ-�,�?,oح� &k���Á�	�GI�F���BQ59�ў��R�v��i����(��$<7��r�p��v�8J���eU�`/;�� EBwKAh�����ݐwi%���f��Η��Ȱ�+��x؂��ZS���U�����5�&��yY��t�|N�-C�����<�VY��0���'F�ͦ*�B���b��ާ5w>�9ؤn�S�2��	r�Y��%E�LSU���
��e��ρ�4��v%Y��=J�{���J�v.�~�2��C�{7>�f'��u�Ӑ,-�[�=�]X_w���O%��C�)i�T#3��n�;`���	�hã�g|Z=���r��!�5�qJ��f
�q�O���$�bG���\J�Aඝ ��-*1L,8J��' ��0��2<����|4�T۬�9��t&�Nل+�K��Y+�ܙ�*](��(F\d��m�j�t��{$1�x���]v��So��uƻ�͘P7Į8`T��٣�糐#��t���'��[f^�XLY�F-���.�7x����W68gYd�2��w\��L�z��5��G.,u�
+��g+�-��i2�<��%r��}�.�x��{%Z���3y}�ѭgrWP��stJ���Sָ�*>�Nv�{"���T��Nts������:��q���l��%iE��l���$�^�AV���W)m}t*,�|��z$�X/�����N�����j{2��K�|p�_<�M,���S�ξ`�����s�8�YQ�\]��Qs�f��[ӞT�5dz,��T�Ɖ�#X�	[t�OVWu�莜ٙ�}���B'�
O�c,`U(��#��ac��p7���*��͋���Y}�n��YJ��RQ�NԒ� �%�]T�M�ǆab��o1;�<)�(>�޴6;z�&�;/��x �))������ᇐ����\����0T]�!^���𱠴ҹ��@|����&ʱl�mߪ�ic�H��g�Q�<��i�:�P��T"�׷p����i�4u�ueӭV�\��Cb�`���q,=|ZP����L�`.L���2P�&�(ht��$��6������0��9v7��I�s��9S��׫����T{�4ֈ_^�X��͚4�ԅE��F�x*��W���9�+M7:5;������C�T�M�� ݺ�"�/l'�Wv���M�V�.�{�x�+���N�5u�3-����%��SO���d��c������G8gY�<e%N���v���YN�l:g-rv`A�(s�7\eJ��.ĭ�͌x�EZ���c�U�=t�C?gl��s�yU���Kd߶P��j��Of'#MΧ^ӥ��g�ܬ[��������Mƌ�t��@�QjY5�R�7��;k+�����=����qY��ċ��C	z�=K�l���( !�+8�~n�.zM>���9��>{hWKR�͊�\�<]t1Ƚx�j�A�c`��pWY�Af���Z��#���7K���9��X��������p�pX_i�����Ԣe�˹�p��ĩB�U�p���'բ�Z�x��:\a�:�e9�0�O��P��a�G1.�ME�8��w�R%0�cz� SS�ࠃ͛�7�ucCN��6�\���l��ќ��D?At�]_t$ӭ�/��/.���k���00�9%�L1���~���x�Z��Vk2���ΐ8!�Ϊ�1p���l�Ӟ��꺦����3I�Z�Ĩ{�f;�Z�n��&�˾�̋f��Iĭ"ÖO�LVa��K��'�����h��D;��0V�W��Ð���j�S���(�lA�G������<߰��Q�[���X9�HIw�1r��yu��Hu�����2wS��r
�Gky�(��;�҂��.y�2�B��R����e �-v���/OpC&�[��ګ3��6���[M�;�,߾�����	*͂¶�@pE���0�o�w-U�
W�P`!����t�����v����_���{ׁ���p.4�����1�D�t�������הiw���.A<��Sj{vze~����As�w=R���2��,����UB3:[-�y���q�z�J�Fޞ՞�r�n'���=~:Ai/q���:���["�Pe:�x�\�xcU-o(��J��<��uᒼ[�#����x�چ5O�ʬ�]B�yu�\<P�L'/��kn�8e)�zv�*b��j���,�u�h��'�f��T�<��B��6���=��k�u����)�&�Y�6
},_�t���>θN��r����t�'͉3T��� 1�Qi�r�g5�I�N�DmDΠk�9�G�>����oτ������J4�6��lV�/4��컛�}ݏ"�@��I/�����Px������y��=����à���n�B0h\����T���t��r'I��>�B��]J$Ȳ�S��U�w�p���¥����èGИC�R�fn�p��c��s�ō�����K�[!>��S;oR�⺅T�+���,vQ[,�2#����oޒ�=1�3�ӄ��|��Q�8�F���Ņ�N\����:gVM�(��.��\<q�n8�qڕ�`=kOwZ㝣�~ЇX�`�(<�m,��5��JǍ�C��g<���T�4���g�'U��L�ȡ�+ɷ�0u��E<�L�=��n�K�����,�p*^t53��.=]���2[�ᡒ���n�􂬱�P��%�uj�lȃԌ/o:.O�׽[�=�3�[��6e穀j!O{���.�#��p#��N��L�-NT��mW�O9-����"~����ʇg1ͅ�rI��qPR�p#����),����j��7�Sݲ���qDe�K��qW�xp���:jv�,�73���\�W])ȍ/Vuħ�8hj f��%�[>�*�X`���6�V�q���F�>�$o7d\F,��9	Ύ��t��=��>�7�~1U��
T�z��iA�Ҫ���T�SL�S�עz��̲U�LFʛ�S��p֣qW�t'b ��(A�o�k��T+�V��q�7>�O*�2�za��b�vǶ�V^O]��Kڎ=�#$��8:�+[�QړUf6r�
��HWc�*�mS3�%��<���۹�\b���w����۴�w��#Bi*�kͧC=��7ך�:ο����V��l��0����M��I��[�h!B���ָQ��|
�sC19[�S+tU��o�Mjﷻzwai�V�5��� A�����IZa\T��>���:7B���T�e&v��>�n1F/e���c�L�WN�Ur�#�gc

���C�a�^�.[ւ��2�uZ�P1��ن*
�%@�W �[.�.Q5��n�=�"�F%B�I�^��2{�gE��=�N޺�7�J��Ceg�4)��l%�j>�[��*Wj�,_21Ӷ�v�OT+w����UX�~wHdXQg:��D�q{hPq9k������^V*��FD��q�[�"��yM1�$����j{2���_��(�%�K.t�{B<�.�ݛ��x����!�|*\����ΞT�5g����n]�4	�#Y/E��__�v�Olv�t��u�X�F��\�R'�,�c\^8����J�������<ñ�:�*�V��T�44<�MW�Y����\*�vxAv|U� �~�	%��u=�
U޵6z�'ᗐ]�J� h�i��5�Ny�D�7�r�nU1��w0�E��}�ۃ����WelIam�N�,X�����3�I�&�xha9�+u&�u���A�n�Z�Sm�V$�m�OG��,�YK!���VK�LNn.�C07Mٜ�\��7sR�'m�zWdlR�T�F��]"�3�K��₼�d��2�+�'���e]w��΀,�JZ�X3Wy,Y#e��s�� �q�JMWپ�FF��������A�r�<9Gb�c�*
��L�y(i,X���!�mЮrs�	Ԑ��cB�5��ܜ�u��Z�z���806�r�s.7#e�M�,n��[\/��N�չ�YZ��K������9Z{��xu��q���LZ2�،����騾�I��)���cVq�ߧ�`.�팻7�N� �*x�P+�d�-�{(@��n�
�h��u��&{%��yByˎU���n��Ƭi�6�"����,�(�r�&��b������C�vu�5=���>��/T�R�<��CR4�\�`5�U}�z )7\v�ܞ}�BOV���x�psq��U�ev�o˨�h� @� !�moR�Ը\���y���<n$G��|��SV�T7���g�l�����Zm_��@���E�zD����OR�ܚ"���b&��,!�%��C��1G��	����~�a:<¼�~����(�o��Y�)́d�X)f:���&�:��k�T��~��Rm_�C�c�u��VҜ��`�<��h�J;N���4��+�9���e��6���/e��m�����
�ŉ�k*L��66�l��71Pօ�4�Z�P�N��um6ȫ��N���dT�5�@r��&ê=x��<���<o^�t�3�����o&3Ƀ �h ���1$/�_%�+��|߆��������V��-�ԥSL��'�qs̰ˍU�ӿH*�8�����b����̬=�-��SV^��-]b���֤gM�x��pW�����g����G>Y>�1Y�:�b���<6�)�y&Aޛ����k�˜%�{(f�����@pE���|��Q�.�\�05�y��&�s�R[�x�i��x��h��ᚶ����C})�szx��W����v%�_	`R�9���ܞ���|��cH��chv(�B��/T�E�g�j�F^u6(��8���&F�)�7��9u�3�,.�F�ӂ}�Ǭ�/��L1��~�4��2�{�L\<���KQ!���^{ܓ���xz>�<��s�xd��G��k����1PT��P �N�PKk%�r�X�r�Qj�:��vX��,w�T��ۦdS܍㚱�� ƈ�{*���-�����S�t�,e];<�Ő�E�SʔR�fLP�wZ.�n6����MX��D�]��Ɠ��E�l[�� |s���4e�&0`0#���[2������ T�q����WI����xa�uN�K�|���œ��#'�MÜ�l����W�,�5e2�� ��X	���^�N��r��[�gqj��7g'Vc֗SZ)�U\^�"X���!�ڴ�&;c�8<���<4E���f����8�\��ڼ:��=SE�ꐢ�I%*d%3f*
�y9�)W��W
�� ����& �t�3��m]/��Dv:�;���	GˆJT�y�\ϢZ*G�Ê�n��ǁ*�B����>Ovu2�c�Xr޼ӰM�ŀ�u�Ar����;~��z.Q,W��t�E�l*۠������>�8/\#Lp�X�5p����p�r-$�y.�X)s^�c��D�X�vP��jΫZ�E��'�:4q<p��.5�AVX�C��	�:�Z6dA��X8�]��}�g�z�m��>�ڎܖzq�ٙ�],G_��p!�N��L�1GB����R�����'E@���5���]��<�^yo=J�BU'!$/xU]ڻ�qX��ݙ��nD%q�l�҈�3���s�\"�t�fY�s�֧`�b���Xc����ê�9si�n��ٳ\9j�ƕ���b�
Ղ���$�ZۇV���V-��:,]ˋ��ٮeGkDf��{^� �B�����#}o�f�R�v��n�v�u(����خ9�j���D�Ǚy4Z4@=���U��h�[��1��f㩕hM)�U�-me��]���,�I��.�C��](�ո�`�@��La�kC��*��Z�g����j����N��(�
�q4�Ѷ���w��6����hR�d�k}.0
�xt��ʚ�
6Y��~x�6SwSe�u��X���K���@�+��ݔ�WL�fp,uY7C��4u��av��+2��W��Cz�5Ħ���$����e����?-Y��(̋`��x��E�8����WdA�9)ѧ���:���~޸n���u�^�E�ZޔR���H��G�6�,I��v�!�kF�j��ԴM�r�r;��M'�8�C�Ml�[�_`�U�)����z�J����9��to*�	�y�ڛ-���5�-�� ��k��I�6�����ץ�l:M��̗p�p,YYyf�T�;�D;Z)����*+Ü�6�@R��Uuz��c�˽�*z#���$R��^n�W�#=f����a�����\���s@��0���Ad�t���X;˵�9�'ox��wnbge��(�|�Z}]��Տ9��ۥ�]���@{�?t�5uփr�8�!�(l԰N��w�],Ksa�)ӾYl�KV=
�P�5X/�f5Fy�^�J��f�\{:HI[ӘJ�}P�*���~����t�4X�us�̤�;¬ZX��;Is7�G����
��t�}i�~�vt9�i�B���C��PdR�8>��]�.һ >9)dE�[ɧ���i�[��d�XH��7W���od�����X�*k��k9㫑�T�������M)@.gnV�Ԕ�ر!��u돹@y��[u�s7��	�S��XD�*B_m�v��+LRyӍ����l��ϝ�@�R`�����l.��6
�<,�B�k��[����D�V�$kX��3��Ͳ���SuoN,�˖�*N���!��M����;�5kB��il��9�0q��RPm�HA�-�7SM:�\{o�ݗa^�wfu��`��ck�Qت�ᚖ��J�7�[v�B�}�ɏ�����t���^ �wϑ���66
<��{)p�er.��z%
������R��7�{d���o=��9|���b��h��Z�Ú�b@]�#s��6��So��V�l@i��X6�Q��v�s��`�^�޹7>/���ʖ�д㕥�H�8@�:�����9�(ܹ�N��B͝8��vH`�+t��])�&>׵�;]*�d��ڸ�Xgd�\�	)oZ;xSP�Wy=�T��OR{�k��ۘy��v/:���Qt�Ht�C���i��aPD�E�Ue�fc0�,�B�EE!�UD�QT�QQC�a��T�CTda5LfM%-TՑ�fffSQCESDEU4UTe�IVeUYAEQAD�EQ3QU1E4DLT�QVFET�EefE4YME�U0NNU3PY�,1f55ad�e�METSEPDQSTU1DDAQLe�Va�LT�U�3TUU4L1C6SUIMSU�Pf%Y�LUY�4Uf9QAFF�EE4fbTř�U4�TM1L��Q1VFAa��3Y�EE1UX��a���55%1�CQPQ3f5�dd��@fdE6fL��ANNe��eLKQ�c�fbdd�bASKETMQM�dTE��4�U�eDUI1EI�a5T���M4QN`aSAA%EQ5�d��	RDvx9���+7��۟xP0�}]��O����W��a*v�w�.y�i�f�.�d��+��QJ�a��ۋ{��;�H�b�ɷw_�ëAƤq�}Q;	�Κzv�/�U����'�}\�ԣ\w�j��3�%�h����ݑx�t�':;�+��uJs��j�b��>��B��l��n�Y&�y`�Gyp���N��!��[T�l���u>�����G�����n�wQ���zv��<˳��*��1lQe|�P�ٜO�M\�nD[�=��Yx"�4k��=�.�+Z�+�U�q,W�b�\X",�H�d���T��>����t.�P��6 �͞|$8^���u�w�9�Q*hq��t������,oD��#}�OOM����gF[�>�5�u�И�~�va���IP,��nL�WR�YD���էf0�*�p�mfB�$�f���p�ݾY�@��L��k�0��o乭�_�n�ν�o�>���᪂���S(�9:.�<��иw�ؼ�B��#�F+c� h�^��$=a?`ܙ������6���c�,R���P�I��%����M�p�����3J'ҡ�\=X"�t�=�Ջ�<l�;8�Y{��	+i�9fJ��F�9��d�[�;��ZB�pn�7�3���~j�x�g�-;&���W��r	��S$=�9��p��ۄɒ�N�t��2���Ͻ�ח��3l�N��W��b5�5;y��/�1�,t��{^"���*\�$��h�����u����K`��=���&�]S�[D�<�].Z)?�.�,X��*u|�yJgî!� '����B�ϖ]$�#Zt�)�?M�C�v��-H������Rbp��0���m�G�r#{'s���M�*f��|���
�M�D��o߹y�5��Y�˅��߅�"���YMtFvl�����ݓB�P���ʱ{5���ZM�"}���E�ӷ��6K4��}sU�;�蕝���Iⳤ�3:r���(�~�l���ׅ�<��#��x��<�����{8�$�4�����7��
��ys��͖5mS�}kk�d���aUƧ�;>�߹37�<��{D%���ʜ���k��Ύkyʾr琚P�\��V)���f�g�_'��=o�`��tV	WGȹ�..���x�x��o�(AA�=S�)�y�]ڬ�c�&n-�l���S�;�0�l��#b
�R�X�G*�қ�N^%p\�w[Ւ������8���uu:9���ǹ���Y��
4�[	���M�2�G+�ұ���r�;t-�7y����4�&qޛ�"u��)V�P���]<7�y�z��N^��mhX�P��5}Z~zĔN�{��g���-�Z&�y7�*�UV���Y�T��(�ա�u��Z�yҡ�c�U`!�����J��n� o�~�~�t�������kvS6�F�W�.���#p�O"��yFPd�x��UҊu�RO5#)�>��U�$B��0�"Uv�W�5�75�YϦ;d^t�{V�ھ)^��z�WWW��Ӆ�s��w�R����B2+�¯ד^%͜�|�G;�y1`�	�Ys��*{4n�%���[
�^�A�����^\2U*^�*�SXM�y��P��HvD�k��nu.���L���$�Enn*�{d���ir����c�'IB��;�LesGVw�\�y0�`�63ܢk���N��1jp��l���Z=S,!� �Y��gw�7�[Y��+�۲DLZ�5�m��h8	�XF�:h�4D�0�����n�[{kC�n�J�qST%d��ê.���{(f�	*�,+̀�Xx�`s �Z��Gk=7}J�y-���!�xՏ\O2��/�_�ǣ�f�WYI�a^>ȗE�y!�{c��su�Ɵ
U���(��N��]�^��~��M��,F����_Kb�+Y�T75J�OK�L�x�ќ�r�Ox(׺;%+W��а�,�L.���aㇻ���l�x%vJX7R�:�֌	b����w�vpZ,��R
nh�|�kuG9�wK܅�ÝÈ���/���1A�^��s�vJ�٦^B�ȿl�t��Ҭ���M�io��`��]��8��v�F��^OQ�шN�H���M��n��x]�be�n�f��Ј�A�G*�OM.wg$v'�͝s�{%x��G��k]W�j>�������8�Q��e���{��Cb��/�ǔ��Z��9u-5OOm�avS܍޹����<�p��;r��S��b�?M�ć��c�G�2�b�},�a�>���f^K
ªR�䁱��ǩ���l����Ip�T��.�]
��c��_�1a3��>�DWg
ܫ����]�a �n�!׷R�-ԇM��T�[3[?�-��úf�|R��#�w�"~�-��;y���Y�����]�z)'�/(i��عT]���^*zΊwg��)Ө��qڪ˥u�+N��o|w�o�`3Bl�A�V��\װLJ��ƕ��;��S��)V���\�[�4�vB4��X�5o)�Up	���+g��r��8£�qK�̻������8<��q��m_J�X������'GIWI䅽�_d�<w�^]k5�S\�ܽ\�<�����D�,i��a.N���U�uܳ�G�`�m�&s�¶���uG�O�幹��7����g=��V�#��[����3Ӓ�4z�����|�s3֮*��$e��J�U�0��H�o��M�{�Y{��Z�ZZ�ىEĞjo�x;��	�'O�=UV9�!��wΔy8�N�і!j�MV^�8��#��&�'gEA\1�mh�2WKY�V/<�3�*BU��r	>K��J�l�IMP�Ĵ�i���E�8|d��Q�J�EN߇	Wi�ʿ,EoI�{/c�~L;��/�;�H�u�S��p�ׁJ�dXX�Ô|�X���ճ�'N�y��I�R�)�Y�.��"�-�Cup�^/��pzy��K]0�c6q�k
�r�h�n����Z�*�2]�p���i��KXtJ�N�C[ڭ���e�s�kC�+D��<V����>��O��Ĭc-��[�%�Gg��u�Ӟ�c�*A=�.����togK1=�h;�=Y��6�����X���a�jJ�
9K��3W�I�nD�[b��,&tl��4��Ei�SC�L�r��r�"���xP[�"�U/�������~�Cd�H���\S�P��in�g��0�N��h5�^أü��H�w_s;�Z���+�a!t�B�_m����S�JY�@]L���/w�Z;fLxvY�Ȓ�FW�8:u���ܲI�y�:��X�j��郞�.!����O�f)��z%�Ny�1��]�b��%@�W�3�\T�(Q0���`B��;��i;E4"��J�P�[���}�#����
 ����'�޾W;�S�s����*��`�G�L�t>����+��]1i�!v�1P�3ݎ� (@�saɯ#�ßXei^��x��Ｌ�C;<���~mTp�]Oc�b�u�H:(_ͿC����S�^���Ƹ����>crبUs�f����:�Y�n�Ce�؞Tkw�[I����3���ӳq8?+��K����%�Ţ���c�ōqx�|�yO����,��x���~����UM� }D�s�yJ˱=��뤡΢�̪^Z1ϛ�J�vxO���1�z��T�^��Eޫ����lM��"'��r'sP���!+˔3fX�U�$6_p���#���y���ߒ�DT8��뀣a�L' 3Wy,Y"�ٞ��jy�kʪ�-L�T��x���q=�V��=I�s$��6�T��W����a��%���-(p���2�˻ɿ+�)���i��L�8]=��P^>N��Nl�f�ܳAYݰ  �rU�O�@�6VPjv_f����V�U�S!r��I�%i�j
�'j�ЙO����6���ֶ:�Ԧxv�����k(gu������,A���u�F-S���9��K���z^��X��ʹb�e��a�
+&-���76Xd�E�Lw
�X�����]�:�u�k��W�4T�Zk���z\7ji�q:�ʮ2���v����=쁳^���k�BE�Z2Ke�m����/Z�W[*�W_u"'�H�@��j*^F�H�ڎJEev�,-���/TЄ7'��C��Mƌ�'jML�]�,֣k�紃�s0SY ����m$��yM�e�,3�����V���.����|	<F����+���9�*D]��Óļr�ݖP�uп71��>Ȭj�A�b�o������Msǘ���d��+�0�Ǥ�_���g�.jj��P���g&;d_Jg��S�9����;��.�o���Gp?�oUr ��u�[(v���Մ���:\g|��g�|�t�M�"��8.��+}z�av�����vˣ�eJ��K�a�:�k	��^,:ϭ�+5\����Z/�ucl���刧7
��$�v3H��(m]S^��P�&ouk�Y�6|�ee��*qu�z@�&xJ���G7���.Oq|��}��^�}Sr�7�9�������GX���\�G[�pykV생ek��3:ʭ������R��*譨p�y��ﱄ�^���5��f�j�<�]H�����Ӵ�%F3;JW֬�_���l���l8�\E�A�s2!�S�TkfV�-�=�FJ�#�w��j���m���Dg-5Z�tTpV`6:
ZG97�٠ũ�f]��z1�t� t�֟wR��T��^K�,:���/�w�C6PIP��a7.�us�O��]ː��kk��L��C�0u�2l��,vl�2�]�zrK���vk��^�V��n��n�s}�va�k/9Kg��Y�"�^��,{4�s�vJ[4��B�Ƚ��4�oUۤ�Hܧ�f�'�M���q��B���׵�h^!:)�bO������P��Yz���Xu�2�\VV�-L������N�fz�z(�v��3�w"���f3����[��>���
�Ƈ��G�wJ����q�XF�iT�,lt��	�zz��ک�F���Xކ*�N�f�7u���T�3'\��Q;���Y�Q��A�	��e:Z_���F)E�K
�0�Qʼ��][גn1�;�qˤ������ep5���q�#P��и	�G=����^Z�D��*�
�lī�.R���K������[�j��;:�>&�����NVrnڥ)p�
�BX�0,���_�yx�s��0R�^��9�R�%|=�GO�s��V�5�O��i�扼*S;�'U�����ף�p6�b�=��Z8Wb�P����#8�˖n
u!ł��s2���T�*�i�[�W��-p�����m�/���ޭ{�;���s�zu"�"�y9rT.P��Ġ��Qw3�,fM���22�hK7'�ei����9�bEC�K4f�R�a�X���k��+��({�vJY�Z#�5���i��	�Վ:i��%�18i\�,-� E<�L��9��c�<��#�s�;�^���$k�*ԝ5�F��0vB7O�Cb����>�/0�V<��8O��ٹ~��J��Hb���B�;E��څ���Ml�ꪾux9]�s�y0��סi}����o�^b�Fǫ��OO��*C��X%��,������ b~��e���b�����	�ff:ސ��mH�I܈O��6}����R���\ӷ��U��;�w���[ut/�J�	�To+ ��T����ӝ5��5��_A�U�uS6u�Y����v%Q��U�1�~��� � `�g7d_��F��Ntu�=Y/������ޝyJ��-�a	��1|���z�׎xU��e�����FXOEF��Z��c1�I[L�^�K1�-L�ӆ�4M����Y/����(����2Tdu���[w;L��,�u������Y��>4�����ɨZ%!|2���^wr��ygwj�ib*����yp{L��N�-;�qD�uB5�oj�®��t����$���ǣ�q��2��{T�V0�=J�=U�����f'��㮞��.�&W=��Z���/�e�}U�f�~;qS�{�J��讖 �� z#3^������"��Q�٫(]�e�ƣ���e>u�s\�Y�ɍ�"�zU?09�^�C�U�csx���y"��]�r0/|�M(G�2x���vS���RT����L�WR�'�a�ؑ�|U�V�Θ�:J	�dn�y�����>ѱ��#��y阁dC����˰���>�h�xY/=�o�ѧ���D�ǥ�]lz��+��]1n��?9�G
�+i�3=74�����.��t����3m
��4%�w<�\q�����a߲g�jyY��Q��K}�<fZ�  z�sZL��*�t+�/���qiŃ��V�?:κ�+uϚn�O{o���g��ML;^���t��~��'G�N/-�\0!cn���W�����풺�����+eu��U�%��Q�8�\�o�z�Y��0ZN�v\��C����
�C��)�r�g@xչF9}ke(8c'R�E����j��U��G[x/p�$h��;/�
iٹ�17�L���vH��wFŠ��ǷB!R�(؎�ǯjI��"��6]�@o.zu�z�x��#*�x�;�����¹߇����{`#T�<�v%]ҫ3���1L���'�����2�C����%hc��`��ibsk$�(,�b��'Z+M��Ԩ������VkwEٺ���no�JD�v�\����k(e+M����1�]K��tt���R�up����Y�ư�N��9k,˩6ؗx��66h�F��C�����{�y�x�3p�{����LG1��	��P{�gsZ�=��+�bQ������f�[J������L��#�/.�t6f��eR�CK$��ö��[�+��,��K˽�ҍy+�t���i�U�o+�K��k5��Q�n��w4�d��XѶ���t����e[!]��@�ڮ;�7yW��8P��zx���2�Zr������+K�XA9�3�m�)uDWfk���lN@�qSyyoe�	\;/tц[��{�c��s͖��`�Z��R;�mi��:�B����­�e�l�g*�ⷋ�=�[ٚ��c�T&�� r����ԡ#��m����	I:6�X�h��֫�f�C��P���j#��#9̛r����T8�EO�_u��7���0vly=}��4ڻOb�G)hVcK;ʊݮ#��ϡɷ/f����@�|�j��Ņ�\��m���7��uC|+�)dQġ�<㓫
Ň�>�|i=��
��9pw��YQs:Vl�72�%�t
�?.䲼|/�������f�=}U���%�'�,��c��UO)�V��2�`���39Ӹ�m�;���)�YZI|37�@s����FR�+��o�(�o��1w�)QKk��eM��N�]פ�F�:©�ū�M!h�ps�%r��:"��A~���`��lܑ(z�}6hwcLFiR���]�Q-��W�K(�My�eա%�D#-jB��6���b���٣a9�����)E�nm��ô��SpV�炚A���-��&�kR�fk̺����-̫{���y�5[��ǡ��4��*%���gdN�QA=I]nspr�}A�ޗа�ܟ,X�/o�'QJ�;���AH�7Y��L�VԖ��zn�w���ӽ��;їW�r5V�E�B,=��jp̬�|������i6P��7˶�7��L��E�u�kKZגKW����F��n0�0s���-\���t����T�|�����Q����WH�G�Y��`5�%�����Sr�ٞ����n=݋����=�X�<���ᛃ�:��%;-m�V���ֻ��u������ud�FT��I�ITD�Y���9�D�5D�Pfee�C2Q3Ue�SD�SDLT٘�QTPPEE-4MU2�QD4%PٌfRUEDTPD�ED�QM�1A��D�QD�dEUUDSQEMQMQQ34S��d�UQUSUCTD�ٙE�e�fc$�TUUQUQ�QE!I�	TіD�Y�eSPUSIRd4�EL4�SV`8EDER�4aXTSJSU5Ya%U@�DUe�Ue�5D�TQQ9��S�TK1T�Y�AARP5EQED��QNEEMU5L�SCM�TTUE5D��A��CAI35�EfL�MEQ5FY1-$AA��e�A�DTQETES$TQ��SQTQT3U8T��%R��I2�9aS1Y�RE,Q4TMY�RMT˴ TD�g{�u2�Y�'f`��F��^w��|�vt�
�x�BrY������ʰʼ����@egk��&P������H���X-u����&z�܁3�>Q��}�'�r����o�(]���Q�;�����jN�.A���� o6���d
N% 9�/ʸx��ᇈ�Xn%����1\_#X��W5�0A�pr�Öx`*���n{�
�+	�tO���H�zv�ˊ�#+y���I����� �&�7���Mu��Z:�)�f��*#�S'JzX��ov�j˾2�s�������^;z{�9�[���o��������V9���(bKs�� ��^/؎>hξcyc�_)�/Ϧ8��'��A��LZ2�ܝ^��e�L����ML���f��v�LWxs
����r�u�ҹJ���gk*�jDJ��j�`�����c�\��ҝ\E�v�맨l}q���!~���T���V�V#��-���)��Ӎ���s��`N���3'���,3~�a�7Q���R	�Z,kqU��*
F�	�q&�trV:�+��hꡢ9�"����~�u��b���x��_���r3O�h�:ee�Au���c��U~��s �ˣ�{¡�҅\��$�.�ѱ�d���wM��om٣�{�#)ֽ塅�3�6�`�V��WǢӠ�ݭ��_]�R�کu��[ڸ��G#}���!�w�m��zI�E�0��x�	L>�@t��+�u�t��*[�O50�k�)�+�~w��)��[�Ƭ�����kh�Z\oq�/��
x�Q ���x�ehzmZ\^���q��-GL�a�U��-� ��q���7�r~�:���{!�����b�ᒕ/uQP��5k)�[8�ޜ��cy,ʮOT����r���Z`�ʄX���d�Đ���$��T��[k{4����'����`I:���8�$�����3L��t��(1��C
p���l�ұ��qd����u�s�gh��|0;��K�EM��3^�̋�4
��V��@�.�p��N-�x���Ǌ1�0������+g����g2*�~TIU/��m̀��"���)W���a��^ӠX�g\�Jf�tҌ9C��X�L���Ō���6)U��ǇS��V��|�����`�����{O���1�ǳMAs�w=R���2��,�e9WBr�7��{����^��#s���P͛�s�[Ǆ�c+=�YbU�X)�bM�q��-gmEX�M�̿s��Ҽ�l�XQ��u�9S���00r��^���m�`*���gui����x͕��>܄oG�Z�Wݻ.&�LO-}���Z�f����rk9�&*�zg�޳=��k�
�0�C�w�fZ:���'fWa=Ŷ�wu��Z/p�0zS��q�WLú>�by5�L���7�/�tΌf}1�w�Ԯ�G�o�eP�P�EOTF��+��D�vXΗQ��T���[�e=���ŸQ���yZP����|�d�q.�\��R�}��hr(���	��t;��/Kϔ�=R�k�z�I����B���q�{�x���x{)�+]$�̬7�#P����j�d�ڈ�{�!B�YC,��x`��N��囂�HqpM��T�[3f+�O<�y�ub�͸ʵ�gF,}�"��>Sc/��:D;�fb�T�����B��]jW�ˁrCs���[>�oL�l��헊��p瑉��ћ��z��`�(<�m,��m�H�(�17�Co�7]�^�{8J};�#�ݎ�C;�80�᭏<�-M�o��扼v����{����90}H�q��,�P��Լ�Ҽ|p:�t��\kdcj}�^Ad����MZ�^__?Mƺ���Yd:ƶ̤xn5)���J���N��O���[8���z�AMV!���u-��7���u�YD��w��}��q����`�����xK�ͭ�ƾ�J�ӿ�=W7�Czկ���9}-�9�I]+�v^��ѹ�(���
S|T,��=��a�ޞ��u�c�^��T"(���޻+L�$�L�G�����&�"�KC׻�<>�r���҈�+�3.�����e��+�D�����޴2�9��ₜn������|�h�j�ճ>��j���ºV0�F
ː#�I�]�w��*�Q���x�S��x��9�S֞���UhÔ�wZk2s�b�+�I߳g���awѶ�K��t�ֶg��+͢%�fb]��I<�N̷��d�Y��+�[K��uv��V��ȥ���Y�5pv��N�ܙ���=G��AW���մWz��)<�F�{4�^��Y�}�BoV�.�I��J̯Bx�n#6v���P}:��HV���p�VZ��v��=Y���1�e��Y֛ݸ���+R�
��u���Ãu�Lfe���йd�@���s
޻	��<f��6:b�{���I��)��m�4Z;o��j�z+C�Գ�z��\��:ݑ�w�ȡ�.���z�9�a'c"�X� ��W�d)���A�];T/���� '�i�0p���bh)��:���n}W���Zۻ���!�;{��2��Gss��;��Ӓ\��`퓟%��˚�%�0P�,mQ��4��� ��a<#���!�+.�.�v+e����"d����B�ՈO|\.�؎��r�u�Ӟ��xz�{V���9Q��zA�լ�/Z�i�!��=C_�ߡpqu�=����[�ǆؓI��u�s֐�~�����/~nv�[
}\2}���K�k��h�k:K�im���s3��5ut[���<�l�l����b�;�<2�}�YAd�?Cy���S�� ���;GI�J˙�Q��E���Ӛ55z��z�GB���7j����d���A��v�poK��r՞?Ap�8n]�<�G��OK���uZ��)_���P3ݍ�y<Z9�n;�A��]g]L;�S�������c��������j�%Ee�������Z�Ln�m�{���t{����/\�f�S֝y4�{5gV���Ξ�zG�)R�L��^.�]��=��}��G�j��B�O���=x�t��]�(��d�v���+[�RBuܼ��g>v���v>ޫ���$K`ӭn�&�Z��y/�y�s��ս�U�j��}�q�����w=�)ḻ�n�,�Ա@���X�S칫�>U�|-�J-+�;;��uW�Wfsz�a�y�6oR�)v��)M�WU�����5�M�k9-���*x��K��＆\GNy��/%�՝��s�7��'�����j�S}�+@V�nA��.uV�3n�J�k���75�M�B��I��(zu�娻.czu]bY�ײ���7۽]��faz,�WTJ��Zk/ؒ���I����u0'�7r��ES��6�Z�;���4 ��ӿ�ys0l���qʩ���V�)��C*U?o%w��r#��]y��*�yu�����崤��^.��۟y�x%��%�t���ׂ:��v[��b|�Q�U�w2�{�ܼ�f��]^lC��^�x/*	{C�a��c><'y^�r'�<�مߎ��͸�U7
���+.q�@�J�ބ��E�O�{�h#;�;�,W<���egjU�~�X�,t���@]�.5�>���q��4Oa�4�SW�/`�������p����:��e�V�99F��ʵ��7���NRg7��{�WJix�ݨn��ö�0��gu���",3��ц�SwM�-L��fҹ^�	���=�B��:�G��n�T�AV]�����|cY����"��<�҅�����3a+7����3TVH�ت�鳴��H8n6q]���u�ʺ�K}���-��Nr��wU��ø����'gx����Z�ŕ�þ�����+jCDR��7�eZ���9ɨ~V�r�����[���oTs��y�=�*�xw&�BH\�a1�W*�����x�tWJ�v	�OOy�w���$��TN{c��S��P�]`w�~�B��|���'�+�����{��kQ���zz��<���bxZۋ:�c�Y��E����5�@��N�MT��Ϥ�Kl,��.��H��*r��^�=PW	���� gNQ����{U��Lˎ�}y�#:�)`��皓���;Q����x0Ng-4���fm�sw�;�\󾏯�~Oe�&8�������V�W��/�|��qE�c���{aҙ���oڥ�p��$&�d�sH�ֹʺ��^��\��t�8g��p���d�pS�o(uZ1�{j"a���b�m��Ȥ^κ��t�v���� ��E�]�"*s�O8[�")�����]�I#�T�z�gm�̩,H��zL��}0w�i�(�,��pi;�L��>ϫ�`C�g���&{�ןS�$�^	�v:�G*���T�)�v�NŚvtx��kا�*z2qf>.������L^f5&8���J��K�k^����/p��G��2����s�XL�k}��.ɨ=7��𴱻q���W�X�	�:]N��h��{7)��*�U�;���ݙdͽ���]���C�8_A�6]2Շ5l���Z盕�!e�W)�-S��y^��R8����9@�Lo������;�\���1�"�-s(���IN#r�b:��P�crWÜz�9/�|:y�sZ�'4[پ�����7�s=E�����Vui^Q^�Ry����[O�:��,%!���^���E��A�z�&�W�F���J�^ҝs��Wm2�c/�DS M%�l��s`��R7z�)ǳI��A�.�]����O���7��}��&l��;�P�d� ����f�J{�{D���:��}{k6����&��K7��%SǸ�)�R)_*;jٗ-���tw�l�Tȍ(�3���}]֞���R�~��n"Ve'�v�3gCᔢu1��H9ur-f=���J��ݪ�syqBθM��D�U�JЎl��ᯧvPt]�<������k�H�0sח�jU�w>V�<�|3���EE^�E���i+�=I�ܛ�ÏC��>�/ؔ�^��{ܘ���t#7�KtCJ\�kݝ�~T &�;m�1ޞ~���<�.u��]R(\M�[�V�W��囔D�<i�Q����l��f�{ u�w8��y7�����dǬ]K.V�7���v%`w&�O"d���]�U�X�ɀUu���33��s��N͞�[~m�E�{P���#dN�xW�욕�uz� ��e+��Gr����C`���� \jp�+ɽf��8C�:�����2�e6�M`��'i�K�]�=ᵽN)8X9��wN�6� ���s-��8g�;LW"�ə��C3/Op�dw�(��Lu�"%'��%�M��NYV�y�Uk���zY�����Un���H÷$���O�'ӄս;�rW4q�[�	�q�f鉸�]o�Ӽ�.�k�P�wL8%^��s��z�Ԛ��L�;���[��R�x�f����<Z/�mʊ;�3YOݫ�
N���N�ku}
9�+V��%�[H��(���8��e��$�|�;�_Kp�|�j�'��OZ{��6szk%E�Q�k1�ɚ2���u�kzF�>�4�R�}�K5;��׽3V�*��_�����lWF%9��O�Q ֹ��W~���4�7�r�)<������|W�\	�K��{��z�z�G���3�P�yp���os�b�JV+3��
㣻���n�K�)�̞ʝ�>����B�)��;��=���ԎwVqU�FnV�<�9�<e��*(>��:�\�\2-5��L+픟-�nrET+���z�p���O�{��鶸NLxǶ}B�;Q垞'��5Jp��
�b�x���г:��4�9��	�R����*�:)�k�����TA_�Q�Q�"�
���+��TA_�"�
����+��TA_�Q�ED����+��TA]����"�
�����ED��* ��Q���+��TA_�"�
�"�
��
�2������A~�������>����-��>z���	lUJ�P�*�� ��
���	J�Z�V�UM[Ik*I���-iJI��
�R������;54j���հ1�clլ̵)&[kc-�M��-"�MV��͢��fm��M��d�M�!��6�T
ۮ�����l6Ɲ�z,ͦ�"�T�kZڲR�cQ.Q�$��ͭ6Ј6�	�l5l�j����Z
Y��j�#+U�0�-�m���3.��{cm�2��  �H
��]ګ6��Nᦕ�8v �uv����Ӣ�X���C�7)��]rmgL�.��A��v����\���������ի�  ; %��FtlWv۱�Jt���ƻm��ݷu��[P��5�E����檀:�t]]�wk ���vmu��p7�B�P�z�M`���L�li����  �h (QB�
��( �@(^�g�=B�P�wW t(P
(���� �B�s��P�ty=t�˶ۘ�-��S�C�J�m� :۶��˕T�j�f�ҥkkTjIQ�  �S�Z7mk�v4���[m0�ڭ��N��MqJ7r:�C��s�j�f�7m�:�8��4*��n�a�]ԭ�m���-��VUb��  v�umm]Uݶ�k]*��:֍f��[��u+�wm�v���-�lt몎�uu÷n�t������[w*�j�����`���:�.��hx  k���B�9m��K�pWTsL��PUb�`��(	븠�VU �pk&��8 ֝�li�j`jҬ��Ui;�  w:D��MH-�� 3\�
(n�pݎ]Wu�� ���@�0�9��)J�2��dԅlm�Za���  a� ���
)te����ؐ	�h�� e�QC0�֢����[!D�;�6��m��me��x  �x�*U��y��
��\6 5��5P�8�iBt�:�� ����'M#��u�������%E;�  c�^� wk� ��4�]�n�'UaT��º8�Jum՗Tq֨t+w��(ݗ]n��V�=�   jm�%I L ����"��b�D �     �~&BUIF 	�   && ��%T��'�`e0��EBd	�CHъa����O)��A&�Bf���# ����j4ã�Tǧ�q�z���"&������`�R�a�2���u���g�<�1���I	$M��t�yQEA����Z�*���D�? �QPF���?R?R$,Hp�b  ������*��0,��TUoÝ�O�k5����ջAPF ¸�KK?��yD��:��c@��H"4�m��f�p�)��,��5omn]'�4	�mRе [f˻�Y#`�{.��5o+!�Q���x�S�ۢ��
�g$wh6�ˤ��jz���+��yI4Z�Y�v�k��آ��D*��P� ��We^ ăV0��u��axd�Ў�O[r��ƣ�r��;�L<Hz��c�!�u��>
St,]+0Q�R�!�CV��XX�#	�#H�R77r���w�c�vA�f���H'�CV]лQ���6QSr+�ǆ#����Y����0E]FR���-a���>�,���\��)�nL33N;��֫�CX�c���Wbn�(�,uRx��Cq[�2�8DQ3��_^����o-��hw�i�TlZ�V�3u`r��ԭ8�v��V��P����%J�yP��O6���w��k�+6mk���U#����X�wN�p�uu��w�h��j�[CV��y-�v��x��4m��Q7��+����w�!eiW���^��.��s�hm��Shv�\�����ͺ3,c8 ���� �&�4�:]8�`���.-e%���EM ^ѷx�L�W�ݓk#�fmQwl^(�l��	v�32��Z�E��4��w�����΅�@��,<-�Ӫc�ԧd�'Q�('�����X�QJ����f�3Uf!*�L�F�{�QSwBƺ!bGY�n�Z)E-=�q�-�qide)3�2�&`�k�B�Ў<N��pR��)�-k�B汆[z�=��E-Q��,���8���n 
���5�E�!,�
,w��"Ч�N�fR	�n�]�p�Tu�������?��f����[�5����u��4�Q����U�ä���[
�����%�5/�1��ޫ� �a�(��S@ޒ���!l�dA�"�F�؍��(6j��\V���LP��ʕ6f�[˦���M��#�w.�ˊ!���]9��1����1������!��4G�
ًv��� 5�7i�y5���f]�Ґ�W�J�[m\9�`�fR��!�q��v.�^ӆ:��N��l}fV����E&�D(1���6;Lާ���Z��ض��b�b|3M7W��gMH��W������[�Yf���冡Na��U��H=�v�\Kvэ���H>M(��R�����v	LkE�gDP f`���n�Z.˫��Q᧎z�ʖsfMb��Ȏ��Z�xe8��6�l�0�%����eOP6i.��t����V��u�;�i�"�ՙx���1�Z񩖜�4cJ;�X3Vۗ1�V�Ӫ��/m]���{q���o�!�^`9JaGJ�"]墛P:�e��]Lg2ݘDV	w2e릪���xY�v�b�svf�%�V��L�S��
�w�~��Z��4"���	�b���\ut�P������mXZf��2��@,R����GD��L)��r�k`�g%,�H$WZ�3�k@ G`q1Z���1*:"��@k{�	���#�`�ՓG.�su�;oT�s���6�V$t�\�L�78�cɻ���⁔�:�U�v�Z�Ӣ���L��x�*�ya�*if�E���R��x%�;Fh7X�:��wI*%����u��r.�)�G~̈́���{����X�l���m��AR�P��(^f�(���m�X��5���.&�eHj,#vi�Vl�K���#��㒕��N�Q-Ж�5����oVںL
P:��M�=j�:˸�&�"�7��Jȭ�sm��oة`HșU�z��/���Ȍ�u����a뷔�AR�X֬���1śZj	����Cm
Ur�����͚3l�FdV�sMt��\�+S7��OV^S��p]�3]f���{lV{	61m�j�X�w���q���N�XuX��C "[P��TC�I���G�I����*�7Z%k��uq�G.�#��V��fVjW{L��L`�����֨��-�e!hYw{�R������Q�"����in�F�����b�S��d�X�+/M��Y�o.a� l2��9{&:ct�u�ݽ���5���Ͷ�:�Րû�x�b|��yj��X)�L�/j6�[�:��6���:�,h�[[:��.�$�Z)RݙB|�5yY��
4�[�֞��Sa����,�p��f:�{j����5��M@�cU�09`��]�Y2�Z+!T�y��mh��2���kw�����^P76Ҹ^F��,�*�-.�`�U�H�ɗ�(i�d�����P�EL�BZ� c͊�MG��zv����kVR	ӳ�X��yA�а Z�r�趤82nfn�[���.䛱�� �x�����ܑ�4r����q�q�#l e0�e�";[�-�����d�u ����/�n�هt�� ,�.�c2阰�/�G
.�T��*�A��P�R������ɒ�n�kzD�#%c��Ǘp����l�I3Uz�&b���F�a��AH��Q�ܨ�@^�*����ۼ����V�RX��ʷNZ�OAbÈ	E�zYZ�W��l�Q7�2�{a��V� i��(����ndytδ㤞ܳbh�� ��5o"y�lۨ��F��.��C3[v�0X���������W�Č֠%��2kqm�֊��,��xaCa��4�Cn�<ZM�e�b�8��{E�Kt%m��ನVe�݌�ǳT5	@��uwFC%)�
Y���[��٦)z�S���$*�(���l�z��J���GF�����S���x�A��\ŗ����I�����P�°�̗�J�mh��4��(���%i7�5n�-$U�nʟ#(��5/n1+0=�,Q6�J�QCn�h��k3i!�6�X4Y�r��Gf�Ak���g)�*պn�
���|��F��5`Mjk*�Rz5�(��l��Z�ug݊�*����I��d9�HUE�V]mm��q&�k��,i�a.��X��?ǻdї�隒�T�^B�:[��[���.����e]\QL�M��F���+�Uڈ^}�;�c�����
M+j�[�[�K�2}�-Q�@���Zd����Lե��\���iV!�݆5oi�X���y-b۴7!K�4�،w�F��-�R�j&.�"���<w������b �.��⑩5����D����d�sW(#��I����4G�Ud�3m�t��MM�fZ��ɢ$`zE��N���ܖ]k�)C�A=��C{%Z150���T�wM�m�wnK�B崨���]�~�e��s56|��^U�>;ric�i��]b��k5C�������Ħ�<��U�b�"��-���iO.n<`'�Y(���B��SC�H�(M�
j����wt�]eE��ۡ�v�����F<F �Cm����m:;m5ˍTP����[2�V��d��++!� �w0�Mo���u6ĥY -4�=����v��<�n��©0��Ӣl�؝p@Q��LKV����Kt�+��ym !��9J�ÁP+[�z���]wʒ?>y�J�p줂����Ֆ.�!���z������dbGN�dۥGc�r��c��=�w��W��#z�<���2�h���M2�#�V�1�8�B�i�QȜ�1�Y��*�AS&`�zPw��
��$�Y�n�2�qVbQa-�1YԐ�Չ�n5-e��+Ae��j5sC҃0���$^l�o�,�JL�&�����oV:Z�[B�,�JK4q���( F�j�xB��P�L��v��b�Y�B�3lB�{��$9x�]��IKUg`e���8�Jh��4�2��9���wl"R�a5��4���w�{MՒ��YD��V�E�p^�0X�EfBa�x�5%�{Y7wB�1�D���ge�5����ʐ�̣Ek���X2�,���Y�!^�R�&���ǒ�ǎ�+��Vd�l��l�3��Y�0m@�t�p�6(J��K^fc/K3"�wZwK�5�f-m�&�޽e:&�µ�^X������S���!��TY�V6Vޣ(&퉸(܌]�I@�=�x
AΝ{6��N�Mn��3R���L�#ʰ꠵S�pi)�'����6�lV�l˭Ae佤��d��P�?\m�
���dآn�٢ ����&S�XKnV:�lW���[ۨ�ZY�-m8�^�u*Z*�0��2�&MJ�ӻO\��ۣ�g���7"�Q�MP�l$�BT�g*!e�0[� �ct,P!˕y�VYqª��\�I������g-�Vֳ���B����t��-(����I�+^T���B^�ZwQ�o30V`��=�o	��lӷW��֩�6�۬M�W%潌f�j�]���$5މJY��{KB�ui*�4�7�	l7J��x�kLg`��Z
�˲�d�FLX���ڛ>���jyR����Vb���
�����4�!��*ɥ�,%���F��ԛD@Y��Cv�� �h]������+��eD��"d�z�+F]l`)�W�#e��,�i@�v���;ȯ-����5��R�:6��bTh�U,�T~6�w2n=�y��b�ֹ+%���i���FM�K�D�uh�0���n(]��6.RR��:r��&�mg�j�U�.5�2�ջ�.�i�GDpl��H�5�Z�J�,enktȓ3%�ܸv�sX�5 ��bA����O���M4�V�
�cX(i�Z�7����fQ��B;��L�[Y,��	��jh�/n���l0��q�Ԭ�X6�jn��z]�VN"U�E����4����N�F�Z5M�T���v�G[s�X$�O9Ͳ��9���Ր[���̊ ��.��Ȗ�!:=�n�{�� ��z��)��x��m9{�GV���^/[Bk���k$�Q��m�ݲX�3[�Jl��';N1O�r���1gke���r�e%��%]!Kʚ�����֩2��t�6f��V�b��Ɏ��(�
V�[/�����u�m�f$K#3�5�(I|�u��D�������3X#ӵ&�EIjn]�NWw��n;hˡ)��7j��@i�	�0<�!A��0�t5���ۘp��}{�^�N)�������ֈB�jղ(�gH��Nj�)�
KU�qP��t�C����P�;j����լͩu#ʑ�!*�<�aFc)�-����;�1�l�S�L��VL���Gc�q9� �,V�E�U�Z� �j�04KÄ$̨i���z3 wD���"w`�!Xm�1�!�I�c2��[utSCXeh� �fe���YSji̦�жz4>/ �h�Ѝ w��O"/E0�
/��ŷO5Y�C�6��4:g�|���tX�˫�����Si�;G0���EB�+V�v�ܫn�֎���JJ�ku�%,9�ޛ���Rsx-'�`��c[N��V:0�yC �d5qH�n�� �Y9����eBK�*ɖc���M�ӎ�ă����n�X��ɟ,M�[ю��Ui�ϝ[V,C�����s	�W�q��˘m�@7m4��P�� �2�,[�,ڷ�5Y��4��o��`F�K!�fK��b�[/	��-��!��a�.���Yxt��t9s1�롹P\�`��eZ�b`w��ʈ%ekϣ���L�[Mh[1��{�V�*�۠ګ��9iĴ�d
ѓ�Fչ�j+�W����VM;�mѻZ
��)Q�)&�Ƿ�Fh�[�V]nD2�Jj�
�J�diT�\nm��ބ���j���t��n�pAfYo�93\wX%J����0�*�%�lW8�n�n��T�0��u�3k6})Ӻ�2A���S�O6ޖ�b���˧N���6wj�(��V���h�R�B+yr��Ib)��7%�;�N<Ҥ�ߗ����Z��)��T�.@�����ɪB�(l5�m[�v��W��ʄ�}�Y����J�}�+� �=s���}v��c,Lðl.s��a��O3]ʤ�e8Ԩ-��oKr������Z4+�)SJKX�X�7h�j�YLSxq�a�p�I����g�C�o=�R/]m'�	w���o�Ώd�f�N��R�1��M���0��^�}t���I�pC�%]HE��%Ch��t��q f�z�ٚ@�F� r��H��Z�aљ�S	�wDi�����DCu�k�/��ā��O#�*R����Qq��D������!&�i�8��B컡b�S�%J���8I��nٵ�4��]s�-�������Շ��Tj+ڵ\�.�:�h9Kw�ʘ�V���&�,c%����x��������t#�y�eGΥG�溈Vg+��{'U���.�£��ܨ�EwX�F܍v����a�C�0`�n»���
D�E>5��X<�aO]��4b2��
�����Ȅ8�
�v%�܏*c4�Ė-ܢ��C�[�WD�ܐ��u��T�U��i�Q�D���Y��si�568A�9	��iy KO(��c+{aҹ�X�B�ec:c�z���5<����O-lVj�4ʕ�Lԥ���ܺ�pK�{��Y'Y�35�%��uL��̼;	#�������j��8�(-B��xC�a�l�nw�fWm�/��d�O_�wK�*�%K(7�Ɗ<湐"��SEXB|��`��[}�U̠�����s���^��3Wl��E+u��I��N]�oK�9ewN���ZHV�=�a:#���2���R-|. �E��]v�K�����U�:[�������L�2�ome��z/[9�n+�vn�jr�WM0=��j�(��I;@0PB�Ӧ�家��fʧe�M,�%돺��]�n7��ٔ��]��6�U��Vv&��N�|�_)ݗ���gK���OgRx�v̙L��i��uh���y]2���z;M9\�m� ��@�<%7��B�Y�i�]��$;���4��-��HT8��{�^��5r��&�儻�B�VZ���ݜ�������d�ۉe���u۳����!�}S�)�l�s�~ʊo<�iW_��P�l2�]o�}ti=fm�m�9��waԎ��JJ��k�Tᇎ�\q��	a��N�-�hs�nAWā���m�=GX���k�rqT]u���f����I������gk�����V]�QB�|^��Cv���Rm�$�� w��/�&t 4g;��p��
�Zs)`����X�:��֢��P;�����^p��T�O��T����4�K	VU��y���F�U�w���%C����P��s�ca��<K9x��mj�=� Ql<���/�oh�o1�g@��y��!@Sn�Քk/���P��5�l��OL���ݳ��z���<�aw�铻$h��Z_ �U�b��E���[�O*_��u��u��)��p*)�m�V�c~��/�=�wQR���=�
n�Vu�.�CzX3�Β0�AY�[ZWTF� ue�n�.����/K�N[�yb���fD�h�V�����Hpv���k����8�c��B��R�x��e��m��y�М�\�w5���%�(qOR�/����0�^:
�r;�pf'Sxl��	��K�qN{��b�����ha��se�eF�7x}��ۏq�ס��C:(�TQ��0*<n�,����2&8Nw';�K�ho�Iُv2��m�hd[�wk�j�<.��/�^o'����Hs{%��MY,�y��9�]��l��F���Fko���!�M��W��`��P�A,��@��x��|+s%ԣ)����@!�ڃԻ�s�w��k�7V'	xmG������ޜo��\o
B��f�c����%�j����v=��.:S#�j�Z�muih����e�x3C�h�WGr�-�K�%��#�̦�n���n�wcv9Y������O�ӠR��;�#���P�W��btc�A�q`k�N�wk�/��c�*���صE5��w��gI&�T�Y�b�؎k���k�����AǞ#s�z\p%��4l���_.�!mkz�I%!������Ke$�d۴��3(>�emx��a�� ��e���ɠN�k8�fA�󅌖&����P-sfvJ�x%KE�DEà��*8���g/�YLح��`iS�����퇮
a��;���1M�T3����1Р��ڙ"�Z�d�v�O����lvYy�mL
�pV_&��̧ҥ��J�r���A�:�$ɲ!1X��j�R��k*�J �8w�5��{�Pnb�+x�%��*&\�ا�� ���nel�D���v]A�#lX� v㏞>f�l]f[3@A(9�U���w�NjU�b��é�溽y�����U�Kzf��:���ę+[�퍕.r=�9^�{��7L�m�	��|hI`1'wR�q���ˡZ#�Xo�W�1�Jr������k�k��P�b��l.Zيa�B�T�5o;_U�殝��$�����X����M�s��\0 �r�8�u+丵V��0*���U�̀OdXF��s3CEB/�P���N_W@�NZ5�^�ۧ��Š� ��Y��^u��ӽ$�^j\U.���:�Rd�kM#�X;{��ݣZfI֨Z�b����f2N�}S(��9�1mk�4_��W0��������ȫW���sw^�x���ϸ��Ӏ��콰u]f�ܘ�)�]o)�-�co�S�\���bk>�(U�CO�y���}�7��`�f����v�G��.�X����Y- �%���������V�ԅp$�v/.t��XAF�-G��n���&��4�Kx:�����^L��$��R v�ec�Ք�opţ	�֙t^:�.`ۺJ7�5�{#���-�e�K!@���:�U2��u�VV�|�^<�"��YQ7{�l�;x�)>�^�8jΐ��l��1�OE�͕��3�o`9ۀJ;��R_d�ܩh�{GL㯔�3�fY�^s����ȅ�U��4�}O��'�ܳ�����;�d�,'yn��KV��cvr{�R�TNmvfN��2�G��^'��2���@R�qAS�3�48�*��,Y� l�!��4�h��=B�eeH��]��i�_�E��{a�A���2�]��;r����*�%�VX���"�¹��ܤ�`�d�e�.�MǓ�`����ګ��+vS_n1qʳ9�ynnkH��Ĳ�z���>ܴm���;�BK�]�+�Ի�bCP��ep����jɠ�����;��8JPU���A���X��N�ڽM]m�C���a���#��K*Mc,��SdU�4�l��g�KZ:�\9./:�a㛶������$ȶ���)4���"�H�Sџq��tʷK ��#׽r�\ �;!�J�;�[u 맹��g5+1�e&�1ΥӠ%f鴝ꘑ5�.8���/! �1¤���o+�*�[��i���bK�ְ��@��iV-:�R��A�E�#N���ަd[���xU�BTv�o:��}�kt�`璹Ւ�l��Y}7s;�����F��k�V3^*]��|7�j7���,�3�Oj!ÓWJ��Ё�˼���
�( av�HT.���O�=�}�N4f�"�\du��ӹE9dF�����h�{��Wq*rdKd P+KR����\d� ��(�����ns�׆�ui����ȷ4��5�����:�X#��#�#xtX�eM�i�}��Z-�E6�v9�3�xbTR�1��d��U��{/5v����51jjW,:�9b#�'��(_;}Ci.����Q�����}�uy-�m]��:"�-�RE���$�F�&HbB��Ӹ�@�oE���e�q�2f>�d����2���=�;ef������P��y�Z��7�ш'n@�H3��h���7Pz�R�vw8�0�K.�px2��)�It�"2F�3F�ֻA���t�O��u�+_$y�$*u���ȩ�u�e�2���oN��ZY�WzzUʽ��:u�}]���R���euj�7r�ZAuY�����}q���z$`�f�	�e�R\Ǝ3�2�(�"��tТzvVv.VQ�wf.��9"�Z��:��;�R/ �ݴ�Y��FD��,c0֔��7ws�\�T_h�/�}�-<��52"&ݾ.��`�܍���-��:�l�N֋�9��dJ���[��A�N��T���7V�!c��4^�{6�����b�t�C�7#���		��&x�쨵��ǬJ괯=�\x�Ϣ|��M�\�SMK��b�/�r�o9��T�$[3�²n���T���EL\%uRB.�גF�|zf�9�*��R��bҬ��v�O���hz�q�2�4�������mɳ�U�W���n�Q��̥#��V[�[a������2l�G5�\\�TQ�p�;u6_.�lK�'d�CƖ��w&.7*�]g$���R�隖�>�7.��&�u"ҩ|�ۂ��.JE��b�./0Y��yf��n�d@n-���+�ʱ�M��)��|݉@�;,oP�Ip���H:��d�a8FSt���n�Be�,����Ƭ�K4�(s��HI���hJxe'J�A��b����&KR��ك�t_,�R�d�p�L�,u�䋡�!mᒷ�uJ@Z{��0�+h�}x#eԫ/�r�3(�Ql9a<�� �&�z�}x;+�Ɍ��AJG+�t&��ʀ���{϶�ҵHe@�:��<�o�[<�����{�i������-+���,|&��������s~a�*���V�fD6�u���S����c}#c�����FikH�nj��hs�HGQ`�}�[�R6���I��2=��R+��Un�w�r�݇�sS1�Ҽ�E�lCV���"M�3Y/ȟ�_�]Nޕ�oD�f�V�ܤ(����r��ϵp�a�3�wkoCj����kt��˟u�;ڰ^��[lr�)�d��d}ukm�t��-ؼg�ue4�vH)nv90�W��J��K����vU��7j>�6��6r㚑��m�2w����DZ�$���1�0��;y�wKj�EG�y��1��=��bк�T#�o�"fǎF+9��هOoQ�ɩ��n���Y�DV�sU|��=2�^Ū[B��{}W����Z���8=�:��֧k�����_Z���=]�hd���']ى:����.�;31ɽ&�*��pUٛ�.�
�fNj��ٸ�ںGtH��o�Ӈs�a�77AWH��y��U�!Yy2y��|�� �Lڙ�E��[r�Z��r��Ur�rG�v�R��ˋ�n��s͂�E
@4ۢ�WX�t�C��Z��"ㆵ��b���o�B��(���g9���6�5����V�ZF+64�yxŎ�&_WDa�P���w,̻K�5Ky#G�
\�5�B:�B̼�k�{�\�U����%����J@v.2G�m*x�T��Y%��7�j�{^E>[�H�'��l��=¤yLZ/�X��ep�fn���[{S�������uo�0�f��i|GWE� #q*3h\MX�+��+��FҖF�3��L[3AEV��Gg�P�����7AoMv�e��u�I����X�u�D�?��/vu���o2�y�6������ �]I{�tފ�t}(�m�ppX�\��H9��3:��>w\lTLɸ�Cf\s/nfJԁsZ��Fe�;�EfnВ|���]	18�w�������3�vїUx�d��=\�ӟ+��ٜ�X�^���Gjk���B,ux��15	�՜�<��2���b��Ð�A$�7���-�m]��v^8�n�/y\��t���Аf����2�����Ғ�0��_a��a��F�m�o_���U-Kb�qoj�:�1����`���Q�5�Ei��p�PaK��.�gjQ5����S���_,&���������r�����
*�Ԑj�2�"#��(t.'0Ȣ�#��^�ɭg}f������+����t2�j,I�ϴv=�:�������Q�{s�9�!7����q6d�i�)Fe00�R����
��q�6�,�'g\�]@={��ret�pB�L����!�Ⓢq��ն3�E}¹�t�g���xOJ��VX�(��+y��X3��i�c5�bmqu>��w۽�+�+`������j�n`��i�H\�ƫ.7�"�uLz�'����qN�m��m"���1]Y9�is6�Oo�5�lA(�r�G�����u�ҭC�Zt�2H���[2PZO��O.�^������9+�H�8��q:��F�3dd�]�MM���\�'��v��S�L6�8>�ج;�.P�r)������UC�f\��.me�c9ӽ��ZU�Z�����wz�źqp�i��#�r�fq�2�u�z!�{A�*�4Ma�N�O �2\�
�հΨ!�7�ɦ�2;�'���&%�8�����)��jg `e�}$ވ�8{���iN����>�4�v �Z��,4�C
�j��mYVxM�@f��v}��3Z�My��Ƣ�x���ֹ"Ǌ��c��TYc�īNj�۵�U˟g
��mxk�[��L��.�ȭ�� �^�#8ܘx�#/E�;����.�ݙ�g�Պw���w�$hu�)'�)P�S�o-/mv�ׯ�� �1h�%*]��$Z/�o0�L68��dʰ���N1�"�5Eq+њU!��J�^�B{k�`�
1\�ʴM� ��`�}a,�5��`��k�BI��Z��sȫ.������+W�&ãJ.���-]须&V� �[6䥸��]ћ*n�;M�Y�����@>��ۆ��J��t-�shT­�Cy)G��Hb���-�f>���΃��6�{6�5�Y}"ݽ��x݋�n7Z��J,*��+U ���V5h����0�$D����E��oX5�:���Wg"I�r��E)�뀓��ƪ�ړ�y��b�O;�Q#��2R�l|w���&po�Y�˓'^��.GOp�0:�OX�O�ٍ��U㽔5���`K�>	%9γ��Y���C��ۥ�	��6�a�0�����f33m�"K�B�[T�=���PTb�C�X�Gɠo���p.�Ga&�mԦ�`ɲ�u[���;�%�{r���fV�;��B]+F$�ҩ]X/4W)B;�噵)�1J�A�?N��*!KT���ÊV��\;d��&	�;.]Ⱥ�ξ\Vp�Cz�yZi�
�+ELN|+��b��˵�ﳩ�%�D�r�@k�NkD���Yuv�]��͛��g>׃.<�]N�E�e��6k3��hQ�#����@�ԯl vv�Cee���	�(��m���c�J�Z��+6�ә}g�`*YEk8;�-��ߴ&���TH��a!4b�)e+ࢽG3lB\l�k�	vxH�i����h��t��U��YkyX�d���YW��(�0;P�	�ew�C��CS�V�5[v����1X����=Dmb�BIm�M�q���7����@��n����V�;%����j޶�XmF(�ȍ�c���,V�Bh�7��s�䳜3���Ƥ-��v8�E :W�Υ�F�z:�8K������:�X9l���W2�g\=0q� �������K�
B����0`���@�o�j���kR�f}�����ޫ
_5q-�Ȇv�0��6�j.e�s&Q���6㾮���fq�\���L�JHmGhT�,rP���t�]<ki����r�84�Z���+b�����N�u�y�O2��|�UƲ���_S<�3㉾�-�q��]�{2���_A�v[40[s�+7��ͣU�o#*pݺ�G�F�u��lp��D�VY��v�hY�*|b�W�v�D��W��s<,*�B�b�)��[ru銲�Iw���U�d"�{Cp�d�U��WMg�/�6I��QV�U�K�ao`Y����^Rn�K�y�䧯��87�ֵ��2]�9f=�)b��T{��u�^�{�.�T#D��r���=;�ɂP������
�=M�9RW^�=[ִ�GM=�*Ց�����jqx�[���oR4���e�9ٙ��>���\�K�� 3f��z��gqzm��"�kl1*m;sdz6�p�b�V����FI���Aۑu2�vDB��@��c{�~%��m�<y|BL=�B�GC�Q�Wz�z�V/�<��):a]8�3Զ����r�-�V{��D��)�u�zWf`�ٵqd�8Z��VH�M7�%
=kZ��)��˨"B2�jSU���
�Jt�;/@싓�M�fC�7+V]>NB��#Τ�[�Wf�vM�)#L֣��w I*�� �p����pڲ����[y[>��H��'4\�*�u��Å�%����u�1���rv9\n�����n6l�k���z^'3�K4aM�71�]W�]#/驉4(3$쬭��J<�k1$1�-`��QKݤ�q��6�M�r.��y.�F�n��1-�����2�M��F��H:�t�w.�M�.�f�K�`7ae��ے]ltD���Gb�䮕�CM�Ư�S�cM��u��9NL�3/g2�d�#�i�jA�����Ǘ�n8��f�s�_@��g�]�8�m��;x�jP�R"�ٔ��v��1�1�Jc蹄���:;F�9�rX��8M%��Υov���tU�6�N�,��E3�+����`�L�.��r;Xn�2�EyB�J�]�|�B��嘑�q�j��g!�����0;��2v��.u^V=���l�6�*�����]s{��^��̽���ھ��nb#+d��L����s�a���j�W8/�,�q ��Z�AY���:~��0(3��2)j�w��Ή��ʭ���{�6�u��qf��T�j����	`e*n:]k�{,���^l�;��Q�Ԫ�w�/i�U���5��&��4���;IoI��y	$���Mj^�U�bxr�#��.\5���%��S�9���=wl-�Eq׌N���M���*����[Z㥲Ptkz�C��4õǟ9B��uuό�I�[T�Λt],� �3��.q�ui��y�ݙjhlHjo�9�n�����e6.��l(/H�uj7��+��jm*Y���}�cܙ�ʖ^��3���*h.�@bF\�%�}��Y�t�u	�J��#T=��s���9�Y�3J�Q�P����㹈�ѝ'�0��� �y�y�鰳(�����nY�W2����oo�n:���'��h�j��;�!�t�l�#,vR,r3L���چ��b�T�GuX���
Ss:f�'g" �9PSX�fCR�|T6�,��Ҝ�%3�^�M��T�ub��A\o^��C�ӧٛk�����䃰f�7R�F�����s��q*����B��"q��GXa�mAz��(������d��ǻG���2��8y��F�l��1P�vmW4se��M�kE]ue�kzR��\4e��h��h���5�v��mO�{u{���nZ.�����s�#�䓷@���Zc��0VS������C:t��e�+C�:�J���&ݻ���쌡\����Qk�i�ݭ��r�����ѕ�����Q*wo�y��8ݱ�x��u8�1�%�.����]���WA�.�*Į��"r��kf�=G.�+U��2u����$��S)eb�@S�n��b���z& ڲ�#y��o3ku�+�ْWn�J�u��d�܎�u�/U�$*��Dҧ�K�НF���m�zl�Y\<xk�K���ae�m`�])EJh=���+:oL���78��7𭣐 �EMN�uyv�e3��З�[��m�;E�V��TF�vن�{��yOC�	F1��)���#$�����a�	����$��V�"QU�����7p�&����V���ۑh���	A��������8��/Dɐ�Hq��ʃd�o;Hsz���k*�Ԇp&�z���Ve3)��.���h��9C����n�^�kn�Z��'\���0T��oE����y*��^�9���AD9�;��[���L-�ە�X��5�,E�v��]K=�-�;D�y"6w[��p�ͅ읐}wkim�
N�������f���袲�90࿂��[����1�/�#�'���ʊ���\K��W�PQ���t
T���n��ycJQ�K��V��V+���E�Kf_W\'El�RViua�/+`*%C�aܧL�ܱ�J���=��Y[�mRJ�,���3gY�L��ڹ}Ր�TCtA�^͝�"�!��٤�\s���t,xf�Z��	Q<���LZ���Ҥ�'d2ķ�^�V��F��՗t��V�Ă��*8Njeon
��ۗΦiͭ�ʾ���rUv��6KţF875�8����s=:�u��R�3����mup=�D���ut��$���2��q]4c�{p� �K�mͪF���%Ӊ�X1fJ�5
�r�n4n�)��+oD&인����}6�JKܝ*V^ɔ���W��J��q�L���W>�oG�7�kOj�f��Y4d݌vyX�9&��<Z�F�g���R�{*+�+����l�A�ӣI��i��d��	aI�t �G���`�V�'f���[��R��&��	}�I�7+zÝ1I�U���G�yIoK��ߵh{)�&cw>��K9�ǉjx�%z�KRXti��\"`��uf:붪��]��[�Q��+�
�I�V5ɉ�qȋ����ޭd<˷���5�q��Yr��M��<�;p桋���{��lY�0�]�,��ֆt�1�V��}%`���N����u�vĳeAYyH���y���8Tt6�6���v�I/(����wg�m�f�抟;ϣ��)�ʹA<�0m���^#�n�M��o:�?��E�T{��7v�ޡ��*t��]q2��g�v�]�fv�!��n���񱷘����;>��M�
h�%^�#3�Gm�e�j���j#&�n�m�rY�H"a}�U��䙺�^�ƚ�d�Z���k``��q�|lD�]�QN�5uҹtԹT#2��̲; )��J_��G���8b�>�݈^u�į�v�h'!���Չ�������x�LKY�1ds�!����Ţ*)�u 9=�滕*�T�y���N�=�c�v_Qo���U�ݳx����a�ᮩ�ql�p'���Z˅�ͬ�$��\�h���%�̣�ɡ<����v�����޵�k""��@ss�*.ǌ���afJ�����j�m�.ˏ�V}Ư�u7!�0MD�B�t�,e�+	�r�볆-Q�|lZI�r���[}�L9�:Z�U�b�.]�pSb�W�<M���.���`e-�j��$E�n�[�K������Zjq�*N��Cn:=(ԧJ���[��GPl��ͬV:�l�8�A�[t^jD^��*�2�9�+m���.*���V�
x���.�l,ϔ���s���ɣ�(��uq�|�h�a��M�^�z���N�q���H��n����O�&����H$Tw�R�]O����I�JN�QLl#ʞ��]����q��?�ۣS� �΍w�ڗ�x�iy(��H���{X��7�Xr���5��	t�ks]�Za�V�mL��p�m���ތ�nu��:)������uMΎ�b��i�|m���SF�r�~�gR&�v�ߕ.��Y6��|jo�hvs9ڇ���٢�PxM�|w����&>KWv��B5�Z��q�����w0 d���$B�][ɻ6�0o�qp�&X��n�CŗG��_	e��$U���h��|�(`T���ؠ���q�X��wvk�	*�:������ˋ��F]
�7O9���Vms\Աx�up*�OD�C{�6��{����ʂ�Iv�r
[��1C\��v��.�7�p�S�,�@%Zop�|��[�Z�Ň��렚O��,�K�}XL#��Wa��,�`cz�b��6�Q�M��H�6�LK����!VE�Bd�t�	�� ��Y=��?���<�ލq]�
9V[��	��H�˜.ӎ���لT�n�`�)�,���[��!��:��lG���ۻά�M�ͬM�dQ��m���BM&��R�	`7D��F�)5- �+�4��h������8ZvN@�q\2z�n��vڸ������̡lA��xp�=V��ͽ�l��÷Ge�^�s��T�gu,�G�ea�]��Vhv��e˗dr�6��aO6B���yW�:�����l��I�A�,�4��*�u%�x9�
���`ʉ�|���ȋ�#|�&�e�Z�e�`_hH�2y��]B-�����5m.����XmZ�.Ot�w y�g97-�iRV����26V��ʉŋH��7+�mmsA;����b�p�n�2�5��ܺ<-(��l�)�A]y�k���e:Ke@խ��IGz��ֳ5 �2-9�_5h^�`b�*�a�|��)v+T�r�xyn��)�w���`c�J��VѮ���*�]�f�t[Xya�cU��{\,d��"m�U7ir�݆�t��.�4�]��v ���3�l)-�շqI�}�[f��/��gw�9��YA�bP���1�T@����]ؔ}���*����2�J���P��3(�Q���eۃ"��qsl�֦ �"����J(�	\b��Z�*ш�=	���-�+3)+ڃlYvֵԬ[j��5��G3�-���X���5�b!�����r�ˎ�
%b��)�\W]d�2�������a�U-2��d�j��7i��c/M���e���L��kTLf�V��0��+�k1k5��F�f�\���5�B�]�\���vȳZề�TƹiZ��6�7K���5*�s	�����D-L�RfZ[�k��X6�r�\hkTL[r�1-�Z�n*�Uq�ۻ�\���Z�ʃj&��)m��m]�[J�kIR�E���fUs�*�#��V^O�>�~2ړ�B:�閙�M��](oY�5�8���{�0ʚ�]��Ni5p֞�oM:��J����RY/7�T`����PԖ�%����R?���,��-5�}"��0������3��i-*pT�)}�?	�Vs�*P:-����^��ܪ�n�$w@��7��(K�HZE�p�nY4�'Á�"I���Uz���6C��6���w��m��IP9�X<Z�r�;�>�ˁ���됆�"����D�Sv\�=7MF���E�1Y�0��c��$6TPS,E4�bd��0�f�+ww������(�N��C��{ ҝ�Xd(�a�-��;,G�9�"��-S�A�U=�UE�M�x��
d;*MF^ʉ�ڑ=��� !="�bD�s����y��K_j�ˏqiفT�((���
����5�ϵ?�Ǉ�9c�f���!S�p�ݪ��$m9M������$`�2����������j�@;�x�돉TE�]�As���o�����U�A!!q��d(�'(ס�??�"���u0zr��ݩKNe�8r�z�!�mc��F�aե/5��[�q�EmE���q�MYI����.�?��[����q��m9:ҭ۵����X�M��]Z�b���7yR8�tG�t���[v^�����a�
a#4��VG#ꋵ"��{��	
�~��R����K⟷ ���NJZlSFB� S0�>]@ut6�\g)�/b߬�ܽ
�9���y_��뉩Q��95��qV}�4á��20���C�A`K��'N��Me+x���C���z�ng�1����ߗVk�x�,T���\�K�����BQi͞,UJ���ё��p�P � ��/
4�����5��� ��{Wl�[��v��c�B�Cvˌ�9��5�G(`x�~�T�[��M_c����VFã�Յ^�6�XC�1V�\�n\`!L!P��2�s]���Sx_V�k��,9��������R�*��t�>��S�b5%J��ч�[�ܥT���-C}Q�fP�lF����J�Xq��m��W�U1��A������e��^�&F@,*�QL�I�ܧx�Ŏ����@���бHk���ޡjk{�$Է��R��Hp���q���{�t��vk��zu+]��G�L�.�=����4�ہN��=ǳ
�NbW�s"5,n�a�br!u���6�:�Լ�I]�Rr�l�ʾ���v�ИX�����5�*�P��ʮ+�n�/3ε �M��C,&]���t>3@~�B-��E���'�#1p*�C�Q��g7Տ^��q�[ɨb�LC�.s��MI��LUx4+���9ěe[�L�ž�uO�[РoL���>�1^ٸ�+���ھ);:Δ=��ڐ�:���͍��Ю��X���}^�!���D9�P���)5�"_8�l�\]������%���Wz�E�-�1��:�n@��J�l${����+�f��༜�ܡ4�����b�6�0S��1/
���ô�ۋC��0?#�U���(B����ƹ\f�牡V�ϑA�"�:S+�;��Y�箵:lE��|����3̴	���Br��z�џ��ET��� n��x�p��bGy��豆��n�Ey��Ys�Z&:��AW���\�St�%�ʧ�^�����u��-֌�,U���E�ZM�b�V�@-
�� ��}�)Ʒ#�Mв��{u�����G>ݪ�֣�K����G�j5�p=7��f�^7����2+-̼{!�}�4��hɬ����X�㯧��^0QkC��F�DU�W&�R*
q..����՗�]nk������|��1�:)S�������.b�rfK�T3��u˒��čS�����iT&|t��xTW�8˾���tv���37m+��y7i�Kj���V�\����²dC3�@��l؏dJ8!'AS���\���m�s�T�	Apy�Z$�.�TP�3��L3>��M�t��)R�3�j# L�Ǣ��0�LA��w!Êj'�|�8�1!Ǝ����/p�W��
/K����M̶xi�B��'�[6�G��0&3������u�\ޡ�cJ��a�*r72E�n�8B�i�/�(��HJ[40K�4�ZԂj��?��4-E�5a��x9���h��Y�.=#B�\�Y��:��g-i�7g���W�H�i!�:�T
$�D������孡����k�/���@a;~A��\V���Xje��Y��d��֭���՜�Bxn�e�4���M��s�P@)rJ��X�V�hƯ't J��6��zlCZ5��yc�]�<�qK��Gr��(�t��2�\2����;���ޯ���k�M���u�	C��e��i4������2���E��&{�{jU��g�L+@T���l���z�Э��?a�WA�w]L��y�V5�P�vo��JcO��%��:'ܖ�+��?�ρ��|89���>��KV�ahD[��Ǣ:�zE5#0Κ��T.���L�+f���ƨ��ip@��J�*,	D:;��]=��b���H|k~�l�4#��u��B�p`k��+"DA�>�G-�3�*C���k/5X����O�c�Ķ�m�Ȋ�*M�&���#��!W�����	r�.f/}�e=�Ox�<+�X'�~s����5ˁ��⃠�8��&8�i�D`��'����wj	s�9�li�Ɔ��$6TP�ߨ]{��V�xR���g
nN�=�z�MP�3�H5��ف�QXbKw�&@�b=1̱�&L�o&��p���=�F�j���S����QHޝ���Z1�]ӭ͸pvs�9��̺m�8�v�U�maih�
�z�<�vO%�{�B�ݺ�g0^�d���:
M�ά��%�+Ǣn��D��2`�Ey�Ӷ܂�s��.A^U�^5�b,e�pB\�I���?��]J��↱"�N����5�`��u!U;_��_g2*�x]xX�����}p?�y�
��L֛�ͽ}�6���m�a�Ȋl�Cs6�Dף��#�V�1�'���^d?mi>�N.7��Iy�����W0t&:r:�j��auY4����t���'(ߞqf1n����C3�z�C�B]�"}�}q^�\��BU�ok�/E^yBVj�Vf��z�8_
OU�Z �
ʾC������o�Xʐ�.,�����sz:Kv��?Ae�������fl�zP�퉤�H�=�*���u^����S3�Sei{t3y�pG󪊖ሡtN�	W��ٮ����T���4ߕi��xu#+'GA[f���w�:6� �Pϖ��-�EǸPT٣T�N^��c#�%�K�`;��ˍ�/Ȏ�!l	
��"2!���s�L.����44�l�4�-Ǫ@�fj<�wR�6��M�����lJ�W��|�d�z"�D�0����eR@k��<�ѱ�$:^��L�4<@� �4b���=�YY��CĒ�R����������W-:���
��I`�����GA�~f��9�u�t�=eC�1^����o��ߏ@*`i
�^�owP�{̈́4� �>�(�vˁJꃞ�g��rBfbD�PO� aFV���[�&�8�a����v.�2ԍ�R�
����\�P���Xb�A��]E8������/	�J1�X@����SOt:�����
S�E�!p�p�f�	��D�)�q<kW22g�Y4�atP�Z��<LQ�9=ݍ3b6�F!����5&2M5"���q�6�Q��A����_o2�y���
��'Y�S������8��MI|LNy�]	�93i)F]z�J
sK���g�GY��q:S3��蕢�lU��؛�T�o�9Y�0���7'!о�e\� et�T�@Ʀ�GH��w\
|�x#\!����-��4�핕;nGE2��Pf��a"�1{B�-�Y�kKGI:n�� U�L]�MG�j�v�Si3��y�v� �\�پ�~�˫[]�����Z<�{�#N[Uc��t{v�&v�aD�p�##E��8j1\L���R�ǐz�T��ҫ����O�_okLJ��_H����|�]
lMa�"b����h�;-�x���g4������n�A�g��\Z/b�(U��^*ms�0�"��T��PgakQ���y�a2i��׳�;���^&��=�>�
}�+�e�	L�l�k,��� 듽=XP�ת7J��D^��JDW���G<��#��������u@�nQ�^M�+�@��;�}�;^�&QI�q�H�}}�h߹S�^����S�^zW����yP��}�:#�K��	U���;��l�(����a���$�=H�U)ImMD��:�Bp�F4�}CJ�O�<�P�0��ຏF��gp��bx?R��]H��/���ֈ
x?�{��W.������NY�E�,O�{���#h�=R�*ˀ)�Z$إ.*��p��0��ʴ'dꚼOX=��KK->��x�C@��|W�S�S�{�k]���Xs;	]�����Y��-������Wa�ⷮ��0��J7݀�{Dss%a�*��"��H�*��[��׳�y%�������g���BP�h��k�I�n�24�K5mj]����-�*�Γ�93�ō5*g)~#`��~W���M��i�� ��Kfو�����O;���G�]{��+ҊC�m�ݕ�V�zp�#e�!D�gٽ+7�t��U�x\�L��
�g��j×M���|4]c�^*��W��V� R��a��uz�$�he�I��ή�AU�ׁ�-m���Ft�Օ�+_zMNU���>��v�}6��8e��%r�2+�6M�b�¬�ɬ�yM>�
����#�������B�q��Y���Tn�j���?uz��Ln0��;Z�9p��:řt�>�=ƽ�"��u�'a"�8�A��7}�W�]���9�ѣ�q��KG�h�g�A"��C�>�WK�Vt-�ʁ��7U�>(\�AM��K�<TX��v	��+���Ԩ)2�������A6�Ǻ>7�w�й�_�sVW)�̼�H�#��F��q#���:%���n:o#���+p�P�[T��[�S���x;w&��iyQX�Z�<�q+Ǧ�Cb�)��j�E�<�P���m�b���5I�����^��r#J���a25�c|F����]5}t�ec����?<�L���H$����Ϸ535j1ãh��*d�ܐ���Dkr��+�Eд(��af�&kׯ�|;c�[�#���Y���jj�m�Ul�|4|�.�x:��!��n���w�1�z<\)�TDΌ.)ߺ�3�*(5LCNv'�Hp"F��U[t�l��J�&��k)G���"	oGP����̱zxh�M�����=Q�Z�����5�lIU=~_�]����"yӱ0���#i�H!�����z̄����P��n�W�&�VE�wJ+L��Jx��y��#q��!H��6l7"����Ϲ�l����]b|���P�r,���ڨ��v׀a<3JC�c\<�@��\
�o�_jd�Q��D�ػ۬u�t��Iczx��L�B˄"�l�w�Y��ϕ4U���|ٮ��˻����2���4����v̍�@�Z�f�.�������by�#��D��1����J�����wh�A��VU��4btQ�m%�J%:Ǯ��ò����J�)�|\Eb6�Q63zE��J�R�q%�]X�ӹ� L�.veo!xyT�X{e�;{3o$T8�Έ��c�ՙ5Н��|Ѻyu�MX�<9p�:oN�V���Q�F�<���du�Q nB��EϠN��C�e����kS=n��M�����X��5.�?���a�\���	�f��)e�M�i%C//`T���.-���O*6��7'P#HԖI��a��Kg����+3`����F���o��[u�2��x	״�E��%r��-r幹i�WE�1'mQBH��-��v�^XƟ6�8��D��g%��a�Krh7:�0�D�P�dOxj8��H.u�[s씅�ꩵ�̄�B_����tu%���j�f��K2��������%�P�� b�.�^��N�,�p��_3��z��n�
�h̾7:�K������Յ�r$�s[ܾ:�&i����Ṵ���4C�Jnik巕�Z:����np0
|hu�r����%��r��Ͷ~�� L�&;�MSsr�o�L����}�����v�v�u��ٵ�v��qI��ڝ�s�Ӳ�.X���E��rc��7�'����z��˴�4���Eyh	E;v���7��#��!��eJc�;w��}ئ�ȡ�#L��ZDe�f�����\&`��R�r�P��T�β��nH��M]���j�����PP�\[��>�v)�Y�� S��fdaN���ˉf�t�+��H-�U�����Z�\R�ĸ�ئ*�H��Rb�`��Q�j\��#Υ�	8��F�l�UB	WQʋrm�z;5�;u�0r�R��le�W�XZ�o:�7;6ѩ���Di��j�,T5n>�Q�v��aY��iP��(>WNjg�0w�'��}��=� ߮�BN�Oji�y�v�ޞ���Ғ�X�{u��D1kx.��a�WV	SH��\3��8����	fhPH�[����FV��XLu���ä�^Ê�(dۙ����Ԝe�uCJe�玔��u_�$�����^�#�EZ&b����%�{E���a�a�bp�2]���!�VP�t�<7�y�I����e�&��^����[' ��rCo3��ͭ�_c�/�C�GJz�hwua#-\�t������`�����pѸ�.�\sd�Lg&!���
0İ�b�(vB4���ѡ+������b֌w�YP0�I�*b�.D�P�����	[ؗ��?�� ���˗"�!���PG�G7(cr��Ԫ��2�fY��b�7suq�8�����b�wt��1mݷ&5�ie�-���
��+��3t�G��n�-,1-�ciZ&[.V�7�&����ۛ���K�I�9Q�q��[r�L��[J.�2[�\kL]�)�3w&��7J%ƀ�Eci����Ա�����ֵ��*���&*�cw6�l̹�15�j(�mQ�����f-E����jE�KS6�i�qۘa�,R���(¥1��cQv�mZ"�m4J8��[& �iP���e�K�[F����D�i����F���Qu1���S)��nn�Cmݱqm6���06�p�\j�փimV�̡��b�V��swwV�e.�i�a���YSPU7n���2��-��u������Һ����a�P�V��AG[����,1��´B�bf�cb�ڶV����0I�&9鸿�s�!�;n�""�����x��ޫ�l9�DҒ÷3�+j!�NW:{9��JpE-�>�/�;}?)��=�}E���3����z��Q<$@�E�lH����"z���MEcx���
����:e@=a;8��{�N��3	�q����^�PɤK���^��#���%�"��5!�%n�;V����t(���p�#���˺��F���]�FO��>�kT��Î�=e��$���[B@�'"�#7'��\�b�Y*��X����^��zʇfbҚ��pY�ڋ����j�^�sH��3BH����[5�וE~??���5�(*���C~�cd��߶QQ�y���h������-�d��8�wR6�nF�ol�]6�j&̣���Rf��������^K�>�U27)D��N,p=F����6�Me�i�5��Q�
p"�v����u��#�l��ddH��a�k�yG��!bW<�\�eV�a�D�C�B�\t�͵&2KDJq>�8i��9xdWU9�y�i��\���_u���s�t�_G����+�����F{j�t�Ct;mJDs�ܑ*�vi�L��6�~U�g��	�uoՏ�|�ڀ�ߎ���fRj�D^�~9ZmKT�+N��|ގ.�U�e(�`g�A��&�nlޡ�����Y�h���!�!-ϜcQ5&��1TЮ������[�1��p��9 ���}V�
uB��p�x�FOR��{k�5Y99�Q�pS�[̓Z,Ķ��0t���{*�!(t�P��H�Už��*$�p5.�2�P�"XN�K�6}��9;;eI؝�����A�����f��{�b�1X�u�7��W��ڞ����u�Oޤ��4��-M¶-�e������G
u�﹈��7:��Ё|�^��P���P�<8TuΜ�����^)<u��hU��M��Z$�F8� ;��ݝ��u\��Ltd�G��b����X�;��z����Cs����F�EgH�)���U�P��I4hfŜ����WXڞ��X����Ip�_W�����)`tN�DW�{4����*�N/s��ZE;YV=��
Q��侂�5���?=v�*�ב&��MmȖ��9��˸�)lJ��h��A�{��Tb�Y�E�����J�5�c�:���nJ5p>w�r��N��xF`�T^�	��cޥ�U�۽�n��3��[�VD1Rvx3�δ�L�TJ���Xe-��Zt�n�pWEL�!p6i��������@ƕ^��ң��xTP@�.����ǭ��[\Ў����(�2�ۃ�"���*��������J����N�hVXr^�wP�>�}��g��*�� 4���.*���p���Y�EE^�%����Ȳ��	�\�g!Ģ �T`%�� ��=�|}����΀ٛ�ml����E:u�b��gƔ�s*�64�! ;�bOs�g�sL)w�1M�������g*��pd:��̡�BӯM��H�L�}!EQ�OU�ا���-�SQ�n��NZ5c�o��~�"�[*����%����묽��hGR�	����y܌)��e���nF��E.�D�.Gh*2r)X����u�aEl�����Q�cR���ޟ:
n'{��Uzj.2<��`lPȨ&�6]������u4��v�Z����}�����)3���58u�s	�ytn�n�}S�'�\ܶ�7��Z
���EY�d)ê�s�;|�k+0�|g-c��[ǖ>�C����
��ճ�p�N~ӏJRz���>��c���(�N�2"NY{�-`�)ԡ}��fC��[�����E��YG��M[Q����}��"����"i�3����k#4�2U�:]a51�XT����è���(4x*���-/�Є8�J�{�>�r���v�;��kK��"LJ�4��'l{i���!�j��RZ<�.8`��O�u�����Ƀ7E�y�bj#�,i�TbR���"��G�r�' �&jtvN#���sq�#����;]�:�Hl��*M�&��$p1�H$^�-3{�FHڕ8e?Z5-__�hR��iC�&�������ǪT�"��Pk!�
�9�VŽ[�����"!8�dFK�a��(����zd�ʊST�4�b^��[�Z�c�M���q� �e(�B��[��3��z�)�����ދ��n���'���|xAV�o�1/���B޻�E����][�ɔ�A���
�m�v�Qm	��f�G��VE7<x1X/Λ�«�x.�=o��L�7��{j�r#`�Q�t
�t�j��:bV�:��4�<�㯆�@��Nu �f��؂Ʒ�9<9�P�4G�bm	�蛧�3���4��\R��]�K� �����ON���H��gk[�aJj�<��T���cW�Dog��lz���<]	�%M�nE ���z����NZ���`��I��P���g�#�ܸv�"x�UգN룲]wR�uQ���y��.9����|E����Q�E�\!���V���ƭ+e�7���O?��μ��Ө�+��a�9U�E�'֦��˫��q�B�qk�*��v�/R��OV����u�N�?�O	x1���yԺ5�pQ�1X��ob&���
�e#��L���)�W�EKp�i�����_�f�K�a�����7Y�M��:\�F���4���Ga	AN��P� DT!;=1�$qX�� z7��}�|��]*:ˇCvˍ�/Ȏ�!l	
���[:�&��w0ƥ���WOED�:8Q�jïl����*�����ߛ��RYT���J����V��4�Dk8�	"dFϤq�[9e��uA�M��\�����|�o�1֮�q�5� \�*ė|�穊���ps�t��{�s�+r�	�$�ȳ�+�[}]%��Jת(vz��qr�_����.��|?�X+����{e���3N���7I�eIS�EX[:V��g~�z�����Xt*���FG�h䐅i����N�V/
a���U���|�Q�Hn�A����Ɯ�ڪ�)PR�1*,q�;��b���<M���0�p4O�j�˵���]#�)b�%�ЌC��XB����{��oe{4�_%��r�{���/����"Y�b����a�jLd�jERq^�:i�Ҥ$��i�}��-��P�
%�Vf7�5X�r��n|���9^d^m�����-M>O_��J~�@1L�\��������ٸT:e��'�Q��y�&��ƱF.��`��8��^�^���BV:B(@Q���<zOV���#ˢ�S�AUNf�γ�h�:�m5�ߕA��U�Pe,���qp�k!�;i��Yeǣ9��8�/6?�W]5W�RxH��Є�V
����z/Gt2��������������Ѱ��+�:O��
��ӘL��L���9�MK�k�MEPݽ�;��d��Q֟'�K�}�����{:���P��㋔�wE�u�.XU��p+�bZ�@�Kd;C�Cκ��}a�-��|�A����wi��O �;8N´]%�frk�^M�k���A��kb��#;�q�� ���7ka9�e�Ltd�G��lW�":�A^�Z��!~ZG�'��L�.��yk��Ey��p9u�\���QQ�"��L0P�d
�*�Ʋ��`��k_�ǻ�dR"n��9�ֳn�V�.��K֩�����B������*5CU@�N�&������t�\���l���%i���W��\b4�>#J�*7$FE���\4�P�����Y�;�׷��#E�zdB�b3�W�q�*�D2�l��U�<�\��`4�#q��Q
�����.�����u�M�R�Ҩ�J��a�[��^��Ț>`�fC�Bl�G�ǌ7C�"ge��&8��O�[���Cz]�;�X�PMAT�1�p���ߕp�*]��`�@ge�0{P̋���^�NЪ���g*�|Řz}j�.���'X��`^>���v�p`���9^M�`��V%^2�Ѥ�t�8���*[U���C���6ވ��C�XF�\�_5���ݟ��˹�*Q8WV���d�P��g-S
w]N>8��[�t�Zi�CҩO��B�z��Ƭޏ�������L3�T~����Ӭ��u�7��
�h��A��6_��7�.վ�r3:��r�����`f��"F�]Xaq��H��R�Y�VI.w!�
�j��[�I=G�e�F���ؾ����T3}��ME��D�!>��
�IO�f^v����յ�c(����}V����>L�XV���o���N�<�_�ò��!R������R�_�1��x�#���)L3�{��"����W �{�Y�+���/L��)��)Av��(���"v=~'ap:2��XgK��˦v��O0y�{��M�W9S��J���y<����������1'��;��+3����ZG"��H����Y��DF��>�����3�����T,6'g��؍���!a��˻���ے"��P��&��'��#wz���X2s_0�@�.T�t9V�0{�V����h�M�l��ja���xJ�0��q\N���p�dTi5u�j���3���X�,A>9޽W:��^^cȢ��\��N��V,]�s�jlG��B�Ԇ�u��.�җLu<���)�e��Kփ�z;Y{ّ�ؓw��[z)��]}'Z��{�
�G���b���0Ȓa���9L�F J9%����!����� �>��O4�M �^��R2$Ë��
�+��������G޸�r^_N��ܞ��b�U�v�@l#�^W��5�V�������]E�;H�$�賑�^gc�ad@���mr�f�(��j�
�s�*E������V@ ���u��옥��8��[�֚�p��8�.�"R��DI/����+d������aj/V#��տ`�L���S�0�*��/�m��ba�+8�(����Cn����׬b���D8�9F��dQ>�N���U1hu�����SEm�a��+��C+7y"���/����b��b�j��\��T|:�*�C�����
,�Ν5|��x�k,T�X�a�؞��૝�p:�S�����������]t�!����;��&�:ES�Ȯ=��G{޺U?���ٛM1�����ˆg�_�`�p�u��/����k�|�Y�R�z�sy����,c�fr�-C�i��\�x����U}�Þ���;b8��W �B��=����Q�0�ѹ��U���X�S�>�1Ev�b]�Q\h����sk����sX}�Y��
�V�Xdv�##���*: D\!s&M-.2�]؆�Q�lW����À>�u��)�q�B��@!H���@�O����^��h�#�OD|jO��]N*�2:/�r��{4�;���A�+G�)� >�&M���5��<@�� ���u�a�=La��H,�a�
)�a�8�C��1�2^Y+j|��Rq>����d���:�}_�s|�ϯ���=�!����0�E���aP�s:q�Y�J��Q0*|��T=�'�_�
�Xyy�O�T��{T�:��Qa��'��q��:����:�9��ߺ��o/�$��p7!��$u����qRT��sE��*b(}�Rq
Ɍ�������}��,�>eA@QN2t~�:O�*MB�]���E�G��/����7�]`���[hE�;zd���Öc+%2}����
~@�i�>VjA�â���VT*>�0;k+1�s���R���XT�B��hgV0�Y��AC`x�V+ӝ��&��7w���2=�@P���k��$��yf��'y�@�۬+
�d�)������8���UH)��18��8����t�a�51��ɉ��}̕:@Q@|������w���w������b��c�ݒ�g����I'E��yd����aS��c���0�QORc
¡�~��x��ě�gH
/��Ā*� �>_D�
ug��DO��yHV''���I�*B�?$��NҢ��bv��:�3�T����æ�$d�Y��E����S�1'HVO��g1������.{�#���٪��],u�Ó&2��T᧥�w�2t���;��h���J���E�n]I��!��r"��y07L�1�Ɖ;�Ք�kuӰ�.�ݍ���J�%G�u��fJ�{�����m�zl���ӝ�k.�8K]����ܔc��}�!w[���fܚ�Y��m�&Qv��ol]Y�H4�';�O��n����듬;4r�mh��wKD3���Z�B�Ov��
��JGmZ����R��w7�8z�j��,�/%��[�>Fʝ�ic�%�c��A�b�B��Y&t��z7r<gc1�=�-�cG���%%0L$Pt)�[tTTz�(лG |0���y#t���J�}�͊8f�i�HH�8���j�Lf'��st�G;WZK���	�&Y*���1�Wj�hӗ�ܾ�J� �V-ƕ�L4�wz�ˠ$%��hT�}wYK��U���<�]pa,�)I-b��Q�ƎS���E`�΄/m��~_����3;}<*R8��oW,'�S�xtGZQw#}9�׺6W�E��u����_Wa�Dm�waGSüj��W7Y'U��,Y��ĕ�B�%Ӹ�g5|�wd���37!�]V(����m�L���{�S	ݶv��wd�sm0�J�<�ͻ�}V���[+v���ޣ �6g��}]d��ޛ��%�ʕm@�Ѭ�[r��8�vjk`n���G�Nv�]�[\�1yݢ���e�o@"�F����f���v���G��Kq�]>"*�|9�\q"�h��:�s�*#Z�3X4�k{��{�&���A��o��ӶR���w}sE	�)ZX�]Q�#y�;S��g`4��Р,��sG"�˸y�0����w�u*h�U�[�h��:[)�"V�j��
:c�P���w��vs�s,�lg;$g�j10)EA�3#����+���9@�+�B���h�����(���g$�5S��e� �]RU�����E�.���U4_ni�u�l[�⃃�S�)=��g�� �L�ϟf�A陛���7��m5�v��i��*k}��B;�Cy֦
+� �<-��,�=��,��n�B���)�*6�Z��Q?1,�
�t��/��Ѻ[��09)����MW�j|�vC˚[�P���I�o�\��O3�3&�Js��|jn�� ۼ��B���X�� LDM�/(�D���]��iw2��%j}�V+�����_A�\Rئ�7����w�B��	-H�B(X�Syj�߿�0w�^�ִm,��![C2WV�1��j����s*���)��
��s�6�Ҙ��
���*�+u�jnQjS.-���nL��U��U�1�]b���v��ۉS]͘.���r�L�eLVa��a��4k��VKw1�t��we�5�c��s*�ZR�YbE+T]hkZ��YivZ�Ɖit�TP��4i��D\�f.�Ql���T�T3rb�fe�
����q����h��H�ᕣ�1������˛�5��bkn5����rʅF�misnj]iSYD�6�SF�s!�Q+XWM�v�q�8��A��̰EM��wnb�2[��Mj\�s.m�Y����2�M��*5Im
���Mu55��f��K�3(Zښ0��]���F�Gm����Fj��fen:���1,p�e��,����ɍ̷0O��_�����*Ԃ�1�ܘ����W�c����5f<zr+NBUޢ�%��yRh�S�B��������=����ώ�� v�Y��O���E+�/I�'�:?}֘��HT�m��k����Ͱ�x�^2u�:ؤ��)>VT�ݞY9ՇʅI�h,�����s�Y�b1���3�"�^N_��v�C���=Xq�"�z���
���:q;d����*Mzu�i�g�N���՚��
Ι:�i��T��S�o}s9㸞~�^~����<Ag� rr����?3��� �_����;@QI����0�I�<������t���I��5�ydĝ�LE����,��O�V��K��YϿw�������瞗��1���p��M0+8�s����񁧛��
��=�v{@�ԅa�ζm'�*��Y�O\I�Q����c��s0_��"=a܈�q��Lx�U���[��C���Y⤮2TY;eO��Rz�d��2��&0�]H);}d������x�R|�l����>�8f9XW�MLg^��k=d�!�<�*�?�����/�%}��"�@��"$�YR�6åB��d��eg_P�}\OY�I��v���v��
3�c�zɈG���<b�@`}���[	o�s7�����8����s�32�Vb�e�Ag̞O�
����ܲ)�8�a}�+��߸t�R�cɨ
,�m�X|�C���`t����`eO�F�x�b�3r��;�G�ǆ$��d8�L�l���P�Xk
����3'I8�a�u���@�>aSg�Rc��Y�tm��(��TS�
�f}�+<9N�s�O�T���D�Vȯ�RޝԳ�#�#��L	�]�H)�'�<��?!R�:��Ӷ�I���@�+1Xs�
,��<>んRq
�_X�-��1�ɌĂ����>d�
)��=�o�zg���s��Er��ꉀ� c���'̟����kXW�N�;�c?2W���)?!���	8��w��C�Xj�^���`cY]��T:@QI��Ĭ�$��xw���B�����u'�Jf�7��?	s=�r��̓%f��<-���ݶܣ8��C�If^�>�9p�u��f��d��hZox@�9�ۛf_��|0�,�'.q7;*>X��ˠ��y,,,[҆���b���_f�f���{�ˆ�f����$a�O����
�P��L'1�TP�%q��u��Vq����cXVj~�uH,��_f�IURD��q����q��}�o)��VF���ew}�.�� �VcS^C,JÌ�<�O�ԃ�N�Ś�a�ړ�Vo�LO�H��T�,���T+M�f�a����+�c~���+JfzFe��.e���@�������
���iv�~�+�{C��I����OI�)���O��0_��oS�'I�r���& jV|���N'Y�}������x���ߓ�RT��Ns!�:�|Ɍ;q�T�ɟ{�Y��M�ۥd���gf��O̟���ëa�
�d��jAgl��NuE ��2`��|`y�J~�}����&�/�8G���ҳ���Xk���!�
(}�&'����Y��C�TYXT��<�&��Y1�2��i+��5���+8���ξ�a��e翹���|�9οpu�m ��p����*��SP*|��8�큞R�xϓ������Y�>L@_���SXc1>��v���=3앋:La��Ll c�Ͻ��毻&6V��_? X~aS�����|�aߝd7�(��w���W���'������Y5;@�4��wH?�~��v��Rt�{�d
ϒc�l���R�)Es�������ߵ��z#c�!@<K_(�þXbw:�b�g磼�j�&��MO�IR~C�7$����LN�Y�H,6{a���P?f`�̞8��_'�t�!�z�ӟY���������ܿ~��W_h�H,�'�鬞���e���NՕ�H��>����RN��eg������0���H=X|�G�#�<�p��}Y��«:I_��&3�nCQCĕ��=�I>B�zw�/_a
��r�'�H,�,��$��*<@��=�T��!]���:H(tyI���z=������7RK�wJTL�|�u۵@n�J%���㬳�%�z�%�~��~�4x*����j�#�~}o�%t�g�K�3�P����	s���9�� ��iS2�ʕ%.
��8\���+�	֍��J�k�|"�[����H@�����_��� �L:O�����1 ��̇LY�q�0�sr��+3���:H,+y�g�I�����E���r���'[Mg̕ �u�@������O}���g���9�^��y>C|�)9�a�2����u ��=q����jAO����=�\B�s�g(&0�P��H(*|}�*�Ԃ�Oh��RT��ɏ{cğ}����w����c�I�K����@�!���t�P>>I�'��S�I�O��'�y̟݇2{g�%V}@�!P��2�}ߜ����w��w���~eg�1!ə���a���!���솢ϘT�)�x��N2g�B��%u���"���f�C���+��{�3�Ne ��fg��x�@�TD��~wf5?d
@��<��+�A���XVz��R�VV�!���
k�ɨq8�$;���f��1:�8�g\�~�t�Xk7(�9@ğ!s�|��;�y5��&���h���r#� �WXp�p|�P>�c�
� W�l:CΩ�ͤ��2��hbAf$����'�:<,�u���C�i�@c��2���ǆ"��1���}��Ԃ���nO�%H,���bq���Z�2v�l�s�;a� �\��d������8�!�bN���'��ιHV½��v�$k�~��뫏Z�����F|=1Q�t	�{�����I�O�$H}����*�X{�:��!����Ă��o>�I�T�՞򕆢�0�
��H�<�p<" �1�F����O�w;�:I����'}{�+��P�t�̰:��풧*�C��T�4���=$�}��Ì�cӜ�H,�&'E� �5��0��ɨc=+c��6#d#��.Z_��O�c��Æ�����:����Aa���5>�~O?SXt��E���!ĕ�~�ɬ��hc��2o��I;C���}���fP�=�W;»�[�8�󿙋����i\�Ho`G�O��`F��:ߐ ���7vܗN���YO��h�:�'F7���N���4w:w�:�1s����*�s�
�sZWѧa��V^S�7�RKO}�! I�o]u߿{�w��P��Y�{��I�TR�f�x���N���P:La���$�nϕ%@S��$�*|�Jμ����-�����L<aP=���Y�%{�9��}��w:���g�I�)�&����I�?!S�ȽyHV��>Κ��bAJ�ɏ���1%N�(���y�R�B��P�<;�|�+8�0��1��Q�X��H~Ŋ�����n������Ρ��g�+<9�I�~I]OY����(�P��k^�1'�+�s�N���*�����'���z�S�+ݪAO�7�8�A�@S#lFJ�Tʾ��W��
<�L{�,Ă�a���E �y�l>f!�z�0��r�%b�OY�S����]�/�&�(����a���$�ΰ5�L/�Y:۬?0�q%w0�<؞����{7�˱	���8�G�` �`T��'�jN��X
�HVÙO't?!��3�}���N%E��fE=d����f��&3�R�a���,S�RT���򜺾����p���'�����a�5��[gY5�T����������'�<}@ğ!S��,8�R���,��N���q��2nQN}��� ���v�͚�}"��ە����p<>Y8}c�T*B�Ʋ��c;6�H)�7���z�@�gV0�Y�
�u`b$���g2N�P���{~@Ğ��k8��n���X����0��v�qt|2XQ�T����Mg̕1�Y�*�AO�7� ���u�a�=La��bAf���@QHo3a�bN!���ɜ�V,�>{�T:H)8��ީ��+��9�Nf�g�ǧ��0 �y} [���1�|�0�h���}���T1�G�Μ`Vq��V�E����bLIP�,�~�>�+�uy�O�T���OIĨ����γ߽����߳�����_܆'����~NuMH>P:L�}a���a��⤩9�1OSC�ۂ��VLe�O�²t���i1 ��nPPS���f�8 � ��i�i��=�_���y�z�������#[�WJY2��{o���:�f��m:U���P��\r��\o
�:�9��p�x�s�/���;�.	�;��Ҭ;{\Ɯ��p��814��m(�pB�.C3WNH�Hj����{� oQ�[�����zꐨՆ>�t���++%~d�S��0���(�+1 �`�aͰ�P=��kƲ�΃��5����°�8�I��3�b,pe�+�NVY��[�>��@�y|öL@QC�i1׈����5�d�>��u�aY���|�YY*q�{f�����ܚ�AgHvs�B���}dĂ�M�:���w�0��<�w�����J� (�|�1���:N�ǇVyd�Y�t����_�+7�& /ma�*s�|a��X_����k
¡�o�k�f$Ӝ��@��<����n�K
��� ��|ĝ!�a��d7)
ä����=B�:��?$��O���ɉ�'�0�w�� �@뾰�9a�Y*V|�+<;��Y8ʜE:�CRv�d���>���u]��G�I�67���zc¢��1��M@QJß~�zL@�?!���=��
�m��k������c<d�̝�pR
v��za>VT��yd�V*&~���9����u����ﾯ�������)��As��q�I;B�߹�z��E����$+�����S�>¤קP1���5��;ϲO���V\{�3����:�M1Ay���;|�߽^��T����Xj|��� x��!X|�&z �S��l>N�Rw���0�I�<����~�V.�w���� ��QC��1&%��1�`_�ޥu����z��5��7�v�a��9��5��*w�&�0+>C�������������r��@�ԅ`޲m'�*���Y�O\I�Q�����g-�*A����S/�Ղ��KP[����ǀ��bVt�+ɶLE����;�����þd�g1��~q ���&�(�����S�I��:��z��9HZ�z½�jc3|ܽ~����wߜ~.rO�%q���AORu���=VT�������P��l�������0:@Q`oW�z�z�{<�3��b)��H(~g��5�>~�
�k{�m�2��%JY�r���z�C�}�8�̺��KD�Z+-�\2Ի ���b}/�/!z���q�'���1T�e��lv]��_e�L�[×w1P�-�{9���R�G�M�=�3�������{�����6����ߍ��ԕ�������t�̛��y���=aY�o߲^��2t}�T�U ���dS�q���!X|λ��
Aw�k���:�$���q��8*E$��YOX�wY*|�z��bAxw�C�:g{d�;�}����L�ó����B��9��P+�T��)1����:�@Q}dܢ��T���ۤh�1�F�������E����( ����c<I�ğ%��H)�'�=�ǈT���>��;aͰĝ���t���:����%eO��I�8�@�}�<]����B��+�տ�c�B��Z2��=f��R��\�1j^���7�}릵q��;Q�M�V@�$B-Ed�n=�+&!�{��U�te�ӭzm҇��8��tv4�Ck`��(K3��1�F5Bj�R40��l|G��/�z�!<�a=��{��EL�E�L!c�l�y�AW��q�o��E:
��g �/7sv���l����Q�%�(A��Pͣ}&�1��\#�Z����͞ώ�'���w������!�k6C�Y��/��W��/��<#h�����)�ܬrl��k�*�:T6��G��jf��kR2.%@.�D�.Gh*W�ӹ�9ɳNpy�7{b�����8^D����C�15R5\�\$j�����Y��1����쭖t��#�EW#��1Kw%)f���=f���WQmu��[�婓gr��V�O�ńc�ҹER�̘�[Y��w�EbY�k����W����<w����h��%_?����EP��6s��W�q#����\����Ep^�BEÀ���0�Y�M9B6�����"jp�k��"��8��q��ԛQ����]�+UNb��t.�o�:��>C��ȩ�}�,t�i��}���:s=�t��;~J���@#�Z&v= ���i*㮩f=�J�5:�W�E����U�D&�S<�n_п��f�ЛIh�|g��W��^>]����Hک�rԅƽ�}���1A�ve�4"%l	��8#���n�`Ƥ�5�pCk�1�ˁ"����Xz�Q��;���P��BԨCe�'b߶m�\���(h�D0H�5="�#�9��6)X���j�m�dU��-Ϊ�1�7���	s�E �(:Lq	���T<��u\@����� �ܛ��,�j/\�C��	�)1�ї�	0������fGt�Y.=�� ��G���m�I\�R�>fl��o���%0��ַ����L�~����G���=�.��|�������Xcʶ�J!��=���.l��tyOM�S�`����:�3[�S�4G���ʅG:��W^����!mBJ�}�{���;7��31���Й�b= G"�Pj'"&�V�T�MFy�bO/=��аیf�oyD\O	jV���t�fu�;�C7�Q�2՘\⃊��y�����GF��A�����V=Y-�;�S��Ǉ��:U䩳mȢk���.qer���c��atv�~��V8�s�2��٨��.=�Yb��� ����]��c�ڗ'HM�%�)��	�!E��5�D��B+6z!���Z\^��s�{��2nGI��PRq��(�z{1�A��$Z�d'z�4�r��o�q~���E,O�A+y`Z��s��uZ�)l�4z϶�*�f��en�:�������[@a�W�L��7t���*[�cLg�j]?o���5�܋�OE���5������n�;V��%��L��-��V����Z�R�+�N�Pt�x��QU���E�Yp��Y����+�-᜾���*}�[�p��z�Oj�v��x�����m��g���¬xx+-*��m.�*-V��C�w�j]VQ��S��g"�Zk	��e��9zH:X�������{�x{�����䢕N��0���=p;/Ơ�pw]y��3�9�m��Tv�w��,�o�<�4r���J�B���RD�l�Y�[8,���cj�^�
�͊�,��St�n^�W���������A�'FT{aM%�<�yh�.�A��|����l�"��F�:ʩ���lJ}s�Q\B�ø��P��WVc\�tl�a7N/A�9���!��9�Ѹ�[>�1nyا$ۙ��m��dS�'�����9�.��Y�1�q��h��93q��Ĝ�Yy�o�Ez|�鸹7����Qfa��a1t�!tz�4;��'�����cQ1)	��wN@�6�Ǫ�)Sd\B&�p��L��UlE0s0ƙ�{���M̳1C�=��U�!NG
���_��Z�
��9�6km޵v�C2!���C�\itT'"��8&�G�k�DO/o�ܻ�֬Q[���D��v�X6z\q�#�� ��&X��� [��N��Z e�ɝ�Mn��A�9�k���-^p��m�V��_7%Iy\�Ym.�vs,��ΆN��K��(ꢣ�U�+�%� �{V]֮\�QB�t�d�9	�F�+��SXj�O�B�6ٳ	Hm2O��P�ǽ[գ��ۦT����Dh�_,҅{�I��Δ��\��LrԞ��u[ʌ�� ����eh5�\	q�V��ı^x�г,ۭ�]���b#���_����~��V���Q)ת;��fQ�i�˜���y���Q�9Qh�����29�\����x�`�Wɭ;�T6:���Ib1���!�Cde�W&ڑPU�T8С�(������P9��K���ʋ��-1:��0(���>پw�o90i�� ��
T��F ��e�1p��k�!�Tzaaخ8˾���tv	u��!�"�ȄɈ�܅���˓����|цb3Xz2���D�(:.����,F\(�/jg����mb�e�t�)���:�8�W��q�lT��aqH���	c߾盳g��]�����-*����2��E�pӵ{.°᮵O���r�]:Z
�"�7�by��[ǩ��8�j�2^�neNz�ݫ����Ưe��"���\�3K�^&��8wb]��wF�t�r����ܬ�Āj��[����'PXd�☖�>w	��>�s��\�A"w�^T-�k��MJnB��E��w6�\z�n�G4�nö�3�?�]�+$�>5e��>=)�Sx���J�t�5j������]2A�휱zQ8���0��Ž��RHǏu�V��Fz\VTz����39�oo���WJ�rZ��ժ�
 ��,�{J}cn�=F<s"�<D�]ѓ�Lt7����4�>�\9#rrc�|4Ѩ� �աX�aʘ��p2֑ǂ�4�ϠN�"��!�m��60T�ۺ�a�S��cUǫ%��l�9X�#x�ү�\��9o^�uɆc�}*Qwz&�r.U�wk��3(E^q{,�.F�ѳ%X��ۚCt�4�vN��Ꮀ�j�3��e��5V�S����8h�;�M���p	\����p��
�EX<爫oP�༛�ͽ*�:�u��cM����b��r=F�!di���k\i��2�S��W���O��x�=7ک�ѧϦ!~a�C2MFg��'\e����aQh�3�@q-9:]��zBŊN3.��ӓ:˙ �u��a�=#5�r�m\�M���N�N��T�f��N��Z�e7e*�)��X��Â@��V�4�0藱�SyY�i��
*u�n��ɇm��'C�^�q�ץA�ˢuԠ�󵉰T�gM�B�=V�C����*ȵEF�wcd����j�
v���g)Muf����C���w;l]���M����2���J����*�E���= �<Ú�6��͗��V�6Ճ���1���i��IMQ��#]C7e���xP�
nh��#�ҫ�<ک�;^�¶���b3�IBf��X�zq
�5��)xՇ��*�r�O�����ɥ��f�� {��龷H�Ѵ,:�͵]u�݋PF�Iٹ��J� �N��Yo0s*�ƕr�}b�Ț�>o�Bj���9��q�Vvrٮ�&��qiK�\ �OH"պ���Q��`���;�zI����td��� �{�o'"iqp��k�i�K�";7B��,��D����.�5pa�'|�X��u!m�׋��.;�����cWS���Gr�!\�U̕�!�$��IY�pk.s��<ΰ.f�:eY��J*�n97J�YE�b�V�s7nEƪKV�c��ICiUE�D����r�b3Xc�5��Um��f�c�jZU�E�j�nت��M�Cne۹���u��i�aq-w&�+�.e�ۙ���l�Q���E�Ըv���9U��rZ����th�̹�lݹ*��s26�v�r�ۑ�����
�ۉ��m+��()]qr�\��w7��1X뙙(�q.B�u1�J�����[��#��;�eʴʡL���]M]Gi�m��n7[��L�����Aqk*�Z��۠ͺe��"im�1u���W\��s3)[V�r�DL��S7Eܷ.;����[�b�55�j��V(;���mƦ�Up�Ļ���k�fS-ܣ��T���q�m&�v���7Mu�\ve��;�#.�\�R&9�[m��ˈ�J1nY\�\�-�29b��i�Wr�v�S&[�en����1.�e���#�f�T�faA��sp�k0�m�ZJ[1�7n]��Ҧ��x��bp��,[�\9��*9����$y�re�{]��)]�j��Z��rQ�+�b0��mh�[����xk��T�C"�_��\�����-ό�� d[���.��c���nbh�[�bܪ��G�jL	����!�i�u%�}�������詨���KR2'"��D}!)l�D�>����v�cZ��b]T�ږ:�{����뭺�����x�c+}Ν���(��<SQyu�N�n�kX�	���;���ʣK�GQp�������C/^�'q�E�7i*�o{x�j0�!>t5���٘0�Y�S(Fg���>��c����
�e��s����;:=�-Fv� VJ�1��V�L�h�7��hln� +J5�2�ٯ��w��%BGB�m�N'��bkMGIh�Q:<<* ������Pk7^��6.ϥ��@TT6��WƽΏ0F��si{
�Ҏݾz��Q��ӱC���w}�Ʒ������n^x��[|�q��eɭ5t+U�Y����	6�{xj����*���� �w.\A^�u۷���������%AO��i�nۏQ��geK�q��#V�)u_U�\��tʆ�a+Sh���\}�lpc�ou�Vt����<<=�������8G���tg M�,����؊�;ب.�ȡjT"7Qf��I�0fd���"4�H�5$L�HاR᳖F�+���K�q���t��H}I�W���Ωr�=��\��H�*����@�9"�~-]�<�o
�;}̣����ڦ!';&;ŏ
�H�,�m$<T�t�U���^a�p�%�=s�{G��z�S�y�L��l��<ո1B&��2ʺ����{g�#c
���1q0ӷb���L@S�!��'�9�2z�����(8��>y9;^\�zz��<���qӸ߃��nz.&=�b�t����2z]f��BW��Q��mE8�r��q�>�u�2ٿa�B+�rً�ȑ�8*�m�	�w;����,]U���Y5�D����$���&����ԡ��B2C�הD��A�ܐf�!��\U�&ie�Ц3�J���f�#*�*���oj�9�+�`�X���.�mVp�R��t�v�Ϳ��� �SϮ�@ǅ�*�7��.�����9n��cdJ�{1�V��e��b��>fK����&����iom$-�����ȸ�^>Y�"ԯb�:V������6�o�[Q�G�}�oZ�q���+�.�B��"�Y;5�s�z*$ˡ��w·u�v�=�c��v�g6Eu������*��`�(��R'��Nr$n����e�9B^J�i�Ġvk�u�B�\^����Y9H�}۹-���*��:]Z�yQ����R0����n/�Fs4������/����m�t766�*aI"	{y	�^�؆hI�/�t����$xwJ����W�鮢������pT�A�P�f,{பm
��YQS�~�>64��<Y�S]�nz��)�7�Y��ߑ�4�ρi�D8�����EnD=�KL2�2����s�+N�$b5-��*�"� �"���yWEkА\�WC?,�������;O@���#�:�޼��X/��ۑo�e�����D+1&5Vg0�*�و��ш����xsf� =��N�uf��|s޸i����/c�0��4��y>uuN��� �Q8Į������t�팞XP�N�˳\u�����Jq/�펤���/����9��n<�y�w:V�fusN���r�cۊ:��d����|�< `�n�0�]�?'�-LO����#b�?sA��|i�C�7ZP�]1A"M��J7*��?������q��{�~�cI���k&;�@1VtY�ϩSf�B(��ȩ�u���aXؠ܇#f|P���g���D:�G
��R=�%�|-gz�����w�_u*
�.�!�N�U�i�PQU5�/c8~{h�q�b���n]����}X�鎸:F������Ƙ����9<.���)�o ~ L�1�w��ݾ���$Q�M�gl�v��ˊ�n���2��ِ�֢��Ю7{�`�a,"Ρ]�阱�k�:��>C�n�A��r8b�d��y;&p=t���U֔Ʌ;69ʃ^x+܏�94#D쨊��	��:D����3�;q]bj#��-�l�NT[8�'�0��@Uj5<R::�ފ2>�0�*�b~�ٝ�� ���\$
���^��*\�T�@B~���]����W4�Uh�ש)3+~��j��Xi�F�ō%wTV�du��F�YM�����#Z���|��\.�X���c��>|�-�+��(`��+�LS�� ��(wu��oM��u���H�V�6�~��ޓ���1�,!G�+kQ�e�qc�F�����&�%W/�ע%�	0D=�7V��_v��F`%���������Yf:V��:����zd@T�و�(D����gf!��ƙ�"4�8��\�o��U���0#�:�߹���>�/Rz�Vn,FQ�,*�QA��f��"�4kqH�x�s5m�u��Uƙ���=b��#(��b+�D��.�w����ӣ��mx���9%ڽHFI�,0f��� w9�\DTjL	jcK�eɨ��3E@��o�r2��zp�0�,_LB����͵"�:�DĎq;'\��Z�t�������Z&z��R�ηJ0��{L=օ�/�v�D������{�{R����+X/q��s�2e^�>��?{*��s+�j�I��Q]�Ҕ&�t�!��k�>� n�f�d�+g�NP�TC5�*�wm�:�n�aOs ��{�-��C}K�|ÍAt�a�Y;�1��F!�>���\�|gƛr婛y%��k��Gڂ�x��[�벻AF̼+�ѕ%��%Ԝ2��N�5�������e`�XcJ�C+E��Y���������N���̅�#��<�z\ő����d\{YU#E��}��F�"�=�Y�[�|�]�= �����tᣡL���Љq:0o�VEZ�X�Q8=�ǌ��v�ɽ��=29l�Ȕ_�K����5A�~sՑ)D���@��⾐���D���	�0�2�է��#�3���Ph���C_��xe�5�aG'!��\�J�W��(�M�Ί��٨5�`�8��-�+
���Tf��tc۸�B;0zyB]{E.��h
�o�i!��:�^�F�#��Gv�A�+*Sy��[��_T���x���qAҘ��#����8��S��L*����n�0{�E*��"G*�"�N�LDÁ�d|je~��WJ�R��\�'~���3ѧ��v�D�2�zc�b+�ND[� �q|FYB�ﵞ�3,�K�\�#���֬U��dW��#�C3�O@�!�\>���\V{ؔ�e��7͵8�fHdb��ʐ(�+��M.�^�]`��7ļ]����yӗc:.}��}��Yt.��ޞ `[������.CH�])��7{u�4��Lqd��ibp��;�e�WÓ����+���[�F�E�y_��� /z�����B��a���{"�*|�1?y]C��� y}SΊ�~��"��$Gf��]������hZ2����c�|��}��C�^��A3�;��z�9��PX	�@��VM.#����l�	|l{��P�<:��Y�Yf9m�х�M��3���&ie�S��iV�(���G'�[Sky�x�g(��us���"ᄦ4֟'@*�����:އ:?��b�:����<�R�C(���՘�c7#�]#�������i�Ҡ����O��}ƊǸ󩦛R���x�{Y�2����VC����"D�Cwh+ҷ��#��ّ��a��rA�WU���W��FP�0u8���\_G����"�8+F�bx
�<� ���B�w�W��+���[B:K@�t�ܩ�J�ZkE�T�KJذ�C����-�F��Q��0��>�j�ChT��5�l�|q�+y�X6�x����weK�Yp��X��m�A��5E���hiW�����x=�*�^'l!I+j��d�w��9-���[Z���}v��cJ֖�B�+a�p*3��9���w�ɻ�6���1+�ԝk�{����ƣ�����}G .���]8���y�p@үs�_x0<�G*J��D���_>������e��;��	n�9T�1��"����%E�P���\��0��Ǩ`�wO@�S���;N��ldu��LE��lD�������sb�2�]Ё��?)�36D��Ї���'����. �*�J������u�}LU*�ӓ'��NB�B�شlR��h?���X��֔:�[���������VG�����U�o�O|m�!��?[��(��5NdT\�_%�!�2�l�=2��y'^�j��Q�d�6n�t
;��zi�#:��,]��jG@��b4<������4�&�6~�
F�������a�{�T�f�M@��������`��j�L����+����o�1�K����9],z�ԯM�4��n�����?u���}�Q`�i���R�%.���+B�L��.)����ԥk��[���!�{�<7Eq�ɥ����n���xV���q�H�m���}��I]Sz���z��0L�f,˹+��Ȫ�l0�G�\LN�ྲྀ�uFQ�'+��Tror�r�_xy�������r�P��xN�F�$8T,ȚS��_(�Թ���}�
���	p�=T���e�u���u0���p��g�Ҍ�sϠ4.��{1�Y8C욅c'���&�\Llq�QwTȮ�4C���.Nk��X�,�^v�蝀å^0Y�B���!bu�m��F�HR GD�Ɉ��n�>tvB�?��c{�����C���\\/Q����7�ܛ�\H���lmI�����lj]؂����Xz+��.����S�zM׶�*&\S�c/>��i�*��������0�C-���D����t�V����V��ͮjӔ7�� �*�7J\1*0#Z}D�3� ȩ��7��鱜j���L��D��N#��L�5�T�!�(��3�����x)���w�0�������1@���b��Pͳp%�"��a��d>�|H�[2��NF��O�P8��C��Bw��pre�*��aXqǃ2��UiJz,XzL$t��3��GÏxt�7��8�v�'�S.�e:�m|XC��d�tt��:�+dLш�ٖ���YHU%�O�U��ֺ��{����Ĺlrܡ�}S����}��b���}�O��͆�Q�^���C�Etc�ͼ���atn�rB��A�ˋ�M����ӆ��|r'��L�DY��P�{�� j����@�M��X*�1>��Y(E�Z1���7�!^*i���]ȱ�25�������$'��O��n�j�3���Qݶ��0*
����Z�\ �%]�����.�5��ş�UaЭ��VV��������i�\Li�ei��K�u�M��W%Z���~.���Sk_�w���X6�DԤ�Vk΋�\r<V]lMPl�sՑ+�D�'E��Ἐ���B�X�V��xE����g��ǣ��4���4W���W����r����[sG�8w"^v.a�5pa��O� `k����zg�Ǯ��c���
�J��sbbVe+ԡwB�N��%EyD�Fq�I1�6(:�_�2�Y�UZb�ޥ�JX��ǊY�Bc>|ƈ�M{;A�I�mh��<�,i�.��!�3����-��S 饘R����sge.���r��@�YIܣ��! gKcv�J�u���r�;9	b0�ڏh=��}%9z�������L>;�G=�.�X�ukD����Nu{Np�u9�]�`r�\����Y�t�[��d�*V��姂�ۆ�
��i�w���@1/L��U�?�&'Dm��,����Yj�}���²𱔎ֈ.��B��z���h�.tՒ_��^r�5`�SC�	kׇ���5EՕڭˮ�1k��� j�wi��#^�u}�NY8�q��'kׂ�%���.)�}�Jh����(#W�GX��p�1����� ��Vh���S��P��/3jZIp6�����w�
�c���;�Ǽ2=k���m����KƉ�88�S�}�&V�c�̲��冴ju&#2�&�9���dռ
�!��B�Dڝc����[;gg*P�V��Uٰ��b��)|4�r�#\�3Wl���M5�D�\;u�Mw��4y��C�Ur㧅�i��W�bukQ�}���ې^�>�׺k���wSbй�1�����`�.	r籪��ǃ�����Q�����hG+�ZU���;/��N�e�w�.]E�LyzD=:��g�eu�
"�6Yf��)hNܝ��a�m��0�"s����MЩ��ʕ��;3{�5��z���]CY����H(��'c����:��$�Y�ͩ��f��t�{m�gG!��������c(\�7��5/GsK(!��]��6�.�I��id���U�Y\�dZ��.�7.�$�R�Y�
[pGt�/&+����˝ձh�oT�uNs���:���(UԱt>���H����1wL"��'��y״�j�5�`��� �7f-�s;m��d���|$.��}BșJ���7��.y����Ju�!����|ӀwgL�$�G+=�f*��`�S�|��ǅ��kt*�����'s��
f��>3��Ֆ�1,��ޡ��$�v�"�ʗV�u}R�v�]/x�R�t|�!�gbž�M�Q�Q�n���C�;��}�Gv�o&E{��;���9z"�� �5�;u�DC�he�[�0�4�X|�c��Ê;��U�2ޭ���&�6n�0���N��BcW!�����3�pu�f%ծ'C�`\-t�9\p|�s��R��jj�ܶ�I�:(�d�5���.������7q׵%�PfJ��}��y��g�(��$P�\	D�2�Uٙ�bcJ�����eX��*��2�G�i+m1Ƣ�Ffeʪ��8�G2�W327*Y�\�ݖ�Y�f#��Sͦ\+5vԪ�Db����2�7+�B��Dk\.(ܕws5�Jڢ�������̹b"�53KJ"Ƣ�DwsjQ�\j�j:�ۍT*jVnn関+�Y�V(�[���.7)LJ娕�)l�v�nۃ�.R�µ�++�3��jj�K���QjQQGr��na��.f&���[Z��qEU��[Z�&aX���KK��mL����ʕ2ŅU�S-0�-�p��V[V����������70�F5���PS�kU�)�wK+bڨ��W+ejV�f3%��i�2��Uq��D�DK��	�
#iB㉕LeA�\*4�Lk1�r��m*�`�i�a��ܢ�B�#Tj�J��}i�	�N�W3/�&�Yǆ5�՘��O�$-�I�l�mr�� �8��:�c�*$�j�����o��c�y����u"���EA��y�!���/���^{�j�=y[�E�@�/�'b��L�"yU15��E�
�H�ss�!� ^mzo�>��V������Od��R?�*�2�zDs,E�"T��0dS�&�`��lM،}�f�"��^z�歛X�������㾣Q�c����XX"�s{
V>a���m��1�n�W�.�S�\�O�W�8��P���D�ؽ4,�ʘ�3e�*MQ������z�S����i{��(u�{�k���OC+�r��(
˧WM�����@h�L����N�P�<F̄��t*�N��E��l�C��}Q��G"���]�lc��-*:v��`27�Dj��{��Q��=#"��0�ǒЫ�zՌ�U9�kЂ��"�Y�//&���uʨ�MU��踨�>؟W:j�H9
-���@�S2�?{�_+���Fv�-53P���V�Xt�<�Cu�a��6�h-���֭�3�z��i���GƏC&��D�	p,Z2td�ʗ3�J��խQ6��q.]tm0�us��vk=7�g>	9�87x&vz������"�����F��^����J��%���QhB�.47v���[��1��	���'*�>�.Eq��Ms
�,H< O��B(IQN�?�/���iyi�ܕ�쐌���4c�K�S.6HP:��!PBtGW�΁�G��n�YXkў֜�`�kN\��3�Z���Fͳ^���JjT�p0+����*�wŚ���W�W�5�Ќ���9�;���uӌ����ɴD�����qQ�vyp�
d[��Cu"��Чx�Ce��;�T��Զ�\�~�u�U���� ��{[���s�d)����(x�ƈ�S�i�tkÈ�\��鈅�U�372�A�P|���
5�Y�t�x���'�!�]�-ʈ�,�^l�B�Moce�j��R�"1��Wu��,�[j�*R"��0ٽ��7D�ج��h¬��C���
S��1!���hV�~��v�7���Zx)�o^�뫏L�
��;�����C����x��ނ�=�K`l��դ��%�_J{�����#�櫊�YE{�a�����J\Vk�(��y�չx@\ٮ�f�Ǣ����ׁ��R�$�/95q-�K��=�蕛�M�\vi����CB�Y��s�mW�_
1#�2qv{����윺�C}]��Z���
!쀵���D�]W��>��6���u���򼵛�Ũ���.�L�l�U..�q���|��S6����q�{���p7�J��M�"b�TG0le������b��A���k��iǹȡSU7�"����\���
��^2���ȴ|��w����q��];�u9:R��x+܏��;V"�;*"�גcqpŲ�e���w��f�!�g��w����W��z�����*��Y��B<~{������B�J��]uz��9a�Q8Z;��I��T�D`* GEns��B��CdF���#`���r�x�$=~�$3�>F��|GHr�!׬�-WK[��'��H�a�r�������UE�LA���zư=���u�V5��v�8����q86��Z��t�snT����u䳇��}���y��v���j�!���)��sx�	�=��tǆX�ò]�.T�æ]s�1ά\�v�R�;S{�n=LM��u���&�hN_'���_}K��r7����������.#H4����{���:��踺��0�c@�Ӷ��=�,����'[&�K�ATR�F����dn�4CE��َ��s��"¨�,G�5^꤫WP����/��s�|���_c�[�B��LTnb>��ʷ{�p�/הѽa
 3� Os�f�����Ɨt]S��1�RC���
���α�y�^��$a�X��`���Rٶ�Q1U=�M1�y��DV�#!��Ԛ���ln� r��[>�c��x�bV{�cV�Q;�їK��z�b�3�D���Q�%&�}*����WM.�^����U� �|�DmDr�z᛬�ڡ�3j���Ĵ��^���+&�dK(G�^�N�=�Yi�}�i�Ã�ɨ�_8Q~������0�m�YLdm��o+5��=PӘ��gpҚ�F}��㼕h3�t5�8 ��"���{��n�T�~�=A�O[�X�I�K�ٓ����h�V��[�/N;�8�+t4uXV7k��k��;��bq�X{�S���%�WPW:���<m��hn�Co�E���x��W���w�d#-̼z��6i� =�ۇ5$X����&�h��"�WF���>�^��
��ٷ=Y�W���|>|�&�Jۛ��a���|Ab6�q�'����z+�R�go�ѿw��}~w� ��j�tl��X��3<elJ�>�>B4C%��ph�օf�g�Ǽpa�ۃ	k'GV\����2�B��B�*�\�M�%E c��Fq�"dFH�r\6`8щ�8/���|7F�ǹeV�X�|�X�j�08:�QA��|ۤ��܎��LFFT08�f�d���^�6i�}W�∸2�ta"���S�-��j�T��z�Xz�M����FϤY�[�ulUL���X�jr �j��YGL>�핓�^0���C���#$^҉��t6��vEi�zD3#X���0���	��F�+�������p� �m��+�I���~�p1�@��`��=Ѣ.�ㄆ̂��w�H�#���1x.����a������^񀎡T�O�Y��ʹ������u�� 8�<�EhɵWB��J�F���QL�<Y�>Y87�V��{��#��ͅ�}���˚hbT&9L�8�V�Q�/
�78���[i���T�e�3{��x5�Y��3
����s�:C�*�
]'*�PU@AJ��?2o���X����z�7�:�]7Q\ 0���������}a�Uȧ�c�������\�<v�����&/��~��:���E	C~x�i����e�:އ:?�4�6[nqq�ڵ���`ٛR�E�g�
���]�+5S�Q��轋��Ҩ�[ĉ�7ݪ57Jz�D�E�I`�8L�����@�@���t�kS�R��d�i*�t�XG28��N�9EIQ:ؾ>�>Zco�-؁��)kQ�S*:�]�s�W��WƠ�]�W>��#�K@�t�ܜbeUv���:�Զ�/U��2r5^�ٴhB�Fb�Ur�<�\; )SB'8�3�]u��w>C�pCO�������,��9/#�iJ�ρu�9M,���]��R�m��Y�^g֊���[.;�P�1���o+�"���!�.�ͯ'�h��W�{��i0J�X��,�ʐY�Y���H1m���!;w"��vh�'��/Bp���H=ԫӆ7X!.��D��j�1�m\N��b`�7I�Bt���X�s�=4{y��)�ptY�W0�o_�=� �6�kP�Ϣ#��G�8�S�W��^���b!��#`C#��%v��YY��ܡU5b3vr"K�>�U�
8S5� <x������Y�X�%��"_D@B��0��Ċ=�܁s:�D��֝�Q^�:j/�n�U0+@4iѦ�㔶{�}%�;kG���:b�ue*��Q&$y�����=H�tU�xm��I��O7ޛ�P���s����F@p��t�3	9�Dץ2y(+��3���fjCF��+�W!@�r�	��� �j�"%4:;IV8U�r(@ỳӀ�����h�;t���]Au�Uc�^�xtwb�>_���ڹu�]�b�O�K��_AK��;�׽I�t� ������x��d�t��l��Z{�6)(`AJw>��@���� l�B��٨�$8UfD�S�,vBys�]���!�=�|��讙�Vcc'f�jT{��}�\ֻ�t���ǘ[�a�]� �)�<�b�:���ڈ�(.N�����A��c��mnm��`o|ͺD�Ou :�`��������^޾����vA����tA�[9GM����#Zlu��E�QY���G�]�)LK���ۅ�7�0To�_Ve�^���y-�QL��������A]�j}"Ճ��5���;����
�ӯT�g-�Q��ش���PZ� ˬ�;o^�K�_C�������KU;��1���$2��k�x����F���9���Ѽ
����U��m�:&��0xg���A/�}fhk/'�z���l0��XPثR�ȋ�V�b+���&������6>��4����μ��X�)�ت��7`�i�ɺR��
��P֟Q0́� ��%�1z^�kwc�Dd	���z)"ޡ:X��L6b(5�-S�`�GlT��kr� ���(�+��X�M�a��$w:�l3p$5&�<�^�^�\^x��1��(m	~��p[�o�fu���+�Md���c�B�>�������:7+1jU�G��lNɤk䫛\,n?z�eD�ʰ���c,c����T3
̽ƺ)�G+d*�OA�������"�ţ�;���{<�I{�n��&�xGfrF�����X �,���ݘ�;{E��|���LJot���ç�z��n�!���-\��>���^����RXͅ�}�EK���T&}79���܌��#0�bld�ti醺��a^��sq9ʆ^*�5Dd"u!>�|+���ٺ��8W�01�{v�m��c:����a�z�S�2k�u��,v4^
]闣���*���M�JU�7�y��`�d�Z�|;��U�˯z�'���ج��Hti8枰�,�����OC���-N�i�9+=u�5A�a�VD��{^��u�D��Y�5���2d��L�zi�E{�&��*����w��NUrl�U9�{��A��Ө�K���)�о�5���q��k/\!sW:�:�KmX��
ȴT��`�����@T��HEX*���h��|q�Gq~�6+�|��ƥ4�}l�y�R��qA�
c���H�̎�z˹�]�$}��� >4d��S�6G)�#<Ӯ�j	�0�dj�N7���PK�&��$�"�HM�q� ʻΟUAs�2�篯nč
@�Uv��o%k���Sy�!Fۀ��:�����Ieu��+���B����{s�S�+�ùǯ�#�Vν�%�+�SK�������x���L#�J�н��>�fn�V�T��̱��w7^H�����;���\��PB�zQ�#$[�{j�X.ȭ1�����?�.�EF����G�mh�:=E�W(��ȧ3�j�[�QXe�`a��$����t�;�q��T}X��n�:#��>��D���p�@�U깖̩�b���{�0;��|�F�F��k|EŁC^�p��2gJ
���Na�m,����<�u��w���jP�=Ck����/�:���NvU�+6֩�I�瘣�:0uw�Ҥ��!�����b.-e�O��*�����'���^����r��iۭҥ/N��c�z���K��Y�00������OhT���٪Hd
�;K�TNf�=��R��p���r�0�C�p{�Ġ��[\]��@Ս,�Y>\��":P�p:��i,6t\�����T� S��������Vu��~�����UD��{jE���P�DvXoTҌ�Hs{B�8l���)��gX-r�J�A�2ʆ���컓�Ηb�*A�d�@�
ף�+Y6ڷj�[{&]
��f�=�m��L�w��:Z&��6E#aH�� h��E0�ȩ��0��M��)Pmh��Ꭷrz�����9k�s$5n�k��2���ggCk�O��M㸌w�}ʭ<�Q��
|��#6»����U�dɊ�O	y|�S�
B��g�W@G�SMem�|���͎Z�3��Ŧ!�� O��ݫuh�]LU���<a�l��l�-�N�D��RX����gb�׹m]�{���,��V�n�m�๞g�8]���h���Sx!��fsR�����vK�V���6���3e�/(�`�q!����˴�`]e��%�K!�dFCO���t�bMĨ\{������A��e�c�Y���&��^��J��o2 ef�I\��;��.ݸ�E��`g1�zkm�m|ql����[q��
F�.���7q��Mܽ�ͦ�Y`V�U��.闽se�j
p���w���5Z*ry���v�
��"��Ή'�E�ۈ��8Cj=���=���幀��@���ߪ�99}��98��+f^M7YN�,NCn�����̚���E��.�1�nL��)�E�]��`%�}m��@j�t�ȃ���ڎ>ǖz]E��C�ӷz��E	!���6�oG`A9��"��h5�:Ӳ�V�匁:,a������cA��c��զ�w�yB�-�R<���>�Ymɛ+�c�f��{س��{:de]�8���a������\��Y|�����_�Ѭ+7����Ւ�-�k@z
z���wsڕ�>��X>"l�I�cEd�d�;��C=��A[���NSY�"��VMM �C�4��8���k�i�K`�խ�����%MKx���5�[L7xi����R�'Zԯ��sM}5���x�[��̫�1+G�h�N.7�1V/u�U(F���XR�wc�ǃtn�PУ[�]Èط�S�/�,z�v�c��cE���w��i��Dɻ}�#|3��źC�i[:z��k�5�f�a.�N��DEi��f�����ȩuj���-㍷�5̹+K���>�D�I���[��+3mT�OI��cj�Ugf�xQFl}��d=���VV5�����%Օݙ�f��*q�����\�\�͕k�`)�Nb���d6f�7��~��^y�S�"�x����Yi`���L����A�1�.1E�ԣ-���a�̙�Y�u(��Ը�c���9q�\j�k����2��n�`c\��iWr�li
��r��]��[�m5��SV���nY�Q[Dhʮ��E�r�1�̥u��7n�0h�6��
�KL�7i5�2UsfZ��e7�q�E�A�bMm�DF��7vE7)\��a���2���]n�±A�n"\��n��B��PX��E�.�G�"�a��U��U��*nQF[�Ԯ3�b��L�,ƈ��n,t)Z�����R��ɹr*մ[�wv�m�S7r1����7nn��M���M-�U���8�i�Ѫ�0��(�̣3[�S��v떅���Wi��4k1%s)���]ˍE���5�Ѭl�+M���k���cK��)�M�ܴGj�6�V��]Ҏ���KeE�՝n�]������mk�����*�5�#��3��m��d��@���_Kř�����rs]��R�;-���^�w�y����йZ�C��m˜�v�FG�O�쐨��^��O�[PS�1Y��R��xJ���$�j�gmTtb�b^�㖄tٞ#��������_8y�=ܚ�<��g@
TƐ�-��\�ki�4���>�2�E�*S9GN3��*�&�O���,���m<AltDÏ8ٙq#OEP�Q�ˁ��F��Ku�|����~�KR�ݴ�0����DAb�P�|��*[�A�S`i�thq/f���F���m4��j�E�u���+f�H=��¸��<�s�>Z���wWzx\Wk!���(�3l�jLd��iлu���q~�p)��6�/	 ��dh'+6xa�\>҇��@yO0r��+�
��6��`VtÉ���9V�,)�/���WV�P1�8b�B��,�PIצ��D�>a7.�:1ە�����:z�]��>�!���HEEB�tPZ��D�]=�-����_P���_;j�Zȫ�}j1f�#��Iq�ք�MZ��;*`Rj��[��^���r0"�����>�j&K�-�+�����3^!��ϨZ�Z�������.N���!��9�� � ӕz���a}�_d�������3��uA��8}K�jI����"�۱�~ʐ2�[5�a#qp�c�K��Q`Ȏ�X��uU�~�a����T�`lM�I�U	�Vg"�-��������x2x��[�랜���0����W^�	~5Z�S�mjc(^�YT�.�d��E�,U.|�(��i�Q��t���;�J�p��;���=�~j���k%j����6��.^�vun&�?�;��3�^���%"*)�M�Ș�3�:�х[J�՘���0F�ca�O@�.��^�(�!E�G!N�M��TUj��'l�W��:�z�xD(��V #K�@����Vzf�K���w��-qD�L���Va��?L�5�� ���)Da�� �>��`��H�:��{��N𵉇ȫZю��׵�����
��|���pn���a��2ٖ���2��+w+�~��a��*�OE�7`�rK�.*�QA��D�	1��G����T+� ʔ�up�`�,��ZBsו8�[���ZvՠN���V��FGMF��jԜ�E|)\o����U�&j�@�w
����E(�N
��/k���byJ�V�U��I|=�����Z�� ~G#CؤlG�'����ux�l�Pj'�Z�ć�Nd�ByQݚ�-�7����>3�v�z�@dl���3��\�>����[ADӾ\����x�h�|��*Nu�z��**��x���(ϰ3��uWWouSYXy�����H�.��+���?z�`���l����<1����c��ЫƳ/ҕGG�BUR���ό`�%��7�w��;�Q�1����Mč�C1MY�;��Dϒ��W�@�6́Y5
�"b�_SM�D���
��F]e0��&�}NCر��7��W�^��h�oaհ$�}S�h����!����^Q��W��
�	��W��;�^G�c�sne�~�^�L�u�3��qgY�Z��G�
���Bi^�qb渦<��j�m�BAޑO��Y뗕��>�̽�'b2��/K'w��6E�zWh$��7��a�k,��_�ho�c��GwŒkN��tޅG�M�3����b�X}YJ�k[RQy`��J��@�w�*s3��	�β�\Ikij��B+�VJ���{�}�^��S9����/�]��!+�e*{^!3X�	��N�h�Tg�sQ������}�Ѥ��6�^�R�H9�r8���Ñ؞���dO0�k�V�9}/8%L�rF�P�41D�4ޡ�n'���S0�}�ۯf:v+fKs�Xi���0�h�m�v\�X�Y�Rgq�N�ѳ6u�2"9�Q�\�u�����w2�CO!WӖ�p�SfEe)�����΢���5��9��h׮,�o�k�;n�7�v�����I���i��9�
�	�\$�PK�w���BG�����)�����QＭ8�������m���V�����6u*���:t2K=���է5�fS�Ou/b��5u��S4��f��n�v�9���ۻ�;�!m;!�}6���qs˜��vRW�*9��ۊ�0�
Mr�ъu�ZΘ)��Ǒ�+���謕�0U�+<�b�Wv�gN)���x��-���4���a��4�[z�P�K8��{�۽[����Q��T�ĲJ��^�"���ys��5=�~[�'`h;雽B��oSU:��1=k�����Nl�v�X���[y�E��X����i�O�i��G\D�8�Y�ϫ9�-\��>����Rq�L5Δ�v�<��0j�������&�0��G.��N"�q�8��%��N��G�V�����9(ڳ��u��1X�L��b��o�me�F�J�p�^�S6&jrk�3����,nƦِ#z\��XՊ���F*f��Hlű������R�Uf�P���	����3!����N8mc7��~�ܚ�6��p��&����NB�kAq]cx0��/k��(��}��g�2�ak�S�c"��Htٺ�S���bA��f��W�hؼ�4ӌ0�gb'gvlq��<S���߀r�ߤ���)��Y3F��,�kQ�P꽣G�Tת1�Y��ݵB���v5��t9�q'AT�7&7ݘ��ÓzN�e�h�C�s�z�B�����=�kq_&#'k�U��j1͵Zr���f��0+��1�ky���	�M��J83�A�smD`}!��\,�y����G���S�q��ޮ\8�>I�jc�kx�D���ʔ󹈭چd��X��YB�ecBFR������=�"v�Nv���U�e�NC轠5�9*���{�<2��ԯòV8f.�]L�_+J�A%uyY4��}�i	��ɵrz�.�7P���Q���i_6"���;�M,��}*���|�o!ׇf��THη0�a{�O)Eە�իǙ�M�L)6�\�K�\js۬���c��'m�;p0oD�ޮUz/iW�.�ջf�tl9�=�]7V�R��Z
�q����Ov������l�kk��-6�������֩.�).�=7��#-X�X����WӼ���>/7	�	cכ��A7˪��˧:�4�ީ.�{ZkP�<+���unV0j>gk��)���ܰM5��u�	RT=���r�!��/���n�5\�+�q���O�(㽎^u���{8h�{<��X�rp����_:"�ۉ{��`j4����+��z��=>��[o���[C�:���Bp�!��4����J�ىj�q��4�dL�ҭ~��H���R�#
�N-)N	��z�Z�WB)��g��*��q�:��د5d4�X⮐up�U䶻]	�v�M�ޣ"���oD!��:��<c�W�J�7�qŧ8��-��Ϯ�P�Jp��Sb��խ�:f�\s�_�mP�0�A��4�̮�f�]��|j̒�(���H�ͦ��f|��}UҢ���ر'�u髼�붚l��n"�`%�5=VF�W3ء �)���O���xb�W��H���@�ō�ق��S8�M�d�k��ڥ�VaG�
*g:�Г�
CO�{*�Zċ��w��엦<sjI��97���9�ԥֆ�;h���3:��ł�r���
��:�9�_W�^��y�?��̩��o��v�����yfąb�G]�J�ڋX�XZ;X&��=����ʮ��f�$P�'}A������ŬY��p��҅�푸ɡy��}ş���VE�2�dpggmk+sQB�u?"��G�Bp�6-zE>�����xAŃZ��x;�򳓈�2�N�>��o�萶�!�Ň'zkx�*��er�j"�,`V��tu��bvjңM�����Rv���L���X��8^��֯ջJ�L���%L�rAJ9¼��[�*rX�V-CEs2��nHb��r�V�7c��^i�49u潻�*os5B8Q�o��kѣfl6�v̂�8�K�{Q���P���!�Z�Szr��l�e)�c�Z�9j/�G���}FC׻z��i�-d�� �gr[�ĩ�.]v�Kr]ͱڣ�n����2�n)d�Oӏ(*�W2�Q:w�i�NAxf̛�	���CN@8�_'K����=�B�W$0�����;�gVE�#gV�~���_4�<'�б�%Z<�x�۹���"����磦d\��������`;�+C�䛠�I��&G8��}sm�5]��s)����!B��װ�r�ͳ�L�V��®���#ļP�`��{�.g��yr�V4'r:�Ʈ��)�wbV��\-�^r�L�ȹ�z�Y�J쮕�R(�E�6���U|�\��l�0�[`՜�w;=B��7Չf�ہ{�.+D��J�a��Ƶ���$S��9T�K�s����zu"��{8�{]�SB/X�Y��盶{.��aux����շ�u��c{��Q�ϟVK���ַԜ;)��[	p�yޑw��7�0_WX��lU&��m�NO ң��_�X�˕��%�2�6|2''�׬b�iE����ދ*�ٰ� ��h�o'+��4VR2�vi��8�>ɬ4}�$��U��̾�ִ�`���F勽�_l��3qed̅gk3���ۇo���Te�(I\�������[�l,����\ϣy��X��>��1S&\
ԅN��.��9��Ϣ_@hj��CžC�n�T�j������s��{{�!�%��EKH�P�
xb�C�WX�*&{���T�]���ᒘy2_H�LSO�	N$0F����e)�� en7'�S�șc�VoG}�t�9�j,�N�)�>��4�r�f��^Fn��,���S�-�҇z�w7MD>�q���S�}��\ݫ��5Q���o$]���s�)��8��i-:"w�������MVz�����#�n�P/+�Б����
���B��oy1)#�������R���t�7�.xecvs7��0wkR1״ó��Yx�&�O!yA�Y^;6�IS�8���$��x��x�;�[ݑ����`��v�U�O��.�<̅�Yau�GZ��*D��YP��ۧ�h�����T���ѝ���7t�S�p�'��w|۰;J�2���nJ\U7ܪqS�'�gT�A�[�쩝ʙ��dY��[m�{&�I�am�ٕ+iT���ֈ3+��׬�K`��L��֥
ݡRK�×�ua$}�㝻���%�ֈ��`b�\����L����uNp��G�ws.�S�D��m���Q8���K6:�JB�E`�)�-�Yb����ZjQf�+t�k�M�Ǒk @�F��bV:M뮺*��)Ou�H�g1��2ٝ�*���'a��jgN���Wr�n9E�o���mr�;-�ͫ��"�0t3]dŬ}�lJJ�#Ȫ4�8W<�9�����$�.`��HN����״�.ZVtx�3�h�5x	��J"Ӝ����W4N�L�ѵ���ҷ\=���;ut��N:]k@�S9����<��������ei����ˏ�;Bu9Fa!������WGn�CO�t^�+x�x����X"pfaP=�Q�ʼ/�*ҭܻ��Qq��+�l���enJ#�Nr��ha�٫)㆝�o�E��	������:*'6Û(�`�p�٢��:u���pWd�c��՞�,d��.�5\ X�R�wER�3�������[=Ȯ�����ZzqOP����k�����:�d.�u{e�X/m�����9t��j�b��%*�!�ڏ�GFS�"v�f9�ƯoM.m�8+�A������T�I�:c��;u�Zy\�K`������(E���C�v��}�%�-�ޫ����xN7$}x3㶫s| ���R�ղ���)�@k3�k���s���͹t�t�5e�cY�Fw&�;�r��{��z�#�Y��Ō��IuT��Id�ݺA��N��e��X�͠���ٌU�[���f�-���M�:�3��u�j�\�l����������.�7y��k_M��GE9[M�W4�;�U�W!xR|��/�e�hք�Ǎ�qVE�e*�HBe@6�X�	��]l�W�����D��GJ�b,<jLԭ˗�䣑����۳3�����o4�Q�Sd�҇�Z�9s�r���Z��$}�j���A����h|貦�@;����d5�W$B#�l�xut�ZhMm�}9�e��yx�;����I���N���ҁ�L�j����Zq٩��`yu80p�}-���E�k��v�-q�hj�9e��L���U>.1{�e����Y��a�g�PU9m����}�y�����`��>�GGw1X��ff\�B�Vbf4G2Ѵ�q�ZqY[p�0Ct�Ԭ�`��QnYX�es#L̘"1���nDmhc�8�l.4�E���SP۸n�ũi�1U�r���̕���i��e��Z1T�0��� &Zµ�2�R�e-HQX�l��u�tr�-�.a�X�1�jQ�L�@�\����mE�72�(�Q
8�fP̰�����%f�ְv�̦R�X�Yr�ⲥ*.
�d�V�Y�1�)�(�W.&,cZc*��¤��pmZ�P�egV�:�E�2�QI*�D+V+Jb-�0�m��LeclR��e�YY�2�#�V11��Xm����+����*b��&1-3
���b����b��
&1b�f�f�W.���X�m�.R�p`bU�2��
x1��s�s���	�k��F��ӻ8�\ǻ�Y�Eʆ� �W)�J���vr�ى�'�}�}Km���n"�
]��\��F�Y���U���9KXGi�uV���@
Dl��R��� e%��k��6�
M��o�����ة0���AhV���Ot���P���w6��7
��s�1;y��nJ�F� ��@��=�&VW����P���+�6T���bV����׶|�:�dw��L�����{�mm�E��F��_�鎂���F�*!� w����{kг�)�8�]�ջ"�d~�k3�X���=�T�<!J!'B��r��螝��ݨ.��^�ѳu�]{�a���<:%8�0�f��'�M;���1�R�C!���`r�C}5��-��Q�0n�
v�\�
6q��`ְ�\�9|k3�ѭ�vۭ	�}�H�\�b|r����J�;��c���b��dR��pyO#�s��=�y͈x_c,�F�y��Y�[DaSz�O�Nި�v�c��(V�u� I�ۋm݄�7B�7���5'u08t.�)9�O����ܭ���J,Ψ�Hk���j���Қ�r2�-�4s�"�/y�pK�7��%1/�L�1�=��Qo�u(d=��X���}�#oC����W*qFJ���
7��b�¢u�I�x1+�����躼c5-VF���k�D���º-e����ܯ���nT���k�����i��E��'+�݂8�_#P��b��\���6P{k���H��@�X��������M�8�)AZ�S4��Q;D/���8�bg����cn�i��e�6��5e(�^N�m�hF����APe�C������cc'm&5>�c��h�H[Hh",8�DmJ�ʅz&�\����ͺ���w�v�vk֕mć��j���s�3jw�ߏ��>�~�"F�`���OU��.n�;[����)���ԏ�^ݘ%t��51y�C�<�5&�oS��-�W�QkU�ppZ��s�+'^յ��7�,c�|�]��@��2��0���8�/�����y܃��$��W��s�*^���E�Ӣ(JQ}���[q���Al!��$p��1ӝ8|�;ۯˮ�s�k�y�?:��;�R{����ѳa���f�o�����ڶ�CH΍�Ƭ��Szr��p�Sfk)Mc�m��B����}�<�5#d��#��:j,�jg�k�gm��Mڼ��W�C��J"�rX8��s��t�I�>��q�2���g4ɾ�}(vk{+�:�tء�u2�]Q+Dm��ū]�%�j�,�6��x\���	���q��}Jd�j��u��{�̠hj�[cvV	ɚ{M��9�J�
����6X���m��X[ЬU�&��n�g��vi��J�Jik3=ghߺ5u^�n4_ڌ:ړ�O�D�#YOP���l�쀾,+N��b\���n#H�ɺ�1��p�r�\�W�Y�,q�����fQn�u)�}wks{{29�<'�
���OyƐRpX�6>O�ﾪ�ڛqw_=:k������&�.���&����
f�F�]�7��]�97ڏ����7���C�Cat�b�ܨ���^!�;-��2V��8��}j�/��B�[�䜹�-��hU}�P����]�Lm�U$��m���F�TQ���uHt�`Ʉ�ccz3���a�p���^���v(�i�>�^#�)Sŏ.�58�'����@CĆ7���Yٶ�����ľ:���*e�׻��O�*�}���>!�����'�k3�{ΚQ-O�{E)\��Df߽M;})ĩ���C|#a��[SS6���z,��*͕CO�^���QG<ӪS���{�P���Z�W��5�+Q��sY-�҄��b�n���ٮ�fn��M&���~��F��Ҳ�ZO��-����iem�En�6��:tVi�wo6�:������w;"����Zu��5���qh����:3EgN'���#+�ܣԵ�F�Fs�u�2�+���\�:���]]�����{@�㹼���m�d�9M�����Z�L��c%���!u7<���8�L��㎩]k2�s�3�
���{�#v�r���t�<��eQ��Z~��*�<h��?]<�k��罙��k5�s�+��r�ج��n䩋�-��ؔAqѻΒ��
�c��^�y����4�3yt����r�퇳O*�R�^��N���"�z�
.��[5�����&��/I{��~�-4��Z�|�G�m��$�Z��*ĺ�V��/-��:���P��M�'
ڙG<��NDԏ��K��fa����13t��c&m�Vy9-@Bע��eEG<�[/�� �5Z<��[�S2g(��b��u���J�mƽ��Ί�GQ}��y�Vw�k��/n�A�Z�C�6�]�2�N��X}���M���9Z/[�bY�ܖ)3�v�s�_�!�x:.��cfm��ɥ��(�n^��ǽ�r\��j�3��r)Z8[�˷{ƞ��I䟟}�U'g����dN���ݗ8׍=�T�<#U"��j8���rf�?�h�j~��V������-�FX�4�Д�z����uN���[Os3�o�`r�Cz8�c�ޛ�݃w�sx1�y[�0��-̶��Ѷ��(pl�1�M(}��(�^l&:C	��qE(<��f���-Ҝ/"&�y5ф�k9�
�a�3I6ч�q�3'��U�7+h�v�����\^�S�%<�>֌�])���v���R�
Ѝ��a�Z�1�XY�GEմ$f�+>�WB�\�v(HV�������zo�m�A`�]I�Nг�ICٱ��1�s������[K��3m���P�����q� ��%#n�����X�9��+;;���N�1$��9�X6[�e��� }gƋJ�ĺ6D;�vT�q�je3\����Dt��8�2��_qp����Ü_K��9�Tl��t'+�Nu��*
:;]�A�MJ�J�IOE�pY��X���Ⱥ��_{��ɍ㶇H��6$�i�%�=�����sn�ժ��GeSi���3�U��(q�c!�gzE>(�pIp��,�^^��&�N}Z��w}t�����7��-Ӽ1���.6��[˘�E�r*w�%A���]C�iI��H{M�*��nV�j����H��t۱[���S�	S4-: �
��S��4��i�P��5
Xޒ8뙇��ڬ�N�l�o���䡷��Z�q����]ta`�ͳK��ϖ#5�	!f!�s�,vE��qG�2��k
�|�'Ӗ�NSf�e)��mTfL9������,��j(�jyƽv���ȹDDp(�K��LGE��&��U�(P�Ϲ�I���}<�j��n�˅Xj�J�{S`�M�v{�uR�M�,lN:1�:|��&�!�:�G�0oA�!<�t�x��z��4��:e��u�>_).�款�ڜ��*�7��Y��������{��gI��srNS���V��ҝaB屃l�Lς�g˪&U�p:k��^�k���kD桘̛7�\�����McVYΙ�u�r(���,MfL����Y^�cvVzri�/����t�E�ODm-O�[m���g��r�r؛�rm���Y٦��ޗzo��s��Ew0�]n�R��zz���)�(�S�w���9tܬ�X��c	�c>������v�a�]��F��KcV�0�Ҟ&��΃�ޭ]eg{;db[^o�[/Q��'�ʹ��;�ւ��8!��X��{��u���*��&�Cs0�ۡ~旮W���;>WP�)B9��{���+���C�6�F�i(C��M�"|��N�!�A��R,C�j�YR�L^4T�v��s~�K*��O)X@��]�G�dn��֬��E������Jp�wr���KyJ�ѝ:��ьy�� k����75��{����[����[�������O�3�u��W
��ƆC��9V��s���6�����b��#�w�j#���N[���%��ux�h���9�A��ԧ�6.z'w��..:yjpƊae��y�U{n�u��G7ME���/\����b��c�7.��Ȭ�>�Jh��J��{����_lB�uvn�b�!���+�˺�I��2�g�NRҶ^��KE\{�W=K�9|�'����q�@7u�'ݬ���1�Oc���йȫ珙�z)S�r��{g�/VR���3���X7B����\�.��c5:Vw�f)��آ}�^Sb��ٷ��]V�)�-V��4zE-Y�L�A��I�fד�^�W��童�]-��ܵ��c&��U�����y���Z���Ӭ:�^ʕ�*t��ggd��3�wji�Uz�y��M��b�g�/�w{U3�,�����F��{˶XS:��n[�m�����������q�P�(�A�M�T�p;!��e����S����������D��Ё������9�;b|u	���J�s/iV%�z��ٿX"��.��T��˞��n!J��޷k`N~���W^����w���X���n���6���ԭFy+4�7Kv�<L�$��-Wc�f�u�#�o�:-*"�n$�;��o\Q�Ճ���z�����O8�T�[�+�k�Ohr�i�
Q'�M	�G]�Y�wb�4S	*�ְaZ1ˮِ[T�(4����a���;[��0ga�o�}�m*�Cn��o����mv�<�>��k���)��9j��O��"���n�����n�]9V�"���,������A(���>9n�&�n�P�J�l��J���Qz�c{�2�u�'τL�2eu�`6�U+��_E�g}��B�v�3tML���Qs��ݮ�Έԏ��fg!Q\;KS�+�Oea�e��>�n��4�t־��1�gY�fY�OmX���u\��rA��Ws�zu��f�\�5'q�F���.Zɥ�/����{�	�.�mWQ��f�W�zoN�mZ���-�5ݟYX����Nu��z.4_u_r��v>�񨁊�I;y]��$��Ҷ	k,㲃����l���o�f��V�u�	�1�t�qU�r8b�%a�na��Z�*ږ�T��Ec2}����7Q��ɛu��.��|��%t6���⡎ձ��L]JεL���m��Y�+yZ%�O*��aR�.�2����J�u�>�1��.n�3GbP��ĭ��w�=yl�,�c�kar;zշR�x��p(�������7n�����>���c��/fú�R�l��/0�psq��iWWf타�Χ*e-]��1"�ժ�K�s>t'<'�S@�ֹj+l"ho*�a�v9�{����R�j�A���[�f=m	�w�����v��kF�wR&.Y���k��LQ�;+s͸#M�&�np�y�7%oX���=0)[N�����s6�������r6���t����ݛ�4]�n��+�J6㻴����[ [�Ȃ�ӂ�Q���'�+6�Ǻ�m!�t)�.���i�un�t�+psθ�+��;S�L;r��ٖ�zn��׷N�^ؖ0[�F�+/��66�H.�e��8 '�^k�9W)˘�����;�sQV  ٷP��V��L���T����s[�-��`�CWͼ:�����:�!�i��Tޱ+����C��HW7{���s�2�� �:�efvlܐ�E���!��U�bV�c�.	��pک�%��`=�:H]+�����_`�u��������ۃ��'�{�i��8P%�B�C��+h*���{�e,w{�.ެ�]��:&�@�̳q<�pw83���C�^��"ƶB]�i�ǈ���Q�o8�U�Kr���k=z���3&_�b��ދ�_v�V�M�+!��I:iZ1��΅��%	-�+,�*�i}��=B��762�7���n+�s:l嘌m��EºSx�/��V�iv]�]K5b��	���gL�:6�t�,]���r�	����Ф�� �-���oyu��o�u6�4�h\�i�cF�����)�� ���.vԌ�w�Z��;���oph�;h��|��'{Ϝ����Rf�97��t�x2���58��c�Q*6��)Z�`���.��k�%���)(�J�V(,�̸�&U
ŬYe����0�f�2�r�b��Lb����[Z*�1�R�
".5ƨUm�m�����,v�Qrىq���ȳQ�
�Wr�c��TT[JA`��VT����T��jݵ��Fc
��1�)pJ��C\k+�9��-��as3
%u�5��QUr�9eFڈ��ZݥJ�m*,�2�s(�Eb�X[H�Yb(֮���T5ͳR#R��Y3*�)U�ȱE��M��XV]��b��(b(6�%C�(��h&aUIYr��Hܳ&�b6��"W2�ԋc��[Sm@[sҢ��m���51��ہ�,t��
�P�MEĮ�����C�r]��4���nP�l���᫠u�na��������9�|�ٳ��ݤuQJ$�:���Vv�����--�}F�=�K���9�yf��T�+#��Y_nKzT���w�X�\��J\������l�')������P����(�ૐ�����W��h9����>�KsNa�NCy����s�&����=b������tu��������ˈx�t�T����<�K�{O_��㶇H��6$sO�R]����N��wUom��d���sn:���D��H��bаw�����j�M���cX����m��.�v>��.��[!���;�x7�5P���o`���u�=��Z����Ru��H�$��[�8۶@��}��#/zS}�ݥb��{^J�ޓ'u{c�sE[��9���'�5@��3$p������IWԐi��p`>��m^WvV�'Y29�j!�ȕe�N�b�l5Q����S)�_�۞>�m��Dh9Bw�~���f8V�ݴ�L"*�;�ܮ<��J|��ڄT���j�\�]&��
R�Xb���{�97r���*�H��L��h!������6hS��*s��;�9�xd�e��O��+��>iĀ����s6D`Sg2�	P��q2�u*��X��s��2��zgm�<�ܵaÇ���0�[ܑJ\�ov�
���&騒��r��h�f۵ڂ��#�ᧂ��\�XP�t�ڽLʴS�.�[ݼ�%w��&��WG �Uxښo*��cBq=@�rQ��>i(=I�`������x-)Y93Og���A�	��qk,���Q{L8Է0r�����b�7@�ۿN�P���Mp�&��	�os���a�����S�=���5P��*���,ڷ'�5���u}�.���_�uS�m�Y�]���b��6rv��.`��ٻ���D�ߟݖ���ƭ$��*tm� C�P��n0�TYA]cX�k5[�yRo�Lԑ�uc��=N�����ٶ��Ǭ�H��{����2>�681ȷ��+:Nbdԫf�C
`��	ݚ}�2^�vφ%��.�e�l�a��99r���iC5)W��m1�V�I6�ٯ����af,�9�Y1�W��*���R�����γ�1�!�ʕ��D��}��H!�_�ݯgS+	P��j�ڍF���i�[n�7����mP�P��Si�@<�H���,�}�\�s��Ҭ=C�C�d��ئ�Qt��W!6}tC-�i��\άN3\�s3YJ�9X!��u���騳�`����ģ�n65��-���W"�3N��oF�'�>�"�LV븖mR�qn��S��@��>��Γ������P�A��[F8TT�D7}�r[(��漕�m	�Qn��c}/�n����䨚�(r��U�2L�Y|���VEj�Fojp�*X�L�و��	ggS��X�ዥX[�S��1�Ɩ:2<]�K|Ϊp�"��5� 8�T���Cq>y��_=���(�5�C�ŗ������p.tw+X��z�Eޏ����܅r���9EnQFNJ�7>HFo�yWMW$��)��FVk���+5��:�q^�z�����G�9y1�u�b%��8���g�qz�W9��A���g�z���#����׭�O�
����D�����ҫ��ѩ#5������7�n�B����.�#��!J�>��mw}�&�|��:.᜝�D����/.*��~�0R�}�q}����-�m�X-�j]���N�~���'f�t]�A��t���q�<Y2J7�x.k^Ѝ�G�_�����:�o�5iQۇ�,w�������7��a�eHY�m�ݥ:�{\�է�)D-���B]���q.�alf>���i�·��d��#,i�,X�Q2롅=��u
Jr�.���"����J���m��q穳���ވJ[�9/��z�F���7L��kkC��v�����s��9�,���QV ��a��`ђʾ���r��Qe�=���O�3%�ٙ�j�G��I_JB*��PC/x�q�s}ӊ���mP��`��qZpts��uWse�#=�TY�j!���V&��9��6�z���J�y{���2C3�c��5Z�mtr�	�����W2/�0!5�QN�}�qz�H��>��k�7^jbC�<�L����DFnmt�I�C��۫�{��N�^�l-�r<�=K�mv��;�N�J�|<�p�k�,]hf��gy]����P]*��;ړ(�������rU�঄��w��A��]
n�8u���(T�^���lHV/i�YGf��Z�;"�}CF�bꢹL�2սj#�Xov-%�G����D���6�flH:���:�ź��j#bi�9z^^�k��{
��D��!R���v�hS|�
�Z�����˾ g^���=S��_IY���n=c�q�l�&�9IN����+�z̎�k:7zŊ��9Be EmL�O��e��>�۶����g��A<eaK˅Y�ε�u��m>��~y���4���>���}toQв��%��#+tr�ը`���s�� T��J��du��N�ZTNF���L��p�������� ���[h
ݥb��{3W��V�Bj7�������k4{�>�B��q�38[[�������e��)��T�y=�� ��(*e]kHgۈ�cp�T�y$�H���hE���%�p:G��D��Tßt嫜8B�g3eg,lGE��9��U����p�5Z69ƽ�+��}��w�U��	��v����r��C83��
M�j$�ys�[�֧;�P�̷s}>�yW-�'�M��:�������w��-:�b75G̘�����@cC�x�c(o�7�5�"}���"�Y^5�z�W[wj��֫�l\w���&Y�-v�e�v�>�c1^����;)h�d�ĹO� g�%&�,�ڛ�ڕle��W;uܜ/�����ݐ���|�QBԬ=Ӎ�B�z�&ڙ��"��Rݰ�)����+(b�1�+=92)��C6k�b8�{DNU���Va��ޥ�����ގ�rbn�M�����uBx��Uy��g�����~�^SA�S�?y���*}��쩁�>Ѳ?Muxo,���<�5��)A�7l�]��Aq㺛w���+�Z��q��]"��G���������2���0��4t�A�5�{�I+}�}���ܷ�X�,j�o:)Ç��s��F��y��b�+G�>��V���4�<��xeN"��(��(j�#T�R���<������Cwh����4ZzB�������h�1�orh��O�k�������%�CcOA�N+��Y��e��W��*���pޫ�{Փ��5�e$@�6���c'~�-��z�޼�Qs��G��ǜ�>Ӯ��}ə�#�)kD�r����7�x��7�%�D�+nsĕ���2�q�]w�pl�&�N��,�:T�~�\�kQ����P�[��1͈[}�775PW����\qi�R�R:v��Ȧ�ӥ5��(O�X;��?+�!�#�����B�4����^���M���0�FGm��;���0�($Ɩe&��XU�jxa����}7���Y�`h�7���Q�݁����H
�]Q��8�C9~�G%��߶R	�<
��r3R�{֮���b�B����-��|�5%**O�C��h�pvIIs�&�!��8�_=pp�g�U�����.Rt�t�>�e��ؗr/q3�a^��e
����;|�H��)��B�k<�L��6��OK̔9��$�}T�N�jۊ��v$qʈ�ю��"���yqp,`�̱=��Uwx�݇1D"}�J��n��K�H�R����:g��N�]i����g�\]�R�7R����7�-��1�-epS�ȣ:����ty�[2��r1Ϧ�|�/���fP�nl��=R]�s8�^ϱ-��N�6�� ���0t[��&d�����mnr�7z�'q��Э��پl׭*"�n��(��˭÷T�7���k �Tȍ�^x�ݥu�)�)u��ͩ�	��)����!2Ha�R��r�P��*�ˡ�2i�{�C)���He*�I�2���aO�q@w�m���V�쫌�����|Y�a�r8�	E�9�㔲o-���y��ůH���������425�QE�8�@庚��)ܻ���Ǎ��96S�lW��M�jbCud�Zܫ?8��g-2��=|�{1nz�=��-�ϵ�*�M.��7uX��T�zP�A���{�'8%nV�Q��_3�ͨ�/�Ҽ3fF�}c�M<����bWC�U�P�Y��QѴ|V;2�&s��z�S���.١���qO9|zߨ��=�w�X	����t�	g?��{|��B��u�쑚�%+KuMxe��u1xj������ȓ0MfL��s��T���B��C���u�^^GDmbơ��[��OSͅb���Ƶ��ϩ�V%�\:��+W#���f�"ְ˜{#M������i��l����M�ܜZ���]��{���]^�k��{
�z$'
``�&,yӪ�QM6��!k�}��.~�s���Ꮾ�o�z1�
����M�{ӓ�=�2�|�P��hy��3Xg=Γ<�{t��ؔ��RTڛ�/�� ���\����Έ�#/i�n�v����
9̛Sjr����t1�gT�wʈ�J'͆��F��%C�m?rj�)��Q������`�u'�ɐS�Xi�2�+��P�jԟ>����W}�FD���6U�0�X�lSV"CN%L>9H�������CM,�s��/�38���Z���3+tGX(A\�I\:�ՠѝ�@��ܮ���έXvi��Uʿ��O�=�R�z�k�9!黺`����l]Ґ���e+[�/oBx:���'�̣s��c'+���I�],N����X��� ��`닷���S�id[r��n�kj��;�:{Nel��Y%����@�ڴ.��f��@����PO��v�W
�%�����%��[���u;"��V��TV�;���<��Q����q�=l�T[SF`8Z�x�m�Ut/>��ӆ��.�����r�[Е��[��V�wt���uH��|�z9�����c�k6 �k劦��Ҍ�e�y�-�Y�72j�=�Fu=�*gSwT��3���n6/1
i������+E��{y�mU�}:nQ�[|�\z#O�v@�ƳeX?�a�j�:�9���v�Y�z�Z޸X6���RL֫�g�cҶ�xf�m��}M;ظl�;�>�ynޢ����.������x�K�jQ�g�t�,¶��k,oVm�P�m�VT��Ƴ��*i��Z{'�WZ�wO�L�#c뾝Z�F�@�X��:�*�Y/�f /:��oO`#rnk�7�/����N�툪�E�1m[,nh�f(	H���F5д!R[��"��<���Dƹ�:�E���e��ڶ[%�L�.�9y�P��θ����ն>,;����^)6��k2���c*��.�&�K6+��Jv$&U���,�P��釤��-A��֬����h�)��)�^2��?
���u*`��v:��������C���m<�v���H.��L�JY��f�3�Te5�1]3��l�e s�������tO0�֤Ь�<s`st,�x��۽��]$�7#���\�ps4����ۥ\�'mӜ�^f�x��W��j_6�
���>�yu,��:;:�/"���sn����$�tA84n[\��aG��Vr�:�Wd�����s�Mj��׽3�7��O��z3C<�/(-��/p�ka���@���"U���اZ{*!�"	��o3����0͆�[CE�2�d�fe��x�V7y��r��8���i��#���k1F�s��-����#��i���2�p��G+O8c�:1������]
�{��~�goՏس���щ�Q�{k������q�̆�-�.��K���M���Q��h�';{��PvXG�c5C�v�Ӭ�)�p�I5�3�Uf�.#:Nb�շ7n&5dQ�b(�\l2�����Z�Z�K���Y�M�����c�KeH���6��R�u�Y�S��ŁP��E��d0���LAV*��QۂcDʡ��`�H�iD��� �!��2������j�Dԕ�IZ�"��ɉq�*��b�nU�F��"����������s&�UiPX�Ę�Y�X��X)��0Qb���XMd+UT�33w1�&0**�"8��CS2��Q��*ʒ�n\dm�P��mb8˴Rk�J��,PAA��M�l���
%ne1;It��ڢ���JZV-a�*`�f&8�lU5�1
�����H�T ��L�E�I�7'�V�2��3�{��iq����%-[҂�ˡ���d4>�/V
����C��k��t�h.G}�t�0騳!�m���噋���X]��ybo.�=JTйoh�������#���$��V퐥�5h�}�6�ɻYe��.[6�k%�8u��9��/�>25TJ��8�̨���U�^Ɔ��U}��㋆z1r�H��*]�}��T꒏t��,�G��"��iWhy�ڼ�K��[�)S�R�<����^��B�m�VM��	��K;��.��77}5���NA�C�2-N ���w�����s�V1nr���Ok�v|)��3���^��A�7l��qX�iot<M�~�rӦ�)W��F��|�6�\��5}��b��7�B�u>=��=尐�w��8�V�d��ڽxC���=�W�N��yV�����O���s}���f�D쁥���������7�S��p��4P�s�wȹ+F�uݚ�wjr� �3���v�zL(�e���U���ۼ��W`�����������u:k��F�TU�}g�����f��Z�
���UY�����"�sx���#��)gVIQ!8X{�N%�Aܰ��H���A"�.��fON9�ohr�(OHS��,�0"ڽx��`&U�o�d�����}���i�3��]�eHuy��Y�0Q��4�h�J��Vox5��Gb������ۅ�Fef�x<���sӷF��9N���n��q�t�H�OՑ7ڸ��Wb�]%_DϚ���5�.�E&�R�S٠ԍ�Ŗ�����c���2M�5Q!���4���zq�F*1�����{�*7����c%�u=R�54�r=�/R�����d���rSy�(�ig�ew{˔�SSٽ�u�{8=4	AV�J��gj?�|��m9����Awuް��F�7��
���/C�*�`����eL<���I����t|��[�n�GvG]|z��-��]%�:ݛ]�<z;���ԩ�;���JoyRKO&,��ԗx�b�w��^�2�k=)g?L�C�4�*t"ۚf�p�՚�17]9���i�}�ڵ�
2���b[�`�v�ڻ��$�D?W�^��K9�!�2���K��A�Ƌ����q��)P�]A�n�7
��c�r��ю�'GQ.�m��uٽ��a�ڙx��5��N�6�D�;��Lؖ&�N�I>��'ޡ�Zc��VE���Q�m��ۋ��(��;MG7�^0����7�<zfu,n��ҿV�4��S��Wك�@�4�J��\��Ho��CH���mא�T1ˡ�<w���w��k�CsXftjXtJq*aON*!��6�V�8f�i+8�k2qn>F8d���r5e�!sӖ�M�l��-���ȱ���d�X:�8��J�=M}�ޭl�S!�#ϊ��F�"�e�o��/͑��I�����y3�"h5η+����-�F�"�濲m��I��]��;�G��j9H!o��FF[�2RfD���%��	k��u���a�j,�Q3�q���v5^��u3��Jwˡ����P��42\���pDqfRn�jb_D�4y�=��ĵ�х�yV\�T��{�����u�h��+|yr~��-�50��+����W94�
(]hf��t��%mR"O��S�ML��	
�|*cv�¶��C-3��pu桋�W������4�3����
�ny�Y^;7GZ�;��9qܓ�P1WZU�"�m6�!��J[�V���>��:F�\͉�%�ږ�YwZ���׬m�f1]�C'��U� 5��=�XG�Bp��܌��dv5ݨ`�Q�?uݞ�)/+�}[�ݏ�[xXz�A�����q�k����L�T/i����a�3�{�S��
�0]���:3OgSi�qB�u	����^�.��P�-1�k{�,&�k{o)����mp�'Xq�7�r7;)_e��&ּ�fXo�B�u�tM����Q���DL�p��Y�����;S���I0,�Bu9>�g��b
���u�K�	{V��͗-����:��A�L�m3R�{��zӢ
Q�N���hCΞ;9���[��Bw[ͥb�d�<��="�3>S
{�̬��ӹ{�yw1��ҭ6{�2X��sb�Ոi�0���O��[�����bY�s2+)N9X!��3�p�5q^�:"���<H15o�F3��o&�M9SB形���D�BQ�+r�|����I�j��.�mݫ��aBn�
�u6Nm�X��rL#v�3���
��38i�K�_�/溦��-vzA֩��.�+%�w]����R�D�	d��aԫL���O?P�|ڮϹT�3R�{z���Y;}�%X����CI���:�NX~�B}���}ӦF���/}�]E���؎��\�����̣�K��H$M�Gz���^e�[���W|d!"�ƺ����"M�i����[��9]z�t fL����,Ow��t�ě5>���O5����]!��yM+ȹ8���3���S�񹖻�׻ �#��Ѝc�9�i%��_lۅB�s��!%n�R��q|�O��|)S4:Q��m��ŕ�j���%���3���h�.�萶O�uz�,Z�;C���ӎ�dS������ۛN��l����!�3��/"cf�݇��ǚ���ø��]o�b�h,�'�(�'��VřpvEѱ6�[d�6�n���ǅ��,m��R�T�g;�H��_0�A����X���U�ˡ�3��x�-N���x'*D����{��y���!cf�)P�+7�T\�v��r�=��uQe'8��f�i�"�)��01LO:6�IϦAT���_<��xG^Ю��c~r���ANpɯN�/�����ǚ�l�P8e�w;#F���rڵ�䥣I'�"y���|8���6:Ö�\��P��jשE֖JS��j]�5{����O����h�:;��M��{jbE
�EUkT�E����Rb�.�i&�j�_�o�w^��Mq��^�c2N��P�a�r����47�H>�֕�9��	
�����i��u-�vY����b�/�K6lV-�Y���O�I�G���Ē�#��ͩ`���M�vmܕ"�M46���ޙ��bbɚ]i�Μ}M7s����l����4,j���A�_q���n�[VN���t�]ѩj;�ZQtuʧ:��Cz��~�p����׳v��FĨ����jۊ��v'�r����2�؂%�ˌ쳘�-`�-��Փ/)���mbvh��b�7pr�2z�8����Cg��>�L����R�U�x��f��fϱ�Φ7�f�ܹ�5��(�[S��}r�kg��Kv�ۍ���[�eߺ	{�Q�ΦѦ��W�+�p�{�Cx����fT+#��2�h����-#q��b;Y}O���І{�#�����v.��m�/ٲod��!gS��ۻ�k��!~!LԆwӋ�Q���B��0��CO�i�0۠�J�\Tkf \m����e�T�y���I=4���k|C݃m:�|n�s���1')\��C�qlSQ���Þ��bo�A�6Q}=��؎�-:7�n���gX#��A��-D���fA���ꅽ2��0�m���w�@^Ӛ�rSb�.�R~�r��<o���.�7��^	�p�N窝X�oog�Ky���"h�nho:|�b�2XN�X��d�W93�nh�um	��U:1�6�ܛȆ�������yW3K:%�{^|*cv�ª8�Pu׼���(ѤV���]�%2�d]�8�ʜ���՞����^�U,=�W�Ε�'��ڬ�ȵC]D��!%�D�؋�%�P9���g���M>��%*�+�f�Ӗ6]�F�{ ��<iTac�e\{�.E	n�2��3�N��V�vEݏ��؆8�SS�z'JS$�}���(�>�������ep�>b ��G�����J2e\�#��5F�/���}[����x��T�7͸�=ѱ�g�.-���{����H7�].��O�^W����ﺱ�����Y�T�]��E��4\=����@�H���JΜI�;wFQ�疢���Y�rt6���{T��I#6����ou��i��7��؎�t���%L�rAJp�!�|GSQ��Χ��k��n�#"tm���]lϋ|���+ʙFZ�Or&ۇñ<J�L,F��F̋	��lϋ1͊�V"yCE���!;ٝ��Z�l>ۣ�f�{�<�Ap�7Dj	�T�v���]͆2��s+aON۹��]��9SB�۔+�[=��㫫*<�q�,8�9D ��P0�'v��6�����oMC!j�L��η[O����	Sl�M���7�-mpƆ�+sM�4�[T�Д�{��y��0�ÇS+���7J�H`X�W�>�y��[���y�R�1�5�I	��o���]C� ��Q?2u���f�>f�LcfU�+�%h��b�s���y���^����}m��}�/�~�8��e#4�$+)h�'v�������E�\�/�W�
�Y�s�ԕ�R��'o�D�b�x�t�;��&9������7��}�|^hG=�!�^|Ҽ���9?���ş!��Ғ����\x�>�hIĪ�ϫ�P�7Ҩn�y��4�v�5�b�u1�a�}��#������b������7��O1z������M����R+��qP��U��-V13��s��贤��������JΝ�/}ѩ�S�ߩt��N�KĮ���}�YՒD��8 �Ff߈�A��GM����]	0,�]˺j��|1pB��f=�V��n�����V[�8�ۛ�=����|��\ͫV��5��L�I��H����8��������+�х��a+I���w����)���]LdS�,��ӹf�,V:�^�TX�mԄ�㜪Ȯr��4;�`��:�+Q��d���.�7}|�%��|D�������I_7�k s-D��0�=���)�'�#��uMzf�e޶8oV	e<{���޽1PtF��`��ۙ/�rEWMTfam��D��{_ek[��0�����Qd�ĭ�+&nѫ'+W�cYt�b���<0���X��&��tC����S�՗Y8��&�-��5�S|�>��}sh�t�h�/C�{x�0����v��pf�[�oimӬ��E&l��+%ڙH<C�2�ޔlM.�xlՔ7Y��#�S����f=+f_%�lw�k8�o��0�F�Zp7	�x���%9%8G:��c\Ow���*͓t跹�۹�61���˽bd�����|�dݖέ��C��d�Dz��VR�y ���{���Eq�O�F���qe�کrp�	c��}p�r	N*���N�5�3%��Y��3��/*�&��w��A	ӆK�u��'׺��K��q�af�9f��J�!�����z�:z(8�u{:���u^s7cm�ٯ���%m��u�n��]Ʋ�JTj��c]bQ3%��y����pӖ�r�i�_;���6뱦�16�mF3��i�{�z�f]t+�E�u�u��Xa�N��U�ݭc���TEe��\�v�;�#�{4�lR��[�FG�b����F.����݉\�ݡJ�h૑;�}o��K�%T7aŝV���n%������Y���-�8Rѷ��%Ye�D�x;�R�l�e�[��\j�0g��$��%�5�.�ό�S��P��dl�m�%I�Ͳ^)�SS�'[ky�h�ւ�9O�Z	{��pr�^�'TT���K�]N���m���\ɡ/aΎ�C3N���6��KB�ރ���z̖��[mY����)iC�f���&v={�1+����V���'�YѮ�ra���/9ڲ�D3)�iɒD:�1�H�8y��_^�pͺ�lKy{�o�V��+x]o$8AgF���w������(����:�Ψ�f�;��Z����*���G�����#��E����Y�~: �"�,�Ј�ϴ�J�6�ڊ�UL�+-�*�(�[X�j$̢2",�J�2&�֫E�PX(K����uX(�k3.���ef�iZ,ܦ%j,U��Y�����eefڱA�`;J���J���m��K���iw2��4˙f&e1��*��-�.\��h9qEv�cXPBT�E����&+��*TT`�Ԇ�6�]�TR�k�f��Ī��d�GXK���(�J�6ى1��j-AA��\�!�"�Ԣjc1�bT5(�5��ʊT���b��ԮT�r�[iY�a\�u��h�멉��h�m�D�1�q���i�*�*�U2�ͫ�р��Y�7.ZUAJ�-f ���:�b���̮�Ww�Zm��"���fn:��E&72Ma�B�i��T��&�����߱9�+r�_)��E�s�\�^�%*u�V�G��qz(D0�MfqS�=G��R-�:�Λ7�j[�կ�x}!���vM�-�T�ZzEi�i5���=p����1Iw���V�]�0��^oơIuozP�����j�M����V�X��w}K4D�U%�o"�	\)�kJ(��7ӷF��~|�l9M�y�i'y�'�c�ë+�����1�L�1���bo�m_:��s�Y�ьs[5���69gd$ܵ1�>qƔ�f�j78��;�w����=��ʹY@cBr�u�j��T�ꁗ[��"okF+B��⌃��鹮[G��7#5*
��_Ls�8�׫�&�%���+06+#M3}G)����ay���n")�mC5�;����7���!�Gf�j��%�Gm��D��wq�c�O�e�k�Kw�������y�c�������9aJh�^�B:��6o۩�w���B������P�ɝm��/	��'\�WG���m9���r�p��$-��F�DQμie�E�o^�:��l�͋����U/7k�_h��,�<��ς�!J�E:e�&�w+`�k�}p�J�[�^m[�nqؑ�9W��َ�a�\#��$�C{}\�ީ}S/)���n'GCn��J��VU�7ւ�����As�aKΕ��f�+��Y�(U��Hb�]����>}��gI���0���t7v����ۥ���S�=��;-����)R!8x�l����)�q3�.x�8ݴ�픬��PX�4�ԧ�0��݆ݻK�{���șc�J���^�u��a����(Þ���Ot[ɫ���RP�V0��Q�m��P�825����PW����{k.�-atj`ySW7}�j���s�ء�t2�r�F���}��DoR7{R:�bfS�7�]4�]����E&�M/c�FP�������v���]ܙ�d�ᵔ�Z�\�f��V𧛰,`
}A;c.K�~�����-뜦fG��閏sn5L�@5*Vur��e�2���P'+3PB�a�pM5h_q�,ɹ��Z��]��|�d�O�A��D�cp�ݢӮ��'ˇN��&��rf��B�[B:ٽܶ�T>V���{L;9��֪�{jB���Cv�	�T,�K�ՕSf�\o<�\�.a����q�Os��lHV/i�YkG:���f �m<Cn���;��0��᤻��6���˛��B�t�^v�AhY�L؄���龕B�K\ێ���[b������p����" �	zi��J����V��ll�FXȁU���|P��ŶS�=�R�bÐw�V�Ԭ�I�MB�v+o&�C�����ͥ'[q>{/jÝ$��+s�(u�X9��U��Y��H�=�%Lд芔�{�˫8Vž�ڼc�_�tz�=��F&��*�����^��>��c�_��>���}F!�c_v��WX��r���g�<O8�.Ύ T[K�1m�n��:]y���t��v�Y%:�osY ��t�Y�(��&ε�g>Gy5*#�O�[��.p�nyKzE*eS�T��73^�Z�P,��T�b�(�p=F���q|X�Ü��"	����S˘pg��p�7�r��pִ�D�h�k&��.��Y�b��9N��ә��`۽J��T0�&.K�9A8�-+�Y��7�WC�q�ex�(u EC��n�n�&���1ܨ9��	A�/I�M
��7�f�@��l��e\V3����ӈۍ�\ �n'Kfb�q�F~���Z�00o
+@��k����P� �����=��GY��y�>�W�Lh�.�t�l��i4wQ��/��o��Jq�;�Xe�V�)�}���(3C�F�z=�J��͚�^P+Ƕ�%9:����q�pa15�䉋ۦ�1�XV�~^���Z0h��`���>OVәG�)羭;���.]8ik1+ã+��:�S��Z�u��v"q���Ẏ�@���y�J.�)oh�fl�A����\�_9;�o4�.�ԡt;�{V�1^�=,g���5rK݂��u)e��ިt`eN�L`,�VjN���E��Av�>a�����Z�`��R�"2�i��'҆���:�<3�nC�$A���(����hT8����Y��-w��3{o:{S��Y8C��D6z)r�d��
��� *�5�⑃��K�!��[��=�v|��-�8i�EZnѿr�_��.��Pຎ���q���1�oz�(,GHدu:ؘZ\p�1���خܛ[5(5^��(Qӎ�^89y�[fF����¡�}�A,�3��y���:�6u@�_�e�)/������P�� /���ZD=%C��@��l�{"UeD:.�OEt� �kj�'V�C�C��@o:�&�K�^U:X�3�n�й�.)'7o�g�7yOwcH��D��"g%��C�j'�{�����ׅ����E�o���P�֢���C7�EČ�/���0�#e�!n�x���j"��C�a����5�ev���KYa-�o�dU��M��Ne�!F�g��hj��>���#�S�yaQ{4�@����0�fGٽ�r�����S�S׷��D9�y&Eu�T.�wώ�F�Be�:���)I*�iy$D���uæ����|n𽓑sE��뭝�&�=��G'A)ìW[�o]=' ����r�T�������%�`r�u�|>ϡ����LkT(EĢ���$�ĴN�����5b�~�2���(���J�W�$Su�~ʞ�\8�oO�)��a�â:�3YC*����^������<ء�P6M�0GJe}~=C2���z1;��+ֽ1R�I�uϛ92dv��u�S�Pb�C��~gU]T+|yՕV�ú(S���|�2&0����8�z:�G��D������qJ\H�	��r�n瓳�b��'�olX����wP��t׬�U��r)�3pU�D��*8;��y.������/�A�*q@�i���|}�'`�eї���U��OM.H!4"n�B�q#;��>�:���˻����C���i��Dj�ERI�*���`��h=�"x�$�zjzET)�CfƑ�K�1�,Hu�uo#K]dm�wU�/��T��ALq�Lq�i�ϡ�f2z	��1D�Z�2����r�۞���W�����|nk:�>] �ˇ7p��������i�U�+�W���פYMǸ6�*�¹���(��� ��v�K LZ��c��'�hP����yNv{-�*��/�Ü�9W���W�^|n���ST�_�u�6Hp&t܅���f,����\��р��(�!E1%>�pl��p�`j$d�N=\`�4DY2m��g�*�/�Ո�#����N�["��8�f��;�C6!G�����3��%u�A��`kn(lP��n��qw��g��zW�<>��ʡ��`/kő��3ٚ�!vf�NEBzdr��5' WX�85J�B�[;�5"��p�<�z�
:�7�����Goƭ��&���� ��\��B"�B�h�r�+��s�<� �C��[��<���ƚ+*�>�u<��ŚfOa�9f����T�Mʴ��{�X*6��%��?j7p�<x�;6��¬��ѡ]E����Kf7�9���g����<B�{+�u짿
�Z5]f�>�p�=�@L���Eb�����Og���7>��R��YT���˅��6��1�Uj53�o��0H���n�W]%X��q�֢ݸy�%'M������&�eF�db�{�Z#{;ʹ�e�����m-�Kw�No]�\�̒Wl�b��ȘF�M��Z��
��)t�a�9�7:'���w��(mHOc��`�%!�[��{�l��X�N�-�T(t@�n��:��E���<9��K�<ɜ�ټ�R�¦&3T���S�l�h��+`HT�舌�fğuj�,�5 δ����^�<D����@�zʇfb�*�6r��; )�!S(�c>"����	��ɑ=W��a�G�=��#�6ϩ*�&�	��Fbx���u�7�Ჰn�.�Ήԭ����.�
�C%���CꑴKr3�Sm��!�T��
��-<H,�1��d�*&,^*q~�z�DCgx���鈫z��Ө����a������W�i�k�U{��
�y�^g��4�dN�Q�sE	9�;�@�!�65Ɍ���N+�8Λg�7j�zJ"��f�����+z�&�cL»Ȱ��9.����Q5&�I��Ю�'t�M�3¥eY[��b_�9� ��!��>�1����f)d��]^��Z(��S�+EZ�n�I��	v,�\|v���xڛ[Wk�.������Kl�m18j
�]xz �G��/lo�)����]Y�-���/����83�t�������]��,[��$`mvBU�&���I�&��������5��ͽ�Tho�����m
ǎ��C�u }�U����(G)4|yԍ(L�k�^s�
�.rU���ت�:*ԁ�J�v7��J�`r9�D/c�ӣ����ɉC>ۤ�{�Ԯ� ����������Yc��W�����J����%a�=~~1�)���cÅo*Z̤Pt-��e`bx����<��7f�����p������> Ah��u�S�3�Ш����Q)׌َ�.��Ք�����G��kH�R6�R"���G�[%�GAж(*�:H��]�g���������X}^�
��Pe���4�"��W&�SL��~ו
&�3��fֵ�oE&���ѯ�>rؑ�t[�[�+K�F3\\�b�rl-���J���=�'>�a���1��L��.="=��<|�h�P��^��u�arqB�9��(�W��@��M"�ӗ���«�"�P.�[6#��eD:,�7��gN�{T'A��zBŷ]8%������l�	��}��­m��v	Z�o�D�4Dn�`�����]L+��Wut��n5��/G�Δ�-���ڒ=�{[O ��14)�R\��L�:c�*$���[7/D5��.��=���|��(V�9�*S�T����v���)��m6"�GYq�WTAJ:�<�_^��w�0���rp7Ɣ�����t_�	��YTѿi�B w� �ql��x���\l�QLt_�Wt����826׫�+�7�zh��dK,q
8AgҔ�j�T,��2.럛���:�6"����ԑq]m�����|�G��A�����K_�9��^���9&�Q�CNE�\���1�*�W�&�����7K�O��xx2������{����O`�y��ء��&��3
��YB1�\�4�"�f��S�y�؈}���MNi�k3ڠ!Ь�Ә��GU]+|{n�>��2n�<}�z8r1��γ�D���;	S# �T����
/�#�X ���p�o�k��Q5��8+B��Ӭ(&~�����s��d�c�/��U�j�����?��RS�
V����.d Ii���$A��!APG0��E��N	
P�cL)h�zjP��c�&1 V�P	�$Ā$�G�;B��28z"CT8�*�*����� "��ubR#H�(��m����K��
c���M����P��`1����!����|���nH��g����+�J����u~}�iǓ���EA�B�*���,BJ��3�E{S�C�?�_"Ѓ㪗��8'a`�u�IǸPT��|�h>Pva�@�낐(�o�f�l���ސ��@����w��q��#J�P,�� �2EAƱ�%q���F�Q@�*���U -*D�"��a���I��S�0�˦��jfv�
�:7����b�w
h���wn�!�h���525�*���-���w��%#�-�!�
�=l8��׽4����k��'���������rJ}W!=��9�=�/2�ܼ�!���v'L0������g�q�,ЏZA�����#@���(*�}�X7Ž<�BW} �G�:T<C#�":��_]A�6���2`����~'�>  B��U�� Ά�`+����kLL��P��-����e<p*Z��}h�`PGQ@��s��МA�Z�0�ck�` ~ǳD�g�@=�F��5����o^�:�=�4�rC�}O<��<<�ԧ�~�)��x��أ�#��N�APG��T-�#���c-����t]F�i�vඨ^�B3�J��A�o��pp�0�+�@������0��9��W�,(*�7k�6�ܑM'��Bc<�^A�ON���Tۍ�v��P	:X$�
B��#�`_xC˵ ����:�EA+���%¹�8�Z�\%q m�%��t �ʐ{� �R�l.�w$S�	�-0 