BZh91AY&SY�kR�s(_�pyg����߰����  `�>U@  �  �O:��d�  (��g��              � ��
ǁ������   ��n�=���í;��];��n��z�-�����fG����r�wx*�Y=��m]۪������{_|>���n���V��ݽ1׻u��>���|   �p�}T�����v�]���ͺ݅�;�=���޲���᧼���{n ���o=�K�x�ޝsd�3���j�^ݧ�=o{��ڊ�E)x   ��׃m�çv����;N>��ػn���{��;{�w�k�s�������];�oF��ZlgGst����wy�f�����  {W�ޜ흲�}�p{��gpz�n�������π��G�=og�p�ٻ7W]�;�����޷y��������W   ��
����uȯm��k�{��ͽ�v���o���o�W����>�|�;�]���^���yݏw]�׮�G      �Ѫ%PUT� �H
    U?H��J�Ra0��1���S�"$�R�`Dѓ M20`	M��%J�b`L��i��# �Q ���F42b4�"H�	��
yL���Sd��a��1Tԉ�)U)aLLM0 ���匞ik$��X�y{��(zI�rza�1)�EU�2Ĺ?w�TA*��!�A�G�U���
�����_��ݛ����è�$�"�PU�P>���z��J	�̈́P�U"t1�An��ڀ�!�~\�r�o���ϗ��`�k�M�`���5������k'���W	��V��5�q&Ȝ�N����[*��"sǺy�{����B	6����%��H���p�ғ���H�K=���{���D�'NlNèw�ԇh�/Z�Z)ڝ1;��E7ݯ:p�8�&��M�t�u�u!�I��2W ��%�2s�:�4r��M��&L�z����Ό�,�չ>փHm��:��z��#��Z�վ��G�:j��G�\gD���'����tD~��䇾N"y&�=�J�:��$O|�>��H� ���D�'�NQ���	�Qx�pzh���;�pI�<&�t|A����Q%�4�%Ĉ�K����$�����l�&����DE�(��Ϧ��R'v�4<�O�<Yn��?Ak�D�D�xI:M�&�"R">,�Q"'�E8P��-<�P�+E'�??,�D�$O�|��"n�"Y�D�Ig�Ⓟ�Ђ�(֒&���DJ�N+�"'�e�A����C���h��DzYG~�"u�>Fx�h~ؑ�DD�6A��%�&˴��Ot�ɳo���Dw���$�i:y�>ttp���֒$N��Ĩy ���:%%�焳BY6;4Qq&�N"z�}���4t�<D�-)�&��M��=���'�茞7S�78mӖ&���������'���oSD�P�7,M؋ڔ?'dH���މl�g�l����~v4O|���r�����{�&��͝Ჷ�G�y�����ꊓ��o�I�:��g4&�n��K�'����zUץ�픛Ş=��������zY�8��2K1���<�,ݞ�vW�+�G=8]j�&\�9,����˞3�Dd�t�O\�8OD�B�}��Q��F�QD�'�z��M���s����A4z�Du�{�; ɢ�D��"&��(Е����q��,M6�J�n��i�AU�M-J<Tj|���"�#;S�;jY��FO:���{�ϸp֢#�DDR�g�D��v�p�l�'jY��D���R��DGmO)$�I��"<�Dd����",�7�TD�Z�Ag���z�J��D��Q:oMJ ��#�TD�ʔ#=Q�jY�AU:#�����6v]M�u>Dy���ډ�{�DN��d|�4���":�D�5(�hu>DoU7�T�ꈜ�R���5��T���TG���#�xj0J<{q=s�m�䒙^�(������%m��n'Q4h�!�7'M���rxׄ��9�;e��lI�bMDnW�ڞ�5��Y�ő:'Y<C�u�D}ɧ�(~O5<w�:[u6=5VS��T��IrU�4NN'tDM��h����(�jS%ZRlM�lM��f��e��f&�{%{%p�b{��/�ewu(ݎ愾�6W�Q9��O�����h�����D�Ȧ,ߙ��{��S1e"�b|�$����~d�2w�O|���{X�"�6-�=�{I��;�w��Ytr�+i��0_cg���}�>������l9�e�p���;�`��3\N	��[1RH{��u�N��[�J���]5��U8=�f�t{5���&�4���N�}�6hI��g6$�X�A��ƧsA���k�2��i,G��}��ƫ�n�Zѳ��oN����)�S��K���">�,���Ϛ����TN�ȵ)���ԮG�������W����1�l��ϙ�U��i�y���=��>c����=���3���<>���CU �n_̺�c�TX����7(ܝ�N�)Hq$�Hl�'*\���Ƈ�i�L���}C���;�N��˕��ӗk�s&f�)��N��GL�?x~Np��O:���<+�����N%&���[�)*����}�:C�؎ګ4?'D]�x���(��<5:�R"'/�6;ܭ�nw�4%kғ�jX�y)<:����ʳC���H��I��#ȉk+��G��jW��%~�ᨈ�G�MsR�8=���|�ڕ�4�R'�D]�ᢷ�N�"_�]4w�DG��d��G艱�D{��O��R�4�R'�"�W�rW����V�׵*��y)k)8oL���r�4=���+��?D��e|���ѡ��Q�%&�����JD��';��͉�D���Bb%�ؚDM>��7�W��%b'�����.g��v�Z'���S$Gr	o�'N�*��}UO�+ޜ�N�t֧NI��{�F�G�8%�X�=櫧����rhjYkӥ`�5]�w����y�V3a�L�A
*=� ��Q4�}_{��DNpٱ�E���+��<#�J����OMrM���qz#�NIcQ8q�W�2:��}�|��'��G�>�t� �����"58\��GSG�u��5U�u�}��=�]ۈ��d7��;�5:w�wq���OyƷ���a�ۨf�!�	�)xzi:a:e;+�T�j7	�K�����v=��5~]뫽�]b��}��k�=��uu��ٞ��_-]��d������G�6{�o���S�}���O�}�Y����g�+Q��ž���V�T�������I�M����;O/���z���(|����Q�W��l���Ke�\��Q9��!��Q9�4h�+A[T����"���{����s�nuI��(ζ:䵖���h!d̨~|*��D�j�~��T������Ko���oY;��}� ?G��1�d�ن�Tv5B������=>��W�]��a��̓�h�pǁ&�6� <�}�������++<]����![��N��7�8v5�A���}p���e�q��/��:=��}��!�NشV�cO:p&©�9B��:|�Ϭ�n���o�ն�w������_��p�L�>2���}����7�5���zϟeY{@��Q�Mb�,�8~�����0���AM a��=ۛ���d,�n�
�\����0c��0����:of��ɒ�S�˰7l���vn\��&��ܞ뻲:^�wB�I����_Mٙ�6=�N��>��Ͽ��~�~g�=6�_c�`���'z��&��~���x�}�nK�Kgf�93�����d����6���kޝ��'�v����b۷V��/nb��x��{�yz����{:�gK�������m��9_�>��}�?l=�Ο�����y��w�?��w�N�c��e[ۛ;�7�1{�}�Vf,�L��)�?#<?�ry�Iٛ�Z��C
n�x��x�q��x�A�u���|���]��N��Sl5c1(d�>״ZM?_����zw����v{�}rs;�i�Yc4f��e�vɦ�z������.��^
k�v|ot�&�fe�n@���.c��[���x��>"g�����P�H�>�vY�{�HΙ$d,'zY�XT���f�V�޾�:��g=ּoXz�HL�յ4�^�f�ɖgg}�w��H����!�׋��h6G�y{�@.��n:�e�Q3!���L�������%:;F`�����ӯ&��3��oL�z`[��mR�E)�Q�m�-�f~����P���1��w9{۞׫s�g��{ڷ������ό��uO�ڞfǎ�S�}�*N���p���r���Y�gG�����9���UYoy�n�E�J��{�w���!��nz|�'ۜXr��wZY��w7߁��.̃S�#;�܊���]z���\p$B����gEj@�����F�"��O#���}?g�龝��Yc�&�G�tb��2M������[����/Hk�P.���f����/�w<kD�}����矶ݐ����;��L�_L���\7N�
{*���{�qB?<׏{�&��%����n{2����XJ��L6�#v�Bl�����Ͻ�*y�j���~�jd��o��x�|�W��v,U���?�31D;#{�+��`���{g�r������ᷟ��y��}p�k�׳ឹ>����(�2��]�F��:��l�!�<yV?�kb��F<���OKՙ[��ߧD�϶�/פr�?k���=Gs��q�ϱ,��za�!��϶x~/Zç��|a�'w~��%_.�zw���_g������u�5��.wǬ�ğ��;�%����@�H��lބ�fz}�oH��4��&�]�m���H�-n�q�n�d�̝��g��_߼+�����h�I��p1y��6n��ӽ�ly��4g���>��2T�ڷ��J�2'�*ɒ���&ʝ���j�wo�{x��o����tsT�W�e��%}�=�ںw��;���O�%��������íX���]�Zf���_���k;9���D��v���hg���F�b5oo333�*�Au���`�!�ɝ�G��=�s&��F����X���݆٠v},��������N�3��z�c�2��+e===������R��:|q|�K��{��Jr��6A�X1�:q���B������}ܝ���y>+ߧ�쏣֜}�6�����v'�*y�饽�N����=���g�C;#�S�|ڍ�O���:������-��nŷ�AΘ���L�/}ܪy71{3�dА``fN(�+�d��6��G���n �ٶI����nJ�{�4���z=�
�����t[��߲Od�Cl��w��ӧ�w����M���(���H��gs4f�;G:A��M����l�����n;�$�e�^�|q=����־�;z鸳���w�ˑ)��|�>�������S-�|sf/Ӑ}���g�TX�>��L��He�����·�va�?oF|^�!��s�G�7���gU˝Y������t�7TFיW��b`����/�݃>�`��/�O�	u��W$�.<ަ�јk�Ʈ�b��zZLci�j;�gd�]ޝ�^ͻz�������Sbx�;7^s��ޮ%��5y���ϻ�����&͐�}9���d�_�����t��$����ua�ڷVt�e<,��${%�og�W�bm��?_�ޕ:�|L=�7�?g�,�nۛ��<<M���M�g�g��?.����~��~ثw�6�T@�rěp&b��?	��]�ޙ�=D��\����3g{&�C3g�.-����0�=U?{��y�`�>-y���z$d��/���y���Y����X�@�x���ྟ{vn�̯g���軙7{�[s�ty7w��f�S{Gz.�r�������نF>ܘ�����=�ݞ���쓾q{�����{�^[�V�#�{�~���}#잒_%T��wgj�;�*��[��/��������H���>���>�e��fi�p�N#�w���Lv��7a:�����G�=���I{��^ֿu�y�tc�>���^x{$��v5o���|��Zc�j9�(�gf��4��Y�>�g���R[�x��i�X���Ω����}CO{ۥ������{�����S)��Sz�|+
�7���f��L����/�������_l|�I�BB�!n�<��M��Hy��48lZN�l��;���rw�-E�:m�4ڛ�`J>	V�\��Z�Um�h�WrT@�E�%�Z���E,n:�@�L��_����P��T⢒�+�T+TU91 ��PT����mA/gs�ȯ
ܕ���tn�1�������<2�T�XK��H��Ӎ�e�Ð��p�h�D9"���T�C��7TmJ,1b�$'$M*A�Z�ej
��D��NDZ�n�V4�R�2H��
�%!clT��z,���vLx�P��� h����#dvmH8�A�Fr�1EJw��GINRp���F�J�d��G_Bs�J��++�+e
X�Mi���na&&ꠘ��|#Vrն+f`H�c���Yh�/fc�R:�t�W�T+D:&��2�[YaU8Q�G��v��,�|;SB���ʅ[�Y��22�FJ���c�V��D3X��"�O#Fb��q��p���X�L���J�@�����8'R�R�YF;� ����GP��KcT#TM�R�YE�2�R8���l���mn�Ư"�ݗx���=��c��������-�Ĺsay�1��$��j�8�|���\�#��Ews+h�\*+CH�jj^&*��"j���78݊��,LM�o�i� lU̪Z	���#��cBF��o���q���F� �k1ȮT�քȠ,��(�D���	��1�(�.V	�Z� -�շ	��[�ƕ��Z%��hG{)�&�%�c�D�%��cX^Pj���Ue�w&^W"9a���CN���%����NL�&�Q;l$��1<���qN0+�R��'���s+L���dU+Z�񱦵�"���A`�ò7�WAյJ�l_���U��k@�C��,;��^0:���&wmbŐ��L%)[Pv^Q[�9T�h����=�ƔD�jh)�� �
��)qe-1EH�ax��e�fǜ����Ux�k�Y�-��j��Zڽ`��5����Wց�>,��� ��[�;�'VȪr����x�������_s�?1���;�N�HH�������L���J�����UU��U_+J��b���UUQUUV*��ZUW�Ҫ�EU^�*���Zv��QUW�J�w��QUUU�Uz��Ҫڮ�V�v��Ҫ�d
����	��}��"�AaYJHC�$FB(D�Y ��)I���
Q!?O��O����V�;�WʺU^*�Ux��U⫵V�k�x�X���iU^��UmUmWj�j�V�U�*��iUګkUV-�w��⮕W���]*��b���*��iUUQUn	x,�$!h�U�*BY �$�Qd"$���RD`(��#	(`��{�*�U[Uڪڮ�U�UW��UmWj��[U[U�U��UU|�Ux��]���UWȪ�Ү�W���{�ۥU�]���*��*��*��*���������O����H�!
�2
SB��JT�J���������w�UU�U_1UUQUUQUW�J��ZUU�Ҫ��������+x����W������j�X�{���*��*����W��U^+J��WK����{��8�@X)A�B	)��-D*+QZ��!�"H� �
���!@�Z��-AJ�� �V�P
�� Ȝޑ�K�J�㻷�|T@`BI�}�o��}���S����<LS�Ͷ�Co�8�K�un�Z�mn�o\Y��N	d�M����:AH"hN�bxDN�i�lK4&� �DK<'
DjO	�DO	��p�,KblК��ДFB���6 �"Qg��,M�١4A�B""pDO$�"%�b'DO���f�CB	dA:p�&�ѡf/��/�~��s�� ��$�ڀ��T��Ň1lH�%rI6VV�DUQyUdl��j��2�֨��ʱ¦�kRI��P���e����m�G�-nQW*��ѫm@H���-l��ʧ�l̪��ʘꥊ+�Y<T��ҏl"V֙\�#�-�����[P�\MFKk������ʜN�Q�@�1X��&��r����~�˳R"�YpM���p�9i\W��jN�؝+��Dr�ɂɊ�����`KSFX�B'%)
���@��'G-u�T>H��o��2'e�6(�n�8+��J���젛�[(�V��B��U10�#�u"��ȝ�ơ*�L�8�1E��EJժ؝�����y��AQKG\�X�C��F劃R8�c�
�[�jz�ԕFp�Q�✶H�Q��.H����=Y�6e����'l�RFՍ�bm�	�����)cB�n���Ͳ(�R9m���iɺ��j��żz(�#��Ђv*�%�Dlt+��UF:��6��E(�uDEj��햦�!��X�u�E,嬴PU��eL�)G+�ƪ�F�*��Z�D���TISUIIA6	���Q��B[�┱JX�R;EKd��k���h�Ik��q8�rUa�*dt���jq����J�/#�0|��2���*��L�iϱLE18���|��|�U����>VݭIYh�ҤM0��R&���H�l��Dh����8��6.h�L ��E��)cQB&���B�:F�rF�r)�ڵ�b�ChZ�߷��X���������̙����X�����>��ə���劯.��p�̙����X�����>�>��u�q���vKun-Ӯ���S����(��A�}\�[U��r�qƭ����[���d��f����YH�먪�M�2�ʲ�	�%�Xڈ#�6E��v5H�m�኉��P�1�\��+�"�����T* NI�L-����dmW&8�L
� ��'�Q�g��)�f\3{3�NJb�v>֣M�u�^����xLlS��b2%�����&�M��5\F��0:����TJ�5�����/]�k��۽���	uW՞�.�~Fr��}VS[!���[9�H�+,j@L��?y��e4�I=w���į�q��c�ֶ8t��gN	�E��[E)ΕV|�Xr�\���!��T�Sfr5�S�Qɞ��	��15������8n7'&ttED�2�No=���۲�H��L��R�wi]�ф�s�R�od��`�C����̛2���un�źu�q��}�!X��,��b��37.XX��ܱϴf�fr���=1��=7��D`s�}�*V@�����/����\".Y��V]n�+���J35�ԩ���B�RA��%V�-:�H�+�a�������m�9$&Us��M��uoV��ۮ�պ���Q��;�u��x�Z�;Y�pKh̉e�2h�!�s�z�\��\n*Ֆr9)b�Cxd�߽55�UUU%_�'\���Csd�n��]�n�f�A���>ȹ;�ʮ��bM���U*��j�K�.ץR�I��b,��X��u��ո�N��6���~H�V��W��d��Q1V���2����m$��oF��_c��4�A�$�8�d��"V(��F�e���bcC&��x  S�C\���Պ�yC���vU�@�ȖW�2��L��u�o�*\��K�UP]�;j��_%_N91D*�r�<+�i�K�t���PoS&<i�#0&!��`��B�v�7�j��<3׷TUw|�7,����t����d]Çh�9�z衣��{�$��SC�6�d�"������ʒ����r���=um����V��:pM�,�h!n�RRK9\n[S98���ˀYe��Sۻn�J���fM8'�X��!�&J'82��eyCr�U���"Ү&��eh�|����'-|�*��������� �ի�,72\����U$aG�\ىe�਌^����.kJ��c�n��un�źu�q�̥#�[e��*�wB:���|�u/�0ٲW�
$(�C�CFNOuk���|^R��Tb\��^�����d+�F����N4��=76t�v���S�����vp�Ú�TWz�f��[�Z"5��w]��ktӔ�T���i����b�:�V��:�8���\5^$��^�UT�Y�s�rrrLNNΖ;oU1�W���B˕d����s���<|��]��xH	�O2r��C��4We�6/{�r��f� �:Ys�(Ka���w�wap�2t�e�����n�~[cn���ո�N��6�����T$����@�/y��֕��X!9d8��ir9,%'�,t-` 8�v��g
��\�b�;F��HD�;Tr>Pj(Z��Ed�0� 5s��bÞ츞F9]�87���`�4���!��6��F�w�uj�sǼ-];�jݒBQNjΘ]pRg4�%(p�<�52\;�՘fC'��M2��4h�T/��2d�MK�'���R�Z,o]b[�7T]]����(��$����Z�~ckun�ո�N��6�ޟG�-h����d�k�Ly4 &
�l�"���^����f������3F�ي�Yp[J�:Y��&e<9��g�9��<vvrj\q��O�Uk��x��ہ�n34l�k+�9�x�b��yjt�PL��fin'�B~���Oτ��T蟞Z���l�*p|'�Ҍ[N��-�kk�	i��5�lj����i111�XƱ��11���ZF&4��4�>~k��8�>i��m>�bc�V#i���O���ש^1�<�>F��'Ϛ��k��1-���0����LLm�z�&-�E���c�nLki��X��hk�	�,�	_�Ϙ�RP��#�F�Ɗ)Y�ԧ�xM���Չ�8h���hr8=Rz����:�<k��X�Զ5��&$cX��f�5�5��jLK��<r�G�Й_��3�GC�Gc�g�,M	�(|3Á<`�����
��k��i�n"����������/ɷ�\���fe}���dF���}۽Y�<_a=�����%�xw��s��w�^>ΝDi�>�f��׳���u��[��3O�_PnW�ּ�w7}=>��k��3��ȫ{���g�ٙY���g�&f7��j���fefff9�̬̻������fVfffus5����y����n8㍱�un�źb֎�q��RѧJ��!�VV�%�4J�擜үI	2������U&-D�)wVR�kRR�0.)0�(N�)xh�)XD0�!	~b���?}��G��$jI�n�U�������xP|ɨx̒�m��7,���9�@�c
#S3�(��EI-=Jd<&	e,CI;,a�∌r,�(�0�9ܑ��%�	���>]]�Y�h��a�%@D�020�K��jMD�bT�,���mo�u�[uf-h�������⪪�J!] ~����$!�v�M�H<�BX��J�hC8���qj-�캫T�]d��'L>��"�q5xC�\Æ	�iL��Tt]5�1;1E��&��.�l��`�T��ɬ�Q����b	2!�@)!�)2�`�x�\d�6ٜ0QYP`�z���C12�7й�������&!esKR�11�	P8$2�JBYe�=��{Z��N�1�b�[��[�qn��!��M����`��8�"q�#Jd�m8:���Ǔh�Vml3](X�c%�0o.s*-��a��i�+��2Cq�5��%-����˂��Vc��D�l�YI�q9\咵dN�+ ���.$r\n�*����2n�/͠_�N���d�D��7���eb]�'5�X���J�֕�o�]b�W3S�����.�5���>���=B���;�Wh�Y��ȡ���+�Փ��C��BX�A�Xk%1#-"�O� �'#bM�X���0A����IQ>��mED]���:!�`Q�̸`�5�Z$fգq,CF�MDpE
�"6o8�jˌR�������"�	�rgй8\(�>"e�C�� o��?Wvٖ�#x�KtU��$n����CҪC��\�P؝=��0!dI�aP5.,�%����5MW��-��_uUY+~m��m����[�t���:Y�*c��ɢ�UTJ��L�.!q���H�:��B�A
�2C#!" �HY��&D�"�CV1Z�#�t�i2C�r@�$�f���*�13�CamI���j�@�dB���ku��2Ĵ�����v�}D�~��6E�"�L]��!b�/ +�j0:i{,��A�&crE,-����"g	D F2`PKИd��<z���uo�Z���:�uǯC�}	��I�Dh��kʪ�I�h�b��2&R_���t��1�������J�-�rèkpBTAa�@Qс�:�Eˍ�����2�(��)�.(lā�c*'D���u*�o
urF��Ġ��>��B�$��0!䅐�0T�L	I���*	��RM�TJ��4�Rla���LHo��c	�FN��
�TSE�R/IKA���Anc���聖#�t����y�E���8����,a���[[��uk[�t�i��uZ�$$ M���F4�ąb�nZ���DU�Đ�(�B�	��~2�Ig�P���$���*	�1��ų���Jzah�e��߮���R���)Ah���a��"&�"1˖���RUSrr	�#7��n�М-DZH��N�ؼ]h(�d�Z-��"e�@���.P!Ɖ�a�pJ��H�AI�8HM��/D^���rM��iaR7�#=u)�!D񊞉�v�����b�D,"�u��U�����i��|���c�"tO�Q���eQO5�֍j��|VȕD��>��E�.3�	8\��J��m����,N!��w&�"�m�(U�c��ƫO0l ����E�|��Kbr
�[��0�Y�_yj��!�ֿv�4�����u�1n�P�q�]s]�[������:.��њK����0ٹ@a�g�F�+9Lŕ!�T��e���R)i�ѱ a�˂��rFP��;�D&�{Jٳ�9�IdtE�@Rf�I�JlW�-|��D� ab�H�.�R�"���9L����P����6�;f����0�"}�>P�L�M�$G#r[�7
����UB�d�]4)��%��t�"0��L�j�3R`L�><p��>uk[�t��\z�)��dF�ha����UUT@�$h0�v�D]Z�L�1*�krr�R��`�5\J�GmD�jv6��G
�4��P�r�h�D���V;Đ��Jq�,@���
��7�a�&>��nZ5w�ŉ�G%�Q��WP�v<�����"���8p�f7��D^8J��(��D4b���*��SS��Fĳ��u�|�խn-Ӯ�q�ݥ�/�L�UV) �+��4	�F7K�`h�Ds[w�X��DL ��CLɑ�\J5��PC�`}�K6�B�3\[��m�c����b��b�6�4�Y�J�4'�\(>�C��x x�}ת�e@�_�Uߒ�\�@�ݍ\��x���\4	ēB�g��F�Z�f�����ѻ*éPf��Ka�c��b�f�r��EW)sNM�(}�-\�����(���8��:ŭźu�q�=k�'���*B91%�2�FY"]��Uj���E@�1_*��F˅q�2rш��Go0�Ab"0� 2b����!ϽU>�NKȖ9��.Y&}D9D>�Uj g�����8%��0(��ԝ�|�IL�$��䡒�!G
�ѐ��鲤�P��.�O	𚌈��ow��SW�l�NH�H�4@���J[9+.px�!�7rh�gD0����D6��CBb�I�-O�ޣ�4�+-5]N'���F"��4ŴŴŴ�u1ռba6D°��"Rx�0�Ʉ�F<������Ĵ�i1�14Ƙ�X���5�$ŵ�X��5X�q�?4��M���LHƱ���5�k���ŵ����bc�bcmb1:��ϖ�4�>[[Gɴ�����枦'���1:�G�R���О(��t`�~*|'�SG�|3��>��؞>(�W�4L'�0��W��>-�3S�Z�5����X��bc�y&&&��&/RbZbb�m�6ƛCc�G����UO
'���R-�Dz���bz��Z�X���{Y���CXh�G�Y��?��07WI
b��ן�o1������n�1�،�j�U&AH�^ ݓgu[}��R�I�v�a>��-Q�>H�g�¹�;�*&�������ܱb`��]ڦ�;z�^�t"�׏��Ƕ�Ͼ��=�Ԏw��(����	2������ek?G?=�����M{�/��1��2´��#��L�QS�bcU�Z�YVH���-y�L�L�;�����^�o�}�k=�X�*��!oK��;;��s�;�~���]����{�'ۜ�7��\�}���`����t����q��}�E������k�H^��gqf窷����N���+��ЏG�fw��?O�K�L�}M��%�~��Q4���E.\i�l[������n_u`uP��aΘ��>N�7q�{"Ѧ.���8��fy]���kG�}8t]���u�s3�q�7.�q�P���sc�)+��EqD)���tW��b���qB�k!���D�:'bjG"v�-�Z�v8�q8�+�i^YV (�K����B+#�5�j6I%�V>Y�8Q�l�W�y��G��1`�)��	�S�O��+��J��H���*���7mm��2�̍��I�t�p,|n��r�����>�6�9��^���335����i\�.�3=�ff�338�+����g����ffgt��o����_�i��q��:ŭźuy����p��!^@C�r�'%s�;b�"�i@R8�+	]�e��v�)����8aXG��ڱ��89[�\T���4�A��NX�4㔱G]$d��2�c��y������X�	!T�UUDF�	�V�O�:ZUe�Ș�i���[Q8Kz��]�]q\��lm��UUR����ޭዧ�V�2N�	wo{�ou�Ղf��3����Ž�:'�).��^li�d��b�L�bh$�<��Lx$t@�;
�8�F�;|(1�LN��%���7.XHD�(�����Y¡���9 ���4��,�tG���f5U��N�!00��ed`���.lCbM�d�+���|T֫��]Ա.�@��l�g�.1Z�*/�U��bY�m�9V�s���C.�m(+IIJ�֊S��&9P��J�+֯g@�ꇏ��l���-��kqn�uc�Z��������UT�SD��Ġ���,I�}A�Fꉓ0C0�5 O�Y�>.POC��E�T*ԛ1#��3),:�`�L��ӓ��2�֓b])q�)��%s
C�&�t����	?墩��Y���AZr31���h5�B��GweP�*�j�]��K�`k `���K8��C �D�G����S=����%�c�ξ[�[�kqn�8&�1�e0njUҊ5af0�*��@0쐍��0�N�\�8-I��wCI��\�<0�W�1��Hr`(��p���u1�T3%T��,D��(n��Tڥi[�ŉVS��A;oV�b8�cB����P�(�t�L��-R5�b�����>�C��w5b!Fw��R]����zƆj�B2BD=�����tc��_!P��S�!��Ň�V5J�WX����x�<mn-��:��c��:�8�����kZMkěOz�UT�}R�J!+V}7-o�������=��t�L�2��a�L;�vB�j�7\�Q6�9S�E�]Z�%vb�eyG�'��7�YF�t�(�m�g�k��ݦ����Kj:J�Uy[j���S({[A�.>�ƒ�vjb�Θ20D:!�U�CZ�L��֪zd̐��0�xF7�����R�F4��h��Q��͉���5DBpf��Z�mo�uo��1źu�q�*�Ǘ�g]���D)�[#��ˈ«Z��+,�VGq�� �!��Sb�� �P -�:��ʤn.���HO)��G2�B����Ĝc��(NH�ژ2�8�؛���m��jf��#vg��{�<��ݭMݘ�S&��X�d�dwV���f�����Է� >o&���y�{���Q+E��.��R����rT�nf�ڎ���yL��R�J2��k	@a��#�B���P�y]�C�wR��d,��5��Ё�j�hɘM�X�.3!�%M3	8T��3�\�ٲ���5ʊ9\��F��o�W)e�&%X>�ue�buT�fbX� `k��1(�/�\̝*Y�ώ�c�c屌q��um�_���UURQ[�?v��v�����1�ګ��2}C�0CY� K�qp�A���*}�̳�UY� ��f�⹙��ь�LF|%&*`�wJ�"AR��2l�Qوh�PЁ�7.jQ�BʘTт�;���"?�K��R�qB������P�T��bK��a��l�ޔ��Z�ʚ�eR�K��
�_�RU
Ԗg��p���Ξ:d�o�[��c�:�8��5�r��C{Ҫ���D;F륕������.o�
�ڢ�p�%OA)�9�B���*n�S�\q��p���dLiS��4X?}��m�Q�呷lr48��~�^{��Ӄt�6�oZ;T�R�UWNj��kCP���.4P��9n�ve�-�n��.�XK�^]QBSY��7s�7W�;x�0�>��}�V�m���V���Q�V������>[���Q��=\B��TQsX&����2���`�򪪐ܮT�D�%�#b�t�qiJ1@����X����9q!�}�ʭY�'�m�0<Ւ锢%%���.�{%̦�&�T�F��1�J��[�,�71�f$�1��1B��i�2!@[r�7<y4d�!�;4rb���9�=B!�*��f̥>0��ǫ[�c�-�c�t��o��Z�2�&L��*�+�����f�јR^\����P�Rב���|�8��?����pc0Pu�j�B���IVO����'Ty&�*��z��b�"^^[�	%n�4eQ��I�j�6�n��~{������fb��>�����]�%xbSs�x4�MnNV�ó9nV��K2ҳ��%RxT�54|Nr4��C��(��	`������4�����4�p3cH�Iy$Q�M�����YbY��oS7�їm�y#1�̴jU�ep�ަ:e�a���������׾��)�V����|�lcc�]Gx�5��T�@�e�F��k3���UURUj��}U�!su��ݕwT�՚��O|x��I�i��tp�;�ə��Y�D�!�Q�;6�x���(/<JJM�ɠ�6��ڱ�3EO�}��n˺����.�~	�d�b���G#������yO�h=T0�ʆQ��'�[Z�r�G���};�уS�\�)��4Ĩ��#�w��+�o�~3��LGS䯓����F%�ыi�kщljұ1����%�o:�OX�LLc^$cX��X������ZLJƚ�xƱ��#$��X�Kc^���ш�Zc�O���~�bz�#1�Lxǘ����5��i��i0�Ʊ<cX��XƝcLE��"Z1ֶ�ޤcmV?5��=|�y��Q�:|`�K�C���D�D~K���-xO��O��u=G�F#�4�8������)<WG������x|p����%�bF5���-�i6Ʊ�LԖ������lki^���$�0�$�X�F$LH����b1=C�0�O�}��/�}��þFs[��q��x���{���y꛺󴙎̋�V��o����I����v�7��݁��\K�AM_���9Ǭ��E��Ws�����fe��g����]-�9w������fe��o9˼��ffo33-WKy�]�ff.�[U��s�y���N:t�ӆ1�c�:�8��8�{�kZֵ�$V5�m�$�����r͹#p�`�b��B��|,��km�WuV6V&!��0���U.|L4l+��kc�$M��¸��	$M�{�i�����'~�9�X���*3P��F�P*\��m�)<=�>*�*��3(���:vV���f8J�Kɨ\Ǥ�j�~:�ƞSǫz��6��q�Ǐ�����!�e�#*�'�Z�� D�Ä�hr���s%÷��W�����G�2.A�,/ �[��d���5Q������%X�p��˚NF�(-��m67�tØz��Q�MC�)���h.ፙ,>�έ{�W��.����(5�m����}8r|'K�;��[���k��4�Hӕu��Lc�|��qn1�c�u�q���ؚ�i��!�ckW�S��'3&f+`�1�T�����;�4f�tY�2cC�`<CU���CV"��rܗcdFd�Y��l|�#a�ڧƄ�dU����r��qWy+q���"��B:��c"���*���UU r�g.�d�3^�H��o�٘���6,��I�ɽ�����p�k�6�am�`]>>���H�����t�"D}�t�n�BB*y�Q�4�>�8���8�Q4���`9h+�E5�IUI��a�-����:x��,�.V�L5t	Y�n�z�Ӂ�u,���/ȴ����gC��Ķ��U�vAdXq��)kE
ª=���!{���yM�V�'�Uo�[�[��:�1��e�m�oɨI����ZҪ�;[���D�9II��_��/Ga�F���~0j�N}FU*gP�'�g⟆��R��&憋C*J��N�������<�RLp���v�ə�y�6-����>��������kO��O��Fc�����>jH������5��o�>c�c�lc�YkG[x�7����*M\F���e܎I#Ww�UU e���h���Q��iUVE�!��,ߗ'��,�t�*��e���C���a���m}6Y�Q��w�ST�j�BF�%�G;���^�Y�~檠l\�%�坚��29�p�=N�2˯����@��|x���*���gܢ����4bn��]<v�ʑ�V��8뎱�ص��,���<X�Q9��%着�@����5Z�	���r��aS�MC�ѭ��&>���Gtyi�21���d��0��t���Iu�=C��,MYg�����'� ˌ�2fjYe��i�%l,�͛1X��s
3�B��}l)���M�"3�0YE	�(���Sf�����T�������9]SM�Ž|����&&0A:h��j��pԭT#�Kc�LT�JJI�9m,�˹��)5�f�S5�,qF̤�F���W�M�*Z�j���j��U(a�f��9�Iٹ8�'�&�����um;��U3b&w3Pj��b��!�*��(��cʃ�Y��UA�h�h(C��������SBZU4+R�D�>�P���K8f)B}&�n5�L�6h�h�]i�]�֫�lY��#�J{������.���uT'�c6�FJ��,n#x�6z��{�,���+q�zܯ�o�돜u��1��a��:p�a��d��J`�9�*���������;G�C���4p��e60���ۣfN����dU4Q������5}���2&����]1G�e�����6�,J9��39>.�
9K,G�k��yd	,+�Q;i#�&�1ƛj����"&
1�1�~S5.ׄ΃	���rNlt��pM��G�r��ڮ�����u��bϏ��><<C�/ �!z���	�%���Ș;��[m��`И��OLC�we���<X"��2W��X�͇N|�5���`(g�m�%�֛�V͞L�c�|YeQ
2��fA6Q��&K���	g�ơ�\ѣ�����Ub/vdMI�a�`L��:,�9
>b��K����G�g���~:l���c�]:�8��7Rz���d�����ɜ�����{�UV���ڢ���c=T��Bb	�(���Ye��>.�-�	,[�5�BEQS�3���|x�ga!�Y��e�4v(�4P�3�92C���n���CEC���78T0`-��?\SbCD?lMQ���$�vyU�6]@ѣp�'�YVS�W��Q��z��i�q1>G4u�:�KF-�X�b�Ĵb[�1-�"[ŵ�k���0�Ʊ<��&&�kI�5�4�xƱ��&#��ŵ���l|3g�2x�#���|8C�O�5�����X����0Ʊ1<cX��b1mb-11-4�c[c_������z���'�cƊ<%.�Z���E_��1��I'�1O�X�N#���|�C��q�Ԝ~k�Čj��[_��>8W��°x�|>(��+�Z���䘖ƫ�mb�q�[��=O�aFT����H�O	�g��G˂��*c�G���������EG�=�תb�js#�����i��cbn��v2�*܂9���^��t�ks��Ra����U �ə���"c��Z������M�Y���ٸ����;�C����}�=��a-��l���zSͣ��{;ߠ�������2��Ϣ��1�dY�ﱫ�'��p�����Ko�*x�q-�ʍ�/��&}�4z�[~��Q���2���v-�w�mU_�ޏ|׳�ڵv�:t�qM�O}�?�3~n�����N緞��/b$O�e:�,�+��{�_I���'���ط�o�;�έ�&{3�����=�k;�9k�S�u4�	��j�o��׍w/fb�%X�z޳횮�>�Y����ǟ}ޯ����{>��F��__om����
�]�I������u�܏,�r��ߦ������>s���L���羟kAǩߖCf�_���?��1�8E���vGyj"��,m�%���BX�pvQ�%8�v�'-m� pM24pClU�bL�
�A��u�(�b��ۃ��n���I*��¦ա�!W�USƱ7�[n�p��[,D��遗�><i�Z�i��rK!,lvZN�O+��ʙJ5��5��!+Z����o�j�[���fs332�36���r�331mWj�ۼ�/3�ŵ]��n�9y����8p�1�[ź��Q��?z����������b��U�m'%���;]�C��#VX쩧��m|%���ҴU�R�\C$MI/���C�:�2D
�bR�'	c���$�E����
ڑ�1�N:��B�(�d���v��rQD��jQ�n�Z�M;�Zp傃��9&e�"̮=UUi!��[}����Z�Ȑ�f,�4�����Tʢ������7*��ȉ��,�}B��Ѫ;�ȕ(��C�:U�dDϢ�揧}U�rz2P�Ը��1�0z���};��B�«b%Jˇfz�pd�S(ؐ!���!����˻��٩�|���&�M�V(�V~�O@���c�,񟎞�g�%LIBbQ�dko\|��X���qo��1�uӧHp�c�>��P�I�n��`��*����
�f�u���{۹	wH�����;�TOCSS&��^e��䁠4l�hN��!��d��zT�T=K�c,StP�%*��'Ff,����5���M�Dn睱��@8ǩ��-�ρTxtM��3.r3aTD�g��4���	�0CsJ�|2����}�����c���b��-�N���/ �Uv���$�{��T���+�`��&�F8�agL�U�C)�i�(0��Ȍ��f��*zPP���C�w�vj��,̬�Y%�%vg��L_���P��<z���#
�g��fX��a�fM�9%LB�bbjxB�`�m(؝�H�NJ"���V��G��~�:�[]?=�c�[�:�Ǐ����::C��3��f[�*����Q���tH�dܣfYv�G4v6hDM�ݻEKi�ʬZ��J�-N�5�B<�qٹ�l��按�Cp���l��'�O`��䌩���J�Lѡ6#5FrO�m�t56q9�X�#�n};(��gXZ���[�ʔP�XC��(�9=��Bk�,Ģ��޽Wˮ�����mn:��c���^^B�����+h��*����<��#��)���Ac@�g�f�V�V�*��p&��(��q�L"��Z�AZ��q��ѫ+,�V�`�b�X�H�+��I	�4u���a��ݿ��<_}{����ԉf��lG��.��{�;�Y�����d�*w1�q~B�O@>����dLA&狇��*tщ�z0&��(Ɯĭ��21�CI.;c:Y�(Й��19�4���"��s8L"�.�h:4�,�Rr�(��֊!O��� ��J�,�⌺������9U�4x�m8at��{T�V���'�r4p���ط�-�c��u�q��$�iR2j%�B�$3�,�h�l�4�3ӌ�im��V�M�^L�E
�=(�x~�U�X�DA;3.>��ΆN	���3
�3֟NCG!�]X��E����$$Q���A�[�L�ժ&�.���N�ϰ��(D�� ���lԛ�C��B��a�O��4������c뮝ul�A�=���*�����Y�ժ7ɵDX�`ؘ���l��(�8"u̽UU���ޜ&���6䢎��o*hY}��6�m��Vb�x�l(ɨ{�&�R�C����J(՗7!D��ke!�<�B�e8pd��PԔP���U����""v�*M�0B��yv�Lc��dٓfK&�mn:����1�:��Q��.��0㐕$��j��$?Y��Y��Ȉ�,��_�0hMv��gZř| I[�:� ʚ�Cg޳hK�>,�;اM�Tѡ�`��5���}"#3��b{�Y�6�����~�e bj��C`iV=���(�5�YF .،�0P�BY�;�h�f�8�n�o��-��N��6��}�s�*���Zt�?�f,mJ��m�+j��"�8M�*�-�V�Y(�!t9�l����`q��%�.��,��I;�s4��i񥽷u��Y{:1w2�NnuD����7:*�s.�˳e���y�v�]�E�**�WB��͚2!��s�捐J"P��r�<�N�S�rn&���`L��U����U%�{�E�]9��&e��a�D��#P� �t��Y�SB?���G��:-v�e�s-��w�����Iӵ�X��șo��O�}*�����ξ|��Z�-�[���:Ӎ�y�En+U��"U�SP��њ��/j��$/dZ>0D>�,���y��]c=~s��J�~G��i�l[���B'$ON���5f͙�*\*0�&���nF��`����W^4��;�F't;y�|pM��Xh�8x�L�P��L�143�~�)Q,��������V�u��/RjkJH۬[�km�[�un�պ�V��[�[�V�<Ym���:hB�H"hD؝�'����,�f���DD��L�#$Dw"#�<""t�4X�&�؛4&��(J!I$���4%�mǍ�����X�[�c�X�0�4``�DM����"'D8X�l�AAJ)�6lM���rUÝ�r�|��eE>yϖ��(��Ţ]7�?l�4��?��&{���fs����=�𳺦�c2�/G���U������C��}���jt�.G��ۓ{����~]�o������x�}դ}�,��~sc��B�Sfd�'��A�K�c?��g=��&�O=�3��Uv��r�333��U�wy�����^+�U����ffff<WJ�wwy�͜6l��`�&x鳧HtN,��hֶ���C�h����i����j���/�~t��_�˶�l�vj�	�;�w�W��;Z�Q��x�I�v�H��v@q�7ƛ�G���j/�S�#<pM90B1ڴ���0!��0�1ɨv�bT0`S�vw�Ї34#'�0�#�����fn	�ϟ�>m��lb�~u�u�+��to�n����J9F�I2�n�3�39*p> �&��w��!�+�$xF���g��X��U��O�n���1�L����?j(/�넇Ԑ���"��i�BsB��`��pѣ��E��&�\є�6�	�7�IEӗAt��ъ��n���������h�9�MUw��[e�p�br�����:���u����lb�~u�^Muo'��#M�
Y�Ҧ�	���j]3eCW��7�
���ۍd���Ԗ�%b��"�:$m��#�����i���'�t/+v�m����y	��|�N�~Su㵽[�صm������L�[�2��un���i���s�W�y�}3�����,M�1�m4�>8l��+����Ҽ_�J9�3�a3,ż�o*��'��=���Bp�¡�ԋM�4&!�T�	��/'��1ؚ���d����.dȌ�n;�2'߾��ՙ�D�2!�w��#�^j�Zi�b}=R�|%���X���Jn����<|��ͱkb�ź��:'�;����r��1�<���	y�Z�Gfxx��,L�3u���j�a���h�>�*����WoGeM1���?"%xj��ekm"��<3b&�tɳ&�5L�w#�ɑ�U�5[�w)+��&�x������h�q���pЉԩ#5X�pX��
J���h<l۴q���ξcl|�X�-׮��D��u21��ٜ���kZ��Cw�յ�V}UUi!�@�m�W_I��,�H|C���Y�	B$3�r�C�Fv0&�=���fMMB���;xiqWmP��7E��)ʜ8/��),]����*H�,�B3=1�~�ep*8P�g���0dNe}�V˻�]��af�H�LA�@�OC�a�(����畏͵]S��uŶ��-n����:C�p��{��j�o���$=G��{�j|]�\?1{[!�`?�p�2r��0"9~��M���!�8(����M�}3'̕DIiٱ�קg�&�S�!����3��2B�MB����u�U��7g��T�롪��3�Ț�]�T��bd�%K��9���3�CF��)V��eB�	�F�:Va�-��cl|�V�-׎����n~��SFܒ^�P�"lF,�%��!�t�3y�)ʌ1��b̘�ә4q����%�@jcjW�NY�r<�m��|hZ��֒��c����;��75w37	��R�ٳE�F�ky&�C�G��Zi��!�B�쫲�x^�0'����FC�p�*�M�lG���F��aG��.}�:���b!C��b\���0�
�:v�
4�&�Q���dș���\����с���K�YrZ���-r��[9G�Y�g�J@j\�������FO�8|��c庶1n�u�u�p�Ud��]Q%�uUU��hK,�J,��Vu�xѪ(I�MO���K2%��&E	��χG��1>�L�h�,�x2a��ɢ�'	FHt���ōD+�~�����[b��굺JӣSZ��\�����{���	�;(Е32VLC'���cI�\ލ	�)�=�x�ZV���:��?:�z�ͭ��>[�c��]GZq��\��}o|UUhOt��3U��V��6$r@�=;�,�|�s���X������������vA�Z�X7yn��&�u���9�4p�F�~/��`Yھ�j���7CF�O*=�A(�`4��3�N�.�5i$a��D#�����/N�[�]c����[�^:�:Ӎ_s�7�~�_��q<���J�q��ؚ��Bn���g��M���30�x���O����N�}wV?^
�Jੋ�WLJ��|d|�'�A���كA��d13��AeK���X�*��}�<v�6}�>���]7w�х@�l2�����V,��7�`���Ԗ������e�4�b���������ǯX���uŝ�D��<'D�<tN�P�D؉b%�4 �N,K�'���؉d6hMAB"'DN�D�"lDN�:X�%�lM�BP�%	D����'D�6%�"p��.ĳfl����-n�Ɩc�c��p����K� � �"%"lM	b��{Z�V����&�f���i�u��u�涬C"֊���Hƣ�����9 ��X��h��]�u[�+&�O,��Y-����n�O���	���,��������<T����0���U�(F� 3��N��:�m���1:��X�v��⸘��eW(�����)[X��y܃�7׳mT�g�����/կ��f~���v3f���I��Y毻�����;leP�>aϫכ���S&9{+{~յ|t�<�ӀڟV�p�7*����y	*o�ۃv,��F�	53�s"��ڌ̩��t[[k�rL`��,�B���ւUX"����&�;c��[&)]p*���$��S�V��YSv^�*���'
�֯-�T
��*���bf8���PAv��JW TX6�U�W�r�
QƇC��H�� ��m�0���T�B��'�J�V��i5���z����k��x��V��󙙙���ZU[���ffffb�iUn���33331�Ҫ����gK:p�Θp������K:t�DᳵX�	�7X�r� ,�(� �+U��+e��(��늨?Ip]���6ݰM�S��rK,��ǹ�0#�j�i��jA���R7%cp��:�e��-'kܸF�,#�9&q��Q+jJH@�9C�r	����dQ�Q2'�k3�����h��jд�f1w�UV�޷�L���}�<~�9g��d��Ǿ&Zz�fٞ��P/to�܄���+�I���C�(k���L03ډg�'��]�t�F�ǩ�e�S@�ҕ]�ǐ�.�S��юEZ=&P��nfBC���9��.�ڞ���ÁA��
�vaT��:��!��H��iQ��,N^EYx����ܦ�t�� ~����x������[u��[�-׎�!�8lp�E�հv��ЙEѺ�	�������:����U!�µ��QE��2p��Z*�O��	��v��
�9G30�d0p@����_�4ϾUWZ�Es0Ń�&�u��-t$��Õu͖Z5^6k��LX����6�ͽ2>�C3�����`����kW��2`Ƀ&:����Ÿ��Q֜m�_L���2�%Ea|�UUZ�>�W��郈�Kɔ4hMb�|v6	����12Pѳ�E|5�l6bn�Ôk>���e�S���2�"��������7d*+n�H̉��p����N�N41l(c!�<u������asf���y��B��h0Q(��������
���Xe�G��l�`�\�r��p`�������O8YӤ:'��lb&+�UV��-l�e4U�Gh���?!g���v�3.�8ܼ�p�ln���d_]��fY��9��1>~�ᨘڞ�,8x��E�f`���Lr}��C�!g�ɐ���%m��Z8|r]����03gE�Md�)�ETt4H���N�SAg#PN�7
�`̀��T�f��
S&�m�X��q�ulb�x��N6�:�ߛ���ø����3e��XDQ�,l��.7�1J�'�����{[�)+ʦ�c��mɋ0U�)!i9c���f�+�u4�2��ʙ/$����UV��Y�_^�z�y�]C"��f#1�|i�V�ǚ4�{w�{ӗxT�g�$��}V~�Tv����46�z���+�i�i�O���h�`�s����ς_�,֑LN2Ό�X`�;�(��EV�[<iS}\��:l8y8g��2U��th���q�x��9y,���h��a�Mk���)����ط�V�-ǎ����c^MF��$����K�sY�UV��Er��!���3鿻K������Cz,0]�.9������U1-.��fc�6��v3s��3�U�ER�v�5Y �����Ɉl`�<r����>�V�u�e1U�+tRE0���t�NCBX��+�[!�Xh,m�zjb��ɓ������;uŭխ��i�Q֜m̩!$>bs}UUhB�%U�D?]eBm�xoo�m~?:#��v�f�5Q�ͪ�w�:kqj�$�*�F�G���m#��,��&��:㼱Y�B6�V�G㧍��m�U֍V����K|�k��_�Ԩ~_%U���5�ޓ�Z�6{�AZ��p8p��z�5M|�&~|��mo�����g���˃!�Iޕ�e�7$/QF���uUU�8lʪ�&����Ü�ID��ǲ|q�!���X�@Z��<Z���2�����P���b�\��%�:v��&$0m4X.Y�����29nRa:�y>i�C���97�w�pt�l�2[�ܢ��`���L��W%��L::8�n�n��u�u��f����si�Z��O�eŒ�7�rbu��p����,�b�u\�L�Dxl��DC����Oftp[��jȨ?G���)`GaWј��8�G��lVݔ��D�+ �ڟ�m���|���� ��&��E��f55�-jݖd3RJ$;WN���:lў�,4z�n�iA%u��-�U���l(Fz��Hd2f�:f|`4h�QG��|t�Q���Qp�ӆa��k��5\�o��OȖ���m�j���ON��¡p��A�v��`�n���'�M:����|�V�_8C�HtN!pw�i�d�����:��Л��U|l6}���,�32_�Cu:}4u���1���&�&�'I��:��E�D�d��Tm6��(�trm��?5�(� �ۥ�M��\�G�0�����Wq�O�jd҆�����<b��$G�������x����[�un�պ�V�ֵ��:YB$b"'DN� ��b �<'���&�؛4&�""hDD��B�DM����"'Kı6P�6ɡ(J����DA:%��Ŗ"p�!e�f���	�0�O	҄ ���c�1��0���0��,�AD���"hNh�+�Nl{�=�wV��{��}�_y�{��$�0A��-��p9��(;`&o|7�}�}[�s@��������Uk��-�b�>��ߋZy/^}�}��?���'���+�ϡ;�}�۽>���u���?�or�wݿ-���ٲޫ\����������}������Ӧ�K�l�g�Sɻ��ŭ���rHͯs ��}z�ޒw���z_5��m�w�V���33333�U[��������_1Un��������|�U���s'�,�Ç�a�����:t�D��k6�����\�����$����boK;b㦒h��'3���s�}w�\]ݘ����k�Ù��3�Aɰ��J�l>�2nvns!�S��_Y�A�u4�O�C�SM�W��������|�_1��uӧ��Âp������V7�������{�6{A�%���̄�K�z���mQ�ڤ�bR�"P,/8-b�Ės��Wd���Q1LB�$8Q�t��>�5��\����Av틸a�����FCf���䁔�_�=W��{�kM�M7]z����|�庵���u�u�I��^s���bvWe�IkA1d��"�LQ�+�(�N)�+��2fI�̵[�w"��8%[�|`��XS��%"��-nUZ��J�R�"T�r�K�Ͷ�o�'WKgL��,�q�yo�j.X֎�[t����ڋs/P$
��[��Y���2��oՒ����'�ؿ�1�4���R�g�3)yUIT�gey���ћ�x�B��r�X4�i2m�G�4�����Q[	�JGֈ໷l�LOtrCǡ��A��ӆ�6�ؑ����κ�庵����I��D��Լ��~UUh�Cjr36)�2|O��� ��_������a|�vQ���Ht�y�5�5��ԼiN��Fh��א$���a#Mv(�s�KZ��ڊ1s;5I�p��-W�!ɺ�y��KclS_C({1�|��V��V�X�:�:�$��<��2Z2T�	�v�����?�a+�{��H|�=��f�U/��^�c;��䵿�g�>6x�_��f��s���RFYC&+�ȕ ��BaQ��F2�c�D�������r�p�q����M�a�f�
��&��C|q[���ח����NS{4�5M����u�x���9Oclq��\|�V�_8�����6��;��k�����p���͇�G���=Y�| �Կ�����A�KB?UŸ1s�l^�j�涢�<'�.���b�ِ��%��Y���$����Ly_�)o�-�u]�2��nI낧�E�1�RÓP���>��[O\m�X�庵���u�u�I�xm/�/V�����lp�m0w�#�"s1���P�v��v<��j#S�Z��1`�b�����cP|ad+R��J�3�G#�0��ʕ�m��`K�UUZ7G9�}����31����4ޭZ]���s{�6^nkF��wÆ��C"��Ux�er*��[:�ĹG[dးI�r�Zn��C����'&�!���溾��97'�J9l^��v��h�Rr���k�v������H��Ț�Ƭv1�����x�ȸdT���V�W��].�o1o�[�[�[��G]GZ�{a d�%HGj��%\%Xj���ZUQs&M9Ƃ�˷0�Mɰ���3.l2XP{�Z5R��X�v����pw�9��|;���U�Lbg�5�$j,v�KdQGg%��UH)E¡Ṱ�s*��y�o�S�Q+�5@�EF"̯ߤCG���X�\Z�Z�c���\�nIr��C��w�UUh��	�8v���f�����2`ܩ���tb�h�>�m�z��Ͷ�V��q`�.j_��.7��W^��ixL�ā.�K���S+!��Č�4a9�AE�I`ӧy$�L'T�\b1�-���|�[�[�qt�G��%XJ�^^.dv��ЖI]��O�������B%��G�}��C�����
��[Km(�*��Н���aF�;���ِ�qx�K�C�E�ɒ���k�YA�l�L(��T��qTWa��a�~tEWF����se�w���������:��^��8���t��~c�hO<'���"'�����M����҄��B&�OB"xN����6&�	�""hDDHxN� �O�'�DN�%�blM�6&ġ(J#'����B ���:Qb'N��Y�6aF$0�<'
D�"lDD��Z��8�c��L0�,AD�4hDؖ�f���54M�5�5�\!q/W1��x�j��*�I���XA���HD�Vcd��Ci�<�������+�O22;���d��u𢛒�A��u0)�/�ۭ�B��"�˖`�1Q�aimn��i��V`F�k�����:,�c���=���l�\f-����E���1��o����S~��́혾qg��0Uswk�뵷:�÷�ET;S{�gyML��K0U\��s!,�rA�/�����k��W�OG��r��Z 	�(�쵵)����%�/}v��ӵ4^�Y0R�'0�	��Ř�ۂ����93c��7-Yq12�(�c$"�1:�|����A�#�¢�ʤCEr1�FEEHT멑Z[#��!JDʚ%vKtE����"T!
�Um��+l��ȯ:5P��4����+S�8�����< �	���X�C��3(�tj������u����e�2F�Cj&[a[Q�8*{����ɞ�ￔU[����33333V���������EU���\�����QUn�����6�8�����G]G\,�>I*x�Ǥ1�5i�����#��9��]xBǎ��« :����m�rƝL��m�#q���
�$����0��1�h�j��-̛Sřx�VFKƎI��R:)%Q�W^�6f�V�L!�u������j�<yUU���������7�xӭ���囗�ku��E��Ӻ��1f�9�.�0b�9C�N�����D@�����ɥ��r�!ӷX� �M��\�2�%	��B��z\���9�!�v;�����M5R�����罹����j�K�}=>4���m�|�V�_8������2r
�U�D��.�f��IG�F��
5���l�nTca�T������}<�g���O���щ��T=k��K>������ƘrY�T���+�0�#�Q�J-(�h6bs�{���0K.v�OIG�2$�+��}�M��V���庵���u�uǎU�i��*��U`��؍�mX�gf�I��&�;�v��I�҃�⍆�3x�2XrtLN��S����ݥ_0v۱Z�ߘ��'�P�{�{V����5\3��es�V3�3p�3���J2M%�y�ː���tɼ�A��^�|��ط�V�[a�Q�$Te%�Ua�:pJ�L��^`<���C�YG
qZJrF���}�R�նۻC��������a��!��l;��d���286 aD0T/g�j��|Ν�
���H��h2t]n�$?RCA��j�ɲ��r����X�.p�����l[�[�[��������:,�T��D���cY2G'��S�ז�I5�"5�T(�V�-�ڤ�̷^�h#U�)�ڍ��⩡0'$B8��ܝ� ��+� 8�[�]��{�ܑN�;�N�̽ћ�����oTk�v��u�����x.5B��&���t�1%MOO������w��d��|CP��ɼ����1E�'oF��*\�)eeG�,3L��W�,���*�Գ�V�B�g,���b�U�'�Mp|$��׏�q�θźt��G�����%�w�V%%4�d�5c���q̔�i˼nY
��C���*K<M�
�M$�_ED���((:z��<qxp>ݵ�b�8(;bV���q{������7�A�	���wtPzfjN�U������z��J[奈���#~>~q��Z�|�V�[|u�uǕ�=�Gl㣃TI_@�q�x/����]ɿ�3<j4��6�E3��so�N�M�M��%�rD�B�f��3�E$��B�o2�X�C�<�d�v�T7<n>*Y��"zb|�:�*���f���`30eX���2��ܤ�*�4�\�������z�����q�uku�t�6Y�Jd�5%"mUa�p�P�7Rk*���)���y��X�\u[�dU�1[�'�DJ�Y���h�}.�UX�{'!�9�3�pv���n�6{YM�d�oG5*�Ӕ����q(�27>5��d�fM��jh��ȜcUuA�j��*jp��8���N���6�\b�Z�m�]G\yS�i���U�d�"Y)r9p����N45�IIwp{Rm�7P^=4��%q��Nczܫk-���qR1GU��I$��T,t� �ZҌ+�@ހ��;`�+j��=�=s-���`veո8g +y+NW�ܪ*�`�B���Q����4Q�FtGf�Bc9���}��5LL��1C�1_"�=����j��i��dr�5�4j����AW���TJ?W�Ca|0��d�rV,̖NB�B$�s�Oⱶ��딳vN�8L)ӣ�4�ђ��lm�q�uku�uq��H�T��v[{�����[Ef
��V�9y��US�;�������&F_ն�[��!t�����F�Xr���(ٶ,��x�:b>�2a��|��o�n�+G͟*n`�s!p���
���w���(����ƴ4�;C�U�����ٻ]�3�Ǯ0���o�X��|o�q�-��'���xO��:'K(DJ6"""'JD�B&�D�<tDD��:%�6&�٢� ��Ȉ��8P���Dٱ8"xDD�bX�&�١,ؚ��2}ϙ>Hl��8!k[���=x������1��a�xN ��"%��<"x�����=<a�a��[��)�|��1�Ew�G�:Z��{�M�����Ǖl�v��������ʹ:���~��D�]��Z�^�f�g��c��z����bx/x�//�e���Ր���yI�]Q�_;�ݖ��ux��ߧ��~-��2���=���xgw3o=����sZ�I߮��}X�M�f��e$�<o=��~]��םO}x��U�x�yI��Rd��gյ�����v�ܭjW;~�����u�8��{��V���\�����EU���W33333Un�����������wwk���m��Z�Z�Z�m�]G\x��$X00t�ј�eA��j`��7t��enhČ4�p�cB��.-J����˰H�e��A���hur�l3$
���fe�q7գ!���&LSIUY�MI�aȗů���>;.���m�n�󯘵��>[�t��Âp�a��UV�\8�r��\h�0���Q�Pv����.���+;l�i��Q?��	��G&Y�o�����fT��<U����Z2]��ۧF�L
9�
v2���a��gzO�Uc�
��!�N���DQ��E6L���M}�ɟ���gnCl�Q�8���=k)�޾cb�|�V�[|u�yuE��Ux�m����*vW V�R8E_+���dfR�c�D�,,�1����3�br��x�lQ�m���Bjڠ1�9j���ڥ�� �$���~ݺ]{�eڜ��c�Ĭ�[�9��[���Dnp���'.Ë�	�l�VVp��`�d��S�C3�G|���&�f�X}O��j�
0c��,�}ݞ�r��a�`PxP�УAE�P�Z%����v��m��%R��� QƫP#���P���pB�/�\�z�z�玱ն�\b�Z�m��Ht�u��J�Ua ���"�:T�p������jå�(�A�R�s[Y"ȰHŀ�TU�јl�u~#X5f�!�P|���7�Z�O�P�����Y�	Yx|���iÍ��ʋ��G�#�K�a�>�`Qp̯}4�)��5U�h�/S�n�����ʂ8�';(�[q�n��\b�Z�a���;���!_%p�MZw���|p��c�<;����	�����NJ5�%#�����gMLиЉ��������deFY��iѮ���J�5T������j�ewq'tY���F�gL�6oe�*'{�`��.���c�co�������#f�(�h{-B���J�7�u��4$����٨r:fL8~Qj5f��"$�\�++h|&R�ēL�����+�e�(k�Q��S�Q��X�=�l7>��/�4�Z6H#橥ixb�CF�3���g?N��e܎��WO�������57>�Ypİ�f�<3�e�J9�ǔ�6ӯ�|�ַ�V�X8C��'Y�z�Zz�"�u[G`��7��7,*2c�`�~�P,�`�!:e�L��##����5T��[hRԅK�Qt�:A����V��[n� +���~����4n�ws�aw��&m��j+�Խp�a�מ���B71j�G>��\M4z,^��EJ�!��JJva0�t�U��US�dN�7D���������S�l�E�6r��C�Y��(r�$_�L!gn��r�}�w��Ż��m+�Ӏ�
�P�o3�3F����fM:x��Ǝ6t�æΞf���$i˵dmR街m3
�=�;\�2h��*�\V�o�)�{��%��߿�H�r����44s�j�t�d�I�4pO|Z�|���^�褕1$v���8䪹%\�m9V�	u�>2��w[�b���Maf�fy�(�����B���Okׯ+���|�q��V��6&�f}����0P�Ubp��sй���2��a�
�*eQ��b�N�l��"���o��k��Xq�2�V� �a1TU��%��fMό��-��<l�j9ph5�2�m�3�T2d�����Z�;�T�a�`�,F3lT���>��ckcm���V��uu�TB���H����\ g�Ab�T�y%<z68����/�FH�U\�25yB��ӑ~Z�j�p� �������.l4w��3��tL�U{;�e�����䩱8a~������Ѽ0���ԗ�Fd�f�����.�{� ��<� �B$�I$�I���4Q�K���ϫ�PI��['4QDA�QK&'���t�d�-�R�� ���(q T�$bA�H�8�D��
0A�0H"1#b1�F � �� �b1$�A�DF0B1"#�"DA �$��������ȒF1F$B0A��0F ��D`�`��H�b"0B11 �#b"0A�0A�#bb�H� �Db" ����A �FDDdF ��D��Db"1�����A0D�A��0A� �F	%
��DF"#�DF �1�D�����D`�#D`��DH1 ��bA��DF"�B1�#A"��%�Db"F� ���"$� �`��`����Ȍ���"$"2"#DDdDH0D� �DDF�Ȑb2"#b �`�A�#�"0DFD�"�A"#"0FDD�"""2"Ȉ�`��X#A� ���"0F�0DDF Ă#A�#2"$� �A��$"#`�#A$�DdD�"A""0A�"1�#"#DF��"#�bH��$
b"0DF �A���F��DD�`�#D�#�DF�Db"(��F��F"$�#Db"$ADF"1F!��A��1 �$DF�1F$���DF"#� �����0DF"!"#���D#b"1F"#���1���D`�""A�"1"#DDF�� �#b	1���$�A�!wA.B AT�EHE�EHQ�AHP H�� BHU T�ABH%(�UQ
�G��)T�`�H-A`Q�JR��J� �u�x��,X�-$����D�@e%(�PA*�)�����T��(A*��T��(�U@���! ��� �� ��"�U ���!D� XT�D`B
A)PJRR�B�TA*�%R	B�	T�UJT���E@�R���"�"�J��UE"�EJJJ��R��H%R	MRSB�i�) ���H� �A`�10@D� �`RP��J�R��D%B!)���%!�J�RH!@ �(F!R��D%!�P�H ���"� ȃD%T!
�%�P�JBR��!	P�BR	U�BR��T!*��P�%T%!�P�*B��%B�P�JB ��(F �D	J@�%!JB�PD!dA�b	U���!R��% A ��2 �2!A��!*��P�B����"�2 �ADA�dAdA�`�2!DA2 ȃ"�" �2 ��"�2!T!	HB��J��%CHBR�D%!)��B2 �`� �@�
���J�BT*JB!*	P�%!
��T%BR��D%!���J�!*	H	HD% �P�%!�HB	HB��%!)�J�BR	P�%!�@��A!J�j�J�T$"	P���D���%B!R��J�BT!	UBR)	HB��"�JB!R��A*	P�J���*	P�	H% �%B!*B� �JB��T �b�b�D �D ����
 �# � P�B��!FFA�	H% ��JB� ��"�����%!IH%!R�JB���%!R��T�"�B�FA��� �#" �A�1!�� ��F! 1bbb���1F*�� @b�FF�P@b ����`�1�)!R��JA�Q�F"(���`�`��%���� ��D ČB0A�F �ČH����h�%gخ�.^�R��Bs�N��b !$������ Ry?e~�3��5����yS��ҹ-�����\�������������;uمտG�g�1����׷>��m�Ǐ^B�<�����}��v���w��Tv*�����ݾ | ?ރ����	�/�"���4�(�~Bv��>���C�H`�bP��'���!���y���Cڀz�AT��O�|�~�T$����HX|sH����w�{r	a�1=	���LJJO�k�^�@ן9�Mx���^b2fw\��p��%�! �}��F�)�R���aE,�b(��f��
�"�$ ��Di��� �m~
��3��	V���}���|�������T(�RB"�)!*���B� B * *(2��}a����M?��k���G��G�>@�W �����������-2�y�U��hQ,�Ͻ}���^����z��N�A����d7r��G��}f@􇕸}�\}�D�g`C���ú��q�ߪ|Ə�O��*������~����W��=G<�9>�{���7'��PU�<��V+�>�(����0�F�n��p};p�SF��u "	�^B�Y�G�,�@P@���|2x�0�� X`s�U`i%%�)O�Q/�9\:��6#h,��z\^	�x�����`ﳿ���Fzr���*��~�~�>	������_�}���=l<��"}�,�l)��'��zڞ���|ޯgC>p|�=�?����/p�%�EP��j�|�+�����(*����9�����{;�g`w��/��g����$�*HB�y�G �r��g`�W���A���ݠ���lKܦ{�����PU�}�����SI�G���E�.�P�����tyjq�O9
�K�aR��t����N�!A�S淬�
~��	�z4�'pw%ҹ������g3E'��u�0���+�C��BH�5����rE8P��kR�