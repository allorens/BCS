BZh91AY&SY~j$�	_�`qg�����*?���b�  ,   (           P      
                B��` @   �    J               (           ��*ER�*%@T�T�"�eQ�R�"�JBJ�%%�U
�IUTQ� �$)%	%*�+a�H@� �A�Q"% *	)%k0����;��@�h���@��QE�Qn�С�F�rsb�n��Yȧ&���@  ��   ҟ}`�zy �B���s ��ԡ��(=�QJ�۸����T=<�P姈j�p P  �   }�T�$�Ԫ�MaJ
�B�������<���zހ(]� � �Xy�@�@n� y��X <\�� 	=�4)�X:�  �   �S�[�>�� q���=q�C����w�=iŠ(�)$p���t�n��� b�@x   ��  ��J��PU(�UEH�J< >� 9���C�� q�*�WW�s�r5Aް���t�'@��B�[���t*�\�  |  ��1 <�� n�EgҀɠ�U������U<��[��ڱސ*�zz�=�;��k���iO{:P�����B��   �|  �TT@�) ���}5Z=�u�[R���^CWz�@$]��+֘w��U�T���3T�y����<ڻi2�ִ5��"��T�m^Mi����� h �  �5}��P����^���������j��h�ҞmҴ����7��K��n��
�h%V��    o�  ��R�0P@U*���AC��wc�U�QP��Ǫ�fJ7J��͢P����U'wq!.�V���%+�a�� �� �Fp�$e���P�U91�n��s�25R�9P]�S�EݸB�#v8��    O@hR�Q�     �E?�)T�       D���RaMBbM�F&	�@`�d�M1IJ44dd�h MS�I*B�i�	�A�b4��� 	Rl�I �b"y#jhz��O2|ϧ����v���|���zKđ�����O��<����HBHIp��	$$���$}@�BK�_��!I	&��/����?�~����~���>�?�����������D		!%�&��R�0$�������G�$�P�%���KC��@�b@`Ѐ��_�ąщ�H��#�BK�I%шKC@F]B]	tb�ЅѤ�шV0щтK������F�GF��� �Є�x4 IB		#� BLh� �B�I	F����AѡшAѤ�р�K�I%ѡ$%ѠI"� #�	.�!$�F���F  :4�F!.�B]$�4��4	thB�Ѕр.�:1 /�����>��GB\��OF��9�;�C`��S;mT@U�k>͠��k80���m��Nl˔���Ӝ�{,>����{p]^`"��M
��'>��{���R��Nù����rb`���j��@ne��5o-f�-�A����a��Ktuk��V���$vƬ{Qjݡ��i-�f�c�(-a	tb�ڗ�oH��uO&���Z7D[�f`��W��!���YS+M�+V`S��cf +&���m86���C��mf	����Q͂�kTd��9���#{t�u��+W5iĵ�f�M�*�O�����ʬl՗$:�t�aXU�+�)`�@�Y��M0�㦣�n]մ���v��1 �Ӣ�Rc��Ex㎷v�qɹs.R���b���(@���L^9���6R��{�kjռ�z(ɕT�,ǭR��i���j�aك7NYL���E��R�����K�H0)X�j���Wk`ܔ��2�4�U]8o��*�����Wf�d�U����jnM�-�z �E�.ڙy�X�+�Q�6Vx��W�e�̤�24�BC�he�����F�8e堅��Z��Tq�DR�T�U���ͻ���dYbf�j��t+F����;2�+q�^VҬ�Ԋ�]�V�1y��n��t�Zƀ��7R�(Ji�4�+���I��	��J�-TQ5���;���VPݣ��)Mؖ�Ǚ�a-U�T[1��$�K,^̧�$��4�V�V�Z�W��GN���fO������A�Y,�e�k.�F5�lKulS�I�v��*Wp�N������3P�F=���SA�5�`��A�c{u(���EZ�±S�t�Tj�`��N��4�1��U�mѶ��k,�̲����w{��w.9F�5d��+��T��+f�V��r���]fǭ��[8uʻ��Ơ��k����,��w+il�rm���c-ն�^��q����z�×���̫w*Y���G%nU����[��U�'�I�H����v![6i���1���#��%7��Ôh����Mv�44�&�D+i���vr��ƭ�ׄ�_Y�y6ؕ��ŀe!`�"��e���{[�rӣ�/#�j�+ז�F�����7GB'�NM�'&e��4-:�[@Ԃ�6�������w���1�������F���vb�BV��j�WwM���mԥ���#zb�����D@�ڔ�=�&��D�H�S���ڛ�b�ɖP�D����é 1@7�ͱ��р��Q�ڶ4*��wJ��Æ|L�+N�hlB��P��`�¶��\� ���,U�,dڃ��T@�wAO0mEci��Y"���;K��ə��:n��MX%��5@TG��:`9��b�J�r�:�!+I�֐b��u�B�/kte��AM�r���n��R�g"�M���m]m��dj"Lt��w��4�&�J��T�u4��^�NK�2�ٗQ������@q*Q�mL�[�,��3)^m�ɵo5j�I,�D^�i��V�aUwf#���2�Y�+oi\�H-d�u����yD
�(d��fN�����B��l�,ޭ7�,m,����!$U`��YܺҮ�Z��(ұMT�b0;x,�Wdi�˭�he��%[�[������� m��r;���n^�ׯA%)Sva]��uvԖ�J�ǌ���5x�ލ@�p��B��Tl��wf-�7��^l�F�$$�)�5�@�o����lf�f�t:g,[hB%���&�j���,�ca��Z��YWQ �2٭�;�B��N�ٵn�nir�̖j�tɴڼј^#�ѭfZR�Z�Bψ�6�����#w�,��7YWSZ;	����WV�ț+ᠿ�n��/�fA�S8ھ6�n���1JV�k���VR��-��O7	2M�`���G(ԺRa�*���f�����t���ĝ��^��{yNQݑ�x�]#��JRr�U����隯^J�����^�}t�!gN�j �D��v���mȨ�nQ�jhx�y1o�]-ͺU��:�h���a�'PV3Zun���[3,�O$؜ϴ��A�6*׹tܺQ*GN]��۫�f7XU��ڊ��V[�Ię �X��ei�xt�z@�j��$Q()Vlywr��3`X�%Ѵ��F},�f�p�Co-m��-@��J�LR�j�A-qQ ni�m�zء(h��!��]޵[x[����ٷ���pi5rJմ���kQO����ap+_f`� ����e�b�F���/EѸ-����X�f��I�*��hc��%ث)z��OQ#�¿���T{���-Ѣ/V}�e��Ov���J徖�%%m�Q.j��zMY�F n�a��F��V��W{�G��߭i�.�'�(太aXX�-7[nmK�&�%V�U�.��/5Y�r�ikicXM�d3f�;b#0�t��6��R6���{���5o�k̂�� F$�4p��f�nbJ�4�kȄK+ǈd�Ah`�*�x�K2�U�*��!�J|i�+*�S���63�M��E�͓Y2@�����q�;���wx�X��SO	P�T���m��4�E&�����h�.�9�fL��P�4��^ѱ���E�7m:��Q�U��o*�,[�/or���҂��siʅ��9�kt�L"�Jh�h���-�2�	���n�yg6h#F%J�jN�	��rJe�1F��jKq��Ul��L�7c��7jl��r�2YM�m��yq)(�T�ȹ1	ܦ�I�pb;��)W��,��,�^����D���t���O
՗h,�^7��,�EH�>κ��QX���هB��M��"�W�:�u��sU'bȼQͭ�O70A��H���NTSs/wK�����n-������0�*���Y����Jr���i8U�h#���i��2<��qջzV���q�WF�� �r�jQV��{O--4h!�u�G�sN���b�LB��Ǌ�#{�`�
����S�n�,�m��I���vr�4��e�5F��jd5b�9lL�	�2�tU���#�ڰI��B�������ץ�ٙ(��)�ۭ��J�om�6�ʒnG1���U{��H�xi�������ǆ��V�xNipQ[gܺ,�f��N�1J���b��`����#Z�U���j�X��:
��[Y��b��~�*��{�%J��Ub��y�n��@�-P�j;��޲.*V�w-L4[�ե��R�/Iϵ�-��%nK ��ݝ�욳�����ֶ,����x1KU���Z�1����G.����h��(�L͈��{Gv �۬�3c�1�Ww��ʒ�j��l#�i�E&�V��XFړ[�ksk�c�S���f/��wlO�̴���V.���Q֚�˅;ɲгAlrἠ����4ۜ��}Ƿ��B�)�g�n�h,y�mZ�v�9�/#�wJ*-8VX���ᙆ�ʍdz���� �a��^ıb�����1b��+�헇7��WF�`�Om�̽1ǵQU�ݙ[x�z~�ZЮ�]3eL��ثC�z� �H��VV�T��՚3j]驧*�i�0[@CI,�$�����eA������a�݅�S�x(�5��N�V�U��`,@����1W&m�lk���ۉجD�r�L����5�[�1T�[�u��]J�Ж-.;*+N����ۘ�$BUɊ���9D�*���'c�e��2j =�J;���JěVF�R��0�Z�ׇ�I�F4+/1�N�қs)ܰ^�%ʣwf�Kf�zinaV�!�p L�E�ѡ=/N`�ɗ�cB�2��V	�0�+T����Z�[��Dzv[xmʲeCcB����R�kE�޺8���7{w���uq��O/kV������̛�N��Y���W���r+J�;��Vؤ��J��#r:�^(�ѭ۱�V��[VVCA�G�Q�`���ٻL3`Ճ1��%�'F�W7V�M�DJZ�
1��^ܺ�+��dj�ۗ(¶�A�N�L@B������*-m4�PR�F�[e��]doXN����*�X�-f���ѥ�V����rX�n��	Jބ����u�Y��n��T+A(1��.��su]�t�5Cu��Ԟ�e\6�7K350���^ғw[m�B����e��/ �6��r�6M�dn����v��t�ز�U�*z2�d.�.�P�k[��'쬰�ٲV�;���k.��$��:.�觌'N�O�cQ�m��܊}����tB�����̄�nV��Dn�;��ێ�⛪�^��[��*EmSe����W3r�,��.�A�8�]��{�v�R�8�I��b�n7�d�õ�tR�[y��⡕6�j���,�M�/6�9N��6�R�kZ�*J��ܕj���f���`�wMIq���7j�����>��Ct�i:��Z�p�ՇVKնmnf�6��hlŏU*���BSX�ӗ���ہ*��έ�Y�r��n���stf9�ك����	�qР�R��BՆ�ڔ��.��P,���d�/0*h��\H�)��^U�$(��%�X�Vdah"�0*�GhXA��)����ɴ�6^�+M���&�B��n�#ͼ���B��Ou[d��p��P�j�=��Ҽ��W��n� #��
���^�v�2��l�T��L\oF��g�!Or�[���ol�/�ͫRe�dF�
Ŵˣ�K�:�bε�k�wt���=���nCmc�e��3ʗ)[�e�v�����mV"U� ٧��mf�H(�[{�9xof)�`%-Öj���*d
SQ���!d�ɤB'Pmk�[�xj�܋YC6ƽj�;��0nJ<T*�4�ح܄�2�&�3Ud�Ha旂�pY,�4�(ʖ�R�%n��g�4v��m��B�fX(c�n�Q�Vڼw9{BҬ�6�VU�E��4w����s�jP�149�s,-���SͩM��m]d�ИW� �#ot��v��SkR�{��0e�͈�YV����=y)�qb	d9����/^��C:��Ҩ.F�n�=j�^�,o6E%)Y��3�vX�u��{v��q����9#v�Ҥ���a����8�Ƙ/P;�636*�`��Tʫ��cU,M����NZ������ݣ�B�7uo��V�8����D��ҫ��َ�Xf�	��D��H���-�y�D�W�P7�oq���+�ݫ�kn�p������FJ�����fU�ݻ��F�s����b�Tu9��8�H�h�c�5y�J��o��^M����؍jĵ��̕���˥�r;qi�:J���ѓU������Ȧ�JF�*��ܳW�M!J]V8Z�WN��|*-�Y�0j:�X�N��t�(7^=�fKtڲ�$^������x�[.�:v���Ŏ&(��s4�u��,a&m��U�w�e��1c;�=����sYr=��iùR��ou5��C!�Ʒ���w+�^���a��)�=��\JH�����um
KF���@+4���Z�c^ֲ�h�a.��k�����iHh"�L0nMB����ۥbͩMfT�%�l]�"�u�(Jލ�uIDU�jbbY�4M2�Ѫ�b��V`4�����+E�.A�Ԡ��G��	Me�Rn+-�Nn0-7V�RV��4� 3qdˉ;M�I�X�6�fV5Z�X�f\W(c��ɕ�M��Qh�)������j�ޝ��T���o-�ی�$e�yvsm��'L���7HF�=��F���R����+ti�k;��Oܲ3/r���{�xd.�M��A��%�-<P�T���#�`��SN[�dҹ�����\�/Yb�X�*�@D���(Ty[��ݙ�u�dl��ԡRLߝ���I�:��d �^9n
��H��.�mnXӏݗq�:���*)�+jV[R�w�nݓYYL�+J���V���(�]�E�w�iZ��0�Z�P���Hݻdң�l!�!RSh�`ȴE�5�*�-�qˠo.��YY6A2��c[vN�Ѡ;����T�a�yX�ǋ.Á�aʛ�b����Y[�n+C94\ڑ�NҩYN�,U2��"�xm֜/.�-�yj�ג�YKf�_2�q��d .c�N8�+MG��v�E�vqd���&nޕ1��2,SUk���76FCq�i%�kPm�˻׹X��9v��v1�V�q	R<T,��B�;�-o2�r䵧p
�ZY�FB����:fkh��WY4f��ŵy��.�nMx��	��Or��#�hjܶ��՛��*ݓ���0+S���q�r�;#�{�*w����F��oTP�$��C\v�Xbѵu��w�7!Fb�s.n�u�eݛ�V��^�Q����B]��je�Wy�l�����*&�71�Ӱ�����ªbڭ��MhѡX���ki<�i75Y��]nV���+v�ɑ���ؠ��:m�c�M.�ȳpa�
�U2�m��F������J��%efջt-��:hsP�Vc�f�ʽ�ě�r�5 ʹF�X�-���&�R;�.ؼ���X�WmL m]d/Xej�� #��n�׊���ܬ�Qf;w�1a0���X�2AF�Y(=%l�,ڲ��6[u�L%[�/	��f:4Q�$��<�Ғ�N�#���$��X��uj���n��lxe'�Ve�T�6��;9{QS2�9cv�[cJY�V�� �ik��#��e��Y����p�Y��Kw��j���J������nزp�v��oFGy(((�7�n��IJ�5��
V�v�ܵ���a�&�v�O�+���/��0�@{�a�a^�bb�T�7Tj�e\j���Y�@B��I���R�b%�;,i��Sp��\*ƃ��жȬV���u�!Z�r��w���U��۔Nh.Ԇ�f�=�+/���<h:j�rjX�̲{Ul��	��U��G1Ջu�rݔ�a��"�]�K�
�Tݭ����E��qd�c�[�^Y�}y��������߿��xx^s&�/��C`�m$!� �h؄�m$�HI�$�I$���!���h@&�$�I!� HCi!�I^����9N�;�x T! lBBl�6�6�@��i���IM�$�$��HHM���ВmI	�H؄�6�` m l!���/ �(/w �-!lm� �&� �I�Cb�؀I �hC`�6��l@�h�$i	6m I�`�B@�؄�&Đ� ��HM�$�`�6���HBm$6�$�6��!$���$6!!��$6�	6`m BM� m!$&�hI�h��M� cI&�lHG������I[z�n�+��6� �Ё`�@��y����	�d+M]eY��3)���饻f�c4�H���wIӧw|����w$I-�{��_���Ą@�I��~��?�>������g�^}������=l��;�,�u?�����9�����d�����O�RӃ�j��mm$p�5J�m�(�U8�Z�۽���;+WL[�����e��<o+s�%N[��_3�#ոw-M����aw��A��n�̺�3sv�WcUʻ��X���ǹnf��� �}���K0����j��ٽe�E4��&��ë+e������C�c���Q�љs�&Z��{Z�����Y�i���m�>�O���Y��*MvL�}-�Na��gV^�EM��Ek#i��JE�Ց��w�Av*�2R:n�,wd�7;"��]�]nv��m�7c�xMܵ2�.�E���9J=wv+������=�ʈ�/#�!���o;W(������7#':�y����Q��jXz�n|.���a��}3/)	�%	>��Y����6	wj�
��kU��e�׼+��f7]ر����7���J�tc��ku�P��>��x�
�3��@���dʻ��՝tV���S{yXu��s���6wvѵyg�������kH��s��1tx^qk�R�����jƧ�a��[g��fv��at�
j�z�p�w��p���Q�K[��aQj�32�Y8*�"#8j��l�͘>�%e�A��pE�6�eի$���8z���h���jﶶ:���!V��h���[�`/4W:Xb|/NV]��C��{��,��K����o*���+���{�y���-|m���ZDٕ�6eK�uλ���زq=�K�l8�v�9 �y�7��[�wk��Ra�}"�mǧ��������Wb��Ac�fX[7��O-���/�W#M���׸�W�YO��l�+܈/�x���^�p���$z`�u���ԑ�*��v ��v�U�];��!Gt��M�k�;ߗ>�wt����b���F�y����HK	����v#���x��.��ՠ���I�U��'�7R�*w��ƶ�}�����é^J�3���`(��lr}]�ފ��d�Y�O�̼貞u��s&��dv�fa�ci�XON��-�\�� h����/6K[/p,̺`��RQd:��^S/.��*�����ˮy�s%�(��[�׶/��,�0�2]�N}X��%�z̼ 8d���ӧg*�nj޼����^Y
�n�ٴ{��2�i�:����
��Vh��2XG�:FR���6�^���|6ë-�gh�D��h����	ʎ�3�sB&�|(E\�ϯ��sf���|�ӷ	drǀ#��K���>�#����@ݛ�u��KCx�׸�;љ��'Y�Wz�i�ѻ�Y�N��_z��mӺ\f�ڏ.��f$+�.�r�v7��:��߬e�t��&�R,�����ͪ.���.�����ȨE��p��4@]���;��*̍k�\�U�`���`�K�9����W�N�U̔��Ww��q;�{:�ܙ�0ɽZ1aݽB�F(��R��{)�R������Ӷ�������:�Q�{�d����b���3��sU׫ٳjmjy�QI��'�������^��%�۸�[7�ɽݛlh�ʸ��i/���8e�:ʱc��e[��}Ʈ�l��y�ۢ�
ڰ��CY6)�>g�����:�o^�@C��v���	�9'��f�Q(n��|���f<�7��Ըu^nG���4v^/�9�oc�2��!˄�.Cx{������xuL6�o`�N�*����Q���C:�7��]h�W�2�^���kf��}��52��>�n�R���;��uv_o6/��ŧ���o
'�bL2�9�z�H��|�v�V�5k�Oh�7@,����J� |,���1އ�6�wp��Rw2]�H�%��奱H8�ї��z� �st��N����Y�롖��٭������7P�ZS��iθ����T�4�t�ݤ��|tVN`v�X�LT/q`:^e���5\3���b���q�X��c72�69����ۗ����:˸�a]�U�{��x�ŗ��y�q��f��P�����gq�Ax Ϥ���p}2�s�M��:��Æ,�G(��輂ZC�Ƹ��U(bB󞓹{zY!yy��d��-��JZ�e,Î�̥�q�̣��0���2�5<T�k�X�fI�!�%5�؃Zd�nT�XK������ydY��hYܱ�Q֑ܩ캱��Gg#�ic̮gL�UA�R�Q3q4đS$H44�������ȕ7&�SnV2�ψ�(����yYo�yRNkV�z4o,���^N�:�ә�X����:v�nȩ����b]p���i�]Vy;����3.�m��=�:1t��	�Ceu��/�Ȓ��r���Xru]m�@��R;�&�.�p�*�e.Nn^-3����]�k[�B`�Ϧ	2˴cxsy��1Ώ�9C؟Z��"����,�Gazt�r�p�7��W������'����r��F�����&�;]@��d����b���\7��E˭��t�K�.�9��]s��2��ֹRQ�嶵5]W��k��a@\�k,$�q�
�r`���c#����#�����D�fn-����jW�a�r���G�x�Z&a�x@��QΣ�Y��C}ֈͺ��[�3�����;�}�[׫o�Yy�b���rb����o�2�|�Q��V7e�}7��3�U���7�ݮ�poqӘo	�yV�I77��uuCvf�D��¸/&D��$�V�SDen��������ҵCAu�J����p��N�_v����e%�
�|��z��)�n<�m�4��z-�g�����h�*v��А����b������15R ʠ_n�{
�&M�Z�EWJ1���'�ݡ���[��K.rv{�D��m|�Y�-l�ս�4��/z�uX�W��#�v�N�����C1ft<��e�[�6޻a��8�vm�Qc�]��呐�
Gu�:��ܜM�����,�PV���qt�x���I[GB�{�Ԡ+:�񂊳��3K���]Q���]���F�
�w��y+wW��ʇz¾���`�ݦl�����9Zx�`r:oNWP+xm4�'�q;Suvm�x5��]�Gwv^_6�3��q�zk;6lZ��>5��e�X;8= �5�Z8�W%O2��u�,ۃ��*�˷sjN%Նi��(�eg �B�t:E��7 ����m�m)Zcύ���֤u�L�1h�B3{[��XXN��}�R�m;Q>��^CZ,�	�x�,d��rn�W2�w=1>΋n����6��i ��Ԯ���3di���ԥ���(XN�K�9v_G:�@Z�>5qT���2l-�n�=}��ed���1�q�\6��.y�B�X�L����a`3kn���Dr�1��q 2ٌ�c�<�v����ۻ��t�<*#�|u����Y�Vvz���:F�W��lS����7;���$YJn����-d����|�@����n�lswHd�;B��fY�&����E�k3xJ��Cp��vBb|��Kx�˗e�_s%<z�FZ�L�eh��o��z
�+������@��W&jw3-����c�������v�ݺθqR�<�E��>ܾ�Lh����J�3̔�Ѽ9��T��d�7��D�^官u%�v��шIϡ�kf�H-*�
�&��:�6m�LU�l��.�)o�u�[�(���$9�f��1]�&𱑷�����J�{���nn@���|荳������nZ�\����+2��k/����ۼ���z�R��v/�S������b�le��Ictͻ-㝦�W�f�[�34q��/�l;� R��j�&;�QfEX��㲳�3�3�����b6�����X�+~k[���IR�h
��:������9��P,�����[ފ-MS����0��Li{������,��
��c�T7���Ne��B�s�\�Pg/�jN=�.��[��m��3���6f��8��s�R�/^}��]Ӥ�ټ�d�l���&M��2�8>�]�8���:Ŋp��4:̓�+��E���Jy�>��Z�;e��eLBns;��ik3�d���\���r���(9��g/�jP�k2���` ��-e��[֨2�p��q0L�7:�0õq�m��(ea��z��e>��¥�Mn��D�cz�.n�)�X:rYZls�C��w�j�	�(;yIu˷��n�gl�L�X��{�}�̔+x���{��Z�E�3V� ن�I��ͣZK���u�v��фϰM�E���Whۣ��*Lܜ��P9����K;q�K�ܻ���.a�����QbF�o��iX�B�A%�F�}k�}���bX���Fb{h�Vc�Ó�t(^Ya�T�H�ɪ]��M>�R��]��s�+���J��WLs7�#�e�������r�en^�jT/]ڀ#tP줏�z,(j��V���;��T��p�_sj��+[0��G�du�h9��M����%jKYn�|��n�̽�8��D���{��WW�Q|��	{��;0����;zk:�sΥ��K�u��e�Ҝ��]`�6C�Ib� V�6��S6��c�-k�6�t��-2fŐ�(�8Q�3�Դ��S�Y���R��;�)�ժ�u��l]f��*#:$�	����NWk�ÛGC��f��Nex�U��N2�K�AS�����X+;��dïXS.���"1�'f�p|~���䓘	r Zݤ��Q��2����͸ �@:����e���f�Ux)4�����jm���{K6����Wu�L�ի���:�&1e�Y�WTc�S�8�Ѹ,I�3
��:�g���)ѱ�oT�,����o��ݫ��=�	�Q����t���Zӛ';�s����h�����E�V�^G��$S���� Z1mQ�t��w(;5�{��w��.�6a?q\��]�J�n����٧���W�ճ�:Tn��o-S�]OGs��s�Y������;;�a��"l�@��U�YՁ�V)�X��f�s����A��"��[ZE���g�����`5{�3W"H���]�wFP�s&
t���eB����4�c�wDu�e��)�Sxƽc(�lZ�v6p��.��:?b�wy�P��*��dåM��R��W*j���hޚh��ɑx��ćf���{�"�.��Wr^r�ݬ��Z�Ϟm���Ƃ)k��!ܹ���nv>͍k�06�_mo^6w�R"��p��"��p�5C{q,w���]-�r-�WdY��u���P]��V��'[��p����&�EU��ݍ��e�!9n�t��řq��%hC/�`�f�f��Gw\ag�1��6+u��<���'/��Ƕ���u�x��*LZ����eq���-!�v4��N�[�u����Dd�pp���|w;>b�S!��Ӝ�ˮ�ʥ���{uwC/���<�6�H� �{΃�����9�6f�Wr(E͸�O%Zᳺ�C�e0�td��ܯJ1b�ۺ�Jf�29٨����=jArP�{���X�q��Z�q؆�����뽛�����b'w<v�qy����qJ��.��	�+}��7�U7��*�������*[�\�Ғ��ɹ���w7���LݤV��Kо8�)v��]�v��"6��2�ɴZnԐb`Х7L��wv�w���SC�֥s�{�U1�
,���#;6fఞ��su�I�eXG��zZJ���	�ϋ�{�k/B��,��A�_ �T��`����\�z�gb��Y�t�ܡܫ���B�Wc7OR.J(�)�ŧ� Fk%7Ju���]]�eg�ov��ꝘZĭ�k��٫&��}��F�%۔�|/n�(Wka��ZCs�/h������l4T���Lַ��'r�;���:�1��w�|OI�������6�me3+YV��J��\�B�8��V����A��6Mr�`���Y�Dz-��.=���3*O:�疅7���$X��r���/*R�K;3Y��tF���9^]F4�Fq/��X���ҡ�볎φh��&uD��Vd`
�٣�p���5a�l���I]hj޸P$p�U�n\}y��4��0����՘�gqk[\ņG}�8>�h���XF���[��Ƶ����k�'f\�&��t��Bq<���CE+�����) ��{]}8��u�í����0�'������-*����� iQ[�� ݬ$;Vz�Mu<5���B��Sjf���5����~�d�cXj:4ە׈
Z��SJ�֌[���h���(�|���'��N	ʆ��b��1�<���u��a�J��PV��[�Y�:�AaK��OH��cU�[y�i��Q�h���nx���d֫5��%"�^oö��d4 �����ekW�L1VU�ص��n�+��M���Z_̬@X�m��N�nJ���C/�·X����Љs��N �o�z��4�MJł�-^��fKޗ�P��GQ�;8MB.�e�e�C�-0J�#�B���n���h�o,ˮ�\�V�={�b�:�۳�m���&J���<�"�+�&ūo:���t�q�eʒ'������*�,��[ϕvn˙o]أ��m�,���wY\��&$2�;��Y����^� L�8�кWεƥ�*�e�%�^.]���;�M�#�n�;�y�+D4?�nT���k�e��v�s�����F�R4+F�w�oI��c��il���9�'�M�L:ɕ`�HG*_Y�6R���J9����R��)X���YZ[��/8�C���ު�5i=Fdz�+/uc��^�}[��xrʺ��JU׹�';��|�N��Z	���8P&��LL���7�fj9���qNyC(u^�ޅ��"����G0�wQ��7��.�@�3���燜n���PJ9oY��\�pV�Wtu�`��7���kZ�R�	 ��X��{����7���ݥ�=��t�fJ���X2�*�zn��7_oj��3z��S;�Rz���m��pC�Aw�����y����&6E�`Y)̮B�f-�������X[���zyq�����m<�����>;���7v&Չ[c:�gY}kM;�����!	!%���>���}����� �}�����O�����p<�>e�&���IZ4��'k*�R܎�S���^ur��ܓ�W\�n/�~i��S�k�q��Lb�2Z\"K6�ì$cqnf����3d�F��Lr-��\�f�b�0�nwDx���<�/#��5v�G�R�#�"��8��2�}\!���6�e]��n�{)�/�]T�����^ta�����iXsֺ�MA�h�e�SU��O�<Z�q����R3m�`,P�9x�VN�y�K���8lں��"��d��1{F��Uɐ*ܼs�7:ȓc��hZ���f2���u%e���� ��%��X�3T;l,������#�ж����]��;E�\��X���w@�tz��B+g!'��;�DN�`@!��ջ��g���\�]tb�M�Y���I�8��6�T�͵�M^�D��,��c�3,�lfv�B=	�ksȸ�C�2�vbU���[5�k��Ylt�R��	�r�M\�;�)��n�:٧W��^����j�1�[G.a�w-�t�ɲ�Ek�F�捖�ȵ�1ef���ڻ0�&H�6e��٘��b�rq�����n0:v�3W�̶Ƶ����!rn��`�Y�u��^�����t����p|T��<y��r�l����)�O���3��q灇�L��`y�h'����M�C�{[9��q�S�z��u����`�=ی�	�v|k�+�bX:�YX6�9�aUҩ��uWp)��qj�>4�\���{�3��bL�"Pef ƨ㙚������	��s����+�Rp�*�m����6`{��:@K�/,�P�Y�V�����m�t�횛v��u��+�]��ۂMbl�.n����oq�8�\���zWZêR*��1�H�SJ2�m���-�{wg\��780s�pls�������m�u�]L=cVW���������n��#q� �u���C�9���&�ZͬC�.�,;S�e&-�юi5Zay��u���:\SP�ō]<�gn#�^{:'T�c���v͓�ns[�:�7@^��F1�\����E��p�S��Gb1�2V��rs��(VX�F��KJM+��������1����A�!�7F�{s�u�rT�d�	[u}�P{�W[�E�+�� ���u[M!
8��e����Bnn8��0/�\�ъ+Ao��]��RQ1�g���"Ĉ%]���M�pmt��a����X]�/Ohav�:V�l���(���h8�X0][[Us�}���5���\U�0 ���9�M<������J�^G��7�LbI�Ǥ�5q`��l�u�c���:a��	�h!&]��QښT�%���ĈwV{�y�<;g�eF�����֪��7�;��2C�[#�w��_j=s�iv��:����a��xb�6��!��;K�����*�j��d�q2j�z��y#�Z����>^q������.<�z��ܽf�wl!�Ma`Z�mvʭƮ�7���Ì�x9�n���T�瓧jU�� ����]`ۣa4�k� K����4�gG:�1�^î6�t��J��
D��yt�|g�V�ے�=�Ӹ5�b�������G�*��z���$Հc��f#4���h	//&��t���M��vcm�c��C���z�٥^�WK2mX���$b���Sj0�RR�켣�[6J�ӬG0k6�� 2�6��Urڸ�ʚjض�huU�!��=���rYbݸ�(�&yƭq�3i+��r��+��pC���.m��iRy,�m��u���K�x�|�ZX鉱�;;f9��m�At���N����6ŝ���L9��+5�kvv�1�4�ƕ�v�s{�7\lV���
4�=+������ō��0HwmÎ'zc&����')X޳Ƈ=�1�.z�� ��v�Ǣ��W5v�C�utv�cX����.6�Z�\�ҡ��0\pY۴����=i�Cv��mm��1��klb�6]���H�vr��Q�i���5������Bx�m���Gc�.��]�2��K�vsE���6���`�!,�G=n6�%��Yp6��� [0��بWI��H6Rm)�;��>7�.��U�Ј��I��g�����#\���[6��՚
U;r��L�I��Y�;؅�p����k�;��M2
��&R�n�0mf&ֻ�z�v�$\b(1��]6�n=7f5X��.��ѵ��֚�fZ�펀E��ㅸ.Ò��v�:���=�p�x��7[�D,su��ϵ;K٫�
lӑ�]z�p��'�^χ$�:o,Sp��iE����gֽ4�Ƶ���&��Z;\�n'��#%��q�5��8����8�ֹ�jv����z뇥��
y<���6�]����̵����n,�4��s��kN9�U� ��=z]��"���g%l�f���]Mb	eҎ��Z)fr�G�v��m�c���;S;�4]���J�,Ԟo;��|N�Ka֙v�-�6*n���J+â��v�Y�#v�Dӱn��,m��׮8e�[q�[��S8�eWH]pF{GQ݌�<�΅��v��GPuo/���ģB�N2�����v�ku�� ���7���e�{;Aڧl.�̹��l2ʷ�˕���7>oy��B]�C5"bݥ��\��P�;2�cj��CJR���=
���M�٪���i�{As�2�7$Y���$kh�r:b�:�tq���ᢇ��h9�i4J1�d5�˝{\=�B�Y㮧�;{ыc&jDܨkD0X�e�6�l47&�3p�,e��3���S�(LF�e�numЎ���CK��jU��8"�iF���h��kX��݃Q2�����/bh�v����%��6�}�j��}��n��z�s��$�[o1=v��+q]7<Ʈ�t�kΔe�������Wv��
�y��n�8x,F-^�=�;b�M�=�ff��hB���(�؆�@!@Xۺ��hf�q�:G���Ouͼ�:�IƝ=��UPr�wb %�wlx<�>�만�d\�+E箮�+��܎��'���h�۶얱At��ݷ'b8^�9�;m��e+���0.Zr]��W��Dv�����YCT�{O>E�m�u���G<mv��us�+�m%iGb �$帼�Վ������;L\��1�.70�LlN&<��H�Y�۹@Z�����y�cM�Nس9���tyH��f<V+q-Έ�w2R�'g¼p�pu�	�^�5e5�cl�/7�ȍ�h7m˱
�S����1��j�WJ΄g��]�	�m�R�ۆ�������Ca��s�L\������ܘ9؃�+�f��Ώ5�сa��U�u�cu{.�Eɥ�^�A�RݱΔ�U��L� -o=d.�;\��Y�a�{����EE�j
�l��T[4a�b���1�0.��dv�4jof�"��^r0dNɺR��ۮ֯f�G�����Y���1������熞9WeȽ^�^.t�\p#�]�ʰ{^n^1�/<�<#���x7O8�e�[u[V2��4=Y��Z��y�]���[v�^Be^<�<nYݜ7=���q���*����lk8��)���9�Q���۵<a8'qm��Y޺�r��\�^,\e6�)���2�m��x�KOL�2y��=�.;��NF�Đَp�9��*�շ���m=�����`��yM�p�-��"/S7m��������r�M���ci�0]n��b���s��\��'F\����Łfu��B&�]���QT�-q�,����
�,Wd��R_<���	�	������-�g��"ũ����ǉ��NQ:�b6��=`۰^Ɉ��է���9��⭎2��L��n3�\�mr:�ǒ&�V��n��rq�ny�N�s�Һ�<��vH {���+��;Lh2�F��D���|�|�Yl��� MEڶ��p
Z'��uňb�=��ݷO����V�ݮ��+Վ��e^aPb���гD>�`���s<v7mV.ۑB{�:�%v�mqn,�Xn֋��hႶz���m�Bk�������&;Y��ʓs��[�MJ����c��nT/C��9	�3m��H�k�\�D���g�b@��c$�����V,ѫH�쎖՚L�cn3y	v����h�e�K��0=cvĽ�����Fě4ѶlGF7h:fm)�#,�̜�V4�&�fNhf��uX�N9�*vڣ������1��lC6#��˗HaM�Ux�X:mczG��8�m�ALۅi��M�73�:nl7nۑ-]Fq�jܐ��M�k��QR���"��]��)�V��z��qr��CC�q��7=����g7�wV��*G��`ѵRm��H�-��8�{u�>,=<��\��z-���|즧>�G���K�Vl���'��KX��rm#-�dҳ@.�	y�\.���ƍ��kU���Qk^�
]uҬ1�	��Eܒ;n#�ヰζgU��.F�<�n��Ol����q��m"8皱����l�fk�kG/]��97���Д��lO�j䛞���GN{V^49��*��'��b轞`QIeə`i�����%�u��xy�ylWm]9����N��Lr��g*�]j�lڱ��qѭ������Įzp�z.-	�:��_>|�<cî�8{�u5m�%�s����r��5&�z�O\2�ղ7fz�Ut��8��^@�[�y	L1l�m�5��<�_]c�p�'c�e�vN�V��):M�oa�i+�����#c��@�k��[;8��z�@�v`RŎ�'\m������j+@QmF�9ݝ���<[��w)s����nu����=��n	��ʹt�vzz��G��	l��j�pD�n�n��FE�ch��S���5j���*�i��ӵ��ڎ���Xz�Y��r놦��Z�u��,-��1z�@�&}K��;�qv���2�E4�f�����ǞS&�*�ە�(��V�?���� �ʹ_4��Y�6����wؿ$%L�e\�?lc�g�>�'c� y�G��缋z��2�|�a���5(��s�����y��_��U��� ����a(��'����:Du�x߮3�F#����'�ɞ��ާ�g�oV�e}�\���/�1$�lt�ѕ�x�� �ȵ:�"��K,��ǽz�6,�%
�	u&�	TN��
KG�2����"��.��-�y�_~�d�O�=~�خ�6���kf圍d�Y�{��<�t���J���o~]d��z�uhu6�F��^��g�ɴ�Y^+�yY�iD�M(��Eh0���϶7.U� ��Ȕ��,�4�M�C�ͧ��@����4�".�rn$|��K��q��S�[x"yY�<��j�G۱h������uU�DB�H#��T6�{ϯ䇲\�C]�\�����Joϼy�Mf�a��Y�OQ��FL1��׆h�k
>�t�~������.��)�5�.�&��h�z�'�ڭ�.��]ţ\qm�uծ���sB�*P0�lś��A(ѥaa�Fh��Zg/eiQ�d�F��1��ݩ�w8N�
u�^u&���`�i�B*��:�X�,�K4!1B����{����-�6ż�$+��m�;X��
j�vmb�aX��1WMFv.Y�-ձ�7C-��m�q*ٻI�]���W@�3+̹�X�2�]Nڰ�K�\7E�e8܊��zk����s�<��̽�iC��ѝQ�*��3!�;���.�Y���h3c`�j[�WM7F)��]�,l�rU̠fvwj���lx�ȃUƻME���jj��4�+��s��7ux���Fi��,�&�9]���Y�^dŎ|sm����:v3fP��t]�q�ޔ1R��n���f��]q׋\Vu6N��^�wÉ����2�귶�@;ی�.�o�ã&x�ҁ�e��Sc&�����d�v�s[����m(�.3Q���y.+��QIlK%asE� 6��2�lM�C8��s3�h�l^��r��&�K-tL٫.h��2�R�XE�[K΅%r�ꑬ���茼[�kG�[�u��ይ�&m���6����H�Yvi6k�����,�.)V0���Cgf8��q�W!���r��x�g�e��M�[�7cW������8�Y��Y��lc>`-W��x�M��e��Q��U3��i%�E�W�Q�����,Z��F����zS]h\imڍ��N�uB�ORl�-pT9�G�R0�lfqf�e��g����Sӽ��X��չͬI��mʣ-��0y{L.���SGK�f��欏\,{Z�7m-��Vc	[ۺ���1�xQg�r�]��ٜI�^p�I1���CJ84*�*i�S\�1�����o;8�psP��6ds&�{$N<y�z)��Q5�$��/�b;i]i�4�fl�r���I4�u� ����bF�R� u%Z��^֩�Zc
�ʻ���ŕ��LxM�I���9�L��Ef�.��v��X���q7L��E��\�Lg�m�v�m�3�h�d�DӚ��&ժgi��
��/l�Ƨj�'kjq��,b�"!Q��l���`���>�0>/"����tI����e���%��4�+����5]����5[�T����7�4�X�Q=Wm��ɼ��f��H�2G��3�PI���3+9z�8�p<9�.7�,*�I�v;��mF��{?r�?H~�#Uk�wh1$�*'m`��!B��x��z���ԑ��=�B�ߺ�nT�7����d�c6��Ȫ9�g
��rY���2�?II��
��Įa��v�r�ڗ���!�H��/���|�ҧ_S��[F�a�n�@v!��<旞�1p��R��
�6E]�v-Y�>��CU$UOW�;8/tf<HP��K쇄�b�K:T�&=��l5R���):�yR#���$=v{R����7x*��`�ǣlc��7�\ޮ�B��L�,ͷ��Wm�ZN%�֒wl�e(rWz��f��ۋҶ�}�yz�G'X{S�NE�G��3x�ڭ�$U!��m�T�l�?<�<Ӫ�vwX�'T�U^���]fŨ���W-�����q���z{��"D%�<0� �N"�w6XMwn.�HjH���+�+�Е�&��ײ9=a�O9�$��I7�<}oD��Wa!�K��`.��JZ��IP� ��F��\�8��ũɈ��$�7�L?}骤5R0���y;=�-	�/�Xɝ�o�n�}�z��5R"��f]`����Ǫ�k��^>`�0c���B��<7�'vV�R�@ ���}!�$�&{�Gt�GYr�T�͚��&��+�1rP��"��,�N���ŝY����J�#.�ۣ�6���c���aEb��"&*���F�f}<Tܽ�����UHd5$U%�Og���
#.��r��U!��5��ד��vQ�R�Ux~�<l!2߯�6=W�O���H�2a����%�~w�����}�_xu�ʹ�=��lR�"�웬�ǔ��ZآD9H*�(Z�EѰ�f�k�]=�"pq���wVƅ�R�A�H�F��ک���/�4:��Խ�#��j6��z�|�^�j}R��H��꧷��9��}�5^�䣿W/^N�u�FmK���I%�mP�[L��Y??K5QꪒK�!�E��f��Mз}���U����Bj�����p�!�*rɽ�N����V�z9���۾W�Hg�=��-Wq}���h �t��ϰ�uw�Cާ�8�B���1,�*�^V �3���fI�^y�Y��]s�` �i��o����5V�����,�]=U���2ER{M[6�N��]�c�˲y{��=�/�^IuRERW�ܫx+�KY��HPE_���j�;��8{at���];�S��C;,���[�I�~��<F&��wzr�mf��ء�B�Պ�!6�7}�v��w.��$�y4�U]�}��y��a��}$URI�SܯefߝjJ��˒I�X�_X�㹷�<��:����~�?HjH�C!���=w�"3̈́��U�5��RE^<������鐵'^cB��N��A�G�U�d���!�%?ea�tn�~��{���A=a��}REN��n��E�0��~�J����we'��]�$��Uu�m]�&b=tx*}ui�7�<�_:+��q� �Kj^g�����2�N?qui¯/�����F��*��h�Ŏ�a�N�\���I7f]6��h�iH�c,�U�`6�E٬��KgE;��(�)� ڇrY;H�ó�2�s�u�u�����c/�۴v�%���c0Va�LDbv�χnn�pj%�k�v�ò���	�g0�n.5�Ȝ�����l��-�=&m��5b.2(F��-����͎Gk���[�����S}��t�u���l�\hq�*u�^˵ڒ�ىx�������|�ߒlO^�3ף��GĦ_��~����ڗ�{ᾐ�ꦲ��BN$�$��U�A�#r�C�k\&�[�/#\�&���`&�
��[wB�����]��?T�H���I�d*���b��"u�جF&�Е*�H~�)�;��KrW׸��jC�L�0���.�6zT�}��"���qK��n/��d?I��u���:8f���l�Է�˶T���m�7n.��u��>_W-���?~{H���*�������8`ǃHS��,��Q�g;ucRa]]������~��צ�C\p�n��	�+�M�Z�<��u�{6��O\�Hd4v[���:Hh�eu�7��bJ$�8gJ���K\��RJB����;,Cbl3�/,��㝉k6�[�k�ܥrTlI�'W����~���5�(��>�<{4��R�W��$���Y�9;��*����yUHjC�����9l��F7���^�=;��
���6�v��5$N<�W���U&�3���	�8MV�o�uٗ��ظd4�U!���II�q�[��K�{�4�)�ڋ������:���xj��`�&م���KG����rv�ڶi@��Bm�F0l������og���l�U�7b՛�T�WӍHd���z���'�i<�լez��3k��E� �x�ӏ�92�4抎���#��\��<Y���x'�𚭺�MjC��ޣ7����4����E!�6xh�����J�}��L�d:��z=5��)s~��Y^oZ�=��U2��g�Ó\E�z��72���V�g	\�FV�[0�d��i��J��S3����;8��+��I2���!���Ç�����]ۄϔ_s=7����V�﫣��3wŬ�>��$��C$o�^Ƌ�	}�s����'�𚭺�n�!��RG1w�"��&�]��R�+�Z�m�ܧ0�]�؅K[0ͅ���ue$�hn_}S�5UH~��Q�5o/��ψ�u�����Isަ���_I%�$U���޼��`��U��Zo�^��^�i�
��*��s�j��l��6�R�1�v�v�$�B潛�u��&��bMAj֤2�H�CY� �"Fuz�޺�?/���C����V�w�9�ι{�?U�o����b.pٻyz|�@y�!G&����r���d�_�1q���wb�p�=�yv^�oIÙ�R�^mZӄ�-V��^�~ǋ�|jC��W���Ul�̢��8��5��a�L3��P}]��ؤ�3K�ֽOl�!D� @�t����.��X�r=nW��sg�uc���t���3nX��u%^I��vܵY2onƤ�UZ��z�)�/����H�C�/gY}hϫ���<����<��ψ���(a?Hd��Gu~��kު�~�4��Rv�IY��n�;pb�^�Xe����Wi��q}!��I��k,B�rr�CU�.ٯف�J��x�}SqU�ǽ�t��le�@_�~�j�C��$�<L�͍�:gy��g���{��ψ}8/U��I&} ��Th�C^�*��f�1��5���c=dd������1t=Ql��õ�ހ]�{u�x�<�XP�n>�ْ��o���/��%R;.����N�0A�v��sqՙ.f�7De,��hD�V�v֚�Z}l��=rf�3zG�Mv�8�=������ !��lf�U����Er�f*M�aQ��K.�L�.}�\wiP�Gf�ul���jY�nqvƦc��c���׬�h�h��Oc�ѩte̽���c��Ύ��?�D��aH����*:Y[M�e����pSC+a��d���7�;��aI��śu���6�\toQ��X�I+\���Z�VQ<U�*��R�%x�=}���������O,:�n���wswe ����?�a�_R��'nlm����R��o]�O1��/M��P�0[_.?UI$�+��G��쬔�y�tӋ{�>">��^�5RI(ВzP�r�seI~>WƤ?I��.{�����Ptxfk��3��x}J�z�n��޸j�5$�/,�䜙/�:0�����}2WM9���S�UR��M\p����|�i���}`#Ifx4�Z4Ú��t�*hl�d�ꮕ�$
���V�������)�>�r��^��">⧤m����w��g���m�y��i��N�BN��J�jd;M��G<mk�ڵee7&�b$gf���p��γ��5stn_+ �7�pض;���OJ��f�z�_l�[�hyz�T���*��'��%+�K<j��O��E��oGV{�@��s�J�71���q}�C��}!�ȣ��Y����{%'�!��ݎS������G�R�5�Ulu{a}�*[�=͹�k�p�I��H��86��c�=^�-�L,ݨ���VtM�n.�]��>��_�g:�i�'hcrV��8IL�zAu�{����a�v���|��]�K�E������-���S�H�v�mԥF�m͍�h-oUO$Ț��01�]�?=5RE!�CC Ol��n�{��{�J{�{�w8�������2M���w������4��OzL�C����WR��mJ_vT�����q~Gl��=W1˲OҚ
��47��z��G�g��+w�\0��&�\���r�-�:��2NVٙ
Jg�CnL5��,g`�N�Q�xgI�!�����[���B�2�^Qˮ5�D�K��ՙKWwō�Q�Ӓַx�g�ǐN��6fO�E���ws��	�ۃ���4N1�/9���}ۘ{�%f�U˷��D�uKp�.��b���n�j�b,[�3���X�wa�J�H����M��|/y�)��	J�r/��Ӌv^��vq9;Cj�MƖ'|($Y��Y*�c�,I/��B��h���̬�R���*t:�����8�.'�]�̉XtoW�t���Ϭ5�InU��Yf�(eu�M��Y|i�J�Y9���ieuL��]D�D���H�������Z"��`��X�q�2�`m<�ULӒ]!p>�Y�x�V�Z�.��4�:ݚJ�R�ǡ�7���d�W�*����2��oh�C�qv�Ts���a`���Ս+ű��㵗W��r=�;m�S+oq�#�����l���T���Z����μr�������T����*��<\��z�g
�]mp�]���ʷ�NX�u�i�Z���ڽ�k�=�M,�O^�s���[u������O:ﳡ��{Z�Pɪ��[���6�"��j�&(s%لJ]|l�#3�j�b�2�n�U�B��gk�+&`^��B���]:��z�R�yg23ХghXc�ՁV,ڦ�y�r����ޞ���d'�9u��DoF�,���J��;��۩�48p����}*�@�,{���_��G߿��D#�y���͈ʙ�nR��+<���_������d�_�A_^ԋ��+�vw:'���x�ry��/O��/I����1�R�F����C"����&Lǋ��X2/��*���E`��A��ɮ�k��xg�Υ�b�c<#g����>��Ϝ�/w���"x��EZ�蟘~��ߓ�蕨��Ϙ��6��W/$����G�Գ���|��׵��EP��Wd�E�S�O���無��w���%E�I��a<��v�z��Jc��DfN��&T�Z'��ɑ]���<�ﱄ��ȑt )�8IQB�I���=fx�;�%�+���ˢL��,3t�|�>��"�! �����Y*������
�i�V���� FYFX3%��II\�*�f��Ck�֓���v+��TEeQ��ܷT��|�b�.�쬙�$G��=���5uW<���'dEM$�u�7Q���<���f���LOJR�<�(������{M�U�"�\�\H,�|�ǀ��F/s*�0Ո�	��4�� 1��h4�e�D���PiY��Q��Tr���Z��F�������FGCu��7
k�7�*� "�K̗O�����w�F1�L̨�eJ�(Y<�#|�9fx�;��މط��S�,����AI�ITx������u�oٛ��f�!�f�K0a�R��%f��n�+�5�֘�`��|�{��~y��\�pRg� ���θe��ul�e����Wc*���;d��f ^l{��Rp�$�@%&F0�2�`6���x���#�,8�{+#'�����5��u���1�x�L�-���� �Gk8 �����$ ����կ/�C*-�1��K,�l�G��9 �� AJ��$�$�C%�6ktX4ƾ;�8��{�ϒOl�{e��1���p�nwX�;���u�ɚg�"Ri��.I�
]-IG_on�M���p�Pv�ݽ��3բ��+`�#�Țx4Τ{u���W2Ȧ=x����ǞM����\<f8��A���z)1�fB!��#�{�+x��=��f�qCzq�5�kl�=Δ��	�g ���v�A���xM�dӀljf�pCu��2%�ۮƫ�8�^z�^su�k��$�sn�
G8��2[��r��H~ڻ��{n�e8��;�1�2���B�	�kk��f��Äû&=��s��pROl����s�{��7��uk�}{e���[��Bf�9��쾁 ��ە�gM*c�a8(U8pD����
NI�I?�U����k-���V��Y7	���I��&pA)'�M�#(�v�oe�� �\+X9'��vw%�����,�mG�0pF>�٬Ny:}U���9I��$�A�O�&�xi�^+��wD��dc�nw��l���	��p ���$!'��ov{�gY�]��ԉ����\���~Y���j��wt�oz�eit�t�W��˟<�s5��'��o�čem���?��5},��6^y����n�pf�p�D��&���ڌd\�e��&��c��^ �=M�q;�M���� ��o`!s����$���vb޸��
F�-�K��1�K��O�7V����E��|u�u#�6!k�q��v�B���lt"-�����(yD{f7vy��CV���=X�J5P�ڋ�$�F q�\B9� ִ9z�t����Yt�~�҅�>T��5��u٣�)�+m��	�x�i�u��s6���˚���r˾3헯��OI�!%�>��N�x�\�U\ɸ���aA�[Mf�nq��'_�o���	3�AI�!������3r�o;�U�6ɶ��S���ڇ�`�Ǚ��^�=�]}[���"�+��A:��	?���RO�4B��\��ف�1Ј�ţ�n�pAԠG�L�pU���O]A�a$�^W���$�}�ֲx�_]�ê�d�A��I��"w�|�L�ֹ��$�pR`��z�Z��׳Ca�8~���}�؞c �w����M0pA'BJ �����N<�d"��*�д� 5�Ŏ�"Y�8m��X79pL��E�a�uڥ�e���'��m?�q��&pC�$����fwՊ!���f�7c_�����V��$�$�@ ����׍�X�����c����H)�8NvƳd����c,д��e�z��u�������;P�2e��*+ce<VQiBm�Ze�� u��#u� n?�쵬�-��V�ʫ�7�@ ��p
M2;-�t�f���<'�I�)0pA	8|9q��6�~�����f'x�9����D�!J�)?��&rw"���Oƅ�n�?�;��@>I<c��;���bxg�����s8#Td����Y���։<��p�$���9'	,��Q`����2o�l�nN���xeƯ�f��
O�&p ���Cu���~��V���qcم0Jil�	n��Z���ˑ�K��u�6J���t+����ܲ��	b�
L���}�P��rv����ێ��k<Su�0/]B<BO�&��l�w���ƙ!��z��z��s��9�Ý[�;T���'1����G�a���:u�)��na~"o @"s$�Ȥ�����w�?�/eC�4���E��J�㣃���܉7fYC��gt��nV˼����+�kwe�� VwiN����\���]�k������jΝm~WV"ֶ7��O�	?��8 ���	7�Q�������|A������'��v�`����3���#�L ���lRi�80�����ۭ �s1����r�M�=�>)1σ|$��x7egwW�8�c7��A��I��Rp�~W��ylv��砫�u�٤l�Y���0���q=1��9�:��F
�T��5�]+7f���#rffiG�O��=/k:�ەՈ�����UU�ܾ��;�ߞN����Q�y�4�2�)0ru�i��/����4h@��8wݫ���'h�9����� ��?����۾MZ��('˨1��2hc3"�&p|�scOM��\������#�����A��
LRp�!%������o�0�-����#�Z?Y�{Y��ܮ�D%\��|��u�K�	D�&U�ml;��[��l�_A!�`0��5r�s�'\�<Kx�O�VҠ�
�sM1�Xԗ;h�sk�ђZr���8����f4�1��fc��)0�~����^
{���;��݇k���2gz�8@&i�I�I!!'���;�����c �ghghqL/Ok��G���6�B�82v�5�)h��{ﺫLc�{4f{y�4�2h��ں���v��ы�3p"��`�M;����� @;���9	(�JL�>��2Ρ1���>"+ G�������]X�J����U?�`h[�Eh�Q.��;H�y� 1���O2�k2Ǵ][�f=\;_+��3;أ�6��>IÐ���	?��9�@[$E\^��֐|�x�x����J2�3�3q ��`��Ê���sQx�4��r�p�$���L��9	#}���˂�����8r]-��n�V!��ln �T�!'����A$�Ǟ�7���yP��|s3u�1�=���;Z(^��G�[�N�:��u�lum��;�:K��A����o��[�s�c'9��7g�E���+?J	,g�:�Zj��%q˸���w�I�=ղIԼc���[t����v�ݐ�#�\��p��ت�u���]Úq$q�W�۔�f �b!)-�Ema������Ln㗶L��F�@K��9�1s�,:4ã��m0���H1��vmc��f�-�XK�=Vn!-���Kp�$��I��b^��WX4h�z�5�ny�ҳ.�`e�g#1����?O��X���҆ku���g���cVoVn�܊�(�]-f��o�������G���#�0�
N��õ�#3��8@Q�e�j�Y�$�8pEj�!'��A)'�"i���,9�c9�$��s^>�s;R��Ɍ��}���ۙ
L7vw2�[&�c���*Tz8�	8pBJ#�7�b%,hwm��毩;mJ��kcp �T��
O�)3�AI<x���"�0˵�V���ft��`$�����d;_+��w��f�9s|����4n�U�#�S��I ��ǈ>	?�d�6#��{�E�j���ׁO6�Ͻ����)�c8c7e0����jUB�w*مl���%T"�*�nL���;���D�fmR7"��]n��qG>��Fn�>9���Ð�$��և����b�d�[�F�^�3Q���A�8;���RO䚈>)0��<�l�4�'�ԿN	N�]�]�҂��ދS��b:)�{�Ta�X�{��f,n���6����N���{,�]�:�B�k�e��J,\	#+�����|����}|�䘼�^?z3lx���!��U�'ޛ13��}?�5c@ �T�BLM AI?��T�a�/M�ii��ݩ��5�9U�Ɵ7D�w�42���DbI��z�����x���ݱ!'�i{[����:b��cw�>7T�A�-���{Qo�ɤ�ʌo2�Ǚ�4�e�$l���[�W8���sC^�"�&�;؟��`�$�$�<BO�m����O|}��XɢUV��zkTBBh}����:os�9K�������ڥ�#L�>��e�����������׍kl��wze��0�c7"ҽv+[��� A����	0p��JDy& ��t	�O�-�<}��|���l��r�S͍�L�<Rpj�8�0��0�[�g3�A�=�BJ�?�!'u�0�|�z�t�L_�n�E���Sm��rJ'��w~O����1�9��}ru
�5"]�`xQ�PD�2����O3�#t.^g%��7!��Tk~=�㑔�u�^jM�-S�{� ��!'BJ#�'&�C?"�������>R�M�9�	���~kl��wze��0�c7��F�,��]esd�{�Pv���̆�e
,�A��Z�C�/Kc݇|�[��Eʍ��-�!S͍� ��x��
L�>I>�L���f
V�?�:܏ۏ��ݘ�y�gc^۶4�ԗm��Y��F�ʚ�N����z� ƹ�ѡ�Q<A	8n����n{�l�j��b~��,Ì��;`��Ñ�G��'����A)'�2e�<:��#<��<Oo<sƵ�n�s�2�j�\1�� �0dK�	1��s��:���������PE�����x���0O��׺f�sȶD4�mV�7A���AI�I��I<oJ���]s��gg&a$�����Rp�Ӷ����rM�MS��OޏU��a����~'�w�R{{��l���^�#þ���Q�nk�]��qdWO�Zi��gJ�sP!&��ic/p�{�x_��ZL�b�̨1�̆�fdPy��(�2g�f�d�pV��=�՚s�ie��0�c7 A9L����W�)893�=?�X�<���|�_D��:��Z.���3)�i�p[��dtx��M-a��W�??=M,�����ÂO�	?�V񝌜�/�bQ�U͍�PQ>3�E����:������	0	0�~��p7��/�8}���Ƿ�卑qQ��O�5l��8$���	�o�sܾuq]���Loy�@��Q<ʇ�'�y�k�':��o;J�ie��0�eW�|�1��ѧ�DLy����6q��u�;0��\9&�b<�
<8�d�o�Wl�y���n���̙�0�m��R� ���&�|� �(I�cި=360_8��{�{y�X��s$={� 1���ffiifR�~Y�A
,��j�yn�����1M!���Y��X��5�r����a��5ݛ�����	���^���1�`���k$�(U�:+Xw���>;K/���-���B+@e�,h<�l�X'��T��&���-V�k���w5z�[B�V��j��Uз2�&��w=Qe�>�Evc��i�������E�vO�r���].���W�F%48�Yu��ˌ�g���(��-h�˳��]G�0�>л��m��R��.ͺ��gx��W�w�78��n�ff咭��﯅���J��M�Y���]���j���W��E9Fb�Zv�k{@y�J�XV��p�x�F�U���	XP�|k��C�ﻭ�u0����w�Ngs=�]�����.Rwu���
�Ӈ��ɂ�.��m,\6��w����ޫm]��f�>�},�o;b��{�����M,�-�ǝDX���_&�RZ���E�۪O�!JӼݱ1����-G�����y�tᓞ�R;r���S1��]�֫(���5�pp��;j��˂��������VD��Q�B�˔�+.�L*�N�wa��ܛ�U`�8;n����LJ��7�g��{ �Vl:�CC�WT/��:/b�w�s��Ewqݱ�*)��&��x��Ȼk�Ҋ��2&/�2�1J�sS	:� J�[xhm��Qɑ���⦲�[Ga��;y��0+'S�O�g�%gʳf�����(!1е��>�`�fQA���{��c�k��)�U�� ��P�n�
ۭڗ#Ʊ�s2����nWm2�i�;�.��3n�<�S����Ϣ��S���������U�G�V��No�L��-!�3����vT��P�%��$%g�y[��ƺ�B@z)%��TS2�2�Og��9˥�E_��u=Q�y�$%I�!�Y�&r״dT~ע��{&����I��V�J�+��P�%d%�rZ��"R�����{�y���w/}뼗�n��3��;�ؕ���WH�	�c/Kv�G]vN�T�\Ƚ��|����P�GSʫ���w�a��bUx��l��o(�����(��=h`&rI�'���eW�*,}H;�4gt<�3��ۼ��[U+z훑�'�A-Y�<��&�|��z�TE��A�Ⱥ�He��%"�嚡����n���Ȳ��4]S4�t"z�ɜ�\�B��{�\�����}l��p�=��:�Mʉ��{Ǳ5����OO�GUm�Ȫ���-�7WF������"#OL��;Tt<�JE<�����l��5t?�i若u2W2�m��Bx�o>�f�\���\��'"��ʞ��;Z�&�ki3E(�3����u��wӾ�4�\��@�I۫�����:���<C�J$�lx;�W]�^ݨ���lcmo�&�բ��N��(ٴ�ͰL�Mp<Sd������l���k��t�-\mha��A#�a�^֨r�i�T`�8�pX��.�P�m�!p�*s	��4`�c̣�N�9�F.�x�{v���M���^3Z���4�*����6���'d䬅�N��I��[��x��K�ڊ{I�nt콍k�9v����כh:.5�̈�F�rpxw<�t@�t�72�8E�e�4W\Y�.N�c��3a��"Ҳ�-�����;�!M�n�c԰�m��xۇw\D��v.ԕ��M23Y��PNp�%�����o/{�c�Yb7+�3>��z���6ݥ0��Y���C$,�<y�@�>�7�m�޷*�S���+5Uly,"Y^��]���8h׆��SR[�Ԥ�X�����gY���@:gjf�H�-&v�sID#Ak�s7/SW���{Gf��R1��WBP��R�lXS�O\\�+�gU0�W;ucojaT<�}kz��(��Ǟ�����E�,#�#KeCi�=��%ೈ�h�gr��E� ��(Z�YxC�'1Jv������/�d�:�3"�X��3L�A�ИY2�mI�8��r�ت������6fhG�лMb�p0�[۷]u�,���N�S�w[���9�b�H���_>��.���9�Y�٨�q6v�]i�t]��1xz7b݁�4WnUݬ6�WE�F�ѻ��úժ4qr�S�ܤ\8���������X5f��Қ	hZ�1[�iv@��v,��>%'3�)��s�n6I��:�E�<X�]����s�����6�}�Ő�{fI����y�A�t�mr+َ�	�4ui
��/Zh���F�o�;��n�ۊ!:�M�m+R\��6GeniaL�8Ǝ��8�9��7ۭ�^�b�A7��=v��գ�B�Ž�:n��kM��^��t�O&/������W]P�ŋ�������Lʖk[1b�J�!��ݞ;uۆ(�A��az�ɳ�T������.��Þ�4�֜��0�����]���g����6��qd�6f3�tR5������P�([��m��,�.Iul�:�1�D�v���n�l�cm�l�v�T.���fy溊����tmv����W���=��;[��]�kc1���}߇տ̈́��MW\O[7H/N\�v��nl������[J˰ms�����?�Aj�е�I��$�2#�����ye��0�c7 P-[U�`�oN�0�A*=�¼BL�$�@%&2g1�:��n�/uq������gk^L��~v͓͍��t�#׎L��[d�޼)�f�r	(R``��V�]%L�x���|�O�����@&���f@�ȷ�y�UN]V��7��pc�\�����{�����1�ah8�>9L���HȺyg��Z��0ILD����IE&�N����}e݃��ƭ���~v͓͍��n���㉃�� �ucg��cƐ����8���l�:�=���4�gQ�fn%��u��kc08 �0�Dz� A���1�+[-��>>[ӭ�'���)��;6x��9j#Ĥ��2fp ������b�e����*���MP]����d�6�wM-R��Kz�����*���wXpS�".�Lօ.����IXb��h��< �K��3�A���x�&�t}�fc\��cp�S �̀k��}
��Ç7�����ȴ�$�G��L*��X�L]�6�*���~V�'��A������9�����v+��G-�È٧GcY��s�-��;f[S��'� 
�pEa���nx�����#�b<A�`������y&,�^�M��/�9����fc\��c7���F渀BL��Wim� L!�0�������{g��\Z1۞���,��J�]0\��F�e�������������	(�
L�������/V�'��wlr3�y�Cu��������p��Lwu��%ۺ��!��c�螻�o�|�+Yw�?hc7u�̄���w��Mq0s��+�����1��"eF1�d�\9�u>��_C�Kt���	|+/f*�Y�
����v�ܮ}���h�v�"p���� ��������%a�e�̪$F*�fU�����L�U�7C�,Ms�|���;�C3*1�@�͚ �i�n���h�a��0�yS�I�h�P�������cw��������P���������p���F�(�z4;6c,�]��S�� )p���^�澻�98�W{��L�.BLJ�x���S���,����Cԙ\f�XۯY����(��ꎕ�V۞��Ak6-s�e�V:�>���Yz�������&��I���7Gpy���apE��I۔�����C�g��h�7PrN ���Mu{;��"%Ѿ#n��̈́?�J���xg��c�͍��um�!�Ria��d�dX�o L�,�� �i�x���Rp�F]vU���=JYt-���L-�c�zM���!%�"��d^B�'~�xix/ֱ�����+��%$�ϡ�7Ghi�yo.�Yn��@�~l�a�_��b����R�FQ�B$=SGS���7b8��%%i]&�M��ه/��$ɝ��i߄\��e�R���f�O,�nXnє�� =�����}���IG��0
L �s�ѭR��4u������q�W�ggc���j�����	���b?�L�>I>Du��V�x� �����
TUj�4�@�.��nԎ8L��ݹ"`�&�+c�*[����lg�>�e�1����
I��O]�k6��������ft��d�;��������O�)3�AI<[>��ݒD��3�	��5�C^n��i�W�,�Yn	�`� ��
(���͎Y���Es�N� ���I?�&DEN���v����&rVlC�M�9��A�#��L���	7��^iM��p �A�NlMm�kk������n?@ �0r9�k��x��%�a��^?����pRO$�$�&#3g:I~�J�x��Pl�Ѽ�1
�\7|v�?�ۙI�
Nh{�؎��0"�$�?D�� ��z�q��k-����擳g�w����n��8dv�h�&W�7�e7�Ρ����+Eх���[N���'N��ܾ���5�,�܂ݰ�%�
��U��o'f:��8,/h����Y�;j\ס��րCW4\�=˻�������S�0�:x���m�ؑ�۹�u��t�k���m�1S�X����v�5��p�s$�G[�=[Z���1۝&��/��Z7P�;G�����ä�>z�v��ݮd��i�������d@cOdv�]��f6��Ͽ>K���.!5�M"S��k�j�:�i��N;�WFZl5�Թ*;g/�=~3�SN��G�I����\��t4<M�9<���.��-*�:�o��:dC��@)'�G�0���B�q׊ p~��E�u��Mu�kj���9���w���Lfd"ff*���rx2�-V��)A��4ǌ��*1����ߛ.mY=w����31
�\b8���#s AE��8�����3H��q�H�p��܏G�dE,ѕ:���&윭lop7t�ֈ4);i�ݳ�M^ �����0 �?�I8�QM�ͽqN�!�
�^]�Y�|��+���84\Rp�$�Й��!��1�S���P�a�a��#���٬�l&���s����p�����`�'�G�r�8>I<c�1����b!a�u���b��G=*T� =�
8\����qE|1ߞ�u����v���Bk� �y��8��5��sr`��k�*R��w��Z�4��d.MW�9�uΖviY7즭$�����G�Os��ki�_|2�r��n���M���DS"�s�j�5�SB-�m�����MC{�?�#Ԕ(����l�P�S64��m`kP��o���;�M ���IDx�ȇ&pAi<�5=Ի���7�<ͺ�|�xǎc�����!a�u��������N�Zh����Q�<u0r�p���I��Rp����Py��K�����
�S�\:�ݓ�̛�%]?�'�9n�_����S�!ʁ.�4��@�6P&�b�i��#a�����Y���Fc]ma�AQ�}Ͼh �0r����'�5ו���r3��{u��������p�^�nlG�NM� ��
s6*�Y���y��=x�;��c�!��\1��� ��
L.�hn��.�&E-f��A	8pBJ#�$�F�r{�iE���<��;E��u�""�nXXV�u]�kݼ�q��,l��k5\�Vw�y��y�]{#�.�ӧ�a�6���X7c�?��W���b�[e�LM�9_2o�'.����Rg� ��x��38L�ZTp�������]��A��u0pBL*ko6٩��	XLW{5�@ �0r�wcB�!e�x�?�2MRO���rj��t=!&+^=O�.̓�!��\1��'i�q����t�M&�h���95�y���?��))�6b:��]�.��nX4]v�Cŝ��9
�A�Z�urg4����D��Ѥ�O�������p���r��zZ�{X����M�o�%$�	M^ ��9����b�s ��Q[Y��O��J�b�ٯހL�L̜�b���F5��7�X�O4�A��'�y�RO��Ԅ���ŔZ����Jь�>��`���#����A	8	*�R㝟n+u���\8!^���՝���ؚ8LM�9Zɻ�r��7����L�F3oS��O�����nl�3!�x�5׹�L��r�us��yְd��ylkդ����pֹUǚ��|$��;�_�u	]��!&AI���q&�+��G��&�!�P�!J���mMָJ�b�ٯ�3L�����O�3ېa�=�M澉>~��P���˲R%�
\��KoO���":�
�ڳ9j���fr�hd����_>~<w�Rg �����O�DC�8Ҵc7Y��O������0���aDpUI��:�F�{������.��!'���u���J��b�W2n��]<
O�)59S��m�K���>7�%k �%
L@I���s�;�m��s�n�ER�9��w�]� f�8 ���I?�'��Gd�m�BC[�k"���	I<�m���DC�8Ҹan`@;,x�u|�p�$H��7�xYFϷ�H4
N�<QE�!'IK��a����U��{[�G	y�c+�7����<���� ��G�L�F}1\(S�Q1��<H��ݘv�S��Y�:�O˸�XX�՛H�K�ļ�Mν7��7�shЀ�����2�|���&#Ws�m9x4���uCJ� �=�{�yT���1���.=kl]-��n�zz��3�{[�u����5�@�X���L���f�\ư��n-Em����5����D������\�]���yu¾��<m�9�ܘ�i�	�2ۍ5�n�3&��1�85��c����t\�i4q�v�.�-781er���k3
�t).nS%3�bx���q����w���w^���9ݞ;Q��k����~�0W0���K��J����[��60��ji]�;bZm�9>�~e�{ww�� �9�8����lN��LN�5��&�j�%����>�v�����&�Rg �
I��Zg��ѹ��oX7|����w1���u�W{�pN��s G�I��sP}�-8n.qDo3�BN��#��e�;�6��މ���ʥ�F	yB���'.��
L��A)'�(�q8��2_,�a@�8�<t�BNlT�#��N��LO{5�M`�]�]��x���olG�����O"��Rj���v�󁂁���4�^܎�"3$��ᅸy���>�G�F�$�V_1ܧb��|�@�v��C@=u�nt���^3;��b�c�;�ub[Z.�;"�D!�گ�	�E�G&IDx��]ۏ�\1O	�B�����Q�z�SJ�SLg��=�x5��A>j��9DL1=�!>g�p��zn���U׬��ˮջqcq�g��s����(�	���t��k�9���{R�ˋOYؖՁr�-�Wn�	���v�/Ǉ��{ö�������z���co����_� �dӃ�38�SX��S6;޵���>�DA4�� I��)0	'|@�_k	��敬�3H�̓�9���vX?�;�
L�����@���I�Rp�ZQI��wUp�\����A �����5��+�>�u������2�ƞeA�J<�Z�-q}=�����!fn3������-~	�`���!%���S�g���e��v2�5��i�M�.lj#0l<��]�a�H��ra�}��I���,����
L���RO��[27��̓�9�����X�7/��70{�7��p��� ��i���LwV#�����������]�OFS�E�⛈>9V�A��pRg
(���������Aۺ�|�4h|�c3!�ag�����aGӱ2)Y��a�F�\�E�r��J�ř�kbR�J���j;��WMt]�r�yά�B��r��S�;VkM��Һ"�+^
�f�iࣕ��)��;�+�e��Ǐ]�����ٝ�͍9�۔z���os)t�E�B�̛hV:➪�ɩ ���!ބ�)��q��[��}�J �eǕ���"��eV������G��{�&��j#y�R�G`��l���!�����F먕��@�o;ӏ��m���٪�;�t�e�׀m��mm*;nR˥�I$h<���aE�V���-B�Z;݅�ݽU�[3$�n���+���q��uLȥCb]�v��.���r��.u� ��rv:�C��36��q�����0����c���UɅ�fj���_u�R��fes�tmi����?k��:?V�-��7A��Q��n\�{�U�M��[|�#t"��dkۊ÷�}.�nç�:n�C$�w�=��a�m욇Ev-��b:�|o�7�=�d)pYS���v�bxWV�	�C$�PS74� AC���e=�*���0�����v�Lѫ��
{D����m�dt�(�A(f��9қ�/���[��`��'D����u�ڊ�XQ|L�+ݖ���7��E�" �Pé���4�څXy�&S���+���]<����O�᫰՜;՛�i��
�a��s�����(>5>���5˯+����L
�κ��"����t.>	�k�'i}�o����VrVbe ��)Q8X�z+��;~�qF��"jQԏ/<�ia4�4M+�4(�8<i�$U$�?��AW��O&x�h]�K���G}��ɹ6�m��K_=��?m�Jc�⮯XFE.N��/:+cf�?P���j�Z�W��^���/�Gl`�.x^66�Qfu�*���y}���Q�t�)W�ۤ��*�	�Q�}��"��,�̧�EA}��CB��]�R�WL���X�e�����E��T<�y�.e�&{������9�⋊.�'��H/�b�~��i�`gù��K
�v���W>#�`E��_��{m�ĊL�*���E˲�'a�%���ű�U	����Xg���7I�7��#�'�>��.�|�P *g�e���r�z<�V%���5O'�C��Y7gh�����@�ٵaS7������.�ّJ=�EKsy3�$sI�>Bk����m��ӿG�=Y��7�艏�=�s����)O
�rA�F��6m�׺�s����x�ٺs#}��q�8c7A����^=o;�<��羜~v�������,� 1��DĒ��� ��}�O�[}Ϫ���F^,g��o��������>��ϧ⟴�2���X]\�� ۷!�Z�v��sFu��<��c�s�)2͟�ׇ޲��𑗹I������͓F��΃3�Z�!�[�����4ǽ�8��E�2(<ʍ$�Ѽ++f�� +��>=��d6n�Y��|�8�1��>46�@ �T)0������^�r*T�@�����	(����Ƭ\X2&E�l�D�p�qX!��qM��*� bp�ٍ�����cP#vh�d��7;m=�k� �9@�w8p�>V�6Mރ<�yc���HUg ������˯j���=P+\_vM�9+���x��o0��eF=�u.��GC���hA����9�g��5���7AԊ^�9�g^��jenS��lB��=�T�> ��<w��͘�'31��)4p�
�S)�o�xi�߰��#�� ��p�n �����L+��${��; ��LY�DX��[�N�v���c�yՁ4LKt��t-Q+�b"=N��	\��Fs ��G�O�ջ�����V3�o%��T۾=x�7_�k9��<BM��I����snۤ��Xh ���[�X�ѭ�3����?G��8bpE���z��^SSH ����NM �RO��C(��;��&�<f�f����E$��	(�/FIV]�k��U�1� �E�r5s�<��Sf�޴����.)������mA��\3*�d� �3���ǰB,Ex���I8��2/��gZb�fy�zζ4Ѯ�8L��c� ���BJx�Ȁ�Z�~z�hy̵���!#xSy��l�6�rƒ�w������9�ʆܗ�=��M
(��}M��nnyI��v\�&1�f�5'�R��N�����7ɓ@�W$��6G���:\d4�E�Y9�6!pUc����ք��R�;m�;��t���k��h(����I��u=��St�j�W.�k�\k���6W�b��W<5y�8X��`�nm���:F�v�!��qz��8�WQ�rݮ�a���h똲��*a����%)I��Ƴ3a�Y����\�3Sk�k�Ձ�\H����v6�M�c��Si����氮W���q�n��랸��Ӕ�ع��39Y�h(i��9Y�2=�����̈́9I�)C�w���ۚ�����ᅸ0�s��Ѧ�����<Q����9	(�y}�Ӛy�WK�0ph!O?���Ewͺޤ����-)�N+�$��p
M��ls85�a��Gp�����)(QE�'��P��{����cEOy6w�&�Lfd ��֠��k2��^Z���e�,�<����;��ROw���ۚXs��w���Z8b������@���7��(� ��$��QS����gH�F���U���j�Jn ��++��Ct�B��O�#��r����7��t�ʷZ�dYz��i�� ༉�j�7KMI����u���c���>���	o�>�{܊4BL?U�Z�j�z̷
��lq:�#�Zx�Fk�#��G�G�4�$�<D۶���h������a�E>C�{�
Hw�Qf�ކ�T܊[�2�a>�W�a��]�L��+���ٝ{��+ci��+{ֶ��OG�ns�n��� ��
	�3�� =�I���R��;�fpm�,>u�!�8an`NK ���QF��V�a�z�X�$�o\Q���I�����Cy2 ��x�Y���I[\m�����F��43��T4QO3&�7�1v��_��r��9�g`	�� ���٭�&[4F����� $1
T���ʴEL�����c"�� �� �D9I�7��n�&��}��,�b��]fx�X�%����݁ ���@Yu���x�~���r��Z kM�BQ�Nvu��m;cի;�:{�2h�,�-@���<��ie�h� ���!%<BdC��7��y[\u�����7��;֞5��H�s �z!���&�����.�I�E�!k��|�����FxT��g@&N ��$�7'�ۻC^7׍��m> ��?�2!�L��RO�ˇ�ٛC��A�#b�Bu-�6��#ܦ�i��|ߠ7nT3��hZ$b��Do�L=^���r�X������=�8�7��3Yì�O���0>9,�7v�.	0pBJ ,�^�ae�ى����(��4��9[\m�����������85]��͂,�A�׀B)�� �	(<QG̦�3n�xh���yxx<�6�n=�l��N �N��G�L��PY���8|X�?BVU�6lл6iY����x�+kh"�vF�e�7hX��f��?<�>�-����GH��� ��xw���۝�]�Q9�pa�:�m�-p��` �d�{��|���� �8'r���0ų�{� ;q#u��V��[��㨵U��7A�o�n7��1�d�;�2]�M�*c��ffCO2�1�A���ȕȷs[*�e����-�+���8�#�B334i32(�eA��;n��[MYod���pA$��ٚ�8��TNh�n ���ضĸ�͎.�:
�Jņ��;�h9s��Q.������/�ޠ�^k61�aݣ�'vj;QV��2��3���b�.1`�*T���������a��y�A�2��
�d�S�,ƹ����I�>�JOQj����A8���'��%$�~Y������g����Q덛c5�y��4^-w\����6�f�A����?��;���FYd�� ���A�N*�O[�gDV�=����R\���2L�9��fV2<�pA�V�<��P�x�pe�1[8���>�f����`ʊ�[������E�=o���5Bc+�X#Dɼ�'$�&��il��o�m%2�(�E��7x�r�ǈ'y&�JI���8p_�g<[N��P�f�A��!'��\�h���<'��{2x@>NTLֻ�樺�\�/�ZM;� �*1��x�0p
L�d���'���;����ᯝ���qY����K �w`G�I��|���1�\y�܋���T����e���,�%G����V���vk���弞�]b�6�d����i�fΠ#���oU?��x
c4�Т���t��{˂�e�pQ��5�8kR�p�n��r����3A�B0�tI�͒P%ur�z�����ب�o<�����"Y�y�lt�7��F��eК:k�k����M��mȻ�f�%^-];\��س��:�(�*1����n�[cK�h,���m�5[.NX�J�ckK�4�8���z�]'��[j�m�]���[3�����]�nE��ڦ�>~υ�ɳ^�%��^q�MuvP�=�*�!�4%�.62�6���n�����v�����Fs!%<JL6�?v�%P�h�Ņ�72b^�w)�f�� y0s����=!������3M����{|3\8}��ƈ����=�ٓ����I����N�90����zX9�gy� ��8)3��I;����t��`��9͓�^ֆN0b���7�pA�L̨���D���4Q�s�gO0{�1��	:�#��?��?v�%N���E��7�V�A��P��K��͖V3�|U뀕���% $̜��c.��5ýM_�5<�'��{2z"q�BN��z<AI���h��#�x�S�3�$3�Y%p�7�.�V�����u����M�ke�xwq���v�'����8 ��Ǚ��7��pd�(��cp.�mԔ1ja ���@!k9	0�Ff8�3�s+my@�K;E��2a��F͘�4г��|۴���6->��nj�Wӑ�:��|��7,oI���L���8�bL����<����='u��������u�����V��	��I��K;,��ܚMo��O�Dř�4��fc��h븧������9���2p�!&BJ#Ȣ�&��Y}58�N/�j!ű�pA�)'�}l����̜`��0���zU�p��-;�x����	(�"��'I4c���ji���o+~��J�_Qz��nr�ǈ8ȇ ��A)'"c�����׍����ճD4��m3ohǵ����9�sA��Ơo7XBll/�_N�H��>{Dx����8p�Wo�DEUlp��]��\5맮�=&=���ii32(�e(�O �����M Aծͭ��]o3'1D�f�NK�5�����0��T�˸��0ć��o2#��Nvn�:�4�j6!��QpT<���eo^0��������\]��ΧCqW-���,F�,��"���W�
Aq��)�M^U�H�f��I�xxxyl���Ԯ�g�����9I�q?�x��A$��g#CWa�t.s5�<��B́+X	8w�|�f*�c��
�dg�q��U��Fg�a��,o?�L���BO�)3d��0t9A^�~n�����8��'8c7d�pA�����!B�uS*��{�����x��h�H�ٺ�}\��ܻ��zζ�Au�l���v�5�)�mʮ�"84�	�`�q8rP#�'��_FwbWU3��ZSp"ZrE�=t�,2��|A�9�g�$� ���GMC�wn�^�X�Ȯ����������ޓ/»��� ����j�8�4>Ou.��SzA�g ��>I�I��$�#Zy��Ee���{�b�`��1�� �����R`��p���g%����_0�z�9��I�C/��7�+��N�rW�A9I���T���/��oKsA�S{�D^r7@�Qwu�;�Y�d��3��{1���T���n�����f^�.����Ӟ2�r<�7��;F��[hڨ_x��D}�r�����A3��́ ��OL��9��h�pﶵ�`����-<'���8� BN�BdGa�Z�31BDG��e�=�Guv3��K3�x�ņ���l��'nn���X�C�CD:�l>YO ��C��8>ID�ϝ�S��s��0�[Tc�;k�4��� cvx���!&!��02QpX�+;6F�<�V����i�|��ڦ�(�ؕ�79�	�ȇ&k.wY����!��^���ܢ&334hfeA�fB��7�mUN�=%L�d��ܮ	���p���z<|
L�ޮ�ҹ�2��G����h�x�2��~�%8����n�D�朙F�m����m���<�.A�N���3@a����1���o�ݰ�z�K͉\Sq�ǂ�D?�LIϼH"(!<)�b�WgۣzXi�����3f(M�*��(�,�K˝���\qNkK��7������΂�u��`˵vwA�Va���|�'k.�jϧ���[��-K�X�=�c���b��S�iպ�i v欼���&��rcS4m<��;�	��U꽻���vU
��Y����nn]譠�^�}\@��ԃ�upX�XH��6�	7�a�u�h���'�x�
k0{Ӡ�R�2\����]��l�z���̟�^Eu[��������_3�;2u9sz�_a�����ͳ.�}!�(K$L����nv�+n�����W1��(�-�.;��2謃�`h�SB�ꏍ�&1nS�;l��)�B�tď0�mbgQ�YL��\_eʕ���B�^�˧��.ڳ����-t��w5l�0���eD±�*�크��#�F���޺{Y.�G:����1��д���^��9Q��X�6��5��>s�� 86Z��)� �mw�����D�¬� �D�R�|b<���)�A�Ef�Ѧ�M7T2��Z\+�}�C�C[�n�:�T��a�(]�A��s�����5�wLʓ��eM���]��{C_a�-n�f�8n��>U�|Diҭ�#����*Z ̛�.\�\L���.T���OW\l�[7W����ޢ�Vɸ��z����x9՝Y
T*�U��v��>x��n�����y�l�mfQ�+2nR��=Dp�3b_}R9�}!��ւ�\�(M�
p��K��v���Gek[�C�������U(��X�;ߢ�l8}��
KzR�.�����-¬��)����������ڢ.{z�ʟ_` T�r����1�H����T��;�_=p�$Dgފ��p�=�E��$�Dڽ�*��+B3���"���~v:���FnQ��n�xSή���i)�K�*�D���ќ���D{]m�(�=39��x��QTU�!UEQWR��y�GQkr���\J*(�<(�
/
����ʪ���J�TU:K�UQG�O�Q{^I����(��"r��;�O$���̺�^QȽ3(����:h�jyDyS\C�TQ}(�as+�*���L��+SƂ_��hG�PxDW�dJ�A'��=�J��ʈ��"�
�����Z����Q���z���A�7�_x�Iy���.�G�%ʎ�O]��bEL�
��QN� ���]B�*�J�.����U�����yY�Q�>�A�)"������;��2��@5��i�.����z��zG��:��<�1��J�u�(� 9	�g��	i)v���v�)�MϠ裳Y7%��e٭��D����=�v�<��"��3͸���Q��Q�v�+�Vq�t���ŧn�lr���Y�!Lqb�vXY�Y�hƜ�Kn��,��.�Q�t��ss[k#e�ٖ˓]�`�ىy�M!j�R�H��QٺP`¶w��Al[=S=���\]sy�u+���\�{8�s*�k�̘Q��V6��IQ�5�h�
b�E��e8K1��:�#�e3���;9�;/H�Լd����v�.�!��ÍiN��ϣ�U��a:�ӌ�<����r';��S��X�q����c�ùP|ɍ%����rI=]�Ē<Te�At&&�*d7]�x��F�����|���L�8��v:�@�Q�fKdF�)�.	x��B�,�Վ�8�lU��Dۃ:E���^�%n.Ɨ�
�n���r�&�f�o1h����Ў�ҷ���c`.��ډ{#��,��;�[���ӝ���Փ�1�/lq���t�C.�v���q$���V*�E�>.�ٗ�Ϯ#�Y��u��.�CM�kq���#�n���")�e�v��vk�Ƌ��r�q/���t5d6�F�YG���t�pb��랹�$��rZ�dO;j��u��^����預�#L#�.�A����0��U�z�C�V�cq�����nR���>�����������X�4�0Bu�z�Z0o���vh��$js��jݞ�W<Ғ��
Yy��
	�S�Sɡ�^[���ʹ#v.�uL�WYX`GY��Ŗm`vn����:��Ogq��%"i�Í3k��Ub��Bs]]=r[���u�z�	� &����V%x�6��s�Nn9
+a�׎+�ŝ�P��G=W=qTՌ;zMӹ�u�a�nJ8��͆�]����E5Z07n�T4�m�h#uu�[����qkuW�t�R�g:�f�9����Ӻm珜LJ@�\�3,�Le�g]i6k���)z{F�l�1�õ��=L�kssa:��]��ɤ�`ܼ�:�۠k�v����I�9�ٝ����#f"jBSD���ɇ��&�1q�n��I�j�s�8ɰ��B���[r鹱cu�ӑ`� �ݔz��$b��Jm]j�5am��R`¼�h��Q�+��InDӮu��Q�v䂆�1=�����f�.+��Uuaf�˙�Wu]�%(]���f2�?���-�茳���AE$�C��:mcU5�����w�D�	�/1ll�n�r/v ���� ��B��q��/Xe�Rm ��xw���g���ɜᅻ��%������
(����rO>��|�Ñ�E!&BJx�N�O�2:�:Jd��;^�%
�qy�+�n �8�#�&�ǈEYvp������ݩ��}أ�Q�AIÇ��t�ƪkz������d���p�>��Wz82�#�6�$���I��Q�_l�_esG��w�4���k��4�q�2g4an`|rX�qE\Rp�s6d6I[�y����63ip:�F�3쉘�5�Њ�#n��l�	�MX�v��ߟs?e��FYg��d!%�Vַn��{x�ġ+Jn ������Nkψ5��1��
I��9���c5�_3�0�����&q�PS��'m���3�u��7730�u��;\�Ff�9g��[���y�Y{��	1L��s�h��U˷+�Ar��i��L|�H	�z|>(�y�I�n�5�SMV����{�[�	�`����!%�g9���y�;V�+��T��N.x ������\^I���93������������s`G�L`���@L�}�y|�y��s�[l� $�z�����W׈�J���@*q��U�1E؜Q���g ��O �8�%I�R�*�!�03�r��ӭ���U��բw�[�q�I��Q>	?����ns;�El�b�C,a�ZAut;X�jα��l�q!.�C1����wSv46m�l �3� �����ǝ��{���&q�#'8c7r;��[��!.i�)�{����8!%<��c�!�n�!,��-?�
����nW׈��|����@�O�&�AH�̇w�u'�Fsy�����̏$¼A	8�gPg��M}^�l3��j�k6�=�&����)M!�@fQ.�:�]��m�E؛s/����VT�z���]1,�l�(���i(�l���� =�&�Z�-���c�V���[��`�N�$ޠ$2M"{s*�AQ�j�����gRN�͝ǟ{Bg22V�f�}�ȶv��:���K�HFff���2���K2 �Ks�4�9��=�_�nW���|����<q?���A)'���ץ>��o^��8!j٢	�����p㠼��p����խu�#y�
Bk�W�=�,�~�F�>�� ���'���9���ۜ�	�nۃ�]�"��)��Z�n��	?������#2�q�k�{Y� �s��ټy��q�'%p�nь(���sS�^�ΰ�["�Dw�IÂQ��L��M��^[y��jSƵ2W���e	�L�&�<F2!�I��$���39��0������x���<l�
N6e5�kSMi�zn�ݾ�L�.@���b3��] �.���3&� �,���ٽj��gn)X��#����k��v�ݥ�2��cR�d5tq²lf}� �����DzO���RO ��$���Y�T����~����Lbᅹ�q��F�.@Jtn�T����l�y��N��*빵�47����ϓ�u3ͻ��j��MMMwC�ߺ]v��B��-&ec
��=�ܯ���|�����m�9^?_$�i3��G��Mfd��x��(��"�֍�kd0����78l�k��55��������d�pA�p���5s�:��\v��i>�i ���<)�Rg ����gMd;�f	�3�kc9�;�ɜ\0�7�9n�(�� ��8!%6�K"ѷ�c��#��������p*���i�}�o(M�f�U��T�ٽ���"�kϵc�!C�� �q^(�]<yN��F���nH�������p��SCy4��mgz2p��J�x�DG�En�t���d����p8��OE��Z��ܽ�^��|�
�;�[� ��Y{3�7��_ot����F��z���P�;3p��y7難;��t�!���J�����e
�Z�[\ �C�&�6�����N;��7m�F��A��א�e�X˚q���]m�]�}�f�=�yV�1�E��4��76	Js3�,V���;������ՎQ��	���{/[.��;8��P��\*y��L9{c�uh�������M�j�9�;��\��[�\�%�`����٢卸�6S�cR�cJCZhmk�g��|��c�����N\�Uv���RMd�3�	����K������~Բ�߿� ����I��RO�w���]�2qp�oE?-�uN��G��>IÐ��@#�&�������	b��jo=Nv�gWٗ�o�0�F�"�2�h�V�i=�ɦs��̢&0P �8 �'�6�eé�g��O��2��=5�� Ǭ��y2�(�$_/���%4)��?٘N��檧��S�g�;��,��p�n>�`���f��co��Su]��[#u���� ����!%�5D��3�O���Ƈ����h�K���(��f�}So!&&�䓕\�B!�g;;!ȈL�\@,���Y]CBR\�abnhK"Fh�cR:f��T钽1�(��4i<�#3(���J4=M�,�#���&�tF���0^ �2e��4��O2�1�3"9�y��'`L�p�
5�meΫ��0�1�n��� �����Q���an���9ya���)�%���
]�#��M�J�z�&t���Z���p���g3�=����sY�A���|>�<���K�3q�0rհ ��Ef=�C��J
f�p�=������������ȴ�ȭ�4�G��M�uaܙ��e�u-˧ɦ��^��.i32�C̨ƞfM32�f���s��t���ha`�*��)8v[E(��4;������p�@3���_n�e��.�:��
L��x����3�"汭	堚\�����6x'����3w��0r�� ��?�q;����іm�
{�#t��[�s���[�Ooh�������N(kvV0��m�}���v�_ߤe�S�Ð�Dx�����9�y-WO�M7���I��h��O����r	I< BM�&<Ck�ih�}}B|v����e�ED�s*~���@>3��^8rW��y��}ޱp&���4ǙÇ �����n�Ŷ��r�u����w�w$ Y[�Vq��V�N���[�Y�F�V�����״A�T�զ�9�\�ʧ`EҴ�]��4��{������в&3f���V0rհ �8!&BI���Tu�������\�m�G�OꝎӜ'��R��i��n ��xd�g�Y"nW�ķ���	3�|R`����&��s����F�����p���i�l��0r�$���O@����[���A��v/<��2��.�NkNݘ֦⽮�;s�2��,���֙h`;�3C����k�=��$�X$������<D��b�޹�ػ͋z��Pӷ�aD����Q���������2F�����T�n��<�"�eSM�q�x�0`�Bj��S�noە�:=s&�-�*�(�h��h����]�sA��(~hyB�jվ����e8�'���!%�"�������]e��h�D?��g �RN[No�=EdL<f-[�V��k=��DNj�5�Y��([+O���Y;:ȇ�rg���д�����B�l�7�jǓH�/���+T���ǅ��5	��aJH���{�-�.A�p�$�@ QpBLJ���ܺ����8����]�J2���ٸ����"��A$�$\�t�j��X��]k�׈b�c���5��q�Psc�!υ��EU����XA��w�ǻ�=,���Q��f@����3���s/=��s�Y����9�8�����u��y���2he��PDT�cOvE�s�xgӛǷ��FD��bᅻ��k ��QD����#��Yn��8א#Ȣ����	(�QbXe3�8����J[�J2���ٸMͼx�!�M�)'�B)�ٺ�[�ȆEo@�<\���m�d�L���\��{ep�L�>���pT���FVG��&���3��$��
O�&p�2a�m9����q��4�bjk��NUz5��	�Y�y�A�2P�ڵ��kC�}׺���4��K�?d�<��5�$2i=��j改��U��ȯnL���9��>��C�Kf�T����TVM;�[7�|!!r��r3UjG1��B�֛�jy�v�]2�.�h˫��V�������mu㧎8��M��:�G0W�z9s�];F7'6��n�m'&���%��is��D3ź���GkEV�hm��Ac�������;9���f5Ե�qS�$p)���Λ�����:�7A�-Je�M��{�_U�������&�7�۵L,��i�u���k��~8~��m@�v�e�r��q�ְh��qnfc-������SJ*�������U�~KCy���ȵ�<�T���<��eKM��z[$=�i�����/�(���CɓC3(3(�њs��v�`Z����"�Î|�N�T�_[uԼ��S�q��E�!%\rbc��|����nk�	7�8d��ROJg��f�|��eY��M�O-��c7��k�V��R`�$��	(�ݓ���u�+p�b��y'��T��\����Ó��I
	�_�)ܮޚefe�f�5���3*&7�Dc��y�NJ��H���~����W�ήb{�+�ӌ/8!$�I������n#�I���u��fQ�Յ,�ͱ�3�7�5��7�يA���x�h�즿|{��X`��1�A��-�;��m6e9��ţ����k�E��`�e��c^I�ITy&@�Ms��n���P�4�K�Fm����Fެ^Q�=���E�[>�67�R��k�'h�L����YX[
�r�zrfc3/3��  5���O���ON|>�<���CM��q�x ���e⼢����Ѿ1�����u����G�`)'Z���!�z}�ƫ����'����h~r�0�Pfd[Ȣy�k���c����1Y�/�^�����U��;����X�Le�1p�n٬�V��=M��������32fmhi�Q�!	(i��-��<�o�]�i�M��򢼾�W���4��dQ�T��2gf�k�}�g��tk4��JX�p��܂�\cpi�u��n�!�P%�5�+Q��{OR�%��H�YI�Rp��N�n�U�wE���l�Y]��v�������b�!'&�A)'�����cM�o�[9�׆��7{�#)��f.�����>Ր ��8�!wP(H\��"��	�`� ���IDx�'�A PB��F��p���k��7V˃��8��Y�6h��c����j�R�nۖ+����#��U7�3v3n�<�y�s)�^��C�z�42]e�K���5�t�MO��w٠	�+ڵ�غ=�wrV�C�[���f����b��'��Y���v�v8�\+�;��1*&RW�؞�m�(�9�&�Nq:��8{%e&,wZ�:���n��sja����|k���*�p�%�ϻ-�`�W�3�$�0YxZ�d�D�71��֦�Sn���|rkƳtqu�
{��+FKGJ����X�g�W�s~a��}��H�e1Y���$f�R����5�ƛW}su�u1����_fdn�gA COE����2�J�:�P[Kw{-u�95ז�5פR/����^�ֲf���T\l�ָ�f�����T�J��3ӌ �U
��]�z���[Tt����,�M�̹�)��������S��]�.�v.(ۘ���掉ӝ٢�b�B����9�ݽM�u�.���9>�"��E�tE]��a7��ӈ�4TЍ����b|��z�3��� m�3����3�f�Ԇ� x�(���Λ��w7F�l�I'w�����"��O:�7V/�S����:aݙ� ���֮W�0���a�D���`��1]����g=�W�VJ��P�>y����E�cg}o�y.��zy�$.�B��rGml�]Ө��
�	H���Is٦_��$ �-���H�U�VeE��t��'�\[�S�8��r��Pmoo$�,����N��/C�Q�����m�/~st�xt�tkʤ��USll*��	!��+\H�0����wba�Y�.Vb�o���"���p��<����$��!��h~���W�l����/�7y	s$�
'>�DVx�mH�#,�$�.UFmst�ӕ�g*#�"#z��;$���jQT�j���@�g!�u/��y�jI�Y!U��{n})�G�V��ɢ��F�xfUd�U�=^�����½����J�!}t��y%�"�K�zm5r*<�!4]�/&c�Q����G5"������ə��İ��(H����H��!䂮����^R�znR:!>�yC�EO+�7�2+�j^f�g��Z��Rg=�]�i�Q��<��
���й��UyZ��)��]C�W�!��[	x�ڂB�e3�krthu҂����Ϭ�Qү���2��(�����{ǽWyQy�� �M�r��������"�Q�>��$�f��>���)��u7N'ʆ��f��nm��y�I���'�h�"���U<ò~a@��v0�`���t�vڮ��-<�{ep�|g	�t]۲��֦���z��I��$�I��)3��՜ú�iKF��x�>��;��2�x�\1���5���5d ���	0�������$ߟ��o��ա�&��5Y�ٵ���ݷ+�[�ڷW
0��m���Y���/��FN�BJ �"�z�9���#Ә�F&�ٸ��6/sdn�kYq3�JI���)0��m�+
���q��X���:ͳW��-=O{ep�L�.1��Kf�K��Y�*���G��>x��$�A ���mgv��C�3+2�x�Z0��5��ud�E�	0rQ���4n"��L�C\���E�BdCԩ�ݧ��l�17��� �sO�27T��"�*R痢�0�qe������-3Q��^���~V�:׽�M�w׋����o�5�t�a^cۢS�st�`Pm�a6�A�S|�x!�)0pI8��?}��_��E	wOI��t]���U]��2p��7���G�dF�"��i�����)>����Pna.6���ӂ����=��1sӠ����<;vƦ�@3)�}��$���I<�ݧ{�2�x�\���3-b�v>�P �!'I@	I�m{��q���p�uO��=*�����9�E�u3p �sO$�pRe��a�IP�/׋0�I	'�L(�dp�7��6T�2�]^R�U]�ހL��^8	'�$�t�pC��fgmk�y ��v0	'<�o,l�̫�3�f��l���8.�������R`�����IDy&BL�$��V�Ҧf���n��gm��wG��e������)?����I��9p���w��ل��w��W)�Nj�G-�(�P"_�D�s$>���R�g
�5n��Z�����颍Nw	n���	1�b���ṐC<��a��)���e�t;�jٸŤ�aL㮚+l���l{n�jQE�*y��;U�\�N4���NzW�2��l!sq����#�3�y�ݛQd���-�\�X�]&Zǋ���bf�
LP��nc����0�&�+���i��Y�a�C�n����*vE���v�[mϒ&����������n$��ME�׫80AR���������f����9����[f4��Y��s����s���3���C��6�� ���� ���AIÆ�4�3����M:��l.��w�fi��C9�2�ZMfE��4��M3�7��pOb{b��Sy�js�3�5��2�5>N-���� ��I�v���%��B��;�����(��2�����"j5�ĸ��dMG4��,��6!M+��� ���<���L��$�I���RE��7��<E�8��A	8v�5���n�zr�Uw���	���q��7�k�G Ef��Zo8)3�$�����ĦBM�۔3��˷8��ݱK*����h�`+qG�aD�����Ĉ��Y\��P�/n/��ղ��"8Iq���+su��f�+33<���K�	T��"��IP���[��gp(��bҺٸ��٭���o^OF5�G��ƞfM32��(�n�V_Z)���B�X��F�˦����&"!<F^(8���J��x�	�SK�3R�%��L�lS� �����8��!k��k3�5z��U=���LV�ȫLy�v�*<��{b�#=�˯4�ʉ�]��(;��&N-sq([P����1vD��O�����7�"c̊���!���C^����yd��]�<0�6�=0�o$ު췥���Ӎ�SJ�f��EX���(���:��7ܨ˺���+�D��z�~>�'� /\?�8ֿoI�u=���y�Lw2�D��/w�̕]�m7�W��M���˄���8�hJ/c/tl��#�Ԙ���t;D>�n.����V�����-�މY4�'3���7I�lw+�/Xh琏=�&;�F]���]�k/(�F������8��k7�\�N������ ��r�?�ݲ�����Aû�+5Ӯ��~W�o.�e� ��w*���V���O߳���q�᯻8�L�N�'�
�VL��h�X[-n��$�]N��t�����.��K-����,����5fdY˪�ܺ߇��[���F^k�x������A���2�2�(휄ι��En�ؗ������󂵜M�?� j��蕑A��s8noX�0��~V��j:o�X�����Wt���L�kHffawz���J�/;�͒��4.�n �%�i��i	뷫���Pn��g��6�uD�=%m	U۷W7k��X�v�,Q����p}���1;��� ;� �]�Vq�s�~�j'�¹�=s��NƷ\���m�x���&{�&����W�?{��\�y�9���2��;r�z�/�����oϒ`��|"�T.��An ��C���#.�I�q�]�Kv�=;�����=3��ow�K?�)?�;�������3��{V��j�׾�\��7niM��FZ��0�w�]��`�PnZ�i�ꘉa�V��������/�V��Ό�{S^_e��e���c�+2lIـ}o����VU�wD��s[Q��j�t|�-����<��<����b��)GwQ�wt��Q;������_�����\__cw)Ǩ2�9�1���8 ���A."L\���~�zE׶�8�33,������Lp�oV�"z�]6Y��j�6����'��썖O~�=z;�v�|�J��7�<����[7�pȜ��|�*�h9��;�����c��1��ɳ������o�8 ���&Y��ڊ�K���pA��U�pe�Ѿ�l�;]c��a��2 �d_�������u�w����3�����VS� �fB;�	w˸R���s�7�6q�+�����/�.4������:�f��r�&q���kg7��h7�X˺PwtF]�w]c5��+���W�6H����Z����v��^��ǻ�wL���_�Փ<}��:��u.ͧ��:���B��� +om��,#M��㬒A�nh�S�:��K�u��Z�k�cn���������N�|�X�=�@���]��N�&�=v'���(��e��TI�%��c�k-t�4[eT�.�KZ;:�73Pj�ltbW4��GT>9��+6����g��֞Q:�٧��'b�޷nE縃v�8�㹸�ޢ'���wUt����8簏�.`�q4���sU�ۍ�z�$��8ńe�ˉe����|�%��孋����lq����@�U�l��6��������v^�7mnݺ��c��)������=������Z��u��o͵�э���H �ݳ��ݧ;���ȕ�1����5���|���)�[c��w�;�#-{����޲�y�������+���/2��܈QJi�m�qĳ�BO��a��ƾD���`�0{�**b�T$4�
�S�����=VB�2�NK�S�a0r�p�]�'wwuF�����`�w�D��͐/4no:�i��+8c7M&�#��y�Vm=]1���.��"퀻���������?�$�Z8vD(�4κـxop	?���v��C�������Ͼ�}y��a�6�]�6Q�;v�<��9.J0 'k�vF�t%	u�tX�a����}��]�;�i�'�]l��>�`��}����-���"�Ñ��qwwu��A���sr��{��Z~��屃v�T��v^����9�͓`2��{�Y��S���q�i���:Ee��}3B��Sv�q[��{z���� ����A ��������!�FG��NUz1���fd �袥��>�e_�U!N%B��T�UR�E�|�x�:�쩤;��WTι3p �ĳ��p.�|A7l�]�����^%4��gc	 ����N?s"Sjڵ��nc���18i�A���3ٙ�c��S��T]Ȟ�)t쯇�B�?*�!���\`2�h�(��.w�d4Hȕ�1��&)8sv��
*Xۘ?!��HtNx�V,�j�+�d%��.e�SB��Y��"F�Blۣ�l封(���<��<��Q]җqE�3��O}s�%]S:���vfu;s�ni�R9�g ��m붟|n�9c�g^�<ᥪP��=n�j�FOq���Έ���c9�Ñw���3ؓ�8��n�ԑG�Tk�Q�]�wQ5wJ�����7��.6M���7/RR�
�{�<��w;jtN?���TX���+���۸ ����vu�iɢ����Sw;�.$)c�
�0��e��#&V|1��c~e�fB;�"c�F]��k7��S@�ma ������ݿ�E�g#�.%]S:қ�&%���m�-�z�s8 �ߵwQ�;�"cWp�wtzV��[ެX�f8>m���޶x���<ь�z���o]���OB�ל@�-� �\uJ�������\�s�W�s/3A#��3*��4>ηl��E�y��g ��p@խ�ܟ�FL,��G2,�T5F����j���#.艗qA�wDL�]��f�\��b�V�U8bo?�E��ü�%]K:���9N�vzPm�D�� �;��Q+}�!�tA��j�w�>tո�yؘ��V������pLc ���?���A��Q���2X�s�cYe���A7l�-e���<Hȅ�1��9�0;N�qf�ul��l�lE��m�nS;B��5x��lR���c<DڵX[)>J��*�]�mc�2�6���RW��vkP���(;���=��wDc3!w ���]�2��s^���$_��󉠖f�o�k"R�g\���c
�B���	ʨHOw!���t��斞��?���Vi��]i�i���9��WY�b�;/ �\rr��iV�Ã��N����2����^��l͙Mj3���*{9�2&G3���{y�]��/��wuӻ��}�}̄=����A=�y�-e���dK��1��&m���i�v�{�f�]��#y�d"��#.�.��._|�����Q&sWQ
.��u�dJQl�7A�g�-��oH7l�]���5`���7�[uS ����ݰ.�8m�d�:��+���@l�8&t�+�Q�"��bawN���1��1�u��u�{j+��3��Z˻��Ȗƅ�9U�?7DLe� �艗tx�٢X�a�f��2�L)��̒�9H�N]���T��a��9���*b�z`PR�#�B�Є�w}DiZ�36����*��V1�wCC����C� Tw{ se����96;��K
3��D'R���piu�\�ރ�*�{��Uo�_r#n��Z�v�v!V�7.�*>��E����:͂;�8;��2}�`k2��Ak:����t��t{2���"Ľ�μ�r��vWqS/�0n�`��ld�{gb�Os�7�Y���.ü�R���[�U.�V��m%Ԭ�&�6f�q�����9�\�|m�n� `�P��|�����l�r>�f�bq�{��sCc�v���F��5�/7�=;C'N��%�^]�����uƁ;�Y�W7Ky؈��X`�(d�Ona��^+Gn;��;``�E"��z��0Ѱ����ZO<�V�t�3qgn�O�#(%���8V��<�0^V`�\%��"��;���6�Ѯ�v�;�f�w"�b�����;;�S�bl(ޭ��2v5�`'o�a�R*TP��e�:	�vb��j����w]-J����%����]����Ӂ�j�X��:�Nae^Vq�����۵����=��ޣwl���ۼ����8��;@�[�+q��F��YGl��݇t�qbmΥ�p��h�i��P�KK��ae�Z�';ڇ���'ua�P�Қ�ۍX��ͮ� W!�2!v���m4�l�A]�I�R�V
�����n�;0e_	a����ld�n�4���u pUА�[r�΋�;fZ����2�,o�>���ѮW���+u��:�3)�TSMTg�*#�J�$���W	�&�^&�^S7<͙�����>Ij�в�E�I*ОKD$���9����+��-�e��ȑ�n�h}dt�y�=��O�PUqyƒ�"PY�E�n�*����>|��O&҉�.�=�Qg�2:��F��5*b	̫��Y�I�
'��y槔���Ȣ�%�2J�pѓvc������(�!W-��uK��
#���f�Dg��9��vDEUZ��J2�44��ؒ�W�xTEU�`ν�TfA^��AM�yyD�9��L�¿V�Y^Q$hI���2��$�(��#�eQ�xG��D�����c"�KX��Fa�f$�U�<�j���yD^���S ��A{�W�k�<���jUy�Fa{�����)�Έݸ+�uM���Pw��[�õ��2)�Kk;�G�rZ,d08��2s�q���P�,����	=�8玮��#�u �S	�;O��m�zx�Z��CqO��nό�/�j���ضs� �7n�0�4��٩�E�H��&s��C�#q���t�h@���1���i�bY��f)�8�0��[�&�����/B�5�'0�dά�Į��Z9�'8ۭ��&���7-�۲{8�������)]���_�a"_	s$^֦��%0�3[6�f�-�M�gYdg�4���M��*<����ggvuu%u��0
\�0��P��E�q@�ۍ�w.�-w3��n�v��sC��p�4����]�/o)/����m���ʹ�;'t�M�]��P	�.�{���<ۗٰ7V� {��ƕ&9�����u&�s�Y�v�+���Y��6��1vhYK���sDa�<�}vT��l���=^�.�P��7���1�8��	�9dm1�X�W�OKj"G1�&+՗j� ��F9���Io�]�Kv�q<��n���k�W[$��G V�7U�����O�\��/2���nC���Uv���O.�Cƭ�褸��D��4��CjhYj���k��74�L]� ꍦ�XLf�P��H����yy�%s�m���%A��tl�8���� 8�0W�D��5ت퉥]|�ĸ��E�^`�q4����P�ɥ��<qx*���f��\��@�fC3vVB�W��e� �R�{-�G��n<mn��"��Cm3l�^cy�����幅ѷ��k^��5��l���:�R�s��݊�ܝZ�i��n͜Y�f�ݦ1yxۃV`OA���;��mȯ������5�E�O�<�ƣz�v�	�ڡ.����q�&R4�F���$�����1�)wF�˴��K�jv�o/H��epҋٹq��[�y܌�.b����u�[44fل�����Z"�2�&�u�q��p���ź8]�����O�.�]l�:��Z�\{���;��Y�k�נ熫v�ZK��8ǻc�޺,�ec��":�����b.\]���Z��u�<�����:��/r��}[Ӷ��g�u���4���'<g��㍺��H=��s-�n%|�6�9��n��1Bf�簰"RY��ip�q*Y�ͦ�e�c+�*i����h� �'������{]�i���xP�f�nd���/LEd�GfZ����:���K��Pn�Dc]�"e�"��z_{��o1��J-�rf�wzw��o��]��O�Hj�?He
CJ��w���W
 ݰrۇ��(ή�����lP88&��Â.�E�1�ŃA2�ԝG��Ms�w�4���e���w�˺{�w�;�{���D�2���}���wtF;�~C[���]n�1�d!��|.����q�g����3p �xUP��-/�:��:z�x�B�HQݰr���l#�)�32E�v�-�ݞ��y��P9�	���p�"���>�hJ�%��wz�Il�Ú�����t3l�	\:-�]�j�=���;��'X�k7e��=��Z�j&4w�A��c�B����-�N[ �9�������0H�����DOy^C��f���{׷�F��?�3n�n��b�Z��m6eMU±��+,�V�=:�б,��k\ǵ�r���X[�����Z{��V��pj�����f����o8�v����σ]nm�[�'���K�]ʄ��V�cz��J�9ʉ�ecWp����n's��0���T3	ꊹ�/Y��#*?A�e��]Ȯ�GwQ3�G��j'�����?�>;�?������[���A�99����0{`��O��r��z���.�]���2.ֶ;��Y�/�*�[�c�DUe����ge��ݳ���T�1�����p�(���[ -�R�f'4v���r\E�5�Z�5]'���q>���נ9�Æ�j;c��vR茨�'�U�b2����0�A�p3��.��n��>�g���޳�ö�P;�q3�@7l��sq��'.�%cNp�n �bX[����ew����^3!�������`�]�����c�ñ�nP	1�U_�����o�S�gW5�����4�{��3ģ��u ��-� ��X��6V�bЛn&�>�q�F�1�dE\)v_c7��fY��-��ij��E�?�U�c&��
"e���v��t+Q��+��De@l�8 �`�u_X�j��&��_iC}�;�������('v�=��7�J0�{: ����]mټ�������NU����GwDL��k��������|���~?��6�hh�.vy �Ӱ��qS�:�&��M��;6%]�O>�����v�{�����_�LUe���U�t@l�",P��_*B�	� ��"֊�t�y��h�����-p�hЭGlO���ʐ�Ϡ8�<!'(�ѲY�r�����3�8��v�]���Y���0��W���̵���#Xep�n ��A�p�7l�v��l+V�?
+f�:uK	 ����w�����Mލ[��&*�K��f�LK?��z�7$��Yau���@�SV��a�sBt�N/=��f�F��s@^FY�����ͮ�[���<�}�6���N{�O��d��?xU�&���8"퀻`&�Ãv���b��F�*p�a�x6�s�xL��ǌ��8L��j�����VB��VgUQwC�E�Rs�m��Ԝ@I�/m�x��9��G[*f9�2�����c=e(_"���QO2���޾g{� ��\1����U�Y��s��� ���f��'wD�����ㅾ ������:���K�S.뱘����L�f6( k�- |oR�wtD1�p���o���s��Ug<��'���xˑ�Ì&�v��m��UHpT�w��}&j�\��N�P�(Pl�n���P��k��� ��b��}�9��#���yD�h��r�"�Ñw48Ɨx������V7/�8d��2���-,���o ����ו�z��گ�_�I*�^�C4˼|���<�w�&`{v�ە�+f��i={%\{:�u��>��O<�?���GT�(
�Ѳ1*9tj� +������v�!6���o��<<&ޠ6�O�oV�����/��qæ�/'�ѣ���� 
�B+]dl)Re60Rؽ]��P�Rpl�s��k�CZU�l��G��ӵٚĶ�M�Ջ��vD�CTOk�j��K�z�X�,�G�P�ZvH���`��mÑ��4��n�F�>���	qEV�t�`���������������뭣sN��x�5���y+f���Ya4�X&��U@Ã�=��Lbw�"c9�A��;�EYÕ~�^xD��ǌ��b�Z�̩1U0ܢ&v�D��]����d�g)��v����s\�A7l��Җo%�[cJ�ܚהA��wtkS&���L7�awp�|�"cWp�n�D��.�S��׺����p]V6`ɸJe�n3q��y�V�]���v�5z�S`Ό�a����`]�v��ڳZ���ǌR1�?�0pB�en���ɒ�����YFCb��U
/��ﺎ/�o��f���g�osoo'4����p�nbX�c����.��k��g={��8���s��V��b+X9	�*��Y��n̸�j�Z*��kZ�֫�YK�Q�a�@��EwK8�+o[8e�%-����,�l1�x�5����)G��g���]F1��+r�$�޴���Cn���g3Ps��d�E1�j9,��G6�m%����M�P�.u��3D}Ƨ%a�y�����CF~<Gyc��'�����j�+��y̑�Ì&�ۇ]��=�W��9V�<�HQJ�(��@kwU���~��D\>-�ː�[�/]��[cJ���bXE�Wtx1����,�'js��o^��.�hN ���._�;O"�s_�\JR�뱛�K8de����z�h9Uc}��.�c��&2�;�3yv��%X��빛�����2?c�Q� ˹E�Z�Ti�g�j��G&)I
t��@�VR7V���M�M��Yt�;iXm)	M��L36�'�=��6�z3�|A7l�6����+li\1��"'�v�4��n�]�pv�;�.�9n��`�!�����}�5:'�];��?�x�+w5�bR���f�A�V�pn�b��%��d@�jh�#i��S]�wG�2e��z��o��o~�,��K5���{�<�"�h��\7��u���c�����ZXU�j�u�U�(�'g��&_�Z��,����sNf�O��(����p����wuN�<�GLN���z�S��V��7l������a�9�W�P�^����sc���w�@c��FfQ��A�A�z�d'up6T�{.��-������J��뱛��8 �9�g ������G��B��Og�-����x�n;W�'W1D��f�Tiɢ�W�li��#�b���;���u�z����9�1�9-w2�����s��cY�D��Wt�;���t�T"��幮co|�1�|jٱ�Yŕ��[�ru����1�T��w��WS�=�L9��p �9AwG�.�.�\�0mW0㫢ڞ:�,�1a��7xc�Q1�qGwQ��һ�{�i�]Q^w�bc;� �@cWp�g�����vsNd~��1��3l�֌>�l�Sđ+2e�&���i�w��-�a����Q��D^��&�\�6�ndp���x�m
KN����ճ��(�,�d�"��ٝ�̑������/���zA�o9�o8�p.��*���	�}L�>㫹75�]㴮����>�p��A�q	��ZK�ߙ��s]�?�Z�p�ƃ�i�.5�x��^-X�nn�Dj��F��}���4<�_��.�D����ɝ�;��X�TX����)99�c�3)���6�B���8(|$4���p�]��3*#1��wk�f��
�3����AWp�����*��^.{�A��Q?n��� j��A�i�G=8�Oeu�V�E]�|a�9�����B�4�HiP�#�%N�|B�[g��%� AX��Es���y���[��Ӕ�B�*��]��V���x���K�^Gu��&r.��>7l}v��`lrF�ܙ�v��&����^w��sG'�i�D�n�]ȋ�C��$��e��S܈1��7l�Q ��`+���L�9Nfsv�tC�dD=x��]�{f�V#q�K���������I��=�.�A<U���-��[��3s�;�z��zc�ͦ����f8�u�aL]�U��L��In%�,p��Z��l��s�a��۞ef�SC30�m.]�c)H�D�{q��y�P�@�����n�� ���㈣I�+N*��e�@�Q�]�jq���y��X��f�.|��kf��;I����\@�n���MP���Ͳ��f6�u��'���'�e��&�CF¬����Y�{Y����7E��v���	I&�^딾�PcWآwu����+V�]L�w�Ըc7���EF�F>���|�1�p�.�A��9�.D]�Lc�b�F�a���㻃%���9I\+���{�j��>V�pn�$_x̲���Uk*o|�2���95=^aܫ���cZ�Kx�d~	��1���r'w�D�y�o~�h�[]Λ�L��v��p�[�u3e�����,� �i���z���M�8�n�3ܢ��]���w+o�~��f��y���'�6os��e%p����� j��>V�]��	�fz�z`�'��gP	�\2F����c������-��y��sYGi+R�U5U��X���#��N�2�34��h�J�q����Llk�hj��^�\��8�w�}�;����҃���_�y��ꆕщ�������,�����3��6��S�݆�l�'2G�1��V��m�)9�G��w>S-c~;��S�����[���l����A�n �6��A�p��e[;3�ך�3s�Y�A��(1�P]��e�Q5v��Apqg�biW>>fV+��/q���l��*��$(T��X�{�̨|0��[�`�v��>����.��1�����*Vt�3�-�R�Lˊ;�����]�w^d�/^Q���ȃT�x���GKv�uCe^3���oz=n�Ʒp��1�Ý��m��Å��}~�['i����]�ō�16�ͬSfk�p�efns���Z�55�:��������w�>�?f�۝�X�ؾ�n!�Z*�l��m3̥��wPe�D5w@�K:ߔ3�lk�����rpk�
U���1�8& ��Ñw{4ۮ�[����c}�A�tt�wu�6a�ʕ�g����*-�1?�]|9�$��=�f6l�g[
�^Xu\���]B�B-���uuv��&��Ϭf>[Omd�vP]�v��A�L�uywe=���\�R���N��fSx�[��0=>�&t�<�7�4C����^>!������@�,���n���M�n��0��*%�]��j]����Jr ��[C���ث�z+kk���fZۮdC�!��Mg&l�4�V!xf�ޕ5�H���h�ϲ�;�m1w���ww.��ώ	�r�����/+�o��K�Pݕ׸ove���[5�)�ݻ2NLTo��2�V��\I��VX�y����N=�j�y�Yk�#���sGJ��ל�v�;���j��#R�Y�($S̊�V+�|B�(���[�lGגKύ���'yd�#c�nu�b7x]�
�:���]�:���x �O�d��،܁�6�Z:oYi�n�&G�X�\�F���n�]Tp��c�~s;[}���S]����v�F{@JRl�7Y|F�Z;r�Ns��ۧg,�Wv�.�fj�����ܼ������;o9��ʴWnYB�X�ĨF)�2V,3p��RV��b�f�G�)�b�n3,�l�"΍����W���f����-gB��3���A�1s����r�M��X::N̡���6�VB��ʹ��]�om�m�u���3��,�W�k:�X,�j����D!V�����ت���u�m�ޕ�)j�%�k%0��+Up������)����u��8�Q�/.���|��S��C���UU�(�U'M:���U3r�d�{���S$��r�ܔSĄ� D���FmJ�������Sԣ�(.��2"
�h�Ex�/�r"�z�HS=�<�ȪT��U2+ ��(�z�\����eyR�U�D�\�L��-BҌzxv�b��D��!S2�A-�)��I���PJf-�U^2��x	�,K�u����j�I�jUyg�
S5�)��M������K"]9�^GGC���K�"�gh��hY�U�S$�j!EEEx�z�S=�e�aA{�ΙzE:���yW��:g� Q���c��e����$����c�E^^䮑�I���Eme�T���6J)Ӧ7%$$sY�w�OC�^3���o���[�7lx�!R%N{q����{��O�
ةP����z@��vƾ�U婛����A�o_T���rGz 9,� ��@!��"Le�"wtj��u����5��'�o��lp�]�в??�0p ]��.�Wt��~r����{�3��Hʹ�X�Ol,PE�V1��B9!1���0�3���&��][��Dƹ�u�Ɲ�@�Z�o�o錬L�|1��F�\�dTM\�c5p���e�"e�Pc��3y3�b<ɋ{͘��?���5�}�ILؾ�n ���U���ݳn� ��U�r֫�S�R�t�~�1���}v��%�;b�T�k�+3��@�a��`���"�����m ��b�c�.����Qܳ�F}+c���3����1L+)�f覶��	��R�p��U��z�i�.�;\9F�lY6���]�_����=Gf�]Yԝ��uk%.�*�d���t�=�е�$̩[Ĕ��z����~���8"�Â�v������8!3�s��2�(o*�F>nV$�l[��op*�ǈ)8m'�lU�ŷ��u�WC����o]h�N� j��9���8����kkd&[����O�&����\Lc���Wtx1���qܜ�¥vs:��+b*��30���pQ2�(zU�elo�n�.���g�ճ�n3��'nSo���Ϋ�3p ���'�e���Y���A��Qw2��̥E�]��f�kanw:5�'1%b��p ���U����|n�Ȼo7�5�Րs
"y�x�H�p�7����*Wg3�@���('�S���h�̑3��A�
>�|�HZO�.�{���i`�v�td�gU��T�pA��,.�Al$Mn�����e�����Z{�SaI�1R�Y���(�S���Z=j�)�^��n�<ї;��>����+�٧.��ͽ��h�%�]�QF���=LU�t����A�V.`7\띢��ر�܂�Y]���Ռ
���;� ��n�*��lƷNޫ��۵,$�S���|ײ,*\�Y�m{u��N붞�h���h�Q֘4���aY@���уnW�]����Ei7�m����f�b�fk�ҏ(�+5�0�9+��K<"�pݳ�a��C�3���Ҵ��,���k���z�~O��kt[����<����S�4	�Qښ�4۵�m����z���/�`bp.���.�θr=��;�)EX�8����}��+r�1�N5�})��8 ����H���!U�E\I����D�s �}��Y8��J��{��8L��Ǯ��p�e�fP�/l?��g>V�7n�H ��Tk{��6ڵ��2Rïu�9�3~������!�e�v�Ȼ`��&C�6��H�O8��������t�lvd���|q���Z��ƭ���,�ț��=��v(Pp��A��#w;�$�#��=��B�<)Jl���xԮ�g����� �����^ֽ��^��r�j�WJ���K���W��x�؏��=�h���]��}�Pqp�'.SZ��+�|��E�����5�u���c�2�u\1��Ǳ�����;\���1�p�.�WtA���)�WkgĠL�F07�AR@[k4D�G�m�&��[ {���h�z���;-�7�z�R�	��Kk�q�0�Bm�7���q�`}� �D㿏����>���|��Wf��p>�g �o��n�	�z���՝UU�l�ܭ1�� Ǚ;� �.�eʤ\���o��h3g�����W=������p��C����]�e��}���:��ّ�o�� �63�5���c�2QuZ1��&���7�ԫa��������g}�&]�;�#w�vk����+�:���Ӂ����%\՛Ӎ��pAV�U��ݴ�v�3~Ϟy�?u���]����˛����!� S��\��YmC[af���Ã���:���e�~�]��A�p�29�f1��]��y��_�u�:q���h�c�p���;��;��z߬L\�虗��1����V�9�u���s������L[ ��Û��r����������:�IÃR����<=�Wg��%�����m�o{�U�� �>�x�(v�{N�WH�=���N��/H�e��ӻ����9�g?x"jγ�܅sVo���A~r�cˊ;���wu<��2�gMyZ=�9�-��L�e������`�]�u���1�?5B��{��	�g!���]�zu�v�G;�J;���t���gݳa��y��s��*r�t�@N��f�L[ �]�ۋFw�҅��eI�G�1���`'�ֲ�C�uE\ܦ�29��Ϸ3�I֧���I��9���A���r����]��݃Gvkk>��W5f���>��6Gi�g�<y�M.�P�_/�x�C�!U�!&��9�cm��t ����oK:�c��Q}��y�����ðo]�{xRO�ɡH��Ug���j�?eH�B[?���<.�R�:������|���&o�*����̸GwAwG���7A�>���鎭`�A�p/g�����ݚ����U[^�7A�g"^ipD�ƛhy�Gw�ee��e��'���I��At�̸�٫	���xvs��X{�Dq�'�ХY�.rKP��ۡ	$�ڧ�W��Pc��x���1�p���!��çD.p�!�w7;�TZ�/\�\����E�E+�Fj�.��O
��_����v�C��g�h�WV@7C&Ѻ�Fd��a�T�E�0�t���h�?Og޽����9�g���q��ús'U�3p#_��q؏���]���]����>W�3����	�q�8wa�;��U[Z: ��U���Y��:���dvt�����y�3k�lp�oM(P�*�3˷Z�/s�uowwv���2��_s�C͔�j��
���ŇT6�G��p�U����QsK��ߟW#�i�<��d5$U�OvP6��ˑ]�'�4h�M�u?cE�{�tL<���.�'��x��c&�[�<2���']�dȩdB��[S�6֢B��]�C�0����ћ-���꽨�t��{Vd꼭�+Z�wK6�מ�zyI�-��0�m\R�����:�Z㆘�b8�1�ʩ��i��m-�GSXM*㶍ҕ�,k�pْ�(�az͸�T���ˋq�m����&��W;��!��s���-�:��.�B�K%��:�ɠ�ܲ�!s�i*	�\\����oX���X�;�;v��7"�cp5��\�Qƅ��p��!�����Cm6��4ً�5�H�����Mq���������-�y�H�����fNn�j5[�@�3�m��A���WB�?�%������m��0�cs=;u��hÜ9��9<�I�����kwo��o?�x�PzhƲْ!7���T6�Gq��p�]��p��ԓ5ÿ��=�-d�~��w'��G��Ecak���{Yq�����.�����H~��3cGFz��7톷|�5[�e�9��Z�v�������Z�1��u��ݰm�wwxuu�F�vtҶcy�w�}ʵl��醫a�)ə���n�3�,tL��$��cv��+���hTw,%��GD4h����#DU�<k�����uÆrmӫ�!�T]��3��滍SA_8���lݸ��d�����H�kx����>�L��1�;lU�T�<�bq�O��o-j /�K�E��� ��e�Zs�]F�����8ˤs�@~���q�u��ɤ���^X?m���g7�ݿ���ü(�95ݲ^��b-��	E���a�m�qv޻oa2#0OV�ȸ�ո�������_6��ϐ�T]��t����Z1��uYmX��@�ZIH~k��������Rh}Ea����p|��av�wjj^��""B�`p���v5��[���tC�3�n��V۩�td]`���^!��M��:�o]�N�f9�6xn,p��=�[��;8e���L�8�k���U���Y��U�iQ�ݼ�����n�Ȃ�E�Z鼫��fO��?_M.�<��k�v�]�ݎ�j$?�5ltC��K�R[�+刁��ۏ	���R<̛� ���X��X��6��զ����
��5���o��^��W}�ʽ��l��Ⱦ��[H~��RI3�t?,}d#uհ��c����w8W;�њx�t=e)r��'oݦC_I������/'u�fZwWc�˨�@t�W=�x]�pFD�#b�@m"��rM��G\����vw�Fs�vJ, /<�:��f���̛tMీ��	���2���^��/� ��;��X��{�q�"�]�ت'��4���),���Ls��Q�X�\�=���m�f�L[_i��U���G=��x]ۿ,�%yc8s�c�˨�C�W=�z퀻�H�n��׆`6v�|�nq�H����W��Xs�[�?�j%��Vm&���.�r��15*�yF/���K��\�n��f���O& ��$fUCZnU�>�N��%�շu�7߽RII���Ϝ>H�G>l���W*�p��+awovF����,��д,�v4��A���'[���kn`s�G֗,Ы�j]s�/��ϛ���N�逻�4�c㺻]E�Z�Z|�6�����mwn�	��g�g9�6gu���L:G�<t:��jÜ[�wwDar��5�7�7�\��a��.������+��{�F�������,d�#��������]�����"ʢ���p.��a��9�uv<����M��T'��o�:6�l�I�!��O��?�����?�3��Ұ��:��jÜ�Э��]�w�{�R���mJ� �]\���4��3a{��5�TkQ���ݴ��U���fw�*��;���:���p�Ry1��'4Y�y�9�+JԐU2�:�(R��+*�,V����mgA�Ov��r�trhWaIna�l!��H���j�	k��h��0j��3���Wi���O!��n.�ab�Z�n�"�o��j�=��u�o�c���[��q����u�<�q*O`��S�vj�V�\2dnQ��b��$;�-�%��ެ���<��*wޡ.�WG]�v��[��ϱd�ջ�y�i���s|�����+�w��~r ���+�R٭����gD�E��q]��R�7\.�yu����V�W	�o�S�����Y���Q�)w	d��q��l�\��5fP"�+�m�;��)�h���m�PҌ���D�]�/��\yLi�`�f�׻��7�&˕A5c:�h�w(���4�*�t|D���|��A�AQfWlrޘo����̝۵��LeQ�-���oj�ՋZ�k�����;Hc̓����}��܉z�}x~"mvڛ�0�α�X�>>�|�Y�m5m���f���j��L�}�(ۼ�Mf��YVjL���B���CT�N�t.��c�j�ñ#<�̧.:Pv��y	y��]�-�K��o����WS�/9�Z�v+�w[Դf6�!ݳ�[�l+�GM(me��'S�Z�:�1k�[`lu����Ӂg`��}{�܂�X;9K0<��o9���7��v���Mڽ���#����ު]�i[��j��,l� �|���4���A��H�Ͱ?�<��R[(th��'J�+���>v�r<�K�O��%�b�T^���r���g�D�����"�!\���ȣ\/���"��)<�4�Jf�	$�.G��y�WEȯ%W4JT��OR�{\���)?�NǮ%g�xEVJ�����U<B)��Ģ�Q//(������<�*���(d��hʈ��<��]��Q=I��#W(�Ф��+��߮?b|�eM\����ʊ>��!����|��yx�,������zzRn�&�+�l���Й�&�ʽ��K�nD	�x�/��W���y]uɣ�ү�|��U���U���"��ȦxPˣfE�^}CߙS��e{�J;'baQm�2�-H�"����9T^k����_�6W߼~�6�,M��!w8OnyU5��9�!V+�n���l�Rⶺ�V�ۖX�Q*�f[t�HkKt%����il�����5N�t�X�)��j�ܚ��ٯ ��l�x���	B��Z�E$�Ϊ�jx�M�K�l�ؚ��	���e�.�� 3�vC�"�˝7�e�̪�/��h��@LQ��LA�LJA�;#�C0;���Q��;.�'�m��-�m�.�U��g�ӡ�Ғ�Rj�4I������o�kƽ��P��i���2��y��3�&]%�SMxݧ.�ƇS��.Î��&��]��"��wpjS�UӮ���g\�=l�8xr��n��q��\��V.Ŏ�I�۝)��hg*��=�Dz�J$�+h3R;]M�l.�/	�YzQ�p��q��m������J���3<�'
��sk����f���u�=\����o����GkVW��8yW�[��ӗti%.���{p <n��D�q����ܗu���X�9�F�[��!�X��;;��Uh��/Y�7+�^��B�c[��m�nH��x��J;Ǥ,qX͋WnC{<F��/Clj�Q�>ヵ��[It�܊Ŕ�^۫��@����C�YU��g�$��5��mn�c�h�[۶֖�.Mפݰ�n��0�ݕ;F��Y�+q��I�v���������kXh��yG9�Cv֋�8T:�z]��m���ˤ&�����Q kx흫�7F^�XHar��6��*㌼9�i{Y%�4�&�.�µ�ʚ�W;$�u��<اg�0U)-���s����,��:;q��BX���wrqG�1�q�YfA��Chkjm�h7g%/hc!E�,ͮx�:�n׆jnv^�cB�ے�q�W�j4I�L��s�D�M,iUke�� a5w;�j�ۭ�HP�`ܬ��+�U�ǒ��\��$m��O]���mZ�q��
���+��t�;J�p�q�6�p�W)s���l��N,u��^mu4�n[�ƶ�n��L �VnKڐ�Ӯ@��j�O\��x�3�qxwFz�n�p�T���GB�
�v�E�y��e6�1�rm Vlq��^���+���7���pb�.�7p[c���#e��g9.� uם�X�n�,�x�lj�bx3%���n�9���P��K%�8ȃ���L���]3u֖Xb�k8-���O���6�9�����x�kb��kw}W���8�X�[J�k�q�'���m���R%]Ф�J�ݨ�C�o�$�H�_��ޢ�,kR���3g!��U7����]�ܷ��ja�]��k���8�Ǌ��M���eHa!bOl�c�=��ꮆ�?I�	������N�1�Y/`��Z�������_I%ԑUHD��NW���l�ɐ&u�k]�;�����Z5�V{���5�? 8�u=��˚�wov޻(l���n�Q�Z�g(��{Wc�˨�G]7�sݰb��E�9����L�\s)4x˜�Ku�ͦ�{�f�:ӝ��n�V���یmwn=vû��#��=�x�a�J(�?;��m����wpf�IuD)�5T�aV4�%��1=RX0�1�]c�'v�-�5T��z+��V9�/ 7KM�;�J�#n:;���¾�h���0����٠RL�j5�;�\�ǵ*�pm୅ݻ�#�� oG��u���]ݴܮ�/�D���f<
ʋ�{�t�]sݰl.��A�C���vv�T��=��.�[v�4$s�z"��+��q�U(_�KÒ�|o熅�I�HjH�����2v�$0���Y��e�eʕg��&��H�BO���y�*W����	At��7u�ݬ{bB�����r�ۖ�M[:�ilZ!�25�]�v�-GFq�]����?���v�ҩO��T����8je�0}�J��X���,~y�W�Z��*��G�z���W�yO��"�Ԕ���~��c/[����\���n��x�	�C�nfV�Ӧ=qu��`Gp���xQj|�P��̦�N.��R��a���$�0�|��t+��nl�U8z0���k�*��fί���l.��h�3��숦ʋ��{�'&���<��l�L=��]ۊ��k��o����r0ͳ��1��x��\<����𻼧�{��U�HI�}�-u��zQJԢi�O��<��wOM�xCū��9�Uu�#٪l�*!��~N�՝>�avS6�s�vu��eʕg�ZZ����u����n�p.�]���(e�o�2lW�|�\'F�����zl��G@{aQ�Rx�V����=쯺�C$_I(>v�2G<�lY�٫q<\)wW�Z�o���C�T�T��W��A���n��ͬ����Q����ϙ�*U��.�ˉ��?o��uڠ:b��CiY� �f�떾PiU0!���ǫ�o��7�Ⲟ�ׇ:W �WC7���é�_�ap��\�n������Ib���eW(���s��OG��{%鲢��u�v�R{uz�����!XC)E�j����Z�we�r���:�eB[@Fkc\T��)��������A�wr.�wY��x��,�x��\Գ������_ +����A*I���˪�^-ใs��k�vq�Y�J����k��Suò-i<��C�|�]�ww{aI�>���p��ŉk絙/X�ɣɚ��)�H�*kէZk\��k���o,�e+5�W�Z�u{�_Ay����|�?}!�H��������=u�q��LE�����"����߾����o���O]Q*���֚�*�.Ӿ~��%���ŌC��b� �
8��Ra�ũ�7k7n 2���K���_vѷ�z���*���;(v⫡wK�Wa�e+�M�\faB��(�+ 9����Og�%�^!���h���݌m;�l�ϧ��kg\ж��c��>ݴ�����ݮ'v#���-���0�2F�MÝ�Y��ӽ������)��޸��͇J�V�A́Lºh�*�CJ9���4��8WcqY7�C�Gwk97sv���(��6���e�1��D��n;Wj����|��\��w$���vuR7EA\\f�j�*�#�X.�&�XCÇw�7���n0�awo�'4cv�o���K�G������{}+�O��?Hn��v�zad6�FM&|�w0��e9����-xWyտ��]��c��5�]4ǽQ�8��RE�A�'���{f�9���-��m�eڅg��m�wr�����v&�Gn�}�bsW@��g0v�\'8���zˈ�GC�*�j/D
�T�Ս�-��Mn��M����^�g��>���w�{Ŗ@eХ��z��9�	3H';X�6�qp�>�=n��Ml=�V8�G>q��Z�,����An���T��)Hj�$<����
�K.����=-{K������u�.亩"Kޗf�܅�M�"������x��ּ��h
^C����7�U��c�m+�|9Z��i�;U�{B+��I�ݘ"�t���n�f���9�h��s��{%�."����qw\ũ�A���yWzK�*������{�/.���مpuoV޻k�]��'7%]u���s�+�f=1�љ\Ζ\��=ޫ`��㍾T5������X�퀻���7;��ｏl��+���}짬�����,����+s*Ǘ��P�(|	�vJH�ݸc3�F���9�k������s���#]veck�wD&�.��7n7�6U����7{ųp��(��}n;v61gPR�;�ww ]����_�n���A��i�Xs9َ~�����^���8k�HݒݯJ.�5�iC��]��aw|';��gC�}~�E��P�N]~t�I�{I~�'%�v���a��wRz4ݺ�f�D�hZ�Zk�|z��{B�6gg>�#�oW�M�܎c��Q�vξ�_K�+}U�~��I�7���-n��x�ܛ����m�fY{�.�
������	�P�Ħ֊,=Y�R>�U$R�v��
������%;��V�B{��p�[R`.����m؜�9J�;�|��ךJ�z�/q����v�!�c/%������hs�AF��퀻�\'����ՕV3|Ʋ��ɵN����]����o+nv�[ �5[Z�u�g1[{�.�
���
�[�=��n�^<��m����~pԑHj�;����T[K����^���{ڵH?~�հ�2��(j��f�48��@��wkD��ܺr���ܭ�+5�C�1y;�{Y�)^gW��E�ƙeSt�8 �qc)��N(�F�Ǫ�I��0ɵ����'��_��4��|��
�=-Y��C��I2�C�K|��*O5���v�:�dח�-VO���9n�	0�����`y<5-����~�,Ѷ$ɶ�W2��`\N�������7Q�����ȫH�l�(���KR�Oߔ���M����t�=���oD�8���M�I��M�q������ĉ�;jc����=���]9/�OalC ���{P����da�Ƥ�]���I�I����S��L1��.��:�S���Z��!�H�/k�=�!�e������]�my�����x����U���ٱ;=���^w{��ݽ�]�	;����(`��]/�Oah�o*�l��i�vy>T�o��r/�Ň��[�u�mXZ��V�n��x9.d���v�ov�9k
�J}�N��醉���w[faкg�(iY�8bҪL��16e5j�:�!�
�9�ׇ'K����č�q�]X�z�ۆ.c�L�[k,�M� �Z�=�8����z�sv܆��7OnOI�s��]2vv�Gi�u#j�q����28+�UY��cv�Jv::�6+�ռE�yU�v��Rz�6�K2�T���s+�PV�۩�48q�WM�f�n�eڻT����{�����
Ț�������;VZK)F�֨�օ̹L7߿y&�w>����zݘg�ʰ_>�ۏ�F։�u�Y�v��{www뾸s��5��:��t	���0L�/��z��z�����v�"���
��h�����wq�w}23����E8�Av���ʧ�H�*���z�J���L�_2��7��ҹ����ɘݗn���_>��U=�'�}��_��޿Ys��HjH��,���m1-��7=�y�p�8?e~��$_I꯹���#�}ϟ�g���b�X�;.���\-	�6+i���2r�ro]����`��soeK�j�����P���Ww/��*�5��#��}�LjL4���l�h��زz�7����<5'Y��}@�YxK�sܕ�a�hSF&o)õ�8��d��٩[�3�f����U�WOiW��K9�0Y�8�[�%��}��Sݷ����8�N^E൮)7�a�]�����m�����i����o:�d�T���$Rn��ΜZkLݿ�FV�Ӽ�rTU4V���uk��mwy��K��ݽ٪��:�|4e�~G��C�go/KK��[s�\*S�U��aw|�u޶�v3%l�y=M�/��VQ��7��316k�cSq�B�2��a.���dm�]q�ß|z~�?~�d��׭�}��֋�ӫ([T�7frw/�܏8���qv�"���m�������h�;���3���vd�)�h��� ��]����qi9����z����}Ë�yGMK���yB�.�՘1�����,L�߲��q��B�)�Hve��,�E�oh�P�Z�t�-l�W�v�

P�]�T����\�Bs��}]׋����L�u}7xsށ4Y�4\�ΔCc^���\@��"$���S��M��|�G��!�*C�Ȁ��0��ޣ����fޮ��͑��� o5YWL�W,������n�	�};Y��Mi{7�Z�
n5�B[��:��c�6}d�+���h�l�]=휝5S7FDF�csfwJ.�m	�a�x(��d��<�z.�ӹ�H�b�\D����Tp���+3P�]s����四�ďnd�F�>��%$/+N�\�����w�����9�6��5t���U![6���/jP؆n�]*��F��6Õ�`Ki�f?�o*G��dYٌz��G+0�n�J��:N3D���E�P��4�]��o�����nQaS���%iުa�ͪ�ܸe>��ۿhg�ծ׻��I��FC���t3�Z�SԞV���.d�k7G�7�޶(ݻӍ�h����	k;,ֻ�v�%�n7׮�}��!o^U�,�59ft���`Mɑv�%���m�`�e"�d�g�7�_�����dP8#o^�^�箟^m�{��Ǜ�i�aj��,��x��ބW� �@��5%B�Z���:GV��eK6�v�qǴ�o#y���×l��\�[�Ƙ�Yy��v:ܾwDP8,��;[���M��Bܲ;��EL��˺�e����e��y�O~�uy/�����%�Py{Y3��rs��T�ߞ�Ƚ>{=��D}Qʂ�<�W0�p�
5Џ�^|J�ky�9���7'�d��$G���N�Z�I=��G�nًlm�0��R�(�����&�M�ܑy�G�;���#��{!/*.��$��9)�m�_��xr�\,��ڹE�0�T��(�.F��nu���UAg�)�[���DQ'&�W�U5k���lA4�̐���M�/���_���'��Ï��66�UJB��I�@��fD�<��hOĞ"��<
�y��X�zϚNn�yS�O����)<��ۡ	e����R�ՈL7����ѿ^�`t��^�W;��,���i3�e�U��ny��؁6�	���}�=�����ٟ��E�o5���{cKq2	Q�7��u\�;p�G�|z2-��Q��aɭ�jEy}��ϗ��yx�ظQ��z��]�9hU��e�8
5t+�=�Ii{�輽[��毩��H�.��C�F�a�N�l�v�����)�ueu7��M�KA©�e��$�$�&�ۧ&j9��@nÎ�/{y�'*��,����l.��;��ޒ���450>,�-�c����vgζ��lt'E����]v�ő�v���x!�����n��������ˇx�;�oѡp�n�>���d�@���v[4)����㱭OR��L�OͲ��VP7S|�=6�&wL7	� yaB�՘�I%�RIgwe������`�)�o��c�wb�m>�����v�lݿl���/��������lm��|�x�r��4.��>4��͓Q|/��q��Cl�;4kD�i��v��Kےk���ݳ2��5fn;�(��=�F����忲�ٳ'����° �2q��!�+n�
�w^{`.��w֖�-n���_���$�ά&�����L.��.���f+�W[ �5�ii{�	��{n�#�$�r'�u�A�y��ôz!��8I�齛����օ�7w�)�T��^�xl�yr�!O��.�R����\1�"s�u.׏������u������л�8�mw�K���b�u���`.���]�讦yE��m �;;,�_�ogN���?�~�*�.�	����bv�2[�����7w�*�.�^BO�ὁk�6���]�;�:����!�J�y,��{P�^-��Q�����?>������m�l��|��4Ul�I��a8̎�m�'��r�A9!���2r��y'sN]�q�t�w����K�+in�'*��m5-�<3�F����[���� v�ݬ�lH���ŉ�ޥ6��uQcN%��d���!E��[����2tQÞ��N��5v
i�c��ls��շ�1U��d,ҹ��˫3�Gv'����;Jq�`�Xa�y�e#�QN�#�.���=�v[�v�S�j׫���m���5_�㯎�1�u��q��U�@g�.v1�1�s��Z�;ACFo�~A�~�ߎ��,�X
��L�u���b���rL�9�U�q�����l��g�O���^��d���%�m��<nhpc3q��SOϵH~�I/=[J��{ާ�)ӛ�����ǜ��Y
ߞ�/�]��94��	g��c\$�ww>�w�{;��B]�Yǎw_����S��K�H�3��o��]AȾ�{�?k]���jvKvv"�s ���ٮ�{e7ޕ��R��$U!��(�k��X��
��Y��8�v+!K詗�l=w	�_'Eh�A�^P��1L��N������T��W�\��{�6��j�lυ-�;��hl~W�cx]ہv�cVv���y�֜���{�c���S��o7p�@��!�-Գ�>w<,�V�R�x՞�{��eO���u|�eBҼNCɂ{�r���J��gx�Ø�C*]�4S���&dE�w��s���c:Y�v�6{��&���F�F��D���v�m뻑��wh5�u_l�F]؜�/���x+�lݸ׉�c���_P�S�Z`�_�l
���ئj�֜��и^SB�z���������CR�*�u��έ����.�x����.�d�[?T�$_I[��K;��e�23���f���g�LrI`�����\�A��j�&�m� S#�ɄM.ĺ����o~>ܻ�]ۀ��7�tc�]	ɹzy�����+��{*CRE!��w�2߭]��{�����*�v)����c�h]�^S�v�j
q�,��=tk�gÓz����-��-tdw���,�9���EX����S5�(��˼ޛM����m,z���|f׏�P�v�}�������ɏ����!ǉwwT���~Y�֚��v��D�8MLrY�R�V�Ww;�p[�;���NM����z�6�Op�-~�n�"���R"W`.�;�1��.��i��+����mv�M��o��������ċ��W[��MN�8v���Wl;Q�E���h�[����=���m��Q��Q.��\9��Ɵ.�kxB9��\5W8�k����jFJ�8ƞ�t��������Brm��E�����]�̯{bc�}	7�L.���v K�VF�w���4�pە����師2I3�۞���r����ʥ�Ҽ���S0��\9�����J�&�0nՓq-oO0?��䲺Ě�Q�I��"ܯM�������q{}tY� ^��T��uP�4=8з�"�Ȇ��*7�(�S.֠F�s����awn �o]ܲ�~܅fU��k��g���ύYt'&�tD0�W�v޻{��ڞtʷ��	j�d���U�xn��m�O���N�v.p÷\c-�3�c�~�`+n�n��n���y�R猳�R�ғw.���	5ݽ�]�e��M��~�m�-���/;����͞�&Xyi�Y���G߹�/δ�W���Hd?I7ou���T�Us'o�dce�	Qm=����C!�rs��g?	�g�;6��I�6�gf���l��<e��忚�o�p_k�J�I�!��ԑI���n������|�ۖ���B��U^�jH��t\W����a:]-g�`dC�VD��P�ۙӪ�Pp��Ã�$�wH�v�wm	{��@�Ў������;7�E<�w���v�V�nq��jNP ]�>1��i�<�6K��#�K���#Z���n~�5��A���g�.��ev7e�ѺKjJu�ѐ������Y��W��R6��͛,�Q�m]��"��z]GY�z�uX�y���H�K+�f����9��aᙬ�ܻ�͹v�:k-��М,Sm��rk\�tn�%]lsۊ�����8��]i4w��~;��x:f50�);*�@���<�z�S��c��� �p��`����z{��.o]�ݿ���v;]Е/�n5i�,�K���2E�Hc��yuz��t��Ս㔛w�n�O:���T �y$��bx'����3sհ�[�{���q���ީa���;Zx��Y�a�U��"\8��]��]��xoK6�Am��g�r`/�]����_{]ȕ/�<7�pE��bޕc�W��u$_Hd?I	�{����u�a�&{m�um���n�OZ���\ �p��o]��c�����QfdN ��lS�� �ۀ�9؊:�ӳ0vm�ډ$�q�h���5�"�.�2~�nOs��&�Y��-7��l{�P�i�{��cwp.�W	�Y�ʰ�zK���hCM,���;��ʖo%Yu�,��0?tj���Şg+��{�F����tg
a�L7 ����]��}�l\�X�gq}�9w"T\���W�.�PԺ&"*��l�)���V��T��f�آ�]��gx��r�?o����N��5!�I���#��zBu�@�m��o=�l}�n[s��&³�"X6̈�n��3�s�������]��q�'U!�ﱊ��/��I��s�Y��g쫐�R�{��vr���'�ݞy��R�z��f٥��-6:��e<q���C�*�6�� �j����f/ު�;�I�/[��3�֩�5`M���'�.�m���v �$�&&~���˻�9�Y�f3j؛���0���D�����O<O`�`�_g?��]�wQs�e�aa��g��A���6W�i�y�u:������v��Z�Wقt �Yc�[�XzL�Z߭��> �H�y}N�
�9�$ol�{z�L���^�gg�R�R��g�v����8�a�V����*j��Xz��U�o�`������퇮��v�w���:M�]Y���Z�ˢnr�ØV{��D� �%>��ŭ���$9.� ��JL�i�V-�mi&t���Q���Ѱ�Ѡظ��k`���`.���k��͋F*�*��̜Y+�ż�q��ww#�rxl�Ξv��Z�v��k�)j��Xxb��k���kqu:-sƷ�����l.�kzw�ù;��CN:�J�0D��g��%�@{�q�l̙��wm��܀�}�߳X��cڸb��K����mC�9m�a ۟e�؞�W�cr�J@�S/@�N�]������;S��v��g��SS���3�~�o��~��^\
��Q�]������o]���v޻���=���w2b��1���^uS]����.�z�v�]�@�i��A��}a�L���3ZA�}%E�qnِ���]u`Ü��0�-�:������~H�m\��k�ܵ�_br���2��	u����55濮� ��$�pjw�Z�tv4�2#*�Y�R�c׼1L	P����?)闫�bS⮷�N�USMT��H�N�X���}����;a���?I���$R��?^Y`�,,��گO*�#�lr;z�8��<9�g�D�[6|�V��UNI�?}�?#�YYX���&�V`W1&�����Z�����~�����#��	I	*�� ���/�3��H!$�W�P�lkl��  1��I�BI1�I&=1$%C@$��	&4$$�$ ��H����B�b�B@��$�cIL�BT0�Hc@���BLi I�j�!&4I�Hc@���BLiI�$�c	1��)D�c@���BLb��$�c���@�Bc��N�HcILb�HcB �B��BLb@�$�c@���T0��$�$	1�BLh�Bc	1�BLb@�I�EBc@��c@$��x���{a�g���H͂BI!1���4��j����_Y����3������a�.���ꨳ�:�+������~���Q��G�Ԓ�^��k����Z����u!!$$�����?��}V|��h�0�C�_X�p�������%�����@����?xb����'��޾�K��!I0�4$$�0��M����@� B_p4� �$Є4����bM ����:��~P�!$�$6	��ϡ���M��~���>l����������W�K¿y�xQ<KK�>���6p4|��$!$$�i��%����Xc@��^�I	/����};=(HBHI}��$$��	������i
!���_�U�|���A�Mz�6�/������|��>��K�>ϴHBHIiX}eP���˳�>�����������}����	I	/������$����Q6X�/�!�	�`�����5b�����ؐ����~��m�q}�оjХ���x|p_B��������߈BBJ��x_�F��������e5����_�=� ?�s2}p!���                                     } N8(��(�P��TJ�	P (*��J
*�E($RP��(
P$UU %T� P���$�*��R
A��R�R��A�*�J$�!D�U ���JP�$�*�UR���*T�PD�T�� 
5I*EP�E(����� n�� ��҃��=��S�-lq�U�S�U�s���{��z���pw�M\�=�&��/xU^�{�=��[��5J�@  � �`  |����� ���+� � M�� n` x� S�g!AAQ&���W� �{�^�י�U:��z�֙��z���J�8*�(�QE|   {�T��T�UHD*�}��T��v��*����Ѧ���{f��Wm�<I[��)�����]��Z��Rj��+'�)J�ԪU�w^�R��ü�$�HC�   wWK�{ԡ���^䔅�*����֮�W��{��
�۽��3C{��tU{g�K�R��k����˪e�w�=��b�*QT�   ��E
�AQT��R�黎=���S[��4)WvZų��/Y���$���Swux�j{�=Kҝ�����yڕJq�T����5y�]����KڥU 
���  7+�w ��J�"�
92 ݀l�� k9+ f΀7Xrv � ��
�   y�*�J�UAT�"�| �� ��  :�T�X��@���� �UJ\#��((*�   }������r)N H��Ä�#� NB� c������@� �� �>��*�%E���$	UJE| ���� i�8�8�� V�!Ƞ[� ��2 ڠ��}�8�}��	)DJ$��@ (�S��wX 8΂�� wwPv�� �d ��J �`�����h2RU#@24Ѧ�S�1%%T= 2�z5R�� ѐ4�*@��   J~�%Rz�`4�MD�B��� d�O�������S����$�!�Ͼ?�(�(92��~2��4�M�� ������� ���	HH@I?�O��@I	HHg�U]n���k���_�Lt���:9��^ܐzt�l�%�[�5b�"�y�M��z
�
��x��6��\��8�mYhꝙӱ��j���:w,���B��2%�81���m.,ߴ�����ӁƱ�$�f2�w�*'�������o[ҕ^�Z ��%3xww9���ӧ8���˕3�v-6�A��`K/l7�b;;5��MZ�k�i��!�ԣ{:�N�7g:�Ś��3���g��Y��@��f7���@7����%]���T�X���v��mv��o6��x�p9ӡ]�q���V0��Ń��!��v�
Ր����[-0b�fvU1�ލߖ�w��h�<rrL{���R�Q�S�ӲT�$9זu�(7�,�ou�{p�U���^�*���z䰽�׶[�U�z񫆮κ9�@�Xs�gNE�`Z�0r�B4���v��ɼ�v��o�^K��sXd"'���x�em��Z1�BG*�ƁY��7����[WL���fo}�xgM]�XgA]�Cs�t�m�������ۮN�+��xM�N0(n�Xc��n�<5l��9Q����C);�X]���v�qyNNF�<u*+i漹����d�ߌe>�D�U�uWnn��l`Tq.�+��OA<��`��z�,��+�X}ȘO6���pv�໴���>��`f��wt��/L�&��G>�x1�Z;�ܮ:��v��A�1�wU��@��f��~�7ol!�,�ӹ�$�چ��b;ȹ��'oA]�.����(�1R��غ�D��ɲ�����f�q]$T9��{v��ǌ�5v^s�&�Ƈ��Ҏ�5&&�.C�[���6n��V���bxPz7�K���Z��k���c@��a��3�s���^6�?w�d�� �;�*5-A�{sL��y%�e���vW1#�E�yзг�T���h�v�����ܚ\b�Y�!# �+y�.{t�A~�'�r�pb�7-=��3�=�77��c-q;�([Ǚ����ٳ�B��N��vUWE������`;���r�P�Tz��0'ٷ�rِ��4����*�#邙�l������j*\ܳ�j姧�u���;'{w�	�7����Kv�r�����A��J堜��L�= ����g���im9��&Au����J��_<1p{G%�M9w8y��F�2H7nY�9׸���E޼xC�ĵ�i=8��X�����cl��nv=�K�;c�'oL��z�������;�ua����z,�#�jw�n,7���р���^m�2i/�<{�Lic�f� ww:%/�[m=6������B2��%3>4[V����'W�G�e��4�ݥ�3��*�*�4΋��Q3����R)�N���L�Q�8��j#�:JGd�9@΅�G��7Y1@GWe��1��[�:������͌!5$L<\{;yT8���e�7�̈́p��i��~�Q�od!\z:�X�ޤ�7�e�K�a�FMYFC!;0�a6p���-7w�T��XKmew�+I�YgL�����ɻ�;�����x�	m��߻8a��^����:�M=���gۚ�8�
���PC��8tsH��JV�|�r�O��W�r]w�ň\Ol��Z+H��E��&�!rP9���ٸ�@�`/8L��X���뫴��VS���8mV#zF�A����3��d-~}��0sG�����+�]�D�e�Z���'l�3K��H	�.SJ8
皻%��vԃ��}��S;&nw<ٌ☺$�k�ӱkx]|om�a��k;$S������K���;��C��QF���9��Žޑ��C�)�j\�C2PDx��_=�h�ۜ����3[��l&� �{����&w��Q`�n�R\����W4oH����u��>�p`-lLuo�1lW�wDnZwy|NQj��f���ˋru��z���s�.�XHmjH��t����:T�Wܗt4u�W�J8\q�Z"��cϽ�X�i�f��L�Hp�$�2�̔Yf����̌B���N
Q�$VZ�SY�X�֯W�N�:����<��K�쑼�0lj��7�f�n�X۫J��ΊĞ!rHz�c*��InZ�uV��Q�z�D��dĞ�58s�h��w��F�G ��}�*;�t��v�D6��q:s��2��q)�l�(г�вP�����ɋ.��)�}r@
ִ�zh��s�.
��vq�w��v,��A�%��/$~`�I�;����. �	��S�t�Oj�[�od|��Jq]�${(x���9RU#�GB�A�.����&b��IԏQ�逎���Q�f������l�n�KC���&�Y�k�(���KUl��wLo+;Fbʢ �e�L��9L��N��ӛ9	�Qb��[ܻ��-����^��ar����ݜ��'y��_�#��Z9��/jo��v��r�7-��q�׋B��u|B��@���wD�n�����=N�t�׷�[��t1��b���jٛ��[2�4C�N�p&>�@�!��w��R����U��v�n�V�����"8��N�;ܧ�0ͬ�øV���k��O�Βû��T��{.4��;�\ٚ��{�j�⊁87�x�o4���&U�h���2pAEӰ�Ά���;x.{�e�Kc��3��0��q��)�7H����/�&O��x؛C{o<��f��qD��%\Ӿ�W+�.=�%;p N�{tu��"rjә�J��0Y��5�1�{�:��'Y�^򸃄a��gn�p�v���rp*�BqO��B	 x�!�he\P��mI�7;�\�#�s[�'�Ԑ�Zn�2J7Frѱ�4��z�o��'��^,J�%_ P��fo,��=r=36�yejoF���@Z3]�D�r�<-F�l�K�ǖ�gd���j��ӥ���-]Qg^��7�.��^iس��<��i�i���N �-�vqgd�㱥�dv�9�H�5�����B�gj�z3�p��sJT�i��쳷[�'s�'�S�nȜ�w���!W�o)3bɣuȘ���n)a�6�������}9�_q8�ѳ�E^Q6�w
��8���2> ̓��E�i���yv�å|[�Ū@���Pd�짫�/4w��F��1X��wt]�D��I�f��TV	�O��]�ΌZXl��[����ƛ��μ�r��:N�rf��χC�)�3fY�x�|o�%�a�c�5n�J����g��]���Ѵ��Qr�!�Ɔ��oL��gzp�{F�؎�\n�֩vt�����>Q'YͲ���*o,�u�ae�}��'��gXTA��ww���k���WG,�5R<�/��s��s5(��v-�4ͳs�qW�����:�mkK�Ð�z���	���,�Ê��9�|�Ԓ�Z���c�C����-ÜuA�e�|EMܔ�g\�n8v�C�� ��{��.���fU�J.aѓ�q�i�xvU��ѕ �[н;2������=�E����[�v���z�	Nu���D:�+ �x齊���W%X�IyRr��a)���8�����T�ı�d�$���:��)J���{AS�K��0�pќMX��tZ@kWvjÜ��%����Oc��ڛۼĞۜO]9�$���*[��ե�E��u!QVi:��A��g5>z�Ut�)Wj��Y%A����J��싐Y�7O^�p�<+�˵���4�[��g^�E:z��ɛ�c����3_p�t��^h��UR��e�������^�۲�()�z{9���-��f���ם�/N�>!�m��8[�6W������<�F��T[��
8 ��"Y����o\��a=� 6�wQɥ���{{�X���^#.��f�ۋ;���}˓₤qXg-�32nG"�s��Ӛh����=}�t�'�-\!��3�ל��[��坽JS����M]�/����%5b�$���������7X�n3իuJ9e��M�ռ��7�����]�[M���Fv��3��x���և�B#8C"�]Mz�k�h���^�_p��%� ;6s�)��3��oq��<4��	�.�N<�3�s�4-.�N�i-��2��۸1�U�(�<�U���8w6��Rq�ř�p���;C��>��N{u��T3{	;��8��@��c�=��7pE6�l��dȴ̀�ܩ:�#r<�A��.���û1s����1��aS��N�Z��Z�ːt�WU�ax'�M��b	�Id�s����-�p�`�v��,tzя8�'7~93V8M��J��-��Wh0H��6.���W��QZ���r8�����W.ŭR�m�n�a�.�9��I�� ��Ӹ��q��괧�꓉}V��
�hHAa�9u��v=��ȧ�G�wh=��Lf��;D�l�/&u��C��c�Y�(�F���6Z���N�[C�meo^ރ�F�:5����t�bieŵ�/Z�(.o���3���nhx�=�:��Y=k{�E9�$�A�����p�-7�x%�:�f�&y�ݚ� 5V��c)�M�������\����:>�:t�]ֆ3���v�|��Y���j��Q�ƅ�'w�;�n+$i��o��YӦsu�����b<�I�K{�2]�����G��8<QtmP\�su��d]�*ƃN��z��\۸�>[�K4���'7��=�a���o��ph�h`�{��%�"��e�8NzԦMTq:Ƈ�a�.0&�Y(`��P� ��l�-K@	vs����E���"�f&�� �ƒ4ë��a�H2Y��w'V�$]�w���3�N3�ǯ=����p��[r���5��7��Ҷ\���o@�|���U�C�<��`�c������"G9z�ݗ{����l���F� �5���AԹ�����Q9�5Ѽ0�4�y��o��ٔoسK1�{�=�1��Uo�:�iQ�U�4ݿRv�ʰq����v�Fh�2��ݭ��Pd�m��"w=�t[���nl�j�s��f�Z�9���JZx�r�ɮ��g�:�Xk9��pᛀrtD`w^n��j���%�0��0wf���ۀ������3ZM��v�I���Ixx#�_!wr9pB������[�E��^���T��]D��ez8n��u#���q��}��;v߅f�W{Y�����Fn��!�gc돮���guy{�í?���.8ES8gÏl�y�U�^*��rgKu�f�X���L���)F�ޣu���w]��G�E�Id ��������`-昵 )\J���Ah���7Y}#ܯhX4hC8hT*��쓗j�u֜ө���^ѵ=��u�V���Y!��U��-މ�9�rˤC�,��J�����b^�&&���c���uKS߫�<�ש��U��=lU=�P�B>����k�f��z�,q,-�ջ�-O�8.�F����0.�4"�Ǹ�9d�z7��6��N��uc�w;;����ھ*�����į>Ap����`�B��V���۵Ekᇭ�m���W�m}��q	����<���f�L���=�r�b4Nws��j���#� �b�+��_w �󝆖�C5�����v��)w��c�o23��&�L�,ANo"����wU�I#���p��U�)e���؎n��5�9�|3� ���we]0ю"n��>�>K_%j#
j�ؕ�����2���Y��1����V�����V���#۶�Zf�'T�3^nl�qr��lY�M�,
=pq��K�;;[�P˧� ���T�~�q8��J���3�α�ӑ �$_�vqt�K׽�K�-V�"�![{���J�9��Eծ���5=�0�ao-ĳ���ݸ�L���� �}���˧gtq��
�k���m���_uvZ�ۍ�5���Y�*���D6�f�l���D��"�e�˱�h�1L�`�jK�1X�ۑ��ޚ�>�f���N�`�oǾ�sN��u|�؏掵d�n.PY�m����bx�׽�ɗ�����J�GJ)�$���s�8��imCm}���T�7����\GZIviSq� f�Wy�����loHz#�wX3�dF�3za[�C4U9����Gu�)�N�f�o���p!��n�"7�-�S�z���
��J��uوM�sz���Ns.J�DkG��2���;��oGF�6��Y�* ���eXgX�_N���+�%�]�nG�
�v^���VJ'`�5��ǹ,m�m�4����,�Bh�A��%<P3��.w(���<'>1��C�uq��;٫
X�ޛ��k���ֈ(�$�6̗F�$��$w�iP����v���r����E�TZZ�]�g8��w�䶝s=��L���Kז��`:,@�6q�7a�v�gs�� c�����v��f��'n[ޠ��z��iGW��Z��*
+nX;��>�y����JuA�N��ܴ��aɼ�vt�ĵ�zy� 2m��D�L��+ŵ�p�>5ОHAd$	$$�P��WPU�U�WTwR� Y	B
I R(IBH)$�
@�Ba ��d�IH`I@XHE���E	"�B(RA@��$$	d�Y$
	����,@Y �@YA@� I"���E$(Ad���
I"�`
H,����H �	$Y��)$�Y$$�,��R �(�H
I!I�@)"�BE�$�  ��$�, 
IB
X 
H�,$�E �d����$U�u�tutwQutu@���)� �@PaE���@�HC�����  x{���2���lEFe����� �{�Kh�Zث陈����G\捅!
Y��t�d�pہ�̄�l�������>=�`�z��6�A� ��R�>��k�j�q��kxr�������Y��7Wi��ޯڵ&��y�oy���.���6�}՝Vü!�:��ˏ�rk�9��9��E�ͫ�#
K���jN6c��A�Y|@~|7ux�)�}�t� -����Ù�<x6k�NcM3���AqQ�˕�]��y{q�ۯ�����Z�,�֬��yQMM�=W{3XT3�L��������i��摇ؐ�W��	���+�0���Ԓ�3\��dF�
�c:HS����j��|�קF��_�wn���	7�B۱o�_t\l�|�:y@������{����a��ٯ�3��w؇���u蘝EDC��������P{�����ha��-�$y�L<h[	���Rn]�����8/%:[F�TK�8Sgm3�o�2��/DA5�ȻJ�MA�ň�Aj�yY�|��X2����g���i;�ܻH�r$U;�Y�j����T�l��.���^B� ��93�y��q�<9y��)�[�}��p�ؗ,Z��;����==�[}}�ѥ�Fd��������=���vIٮTOLʑ67��>�_y�����^����%��бCm��mK���F�cH*q1l��7��J$M��hS�:�єi��yQ�qw�p>=�Zz4w�X�轸`�P��w����g	G�x���g5���w���&6=ȸ����
.U`�_KpS�Vc��6p�����z�<�ᾙ���{ĵ������	�-k`�=x^���xK��r�Y�r��-,!�Ǧb Qx#��=89[ڻx��K���"ǝN��ԽC���h�ՒU�y5�L��;���JS�%��%�`����a]|��W���j�����@��p ��cY7}����Rvɧgkח��=��.ގ,$8����T���s�{�i�{z�=j�(�mj���j��Aq{������/��N�L7	��A������3���͠c"�E��ѻ��J�y���u�h@|gk��G��{7UFo,P6�nݳ�̜�Q֢6ĸ���n6��u\�3e�r�d`�Y�;2�K�i�����&/��D�J���s-��[����)F޽ټ۹\�M���ٖ�x`������d�zȟkx�������b�eˑ:]$�P)�]U��Ṉor�v�tf�� =�ѵ�i�xJ�h���|�wm��/|�R�dr��#xE!|h�$j�sm��lF8��eύ �j���U��c)�W��K`dR��=�T*�DOs�@�#�ȱ�}=w�ۆ��u}si�d�z���v�KNҢM��G6'cu��f�6b�!���e�p�
Y(�w��^w�yM@.���ؾ�n�[�qm��$��#r]9��	ݠf���չ[��_m�� �� -Ç�V�Ѱ�7=EX�x&Xː{M���ݽ�&k���4y�G�zn�c�Wٴw��p�|��'�����ip�k���T����k;L?s\�} g�<Jn�m�<�U��U��|I��il�Ҟy�9��B����_�`�&D�i�=Wr�5܉x5��3v�f��537��q���tO�η|t�B^�r�9b���8u��8�!�zA� a!DV�H{�3pnǣ��}��z���?!��6x���b���������2�N�����V0mYn����+̄��Dc��H�ةj�{���~�5)�÷Sf��d:��hi�1'u�x�=!����F���ۯ���7\����~�7��=�4��-+<��B��
����o��sb���z�9�c;Ճ8��r_c������Oyn�:z��c>�Z��h_?�E� ��{����v,ܣ�~��>������b���{z2�	�� ٞ��wt�38v5n	NEC��m��
$F"6�SmuX4�5UB,�X0y���J��-�˝���������~�m�����V��޻�7(���5�o\ߓ�ћnvT�| ���KW�)���:i�En3/nD��͖���WF7f"�Sˤ�<���7.XZs��{÷���E�ڽ""?j�Ѽ�<wh�ol�Ѻ&��s�7�{t=bI|@�����,&���ѥ�E�7�v�^��\w��A�!-C�k�q�iXCDѡ:m��s�U�ě"�f+p<j��D����ɯS�M�*.���	o�g��ɸ���'�]�jwP2�ɼL�/��zҀ�	��]��AXq�%%י,Pܑ��Ͳ�j�zo�n=dl�|��?{S�GH)q�{�{x�Q<�a����/�Nrh~��מ�X7*���1�w��WfN=�������m3�e�·�{�\d��U���m!G}Iz�x��i>�xQ�lf�� b'f4�����M����{O�ɔ�W��2n�b'���}�M1�GI�x}���Ǐ�{�g*�ؼ�u����(^�W�7۽7.�G��SD}>�y�}���i��c_���=��^�S��}�c�;����5f��Ҏ�r�6�99�g�k[����v�f�;N�|0i����wE�X0n�B�[Ol��㕕
C�2[�
������a:����SI�w�G`f�}����}�����hGAn��Ǹi��{N�o�]�n)�`��=�c�I]�{��+�r_*ѐl���w�^#�ԻY�aa���sۯ��7X�B����E�b]nm�N�Jx�&<{+�/fǪwG$`������IP��ӭ��^�'��nn�^�	�
!6��w׃p����5�s���>s�W���ۍz2��`�Onq���pq��=AX8}e��|#������w��Ck�L|�������zxg4\�d�Q�e{F���[�fQ�m��h�f�kͻB�o�{}��Y��Ttz+u����d��c�h��C㾾P{Y���u9��f&;�{���H��TS
9��{�w+�%�>�`���,��!�'B��|��K�,M�����G�E
����s��M�+|�"=�N��j�X�J�ʼOAj�)ub(}�d}[G��Og;��Vs�g�=^2���ܘ	��$a�]��}���=����3ow�����p��p��r�"�7|�;����|k�]�nQ5��K�LQ�^y*�wA[0����Wm�f[Y�U�*��B0�@e�Ufe&���7TL�jͰ�U�T��_����*Qʘ�pR�	iƎ<��3��AZ�~����ʦ����o����
�n���QP"f�f��;uQ�z7wb|^=�	�L����Ly@��u]�}�Guǯ�@�$軻<�۴Fjߟm�{ֺ��S$'`�������WhɈO�@�Lp8����@�K�zk�V�����% S�;��UV���l�fF{C9����Fj�JkL�݇Z������&�����$ʈov=�[>
c�b.�k�5�ső'j�Քޭ�T�2�v�f����M�RkcW3��]��M�/DNrn�<;uhM���v􈅓F�^I.X���wƪ�*VnJ��}z\��=����B�����hf��=����C�tY�g`�n���l�#˸(bљ�Ȼ��7��s��*p�U������H��{
pM�5�TC�v䩨cA�,SĪow{}�g��s��=Y]
��nU'�
�|f�f�,_�9}Ӹ��ic��X�;�������n���7X[X�Kupk^DZ�i�9d`ئ��D�fF���T�٧%�W@���{��^ S���W�}��o��;l�Œ�k`G�5���z����F�>��~��*���x��W��7�>>�$�m	Y�o0����� 0}���O�^�6r��T�a��F�8n�PD����� �b��o"u7�����|W��&C�SznzJ:S�ׇ�^i���Q��"�T���d͘y�)c��;���ž��<q�v�7�8�G�Mw��<y<���ٶپ��)����H'���473g,�����!E���u=��w�X]�}�����z6��^Q2��0���a��-U�]Dz���r�޹��E���ֹT�3kjl�:.ֆ")��c<��ʻ���܈h@0���g]��E܉cک�ѹ�ݪ��TZ�f�'0�v�C��O]�R���cvUz�}' �tԸ�0&r�έo�84[-�>մ�T�w
ዼ�E6�I�ւ�XSGg6al�(�Z��N[��`Λ5���h�p��gbn�(R�3p���� ���w����{{Xu��ݳ&��V[�<1m�۸�㞎ۆ�wW�4�c�9Ͼ�m�z�gv�5�<���?%׮=^�Z���;+yB�k�a�<���>�ow}J��!�����o�d���<��/z{/�m[�)!f� k�^��r1h\�n,��H2�p2�]9�az�f���ܣa�暱	�z�1ܶ5b�c���O � ��5����L���@y09bP�0"�F�I܉i��.�i�yx%�I��eӨtUլ���1����ao:d�{��%������M/z���wܝ�{ʞ��T�({]��l�e�tbk.�j��tOo��~x�AU�}Z���tW|�|sz�5�ѻ���x�+(7=D(����a�-w��9'���k�l��N��<x'�S��Q_c� ڰ��[��
Q��͉Q\���r۪܈>ѳ'��ܳ���4v�`�(�}��
�=K��e��XZ�{�1C�׍���Z�Z)�Q�dͽ��&N=����	B��^M�ؔhC�O/���<uZ�CGU�%wK5�Hw�xc ��~�כ��/^˄�k�j�3�qڜ�pa�B/a*�w��	�z۹ڲsz���v=��vSϺ@)��a=䶕J�\����f�ȥp�l�o5���ndI�e���xy���v��|�l�Ǆ(�tk˃ueG`���$^�ü�#���� �$:�v;\Ď�&w�����N�f#�/�Ƕ�Ǟ߅��yܾ�,��/^ �����>��{�#������3Ч�Q�n�@�]�0�uK<�n%}�����c#j�{xgb�s�ۼ� ��@�[1bSa��[���'�4}��O'Çq���/M�ݠ��*�8�_���|N^�vy�~����[`���3(7�A]!�{X��z^X�Ȑ�S�G ��ϟ����s���H��^��xN����^�9�+�pgt�_8�@���nt���拦Q�7�U��(+t�{w�kB��=7�}�p���w�:�{�v�'x��]�g��ᐽ>�����\�^��Df�_8�D�;���LLe:p�e���D����`�XZx��@��}����גfb�^�µ�y�N2��S���j������1���(�IM��z.A�.���X xQ��>ڍ�Y��]ב= ?17w�H�f�P�|�o<۶�-��7�t;-cPnI�U��A�Wo,U��3��v.���5�Jf��-���`�%;�'rr���V�;�٣eUn���G	ũN��]�m�={PY���[i��d��.�����Q����OI�w��c½��J�Lb��fb�N^P��� ��1���j�s�@�� �+�c�E�,ɹ��0���-��;cH��!9�gB���=�to����C����[GG�� ;wv�����F��W0�����Na���uOn�u�j!U�����A-�0b�[�6ݾ�߫3��鱋�>�eF���0�<,��<�y��l@����Ox9��p�ݾ�p��`]٧BnɹW�r�gE�E��8>OM$�e�y�}Ua��]co�Wl�'U��ܨz%��]o;�¾�z�"���������!ܹ �x��)���练}|.��õ�&�(7��m�}MŜ�2�&�؂b�Q�3�x�;�eCwnN-:�����k��|0m��_z�ѕ&�ș����Ma3RA��w9[u�1,{.��MlIZRL��zb�[=�Ƴ�;�ٓy7wk4��C���?=��{���U+Ñ�=�j~RqҵAg��*��)�ĻaE)�<R9��^�}�ե�3�þ��R��R����V�pVI�׎٫W�"�b#�E�\������y���ި���WSTULq�N�[T
ӌ��C0g#o"կMf&4=׭�V�
��N�n[=B�m��v���#�{8�كy� YY��Ȧ�r�N墡lWHm޸1�WN���=|���)��ms.�m5�^��W����>�$(�O�ά�V��1��@�u�W�>�d�ۺ3I�e��v�?f��kޯ��ϭ\�p�WI��c�R于˳���� du�|��2G5�g�#uS��w��^Z��;Hqd3��S�����׺pc�|�����s���Gu��}���vܝ��Ab��y���Ü�9�xh��c�� .x:���=w�w@�jk7.�#S��_w��w3�m�b =��٬#�M�'�q��8�zLHf*u�#V���F"�R����w{�2�u��^Ay(5M��'�:��]��z�c�o�{sۃX�B�Y�T�k}�B�on���aٚi���za��z<{���}��A�0�,�	�Q����(�2��=v�)���$��=x�1��$�T�˚Z4K�(�iQ%�d�g.�s�,�3�r��ٺ�aE(�:H�؇i�-���Q�V;�W���3���ZL^��o=	�7)��VjJ��4
��*��]Y�:ک��bܔ;˼����F��T�c�-UT�N|�\�p�ҩ���1�a�TI�{W0�n��p�܂�ʽ��p�����/z�A� -[���6ə/��p���h{��U�7
QQF��������uw��Ϻ{��`$���UfƯEkKZ�:�B�k�vYV�8]�̬4E�	���6c�IL���m�1��,u�AѥΩ.ȱ��JV��vcX�.��\B�np��k3� 1GFk6�lBj�B@e�K]m,0�։/a�г8.-tم����Vh�B1�͂�6l�tĽ��	�]�z����0�ΰ��3M�y�3A��G%�նX���`-�:�Yn#��-ocM.���a3���inK�!dv�F�F�;��	t�ڦ"`�eŚ��6Y��L�fMi6h���c�D*1�,	Z�4�Ӯx�uؘ�a#1Bm���4�tl��#��j�H/gBܗD����`����A&#o&)5s`Κ�u�H��_�hMCɣ�14�T���������.�R1m�m�@�v�5[0�˂��� X�af`�G\�&��6l,�� !��J�\��
�7hQpk��:kTn�6a���\���jM5İ������wb��Q2��¬ô�m�����JZ
Y����f��X;C��լR�*A�p�ۅ5���m���1\��h3X�n�f��͇Wu��-��f����T3�1��cFf���a�	����mQ�����ـ5ĚŬՓLb�WLfF��^���j�ך8;8P[��X�v\� b�e��Д�0CUͰ���6�f�
��ai��j#���
f�4�/l�&�̻Ո�<
m�i�d�3T̋*�[M����9o�bچ�	v�R��Gi�X�"�"h��&	f�4nyi�kp;�1�
0�j����@���YSLT�����䖫��p��ڳW�@��2݇B���/V6k��Qgr�U�6۶si�aV^&Wii)��\��TB/f����9�������d1����mZBVPh����[et�����1�SX�c0�ib���.S4�-�4됰��0&���"Kc��Ve�.5�U"�bYt��V��W�+]���nr��q�0ӳ�CJ
�1�d.��;a�[��6�h:1i]r1�@63��E���j	��7Xmc3M,�X2ҳ:-̎0%��Wb�,��c�9٘HR��ԇh��+jb�L����v���J�hB&!1�0����J#���z��(X��*hb٫X�6�2\��X�#Wٚ����\a���%�ŗf9�P����H�¸q��M��5Avf�R�Y�Ң�V6���ɘjE���L.Yz�4�Iq!7b��1Fj�`��b�ڷ��]����+IP:�*��kt�8�S��.�g0�5�F�0Y�-�kN+��I.�����g��&�Lk�˫p�%�c���\��2�n��걭���̫`̱�s1��L7ZB9���%�HBf��%qtIiie�aC��Mc�)4!��3.t4LA%�č]`Y���m.��:�#k:�kg	Y[�a��4q㥙�$�ȗ�L룚%��2�AX#[ĵ%�f[lwR^�pm���m�\063A�s�6R�C���V�X���ي��hf-�R�� ܒ��8(nX�]i�Ut!56�6�6�p`겣@aJ<�n��:����X5lŭ�����hN��b�uRl+k��Ż:��-i]RdA�c�r[v�+r5lF�7b��u-�kGa /]��T�[��
*#1Ie���"�h$4�ԫ�u�0�NK��qk%)�͵�e��),r�r�P�6L:/2���l��^Z.�P�D&)��y���⎻,��5.jJ �@�LD,��ݱ^fp;"Ю%�`���L��q�KfXԶe�\���ڈ�2�W�U�%rT3�)[��3ԥ�2���Uô����i4����5�%�"�{+1qr�l�cv�DeЦeUPps��f���u�ha+CM��\�їY^�5�	��Ѻ��G�f� jۦ,\�f*5�kjYtcA�`*���4-�0�GR\�ۃp��w2�$�ɢ�dR�`�c���!�A6llZ$"R��\BR��6��JiT�b�a#�ju�gB��j`���b`�0ܗ��.#bb��H�FiB`��rU�A�7:�d�b��[a�D�F��F�V����2R���<c���n��E ��j�"n�!b��`���VUP�W[D��M24�uRUs��ULv���4i�Xi�ZKsZ%���5��͆��Q%R��ؕ�A�s�k,	j9$۝��B��K�#H�B+ft���D�N �SQp[s��q�kNK��l+���	��-�lb�Z`"]��*d�Z=���r���aZE�I��\ݒ��f��h$l��c�5&���j2���Qu���\$�I��j
�aV�1\��(�	��sk�)��F7���:��ej$�!h�%�f�L��,-�blZ٨�
�m�����2��!��]ά����P��13�V���)�%�֢�n�5�kf�3@m2d�1�s�Q�tMM4ʤ�I�ik�fہΤ����V��c&��I-���ȳI�kie�h�B��j�Xj�-��z�P&�"]Nۈ Ff�SB�t(�Zbfi�sRۘ^ ��(D�5�@u�/R�qZ`�8%��ͨ�A�b�m�J�dݫL���:����1�T�a:�j�Z�6if;����b#�fc,Ύ-h�b�6�/]MFZi���aZ�ʆ�����X�J@����mmM6U�9W,�D6�Y2
G���W4e���҅��0P��t�0-"�S`�t.*�e� �VRhm��rU",*KVm��<��� /X�*gK.��j�uK�\81���k8k�B��]fu)&j���uJf�\f撰��X�jnE�KPef�E�݂�m�.ٕ���k���*��#,���1f��6a�C^�Z��jK��n��e�������V \��ǖxy-a�P-!il�(S@�ƥ!,.��XLd�kB��%�p3M0dX�SqO^>K'���-D�c����'6ڶjIe�c�&��������5�����f�k@ַGa�R+�g][
�e�fK�R6R�Q�	2�M
�J��m�J�c��꡶�&��S*4��0E˫R�uP��Tp��3��h9�PRX�0�6�P������b֒�q�6��mh�D�g��Ƣ�YV���u�n!p�K�]����h�F�eQ�c��4c�u�+\"�Rل+Q�ba5-4�!5��Y�91vn�G�ɘ�J�u�"[X��#��Z��@�L#��xkv��L��^hs`����f�LCDL�H���ڶrg��[�&�],Z�m4i����a����rhD�n�Y���m�a.W;�]c�e�S�G���lRn&IU�]0����+-��q]��Mq[)�	
gCR��)��WT�jgj��Sf�:%�F��n�$V:����%�6`[�.���e�iZ9	i��F�r֙)5�"���M��q��-c�6�+A��Cq5��͸�	�K��_8���9��b��[�a��Z���c*ٻ4�9a�D2�	��� gj�i6�髥U�Ҙh���7*�[1���-�e��j(l#6X��;b��TiZ莸3\�;`�#w	�T�%KB���GF�fm�y�xJ0�S[�.\u���V�P���aVۍ6Lm+�����c���]ɊZ2Y���F]rCn+�T���a؉B�6��o.��Hj0ئ�r��1�m�:˖�i�$؛:��2�)�����W\�D�E� �Yy���̕���YrC�u 4�@o�Į��tCj�E��jݩ�X�m��se,P�����5e֝�H��¡�Ku�<�0�i�+�7uWF�f���.��"�r�SE�Ri��-n��"�rԴ�HkA��̵lZq�yҋ-�s5�d�֨�5m�fUr2��e�m4�k,ƭYs�"jd٢�e�k�GQ
13d�%�5������6��.�H͇[��X��mD��SZ����ˮ4Κl 5���8N�5�aܲ©�%ڕ��]MmM��ˣ�f�*�R�rڴu%3����̷�,�#��|�<l�WEJc��m�-�Klk�63n1-Uaa��q0CEh��ij�̻۬)h;K]�i��.K!5���MT�ۮayQ�f�:���31��K+���\!-�Y�5���\�5m!�]����Q��U�d�ۉS;�"�B�sl�R����:�!��2Aح�#��F�T����iWj�X���@����e����rm.P�x�� �U�Kit5�X���I�Z̶�)s��R�ٍ3����!65à�T6"��ji6f��53@��@����bYj˰u[y��^�7�A���6����)�vPt�f@l$����5�r+Kh�3��� �j����^a��Yg�*�)Mb*il!�yj1�К%�:��`��e�8����f�_6�������<kB�Rm�e�(m�fԙ���6� ��f�5
fm0.�V �`]�ZJFΗ��e3r^WgT[.�f�6�C���6c�1Y����Xn!b7���vL����V�3L�K�c�H�p�tf��:�y�|��4BS&ƹ��7&W���F�ɓ.����"uF���R�[b�P������3�+lh0��cV�Q��Es�Q	B�;\�m�@f�1ce�ӵٻ���!�k5�r3��ĺ$f�)��;]�6��F�Ϋ��ك��/^��SJ�	K
��uP�Į³t��-C^ˌBkoXV�,�Um��(L�6������#��Q.��d�v���g��eY``؛A�6��ŵt6����bWMl��3���eisZ��mvlH��������1�6b ����1)�η���b+��iU�.�!]Z��V4�s���L��.P�G�&Yn��帬��b��R�llѱ�u-��7LL �Qv�p顡B1Dլ9m:�FcV�X+�2lfЃaGM(:,��k*l�k��f�f�Ũ0b�&*6�ʷp	�A֔ث]�:��K;M����?�k��2�����:%�6�9�z�f�9mY�\[h��ud{�f�gggi�du�Eg�����١�67E�n�m�X$)�g�N���M̂[#�ѷ�y3m��%���w�����X�e�M�m�&��6��4�7;0�쩴u�e�,l�[X��i�Xۡ36٭���[��\�/-�[�U�A1�ޥ�m��k�f#L������!�6p�9�%��{n�M#����bm�n�hA��lj����(ɷ&�FegW������-���f��@���[{֖m��s��;laim�;=�ّw�Vs/{��-�48i�%��Y5�޶6^�痹���[k$M�knJ��'7�F�T��I'��0m�i��i͙\C��а6�.��
E�[A���]�f�J!�����L8f�4�3!V�^&�ى),��TP����b�q1]]
�u�]tY��-$v�Df�#�%KLh[f�4����	����{]Ņ����`�`k��:��)�����AtZ��,�Y�,ff.� $��6�v�k)W�˦%�r����eZL�@��iĬ�[5��*�@a`���B��fZ��Jp3D�e�kn;+El��R��t�y�ak�P��1i��*7K��h�1 6T�T��1/[(����9i����%�k	�-�a��j�3L�)�.�Ź��E�t�-��Z^�-��cKmFT{L�1u��"�3`���δ:�j��rA��r��0��K�Wtek.��\�7KVk�Q��6[c��1Ya�����ѯbeBgA�M5�S�_;��Yc�y���\�.Y�P�Mt�a-6i�z�ũ�iAB+�u��7�mk��H�k6���լ,�,,�ղ�.̧L=��0&],]Il�(��V�U(;#s����t��b�#�� Ů�X�h�`e[P�:m-+�������Gb�6�;�B8n.# ��h���YS0=�Z�F�U��Ŵņ�1M.
qfQs~W�-�
�LW������+1���4҅iK�bY��bmY����MpP!���9�Q͹s��R�&�ֳR:�.B&���ƺgM�2W9���32 ��04�Xd����V�	s*:�3.�V�(�a���hb뭰-��k1�, \�pfS-�k^�Ų��j)��q�$E�
�m2�� �mu�3Aղ�ĵr���؄u4V�4uΔ&�e��R�63�L�UY��V���L�5�]��9�3��LU����2jpS�(�V�BR�P�l�sn��4��Jʡi��I��V�fcp��Q*m��1���րWC(�a��hΒH;XÔ-��5aZȲ4�*PBE��Xޣc�6ň�@���F�Hr*�j1�b2�6����S��B����#`�mUjZD�j2��V���m�y�"l�{c��m`{�-���Z�ධ�Z�y�z��)a�aՒ������Z�iRn"� T�)*���c�_�?�?ʿ�Uc�y"h£٠k�S4.�h��%����VՖ;d���*��{4`�>Q�����+�����8�r7`���t��J�#��
��g�DBH��
=T��W'�����5 ��%I��
��싘x��@���D�엽)"����ǹIH��������n�oO[�̨��y薡*��>�#�� @�@���!)�$<����%�nU�^�9M�y%B�yН'�o�2�v�$a� C�"�-{;��>�]ȠOG�����JA�H�	#{�т�%jg��\����Lew�c싘x.�*ό%&$�^���9Q*��
���qP����յ��ti��3u��˪�4^�Bh�ף7�y��М�\b$Al��J��yB<*��=ܝ���C��w p� ��5 ��	|�"�r��#vX�U�ԗO3fTӨ�:�s���s��~;@�zJ�}�ROw���,�?o���O�B���rwV�8���2���Ꝋ2��+'�G���z8��|o�+��H�=!��� %<T:��n�%�1U�D�܌�ni�!t��	H"F��H�ׯ�{�4E2f:���cy0(��O��>0��J�@JLk����̛��U
���BDe�މ�<8�G��g�wH>��#��R�c�ʡp�5���+D$��>"�)r����[n�y�R���m��qX/o2F����P�#��X![��r��ENuN���4.H82�6P�	���tl�ե�11u����U�c�`jb}&�;d8�"F�=	H"�%LewCy슘xV`L��!/��>�$�P����J}w7�=֧��{,G�o@�9�H�����g���@��BH����&�*���d�"�@H��R`G�T7g�� ط���ӑ�{�xbg��C�����T��J�{���4�?JR�1�^a"ƔOL�d�Һ�&�3�u\�ň��M��g��>}\?n���gxl�u����}$@���Jr<��$r�+�+p�hI2/�#ѺϨJA�%Lgv2�&(v�L<DB|@�ޛ�8o��F����	I#Д�� ���Qw]q�7�+��:�Mic�PN�0s,�F>������r�"�k;��ݮ��>~t}Ye��XQ�R�T��T��vl)+V��Șʚ��&&&�/�~~e�}~f������J���4zs�+&/o d��"N��y1[s���B�r���b���F�q`��E.Ӵ�'�ظ@�	H>��S��w�6;jfE��!> Rg���%!�(��^^P��jH $��z H�����S]Z��ih�J�j)A�1Y�zz;��F��% �DL���|�O^U�C��	I#�*�΄z�=9��^�@���12B3�̇�������Vg�H�� H����{";�P�;�A�|i�ܰ���{'��ozs�A�i�F���]�Hx²�?��G�H"F��H$A���.ͪ;��L�44G\��'�3_l�Ȝ�S��)3�!)0 $�[�:���ūau�����{5x���	s1i&�� �"aԠ�d�:ְ�u�.��
�^�]����<?�V�绣I�P� e�p��WU*OY�zA���sѴ1��F�BR`Dn�"�"�Pz��6�n��w�O�����}��wѧ������y�z<�O�C��sATD�&�H"�% n�bҰ`�i�wG�{�77��q�yۗA[;��>�XǾ���\�2�#�e��$@[E���-O.�܃��G�n�F^Sԫ�*FO(wS���=r�^S�^���{���Ո��,2��̬C�2�ܽ�N�{!Kc�*����g�:��}���9��'ye�e[2�\}08�(�,1CU�א�wlUxd	��.>>	�v+���1�m�{.������q�a�_L�g��^o���^L��۶�؇��n�A��V�:�4�Nͬ64q����.���Et�XW��Z�l����Y�5��	t�Ď���2��L�&�*³36h`JJS�Z�uM���YK*��h�XeU�	�K��J�ftD�frF��k�k��T!��kb��!���6��!6��J\�T��7v�v�"Y���n]��J�m��F]v���Pp;߿�~�f�@��[{X����yb�D{g;�0�(k4��g^�SMV�W�w�X&�E��-̢�J���^A��0,��P4�GMm�ۣh��{V#�e��V"�T���k���vI���O�ш��.a֞���~�U�ޢ�'9e����ڷ���p�yE�����q�a�_#3,��J����.�w�?����2}� ��hü��2�c�e��l_c�(�������! ��'�"7dWd����:�ة�g��C���mג���=W��>ʴ}�,2�2��Y`��=�3A[����C��B�X�H�����}�9�,ʱ��V����S���ߢ5~k�Lf���u����h�g ��j�Ա�"���!#�J�w�hC�&��v��&���w��ONw@��7�.g��ؔ��.�T��0��@#ۤ#vH0Zq�1��}��-'}����d9�2� �s�kY
SZ����?�^Ke�<���|GȨy���s	�$e�X�	όf�>���g_Lk���S�H0#Q��1!�d���VZgj�{�q2�2�c�g)�e����k(GV*��᤿���� �����Zs-x�;��5�⟤g8g��$@��Anw��ONw@��g$\�@�}>�v�00OjGd8d��yiF���7d�}�'$Ŏ�4r�BΘ���tΟk~r����XǾ��s���9����}��}~��O��V�T0E��Uθ�F��6��5�0$,Y�[���\kX����ʱ�&e[2��]���wy�/�usށ���g1�E�od13�1����2�L�-̢�{�{��f��=��bX�̃귥�Z���Kr�H�� C�>�7f,��q\��x��1���sZ����i����c>��'?mT\T�,��N��ߖi�اz)FL�����G�zC�[@��7`����#��ul��{PZby�P�iF�����X��70,���@�\�2��,Lʴmֻ�[�3��v"/H�q���,��|�s�z��}ގ��-�N㤡�bI � ����n�>���ݟmf��u)�*"��t�g�[�X��$\�@�}&4A���j��)�8E8G��4�3��b�恔�k-n�hWc1l+�\�ś-�8���^�ǵ �{ �ݓ=��s+u���΍��{�;y]H����b�P7��}>#t�vL�n�1'�w��SԱ�3�#,���a��»Օs� �D	Dn�aぽS�r�wH0-?,��e�;z��y	��p���M��k=�����t}U<��q��̫�E��'Mv��ޮ��Ξ�f�s���6RɅ���jgF��<D} �o��H<:�r�@�I�E<@E{|����̕s�st=A���i��*�!1����)�j�h1rri�Z
l*��{���U�9�s��U��E�;,Ó�خ�3�2-�b5,�����˺����i���V��;*��������|��υ��!@4�,(��s[iu�бm�(�-bm��	B]q5!}O���#�Y=||}�Dt�W�z�����V,��3��w���ed=�U�� V�Dr�ݓn����gq���#�ϧ#��!�Dn뎨j_N��	���T��i>��~�&�����spc�`�'�2ՙic�j�=���(q��{����*�>Ͼ�">�"g,�2�"9�ZfB���j�V��@�7�2�|D'$�^)u��_z�VNs<#��D��¹�G֯d��_^X��i_�Z&e��+5����k��#��p��^fu����~�e꒾���Qb9˖G2�Aj͞��,��,�Ś>xtm�R��1_�D1���g����Twڞ���6�a������R�1����|E3����[7�ެ}���/YXj�a6��,tD+M4jָsf�[3��Wl�g#��r�y��j�.!�-f mk�f�A.�f��̔4�m`��&nl�
@��X9�8�mU��eU�\ǈ�KZ��ֵ�<�MY��Yx��.1`��4�Yn�$b���.jD5ai�M���^�&-��LY�4C����&���r�ZM��[��2�w��H~���X�ЩK�(J`5q�%��uۨ�XᲣ`��mF�j��W���_�~�Z'�a�A�� �,����]X��\���F�/b��ڵ�E��D�&=� n�"n�"���g"�Oj���"Ȋ�������X�'����&R�i�J�f!l���lߨ�s,�9�`��G4���|,ODWv9�X#L�D	�"#�@ j nW��e�3*��L�z�\�[�r#ݐ7f���e���Բ��\.-VO ��Ps��w<7��ɿWv�2�N!�ՙi~k�R�?��:r�w�Q���d�3�";��H����������>W�ZQX������7�7;`4�������]�	�&m^M~�o~����C�e��-̢���7�ys���f���gWId��Y9�U�B5ό=� F�@ݟ�`elFsZ_C��B$췂����`��1t�d���ܻ)��Y�z$��<2pJ ����N{�HC2�"���i�V6�ۤ��JF)�2�މ��:��z�VO������o&,�2L	 F�5�0#ۧ�F�7H���
�r�J����i�5�ݎ��/�V����c3*f�V�-�p��O?�?�~9�/�,�����n5�ld����	�@��r�~8�T��O�F���x�vH�n��vmov�y�$$f��0]��J2߮�d����	O�d��wG����?|�k��m���9 ��,�G8b����ق��{C"Z\G�kه���=��B?oF�vA�ޞ�]�Tb��"2xG���� |7޴���{�ZqJD�.&�<k�������0~��E��>w���#m�O���7������љU��LƷ�ᗖX�}V��*��-3*�9�!(�����U��y|��=ڃ	a�.8���A�,�tj�u/y�
ܞ|�9^x���Im@i&A�����=)!�dK��kLS�G��
^�6f�ֶ`���L�:�@нU�־�}���mҶ#.�ɒ��+`b������9�&�[��駠�����U�
�f�0�>봻r���rx��M�D1�&��vq����T�RE�Cl��.�޻��˼7G���ڝ;}����^�O��f���߽�ekJ��R������=\�l��x�/{N��C�i����/3vd�&�!���n2�v���.rL�E��E�%FT[q�a��Z�)�@<nBrA���e�Š��[�8�U+��a\�m��:|o���A����p�k���i��M����*w n�z���F�N�V����v��(��^nvM��V�,����H���M��'Ec�C��I7h��Z�Wm�\m�X��n��^���}���h��<��kNG�p��vm�;ޅ�h� ��� 9ꗈ2���ϙ܆�8�����Lj��=��=�u�j�c;=��x"����!eV˄�����qS%�QR"��
�Jv�m�]	�Y7��]�8���ͬM.��s��;�6m�x��F�j��+���|�����V�kR(o����_]��e:��gS�Qv)Z�kG<q��ww��#��K[���X��<�<��<笔,F�'x��ץ����t꾾~xÇπ$��Ay�`����e�,�kz�H[ZV�)o^N�t%��9E-mm�{�n,���,mg`�Fn��ba���m�W�ۖۉdY�bٶ-�緽�<�ȶn�����n�B���-�i�Z�m��0���e��+9�{���6�C7,��4����H��tw6��d۳�i��km5���d�nn�چ܅�[v���Z�e��[-'6������k.�&h����b��񭵸S-������j�嵲	�4���Q�5�b��fȲ;e�ɶ=�9=&��5 ۶��͘vѥ�-��5�oNg9m�chY��bf�� ���vV�,5�g.Sl����vJٳ{{�G�ݶn�:ڽ�^[e�����9�
ڹJ䋿�� ��@�Y�2S��p4	) ����4�R
9E�؅$��p	I�9A�:H)�o۪�+���E�B�RAs�p��)�}P�j2RA@�(���_o��������~4�5���i ��a��$�!L?~�[&�) �o��ߵ�|��ه�_������A{��
AH:�s�CI��9�-4�Y@�O9wCBJH,+��i ��
@�(��ž_?7�����є���]����{�u���W�����A�:H)
�@{��u(�$����ЁL9ʅ�L��P9�- ��k�׳���߯��Ȼ�Y�q�]���\��)ۈ+�睢mu�c��۴�R�f���:�i>�t�褡
a�T- �z�H,ƒ�]��TAH4T9ʆ���w�=?}��W9��vk��<��Qi������ƽw��GdӜ�������ᤂ�L)���hB�%�����i) ��(4� �r�H:��[�k����ۙ��o]ߠ) ���-�d���AݣI����׿[�>��Y\�{���Ao.��
Aa��d��H(w�i �4�Ay˸ߟ՛���V��
A�P�چ�� w�ZAH,�d���
�) ��rᤂ�DaH��HRAd���p�~��^��|X��Wխ��~���ׇ�i��A��AH(�E�Q
H-s�� ��
a�T- �4!�Q���L) ���j0���>��߽����o>-�׿���P�O�RA@�Qi������J�
A��9P�Au��>;�����}���k��<��Qi��
A}���R��k���r��꭯����h`g��j�}L;9��\���u�=�tz�{J%Bh�5�oV���Ѣ��3�v�7;�ܢ/��v�+���"�ׇo��WϷ���H,<0��I�B�%2�ܨ�Rr�`� �(�����!I�*�� Sr�l`Ok7W^��|~��*�� �����F�7��� V��`{��g9p��3*�&e ?�^~;�V�8r�~)��[d��k"\��*�J4ҭ��lGY��*�i0KkǠi���
AgFJ{��ZRAaA��i ��
@�(�����^r�Z���o��}Yݿ��H,/�ä��ֹ�Z��t9���>��}D) ��p4�R�BٶJH(��Xi�$���a������B�
A@��W~�;>H,4�^�ZAH,;ʅ�7i�����-¼x���@`��)��hj$���ᤃ �߾���Ņ��Q�R���m �v2�z�Z���C���P?v�H:(�$�ˁ���@��B٦JH(R�H,=V�� T���/��qY̮�d?0�AIHSިZAH(�l�A`hi ��@���uP�*H.��9�-4�I�[���ߊ�~�~���%$f\4�XhaH�E��!I ��@�O�er��V{o���������:H)
�ߨ���!I�o�}����}�H)�r�l��I
Cߨ�Aa��$����I%!L9ʅ�j2�
9E����T��뺫��ܫ�H)EC^�i �ߵ���?w߷�v���}��>�-?�YC%>�P- ��B����Qi!�P�L%> �f��ڋ���_�'m����Iг�wh� ������z>��9��F�J�_��p���J�qc~��7h�O���w9��bvWUOT��]s��?��x��Af��Ѹ����(�P�P�MT�-���j�E�I��\�W�.X�Z���.*��gZ�&s2��	Z�+(�ic�u.כ@*��x5Rg3-���%��n,W"���m����֨6��,
ݗ	�uz�[�:�6\ Q�T�ήF�uC4�%lT�ԝ��*��5#��&�n�e���Y�8e�,p4+���VT��?C�)�˭�KMk��	Mf�6�Ga.�-�Q�uZjWM�T:uZJ)�H,2�?�� �*���u(�$��j�Rr�l�%$r�H,5�3��ǵ����ھe��~��yv�RAIw��uߎ`q�z�i �k�ZA`z4�^����)���T4�]0)���Q�*��p4���_=�r��k;$Rۢ�hB�%2�r�����ˬ����=��__�~6�Xkꅤ��?~����$��j�SB0�*˯Q�k]����H(��H) ��v0������B�42�
9E��H/9wH)�9P���׳�z�u]^�埢>ȿ��\��W��� f贂�Y���~����%$w�$�)���
Ad�)�.�(�r�@� �>������v�=����Qi ���H)��w�f�) �B�H,5�3��Ϸ���~�|���~��ywH)?
a��d�) �{_����ߌ�_�Z��$�H/�]�R
A�T?z����`R9E��
H)�.�(j$��§9p�Aa���Qi5��������'FSyw@��?z�=����U}a��Aa��?:H)
*����H) �wZ���Ü�[62RAB�9�4�Y?�gￚ���>u�~%kM@��U��
چ/ЉWX�w8oTfX�Ӏ�k�~�l�o�k�)'�)�ݨ[&��H(��H,F��]��TAH5P�*H1Ao��C�/��eʼx��� xY��ʷ����{��u��[��p4$��¿zᤂ�L)���hB�
Ay˸
��r�C�����9�- �RAw�_��k�U|o_�����G�PiRHELU������)8\��hcn]a�D<���\[�����U������5��������.�&g:s�}ڣ��H)��s�f�%$)��$�o��ߟo��������������R~B�~�B�42�
{E��I�.�U�82��W�l��rJ�n����`Rܢ�
Af�)�]�R
Aa���i ��9�-&��Y)��p�U�W#a��Af]������Ă�_T- �?U���tQ
H-s�� ��Bٱ��
�9F�
AH/9v�) �����v}��Y��ߪ�є�P+���A`i����*�)��CI�3�~^�~�o�{϶_ߠy7E���ђ�~����$�����C����Qi4!I��S���P4��Xs�t�RT9E���]NsZ���Ü�[7���x�Kw�IԂ����Aa������n���ߎ�7����m ��a�aI%��ꅲhe$
;�4�Xi ���URT9ʆ��xLf~��9=���U%�YlN�V���]�i�m���)5\Y�!3j�k���I=�1>�JYL��p4��
�ˆ�
A@�(���Y6�y˸
��9y��m{������}A��AH^��_?g�߇�_�ZA��RAk3Z����ި[6�I
�(�AH)�.�q�$��0�*ɡ��P+�t�Z}��$F��]�R
A�P�jH.����Z��w���Oy����@��i�@��ʌ���wCBJH,(�.H,49�-%���u\��x���ɱ��n�(JH,9���
B��;�- �Q
H-s�� ��0�*�%$r�H,+�to���{�5m+�#�sՎBOX���8����,t=�'y{t�Y���'�P�G3���ލٌ�#=�����0�/��q��� {���w_xd����G���
a��B�4�����i����]��Q ��*�]0)���H�Y����sy�ޓ}wC�) ��۸i ��?z�I�) �����k}�^~�m����u��~6�X}��� �*�ߨ����RAl��7�����ν�
AO�)���-����P3�ZAa��^r�4
JB�s�d�) �T�,�A`hi ���
�v�U��S�$O�t�T�����{)��:������3tZAH,��O��p��Xk;p�AH(��pB�
Ay˾��!���^�����~�/�,Ms\K�vP���X�2ۙ�F�rd�ٻZ���,FJE��xH,?]I �o�ZA������j�Rr�l��I
A)�#³��_f||����� xD$��`xDw}�ɯ���'>S?|�7���~I��f�
AH/�]��Q �P�*H.���Qi��
Ay˸
II�W�^ʽV���/ކ����E������2|@;Y�W�A���9hp�Aa��?�
B�P�QiE���;�@R
i�s�g~s���kZ����RACB��$RAy�
AI��0�jɠe$r�H,4�^r��Rr�i�;kr�b�vE^l�ٶ�z嬰o�@���) ��J~����ü�ZAa�� s�ZM!I��S�]�P4��Xs���
B���o_n������QiE���~֠)4 S�B٦JH(��c½y�O}}��=�R������t� ��!L?~�[&�RA@o|�k߷��G����bZ ڠ��ѽ0P�m<�v-�UQuMބ>���d�a��QҌ̉��e��&���r�M$eZO_u�c��^�����$��é��i ��� �ݣF�r���"s�ݙ���}�Z ��~pԂ�x�W�Mt��b����Q��&�/���߿���o�=��qDqV��%R��BS/j��ݍ��ZJ�\Q��cf�m#�`�e���!"�n�t�i;S=��7�Z��\���]�׵E��T�+�`�Qq3(�F���.�ހԿ@��EZr�������Ճ�� Gt����S�S8+{O?��_s?<��O֗��Ӛ�O�I���ޞ8��UNns�U����yfZX�Ne��3���LYw�y�2��Ԙ����L�.�ڎjv���@��-gMR;��d!�Ɂ�`n�>�����ݝ���]�]t(0.�5�e;w�tB[f���� @�&$A�Nb�a������K;�<�g�m8�H��(��KL�Bb�]�+�r�
Y2�W˦�ºM'x�AqU�~Zp�Ҟt)�����ި3(7�4<�
�Ə_އ����ljZ\�m�i�l�����f�V�B��f"ii�T;7s���ec�դ���c�F��KfIE`�72�muH�Nxݺ�
Y�i����Q8�H@�hv)tR`-q��4YD�̄�$0��uAم�iv嶅˨�[�&��JP�����VГ&�9�ĥ�6+mi6��*�`MP�vu{V��fSHMy`HU��b�)-2fj�eMFT���aY�͘�[��±�.X�V���u8G55�7��:TMh���,�V������7�-̫���K;9E(��,UH뾭�k�b9�-�*^e�&eK�eX���3GN9�s-M� WI=���
o�^h��;O.z�D���ǳ�_h����Yb>�#3,3+�s.v���ܿ����צ�+��
�[su`�@��>�_e�|2ՈZW�/"���r�G��C��sp @ݓ뷥�Ӆ���`��������M��y粧r�'{E����K-X����c�tN-��Y�ߴx�޼�O�M<�����@���`i���8.?�{=ɂa�`C~H�c6�U�"��6�đ6l���5Ub��Z;-�5!{���DGd� Db�Dnψ� ��s�yë�ػ��\�ָ��:�ծ	wI��"�{�.9�3*}2�30��ݡ�3y�l���M\��)�a�y�bPw�#A�h������wge7aۓY��5�D�PF��BjZ[5�d�6nw�_�3ћ>0;����J>Ӆ�{7�`��DGt�#�H F��誗��zq�Ys|�s2���fY����٪�_+����vc����<#�:�n��0s(3>,�1���F�9����7H���^pn�Rػ�s�}'��=�1F�&�I��X�nO�� �7d��-8��b���<._�����W�8�,sٽC�#�A�����7d�fX�h�`�y�˭U�M�*�j�	p�ͅ�`K�m6�Q�6y�e��R��P)af5�;���Y�r`c�7d���g�Zخ�{3K.zN����ƃ<�XA��"N!��X��ai�䚝��/����Aޅ\�;��-����=�!��9�,2��U�}�����w����b9�\s*[�EP�+�e>�L�k��T�r2��R�]U�g&�79g9���b���v�'t���ۚ0,o��ưm���6�2/W�������d�ےǻ��p�z�b>��.X�T��e�ez&:�Ӯ��7=�A��H�@�"�_)��kvM��f�T����W�%�,��w:�e��e��Zq��Ol��i�BZ&O�k��s��<���^F=�X��,3+቙s����tt���Ϳ}~o�:��	[p�$�D�z�3���ٱ*�S�쌴�04j������^�������\n�"�F:�X糚�]�-�ZG��~ߟ'56q��������j�2�`DnɁo�j�ְ?@�$��5:���|�f����YS� C�Dݛ[��K�L�Sr:��U �r�wHۤٸ��0�V�<�6a�rY���K�y���3���e�1J�J�a-������X��P�-8���֌vF��p�H�#��{b 9��#N }���|����ÜZ��%h��ؼ5Qu�1�b�Թ��K���]g-�7��J��ibz�"i�w.3kn'�ˮ�*��ʱ��:��~���������=�ᖔ0O��Ve�����:r��DT���,٬�=�YS�"9� @�->ݛ F슾�v��1�D�
��Ti�Me�i�)��l,[��3*G;k�%�!K��:���e���pOv���b9�^��
�ٽ�sr*��d��M��T�����:���b�[�V";ʆ�o^�r��]ˉ��u͈�l�.��/�5�y�X�k��� �5ݚz��अ)��Ds*�̠�W�s,�s;���9�=Y��S�K�͛�梖T��@>ZA�n����Y�y}��G�s-o�X�e�^�#ۤS�����^V�Q����3�7��^��������eZ.e @�>ݙ��θwq���k p���An�+B�0�p" �����n� n�>MթewKoX���8���-��h{��w����@��4J�����Umⵅ�lE��o��ݞkbB�+h��-{������~�߻^�rv���QZ��6����t.9����D=��5�l�eP�'�Lu����wiƘ�oj�:�U�������B��{�QB��b�gu��J��u6hق-�����7���*�M��]8#�q��ȧ�[`�vG�P\3�,,�,�/�r3Q�32��	��N?qʓ�7dهP�K�����V�-t.f����q��u�֠���,s���~�Џow-ژ
��8wvmܮ�-��O`[˱���;g&w�,/Q�Ԟ<n��!0��̚:���bZǈ� 7W�OC)�^+Y=	�͗3�痼48���$�*��i4oV.E�Фf����G{�|�^�yi�{��f��F�lbAIКZD����]d�S�a���V{�xk��c��By����$x�qg��bzj�q[�,���]�t���S�7V�'w/
3	�sĄ�-�Pΰ�)��
9�Ee]�*�k�%�x���`��X�2�8�{z�Vo�y�� �nuT.����x�-lȖ��@ �k8�Âg�~�^��.�b�8�^������j�I2��m)���rvDc�L;qP��6vD2�]����O���3ڶg����:�{VS��L��xEf��{�LL��{I8�'�[�,�=m&������j��m��!h��KMZ�L�(U���Gm��{����p���� ����iv��Yd�2�ͨ�m�݆��C��tp6�D$�a��4�޼�v�Dm��A-lL�7�z�\���{u�S���H�=�w��YLi�l�gb�r��Z�2�L�-�f�9�Ġ��5����6��\�����u���-��e�������¼�n�ͯ{(�֕�^vDv���Y�	6Ŏ{l�G{v�jkim%�m��6�v�3R$gb[i9�;[`6����:����k�gZ6đlnp��6m$�lFش��m�����ؖ�K2m���-6��:��+�̬�[a���g[��e�N���ڷK�^�����,��5i���)��;2�öܳFfp�^jSӴ�K�ݞ6�8�Z���D�ٗf�sl�9�n��tm���z�W���/l%�����!�Q�������=O(�sF.��ҴN͹݆�M��6#��kYh�b@�M]��ћ�N�B\j��!6Λ]e�F��@��kf�#�3fR���8���B�h�5���j���(Q��,��X�-�����e�)$Qa�U������k�/q���6���j�l�#!l1��b#��1�bΥ�і��0`$\.Ś[�&sBV���f��($��Ї,��Y��ڃ�@��H[�nЋ�FY��Ԩ�İkq�86H�t�S%c���L6�7iRpdEH͕�4����Ͳ�]ke(�d��3RF�Wc��uF�b;+�����ӛ6&��{$c�`0��b�,r�[��*���[p����-����vK�k�1�)F,�M�Ĭj=e��qײ��:�,45�^���*l��@��mY�ke����g�y4nf�!6��ԋF˘ Bf�;Z��U4�9�lт�A�
8��.�ˊYQ��I��Q(mbPseV%L.�	f�
����Cm��s���a��!���Y���5�%�c���3.o6:�FmK]��Y���[��Lx0Ֆ��e`ʈ�w̽XT��lq�L�Cَ�i[�L�+�1�h�X6�h\;��*[5���2u����l����6�l����"��D�jZ脥�y���0ib�hun��l�J�%�D�#�)�=�vn���G2Ԡ�6��P��n�̱���`�&�!m��gq�*���E�s!��� ���r�l1�F�bʧk�<ҳOZa�2V�f�fmc�*�@i�����`h��mV��j��9�mU\svs��ۜ�\����t���1�4v&��XF$va.1p95�;Yrx$�.��Mq4&��x/;��t4ر.,)�ѮH�h�8��Q�W	�H�Mڭ�QnYT#��2^ݣ%pv����JUM�2����u����K�m2�Xҍ��-�q�BÊ��Y����gW�;�K�+�z�V���]U�M�����W��Wc�E�l͘�]Bm"�]��d�ˡ.�s��Rz�rkb���F��7�hR�ʍ�b�b�GM�y|�+D�JA�����F�с��F�S.���iR�H���wg8Qlj0����t���������B�CkME`i4���.�Q�ih����Yqa����5�c"���I��F]��i�׵�@�3f�X:t.nTs�����ڱ*�ln3�1� cX���&7P�F[t�����H�5W��T��&e\c3,��{������/��#��;ft���q��d鐽a�(`�Zq�/�8�f��37�E3�^��>��Aޘ|�7�U�nE�Y^��}V�,��5����n���m�\;��;�X"G���-̫DL���e�V[��c��i�jػc�8w��`7'�稴G9E��bfQl̲��z���O�H�ZO�d\��7˵d��{]B;=����ՇyVtw6�Q[&��,�S�Zq�O�~���~�+�wi��f�
��ȣY�����0#�"�Z�|-YX���f~�b��x��T-�&��.�90�uX� jjX�܅������ݬ�0�O��s;�8`��֖0`������c�GC��c� ��O�#�Ҽ�D�2ǹV"fYi�V�9�l������w�x����~��{�� ٫h*ДlZid�hs���glY鉜�8{=,�,�Jt��]���}��m��Vh�����_�o�ڲks���mO��$A�<�<�!���}<�T\N�r��(/2�eZ32���Hu�ꉬ79ۻ�+2��5�.}�I�9�-3*�3(�̫���w/3YwI�]\S�1YBr`G�f�>���Y|��YZ������oTF#VR6f���&�2�E̫FfYi�[y�w�B7��}�ZA�����U{�a��>���(����_��n:�gu~�޾{S��yt�4-z��ƻ ,�n[p7�Z��,U�f�<-iJkv%;����}3�O{77H"���n�
ËbM`�����s+��Y~s�uS��Xo��ds*�FӋ��R����y'<��Y�R�grW���v�1��"9�0#��\s*�۪{ݴh�����YV�=�\�v@��FxO9�S�s�;{��V�u=^��^�*����,Y�����ld���k����̢oݝ�3�N�^7"嚹�[
!��V�����z��u �6KKrډ�x{��W}7���W��y������ʱ2�L˲��}���_v^nEq�����b� F��<�u��8�$���>���}�0�������Υ`�C�@G�Œ,Bom	�n�o��_��4�a��v�1�� G9@�k>"7g�n��OO]�6�o�����w��F�4���jh�]n芹�	���m��rm����w�w����!�ۡ����xn�E���o�3t���+T��k�^��VT����Ƿdt�7dn���u��S� 6A��<�*N-�9b�zzI�H�̮ݾ�}��f�gӞݖ��fQh�cvH�7d{�㛇�s�Fu�p�L0�n�&0�D� �����ݓ�a�a�_37�o�r�;[����j�3$��S|���-�=��>�G)Ԧi���q�N_Uc�������8����a;V0)�/��\��ݬ׎I���S�x�$�����}�};��P�±⿮��;}���� @��~����gЈ� ��#v\��t?���E��ǭg7��-3�`���>������Dz6��N����3��D�"u�A(|�f#.�z��+v��[M����a�,�0� �R7��~B{� �[ ��#vEۭ��5�v���׽��kv{�hG��q�U�3,07d���������Ҁ��{6A�ζ��gM���\����z9H0 $Ae+�<h�؋�h;�>��G2幒D�#���]��j.H�=�]n��:�2�|^�ȏ}V#�Yi�V�3,��3ߧ�"%���-�x���`�iŞ����+���Xu�$p����ӿ^o��vl{ʴ}�.32�̩a�e���$q�g{+#q��2/YĦ�ޛ5���SU�����O�BD#vO��).Sufg�d�2$h��WP�>}ϔ���Xt�(��ʡ�2m���җCʸ�x�͇�/��@Yy�x��Y}��&���}�u�I }�8�TѢ�5��6�Ωk��`&��7 �5����r�h�X�t2�[��ɍA5��m#[�3��k�kF�L�+)H�s*F�)e��E!f�,"34KMr�s
C2�c�#\��a�mm�!ځhv�\1����n�6a˱F� B�F�W �ܔ��k�KW�ۑ��!����
��
�5��� :�:������TMd��G_�>����(��Zb�8�%̮yF��ck�{j�*$�� �B�%�~�\�Q`��Qc�V�e�kۮ��uϻ&���̿�G+�ؙ.i�\��>_��t��`D�0#��F��Z��n|ʷ���+��lu�:����G���Z�\u�߻��Ttf�E�9V`�N/�֬_Vt�p���э~��:-����_;Y����3�b�>���k<ݟ���?�����C�L���KF����j�i���D������yk ta�	�Dn��`�_j�-:;:����6�B�=ծЮ�1�ְ�q�9$|DnɁ�"$췝R���FE��M}M��F�9��٥f
5l���U��\�e�]��vj��t�x:�"<ʸ�9a�_̠�����lu��q�T�����6�}6��y���y�(0�,��h���X�ev����'��߮?�x�ԏH~t��
SC�4�{M�sM�P���T���o/�cK����0
Ի� 캪�n�FO.�.����X��������/|#>��ȧ����ͻ�T��2�T�����,�̪߳~��둕�-��b Br��F���ݑ[{uz�q�S��Э�1���:�}�"9�"$|cvH���D��c��f\��A�� �El�)�ݎ�X��T���������ئQ)C`�s-k�ӈe��F��Ot���u݅�A���k�����W1��oU���h�,�̫c�s6kc��?���{��u�Y�AZ�\�L�e�5,�+�3-�.B��F1�f��}�d!��ӟn���ݐ}k7i�]nb�{2u�����I־���Gް�+��,Lʸ��| mH��0�ɯe�ˏ@	�[/��n�]V0�5�>�ސ`BD�<|�csGzxL��Ń8�㘲����#t�f�ڊ��yi^����{�P�����\]%^D�Y�Y��H��Սw��b��7#.���h�嚘x�'Q����^�1��.b����33��C��%��hѤ�r���#Ϥ���vH�n�c�R��3>���Q�G=e�}V�s(_f�hW;�;�Ń|��"���g~3w��}ڛ�D̫��eZ9�@ݑ5G"�]iX������S\�:���T�܁�G@J}�>�ݐ��q~����\_��bƀb�6������f�dL�0���:\(�-��c�>|ğg������A�(�U'��uMU%��0��G��t������l�'r��̲�ʶfPn��F�Y���!��iƇ[���}�:|_ޖ#�Qb&r�2��j����Կ��Nv�E�Ո�Yi��c�se8<{�:ff릗lWe��SWs�@�G9@JA�>"7dt��wxW��]^����p#,��r}��=tOwꚪK'(NO!t�0Ȋ�����J�����wػ������u]�!ǫ)�l���^K�����1�G�W~����L6�!�RcJ�'Xk}	�8s��a���Ov˃�V��-3(�->�4�)���8��NS���٣�f�>/��r�D�\�2�̳3Z���������B�B.�3:b-�WE�4��0&�J��x)�������e����cg�c��n��=����l[gd��@�Y.��u�q.9�Y#`@� �l� n�7H۲�b����웩����Et=tOwꚚ���8��LZA�n�ú�ָ޲p֬����A3�h��3)�3-*-V�9w�5�r���٣�=����%�>��9�.9�,3.�Xuq�2J�Sp"���>ݑ{-�=�x����7s�9�Bs�yo�� �) C����E��Ac�E�����{�+oE��Db��ӧ��b�Rأ�"#�0u_e���},9������d��Cݻ�q>�e��Q~mR����^�{�����Ӆ*f�%L�.�U�B7��y�.>�u��xxxWoG�X�+�H�v�r���˓���)M+�퍑1b�e��WK����L��1����j�Z�С��6,�K���T5S�)���Yk��&��f6��ٶ��Wmh�ds�c-m�(�av�ج������i�e���,ʭ��]D�$%�q.�J�X�J�Z֑fL)��Z��E&!	mvq�]����+��L�|��?��S�R�q��i#f%��&����MR�WC:�s.���l�W��U��3*ӹE�eX���o�Np]�zno�W�{O�a����X�q�,fe�1̫N�e}�od����ׇ��{=��l��b�:M���r`G� ���e^��sQ�����eWj��]����.eeZ �#�sC��9Q�f��c{���lQ�o��y�y�X�˗��ʉ���ر</�Lϳt��n@ݒ/��U;�f�}�#��A�C�F(�\7t)շ���joմLˆg�.eK̲٘馲r/7RJc	���y��;}W\)3���y'�V#3�3+�����ܪ�}��[��ZXg�7U	]4CXS-�����֦�F71���`���<=ǽ~#�Y~#��ϷdX�Ӯ���QT�(�s�9�;W}����&�p�~��˙�����bP=8�v?]�����6L��c#એ���{���	��~�n��o9���N� �����R�!bB�����ew�Ϸ����ZwÏ�IkV~���`���I���K��U;�f�r:9H0 F�F��Swb�j�z|)�!�"��n�����2��J��:;�w�\��������^r�ʸ�fT�}b�q��R��@�JA�-���+�u�uB��U-�>���I(�k���Ή�:>����s�3+�fU��E�ek�qJ�@@͓W��I�:�޳9�P��=�.#r�ʱ2�f��wN������~OC�Vh����kQ#e��$-vK����40��j��;�}v>�߾�Y{��={t��=�A��g���&�{�������E\��\AI"��vE�ݐD���z/#gw'��`=�E>�u\)�î*��1����[ lh�'���sFO��v�"GlL�.9�傊.}�?u����`������}����YP��ӴմA<B�aО`�Nwe�h����j��'w��l��(��������.zh�5]��Ky(_�>�M� �����8q����x��k� |�����?mZ`�ֲK������x^Ǎ�7%�"�j��.�]@?(F�ص���Of��Xc�z���'�g�qi{|�ūFN�`^[[i%;I�E,leۈ]E��͛kA!��Ygj�\)V�A��n�r��l$��{ïz���W�J�N{/nݙ�隴˄�cm��ųhN8��h��Q2�V�E�Iz�"g�a�(��hz\�5����X9m���Qf���iʷdnO	x3ssTM _ӥ���t�x�����gX���M;�Kn�x�J^����lADv��1��N�;��ײ��s��=���nX�y��b2���J��q����3M�A��<Ԑ{^p����$%�OL�i�����]ٝ�7�Zfo�iڛ �G�jF��^���,:[��ZO=&hsެ�\��=��LZ矬�=�<Ԛ���|4y�ٹ��ۻ�T�{�5�w#���aJ��������)e�u[nЌ�F�n�)�BVE��l �c3*��n��^Yۍǰ�T����Y�<܋����&1�0���u��QTM:x�H<B�)���&Uk*�ԹN�7��ђ�9��R�y�8z����+� |���u_u阮KC�����0�u��p���H^��k�S:��>��M�/b�a9����	�+���5�'�=��~;���\Xs[�,в���Vi�Z��3	3�":ۉ�)��-�'-����%�m�f�!r%m�͜G$m���dT!$綖�7�nŖlCm�a�H*f��(��kr�$9���m���mlu���rJ,�#����h�ə��{�t��7m��2�۬�9������ˆ���,�������fۢ�ᛜ$�rm�B�m6�)�oz�N�m��Z�"um��9i''8�Ҷ�k;m�cm0� ��ݝ�:�'6��78��kI$Ym�6�)�&[kedsl�6��Ea�--J���Е���D����r'4�Z)"qJ$x�ڱ�tN�ݹV�ц���XٚD�D�m���Ռ��f;���v؈�5������u�Ns���ͺ6��"��p�: �gom;���SEV1@DY��!��9C�vu�s�W��@�)P�ʱfYi�]q疵���V�'�e�ϣ4���:�o,RyD��yiry�9��������}��Z��ݐD��cvpH�\�c�QܧN�\+�Rآ&3�"#�����G�Ճ�g�f���}x��3n#:����4jp�-H2�-
E����*,g��f��j�U����͂3�e��b#�7m�*P�L���$Uq]�%��
k�������9V�e���[�S��t��GVA���q���Q�h�T�L��
{�����$��D����cv���ee\G2�w���CM�������uC�
>��Dz9ɁH G�I����"�"���vK}lD�@�}�`DپnJ��I�팬bA�Dv�"(�}W��oWx�:_n��Jｈ�S6�Fo��lq�~�.$P����ҌL��Q37zEkq�)�5�$�6��g���}�??z�����v.eK̲�3�.��Q!��R���$��QSٞ��k��W�W��}V�9e�eZ"fW=��y-��b���h٘�&fb�<DMLk5�9�J;R	`�riP��嚬!����^�_&�>�A<�A�nɁ�Zs��.��\0k��#Pt�!U����Η5��}�>̟l�0m��v�����[.��+Ls�&�ÌH7�v�"=�A�n�
��]�VA�Ϗ��7O����v}	�%v%��VՕ��2�4�L��@�@�>ݛ���>ݲ&����cEq��j2�{�|�o�#t�NuuE�ޛ�b}g�}�H�5b;��2���ь��`�2҆Z~��@��\����N#�:ܝ��է��&�9lo��l�=��۳���s���$9�a��E��d���S��lh�5&���FU���	��`��_ި�ۯ�����̝�ȭ��x2]�3c�:?���B.iuŮ���ƔmH�1�˚��g�)B�-p�k4-ȕ�e�vZ��V��ՠ
E��m�vnBh��6�KS.�P�Ti\lP�HJ��ƋA�RjB-��:1�۶4�ƪ�k���9c�L:�X$���;L��e�0\�\	۱�d&u�-�Rf
gf���]S%��T\D�v�qS���1cuF��d�6h��,�\i��_�?O��T(�K�7a�e���ã�R�fGj�G�K�lrF��w����!�����i��$G�n�kr���Sٞ���N�n��aE�\�u�v�����}�b.e&eع�^iي�	�>��'��6��:������(�3��||��vV3+���Mz��~�Eߨ3*fVFfQT�����u��<k''�Y��-�ϞH��3+��e�̫��k��t�U�g�h���c����\�e=���sI�����`g���a�챀F����e9�Z9�,s+��{�V��q˳=�ө�[���B��==��- ��c/{�O�����߉���T�Р��@kal���Yl]�GQ��fV[��J5������^�@�D���-�F�zVJ5��A�!��ڪ�!z��	Ɂ� ���b1̫�Q/�B�޵�,�|־�[~����+c�2�?�	"q.sn�+2��E��[hȈ5�I��*�:�7jH�&'"�rz�ʌy����x��c�︃꽮��)��w�������@��1�%Wj�V��L[ �>��PY�r�2�D̳Z���dH�����¸P��Da��;��i���ՈZ~��~Ĕ:��9�8pL�3$W,&�ga�s�T��A��ߵ˚u�C2�2�E̫D̲�nȹ�z�����$�z�)��36�uW��1���s�[�V"9�]���^�=��{�6�#le-�5PnH�n�V�2���6�Ь�!�s�m=y�,�����2������]��8P��Da���}��}��k��|1̲�2��e>���pk�����A�IΙ��So �|}� ����r��疿gjʛ���eX">�ZfQbfU��8S��2!������H��j.��U﷌9�uր������=X�)���f�hE�ᱻ�z�0��"�Ne�d�iN0;����=�O7��)eI�17��U�#z��,�̫Ds(�̸E

����u�9Ϸdhޞյ�xP��Da� B�"d�i�]����wd�l�@H�v}`F�F�ѻ5q�au�`���#q7�1�����yUq����#vL��|�j�ۢ�3=P9qf�EiJsu$�F�4H-�0��%B�Ekk��e�qF��_���ճ��07dǣۤVu��W�]q���V����y�x�~�Nh��,X'�ݐ@��|Dݟ�O9fX�3���C�"�O;�eյö(U�2	��0#�Hu��}�6��H0�� wO��ѻ$vf�oޱ���	{�o����EW;d�ݓ����Jqe�q�c��#��#ϧ�n�w:��n�*=0q33U>�@��M�ۺ}w[j��Z!FT�a���T�*Jr�:�� �=�^}3�=w�1�	�.�۵��95</gY�B���՛�{��9�	 M}�����A;����i�0|-8��׿�ckݸ<�+�T�]�ÆЫ�g�x�L���%D3,ώ9���ֳԉ���h�j��l�bܬ+v�YUm8�@;v�I���"���ͳ[ſ�z����2�Dq�ϻܽ��W;֮߯K� �fG_�Ɂ��
������q>�eZo���:��>�<����޳f���wԷ)ю3&���::=�O�2��]��}����n7��c�����шZP���'~���x��y0�.�k}߳�S��Y�0�PΧ2����>��"�f�j�-=v"*.@�7>�rc۲�ӕ(�u�\�pA�#�AM;�;>�o��Cy[ݢ�2�̩y���ju���>��Ae>�Kr��q32j}�;��Dݓ��;^����YeԪC	'j\)M�:���1�d���z�Nڧ6�� �j�r�w���0zȃ�¬b����s�~{���I�;g�o���%W%�ڦem�jkJq�Qe�Iy��\Lm�0u��h4&D��T�j��tP#1R�`�m�ͱr�p$�[6L�,c2\����m����*������#
hl����2P�]��s��9�	v��K1H�%�2��M����v���$a����q�]*�d �E4c(�"��+��ؔ�i�E�ҹp�j�c�:#�Pq]�2�S���?[�c[FL�9�LK�ȥ��knWZ�JnvB�JHR�^�>���r��~7d��P���Y��0E���K�CF8q|3�C���F�#vA��|��A��٣D;��#vA�zr��N�U˫�p"=�Ϗ�vyh4ϫ4��0�`_I�_�0Z�����՛x8ӽT�}Ks��uF'S&��DwH"j �ݓ� Zs-,5<����i��~B���-Xk����<\�{qC&zB�"8�6k~��Vx�ղ��ߎ&�V1;�X�U� ��,�V/���w��H#��=��$r��Q�ysVH5#�v�"�|cvO�n��nC*MQ�+)�����e����k���4�\������Չ6Xm�[c�5��:|���A7d��싹ޯ���VOQ��s&��w��N�&-m�)ӈe�	�i̴��Zq������؂�b:�Uq�Lc�f/Hdܨ-iS.i�^��m6����wBA��k�B�?�hΥ{o�_,�R(��̮f�9v�$!s�O���C����o�����\.�����@������"��l�6w��e��V��h���e��`G�vD�e��Y��둧5f�׬`�(,3���fQbfU��멩�{��� @�A�>�nȻ�T��깞�9�&MO�t����q��O�|��h��(�3.�̠������/�N_���L��^o
b��h��>s�pF�-3*�&e��V�5�˽w������=�� n ?gC�"���XL���K�-9af���Q�9��[��٠!�F�n�>��r��"�R4��k�
	$ \��"�� 76 n�"2҆��������.�P�x�m5]�-;��3��d�����ѻ.;���ǽ��wv\�h/2�2�ٖn��}���]Fkt�Lӥ�d;���A6{z؛NS/c�W;A��͉��7����֗�\ ��꽆Oc��g���2c���[Y1��� �/���\+�Z�XY���1��w�,2�fe�J�	v�"7�����`���������ȧ5D�\��`m|]veL�˨9O�ȿ@��"=�`n��.��r[����O��o(�2hV�"�������/BҰ}E/�%5IG锚��+B�f�����ݐ��5.����Ħ�ۦ]Mٶ,<��z�f�>_�ǿw�t�����r��
�U]h#"xHS©�o����n����Q�Z�`��/�v#-����A���A���T����u�"��5>nG@�� �ݛd5��e�k�erÎ|T�*�L�-1�
��FUj��Qa����5��徹�+k^T��Ⱦ|�g(�2���3>�>���{�gj��ѮH�t����h��~5u����$@��`*�A'3'l�f˒���7�]uo�t���l��p0}}�#��v����VG^�A�"���@L��UÔBP��)P0��/1ӛ.��k_s�$��{?&�̳=e���|#�}�5�ǲ��슿����R,�e�B�����֬�x�}�,Fۖ�U��s�g�������8X��� 惺��m���P��$�m��ֱ�C3Q�ʶf�����~l��07d����-S���-f��()��{Q�}l���&=� �ݐcvA��!��κ�k"���TWI��Et>CY��`��#&}��J;�&e��;��m�e��uh�ޡ��?1i�9�/�Z����~vkZ���ޢ�fv�eZ&e��� �I���n�b�?wU�xy��k�>8�ܜ��e��8���S݅>�z����>�g�6&e˙�X�ec3*�9jV�S���qˇ3�8v@7u�FD�wO�2�ߧ۲,N����U�P���'z���x�� ���w��x����_n�{e5���M�uc��|�klc"�f�/�؝M��Kg:�*��b�as��o������m��a.s��q��

g�A��y˛�fd{��$vy�壐�;*jﴟU<��k�>�=u��z�e��!�{�eM��^�N�z�na�!���5�Pk!��e�&`>
zo���e0���M3���F��1ү��Mw���>�s��s�^�����p���Wٛ�|���{�mo=�e����.��9��H�����p
4N��m�������(ю�3x�ի*�Y�ֆq!��Ժz�U"��n�\t����Sb�*Q�"���ַ��5�=sUYt��a8YD5�n��
j��&X���'��7��݃�����a��?wwz\�ȍ�I)L����ۘʴ�e�h�{��yE�d�H�kaN��6o�<�3����"�U�a��˞�@��s'�E`��Уf-���+TT��Vj��������<�a��}9���íd��&6�Ǟὢ��0u�C}_K��}��t���vb�����춧H��P��-�/GM�3�p�@u����n������ElH9["��ӹ�+�R�e�7Ue\�����Ӥ�s}�Y�9�7�g���b8d��Eڣ8��A���j~^��h��֦�P"��@'�U���u@Y�nQڈLoS~Y��`�1�]I/r��)�����
������792כ:��])�93P�3BN@�H!���g8�[o�%{��ץd�II6�f8�&�����9�iYif���J��k#�C�zբ�{n�99�98����83;;�yy�\�<�۰@J:A� �p�6�NW�s�ՙs�vt��"�۰fQKڲQAyدl�r{bB���&Z ���Dqp�]�6g'�N�2���;kH�ڲ";S9�=��f�Ӊ�����9Gמ����g`�=�{��8���=�_{S�H�m�Z��#�Þ��s�X8e�h�76K;&gcc��,���H�%�uﾬ�Țζ�Fۭ�rq$fAIM��&ݧ(���x��r��3E�9�h���"F��qə$"	�su�Yo,$y��o�@ON�D��L�m�ٍ�;��w�����6��p�m#��I��BJJe!E*�T�TP��쿎�k�gX˰�4j4N��kn;Z���H��H�-�*Ɛػ��*l�]1i9��LU&�唹�lc1�(��ڃa�B�K4����݄��m�чn7j�Ƥb�K�֩3������,y�*�F`�z�Ԙ�)�(c�a�۲B���0gL���.r�mF�(�3N��Y��)-Lq�����[sf2�d&�,SY�i`Q��w50�Ԭ-H��l\�؇g+k5l\#�l�4k+QB.�{�f۶��k5jhDsA��F�Ej�C�D��-z��Ѡ2�h�5�Tk�K	�mMf-2��)^ \Wl�j��KC:�f0��]�l�XݯZ��\�al-�憧 ���%m�w�m�(j�%\��Y�ƛ5�f�0�4 isqM�Q�bX�lt:k�.�q(����̳c"���j��e1�IX�&t5f��1����D/jBۙ�e5�,t3%{gF+��F��lĴ]��4���P�ҷ��<���-�),���g!�3k�b�&#u�a�b[�^Te0U
P�L� 5�ƨ0��TKF�&�d;i`�#k��75��Xi�F�� ]�[h�[S,V���ņ��b�s����I��6rUζ�B,u\(�4�ե�Fږ��2�A!�m�j]L�ejXH��BY�2К�i4�4J�#S�A���i�������iy��$McE��ݦ K-\e��'h�6Ę��qD�l]j6[�ְ̈́�1mwR�֎��m���\���ո�l^Xf��1R���2]�\�2����5���i�&5��Vh���� 4�@�"��!m�J(0�e���;DR�q��5ix���M�[����ʶB°ƹ��"��uQM�Ne{F	��	���U�Z��XR�$�p1l��k2[Ha�]Y����؋� [:��˱2lB����"�e�b*,���TjP���s�Fd[��tmqa��0�R�:�FV9⼶�*B���|������Q��ӧt�Ȳ�GPQ6��Dؘ8���.0ɡ�sn�нY��E�n�:/X�[d�*F�%�a4�1%m����.J=t�&m�1,��������̰vW6�X���.5��J�����vݬ%� ��r�ٚ���x�x/�y����
V.J.2Zѷl�n�ɱ�T�X��Ḻ��D���\�;{,���@�V5й�vt%����gF9��������K�qs���h[��
�R�Ki[b�X��V��c���zuQ��z����ʴ\q��{��lB���vEUU�M�F��޹�#���jŃ(�i����WK�V0Ϡ�vZ����[���d��@��F실�^$��ݽ�m����<��3�,c�PXeb[�V��Fl�顉�b�������HȘ#�Lr�li�n�1�>�f��b��� G�gM��ط�`���n��Z�Z��}�-6�=[���Rh{�b9�X��ЎeZ32�Ls�����{�d㊙�oi���VO�!"nɁ���V��nftR�k=��E@��6�%�Ff��bM���%����6îËk�1AZ�kV3���%��3(�>��v��/�ïn����E���B	X0sX�Q��2����>���γV�ֻϚ��+K����f���a����=�G���t�sC�[V�g����hlN�m�ǚ�Bt!266�E~� 	�Ϥ���[�&~�/�۳qU �";�ˀDnʽ��/yu�P�D`H��7Hs��Kv�89��%W�f���;|1���������`���,i���L��QwH>���"9O�� �C���9d�U։���D�1���,@�F}�e��b#�2�,�̫;��o���4#c#wt�x#e�;vn*����@��1`���-Y#�� Oۛ�np�����&�˙E��R,+����+4ԚYkh�YJ�[M^�U���ϺTߪ�s���Q̲��w��bj�k��w���.p��5�"80�zBR���2�����o��O�E��wdh�rD\A�w �-��"E^�O�{�@��`@�A�n�T��R��}ۙ��'{V"�X�U�&ei��n��L��L�1/�sT�����-��݌��6b� �I�t��vj�]�W	��M�.�gP��f��y���u_As��q&p�'Ti���{o:L���+k�Z����>��;E��h�Yc3.ͥ�q�>\4����v\A�v�F�]�T]�&��u��W==�L�P�Mkܯ�׳�ޫߪ�3(�̢�=���D���ˈ3'�s�q��t�ƽ���|��Q��^���w̹��퟿}��}��z
Lcv�
���cUf�H�b��bmiu���rkn,R�ӛ�տ8�={��A�A���7d�}ѧ�D�{�̻�����sۭo�z��F?z�r�D�X�}i���m��D��N�v1�S��f�W;��j�9]q�-��@�@�j�~��m=Q;�\�Q�#6 u� F9`��B҆Zs�$iy��rL���fx�x:~��M׬^��Fo,�fYq-X���~�Oj㕟�X��-�}zrc\�O2��k��@����:���۵g{e棤MH��ެ"��C�5y�U�[V������G�u�����o�����w�%��T]^׽���n�����G�3.X�yV��[7\�S�z*U����� ��3�E��&��a�ws� @���v}p7e͉�r�����]-�h����r��C$�+6̷֬9]�*��JD�uE��6��|���/_�H��"�}WJ��+�EE���O�O~e���C��\L�-̫Lʱ���g6c�g�&g�%�@ޚ}{ �)\��X5"����F�7e�sn���^7�.3��|�2��3*^e�O��Å�l�:��T����d;=���=��S2�3*���f{�e=��[���{ �9Ɂt�-�K����"����&GGt�\�ۭ�{��ċ�?/���b���J��-_Z{�����tv #�RP�a�{���5"���!t�c\�vn{t�k�f,�����n��n�ٜ��y���8s'�Yo���7��?��3fY29�w=�{�I"X����\�Ș�o�v(U�R�����=~�=I�������b�S6�i�����5͈��t��-�
A�T]26Z�a5`Yq�m��&��Fm��un�F�!������\�CD�c*����X��B��n�i�4��hg�f���Ûs��A�]����0�B�Y����r��6�[�FkiAճK���8���p�R����z��`mB�����]
Q�fYp壚(��~~-?Q��Y[m�60ˠj�L�uuFذ,lY�-��l{@�����ocۧ�ѺA�U�34�=��]�5��zƑW��ק�����,@��c�Lʙ�|9��;����*���b > �M.�K8VtEE���O";����n�����!�|������ݟ@ݙ�B/�Q��t!��o9�E�߬\�C�������n��|:ܭ}��b��=�X� �*����$�lN[���;���]�5M�;���o*�2�\�,F9�X�V�z��S�6Avkjmv����q>����`F�=�G��d'���C�̇�א��ġ6bg3B&KA��&ڔ/Z��D1�)\����֩��7Q�]z��*��Qps*�< n�'x`�Ej�R*��.NN����<w7GϨ���̸f|X�ݒ N���y�d���G6�Uf�?0U��G}f���]YӴ��&�WПn���7c%�n4������+��"���]X�����3��}���}��"��k~��I5ےm��t�1�/,B�Dǿ��߱qx3�Ń�`�X-?ZqiΈ��3��� wz}��񪯹�Su��}Ꙕ|̩s2�e|���]7�;u�3>�������z4�GM)Z��,�U���A�i���:�N�Tp��V��fYs2�2�nΜ]Fvq��A��3���I�}�6�O�L�A����٘i\��>o���|��F�ICH�1\�ViiF�.�0�2ڨW�GP+�Z�Qݍ�6��M?lЁ���͓vA��qv��TLZ��d�>n���ji���2|1_��n�cvL��0���>�ٮ�̱�*� s�+�4�Úr�WlX5 ��A F�E��!��������X2ӈ}j_�0NG�CJ`t�]������(H^_��0{��������zl�o��9}�_c͘���z�{��Y9Uv���*�Ȫ����z�0�wcM������������nfT�����dV�w\��9�:2�r@��])r�\��&-\HȞ���"D��%�Q�N=���e��q㍂fQn�d���&n�7!�y���r���H��DG)a��ݓvEI�u������,�T��,ĺ��Wm��mˣ�C\�"���n6l�j�^�U���9�r�#3���#t� V�G��.$�[4]T�v�^q���i�D�\�Wȸ�3>�1̢�ɑ�24��B� fȵҗ+;�/F���?~�C'�+�8A�a���w,�7W�y�X�U�8���W���S�^��r��cA�\�� ��.G2�2�Lq+�v�}���ϫ�Ԏ���O�d�2'��O-�.�z=� �$չ@�h�oƱ�}gu�����$<��W'�'<|�t>�\���!l��m�{�%��񏗺vv��N�2��X�~��;h\gI�A��|�ݐ��3g�b���5���H;�)s��FgT�q#&{� B�"��؏F�_W_tu8����D	�d]4,z�aj܏%V�pҋ��V�[3�c�p�*%���}�^Dw�X���2���Y�}�y��r�Vv��k�UnZ��HA�(艿�[ܩp̰̯�2����K���3o�p+$�G��
ܩ�]�TI�H�:��wH0 r �ݙS��§�^��kI�ˢ�{�X��&eKs*�=�B��8(Qu5�*����5��ūh�T�<�K7�X��lL�,s*�Vs���zlnV��8F��ݐE�99��zt�툭�k��j��eלE�N:����\LʴG2���\2��#�7��N�v�B����Ӫ��� �� F���쌞��H���9���U�D�kB���2���Ć��9&�sx��>�+��a�؜�x"������=��6{�67���@��o�}�N}�z��)V��vݳm�en�X:,�B��.M6f�nܻ;�������t!m�v�s����,�m+H�gv�(66�[6�.����+�ں�1�KE��^�%�8T.�u�h�l�\�4#�*M�Tخ�hB]h1[b�[u���SmZ5&��V볉�*���D�\b�4�in�T9t�����|-�t��.%�;c���D�����~��:[�[�0ԥ���Dն+���U�v�le��5�f�q3lX|����0����nɁ n�k��n�r�Ψ1j��O�_�B8��c�a�ʍ���X�E$�n�Dnψ���:���7Ip3�F�� Dfȵ�n�3�����S�pA�P^v僙[�|����ָj��&��}�D̲�̫bfY��?k���q\�i��L���Ӫ���� �7d�F� n��0v�MOB槤�#���&��nW7r�FgTj�FL��@���R��`�;$Ӌ�P.�������i�2���%��O�Os���*p�o�)�+�Y�*v���ϐ���Ջr{.Q�	w:�H�t�
պX��T�p3�a�kb�hbVl�%,�(���/c���K��-3*�&e�N��W��蚓�#4�Oz�W9�3������e�r�"�PfQ�A���]Wu�k��g=8����3�y	x�E��*g�����CړW���N�����s�	�q8˷27�W�-I�qx�����z���D�"��|�p���1�j�L���}�`llr��)(�[L��kv[�U�8��̢�ʖ�gw\�/���v�k�ǦVg
��k���X��-̫��Yi�]��k��EK� R d+��vA��˙]���<�L��������n�շCn��!��_	N,E�Zk��Y?pw7$U��Kp��ū��H�]$',C(����V/~���g���Q�f3-�B70�c�)U����a���┰r�΁
^��5^��y�b3}��_D\q���|�5��ͬ�S���[����; I�>ʗ3,��.P��4����7Ͻ�^���@\-�G�H1[9fWv�U5ʥf��G������ѻ1#6�ʞw-�||�8�ʞ�	�%��q�=���h�׽�����T<_����_Q�L2fT�SS�E�R��M)�����^��=r�F����������ۤ�lE$ݹ�X0�Q�&)�4�`�����wP�_s�y�*l�-���lz���R�흢�؛�{5O�Bq�T:�m�v��j��$�����x:rp~D�<A��7�7Y|0bͪ��͹�t��a%;ǡm�*fx�S��,{/1���7@=��S�[s����U�s�R��>�X����{�U��%�I���?����9�S���;^�&��<!X�����5m����	��݇~�c�ǋc�3}�4n`����N��˫|�<5��|	M�=�b��CW_'��x���t��(�b���>�V�pw{�r34�ѷ����lQV�{������}�������lL���3F�X��9u-��{S�?^Y|T��.��ٔ9�x���q�����ȼ�=h�m^�l&���w��$n�9n7��[
�f��n���f�ɪ��U�,�ݯ�qŶ��l��AT��ݰ��N�q*.��(�<F������Z�C��|�Ƴ�2���4먝u�-�u:�÷0S&���9X�������;����'w��~�wx��/�}<wγ��4�k޸��ۀ0����[���3Svi�k+�GG�:�n�~����j��8���G��K�]�{��$ͺ*n�F^Pfu�à�&F�m��m�LQ�Zb���c��n������x���;n1�O���]�Vxg��r��S7�y�K�m�#��e�ێ<����v�fY�2m�����ޭ6Ŷgm���n�p������Ӝ�Lm�`��QV��ZNIÓ�;cv������ KkZ�b�L��^YZRQ{�^t�'���9�G$�6�۴�wfw��ݭn��8��N�m�����k9���f�m�m�:r��a,��,����kL���#���<�ӣ��4��g	��B3e����#��R��{j/��gd�9%�Y�ݎ�a���d������3t�V�M�������{[�{[;5���{�����.VnG1�1���J�8��kD���nكq�Ŧ��{{�o5l��t�kQ��,ƙ5��ݹ";*[w���R���$��rw/���q��$L���
i*�i���B�W���w�����>tm���U�f�e��Y�e�J���KEx&�gx��(JH"66nܞ����/O����Y$���o�~����@ݟ�J2U�ᖙ���q�|�_Vf���P�5ʥf���KS����B���8-^���'����^�$9�.��j���d0�t����c.���Đ��Qߴ����ZWx���௦6\�_{F�����������t��ʻWKgڑ�������/I��@էۮ��m���,�"���l����X�;�q>�H�뻕�=@��U(Ԟ� 5;�7t��ر�@����R�7d�J��௄��Ⱦ�콜�R��ř�j�W5�)h�b�`;���1�U��ۀZsqx��B��^N:�Y�[�D��`�ir��oj�ç�<�7��ݐ7t�vF돈7Wum��ws�S,g^-���7	���Yfe��{m��9�f��(��Eh�Z16��;8��X�� �rLM�`!��es��e��|��>�7�wH��٬1�}�5ʥ��q���p��Ĥ%;�F��n���|a�uv��5�9��m��|'Q�̛�ڨ����œ/`FR2�W����ל�)׷=Ћ�J#l9Y�V=�3|;dZwd�#wH��`�����A�����Ml�0��g�QF�����,�Qn���v�N[W���~gH��:vJF�n,�mjʞ
؝F�ro����S�� n�r|�dP魭��rWY�G#r^��|*���N{�ӽ��[�J�g?_=��N�dFB�&C��-�ffdl%!Yʯ�{����SL��4�,Zn噺�-P�:խ]Bu���isi��V[n�����.*X/n�te�:����ؖk4Il�� GL��M��+i��e䔖`eJ� Śm��F�Dm���h&��T,����ht܉X݅l���YL�p�+V���mK��̲�j���lm�*�+�7iE�K*��v&��.l�
������j�4_>}�@��n���e����FҺe�]�b�a�!B�;�77I��3O�s���O�mY�}�;��k&J��o̚��4��6I0Fr#\�۲7t�u*�	]B���u���^�����k�[������S�����:�!+����wwo۳��l1y�ҳq��Ql��ʾ����;����w�O ��2��~���8�Q���5��&�pʛ�ЁY1JՋR��F쁻��P3��u�`�,fɰq=@��ttԞ���ݯ�v�C˜���=W,.�k�a���ʦ�r�V[34q��v)�̉�"1Q"�w������9�i��Q|
�ʺ�PMOuq2���/+M�>���L>�ױ�j����۽_�-�����ƺw����3�� B�#*�V}r��Hj*�1jBP`��跺�˽���r��k~��诰C�F�Xd��ɪ��푺�K;x�n��+���%)#��cXr3�`���PsV�&z�5'�}��3��I<
�a���6��MvN�L�r��PUK*�.��CB���z2���i_�G�"��YV�8���(�m̋Z!8�Բ�ջsUg�'ۨ���SOTt��w8艞g�2�]�n����9P�aY�Mef�k,�b�bb��32FVv��)"H��{P_=`��ttԘٺ�^����7x��BH���K7��q�cR2g�4.�S��m��W<

�e^��7)(�s¨��K���~�BH�)�I�ˇ<_Iq��'�&��Q��h�晕��T�u�:����,$b����)*3f
y�q��W���M��VP̎�^���������{����˓w����vH�D$�RDEԕ3������Ju���Z"����n�5'�;� ��{�nQ��w�<�>I�I(�X�����;�.E�;ɳ9��A],�໏��D�eLШ�ZO~o��Q[�aɞf��8�H¤�j�-C/0,�u��b=P"�D��3��X|�>JG�Fi���2��A��j�JWNE�`f��m��$�	#���=�4Ƨ��-dU��|�ٞ�uHԞ�>>I�%�+m�H����/��$RD�8̙�����֙[�IƮx�˾�]���I$���%KɈ���3-m��SOv����\3W\d�������d����@�����5z7b�P^�duJ��.����^���=��ǃeUrq�y��W!��<��?e������|#��xV�O���I�$��}"��E�t�6�jŪnz1�*�<>!kJ�H��+����^�1k�z�@6=H�]�&�lK�J�
e��tS\��A��l��g���|��qI����+��t�,�gC�?^�����!$BRG�ד���aán�SuD�n�4�GoL.�@��5u�쑩$��*Ǳs��l�X|�!)	#�F����F�n����t�������)"�[���Ի���}�����+y�9�Q�J�̾��5�������H�H� $��"FZޭ�bS�^�<g-z�U�n�c����>ԒX��Vɚ,U�2��+^��.�*D9�
�wLҋ����/ճ;q�"�=<�}Kcs���i���j������[����:�����g��bnfH�RUJY��6�wSe�fk��(���i���-��2ג��k�h]�b��ZB�k*kW�f�:#-�,��@��,��-\-�� ķM�-Bŕ�n�m��E53�A�e���n���6��,�cVmAL3&K.a �$5^#��u�m���t�b����Yp�q�67b�<⹰�&] �1��"��es���m�6P������Z]Ff��o)c�0]�d`M��K�RlK�v��r.��R�B=S�y�@ޔ�	".�h��޹�#Ҫ����cMq�W���� $�SA�۞�=���)��[���َ����s��܄��pwO'"5���#7��H��$�4���*na-��V�7�]WxvN�|�#�H	"�M��Q��I]���j���n�\����jI[�f�Z��|�>JBH��In$3��j�V\��=�������|[Z�$�7�����|����[AHʵX�	�ተ��,v�[�4�8��6�EF#�1���~����t����1w��"O4&������~���4��q��>���$��H�Ae;0�2L���Le����Gi]>�(g�Z2ݪ��T"�kro�n�4I�&�w+k59ZQ�8��[3h��xl�������}kT��iU����l��Fjb�/GZ��J�]~I$��>ɬ�M�^��U�����d+���9����$�������;�h]�ˤ$�]��s���	�ȷU�윝�{�GT���q���$|D%))�S�4�ըL��3����u���<w��~	.�:�:��b���������,A��`�֑��VS�E�h0�ue[������(�?�}�?n��������y.�l��R���Υ�J7MFr�����J|Gj꣰�++LZǻቐ.m���f��9���ݒ�In�s�f"U�O%#��!��l��$}���z��������*�����_�My^�J8��ޥ7�ʟW�^_l�,�;�L��9=�����J�Yy�17O	��X5�;lUE��'�������Y�?��)O�G�,Ρ�����;]^��`	H��Ӽ��,���VVw���L�R�Ei�l�kG�JH�$�	KH�wY�k9�
L��X/TL�hNvE����d�H�$BSI�S|�=�f.��%^��k�M��Y�.�k{&��KX�Ff�[έ݂d��-HI$�v�����:�,��H�Z9+`�����|�IbS�]3�qV�ٕ�=��UvL��
�d�k
�f_ ���H��s3��Y	H��I+	,�;�Z]�H�Gy;7n&�$I%�%!$X��Y��T�_kl��H��p���v9ՙf�����-��t\ev��5�Eٻ�����pX��p����*��	D����b�y;�"�ى4�D��Bv�w^y8U<�f�b�� o���BH�#�"Y?jCAӰɿ��<5��և:�U�6�f_x>����r������ˡ$�;��R �Ӻ�;S"�L�Gc)�x]�m*b6�7Dk-�k��>����>JRDYy�:3�ڛ�k��=�d���yq�JBH��v"q�q�ٲi�g:�l!{���wf�����|�����:i=�|O��)"5l
���mJ�u�%���ER�+2�y�'!$|�>Jv���E�ESXIXՒ{GQ�hv�ݸ���/M���.6qGh�dI+	"����n�����4]�R7�نj�{�����I?	.!�.��ov�^�*��5�b��[W$����X7�����}��ާu�Ѭ�1$�����d?{{ðQ��ISCr]�,ݖ+\n)L�ѫ{��J�R���y���ax.�����Q��U�xw��li�
n�{�&N����K�����E��ERg���8OO��J�t�����_� ���׵�
��^��� fQ��t�Y*��^��=Gy��;}y�/���0ۯ �%��D�
&P;����޴������c�-ȸ�Hә���N6/"*B�\
�rh�'ҋx�q�Fp�u���w���w-k��m�XA-�"�n���F;047j����
*����,����y}�Ƣ�\^���o��������Z,^�q�%���2/w����%�f/D^[ǻݴ���E��zv�]��lo7Ψ|oNٞ���݅����N���J�
e���9��<�5�8��С ܜ��Ignj۫O^=�o�/�SL������ይ�7�ӭ�xFr#Rj(��w&u���۷�lr�tu����WxC���:�����h�7�r���֌���%��;�n��4���[#�� ��ƨ/��gnC����fn���h��u�����p{��Ʋ��1{C�o�G�ST�O��-t���<��������a�w��(W����ۅ:��wm�Y{XEua�Kǎ�z�ܗo�Zn�^�ל���:xo�ӻ$,瞯j�Gsw_}�n��g���}ks�z�¨�n�'�q�R����Ќ�l�Wlk�٢��6�L��.к�U�TNgh��,���9������������9"�"��r�;��d�K�Af�0익�G'����5�(���n�d$�!a$�fG�icg)@DA��$�m֔��)ƒ����!o{�{γq��8(9	�9�����׷n����)D��D�M����!�Xs�!���,�9[d�9N9^ݜI�����:6���.����[�C���'D���\���J��r�����;�)p�"e��鈢Ҳfs�@�� �8=�c����QD\%��ɖ��:ma��5�$BdZ99�l���ki�m��4�$�e��#h��y�6�.)��Ľ�:۷�l��ϱ�,̴�1)c"�W���ma��x�GM�F�"�캗aJ٭�Z���\B�A��Z��Ĺ\�.��&ekE�w 
."ׄ3��l�[�6e@�l:���Ղm�.��R+��Q����jQnNW�؆�VQ��r9�,1i{,s)��5���f��4����Y	cpX̽�K)*K��XJ����^X�畸��T*��Bed�S��c �Msb��.�5�Ѯj��3�:�u4�x�f���A"ka^F�Z\����-� h�e����+V��le@�`I����t��܉`�V8�/i4%M
�Kc��2͍
�Y����8�����J\ *M���A/��� ��j୶^(�	��UKm�e�:�ҵv�H1� <	m���1�٥ʱ���GJ��.4�[��k1����ek"�5�*B�1KibM�Q���V�y��ݳtk�KT���,m30�«1(�&vs��ij�('4��Z/k��-�k��a��c��y"52��Bi�B�
$������@��\��.�#H4c�Cmq�2TŘ!��:�A*���[s���� �����W�[���͢�bPZѤ&nt6��m�b-	��2��m�%��˭)�
���1��r���n��7O(���h,1;��@ƛMf+f�P!���E��c�W1�Sem�{3��(U����f]"av0/\�ka�2e*9�oc]�nH�ڬ�,͛;^V��%1*�#��̮�a����b��!�K�<�&����"����J�@s�ҡ�Y@R�b2���%�3hLe���э�!�s
�I�a�1�����#�LD�5��,�&.֦���`����Fc���Օ�5����2�R���s3[k��gB�4,�
 L�v�6Π��Ŵ���3]�	
�-0˔F�3�"d"D����fA%�W�MX����[x�JZny)��為��)ek�]L�L��6��Ι,�+������EnC#��ly�'�y��jA�uY��%z�i�&����9��WX$4kh��)�e�[@خoVQ��^ACB��y��V%.����0b�k-r��b֨V��1,�t�`�����3�� �,���30&8�IhT+
Kn˴,ks���V�1��`��]w�+a�j�
��[��{ky�[m�kBL�+�P�5(lS5�֣*��������y-�a�3�vXm��e��b�1٤�,�ڈ��Ԥ�$|��Sȕ��슥�jVe��_�Z9\�_H����!)	#��J�b�ܼ�7Y��{GQ�hv�չ���5"Kl������w6�v�. $��$�&��F��䱂��ݘf���Gk j��I���=o��_����"qpr��.R�/�q�&��j�8#Iq�݇5�~I$��4��n�̃���>j���K/GmѹsUº@Ԉ	"�WvT�7c[��"&H�QQ ۤ*ԍa�LQmmR�m�])�ĳBn��=n�r���|� �dR�#�#W\�E/�����3T]Ȩ
�7�@��$�H��O�ӵ�h;���U�}�.{�I��	��+{�-�k,h��7}���%�>^^b+��'U9�s7:!��1Nt�-ו2� ��y����0��vV�p�'!$�l��OFwbȦ�3�ϸ��"���J鬘Y8�/$�N���ٲ櫽]#ڑ	"<���"��8O^oUwiһ�X]4�+���]C5E��ތ��S}�Y�fNw��S��)%t:���ۈS�t�s��[�.enW�Br<� $��z!���o%Kq�"$ɃA�0jʖ-hdCi�4Mfc�qp�bQB٬kX�!���Y���%�XI��=�x���͗5\�U�s��u��W�$�����Z�Jɺ��<�W\�Es�#�˨f����;Y	X��yӉ�ާ�z@} $�H�$х������Ț�\RJ��;�oL��Ѯ+i]Q��D#K0���Ψ�~���)�*DS�� ��ɋ���J�p���8)̷����LGr��}�VG�)HZ�[�{�^v���$��2�����\��6\�w�� bb�HXxr�صJ���j����H��)IfX�bN�]����Њi)�e94k���ݬ�)�H���Y����B�*��� �XF#Gv��#�3pĄ�қ��SQ��&��Td��s>I��y8yÜ���Gr��]��U��u�<���$�$coqC6�]c��嗷:��f\�َ7Ş��m�S�ԏ�Jc���]��<>��>I�y7�i�Z�O�VsRy��Ѯ��=��J@I�'����e�sQ�-��Jz�	�xn���++�q�q��19M�f(b��b��Jm;0bYu����fH���M�ul-@�0�e�펺��C7�J��+%A��am�tؙ��]xՒ!8�g4�����$|D%f�D�V�H���+g��S=9dۊ��\�G�"Y�]�������`W��Z4����gah��ښ�Cb�<A�(TС1F&&��$���>j}�IU��#;���Ӛ�P5�@��yـnji-�^JB��	U3��G�O��	�{#xV�:��p��>jRY��v���Q>���}͟$��RG'����*��'�quj	�:�I%�$��Sզ�خW{@WK|BH����;�T�'�n��� `9���)�����ڒXI$�hfdTv��F��m9}u:��Qܮ]�\�$BK5�e�fJ����wB!��j,�樈2hǬL�q��njX��/��W����n�>3���j,�T�8wخIb�}H�p2l�B�G�k��Ÿ��ىV�m�
�a����3M(gl�E+c�3�G&�4A�����S8�F+0m3f�ð�9&�R�Cs��GWlC&bً1.�ix�,Ζ%!�&�m2�l;#c.\���z�\��1nke�酩{(0X�'3B[,3G.VV]B�*Y��,(Yv�����Տ6�6�ه^�BY������V2��1uֱý|��R��!�:VP�[�����I��7wkGc����͌T�\���4R�$�����=U\ﰋ����95�Uo�[>M�%>IFﮡ�5u�G6@��]g!:�Q�O6���� l�%S;�����Y�H	"�>K#��ޫY[OT�].�@찶w ���R�>I���ڪ���ոWO�H��,��UW>�ɻ�PO��%��b�J�H����� %!%F;"�Ҭ��4�5��\��;�th����sd%>I*��2	�E�Q��3@Lc��4�ґ�V�Ś-�٤yŴ�0�n��-������ n�I�<��s�մ������})e�г�zp�ܧ�!$BRH����{�s���Q�Z��0�����*���4f�s�V=�u/�E&5�P�G���<e[8�S)��b�D����*u��i[��#�e�ٞ�]�n.����s�H���Y��N�{\��F4|����Ia�2�&��[�z��t'{e���;��sd%!$BI�U'����{��<JEvOmC���i�9G�q�P:��vu��$��I!<�i�t�7=ݝè��U��uqwv���\�I%�k�Y2�l�����ty��wP�p�F�s�ŋJqY��VihK!&�=B������7�IDU�s��QН�jk�[��L�{o9	"G�O�=����O3v�M�d���1�]�]���{˸�RY�l�E�ݧ~��$�S�x(�Vz���5!nb�y�,V'Swp�rڠB��3׻i8|Q>ӔKc�����~��G�5���I��{{�����h���q+v�*&���U�Jg+m;�����\�D�	HIfU��������[��$j�9��棡;�,��{�������#i�y���܀��J|�IdLsc��.��ɻ�(y�]p2x^NQ��ܧ�#�$��x{{*��ցفɂ'S
Q5�h�[4t�6��E�foԷ����5��O����������կ:���A=�ܩ��L��z,e6BRH�%��F�p�v���u�u�wX؝Ű�VT���#�v:dͺm��H���ɵ�i��s�\�Ú��<����F����	"�Ј������]�F�2�lORy�vZ�G���h1S\A�l�����Rf"��[�M�˛��x���Bf�X����]����iA��WT,�w�*�T��!�7r�U��K�$R��;��S�ವ17��t'ye�����#� %!%���jvBm
/1�+��JK,i[�4�0.�n6KXB������&I�1s֧ʹ���tuvuo\Laᑄ�0B���@Z����%���L�N>R;����=�=K����Z�7�r1$�i�ب��%Mk1w�s�>����I<�x��j�p*�v��ICR�2�Ԟ����JG�I,�yT�kY"��%"�����=�.g�'S��T��ou�k!)�H��K)l�˶t�Cr6�lK��[f�Y�/��8�	"Kkmwp�єΛ�wr+i��O�������k��=��;�/?z���o�1-}?{10G)��+p��f���O<S��Z	`>�b�6{�Z��i����,΀��]]����b�Lb#���nԛԱs��f��$����O#7+������[DV��:m���g�ĳI���Bvk�K-k��3�k��6�!,����� ��M\�jA�� έ͌j�� ��M���-�E�D4*0I^����	e�1�8Mi��5j"��l�$V�׃f����ͱ&��!tt!S�A��ð�]aZ/���~�O�t�:V\"5��,����i`ȭ�C!�c
��z�|���=�~$�����b��Q�X��JS���X��_R<�)#�o7MN;���ԋ�ӣ���p�8x\a=����[�,cj�ڷ�<� $�J|�������:=�9�Lm�,���5"�>	JH���[��sY���[I��I���<��R�V(2{Ϻ%Q�s�K<��$�;	syO.r�\�fOՙ]�"���{˸�ܥ$|�j�P�<��ɢC ��t�.�n&�$]M�Ֆ�x2uM��;]$�}���IXI<g�'�ͩ����Sӳz�	���g�JH��t���W��Z������S��;S��o�'| ,��"I�F)��@	�0'H�s/j���Q�%15vZ���J��+�ƆD!���`���"���ɨ��eb�'�}�6BZ��:������ý!$BH�,��i�yq)MOd�{W��dfO|y$��$R�k�7Q!m�4����Cs��/Y�M��#E���9H�$���y�u���5HI�!)%������)u�N���JD�b�'�� &�R��h�Bo��*"��	k�J.�I��˨f�A�va�:T ��T�V���D�hL{9y\��>I�����vs�d\���و��뢶�X���"S��"ba�ʨ=l��r�T0�����E����>Q����t�E%��u�E������J���.������f�E�����B�"F*��[����UF�v�܍n�N�a�%����"�
F����4P�o��ٶ���Zy#+@�t�gzv'F�x_[��[<��S��V0V�!^�sbܷ��h�ݍ�
�_m=��c����Ѽ���!�/_[���D�v��z|
fb���f�{x����G{�&��т�mf�{"<��Wy�Д��� ��P��t?{7]�g��>W-^���I�[�h���_7����F�XBEƋ�1�\�C�H���&�GM{�����<O��[�c-<����.���s�1Մ���.��y��W�G�3�����x�<��B�ۊ��U���t�\w�O	�t �,�6���Q;��N�:e�6�f�a�|2l��p�*������c҇���y���ٝr=]_��x,�z\!�Y���}H#��=I�{@#�;ھ�m��vI=��|4�k��z�3�H��/m�*���f����L���֨�U�[���iP�X������tx{��UOY�ܢ��5�ZS����9�FS�t�Z7[�t�	.3
S�L9|_�w�q�h�z�}��k����ܛ�@h\�Vuc0@*\�j�6F[u�)b���͸3���B�n)������S wp��^p!�ھ��p��W�Q�pn�h�Ȼج8��w�^��	0����؄�W��o�����VƳi�Q�\��A�ײ�OK�|�`�ɣ�J�.R�ͻ)��䖶�̵e��m��:B���Yg��;�������C��m�l���R�$���۹+,����H�G)K�tp����}�{g`r"f�	3K2+�������^i�E�}�����5���o(�p�Np>����f쳬�s��K�"���"3[[�//z��yX���g��X�3��}�����{����qe�D��پמ�-�;o��yi ��R�m�
p(�H[n.D���+;�y��i{_{I����mbs���-��W�$�{ק{ܝ��'kRϽ�t�ح���N%8G$�ҷy��KڋG9�8':@�m�y�7��yE�3k��)H󛬕������%���)�m
�3��l�s���.�Y�d�}��J@I��Q|�nBӕ��Ϭ�ϒ�]�\fw�<6�h��>Ҡ�΢X��4��JRG�"���\c�����'���; ���O�ԈI��U���������zE	��V�̺se��6VUq)+�i�C^�4�1�s�'����ߛ oH	"H�\�����J��2y�2'�V�\���z�s�	#� V�}u�x��U����;e��C�L��;G�9����1C]���;��	"�����T�ؗ��� ��O{���Ԓ�%!$F�)��&��NL^�`r��$}ur�1+�D�̓'��ك��H �lNjI���K���C"�b�Oȧ��SZǸ��}��ޣ����<3�j�;6��ޅ��+�<���������$��C-lr��*�� �r����F��˝�����BH�jF���!Ļ�ާ�=|�<�~�������ٍ�!R��l4�fCu�ĊS��D�&�*�Ԛ"r:�K\R�DvdE�؞q���j���F�F�dU�@VY���	"&��m=�"�=dY���"�QҊ��2{�}�̤�I�y�/����+��I�6���٬q:q1������Ƚ����}�BI%�)���VwѹYP�-"��%}�{"y���~��w��S��mT�鎮�d{��$|�>I%]&��478	%�υ�at"��L��� .i_�CWT��I��l�#I�5=JJ%�i%5&�Nf�f6��e��AP��^W&x�B���ntb�1���>�>FQ��:l�RҸb:�A�u���۪�V\T&s�i�R����FPl]m"���Sfm�X��iT�W;.���Db�1��a�Z\����Cl1���,V1�Ys��bͥԚ�����űbnk2�I������H�e��=�.��lKk��
�L;0�sA�%�9��Th�rj[�kЉ��p�u ^%H�F�m�5�`�@v[�ڃ���~��<�ccR�)`łTݍ�X1�Dq�%�p9)X���E0jH������%"���¯�=1�j���(�/)�vg_e ��i"��>��1Qq��:謟�G��&�lO8�]�|N�It�CiT���6�e���BRG�	.q=2��千����#x.�*�$��q�J}�I�Văz�/՚sQJ�C�W�����j��]Ǭ0E����niW}H��ҿ$��D%x܃��R��Dչ�+"{���~��w�>���Y�Z��UW7�y5=J�n@��ae��w$�,3M�nє[ck����"	��EH�2[Z�JH��"��>�!0�0��I��uB�1}�����6��$BH�%�XU!et��*:.]��l4�8�u0�i{闶�6��V2����j��-��+y�6�˗���~����ߪorM~���ʣ�=����E���\�]>��e��B7�Z��>�܄�7fS�����eφ�|�>J|��Wx���X3nd��s���Ub���j)"<�J�'�v����r>I]�=��j�'n�L��|@��Wz&�J�2@z�H���$|��/v㜎�*��g����Q�"2�Ox>���J���Ż��ov��{4A$nha�^�CG�kڌ[6���X˩�h��TLu�{�~z~}���H�>nf�lJ�W��V*��ڸK��ԍQ]U��	HI��F-�+C�K�]\A��#P��v�$�����Y[U�M�).W�0���y$���^�~[�����Os5�����~>��I޿�m�ô	�vO/!Y(��g��>����,�7%���h��QÆ���
��h��
�{�I�{�GTF^��}���H��)4E�^���+���F�l�Į}Q�5b���D�5OeК��t�gHפoHI�	$���i5��':�VDS|��N��=����	O�A\�*��jxڂ��pKYH���b���շ(ЭM��-��fK��.��`�M	��߃�w�I%~���}�kw�L+��x�j0M.�:�w��RQ����������7}g��W�U���bE%YK�q~��h�-g�)	"H�t��Cz!�����;��d��|@m����K�{p�k��xwY	O��t>�;��&���<�0�S�T
"e�l�lˇy4.U�x%ޣ�we5khߣC�����g�twe/�ʶ�%�����dS��%זK���,������W��)MA�ܾ�wP�+a|; �X��y��bE$|�X�4{���bbA53"&�"D�YV�͹uqFZ��ۅZL'ZV`8�]���o���O���%`$�����s�M_{XL�����p��F�@_s�|� ����W����������/��@Y�W�|�>��~�����	��.�TO����P ���N��~y����6,DL��DVQ���� mЯCrD�~�s}�_�u�0�}tU��$���3>�>�||t*n�zd�B}q9�q1}SM_�|}���^����wk>'6������}�����2�G�eFޱގS�5: 6�P�nL���U�j".�T��~����糹�|$"��T~���P#���Q�َ��r��(g����v�Y;���_t^��}����w��*�If*�?����S!������r��O8�׺ 3`҉kPb���_g�Bхe#����v���3Xe�.�nD&�@����
���n�[�qJh�tu:���,�Y��Ō��r�d�&6+Wvqᰵуq���Q�M��E�L��R��m�l��h�����ZXnHW$���m��3�̕ى�K
�ݒ�A!�#+X�u��
	��*�kk�v� �%\G:�\��Fٸ�V��.`KQ��]\�6�8���y����~�Śݣ��٭+p�
�ZZ5�nX�b��)1�,�#�\�g���^�(@��EnH!�C>ٛ?l;�e��MT����X߾�7�:�Xh�;�[�+� �ClЁ�5��BQ��tl�?�ށ����~{�tMl�sNI�k�#���(@��P����C~�>�G7B�龜t(@mЯ@��SX�?nQx�w>_	��U�����m�P�٨�T>�����2�L�c����B���0#ͺ��8~Q�lgg�T��/>���D��ޭ�Ǔ�g~��o�z<� �m�Cl��d�8�U��VX��#��ٟ���4��rO_|E�]^npۡ�\��߿��~�����6{j1&�ce%�XF$<�q4�&Sv��������%�b}�����Y������o;~�_dn|�0w�>���:2����V\�m���٨�Dzd��×���af!H<�����+��>����I�n�E*zd�@�;]� ��,�����-��2��'!L�f���r�b�p�������ϩO}�������^}B#龜	�*l;�:F��QGwP���� ��P"d���y��M4tmϏ�7��eR�9�$�|�� W.�P����
n�C��75���g��/����uW��o3���6����]�������	��׻���-fq��߸� G���6ȡt*���zl}tF-Q8�O}����4f�xG���@��B�6�����}����"�����5@D�I�FR��-�&�V�̲kB*a��nBmhJa�M���� G�3��0�4#ͳB�韞���)�朓�5�#}��<���0d�=�Aܘ	"(@H��w^���v��!�3:�^���/3����}0�P��������!�rz>}2�$}zh�"4�ۯ7>m�����*4�*EU�j~Gу�a�W݊{���ltt���5b���.{7�<��lo-�cJ���V]A���� Aoi�D��Ũ���z�z>�LmС�}M�a�h�ڥ(��߹�]������5{�έ�S�V�M|*�"w|E�o3"���n�������CrDmШ���G�
蒣��H���+k��|�B.�*�ށ;�>������m�9Q'����}����~|���xai ^�����i-!l���V��M���:�b�.&:����}���,����!�0dVv����}�?�&���/>�`�qy4�I�n�����>��f�@����s���#7�d|8B�5=.4/:gV��Tݩ�+r��R>��+�P�nI��)� Gٔ+�ϫ�";�0 6�����:^}���˴ܽ���\<B,����#���;��g< D6��E��ыX2���sć�"�wO�n�}�?ei�'�ۓfo�^}B}����ߪ�����h������H�+&�Y}[�*��80f�� vf��s͟�����������^�T���39��U����p-*�C����!�j�"e��kʘ�h8{F��ҷ��9j~�ܩ��W����{�P�nL���EO���57���cL���5�0m6����MX��	X��������R&��cҨ@�}����@m�7#=w�O�]��ɋjc�����'�ƃu��7 ���� Cl��Ͳ��υK�k�}����fv�������nN��f}�}'�#ɺ 6�Rfc�a�ΐc7Mzi���6�@���gL|�}���kTrԼ�ʚ�U�"!��P��ȯCr`@m����H$����P!|�����`U�O�]�\������]�#�����L��^�h">Ϗ�>���l����nU;#��l5dc{��/���rp��#3�B<#���
�۠+���@{�z�w�y��?Y��wu�y0����n]���| ˾K���	k��Ph�pU^d�ꉕe�!�'�cH"ɿv���	{�@��M��}F�Ɠ�r���y����e��0\�Yv�=���d�Tƥ��kQ�����n��wr��<w}�3I�vv������Z3T����_a��^"�o�Xq㽱�)��o`w��/j=�/x��yo`��+rK��?f�/(C]�$M&/�`��,��y>��z˹�s��s`l��$Ǉ��p�R��Χ���
3�m�7��ɼd~�kO=�Wއ��e�r�PB�[@��+��=]�g)�9��R]f�w����4�OO��C*K�N�˻�kC'�ɮ���.��5{�gOp�K�m�l���e^���xH�F�t�o-}�+��^��&���#����{�m)����""��^��^>�q��79=�L�4��<'3�{�O� t<}�(֤FR�Ǥ�+1�/x�ӏ���vLc��E�X�]d�,����c9��d�;�k��k�'ǌZ��}���N�'vܢ���z��2��w�ey�Z�sҧ.LZ���z4F�Cg�xfx⟳�^bL�*Vњ�Xo�e�D����/o92��ٳ�H^�Z����r�S0�bsNT��gd���t�o�W}⮒<F�����7n�x��:���=�i���8o.�^oQ��8j^u	�F��	�V3u��tJ���� �j�#���[����PE��w۸;��y�T��B����	�  ����	��?%�����JRW�p^ZW�{7a�9���b���-Jt%�hq\��ڛ�Idbm[�����k戣-���Pd�w�m3rw����l�r9(�Ĝ��ۋ�׶�rw���s<��i&�^���X�AfJr��б�yzb�j����=�"R���<m[޲��^c�O
���������v�b����D�e�L�0��e���!N�1�^�m�.{^�m��^�����GG/Lvٵ��ٸKtȾZ�|�ڳ�yi��j �"��4�	m�AI,�-�P*KEh���e-��m����[�Üe�(�Zf#�f���$=���n�+���׶^�s0��/�wƲ��|�З���9�w�ݞ_2(M�IHm{�S{���r1@j�`����](��[��b�ٌ����y拡491�ʥ�U��p�.
M�<m��5��fh][@���TΈbaHCZ�-��c��.���m.��a�e%����������v#��sb�k����<��%�@��`MB,�������v����*�21�X��,�"�\���^i[��� ��f�Wc�e�-cfBؗ�[ͥ��u�c�*����G��҉���L�±j�]"�.V�@�b2��e�԰ڛi�$u\V`��8�m�k��jL+eWEsYe���tkGS#y� ��k�,�4� j%��d���`d�cSKBT�V�P���P#�+�[Cb6�k#-&YKke�����]��Mo6��,ː�в�K���2��ٯX��q `�L�S��1`��J�\R��ə�E�G\D��&u���,!��!�6�ˬH�Ƃ�+�����fɘ���1��5�QYJb�K�M�	�ܐ���m4��"�pP��[C&U�f�[P�pZhd+����+U1e]a����=�1���lMvL��:�E��Ѐv�-ջ���Y���-xQf�2�E�)\�[����K��̳h��R�`Vl��&Ż6���RV�cb� 邲�Z�h۸�L��u4�^tj�k0�!�L�5��6�9��\���H֭�Ѵ��i5���KX�j*%Yb��d�õ
L�$�-�%Za,hƉՃ�7@��B!�Y��r�m֢XF����S$ Ƣ�5c�0J#)�.����*4.��Ғ(c�*F0�0Ի��Ҵ�EZ�X�[at�JZ�&�%�/<�J�C9����a���"���]- Ebe��j���n�`1��S�Ԃ�mspL�vr%�!0��d���`ƹй���J�+Rj��+f�Ɩʃ6i�݁R.��V뢺���ٜ	`�����j�R�u�]�q��mdrn�f5D�f�t�P3	����mH��*=Up�����v����K[s�XQJ�j�̮��t��mx�І1�ח��Y�,WF8����j�L����� �b�42T�Z��Wk��V��-�-�(�,�æE�bd���F��:�*�ͱ+�!6�U`��`m�F���ȂWLVؼ�;Q]�B�T�e��"�\�+��,�ioq6NZ+)W�Rkõm�^W��
�׌�ׅD�q�X%�[X�k�f3[-ne�0q�������`B��"�uFnk����hK��.�Q�&�J!�5U�w���=!�5<� �m�"f�yӥ.��r��*��_x����Y=ݦ��F|����> 6�P��"�7&���"z�;q�t��P53��5y�Q���������]�#��Bwa�~̠E�֯u���~�x��"=�t(Cs�t:�T�w�D�Vk=�8f�y���}'�#ɺ 6�
�y��5��bބ3*n돫QB|k�"f��N��_N]��Y���}��D���˫����բg��5�ECrD�����}�],�q����O卑�g��Fc���>�GwƠGqf�y�i��_	]���eo��L�թ��$�L�d�K�5 �m]If(gAv��VQ�M����>���nH�m�϶'�=�؉���7�/>��s����2��Fc�^5:�z �m��y�h@7k��ȜI�7?5�.�oG���Ӟ`|2->�h����B^Fi��z��l����M�?���*`�iA�����|:3�5�#S5y��_u�b�r����g�D}����P���}{����Ɨ�+�>�O���@�� ����v���w��m����F�9��t~����6�@��^��}=
��C�J�^��ȡ	ψmЬ�b~�G��?nN��^|(@��D	Q��O>���Z�g���(�P�Cdm��f�CdCl˱.RK��i�23�GWƃjw���[�`�˟��|G��Pܘ���|�+���~���Ȼ��)��a`�R�&#Pph]:]-T֕ՠ��%�r]�'��/K���}�������efw������T^�{+��7���0�Oa�c� 6��l��"�<3W��8��0��`'�W��'�{��G���9��ϨD}��z� ۜ�8+��N�����XAY��D>g���f�D6���|H��Xv�h�`�'����>q�d��]���/_ޟ��M@�j'�1M[w��n�٫��t�MF@��.��z�r�j�-y1[�?
?x����5=�h����g{����F�V�wc}��~� j�wo�����S��ϩ�\藱���@���S�RI��6Y��b/�Ё�q�y�"dW�Cn�nf�ll-϶"��T��P�s)��?nNτ^�}��	2+�u^��u���'��|����[��q�]VT��b�.���L�p��b3r���fZ}���,����Q2��h@�Cl�gȪ��iW���ܹ�Q��1P��<��j���;v�C�||ۡ^��>nr9�Ij��@U�@�A�Ͼ.��ϩ���^�����������Ɵ��~�g�@�H��� @mСϋn�X5�eb���,UU��Y^���E�� G�I�'B��}^�6�@���!�#�s;<���>�m������ʽ��N�����B�������nO���V*M��'�{�F��]�8oj5����N�!s�|Պ���ȯ��W.�!�C��nyx���aŌo�v��#��B��۪!�0 �
|��w ��ށ�A�}���ݟS5a	{#g�!����A�>���������������MSBj�KB�ʵ��"ⅶ�fF&� �B%�l<mM[�bW"q���78 @mС�8_�O��F��3W��}���������4e@����/���6Ϫf�d��]��
����ދ�4 D/�5���]��*��w.~~"?�"�G>�Pܹ�!MP��~C���z?��t�<ۡPg�"��3w��C��nU�x�5j"^����@����m��f���G�P�d�[��hG�#�@��
�rD���/�}����s2��{
}>���9'~�蟾@�y���s��ٯ@��"f/תּ��G���>�49��U���D�۟����+��P���ۡ��ĺy�6�����G(�H�bd�{=uz�8�#+QQ�v��+r�6�J"�S5l��u�>Eo���g2 p5�뢔<��>X��z����1����ѩ�Ж��V7eu���!��4`Ʋ�����Z�ں趶����A������j*�5���U�#vi�cT²ͦerj�KPx�d�s��g���@#��.&�!��%������&�t��ٶ�F�cq(#A#�6�{g���k3`�s3k2A���#���cQ�"�\��eZʴܭF�W4e�6n��j�����%�b����2�)ږ��:p]0Q��E%8��EȐ�R9�����K~�� _: 6�
�r�Ͼuo�ϋ4�"^���������ҏw&_�G2�S56�zd��� ����d�,�oS�C���
���/��?n��U|.�#龜��^�ۜ+�/|�H>�\k�"���d6��l�+�-i�q��R��H%j��s���"?�"�@��7&y�B�6�P�1����*}y�B?�
�r�ϗ�o��],����8~��[�o��t=�X���P��Ѐ�"!�E@��
����.����
�Å���\O۳��_���#�>�O�$Ȩ��z"��8>ߣ��?ɯ�+� �%���L��[�69Cj�u�x��Y�\�Y����4���1,���zF�5~�}�@@�m���ڮ���c�wj~~m�7_��)���z�_I 6�P�۪7$z>�U�q3���J��e�mk�xN�d��x&�<��;l8\�~f��ԙ�4i+8-Ս�+���Z����n�{�A�o�J����1SK[�|Z|�F��}o>럧]�y#�����P w6�4O�:>�#���>)�B��l�M�k�������Zk��������龜t(@mЯ@l��m������!�
�1�;���B�L��!�kכ9�w��e평ݩ�Y��|E@$��������BR}<��@@m������
�ۻ���l�X��2V���}�F���|������ �i� Cl�
�)�r~�y�xun��$�њ7st�4�ו[e�V�,iE���	��Ŀg���}��e��B�7&l�̈�_�����6v���w�
�MNVͬ��
\��[�+�9���D6�!�k�:��ݿi��o�?
w�����پ�����������"?�"��wW��_:����ΡB�P��n����ds�ݭ
����|�91�*9�/9��_Y�GC�Q+R�%H�J/�����%sc��:Q���vb�b�$�LM;�S�s�(�2��uuQZ������u����J-æ����8~������g G��h@nB޷�>���\֑�y��P����FfD|/����ٳ��_���G�O�jK8�\�9���W�y9�l��٨>m�k����f����-�����m؏�����G��P#�P�nO�6��Y;�g�&��b%�Y[�Jņ��E���t�IB�W6�ԁP��$��1HB���D|Ezn���{���v�*tl�8~��պ��Bz��w`�٨� Cl�3���u�����V}�k� C_P�ȏ����멿�6���{�z���0 �
��Y��ߏ���?H���y�Ƅ�dm�T6�}����.���M.6�G��������9�
ܐ @mШ�#���+�^� st(@���l�*��o3�}�:�?*���@���Ɉ���R�;ދ����M�p���ǧ{����=�3�޺RgU��Krg�M �,��'���ْ�v�7�A�.��f�{�Ƅψ�Cl��mЯCr�Xq��g~q�뮡^������o�̺�U�G�I�IС�}M�iȬ���p�3F���*"�T4�vԙ[1q@�6Ѷ��Lj3L�B�bZ~޳����ׄ�A�٠ D6�fl��_��1]�}jv~_1V�r�s���ӝQ�����s�#��B�6�P�nH���>D�����ܨW������+�������^|!}���6�[�{O۵^�.'~>�`>︊���nH���]<+Eb�s�x���*�u�ߨD}����Bl��dm�ˬ�EF_i�������Y�������۸��N��+��_|E@|�5	W_`��b3g��� ��P�ɀ� 6�M�騝�?Wz����_<9��BUN�~����||�9=�`{���Hʯ��N�e�_��]	����V��.oLh��-�Ԩ;*�Nl#�FeN�b(^<-��V�f�R�ѷ�;_'����Ȩ����0e��0䢪Ĕ�jS����z�l-�q ��͒�l`��u�4¢E���d-��CT�;jTи���\�s���;-�k1�ɞi��/e�s�J�;Q�VhneHp�R�kx�X5�a��0�#e&���Ǜ�����צ�]v���bX�F�.�`&Jf֖�d)u�SgLuUL�MPKv)6[�]�4��f�k]���� �Y�KS�iJ����f��6\�2�1��^�3�qm�TK��/���E��Ϗ�t+������9_
���>�Ҿ�2�@��P5}^�G� �l��٠
���ϫ����zGs5��}>�ͻ�����2�D/�"��wP�naf�~u[��cGb�BwB�t(@m�W�"�6�1�ݚ���9za}������� ������١m���!�����-���#� 6�P���}�~��3>�+�W�}}>��O�\�ɺ����}#!�hG�f�����;ݛܡ���	g�\�2��"�Q������(@��@Cs�۠s>��e��?�IA��!8_P$�z���������4I�=�ZZ�ۥ:~��м�X�zÜ��H	E�pJ�F�Tg�瀁��"y�t�~p��r���#ͳP>"6ȡ������������� �	���[5l+<-��1�Ѫc�ț����^T�x�?�~@�꿿Q���Io�����i��nlե1��Д���0p��O�\e�Õ¯~����ۡPs����IT��o��"9��Gs5��f�@�6�y�L�Sp�����olX�Q������.����B����ͺ����q�������@����� ������{�J��Oۘ}�/�5kcz�T��Eb�.C�5�DCl���!���#��h���Y�Э���2�؉ܯ���P�G�I 6�T�^nF���������̵��[ �9p�e��e@��v7V]��i����Ssrn������Dj�P#���l���5c7��_:齱B�Q�����^���a�iu|B{w�}'�l���
�nH>�0���aoDq�\�w:�zdZϾ������%t0� ��ƽ���uc�;�٨��̊#ͺ�s�����Ul�|�r��v51�2��;tCt�y5v[�^'gC�}��ɠ����80�!�~�>l���v�][��+)e�6�)�ܠЌ�E��x͙��W��	����NLf�;S���N�=�N��gk~�I�6b����6ξ*<�3�FRڙ�A��S�`3=��q�2G��Z�m�8l�g{ӆ��j�*��obq��F�EEE�����A1�%�sS����s����i��m���g.���p�x	́g���TT?+���B�GOpnk�wOd]��x�M��M�����n�4�>:r����lY��V����oˇ�e���{BS�&Q���Օ9���,`0�n�7��ݽ�!L^�57�*\G���|�ok}쇕}Y�pwi9�o��c5��� g�����y�iU1L��{��VvF������a��Mt"b2��E�2�����:Z��������A.2s嵦ۼ�X�d�Om{XٷY� �\�TC�gP���;�~���.xa��ۊSKL����	p�=2wf��.�[���c��Vf�+��ѷSd�m�!fS�`�P��}���������ލ�^r�3sn&3^R����:A��'KfDG��pGSdʸ��&m�꓆e�X�&[�)�前�6��<�ܬnu1+V�Lm��6!a�I����絍aoUQ�1��x�z�=(�$YJ���~>�ۚ�����u#O��E���#jL��J��mOD��ٝ�b~��s}pz�a��-��^K�K)Ar����)�Y�+u8�;;��Y_]#Rб��B�ad��J��l�F���H�<�w�q!;�ݵ���p��m��=��,���ekY0t��I"R5��9!�{F�k�y�N2�;����6���g��Ck^�� ��������bv�/4�;�i�=�^@tQ2��t���"_m�Im�tGwڵ��9/�Zt�ڲ𣓣y���6��7'Ͻ�Ok8��C�"Dr���������Ҏu��z�Y���Ӭ/m�����ݝ|�:m�_m���$�>b�Ͻ�&�Jq
�[W�h�f�ٯzk[Y$͔}��^�;۷}��+ӭ;k�E�����y��&h �B�,�y�l)p�S^z����ؼ��g,���{ޒK�y��̋t'Y��,�Ƕ��o{{��
�b���'�y�e����0�޿��z�G�I!�B�6�
�y�6�@�W�b�9�k1���}3Q�ٯX��~����B�Q��ʟk�>2��y���>�7W���N��4/{W;��Нnn&�z����>$M'<��g������oޏ/�>�> �lЁf���'s����zA�:i�ݣ��R�fYEf�le�ai�қT��m�1/��{{�_Y4���wߧ�dP���s��yTi���Mgԕ=A}���
���:�Cdm�#��5e�1�N�w�W��4 Drf���߾��/p]��l�2�".������nr鏲�U�D��^���(DwO�dd�
�6Bꉊ�?*y��f���3Kp��u=���@�_||�FCl��6��>��`o�"����B���$@��
�������叆�^��j��������\�4�(����r�̇7���C�Rb��e�>~��M�p��\�Q�{��{��ԯ�rM�T� �=�sỌp`e!'��1��{���f��܃�i,�b
�}����k��7�uг��F��+��|Eu
�������|���?��O�30�liZ�۶��.�`X����(�h\����u�6����������(@m׫�dn}��W�f��$ni�������	�-D�{��O�Bzf���Cl����9Yq�Ic�-�{����}����G{\&��P�G�I��B�6��|�vA���ݤ����Ё 6A�4 G��h�Q�2O^]e�n~���Q+0_B�����G�}����!�>��"�6�P�oM}y�޷>_i |�>��;���w�d�}�c��?@��mu/:��y�jd��n�z�����n ���	�M�
���>����4U�|&��B#龜ӡ^��>�6D��=�y�{�R+V;r���;Yi]��;�|l����W�iH��?n��vڗ7(�V��T��B����_c�o�%�O�����?z�=��� ͩU�W]�����d."ݎ�a�,�V��t�[��Q0l�HJ��-T4ѢX�wn�#[.l� � �j��m\*2���F�.-t�l%�i�(F���\�4���˅����t֏e����5������]B�L�5 &��H�Ҕ�i���ff:��:�:8�V=G,t�����PiWKq+�Z�r���\9�	���(�=��K���-�Ś�u�	��:�5�ҍ�Q]SU�٤�������_�~���l�D6�f�����+0WЧ'�u�#��~��²��OT�>��"�/��ۡ^�۪����z�𰢶���y�~�G�d^��ъ�>Yg����^�� �l��_ۖ+����_�|��
�mШnLm�z�*��5�+>�3��¶���U���`CN�@mЯCd!�h@X�P]��X��T�|��G�f��������M�WЦ��u#�_|Ex@�7�"�Do�tvI!/�P�ۡ^nH#ͺ��?��)�h�A�}�S�ȭj��]����>��A�5 `���������g�i�	�!�[m��p�%�ì�F�W�@�n��Ȕ�a7!��a����E���s��#ͺ0`��=?V|(輿�5��*3�+�<>��\���m �����f�ͳP+��ߑ3^���</���X(2�1�ɓ��,�n�V�)�[hܬlUQ������(��d]�o��lt�L;�{�{i�fr��~��L�n�g}dv���)��]|�_|E@o�+������Z��T(@������
u^�6G&���r�?M��}���A�l4S�����5qCl����r"�gG�ۚ����E@��ЯG�>-��>���?O�3�Z/+�&�">�L��5&�"�Q���ខ�*�@��D6��m����ف�'�����xԽ����}F~�5?��DB��*?��z���ﳥ��2$n��@�B2��k���;kvvq�^��1��3@�6bI����P��$��Ш����l����+��o�5��c���@�?��������>�f��m�7�Rky1B;$�y��X3菻Y�~����y	����� @�%�(@m��9=�u_�p���DE��G����D6�@�Cl�_9��ύA4���FS��4!N��n����qPc��e<�kD��e>>�r�dƮ�nk�{���B���L4�l-c�]<��<w{��ɦe�V���3.��.�}�"����@6��VT[�
��B�7��don��\�3~�S���z�j^�Y�[n�^"�>@�"�mШnjv������t(p��k1���+�y	��P�G�I�K�T�W�6Em���f�U\��$80Ka�d���:�&��	 uˬba�շ'��O��Q3�.=��P!~ �lЏ6�{3g����2�g�SS�� �P{�о�!@����t��C�ۡB7&wH��ix*����~������s�����+�����^��>m��Uί��<�ﳻ{��1
�Ё�H�B\E��
����Kal�_��T#�pW���T}�?@���@m׫��0�4��/��_�a)ϖ����ل�|h@�Cl�l�{n>S���MO���|E����}
k+��3���F��0l�U!-g���	�Y��ev�;&rӔħ�(r���W��9Ҽ�vk"��Ѩنvk���R`BN�m�y�0 �
��G�͌�w��u�|7�ۧ�����+����h@��|�96͕����Q&(�F�(�d�i2�Ric��jŽE���&�V�$6������'��F[��E@��P�ψmР0g�D������"��U��f�3
�J�\���=��T��+���l��6ϻ�>����ُ��F�k㙳�=���L�
jx]|�|E@��B����۞]4��1�SG��7(T�С�H�� 6�l��/*��?�2�iE�����1�?��!��l��g�� ��vO�".���G�&6�W�g|'��|G��5�𚯅{����K�Jv��@���l��BCl��Cl���ӿ�����ˢ&_A��EO�����|Ez ����ۡ�
�(U���M�d��@�U��>��p���u(�=��hC�=��W
*ɷ]*�4��+fT�[�y���ܶ��'7͊��sI �Y��f�Z��[-[�B̍K]L���Š�Ԕ��hrhjCeBl7J�̭�P�*]v�d���fնc�h1ԋɦ��v1IVF��R�LJ��!J<�f�+��ªt(�;J��1�4SG#e��-�B���i.#ix3ʮ����i\�t�͸�k�4%!\�@Y�4р��L�<�`�]�f�Z˵�(m帮i�����k�2�&��Z�B�E�IcV��v����S2���9�H�(W�#�v���g���;��Δ_߳��1�+?�ߏWܧ���<�>��}�m���D6Ȩ{b�|����xo:���{U�$}��Tr�k�P�龜����b{����a^a�G&h@���l��m�#��)n(���lš��T��w�J�!�T�.�" ���(@�>�ɀ� 6ȅS��2��ɏ����3���+����������׽0nX�V}��>4 _���V}㵿����Fo����!�@��y���Iо]3�,d^9A�nt���G/��}^��#� k����l�_���Q�x�8��m�(�]qMFV���4�mi������f;:���u�0З��ӿq����� �M��6�f����p���"������s~�����,@��m
�����
���s��_���Uڅ�Q;3�M�"�ܼQ����9P�Pp$���A�EU�o<��:��F�"G�?��ܭ�s삹���ӱ*�z�Uyt����p��~�?�>YdL����ف{5Mޚ1�0�"��!�0 6�\�r�{��eoc�J������ G�I�u
N����l��}��VC�������#��Bzf�y�2�|��0>ȩ�]}� CӉ�p-�C}��<ӡBn���۠|���3k��Gvw��+�i��r�?@��נ@� �m��6��|���Չ�����	Z� L��ٴ�	(C2)(�(
����!,l,��?���*�������Ͼ1կ>�/�,����
6;6}��+�P>N�y���5<!�j�x��O'�)�=�jG6j�fY��Qq`}�S��#���(@���W���+��IHXuE��$���r| @mШ��l�Մ�t�����Pъ�>U)�aDb�N�_���}"
{��9���
�.�S�����W��7�[��-^�(�gάV*\�]]�u�p�{�m�A��X�c��?z�Ё� �m�P�٨�39,F��Z������6�Vg��ןI����V_|+�}&X�;���ϧ����^��A�١m��l��m�1�0>��gZG�ή�g;�
�u슞_x�|@��!�0 6�_��������z�=�}-3���a�4�@\M��\L�En*%�JmTE��	rm��>߿��-ϊ�B�6��6�~dm��o�+�C�g���';�V��a���S5=����D6ȡ�����ʯ���E�$�W�|eּ����|.��w�`G���y�U�Uy}K��e�A���#~���Ͳ��em�#��-�4M}��*��T�	���|E��s���B��T	ߏ�_A����}��ݵ������B��>Jk�C�g�>>�	݌�:��ع�{�\�z�����E⩡�UD�a�oX���VL��/lz4z��X�E��]��}�+�*5�U�QW;s��%]p�7>5����dTmЯCs ���[�����O8�w�F��|.��B}����|܈���D���f����	b� � щRR�<��������+��&�O����K<s�ڇ����d���f�����m�晬͖N���u��"��u������/������};��t�����ܑ-�	�^�X&�郳o�|;�>�>nF,�~`�L|�W¡����}�h@����C疦�"��[>쑂�*6�T7&y�B�+1/LUfQ��ܪϳ�u���y��#���"΅@m׫� �m�W�RFo�"�!6hG�f��������G\�.~R>����Ɣ�W=��z��cD/���Ш��7>>���r��jf���2'�<��E1������#�v�h��9z�r��I?� ���@O��@!$�$��	'��@I?� ����@!$��O� �BI��$ ���I $� �BI@I6H �,	 �$ ����O� �BI�$�O�$��@I0	'��PVI��a��΀�ޗ��Y���y�f����K��X    �@@@ �   �  � @TB�	(��
 J�@��(���)@R� �3�@
�J��DJ�)EE
"�U%$�D�$���� �*U���JQR�m�+�4hhi�oq'��F�@+�&t2��"���@(Ǫ�2�4hhk�>� �p=�}��C��� ���@(/� �QI%T���P:h�0P:4���8(
�I� u�h�Mі�F� ������A����@�R%T�B�G�����r��  � 邀Qʩ(Up }ǯ�Z�UYл]@��@.�=y�0�d��tM�]
pPo�/��U �Ot $=t P{�;�7`z{� �th�I��:��"��zD�m���Ѡ�F �@h��7X��Z=#J5�}�� U�� ����
��!���7av;`&��5F��^���H�t@�Q)Ǡ%��G�A�y0(
94ht��@P:�� �   ����*���`�i�h�4Ɉ�F�LIJR�dф � A�� ��T�e$�      O"�L�J��`       ���R@ �M0&�&�A� �!4�@LBy��ɢ`M��I����z<����=��&2c��㗎��� �?��Rࠪ� (�X�ć�J����	�[q��{�~a�d���]���j���q �'�EH�A�T���ߗi��  �;�S(EF(�!�E@�3���׹�p_���??�����yc�q�s��٭q�j�ֻ�@q WqWqD\�Q�CpU � /�DqP�wM�U�@q�cf���Zֵ�wwwwsww^�l�=���C�Ϣ|��9z�A���Cg�͓��άk��K���Ň��?��+��0?�5�0��*�e\p[�<e���iދn����1�
��q͚m�!�r��svq^<�k��`��$y�pI��.5��m�^���rœ:'������X�j���	sr��B���V�Q�����yr�-�lp�bJn��j::��{D�a�ޭ��G;�����{���S�D8���jn0�-n�OX�n���K�4]�r!�T��n��&��ե��7d\\��D1ڗ>�҇`�e���$�;���7�L��4�]��0d�I� nS�)�Mgt��b+G����1j��g;�H�@���u&[�9�� �_t<7w�h)l��t\��u�OOu��S9Շ��L�B+N��,+@/z�1��]���dv#uFQ8��a������y.0y�o�SlɅt5Mםk�7�jh\�14;g�BQ.��u�i2/�<��M�S��iY�]�ɲbe;��x�A�����L�:�]�89G���`-�����ɷ.�]�9�UBC��N�lp���	�p����s���Z�ڤ�����h��Ue�m�
�2U]5�[N�`��@#:gZf	�]�^	��� hź�ǻ�c���!8Ѷը�7�NN��{h�7�{n���ƻp�ƫ8�-ɔ7��6�H.V0��7�-��Ï�6���c�$�"d�����ĕ�	%M]�����IE�z��96�/:C�Z"�X�=�>�m�f���a�J��yַ�3Z�z��f�	Im�Wj5D�����NR3�E�޵p��6��y�Rn������*�G�
�o �F:�܎�(ͳ�_�Vi1I{mgp�
mǌ�D�[}��+ihtٸ)���d�|Ք̫隱����ٵ�]���1��p9wH�W�z�R8Y&�<��F���5���T���yK��s��tɻ�w�S�ܨ�q�Y9<�N�xd�Z����X3����8,	�p�Q׭�7�3�V�>����]�H�`�W>�Ɩ�K|��������ܣ9�r��6�;h�R�9�9n)�iP-��^fSX�^T�vF)��Pt9E��iW�j���9���ݘz2q��Q��[��8ȋ��ӱkIwKS�z~��Z3+�Su�̓�®����b����t[��+�/�
���qT���uMm\V�� �X�"g)����z�9И�^ƕ��m0���D�U�;DӸ�;{_�H���s�913�$(�%{X�
�Y����y�nf�3�;_6�y�o�Mj]-�L+7.+�V���\�d\f!y�-yG§͝�*E�Kx�x�������b�8c[�X�y����tP�eg :u�+cx��ع�v DH�(2�P���)v�22��ɡ�r�jXG[���сV�1u���s��_f� �T"v�������m���K��7Gi}�vW�r�}�B1]+���>�7�#���(�ș�����p=з���-�\�-X�"��i=�6�VR��
3�Q�R'�At4�����N�p���	�n�qP��z;W`U�V�h���#�6���i�rI�ʈƛ��r� q.��f��zb�7�x�%�Hoc��n�'=K
�7�����3.����]0mI`~�/J�����w7F��9ˑp�0iЫ����A�J�m�wIڛ3��2�!c[�fv�SRv1�];M��N��VI�V��M�VZ�3��:V��c�E��r�� �#+Z�j�F�ݪrպ~�.��;�����w�Kb<��lU�_V��+���/,]�K����6�^k����5Fu�Nw7��s]qo$;_�@�����i�oI
lX,�a���d�"ۣ@�K���A�5����/ b�ŗ�����D�^��&ԝ��c�!\���]	n�\3z���6w.�_ w���P�� hI0�bG�� \T2�ׅƋ�#�B�UaM��P_������N����-��N���M�Ή�4�Bm��`\�/�8P��U�"�ˑ�p;ƻ-�NtAۗ��R� �s�8`�"��f��<�;/&�Nc�Q��p�5o|�h(�w>!���8�A����q2FJ��`YneB)�lK%Ï~˄������L\�X�j���q��7���#W���ڢԇ>/>�+���kf����{��,	]�~�X4���B�X��hH�1�l�sw�+����x�dv�%����[�7=� ȱ����Q3+gg]ߧb�pǤ�VLԔ&�:��	蚝��^U�Lc�mCI8��|uˀG^9��0ڠt��Q��LNu��'e�Ȍ����8ZNu�,��.�Ϋl�rr:�<�ꍿ�V�WϷ(�S�msQ�vQ�-m�!ޛ%��n�V���Ü�M(9�1n����wI�w��u���|l���U��7��y=<��*�IѹSs5h����������]ևۚ9jV����:���6��+]��G��..A3,w�ݬ��$PfŴ6Mq��>��?[�����ݝt.m�*}[��La�Ip8��e�P�l��㽺��voXzm�x��u�;Z��5L�^��tg+�2m�'<3�^2bl����7�(}({�6B�yf�#�����Y�1m;��R�o'�0;FI@ŬQń��.\�Ar؏.p��uk�[��Ԓ]K�]gr�Q$u�FQ�I���H���i��;�`޳�^[���܁M%�x����{㹦)����[Sd�8��ra����N�Rt`|n���2[�v�L���1d0i� v���i^�Ő=ȴ�!;O���ޠònW$N�s��'=�;��isfh׋V��s� Xȓ�H�Q��.��ٱGe�k:���Uܼ�h����_NgP�	��a�^�����N�j����Ys�C����$�w���ҹ�j],��C��I�'��3�X"z)��/a�OЗh��v��zC��5T�H#���ZY�ݽ&�^�xnW������h���ՊmRә�+��j�����]���9�R����h��g-"MQ�xF�����4�������FU��>�%2曋,һ���y<����s���ed1c�qP�ٛ�6�UY}6l�ڹ���zf��G�n��Z������1jYZ��/c8W�U
.���1[���uc�k�j�iĵ�.���"��ݝ��{�ǹILo�9i{�:L��V{LZݿv�՝����Y�ǓV�X�&捨��IˡL��ç#�1"[K�I�Z��K~:L�m���:��5�H<~���bS;�A-��s��廑���b��@�QwP�(׍R��2f���Ѷ�ivb��lX;xM�&�m���UZY�=[Tۏ]縯A����7�q�rӸ���rv����J�,��\5E����w���-�E�iA���(�)Kfk\$׉�:����=��5���������یwhg`��7��u�l���ZI<�ǯ�o&]�9콸�yV;6�l�T����Ï(��eh���N'a�K�SK֗]Mv7��z4u��/q�s�f��$��K�����0��u�F��o�ut[�����({aQ��
/�=R��Ǉwh�@��\�W-݉�����i<	�j;(���4rvȠ>qQ$@Y	�	FD$DRBDQIV@P	 I@�UE$@$AF@RAD�	FE�@�d$	Q�E�Q	A@$	P�d E	AP�T�$TP�I�UT�A$QFE	RAddQ�T�BE  $AF@P�REG�V���+"�Wl�w���f�]�������I{~� T �ؒ�+9��D��ӣ�W�'î�ڒ�a/���dTP���Q?�����������������c�wi�R�(��KxT��ޯz�5��&;�q��5��=� ���{���O�����ɏ�-e���=���Kɼ�MۗB�� �=�h�v�f$@�vቭ��R�$ ��Bݶ4�����u�p����Z�?"p��sV.������;�3�at�o��|<�In������vw.ͮr<<�U;z]��0�2!�T�iZ���:�S�_����4�J�������������s����dY�.'F�9�q#DQ��3������ڍ %l�/Ë��N-���X�j�dR\ݗ�1���.�X�>>^��l��q@h�l(�����gι�=�\}���Ƽ}ݷ �y�A�L��f�{���Í��ǚ������z�q�>ݖ��1��٫���O5�m~1��[uo�ʮ�ܡ<�t`��=3��z��[���O����M�Zdd��[>��8[��!�8��]�soq����9p���d�EH4G��T �):l��<)���;ks.0��!�k�{�dxyp�G��k��y<�*N��P[����^�s�*���'L7Ʀ������k]=���R	��Q-��>m�~M�=���4=�ս�Eu��=�%^^½�1L��ˮ<c��wq�Թ�h/*���4�Q����a�;�J�웃��:2�ִ�^ο����ƹ%Aݏ��Aſѹ!{����ƺwo6U�w�kc��i���["�F���!R��X����}�t[����;���[��*&��}�
�����)���x0�O]���Ԗ�����J����g�E���������;ϼ$�P�}�cא��>nv���j��:���U���ؒ[�ra:#�
��^�{���pܸ��4.���Hꯉ���^��%�^���˳9\s���ϳb2��M)����^���X��RR�xz7�;�(/��=��Z�A��)m:�^Fmf�9;i5�)����E꺚�=�ჽ�i��)�2P��J}p�����3�5�<�h�$X;��oc��>�E��ݝF=��!�pjt�(��LZ�M� �6�^2b��fb�^BQxA�w�e�9�L��F��V%�l�r���ێ�b񖎆����bF`,��/��1:�G؞w9�	�7��8�T��[W!Y:۱[-�0��x�A� q�{.m�s��V ��l��eT�����r����M������+���y�	5����"��t�����M]����udKOh��3�0����IA�x�#L����b�v�Nt��CYw�}-Wx��Ԣ��)���cKä^+�bƲ��TE���{W('J��l���;�@������`�b�-�R{�=����w'nH�䧵t��n{ۊ��p.��J�w�dN���hRxܛ�I�b,���Ñ�o5��zV������{��@��UP�z��O��r�˼_ҭ+|�;<����ny ���K��_;薕�o@�j�E�!�׹�h����<���<,dE�N���< ��W��>��!�ݾ��>S��cK�9�7R�t�����ȬҖ�ה!�N��9�b��������Z,�t��ў�H��9}�ǜ�o{>ݡ<%�ץ{.1����d'��]��λO�O{/���'���7=��f#�;b˝�w��+NK^R�5v�z`8)=��d����)JW���k���ґ�Y�A�n����6k%u��&��T��7[�8���q���Fۂ҈:f����y��p��M�<�����g)���=�B����c}�OD֒�C\���^/T�)Р�Q۱3�WmX�$E�x��o,� �Y������c� ���/#�ss�Q��qn�q8X�t�ge�w+i�^s���Y����⛿0�l^����#�	,��xy���r�mͤ�Tf��Y���=����,Y�N�d�f�����>���j"�����ڼ��K��܇oz���7g��%Yz��rxdE��P�nj��b�;�c��5�2�5�vuŨ�{!����X����v�!m��'��;�Xs\��d��=Ԗx�{r��;W �a��;��8F�ht������a�s�.�nL*_Js�~{-��4�sͺ$���C)�@��U��;�!y���qwg���t���K�d�ށgo�?g�O�9{_>��ݩ8A0Z�[���S�rKY���)�Z����W�ְ����OV�۱9^�ʼt��/�:����p%�1�p�]�>��p�-m\����b[����ň�Y�z�5�a8��v~�.dM��3n;S��3��)�m�?O<�:����r�7IslV�7��-�A�̗s;��=pg��[����d�ъ��_ܪ]�7����2�2{��w�=�)�R��RyX��	<�h�&H�<;W�vTߴ�f������yk�r�בJp���f��y3��9wM�b����[���F)s�b����ז�.�O�*�^�w��o�kw��_K}J�vø +��ك��{��/��������IL͆��������ɵ��	�hfi�Ġ�	jf;��[V�~s�ƈ��|��oh��F��/���/n�`����s��Ӱ�.������d�m��ToF���#g��>8S��\����t��o�U�[���]̺S+qz��>7�s�Op��ܤq���
��A�W.���HJ�a�N�C�na�\�Ꜽ	X�M7��_�{<P��ۣ/��F��_��F����X���p���A�kSu#m%:,S�����oX���MIv�|7th��26,+-g��~�yP��K�yM�w�\��9=�x:=|Y��kү�|���n	�On����V����ob�ͷ�E���0bg{J���@vz}��1�M�M޹���cۻuR�sa2@S�=��_g���Һ�?���f�uHG]�싏�)*��N��v�fݝ�cZ�ZK�d+��_�e׶K m+�
ǳۄÇ���s��
{o�qlH�q�.�Ѩ���C�{�
*s+Nn��/I{��|�*�KM���_?G�"+��<���a��<z͂LՔƆ{�΃�Cݾ۾��W�8u�0a�%u->[���!q��7��V��K�H�N�r�
�;��p/o��	��m�-�g�ɶ5*��z�_�á�g��ԧ�ٹ��u��#��e�\׳�l	ɻ�kw͖�j� �
�B�/qK���hU��=��8�������֟W���˽xL=r^�}���CQp�;9:�٫�We���Kr������xG�,����靗�=z�����}���`ަ�ނ��(ߔ��Sͼj��q���#��+���u7h��>���zl��~gA�����]��!:F�A[4,�y��[Y�o�ci����G�M��gu�3Ds��{����zx鷽��&m��r���|����*��i88��^�5��?B,��|�;�z4;йA�R�nly�g0�����x�F��*�Ǟw�qy��7���'�sX7�>�]
�p�$a���x��Ԯ��wB��7��:�3��N��+Y#BZ�r%����I� .�y`C����z���m^���p�%�#�x�[�yNm^���aCr�Fi�S�������I�������	�1�m\\��f��~��-G={�� �)��|�Z;����`���+fڈ�A�k]e�TE����x=�6\���<�0��-�:�2cA�t����o=�W.���w���0���#ڪ��ﳷ�̧1%sV�ƬQir�[����>X@���L�<�e�\ʀ�\ҹf�k�])�����r��ik�V%�6���f��ٛ�0��FP���3�k5�ζ
�l�  �a���z{�<RR�[]v�62�ViVb7L�[-��+p��-ɶ�d�X��WD��b�ը�X��S8�kKsi3ڶ1D-�qq6��Ԗ�.h���qi!��͛��f�q�ĺ��f��au��\�wC����t��HY�Ff3�*$0��6��J�@�`G�/Z�r9�1\�ڳPX�K�1�;F\<1-��)j��:M6�QL��Z;6���h�c�w�e�F�9����j˄���hb�2�eŦem"���K��5��0m���tն�r�U��51�j��i��TZ]qJ]J`��kJ6ڰ��d��M�m��b�
ˋ�k�MG�4
�	�t����Թ�Ѵ&s6�K���ϙ1il��4�u�4IiJ��fP�b���U�ѭ�"]��Bm��W�pDs�,���������e�-٦u�Bnk�Aq.���������� "�U�@3�<]U�;]v\k!r�l�j�fh@i�H�A��n�	�lWE�.G�[XV��j���!\��%X�5Ԙn6���e��f�"�� Ջ�(�X�4�����3*��D6Դ�NtR���.�\XlSlH�P��m�F"��-wXٶ��.�-Z&�#+���sk��.B`Ѹ��*GE ڍA��n[87h[�T�B`��*4q�6�\�1�0
m֒��bʖVZe�o�Ś�2ݖ,lMZ���U�V%u"9cv���A.�  W��b\7 ������YB)�[K`�)v#s�M��A��X8��
Ь��ku�u��`���#�[y7�F֓"�tb8����MXA9���D���v��GLc��c����e˲�I�:��St��
�E��MtCY�Q�V�2��QBb�^a��p޺�=gC:�`"S��&� ��U
Z�Z;:�P��,��a����m0��1δ&%&��Xִ��j6h=� �eҤf��f���]÷j��i)j�=�Xy[�M%�]l^&��%�(�tf�XܕCh̈́�B`�sv�]M�u1-��΅�*��&e��˨i���虷X��+���}�fD�ea4�˩[�,]	lB�&�q�%�9�ţ.��ԫ1�[�릇��6Z����ٌ+up	�
fS�r�l�K4�<t�A�)B3C^X�36��뱹�2b`�8а�cf4�nEn���Z�a#�ё758�(+]2m���[�5�#*h˘��e+Z. �MtK2D[h�]y����k��!P�j�C0Mz�i1��L�K�8m�,eo��9�Mw�^�}VZt��lU�m�4�-��-������Q%Ω6JUUbK�sF��G]�	k���عը�D9��%��xgPA�Sa6	�tږ��-EL�bm0b���̷��Y�7�D&�̰dk��vԍƻBKP��������H�\1p�^\��훖g2�()�&E	��r@��.����� ���uB�Φ��n4��5`ۥ����ݣG���3\(3]o��%b�C� iQ��B�0ʠ�YJ�6�s):T�@)SjD�m4SbV�]�G�3b��Xj�E�`����\P�*ˆ6�LE��L�m���(���B��l��FL���Ѐ��<L�16��]��$�7-���XJ�mT�f����c��ye��,c�]lѦ�����5̓5%���5e&�eҐÂY�JǃCKWuD&s��\vֺ�umʓh���H�{j�K�K6�al#�ĵ�x�mٱv�T��[�IU���K�JimBѦX���:.���v���Z�4ԍ��K�e[a��
�6n�d�51M5����]5��M�
�C�nD@-&�ٸ�f��iCJ-&퐫j��22���Y1w5DV��i�3b]��j�fcjV�+3�������(V���i0�#�"D��K-ًfkRJʕI^9�B���]R�tbi�2l�9&���6�I������:�:�1�B�K$Κ��Q�7�m��)2��K��+ ���������i�]�t�lXp;%��.��#��]�\�+rh⹐�)*$�.�!�Ҧ՟B����в�o1�\�p��N3C:Ԕ7Kt���P���n�0�ti��+�!�,.��lF�Tɴ��2��Ǣ�oV�T���2Lܵ�3��b��-{KM5�.4���	t�b�k���j�yc�9r��[*h��M)H�m4�m��q��v�Z���x[��,��D70݈ͥv�����F�K�\1�911!a,��-H����J��CF�¬Eġv�J�%�
-@˭ql�fu�&�<��m̡��A�m�#�k�8��C��kx�&�Yh6��Pp�<��s��X�ggr�ĺc,�lk(2�13��c,���f�ƌ�b�X�7+�$��+.�5L*�UU�Vt��Ebm���Q��ݙ���e�n�R��&�.��H0��ш��pf���gL�hZlFV-���(�R ����]Q��5�UUUUUV�容UUUUU�)T��+���jF��aT��4U.(�X-�A�&�Z�/��̻��h�7��&B�MSf6
Ǖ�J+�R�	��3�(؛d4����Anα�mI�6��/�֤����"��ˈ�H �������*J 5�m�[$ZQXC����9�>����EOZ�E^ �����kEݷ�DEq Ҏ8��4-*]��0WiP۫&1$�"�����%�)i�[��7"+$���Ec�����Ƒ�͗�a�ӊT�X�
t !:��XE^x����x��e�)�	3�P2�	��<Bb'U$��r�	R�n9p��"4��@8� %��G� +=��TU�E����/�UAܓ�r�����e(�:%]��,Z,��6�8�\I�6T�"˵B�2��44�T�\��	M[,y��j�C�M��Q���0kL�r��m�F#�+��%���36�q�cMWT�挂�͠3cX�hG:iQ%Λ-m�VR����F�lR�����#,e�CS���.Ī��`�ԕ��Ն��⁜7%it�nW��\�a�5T	MQ������`[�V�&�v�.����捺���	��@v���B幖Q�1�݈kE.��!mZ���ڹ�������3�+��CҀ4�1�]/R�*��x4��e�8��Q����fqFe�ꖳhE!tymP��%��-�ʛ!�7��7P�-�G0-�mM�܋�b&��q�4�X�[V<��X�:4�]���-����-�q��-l��B�2�6��h�^���19��s��R6mjǍ�3`eƊ녺%���h�K���0^�.	m4ŀ�J:`�ȹfW��I�-��*2���-��ZV���͇it��ܗ��'FP ��m���mDZ�-A��J�jK�����dX��l�[a�"��m�� ����ń y��������@B�1��v�.˖�����~
i�rMq�GBiA]�":�v����l��0�w˖u��H����8"�i�z����ȅ^������ԏ{7{1N���2����y���-��}�f���Cyڏn�A�wtuAG 1d]�,�ӊ��*�x��ve���G�b��W
ΫJ��4�y�L��m�e�b�X�A���o"��^w�v��]њ�R�2������l��
���t�E�'{�����j���O�5��lDV ԍ���Z=��w�G�oP��n�胭�n�rWP6��7�_R7|��oN��S��Y���m�������p�j!_u=�!��!��*ӛ��G;:���B�!��Sz3N18R+��nX<Y]��e\�����>fj���6�����=>9Q��k�9!�fm.u�������w����{�Fda�fr��ln�'T�[	��Wq-�ע��2�R���:�3vA�3u��僜�q��ù
-��=h�L�I���v룫�&N�C7'1�ۀ�Zػ�Q�Y�ۭ��U&C��*z��v�Y1��l5"!6J�WKV���6[�ߟUl�b9����u��L���5F���뽍��xa��뙘�р�#q �>lvt�tOueun���5I�ێ��)zRq5p{����[�GTtL\-�ԯy{�BZַ	���#_�����@	���g/�r��Ci�WC-H���6����Ck�D���*S�(��A,���xՔ��.�ϛ��y�{�۲�\�A���6�fezg;�	˸���;���{�	��u��S�qйVfT���T^��N\um#����f ��TUL���f��G������q{O�P(I��\�Z�/s �o[=ܦ�&j��k����J�uoU��k6q��M����~2'&�Wn^��9�hZ&i�fY�����f�R�M���Qɶ[
�.�)DL6��*�Ԙ�K#���v�e���p4���_��OP/�Q%�cK�Cp�]L2��Δ�;0+�m�.tsr11�߻����t[H��CFgS!J#��HW���:�׎���:���Y��_Uk�3��2�t�U�%^�f�wL�=�Z�=ȬKHF5n�333�*�9;Pz�m��Bj`L���*��ʌ�$�뾍��{�u>����p��e�̰�e���Y���2�f�L�����������dٹ�%RĲ�#rDG@~_��O���]/>�_{6��i��d	�*ezlô�Ff�=䛵�5X��WVD��ʊت�}�-�{�u5�h-e8r]`�nx̼��c�CO>��N]l}_R<7V�3d��QC, <C�+�}3)εö���feÄ]�Kr�T������Be7u�{z������׸�}�[?6�d��wϟ�*�=�ΙC����-���t�Q��#�H����isƑsr�A��{ۓ2���n�t̢{�P�^������*�"+�	x�u��w���ޚ����O1{�Tʝ��^{�k$j˪E�DR@q�]\�O���59�����W�w[H���(z�TQ��r�l`�TD�yY���2�=���6wj��dL�37�κ�X�!ooS<;��}3./3m-�}�������W	�+���p��P٬��35�c������6��eE�����w]f�n��=�d
�3��B�BL���g
����f#w:��.[a�ڋ��ƃ6�wo#k�p�h�tF�V� �h��!�q:ʌ���J�ۋ���RU�^q�N�}�7gD�G �lHw5����ޙ�x4��w+�˚Z�M����bl��E�Khǚ��p���365��;s"7���ژ��-�qq��n�.s;���Ԟg"g{���m�p,��2����ݙ�xY���#�zfl\�Q��������Ό;�F�ۈ�˜Ñ���ݔxn�ig��D���=�-$V��4�A}�g�;93Ǽ,X��:3X���ky]��K� ����!	�m�j�f3bd5a��+`���	��!Qۛ�g�0�T�k�W����hh�K����֎��к�ddf]u��n�6W�W7k� �BjM�rLj[2��8#r*�{=�|M �ڭ�ËB�2���m��B�c�N����f�L�=Q�v2M��@m��
1�/LM^k�̈�ݦs�^RL�v�D	n�g�����dw]��hv�%�k������Η(��:�(SR�۬#	ᙕ}W�۴�{L�oS��Sv֬
!���Ã�1c3���Z�`$���H������&�L,��E��Ƃ��A��'�����ݬ���x�Gq���\�UQ�]���&r�l�۫�ާ(��M�%�vnf�6�<z�oTE��3�H)�[�ya7i������#�j��t�#��yꙙEj��ڝ��Χ(�)�Gmة�H�vO �D'�"Âd,�*�f$Dt߿_{'Ǜ���L�j�������׳�X�bg���]�^�Gc��qE�� �^���5�?���/��F$���]�g�te��qD7_�H4�ݡ\�]/ج���ܐ-~�<ωJ��$�F2F�����E���)�*؋�z�R��;�m�5j�4�r��x��̪f����N-ښ�Ӛͧ[�UGa�e�w/�Īz��5x��T�6�2��v�Z<:�ݝ;�fn�`e�������Cӯz�,'�PlA��т�+����9&F���+MҞ��0g��G��Oi�
����=8J��7.'<�wvR��w�{%z������v�8vx�l��=ڼ�ec����~�{驼x���-ɾ�w5<�͞�xp��.v�B�G6��n˽o4P�D�&I6���D�Q2�D�Tv)y���:��bþu�j�q�����p4���E�|��.�]�ΦL��+�C\;���	�޹i	����U�,&'Zq�T���>��d� ��|ytF�X��:.N�z.Ȋ��Lr� $�z!-�����1�`T�X�C�G���)1�	))*�V��y�U��K+m������lԳK�i�xx��PIgKy	`=Z�6�V��
2�cN��K,+��n�Ɩf�Q�b���d�@*�ĄX,B԰�Ym�"	[��Wk{̵8�"����T�0�� �bђP���a..	�ō����{�H�5	r�X�Ԋ[y���6|/��y���G�!2�$L�|��U ޻��#~ݦ~���IK32�ϦbH��}�c���.w����G�Pրn���6�[6�E�!�t��m�\�JKX��X��D������t�N§�V���D���lA���=�ȏ������o2Ŭ����3�C#B�y�Ϯ��>�f�;�ڻ�,�Uu�}��G�f����y|��L(u�}�r�g;��n���ƭ���Tbܩ��7Ob)���wP���|��A��4��M}�ﻥ�}2�U<6��<�G�B!�`Ci��2�s��c���w>K<�t�"bf�3�]�o�R��4�m�����l��{;�;�ݣ�l��5V.n�C!��I���ݴ�{��\6�Or;��F���3�ݜ��=���R�a�� 6�-�C�u{�����-��:xO�j���}��o l��Zf���Ѻ�j�(��+����
��y.���z��u�B�ą�[l� ��9Rm�����]�� Pa�\����KR@�4vtιÁ���0m�l�n6��`�i�A�lfҋ�X�i���@�/6!�Gl�MA�lf~y���يT���(]�ʗ-��m�j����t�>Y��mG}ۑ��3{=���j�Hd6�����"��3s_]����h����P�2�ݸ�C���3�v�Y��e�3g�����h}3o�؎�z�����55L���2ooR�\�U��nk���@ag����;���՟'Ȯ�]��\T�텲�}�޾��>u�~���=��#R���[�צ� �Q����[��|\ѵ>�tSĲ��q�L�\�&�T���5�_/�;��b>�6�ߜ�$|�����R��2O�|�ģkv����n|���y��#���ϙ瑩�6~���Ωy#`<x��!�(֤��������g���e�GN���QF���K�T͡����b�C��߬�E�=ۚ���y����!��_�UR�	��&�j���.6Cwxo��b�M��ߵ�/����ƺ��6�������7v����i/���IvV,�3�[��������lGf�3�|f���o��tq��o�������}tw7���P6(Y��~����Y���n������n�D3�q���""B�B�)V�鉁���>^2ډ����x@U�TuV/3�~��=�ZoO�[�Q;yz��=�Տm���pýV��]ӱp~φL�m|�&yFVcK��g�dF�m3���{�~Fzk�~s�?Џ{��y8A��/`���;���ͪstVd�dƗ�A�ީ��
��*�i@m����NkYAQ@����{�[�\q�@舒��6���D�� !�k��|۞5���u�3ř��ڙ4�U�r׵��@�osH� 8� � uu׿O�}�K�{փ�ϰP^b'����� �(�N*��\�L�@(�����u�[|��/�
���DD�i �C<c�-X�� �(.A\�j"bTG�,DD��un������q��u�q��*Q[�lDMDJ��Q@�)� �A�ѫ�n�Cp���%�;��}q�������^�:`��5:̘��PqH��x�m1*#��nwZ���<s��[�u�����LD�i�D(�8��]:��琙���G���赳z�*ˤ�l�w�w퍥\�c���\��|zQB�.hp��8
U�Kt�*Z�+���-�33͗ �B���������f�J��R[��:�@�	�l��9%�;S�E�[����˂�	��J<���h\����a�~�=�
�����<u3�0j�5�I7�'�%��`���c� b W�9�[�:㎐*D�ѽs��Y��9��D�P���c�� bDHD1�"KuU�V�z�\�`��!QP�x�x�[�V��/T�s�"j ��bUrb��`�h���(DI�D���(P̅{ɗ�}˼�=�n�u�/�
��z��D�i �E�L@
b1H=g�sW/�p�:��4	Qj��q)���w�����
�=n��D�8�W�d�(��y�Qu�@� �
���bQ�K@qѝ����� Vw�g<��:�z@�R�G�"j �p��#$�??>N��ʆs��Xdu�E%Řq5ʵv��"I����h�h@�E�b�-}�z�������u:θ��'TG1\�� b ����ANy�u^�ί�u�w�n���.��#��o�?.�y��y�:'uu�|f
���>� K��� ����z�[�\q�@舐�kt�$9�A9��1|�z���@ f
�
� ��"b u}��Щθ�=s����^���4�I���1H �������j��H' j � s}�:�oֺͶQ��Q ��5G�W��9�Db�m �(�Q�(Z�~5���`�Y��=k㍠TA�kt�$�@,�b�:��ɍ^���]�c��`�c<�Va`�|�H��C1 �@1�k|g=s��g��Q޳-� � Z ��1�!�@b�B [�&8�J�V�']DZ��R��9�s~��m�@�
�LD�sdKD1�0�� @�DI �+�c�x����U���S�3���/2c�5�6�3׶�\6>-Ų��g�Cz}�:����f1��ֵ�u� T�"@�kt�[�1 �D�1�@1z��(��� [t��Z���x��u�s�w�u���A�D�P@�:�Z����6D���lALAqnz���c\��T����Z�9�[�6��Q��i�
�8����_}y��u���1/S6�V���/rֽ�Z�@� �#���%Dq��@�@�w��ַ�u� T�����w�f�䈝DJ��Q@�)�(����4f��f*䉘\s�s�:�:�z@�R�G��5H�Dq�Z�U��q�Pw75�@�"C�DG
����R����u�c���f� ���Cq �@1pD�@1���6s�_|�s�N����%��4ȃ�����<�}_Mw�� 3P���օ�>��C�Æs��/m3��'F�G"�Y{��j浌�8�����}��;":�TA��,@A1��k9��i���z�~}7�cl:Uu7>�'r�""�����7A�.���":�>�SM�N�M?���bu���>m�d��R�p�s?^^�M���US{+��^q��U��n��MA�cm�%Y˸��m�V��}�p{�o����6�-�d6�s6�RC���3���f�m�;����~�Ѕ/���ú��n�0����4ToF�F�D0�n��çww"��N1_5쌷��Oy�'��^~��Q^H�0�N&�����4.�S�j�mwsŎWRۛ�*�"Ł��m�p����*���^�|�O��9K�J��;}�կw} X�Y$r�m!h�%���u�'�Ȼ�%@��� dtEy67�}y�j��� %�@f�W��m¡���77�ژ�2O����@�&x��~�=�Y�bD����g�KZ��b_^Ӄ��-��C���M�ַ��x�ci�E�99!��ܽ��.��e�w�?z��u�s�s�����-�zzi�ˆ̾���\Q��+�q����FWʚt5�֡��k��{��o��o/!�h�͞��|��ឯ4��j��)BttTҏo���u��T��m��-_����~��!LO���u�5�9,b�K��}���>�B�(E`�ҕx$��!�W�$e�րLj�2�k[uൔ�@�C^IH���Ù
I�rdHȴ�@b4B���LxezE��g����̤�A�Zҋık�I��0�% tHH4�Сa!���c*֋U֔�E��c���1�	0�MyyҴ<m�2�3U͍2����{K8���Z5{��P����(�D$�4eY5�eFҼ�]a[)F^����jd�4-�M������:4�xs�4��[�b$�~��I�i\۬4���
�g�bKbb�Up�V]�MY���U�50lYKQ�,f��u̅�n����f5/�
�D�a)�Wlb;g6%�i1B:�1�ѥY\�G)u��ն9���-��f��$���wL���'7@�X���[��Ie�vtR���v��n!�DSL��8f6�+5�����6���65�7�^��\Z0iF4�S���f�XK�VR��b6��P�� i��3̈́���15u ���+(�����їE�93+��.�F�B�Q�����f�4�;U�tūvSK`q��6i����[	�я-��K�^2��-�\ۂ����G�v�ɈY���n30���㕎n*�ᅷ�Ŗ��Kf(9�lFhl�"n��F0�#5�t�ie�2�ʦC��!��C��٘M��-�`t�GHf\��b��Le�.��\d
�����0�\�Į�B���̫t�`��(��Á�9�Sm�&#�r�Uh����n�����E��2���1˪W	1��Q.5Υ�p`p�;���З9�i���ո��b�l�D��6.��L&�CR��d#L�ܲ�۝�.��)����q��@�ˊ�l!�[�mN2
���\����̉k��s��LM6�T����Q�����{�����)~��a�̄0cD���d�h��8����{$4�+��5����w�>�m��ێ�=�3/O��/��g\���u�k,>����2��`����٣٫n�9����,������n;T���!�0&P�7^Sx�wvi�u��Q��v�q:���8~)&.kjݨ��M�r� �|�S�2�����ή�2�Q7�V�l��[��N��
�p�K�tƱ�v����ʂ��ڙ̓�m�r�ɪ�gV������W��~+�Uo��p{�y����*HmԞk��sӯsm�&�g̶�gpiې(�v.z�:�h�m����F�Ǜm��5��������m;Sum̅���r�����,Bpх��mչ�1�-�;��<�T�����w�	�'ibCm��Yŵ1��zj2z���h��Cc!�=Mɒ�g��x�����3�эv�ӼT��卓"���	&���Z�*�H����sy�����q���,��]Ue,>�US���{�L����v�^s0&TIJ�Uv_WU�jYo�/c.�O�b�n��nj݂۠�̹
!D1U6ᕮz�7��9o�ii�Cj �]8�^"�r���u���*��0Z0�ǔ��=�����uQ�Ս�d���wwO��=7����~���3�ٿ��b/��T�?��rU�+ޗ;cv�A٪�g+��x?���Qm��3�;b�����:��֏>�n����Ϛ�;��f	��dq3�36"��@�E��ٮ����&���h6���sg.p-��gک����;G�of\+!��l3��GlR;�b:_t��=�U�Cn2�b������35ד�Txf�7u{@�C���*r��UU���N�������0㿷H�@�%���b2��ʃ�=YX%#M��sy0��n��h�gmh^��� {��B��,����YB�m�Y���$��	�!�Zp7i1c��GJ�����ԨcX���3F1�b<�hF6kf���Wb�Un`*��iXK7lc*,��oL�+��|�)���t%M�t�nR`�EGA{�����z�v���u��;o�T6�����5U�6��o�ﮏf�{S�:7J[��gLE�/����S�xq�ἙӰ�Y[Cjn���u�����ᙘ�%�s�5�m)����޺<3V����+��S�Li �.�ĭ���浅G\1�X ��u�T���ާh�%�
��u����(�ޘ�C�%���3�����7Z�t8|�ȧv�Eg�r"�,�WZU�.G�=� 荒�^��W�Ol� �T=�`��D7������٫Km�J���n��Y3s{�n����*�f)X�-6���H�-ɾ�묭�{H�M�k�=����2�i��K�����&��Ј�a�\(�p�UW��rxʠ�B��"�m�qqȈ�{�s#
�����v���fA��B���ly����a߮�R.��2�jF��$2�m
���ݮ�'�1'�}�/�,^S������<<=�Y=w�mu��6���yKUwp���Ws޹<3b�Z���u�P����
�
�9��]���p��l8}ϣ���b,u�4K��-��]R�	����59����f�mu�c{F��@k���'{8*/1��.&��� ׺�ގ蝘�o{svF-���Wd�� 6�8���V�kvs������߶vaV��f�4~?@�'�ٛ�?e4���le
���
Yw�{�mz�\�O�{�����>-�۬�t��>5nro�;��f�,���Md@z`�t`r�ViX:�-r]�C9�#�� N�2�&z{7��Kf�#NF��l6���fb%��G󯺳�묯���͹Z���Q�9�;��;X�zc�����#�O.U.n0\L�voE�=��㜟���s����ܩ{�.Sޟ��_N�s��8��'�j�#eD��a�3�	>�H�ѻ���W�x��p��s���%���chu��Z���vbZ�9�2�������,�hӁHM��Jkq�v�2iJdխ���9l4f����1uK�nn\-�&�i�:�6�u���(����M�ժ�+B�������4f���܃n&vbE���D<?��E�D�Oc����;�WQ�p�]����&&j�w��F�K2���};��:̞��s��L�[D�����jvg�gz_��n�����FL���.�n*�w���N6q�;��<�;�)�[�2ܗGA�P��[�ۆ�7Z�Q���͹��'��72�f�d�T	>��>Զ���_/�۷�.b:LL�����>ɘ��^�Z����xx{�O�+�ED�V}3���j��췙YD6��R�Nw���z��2�i��ܢ{:>n]��t���q����=����[ݺ
��������5{Z�B���1���`���&�y�a�ۆ2�<��3^����.�jmNf.���mĆkjwz�m_s�쭜��xl���B�N�Qd6��_{�����C$M}̯��*�6 n*-ɧ��"��1Ks�G��o9ۼ>=^�&���E,ɦ�����â�|�����Q�{V��?Nu��>�yC��N�Qm{�lѦ��H��菒�<l^�%=�|�nr��Yb�8}v�����>#9��"ϑ�^��`a�h{�osr�\B���@�H`�������Evz�q��tk����@���l�7�Q4��UCX��N�2f�bWѼH7�a>�y\]��cģ��D�R�d]O�70�c=��	ݓ�!��'e�Fvsm��������>���������L��`t���Ŀz�?�V��&�,3Z:��O�Q[��7t3E"�mې���E�K����� p�穇,W�:��+��9��l���F͝9�a�e�;&^A��K@�B&�hͣe��%{���I���+A/����}S��pi������aG[&���:bq`�����n/j�$fՉ)���a��\��1H��" Dz�F�Xa̎;�j��Bǃ�&����8�g����I���A�R��YF5�k�`\m����ma8�P�3@�e��6!3,�N$Qo����zȔ ���8X�ů�%E
$!�[���mZ[�I( ,��X`����*��JF�F�BG�
Du�^X�0N"�m�D|�z��C�i(t[��Ͱ&Y.��,9�	�� �^!P�f-�Ʃ很�Ī��2���u��KY��4����"P,a[�:�j�D=~~������w��g����٫�s;_��z��n@}=9�t]�Ө\�]�@��E�ڕ�r�k����{H�<�Vڽǽ��q4�p��Gq�u-���@1����n�����o��6)���i�uE�N�Wmro����h��sgy�6�ų`I�&w�c������'�����6�3n:2����N���w�>����._}Q�VG&�d�}FlfE��v���ɘ��݄ld����=� ����g����&����FVe������!���u��P� �h�5�[�i�9e��7�����ݗ����g���Zˋn<���m׷n.&믦{���0���ޫ݈��יq�t�Tfvov��{ۉ���#�2!fO���=�wO��������$3�1$In/\-.�/2��7�5,���_���j�؅��9�6eh�b$}�%RLT%v�Iн{{j�H{V�z�+���<_Ȍ��Ի�`�K6n��2�Ѻ�F�(�k��^7B6� r�T�s����s
�"�⠷[V�T��Fm+��
�K�!�4s��c�v�p1���rJ�&�Z��ehU��������3�ex3(�4���k6 Pg�s�:���uUכ��ڮ������׃u��K�dK��s�wM�����j/X�A�[L�m�{�/u���x̩:��[��o!��3�}����ҫ����e�6���в�@j6��2�z��9�;#�C�o�:׮y"2�J��9�&vZ˖@z�g���ם��}�|:��(��d9�񃣰}��M��}�5ܲ�N��Y|/�тVX��rB��� g����7_^���N��e��C16PnW'�9&�`�WW�ӶNvb쉗��,��b�)�$�ɛ�ؿ�7ي�~�!�Fbe�6�DeW��f�o:�xi�ػ9(C�e��M�0�:�A�6��aH��/v�!�&�3+���ؕ�֝{�[�h2��Vd�c����[��0����1{������:[�����=�V\�ysk������Q�DL^��.�%���񼹻��'���nj��E�Sq��f�.og���ӣr�S
�e��d�p와�:.��9���8co��ҽ�߽}��5ں���0��/-�0�)6 �!�9�A�M����ފ�{in��|#�sm������{5���=d�����&����#b��p�o��os�����iԚ�BH���xq��=ik�������²]��^R�ef�39t+�f�9ջ�e}�����nV�m�������)�gd���L��.b���y�0K�ɄCk�"N+c��[ă�P(����y�]y�k;5���F����so�ȱ3[�[�}�4O"�u{�f���X��E�͹흲xiNm;��Y�	㝻���Ѳ�r����D+	l�ZgΣj�o���e��3�-��#�����{�|ȍȡ����m}�\%S���z�:I:_����*�E��h]�vE�p�Y�ZR��6��,��$ĳ9�ȉmI�ػ9�`T5��me��HT�@兵v���,�Z3�l$�u��R���-Vc"�j�*͋_�y�`�a4B:cj�u�qur�͌�s?][m��o\�OY9jĪ��95e��̬���L]ߪ7&�o��o�V�϶KO1Y�pd�qa�]V�g9�{���1�nP��Y�٭����'��Ś��=��qI[L��n���Ŕ�.�9���v�ad7��Qw�K��0A~]U�E��A���A�w���������4O)�9bp<*k�V�9*g��7����I���kL)bqF���^"��*pER�r?x{������5�}Y?Y=�#)��hq��4���m=�ث<�7�q���8am�����H���5�U�}Ψ��[��r��|�n�^��9������{��(8���>��S.�m	�	vr���t{��m�c����j�g	h6��#;gOi,�N����uD��2fsFt�Ǭn�l���1��'����Cp@�oI(���Sˍ$���r{糦�U��������Q�n�>��Ͻ��2ܤ�B��e�r�V��y���;B��2�m�1�Ae=����TOxi� ����Y�~��ZZ4��mX�TH�D�6��,B��75��Oz���ڛ,���{�]gv��C�n�ϛ�w!��SXS���ۆ�����T���s�'��m�=Gn�
�8[��ާ�d����ގ�|h|Q$h�)i�{y���O�=�q6_[���G׸{�{�,�6��}M��z�!v�eV}x�k}}���Y��hB��i��� �b���/-���U�����H3�f&��w��2�u�T�,6��QG�K�S]}<����6S��3(am��:���s���7ùm�r��Ut�CA�;[ۼ�Ὣ`8��F�,���I�-ʼ���׽d���C�����߾' ���q-ȭWAT���joNq,�ڽ�2��ʏeS�����ϧ�ޡv���sۯ�����2�Ѽo�Q$�5��>�s����l�w�v��vdS����������Odp�n�Ǟ������OsǶ�:ŭ[���B�y��ޑET���ڼ!lb�2�V�\��֮��ި{}ހ�9�����|�t��oˆw���p��\B����O�g��2m��;�e	�J�ܼ͡�{W�3K�p���a��iw�Z���
6�V7��C�g��L��4G����WJ�WNvL���1�{�_Q�po�~T�k�p,���\�*\V�1n�g��)Ax��������%�d������y{��J�����k���F�x�ui�Cv��ކ��y|�o����7���ߦ��O����_�����!�"��沰�Cm0�X1���)�`���A�XZ�Ɖ�3���e�1t�޺�g]��^\݂1[��,�Y����Ta^OR�7��I�Fˆ]h��zp�`!ɋz6n���7Wg_n�޳�	,�cBc)DF&"a1�ڍ(�ՠr�m�j5���3(��G[M<ir���d�S��|��Ȱ�ZAMz��a� é����I�,+J��W7 ���K)X�d�� [ԇW�f�Fʤ(�V�m��i�c`vRq笄�U�N���"�:Q�� �++ć$Z�JF�!V�� �d��>6zX��m\��2�3Zb3hh�q���Ks��B&����^�U��A�ɠּ�^2��MF;@���Pe-�3Xk�j),��7e���`0�1!r�s.ە�4�%��E��[es�a��
2�fg�(mK��Jв���!��F�cXQh�Բ�3[�/j�Ѻ2�!XJ�W4`��0q3c�lq�����)��\�+tm�Ҵ������D`�<܌&mK��׉s�0�pQ �I�������ݦ�R_�t�:Z�F�l�6���m��%q�a(�͙�v�̛l�
P���FL����串�ٶhS���u�5�*��V6GAK�c7	u�4R��j���4�;�dHٮp�ōv�\Ԕ�\��2�Q�Rmu��tA��;���nBYe��	��.K@���[N1�t�t�3c`Y\�P(u
Zd@�%�n��[�k*͍[Kİ��".�[���eq+�pܑ-`bK6̫nKiSM�kе�yUm���+Z`������b��-r�*e�sVWf2ׇ-5[m�.UUPfY����m P�ح�)�&�p[�;�����g�OZ�p�/iX�2�1�`���蔢L��InXl�:-��J��!��
�sv��l�:�[l���!H�ll��苕ƛ`V��۶�j̐-�����\�+p�LZ����_�Dm(.�fGU�$�|��|�.|�{���Zj1>���h2�qQ�]�f�n��y��h��MV�� ڙ��5y{6�N�e���٘�6��my��[y�^t>�SF���8�b�Ci�3�lE�ooo;�xi��ո����%K~,f[�xM����"�ce�ryJ�!���˞��'��հ������.�7�|�đ�~R0oϡ��f'#;)�uY��Zor��q$8p���ȩf-^/�����������?C��0��Y���m��6ּ[{ۮ����ڈ���M���ܞ�������nY�3���l����n��d�>�^Ǣ��:�3��{���L�+�.3j��́��wy:��]y��>�%$Ⰳ|��%���M�5�q�!{={���h���}�U��4U,q��P�ka����a����ȏ����kf���Su���56�f���<�+s7�럡����C�*R��໥g���3��������kZ�SeK�Gmr�[Sy�s��h��d�7Ԯ�� �]B�D����yn�J8j��!��"�h5o+r�z
�:;�Y�3���9J��D�wf�'��Y�M(�v�d6��m�%��8��H�p�d��Axj�USW�o����c>���P����}0����F�L%���������|�7��1�Lď� {�S����ow�z��d)ڽ���m��!�.mK�m��p�"a�\$,v��me& �*:|��τT�q�O\�['�6\6��%J����5{���{;�RsF�
N��.2ݗw9W�sh�E�יnt�A�E�ף6�q�O\�n�q�3e�d7n$-٭썷�;߱���������5��5;�9J�%�`���q#�f=7�����{��n�B
N=	A�,.s�X�
�ĺ�l���)+�r2��Ŕ���ͪ�K�Z�YQ�;����u�ih��:��HB`+T�݈˳�xI�1�"�CF�ͺ��Ͱ�1]�۽iml���宎Hp[C�� � ڙsW�ݓh���P�n{����G��ٖ|�D�v�ޞ�;�/j���{�4�NC�3V����}oP��l�$v`��a�#���gvM��K1�Т�my�N�NUv�Ν�xq�^e�t���1��1���UԷ� P�o���Ϫ2���r+_'o��������]�|��߄��;�V��꿙���X�.vF��ӑu�TTYV�� o��\��_}�h��-��jx���l��U�Qݓt�'m�rW��	���+02���+�'�_.}�j�Ŧ�m3���B�̾��G��m���zw�6%����l��T,-%L��"��$�ޮ�32��r��������u����fFj�4��+��7[ٕ;<���3���F`p����-lkN����ƃ�F^�T��sB -Kƛ0�FhY��ˉ�� ӕݛ�V��6[pϧ#��۞�8���o^�Nܞ�t�s3%��e��\t�Y�]�]S�|�4�w5�/�h�j��Y0�-��"!�C0�a�A�c�Ǚ}<����mݳ��L~0�a���eG�ɰ�ϧ���ϧ��O9/�[pnU�Cn:Z6we��eODw�����dt*@�T�D�^�u�#�ߢg�h��z�Ne\T��g"��}��Ǝ#yԽ��aGSg`��T�=��=⫗����i.�}3��_Oӷ'���(23+���Fy�7D~7J4��-F�0��o�J��_e�T�FuȮ/�(6���I�:����޺�s���]J�!�>�M��v���n{�����&[t��*�M@eV]�et�Du�B{}qRb�p�{�S�n�//k�����i�~SN���O��?fE��7p����#6�\��~{��F���F�tb�}�x{����A|�Ee���G;CL���r���҆llеu�h"���6���D��E�ؖ �@L�#��8Q��$���-��)I�4!2�j��#u��p�Pc��f�uqf��"^����� ��;&�j�X:ĺRb��h�{�<Ӻا̯�쟶��kj80�I�S(NzFQ�")z�����ٞ��|���5�1v(��6:wUn��ڼ���Í��ѭ�����]۳�WG��C��]��qm|�h����72�g�+xcM�p�Ө=zn�����ؼ��#R�I�bC� A�.
gr�:����蛘�W>e�6��o2!�up�1"-�.������Q�$F���x.6�%C1�XN2dƬJx  ��Q�Yݳ�U��ʇ���]3�ȓ��ΕTd�}9�];Q���䉗�t�P�q�o�/���5�`���^��i��%Y8��`�Cow��{������qܟjb&!tܡY��V��ă�,����d-�����F��:�����6����2�b�콾���Í��hCȫ>����|ۥ�)y�-N�}'�k��<�qk�ܦ�@p�.�SݵY@�t1� DM]ݛ���g�DkО%��-��jIc쮒�mR:'7PR����j�/=�+݋��5ʐ�r�l��@�^d�f�KBv�7��M��* e�h��;f���4j�V��g����C�>Αjx��4��4��nb�و;�[u7snK�bq��{�S�3I��"������G{ѱ�K��f�L ;�5����-B�u������{f�̜��s���pl��TEݛo\�;pZ���{����#c���6�'z�
��#Y�4��2� d�m{�4��`�� �ز{"F�2�0�;=we�Ǻ�E��I�{up�w��λS�x���-�/l�'Y�gl�H���^c7E�+g��.��X�zg׍��>o�v�Y���6Vŝ���� �݆��E�TԹn���������0`  ��8TDD�8"��R�舐�<ʇ���EQ��01/�R"
0X$� "�� �"��`�0^B+%aB�P��sX,B,�%�� � �1�B1z@*���A�0%l
@9XC�֚*�!D �p����+!	`Ă��"�:
tER!�-B��
�G���"�UB<(ÎE�J�V
��AV#ブ(�$$�P��ǴE5�WZ箱�g�v����&Y{�',��my���ά뤻��q5o��m2ϛb�;\	�~·s��������"�Fez��9UH'��QQ�m�)`�/7�kT�]���#��3��7k���.Q�fr�>�'=��&�a�%&B9������t�����J�Yٵ�t�A����=޳�ls�X� �k2L�� ���F7��+��K��@�-�K"H��<z�-j�>��$j���������}s�:6���Vg`͝�S�9#sX�ӳ�3ijr!^��ae��9������,>����%'�+}t>B�#�~[��Y�Kr��Ϥ�d����O�:#�:�ƶ�t�0�YJ��	�1���K{���,��"2�����s�7=�7j�,��^�˂�BӲ�����2�`��=s{ەӷR:Qe@�E�4ER	+�� �A��2YV�3y���t�G	�@E���L����!]ґ,�h
>~�Uf�n�U6��4�p�x���zua���L�>"HFH��o �,���wk���#�>�@>^2���w��뿳&3��I�C+stc��ko�*�لܼ�2�	��
��*2�v3A�[\�)a�T���6��&���3���hU�˲j<����LQZ��hCG� � �{,�piE�La����i��7KrbQ+65��33�]5�����������k�[4�Tkn5��;%̷{��@�O�0�����v���#��(���؏�d^�L��@^���+�׽X8����n�svw��RW��9+2y9fǌNJ�<�-^��t���̺���۩� �D���(#2��u��:}��7* ɎU��Y�kr�!-r�����5}&30�$k�뽜�Ԟ�O�G���KE�K|iΗ5ie#G]Wn-�3KH�S�v�1hA}'�(M*��������Y£3��zx�K�Be@ �(�����:W�k������.���!�hS6�`��j��k:!��kݗG�� ���( �(E�o�mo�kr��w�f�7�Zd���!��R��u�Z��+��H=�0�fT	��
!��6)Df $46|�`Q��ܮ�ʐ���"$�۵{8 �Ax�A2���"PFerj�a�WݙY�kr��A��>�3i��D���n. O�ĺؼt�#R��(=Ϟo,��p�/(*uۙ��U.'�,Ui��:L�J"R�SV��v3��Df�ƫ�r�w*B>����[s'�!c�>BPFeG�&O�WK#�m�OZ'�����5��͘1�h ˞�'I{2?x{�OnmoM��	�@Yq��Xb-���Q�&r���!=�v^l�T�K�'J"�먛u���ԐA��>�@2$*w�muoB)�ٻ�]=�!a�2��D��(cժj� %	�qvcð9�s5�f��h�� ����e%j���ΛXcRg���=���13!bcX�k��@�H}V��[��;�0��	��"��"���p�!� �! d���"{++U�W}���R�t���	>r�3*
�s��Q7��:�3k���Yݵ���\���#�<�����&oo]���@N��Pn+��uS��UcU�-�YX�?{�2>� ���/ID�D���EG��_�ݻ�0��������G=��#.�Z�ER�ե�.�A�QY����7ٹ�zO,fJL�ƫsr�w*B��!p'�x�g�� ���@L�A2Q
�H)�`�Q�4c�nn�gY��z���>��@��YD�I���'��vn��K�����.TL�D�є�� 0�8}2������ܩ����P�16�h}��2���|���͏H�l������8y�)d������̾�l���Ɯ�x�A*~ZM�#�P
Sc*���o=RY��"Y���'�3{&�Z��MF��e{0v�m
0�*l+A�����5)�r�+5tM]n*K7p���1�p���T5C,aIkf �le��6�`!��Zj�#�!l��TV�m�,p<F�Z9=����R�Uܸv���l�q�A��M-��N��D��!c��Ν�ip##��\YG-A�DI�^o�"�{�f�>u1U^��ueH\����<��O�ȠnV�a�/U&���ٍڝ��8F��z��ci�L�	%��������,�H�u��ӽ3/q��<B1+��L L�2�'��X�B��J�;[��=�u!a�\-x�CQ�\5R:�:���Y�l�eb�2�m�]mC ܺ����ol���wf�u��R�v��Y����vN�nu� �Of`@"R�D~���*#>fj��}x��:�����}׺p嚺����L�KO��S�7?T���>u��ӿL�K�t��c�4�[�wz>'���=��d����q���f��n�"8��Rex�^�Lʧ���FH>��@Ix�z��Y��/W #w��ۂ	����% L�D�l�ǻ>��M�M�Nt�4�N�A�3* �YLZM�	��Yx�\�- T"&h�����B�2|�������z�B#
"0�E[�[�}��H $�e2	������X���Ӱ��k2z�}:���{�PQ�D�D��%��=Ӕ3C�U寻N�A1;��S�MÝu��
::M@��Σ`)T
������x #jj�'zf_x�O� ��PA2Q�у��H�:Qf<�y��z�B�^�!���$�5�4�0D�G2N��&�ߑ�S�u�=g�	�@Y%���;s2L���ȿCa#b��٭
&�Z�����|��m�"�v�l�:��Ӄ0���]�$��� �U��S��}=u!Ǐ�ʁLH28O�k�)����0�2��sKu�U�=g>�C�B2|��z<D���a� ���)�(-u�yӼ� ���~�zL��;��i�fi��C������C�}9'N�Л˵��nM�ٶcn��V���P}�)ze�&涍�B�}O��}=u!r>C* ��%|����Fu��&!��p�M����4� ���/��A�#��S �%s���ݞ��~�웿~=N��#�e�$i��ɫ�� �>�"�wם;Ρ����b��b�E��"�^�@D����A����Ve�������ʁI�3+��l�i�IT�v�g��GӨz'/z��y���X��5y������U��Wu�9Ρ��x��e@ �2m�ӿ|���W��3� �M������$FK�Zm䏽����߁�25�Ν�T�M�>����-΄���ƏVy��fc�=��^U��w�F*��^{}��5�ݾs/Lz=!�=֦o;�=j8�<��J�;f	�y�t-w�����oۤ[��S{�bU47f��<�Ow�3���ڄ�>��d����F���O{T�
�޴��}s����|o�<3|�ӻ�l���	�q.w�j>�J8�X�$iVWf�Y�|��dҳO^������e�+�>7�g�}�����^��ܷ,�z����<�kAw�m�p���������
���3`鍠�7fg\�ك���Sl!Yzõ�Kn��ɪ���OH���ɦE��~����`��3j�1���s�Z�3�>w�g���Mr���^넭G��P�2�xȢJ@VE�4�c�"�PyXA��  �`�b�
��G""��HT�a@P�b�ˢĸ5�F1���,`�Fb��-�Y�ሄnΌL!PR�UDbҪ*����U�%�hP�q^H	 H-%�p��� �p� -���@�B˲�r�/B,Dl�b
+!Z�hJFIB�� oXYj������@�Y�(��D��$�"-HFJH�=�>k�}�� )��8����mJ��,!�)�@Ѝ�K�j��	�����*U��nͫa�f�X$lK���]y;\��քX�Ї5;�Ћ��Y�y1�r�]1����@�tMsa+rЗ`X��`DA�V�JX�Ck�p�8U�$Vƴ�ö
�6�4X����ؖSit�aP�
5��G(���sq�nQ�����=s6�W9�u�G���d֑�J2�C5Ֆd{eW�Z0n���k+���]��f6�\+[f�efll�&�Ќf%[��/Vƻ2��(�b�`hC���H巘&��Z�L��׈k��H�+S)v�p�*c΍�7Sl@.Ж��H��ad�J�9�ۮ���6����R��.]J�0� K�2��[bBhJ�˓�'dVj�D�M��P����Py�L%؎���MZK�� ^_m}��Y����l�i���Ƶ��QL ��,���]LF����;�m�U�ecv�4%��i���6� au��i�^d���i��S��-��`����v"E�fu��[��B3*��:�:�pM����l���\.n�rn��������͈K�Q�[P��eN��b\���]x�0�b��u�X,�b[�" �v��E�nr�RlY�`�!�0��#s��-�v��[z��GR¤#�<��X��Z�Ƴ?�����k���	n�ٚ�;M`MEf�����~�-�O��}Osu��ԄFJ�0y=lG^Yi�JƳ%hi[����Z��͵W�[��p"8� "פ��v��@�>�@I���dr����t� 4�FeA�J"H����ڌt�� �L�Q�ݳ;r��	∓1��UB@a��̯A��}2�2�dA��K�Y}Y��p#��2}2�]U�Dz�v�=�=�U�њ���7
��$��""C@�>�@L�I
:�o:{�'�1P� ��b�(�K�(@#������|�������e޸�;�5�6.{-���mY�Ov,�4Cy,!u��>?!?@������3�,"8�D�D�F^-�����%eze?L�,N�3k2z�����&�B�%�n�������(E��gOk��{���s{���ǧ3(��G>���k�{}��;m����'�J罰��);���n&bU�m�KV��m� �����{}�ٯ]b�d�q[����p.F�y�k�}0 �AzJ!)��b-x�B6�+6{]'�x� �����b�Ar�(#%2���x�R��`}���DF������;�����~&����0�%��;s9M�˚����ssfz��O�t���%fT�o����(��Ge@>���+�����|���¬���3vX��q��XfV�������v_l�;N�>C�S>�ӣ��g����y���EYNl��@�7�6��Ơ#ֽ'�3S��|���/�r�̲�7� �K�W�S ��@���׳�X��A�Pl�0.b�����`\�I#HFND�ި!�@�5 N�A0 �K�P.k�ٳ�5�p��,^�@I�$� v�������@�&`<���|����߳�韐s��O|*b�����3��7E�O����u6�y���6���v����>"O� �ʀ}%x�!������Ϯ���`\�3�APFJ&`!߾������V���K�r�&�P0�n!��4|��	(�('U�y���8^9z�>�H	>r&e>�=��h��ռ�{p���n�A���~�^�^gJ�T�T�����l?�v�j��|��A%f`@"W�4j:]�.W��꽬��v�.�|�͉ͨrW����L�$^��al�^#2;̞�}p�,�>�w��>��15E8i��~�(��^
�e�ǔq��`o�)�����6z���Ð�t��������JM�vZ�]�P�4���9�i�Jڔ�u�,�f����	��0Tt%v�Rjg 4����chi�]5�KQ�Y����l�37*�b�������!4��D
�g:l����e�;��&�"E�ћ]��qr���>4QB3*>2W8����X3�ɹ��7�kp��"fYt�%c]�w+�Z^2���y���8\}���+�L��L/M�^�虀���N�";�0�A��I��L�vD�e�f����>��u�]�]�����/P�p�E�HT	��5P��M�ؠ$b�][���8\'��/L�A3t룟>{��s��ڑ�ֶ��[����ޏ�||2��bx�y�s����0�!V7`i���>��4��A� �J#�3E;��#�1x~���͹;���C��u;�aا��P3���Ż��C�=����u�e���`\�9�Aڽ&�2gd!{� �H�5H2+����1����~۔���>C!�� ��}�ч�0����޷{�c��}���"��@�(�^�L�(ezeB���jows:�p.^�E��J��̳�����޵�.�F�gZA�� �#�v+ (:^���� �Ax�
:�/9�\�����ţ8�}ڛ^�B2��;ni�}&�n=۞�1�J���Z��b�~Gً>BP@̯A� l�
��(�@�=��sw�έ�4���)2�)�0�ȷ=ٶ�f{������ڻ߳��#㼀���3A7�m�a�Ay��$E��n��i��<P>Zq��;�3��8U!P�5H��9�ۆrn�X��5���P�q�J^"P�yZ`S�5�44�7�p�EXC\QslX:#�ݹ��u��5�P\dW^��U�EܼFP�/i�L���2QB��[ i�����#r�i{N���S�\wU�>��h	>�$����s캳��"4�D�_���L��6�ψg�h	2"���m��`Dq�@~W�>��(��"m}�M`�	�����<y�-�c9qp
�^�-K-̡5��>�����>S0 ���ݞ�4c��3_u���}��}2��8S�ޟX̐�nAӈ.xf�JE�Eg��e<в�FJ"e��lwR���3�n�e�#eG�D���}������(GMNwV��X]�	�B�2EM��ʨF���A��'�P�5W�Ӗ��H<E���^�d��#����A��A�[���"8>kz2�!�E%�1ze3�>R�2�[jP�l�9S{��7Vy{�}&O⪠<�o�&]5�I)#bܶ��*�����u����s+��]ku�Q.�*����h@��)m�.�)u�Q6F�����3f۴[H�����捕&�fDf��M�WZ���.,��4E�
M�%�F� �$ĩ-��ծkp�A�oT$u���7u�؈�g�w�M��U��f�ͭ�ee�7j4���;��n��;!gIzHQWy��z�4��TOu8,�٫��DI̡Jfu9��"��h�����L�Uޗ�#5������`c�=M�+��_���v\�y�'�0D̲�1=3�\�<NbEI��o^u8i8(��Y ��QBe�%���:��ѱ�p	x�
�D�I{k"r#98m�F)��܉7W[�r�D6 $�O�XA2SyS�ӽ7V!��GmI�@Q��("%��%?<8*FOwE�Ʀ�T4G�_�.HU�� �����U��f\olV5�x��iE��f����OA�3(�E|�j��MBW7D�X؎e�5����746;n��j`	ax����S}��qs@2Pn�{:w���>�C�B4u؞�i���%�A��(	���GF�u�OSm.�PY̯A��Z�3��.��%7�NE�n��p�Lй~��4��ބ���т&P���s��u�$q�R�p�U 4�%ze'��s#z�q�^�ž�}��7VO`������Y7����B����\��D��TE�3��?2!.7sK���x���/�}����ܧ"���;��..�U����S�u��x��K�Oi���Ν���jRD�
?/*:])��Q����o�d�a��I�������R!,mf�s��7}7���*B�CɨS��ɾ��M�nY���;��O���:��`�E�����Ǳ�!�;�!@r{���_C�;���y��^#�N�t:@��3Y��a���I�C�4p�8���@K<�y��$_��n�Hj�������ݲ4���7��e��d֧0&���� :�E��h`��p�?F�	Q�c+T��Ѧ>[�s��Py�=�n��W#Խq���Vؑ(����N*��`��ye��y���Ց�i�?v~��{�ڜ��<'�7W�rY�\\Н��lj�/|2A��Ė0KK�ij�d$a�'�ҤV	��È�ci$���]ح��DE��"B�$�B\%�D�"�b�
�*�88 V �-^�R�,2�XqAX'�,��X��
��$�!)DQ#1���JTh�A������ (�ZE��#Ȱ!�T), �"ǂU,z*ղ��V��%xg<F�C�a�E`�c��@�pp Kn�0I" �d�K��](����Pe�6�-�YH��@J@"I��3�ޝ�����i~ �>U�G2U������r��Jx��V�ё�p�>���7����di� ̨ �(efV?����b�7~ٽ�ޛ���! ���}2���&�2{���#5�5��H����.�/�s�X�Ԭ�;�s����m��zz#G5̟\��J�AJI̠2瞛�$+�� \��h���'J ���#�,`N �b�
���X>a��1��ݷ�?y�p�"��-���̅��ް�y��DEG���e7���vz�i{�G�C��3yG���i�S�n."�,�;sIQ���e6����|�vm�cg�����K�(AY�&y��T����Ӛ6;�	$q����
���JΪ���#����̻i��-���h�Pp�R@q��L�&J�N�N��X\5|�S��BH"פǁf$$�2Qݖzvg����>� V�����6��k�q,s'{�׷���;W{̞�虁��U�]�p����$w��!S I��^�%�֣vl��#���Jojs�w�����rC�8�a������$�O�BA���G���"���'i��	��h	�� ɚ�ȞF��ю����rc���Bh�Qn�9ɩ�Y��&�l�<<��F
��!�J��Q���GXU�s����lse��u���hI��^s�6]�rY��8�������R�vz��,����S[u �ֱ�ea�B3J�"k�T������:L�s�￑���U�4W�����f�ؿ�c��,�d�e
u�1���ǜ&O�n@�,�J���2Q�	��B�^�%7�=�;�uap^�B�?�G�_�S�l��D d�&P�D��$<�\��罵ۓ��K�p�Z���J"H�\M�@���4�(#�D���y�_u�$q҈u#������O�W��@�!�cX�����sf�����I�A��KUvL$�-��z�Tn��6��tJP~O<̢�'�	A]��fl�Ciq	���F�#O�� �d�afP���������m�_��Gϖһ�/w4,�ol�qE���Lt��<��~����O{����^҈�@M�ȅ�^�B���� ���g�Q�+��1=�5s�7V{��F����@Iq�v��� �^^2�s}ٛ=P�^�ҰIG$P7H
,�Aze�2vz��f��;�;t��H�x�� �>R��TDp�^���cb��cu��UB
��U��E��ʃ�-�<Μ麰�=��&s��4��L�&P ��fZy>�Aٽ�͞�m ,���L�=6sT�!˕�B�0D̰��'��A����C�s��bӚgrK���j)�ۍ�Q^:ͫ.π���=k���`�a����IS"��p|����P��t��s����	�@k��Yf�R�4Q(A#�Cv��!ݵ�w������L� 3�khu�S�s��rFղ�gX�0´�� �a���ր�^�虁�Q���m�H�"�Aw��$,UI�4W��u���՟I�3�9�N�7V�܀���g�s�2�c9�O��4�Ư�/g�K��Y����>���Q՘� ���S\�rm�H����\��:nT������N���SI�@�[F� ���w��vG�Jk���KE�#���I�}yz�ꮩ����Յ�܄�#'�L��"���wɠ�ٔ��q�q��Q!�H�G�r ��(/f���l�Ciq��˦�͐F��nT�($ fP�Cj�\(��Zl��n��l>�G���5��+�kIm�Z ��g�Ό��>|�{9��^�y��e�מ@����fC�r�&�K�&5%�7�ٛ=P�\���"A�^�e+��(��=wJ'&�
��y�]�w[�n`	k�A'v-D�\�\�Ɛ��wL�rsZ����#@9֔:��v,6j����%��x�eƩ���[��vڒ[��+�I�p�8P�H�XQ��́�H��ي�mu荥��-�l�2���1ɋ6%��̱�H�(CK�y�i��Qa�t�V\L���}�[�;e�:���M��a�h8{�{���h#2���o*{�w���!�7P�4�p�e3��>SG�J��Db^����͞�m. ����eGm�&�1Ӭ}P�v���>��|h��m��r�>�A�+��J���a[�(�+�I�IM�mwN�]XDq�@^�]�ǌ�$�k2oFcs+z����������>� ̨>�oa��q�]�ᕛU�D�]X[�Bl8MClN Lb����B*j������x�� ����+�(	2Bpθ�|��N�;&�F�R�ط1��C�����/�P�z{���+�p�겷������� yd���۱���H A��5P �>R�ݖ�>�ݟ���A�"�@̨���I�HH"�FJ�9y:qvԃ��Q�R�:���"�^�(��ǢU��1��w'7+:zjh-@�� �9d��|Yߞ�|�fHֱ�nڣv���0�A��b����_��;�uy$H������m�����U�P$�5{%y�Hd"�y*�UP�ϓ�WW��WuH<�8P ����Kޟf��Z���8Ce`���c�rw�yE��E-k�ܦ���T�F�,���h�� ׵Sy���6�]]���Յ�{�����|�X�2r����G��bG�!E�����6�O}w¸�4�% A�@D���R��h>��Ӌ���|�s I�/2:�p��Kp�N�u3��D�j��,��$�O�CO*g�kwk�����K���8��[m�,L�G�|�s��q��#��orz�iq���e	���:��>����1���=�zQ����ǋѸb�f)�*�1G�G�ߎ5��k�����rFk����.gch���7P�b��o?LX<'r����>�C���2Q(	x�h��]�]�n��m/q�"�Fez�Ʉ�o�e8�e-�[�3U�h""C�Hö����A���y\uwT�}��*�dp�9^�L�J"�,x\�㘠�p�uӽ��uaǹ�&br�nC��@�>�A�'�F��0�X���p��|��1j�QDJC�z���B���&`Ggוڗt�N~|��Y��p�~?�l�0F0�YW>�2��7'����'";�C6Q({���@1o�ld}�MLM@���\���ݏ[TjP��&�j��4B��qn�V�с�l>�m�w�{�L�pwN�ȝ�f�XY9�3�r2�����g���:����_���-sJQ^�^����5|6rj�?L��.�t%v���s���l�WLp%�bsh1�S/X�7VЛ�;��N�8�g��7�
_A�H}�{��^�����p���b̓#',���kG/=\��h���cIbu���_˞}��xNۀԆ�^8�!j�D��Kƙ������v/V2�J�)׶�ܙūv�՛3z���.f	�-wwUkH�̫��;#�\n��jk�I3��ݚ��F�$�\�3�
�IT�9�Zɽ�TT����I瓢<���8�9{��0�N�،�n�0�2cj�6f�=ٙ���F�£�B(N֣U�`���-��Q�h��7���"��ZcwQ�a�X��Q��Q�Y�@�+��0�<��)"�F�
�#V�2EcDTW����J4JNP-�F��(Ҍ"u�Pus3%Ib���رQQ)ń�R 2�������%���Ys-���P���,H��"A'"�A��B8�kZu1=yď�XB08yx<��@	�YUXIH��( ' U�ռ��H%|D�� ;,��kF1���t�2�(`��)V$���f%�u�:��o�`,���u�5��ff�rae*MQ��Ҭ��6l��qe�J����5��KKe
�D�<��X�"id�\��R��ؙx&�y�-���p��f����x�k�\ƛ�Ezٝ�.X���xV��Ti��$6�n��h���T��,�cK�VgMX�3T�U7������V�%D��F�m�V��L;s�#wT�0�"l�4ƫ�GL��J�1a��Z]1N8,��5ᘵkr��`饔�Q�Ћ�]r��X�I�LB�erJR�&��0��)���[�l��-�-��L8r٢��WL�;i�w9�L�P�Gj�.cKft�KP��[�*8�sa*U9�t�Ű�Me��+��|L�F�jH`��K�=I����)&�bb���JF:ۆQ[R��j��V�L�eX�F.wb�!Z�2���%�[�-�f3͗R�,c	��e�����16WP&Q�Η/	�\����ja`���+Ò�����y�]�Xr�ٍ�5*�@qvV�sZ���*��9�[v[��`������C��[�=�ۧF�Lb�����S`�[��if�K�)�m���٠GUGi���֭ųm*�*mW	�0G�JLT\�lp�9��:� �;��kM0T�m@f�.�.3U��+B���>�����(��ma4�yc�R D4	>�@I�!v�m�9��.#�e��D�G\���L�G2�Υ�8|� F�fV�]���	��(	q&�sF{/n���'�)�Iuu·G-ۗ����uar��I�&PЩ�Y$� ��ļD����u�K������S�^�@Q�D��J;��vU:���uv��L8����'�GL{�w���澶]���̴n�+��.�P�h菾m'w�/}��\�}�z��._��G�`���I��5�\�K��^;��E��zn�=Hd�"C�C�q��U�)]�.�<!*dGP���1����s��.>��-zeFr�m����!ă��h�+L�K�߷�\�+�.�`���70�I�kڣ.� �6�A�wg;'����	�@��y�c҄�� 
!�G�(2%�m���ww\��K�'� ���g�iUkcIb�e0XH��-�f	-�2l.+�g�����gw�Rf`E^�V�]����{:}X��^2�2���I㵷S��p�s�[�=WV N�F���S="�`~"��eT�����N�?G�o��A�7*TH��3�g:�`Z{�oI�G���9�a���W���n��N�B\A����K"H�:"r���(��f`f�d�%�L;�,0F�=����8�H�2�O��e��eM]�ol�]XG٨>g�3 ��G�>�>{>}P�)6m��������C�藢�~rV�"{�,Ljw��=1	q�v���Y|�&H��=��n�W��AɁ�y[�oK��D] '[{
����>�^��efTx�d���j��ڨ����꺰�{}�~B53,����k�mNC�d�����˟�9�W�Ά���CZ=�}�Q�^zUT��3��DU=��é�N���#f�W��x�
"W�&e"M��T����[,�>�_�����Ͻ=߿e��s]rS-Q�m�@	�HI����A�A���O����]X\�E�W1�a�}s00�>���R�aH�x�
+/�v7��$�p�3*7���{"���PFJ�bUY��%�r��`���!w��'�+ڠ)�ta2A�.�TNt���]XG٨q�>���#��h0D�	���B��K���x��W���z�@i��Y�`~;.�~��Ga�j����Q}����uz�Y�n���ù��ӫ/߳a����6Z��ƹ��lˆj�b�5������W�ƣp��Vf�B:�t�8L�K�Z�45�R0�P&!Ή	N5:k�a4J���i��)BVf\�4��&V�Y�k����-�gdͩ-�f�������[,�ܷ�H#��L��Փز:X<�5e��b��|Y�����ot�:>�~M�;:z��"8� #�^2Vv�<��30�9^�f�v�NjΪ��	��>�RA2Q�Ӑ�A�,�O�P�ڹ�Ȏ�� ��GwP��*�K�B�2���J�ʮ��ezN=͞����G��>>�L�����!<��[-��hnQ��!b!�u{
� �@|���n���'����NA��@I��� ��y��v�o)
3\�y��b��u���d)G2�gCw�U
�����ܹ��|��	����o�33�%���&�"O�Pp,SW�۷���a��!�#%&P�$��wGj�Q�ax�{w��:�\'��1��t{mi���3(	!�&4Lm-����s9�H�l�.Ђ$�H�I��I�@�Qi�·bf�˵�!�:#�ͼ��(�!��2TNV�v�VU��2�i��H �I�f`	h'ڥ�Y=�k�g�Dc���[�P�x�!����v�(�!z�'�`��4��v��u�*75-��N<��}�����Պ�=.
�ٯ�*;����8|���p������|>���P�{&�vWVՄ}��VG:�o�#%x�� ( A��A��N��5s�":ko�V��TDq��FL�}&n�5��*RUa�j�4Qƭcl��.+����6�jŠ,��'��0+�vc�0	
��l%:}���^>�����F;��<�{A¥�M�mt��\����I쭽3R����/i@�3 I�5V��}���v�@a�A����D����� �"�G
L�t�7vy�����F�I�E�b����MVs!8;Nr��WƩ3dZT����&@��"Lʃ�>^�3)kY2�ni�vWN̈́Er�@2��2�[Z:a�F��6L���c�a���0�H�0(�3 @"R�:���urOD�V���P��7ɤGl���-F�&//����������>��]�%�X��5���	A fW�2a舘�Tb���mt��G٨qB�X�1���gC+9�}��={9o]BK�'J#qd�O��>����A��"�Z��.����S��(�� �K�P~����hM��.�&<���S������z<���}�1�P�͗p����Q��iDs��R�9V�xjXhKbfn�\�a�c��͋6&R�]y�,f)��66*�f.��e�fԶ���p�ɪ�������*�qZ��6ְ�\�@��e�I��Y{ޙL�J����Ol�D}3)=�> �A+����̔E�;r���b���+u��˺ɥ�:Qؽ2��Zz����&�"�FJ ��1�4�7w���8|��	>�8̪!���Q�,��0A2e�_f�>����s�[R��ô��}�0 �>� �� �!�+���nvr�ix(��"�%{ކk/Qm�XR����"ѭ�~�H�d"8�Y@�FT����4��aҏ��DR^"PFe%�Y�b�����^��s�ytj	��䬙!����a���������sv�l�Dp9�!�#;1�Yā�P|Ȫ��7yoe$�	��"ʏA�dSUfp�UHYj����7;3���}���ʈ�V��CAz��S �%efR\{'�rz���{��#�r8�2Q(Z�3|qdΥB!��C�CJ������nwy��'�D�O_f�줒�Fel��&��B;��d�$�g�����D�K�ِ T���ߢ���t�.Ђ&c7v�e��zϞ) �����d���5�.Y �0�F�/��b�55'�w��QM��C�tT썘6�Jѷ$����ͥb���mr�4��Ϧ�^��`���wc��T��TOQ��G�VX����f�6�N�/ohzJ�w����'��BW=����{��"��2�����9��`�%��Rm������9��`�]p�����*YC���rOo� p����zn?y��鍀}�_f�lL��� =���1n]��/B;���nݝq�X�ԗ�g7�5�3���m�Oz!�v�a��_-���+
�Tc�Hr��������u���42�*e���܈��l�j�b�T��N�m�[�����N������;��Ľ��͡�s2�z'{7�-�{%���%���r>{>Hͦ7*�ً5U+`l�a1.��u樨`�a�<1�Ɂg��d`�G��h��s% ��P�Nx�X0J�z���mIJ��Ϸw�ޯx����BpG7��EZ.E��+!j �H�\F)�"����f�9��FU`C�ޭ!T��,�Д���G�1�_YE��H@�d�c�(� C:��b�V����$	L��`�j�C���HV@�q	@�����هTH�KWM�AdR
+H����*"�$--,b$�é	�)�ŀtR���36�v갾@���d#'�f �(���P��$F�i��T�����I.>��T��ק�N9
"R4�&+�6�;{3���}��7p�I�u�M��-�	Q	�(MDB�tђ�fI�tG���ϛ{y���e@ �%K̝��{b��*܍��\��Y��2���2k7{4&52�;{z�r�K���}�g���mD����P���)��y���R8i�L��WDԪp���s�
��^6��}s11�?zg��>��,�Գ��p4��sEة�s;�(>��&eęjh����ge�p��T���S<R�)�ZCh�����@cm�+5GEW�U4ڗٙ��"��{��[��qE�0�ٗ��#7{`���IR�;��Ci�7
a�/.�oe�p����^�f�כ�y���#�������nob3)Y{�rk{snoj/{��l-ww�xb^+��2̸���N(������#k|`�T��"|`��h�s qѡ�t�G�g�V��<.C���)�8��p]��sR��)�R��TˢB�Y������K,PhMeh�1��:��%���k��Fm�k�����V�f����y���4�b�d�f�#\A�"!8,�aC{�A��]U�-쯒�g&��=N)�\���=;54^��{�f��T�����,%f����im�;��yl�&;3u�T�o0�l�ǡ��˺�ս�O�}��\M]�YM��g��1B�«޽�ފ��Eۆ�2k�>}�S��0l-r�6ְ�TnP�ff�7��;p�f�����q��d�I����"�hfeձ�~��P�
�`0�g Fb=[o.��t��Oej��G��!��DT�(SA��­�/��՛�#�]�>e���eUu�4�8��1�ݨ���Z�v�3\�8��"]emj��G��cpΪ8�AϞ�@��M�LW�ٖ��L#�ܭm������r81r"&y����#����]�37��B�3ӼMwo_E�d>`\M��=%P**��R�^��3�ܛ6*���Kǥ���G��[L�G5焔��JN��Ԍ�my�B'[��u���ٻ��q.����O0�����L^���^9�Q������B��׈>R#(lCA����hh�h�3,D�ϟh�M���Ջ���rhN��fۆ@mG7;���H��ͽ�݇#xU �b���yB[t#���«�Ev����E��1�a�/�g��u�����3ް�ʙ��]��٨w6#r�e"E��\�UC5E#IH1�/n�D�t�e��,��nC�nw;{���U ϝQ�~;�	f"LB�C\!4$��$Dt�ܟi6ڽ�V�;`�˜��vz}dQm�S��U>����m�����7p�y��mY�o�u#�W�Y��ܜ��UC!�6�P�v*�q�}��;`��GKWB�a��m�vn��W|����#��qDّ�(�<3����ÎP��ws�����6'��|!�Y~<|� Ļ6�3]�e�k��,m�3����{!�:+n
7@����%]2熚V9��l.�Aqb2�JM��)��$�i�����e1۷Ra`+�&m�WR#r6�&>��]�<Ѹ��j4����@cm�+̮���n|��j^���r�j���j�;0��k̺1m�H7��s�}��"5�T�*���>n�zra�h=s�koq��Dʖ�GѶ.&כ�}y�n���A|�2/��i��I2fw�6�l�U��������](O�\&D�☄�k��I�z	�&P����U]r��F�r��Z�,���7>w��UG6�璨_���9�[Yܾ�B�_u�k&xD���5�{�����>�A⊜��E�!� :�{�r����݃��@Q����]C˂2U7;U��o����]�Ә0��w;UOE�S�����c�������=Frj���pa�P�B���u�a��5M��޻�/�8��z��l�4�dT Ӏ�v�#eг��]z������+�����wQ0�wq�����14V���zM�����ޣ�#6�T��i(:��z�oc�ڧn�o3��"�2l�hOZ�I�pnV�}��{y�p�3i9�)�3�ہ��ۊ�[�o/V�Z6/�A�D�}pC7V2�K61��R�.�C7Λ��݈c�ߨP��`�m�61���d��⧯n����O�H7.��cpr+[����֏>ƁhC��.��,��;g�;���E�;��WF۩�C	}wqQRC���.��R�:8uX�MU�[��pF����F����ﻢ;{`����E�糯�>u{���38ڠC� 3�>^u�k�^u�ߟW_R=�ɞ�P&�:hUҊ\��\F*ٻ���8>�}"hj��|�m �v)�u��7�`��B�>m7D�}��NQ�3Ϝ����G�Z���*�>���n��T�
��wn�Hц����/菢}S��Y��^�i��8��-R��(U �(��p�(��Bua���AzOщ�x�p�Sb���h�.%%��~��.��81z�cdu����*�
��@Umj�� ���D��P?7�˂^�֌�Q�( �҈���۵�hT�T�%(�����̰�դ ����D��G�0o�D��@q�����II�C�6�� �R*A$;I��]�Üv���=�~�)��`0�A�Br�0cO�01r���_!�;ut�Q�d,��UD��&�HVO�'>IC����0�=��0����	����e�����м�z�Q@�"�C�"� �hE	�l>�=��V> ���z��?��C�$�8^�����������9hx��VQ�}Ȩ!⾥?]����z��D�`��	p�>��f�O��LN[#D���ʨ4 �/�c�z���Qk�/h���U�c(1�|}��I��/}���!�k2{ύ���7eDP���)�,Qc������ 
���S6LY&)��Q��Z�##+�������X*���?NpF�xf@�����_�(� w(""�lJ"�DJ#$��i���#��{����ѣ�x�{�����U�W����?a��S!��W�������d�|�@���_��VOXq���g���@@8>��#��y�}���?p��H�����p��C�x��m��p��S��AG��|�~��2u�����x}��t'�;��z������?Xs��{P�C]�y�2�G���>A�;����~ ����%j���  �� ��p}#��"lg��B�(O"�\6|�c`�0.�Qݠ�X���L�� 8�-$H�f�xP�?��c��R "K�K�����|�@r.@���]�@D�D*�`�Ҁ��9U����XN/��x�m�H��.\�L	6�\*� (Ճ��wX�����B<zA?� � �g����
���}��=�-s�{?���<G�����H/�{@���������%�OI�{���B��<�|
�v��:=�>(~�>��}�N�=�m.~��
��xz��X8�<��2"�	�	TЁ��?h�H�QP
Gـ8>��-��������ˠ;��|Alw	�~��L�1�"�C������7'����wo�!����b�Or�ӂ����'�������,�����P�X��2�C�,y�gy�}>�!��h���Q	�����`>���顱�'>���3F��e�|�O� 3�z���TP�A�sg��}�bu�=$>���O7f��o��(���<�G�Og�����d(LC�m�XO���p�zH��AH���?�@�a�+�������)�23��