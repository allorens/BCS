BZh91AY&SY>����ߔpyc����߰����  aE��B}�  �S        �h5@ 4d� �   �              �   AH�E*�;�! ��`�p |�
G÷*}B�f��1��Xr;"�aFmvM�:p�f�;�]H)p�<�t  ��8 i����Ѡt ��}�����hG�  !  9(�wǻ�x��@�9��� 3��������:�: ;�� Q� r�
DL�����ρ��{ w8 ������ �d�ܓ��`WC����� ��4��� $�|{r�� :돰y{�4��:4u;���(` ���� 	�
ht��C] -�.�@�W��P�F�``�
 �_��F��@��N:�;`���;��n�L�8݃���r����Ӯ�w(�V�Clt;���c�M�u�t� � Q@���tx�� ��`�uA���4튣F[�'T6.Rې� 03����k#;�)��Y�ˇm����2���                 P�H   E4�G�T�U��M��10LM��!)*SQ���i�� 2h �����(�R�� �hd`h0 � JR�##&�h 4 �ST�4 �f�M)��M)�=CLM<��x�*���J�& #����` &z��e���F���s:=�|3|?o[ƿ��!!$ j��b[](?՟��`�0ެ��o��o�9���$�
��U���p����e:�7x��xmjҳ7�-�v�l	��?�sb�U��P�`w,�Ŭ�e�)�v�����t���v�yX�}�|	������ϧռ�O[���sǒW4濲x������DmqmWK�5��鮙�ac
&G}2�eJ�NȺt�q���\�F�Do�r����q�W���S��E�?���p�<C�Ft�՝5�d�2��Z����]9���ۻj5��ϸ眎�����s�Q�;�p��1����c~S/c�+?aM��GiF�XN�6�Y�Ue�+.a�z'ZVT��갧>�����ѝ Μ�NU���1YҶ����G��XO��F��;�:�l��yR7�Tr��O��55Z�������������}DMW�{(�1UTDu��<�9U�m��i���E4���:Ƒ�G���]m��DG~��}�'Ȉ�DrW��H�[q��}�j�:�Dou�G�k5��*W��b��ު#�����c���Er�#�J�O�#��ڒW�c�H��j#�'>���TDFuQڨ���Ͳ���+��y�m�Dv7���-J���FyQ�eu��R2�v����e��"73X��j#)���"�DF�Q�T��f��'+��j"8�kh��"5%b:ԭ)��Q���G%GYzU<�f�lBz����}ϛi_y�F�Q�vWO�UD�G�{��3��Ym5���'*8��#���u�]qagcѮӳXt��9������V��uG�C�mçGׅN�C�u��\���D��m��'k�4�|���)���#9G�}�U�gh��΢=����ч����xG��y<���q��8��r)�y�WQ�^q�]aǾ�E;�u*��<�5��ʤ�;�'���'���U��|w������%�b-V�M�Mw���㥷KN�:}*�N�>�����t�Ŏ�a�R`�H�*|���3�tql�Ʌ�Ҩ�4��Nk���g3�|� ��7�h���B�;'MS�M���3�E��65���`���Kx�w�x��G�I����WB��5շӣ��͖ݷ6]>�o�OKO�k}�7PfBE2�^��9ȉz:���EG<���yƜgMFX�ar)�Ǟv;�<�u��n�f3�F<��z+�m\q�Κ�:�~�oD������JR*7�r;{��{ԯ}���܊�Gr��L���Қ�3�a�5���v��2�y�Vr���0ң��c��^����n��c
�ʪ�S�N�w.a�7���G:�Q�"i��}�^c)��q��Ne�0�L�P�*��a�w�զa��cH�GM��#�먍��"�}�TG���=���r#��Dړ��9�}<��艦c?q�G�=�~��w��i�]N8�w�˿De�Dy��'��'T��m�Y�G0��Ǻ�2�R#��za0��(�������e_F5��#/qO<�Dq��ԌR����"9��8���"#1M)�DG2�Dy8����Dz4�uH���a�aO��#Do����Ȥo(��Qb6Ǒ�#̶�mO6�e��Tq�#���c������O���Q�u���G�6�4���=u+*�,��EDw�'�R�瑶�#���*s*i�n�v"{�6�9i�EF��;�R}߰�~�VT�i��ǑQW���Q�C9C�JO���o�j�=H�1�q�#<yNǛ���j��\W�7�:��F��1ʭ�����D��q�F���)��)�;�*7�:��k�"#c�3����a4���emߢ<��O��YCM"r���[D�S�S�s�#�{��֓+�1������v=�9�\�-e�y��yM�4����FQ��T��DEu��˸w��j#�EGL{��y?�Zq��L-m�Z=�8�5��EGoN5uܶ�"}>�jӈ�|Dcdr#�����u�oz��Fr��*:��5�DwHD��g���q꫈�y��D5B=q��h��"'[c
JR<�"&���"}�ⴤF���q�EFѨ�g����+�4�DsȌ'���R&j#�G��iH�#9De��2�>�6�(�""}V�Do��iH�������}�W�g(�9�Dq�Q�g�XG\���o�S*DV��"4�R��+��Q�0�y�6�H��'��m��Qr"&��3M�F�<멥#��x��Gޔ�ik���m�U")���uQ�G�Z�ꩴj�>����[�/#q����:�2�G�Ƕ˜�e��߰��k
j0��8G)�;�1���w�>B'+a��=�;�7�7�"7�sh�Q�{��g�uG4�#�qq����#�1M�Q�Xz����g�cޣM+�NDy���!Ϝr�L1��B�Cޯ�4�+��aI��ZDy���;�o�$R:�V2�(�y>�<��6�Ѷ��6�9s�����c�~��#S
�G0tݝ%�;�gvL8svC[%�j#c1!��=���Ҿ󴇩�i�y�5�j������(�a�1B�K�u�h�{��b|��}ǾۺR3�i�sH�NDN=�]�neM}��n��k˺Dwq�U�}�Tv#��׶�+e�2�e��q�Ӫ�q���7�h��>C��O#�����o�}֢9[�s�G��z����YTk�6�s7���#�qU�b&jv��UG��:�c���+jVѧ1ʇz��#�w0�S��Z�{x�6�YG��N��G��W��](�N3��cZ�l��L��Ύ7�w(�ͳ��8m��m�:[�:C�2�D2� 2�mtη�~�+m#�G�{U�cL�Y�Fv�za�TGX���*<����W[e�����JO���S���-=ULVT��a��<�Dq�D�<�Y���4��n��Uy�X�DDwu3Q�Yj"�Q�������l'Ҷ��j��)��'j���Q�DGj�&+�<�I���r�#�ch��"5��Z��0��Dk��e�T�'kjO�Q�Q����#ڨ�)��=�TDa5Xn#��y3^q���Dk��m�DF�Q�SR��Z��r�#����*��4�r�դa�VU��m�c蚪Ds��vV�O����G|�H���e�j��f��?u9\D�q�|th�3�g�A�gȰ|<����>��2�T�
�بF)�'�ck�Z1�b�#�m�TDO#�J��u=^i����+5L�G9�F"}��f8�����n���Wj�Ԫ��U�uWS�G�����b��W���:׫�J�uIڌ:�]q1Q盍9>�E5���S���$lͶl�i��^>��l�"1�GKgV>�>����Ɗ#{rC%>�܉���)�{�g�(��r t�(L>ؖ	��i��_�p��{Yw�!k�*D�?��!�F@��_�
��a��V���UP�O�����1aGH!��P���H�z�SeH,�$�f*�������<��d��g@����'�<@��
zR3�0vv2�����Y�[��I��۔�z�λt-%`�I/���v;��~��T�gD�v��/�9|`�n�����}��Dru�>F�w�4�[��<��˛4���[��,��+�X�As��u��g�n� #�Ott��M���O/��ޕ�խvt�����Y���9)��ӻ�6�ǍV�����w��h	�<�h��&8{M�ɏ,�a��"�5w��z<�.�qLp�[������u	��7��3�ͻ��]���yf�F�ai�*$�8��a���ǘ�y;$�7��_|�s}����v�\��9<q����xؖ_sn�G���H>��	�zn\o�T���Y���E�[ݣ�[`圅�g���t�_濈���	���U��ǐ��
|�r){��=7��a����k
�x����Z�}9����2O7ګ+�$F�0�Sk�;�������U\KR����f��yJl�~z��앷.����W��v�u�'��p8[LW�O��>���t���Tg�����ns���S��Y��:��b��NN����V#҄�������z^�#�ؗY[�y7���isu��0��K�fn|Ξ��|&Wݚ�(���DES`��ޘ�[*HV�OV�0MRq�Wg��H�6j�7�Y������s�-�O��e����B��o�Ӳp�7&b�{��L���.�3�Қ�����vg��$��-�x1
���������r9E�}�Ӕj�(�%BP�Y|z��6O��ۓ=��=q�8Ȫ�M0i�kP<H'���	o#	4V3nˈ@�AU�=��X-�+h.�fIwP�)�{�=��,��Y.΂�X�y� ��!�3
�êb���o#��������<�4�[Y�;�P�e��>SyOm��jY�e.� ��a+����r4�c�㵔$����F���za��ni��E��zo"�~��$��A�=��g,6�^���),�y�*��e�M۶؞��e��n"���nҫ�:�p�uǵ�W�Z�t0�Y�f���&�۹�Z���K��R��Y� ���Ή	3��<����O$����\ZB��ew�HX�8�bb�Z�b���O�֩��3�e&6��!�3�ꀠ�9;Q��|�m8���Q�Sd�RuD�������I3�����n���Ģ������=�Բ������V2������~?���[�p9�as�ꆔU�آ$%�u=�P)�л�o%��x��f�?%�V//�g;�բ!�bEK�W7ok�=�ta���<�����+�
���0��3�5�og����G�aoUUt�u��R�-�yY��f���/qy��A�n |�Y�r�����y�s�֠���O���Β�_�4�9#.1��L�k���wM&��u�M���z攖���n�Q;��|M��Cl8O"���PE3��[�Ė30��Y9�:y�=��	�:n �Wݛy��Bj���Y����I�(�ΟM��=�ÿJT��{~���Jc���2j�	�P̈yE���q�BzYg�ވ��2���|	iB��h�o[d�&Apfy�o���:!���FhB�ܫ.}�`��2���8�Y�fb�x�XM�r�?a�;����i�߻�Ͽot�u���?y<������b��˛�{5z�׈�K�?k��Ć�Hn�o=�ә�(�Q1t옣M~��ļf��N����v�?O_�R�{|����[�'����5�8R�C�;�W.ϰ�n��2�]�Or�\]�ل��1��if54s���%�2k��/m�˱wq������_�f�������?`�S�6�٦-f�L`��{��w؅�ғ���AT������?\��?|�3�1p���2o!��yu]�M�1��[19����/
��<X��zd��}�. �׸X�vi��/����9aJ��2ZE#޹��(G�Ar�%����+�inM?���2>�(a��x������|w���a*��
S�-i�2D��J�uܻY(C�P?t�����s*�oy�q7���s|w�[�8�l�ˡ�z��;V:�~X��c4˛�#z���1ŏP����~ǻ� V�"���Fg���@�!O��L.q�b��z\8p�Җ��-���7/{}�p��Λ6��x�:2ж�rt�An����_�f�ܑK���;�k�Y;�W��<l��'�1e�Xq5��0�lu�;���à��2���ձ~Ŀ2��<�������E�!�n�_�2�RAT���D�kl{�3��g�B$0�
D���ؠ��絭���'�)��q���ܤG�"�n�C̖�4����]����G��^J�+�4r�ضGQ�1�R�����tz_p�g�'�Ɗm��da[zn���l�g�֚�F幯30j���Y��H"�;�B1��߮��]͍����Q|0Kxa!6_C�M�͍NR)��9c�z2q�����s	驕AT��"n:$�&����T�Z�g ���v���gV��[0l[���N�6O����՟��(.��~h+K�+�:�՚��#4�Kأ�[�w�'	5�M��`kg�s��pM�hv\F���V`�"X���a1S�&YV85_�E[F6������mjc"�C���ǡ��tR�ffc�T�L�D(p��ջ��z9�D�3a��jfd��o�"c�5�Vc�О6N���3��O��?�?�#�G%�����Oci�:+
�l�"��v��Y[f�o]�W���:���
�����i������Y������d*�TwFn����L--Fl-"�fɌ�ѬF��� �2�1h�aP��J\~V|�A4�f�\�zN�c|쨒Ue3����6͹�a˯h.E+���qve|���C;����������?~�#?������f���f����
rk�m�C��2)>�6�r����j7�B	I��q幓�,W1�Gx�9�Z�cfi����t$�ffьD1���^W7�Z3	�d�K���a6+W�o�����M�����u��2��0۹G�i�<ؑ�Z?*�������]E)���c�Lͮ��Oݰ�m!��{ߛ���E���)�~�M���p�'����L�+ϰ����e4ǻ◔�z~��V�]
��YӁ_��9���z��O<pش8���bX�-������o���C������o��t�b��L�3��^�n�?c|1<'r6ү,I$�䗞�'y��~Ö�`�~��ta#�"
bN�S�3�y�JjE#��U�N��H~��+����o�KR�,ň/һ���*�<D�q��**Q8�����3�bj�
ӏ����@����%��˖�l��M%��kLSb솉61��nQ�0��O&��4�fS�տ�|x��ӮS��%����"��9����v.��hņl�|�ʰ��(�r����4��b����ٙ;)������}p�?��;�^�6\��_�t+_�y����(��#��.�}2ǘ]Ό�&�[	Sy�K����E��|g�|�B���X�pl\<��W�G��y��x��u����{��}�K��43\y�P�V�{f�^���v7�?�p�'�o�ܸ�w���;�<MoO�~��[���;�ܿ���WG�I��y����~`�?�&���3�?��v%��VNB�+�����$�e����</�C��OD�n]U@�;
�9{��زw�k�����uX��B-K|�י�!~�6J9�A�5�|��F-̾x}��^}�a�G}�E��7.&�XB"l����w���3���/O�.l䌇ۼ��j�A�gĐH��E�xc�=�xh6�-���H��OExӺ�+�r^��s���A�
31��_{������<���֣����b���s����w�l퀹W`0�"oL���Jy�y,�_)�8��{��W]cZ�Y��˄�� ?*�ȧ�9֚)Z��a��3P�ܚ8Zk�H7� *�wY�wr	I������"������XЇuj�C �ޗ1o����P�&�7#����o�M÷!t�~�i�	z����<$i-^c���9�Qg,ɨ��9\�<��	D�%�R|�ȓǫ�S�?1)��;�n�D���|��
FŘP����v�N�3Eµ�M%"m����|�;{�}'')�pe��ܾ��}G�����#d.��}���M�ME�ڥ�
(�F���6F���/dݴ���ϊ��gd�����QL��.@B�c��$b*}���~��aH�qP&m�c�����S��� �'�S���~�� Y-H[�2��*#pˉ��(�]�ӌ̊8~(����(�hz]�邍I V����Km���p�ݣ�r��yAt2�!�z@��Y�b�=��{��3���&Č?q�T�tvv��d��n�`�0�Y��V�j�h�T?�I�:�b��R�H6DM��w
DI���e��~��E~�<�l��	3!���<�p��b2A	ɗ��cNX�����3�y�>Ͷ׆ulj�[�4��fk\�]�ӳ@���4�,���a��6�\��[��U����$9*�-�e���t8�6���{G�܈���bl���O�&��8��A3�}�s׍��oG0 .DĪc���u+ۍ�k0���2V&�a,�&���	�}U��q�K$gМdƑ�ϰ�W@����#�ԭ?b8EaϚr$~X��Wz��;ޯ�̀��pnaV�R�?>|���X[c���5PmGu�	���2��!�{k�"hD�Dz{314�"��Q&!e�(���������m/�	D:ƍ��$���;LLM�fZ5�?�(��`��*�+��> ������a3D��i8��� �н1�{YhInO����.�P��Z���ow4���Kmд[]Ǚ+��v���>���,fCK����	�61�����@�6�Di���}�z�_i��k��k-��kv��V�(B3�K��T������}��v�)f+`��b��]3��8��b g�g>��1�9�
Gu��e�묫�˜4n#�˹GdF��8�k��O�@�d��?�O��W��h #����n�_������M���?��s�?�����ݿ��g����Z����u�|���5���9�(� �4 �z;�x6�X8��M E��x6�`�l E #@<���`�;�c��{ @���@z��\ֵ�j��.���YB��e)�Kn���4�TM��Ve
٨��8g ���mYY�
0��KY�gN9]u]A{羏`=��l`x�`�@p,Ӱ�����zh ��g��a�<4 ����T (ӱ�����,���`r��V���ֺ�������VڳV�LPD�LP�1TmT�el-m�jn��Ś�囍`�+Q�M��AM��͸�Q�jb���liHj{x���=�X��X�`��`=P4 (�����<P �hӰS�a�<��@<�����z�]�� �� POJ�I'$���X��+��*�R�mZ��Օ���ے�Z�f��e�+2��ըt�q2��W,��Ub�>5�Zֺ�k=��y� #@�4 � 
 �� ��!��@��`����� �������� �l���@���� � �Ps���V��k�k])��d���M�dZ��(ܙ-��Z�F��9"Hl܉ 6����JH���#jͺM��ۖM�9��S:�M�:�VogZ�,9�9crձ�k�N�n\�}���ۖ�[�-X�,����k{�`D����~����W�����l�=/R'�=�=�s���:����ʐ��Di�m�"#��#��"<������0�!�ee�e�qGQ�G��QG���yy��"#�""#O#�")�DF�����mF�q�!H�"8��<�0B"0���#��8�8�6�4�2�e�R0�iHB��E"4�GG�e��y�\u�!De��Dy�u�m��!�8�!��a_5�W7��t}���O�+!��w�F%�Yk��{n	�H�2X��b�R1�Z���0r����rahq�\�tS1�~#		r�`��2�c�S��S���A��ρ̓�1>e��Dx�UM|��?9���~1$�m��,#h#'����W�����}|f�OE��f;��z���t���2@�l��\�xЙ��@��˥���^�)�mЅ��+����oy�|�x�T�4,/1iU�7�a��%,)�["b�C��z�n�)5�J�	���q�\�~��!;F�1
K��%9�F���4&�����f7	i
練"��3}�+����I���uE���` h��g�����M����sWDJ���E�F�r5˔fW�0�[0`$��0�"��Lu�
�I�U�-����&?�Ul�q	c"����ĥłg�ڃ��G���B�f��(溜
k�TV��2d� W$�����	j���,��Z�s��c�ׄ�W�z�ݒ�Mr���8D..�+`���c-T�'�'/��aC+��JuBd�$�1!�ـ�X>�_� ���!1\��{��̙��]��u�U�WU��L��P.��+�����&zh(ww�W]uU��3�@@�����ꪕ�T�R��eE����<�:����>��=�
]E�h����]��'��w�pƔ����ZX2f�`f1t�n�m֌��ע����3�_���c�T����)�O�����h͋mw�{�����I$����qtP��Y!��a���~�d�D��N&�/�����A�)L8�p�KQP�2�0leC��PG��-�㥔�A����P_1��;�kcQk���[����{"Ѳ�"��1���U�9
�k�u��|^�z�G�4Dw`�2��OQ�;)���Z)!k��v��J�OKT�u&�RT�%�.H"B4��;�?}����@a�7û�ª�_83�
8Q��-�DyGFyN����]�5�uy$���f%��$�LN�'�"&�%�.#9�eo(Gl8���3�,�-��޶i5�>a�7H�6Ƿ]G�D���'�Yy��M)]a�j�UF��{m���4Qա��Qy4k��ۭ����$}����:�7�t���v�x1���_��fƓ)�^��f�E�]Z�Iu����oGj���u��tb�i�4����<�qG��Q��S�1%yRg3|�)�k��hվ��$�H;��D�?���h��`�
�3AB>�M2�٘Y�O�߈��`"�M������f��]l���XD����������R���z�CY���f���#��%R��a�Ѥ3�z�M5�p� �ڵ��(p�i��VogN�R&�f�M�:�m5T3�
��#M��	�a�aG�9��[~M`gN�,��P�_u�a�)���(Ө��yuy�:��RUo��f�54n6�l���'m�=�7���u{��d6{��u�,oo�	�Z!(�I��M[mX�E�����⬇15�Rgi�L��w)9�m��1�"jm��ν{]G:�!"�Ю�8�v���ǬM5�Q�jYF���p�R�[�5��1����7d[YV(4�t��Qkj�!�e ͖Q��iգ���<�:�<�{;��&���I�oO5�1���^�6�8)��u�l��k6��(�w�;�Jw��z�9+]����/ǽ��g�gq	ӥ�H�lN�'����p�I�[k�Q
�R*0��yjN��U9�����V���\�&(V�T��%k��BF�<Rb�� Y�-�%�.D��ʵs;���J͐ٯ!�W�Z^4a��J�fsp�B�j?|<�վheKd�������pO���?c<A>bm�AM}�j�B���P4Q�cZ����f�������8��A��2�kE�Ex~.�c7�Ǥ���h�
��	�wC�EC�J-���`�"O�
�6o�A��,�)1j��=j��#
F�m�ikG�p����Ы�WҴ�KQ$�Cm�H�e�ތYK��E�4>��[�vr�}��E�p���`�Q��8b�N�)X��F�Z�Uv�yC�֜��[�N�M���9�X����V��k杏"x��n7c�Q����ׯ|Ehl�p��5(o���IF��Bfŭk[j�a��/��+��@�V�U�uuNܵ��2-F�a��SM2��Ө�"#��:�)���n��ʦ��[���7�/�&�I$&R÷q&Ba'�<E:t��4x����f�Z��=��&&����x0�߫~��s�~���@�3��O����=��,=v�G,�aeUP�È���:�\z'N�Ûon�c{"�f���8��P��[C���#�ןvl>�U�r�mw	I�f��!x��Bn]�L�u9����֥4~C�1¢ c��x�0�a���T��%ŭ���4uh8@���y��y�"<�#���yF����S���m�c�ίZ8_�?HW�ɡ��<i�X5�Û�Ӛ6z1�������_Wi7��ߙN�7k��k:\ǭ��P(iE��2�sT{fS����l�e��w��R�6{��E.�����>��$�.,ɻ!f�4k��ҳg	,�f��6��-h::�m�����h�GS�G�I��Ϋ6O5�Q��1:���S�XSM2�/4�#���ӇM�883fNC��b��
��޲��/���2�y7F�a��\8�Q8ˤ�� YC���7�ڨ=�E��c����		`$���XD���e�M=s���L��ڀ؀�(eyaz32�L�X��I��?:Y��W#/,�A��-d$0Ht��6e��t7YYza2ߗt�	�=��}�Cx�T�XZ��7N�-��[Pl�e�FD3n�Ok��׍45���}��,3��
��o�^�&v��qr��	?�`���=6͚;�������\P�Ǻ04G5�	P�ș��R��D8X�-��fi��N=az�"ˡ��+eU?�%=��R���[)�L�p��Q�L�:Cf�Ѻ�(����f�6�l��3����2�3�2�.4���"<�#����#�q��H�Fӂ���Iǆ}���Ν8r��X>H�ƴR�ʫ��5������픘:|�!*�6��O�y��m����ȣ�.�X�(���m-���a��5v��ǈ��I��������ju���64��ejp����!?K3g������L�w��u��F���P�h�GJg�5q3
ٿ*(�(��E�Jl�Pg�(i�Al�^C65�0����?�������y�U�Ū�kaձj�E��Z��ٵ[,Z�lq�-O*�j��Z0��<M`�<Fx�g�����ݐ�5����xd�l���(��[Z�U����8�>�y^U�尊��-yl-QKTU���n1�ե��:��­V�elږ��U��n��J�}l1�2�-ZU����ŪԴb���?> |p����k���%����jFX�c�c��3�_�ձ��0�?���c+b�n1j��jZ�]W�8l�4=!g��a
<H;�!�QC��<D�����?���3Ƽ5�xd<E���5�d<SN�jږ�*4�TTW�y�U�-�b�Kb�l�j���ͫ�ajEZ�l-^W�ڲ�R��)f�F�דl�3�Ix<L� {�����[
�q��L���,p��8~��|p��}��x���B#��(�щjB��vW2��>d�f�������dx���)��ҩ���FC{�麍��k�'�����1�����Yߣ�;r+���n�Rj�v,�"���\�,��7��c��7�o�㹜��w����� ���3>><�fffL��������$ܒfx;��2�37��UuU$��L�`fL����{��U�RI�$��v�uww��7���<�m��y����yG�-y�:�ҧ���6k7��{v�kP�BHa������[p��L�Ҥ,6����6G!��R2�Ë�(j&�4� �����ɉa�1�-����c,҅p�@pf0��(�j�LP�2}��)���6�B#�^������<�D�R�8<��2j�5N��0��0�H��_^����ahc,ڇz��\��lih��E�5g��UՋl�p��GU%C�#8r�ֶ�x��4}G�M��t��e���10��l��2"6��+�u���/����5�%�����=h�e%��2�K�Q�c�5�@�8�=��H�cG�����Q�m)��[(�ַyםyǐ��a����X�+|�5�:�s��BHa�u��%�g5��;���o���2(�	�a��S�"g
P\��$ta��y����C������R�M:�nH�;P<2.�M֮��Z6�Q�Ѐ�� ���xߛtZG}�#����Clih`�D�,(����ba���k�����8_U ��Km�#3���ڐV�<C��A�F�:���A���u*X��:a�xg��C�L����4�Vt��,`��%?j�qA��> SF3M��K\1�Dn��0��ƀ��l��>"6u_c�>���Q�6�eF����DyGQ��-��k��L��'3�=�u�9���Gް��wd��,+�l(6������̕V���d���F �!�3 �H`ɏ2a�ɖG�)\ur���T��!�oE)!��&71+�R1w֖-gt�c���0�_�1X�VFW�勇0�D�Mܪ�R�ܕ$�4["�<3����83��5����܎N�|4�M�F���g%fKs�J40޴9B���i�b6Qk�Mty����A��k�$S:�裍F�1�>1�>4CC�rՆ81m5C>�ҍ"=ׅ+�}f�+
]�����Ѵ��0��w���־�t�d��c�ִ�&3�_2&C�-������n#�dL��r�:�i4���>�8h�j&pgѫC?��o�v�R(bLiq4a�v?��������P)WO�70}h(h?|Oˉ��Xұ�X����}��-z4��>�uE��|�1`l��0��i��DG��u<��y�v��3T4�e��5��Q�O��ĉ�v���ԭ���$$�� �C�-��cC��L��Ό��äy2���9��|RV0��J��`����ߣw ī�Q���"��h��0c0�l�{YHl�f���)��Ϊ\e�XR
s�?��>�4/3�:rOO���	xF1iZ�V�����UD�Ɠ<7���%c<΍P��L60�I�/�K��45���e�g�A@�<0�^M-T ϓ9�gU��B:0�oa|�VIW*��EJ�D��Ґ�t|TD�Pp�3qXRX31��)�-���La^+����X�hp��T;���3�kNT�a�*D<P��@i�LQ���cA�CG"�D�b3��6Z��4q4�pkm��]y�师�"#�����o��y��ˋ^�&���$�H%F�dKɘ2�YH6��p��9!G�e��ex�WG���q8m�ډ�J��]#a��n$gXD����|�ԑBEH�cٵ����d<R�6@�SpM46}�b��0�	�#�!������� O������5�F�4�b��Ъ�p� �#La�!4R4�k��F��͌=d8�5i�|�Q}PW�B9zm��������Ѩ`{O�i���aQ���f_��4b�p��M��I�Ki����͸Q�YI3(��tb��}��P���}���B�6�Hy	��D4�&�QG����08ч!
��*���MC5��B��0�J�P���(�줩�3Ҩ�h31��.0�g\S�l��?�o��"#Ȉ�ӁÃ6x��G��cys�Å��SOx�k��BHa�8��C�N�ѱڤ�����<�ۤ�M/�l��Pm�����`Pφ_�g�D�
:ű��61X�*���O�m/����l�;VU%[A¶+�lre�Z�������Imt�F6i��_&F��נ�a���u0���Do����4�&*oy#)4�S~�'��AL��(��Tl�Q���a�43�1��7��`��᠌6\���	C1qdA���H�C��J�xDxe4ٖϲJ��a���<�Sq.�����3G�� �64�0�0��AA���&���Uك;��d�ѭ$�B,il�u�>L�.D��*|1P��!8P�"a�h�)��}m��	D��lfQ⍞0����#Ȉ�<y�:�2̙�i���f�٧�z�	J�=�%��0;��n�*#�$�9�3($�Կ*\k<�؍Q�ũPU��E!�tւmN���5�t܉��A�������(~KL)�H2��������xp�{��hD�[@"�w���n���?'s��da�0������[a�-��R5|��F���>�A���[L�">�p�*D6l�-�;CpWx7AM,�{�����.�L;��:�i���Itb��16c#I�@������Ő4@�:��h���`�Z!�&Ǫ8�
|��ӪEe<S�̞I�X�Gu�G��SEx�3���!׊<�V1P�C����p�11F�8��)��&���1ha~���6��PA��F��·�}w�٤XÅ60�t�ݼ�<�U_{��t�s�觞��F����dm�Z$4���3.�����K �:����xi{-�zs���^M�i�d44�2�
�pfQ���7ӆ�3f�H���ӥQ,VUC!�����8B�V��P4lf�2���Ϳ?8��"#�����ܭO.n�x\�KT��r��%��G�i��o�͏���	!$$�����YۇaN�ʕw\��w����h<0�UG����*GV�y���(m0aDl��C�F2Z�f��s��m?�'"���0��d;����}XZ�!bȱ!�3M�g�kk�1-7�EigLV2���[�����T��trΔhacϟ6�0h�Wc�sf�Llz]�S�����Y>BF{��}��@��~���vm0�HН�c��^�,u@���C�x��D�0����3���D�!��b��ǯ�ͩc���S)( ��9M����)iw������E�J��4,�م(�6���"<���ǞS�z���f\��N�sp�H�0���m=yC0�?�����4-JE��D��{?��)���Dt`A���T��-|N���d�XYÅ+8p��ѦpavqPp�����x�Lgu
9A�����xRѽ%��G /-��x�-X=��n��}�m�Y�)?d\)||@���cMf��0���֋<�C�1�4AX���8a|G�i������ekC���0aw�������e�<�l��,��p�h(a^������竫��LN#���*"h��cԟUT���^� a|O:C�pmW��^Og�v�)�QjSm)��u�����"<���ǞS�W��{����V��S�޼��8� �Ba�)P�o�>��Q}Ҍ��ãl����6�g�}j1�Dց�����&+1KN�����a�ߜi���RcS�P&��8��0��u����8n"V�-Z��Qa*N�5c-VϷ�#Vt�2�)m��C
��yD�pc������pa��������n�SҜ+g%��{�;zO��GAm0�'��C�0�q{���B���[w��n+.+DQ)<1���i�����c�y��i��e:�|Jta����3_�b<m�Y��4��C?]���(m��e2�h��2�xg�_Eg�0�!����C�Rص[8�b�Ū�b�jE����[�ey�b�űb�V�U�х�È�ڙU��e,��]W�ae-JU���-L)juZR�c�-���ږ���������0��E4�+�-��F�Z��Z��E�居��ilR�V�2�-V����j��X©�jS+b�jڭV���Դb��W���un3�Z�U��Ҽ��­T�"���jZ�]Z3l1��YV��Z��-V��"��Kx�g��l�4|M�!��V?�G�(����G�/�B��1��c:6?cg�:5�����/���j�����x5��}.>��I����T[a�U*�j�X��j�صii��TU����u��ڲ�U*���Z�K������U��*}T��򿗛'w3c�M*[Ɂ�H�LP?�ɟ�9-{����7�/�^�L%ፗoΆ~:��5�^o����N�I����g���� ��t�A����O����V��#b�p���㽴�ҝ	�	?Y���U�F���Ņ*��UB̧(VA�j2A���U}'Yam�C�#�oQ��d[�RC:?T��a��SE7[Նֳ$R����"v�S���ey�34��4�5�!8j�R(Ĝ/cdV$��b�cO�� L5��J�7��3:*�q-E%��Ӆ�H�D��[bc$Z�_3�Pϣ��D[��?1�c_Q�
�[�ɱ�����?����e�Z�YC`�����ȠMda�k�oF*i��5�����M�(�b����6�PU	䖂[4���x�0#$���a�*��?�Ə�"G�a�M��Y����g�-[zG����̅�`�6 dI�C�MGL���5X��yC�L(�[���N��ML��n�zͣ7J^�]�,�X�l�a���ө$�T�e��s>:�h���
�45��������Ez���1~�:�9���>��}� p�}�}u��駿K
��6�v`�*�{]� rB��b���%�:��""&Iqw�n����t��c}��Kþ�����)�A��5
1�R6�d��2��d�_eN��3��#"YEd��(*�E�T]8t�t�2�u�F�z�>���J1C>�2�<m�n�!
QL0���uŊ͛���~�$u���}eA�%�8��	N*Y$'XaB���&<��A9����j�vI
�F5�sw��ﳽ��{��fr���u$�䙜�ᡜ���RI.I���˻�uRI'$̰�˻�WUWZ��Z�QO6�̼�k[�DyG�<#G�����_߷Fl�A���*�|joe���׮:9p�	j�+J)�D�Ũ��pI�(��h�ܹ�v<��(����cC3���狣W��l�B��ס�o��$a&��J�^���v�U�J��u�����t�lk�DG��J�4�})�hf�O�E����Q�f?|�clqO.�+��d.�k���E<0����-i<�Gc�����kd�x賍�Y�0�߾���|y�4E��ur���Ýn Ϊ(5�"� \nPlh���-7�-uco���WJT:p��[i�Z9ѵlgD� `���g;N�>��1G�L���w�PT~�{&�0�l�^"����o�~��G�E*�����߇���uC�g�ղ�d�>��ap�=�����V��#Q�������؊:i��m�Q�~m�n-�Du<�[�6�����,g;U�ꍴ7�,��Ǩ��(�@���9��ݿ?<QF}�>�(N�������Ҡ�0��:����X�����|`ta�dK:;�t��XJ�aŵ�7�+�
i�t��4���Ѽ6���tDA�ч�
�Lsn�f���[��o/�k^,�,�-D_�z���R7��A��@.~���#��Rl0���]��_I.L4"�1��Z������0䙌�е��ֆD�·�u�h�\( ��5h�*�ʼ�rQ����؃�
aD���uKa�;�x�80&�1}�GZr��/���G�g|�>ɗa��~eכZ�Z#Ȉ�<y�:�q����ӽ{������=Z��(��  @ ����>hpq=���6a���{�p0дP�4y���-R�`Ã-R;Kw�:��F�cY�����y5~�����h�e,
>>�( @�am%Ym%�]%�%v���ۗ�J�l	�K@��:n�����	ӁH�9.İa�>�T��J#~]=Le�ޚ��"���C,h�A��D�V�걏6���+��`�68���[_/������X��:0��t�o�ϋ]X`���T�@������s=�?��&v��Pז�g�`F���\�h�B}U�>�h�6��E�����C�M�883d�:���5.����q�q�aͼn�a���o���[^�j60ߠ5�wݯF�֎DUH40��ɓnS9yP�S�9e�zA�t�[�֝���%�7����|�Qlfx­uDY�c݆5�p�W����8|q�z�<�Ҹ��K/A�ᇓ
ê�=��-�������æ+a��@�#�1���r`��y�ٵ�l�D��]3^o^"�:8e���U����|3�H�-��0�e�UXR���y,"�x�V;n#EV��v7hΣ�F0�"���?q��O�cJ���E���n�82{}E�|�1�S�E2��H�-����yG�<�Q�W�;>�n*���gT��7�0JE�L-%�WrE�SW^�{�����D�k������~�Ϻ_��i��l�����G_Lݸ�hf��퉞�ɏOOx�jJ�!٩�Ȍ������g �#�fe��g�v��;���zW6�灦���'��DDDII�s=��%1�Ͻp޻����B��4�{ǋ)��g�{����� �kI��E�li:L�촋楖�C������1����$V�*1�'C������m\pnH� ݌�HfDi_�8Xha���j��G��8x�/�y��m�ٳH�a��-*��p�����L���Z�x6���<�>J��h�C������X�1�sz$�+Q��9J�F�Q�5�%�~�g����k����f��4�[�[�%�Nٰ�v?Y��E�m)s7��Z(a��"Qi|t�\��c=k�>�}M�=(43Ř�4��G��yG�<�[A� ���}����/��G������c�$�{��k��w�&}��$a!��E�I�h����E"�5ָ�3F���Jލ,��i�E��S�la>kL*��x�-tS�ʹώ��pa�Ү#Gu��g�H�6��ҐƱl�;�0�~�h֥/��h�f�v��A�u	4��qi��{��ژ��
��5�͗�^��Ռ�"Z�J>��V��u�	Z% [D��|B�;��2���'��9!{�Vo�����Qщ��k],^:].S��heC�fĥ7�7�0a��:t���ќ=4y����2�ѤY}L	�gHaA������.�|ꥩEZCdR���qe�>��i�i����֏"#�������x��A�컽�\��=��8�0:��ҍ���j���xs1����z���#�)jԣ��$aD�^�a��l���Oq�~�X\���E�_��0��/��g�A��C'�	�60�<���R�x6�q�$��6�!�%~,�|�x�`ǘ���}�]�鸞l����1^���V�H���2T�h�گ��V�0��5Q�4Zp��_`�aی�������s�����F�Yf��l����f�'��n��2����^��(�u���[���9},�. ����L�v�|2!�W5􍶱��
����� R��{�R�Z�	��񥴍??6��-h�":�yN��>�4zo���9�}�Ҋ(�� !�a���{P�!�p��)ʧ�E-Ui6�k=g�w|��5�5>����[��fg
�3XC�X>(��Q���:ah���4K{#�T��H���?>��ܮ���$�Q&-�e�-��6��CKepцȢ6�����M�t����mO��.!��B��[6M�jM�5�ʆ�M��c{��^Ɨ��~�D���.�QmE��m��7�I�xi��Fq&��n��5�>�)��TU�HS�:0���Ԩ���eRG�"!��4P�K
(mm�����	��3�"�T��C�V3C<�
[l�Egu�}D�
��EC�%������~i�i嶏�-h�":�h@
5��2[�:��)�\@�P�N����	m_d��Yc��Jx���R��f9�"	-;Z0�)����T"��߿���D�p=(��%1�EM*X�B�m�邥6+u�|��Fg����N/ǤR\]��^�����(�G�C��8�C
K�7η`|0��$�l>9c|c�g��0c�Ĭj�F��Hq_T3� �æ���zSt�T:,1�(��<Dq��!������oJ��Δ�Z��u7뻗[70���T��EP�Q��������gF|:Ce!�C���3�
hz��Ά�{�g�0kZ-k��40��Tlm�a�#�џa0<�6��xa�>wEUU�e�ΰ��xXD���լӼ��Ʉ�hlc0c�FaçJZ0�f���ʡ֝O������0�����&,83��,�fό<|h���Du<�g�b����+�*��!�Ba ��'�}���x����8� ňg��7�������8d$	f�(�~8iV���������*Qü�=������]8�p��2��w��W��}���Ϝ�پ����T(�#k���,�j<q�X]�t���O�^��`�4�����h�)��}FoZ/Q>>m��;���pz���b)gHl�1��¹��ݚ��mp���7������}�q�_���?��<�͠�4
*	����6��(Anƛ�*�,��!�&�lp�ZgƈgV�KC�6���?��9%bҢ��۲��n���F+H�=� �C	���������cxV'��6W�t��h��?�-�Ā�w�C(e��A�E85���,�<@��0�����p~<aj�qV�mV�y�U�-�p�R�ŶŴ�mV���*�l"�V�!���M����i����i����jR����Z�ⴥ���[Sj�}���-]R��Z����)�E}h�х����-�R�aŪ-��u[U��j����n1j�Z�E[�0�[�e�+�i�U�j�Z�����S�"��߉��4CF���zˍ�?������U�ԵylYQV�U�ūKcKbԷVͪ**Ե��Y��C�	m����(�(t?O|PS��Q�d ��L���φ��|8?��k���k�c-_eh��jeQ�Tc�صEDc�-�ͱ�~U-�[[U��b�i��TU��l��U��mYU�j�<�m��m��6?o}v���#Pl��&8dQ?o�i�й~��N1�U6B�tu�	��I �>�{�E�f�FEm���Ȓd��b�n�[h�F֙��������q��B�c
|}}��YE��������u�r矇��/Ϗ�aP+.bt�h�$���C�һ�ڨ"�qe�H��kM	�ƃMca�26�S����!\����QEo��z���1�Nt��u�~2��&k�y��k_
V[���n��﻿={��.��g^�<%~{��$�W���Vr�[���m�=���	��'�uZ���>9���a�<4/.�.�I$䙖��y˼�$��fX,���˩$��fX,�w�^G���S�<��<�k[�Z<���ǞS�1�c?����e���[�Z�ϛ�q�$DQ��~�x�Z��e*�a\S��N�u���"4|@�C��ݣ�EkP>M[�ᎺNڶ6k��}up�*[�,�|ۺ'"��C�Q�k{!�������E�z���+.^�VDVK�5����Hԣ3��4�_l��C�\{�.D��aA�w5F�Ѣ��~Cf#M���
�k�4=��H~6���*+�a��E�=xغ�7%�vFq��3�{4a���z}U(u��US��S�P�ꣃ����#{�7�4ѓ
�7h��ƅ�0m+���)Q�T���|=-�-�*�a�͖3�E��?-ſ8��Ȉ�<y�:ϊo�޷�����PI�I|"��T�#챹F�E[!���w���4z�<5�6�QCH��k��p�.!��D;�B!���E�+g�����'�Ok���w��KzG��eX�����g�]���/)�KM�3���ϐ���+Qp�ٺ.֙CF�g4���wm�V���HB,���M��vx���-,X�iĸ1���l��!!��sTgˬ`ȋ�ҋ�WL��� kH���W��O��(83ɫF�P�Xa�����I#SO�ɇF>�ݬ��GI.��݇F���M�X��4IE��!kG,�A���!ǎM���Ȋ������!�et���-�ŭo"#����c�:��_�&�!����Ē�I�	I�k��I�-x�*�$���
N�H,Ʃ
`��d"�!6�l��
�2�~��eJ�
RU�Z�LPX:����焘2���������
�CDGl�RX�]�lgI��v{wf��?߫��yq���Pt1ܪ��.;�UVl�p����e�th��}��+���`�bcu�p�G�P�yi��9�F2�EFݓ��,���6֓>6y�/L�`tc[������S�F2.�P�P�(qH�aw�gKZ,!�dF)�~0��"��Ӆ�m�X�4t����2ה�_Ytڇtn�c�᭪�44|x�6>=t�ќU�T
�����C�"��g
���iÉ��-��Ϯgo3�FA#�M����0SH?	߀��"�q�����D꣑��P��Xh�<v��k#l�<1��H�CMH
��l������ַ���<y�:�+�\�%+�Ȯ�V����6�I��X��a[ ��hll�ۀ]�G��M]�J�]�m�b1�5׍o2PU�,h
��d���bk��q@~����G�ĩTG�f���!$$��f���-h�]}��B�[�ƏG2�*�{5/��o���|f�"�|t����5cj%�^�3T64� i�ƶxg�a�J/��!'�'�<jAE��$L��u�F��������`���2�ū���"��[i-�m�r�(2��[al�lD����>.�E��e�*��˒�ZgU�B S�a�k���'�J������؁{�N����G�(Ӌe�m"�MvJ45�Δ�\�Zl�2A�G�4�3^!u�* ��D{���X�(������4�0ʈ�������*�1�YwL�L2�-.�lF���iZ��f���c咒7��,���|�����3��-�-2���R\�2�k)�����08��][VB���������l01���9�J������>0�	�;�Ɗ�a�O����̼�8����Z֋G���47������`w"�L�{��	!$$��+O�E���65�D!FA00��ܤC:v�F�HP҇9ܣ师3C�3DF�2�(��:����8},���[eif!�!c0�4�+ڣCC�l��1��o�����?��'�%�wg����H@�[V��i��"M�����m�1�,��E��E�Lf���z�o�uM��k�2�?�ύ%���y��4C
-�h��B�ҪM��Z>��!�����){3*���s�h���C�^,�;����8aH����>k�ED1�����R�S0�εG�,g:�h��3�7�3!�G��}�����#Key�庵���M�883c�7U���Hc�k!$$��d�q>kc8^�6P1���V@cW�"V4�Q�=���+�D`��""���������m�B١�v�a
��3lm����;Q��!�g�:�F�FX��(�c��F�r&|��3�R]�F�l��cF�񓔜��Z�~�3���W��g�Ϛ�g'�r�8W�a\1_|�����&lv�67�Ə3�s�UP�eU�F4#Q4|0��p�>�C�祤kƆZ��/j\h�.��b�X�5��A��g����Z2����R�4iD������a��T@hh�|��0��Š��!�Zq�_�q��խh�����4tkE�� DX1�#���G��צ��&7}�쨘�@���տ��Aeޖ�5��'����L�O�	0�P$NP�a-ȠN9�]@�-��A�Z����O����me[*�n���b�X�#	{y�|HSh{8^�ّ�+�70�l����)+(���%���B*��H�&�o��LD� �4�ͦ�d�i�1��|#���q��[m��7�{
��4Y�14����j�P�2�Z���y4�d8aGK[>}׫�GUt�Ĭaᝌ�U-�K��L���C8||����h�.�0k�n����/Q�VS��W���F�/��*��J(�E��bc=���H�m�jo�3��M͒�H�g��_t���:�_0�â�(3��
I�r7�6�b�o���e��eoθ���ִZ��x���V��G�H�fl>C=͟�a��c�}�wh�����H$�K��	|��4�4h�h�W����6݀�|Q��쑖Yh�K�q%Y�#�6�V&�=��2JnT�m��T� ����o�-Ҡ�8+9xч��GH1ș:Phg�Q�}͒�h�F�t�pg�����~��������X�s'�� >�������k��>:5hc�_���c�y�;Z�!��q���r�V^�m��g���6�4E���a�F��>(Z@ѿv�F5�%d-鑕R�mt���*�ph�����-�R�F�QveP�:�j�����}k�n���0ʜiƑ�����ִZ��x��w�o������Z_�H~c�2�J���y��	!$$���K�8��F��2�׎���9�^��>�GJ��A���[�꩙>6p�5�oo���I��6��������)��z{��#h�) Η��ꬼy�Wq�u#o�R�E	�!?�?oxO�Ќ:y@�Μ")yDv�y(��2BH�-��;�Ɠ����GFϷ
�b�"�`�C>��z���s����t���hg#�I��O�USxbٿ������fҫF%�Ŗ6�v�Z4�u�h�T�63�m<������kE�t�q�Ԯ�Һ����}�	!$$��-H����
��5@�p�E4|>���>��#q��1��TF&���Q3XEl��6��	?`~r��PYP��n���kI�!Ӌw�4�Tp�"�3t7��x1�2k� ���7gÈ���8��6iE�2��a��L9�d�+o_l��q�s��ۓ�
����F�9�Mό4xpaє��8�S��י�E7'W/`����E����,ሳ�(g�E����="��6E�����u���cc(�&86:���,�<C��χ�,�6Y	����W����v�y�^+�ilR�V��-�:�U��cj�E��Z���*��mqy�I�O"�U��O%/%;1��jZ����Z�W��Sj�-�>�-]U�ձ��jyV�TRч��֌Z����<�R*ԋbыF:�WbʷXZ�j�Un-���W��-T�Vl�j���Z����j[�Z�H�N-��\U���ȴ?&ǃلPg��+ó���U��-�U*-��b�U�U�Kb�ǖ�6��jZ�����an)��g�x�x�3â�Q�/tx�^I<�I��Ry)<�䥫J�aKSj�}jˬZ�i���2���S�<?��||N��c���	�����O��?0���\W�+*��R�Z�_Z�g����v+r꤅]Q�ߛ	,_ھ3EMI#%���";(��0L*:��"MQL�Sl/�#�*<�d�����l���{-� %i��	Y���6�iP���1Ä@eQ�0�Q� p�n,tD��ϨE�Wވ<�z�I6���O<&�kA��'u��pK�}�n�i$�,�>��-+rV�-d�D6DeT�B��g��O,�b��N����N��$�,HP�K1Au�A&���T�s0�I	K�O8�hb:��F}���o�����D3鈘ݱO���Knq+WH�8���:ؚS��Ļ �MWXdBM��*U'暕���d���S
|�eV4�u6�0�.�lb��R�Zvl=���uգ�p�Y����������B"����,�*J����j�Q� ��D�f:�d8�6IIT�j`��bQb�����f��-�λ},��LRX�q��ޝK�*��b ��O���2'��r���%��8Q��A�b�E���%f�z��?��0p~��4v/3��lo�tі���[?'�iI�`{�β�������>�E�Z�$��8�W�g?�`��:<V�͞�ē�ҭK��M3�w��f�z�8�����s[��́w�_Z���>��P�Y:�������ͺV������d
Of��q����3�ͯ�+�SX�k��nݸr�V��Nńf �#B_��ੰ���h�,��1N&?�������||X,�yw��I'�3`�pv]��nI$�L͂����9y�$�y36�k�����U*V�i�i�qkukZ-kuӮ��F��RMc��J)"��%�\h�k�����Yڝ���2ҮJ�Rʴ��Y� �pJ����1'�E�s����R�Ɏ`�]w�{/[k��oJ�S��+��0���k�yZ�m�7AWQ\-ۧa$X��G�;�rG(�5��M�E#��R+~�ӻ���8mX�C6v�F!�5�4R�qf&�h�Cem���89�K�"�l�J�C4�+����4�Zca���$����c3ayK���4t�dM����0G�Qj���{���͎L��#}<a���H��:�N���Z�@��\B��dDѓ X�_2���ήƈ$2��s�ţE��0�85��7�UJ5wl��;��J��[g��Z[N�����խh���N��c��w���9���}ʄ��DA�d����<\������i%k㸟�ڡ��m���]��8�K8��f�h��Dg}�K4}T�GM��9�J��������c�aE���"�`�Pf�6�>��7׏�ڭ����ڒ��饪[CE��*(��Xώ?3o�Qet�X����5��6�$rv5F��<!�ъ���lf��[���q<��,s����<���!�y��<�yx��2�9��!J*������Z$�8Ξ��?qRJ[��q�e_#�?|�����g�T�#N��m���V��ַ]:���9E)[Ü��+�,�+Uy\*Cf��P>��c��vF���o\7}��$���"�{1ZZ4�h�֑
�1tû0fI���4t�~1pfg��8B���ȉrc�45���?/cp�:�j�R���󓰇�Ą�O�JJ_J,erޝ�ՏsB��@���y>sK�R�ϟ	>�ai�hڱ�p����
8�DQ:�

�ED�ZÁ����KU�ĺ2���a�d|L�=�h�"P42α��Lh��mѴ5�||��^�9H�����^�x��Q��Ki斍��ukZ-c�Ѡh�F܃:~׃�c��ݧ�{��	!$$��<h��--#F3���Q�}-\:Phe��p4��QC_V�mi|Z�o�v�}M���Bˬ��9P��["�~h��Iχ����MV���V�C�e��������<3
k[���F؛f�hZg-�k �ьу��כ�a����uQ�7"�p��oû�(q���mO0���4R"�2v��Uuz#k�6VȢ��cc�m0c+���t�y���w�<4���Vt�߆�Z�Z*��n�9���NN/�����/!�=����4��tѣX;!�b�!���N��-m�պ�����l����6TmʩQT��}-�\q���J�޽��R��-�GB��:�˭q���mU�7,]-�{����'�	&r���̏3�f��k�vv�:���cR.���^�T/E�bm7-�?X�V+���O>#qNWj9.�Qt�mҌ��Q��&&��n��6��"��%J�8z�������þ6Rf���;���f��z8�R��{�������g�c�5�v�$nփ�,���Q�\8A�_��`1�-&�[����-@���ہ�7��[,�\����{}U<��uNZ�;U]�Yj��,,�L��m�l�1�p��>[�㍸�F�0c64H�r6ۆ�F��3�:�4�Ϳ:�V��ַ]:���oUN���$$��f�P�7�h����z(�E���j�Yc1-yB�c;3G�i_M��F�;/O7�N��~��gM��<��Kg{c~8b��>6�G�|�*g�}t��� �-����͖3Zl4��F�g����|�\;
�.z�/nn��;tt���Ac%�t�C�n��79$$|�|8�:|�2������Y�p���4p ɯOwvM��_��o}w�V�WMVws�C����e��S'��G'�#FS�F��iO�6�4��h��Z�k<l�l��c\�e6����m:~tƉ�E�n�����y2��O�}N���b�X�#	����N�vQծ#���dj4�<<���"��Vx�P`�1{(�G��m?CzmA��xg��R40"���P��g�țEQi��J���v[)�#eY�}�o�p⵰�����4y��
\\o�����C9�z)]5���:.��%�HUJ�Yh[��3^O�XJ�)Y���|��$Pc���GM�z�k<�᳋�t�SP�񠡗^JDl��,�ag,�g��"���ִZ��N����o��%d�W�V����!$$��gN���~�G��i]�}�ܭ~�:e�eO�T�ku?~uZiz��ﴷ~pʗ���)�{0��icEH��&�ј�I����*""0�;}�hg�kj�E��������h�+ŭ�3��J��1.�/�	���eH�B�	u�w�-��Utʊ�����mJ�>�Z��ǂ�A�����|b,�g�����A�٢��a��k�7�߶t��K��}ǐ��gl�[��k{��|���u<����C4aFl��έkE�t�q\{�j��5�r�������w���a��H�my^Q�q��+|RJA3׍�D3�i��.m�: �_�u���T�V�2�����"�	�M��K��8���EG豟�0zt�����q5�㫡*�G��X�W���&;|S�Y�Ŗ-2��hѶvpў�����)|l �3gk]4��܄U\m�8l�G�#c<a
��Z]0�n���QEb�_����3�zuh(f[�ۥi���m�b�\���xfkV�5�h�g��;�/3>�E�h܌��q���p�Y���7�}�W�z��yp�����ݽ��ۃ(���ݴ�C.lqo	!��5�+��M�lLg~��E�W���ܗ-��[^^K��Y�-�KDun����u�T�C��z/�{���~��?��BHI3�F?�~:p(c�m�f�Q��g/݇��1�2-��Vf^��Z7`��m�.g=�
�c4�����}ru�q�{.i`3�:3��{43]0Ԛ|7ㄓ�C��_�~STu'����L�^AԽ]��F�ٵ�6E�x�d43ѳ�Ϗ�����N��]�t�+�kґ��ɉ��FA�1y5G�6��Ϲ�J�E�M#�>5�kaG
0�N�î4�/4���el��"#(���:���"#�G�GF�a
B�!#����#(�#h�#��:���yG��yG�G�q�<�u�QDGZB)DeE"#��#͢6��ͣn��JB6��"#����E#���H�!�y�ѤmL�2�2�2�"��!�<C*De�"8�#̴���O<��yky���-h�ֵ���ִumi�!Bt>)s�so�}��3۾��h6����_�Q~)����>^���yT#H��V��׹\e�d���XטM�6s�3UX�#H~+�1�G��[T_"	�!ۄvc$ء-!Fc�so�M��-J�ܮ��R��X�&i^��q򩥧ڇJ�rNx�9oF�|t�7�.9������9������5rB�{{(��a7}�9^�4VyOI���z�*��O}��3�`p,6����I$�Ĺ������I'�3`p,6����I$����x6�kV����u��iխպ�ִx��f͌��
��>wz�7��z�S�w����}�*BHI;
G{V�(�Y��cl��1�G�0�Yh�f�).�422�s�[G|�h�Dl:`A��՗�U��z��"��?��AD�����M�~�~,r!��)G���8gU
�(�P�gWW[o<x�c���5�}�i>A��czﾭm`�ƈ����:��><R׬�Ef�Ֆag�|f��>/�ޱӎ���GEh��:~��o}OmL��2��<�u��V��֎��a�uwZ�5X�:�]jBHI��m��3F揾ٱ�̭G(��]m�3��C ��i���?��!�/#&:���xgՏ��p��3��Jڵ��ԏeb�3�1���P��C�}���4+/3��dj��)k�R��G�eoO���r��E��{��T^�!�4��e5ݞ�/����U_��|t���,#)Y�i�E�����a�O)�u��i�[�uխh�����Xq�5W�g=޳��:|�V��2YB��j�Ք���׷��z�]��&��T\��\�lJ!cs����i{m{*���:�n9���$/͉astg�>�W���f�p���3Vc%�*:ی�IeR`(�o�+���zW��
�-����hv������Q������Ӆ�[3�{��zf�K��z�k[��������������.��1p�Py��O,V\�w.Jjhe��13�0�%�^L�Z=���*��%e��G����k�έ�k�γ�ƃG���i�K�"y�kE��S��A��!��z����s��s[d�;{Y��yu�퀗������mCg��*E[] X�z��6F�߹T�h�Xh���2�x�M��?-��]Z֋Z:�u���C�!��^Ԅ��DC�ZV�,��x��fc|7>�_d�F�8���C_/w�W86Y�ٗ��KR�Û6a�>�+rN��}�C���]a�N�!��Fn�KHK��
4�T]�X�P;#�)]��l�	�ZZ�,0⭍������fѴt*���l�E���w���_}��aEӋ�#&S��*���//��CtÁ�A�t߲�$e2�l�a��]5]�ww\42+;��B����=�S������������>a����[F���kE�u�!�T�26�c�h)�QN]1��1������	4xFu����N��a$$����QH�{��h0����	��]Z!F���UUWn��ܟ��g�ݽ��A��ndІ���sn�p(g��:�p����L��uW�<�l�>ۘ|^��Ω�F�Vk5RU�VM��N��5ׂ�-�N��e����[P���{Vnm���4�q����U.G��7����n�v1�Ӆ�(0��e'ަ���eq���ͻ!�ݸ��L�ehn�����q`]k��}��-��{�$��0fυqQX��&W�A�C6C�uƝE���Z�kG]uN���[�rj��U�ִ���HI	"!�(�Ͱ���N5ËH�ͣ�!�4�1Y�텪�ySꍌz�FBK�
��BU6FXʫ[~o�����C��g�ֹ������7@�_�z������<(xᮔOf&��<m�|a�w},6|z,�&�������3�פ��,C��q�-�h�s��Ţ��6��^�ےp���u[8b6E����:G--��A���̸�N�:�Z֋Z:��|�Fb'�nrH��\:�}t�e�f��l�r�� Mu�:��[��Z�v�b�&$sҐ�؛~����:�����"�Z�:8Գp�Ml��h����=d_D�Xe��+]��k��L�l����+��3w��g�e�k�BBXM�#I"q~�>�{�qR��zǆF�#g�\n1�Ά�z[�9��ת��O�f[���]6N�A�������?�q\5�5��%<\8���C3g̴4R�S|��i�-���5[Qhl�,s����u$r����1^�9�F��O6��ÇƼ�˳��:�&��(t�e̷uƱ���7��
H��ぅf����pڋ���#�h�>�S��.��Q��r�X�y�(gl�Gx���񵼵�֏<�a�������1�d�7	!$$��n۞\0�ےQ������<�X�G��o�6�Z<��;[ݳ�"�a�1�6ڔ|�å\=�o��R�ycn�P΢�ģqm���F����YVǨ�l�Y�5�}T�uT�.�P 2�,�F�4��C��C?��۾2�)�iB�̠��q��Q�f���
;�sEt��4�z�0�C&:����8����
�=��dw!(�M�mY:h��ZS�4�/8��?:�V�֋Z<���~�R��qi�
�R9��'����A|�LW��v�$$���Q�7,��~����,�Z������C���f��>G�zZ3F�>>��e����ki����r��?˂�w5��{���3�:w�!!��OP�Kлo��N�5\�1���#**�b�&̊�v�!��ê���L8C^Tt�l�C��c,��qB�����<�%F�TQ�V�x���C�>�Hw����Jg�z�G*�Ʒѝ3�+�<��7U]��)n�M3�>ɥ6ϭ�d�j�3]�!UWчtj
��t��Y��l~7�`QЅ�(�<�ο:���Z��S�8��<u�9y=����DB*(�K|����TUGTTc�^:�3�#G��,��(�������#�aY��$��3,ȃ(U5]oeiB��T���%�qB��Ed�*
F�x�Ç���>$��Rf��ڊM\��ײ9��EgA�[&��||x��g^9EW�T76�3h��uZ4�3a�#W�o�#f�ce
��0�-#5f����3�h�e0�_%I�\�kL�3V:'�\nL�x|yQ�<|X%> 3l��<Yf�8a�g�el��"#(���:���"#��"":�<�8���B�����4��H��8�#��<�Q�G��uG�um�E!F�DGQe�Di�FȈ�Ȉ�h�#(�4ˈiHF�DDu�P��Di�R8��"4�8�#JF�e�eR4�!C�!H����GDy��u�]u�G���YkRֶ���#ȵ�o8���,,����t:���)�o
���*+%L�dĩj0(�C>�T�#+20�D?�c*`B)N>s.Ʋ�A�(e�n1���`Ag�R7>����>�s��ƃ���
"�"c%��l���IV�/�!����W@�H�����Y$R6�O�H�_2H*� icb�~(�p��АʰJۅu�H�:BEŋx�_�`D�mط4k��oz(���Owu}���
m�K���Ad���(�;D�c�D��
DqJ��-�V~�Z�i`��a�j1PU�򞻡B��첦m3"J�	ݏi)�(-j׆Ӟn�qRw`�����ճas@ߊ"5]�C0n�4��g��	(�t���}$��[s*���jf�q�Jo:.6�̰�	%�,A�[�~x�nc�Y6B0���[�4
�exIDHD^ט�0�a��Fo�0��cj?�q]��_���<z���]�ۣB��I�������",����y���})�0�5:���Z.BR�2�X/��4P��)�v�n"��P�b,�}tb����y�$&LΫ������s;�Ǯ2���=�nIʟ�u8=��$b���y)XŽ>����;�A���3g��&՘HL�F���1�I¯��j�%� �E7��V""_q�J$Z8�m]��;����t�
N�N��J�]n��4����fY��f-İ>̷5�G�E,�SJ�YN��E�ݭ���	t`뉮�֚��F��3}�&�(�݉1u(���sq�hlZK�mt�wl�!��O~;{��z��x6���ԒI'����lww��$�Os;��.��3RI$�3@<���U�T��ˬ�����[�Z-h��A�^���#:?ؙN� �c��v�����ƛiو��F�!��C�[��H�2Y��B��Ʊ�p�0ڦ�q��+�v��t�4f����r�9�_��������X�W��'�S�HYW(nԒ�$#m�f��G�퍷A����-V=�6��UY�� 3�n9�u�Q��P�Ƌ��[4�wʕ��\9ÿp�g����o�r���~'���J7��3��c�������57�S��ÁTt�SX�FqR�e��5�8��%�q����>��T3��i�Pf\Q^yێ뼼�eN�Wv�!����N��t�Ͷkd���o�|o�㠊7�e>��i�e���c�T���4�a��Q����Z�ukE�y�:ËҘ�v; �]�HI	"!g&���]�!eY��~TY��ؾ��<D]�	��w;T�����v�h��Z�^[[�㍲�?�sa�����m�%{g��%�p��0���i�l��6Z�xl��Q�\t����hi�TaC
;��w쿴��C/NفѸ�֐����2�s�|�.�p���>9��-*4Y�)c`�5�u�A��������ti�ˆ�Q]o67M��#Fpс���Yju����㨎�-�V�Z������~��XƛM�&8ۨI��oG�p�BH�5�j��^�N����:|����n�������t������T]���nBl�af����,���=�~Z8hxom�q}��A���1���f9���Em|2��ޖQ�~�0 W�l�N�ȿ��������Q�lvg6F�q3n6�4txxZ9g�e�h�g��z4MY�����{!M9)�8q�ǁ�3�L��:��q��g�W4�QJ��:6s�a��cp�C�oN��B߱|t�N2�Xm�\e���ukyŭ��g���jD��%Dm�6;��m�i�^�g�BHI	"!�����v��R,:t��~}�Wl�@϶���>yqO�#���aG.]&��v�1�n�#���FBZL�~�a`���>�(B�WA�:a�O�6T���G)��O@Ϗ��&�4�$ulgK>�G%��dvJ��62.w����W�f:=Y��͏k��kkЯY�?Et��W��<FiT�m줪�>c��q�<5�h겑�ѣ/��m��aM0�̭�]y�խ庴Z�מS�8�ô�q�x���٣H��]���R�r�׽�tf\V�W��t��{H�YY-���ރ��;sXӭ�G�"T*S��Q�ʛ4��8Fؚ�EnX�^S�RY�\�Sm�{I�I|�V�HK���УD1#�ܐ������<�CEp���γE�7�l�z�g�N��o �T85����~d�����
e�XY3�����m6qY��3�w�fsհ����ՠc�}ly<2�`R�Υ�P�(g
4t�T^��<��n��T���������%�p6y|lc�S/A��V�����U���]|sэ��٘�1[+.�:c�ʍ���ccL��Fn���i��b����,��,&����X�5�eL���FV������Z-c�GhC�n`��_!�c�����DC���#J���g>�κ�M�.��m��pᠣ�}5��Ƣ�#zi�6=:g[��N�cHo���\4x(��-a���I���c��
�9�86�#]lv��nD�`n�����:�h1�J�?��?�5#�]��]D���A�{����t�\E"�4f�>:�Q�k�hڳj�����R>�D}>�}7���C1���ρ��n�T��F[8s|�t>��S�:�ˌ�:�����[�E���GhCe��-�����[W�I	!$D8�l��W[o���h�dL��D�ۣ�4a[��J��K���6��_zU�k�&ݬ��#������x��u!$#l���"�nDI-c�D�?}�hdg�2��a�9�q�a�aӫ���(82�g���hN	I������	(�� !Nh���,��6J����gU��AVX�_��0G8m�kE6@>>����ʀ&Ƶ�j�6�~��;�@��viu�)ek���͏6�,MR5-�Jr٣쓨`/�1d]�"���A�Bo����aε���Q��a����l�/�Z�g�ǎr�"�b�)��x��8_m�6�(��a��^e�y��張��Z:�Пc=4���~dD�2��y�ل��q5H)Y�wۢi9r;�p06�F	�-��[�E8�ȔaM9-�1Pj�aY l����;am+i%ul#�l5U���m���!���7	!$$���=��Gcc�##�ʦe�҄��	S���p4p�3Ƶ���CT�ʃ-d����֮q,A�ER�qT��΍�����O���p�>�)���l��g[:|aӋ��kC{�t��7����o�m�hf��gOy=�=�i��q�k.��}��q��#��~�u���d�4�J&i0���w����3�D��OI�<�M�y�2�M�����GV���QkG^yO0�wZ�U����F|�O������I�2X�gs"d�]ޗ�t��6��I�N_�=���
&���n�H�]@�I�D�$(��o�	h��i��w�g4&T�)�]R������=��~1X�W��{���*���[ku��!>�bf�|0���P���d���^�#��l4Re��xkKͺMq.<����B
]�Y��C�[L>[6�v}���E��y��T�[��d�u# �bgh�7�Of((����=��4qP2�����ݱ|ql�.�Kxj��'y��/�R������_P��>zj\��5m۶n�;�i�.e��O��ZL���Ə6yt�:>/ܷ(�C�6CG�@�c0����(�#��yku�u����<�h^^Y�f���ڂH$�K��8r���M1���l(�jA�}Tl���Yu�vh�f��O��c�G�B��!Mu/.&ia��qY��ua-I���c��45�o���[���%3�0�B.{�:��%�IHM�%3��T���{v��r��e�]0�X4kF�|>�5_n�)�*�����|A�=7��Q��%�S�����IT���u^)1z�)�8ï2��O8��m�q�"#H���:���"#��"":�6�����!�!Fц�#(�#h�#����<�#ͣ��<�#Ȉ�:���"��P��":��e�GH�:�����4�#L�.�DS(�""#��DR"4��0��":���ڑ��eF�*U}B!����e�a�Zu�QE���Z�������"":�-Ÿ�-�,<B�W+u9RTZ�˳TF=ϖ���̝-��Os�X�4��j_�D�8���8���!*�!r
�A,�u}q}��/+�&2�$0Ce�~���0�4��yd���o�����ǧL�6�L�E�m7��[��s/�6b}9�I�@�LL~d�	�J@�O�>d�x�ѺԀ�"q^u��S�j$��o�>�g�\,-�0�k�F0������h��h-�Ϲtl��
e�_T[f?\㶶� ��`u���ۣnS�~Bu�L��jW��������l�ѫ�0{|9�C}�a;7<�1�{�o���O��L=�F��3ɑ3@�����RI$�3@�����RI$�3@�����RI$�� ��ww�^׵�묺˭:�������-h����q��SNJ�Rەb���$�!$C7f���/�ݲ��PǯӇ��5P�s�>Qtӛ�"���~Ώ���9P�RΞ(��\m���Y���^:qw������w��C�'ͥ;/jr&v.}��q�r�җeH�R����GҬ���a����<jö�Y��m�(pޤ0t��z7�u�<��k$WO�F����א2�m�#|*cZE�����}?��Vr�$_��Gt~b>�D�xx�v�,��d6wcwGj��@�C��l�h6w�O5E�aeY�u�(���z��L�e�\iռ����Z�G�6p��(�6��H:�6ߤM�����V?0�ZV�<�����{~�BHI	"'[��8l�Ӎ�UP�6�&��I]�l�yt�<Qf���^l� s��{r"D����ɩXfv��Yj��m�;?���~>[[z�������C�͘��f����6�,���m�J�R�m�~EGƸyXrq`�6{R'�F��e#�_��C�rK42h�>��NB�/�R���KФo�C,!F`�h���$	l(��i-�ମ�|�у)�q��]y庵����Z:��y�Q�g3��{�W{�q�2��$�
�L�Z���b/����f魽b�Y�K�-m�tx�j<�{�����D�L�Ԛ`H
dj��Lu=[���b�y���f�R#P���[�ݬ��+��z{�Ӷ�i���5a]K���* Ͽ�����^^v{��"�<��00{-�+/]wq6[���ߚ�F��*6��a��Z��	��f����:�xl��<h��F���Z�{�E�Y�L)+�ˁ���q`ȝ�uQS��]�l+f9>u�8h���Q��������n2o���mh^�y۶�-�N�v�'����c!E/�|�{[��^�<�*+��]�=c>�2� �x?��UV>�0�j̼��[������V���QkG^yO8˚���y�rL��Vg���BH��"$�|nC�|Rً�'��6����n쎙N����^>6���`��ݫ͖�m5���2�z��.�weQe\��4��8shƭ�U36�;.�$��Q�D{a>�������r���U񺻊���h>�~0�j���5�||P0t���f'd�ep~�	�,�Dʻ����R�����^8h�M�XipZ9�'��W*�EJ�\!�����0�6̹�����(���0����#m�Z�n��3���6C�
6e�h��-��Z�מS�r���n�3�� �	 ��JIc�`/}|Lf��J?1��)���dG�--���F�����^��k�p,:aҶ�P�[�:3�^�~��]��hN��Ņ8��pQI���χ���cD"�"���=O;�F烣��ƭ<:l=��)<�n}�GF�uN��^����Jǈ���4ΝKB�o~6�1�)h�QQ�\e�E��[�Z:���<���`/��<�!
�{���4�e�c������Ŕa�a|E����;�K[ʮ���m�����DC��u�ʝ����t�F���Qlj�?O�+HB�g��
�Ȭ4Z���v�P�Q���}A
1l�ׇ�3N��{Ƙ}�&�x6�����xg��jΖ�t7��㵊��O�T�}GM�Cz)x<k_HߍT���1^,;�=�\lt�A�>�./�9Ug7KO�꒡A�C!�X�(���e�pa���J��ey��士[�Z:���<3��*��~O�!D�G$nJ�?{0��LS1IJ�Çͷ7b���r��/{7[�D}N�@�����tt��Z����>�{y��q=Y�ݦc6x�kZ恶�b��%2��O;i��� �
�y;(u��Ӟ���ڮ'Ll���I~q_��z�!�P l�4nw�]U�t]]��6t�:�]W3m���lo�����rJ<����w�?}<��+��G�8㬳�R|��9���c������8�nH2ɣ-/��p$;�7d�E�����#��6Q�h�у�>k��s�{�0��ݚ_[����ԧ-:|�x��6ATǄF�[}4�j�a���p���B��>(�F�G�o-h�֎��q�<���}ԧ5Y�ww	!$$��K�������ut�(�䯳x�K��ߙ�js|��Yj/��Ha�,(�F���΍|�\G�7���vI=��>*�&��Lb�ӆ���ͥ��GV������3������������Vl�&�||t����r�Es)�	(�JiF�@����HF|�@����д�޾l��
;�8��کU6����xn��a��7��:���HxQ��_�k��Q%G�C�kB	,۪y��e�^Z�E��X�<4p�G0%jϩ�U~;U��-��BHI�8Z(�}�C�;�>�á�F�x�A8bၚm�o	%�������9r��}gWWD����k�����\
[>��U���F�޶ L�hT�������ߨ�����p����l5������XÃ˥��CPᣜ#͆�ms��/��ma�
66a��څ�Vi}�;�#*r�z=��㪾�|5��O�RߙFQ����Z�Z�Ş:l���4Pךj�2`��m��<@!F��h�����=��	!$F�QZ2�l���p��vyx=ͽ:��?<4_Ԧ}��$>48ww�����e������{�;Z�?f~��u�������G`��:;�D �')y��R�ƨ�㥏Ln��Vq�Q�2��6���!�����Ӈ��|+:�:�|�woD���G�8���Q�::�׈�3E��N���޸h6=��e���#�6)�4�:�Ѥm��[o0�)�DG����Di�y�Ѵm��!mB4�#,�4��(�#��:��<�#΢��uDDy�u��F�aGXB<�FQ�S����8�#H�4�uL���"#�#�!H��"8����:���4��)�aR4�!C�"0���M�8�#�4�κۮ�<�u���-kikDuDDq�me���ͬ���;��u��G��U�Y	t`{x�d�C>_�s�$�UG���	 `����)���N��;�A�(��U^�Va�uչ;Y�q�7�3y�x�?t�wn d-���A�󇆠���fS��a��&�V��3.D������}w��{�$J���T��Z�kf�R3!$cTdjg�QadI(��`���;�a�RbN�	�a"4����_jǎ��?�J)v6�jH~�D�bmX!�{�:�G)����ت��F٬!o� ��ry��
%
��	�����ꨬ�䎺g����A�]��ɸ��*�	O����Hύ<��qdh��(�G:Z�z�"Q@O�d��a�\2i��5���~�g�`45�N��X�Ʉ��%�3��#26�չ]��A4��Gb��TX/���F&��f|Z��.O����q�YY�!$3&B�k���oI-,кӿ�d�`��� ������58�G[�c$0�i��e
Qj�#e��>�&$0�5�Ċ�4�T�io�h���s�K��X�|�O[+N�eK�@��o�q�������m���K悧�O�>���È���Aq"C(��E!3e���wkː��a YP8�N҆Y���WΓ��81CI$�b�܇H'C9A�gu���yk4��"Y`<�<.42UZ��Yz���:��e�-�m+�Ƨsa����$4�e�͟F#� �t����������Y�Bћ��9��t~�� �9����5��(]˭1�b���]n�u����������:L�2||(Ӱ]��*I$�1@�.��$�I��hwvʒI$�P4��ʭ����^׵��n��:���[�Z-գ�<��e�N⯋�Lʄ��v/��X=�w�s�z
����壀51��]�n��*���Z��/"J���O���ʅ�V�X^�V�g|ݽ�W����y��b����eXr�p�v�c������"���{����:c����6(�b�w�K�C�{Og���Y��a]JaD���ix�3{�����"ͨ�y�X{�]?}�y0�^&�W�^������Z��Z��Z��'Im�R��P�L%A�?�_�v�_Fbm���KG�u����a�K������:�+eƖ��E����ԩZ�^���)�^���H���߾yl�c�lm:l��N� ϕ��#���C����]\�	+�y�&��(5����I��.aF��m��,�;�5̿Cg��R�wdq�T����	���P�h�H�5ϲȴ�-2�xĵ�����e;���v^L�^茫����J����/�Zǲ}�g���D!��3��D���Ua����ֆ�a��龖tx�]1�^4`�x�4w@���<Q��:�ַ��[�G^yO:��7��1��[ԽI�]�C��e�,�-t�TU��utTpj��N�[>]:N�l��a����᮹(���v[\d�����QF�!�fчB���H�&�D�1���B��� \gL����^]e����s��IִiaE�q�3��llѲ�bg����>z.���Su��8�i��C�*oE/6C�u�Lc,׃VBG��J�1��--���φ1�akG��������L���q��8�����מQ�e�SM�5�N�ci��291ݚ��Ȇ��?2<�/��|�F>���n�p5Q�,d:X����e6�,/Y���`�5GN��a���e/���eR�+Q7�4�\R�CmʖDU�Ͷ�Z����}�]���q����~�7��K��������"�
9Ӂ�M�0:��h� w��v�q��ф"��z��Wӭ�����>!�����	%,1C��YLw�g������>����n�~���Cf���sKkAÃ,�F�6Yǟ�Z��֋qh��)�Y[<��?E:&	!cx��[��I����2�^��6iI	��&z'
/pB/^�k�s�[`�������]_�}bdT����~�H=��1�uop��g���YbF�7C�嶳��q�� rV�ig=[��@��H�����!ʠ��g�h���# �:~7�fy�țl�m���tp;��P�}�Q����۪���׷#l��҆lzY��L�aҎ���Ϙ�|[��-��]�;��p�&sM�4pލSG�&�qx��l��7��m�J�c��3��[vp���0�o��kٮ�>:�=�ߴd���lo�'�c�H���r��%��-�GR�_���2-c*����7�uwCT�6S��fͲ�/4��-kykE��u����*O��ݻؑy�Ұ���OĂC��Y�W��F�43c�g)|c"�[
�����mL7��I���kr���]��;]����G�&M�}�dg����77�=�]�7|0h��e����ߤ�=���y��6�/��l���A�� ��/��`�D�	�N\���ߨ�ےH8u.��t�5����3HáF���v�l9����zv���Q�FD?�82l�O�ҚF[e֑�q�kykE���g᲎l��zƬ�yy�:����k��xaS�g��e܌s�e�/������L(�<�����d���J�d��3�Z~� ���4}�?~��g�����*dP�2���A���vUI�|CA�n����Wy��F�h�ӊ���a]ʅU9Bp�y՟��3�M�9���vEЊ�A�n�g���&��F��d��	j�
��$��,6p5gZ;�2�/}�#2F�ˌ�/4���~Z�Z�n-y�<�,�R���UX�3��!S�s<o�ccca�/�Q�|o��V(�TyVC�}­te��|W:�8	hze���B��"�����>���������S:!w�@��z� �����?��������8w]���F٤>sB�d<��5�J�:�+Xp���N��D:3����p;^�y{��t[l27y����4w�>�6Z�>�P�`̿2�(ӯ�q�kykE��u�p��%<2�f���6����8�^��1d� �j�3�K1D�T�IUJ�u?��BH	Y������uc����p�*�B�I.�?Y�_���h��-)�X��`�PA ~��u�F�HD���0KA��ik-���mF&�Y�H��� @�'}���^6��iu�ݱj��_�@�q�D����Aߋ�{6I�D�~oƺ6y�������mXup7�~�8�G?��<ҏ��+X'84`��v�tʻ������s����z8�m���U�663آ9�����Z?{��>D�ϝ�Ho$=?y�s��ul*�pWX�sO�z6����6Q���8N�J*���QU������!�T󌭔i矜~E����Z:��y�U;y���O��P{�o��666�}�~>��kF���L�"������Q�|l�}z�U�.����"�Y�Q�a�ڽ�9�IU��۱�g	ݶ����1���?��6 4v��X�]�5�z�����=?�M��X(��e��
/��]7��fI�%�����Z�)��`�����L_�y�p�*j�#�(� ���n9%�/�]��u*����/֛�U���#qQF�fݜ���}l4�5J���.���ǵ��83Sl8�4��[�6���R"#h��#�!DF�Dy�u�me�}B�Q�2��H�4��h����Σ��<�#�yG�um�Da�DFQN��DF�G����mF�i���e�qqa�DF��G�G��qƑ�Q��W�F�#JB�8B#�H�8��,<�먏#�-e�l-kmkuh�#��h�6�B-M���8{&�߯�YI}����k� ����h$�ԉ��֌z9�ѡV'�9���eŵs\E���Y�W>���)d���=L ��&zA8V-��RZ��l~6�Y �g�9�eKRҎ���Z'��*/����tq/��|:��h?c90�!`��<�X�ϼG���]����;�|��l�Z�Q�23(�ݲjI$��@�wwy���I&fP �]��&��I��	$�$�Zֵo��u�Yu�V���kE��u��uw�ֽ7��֦�Y����ia�ΚE��9�r8p4Y�(�ia�y>&p8@�����n6F�,��mC(�����l:e�8W���6�cz"�u)�qӪu9]T[�����{������������t�7�|��z��63˭W� ��k�= ����4l<S�z��&���眒&wy�������Æ��ؾ]X��Q��uh��:�Z-���<3��*�ol�-�����`͡�=�.���#m�iiN���)p.��Ø������q�[�7�v��EP� [���l�|A��M�� ��ᮑX��uCg�OxU���]��w8o͍�A�p�9��e��t���P����΢��Mt��g�W=t�e>�]dɷ��d��,�X�0����e�?���>\,�c�wcogN+��G\S.��^iZ:�Z<Q���e��Z�r�5++/�PHX3��0��
�;��'��X�k9UFL�	[)H18_ʱ[1�dy�ef����@��6M��uy�)�g���W��V�/{�$T�kd�_��t/��	� DP��G,�q������y|$�(-��)�(D��u��z=���� ���I��:#{�.����3l�OK�z�[����C�>!p����a�ぢ�,�ZAKF�>��Ƕ�P�
!xrȭp;��/���h�X
þ�I��CwE���h�r�a���O�V��<n�C:݇ǥ]�FI��E�Sq��5�������ln�&>+o�(:���uh���5�W#����vp�4x��,�����Z�kiy�<�*�w���)b�l�$�Ho��/�ȝ8��t��X}w�6��P��>:Y>
/��p�,G��ɮ�+_f����2��O��L��*Iu{udj�cf�����u9B���y���V���n��%���!¶����Y�T�E����q��j�5����k�w��C���2�PTr})�I?x?h����Tx.�\4N���F��CtgC���]��Iz׊0�=�>_1�c2{Lc�>�f��*i�,�*e�\em#���:�Z-hۯ<���9��(�O�!�2�Y�$�H�S�L�<����A�wTS!�pk�:x�M�5^���Z9�N�"|P�4��b�_'����R�9ܟD��w��륚v�e-[t9�g�?��g��H��Ϸ��/d�nxڃR�+�l���Zryb�������P��$p���Ń2@��{��EC���T�h�Bώp��F�C˦�N6��u��G��Z�kE8p#��'������p�%�6�����m����x�qQ��dH�m�Ћ�c0�Y�{6a��
��6>Kqh���H�Q��b���q���!���.�R���K��Ep��}0�Aで�9;�O�7��4oLl�f��ᾜ"�5�x�Q���U8��wE8;��'�yFJ��>9cm������!�5�����뗗���ʝ�G6Oa���<ˎh�X�4��gK\Dp�UU;��a�2�.��O-n-DZ-��u�^���{��s�H�e,"�4�w�al��Ȉh6�ۙ�
�HESi�ĵ�Wʂ!I}(���PHTQ"7�9�ɑ����L��%11d&`H�E��0�?�#�"�r:����E�X,9b�#����e�	%�	_K��0��5m�nik�i�ڙ�� ��������R%�a3����￿~��>@`��R(��<����#�H��gśŅ�����<���t�3O�5ٗ%�����9��υ�G���j�|4�y�:T�﨡�3��-�(�j68Z�Q�x�o�%��n�/�]GX�7���em�xnQ����1�	�C(�υ+���D_.7��p���d��q~ׂ8�y��_�E���uh����A01�{�C��y�=�0��I$��I&C�F����=�Vm��鳛�JE��d��p�ВAp�O����l�Hх��1�U.��a$'C��t��ņ��Ҏ��I�έM���D��}__��.�g0���k��j��1����='Wwn�n"�u��#��8Wq�a�O��U�({a�Y�Y,�YF�ZnIH���QDY>A����޻Vfs�xgó�H�@���5�0ҝu�u��[�GQZ�[/:�\e�}-�5R����c��+{~$�H��+��χԞJ�=�ycz\B�x�u���\.��t�ㅜT����p��X�t�<M���L�V���3XbC2�h1��j4[MԶƶ��*-��K�FlÃ����ra�f�Eє�Y�5��[��|���v(���ѐ�g,^�|O�o���d5P�b��tʶ���=����Z���Ui��^S��y�Zy��G�����u�R��s���Z�\�J-�Vsm��=Ѿ��!G�=�UƣlF4~�ܿ?��x�^�/��������oí�b�Mm��(B�Zuյ��;@�>򓲇y��.,o�k�c�*��(��*��ia�Yw��C�{;��+%�:U'���&p8���Ge����OKA�A�ZJ�nM,E��'�ϸ�S�F�Zo9�y��w���������e4���R��M��.'ݽ��}��y�u�����K}ǝ՝��Î���`�!$�'����"b�����w�bCf�`�n�A���MdŐ��y�2ɭ��bд֘�օ�-5��֘��Z����I���Zb�M[D���kI���KE�$���I6�֚i�h����$�Zb���Jb�ZkI���Ŧ�֔��N��D���֋Mi�Mi%�-��D�ZkE��LZkMh�B�S��E����i�1i�5����ҒIh�œZH�$�"KI-,�ii"ȴ�YZ$�-���Ih�ZH��ɊIdIiȓjIi"�K"i��$�I,�ZL��%�KI,�DY$Y$��BI"ɩ�MMi��Mh��I%��Y$��h�Y"ZI%�I6��I,�K$I,�Y$��,�A%�%�I,�Ihq6u�qd�K$�Y"Zm$��Id�d�M�$��Ii$��6��I,�Ii$�BI%�I,�,�mm$��I,�,�m%�I-��KKi&�Y$����&�Y$��%��Ki��I&�H�KKi!�l�Y$�d��%��i,�$��Y$��m%�I,�[I$��%�I,�,�Id�%�I,�,�[I6���%��K$M��!$��i&�I-$Y$�H-"Y"Y$�IdőiK!��6F��Y����dk6�5��#M#9�5��fF�h�4k�#M������g6ѭ�o���F���ё�#XF��^q���qn�$�&!�3�F8k4kl�adi�5�k4k�,��hѭ��#A��̍l�a��4�5�5�4�i����F�F��i��h�F�F��1��ѐ�g��m�h��di��F��i����F�4#Xѣh�ѣ#CF��CC��b5��6F��[4km�4��F�!��l#[4k6�3F�h�:#8kh�h�؇H�m��6��!fг!l���d5�B؅�Bƅ�Bl���e��nKE"̅���!m��!6BƄ�ɲ6�٦�����&�&�5�k2i�l��l�bkhi�&�i�ɬ[i�[M6�L&�Y��&�Mf&�i�ͦ�M0��F&�Mm����2k�m��d�bk�4�	�&���i�M�d��Ѵ�ؚm�������M3M�	�ɡ��&����ƚl�2i��d�4�km4d�FM15�km6LMa4�k2k4�i���M	��x:��ܛs4�i�&�5�h&�MbkdѦ�bkm5�i��i��l��5��m6[i��[i���i���i�&�M16[&��[i��[i�&��Y��M	�:*N72h�ɤ�qƴh�ɲMi��M&�i4��D�d�i5�I��MZi6Y5�I��M&�Y4Mi�D�M&��i5�D֍��k&�I�5�I���g&�4�ɤ��I�kM&�e��kMY4�&��Md�&�Y4Mm4��"E�e�"ȑdH�dDYdH�&�DE��$YD�""Ȳ2!m,��"E�H�D�h�"�$Y2E�"�$Y!2�$H�$[D�Du��tȑ"�$Y�"FYD�""E�!�"$YD�FH�,���FY$Z$DP�6�kE��$e�B�d$Z$e�dDY-�#--	D��FZ-�,rr�"E��h��d��DE��-��i�,����$ZD��ij�@�B�"Б��D���FH�$ZDCYE�d",���$,�dH�:pt��3�$Z�CYD�B!4mdD-���,�B�#$DHZ$-БhD-Б��і��^gъѭc��Qu���F�6�5���d5��Z4 ��5����$Y5�Bɭ1dZY&,�ɬ��$Y5��MdD�ZM���Q���"S_&��F.�iGX(�c�w���d��6-7u��kz:Gw=?ß�����W�����=G�7~z�����:=�y�{?���{�������y���g������w>�܏S��ݳ�G�OϞ]����קR?S��\(�\G�$���?�)�~#�,�{�����3Ӷ6��sz_w���o�����Fߛ��>��l���x��ka���B�l���f��������|�f�����m�ߖg�n��&������[��}FϏ��m��{so���O�i!����to����~߳������n�YgMm�g��w곙������c�=:|;v�x���{|f�>���Ѹ~��e �[N��������t���N���l�i�t��Q�m�L�cm���9���m�H���6��h�u�S3k0l(�HB͆/�H���Ҁ�A�C�JPEA�N����%�S���^f�g!!��$�l��1�0�ٳX��l7 �s�3$6�P��5���c�����5��;��}��A�o�l�|wn��޼yo9�8ww��i����w���6'��?�}N�m���5�6��|��^���7�w���?Hw{�K��~�?��癞o��'q���<�|�~�v�.��oyտi�����<�={�o����c�ߌ��ߗ��G���lS>�mx��>D}�ϳ���_���<��!��pݯS{;����Ѱ�������m�/����7�p�t��:�yo��z[�����q�]�A��3�C��$,X�?d`���L���I���x-�؍7A����wm�=�P��B
��h�:"/熐���7���L�+(���X�&xh������Ͱ9���>վ��尾�����ç����#��z�=������Ǐ�~��}[}秮Ѻ�>Y�t�y���oi��7����ɶ�ם3�7��&������۫clO1�6~#Dc���'���l6��7ñ�>/�lA�|�=y�=-�=F��g��ݍ����͸v6���/����-��v�X��A~��
�C����/��<�A��~����?�h���-���w�Ť�I �O� �@���\�r�v޷cz[�y�@�y�ޞ��ox}>��x���|�'�L�Q�n�Vwp�;��^ݛoG�oZ̳a�s[o˺o���ݞ�?'��ݳݼ��lަ�l�#�|6�>n����{}�ou�g�}No�+Oǜ8��h�m���������w$S�	�.a�