BZh91AY&SY�[�_<�_�py����������  `�~��n���P)A*��)A@PP���
���(PJ� �B��@P  �!�� :   �>��0�� ������݌�=����ܷ���f
;k� �w��o����㹐����1�L�[�]� 0   |l�ݝӜɻ;���\��Uf틷v,�]iݰ�ڏy�κ;��j��[�UB��cs�v�vmp �  x�<k�խ�:��aw\����m�;pp���� 㯎�֫'�3���[m9tlݚ����8�  6
��s�wsV��;{iWv��7:ݝ1|�o�g�v�k��b�mݺwu�����9�u��i��  s�>m��}���ۯx{��z��ۮ��&��ӊ��*��zwu��Yܷw:ݮ���;�tͺu8       � 
P� ��L�T�z�Q�z�	�ɦ@�L��i�HI*Uz��0�h��0FC ���6����� � �i��j@5*� 	�� !� 	� D��M52 )�M ����ЏL��(
�i*�S  Ɂ4���!���ϔ��T��~�>�.^&� 
X?���H$h�?���G��R�����0�Z�����0����D�Hj IU񔝢I$E�T����fU��l#���RO&��UUU~�0�H���ߌ~0��~/Ï����Q7nI�ײ`��&�rQ���j^�1P'j�5��T$/4)bp�4τ'ZݡP���L��D�/ZB�'bY"bڴ�"�[��-� X�R��Er&*�jQ���B�'(�	�5
ł�o�>�jiU&/R�P��S5j����(� �=���x�(�b�w.q���e��4*oUk��R�̹�+�:�J�����s���x��7<\5��[�b���,��ϕ+��a�嚜�}�ov�%5�,�ܪ�;��/N}�j�X�^�JM��g� �C�d��lY�l��Vkn-����F�!=��7�S-8�cnF܍=��6R+)���ۍ��w��T[z"1��������^cu6��5n!�~.��ܫo��j>1���dSy�7�
��Y!��7M���ך7�h�C��}�x2y�������$.F� �[�η{kghK�ˋ�y�>���ʸ��F��u������oI���s`�Cz4F������0sǧG`�k"�x=�<�*B��\�t]���asÐǣzy��k���}xDKE!�����;gc�"i!xfp.6�m���	X5dV*� B��ߛʦ�P�z�!)�3C�@�3X9�ÿ��8�wn��nzc�m����ѻ&�@$	��K:�4�O
h�*��������8�r[��f8��/Scr�7l�2�AP�-�r�r��^�l�=�d7�h -�B��O�oĸJǃ�]����dEg��x��;��'f�nꛕCx</4"bj�PQ���a�)�i!<Hj�66�1�d�y�}fF9fη�����m�ۑ�Y#oѷ��:l�n�Im͡�L��}�3���q`��Ũ���&#nv!�Ԫ�r�,�nrq�r7ucu7^^ߴlo�&XI�V"��i�l�1���z!����uN\���<�y�ڀ��C�<ۮ�qo=��H\��0n=���-UN6�sniڱe�ز^��2���	܍�6ﭻ��d<7���/`�T��p `��O�vuL2��S���	���~d�>�*�!��V:�T�)�NQo~���}"tVxQh������?2�����<OɀU�q��n^�EX;"�H H�t7zߪ��P�z )��������hqc�f591�=1�[�P �7�?�L�L= ������cA)�M�!y������qv�;1�l�屽o�hƬ�5M���n�]��6�h߉�{��j����*���kJ�c�]��v�2"͈�b4�C���7��P��n�]��E��PQ���e9C�&�M��ηke6������žr�N����P$m�ۊ3BFߣo#鳭�M˃[c��vw�:<c���sI���7~����
��!ı�/åP�V������MQ^��y���{�>���|�MN.�(�
��M@���Tjs:d�Tf�[<=�+Qv��mKA0Wê'��:�����6�Ncu<=�,t���z7�A�ށ4[Yp
Ydj���EJ=n8>E�-K�r�Zoȶ)F91����v�=Yqh��m�*@:��������Z�:L�ډ�*���8� ��yT�)]�6�p��ѷ���ߜm��ۊ�W��*Q�q���b��>��FӘ�O.����^�oЃ"[y��h��#f6�qc�E������
(-�ھ��Rͬn�Փ�������9f�y�ɍ����n`��Z����G�ZD���
����tv���X��Z�E�
q��",��&+F�5�*D:�qHW�]��v�v>N)�9-���U1��6� ��/FߔdZ�h��q�V:��1_
Q�q����\q�pm9������yj��z���
ɄSM�D�a�8�'���PO�77����u^O��J�*��l��ʋLDM@kQ��TDY��^���cj��7���h����GyE&�U9�(� ��ǚg�6������Q�ْ�+BX��7Z'"��(�)�.w�X>�����P[�u�_Gi�n��E�T[�a1�b���-��؉�f���x�j+�.�j'c���O�B�<���T�ڨ
��ÄY�5E&l���*�Դ�_��v����\q���s�᫴E���,Y��Vy��[�7D������CU �"����e��G%%t�JU)
��1�cw�&(R�-O��(nP��Jb>��v��9Q�~�=Z�U�b߅�j��[D��J�[��sbQ�- ��Ǡ�B����z�U ���PB��P������D���c����̒�ܬ� �����M{�c�s�Fq�E����W�mƍӲPT�5�]3_/$E9���U;���iʕs��0��dt�sD��ټ�o+v��勼��6չ�G��
j�>��"=7�^ד~���<��u���m��oo}�����`U������>������ �z�o}�o7Q1�N��y0ܸ�g�v����Yg����ג|���5�/7����p�˳�	�ſe�5q���ܝ���>��A��>G:���Vҟ^���{~�{�SI�-��]��y����a��.w�&o,��xz��z��45�����mS�j҄��߾�rs�w�T��[����'��YDP���gު��87��m���������S\9����'U�I��ׅ�w�_����6N���C�Ʈ&��S����vt��R��UהK�l��z{�b*=<�v�}u�?M����z�\ӌ����U΋��M�7~�N�4����W��_f��j�c�s�röM�G�"��NM��}������.δ��~�p��rY+'n�Q��y��\���9�vE��Dj��VDV[�S����L���Z���3)�^�Ә���)�c��U�:�H�8�����w���͎[m��Z��g��sIs!���p����8ػrN�r�b،dڙ���v{�G���_����٩��N�{%g�ADo�ez�����S����tҞ��%:=���{�}�4\����z��"�α�sO�iY������k]��g9�&�{��܋���;��A���6�(v�_0�>\v����v�o��9�HU��[ӗ���x���K���8��pׁ���o�q�[��k��qӷ��a���x�$��v����z����!
��o��V�	uv�x�r5�j���j��0~���2-9,L��+�^A�����}�^�����{�w��~��<>t;��]���s�~�}���E��6��R��E��͹~��S�ׅﷻU�}�V�y��n7v����u���o��.<w�9�7��Q\��r���������9bq�}7v�~�8�;�{_/�����Ъ=n�9��y���]��x�N8�7mW��2�ݶ�TV7*�UE�U����}�M٧����Ħ�F���{�^��y��+����ն����xp|�A��*s���u=�ٲhE��͔�zξrl�}�>ݷ�]�{�.�/�߲J��m��g���ُ^��L�w������^��Z��6�/6B�{)�s����^�LZl�8n�W:���5p�>�p��޽����զx���<�ܽ���,�?:w�Н�T��wˇ��ˆ�^�l��y̶��tQ��V���ƈ�/'�vJɖ�W���f}���ڷd��zלu��������}������G�,�9v^p��ǳ��/���]>���s�T}r�}8K�����G���O�W��\���w��G���r^~a���-`!���H/��!r�k��ܻ�M��9�Oz��cP�{9ge�ع�ݗH��[{��z'�5��)�$���+��G���ߧ:q";v|׾�>�~��_t�\6g``��H����������ӧc�P�0�;�/Bvl�¨����뽝����Tns�H���nc�M�/�(q�>����~������[�UW�a;���Z�T�j5����Ox��te��t�ݜ���TF,����	�N�.ɾ��l<5�Nݑ�U��[g�zU���5���c�;�p����F���[z��7�� ����=�)�ͻڤ�����vum�9Ȼ�C�u�y'8�t�y�~��6d\�t|���`��!�9�����'}���Z����Ƣ䢇9:��a�{�����{�k����qm���a,�5W,�;��jq�o��6�ǜ�_+���.�;����������'���75�*�_�r�)��ޅ5yŴ�%ݜ�ޞ��
�i6W�����
vo�Gͯ��kה�4������r�>���w���κ}s=�M�n쫛w���rp;͌�-웼�K�ۍ�CW������7���,���09���i�ګ�L�Ӝ�<�_���ܛ-8���T��+A�x��j��Iy���7tP�w���sM��f@G�{y��ol�o{���@�8�S�m����_9��yF��������������O�n�7�j~����$���od�qοy�����s����o�h�y�>����oGϹ/�W(����q�����쑵�S�ޚG���ݠx:k����_�QӜ�	w�+��ֹ~~����.�m^�7{||M��I�f��ƚ�J��j#��b<eѳ����/�Ѫ�>��*�k�u��y	�w���n���v!�&|�7W��\�V��Z�CL9��!�Lz�{���P�p>�^~v+�ԽDW�-�c)�������2��n�5�S�V��*��'�V�$�|V^�WUҺVW���.c&U��9v�������^�ɯ^�-a�l���K6q�b$���.��ڎ�����|������s�����+\!Qc���m����~ׁ��Փ�ʹ���g����i�����yF\�C���~G�����m|�>�^��!����6-!����H1��������
�9��� �s�����$j�P����V��;!km�vF-ˢ��Q�L�<qA����~���[I%�:�n�l���9���ﳵ�BL�V��h�͚>#?�vn�d�r���[��{�CWk�ժ��U�k��G/��;Ȼ�\�ׅ,n���c��A1(ժ R���ҽ�a 㶐#�T۔�$6ų=���\�!�NJ����;����P�[d�T�Ae�,�����d���A6�/Ǘ8��{����P]�ɭ�
�$spM���q�Ԙ�"m��N�dhdj�S`Mh瞮����tUc���;�"T����J�k�҆���f���b�k-G�V��;µ7��h�>(�+d��TL�[	:�VZ��US�����RZL�����j�M��T�c$�XԥJ:�FZ�v���8����E<5�9*��FN�8�'{�y�jqcɑЈ%���4㮔v���F��|�x��{�R@�o����Z�2e�K�Y�6Ѭ�­��;%B��Ɲ����T%*EQ'��uGFc`���m�7�C�b�G�QE"j(�
���/������+H�|�)�s�� ��-6+��hE AD6��[U֛��lU��X��ⅉ�<Z�Yk��V"��Un��
6�N�t�p��zn���'���@S�Bj�D&Yb#��Ӳ��7��[��Q]�����.ż�em��$�b�ֽV�X!�#��A�nۺ��TU5߸�Q�ǀ<�;fjȊ����V�	�Qb�tQ;�ᵃJ"c��2&*z��۰�[|I�7�����#������*��
�J������&�°�'�љ��@�Ϡ}�|�hI��U�PG������(����&�~a�`�_��O�?��}H}I$�����/���_�����bf?8 X $ � �  �`   FS3  D      0@
� ��@
 ��wwK�_�����$���I�^T���o�{�ל�9� `x ��< � �`  z�@, � h     �  0 , ޭ���4`\���UD�;�I�s]{� ���  h� 0  �@ H@ ��  H@  � X  ��  �  ��{��|�7Ü�Tq\�Z"�i�w��}33<� 4@     �� �	 (=��@ H@�� �` h@ � X�  l��nZK�M}��|�(�̀x , �  р@�� 0  ��� `x �@ H@@  @H@� 4@ Y�����I}���m%���d��� P�x , �    h�$K�{�   h�   `x�b@ � ͍����$���5H2Ao~'��?ATH�H��������?`����>�Y�,}g�?��OO^������O�8ڸ�㍱�8�z��GW6��������oc�8��<q�=q��n6�tS��Ѕ�!J!	Z!�P��Z�!
֬B�R�-B,V�HT��N1\m\8p�tӧ�x�\t�q��Ç��mi��>�W.[Ϛb���l��աۛZݵY]tT`ۭN�O��X�z�+�ah��$2J�evQ&�Tm��,[hUu��ad���j�]bbi�V	���NKM�iG,xܬ���T�ڝ�����鰒D�R�ꏺ����8�#�E���⍣knV�X*&���7"p�J�N�ʚj`QAK	����[����	8��R�e�����4��&�!%�Bc�U�&J�2J��p�]V����펻�CpU1�(�S�j�KV��&��Ok{kj�v���9�b��mj��Ӟ�	U�y�'ƞ���$B�x��֣f�U�-�Kj��6�m�:X��Z��:��Z�#�:�ze�PdcؙULn!R�!ʮ4���5�	G�1�"�ᒼ��R��2��Cj(�P��q�Ut�JA�X���}Sǆt-�M>�]�/����l��7D�S�q�`���RZ�Ur����ع+����c���:����zֳ�/�M� �ww��kY͗ۦ�$���]�Z�l��7$$�[����{�se�鰒L-��/w��Y���H!������ʵ��h�M��q��;K��
��5�mAm+��IEkR2F������h�U���)W�H*�W���#e��L�⨩�H+vW@��AJ�K��F���ڃ�IlJE$D#J(��������DH��|jf� �͒H|[��BR�Bퟍ�A8a��F�Xw�I�qK�0؜r'���T�ʕC&�i�N�!�F=�T�LN�#�6i�⪽gy���8�&a�|ð���=U�D�N���፝���ə���-�0/@L�g�޵r_�������Ym�TZ�TH�v�q�W�P���J'aP�����w71�⪼v��Q�� ���ɖa�ل��i�Es��%lX�p�a��A��2=�C��p���b3Z{i���b�c�G!#r(���)���;��&�n*�,2�6LI׌�%%z��2̸0�7�����Ҏ�P;�(((�8p�E'{Y��4t'�����Er.��!��5�
}f���2�0 Q����A+�.���qLxY/�26W	��@����Z��n0�\�n�Mȗ5�i�@�q�\�������M5ȮzrY�kL\��,��"�Q�H.���+�n�4L.��N�xJ�탦�v���[�Q�*���̠L$�ch��`V��i�#"�M�⎊i���`>*��qN*R[r����j��֖���v��i����hE(F!�z������mDMB�ϞwD<�/X�V�����*�:&��"(����4�cU\B�aM0�UW�c��Ɩ�%!��+���1OjQ��\媥V�p9�)��檸�:F�cx���aZ��Q�fj�Ub�XUmU�T�X&6�fL\Դ�:����̋[e���ˏ"�]2���a�*�oZcܷve��d�P3�E$���jI��%�T��(�T�Κ9�3��9���&1B�6���U\l`�@�BX��p\&��Tʪ��)��[P�L1Ύ-n��t��æcEv�h�=qT(z�0sa��a�P�����QZ�Kd����rͻ���-ݮۘ���w-^��' q�m,�44�yC����J�6�v�!S�DD���3�:���M�$�j$.�QE�P?��[�x��\ �x��	��ʛ˫u�H;G�c���Da�8D��(�[���f��U�#'&m�5C�����.���䲵S� ���BR�����-��.Y��L��� �hONN��X8	E���=�����&T�]m�i��\K��b�q	|��"9�	6��$JD%��b��<��~�N��ޚa�ոd�tW4�N��ZyXJkA&�p��r���hL^\N��4�� x��aS˅��1Xg|�;���5,��MQTP��ƨ������Be�Y͛�h�L�8Mo��c��S�cnZWQ��j22�;���|�4%�Y��E�c�آZ�؉�T|���KlDKK|)��b6"YFJ*��VF�>+���'�J��G�`~����M��D���Q�KM�R6%�ȝtQ��4>�(G��+᭫��;���\ǣbX����Y����X�أc,hK]c��ݭY�h�����1�UUt�\�՜������k�e�b�MQ���ޖ�]9(�6�6*���-�*�UUålokY�Ȗ`��|�ǳ�~����a���z�7_��Do��~^r��ؼ������:3Z��켃T\:�Ͻ�]Mv__K�կϯ�Z_q>r݂�K�þ~*:�yz��ka��R��y��x-�\@_ؗ�&>/���ˍ_գ��G;����8Y���߹�o�������-������z���/wwOe��r���7����ww\��"����ww\�� ^o������wt@��T��0"`�%�0`��Sm/0(��)�?	��'��pa��I�B���Gc	pI0�0$T���Ȍ��+Pu�r����D��OA	�+B)A�{|�#h#`ڕ,��4��E�׎R�+f����A�(���S,c�D��2��B�;L�$�p�w���;!\�S�+1<�x�`p�`�iԔ0#��'�0`��"�(�����1�3|�+9�T�\�Inl��kV��"T�jk�-	C� Y"�#،v��6"x)B�:R�vЌO�H3!
W)Ͻ�U����NSk��c���!�4�k�4э�G-W b;�>|	`��Ͷ�a\��p��+0e!�WL�pR�ȱ:��\C��C�Xv{>�4��vW��i����ѥm����۰���R���X�Ͷ�¨�VQN���<��֡5AٰR��YH�diH��i�n��|�B�KD܎����O�y��5�wXK MUM�ER�6��5T��[V�ڪ���$� X��$�$M��B��2e���R�ㄊn/��'�nW8�N���$��/���4dԎ���Ǌ<�P(�CՐ�,�#@da�øcL��a��a���g�̝UK��BD����-Ċ<Ԓ��ĕTB��F��N)p�cIMS(]}���GkB���$�J��L  J��;M�����M`|K叺�,zt����,v�'�����ُ��i�o��z���k�TX� u�)�T�8��ԃ�s0*XF��D��(��XG0D�� Y8�n����Q�x�j�WQ5�懒�}L�dn�,{gqG_5�fk\���^X���)ш�Gu@<KP�H�.��jTa�]�O$v�w�	B�6�i�Sމ¡w&�%�nI(�I1�G'�h۵aZi�l��m4�o�ۻ)���>EU�P4�@���/X�����bʣ�3��y�Y���
�K)~IH�s�	,����d]db���$g��4�M��J�� b�S�J�@2X�(�zf�M�Q:Re�z�+�%�R��Fa@���M��P��w�UT�U�� �K4�%�Ҝw1���,\��h�
����=v�M4�V�2�K2�Q֕�Z�l�O�G��G�1���"ŚQ�uw��c��X��8���&�5;*[8Aa{V�0�n�8mQ�&Z�Ā|"giHթV�-���*���H�y�e��V�d�Yq�o��/.�fPc��"� ��! Rr�'��Y�����3l����?8ٳ�+
�Lcf�v�M>ﯱ��̺��D}Nk�����m���U�
��*D��b�Ri�HEZmD�MB��VJXH�r��4>G!��+
�Q�<�.E"
�j��X2��1Hp�Z��%���K]���
o)kh��(ؘ�qf��7L�Z��L��Q�8�j�m3`2�@�^��h6O������	�靔�>��bՄ�K����.Uq}�Iq~���%q�V��m��"I-O7�qw����2<^r;�:yq����4�6i۶�i��V[�-�U�j-�U�T�,�Œ�v��&!1��'���j�qjK�w츹�����t>��?7S�c{�.d��[I~Q�Jƒ����_�bu�W#V�9K(�溘�`��$�K�5�j8�<w�_[��c�1���U�i�1�O���n�VI^ad�&O}W�-�/c�^ƣs���iF�<�~&˒0��<�d�&��i*�����Q�q�X��"�L�f�Y+.^�BX��!.�	�a��6�.���x�^:c��7cѾ}�b���TO��k�77w�0��aZi�l��lcz�u�3\B���'�&/gВ4B(j���E$���%C\UU�%�}�"��(�Ij�*��f(�!d�yXY�����x�bJ�M�ލ��a8����ZK��&��宕�� R���3�ۆd�i.'M�e2[E�:�p�r��J�h����;<Qe�%҈؉�Q@�b����2��F�cBX�eK(ы��,lt6%�*��eK0U���2T��g�(~�Q�Q:|T�L�D�����^�
�(�z���O���>�c<6=CfJ��lQ0	b��4YR�Xಳt�Y��M�ׇ����8���⺺=�Ჸ<��+�4X�lnƼ6t�-���ؗ���*̔Y��lQ�F��l������}��gJ�ކ�6`�f
���V(�`���Q�b}��E�����V��Nh!�C�5
��.�s���v�?�:���=��^�;�2�G�����~��c���ؽ�sv�S
�vs�9����qٯ�U��;'����mp\�_HqTw�\�_�p���x���#��m[v!�¹�|����o[�w��g�'����N���Y[5R���[Y�D�;;�W��z��q��=��{��X��٭��kRF��p�]���bj9�)3�%Ol��	���/�W����5�ݦʂ��QNm;�%o��q�W����k|ݍ���xf�lUNOD���T[:�@'�>Gg�M(	� �MӨ��8E#�.�(��%)|Y�j���]����7�u�׷T��[y���ǡ�#z.���<"�$
�-\j���p�>.Y�N��'+V��V�^M�+�暺�/?N�,^�}\�Tֶ�O[�~�3�;ǰ[|��x&Nmd�����hůX�kcl���Ī;��`����kRT^��j��G�Q�ƝM�\nV [�-�cV�Є�U��s��cP�)�j�m�5#i���R(�n��e�[(����\9�Q����eU��b�L�H����D��*�2�+R���7�ER�L�w5�B�pEU\hB���v:Qɱ�����=��
?e/y����V]�~Eߎ��7���U�w|��F�}���Yww˹�o��wwuV]���}����ꬻ���������7��˶�gJ��%`�E��kϹ�G$"�Ij��V�R5��j�G]����*���ʥ�t�#*�<�i��cI��\r9ۺ�T<�50�<���MURVJ��U��LA��՘��H&6���qJ@n[&��6§ ��^7O����J)\�UL%L��s�Y�c�S�=tv�Z����j� u4�i�ݤ ����Sht1�9J�3�/��F�O�{��ŹR^�?�@�L*����	b�Z�.Z� �ۤ�o����A@\�Z���oN��CNR�2P`.yXV4�ح=v�7�F��k˱�������2|<R���������8`�F���f�m���J9����Jөȣ�׋�G��t��a����I�z���y%����rE+$�MƇQ��E��s�%�uy֤���bD�Iq)p,zK&&�m��u1,p����Mh�C�׊±ZmU�n�ōWٖ�yL�a�kǘ���F���Խ_&@�g|kI����n�	��ozI)),���3���A}Ǚ����Qbf�=vQ�pъ�4�+��x��.:�b�n`�M���$%m�h;��h5x�|������]�sL�d$3��Νٶw?9mV��4���갦�B_.&����?�)���눆F	���Eg�&���{�j�s�D����j5I�E�ӓ@FH�,�y����j�S��N�Ip��wR�����ゟnQ�8/횆���uA��
�+	-��H�.�OTnZ�\7둱��g=��RcpTMy_Bf�Y�WM�6v�XV+M���1��4���V$�d�K�4�pX�5�H�
7������<����Vv R�M₰jH�(��p��ы���.���
�D"��%�l6`�ˉ�L�M!<w�b�kq�r�� �d�(�.]][��{̥�GS�ja��~�w����Q\�C.ۗM%��
h�s��F��;�¥FI(�]6*�C��}q1���V&CI �m��	rK�N7�0��D�zӀ7᧌�k�eES$���bi�V��$����)��|�3q�QjI���Q��G3�?\W-�9�����P%	�"&,��q����C�[%I���v�I#f؅�Pᩑ!������ }b��(d:�p$��v�ˁ�Oc�P��`5�M3D��wލU=1�Q���TB�����怉t�]���Ҧf�&�0�Q�5�0j妒���o�q֝1ѳǪ±ZmU����܍��y���*�5M�Ӕ��2�1���f��ټ��1a��X���ϑ��S�0jB�Yc2�Md��Z͗M���j<L�z9�i�3�Ew5EJ����i�D�c	��Q�ݐ$xL^Q@^�mI�I$.���������|'1�����;V��j�>UWV{�ʷ�`0��a�3ة��sz��]#Fi�a)J/"�%D'k��փBT�Qaa���Pq��̹\��Y��^G%��~�^9d�����d�>M�rm���h%�Y�o�)�%����ra��#VI�,�NNGC��m�y?}m�<ióo�M
*�����?֑U@Q�-n���k�ݵX�\����Q�����b�(��Q-���
�,���)$AS�D��h�n�B!Q�*q<M��k8�(�B!�Yvm�4�&���bScN�~_�`�+
�#f)�ӴS�6�%�ÞK%%6�bp���SfT�|��[{��F�_l�̓�8&��g�w���\���Gqñ������Ӗ��-��]왖�{�m*��0M��E\5�*a�H�:�u4�f)X���e��o�-� M�͛8�+��Zv��_^���Y�Q*�I4	��<��ɴ��|']u�0�4�:�)�,�
��Y7ݸ�&�j��aN���0�`��kN���T:�]2��[���N'@�\�̥�� \"x4�:�K�w�<`�
%C��:vj��l*����N������آX��DlD��(6(؈أ,Q>l�6U�K*YEX��U�c��,�V%�F�(�<6=C��Q,S%X%�6(�΍�Á,DK|P��O8>0W��r?á>ώ���	g��<6'D��TlR�A�(أc�,e�K*ƗC��,P���G!G+P'�P+��B�'�T�j9
94'ɋ�	��\.��elrYFF̕���P�6(��c�lrY���譎K+#c��-6������滏|U��s���{]��y�������'{|���z�Ր�ވ�)x�\L=�����jdySW���5�p��5���:~�������)��[�U�w���>���������w>���������w>���������w7�wwuUe���o�����UYw|�����|�+��Z|��#��8��[�I��#��e�
�F��i��]"i('����:ʘ�/۵�ZUc�^�f�6V���"݅`̙�wĿ��U�T����@QǱ�6��q�Mu��U�$L�QTUST7 t�<�bh;i�C���#|�0h�ⰬV�Ui�Y���y���J0	��M̙��B��1�1I�؋�7*J&V3Ča�uX�W(��Ʉ�Re4٨�,�:�1��Nt�E���[�O�ORb��2I!�0e4��7�L!M��!��<���9�̛��/��sQ���O���a���g���U
/(�k�����-���F���[Ӛӡ�E��;�Z�["��J5�*.��&�J4�-dsE�v��M�k&lxJ��ն�\��M�)������Y�u�7e`ӎ4W[E��yr�,n���@�+>Kn��Mmj�Ș��"��h-c"��E�^�Wj<�\�54zr���1J�vh}�ڢBF�C�Բa�\��9J.9H�R\3���+,:��|��mɏ;��߱;ڵe�_~��� �K�L�:�@6���I^N�`�C+�������i�0Q��b��*��d0��g����2���Z�i�N4���Ұ�V�V���;_��T�&��$:%���3�%>L)�ɰ*2ɴ kA��x���*������jbz��t���`J�S�0"#�h�t���&�I�a:)�`i���0؛N!�I��g�+
�~mZq�1�}�4�L�a,rL�L��P�c'%�g!���2texYUGN�͠{:�����V����H7j(�+�v�y ���|gTH5YGI����r�C�>�����Ys�nF�/�P�=�!:�ǣ�|� ���v٣o�±_i�������@�^͊4�mZT���l�.�ld�>�񸲌���jŹr��U/�J�B�n�4�;����۰.�!I>b\8��M�)<a���3Lۦ�����w6�6��P�,�7�Cb�I%'�!�l&�C�M��?4vv�XV+�m8�?����E��[Уۄ��)V���"m6���O���`@�c���S$�;-�PBv֘���]��+P��l�(�R+T�ncՔ��Ħ/+��BH���s4>0�K<	����kw`e6���MrI�������ɋ���q��:��Z��-(���&�B�!W�i37;��qcR=����Ԫl�Ұ�WF�~(��{}-����kZ���C��&�&�@i�G{ O9h��	��U���P8L>n��̂[ �&�2���i-g=�G-��2���+*W���J�p\;�8\>�@�����l��F`ʅ�=¬J���oS,zن�+
�tco����d!Pa{�.�E�y$���"���M����2�;uUEy40�L�	q=f�� m2xb5�B15$JI#BdN�#1���8�.t���ᘟM�@a.�i<�o �e���8����N�I!,�����ψّ�'��c���aX�����Q�����e?�2��œ.egdc�#�����☮b�?l��#CR�c��]�K�S/F�e��awh㌥I%ޚF��T��1�U*S
:���Q�M���e�c��j�l�H�K�B�3�)�Y��(�eV7>r8������������W�X��Q��|"'��#�G��F|*�*6p�EҖQV&�#cbd�6Qfi���S,��8].���F���lQ�<R?�2�U���(�	��~�K�S��Q�E��<'���t�أ�6(أb`lK%�c���V6p�Vʳ�Z����4��ǃgJ����<U��l|Y^:W�t�[�VD����+T6�,��%ptp�����[�VF�xZ��F�,ʭ���]��FӖVn;�Whu��=j��9�~��3M���>���4����������n��������B������I$��ۇ6�zȗ0���t)��.�%�}�.���%�۷�&r��۪j�$�AeBcG�g�4
�r�nȣ~�5���
��5�wo�0]���>r��7�|����>-F5�/ST�闲pOSb�����Rυ��Ύ�x��|.r<��T���e����Z��8��]۲D',���ⓎE����ϥ�S$�w���u�VDږ^W�=��ێ���kFc>��N)�nUz���qґ��؜۔��4[�'�hꃋ�֏53�w�����lb��6i�U*���\��P�U��-WX٢M:إm�D�nW��A
J���۷m���b&�U�4
���'Ib�ʔ���j��bچ7��%e	THL�GJ�kCB���icn��n�i����6�#�AFF�M��Z��لF.ĭT/��&��QN1:�J���s|��wwUUe�.��[��˾]�����UU�|���o�����.�w7��wwuUV]��\�,J�,(�E	G�������E ��D��4�a"y���O%�mB�B�R��1��7H�=�kQ;L�a�p���x��EN�D����Ț0�u,G+lF�v�l�V)��:�KJ�-bZ����K��iIF����$�.,L�lS{r�Nh�0Q�!g	�ɯu�L��1������2�ɘ2�]�R-%%!D��9I�o���q|�!�d�E�ng���+��1X���y���W�ʦ��vN4a�O��ۤ����l!��i��C��y�'�� y9O�%&:B�ӦI�p�1@Xq '��)�5�FH#>�XU�e}�a))�*S�i�@,���v�MdȗJC)N��p¥ʛ���w6%ýj�!�śS�a�W�8�co�ve�Q�L;f�6@�����5��9��6`b);�ԔB�ˤ��Ô�n.��~^ E��ǟH�㤪H�+�SJ)��*.��2OA�K��EQK���$;�і����ɽn�$-GS�eMܦe�q�U�{c�����h�l1���Θ�:>Y�T�	{6�G�q���\&ܦ�i8@�qj�����3k�嬶5$V��jܕ��U$jXےD�1~��[��5���s0�mb�x̨>���Y��ݩ�1��q���/���aɀ�͓�<��b�5Frwa�h�;UHS��\/�"��m�^�i,�1;�����b�;x���z醾\��D�]�=�6��)����3W�	'k��M��h�'%%��{וsF3�%��7\�U�hnrR�TT���_$��k6���kUKرk�)9���	�M�[���p���%@�^�櫵TJ�)d���K�ru.-��m�����i.-Af�F�M�L�.����!\�Ž@
%���#���#M9(\Q����L�l4�FE�1<v���c�i��L1��U�+�7����!�(��>�j}�n e.�L��)�C-I+a|�;6�4��d.�9�Hi<��e�.ۺ��ת6&��
���3��
��2�Z6Ot���7�����i�yrg�!ueQ)�Ź�
�8�#�Ι�ͧ���c�V<Ut�uk�J���] vn�M{'g!���@��f\�f��P̤��RR��t"y)��'R���sz��{�֫J�_5�b�\o���.��fX�q;A��V��t酷���Rɠ�~,x*��ǑXM�)�e8��q�Xц1]*�ګ�7��j�4�,a.;{�M�̉���f�m-���l����7Z�B�U#M� �rW&c�����C&��zۆÀ)�&��p���X<e8�<��&�w���%��B14�ci��v%�ż�F�Y�z�-��N�*l��
(N�lD�֚ٗ�X�4.tcW�P)�xY���+p::���n�\���cj�[ǯblE-Bam\��h�	jW�llT��+C��7ci<�qD������N��-_�K��+����Qk���`�0���R�S�)I��9�]�ʵ\:�����xκZHY/�ۄ�e��H�)6��K��{I����T�!ͦ�-i����ޓ�J��(��&�`� #M<��$�>�15<��K�cɨ�ꦏ^��+�	��	�.coW��D��f-(�b��Z@�9{c"`5I�8�6�p�\�'�5�Τ��K�L��n��	��Pd�)�9�>���0���b��8��&��O����[�5�m��;K���JN��x��჈��k?#�0�U�+C��%|2�G�'J<"&��3W�
%�3�U�F��EX�(�C�,lMT��YE�c��(�S�c���Q�F�E���6!�D���E_
=�ѡ�x?���M�|<��O���<'���t�أ�F��c,MQ�ʱ�el�[8W���Y�|9:WS��Y�)gJ��l�<`ŏ��<Y^<WS���.K+"X�o�,�llQ���[8W���t�K2a�j�)�M��~*���G&����9=����p�ý�gA�2����������]���xx�"��^�2+�㝇6-ٜ٧9Ŧs�FU*t�󬃰^��lΗ�uM�S�d��w����ݘK��βj�};v
���U��ٙ�U�)~�:���.�w7��wwuUUe��o����ꪪ����S]���UU�˹�����UUY|���]���ֵ�n˵΄,�����?)�:NI�*��||_I*��,��ɔ�Y�a��Ih��I	�����1�σd�����l��u(��EUZ�r:ҪQQN����<�����ɷ)�ki��ٙU%K�4������4`3�t��f����a*뇉��%�>0ђ��`�AE	��F�c��H��1��3��J� �����">M�w��q;����?����+ J�Lv���S�����	��.g��b]ɉՊ4Y.5J��Ǔ���!�2�\��a\�I;$jS�˅�krƧ"��s��q���Ҩ���$�B����FO�#�7���#�Gt��f�Tن��%����;��`�Wh���*�|���z<EETo+��.R��U�Ũ�z�RH�7k��R�l�ղ��C	ͭʍ���Ur�j����a�� �YÄ�a�G�$��+xM�w�-5Mk�K��f�P�,4M_��UD�Cm9�hK���Z��6+H�Y ��V�0�1s�s+�;�b���2��ʱ��Ǝ�a�W��|��z�{�]�3OC���S��`�}����p�j��B���<K��%�)���UB��Ap��K�6��R��QԳ�'��S4�g�⸑��'�;e��4��+[Ol��C/�<��lL�v�.4��J4�P�+�ϋ&ϋ(O��Bk�B�v�6�F1֩��SS@}Ha�XM���J)<�8��dQ^J��g��+UFx̲^�˥bH��'��ĭX��	�:�v��֩�Z��h,�J\�8��c#�~�6��9j�Q�����+�x��j��y}������.�"a�AE�OK��L%���7֩#��KA�SR:@F-��Y,JM&}�	��W	$1*����xsČ�q�K02���=l�[���P�krK�޼���l�ڏ�Wq��R�Wʬx��������N�gT%���;c���5Ӎ�U�*riTݲ
G�rn�6���"���+4Bݼ�ȇ�e�*�F�UEB���y$��n6�ޖʕr9�!Ll�=*��)(bQP�������k7O6.��m(�bZ���7M;w��1��?7j��Ӥ�C�>(>���}j)�\���h��	�,�Y�����iPQL5MRL��N2�`f����r�ij��Q�(2 �b%1�h����ɕ��{�#�����l����K��I���7��έ+CgB���x�/A���`U1�������}�xj=���r�Lir��Ѥ�Hpщ!`��O27K��%���ަ椯lҕ�t�Ǌ�����˛�[[;����s��K'3�ngcu��i���5��]��H��킘�_�s7�����_�UP�L	�`��ɵV�f�N-�c,[4�}ܪ��*�dy<��Slt���+�qU�ʯ���Cc��#�QZ�o�%�!�]I}�����!/<3���r3���4��"G���rI$r+�%��
z�9�������=|yI�6�B�FmǑ"o:�jT�QE&�����m!���5��Y0v�>��,��xk���~��G¯rڼYU�՜+��3�W���|	���*�B6'��S⌎F���e'(������	�����e�(آX�ʱV��3��O�¯��(��|9���>(�z|T�O�ϊ��N�Ģ�Q�G���6"�T�E9,�-�1c��|t��K*�X�rt�+cg)�Vt�i���V9=M����x��eY�\�VF�^�E�F��F�8<0V��ô�7K��2680U�i,�l^=���N�}.�b	����X�b�V�'�W.��4ږ+h�:m���~����'��j��W�}t��a�$��*�� ��*{^��ܑ{~�����58��go_ڬ������G����u���g�����z�
�;NGo��9�i��/{s�6�/c�Y(�֩�X�$|���r�#�f�89{�W�8k��y���˵ݒo�i���k9�2D�[b�$mv�*M¦����}ص|��O۷��\~����z.uu��wb5��8.j�B&�kE]�a�Dq�#��)�t���)nY Z�m:�.�¶<�U��(�Rl�p����"�#"$oEt%���S�L�QʚV��&�[�1j��a�Y(�D�A�;SQ�Tf�\���M-6��J65M�:���d��B�[6摧b��w܈M�|�
$Ȥ|{,Qj�F4�'lhM�R�6GZ'�E��UUY|�nywwwUUV_.��wwuUUVr�oܻ��ff{9w73˻��fg2˵ŗww��9�Yv�2��%�b���!��CÅ��m�ږ�V���6���E|��X=�����!F*�njf�ф��V�Š��Șؘ�>&��"*n|�QQ!M$Z��q*:�J)���Mo�.}t�U%c>Z�1�{x����GRiw6� �[R�cF��5y�V�p��� �bZ�b��b�5�q�8�'"�nF�QX0`�c��(�0v!����ٵ+�Uc�W:�_1���k�����QU�{�kUH%R�v�(M�� [����-!8��Y���&͖�{f�c.��DޯQH�a���CqL�1L�D��s�
��O��K��vH�XiX�œ���G�W��U�^���G`,Qx� [)���L����c�5n%�*�T��8��E�8�G�����Ecɸn\����z��*1¡�cƚ���<��ۄ�	T\=��c�(rB '��D��&f\�kh�Q��R��z���:,�<�L��=�Hv��*��b��LRD8�������IP�}���t��e�)R�G{T\LA9�Q�l�Y�PK�P���,�_�ʮ`)�ɲHB�Z��M4��[�KS�o��}8ζ�j���:��-vY�ii"15���R't��@�Ńr���#�mHZ`a=�����$�ց�\���)�Q%���"�Y�ܱ��VI]�T̊�rUELx�-jb(�p���ĨT5�0�d�"��b�)P�Q�&&yIW�*��(���m(��@�Φ���m��#�X�q��c���qv�����;�:i>UqJ�OX��(�T�x2זЖ&Eˆ�	r�[��l>#�bi��Ÿ��HQ�����.�+)��t�wd����
2�s.�m
<W�Ԧ�6�i�l����{1<Os�*��g+%a54�%\��w����/��S^M4�C��W�r�r-��>�8`ڽ��n3���*�昭�1Ō��i�nc�}<�k1�+M0vK� nn�����e�	��V����;ҡ'R&��!}��IN�']%���d��9%��j,kq�y��i��a]����w��XM�P�7|w�4����>��:O�M�՚J*�Q�"Ʀ!��F�%����k�Z�D���ʏ1UCT*K<!�	Æl�%[�K&S=���lY;��U%2��R�,��Q��L�7��V�ei�qO��d���bw�kZ��ֵ*r���M����rD]�UN�8��I5I^J���M<�=�h��5Ș�YQS��H�SR�acMX�5m�Pc�VE
X�����7L���(�i1)3X�29���wj�\8h��$���j�%�(����~���.3�]<�[Q$��g�X�kHU��<���IE�V�S��5 L��<�?e��Wd �c%�(� 	�q�+i�}�%i��Uv»S�(��挲�a�	H#�Jy��pkL�P���4o�䠭��U&B1�-މ�)����I�;N���sK�Vj��!C�!�V����C&!�t�-QG��`�=��*=S���zǮ?>t�������+�8q�q�㍸�/c�/�8�\8p��j�������8pK,�e�,�g,l��>4l�"rBR����(^B,B�-X�b�
�^R�!Z�!j�j�B��N�tӍ8�p�÷۶�����N:iƜb�q�p�s=����(��ov�8X���^J�ݷ��5�z~��U�z.������>�+.bg��2��Α3<��U�%v\��a���o��u/V�lT���Dn�ޮO��-�i��`��.˳Hgw�8#}յ����w���u�
�~6&��wY�`����p��e�`�ln���~��=�[��B#��u�Z�����+�6ff�]��.���]���wwL��g.��˻��fg��s~�}�z�s��k����Y�sw��ѐ�,�K��(�����	�:q���4kip&'���n�bT�n�Qd���1
����ڋ���~^��ޡSs'au�TLL7r��硨j5�y��q|`��-�f�ٷV8٥W�a��U�=c��r������W�Q���(�Q�;3.1��~�>/�.��l{V�5DƋ�S5Q\���vgP�^�y�F������XJ�q���G�(�z�K���P��ޔPr�b�Þm�vt��c�Utǌc6�XI��r�Q�j��P]ұ��c�RW��(W��Hڶv��lf>4�d�#��k$N�m5T��4LMC���&��y,�pjI&�R䕩`㴵Vۉ��Em$ًqRjA3r*�������l�3�7sS;
��"� ��;�`İ�Z�ó�a�Z#�c����3��!�kn2B�-LlB��Y���K�f�|\5P���
,DM�x��/�k�W�Fs�2UXJ���9�&�3�Q�,���kȴ����}�i)�к۵�e@�dʭ$|��|��,Z�_�QI%��x����#V�^1~�B���h�>�;�Vd�.��f��
Ұ��UtǬcɬ��W�� �&S	u4���`�p{��'Qa�2`�5�C�ɬ�?[%���r������$b�&-m1C����|����uxF'��Qe��;:06K�2ySԊ?L��ۨ�+�a��U���m�JMt�IM��I�N�'*�(�� �X��v��'���!�_��c����:�0xNl۴�b�r�eI��Z^��gqZ,~�Xp���.!Z��M4�F�r�K7m\�^5^��f���u���Wu�U긡�ƛ(�I[c� ��E5�
��
�u;�un����E��b�4�QZ����4��7����M�z��I%�^��2����CJ���>����B��������2x�1+Y�N�i	�Ӥ�gk�46���Ed��*��y"�Z-�fg��n~���1��=a��lDN�YE{K�,�d�K$��	sm8�wX�
�D=H[E,��M�ײ}�]ǝ^�_;��g��H�!K("H��g�ί|�߱n)��ÂNÜUK9P���T%*�Y�N�Xa��U�;c=��7t׹��& l䖪���ܻ�sMF(x��Lʞa�zz}��ţ1U0%�T�*L���K��,�l"S�e,瘒HC'��apK�C�J�x�hi��U]1�ƣw_��ذa�f2sʪo&��\4�u��0���!�VUe�8Ҙ���P3�8���j�%W�Ly.�3I��q2%�
�ֵb8�c"nD��q���8�Rc����4>,J�d�E�,�:<=6zzzc��8q�tᡱJ��B�jh^M4$$$$g���Y���,��d��8|����;|��>>4p����M��-X���B�B�K�P�+B��q�\z�<v�q�i�+�8��ݶ�ǎ�:q�N4�ĢQ*I��O��M�)H�]:��t%c�&1Wlm_,<9}�|�.i����ƹ��j�8c^9�>F�\����ꠟ��4��k}���qs_�w��GU|�&�/�UrZ��������,��N�c�!�K�mƍzƋ��<�syE෗n��ը�]�ro�l����F���%�U�Z�	��u��G�Y�{~�����s�/��'m�j��ȶ5����5V�id��]VB@�����yY��;�ǩ����.��Z�xO��m/��Eï���v��imȯ�n�kdU�Z�G�J�(ۂ�ٲ�]4vv�˄�77Z�w�_�xɧMQ�r��n^��g9����J_�r+�uE����:�؋,C�M�N�mPA�����ϯ(�`<�X+ µ-�*XH!ܵF�`�R�vA�kP�Tyrڢ�(`�lr��TB���]C(��kWGk#�j�%�r�I&Z��h�آy͜��kÚ���OA��بGb#���4��ʷP���P��%���~����?x��߻�wuL��k�o�ϻ��f{��7����S3=����s���}����wT��_[�FB��

,DK(��(�.^�/�R7���\#�LTL�%�25*��7F���Z�F)�('+r;�2X�r��KbN���؄	ĝ����K&sR9��e��bض�*1ki�L�//BK���;�a.��-�ϭn�h	YN�5*�t�D���N��J�+�zn�0�UT����J�.�SS��|�IiZ1ʭ��i=9fz������;�G0�*��F�(���Ld�Ԕ�i1o-D&��Y)(<р1cQ��QF��P�3�}>�Q7��?L_ؽ�����##R�U*��U*���Hd�oń�R�cdp�7��c��u���Ӷc�Uz��4�KH1��)8�7�������7,0�JM-�:��u�$��z�ָ��TCrZ��"y�1a��9P�f!Ϯ��;�[��o�TJz�L12�ɼl.�Ȇq�NU�UTҵ��j:�V�{yߍa�Z�!jkɦ�jqJ���Y�)��&/��X�L[ŵ��ծ(=��V�r�U�Wz�x���ǆL'l�5�e��r���gq�ۻ7����*LyQsy�y1
C�k���̻��)��1�UxǬM4%ؙH'�B�N����|d�(� MN�+7i�c��i�A�[���^�V���?H��는�IH� �1���H��eV9m����,TT�(��x	�D��UI,�M'��ɮ%λJ����d�h���M�QZ��&����>v��l�wh�t�S�0�N�rr�Kh5Q�,�Է]F��?-�r��\�c�f�Xa��U�8�1o����Y��m��/�GJ)�]�̸YK���yc,6��b�<ʪ���m6�M��&ڤq>/��	��H�L8-kH�N'��L�e�}Y�E�ig#�a�:Qe(��]��R�R�p#L�R���Q��&M��پ�z�k��zMbp)u�Ta����E�H��7;
�}Z�'�aszȩ.��Q��t���Ǵ�w����0e8��)��1�c�1��ԑ^@���&�z�9T@2g���1�$r<c��7$�4����us7���X����ʬ��x�6V�JD�I�t��n���z�:�jJ����O'�����W����AAGH"h��(��ޛS��)������$�<j 7��x�ZY�ʨ4�M��e�x7.�M�Z��j5d���B.6��
F!�X�[<V%qQ1�,�7�4�Jj5�c���51G��DO���Es1�
��I��tn0#��(��(���k��UQ�~�����T�DW��^N����N5���kS������(��[:�yX�A�_�+���*��]��M6�j�ǌ6f�9�s>�ܻ�����Oa�aԖ�58�ŗm��_�Q�!I���}�S��1UB6z*J��x�n��F&�UY��.���Ü
��ӷn=qڽ<=6zzzzҾ>8ڸq�m�\^7��q�i\1Ç8���:Qe���66Y��<p�e����ϕ�8��N;qӷ�B�K�P�+B�(B�-B�!z�ێ�tӍ8�Lp�ÇӦ��j֥HT���(M			l)R���ڮ�4^pSM��oM=�>�q.�e��7.#���]��T;��j�zdb�O��蹕�7�z�1Z��#Յ���N�_'�'��:s�F�+M����ų*#�*�]Ub��\R�K���cǏ&c�Ђ�w���z{ޖ����������2*�FS��Sn��b�j�g��r�wtwuT��=�]����˽����S3�������꩙�oytwtwuT������a�8��1�1��-2�����`�]��p�1��g)p�+\�����&�m&��$%jѸDc2a�����b�{�������<K�m{xH`�q���"[[��U*QI��`e6�2�4=���a�*��?1�qſU�h����MCS3N���;ʹR �p�UG�C$�	�m�jY@ʜP�#�!ɨb�*��>�!����8���Is^�ۓw�!9MIY,&�	.�<��{yj�M�h�!�7�Fa�;UWlx�0���Z�h��k��Uƶ��tkMm�&-Z詺;]�,vl���\#�%i�8�$kw V��N��t�m̊5b1��P(�H�EUN/%����:Ӊ6
<���En�g��95�r6�,nj1�_ƻ�$i={.�\�HOv�(ll��a-���@����oU��p失��핪��z�WZ{5T�����ɳ��I�$LQӱɒ�X�h6�t��X�cO��5��='nM�,Y��N��{R6,�UmZ�(�A`�ě��fO�vx�����7���y���~^��nIkAm�\j���Ё���n\\K�c_�ã
*v�ϓax�J=ú�;j�X�1�Ut�Lc'9f�5�P�����+!�n=K�܍�]�]-���x��"m@C���bD���zYp�3n
��Wa�t��Li\�ы�mu��<=�j�b��a�>��0��U�1�Q=��#lR(,�E�9���Z��qn'���{����2H0�eU^�Tr�4].�.�M�I���1�E����W0�:^�!p�p4�����x�J�D�t��j�a�6��X��w�O��̸���M�R�ymL���nZܠȨV�$#�q�Ur��n���++@H���e�c��XƝD�i��Xޢ�ǃ�x�.��"�nP��0J�l�������b�UQp�!�W{�_C	"Re�%B�c1��I�����'|���b�k��۶�̎��e+V����孤��Oy�q=��	���a�*��;c��m���n��oL��VKN�o�z�zO"�m��w�J�93ݪ���&w��z��(��I�D��7�U�1�����&��UW8�<�)2���mP�E�9N����¡���cE�u�p4Q�8��X�c�L��q�#�:�4���%��+��njY��l`óp��ڼ0a�4����a�����J�>�UrU���,�85��ܖ|�(�e1�D��h�)v�P��N�2�I;�擳a�*�lz�1n���`�NcC��\4f�ú��]�!�_�{ص{<�t���\��+S*��KUT�V��J���$0�υ�!�C�h�;��"��CSPr*���˴�a0z��:���I�i��A���>�R"��UUXFI$!E�~��п�l���$����lX�����1J+D�08�����f�f[
Ŋ�VR��{A�JE���JE�R)%"���IH�)�����D�T�Ia%�%"��(�%B�
,���EHQdE!EJ��ȔT�)
*
4�b
*B�"�"QbEDQdE$QdEF��jIRE�$QBQ`QAE�QbE$XeH�%$Q`QbXE�$��apY�2(�#��(�E����-��E�X��,Qh�E�Ń*FQR�E�,����.�j����?嶤в�E������V2�W��*�u#%QeQh�B�b�:��F�Qb�(�,��,QR�R2�YE�YE�,��(�#"�Qb�E�Qb�E�1H�EYR�KEQJ(�I,QR�YE�,�y-�бEJ(�E�X��BȢ�YE�YEE!e(��QB�,QeRK(�E�X��(��YE��DbQb�YE�,Qe(����,QeQe(�(�E�Ie(��YE(���,��$�E�(�e(��EJ,RK(�E�YE�X��,QeRK(�E�X��,�eK,�b�¥�,T����T��,��(��(��YE�,��RKYE,��,��,��Ie(��E�-(YE�e�QR�X��,Qe(����,��EX��QU*$`��B0H�#0H�#,T��YR�K,R�(���K�D�K"�)e,R��K(��e,��X���R�X��K���K)J,R��,��X��YK���YD�K)iib�)JYKKK)e,R���YK��I,R�h���J�K)T������R�D��E��*�)e�*�)b�JX�R�,��Q,R�U,��J��X��Y(�R���JX��Y(�K%�X�)e,��K�R�*�b��K�X��U,R��E%,R�,��J��Y(�(��JU,R�,��K�T�J��X���%,RJQh�J��U,Q,R�,��D`��$�`�D`��2#d@���*�Kd���X�UEY*�X�%X��*�XR���VJ�V*E��J�Ub�U��*E��J�Ud�Ub�j�U��LI)	H���dE"�)BT,����Ĕ�$(�$�E�%"�)H��H�PR(JE�E"ɺH�)"��)IH��I)$�TE"��T$���/X�?�E��W����)Bd�9���}*(��$����$�b>���O�������o_.�G��'��.� }e�����ϟY����[��u��X����_�r6O�������|O����$>Co���}E��?���u>�)>���y��G�EU������������������@���*���%$#h�?��?�\�����~��$2�X�)K� ��6�x/C�p���B���|�~D�?���$�	����?$����C��H�4,������1>�e���RR~���������nM@�	�'��s6�\�V\%�X����o��䍲ST ��B�Q[�D@�C"D�����	'�7@dDK�~uYi��V��jm����\��>_����7�Ц�J*������(��@D@!����~0�~���v��?�~d��h�� 8���l��P��?���L�?�A�*���k@j�e���͟��q����.����_�h.�pV�~����� }����������D�g�!� �ꯓ����?Q��X��*��P��	�_���C�x�V�i������C�e`!��K��? ��'��ެW쟟?����X�`�?Y_!�h�p���AJ0'��
��_9!	��ۓ�,��XH�))`��>cdL#�(c����)(�����L��ì��؍�\���.�M�؟�;  �Ϭ�'���Q�gֆ~�*�����H���~�O��C��?���G�N$�4�5��1�O�~��ZO��?����ڐS��C������G���tUTO�H�|PB���އ�"���~��ϳG���?���/��'����R��ܯ�*�$`RB�������\�b��Ώ�ھ���E�����O�Bۺ`K�)��ݴ�7�~��TL��'�~C����D�'�� ?!�� _���?1�?���v�S{H��!Z�q���?�~tا����>I�PP
b��ߤZ삟@�?ӑ�|ρ�A@>a�K�@����R����I���\������C�%P��;�M���rE8P��[�_