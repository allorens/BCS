BZh91AY&SYû��H_�@qc����� ?���bR�         7���=��M��J$ ��V����
h6̨R	B�hA��"@M�RTP����@�m��Q�R��
_w�)��6�5C3
��$���@��Y�kj�U%$�SM)����iV��RV�me�S-��نƉK$�M4m�f*�g�c&ڨ{ޯYm�Dʶ������S(i����4J�V�&��R���(�+ZkEA���
��45J�hE�he����V٪���ڭb�{��5��Q�Ǣ�    �z��J�� utb�C@[�C������6���C�M5�n���:�AВ�Ջ�jf�����T�D�INa�U�&�#X���   ��_J��U��ܸ��ݻ{;+��T�S�Ξ��zңe�z�w�MJ�*��z�������D�U/fJ%��{ޚk;wq�z=����fR����G�J����}���iZ�ZV[i��   ���۫�����{-�iPR���ޖ��K]���띵GZx;�}���hK��}TUW�$=��Ϗ���jGm9�Ͼ�Q��2�'�{�)(U���|>�U��=�	�Q�liT�6�5�kJ��  �ϟJ|�KR��>{��2��z������T�}+��_U�km��}O�zR��^�A�����}Z*�Ϟ|��ɪD�=���E*=m���������ԩ+�z>{��֬F�}��CT�Z���ƳK-�l�|  ݜ�O��QJ�r}��}�KV��������٧�����K���ٸu�)�3�wl�כ����R�Y��}��>��ۮ�;����O�$�t���y{������|����%��W[f֤��Ye�[&��ѯ�  ;7��W�o��k�T�ʧ���ޯ���W����x�N�{�>��_m��t���f-���n�|��ٶ��F��c��ڲ�ջѾ���]-_o{���%��Z�/���e2�ֶ�f��D�4�|  uξ=�mRWu�����NZ�w���χY*S�Q���>��i��]}����m��kG�=�T������\PO.{���>�
���Ύ�
�*�4�H�Z�HSkj��  ;<�4�Ek���������� ^�9�[�A@�{ٹ�=n�9� *.����>� }���AG�^���Q]8׸i�n��yR5�٬!5�SJ�|   ;�{��P��WG��n��z6`���c��+�zn<�F��G:U�pAO�ި��z��=:k�އH����*��4�f��-��mj��  g���|��J(k��n�ҫ�kx���J9�d�T�nO\��(3ҽ�@j�n��PP�^�/j�1�� |   P   ��2�*��z=@��������!���)JJ��i��ML�dhb'���H      ���J��  `  #������T��0�j1Q��HM"J5'��OQ��3H�O���}�������9��z��0�2��t���X�7&�R\u�!H��S�>�|�����BD�$?P�		'��?���		'�����y$�'�������O��!FΪ�������`�@HI7������`���I����O�?�IчD�	��td蓢D:$蓢Ftd蓣�'FN��:$؁сс�'D�tI��(���FN�:0:0: t`td�����!ф���������ћtHtHx2t@ؐ��t`td����D0C�D�FD�FC���D���!с��N��:2`�FD��:080:0:$���: t`x$:2����: td�����!ђtHtM�:0:0:2N��FC�&td:$: td������@���td:2蓢B��E�N��'D'D'D��D�D
3�	�	с�!�!с����td�N����N�OD'D�aс�!�!сѐ��x0�`âD�D��D'�D���'FC�C�C���!�d��t@:2N����聃���'D�D�NN�`���N��:2t@蓢D��FC��FD'D�FA!�	�E!с�!сс����@:0:$:0:$:0:0:$:2N���!ф��:!:$�N�<N�%:$:$:04'F�td��d�x2<82H &@:0��N�	���F��$����tHHtH��$:2$�	!'FC��'F��HI�I� ��$�<���	҄��������C��$��!�!$����ѐ!с!ђ�$萄�萁��F�:0$:2H@:0�:0tdtHI� �!ф	�!	�		с!ѐ�с�!�!�F�BN�$:0�:2BHH��F�F�FHC�H���I��B�$�����	� 4!$����!ѐ��!�����I:0�:!tB��	� ��@��C� C�	'D`��H�ta td�!$�$��B`�@�N��DI8$�:! �D����؁��FM��lN�h@�ѓ�C��D�:!т$���ѓ�'D�:2td��	ј0��'FN��8 t@�ѓ�D63�D�	�:2:$:$�N�d�����N��D�)�� h@�������������FFD�:0:2t@�d����ѓ�'D��N�
 t@����D�:2tHt�Ht`t}�����<������o�ך&���ȷ�}�rM;qX�V����d�+(ѡ��%���$��,��?ݱص���� ����i��e<���m�	�Ζ)AA��mݗ�"έ�c*�(��YÆ�Y��eʜ:�%0`q��ؙ�;Kf�.��YcH�hA�S�钲*��,�6�g]@W�ŶI�c{`ZZ�����/i��ۻ��n6� �Zk�!0u�)F��j�e�Gw-뻡�j���mЭ�i�˥�����[�Pb�wd�ܔ�M�05�!�d5r��E���gVz4c�E�ݩ�4D�б%��7�ŵ2���ufnf<j��oc�m��Wy����:�JSN�Gi���tsFni�	sm
T�*V�yqn�u^�-������aŤ�\�`9�a�� ��X�,�`�Q�,�'�/jG��W��dd9R�ba�8�Fݼ!�,��6�74�!�������@�����R�9rneG�Ţ�эڱh-}��|�O�������T�֮��ָt��4[��75���qT�"�Vn:�{��~����W�����&�b?1���-��QZ�6ͮǍ�h���y����f�o$����=��E�
�#�2�*���w�Qu���A��n=�R�<�fҶ�'�X![e�j=�u�h�+)n�Y���Pn�T�����7x%�����=Z�&��m�֛���v9n�����z��5�t_�e]-�\�R�Y�[E���"�H��⳹�Z���0�Bmh�d�Z��b5�5Xkhe�F<2ջ	�� ��hL�0���,��x΂Z��]�SR��Z�6(^�o��+/qZgK�dZ\�k���A�F�U�����4��$��"�؆�6�^'n�BE�:b�.Mj� ��`��Bb�b���B7yQ9-��@У��	�.e��iLِ
vg���G��GĪ)�F�]��`�N�kX�-@��u��`�ۙ���
���"�WW�".6r6���lQ�#Z-��T�F٭M��0�)S�z��F��-���X�"��cO,�kh�X{�fa���U���s��w-&(zFvf*�u��iș �Ql�����3\�6��pf�Y�]Q�f�-=���73aE�C�{sI�v
�1�{��ܫ;n�jm��Ve���]="��TEA�S�[�X�,S���{ip �SoA�2���h�V�=�4�w���dy�;�
r� 5��(�$S{��v�j�Y�/R����F���9��r�V��)�v�dJQXi��0����Ѭ��7R`+N١4�fHּ�z2<�0��{gt]<%)y��̔�([s[5)�L���K'^�kc{�U�0)�YK1
��{��̐��<&���B;���#4�����Y���uwN+E���L�q���wr�^Фf��T���o��:��[�ba�wU5ؽY���n���xuf`R��.�Ǆ-nkb]�I^������yu�S�	��d�=tN1yN�Р��y{�1�2���,L#i���ݧܽ���2e-������ZX���Y.��?f(*�5=� �g]	��Z�u-3&��i%�n�	F�M�i�0�x7Zɞ/l���W2w��`��Vu�v7�WAY��dZ�ڒ��ӂ�M��)��������W����� ̐�.�H�9�l�v^Z7�ܩ@����ٴ��3I�#6acSq��Ӥ�+�6��-(fխ�0��MP��ݓ���n�4X5Ym卻�c)hw�#ˢx���)��su���wV�L�-!l<8�ݡB�������N Q.�lۭԍ��{��t�R(JЙ��9��/F�3P��z5�k���%<�/3�&`����C�h��)���5+�x"{ �*�\�s[�^w$3q�x���q�Z���#q��b�m-��=(;n^Gh���Oq�R²^^V	tԈ&h�y�V(��Nl��i��t�9͢�d��`s�nl!�r���uz��X(!�@^������C�e�X	B�n�m�+r��:.--R��R��kjzE�/6�2��:�t�t�P����e<���H���F��GSS�):��t(���3Fe�or��	�����/^5iH�ZE�: ���{��:���1��mE��fCy͂��Q�Y�q*����p��ɑ޷��M�#-\�/]^$�����B���� U!�bbiU�F�-�*���3�bf ����d)�V�v��ktgr1�����f;�J�Ƀ��2��ۀ�:
�,q@�W�kZ�քk�M��O���u���w�q�m�S���T�����,1y�#k+\���e�j[����m(��	�c�+A�!�UnRu(����h	ukw�J�ST*	�`�v�2��Qs[�X�D�9��n�[�[��m��P�7VXֶ���4�c���r�:��9ڑ��t�=�a(��!��!��$oY�NU��Ҷ�5��<�J$J�k�m�;@�8&��Bn�]'ccr�F�P%tij�Y���S�c#"�`�����s#��^�hڏ^���n坭����l-�f�6ޮj�.����]��GM̠�E�å,(�e��P�Z&Z!xm�ݛx2۰dEލ��OfitM���$�B��  \�09{yM 4hm�b���4+K��jE؊��w�K>l��4K0�T�Vfպ��=2��m�J�܊����uU,�����yUb֮W��%b9�ls��A�va+O+w#�@F�ء�ۭ��A�O�ٮ� �f�r��w#�ѿ�J�;%������:yQ���0��2�Ea�;n��(B���
[sp�奧̙bb��k0ц�Ax6�v#�yL�v���Qe6u��w�6�I�]����~.���f�o	�=V�b��څ����w�����y 3=Mm^+3n�k���	�4�7p��4qf-u6��+դ��S\�ʷI�e)�l<ڧc`��]��6�6��[=��@������հFQcae��H����M��f90K�!�!FH�a�ܑ�R)�v�byj�R�n9���r�/hH:�j&`Hd�8�Ɠ�a��n=8d�ݭ#5�"��K�l��6��S+FPA
R���]�E0N�2��m�i�p(�]��--�S�^�!�Lf]���:�Z6Ы{LKpf��pS��^VL��*��歐V�M�l0��E�[�W�4qLw�]'r�y��.âUdx֐wr���7'5�ܼ�-E�ŏ+E�1��iP�h�:˃JeU��ϊ����jFG�r�;��-g�� �'7L�p�����"�;m킕�K9��j��5�6��'�:���+&�֚�C��P�YwV�kKw�����&���T�:�{���x��ވ���ɔ$3Ȳ��r'b
��`+���,æV�4;����U��	l��-wngqv/�\���K�Ke!sYp`FKqf̰�UF^�Όv���[��4�\�jv���
"�!V*�����%n�Y�@ �֫7^f��T�6��MCC5�u�H6eC��QiԚ(��Q�W��`�&Cul�ǋ@u4��m�Opi���=Eo^�7��e��:h�\�`�f���#b�I���K,j�Y���\˽�m%mI����T��&6U
�W��su�D���,�[�C��@��%�3DɁ�����F�l����R�9��Q�nAcA���̸��N%ֆ�v�5���h��^�h�K(M�Γ�v�X�qm��'���;Y-����zfTn�:ehX����Lhi%�6�N�`qV1Gʳcو0N��3R=�L��m�Vv��`-֮�9x�1�
��u�s�蹓[V��Aq����T̦m<Ѫn¬]�dv�dz-Wvd(��ީ���X�T6ZaŔ�y��/�8%ea>Gh	�3%�@�u�R���j�/J&�tۨ�48�aKM�&�Jdt�Y۳�lѰX����q�̪��dJ��H�7$M�R�*� n��RԨ�ZHb����ֱ޴�V���Z��[���K.mY��vތa-�)L'J0��^aa�-��t�bi4�[Vs1i���˧���x���Q:�.�,S�n�sB�1*��a��d�Q���N��+�Fna9������[�[ԙ�fװNI��OK��l���[�*{0L��j��[�!dɡ*tżÎ0����I��Dj�aC���!�#�u��+Kk!�Ľ��v��'����X��v\���́�Q#Mdgp���f�r�&��Y�	R����ڊ�K���Owk%�EVz��h<y�������;�\٨֣Zv`ֳua��;)B"VP�t��]���aXw�=�6SXذd��Ep�n�.�!�9@�h�d�t۳F�Ī4��$i�ؠ%h��,��ܷ���Ͷ�2�d���E�'q�t�]�ǭ���UYB�h�𭦮(��h7�,ܭ�|y=GO��[:��w_ֱ�sUY���
MQ�����Bnjh�;!��,Y�U{���k'���l�u�=�BP3`{�U/m����,��	�wn�7Y���q�4乛�˼ږ���kM�r��q�z�и�!{�����Qvu����$��N����m�E���
�FU)�����p��e�ua��RU!A.����@���3t3p�^ZEnaйV�{���#E�ffa;�2�=wL!�R0cנ��kS2kz��V6��l��G�Ca-|3$���lt���B%��j򝂍���^##4D�VF,����2�-4�5���B֜�ӛ��cqF6�X�@YF*7�ƺ��C�Z%�[If��Bo��2���5m�����2��7�լ8�9�*xu��Xw����m�����D�g����q���tH�vv��H���F�z� 휛b@욎���&k��ucKŴtV�,co"{�F��`���^b7#v�")�pU�n6��V�T�gčM��"����ޜ�c�&�ĲQڳ zEh������%݋1�ó3eM�k'�,C1,	- g�7S^�a�&������Nj�Sh���36:
�h`DoS�Yc#e����=%6�P�˽(c9eZ�ݨv�5�U Ӷ"1�$��b�(���o^����a��mS�i�um��F`x��ݜN�:5z���˭%�kf�U�������R�26Z�D��˱�+ި@+-�F;�t�����Pf1w�SG0X�n6�B]�-���0৊e8E����ZI�R�f����7w��k,jۚ5�K��@�]CrI6��#�U�IF�l�c�IxV�o.�7�J@l�����̩�U�[-��ӳ7�l:ð�E�t�=6���e�M���!e&��:�k���|C��Ϲ3ˊ�5��(�9��v�Y��e�C�J�s+`{�Z�+ZԀ�TڱL\�WbYӖd�v�܈��0hz�̚��&�!&ތy��2��¡ݬ��G�����9U��e �g�&��;6�J�x�ݞ˴��7��^&�<�+,n�`gp¶�_�b�8���6��U��e��Y!,B�ǳ76����]0�˨���p��ziF�g�ݬ�F�v����6��6V�+-�	=RḺQ@�i7���K�Ǆ�d{
���K��i�o6��ٍ�wBE�]e���lT鷂+Khm�����56S� �f��ñ�&ѹ��r��W�K%���f��ObHB�ڃ�O"�an�JΚ,槯ƕ�0��/̢�2@6ԲFpM&��e��f����lm�RF�
yq&+	�!�6��a����<3pݡZo2�{���]�%z�Jr�5�u�io�s{w�km"c�¥U�sx���2�(��s\�L���AW���U��Y`嘬]�#в�ضp:��jUk�fa�O��4Pb�����!�D��5n�22��i+p v�V8v�z6*4�䬷�	����ic�M��۽ܙ����`�l̗�f#�1�3J��M]a��Cӑ�G]�m��r�P��Xc3E�lЉ�[5�GS�-8��֘k%�J�ըLveB-�QX)̤,�L'�x�[S��n,�̩%*ف<Ȳ\X�v�~�Ȭt��6��-���	�NO������(�Q�1�JE%[��g$�n�ѾOHY�EO3$1kgs�4X����f��«3]�e$-���Ė��2Gmn�0P.�DK�2���jS9E#!�{�R[�v��}��ļb6�׮�4����e=4sbYxU��;P��bg�H!��&K�����[[ݦ��ص��I{�����Z#ʗ��dT�����-�t'�g|�lv��<�of�6�����4
5��ZН^<���1��6��(�	V�ծ�b��
��I�Ό;-i�4v��E�Fk���5���Z×m�f�/Q���Ay�gXu)�<�#EI3&�
lRY����rE#�@<;����A� �x
�\v�X��4��9�{�%6(��{u0�,3�$/h�#'-:���.w��T
�i$�i�
Ƀ^��5�'�v��7eQ���Ux����B<�ә�Ӕ���	c	?�N7�)�C3N�ۥRЁi�~u��{w3KD�	FF,0>���dގ
�]�Y�O^\UdG+qc�[��6c���j��rϴ&Az�kT�=���I0���w0Ա��1��/�E&3ICSn��t�򨝸0����.���4d�	h� ��0j��5ts%�\Oma��B��+^RX;iɮ��V İl�j�kʢ�
�E4٠�Ĳ�f'G]Ck�#{���E�+�l^ͪ8C�FnNҷN�S�d�	f� ���� c ̺C1n�ئ������ܓfk�	g7D[(��d������tR�]K-x�MS�4�Bj%�t���ޑ�����������?Ϗ'��]�8os:��T뼊�,H��k��m���	�GY���c\������v�n��=H��&ڊ���b��Jb�����?�n��D�N��}2�ܶ��|�w~w�w�EfQ���Cq��YP��[�UT����o�d2�n��B�m�]��:�*Nژa���E[ƩK�@4D��U�o�j��K<���Yt�j�'HQ�}n%׍�^b�(j�+A�f�B'!F��:��Z�i�;;c��Y�٤4����U�9��Nen_>f���ؖ����3���Fj+��� ٗ3�P��y��9��]@\�՘��Y��˧v��*\(*�(�*��UH:�~��
��!���n�}Z,�{4%�[��i�{٢�іKC��@������q��ֺɔR�A� {�j5k(�cP"�t�N.�U��b�&��Щ��YiJkG�ܘ:]k SI�e�U���皺b������;�tv�hr���	�!4���� W��ݙd�h!�D�[}Ցp쳝滶������R�ܩQ
栬�󮱚���7�uf"���\�\x��|���'�T3�e�}�n�ӡ.�w�]��sD�D'��BL�U�'�{kn^�$ǖ�.Tf��!68{�#���e�����w%�ŝ([kR#�3�SӣINu�c-:���3 �����T��՚A����C��e*��x��pό_���}��e�c{o7��ˮ��ؐn)�;PM��W2�#�9g��ufz��^fg 	���%ї���?_5Aζ�誆<r��6w��,[;�2�[����-���経�;�S�_'���ݬ��H%�Ɛ��pA��X5z�7�9Q�3�$Ӫ-�t�p��W:o^Խ�8�]���+�%_A�jU#yoX�]9�R2��`;vWnE�%i��@��]���"��{|%X�e��ZҨ��B^!7r�YJ��������5��'=f�>n<�t[��+���	��Q�w�֎�Qr�eDԸc��a�q�õ�׌�,�E�F,��i:��R�0G��M�t�$��ur�V�]uu���?KVL��`T�M�J�qQ��X����YG�--c�Y�m)CK{9-��!W7�t;�z��JQd��vBvH/n�B��t(�ƺ4�438T��78U)���|6o"�R#���U�^r��0�� o�]��V:ܸ�A,��,9I^3C��uV����d�͉K�ؐ�ܧ��$ǵ?:�a�(�a�!]v$#;&�i�)�+�q�v_.f�r��D��ݖZ�Psr�2�s���oft�u�ăݐK��<�ݎ39��b��U�Lh]h9�$�4 R���p+�[ю�kD���H�m�%�炛�74�4�*�ѭ��t�خj���s�'u4���Y�L�%�-b(#ԡ�xQ{¯���\uoX�4�9F��Y���ѼaE�{n<���	�f�P��t�a�P�b�ϫ�F,k�@�nIκ���0�w��h�W���!�&�Km������Uq,
k�5.E���wz�h�a曆��:�A��SMo`x0oh�y��a�����u��i�R�Bt�r�^5��q\���G��_K֝��
QC��[��� ��Mx��p�7&�+O�,�ġ"�j�=�s�JgdZ������a�/RrE�.^U��-<�p �H/���S�3(��f��p�vN��Fw�ox)C�;�5���/�F�R�;��b�h�j��·O_)�Z�n�ˀ_��Y��;s1KQf�4�]����f�,i��d�}ѻ�J�}�j��Kʕ�(Kp��9\��bƱ��WZ�XwK�e���F��;&��H����I�[��	Lo�Qi��T�b7$�I��B_�c;��wM��A8Z`�\�u(�����u[d�m�o{24�'שr�S�4�Q��]����(=Kn����{��O5��D��z���s�17Q<�Em�c�|0�+s^��m�6͡,��
S�GsS�Y�t�Y��IA'oq��|'Ҥ�Ou�z���,f4(��d7��{p;�I,n�Q�3/:�j���⼮�/����N�Vf'�I��kXdz����k�ͱ����C��;�Ucm��-�\p�-��C��%yv��`�Y{&\�����eɢ֖N��S��
�K}�!�����_�}6J�j%��`�FD����%��7���Z�n���겣<��V��HSĻ�.�Y�|��,�$�X��Hn����7���uE�y���}:�K%��5��e�B3Xؘ�(�c���(��	Z�b�B�e4m��6Xm�qwcn^�:
��;z^��
�9v[|�[b���*"�i\Wm�N��Sf��B1�o͌�Z�Ow_`D��֦	T!�7��Y�2��ײ��n�
���ݐ�W&T�ӭ�)���^^\�A�n^�˷U&�IsH��!�\�kS�V`���j�X7�*MȦTLC*�+���㸮թr��7��3iN��L�4���(��\�c�|����U֥T`J�Y�qܻ�B��A�f'���6�B�)�Gm.����2_e��Ab��o;��g�ʛlI�Z*��fmІJ+^Kfc�R��q� W��ү�>hg^�ٯ���w��+{���v�xk;C��M\��P�r�n���&0)�2f�J��4�C���ү9֛by�.q8y �\NXu���Z�'+�4�f�F�sli��ʹ�����Zݒ���h���2nv�/z:��4��K�uZ�),���v6��3��{�}-��X��Ydo>��vv�"�[=.j���\j�����oz�j%[G����d�Z/��r��&2.+��m\k��0mnkD�����
2��u��{�{ �܌��Q��
Y\��t|v�����#ȱz/r��}����mZ@ٞ�ѣ�FM�')^�d"�k]����u��G�aj�Z�xUn�MZ�'Ov���L1P��k3�b�`H��R����͌���aTi��#S*���F���NvM̾��)i�l�R���X\�J�n��u�f[�Qj�y�Lk��J�wM���2�w�E�ڹ�� �g6����gGQ1h[��\�4"��<�#3kU�Y��0��U}F������ZYR�3Ei�(��ڴ��yu͙�F��r�3|��������WeG�R8p8[�V`�q}����\�^�|FV�j�&5����v'QWZ�.����K�/Ǝm*�ݧwls�+,��r��l�݊��M�q��yWL� �w����^-�ۛH;�Q�7�M�4H۬�d1J6�bV�}J�w�u�W�����3%����ʖ�N�4!b�;�G@�� �>�U�'lk����e.uU�s#F�$[��;��Cy�U�T�r�v\Y��^�/�ᇲ�z�����P�Yf1�����1[��*��L}��]cS(���XZ� �ɔ�'�k/��b5w�]k�{U�jH"�:�3;�=Yj���(�r�ޓ�S�c�9ð�ӻ%��ӕb�?*h��i���9P=v7!D���W�O�*�,�	�5$%iv(^u�M&�glȹb�Ѣ�p\4w��$��kh9�x��U9z�݄:lF�dB��]�2/�YW8n�q��]����@�MX�v��H�Nq L�;��$�Js7ֻ3����>k���t6h���7Y+�i��g1���%���kLFV��D��tv��r�h��7evn3c�R�L����{��`ͭ��qL&9�Y":pefD]\�:VCXlm}r�ĶѲ�W�E����S,g�N���oz����E�;Qr5�P�U]�&�%���w����btx-�&f�p�ν�MB�l*�	�]lGFb�G�<��\,\�ۭ�$z���*p����t����*k�T�zW���'�!�$���� ��z��znm1mLg7� "�)6!Ԟ�P��<�9��\G`�ǹa-��$9����з�e��R��An��I�.^m����IZFj,�Wq�o�f�2��L���;�QE	o_!���ɨ�{����@&D8XJ#�T9Z��74؊Ku������j��]7X����*���$X�-�	�{����h.�N�
���iRb�+Pc:mv��y�sbՅ�V\�s<30��Ktfl7�����8�1M%i��v�q�6��-֨�8�0UJ�kŷp8����/0�[Nf��^��e�]I�o+3([��e��ۯ)�'�j�ͼ�]ǁ;�4[���:	/]��Q�vv�v��DYѳ�2	�9�Z�wy!�ʏ#,$�qS&ޣe�v��Sb��W��-�܈�ɚ�EQ_N �vQ�D͉i�;���]0Xj���Т1[[}�B�J�ꉵW����޶�Rf�<���6�3:�jL���^u���5���-����Ýv���) 9HN����c��v(>P�(��;9АrgeY�j�ȇ�蓁CFD�W5#�y�m��j�Ӹ,KU�.K&�c�_,6�����{m��ne�(Ú�y<JV�2K�7ҵM��qH�5��y`��ݩR:���Q�A]gs�[�Ų�
��@թǊ�U�l4��Y3n	�3��8^d�]�!��L���d���^ʽۼO�� [rn�};F5�'��K��/Xu�-o��k\<�3���kf���B+4E��6#�h�P�نJ�f�
��{��1^A�O��;=�����ő��k}�R�XDN�rb+O	SB����z�!�@Źvswd��Oh�jX����-(SN\Ë6�H .���PB����(�2������n��n��<(�X��Z�z�L(a��ʤFS\����"�Kk��y��(�vH���-�`9����];D}�oH�7.��E�$\bmu趚�er5���'Mܢj�A�����|��t�S����/�D_,q��sSA-e�[*Y���G	�ʰ�1h�r����5��=��c6F_i�Y W4k�搗j{�Y��Ӫ����R�@~yk�ࡵսR�p�+���F�۷�EXdm;�2�!��'q�
�q�Rv�=J����<��8Y�����֮ɫۂ�*��JTj:�k�>���&��>�@�#qj�7��3�%V�d�!�O?VG��n�/p�n�-�LD����7�5��;ڏ���Eq�"7]}�t�廘�{�Uq��R7!�&Գ3&k
�#gݧo�S#��p����.�}z��o)0����`9+�N��E� QV�2d�1V��+�H*�T�I��r|*Ӗx�e��^sz2$�}!��ɽ��t����v���3T��\�K`4�8:���u�J$��U���G'm=��Dp2��*�&P�IWL��%C*��ݎ��[���ީ[�#ir��r�E���7�3���Ŝ�?+�z0c�I�3��̹�eE���YG9g$��	An���u�#\o��K6D�g�����Z�Fp�j���i6& �dI�v�ùbL��h���y�L�x�+b�Z��Y�����ka���w����k���y4s�w1��1�t$�^�̦EG޹�{�e�e�[����b�siq.�5��h�҈bC�W9����_!t�61�+%.i'Z2J6�z�wU�Z�h&=J9�2<�Q���g\�y�e��üe���Eӣ�{�7Z暠�9�t2ٺ�K��,$+��_*�5ty]Ml45��Wn��S��u�ut��O{��=͚��f�4P����|�������	HQ{P�ki`c�ޛ�A\��:ҩ�B��G
�F�|��f합_k(bD���X$]-��v:N�j����Վ0��_����'*���W*Q�JI�/��=OHA!oU����U���1���N5��)=9C��8���YҔ< Մo�Y�Wt�.�]��ڂ�H��5dѼ.�wl9��ZO��,5��<�>��ݸ�/H��z���=v���fH�<�L�c� i�������R��w��:S�/9��U˘�����|��H�:����/�仺���s橼�NTڛ������ҷ��e�hy>+j������8��}����gΟc�"_b��hUb���tGI߯&B1�\�6K��Ҍ��}���FA��C�f���+1�CFL�g:��ev��r�n1.��l���>'1�pTj�"�&P4{h���{͋֘�R�o+(�PΉO^����TK%f������\ɑ�a�����fp�buqj6")�Xp�T���vg�2���"���LC��(�9�����r�]���R(IE�K�#n�i�kv��Q/���Z�uv�{��1�u;6Spn�Sr����0A>r���)%�e����乸f��Y�(���%ܑ�=�)&�f�$�$�t�	�I$rI$�I$�E!�I$�H䜔�ʓ�:�>rq�;��H��J�'$�$͒L�9]&A��P\�n�_n�r9�fu�6G*��ts.�X]�;$�:���T�I���S����Ve�=Ԧ���э��* �4��f���,R@SL��Z�%.e+�/36�do��q��!1T2'�1��6 &���ۼ�m�@���=Z�e�]:0^�ὖ�m�i�e��48���5͆����޹��x�̶N:���p��	���%�LL�գEU 	��d�A�X!pOӘa��K_�H0ˉDXJ;���AXS����-'���l�o$��Y��QˤY�*�M��L�o`�
�`��ư@�v�ʇ�{O��a�0Ф�m���L!��^@n~�N����2��6�W4��0�o7� �y
�#D�RB#�C���0� $��U��G����wn��i�����B�#��&Qq�!��ɚ�y��=T5�4��v�ƫ�r拪�R�T�`���f��L���Qf`k3ZBʖ��d�� I�?��`H'�?^��?�~�>�$�������7������M���.����#/���u���pJ3U�.u�:-��y�J��H�Z�Y�K++v��Z�&���Y����Ev�e�%����*��{�N���*��׏qR�Iwu�V͖�85��	ʰ��p�ù2.��x]�}A���L�9�n���� ͛~�6�R�wz�Vz\0�5�3�x�r�sND��㉮%ܲ��u�acߑ5+�sS�m����cN��uV<.�#� �9���wLi��dƓ�B�I�8�i��i��a�.Ӳ��g}��Y�r�رX��mvh�9��wD���dS���|����f���>�+]�l��m&���Gq��a�Ҳ讜9�N��\Yۂ5����v���I <YO��P�������v�1 ���й��.DT�7[�G�]j��"�q��*q��|��d��Yn��β���t��ǆӣ�9��WwE���q�����sB�/��������r�AZ�<���=XJ{�;�-�v.y���Z�;:s���Q̉���#J;�)`��d-�[!��x։�YL;#���xM%��SĹ��+���X�Z��Q��ot��F�_N��j�n����&VMgB:#���u�]��� S�۰a��f��[}��&r�Ml�8�V�4g7�vZ�$3�tC ���� � B� �A ��P�AAAB � � " �UW�ԭ��h:����B��&����f�4pV�����f���8c+]J�H�G�J�o��v��d��)��A���뻖��o���r�j����.-0!D-'?�KiO�wLG��֗1��9��}��y,7�CV�BuR�#�b<���R���h�jl�2;�:݉%�G֮f��nۃG(��2���}�GF�Е��G�TZ��a�jś��3.������i�*5���SN�cU*�ݚ�Kö��ovȲ�SMڸ�WBlkx�Gsn`֧=}+�9�b�,2{l��]�5�%��N�3�
:\G>�{�4��\Ku�Y��YՆ<K6�;�44�J�keL����
f��L\齛Z�CV,��)l���w�]�m�x����i�7��)i�A�Ŕv#�}.�'����[Gl;��M���\A�XEӫ�*&(�B����y��	nL��p�Am=g�uv+�<+x����5�n��IJ�A�z��7ym&`�������w;�5ѠoC�4��]�S7n�8iX;P�x3]$�4��Tљ����X	����wt0+�@��M�;IN�$9�c���[��X��4�ݐ�v��%����a��� h_��{��=6M[f����|&�3S�)���6p8'EF��$1pb �AAP� �A �" �A@� � �A x�hƢ����!g�>1JZo�a�x�V�m��|�,�f.�-�ls��;����z1Q.\z'^3�v��s�O�f���3}�R�0`�.�d����ٖ6u�|�ޒl�8w(Ay�b�Q�r�#fM�c���ƭٛ���Y�Q�eD�%��尷}�[Ӊ���Y�߱z+n�ݱ�����{���B��H����2Ƙ�e���nJ��c�{.�1.Fbim���/c˲��<ǹ3��.=�+���JZ�FK�wav��%�%��Xr���)Bj
e�ڝ�<�kM]�;t�I�?;�T��hI��5uyjt����7�K��SxM��B�y�8^�|�ͺ/v��yr}���Ŏ�֣��We�����V�5�\��$���=o;�V]��i�joA�f� i�|Q6���!"�ؕ�p`�Wg�;&r*d��nM���*�MA������o�u�嘗��ǐ�;���EJ�
t����X�S� ��޺�r��5a���{HՀ˚�%%��v�m�,����hDa�ym�Png��+3�n�9I&��7�f9�#sب��K�����Ń7]ﷲ��Tl����=S@u�~%�� �n�i��^���0 �S..\}��˝�M��Ĵ.YHy��8a7���k�)��f�)b����=���f���A�AB ��A � �DA ���(AA1 � � �]1'n&:�mJ��QA��J�i�����B頎�mtY���0�r_Ym0����S�<���c̭7c���F
cj��-������F��,o���l�rX���\Ѐ�j��q�X� �F�-ظ�D����:�;���ϝ�qĠiJ�u䥗�J��R�Q�htu��u2�{H媖P|�9�[2�[v�pv��;'��;�wL%r���{�ڜ"��]=�	�mϺ�:g__'0؉�vˋ6^�����-�����B��lv�X;j���U�:�wm�7�1�Jl���o	�F��[a���]y§��}���07V�FJ�里3Z�0ر`��"�ȳ�)�c*��oe���	-���G��a���譨�������5��ь��\�5�<�]�a��o6P��{ol�âܼwb�l9������Zݮ�[�{+���s��;	X�VoQrӽ�p��3i�:�r��$�T݃�S����]��>x��cj���o���Pj�}�+Ĕ9�y�Q�3��X!Ζ;'ǅ&^ڮΠo�
+]k�S8UUN=O%U%�5-�[&�rJѫ��C�1l�;yd���Ũ�a�]���_B�C�s����W��[O5�|x⼭�z�R�`����S�_fZ�m�8��0�0&�1�'X�`�3�8L�'A�L�S��hq��F�t�5b4p��@DAAaA �X� � � � � ��AAAp��#�ܬX5��pU��*������F�B�I��(G�u��)�j�@��T���]η2f�X��U,DEݮҌf��5�]�×�6�
�!t�����լ.�U�-;7��n�DXy ޶5b�ZN�J�ײ��d�J�Ow9�n��䟚=yӖK�p��1�`��/%�^��5������j�16��)]�����Xg7��ZS#PI���޺�)#�=��ي�Puq���#Ѫ�݃�>��������}�D���-�]O�A�R�ڥoK��Z�:
v��C+�]pcuq�ή�w�ҷk15P$OP1��I���6V���{t��m�0k��-'t�2��[޼R��c	=�[�Oy�X�`Œ��ėJ�?�殊UQlb_�Mw-艃_^�"7ĝ��G���r�V���q����fWtvR�>��q�!$z꨼���iH�b�
��� ��
Y0+xc�Zћ.:x��������nr΋#��t����k��"�������_07C�ռ�4 �-�}��jwF�t�{�K@z�t>������޹�:�\��U�-h��#v��,�]r+9e�4���.�ҧC�N ����Ty�HB*�*�Q�[JgL�u}ӃFB�����K]t�[8P���s�:��Z8]�_,Ƌ��X��/0�]xyh��#�@e��')�WU�pc�A� � � � � B8X� �A`� �D@DA@�A� �BS��P�ͬ�mD�-��FU$�������6��7S��IΥ8�Ŧ�U�d��Fnٳp�L]wn�ȧ« !�Xo8KYZ��w:�m�׶6�'B�^nu��L0mv��:�L0w��,v�8�¢�����(Na�7�HH�a.�o���t�m�/7TGȼ�Z꼣� +�Wv��WO�Fu��7.F�;�0󖶵Y�P�R�Y�uE���A��Z����b��j���$J�aW-X�2�L�D	%p��{IBa����>�n�Iu�7����B�]����k�i(��H_L�S#�sN���Vsw�R��͊�W���)H�nf�yZ�ˌ���#4����t!��;#z�c�f�t�eMSa�~�Jx��෸�`�v޽yؤ���r���F�eLh<�.���_*��E�-�{��G��{U�ա�B���;42�6�t�ˬ�U�,D:���g|�&�����[l�z� �a����k�w���Լp��r����3.��d��y�����H2�,��u鉔k5U̥����lj���CA�X�;d�6z�f5|�ҝX�jU�$7u�+:���]SL�x�����
�c�����
��	�A���o���ӋK
�X��3[���+sut��<Ѽ-冪��C6՞y�=���A��D�G��ۑX�@ΒZ�ܷ�;&�N!w;c���T"�
�|�m��^W�R1�CA � � � � ��@D,A �0AA� �A>]!J�row�:m0.Y|���^�����CO*��rZ�-n�[�}�����1t<g�-�\� ��.$�*�G}�h@�a�����x���gy��n���rZ�f6�dɜ����pd�fT���[��3eH�[�h/�FCev�p_j���Ւ��]������5�Kg��gi�n�*N�b���y&e����T��Ym�Π�(��W*S�e��G�[�Ko��N'�\��Z�Ŝ��ech��A����;�od6e�D$XJ�� ���&�u��2�7k�b�uB�ٹz2
s���s�|[Қ9@.w�ü�]�k�Cr�;��S�r����7-�Z�ᣪ��+ۦTOo��}׺�@�L�V�ҋI���F��m�j>Qӛ��y{.h7ׂ�u�R�o�űG�-t�AK��Y� ��3�Mwi=!
��Ŏg�L��f�>.[�hf����>��B�km�qR��a����ۺ�.^e�k*R*�mŋ/V��x�'v��]��鷝�7���d]�s���C{��?�
׼\�ޗ���{.�tk�����]�e�mM�ϝ�bvf[�.gpS��[�%�8�%ju��'GZ!.�;�~��D����@K��������W��s�X�*f�U[K�}�N�!MS��Ł��9�՝��y۳-��	|��Χ�Xm��낗.q�ٸ��߂�^�����朜	���\A� b�Ah� �A! �" � �A� � �A� ���`�۷v�}����3��[�yٔ,����e]*^�sJn�B82�r�������e��q�.�Sv�ۧ}�����'F���@�&qn��r�N��'�ע��]�u#V�|V#ܘPA����fU�wE��J�s����7HZ�WcF*��!;��rK�/�q�OQ�J}ͧ�����:��:��{�?�8�,յۆ�܁�p�m�I�v�D)�5�/]�ΰ�h��⃗{�.Уs��6� ��;X�i��:�-��!�(e��&!&Y�����j(G/�`�]Cu��x^=Xm.��ȝ$��ͷa���ok!mh١��^F�/.Sπ�,���zkj�@&�7�Z��tn�c)%b�?Le��F��P��6��Ra�,�#�{gmm��˖������`"՜w�xU���cl�����Y��%�2����Bk�ԯ3׸�0�,j�%\���v]K��8H��v}�d1�+���eP>\I��PG�ΝT+Y}�T9�q�؟�n֙[�s��P�8�$a�Kn�8h��z{�n�KY�P�D!\�^��4��gۅ
�W�hM�J.�6����@�9�f_-:�I�C��ȹEp��۶N�[�'6�z(�m
��_9U��Z.$Uqz��=��5�װ�5v�&��w���{��F�ʑ}�y�n���Q������M���P�Cf���Uhf��_�f�nf���,+��Y���\KK��w	�W�a'�K�x,A�C1A� � �X� �A ��X �AA@DAA� �wϺ�u8fb���\*m�yJ
��F�-W��;-Tǎ��upC�L�^�C*�&w�3�5�=��WmWR�k��w�m&�/�8�j���k�%$��f���������}b�:�R�H%+����w�ޜ���b�\j��w��t	9 �q$��������[M�r�ܥK������ڴo�������#�Epuj�b[tC�.8��*!X����⏫�
���\N���晟�Xc�2�s!W25��W#d�[N��ו�y`�־)F;��ͅp9|tU]Yi���7��e��q��Vl3�Yv+�N��fe)?b݌��n��ׯ�l��*��e��N��j!;ST�@��n\�N�����r
;�g-҂�QvȦI�Km�$m��ob�ڃ�'�:I�x�*F�u_Q�W_E��F
w�u'uX�s��k�+e�4�7 8��z6��X�c'�߻7�P��q��naʧ|�Off�݋veV;ͧE�#7ܶ�Cs`���i����"��6�es�|,�M�a�0�Ŝ��#�m��`t_J��Z���[�fjV�ndDi��������;b��h�[P�6�VJ�2��2��0=6���f,�|,:���2�.��
m*����.֗N���%��X؝h��6uD�Қ�{s��t�혳�!����r�Φ� f����&i}|q��Qf�VRb��a�ɓ��w
am��)I͗��-c�V,�R+M�BU �	�x�n�SڪX ���J.IC/����)�f�Ver�7�-�ی�kJ�W�����0�����w���6aA�O9�|Vm��n7�lq5ƞ�+i���5�S�ks\��F-�2u�F
��(a�	�&:�`1�K}	85\UV2VNA��5�&7����hZ���*p�[:��M�B�;&p(m��.}�7�CFȺ'�lV#Ks5��������YPg�DQ�y�����%[�31õ[B)[��T���Q[Rk�v��(��3h�u(����l4��f�Ҹ���#N����#=_�b�Նl��$����R�;�η�_lk0u�:Y��y�����]>`U��ʵ��פT�l�s���!���Ik��Y�e�|V��(� �K�,�+3`2��>���Fn�2iFʾ�!�:�ow�������]Oo_�"�YY;g�A[���u���Wc/���v���/�3P���*�t�����n&������X�ac��Zf�i[�#�-���I;����1��`ϭ�֮������E[kr6��5���a��̛����|z��F�O^�F�|e��`�uǳV=�C$n�z��ΎtT���~C3�_ 3U�z�<q7Y׺f���=�����c?o�?��!$���?�������?�x}��?P���?[@L��~���TL�'2�~��7"���c9��ը�gE_�U�����Ʃ���u�7,Վ�9|��ǃxY��wV�c�/-]w�J��8jr�U�Z�7���lB��qxuJ�/�c(j��D��zb�x�L3����q�N�뵌�٠v�3:�n-��WDJ)\FHL��׵7 ̢L��P��`��v������r��JKIh����wi��r�]S{sS��ک+'9%�]���3g$r����;�\M���p[�]TL�/SW��U#��+s�k���XozcMS��Om�}�]������zNœe�q廗@>�".�o���v!4���OJ��so[�;���6�84��Z�1�w6x8,��k��:+Uf_`��𘝎�c�}F��x��C�o��YN�UT4�����{V��g�l�����J�hb�B�[����h�ț�l���]_
�{0�$v�c`)���qN�2אP�Y�*�+d�I��;�4�	�/�R�SDV�� z��^���a����1W+�/ܺ�s�������݉9Avzk����^��%�V'eM	��t҇npކ+Uc2���_���*�:������}�yf�q:#��x�I_e*�v�m!���I"��������a^RŴ��
�I
(�R?ą��TL�
�)��	��a0�m�H�!�҉�&a"3$"��
H��.�b�Q�х�Y����YM73�i�M!�%���(�m��� r��� &b��aD�a�H!�"M� ��ܑ�Ȅ���e$�`�d�ji��8Q�e�e��	��n���
��eբ�X��we�f�o� l���̔Qb�"(�˦�a=gr��3-F#�o-1ֵ���,)��Ӈ0^%x�A�*�A=�L[j��,�L�EUQq7�����$j�0����oR҂��Ъ��-WT�m�E��0S-E\kiiV$TZ�,�E�L4p���E�X�Ƥ����c�UG=�fAE�-�(�V�MڱLe
�"����g��<j"����V*e���]2��9j�*����TV��֩���"�c��,Ç���'#�����D���b��q�Z+Ɗ�k�\lЖ[1�h�[J�2ڦfQ�j%B�en&Ln4�a�g�8��2R��UF{��2�+A��d�	��r�8Z��T׷sE�aL[J��T�`%Ls.�ʚkZV2���V�[��FA���)X��	*cM==<'�>R�%�I��`�J��8&a�DL���PV���-(���_K�Z��P��L\ek ��eZ���A��QkS2�q%��DaG�8�י��6zzrs²+�"�lR���ڷ2�"X�b�i
ѵQ̦-YLpj1R���&[-(�*�\ih�yq�+t��[K+m1�"�5�+Eh��-)K�aKh�&�1��`����Y�U݅UQә0�`�F�ԭW��TƮ�..ccP��Y���-�cA��,V#m,eA(��~C��/˫�~w��}��!���]q�.Ţ���|N(�����\j�����Ua�,ۤ#�+�㳬rK���@�Ȥ��(��A�`%��NLh���1����9��8-��?���Wv��E�&���֛�W���}����Ry�xf� ���7�������{���#B26Ci�I2F�ض�72E�P�:���vϳ�c����06���5�9�wP׎$��x�Q�l�42i��UM�yk�fؤ;�.88z~�_<w�{�7����P��@�9���6<i�x_���l5K��@�����~|5���=���w�|��Lty��Au�Ί��S�g�.K��"�����H����_oi��sD'%�%������5+3��{�;��Nm��A��sg�Ah�,�۞t��	K�_��'n��y�n]����.�>��ޥo�n���<wr*�z���>C1Ɉ�>��4��>�ӄX�n����T�]^:�xB��"��LQx�4���8�͕7|�����;��EЦs�5�,(�,�h]�o\2�=VF�YV[��kiW/d�)�l{�� ���F��=����0N�3���B�n��zE6T��^�g��	u��b��=�Pn�-�gc�n,�J�X�◌�����ܗ6�Xb	ǻu�zܿ��b��R������EK1*���k��W��g�v�(xE�(��/�氷�l�o�������|��VA�X���TF��������;�@1;��c5oS+ޢ��Q~�z/�AA�8��a�﮼4K�Pc���}�w�����g9:������į�x^>���<���o���\�m�,�Z��[�=M����ɩ�22�;I]�w�Q��ޝY˼��]�^�9�����S�a�6Du�B2#�7���i�Q�V�uC:�;^Uy�$�"J����Va��9�U���"��V�p����A`�^t��1"�@�ܬ��w̑Wfx�1�[&�m1�M3� �p��`V�r8˂��¢���Ƀ�����!�E�����߁:}��j����:��v�m'��~US�P���
�#7���Y�|�b�{{g�/���^X2�D��<�����C��ٵ��5��w�)�<=���#�ٳG�r��s�7�얟��2�I9]���НJ�x4��*��uNۮr��j�aǽMYf�q�L(��`���чx4��v�_m����IV�ݮG��^e�v}�"Z��iP�'l��<~�v}h+�3��K�Y������E�O�D�Y'h��/dO�sj��P�VXuQm��G3�]��K�v:x�躻j��l/'��5&���w����Ds.׈v��owB~���پ����[�d�_��}��(._Pa���au����t��#��L__t�Á}U\~w�M���c_}�r��;_PAу��g�{]�z'�)^�{��ޞ�޸%R���𯼽��Q�bU!�-�վ6+����y��^)��~H%����9�c�,8��Cc8f����a�Y§���'kHaA���ĳ�yrj���sN�h�~�.�����Z�hժ���=�p�=/�����#��U�&jw2��#���dx�o:�|�|k��7�5�����*Ob���P~��W�	-�}ή[�Ծ��?�u<Xu
8�]Y:C�Z}�����0�{��=�שu:(=3��.�J��H���cQ�d��n�7�[�M�Bw{���艽����u�.��t�p���9�m���.q\Y�貁y��{@ە[�m��:�o%�y�s�K�1�U��&�#���}�`�s��ϧ��8�>�I
�gAPm�x-%�m���dm|��.�e�]��S���ނzɒc�<v�[f�ͳ��nX��uy�o���m	��^���~y�>&���q4k�x�>\mә����~�ٲ���E�c�P�࿋�1��c7�d�c��g��ц���r_o�L�nb�
Zo��_����c^�ƻ�	��ד����Cnn��wS7���J�~�C���PٿT�t7�-���]���M���u��f�����$�FH��ɽ�	�b;��U�(r�ξ��ǯ��T�Z�ũ3�Rw?;���zo����W7V=�W�'����.��H�|�1y�;=��{�P٢\נT~{������y`X�v7��h���g�z������"���D��$^���;7^����}��4_>O*�+o*���J��aq�7c A�!U�*��8��[��%��cv��`�w���E�3��(�ͭ�ʰ�t�v�b�]l�D���n�E�V��!�.N��5�άEf��.�F�a���RLlo)��]\�(��qK�
_Jɻ)Uǲ�K���F]��i�ެ��U�!�p��вz��U�x,U�{b{�9R�ϴM��srw�SYL�'�����T��e�l����xK�:Q�}��Ȑ��g)�^YL�x�'s9��5�"c�z:�8o�ޙ�8��\«���̻��mgS�K�X���ޞ�;O�mƾ�x'���5Q��Nv���O	Ή�\p��ێ��GQ�}���o�Z"���d�'������h��{l�zØ�E�[�!��vY��Ѽ����Pv�ۘL�6�m��E�=�;U�s���:��H����r49��$��~�;��u����9G��7-zU��;�<<������n�k���u�'���x���S�uL����\���㵰��3�u�3�,_��B�>��e�Ԟpz�\>���z{��y2�L�(!�g�u��qί(���>�[;�:孶�q�߶
ꁅ_g��[gJLU�.G��Q�1�]u�r����΍G˃�q�4;a�6fW��شs�;��
z̶�&⬭T��oA�ΐ�}�!�0������=V�:Ő&re�v�_w^�z�)�g;U;R�&�o����:i�PӁ����lK�����́�MW�L�ъ�Д�V��r�eQO���^����]ǂߦ��d���7/����;�Ae;��=rmkQ��SDlfg�`��Ϙv�,�gQn���g��z3���v�a������#>��,{)kl�5��m�l8��7�kϤ��vl]��Pk�9�����Qw��L�*]�J?!�`��G�ï2�yn��[</���q�A��}�]���Tf����s`zy�+��ߵR���(��;�A����RA�ʂÇ�tX�wi��+��G�M�:�B��ټ������h=�R�Fod��c�AxP�y�U����m�)�q�H�K��V�ݷ^���K"2�|m��<:/	���N�)w^�S>�jl���vݸ��}�-ℋ�a��==Bf�|r0oEg	��𙇷���2\�}����y;���)��>�Ӥ��lʒ��X�'I\�e���E��2�_3��vu��}��՚j�dW���df]��
4�N-���oCӽL,S[;�&�c�y��C&�k�˭Do8/՛Ij���ːP9�܂���Ӱy�Ӌ�VW���t{�g��
����2n{$��s��xL��DU#�4�z���z�J��y�(1���\��>��ߴBi��$X�仂�WpCù����7�#&A<j�/g�t�u���zlQ�59<��$㡖~��ϼl7�����>��y���M��2�t���jk��N��w&������&��n���h�
������=֛��z@�3��J���U �%k�l�-q���ܡCj��_�g��Z8o\�9�d 2ς{A�#�e��~�-��ov��*Ʀr�Z���ꥹ��zI��څ������}��!z}�X]I��7痠����zx\
������o�<F=
�x)�_R�N���y��%�72Vf�����}���`�^���}�[��ɂ��k�i���/���;�D�5�x����^���^�u��٪=�y���W���_�]U�y�yN�	�L�;�����0p����g��b����V�_+q��j�x�\`����r޻c)ծ�s���۬�q$:\���6�Y�8�Z���SrK�T�Q〤Ė2�0-�s��zbT)_��]SMSᎱW����]w�ʻ��������3���ɠr;��q���� i��6��s��b����sE�t�d�>唃�Vo�5;Y���to����Fv���;�/�5�z1hM{;i[�#D����`�f�;�kb+Fg��98_�ތ˦��pE���\͞n�����B���"⽩�s��������A�tuͦ|���VL�v�b\�6P�<.�H;�a���0�O���t��vu˂y����3������7J������,�l��c�Ϡ���׈C.f�O	��6��g�0r��ř�����X^t�o�X0y����=���'��C���h"͎�\�54�w��g�p��ɟ��:=(�M��~z4c�=�r&��N|���8�MPt
�����T�4��C-��&��g4�J�wx��,X�o9����Zο��{Ob�:|�;��%O��F��4���WMi��xT��b|_�O!ø�Ie�Ǝ�"�q��L�Y����J�����wgHK��2�b��iY.��ʘ�����i����*�uX{n�����=����]�-�Pk�`j<�xnᬠ�2��w��9��\3q}'�}�o׿{U��X�*O�B���^L&���Lx�����.�����r`��5=���sڏ΄���ߖ�����.[��������"�<�#VǊ{���˭�w7�����Z�u��UV���Tf�xz�4V���{9R��|��}|��&X7��'��^x{~�]����W�7�����]{�0[�ds�vh�&�v��ި>;�8����ا�Y��"���A"5�kd�Ɖ��?T���u�/���x`~�ư���נ��bǠՏ^�_�I �˓����nۢmG@��j�����ˋ�o}�vh�v{�XǯF�<?�%���3��c�=�ٸ��j26Cou�$Ϩ�����k�/lm�ۋ�b��C�R>���F�Y��c/��n$�{I��{�fn
P�Eq{�ǂ���ylk���;l�Wceg�{_��yV��C8�1iB��A�x�A�mo@�t�'�nc��vgS�1 H��]·G\�E��e�هJ�Sc��(�2����I�F3w1f�f�-߽~Yd������� �m�kA���r�_��SY�$���./7���xj��;\�FuGT�շ�8ן���V���EI���z{ ��+t�.�Pz���{S�8�.�ѱ�]���9�4�<m�N}�t��⠍a��û����'�n��@�ul���f�tvz���[���Gh���L�e�NP~S��m������CS>�]�ϭ����'����{�oݡ�}�r3��{���r�Kh���}y@���Dл�3��-!=,MF���4�����Ǜ_�d{=��S��/ En������ޝ&�8��p�����B����2h�1LJC�@6�h<�گUL�T\7���vj5�GY�Y�-Y>�pOH���$s���xH�� ��ec�J6"�,�������o�K��Xo,v�uuoc��wEC:���)��v�!�ٷ�ࡁk��`L��e��V��n�=�48���/�B��qGûO3������{q뤊\6-p��p>`θt.���]vdX`P�턆�ő�V�����z�^gX8Bn�s9�ɂ��,����x�8(�f�M�ڶ28��ܮu��"Tqc*���Mn㌻!>�QYƶ��_)k��RP{�"J�%
o׶��:����i�Z
ⷂ޺��Ѩc/R����ٳL��g�C���m�ww�a�9Y|P9Aj�|��Eq�:�[���02^�@a\�-�+�%�ר�)�%��\47x{�ڮ̧\��y3:.�Z��c�����f�R���/W��<x� Q�wz�x����n��t���֕Joz�K���sx��n�e`5"��W����Vdk�P�m�H�{���̀���.�{J3����T�6�G��x6p媹d=tԁ�Wd�
.l]|�6�<Geb/�-ۇS��ŵ��4��w��]���W�l^u����U�3���e���\Wo��X�ۖ&Ҥ^���{�	����7Mq,�7m���-��B�F#V��\�e�LoNn� n�ĘÂ�\�C��P@��\H���!Fr���Z��`���x��܍vC���s#�ɕ/k[�F�;��#9zX�ף�Z�O&V��_;�CӤ���[��0�K����JY�b�/ߍ�;�;֎c��۵u�*�:c�u"p%�ي��e]��;jss���T8-���夷�R}�bv4f8~�;��������Y;�z��j��02#U@�6��սR��w#ˆJْ��Vκ'�θL�v[��v�F�D3*�j!���␜�+���I��\Ф'g�sF�*�
v��G�K�Yu���꒙�>,A���t���8�(ݦ&�{��&�cUu6�+[�f���ݮ�g���B�j�A��X��D��i���Y�j�`Ѻ�E�B�5r;6U��M�#���O�e���̼�hw{Mgi63z�C�V��<{%P��"��%���\��s��u�)��Sq��ڬ`����q�N��P	�!��v�Aԝ�j��Vβr1�ʸ�_֌��׵Kn�:ֻ������uZ�m��
�{UH�4w�sv,�U���;�rZ�g�h,M	�;ǴX�[Y�=c�ص�1
ib�b/�����rZ.��Uؙ����dͭEa*Z�ܐ�V+JZ۴�E���2mc�w01�9�t����Wp��f���ݻ���T����T�+���ە����B��B�=F�5�p�^^5Ho+�ω]P�V�P滑�rq9�P���HA�@T�K�I(�d͜������4j�{��4yq.;K4��,���ӂb��Ym1,�&AeF�ʖ�j[(+h�Z��i[�E��XX0X���eQ��F���N)�*��Z��ㄶ\��Z%��Tnd�����W{�+r�n�X��D�b`*açM�'%��|����";�Q��uh.�Ŋ�D~o0D]6T�D�Q2ݵVED�4h���y9��Q啋
�c"��|�`TQD��hQD`��vc�+#mf�#���|Jh�ç'#bqN\-*1gR�T�F"�>ڢ�A�����JoZ�i���ak�DY�UH���M�:t�q{�x:R�
�R���)����L���Ŗ�b5(��F&P�b�V
Kk�*qٕUf͝:p�
��cU���aDY��m�E��VE�b#�P���xxxp�=eFEUUQm���|��T��׮�c`�R��x*EU���FΝ8q^RV�G�Qb*�U�UA��(�X�F�̘�Uv�� ��*%���b(��ȃ�swHE����lY����N�/�}�����5z,��E�jE���6�-U�l��+U�d����޶���fg[�R�0��\�l]����d֛��'O��m?����7��ٳ�!�oA!�q��q>���B+�k���dE0�5�g5wa� �cڣ"�	�����_
���"���n�ћ��[�%�4
�W).��ٲy��Hl8V\�X4��V.�n�4%�-a��q��AoO�#)��z9�r=m+�$��ge5��S�3�c��S�8�m�ocwT5�6���Q|}6f�썁$�`)�2�Q���%ӱ��Cx�M�2���3R�sST��N3��ۢ���0>�X�Kj�vŰ�{b�ר�h��d��V\��Hyղ�s)�4�*��r��'KE�G�F�7��GB]IL+ʺU��Z�C����+I��2���O�Xe���,�����_�(akׂF��1�d��)��
��YHK�55ˍo5�z��	W8���i]<��K��3�Oj!��PAif���}�,�a����$��S���"�U�9��������o�V<Dս�����h�4!�!��a�6V>�����u�m�7�j"-��A/������3c)/SݻRf���׆t��2ýC����D�0�<g���Z֝����+.�2˷������lvUt�V��]�n��h�*-�`�m�R�͛ ��[M��u���r���7c�����7�M>��^E�e5\��Jڂ�7J��Ƭ#a�u��	�K
hJ�NR����9�(��:+Fv��\G{D�r�j�C��	���sr���bC��4�DP�k]�5���� F��}�c0䅵SL��^���J��7!��3A�υ�n�Zv��P��Ђ�=f����O��z���/=�Չݚو)ٜڛR+h�l�>2�OG� η��KG���v����Bd�mҎQ8÷Q'9���P��X��n�κ�ғ�D���m�+���c�OS$m�rfa.���m<�IVX��O�\�_�X��H̐Aǽ��'@�4]�ñ!��w1M�,�NE`���t��j1�(���@������}b�"�����o�&�dD�Gq�f�XŁu=��7F��	����!���E�7ȎN��`D���|mY����N���D��+R��n��[�3;�k��vAc�C&J��%�Lz�c[&dY_.1+B�/���v�>���4�3	��M��B�#dv�I���'@���렌�[�}ܶ-��M�/Nz��oX~��O5����/բ�rR��V=h��l�lck@@NO�=tB��d�$!��)Z�,)��5�G��"N�!�b�4Mx�÷�c�U�����<���t�[H�}T�
>�je�KYb1�4�#�:���U7+����X��e��~��f�oZn�l�:;�4T3�J6y3º��]c�{��yt'��i�*p.�2	r�'���Vt?�j~��X-FJ� �ʽ���#�A�F�e���Si���/B���y�O��-�$���9��:�#C��?��AXu
JqP�X�ZzA� T]�E�fakU�l�q��9�ΠD ��H�"��j�2�#�*�dY�b�bMNvh��Y91/q��[�*��z��7E�B�ލ��,��p#�@�t�e���	��h01-�z�k���T:�м�)��:�78ր��;bt�:�:X57�`���ه}��v$�l�ڇY5��@��A^=i�5�͕o-j�q���t��%�&$�����> �l ���ʘ�|�N�Z�su�V� �|P��Ӵ%l��,�%�����6���������6A|!�J�\�ST{��Z<���@P���5C[X]Y�VI���ǥs�T$�-����������|�y=X�n�E��w��L)pa���b����3,�{E����&���eӂ[��O�j��ݞZ`��6K�n��@bqz}#=	��80br��9%"�<�յ���Ɗv�A��oz~���iK�����v���� k�o1�����EW�)���`L]�0��P��Kz�g*ǥ:+��Aϕ�f���X,�y��\܈�����\�T;C�͏e<�A݋�k}�V�ϻ�÷<[��}�Q/%�d}�`�5t�0�'��=�-�x��H�ƅO����Mӌk�bnk�DgW%i�0�br��*�MI�� �kܬ�z�^�@���r�gC��{�P,4��i8#�ʺ6�%��g0$!6�5M��:N\yu�e[Oa7�qЗ���;#o! �ݏ�0��ȱ��͢�(�4�����X˲ӊ��%�!���thel�,-����{��j79T)�\�ΨZ���x�:��zm��P)o�y��}�ϳGZ�Ý�h~8f�?�h>^Շ�mC���D��@��ʇ�*�sZ�1)��TDF��|�ez��v�zM1g��[HN&�+� %,�_W�n���G�'4g,�qP&�kvRf�W�y�XP��w>�8�E��FɀQHa"� ��+D�+3)M[��k5�2�1��]jw���V��ܗBb|��/\
�Ӭ�f��� r�--c���u6q;���ۣ�����շ:���)��a��t~���[=���$Fy�:6���O%k{�������ŗO��.Ucz�{M'qY�z_�E�洣ō�y.5�"�tݺ�h�������(^`��a���PD�a�9{*���`Z���%O����Gs��#��36��N�]r��w�N?�׸/P��vި�V≽���|���������Ex��,��C��6\"U���ٍ�H�Hx;q�A�Es}�Qf�l���yW��GҥP�'��曤���-�;L�
�qg'5P�*Vq�S��Ύ� .��~�OR�"��P!�?�
<�,1��{�%�P�����Mc
�ҵ�n֝0�0Y��r��h��Ց}\�i�]Bv�;!t�+�`'��������h��gK?O��)��h��^�U7�k콠8ϧ�8�4��,Ɓ��c#�3?��!�`+���9�BUcZM�iՙ��M�A�w�"�8����=%�C�@�1C�P<"ڤ=t-��A.���z��Y{��Zآ����3�Ǯ>BY�CvCl^M�v�>D>�D[�e�}-���үVu7B�tq���h�Z�X1Ɛ�`N���6֌4���n���ь���kݒX�B�K��ІHh׾��#I���	�^b��a�4
goHC�4�tz�S�z�i�*f�Y�A������0���Nx���8�����A�/"�͟MR�E�q`�R#�v�Mh!+��ϱŲ���1Wd&�l��i�7Acj�M4�J4!l[	�kݙ���f���A@�5�4���	���?<����-U����>l�6��Dh�!$�A.�eJzSU}�m�i�Q�G�K�^qe��'�����2���GǗv�ϯj��x��!r��r���{�(^�p��ٍ�,X�P�~�yK]P�4���XU\/����.�����f�X�ܻ%��Yn̩p;�·�>[B�=�S��:��G�n4��AJ7��u�T��l� ��x�[���ԤF0���8O����x�I��Js���$i5��}f�.Q�4�[3 �KKmR�N��8�1���=},�H�a���4��.�!� 3��YZ�X��ũD�,��ٵH���߽���Y8x1��0�	��/e���
�i�2���|�ӓ���&��=8ѫ.��,ڄK����ADp��j���xr�E�nx�1�=[�����6+Lw��ږf�4_����(.}�>F��K8Ƕ�`��t!w($|{� ���yW^�]*5���t��E�!��m|���8��y�+�����v�;���x���7��_��$Iw�l�w+�w�+�[NB�"���,Pc����^���{�����Վ���3^D�R���m�v���Rۚ<�6q�-&�
� >^�DpZ��qhA��*+ũ9���6K��ǝ��U����B�{����	�C� �����~���7{}`K�^FF��ٓS�y�k��b��2��>)$}~;�_�B(�P��D�z-�a�䊸zk�׏쫭�#^�^���3M7
E�T 9r��.}�.��L z����wlT�U �Ɋ��J��=�/�1��dLu�*�*�c"�>��g�
�����T-k���y{u���U1�T�S���u�#$���^���e477�Uۜz�,X�l
F�}�V�m���'"֩#d��M�a3� ���o�"���$ݼ��cG�>���~�4hٔ}�LQ~��$�9�G�{`�i�\MO��v�C��ܑ��g�X˺;C�n�sH�q�<�-��E2�n)�Q�2L`��$��0�=R�Y̷�]]��O nPp"m�u�GZ���d+�,Xэ�u�6K�X�>��V]�[S(MfT��^n�HR���l��-"5�0&��\x�h��̄��%"X*U%�5.��c��e\�"6�wK���{^z<U�>��|�����5��#ͤ�H����p��R�c��p�#a�z$�A�z�F��:��o8��m 9H&�U����^��O��Rd�0�,�%;97W3�(�]��!�z�T�/A4��/����a��{hs��q�L
�%�ݼ��S�6U�Y���Ӻ��[1�u	�
�m.�2��'y��zk���c����r��h�t��e�%�C�n�f��Il4,��ѷ"r�jSy�e\"5ᦕ���n��%�G��2�Ƿ�����k�P��W���Y'����yP�`Ĝp,�%��u;)��q��5G�����\�e���=� V��ݷkd����GXr�+�$-j��R����-#vwe;���p��shN�� <��:�Pw������P�[��S��8��7�׭���2��x'�S�&H��2�Mْ���9D��*��m�U���{�Vl�-���ӭi"T?S7�����`鹜q�Aףs�Z�	��8-}¹?q����׻.�E��{/{�u*-Cf�Yd0HX��u�86�H�fW��a�7�H�!�xM+s��Lt�FWF���:ra��]��{�:�|$l�0p]򏶢H���l�-ܭ�=Lc���&7zX!����N[�fF�C�hv|��+��B? ��(��a�Ҏ�y�fت�Ŭm�t�U�3*ޑ󉡽A��H��9t�H:"�P1鷆U�!�D�2)^�`F�!t�-1��AB#����mY���ߘ9[�x�(j��I�)����V�AB|���U=�G�l��B�(F�ڂ�(�_
���2a��ǔ��X�ʔ��\� Up���L����+��*��,X}���6)��9��8&L8�y�c(ن�79���&C4�f�U.t�;�N��ԣ���ܷNx&lzy��}_\ߍ/�:VB=�>��6�k�6N�;�����uu�O�
���x���V-B`��P$�mTm����l�4�R�C���J�Vn�Y�͵c�%�vƻE����!�=�h�F���i�ۃ}F�V㩰j�o/����1���HsO1�j�{�&�KX��m&Oy�x���ْ�I��x�#ۂ�o�'��]�ho&9��yt�6��ݩu�H�F�eBL�������{»�9vW�O*�]0�,���L\R�����|�+��U�=?����]��x�pyWZ����Y'�vR��Ȧ���l���&�^Ԏgn���%�a�d��\+�q�y�t��f�2�vni�!7�L��E�F��B ��]/V�N'���ņ�.�����Hi�r#\��BP�j4��N��A��.�|~ib�
�
R�v��3I�I���چ�5��m� �Bi����p3��~���s,��A�;"AW�������V@�{׺D��m�7μ�^��
Q��sۃ��?A�P��
x>~l�_h���l���٬�MwB��^�c#[S'�7�4v������>�;yhp��h�_s�2�*hӵ��6�k��v/�q,��w�C�0@gA��c�tE��@:pǅ��<�4�-�5����P���T ��v��T� (�C(�6 ՝aۮ{6��4��$=D D�=NŴh��fSV��K�nY�{W��>��nq\f.���4�"�#�f���ދ��f��X+(!u��m�أ�ɝ�vb"�ob��j�]�2��l�HH^)��.h*�����x6���< U}�μ�*^	����w�9ݛ�[4����yn��C��<�[o�egUt2�)�a�����X���U��o!����f������=��+ٜ��䃼�? ��x��w��UtR3�(�z0Ȓ�AM->�.STTe?0�G>ȶ��S6^�&8>jw���K�N��޴�����bћ3GΤl	&�
i�WG���S�A���\�K�������.h^b������ބ4�J%
v-��3F�Fh�y5*��8?Є-�~���^*��WF1u76ۑ£:��?B	�1,��%�,�)�MT�m�;Aي12��ޢ���砧n��qhT�>�m^���H,!	e�?D�,�����ƩʂF�_��nO4E>t���ה7{7��b�>�1�_.�T1��C6H��ʷ���;�ϑ~������et�_�V��6�`��u��F?9Ә�@`��Bn�L�7���NuD7z�&�wR�#�+|U����QoX�H������R[
�t�a�C�9Ab�FlKm�6�ĠҒ�{��{J�F�Zޫ9��y
R1�́���Q�F�r[���6�0;��Gz��Ɯ��R�17%��5 �i��5����Z��'�lF<�+�@P*�e���wf�q>�B��	 y�����K�͜���2��/?-
��ڧX���ӛ�M�L$�ǎ+�\t�D�4H�����I=V1��sk��V��Z��1)e�p����<��+�(�sGZ�+]�+If�r�Tn;����X ',�Rw�L��7��;gN�Zs�E�,���r�5��}ʦd֬Wj{�]	h�8�w�eK����H�#n���ӐA�ɜ$ی1H�cݗ�ê�d��,i��k/'[A��'7�4�w<�:Jە����y��ٕ�|�2��V��L�q�:�e�"R9D;��;0ep��ɾ�@ř�֦nU�Y�X�MdX����M�'֫�	Y1��jY���ӱN��
˚��i��w�<&�Puׯv+�MA�{�4^��fh�fӱQ���n'PMع!���y�����<Qǜ�Zt%/n[x��Ȩl�#Զ6�C	�P�4WV��Nt�p(�]�:���f
OuM�*w� �L���K��A�hu�Hƣ8(�#j'���L��NV~����.������h����T��-���t�LcXcr���;R��A�";�x31���;p��c�{�����)��s'	{*��%����N�N�˝6.^�ș1���r�C�4w��C���{�a��WnQ�_Z��5ɍH�X76��,^>v�.w}TV:(�nܓ���֛�+0CE��w	�I[WG`��u^�M����|�/ݧD�yԝ�n�#�g_F9V��6� Ȳ�L���Lh� �7S**��)�Î������!^����N^`������j�k��t9�E���x�b0`��c���uu&뻮��CX��XN�j����#�(�f�M'�T��ܰ������M�l��]�j�\�T��dLuO���K�KOZ\(vA��P���!e���(�MYu���E,�`�*���g+S����c,Le>�6����0�ͻ˜����l���4����xV1�a<N"y��Ŷ�t����t��D�C���Luj�Z�Y6������Mn+�qm��h_n1Me�;.�nt(��EuF��ڏ^�<MZ�*���p�hQxa�ꥮ�L��1�/(Nu+�Ź�&�#q�B�\�F�go&�{����C8cks��\�f����	������{�Tm	��p���*�\�b�C2����˝C_n���K|"��J�X@�~.k.T���'��Vi���Yce4�V�w�%x���`���*QN�Hɇ�Y���0n";� ,�N�V:�o�����k�@Tn�S�Zd���C���1͐c�鲙Ѷka����+z�u`��%:�Y��@f�^�`۰�Nt�:��{�:�K]"�v�Ĭ�@vgQΠqO Z�����)um�틇�.��I�}�[��$w��Ծ4�.�+᧾0��HN�*��d�I7.f�Nm�I���KFlª��X���&	A~1�\B&�H��JP�cfF�l��n1JڣV��(����W��  ��zCW",QTX�Kk��AEb����*/-�lDçO�娪)֑Ki�DQWIDW�TEQQfZ"(��UQ�D_DSTM6t���QUj�ŶT����*��2�UX�B�V1�.�R�s0ԵY�˦UU�T)L:t�Ê1d��F�D�Q�TP1*����UU�ݪ��T��S�:pǈ*+�P[h�"�ȵ**[e8��EYXfb����<qX�M6xxp�(�z��_YTަ �E�F��,`�IU����b;��v�X��:t���V0Uyh�����k`�>�Ĉ���Ei
���OmX����:rp��E�VJ��X�i媣d�QgZț��Y�\ԥ"1e%��c4a���������ֳ���,X�^�QT��J�(�Q

|��Q� ��X;lE-�l
�QT+Y�Q`�O.y��_;��<�R���}�a�gos��<�{*��|�}f R=5j�+j<�Jr���:[�X��	���2ڠYۺ��Ξ�77t�q�.�L+MZ�n��j2څ���� �+�z�}��o�<L����b����s��*�̖��V}@wlzq�5�q�Ѳ��%���N�_5��*�6S^�a��&ƀ�i��d�>�T#p�N	��,㯼q�O5ҁ�'�+9�������!t���#��.���bσ�عVyȦK}�@�;=Bw���(z���SQڽ�W�_;1�'�K*O��c��]H��
C����?�_\vr��6~�*���[�r]A����"�v� �!̞vA\[ �5t�6Ԍ�/�2��9�@B1���E�%�lE���(a�kEȫ���MkOlP91j+&^(α�yeDKht�Ɖ�d[�2��_�(�rv�ܮ� ����UA˃>�3�^��t��(#��Ct���3�}�m�/NJ��uQ���ɫ̥���̄����6E�<"�1FA�g��ֻ���{y�PtR���0�4��FԆ���D����5B�%*CD>��m<k���
b����P)�E�e�3h��M�:�#\���������blCU�3�;�lJhJ���|�a�e��b��8�Pt<���S��:���D�j~����������t�A㬹u�o����ܪV�tb��Nhtj�`�4�ۃQ��Ў�s�HsY�j�s�������Z�|s��+����y=HL�;T}����-�o!���1P�4�t>5�s՗�l�'W7ݛ� P�e����(q��Ʊ#`O:	q�o�gzw�xa;���슉��N�nF"gĩ���Tnj:햃� +6]�u�RQ���ˊ�78֏,�$v��f�:li��q�fe�
bi��}[_@sW�)��2$�i0����֮Qy������0���2ɲ�:ջ����51A���{H�L���R󮣌�;�2q��*�
���լ�a �~i6[��L��Y,c�F�p�𨂀�5��S�74��	�b,6�ϯO�Z�2q�XzV�NK�(��x��}VfLԲ��ͅs�R!y��Tk���ǆ>�h�eSq�-��)�3�{���yx���\\�@�\���������x��_� A:8�#�]�u�2EN	}�<�@�n�Z�;r�I�^�÷c��iD[�F4q�0J��h��ii9�UZu6]�3Y�Z�00i�n��
��x	�4@b��H�uCQ�ʆ�����n�֢L�m4���q<!A�Ȁ2J{��zmǶ��$`�n�,���B�|��|�� �����/��%���C6bZ+Ϊu1�8c��l��iA�A�WN&�L����
T�^m<�M�b�+������2�<'�(�=�9Ӌ�I������n�w1����)��ȹWc{v�S�V�^��.g.vfUR�j��K[ޝ)S���1���=g}��SᮊcC��aw�!�������'=R����Bװt҃EYB�7.��~9��:U{��O^ �Έ���Mn�R��}�i��c�����޹�r!5�z#]�dK>�Z��A�ж�C|w�o�(R,#�Ѭ��Z�Ճ�d9�n}���I����b�J��0Ӛ��������P��1\�Nx>Eٟa�.�5�bɒ�+���6��!�E��Zf��*��g�3b(�����-�t&u�H�j�џaƷ����-���Ӌ �NF��3�:k�Vv���j�0����ֶKu���Ķ�uF�[箢�幺Zz�4�K>d��|z�=��W�����]/G�5���[��鬋,�/{OD�`[9(n��>W��i��jbK�����	�J�/"i��3Dq��{�~.�S4�����_�n@����`�Ҙ��w�V8C�����T]���z�	2y�%�U���]Bw��@A_�s�w�'R!���ƛn5�ر�m{�{qBC�gs���Y�j��l8��o�B3['B��m��t]�ff�~��V�f�mq���YVm�N��H�Z2���S��r"it�b��+4d��c@gv��3K�A�V�Q-�:�q���
�!Ӷ>�R�9K�nNs�}���U
�@һ�
I�3V�Y�m��� �f�9G�܂Ϭ|v��׌Xgc#�38�`>n�����˺�$پ7�z�(�P�S�un��v�;)���>a<����z��0{C���>�؇R�_r�x���m^q��X4����<(�.�e,����]O��x�����iZ.�y旗	�DeL���5)Ɵ!���[�A�C@C ���$�/Dd\_�hkH�Φi�{�K���Z��|����k��$,R����ʿr�������0X��z�ٶz�c��F��lջ"b�T�R�
��i�G]�.�6��HeV���Pz�ؼ����F��_��q@�0�ѻ*�%V``��M�.�a���9!<�c��ɦ��EF�0�׫3Fh���d!..s5���P�IոN�	��[��1��A�]�:�D�QКu�h�O��b�u�����5�|���چ��"�`d�x�͓�~`�V�h@���>:��O��	��~�"�ʒ4��:�ՆD�s*�6&&b���NT������N9���a�(q�D�=8|0�(�v2����LSʂ��A�<�Ȁ��C�u\�E.rl5�4M�3�:�&��ok���Z�c1=�f�s3+teҊ��wa�%E�Wt)V�a&��D���g1���[3h�=�:z^u%����eͅVUd��fd�M�9�~kZy��g�y�.~}�IJ�(�@�������ǣ�Rb��R��p���w)�i�{�����A�p4�����k�}Fo 5~:��Lnl��fhB�[\?k�?�AӂySG5?��`y��RX�"]�K	
1�p�)�,8�clU�����-.����oj�8Ա���ۜ�$��Q�Pn�'�Y��5������`��u��+��9��eN0H�ۈٶ��H�R��0���#��K6@�>$?j˰���|���N ��? ^��H�i��dR�2Xu1��잟Vܚ���c�?�}��ꙻ���9��]3��wC�g��(X������9ּ2 �7���/e":�ˢXO���ئɝK�a'����`�?s/YB�4�Hiv8��XG�"ac��5����#*+�k�gsU��Γ��K �s.:H����t��p�א!�0�֏<:ET=5���/������(9��nF�W�JdD��x��Ql�H��Z(�R24���@�ls��#%bCm�D�}ۉ���ٽ}&[q��^������r4� Ũ���1nȼ�e>��k�2J�6*��N$Yݻ�Ք�?��B��M����>ܽ�,w��}p8vڙ{�_5l=�[en�v%�7��q�!D����v�~~V]�^�M��?dM�u}ø�5a��<�0g>]�Sr1�C,Í�\�0�Ӆ�3�����u�����D�������7��*D1��s�B�,G�7fXHx��E���^}~�Wc����%�����,8�����aْׅ%Wg1�K��̆�6�.��/ŷڐ�b���/�fd2��v):ĤJi�t��;���}��0UglA�RZ���e��Y�6M���L:E��E��kO��2F�0��<�R"�&��3])�hT-\�)žŰ�vE�.�o`�c���6&��h�jbղqO-�0j��
k�����s��HLV5H^��C��/��t]�{-à��C���3Ax��ʑ6�'m3w"E��%�ꆑ�R�����\U���Z�0d����E3�.�酅�-��A��]�o~>�@|.���:QI͉�B�t��%q��.�ƥ�+�]�bHݔ�3�T�l�}��-�Jj�0)����u�U	;B��b-��p�&/�us�u�`ܗA�&j�>�)�m����Q�,�� �����y���8N���k��t�TGYM�D�U���b�ka�ti]��F��"B��<h�C	��f�Z|��=b��fYS�1�NH3�t���Y�1W������[͔�r�oU.�ea��Vs��am�"ܮ=�p�����C����@��ze�A�_u�˘"5�F�H&
5ɤ.�hա:�%�3���Fs��F�Oo�p밍;yS.��μ�4�^��yӣ���# D�$�FDdF�����~�|���<;Hw�Lֽ����f�O@��(̃"]぀�	�Hx��)��k�eqwL�f�ֲ|Lӯ*����YE��$��-�doD;v-�D����C�DJT�]M��o�}��<������3�5�fK0z��19�;��$���@���\�}�^o��>�� �+�2�v���H�q绌�^�Ve��5��D<�vAʸh�k��UV҅����X�-���oEp��g���P�E<0W�"!�x�pcrna���
�YA��u���h��F�9��2��Z�ϱ�a>%�.�ש�5�[�q�^��#c%bv�,\�y2�
��
8M�8ڀ&AeiH��+������z�"�.�A�L�9		�^�\_D�ll�\w�U/hi�}dw9��Rg�/��	�c��NȻ3�,�3F�q �n��;\=��ݕ���Q7נ�찃9| p�3�脜��c�SlSH�`��"����Q���VD�Md���T���vl�"<X$��7`���X��>�.�_*�]`
���S��^X����퍒i�ᛁV��ჶ�f�D���F��}�i�t�~�'�y,/J�}c�qY����pK����x殿h�Ldt���'�YЫ*��>�KN�Lz�t�N94X��q��M[R����׼%]���-�1��$�	�$ #�$��# `������R93
t�|<HoYpL��3cO��&���M�/�
7����8����Z~bXf���OOMf5t�)�W	z9�L��h���������>6�!�W���-^�r��Ou�j^+����gR՚����{�=}=Ʀ&�A[�hd��n ��a���������\כO����Q�x[��v��20mcZ����W�ό����&d�3�0���>��W�۶�]L\�V�e{�I��',�C"�,�������/z9O���9��3���@f�F��+���0��$����?_-�����'+_�������-���zN��-4^^���뫴��"�'b���"'����ā�6hD�㥻!��mcm�9!�8s!ǧ4��K�3�P�l�,reG������H���L셞l}L���3Fz�d�k��f��ny���#�v�0ŋ(A.��<�~�]�a�/A���鍛��3»��{�@1�����G�'�S������u�7H�Ú@K�A�ȴg�f��I{S=���E�Biv]tޡ�w
�&�^8��Cu���+#�Y�X�5�WְӃ�>�1�}��g��v%��w���R1ά��0f8�]61�C(B���K��(e]�����y�r�x�
��s�k�K[O��!l�)�c���/6٘=�bC�e%Cc�g�/��֚5��~�#	$!�AFH����{wߟ~�yQ���&�"Z�
��v
?�}Җ��3��׼�2�{ԔR4�[�4e�L�o��h������HW�������)
�]��t�	{:�㮂"��I���+
�,�&;Z�J+y٩��	���9�{XѶ�x/	
 ���qi ���@����'^H߹��P%����T9k���/h�=nN���uML�\kI�,����`튎p�0XrT8�I���x��Yn# ��כ��f-�e"�-�a�@�����80����V����/b�x���K�y�!ow2]�q��{�Z~A@%�s@Ԍ�	=�C�C��9�o5�����""'����**�[hnl�U�%q�N5�΄�t��F��K?�1��!�:��r�r��Uc�,).�]�
T"a�&6D6���5f�#�޵��b�G�)�#�dȺ�̗G ʅ�1y{�u�L{�������3��_@���sHm���a�͏NT\ٻ�����i��(�tTԨ!��P�c��0t����� �n�������Y� ������atL19W�Z��hmc��<�^��S�7�U�	��R��AP���%K}y�ua���]�O/��6�a��6������&f���C��
�<SA#��U[s���"��)M�:��E�Z�3��[����/tD�by��L[���ָjuWg�}����kO�͙�{���$�$�F@��A D�d�#!=�=���Jt6h'>+�u�#c�A"��b�����4'Mxz��!ŲS�!��4z���U3
����fɌ�B38������ȁ��Θ��:�H�]�X�昘I�./G�3b���C��p�V�^��"3]imJ-�m\�MmPs��_� J���Ր���M5�6�N��ጣT0jx�oq�+v������-@���3����e� [y�۳��*_fr9vfnƎ�PJ��6Z`9�2�^*u��f_�6�;g�SȦW�Z��X�Z&ӈ�iP�L��Kӝ�p�P�.|,D�>��-T�9z��':!V��1I�a��j����
����Z����|A�x�{i�/NUp^�p��p�
�C�Zd'��6;+7s�k�/�ϴ�����35Ί���)žŰ��кD�{=@Ċxd��be�Pǝ��e-�!g�h��6��7ٝ.�5Q��ax	���].2	�8_���H܁#�|J�T"&���Z�rT8��4�s�m�6ԻF��#5��x�na"��f���łe_�h| �o�sP��*�7#�Ħ�:��ޭ��^�`nQu�0�|��`~���gu��LC]]�h�:ɮ�f��f�]D��Q	dt8�hc�:5wj�u{�J�߶�|��Y��R*np��s�j*�l��vm�*] ���8��r��̡��i:�+&�����"��t�f�r��$�%[<r���Q���ؾc�W(ju�*ӧkR��/"�-��*�{��֗zM�+V�Gp��CY�Nv�Z��tp0%�fvo�]�(��-ԙ�E��I��/��v�i˸���P��Y+h<(༼}ۨ��iZ�7)E�	�PF��CC&�u���U�3�/��P��K�7|�d8��v�L�G$�����Xb��j*UB�5n�N:�?=v����*`�x�S{pB��p�z)�0�x���h��u�|�T!���F�`�wOq�*\e�1q궲n�܉��9�f���[w���-n3N���6�f�E�h���Q�ty��Ζ�k�m��TDꕇi��,���� �s-�hm��t��4j��+2���'N�ᣍ�v��&#v�3gUf!����]�ĩ�+ݝNȖ��e���-��͚ō���!] 9�-q���6�����+�҅1O*��:���Sq�;�:���l6ҪY���rw{r��/g�=u:�Qo��\v^��8Og+��x�/b*~��D�̀�9[۫5'��r���*�=�~�z����S��K��R�G`��Z9��Մ�����&����2�bW�Cˉ�§��k,*�y5��lPj��\j�ln5���Kb�%yb2?=����sƞ�r6�'�ず�h���a���Vr�5D��H����+Pŀ���/��$űکհ^>5�ʮ�h.02�d�w�#��3�"[�Q�,iɷ�W����qn�3VW�٭M\5�u9b_3��fS�����Z���C����9�y���4	��
�섴���v�w4L���Uy{p���V��兹���[ʻ����{���<����cQaB��K�P8!}{��O�VV���v�`�t�
�Eͮ;��ثWM�S\��ωPSW�Z����e���wcG�c�J���޴7��b�w�����ɗ�(�� Ŷ�d���E0�=�^�,�u�.G�*��~�ot�ܦG�\Y�T�����t�+��N��pk=LW�d׳�>�Yu�!���5��!ʜ�Ch7W�YۼsD���G�,P�3S��
�|]�����p��aeR�����;ejj�Z���6H����c��r]��Xb[|x���5k��;"&��	��g�Q�S9�!��i�nM�@�WJQ�-/���X��r�vvbկ�.�ڷ�)_��qWL��}�%Z���AJ���ǚ���,��[#
������3׎����v�
zK'��g��|7��w&R:���:I$�Cr�>��[�02��ghU^��U]�=�KVZUUTD��7,��""�R]X[d�b�h��Ӂ<a�l�$�Lf���b�r�"��ʒ�1���RDч����6�x��O�+Vi+
�LeIc!D*����6�E�B�ç�N�QQ��X*�QATG�UA�,����EX+UX���:t��q��,�TifR�T��P�(b�*�V�*$J�E-��ܴY�O-�U�x�e���� � �E�dQf+[K�b1F$��V�0������ƌJ�*���,�T;i ��|���U���ƪŋ>Z�&�N��EDR/ZŊ�eJ�b�E��X)aVm��
�`Q,�<8xp4��ba<B�,Y4r�&�c9l7i��X�{M��4�m
��u�D�VLM:<q�J�P���0RtM� $��L(�Zu添���9��Y�v�׵�ȷ֥@�ݣOc��Iْ��`���L�YO�}�+��Z(�Ն��z����q��HO���H�FB0 # d� 	�^}���,ʮc�<.i'�����_��ƅh4�aT���=��E���,h#��,8�D7h���.;	
��du����@LS�F��'���t�:��aTX@�j�_1�V�..+_$Ev�����z����{`��Pb�9������	�Ll�{��Ŏf��?q�����.��c��y�O3mh���%9��^~"|�P\k��] �\�W�_|���� ���C>;�+�Y�\u���@ݒKj���lM��Y�x�f�څr��W���1Ç�������c\�h�{�'�Ow)רvm��3g>���,(�I~.�����UKP\#W�5D����νN�{d�>=�O���$k�aӳ��v��ߔ��<C����#�E�[b#��ۙ�y&����(��j�3�!�D���A�4���Ɵ^A!�ݐAzd��B���yUwR���#[^��vD7��ʝQM�d�}�,ha��R �<q�L���Eءv��<�HE�I��2ۜg��;��RWr'�j����0�P��X���Þb��Ol��b�
)Щ��e���k�Ҵ�Vu�i={�E�e;��J�I�q�9�&$���z����NZ:���-���$�#��&��^؇�b:�{E,���Ԩ�]ousD�(Iq]g�&70���s�l�������uI�SA���4��Ԧ�=�<�ܿ��?CA�B"�2�F@`=����IP��s[~x�	��d&T-*�Į��y�̤�Ҳ��yٟ!<������[Rf���~%ې�2���tsk���^$'V�s���EW��]�Ö]l�K�N�ð�M�n������,���!ƍ1Z!Z�כ�\��qH6��%Иm�lޑc����J����D��#3�+�y�@N͐�iv�ۗ�D��"�DQt���.����Hn����E�
zˋ�R�.�bC��f`�}�%��S��BxӁ�����;�+��Q"z�l35�Ar�-*��l'�,�>�<�a<�ZQM�)��]�M� G��bK������ӷ��Gj��/-"z�n�hi5����̑J�s�Y�G �n@�7?�3��y�v>dv�Y�[x/��Y%��)5�+�J粣�W��N?8�����]:
9�_.�ݸ�v��0�����6�h�����f�X���1�Pi���[�(�4��Nʼ��W��YM1��^�J�h�A�P��Xva��PZ�U�-wY�כ��_�:s�*+�v���gfT8�l�9!G��B2��w�+�.&,/�����L���T5���nv�ي_6�L�z�*�.����T��Ȱ:����A�B���.ί�4���GO!W4�1R�����B1��V��L����/��3]�s�=�{�9*(�� ~		HFHA$�A �����3Q�|8]���ѓx�r�hXž ��m��A��W�VR����l����۪*o�*��޶��EHӲm����5�c�1��a�~05g�EV��7dcc�+v�cnL���m�*�4%��9*��j�$ǔli����b���C@A>��px��ZA���K�)��i���*f� �ƅ���7!�fE�6f��Iq`�jޖ�+M�u��w]l�O�����mA�h�>�A�V{zd� ��Q��b�v��tf���a�<����R,�mc���͉L,����%�N��레��X�J)�I��eE��7�1�kws�U�^Ǧ(�h�E��bԈ�	L�� U��נu���;ƞ�� ���%�B�i���/bT�����O�p�s��b�~";�s$}�vO41F�Ȧ��+�Z��a��*��b(�X�"�ymsj���}��l!#��Bnɂ�r��kz>��Y����s��O:�3"�&�z�Z~X�A/��y˅�`K�:�l2C��/��e���`ˬ8Ļk�a�������`��u�{ ��P�[|c��^׀0�����*ސ��p�L^n���ڈȕ/��aw�Z�1���X�h+uuPWL������^��Z��)����Z�hWoCK�m���W�^��_�
�H�D@$D HF@" I$ ��>��<������tyOɅ�0���nۄ�Ӷ�L*P1���O�SZC��$~��9�YՔ[�?�1{G*B�����%��b0��l	m�ݚj�gJO͈���Ϡ*����jI�Ҏ�np��gB݃`�q�尮2�k��B�,;�Ʋǲ5�� ʷ�!�b�Ф�eku�~�};A�?���\S��{��!�����/���vw��Q���XIj����1n뜘�`�"�ry��_��j�"0C�/���{B��"`㛘�v'���^t#�����k���T&��.��Ŵc�ă�-ǝ�������e��S|�v��v�m�[�c�T�)�m�7�>��#kٰ��&z
�����-�� I'׹���1|֏s�=�W��A��<^f����mB��JA���J��ЗE��g��q-DaL2g_��i�Ѵ3��j��rP�<P8�L����1�7f�TM�&��V5�B}c��r��х���A4�I2v��\۝�*ثuF�⦷-�|>A]X��2��r?s������}��2�ｷ*W\�w%�yr������+�4A�]�h�moJ�%�1h�+�%L.U�hfe��¨��A���ƭo��H�b��D������1|���#�u�WE�.�ܶ�f�2�5rv��C/N��빍��=Ռ��rَ8&��f��ݟ�}	I "HA"A$� � ���2�N����ޢ�ć��K	n[s�e�ʺ{c �z|��T��h�f�[�Ύ2���8�S�u܉��L�G7���U������TS�������ȶ�^���H1�Y&E*c�=�S�I�r�5k7p��^K6��}��>ޥI�h��QzH�!����|�����@<U	a"Ɇ�ـ��od2tq�#F��k�e;���vT��`r�d]g�������<������z����/�$�wh&����A�p4��dh;���5"7�CQͪL(�.yn�r���),a��6�BO�ǧ�t���M20���5�P �� `��" ��%�]T�f���d�,!�Z4�
�:���/ֿ<�?pEk��<j��+A=@��t�~!i�����cNJ����˰�W�u���B7W�;������)�zhO�[Bu��;�`�8?��j�L������_/��/ws)��,ի.�j�Ul�k�C��5-�^�Yr��x������C����la�q.j���(`�x�.�L3n���v�����Y�&�ߊ�c�@��i��Ƈ@�r����{���嚺O͑����4�SBw��w]�孝��Weq]%L�{��^8;�ѯp��ͭ'0�k=1�p���TM�\��r��n=/:�i�Z�O+�`�&�̔򨨊��k��W(���N�~Cgw>�8�<�a]��o~��~�����@��$�D�0��FBII	���p�K9&C*�?�,��0��0i�`̖`��LH́��� �5l����;fW���[&����^(�\�b,'�"Eܤna��4�*߸��+��8/�I�[/��s �J����2�=�֝��=:��60�@�D ��yH��;EeÅqt�]d��{<mi-�Yhf�Fd��K�Uv�r3���q�^��,��?�84G���z.��z��-�.�X}�ꪖ-A��M�=�2�]"Q�np5ߺ#0Ϭ�h�����I�.u�3��z:3tV�~�B1�L�#���v�-�P�ce�(X�����o���7�z�Dn�������]+&	d��naƄ`� ��5�ze'XĲ.�<�K��l��Sze�u���Q3(�����H1�l�X.xb���D����]0�U+���^d�p�!������@�mVԖ�vTr��2����
��}m� &���l5u��$K�#1;�s�H���ok1�U{��ƒ~n��Q��J"	� �0��
lh��~��)�_+�}�m��,�e�r��ۃ+Y`�Ѝ�ʕs�"��fS��v���/+I����i����m�X2����<%����4�h:�����sՂ�&�X0��������}��p*�M�IEvn���ǽ)��e�L��ަ)����@	�0� ����J0$��	$�#�<��Uړ���`I�!Cl͸�K���'�=*F鐭Ʒ4g�nt�`���E麕F�7m��1�W�ķuJ��a�	&��a酱~*	{��^~>���TB�p���As��J���w�_~��� ��q�4Nڂ�G�Ye�UceO�/�z��s��}R͗��G�Qnꮍ;�j�;J�@f|�ĳ�9���\����h7?���-�8ȄZ��am��0�6)yaM�i�[�s�.������C��{���E���UL�0e
M��l�.8�>��D	p�}6=[pfmዠ����-���#"ٛ�V	C���P�Z�[Of��B�n�K4O��0��B��m��6a�a�A��sKe߃%��e˟���sU�����}:�=��]K5�;(1�jq�j�G(=���6f��Ia7�W���7j������A�1��s�@�h�y��%6X�(2j������q3���� ޻[,��*Ŭ�*���Iq��\X�ar"!�[ ���j�k�~��xD�NiX5l���9������U��B�����{n�Q��+b��m��ѽc^���btSF�����e��n�ޯ5�w�d��j���;m��2�U�����HIÍf�q��u��jʄ�Z�L2��K�K���z�����^[���s�~@�~�DBF@"!!�#"�<��<<<���|�*e�uʶτB##Z��1�A��		�@��,�>�L
��V���G^N�zNٔf2�s���l�����&��ܞj|��U��`�ơ*��jc�)��`��[������H�wvp0ըÅ�����b)9X�"� �����=�k>9a��:?��t��R�H��^�k6��C]\cO?gD2�	��(���̤����F%�����E�-�
!�m�H������m�s!����О٦�����"�J,61�^J	z�d��#�Ii��78꩒e��Ȕ����e,qP��0�S#
�[gϻ4՚�jZ�&���2�yUSf��c��S����$O��5������`9l+��-��:��<s���Z�mId��] ���!����/
�L��/��=ȂF��g����֜�d��gH|�]�L������Lb�#n��)��:�C�E���и�c����9��fbǀ�f�N6�w�!�W�(>��${���噢�G�ش�Ѓ��1_�է�I�g�����߯��y�S-.�F�bm�����3�bٔrf2s��h��y�iйR[I��+T�>�.�X��:�#�SF��}]�Ɓ���#�u~D4�R���3/��`�5&+霓����s��\���`-��1��d�wlZ�m<�(0�^����y�ׯ/��{����$	�$$A$A� �!@�����S䫮[�%�>ؘ��u��^Y�;�%;�%8�5r2�"ȍlNK�}�]wx�g��k����^���Pa��L��f������6�厐"{!-@�C$b��jw+���.���AZ�E��-��$�D]Xu�<��� ���e� ����!��na���7��0
�����4��8�|ʄm��^�zr��3 �W	"`�r�Z�[ɥ�֒?^z{0??l�c����F�0pރ�\估-�L�(TXSP]s�����ؼ��<✤[wh��r�踇R2�"�9��i����Z� �Of"S�IP��
��O",����H0�$s�l8�vԵ���u�)t�ݤ�A͆��͡�L;oJ�� ^b�7H���@�t_�a���3li	���7�[�� �`�i�`�:�P,s�΁,�5�0S�(�[=%z|�Aj;F��C^���CM�^&ɘ��(�m�$c�@@���ˌ��u� �_Ja=z!q������N1u�'H��๛T4�kjG�rFY6X5�``y���xߠ�1�5>�~_a��~3���^\CsC�������t�'l��;l��Q��7���gB!��{�^�3x٘1ӝ%���������u�]28���ͤ
�A���n���,ν���r������m���5u��3���į뙷Z�Y�5Y	���)�:wv!�C���� d�#I 2I�H�a$�o��׾���u�}�~}ݍn�T���Tq�4Aa�p8z��?��s5Uo���:�
J��=�uۇk�e�6�jeҵ���'�H�i�@��k�C���n�<���&��`�G�`
u�L3vڔ�[}�Ug�V�������A�* yX+�z��Q�ڍ�kʣa!�B�t(>0)U�\d��۵��=�;ם��7�C��7�lP��l���������e��Y\��OG1'�ϒ/��ਖ਼�Φa9�z� ����&��mOH�%@�ټX��W�R9⋲�c���"C�ić̊F���e�k�[��4l^�,٭�yG#/P،�
ŕj�H��O�6�5{�.P�x���Xt�L3*�̾����i�HD9��jv�f�mŭ��>�u���|�H�ĩ,�O�� 5�y���~8f�J��k�@MUq�J��9Ɵ�!6�0ŷ��M�\@L��*��vP�=;�^f��zM1n̮�.����;e���{{H��ʰD���ê=c�4����8�"��G0LW(�|����P��F���g�I:�7B�ELY|ݗ�Q�wtV��h�]�Y'�k{x��59��`e�6bn�n�ے��;-�r�A��-�Z6�S--��vl���s>��4х��UK��P�]�����h�rL�\��}J���Les��s�tg;y�usw����$�<�b���w� `!]���n�+��1�����5P�k-$�_mi�1`�;E���g�:c�V���`�/B*�r���+�����d�6�c�h�Q���,�����Wn��E�ș��(K��Ҟ|1�}.HŌ9��'���6l���d��$Tz�g�v��]Mn%����5.��L�N[�ut�y��5���c�ի9y����zb¥�8��t 9hc�U�����sz)e��1,���vu�|�;�*�e4�9��=J�)%/�������hW�b�eco����dM�A���(���9Էt-����9g<C�S��^w���(����i�6*�.�Y"Qp�<��$�HJ�v�V.��\�˹ɣ����%���4�๩�5�PX���}z�e�结��(k���t}��I�Q9����,�ƚ56�ZF��?-�>ީy���0�R�de�ы�b��K���3^�ݼ���ɝ�]:�]�IMf���f­`��\���zQ)'H��m�n���^X�6]�A*����K��{��o_{h⧵�0�B\�wԞ�4ְl���}��ܔlF�ƻ����LU�8��a�8@�HPs`�w`��%t{FJ*�d��>X\Й��q������&u��"N��L��GmJC��B�XFU:�ݤ�\Z,�Jfn6n�KL���T��t���-Ბ�
r�v�T�	��SW�vv���c�ɋ�'��.=�����)����㸭�5��!Y$&r�\����Z��^X.�7�&�N"�!-^,�Ǭ,$���۠Fi�{J�?))��i]����l&�n�j=���wm��u��1>�	���ݏv��՘�؀0F�h[��NoI
}��������zM+2>s�_:�Ob�lY��9�H�2��+�Mg3��[Ub�/3�o8��@tb��qM���	�Ȋfn���wz�=΁�ti&i��u�e�1�}�]���OX-A��P��ЋΩAR��"��nڡ��A�����e�����ΪD�cع�z0̮�eE6�OT�LL$���'7[�؄�90�G�W�a�V�_5�:�s<яS�7B�ܮ�.��F�p#���7V�V��f@�1��h�O� �	�u+9���r�(�NJv3����������\�|	
m!��ѫ:
攳V���n�'�x�9B]F�l��xZ�k�,�I%�[��Vfp�l�C�c��ƭ9�r�ٰ`�{t[�}�Rɔ^QN4̎�����w\6Z�w��HD��(�sR�jqo���V�I$��{�^ϱ���6E'�K�MF�Mڑ�0���U
$��,�z�p4q�u�b"ŋ&ҢcI����1U��bhϖŊbŌQ�B�:t�8N<�(p�qV�c�Aa�LU �giQ��5baӧN�+X�g;J�bn�USZ�6�AB�wf*���ڣ;k�.����
S�f�Y�lT�$X*��Ne1�dV���A�*�*��b0Mxxl�x�f�jE��-db*���*,�Qj6��e��dU���"�;0٣�Óhi���������@�oVb���.KM֊���
��:S�8rlTb�)1H�**��ݢ��4�#���-�*��ç� m�b �	~:N3hx�i�Q&�̪("B�,wJȠ�У:S�GNgmb)�,_bL�ŀ��
�Z��U
��
�b"��T���p[OS��V,Z�"�,X,ݢ�SXX�x�#��$�PSw�Z�5�hwԣ���j�G!Թ�L���g2)oO]7��&�Ǣ��B�fen1�Z�g3�����9ɓ�4�E@�P�A�Tm���ĒJ�����i�B����$	$�!$D� �$�ߝ�{��~}�ҝX�T��J2��N��I�(���!�	��@Hƽ���\�T�<�tS��9����8��q��Z:�A�_ n��f�1�̜��#�U�x��B~��K�����c�/�W#f����5�:պ[h��i��u��ۼ�'��6&ZP͍>���L�7ƅ�7Z+e�6����zSp��]�5�oUt�z���B>��O��s'/����ؼ���[��}5��s]��z}�+xt��M@q��	���h�2�j;��ҡ����q����a��� �}�67nß ��$M7tt��\�V0�]+���f	O�T�6O��с'��$٪����������~�Y�֯<-�f�b���M���M�У�fw�Z�<I�s�VC���9ל����3{Vņv2z2��0��PY�����X덎>})�\�8Á��)�,Zo1���Q��P�A�HM�eAݬ��~XP�o���ƠՔ�n�m��X�Nޚ��oG+y�XC.�����D��v�_E����އ�y�id0�[�,�r��B/^}���ߤ_k�A���>���Z����:�/Gю63a�2����F��8o�/��x��T���`Y��C]W�*��@완.]�z��q�tN�����r�ԟ,���-bٓm�m�x�UT�+�����f�Y:Q��>�����`H� �0$D�a F��"0�)	�����<S�h˛푍�nu3Od&�VPB�}<�S�쿕r���T)���k�������,"6��˝�k'��7@Lǡ̋��J�k��2�����C6s��cռ&,0��@λ�FU"8�fL-�����
}
o�|1���׳8�� ݶ�i�W8��a�CԖ���Tí����dQ�\!�.ň�q �󚣨5Qj�sJ����>�?n�P�B3We��<��q�����M��i�i�<bM�9��!�8��������܍Һ��V�L�u�W6�OF���
�Y%КX�>���!������N�|ʩ%x7H#f�EY\3K�z���0՗='Ǩ�O�"����)R����az|�>�p�a>A��vمgD�f�1-�t��VL���P�&����0�]1��1i�g�h�K�P	L�	=�-�v���D�l,�ܾ-�Ac0�և<�xn�^���͋i�u��9H��6�:L���gr�������'�z������A���0�τ;" �	�Z�&�g������'�b2tdS�2��ء��tِ�d�$�7x!dnA�Nm�*V:]����%giՇ]���حd��;.cv��,��K����/�}<�˘Y~�qeU�Hxs5kk��
���:[������Q��Z���8k��Zk0LR]���Z{�dN�ǆ�oA�������(}�� #$�0$X#!`A=���x�0����6�^��fA/N��c��u��;�<尮2 ��+,u�����;j*�#M-E�T�YCU�VX�4��dl[k���:�/��sC�k�>�����m�{��N�vh�Ʈ�ùЎC��87�Fi�-���><)x��HiE`ZQ�0|�M	wcϬ�"͊&�c�7v�a�5���A�����ޕ�k����>П�ܥ���`�/��Ϊd+��d�٧�DI��J�c���ɋl��fό�a�4	��j	E����Q��nF�m���e��󵽨��. �0c�{`朊=ƽSQ���p�m�Z��A�JW��^#[�c��N/���:_�V[�ﱋ+�6(�9�G�:GC��,ӎ��y�Zx@Q�Q�ժ1�Bk"�_gO&7t��}�~�h��Xhe;k�A�l|>c&E�<ah[ɖXhlS��MVD,��&-��(s���47�QUiH�AL�	j]s�Bm��!Ռ�g�H[��A�f1R
���[�R�w��YU�6����wL��w�]RJ����N*�}�d+~�W��}g�*Qx�ۋ�ռ�+���n��S�gk�:9��[��a��5`�L�sK���l�������A�[�<��iZ��e��>Xܬ鰪_b\��u��WD�ǽ�6ݗ����ۡ�3�q�5��!V.�3��C2��+t�s����!��ڛ��>�� F�$ � # � ��߿>7ϯ�<�~}2��"�l�9ˀ����@ު����LU�H�����'X�S���Sa�̺:��_e�V����8!��t�LhC��@�T;COeIO\��H09��dCu��o!Uٴ�nd\!�j'�71�`�L���s��|f#�#z�4)0�;+Ľ��Y��k�Ze�oZ�݆�=Rb���.�rC��� �6�w	���1�>�	�S�����休��y�������h��Z��3�M#|�֚�h'�W�����1�4�+����*4�b#���H�)��ȭ^u'\u��Jً�����Q@��-�6���(����I\G���:jK����@|$B��n,5�a*��]5�|��s��sh8:F-a<f��]k��ܷ��0�AV0bUȓZ3!�#�N�a`��
�n��N7��n�&2_G>�.���!kb��Xُf��0�1 �����4!��?z��C���z!�bԕ`YN�ؾ��.��h˴�ly��3�0%���p����fZc.-�x%�Xٰ]�ta�G����ޙ9���G�����g��F���nڼ��);��Ƈ����g^��f�S8��!�=�k��a����N��
U�^��IUd�-a`{�1��}5��Q�61����8d�x[�4S�Ȝ�u�A�f��N�b�d�q&�}Y�}f����? F�d��� " #$��'�>����>����u�h�0*�73]!��4s�p��1�|��F�ӕ��<�C$G=TO�V��etg"�]/m�=R��L ���R̡F�Ty�׶GU��&b��ıH8�-�����Y�J�peҘc!CIz�3�VOT�j��8�L��.���!�=;��4��Pz�jlږ�1w{*w��>��9��>T3*�@/+�4��<����6^%:J�T-�a,��.�'1����=�9e��$��0�>ӼH�8Ǩ�'6}�ǹ��>ڎ��֗W����)o���ӈ:�W���?<�������E�z_'�c�����\�.�0]&�/����8)��6bX�v��x��-N�٩���GM�0u�kg;"i�JX���j�ۓ�	�jv�I�jI��qGƾB$�X[���:jw�t�����܎o���5�zT��	�c=�'�=H�*����H9d�����Պ�f�3a�S��#�]�d���:�E�����|PmE��u	�o��]�e�X�C�çLy�u(:�=��V�#s7�\�`�,֝�T:�Yjݶ��:3ٙZʮ��&�1�w���{7]j���8RY�r�
��t����]-e����29���|-s�����ɰ昆���J�n젮=���	?H�!��a$��]��oߟ~}�����	!�X�
q�尦,͔job�S���5���fh>����E�Z�F2�^�0���a�(�ǂp_�x�1'N-��t���=[������+^&ﻡ��}t�"�P����ź��v�'<����&4R��^�VV�f]^5��ª�ug�Ks�Hﻧ�a�O�Ex�S���-����/�&��-,����j7��]
��l�_(m���y��v����i�vJ`h���RR
�*�-35B����.�����g��wX�Ml����de:�����nE��J��� �����$P~ޝ��Mc��ϧ��
:Yݻ�j��"�{5O}�$��E3������u�-�>���^�ɸRQ(���t��1v��[���
�W����dQ�x".�<0���1d���ZN����6�`��"�rk�7j�����r
z@�	����_0�+I�c⼉�?�����즊�Y�iy�eqU�N���W�>��)͕ S*	Mmq�"@�9.��0� �Ƒ
噰��v�z��s�<D�ڳs�1����4�0+z�*��**�y2cM9[���9���`��s�s��N�#��I��CqY]��Սz䪙}��٪��	�e-1�`�ݴjY�B�͛�(�Ϋ�̩�"�/��#1�ҏ�hLJ򸷟�}��_����FD`#$���H����b�8R��gòzH�I>��Y��6եVÚ��=/�l:��k4�\m9�Nիr���cCl�Ȕ��!�_Ae\����R9�f�^=4®	��1i�4��{����2�����|hti��oD�Wfș녦)8	�C��}��,L4��2��4��tܶ^a9"��ʞذq��/6�׏z��j��� ����{��2n�m�j0Ů�۪�����8����ڏ?�Q���%� �8DyF���U����4-wm��E�E8��|��5R�Fx{���O�C(�~Ǣ�<wB�����������~/�����������ՊJpl2��0�ɠm��δ�;G�}Ɓ#P.�:��mU%�h*v��Yw-��T$:'��e��š=�Q~ѳמ5�Oa`�߯�,���z��J��U�T�&�U����6�a���.��� q��o��̀��/�Jޓ����H�ơ�D�]S��v��e���5	�x�<����a�$O��>ƲǙaQ鱙8��q�vAX�V(k��\x��ܙ�v�)�ݔB�2�,x%��U�r�n�1p��=w�*gwn��7p�&�n~)�����N��8��ݞ{�[:>T�*C��N�<�͢к�������V8#�M���^DX�'c�l�M����6_s��'�"$�$�!"B""d!���y��~k�w��������)�u�1GZ	���(�y�Q�֢��,��%@�һ'�>
��ټ0��Y��:8���-�!l��=���`���]Xs�@|���~3�l��߷L��+���41öP�~�֧L�(��Q�}sEMX�YO��]�4��3%���7rL��/�Z+`h��M�>�t��;�)%p��q�Q��j�w�M�n̞���n�6�B��G����~�V�7���*�,/1V�"����Ոʥ8`��[��uB%����i@��v)�	��y��,k��4{mT�!�ϡ�����^N
���xAk6!�����]WŘ7h�Kǟ �M��P�j���Ү��Fe�@��fq�h�v���N����Yv.He�� �1���6i�A�+�cC�G��A���(����g������t��c��d��W�:g*A<@��
��P.�����?a�_���|
�*`st�T,ߜ��z9O���ң�`��c��3�A �7�n���T1[�����if$7e2��&��Y���7QY��u�������b���ʘK���f��qۚ�yq Q��0"�J�&�n����O�+*��3]奃���a�o��y����|��\���U$�fJ�XFٻf�{���1�iJ>�k5���6���ф�"����# " ^y��}�����ܢ�i�(2]V���s� :�verf�LXҲ��2�{��UK�-�i�LsatN��`��@J���p�*����s>];N�P�'�<tOY��s���K��5wgÜ�ૃ�^,xߴ�(q�hj�(3N�ޭ�'�ݖ��c�r�y�	f�s�T7__/�P+�\ph]�[�j^K�͸f>C�Dx ��G��#0f�;5�e,�cU���\���Z��Ҧ�9`�/m��#��But���(����1�yg����d�Mv�q:�b����L亻+�.#�#na���u@Xk��e>Wt=��ȶ�^�宫M�n�S�n��t�%����X2/^�uɆ��%6_	���'�]�����x�������Nf���X^
q�>/l|���p��i��;�W�����%:���	���P��YIh�9]� �[h4���]��LQ�4L��p7>��������؄�����w=���1����Җ�+بE7%И6�N���C�5�NSz�Ep��| �︯MB���VY�6�vTǩ���i3�Ԣ���d}�iO�{� V���k)C�92�]u�:��SU�:�)�EWˍH����fv��!�d��;�����V��4p�wH�e��_#Ǖ�����}�������j���y��F2�"@Ff�0oy��n���$�Z�?��\��T:◛^YM�����y���\�gA;5��>�M��x\��3��!�CR��la!xp����='�A(,hj��ZB"p��?�iqȃ,wu�9��@�Ce�&�x���XsP�YB�F^���1A*�AH��9���<�uX�jXEsA��a��0gV#Xd���*�jDd�e>}٬"�uB�\����(�W�L6���5V#Z&ޥ�3N*!n2	��a���(���D��c/�2;�H:���Ųf�;�ì�{"���J��e�a��[p�i���Ɯ�_���c��#qވ��3z1�U,i�Fߗ��Mn����<s�4_�s�M�"ƅ�B>�����f�7m��>�M�����X�<ӽ��	�=N�c����QkbY���6p�r�e���݌��Ps���q���FEŁ�^���f��,���S�	�1�ʇV�\%�z��>U{[��=��ʁig���j�]��~����*f8�1������`{�q��<�Eߛ_��O	�=��5ó��j:��n��� �W�F9���1�eiΌ��쭱Ћ�[���1�vA�oB�n��,��6n�[�rm�F&|��X����2�ޑ�)}ٲl7�jS:�sM�%4�+�T[���tC�*��)^>[SrM�bTkw��:vk[V�*ͫ��&R���.��v��X9�`�"�t�2S����o�!����l�)ɣ�i��)6	��1�b[��w1;�x�(���R�J�g2i���A[�
E�4�f_q��P2��N���A�u��v�4�Y%n����Q7�s2�^���Ҳ����YB<��9Q�.qCY/;4��ٺ���ͧ��!u�[�0���B}�oK.V�K���oeHn��B zf��ȭ�Uy���T;�ZXcFSu=��"�[�e����}�gʭ��L�PR}h�m �tQK鎹�W�t��(tf�MV���*�ɔfSq�Л��,}���R��6fb��P���6������ᬭ7۝����qv3�6'Yx�H�*�U����n����Sj,��Բ�6�>�V�;��<P��f�xhk{��� ��b@� �U&U+p0{m3ٌѫ���!�_[�du��֞VQYv����[�-�����5�5�L����n��^q�z�*�Q:�;7k^ЙjYd<�Vd7i���T�W��xw&0w�e�}���,|]�' +��n��S��r�@pY����S�[G�g���<>l����9D��`p�U������;�p1��Sz�V�����1gMU�] n�nP���0"9�ʣk��\�}��W@d�7վ�u�rc�8:���nocn�=}�Z�K�ts�h�cj�	�7n���ɼ.�P&�2�AXg7�n�&v����1���� 3.�[=�r	���qcs+F��a!�ք5n�)�cM[�	b�5JíB��
����椸:��9�&�c�;��GV]���i�X5�wjQrHjc͋(mp��7�.�ef�U";�UF�g��m;wT����]����D\�o"����`�q�H�8IƬo4X��.���VR.+<s�G���{51������V�Cbtc���]�����0W嗙G��83�=L�rV�V��٧�XvX�'�o
w����؆�;ͯZ9�>�u�\���mZ��Gj�Ob0^�Po:�`7zp�2lyU�s����!S&�c�{��C}�*���XwV�ݨ�kk�r�j�64.��Y^Ac�`�V����y�յ#����!�m�[�L������l�rb�����u��9R�:�w�e�;ZFuώXēotڏraF�]��ŝ�.P��Ш��m7��,	űpbIU�I$�Aܛy�\I���ZC��cQA�e��ݳHjЍ���V�f%t��(�5���ڢ����m��X1QEY4��U�VZUGt��W�DV�xp���É*UDW���4��
@X�"A�J���Ç ⡶T�Q�A�F�D��iZ�A`��j��PV�`,O�<8ruӞU
�������EI�AQk��ձAb��m+��'�M�8*J��1G�G���1��
մ�|t2���dȕ"IU(�T�gN8�Zx�-�X�au�"��j��h9k�K���ډbDTE�V4���6��	�g�M<�+4�n� {IF=e�"�dU"�"��]F1�S�ueO�3
��zl����Ŵ�.�,����lX(.[*m'Y�
¦!,jT1����SIPP1�.�(b(�0*T��(1��(�+9�
�?����a���A*�G����h�}]ز���*��Fd<uT�YWՎUP�"6ř�S���9HmE�X#��?RD�!$F�1��`��ǊB�dJ����ߞ2)����K����M�&1�ظ�M�A���jԾ'��������V��Ai�aJGEY�Y�.��,��0��i�C�^@�l�����:,Q���0���*��q�]��	tK*S�%s3?0��<Ŋ0�K�����S�t�OD�Qy�*R�@��X7Pm�����$�D�6T�eA#I��n{�.WG��m��9��έ���RfP�dWK0�����RO� �V�"�y*��Laz��y��;@m�f�,���+���`�@t�cSd^Ȕ�ئnDI��NS�������.�k�Wz�D���6fak/]����郄�C�Ab�qϣ:k��j�G!s�(	�<��0IjT%�՞־���͉�Q�C�Ë���z�]�c��(�ޯ�	����W�\�<9�O�6���g�����*h��cx�yTy��׆If�e�p6���`�]�{l��j��^d�Ҙ�ZD��(dO0��Yk�=>�1��/��ЄwQA����s��ޡ���+�toQ���9�<Y���A�\X�vg�Z�$.�o�l����u���=��(�B���1�F�3�X�Y*������nъ�jWYDG���jٛgv%r�S�#�kV�X������Y�ߣ���s}(�I�$F��ż7��{��[Aa]j%��m|�2���"�P	�V���������^7�a ��M����]����v^���ۘq��d���ގ�Ŏ1����-�y�Ȏ���d�)�ل�^�wV�S;ς�1�&�΅:hx}F\�R=W�'�*�dD��ii�Pl���D��	̅�w��iy�[����yU���#C�4�ˍL�zpfE6,~��䞍�%6�q���]��O��V�He��VE2��)�1�IP��#�w�za^��	U3�O�]��B��jba�qkw?s�v��%�լ��c��T<���r��@y�,v]���'>^O���}3��z�F�����ܨs�c��	��"WzUs
j�ec_H��3�4�5HsO����M;e��,o)~��!��v�{�m�7������I*
��%8���a�5)emΊ���r$gkEؠ������R\3 ����b}|f�PޣI�x	�K��Ꮁ��i������v�>���<��I�.�ۇCC�C���8ᦴ�eco��n���f����{�X�����j���=�<�}���d�Vu�O3��yKZ��}9�@��������1@�K���o>�*X��z��K�Lu��M<�M�r�j��f�b0��Ky+���3x ����SC2�;1͝��W9y�7�=��{�妇�qu�4�C�`�� ��"1b1C��p�l$�hn&`3D4��X�o�2���t�#�'L����
�9��L�
m�/�
=zC(��/���6�"v�aH^�醚�ƂO��1t�rC�3��_H|w�ދ`�
�z�Ř/H�".o$vtm��J�½k��ʩ�o��3�*Aa���ݭGPȴ��A9aC� ��Lm�^�W��N8�ǥk��1��A��GF[&�u#{yCSKt���]ɛ��b&V���ܠt<ମAﾃ��JǿrBEm��X��,7����9�TTԺ�g�=����郂�t}�!ْ|ǐK��h�ۨD��w��(�aEa�`yn�k�b�0JC�9�^��)ۿA�����>Φ�J�DgwpV�]�:�A��׹@!��K�0:Ø1�/�l�js����E#g3v(/K8Z�,�ᱡ��� ;#j�0��܅ƅ+�����Q�)�\G���������Ikϯ?~2�"N��L�A�x��\R2�0j
�C�eAg�(8��"�m�T9�hKg$�՝��r3��78Gwժ�ZM�;:�����y��"�>[{���qvK�G���\���vt�:j��gZ,fh����Kgo[�zʒ�j3P�-�ǔ�v�C�j�3hUMf�:�4yvW*��s�����۾ַ�o�{�|��Q����y�`�%��,˵K?� kF�i��@��_�jXO����Rm�T�dB�B�ܞ�p�qV�K�<��o	��2���4]�l=��m�D��gO�4m�֐uM;���s!����e�1�,%���U>E�Ɩ:l	4K�"��:!�e	��&�| ���^�Oc9��~<��b���[��]ģ)�?EqR ���Rw�!a�:]��l�.YA�<m�8rͣ7�E�
�0����e^��<�G�A!�����3ε���wa�`�][06����L�;����qOK׹E��JK�Ը��Cڂ�[�9��N۽ɺ�A��ޕ���[
oS�ҟXk`�W"�Ī2��Q�b�����3��G"d_�܆\��&����d���?0���n���C�Z��!��݊ay�G��5ʆƓe���6saB5ݛt��^��!���0���ޜ���m��_W[ky6���դܩ�kˣ���.;��P�0��	CG0�o�}�Ni����#z��[	kg�U���{�s��^R�s�ї9�;���M�*{�||�.-o���*tb�|G��*�Ak7�^�7tG+�v V���*��z��a����k�Ζ`�*�n����º�$�4�M��R�.�Y]%G��η|�x�\+d֟�B�(TX���������?_�}�+������o�����6��~��"�ڇX�g����c��b)@�^��{~s}N��vB�t�6��ݠ�#:��4�{z	
���O��|tR���k�*�Y�H��6���ǰIf���`���9C�kO|�KսͯE��3MoIa��VPB�Iw-W�p�*��nv�ٗ����6��˟�*Qxo�Øa[�.��|��rT�G!4
�`[��l?6+��a��,�<r�Ϸ�޾��=Fd���:�R.����)�ߧ"�+��ة��e'���wwxLnl�D��r��z/�ȫ/&}E����H�d;���n@[5 ���i!SdY�3s9ɋ�,�pay�)s�%�
6������-LTp�- �������jյ��m�����7��/U� Wh�� �H׹�6
�̒2����wd\:�ty¿bQ��M��<�{`_P6^�'�:�+�`�rzOuI���[t�T�sj&0���/���(f���z�y�����p:�BCdY8϶�;E�R45P�G����{��]�Ǟ�q!����.6&�N-��n�[ћ:�_n�V=�������r��N��T�d�,	�����d�2���\���Y�H,�B��Lca�ks�s�v(@�F�"�
��ꂴ�C���[v�����e%�2t���N��[�)�Ν�� �Cx3x7��.���F�Uz���a�0��[C(��t3�xމn�;U
�����{�7�d]�8�]� Q.V'�U�ă�i1�D?�1���/ѯ�z�WϘ���{�q��^�j�sOC�H%�4�Zd��t�z!\�*`e�[�63�C�>��;E��yǱL��rnx=���b��/��Xwh�Z�˧�A�i�����;�
Ё�_g]�$0KJz纬5amP�ge�8܋�a��f��ғ�a�M0�M����r�^���5�#6FͥY���%�A�=@>�ߩkC��3 �1�y�F��:��T�N�`T}�.��g�����
v�GZ���e��e]{dN�v�g/6�cd�&����7�DT���,7ʿR���P��$ ]��?�.��ٝӍɭ��my�ml�'b'Ve��e�1d�$�����ٶT:�F�%�s(�y�іJ�'48Y�؜��CqOEco�AO� � �n(2bUN3��q��*��f����O��=�s��5/.UΕ�����l��ګ��Ve�Ot�D4�12���'v��oL���~�#!�j�t�m7v.�����L!ܾ*�> �vH�Qe1W ��^{^�ŕ��v �(� ��Ngʨ���ƽO����.�����y���uLo���V�j:�u��H�b�,s�y��N|��7���ni�s�|"DƻV��-Q����A�=�P�U�B��U�)�\[`ꋇ��4�����f[g�#��6���N���; �6�B$o�������r"���y��x�-ڽԤ�����f{��4�bm ��@�!���7�{�'zU&Y�����܍�NvLt��5��g�s��RU��'���Nn��e�t{hs�sCÖ_1�g�������S�O��p��X�&��0���H\^F�D��Caq�����36�7��p�����ng3��B5_���J�Za���/a(,kQ�a>HB0Ѣ:07�[��
i��x��9E�7of��]z^y���@װ��`��C�#%�~��x���a�
~�=����=���Z�ͦ�"���'���8�
�Vt�T�N8�ǥk�PK�\�����e�VHiЙSD�=%�K톪��c!��pr�feU7:�4�Ԥu[gQN��S��M��l���V�V��'f�^ˀ���'���C�yk�2~�Oٌ��X��6�X�9��Y+EA�w�2�7����f��vӄ~.�b{ǚoA4g�;��=��*����{s�����#��~�(����xg�@�g]�0-�ASem����z�ʆʠ��+�>?Җ<��>��O2�wb=�V����}�h��E�e�$m7��,^������UU
��W����/��wRs��Oi�m������-�5�1���C�?��bBr�^^�sU-.g��+x[�O���`�^��pT>�	�w����;0bt��C 3 \BV`2�bU�t��216Z�p��[�����P�i��yj�u�G+�����@��*�l���&�t����9�b�(��݁ q`��>��qI�\Bۘ���yHZ����2�f�TvoX=�R���ޘ�7����J�<��tS�ŗc���+��u�?k���%6!&Bd�H���TbV٭��H��{�I���v��V����j�!��DD�Ux��;�7!	�Ն��[�E��R�n6Cp�+��l9��r�G��Kt	4K�"�2�n��F+h465N7GWRe����t�Cmr��=�Keǖ���r�L$y�,��u0ha�� o�>�hd���x����i�����9HkB�H��bb�tZt��U$�bAZl����y��pI�Ih�%�vw��_R3�8��������^�5��OJF���PiY�gڞ�֠�� ���ǿ|�������y������)�wO�W�w�f��+r��ދ�&r��Nk~:�6��]���Y�͗E�jꆬeQMڷ�h�1����6bW%B�S�E�umsu�g5˶[IN�$���ѭޡ�>U]
6�X-��O��yC �s����vw���� � �A�������3Ͽ~���~�r�G������\ߦ��sP�YB��z�C7<�#t��	���"���֢�e�
��d���p\p|`��5����vD<5����,�ݚa9��7�ٷ���.�`��s�:��u�]���6,��k(0`�y���(������t5��~�[�K�G��-��4=0�|xr�Y`w�銻ό��&T
=�C�/���޾+q���<Eb��f�n~��w���	���IW߷�G�_�yu�?�����򟳴:<k�4^��_�lbN�����uW�{b�(���#C
����
j�����`bǧ�C�
>�c����lJf��d0x2��bkX�Pp���t��6�"ў��MN���ls�9`�P�H�4�I�_�b-@;	���P�]� !��"	i�[�s3�}܈�\��Y�A��n�
�ij�z�"��c\_���΍,ո0�Z����^��LT�'C�am^�UO�_�t>�|�ߒŸ���E�t��ݣ������pb��Izt�
=�V�n�E��d�,|�0(E����+z������8F�ϡ6hqŶ�'����qR��ï"��d�u���bh2(�v'��b����y}�G�*�&G�j�'�/Oۧ���`rH�����	�e�u�T�eWhw�U)H�EF��*\��|).�E�Ò�Ќ���!&o�����*#"��F�C3X�mD�H5�(�N���!:`��$���d�`)d�F�t�bM�9��ϥ��9
�(��y�⠻^�a��
ˏK�&�x�Gw�	dE����>�t+ݱp�n�ȩ.Éf��\]�лc!�"Y㌷�D9�Ӑ�62�\�ݕ)��r��`J!�~#�b��oguѴ>}�N����tک>�(����~a����}��+!�B3�h�̑�OH�����6��B���O�A,ڄ��E�XX�m�c�����>49�G��,3�-���LB2�:��N��ݭ�h��0����)p~��G	|�OU�Ȇ4c�DF�=�M_T�1�,���*�-�-�m�<D�$d�-t�y�dW��_�-ݛ�O�8���3��n���YVo7)#h�?6ϭ*��3E�S�Z��]>��:�^�N�r�bm�ٲ�UP���N�j��a^�����6�"i��fCra-)�Ͱ�q����sQ~�-�w7�&}���
��S;�V����X|b��8p]���	��3$6��0�5������ h���ř2���&��$�đ���`볕�����̘3>�*��v3����0E��^�]#̾b��ť/����s�k������%�Wӑigv����8�p���=[s;E������->��j���6� ���;�b��l>K�8u��K/qAN��'[	�#-U��;����40Z�`��՜̦��IGnl��ͭ�F�6yst�BdO*����}�/=�9
�m}~�R\�<��>�u4�c<�{b��&���:���S���ُ��5y?%��h�-x�YNtǘ��3	������\�w�%^5By`�,	cFTzLr��ڬ���V`�v������)Mॱk��pi��e[�s&ڮ�.���O�ǩ��u�<�Smˮ�m塗nb,�shmS�m_�w���L�	ݗ@��!h���3�Su	8�^��%�ۜ�qV*�Qθ�R�h��4�jOI䳱�:��[��"�Z]�[�Sӓ��(���+Z-6�F^Y|���Cjd+���OE���C
��V��0�O�5X��*Ì��ື���蹐�=3 ���/V���+0 3aT�fG��W{EP0vPyN�y�+����9�c�g2cw):�0��uӖ�wKF�˖��Ct�rda�f��+��u����3�˼X����Wu��ػ�;Z��n��6�mF�C�:��?%���gf�D���\]C�����S�K�J3CNf=q�x�DP���A�d�l��z��w]Eފ�xs�V^��J����e̛�ip�1���;���($h�Cp��4�`��9.˕B��.��qP뮥�N��X:`���o\����S���Nrop�g$!��ނHg�pU�#*7��p^d}�ʗ�e�Q�� ���_K�5o���Y�^>9K�p�����g�ȆP�������G��8�9��T��7���3Ӹu�&�mŬ&��n���ldK�l�K���]�&��<KeX�wL6:"��ћ��f��y��W�yʆL\��v)�= �����x���b�]����>,�K6'b��ܛ�n2��������3���$�@�z	BV�V×f��R2
׵�|ٻC"vc�Ȝ��<�%ypU�inN�e�e�O���]�����#N	{N�p�e�6����YR�A��JfERDv�o��d��P���s;��DӜ�,�Wj��OF`�S����ê|���n�lv��.��:hR�d]�;3�u\OoENص���L#��*R�Q.�F�dxmR���m�t��2r;���/2�{��oЎ��x�<�^+O5����N��t�ޡr�'��oM!R���yٯM��d�y[8�\�9ި8��e^.��@��M�8 ��\�I#���y�s�;�J��~�2�a�в�qă5.�xP=��&
0?�Xy*��:o �,E4�MG��(�AB#!cn��Hq	Ě`���1��T�x��(\�%̘�m���T�4p���ECC+',�����t���ʪ�c2�Y���M"8��<jc�Z�)Ӈ�8+IP�Q�K��#hT�T�3z��-�K�.i"�J��8�����2W'O8rq/���1�i"�A�[v05hm%C[�!s0�-�s��)=B �N�=<8}x�j�j�8��J�"VVVV�7Hm��Ҥ�i
$R(�4��çR`���%I��|��fe�j��c(�A%E�ڱq�*	���Ç$�����b��`�N!���s)+�TP�Jɻb��S-�edی�f&&<8xp�8���L\����f3M@X�uBT����`��+6��0�w��0�����^2x»2fyv��ʍ�@�x�4���t0�t�
���kA-*V
�2�X)QDE[i�DLd��V�)�ES ���?(}D�	�i���� �ʖ�����{�.�Ej1�g�껶�S��1 �c7[^�:�{���;N��.J�S�l$�6YI��M� �ADA�4�(�&6��
�
R���",F,DPX�����ߞ��ڝOc����UWt�ϼ��>��W��Ó��اր���ԏg�#�u�"äH��Һb�ƨǸ��/����v8��v�i� ���}�(��F�"#�<f\�2���?��ԏ�p?�A��}rg�X����v:[�
�!�0oep�:ㅗG�˛��Ń��38�����4��θ2����Qo6��q�v:�!۹d[��"*\��l�a��AE=�����"�÷c�&6{Nw��΢�u%"UP�aM]�ƷK��ר��Ve�}٭2���d��3��>~�*?�F�8A�><hs��?��N�%A_mje��F���9�e�TI����m�3�ع>�P�b�Q�H�!���17�"w��e���#=��j���\)��exϗoH��Zg�ռ0��"1�vԤ�b` ^l���U�:jK�,��:������{��(�E��	�,�'�'L���\-�� ��m�Dr�O�ò������h�Sy"y4XQ�\��j�I�V:���w$>�0Ai-uSY�B�`�bs�6q�6�cʊ����w8^�s��N`A	���sS�+�e�K(�S��y��J7��u��ޭZ( 5�s+�2��.�,��徍�tK�ݜ�Ҏ��7�u�\I�h%<Ǟ���[4��a1��V�������l��3`��3`0`��+�4��-�a��@�I�K�~�<��qvJ����f�
�����2A���p��ܔe�V�v�]^�����|n�~���jÙ8���~*	{o\��b�c�E(߾�O��~�����@��Lr�Q39�G�D�7U	�����^T�-���s��ͥ�kNI]c�F��t#%�3��%F��`��L4{��fI�fC6\��']���E,�M<�)`�^�Km�q�6�"X��	p�8|��ti�oa&�&�KVW3eUc_qY��k�۴Hw�˙��}�1�1�g{�0{��I��	��1;#����_��ݭ׹S�XBn�Ϡ�i����E�"[��~�Y!�O�6�5t�9��z��!ڦ�M���:�8�X+{��|��۔-�r��� zi+2��T�p�������3ݴ�����E
��/N"7�t[<| [X.[�����H�v��oMY�2�2�/�<]����*�/�p���m�����{b܇�ׄSd������=�y�i&]�C�w��}��:�o�#.�卮���I�YF�f���S,e���5��^�,s������0]H+�W�z��h�[���j�N�s>|��d����MWu���s+4�Q2��ۼT;���V��xX�ң�쭔{=����7f��"��E�Db��ᮞw��_�kg�j�{���:�h;���LQ�4K�ɗ;=ؗ	���v�±#C����aٝ����)��d^��n�2�1E�y�愘�k�~D�f�z!��m5N�ܓ�{F@L�lt*~֑"�����K�ʦQ�>n�eX��߽~������y��!Z���q�^���#�D&509�oz��xi;�8�`���y'����ֳ�F�w�,���K�tdF	��J@����x0/5�%�$h�j��uSs�9��ȭ%Q����(�&��
�w
oG]���A,ڄK����H/��q��a�b���<5��l��DX��=]�q���y�Y��*��\�Ơ�"�s�h����\?	�d9l+v�^��1��Q��iW�ڻoF�b�:������q�s�f�i��v���f#G8.���5�N�8��)�3[-vߓ��C�[�� ��zy� ���.,m��_��:<kl�{^�b�WAٜ�I��顚�� ����m	��K�g��@�Մ3��#�h@28�;I}�΄��}Sn��ã����v��g�-L��v_\tm3���(�g�W\�rD���7�����Mn��9���b��{��ziv�x�F����1��NZp^��VA|;��*I�Z��q�C���H���n]��s��J���ۜm��@z�^���z~�� �"��R��}���~���"s�O\`p�����3�5oF�k�//�M�,:�YA���,�
G`Z���B�zF|�.���3�A�C@A8sOH�C����zhZ��J���w��~#�L���༘*=��ժ�V�V�{܌Fp�� ��El7q�=��<�)�mT�(�[TI�v�g/]�p��������Bh����aD��)\�S���.o���"뽫z��[-�<����/{:ޑ㮂"F��$i.�e^S�&S�ii�p�&��m���B�)�on��!���dz�HBo���~��=��Nl"�P	MmO� ڟuO�:K	�uy�r3��,8O!��-vls��)=�@q�@݅��=�O^qw������_z�1��>y�,�"l?��!��l��c���NvdC�%����w"����Q�z�H-+y�m�)�t����#���^�i��Tޔz��D��M�����i�FV�(^���t��#�u%ٸ�/f��p���6H`V�k�~�|z~u�`���-��_o�.۰���eug!�r�ю<�H"w%�xg-��W�t�6a#{2�2;x��16tg����;Z7~Ug�_d�n�9���G*����� ��\��|�K"�Ev���-gm�8=w׽��}������Y�~",�"�DF(�&�}��ϝ�s���=׸�[�����?�\~���7c�{�D�KcQ���s�z%���8h�#p[	���0�FNmIκ	ܯ9k=�D���ޡ���Y�uy�k,{�}]%?��瀚���	Y�p��؂o0e`�"��Ƈ)���Kq�܁�t�V���ɠrS�c�݃R'i�*����ϖ���	7�e0>�0y�]�r%��^�H����f6m�k�*��l�ǯ9�&Bv�Ac됴�zi��L�C�����F����[����>�O,���-,r'������ځR>��0ya��I�6V9>��,"��{��b�h�m�d.�r=q��u	� ��\3E������u>�g����C��s� �82Rz͌oQ���� �Y%��i=P*%�wN�֩�����վ�{h* �p|���\������S���B���&� �꣕-���f�����L�ע]M3���n����al딑gIT��g8&���ګ;�6�w`�j�l��� #���bs7��J�ɗ�{Vո��P؋����5���3:+�U�«̞w<�g�B����S)��#1݃j��oט�꼁��������{�I�yuz�ζ�56�L+.���>�@P�A�`���7��WE�()}���3�o>_	Mێg�r<$[�B�QZ8Eoq��8V1����fn�0���jT���$L�W]=����t�`�zf��6Q}�Z�0^ql��e8�Ν����-��OO�h�@�*9(kx`�slR��v[P;�{���0h�+ío��]!-�����י�\���22�]d��baY��#��9g���"=kq��үiCN�4۸狜0���"i�&`�a�:��>�4��M��V_�\L�=:�����y�נ�`�Á���Ձz �Gԧ�� j�
�N��<��)3D]U���tf����J�ތ��~�o�W�	¸x萌���)��f�i7^EGHQ�^�qv����*L��u�b`������g@貶=�"{Y����TY=�����[�cז�3O	$�<y��י��0�����,�؅"�`�ˆ��ڐJН5�ֺ�y[�;�+9�]}\d^�]aRdO���ѤD��3���-g�!e��kD������L��c����oLNu�c͢��n)�wS� �u�p��P���9�]��5�#��n���vZ�z�U�[�������Pf�bDg�ˡ�3U}C�<��DMOٗ���4�a��di���{kZ���=�ȹ�c
v�X�U�E���pj����saj*�u��� �;���ٍ]nF��n��>�JE�>��g"�
ߦ:z}�R�FDATz��_f�[U:�l3�t�|�[�LZF@;q^��,*���ʉ��#V`;7������n�.�)�m�͙׉䨉J*�n��L�M3�p�T���u�j�g�{���WV0W���4�_��4�L�Ăʃ�t�ӭ�y<�G-�薻�{t� ��kq�>ck��24��G��7I������5�0�і����&���8 !��~��oA���+bFi��1ݴ�Yݽ�"��*̝xɁ.�-��Q�m�$�F�v�\���bb�ߩ��CI�sz8tԹ�ÚM��i���Cz�y���Pr�V����ZP�p�]�\�z���i2^���U�W$7�M��Y#z���2~��&�w�J��`�ږ��1;�O�p�jF��$���疖���`����c��s�7:��a��%b����l�Y�7{�����?��ꯅ
�oa�����KV��_��'�&c%?��Hn�/���x��G�D�4���Y0,F�kWp�հ.�k�Qyk��h��_�x/邝�(�+��]Z�M�����^m��F�x�����qX�>M�u12p_����E�5��<˘�W�-��k��|,J�0# <+5�z ZU졗�/���	�lA�h��v�M=Ӎж)�m�x@�B�y�QW=^�qW]2�f����a��an��݀�,��[��FK=���F��OV��rC��D�V�<]t�"{a�pf�}K��8ٴ�ܶ��g�n�ĭ�cÂ��U�A��㙫�]��B�$,�H)��ih=y"��!VӴbۮ�ӄ��6����Fp�ofǍ,�؇-�-	t)
:ģ�J�MX�kV<��Uw���E�}0�������0���8��j\��-%�����Q���[�G+�o��9���$n�4�9�me���뼮*�]g&,{�uC]�V�O�N��˓w�gՕ(��=]_�u��V�f%�R>R��A���w�>�l������(t�������-��N��3
z���=���y�uunkYs.k��`�X�Ex]oVN��o��f�!Q<X=d.H��v[�߸@�$:��(���sǇt�J9����Vٹ�3��A�m�>JT8d6c�h!t�T:䎁}
A��Dpk�Ȍ��o0�<�w��W�g*dq^P{�uo��΂�\p�%a�p�5�_5;���xC��n^����QHƄ�`-�C�v"��B��C��L��>�nW�x#8�wLF�����x+]�!b59����F�<�Jɺ���u�����f<�.�q��J��ǩ�]`� ���[����#ь�ۥ����A���0�d:�&ʭ9|������
V�d�e��{�<����7�:�("����4+��鄖kn���'�p��{>V���f֑Uޭ�uO.8!+e��3�b0_G�h�"q�x��iͬs٬v�]҆�\#ى8��g���=z��Q�]Qr������u�m5U�:��F���+V����3 �V5|]��8'z�J�{��u��w�0$�TB���\1VܭخT�Z�S�U�VQ"��kZbtl<ka�o�$8A�$z��3*��;��^�:�sO[[�@�ۭ����3x3�Qį�2���U�qؐ���%Y���:���%i��b��S�߅OA$#~���B��\NB/ ����a|�4
�i=G:LT�bg���Y�k�u3���!C��v1t󐯓z��2�:[�ӳ[��s���}�JNQ���'����K#���>�N�iv�@ɔ��^	����f�a]W���5O��H��%Y���p���(LV�P�U����T5tWT4f�p0�]���}ΑW��2�6vک��?�# :]RC���&�8��ٺ]��Y���,��*�P1'$�T-T�<�NG�cc�,��wb�<��^;�w��:�h(-����z�|�Q��JQЗve�CP}Q"Y�otSrջ�M�K�6˵`�Jc��=uC�r�jGq�Uq���z���%��i}������YϮX8�8am{e�<����n�>ӫ#�P�����8�PE��a�Iw����N�E��fV1�9y�O[��wK�t]��6}}��ܵ�sԦy��PP�U��;�5*�n���2��EvJ��[7�Xs[�n�r��|Q���H�����[�Fcz7e-��X�˧3X�쫼���PZ��1���c}�`�YQ	^ޛ�G����TӼ��	AV&�)]�t�Y���Mևq�b�ula-2�Mv�\l\{��*�7xV�i����Bv�� y^��,��4dp�s)R{7w5+��D
�����&2��^����L�lzHh����bm�}�Vs�wk���y���PlfX�B�n�D���**Lm��&��f�&@4��\�����WfU�i�kε�@ڴ�q���>�εlJ���=S���W�b�u5glK<��d���♖��L�뾷Մ�#њ�P�tͣx��f3�� 5o.�?7Ft�ب.D�K.�)�lu�Tx��c}g:����[k�$�v'\�`:��L�����^�zr��Z�5ٚr�\1��t�Iav���X�\R��1r�6� �4UX�*zQK�e�R�v�1w1\!ȹ+�u1s���r��U��zT��,@⬮��w��n.v��ě(�Un���,h�.�>б\�2��,OXct�ٸ�"��4Z"7x9��vD��y���ў\]ȷG!-K`5k1]CN���ՂDZ��j�o[���$��J�+f�V����B!�N+��.��Mvs:��z�
�j������u[߯�7MTq�c/|_U�㭇*.$�՘�\�ד/�?X�݌<*�6�!wLs��&�R|�]�5z.-q���?�S�$>��-��bm8������X��\ɱ�iwU�{�I��i�i���J�ּ�v��!�{��5�ܳ�E�S�}[�',�R˶��ko�v�F�} �c���Z)=CUb�4���
�77Ewhn�	�����;hܝ�B�]8�u%s�<���)�fh��ybۗ���=�y��
Q�]��e�}Ä��s����O����:��Y8�ro*s�yP�i3�Lp)J��ڝ��
��5�:ɻI�_4Ί�GX�ݹ��V�UB�r����XHԵ����,��\ۗ�w1�����ػ��n��.�k�W��P	2��V�VP�Cd���]�����V^�j�,��`��R���WCa�*Lȍ�p����1��v��-bn����'i׵�(8��Z�%F��Ox�Y&d��L���9�]�֛��aPe��4�f�Q�u���	��X���RlѬ���Ȫr���w<ql���~��!�+5�F��C�e��FP��PzP�9�P7�7;Ra������q__VH�]��"�~B�u7/9RLu��kv�Ǳ�$K2�4��@��C��0v���v�8+��$�G��2)&�wwf�_��,=j((+`�aP^!\g��Y6��&D�������h��P�ysT�
�4��)�`��1�t�Z�jE��t�Ӈ&��kV��=q�.wP��T�\�(�Rc�CF�5�SE�8�ĩQ~8��6zh�����`oUO�.�L`�&g�PY4����`�\0R�C0���([� �h�:p�Á�x�B�i�K���UHm8㧛�b
f�����Z��Hi &8t���x�����i���cRc��b�eW[�3VLG*$ճc&�OOO&���,���-&=��(�(V���Q@Y��n�oE~%�h��V��P�M��6rR�m%TUF,��Ҍ�F���Ub�l�̋*�g���J��Z$6��嫕e�V�l��J�YU�E�W"!�T1��*[E��S�Cq��U@Ŷ
G)��&�i*-,�X�1PQdm*����4�g�ٗ^��g�ˉ�wW
�mIv����2�]�H�"�!UqՄ�*�qݔk��ʭ�{-mD�9�S��4+������0f��I��,������I�͑�ԃ��y�t8��<_r/{��a���Z�f�-�0����X�%~�@ǐ��V�=Eްmt%����ݪ[�����k�B�����o.0w�[�G"|�=t睴��n�S�\u��إ)������?m�m��.6�?{�d��h�g���($-�>Ρ��F0��0+NkT<Ll�́xxD���VD���F��UM8���:�>f*j���
p���!��������ѕ����Bf�0��%��&�S���vH8m�^R��u#e���XE���bUơ��c͵�Hks3ZxMм�\R�	k�#��wj�̊�@�,�i<4��Yr]�S*ʳ�5U���f:|<B����N���r�(T��A��~��ֿn����?����z��߲LIX/�d�qr�����޷ ���%H�l��A~M�j�U ���F�7�A�j��X�z�`��w\ڠx�t�6E�z8�EzN�}��8M��y�D�ف���b����8�4�����.���k�`ɭ�v��;�c�Φ�!ܡ�	wj�?U ��0V�Iew��v�/r��#+�2�����䯕"�7X�CmC���Á�,+�:��U3�X����7�#ek�c�SA��:h��if�i�.��5�y�CC�u33x� N��0�g�d0V�F3r�=���3��y�'�
<�6�@�@.��ݟ+\e�m�f�6HY���M�;癵�e�Y������6�r+h1D�B�����:�?�����dUemmʤo)��q��E��~Q��^��q�z�	�4u>6ѻ��布]u��o�%��/���X}����?W�c��>s�y���S���L8!k����Y��~h�c���<5�������"A �M��ǵbd������X�4`���nK ��p�k�%�o$�_`��	�C�a�2�Hy�'��t�r�-XD��2U��s>�g�B
���Ԍzg����i��ۻ"[��U�3�M�%����mSWZ>��ױf�P�e�{�i��Qe)���%��*��x-P�y�j���M���Zs�oP��zX=U�9!ھ�1.�mu�{��7=��.B	V��q.̾b�ִͧ�Y�2�i�wX{�\�����'�{Ҋ�_��M�G�~33�d%�����8�x����dv���h$q�ٷ5�]^ X���2�Z�
3�޳���Ԫ��.3�z9 ��w�v��i���v�7������,x�B�@:'N��{]#]�2��Jp��X��t޳`���^���Z�����&뽟"�B�����T�������u�vJ�2����7 ]ӝW �:B<�N[�:0oJ^����7�7�A��n�.�L$ϑ�������܃�2���>럄Z�ש��Y��î���5�-n�����c��q�a@n��Au#A�Ґۘ����T����4��+�G?K��f��a����ϖ��>��j��"}}C���X�z.�h~1�P��Z4gC�OqJ�銒����MԚ�%r��8�w���\`��u��Lm���~�'�.��]��Iu"�5������'�^����0���m>�e_G�8���2,�݅ޢ��׸;�I�4�ز�1ۥI�VzҶs�(��2�	w���`t��h� K�NK�B�<��U�A���+������bۃw�u�Rf�wӂzn����c��0`7�`��0�e���T��������С���E���.�1�S�m�Y��/�6%�c�haR�{��d�xj	}a����6b����,�ޔJ!��-��g4����}�t���� �"�G59�d3�b=����)=LR�L���ĳ>�,t���I���o�iց�-W�E�xxϴ0�a^M�D��>nR��w�c(�H=䃗UwT.��� �V��[< X)h��cU�w����3u�ʕt1��4�+����d\�rY]�iJ৶^�u���M��}���\z�#�}T15@�
 ����Y3._9+ܓ#W�g��z�"��7�8������P�:%�Z�=DK\�B+xF��CzsH��Z��7���!$���I�Q�EF���I.B8�N�-�"3��	s5��]�1��0�B*��K����^�23 FR���i��"`_��	YPI�Rf���B��<�8�}r�O�:����Ҫ&�%�#�iΤy���Ƀd�0�����h\������NG�#�Z�o��;�C�,��n#]|{V�� �q��\�%�4�=����u<��s�>����]�_�3�7���_�:)V�^}��GO��4���a%P�+���,�9���L��(�����r��Y�XU�@Y��%0zq��X����T�	0's�{C���y
�sP3318�V�ǘ���:&%H��K
��2�ݪ�]�%:��[2�y�Tp3v<ͤ8���6�!{�a�%�����&�[�=�8{h��$$ξ^$�����n��m�w��g#zb��r.�<�K%�1�H�;��<�tާ����a�@�c�{�l�͡�;���[�:5l�Z��p5�j������MBz����޵�s!���T�{��}��bz����'�]�3o4o8p�OhiPwM�Q��6%Vv����i�δ�8҂65�$(M]*��(G\`eC�R���-�y�F���sgl3즞�\�_��{�$�pb��b%b�l~�{�Uwc���cY#6�G��S-�>!���x��L�|�+�!�Eu�\�g��o;���^�7�\�?���&~�o]�U����U&a�F͔��蛃��u櫜49������6�3)l�}{o*iܭ�9� �UT}B���>NHD�X���O7�6�/-M�:��p��A���,�-���;>P�q�+Q�z�u�۱��X�w�{�.��z�H�g�^�d���;\�n����&�ZwhnAX�2�Y�B�����qkí�Dջ0���G"�"M;�'��*U����лqƽ�)Ra�BQ�*�<x���T��sL����{��w^��ԇ+���Q\Rq<{�N�S��n��b�^���<�i��ή�ɶ<��pY@F��ޓVSA�L�C�h=r��ޖ�z��q�E�|���m���0N5��X�{�w͛�0��9F)ަ�6��ܕ���Q�y't���?�������C�M.�*�n��]y�.ܜT5���U"OC�\����xm���[ʶ�����d5j����VJ��!��h���G�ȏt�������CT���ӳ�'}��/����'��*�@�>ڱvh�{}�~V�	ժ�S�I�K��E���5m��f�.6�Xy��+��:����c/�$���R�:L�Q}:էj�xt��ղP,��E��}Wir�:�)R��	�m����Q���߿W� D`�&���{����<��32�T<��ypΣ�b���e�2�>��2�d���G�Po��}�Q�g��f뾲������h;�#�{A0�����{}�H3U�1�PɄ+�8��� ҄�g򡂲D<�nϸ�k��J��M�ś�{*:�5>D�\vb�����{�@�k���P��ZM� �k�:*�ْ}���6�A���m�i�m��N�t�`����O�"i����Q��=�����B0��A?�GHv����r+�-�ײL.���vÌ�0B�[F!�Vy�����$�(�M������t^M��US�m[�����X�V�^��aFy���X��jwس7g8��a�;T���+UA��7NdmA����
kG.���`F�p[S�̅�7���m�!�z���� 6c��p�Bَ|ׂ��q����\��lmM��S�;T����W�f����5�̺��]m^٣���ڻ2)|�\�����h������R�v���x6��)>���-�9U����@�6���o�[���ͭ{M�Q{٧��̦x)��?=�s[��o�{�w�����)�<d��x��ܡ�Ρ,�Q^R��9��吣ۭ��!���o��̚fn�l��kkD�K����0��g)���(�ϾKv�~,���kI�0ډz�.jk�pO8
�NτF���:�s�Dz�{�B�51�1���O#�X����c��Hj����	�8(ȍ{jÂ���OSYC�uZ��\���SC�`��[���
GPc���?b4 ,��c/R霁�of�N<m�i71+��^���d�Pc�in��hN�Ea�F��5��%���\`���O;0p�6�8��b�$�(�Lq�@@���2��:�8���ُ��\�5T���򅙡���3����׃l\��䡊�\�0�i�/dV��w@�l(jk���W3��$v�H�Ȑ������ID3�q3**Wf��V}���q���u�=B2-rW���&e��l�b�G��Z���:��xI.g")NT�b�wKJZ>��v�n.�s[1�A�V0�U��(X4�)}Om�zl���kuEU-���TuZD.� [
���mھɥR��6�	�g#������\�vi�OrA��^�b)S����x�������B��}.��i����u�;s��/V�4ϙro���v��ْ:i�i� z�HEkR.Y�#(HSQ;��y4�ޮ.��I$+��yT��yrv����	!O���5�l�]�̈�4[���d�^n�>K��6�ϚE3��d�כ��Y����q�؍�m;�BE��çT�/�g�J�5.[ϲz{%��e�e�޺�V-��=L2��%dx�ݏ?l�>��3ֵ�J:�utw&(ٖ=x��b�mK%��z���m;��p�&�T�ܹqj혰k��C孂:z�2p��c���-�����-(u��B���^����f�VH�XwWexq�`	\��M����~ �D1����j�H-V�im�YM��#�+�b(יt�O��}`;�$qȋ�Q�j�w�`v����u�vkU٨��s �~[���xZG�4Z��>N�3c+�uӜ�`��`�`���Lc����@��]7���m�_h�s/�w$;�a���n��a1��a�݄�q4:�m�+�d[V8����.�E���z�z���o�݂!�xҪ�
��Ď�2g�X��f;u��m��Q�e,ח���3�U�1|�X�8�L�H��������3O	$ǈaǚc8*����C�	Iw�sO��� W	+K��D|Ļ`<
I��3 ^>�={Z���Ȩg�������Ji���O�;��>-]�T����#\��m�/?%�os}��Ҷ�x6�R��-�-He���F�D��u�l�#�0+�ե�X���|03�p9}I*�u׀������[8��A,�U��j�>�!�~1����?>�������O%P���ne��T�U�=�i�8M�ڽ-�T�����U���;��Iw�°mD���q�m�\�i�CF�RӼf��r���� u��䢄�b�(�/��/J�C�uB�m�̧�ӱ�F�m��\���̛EHA�pX��/zMYM��=�F��jڷ�椁#՚�$�e{�k�)mT�آ1�-�u=x)��ױD�t{�Y�=��/�H��z���ܢD�ʹ��Ҳ���o�7}�����c�6�0e*��#�:qDe��zy�ыyYq��T��S{�5񏐽�V�:�t���%,dk��x��*�KT�ٶ3��;P��R�T�$�>��&^e��V�bѲ�U(����s#���ʫ(�X�侫���p�;kS��n4�5�=�M����TR���V���
��3����)-��M�m���w&wS���mcm���'y5jU�#��r�R��m��b��&�H��ɰEk�,F��ݣm��e�a$S|�3��A�Wل��m�wJ�43*�!�y�a�E�Һ_'�˾oo�ßa�	7C��E���h�����Yn!ht�������^���y�E`���oL2q���Vo�P�p�v�4���n]i*���Fd�fi�ϯ̄�aʰ�%��Ew�N��ou�h1��Z���l���X������x������'Oq5����@�ʿ�lB����zI�smH�
�p�3�!����Ӛ �H�R�s������E�d�b��C���p��9F����&�R�c��h(���F�L�,���Kz#sGKh�I�۱����!��f��G�����8�V�+M��ڃ��w0�좻n�1J��!'DU�"oq'����)��]�g���w��[|n�XXo���1����̕��a���w�@ޠYb���e�h'$i�t�t�}�8�+r��;���x���\7v��^��r_7�/;xVJ2��qb�ٰt\3i�}�dU(�a)s��a�h�\%�mf��J��OU��[��F�.�Bl.s&�,mup�6ݔyWb�F��foU���r�ڤ6Z�l�1��em�v����*�) FΙR�s�p�b��q�����QZ���0n������2��Ŏ`����� ��=��Դ��]�]]+�]�H��ܕ:�	�j96�i�T�?Ly����Ĩ+�*�W2AK	���c�Ĥ��+�[�K�!ك���#��X�����l���]{����q�L�'%[��
��9��\mS��	�M�S)�ys�jg��1���B6�v�[� ��2�a���՚ޡn�}�������cA�V���*�e.��<}
��܇�g"�(̰�%e^Z���b�-�en�e<ݷ�맠��Wy�,`r�׃���7�mR[~SoE�#\��:��%-��	���DNBwfL�9��Ŏ��m듴P�6��0T.�{�]$��aV�+��o�p�S��|d��AS��rF�i԰����r\ܯ0հlF�e)*M��RsPL,*���k�V���o����@�,�9��.�;�0ʓ.�t��C��ڝĦ���(v�4����2I$�@ne̊D.�����\0<�;�Y	Y/�Ȩ�Js���A ��9���;3�,k�4�wۋ_wS��&j���m��E%>9�e���[[F�(�Y�1jQ�)PX��L4~��e��Yr���B�ѡXylP�R��j�4�!Z��VKhUB�(S8EyF���TX�(�ڬ+*��̆9�f7*#hբ��"��̚q�DM7�O�jT(�kUZ�(��LD�YbZQ���i�5���R(�6xxp���fK[��-4��h�����T��mAHڵJR��(Vu��*�4t�ӆ�Qf�
�"ѝJc|�)��B�T����e�8�c*�k@Gi����m���Ԧ<8rpPQ����lĮ ��b�3[Kh��
""��q��Upa��0�ÇZy�UuJ���Fb5iiq�����AVTD.�1��J[
�Sy�Q��G��s�q
&-jԬR+[�X���E�e2���qh�b#&����5�m�4���*;,/i�9j��UT�)iF�ۍ���R������Z��嗗J�5�>�w�>f֪���sݙ�;�9sM������1d��o-��ǛjQ�2�,�yZu��l�㷃oRZ�7ݚn�%,���(��bI"�?��[M8�6�i�qA$!�����1��� ;��o���8���)UU��%��e��&�N�܌��a]4�~�b��y3�`6z���9;����a��).{�[/$�ύ�(S���TސoD�l��\;�f��gl=�� ζ��mx�p\�'�S�B�v��0���%��]F־�M���+��f�?-��՝
/��ϧ����f���_\��x���I�cO�Fl�p2�e�=���lf�Vii��E�p�&����9ȅ�"�F�mfC�,����l�a�-W��F�O+>�=����%�:���v-ؠJ�u%!棣�.]�s!�t֖�<���ܸ�Һ��t(r-Y*�<��.��q�b�kv���C^��^���x:#��t̪��6D�$CQ�	U�BG}�L�:e�5�V��٧h6�m<�J��^nz-q� ���$��t��T^w=�b��<""n3#!����\��L�?4+�ֶIXװ��[�ŋvM�+1�!*���rM��p�2
Zo4�= &�� kk�s��d��v�ˀ�9��m�̱	i;eh賝�үql�\�xh�Lf:[]��!UW��ttˉJ�z?��yW����U�!���!\��ө�nk�Uq��%*u�p���6�o�̿T�����ndU��^'50�&� _.�k�=,�)�+�Pt��5oy��QS��PK�ώS�jJ��\uX�:A�`'�u��W!�r��p�[܁���#rw{��-��N��p�lǁ��!lB�x�~�9mR����6c�b�ͤt
5r'�t��jJ+�������j����2 ��햶m�4�>۞Py�h?5�N��=���L���"��fB]˱�4����[��C^�5]�w4t�.횠�����B�.�q�]u]�p�]SR�ME�T8��t�d��%����������Ć��	���O�����a6#зx��]��#�:��/+�y���ztuO�n0Fe��sZ�)�����*��,�4�8Cnʯqn�� ���	x?����t�Ů�j\k&�kqM�R�_E������})X�u��W����~������ux��s�/F�d�%wFlm�6&UE��8/Y:ySA$\˂c/�p˒�]WN��`�ѣ�θ�����W�;�%�Ec��5�wt��&:�b��[��#��|�W�4}�/�3����f��Lv�i�q�tQ��/� �xy���h����,Jo3NG]�X�x�h�뵢��$o$$D:ހ9e�b��<j��y&��nФdz,h*C�i�s;wY�#gp ��I�+��5�������Was�?{v��2-?�fce���l��8�|���-�l�U ��>pg�eOiR|'�z���т�V�q�ňQ�s=h����y���4\�����&�^��d���I�t�Ήw���G�����ۍ:ۨ�䆫�}Yz�5�J��	RIK�4�Kn�p�E�4ی����=�d#BН�Ĉ�\^:]��I�L���ml��r�X��$L��*��gR�v7sX����C�ĨC�������`b��M�
T����L�Bx���NL�d�
-8@�\�ly�֮3�|�P8�)J5X��Z�o�.ҭ�_X��w"��%�Tƽ�1��u����	*�!xȒ��̭�R��3u�K�wm�����������j�7S�V=;�ӰB�i�):��Do4����ūN^t��4x6�m��m,��,y3�^&]M���k���9�Pŝ��,Q"�tG0C��3���A,��M�*��l�5�`rWmz �8�=S��>���{��D�M�$w�+v����a��H�a��l;m��3�"°n�L*W\�G�����8��4aӜP�P�t,��6\?�sσ[���2�Q)�x�����:�rRX2���o��;I6�
�"L�ͧ�rs_p=bX��<+5T
�r+	5�L�n��>|�у�%N�����c���C?��Z��nn*ѡ�6/-����D�$���C��C�,x�>�\*=�/�-3����)�@\Q��Ce����{��[7��}�y9����%���)?TxVR�{^K�c����M2�b!�;
�X�m���4���]�����ځ>�fB]myK��F�!��Ō̉I���f��N��2�t٠/PN"�٩)��)\��3j.���[-�2*]32��n�dU�fW;�2kUBUM���<ܖf�֍�dCU��p��3�n<#��=-���P�;w�V�<޹�n�*oM��O�L�63I��-�;�m�j�lNd��13�p�\�l,G�\)Wb���n��t�!3*V�w�aQyvC���Q��C/J��,��~���6/w�;y��0g��T�B
8�p�� �L#D�U�m���7L^:k�����8�n��+�#�$D�89[��;�JN]�,��ז'e��Li��m������%F7�e���МN��k��F�
V�]6�'4�2"�gv�z�,g�̍��u�M�ԡ�vf��nx^���7[��,�����Mnb/w"w�L�E4����w��������'�f��'*�(���y�ɵ�0u��=xn��{h�j�W�h�ͪ:�,:@8�g�r<�
<s'g7�O.�y�@�z�G$��	�En��n�m�u P�pGb�Ou��<|u1��jsP��z:v$,2�KW�W��V)�Pǀ���^Y�#�\+�-{z�S��k!��;/+��8u4a;
|�Q���5؎��˴����@%9�,TC=�#�Ѓpm���0����ҽ��a]T��a��U8r��%��ߺ��`��Oi�6<���>5҉��~Ϲ�˜�x]�٤p�A`�O���V���E�Sf�[
<�&���[�n�7%PA�b��h�NZ�.��m�q�ٚ�u�ۇA4�a{�P�B�6��7���,;�!\ܒ"��bD��d[3�H��-8na�����F�b�E�
�S{6��*$H臙2��
��q����r͌�T�_]2�Pܳ-�z���iP�q�(he>�eZS&��zys4kpp=��B�m��Œ���q+�
���:�]�L'�J�A�=,܎"�#d������(Jy��=�T��l�U@4�زZ�D�-t��tć�̓��e��̅�/+��ȫg��1�w\�VZ����5i��X}g�ּ��CWx�7�x��%�d��M�*3��u9H9ж�vSⓃE�m��f�����O�Ʃ+�\a�hvx��Æ]��!�����[�d�<ܢNr麁xD`��6F�x�oɞ+ܩrtxn<7!n���[u���ܙ�K/Kl�Ї!c\x��Y"#�czz��g`��)n���9�4��/l�n��{q��%��O���5���r���j:�/���;�tX���T+���&�J8��:Ԯȕ*[1�۰&Ȼ�Gx�̴�򆯥�3�Yz�4����q�̧]�GcO�,௘���vW���?n�0�j��o��'brY�����H��>��N�Ȉ��g�tu�w%ޥ��ە���<D�3k�i�w6�B���`��`�f��	6�ҧ�=t�4�g����2�9�m��'�UB��r�H�dm��opF<��נ,T��}�Qpov�'H����}*�;�G�h�Pc�G6�e=Ꝉ(��N��9������ٶ���L��� �x:(�SǀmM>��^�nT��1�\+R6��ly��H�gG���H�$HH�u�ܲ��-�*��Uo"푑hF!a���(^��X"�g.�	��r	VE���&y�FNF���|�$�?P"�T����@%OU=^��ϏV%���nj���|��H�ܑa�S�vS!�2\�
����r(3����n$f0�G]X �ή�y͝l0�C�S��*�i�cٓ�OL���E���(���fvJ��pw���f<��>}�����^�HpN����\��@Z�?f&c���1�=|��d:	�(h���KK�����$�]�@��sYʰh'+���y�y ۹�Z҅s��u7��Ua�)�讶꺭ԣʚ�d}͏� �Z���tf��:�n�J��D�I&;�j0����]�F����$c̡(nT1Vۻ�%�����ЄV��(߹�$,iO�q��[م�I���xOnntD4�F����#�G���6i\-���8
����p�����f��y�0��<�?��OHa��#����YRl�8�Y���\���!���m�1��6�Y"�Zl��+Y���?O[�HA��\��s����"z�h�;�U��[�P9�������ކ���)�W��lFÜ*�8�_Xtq
(�P���V%t-��:�ݤ0��Nia�.�!��}���a݅jqu�Ĩg$i�H�5NW��76�"f�����n�:��b(
��3�k����}ź��a���Rg�y�ۧX�q�t�p�[���H,��U�iy]��tcם`�9�a�N�/������ݐL�,"�I�NZ�&ߘY���v�=�:�����}����3_#�N�������+PI��;u/nd�(&x���	\���Ľ]q��g^���+wke�k�ٙ���wn�^�U��"P܉7�yK.���3�J�D�I_�d�L��;s��P)�`uPTz=��PS�ZA��x�1Y��������j���)�:�7?\���s�0���zI�4�m���E<{M�TH	C_��K)lH�����Ԏ$>ik�r.���w%|�mfĦ���s#HB�`[C�)���Y�燻Lv��5!��{5TdFr
�#�Pz�-���;x�ꝴE�=[��+��@�q�*b����ڂ��F���Z�t}�'����q�h�����h[��g�C&��Eo�H�9��|>�{(W�.LEc��;|<�~ߌٕ�L�!�@�1���Ep]e�z�\]d�Q��u��3#���y���	^�I�-������v���! ��rqfx<ƟC#('���0���������'z�P'�����ǙL���hYkm��T�mJ��[3�'�ub���]1GuE>�4�T��X5�p޺�r��ꑧ/��Ϋ�z}��3��	�W��."E��Z��[hf�sMѫ���&/��.�g4q?��\�V�	BsT���H`�G��h�}�:W~��8��CԉkE�K-qJ�w^�˹NA�|�m�R�*I*s+�w{v75�ɱ�R�����S����[1��6T�ݮ�K8MEJpf,5
�b��GY�t�x�O����������r2���w1ݽ�=A��Qq���|7\���+H[�Ǳ3�	� �>٘
�����R=���D���1ո�ܪ]��F'ͱ��
=�JS�v�
�^�R���˶�S��������QDH$ӭ�Q��~������	���T��æi��i��Q���M&娝�=@�C�l��o�K�ϲ������[�_=�����X9ڨ�L�U��K�BGZ#������.j�ff��p}��Z�c2�s����m�n��N��]���2B�\�AD�6��ih����wg6#bi ���D��!��2��va�Y�@�0��qm�(L��F��4�WDg4g�|v�u[�l�HOx]	R�^�=��6��Ӡ�����%���m��5��soD7�vI��[�lk�0�_`����zt�T��6n��{C=�*���q}I�X��[�B�r��Ҳ�.	4O�/��;9���:�y� J�B�e�+:���&�}#�8]�*�m�����;"�R}i���tV�����;�B%�&�V��ڣ�nnn;���[r�5���C!ˏ�M�vήp�O�\yZ2ĵiv\�:�V��ڸ�[B�P�2N�q5�����P@[Ы�)8e�8]���'#Ͱ�/q
*b�*�v:÷��w�:�YN�6ĕ�y���}&gyQ\Of�B9e���3�6p��y$�6�M�TL9Eq
�'k�&�k)C���r�t�.ud���뻭��N#$�rt�dgv
/J�ج�:�:�V傸 �E�K�����	����'Fd���lx/�>��J���ހ�|��U3�� Z�aћi�v�/+��Yy3����H�q �1���k�����]�w,��"�R����f̪��aF�=��(�ƄǶ%`nF�ϥ���p���h��]�S��U���钭������V����h�89�.��]����Ywl�Pfn�r��W4�K[�R1�wٌAw����FIsOrp7z�\3��fc���7���7I_h�e���*��-�;3k5�ӆ[ړ�] ���.�#3�e��p�v�+�kG����BULd�p� R��a�qe Q��9���Hy������(>�{��Y���#ZS�c0g��0���[�Q���A�3XP��d]o�]ڳ��\E)G���g^Ǯ��ţ�JWvD9�%M�Sk��Z��	9��X��Ւ�A��fJ����p���� �1�eP�.Q\��+���Vp�Ƴ���zNg3�qk�NPmfo#zܺoS�^�4m�̻e��=<qlUd�32)#�8��T�>Ȍ�uV6�]V���:K�ks�OY���+)��o3�a��[ݙ�/��N���\�m^'u-��ob/�n[*���\:���`�.GϹ4492�*�^Ͱk�;�X��+#�{�^ӳ�����)�¸S�s;_:ui�T6,��vN�	v�R�M�an�;�ET���%��E	�9h���{)#�۴	�3�bI|�����jZ�3����i��|�D�[T��xcY�ȹI��7�	���n���W.V�z��6](%�ZWL�Mޒ�h�Qʠc���p��}����,��MtCC2�1���ԙ[w�1��eZzC��	G��̜�U�cu�C\�O�:�s'��z2�rD�R}��>k7"����.��|���o݉�<��C��w��7mWU޹�j�٦�bv7�sD�Wg�8
-b��
')E��`�+Ow �*S�v��}�k¨���y�c;�;}�k:Zז��7m:!�O�3(<�O�Ū�Ӯ�S)�X�i�,��	�����/��I#��̙�Kr��^9��4sOl�]�8%��j*+�m��QDTP��D�4�--��QDDe4h�<8��j*2>U��Ĭ��%TJ��U�8�b ��S-�(Բ�xxxp��NR�PPx�ի#5k1(�*��GѪ�b.c��n�USV���\�pS�:t�80*�����W��'���P�X�����-U"�("�n4�m
���
p�ӧs�chS)b��TƊx˛)�lʅ().eq�X���E���ю4�t�f:p�/(6� ������<i�St��XJ5.!\j(+�`�,FQ%
açNC�`���q�%�Z���n�v�b�{j�b������jcV�����GN��M�ؾY@W��-(�{l]eF.e0�&�LaAխk1�4�"(�ڬ0�GN�'mUEUDE-G�J8[D+�QE�QF*"�*�����,v�TKh֯�3(���V�%���+mPUU�-��m3,F"�*o�]��١Hr�ng�r�,Vވ*�}�Z�g��b<��9<\�嘭T�.���X����l�|��&r���\�o;��#h����Ę��j��SϷ�%gg��15B��6u�i8U�f�q'�al�vs�ޔ��4�=$��'��o�x���D�͘��ǳ���G_��ح�#l�i*4T�[-�yf�O�e8[͙�����ʁ���4u3zO�]
DPP���zz��ɵ�"�F+�w�e�5ÉT*���cꊕ�>3^5�ؼz@s��ƚ�u]�b�s��f�<hGE�=uөTe���a�k�u�S�S���V�D��<�2�90�R�����~�i�_y`X�X-���� )�����,;W`��Ζ�l�]�Y���-�&�1�v��1�}ا{jt���!�W��Es��G�:o��c����������U���LK�}��}{֒�6���Q�Lҍ�*�v��o.�Zwͺ�m��#!�k!�	�Б����.�&T�Ô�tn��2�SL���.y�q�c��z��H��8��>�N?�!X���B=y��.�����|H��K����4_G[�|�W}�X.E]�g"�b�5t"+j����7�y���Otc��:
 yHj2oB77�" ʥIʹ:9�AFŦ*k6��pE�"��}����g�A(z��%]^|{z�j���)B;lc�ۻ��b��M�Ac�q�O(��,��K���gA\X���"�¥��#���"�1!�Cq
�rT慞�^���]�M<X�P\��vT�,��J�;�f���f�;���[�a+S�<j�-h��n�)h��kY�}J��1ˑIXǤ
��"�G���o%�7I���{��NT��.�v2&b�rT吇pyl?y΅�_}��*�J�M����o6��曮��K6�B�u ����2 T��]"Eq��}	<�Xznc�=���K4]T��q@���7y(n��a��}[�x3ߵ\�w���]��C��|��s�G��B�q�HwpY�e���!�65�9��|���u��/c�z��Y�ܬ��Y�7۫���u��2k���},�^�y
�uZ����J��y����kVt�WJ��'AYS������j�Qc���&�x�����zv���-S�W9�;��[���j�-צ�HX������g�Z����Vc���,4�9�^��X�ӊϸ�R�O�d9�;�2�����g%r}_�~���
�����	�ʇjF�.�M�����4b݈�W��<�:L���E�a�z�bX}^��[]��M{��8�Y�j�T۽ ��[A�wg�C���N���Eo�3��Y��F����"���1Xv�ǆ3|4��㊑ظ%��ィ�`�
�(s�\�BXE_�b�\��]HI�+������@v � i��{k��?�,B���B�V�Zk1VK���ut���Tp%��y�][��z��U:��� ��X=�w�� �a}B���d@�!^�J��T,�n�9��ʗ���W��oD��X|����vX\�#Vְot���7��@ڞ��̎Y�����۱e�i �5;P��L��F;��"�"w��җˡ���w��=�c��z1�Z�-yQ=GV]�OFU��KK����uSL�?IhO�>��{��L�9h�֧+;��+
X\S'bg�:���u�W%���_����w�x�O!r��m�B*4�fU��:���G�H�%��N����3���-L���:(�*Z+�<U9�!���b���U�U�{g��K{�[F�a�����6-�S�M���x��	���Ю.aq��F̽q.ǆ����5�%����"��K�-Ҍ���a\�g��=�ɜ�:�h?5�N��a]��t�b�s�'v$] �;e��~�u,]`�V�����hh�B�3��1bqW�eO�v����Q�g�6Fxn��q�l�I4�!o<~�h��* q�f�^�nY�ح�↚�<�o[� ���#]˂t,�o��:m��}�d��ɀ�2�c6���޻
u8�O$��O:�V��CKm��l��WG�Cd�/�u����eH�&�i�bsw�wb���7�f�"}Ō{N��Fv)�}�c�S����n�n�M�L^��>W]�i�"�c�W]� �K���_�?ʶ��y>��#�h��o�n�;�ص�g��C$1+�K+�j�z��q���wc�G>�Wl8v�<��{u�ca֎R҆dm�t�i��K����:R�&lZ�q�:����u�t5���b�}�jK �/���^�񞞿v��m�[ïwެ��/�ѩ��z����h�3����јVF�w�!=hl���I��[��a,�\�R�V�/�@�n��%�HOMc�]�6M��x+�H&�"��+c���}�ӓ״�-���*Xp4�̃�A�C��>����l���h3��AT-/�U䔪S� �\�P&�[�`(\2.޷�ܗ�@x/՝87`��Lz�L��=��z��TR*y�����q ��2i��{�3�ˡ�a_
��x\���Ù�.e<H͆���NGR4�l�#��I���Tj�����9	?�V�DM�ry�+U2��.-�M\=�dT_I�l�m���smLΫ������oH�DuO8Tl�;=�+TU���dD�
�8��83n��k^-��[\ �l0<ˍ�b������kC���O�����K4��d�͒�*rF��y�Fi�`�5׹��p�:���>]w�&�y�Z��j�3$�ݓz0dWڰ��Gy�)�m�z�kIZ�Ca�W�}sƥ�og�]�:x�����L>�jyhSz�.�u���ɱ쫶6W5�\���q�m=��Xi^;��gB��D��Zx?�
�5x��>��η�h��hr�������w�{����}�9�ͻ�n�Q#)Hڤ�=|�S��������H�1��Xy�����^�M�ѻ!�t1��'�$�==!�w-��6����ڧ�<,���������{�,����l3�9��E#v��FOD�x�>H�dcF�l�ꩃY��C0ϴҺ�1n��
!
0
��V"�gn�	\��1#�o-z�gKL�`�g��^=��T���A,��O<Y⢘���ْ��-c�۹���=C�Z�4]� �@�D��,�A]��ʕ�b�W�̝��ݓ�"��{݆�zypM"�I�:��fP�u[��m9*�QcbFIǸc�y�%PL��+P����딕��#^I)�sƫϖ�L���!��T���0����s�������
 �#·�6
7�t�e��c�婲�����6�k�ة�Qߪ�^�_X����x��i��-Ka��Be�K�z��g2��������Z�tM�/%���wL�} ��L\�27�F�"�G%
g�z�����6�#F�)��7�/p:z������s�����f�����8�!m�eB:�5^ť�mZ�9�h3G(f�J���R�*]_�FC���0�v�:�B�2�.�����n����+y�i��cp������q�Ҙq�(����n�ʖwtV��h%�#2��+p�X�c튾��3��I�ރ���8�^��4G�^t�uȮ���w����XvS���7��TІ{���F�j˺fy���&D$���M��:���R���m���b���!��
����^>���`�`�o�׻R�NV���xF�J��= �S�N�c1��=�*j]v���f�e��� %V�u��d��"�WM�Y��_��6����w�g��u&���"b�EZ4�}���K��ݖ��.U7�i�	�V�5N�0�Qǚ
�y~��t@B�x=%[�3nb��
}�[��p�^ܷ�����h!C���^ڟtS��=��!��X�0��0cG㺶��m�R�\C{���M�{��.���:Y����Y�g���� �c���\�]Ѱ�/H�R��T9� ���s/-�j�o�H���ۏ��A�0n�"Q��� q�b�(���sEl{��klA�'/���<Nef��RB��Mצ`�ˮҕ�C�+2�[H��74�DF�5õ4�T�ݰ�FX��`ŉP���B��IZP��ч��V`dj��e�������D�l�nd��"	9bع���d���(�v�0n2���6xPL���S��^�t	���@�2D%��i��i���Lp73ڦ��cj��������:{M:�5���|��I
���-���0g24F��0�^���� �!+��7J���:`���5��U1�B��d��vx �D�^6Si�� i��"O���5��l����ZM�Ψ�f蠝y�c��rqG��n�d�W�����Yywd���i`���Y'N=D�x�cO����H���
���P�K�MD.��&�_���6�]3l���Z�wz��!!�k��ђ7;�W�>�1^x�q5�n��;���}b�C۾��VP��{���I"xǌ�,�f�>�b�uY��
z��?��8]d��3��j\ڹ	gxHrȻWEG���fN�R���0OM4��s&>o(�J�湅�R���ͺ	��wm�v�0ʼq86��R�v�5��'�;��c9�sH!�l�]�������4d]6�1��1���S}�;ͷ#z�����9�;��"a[A��є���jow��2H�Μ�dd]x����z��W�3�w�諷��,5Z����j��\W.Vj1O��ǫ�����	�C��~�M=�^�&��w`���k$�N�(�0ii���=cݹ�!>�C�q�w��LIm��;R�~�b,�]R���b�=aw2���brvG���5]�`�ے�:���ܱF�t�;v��P�w�A�0(G\�_hp�GJ���Szi�鉫�rb�8iѪ��f	�P�lv�u[���Ӛ}��2V7x�9SV�`�y__׃�g�9����s��*O$UP}��S�ݍ���\��`������l���pW?´J���zJec�B�`6�H'�W�«���?T[����{�&R��_��-<�";w@�2Ju�����U*P9l嶵�!익���Ҿ4����eW��s�ne2rS�
�������㸮��}�{�25Z�A<�>mӐ�[�c�q�Cvhj�=����p�2��r!;1X��L����=y�m�?h}���i��1�F����8m��3��\J�R�K#q��X�ڧI��u�2�nq��z�P[Et�-�ޞ�|�z��� �@ӆ��[�{���I,�B��1oB�.��t����;��5��9[p�a�f<��ڪս-Y�$���b
F�7�HA�!�������ʯ[4��5f��r�uf�]�B����7Gy�Ӳ%̤���t��޻�֕@E�׊���.���ݜ_��X45�4�V?�t�yDn5�=�.�ѬY��6A-��v��*�m�}f|_cټMq.Sss6aZ���3N72\=�� �1�:��V�if�嘟oa�
�[n����6A�H��pd�\���.-ԍf�]
�:�QW2:_�M�@�V��kr_o�"'("h$��j$φ=#����A�����_O��������$$��2�O�����d	���0��!$fӎ�DdF#D��!�$�		��!$�HI
 �$ H��B3|&�n�K $ �@ �  �  H  @ �A  @@ d�I� Y$�   `  @  � � �(� @ @ 3	H2  � ��   �0�A� 	# "�0 �A  !@�IPd ��� $a DQ@Q�   �DQ$ ����1 
�� )  �0AH� ����$b$ AD� E��� (�
0�
(�D��AQ��1��E�"���B(�DQ�Q�$��HD!D	$���CQ4������! ,	I �~:����_������|�����#��_��������p��#� L�����w�?� HI:I���������$$����HO����'�g��,?�����P�		'���'���ـ��������2�#�?�L�ퟰ�H�����F0 �@�F E� $�RI �	$�(a	E�	� "� B � � � @@����  �@   " Y ` B �   Ȅ � 	 "H $  � @�  �d �A�H �# �" ������ �H�#$��  a �I#0� A�FH���D��"@� 	2H�$I � �d� �# @@$H�$c 5����?���`��� @�@	 $�B?�zO���,��~�'���?�����		'������fnL���?bۑ8z?'� HI?��?|��?����:��$$�aO�O�C�'�$$���d�d	BI�$�������"Y��|�߰���&�D�!BI�B~��~�?���B��Sa��I����������<����}�D�T�RB����� HI?��=��"��O����F�?�����5�=�3���됄		&�Ȩv00��a>���O�g���B$$��MO�Y��sp�		%�����n��JO����
�2��9��+�������9�>�<�����R(��U*�T�%B�*�$�*�QT�
(��PEQPP�
�R�� DU*�(��%�(UBR��*��T$P%T*��IB�J�I*P���(�RR��(T""��P T�UJ/F��*H$�(�� ��D)PE*D�I!T*�TB)J�UTT�EUUI EQUU!IUE"�DU$R@�I*��DQR��V�R�T��x  +�YZ�5���]�Ѷ���	M��)�-UZ�)�ܪ�U4S0ʣ�[��S�)�wj���k�Z�C\Me�@�Z�n��jUTH�)(��   X�"DK�R�HI*���)%Q"UB�E�����U)�"DIU�:�d$��^��3��A�ۃMl���cv�S�Sk,�7;�v�B��VZ[MuN����H��J�TEET��T*�    ���MW]���c���]��b��Gu-Ӫm��T�[lw0��V�[*�-�R���j�]:49�m�am:��5w��
�`�Q)AQ�U�   ���z�Bꝷf���FPѶj�K'e;�R�VU�����Fp���P��L���]u�\M��gW5]i��܎m�E2v	U ��)@(��"/   ;�7v�n�w�jٛ�wS���qN�S��U:��)̛��V�v���ȣ����-e���֦�����fvΤ�UIJ��U@R��  {ګB��s��]iw���j�'q�j��Wu��]�ݳv�U���U���;�ˮ��R�wf�U�Jn���u�P�*��(��*f���   �S֭V���홭kZ�Ů��kv��uJnܪ�+t�U:d3�:9X�'A�� ���m:�93��0�P�@U@�*�   ��@ j`J�3��� �E��t΅ )�,�] зv�4�(�ep���L � gF��;��JQ%D@��QU*��  =���8��P:�� p�h iX�JҘ�����X ��Ҹ  �i� ���U��P7vd��)J��JJ�I)<  ��� �]ʸ@p� I���um�u0 4`A� �W 4  �܆J:)ۚ�T�Ѽh��@ h �{FRU#@24Ѧ�S�x�CF�  ���R�   O ����4@�J�b���A����F2��b@���������T��V%s"4����Ɍ�饄d(ɍ� x���y���������6���m�6?�0�����6��1�q�m�6={��&~����h�h��h�׍h��ܻ�;4*�0��K�g@ڔ�:u:u��64R{&i[�B�9Q!A0]��]AvP���ҍҙ�6c�Kp'��Lv[�/B�ۙD#���}�W�ud���]K�m���˕�Y���GpS����v�� m�rU��Fҩ��S`]��� �ɴ�wb�=i�tZ�iR;��9ƃw��0���	bR8��IT�CFC�y�4�A����Jt3r*I�qYI�H`���W�/S,,`	^ն���^��##x�P^V|�`��ĭ�1�N�HQ�7�5��3a�6�)��Î��#U���dE�����򵝽;o#��h&D�hzL�m����&0v�F� 5e�6���ǣq�Q���%ə��Vc�eI�GV��&%*�־�/�`%=k(e��`!T�fM�0`��/.%;iB%�s,]���$��M_�,2��J�o4R�yYw��ALX܄�3jD��R���B�E*�WF^����s�vU������,U�r���p��6���/B�kku�0X�J�;�W�{r,�ͬ l�t��t]
�Z&��Sj�-P,1g�17;���Fw��M�V R���+wb��
�h� �eM���Z��b��LE�R�(%2\�e<�Eҕ�U�{�R�T��VњF"i���E8�i�%�ݫ)��]����^�� ���J0Xw``��b%�ڻ2�%�!HY�aT�mb� ���X�NZ��diZj:��ʻhڏ��U�&ź-��V�thk�l���͚�pm�N`�L�`���RVK!Y��#�u�V]hU��
���[X���7&4
�LL3@�7�-�&�(��I�u������b��a�=����r.��լʳ(�U��[I2��]a��Vr�c Z���l
G�[,�eeq�ˍ"vfԍ����Ч�����m"��$�Q淕^̻7��ǚV�h��r�/l�uX��*�E�ϪG��9F�N���FeY��f�A�j�+KA��܇+��ev�w��͐�@�hR��P���dݖ�m[�:���m}f�-b��f6̬���M)i�������[t6
߱��L������F��XIc"?[��������)�cu|n�X�2�l�9n���u�F��1��Rw�A��ۡpɬ;D55̷������n����-�Հ��D@���G�f�7�+�(�/I�J�K��S��$1��nԬm����̤�ж�YV-�jj�eZ;�m�WEݬ��ǡ�p�yJi�N�ۻjի[���t
�A��:.0�ǻ�+k2(	y.�k���#[V�l�qT{7.joѥ�6b,Ф�jKp�L��=�����V"{�(2�q!E; w�u����3#�k(���ʹ������f� ��X�	�#9'b�l=�ѳ�� ޷ j^���eX��Ϧ�ߥВ�A-u��uj�8��e
�d,�С��u���Q\�4�6��7��*�� �n�4n��f��H�Ĩ1�`Ĩ��((	u�VY�4F�� � ��t��3p�C�d:E0�/fb�����*v�*���oan��v����t���W��r�4��c��)��jֻ���ۑ�J��풯N4��KPoY54D,e�n+��=�~��MҚ�Z1��I�XF^&K����PS@�Uz��$�1����F��o�Ц�L�`b�yb�ۖ�B�^P��Q�K�������A���h9��M#tJ�`�1�/u�;ǂ��c�ad[Y��H>;WL�j`SR�l!YRB̽��������#d �ݕdY����Vr�`�yKQ:�M����ϐ�op�2)�-X��Ii���Mnn�f:�`3,̆�/��W�F�[8�/�� ��f]��r��i=#+K���96��-�>ĚX��6AE�ջJŌ�n](���q���i�tE��bW�4m��Y4�ǂ�P9eq 	�]�����D��
��������!�B�)�%b��F��5�v�+��*9�g)�f��fceP1��Ɠ����Z�F��A�n�;/V�k|32Ć���H�S�T�0�#�Ԟ�[�U��񷀓X(U��:�'lٽ��Z���daZ�JKi��R�[uz�t��ę�Mř�k�
`��ݵ���nˠ�U���d���ۭ��B�]��FSpj��T� x�4�[�x�t��rW+.� �Xp���q�eb�V�5{s.��*퇸�.Ԗ'Q�,T�X���03Y����7�6��gf��eqw�-�H�7�>�	���Ǹ�;+%����sU�p�]̸�So
wZ��@���5a�J�u��H��8JFQ�v�*y,�Q��G�I��ͭ36�ԢMMB�k.�n�ƝZ�z��x+U�&���S�?+�cr��q�ɮ�C\���N�[Gkj#���t�m��Ĉ7h���f ���P� �D
�M*WW�i�۽���#�J-�*��-K�� #�lZ��nJx��f˻��w.�J

�EnJ�Ah_+�^UÓj�m@,��i����	#Q����Wbi��U(��wB(��f;��oK�#���A�!B���,r��`�V�nc9w�f�0Bh䭖D�W�r�P���KRIB��-�YN���n�=jT1iw��:��,�2��&��Qҫ�q-��٧�]��xl�P��]��F�+{�D�icz��/�q��V��x4Lj���Z���p��ĝrSL�M]��Zl!��)I��˔>��e"`��>�A'e�f]ը�j�Y�#�[�̺�7[܍ڀۥif�����ɲ��DFB�IG�Z7��E�0M9��i"��k��fT�6�,X"��U��U�@�emm5.��V�c�j�ݐ�^���16�V!2��%�`����]f�6�"vG�)V��̳��+Y��hV�2�*cF[�U&U&.AV��s�
��,ԮS��V�:(ӭ��!;��3af�(�2<�ӪLWR���Ӕ��Jh���L����'O]�[�.��Z.�dhl��ȴ�������,'&M���)hm䨫K*���kV]!v!���xK�� t��0�ym;Eu-UY�m�׵&YC��)=4f�d���Ǘt��X�n����u�KJ��V��m�A��PYr�%[�n�JʍDJ��Soe,KT�b����8(5SU�����X��n�;G9���4i輏Z��r��O��F�ʵ"ߴf���ĩ�Ҩn�$�.G0l����A4D��f*%�vvY��u���fD�5k�;��%��e(�يc/^� sf�4'YCN/�S5�6�jYX-�`�!0@w�i%�*e9� 0�GtغT�ܦ�?W��Q�&L�v��\�G+/réy)+���{up�y��g4�ٰ1��L��i�B�QS0ٰ/[Xv]5�(�LI�-�N�'c�09��m]�-��Y��(*����5Dfi�}�sH˒���ۭK[XڙB��lS��vU��ƛ�o)�Qw�:fQ�t/��j.`G6f��Y��sA�Ō�lu�|f����He���wh*uh`M��N��bGd�����N��@���	�oA�q�&1�%J�eݵ0Z��iXX��Bz.�^�{��Q��ZI���'L`�6�n-�*O.�(��急@�!f<�FJu�r�!��;�os6�ͣ����������`�YǐJ��1h�iU��]���{TdYNڻ��!&�2����ᛏBĖ�Y�S��X��2jm5G/�&�`�����<!�`��VT���[���z���;:��+9S;�&�
V��.70m����lr��҆�t�%4���VqY�8�ݖ�m4sv��q"e$�lҲhݔ4���wR��,�� "+n�,ko\?`�ԝ�7	�tX{fS��2��H�e%VV��l�� n��kiF�ɂ�F�A|m��T6�˦�(�*]�b�Z2�mL����h:B1|a�/I-��	��x�uoV���i[0pQXȳ�:5᪱���ȿ����>:�B�4蛸�ɨ�
;[��D굵yŁJ�Vp�n냾^�ȱ��i_\8�mZ��m����dZ��%Zc�^�G1�dScۚUX�!��|h�$��NK�@4���qJYhC���$��ž�5�k85٬Z�c&l2�l��24$��	d��1�X����v�<G����#M��E�^	IZ�d��@��f8u���ɲ���S�VZn��&^�E��1�B�è6�����n�l, SںA桇@ w�% �E��j��kV���s͹�|����e��G"ͽ�P`�d�lb��A���hhOl��OV6�/��X�#(^��iۅ�a�D�Z��V����a�쭌f�n���7�Q���k�ʷ�|��u�V�	$Q�b�U��RBr��X+F����җ��yG#k�w���l޽rD���k�Z��{W0��\��si��"�7fա76��aT��2GF[�h͊Ōin<M�ܶ��f�QT<YA�2CZtL*z q���� 9����n�;X�XkJ�;Z���I�SFD��e����;��˿��d�B*�ݪV�dV��2�1ކc�o��2!PI��o��+2��l�e^��K�'qlhDR[+0��gfBmAK�5��iF�j�e���yV^ʰ7%�(RB������VB�Y*VJd��˪�VU�yR��
�n��:��OiPթSk�i�)-ּT��[��\�YS/j��+0���T����dqAwl�1$�n:Yn�\�L�˫���;.�H�[�V��F�C2�����¨�ۡe
���)��a��u*����b���W��w@���Z/Cs#v�V!�(����{�Ol�
)PjȤv�J�V�t�ۗ-b�e�٭�u/vnK��%8֓�j+ ���O-�	t�8�5���c:4�t(��v�e7O�U�e�6�8!ɛD�j��Nʊ�ݵYWR�L`l�������ҷ@n�6ݸ�+���`�0eI����v�ɵ���`�F6P�A�voi��6\1�4e;s*^*X��n��	0!V�szW���GS��T
V�
b�5ѵ��3bncy�j9���)LH��F�\(���
n��[-l�p�{sFf�t��;R��-
M<���W1�i��nE[xTWY�i`E�7te�F���
o�;����V�E��}h�i��gRY�Kq�w;��W�Cq&��^�J݋�F<����U軅%㧴�S0I,��fM�%V���JU�;әz�Ye���҄ҫP�Hn\�Z3u���p��lۉ��V0��
ʂ�p��ZT]FV-Ī�f�
O�%�K��)<a[#kmSU����K5��̸C)�pc	�4��ƙ#n�Fr`��@fJ���Q���YD4Y�U���-����Ǖ���Ц�2ˡ���i�6�xUѼ4!���A&�ʽ�2"B�^�q����n͔T��U��O����џbE��РVV��D�׌ұ��w���plC���3�����ȢF�� =����'fLK$"+ņ�Pl%�YaC�q�P�n1��B�B]T'M4��Cs661S�vJ�+M96�PS2�=t/M�{2���jZ�zB���(�u.'��V��T��/fVj�lJ�H�b:s&�F�!�q�wt�i�HkE��U�� d	��*@�Pϖ;��GXn����7��7.���r�n|Ƌ�wZ���z��tw��\�Z-��no>��)lV�U��ohi� �!��3��j+ 3hbτ(E�m7�a�&��i�pޘ�BK�u��.����
�ޤ.�5��1
�a�An��a�<O&j�r�lX�Uc1(Vi[B�[����a�U�7�#aT���g#�$r��P6%�M��AI� ��GE���*�&9z�	���5t3�n�U�ܥ��[-��L�䲦L��,�\�A�#]�7��(�D�YNd�u%��֪I����]�ܶ3hl4�ڕ`Pǚ-�6@��n%��;{;Lf>�V
�1���`�i�nU�!Ƙ�kvü�Q�l]��P-��-�c�wa`2A�K>Rj�S�9dV�r3A�4����X7L�����n�����̖���97�"I9ua�����^n!3q������em�nRq�(ݱ���!iE���C-"+["Ȍ�-`��Bf�
܆!�Gx�G�e���ڼ�O���[�"�U�x]���ĥ\%��1�������2�J��z*(��Qů,��`S�-�5�X �Qf��ʏ Ֆ[]
��5L��$����<��s�ҷ�[u �X�&�:����5��0|�+y��D	M�{*^&9(�ʺ��@DܧvZ� �����!A�5r�PQ��3`d+��Zj��֋�d��I��'��4U��C)�ѩB,Ėj�sF��nK��)�S��$��ծZiK��r�%�����|�H��)-�;*�V�!geU�X7d$Q�<H���U�`f� 4ǩ�ߒ���0eN�9���Q��-m=�Db"8�3w(7V������"DfV
)^ 흺���2��a�e5�h8D����L�ݚ�ĤjՔiV�ϕYFSm�u�v)�2C�Q?=����dmfck������դ���#�(���)[�����C�b��"8tSܭ�-٣�(emj��#ZR��r�Ai����_��S⭁ .�
Y�����2�۹�n�7u��87._P=��:p!�sNnq*up9�I��dml�G��٤&p���!��;;c����s;�I6�>sZ8pm��2��]�� �8�.������K�c��Cxx���J����z��Clw\�%���C���h_�r��u��K��!U�3)_dU���b�;��[.�.k��n
�/�9��	\�r):�\��p��})�7w/�AƵb�+i��.�ᥧ&�N���dJ�V�]v+'@8jT	��ea�q�O�����	��1��V�����Me���J�Ku��f����Ď]���+{(�p�2�s������+b��>G<���:WX;q��ǹ��q
���d�z�:7�El�`���9H���ښGN��6���u���DI����dh�3D���z�D���$�n��B�Mfx-(�i���Ĥiaε�8�FݥP�]
'������Mx{-���V��1�v:��<y�,N5�$�.Y��«�xbV�����Cn�ơ�!�i9ɮI�<�R�)�k���-ÄuŌ�x��Es"��n��:�p����K��!�O(�������7j�/M݄��ވ<;8�'��l#��K��ҵa�2O��ʽ&�F�=�+�EE�ƶ69fW%�V����sF`%`��#��^�[�h�AjU��f�r݉�0q$�tNe�L�P���yRkS��<�zb�IS<krw��9��q<���b���Ӓ[�n.���:�!��[��Z=6E�l�PuZ�np'k/FΧ&X�\��)���Ǻ�kw��h�r�J��}mN��Cs��ʙ��m����nҼ̯[v���l�c'[��i�d��-��v��:�8#t��yݤal���*4u�`U�˅n퓮whл�:YKE�c�������6zN���Ď�K��GI�;��U�d��jU�.�]�u^�NpK����Le/��e��ٶo)7s�h-g7�|6s����Zy�#�ujy�C2P�ۦu��3�f�3��p��s��Ö��д�,]V YG�z���H^Ǖku��WP�h�s;�'���3*!W¶^�*9��o�U%R*%�t����rA�N�*<�_A��z�/�Q�/�,D
�O˺�#{2�F���׳���*p�o���n�㔇ti�T���Ws�͠��)n�J��wx'��ޤ����n�#w�ۯ͇ ؞�-�&ћ�hL�{�Z�pu�V���21Y���]6�š�%ȳzPnM˗�ʤ�M`��۹�oq�W@I'c�D�k�[��*��w���b9[��ؐ��U��9Y�t��B�@5�M�Fp[�WM��av�lp�����U�k'�F��*Έ
� ��� �S� q�'�a{:�"��ګ�s>���N�'��]�rJY�l֙���Q�.�G(�Uj���j`�'-J�v�����If9�C��^�j��7��u��X��X��̓��k�����b�5��q[�����i��+��"H�@�؞.� ��R�o/������zQ<��%Z�z&�Kp�X��&�y"m��|]3�Q���_q�ͤ�)[��Yem�kAy�#���.�9���Kv�B�T����ʳFV]nӍ>�o�������G*�Un�t�l\�dܳP��_	x��ŕ;�+#�v�>��a�(�����9�=^��ӵq:�+ ����+�L�X5RI�Ώ{�����zk��YGb���۝!+GN�^u,ň^\4)�C;�z�tK4VNfTY�ϗ����aֽ���v>��i[��_Cr�l�%k6�cU��E����X���ov�.�D���_M�w�=F�{�0qOC���g)�[m���r�T]ˁbh�ޗuI*��Z������1>;��\��]����9[z�0k^�!��	]E,�B�vf�p��E�VWU�ϡ�O)#+Gu>-E���&�5f���%)ׯ��W��w=ز��ANe@�W]nX�O���f�:Z���{q�@�ӫo�t3L)n٧��l,,T0�"�َ�npu����#H����!u�:�C6�vɽ�л{����)�h��ήǉ(���qLإ����g>s�ս�Sop�i%W]�닥�J8#W��7E����B��qӕ�S�[���;���|��sq��ܫ�$�"�b��:N��L+\,f��Bg��j�z:a���v�P��������65S��`voZ��,�����ZoS99:�ҷ@-j�Z���*�]jh�w/�����_k�cb�i�/��'	�r���D0��|����/�v6�V����Bgpc���!B��0�67��D�y���D���5aյ.�o^���f���
��ź�Q(Q�&C�v���(�v̶I�� t��76oT�ig1�=M�,�����o8?�ݞA~^C��^�U��;�_�\��J"V�_[�ܶ���=O��M���@� ��6���<�mB4��q.�k���`oP��E�낞����w$���f)����Xo�y�]]�>�(�]XX�Gu�qo9���1o0�	;�Ch'-^�t��o����������7R�#�c���x_Y�3I� [۔�z���+����e ���	Z&���fv+T��5*�X,�У°k&P�r�x�� �{��p�Is��:V��n��R�K�n�1h�jmH�[8�s��%F�c�V��C9]���>�u�b̧ї:u�+�͙yW����h���i53\&�	ͼ����Ŧ�Uה��X^�։���bu�y�Y�����es������c��]_gQ{��R��5p�5�*y��E�������c��ƝsV��%���+�Eٻ��;U���엍����t����t��7�hefDsl�A�ڕ�
]�-���Y��z�n�83êV�a<�N9L*+�qs��P����5��*�Xr>�[��*vr'u�Ѿ5E�ƠeE(�W�;۹��^攠yJ(v�|hRH[O{;�^m����\HA�4n���2���Dv�>�Z7��+��ﳆ�����؛�������|Ы�_ǂ�w�b;J^G;��5h�S.}4v�6��pK+�`㸈��m����g��F ���8w3�8�$G
�)��n�����l�qR;>[�p-����]�CzdnJ�����aj�]�9�Ҝ`�WV:e��T8v�i���ʠڵ�);���<�[�ޭs�>hԹx`}��n�cOX�p�-�ӡ�3���EL�o8'G�J�(�I/�i"�X�*ϐ�d#��1}.�A[�p�SGv����[�����9L躕�Y���1�S/ὂS/�IOj�j�ɻ�}�]>j���k&�t���MV3s�fہ��rq�?Hj�$D�Zp�^1���uP�,�u`�� ������!�ۋ,<3�=�r�f���Ү�S��6V��$��}G�mu�D�ŝ�1V�@�ɹܮM��Ż���x�#ε�������U8 �6ΖI�.��V��]3����� ũj���;x�)pýo��vG�,U�ZvNƳ\�䫲�8�f.ʾJ��XR��k�]���/�"ڝFo,m�\����唖��<�i�'���ڱg2e�)�,�^���wZY�`n#�]�;�)���A�m�����wpN�k���.�6.ޤ���m��_VJH�^� ��5�GF)��̃��B�Q�>ab/o:��PmY�׶`���V�}j��חѐMN٧��(2����G�+�0N�2�,�/�����Y>�����kG*�̘�[���0n��U}���ya(�W5wrW��U�u1`f��i���A�A��_Fd���Q�|p�ߑ�2�T��,�O��Kĕ�u�c	�^r��a����^�j��yj�&@��}$�8Z�%
�.����#i�e��;Bǉu����U�A���s��S�3^Rh&�>/��j�n������m�;.�[�\l��-�
_X��ԏ���I�I�$!�z⎉2^vP�8ek��2:�j�_Vm,vr޼�d#��(��l�-kQTE��SӺ
�+%v�I�}��fg�(u<�/T�k�j���5}/&��pSb���s�('������T���ܛ�z�%	��cs����D���F_���c�_n�9�V��J�+����MN7I4������6����^xī��" Va�paBŤ�=�x#�5RY�~��p2�;���K�c���(T8V�*����mq�z����fG:�d���#�{
�F��#\��7�a���p���s����z���[��i�r�&��V^�D��uύ
RX0fѣ��+!m�H�D���c��ݰ����!X��~�0�r�N��W$"U0�>�Ÿ(d�׎��g�Z������鶹^ �n�q�U��}�4C����˅DާؒF#>,�������^�ŧ���;�NN�뛨�hs\�t�tĶ0�{g�U���/�1�mƾξV��V-��=�f�뻹:�ŬL�a���K9n�:`��ք/u�.����c&�dy6��h�(��A�P8h�E����CHr(l7y��ΡqI�*s���Ļ��N�.(P�*]��i>�dd���ff<��>Y�+"�Mm���p��T�7��ʓ �}R�ھ�o4Tw��H^s����A�
2��v7�t`^iR��Uh�.�2��v���yЋ9WN��za��;�B��T����f-�r� �2����7�I���d��w0_P�E��c�=��U��`�\���F���	Z�mgu���;���/������}٨[ī��Xl�¾�A�r�	�ݤ��+��33��6�K��]r:�|o�ݎ�X>�P�^���|iwac���@�L�T�d�Ŗ�+r�&��S��W%z��|��9˷������ M^#��;\4=5�
Zi�|�C���k[=�fN����rfV��eU�*��Pȫ
L6��Z#<�I4��j�����j�@V���lH	݄���z;`���Z�X9e
V������2��_:7ً�`�!��XU��0@�t
"�G�wvEݜa�x�m��g)>9��j�.�
�ӵ�-��L���O�f
*�{��j�����h�ɗ��GF��'��uec���O�J�[=Y��+7��T͔�� ��ʍ){rq<�Y���{�+� 0}{ԭ�!�:vl��MD/�[[nPV���/g7ёHnrф�:<�;��f���3��|���.n�K�}]���lIa�篥N��}��}�]��{w;��Sz��;���0��P������µ0@��`��+��i����:��z����˜��r�+�+RՌ�8�E���+��z�IK�/���R�GV�:�ŝ�Qc/kP-c����6�6�8{�g7O���	�^�*�J�����I�AZ.�K�����k`���:]��FoCtRZ���DI��&�T��^h�឴O�j������\�^�A
�J��DJv:u|Mb����m\�e4����H����w����,�y�X�z0���O�əCM^��c����^��|9��L�'<2������R���oR�"�D���7c-Z�Տm&C|�<e��;��$WF"�����o"��;�8cZ��i���Yܶ�yep��7��]��HNf������X[.���%Z��h9����l`a�"t!�ښ��Va�]�4���D���5��dʅp�Y��]Z�rsS�KxP2%dӽ���uù���eJ}Na�m\�Oݐp��.�&��ɖ/n��+D���At�ywNRͧ�������u�T��|�];g�-B��)1��d���cz����g�Q��^u����>��먮L�k���,�ǶƱ�C���We"����rFX�@�� �����M�`��5+n>bN�z(D�ł[t�7��ۋ��
@o"�����ww����H+a7���6�_�}Ln����b�P�]TiDF]J-Wa�[�-�]�r����Nv�>��b� [�O�е�k5���Rb�-�{���!����{I����e�^mg}h�~�\�7��Q4��v��0R�(�r�B�ۖ���u�۾Q�J��i�p�����m�D�js���65�r�3c+��3Yhg��N�i�q6�����ɋ4ۨ���x�ұ��� v��:~�t�U�!�K�o�Z��S�қ���Ża�]9��ۮ���e�7�!�
IT{��,�=z�{@<O�V�MV�U>-�f�E�f�5Ra�E�jkN�
x�'[��������Y�6{9��*e�J���s�p�,<�2��̟K{4[X�Z�E�i�M�b�B�C��x>R��P��w��7n�i��;7���cbC�kvB�x�A�{�l.�Үqw���}��n���o{��Y�i�LrKU=���۽��P��N� �[դ�V��:��83��T�+0���2�\�Nۡ!��R�J��n
QUpǅ&/�]N%'
��k3��X�o��%�p��;F�Z�ָ4 b����B?�t�C����찹�n�cٲ�6�m\�KI���#1��
S��t��֜G6�4=+g�hWc����Q�Qe0e^��L�9`В�[q�ݽ@ev���ur�O3�o-�v��R��dnm m����͌Э�uFW^g9��OU�8�������˶n�o؝ʏw8�Ŭ��ˮ��q�;(>Ő��X�����o��S���:=i��O7ZI���y�#h�ѷ��Yw�E,ܸN	ls�a��Z�˺�Q� �j�o~�'T�8̴�P�ۃ��%�M��[�go+v����>�g0�k7�h�.n���d0�mh�ö�o�%񤲣��f?��Z�*�����XӼ�����تZ�.�@WN��z�Z�v��L�/�$�i�}4U�>.ۅ3:�=�;�.��M���NoIx�RWK���j��Q.kYݷ�}�w�z�uvw������x xx{޻��5@�n�����µ �_�zڍ�.�@P�*}w�8A�b͠±I|�/�:Ť�Y�S��ۘ���m��b��t�^'t�[8;�G ��r2�J����ӧf�oU����hYJ"��6�˥IG�g�H��U���/tC������nv���n�l%4u���p���;�=J��
����u�A�wm`ô�Q��)�Μw���7�X��a�z{L��V(��Г2RF��f�:�n5i�NZ�1�E�����K'JM�5{ݮ�Ǣ]đ�n(��S���>ڲ�;�|��B��)��[��)Y��n�,ї�Z�2�g�2XqR�)���w+{H��YW�f�$� XS@�y,F=�cw[�L��8S�	�n/�6�J�28g׃�^���%�Ǽ/����s�t/jgD�b'+��.�p=bQ�\ }�_T����%�3)E̜�DI�m\�P���#���5f�Þ�{�T�G���������X��wv�Z��m��<����\�����㵊���Jm��@��s���j�C����) V�[�-�n�Z�^p��C����:��nn=d�\���feo*�5���vp3I�ŕ��ً{���N�RxH����i�ALE �Z�ܹ����1m����#Z���EP��6	Ӎt�6��	֊c�[��_u�u�jh���:v �սZY{7qh��9(TU�}�9ػ��iu�_ms�e�Es�����g��|Z�뿄+�ظ�7f]k�P��{�V��Dz��H����\�ƙTM�����ݎ��m��*��Z�@wW7oW��w7s��P���j�Je)m���g&��fcuLu�']��u������ރ���fP/����5�|�b�ܫ�/e,H�=:є���t�	�s��q�ql'i����;���[v��G���S�X'��i_�nj���k�#��'fkY���^�Ƈmp�UuvÙ��{(�W���z�X�kDmo:h�^[�K.5Z����41�J��xw#�Z�{�,�U	 K�i7�m�[�wK��F��2�Kv2a��&u�Xu��U��U;un�fU�1�ͦ.��n)�;�*өCE�9r��n����VԾ�,ѵ��qhn�]e�,�:�$�ڨ2��C�5;
���`K6՘��[�����-cC[.P��r�]�}9��O���S�fL�E�o]lި��Ƹ�D�6��ۈ���6hb,�ōGs+m,�+/wQ�s{�r����Q�)ci�����(a��f��@ޗ���K.�L��&5fh\.�7��u�H��Z�[��}��4i��NY���rPq=B���)T:�E#�[]͊��p�7�e�u�����U,J��@���W��=��Jh9�v\�ϴ+w���,P�� �Fʧ}y�����b�ٜ;��$��k�(P辺b�r��B�r�]�ǅpݤ`�XZ�]]���0�!GPpjÁoh��49��͊r�B���f��K�y��� ����2��@������y��[��k��!�&�O��.�4r|�XN+4�+?mж	�w�_�lG�U���܌
�,[N�OhE�E��G_C��c���[��ZF���/P�%��[Z��Q�<$��e�b�2����;2Ƹ�a�f�o�zW&���2����P#9�ث@�"��z�wIP*�1�*�.�@k��;q�{� :;�At���&fK��r͗�Q�����Հha��0��R�⻸>�q�,�]�tsMwpf2Tl��/g>i�,V!�G ���XR|#��!na��� ����nu�}��c=F���Z��R��(C�;�/:�F��$	ʝKt�Ӕ5����3���Y5u�k�(���5�L5è��m�f��=}l7���A�ܢ)!1�¶�"��y���w��"����j�r�κ>\bHWk�V�],������ߧ-(����˰]lG(�_gtV����=�R�,eW_��)�s��i,����2�4��rU��c�0,����yD�v��Z <�doo^#�U�b��v*N�9`۰�č\��/`J��	Ӿ����+*^��;7z�����-�p�۶`x���N��F��&H�s�)�� UƝ<g�v��Z�����i[�˳0����_�:L��ꙶi%��uv��Y���ؘx
��8f�N}>�珗+չ	��P�M�)J�In5�m��v��4�.v~&�x���'TɄ�'���ƻ�f�5�/Z	J� :�\\F��Lh����6t��IK[>w۠�:�x_N�T����71��i]p�1Ы��ϤyX2M���`���o\ۈHKRj{�T�d�\����t=�:�;ǁ�Q�,�Y�q<E^�r�g�tg�X56�f�f����jp���I�-�0�Չ���N�=��s;���)�C��Jɫ�	�WY��9v�|b׈Gw�{�N����(+�y]��gh�a��!u(�A�爜Gn��J�0�)��Y���u7I3���SnE���3�������#���30J��_�fQ���T�������������}��mm,9&�eR`�B sR8����t9\�����s�b�{��|��r;rL:OuwK»-9��N�<x���D�}]�փ��s�h��2��V���J�A`TŊ��\�y�=}���j�^5��ëe8�/
f>np;sX���=X���kWl�/k,�l#�˩�^��v
�vh�>���E�)��\9CQ��݃� ���q�B.�l����w���e��^7�Ev9*��	���6�;�[X�&
0PT���a7J�
��&����5�T����,���q��s\aL�����h�Y�4�z9��|Ax;;�<��ml������>��Zɀؽ��ۮ��;����f�VL�t���3,t����'p&��Tj4Î>[{Ko9�[���4�Ũ���Cq�"�{�խ�Q����b�ig^��y$����\�#q�X��r��m��`ڎXl���f��M˦�nݎ���{l�P:ξ��t��{�_el���;���źh��,e�j��b�)�Z�-�-�փN���F�ve��T�Pb�ݗȍ��?��T�9���*;/K�m5ը��+EѳAh���������� ��f>F�r��6��>��q��lP��2�C�au<�̭��l;\۷B��V���{�]�6�����'����&|/&�6�^�M5k���D�P��W�P�`ϓ�ݺ���<w����;���םv+jW%����ۡ�(W�j�8{.�x�n�>鐣��U�|�����s{G�%� L�0]�}s��[�6��&�-�2��*���+�A�\����H��v^i���T��S��y��T7sN��N,�2�V�����N#��f̻���'*��C��86,5�V>���ƭ"�l���+�D�ߏ(X1��7�^�p���ޮ�u�T邍.�7��[���=-��;��uaM&�X����A�Z٨�U����k������.���%B�h�Av��5��X��|o����Z��W�*rW[�⻞�x�4_)�;e��aL]�e�y�qm��!�u��@���J�����1۴��w�6�-ڕڑ��8'x�9�YSz���S�*}0��U۾��3t���"ۺ$ ����w�f�Tҭy������8P
w}]�Ρt��y�8�I) ��dX(Xۋ7DHh4�9�3w�Ճ��]ضo��3��k�4�U΂�: ��B�p�����Vr�X��8�7[���v3n�]�Z��Sx�oa�����ŵ�=^M�j��rMk��m�AB:��vl�7p��.��h؃i�ƙz霩�rƫL&��I�'Z,��o�)-�ġ�tO���+�XÍ�Y|�����i̡�:��e������A���ʹ(��ס��
���\{o۝��
�_%(�Q�
�R��.�
Ӝ��)��ro!�»��]��$�sv�:��J�u%O\Mf�$,�S�������6{y]fq���v��D��F�L��Ӷ��Q,�$����.�n���\�]���,�]�HCU�`6���+�A�Ra��B���=l����3�uXd��po=��E˶�x�o����փ�Xs�q��p!��]"5n��=�:/7]aZ�P��73���c�0�}��T7�X^Q�34*�V����i_G,��P�x�]��T��t4/�s[�����Y�K9�*o*�Ƅ��^��0,;�<CP�)�;��4���(@W���uֹЙ��R�KB����1n�v��뺔R��6)F�w����ͥ�7V�B)S\�<���ތ"gJʜk3�[X�YVb�h�$c�pX�X*�!KR�*h�"���P�(XR���5c���X6+�ܾS&RT�x���z�n�h:���]�O^*s���NAM�ڴU1�Vs���XW8n���[��8��V�V{U7m��}}��C.mڴ�QC8
]���iPB���eGmf]m���p���v���S:9����f�z��)SEoU���r5�5�m|;\��u170�`o)E�v�G�jݗ�@r��8;r�oF��e�Gn��3�}A�V[�Va���#�
�\[6w���\�i�W3�j�"d�x�>A�:�1�J�w�j�u�ha��%I!9�Gn�*����t�o^������g��N�����U��X�Gx�����:7o���m��m�eM��b�I�ئ5����`�����ek��M1����y2�J�0�T�h_n���'�,�[j5��5	R�'+�:V6�b�v���v!N�6�s��n�u��v
���녑j	2>+�N�3��S;VE3ī䷀��#�GM2Bw|b�Ԓ�x&d�':�]�CS�s���)N6���=�&�����C��'{�����qi6� #�pt�o��&Q\�P�7��pqɭ�u2]X���ŵ��K��ԥ%6@���6HH�*�(�$)YtDK-�m'AZ[q�ҙ&�0醧L�ĩ哉.�)�u,wes� (����BV���S�B!�Q8�nQ����c=+
�J_��{6Xײ֊W�Pc'i�zP՝�s�*�V5�򋩜ڮ�+����C�ښ��auctk��6�z���:ܣZ�A�Ӊʻ���ԫ�;)���P�7 ��N��0�Kw�+~\�A������[�ҝ[��°\*�"&�W9�[�l8z�ӎ�v�w`D��n4��O�^%o��R���˛{���.r9bB�]��{P�COv�%ȕ�U�$��}�F�a�/�pM�h�Ͳr��A5�P�d9�k}�sFo*/��-���F�7`�2�nTt>�:9���i�A�t���'��ӓ��WF�Y�PU�4f���_��L-�����m �^69��V��]
|&i��ֱGtxz�p��{�:2nQ�ǞC�rj�	i��[-[�V	>����y��mx����9w��9��oEvJg���%����7ڟK�Վ��yD#���_Ơ�OG!w/J���TM���s��wI꾥9Q:�jS��Y�z&e6V��r�G/�5mqS�V�%
eeޭ�X�0a�;1�7-+�Z6�˹��ޠp���	d�x�CMjn�����*�8��w��O*Z2ݱ��vIb�Y�]�^!^um��|(�i��̙�76�_+j>#�&��f
�&�b�\��;s���ϕ��h]�@�YUd�I�Ò��ɫ�6�Ó�V���j��J��n�Ή�Nq����n�7q�<\|^��m�%m+��U%"4��Y��tݸ wVweѣ�Ñj��y��=Y0gZp5��t��|��r�����\ܖ��1rJ˾�Y����b����	��f ��R"�!=wE�1�_A��Z�>H��^���"â��U�L����V��q
JLh,�J�~ç��:vm����j���U�7�娬
�DS�p�j�c��4Q� י�w�oe�M w^�1�O��R$�N�i�2�\;�7�����ǥ퐯�����/[����S�� `MWb����J�ޝ��Mr��G�Y!�{��As���6�WNx>�ki�!}���YՉ_TGM�*՜{��9e���ч.� ��֙��=Vô��Z{���VrcP6��;X���
/�]e�\���R�4�E`�Ź�x�SC=ٹ:5�B"�W4���N�X��G�ybl��8LQ���Q��q[W�ҋ����V-v��sU���X/.K��V�$ʺk&���D�"Lͻr�<���	����Ĵ�cq�\(�����ܔ��CA"��ڢ4
��^��ѻ[:����i6���,}X�M��E�.���ؽ?CX��ݾ΂Y�o�؍�G�n����Z�$���"b�:ô8w-�ʛ0��u
�M�+IWWM��v�]�]*���!���·\�S"6_bt�(w�=uu�i�G��p8s��z;j�(��������x�a��,�S6��ڔƓ]�v6�u�+�����# 9H+��L���[�Ôz+Rd�sb.�Vuf��k{���v��z:������X�p�ǉԎv�
��n�n�h�F-R����1Wl4���H��O����s᫹�(�n�,�6B�|v;��[��-��?r鮖��$LG$r��nrW�t�Y��1	CxR�b�Ղ�^8�6�t�v]�L��f-bP�u��h�	9;�/��P�����I�0����O���\�k ��&g4�:L���f,�@���Y���7i��.8�.�#+G�
�_:�3�)�:U�E�0�YR���:̧P�8�z��&Z���mQ�N�^Eq��'�4WM��I&��J����y�s,��9��_SJ�4���Mb�� �PEQ�]�d����c�"�TL��< ����#�ι�+��j�\��V�
��v	�RXʇ���K7�;Oa��a���ӷ���%�*�S�Ә\�G�C���t0l���:%��ٚ�4��ў�/����]0V"o�7b��
}|�3��s4s���;���R�}�����9a�<�iĝ�S"�t��Q�˔$��6�u/`�[��\��xԖe��XfvaGq��Q.�p�u�>xt)�yk���x����I[{��y��)I�X$�[�a*�'i��ssj�6Z?�O��X#o]+;A�Ә�Q��U��`4��)�P���;օ.ә|,�W��5ܡ�u��m�WفR�K&�v�S�XΠ�����N�gd�F��eG��]f�0`�����z3�w�V<Ӻ�A֔�Wm4�3�I��o$��C;�7�9�o��z�gU���W����6���O\�ل��nަy�)���n��T���0Е�����mm`)�]D_-��Ί�E�5_w_wQ� X�����y랴��׆�`�k�*��ށ��W��/z�x�Z���ә�	��m�ܙz"��eoGݒ�7oI���Ls>*��ܙ�l,�r���&	ى�Uz��y�����]�9%s�9�W�����\�ԍ��jݹG3.6�J���m ߗ�%t������aj��ٔ�/�c�@�I�@3��+f��4Us�����\=�%4p���uw\*V���"���z���^�
��]��Ji�H�R��R��]��6�U#���\!��tˑ�R���^,�s��'V�������0<�]�R+��x�z��C�'/P��1=���RH�p�=��ܜ�:gO$�w0�wws	w<�<Ξy�u�$�n��7\H�I�+�8Q��N��x��E�t*w'3w�' �d��\�sq��<�n�����9�����;�z9��y���!1\��wRr��-�Bw\�7+%�["�nV����ss-T���뇁���K���<���g�]�d�+���RW�*����蜝GP]ܽ�$�s�\�\��d�{����v�[��5�=n���Ea�,U��ܗ1R�\"�b�Kqu-�j^�����wH���yYE&�T�2�LP���B�(���]v� �Ts!3���V�����׶;	(EdNy��c;��7�N�I��Yw>.�kf�W��@��t�||��pU�]U�p����Q�we
�K���Vo\�ݭ'4DU�N��d��-��'z2�Bx���j�u�?vF�)���E�=���R8n�=.R�Q]�j��W�\f�}������Y>�d�}�֕�!��C:-{�*Y�Sږ����UFA���M���ش��:�H;C[�79��}K�|j��ճ\<�������m	l�|ſ0��>�^0�F��]�]ʽk���Q��S�܊���S.����k��:ǁ������D�F���թrN����J5��ߍ���ߝO�7s��<*ei��|�9���+>�p�t�+�8+����v��Ȣ�E����p;�FÑ׷�$WD���[�ԗ��6����[����"�!GO�BT�C�Fn��N[G�qa��Z��L���ڐW-\/�u��i}�'\�])���-]v w\�nS4��Q8�{���q�+r�U���x��'��������p���	q#V���EM<��S��l,�u�p�]��vV��S��sP`X ��Z�xM��բ�[ql,����j�m��wc4	��=�s7�]�3/G3���T���Wn㫈j��F3f��q��K�}Z�M��!Ո]�9��k;��גּ�.W[Fwp'm���Eǝ������[Zh緱�r�pqmzׇ�|��u"x��4☷#����h]��$�t�ZY�/Jdh�s�Jo��]d3�9��T�Ab�*Z�\OI�Z޷�<��|7zcԨi�(>�d��XӔ0��5H����}<x��B�f���6��m�	���~Q5Ŭ]���v"�	������EvC�r�VM{v��_p�}�^�[u������SßO�������������|������aƻ��[��݁`3^�.E�&y�{8S���?_l�.ִ�o7$�2oP�����bB��$h�k�5��7������o�Ou�X����+2�@x�ut���r��
|��nV{S��j�x��2�>��Lu���к�_F�j����$(fC.bbǄ�������q��_�p1�%�}�Gv>s�=e7ľz z�gޫV�\�x�&l���$�[��P�C\�{){�n@�CrKC/�"�-r}�l�����}�I̅V������)w���b�����!����I�QaBx-�O�T������W�k�y���h��4M0�m�z�olJɻ�Yb��67���~�2Ujnk�^䬭[f�!b&�ȊB��	Xx���wuvW��!8���:�k�gZ�w�@���6Iw��Zk3_R����FӒlq_݇Tع���>�9᲻\���7b�]�`�^�F�>'E�K��+l��<�j |�"=�m8dA��9��ȷ�Ru�ܻq�y���H̠���������I	ir��Г���ݙ�*�K�}Y�a/c�"Ӟ(�<��������J��M/��<[�A�xCW���ݡ����`���"�z�ׂt�_��u����L���<n�d������k����G�Ӥ	��t�;x�o�ng����Q�^�*�GK��^�'˗��S�}�Z���CC��?bm�;��g�P��3����]Ӊ�uq�a��"���i��/Vr����\�:��W�Y�s��f�{ɏ��'��z�*��N��o�O�Ȱ�o�d��rGx�k�$z��u<��U����%W����H���ڡ4w���#ج�n�U�lT�q$��*x7M��sw��,Hd���+�C<�SI�=6L�O"EG&����c�)sn�l��qn^Q��'�s#��$[��C7���L���)T���H�#!ڄ��Z^�X�O>�z+9u~Y�'B�{����|D�ł��<���b�k�j�be��4��p�����L���u��(�`�:%�2�J&���\����Y�Z2�ԗz�Q<�\�hu?���Z��Ur$��={��f����WH���O e�p^�1��T�j��a����W4W�=�f�g��T��p���w:�<Y=���R5��اՍ��^���Aee�	굕%����$�mG��7i�4��gz!���򘬦�\�=�E?/t���^�F�(V\و!�k��*�5^Y�:�ܾT��,�)��~l�돫��'��Vmzw�.��J�*u'���;���H����^��#S��4ꇡ���m�Z���{g�x�fs8gd��.�F�(�\�Nr��l�;��f�^�7�n�_jm�댅�r>��a<px�c5]b^����K\w�EC`��Wx�~aZ�>!��d��u:���*%�mޙj�	aV��$���׉�|��ے���Q��1�|?tK%d�C� H����,И��"#�������61��zܓد#j�#���]������M���r��h ϘG�:��D��[`���b�i�Q/\졹��{��P�t�ح�#|�}̪K�tsb@�ĎC۫-Ğŀ@�"��*��⥙�[��F_r�콰���<Q㵒��Z��.�ݹ@�{C���ηw���>'�kh���S@U$������c��X�����8\��-4Tޡ��㓉�گs��c����6�����T�B	pS�ꉥ�L��9V+�	��`S�]%�Q�f�T|�X�<",�E����s�FSr�c��S@tAF��÷I�C��;��ׂM���1����)!�P�V�4��M�L��]��Y��WB]SPy%�L"6"}��5Gw��^Oٽ�QFu�#�^4�>=�ٽ���era!\�W��n]��L��:3ת�s���/R���%W��[hL,.�]�D��Y�PYb=��ZN�p����_u�n��5ts��u�Q/�Rb�vէr&;g1\������'5�3m�Ԧ����ܗۖi��Y6��n���x��il����ڃ��Yϲ.��9]ʰ+J���9L�ȝ*!H���S��#X�ڭO\�3r���yTkS���M&tR�dT�}2�Qc��q�� �>�x����lN����B6���$�U�\���_WVD�a��W˲�e��q�2�Õ�Ԯ�g��e��͇2�J�^�7"���Q������][��N���FO�_o_�0E�f}5j���͑���ZQ����o�̶��O�Fc�AJU���{E�$��}��[D
��q���I0F��p�Em��׼��~��~�U�z�1���������B������iGr.JjR�Ӳ���H���'f�!َ�����ԡ����]qͭ�r��#�+�.��ޔuN����%ga~דW�4��G�ǒ�8��X��'�Ʃ�Ȳ�G@��n6���n�Мe�+��H<���u�[_g��~�UF$�#�_�t�a�F!��S����e��K�5���������ȯ��=,厛�=eRC��XH{�LG/9��ok�G]�s�ƺ�&�Rbu�z�k���`b���8����0/��Ok0r�ם�E��z�@������>_!�pA�|�O��a�V�>�������=�]��%oX���/w�Y5MA= ������]�Q�O���b��x��g9�bZ-�D_>�;9V%۹�{/�E3���eWCu�Ą�;*�.������}\Kq�V�|�����e�vq>����Z��I��8MC���B ���+!�V_@�H~��ᔶ��O�=ص�ar��t�(بN�'�v�I�@�z#��S���o����v=�l�>���Sق%I�̕p��[t���̹�(�A��֔�ܓ�8�Y�)%����Yf�B#L�g�Ҽ\��CM��
5Pca�mͧ9�&��X2���P}���Qg/���А�}���;�zSNL�dh����U��m�loP���8�l�9!r�.�]��R���CbI�Ջ�{����[Q�t�M#X��w5:UĬh|��.�^����01��Y��9Њ�h�s�'�1>�p��Y��
�03j�;�u\���<�K��c(s��Z���^�	х��5�V���b�1��/�����fF�N$+28�l�Cz^ر����<�@�4f���#.A�M޼XVj����.K2������x��eU����9nC4(k
�r�Ce�S�YZe�v�/-<�eQ���f��܍	����QU�]s���ê)sKQ<I�V��.���-�<L�{[�7$�
Ę��n��t��tު�3ҙ:.R]e�X�e?7�lU^�3���;�M�	������@�J֥<�{�;�3��#2��d^���B�B����g��	������z`S+�ͼ@��l��Ox�[K[��[�^���xK��k^��q��:t�+<�˶WFb2t�ʩs�Ԅ�|�P��N�^��L���C�[a��I�M7y�K��TCI�� wIƻN��>��^�4t3f����_�����r�+Y=�-���}�Lp8dz�-/��f�P8wN%^KZ�S�7�dBnF���k,cݫd�Y(ei�:wm�Z=��]t��\������P����z�n�=�2���ѧ����������)d�F�_�S��]��v(ɨ�_m��Y2Q�\s3WMژ:Iy2w���Je�:_&7�Y7E:[Qς��#�<�����ә�8���C�ޝ:�z�n@q'�H�Ѥ��Y �gS88�c�ve<Sm�1�6T�l����w6��Vd�V�!�a;�*�7XM3DD�B\g�0�b���i�Q@{�	���!��s�tϾᓁ��3{e����8����d�H��$D6�d�Q:US�)Ec4��#���^8��4�!���Z�1�)$�j���Rs�CMMv^)w׵���^�V��;S@+1���	]ޑ���������|�*�P�/���C=܅�6�ڼN1j�`Y�漮�ظW��g�-����Q5��#zm1[[8N[վ	Y/��L��l�
vx�`��#1Wm;~�>-U�Vc���^�}s�ӎrB&=���ȴߌB�J��C�o�De�^�w���Vi��#��N�°F���\s�h6;3a���%��=��t��M!�9]�?C��T��J� ��:������)��78Vl�Ӟ�"�4�$�����ڬ�̜:®;�"6{�����ixZw,���9SrjF�`XN�)1Y�`$ɦ"�A��V�����"���<���e��]zL�5J�y�-|�������To�gTR��sP�/�7;Yh���wj�j����T|��q��!u��:������7w�u�:�1�R<�1<�/�EA+����>c�]aL{�bu�d_<Es��۩����b����G�o7/�<�Dd �cUR�>|�F���n��L����#�u�A���q3��o���件��g݆W�z:�Dx�:I�EW��]]�o�)x��3餖[��~��[�t�o�4���Y/��/���Uޓ�Pd�� f��Ǡn�q+g]���W/ݞ��5i��t"�C;����.h�{�n~i�y\�"��÷�@{vLc0uw�V��@� ����`��u�<v�9�hZU��_��dH��+�%�5���t�Nʵ-�p��BL�朢�y�#�lI��5�3��ڽ���x��SO�
亁s��F^��h��1���ЦpC��t���6�G�~�ڄH��.����E�Ǥ}-'8gD���1�ભ�r4��g�Lk�#SKG�XN�.��Y(3q5t8��wL�t��J���N�*gu�r3�@��������W�>�3�M��1�a��cAh�=*��<Z�ͫ�n@���L�)Gw��9,���p�Q�����=�����G�o6ā���z�x<�"�K!��wDw{s���g;�泗]u:-�\�q���&��{6��>
uK�MZ�uk��]���-^R;��%}Jɕ��]��h�bj�ݚ���Ҥ戣~/�3�&k�\�7+���U��] ��
��)�Y�h���6߬9�j���ŉ�9�6cu,Ln�5Cr��C��+[�w�v��c����5����ꏟ��%���^S��&��1r�X�U~��N[���ˠ+�z������Y�DU�N}�k���Ω��9�1�*�-^��]��q;0�`xK5�)�45��e2�وm�q����7um�q�����~��kK��Ҿ���x7��צd�+֛Hޛ��}��c;+X[�]�wn�z��
�%���uϟm�2TXI�>��J��H�Մp+�B���x�t��hov;.�����L^g�܆��=,�󹣬Mp�I�K�C��VZ�����Տ���MǛ�e���j��7ń껺����_�{�O��4E4�+�N�Y1W��ᚚܞ��{�T���{f!����%6��޷=���ŵ�\3�!��:�/�4�u���f�3p>����VOqD�#�"�ױw�Q�Oc�:o��W�Y��ԏ�=�����r�S9JK�xc��R�{d۷ڑ���҈v٧ƍmo|�\�s�Z�X�k�u�.���%�S�j|����ec5b3��p;�� ��l�PC6���\ۦ$w�_i�����`Vj�G����=�Gl��>
�|
���mvTՅ�s�����G٨�zM�M���P���PCiT=���J�]�g�z�4��w�W-Ts���Փ���Ϣ���>�Ms�=Qf ���$��_F�7ti���Sa�̬��Й[Ѫװ�����^�.~>�/�}w���Why`�J��]�G�[�� �qx�1a&�D�%BCʂ|ll]�E�,�2��b\��^r�m��2e�'w�o�k&��ζ;i���H4�۪�weZ'��E�ƶP^�Z���&��w%�Q��u���Heg6�r!hd��C�u���)E�;�a�w5"�0`ȝZ���LӜ����Y�!��ީ����ZsA˗�2���f��s�i��A^:i�X��W'�>��ȧ+��k�cǯ�A�nMٓ���t�^�0� ��Y�ifH-S4�2��]&����;�z�Un�/����o'��:c��
1�5#.:Z݀�eh��������I���C��U�t��l�}l΋0����"YM
̗Y�о̾d�5S(�q#�Tgsx4���^ev�{B�N�)+�[H��]n�����Q]N�R�z��]�\�b;I�G���B
X���փ=;vջ�V��p�t��캹���0tC��.=2+�qwo�Ӡ�<��J�r�SrV<��#�Z�iZ��n��]����9G,C˘b7O뢶���hn��Pe;��;�T��m�X(ڭ�;2�J}��Ѱnv�	�l�T�ok)�����frK�	|����$��41X���Ww�}��`
�C+��%�3V�s�{q�{���"4k/i�k�d���w�).��-��=cdP�W�0)�� ٫�/^sTAw��e��N�귪�".����Ky�u�vgn#R7h֜;([��G�Z��
�뀛ࠦq�/���o*ъ㶻;�wʌvֆ��W�!���=�&�hH��B_�]�v"�Ε���ow93���#�f�I�u�Փ��=�Z[X�*�]x�W:SsUa�	=�٫b՘���h��l�ljӂ�c����G\ݙ�������Գ�_ѽ���Ժ�-���	P�}�aucY%� λ|i�;���ɯ���x
�zU��|ٶ0v�4���os'�бI�z���[�4�[[��nf�}�M� b�x	y�o��e��ܡa2'H�+Ms�X�[���m[yO�%����q�]�(��thG�����7z2֫�ۍ�b��}Z.�&�ȳ��t뗋�]��.U�^Q6R]݄N(xvX�S�K�\����+�'32���Z�fk�l�w�T�2�ĳ���ʈ"�"��«R������]��Q"=J"N{��f���֕k	]�Ȭ�^��]r���q��ŢV�䃻���w͡AW)�F����������w4�B�R�r�p�"N�t������H�u)q�uss�HW=��m��øE��.�xwOv��`�hT;��jӹ��'�w"t��N������u	�"" �YE�d�h��Uʲ��wS��;�VjD"U��ࠦ9	��Y{\��sw%�ZB����NI�i$�Fj�:��꛻���q�S��w%�+7]��ub���[�Ju�.K�=L�!Tt�;�s���pr�\�C�ʝ*B"�3�'TKQ:�\�p���d��D�,�XR{�E�\\�7Ue��.sT=��sB*/"D��4�L��)��r��u�c�z�d����qC9tɕ/���v�U�ޮ�W�'Tҥ��F ����mr�k�<$��d[x�e�Ӌ73�k4�!��;�޼l�
�pBD�?¶���/�vw�<ݏ/�90�y�c�BO�ro ��t����ۓ��<G���~F�!�y�ʟ�����o����>�z�ܓ�>� !@s�}�l��y+5�����Gc6���? Q��AI�.�&��v��'�߼����j����O���]�=�=��P<|�W���9�t;x�����<'��S�{<� �����_tY���1��o8<�1�Uҝs����ϼ �Dx@}�����xv�o߯���������o�N��t���oHI;��<�~�'rO��}|>.#nv�}O���q�O�'�}	��Q� �1+>�cC����~��a��8�@� ��O����}c��� Y��|�
#�Bpy>��#~C��.��>��'��>?��o	�!!����ۓ�s�)#����$�p��@���>�w���EE��5��0�x;z�_�G���W����w��o�^m���v˿&�y�o\��<	�>��� A��x���������i��\>��>P}�/z%a�߻����w�j/wv*��� �HG�X��!�	#���z�»۴��<����n�u N�z�H�G����0����>��Ϋ���G�>��O�I3ďX�� I'�=������j�o�Ő�+7�|4���~�0�>D�������ߓ�r!��<&w�>�{C����<&_����y;�>��n�[�����7�'Nם����.#�D{��<��j*l��N�1Y�tou����=ǌ�}�����>���|N���ǅp.��ޓ�yC�k�o_ ���s��?����zw>�?;�S
������o=���ߐ���n��N'y���>����
���_|��S�߬��G������%�y�zмH�8�����?����@����{���������ù]�$�����^������txw�(�}��H|E
,��˽���_e���{�~�O�H$#H~1�'��N����n;rs��Ͻ�;��n�㿃�E��I#��.B�����i���+��N�}��{v�󿝯G�7�v� �'н�#�@G������)��OL��Ðd��9�L�,S���4�M���t4A��-
<������γ�C)Хr3E��W:�J�B��͇+�����7Y�z�}q]�Z{*�Z�ޜ�T���کKP�}�x(H���u��v��a3\8m20��Qt+�{n�(��v?A�x#�|$���s�<&������.���m�0������yw�k���Ӥ���oiϣ����ߓ�O����?!�0���[�����9���� �/'�nGcw�︻�^_l������#�#�!�^����z@=��:9����{��|M����q�<�}� C��S|M����� q�������@�,c�?O
��uO�_v��Y� A��@Y&������nC���{:�?$�q��>?�7!'���7��������e|}��a�y��K���t�nӽc��������7��}���|�5����8�޺�#��L�#�j�7��?pzw���]��P{O9��&�@�(������a�l�I��M��v��=�nw����7�����0O��ʱ�C�@�<����y����s7^\�辘��Q'�}�|�QG{La���<&�B��;��1ɤ'�~?x�yK�bw�}C�۟����9ӵF���`S
���.�v�2��i��>#�^�C�3f��w�s꿬�}DY��>��G� P��}#�Y�d9���ݼ{�L���{�� ��]���-�z����#�^Hx"=$cBH�n{�b~'�nNM���w���Nȏ|ě�q�q㫷nX� �3���̛�zNC�k���݃þ��܇����990���~v����8>��7�o�I����Q�!�����ǔi8��<?]�7!}��ny��s��˕"D�ʉq���W���i��<�!���<�۴������N��>k��/{����ޒ<ϴ��o} T��;�o���90����}q�=8������7�?����ݼ�V�x���Yd�C_ZV�᷷����6G��������;�[w�k����V!ɇ����㷕w�iރŏ��?;{y�S���o�O���<yL)������޲.��G�����^�2D��*t����7@�=���T��>��_0�~��&���l~��xv�i��S�r8_IɅ��������raO!�?&��q�q�͎��'�t �G�}�`�O���G� #���gt�X�!�q�1����%5S[����wmk�=�zr5�����ם�]��=D�D-�N��*UiR�SWpIj�����]�mvp�t��������#\���{��$�`��"9-�}�dܾ�)]�C*�\H���;��؝�ܔ{��ڊF�C�}� 
o�ϟ|����������I�7�����8]��C����yq�Į<���}NNCۏ!]�1;���'���0���y��yw�}C��緅>@D{	��?(�b��k����Ʊ�o��ei�:���Y |B>�g���;rnO�c��K���w�o(xL>/i��c�zw�����nt�N<����[{w/����<�����x#�|b�W�@�
#�Jgq�ϳ�'㏮����n�������C�����	$�Ă@��#�G��{�L�������ܝ��<bw��n�������©�?}���o�r�����]���� $A����F����v�~ͭ�ܤ��_߾~��o�'Ӆ99\
on�/�o)��x���+o������o��f�*|H�$��D��h>g�P�p ��C>G`��qG�>�4�����@�<
�VF-s��1�����߼��i���.Ϩ$��>'��>��N<��-��ɿ!>�Ǉo�������<���ﱿ�9��������x��p�v�l)�<8��W|�=${�>"|�'j/��>������q_z1}D#��d"�$y�������q�ՎWo�r�~���z�<?��}I��r|~;s���yC���_�ޏ���=&�Z��{�G�}�|�������M���;s>����"���Y��: �<�������7�{y����zC�������9�S����s�8���w�ׄ®�)ڏ��L?ly<�;þ�Ss���v\�#��O�ޅ�b �3�>X3������ �I.=��=d#͠!!�ە��~���(I����׿�|v򛐟�}���7��ϧnN�`�}�:v�o��xO;�;�A���G�$�nY�z%��r���/�Y��x���Q����]}�q��0S�G�G�>�,D�>G8�~�I>�4�q��{����e�O>�~�I����py�o�ܛ�z>Ǉxv��	�^�#�i�@%c{y�D�y��jv4-Ϟ����yEd��]&Y7�{Nq�į��)�'��>���<�!�����<�oH;���P�����\{Bq�������0�����Y~>���o�W�]q�4;��XA7��S�:C4D	=�m,P��i�*ۖ�*�I_(N�um
0Sb}�S6�\��W��AX�mS{���*s�S��g��v��)���K�����b��}@�hA{��������Uǆ`Z�f��t���-M�o��p7s�5�fޘ�{�c�B����߷����M/�qG�xM�H7����o���]�÷����z���x#�^����|#�}C�M��	��/���_.9ߓ�~��.���s�S�uG7<�W���5��tbj5����]�y��<��=&��A���τ��C�o	�0������7�90�O���7�9�|�w���������@�G�޽nl�O����l/�}�"I> �;q��N�|�(gt\���������;rw�o����|v�o���^yL.��Q���.S
��|�ɾ���]��=��}�����aw���>8��!�=�lr��i���z�S@"<N�.�r^ۿ��R�e��u;���2 d#��>�Z�z���H|���D?w�ߐ�v�{���s�;I�?����y��t�����rs��y+�3:�L2-�4���u;���,\�jgM����j�1�ly�]�m*�E�rK�@ܮ#(sʣZ��]aT3�Sw��-��;\��1���p�?}K���ꗩj�n�j��uz� <B����]��P�Xk%J�'����3:�V7QX�$1�E����b�z|a�J�^����<�]@��Y�s.Mn��ޜ��}Ӫ�3h<���\�7e5�=���������,� �oMM~�_�J�������>��oK��̓�[,��Zg����W�#����Z^N`w^��#�θ�>�z+)�d_D\�]dwtn[���xa���ذ����,�o�+�t�C}k���C֨Tv�f�l�6�rƙ;�r������E�{%�ޙ��BfH���C�vCV�<��엚7�N�w�9X\U&MW�	z�>����JH1�<�(p���U�[�"+�]#�{5k�����]";�eM?ggocGkq�`nE�D��d����LV�P���ⱋ��պ�A�K9~����B�,),��$]�@����֥'p
c `�3�}�/I����OVq���8�q�J�b�y��0��3��_h�d���K��Vs�V��4�ǣBmi�C{w,���>���vx� 7ջ��]�<D�0�Ha�Q=^(v$g�kػ���;�ҳ�����E-u�䢶װx��LX��ԟ������� �{Q�A�H*[��f�z�]�:Q7i֫���Ʋ^:˚�}X�WQan�HP,�䧛�&�:v"�	��ݨ�G#�\��ڲp��{q�y�����cr^��sy�,�R2�r)��Jw��p�<h���OD{
<ԅ��p7�8cMQ��T/6�l���!yl-�++��41)���:��̛��I(��6;�e_t�
��|2��A�=)ymF�~��6jX���k���,�<e1U�5w����u<�mK�^aX}Uf��"��`Y�Aڳ>��ąfGC"M�kz^غ���R�Κƣ1Mo���������ˣ��e�8%�죜�=�w�ͳF�{�҉{�ۋ���*��c�-C��Vp�s��M#���蕃�5f�'ֵ�9v��J���!�L�,�N��x��� ��/^�V;����e�Lk�7�D�%F>=���\/���E��|QVlķ?S���a!\kr��R�e]^�g�nC/����y�xuR���y�^�=&���͹�������s!U�Y�?��â�x��Y�UGr)T�
a:X��9�/l�%�r�#Aː�V���>�"��7���Җ�frT��\��t�xƱqo&���Oj �X���4��\��S�8�q�fS�oUBÞ��
��:&�c!��-��㽠%�nc���R��7�\�Fؤ� mR�ex�V����ٹܽy#_lܐ�G$V�(�A�KcM�Þ�� �z��>�a��'�eOl'H�P��;�I�J����W�Ƭ߯80N���;��T|��͑��}ס	K��[ci��/y{��s�1��zvZI�*��Aߍ�jA�̀�p0t�T���c��MD�=�;{�jT��N6ً���w!�7(3@'R�fs�:�z�P�Ɏ�<���8�ʽ��L�trf'{�
��܍F�
���E��Ҥ�iŐڴ�l���	���	q��]�_@���䓆�=zqW�������Ev����к,WaN��R�wpPK[�&�tm��Y�Jp�.;�S�+�ɞ���GI��cC|ě'l������y�NID�G�ᮼ�Go�te�p��s��&ӪT�!��U��r�,m���W�u;n�#x�WJb��������	`ʈ�!v�7cw*ũ����sCK%�乀zl��H囼�������^�HT�By��+Pf�vБ{�5��4�!#_:R����Wu5w#�{������é^�vQ88�ʡk�`�t�]X��z˔lpǛ'�{�̘���[�����'"+�	�p9�*�J���n�1��0��l�!�d�gtXE��z��[���"�F�A1-��y�>�9b��Lki
�g��@��#1Wk��>��&Cǥ���Q�8�>���K�T3+i� �'�P�~�>�^���Q��6i��؝�f&ީ�c-���.\Ϊ
a�\�d@�d=1<�K�����{_Ej��)]����My~�c͞��t@���KY�!�[�p>�.�f����q��/ ����R��u}�J��OD���S�4��P�IQ��zb�h�K����ϯ��"W��w�:m�Y:�.C���_���`��3����yT~�Ek�)��i#�]�:A\��X�ù@��꿯4�`JkVA;{���#�8���e����>�S�D���^�C|�S�~�7�J�y�U�
�i^���Q��5�[����Q��}�#��҇>g��[]Q�sN�S��Fe�&�k�ոv��%���.vP��&ǥ���WN�Lg�evc�����뺵.�(���Fjuͳ�'�h τy��hc-"	![��F���&ov7�Ո��+5zSr�kE�}nI�T��2}ޓ�Pd�� f�8����v^u�m��sdz�[��~�}B
kuo�@gp�yY=�D��s��r@�O���TK��i�Z�b����/������(j�E�Ν��M�iV.�a8y��}���S\{y:�5�Aid ��Q�b!#���|���i^i�ol����qsQαj��p���[�H��~�P��ш�cm	�� �h���p��O��� ����S��b��y�̞Iߋ�N;3�&9�y,�����틵�Pf���	��go =��cu��!��֞}+�6�<g�2q;�(�t��M-���>Wx� c�ӯW;�t�շx�����-�&}�r:���_k�\��qC�U��] ��Uv�q+0'Q���{ol����EN����0o�`�^ܣ^��X�&�k�Ϫ�mF�nR0֡Qh���JZ���N�R<�P���8i�j�5QXv�)�t�P�ON��yA�t�e3z݀����/(�0])F!���׍��z���z�\=�ufdy����w��Ɖ-v;[�`�]z�u����������mZ|a� Tqvݟ����w�p�[�����jB� �A��Ю��54��8��}a�e�������t5jg���N3�s����Yv�ƀ�eW�i�Vn����+���8�s<C4�D����?8��/��M��x�̓�-�\{�<q��@������ ;��ז���Xh�Y�ݎ۽8C����n9���dk���S9��ܶh� 1�'�������ff;f��<�פ^�hh+T�:��\;]�^g����㡛ޛ�=~*��
G^�.p��Ӟ��w}��������0�;�LKZ-<O����b��"�AB{�9�����Ѝn��K$�#V�e>��mL�N\z4��f��F6�|/w �.d98�V�._p�}jcH�f���PK��bFRױw�Q�v8Ӈa��t7u�v$�D4�{5�yF�}ꝲ i{ƃ�o��A�z�=�bB �s��҆u�Gt�k�Q�|����<J�f��o��P�����<��np��؂B����#�!��xѮ�J��S}�5�4��!=�wT�*�����.�	b�Y���jp!n]oC����摃e�*.�!��lp��e�Y��nGǩ�l�z7�F�9�G;*�oYy�8��f�[�U�1��=�y�J��aW�"4V_>���殐W�)�h���7��\���P��E>� �˟c�{�G�8S�nt�`�d�4x�1�����8r���x��\��KFA��I���nl�1��Uxn�j����D��)[��0\ɺ�I's�,����2k.�C�{\%\5�ϴ��cmzD;�f��W�R;�s���8N��as@��[y;'�՜��@�DWJ�`Aڳ;]8������6Y�oK�`��0�]P�t�]�è1�W.���@��Ͻ�V�r���j�4��~��w��c �n(�vd4oԄj©�z�>Ps����T��,�
Z��}>��4��,vs[�e�'�n�Ηױx�"p���納{e�m+q���z*{��z�l��).��>�=]~�s��7.i𧓽�$S\ή����I������י��#2��d^����j��}��T]��/\�H0��0�D�Uf�aw��ˁ�<����J��m�Εtq!!�͔��`؏�����p�\	բ�G���\	1>�tϨcx�����%��S�y�Ϋ`��#��l#@E���k5�S6C5y�u1��{�M}"�N_,g�{7���j�u^T�}@���mI|�fO�~}��b+h��[5qZ8���,������QǛ�6J}r��f�/]a]��fؑ�wS�Y�-��[2�/�����&�3�s]v���{����=l�������em�A�F��Li.�AY�� :���̙g��c��b���㇧F+�L�<kJ���f� ��Q�u�w-eZϞ^�=�dl�z&w8��\g��4��M�%������+:?���q�f�ˑc�����m�6����}�n��6X�zH�Z;��y���Hż��6���Wa�+Z��f��u�4�w_fq����/:�ӊ.4	 R�-s���z�q�)&�&hKf9Eh������Z�V�2��t�gY.3iV��ɶQ�p��^M؅�f�!gw@��f�G
i��8{(�hk���@�Ɵ�c�U�]L�I_u`�T�UӼ/��na����g16���$��Au�]*�t�x)�2�A�p,ј��/^ɪ�����{��VΜ����<�=���^�a��3���q�b��|��a�(>VJi^�A����:��Cc�cL	�X�4���)�
W*3��oA�xh�S�V��vX�F<�75e��EZc8/�;��R�V�����kͧĠ��t���h1F��.�� ��:��HR�c㸔]9�U+Uo�� 5���H帯�W!�G����*���,z�Nor�������>=����������v��V�|~�)�BY�UZ!���������Nun��ˍ��P�a!��y�2�Mo�[���]�V�'ݡ�mo'�iĞ��^m`��K�_9��қ�rbWȫ��f;�H � ��|�ţF[�5�:��nK�c�N�ս��ܷ�U�7�23��́�}�R�0#�k�����|�h��I�w����\Kns�œo&�%*�����4;�Ļ�b�g1ȍ	�ā�{iU��4���X��rV�On���Q��|���.���M�
�1S���B�7F^�����F;d�J�8�ůŔ��e%`ӽ�[�+���Kz�qo�[��*��ΘF#�T�C2�Gk#��yذ���u��c&�ڰu��� x�����1���U79���	������`�|%q4S�����$M�)�t�"���n�������iy��6�}-��;GGR�d���%ӛ���;��ް�Md^��y��!�TFS|u�f�x�Gy� �5����������s� d.>f�v�:k�P�l����%�yQhJtm*����L왢�Y���50D�Ň�u�םz�a�hDZ�+�)cngRY��5�a��`%t��#n0�'*�S��V!��:c��;�3;s������yP[�|Q�(���ۡ�������"�za�N�Q�usr�z�U��q�C�=�4�]pw˞g��HS��=MwO%E�<n����u�˹�P�jIY�8������7hxe�x(� �x��;��^�䊺V.U�z��Q�$��*$!&�
�B����1L�����R��r\�Zd��^��TE�2��L�2�J�b�V`Fb����:JsZmKK�3�6�Q����ʬ�����@�E�Dx��m+����l�<��6N�)ȫS�%���qL��8t��wwp���tr=�;���(�T��xb�y���fnn!h���囮ZtE��G�9���A���wU��D�(CI4�,����d�E�r�Zi�-�/]��J͚����Q%;���QJ%憒Zk�A9'��"��^R'E��K�VK3*��L�"����"����&r%Z��$��*������*�1:�JVf������J�"FQȶ��^����eK$���衕/����w��W+�����gb��:�*��Y#�s9ćN�La��Dc26�6ub�� �R(޸�hWig%]��u��x'���M�^9��tN(�{�;l8�h#�$��W ��C>U�el����
�6?s!�'�i��*R�o�Ý.Jߓ:U��N��nS��
�q"u���Ύ�S3A�n����vzn}E������WT�Y��N�mkI� b�;����3J����KBͽ��*�mߡڧ�ڧ�7��+N,�Մ�l�nl�$G{��0KHЅ^Z�x�%_t����Uع����+W�9�:����r��!��qM&:(�z^o��:Ԭ^^����P�+����`�,�7�بf���ƙ�$k�I�ԏ��u���ɱv��2^���Iv�P�l;P��SKd�{$�!1�"�A�bk�_3f|]A��ʇh���I����͛��gIȆ�L)� c�����I��c1y5t��Q�=͹4Ȉö�_p��ʈ4X97hs�dW�����1��*a��4)��n��1�VyVsRr�9�߯��{�z��;�f���C2���K=�,���T��������(��W�lз���7�s�Fe[�ɑl�V��˶��ʴ���4�f|�^d���vѱO�0ĺ���-�d�v��H��I�58U��V��"/z���ׄt�a^`pڹ9I����ĝ�O���.ةffu&d�F���GU�����)�Jf,�҈���oa�O�i#�R9��}�M��x�#r �h;��X���}^�}7��S9o�5˚����S�� ����>�/3b�{V�wVT�V��n�>�m�t�w��{���Jr�)�6\~���RC#t�3@��L��OI���Q%��N�K���%}�>�}�tB�!��r�����
�$v��*� H���[�b7E<�N�ب���(�p�X�n�˪�1�[ՇC�u�'��μ�P52�Y��~� �3�~��_�u敤Fj��s���Q����4T���`L����-�rOb�{(�s��R���a�H�� T�eF����K�#�9͚/U�>�5�� ���pH�nQ�:xl��A^����x�s���,]y�-rD�x�> �ZFC�H��ӫ����U��X	��*��1���#7+L�]�]T��cuMA��������b��4'�3t5C=K�{7�Y�ΙZ��6��G����[,�(�<j�τy�t"�(p��@�cm	��R%v�N�����7ϑ���W�v7S[����%5S�q�#��k
]ۈ����zC���3U�/@;�������{�q����;KU��\����$r���uNǹ[ӕ��9�³�1q�\wu��o6�B}��Z��NoD�cWP+��f����w������N�t� ��s&<�CI�p��~3�'�@A�=��_!~9K:j�ԢR渤.��d`��q�}�4�]Ȳ�wL��2���'��N'�A�N׌���+݋��իϔDvA<�e�h�9j�3늻�n�a�0V��zA+s���!����a���뾩�$3N���/�V<n(���O���َԱh��Pܮ�rA�،彳"2v#tN^t&r�����jZbТ�qi
�8��=Bb�z|cSJ�׳���}a�s.��z�^r���*\ϲw%{ *f�~�q|(��ٮwU>P8�!�����OI,���'�8)4j��Zi\	����6�æ��o���k\Ǯ��t��1��4��(�p���j�2�o8�=,;��q���<S'H�\�7˛��;�F�s:Y��>�ذ����yT�g�{3���%�De�F�M�U�N^,>g���!�l�f�\ۊ��r1L�JF���)+q�n߄�5�ɀ�O�wT���OU��>�X+����@�SY2UP���z��U$�ׂ0���W!+�����B��%�ֽ��te1��d���E�l�(]K�FV�)C�K?qJ�֯l��93y��y�ly��E�=�q^�탠��qI�A�Az��U��J���%�>�Ҽ�EȪ�7�8$[k��������+��:�<�|��TW&	:m&L�*AO�z��J�J}��׷�ӊ�2t=����1S�q���+~�g֜GK�M��(v$d%�b��Tq��:t��tSK@d��=���_5��᳖��9�Jې�l�k��P5{g�1!5�e
���'S��pr��s��Gf���p��x�M�%�d�Y�����Ѝ^�S吋��R�Y�5Q}Yi��͙�/M�'��D�W��eX�:��<� �%��S��T�+��{+;<rpTݧ<݌��+�ܞA��;Uo<�7� �,iJ`srN�̛Ww�=u<;N�c�W�����`4�B��s�����u�*�v�f˕���8״��^� v��ӝ�j���$~�n��/+)P��E��	�Hv�0,�
���`Sc���m_�{�a|Pmy�C��}��/jN�{�'����}sFN��C��dgݖ�+�:�XUntUUQ���K�/sǛ]��/rC4P�@k����;����}uS�4�1��_�>�^���GZs#stM ,g\�J�׹�`8�XZ�|9.��X���uө�4�W��G9���Ֆ=z��"�`;>O��$#�ط��\s�s49�|��iΠ��dl`u�m�7q�לºǑ��Z�{��gj�s��띌gq�G0ZeC������}�U;͢�Ǉ��Fb[p�$���;�_gj��z*W�މ��i��tY]In��~�y'Iݣ�;j{��ʮ�~y%��{z9�����q�fS�u�he����z�puݱ9���p���K���ݮ�_/nk���.'�ڦ� M�����q�hfi-�7w�(ϭz��|[�A�x	�>��Z�L����T�wޞo=���S<c^���N�y׹������������cܱ%�q0V�D�;VxmT�o&�hٚ�n�Xk��뻙0\di�@7r�hҽ	�*�9r����iC���8��v�{ow�#�m?=�X'�o��w��0�'���q&-�&��$�ItX�I�/�f�6��w�P��op�q:�D=R/�O��w.8�V�͕C��&���"�f�q�js�.���P���
�	�ܴ��ج݌Q�aԅ���r���3�8����<w�q�Ț��^�,\KH�ꀱ���ٳ":0C;Hm����s׃�33xg��.i]5����o��`�u޾3Y��R��z�r�.tt�fT��"�c����R�|˾3�i�j\7@~3�ѱxs�#tRjޠX�y���ٱ����{�vڜ��z���f�]��3�wˊz�rV967��Y*7����w܎������͜��,�ʕ�����BFC�	H��h�첝!";dY\<F�Y]o��0z����AP�3�d�MnL�~i��9�&� c������T����!��m8+0��֋��zu�f��z��^77�D27��ji�c�)�yS�F�?��6���h>9w�]-������5����U�0,�4�6�2���K��+�H���/My\0z/|]�8�p.�j5S�+��ҕqe��b��;����h;1<���ҍ{i�¬']������������HkGq0�K�A/��#b��=��Dq=C�������h�O�r��s���V*jq�s|��*ւ������/
��q��I��W_zu(��[ّ�"�ĺ�Ӥ6�Y�:�/n�*���q�h
�~�V����R�k�9L���#sloV%�\fL��bn���1�з$�P��Dƞ߬��� c��T�����k��Ѥ�AYJ�]P��J�^=��kE�l[�{��oG:�:�T�TI�0x�yr���*���aG]�eӁ�]me�U��VS�KL�F`S��ο����v.���e,��kz��4hn4�!k#�9\��R�CD�(E#���GY<&5GEg�e�r�S��C۽Λ����p�����鐚��I[��/�L�{����^�v��I���q0@ֲFt��V'�P��Uytw��2E7H����T�u>4�3xs�����q#��Dú<A洍�j��;`G:mgrΉy5��^Q��{�Mfo+��:�!]K���\�#�6��jb>U�r�����w7�3���3�8�BV��N#�G��~߫r�G�n�;��Baap����Ar�N[Fo�����O���5~��l�kI�.8�Ϩ�p\�H*Z��C�O�Z�&�8~z'p����~(�#7�Y�7�R�h�29�'�Q&�'k�=��Ա�!�;�Y�VM����Pxo�f�3�p}�N��W\~�ΫU��$�U�r���s&��`h��;�_19��QE���v���"��َԱf.i����t@x��#���"�{��){}*�D�"���QT�$-���BՎ�ճ�O��z��t�#i�"��}�4Vf�;ړU@1��,74wlwVr컘�^�	�(q��q��ٔ_0<4R���!u�L�>���/s�HH?l��+�*��6C�~Ww3�Y.�(=�y�^dnj�k�3Z!e�mӝ���<�M�1�6𽡵�h�Ғ�r={�j棫�r����s�j�kT7Ss���q���B+��:�*�h��g���2��n!g��x�簞i}�lQ?	˦Qp�׉S)S��u�7&4U4#��=p�lG�x�\;�v��w �/n�(7m�^��Fo���u��Ζr㮽#��-�� ƅ=����������z��Q��3T�`�S}�C�S���y���k�}�����}��T�Kɽ�
�k�i)2��L��#��d�Z�����֋O��8qeDD[{=�d���H��O����8����� 4��;T��tz�ڙ�Μ�kME>���B��t�0���*�r.w^�pqm\3�!��:���:9���(v$e-{cTq.e�L4�DIy�c��]���'�Ư��[�c`E�e�^�-�=����F��Z�}�Y��T�򪓭�ow38`n<t�;ϫ����HP,�䧛�&�:v �н^:	v%S徙�99v4l�I3A�#7*���[��3��R2�t�
y�Ҙp�6G'�g�Bνhv��ʫ�{����٩��0Q�-�@�l�&������7�W���}�ҕC��u��e����ͺ�7Li�Q3B�Q��|2��g��!]`;�R�	���Mi�{W��ȝG��y�"��#/7]�4G�"��]�+�>�!�>����*vǏL�#�K<�1җܝ���n��y�>Q��J��+u�|��+5CIb)��I諌n�~����N�TW>���p)%�q�tmp�< �kl��u�f��뎻��O
^ô��^+:���d���?<^�A��T5;Qj���jmz@Aڳ�щ�dqvb��E�.gv�w�т	�rW��c�O���}n.������$+�W�9�����Y:�O�h�Z�uq&F[��{�5�V�z�[蓺�=�􋪘5[,�P:�R�!��bz�R��2�w��yÁ�|���"�0om#Ce�m&�}���ӷ^��)�6�a��y�wk�y�+~J첹ף��͊��eb^�П��4���;AƑ��G�vg�S��=��r���9Z:$�I�O�:	`�����9�j���Vy�0�v���o�[W;ȹA��(%�s����������G�S�A�x	�>��Z�J��+������h��T�>~�-�ً���W���L�Y<����k��d�09bKeG ��C�>U�S�w��.`/;�?�z7c]Z��v���p͚����cF��p�\9Ӡ��&��J�k����[S�,��=��(4O,X�8l��bs�������l[�xS�A��A��o��^�\n�fYYֱn	���V�=��ń�s|�I����Q0*��Sb�ޞ]]e�Xc�]t�÷�����r:��j�7��(�w�����l��:\,9��`�i�����"�!�OL=W��:u*�rI���j�(��&��1��^I'�~ 7��P<]h�ڶ�T�}�����'seP��	�6�xuD��7�"�ސ���c�;�(� ���N��6.ǱG5@bԆH��r�p4�u��q��&��� ���̚L��`>O��*X�5�;6dG@fgi�֯Aj��cN�"�:�)���
�o��}��BFC�	H�-�n=�S�'���Ī\�e�yk��h��Y^쳻[�n�u�^�C[��\�=#�2ak@^:�*E�K$��3�Ptw.��%�
{����qy�c�>�dv��q�^77�D2:�RÁ'�#�pmT�k��TҜ�[~�;N�����i����N�q�"���5^̭�l��)��X}R#�Z�JT��77Ls[����/$�O�E��M��0���r 
ײ������:��{[�}z^�����ji�¤5aq.�_kK�؅�/c�{�HQ��8��9�\R�O'�Wd�S�dĉӊ�����p�ݧRunn�i�`��B6��۲q�ʚ���K�d4`�n��&��Y�k6<E�;�x��<����[F��U�m]_c��uF^\�
V
*4f��Jń�_�ĴOM�i��B�5��jw����pN�oZ�D�v�Je�&�����W��GSIݣ�f�T�u��n��:`Q,W�bq�N�d��ϓW��c������Ѿ�Y�u�O�����z�N�����fb%d|w�Wnj��Bw|�ߕ#j�>׫���P�yRO���T�8^�mn|w�����8AnF����*�w$o�]�Sz:�>��G�#nT��,s�mIt���s�=��;v��:���4�oo1���j��ɟ@/��ϵ?�3E+�u����+��&:��du��=��P<��L�a:BoRQ�h�萩���ܮ�>�4�;��ti�Nґ���e1��u����B�)��L���lm�Tpfp�+�=g��b�����T7j�ƍ�F;�=�ͩ�eu���4^園�ba��7����Z�%wRM�ھ�����v��d(�n�jOi8�4�ھ}]{��f�cz(E��`�u�����ij�u؝WB��oTi�r���󥭔����Ǻ�Ԏ^�@�l�O����ϱT�}��ӣ,��aD�ůX���U�\����d�:uV��}�u����>6!au���m��y6���۸�߳H�q:&�'����8�p��1I\�wmv靠­�h�X`��^R�@�.�ѝoV�NrL�C�����V��}\�50\��8�a:�^_U��&�n���V�Mv�nb�[�8,nŸ:e�.���'Eح��-7g:f�b�LέOK�#���h�:����U'�s0��k8 �ݠ;�r;@t�U�q�X¾�ޤ.��dJΖPhaݏ K9&���㒹�1��=\�}(���!���egG(9���)���Z��uMk�Z��V��b�eg$�W}�Y���f�.�F��k�c����6�:����[��A0X�Ի�ʕ]����ܨ�K:���Fi��'�¢��A�u#�w\y�F�AQZ����� ;��6�z��΅YΖ���!w���);�2�]�p��
ZG��Q��Q����d�S�@]p�6�y.������sW\ԋ��:a���Hm8*}���8�Ǯ�w�s�/C'���tC��ی}c��;e�x�b�\��*땄�<�����ocH
,�˲3��}!�r���{�!�>JV^b���5i��.Z�����C�mu���h�ݲ�5��ʷ��� Y� �A�ww���]��������L���Q<�Wv�TH�d��\t�T�S�O��r�3�wLm%w�� ��wf��Nm^����Iت�3l���F\��� f�֮���.�c�.뒾�EQ�u�PIۚ�Va�ۨ!s>ܥzwr��%���I�>'�h* A3Ԏ���aE&�#��s˥���lҳL�L�CLڑaJ�N̉DK4�£�5=Bsd�[X�n�D�d���j��e��@�-3����R�Ujd�z��YrԊ=]"�rB�/v�FH��d�]r/i�ջ��t
�n^��I%\�V��B�q7<�i
�^�N�V�rwAK�+ա���^QR{��"*l.j*IԍjҐ�W/v�P�2)�6��\'u�1��GQu�PU2N�l��J���g��Y�Z���2s���J�$B��JJͪ	��WY�J��f���J17=�QU��!ZZ*+*�9[P:�e�:F����bYiU!D����*Y2R�J��@�ID��J�$[0��V�����P����h�g*�Lf�
���Vs$ �ea����L�Z��3Z4؊�R��)֎�����(�%�XM���Um9�DæF�ӈ�I'"gNEI��U�IJ�	 A>Ȅ�����ي��\�*��Mgt�WK�sP��sa��39ܲ��u���Bv��fR��įGi���	�w/�M����W��}U��z4o��c��w�"��S}�\*S6�+w
�(<.�^���q�1"b����uv^i�~��L�a�C�6��N��	�0ۘ�T�##���,�����۫�^c\;����PTB�1�:�:�&�0��nI�μ�Ӳ�W�pp�� �Χ���ȵ�8��9��z�����:(���tsm�v�\�[�z֋{(�s���� �Ȣ�t[��t��Q)C��%�L-$rH�Y8�j���"����Atw�pH���GE��_(x�'ju��(�S\�� �#B8�"]����3�P��;:�mRA���"h�Y)��2��r�q]+���Cn�ꚃ]�O�Q�b ���-���xp��39K���e��/'��z����̈́�Rj�B�.�\�@n]��-���^����Yj�#I*6=�h��]���k��c���cӯ�����'�>�`s�#W%�T����Y�'mg��r�:ws_���W(i����`�wLߛ�B�'��p���ܢMד��q���ə�_��Z�o�[Lt��Xxr�a������fЮ�n4�+�K�A[ط�D�'��T��ѷ@B�W���Ņ=��$�3U �P�h2��n�����'�8N��Ök>`��e+ ���K.����q�nm;e�-�������3�����11{��4�*@���Cm�ăg=�>�{�X����0t�X�5�W��V<c����C7�Jfk."� ��i3�ǹT3[1ؖ-fw��3����w��=Ɣ�eɛ�Fx̞��w�v���v���F��-5���j�#h�>&m��<��ai~/<]��~��ƨ�1@�f�r���G�k��@]�*�*�<�'g���W���`T�)��'�b�֔ke�e��O�7s��nLj�I M�>�z�D�Y4�Jf�5^έ|"ߓ1�GWI/�j�,�-�v�9���dm9�,��G]z{n`�h�F]����&�Έ�=���%I�VG� �N!��S���õؼ�][��祜��q��=W������Y&�T��XRX��@��З/d ��4>�z���đ�n#���қ����{�^�5�#KqӰUˁ'M�čZUx��و朸�a-ɡ'ѱ���yn&�E��Rx�}���pqm�}Y�r8��0�HЉ͒���	�wگ	&���}S<��.α�1ʱ`{��}ʇV�t�8e��ڮ�m�nӃ�v��{����u٤�
,Vʔ��\���Q��7�<��]�v�KV���	�=z�).�#�^J�	���NȬ��wt3���Aj�l����T��C��]?x{���n��Wk;����^d��~���E�G��wR�n��BT���-7W�^0>/�Y��poK�����H���B6xo>�%��h�S�np��N�PA4(��gn�=|����y~�G�.3geW�v����:3�H��C�<��N�r�8kǍ�t��m^�����Υ}}��֧���7H����vk��T7c�P�y^��H�#�5�+3�sH7��ɛ�]�q���0rd�t
I@�lO��>,�p�חT3;p;lԎ�2���u�t��x�V���ݟv^��N��ei��fV�U��V:Bՙ��N$�[��;���]�w;2��q&��/l_k��PyW�4d�Va
�	X���B���<�˂9�}}��/؉�eS��22�C5�«^�{){�n@���ډܳ�I;��ؓw��u����M�Q�5X����<I���F�\�ҷ�خ}:Ey�ΝiR{~�����]��4��@�>̖��#����`�y&�S���w^gl ��4���C�d�e3�3��v[�pi��KM��C���Bm�9�PP�(`h���b����ڥ%���Ams�.�(U��E�UE�-fm�pT��ޱYϻ�2Q�j����U���c�8���9������]�%��:3�fk`�Ӡ��,&s����3Y2�4)�|�w��J�zb82b$�=X:SKڪl�����lr�OF����u�3����^��$eJ��a�D��z<_�� |+����d�ϑ�)F�S
3-���n�L��znNO����v'�O>���&��$q�-�w�$�b�ݨ��:�Զ��Q��GJ��І�4�g.�[Y�g�����0��7�&#4i���p�F>�� �nI��S��>�"�����At~ә�z4�~T��c�_�N���赛��������ƢM� c�¨����ڧ�g�7��"��.���,4(��l�A�:���Vz������N��/�($	^=��&b�w�9��!��.WL��e�X27qv˹ǶpQZحI�͓=�PHk������H����xLh��m�7nc��{N�VM�Co��m�c�^97�A�� ���7�����gV�5��m���6�o'��w9��c�G6N��t�gn]�ɻ�^�����27�];1٦�`�+U�������!Ջ��!�;���D<8��MD:�o����^��{��fF��,�vV`�ӛ��b6a|�7
��j�Ʒ�$ڧ�'o&s5e�B.���) 7�gTj9R��M�ޑ3wk*g{(?� ��ט��E깣n����mՙqKHX�q2�eo�N�7����M��'�{ܤ��E�I^{�� �ܵ�S�:��B�ԱiFCi��2�u��}�is��gX�ޖ���n�$U����3X-Z�i�)<0&.��/m5�=�rj��ɾ�M1��r��$-��w!uG�͘qrc�����4;n�������Ջ����1�)%�H�]���]7��D��!uG�Α	�Jt�l��p���l�q�NK�Ydn��%��VP5����v�w��9�S|�S��������©&M`J�27V��EY�L�����;�ت�Ok�e�ƻ$Bջ0A8$�����Lo}K^�fMX�ݵZ�3u��Mt�Gc����p�ܑ�{hG=R�����*��#�+[��ꡔ��f�̸���o�a;��{���F������NP�� fo�����޽#`��ۏs,Ne�*C�RR䀎�8��m��۾���ӕ�rϴ�y`P�z`ZA�n�VfpK�1�ŗ���)u���&�57��圢ێ��Tŷ�9*����Y�`�Ć�+�!��Ҭ-P�Wr��<rv�۪?3{��y���4��������:��ّ͛�Z�z���(-{�ө;��ѓm�Ω���Wݝ�Ž.�uǨ�7_&�J����fgd�٢�nj��.Bݹ������2[1-��t[�ǨG9�q�Y�Գ�D�ڄ�-?sc=��ςi��Es�s�Ƽ�b@�c�@��:�;��k�7L!��#�޾o1�(ĝ`�d�u��X��{`Iͬ<�{g?W�K�f���Ǹ���{A�|����Aڧ�V}6��|UM�n�9�s���2AKQ�t5�۬pjw�'�4?2��������Ëj�z�R�d���������w�*��}��������)���Y(qʿN����Y(m��^�`H�~w΁���xΗ�ˎ�~s�����,���v�f�e�ɓ�sa88,��K`�j�O-g��-�9ה��Z}MN�^Y2fu�#9`����9x��
.�\a��me��ax�,��m�y��\�� �kf]����8p�iҍ�=HT�U�66��֐�f�2�+yY�Y*C���Lۨ�I�h	�{%Yk��P5�9M�B�vB�6�aMB���vi�7|��� xy�޽�O�&��,�����h����t�bn��}um��h�#s�֫���v��˿y>w�S=]�b��H��>Ʌ�~}�'X�ȣ�z��6(Ê�r0�,rii�e�<��f�\�!�n{jy�{P	����V�����!���^n�m����d9�'�}�4{���h'��xd�⪓���72���[�%��+1�'��(s~�t�A��.22yE�q��;���qV6�g�tf�IgK]W�Qy�J�X)IR��h�*""���ެ���ǭS�p�7�͙�|�H��:�JZ�&�fˁ�roz�8���]�ce���'b=��.��μ�7���sS
"�(`���ˌ{�r�VX�c��c�w�	��>�Ȑ��%�6?o��,y�E�����}���8�|O�;��T�gEv�K��z��p.���{�~X�Og,�5ti�fk+p_%(2m[T9L<�N	��8	����0D{�}�u�^�	���t�+K����jp%�ꚵ	�r�4B���8���jP�}e(*%�����*�GVgn<7 �ydWEv�a�?�=�����S�̹������Ӈ�/S�@Nz�Җ���a;�S-v�\��k����_���/x@�z�����>�׵�uJ�Gח0ˬ6�;!�*H��3��#K�$U�$�^�Z���l"�ڜ;LQ���Eҡ��ܡn<�4�}��U3gУg�%����̈́�}�������Y�ߖs�ǐ/}K[f�˶�A�w=V�_���v����
[�w��/ g7��%�X;n�o\:����}8NBa�T��K�N T����11�X2/'#������ձ� s��] ���' �Hź��F��Q���n@su{0
h'��t5��c�E=7��h���VSvV�mc2��7��}���D��s�.��Ǽ�ݠz���M��a�jzʌ������Q��H��Dݳ'[��o��o"kΫ	4����v��;���Z�pDhh�D9P�.�
��|��j��uj�����4}�'���f����T�feC�#�%Gkq��҄\n������:{�{���r��;���������tR/'}��KUpn�����dP�E���;�4��j��sї�{�����u��?
�r��G���|p�c*�/"�{it��w	����~=0��/3���P.���6y`:�N.���Y*�y��%Cn֦{�����[ى���[b�����e��2С�ka�0/�:T*��ͥD���c�G62}�1�5��X�/�"B.�.o��]�������֭q��v0�@w=�ᱶ��l��:�����xl���i�x"�.�S�Y�.4�B�mKQ%R��!h�1��m^��B�T(L�G�Z�4��?Y.�7�kKCV�}��![�6�����=���ܚ�������c�ʙU���B�͐!Ņ��ȣbbKBSI�sxv��=�t7�t̑Li{��Еo�����>��چ�Y�FD��ӯz�u��`�k�{(���{@9ו�ճ�j �&�H�9�쳗��s�)�lN�r�reE"��0M�ַ��H۱j��쎲�M�#3��:x�:�&O���x݋�O�#頤v���U����}0�;5c�R\B01����ޭÎ�t�|�sn���zU���ƌ�"O\���b�{�o{�`���VV�3��h���&�%v�>�p��X�i�5�5z�l�ڗx��n���fz|��kGǸvwy�z�̯W8"	׷�ed�}���N��=o�uΌ��f�wٗ@[�u��C��Y|vY��x��޻܌���M��3��z7٤1݇y8w&ٽ,���^.�9
�◆aU�U����-�N�����8RבS�lG>���ɥ�c[��ݓ8m�x�}�σz_\ds��k�[�v�ɾ��]pƧ��}��v��D�^tj'�n&�l$C18�}��t[�H�:n���ʬΧ�[�ړ@��eϓ�}�3]�o�$��=�S�T���9l6�;`=��+�!yR�lF�xy���7�iv�5;�:f�O)�
�+��q�Q����Œ<�̌t��7��dCw>��9Y��x�@��α���K��v����3k�u�6F�B��lMO��Z�T�B�V�K�7��r�%u�"Sh�!�y���)�C��J.��g\������="��̇��:�&襪��rnۡ��_X8�v��O�o!9E�no���d�;���-�'m��Ս�v��,��V�9Όf<�c�^dց���o�X6����|��F "��s�4Dw��v�b���V�V��|��7k�k�+�ʑ,�{Ko�u=��\|�x4&T(q"��/�U���p���6��6�m�32�*R�b7n��2�	��E��u�q]'\�ޛ�1T�VrP�Yʱ�nL鮩HgAnϞ��B�Tx ˂k��v�.֧u�.T�E�B�X���A\|\����U�z-��w��Cw��+���Tx9-V�B�;���4��|���zt��rxH[46ͤd���y�'\��E�@Դ.������3��6�I��TL\R�Q���ۗxn�u5�b�ҘjWv��՝�u{�^f�̝�ٽ�[s�YU2��\o���sh��Xj@w��]p���4.���r�*��xV�Ƨ�[�p#麔�&\JTģ��j���4�V�C�-e�b�Զt��r�"cT��pR�DE��ڴ���:�S����m���<Y�u��-%Ә�)M�n����v�*n��s���|������0+Sq�����4�qu�9��2���vn̎� �9����{�]h��r5���I��r!�R'}ȫɅwHh��ůpb��ۚ��c�&ԴMN�L9􆯱�ɖ.���[�|�S������ⶺ:�����>�3���-�[�C]� ��ᮬڴT:�\Bu���WyI_6��g:U1�јsr��wE�;m�ô�j�Ӕ� h�튛��4m�_Ws8kM��u�}WE��n�kq2��]Zӧ+�&���U)��mv�2�#us���`����/�<o��q_f���MO�R�0{��}ԁ�,ne� �u�ڢ5�׈�PS��&��h�����Tb�`�Ӗ[r��i��8[d9�@�V��셂�;�`Ř�7��@�nv�i&8쑄�d�{d�V�3z�)��pVн�ufWf-+;��cıí�����<S���1�0�j\����Զ&�X7�c���-�u�[�
��%�S����t�7Kg�|˧+��;78�Y/�}@�4V����r�����%n��λ�t�w�1أ��AP��(0�+�=D!���#/.��G�dB�Ug]>�n����u�x�j����\z�5�m,�������]m�XZ�Q=3#���s��k� �eѧi�s���8������;U-졆j�vS����2P]�M��T����.�T�ڢ��^t��S�m�n�O��jibu�*��B7XUkAu;�u^��4SD��n���Yf�]uH��D�K	#�T��aR��"l�.&%�*�ws������!zh�fbz9��8(;�������5#�wIʌ�L,T9���Ш���r�0�b!��asB���I�U��y*��e�i�J�!i[T�U.�^�YDY*$��+B���Q�HY������29�����J��O'r1D��:�52�t���IUjHDr�B�C�e�D��Α'�9�*�*���UH����LٖG��z0�ԩDDBCIR�*��,�QV�B�٦bX*4:�J`�!��劥Qi�s$����L��$+DP3J)%�D\�A�!Ҍ��fd�а�K� �&(��,�dr��a��aj�Vl����T�Ql�u�#3YF֦�(�U�TJ!�AK$�:�3�F�3Q�(�IR*�+6r���Z a��*�t.\�ƨ|I�lf�#�ũn(�it�����\;j�����a�V[鸍�Z6�H"&)՛Fu)ک����6�����v{����v-y�n#g欃��mF���YpfD�z�a������Uyz�;{���������e�<~���l��;[5]�Hʝd��'�35���GMM��y��M�~��VQ��S�ˍ�=̦�d�X�mp�Ԏ!�l��s�{3��6��=��X}��y���Z��F�0�7SW��;G2C���'	�O��t�O�t-�qۉ����Fӽ�\ԘՒDno%{'S%5���UG��o4uZGՏ݂R//�Q]�,�c�[��ɾ����} Sr9�ey�6 ��̀�ۦK������hB�&ܙ�c���R�df��$����D�I���}��w���P�/�>V^V��H�8sd�f}ͪAm���nӚG,s�3M�N�酮7h��]�0dv��LΜ����YњQ%�bL��sv%\uK�#T,*���TC7�X+�����0�o
;6�wr��s3qt�R�D�:1ս�Rt���J�qp�Z�xeXI��e�VRgo��0�okzZHAg!����x+S������k��\�G��$&��7�s0����]���b��a��{�{�ʻ�nޅ2:��7ށJ&\�f�:/N����g~U��[O5'�\,#'�þ��k>�/*o�X�<��s��>O�=�i��N��U8��(����%�1����g�{Hd��e�l�;�o�yH�9"�o+����ѣ��9�φ:Q��'%��^�@{P��2�KZ��}����9�~n~ڦ�zp�s�{|��yl�T�qA�ss�_sȗe�N>���1�^Dn�]�ף�޾��r^V[���F�]t{���}��k�7r�@=�UP5>[�N�:I�Y�V.�n�1��[f��{���I�ն���hq�p�uzC�j���-�{O}�4oqz��f����yr�7��	쪰�pzm=��ص=���>��]�k�ٗ�>����z�֨���|'	�M��U�e�x�dBBQL�x��#3g�����f�M% �[��T&��4#{���u0�G�RV�n6�v3���.��qϻ�I�����Gm�}���aK�v�������@�N����oV�ߩt\D���[Թr}(�L�zu�5?�{��31)U��,��^��gckƔ�YJ���wV�d�ϞP讐`��9zE�w�SZ����
��d
8�jA�9���^�;'������P-&�){3�z]ޘ,��g����go�E�h{�Wo�������P�z�o	�t�-u�͂���}"���Pt���o>�/�d쭚�;�^���v��m܄����=��Dm��b籤C��U5s����uV����m�t]q��_GF�,�V�*c��m��9yɹ9����.�[

Rٍ%:E��sLT�i�_4����C@�.Z:v�9��/�Rhݸ���k�F�J��6�Ĕ�'ڢ=���;�e\뗼��vQ4��o`-��������˛���ׇc�E�R�c)B��+��cj*߮L��r>�w�O-]b�^��e�����0�_U�q��;�N�����ck�c����VVu��cf��fԤ�����n��a���%O��W��
j#׃M��3����Ln�L�u�&u'�%4�Q{V�#3�� �R���+4b���lmv*B�IצU_n�b�*9��_7��ox��k[J5��ڽ�}��䲢)�H�~C��Q]�.oVv�� 57�����ِ�|�;�׵�5�okнD��ɶf�.�bz+--�7E���Fv�1[��^rwY��g���x�,����i�F��0���z��9����-����5���5�R[L�VS['l^ې�L�	���5��]��I��ܘOg�<�Ƀn�+L�գ���|��ۧ��i�
뻆�v�QB1�J�Ѐ/5כR�A/J���G��H(J0-�%ˈ�wC)�ܹ�td��l.�˵�
Ѝ��(i���b�W�dML�n[�b�5���I�}�5�݄<���E
����f-[=rx��R�}�x�ήwfy�sZ�zƎ�8^���:�^�Nx���H��Q�xL1��{�j�����E���&�Ƕ�{NM̅mh�惗��u���%
c��2��"{��|uW]�n-�-�����5Vޕ��A@vg;��$�Jvá�Wj)�t�y��`Y2�EmϥM|�z��X�̧0�P9�����H�ZDk��p9vU�q�����n�9zC]xj+�J����1�N�s�������*2�V0�Q>mE:�I�S�cb���R�Ӡ,v���J��K�S��q�ٔ<��nC�9���v�/vh�Z��';<�U�K��Q�!�jy��ŵ|{s�mb����ڢ��|��/S��T���Q+[�n��|�y���J�c;�VȆ�D�v���Eoh�Y����e��1�`�����UO��E�C�k�m.���$�x��2ڶ.�򻶏n+����c0���?z�3յ<���:��$N��͇����t:܇�O{���[l�礡k�V��O�<�H繕��Z(��v�e�{Y�Ux�m>�V�ˀv`���'�'C����g7������B&�cE;���Z�%/$\�7���P����~[(M���=ئq˳m�"u�sH��v�y�����a8xg�ޘ[i,~�|2X�Ϋ�t&���a� �M�|�y�K}z6�+(��]�����q5{�ip{��=� �~�:e�ŧ�qw�!�6�P��Z�����Tָ���|��W}��������o���G�+���K��a�Mӿ�:��T�v�2c;��b9$/lv�x{� uf�9���*�1ոr����RcrV��QIW�\��T:��v��!j����ڗ�{���r�adKU֛Gq5\���JI�ys��4�p!\�uS��	�<���FNc������{�S�y��5��\%,@ms�;z�v ��z�)>�v:�h;6td�D�ċ�/i��V��{*D_+�?�MF��|KZM��l�-�D�^f���'N�"F�P$J��hY5��r̳�l9:8��债$�]�>d�2�zWo;w;���1�ǹ���c�r�o�k�9���F��W����;;QVn�QD��6�ĔB��s�Q�g`�dN�r�Ժ����=voaV�/T�6�T�-�n��eͭ!f���:��o���l��Lȗ�}y�L�`_�Ӑ�LS�1�n���9s��!�o_>��蠷A�PW�`n�M��t�h��W��ƴC:��7;|)7��6����3z��� Fqc�E���ۥG�k�q�wR7j��+��ڑ��l���W��z}��ȹ(��K�k���V��ۙV�u�X�ч��(�	s�c��v��8��ܶt�z�K�ﾯ�����7��ֿ2A�d�_���z�Z��͑Ӑ`�$#�{���Nt��rim�W�E�����r�9��[W�^��r��~��;X����c��$���1��˔!��ɵC�X|/җC��FFnP�f6b�h"�Z�n�Kk�u3�f�B;�C�4ۢ��{��>�3:���K��c�v���M�l7v�^�Ee�5�(��-�6�'w��qL-'e�P��G%���!I�� �u�L�P�;$S�x�1��p���뷰k��Ga����=�#n{h�S{����v��]��ὸ�ުLV�rʉb��6"q��V�{Aٳ��Qi_lN�mC���c&X9]��]ِ9�r9k����퓅�bDv;��wڶ[緱�tuֳ��o-����|�����zR����?��V5�ה� d1��r�E������0�,T�zi�2鷾����i�e��7բ��ަ�H��=6B������67�R���p�=W�[�.���.w�w3��]2v��2q�GXz�e�
w@�ǜz1ԫ�/-}�\��7�'oh9���"����0M�W7��oNi{M��[�2`UT��l$9���s,6)���Q�9cP��rv������9��z��M#U��6���$b5��1,RlT�"+q�f�b�%��NwQ^}�~�7�e��ћU�KV��U'6��퇟�ـ�n���CՔݕ�u�=h3����x��r��Z]�a�ټ�o��OXĦ�nd������(r�un��m����b�$������ȡv���n�(d��t_[�/nÜ����8v���e��uB�K��L��܏֐����{#�0�������gK�w\��}�'U�STA�o�J�8�b�Θ�V�Iӷ���E��LN�F�-6g���[�����]Z&]@��ۛ��϶b���.� �s	쌞�_t�t�}i������F��qV]d�Z�5U{�zn��0���<$��B�{0�<#�T��x��1<9/v�gD�S�ٰ�<t��$Bb��eucOk�gݬ������o��6��Frm����%�_]�ϳ�Sk_*a�VR�Õp�ݦ���iN��}���V1rɿE��������n�>9YWY/L�@qB��T���t������f�v�j�w�o[o�KN!)k<����-'tǎ�N9楖/p�YvVǑ�w	�"��}��^H�͸��'�}�A�{��ީ�m�ȱ-��<��[����HhyL��Y�-I=ϡJ���UWN�	�a�7���_��Y��t�]���E�.�uǛ���\���}�+0Fg/iP{ũ�����ջ#�mg5��Gܮ{�ĎoK�[�T�qB�V���:���K�A�3�@wO��=�#]���Iy#0�=4����nI��-��;��5#��`�]�ݮ�-s��{��~�ܻ{hlYe�<vI�l��8�|O;��J�c;�d��C��b��޻�k3uwV֝~��˛uU;=?T�/M|���H:����*�7b�T���0�f>nu�p�$�ҝX���+sϡ���k�������J��a$-L[��rի��I�'�	D{�43���,�P�~��tz����qfE��f����r�}�f��w��Y���c�Ȕ���`W՗u��2��j���	Ɉo,�ЎփD{�t�[�gn�M�F�D�Vѡ�7E���g#*����7{��y�ܤI��YD�����9������k�oi����a��{�%���nnq�E����e���CKik��ې�shC��2x>��m���w��-&{��o�Eig����[}�ѯldc�X�q�`-�,YRA�YEF�5��*�Vda��uX�n��[L���1[#��H�'	�H�����g29v
E��ެJ��ɉ��V0��[��{�����c�`�Pñ�H���H�k�{�3���R�9�J�f�h��kɧ��n�2Y�s'ҜYw�^��L��a��kOn��Bov��{�9��z��W��D�,����](go�z+�{��=��j�}�7�wX�d�P����ɘ\I��):����yV�o���Δ���L�_1=��k1K��cN5SΞ��b�8�嗠�`�X������ۇ��йDB��%�2�n�t��0�T��j����&-K{�c�a^iUԷ�ή(�:^>F��#��r��l��Ӥւ�u5p7!�#�{�{ύNd�3o���R�ty	Ǵ��ge�\FS*EQ�1���+-�]u������� �:����M�}}Q�x��pѲ����둧�8�]���%�v0+��j�|�T;�z�'r�oeA�\�D�s�-wg<�r.�uP��tډM���.��ڦ��:"�1���v2��D��ڊD[�>�D
���[�����B�qC"�&� ���i�+�W T٣��К�b���D���/Cϒ�kS���ޖoP��+F�1n�^��9}es��C����-��-Ȍ���^.ٔ��Sr���d�Uʱ�u�x!d�Z��uu�-���'gw!��s��W̴cm��v1�oE3��H��NvtFo�O&�`J޷��9]�ջ�r] k&�.�ɝL�*��g�(2N�3iP�`���q۾CZS*��ƹL��6�s]�a=�c]N�5�\��me�}�M��Q�k%�w��j�R��Sna�k���Z~��;��_J���9K)!3ĕ%��m��ަ��"H
�*�o����䇣�]V@���9%*k�1�9y�K�&<�U��2E������M�;T7j۽��i]�ظ:��f�S�]��΍԰��w��ݗFt{�ң;A���
P-1on��9��*ӎ[W,�p?u��U�(rǵ�U��͗rgs�"0����޵�p5G��PD��D�S��.���۷z�� ۷Lt�31Z�h����pDre��g+�f���Һ%I�/)��Y�#h_
����(��v
Z���L@�	�R�x':���
�*3>}m\�YkL�{�n��*��s{���A��hs��t�ul���5��u��5��r���<�Ҡ�A{̬w%<��e��6��u���ː~�[�^�AB��zD#��2�o�w�d�hh*C �B(��%Zr��b�r�2�+ofGM���)�EL�X����e��^=f�ȥC�l�i�6�׌$On�G*T=�Mt����S!�No^
DJc��&GBxumekǱ7z���)�I;o�I.>'�*ޓF��:q��×��m��EL�l&%��V�	f���c�*/7�^��I)�����s%t�KW��f�qI��<c�Ok��	ety���^ag>�V��}]�x���d|c���i>�n����lʢuj�EA&�"W�XHY�c��TF���Wp���ҷ�t,Q԰�y�u-!7��������_.1U�K�e�)�o�\y;��2�`Jeh6��x�6T�����ڙ�r�K�	�Co�ה>ӠZÄP�~o9OL=�Q��ۤ�ʡ�S�/��lEL��N��?c�S�i�9��K�}v�����U�7M�[��d�*0�����h�Dl�6�Y�T�"+N��A&*$D���t�Xd�����"N�%��H��R�YHJr��MR�Sj]--��&��"(eE�Tr��4�UA�&��Q�Qȫ-i�r��U���R#DJ(��Q,��BȈ�Ce�UZ$,�Z(��u#�aF����HTT�˕Y�UV���%ʃUP�%,�3,�Y�VU�%��EuB�h�J*.�	U�Ju�*(�-���VQh�EFq*�A�YЩT:r�bԐ�,�:.U�I�\(�
��Ե%)J�S1P��I]"��R�K��J鑂U�B���B����锚hl�EhAI�J��gT��JBP.TAqDB�����T�,��*�T�fb�Q״���Y������*)��$��X�ܗ�6��7qGwu�.����G��@�Y������U]���S������ڰ�[u\�_׸6X���i,Ć��C������$U�gYƹ�^P�b~�:z��f��{T��1 u��#�$>��c�c�Η������y�Buۤ۝�U���fyy�T��˛t7��{��ʹ����wF-\.8���܅�.qps�%��ϻ~������\���,[dN\)ك/z��'�N?/A���F�����Ƽ�a�Bz�:�����
���|�Ƕ�w�C^�H}�-Ч��C�Xs~�bګίO)���z�JPS�	W=&z#K���E'�R�Q�̯fold�}�f��a�^�uG�R�=<&ព���Ʃ�٥�g´v�6�ӝy]�;it�p�c3��k�{V���W����׍�t��>��h���;$s眧y(=��a{%��u�"n��2v<�#��B��ڐ���rUcjdr����x0*��Z��c�~��L|U���evzޘ��^�Hm��ժ<%��u�R=Œ�m���o��Q��s:��vm-P��箜s�T��Xd���8!]֡R�3�+R��},k�u���Z�<� ��Iu�w��7�:�v��O�y��mX�[bMIE��UF�zt}�`�g%<����ܝ�+D��Q�cE�F��m�:�oqd�1��y>���g����f�2'\�����pɥr ��6�6��uqL,�u��;��ݙ���9jG#ڏJv�OL��M�ͳn��W[�{.��wd���ٷ�'{_P�.�uǫ�Ў�5��q����X�[�ݝ3�S��1�7q0��w��N|��H�ˠ[���(�>����ձ����ڃO�s�*˺f�n&���T���ci����H�*ޮ�oa�܅���V�b�#߭<�[��I�~kW�ّ�u��6E�ן���4��)�����_�e�M�����3���y�������K��ѧ.,�m���M���+���*[U��߲�.�8����Q���E�Թݪ�6	��}M��]-Tb
N��iS�Kof腳�-G)\:�=X,�mр`�/�WxQ:�:�����M�����}�7�b�v���sUn#�]�9�ױ{b�Dc#!�aD���ʓ��f��=�r�^��GJ�j\��"��|L�Z�vR�j\�{c}�S�3��}���o��Df��H��W���跢��^���8��l�;�{bwY����퍚�)����j�k��VQ�0n,��i�T3�����,N8F�'^�R�fT�ה��{b��[���.��ȭ��n��0�4���%��&N?�b�{��.���J�:���fwDS���V���d����]ΆԮ�Gv�V��tR�,����z�3w���z�����St��f�\;��:�7��O�)	"��'�ʫJ3�P��oc�1�ɦ�Ϝ�ux����d2 H9{��$�Xod�g�ڤ͕��]V���zƅ(ID�	��٦��ȻU��`;�<i3�dO�a��L�Ό҉,�k�uE�U��3���`�cE�
e1I�m��I��Qy���Y#�\O��-�e�Q+g/`���sEH��h_oTy���=���Z����+�賜�v+G�rJ�})���:_7�9/���vh9Ǫ])�l��9o$P���y�P�\՛�rT�3@W�A��Z��Q<F�k/���Mh���Z���:�o�`sCT��!v�9��6"�X�+sk�R\-vPX�b�ٗ�q�;�%��_W�<��v{׳F�*�L|cQR1�07���$�Cn��mB�ͺٷz��B�tպ��5�^]*���5���8��Y#���S��x�h���Z{N_P��\^v��:d�~n{i�^5;=s�Or����on�5|.�s����=�̸���Owk^���1�^Eh���)OpV�y�=5��M�[Zߥ��}��uw.��OGih	�x��&9��Z���S��9��}K�=�c���v��Sk��(���{r��������E�*Į)�S�H'3�G葽��t>�߸�Q�'	�Z��^�O���A�)pS70q�G�/>���x������+N��O ���{{���t��Z��Oc���깑�E��W�27V�������%Ld�v���>ț�Q��������Zαڎ,ڐg�ND�U�j�v�^O����ܶ�C|2/"f��H���=�k��3�iȗVp��T]@��VJQ�'kF��	��b'V�m���* 7��+�-,�SaX�-�gr��3"o-�zq�5�lR�q%���oQf�+�>�l��-*���kNd*������e$�V���筆�z3_ʪ���ZX����6y��V�h;>��A�ޒ�}�7tO�i꘵0��u!k�a��O���������:.�?�"g.5+c$�ݺ��'w��3���Jħ-O���� �K���;.��~;�����)�3y,^�Ub�+3b[z]x�e�=B=��6yd��l�]�78�ZcFs���;P�����Df�x^I6*�ؤY�������Ys�*M�;Y��u��Gތۋ�x͛6i�S�i�II�O����E�b�6+6n$_���lx��E�3�V�S|�I��?�g����myhH��S{�	����0�R$���4�M�H�{>1�n�{�r�]tC�q�9ʘ/�<�*���w%fC�}�����_�K�ҽ}j+ao��=@(՞Q
>ǈ�Vr)DmRk�$��å�F��E�z�2�qk��v������ɯf��3FeJ�g�^ס��H�YLy��C�)��|�ao<~F֋�����	�m�AT	�&�D����)sFo.������o�E�5=ї����jD��Ԯ���͡��XvyƧ2�d�aﰴ��q�%���̽\���f,�Z�O:JOL�,�;�Uk�w�&�3�ˍ�{���o����FK#M�6}@��c��d��S�(�l��j��p�%�ʬF���z^c�L��0i�hɦ���Zd��+M�P-�j�J���W:���ͣ���]�r=A֙h�6ԅ&ND�U�6�GV;���Ԝ�g�rY��Y=7���ޟf�>%=9;,�rt�y�bL�OAޛm?z��ʿ5m��ۗ�-|������߮
'�*�w�s�.�F�wy�m�U75Wg��3{�j���Х	b-C���G1�e��y5�]Ï�og��E�[/��_ok� ���.��sK��TE�	)}�+j�'<��_��ظ�{�;�o"��e׋b��<V�Y���b��'��u+������=���i	㌮{Nyx׽ۛ\�]�8��=�B"ɤ�HiB�[Cm�ߍIt],��л�I����b����^��� ��*	�����;�c/q�1�\r��w���5����[ޣ�p��}4N���/�bht4,.�������_�^�i������O-�bQ���˞u�/���ҧf�;�����E�N��f=��f�g�Y��T���\owv���:s�k�-���uvygbu�Ǿe�xj��]�S׫�[=N����'�tY�w$\��B�I�i[#Vc*"��=܅��f�-�@:G����=�]�b����|�6x9��qw�{{4�gZ\���s]^���wIy���C�#C�Ζ��;��os?v�����S�����v(:�/j�v�8�U�2�
6rK^�ۤ�d��ʒӍo���Vw���f����^��ވ=�]���i�@[9%��&M`JŘ-�WgZsN�k݌΍�A��}����3�^�g01|z�����J��t��dO,R�ׄ�qh��?
��1��V�d��ƥ�Ow�mw�L�]��"n'�u�J��i�j1r�w;��+D�[t�q�My-I=�7�(A��iɥC\�is��B��^]�+{)$rf����r'����P�@��r�#�BE�dV��8��2]�GRn����f����)&ӻb�y�$���.����Ml���:�A�Ĕ�ĥA}�v��\4�
t��hfk8��ZhȎ�o�������ݸ���uZ���ݠ��Xr��yjI�aJl�26b*`�\�Y;��ԡ�x#�*�͝����_ ��*ڋ|3S�}�fW�����㮬zS��앜�ks������ܭ6��q�{1�ڳMQ�U��vuζ�w���Zt�ַ:�#��ֿ��ӫ�V챹N�w]��;�cG61��>�d*���t=<v�ח�s��V"���i�٨�k����%N׎&Q>VXd��n��~~��zYk�y�驣v�y��/Qz��n�,{�6bS칵Zam1�ڍ���}�x�w�m�X|=��q�����<*�O[0��^�z�'e�z���� �v�c�kcw���{t<�l��'��z���3�k�V���=c�
ø���i#}����J��}JI�MP��o�-�rÛ�ɯz�ŏWM�'�aG{޳V3�Z�,z����G���X^��˝���ot�P��L���=qTtɇU\������[�OV!]����f����N���P�WY�L���_.UÖ��b%����J)�ln�۰�ї6��w+��<6�-�N����o��]M����vb����s^>�>���.�{Z������p������]�'�/U4װ$�I���Ij��|b�N�38��ZCδc�c�Q�o����{��?��^�3�e,�bdn�1�b���J�\���P�٭��d��ƻ{���v�	�+i��)2r%�*�R9i��-{����k��u�ܻ�="w�X\=�g޹�L7�]�6��!����j�u���j7b�4�N��j{�R���|u��'�)�8ZΌ����n���enXR2e����vy����#Ѱ{F�cFsJ��C����1�]9n)�3�!�\ι��{�$7�'�ޗE�,t�\wg��WJ�9�e�)�M~5�-��geć��o&��`��a�-��#�X�7r�ä�I�	\��#=U|p&���&�Fl�w8��6����EI�U���N�2�e� e��$�܇���'���Vݚ�&�i)����*��Y�FY�lu��6���
	Z^m�qu�_mc�O#8mTn�����PDu%�^@$�K0u��IaL�
ܔfo<�Z�7��hE�nV\�+����@�)Q���KWmҾ*s�W>bȿV��-��қ�Kjo?E'���Ƨg����v�s�\�ݡ�~fj��ke�����R\���y���N����h��!���ͣ=�8��ݗ�:w*�v��^i��H3�f�B���Qak;d�:�v�B�4��rNݲ��L�
N���������ZZ8�Xr��:|m�50w�s��0b�mz�g���Ň-�{�s9�m(��\����w+�OE2�h�un�`�i�$�e��b���YLb�6�Y��6��i{ݭY^����w^6�ut��|-���� �ã�j�MU^�=6��c]��vޟB��ڐ���rUz"I���m޲n��������r�=������ݨ��?=��å��^J��<���w�.����٬���z�ٰ݆��^V�G��>PVo`����K�n�6/�-�¯�����m���c�N�����5F"�M�.��7�T�n�_;O�7/'nK%�� �8L�ѩ��ڼy��e�\��V6�ŻG��PnR2���;����Q"ؗKm��pU�J5*]6
}+WjGfԬ�5�h���.�G3#��
Ӵ��,O�Ig#�E��tF{���o F�]-tU��Ds�.DY��G2�n�����{i�-n�4�-*��wO����6�pˊ���-���PnG2:d���e��D�M-�0+'.Q�,D�E�L-T�_Q9fdf�£�RLѲ^�%��BX�V���[���)���ݰ���D��xE�߆�R7�f���n<{�-s����|/��X�E�[*w�˽�#�[�����Mb���Y��s��"��]3�K� gCpQ�	l*�Z#t��zȲ��ū ��:�Z\/k�yE
���% ��t�D\@.O���Ӵ�`Zb�pQ��u`/s%]<*�[�Ǥ)��GU���msCUYb�8*Y��:�s���oalT�Cm�vr�`�X8��+����h���,HzwU���j��^B2��r�7�+�o�n�0L�-و�)��Z7�HcY�mMdk(a�]��x��\̧u'b��m=(j��n\Q���He��==}�~�%>�J���=s�dY�.k=��'w&�����&�r]1��i��t�y�s��:�YA����i}iV��=ʏPㆱv�Ϝ{��R��4H�����T%�/$uB)m��V]��Z6q׸S"Ճ�췕��9
T���e��c7���w��i%'u[��M�8 <�Aq�uVf�#%�Cf�[[��j�P�GU�c��PQVS�!j1Q�7�'�u�ݒʚlr˯7�*����]�%Ns}�ގ|s�Z܊��8�֍!{��1w^U�t��k
��g�������Z�7k�K��W�3"�3�����1f=��.&tGvq.�������Z<��u��!Co��`r�-=Nļ ��	Bi��z�}&��mВU�蝭hTm���b]=�Z<sP�p�������mfj���J�Vf�ց]%=�w\rn�*	c��*�piࢻ���{0��v���o� 9�S�]��̑ɬK��3��
����u����;���ˬ��v&]�d���;��C��*���S^������D0��3����G[���Xkrf�M����lɁ<��`���m2�0>N��$�.wc������Ljtq<���l��]`��r+1�Knk�`��'e+�6w�5`�]Ɏ�2�4����TOh ��:nS���^��٦���״٥���/p]���αCQ|������JT�#���;�i=V�1�Qھ����>ޜ-i�6M6��u(Z�.U�O6��張iUϢo��+��C�-�fGˀ	S<��5��
uE�aﷹƶ���(��� ��_>��^_Ou9_)DՔ�4*S���.Rj	"��R�h��r�C��$TAAaӪ��J�+���Veւ���4P��EPfDQ���(1"���(�i�X�0��4e$�L��±hWj
U��L��$�H��DEE��X��V�F��Dh�W4�	P�r
*�iU���(!̒(# ���L�I�
��U��A\�����T
������
��36��QH�R �r�(��3
,�R���5Q""���.A��Zr�4�aTU�Eer�UG�-H��2MZl(�af�L8����(9QW("�˕�*�Eʢ���e��3#�(�鐔UjD�J*"�`��(��]�E-*(Q%�NjBt̲jr�D�
$�����Ihi&j�"(�I
Xd�uA:E	&\���ijB�r��̩U[
+0�BQ9!gQj�d'%0�
W@SZfV����D䇧�U����ٍ�wuײ�{�\:���r�5�v��j��E�	�:��ا����x��lVѝ�	�}�'w=��:o��B;����]���`�-O#�6knK�T�{�}o�{[��.��{#��y���_�oK�]q�.�{��c*f�h32��G{щũ����}OM����Ky�ܜ����t[�5�N-���ov�٪��M*��q��[�]B컨�q5g'5Z��������;;F6��NŽ�42�pc���c�c�����X��[��~�ꓛ�Jx�h���LJJV�S����흯<aĻ����&F�U#����R\����;���OCVeO@Mmc����V��,�ԛQ��2Yu��v��+��Av�F���1����l�^>xZ�W���j�1'�8v���[qn���M���EI�*�{�	�|�Z�]�b*,.pZ���S�ˎ�~u����;����:��grz�>C���쀝�BnG���z�fo��};+�e�T?�_K������2H�0n���ר�Hk�âL�<���R�B������9h�_˃��Gd��Ρ�{�_rǊ��'V7\�y��-��}V�V�]��B]t��w]'��Da�ӻ�ǽP�����Y�$vR���3{+��)Ft�igK����g3��]x������X=���&N��'�x�w�e��Vb2J������W�+xA���������V��)��>���'� ��oF����ؙ�Lr��BQL��<}����r�)�bN��5u½���/+Ƥ��� ��{m��)�r�p�ġ�sg��K��/u�H�w0��׵Z�f���M�U��j������ZLn�u���tx!�
%?R7�n��u�W���]�,����M:Z�I$Ml�mݘ٩I �����c�!9�<��v�4�Lv\Ks�O�7�}O���o�����h�y�]x�-׏P��;��\��@]� ��.��ņ�;6鹼�{��WLH��bG61�(��h��]�];��W�[Y/7��,�~嘟K��󙴔z���q�c%��9��:U#�$b�׌?;Mz�(�Y�ZU7�5��r�
�<�I]�Sϭ��)��"3��^�t|Κ�k���&��89a;�r5�޴ߍ�����5��$k4Y��R:Spq�T�X[�O�a��WD��=�Wt�Sb�OS�F6CXAe◝�Qf,�҈��*�K��k2��VrZ�a����#.m�އ��ƾ{
��Ȋrn'PѺ�5�c�n�ůt�ϓ�7nb�I��u{����tCí��I㝤���{OKӎv�׾Mv�Aک�KG����]�:������%�W~��{=�m�]��k����M�P����O�a�B���,�)��k����#`�-�{t-�J�����oi��S����|�Tw�3�_QD8{p������z�l�:�y���x������1[,v���wƫ6I�Z��o	�NXd�r��l�ʂd�cYK+#u�Lp��|b���i�eeo$���պ���q����w�R��t�A�u��o��1yBL8RN�v�7�}�8c�{��]�j=Dwa��j���|�hM�X����#
��9L��VV�ǖ����,Μ|;��U��0t�S��]ѫ�NSM ���p������L��ws
ĝ�b 1ѽ��u�gZU{�M�^(�)�̠q���<U�_a��s,�h�\�s��kO'f��63Q0w����oN�;y�`Һ��հ5�y�H�]�Pf�u�wJ��g�+gFGTڦ+3�X݂�̎nħ-O#ڜ���&D���#��Z�i'&V��z�{1��t]2�����,�
��U��z�Z��2l�%"Lk�P/*�d��Ӗ�b@��a�-�P�t���5	��R�9K���4��'��5q7g'6l׉S�i�II�E�Y�i�z��ԟR�}���1��x�n�;���{cu��.m�އ�D��8r�b�J���ܕ�x^,^��{�P�v�Z�=�B�)�tX�W��3ϻ��bޣ�e��_DmS�;o�}+$<���U��9�TKEE�a�ġ�ayW3�0-����|M�Z�զ ���p�3wvs=J���n�˩qUhV\�3�/���ק!�Pe�mX-��
y�RzR�Q�̯fE��b���H1/`�=�3�[
�
�@[�X�l�3XI�5�%��Vd�_N�zU�b:ݝ�� ����>Cup���&^4(gW^sB�����t��%���Ϧ�!��C�`!�^�ByhШ���j̋���5)��Wwp�OC'�H5���2���Ը ���
cS7�
�n�F;o�oN�����^���%Α�y�\D߫]������*1�&�%v�*��m�h��;�n�Ee��FO@�'`�x����{jB�'#�1"�����6�mcڈ�+�Y,���'Ե�J�����k��9:A���03%���7چ������1W��7.g�y��l ���%U�̫�@Y��]{�W�L����ݦ^uY�~.�χ6na�S�G������p�,�sV[�b��؟B�u���'�u�oK���m'g�|;tB�2r�o4E��<��#�u<C"�h5�v�H�HG"i��~�J����K�S�rӖ�j�nn&W��@ɻ�=�\�2U��H�u��;,�h�r�le��xd�K,z��k�ZΑ���&��(�{���R�f����u���{��q,c�2��h�ꧧ0d���\1��S>K��GR0�n���׵��g���[���+��<��r�Q����q�[:`�̶��*��v���#��������>���
��fIt����w�}��q�V�v �<�ڈ�t�52��es(�:ir�Af摷91;��=Q.|!H����r�	,�-8�r�N�;@?=z3��v�ɧu�_B5�v���w�u*����7���:��I�,O������{��}&w
fܣM��b{CY�i<����wB,W�������E�Q�i:���v�+)��,��? e��>6����:���O�l�k`Zv���\Cʜ���coY �F�b4�a���&�pS0�.�q�;�YT\9�]\�{�{�«j�3��LԎb2����S�h��>��ܔ�n#F� ��Ĉ�eM=2E6җt�����A�J�Ȫ��P2��D�s�Z����r7��to����º.���i'K�{�Q\�ѕ��ؽAx��I���v'�오�wae������^t?�͝M�c�G>2����P
YF�f!;�d�b׈�i9�S��#�5�
��o�e�Ɗi�駊ԫ���h��t6��y��&�_XQMHa�>�g���R�֌]����~�p�kc�M����zz����H���>��^�A�«���{�������F3����8��^ �"��.���;�'�״�WF`�]�*����eP<Z�0�*Z;�@"X�gE����dC�zD�X�C��ʓ�y��û;�9
2)�2=�����oZ���}�6��	&� O�1�D"�[����'�j�񺱉Ezނ�J�j�D�Ssn�x�]�3��bP�I��s�V<��s:7_Mٙ׻���nڋc]p�9����]4&�>g)�6���P�z�=寢��s9�r3wt�4uu�W�GDg����H�iFMn�̙
xnB�e[|���1�3c���ё��\r~�w9����e̲���F��*]g����P(0�=���aR侢z��۱�)��YW�5R)��w"�t��[!2�L�� �@�3��Wu�5&�Ǭ�:6��i.��zahǩܞy̎���YL�.�!���OH��OL���3h�c1�U�܇�y�b�/����e͑�v`�ǣJt��Oۓ6��T�-�sб��<m����8�K0d���Dv��6]�XO�]�0��/��zn{E	S�3�w9|k��L�2�����^G����c�u+�U��r����lz�2Z�̳�H��C~��,i��pP�O�b��&��o�Rˌ��w;2)Dm�~��I@�uKj1k��6ܲp����Q~'��n��])�o��63��Þ��k)B�g{�GlAu�����M��Q�ݶ喜�h��� l���h��dH�U�{O�$�X� ݆2a�E��t��~
������7m��"�6!	�s:�I�:�c�����8�AVn:��'wG�r��vlm��8�%��:t��=y�W�mtω�]�aO�6i��נx�[��8��/lGY�(C0��LoT���g���;��IyO�ܧ�<��ܯ&�tn��#�T��X-��Nt�ƍ�+�ܣ���I�7�U��8�5�:K�mT�P�D��b��׿o7J|·C.Tݳj[-�/��^��aփ_3�%�h��9ݜ��t$b��KGR�z��.�}=���n�Վ#�)�'h�f���/��g\`����op8JϦ|!�;�����Ȍ\e���N�K^S�黣5i��d�?r��n���)��C�t�x�QD��wF'à<4%:��h�{x|��h���+��*����[k�� �+GpC�q�2�w��L� O&`#6��w�{ �ng��
�o|�B�^�D��k�.@���E��)�D�MB�����3$;V��˗�Z���9�w��m�6	��PpI�X7�za����mb�P�M�Ͻl���4�'���[�7��(� sP�9�1�:БvV�b��g4oUaf�UI�Y��`�k�S��z��xmkq��~��Y��	���/W��B�{`Y��?Ә)�B��	�}zܬ�u��pa�@\KiՖoj^���T�M�4�v-�l�׍���d 2\[��,���0�j����LXW�������V���V9��[`2�h��u5��"��l��,Y{��;����	M����7�סi��O�}F��[w:!5Q8Pw�e�J�{�m`��gu�:¶��\������u�W�U��;Vf[=��4�ՄnK]M��>sc�?{�g���s�1��KF��k������8r%�,�X<��~y�ۭ�?K��{�����3 ������(�u��\8�@�Rۧ�oE�TF9�,^p|nǭO,�4�j�����zh%�>c%a���ųdBw4�s�b�p��S�6�m�]X�jò�g܎�X��'bo����0��,�4sצ#���.��m/��W8|MО������G񸼶17vz+��;"oCS#sU l��\Om1���O<�J��h�y����1e������*��;����Sr][=@I�Iv �0`/�C�*]c��G�_��׆��2�әS6������y�r��t?(�l�wZ*��|�]U���,���FBd�n~(aj�������I�7�T�ܚrE��M�H�
/�ь��t���T�L�!,Ń�=�7)Q(]D��[��9��S�gG=�E6#%��RA��^�CtfL���W�z��8k����l�T/���Y[��ـ�Ͱ�r1/Lңxe���}��s���hp��R �ܬx'u�K`k��N�'�FWW �;zFf�YK�䓫�(�p.b�¸��k\��q_Fk�𒺵ZGm���5j�b�}���O	�a��֜���6�B�i�Jq�Gge�]w9A|�t՚�]g.�����)��!��ٰmr{����f�$�|䗮��qou_�yR�U�~Gh���a���!��l2���*��w�t�˰��[h�ܓۖ���3��9���Y2����t4�|T����'�����ה�B/R����5�TLD��܎S��N��FjE7gK��e���:����ʇ�8.-֊ꧧ0it ���@άY���_I�VF�Gh���eeuQz�BovT���.ۧ�:�.����������%��5�m�/���ӏ�Ƨ�ͻ·(�u���l{�O�j�6��+4Sp�"�}U�+p��ɉh��G妢�ep���1�=1r1���2��S����Q��&�@��|̦�g|]6�����vP�K^{p7ͷs�4�̠�;�&s�q8�K�~��;Ϭ�.�g�_8�X��}Df�?nNlv��W{*u�E���n#F� �����g��$�cT����g�~���"/�(�da��A��Q����m�E���]�G&dhF3@<em"8�k�J�]�4I��ݱ�Y��:ɪel�:{�gC�Ym�M�c�G>St][�?-�t����X�2?O_ᡈ�ִ@�WB�c[2�9����,%a���WNBk@��V*�U�x�z���"1����!���іhn.w5v-�J�p�3����5��du��Y��%ur�_-Fk�y�{X��?uvos]XD�x[��x3���Ǌ����ts��Y�YW�{�U`��HJ���5��YWN]�v�]΢%�Ɩe���<v~�����z����[:�2�S����ޓjV��+h��+�B$׆��ա[�9�SU-��6t������Yv�:޺NB�-���1q����7��zi[HZ�j�겏�����{(ު�a���GV|U���P�9�&����pʙ*�!+ט�^)yXhs��þg�։�(KV�j�þ�:� )��%��+�)�DvZ�a����*���=U)'a�+3��M���1яD����1�F�o�����E_[FB.�k��	'V��u�\8N�V"q��>�X��u�b]�|V�^���SR3�jvw`e']ۍs���P������Ra�(�����\�����նG6o�vo��2��²�_PH���v�1���i��2�es˲��\S���ki(:�\
�U�zI��s*��x:����Y��f�����Yn��`������ԫKu,��h"���#F��
��r��\�<�͏�o`�����v����9��ܨ~gR
�b�+"Py|h�
+�؝�B��;�=�u�pT@�b�$+�NZ�.���#K5��Z�M���c�\������pt�4]������d�B:uɛ.-tz�w}��櫦���9�V��i��S60ٸK�k���ѐi�au�(�0��U����٧m\n���;L�'ns�u��ɭ��]o����+�2�ky�1�8.�!n�\aӗ5^�z��Ӹ�Uq�[�K=����ک\-<2�Z���\�À>�9q4��`�˹^�Ԧ(厛�,w]��t.L]�-}ө�k^TW:%�<R'�E(�s;M���+mRt�Zǻ�,���ˑx�n<t:�4a�oR%�HEqAX���{+����B�h闠
��\c۫��Un��;k��»�>��x�X��͘9�jq�nelḉ΄Z%���|1J���a������Z�!]+u��v�<��K�lE�6X�Ձ�����Ѫ��ڈ��p��3/��UƐ�ڜȮF��I4�,�`��f�7�Z;�ԭ��Gv�/F�E�L!�`vZ���d!6���t[ܬ�뾒�A�W+N�� /o�q{`Ɔ���3�E#�C�>WN[�]a�Z��yHJPsP�)խ|K�qNR��M^;WԹ*`��r�rL�{(�%ǆ�[�:�Jj�o$0�vs�b�ZZ�dT��2�OL��릵;�-���ZE.�D�ж��mjFZ�J�$ZN} J|-����A"��u�����j�:��>?!lޗ�F8�:Ә�	e�h�"�,��3Zԉ����ʈ�+�]E�%E��(�eXR�)2*��F�eIm�2�\Tɩ!T���BD� ̹WUt�Da��B���6�Q�eD��JH�b҂�)�Y�r�E6E�YBp�Z,�9UU�.�&*���EBaS"QV�$V*˄AQ�F�4�R�EJ�ȫ6&� A�(�Q�EUs�L�(�H��C��L�Ԥ1(��IUJ�*)5�i!e4��UW9PTQ6�� �4ː�B ��R��*�D�*�J�H�""��&jAP����Es�1Zr.ET\�L���DTTDkB�!��tR9��ӈDr�Z���J*�J��0�J����d*m"IX�re
RU��eK �+X�mh�t��TT�U]M
��P(�ԨK@�.TUrH�!�!$	$���䋮�U|zc�OWt�]7��3-��2�Φ���j�z.��a*��sJ�ռWv�̾ή�	�״�[!��4{\�L�m���_LA�׵u1R�x�ԫ�^�?�8:Z��-������m��t^Y�3��F�&7~�TV���ϫ�������K�{���=�[Ԉ��|^��a�ْ(�z~���s9����~��|n)�"u�K��I�+J������;�'�0��O�{��A�]�r�/4��9��0�M=J�)���������슐�v[,�b7�``�IXϝЫj'U�2��� ���-�˺qޚ:��)DtAg���!l�iFL,��e�Ku�s��M�/pCgw�˺K��?O;�u���yS)ı�Q���S�VF�Kb����{���m��y�Z2E3v��M�e7_��T�Y��L���zЙ{��ȁ>0��~}�*˲�}��w:��{k���-��o����kْ�Si��V�Uַ�zEvBg��]YB)����g�&�J��X��0/p����i���^4�@�m�Oۓ6���Ok[��dW<u.hu��ONّ��U&]�?r[����ߝU�b�kT��a*q�[a����5�8zh�Q�.�f~ܵ�6Yf��X��de<���M0��D���YА�0΅t�g���{������c�hm3 ��i��p@��O�݂Y�J��	wWf���W��
z�_}��Ժ�,g1/5[�{mԮ�*�UY�y�?9��Ν��d�2�{�v���Qq�L�4�n9%�!����BX��YS4��
�)�ؙ|�]u6���܅�����:��t.��[Q�e�K��^��.���z!Xq��L��B���;[pf�3N:$s�g([lG3�����B���-�57Q�ݿr�OM�2�z� ��� 5ý�h��[Ֆ��j��y�3�'�i��[]/
+M:����*�_��k���Tݶ�l�U��^�2N���h�;=8"G3W@)�
4�w/�Lt�S���nh�W>���t��ΗCo� ���V����6�ukI��h75��p����ɽ��R#�ӽ2hCV3ABO�lGc`���Ȯ��T�������n�p�L�w��bL���`r��M˲��fzW]���Ò��9����ߪ8�>]:��@{֞�O��b���)��^
��P+%�7#QKEW,���%�������0�qK��޽5�)�@	��`ܵ;���؃sR,l��$p~�r�y��F>[h��"!�X�]"�G8[��:�M��(��i1c��o���~�g1��=*e�B�&�ж�Jv]v^p���N�53DwgW�&��Ʌ"�ډp�e`�g���䀽��������uX]W�m����.'f�!B�u��4�\�ef��]K�9���nlӢ�Ozj�w:3[�fv�}��~���)U��5�k��,G�	;���n�U!�]"Af�gތ+ً׍c+�-lSr��d(��|߭et7�����2�o��i���S�n���UK��U���Ũ6�b5�2z,������-��x ����O:���jzsx�-I�|~�ٵľ]��M����W�}Q����ٔGoC��ɧS�k�i���=�B'�-�
a�,�nx�p-ݺZ �9l��M�^�Gj��&y�)��ُO9��3��Ш�9���cC�6:½I�vػ�l����O=��&8�E�Bg��ƛ��A���Q�\���U�S`���]XK��O}9[�8r���/���%K��D's^���S+�8�n��j�6��(N�s#�oTkd�y#�CY��@�M�g�=LGM���W�����us��lMҟ-�Mj�c:�1=df��6;4W{*K��Cj70���5�.6��$V�O<��t���}Ѣ�mNi7Y�}s��b>k,�I{O�g�W�7<]�jS�%�/�C��]��IȄ���#U�����?W~�����w��C���9D���<⚵��q��7�5�آa��|..��i��ñ���)����R�T�ܭ=��e�X�k��]��n8.P#�K�����P-噡D���3�vb!�ĸ^��Xʚ��fP�Ÿ� 'dଢ଼�;j�4X�mi��h��lz�m�:]֊k�!�Us��� ��cw�q�t�t�����ۨ�.nl�q��M�ɧ�.Wh�Gu-���tc.���}�)����o(�V�n96��3��5�����+��3��qL�p/e�"�ƾ��Hn{I�v�.�a��rݗL~M~��J��h�B�괎�y�;��B��%�F��b#�Sb5�Q�t�ø��"��mr������\�-l��D�
��1�A����n%{��J`~g���{�[�c�b�$���>'>�]&C��
���Qx�/�X-����O"����f�Yzh���m�s|�{���jE2Ηu4���GZ/t��P�� �[���r�e�������i)��_�1��s�puݞ��Y�lWU~[���)�*S���zf#�"�9�fVf�
�Wm��ܯ
��y�}��M7%�jV���ap�nQ���)��lW4���4mw՚>�g��k�i���h������FFTG:���U1r1�I�-��y��m�jeu��@�KP���
U�X�n@� �s1�.⛼3��]�u)�SV�Y�Ȝ��i�ǎn�cfh�,�15&�7+]��G���|�N��Wp���.���xe�[��+��ܔ�������U�E�����h�Z\���Ȗe�C����q�Mѝݓ�Yy��̧zq��<�?��E��������ڼ���uf�BT���)�l�.�R�j2�v��7�����Ok��H�����K�aɍK仨(ԅ!���m9%�-39E�Ig۾ہW��v�/����>p]щ��y��U���B�/L�L>�F�4K@<e]� ��;�]a���]T�����[gC�Y~Φ�1ң�
����RN\iIjiX:e�/���{-�?�.�!�7SSJSOڕv�fއ�[gC��|i��tM�쳛<���������5�:�@���\k�9��\rP^��J�s�%�z��ߊޤFoC��z���tԠ�ى��Z�0޺�A���;������@1vD'5���{��I��N��\*=LUKfD�={�+��;�U�S=]M̄$�gF|�4A���G^�,��h��)��lK�i�rz��߯t�=��[�[�+˺qޚ:��PqDH��-�c��~��ɍlI&څ�n�����x��s�r�H��%��5�+˺K��g��wηSn��e8��.���E(z��Dm�ۚ�n�S���f�3�X"R�p����GpJ�уz�����e �W+���)ڔ�v�)�n�!�m)d����.�e�G=ż�o�\r��̨ݵ��&��q��c�����n���z��.2.��9�w�I��҃�S�
�8N��Gt��4Ƒ���[Oe7w)�� �)wK��x��q���&"��Yu}��o���J�6������=3Od��fJ�Zk)��]TC_��OH�����W�\���+�F�E---����#���;.1,cvY�mʬ~r���o���p�ձ��ь=v'�ܿV�0��;t�C�x��Uw�B3*����^6N�����$}�9|+k��&Mk����)�M9"�䗦˹���2�C+8�(���Z������ɔo{tǍwz+d?�]�1����\���r\�\����D+�3�T���=u͓&t����_9�F��L���b9�V���\;q�黁��4۶ܲ����<�ݡw>N��e�N\���%�����}�(m90⽎$�JS��.��~��m��7kD�z��UOZ��;��l��b��6Dx�!<�zTZ�4�M���^�y�S�OX�`���OD7I�W6�[c��7[�$5�.)�Ew$Oɾ�u">�N��q�#��o~�oVC��g
9��볺˼0�i�t����tꇬ�7D@ѝ���(N�gv�ݣ��g*��$��|ﷸ�a����ɶ'0Q�_D����W��ݤ���E���
�o��d�[�ޤ!fWTY��Z�ֲ�m\빯s�v���靺������b��{z_�AqcWWSu���ϧ2g�`����Yۍqɶ�3��x�쩾j�޽�M���W<F����e_�̌��I৒>O�܀(����UT�.tm��^��	dE3b"[k�u$�h�	�d�]Վ���\"�@��%�;�')����v�e��I���y�L-�m�
�"%��Q��L�8���t_��m��c��a��4Y����~�����3��7��4�M�V�=�}�j�1��$*eQ�OV��s{�U�Q�Y�����u�X�g��=�Z���_Z�����V~�ˬc�����l����3n�s1]��񧩡�a�q����}=9���B���&٠�=]�/�s)C�������.���?	�s9dK�{��K�ufK,�k.��!���"b(��}ȼ�~Z`9���[�k�����g���nU-Mۗ�J��]ls�x�9ٔ��9:f�xֲl���a>���
f�y���x�u�@��l�9l˕17�U�C{��
���x�7��S��l'Ԙf�:���Ww8=ua#��msś��3T,E��|���*�%�֎W�|��r�zo���T�y�9⺙U`����L��|EM�l������;���8x����s�7G\��	 ���"�t��S�p��/�L8r%��m~g��1���b^�J}0PN*����4k	�ӯ�{�6�w�kjÓ)�p�0��.#Bx�ͥ.������us��7�ٕ��9WWNñ�6	��%�mD�^F�����,{�es��.�6G�?i{�?-���qݎ��N������9��ft;�+�?j��狿����IqA�~��o�v���M:�S32e�c�����|�uM+ƻi�%=cOC�Ηu���{�e�\�l�,>P��b}5��q�-�,+����s:���Y����3O�\��u4wQ"�tg�C�ھ���SHOF�	U���뫱Ѭ���c;�@w�~����dB"���sp��~{Iaю���[��m�|�����֡�
��" ͱ�i�$<@���1�V��l�C�i4�;�/�9��`v֑�=s�m�P�,���-l���Мt/��3��`�:FHG"i��~������4a�sg���V�>�^�T�7r������Ω��t�9�q�S�`�2��08cs����4�Y�A�=W������еߢ�
W��٣�P۵^��#��۩�Y1x{@���*�,���l�³��zR��?$�:(���0^_��ɺ7�����T9Al�]�^�q'��b�G��޺�ۮ���7\<����j�;��|�)��v�9�}/��Q9�ك�Wes�(��t������:��D��6�T8�g�Z2������Sӵ�K��ޕ;�$n��I��^ܬ�Et΂��ߤvL'���t�G\E�qQG�X�^�tUe��q��S��o�7<�f���.۔i�����+�7��h��H�3�6��e�ZA�*����G�/DX�p�d`��ϑ���#���]�N�/��=����=��95���4��D����ư�ʨ��g�\���4&�qP
\��_�)d�����b"iT<s"�F�8~��%i�uOp7�%�E�d��91��pІV'�#e�4��<l�]N��cϮsu��gs��y�L�u��!�b����s�ǦK��t^�ɇڨ���xl�'�;�U��;Zg�82�tS*��1)�G�:{�C�Y~Φ�1ң�
����� �y����s��RxU�;��S�3��	ݭCm��.��ڙ� ����%]��z��y��m�X�kj��S��5y�vo���
������#����9(/~7R�[4�Ix�����ⷩ5�%���ur�m�b�z�7�v*���t�8�WpΎ��r�����ݨ�^S���ܽ�&�<�sN�`��&6��M-;�j-��&�a�tn�x�7EΑc��������2y�%��Z��Q _+�ݽ�B���'�eNn����.c�p�*��Fi���}g��SuUpeop���L�w�g	lw<b����u/6�h�z��ww�u�n�j���d�?xT_q��t
��a�����8g�vte�@h�Ӳ+����ޗK�#��h���Si>᩾j��n�>�wr��úH~~�t2�/��ҞK�N���2��0��/ƻ��{�\�ۙ�#�^��e��B[R3��t�~~�w|�QN�̦S�1J#^���W�Գ�QTK�?Zs��E�7��sS�H���V��n��UR)dE2�}�QVxt���Zy������֫Y�tT@��(�p_X�u�0pcץd��fJ�M���%�:�o4��"磮V o\n�cЩX�x��U���d:�X���g����t&>ņ���R�vY�rf���8
͝i����×�S����.T_�b^2��ѡ�s��Wxaf ��Z���N����7m0�|{��;�s�k���-J~f鞭pz;z
�4��^��a�c�̡�H�,���G\��;շ[X{��壘Ln�o��YF���]�1��[Q�\����^����ڨ�����9�ô巶U��MT��߿v��,��a�]w�7�pgj[Ǯ%ƶ��<��<�����ܳ�<4{�	��R,d��]׎��!L"ʜ��E�PuW[�ͣ�k�N�t1*Gt:JS�;)�U�ݱP���o-��&b�����W��F��"�Jy���K2�ۨ��l$��*6�l+��Uj��ku�R���;c�[�1���o$Tn[o2�/hfv�;���J��*z�F�S��6��
���!L��{n=fa���{4N�O�kXB�]�^�ە()�l1�V��P�G�Q��*�ޤ&,<��\�]�8Q�X�=���i���N�L�����l����G-��Մ,�W �s�.O��w�R����'��eX5�,�巗G>�w�:ة�@Z}��f)6�@��a��e���:�Hv(6��d'}��ՠ��3������75�Rl�45���t,�Z�a��'L�B�g[[8��b2�~�4�-<�R�tfe�e�<�f�	�����$f���M!M��C�i&i�8�Y۩���jQ��,�z�sQ�kڲu5:�d{֞��<���=v#��2��{��*��q��;��k�^[2Ӆ���y��KUy�+���ܩ.Ф#D�&����f�U��t����%6��D��Ⳳl9��ou�	��W�j�[��f�;]�'v�C8@���l˩6�<'Ǯ�g�p���Q�W�n㴘���D��p+��3M�k��&��(p�5���b :\�]��V���ņ�抐�[���o-�7x,�y��b*t���:�U�%^�Z;l]r:�����elͧ]����?�JKy|A`l�������������g{�|L��yt$쉄۬ٺ:�����+�m�-�7a:Wf�F��5Y@�YJeٵ��.!����N���i�B6u����6�f۝��oBn����ВEԏ:��IyJ�����##\E��
X픓���y�/`��}z�R�L��n0�ll��ae�Wj��đ��&pHQ���4 �_U���v�]j�&��oaE�܏�vQ�/X���v�N.f[UqY"��ڄy�^U�[0Z��<c�#n�q�6�鵵\��P$��Fu�rv]�C�ol�T�7ݤ�9�EN���}�e�g�V��v_B���Tǎ;���Y�]��Ru	ܹ�W}HvG����[� o��)A��i�0� .x#�T���\�;ݹ�қ��r{\��8,'Ee�)�[|0f�$����2�2�T�ef�<)f,�/^֞���n$; ��]�Y��Z�c8�G2�f����л��ewWk��x��VV�0�F�:[3	���9���s�R5ח�{:�Rr���X�iu;����q�*�".2�rU[t����i���	W^�w:�^I͇T�WS�OL�`'�nrQ�JIȅ�=�5��v^�1,��c�Ls}a`κ�ӏ%�GH�XR)��f�Ⴔ�-w ��s��
�����\���VY�Nl��,���Ȋ+�%s0ì���-I�sr���U�dT��QV�Vh�F�*�pKGuΊV,�(Ȋ��y\㆔uP�����L�*�wO֊T��n�I�S���)�D�	���\��8UgK2�:QYem�I%)imde�E%�*�̫������i��r����nc�QX�QR���ZV�Q���Ӧb��L��ȇ�R���I�wMQT�甐�y�n����n�^�P��<*��2��s���Y+H�)���V�T�n�������%��W�����,�V�p��e���s�Qd�W$�M�̑D�w	�4�6TwG<�R�Gs
��\�)U\����"*E���35dPU�Q���VP��p�9z��翽��?=y�3c jv�܏%�wosF�2�+tm�6;y���i��vM]��q�Y����)G���Z��Jx�d;�d}�[i�&P�m��t��b9�V��T.��M����n�,���0�j�b���U�&�'b{ c�5t �'RF��LG�e���q'�brʡnKG�Gp=M��g�]�n���eWeD�j�X;��)�`8�������K��OJ�V��i�us�����}���M}p��CGk�a�#k�Sv�S|��pO��!;Â@y	�u-��T�V&�DTf5�mÑ�w������y��qm_��b��}C� �/�$�P0������9���n�l����њ�N
��,H�\i�w.B��7N��M}�'���
y#���=�\���	�	��/����չ���}6�eḋZ!�1]I��?\[�]Վ���)������@���R~��衰��M0�c嶈\+�LQ��^]@��+������F�P�����DԒZ����x�5�!�1�{hQ�%駠��0�a���q���N�6�oYӱ��o����th;���X��(K�K4�����	�Ƕ��i�2S��<����l6Ƹhb]_�鮶k]����:!���w�^�[K�9K_QSra(�u�#7��Q��Y�r�&�ܦ�Y+`�Í�R#w��-;���U�u	�u�ܱR��HsF*Y�0����o^v:�5�TC�gT �a�]e���t��C��bw�W6GF�QF�Qr�vf]Z�3̺9�6�������0���p�i�01���zNN�48i[�v�cv�&���:e>>\ܧ��s-�~^�u;˶i�TCն/���J�i�e��ҚlN��O���j果!�vcw
ܣ\��f{@�c��yF7*�����+��}AUM}9�e]N��h=�?cM�� �k�L�yKr����5l�SV3%�9A��=Q�s�$A;�=�1�5�(8p��]�tk�8%Q~c�+���ΟL��9���ras��a���͕�۷�Ո5aɍ�;�	�hO q�J]�!�RA����
*�VndgD_S���R_;��jn�/�~Q6CS#sW�he�2�"���$A�z�F4!��[qg[��k�}�f��k�M��h�c>�^׃���S��/��MHkR]*.]i�P������=;�w �\�#pj���
VKJ���[��y��U��^]U����Z�͑;
��7��م��;�Ts4�ې��xn�tE��M�H�
/�ы��mz��>L��0r���������>X���Vؽ�(�b]�,K�>th��A��=4S���?aTś2._e^���l�扡��24r�]Y���+�R�z�"���#���΋�u�͎IV{�P��ˆ�MTK.�x��ֹ�F�Y
Y����������ޜ��KS�\AX�����" �ҝpθ��hM��sp��l:���y��3�]�3t��+T����B�D ��d<z����㜬F��-�ۖ��*���7Q<ilS�[���T8_�E������uu4R�<C#Oa�=7�����_>S���v�l�ߧ�$��I��v�^����w�zc�x���|��.��!�T�4�AP^*�����Ol1ɨJe�3�Ų9�8����Z+J���5!gC������98���ʇp��T򉞭S{uN���i�ǉ��F���eBЈ�ah���elWUkz]�EvT����t�^�7}$a�܇�7��"7�5����>F?T���1�Z�l�\7$�qe1=����a��I]�9e�����[�dW4U}6���ЋG�����Y�1�4��ǡ&~/�yl�6����\���Ob�7�/U\���3�7�%�5�*�0@]�es�!=4�N
�ߎ��P�`]�v���V�չ\��9us��HouI}��p^��0.P�,�����Aశ���ɶ�&8��E���^�b��i�؄X䭠�4V��"���>�y�eUn�c_�B������FBRf1í%g�w2�zs|�Z�N�'B�v5۵��c<�J�g	��X���Sk�����������A��!�2�r
�s��A���_�#�4eܫ����W����b����~6�T_�m�]�ra��� ��S�R�.JY�zݣ�ɴ���6G3����=�����[gSw��<�jn��5����7�$�nh-N��W�_�'���w:�)��*�lmq���ܕv�m�~E�C���;����35���N��SVsdM���p���L�N�AqN9(.jap-=�^)�z���f��kw����۷G����*�r.{��k��L2���d���	���-���1e�s��vRQ�s-�� �Z���S������t�5��������Ό��@h�Ӳ5��,ξh̡2)�܍%-\D�4͜n^��T��wI����K�qޣ�����C�.T߭K͎�����$���nD:"�7i��HKm$k�R���y��E;���oR�.��I�'V^�MD[��1n�<�� ����Oe7_r��^Y�����:2�p��N���2$�i-
�,]D0��	���-��0pc�J��̕���S+d����7=s��
#D]����(+H�Y��K��#����|<i��*u�Ӽ�FP����ڲ��U�v�e��zRBs����0u�a���L6�VuZ��z^���SyS&��Y��u#6��,I[���G�=�j������=n�N�ˎ�7�Ws6k����d���^��"�6� ��24ϓ��c�c�Q�f��~��֏Fs�l)�gfE���{~�(�_oK����+��n�,S6K2���A��	��V�F�[P����	���.����\��g�\�ރ�%�Bۍ~˹��8���V-��D�]q0���jt��i�����`�wyk(�zf3һ�cuKj0�F���^�\�Mmw�ʡ�ٛ0vp�$>�Eؖa
[�L��P��؎gT�:x
f*�����f2���S)û��^M����ͥy:_�F@/: :/���b8�l�xQ���Bq���8���g~=ҡY�$�s٢�rX�3tM�H�z�[!C&_rf��Oک�\Xv�J������\��u�6b-S����)����eʛ�������d�ܑ��7ћ����H*'L�/'>cMX��ݲ�㻦�|{'�;��0�_Iq���������ϧ<!�>��(�;��ựy������͔�w�Iᖎ�ƚ+��l��s�n.�}��C�OU'�^H�C�h?�yL�Ld�o�"��J5���i�b�Oڶ�wt�13;1?���C��5��	�v��Dz�靎*�aɔ���Qc}�o`4�i���'iDxҘ�f����^�Q���f9���t�w]m޹غ봥H%+��IZ��J7x#���_j�[�n�g��~$8�-�qL�+/�8���b����z;�0�qL˺�ަ\@�G�d�Y֋6u�U� �0�w��x��^`-��!p�lDKmy�5�+̺8��v�쉊����j|� S\S����B���c���Q�%�z	��+E{OL?D����;wz*W+ا�����BE7ts>����6>�	qinx���Z	�M�k�R2���hӭ�H�ۦ�=��j���uT�,�u1L�9�6�[K�o\Él�e����`c��u�oZ&-����o���2���s��}zܬ�{f*g���/�k�i��~��붅���r_��ޤzs�N񇦽���=��R�^��E	��`�0�W�(�:���7ǧ��nU-Mۗ�1;m�j�n���a1�:l�X����SM�� E5�&yk<����%p�3����А��&mhi��'�k�:�T��/���c�]��g�m^d�S#�%K��D's^���jޒ�u�Y�&M�m<mOѣ��a�t�ߏ�{�j���MC�%�z��=zb8��R<}�v~=��rw����csToK&���R�嵧1\�����M]i1\;DH�Ց��8�yk�B�b��d�%nqz�roM�����^����Jl&8�Q�*%�N��h{��ޛCVǐ=�69�.�
7fuu����RU�5�֟gh��]�.�d�7��5��y�m'L��ҟ-t���Ehd̎L!T4��p�S��������Q֪�E,��_����y�W�N��wV=�4w�Ηu�˩?hQP]z����Znp�P̮�_Qh:r�����l�ԈDq���7ʖ�MBU�-�C�·u���������J/O]*����t����bZ��P�L�	[�N���ZwQ"�(�Fyt>�͚D��ʋ���c0p5R�l:�i	���,Aߩ�)��z���d�� ѫ8�^�c�؞��P�I��uك�����eOUp��(������>�p�KߥF��"9�y�~��o72�Y����W��׻E��w,tZ[����OKFy��!��x�0�zDJ���){�}�Rۉ��}��U��fe����;�T��-����Wg��V2���;�����_��}����m#Hɼ�X7Oes�r��L���M.�w���D��oeC�6�C�}ӡ<^f�5�+���p���`���ah�ܬ�VWUl��ߤWeJy���{�����ŋr]�w�!��d�`�}�<�Ce���c4��h!]�ͮ���ܤ�G6�"C�,[��s2u�{ WKz��u�+��}� �LuziWm�H۽̍ɷsW������+�ر,\�xpN�u:��TqpAX����c�����3�x�{]]�+��G:�O�2c�l3���;��a�EюpD��sO���ny�J�4^l.۔i������n��آ��.��v�5���E�h�n��Ep�"��#)�9�l�=1r1鄙��2��M���c�c�_\_Dm&��J��g�b��u��]�`�!�B\��O#�Y!�O+o��3����͢K���.�����=��uI}�mݒ^��Ɗ� ���-���M;�vZ����sd(��T�ߖ�C��;�=6(]Ѹ�s�ǦK��t^����졄tq3���֝Π�h�Dm��l��n%T��t�l�~/:���J�|<L�&껑id��ޝ�a]/|�(k�7=]៌��������`�&%�9*������q�2���D��b7\�/��2�����!,�;�p���㒂�n�p��/9�[7n�Pgz�bn�����O͋z���ak��2�-��$�w�,!ߡ�%��<b�2�غe���h��/�jmS�6n�9{��I�u�'�eӺ_u0�=-�%�vtXh~f�-ն3e��@����+Fq	�S�y�-Af9v^~�~�"�]3V��hy�]E���9�y���V�r�uS�h�	��!�e=�n\�������+ΜNK4��H���_�k��͸h��m�	*g\�̽��+ghr��krs���9N����h����p�J���>�1\�=��t�9�S�t[�ԿO�Jy/�GNX�L��j�U�ua��l�y�;���4ɑR�Ne1�L��L���L˺K��g��wζu6�d>%WY=SG퍺��7�F�3�`H9��y��ǚi��$S����Su�3<)dGws�ѷ`-��7qֶ�ݑY��\�2�Lc� I��bX\'�~�~����d��fJ�M���\�1�ՠ��\R�[6��Cs�T����M�M��E�f��{�E�1��vz�:���`�ߎی��F�P�׵X��t�[����!���+����X��_2�!�ax��-{;:&����h�;:�-��;��Z5�~e3ծ,���Xܦ��|rK�]�=ю0��̓��������Z�8w�$>d6EDX��l��l�A��J�-����[�Q~�4*���-��>/�=�����֍���IhTqVȗ3����f�0z}i�J��sYn�6%%�~y5�U��)�%��W��T�u�_k`��x�u q��m)xQM��X|�im ~y�O�:�1ͺF�(�J��
e�ܦ���'1�s����S�:��$o�7����]G��uښ;uٴX�+����Pd�u8I�	����N��r��bj�f��CE���&�,>�sB������]�`��J�d�X�r����v�tE�fp�̱�4w��@ߛ�Svډ�+̏Y^/IA�@���>���#����#5���E��`,l;��+��z��}{m��O��.���M�aM�n��K!�)�rD�,�>K�FM�\������*;.��kҺ����Ƕ=��ޗ��}%�
e���l��wg�S�V'ޮ��ಌK3��_M�@v�Kq��4W���wUF.�}��=�OU'��,�\�v��'a���Q&��IߜiZ-e��-�t��E����8�`e���V���6�48�����s5�H �0>1C`<B�K�4�я��p8���(�H�����T�e���Qy�oۀP�@�~�w��@<���!�S9�y��^�z	��+@*�=\V=���q������J�zkrfCwr�+�9�zБcWԡ+�Z-�}hH��Xn�^Yum��P��ŷ%ξ���b{6y��z���.���Y��b�G;���iy޹��e����j�kx~��c�t��L�
ꃣ�\���Y\��L�����_�����\"Bg�Wc��^�S=�%2��ާ:��L�i9k��-�J�Wj�doq�|T\N���X��r#��g��g���GF=7����y&��w̠"��Y\O:��L�۽����5������i���=&�[wF
w�N��:�f�[t�z�|�]1�������f�h�7����E�[K���N��X��ǈD�o�bX�ݩ9ܝ��(��̲�,N��0�	�L����̣�6�n�ً�2�%j�̡�R�c�"s��9���Y/E\a'ٯ��O�-D_;s6���.����r.��b�p=�b��x�k�rk������ܡ��ܥke)BcأQ.�p��m���|�;	f���hG�ld<ɝ���:=��};zg���\2mZ��=}��]X�e\�V�w�qS��TY�����@嫹�k��U�Me�ft᯻�����'+�ɔ�5vҧ���}�`�
�p�.^V�^�|Ơe۩�&
ۏd���Z[	�[�Ĥ�thqUf�]u��~�32�ä�M���������L�vՙ }A-twx��A���u&&o9
�om�C���$_<r$!�XNVm�6$�m�,���{DD�!�o.*s���ٝ2�.V2��]}��3PD���h������۲�����O&� "�fL�΍��mZ�JY����dZ5e�f�2]��U��!���W�6@���%��5؅�w����zT*t[@)�>��B��ݢ�\���!3Br�W���KQ�C�v���DzN��'UzΦ� S��rj�pi�л��z�,yh�j����ޮ�-nd�6�I�6k�����[�z�HL����s�J�9O��kv�ړN^����a��S�c�t�9�
sjbVc8*�Y��
Z���]�*P�\�}��Q��1Lp.�ڣ��K��!�v�d7j��-�w�e��X��)0��-��秈��}���m�V�Gok��Zl�D�yx�]yQP����9�K�V��oa����V�ˎN�����C	+pr
�6���l�5р8<�n�-���P�>�u���:�uu�(d�U�2R�H�Yd#����R�`Q�cv[�T��e4����B�#��8M��:�2M�Õ��l3�-�b���_v��v�&�bKY�t��ݺ�JS��-(�k��{Jv]�\�r��2�:[����Ⱦ/śu Pι[A��2mIW�dsR}}�U�Hc n���peh��j�;��w����X��ez7>N��*Ig;I�.��S�}�x�X��"}4-t��~�ۏY�1^nk�Fr��)��6ul��
��LM�$f��Ӛ�;x�[�%�H2��HY�N��j�i���x�6f�m�b@�� ��T����o���R$ �(��T8�q�CCy������wM;fm�hI��/r�k��x"U0%ʖ,�w���\zsm��(Sw]�Ճz���"�[Z��n�{:A�A�(�ci/�MQ�x'߮�5T��K[�t3uۉ;��d�uNDG�z稙�����B̢��y�BYQ�t�B(N���U�J����hR%%DI����իwr]�LR�,���9-\�r��y�EW�3'R2��w7\����e���!E�S��=n�9jsE� ��i�h�N��Q��	bG�y'�Ј��^��DFNyG��{�J�Ԉ�JQws�ȒI<�qԊ"�h�Z�(*�.��ʪ�LS]�t<��I�K����,����Ng/wr�4Ē��!�L�ۮnf�z�������QN̈�D��tOQ�Z�RN�$�v�j\L��]��������(����0��J�t'K�b@M"DΉ���+���<E�2����k�X�X��ۉf[� �;c�c��/���ȋۋ�+��{VXt.���OQ	� i��K]�����~�V�M�L�a`/.�g�����O9��2�Y�Y/QZ�D杉ŏͷ���慰��U73�����dBg��ƛ��ĮK[�c�6�)�aى~�8����E^��3z;�F=��+�x[	h��_��(�1���^�<@�z]��+KC��Gq�ȥ���[)���!���n�.�A��rcEP�	����hOM1A<�؍.X;tL��$V!��g>���{W8|MО���۪K�߂�!��B�hg�p���m�;��꼛=�'昃��UIy�ej��^��ǿg4w��wZ�S��3�46`�6��cV�n�������m�i�񺦎�Ki��*�����o���U���F��[�9o����M���;/\��ŀe��z&;å,��	[�N���Z������)ا��k�tjr7M�f���_Y���5�i�C��pGWH�'��nt� ���w�*�K���P����C��̮���f3��s06���aј2�3� &`:4ϲ 1/R�xft��y�F^QPB�Y3� X��	���e�*�.�6�� �[Wۃ�SYm�m�'���V8X�`n�P���#b���\_c
��6,X�w˦�2ԫ�4���
8����g����.�=O�ʺ<�uӴ�ͭVJ綠8�U����X���#�����W�o��r����?�=��C��/���>�d#��Ǎ���Zm�@��A�uu�y �ng��{���gI~�J����K�S�sp�{�R��ze���l��
�dP��C8�����kĎ`�Xf�XƐxd��2�M����ԅ��J��}l�K�+lॴ�~ݣ�U���N���e��q�
���_���3���ݞ��YL��oK�H��%�K^�͌��O"�mH�/7͛�O^C�"�s�7���>F:���|�R�۰�nI�궜�l�v���]D6�h�7���w՚)�Z`��Ȏ��#W�.F=0�?���-�U;�o='̾�Ygk�߫s����2��q�9Ĝ��՜�{.�1P�Y��;��!=N_1g���n��壄��ǎw�YT\=���3�{���/�/��%�Lh��	ۮ��h*r�C�U�=�s������&P���t��&_�^�X�wF�\�����p��ľg�ܫʜ�Ӽvb�>w���K@HK2�R#��ڄ�SbUL��t�l�~/:���Z�]Y�_�[����G#<�-�.G��=Lu{g�'T�����F��,XS�Ӡ.��[i�0�Fm��Ή�˽m�w�S�x�������UM�I��ν�S��mv�������[�i��v+J�� 	�(�T���ҵ:��-+P�rv�NA��cu�S�w5�f����Q��X ~߽��]�e���56��RL��rU�/4g1h�U]��4�p���s��9�C��|i���}��)�"w�d�����㣮�p[�R<�4Ђ�c,�W}/<�9E����h�c9���e7UR��� Y���w�p��t#�1&{D�T�̍����#Q�ʊ�\ױu/mʓ�����3 -}��OWSEyK���UƉa)��=L��v��f�� 0�#����n^��T������-�˺q�t�44��DŮ+��F��:j#���P�g�T��&�i�HCf�F�E2�W���'>����x�Z�2�5�ɚ���}d�.g�tW�JM�]S��8����\�wr��5�Xvz�z4���E{�*-n[��;�v]���e����x�uF׆��X�)�ÂS�?��ƴ\�Q�D��R;6��5;�Ǜ�!���zE7d&x�]YC_�Em�g�di�q�Lvyʙ���E�n:	�� 0�v�V?=�S�������x����F��b�b�((���Lʙ`�oو~�vmN%n��/��ӂ�o�pYJ�	ܘ�bHv`��pYU�x��D�V]M�����*�S�b�Κ^��3u�43js2��.o䵼1�G7kXk�����	R����5�5l��J��I֊A��jc0�w:Yd�h�e��(Pj����zq�[a���͗ƹ�GN8�=<z(����$�6]�=�P��)D�N,�@ip�C�)n���&;�6�%;��F���]�:a��r�%��37<Rw̛�� �ǜ�|"�j�|���"6X����	�����u���iP�v�k���V�8���
��k�W9-�̻-=a���U� ��D�1]LG����qCI�����n}�����/��^ˠpw᩺�7jEk]j�V�+d(d�+�L��O��q�]��u��=�I�qԙ8��k�fm�溹����=�gK���ʛ����{���5�.�(d��������)L�Y=�{�0����U0��ҕ�Ä�m��d�=�/�o������������'�LkՑ=��;=S�,�΁@��".4�Q�l��s�n.�}��=���wT&'�\6�����9kC�'����opw~1>�2Ju�7�-vD�"���m+� �E���&�b�I��d4^�{�\w��c�t�!5�s #6ǡt��i��5��}��mi��x=4�<>�k[�Kr��ӫ���1�ѺG &��t�1�ژP���E�OI��F�T�?���b�#�훲��m;Xzn�8� �r��d���u%���:��}N���hҩj�a�,�\U�@oV����{]�V,ۙ}YI�9(�G�Lz�m~Z9�cP,t_��Sn��% �ơF��=Nf�Zo	z��k������{6���7uۂ�"{��Hj���$wg�OL�c�@Bg�p�k�a���+��^6�kwk�/�<_�z	�fI}��U��iuT�2ΗS�;�i�i}�q~��6���`��zk��;i�y�Pn�cGh�L�����*g��[��&��4�vdK�)���J�Y����7�qC�f0@�g�E�n�M�^ �xap��5΢#�=<�aAo#jYUC�^�<��B����2Ӫ�s��
��uSs:+�`�^D&{<e�_u�>tvV\$ѕU�s�m��]���i�Kn��z}��,��8rR^�Z:5���*_�P8��em�����w����y]%���Rl��n�����Ɗ��L!=ϜF��Ӵ_t�q��Z�H��+kV�a;���D�+l\��؛�>.�᫪K��Sd5#�SP���	�U�����ۿ�k�,���]�����d�a3�*ٕ��ez;��;�[gK��f]I�E�M�th"x���^���2�y2���X b�U��%jWKB�*>���BJ�����h��X͠u�����ط߃�����*s����U/;��[Rv[����a�B�˛I����i�7�VY�6v]]4{���Z۔��W\E��xJlZx�����o9�YܳsZ �ٮ)�y�6�ǁ2�R! ML�p�*[M5	W`<�bΗu�-X�y���+YD�O"�x>�fU'�z�w|0Zw�t��Y�#w�]eq���$����+���l��=W�;hb�C�ھ���4��q5#�:�}O�[�*�.7�2���#�R�k^2�vB������\��R	�tfL���T�Wz�I��>�x�xĸؽ��N�bi�P21��D�Эq���ơ��5Ν���â�	��񻫩����XD���(
k��=�.V�J�%#��rȜ1�،���7q����x�?G;�[�kw�]T�]=׽�ݓUy$�&��t�|�!�
r��[9��#�ɯ^S-�{+��ܦ�,�wRYus���2J�E�9���:P��?[�feC�� ˋu���E��������|L-�YL���##{آ`a�����I��r���Ƚ�ǜ�wm�׈눽��aq�i�#S4���xԭE���b-��
�=��v�r��F�5�dĭ}��x.3-[����HE#�F��y�1�+���	6��/��6o�3F�6���<�+�2�t���"ת�
��Y�*\��0�{�mL.���utҾ]�^跁�b��x��8�Aq/����t�!�y�}�ra[�ť�ƹ�˜�5]��LI�ٔ3�2_u`]c������zG�E�z�H�w)}��)�/�79�]l��3�m�SO�h��͗s�.�2�;^%EOzF2��/�Q�_��H������y�Zʢ�������=��T��ݒ^���ƃI�s�A:����Zj#"�쎅�3��!�ĈR�M&d��Rh�~ux;�=b��������>�'a���Y͞�]�%�7�:_�dÚj� h�X�,��GM�	��Ī�[h����+��:��Z��=��sf�v��}�����Q>yh$�K�!��z4��S퍮2�s��'�C	ռ.�:,��Vdو�Hsb���/:�k�L��W>qN�L�τ'xs�?%�N�Ψ���!�-��,weU����^k��E���DcoC�ھ�a��UH2��O�}2��2����eZ)OTfhq���1w�9�-�.^�Rw����˧t
��a��z��)�������_�q�e�p,b;t�;:�x�=��)�v��D�U��>�\�:f�@�~�t.��{�|����pF� ����ְ��Dsp�DW��x���!hɦݦ<)�!-��t����<�YOG6e��w�kgb4�a�'��Wp���Z�����V��k�'��ٻ����/*��WgN��n�ߌb�6{:�G�6W�q#�8_IOror��W	�b0;/u���u]y0P{��m������㴢Vn�ud�p��]|�x4_rJ���uݣ�ޫ���ޱ,b�F�y�B��S�-�y��\�;F��n�ǹc;jb^�+2;{EN�{��ٱ�	��.���e�:��� a�'�~�~�p[�zVO<��kU@m�Q�۫.�,u�e6�x�U����;g��Ք)�u��^��f{�F��q�OvxDNQR֤m��qx���v4�ݒ�^ܪ�粧��އބݱ/L�����Ōr�E���SF��*v�5�w����7W���&q�a�ws�ƹ�L�k����Sr�rE��I~�y�l��P�_tcj�A·<c@�p�B��Qq0L. �	N�-ec�w@M�-���V5p�N�v_�ۯ�����ٹ\��.�����6X���!3��#��6����V���M�j��.�T��ct��e�9�qc:2�Ԓ�~	iv&#�Ci�8�dW5K��l�;�;/��5��⯥�8-���n�MڄQ��B����a	ݟ�Nu�W`{���\Q�:u��ʩ2b����b��׽��O��.��.Tݶ��{��� ٩�79Ɗ��W�o�S�ę:YV�wl�f�G�4�s����Ԟ�����k��V1���{�u>��x�K4+�mbw�������S��w��Hi$Q}�-!�Gp�ٰ�p�lp0oni�O�=JV�ɖ� N�N�jǇ^��V�0n�xg0�P���u1N<�V>�e�_����ރS
�xu愺��\r�c9�����z[���&�{����e�M^��G{C��Yߺ4 �6^qq��f��e�����u��7_;�Ptft�#LUJE�p|�k���F ���İ���N��p�u��Db"[J�H:~:�a�v.��g\��?]���'Swuc�_������|��)GQߗt״����\+o����J���>B�z��e�j�s_z�h��@��t_�Φ�Є�7E���A������,IW��:�{�}�g���l�����j�1��$7ts>�����b �!��p�z�ct�8$�}*�f�����{i�8&��<v��U���U&�}%�PG����I��s7�DZ�q�n)�
�;'��g�e�3�9���v�$�>>\���Z9oK��u;��ۛ'�M�۰Z�
����e�����d�U����$:s�P�Xl0�SnQ�u����ݽݛOo�t���Q�F��ܛ�mU-^�Գ�?L�a�hy��j݀���,I��3������]yR�6Q���k����XU>x�N���"R�մ"ʼTyH0-ö�p��1�jҮ&�$C:�EZ�gX�H�$��o]�˝��w��uܕ�|u��
Ś^OEvþ��X�]N]Z���HZ9��v�R=-��qv5�fC�ɉNP���\���nU�c�Dc�1�2�!=��k�i���d��k���y�ݨ2L����lAwU�L�J	Ū���2ً��kۈ���8\'��n�yc4��Ʋt�{�'z0'�$)P�8��W8z�&�O��{��uI~�QD6��M3����<�qUQ��s�|!�)QӦ��}ʆ�K2�;wD;W�Vτw�Ηu��?`@�9Z3�D�2�w5�}&�5���'>
��:��m:�-��hJ���C�Up@z�bavN�f���;�vC�.����K�N�"ɢ܃%w-�7��X��P�g����ח5e���Z�;��m_uΘ�'<� Y�Aȇ~d�\_�.�JɁ�A�d��"��}�S}V9�vy�?VI#�F`˺�e4�Wt @�G����[�dt�~͓vZ_�i���J%�r3F_�T؍C�1F��߇q���E�t53�uu4S2�g�ե�n�)�펻}m�;|�)�Pi��� ����`��s0g_KIߋ�NW�E� 1���������0��1���co����0���c�m���1���`1�����6��6�����߃�m�0��ٌ1��L`1���1��@�co����`1���c�m���m��b��L�������� � ���fO� đ=���(��H�IH��*�
� ���)U$*(  �R�@TBPNب�J�IJ�D��**!R����V�)IJ���J��!*�"��D�J��R��;j���M��TRR��	$��)��v�P��Phj)�PzԠ�����*D��U�Of�"P���H�Q ����j�AT-���@�:e)@�T�����T(�@T$Ѡ��UR��   ]�y�>l�ø޶�׻4��k-���Z�Ӫ�֧F�-��Q֚��tP�T�`�S�4��j�@:.�6�P���(TJ'�  ;;�Hhi�5Q�k��A�5�  �nϯ�����=N�(
4h����{�  ��X   tPξ�tQE�U�����ݯT�B�k"��e����  ��Xj�7�]kTjtnۦ�Uۜ1T�53Q�j�>�=��s�A��t���r��M���J���TED�
��>  -8 U&��z2i�en�t5N�wݯ[�宝n�j�i�������ס��k{;�o\�nδ�h�͐�{�=�]�b�={n�N�P.�PPJ٥��+�  G)�}imO��{^��{����ΰ�z����浃�:S���z��K�훮�ۄ�ޔu��m]���v��ݯy׭V�6޶�����ۧ�^���ݸ�Җ��灶P����J��֙�   ܻ�����{^��k�{m���+�V��cW.���o^��/w��C��m���fn�هl�v�v�{��=��l�nu�A���V��ޚ=�u�v�1(P��R�h��
�$   ��}دv�����jr�kwGhv�s��;�n���W�vנ�gA{��ozzǰ��r�u{�q��Eݽ��e��.�ն6�4��o4��Rpf�^��
D��J�U(�N�.��   ��t����V�k۪vΗ��w�{�ikmYn(��^ݦ���W��{ow��y�n�z�ۮ�el�v��=ەv�kGt۽<=ۮێ�G�۹���j�1"HJ�U{jD]�QW�   �}�Ю����'�5;tTwwb���n�{:�{�9��{m:���S�Rv���G3�V]��z��wg����e{ݓ����m���{���Wm[v5WuZ�mn׻Z�FڥE�HI	|   }����j�{oFν�����5L�;M�q�K��qM�s�n޽���g����޻$�U6�������m�r���p���m[�ד��c״ӷ�T�"ڶ�������fU%T�F�"�ф��)� ��)�L�UM d��)� ��!�d �j���*2��&��M���FO�߳������-�w��/����߿5��k)�83���z�ߧ���o����ٯ���$����IL$�BC��$��BH@�rB���BC������:�^��+��.�4��ZH���o(�P��r��lIX��d��f���rJ){�e�Ș��+��N���ķ\���mdTVآr�H+F��q^Jߦf%�FT�鶖 .k;DoPLmZ����$FJ�[�k��j�VVhYR�ʺ�e2V�u��l���X�t�3�V�T�RJT�ݧ��\Z2Ef�,*CW{g7٫�b�mm�%R����W��s)���@�j�Q�q\��o�2kf����iK#��'e�,m���e[�
�%dM\�f��UMksN��X�S�(��I�T�vqJͷ,�C 
�VH/��H�c���e0S��l2Mٻ�Mk���{�3k �#�b����5�lUӕ����������5GoH�{�MKf���/VR�4�x^�PX��'v6�0�bwNķ��`���@����Teu�i�LФc�4��&۲N�Ba�x�w���&���M�R�Y��̀� ޵n�Ӣ��T��f�MB��ٗq�y�3��7��U��bz1Ԣ�N䣒\
P�����I��h�r�o
�z�#i�!Vl�tf�����V�Q�n��A�̬�+��#�I@u-�٪�]�������
ܩi��Y�VKm��m!WjQ�Z�ͱ�h�A r��1Ck�L^�oc��Z�{���*�Ȗ��q��Z���n�u�>͘!"RV��)*Ц�3�(��d^��`TNFu;�tau6�3
� �����Ѳl�fK��%XU�R٫�қfԧ�j|(n�j���$!�6v��*aαjE��aC�`r��m��)��:�`B��1�V�]��/M�X��A�6<g��J����K�P����ܔ���(�j�{�u���;��I��N[M�Pm�K��m1�m�t���[��Mqe�d����h��(h;���n�z�I�rV��ql��k�����RA�-�e#�R�j[6��j��Ѷ�k,*�Qƈ6���|�6��Ǵ��9�S������GIl�g]�;3BN��괞�Ckosp�Xi'
)��k�GI�o("�X3Y��J�����F��! ����5�RA��ţHu�2���,�`�YǴN�F��˷A4'{�K[6��q�Z.0%��SA�z[�T���K1�u*DbZ��U=����$�m��WV�d�$��S�2J<�N컦�}�6�bb�ڒ$��o)�x�c+v�H3&��M�����|��e��t�� ����ѷ�κ�"��t*&"����$�a˻�VcKt�
���[5čk$ޤ�)��J�g*Q�TX�k�X�����6*����մB���HM���f�`j�X�2����diܶʩl�-۱���a�g~ɭ�:�ш�.B"�(ˆ�C���j]���/DBX�yc�Yy�M[2�.Tg���b�sGL-=���2}mZ�c*�ų[�	��!�� )V����f�2��z���ӹ�#�@\;/L��1�4��(`�fj�jB2
���V�vP-Z��j�a��%+"�ɘF�ff��e�N�TձG+
vޏ�mI(�T��Y��T�o8�k��̴2k4s-r�{���in�S$ʻ4״UZ�i��Rץԃ^X����j�S��i��`j���/`�p-zĄ�S�W�N�l�+)�*(e�31dS�QѸvR����ٸ").V�^����_L�bD�;��u�0�2��I%���A<cdn�\����d�t�6���a�`_�!l�.�2
X��-��m�K�6m�I۽-���;쇥g[{%��r���]h��̢�p�a:�n f��ļ����6��a2����t(��x�dH-���N�k:��Kic!ޡ �͘�F)�hn�1�]M7�)m�bC�DF*���UY��I�/m=���p�{,��%cE��Λ2�pҧ� q����(ڣ�]ꀌ4RTP�8&�V.��uc6�0�B�mD�ֵ��
�M�%F݇YR�kha�յw� o()���m�uu;�U(eE�r���,�{���l(ګ�rV��^0��UqiҨZr���$���V�/��L��ʽ�uj����J���iY���,2�������V��Ÿ��.�����7^	[���%kV��x½��x�f���&�A)�I[k6f5�Zգm�b�M1��㠶:6*�6ci�Lݨ�X�̣stT���{��cDc�TsZ�.��Y�7*�y1k�w2k�C�qT7Os&��`�(�ŭ�C´��E��y�!��[��W��R�4 j^#�Y�W�{0Z�E	�� ����`PX�&v�w%k#,�Uhj�.�Gt��N��� ����۫��ϊy
�̸��֚ak�����V���6���z��)�	P5�w1�SHӭ���A���A�6���A�H�r�
�lDC�L�e�
^\A�@sn�^�k"*�h�U�C�(�й��͎d0}�+ �Y'i��-�#bQ֐��:��6[����7ӥ��4n(dj�bS�0�������qy3&��yRީ	�8eD�;wWr,F]<"D��@qZ�ᡊX��]��@.���7jC��"�am��f�
��(<˦��w����(��܍+�Ð(wN[;Wt`����Uܸ�!^5{(8�&O���3��V���ں��P�A��yt�`��p�EK��80��Ѻ��W�*�VR�!3��Gq����3Q�N�.���
� 9<ôi��5�5�4"E�/��HڃomRiZ*��2�����f�LR�5R�ܗqbck]��٨�]�7Q�r�5T�O�^�K@�a�Ϧ�N�%��[��&L�wH��F���E@��q�4	W�mgg�F���A�Yj��3e���+����7��YI��1�M-	��D��0����T��^��QH*T��we9�R��U.ӄ�*�Kg�o$6�ܬ��n=�xҙ�Y�6�7Gu���7���8ڛw�D�;�%*D�V�[p�,�`�D�'�t�Wa��ڵX˔��W�c#?e�2��w+a�ZV��2�W*R/*J˫�i%�+z��/�-f�RGr�\ʉ9V@%�NJ�	`��:TN�����;��-YE�"�utE?���a;oDt�b�e�и2�G�u͑�Ι� �΍bx�
��""�����FV˺��sU*/V�
d$�6p^x��}���hJ�����5t�����-�?�0�&���Q*�pe��I��Gb��1V6� ����K&��۽M�`��F>a��@��C&��Sm"f�+a��4M/�<�`}��X1��`�:���3`����x��n��"��M���%%vY�J�J�v�LkQ�P' 9b�S �����Jx�M��N��:ǎ�7wBZ��f���8�ݍҐ�t��Q�.�V�P[	F�Q͚��wf:m�1� �nm��f8�uj
wT��66���F0�۩��{��+U��^�pA�Et$���#O
�5��h����E���Yǘ]����l55d  uH[�yImB�����Ka�W�Ǌ���v�YaR��^Q5uaS��f�t�k�I�,Ǯ��q����t62-L��d�mdX�J�m�H�e
������\�p�����bN[u!ݚ���F�ml�,��d�/NGs5��c&���῕I����=���m��� $m�##��ETtiޱ�iU�#�J�{m��Eyl���F�O�ORVa^��2��]�߷n�v���V%P��-�:�4� -�P��l��В�l��*(���t%��0�l���D70/h��v�a�@y0�'I�5�������J��`
����f��IV�MG)m� n��%��scw��,|v�,-�l�r��yw��۶qe]�J�r��۫�&�ڶś�Lubҩ�e�+9G�Vl�d��p2 ��uۻ�s,�Y�t��LI��J��r����^V�{���d[�j�!
` �D= 9YE�q��u�̱N�]��U�޸��w��ě��m�U��"�)��.���s�lؼ���1����-Ȅe��<�`�v�TA�J�C`M$���q#+]��Ae@>�9jӗm��-x,�0�!�Y�H�;�iMf��S^+Cs�t����y�F)U���1M+�YN}q���c��X�T��6��n�t5GZ�1�:YG'�Ӣ���O]���æ��r�j؛�1
�M]����	N���OU4�#SYC�Xg�fC�܍9����f*����+�)ͷ�Q���g��t�`qz�4C�������^�im�`6,,��f�����|�r}5e� ��۬�5X6�ܷ�H)K�Fg(��Po0�u�V��J�H�i����Ǜ&<�&�h*�գ$���[��zt�;2��C�´=�-Uʳ�qP�7(V�X���̇C���`�V�/kU�,�⬊-%��7J]ހ_��c�H!X�XI��f7��cl�2�Gj�(�MQ�-���ǔuˎ��E+m�yY��ۈ�ur�fa&Vl�RB��M�#�f�ہ�7C� ���A!Z��V�J�JJ�� ��Mm�jD�Pdv*;�Y��c����2&L$��7�j�PT�_$f�ut�e��C{f$�E���f��"�nP�z`�v��Th2\�c*���U���i���k+��Sf#�]x�1ҹmZ��t�����d�Q���u��3j���M3lQ�ܲ1�IӧF��Rk~{M���ȁ5s�kr�gp@��r�n;�:��3cيT�u���a��z^X�ɗ�6��1�)�RܩI��\B�sjQ�Y�iG����y��W��W$�������U��,ݵ�X4��U�w��1�2���"�e����7Q��L�1v"lǚ�y�]��F��b	�u�aP8oCu/�钮��ZU��$�SHyQ�� p)��n``�q���cE<�׸�n
���d �q��m)`f�	fF�^�q�PW&�%x^@m�R���Q���i��cr����i��N�C�09���6|�Yv�{�V�M��Y���v�`�#b`V¥��E�ͻ�2�6�Y���X��[���U�c8$ٴ�A�ۼĜ0�V��	N�FеY-*�V饑�o�m��xQ�v��o.�
%%���<.\Ú�mm�F��߰`�nh�'%H�Q���*�4S�9��Jbg�,c�e�.�׫2�fXB�4�G����!@�L���mVޕ�.�����iVK�f��x�׊ћL���]M�ցz�gi�A������4��Th�2]1�^�RRt.���7r<X��7M)Y��̹CK+(^ ����9B��wLCN�8�n��ٳV�T�up�,Eq��X�v��0�՗�����r�.��>����66&ĳ-V]�X��%��j֏��]f�8���sm��UwV.�s��ͭk)1x�Q
�)�v��X���*Z��b�q�r
{J:���St[���9�BwWX�z^ڗ�apz2�N���զ��w�um;�鬩ux�3 h���˺[LӘ���`���h}��[j�d�5V��U�ۼy{r+�.DvZR�]U�
A0f��Sm�H:/,��
 a<S�)�afc�E�m=�G"7�b(FX����S%֫{�f���kYc鶶�&3Е�V���D����)��U(m��F��Qó4[h�iT�T�ռ8ƭE]���0�=فջ)jY��4^��x�o����G��O�X�n��7Y��٣[o@s��f��S#g�d�.�mn�O�a]ݪ�GԫE6��4�YH��y��Z��f0��J΅��9`^��ܠNWu=����ĥ�y&<1�45��Q%{����h7kP)��{R^@6e�ZQ�� ջ.;T�L��ͭq�)z]�jP*�]��(#Q�X�N��VaZ #E��:�VM�4`d,��vC0�VcF���	C)��P��l`-�[.8F1�w]�t��q��ff(@���D��klޙ�ܩWSD+Mb]%��H$�o^ZEV�T��5I���p��Qk���H��q�Z�Lh��F��[%��a,=�1f����W��f"�ݱ���;���H{b�Rp�{I�v�,ƞf&�ۡif4V
U`a&� 3��.��~YB�3��@��˗Y0��A�
%�b$�Y#�e(B��m	�^��+
u)ޘ�cU��%��cS����Zr�)ٹW���Ո��-��m�����ukY%J��hI� .�h:�A��$��a�j�jN�=5f^���m�F�8X�3abaIt�5�.<:fܺG�.�n�R�ݭ�d8�Xin�x��ch�Hk��5����òn�*|��n��1��n���>r�]�t̩l��B�+,��?k��6�#N�iBɗU{�+]�tv����1�63�f�l���^�);á��R���8:qfz�h��@imKR��#�n� cef�B�\d�{�^c����X��o�Y�)�W�}˥`��hV�8-Z�CL��E�u���f��.%Xɖj��NC���o`0^���߰<�T
Ä։��-lnfb�JӢt���
�c;��NF�nV)�YZj���;:R�ە�O �H��sU6o&+�L[F��D��-������gA�c�+.����I���,�cq$��-v�y�
g\G�:�\ι2Y�LKTn�u���i�Y�*w�L�R���b�͝��9:]�Xr_c
Ɣ�T�� �2Q�u���mZ��떁���W�js�Ǯΰ��Ek�����g5�yA����ϴ.��\޳�����(o2�}:pn���e��������d ч�p���BS:3���f��iC��wq;u'Y�Z[�"���N�2��s$�Og'hu�z�T*�^�}�!�����ϝv��7�#�KaH�r��X��0��?�ގ]Jm�ce=���ܠz#1�+��K[.��yBtǳ	��T;X��_k�NQGA(>4
`��ギ�}J�� ebyS��UvQ�q=XT�|�'��[�gn�2��g!�ew�2�͆-��	Vi�����5�t�]k���vBql��тB�#�xL�<�e�� ��T3-νѻ�X�����V)٤]huc�eW�)��QKi�����p�|Iq'i[��yڀ�I���[**�m��� R�)��ms��で���Es/���{m��ε��9}�¬���](Vd9�el|r���C7p-���_�d�s@R���kf�N��kl7���h.�ῖv�%/��\ݳ��U%n���0�w��m�]g ȝ,�����ޚ�1n��Wp��98��!y�� gA܊[�]}�sV�c�Q����U��W��D�\]�t_	͡ϵm�v��rGE7k�iLf�LPV>��9�n��Jb�M��$��V�]�Xۇg�J�_S΁���j�W�h�c�6��K"�Y�a+�WƮ��̬�D�����'P��wh���K;t+;E�ԭv��d\w��^�)�b"Id��� �]b99�^7,j�G���oRT�I!�Z���=�b51Os�fY�#oL�E�R����2�_>�֝�Q��J��ur`e�MU�J�=�B�̕��ۺv��@౨a�k6�sZ8����ae���hᤜ�����=������O�����D�^�TED��U���!"���9Y@4�;g�us2.aQE��������[W�m�V��ˇ���'���sރ��vF�9�@�kRw`-�2T��'L��,��fn���������d4�d�t2�l"�k[��4Q�q����&�!Vp��k[�]�aŊ��q��d�J�ӆ�o	�lW��!��J_Qb���o����R��#�-�l|4�v{�6��a��X30=��*{'�뛦1�����)��e�9�[O�.�b[KM�+�/@ۡ�0]�9�]��m��:a�2X�'.����G���ϡ�\�Km�:t����+%u�[�2@ֱ�]�A|�9s.+Qi5i0vU��<,sq͵k_	�ΐA͵��f)�b�q�4l}G���=��>䢥W#<^=7��[�K��*+A�5�;ҥ� jF�W �1�"Z(�f� 3t�o�W�m�'L���m�J�i��Q fv,EU�K�tns!_j���^���=ŏT�":���u��+T�M[u��A{��=�Nv��mauA��璋�o����;�y�Ȋ�:�Aw��Ԃ�P�]�)���6�f�c1Z��q�j��q���˻��u�oVi}+pd%�p6f���ڲe�@�;�P�-ʐ+�N�&k�:�L�KW���S.�v�l������Z{��JlT
W6��T���g�
6;9�l��y{��)M2ɴ��d�[ц˥��ok�G٦A���G�#l��,�#��o�Q����S� ;T�tXo�m����Okg[願!�a�y�սv���'E[s�S�cB�V�g!)jt�+�i55۸����S/�����s�z�*˧Z�^7q���΍a�)Uؠl#]��T�ir���}c8G��%ZR(��o�|����Q��7�`�]`���o�LR��sêG@o�7�^�(cDbW��y���I��s��sO'n�����T��Del�q���V}����E1�]��VPr���8,�i�s}�l�a�p�ctij�/�mE}{��E.�F�Eۖ� *\H>�Qw��zqO09�[��z�ut�����_>)�:#��3W!
ø�eTRq��1H�������MZ;�%7,X5f�;F�C�*m�����&a����*+��l�*ﺎk��oo�DՀ;Q7Ջu-ei�P�u��'A�}�]�w���yٹ�X��#�u��S�	t��㌘0�a˱��hn蛮���{�k��U���~n�dv#QS��U�cf����q����#�F��@�sQ4wu���7�*���G��9�*۳yv���٫��]+�}Y` ,��aC�eY��w�ǋ��њˮ�-�;���d'�e�^�]�rIcYXʻ����X��*tۢ�],mk��\��4�_pT4q�g�S��5��B��R��2��Q���t*}��z�sB��1��h_<kTt�o%��LP�lU�o#���)�Ce��1��ʱ(Ұxu��]g0���
�Z�R�$��wO���`�gf�ք�D�Z�����F�@�坙+��fLm�����}�G��e�.۩��z�u�}˻�Ҝ�o�O��16�b��T[�.�^�u�����,/���f�[t¢�U����TJ�t�e���%�.����NiO�{E�TS�����hi�z7+x�L/=t�à٣I�ݫ^�	9p�;v��W��7p����v�cB���$�_���z�r��M0�r�ŝs"���vl��}x>��j9Q/�(Mz�l���u\��$[��wC֢
v��5owk'�v�L�	�8��]�]�Y[�+m�������DB�����9����ُM���d�rg'H^�t���bh7��a(Ҷ���@\��y�Gs�����5P��k��V�3�wV6��ޑ�<�ǡ�RuuJ��0*|t�p���Ԧ�Ҿ������H��C9��v��Cl6�>.Z�4:�Q]���NJ�������g=(��B��⁺;*+ـ����&���ǻ9i�YB�
�ki%+�3J��6o}�GfP�[�7�mT��uTzMs�3z���ݝRЛԛG`�@r�]�{L�r@�۹%��U���)M���5J-k�z`�=;���T���|-��r�Z���Q�'n��ĩ���2��F�[������u]c��n��dvp�)_s�<�u/g
J��;�(Up{N�e��[�V'b���+p=xf�4:5^G�5��$�r���ӫ���y�U��b���5|;�Ǝl���5&6$a7�{J]����K��)d�&��s�����$H��I�G�b�,�8Qgf��|wQ�7]R����m]���n�#�i��J��]��o�L/2��6���
lV͢R���i�YIs&�}�|NԲXhP5��ODЮ�C�Z.p��E��w�X ݌.b���6� ��]E������JgtqѨ��wnP&_.�6�Ti�����.Fh��r�Z7-;uy�k��m�W�=��lPu�����gk��ǻ��S's
ǐ|f���_Q�ﳛ{K�L�k"=�YեO_τ���-l �8'�s��C��gi�|�m��Sj��k5r���1�f����ko87���Mݝ�rZ��wl��=�mT�'�����K�KY����[��e	'���Q���IE���N���ӌ���`�)��|�)\UCj\w��Y��e��u� �V��z���k����X� |���-��Z˲Eg{Uʕ3!�MM}��M��F�Y�s@n�U��,��r�JK�ƊK�]��Rt[}1v��h��>�b�y�FgSˑs΁���,�J��.��a!��"՛��:��[\o�f]�aH�ǒ#~پф:T��us���irճ�[//�ps�-�5��V�)��o4
2���f؏OP�ī�&"�m�\/����eԐ����
�lĲ�q��͖��N�3���bõ��<*&f���С��1Lح���6Fj�Y���e��ɐT\�YR�g�jļ6�u���]C��&�I��{w��-ƴ������,�a�3$J�P����FK�9X]`�� u����G���	|���"�99��{�p�U�Y�b\QPiN�k�,�r��9
 ���k��&/2z��|��59+�3��Y:6�d�l"�K%ٙ;gWJ͗���W`)��0�X"/q��b��ڌb��%�}c���o��v�M�.�u5��YZ]���ܷC�Gl����l�R̛���@Dp��m$a:�q��A<DMә��+����"GQ�xv�9ե�˯����+��E�gƋ��ث�.��p���L�U ���yR�A�nZ�WD���k�֤��;W�AT�V%����;rj��r��܁\�q7F����V;*����*�En͜^�U�K{�Q��,u����$�6�u��ք�`r���/�YT���T�#�e�7����o4��VƗJ̺����NۘhF��-n�=w��=�}BJՇ^)�kH9�ZF]o5W[�R���	bbն)�a�A�Ԯc�w���u���juk<�����Kܱ%��M3c&|!�U)Z�kU��n���d)1���Ͱ���;��]�]1Г(b��5�r��|9Hq��O"p�3�}������J��!S��L��+0H�;z�<�̙l������,���+c����C1�r˓P���:8�=-����pe`�ML^�-wO�r�Am�����Z���N��3V��Ja�мB^"��3�����m����ҽ�{���{�ֈrbW��t3-s� �ƪU�t�ҹbK�Vp����g%�f�Ӂ�f�.a$ܳ����2�gV۩f�͛b>ƶS�uj�{�'������t�Vk2����X�R�:�F���}}s��� {�I��c'���k�0t�;����;�����(��h��Ei�slp��-��Q6�<�N�
�,m�SuБ@�lZ���Z�aʾ3�-Z����V2��G���0aGz�Ь��8�=��a�*i�.��a��Pi"2��Ս`�����I9�8�������]�ti��+Jg-<��o���e�}}�E�����qss��Sv���#s�$i�pn���w_#�l�w��޷�uÀ�G���$S%�4u�4h��T��A�����\E��%��.��U��h�b�ؾn�sU��(*�G��=x�,5@�I�#P�����h[ˑ�{��#���YY��Ў�q[�]�Zx�k�� ���X�L%W��h�[ӟQ��Ե6pɼJ�:v�m��̷��6x�G��̹SI�N��*�[����n=�C����.A��=���vkqw�'Y�ޔV�Esu%�,��f®�JW�2NYKx��:+b�ѕ��R�݈��;���v�5���ɝ/�vբz[0^�u����rW)=��u���0)��Yǧn�n���(j�_J�cn]vQx7��U��G�-��#[�v�����a���:�q������&W�3; �U�
+�[�ȷ۰�����R���iL�
j�4O>׆��87��
�t!����q�^�n�7������wugt��h���ɸ/8n���>���Y�n��d��G1��5ڇ�R�f�b�g W���[���߁�k�]َrf9�F�A�O]!wR��Q��Spq58��\�|��� X`%�H�����W�+�K'm��Vw���;��I�k4s#�0��/�2���r�n��sz�	ATR��X��tt��c]���j��Չ�1%����UY|�u�ڙj���/U=<�5�&��!+�l_)V�t[�Ԑ�&bO4&�v���z�[�K;_:�wد����-OK�͡�ݹ&U�l4oQ�U��m��� ��^,Z���;�|�{+�.��� ��f۴:E���u����p9��P�����ř�U�g�;����KcrT���d�;���{1�Q��/�Y#�)Wd��y�]ow;V(�9D �u>�|��>���vs/w���������N��۴2EkW�wy&�{��Օ�7S�{��
�O�U���[wF��@���L�@T�s1vxbo�e_ui';-�����ˋ� �+�A&ܰ���,��˻��/�����򄙘6v���g SK툮�k����^sx��x�G�oo�r�� ��o.%YzҮ��%@��ǜ�Q�ö��p�W_[��l����BwS��Eg�3��B� �&��J��8g�ʞ)�v���s*'�$غAG7���*�b��7�ܤveL�ַg����O��ۼ)��a?��L ����d��e:��u�Y�n����"=npX]�*K��rk%��K�#Z8��֩��sgv�^!ݡpu���|:N|(���Y�r�}�;-O�]�2#<ҖVk�cf��f�B[�=6���H��Kk�m�7i�Xs�55XWK��j�z�uK]�t������̛��gK(P,��s�Ԧ�û��W���v๙έ*{�2���h�̂L��9V:��J�㸅�x"�.��k�ӗ�k[1�L'K�%>��՝s�GWs�YE�#�xw�0�j&�V�`&Zh��n�����\�u�3��țDO��n�T�:���f`\�gX���ݨZOyo`	|��T�&�X��C]4���WJ����n�AcO��k~d=F�R�ځ>�n�9�:ʹ�+a��4��+�˕���\jr��}im�bk�c<�o[��,��t�n���x�:����-�d�����S�h,9M�;:�����ۥ��;����m���m�km6�m���y�$�9I't�H�� �$�"2K� W�>�����HH IO5����߹~�-t#5��z�޺�B
����˕�ռŽ�����(rѲ�e!95���[*�J�	�i�8��[I0����6�V!)4�)�t������R��s],�]����S�=�����pFBc.L��<6	g���ݬXj"�<��+�
��s0�	�GJ�Im��U�G9�0�����\�ܧ(e�e�uor������V:��PKB+i�.�AY+R����cvR��b��?�h�Z��uĵgnƱA[�]c[:�ThH�]����X{��Z�z���%"i ��i�,�����~�b�=:��V��5���MBk�WV[��V��ښ�mf��[|Oڙ�Ft!5��<�p�-��Dŷ����R�y��m5t�;�[��5w<�k���m�d�fZ�_E@��Si�]|)7a�Tz�W.3��Ss9�fYΠ5ۛ�q��̩�q���>�
�T]��.��xye�`o%� PHGlϵH�6�e|�c� �o�\yodz*��U��]��5�%���k�ȭ���e���Ҳ����,��\#�,�T��ԇ'�fm��#�y��e�� �f�\S[�­ j[���*M�z���NY�#�W]�m��WEts7�ੰB���PVWp����I��t�0��9l[��b��;�x�;m���t��]7&rA7V�6z[P�ZV���Qh�N�[Xk����z�OSI����J<]�K�;Br�����`V)\�wr0Y���7��
La�-��wm>��e:,�W��T�u����ʍa�7-���o��N�%O��}ʣcc�r�Ӏ9q�������{Iř4&{�*і&!�d���a���qV�,�&¤�����v:�$�3�V�*s���.��(������x�Ẓ��2�H��X�M|j"(!��e~t,�Z���C�[m#�B�Rw\EK���������%��K��,p���8	����{��Mno9���YM`.�R��tJ�c�>�_p;�Kv'k35��)�L�O9K%��+^����kfC���<��3����ǫ���dU�ʓC����-��-��c�Y} �oj�xѻa#�79.��5%�x�rs��p3�x&u�%��i>��FRa�VVvZ��l0����1ӫ6�4f^�j/;H�c��z�������mmՉu�ۘZV�nmsϲp���wۂR�5pG(˩,�A@��׽\���XFښ�b�q8�����T��җfr<DB-#G��=x�.p̦�R�r���9O:+�yܴd�V�`p��)'(d�[�+�	����ݹ��K�:4n9^�[/��W(��"��1@��|��Q��[B��L-̓)N�EV`�'W�����5�ʢG�f��-��s��Z��e]��|�ˮ�yϡV3�e���3��N��W��9{b��M*u�Wuv���|N`Z��*�գs��F@���К�GtK{��u7�ɽ��&���d�4N /�!�kp�u]��Kzޚ�|hq���d1���kѸ"��
%�U-\�8X�i�\�F�^���©0s3i���ܔ��,ᰁ��	��ts\���:�2���FT��r"H��|"�����Q*0+ݳ��.�}��Y�w)�3m뼾s
�5�(Tp��O+[ڍ��6�Y�r��0��;�ްj�-�"ϵ��]�'��N6y�*Ɠq,M�3uc`�	F�07u����qޢ�ټ;��`M�Õ�+�R���wZ��d�2��<҇L=:ݡ`�$ԟ�-�::lܺ۬Rr�(*��ӱ�������G�f��G'C2����L�f#<���:�OVM'@�P	!5�
�̾[�"b�p1���p��˵4��L_1B��������s��ޓ4p}۸9S��>ѥ�3�1֙`���r� �,��C�����=znX&�D-y@��؊L@f�K����D�2ȳ2��üu���m�,��NUn�ʽ5Ii��JPf��ړ�^^���ݲUt3�f��rMj��ɍ�������,F�7nʼU�N7��3,7��Km�ă�sV�Z�d�[R�5->Ә��jkp+��ƌ|�`�WM��Sp_]��[,QZ�Gb�D;������+�pe;�q$���*�3�7Y��(�i5�b�3S��j�n]>��WΟI�>�)��xl�P|`�
���l��7�3��r���w����a�Vz*%��7��}�l��P�{Q�Cyg�K)�ڻ��w*����m��8^ԵAgZO�o5P��׶*�
5-e��ZF��7WkhU'Ca�Xȋ�V�q������Z���-�FgY�ַ��j,@}��ح�}��U��b�j��n��T�n��(����ѣVHDp{{[���K��n����̇	ĳX��S��Q��z�ƐI�Z�#1m9�(�{�H9.nֻ�U�����x)�;[�|�z��
�ZTJ���Ƀ0R���Mt�iY�ې�N�9_*���]d�}S#���;7�Z��J�N�I�
r� g��A�)vb�b	��]���.EÄӦiJ�����f�Eum�ux�Ć�= ]h�m�Z9}�gNN�n�v����7���i�9�<n��In��s3�p+�ۜ���Ҿ��	j#��ɅO�\�`��Ya�bTy��Wn��W]M�df�o{^Pq��9�B"y�DǪ�=z�5:tN�2ҿ�U��鲝�0�9TYuy��Ec����e���f�[o:*7,�̃��_��J�E�<���R�Ǹ��Y��d��]gG��wk#5�bf"�ކkU:�vh�P��NC W5q�&GX���[g4'͓ۅ(����EU*	�^m����˗ڸ�=[����	緻������q2ȷ�U�a�u���=�h&���S�ˣS&D�w=L3%ک�Tw�V9��r�=&�ט�|z�m�t`z�(�vs��v^Y�5��pv�ڙAչ�'g���/c��,u<�S	�RnH�t����	Q�n01һ��.nDz���]�Fh�u�kL� `�L^��H�zHe?����E=K��5OlЂ_N��f�ti�)9���B��X����fGeh��4S3`<�j����y-p�Ǚ��6�䬲�P�GW=�Em�ظ�ve��j��o;i���q
X��u*�c���L���<�}7�C� ����#������j����E���U�s�����v���guL[��Y.n���`�#�8��j3���$q ���}3���G���R�<��2��@1ճ�%�jj��a�Na.�����h�@g6�-�෥K�1�n������k�[�e'�a������p��q7�u��)ĺ���{��[�S>��9[tc�jG�yJ��hm�����]������ �b|�)V���ڝ�`*�.��ˆ��1N�,.��-�cj
����u��-=Ժ࡯�MwW8��p������'�7hb�&��ط�6�Y�ꓛPҮ���P��o�W]]7r��mO��V��s����T&���㡈��@�x����v��ԗ;A}��yyXr�3$ޠV��,\�S|j���5���Ϟ���Ro;���Ҋ���x�vf�S�*1[1�)�>joR��Au���˼�U�Ar����ڊ��.!���n��泇S���_}��[(�!�ڰ*�l���wcz�y�n�i���к�nƁCS�¨P=/H��pŜ�4g��tH�i`�G��l}�e�&�	33���C�+�r�Lj��R�@袹+�t׫�qd�wxԝ@
�vڋo3��Oc��Ӗ1݌2�v��W�*�e���ݡ˜����FR�Pp���|w~�ͩuw/Dg[4�ȭ<�ƨ-��"���M��9l}����*���+��
��c�1�7�HiJDv����)n��Z +��]���@c���'V/K��<��ҺÊgX�IӋ�bc]``�9�WN7iȳ�Ņs��fڵ+V��t���%q&p-7��ttn!���볅�
����Xm�rn�9�yK�?��,���b�,[}v)�b^=����]��T@-��3.�941ǒ�@���.�k�5ju;Y�{:�i�����F%rF6�幽u�1��dy'm6t�]u�s4��C�Wb@=y��\�C���*`�,[`��'SBQ]�M3q�aW��xmM�R�E��|m�0�����NdT�I��t��o"�y$.���S�/� �>.c5軧^�%��K���OGXڈ��ѭ�ΰ�)��Mt��y���oZ�u"\��i�>X�p�l�Ҩ��]ۋ��ǹ�ԙo�Ǘ�������y��β�E+���Fp��[w��!P� ��1��W���<�`�A���[����;�3H�g"cޝɝ瀟��n��vNUР�ލ`�2�d�*�Q|չ}�X�NE�zNvW��W�&rJ����eg�	7U��qj�i��P��KV��T��jm�G�;o8.б�\yXc�
���m��_Z�u�s+�v�U4v�bwXR����G�[t�I<�-�^p��up�)܉�i�[o�L���F�i��g�a=�
��eL�Mq�5/����@H�*��6Ա\�ٻDl�����rҕƥ���̉�<��]rj�#�t;���K%�F�	�77��Gv�� �T;�6��� i����f���"й�S�!۸-,�ئ�������X8����	��XP��vz,�ǝ�U����mquI�@Lܮ�s@a߲���	�4S��f��Of�o���+Zڙ�t)�Gz���ӧ�����["i���Tni������'�V�ab����L��9�CMSj�9���3Av�]���lq%b����v�v*r�$�P�,�����p�c�u��*���{Lp4�ꙛ��s�m���|A}�R�V^P�دjӜ/����Op�#��=���yoP�d���U�v�j�a�tG�$ѐ�k5qۻ�&��Is��#䢽�A�Է�n�c�M�a��uf6�@�u֝���2y��+�J�o��Β�^��^
�x2k}�W���dy��(��v��^��h)��|�UoE=t탫��B�t�L^(p�ǹ9Xq�m��^��֜��w.�¦Z[��\�$���yf
�R哇BzJ��)�t�ʗ��v�����r�J��&�1���ќ��C{Y��-h��g��Z**MqW]y{��j��G� ƓG-��lRW�V��V��=�"���s:�)��ЭOB35�:L�C��������l�5�뻂`�fT�ᢞY�q�ӽ����J�mМwssw]�t�Z%u��4Y�����rz�8��:�;��xT*Euj�Ny�t�oZ6˩�+Mu���iiqqs;�����
l^p�O
�zQ��ttѨ�v�N��I!�r˖2�8�G7a	��hS/r�K �x�['R��;�&�\�:݃� �=a�3c�ܻ��O��\��q����̦���=8�����Ӵ���@�������ڒp��A�;�!N�����.�G{��N��$��L!�M�8�R����վgb;��ٌm˶�؊����u��wض����K���rH�&��T��آ��э�����C9�Â�]*�*���Cc�����䒖�i�<�ו�|�ɝ��YԬ�p�賏	S�q�+.�ޑ��k�*2�C��n����2d6U�ևZ�6��*�'�M���J�U�ɴ�;��z�ԭV�N���>�允J-�1S�7o� 2��f��h����633`j�p���� r��v�s�׉Z%6z���6&P:9�d����݌��Zu�����bMn���=	<����-�[�IL8�<�[���odnݎ��Yg�#�������ǖ�̂k��c)�S�gas�R8/�d`(֐㭻V���Ou31�t���@fMw+��i(��os
48��O�\�X���3r�0�Φ��Y�����h�}Ԯ���>���hԥ}��nL[�˝����b��3w���][Y��6���r|Lz@Y�<�{��m��+�U�-P��g�����iYr=Qӿ�F�:��mY����Z�\��gi�Jm}{N`r�<��]�Ŝ���I��K(oT'.�J�w����Q�	H��En�c8Wi��}2��v1�W��y�V��v��ں˶�u��5>�}���2�[���S��޻��� �YW�j���fhS�ڽYD��eZxbv]��ͧ8����
7�9*�P�`d`Μ��d��,I<L*�D�X��<����G�09[g	���B,�*s�b�+ϲ��M�S�mM#,\���9c�1Ţ�1�j-�����K/�6�Gcy(1O4&%��ծ��
��)w�����R�����Q�ڲ�iv�!�̷�N�ZԵ��5�&���v�.�{��^4i:��i��%�3J��*WoXi!��O�䠟!V���_Y�E���C%7X��I�W��qJv,OU��-⎶�`0�q�5Q�mc��5§	r���p�nN��J�×�]VNP=�j�{x �J���C�\f|�VZB#W��K�,��3\k:-��W�ct���v.�I���;̈��b���ھ�lL)Uf��g��|�=�䣵���*c	�N����%e��6e�|����%�M����`���7lg)�*uM:E0���e�k��1]���t�
�纂�(�rWWxb�9� M��[�Ň�w������h�r��7���+Xz(���dG_	�Q���A��&Wj���n��fA1p��+�����-}W��GQ��V��ۘ&�z�ͮջxr�pTɦ72��3��r{�n�����|>���}��=�b�k�Ń�|���Be�NsgS,���?�5a�x�U��2�ed�ɽvs��h�F����ӖkRr�����v�EA�t�d����[�m��N�٭�R�U���h�;n�z�܄b�N��'���*�3}s����N���j*+G�$V\4*q퓞P��G�{���Г�ǻ*b�$z�M�[�J��"��>厌�L֬�5n���W�w������D*Sm]$K���μ6pN��7�uU�9�%�tMm:R5�r�x��Y>=�9ӌ�:���b޶._dglf��>���2�!2ؒ]�Mϻ)R����R�]�WΫ�)�-3��ߧ[�Sr��"��7�3%X1�*{K��b���=<����	˪>'�V�%�@�s���ڝ��^�-���e�76���,���z���s;YX(�� )},�V7��)���5{}���(^��1�-�-��I�!э5���O\[,{���x)OC���xn�i��Em7iz���FT�*Ý&Y����΋b�{h�m�}�)|��ݱ����/{�*��aN�Pc�$ivf�x�q!��d[F˱A��x��5{YK�t�ћ�ώ�u��*r�!����n�Kҥ��w�t���;S�P�����dmv�EY}|[��˭��ͩW�z��fP<��9��lׇ�5��dͶ�����n8-6��Zn�d�$d�$�I����Kh�E��ZUE��[l�Vʵ�Ŷ���+QTTJ�jZ�m�D-��Z-��l̹A�Jؕ��F�,U��0RҢ�6��+%lE��D���(��TV �F�eKk��KB��[F�-�iEW-Ƣ�4h�\jV����A*U�E�m�ecFTEF1Uj#�V",eh�QV�kKJ�������e�DDPj)�Arֵ��X��Q�Uk.Z�Ƣ�X��4�TF(��Q�*��[J���A��-�lX�T�V�TD���QTV*����
Ա��Z�jV����V(�kkDfP�Z���eEjJ6�1V����V����iJ�R��ѵmTc��*��V%ebm��Q�U1���8+R",U"#�)��+\�E+*	R��	��QA��j,�ʸѶ�dQ���aXUJ�2TS�%���!$�) H6 ʶ6��.Ӊ�Ys�30����q���K55���JqL{.����>�whs�3 <O)Zf��;'j����㪮�&tP.7$3+�T�Xzs����4��L>��^�h/�Qy\߳:߳4U�	w�.5ɺ���J������{�����g|%��AɗB`�U�o�����v��#0,�W����a�7���\7	�}��ϪeBītN�m�:�����w�����k/	��+r��u�>J��N�:��Ϸ��<�:��R,෵Rm�	�k���by��n�6h���r�Cl�ZP��쳿��^ﲆ���O`�p[~Wa��q����x��Xt�g�2��[p�8F�U8	���R�dמyCG"����*z{\�]�7�����.%¸�� �Փ��X�p��G�ۏ��!�'�ﻖ3#k����&([��ŦIvG��Fh`�sV�ޤ#�6��J�g>�t�A;×q~혒�U���1h�>:d��2�a�F����m�)pv�����Ӈл��־��0��T��A
vP`��EϽ��u��14�T>��C�&����R����M�Ǵ��6ՠ�x�P��v�L���eD��1a�U��F�^u��iw�n�]�C��P����|�U��SZz��6�%\ke[]�X.]k�Y˨��A;����L��b�Wdݾsk>0Eݶ�WS���,��ܑ�H�1�/	�jr\�;��t_]�tB]��Y��Y}W[�m����@¾u:�>T2٬�1?9��vmGĦ��#�cݯ1�X��B�먣\d�w�g��B�6kg%M���^H_*��c���˒ϫ������_[����ԱS�P��r�<(�y a�ܪ1�\y�9�G�A�{(���YD���7�:b���W��:�W�0�Ke�"� X�Z�'�L'׃owyCy\�Ln�{�˺=~'y�Ǐ<�t��,9�3"Zs��O+>��DBX ����#�h���^��w�,���`��b��2�T8��P�qf%�����������������ޭXCG�a�7������G�|Y��,��9�6��;Y�o<d�(>1'��p�{'PO���y��zƝC�"��Tlp���<3�O���,v�/�w҉��}�r=W��s�*$��"��h3�ӭ��+�C��^��u�0�<5�dI{�8����[��K��47\gw+�O�BБ
����t�����W;,Ŷ��I�D��Y]5#���K�n��D�Kw*e�t0���N�lqz�#Z�<�9fV�7y�n���i�{��ػ|�V������O��s��-�,��K�ka�B=3C��/-Hjq��"����Y��]��,����E}����k$,�6�Y���Sι�Z˒�ν�s�8/���v�}�%��9��m5	!|�'��#��2�*�Ї��p8�R�hLպ�9a�2�b9�(S�!M��u�<8t6]7�y^��X��h���j�{�##}Yҕ���~Y������v��6�8�n&f ҙZ|B���r=�R*)�F��{v-�b��y��t@{@�\B����^������w���xM�Ƈ�{mK[�i��~��� �M~�����\��?�QY]��֓/��T?7��u���+�[u�lC�3U�e�{�.*�o����@T��p���Փy�Z�z}^�W�s�=���B9�ӎo�y;=`tf��T�ϲSx��T���w7�^9�l��L��];3��X�X�U�P�<^{�����qP�au��3K��.y��p	������Σ(�i�Wz[����NˣQ�6+�*Z�ﳷG5�)�ӻ��*�����_�<B�Z9N�MSw��%>麙'Hw�rP|v� �u�+��p$��2.�ll���/���o����bNZ�E�Q�I2�2ʵs�]gg&�ȑ�����A��̇�w�u�kju�}Z�.��n���Y՜L��w�n�Ձ8��ݓ�Γӯ�[�[ի�O8+�{��Ol��S��j��]��C~
I�!���ߩ촻{��ō��C6���7L�g��5G�����r>2ؐ�	?����%މ�䱌nα~έ�^q{{�}�����<�f׶�Ps�WJ�=���\kt���Gm9�=o�����p�Ջ�Rעj�y�h��WM��w���q�%/
����z���.Ü��_TȀ�ڇ�������{��W�d��tkT��Ǻ�v_�-���5�i�+o��(��ژ���o�rEw����}��So�zu��|���I�o=�;�x�@���y�ZH���j��z���W�;cg���N�|�nL�H��6���"x*\i�{�70�U��%zZ�8FV7w:3O�G���G�q%���t���m�ٕ�B1S��q~�2�/+�rIȣ����Ss{����*֠xp[Ug�쉬X��òm��[�Y�538�yj��\q�X��WB��Պ�D�\諹ŕ�\o�݉�,�F�jי�_vj�O)�W������r����s��^s��V��/��N .�͔<Ğ��%�6`.s�N>�=�j����ۏ���,��t賭�Υq����n�.{z�n��9)w�q˓��Z��_/��<��+��g\T9��j�?`/z��=�Dr��
�o6:�������;<侓�)dW3��/�l����<:�6��䤞�zhxԪ���4t��2-XȐ04�����j��]V�ǗV�ky��f@���~��xe��H�K��扷+�e`��&��{�L�+7m�c�����u�dy���C�97���Gh'hr{��s{��fף��M���
�v}7fo:=�/���^y[��������~�p[=�tpJl;���AOT�G���of﷏ԣ�9�gǾ�>��	1p�����<zs�}~��8��3џKGʝ�qJ�
.�{���(�l_d�^拀ʚU:w�^E |\q�wv�o��eu.�t�ѓlᮤ%e������qޖ�``ÊvP7�Gn|�m��r�05�m���S�89L�v4��JF`�Ʊ���rQ��.ϯ��p�����Ρ:��U�秚�|�N�A���+&v���z���(>?�~�a��,��m��{_�IR��j�{��ɢ8��2�9��y߳��o� ��T�Z�
��MɊ��>�o�E1>��ϵ8�^zt{��G�'���-��R�(�|�`�M�}�{��z$86W����:���컩6Vծo���`��^��Cng����Y�ꭊ�����bB�v֏d^z�+|.t{<7��'r�f7���:tY���>쫗�w�4*D�֖����/��9��ml{����U��g���k��������S��G��s��~�1�l�S{-�jQƐ���+�З�������xf�Ƭ���=c���/����A�y�"ՀL��sEy�~vO����E��MGM���.�]ճ9�yQgaq{�G�tėU춽A6=�B���l	��9�R��aM�@���ⲍ�b=yK���v�
kK{�l��Q�[LrE^���Ml
n���[|ҳj`����C3����p��|x��w��RU�cq�R�.r��)�k�ιk�����F�����u���Hr�4Ml:l
s���<{pz�z��L�럛��~��a�͘i�@=��sTˉ�5��*{-[����[3��>��*o�9o�~?{oz�� �Y[)�V�݇�2�>�T�2�#�<�h�u��e����`�t^�^����=c���8�ў�Y
��Q;�/<�M��g;�����,�8olA�c⃘��~իeJ�:.�]�+�U7��^c���}[�Mz���c��4�[�y�VL����+�Vm���ǜ���^��-C#������p���}��R���=W�t���;��tk|��J󶂸�?LU�,��.���U�m3��>��m[�N�O>�$����Xr�i��z�;=l_�]WC���76�/��>+ �'N��{D��R=`��Q��q7I���`ػ�m�����S�6�˧������*�f�m��i�V�SV5�w<�l��ru���imn�U�ݥ>���F�icը�k���e\�B�!70f�Z����`�Pe	Z�_okL����kz��$a���,�m�JOs��R�w�{>w�~�@/oP�_y�=�'&��N=�jo����9���ݔ)�������>�N����ˣ~�/'��g�3C�o��L�ۄ��Z�y.�/��e��t`.EC�����{��.{��Ux/<�`��x7+յ&�YiMƹ����9�7\�}A������y�O��꩙��CL�5�=�k�������pR7��|�9� �j=y<8�#��%1��[NhX_���2r����H���:�,�������"�M�3,���磯ބ�����bC�6C�t��iN�{��"�kzfP���q�^O=�3��c�b8��}�y�t�9��*40ߟK�}�6^ӤpM:v��˚7�AW�q�^��2�����,W��b�6=�(����w�s�E�Qz�si	`��)����_V�gk[�[c��K�{7�`�v
o�N���B�]B��٦[�3�'�7"�����/�����nٮ�Κiu�EH;�t����Z�6&���ퟹr�J�7.�P��M[x��N��A�M�ݹw�[��ڰ�[�P2^�6N��q<͎���=#���7�'*��m#g=(�l��T���>�Nۡy@�^��:k�F�:���3�M������Ǽm�^�
~9y�����|�J��0�ɼ�N'qL ��`rG�
Om�n�?2������hC�c��aX}��^�g86xcq;�0:��&��ɓ�xվWU���wFd{��ʀ�܅m�U���͔<Ğ�A,)6as�0��$<Ey/H�zsǲv�Y�:tX;\���\�C��}�Fq;u�Mmh�]W�\�}���'dP�tY�0���f�e���ɭ��^p+���̿wd��ڛ�m>K�rBO��9�9]�hT�z�GH��Ӛ��=<wtY�[ۀ�<�L�:f�dZ�dJ��D�u���V���3vy0���_O�=��.�@��9�s�&	�׾�����\������WD!�p�ȥ��v&���{q��]J"����{I�߰�Q�7���蠩kp*����2tקO��k�z�?�1��۾����f����=�p�o�u@x�wV��=ãal����J�윺v�7k-]�0E��c���n��̏ 2ؐ�	^:�ۿi��u���>G��d�o��Yn����8^R�p��(�?aj`yA�]㇅S�;F�\Ϭ5m}�q���Zv��T��T�̲�)^�5Z}�k�Vs��ǧ:�/E�q��=^���C{T"�b]�K�ȴn�N�-5�A���9x�sڷ6!��k+�w�8�0O�\���U���Z��g��0j�B8�<�(ds��=���UV��֝ڑp���ֲ}�=e�t���Y�����:�56w��_�/��ҥŸs���ֹxr�x�U�hT�a1z$������s�o���::�Lfy�m���'G��7#�N�W����[}��$*��������H�f�l����\�ޜ}���
G�:,�j�Z�}�}I���w���၃�:`]|�Fc���[y�v�;�C��d�
����5�K�Z�
}�..����d;�;�+qݺu����o�����@�;����ףI�)���}�a��=~6�:��c��m�E34���4��["�J�T����Br��f�^�����%I���	<�J����	�@ds��7�+�N�'�u�e�.j�8��z�/{���Ū���p�-��K##��b���+wd7PN��|5�ܣ&�D���l�i1TKF�8Bz˚&��voa�2o�=4$��4�̚,���<�YC+��iK���)I�+��yF��J^g`�v��O0N��8�rdj���_;�Q��r�A�Z.#�û؎.�QY�\Bz�Q�r4iG�6Nn·;� �Ӷs\�=��7�*Z�̍����:T{{�<�v��W�o�P�(��dbu�w��Pܳ
��w'�ơAf�q�}��E��>&p��gY�]&i��z��?]Xtb��1Vv�%���t�+��HV�&W^�p��6-b���/纕��YGi�ܬ�N�[�4�,vY�9]��璍諂�T�1y�K���'9]1�����Tx���K�f�k`����/[(���z�ݾ���z��a\����Q(R�A���U�F�{��z;��y�^���eԲ2��jVc�K�9�ӡ��v��2S��`�P�wzS�'��7z�i���o�Bb-�����U�A�Y�yص�▷QҜ/d@e�X��h�p���`�����F�R@+�o��/(6�J9���*q9�ytל�"ű۪�a���Y���@p���"�k�gv��z7Mu���*e:��%Z�SZ���w�%�/��$�����ZގgS=4s��D�o�K����МV���WY��8vc�m%Y�gd!
Ѷ���sLlCj��Z��}۩J>�:���1�N�]d̨�%�����:��*���>���*��9O�v�LI�����R�p!ݐ��W�YY������;Xe%cR��y�6�.�730B�ͺ4�2x�ζ/���	��䭱�u�[��j�+P59ps�AR��L�74Ԏ� c���a[k���{��{� aܘ7���S�q����Ӫ�U8��V����%��.@Ļ*�>��Ljs�QcU̬fjhZ���wi%���{z^ּ�X��rVsŭ30�͸8MS��)Ĥ�\�9�|�<�_�z��yב��bزI̊�:���d���̲�s�0PUa�'�F\�r%0���ռq˗�w�+i۱��u����젚ܨ�����X`��,[,&��8�'W.���2rKn>�۷���`j�[G&ؼC�#W�Jw9���������#�̑SuÛ�ICS�ܳL�&.���%c�ލV;�,,�9C����'��e�v����u�]t7Jע�f͸R�;�;���B)�+��"*�eU+iE���ҁF)Z�lKVV�pC�EAH9k2��q�lq*#�V�\KUF#-U�ֈ�S�U��\L�"�,�e�E�c�[cmb���1(T�",T�,V �eb�
UnS**��Dkm����lZ$Ƴ*�dE*�je���YEQ�[Z�*6��3.$ŉR�R����Ab3�QQX��*Yc���QFV� �Q-
Dm�����Q�\�ƪ��)l���̕@�F��m�EUe�P��b�Ue�b+�6��!R)��(��F
�fY��Q�((+T�VJȆXTTTB�,kAEը#X�"¶(�[1���a����.5Si(��&[,U�!m"� �H��aX�Z�U~@�� ��]\�ܵ�R���P뜂�-���B�tPΊ�{ �/n��m�Tڛ#X.����夠���K3�T�]�9�9Ϧw\�~P��lN��#�ǧ���A�����]��C|�f��y~Wcn}�z�8����6,��x&ob�_l񒈹C��U~#`���R���>=�����\]�t�/���sS��b���9P�ưG��s�6������W>B���B���[3�s^Qgaq{��/�iw��c�����++z�7�m{���������|U�ib������P5�Z�)�}O��.��{��o�96*�xMg�
{.�xb�1t��	�Fn����{��|�l�'����bB��<�vhh�t�=O�y$%�s����3�t�~��������GBLzc9�y\�S٬�%�� �M��^�4A�*f�R��)���lO��⃘�����ԇ�O���.޿_y��aƾ��3f�v�L٩��v�{Y�����=���R�j�Y*��N�r�8�I�LW3��F���MG5ܙ �M���n��'Q�8@#5�����Z{yd�6++%��I�X��9���e����_b��9Ӻ},��ųV�u��3����$*A���{�W=��k��'E`��8rsa<=��Le"����߇+��Z�lgl��s���N׏%W�K���u�N��m�}��4H�o;~;hEy���u=/��|<�cIA��T��#A�Pt��$�s��Xr��6�z���d��4t�P,�^�ד�q+T x<��:�K����Njcy�#�t�A��S�&��&��S�r����8G�0�9���s����_l��_{���վ����O62Ͼ�r���'nL�vsUC�F�ҥ��������u$~�wj/i���ڋ|sِ{}Q|�gF�/�s��[=�O5ӛU9g����=��F���I�������Γϻ�]��}�����r�S��zc�#�l��f�y�~W%Ϫ �Dֳ������V,JI�E�=��ǑA��^�� 2��$7ྒj�K��u�Uٔ�Fb�5��ΰ�QU��
/+O�h�@,�j4�7�,�C)��`�߄��J�xT�����k4%��5�]�����C��WfM�rM[�Rt�!�r�z�l�θW|�e��0Y����Fr��wV-�qN��Ot��(ю���6� v�a��4�=w����ח��/k��9-�O9l $=ྐ��j�y�*���
�Ϥ^�'��;.��WMK���l��G���q��郰�p�0�z��t����[��چ�k�L����{<����U�+����Jt�����f{�t��}c��}�q��Z�����m��P�n���H4���^�)�Ҟ�)�{G�6��6k��z�`��B���ш̺ݼ�v�T��`�F�ێ��3�M���h�I^u�`h,���ߣ���3s2�K¯�ᝲ���)���9'y�<�"�[^{��{,W+���&t'�e�y�W�¾��ns��>u�M=��z�%Fjz��w�??-�)u���j�bZ��bO`�ԛ��&��姞�[��ɫ?>>�>ه�vz�:t_�5U��ʹ����72���^�b�{c+9G�>�
�we+����z�a�7{Yy�g!�z|�<z�
�wJ�=�*�A��u5|����GCFz1�G����������II�Yۥ.յ��h�l;���n橚�|N�[ϓ���U��i�^��eN��T��\���I立������;"��������.>�"�{5ȼ2wl�f]�����i�\�JO��9�'�w{K7RB�,�5�+��>�=`'�ry��y�3b���dHT�������{�(��c��l��l� ��u7�c2��l��kʊ<_� 퓩�'�nwX�|�����[��y�����������XO�y咥I;��J�l��e'Y>d��,'>O!�2u��=��Avɤ5��a1:�S��ԝI8��2q�Cϱ�͞^W��#�~���~���aP�M ��߰'�|ɠ߸x�8�G=�*V��M����N2|������!��x��L�aߨ��M!���&%a��_�o��s�}��]��4�OM������d�S��(q��5�a
��'��2N0ѿrJ��9��d���8��O_��d�!�i�M$�O~��=�f��;߳��߯6kz��8�d�7��	�wxu�by=�d�G;��N$��M�)>d���y$�&���W�I�����:��aԓ��7�޹���3���վa���}����gCi���q�2u��?j��<d����O����Aa>CG�a�N%Bh��=I��2��;�?2|����'P>?{���'̜M�U�է����
�x�s~U>Q���#��~?�m����m	���x��(�d��Y:���XI����d�i�|�s�q*�� u��ԛ{�?2|��<���n�����������Xm)�F�HY�R#/K��^��հS��D�t|}6�"�e��4R���*-Wcã��)�3������8Y�+�Ɂ7��e�Y��L��ɮ���)��=�T!���{�9���j�p�4�Qe�#]wl*Fv�B�iV�N�2�][�0��;>��Ԟ2u+!��d�?g'��T:��O&��2q���>C��J�kq'P��:�d�����~?}��fQ�^�g�9~}����d�\���&�$���ܒ�z���'��'��?'��Me�a6§�T8��3ό�u�^���N2��PB>�~R?��ܞ���7�pl�T���a�&��'�>Ì�I�OӾ��I>o�J�l��h|���!����N&�)���:��XM��p8�Ԭ�ϻ��9|����}������H��M��o$O�o�봓�Y�;d���6I��'~�I����*M�<�>ed��O!l��'FS'�F{�'U�����������dq�ﵾ���Ĭ����;��dN���p��	�;��i4ɹϜ��6ɣ���c$�k�d�&�B��+'�,;�u�q���}�w\�޷�����I�,�i6�MXu<d�n�q����ט�q���}���5��OY<d�}�>v�Ԛ}�p���Mw���'X^1�߷��ߥ�?N~�_��@$���
?O�Xv�:��:�$�I��j�v�8�7��:��{y����?;C�s'Y>a5���2z��uI�x��������~JY�<��^�3GN����G��~��d�CG5��(M�IY>J��P6��6�aa8��y��$�<��a�̝a���Y'�����'�&���{���MGz��y�?oM��Oz��ﰛf�>b�a�0'P�����q�5�T�&}N0��%d�2��dߔז��'����m'���I�߾���^����{�\���߫o��/�W�+�d�9Ld�OP>��B��'�h�rC�|ɣ���$�Nj�R��<aY6�a�N2|��)�,�e�o�"��?�ү~I9����ҭ�qV��N_�Ӳќ��]�9�d�ϯ�^f^��&�k���u�6��T�.�v��8��2��PW;��@�.����Wd���*��q�r�]�p)�(�9p?�h:����]v�
s8ݦ�LN�y�����~��ﰁ����M0���IR���0���&�w&�q!��!P�'�o���ԟ�5�ē�4�$��'O�N��߸�f��~B΄�=���?���D|ΧO,6��!�x�d�R{��<d��y�I�Xs�u�c���ԜAHw�i'?%a�y�*O�<���0�d���M�轥q���߯X��}E���u�Xz�i��d���S�2u��~N�x��>�����N1}�o	>C�59�:��1<y�Y6���;��2q~	h�睐��g�e��צ����=d����I>d��%t�m6�i�'��(u���OXxÌ'�S�x�ԝI��rO��'}>ׄ���r�O'�4{��u��:k�������ӌ�%d>���~d��I�� |ɶMo_y	�����O�2i��XM=I�?g'��:Ì&�XbN �~��$��u<k��3���W����=�?�����jϙ���r�d��	��p�'Y6�����?2|�����+'�?R~k'�8�d?3:��Y�I�*x��
I�����_���ӓ�	�Lw��w�*������AI�M�f��p'ue:�N����m��s��a��'5߼�����g�%d���>Jɉ8��d?3��Ћ�������m/���_�?}���:yC��<�(u�iX�a�N%f��P:��gwd�a��:���	ߛ$��'��I���f�J�l�%wg��`��~{�f7{P"��x���̤:���Me1$�f!��I��o!�N%`k�0��u����rAd�k�;���N�I����p�ܒ~v�~���_�`��/.�'�-�>���2?y_Ұ����
�����u*Vi8���6�M�3y�s���������!�l�����|퓌�'�YYZ��j����F����Wi7v�����o��#ǀ�9X"���|8��*Y������x�r#{�-�*�1@(��$3t5� �>��?P��,�z{2��r�]��E�)�W��	P�����=��o��b�W��Ro��"��miS��f���s<�lgXĮ_v�p_f7ԭ�����~��ݯ����'�s��2M��y�T&M��*O�R,�I�N��,�i8���x�q���m��䇥��a�����7������O/�����gM��'�'o6��O{�rN�=I�����f�5���,��w�%AB{7g��%d���q�i����SL7l���=����η_~5�������4���!��&�'�����OXO�B�2i��g;�u4��M>���dѝ׀��C�Y*T����%d�+'�P6ì�|}��׍�Z����<�|�}�wzי�Jɉ�m���I�̞����q�|�L�I�I�G�xɶ��
�z��v���;;��u'���VV�u�_�o�ֿ.��{�[ﺽ�J���L��ɶM�&�,'Y6�������C���l�a��䒲�����:�9��8���{��m'�h;�!R~d��;�yԠI��~\���G�d}�C�?Q�}߇_�,�}@�e'P>a����Y8�|j��̚d����>N�z����RLeC����,����d�
Cs[��s�:l�y������~�݂�2i*��$+̛��m���_l��>�OϨ��'���hi����T�βi�z���L�a��ΰ�B�����v�{�L_>ן?���ߏ<�]�AI1;?}��M�Bo�i'?%a��a
��'����'Y57�I}��f�)4�d�?a�I������q��~Ld�$��k�?>r�����{�5��d��m�5������}è,'���:�������M�}���{�|ɶMM�>d�d���'�>d�{�'�O�a������~�3�ǻ�ڏ����?s���<��a;?~É�N��zO��>Ci:��>��N��<é�I���I�VC��ì�d��Nj������IY?0<��O�d��k����o9�n�EjJ�N^�*fF�o��{ܮ���e[B�+����i[��ckn����n�s�4��b��1�k�}�u��[0��jZ��싌U״9�eV(�JoY�ˡ�����v���&�b��v��wa;A�O�h�*;�������c�o��/�C����T?$�eO��d���:�ɠ�x�q��S����:�\���N�����M����u���~I�l�d���������]�y���u�~���+&��C���0������~�8�m
�jè)'�8�ԩ�� ��'���Bq�Xs)�l��7�ì��a<��ߧz����~7����?��Ͽ=��8���o��I�I���T�Hyl>J������x��ї'�I�����|��C�8����'Y;���H,�a�g���^{�޾u���?~3��}ݷ��Y'����xɴ�ݩ'�̛>�B�M�G<�+�<��䬟 ��ZC�:��їM��k����n�y$�+����3���{�j��;����������l�}g۲
�����8��'�� ��'�=9ܬ'l����J�m��%b�z��� ���!�N���M��9����2�y��7߼�8�0��ٟ�2o���/0=d�&��~�s |�xk�|�'��2{�p�f�=a��s܄�i�G{��V�jw̒��3t��䬛�5�}�|��\oyӞ�޷��'��'p�O�|�5C�d�Oo!�N}d=�ì����;����M�z�ԟ wVN����i;�!�$�w�d�B�������?&���tn��������@$��>�>�ʓ����'|�����3�hu�����6��:�����'�zgp��Nz�'��a���u<d������҇�S�?C:����<G߾�X�>��IR��}z���+'���d����0�@�?{f�̝d�f���M!���8�bu���=Iԓ�����Ϲ��׊g�߾�����ޜd�C��d*2~Af�9�:�̚;�2N��sܒ�a:��"ɿl2���2~|q	�C�1�O6ÿ���M!��}���\�;��r�i�*�&���Í
tݽ���mھwrE���X,kJ�Q�]�[�eǇ��\�$�;Y���`��ⳬ7L֏���~v=eѽ4�.������e���)��b�y&:��Hi"���;���n�����.uI�>�ޭ��L��yߥ���t/���L>I�P�0�'X��AC��%a���'�Ok'h7�I_Y'5>�N�`y�8��O_Ɍ<d� ݑ�*��C�����FY�(��G�I�oy��&��w�'�*��Ad��=�d�A��z��>eC�}�
O�<���I:ɽY+�I���}g߈�s�K�^'����,��x��gOߧ�4ì'����2|é?j��<d��t��C��è,'�k�0�'�=�I���P����>d����'Pʫ�]}�W�U��}��l����?]���&������gǴ4��Oo��N1@�����:����a'�:���'SL��z~�d�T&��� u����A��b��{��~���~�����?5'��&����M&�Y�I�+<���ɭ⇌�Ad�vO��'R�����I�59�N��'�~��\�5�;�?��oq���?|�?���M�o�'f��u���>��IY=`y7I��<I�T'��N�쳌&�T�T8��0����Ad׻�)8���������J�����k�����o�=I������'X{�ì�0�ÿa�N$��'���I>}�rJ�l����+'�8�d?&2q?S'�u5<��2qk����m�K�+y�u G�J����"��6ʚ=�H,�a�a�i'X{/2u��2m��ݹ$����$�	��k$�6��Z2�|�'�� ~?}?�ץ��b���s�+�O�}�=N�a�x�>o(u��XO���������� �u���~a1&�� |�'�����g̜�Yd�'�d�&��Gx~�<��?w﷽���T+'�,;l!�'ɣ$�'S�Xm<d�u���'̇����d�����>`u���m�'�O=���z�O��xT}�i�YK�����$WvZ�^��:h��͝\�A�\#�ۼ]��8�OA�t��y�5���㗩��`�^��sk��n���WA��'J�%��c^;6|�����צ.I�vT����$�=:/��F����w����_�����%ABd�gP�� ���6��6�aI6����I�~7��:��{y����?;B�β~a9��M0���� �Z�vmw���D���W�>c����_{��M2h�?x$�	�w�+'�Y*�q&����q���ՇZ�q�݆�c�'Xo|ì��w�˞�N��g�S���Po��������M$����a:�2|Ş�;�:�̚3��I�4sY%J�g��
��VO2��dߔז��'����mM��/��/ߜ^�͟R�ﾫ�u����=����p��Y'={���I���!P��4s�!�>d�}��IԜՒ�I=��d���,�d���S3\̏>ߗG��5��߾�;!�����~d���{;�H.�i���gY%J��o�u�XOS�ɤ�AHk��T8���7� �����d�$�M��ud�s��q�!�ީ]�����?7��_�������d���O_���Y8�i�?�<aԟ���3L�C߷�d�������L|;̝I����'�8��V��AD}�}�xf�W�X�b~YN���>����Mj�]$��Ϭ�_̜Ma�I��5톙8�yS�u�I8���Y�'��I?!�9�:��1<=�d�VA��L���{�����滿_��x��V>� ���&����M�j~�$��'F�'��f����u5=��0����:����!�N ���'�?c����c��9�[?a����C�ӈw��l�J�h����'��7��'̛���B~`k��O�2i���XO^��4g'��:Ì&�XbN H�G6�,����v"�g��(���d�Nk�N��9�f�O�o��'?XO{N2q���O9`z��'�d�����?5��CYd?3�N��_��ﴊ#�	z_��?Tos�h;W~�xk�2�A:n�p�&ˡ���v�/���9�2>�y�舦iYّ�EP�V�E�������6��y|$��㼭�/$���ߏ|)H�����>�^���S�v�a𾒛�v��ǡ��f�dB6����ci�f��w��%�̓Ml][ԥP�(Y7m��a�m+�7;(˚�0G%b�6ljE���mG�K�jm��ܬ� lU	��L����8oi��N_̰���k��[��Q)ۥ�:�et8�P>Ջjﴼ\ ��(Vqj��}|�eN��EV�s)P���<5�_f+2ȓs�=�Rq�V�m�fws�k�b2����po_w�*��Q�w���]���l��JĕM	2��]��=Z��Z�y$��Z��@�\jJ��M�-@6�������j���-�Q������]fa@JEV�����v^��}���r��Y�W�~�m���)�n��]*��^*4h��IŪ�96�*��%ukԥ�5���qF�z�!3:,C �@�&Wu���M�t»��ֆ��A�k���l�L�B��\�]�7Z�4�v\u˸	��n5
(Ր�[w	�W�9�OE�>n���H=�p��3E� �̹��]��e�ݣ�w���˲�U�H��G>�m��.��5���X�fҵFd0�H��(�:y+����y�oI
���P\w@����b]v���������Z����@��-H+ni:qv����w�X��C���l�_Q��mv�;%���z�U�N�	�Y�5:/�P��Y�
Qc}-��Gpwۻ:������b�\�]'�o&�*,jj	�5��Q��{g%J��ڽۺ��
�����.��wn�b�^�j�[��pB	���گiM�Q#�84�=7��}7�o*\��w�]�|�����=�')�6��"��x�iE3�R*�.�yN����g��z����*Q�O/4�ר^�h+�6m���O$ 蝀^�,TO�J.�O ����\�r]|J3�����r�MF�Z�R��ty�������/��M<�om%v�Z��4�I$�\�k�ad0�y�,��vҼ.����H�A��r����媪�;�r!�(R}�q��Ӑ3/J�m���JY�dC�� U�Sv����}x��#m�Ľ�����5��O�?����ц����jI�+w�.�*��s�@[��N.�	���"�B^M$ʸw��@Xm��(�]��y���N��y�V"�k�[ڰ��)��iwz�n3��[���ޤs1k�8b)n�=����Zec���S:R+yV�|�\�l��b"��\R��hJ���J�Y��l�;�if!���b�¼��֥+��>{����l8����v3x�\
��ۤ_5�������[����(_���82�h��U�]���p�R�9�f�T�����;�`�̈́�0t��竒N	���ǻU�i���$�~'�
H/��H�Qb��U���-�"ĭb$V#m�AX#��Uc1�����UDAF(*�F1DEX�[
��EX"�,FJ(\a�YUAQm�6�(�1DX"�,U��aZ"�(�m��*ƴQAEc-��U���,�*-��Uƪ���X��R��*���Dm�҅b����kYmm�V"�DV1Q*)D�UV�ª���AH�
�%B�Pr�Q�J���Ԫ"�VTY*��AE�j�m�b�Qj�b"�,��[Z�DJ-��b(�J��+J!VZU*TmR���(�j*�A�����D��IidPFDBQ�TF#Ej�Dcl*
3)*,X��E"���Ah��E�+�6b*��q(�(�K� �,QC)KkĮ&>�oPp�6��n�v%��Q�w�85i@����mm��.N
w̍��vS�2����=��΃3Z����I�s��?o��y�������A@��
M�q+7?sq'P�S�����:ɷ�	��s�a��O���I�I��䕓���|��Ĝg��:���bN�s9�Ÿ�����~��~q�z����RL>��q+P�xE�8����A@��N��:���:���	�w�$��$����a9g���b�Y�O�眏�hg����8���3�)��o���o�w!^c�����iG9�� ���ɕ������\Ӟ=�v�Y�,賲/������t~���{`����o"�'����ڮv>şHҝ��Dg3��8�s�ٝ�O#]��J�ŕbG��m�_(�Sz�s�\Q��g)0M�DEs:o���]�]T_���6t1��;wpY�n3ngg��n 5�E�Ȑ����:�U_�nuۘ����/;g&^[����[����e�%nFkrj��<{�;kīo\k/	��(+�Z��/I�:�n�y���e�����ʻ��ro�eOU��37��*j����y5W:�r���{a�P1�kD������;b��ӽ��{�j=�RU��#�̾�x�-�l��_X�0E�z_m�҅�Rf�|��ux�X;�c�rM���|~��_<��I�,�S.=j�̨����ᚧ�6�u�2gj�2_t@��Ƴ����:�'3��X���w�����  ������v7��?Ù��s�OF-�X�v�y���@w)�^+]��^��}�����>� �|T���s/'�q�侧�by���,�K~����M��v5� ����y�P�cj��6k��(?V�Y�%y2j���{�Ue�3b�|4-�m��;��#�)'��'�.AҁZw��>��m;���}���S�\0^��������)�����s���W��$
����\pR+|k�^�B��}z(}�8��sgy�:��A��z2W�����SG{s�=7)��Y�~[�:�6P�1�ݗxuB�*%tu���6	�����.s�	�ܾه��:tX;\�W5Uw������l���v>݂?��w�p�϶a��_s:,닜<��g�X<������S�7�~�F��D�<�p�O�km���D9W+�r�0�zmxw/T��c�F�뛠�5F���7/�QW�^���*:!���P�|{�5�G�F�A\!�`��S�(��qk��LfΈv�+B��=��뵂���ۇXC6pi{)=uX�7W-��@�䦬]��.=�U�$�SOL�������ȥ�g�ۨP�|��[�H�����{�b��x����r��2���s=�ݩ��۠���郓����f=����r ��)�Wz�ߐ�$.���l�X�FGs�]���C|5 3�N�]�l�L�������z2�A���MBe�,p�{�Ňb�`�L��_>��}��{� ��8�8�@8�3�t��ÏD^��g����o&+Օ�Q�>s�8;�=z���}�ӊ���p�1�΃o��vue��,���$QqO�f��m�\y��c���^q�2gi�緆`����Ad�c"�{�=�[�YZ��/��z�C��v�w����Q���\�e�琯�6=v���������^�
~7��������^��\E\5�uS���
��'*Q��۳�I��d��h-`�.��:�D��a�Q��i�w�bg٠�����:y�&��N�f	�vN}��vؘ!aУˊ�����n�U�J���J�++BV5�k=]��B�T���r�wN�s�I���Τ/m^�V\kv���J��i��&�`�k�H�s3��꟫���
�_��M�c���z4�E�;o�4����_W�����|+{&�-U{���+T'����AЬbX�LǳJ����6�}n�WMjb��9�8�P̽l�O&^�'6w�͕�'�A�Z#�O;y�C[��+1ƆgG���^�6,�:xX>澮v��WG�/���Sy��obz��S}fت\��E�y�5�γ	�j���U��]Od�y��(�{r��ŷ��̔k_:4��r�Տ9 $��"+�5[څ��ݳ6��z�Δ9������N�O�z�|�[Rx����5�7Sj����P>�5�]�UF��y�%����Hk��ا�&��e�'�FP��{�/x���n2�����>�n�y� r�R�@8-Us]!fZ�y=R�73=��ִ{������o�Ϸ�{\q�$zqҸ|�0���>�|KИ�/c����䦳syM:��NN��Ք�
ܓ��B�p2%u�C
�����ջ
z��A��� �-G���t����ַ��z��m��w:}l����g_l$,��	�'{���r<�^�ƛ{�<u֮�|>������/�����}�q�v*,C���.n����+��Z��S��=�ې]�;��:m���9��y5���U�{Jw�/r���_�s��2mc�@�j��ɏvy9_Mxt��m�� �,�dX�.���ϸO�����}�5�M��O۸���62A/6��q�֝k�)&r��7�t�}��w�zw���b�`��m������*%w��y�គ���7���Y����IӋ��4��+b�O&mM��|}�^P���S~|N�\�se1'���%��ؗ���$��Y��Q�ޗg��T����칕u�@�4V�|��^x��+�ꊽU��/��u?8���qp��OB'�ߜ�ֶ���ݷ//~y!�ǋoA�ϖ`��6MNs�ϦG�.��OE����<��+�|������x��jp����rU���6�_p������֝���!C��e9��GRWRJ p%�f�u��vM�.V��S���w�ynoS��s�)_Eq-�Ց���ϴֆ�q�il�����Mv��i�
�����m�Et�������}U_}][36������W�����s]�7��|�E�>�����(M[~��<�z������FS�slc4/�^{���Q���/�'���7�N�݊y��ؑ5�3��-}oo����tM�� 2��[OE;���=���՗kR�/���Gܪ���י�3x��@]��7	S^���CBk�'Wxd���b�:�m�Q;R�:;�a���})fp�5͹��T�+�cӟF}~^���"����������+N'=�po�g�G:�����{N
f�H��qb/����x��k���;�X]�^�ڥ��/`�2�I;Z�I��q�������ٯrV#]{���O�/��ßjq;�	ӽ��?7����6d����8��}H��N�.*�6
�,��^np6/t����t�]픩�A�V�WD������3yXKD����oUd��X�U��{ϧm��#��.����}'9����u�6v��$����#��q^�B}9Ʒ�v2�os�SA��c�gz���۝�Mh**���(�P�����e?h�Ad����������)��Ӭ��^���oBj���q-Ҭ��{�����Ѱt����8��ٜ�=`��`�d��=5����:c�=I��W�D��s�7�8_lG���t	�5^�9��W<�{��إ�;݃�q��o8p��:g�o�ibYN�Ig��6�;���#�t>pP�k���:n [��Ny}3}2-W�V�MxX�8s��S}��DVæ���^�B�.���y�٪�/!y?W����/���P���
d������ս�����U&jj�pSF{i��yd�`~��!����C�OEQ���Ѫ����/�>�Vܜ`I���z�Oo$=���% �a8����j���0�\ӡ��^`ش���Mn@/}a(���8�,=��9�1���o�x��H����7H�n1=����� y�r���=+ ����_i�E=�{[H����l��\6�e�d�7Hʅ��,$L��%Ր��u�N�������'�4&��h�HZD�n�n��.��:�1Ԫ闵��u��n����|>wj�)�_��}�p��+��t�|=�L`�؟Ax�x�c�ޏ	�E27��׾E=F�ڡ�w�^�;2�=�y�+֤�oqFm��O����ޔ3��H�T�}I^v��`�{鎄�c���̍�X;]/^7�C��(���}���N�)�_L9}�m}^����Z>v����	T������x'�wG9܈A�O{�ž~w���go,�ҧ>v��}佭�׽�/Er�s�g��|�@�{S�{>�w*87K�o��/z����;%�iP��*�B��l�9=�A-I����zvU���{�,/[9��vF����g�a�`승�������=�Oټ���zZ5�Nm��[����u�xY#�pqވP�`.k�f�^?p�9���D����'l>S����j=Y3�O�DP��@V�����~㻐.׃Swn_�}ǩ��nP2't��������^�ߗe�m@@�U'5cV�)�IJ0���z7�?s����Ũ>r��:�P�lU�:�����RSo� �L��;�޽�+iQ�X�(�Â�Ӓhv�p�Fr�Y��eΚ�%�rXö�>�����FR��vw�8Iy�ȷ>�4��:5�7Shtz�8k��w%��lo*vꟷ������Hk��أ�w,��1g�$�S9���h^����tE����9lO\4�Ԓ0�o7�s ]Fo�nwzI�fz9���W����7��*���q�jW�E�y�͖��ۤg�r�ܯ���z��=�u�9��y=�m�������YS���*�ǘ�=��ǧ>�lz�9�;<���meF�߽hvK���'�|�(枙���y���y�W�1���y��kώ�������=R��d�SyN�%J�[&�58���o��2���(���'�ǭg��AG�Z�>��s�|<�u.i���$ys����8�Nv;p��}6x����7����+]�^�pl����t<6+���V����/\<��G����_:�\u���՛���M�ڣ����#o���$3��F%j�*�{��L��h�G`܀�����:d�9D��$f'7)����Q�p&�u�o{���1;�q�⤊=V8OL+1���*>���3 �U���}[^M9����4��||�m�;=s�se}�$���[���v=���� �5#����O������G������/���?�F�ҳ�Vi��Nz�vx�wdð�w�f�`s���ԩ��>��P�9茴|f�s���_�I5Z������O�k��5qNJ	����DG3��4(��>��ii��ɖr��=B���ף���o;�%�I��gǥ��h$�t�����T�u�t�?[�q{{�K��^�R[�kv{� Ѿ�9����dh����n�?\�~����}���D��G����hp�;^�W=0ӱ=�|��wmv�D��ʣM�ү3�(��TŢh\/e��d)��n���a8�g����W/	�+\~}oz����qE��9��W�������s����3�_��^�� $E"qKt9��Ԙ��	{�u��;�mFo����8Y:�K�Cu/��y��L,�B>�����L��:�i�1YkE�rf��mIf0/b�mGN���M�E�s7>�d���\V�C-�W�7I���UAY2��&���3P��uքu� K�6T����(�\���w�V����Y͵)�i��ܺ��X��Gj㽔MdJ��s���hTN˺�Q"��eŋ��g�kyRX�_:�[wy[��W:4m����1���*���,R�q�U�pyQu^��[g����N����9[�K `R&5��A���^���97o��'�Ӛ���b�m,��f�|"@)uj�X�#��SX���2�:�>��%ͽʳ]�w������D�t�c���tek��5�j�12��X���=j�+8�S]��H=Z�����t�|$7:�c|S�W*��8�2���B���^�K�޴��$�N���PӷI�۬�g�K��䢒�ӈV
m2y^n<gq����CW�j�_H��v �]�|�$ⶳ�q���Y湃>N��Wٝ���SJֲ۝.V�@+��zN+��^�F�ݺA�!]�R�c�H�-.���e���';3T���m`T�SY}|{��ȱإ2�tm�ęh��D�ھǹ�;����{
;��\JLv��,!6S���kj�ҁ"rS��-����t)�7u<����`�r���{��.f.�1��ۯ`ߘ�2���q��3���զ��6H�c10&�7�f�I:�k����lI��|�\O���;&����g5�f*�&�^r���엿,���8]����1OLZ6!R��b����/�T�e�.�5�7����(J=��F��ث3������G�ξ쉪��w.^<�H{�^s���$�����[��N_4��ӍL�|9�):��h�����33z���M�� ��M�}�]@#=-�Vd��=J�w7`��:�B����y�{+Zz�{z�˗S�r�m�5hJ�0�:�9ɝ���j'�t]8��5x��@;D��cp1��YթMX������.��7�5�6hqH��{�/x��1�-۵JaY�����ʒ�����J^'R1C.XF^�����,9)��$Y����=$��^Յi�9�7Y�:Ă�*��l1�Wl�o]𐎫z9pп��^�q �@��T\��ȥ,9]qێ��u�ڞf
hN�HWmd����J�j,�V%�'c}Ǯ��*�(�t(G-�:�ovCc-��\��!�+7��B�[X ԥ3L�7en�YC�NǨ�_r�<�rw��ӫs�]��:���9�.ŧpE����Ȼ�gix�.�5s��*g<��V� �����鴁{��w�J�Hq��Wr��n]�U�[Ȳ�nwn yofw ���u0�N���E9�WG$�W5��� 4��n�_]�\�2��9$�3xZ��z4�)-��_y��{EQ`�R[j(E ��F��Ơ�%D����
@c
�!+��-�X�!Z�J�I*"��ATơAUE���V	l
�I1�%��m%A�Q%V
#"*��PRXJʁV�#[��"(�*V1kQJ�؈)EaX*�U��Yr���Z�������ʑT#"�`TYR�J��,E��E��2Q"��
(�*�-"�QQ�Kh�*�Kj0��-a1*��f!R�e�YY(��iZ�*��
ČE�J#Yb�-
�����mAm�����Q�m(�JZ�̂�ikKj�Q�KV�Q�1L(_~���އ���lfֺ<~���nkj#z��^���&��d�GT�������^�|�P�Y��ޱ:t�邊�]���W�_}^���s��-E��=�����j���87�3�&v��Oj��	kiW�j����X����d��_˵1�yl�>���/`�3�M�ٹ���:m��Of7��1e�ӝ~�����.�N �&{�k�x���^�5��η'F��I�)z)����M�¯C������AL�кM�y�^o��o{pI�pR=�ZN�)��S;k����X=�
�M�����|�A/���q�!�94zΝ�O|h*2�����J�pW��S�W��}�K
q������Z��;'��<���Ŭ&,��/h���S�}�2���M�<�>y[�<^�Κ%j�Q~��t^)��ӊ��z��
�͗��5}��S��0�Z�B���v�yi@7.���DP�t���{aB�wV�sΒE-c#qW^ɝ�&�̿k���9�7YW|��{"@����{o���^�62�\P�y�	��M6o��LP�k4�97E]`{��Y,�X���i�d�i���U�WQ�*R�T�fH���+ٸ�v�{i���v��]v�R�oW/�}_U}�O�}���K���G��~��������dSW��GP�`G}��v*��Vxs�
�D��x{ӽCvk�Ndy�2ڐ������=�v�����Z��R�ϸ���soS�;���7�nJN&p?!w]��Z��G��S����O�t�'+�U�$��z���^�9�N|:K2w>>�Ҽ�=�/�Z���T��b�y#Ͻ�Lf���s�&8�M>��D�����a�6Q^e�F�>�wj�/o�fǞk_�E���xD��1� �-��e7�t������e���ah���K���:x�M�k��A�ƶN�rM���D�y�]�=O���zO��<�g��Z��g2�7I��vg�7��ٹXhv�r���a�-
x��gj�G�@:���ew\��Ns�|\jx�!&w�>�"r�;*h�轆^���xЛ+�BR;_�YDv�z��*��@\㬹�by�ߑr��;��X�5�	��3�8*\6�;w��ͮ��-uiŋ���rx/���C�bj�,Ɉދk��@���N�[�xyJ�W�}U����{����(3���!U�\�<��9=��XRi������q�9\)��`��1�������E�p��˯���4�v�M�Fd/�^�Vo{W
��J5�W;b��l�d�7�����;.��˫"E�赑����^������9�Ź"b"���U���G�Z�{��Vut�$�����5������[^�"ܹ5
�4 �p���*{
���c7��4��[������'}"�J���9=�#H���ɗ��k/	����^ߕ�x7DH�M�9l!!�~��c4�+׃T̚'�^�S����CWOs���,y���^�E���j0���򒎵�E�F.����=
�j���Z=_�-�9��y1��c&u>��2��e�=��U���|�=8#���!�q���9jހ!T47�k�z%��1�kMq��{E9F���WRn�e�1�%F���u�j���a�we{�����L�/�MV�s��vg��M����K�ő�����QA��[��u>��R ^:/1n;Ԇ��$��%[oP	϶�m"V�����p��?>��>�|ƅ3jH�#v��x�������W�1�{כZ�G�3�Ǔ����r�G�#^�wvW���v�6�u/ �I=�Y��U�9��"�ʗ*�}��pp/x?��F<3�+���0��c�= VR�9�x�Z�h���:�U��|��ڠ�m2P�T���R^�gd��ϐ��'��!�Ǥ���q�zW�s��>>�+o���k�)�3�-��m�tES3�l�8ƍ�{�9�_�q�!� ��N�Ps����wᷩ��Nѳ0���
s���G�����y=�s=��}>�κ#�������~/�wnSN7��m��}����|z>6�8V��:��&���b��v�ٷ������]*��\7L�G�*犳ا�W�k�����r����s*�Th^���s����q���=�F�ˣ�H[�Z��<�������Ы� �&g���h�X}�u0����yqaV�ޡ��v�o�2���f��^!d�,��}\ݝp��Vq��Wҳg��j�࢓j��cy�g�S}u<��!(����F��b�.�Jc�}���S���}Y���G�%i�S�m]f���Z�$�gHS�m<�U���꯾�]������������*����G�^�ja��kWd$n:�V�aǸwJa�uYѕ{DΆ���%���^�s�������9).���n�f���P��ՋT}��I�S�$5�Wh�*
p[ڬ�Q�)"���ޣ3	e!�P���{զ"߼Y���&-���C>ވuS�,^8��2���#�<3���� �W4u���� �ܲN��n�a�Uš���=�!���S��Y^O��U9o��#>�N�HW+ޣ�t���O՜]�,x+�|V��7��D��+Jtp{�(�������5�p�ΓZd9�l,�x2A�R6K񔍊l�*��O)xu;���1jh����|f�\l��v���2H��ђ����®R��u��c���j��/���s�;���Դi����4���S
z��:�T�dp�bHy����})�t��m�{�_a�N|_��9c�N`g�g����Nh�z�ѺЫ��vΐ $$^�Qgh^���=����]��)��ŧ��y9^N���E@��b�CF�i�l���Ѝ��â�������,]+��5]{����f�{"���v�WFA��޶Щ9�5�%_u��a�䶒�i����k� �w���y�瘕6��s9�,1�{�������v�瓭��yW��"/�Wq�<rT���2����,�k3�e#Z68މm��߄Ĩ���߶�њ���e�f,i�9P���l3�oڰ�����G��}L�c�o�Aӏ��T�H�Ҡ_ܢZO(f�>���2�l(�=1��K�ؿO{�7�yV����=�����4K��ǃ�]uʅ
?g��w�b\5��|'rZk���G��ܩ��_w������U�K�| ��.#�)�Y$g%�#�^���`���K�J�[���]i�wY�ؔ�cJO��RZ����9!�td��1#�t@۠U��=Y�>�o�tYX�|��/֋�֡���).K�38��s�*bPxW7^����n��'�/���!b�
��S�v`~��U�Ϥ�����j 9�kf-�-����,MVQ��.�W�����u��\F�bol@E$�\^�q�W��IWg���Hu�
���j��^?5��{��N{kN��ǎ���n���z;���q۠L�Y�U���H+�j�wo(W<O�z�;�w��.)*�@��"�VNu�����%{�U��ӂj��R��*�̇�r�<b���D�UoV�x)b�O%1���%�vΜ0bju
ŝ�X�3C��t`��'U�G1������h���[�6���)�#��t"}~U�w��鲰J�	��x3�^�C���xm�� >=Ⱥ�����<����2���?�"�o�C}J1lg��x9]�ޑT�}���|�.�[D��,ZbƂ�lʕ��Rj(s�'����L�xd�ܼ(k=�/z֨�9�����{���[.�WV]�3���	9�Kf��̠�X����i�0�51e{��r�O��Z5���YTNUiB��tk��/>���9���`��f)5Ն��?oT���p��!�Y�=����C�24��h6�����(o�qM�T�x��މ�0_VǷL������9�39�8冩l��#B�t9�ҕ*�:�G2���f�j�Ǯ����kRC�-�|�y!|�?xzdO�&[+�z��	�ɱ� V�a$�y.��������mV���n��m��Q҅E}���x����ڸ� U�#�[�u�U����r}��.�k(�ڛMm�O�*W�d�����*�3��]Vh֭�\7���E�Ɔ���MQ���c ˎ�ȗ���j�����ob�F�=n�ZcM�/��@^��h�� VȮ���4W���'�6��7��:N� n]\�R1�dr��E�M��q��;\8��D#��\U�����9F�}�W�}��II�C��N�Q8 ��/�"�����G%?n�+w5UI�0��Π��]�CB�.�w����$VP���,���׶"?�?�t��^]7\V�ٕ%v�Vj���t��M����J3�����D���*;���0w�z����XO���[E�l�yŜ��50�|��]���㧓�����9�Oj���Z�^U�Z��p�	�,���DS���bN�|�U1�cқ�t�<�uX=<�����ui�{<�jh�Y|�V�Ǩ�{�ae�KLR�g˵d�n_݇+���}RS�Y"�������j�Ѿ���I��!��V��ʮ�5��+�IG鄖5[3Q`� ��к�~�Vv��R\�Z.����"���`�ţl�.z�����ܪ9�.J��P��o�b�y�б<�h������~��fS2��P�i�����thl�J��]VmO��uG�M�^C�L�{/�K�ͻ��J��s�Č޺ϺyQy������W��Dsr�yҥw��\k*���"���X�L=F�V��P0�1݃OOv���߮�������Cbuӌv�+����;�-}�M���8V�w��oN�|ɰ�P��[��>k��W=�I�T(MyG+:庑���L4�/�s�;N��٧�v�G.� >��sW�I�H����X6��7�0�W�9೟L��_�6�銋<Fɷ.�����6��\�e֝3�8�U�'aU�Ø����ӣ�g]5\H쬓J��~�*{����3�c{�V���rTߌ�@�&���yxޯ}|���B�_��F�b���s�Ķf�:���P_�殁�Tv���-bP��K����W�r��}s,�3Uu�'hj��"��?#�9V����"^���Y��7K��9M�k���\%n!�]��P�4��ެ��\���ߪ�+�`��N�����X�W��W�	��RO�V$ȋ�/�Q��˦��vz��;����ך���g�a�9�_ޔ��Q���&�g��ᚐ/���r��	.l!��������?KT�}��0p̦v�G�t�75C�5�f�Xj�%6�v9HU��a�o����l��R�n_�@{��>��9���\ �Or��`�>�59���lz�[�+-b5��-����WYZS��{�(��Ŧg�$F��%�UZ�ue�U�ѳa�)��jU���^���;�Ef�\�1�ƄQ��e��H�{ɒ<]����A�֪��׎fLg�]����K�k�hV��]0jP�=�VΈ�H��+�y'��־����s���k7�5ʮ=��!(f�wf��;-v��������= t�%sDWN����5٦�k�����}�-z��T��(L����`�yH���Ƽ{oR>�6����Q���p�l��]y[[HPQ�H@G��ژ�˙�ol�GS�)q�>,[�0o��A��)��cMi�v�'�!�^*,�\o��ۨ7�5P�eޕ3�>�~W�<(�4��x�}bS�3������N����Ѿ�|2A�y$�s��f�d��<��,�P>�$�y+o寸E��6���2�G�g>���zP�4���V�kxż����x��<�m!R��ǌ�@�Ƒym��s��t���>Ŕ3���:�{�\Wv�.3!���lD�o��/�KA��8e�>���124�����}�Ά�%Ow�Zj؅{޼Nq-	ǜ��]
�.�
5[ԫ�.AC�o�x�>�&�u�K��3��є��Bkhk�L���a�Qj���y�E��q�.W!����9j|�{\�w����*�n�⟬�f�B̔��$��$6���!�&$aϟ�����f�Q*k��/�v�2H�!��i��r��|B�7�|�Ji=����P�؉�2S��������m�v�fw�]�
�q�Lɺ�GK9@N�T�}��}՛�Ѝ�蘺��Ցv�˳��Rs����A�A�*rJܛ�8@�ǀ�0!s*��=u�e�iC�co,����Bl|i����hE�.�n^R
�60�JԹAwU��7�ʱ�NÌ�MɲF���F�y)�Y�o���۷�J�:�u�U�ng+$9�d�ᓓ]�o��k��l����6>��e�+t�=P�V� u+�XW�͡Ρ%����w��l<Zr�LV y>��!���'jWe��5;4'��1�V_R��t�\)��rԭV0Ωf�P���hl�.�_d眷.��x���r>"�m*��IFg֏+lh�1<�53K.���V��,�k�R�a��$��/������^�;�I2�""rr�!�m�}�4	)�ڤh1N��ZS)*��˝�õ�f��ȲR�Ň�	���E��]l�%Y������.�ou�����/��,:^ē�s_$�ma��\���z��Fs��Q�Vv� W�),�TmՓ��-�E!�K6��O�,�T���r�F��������WnlX�i�}3�)�Mi�|~�0+��(GG+%f�7�j��Rmoi�xyM�v�>�57����YEJz�ƶ��6�P�}!�#pN�W�0���MA�v�G��oN*�iӗڹ��>z�2(�|�)/�t���r��{��5NC��-�{���Qh4��ށ��˹[����_L����p�׳�SΧ���ۥ��J��(�2[H��s�:w���d,u�6H���ڗ;�Ε�@���Wh��k���%^^+�4z[��f��\��,IQ7'S�z�/�%MA��|�*OOݮ�7��<1mm�ՠ�o:K�p�o��v��g4@a��:Q(���qJ��6M�9�h�����o���Y����rM,X.��V�K��F�KC�)0
�i�L�Wm=f�T��P\ؾM��۩s}m�Yv�A%����aI>��U'_n������2���O�Z+���C�Ei�}����וwt��X�DR��gt�}B-��q۳n���#�>�#p��d<�ou�5d/.��a���H2���#��SFJ�xW���U�7ˑ��]�y�-��}�����.k�u/��\�h�x���;�`V�[;�/��4�w5��8���;�s�-o�,,�F��T��o�.k7�6��S� 2PG`�c��֒�A�7v;���XC�w��*�Zׄ�p�s=�|���7�^<�Ӿ�82M�Iӫ�v��U�����qG���?�������D7�9}[��y�!����k/��P1t��N-���W
p;Q!ð�B�k2��F��r��Q;}R�ڑ���܈�٣;�N�A�wÐ�p�s)>����!.��C��`X��14��Փ����X��F�Z��V��
��j�Q��&ZfQq��mQˎ1r�R�+j��lZ��
�6�S2�*�+ �R��FJ[%B�J�4Q��Z�!ET�TKebZ�E�Bڤk[cj�J�hQQE-����b�@�U��mR�+V��,����6�U��*�UaR(�ڊ�eE��,�A��YV*�*��Z��U��[e,+�U������JfY\[EA�2��U�am*Ѷ�-�j��%b���T���F��b��bZ+KbU�afZR�,-��T`��QF�[h4)J�)B�Km�[m�YX�5r�-�Զ6,�ADˈ����EKQRՅ@X�lh�!�H��UX���*��+hڒ�.a��@J�3�����mia(Z��՜��X(���֫��2���
�z�������(���]���J^ָfs�Ko����o?E$�S#�_�^=��*f�ya~֌�ϻ�
�@9p�q&�,��%�Voԭ������I�_�K����eˆ}���lj�poEuO��z$A��5�^�j�{�6�9�[ګ����4�K��Z6}�	���q1�S��j�i��j�S�7Q��Ǉj��+r4i�<���w-$��x������g*�����R����>G8֏Y��s�����g{��\�;i��W��r��4��E�^[M�=���i���;?fIY��Y���Mz�û�G���$�" �I���c�fcJei�^פ�iv�U�<�+uM�m�Ry�Ⱦ���v�S*]�BT�N�6���q�o�t=q(tu������`�m�NZ����S^���X�Yê��2N��L�j�%gY-�ϼ��@��&�wK�X�M���-��6;*}Վ��vU�Z��X|��W�ّ���;���vy��N��ޣ����HEΰ�a��/ܬzb�-28��KA���/[O���3������ǹg����f��Q�>����Ú�|{k8]��o�j�#��R%�$V%D�;��zn��/i��It3��~���<r�|�{k^�d��n�9Q�WRM���]�XB�mꕴ%ѩR�nq���%ɕ:.����H)�5�\}S�}��}���>]<������d��s�#3�ÎXj��*<�@��u.��!�g�)���y]_o��ο�ẓA��ޛ��u�e:�8$c A�D,޲ ��V�NW��q�[S����B���򦜖ع.���L���}��>N�P ��� �v�u*/,|c���G�-%��.�!������fm�\�2`~fS��/�)��u{q�X���{���[I0;��ߟ҇�7�;�ڏV����A�0����w���z�cF�@��#��ݟR�<H>˪�3��>��yh��n�&]�����:]#^�Ү��w����i�*�z�A���<[�t|�IB;����Bg��^��p��S���P���s�߻����.o#,݄�򶏟Ǹ�9�nJ1��B��:���j���g+�LL'=��R(к��d[7m�'Ƿ֝	�jB*�PyX��@t��u\=<��<t�񅎐umh����{ך��|�&a~K�	N�q�P��A��r�ć���O$P�*Y�7�����oJͱq;��|�9�
H����nBѕ���NT����\'u�	q1�Vr�C*�R�Ñ��u�����$�^RJ���p��;��W�
�S֟Ā��Y2��O
[坫�)y���:�A��.�`H˝� �m�0DV��K���nT��7E�������!��s'�mc��TҼ�7!�V�V��h�\.J9��Nj�f|�X'��=���@9M���g�58��$Cp^*�_�[�u�S ����-����V{�C�΄4�<K��I����O|D{0@�?X�k6��̦f^*��!�9�M1�o����M��{�&ͷ��ʨ<ų��L_�i�*{�r��^�`w���mt./���3)W��2��اt���-Hns+�Ϋ�|��
+��}���E���8���ch3����l�{EU#��A4��B.�LP(�)����,=��R��V��������}=��"�=��e4�5�%��W&
:6z���w�Zd+�~�@�#��=&��*�/����@�r#Ik��8߆�T'�Q��o3`�ȍ��|���e>��4xp�]	����x��X��R�|b��<��6�-1}�������	�ڰ���j��S*�ZtJ�Coh��:����^u[Kl�{N5c��V��6�U��(e�l�����{ݐ�rS���v$��rVP����}��hF��ޫ�%��<���?=�l�wo|��k��m�t�ڀՅ�
��T�����6��d��ڈT�(�w8�Z���uy��Xv�ь�F-}j=)���_W������H3g�s=�Yڵc�l�#3z`��Q՞�`����j��H�eu���vVv���#�|{"��D���.�ά�����J�T=���v�b��a�L�`�(雺��3=��#�^۞�b��>��!�F�3�_�&�瑔7�H��!�<�:��D��7�`���,�l2� =mz��l���U����W3ؙ_eiN�{�(�v-3��eq�~�[����bs!��CC>�c�W�~�ׂUa�_��G6xU�M�����E���!�&�Rʬ�~��wM��b��jf�h=��.v��p�}x���
�ϩf��Z]�˶vn�2����Ҵ(���s�_X5c��P󸇎|&���~ݐ���TYU����1z��
�^:��Θ�&\�7LQ�5��>�)��i���jh4�����pI�B�eE�[����^��^j#@�y$��i�:�ꐫ0ߌ��"��(p��4���_��vTw�y4�D�ƕu!N��@�+,S1i��~���'6�å�oX�7gJ�%f ����Wh�[��emb}>�1kV/��*��g�%��x2��}V��3DV�����k�z c�T��W��W��Ŧ'��P܉�����O��F��\P04M�Ϩ��p���uo������m��c���d���W��}^;�N��:xXO����:�P��p�d�.�.��������Yn� ��{d�b�C���wl>��;�vU�-
�޴<"��j<�TX�|���$z.AC�뗯����틚��Tj��g�����C_�fx��w2����LP�	�K"�!}�����4���Js�b���C��봻��C�gk3����K�A����GF},C�LH���Y�Pݶ躻��K�&��w��a|0f�H�_7z������d�{���LYAN�%�H�ޏ�ߑ,�bk��*����r��(�C3V�6ƪ� ފ�Ab�� ����w��j��n�$�fue[CPDʝcNW�Y�r%��oǮ�68:�q����x	�������R#�L���a6�ɒBb�G{՟�Bg�|͟	U���Kδ?�|r)^�b��{z� �o3Tj�R��A��ᛊ�S����g���_Oc�a����6��IX
��T{��XIMw�s:��*�Bi���eA�|d�4�V�a~�="��r�l�*�`��d:[��?uҮ/�8��R���B/gYYK޹{Gju�a�F��TL�_n��U���Ջ7�h�t������ko&�ƃ(<��z��
p�c�,��4��/������wYbL1p�kk�[Y�wv�JR�sE�w$�����5�t��}T> {�%��b�,��.�W`p�R�,Z�a��β�Vd9K�d>q=�!���E9�p��\���U��Uhb�qz|��RKG��S�^ :��l�yٔ���A��u��P'���2o�^_��3�ᨄ��KRؗ&f�W��Q"�[RU�`�=U%�w٣^���0읃{g��ԏ��V�HB��(��N�y�5�qn����N䜸csi���;��g����ޤg����=,5Kg��Ҡ~dh9�W:���lZ����ko��X�5j�4��WA��ޛ��G3�N��	|c B�&MʡYƇ1Z<7{�ze훢O�i{�Y]�^W���	�J_f�R�Vܹ�����
�����ƽ������t��\+Qb�d�Uז�>��X.d���3ޙ�s4o����{�r7o��Q�+t��WEd��ds)yh��.�����`��I�}~���V�g�^vV��g`:��.��.P��u��I�����'�Dī�
5�n�^��܃������Pp',֊EfW���qŸY��;c�N���e��hw gP��J#����ګn������)7{�E��0��]�c�-\��]�"e��շX����T�JtQ�j�z2BE����]�����K��:w}����f�����G���d��\��n�ٯϦe��p[$��[���BƥcCk;(�1ң:�[;���������Vь�:}ے��Ӱ������U�Ǖ�a�u��F�[�_6�{���>����`�E��Y�ܦ<7�X@t�8�W�[;��ǐ�u���g��&_�{��l�՗xx�e��a.����v���E��R���]�&��{À�8��ut1��yⵌN>���m�aU�-x�g)r�q�7¤�ǚ�	9��f1�r�ό��V�c��xt��ީ��%=�%�pQ�_°R�E��\�P_=��$�]���l��9vB{/�$�����`��{cӍ��ELμU��6Du�B���򤆚wN�ڇ��$�v6����-��fȆ�pS�;N{��2����$G:еg�SY㇋�&j��r��Y	�s;2���Ī�����	�d��L��_�e���GX�ά��{sDE�/Ӟ�~84�DA� �AsB.�LZyյ���
Ы�u�����L���됯We4�W)��i����Z�Py1 ��_
����b�>��M�\7�z�}iX�Z��"�Lg�k���Y����=�zqA��Sn����|�n�=O�&S��uǵ��ڒ�o	Sm-.9IVL-��U��'��7�ԫ�������*~>�~��RC�G{���W{k3�:�Ȱ��hW�e�9���/��jέ񁋣M��C�_��p�=Md"��t^�/]:��Fh-�F��r����yW}�&ẉĥ���<��zh��c�ǼbL��A�&\!	��_<UT,k7�H[�1`J�����gh�ѵ�n�Er����yx7b�3�P�V�{D��K�!h��p��d?v��'~�#����]�U��1yc�|������}�՜�`�෵Y�j����mܟ%���'����� F�������^�>���d"��S����9�3�l��h��v���M|�*_���C1[��em�_/���U<�VjP��ܨ���@��P�>�X��5�w��zLP@+�+t��Z�Y�c�w��T�pC����ĄS�w�vfF3�(�����#}��5�9"�1�nx/����Y��3y����`� ij:o
\���K���꩸����;�hg�Q��K�r�"���?]����(�6�Ժr� X,ZW�Cs���Uٸ=qC~U댶�����E��"(0��ND
W�E=�PԻҩ�1�F�l��q�����󶱃$���f��,L�M���!�HYbv�й�l�V1�\%kŨ����==r�S{�}��g�����{�_+�W��U���������ҝP��0�Zz#����ŇE���3��N���_qǥ]�:���
ϯ��F�"c��Pu:�._:M���b$:|iK��9�P-�:C��I_�쎮��h,䩵��2�>Vr�6$��X6���v�Q�˥�A���Z�H��y[
\l����)u<�XYg�S�wT�����m�z��ᖰ��[�H��U X��k��a����p�uxW-�潃a~6zJ~�")�z��ȴ!7�KBq�"���"!,GC[U��ur���\��]-G<��;��0%��nAG���|�I�c�#����.��P�un2o�;G�zy����Ӹ�	ԇ��+�������Y����Ğׄ��тX�z����^d�W�7�7�ܘ�밈T8V����4��c���y�B���"������om#W���2.�h^��v���FU��	��Z���^�p��E�cUC��]P�wҖ�|'�&L�y��3UM^�,����+y�`N�	�ue�2������}��"8�9��f��e��� �lU�R�f6���i5D>�[:�\^Wn��J�X�J/Lھ-�ͯ��/fn�$N�i��M�o�_zxj��ǞXOQ���r��� �	~�ٽ�g������q�;�yws��[`?k��C�x*d��I(�ї����W��[ɺ.���L&��P��������q�^?5�Y��#�R��e��w ��
��ӄ~��}��&���J��~#�6ݮ�h��ym6�;�i٪n�o�b�{��l�(4�g�9a�ʕ~ʅ]h��w��eA�n&f4�V�P������f�!25Z��/:wd�!�\�υު�v�� 2��a��EԮ��RjfC�:�{[��:�QYs�����}�b(l��\+"���g�%��I_�"o���%gY-��;2�*Ww�\U���_�SK��Ǡ=���'�>�k�%CJ'	�2��:"�t~lq됐�����R�#��zg��յ�eV���'`��KՇ�s�~�VG�KA���z�|a���g�ԕ�n�yx�O�|��|)J��&|������^x���T{J����ŧ�U�m��)�y}[JX�ܱEL嶦љp��Q!|�?y��V9���L3�,F�{�8h�I�ʳ���W�����#D�٠i@.���;(є�1.Y��3����_4��٨�\j�7o<r�����Q�.�>�Z��n�<ԖR�p%�7����]u�X^����\����B@�E���=�MnY�bS�uy�H2�v�ЇZ	N6mIF�@Ҕ�i��N��V����o���u�qLv�5��uZ�coO���q\^5\Q�}8�8l�+�]��oW,ٔi;��2� Wt�̀���ue ���I��VX�B��4\��IT��͔�57�w�{\KnE�V�{3}��惃�S}x{)����sN4��F��ә�ޙśv�
�2hј>��gv�5����w%�ԣ���̬W�w¶nP��H�j�TA���$����j�]���B�(L���Z��W�W�ˆ_sG%��:���.}���m7/��,ch�Ӭ6�,�1�0�vugu�-�B�&L��4�`$��Oo@xiGIK���3��f��aڥ���5��*C!��a�wZ�ɲ��q] �Ʉf�'W�V�T��Z��@�M���w%�j�Av�8�{��E�M.�rc�kn��Ǻ������ΖJ�Z��wzݴ5p}��1І�lRF�������ĭ�{��SI�H��.MΡ]p�!*�;g��9C,�\�SCj�����I��8��T�[w�
@��鞼�(:|�dRV�ޕ�x-7��Jr��Z���\���9�/7Hax�<�G����\�5��j����Õ8U�kD������9�RC]C�k0�V*^d^��Q��=s�">�`�� �R|�y��ݑX��B��3�v�L��]�L[��|�Z��,�����ٕl�m+C�k�IvY5�yr���S��,B��_j��sj��z�k[�� �t�Ί�����AO��w�V��8bE\�S�*����B��p1��^�zM�<;�ޅh)v&�K����!�rYw,��,jo�#�K�Q;`��>C'n�s{�i��o ]4>L�r&�G+�hM�Q�v��s���X��9�m��֨gd��V�l~oK�}s�e$�7�2���%���q�F��.�W�t�9ܚ�w�&N�,�]^q}���C��yqP�T;)hsJuu1ul���ǵ�un�w]8���)H�Vj��M�d�F���	�L��/:Q{�/K}{�M�k��ø%{Iw�s�8��Y�'
���U��CոE�;��Ts098�T�=Ṷy0��VrL�v��I��.��r��0w���p��K�A6�I�aUgEL<;x^�Ņ���ʙ��^�<�����Uz^fv��"���$Q�,:������=W�
*��)�G�)_h݀�D��x:V�� +Sy!�.cVv�Y�8�:��x�E6�886�2����6G�2r��vDsAY��`��Y�w��E|^��a�Z��r�ټ�I8�  �~I�0]��ʖ���m��q��Z*��P�X-eDj��l*%m��R�T�b\���Z1��T��`�FR�Um��E�%�&4�`��kTTţ�+D�D�W�(V֕�mRV%-R�a,H�R�Uh�U*�cRd�U��Q�A��������(��T`�VF��d���D��J�ڬ����VV[ina�J���ej�k%EU�XV��`�#A�����$�������6�Z�l�����E�Z�U����F�eUjV+
�*Qq�r�ZZ
Q�4��TZ�2�����KJ���1mZ��e*�\L�[mcj�h��
1AER��\�\R�m���[m��m��5��h������JZ
[f&8��j0m؊�b���H���Tme�("�B��l���
�ѩP�V�
[J���j����]�-Қ�"�l�Jpu(eq��`�{�1�|���@k/��"���3���luC1�[�#al�6������I���?w��f����,����_%+庭t���JLֱ�X����|�W�C鈮�6�k�;Vl�c�,��s��|����Z��\v��v�6�.V\Ɂ�e�8�K����f�4�a�vʯ�:��<.�+$��#�Ur�U��Y���pQo`;/�^˘Ur~��{��4 V���-&ItG�NY�'��uT�2�����A��ѱ��kHU콷�gܽxa�]kz6W	޲Y���O	>���6�bЅq��N�:��7�Tw���υ��~zX��g��q�'����}WcND!��a��@$������L~S�9H_R�^9*�C����epxq����<gP�����o�p�X��#��S�a�K\�ɞwN՛6�Ԋ�b_�^>K�痃��z��Z+�>��q��7�ECc<;�X�7����6U:D��y��/�`ͣb�*�6Z�IX�'�M'd��rQ�5�L���IpNw�.ֹ�����.5�����ץ	)��:��f
�K��gҗ=�P��,�,�a���,�n�����R[����a[0v�*駮}�����Y��C����H$���]Ͻr�k���!}���;ۅm�����9���@�\;���m�oi�Y��[�i)he��X��g�!3��Į'3zT�]���'N�[&��Ǘ��ﷅ�U��B��'���Ǿ����fg׊���6DuӮ-8U��ҳf-mߕ����Aҋ=U��f�D�2!��;V����Ǆr��p��,t����S@��;�=Zr��J��Dw�R�r�Q.�e��0�rsB�L��_�6˙�m�E�u��}.{3{�h���,��i8�\Ћ�S���S���o^R��ZU�.�fˡ�~�o��`���I]馼|�>�rIC�0��x���;��J�HS��c+�6U�L>�3��]W;��Q\E}q�W*内�YJ�p��(yz�/��ӳe��I���<�Ly�����:�Ys/�$��T1V�B4L"Uf����Y���"3y������76�h3�J���̩֨��-:'���Ϫu	vD-k�%]�n:��y�7���DÍ-Ե�>�|F`�x.��ug��X(8-�VF��o�)&<��Z��4x̣�;^\Y����4u�����!\�� �tZs;�L�3��c[\���v�yK�q��=�Y0i��\��۩~�pXJ�7�m��C�t�p�N�oC��G��K���Ҿ� �k��l�.u����kR�v�s��2\��.$.Xr7Z�I��P��؟)�|�"� ��ԫ�������YB��̄`y1� �<�oЯ�=���5(g��nTÝ�l��8n��O��ǘaσ}�����Ux�V�6c�k����x��k��8P�עs�:��=�{QLt�uW�8�O�p4��i���s�x����
���VM�ٽ�	���p��1߽��|���`8=Zy�`�L���wѠ��zE^�w⣅s6�gLj��$�-\����)f�GYt��Q����^�����S�;�x�֞�h�쇞�����)�[��=7��f��z4���uc�W�]lʤ��R��	�SL���^��^��J(�����5�o���B�e��e�B��DYv+�ɳX9*mxl�+��D�yZ��o��X���2��r���u>|oj�J��;��|k���X�bEඃB��ޢ^�n[.�N���_#"ʗ�����u�Z���$D"TO�3�Í�sO�4d�(܏��3=d���%Q�Ξ���oZ��hN��FB��СG`�܅�Ytb�cJݙ3�6]n��7������Nh|1�-;��@��T[�cV_���N�>E��giUo�"���=Ý��4�;�KyfGZB��)%,s��p`�Zצ0�V澮|�h��ҏ�\+��F�v�_z�w�;`��˾��}<Rl�ב_�)X�=�*�э��;�W�щ1��\G��x��Y�\hot�)R�q�4��[\�kՄ����H�r���x�Y{�Ґ~�5�1'��6��㸦`�廓���9�б�+�c>G�y�L�Qۃ����`���E�y���H��|��f�@��g�C�G�f%?]z��F���(�_fj��6ƪ���P\;�V������骓�]T���0vK�p��|���	֍�O�P��wt�� l��ע��_���sak���O��ik��	������bzj:���Uy�f���v�]0�?9��l�X#9=�a~{�Jz��#���_S�Ȅ������~��L'�X�1�q�QO{Z���]�Ve�6�!��$�vTq304�V�:��gޑB6�u����7!��\ypxm����;ߛ�F%�Mo�R��a�����f/+����L�X�T��Yw^�sg+�:���=+°���[���,��Ih���.	+:�l��
���y���fF�6����Dt�;*��Ut�c_C�E��o(�A9K�k`��a=�zK�L�)�*0	�h�C��>Ղ���󰖺�Q8$D�6�p#J�z��Z��K��r�{��"q�"�`U�U�����z\c!�����;����W��v���0����C5p򸄰�:�ş>te����̯;8�T�ls׹sg\e��Q�
���~�{�?!���+ڽ��*�dq�Z
��eF���xpk�o\�����=�'�{�B��<]�
o� �Jyo��^9�a�Cg�wt��z�ϹZp��wd��E�*�kpX��/���m���y����Y]7���9��q�|�ci%o+�_�Z���\�s_� �G�byP�,J
�n�ы�J�_ej��\7k���e��<�cД^ZWʲQ"�Y�I�[eЮP�~�v�h2���U�O��(��	�u_)YV�A�B2��vW�����Uo�fR��I�\5�X�n:Ȋs�_zo	z�2�{�U3/�I��K�<
��>�$�W
����6V$
���{��b��m-�g�mvVoEf��0�B���_|�IB;���И5�f��y3�ʻxzW&f�ٓ��Y��↗�\>j�1��t۔,.��p���U;���ƎѨ�q�%
"`~v�����x�!z�#��<��QIm��{�`�b��@[ CXE����W�k;q���v�R�Q�u�9a'Zx��v���眝A-�̇��8V��;��n��?Y��-�K�˭;Uhߛ��n��4�x~�7���~{;?]�u�U��/ҭ�s��3մ���?p�[�]��5���YK�[����bw��X4:Ӄ����_�^).T��p�|�85_4���&'���5g2.^�:�Fs�����o�@�=��V�-t��z�|�״���<���'7ny����p�&r�^��<��xJS��"����E�B�ʦmq�:��b�߻�R����~�Ts�AnUg��/���'�w؜k0��<="zi�p*�>��̾=�f�j�f���Ȫ��[C��F��ip��_0:�W��]6�V���}�)%�>�i4u���v�Q�K`�*��I��(�y{ˉ^(p�~�3�7�XUQ_��X98��|�$И������Y�h�ƾA2�\Д��5`Q�SV��#�/�ҕ����.툫�t�;�>y����xEt�u�H�c��L�����=6�n�ov��V=jM�o���I�Z��W���5�a�}qӮ�]���K��Ú^f��P�=��rŬQ�f�#�<�BY|aU�uC�R��{�M������̹|�)��mR\�n�nY��i�a����{�:v�wrn�	^5�;4�ga�̘��CT��[�����)�V=ܼ<�D�"v��[�=Kc̀�2�t�x{��i� |ƥ��U@��_��k����X.b���g}P�Z}2��0X�<UT,k7�Qw��WNT��׽}'VR�%!�͠�}ս��.�b�T/�����{%ب�jbm<ڻ�=����;P[ﶖ�h�r��Qۜo�j�3 �x.��ug�"�pS�V��[���ï��;ӯv�H��Ī�l�ZR��ν�'�|�Q��m@OV�,�K#��E���3�ՙ�j��V��x���L~�:�!�J+��ˋ���מyB���������"��*t���o�ظ@_�v���X�W����c��
댚6���{��q�^�`��n�+�]��������v�}^��g����/�R8)��<֊xyy)jw-˱Vc�R�A3�!+��&c���v;�ޑGף%ùx��*�g��F���s;��,�f�Ǖq_X`���E�p�]`�1�Ψx;������$�mJ|t�c�-so�Yt�&��c^�c��\��T23��'��5{�<3m�_���jt�r��f�*M��ۣ��=�����
�ݘ��u��C=Ѽ�f���X���D��+,nW쮭�%�:")m�P����V�r��o:�3��RW�l<��jsCy�,�:�n��9cs;�T����G���o%}������nP���v��,���*�먠	���RKG�HV����gÄ���Y���/�[״�0��A�fY�R�!xP���]H
wG�<\�)���]Up���<�����ϐ̡>���oL:S�XV�(��^0�[(�4}�o��h*��l���4H ��k�ߕ�:n}���W<�������Є޴<�Ĵ/	��W�K��Mc����o��k�d�ӱR��U����i����{���\G�-��A�"�]�&)���n�l��D�^wZj���R�i�W��;Y��������1'��glw^35�i�퍍�¤i�*�f
��!|8V�G�X�Qۃ�9���@�+��*��#x��a��2�=�d�
�X���c�TY�/��fi�1�U{��f�,�ܶ�e᾿+{=%��pn����� �.K)uz���v�doá0�>��yT���Oַ~ׯ�T��r� �}����Y(�'� �}�Y"��/�׺V�ʞVQ�ZaV~��{*S�y��(=��[�} �):�# ]�0n
��;+&^���C�A�8��&;E5X+(Z�R��_AoN2����=��܏��W�L����rH��y�NFu���DAm	����GY2�v��Z����J���ɥ�۔��W�:�n���A�dA�2�P�RW�m�L.U�~�-x�$'��6tו�]*[������ј.�V`�X�"����n&f4�V�|����FΖAޡQM��&��C�r�ݧ�^;�m��UL��j���p��Y�]J�d9F)SDv�Q����@y�.�ߪ*��^{���J=�`|e$�z|��K��N�S�m���=��K.��5���'X�\Ok�	�Ǻ�N���꿪��]`��^]_9pJ�t��s}�cY's��Xr��#ҍDu�e)5կ���fi^���QI�`(���5uGǫ5��gV��w�Y.��b���Fe�3�؉�웜���bXj�Ţ�X>�>ز���|��1�U��*���X��b�L�w=]S�z*!�����ח��&y�{��-��u#M�]8�f9h�=E�4Idq�A'�TЫ��0ώ��<�Х��^,]�*�s2�y�=JVb�r_ӧ�zS����.��Z���u�ha}�uɚ χ�j���N�� �C�X�^<��4q��h�;{��M��,�4�εY�7������[����^J�����1�+(���}�w):ni��_Q�P�ɫ��	,�R�Hn|2���xI�:�˸���`��JE�{��kk���'�����j���9��^�`�|Hx��X��WL��GWEd���G2����v�;����\j�W�SgY�� ��Շ;���a��w��TF��O�5�:�P�j�xD�<��Η��/���mR�[>��������\�iS1�)�l���>j�No���{�|8���㗬fҡы~�/�g��P��X�������\T��Yܞ���)�*{�J7y��{簩��"��S]��c^g�x���V��]edu&v����m,��b6L��z�/Run>����w-�#�r��w��V�_f&{U�%±�dۗ�@7f-ޯY��眸�狅(=SY4���{=m�y�f�X_Y��JJǡ<p��L��蚞!S�L��SKj��Iۦg5��bP��Ғǩ]*�F�n���*��ԴǯW%��5��0��Ϫ�%S�eW\�Q�޺sE���<=)Ft�T$��iz��پ���p`�%�!ua�J�.�~��l�bȆ�s�s��oћ�V�^T����I�z�ʦ�!�Zs�_��!2r�t��Y�b,괵�Eh�n��u�m�3>Z����x�폆l36D��-e��F�ZsSV]��e�)N�E�]%d�B��Z:�w^�-*�u
Amv�G_=��W�wnV�z�Mt 6��VB� ֪Η4fT�j>N4�Nb����u�nd�H�hՐk(5,��K��|^b�a��}hu;v�M^7'@ ��|Ig�⇢T�e�һ����x����i6鋩�1�SÙ�M�2������"q�Ã�.<ohlo�3-=G��܊�Y
�խ��4����N�1����G >�R�j3��o�:�oF�4낺�������d��]��3������_]��WZ�d��v�q�y�(�RS�k,
�7�Q<�1(�'t�f��3��&Z �P�j����qޱ��sY٨��
\Z�j�]�:	Y��0�J�+��7�������0A�䮬���#��κaN˼�o��*T$�R�"
���B���@��J}�z��㘬�n.�iLF�N�B(0h}�k���cv�تG�W@�)m�ř��o�9WCTl�bb��:�,�����Y�r��!�)�r�kV6ZDց\)�\Ψ#;*�C�)�������v�;�`�R.���󘄬޸i��a��'�k�K"�L�`|��;;�����V�*J]@�&��y��ż%��H��8�r�5�B%j�:|;Yzί�w]�]p�	Ӝ5�����q��"4�����B87s����$��e<r����C^R�*��0E�'t��D����s��cnv��po��F�n��J�K��ܜ�gP#�i���������,�ݍ�Q,;�{��;�C9��j�Kz�;:�|�3W�W�`9yɠ[�g`��)�[�o�����������R :.l�N��h|gP�;���M̭6��/FفP[&�Y1���q�s�f���Z/Q��3�ԥ]D���b	u�r&.(��v�8ՠ�����}����5.��Q*��kz��#�R������o�'�2�%r��	��q�O�kT����7L�S2��Ŗ��ý��a����ƊN)��tŜ3ijm��ͶP0c�gQ�"�X��]�q�޲s3��Ʃ�4�C^� �B��5N
C1Ӛܤ6@����Y�:�v�_}�w��@w�*mږ@?|����PgS��u3���چ�pD�[��7�U��.�}G��i�`5��.�]�]��wL��䨻�v�������}�f��-1���H����֝����[X�;vŖ%�v���M>`-��Qv:��E���y�V*.�n�Q���軉����dT�k��M����3��G0NL�0����{���Y=�����02/zP�U,�@�w�p��#���U����'|yq��V5�oC֩c��x�[RVZv��r�v>[7�֧��j�1�d���ઐ���>���-�Rbc)-�j%F�X
6�R�W3[��J�T�J4���B�km��J�Z��J����[j�	R�5������m��̤��cs1��KZ(��������T�30�E�(V�$��Z���e�4�A���9s���Fm*���+*֊�Q-�KlmZ�h��ҭ���`�X�m�ն-E��h��piiJ�Z,�*-B��,-+j�h�[E�Jʕ�XTF��m���6���KKZUaKk"(��P�Q��ԑEZ*V�ֲ�Zұ�U�E��D�XT�bҕ�+D��&cJ�F\̀�T�m(���e[h�[T*�ۘVbT-VԥT*)m���
-��1�֖�J�JC�Ɍ��JЌm�(*�U����lh��E�e�fer�ڠҠ�����X�����EL�V�+TE�V��j5i���J�+i`�T�\n[�D�! R�hk�S��5��pc|13&،��a���/@l�.��S��K��`�Ս��ԝ�-,��֣rM�܁�xl�^w.:�=m������4�+�蟛�TJmafn�L/'<Z9�]n����{��4���h�9Vƈદ륝#\|h �y!0޹��qLM����-q:���[.톈�۹�]�K�`��M*��]uR�f:�YB��J����T��W�,;��Z�qc$8�Fa�������+�,��Tv���-өJ۟c�9��ĵS����7��)u��������3������p�>�,F�����*�zة�X�w��gd���+2�kƸv��|7Z�U���!��r��]4�
�!5�����rL�w�n�Ӭ��}���R���8�{V��7�"��{��6X,i���`�}@���'7o�o*����TXC��H�����8;7[�>��}��.{j �t����%ra( �\��p"*gտG�t��P���������^��y�x��9K�/(��=-�v�`����}�s�:K�g�W���r?'���đM𽦴 �Ҏ���й�lxҲ�O��'�5��w+��vyjT3ؑʰ����$݌n��.�02�s/�r����x��3d��*�-K�<�2z"I �vx��%݉�T�뛻�w���y ùf7���Ft��M�ǅ�Wk�i*�p�G��b�0#|�3A�I1�o�׽Y��Zs�R�#�r�ȟ��],�o6e��8+�o�X���K�Ln&f|��;�h`���ϳ�ש�f�����}%,vK=�W#g�p�䎴3��r� !=�ge�A���T.��1Y��`�M��w���3W��������(��4�,g��N���6�Br�}bS�8I��b�����t�� B�Y �z^R�����Q�:=�Z=B�����3=�Id�����o����~{�!�;��g@�esgK��#i�����gs��K�)G���i���A��
�����O{<W��u���H�%@��uZ^O�4�;X5IY}Ӣa�RѮ/ϭ��������B�7�KBq�"�t*0�:W�=x/vn�[X"F��u:�X�{*UC�W�3�CY�a����7�-y��{y^������6n04x0�8G�uʦ봺�����Ѽ�Y_Iy(;������R5�/�!}�u��/�v��Ԛ5�Y@�$��bc����&Q���3�܊5\Җ�ggR䈛k-Y���a`�U���ϪÝ�'͌�G�k�R�w��R�^w(���KX�s�28\ơ��g�O:h�����{�_ie���1:��og�u�熞�T��ю�:�Č9��D!¶H��4���y�xŮ��%���/l%7�.l�kP���"�<�,�тEGJ�bP�����3����=��QB7�˩���܈�=k����}���'�!k�`���u�^����7��VT޲}����YC�TvϷA�؝7]�C�>�|W�*�~�j�Gìi���my�I+~5�ﺹu��뛣}� I\���)i�/JUW�Z1�G��_���V�����ǟND*q�6(kVtn�����r����w��f��5g��eKJ�#�\`�<vT73>iL�9=��qF����\1��*�ۨ#���Qx�׾�oJt�/.�T�w� 2�eԨO�9x�7�{�j����\`�i�	*kɂ�/
mҧU��hw�b����P�~��(I+�m�,b$�;%���)|d�9o�4�ͦ%c��]��F�o婎�{�ߪ���G��V��YvvjJ������b�p\��aϞ��T�r����$���8�M��Ԏ,�Sm��k�ɸr�r$�c��"ɇ���W��st�J[��U�lG�k��ӀN|6��*��TI���j��a�c7���a�M����JX*��Fh��|rҭ��1���Yc���`�}�OE���e�ں���UBvj]�KlҦ�Ǳ� ڻ����3�mS9n)��S��Ld��H���	�.�	B{�]�Y/�2N)���#A��*`�c�_]3�[jm{�P��*!�'9����Ww����ɴVG��o��z�� �Ȁ
����Wxb���BvҖ}KYT��{������k���g��-m(�A\T�'�D/���-.��\1O]{�� ��Z;��{�D�R�A�.A����v0�F��'T�P��.����h�K��#��p�5TN�v�>�'6l㮓Q���.��:�%�J�0�Rx�x;ʪ��]��]0�G��zC]xL6&y�ઙw����4�HS1�)�l����oah������'zh���xY�_m_�ʾ�M}S5��Y�|մ`�|��c)��Ej���;d��G�v3�L40���Rյ,�kk�LL�gZ����{��idu-�6W�Aj�����i�n�����|�o\��N��w�t��c�10Nc;T�\(c��j�y[�ʶ��c�I��v;*� u�~j�0Nxi���p�Lwv��e
�ŉ-�ӂ�ҩoT·w**���N�M���Ab|�>�/k�Ld�|{aE��b.���گ�����%2�\��]���Qιsw����:2q8:�vv��A$�������#�]����}RS��.��<�\A]+����C��cNq��3(Y�F�`����f��],�'�磀U�05��bP��ײD7>�U���wY���v;��,���YɄ#Pe�W
r���b��EN�`��?]9�ߊ��	C��'y2v�{�߫(@*P#n���Ƽ	@x��˪^bᛱȆ�r��}Wօy������zs�;�w��*,�\o�_UqUΐQ!��:��k3}�	�1S��{�����������Y�]�pHm��2ц�E���h�>4C���4%|�ǘ�'}�5�9���O%�m�*��i
o,U��dbǘ;+$ҡϢ�ܺꪦc�)�����L��^���+!ӔX������c
��W�Fa��˙X.x �<T:��V&'�U��.�{�t얋I�C�	�W]k��yԵl�1&{�T1V��e��bQ���J�.ɖ��/:�����U'L�bP��mtv���Q��L�y	y�R�i��rPf���i��,4��μ,0~�jlmӤt������m��J�g
�l��F��sjp2{7ܰ	j����PG���X�}���[u�gNdL�;�jr�Rv�iK��v:��\FG|I}]v��q�-N�o�s;�gf���98�t��Y�ZB�?� ��m-��Ӎ.Gnq��2]���.>ᗵ�ix�K����.�K�J�Y�{�#���49BP�}i��	f}�pry��9l5��/�7/��oU��:��F���|fS:UNDxey{ T�;6�.#p?M_&�����Y���_*h���ynW�w�'�!���U�X�j��V�75C�<�|V��pf�%W�_{y����Ϸ+�+��ŦJ>�Zf8���N��7�"�g�nx}0Vr�7�܌g�!������-�����K��6�09;+�iS�'m��7~)�cq���3��;
qk[HP^c�|�'�(�S.����:������W�	��F�S���tOk�j�]�ʮ7�eު�hqŎ�fUo��R�qDE���]���rc���郫ҡ._:�hU{���P.���:G�bKG��]����IY4w���n��ϒ�P8붼6Y����,�,�V=68�}��cXt�$m:�tt9��Y�O��qǏU_Iֻ(�A�َ�����9�ع8���뗠
�"lh��:)Ab?vvu<�l���^aB�w	V�ڽY��l�D��n^co�q!d\��Kz��G�j�ѕ���`� kp��A�_��"��,x�� �I�*ӈ�6�"�T�z�ǃcܗ�v��v;�=�~���9��å=�o��^��,�K�EL���V{X�_s�N����㤜�)���!��ɑ�>����鐡7��q-	ǜ��N���y�+4��#!Z���.AC�-�/�ېQ�����U�W���17�<��d^�ً�lZ"SY��z�* �U��n�wk�N�[�-�i�5���^�	�KWb���r	O݆��ߙ��^	BlČ8�n�dr��gb�T�]Y}�X�$��Y��w�����݂���E�s1��Yu�K����VT޲F.�������yC�c�}�N,������Bڇse4�$CA�#�Z��~�eˢ���&c��h��4����YB
�3pZ0�W*gF�V:>�b�k�BHRbzk��uP#
�ɽ�[�×�����O��Uꅜ�[q+):@�����BS՞��}9N�=r���3�̈́�·�i٦��}+*X�V�8x�0}����K��]Խ���d%�q�b��\�+N����%�S�$�g&_C�P��p4[���Z�غ��J<��|�,�O]�O[�ݗ<�o�s_��,�4�/=;��[Ki\�����ѝ��45Cl��q�<A����ʝrW+������r�/!�Ρ�f$�m����t�����zE�|��ݯM7��hĵ�ho�R�~?���n״'bd��b�V�����w�'»L�@��{BJ���ɂ�>�+
�T��Ju����k��.���4��륀%��O�C�M������h�zT+�rJ��N�m����8��/��E�O��Obi�ԕG6ՀzY1�w����azjmt~��e��txx�?#�s'��dY'�|�Q�h�)p__L�.�y7���o�{ɄȔ��$�J�Н$g����0Ы��u=b�41r�sﭵ6�*yC�~����g:���io'��}(�i��\�upJ�1� ȅ��H��F�������j�zJ�㲟���c��[��Gq3[Pգ��-E+���}�|����Z��W\���͊��W1y��-U>��f��QD8�^X�]��b��ΗE����F�e�]���ir�T���m��{�檩:��$��.��)�>�n��?>�̫��<(O#z7���V!@�����M���A8�cN��m��T�nK��@�;���0�O7�K���q���sȇ���y��=��/!�]��.��Է�9-����N���)��vz���nV+���a�꿡���_E-��V�7�U��]�x��V��-r�yt�x&]�����37���0�T�tJd�7�M��џ��d.����si�!\jV47=�W�|)�1S�*�}g|tU��A
ɞaa�R��-w+�/oR\��P�s	��E+v��m�u�U��_�?ʘ�p�\YѲ���^��۩4ɵ���u��S������G�r�~���Ǘ՘���;T�K��4�·ۢŽ�&�</�e�ϵ �`L���)� ��7O�]�ѡ
A��9|��؈�t�CBc�͌W�ד�r��57Q6�\ts�q�������O|\Ok�P��Ғǆ��I��./
�%1軒]b�ϭ�i���ܪ>b���l���8\{c�N7�>�-��-���r���S1SX����4�E�~�e2ꗘ�f�f��mP��ܮ�����'�ɠ.|�����uq| �)":*�˥D�U�f���W�^�<弡��ӆR��t���V+��}�屢8*�,������ѭΣ]�g���.���;�^Ԋ>8��G(r���-�f�5J�u�eH��WwX�J�F/�]X�7�rZ}kig��>	t����o�4P�l՗�0��\�@/x�77���*gt� �2�^�Q�̬�c7
�:�͓�W�x]�,�w��_��c�6�kFy�]ַ��ؼ9���7�+B��u��U�V��O�T�4:���q�w�b�;�xY�]���+�ZG��0�~���|���B�b3`ߢ����+�犁�D��]��P"��l{�n誨-�Wp���2֮��^.V�τX��&gt`�}AEpWl���K���x^�5d}��ez%���|/I�tGw���*�إfs#���<���S�}z�_��L��c�.�I������^ݥ�H�8���R�;s��V���ޔ�M!����;�>��Meach{�����dc,!���C\�Zh�en[8��Ju)��O�����m61�kt7v��I�!h9�3)���(�CsT
��em�\Tn�:4oܕuw��%b>���Ū��f����ܨ���������w�ظ@+�+l���k
�C�m�uѿx*�v���+�\w�ZT��ش�Gñi���<�f����w�8Z�����}%4�7q���
���rԫ�!����z*���ir�73��}hp�YwJ��P�IG]:�r�wjM�G���x�%S�j�6�0@�v0Pݙ�c3��i'k��Doj�+#T�����KЍ�䮛��e-�t�u����{BEYo8V�AÅ�lH/X#<�%��ӎ2���+2�s̉[�2Pڎ�k+F�=���&#oq?@��~������Dn��í��&^h�]'g^�+u3���)\�ӄ�&��Wcʔ%7JF5��p�����>P�U#Q^JR]�^��[�L+��U���Jv<'�����s��S���:t�]A�m��s��c���|���0�ҬMmv���N�X�(���|��鵙uzU@9�{V�$&�ڝ����קdD颦U��<(n�
V���u]�cU�z2�в��Yå��jQ#���s5Rs������Q]n�oL�m
PLWX�,w���k�%Սk�Uf[�1!9V)�3]�ɍ>0\��W7��=n����45.��)��My�l:`���ľ��ĺ*�gL{mVՔ�#�)n��Lp�7�9@�8���5|�MTʟJ�Gõ^Vu Uֱ9���X��]״Ue � ���L�M�N�ɏg������z���PΜ�ɼ�156���%d"m�ޒ�@&�e��b��>�sN�ܪ�f�D1Y�^qX������132�=�7J��UYZ�����w`ʘ�Oh�uGU�ywmo���%<yt���e�t���>�f��� sV�UF齷����Ew
��f����Č{5f�*�܎���<�Ժ��]����ԣy��.�d��ʹ��Sk �H��g�rN����]}���[ۜ�웶�Z=e�z*�fk"�N!;��i�"FRY%��&'Y�aӖ;�D����"�e9��'rCi�B�F��7J���f��ޮ������u��7$v��5�:��R�ԥ��-IQf�]��e7��)�be=Յ�)�Z� ���2�����T%vl?LR��n��L��`ˣF�k��L��%���,n�����p�/��J��uW�\Ư�Qszwos�Z
�}�i�7����.#zOW9��:]Y����R�\���"��5��3WG� Q�/��"��w�����U)��o�x"��T�"R�gCh�Ů�ʔ�cG�
�S�ݰ��h<���f%�޾�j�_	�")&�iuG�[}��o鯞�U�����#��Hg�=0U������.���#�+(-�r�M�SJ������b�w��N��C���=��崙�O��r���Z��v-��/8���i�qڅwj�LY��[��Uv)�=�(�c��۸��=��Ƶ �E�)r�b���[Wf��3��r2h���M�t��� 'Vb�ʘ�3ya��\����%Ά�U�:4v.��T0��z>���$[p���w��z���i�"71��Wwt�Ruuw_4A)hѶЩYc*���["5��r�*
T�e(�AZ1�D��"�9C2��lF��)Z+Q���TVګiQZʌ�[Z�E�Q�Z1Q�V*�V�ŶLLG(V,YR�����B�QYU�*E���V�*�QX�XZ���Z5"�j�hƥ&8��%�E�X-Kh�kK`��q�*�ae��Pm����-k[B�j�\LAr�+j�QE�m���Q�J�kS-��miA�Ջ�U�(�"4��J�m+mV!iX�*"Ya`���EƹJ���Q��EE�#D�V"*���P��TFUUK�ֈ[R��r���m����V5��m�m��R�Pe��+R+iUT����
#.69A��l�"��jʕ�l���Z�Z�(�KZ�V"����U��Q�e���QE��V���*�T(����UUD-m�
Q�F�R(V�"�mFЩ+R6��UV*���W
�b��� �-j��mRڰE_�W"�k��fR�el��ӊ\�`���=ݸ��F�7�+�wN2�rg;{��Q�1m����@l����ʏ�'E`esiw��<�{?Q���W���ڕGn��;HX`��(m_*���Z�i��!�:�c����T�����|��=i�v���{��Qe\/DUW~�5���]n���~M���<����}�}��[.�O��,�S����Nh�z��o���|0�#�!Ww�{��Y�c�)-��s�2���M��e!��Y�R����'к�͝,�#j���z(��%�,�ɖt�b��3-��C>��ͽ0鰞�x��fS0�Ke�!���C��u��)���;��� p�Z	���a��	��09_#B�7�QĴ%P#���[�*ۙ�]י^8��A�/R��.AC�>��h\���c!�,;�O��j�r�ǭ��"��[U�i���]�F��~�Gh�����N�!ll-C`ݺ>��Sz`��f�Ρ�ݿW}!�tJ�+������TYخ�,-�4��壶#^}�b=o�&�.�;�
�r��\��.�`q�LJ�^��u�0��1�U��T;�e�d+��WB�>3O��%'^�z���bΥ|������ˬE������PvA�qc�	)�יuۭ�}N�$���]o]��U�oN�����D]i�VغGrs�]�Yg
q�*.�V�/5����)��7&�˨��z��M����1�6���﷢��@��$A������{��q����WJ۷K)W�^r���;*��zk�&l@��x??b�mׄO�~w	#d���;��Y����~oy܈-YO�ք:�pLY�{�¡۩+�ܰ��ش̧)66��φ[�Ҽ9��{4[g) �V�P�N�w�|n�VT���b�����>,,�굵�[�/�<����O@��<Y~��������:�	��c>���=F��Ҁ=W��ͨ}�y����YB�c�r�jfC�-������ɂ���XWmҧ�zS��6���~0B�)��e�3�m kl	��}bm�_��l{�>����vP����b�>ג?;ڭ�^�r����٘H�ڐ��F�*&wyU��w��)���P���\�dw���di'�h6��y��+j��-�6�*yB=�2j�H�d� �|�ɳ.�hZA3[f{����?B4.��c���
���~Ə�uE�˿sOw25�x6���r�7HS��C:=��W�� <��jx���snG���\������-X�>��!�].�[��%@��R|E����.����KR�Y���CZ{� �����SZ�g�y�w��1��N��4�+��9�ҍה�-�>Ǖ�y3�*z��	�ɰ9�l���X�0'��+�(�>�Ѝ��)z���C�����>O��pz��"��t�Ip�E
��n�[uH�/d�V	��c�,���d�� ���p�*�]2��Q����X⟧���Wj���p�"a�Ţ��K�Yb�}+q�0-��Nq��w�=RY�d�Y�U0�$������ޞ��u��$����������w���� w��@���D�~���ͮ�ȣ�]7kB�L{�E����F�V��-r�r��9��մ`�|����݈;w���:���lϷ���=���~^B��r�0��nxӘ�pW���B,��j-�1�;v��@��ϥ@t����=<�n�y�N��k�+�"\0�ݐ�ٮ�AS�$�����ĥ�z+�}���WdJ�̇��Rd�9߇��L*�e�E����L<�w8D�b�VDM��;�	>�� E�xڗ^��o�)J���h����`��R�1��V�>�m̾T+ue���&�f>`v��KԖ�L=�M���t������n�Mռ�����Fk:�Æ�ɮL���&G���-���Y����b/_e�{�/�9���%9\l7���q)҄X�"��������:-�G)S���7ru(a�
Z]#l���r/P��[�G<��U�����'���o���&��lE�9����g��WP:P�Ԡ����1*���+�4�Z�#b�j�jN�N�C��9oޅ�W��F_�������L	8mo�j�q�*}�̩�ڬ�9>��o�Ѫo 8b�ʬ/��k��_US����\��>�
\�wk!\����������741K�bf0�v.��b�O{<�������~�J�]P.UmU�����t��ζ�_9���yj�*�G¯ �ѣyߨ�����h��;Q���˙U0X~��;��ߒѡ�Ok��B}���L<&z� �hu�ͳ�_���Y�X�~ ę���.�Z݄���hU������^"(m�*���U!n�ŉC�כA��{/7Z�2�T,��Ԏ
�)zM9���/|B��B]�
	�/�J��jϒd^/,u�:�������|'Y�5���;��V���w7��H�Pp[ڬ�'M�8-!��<*�_��w�;	-�|{��@ʍ�x+MծF�_'�X��=|�VK��X�y�����I��lo�� +��E�n�Sy�>��4�v��r���S�9o:�[Lv�;�'
�6b��]+�z�$R�J��Aݠ8^ܛ�i/�8��%*��(P�nn�c�ݢ���k��\լ�c�ԧ�v�P�y��X�-9�3)���(�CsT8�����{O��������X{��L�Ը�}�[���s�!|�Mw����\ 
��;z��C{rI�5yf����Y��r��lD�@���/�J:��@�Dn5��"�X�q�t�����:y�`�=T��f�`W+i@(F'�W��	���<���}����ޡ������ӈ[W�$q7׹.�/<�\���AS��A�2�E�=��t{U6rm�}d?1�ݚ7�la�9-��c	�=����Q���G�Xψ5��u*מ˯j��>�,c=����&>��Jq	�=3xө���\8G��e�B��N�?����M���*��WTFKj3XY�Sk�,�Ye����zP�}��\�\�epb�nw�=GQ��T=��'v[�����'6�æd�+���^��0�U�`��-sS���FA��8|���s�X8}B�K�#���G��.�;6էY������o�}�P�����A02%
��w���JY�U��v�Wjt�@k(�Ź�e�!E��B$�A|�KT�-	�P�!n�.uû{V���=v8��i�P��7��}NG{�69)�a��&s;6^����]�����'�v0��&E��"�G�y���Xk��=�ߒ�=ېQ�w��1�����mc(_����ѵ��x�~�P�D�g~E}�����4��t	��+w�lF�p��d��=�ު;[=�����bOk�Hm����^��Y���;�:�TZe�}��(�u�զ�<�7�'�
�*{���.�`q�	�B���,��?J7޺U�d�H�)��A�n(�Y��͡�{z+�O�B���l�h.�C��/R^a�8߫vH�P���R�c�v���8��U� �a6������n3FL�����m���Ǫ���#��`�eKuDo
��2��BS՞�*�tsј/���^Wï�G�,��H>
߾�v]�pu�W�%/:����R���PP���/���vnas'��o)��Õ������P����Qx�ׄ�zwMYzު�P�W��p�h^.�'H�V�!=�a���S��C��S2WD����OJ𬔠pn�]%�x
S���Я}�7��3��C���\8l����rm7���rT���8�LX�x,2�2�]J��an����*񣊼�qZ��Tas��v�P;n�s�$������w�=F.C.H�!õ��ac�Bww=�S���uybW.�M$/o9cKO�Wl�{��A�I0g��Oip)m��
��!�6�WK�d�t���\j=�^��;�����麘4��n�|�3��xH��ڒ���,OVK&,��Z��Szص�����vZ�X��7��^1P����҉h$4�˧3��^����0��}��5����4w� dm���*��Wh~8o��@����Χ����ʙ�m����^�Ώq@�̃&8�G���4=���++��xG3�N��	Q��UHĀ%|+Gh�]��2v���|߻ݻ�/)x6#w��_҅E��V���-j��Y���{,�%յV�FBS�;ӱ�TE�B8��(47˫��BJ`\Ɂ�ć�,��r����p�@��2 =���{�+\I�j�5�}l�Wl�}*v��G�����^�BE*,yV�㏩��}�ǼQ��u�'�6�����*�˸�V��=��C\�h�����F{ݼM�U��ܥ���o�צ�6k��C��K�sƜ�O����-sx<^s�{cyR�R��I��vf�c�)J�1{u���f%���;^0��	,q��G��j���S�yu&�C��q̧��6s�=��쪒4��v^�����E�)�1r;v'����N��<O}��f��7�ӕo�*�RJ�j��L���};e^^ҝ�Y�|�5;�n�A]v����EyROl<B�u�������u�غ�j��	A��g�y�w�+�Fi��>i��Ř�<����Y��\�����3ހY�Ժ��+�R��+�_vD���x�%�������ܗ��)�nm���K�t�e.�/6�BϳD z��Z><�J��%=�޿o������o�\Z,��X���6Ο-"�	p�*�yܕ^�u5�,'�����d��㕍;Fm�_�3��U�զ�(�M�.�<w)�T���6Y��5�^׵�Re����9�; �Br��}Z#7���T^D���q�Uq}TG:J$:��i������0�lb���7-�O��Ys>uۉ�S� �U�q���0��ە�:[(5�Z�Ɋ�`ҥQv�t��?S�¯��jx_;�K%Z��\2� �*�*���c�ݲTz�T�\wRHzMl��g�Q�{��lp�8̎�5�}�A�Q�z�њ�e���s}o>Ə���j�L�u�b�F��8�%>��Sr��6��π��o	y�a�������ʊ��֛�֤���ZX,��Wq�wg]�*ԝ+��LyA
�o�sh����w�E��;h�D*<{+��C(����g�\f��N���������R���%!��Z��e+Θ�/�$�Kv������~�$v[����X�^��B���UP����-q�uja��إfs#�{��:���,�Oڔ�����4��`��pT0�"��;���]>�XL���O �=�B���\��}�u���ך����X(���d�E#e��a�x��4xm��̙)+t��]��,�}~�ia?d"��ڀ����]�`�e3��<���P��0��UJ:����X��-Cp=+�FU/fA�y�e�z+�U��踕T�:K��#����۰�R?J�^]��EG�m?���O�>��\x=�.�<�f]'K��b�ȑY�=�I֖����ť'V��3��L8K�#���¬�����Y`�K�Z��vo�^jW��Wy�X��u��ք�="��J���Q���jV�T���B�EgraoP���{���SǪ}�B��)�2������G�9dp�%ٓ�7\E?
�V��nm��5_�7�	N���;Q�zu�D�K�U_����	��`��B��	�����1u�nL�GǬ�]/��z)^ޠ�������.Ŗ�lwv����'d��]�VX��vIC.����m.���Q�����t��y�N�r���1���T�,w��9c�*�@A�q�`G�osE��[=�Y�6ʮ��2%�f��X�2<�|��Ѩ�X��]��{����pP��fR��,�w�s҇�U���~i^�t���7��N,^\џ3�@aC덙�es4�<������c6�<�-G���mfQ���T�fY#��]���Vj��Uu��ų[���24��򻾷3�Y�[e{ݔ���x�W[�F��8ey�Z��r0*!�B���9gx��,�U
�W���Z~� ��~�s�ڏ^��GRcj���`��ɐyU� � Q�9��x�M�i�+�73��nS1ͳ0�J��R�EV2��?�ڐ՟�!�&$aϟ�ѰY�$��a�yc<�}����pq� �U�&9����v*$�0U��]AWK}I�N�1(m���b��bp瞝3L���1Z5����Ɏ��Xφo����!hH�JN�U�z������w-YbH�	������4���R�Rc���s)�o�c��Ƙ�}0��W��į<�AQ�$U����W������[t#ɶ��-ǘ�]��zFd7��
g2�C63!HM'�Vwٺ��zH����5�B]l�=VO"3���t!��t|�v��;yM�CM-�P*P�,gF��γe��ϋ�Q���9Q7�[ �b�Y���hpW[�fP�6�D�X�X)ug���s�M�f%��cRG�5��Ov�@4�F��௶�'��N�n�4d��(��;��R�AJ3�1�b�Z����ׂ�ζ������k��<��t'��*΃l�g�1L2�F'��p��kc��!�1#���ZK�Q�����g/�F�H�qr��5�b��)2ʋ�@P�VX$�ȡ���;4�T`ֶ�4�/4
@�4�Ej�����XK����k�h�4�'�ꏃ�!��|L�Y\F���ި�M�l�-dc/$�sL�sb��qoB�@/�����~�����Mk���̈�=̔��U%؎cv�e۱.�@�u�8��o�h�.;�<��-�����r� 6Y�)m� 8x�̷'B_[��!��1[nM��jP��e�ҍ2b����9�����q�i��8�jv��m��|�}X:ր@�]�Ľ��Dm��kT���V��
DL��u����_M�?
��\Mb�������['��ͭ����U����z(5�ygw3隞:Q��3	9'ɽ}1�A��˕�+0(�@"���fN`����f���T൪��9���7Q��Ԅڣ�y�fJ�44��9[3��qؕv6z�[��[;e���J#��r��	�v¥�q4Z�}X��X�=�L��@� <D��V7zW&�����"^�o lo'\���{+�.�iP�OE�ա��"ȭC:[�ڊ�ہr�:�x{';:RĜX�����뷠o,,��f�U"T���55U�fj�7�.��S����s���V��m����r��)ٯD���$��,ؐ�2� �-Qҙ�5K]���ءV
�V�]��t�r+k���.��&ի��X"�x��G���w�����=����~���;X�_�f3�q�o�q����������Ph&����{%���v���%r�Y�]W�k��%"��ѝY�'�,���)��VӼI��j9�ct;xD���2���<�ͬe�6*�����]�A�k����L�(wYF	{X똱�����z��ˏ��[RN�t��>���V����b�>����P�B�������{��1.�|�0��U���F�X���4J��O]u�
�ȇ��LX]�/)_g=�HOvw[D
�;�۱!ѵ)��J�ZC�3�k0�V��5���B�����'L6�EyV���mr��_+��D���f�,
�
�u��8Kf�ٺ�5ʚ<��nfN�W�p��9 y\�<U����$5��8+�C�բR]}�NQ����x��i}�Ӿ`�kTm+l�P1�7��QZ�DF6���,UEQZ�UUmlm�E*
 ��nZ9J
�(��XPB�|˂V�XҶXֱk(��_�ʥVAe�[m�mb(�Jʪ)mE�-�[lZ��RL�&[h֥Ie�eG-�
�+j(�j�嬎6F2��O�*(�1��S�rҲ6��X�d�[k�Ec�mUA`����F�JV�Yd��X���"�(��j4��B����b,b�U+Q��*��*��j�E����TE���j�"(�b�O���Xڪ
(�>8�J[h�EE(�iQڪ�D�iQb(��"
��Uѥ#TF1|�Q�*���mj���ST�(�\b�UF�*)[������Rڱm��ň��|�mm(�2�P�TiEETPX�ZX�Ŋ�Emaj�%J(�[Qe�Z�X�R�h�<j"�j�#s&8�EUEEZ5��)jZ�B�1F�UEbV�'��ޟi�6�5�߶&e�+DJ9Z큖o##�q����kZ�B�=��R(���7�y�6�޻��We�4��CSt�s�%�W�:�]�~��:݅��H3kƚЇ��Lf\C��):G����7ܰ�}�{����{Q�,�����{NT���{M�U=��a�f��4�,��N{i��A��LW�ha}����]S���1����4�V�:��zK�y��wk���0&:|�3�(^e�%,nfOM��+h��;E��uR��C��jfBz[�0d�u��#�/
�z�c�3I�Z
�m�Oek�V˿�UL��(���\$��d�kΌ�&�p�{^��uq�CɌ��˚Ѩ�׏gtx�i4%AU�Z�/��W��Q"�[RU�,FU9`L�&��|��`��=�~���u��t,�+zî�
��!9���wN��[�m��x���+d�u{ORa�z}��Os����!�ԏF�##Aa.��c��j���hɹ����)��~��kRB��jz���++��xG3�O��F2�B��wD�#�����F����~J�
�����g���N�Q҅J�XGx{B>>P �*�&Gf߇�f�ZѢ�}(	il��?\�����s������V��:�ڏʅ�˾�\�d{;��Z�H^��V�X<�f�3������mo�Q�������u�F�<����s��s�WD�t)�ݮ���i�4�����x)m���=����:뮐��v�2��_W^p��2`b]�:�^"���ב�&GFí��G��̫��%_":��yh��K��)J�ڏV�j���axbL�tF7u���_����Ċt?V�6y�^��I��G����^]7\V�����9�H�7oA�ڸ�!����mr�!��L�[$�#�>O-	��^���[��>��Z^V�\���į}1�ϫҼ{f7L�֚����(�Ұ����������Q͵��L�"��{�43_��w� ؐӃ�{�ǆ�+@t��u\=<�����զ�����[��n�	�֦��^�VAw��!��_�� :����c�u����)�d��pǫ�G���v�=C1�\^<or!(����l2�j�g ����z< ��٘�X'�.'��!u���X�B��yl�cyI��Sy�E���K�F��\�Rl��T|�IT��P��W^��ոEJWo68FO. u|�ǧ{��g�ϯu�i��uӣCg���_|�$�;�ʐ�wy�ykVY<����o;YW{��[��Lj�a	\[�Aj�-a���t o��fg:�$m�g��;��BMڠ�5�Ϡ3]^��μ�+6����N)�ާ\���YՍMrlu/*cє�Ҩ��l��)_ ��'
���8��}`Ω:���5�X��9�-dCL89������2���a���K������
���h*������S�c��`�_�لNx,��/{����G��Dl���B��=|�ڧf��z��\��i�A=Ay�)���yգ��Sz�V��dbǘ;+ �J�̥�ԗ�Ӌڌݽ��⦁��rT�VP�+��aѳ֪�\�f+cj��+��q���J�a5����=���2@��bU�b�o���-�-bP��K����^��X"�a^mn��R��k<نc8p�ZR�JN���8���o�]���M�6'��kU�(�O^]����*ӣ����{G*uK�!A�6"����}t��]�	�x!4-ST��]2��1"=&K��m`�K��Y�H�S���dj��H�eu��ٞ�ч.@i�~���f����XL�%k�T;z!�O��|������75C\Z9z�{��uW�����#.z�Y-0i�/3��Mk#�s������Eį���I0��,!lg��.�=�`N^/�3zQ����;��k�2�5;��FosA>���Vׯ	��{�:�펽�֨I���i�}�4�j`�g�w��E��3P�o*���K�.���M�;�I|��f�#������ի�J�h�i��M��O5&D�;a_���X�T?���W��be}��:>W�J,v-3$H���a~�|4�#�uH�\ѡ��v���eW���e#���<*�^�uS������U!0�mw�_=�kǧ.�;��{C�\�)�ؽ�|W��*�������[�/����0��u��1 ҝP��0�֞�l�d=�x��΅��,g�Yh�Y�5�֥#w�/��/E�C�T���R�0�u4��L�54^߫Ѿ��,9w�
w���	dx�\=)�+Z����J�^�fRe���.zP�-������}[حˊr�Ul��|r��<��X,S1i�[A��
x�����N~Ҽ�9%��D�o����9�v���)V�H�U xĴ�1і�ɑ�?'���yf�^J#���~���]�7v��|�Z��9�	`�(t7�H]s��b��*�#h��`�2��k�����[~�>���uF$Ʊ��u�L���@pC#bZR3˫<U]�^%4eDY]Y[�[9��U3��zl�F�=ܠS�1�Z��I����Ա,�z>6�oς2�ۻhl#s��ه�V���c\.؟.��_n7�cv�]m��x�3zq�|�Q��"�!f<z���9z����\{�w]8��F�`�Nv<R�o*��Ij�|��/��!�𘑇���_�kmU��BV�Ȏ�Lz�+�p֎��"ʾRm���`���E��~r˭�q������N��f��4�gN�0e��,�7񇲽�(Vf�/�lj�poEuH>�_H�}n�:��AI�O���Ud�5.�7�WZ6}5xhq�w�c�^��φ�V:>�aW-ϼC=�k�T��߭�*NY�οiZ�*/��^�̸�2��x�+ݣ	��H8}�	���]�ǆ��}9�Ǖ���7sr�i���v�J�ex�Bh0��}�n7�tR��$�D�I��w�����)����/k�P��Qx�V���6��g_�%+��6�d�s��D���R��6��[c�+��]\J����2T:�2`�o��oK�i�rf�C{��s
���U߆BI��,���Jβ[5��̤d� .'�goog�T:�$���M9��eN�t&]�ɀ���V�ш�3~�U���9���O�� �����r�G]N����]�7��0$yu��}�f�:�y�&L���.���7)���Sm���a^~����éKh����	�����_v����p��V͐c{R�vf�[˨�Mtn�,U���>X�xGq�6]��鹜25ݷ,�Z+�*J��QN�ۛ����"K�C��6G�>������8��D�K|���4S����ڧ��t�z��On�ݞ/��f������	�y��Xj��*=��@����Χ��oQӪ`=��/���4�a�囝��y��fW�t�K�3�N<��Q��D,�z��{�}��V�c��#����"�ƕn<k��9�Q�:��5�:�].#��P �*�hɻ&:���|4y&�OeaT`�]mR��K������������}��UA�(YU��z�]�5�)l�p�^e�%��y#-c��P�f���Ϊ<;�*�a��M�w@׳�X,^�%\��R�f�FC�X�K����߸/b^\sw�7��Gz�����c\��ʹx^�ή�V���}�M-�;��%	�C�W��,�*���9}t�������>���-�c�%NdWY�:���C�<��J���;�4/!����Zx`x[�u���Os~˵qz���jB��{���Π:W�N��޹}�r��w�E/4$�fz���Ձ��л��%�#�a���nd�罆SV�&�ڑ�@�u�6��8���l�ԛC+���]�\��ޣ�X/U��:�j��7��{^��/�5
�-,Wg+9r̮l�]�i/[�}���RW�-�{�uf�7Zi�}��ͧ7Dk��m���r]���n0�Y�k3�j��p���dۗ�A�a��������)2�Ku�+��\�|���,�6*��͖�RV:��U9������q��U��B#��Vy_�P�}�ޚ���bu�=��ϯb�F���^���*�ps����)i���:ih5<x���X9��L~���a�6���z���WPU��(��j���	@x�/��g��h������.�UA�-���	�,i������u1�ʋ�����x�����yg/ͳ]���O+����RN'U�k3}��&�г{r������Y_LG�XX	O����o_j��p�T:i4��4%޹��"���f�U�\B\��V��,&�k��6�4�}��;�,�譅`W%�y�����u�Z���+9�X���n/C:�=�w�A7/r�_x!���U!n�k����]��u�����ūYY�Ǥ�����2�!�}6灻����L�B�,F���f���Z<���k�0��=>���O��Qɇ޴�ڍ��-XPh�y��L�t���'Rf�tNCI�rءQ1��Ys�Ƥ+/������@n��Naf�aǢ����M]�w�(:nP�D�ys
e�;@fB�a
�r���ܪ`�]B����i����Ӳ.J>���Xwn樼���-:'����Pë�.ȅ ��vW��}Z�q�`��fN�����=�YjՎ�V��oLH<���e��{U�F���R6Y�U�G��^�'ʏsx�̢s�E�f�e���^�}�7�����-y�`���3��-�9v��gt0lӊm��җ<�A��B�+��ˋ����{"Z=W'd����O��<��yx��n�o�����U��2�Y��ி�]��b&��#�Bk<$!��h]ȼo'�����mW	�̇]�c��k4��ׂa�_�G6xU����:�s��{�ѵ'�i���uT/>j$<����4��;o�)pv�h�3�/!H�4��#T�bǛ�e�v���Я\�&A|egڃ14�T>��C�k�����d=�Uq�3]���m����5��z�.�x���b!�̪@yٕ+>qq�`Tzf�U4]=U���m���/|�>�G�����e�"����]���B�6k9*m{�e }���[�kꉮᴌ��z���ԼQ��!C˫Vm���d{��Kn�`�%��J �6�_1��G�ߝ�mu�}i�=�����%�ŸWb3;B��J�ѵ������@4⳻����u˪Uݮ��Ap��GE�1q{N�h(�=U"�F��"����&�2����h�Ӟ(a۔�wu�]Qߎ�*X�bƑy���`��ͽ0�U���jq�X+��:5�xT�:�W�-V�$M�P7��]l�-���uQ?&F����#��C�D'��^�_�a�k˒П��"�b�4(R���I�}u|4d�6ҕ�}��������/�ʹ	6.z�ho;��ã���e��P�D�gJ$����ԭ[�pQ�q|��KI�b�$R��g�Gi{�X��Pb]�W	��>�!�1#���kC�	{7��(,�+!h��jS>�nx��ef�0UR˄[�0u�.��|.-i�u�<����7f��+��6{H��8l7)��91��X��f�uI�B�~.�f5��:.ۂ�}z�&��au�������yT��>^��πݴ���7�ꃆ�{�(��r��6�*�n�aWLp��]>�f�?��/�ʰ0��P4�q\�w��Z�L1�3�s��S՞t6]��ym6Oc�6m+m1��}���{Y�)��[f���kD�T�ZX��E6�����]��]��G
J���"������V�3��
:Ɋڽ�����Y�go>�f�6yPx�Y������M��'&�iͫu38�{�5^��Fz8$��kRY�ŝ�e,�����h�&��/�jJS>�P�L%��㲠���Ɣ������zL��r�l��X�w�79A�W��y�,�;ު컇j�1b��a����U�+�%��;ŉ��u��k��[�c���������t���,�8�%��������@w/��_:�So�xh���aw�럙99J�P�_��\B[`�`%�lV>|��i�]��_d���WQ�a����ڼ�{"�{�1�NϷ�x^	bs�N7�X:x�
#��Z%�^��|e�r�51���]���Ϯ�*Wy2=�M��Ǽ�N]v�G�o]�p�C������[�lǝ�F�*��ǌ���תyC�~������#2[����g0Y��:�6�e�E�vs������t*p��^W��`l;iD;J�e}��>Y2����ve��s
�ۓ����fU\�Y��.��Z����u�v�ۮ�\QW:2����f$t"�/V{�b��k��H;hAN�G"���'����p�[�p��UQ��"�t�ge����n��\�#v��Z
���Y�S���#ɮ2��C���]R���!ך��z�\�s���+jT�_V�ik1u�s�{zbd��mMV�2��<�CN�Y$�B�4�פU�����ۚ�Ӌo��<ޫ�iqj���dQ��'!��wM����6V��kMb���ׯ�n�aS���`ami��v���T��"�s��mT�J��_1 �z	�2'g�S7B\��l*���{��4Ϯ�뢄`�Er���8�����k�ϕ�K=�7���-�Ԏ�o:��N:�����Y�;ycӘ�kJ�jӷա0�[�HZ�i;���AMSQ����0��a��f��ޙ�5F=/k
�݆us�|Ҳ��Ň���-�N��t�������_׮��3�[�L��0d��s�=}�%�V5�9bSNՊ`t{o>m*�̣x�K:M�W�D镔k:���O���=~"v^�m{�J��ݨh;t�I������l>8��X��ەi�dy������ͳ�񦀌�D�͟t�R9��7���~��6����6��:��P��̰i����eq��Lԏcj�Pչ9R{k��jm�YS�){���_^W��]岃,&2���<;V�s�� �I�]Z�Yr��5��������b�W<Zm�5:E�(�������hTѫD4ս���5z��e_C�*T%\V+^���,ܫ�=w���@AX��I�x	�7h����Yo��8�gz�q�Fi�)�1ml䊙���oR�]̋�ꂬ*x���Y.��.��ά0��At,=��$���ҝ�;�6]\���',�1Xz(K87yWwVt=f�X��;� ���0��[X�aۓ� ԫ��굹�*�DPbyɪT��;y �D�R�tD�*>���qe���ak�cy�99�B��l(��'d��#YQ�z�T�P�����C;HC@uU��ؔ�<�ׁ^�H@��]*:z�sz.��ݝt���Al�6չ���k��nq#�� q��2�N	��h�L�8�h�u+�2�	ԴN"t)�Au�#�:nhw��16[9���������mge"�]�j�Gar?���t�S،�ٻ[�R5k�i�q>�\;i}�5i�y@����`�p=��<�цݘR�_�O�[����!;�=�hF2�\ⵄf�y+ZT�µ�K�3d�vs��l���
�0�.�:�V��
[8�����������x�BvK��/�8U�	2L��q{Pf^@WC���Y�w�i�|�]褴�n�}]bP��ާ:��[ɾ������<2�;�8�On�]zv��ڐ��#+�EK�c:�4-���SC��"�,�[XD+{3	��l}�6WV�{�Pi��Է�Ά����2�o#�,��jn���Efvw�rÞ>}��Y^��5�f�.��(�F8R�;����� P�B�mU�E�h��E��Eb��T���b�/�Kj[Z�V"�m,Km�F��m�cU�U(��m��CP���S(���iT|���J�ƴUb�-�Kj,Y��F�J��2U�cl���KAڪ-��E�X�+��֑<��<�1j#h�#R�b�m++�Y�YYUX�3�\,E*���fQQ�0�1cQ���,b�˔̵-J�`�Q-�h�UEJ1�����Eb�UA�(��QAAJʉU�9��Ikq(�Z���e�EX"�m-��̘���8�ZV���
%X�[(�-r�h�ڪ�(�őV�ՋkF[)n5�Zも��H�#mkE��Z��YmV
�l�3((��R�*��-B�#+����Zլ�J�ҫFX�F#)Ah�,Eke�	kkhV"���b�%-��-�p���J���Xc��QQ�Q-)U��kJA��~�> �AAMl�*Y�{�1��p����2�v�z�mc��j�(��S4h�9��̊�}������胅���5E�{��]��o���!���6��e�N�Ie��\�ׄ�B"a�-*��˸�R�P�����Ş��>^wΟT��f���E��p[$��]�+�-WX����)��>I�0����yY�T�r�5=.��5m�æ�ϔϜj�J���#TG��!�9a����s�c{��ܴK����j��+~�s�e�S�l��:Pq:��޹����d�������A#"~��f�+�Y���v�%B���"5 �`jf���uT��w(��齹m�ӿ`\b�f�e�a�n㫶"*������j�!>��<&舯L����2�!�9�߇��Ok�JS���"J��F��G�+��n\�D�'���t��\����{��nAY]sUOW؜i�m�=P��]A
�a�G#�Y�x�r�S�����i�BmiuK�[3|�&!�0�9���3z�O*/J�(W�u-*Qo3�}�/�B�DoRM!+�u]����0�P�ܪ���A|9Nj�	���G�R��K�MԴ��G���]�9y\0��n><�,��9��:NrĨ%�0��䐊��o�V�9�����f5(��
�9��ܴ0���W[˹��s~�K���6�%��r[�A���M%��wV_'�.%P"��l���2{lڢP�;���ۗ~��D0�G˚�z��G�M\pԯ��+B��u�Н.��{��.�KR���5��h�,nE0��4lv4��nUǞ��s֎����֬��Z�պYS}}����V�<��4�ȍ%��xs��m���g�KC�^.�F'���SӲ�����=�"�˄!0X�⪡��Uz��2Oz��%Z�v�3ޖ&�!���v*3*eBītN����:��"b 8_z�}廊���͋�\�y]��^X����f�B��V'���(�&u����:�2��K�*���^(Y��c]���x`�J,���(f�C��>�^s9�L�W�2����ʔo�9C�������Zg+��9���l�ԡ�|�*�w�/�@������K�8�zb���I�� �~eﭐ�WA�[����ؙYZS��ش�F�EY�{|;�����<]�䙗K�Jou�4��=��	����kj����HHS#�iGU����wz���{ʮ칳V�(b
%��T�:��y��47v����fJ���3�f�@�W�{�/0�����QQ�M��ӈ֦�!�$�/�����;��u�K�pV��ooV�c�1���XnJn
�W*����#��9�f�c 9�Y�w6J�+�.й���G��n� �L�jf�����Q�ʞ^�T�a���#��_1s��0E�5��^n_+�T4|%�>��.Y���@4�T>�8&���f���Z��n*�#�����C��}�yK��!
;�>J�(�Q0�����i��t����}��p��3�T��1�Z�f�zP���(�%`��3>Wdr�M��S��,�Ye�(^�u�F�;�]7�|r�M҃!>�C�k����@�3��P��Ua��)�so[�����A�-�l���iO/�fS0�K�H��c��h*��x,[1�ꦂ�*^}�w+V��l�sYhR��K�h��x��Z3���C���X ��R��\�����u�|����X�7>�ڮ8��P��=ΌI�t:�>��.긐ۻ�$�^»P��]sGy�`Ya�$'R��e}޳����fJR��Q�����ׯ��}[��4]�I19�ڑ��n�dr�0�W�L��nx��aJ�b�N}].
��P���0�����ܵz}�<���껠�h�n�Ԟh���p�Ҷ�.���Zij�dC�+=@�s"��+��.�X�K��Yٺ��E�=��������gM�+.黇8�Ot�<�8hQ����⣐�zja�)�ȫ�ٮ��u>��#+׌�7�}֍�M@T}p���[%�b�Z~�#P�?q5�n��2����V�l}=�Ƴ��vY�l�YG��68:�q��Iz��A���o�tX�n�ƞ_>�M�>� �購�~ҫV�E��`\_��/:ч3s�ա'Kk�����↠�y�����}�:���w�۳K��Y�ym6�;�i٦��|�g�.N� �{ʦ͓:�d�	K�"���㲠�,�WfD|q��\�>Ɍ{��x� �Yy��c�)�l�b���5g`��S>�gj�Ab��eԬ��S��/�=���]͛7��ñk�5�ˑ�~P8n"�JK�Z=*���BJ�%�Lyٔ�i=��n\�����1�=�ڳ�X�V<�!,6&���Y}h���/��ڒ���[I�tz�yþ}c�kp�=��Ժ��é��.��'&GbZ��^��t�US�=���X�i��D��o�T<��I�`��8{Ʉ��aϦ����
T8VP·���U�#.��KP��.�b�+��;�0�5#�'j��b=��=׋�gC;%z��������'&���0�;'�}g�go9P�k��7��3hB�}�[]�r
Z�j��R��ѱ�wFO�H!��٢���*v�ۊ:o	��r�
�1���Vc���y}[JX�ܱEL嶦תyC��!�jX$s9���	Q��8^�C�8�����y�k�}Xp����&����a�i���`h1;iE��(TU}�����|�����w`$+�"k�M�ja�W�+����%�pn�Q��hJ��{m��B�⊹޵��J�%=^�^��A�,���SJ��	������U��I�\4!~>��4����cf:�S�O>/c=~d�����C�:��,�t3���uҶ�'��h�˥������� �wX��x������7��#7��K\�iS1�)�l���d�<�&TZ�2��d�M�Z����g�=[�x�E묅5m�à�nJ1��N+ڬ�"���/}}�	�*�c�o�����ld���2}咂5 ����=^˧�C�>}3�N<�L�颎��ʮ[�X�K�˼+��ab��mVz��흪_d�q�Pܾ"ԃ����6�k��3���ѯD�)�����.@�=�WJա����U��é����E�����P]`�E^,��ǵ;�}Q������:|j>�����)�6�֋��
3�������q�wx2�A�eL��69�-�L	l��k�1������B���U��n�0���%��I�Wn���pK�WF�|Չ�ۢu�sMN�|蹯s���ޗ\�@�S�$���D7>Q�X���m�ZE�����N�$��Ԟ*��ŏ/Uh���;��3Q������w �U�զ�(��u��{�oVcRB�{���_�o�\2�u^b���	��i�9���}�u����%E�(�=�߁JH�MZr��K�q$w���[+��G��%�9೟	�����n�{6��ru�ݵ؟wEv��[�GH`��5���	O�sQ�☧ܴ�*o^RQ薏}�˯J��[~���"�fO%\�=*�+�l9u�H]�`�L�\l4+�M���ם�`�%�2�<�%�ք�Ҽ]s��`U�U\u�ݖh{�wG�����J_z�.�-6.f�lܭ����f��oV�B�>1&{�X���p�&<UT5��u�,����J���v�o}�5�/b�k��!��{݄Db0r�/8� <�@�K�P�M	�9˼�mo!Bgw�o�C�����)�����{V���ޔ���6�6���C���5�zs�^U�E��2�Wo3��N��ݵ}�[}%\��G$�Y��:�X����B���G�OD��G5�K��I$�h��y;����\,Ar�o�ة���s]�5�	�33����t-�ӝq�KS����Ļx�oO���ղ�q�w�4=��n*�����b���,���ˋ7\O�q��dY+�k��7�U��B��`��j�5��k��S}��<��2��6E�z�PB��[a�x������P��������1\�fiN��y��wC�����W��/}e�x+����+��]�s�~癓W��lO��܂��]�{2��K};c2��iQnxxx��l�Va�L�I����{y�������=Zy�j�g53�a���G֥C��^�>(=6��1��[=�8��Lf�5>>�d�P�/G&{���5c��P�w��&�؏�\�>�N�O͸��0^ߨ�z5]� ֊\��;�}bS�L(:�P�/��,��i�B���=�֩�o��4���
���]��_&�gŜ�6��̩�n��^��'o5x^�o��s�`<[�τ҇�}��\�\�(��@�y[
P*�Q�h.���r;�oV��~��\�-d��+�O.u�|aj�Q"h�P7�S��P��^bكx�~LS�)�ڭ��]�7Z�����Þ�*�s*�m�)X�o�:O7���MY�ltbX֢��YSv��VN�e��M�qs�'U��nٔ�Y/��'�Yv9�Se;*�*�t�\,i����Y+�99Qˌ��4eƪSk�yy�flu6WE�B�:r�׀"��+�[�GY�2����mگ(����ET.�L�]
v�6@�պ������2�G%]^��W	໮���L�s�ck����x�� �7���3�9�Y�th�J��r��SX�}^�L��Y����%���1'������oE/�S�������չV'�60O��!
�Z<3�Jg����c�lC���TIϺ\v��ߪ��XM����dF�@��=Z2DN�>���e��l
B�n�d���f�a��Ok
�TɛNMʷ�����M����8�7�C�߄�Fϧڀ�4�Q���&�Hs؎��[���>���Y^=���gX��Ϧhy�I9���������Z��	�Z�����C�ӟ_n�>�Fz��:��nu��b�a��r!8���e�j�Z��j�޼oA"_m~�ݎS�~]�)\���B.	0p��Pf�fcJei�^פ�G�r�g�(��Ku�۾x��o���`u�),g�%��Q�{J�����Yl�)53!�4��48O��W�f��i��O_!�uN⋾:�T����ss���w K����v:��=Fi�}�N5xw�����ξd�~~9�N.4Mt����1@Ҩ���� %\W���R���Tpw)\U�n�1��t"= �%��;�⧵lb9�^��ύsd�ru>=)�j!�#h类��ҝg�w�b��¡'�:�l�0Q�i~��|�z��jޖ&|\Ok��X�W�q	m�Ʉ�-��:1�o¢E�'�Mͥ�j���96���FW�����9`LRk�R�o[���V�4!Dq&%���o��,��<\f��I#˶���à��Ȋ�*�0	�Jyo=����ycUva�O(w���#x!�y�1��"�'}^�ō�*`�\dEp=t�J���eE|0�xK�=�V���O:�N�������􂲻��΁��~��T;J.��x�#�_y�=~����Y��ɢ	T�S�����:K��V��p���}}yì3���`}�l�<�O�ʚ̧֫���	�g���SJ���Ȭ�l�9�W/E^]��83k�.�|Y��Ɲ�<����g��ܪ�:��	��IdS�!(��\��'�m�}r��eP]��A��=�=�A��ܶ|f�eoK�\��Ҧc�\�;���qͯ�Ѕr���r}�h	&�Z%g�ᱷYn����@q��Y������kkk�Ռ���uyB7' �R�	J��U�g^ꇲm��q4m[�**���q-�0l}͝�0\�^��K��@�2�Vv�1Z�����j�j�������-�]5^*Z�]���ۄNz)�u�1����Q�}���s�9����~ʇ�i�|�6P�(�Vƨ���W\n�G2��ɜ�����Z��S-m�
�jP�ԃ9��cۈl��J�]��%Oc�s��s����ov�{����r���fO'~����v��ܾ"�T^�P��j�{�{L1���W^�NU)2�����L]2�_+V=\�����/x�rWS+��t�;�Q7uۇ�3���O���!�7���d�Fat+.-g���A�傱��mL��qs;R)��K�H�~�r�%�-���u[{c�N6��Cw֕u+��2�_T�����k��&׬n�K��lw�]RbᛱȆ�pS���Df��t����f�|��z���^Q�>�o�B�H��9��D�e�.%W�'��7��lW�wd�K�I���|ѓNx�����Y��&y.D><�e�	O�sV|�Ȧ��?|(ͼ���k���XUێ���7���CiIeâS@æ��9Xara������t���$��	!I��H@�����$�$�	'��$ I?�	!I��$�	'��$ I?�BH@��	!I��B���$�!$ I)	!I�$ I?�	!I�HIO�BH@��B����$����$�H@���d�Md�z�'�~HAe�����vB�������m�  P��� R��l�M6�e��\}���^}���'����TthC;������
���PХ%AI�w`
���|�y>�}����8zt  ���CT�RՓ�n��TQB86
� w� 
      hiT�4      S�mIT�F d`4�b)�g�%P11 224ɑ� S������ �     ��"SJ��@     B �i�i4i�24L�i��f����ǻ�	"S�0�hD�����"�$�~5�.+�ᬑ'��xg����������3�3����ۢ?Ŏ¤[V�	� �*aG"3��{5DI�R6��ܖD�V$D7�|}���������lW����ϻ;����n�Ā�`1 �b��m@�@�@�@�@�@��lP,�	@�l�0�0�0P,P- Y@Y@ A�� �Q�J4I$�-!D$�39�m���n�  1  $즃b�b�b�`��64 �@�lh$��@�� ��oێ8�Q������]#O��bSF�t�3����/±���]��j�^��ӣ�r�p��5b�i����%`�.�ڜ��,�CMZ��N�	ۥ�d�%�RjE}J~��G �u-��*�w)]FX Ɇ.�];q��]�hU��V�&#&���+&$����&��.fҷ7i+(5
�Sn�FL�]H���"��($�? �fD�qw5# \�X�.&,���5�G&`@�W�HC���db8Y�W���C7�@ʸ������V��0T��-�$E;���]ӬJa5ջ�Ǔ7���R�3��@BEd��/ .��&�7NIJn��4��M��6 ���7Y�\UKu��8,кWeCU�F��`ۓ�ve��Eft~yeT��J`B� d���r*B��U�9UY8�\�N/1IF%�2��0أW0���e�E]"�*�!s)@�R��<�).XiQ�0�UDN}�dc�P�2rEI�6�1NU�E%nh;�ʆ*&V9t�V}-�B�*.����X����Y��ri�7m:����#&[�T� FE5`�H�� V>�u�X�Ê�9j��ʱ�J�U&nn^�ٍ��ɓ
	��%���u�G ��%J!�MR�B���*fW.�!1a�v��m��Z�>c�D[%���dLۛTD�Ɇ	h�L(�X�b����t۩r�Y�+g�Y=�9a.\�9C%��P��,p���Q�2��!$�SU�
�PK��JӅ��.��,QC���v�@��(d9i�TCl�i�dӕ2�dZ1J(	!I"-���чI*�jA���T/�����#���:���ݴ�ÄR��M7v;��g���-`��
���7�𨄨�`�F�5=�L��R�1ܷ�Y�I�Yf)�nU��K�b�|� "a>��՘Y�3�C^H nb�����od�B��;6A�oIHOARس��%hF�K����N]]���sJ��e�D�
Z"��[:�]��Ӆ�A���P���@��˥�yr%����ǽi%����yǦX�C�TH�̡U��HdMq6��P ,�A��	�q
�D �D���@Ku 	����D@>��u3�V��yF�"�v����|�'[q���3سP      @         ������     �.��m����'1"�q�xX�0�&j%�i��M�NMU᳒����e�nB���[����ڮZ�b1�,��̲�Mz�e�0����nl��3�q�ӛ��
k�L���v�P;,�8��g&s0=v�#g*�;����T6^NTYK"F�s
���% `nMN��A�ɜ���띵�WS*�ڽK*qU�5����[An
�}�C'�|�O�3��Q�;4T�[V-xp�Ç���?/^Η~:��^���k4���D4t��&7����zD�z�zx6ؒOq�͆,�$r�Đ�G��Y��w8W{z���ƹ�*t��-����d�(U2��o2���&���vv���+W�2 B 
 ,� C� h@k�p�0#%���2�cnW�LP�;h@P ��(�����et\n3�*-�%� `  @D@  �  `a���xj&i��
�g���m��Vť��#��f��A%w10�'�Y�JA�B�M6�A�0 p �
" p 0  ��t�o��QMt�R�ѷ�Y���N�<�t��J��m�h�6���0SR�bo���
!��B t`@�� A� ���)��r~��k�SC� ɍ�>j	���^ѩB�^�$S �3I�Oa8D����	|Hڵ9Yu��� �� 42@�� ( �  E���h>FY�x��6�3�W�����1ʝ�������r���T��,�Ξbiw�h�7
 ( �p  p �� �
 ( �2Dk'6g\h����ÁI��h����V��V��͘�p̪9�ݙ 򾫋�v�yYSq7w�@�( F �  � �
�R�g��v���2�)16�B�L�)�"��f$���0��.����d�Z: @$ 0& `   �ݮ!�g�*e�"f5�Ij�9!X�2��e�r�`��t�
�;}n�6S�EM_\��7�
ĮP�rt�������Z�W-�wU���+³�]Y�OY;"	�eT��؜Q�*��\rf�Li��n1�Y�le���a�}(�T+��+��BqB�L�ʨ*�\��!.рC%�
a$�P�h�a��A@!����K0Ja� ��� �j@JT�ƚ��MqCDD�5Y�X��c�g�e��y�K@țB�h�7,@x-��" �eM֬�nm��6�0D;}-����1u�5>>Nf&Ȍ���3��kZ�\��fb2�Ѷ����u�'3.-[~BY-�KT�0Gd� �І�n a�n[���� �&���}MU�О,�j�-5�5В/1��ާQ��ˮ��n{�Ƴ:�w���[y�<{����,�f����0�����D�F����ܧ0D��y5��3��V.Y=�D�ܷ_L�f�C,�i���+�4�t���LJ�+���iaBJ�V%�%-F˄�kQy�w2���+!EO�R\�����/L�
4�0�&Up��nﵳ����Vlp��V&B.�^�B7���<�ŉ�\D.�[J�jEE����(�(�B�Ԩ�`�� ��	x.�_��!`���j4�!,KbZ.J��zN^$����f�@3�eEVf'M���}�n�i�ٓk�u1L�ZN͙�M�Dx.ߓ�D$�w�K���E�BR$�#E�਄�*�9UU����]��.�.�>��+5eԙ>�K��5ww��M� ���8��T��h�H!a�YN帎�$i�P�tL���	+w�EtZD�D*��rfap��GMvd�A�(�BA�B�H�X�YP�^m���^h���!P>���[-x��Vw)B\#�y;1	tVG�n:Wm9iC��RL�,K�H�E��6���I����.�J0^|iI�+!x+cV(���	����(ޝ�9��w9��SVDt^����ȱxDdG���H���
���dV�!%�Su�OK�����+�zD��g��M�]�y�ۿ����:�̸�I�zk��y8��������3�e�'idB��a�=�D��ٻ�#�uW��F�^��{��H����DQ�L�d+[���V�\8���}�DyC=�Pl�w�tw�Պu\`�-9����2�5�x�[����ŷT�a�K�^�*�����,Y�٬�����,���V�,z��6���?��|����*��$��i���@#(� nX��%�8MD��ܽV,��S܂a_7���k�����#����7���Nff\Bnx��Aq^Uff_	�������Ͳf'Y��n�vv�}
J�~P!ꗒ��i�)D0��v6�q/�x����\a���^�لx&7�}WFjKn��F��EU>��oD@O �c�8��������axI!�7�i��|~����t�Ҭ����j�a�&8C�)إw����{���	WV��ޜ�*�-�O�<��;1g����Qy�}��O
p��'���޼m"�=����ssW�㙚�<t�C�N��%���j�����n���}����������N[s���7q��[c.�v=#�Y`�\eW�ݷ��y{���r�3��x�4���0�&`�E�`䫆ʖ��yj3�ֹ��;�t������}�[�˾��p�����SG+��hT�b��W�x\��D���H�)q���/��\`��B�77��8?Ph�����舵Kb����C�vD%��Q�Q׾��}��Z8mf�U��l��I���L�}"��=��e�^�_DCI��_.F���xȧd���Nw!I�y%��ޏb��-3� �p��,�e9���ggDA3�@dA�^�Tk�o�3X�@��;"'���L�?{[��"�x�jt�
2���B��+�&7~�7{�Y=}��~�&7�F�'֫3���~������LV�]ה���*{�i�S���L��Y��" Fݍ�]���M)*��D�Y[/g.1&���
��إ��W�F ̼��cn��Q���ELh�Gԩˉ1& 8̇
@"��	8I@tx[����K��flN��k��z�X�yb �vd�H���Kv*J�cFw���o��|����!:���.8����<�ˍ	h�wj։i;��q��̸�O=�sG�U�e+E&K"�6��R��/�/˙�r�z�T���?�|�'U7�T��bA8T���+-�4�s�����Hmd��#�9�ߙ$��&��7k�dr�'b��ߗ��DQ)D@@��U&Gs.��B�����m�u���#�E���{���([)����{�~���E�UF�XO����}v���s�﫠߅a>�.�f�zҮ��������y�G�y�g�n�Eo�ߞ��%EgK�ϫ�� 6�q���%��qP���NF	�+p#���o�����
��x͏q�z�=�.���kr���G��,3C>�3L��3�ޟ+PUJ�߬��r��DV\-�V{՗7rr�R�3��p�o�#1�^�G�z�.
=N*w�0Rͬ���DYAz*��]�od0�ּz��K�yr�
����%�8�0Dђ�����$샻��^����������#���zq�b\���{�pB�-z�-�T;+�Ez��9��]���w0����c���m��~�w��.�mz�7�!_EE�t�I"��8_�[R:���������S(𔗩�����}��zc�1άk'q���H�3w6�>3���D>U����&0y�x��q���<l"�Ɂڳ�U��߄Ǚ�3Sn5��w�:㼬��k�5��^yy�g��Y��772��#��Tqud����q;�Qe%W�-ټ3' Lҹ#|�z��c���q��U熚 �t�\i��T�%��<Ȓ�-��@�ȴoe�ꮎ��2T�SjL^d]�F�e�Il��ܳf/^��Gϝ�sJa��u�׶Z0��,F�^ �@�� VfH���Ht�UY7�ơ�����K���.�h7q�Yy���h.2s31��n�k33333�UTׯ^��9��#T���:��*�,��ةa]c�8bpy	*yx_�Z�G�0�������G��t�NH`�>�Nm�R���o�#z]�{�U(���y\��^yߕ��W4��\���º-K���V
��7]�HH�a�zG#��$�:8�YY��DV]H|2va"`�02��ߛ�z�w�g}k"�Ϊ߲�<K7;є�6[i��X�%�{mm�+�o;T��/A#���P�/���
��q�n^v��< �h)ǗLN�Nz^O��%.m�����b��ɪ���D�L^�n��i�?2��^f�!�b�R�;! K�K�T�ݝ|���}���K�jf��U�\�g���i�G���m�z��N��o˕�x���BI�Us**�]�櫷g/v��x�^�L�[s�(��VjKO32�OO��5VA;++��|�����h�ٚb��N@�6����}�S�)���x��"ݔ��cvN�z��f��N���aU­��p�/��/m�щ�]z���|s�s��n�zN�/�Z��\�$୉Foo-G����l�+PY�30��i=kՎ~�o�Df^]�fcEc;X��R|ҩ+��=�L�;�:�����D
|�l�5ӤtO���Fe\��}x������ʄ�D�#�>��(�\��uw4>&��#a�V$�Or=/�n��źdm�u�g5�acz��ƻ��ü�f[ٽ�Ӏ�9����tQ��?J4N�(R��Y�{ˎ���4���[bXeE�^n [� f��U�u/������`щ�����W���@���&�/7q9U��p�Pk|fV�3|$���3+Y���WU��菊�������^ǏOV��wDE�{����й������oRF��'և�Nľi���3ew�>���[����
k"w��}# �%�������\ e����b�WD�ȅ��P� 3^��M��sݷ�7;+my�w��|�#�AQ�m6QG�����$��^���"	�K�w}�2�nl*�+����'&�!����.)� WC<H�N�P�F\�smx�68���>w����W����ز|A&1��+�&ξB��{��U԰/�I�'���� ��]�� ]��no/=����}�{��(�$	���0��׏���C�<�i)��^'�H�B��x�-�[.W5��X;��Y��fi�~�w���a�~�}b��V]ם�YP�beVy
 �5�Ҩ�/=�^>��|����{�@+���'������צpLƦ�Bgp�0��^�6R\Ur�I�󆏔oC�N��i�yEW?])|�Ϧ���
'��~���yX���Z#����J�����9�״�K�}��#7\��,�\8=9�D��E����k5׵�+���:�D/BP��"$��!  H@3sl+�+��e��c<!,"�>_��7�~:&�X@ǥP2oO�S�O�.=�ٺ�{B�q���v�p�Çr9�[%�j[Ql-Fw:>Y�U�,��m^ݤ�c�`ī�o�4��T���:w���њ�p ٴ�n">����L�پX&����(��	�(7{7+!�ع��wce�*n%�ܩ7�CeM5wzB�S5��.e�Z�n�^*j.�wP"�!/5 &c�T�R�C,l��c���GZ���]osyZ��n
�����Pmroc{�]������θ�^ym�����lZ��R�M��|��)O�p�W���Q�D �0{���&���*����Ѯ'֬�����߄���`��lUe^t���Q	@����P�Q�z���W~�*��\�B�c��x��򩙥>.E@p9�W{��؄
gq)�/aJ�����|�G����;�z@D P�(Wk��l/ߒ���?�U*IZp�P�/2��Ը�ܸ][0��rg��xޛ���b�/�
g]������ � �~Za�o��H���~#l/�ȏU��=��s,K�[Xm��;�U�9�����O��{�s겋�ʼ�������ۥ�>��ʢϨ��s�;���j4篓#٪��x��QuqE�r%)�f7��>w������   ���`�˞!_�{C�~<|�Oq��:΀���8��A��^�I��0�\g�_�E�E��	n��v�G߄! 	s�ܢ��R���s>���]��҇v�w���	jϤ�3���ɲ;k=�:b7�3b�����ԋsW;�/@  @	$�K]�����eTxJ����)����ێ'�߇9.(�Î$.z��O�E1�my�F�q�j�U�UV�w���}B�D@�$�@D�;�z[�.�A<��*�k�;��k��ڥ�c��I*�U��ޗ�ݖ�`��xuv�.��������zHpߢ���-?f�&p�M;��9��xXqޗ�m�u	�����*Q���[ٖd(������EzV��ug���S�ˆ�n�gQJ�r-	n62�EU��"Y*������1�^F�k�\��������Q@�\6Ғ�惐!�d0͉���!Jb�ɗ�*u`��Q/��}�35s+@Tbe� 5��
��ћ�Ms��Z��������ך���Y��n�n�զ��u���IX�M���In���gkwu`����݅�X��@	�����J��H0�����^o�@  @�i�Z������ed�8kҜ����K�Li�pD�[�AB��m0��rX9W�D��ou9]f*on��	(W��[�*X^0�ܬv�m~�N���f�<*`ǇѬ�V�n��F-|�g�Q��{+v��x    k:���y�w�j��2!�����r]y�n��={Lu�9�+oM�ȼa�< G��ڮχ�Ҙ���o=�]}��� �>nϿ`1I/��7��/���M�O��g]p�`E-�Uw�WE��J7�Gm���.Z���QC���}���@ �\J������~�:a�c��UC��9-p��q7~I^Ӂ���ƹ�$Z�v���O�z'�|�ۉ�޽���� @  ��^����{�~�<���\��A�c||��{.*�$p����3�,�L�ݱ�59��FzEJsy����    ��(��Q��~-y��V���ފ��=N|&N��ueU�3NևV���ô�+f��\g�]\��w�  @� �nt�;*�Hx���(��K�3|�ygA��W�X�ܻ�a��H�S�W�Ӄ>Auq��,A��Veno�� ��\�G��%~Ô�N��i���7FN���р��(��J.qp�3-A�=>^7�R�����1�67��el��n���  -��h7�'u�
���c�%���|͍�I�OdPF��f%s�+7��\��`����k.�U�U��~q�n��Y���oj�:���-�ی�(���%5�3��Rd�e��s*�e�d�͠U��N�1yi�L����*�2� 6=�C�Zδ75a2m@�`������77y��5�H{[���ZXC!S���ō0 I��ՔᷛOowlc C��wuaB����l����
)�!�%�kwu*�%8!	�I72�D	5-�i�����<�<�� ����x	��)^��3���Xi�/�H	�\xB�h�l���i�H�����|n�ɗ���ŉ�}�M}/���t��|F�^�Ѭ��J�8�T�	�Fg�6�f9�7�d��Tt�����W �������QY;}ۿď�z���<ȪQ{b�$͌�άB�-�¨ܪy�9ƚB|aB�N'�o�Ov/F?�x��Tt�/r���w�y{�����Sotv�s���,��X��j�:�<\������}��
���ǉ�w��˷�x�z։�g7:5��ޓ��޽߆�"���U~f�zp=�GW��ʊ����ޏ�����nYim�jG����w�>x���@������j	�P#tO�&�y�cq>�팹>�XO�?�҉��u�g@@$O1�+5P�׋i�~t�D0�uy��S~���1��g����w��F��qq�����<�^_B  /;Ѣn�5*���Ϋ��;VmR��n�|ј#��yR�wlկ� ���\Ufu ��ĸ7c��"Џ�U�����a��;ڨ�t��%�z$Y� �]�m۫�΢sW�KlEi&F�?$�$��z���}���e�򭉆��
i�S�� 2��K��<�Q�b�殮�<�(V+���Pb�}�l{ݻS����T�L�F�5$��=��r���BL�I�l���\ ��ƜO]?�'l���ll�/2V!�#$u�J��B��b@��Rf9$S��܍,ݹ]X�О��]��6ؚi�N*��ڽb@��� �����woD -��F6�ٳ5��z lm�;��W�"Zn�6������āhco'J�ݽ@1�&�� ���ۆl����c i����&�f���{�ōJ$abm��6�!lM8m��/om�( �AK��%�	��m��Q4�9w[�������M^��R�/�[�j��J���0��6j�M�Z��N7�j�H���͟v\��f���4���^�gL%�V�N��o�,>^l�2�OOc/6y��&Y<��.%���y��->���1�E׺[�S��S�c��w��������;�u�nD��7�;�j�Ս�m�����(9u���@��\�j�B���	 �=��T�?uū���M��O��W���|��zU���g"�<\��!�뇐P$Pcx�_b��W-:n�pS��+�Wo�:p!�9��9�[��GV��*r9����~]J���m9��؝�t��]!%���ni��]� ���s+�;�:�uO�������<��xU�����
�	���S���?GA7D����]�#��1*9�3�f��}i���J黣w�pb� �\����/%I�.����y�u�N�8v�w�$���zV4F�z��H�k�:�VcY�9��Ĉ�gC��;+2��;^��z�6C>}�Ϯ��rfL��Sqm�L��#�"cʊsQ�ҥ=��2�:3�!S�wp�6E\��0L�8�V=�A���gi����rM�׌�sr��Y�=�ԢMҟ��T�^�f���E�R�@F�ā����&I�V��dQ�β�Ӟ+��M������ԅ����ci5�kwu," �wwU� �l"*�wab,!N��Ƙ��iU��� �����@���ǵ5����"�;�����ơЎ����S9&e�/��t���&���j�P�^�q����鉆�������y��,�e����֊o/���}��f�.ȯ*�SI����C(�8�[��V�5?zu�*��Wf��aY-k���lVzz��wt��8���<�B��w^��e����q�ƍ�.a^���a���~��ϝ�뇛uJq�\�!XcO�>c=���b����,����v5uZդ;��4���d��y�j�đ�u�[�η(Ɂ3�����]���s����͉�q�T�K��o+��|�@���$�5+��&|��}@�O���ʕKZA�~���"'ߦ�4i��9q#'M�wQ��u�W�� �Le�ytYl�su���n�*o�/�C���	���yL�n^lc��e����>�����빍�Uj�-���y����VN�9���\f��O-~�)3�}����/����{9I�1���ٕ�_xk�=^�J�fW	�~�L�٫���v��wYy��:,���4. ��~������}�+E����⌥��+�U���ѳ���x��=�`�^���Ńm��[�`BD�a��$B_Ԍ'"�i��%��c�hd��-���a�t��l~��I��p���L,��EN!�Pe��$�	�2��I��D�F$L``��L01ޡ�\h�ќ͵a������U��*�QV�Ъ*�(��(��(�.�0,���`��)EQE(��(��Y(�E(����UQb�(YE(�)E�R�(��QJE[mr2I�f�#�����5�"�r�4�an:`k�	0�F$�m��v\���KaJ�Ũ��wR^,u�㻆�v��G~�bƆ�jp1�2���MZ���JC�Ä@x���q���`24��J9�[��77X�ф��9�Ʀ��m�8H�������s�:x��_�I����I$!��M�wԂD��B�b&S�=�t�'6�����!܋�k'=#���~��y<���q�v�rIp�}rA"o;��R>y����=�eڼj48"�ݤ�7=m�5To�&��� �ō,z�����<a�XL5j�Lcf[��������]ׯ���y���e��)��bH�+��f')c^,��kX��+H`��kH��u�%�[
o��Q�8��-��l��`���}���ɫ��o�f��m���h��ܑt���Ce0�F(��\�XJQ�sc�}�����v��{���kf��>�[��;�ֱ�u��(v���d���^d��F懛����~3��#o�oRT�!"j�I�gaޘ�����G�W�:��[40�k�mۆGř�W�������n����[�d�M�j��z�}�H��]�{���{>��{��H��k�d�D��˓��┧���5M�U_��>�ӽ,�$[ۭ�D�d�	�i��c�]_;#�X��̍��2tj���o5�:5�⍝2��l�C����b��fc&�IO���+lT�$LIbjĚ��x�ȝ�A�&�wyUr���aX���`y��I4۝�Q�����Y3S�q����o�������BD��':��c�s��D�� �1�_�֓���S�d��Dyx�O/��ڻS�;]|#�'�:W��4��BG��zd����US/<{^���t<��c���&�8�|�~�?�è�>��a �<^�߫n�}�U*��L �|>�p�=�����F�a[�_y�C��rvs?Y�����;�2�|�wqF��)M�Y�����Ud�I��u��0�v�kG���s��#ro{dp�5d�_��n�����ɪpL���޺������x�Ѝ��K\�.�{��q<[�K
{�U��NGc^d��9�a2�X��-�w�5F�sʾ6ǯp��9c�ĲI�X>s3�2>�B9q�#ү��~OD���z�����zOh�S��=^�&ƺ˱����~~���g:�H�e|pb#�)~����s����"�(H�D� 