BZh91AY&SY�I��_�@q���'� ����bD^��   �>j�Jm�h�IQ�lkII6�T �
�� m�P�����
 �lm��V����-��lV�2��AL�T�ثf*Yl�=qEV�*!R��l�-���62��D�&�BkQ��Ҳ�
V�!J+h�*�R�m���Fl�EU6d�4+5��MNwUv�L�`"�I-%��h��4����V��Q�lԕT�V�M�D�bFZR��5�H"�h6�iQ60IR��R�9��%Sf��0�   ܓ첄=��k���Z :4ցj�*��Y�\�j���7j%R�� +�k�U�Q�gE:�i�q�X�_v�U �dْ�TmU`�/� :��Ǫ@��wJ��;�p*�*�W�P�N�J
��r0ꄨ]�s@HPWn5�J�n� �R ��ꃠ�wG��jՅU�ͶUCZ�4|   վt�m`�.�  ��qp7aAJ��xv �{�Р�^}����O=��@ m���@=h�K�� zR�ҷ��
�ҏru����@Z�,��V�<   �`�cI����q�`S@7����(S�C�v{�(R�.sA� oU��
�={� ���  	���]m��YA%"�����X̰��   w�PH�h� ((��r�eӀڗU��UJ� ˎ�JU�un )g�*� �t�С���顖ʖ�kf�Z����dπ  ��z R����P9³�]��t� �Å:��X�f������d+�M�R�:�t��րu0 }�W��F��QM�����i�� g|r����t �:� �� :+n��e 8q��t]β\�F�v%�E��(4}�z��[T�l�mI61"د� ��4�t�̘ ��  uc@ �+ �� [t� ���@Q���h�E�i�(�M��EV���<  v�� �3p
Krp n��Eӎ
 �)��J�;�@�
����  f
t՛m���T��m�J�  nx( Z�p(*��V  v�8���2��F��78 k�qTG7  �]pR�>   
� j`�J�bh` 	�` CB)�4b���hz@h �� ��d)*R       j��@��T0 �20  & �E!H��0������6�Ѡd�h��A'�J��Ԓ�A�=G�  L�@6�7�+j��{�eiˍ1p�Z�u�+8�m4)�/c���m[,,`�ny��   {�����[l������kUm��mUV�q�x���?#�{�}9��>�����>}�j������[��6�5����>~\�XT���v�.L��O�k_㕯�������[�m��k|�[�k�*�3[|�[�mo�j�f�����+|ʙ�|�k�V�ek�V�ek�V�e��5��~���+]�W̶�f��-��Z����ھe[��|�k�|ݭ|�k���־ek�V�e�����k�V�e[�m_3Z����5����f��-��W�[|ʷ��o�j����j��W�-_2��Z�e^��3j�����|ͫ�Z�e��-_y�����U�5^�7Z�f��j�f��6���j���m[��m[���W�5���5k�[_���|�V�̭k|ʶ���U�9V��-����Z�2֭�*�}e���m[�m��2խ�6�o�mk|Ͷ���Z�̪��5��2�k�m�e��̫V��j��[m���j�e�U�-���mmW�ժf�m�-m�̵�_2�������m���kko�j�|ʶ��m����W̭���j��mj��kV�e�m�5Z��[~2֭�6��̵U|�V��V�e�󖯙j��ݖ����Z��_2��-_2��-_3j���V�eWf�f��-_2����̫|ʷ��_2�����i��̭|ͫ�m��k|ʷ�վf��-��̶�3k{*�2��߯��6�����B�����pKR*£F�T�@�[�yJ����Ѵ�Y�N,`���=Hc����/�QИ�Yļ�RK�B��Av3��V�Z��(�n ηZ4�Y���,��Z������M��n-���$�^X��X�E-�)��80Ʉ�i0Fec� ���A㖍�V�+-�`����۫��n�{	pF3Yc@�Kv�6&��f��Չb{��4��gu��p7[B��T𵴞&��O��8J�"u��M��w���.e��6֊�qЩ%�e��Xú�e�e�V(�5�����M�B���N�b��EX���j�pL�*
M��Ǖ�̦-YJ�l���Q���SqT���B��7.�`�
z�I�d��T��s3;r��/pm�ͨb,�h�1)
�h��.~ph��ܗ1�i��e g죘�b�;љWY�����3#CC���x�7.�ZI�f�9%#� *[�T;H�[�@��xT��K4��=�*����1��Ulջ'�rf��f�s&e��(�Ԩ pR�:j�޴�뮼�e�j��������Z�L�kDo�:�mmЭ��̊4�cu�j�@-A�F��b��V��͖�٫�I̢�`���	-��B�r�*ح�VJ���M���r^�,g�Y��Y7T�"2���q�l�I�4���螕��J��K��t�Ι�������4p}n�6)��}�%�:�4��s
c�=#ܼ�'r�J�ː�4o�i��v�%9.�;�鉲���`��q�ɐM7��LN��{�,Ҧi���Z�р�R꒷m�2�=Q��3wIxvhj٬w&m�+F�M
���n�Ư�l�9����9�[S2�v�c��nY��0��yH��kk-�J2�q,��BYM�x�"��5֨I�i�5YB�ƶ,��:Oj��5�C��kC�0]��A�U���y�5Ğ�X:���[��#q/ہ�Sw"�������7�ۙH�V���6����;-�U�l����/X,A�)dѺm��V߳"ֻ^y\��2.b�Yl�-���e��ժMad�f���Pz�t݅&����uj�����WX63Zv�T�W�A��[��Cg
[!˽K��bj�Km�tB��<�a��ض�o�5���P �y�M�Yujj�a�DǷ���P��a�w!��n',T�w��ZN&�[��QI��H�y�6m6�4��7,��Tͼ��Z�v/
B
)?fl�Yb�	���2ƌ܏]^��.槩\�o����8���6\����*ɣM�f���Rʢ�/X��9<x��h����8�[J��lNQ����N(�o+B��1��j�a�B �\�͢�L�X��k+`t����`��p�*��'6���|8&��+i��Q�<h7E�NUݑ`����n魃X�4�]JYTĚM""��Z�����*��Z�;�jm�7q��4��ܛjd��2����l*�qc�e�̸4:6�b�Ed6�["�L������e]����[�,]
j=u��h�e��j��Xݬ�lx,��oT$Tp�������ܩ����3����Om�Q^��9J�l���.H��w�O�]a�Ƌ��o	 RֳWX�`;��4�ێU���=	m[�ee-W)���a�u0n�^�L,P�C�QV6�ܗu4��%���K%nL�P���W�:�k�i�JCO\��:���nfjN����;w��<�J�X���*�Rə̱k"H�����1a��3=���j��/5-j�6)���{s^eԬUf���J�� :[yM�Ѡh��^�Ѝ;����{�Xnm�{�d��M��om'��wN�k�{�$7��ֱZ��ab��WQ�������7XJ]��Xk2�TƝ�y&:��"T�)�!)"5��Z����ш���ש"���KD��z��Dm����xe�I{Z[��˺�{�ġ#����{YA-ǚ��I*��Ը�͵�I;�rV]��f��G%����mV���&Vhu۹��A7�K��q�M'�;M�xIU�#���Qlਗ਼�#{������0��B7÷�E
�G0aܵR�NHS���7{���at4�Iȑ��m��c�Qم�T3F�.�șZ�hV��0:�.�+f�)�NM��K"�R��O(^a0Cl�S<ʺ(��}u�5j�,�ŉU�.�b��X]��J[d��Z2�"x�e�U%�6�
�T��/"[��!�e^�W��^�(^h�5��!9�]'��K��źik��6����J�J�X1,-�M�o\�.,��$�"р�Kq�Q�6����0�(�䫕�T��u�١���to��Um�*BL֝]�Ѷ����gs$��3Vjm=t�B�x.γ$`����жqEO6SK)®S�򱗚3&I@�q� ��ne�������G[��`U�i��l<��r@qɁޠ�g��m�u ʵ��č���-7�,�Mn��x�P̴2!Q��T�n�"c�la*�M6z!�#Dv�*�/-�ecx�7˱���m�x6H����\�{gV+��d�=%Ǥl��i��m�h����r�5����B�Y!�hW�Z�@�4�n*�m%J�n�n-:�m��y��D@���*�Q�N,�"BN�S�g1ޘ�Ǭ�Uw��r�:rV3��6��oc,`�6aUi�5�ߖ�#Ӡ;Xtl�@h�&�򒞕4A�{�=�Cӭ�n
�O|��dڕ.�bL�yqx{EX��w�M��	S穮v����-�S�W$Z�@]Mڣ{,И׵���Eg1*�y�.m[���4Jx!I�60A���ѹ:*��W~���MP�����5�F�6�vҤ�`��W/�8��X�*�f�qn�2�"��Vaѷ���"�2n�E�K/VPl�.ƺ�c�ĳs㏂z��튞/te͍ŵx�;X�q� ;yF�M���Ԙ��BJ����ìŊ�v�cD�NZT�=*����z���^cʋ!z�iX{2fIg�
z*G�Z������(]Z! �R5�l��/Te�
��4&�!�����r�^K���ʙ��@yH���f�B�uX�SU�M{q9�`�[�~�$1S@�l5����]��U4���N�iR�#2R��r��+Zɹm舰�.�އ6�iU��.�ٽTuF�y�T����-6����	\������L�V(k���#����h5��k�;��;��� ��y�(�tYEU��(Ò̼�-�qfI��{t�T������ݔ���6Dy�)�S�H�E���� >9�G���w�Jh���sq�Y���*T�cd�v*$�tN�]��kՋr�!`�����݀g�o�T�@�kE3�X�Lَ<YR�^Go^��e�f�Ȧ;J�h���8ު�'r^�/�	.�[ƫ1�E;�D��R g�ܔn@�5;����S��{g,���#6:;+BhS���-A�Z�XdLF�Y�[��-l'zK0�+)�te��'���v՘Խde�l�͵s),V�R�
�tb��Q�{`y*苡��0V6Z.�wQO94�����[�3f��*�0?46�.���j;��C�	g�oN��"0އ6�-�D�ɨ�x�U����nM����9�ַ��/��J��5x���m7�7L��LS��P�Y�
�ק#���#6�7Fjj��:�z&���wCF�9����Q�o\Wy1P�ӥVѴϖ�WRŭw����~'��b*�uQ�X�7j=�Y� �pm�e^�Fo)��\l��p٤���Y%�����b5r��fV�i�2X�BQ��a��t�1�Kv�Cb'p������L[C.	m����XR~r��tN���h��F�fK�e�T��2��e�j��H�]�����٨֬�C���se눰�*���۬ծ�A��+b�h�3r&���f+��N�m���R�XJ	��H�ڬ�bO��6Hs(�A�ԑMpcX���-��e'�����tg��X=��NcI�G����hu��ۺ{x��w`��F����C�Sb���I��mRk��Ax�^����de,ʌ
���1
�(T���c�������eᰱ���NVIo��=�<1�8�>F�vV�L���U|rm�bB�9�Fz�N$�}c1�2ae$*���1�f���`�е��!x����]�n�]	)�V�.��.��4m[mOv��x�`��-ؖqH�3v�e �ٸ5'���C�pJR�G2�:9$ �rYٗ�q�BF���fk�
p'Wl�.����)h��c�+m�x����mٖ��*��r�֕4YB�T�B^�gqa���4]kO�[���}�YfP�s7��,�����L�߶��A�n��I����ki���e�?lÂ�6�J�	l���$��Q�W��
�=�Ki�##�]��#1�l]��6N�C9oc���Yz�<uP�L��ɋ�F
2C����ȭI�Y�����i�f�[�lr��`Ɔ�Rْ��kX�6���!nB�/ajT�:��ͦ[C]S�b����y%'�!y�!�Ԙk	�%GQ��Cj���Nձ�&\ &h�"B�]٧����Zˬ�M�,���p�4*�Ұn�˭+SF=�˔�m��r�$Q��p+�o!� O#��uX8Pש*��׋Lm�ĩ�T&Ԏb�
2��2���A`R�ô��z��֮³�Xa�hV���]-���<hQ��Dkv�&&��7�-���0�#j�̕M��n�+��w�8��Z��x��
� �M�q^�����(��+O�HjM�4[$7�����]��J� ��E�Y���]�6����,
��Slf
բ�e��nb,�`e���F<�7��1WP�4��Z�&�E(m�VZwPGZEW����w��i���Čc�轆�li5O���%K�~�cF��	"�j�'faIVR83xcoڪܚ����qY��8�R�ׄ�%d��5F�fwC�%a��dý���: �.=ۮ��Q�lp�T�����D�k7�LmRuy륀қ�f�f�U��s���tJ���c��P�:�*�xU�h�n���n����M�Wa�*F-3e$���"%�z%k
�����1�((��eK�kR箴u�)>[A�*�](q��D3�P�l���t�d!�=3#�Ql���k&^R&�3X5��5ƴ탹�.� %�����Ѻm�u��U�����l�Yg��;N3�����6w�u����X�F�b&0F��0��ǳ]�.m�v�;��k:�w%իBL�c�t����9�n��GSJ�@���7S�����n�����p�{J�A��bv30cF3n���:�c�Z��$%"W��\�
�f�e�ZJ�Iԛ1��m�bș T�E����f4��b��,P�l�AAs%��l1k��Ӱ�h��BjD�^H��G����4�F�$^i�l^^ޖ)�z�4X�N����@���fVc���2`�
��dPrMZ�e��;�VGYR�ɴ�哉Q{�J ��]��E�x+h�na���\M���٘#nݻ7h1B��@K�ШÛGP��zѰst��*=��ȶ��(neِCm������cE������ɲ�ڵ�8r9���vh��ʂ�X�٣E9�^�ZR݌�7�wc��5��"�֭����w��MeZ	���)lX.{_���˩�P�R�N�S�6e�O�w%���s\ZV���0X��F�e#�X�I�K/ڸ�m���(���j
�ZM���e�oX5	3W3Ư��ۨ:f�,�����>���]�zt�Ԇ�@lsm�yj�E�*CiL�Xi9�x�f"��nT&��I�N�-���`���Wd����ۖEܣ'�Sw7,Ԍn܎��
$�Z6�f��zq�b+x5�˸R=eD�i�WYV���463V�������㕲f��sF3M�`*Ln^���(ln����z��{z@j�{lQMl��	gEc�v�Y�(Z��zM*n]�LS�@�ԽJ��W��M�I�p�5�/L�4y*�^�ޠ��"�DlЃb�0�N *�����
2��[�nmf8awdA�l��"�_�	��*��惂�曷���E$2lԔ$a���ʷ(��̔�2&'q�5y�G0-iŷ�}o1�L�D"�J:x
�����v�H�\��2lˬL���i�Zw�A$6uVT�X+y��i���;­%����{�W6ܽ�Ď��ĖV��k%���!Г`���4��2MQ�Jw�V����ݿ\��Mx,]��Tr0ذaŒ���06F�Oo-X�+�m�R�ǲ�2��	��9���S&�N�&#hһKM�W��<�ˑ4�\���E(0��0���ɲ�Z͕�����;t{u��)���65��xo��<�ލ�r�{�Vj�of����V�*�
.�B��j�mI�+}�O"5���*:.T��V^ʈSZ��
0m.�Dְ�2-�����a��)J֪���cViSY�GFå,Jw�<ݠ�ҭt�h�bkM�00ݍ+t��Xr;jJ���@���������hi�B٥�f�:&�J��%1BV6�d�p&�f|�S�K�6w�R���]\����O�R)i��tYl	�t�H�@�t].��m�x�$�|�i���\�W��}�E�oG3$��n�9\�z&�*C���[Ȼd�/�F����9��V4>�~�`<�J��
�l��Px9�tv��L�x���BȽ8���@@	�9QK" v��iή��Eܘ�R�B�sm�R�����aV�c3m�@&�S��' �E��3@gf�Y��X�̣�4g���J◚ejW?�;?ۯ:�~���6�]\��m�5�����O�,�9����:)(L��ǹ���仩�z�|����	p��(�Ӻ}�.�m����S��do�\yZ��`Փ#s \ytu��7��9s�)U�[TvXr��WE��йkՔa��ԝ����B2 �N�2c�ҩ�=I�h��`R��ۄ�[�2�tX㔺���yB%\*k�cCS@Q.��hڽ�6s��zF.���+$�&����9���k-V���쾲J��;dBW=klR�=����әV��U��[^�{�eY)�t�����^t�O-�sv�ZK��:��lV�t%�vuB1�2:r����e����$�Y�-��FT�]�����l���*���صy��&�T ��֖>s��G�2�`�n�����;���Gq;����!]����y�܃9L+�9���9mf֍2�㣉ؠ�YkG���ר���3�����5W��l�����|J���D⫤��fm�G��`��zF�t޽�K��jgQp:�]��hu4�r�a��iJQY�����oF�k��oq��גCn�l��wy(ӓ�6����'�
�:̫��>�6��˜[�{�e��eh0Zަ��jI���No5@d ���;��ⲱ:y�S:v��9������#ndJ��ӆ�c��b�,q�q��@b٫]%����E�ٙg�ةK�-nFc��jȴ��N�ܸɘndY�R�!���ps8�a��5�u�o���E�3n��+��gr�.�n"�k�E�hYW��N���zU��޶m�Db�1����mN������
uk%��͓y��<D�Ӷ��~趐zN奈� �|��d���Q���޳�k]��L�m&�p�Mp�Gޗ�d}�T䃗���V��u��'�L���,�@�B�˹�8TL@�)�zlG�F�3n�)�Ln��Wy<5^c��Ŋg����t�͏"�Vזޅϭ�J�)Ճϳ�ɏ�K��Y��?w�Vڄkvox��Wd���X7i�p���U���'C�γo�\ֱ+P*����}J�6p�ѧ ww�)uY����[�c1� 4D�K� ƀ'FE�$3S��|�ۄ;�ɨf��Y9���^��W�GD�T�ll�F"Y�\]ۙ8��\���g�fs��9f������gL���'��%�|�saI/�M���,(U�L6�t�5ų�%Χ�r­=s2�L�]��_�^jyj<Y�^�BP�v����GF��]�!�N�ڔnn˰�B.�\��Se��+BbÝԵ���2���"U6�v�U��������ҾeYg�nc���nz�a�!�ξ���� �C%SG����| T{������>�Ι�H����k��t��l.�#��7Nʷ���e�]�3�r˘�BK	ݡx����1��K�-����[����kF�nZ�.�su��}����euK��#��YX�;�ڥ�VL���QƞN���6�na%��X1�/g	f�n�&`�;Q�훬��Q�Wr72����ADd�7���,�F�g8�j_A�IKS��YO�Z�;�O�����^�5u���h6\ou]:�*����u�=�!f�8\p�좕%}�����[�2Xx�����w�(�b_]3E����(
ytoy����Г�M���M-#�����m��vUJQ�Rt�,��ޣ�1��
���tT�H\�eʺ&J�|��;`cU;�:��fe�YȔ�+�_'�OjSw)��v�SLz����L�����2�OJs4@xW4��x�J��D�<.���|L�����DM(
�_�K�1�n��FD&�K5��{N���-염4,`�+��?���#f�ˆ��`��/�2�`x9�b�&��`��v�f�����k//]^6;�)�@@�;��X_V�ݝ�����C;C��� �U�4)�KO3p����V��X!֖	z�A��D������u'g<g;&�쇀��J+��n<]�n�F�ǢY*2�%��j�Y�t;޹G��
w=�������r�'��/�].�C���@u,�8Y֌B��k�^W,�y����1L�Zd�܈�p�B���yS ��ڏ#�Qˀ%�w5<��������e�j��]��9�ܺᵄW5��W-'�.� ι�-]��:���f���:����l���Gw�6���M����fz�ŭ��X������}���hZ�҉�N!�$6���88bA�u
;�yy�7r���6#kI�\z! ������+%T��;�Oz�mnF�̐�NwQf�)�z��ob�zun+Y˳$��S���y��7��X\C�z�ݙ�܆[�λ7_i�����ae�� f�:�L�X�Vq����٨��3Q�X��Co�������]h����Q5�b�;��C�;.R��g�u�6p�o0��ೢ���df�����^�ʕ�hӡ��/�3w��6����]s\����^v����� ]����͡�mN�:����K�/��ŕϳ�mJ@i��!��N���qS�����m;ZՋ�M:oN��	Fv����L�Y7oI]���v���c�aV�%Ǚ��	v���Wk5����s��vk��bF&]�9�iݩ�y���\qI=��|P�Y�s����LJa�{\zo,o!2u�픊��VJ��i�݌-�ғGƏX}1;�t]�c��;��$��g[�����:�y���;���OwOб�"�������y6X��b.��invj4{#7���
�+@#�:����<�%�����لҬՐ%Tq�y�)�	��!�ۦs�rgcs�۰���.ԡV5,bJ�2cw7�E���c��]kԑ�Rd{#�L�,)"�Nl!9+���ش�q�ޖ
��0}\��
S�ۢ\8;}ǃ�9�+0-2*�����M�8����Tʙ�hO���a[ې�c����z��Ε�+�gc��͗"��ԃ��]��-wy�trٽ�ǚ�Qz��2���F(�Q���݆w��ɝ��2yt���4
�e��d��@6��Y�M�YĚ٢Y���3cBP��I�㔴�F��1�%)2h,^��q�t�Eg/�0k�OE�4Q��C�����+� ��t;3�����6�����.wtvy�ut��\^�%�Xtǎg��݆,3��[t�M:��jue�0�cr���:`���$"�/A|������i��.o(%$koQ�#�֩��4aO*r�4��y�.�0���u%*Pܜ»�P@�ˉ��Җ��}ZR�+�cB}4n��l��^��o��f���*�xs��hGy�(���ʚ��f��K
J,��ވ������R����7c��ū����h5�;m��\�v�;��[��ttV�#��X��o�$�ڣ:ឺ����˨����{�B�N�#{�˳9ΧC{o�uP;OL0ai�� ��Z�`�D�Վ�X�*�F�G�� eӣp>�4����.[����g�� �Ji�o��&�Z��������/�����}jފGosS�q�,�"��bg+��*]Cޔ�f������
]T�+�e 6�=mb�}.DXH��ޖ���fVM��9Ϙ�+b�,�(�Y�mZZ1]�fB�N��'ooi�P]Jlu�`���	o��tǕ;+�g�)坷���o'�ŵ��Rթ�>(��C�1�!,�U{�e`��t��85�j.2�f�ս�&b�]���6Dfb�����Gm	1Pҝ������.թ߱��[ˈ����n�);4Jk����:��d�os���ɘ��y\��n	s{c��&q��Tխ _3��h�nqT1���.�Z�rƏ+��9V�^y��
N��A��m������c*媊#7��\��lqEY��uVܝb�4-���Y4�͹������|�gz���G�;��]Nhk�c�h�i���漭�/o4h�����1���7�dV��E��:Fs2��p
�Rblre��SCm�a�XO|���5��(�[���>`��锈����+T�>���f���[�8�A���X�'���-(3xpj(VVYrs/�tná(ܥ�䧡�m��Xc��)�����	�{�nʕ�����gs]y���l� �S2��z�\#6�n��f���i��y�9ܵ6�U�n�X���o�������e�N���O^Yvǻ[�sv��A���ܛL*{�f�%�1�k�������`7Ow6�.�qoN[�4��9�](�z.�|�te��U�{�v^˔o�SI2י��dft�"("��7/v%gNҜ�<�d��P����niG�޾�S�wc�-�t�]ҍ]�U�ҧ�E�N�vزD��<���(�R���ͫ+X���}c]ˍw�y��eX���km_#*lT|_`�x+��+)K'�������T���I����R�����5F߫�7�ʄs1yz��
t�N�֪�Xd�o�K8,9��9T��u����쨉1,�FC�ڰJi�ė�j�Я�|-󭜻���P�5�GK\��6qb���JJ����)Ց����;��]	Y/Y�ۥ�@U&�oj�f3��K�d��7
�l�W"wGm�<���Q;��-i0��W,�Z6ؕ�V�#�����	��L�E=��ݥ:w�����lh����Nk��o�+�A����Z���M�
G�������.�ֆ�,��:�����rF�gNWeN�|�צ�gg�U����;$Ƿ�w%Ԟ8l<,�tL_e,�W-�ai�[g�'-d&�d��WI�c�E�{H��˹��B��9�D˕�g���3��OwH�D�u]��F����F�e#�F��*ҥټ��+�R��"���h���LK*�bO�ݵ�ۋ�t����g�ަ�ʼ���RkG5`-���O�d�Nu>�ˬ��P8�]�'lNBt����(���b��Q� ��cE˥P�v�k��s�(R':O�u%��A�ܛ�N��՜��ۙS,�0��Q��5`�/s���Β�	ۅS�3Ȍ�yΠlY��Kx��j�v��1�hKp<�#���FTޑv�Έ����X6[p�8�L6]���o:���%Uњ���n�oWo#��*�y
!�vk��;Z^[��Tnh�ps�Φ�}�;_>��5Y5����5�qU�,���p�6fj{/%+��ui��s%3L��$�"4حx�n�D�7���(����n���bb�rJ�vCV�q�ø��P�Y�k�����K����V]��	�\�������`�٬����kNJե�D1q3��Ci��F�&��<���ʽ4����W,u�-U�~I����"��K��a�D���W����)s +<XJ3@]��͸�K��W�f��y�3u�/jh�8^���%�)+Ү�8�6�i�2)g<�v�e��8��/	��Qqѧz�D�pG���VR	D]5�}��:꙽Q>*R�
�odK�(	8���k�]�#�^۟s�êr�bg�n��Ca�ۓ��*��R<l�+o`����	kʕ�S^�"rUw`����g3E[;�u-$\R^u�M�ȹ
5G:�&�:f�*��9�1V_$�k�m�n��X�oSy�2ͷ�k�]R��6[l.	��(	:�6X+(wR&���-]�B<N�S�nZ�w��o��y�>���3�XS��+F���wEQi���Ղnl@�R��pv��rc����k�f�٩Z��;.��i�w��uu�����n�bԝ2bu�	�|�W���F�[��V�ǎ4#��M���r�ѽ�r!�
,=ՠI�c����`��6_/R�I��NW��W�l��U6^g�掦m�n�w`�`�͏;8��J+nS��c���5��{�#Z�^T�.F�W	Ү��F�B�Ic��K�2(��X�a-|3l
�wl�R���J�ׂu��i�9��W��T� �]��"V�����|��@�ٴ��NTv�C4E�p���k�Q]6��A1S�}�1շ��Y�mܛ[����̹Zc��C�k���ma��D��u.vws��&�a!sl=�s-�E�S����+,S)��4U��aS����;wR�4
�}A,�i3�@�	ǰ�l_��dr�x��W�(<Z|:��E��:%���UM0vṙtíL�vo#g<�f.�W-��-lΕ�=�h�.F܄^lZ�79���ʬ.r�p�g%���X��ևa����tu�k����n��pj��Տd�Z�גD*ff��.�����T���P7xB'�я�k�J���6�������B늏��;]J�Z��Y�V�z<�^�X_Ύ�ǝ�y����Y��K{�\��`X��/���;S��Wuoy��6:z*���6�����T�U��Yy�l�`��'Ǥ�őY��s}T��m�7�1����u����o�<u�wP� �
z�T�n�}��Z�����Gi�w��̈́�kSw��Xٖ�y�aZ0�%���I���u���l��薵����IP����P��Fh"Q�TI$o�yEȏ�0ճ��ŋ՚5u:���v��-��`�~^�J>�L��u%���Z@X�X�r���!9�Rmu�wCD��{;hE� H�4"u{s&�:[�Y��'3M��naogm�Tt@G�_b��^��mh�S ��mPW�����T,Y�WG#]��� ;��T�a��J�(U�r���F�V)���G�r��u�F�wF���kE{��W��^��aCXE.�s��Hf���8b>�� ��5�B����a�6&��I��*����8����a����X�ҬX�A�D��E�����T�U�D
 \݌�i��5��A�0����s��F �R�}����c��eD ƛ����0O�#AQ��_�3������g�����Q�DQm�Jz �+owq9�EnL/��.�-�*�e�毫��ޫuۨ�����J���.����r[���x���Y�A8�Xn[��\X�sor��MTY��Pڸ�l.=|��X�{�\�k��fbW(,sv���u���X}le�,l1S2ـ��f.�N�m]��9v��v�C����}��\wcYHڢ�@�B�����c}�{a��|�`�u� m��m�'��PKddcv;�v�1ɨ��Е{��N�����r�k��]��fr|���; Òl37.�1�t�honp���,�4z@֐ˣX�,���������I+���]rG.ub1��#��e��n��"��yqR��/�pP;��)V>3%���IԪ߳6��m�Wtޢk(�2����
G+���ۄ�$���PL`T�8eܜ�«����0�%�o"m�Kͥ3PNaIl9��7kK�P�W*Y�X�����
�C��s2�2���P�s�U6]����&(
ua�r�S���:�'�6:z{n]wm��h C��hʖ�-�̱�;(�.�O	O��,XgR)��[YM-*�F�mB��:'�b�+���:ejs��ό�UWw�8�V�0%K��3`V���ņ�(�ֵ�}�Z��Z�V���kWW�l����s$J>��ݜ*�PK�9*�k=f�@�&�L��8�[X*�8��K#�o�����87���� Mbr��b�J:ˣ�m�Y}��SG9B��
������M�1#S�譡�w�\��*OM��u�j��z�p5\8� "97�YS1���f\ݙ�å]�R.�]m�w/�\͹�z���H�s`_<�/r+,I��<�cI��\;�|�2��8�B�v�(چ��ݏ����M57ol_�A#�Ikל�՗�D���0��G��q�&�mA#E�v;r�+@�W�x̱U�Ve+�{l̽ P���8L1z�/b��(<1i�"�{e���L���20+f�)v��q.�*�Bh�IA[�s� ��46�u���w�Xj�i��v��/=�70q�CX7�Wᖲ�'�!�LGzA.V�d+B��B�}�
�5b���	��<�NTd�١<��3�L�EY�#a�#5��s,P�@k�<����9Wѻb���zM���ē�ndopO���"�r|�u�U��ST�h��y�k`�쨓,â�KT�VGy���i�]c�����1����^d$�vyu
�9jI�)�n��P��A��T���%�>e�K�nd��Ì��Lh�aEqv^��R`�]�l��ɔ(����J��A���܁� R+�j=�ib��y���=����=z��f��5� {��lj�������ك!���4��;T${c�	��0�2���.k�f�c��;,�X�cV:9���f{B�)��] ���^�3GL�v�G@e�XS�r�]s��-t�⣤�2�v,Ö6�D�]3.t���)���S��v[�u`�;Lj�9��d����mb���h�%���<�Gw)w^�`rI!�}�1�-�Z�Xn�1B��1Λ�&�
醎����Vs��MŒ˼�n����'�}.�jH�n��&��6^1iiԪ��t ���V;�YAM0��\�0�f��7l���f���%����k4�	y�	��b��j6�C���x�m��T�r��C���� ]�lmbp
�!~�9�l�iE`M�9�э�-3��wĬ�XW��ɹ����U͛�:2�%]���X�2T�V6�V�n��d��)�gVa�j����%�Ve(�ћ�=�Ն����ˡ5��EB�XXRb'�����S�;�1gr�Q�*�r�.f��4/���r�s�7�8���)���BNqtb7�lU�� {��Yt��[���Vu�ڙ=���o��w�@L�l�s���3[��{Qu�g\=`�⫻�K.ou�#���	���J����TX��-��C��܁Xz��}��q.���Tm� �iuvf�N��/+;p���
]�xQ
�+�n�4W�Ak�;��� �+���E�s�j�f�z�����T�;��م��T��ۉS��W\$ڒ�ŀ�1�l�xԊ�w�`�w|�)n��k̮�: �Z霅Fn�ʙ�T2\ͮWWgc	w	�8�F)��A̤�P\)�ǐ�;[i`��v�4u�ٸ�D�Ǘ]�b�Z����o�Xu�o��L�N�J�(�ɘsT�V>�=�+�q����|�6�k����F>N��o{r9`T�u�4m�l������8¨�i�7�;Ws2`�3X��V7),�XZ���Ts�W]�
��%�� ���O�P;�N1+N�z�v������rC�L������3���s��f���E���JB�#zޙ�-�����������M��q��c���M����5�1�>\��e����K
kb(�8�Uq�ݍwiMVm��Rh��+�����i�*q[}����;y���V�X�J'[��>̱�ڳ.J�0�LRT�5�Y�Ӕ��զ�͜ &����wdR�ڃ�C�f@`.�ӔC�Y]s4���bJ��T5�����)7u֌O�4�Nȅ��;#����g+�� ��k8�su���J���"K�m[X��v��f��Y((�mE�+%��:<��K6�^�`J��,8����P�ǽ��4��B��E֣:Л�Y[$�La�)/�P�|u��K�wSw.�J�Yh�<���<�p���3c�ړBg��Z:${��VP�&�Ժg	��^�"���g�@7a���ů���;��!ʡ�*�u���[�es�I�A<n�՞M�Ԡ���1�0f���r\�.:Ñ��9�[�V��a�Ӡ<�3K��,Q��z�M�wD���D�I�����AR8f�h�Fը6�]Η�;�rST�s��X��'�8!��1%u��-^:n%f��+eC�qý�V�w%!g՜n�W#p��f�����ou��FTK+��#v���zRڈ�m��(].u��E]uR���iM�u��q��w\��:t�X˻\f<�,��{������:�4Y�r����)�A�)m��h��>���ܘ*�;��	��;7fH!��C78`����Z:�"(�����|��C��v��6��]�5}n���6t��A�}��
X�'���e!tk�VPyס%t�2u]_K�k ��N�,2��k�6w�;Z�kV��u��ސ$z�<ʼw���Ѿz;P� <�)+��GW+ 2b�uۢ��I>U��/r��Y�ѢX9
���r��j?Y��+�wV�żŗ)��*ב]�r1�5PE$u�P�H%�Q�v���Vŧ �o��t�޶�夽�����X�y땲j\�{������s��\v��t+`sJ
秸�-MfZݽ�X�鐞me��F��X3F�.��<:I]��׌`��B�»8�p���ϫNu��*wh�H8��X���ڻ�C��u��X^��(Y�$�����m%H�[����L�}������V�J��+���z��9��y��"�`�v�e�E�Ԯ�ٜ�mA��X������Kv�K�P�Pmt����=���T�G�p��T��D:jX3yS-)�\�
}А��v\�/.��ʾ�^TwB��Ҷ����Z4�����E[��S7�WGe���H�B��\����v����l�/�q÷|�7Cf��t����xev��-C�˔8�==[�v�]�7�X]�zȝM8�v�e�OMm�P�p�F�v�ɔ�\��4�Ou�B�83)���e������&�"-��0K��"� [��޻ǌe�*�+BK=��7-JX��F�v�{�}��T5k#��hK�Ӿ�>1G.�ҭ0!�p̙�h���N���TE�K1N'�G~vj�
�0e���&�\����B���P͞��_G�B�c��3�`sç(��z����q��o�U��ݥd�=$���,�����y�Z�.W=ʊK�P��epf��V�E�D�����]�7rM���Kwc$Ƶ�	�1���!��'�U��f$��)�I�4�)!�ъ���0�ȪɌ�	�C���F�uu������c�a��:r
Q�:��$�)݈bU�6����{*�R�2�8Õlue�Xfr|�Vkzq�{��Kv�	w]F� 4�4.e�.�ܴ��ڂ}ƴ�s�آ̭v�׶�p�N�&�L��Szt/��S��Y��;0ǵ��1���j�j��}ۘ��
��� 2GL�e�=}���N�����Y�g9/��̀'IQ��[����9N�˕������k[���n!B�Fe�ռ�?>��o���n�޶�	���$cw���
d���^&�l~�l�؃B��`��;Y77w^T.J���$Tm1]arI��۵:�!����+�n�gW]����󏒩��)�˾��1��[ߠ��4���a�L�+�Q���H��t'U��e
/{�U��\�rs�m�N�
�L[��.��E�v1]��F�>�(�6�s�`s-��=��h����;���z7S��\�w-=/C9���r˕gjZ(���Z�}`�i_ge�=��'H{�qj�1�l��Q�[MF�C�����]���<iR<r�����h�Z�t.q{+�F���Qe� I�q����ٖ�b��0����*�(u�x(��$�im����/��q�ޕ�(�e�a����f�%�Gj;�Br��EM���b��a�[�2�]ڔ�X�Ro+$Mf���7T��Y��DC�̚ufE��[DF�%��0��[��}M5�P5	��j�|��m2��\ �x%�o43�����Μ�X��xQ���hBo.>
��4l�a�$��3M�נӼMT	�)���Sj�5{r�;IH���	��B�YW��\l��僙��F��elz��7���3��o%ʾ��N������m�[��LL-֧�Ɯ�+��NJ���d��a��-�e��.a�[��%-�s:ƅ��qMRټΗd����tmҗ��Z�����:�X�r��F��:�I#q�,@4@�%��La>fݥ�ׄ+�HEx�I�ݚ�q(�z���:�w�d�����	��'^F�"̚� /��̓%n����M�}U���."g&	��Q+�v�NQb�1)�N��>�p����Rbվ�$�y���2�Z�b���AK�t"<��æ�^�O��49��j�C@����]:��q��7G,�cM��TP�[�yd"9�S�aq*��ڝ)��rl���O�;;��5��:�ۨO*�'o<DP�wL�c�ͭN�=),ε��u�:�Y�AO�2���n�b�dm`�A���7ŇI]�.[Q���!$��;��/^d,훤(�1��yW��(E�x��1��)>�!��S;(н�鸴��Gw+{,kQ1þ�F���@��wG�:+�<�6ز��]z2)��V��.���ov�L�����V������f���84o��ͥ��gPmU,��7�-�V��fO��xl+���M��R�KIbJ��ܾ̠J�:���م�fYN�ӓ���@�ht�Њ=���FX3����Ui����om��}�J��	��5[B��C��s˧RڷS5�[��w��j�����x+���:G��k��TB�iM�\�������N�sk��YU7C�'�jW��FE��pR�V�e;8+'A�|~F ��*8��Luc��J�i�)iҠ�s����n�o���bb��4i�ɶɌ����Z#+w�-.�]���Z�d�P�u���N==�n�A��(�d;�w���{�2�m��)>�P�%�}O�wS�\�A��ّ���!��pe�wM̒�e��FZ��	������da1����{6�-d�\����I
o���/r`ViJ宩����	m� {�b�ݥ��A]@��L�Y�����bh�n�ڛoPg>�u���w+�'�-�X�
���7t��6�6���Ix-��0[�&�sx;�k1���Ly8����N86����9I�<v��T�����E�z�.��ʔ�4��06�܀ڏ�#����7NA��A�G�Ԩ4�4��O;���|�����mH�A��O���4�)Ks�n�`Tr�SB��˃otA��uu�De[+�<	Z�s";3M�Wu�<��m���̈[ģ�:�Ъ��[d�WiT2Z�y�k�F�F�	\l9i�q-B�9lN�-g�Lm��-�B��K��y0�:k���N��]��4&_u(kM�}�e�h:ǖ�G�YN��:��'H����{a48L�ui����,�WN�e��:%G�BS}o05�E]r�$rv�:�hG��V�׸����	9wo���X����To��m�}�w�N�1��F�p bF��f�Gs=�T���& �v�s�p�(vy���I���f��y�Q�zl�^�����رs0L�4@�v�=1��wW. ��a�s�_P^��\Og���[��W�19�M�@�����W�p9LIY)�b�Ӡ�oV�B�Mco�Vlz��]�V:�b]+pn�d3�usM{w�ie`��[Ι�zr�b� {�@S�6�T}�Sw���\�D+����6���d�С��k{I@���Y@���di��
����]����U�`x�#�bw"ΒL�;Q���uwl��,Y�gwfP�a$��f�2H�C���R6Yͺܧ&�rvfG�@�%�U0_3���Ss���Ѕq���[��p4[��\GE�i�M<���e�!j�.na����]ٲ�@�:$��Pٕ؈�wuҖ�YkM�i���2�٧+��P��c�����֮�����_�q�UU�b��_��zӋ���y<�/&�۷nݻw���N#$�K�1X�Q�Z!q�B��jB�O-]�����a�?��Tk�0ZiJ1ƣ����h>F\��N��ţ׹ׇ��i����7��s�=�0�W���n8-��2(�eEx0���7�Uײ�H�do��7�R�;�Ƕ�'`�6vED@�$4�k���B+AhtM��;�޹4�J��5@�B(�<�����}vu��d�k-n's�\���el�X���GX��ѕtY ��H2r8��X׹��i:C��@�ٔ�ɗWr�˃oi�I:Z��f l��ל$c�4��Ub�l�m��e�#h,.Wu��oN1�V�/���\�/5�co9w�z�ܗm�w��N��@v0dP���m
]vm	�C�֋Nu&�/v�r��R���gE�z��x�‸�;	Rܥ�Ѳ%���؀w�Y���|���"':(�c���QU�k%=GO]AwU؁��HVb��X���t���.|f�~��S����#��G�*�`9�ʷ�S�Kc.�t�l���?(��ׁbK+�x�; �{-�V�
hvn=��=���RتI���*�q�ĺ��n��fR5�����SE�U��᡻��ñ=
yO"�Q�qf��[X8X�:fu��*<Ҽg
2�΄���lKowa�'������0�)��\�z���^��BF�%�^L�=W���me�o�f��7��K�;xd��Ь�c�`�t8gu���񕮆'gJ�(ku}�GKk�@��ٵY����C�dO�D� A��14"P��.Pi��D6Y�\L��P�2���Ha*8	,"�0���-�#��c@��D�'t�1�`�VR�V�J��E�����UP��ۻ�W?�Ow܂;��m��:�˔�Ύ�tWw`������Ȯ����i���钅{��B^�ۻ�������%����;&�A�v���8�;��4�7ĺ4����$r��ܹ%�ۗ!4��9�K�.�r�v�W;�r:k����Ⱥ�����$�7uq�n�D:RRd��].2���N�s����A]ݻ�ܯ7������`��=�x]��;�%	snwus�)���w:1p�������:Jsv���"��K��d���'9&
n�7��]ݓ�Lf���ӹ��!�׺���%»gv.�'q�v���YJH.�\���%��!BR�s�C%'pwwwD˝#��&)�wvM�Ӝv�$�p�]���������y����_�������;f��jIj����hK��5f�ҙ�wr]��S���{m�����]CY)u)�zu����W,�oV	ag�
�@�R��LE	����K7�C}�b7S�j�����}*�\^ӑ��=т,��]��ˢ,���I�@����5�;���3���I2�&6粯ni�b\�`{q����mS����>� ��#�[��^�1xwi]��{�y��Tg6�b�lp��o���~=��{;O�U���~"����VԭqA�OT���â^Y�����o�H(ޥ+�z�G�%�+�{��t��,sX屽ݙn*���^�vi�WqPNٌ�WK���s�`�0�/rV-��k�.�Fw�r��^ߣ==S���y���8��<�^�]
j�xTʺŰ�a��)�Ǒ^W]����0��H��j���D�7[#���
v��M�iӻ83�8-Ϙ[�����έ��NNHӧ(qI�5#26�;���W�w[C�"|�3���1���B�*�lGt�f=�N���A�w\�Í|Z��e�r���g_�M�o!OYΪW�M���Q�2y:mJ�hu�z�ك;�p�25���f��ø��T�p��B)�\S&wl[˯w"�>[#ޜMi��:��l��N��Y� onںQfn���!N��d������/mO�)S����}���Z/��p�kC��E�qW����ל���ʊ������9�?WS��zo�=~�쪂bE��ݕ'9��^D�$O#N���x�v!�W�zT����~��?��<�v4��k�gl^Y>��l�x�W^������y�.�7\�x��6C��w�`ཋ�f�6�2n�A=��|�tl笩��G�S�{�='h��a�P���,t�5���o<4�f����X�	���=�+��zp��[�z�膷��7���H���1�8z�Ы��꣜����n�c��3۴�7�7�S��������� .��B�ᝲ��b.w1���x��L���M�����8�P'޺M�֮@�X����m��{Sվ���׊{���0a�l�������?Zko���n���w}�Ğx�ʺ����0.Đj%A������\��[-}p���絿Wc��m�@�U ����٧�h�Kp�*���ǋ��u�;���`�#��q=�t�~��G��o��>�0Uˢ�I�ͻ���6�ֈ��+�oDuu���ÕE\��jz�R�@g����!�8���1����<����c�M}�%<���Y���]=�(=��6�]u���=����x�E�{�C�JǩL�o>5��nC�Mݥ=���U��5y������O������+n�R��S�<hS�k�k��q5�Q3Ͷ��d)�Qv�y���k����?�K��k�)��W|OqI��+�}�zW�O}=}��Lt�g�A���k��cE��fS�kJ^��:��~{�Omw��4�����N\Ϥb*2�� �w����`=��A���(uzh���&7�V;D�����I�c}�$n'���p���{8����5��W��a���#^^��ީ�{����*������F��ݍ>��"��H���L=ܚ��j2/꿽��)ܯ)�����X�:)��*����[ܲ:��,�l�g �O&���������_;��ݾ#���p۔VYf�r9��]֌���c�D䬒�X-U�a��ﹰ�Ǖ�]��Q^2WL�w4	�n�>�0^%�sz4Tӳ��U�*j7���\ll[����u=�)�ǽTz��P��J��Y�+�Cpc6���ѹG�}�GFQn�i�hY2Ltaڹ4�*�c���W_�u��eM�83��X���V�Hm$ǹ����4g�S�@ۧ3qVQQO�F췿 q�K�g�=�O�<�y���+y�:I69�A�zx�vY�bX[э�n �k�\�x�du��u��e��`��b���<q���ضD=~@f�^aL��u�r��}Ig�Sg�ܚf���5��~�s4�g#���ݎl��Q=�{v�mp���;V2�}�T.n\C����^��5MS�9ܢOuފ��1#6XW�y�f�3^<�q^j{�`"T��y��������_���W������W2|��8,̨�M\���/�����+�<�==�_����ho=��k����H�jǩ����b�H�4�dm!ק��X��t�ӷ�N��<ˁՈ�V7�(dNcO���C��Z��::�d�c�|��8�罎;�*o%L����`j�S|i����V�3���f�ծ�,��۽t S�Jz�V�]��.�G� �m�wۃ�+���[��:��ʱ��h����v�N�>p��-sn�����uHgH�w�(�Q߫�[�^h�`5㮝��ʊ�_��t����Bsgg�9�����z0k�⬧��uo���ac�zdr�d�MNomb�L�����7�D#���:x@���.oeݬs��{����VC^i���:m�t�^�7���E��w���Or���N
�u��F��E�pUxPvN	�����^�~�������G�(�����KY���=r�N��ڀc�Ȋ�"E���j���K��D��g�n��SN����ͺ.j�ò�յ�7rEȇ�kD��(=�>��c՞�s�j(��Sb��%�����}uc1����ٍ���<��,���8�\y��$�T�j���= Y���힐��� �mc�UO��U�1���V�u�-��j�^x'B�0hȨ��z`�ޭ�'`�܆�Y���s��ЁTj�n��(���`(Զlix���_X�Wϖ>���1�Ƕ�nH�s����N-r�i��y)-糗,"�^�d���{�ܭۏ���9-S(s��"��'-B�����������|���<�o�t��]�E���^Nїu�q1���W�
��c`U�]"ݧ=�������jQp��h\9����r��b#�v�G�#sdFN=F���:r��TW��j��Ox��T֡�NJt|�������9�0��eϫ6�?��f�)�����gh�B�q��W2�]X�u,}N���Պ�?r�%}����o	����O_�Q��} ꨫa����,�����{^(Ŏ�A���Gʷ%$�X���H���h��싆#��o�7�E��5��V=A��m�/�7���D��Ϙ�E{O3Ee�庺-���I{)B7ϯՔ�>U僸�`e�����A�w�	��y�=m���v���Ok�_SNL5z�=0�'�l�0��s��_��	�qk�7��1U��יf����'�� �V�w�,�ֆB�Re^�z)�����t*P8P�Zu�k�w@�.+m�Y:$I��Ўȗ�BU��Շc���d���V{6�Υ�Ts�s�/vK+�Ba��l��wDCZ�%\�Pm���\�u!���r�N܎ڹ�M?O�؃ubȂa�V���؊ dU�s�����O��Y�����ު*���Sl>���k,fG5��y����s9�p�G��K�ls���'���[-t�Fߠp������n|��o��i�a6Dt����s�}��'�)Q�5}k$>�짙�X^�zo�������_��X�3�L���}=����>�Ro����5q��Wsc�����gZ��.�x�_���7��ݯ�?M�~�|�㴞\��'fo{@��7��׾]~��mP�8?	>7>n�U�7M�w����񇽪8�H�x�x�q[t�})�Js(R�8�2��7��s�gn93*�ˎz��k�+a��ʶ��j��^���~0�ήGϼ����H�c��|_f����m�Lt�g�0b���[�a>vs.��
͍������ƈiu�N�137W)�2��/.f�W-ո�>y�a����G8����N��zaBZu�F��$9X���1�eˬ�U�FR��#�P�:��P2�?�q[VE�a��^�Ut;�+o:[yG�C=��K�ڤ���c�;m�*���̪��q<�k�{���#���@"� �ľ�Oh�qW��ґѯ{���&k��Z�8͝^~��5xg�g:]B�sc��W�ܩ�/$@1�^��l��y��v16{\I�u��ov4�Y�t��h�`�ti��rhDޝr��)V��_s�:p�r�NQl��=+r�d���q�f�=�?U�P~�f���C�����oW����5W�5���I�&Mx�v�@٧2@�Ʋ���3����;)��~�~Fu[��i�m$�<�=D���QoVw0�C3�Q�۩:��n���q �bEy�ڕ��^(}�T���٘�c��L��.	�6y�v4������`�] ��p���U�׳=�`v������+L�ޏ���L����v����W��=9�T��H�����C�Z�0��z�R_H(кN��)����<�xP0����`�[�
Jh�+D�
�o��b2.$n���:�j��
�#OofT��R[�.��gv���H۵��R���1�v U��r��[�(Nw!t{��Na[�9S��K��%��خx�1���;�
4z	�;nAv춿^S�����1��>{��hQ�ɞgu_��S��|��>Y^ӕh=���I�f�w�1��V2�SA�luj�I��>�;'��&���NW��Uzt�����ϝ�H0k�L��u{��M�X���8�Ozm_����?9��=���K>�1s�Nfv�E�zP9����"����{՚u�Ӥ�X��w���+���Y�{�y��V�6�1��r�/�~�U���i@�W~Î73��>-9:���{ޥ���}�,��}��~��d�ɢnd��������$�^���a�ꆪ{� �p���]/k4,v���z�S���g1��P0���Vvqo�[Qz��܊�������"c�+�{���gХNgd��:N��w��d�dl��7�� ٓFw(��=���y�H����N#���zͬ������*��v`7�0s7X̮�n;�s��'�w��kS
% ^�o����ʚ��ǜgd�:�I]��|�d�n\�8�&g^�<�t;-۸��CD���Iq)�5>�ݬɘ�Gk���H�&s+�{�:0튔��Wz��Z���zX���K�\��V�c:����������x������=��W�k�Y�l�q�y�S7��\��!���1�u0a��?Z,������+���0�@7P��v���4�2��Ҟ��y���k���0gy�q�j�
� �-�é��l��3�Y����P�",����=d����o���H|�g��+)�p��q*��fn�O}������y;�P�5�-�s��s6��>�r{'�W����^�������=��i�q��E�`|c���ܭ�����{Nߤ�TN��bAw{2��X�ޗx�8{����۾Ѧ��y�g.Y��]�p��}-G3�܌�ܣ��{;�T[P�6�eJu/{����cx���p���m"�e�%�m�~��J.[�&dU����e<���]�V�e���ã�,��v�ۺ���:�	y�K�3.�1ص�����þZ�Mr���^�a����LϐO厰�,�ml̕�zc�.���%� �L��Q��E� i�{��X��tՏ���F�]�����AKe�[�Ց���{��V�6ƕ��"4
�vc�X�"5j�ѧ�v��+�W��u�o�m�ҵ2;$ˣt<S�����{:����,݄v��Ǭ�j���)�	�V|\��-�_�s�6_]]�K3��WWj�*����}5��}|�5q)�h���avWt��UwLξ���u��y�v�t���L4u��C�a�Xs*�.�N0�0��NĨ�Ѱ[��h3$+�5�RP��^Yt��>�Zp���*ND��_0-��'_GZ�4��I�;�B�vX����P�+N�RI�P���LMt�y���}$�%X�,��j�E#��z��^r'WhV�.N�E�gt�؉�Ԛ.��*`��Y鶐dam�ڽ���D6���<�]��A}�7���zr7�R��yeun�3V5n���3Ody�J�v��*�3�w\q��(K<HM�yy6]�o�s/�L�&��eiw���Tz�:����c��/���#��"�9�CVJ R�򯞘r��#64�lz닮��Rkwn%����p}X�����f��C�y��/�U1>�&�{Dދ&��g���Ԩ����s�u�l)�,62����ǝ�Y`�o��v�5��z��	\�����k;2���@T�#x�$���GŮ9�n2��$>ch�bw3�>�m�v��*�W;fS�ܽ�B����_���>y�3��]N��/\�3�PSaÂ���7�k�*�K|���'����G"���ܹ/(�jzNr�¬�::c��8\�@�Uȅy3��6�qO���Rg�x���z�}d�cGM�G�]]�x�#B�ɺ�R����g1�]{:j���c;:=�2��ۮ
e�Z7K��v�K�}�G܄1Ղ�pŚ�)��0%�u�Kw[�;�ש`
Y�伷��mϭIƸb�C+�5_�{��i��d�pV`��R�Bk��}x�R^=kvV.��GP����������8W^U˲�
t^$b�����/� ����B΃\��J럹c�Zz;��Q��[��+h;�d�j�˝8k�{�K^�NJ��ζ:�wwoe�h�������}�S��L4�'����4%G��aW{5�a1ݐpvt����Rb��K�-7Yɓ8�[�x;��t�pܶ#W�M.g'��V�ͨy���|!K6��bƲ�=�R�����p\����4Hd�;��L����x�\�vQ|L���H��Di��]c�Ӈ�..��,�r��7m��f� ѻ���(�Y�t��A�Ӯ��]��`��~�\��	�ڏ�Xl�Ľ;_lݘ�sff��0�၌Lf���m�X�����Q��Vu[F9M@��-����z����z�4W�����e2wk��9s(��;�]�]u�����!���\�wn�';�3��N�t�"SF.WC`��w��rR��4@���1)\�D�u�E��d�;��q�@;������AG.�D�K��9Ȅ����ۨA/.=ں���d�79�L_NWws��K�ܺ;���N��P���Ӳ�sz�/u��	y���y{�w\{�(��霝��/7����;��]�r.�Nr�oz����#a �a�`��6
�)#��yq���;���=//r�H�n���o{���z��ys���sy���޺f���{��<��v��v�{׹����]��w�p�ˎ3��7�v�8����'����no:s��΅�����ۜ��N��E2�eG�m��-�� CH/gu�sr�N]�=۳�{�o稽�\����H�{�"�t��u�v\�F�v��{�K����|���ϙV7D�6z�{�it����������i*�g!bY�Ĭ��21F��s�x��|$�:���<b��Z2,����������䁛X�K�(H=�=PŴS��"���%���Wn��M13�8���` �(c�V{ʧ;�~��C�7=D�셇RYA
�)9��2�Ӂ��k1�܂��(.W㷾�V��W��dL�)B����Ϗ��&=��ٜ`(.J��� Ȭ�`X�)g��bkUV�����H:�)���V�B�:E;�ojÒ��
g%�j+��Blo7,=Z�v6���x'to�U���z�x�����!������������b��>_l��2u�?E\L�οLNf�Krw�s �A⒉d^�SL�*4��Dm�754C!��= ��������kL�����o!��k�T�(Z4H�(�?D�I��"S��"�P(�`-�6皼��tVU�(6dҊɰN�ĭ�j���Y�N�&��������)�Oq�ZzO��Rr��Ek�s{.���Κ�7]�W�a�����G6קg���鶤�.��0���Z~X�A.@�v�[LK�����k���Д9M0�&C��&���9�cbYs߇U�7_��sYt^����eɂ[،�ʞ5PA<�_f�q+wkuޛsL��+SdQۦ�Ǒ;ϛ�'�598��oWY�I���q��NG����=�0u�\�v*���]]Qp�r�qA�*�;r��綨���m4�B�uvN��׼VV+x���旻�8���4wH��tzz/���5����Ѕܧ�˼�	�Z$Ȧ>�o<o>]6�dVjh�ֽ�M�����>����=��f�L2=���'����^ |6�"�o�w���]ڞ��о�R�u1���O�L�������m`�jeՏ�	b�~���]CY�ܳ|�QK�'ke�̋О���Ƅua����SG���QE�'᎚���DxMy��n"�𨘴l��4��C�;+
LLv9�'dk%~ޠ���:����2�[��5��K(�7���n��X]�6��.��Cm�3Ô�6-����竣L�C:x�7����m��M]�Ψ��ޏ"�F]���>�o���c�["�&�}]~͊���6�f���jJ�����Og#a� �sy����R3��3gV@�t��T�<�L�k1Q�l���o����謲�����m	ثd����vO^YX�ӌ�u�6K�9�p�p��m��[�W�B�)�_$����7��}�O0y���A����Rux�
W�TaMJ��F�\:oO�'��!�r�Jލ��z���־¬@j�W�����w���[�z^�ء�U�t�a��w�b�㚺�pb����v[8c�	C����l=w���Z:� ��$1��*8�`v��K�Wn�&([��@܄�XT[�<Լ��3���EJA4K����_�(ݱ5P�w7C8�s;珽�1�&^Y��/���f��_Ab�ΙF"S�(д�JqM�}���<�0q��K�<ǻcqc+���o`y�D9AĈ�!�_K1|a�4Ҥ�<�LS��[����=+*��l�el5Owo!�{��b���ZdO�1�~��>\��+���ʠ�n=���ث���;
�z��7Ώr�ߏ��3�0m{�r'��e��kȇ!�����N[�(0��=�FtV*�0�a+֥s�Z�E�RXǫ���O�H�x�"�Ǐ�H?���6Y�e�A�)��K����d끞l�*��Z��3~�Z�@Ot[��=�hl�mZ�T�1��,hA��s"�c@OH���"�R��Xeҵ�%�U�Iq~Uby���6g�L��ª�ٕ��w�H	�0BC�O�W�yy�Y�'ѝE�5)P6�=�X�9C���pF�e� w�����̹@����9����x��M���o�9.�:��v�9%y�$��vb#k��
�7UY�A����t�ý�UޑhT|`���?j�?�dh�/0�P���G}NwZ��&�ÑY�5�t.�����3�y��W,R����0�M*2�^�s�λ����{Sȫ�񮯯�S���٩��NY´�R�<��&��j�v33΄*��� p󮋣㛴��K��uG/Q��oT^sD��ݙ'8�����x�Pi��H8"�P�s�w�63�0&P�/��!礫��-�x��me��צ���X��������z�Y!F|�.2�5��u] S;{(x�vj�cϴס�6Y3
|�|"�h��F5+��lj���gaK.|$�~��GT�x^�6�as��¦Vq���u�����iƱ�a4È�c���N��~{�"Sn(	���B���c��ӱlT�ۚ�8���ʹ-r��ƚxk�=��-�'C�	���}^!��so��ɽ*�\�)�P�'&���f�4���y�j
J��ټT5n'�-b@1b���*&<>U| ވ��[�O-����[�Q����
��~L�Ⱥ^�c@i0���)�����h�a�����m	Q���Q{x2�w{��b��'|�׆���u��J.�s�1�����NY�6��a��J�U2k��qU����m9�ɛYF�6���:�F��wBʮ��j-?2N[�.�̘C���A����D����s�K]�?�z���&�~-�'f�ϕ��`Z��v��F�8��%�R������+��v��+���nV���t84,���8D\��a5������}ٖN�\R�Y��!�w.������R+tG�W+�|�eEw�l��[�Ki
��+�۱���nA��'rk�gpPk�幋1!ϒ%�Ww{z�cs;1��c0��yq%/	ft��#í,A>�c����s��	k�zv@���%���8�r�Z�[�6��	�h]iv�=-9٫e�]Q��:�Y�d/o�O���<�cC�(GW� ���ޛd����ו��=w4�j%�OVo)b��:�,�����Nܳ��d�%p���H�Y��f�հ�>��n�|=����0�vfԢ�lc�C���@��H:"�����;�t�ݧ_SLs���\�*���=8^��\��z�oH~9���r����Gf��n=����1�<�ծ]ղ�z�R΄�Ƈ��V{�Bs�W�ޡ�f稙C� Xu��9Iw�޺�6�@2b-�z�S߯������i��
vg��=>5 m9�MO��{��8�L�`�ɽ��o6'�&�lq���ܹ����/6��x\~UW�u�&P�O�R�
�%cj(zo���Q���I�so�ʁ��c1�� ��4�®�aG���[ռ�_z6B
Έ��&BA�j��j��Vkm�� ��t�&��=$'%D�/`�4�ģI������{gO>��xc��fFZ�&^ ��ϽT�ѧQM|2h*�-��:zqn��z���gGH�2��Ә�5s�]��8wd�Y떥�d�I�PL+qo(\���D��\cycR�y��o9b���𹓖,�m�]�!��bU�6RE�Q.��k{:�(U�U����{��:�zo���,|���X{�MIZ_]�~���+עA/��nxN���D�6�ȣ)��Fǭ���.7�i���L>�*2�Ũ׾��`ni�6���cXe�)e;�iRNw��k@�^[\Øå�ѡ�-�y�pF`'��6��0����-�?�9�kӳ���t�E����~��>W���q���o��OT�"�wwr���it����>aG�>1�B=p����G�;��g���9�c
ʝ��ٞ�=�Y�����c��|�!�M#Z����jd.�?4~]��:�s��z���56lr��6;P�(��kFy6���y�)O�ʦY�����ٶ�3��G�~oj�0���,RS�2����n�a��"�:�è1��X�~��S� x��Ph�"G^f�⹹u�U���)�GO�|s�_���k�ʄu4���`�h�9SE��>|-|@>���E��<
PU+�xw'�|;<�7�����}gd��i���o�vF�W�A��uxMq�.��2�X	v�p����ćg��9˝����^O�v;�A�6�~`/�0����m�9�>�yf���~�8�ȍ�����V��.�^u/2B������d��]b��.�+���)�J� �g���^��n����!+2,�(پ��1��E�Xf��!�ܵ��� ��֫��є$��6�+�X�{f�'�iV���sg_`j�޸¦;Z���ɛ݁+�K�M�nߍ���'�W�2�6�cZz��Z~��RLb|jݟ��U���������A�9՝��� �(,��W6�gY�f�2��-�<�Ӽ<3��d��ŕжou���b�y`P��؝���r�t��%�x��g�o�C*.и�%8��C�Z&:��"�Ӽn�H\��qjbu�WN��2=tB��r�N�bT)Z�,)�u�*��;�zCu�<��ܭu�SY��)�����t"|��O}>>:��R{
"S���H���gU� ؜6�����M�8�а�oD�#�����5��1o��H�J�&�h��ӲhF�o^L�fi�ɺEs�$ׁ�A��ZdA���^.�:*,���h]F��E��wd
��y�f�Y��4�摴�p+��g�`�ԃ��"��p)R�׍|в�+R�~����zz�WX�I�*��熫W(��W�,m�a)�ݛ��Ç���z�[,���ۣ:���;&����C��)�P5t,ۙ:���U-t� f��Z��GGh�/1]Pa�����U�8K;���:���������{��)����7�7�K-�}ww�Fθ�ӛΗ���B�eӋ0�{Ͼ����o7ƒ����2�0!)>u8nKI�l=�* �eD�^�5�3Z}X�n�q�CQ�#�m>���yp�g7}��H8leDD|�>��W�����H`�Hym���&� �1��ͻ��BՇR�{p]��^���#9�$c��B}���z=ڬ%�k/��Jᯗ�Y��	�v[C��XsW��@ߙt�8s�*�P��r�A�����z�*��.qE����0ҡ��-�
[K�dG��7�<��רm���qJ�sR֙��R�.��jJ]���l�:"���g/T��  `N����yO�පS����y�zv�Q��Lui�a�h<֙�I����O�g���Zgځ8<�?�������g��hhL��'�Ft�{j/�5οf�A�� ^��W#^i޶MC�.7��S�fkg.�UUpݗ���p�ZW�b9���D]�'�5ޮ�'*[�)^����2�Q��nN�3�^)3>4A�O[;�;M��0����G66���s���d�	ږ��D����ɽ:�wb~���ϩ�"e�$w�~�{�w�M��ᩭ��ҜI��!���}|��
~�GJaW����ﷂ����:�~JS�
�Z#f��k�<*���x,y�H>C8!<y���d_WWFKw��*�P��JMfV_b:�Κ����f8�^�������^ۂ>�^p=ٴ�ޛ]������F���8抰g�+&,|f��q�G-��W��M�*9M0s��n'�ms��HNx𓹵��ѳ���o�:������������9ŏ��#ω�<��9�s�1(�e�":,��>�F���D��loUk�X,b��Cc�v����g�C�o9�b$׬�w�_E'L/�J.�s�1�]N�@�S���\��=2�i�Tڳ[�=���P�Za����aqv,�I�U�=����XIzS+���~`*e�b����c^к�?}�~�v�ψ�d.:`|#[�ӳE՚�`Z���v8�0�-Gs�#�ٖr�sݵ�6���;��tT.ƐW�����s��_j��D��V%X����˲�zmVv��u���b�|`]Bv���@AC�0���(���4w	�op�'���`��&�ֱBW2	�^�G��z#[��������%�5���2"@�	8�j��R�~���v{�X�_m��:~��!�f�I~�Ǥ��-�����lZ�X�c��2����撖��{����[���Ĉ�6��;��4ϳk)z� �S@A��T6�n=q���ZRQ��>�#�L9�!�L���d&�!�z��ǳ�#[�p�4�Aa�\����E����lBߖ�Lي���luQ�5;R�<��3�Љ��;F[��n���y]w�����f��1��  ���x	���p		A@��J���k8�a��2=�"D�VrrJ�y�<L���)A��l��7�M���xx|���Z�HL��Ļ������Zf�������\^q�|�^�N2䥛��QQ�Y^bci.�ٛ�ߘ7��;ݐ/�f|�b�O���RL`B�,:.���V0I�o��Sv��|w-�]���;'��8n>&�cb	J��)��t��(�^=zޭ�]�2PP6tD�X��ՏN�������/�ev!:vG
&��܄��.tSL�J4��]�7Ǆ��p������V�?��km��O�)@TJvl�x�
����%�%:O��Js`j�Lhi5���� \��S��\�WQ�z��P��ǜ@P�m";��hN�U�Y��2�ā��$�E'*y�Z��Dr)K[�gv�q���av��d�D��t�bvx7Vt�Q|*�Y��8�*�Cs1��e����j�|�y	=��uyt�=��l�
9��q"6%�=�\�sz���~[g�)�������M�<�F7C�1���<�E��jd.��w����kk��OyvH���a�EK�;"�hBUmv4�O�x��y�S�T�6VŻ�n�"1	4e��v캷p�,��,��8G�;��.�)`0PP.}�ue���+�u��f�\���98XH{�����`/dN\7j�9+$��\gK Ja❇�@^�c��g-%C�/�j}�\�J��N�cV��i���	Э���0�p
kͽ����'t)֩4�����Lj�s�wr/��ç,
��Yh�;�)�JQ\�����&]��ށ+������SV�C�g=������p��/���4��ns�sk�Sj�Ė�3��Q�͛���[ܷVX���[5;;q��O�nQ�2ṣ�f����L<�(;DM��U��e�Wlc���)pp�mjT�v�:���	;gd�iȯ�����nϵ<z1Xׄ��tb%���Y���	\���`=�0���#2��9����`�o���vr��Wy��p;��L��$�Ů�+D9�N<e\j9r�>\�nn�<����N�ؾ������u֦Ѭ�ٽt:�fF�;|�pNʋ�.�6��.V	F�^���$8o�U���~���0���X�����m��Z���{�-듵��2�r`�k370��#�$��$��*���Pp��T����k6��6W*f��9�σ���Zfk�S���<�5�wf	F5x3�cX�����9��ک�3���EΔw!iu֥)vn&զN����%��3b,�۵҄B��`�R�ݮ��q�7�&p�@7n����+9�@���-���ô^��eT5�@����,���NoM�J�f���К���$�
�R���	5���9���+�ూ�$�9�ҳ�J���ӸD	^����R癒.�ٖʲ���H��/n��"����g�����c�[��:j[� ��u����һ�8�]+��Tb�ғ1��BU���wo�Ϊ
�"�]�噖6E�9���38]ܭ�ղ����)���6K�s#l�W�u>�[� 
ǀ�սv���X��Ԕ�~��tپf�2������5���r���:!�e`r����*受i��b��Y)��#y2���������
�#�絝&�7W�ENJ:�{e�Q�+C;vdo9qp`�"��7zK%�g4e
9��㵜Lt�%>���г|\��v*����8�G���z��W:�ҕ���L5�Y�51��F�G,��af��:�N��:3��@�S9���|�t`�$aK�vU�zU���K<��wAݸ���w�kQ݌f�E��$j�;:�ɒ�)bn�ɽ��9��93�]zt��_@��MS��\^�#۳�he���|f��)\�5�b�2'��Mٖ*od2�3�ۮ��<��3�X��E��E`�bu�h΁��+g;4�*v��H��ӥ�jΩ��|2��/� Վ����r��t��w�T�)��PHi�B^���o5gR��92!�չFp�{�1��<b5W/9�x���U���;U �u]ҝ޲Ej������̰���l��)Q]C#��π�vI��^y{�;�����������R3wN���x��w]�9�������ɑ�p�y����1��)ι�Ng\A�!#��s;�Ns�#w\Jy�w'3=�M�i��}w��_N}w������9�Myqw\s��rv�w{��WuȖf�!��%��:nyyE!zs������ݹ�[��{�7����
$�;�1��P�����v�F�)������DdI
Nr��$�tA����w�p&�2A��We1���f	@�PH�]�A��9�r���䥆"ʍI��4`�(�ܘ��dȋóDIyq/��F $���5ڐ2{��4"ےb��l�JI!MΐJc#�$���{�x��� H��~]��i�c�2�%2wvQ�n�ۮ]$�$~$	������!p7⟯ѐ�O�1�������J�dY�Y5"=Q�YT��S��*��g3�d�ִo%��VF�-�j�bkT����޾�N>��]�:���������ګo�ڴ�JX�Q:��U��;k��;_s��L�0��5�=������5�E��z�G�#β�-}�z5&;����� �aHX�ɧ���^5�>��4#��N	df�+)����D4{R�/˷�onv�����XH092�������Ï�^�63����Ѐ�)�v���\����&�N՟�[������G���2��J��@sͼa��!-�?�__����oO���?e���q�N�9L�Z�E����~v|w4~��W)i��
K��o6=Ų/����|�|�m��N<�V>����/8��W�BZ��!�#:�C6q�{"<�О�=;��`b�����j�$tĩ:�v�yahMe7;�^ބ�_������ ��g/���T\9�����R���b����CN8�]��Ӭ��d.~wA���N�j�Jª,)�سfSPN��3�u���D��\��Qpꀸ�x��
�\3�헲��}})�S�&I˼':��7/�5Ls�������
յ\\]�ٶ�M��m�DcH�H8}rWC1��˵x{�[�G���IL\��T{�4������|�uɏ�H?b��1/�}\�i�n]��t�.��ٙm,T�o��HB�B�Ky�meb��+L�EgV�5d3����u���o�b��vZ�+�۰z~������n�;T���}��J퉲���ޜ��}�P�����������{�zt�LeU�W-n��b�7H��Q4��.͔��qcF@��gb�	��f���B�iܥβs��b���mT��~�6Ⱥ�7\�6��z�3�Ϝ=� �k�u�o���)w����
�o:��NlN�
7��
���B�c��;P�Sû4nC���|f\�������I�������>1�"m/^���W�WB�8��U��c6*�	�C�0��0	�cd��-}%�6�p�K��C�R?2i�a1��ͻ�hZ�R��_���V��������ة�۶��7vY�r�y������j�<������`�#�Ά�4��9�N˲��u�0�@�wT*��vN��E^ws��?v�IT�5�,�x��r`C�ǴBa��s�쓭��8�����+�=�ء�h���K�v�}�3.��g�9�+�Q'�����q�C��-�ɋ��R����s��� ^E��Zd���HG�|pE�����466Ou�x/-QL�vpb�\�9T#9Ĉ̞/sQx�כ��a ��r/@�����Y��^>�@#�埑�T�Y�r@�GL鳭�ުn˱����;�������t��ES��)V,	�����ms��HgH�'K�5i.
ץӐ��e�au�q�#��	���
�W.��-iƪcfe��k�uP�	���(N ����U�2zX[�=�=�5���������=��4�6^Ѳ�b����G0�Xr�L[��y�`+�r���˔��~aTe
&�q!�U��oVo��7;�Q��49�`�s���Ali&H��	�eѬ�v��WB�=�;�ZM5���o>����kv%��ש�E�Gυj��c���e,s�?y	�e������G]c"�����r�^~��ė��2�&���q�x��[	��o� ��1��)���Z��;ݤP.�>���bu��YX"�M[(� ꜆ �����`=����I��瓱�##��1f��=N�T0���w�1I��J.��)�b�v��.X��?K�g5�5�,�ԌY��A��p��4(f,�9n��	�a�p�w�Ut=Z�O�iAb���L4l(&�f1��9��a��"���������zz�M�������'h]��Q������E[��e�l�v�`�^�Q���9�����k|�<�4ں��;��<h��[�z�]���Z�wY��Fw*`���� ����Ez�|`������Os������o��K���@هݖ�����̾Kp̴��j�r�G��27L��(E)��oV�j^���9 +KޯI~��հ�c�W^�9����E��{�<Ѣ���	�CR�̤\�̅wWӈ�[;+`۝��Q�:��"�+&_�G7�⻐�avv9���տ��j5mh��ڵ��>~���>�%.�N�_�&m�ҔĆQ��c��qɈ��w%�ы�K�j���d�6H�\`n�E�zy�+N���y�{��~�V�v�������Iƚe�:"ص�!���զ��,�F�kn���
����ָ���/bv3],h<��m�/���4$#�[<vM0)�ͫ�����z��~B9������{d����y9�-5�v]D}u;\~�w��������ф�$����̀P����\��t�������cǔ����`����^�ar�����ޤ�PJHb�-�m	���i���P������E��q���nxiI��"X���l��z��a����!"%6߹J��)��t��V��[�z��q��J��y�7��t�.�uL����@��"<[���N�D�/`$��\�I��;��?UI���/��'k�њ�˝פ(^�fK�`���A/���xN���T	bWIje+qyGg�����mC���d��a+�z���� �f����{�>�)�HiRO��Rr���$U�>�K���P����'�~{��vGN��-(oja�7x��Z���!�²���t�4Җ��墌�V�[���>��d�s���Ct���-�t���\����v��#0�Wk�5󨋑��]�1��n�f�]?�L��pY�ow��Y�[U�鍶Ƶj-VǼ<7��G7�J�x��G2� v�j�����}��
A�9�jvx7W��ڋ߰�s�=����^���W��l>s־���	u��wM0�=!�e�4�A��i�#\H׆\�x4baRNL�#LU���R�&�u��xV�kzJ;��O���v��gal�w:"�eL28���2�&w�Br�'�dS	�k�2��b0i�ҟB��l��wf���ڽ}I��1���}����!�D;'��=ϴ3�VJa�����˧զ@y�ХOh)3@�вE\7�h��6WM���iO������>@+Y�;�P��4���`���tQ�.�xT�@��/�_n��qs!΅�j=�q�� h�gh�"ac���d�oo�G={N��υ��6���<��T�v֞���������C`�|F�����N6ۑl�Ë��O��M6�ِg9��y9��5}'���dyv�|kO\�o�ȧ|�R�6qS�l7�U	�u�;�Z�P�n��ϫ/6+Z�[rb��Hj�Fu���8�S:|��|���!PW��?߿42�%��A�tr���3��GK=Hf��:�����\g�����,GJ�z: �R]W҈��x��`����6)2ۙyDEǇQ�OI�%�7�mi69��{Z���B��WQ~�����4��2C��q��Wk�n��7q����m3x�
W+�(�� D ��*���6��V����?=��>�a�l��{����L:沁W�جj���Z��	�8�:
��z:�������Dv��S]֦�p��@�����(	��i=:ɪ2=tB��QI��"W�
��f#!X޻�݋�S.W+���5uo
p?���M�?�F�a</���_�2N���m��i���R�y2suP_ܺ��UE8���a=�m� o`�i��C,��|�`�WYf�&u姫slWd�qvEWV�c(	���"��D�6���[���F4�r񽻨�2*z��k�"Wwj�b�-�T�m���oܦ7��	�m�o4���\�%�r ���>����m�ɼ�^z���t!�2�=�`ԉ;�4�UfW<5��^y),i�a!<;�eŖw�M�T�Ď��u�]���sj`���^���ՃWB��A�G\f*�
�<�oԫe�nNj�7RkrK��΅��M �P ����<H|QC����q���L�[��]+_.ܶy�T�ٗ��;/l�&8���<�{�a���a�i�����a�m������m�T�j��8`���W:��g�n��3S;+�T	y$��Sv�L��j�T;R-��-���o_D��_r̡����o��C�Qp1kKi��I�(�ު��Vj��k�o����-<��GE�*���0�2��7��C�[v!��u����~;�������M�V�*��6��֢�k���*ֿ������<^%uf� ~e�X�T;NW���,�+z~�.AP��!�������i�6�{`�X�t\��"��t�o��y����C��v=f]���m�tg/<����ub1����V�5�ӡ<��F1Y��:�,��� ��RPiG�|pE�����/�{ވ���#��kFm���'��1&��Y�~[�S�Vo6=f�A�� \������,��'�MJ��S�;`���\:O,�0Aa�q�/���j�Ɇ���Bװvd�3���������";;�H�CMp��6�}skb��t������-�d�v�����p��(���jﷂ�<`kr
OaWm�Ӛ��O~��v�[O���!�C���:��J�lr�c���^���VJjA�xNx�LPRU�7�Z��	��=!��9�4G^��՝��uS�8e:T�-�^�M�O�̤�x��b�ϩܮ��>�s���Of2�c�e����a>v-h�ڽ�w=	�!�xa%W��w�f):a�aK��LkSߟ��鮥"�yvγ��ǆ:�^�*��;vl� ��E�/K.� �$�P�#&'WZg\[�J�d��l���f��>�Q]j�Q�i��=��Uɕ�M�n�t��׷.��X���f�����B�R��л��zQ��s����9�Ma9gq���~Ow���������V��Z0���a� �Q�xGucj�yo���8zd�cl0���>	�b��ة;���YU��-E��g�
qqى�ښ��/����m�`������G�<:mi���'f�����rE=4�����W�gzƯ�}�9<:܂\͊T;����^V�c�������?j��;4ژr���ٽC�Ut��mb����(#ҵ�r^�ȥ�Գm{��?O�C�s�w�}he�HUTfgN����b7H�h|dl;,z���؂�1�2����ӎLG6��K1/A����;��U�1���2%��AС�0�؝�Oٰ�E��`a�Ao3︴�&+���,r��9$#�B��E���XQ��8N�/�$��3e�ӱ��ggٵ��r���M[����k��̧�w�{uC!�����T?P��g�D����__��Q��w�4�&��f���e����O3}�a��h;C�x��-y6�������~�
c��?����/\��s��{Q1���%��Eg��k;�2��LܶdVN0-)���i�cռ*�H�x[Xd^���\zj�u#/�L5�;���|�������ۚ��ӶK�Gr	��U�����:���5d�Ȝ���Ó'n5~y,��۽�T:�ʚ��.�o-��8��JeCw�w)�Q��+7Zm���{y�<�Y�n�,ĩ��Y;f;'����F��_�W��UUVѵb��U�j�Fڲox{�WgOh�m�����Gj���mQ`��ڊ�o!)��)�4Ji=���O�r�]B�_P�=�wO� ~�> ��՛ՍO��-
,T���`�Ѵ���D �W(�E�$��B2�������j�eFm�D�m0o��T�۪}w�%D�e	xL_	H��^�DJt�D�7�R)�m�l��X�d������H��-L�\�S�\9��@.�mB�m���ʽ�Y��,�w�of�V���N�o���0��9���9�(��a���az��y��l+�!�"mzvx7Vt�QxX�Z�1,\^�Z�8�lv\�rv@�-���O��%��ܺi�I���'X`���t�ݹ�`�:���W��v�/�yק�i�N5p�(�Z��a�(�zO��O�q"��D?���1�:�ϕZ�����vV�����	��ubL�c^�j��2��b0i�ҟG�L�f�;�i�J;b��i:���uf�٤y��>��>\^��?>�q�jà%0�c��t�����f	�����Zp��[Ngl���Ch4rk �����/��~k�yzr����9B:���pB1,y��G
[��V�U�-�2����K���ິ� 5����o��ͩխen�w�`��Nu�6m)��]M@��ضJ�f��,�5�(�X��jb=C�;�nQ��A][�{,����9�65W���G~f�}V�V��SS8*lfN��9�3�< 0�����3kcZ�+lU��T[m���r���̅��*(�'�nZ�{�<3ǴG3�
LL,s~�����z����N���ښz�����k�~�菌�>HOhw�\���`�|��.9�'Q:���3�N��m�ݤ��5O�^Z�i��O;PJq�j��6�֟�)��"���	鶋U���������KBv/�mК���Zݮ�q�91j�Y$5$g{��:�\���9�6X4k�*Uϫh���X�#`d��ݳX��	_�b������vOAd	c^+�Y�_(�g��K�w��lZ�~k�)�]��`���.Xs�2�s����(�ώ����+t9E'U��i�R�
�X4�!��t�Wߵ���e�|�G��X
D�(2�pΓ��f�7Ҙ�Z�bCt�?N���W}����c�*�U��� �v_����������~Ǥ�ow@�78�����Qo�o���7�V˴�F� \&)�^�&�s]��ᆍ���۴U'�o��:�ץ=����WE�#]��E1����lԤ�|��Y�09�b摴zk���3��D�|ޏW�������x�}��o���뚀XS�Ͱ������[��]�n�霫�wbC0-��̼i�At�L<�Y�7�c�����]�Q����*ps5�wJ�V�������*�X���6K�ep)� D;7���5Z[Qܾ77���-��R�0>�:�΅;w���ǳ/j&�/1K�6anԓ5������R��3;�kg|�r�1Z��S�IaP��N࠯����!MA�tt:;"���cc�pq�gEq��vћ6�i��J���pB�t]���ݭ�����R�wWA��w�ٚ	��}O�.��5�fH�ѻ�Q}�Z]V͵Ӳk�Ǖ�(�C�VK]�DeG3i��{�N�S����3�0��\V3k:���`u�]�<���Ōf�[>J��}:
�KC�z�|���� {v���ikT�ʝO��n�G�P�刟�e ���S�&��e�5���PfL�qe�$�,mjQ�+˗u�s���5W/aU���KZZ㦌�)v���/�j��;�P��L����=\�;�~uh�j���7�wf�|&sa��ε[�j\,�_f�c
���j^%�h��]|q���X��iWČӲ�St/F�c3]��ΚrY�YE��:�� H����}x�B��v>��9yձ5	�{ڳ�T=�K�Օ�B J�,Һ��F�9�bHN�K��wg
�d�P9&m>����S��H�=�n���n`��������F�| i�t�N�v���K(E��o�z%��Ez�Rݛ�k��:�hgk�`���=TSo�Ӡ�˰����K�7S]�)J;�ȥɳ5;w�-��;��ﾷ>O�,�ɦS�u� �����ν�wI�`Z��
;�Y�~�w@J!?z=W��x�Q�]-L뚖�Pσ�K�Ē)�����]z�R���=�2Z5�#k�`33x����5�6q�l�Hh�����/�2��s|{�Iqu�gqj�vs��X6d)a�������%���ii!�=��_P�z��7&;Ù��7,�ybM9��+r�:�0���/�!�9��tZ��,.�w���ںy�xJ�����Z:��`�[Z�]�M\͎�u)Kn��A�����q �tm>�8ig�GA�6�����S��u�#]��*"H7:�]�s���u�u�j�NK�{��u�.�%^����/RgC�Ј4eg���C������b��'��js�}�9/
�A�h�DX��{z�1i�Z��nTq�gzYEu�51��ً��jӓ�bf;ʏkD���C�C�mGՈ��rV\p3,���(d�1Y1�r�cѽx�9��S�G�+ ��r�)����)�,"���*��
��q���%��Z�!5[�K�ҥ��b^-���!pq�� vtV�:8�����Pڸy%r^f
��\�0h�y)���te�]�x{0�<�>�Z�Q�{2�U�,>;:�1�\����;l�ЬNCL�yպ �1��J��}�/KkQ$����u2 �9,���Iӎ��$�ߥ�{� P T( ��!����\B1	%%F�^nǺ����;�wq"�D$f2IJ�%b�R�E�9�����d��%f"b��S�"ȉ�Ld!�@04$eg8���	P�� �)��$ �I��wt�A�&���B�� 0�3H�H,��$"iiID�� �%��#H	�D2cӼ�/�\�@A�4���f�E&�F*4���RD�Y%��6baH�	J`�Q�CIAwq�LHc(���d�L�H��HS4��d؂̓h؁(�(�$��0b4�L,�H`�Y�_���{��phuCC�s�Rh���2�H��V{V��ns��kf!��]\yQ��T�[��� J9�tI\�[��ڶ�����[E�E���ֱmh�h�m3[Qh��0�w�����k~zC�/>�A�����.lI�o&B̮xkT})=RX���Uek]8��7mT�̧!������ ��=ά�г~s'\]�TXU��c%���3���u3p�������V���X �5D-<`c����q�S�]����
�=ഴw����~��M�<�u�P��Br\p]by���s&�f!�3���6�L�y�f��1K���n���0���.�
�t�=�i��CƇ����`�Oނ$�y��h�l��.+�A�+��Jq�OK��7�.� a�,+�bK��]��L˴�C���,�)�%�2#��~��\�|v>ゾ��j�O�A��>��D�,^E��!�pC$za���e�4슣���\�L!�%����6�iĈ̔����f���H<��@�9YA�ώ���jo3N,=��̺�cP�:)�0Baa�qqw4^����KcR�!kŭ���<�vi�NR�n����5�9B�ޞ�~ޖD5�P���8��G;H[8� �\=C�����.��Jne<��H2�^W�ݺw�xB�/�V��t��vF'�q7�˗<W{�v����ٲ<��a�єl�i'M�G{����ċ��I�o��]�od�f�v���k���������+�B����{_k����W���.핥}�?����=���U���h�E����m�IUb�b���6�cZ�m�m������|��~?_����ȷ7�ͷ�U劅'�����v^ix\(]S0��0~�����e܀�M��z;)bB�����<��Be��	NJ��1RU�#&������{����Y�N�ީ;�<�yp���ߚ�j^���E�i�I��YY� S(�aO�\⻫;mQ�6���ƚ�O]�*5鹐���$D����5�H�B�'yb���t�<S��wk݊�v4m��Nڅ§-^w���� a��:n��	�7B�N�{�Ut<�c��=cDF��-l阮q�r��\�~j	ĸx`>ϘG���M�pDs���Fb��+[�x=�T�m��}�-y%F�Gs��J�s���^/n;`8Aq�9�a����G�?�?�ݿ?��:ӑ��=������!uc]�PKܼ���u,��L���8h �y������aVI�.�N�����H��m��{�ln
���(�|�S�ǯ3�^;��hņv"��1u��a���l�Z�2*ǅ�I��"'�ߧa��lm���9����Šv�����q�.�w
]��7���\�)�{t��x�B�: p?}>�́i�jCZ0��|jM��q��q���:���cSۻ��꾬�i'9�#Y���97i��s�P/�O�v4�V	�vwm!jk
{4cN7Hٿ�񎷃���:n)(a�+��W�*���#[F��U�6�[Ej5V6��&�6�+��5Ƭj��Z����?�ϟ_���Ƶv���077�u�v�1.�1aCC�q"%M�hؽt��df�0R�� H9~��6���LN&��{���"��&����_��5��
c��a�~05gP�(i�z��V���0���r��(Ӭ8�����}y6���6����@X�ie��Bm���R��"jڹ�3�{i�������"�Of����'���C6q={��W	�[ݹDGC#��<4FV�y�=�9w��P^5X�z�b�>�BSe�5zҚOaWN0�>��9C<����G�K� �ݮ�;�~�u!@�"XvDA��� ��<��p�D�����ee5(��d�Q��/x}ޝ�~�\~Օ�'��'�NdP�*�A/���tD�I˼'$��#15�ޤQ:��m��B[P��Mmq�<����<�|�%L�m	��ʆf
�'p����:1��Q�w��t�����9X<�4���5�/O���=���1����+g�O]=X.�����]�����Zt�������	z\^GP]4�@~�4c 0�)�z���j�����8oߎ���G�CL�;c�22^>yע�7-�[��'��-l�7��x��ld��`y�+w�N���^H}cCw���O\2;3�G�R9Z��]	\�K��,��\w�F9SV��,�K��JUӇ!Z�6)h�:�w��91��^����{ު��jf�+PV(��+f��ֶ���m��>��?Ͽ��Vj�����&曯8ֵ��(�ZcO��庼m!��G�xQ����ti*hJs[^_����2}8�
�V$Ȧ5�&��L$��Y�G���TC6h�J�ΊU;E�O?cr�vi@T0g�� ��a�]�'�����hZe	����r�����l��*��#"D�>*m�����������,j ���ǃ��B��c��ޑ��K�P�kn�g�l�]=�7�����h�(���LZ���v|��сAg�X�=;#Y#�{�������X�I�A˯q�Bi)��C���w�F���~T9KOհD��^�|u���0���ɋ]��ާ�WV2�8;�є��k�d�%8�7#���5�=�碀ſ3Z��{��
��ϼ;j$-�U�B1�!�-���\�f�[+t��吃��Hj	�z͜e��jx7���5Y��4o�K��
+���F��ߔk1Q'$%ӱX��B|na�@�9U�}A����7oe:����VνЭ�eEÚ��f@���\d<s��Ӭ��d.z�c��եRѼ�U;2.%�C��ː��B����A��-���[�%L��R���ʭ+��ݷ�30nӁ��
�;$]����fg�9\'&H���;ns��,J�4���,�sT2K�����T8�AyKF��)��7�-9�#Ut�f�wZ?�� ~�O�Z)"�`ض�ɵk�>9!n��s�d���.�F�QaMAm�5u;k������̛�����s�>��=ܺ��� �^��-̂�-���%9��Jd���5��4-�oD�#}Pqq��D#�{�m��Vцl��v���&Y�0:�+�G3e�;�D1���-fʿ?��{����Z�N�����YU�N�fy�˜�09�{���=5��ZAwzTSi�kU'�g�AÖ�pp�ȇA�������t(��z̮xkU���D�L�h��s31�}����#JH��sb��X~�`������u`�гa̝qvE��r��U�Jwr��B��ݳ-r�L$WAi���L@���i��Oy�}�o��W�gAB�t����z�z�s��>��J����PK�]by���s&��3���"�s�)��W�oK��wiv���E�5{T��Mc�(v��q�x��s�^V
��iP��<�V��Īl=9Y���Bv	�99�	�v�����t�QaC�Iv��]��L˴��cC�Y^]���z�&���}��xk3y���Y"_��t�1��,!� %xݱ���\��@ 9B��Ez�v��{�����<x��!�
��k�\S��.��t�d��w/`{ۜ��R�Q���Ƽ���*��3�\�*\�s5��E�=���GN�}��oﶱcVجZ6�_>��_���Ͽ}5K��T	�by�ό(F��#��� ^E��CL�C�J�D6X�Êc
uGQ��^��1�R0��~���Z���W@�E�����^=���\��	����x����5�f���1�:dwr8k�o�����g��a�q".���cPbr���m�,M�t4����qy;]���%�7%�B�Ru��ޛa"�*��E|�7�?�|�U\�}�K�k��e�=���d�s*RE&���Ƃ�B��U�B���z����v@�3ib�:|��H�=ڃ�}S`���"��7:�xO�)�jRU�ɼz_r��(�ۧ^2�K��k1�ǝ�0�u�>W������D���L�N��K"�9��F�	p�Mt����wh�Œ�?\�t��!C6LA`��zcC�*��w�1I��*�]r�Q��u�]�[�W.�P܆Nܟ��k�mx��@(fƘ�	����H��i;�1a�-��o�������Z뜧,l.��A8�;�XG�<��k?�����u^b�U���=�~�ݠZy�t������_c92�i��U9x�wv�V�6�A��`�/Yͮ�d��*���S{ ��*�c ]�_�;r��}s8���ښ�s�|m��Ė=�+�̹��7�7Ҷ�9h,w�ow���&Z�������߿�����?�[J�-Q��+o �<=�3 =8��Fl]����]�.���i����w=,�|�ۇov�qA��A�G�N�z�������g����^Н�e�$�kd�M��r�Z�⠗�{��UԳmt[���f�S
�Z��gD+Uo�v{���ס�?3�n=oE2~R[������}8��sh�ܖb�P �fzr�[�Ï����!��S�4k	�y"�g�	�|��`Ge�E���=$=qh���������m۬9ڽ�=6�PwnC�]�[0��F����4�-�v3].2�v��
��f�L�F옂����s����Ty�`D�CH��k��5�1���?|1�Ƭ��Ӣ���-�g�UYI�Ud�)��ͦi�rK��������O����yg�������^v�ۗ��
/��"�w�c��{1E=�5>�z��ƥ�S7_���,�`Z�;A�ٳ����W�E;�r��d�O�5���c
v[*�����U�
�دN��9G��&"ҚO~Uӌ(zg'�n��	�wv{�Y%��m��϶E��^���`xaw耈y�A����D �P�Ƚ�% S'��	�Ee�C���Ś��-���vU�����q�HjWL��y���"U{tcy10�R�Q;�z3�u�m\����L�od#����g��W��ogNIfT���o��,Y�-ܘU��ulG�����Z������Yn�:����ƽ	F�ھ�o��Z-�5Q���y���� ���n�u��kp��ۚ���)��= ���.͕/	��/��'��K�'I�t�k�1�銫�w����i�r�Lk�Ml�Qͯ�p�������!\�y�v82�2�h�ey�$"�6�qc�g'�|�8@�����ީ�C�E�*��E���}�l!#<��t�Hb�J��]���Xb�-M�=��m)v�,�n�����	�����u�L$x�����O���4[-�̚\���C,e�8��~/�ri�8����BԍcIGsד��1.�s5=���9u{v��3�R��ȇb�jz�s���ƄW>{�2����J��Q�`��L��[�S�^g�kg��5�ю��O�0g����|�ȇmt^�����q�j��S�1�����v-��)����2�۸�x�������v���8���:���}l/Bv>�q��̗A��Ҷ�rﳞeu�.
�.�`S8��q��^\-xו����cC�>~08����U�j�ߦ+eX�������b݈gP~yŝBhq�.�aض��s���,�y���!�ǐq�y�A�����%��8�����B��H��y=���VX,��r�;���%��	K�ӽ�S��ʚ�5�@]^������������W���7Kg4c%Tyj91�e��9 /��q吆2hq]��":ڹ���;��8��U�92�e�{akJ��Q�t�~�& xy�{�y��{�)b��&iheM�������m����^Y�i��O;%�7.��?[�����n\a�P]dG-�m���#`N�L��S蚹殱��Ka ��A�QY$5 3�⺬tV_C4��Ќ�i�xՌU��t��H�)�1����K=[���'�8���;�&�}�[����mC;�Y��|jQp��fA8�"K�lq1<�>\�\���kf�1[�I����m��j!���Q\�j�(������T\:��g�[Р�5�:N�Y�&_������ͦ��ܙ�!�q�PQ�{"S��J"��qw6�{"�t�z �Dc\��}SU�`xW�_C�#����f����.��4�2��b�7H��≠lA�/A�-�n�>�b�wۼk�D)�#!=��/H��O3���zA�0��U�*���$��"��l\�6#n�K<�;3�۸�(\���n��^w�~yp����Cw=OE'6$�
7��
�fW<5W(��n�.�K5����m�U;�5{rC���2nw	��	�u`��y��s&�<��#�����>����+�j�������7Xa܆�ܔk�ǜL����-R׵�e�\c�L{Oc�F#�[H����M㢖pujW2aH�:s�*��'���kcĚ��ɀ�z�;�`�lMߕ:IB)�N����T��E�+�M�?����x � �ܹ)Qj���0�R�.j�碯񎎇\a���B������� L�����v�h��F-lؚ3��iA��8W�]+\�%鈕�@[Bu��ÿm@a���F�3�=Rp�S��w�;]2t3em�mS����jR�m�Mc�wh��R��@��^�9�dK�^5ܤ�(]-Y�kv�C��`�
l!� V�22�U�.݇$��q�.�aۭɈv�M��k�Wڦ���a���2�B��`�'�g�5<��{s���D1yC�i�P$=�Pe8�m�3��EOgk�	��]�����@�xc@lg�`L���c2R{�Ƕ��֑y���zx�	uܻ4L�2�	�K����R�i�8��o�2�5t���"�σD&a�
5��|:�⽍���;J��Һ��~[8��@�#��l ʼ�(QJN�~ӌ&㦽_��eH�#��Z�6�$}g�u�}oS�ՠ_�_�����=E6_.��1H>���vzs^��V���{gn�OP�z�Vm�ɚ-O��R��C�8���7�y�t!)���Nl)�j�]�ɼu��og������{}��w�����|�u�b�g9�z 0�~�7%��\���y�6'��U7��D٘�j�p$`˨�ް����i�԰���{��^) ޙ�UkH�4]&`�H���f�)r��R��hJ�����#z� p�u���rA�����Tf��u6���s�d	��'s:���@=|��L�Gq�{ ��m�@�d�)]Y�ذ�ne� �:6�3�d� ����b{E�՜w�vR�`]*�*����0�֊��a(�I13aވ�(~e�d�g7)�����G�wiӡ�ė��ye!v��C�:�D-�]݅�p��'֖W��J�;���v{�ظi�)j�A_��z�%�³�2���w��LVY|o2��C�]��J�&jʵ�j�p뇐��vާ/}�,gd�0.��!��C�[c,�W��m���|�]�Z�c��*E, ��b��껩&և3F	:�D�UA��sc��U�����h@�*�R��6�;r6g�^��Y5���v�i���e�b�:��.���A�=9Kc,f�c�C��fse���0�L�4��y��hU̡0�I�� D&n�n�H\�-@C�ŭؾ�Z"�w�y����@Y�Pll�����݀�1�˸#�}�XP!5M������4���֖�Z�@{���v�B��:�jD�}{B�R�+36I��z��U�m��=m\p ��u�]<���wZ�3ufE�̘�HD��N�V끂���z��;-�hō$�޸w���`���p]��41�J��C�\}iH��!�ki��u�=�7��]gz$��:9�b=���.�&�_w.�B�D,�੾Dw[�+�]��w��(��'�n�ZHCK�=Wb�9�q1��g\1)xMa�<r^�������7훑�˛S^��رY��h���d��}�&�A�,4������l�˭��$�EJH��;R��qF�y��4�ʌ����Wu�4s����m����U���&�(c$h�I�R���Z�*���J�dk[el�g�ȸri
;�;�s�ey���x�<0N{�wA+��b�,m�V��l�u�[-o`k�eU�*5;ר$d��j�v�qg^r��E/kX���(�v�/�_.��e�)֭��R6��es}��� r�w4��͓m��ܡ��U�v%��-�����N��o�:6Mi�,�݆.Q�C�O�ij�k|A���7�f�)I��۱���xh܂ɩ*��$ە� ���`x5y��D�����{eg+��հm =�N:��ҜU2��=YV���oK���*_���0����&Q�U.l�m,��_�=��MZ,gP�V΂i��Y�5V��k�'v�\�4l�{�t����Y<P�&�w����mC�e!��[��̛X�6�Fs�h
��(�`����G�v�;p#*�]VdY �A �B?�$S()SF�c��f1��0��C��D���feBa�2&��KA�#.v3$��$R��d��q�*A)��L�"T�0�SdPD�QL�MF�Bh�c���M�h�L�C$,d$����;ILX�SQ����$4��i�4�!&LEcc"ȥ"R�2F����$���Bɉ"�I�F�l�̕�PQ�K%�		HS2i2X,�:S��5R	I��i-!I~W/9�c@l@a&ZLmː��;[���o���v_95��M�lԕ;5添[��-
kO%�M�:ںkE�B��m�_��:�Gl����d�r��>[�b��Z��H��>�P@�) ����U�xU A��;O���r�u�ƸKm$�-�����[�x���2!������B�צ��N��K"�9�|7	�7���; ��+��ՊX'Q\����}h3c�`����C�$J�4��R}`ՙ�׼2cAF�{7	m�y9�j���c^�u#�]���:������~|Ǩ	�	�a�f�x��Lw�3��Ӽ��{�w�U��j-?1NX��L?5�\;��C�ߏ�J����.�(�u����o��j�r���a�@bYB��0��ut��u}�1�*A>��v�l�u�:r��t��R����S��M�:KS.��r�X�⠗�{���� ��K.鉦��u����t���1�G6	�v�z��W�*��(�|�S�Ǣfy��̦�m�zǳ;f��r�dt�/��	���S�S�yX��˳XGt_O��ϟ��t(�ڑ��SA�>~�?>�Ow��
�W�.l[M�v��xA���Se�v3\��7��
:ZXμ�s��e�"�x-���hI=L�-�Mn���/>�>�Ƭ�����D�v�Xj��4��W_4Eo3W`M��f�!,���f7#��{٨�{����R��f�Q� �l�ʗR���^�W�Lsn1a������v�bV�t1dY7�^�+ȷt���-���_+x�ie�B�掠���p��R	���\?Ͼ���æ�u�x�Q�q���*�3p�4��XrW!�%�<���R�3T*��ɦ/��h�}w>����C"�E��Ș��ٜj�S7Y�A�yd�ԑ���F=[����АCE��}�XX�Y�`�C�Pq�C�y��IV0J�'b�#x�M��R�&�ZSI��Uӌ�T[d�T�e]��#y�z��[ռ��|�@��"X\� "Wl�(d�殈A8��!z�ˡ�0���t������Ƈ���O�Sj]E����|j���Qm��"�d����@K�`���A}$�Ew/�.ol�l�殦�7}���:�s`j�Lhi5����S�\:���̛0?���������+�������X���L��S��BTi'�b)9\�$��\Ø��}���a��wM��;k�;����sڙ�M_HZ܄��^�ڋ�¥�}ft?'���y�{yH���@~i�r�:�Sm{��y��N��-�ƾ�z��+�r�g}0�g��N����Q����A�.�z�`����Z��}��S�}�ga�fB�0t^}�ʩ4+���,\����2��_�6�^Tp�?�f��c�^oK�Gt���,�,j���O�,$�|`�'�,�~���p�u�t�&o9��N<,w	�8�;q_]P��Vc[[8�����BH�7�Y���\������k���:n^N�\7i])٧b�2��k�W���������v��T�����d����'f��|ycGW�T'�����VJa�]���\.�['���:���[��%>��Q\�����C�O��+B��ӞT&���>�I�G��9�:{'G3�U��[#4½ŠvW�j�~���;��}��9d�g`cA�*�.voP|�Ӓ����o�z�z:4�ȝ��4]�ñm�������y��[7�~Ϊ�l,���|��c1�۬i��D�.��Ӎ��z=޼�L�^�'��%8�5r2�m�I��8Kb󍛸��p{xr�x�r)�4l	��aql�ؚ��u��kR�H8����CHK1U�	��{�n��l�r�>�b��Aʒb��Z�(�⣿��N�EG��.��s�[b@�50ȧ����]����-Մ���o�YQp��3_�
ȱ\d<s��Ӭ����L�S��9�Vp�Ó܏:�Qǰ�RukU
W�TXSW���PꋇT.1�C��(2�r��e��p�I�,��9�K��,�,�b�:!2Of"S���EU��:`��b�~}x<<=��x��	1��V�$FQ]:��ʒ'�b�'5��"�>y��t|:�C	�¼�W��h������AAl�=���s:�� �[��V��[*¸��9O:�7A�NQ�Zsӡ�9F���v�a��@:�Q�t�Y�'�9�GU̱�W��ϠZ��>L�8�FF�T/����H�]��iRd�� �"��(����6�/U{_.���b�˭��=O��i�9�:�jq"��ʧi�R����:.�5��Z��=��Nە�gz��Ŋh�yܳ�ˇ�� �kϡ�n�=�ؓt(��{�es�6�n�i�T_���Fr��Gv���&S*GjHO���><�|m�&�7�=ά�в�&m�ޜD)��֎5Ϝ�8�����G1�J���O����
OB�1�?������^S	�����{�P�(g��V8�?��'����P����p�3c�І6��7|�QH�el��9��n��XsV��.�ǿr�i��F������XWy��~;�ΰj������4���V�RomsƏ�_{z#���e�ى.��]��3.�Гlb-T!����z��Vi���,YX��O��ϡ�>0�ۜdsz��^E��ZdQٳ�Qt��O7��Pnވd�T9�L��x<ă���,���D�x�+5h~��>�@X���u,t_c���Z���?Z��b�ֽR�Яz�bnW]�C�cqh���˝�V�T$�ej���lI�������$���h�xi��@�3���Y�to]�N *���Aa���"Lց�;KkZ��N;W�7�yͮ�Z-fI�vӶ�����r-������p�}>�Ly�s��Y!
�y��-�WL\:�{ ��,:N'�w4_zcC�T�iF2+i�_q-�0��d-s��"�(Q������	��c[�BksޝI�%�Ċ����<���Ȳ�)�A��޹ږ殄%6_)	�yb�I�ʻh]���{��z��ˡ���wu23Q�Y2���q<(LBo��4��<�B�Yx��L���gf��Te]��n����W�}nq��)ZLE.�V�<��oW���\�/����sن��\k�4,��-�;����`
�?�Z`�'-�������p���w�����hy5ؓ����E����8�ƧU�i�ϩx�@� у࡛}!7T��S�O9���fm��Xk�P��y�M;�E�沠���Z���Af���~:vw����]��Y�g9񃃍��SI��Ͱ-�܊��Q��M��s8)P%�� sH�����8�<�ǭ�b�/���kK����/0�� ��?P��m7=E�����	�ҵ���q~�����zf��ԲG����fs4Ս�u�v�#�]oW��z���[W �.Y�n�"{�̝�1N�"�.��V:�I�RnDR���Dy�f�����2?�}Q�[}��d��������f�Cq�>j�غ�>�V��sVV�e���ѨY�BHk��R+��s�s6�\?�/ϷOes�;�D*�\��xAO"��>;����WRcl����)�㜣��Ԏמn�p)�ŝ��j�fA0zK�m�`<{D"�ѯ����Lжz��d����l�mW���>�����W��D[�:=ba��wA�
��\<(��'c5�9�,��m�x���r���r���0�z�X��S0yh��n��L���~0���[��,L.4�m�u����bv�xע���hsO�qS4�d�^K(!��}�i��z�[9�"���;��S`E��[�9�FS�5>�-�^��R䩛������$v��͜Nj���F}�SWA7O����P�����=a�<�ǧ�U��دH�Jl�2ciI������ڦ1m#upu�j��u^y��5�1��O�D��pH{�Aᒫ��!㲚u��be�a�i�Y�KW:��c~�i �b#��s�:y�=�Ǥ>
$�6P�+� ��x�z�QiC`�����`�N�%הD��|
"S��"�׊5�A���(<��\�U|������|���/��~YD��l ��U��[S0Do��V�+Tu6<f��H^T�u)����X�V�,��*+	'�� ��䭰��U����Tڏ���,�rh�0��d���CWg8��^�%�J;p��u��y�X�#�ֈOF�b/nk{�#z�e4��i�ƌ3^�)�H�J�|1���F�W0��/^��y�|�-�@/��z�;��ҹgc<nӝ��D&����tSI{*��M���-?$�	s��r�+m�c0�8�e����k�'�!���Ƽ9�~�s�i����Z���BԍcIGs�u��[����Ή��9��	��,k҈c���;'+}&�ۓ"��V�ze'�cY�� Sh��=��U�K���J�;GN}v���~`uHNP�i�Y�y����;k��'�����hZ����2P���rWv7I���X�n=���VǼq����=2
B��||l5���Cj��欙N�0��:���؞�0��R��D�C�@���ͥ�[��<�$8������*�?��>�FLÕ�3ST��he,�c���H�*���Ý"h�J�5ވ������ʹKO�|�"�lUp�cS��5�b����8���Ai1���m���z��3M�O;PJq�j�eٵ�eD�w���b�sͅ�ז�P�)'�1=�zF,xo�ī���5ֵ �(�����`(�*r�͑��w*��LV�b���`�/Skht�ӂ��@�Oط-��Z�����u��lˣK#����+�����>�Q������E\��ܮu��蘆�w9K�ŗy�7�G8v�2c�rj����*IY�����̽+{�!�9$���W���mRe_�YVW˟���+��5���	���u�s�n)� ��붻Q�J8�@@�5⺱��c��*.и�'^�\d<s��gKvd��*N^�~�<ݔ{Qngײ�߃t9E'V�P�j�����8�/P�.1�="{�6T���͗�Ύ�*{��3j��,v��f"E��-]�L��1��F������[�S�m	��z�)*�אn.o@����C�#`�W��CWvΕ%��	�K�D�4N�Q�T���q��o=���];��0�r�i�!?)2O��Km���L�O;�m�u���Zr�v�[<R��o!�}ō����%�r��V_�j���=ʄ�Rs�I��I�������g�S�}���-W=�6<��4چ	�ݛq��>6�M�"n/^���Ne�x
�vUVn�ػU�HiN����J�
�OK��H��WAi�V�z�����B�Ǭ6N�Hm��H��=����xN�MՅP�~u+u�˥k�*	{hO�H�n�+	w E�_���V|W!Q���!�{��VP�A�Wx�������F'���I0`�m9qJ���������17�h��@P�=�)���Mp0,�=�p:p#)#�K�ط���7�2־��!��µ:������hZd�eG3�r+�,��F��k�,nU^37�r����(��tr�@�/}��v;C:�j
T��~N��j[��@��*���Md��Nk��TyUI��c���&��X�����ވ�9E������4���*:+ ���,ċ�lS��ڝ��[u���חx<�,"�T��a���"�w৬sx%�9�z��W���ڄ�t8����w�3�
���Zg��N ��;�2}��Ƕ�l܅�Z��fF�CoVB�2�ZX���d�9�h��t�:b���g�兆I��k����b���}��uצ�Z�2a��q���� ʂ̡^��}^��K���k���u#���n�DA[N`��?qm����#��-�dck�-ͽJm�T�ʼ�P��vл�5�{��V�R�5�?>Ѻ�Y/���v�ҜI�0���7�y��҅&Vħ6T�	��n��%���/l-����hZ��λ[�zkw�Hqm	���O��@"�ϳ�fRt��K*��/+v��'~�9��W9A<SH��R�[����ʹqpk''��#�T6��XD�Q����x,A�x�CV�d�fc���+Kav���W�8.*|�lL#-���7�O��r^Hf��<�������ǫ=p�������񶸌�:�2�����·k����u}
�η�W%{S�K��Vk۸�P�Y�:�=T���$���y�'�s;�{�.�����3��ynCS�Q��,�^���N͏���	�gB�4Dt����M�w��c}R'W��w�Ut=Qi���.��A8�O�GS���-�1G����n�Gd�N�e���&T'f���L���'(]�Ta�֣��zYH�~ sO�Ӈ}�q��ė�۷�j�����蕎���,;��N��6%�h�����%X¹t�{A/r�1�ٚ�75a�7��|��gM�f��l'd0d9������c!�q�ޛeb
���GS�cQ�l��z�����h����^�t��e��LXgb\3W��S�SVyX��˨f����xJO��W���oiU�<�e�#.P�ӡ要�@�:"طPwc��t���ā���e�ڗ�Fh|�QjM�nO�ߒu�d9�ٵ�!�i�C��A=0����5Վ��?w7G��TL�闚���/(�e���x�z[�C�sp�4�Aj�w%�J8z����6��U\���{��B뜬��Ռ��DkKhO��FFS���O=^��y�S,��eK"����R�j�V���Yp�-۸e�Y{���M�uR-�oǳ5e-����zۥ/\�L36���k�W2�f!dl>9L�7G�,s�t�����7'J;��6���D���h�oMc�**�%��_h�a�N�[�SA�.e��t{�5�Ap�Ӟ�]Ўd����U��oj"=�;)pu�Z�f0��5gg7R���6f��.3} ��ak�p˰��e'xe\�*�÷CX���e��'`�n�Iʙ/�	�4�`�N�f�/�{��6�C�'ㅳr�+���o��w�	��X)i�� ޾�NF�w+uN:���ib>!A���\K�f���W()w6�dx"����s:	�j6lS�4�r��b�T(����f��h(Tg��I�[b��en=�w�
�X�T�㤫:f��RN�� k�t;�<�˫!n�IoE�kLW��j^��Wn��<������'�N���M�ܓ�$t]X�,'[����[�@��[���D�]b�1ci�f���>�����?�npF�HV�^R"�ef6���45���D�l]�Mj�*�^����g/+�H�5�&2Z�WcYj���k�腗�e'L�����c��J��b�բ����FPZ�SA�Y�/m;�iƫ��x,�IԩLU�|S��9V��ζ��p`.��5հ�&����]�
��}Iq�i���2O&,$��#������Q�]�q�\�=��bfŕY���	Us3I�ŚpuЙӦ��WǨ�h�T^��c�GJ� |��$�V0G'i)�K:�廤��pZ�(<���k����z�]����8k�X��U���[���_����9�����]��ran�)Q���������,��d˕P��O��s��K�
&�ܘ�h[鄤��c�cV0�tN�:U�;{IJ&i�@�|�-��R���,k8�H���	�W*��N7�SW7���M2_vj8���y`9��L�b�TӰ��������ܣW&s��vC���,%#Sk�2#ˮ�Qӟ��U�����. ZL�*�����=�^�| ��������.5�76I'J�py���a���N��k���5)�n,�V���r�7�R|�u�q�CUp��5{g>+L�>��9�^��l��;ٙ��Z��]�1�혺:��b���QN�c���a�	OI���[,�t�]�s��+)RD�{�4a��]j��T�K(c��6B���)�-i�߮XFXy�����}&S$�c�B��!]���ViΥ:����۳73(�@hHku�e�W������ejk"p�:��!�ٱ�}�đv>��9��e	��q��wI{H�aI;�h���	�����m�#u���Ydf�1dGD�xa�H5x%�b�i�8V���U��,�y�t���)����}�[����Bn]Z�ڊ��sgPCtbu��n���3;7�L5``��/���PU�ag��m 9�˝�j�7�����^�������h�1 DDTm���6�����Zf�bSii�#%
BI����D(i(D�D�0E2Lȧu��E�� �I��wp16M�!�����nr�hԔHb���G��ēKD��4��vb�l@h�B -F�E6B��XѨ��+0a�X�;�3@���[��eE B[0����64LiD�,�����F����j,����I��[J2�Y�
������6M�Ŋ4d�!HQ�Dh���>�ofC|V�����̮��	�����.l�k������7�pV�7�4���e;���m�Δ�|ZGz��]snI+ʫ���៿d�T>1�`|O Eǧ�x*�`��دO����c��ɢ�f�,g7]�tX�����z����a^=�V�o��P2}�%�� ���Ed���3�Tm�O��غ�K7}��p���{�Ji��4��o�a����JV�y���<�ʉ�B͝��A��m�"�껩�;�B� azQ]'�b%9�j�Lh�I��F��P|��\�����)�SL�4r�u��s���I���,æ̧q>�J�| �Rr��E�\Ú�E�����TŠ�=(P�z�Zv/�aC�yЍm����Y�mI�v�M��(���@%����.�p�w����X1,mՌ'>��LkL9�}˞���7_��k^E�n�wf����=o�3��N<�;��ׁt�;��5�
!���Ѕܑ?.�N�\���Ȧ5�&��ز��u�B���٬����.JU�خ�W�]K6и�vm�`�B���P4u}�S��#�o�U�ɲ{%kwD���CJu<�S(�X�˧զ^y�����; �q��<!	�g�ֽ���&h�V�~<�ުW�b�՗�؍`���qHu5��_?�Y��vV�VsU�ۚ��x0�9cg:�e���בjb4n�NLne�C3�֞��x�������!����\W7xۻ]
���(��t�v�nu�0�^�.�1Bdx�]ݛ�GU��i�K��_̵��O�{
�FRpHdf�qg|^u�/�ܵ��!�{��:9��M[����c�fp+gd(G�u�]c�������χ:D��jeش�wtE��d�gH��V���
76���f~(�����0@v�.<:N�zq������f�d�Ql�![Ku��Vdټ�Y�{��c�tͼ/.�N��@�����x��7��q�:A�Mtya�j�5|�bmv���&���·6a���X9RV<�^IݳX\M�%����<C�C����v��wr�EA���	�z�	cEuc=�|l��s���P.��q�S�k��Tu_5���0]���b�# ��C,{���Z�R�TXS-��Ψ�u>�s�k��jO���?`���y�_D�W�e����ŨtBd���s�	*��N)�)��Vew��藽��j��M�y�!ƱHq1�C*��bo��H�J�,c1C�Ix�&�0�ro"�픶��&��C��6^��xa>܁#a�O�= ��\C-U;H{.*�z�?��|�;u��@�y�:�^.JزF3N��r�m�{z�M��.��*'�*�b7ι�xݶ�Wi��&��f��f�~ڔ{I�x V��֡Ĭ=gyt���#U��J��%	�6r.m�� �]�=��bn�en�-Z�e�d���9�)�U.��ԭ�hK����nqhXo���^Rץ�7�y��h	b��A�בCw=	����
%��N�M��Y��Ы'�Lxej����(�2ɤK�k,;��y!��'��{|��R�nзŽڪ��u]�u+\_$�h��\�ԫ�O��֠9��ǵ�!���]�$����sT�®Н�����2���	��"��u+p]��^��G0����P���[;�C��gUM;������0 �=~w��5��9�;.�k��XsaJA,�k��E���URтg ^���b�;f��}j���%�<�����@��+e�ӫ���rKbK�4e�7�͔*F��蚣���j�����g�sW��ߩ��&��ݡ=��ۜdw��n
jQ��#'��sR���p<���� ��CL��ou�5�0&P�.'�-�)9�kF��V��k�~d(֟^G ����#�+��.�1��[��t�ê�g��$H�²ݹ ׏q�������h��:��V%<5�*[����`����K2�	Q�^ޜa.:k����r�j�����Ep>��i�{y�JN��n�j	�9��z����;4h�n��vG�XJIeɒz�ESOI���\�}��)u;��[�-dhu��}�dD��2f��׹�6�nF^'/���j�+.|�W:.B����T䞎���M�Y�1Տwr=�Q9=��'���Bki�1�"Av�vq��	ږ��"�U�W��B����[�"
�^������M[��P���熟S�;@C��0�!�C��x��_)�t!)���)�c]r�d�&r"��Ά��܇��8������C��*�kb,�.�|�/ ��| 7ƽnX�z2�:�eN��u}�N9@�Kqu��)�z�(��W容

�?��9�2r ��}ʄ�C��r���Uu�����i^*��mEL,r�E�s�1�b�v��.[]�k�p��'fƅac�u�F��Y����B��9!7_�زśi;��iWC�zO��AcK���Rq.�}�����J�Z(����0{b��B5�lIu�f��'(]�Ta��w9��w=�9�����;��<F-�׶�q�S�S�@���W�9�Ꝛm�,��ame��k
 �JװT�.t�̄�~[Z��c��=ʙb�f���8�`0n �xB
wf�-~1�o����M��Rb��F7u\�p����Nn��z\�ӏ^�U�l�*;�@��#�84?��y��Y���������}n��P���.<^>s)joX�����~]��[k���(�a�׸�����.��N��Z�l*�m������SVI��;S�8̡�����L.�gyL�p� �����uU��侱�*�zhkwm���O��!��rw?X����9N���C�Zeb�t=1n���^�n`}��4���]5��FE��-О�Oǌ�'6��4�0H~,��'�A}���7�XlmJ<q�j�t����"L�����ZYX�-0�Ǟ�����ޡ�9�i�{ ���W ��o&��"-����~�kV^���ș�
P���|:O�#)�Lz9�׳8�%L�`��dY;WHf,�@�o웗���}�ǉ���}1|���W�E;�amV�����V�W�o)�{��0����NT�Jv;/Z:.������/�*3�=[�M<'�y�gx(���%�Ȉ���d�j��`�.��:��ܝ�<�� �p��"���ebQ��b#��s�:zkw�J�.͊{�"������]�e�BБ�}fQz�%:N]�9:�SIb�&����-��^;O���m)f�N-t���72�R��;=�ʆf
}fS��*R~ �Rr�sȣCsj=_&�7D$�bv�
�;u�guy�XAG�Ȏm����C:m�>��mO^���y<�]�y������SPy|iִ-������pjy��7��=�N� lm㠂��o���ǯ\��"�)asQul��h\4�����̄uq����
�-�u1�A����^�{���O9��:4�ǝ�1�u؝�U������O�N��Q��V����h{o�SD�:�)�4�~�q8�y?6r69eϞ�����p���E�n�e�?3=N}S��F���B��=��� s��H��j�.�?4~]��W/����PM��lK�9��;��w�����+��ޞ�'�~Ϸ���RD�k �< ���!�]��*dS�,l9U�Z�wv��+�	�}`:�è1���O�l��^[�~���G��gI	�Aq_T=��T��^~o�����v��@F�����ƭqU�hGPi'���0�ŠvW��sP/�ܵ�?����kKD����0�̍�ߘp��y�=��6>���/�>p�V�����t��{�d&z�/�����F��.����� ΋\o�W=8�ns7�ӛ������&�u��v7`��슎��Z�a�vV�֞���l�w�\E!���01����u�حh�%�::*v�Ŝڶc������������3�����T2���zw�O�B@�Hm�VT�o7z���ӿ?��~���جjA	���!��`q��Lo��}}�D֢?8����T���oz��u��k���{Y\�<��]�w����oYV<�o?{;�\�]r��7p�ܗ+ȑ�u�����a�6�i]��y���3^�Bd���swS�DyÊTu��		�oC8� |�V��`q��+e�ӊ�FO_6`��6�K�z)����7������)����:�g�n%&�#����?G)�6i�O�WD ���):���%2XK,���z�]A!靅tw�Y犯w�Wߠ�Bm����poH���<��'.�I2(���qqw���s�*|-܌��(��AK��B�P�#`�T/����_v���&X�b�$%�W{4"!V�|����"y�w*������q��#a�O�= ���0%�*���j:�'�[�u��N�؝�W#zѧ�9M�.��i��#}�rԸ�S�
���C�S�^�P����wS�o������ZjTy�lgԽ<eѣ^Z�E�q%�G�HO����~�t%��*
e?�?tR��T_�Z�@NE'����s'\]��Qak����i|���Ɩ~/5��'=��F�2��5���ρ=>�Ӡ�q�jéX㭗J�)�zb%G0��'Y]w��3_kvWE��!�W��hl���zv]��u�R�K.�ǎP�7�ϫ���w���f���ne����W��J�0�����k]`L���^��t�9E��y+�7ޞ����7/$��sJ�ɨ{;�X���W\�	��C&gl���ȥ$���Y�A����]�rs�9<�zm]ꅫ�R�`J`�H\ո��w`��tj�Sjv��a�{����F���PN��94b��)P���C"��RvT���?.��.E!�f���o�8˶���1hT}���+��$���ߍW��S�����Q]�$\&�\1˓���ދ��ĸ��?%G��U�6�ƶ3���p�Q����;ʳx�!f:��b{kcZ@��A��~,��F��.2�5��u^�q�q��-\
N��po������
�� wr���Ԯr���r���� �eȓ�Q�t�=8��\��b�hn���j����3����?�h>G����M�x���LU�B��F��|��{�ﻳl�\�5�cռ55�����!�		��x���<�Є�]Y������s]x�1��F�֩��IT-�*����z�%k����P��e�c��e�oy�LQ�l1K'{���n>��%�u��Lh�I�y�+�P<��*�?4HP͎���uÙll|�r��7�6V1���҇�D��4��Y�N�X�R���zccS�.g�ɡ�x�x�^�T��_���Ou���?hbͬ�Xh��`OH�5�7B���*���zja?5���0�ܜK�~��ʏt�Vm&�w��:�e=�ugv����ˣM�X\:p���=I�I�c��M�%�Ѥ��W5��5gS2���Zj�4�6��&�����k��x6+�q3�����E!q\u��6#x�I[ˮ;���}.f��mۓ��"�"#��l�޸ꓰ���#ی��75���ؔ�D���	�>l0�ßQ��n��/Ϩ�X�w���	�gM�,���ǳ`8A����8s��'f�U��-l�BU��C�J׬���qs��?#�S�A蟙��6	{�.�B߿_A�s	��F���x��[��w��=�].��'�7��A�t�aQ��&#���1a��qN��������֪�Lt_��~d'�u��{�֐��c��8��b��DS���\I���������ru�m}���B'�s��f�X8�s>ͬa���ZOT1m���7C�t�������xU�������GT��H�ii�{nO^��ǳ�#[�p�4�AaܖPB��aW4�sKFS���Q�����y��-���de9�������w��UL�geI�ӱ�U�kڜQ��TGN�r��ĝ���i���WH�x[G�:/".=<�0K�b����L�w欝������WolI���Ab�O~U��=[෫x/^��xA@�-��ޱ�܍�^�����s1��X卭,V�d�l���T�V4�"�9m*��:�2:�j�#���-`E|lN+�.��cBSnt4\��x���]��oa<ð�����p�sb�H���̹*��f�j"2_M���Z���W���lfQ#��o!�b��D�W(�E�%4��bQ�Ց���L���@�``SL �2$gCS)��zjw�>�6�/	�U�E��:"S���)͍R)�FUyٻ�8۷����8��➜x�٢,ƽ�(��!l����c^�,�N��(�T��yNV�	効�5�;���T�~J�͖ϴov��d_ ��^�;!��z�M�'g�u��cY|�S�c��z����:����c�*욻l\{�<�;�x��^���(��a�Ϙ(֘r9��Ĳ玨���8ԣ}by@+�V���7܎�Y����(�zO���v��g`��`vy��<���F嬽����3��3��
ݭ��F�P�.ri�#%?6#�eG��US6VŻ�l�����~.�)Cq�J��6�a���C���:~��R�c�¤ì1�e�d����7������X�b]�K���7{��,�P�ni�M��Nç��";���pl23L+�Ze1\��-x�gƺg�ߎdڿ�����&SCҋ�s�?b����J��^1Z�КM'j�.Ÿ���v��M�]Ye��e�]\�V1kͭkoM�����;�-}@汖�u�dI{t�\�w1�|ە�R����f䕋L��z��Wƹ�S/i�D�ė3���(ej��u2��:�k ]Ʀ%H�Vs�V܋��"�=u�7y���Kd)�1o���aѣd��ӃSS��}����em�o[F��(V����ʜ_C4R��8f�J��(�6�w��;��<pG�hz���bep�*T0'c�_��X���x�mŬGk	��y�`5�Noz)�qO}��	��eh�����ޝ�dn}�{��6̭񣷧<Ǘ�!��93�����X�-�ӗCya'���]�.�Y
N�tD��S*r6]��WNd��ޙv���t���u��eXw�KNw_=��$�-u<��X�$^��hgmD����6}���u��F8�����N�p�Z�����E`.ެ�."�;yWA��.�uj��^4[��i�;k2� :��죉�=����S�d+w{�M\L��8:�!Z�n��m>�+ny��p�[�9�\+t�݋��\j�kt�G��B�$G:�[��#���ţQ�^�O�%��1WC�A�&�����¤�]����*�6KO���jK�.�3�E��[��7�mA{�{=���-��	Lq!XT�Ǯ��1݆�GY��r�S݆�ݛ�=~�j�䓋X�K�Ϙ�ڀcT�����6���f�F-wAa�c��J�F��޹xe������N*�֭����9��b��KC�Y�}��P��V�{���v��Ah9A�C��6?^�4=�Ֆł�ǁfr��;W٧!��L����	�K���[��ƞ�k���V����[��p}Е�_ZN��u8����N��ɭ��t�q9�ۘr���i�vl��:[�k�p��a�m��c�3��-�n�G,��]nJ��w�ӧ]~�~�W�a�N����>V�6��61\�F�ۛ�ҹ�^,P���҆e)�P����Z�	��59���-ʑ��oV=��
x�y����y��uS�lgӴs�9FS�ӲvZ�2�Up����;����XD�.��q����pP�JuJ�7�c3���1Wr0ʝ���@ɽg�w+H�;���bP<�L�A�JN)�ۗ2U�a��2�NH*�W �ja�*�w^��{.I������v���d�dY�1��Z9��f<'mb��רZ�]Ѯy��]>��n�g9Dqr�ܜz��X�����I���	k㊤��7���D;PQ�f�Wu���m^S��.ݲ�#}[�%����L��`��٘�Z�@��h��R��zvq��j��b���0�\�q�� ��i�n�:�-[e�]\,��Z��c.}}}j�3+b�1�p��:GA�.��OS�H;Y&-m[�z��Cg8�]����e/I��M�����}=���q��qj�Ftt�T6`�U���ֶs��wt9���8vE��Ⴌ�Ni[~e�m+����D��T!��Qa ��04�K�]1b"Th�Hl� ����*��,�,��aBP�ʍ/5�B���$��a5��JA�T�DC-��&%�b,0�Ĉh�*�M�"LXđb����%E�HVe��HI�f60��Yb2.��"�E����S4���Ɛ�ȉ�2�h�&�j2@c!�����@ذ�'u�h��bɼ��P�	���&<�v���NՒ��(�)��:U���e����淐ԇ_Gxd�A������M�7s�n��C���_A�&n��/�t�Y��� ��� ���5T���zķ�ş/t� �����C��B3�ͼ*"]��F{#���tD���u�z}yjY�}2�	���fY�e̹}��~�L:{ވ�ְ�ˋ���%�H���=!�X��ʹ���K�7�\��Ƥ׽V'zp�w+e�Q�R�A�Pd�ԑ�g͋e��Ξy����0:O�m�����r���Z����9#�1��A	��� �c�K+�Y�o�^ʋ�5�p�051S������K�q!j�N8ʘ�v�ӬZ���!X��):��P�j�����8�!�F�?����һo��|-�L@��c��MԼ$�^��n��LZ�D&I��Nm%B�m�Ax�Y�e"*�f�WUv���M��E�*�N7�B�0��C,�Y�k��liRe�l��ĸO�y镛�K_ �"��4�������}�<��"fO�= ���!��:p@�0�q�\��]�=ܝ�U=�7�f�X��3��ʃ�l�D�\�e��T��=��np~�w���vUݺf��I��e0�̮xj���^m),k��C	O�ۉb���t17G>�ņ�0���/�<˝�<�>�R�3�T @��\�u���mtz�!T(�f��,Ѝ\��u��"'�!��f����]�]40�V�@tu^�r.X%�Y�1vϳ�zM/YT�wSh��ʞ��$��$�4;eZu��mo�uޛ�T7�n���xܳ���{���yu����w���M]6��닞*�
�y�إZ�5�Zs����'�D�¥9�+-�{/�;~2��	`�8/�c�sgg�Ԭq�t,~(%�ң�>�̊hh�o��u�^gM�4�^þO�� !f������eՃ����C.�Ǐ.�>:����7N��;V�nc�+��̃"]�Á��x�����$�z�F�a�H���{�1=w��X%�:�@�v�z�F �F�g��a^Pj�?���C�$Z�ac9�j�i�����;lh��;�.�^E��!�(4�.:����e]ohk��h1�5J�7lJ�kݚC&&	О/�����M���"�T�; �z�K$!C��4���MC�1p�M�ȎOR�Re���u"5��Z��s4��cWd�5��B�:�2!fP�iQ�땼>��H�r�=tw�j��X|LS_WΊc�8�h>F}��|lM�y�t)��HL���4���J[!�v��:�mvP�=9�^ǫxi����[HN$�|a^h		���G2�z�v ��6���ۚGL��8�<��7EP`�r������_�(���u��5���>g�:v����2���Ýve�n\�ך��+�u�RsҔU�m�ݍ�Y����92ή�N�-���pˑ�?� �1mx�Vy�N���*�������=O�n�x~[w��u�ʔ�5yIT.�&�����	���0��'H>C8!>S����J=�d�욃�{�a��	L��x�E�3��K�خp�Q	���A�l�y��5r��=�����A���(��I���t�yT��=�Ʊu;u c��Pw�����!Q�M&,�Z�H�f,�?7d�ƽ��Q�)�OYU�����w��,mt�rՙgy�4�u����|�8u���/76��|n�٢��Ͱ-�܊�^U��^��c`��vd�Nr��t���܅�Ti	���@B5�Ha��p�_�N�6�����+����*z�e�N�Г=U�*o�;x�:��E�^�����;ʈ]��
�0���$N���h~�z�a���H&-j��;T�(B��VGS��N= L�5�,Ɓ��K�n��B/���rYȤ�N�v{��gfYo��I�N�f�vٵ(�[�����D�x�zb���z%����5��2�6ls�4�P~�����f�X8�s9��!��!���z��h���d�X������������E�7vT��|���O3Dʼ֪2k_G���R�9<H�;�q���;Y�n(����`��i��(���"���;�$Ӟ�Ǻ= /`�ۓ0���Lϥ,��4�ܩ�O�����V��X��t^̺k%郃����Ɩ�d��L=��>Ɔ��d&�{d��=�g�l�2�:;$��Bc;&]�ZӲD��r"f��o#V���Z�?46 �4�Nl	�����[`��nM�w_Z�������E�bl��!�3�9��N�z͜OX�o
��)�08���C��^�������	4���B�}|Hμ9=ܽ�DcZ	J���M'Sь4�^=z���c� �d�K͓z4w��0�_X�ᔬdy!�{ �&��܄�yD�/~IM2�F�]���Ʈ{gO"���zaN+�(b��z��~�Dr������`��}$�{�%:O��Jsz�SMl�Q̫
0��	�4���<��UC�z���S/Gt�mN�T0�0Va;�iRO�"����(����bʼ��*�v�JE�h�^�����,"�@@��9�a�6ཞj*�{���<�o�nq{��u�u�}�K]�%�y	=./#�t�	=�|�-��
5���s�6%�=��n��q5n�E���Y=ܩ�%(�U������ćA^���]C�k�"~]��@^ �'eD�l�T��Tݖ-�*vk�.���
�㣂�ͤ%��	�l��o"c[��ξB/���r/���Z�DǗZ�6����M�e8e�|��"��Yx��S9���p��l��Uʚ2�i����|HoL�hj�rTM��sM���R�%�>L��[6��n:j���T�P���M��F��L$�ֺ:�U)�l��wf�XC�r�<���k�Q�sZ�:����ͮK��~}��hZ�R�u1���ܺ}Ze�K���b]��V�Be���vc�0d =3��	�H������t��NЎ���pB1,4qh�^y�lJ�S�!�W�з����F�gl,��Þø�vyBgh�"ac������z���/)�v���X{9�k�^~-��svG/����\��Z���Z~��$��^�|�"a'W����s���=X��SU�ⷕ��gs{�3J���޿%�5x�i��*����6
I���$ߵ�����]4��c7��y��������+Z�v
(� Ũ�d����=f�2�y#���|�٨.��v����
bv{Br}
^�����g"��9	�� ��@�4WV�׌u�5��s�FrzSt�&��;s������e@����q��.�zu�P���C�%Z�J):���Z�+��i�v󚢩�C*76�T�N�2�]Eê��6z&��y9�k�xZ�^���@��ŨtBd��b%9�?���K�V/�鵬?N6鞔�w�����M �=�����[�MT5Vl��N���L� g�1=tv��Vs�ԓ��s�tw��,�C�k�����;rl��\v��y�X䒼Y���A=��59������oPP���OjfwY�7�`���M��z�/9߫_��<+��a>�hT:q� �Ʊ�q>��_C1��˲۞{�j��s-��_ur����*�t�/Eq�\�����w @AƑB~�= �����3���ٯ}8�9���Eu;Z�)�@�6Ⱥ��9�s@�f�ٹ����B{b�o��H���Y�+��q��A��{.�m?B�oe0�,�熡j����(�C		�ݛq���IpmM��99z�0L�S�2"n��u`�m̝�S�ak����XO��֨W��м�c�����mT�З�9e��Mb�ƽ=#�hg�:��:�t�{*	���UjZ���/ zr�W�u����`��a�G����i���e�mgQaͅ)!rΙ�ݪ�F.�Ӡ
�iĦ�G����W�z��0�ptC	���&K�N���5�SEgo3g]�N�;E��K�q�nǢ^f�{c���^F���@���\��~�j&4q�[��ё|qT�0^�)��K��ȴhi�Hz	@A��i8"�s�<1̀̀���#݇����bT�L�E(>O��Ӓ滥�e�A�(5;d�P�����W���ٹ����z����Ʋ�t9�r5�<8)A��@�W���zt�lkWS(rV�g)8�kpp�[���ZSy�y'l
Ĩ��P�C�t�%6���8'X/����ヾ�(<� y��ؚ�Ƕ��֛�$<�c�Ε�!{��4�e�i���1�ZE*܉��ez��ǘs�&
�Z)zQ�ƭIk��)Ł���`���8�17r'�li��vκ���9ݼz�_w���:k��Eg���`�O����L>�j4;��s����Uj�k�}+C���B�m
��w�Ӛ�1������ڜI|����_W�f��&�Xd��ۓ�˙("u�g��R�&�%P��x��������Ǥ8��H>2��vִ� ���D�*�#L�N��d]`�c@�I�k�85M��j�@
Z�ŏ?�K��,-�|N��`y�_�g��5�]�s�r�L��'��Lk6F�F�4�f�ii.�2�R���7�}�3��Z3r��zBcCУc'qVT�?Qi���,kwDj�{���ţ���Y,�Ļ�t�?�Y��{�讚O�b��a9Br9�{g���;F���E��h�e+4;{��]hp`|��:��4ܮ��M����U��e'�8ڢ���<�t�"��ӫ�Y}�D����X$C:����j5w�u[�tQ<�W�S1�z�K�^��o_lI�+�j��),s^�rƳ��m�ll���6&/�R���A�Z=����c�j$ԤU�{|���'\&<и%Lb�:��U��"jě���{�߲xH8����Y��P����]@AC�0�yXh���OnF�d;*�l�K��I�����6�b��'�{Њ�V���KRܖe@ņv%�5p0⾅4���G�S�����+{B{u<�s�?^@v�����a�zHzZe LW��b�A݊3Mz6Bki���O�ûo�_@��,/��z_���5��ƃ�ͬa��<X�=��2�[(tM.�ѯ����1/dS��3�: f�J�u��v���Ǯ�Ӫ��T���ss�I�rm6ŝ3�4~y}P/W�����k��:1[�V�ߓ�,�ٳ=�>�Op�7h�q�fڸ�V�X7aw<F-d���фEm�_we�R!eH%f��T^M�9�V�W1LZ�c��֒pކ���b�b��7dk�W(G�R�q���}��V�0I���{����A�b �dp���|�|L�xH߹��{
�^(�=��pɻ_���>#Z�2�G�^OZ����6a�k���AKK����F� �j�S�2��r����f�J�5�����;.��봇� �<\�!�ٴ���`e{JnPΠ61�YK���h�c�,�s_s�n �eZi3�M�ZV�y;��ݢ��f�@��Os��!����o>�
�e4i����W�Y����z�uj�{���j���2ُ���B�˲؎�&��3-�68p��s��;�y�4�r�2� ��<����F�z��iT֮g�j"�g1Xk�o�ʫ'�h�1IwO�c�v��oG�wi�K��ݎ�����~����$E��ʋS�Җ׭G��*J�H�L6�2�0Md��3x�%J�iH�oK�i��1�\�%5e˺����;ck3"� $�>R�#`4O�`�r7��G���Y"��͔z���-�I�wWM98xn�>�gv桤W����q�uf��{��/�'Ź͑�Q|��N�L~�q�S��x�A�F}�Ndd2�h��<$��$��U�a�у;2rCz�D�����y�ԻXb�9oc��W�B�y���j��u�s�PO���`Ժ���Q��{/��g'�>�RdVjl���SD��Mዼ����%X&�m��ތ�t�Au��F-Μ�iᣫg|w�����Kr�J]��X�r����,,J�L۹k-p��k�R{�C�M��}۩I-�����w��ڻ��2���*��%����Sj�H�h\oK�ܟ��CilF����Q6UFE��P��&��c�O��z�q�r������~"�4{�d{+�� v�5�G:
�R�x��":fތX�r뻳U/r��4�E[<��-�+G�[:�$��WT����n��m�i�wk��x�x>Ҟ�u#ݙ�����#��+]����yj��؏T�ጼ>.�E_<�S�.�<*\ﵱ�C���mUu�m�v�e4���qa�����j0�f�\o��ػ<�G��6��
��xt��볡�kz��M9ПP�l�<hA����UVW<Ҥb��{J�	�ѧ>�RƫO��7X�z_'�?
�^ �#��95F��U��P��b�n�NFkoPk��ww[�^ftމ;L�yHa�
����q�N��Z�</��g6��۸e�Yn��,���v'cI�L��刴�8ՔI����(��v那��t����#��uv^lWҔn^k����V��8��q�b���<�od&���>����^gR�R���C���Z�@��G����6��;an�zb)����жV^7�ѝ(�*-ϟ=P�'Ã�WK�`�F���^vi�J	�>\���j��A�y_]^�f�dV�*�h{���8�L�x��c7Z����X�AgW]V�D�
09ـ��`�2��וوj�u��D����ڮ�e�0E�.˗�G�+�j�ǽ���nK����v�Ƒ�����C��GN��ޭ��o2n�Q��y
���q�����t��!��4z�μR�9��q��*�!>[��uҴl�l�����݃`:$2�LŬ�Ic!�e�x�m'"�ǛRa���X�`��8v���B4��9�I���2Ӯs��Hc:�n��Q*�Y��d�vƍ�y٘�X��ȷS1	�C�jZ���i�7�6`���.�������G:�o����R�On��oU�y�n$#��d-����*��՗Ԡ_:��]�<.�1��ܹ�M⁭��Ϟ-�Z�Ո*1t������I����o���]��y���OQ�J^��Lm؏ˆJ���`�{y�I�w/c��hS�֘��JQgxθ16�7�.>y��)u��@���=����u}(�24[��ޒ�Lf�4�1K����T{K�v���Ú@d^�E�8陼4V�IҔ�s���F6�eվC{Q�/@�1U���ʻ�]��=/[zM��=����|��G�^Tz�̋�	��nu��V���{�z���^Ԩ8r{��=\(�'{���V�0�.�;/���U�R�^��}�,��Cٲc�ѕ`��a�t�J�t�l��Rv�zuoN�7V!ůL��1@7��Μ��9=�Qұw�7Vȉ\ⴡ���_7w��;:��9K�A���\7��ѧ��kNs��ɬՙ̫Ԙ��:��a��U���d"P')�����@��%t��\Olg$��nK�y�{v㢮��k��9��4�E�*Rȼɮ�gw�)���v��56M}L�X��E@�
���onEŽ\�h��aނ	���t��S����	�1�c[���z��d�Z�����c�1�MEb��7�.��s�;ǩ"[L�b��ҋ�a�X��3����Ts��s�j�	��6�NC.�-��.��<��)�Q��g7L��̕���.Uw\Q����z��ﯷ+^	�E���i`���l�SB�:ƅ�|��l�J��e�8��s2���e�]�n됺��\��䜍r|�)��CW�)�)A���剀������/{��J�μ
��+N�,�}K���eX+T"X+/b�;�xmm��p���]��\��E���.���GږS%l�j:Җ�a��eJ�w�5Iܦ�?�����}����߷��.녲1fѹnQ&���&K��()-�4%��
J"��5�n\��4wtW+��U!�	4���4��F�n$	��,PZ1
l�3LQ˖�*�lS1��%ݺ���".[�+@�$���s\�I��� ����uŲ�ú�J6K�IX��#�Bb�r�"Jwk��rђ�ܹq(�G5�F)�[��E�]6-��a�s��(�h�5�w9\ۛ�p9�	<��\��0h��\�<wN]���r'Ǽ#K����%�v�Є�M�
]��r�p1�Xz��ӽ#i��ǳ�h���>���򜱈�ܵӨa�zS��$(���I����56�c���t7��"��3פ�"�-�� �b��׉�ގA�����s�#�Y�l1�`�x���mq�BQ��[g�s�{
�^�m�7ʇ#�g��E��}��:]�ˆ�O=�6v��i!�J}�+��u���!$��� �=泝�3�+1��x͎6��7�'���Q������D`dl�l��ɷ��j��]]F�ݍ�Ӫ;cn}�dۙY�cX)���M�P�����:��z.��6�9/F����c~��i��}�����?���s��O��6�0i�ɨ����`7�}�+���5�iJ�������ә�[ md���|�<U`T��]�`;}ڸ!��!*��ĥAIUO�r7-�[\��40ə��A��v�>�"�p��S�RW������I0������t���s��v2ͯ	�i���d9���g-���]L�t*ẏFȋ�B���iT9战o%X�y�ulˬ�a����Z�^�5G��f̛W-mJ��i��	���љ�m�#��n��.��ňS:���c"�:�;p�9)5�͕��u��L[[�:5�O�I��!Ԕ�]$��*E_<�f��3��X�}�U�3��ݸ,���������5��Ք�4V�:�ݚ������Ή]�Eܙ0�{yt��}�Y߽����)�Iф�u�F�ў��WUgfzd�oc�=�kv@6�M0n0t7���8[2�\�>�PUx���݆0���H��(����jFHI�Go�?�<Śrd4=H�<�����懳ف�>1�q�<�������v�2�qj��[�����K.�"_�`��X^��vo��=�1�#�u��:,�f��+sѻ9aVN�tgU��H�g1G����b]���זcI#x�	u��[����N_i��8E ��)�@�g�,ÛJ��(�v���[���u������n�����Iv��Z��a��B	[��x���z3z�CL����8U���o�6iuO�6j9@��-f�S-�;�l�O@P4��@�Zd���a�����y��V2�˿/u^��M	��@�Y��|��H��3Ys]ʗ2���������[Y̤��������])�"'5D�%�ڼ��[�� ѕ�;�:�+��=�8�&���{��#�9��%���7�����/�&n�1.�iy�cM��jH����(rA+0t��=W�4�E[*rՔn�yS�v��TdB>�[x:<������r�y%*�q��}�]�����x���j�����){@V��ۅ.a�U|�|L��F���&�t(�&V=Ck���fĐ旺�e������xC_x,�HSF�I*�yg��;۝TG]��ɉ9��zG<����z̶cﮂ\ �-��P�M>����Lt���<��I~����y\��t���d�����ϖӑ�t��H��^�]j���u[ݯ<DmNо9U|y���c��`�����;�ON��N�%o�3�t5L�N��Th97T�����b
^
�d�0�t��S���Y���Fv�����������J��������[~5��L�6�n��w�BK�|��X���J�C��%�so��c]� \����fwp��򸱅R�ٻ�*���P��W�v�f�-v�E��v}�nkc�ݼٽO�ケG�a��y�'�3&n�����t�1Vy,]g_�����9�k`:f) û�ݯ��y�7�!�7���;��k-�/�e�1�S���&�v�l3�E߲�ãMG�����=��h2�n:�����Q��^�p��3�[�5G+���-=W{�|rpH%�O��@:(�E9��tG�_3���)���Y�#v��*=�=�9E��'�TF{O5,���3����͡y�C57U� �I:o�����������|U�)v4�Z�j�s�>XSn�M�]e`헾�d��u��<R/oKHW�Ñ�$���#:���#WVI-''���C0��.m�}I����DGq��΂��rFa��vu�\����Ӑ�uƜ�U^;y=4�4΁��[�6������l�n�i�u�j7���z�Y�^3%z�F�HܷSِ��<���>�x������&߳����M����y2W��e�f8@����<�ōdl�]��F�m������P��%ۙ�jhA�B���V
LL�v^Ŷ4W]��m٢�+�~5��C����q�>����V�Mߪ������ّé�[�]bT;֡8���G��[Aqq�Ym�p��^i�C:���p)�D��s�T1��O՝�f�߉�,��2��\q�!��{�˨�ꡝQ���{=Y�;�0�Te���dY���U��ԩ	w�X"��(�<��z�Va���#������#q��gP{%Q�3�g��yr�]�4�h���ϖ�.��m�n��Ul�`��`F�0�`WH��U�i2T�7T���57OVt윬ݯvђz��]dl�7F���go0�^{ee��d4s6M���n��Wr�]7Z��oF�z:4�c28�0#���eM�D(�X��WvT]>7b��+{�{��>����&#݂�|4ۙ����z���ζ���s�s`�"���^��&��tz��i$hI!>G����)���~|Y1ó�1��?�t@B�=$�7=�ٻ�:ΣDt��wf�̑O�UǅNY=�ɗ�_H1Oa����	G��M"�.B�WG�ڭm�0��_��݃)�x�:�w����e%u�B�&(�� ��k<�F˲�=W0�o��xCs ������9��Zme5F:�F�JWM��$��4^]pl*0�9����b6�rL+Q�ZŤcU�Jvh)L�ۈ�9�fTdnGgU;��z[bo�{�-9�8�i���ӝ��!N(#��V�M.���E���e�eXr{���.�)*��*��ώ�Ϫi����7^Y+//����Pc����UV��l���tV��r�P��@%e>U��eL��YUP��Es���0��U���U�2�,��)��*�k�SL��b����n��pE6�ܝ��QE4�%_*EsA��[T�o����Nm�َ���f7���&��
tp�����:�Ք�V���I�{&�5�KvA����]�qi)./ڌ�y�}����@~{��6��M,d��mn��Fv�ݘ�;$`�c�{͓��<n����}����p���2��A���f\O|�;ݳ<c'$9�u����z��?����O�7�GeƼ4�ʔa��l��N�������Qb�[���9D�_�������Vq�Pp�o��nc�d��w��%�b�6����RMIۍ�CY	����������%l���9�%���d�2��, @%��`�C��t-wM�/����ov�QBs�m۽��N�vk{
�s�>s*�}5J�r�y�����:��I]�
�S�5R2%Kt��4re#{�/�_�d������=&��d�	3���"̄Ҳ�֖c���]܆�.����	���n%Y����1����=[�]�ۡ��[qK��w4���)�r������?$��״{H�����㮛*n�������quy,�ȗ��~ا3�{N��C��j�G�wb^h�9��YK�c97�ht���A#�9���L��f��n����A����uYx�+�7���旷�y��!\w���&��1^��f��Q���EA�\��@�#�[�.VκW)F�JS������ɚ����m�ӝ�����O�[8�Ɉ�B�p��d6�y��,�F3�;5��Cvw�����M�c��H� �d�>pR+G+�۞��'�����߲oI�?@絃C���-��4[���[>������\����??��IK5�-ד-d:��+܏7�W��~�����}�^�͕�f�W7������n�2yf�$�TJ�(�����i/����ed�6��/\�u9�6������K����
hfV��uK�-��e؍��:�ɻz��j�i)9��6>��<�l���J�A�G��d�����t��9O
&��9�-(�Z�c���f�k��PK�v>`�ms�A��E��r�3����[����>Ɯʍ97U�)���g�H�QS��5�z�=�׳�����9!ɁD�vM�NJ�e�+�uU��e��&�츼eg_f/-8$�n�w�o� ���F���g�Q���=$�q�����y�ظ�Z	GO�Ϩ�9��l
C:���*u�eu�k���U�8�Gxo7mlѢFk$�A�F}��C: `�^��sèqé��Eh�N�)�y~�]��󎲽�Y���ll[��z��.2%�(�0Ǜ9-C��x������ h�U�p�Uҳ{�TF<���ō������h�C~`=T�z&�tc��l� Rs��TU�ӯ>9�j�����K�X�S�_�2.N�kf7C�s�i�DE��KY��yz�Na��#��|�m>'��9���d�-��{:ve�YJWL��@�[����*N�]�#��Z�e�4�M�0=Ɏ�r��p�.M��j.:lpn9���G�W}j{�0�������	��E�v�r�Z2E�"���G�������(��}/g�#��:�\�H@�b����3T�9q1-3��v��v���'��K�q��X7-��d���v�)�Ic�.�?ev����C���� gA&��*��ϊ��j�G�I�0#�=t���E�fI��%�3�/�dF�3}>T�Jh�.)=
�K�Δ�6�;<vb5�4=p�[�Z����I��0�E�=��͚��|�W��y��]�z.�L�3G��E�Ύ�Ht0~��`�09�z�l�^3Fl�Uo.W�5��� P칺AA���qPg��"�/�a��toC0+�Fv��4����v	W���Ί�M�H}^�kjzM��W@[#g��7�4s8#y�͈�dO44���Yέ����;����_r��4tާ��g{���6�8�w�X��u�;�I���?}f���`_b��G����)o�zt>ǕmA�s�/kH�'md�f���61,;uٮ^_�{��}���U��P{�4c%Ty�i�ىKT�Rf" ˀwOw��.5��۫6P�:����^U�e�$���P[ʣ��ضs���:�ߨd��V�~����W"�����+��m�ntAk�ȽS������:~���|�'������t^Y���H��C�7	w�vm�I��DDj��ov�����13�� �0��{gRo+��Xjw�=��3n�~&79w�x��Ξ���觏{a�P� �=�Ix���oP��a/uwUق�^V�o+$���vd%�ה��s#e�����Nu,�4�+U�Y�[���H��`�x�+���(��OY٫�M?H�e����Q0H��7\p5L�m&��D{o�q��>�w��2�*�i��݋�i�Q����6��X�F."���&�֘��x�#^�= q�L5^��KR�|Yp�B��ܸ-���pEC�[S��Y
�k�J�T��,��J�x��[gr���s�n��;|m�� �n$F>��g\���=�c����������=��/����}>���A�����8W�M�Q�ݒ��.�MѡX6�:y��6
�Y(1Մ��L�/)��w���*Sx)��Ѵ�ָbW��v��)h��s�h�����6��!b��Ծ���ݫ͹��`�,�p�,��[��gA���u\�)(Wel������݄;9+�W��Wq����V- ��Д��1��vi���u��i�ڈ�Ȕ2�1�J�+�]�L��ƪ��Z���-���ʠ�uN���gm�;���I]AEB�9��V�� �\p�{�mnYQ�����z�\�U�aFaCts��d�l1t��ڋ���έ{3��q>���W�+�}��AD�x�9n�s���s��R�Fe3��8)\ڼ1�Ɯɽ�+������6��;i���Qw�yZK�d�k�oB��$VY��q��:RVl�]���W
��U�����<���Pu��������}���n쉝L1O���
Rɳ��MVK��N�=�M]��H\�\�crn6�Cm��u�N
��|��@w4��ǽ�۷��pM�u�9t��˙�qVG��}��VGP��N,u+�q��g"`V/���;�"�Ļfpg,֔����NvI�땡��cXK*ݺމ��S�ƕhMޙ���靸�Y������T���������3Ton�e�ݠ�ˀ��sD��j
5q>ݺ�w&�ȟu�k��h쏝��%��k4`VX�Hb�(.K��:E�d��RIW�P�u��'-D�d�u�{�c��	�)�B�/m��+&��>Έ�� �	�s��$Z{�h�Jb��f�T�����V9E4q�˷�S��ǚ�����;Sܬ�ob�ueA��Xyst�u-&��Lk�Dο�*��ӮXQ؂�e٬Rh�kz�\o� g5�x�u���i��'�s_kbVC&ڌ���Ǟ����:��0���q`<Wg(��札�C�H�V����M�5�@YΨ(L��ճN�7��� �x��pe����ٌ���M�k�S~/&��h�9��O�E��J�}�(Ȩ2f`�X�u��2�����[<����S>u�D��
�D��:�X2s��CU�"��;Z�^��3(�5/G5�s�r=}�̏�l-�}S��(��,Ci��[�u�}S�tw��ژ�Go��5�k�}8�-]��3zet���I�ed�u,P��ϸv��W�c�G���k���3Ɔ���)��H9�﷝N�vU��;�y{�H�.�e�c��M��O��K:�A��Jkg��c��˓-;z�{P$\��И���9WZ�a�RZ�I��	���R�Qz��.�u^��f�IVV��.2`��o=�)��)l��v�!�]0b����m�&��je�(�5�y��5��ٚ˹ɨ-��ՖceRx��3��pc�V����"�u�QX���6�Ɩ�Y@w绽�����=�C_�~��j-�r,-t�H���wv��0�륍r�&K5��y���os�rݖ�כȱlX�˄U��E�6� ���.V�\��Ķ�$���hI7+�\��˹[���A�H,-�72h�cr�Wwk�w6�78S��Xs�����v��6���\�����ֺm˚�Ѯ�\�r��(��sN�p�s��\Ӻ
�ndK�r9F����)7'v�*��˷9r�,r���k�cs`����7]�ܮF��W+�ٷ^�^M�ۮ�������G��ϊd �	,߭c	U���W�2�AZ�glhnF)o�bj>{H=`L/,>p�]S��h��M(n�uf��7V���z=EYQ5�h��8�"2�����n)Ϫ�Ҫ�I%��^�w�Dϗ�F^������~�
����9=_F�b��u"�WmPI�K9�wg��I�7���O�<�Ӓj�C�����;B:zEGu�)gME	N�9I�|7σ�>*Z�a�UnD�`^Ã�}ۛ�+|��݄��9D�����cd��n�VF�c�o4��h�C��3��Y"����=LzM{�W�"s:�\8Kj+X[j�]��u�������:����ث��kM����r&��Ďx5�� �6G���R�lTG>W��t/����O_��V��9����)�Oz��?MK!��*�N�9��<��:�b����覆c���c��9W��'��6�$u��R.�F�d>���z����1��;��(^C���
����U�	��$��㶎՟W�z�<Hv�u����}�iY���3pJ�=�T�X�e/-(�֞��
{/T�b�(�muU��ˮ2Ӿ�[\��S���H��nh�ST���|;U�3̈́iȟc��Yɼod��a�f˥�Ie�&�19k�ܴid�6W`w�EW���.*��pс��)�o�읂z�����W0�@�M���^�(�IJ�Z�z"��;�4q����7�Z���[82���r*}��4_#-�c8���W\竫u�v{7w�\GR�IT�]sޅ�. l�l�
��.�(|���&U�vŜ��b8���s�Zݜuq�:1�h��A�9	���6G6%�׏Y{�'D��m>�5Ţ�%ʗ �mk?�}�HԖ�먯�<|`1ݵ�g���#���FO�����k���)���˱�o٘��{�:꛳v�Ev;(��1B�B*uW��QbnkJSKw��%?V�i��7�e��vK�^g�މ�`�x��B����;�oM*J�e�"s����`�;�v̾v�+Fxώ�ސ�}��0.�$��]g������>�ٞ]4����KĞ�ގ!��)�����g�1��}��	�:��w�Yk�cU�LW������f#]��ŧ�/=�[gA��5רP��9ws��үi�4=\xɚ��/���G�r�-�ͺ��Om16%��F|�oHk�V���k�s#o�@V��҆���*bà��T01l�,��1Byt����r�5�^IKpof�vv(�C9���i�����O4x��:���q���oF4��]�l�<��hi/[&��.��"}��$F�k喨t[��Tf]��3]�����oGs�`dG���<M͋ŧR���'�pT���i��}��F_4�lm��ԅ,��*<�S�g�2.W%�a��kXQ�c�m��b&�q�x����9F��֓��p��� ��G�Z4#39m���T��6��fK+7}�+���I�&�3����KĶ�Р��BA&�3)��L���.�;��A�ײ�.�V�E$_zH{�+�nDH��=\K�5u�F��syQ��3�8EI���r|�� gB'�"��4Wm��5S�٥�o}�]��5c#��c2(Ly���7�_(TSFR���FF.i����&��l5����a�mۂÜ0�!v/T����S�/��+��R/����+��6�$d뾷�����O��o���ˋO}r�]hY�"d`C�5<�A��w��n�z*�dS�pt��!�J�����������bu$��s�ϵw��c�m��gfI�[e*�јX�*�Wm��N�c����tń� =7�`�/��|'{��ώ�I�W�!��侭��l�FhϬ�W'����9wݙ&��v��5b���
�zXW�c���o�
���X�c�����F{_8��'M���WB�=M����ho릓�0��̼�t��|cu���T\�F�a�^6�fk]j��7Gb\�`�"E�
��*o"�q��H�ź���`�R*��M�s�dF��-q|l�P��P�6@B�</����I�A���ji��$MZӝ�}�T{�_m1�0����y}��xH��}p�8��g����fo�^Nu��7�4��Ԏ�x��=�$��?+\�KW��o�m�gW>��{���ț��
Uِ�cK^Z��8�!R("�˅so�,w;NOU��m��J]�Ќ��+�)*��R��;W>��3궟O��?<�u�1u�
���o��z,A���u��_��{�!C<A}+&���j���&��t#0b�>�Y��L��f���9�1��)ø�ZgM��©���QW87YӏC+8QO���%��_]-3�*rO �]J�]�^ɯ&��N�Vg*&�x��h�.h�Eu�R�XG�D���9�R5B��R�)*�ϕmj�ض��<ˋ�ݷde���j"q�@W�W���R/�+��2�,��*�t��p�ۮ#���u�s:���ݖ�Y
ѝ$��ⷙ��u������m��?G��_���p��O�5vuA��dk�ۺ���\�\�sOc��:��eq~F�u�%���[ ?ڑU�Y�-v[���-󬰮�<GM������/"�sωݓk�Ƙn4���0�nF�b�7�e�Mv�L0�:�9�?���)m���f`^J}���>�>��6��0�v���	aڮ5�'s���[>n�u��(���חJeF�]��3�oE�j8��,�c϶f1�M�s�aH�#+k�Dl�7GV�՘ͦ�w4�s��_O��k4;�#o
��f��}1n5k��3����l���s�ܷ���r��]�=G.ILї+�&���K[����Ǣ
o�B������[�L����\�fW�V�u���h�ʸ�9E�BF���������P�����+9��n�T�$�կZ�s�rn�(�f�r{?W�JLcǵ�݂��S��3�t+��s\{s�����4���}sdp��ϐ��x�%d �x�])�rYŎ����j��*��j�+�A�z�CN���_ױ��䄎�:GF�G[6�]2�Gji�Q�nn��/��`+Z5�%7˄dn�
�rB��,:GĦ� .��*�wwlȽ}B���
mN���H�w��g��C��\�1�u4^[���%�p�\c�A���H�hS�S��^���e�猻�y���bMm͝ΜV�}'�ʕ QUO�t�M�"�:B |ඃ�������im�;������̦
[�u�Z;8��=df=�/��/V�������ʯ�f�F͘����(\�r�7�ߝ�Q��K�b�&����ެ���ڵ�b�z���Ѳz�uO_-��rןQ�$e.Ŷ���z�s����S]
֧!��f]}��x����h�x�Tً�evF�/V�;��Nu��Q!���֫�Y�p	�o�G�Co<��W*��x�R�
�qs���xG�!��ʫ���Ax�*M�-}�rs]�+�C��YA��)�ɤ���+0�W�{�ե��h�p��!T�p*��q�:�G5�&괥4�z*r�o��;l�&���NR�܊I��?Ƒ�ցk�)<�[�������+\�՘��:��F�����퓤��=����Pn��m���~�w��lFs�(g!���lŲ	�~�4�eP�ݓ���z�ّ���}�0}��f�bR;Wү�w�Y]���"D�}W���tY���0o6�'��FGS{�4��*��Y6�G�8>_Az����jɰ3\��4�	Y{^9e�O|�10�-GO>�gF�<��dPl>�"��^&��ò� h�*Ȟ�|k��5m�LOZ�s����5��V�GK=�������=^����,q7[[5�֘���}�������z�=�zlTK�Yub/�a�B�[��x�>�1|���
��{�H/�,�%͙4gUP;y#��&��=A}~u�(3�I�T��~����U%��'�'��ܝ�[�>��V�j>n���VS��.���ۮ=�й|ޗn4�<&=�'��wkðR��u�F��M����R�Q1�+p�	P��b����gZ��{N��e1e+h�7��
K�\��q���n�c�3�6�s��Y��RRc�5���uٕ�p�̮Q�3�����??`mk����
�W�t"o��|�d�}h�?���f����y�f�l��?~��
�C#����ä�*���(�Z�q:��z��Iz���hZ[����|f?U] �\�H~�:|����*���i��$3�cyR�u9m�f)n�Y�ώ�P���l��`�<���6�EY�3��Mg&����9��=\��4|	<�]�!n���`�q�������eu6۶�b��1�Ov�(g��ϵj���J�tyl����n��p�۔y�	��/w�+�A{a�_.Ef�C
F�tM��E��l� V�7ws�yx�+��e�Bq,�P6���M�d
�Ƈ�C�U���<ّ��;u���k��8���Ψ،�f�����#I!��|}�7���׌���W�4�nW1�p�zz��� &�^oi��Q�<���սkVI��0�`�ϕv��g�֖y����JĽ�}O��1�}����S,(S54�
}.����d�����w��>u��v:���w=Э��	ˇ;ԵݳSe6�jw<$�����sן�Ty~�|΁��a�)�u�k�3Hr��sb������bc��w6}�ȝ<�}yj}�O�t��rnM۽&��;;M������u�]`�
Uٟ%�ה�\ӝ��*��GFM�;K{��v���(H9�����#D��g�V��K�x�H<��TM����+n٨��"��1���Wa/�O:
F�]Ĥ|���ֳ��Iw�v4��ц��v��m�+o#0t�
�D
�%ƙIX/̲�CBY��h�I'�z���h=��H������!Eϛ6����$>��yA�'t������_�q��Ŷ<BCpO��]��nH�ˋSZzk�r�w�#�y�y�{�ey�`3Ѝ�x�w��43����bOg�\w������0��.}�����k����ߘsU��~�ӊ����7��ښG���o$8^�)�Vꆰ�,�u��nt���4)�صB����r� z����:�-�S^$�^R��^�Ê�P�/A�®e1������og`ٹA��ɋoON�~�j�W�Mz�4�l:�X��'���p�u��:�l�~�O�f�jZQ3%G���v�-x�ƽ�~��O+��L1�m�s�Pr�[��oyE3R7����f��9y�۷�Hm���{G3��>٘�Y1z���ș��t2�Ә�gި[���U��}Ϩ�4:ٛ�5����
��K{3f�LOuV�Ln��7�Q(�$qc ���G^_�d3��κ.;:)6K�W��{؞�@���x�К޳<�,BB%⮔��s#%�BO@�P�l`�Nǚl6�,k���,����	�C�6�$u�i^+͸��O�j��8�>��膰����I�K�#gx���*�/(��Hk���j�nu�k;�v��y>�z�[07"�vO����T��n�.n|�gZ��"%�7zp���W��ώ�ϵ[��hBr*a�T/G{�{�ޏW�������{=��g������}��k��a�<��S�v��z�=ܠ���C.ux�ʉ����4_^,��_cv�����}+";r�#��ohL��t���&�GE�5��8r�Z�h􅖔�����W��ci�AFQw�����35�ȯ�>��w�WU��n��'��DDr��!��yB�
<����LD;��A��geEPN�d�I�7�o���ݏQ5VUN9����9�w-�(-�P|���S�=8��kz��f�짙q�X�EAŐo�1DQ��Lb`j�h��l�¦YG0h�h��j��[��7
�3k�9Y�5�[�WD�]q=�EHU #Vs�;؀���3s�d�#�Pl}֠��l����A�ަ.�90ԗڌ
�n�č�P�Q7D8j�b��;���YV��os���P'^��ܚ\ld�[X/
W�K��:�{��w"�Z,C8�:E�j�ά��O�s!dRW1ktB�@��
�׽ج+Ug�:�.}��N�K��p���B;H]�t���Xl���yr4Xr���[�(�gxtK�t��+�u�*�r�/����L\�oh�q���q�Xm6�m�7%u�c`��}|9qU�-|8[g���5�L�E�������N����=��,���w	j�R��
�U&^Е���뇮�8��n����]�uy*n���ר�ֺ���m���8,��;���!V+.�	�2�S���V�OV��ʹ�l�Jr��Se.�Hm�psʱ8�[+Y���Nؼl�Û :GL���S��z�ѥg�kI�l�5���-�w�kq�ܲ��:7jֱ�8L�a8�B�7ϏsEh.��S}	�{���^re2T�/fupr�T��z�̅\��F�P`��oWm:�<��.S�g�W�,P�s�w7JS�#��z�?<�+����!��}ÄW�6�f4�gV+7��e�U+cm䦦2�5��ҘtV�]{c�q�B�%o]����S�sw.�jR�Ȉ�c�f݅9�I�h � �����Y�Zž����a�m�$n�[U5�ѥ ��r�^��#�+P��޽��v^bh���o���r�Z�8c��n'e�8�t���U�=�YO��9n��Q�7�K="x�V0+j���x�2��J�� �g���d�)��c�����eь�Ű���w�qj�{����1� ��9��$V�d�`�k�@��Ƴb��d�����޹f�Z��3-aO0�h�l�J!�Ngnq�.-dXԥ
����V�귎�e�k��H-�Ҡ���3��)/�J����Ŋ��������/��4�r,�jn���L|f��A{}�]�O�����o1���X뮲��P9��a��5r�����ƞZ�sLW�=e�{ ��Es���G۫�tjb��:�0��n�{���1T왈��nqYJ�Cn�P l���Ι���1� �*�"��"��m}�=�5sr�snk����wh��깹��s�����W;����4\��v���g��[�9]�(Ҙ�](ܺ�9�T�(��rMwtB��e"�Y"��]Pp\�8�u�wuD�N���(c�б���q���鹍��s^^£Šw]0Fˮ�n��I���ݷ(���u��yn�;�e�p15�ј�r�n��69y�4�r�
�y\���vܻ(B���{�jK��w�w����N�\f��+�����w�����^is��<���DW���x��z�Q���B'��s��"׻Ǻ'.��m�o�s���&����:D���^{�{�҃�͹����1��`�HO�RD�@�߻3�o{�iIn��V��_L�8�lǙ|1ҥ���6F�Ek��օ����(2U4�@���j��zv��)#V�s.M�=�Y�o�Ԩ���on�H���Eä+l��m�R�9k����C���e4{L�������+��Q��x�t�����ܔ٧"�H`S>��υ��z���(�9R�a�ŭl��Rg�OZ�uz�� �U�������˪?U	O��M��O@�S"�k�H�y.�3 �c�v�]��M��^�vJq���w6!�C��\dFΧ�'\���)kή��BkzI��f+�n*#Rڑ����y��a�(q��-��ziETׯ4L\�Å�Mt�r(Gp�����:�wzF����}h}؉tZ:�F�N�v3��Os�ɺ��t��>�`�h�-���Z�����Q�5�9gӴ#W����9�8N�G��<�xQ�1.�u:������q��{a�'X`���V�昼�"F��"0��y{+X�
'n�NC�*m��WSW��Sx�a��e�iIy>b�<���'���Oh�i��v��Z����:6�,��B>6k�����`[�uھtu�nk����l��l�������0�;��������a�[�"1i�,�h�aW|.���I��ǧ�Z�E\=�5WW�u��@�!|��m�E�{�͔fzg{���WGU:�t��4��y��ld[�f&�lCLU����]�]݃H6������Op����1 !��_��>�����Ľ�@NB��$dٓFuU��:0폿W���U��^0e.��n�4�6��M���o�Y$����j�{��N�eF��^ҍ�O���3Z���JE�u��F��_"��t"ls�U�y2
���k��y�it�{�d�0�A��ܸ!��� �1]q�t��ʲ�}FR���Ur�\�Nˁ��X͒I�~��\5����L��������Y���S��u����x�zH������{��u�	q1��,DF���TU3��D.��Y���rI<�Z�1@Jݕu���pWս�B�zy�}-��:���,�2���u?�����G6Z���8�&�4�5׻��SAK��r$*��Y�`m�f��o��'sn%�
E���r�����C��P�;���ȧ�ѩ��0������MS��[!n�A���ҜA����7���$��v�����e^�u���P��}���j�N�H�~>��
J�;��dl�7@����ݳ�=�վ�J�&^�����Vw*
F�t��.F�l��d�9���%p�ʳ�ŷ�w�����@��`�#U<e�F2Sx�Z��w�f��-�}C_/u�2�Nÿp��[7�;HEl��������\h� <*5x��u]ve�ɫ�L�C1a/1{Ŷ`�ṽ��I5�yEG���}m����zJDm]s襶��:�Yv�dvt�U����i����S�鸞�qb�J�Z�Nn��{����vsl���=Y�K�AHWfR�i��"��s#e�xRp]�ݿv:��l�"��Q�v#�18���%V��S�'j�7�O�/,�@��ܦ6�F�u���g��d�t�Wa���΂�P��KWl^����j�Ԛ	cc:�vm�t�Lbi�@W	�!Қ�D
�24�I��޵��+H�2��X+Y�� ��0'{��v��҂V0p��>�f��7'��%g��|r��Ǿ=�7���U֏$���:��e
��
Y�/�;q��_�fs熳�:#��z�_<�6R�"9ei�Vҭ�ff��
+m^gKSa�(�e�t%o�^[N�K���n������H�A��Z���8"��;�H��"c��D�C�g[L_\�soFZH�*�<���;o�1m���,R��*��'w����'��YX�z�e5zC�#MV
&B��!x:���;3��k5����%Ά��|�".s�%v��\Qy���N�k��~��gġ��9^�s�E��G�#����ҧ��F��ZQ3+e���X��<պ3x��m7��z$�'��2�q�������Z�h�4��z�f�X'�����L��z[v 2�^&��`6��h搂1���W�*�~ہv&��~D�<�@O�)3�b�h��|Lt��=!�q��bB�0#
�Q����W ����nO�;�{9�-_� i$H�����
:��q��x�V�h����/(�g��g�tgU]�Ǩ�|� �{�W�Ns��\�.��R��nخ�}�����cɆ�ڱ�v�N�V��si�F����)���`���Z��ӱ�[�������7�S�q[Z���������l��.[����9.�w��@K�W5&ُ;�G��Z��pzv�N��wp?n���ѳd�Wϰ��HU��XY��2W$$u��i��c8�ϲ�����Φ��ם�B��x�?�+������X˞��g���l�>+y���������n��/wדsNgޯATP����v�^��\e��6�s��Y���Kz3I0\� v�F�uV� ���S�S{!D�U��Z���p����x����R�QUO�t�F��k��P��VP���;��{��{��Oe~��h�)+�\u������-��%�s�N�yY�|Т�8�����ò�rl�rJ+�.W�[ֶd��!��s�\G[v��+Fi�ݴ�[����X�덕�#�z��ȮZ��+�.��z��V{�q��<oDk#�t�$m�Ǵf�`�q�:��NS�ǰL.5�st��_Vv��0��)T�6�?��͂7��FDH���������m��C�~]Yڠ�r��+���
��{�̚�Z���\���U)P���	$o!ɝ�R�!�"�5_)�mY������Q�ݹ#�\TS�E����z�	L�̾�n��k����օagpK�=�ɀ���jG\M���gjf���0�i��c���[J�-YC�uQ��loHn�w�|�.x����;��K�3��f>��VȲ����vO�s�1�m�HjWd������N��o�,O��}��J��tY���8o6�u���=RY��g��jř�s�GCQ�g����Ŷi�זDN��@J�C�E��/&��M�h��ށݮe+��s:;��B�D]�x���;!j@��%Ќq&ư�GfN�c2����W���*�X޷S��,��;wΕϻK�#B���1crV~�������vp��4
�i �SÚ�΂���)���d�/5`�Q5���k��pUƢZ|���|lɣ:��v�^��Xs�&�7x>��Rjx�݂���1�EiZ�u�J��%%��k��u���Hb�f%�"�Z�콚�|�,-bGw��R�B<+�gB�y�+�z�������V?x#y��e;m��|��.�#ƞg��n�6�.��."����R�I���|��C�a鷻�%p�4��՛����G�'�� ֋�_<�� w�
�N�O�:�]��1'����P��P��P�+qv��!u �����ަ���j4;nЬ���m����d�l6���2�Os��@��+�Ѥu�E1e&��;a�ˎ��m�y�ݸ�#�Ao<�'g��;	p�Y>~�9jz�z������w���XwrԒ/4�K��:С��e����ѓ�"��-V��nwl�6k,�V�Uk��Jݕu�,7���J�-c˳�ӳ=]��}��kU�J��d�Z���W�] :a�����ƠC�;���}�Pw�!�&����՝ʆ�]����ѵ�}s���jc���'3�mv���&��>W=�UmdV�4#�����\�Ʒ�S��Ӥx���5[��g@��f xT_+�m���ܜӜ�ss��v�ͽ��=�$iHO.hkC�_3��,�zI��Η��w��k���v��^��Ú��:M7����l5�����?�/��/�в��N��k��Z�����R��̵��T�U|�1�+��"O?����^I~���4_�Y4�u���|$�&3K1����Q�I�cɎ���5������-ġ��������T��lt��V�[��aޓ0��(�Ԧ�}��mOhn!����t��u!]��]�7��$0[�HsG��[f-m��
{9m.�L@�!e)+J��^{�[V�#�*yݝ���NP���i�����|0n��wa!�D���:
F�\FTլm�8���x"�k�w�����y�W4��Dc�V+�[���6dOU��"��^uu��<oP�&@��1�Q�ˈO�gT?��4#,�����>?g_h� &x�R�\�eco�1m�0�Ah�s7s�w�yk<�ma#4ĥ�0+�^��(�y�GQD���2�u��� �}[����Y������!���f��9mW����Y�N���춭ǖu��^^�ý�_��� `�27懷����y��֔��&��>f�fC��mV���x����\⏇R}���8�q�ϣ[r@��T�^�)�l͸n;�2��	��&�*^�L"p��e�u\��K�$�)N��9.�%㼥uy�h+[E�`O��yd��=��)�
���ת6��Wu+�'[��u#�m6�k1cE�u�υ�;�8��Y�L�Wv�Luj�2w1��z)Ƥ�0��ӹ�8`���>g�?~+}�!�Ϫe[�q�G3��>٘�Ys�/�5��_1J��?:�ܷ�]&��d�c��E����vt;�%�EHz��M��g�b�w�f���(�D�>���x���S���\'��	� �ʹ\�0y�3��GyG^Q��WDD�q�K�K�]*��b�]����z��\:B��`�"�j�hD��^�.HoZ<m�
��f�È\ggv�S-7��05��PW�,���ͪ��27x�cD�W^|�3WSV���E��qG�Ѳ;�x��sNf�@�nxZ�V�]�x��SwénN�i�b���A%*�S�>;W#U��V�
b&�=l������v6m�F����E�jF�<�*����}��S�p�[OEN۳?���c__�0־=�5�-ţL���q֎��WP=eg�����E�$����\��JϾ��?/�q!�q�L��HP}K�<�
��:�75��j�
+g�g�5�gu�����y�0
�;��Py�q�L�'L؊�S�V�r�U���Gx����U��N�f���v�wQz�j%��o���M���31Ծ�m����x�r;dF��Ц�4�$���\����ֆ�3<z����_�z����%�pZ�o_�euꞯ_)�寤SE�پ×s��6f�ꛎӨ��<Ӗ��`�q���]&����F&� Ω���ߡ��Hw������%*�����y�!��Ɓ�4dآ��ksb�{����grWS-YC�u��ϩ��W2}o᚜�ʐ��nw����D:�j9�o��z��R��䂣}�]OPb�ot�n�-��z���}�eY�s�|�{E#��f��Ϳ>�Ǭݝ��߶��o�08�֝_��¤����l3��,ߞ96ͣ��/,���'���\��ٕ�q�ׇ"��t�ٯe��R45��v���߅��=�'E�1Z�J��{�~�͐�������4ԝM���&F�����YZ|;�~�+�҈�  i�
"�����|h
"��O�*T��W�7��WY�������fV��fV̭�����[fm�+fkfV��̵���m���+fkfm�+fmf[fm�-�5�+e�ٖٕٚ�+fm�*�mfUL��V̭�[3j�[2�f�e�el�l��eT�ٕ�5�6ٕٚ�6ٛl�kf[fkfV̶��̪����̪�m_Yk���Y��5fV̭�[�Ve��YeY��5fj���ՙVe��Y�f3Ve��ٚ�5fU����3jߞ��[�koeUS-UL�kU]���m��m��U���U2֪fڪo�_�ݶ�L�Z�[mS5mS6�S+UL֭���vj�Lڪ�Z���M���Uvm�ٕUL��fmUL�m�-�ٕUL�m�6�l�WUU2�m���f[m�*��j�f�m���fm�ٛm�o�v���2���m�f���m�eUS6�l��̪�[7+�ٛl�lͶel�l�l�l�lͶ�o7��+fV̭�[2�elͶel�ٹ��f�el�ٕ�*�V��̭�m�������]~_��}m�Պ�[[2ڵZ�k�/�����[�ua;{~�,��=����gݺ���
��ڔ���r�V}���UE|���}G@W��
 
��|�� �G�>�_z��և�UU�s�9w*�MC?B~��7�k�־�����
���+����Z�[%Z�k[XխX��Vٶ�fm��֪���e���M��6��l�j�jj����lږ�l�6���j�����Y��e��l��U5*��[m�Z��V�W��

�ڇ0�(<�{jv'�TEE�[[E��UVk~���?�������<����9��UUTV��@��"�&�+q:Y,~EN |��s��L���UU�7��NZ�ޗ� WQUTW����ۡ*��CYP d��ޔ��!�C@��
i�X�lR,�UUU���oC��]ꪨ� ��)@/ϑ;��k�o�5O��x�ƀ �|�y�
���l����"�ےP�P.��1�Ӏm h�!	~��UQ\�8���s�Q�,]�*;����dW�ـ�nr�
�+H�{\n��9����
�2��'#Z�3�������9�>� ����	�B�B��I$�B��%�T�
��� �@�*%
TH*(�!)J�"�BUT
$�QE@�
J�U@�QR*�%(]h�R�*H)EUH"��*�	 ��I*�IE"(�
T%$JTUB"�6j�)EJ@$�!UU R���J��TQ
"R�AA�QD��*B
�
��UR�IUEU
�@JMd�	R�e.   N�)��1�>�.��&���kM�����m�v�Қ����h��lL��mf����+SJI-XKV���nkkS$�Z�5H��*���"���   Zá��Q"E�447�M�P�BFؑlh]��(P�=����й�áB���K�� �V���l��j�څ���l�RiT�uҴhh���ڕJSL3)��T��!B*�B!$��   1ݵ[SJ�Ym�K[E��L�mm��[Rg�t֕�ڪ�)Um��Ұݻji�X�J��V6%����i�Y�j�[[M����t46�@�T�T�U/    �N֊�5�e�VԫeX`5�7�C�[j�a�P\Q�w.��v���cm�DimUJ��j��R���j*�D�m�UJ��J��R����T"�   ��J���W���m��1#�gM(�VT�խ��b�[cF�fT����چ@-�J��T�F�F�(Q�D�)E"�K�  �➵EZKh��j�!�wv�wwjL�.�SV�
��U�4����Z��R��dP�F��H��QUU$R�R"'� X�%k*����4�5m��]3Je��Uƥ�TJdVֵ�KT�j��VC
�Q��@+��ΚR,8%D�P�TR�)D�� oJ 
�R�Р�I���ʸr��[�s�@w$��.3�t�@gQn�(*��(hts�pU*�QV� �
($�O  �� :�N�
:�p`� �3�`  ���A��e@i�]�cJt(:�uA]w`\;��P�[C� U�$�B *����7�  �{C@(Y�h֔4�i��aV�Ps�7k���� t nS �Ԭ�@:Ҙ �ΰ�ڀ^ T��eR� �a "�ф����  Oj�P�  "��	IT� ��F�M�2����4@��H�2�H  b5� ��Z�K�b Q|%%���%57@Ys�}Vr��=�F����r�����km���m���n��km�v��km�=[j��[Z�kk���/�����W����U­ۦ�J�I0]L.�\�Z�͓L��-d@!�t������z�f5N��*�Kۡ1�u���4>B+�ĕ��04s"�ٶt��������@t� �0����a.��*�ڕh�m0��7Y����lW#˺aH�Mni��Q�x����]�+R�Ùq�R�#.�#��֡tb��m ���_�^���Ѝ�]�l� ��� �[I���z���X3H !��St!�f�i�t+���"]:J�-�����l[W�W�F�i�Tk ���GkTt�5������c������s&B�uֽ��YP�f^�Y��G�c���T�D `!���EI�ܡV n��Un�5Y2�c��u`@U��Pe&�(���Y�bEZ�C	�	��;ohflU��a@�V�%�6F��ww* �Tq[]L�Q�,ׇ�Q�(���`=+W�5�1X�Z��4p�T2�p�Y�����J9h`��o&��	-��mj��hE#�"���v���C-�7rJ�zC٠B��3u�{�f�ZeY���OXO ̢�6��Y�r�T�բ��T2t��z�^�{t��Ɯ�1��VH�5���Օ���[j����v���̂�ͳ�4"�kBDҔ��ً�ceZ�C�lפJ���7��KL����
��'9`��ϳ�[4-�jݚ[h!+,�L!9�k�e��ȩjx�F�yqb�KKc���Z��VJ�b�k��ݩ���Ø%�H�f,u���n�q�� ne��t����krcQˎ�Q6nC��$���j�J�9RVS�h:�V5I�<�`��~sD�T"�Gm}�j}�p�Ҍ{�;���nä��71�(i�^b��8C����W��<���u2FE��
�U(	GKT��U�@j�FJyW�)[��ͱ�f��N�ݗB�[VH��:X �4~ϱ�N�n�`&���-�)11b��B�&)������3U�T��������a��]���1F�,n��6@Yr�TT�Ӛ`����\7q+Pܥ�$5n����]J���Cjʸ�AB9�s	�r$��f3���9Wv<�s�DZs�N4�f�j�Ř����Q�ѹ���R��k-�6��Ra�{VE"Sn]�چmX-��+׬b�A�!@6D�n����v&h�j.6^B�d� �ڽ�N�#"{j�:EX�B�Y%��Z�f@�#�B��wM"���]l�ǮT��jPF�FdK��eܚ�`ť���N�'J�C�&���e�&��{Sn�Gx�>��*M�x�F��u�ph�ޓLQwmV�ԍ=P���y��F��7d���[k/Bi�7�WE�7WW�Կ���6�s\�BB�=i�u��|��v�к�6&��ժjm]l���� U��L�r����e6�# k�bcv�k��`�(I��M d���e�*Z��㥕g&��f���B(lp�2�Y b���Uw1�8jJφ�i�xp����0��K�ZEa�IT�E���2l�0F/�q�1���[�����6��[c��6[�aM�Q9F��ܫ�z��CUIB�g>�U�Z�����,ޭ?��bV�X�ʸ~����A�%���ՉnIV�ncU]ɺ�&�k�kf�K�J�� -�	Y]��AS8L�2���P�9C�����e�G0�Y�D��Z�%��Ʀ%,�K4�V���B���i���R��e�n���t��1�k"=�u���e��z�Gp���
 �:��!��\R�֬����ݵ3"�v�Ѕ6�J������w1姠�Уc=4N��B��`����*M����՜�}�F�j��F-�n�n�Q9sR噶�EKf=���&�R%�] �.�����vU�Wz^�&`��(�e�
	��%��q��m���^0*�Z�z���ieH��n���JVG��D���u����kY��Y�j*Q�4hh���N�/v.c���f��*ݪ��LՂ�]���C�{��^e�\Ĩ���.��O7^
�m�q�6�unP�&�nG��5������G��Ò5,-�E	����bT��v�@�#�����6�&�:v��V��55[az�ɐn�YB���6ZSBeܧi5�N^�pA����A�Ek6�� Ϸ[��I�@iWvFXސnb
�̰�����uU.�i���nX?�T�&��Ev�m,y��b&�J�&\���ڷ�uxb���6]D�b��Lm�he�t�v��c�����B)hѻbͨ��`���ZȸrH��X�S)�bQ	I(���'w@h�X�Ů`p)n	v�amj��!J�Ao�S�cn����V`�ԅ8�A���ڛ��5�p+(l�Ln(Y�h����7%�D��p5f�L�E��?f�l2/K-��hۭ#V۽��捦�bV�/f��6ᩋSK� ^��&ۼ4
�Ͷ�؏���h�N�*nIR��Z�%���kp�8�K�і�h4�ܕ�F��6��a���v�J�J�l� ��cE4U)x��.�(O���,(���	!��c�W
)���ϊ�ǻ�3ݷ�ؤ�
��_X��C:7a*t��L��[���mT�WtDE0��f��i����1��H��t4��]�u1ix2���\%���f��V�e��Ië,fXJ��dX�ފ:EE��H�R^޴����EP�'��*��t����cHV��;6V3L����W��)�l�;BeMvGi��"P�4���ROwYO+dY9T�E�����!�x�������1b�M\'{��*� 0V n���Q��ұf&�/�c�b{	q��]�[�\D C����XvY��ձE��K҉V�0;B�E�s!4��];P]�D�ԫt�4�'�{���� ��J)K%��s3,�:�l(&%[b����c�q�{Y�#)-V��v%�yab����̏`�.:U)!x��W��+^�/+�f�$����b�"��wor����:H�ۭ"-�GF�$Ɲ�z���� 6'3B]5�"�&��Q��V쬁P�]Ѓl�tX��d{e�D�2BX��ָM27F�um�N���\��"�0�3MCYG˥��AD����H)�9��W�T�(�Z2�̦��#u�fa��B��{��b8�����iz�V������%�o\�;NP�'n�9�D���m���b�6��S��S��h�XЅio���qR26r��$JP�%��ol<Ms�*3]Ш��iں��se��!#�u2�(@���e�*�ʃY�*=[,�n����Y��Cg54q�"j�dV&����5�����a9��ҳ�R�*���<+�0o�##D �yN�&���z�c�v]���%ͦXs\�n`�� ����Ɠ�D6#��M�B��\X�(�R�mZ0"�tw-Yèhz��gCܙOBbL��K 7���+Z�KQ-�&�W[@4���
��ڸ"Ŋ�cr��l\B�J�2�� ��X�m��3ڛZm�3Rcˊ#�aA�PT�(G��WW�:8vA�3$�={�*��aU�V�X�Ӱ�3�nYSV�mT4�Ucor����s ��,���Yۦ��d�D�x,���g~�̌
t1���(ɬ��h����Gq�F[5)hR9�w��U�����hK���K!���0F���Tdhmf"w�# E�)Dpc[�{up��v�:,H��RՁ���:(䷚�Dy{>t&9�$�������
AVV^��u�d���B�1W�I�k.At�Yͪ�Ҥ��*T�X�֮�����O+	�d�6�MչN��F�j;I`��5�ҽ��[L���Ǧ�!+d�K#�X@ͨ)��P�Գ]��^<o6���4 �[(���Y����f5�X��a�ZP]���dJ��t� �)���`�������]�(,.� �d&ٚ^Xv��<��.`�f �'�6�j�U��5o�f�OM�Q�v\Z����j�iRy��ZA�TY�V���x�2Th���Y� ѫQ��É-�S�����F�f�v[R�+�C.�n������I��b��X
�j1�Mm8��/rT���;�B�љ��Mbj:[5] ���
�RclmaJ��{��Y-��Slͱi;����oLjDF�ñ�&�a�n�^�TH�X(�[t�	J�Bz��$��o�^1.��$mZ�9��(����QcC6\`�@Yم�d�n�ѣYia�oZT�v0�k�-����̴��VK��(e�T*P��R�]�Q�t�&�G�&�����e��.�3�F�ՠ.FR��^0�"�C.台�&���Z���S�MN:��k.�=2Ԭ�;��T�/.�a&R۬G]@��KQ,�[�3U8�K
��i@�)a�jb:��A�	@ûN�-a�wgX���vQ*x�C���s0����	Ie�4F���rk�,,�^�Y��U�:��+���0˖v�̒]o9ļ���H�Ȧ[�j�$PCN9�����	��iҧ�^CF�u^���Pb�u��7W��F@�����Xl�B�%3w"�V��T�5A�Źj��31�/)�G1%�Q	��T�d1`Z���=f^�8�5P��B���*�4�w"ٛ�ӊ]�˲`YwL�+5n�F:�2&~1�+"�@fo�MUڄXL�&`�R�J8T�"��e�r
����
F�.�d�d_�c��v�����t��d�wxF�ɔm(��[.�z֕�e�{N�ؑ��V�e=e�:2Mw��*���j���NGF�%p�yl��f��� 2�ر�E2�i�Y�YDܻ����#X��!mZb�K+(�偏[���tј�@i5E��,ϕd��ŹkZ�"�ҁ�c[������V7��j�i��k�[,���)6�E�N*�����Ӱn�YbB,r4�F���������h5���]�Ix�#y���dfe�,�R7�A��.�I�&������
ذ�bѴs]��:�=ϰ���<i�6�Eӡ[��9���,VAb+�w�ڢ&Z������H�t�Y�$v��2�]����ҝ��j3�4��sp����Os+aH�5٭[���N��ӴU��e�f���MJ&�)�����=�Ջ*Q��r�[(���*T�����̕x+**� hB�AՔ%�12EjZ�4�V�NN���F�5v�dJ�����G�	����%�u�*ŕ �v��kq�=��Xԯ,$@r�&L)S����X�J��D�����D���
����?�p�r�&J��m�t�4ɳum�P��F�����ֲ���W��\���M�[[�N��"m�(�4#jT�A�!��-����H��r񛦚c
�uw@U�V�t��K6>�E�%���pYWB
QV�`=�u���r
���*]�xY*e�f�n짺u���K-�On�7[!���L��$���Ի	��T�⠴�x��X�� Y��Ԡ�l�e��ZƖ`��n��n�+N�.�#S6���Ғf�y�#7.C����V��x��I�w*�Lj�j�3��S�jjFb��`�pE-`r��l�EM�˫y�t���v%Ly�{ble�,H�D��V�*,�j�W��XF�tX�5Y�r2�MV� '`޸�9�P=��+�(SW�^;��l��o\��(��;�Պ�nm�(���j��a����Oi�(U�$�X2�C�e��H�L�CwY�81U�^��v�#U<;M��wQ�CU�Z�f�Py��d)FK�����M^���)T��ں�����2;����h��6�6*��%�f�gm�B<�+j�dtB�6�su�Ŗ�15�4��,�ą9n*g�����i.���B-M��ɓ��nJ:�X���t�b����O�F��CR솬���JU������n��j�,�w(}�3\�Δ�)Su�V\���[�����q���m�2��`�&�=�ة"wt�jk4P]����"���1���2�dz�Xܘ4�QИ'��y����`�ە�݄pL�!�(Z�*)I���(b�csEMj�#�0��R�m�{��!i�	����x����C .
��0��Q�ő��u1HL8@��5nJZ�]��zF���֩��H؎^ ���E(�[H/lXX��E�K��n���#Tu�k
�7Sv��pDګ�l�rlb��.&�fE��ڎ����{����e����1�__c�g�q�Cf
�h(�
��BfT��vr�E�dbc�`+�tK+p�wpc:5k�l���6 Z�5�ͬ�i�4�!�*Rn蟮�])*;d��b�Υ�m*�x"��^�kn��V�wA�Qn�o�Cxr���r���mƶn�Xu
��4S ��)�R�/uѭw�Z��E*��h����b��*+cF�mC0��	J���:���������y(��n��P �RjG[�K�9PH�
���rjW���d��C���N��X�/6�]��86��I9"�0�����	M}C/*n|h߶e�7��pG�b}V<�N����IR�4���5�e�2�S*�ZvvE�Z�4E�,^�R�o,�j��{�M���`P��J��kvؑ��0C�������¥f��g��j�,ުqncB��5��МY�Ԑd��-H�gW2uU�(�� u���R�A�ѹ�n�n��)K@	��vJ�te`�0�E���;caI`�5��g.����d^����HR��,X�J��q�ͭ�p���0:�۩�0^'�t��ܥ@B��+7kf]-����P�<��v�7i�Q�!ػ..[�5�7�9��=�J�eolC��Vr�nK�N�]]u��k�v뇀[��|"4!�Z�l�u�ƽ/��3�k�A1�W��+Ue]b��MK�R�zj���Sܮ��r�]�r�w�Y��Ϩf2�3%F�������w'(��ԧ\WhO:�u-q1`���줍f�����|��-�X�.Y�+)�YV�k�ns@	��ھ��pX����wI�`�Di{Vܲb:s��M�5#I���؄F�.�q/��Y΄Q��6��R�]�jN��9�Yk1�_f�t1aQ+��MN��Zɸ��]vJdG���bmk�C�j�+�6��T���[$I�ѳ�뫯���A5!o:��!�YGT��5w����w�>�M���n�F�j����w[L3��6	3t:+M�N2� �[����L�L݆�J&����wbX/[�A��s��0�eL���ͭ�4�;+U�:+,��N�ׁJ�T���)V%��2���>�1`wR�z��Aݘ��.��%�/-c���4W)OY
VE�0Wl�'b�F���S���ʒ�eR�4�9Z���ɀ��C�Y��)M��C���ţ��C+b�s��O�`�G ꊰb�݆��e��K�n4Fa�����Z�v-b�Hv��fõ�����+_2:ɔB�mD8	�W8HX.�j�Jd���7/���WK�_D�emn�cn�N� ;-��{����0���8�VQ,h�|_"�v�G�̠mڨ��_kj�20�oFu%ܝ�O�^��g����|��lq�ޖ:���V�8Xh�y�n�5�g�ʧB�֢#̧��=�|��.���ڦ���S�+.u�W��3U�Y�@A(g-�+��G��)u��e�.C�9���úT|{�r���Պ��Yh���=\�����u-��w-��^�T�1I�2�t�	�K�Zy�0 �1r��]F��%c�����2��G�)N�\���`�N�J5C+�&��k5!��ƀu�9C/z
j��K�9���V���ͳ�O (a��Ґ�J���[�M��rJ�� Z��v8��xɃr����R&�
9xޮ�ܷ���C���V���\���C���<&`�[q���yV�n�R�@��C��eZ}��)��t��[��l���Œ ��fގ���e`�)e�<(ywuEՆ�N+>��<lX�؄�!�}���0�㦍m�7�W��ehm�f�v��q�X��ҁ���t��8�)ݖG)�]�:�}�2uo��r�O;4D.�bث���Ҵ���;��zH�M�y��4ӭ�������`@�9��g�9�M7��8�)x2�������qФ�-ꚯ��c���v��8���V:
c���IW���ڴ�6�+������e��v��[B�1�=�X�ӹ�NB��6؃:��"���ܛ�y����D�W�d�%�O�c9�u�&4�Nj� 
����]%�"�l���NA�|��u��ȃ��|m�3&\ٮ���V������)�.�"3J�/0v��ln�z�[�W���AY�gT��AZ]��+2;�W*�-��"��q�w:W;���k���z�u9z�2�8h�ҷ��k�wY�DqA��=��sӣ79E�:2��#Z�-Z�@[��[���甋1���JJ˧{A=���Rnѥeޛ�����*8�7��+5�����;����\5��O2��Xy+����5*vڴ黦t�Ѓ����Sq����]��Z>�j�A��
�:�D�Uܣ����-�,���Y|T�!�0��7)�0_$����Wӊ���<�����u9�X]��8�k�	�ԟb�z����ܺT.�_N'�S���63�Mm��aDV�Yu��	8m;Ȧ��}���Iz�9L�{��V��k�f�zq�;snfn�'�do�V"I:$���5�]sO����z�u�\:�Φ��:����Ҥ�B�<���^��R֙+	)R�:�^ݗo�SF���G�gEǶ�5yN�'IϤ���}y� va�ݖ�_s¯�߲�C�<�z|��ʺL���;3{��꒜�{�_Gmp���#2��㜨�u��撋ݦ��(�\0v,�|��odĳ�ηu�����7F��sfT�y.�1���~���nG\�M�=T��(X����.53�(M�Z�,�����#*����j�M][�t�A�];�JV�l�����oQ;s9�H��/���au7b��fI�,jY��;x�̠v>y�4+=t@�Ev�َj`�
�K�9��gMX�Q��k[�R�.NnV$��o9:<ġ��[��ϫ�p؈�V���R��đ̙���X��Rɟ]͓w)�r0�YƸ*��P"�N�:�i��@�D=��;6@���R�>�_��vgv�åZ�iA���n:��;5��n���i'	֯�m�_y�V+�
���{1X<O$WVf�j�<���{_ļԻ/�vF��մrȆu��-�)�$bc4u�E�[���b�,�:���8v�ݙ8�����Ǆ Hу�]z���ǻ�%���f�Z��zf��}�;=�D{tpw���X����++f�F��@պ!qC^wpt�Y��x�e���˩���\V��y�]4ཬ��fS��j(u�6���=�L�[/���mS&�(���*�R;����ɞk����{f%[fvVҴ��c5�.�c��Su�r�ƃx���K�VQu����bÛ�wu��p����E:��$�y�`�t��j|t!*�!�F��|QW}���^���|�x[�^���6\�m�e�C%��t����ۥ�^��I7T����Vvm��Sm�d
�^a�n���")�V�K9{��s���EE�Vz(/�����_l�`Ѩ;wM�����,s���f�.�@68���j����#p3�6��z��:[�ږ��:�C)�.�N��X0�ϛǭ��}����(Q�SH��M0f3.�R����3i�U�so�#C$�y�w}��wF�`pg	��)>��g��u�K�]6����q_N��Uθ���^��E�6������������|9<�J��۫��:��{AU�y*��n`�#ӛ�PYO�<[B�����:��x��;�
��AEM��e�)�s`���;n�+�D轝x���+�|b��!�'A�wZm+��G^Y���Λyc������<�Q�K�>�ݺ.�'8�vf+�V�^��$C��WoY̏F�B�:�5�vt����}��r+�7��#�E�w�V���i�"�h#+�r��pŹ��4�b���$�:��";��6��*f)
*�=,]��k`d���ir3���3�*78Թܩ,㮳f�%��=t�9�
� т����Z�T�Bv<��y϶��H��3s��峫<b��Fk��7� 6��M��;{���+�p��2�ܱ]����k�n]�-��d���P*J:��{�O�����]%)X�x��t*���&o�m�u؋����1`/�\3��!��c�����dӹ���2LŲs6�I��s�����
����u��<)<��we�s�w�@����uc&��^3�<��	J�Q�c?Y�:�¾.Ui��܏m�+;U\����U���#���=��ԛ�)�2���ٶ���7�6����Iu����6 TtgT}���n��dZE%s��q���y:��R�y��x����(��D��g5먱�l��A����ũ�|��YYp�3V:������q�w���W�N��2���oJS�8(@m᷷�����ZH�k�0v��8WmZ���v��Z�;'s�Rŷ(���
%	�$GS�U/��Aa��Au`57�'��>��/S�erC��>����N��xx�L�p�L����e�C������݊��.>�CRT��z}�}2~�\;ƭ�����m�8u�x(�G��X��,:i�쾼��}Htb{��_\6k1��Q=�:h�b/;�Uʘ9k�*��n�5Y�_{ϾƯ9��)��Ry���T�۷l(8�k��%�R	�[9� �mݎ۾#)��p���f�)�=Rl�i���岇s-����vV
5P��Ra��0g�!�:E*�4�y$y���D	c4X{�S.t��k�L��r��mJ���t��K��}Ru+v=LUM�n�«*[�^��]�&�����OA����3�����d�A�[c�������;��{��B��g
�6d�3r}6U�����::��u�C3��$+ڒ	Q�Y���y31Z\w�>�i�
��ì̮\:Stp#�]����'�b���;��v=u����M�^n#gg4*��]4f�ع5�c�H��+�Ԏ���z�v	X����mB��o��[jR6@	V���YM��Z��k~*��m��ϕ2�]j��1 ~Յ�^PP���嫱�cշu���7zUkܺ�Ɉ�n㢹�:����mfs�n�ջ�Xo���S�sJ�1i"� &���)Aңn!xkc=ݺ��\jWt2�"��C��j�z#l����X�64�Nn5Pe��V�h��o�Kx�gJ{) ..�G `v�6]]��,a_[A+sgT�r�tw2�	XV	5�ص�%nQ���'\��o;j�QWf�'M����!K9WS6�Ps���;8��uGb:šS�͕�A\����a�/�Z�K�Sz0͛�2���yg��Y��o��iŵgHӵ����R����!J����A���J���"���([��䲄`�ws�juЮ�]%��c���ivfv���5����$;6d]��;��jY��Ua�6��v�;�ڢw�pTV��$%.j���=ۋl}��c-u5�"��Qb��ފJ�c��]L�[ad���������4��4��n)�L=��{��*�Vm�ok����>����{�o\��\k��r����e'J�tS����� �{#}��a�\D�Ⱥ� �o���v�����B su����ʗ'O��j�5k�\�5�ge���ԛ��n>t��>B��4�f���˗��^�UO���0Ƞ{�\H��v(�6fp9��f�ΐ���N0+ZF��$��:���i�*����nR*����Pv7jA���U�;+������y�M�i�fE��V4�a�9y��!&�� �G���)wL���]�9\��3s� ]�KV�V"#[�G(��["�D|7:�� <]�8��>۟\�9��Z���JV�.F���h�;]w]�E2��ϯ)�uN�l +6���]K�;�3)�\�ɵ��B92��,]٥�*�v�J �-ڙ�*�a�b�2����S4�\���a���� �u	����A�io�.;���������"�o��*���E�}������D�vt;�,��ˢ�cU]�s"�2�v��(�u���ԝ�X��<�C�6w/����r@[��<*vm����[���;C�Ha����M<C����BΧ{8P�a���I���U�'J���-}t`��S�*Rj�R��Fi�KN�cHW���m<@`��wM���2%�2ͥ��^s�� Ӻ�>|�����\��;&ފu�h�8IiW��C���"�	�j����JImt�oj��s_q$�������Y�s��k��eJ[%�YY����3��L�nm棲���e"*�B��NY�6��KC}b�e	A3嗭�Զ�����Eݧ�-u�?��Gjܧ]�1k��֞3��7ʯS�3���!��f)�ox<��g��|.��N-��@�� �l�k�Y1IEFs.T������ˮ�UȾ����tx�'�w
�5G�j-�������rp���&�!���}�V�sWg���R�����T+�w�aT �l;�ݻ�X�X1�:��+���Ĕ�m�F5�ڮۺ��9֔@ ���7�_vJ�nPF
o���L9]G�rx�s8Sc+%��5�a�{���^�Q�nƎ�3���vu�\����M`����O��V����ި�m���%s	�Paׄ��MI�2��8�O���j�e�iE���x��}JŴ-ҮR��M�,ՁZ�M����ےqWB��9��Ӈ��[���e����6Wkp��<Z���wC��"����ΥD�[�Vͻ�Z�:X��J媾�3��)8�r0d�~�=�8�q�¬�^�r�h��]c����p�}�Z����A����cC�v���C��Z�ם��)Oq�F�6H�����UkIM��X���O�s�&7b^�z�;3
Ώ6�V)�LI�"[�^�C�+�� �Ñ�ݜ�!VW�݂4��U)J��U���s;0�E��s�v�duחc�����B�>���4�<��c�.��Ir�f��ܭ��B��r����#�7�e�7�+s�q�����&_(��=R���S踖��+F*�ҚhN��L˒�� z���H.
�:�����a:�n�}OG��6��Z�\�zN\�:��4�e[�S5V�r��p*�4#����g5ս>�S��"�@S��#]�m]]���@�b���(yȺ���_#��Ոd�9���Y&)��J�tL�r��F�[�3)t�{��	}�Vy�U����8�ME�t�U�0q
����@�|�KI�f�V���Ż �}�V!6_6�5Ԕu�|����fJ�跔2�n��X̧YՉ�$���ޮ��qp��X;;�]3Ι"9�(N,�G���T�;C��}ܯ�g��:粻��|���_vju3qr����xm��`dL	M�W�9���� ��07t	Fr�ѓ�q����2�3�����{���z�U۹�s�#�)�I,�7y�9dU�r�_xx{�����<=���z�Ê�k�sB�z�����^Dw0	(:�z����ĮK{��i&�z^,�9�E���F�"�*�qG-�2�2�%�U�ke	r�`>�wjYk��%��%��Nx���7xz�&����tPzܥ����Å7�wgc�������Y.| �@h��J��[w@<�Q#'gp��
T�T��۫l[�SyݭZ{ )Zݑ�FP\�=&�됭OZ�9/1�YY�Z
���}s�]|� ��@ʜJ��Y��qn�V�L��B���Cp�C0�A�y�"�.�!YRȫU�Y�s�G5V�(٬ϰ^�<F6Nz��YAњ�Ѕ���5��l�X�RXwC/R�Z��>��2�.'��i��_:�f:Zɂ���v]�$�`7�X�p�Z��p�g�6�#0m�m����|���}S��;;l d���Ջ��՚�3WE5��n�ݞ5 ��p�Kq#��ʽ�ҍ� $�c�Z�8�f=Z��O$���9�!R���ʄ�)V��`M{n聓���Kg-�۔dSAh�.n���9��:] 5hD�'v�7�0]���+gp�C��,��j�0ovq�Y#���ڶn�J�iRtn�=]�h:�:x�"�Ί��g/`<�;���r�ܸ���v�Q9��P���Auյ�.�d��<(�MG/;,��ӑ�������Vu`�5�IYM}Y�Q)L2��Ϲ��$��P�u�y:��8T��gu����ȝ;���p�����V&&�h9R��h5O#�i��+Sfب�ø0 ��h�q�a�yYFa���-�HҐ�$���5o�?)��Y%s�[,u�����QCJ�ZD��\E��C��ҬC ��wtrS��醨/�$r!��	�r�x���gyx�mơ�,p-3oE �>t��[�cJ�g2�R���&6ľ*"�u���j���XXN¾7J���0��)w12�$�gMrM^.����ޟc5�U+U�(+�Z�$�8:��p�h��축͹���S�U�J� �]F�hgv]�X�2��v��r���R�9χ��**WR�� d���!\?^��ҭ�A:r��P�; z9�l"�9�(`�\Ҭ�GZ�4�mVѭ�����^�>h5};k͂�6p"R``݃�e�w�\.d뼫�v6�6�:� J\�0(R��j˖Ԝ��M�u�9h�rl�V����2@we�Ǯ�xLh)<�i1�E\�[KWee��w¢�=��l�CEe����B��U���:����|�d�]�D7���������D	[�u�o@�������@&æ��Ұ��Ϥr��u��8cI�:�y���3b;�A�2Om��q�yQ)}�Y��"^>�w��`광���~�nl6�q�Ŋ�;�#��U\�TwA�HP��قt�RuG�����']t�����|Q�����ub�!��X����O�庱N�]���wOi��y��Y��5�j��YK6��^4i
�[��[�w0	��ؒ����W1�ud��{;�3V>i�����.���s��<�K��d1u%eTgw�Ӆ�P��K�JI{M@�˻�V`Ӝ�w���!q��;H���0G}���r�i:���}EM�5�J1{�8���.(6�^����Y�E�+���82M�`�
wB����������������6��yRh�^�vAyBR�ٷ��Y�
��oC}BM	]0p+��cڼ�:�R�E�WY�^�n.[���V��w(������X��iz�I��ƣ�=jB�ܛ�C)WS��r���Z��^].��
��]%�^<��2�mt��,^�`��Y�3�֯�t��q�'���-kšn���ԧ0�*H*�;ԣK))]ٙg��N�G���1�;��*�������c�
�[!C��J�(��U �O�D���6WP�J��T�ҳW���,:�Xl`��i�lѾS�JMAY��n-��*��Uӕ=�8Ϡ"��^U�wi�t�֩�����W
$Cύ��v8��M�5bwG��)���3��I��	�r�w���'���5ٝ�4�d�L
�N��1�)\Ʌ��sC7��ov���y�(�Z�[@9n��6�W<��zqYy+02GwƂ�!��@mѩ��7�U���ɽ� 8�b�C�w٬�
����Q,͙y�	olA�hQB�Q���wq��U���!�".�m=�X���i`��XGv�o�5a�f�ث��`O�*���Wy"�O��Y�+��2�-!���6���.�b�k���v�>}�\��n,�9�r�T��;��6V�s��{�\.nv��Gn��IjT���o
�"�\�-N�F�Rҵ	�������{�G�p|y���N���n|M�{�:�O��6����J��G�5��E��__ێ�������֝����p&`xѹ��{1}K��/���Y� ${rᅋS�V�M6֌´��tRBn����5�ɺ�7)f���4[�5����7�\�LT�6�DWF <M�I�����2���ѩH�o^��Y��տH��\�Ӓ��/��-*�\j.��3�{�+b |��H����&��i��������pM�ǹ �Mͬ�=���xrR�Ys�PΗչ.���R6��C�_I'C(ܫCX�F�"���1�h];�nd����/�GIWfb�:�,#:s��U>e�����Xb>0+���?E�˒��¾e�����N�n�pp��q�w>�OT�t]=&tA�0z�s��`m�>#Ҫ�����Շz��V��i�:�0T�*[N�n��� ��R����nH���(@$���t�{k��Hv␚�}(;�[6U��E�EսR�q�z;>�mnmܘi���n")���WJ>Ҍ����X9���jCh��M�k�i�ѦP�a� �N�v^�Wu2��ǔ^А����-���4��ٶ�Hj8�`�jձhglŹ��իIح8�x�_,��C��z�5�Vo(�7W�$��������8�]ث3���#I����[��G}�.6륈{ ]��E`�+k0��Z1D���1YL�*
�!��1`�;]�4��_Q�[;Q#�_i���T�@�<nl��	��(
�X�S̈́7OnM�V)���ݼ������_-H�#����o;h�jrt�^�u�c��*�B�pPc�A���/0T�v?�h�0%r�WŞܤ�U��|q��Z;����{/��5*��ܩ7Q���4�ۯ��Ǡ��9G�l�Wv��Hu��ͤ�>Ki`�*��4�=�8�4�j�����x!�+�źj�ek�윀 �GX� 7b�֒��px��%V�n�XhaBVN��m�(��m6(j�T�v���ޥP��ۼLtAOv��5k�����љ���1e�N���u���rBE�Y)�f�.D%,]� �Ҹz(ve6�v@Ӑκ�᱖��aݵ].e
�Y]ɍ.7{��8�*���=��oo�Ιp���S^��֜{o����v�_�\��T����Z�����,$n�v������}np���R��own�)�wn�#��He\R�P=��R���v��KrY[.I�f��xΜ�L�V�k	A�����M�4��$㲜�JX�XJ��+m�}�C`��M��jX�N�S'Qγ�۶UQ5u�� ���酖�:�=�y�:�l�oM�6*�go��sjӆ��
�h������)��$-R �9՘&r�v����RO:���qS[���J��B�'k0ۢ��2P�0�mԢ�L\�A��_^լ��S�����Ǵ@��oJ��L��ó~�s��IN����[�:ޘ&xxn��pJa_�X�E5e旔#]�)u�f�s�Q=/t�V�(M7[��) ��V#B��ǻE�R�凡Y,�@@��{�,՞j\���Ksk6�(���B��-��U.�����-s8䓯J�4��Jp���kn��f�r�ԭ_BX�T��ۦV��i�\Kmj��l��y`��&�-�p�ӥn���b�v�`O!G6�C��w̶vf���n�S�pyg1���P��X��{-Z5�Ћ�����U�EY�*��|�:gjӭ�H�m_vl�n���Gp�W>�gFeg,�wvYw�}��t�]�j=ʂ�>��Wׯ<ĩ����VɭÚ0cYP�_*�Y@�+����gn�H�z���l|h�/�8��)5:�]C 	�<�IYMh�QǪ���wnf;�!��v)v��~�V�v��˥���7/5�b�j��B�=!XWt���i�ko+.�n���W3�k���-�Z�����{S���A���f��n����P�e��nle��U0mj�,1�A�W#糧Y�qP�]���W\n.�-�U�׎�	ѵ|�Obr��:�6취T�p|m�X�[ǯ칬m�"����͕ä{B�X����E�Q]��4u}�Mr�*]rt��R�8�3щyK8l�Lپ���V�����* ����,��]�$N�꿶�̷O.IځIj� �f�]{2�QV0��\+Y�4-l㝑$Y��m���j�l���Ȃ:�;SS�n��	$��#�oV�N쉍�P�)2�4h���b�6%m�ͩ�
Z�$!��孇!��g��Qdd޻�NY�f��o���o�RT�����^-ULg1*	�m	r��)�jj���s����t�R���4�v�tr�^e�/n�*�X�j�@��<�:t�W�!gE�[[�D���x�N�/2����TA���BȤ&���gp��@�4�kH�4 ��$�[c;'@�.�Wo-0��d	>4�Wj��.���P�]����]�Ի��\�e�E����D��#Pi�����Ȍ��7;;i��̧:T����ꎻ�� ]����ܙJ�������I�c�c����Su�9۔.��Ɔ��F���'��VV��2x ����<���;]���6�ME{/,��`��o#����j��R��EWp���Ty����hQ:H�]�Zre!:�|���]�[�]�C�����ئ� ~h���ǔf<�c�Q�uvm\����S��Qr�\��Y�Ѩ6��ne#	�W�;ၶ��DRƂ�9�k�S�c4�9�/�U�h4�앢n�>Yn��*�W����Ҁ�`�+�A�x��25����+��_
4��8��s��c9VS��Q���3Q"ѩ��Fd��!^�4�q��[4J�y��nr{F�n'"!�,l�2����Ϧ��b�w���a뫥�w3X��h|"ʑQA���8z � ��rIt��6*g\��̀Cr�!�b�(�,l9�����EpJ>�=� ��D�C����	38�5v:�I���8���uN��V�݀f�z��Xl�YΛ��ŗ�w;�
�Un���}f��f�F���Eԧ4V�*�E%�.v�7a�$�T�	WA���1?��v+b�G̋��g0� M	nザ-�gGv����:e�$�d��s窺���y�x�:������d�ZT.�mg�t�kI�t ,�&C���@
��D.*ﲰȺEV*AQ�E���w�Օ�T��$���@��`��νþV��,��F��<3}�*@b��#�2�3��W�I�r�� E��7wp�AѦ�oajf]c�U��[zV�I�}��fl���b��ʩ}��8��N"V�7���9�1:�Z�oY� �S3�B"���]X����dZ�6N�qgV���V
xK��*T:�wo)�q5�H�c��}$�;�� +&/��9�l�գN��^��`R�.uw�
��YJ�eq�j������Fj��o�G*8d����O�u���(J���C��}9�Y���������Fp�j�!A��ɹ|"��Hp4,WS�J�vbԯo^i�a7�X��X:B진U=ҵ��L�9�׽ y�V��AH�Y}�ڪ�c�fhUbe���O��)v��b���e�|��:@���Nub��w�&˫Bp|z6eI�g3b嫁���_*��L�� L�)�Z'Cz���}R6T��Wm��f�Eec��nR���hn�����B�*}�^7��=r��Q:�d����IԚQk�Y��9d��n�fQjuD�`Ҙ�]09��I%��2��VjYe;Tg],g+����[xJcC�����0HÆ�d�h�2wU���I�P�Z�g�Ƈ����=��f����,��R� g�2v�*:���X6�m(�7��e����?
x��L3ݙK.�8�$�#lNjD�^��'>�x�7���Y�%�rQ���C��W]��\����{B`�ӆ������nud��R�Lk��n+�x!�&������:�����^m���8�h��K.��;X�C� m�$)il�I�kݘ�T�*��)���Ou*p��P���]EI��\J��+�ļ�J�F��B��ƥ`ni_[R-��wPu��cz���-�[��N���QR�C�0��V���47q:���k�;�\�oKG�؝X��Y��ޡ��l�}���5��85��t�/��.<2��"�[u�*��>�,Ǵ	�Bh{wm��F�FC���E����Z$�n���
�z�}�D��TkQ����G��x��VpR���G�;MVXvGn��yiR�
Vc�W�J+����4�TheUuD��ͺ��I��0x*X�B��Xi].U�HU�9y�*f]���s��	#���|����T�\	o
W\��T�v�1vK���엔�(��.��T-@IY`�t7f���9)ɆD��<�%8$�}m��6�wet��Ō^��߮N٣����+OLX�{e�7K���"����gU�+j�J��,�-M����/�{����{ׯ9S�k�s{Sw3sa�8Q��;" s�F�z�<�ՊJ�n"�m\SY�uo �,=}rh�E��b��SlVL�ntU�Y*L��:�Q�6G�aW6�z`�'�cQ�]�mW@��C������s8.^`g-�V�l�4�֐�q�me(�*͊}�p3/[��O�����pO���������ſ"D��9&H�����b ��;M��'��C�.����nv5Qi�
�be]�����j�$� ]D���t���we�:jB��<�&�Z�uF,�Z�z��RӴ��5���@�n,����=�M��;��[F�r�7V�fɎ�J��=�!׊�,�e�25[D�n�gi,S�2�g^m�30&��[�DM>@�L���SF�P2�o�`t��-)�U�hm=��靺k'�R�B4�*�㾣��<��BFf�`S:���oL�{���W�%��t�'��R�Y�E�W����F������cG��|��W,ͥu����\�{����&�qx�K���Qܞ����ya���VP��?�<���(����O�,������M��R �)�U�.����x�❄���]�ԉ)���-3{w��Q4�f��J�uIl��P�N�.��͜�C|M�&���Gy��h���5{Y�ݎ��l�z��o�w!Tn���d�x��g��"8Ɗ��'��������Z*�đDP$
�y�������U�ww;	�`ۺ���y�\#F�]��`7غb� s��G9�s�9e��
7:B;�tq\����Ӻ��.n��\;wIwqF���u�rwQ��N�ˮ�Bwl�4cF�wqD���wuqݹ����p�Nۑ��8���E��$�WHR���2�[�;��������wDswww'q�R뎛"�]��uwts�ܷwN�;��W1�FL�:�9N�sIt6K�(�wE�]�wu�h$;�r�sB#F��.���\쎔n&�I�5���+��uҎj�v9�3K3��)�������r�	Q����w:ƒ�9۷I�]wut��'w,%�.�l�k��7�"�vᛗi���]�\�L�0�e�\.[��E$�IFH�(2����B�{z�������a�%�^уZv�ͻ=�I�Sm�b��.mɳP�g]l�[Ti+�0�L��1��;E��P��$}���Y���v���ȀU�@�����3\-?��h�[���v��@��n]Z��f���#�"��-✻bz����_����"��1�a�k}���:pu�#�����[�����]H�x���<���x`�=�ؽ>Į���j�ݔ��O_i:|Y�j:K��7Wk�������ÙH��cys�=~��4��-�쪵��*4E0�3�x�[Y3���(�9ki�P�k�uJÁ��>��m�,T���]]��W�����{m���=®k�N�\d8�����V��/Ω���J��md���E�u�Y����}���U��c�'`*�qRhV��Hs��p��1V盞w.��2 �ȩے��*{�QQ�NW�ّ�r��N�;ŕ��X�y0p!E8�*���>�VL�T���hv�K�|�7lr"åN6���GqPI��ʈ�v��ׇ|�P�X�!�ə���כ�
%�+|pr�e��i��(�mN��I�վ)k�w�9��ǻ|����W�0h��)b��?'�4M1b¦3�Ed�^�3;Z���G��Y��ǀ��}�+�72Jͥ0��c��m���f��Nt6�"�.�9��^w^���on9H��Vㆁ�Q�z���IG:�E?��.ɫO:�qZ}�z�'9bᓜ|��U��V��^�l�d_=v��9�i���}��lT�hp1Ӌ��R:���3�B|���W /k&u���)�宺60Kj�u��8']���bt؉d`��^ݘ�o1��v�UTD"��^W�N�$KU�n�GC��b���FEMZ��D�d\"lV����yCj����]��w���� ��ώA����\�z�r�8��(e�A�cg3 H��;��.��fmj��(<����|<,��+O��;�i��a�Ƴ�o�Ҹ�1B���EZ%c.�W����M�n�9�ʨ��a&GH�ѵ9������c��u�+<�o{�r�ق�}^����`����&�ʃ�����͝�"8Y�D��^yV�-�l�DR�����}�
5�.�v�C���\�<��v��*��帆L����a]Q��ԀO�>ya!OsZ�����ez��3���U���F{6�TW3��5������7����.4&&�>*��>��QU�I.�;aW ��Z�W�J�ۺ��i��+�H�vU���c�Ɣ��YvL�m���t7���W#�J�����/mҼ��&�\����ǋ�MG�N�Y��{oH���6��W�-��V��;OAU�rj��u*�T륭���G�@!(�n&�=��`�ݽ\�t��+\O˖E1�=
�^,��z�L��:���G�˄"�왇B�2wop^v��t 
�����AM�V���#b}S�&���%��do�Wx����G;��r�9ܭ���^ߡ�=N8�]��r�YM߶��28�Ʃ`���wc0���#7ݯږ];}U�H���<Ȩ�N�{��J3q�Շ�m�h���Y��͒�bӜY���d���$%jU�3�:^��:*,	R�"��4Fsv܎���O��}�V��Ţ�rp�xs�d8��I�1̬�U�_X���tYwO��_��gƥ��F���ٷ�{�2���k�O�H�z@iP��w,a]�ف}�w���7R9�Y̮��'��j/����	�/+ �m��[��d)�W�#~$D	��BzW��V�C��aki�ۥ�h�.1��S��C�K���/�B���	����{Ύ�}U2�s��}Cba�q�E뗦�:0��EIӣG�r�F�ivd��茹n��_&���&��<��zk��z��M�-5KݲT�;�K63Vb��k&()qS:|k�u�˚r�!�c�X�,i�3��+^}xj.�)�t��q�����T�`xE\`��@����"6��c#4>����ʹ�3�$����b��Τ���a�G9Tr���1��'�;����y&ܸ�k��#�^��T�-\ܽ�8���^���o�x��s� aκ�URFň��q|��]C5�'�۹:��v�S5�WV>��U���6����A]e4n�F@ȱ�)��T���V�*�Y˶���X!������;F�~����DG��٦=
��X�ia����y'˄����l����2��W2����j��Ӛj�2(s��.W���s��{`�2�gޝ}�VT�Ʌ���q
��p9e�N��ꞁ�aVq�����L�`��YV�[�{O�3���R\
����up�iu�aˁ�N[=��t>�f��r,�lv��#�"�y��<E]�_�z�mL�9�>U�J��-��bC���`���y�2�{�#�ߔ%��ŒUx���ԤR��dK����^A�R���ո�h�)��C�z�W{q��>�H^�7�:��@՟#�*
C�^�*�U��]����\�=����Y�`��U���1�i�~�V��q�����c��^�M�ޱj�ۮ읞���X;w�6���?�o��������]`j+���oe��O�Ϻm� ���ڽ�\+�0���A��̏���*]lۺ�K2Zڔ��tK���+z�^�U�T)�eBf�Rv�9�OB�W��)}[Di��D�w?�fGɲ!;�Sp&�o]���+��#�Y�����Jv����r26�N9�f3�=���޾~���4��}��~m��N�3�����^���D6��"+���xHT�M�G.+�6v{�R��=�O)�}y�Y�ȅn~�t�"wz�;|�À�g��j�/2�5��^G�KF��b�/O�I�o�TC���0'N��-8�%un�ې�gv����(K���̪���=�6f�W<�^Ώ=1h}~8��Y�-^']�1�a�~�kc�=���]�|�x���ډ����������*`��k޹�O�+��+B��-}�G�}@�ye7^T�[D��ᐽ�|��rS7��n�~S!�9��SUBumf�Do��J�Ƿ�P�:�y�Kx�D�S�T}B%N_m(��`q��Xp1��<��n�����yS�82�[}�)���E@L�U�P����N�\��8
�Z��
ӿC�l�R�n���ȅX��{��&�S&V���r���#	��hqj�A��5��Df�w�Y[�P��9M��d.���X�{�bͭM��6o��
��bU�mV ����ڕ\�#iX]����y[W��ه�wy�[
��D�9�J5��v�{��/;s�寬z���*�}�v��&�UD$9�G�&����u�
h�:���'�G��]/d�}���O�n�2�$��I�`����Mz4p<_gI\N�:T�n�{]�a��:>�s��\�p�(�mMM<	8�.k�֗��^�8Z$=��{7�"�TTM.v���2�熟(םADE#�*��!Ē�1n�yf��n'�{o����3�}cV��ϧ�g�"��Ǹ9�!������d"5lL�q�ȹ�u�* ߨ�BF��֧tS�(-uѰ[U�!�ˍNwI��0��y�[�Mws�+9�C�UVD��(0)���h5[2����ǡ��{S�ǭP����~��SR�����j2��,Lq,^:؋��#��4vLL��F��)�U�ϔP�"�;�5�Mgq�2���X����_��p�r\��\Oʁ�����aϨ��8�����b�x��'S}�澿XmP�XS&�jb50���@�Nt�zh��8�ġ����c?S�Lo�Q�`"���C��bB���%�)thi`ZTVҥ���R}j�E��{��{.�}�8`�r����6��Q��ɔ�8!vw�F�W���p����Z7��c�� �rnvxЍ���n��Ŝ9����.��"2p6,�(�p���<��^��]ya$괄�|�����r��
�4�w�l���C�&�-O�chp�<9Jt����ߎ��q|���B!>��2�*9��N���{k����E�d��3�"a�C�@�3�DGn:,e�Fs��3�w;Av�o=�(��uK#t�nϤWS~�d��2�j�Sr2	)����<r��X�Q]��Nw�s�Ew�__b��s�Sb����Ѧ��s��+l�g�fV�U�/*3���ڬ�k~��W8ɨ�OM7<��y~q�|F�ѕ1Dl>$������Ң�����{0�n��*�Nd�#qO��t��.!�����VSw�E��`4)I�����r��Ќ\�ݨ��=b��N��ʔo��TMN�zư�Faq�j��3��� [����1����9t/ՠ������!��q�j��^��E����[�
T�������:�ً���*��l.�(m�.J4=��
U�؃�̅^襯�U�v:*iK�ci���ݳ*�_읻˩S��X�XX7_5�oM�$h�X(nDH�n[J��r��wh�����/�ق뮻�el`>,��ղ���Q��J� YIM�L���+��J�y�MW��݀���}LʚxX��!ZDW���X�N<ǰF1�Y�:]���i���p��ރ���p�E�7�>H�z@~���{�>�+��2��D"���`o7���ś_y���@���/+ ��"89�J�Ԥn���}�.��{�ev��R�Y�����v1�2��Fo>�F�NG@qnf�/���6�f("#L�̎gu�XX9A����^�C�K�hB�W����0����+�vh�r�F�W�^'�o��)�Ckz)]h��ʦ֓lFO��;:]��Z����pp��l�p������2�q�/��U�[��-��˻܏;YS�Y=B2C�wO�	s�lu�
�����*��^�xT�x4���/K�kۘ�1�]��u���4�y�*�{㙳�A_�)�~���23�fYW�`\��q���w��\�C2V���u挭�tnW�o�DM>���T+�,4�>ֵ�����=��|��|qUN}A��e���{xt暀쌎d�*�3�S��fZG�<^<P?/U=�C�4��e�+��#̸(;��I�	?��A[��/�z�#��-�q	<72�*S�M�]�7�����#CmF��d�����ct8h�<���F � ̙��e��C5�eS���/�V�Gr:�Zٶ�X���;�4�B� ���:q�
��c��52�Xz�so�Y��ے�e��9�ԧmd�z��ݍ��].����
��G�a�5����ע([��r�������r��s��(';�f�k�צ[Xd" l�����R�u]Nr.ϒ�Ut7J�OՕ�L^�j?�H�kj8YK�����~ZlMN�_���ŒU dy�
��$VW`�qOgч��5�Q��.5��5&��C�d����f�3���N� {V#�!ʼ)�a���h�|�<\t�k�l��m!�fq�9����\b뼀�z��^O�|�"��u�� G=�dI]�5�0^=<�G�p�oz�;%;l�ޖ�2.�ۡ8���tA�9�Qǎ�TF%�;��&&O'5�C��#.�������D6���ŢU�3^�j���k^p'�ri	~,�B&Bv"{�$�95w+���P�|�À�g��S%���+�Y��Skg:�@=�tE*��q���_�R�魅T�W��l�]oO3�K���εs׍���n�||N�ּ.�.#�v���������妎M�K��ם�\F�:���)e�>�������뮡a6����%o!�� lZ{�gQڭ;�d��<*�����wȐ޾5`�JS�R�<
�{�`��ɜ�ˁ�ƺ��S\�X���t�{;8��k)^�,�m����T�0��6�%r v�ݑtz�u�ħ���O�%L��.#�߾K�>���u�N���A���^���tI�Q��P�h��8�MI�j���2�q0*�;�������=�~���CT�1���{�F�t���ԷV/|tlK���~��>�����J"��X`uJÁ��Q��w����װ�����X3��ޏ�9��"�b
���^]tm���8	���������㒳�z2�D�����n)b���QA�\���(��D�u��h�y�롾�|~C���u�ѥ%랂;+��X�'��|+g�oG����#B�\I���y}{R�����MM��D�o��6�cJ��=��X�a�-ҧ�c��5+ON4�����O �f�->Xe�ѝ:Fí��E�D֥o�s�e����6�ΰ��M���n���E�3�J������9�8��cL�}�g�n�5����玗�cOX8ϲ��Dy9�Ht���Ou;�<Q`h1��1"HzLPٞjt#�;�k���ڿ_��ˍ��w�,];WY�߼'��tQv��6�*A�%�XF3.�cc�!�5���b�(G�u����hr����
���d��8u p)w)��LH��en�Oز��!6��ڃg�d�wL ���ei*ྵ)Ij�cx ��s��P��x\���f`f-
�K]�3� hg��C�PTI1�ꎶ�����N�5��-0�:uh�Έc.�m�J��e��ʹ���ؾ�)�go���X�8�+if*o ��EW��0�����{$۳����y��"�2�q֠}���X�vu�IX=�z����9�9q�ۂvͻx'�������A�������4�DX������u[�3N�#N,�okLWӋ��l��]z�x {.���G��s�P��a��]�t����24gc�Z�E�&�W�pY3'";��V)5���p�H34<q�TA��v�
4�5f�yv*�R㧚��I�i�8q�s�;\����s"��m�w������K��4��􊮘�`ŝ�}{���7��X�2���࣐nMgv�t�/v#y����2&�-IuΥ}9��R��%�q��t-7����v{T�Ukx�s�X0�|�m_T��1
�V���8�+L�!n��s�Ay4���x���6s|���A67����v�w{	<ꝕ0_�Tꬉ7��N�쿝5����<�vr�W>�2욕(���_ku��W[3ltz�7-��!�X�$����ck&+�p�Ȋ�&�V�J��<�.A���b�2n���!M�6�ͳGQ������]ۚ��.C{ ����+U�dj.���4K�������s���^࡛�]E4^$z�.6�m�,�!L�X��v���^We)����Ãb������q��)��m���k�ܟKz��vg9��)���u�٦Q�q���F���6%����t�n�g����{���GI�[�}�td8P�=T����V11��K�6>�v���`]����JėXͭBaȮ�b.I���Gp����;-l�����zq�µ��v�d�Q�����k@u)����Οю�u����rum�u�+����C��zfU�`��כS:�>����Υ[�d�}7]oEC{� 6�oF�VF�',:U�� �XMŗ�Ms����WT�fRƐ�����.�v>�	�i�%ڛ��K�jQ2��޶�e��Hɦ�3�8e�����[0�
ɏ�%B���X����Ɵ�ΙJZ���3';�S���j�yh�e�-���]�r�aq:"�f1)�Au]]�5O� E����sI��e�9�63�c�f������x�d�
*x���Ƨ]��OPש�#-��X�{s�hi��O,�O��0`5�8Ŝ��-n;���P!O��钰NV��8`jv�q�Ϋ�V7V��Y��F�=��s�pC�����_������7�`��]&&�s&勄���B(1��)�u�v�
�9�H�!A%��00���Gu�u�L��ܮK9�r�wp�$�Lb�F�3L��d�(�Q�N�F�"�1�ti�n�H�	C�"d�n�&�N�;2&4JT)���K��0�ӷsn0�Ac�]$#��a�;�ӻ�"�M2�Pw9L�$��g.�0$�1�����%4�L�.].s!���wH%g:h�D8QEݷs�;��,��� �Bw\�Ʀr�#&.n8���r�t�����s��%�Ċ7.����g]�g.�$H��CD�HȎnEsu$��qn�:n�&�����F/��������������7�Y�s�T'U�������p�n�����Ĩ����90%cZ뫻�ϴ�q�Di��:�iqfq�٭�^�����+�ѽ5�����z+Š�_ݯ\�+Žuy�k�����o�G���m����^+�����/�����|������o����snU�\���>���dyǼ`��0�{�K1�y5�Uy����}����m��[���1o�s����wϿ}��߭��~o�_����oK�w[��7�E�Qo�:�y��o^u�oW��_�{_V��[��W��|k���m��V+� �
������D�c�!��)6��������_�Oޯ���,/M�m���>�m�ۼ��o��<���ssn��~]�ʹo�sz�����[ҼoJ���ү�4i�;xۖ�����^F�<�:���g�~�/�,l�ߧt����H�φ|y�=0@c���*<���7�ϟ}o�~-�/�~z�kzW5{����η�x�{m����6����r�}��y���ߊ�ߗ�o�m��o����x��z\�m⯋����w�����ߜ�.#i̞K��Q����8�ϫ��8��5=��~��߯ž����o�^lo�~�k�������Ѿ5��|���k������y��zW��>����k��������~��1�3��{�>���`]����"w��^п� Ǽl��#`
�����_���7��*�^������͹{���+�����_����^���}m߾����\�[w������_���o���ﭽ�^q1�8����q�"��w �u�貪���+~�y��G�x� dxT
[�x�����x���}�����^����+ŧν/>���+��<����6�;�����~-�\�۽����m���{�D�pǪ
���.���c�H��۪u���z���@��|�E齶�W�����k��߻�������������7�x�+�_�׋F�������^փ{�u��K��{޽y^�u�����g�U�s\�//����[}����ޓoV���{# z� }~yoG����o�}y�O�|m��~k���_˥����oM�ۚ��ߪ���7�oK���<[��޻W�����r�W��7����m{{W�_�ϗ��?/��o}��*���]޷���{�=J�����_z�7���Ͼ���o����<ޛ��m�޷�~��~-��u�y���W�O޿[��ۛ~�w���zx�����^<m��_���o�s�W�{�f��F+�b�`9Q	�6��C�������u7(
M/�]�p�tE��H���*,<lw^<f���ln���Y��yt���1�5��<��'T�o-�{7^^�ǘ�]u�KL� �o��؊��c߬E{x��������;�j��L�x���g�qk�������w[ǌo������֋|��ﾫ�}m�v��Ͼsr�׋��������}_Z�/���/��Z+��<�~5�������/��&��ߟ���������}���?}z�omsno��m����W�����ǥ��~~�~z�x�[ݿ��W������;*�>v��߫{o���������:m[���~��2]����{�������o��h�ۺ����W+��[��x��~v���湧u��[��ޕ��z�O��/����⽭=w�ߟ>����ە{]���o���ۛ�_O� ������{O���\Z��5�����޾��no��/������\�-�x���|^֍���_��^>+Ž��TE}_���->u�^�;���߭�^+��<�7���ϝo���<�֍�۽Ͼ�� d�5�-�~�z'x�'~�{�����ݿF�6��?�o��|m��Z���K~����^|���ץ�W?��������\ޛ�ί^�o�_˛�wu�<c��}m�Ey�_>u{o���[�����pxL�{�4^�����_�����=w|���?T�t�	���] `��ϟ|��ƾ+��/>����c�������U���6�:���ϭ��W7/Ͻ�_��x�_:��6��η�~y׶ޕ||x>�F������"�����i~�,VbV����v+�&ǇG���t�(`����ߞy��|W��_�~�z�^-�^����[񾷵x��|�祿��}W/���ʽ~u������_<�^�~�k���{|�ꊁ����1�t	�O��(Ugu[���;���<!�>��\{c�0+�������szm�w�k����o�~�y���7�ſ+���U�ε��o�y�zoKţ��������>}�ޕ ��c�����>o~F�}}[𝬮���t��+���)
�f�������ݯ}��zZ7��o>u�������������ߟ�~k�����x��~��o������~^֋+���|����sw�=�O��T=��}|-wӵ�^*�����{o����<_w�����ۖ�w����W��ۼ��~��7��^/�����h��_����_��h��]}[����^5���<ׯ�\��5�����}\߭�z6���@���@�zBt�̽9�JJ��;2�����v�������r�ȑ��q/`ˢ���!}����W�ʘ0w̵���U�Z�j������k��:�p�n���1�MfE:N]����1��T�
�n�D�Ҙ�J�8�A���i0��Uu��LU˒�@s��Q�I�W���1�"�w}@{\���}o���}��*����}��zm��_W��Mp����ž/��4w�Z��W��r�+��-�����7����o^v�k��[�]������.6 �/>��jR�Sa�xs#� J������o�_W5���׭x��V������^�����y����ߊ�����k�{o�n[��_W�����׽�ץ�+����ݫ����+�ξ����s|o_}��7���O.�G�,~�Q��c�}�������^>���ן�U�lEzߟ�}_��Z}�z�鿟V������Z�����u������Š���^~u�U��������m�������m�x���8�T�f����3&�{�}c�h������^������z�O���?z�;�_[z����zW����zo������{����
��|����z�o��ο�<��}_Z�7�߯7��~�����W�Z{�����l��r/ݛ~w����C�T��}��?��}�v�*�����y��o��~w�/M����o?{|W�;<����߾��~6�_��Ͼ��h�۟�{E�zk�\7Ͻo��/���'��G]�Ր+g5��Z���m��c� l��+�_�Ţ����_��ޛ�k�\5��_�;�:�U�<�?�{U�s~_��^�����������?��������� ���Q�}�\{c�1㛋RuK���W��ʝ�����}������������E����ƽ+��Z��n�~=5�/{��x��x׏���-�E�+ŧ�ì�TyÁ���@����}�=�r���#�7#������ ��8�޿�o�[��������Z��}����/��^?>��6���s��+��5�+��x���_��znm��}/K���6���]�Ǧ7��-�������ϯ�Cu2Z�]��ﳏ��|��\߫�^/����|_�F��������x�����V��_�y���^wW,������o�^�7��/�^����Ž/u�M�y��z������?�����?�╰(a���M�����c \zc�1o���|{hѹou���K/�ƾ�����r߫�x�?�[��Z��W�>���꾯���_��7�_o>�W���w߾}W�����~W޽�o��  ���d�&���ާ}����/;7������i5��.*̓��fP\Gn;��}�_]\�0	(�6<��`�8#�ge�P��s(���s�5�kxw�)�u:�f�������)��m9y׷�n.�m��M���C��*���A����靽���f�u�}㾾�Ƽ^>-����zZ��~��\���^}���۟������6��߯���o�ｷ������Qo��}�����wε����>���׍�x����]��p&<&`/�'L%�M�=uR��oG�����փb}��{_�i뷻���߯���wv��-�����u���h���/�����^7���ͽ|����zo��J�._[}����xۖ��}�����¢#�D?mn�H�ό��]����1��?���m�����wo��wm�|}�眴o�n�|�����
����o�uxߪ�wo=u�o���?/<���^֍������k�_�������n~��~_��Y� ��F�X��]�}�YX~Գ+ᑷ�_7���6�ﷶ�-���}W�ͻ�r�w߾z[�soן{�|��~��~6�~wW���F���o��^5�����j-�~��ο�z��\����_[���{G�}�fbZ_��Yۼ��i%ӭݫ?�[�7������/�}Z�5��o��7�^֟�o��}W��6�W������k�׵�=?���5��Z�������ߊ�/�>��oK���󊾮�7*���T8 ���̮Z�{*X���k��~~z��o��[����׵�U����=��V�x׍��_���ʽ7־�������_�A���ׯQ_W�Z}��צ�}[����������o�������W����q�#� L[�;N7����m�����������u~��>�u��._��ݿ�M�m�}o�}��m�x5��y_`	����#�q����`��Xp3ΧxEU��r5��y�׽�@��d쐡R�Z}��\½����(�`xO��Tޛ��N��yK����v矤a���{����yc��c��F|B8��/��@wm��p��<�<󮩁��JR���E��#�-��>ݗ�J?��h\�����;�/��=s���<��v<������M�L���m��Pw|�yX�ϳQ�Pe��U�5��=|�Eb�]�59m�eC�حb�{[�w'E��/=����S.|-%G�K��N�\��'GMY�8y�i�"���=Z����G�RĹ�����ݙ�o%s&�vve#���Յr���ȍ�f�U�qt��yô1�l���ᅬA�[��'\(u��.���YE�Z��z�X�:긅��y��SӬ�+K��(��ΰ��	�U����;�� ���Y�ئ�O: 0"b��fli�g׊�Yt�����9�=��S�lC�^,��.���>9��]�k+
~Rl��b9Ó$��Ɠ�J��.���e�Y�q�ߋ�[�/��#/���&/<{�z��`�p�+�_�.��XM*[笭5�״9����@X�67����K��w�-����`�H�ȸD�n�"�;#�;&$J�tlu�G�3DH�"�g�Y����^8���rx&렼f�Dl_�FDHUJL�J$��q������ɗ�M����^tS5�ѿk���}~mL³̚-�Q���EBM����B4�ދh��c=6yK7���p�T�>����d-4^XXN���|�չPv۽��f��8���Yw�{���hT"���Uc�Eu��E��P���9S�:�k�T9�+\����x��/u��s z�<�d{�B\�8�+��f�g�v̬�cKi����v+h�5$�9od��u�ĩ����m$.���p[wX���L�8�:�<c�'T�����p��,l���ֈx!���˾H��,�O'+�����U�`V��F�R��K�"����\Û������*p���7c�V�+�U�6�]޵�]"�f�"��-+{��G�r�=&�57Ɍ�y����hIZ���k���?�V	=�w-OA+�������/o	L���l����U�:��a�#}E�r��,�u�Kk� ��^��f�_�Ć�7DŃ��X%�Mr�e������>�Y��δ/�(����I�7��9ɬ���b�n�/}��&�	`ɑ�5V+�A"����N8�]�NS*[�gE��=V[�ϖ5˓e��s.���l
+���oc�۶�Ϻ*agy�{��J2B98�5�F�	X���5�@�6�߾*a��c�V�$���P;�H_�d$o�n���tT\�q����Z��e]t)��r������o";LY��t4�PB�G=��Q>*�ns+0U�4��+�Gu��I^]h���������Ѥ�3��O�<��0���`�Ӝ�4�V�1^4����>}�u��k5���$p9�����m�؋r��I\lԤLF�r!�!��P��]��λ2�c(��=�v�����������9�R�疥�E4�� ���eR��DwO���oܩ��kyY^U��e�R��Mm��c����
���Qu㴜f���e:�d��_̙��-D�����vM����=��ӣ��8���v7Gl؍�#k�[�~�*��<��>�/ u�rH
����b���ر^{�K��&��v�^:���E��ZW90�󞊒+�ӳE258*y2�ީ��9_`�e��	�ې]�R��E��OM`aF����m���O%� ���k36�'��9/}1h��+g�@�b�:Ū�a��$���^r�C�w��`�/��f�V�����kYwga�ڥ޺�k�и:k̉��aD���gAݠ�
�h�B�:���{��N�����-�>�W�=�gu捎w@�NF�W��U�Y��챾<�
��v]��vcϛ�Jd���7Ϭ<U\�'"��m_��U�b�X�͇�k�,�~P�13ѕ>{2��h4��e�+�A��S̸8�=�=vkWs�s'��9��r۴k�T0.�p��|�V���K9�=t3����S����<Hb����6�(u3��W��C��qb����x�+_	��~V$?w.lWo�VV8MN�R�[;\%��n�1\�?}��𩎭cӿa]g��h($��c3NBX$�@y($���ƵЍ:���F_
�I.�m��B�ۅ$e��u,K���f�R�f�7v�$��\Dj�p9.�E����E�90�Am�Z��"�p�����}��V�k:�UNo�HQ�1�B�N��ؚ���'��{FWނ������f�|X�e����E�%>�Ξ�0��s��٘Ι� 't�=�)�w9媖��w��F�p�t��2aO\oMP�2��!�a����;���#4�`��1��w7�nEok��Z~Q�s��a]��0B��Kz�; ��0�����dSn�n���h�$�ެM��M+y�e��9�}�&s��+���h9���>�
!�E��Yq�9P(ś\�Y٪�͞qq<M�a�	�<Q;�29�����"�E�if��oB<6��F�S]9��f�'U[>~��d�f\F�����8�tA��<^P+�p�܇4.z�/�U��]�6��46�o�<ګ�1�����ڸ�x}Y<#�A���i9��Yy休�s!]�l��t�Z:�����c��Ӟ\�!Ҝ�q���/�ٜ��t����9"GV95ϲXy��LGO�	�q��K�ユw�����ey�3�����MdxX<��ݽF��3�=n����$��.�s�y��^������_�Z��!�8�0�����n�Mw|�;��bɋ�l�|iu+u�2���[44�w���k#R�ǆ$9ܕ�V���̼��϶Z�i����1sPId���o��^0鸆'�7Z���{=��;�Z����g��tkÕV9G��->&���Շ:�a�rqي��K�)��{vߞ�
�����]��+��i�n'fQ|��,p
���+��jٮܱ�T���m����R�<��w)׳C�>���ʨx�t+�Q�\��F�j�����y�o�>q�=xS&([�n{^S��WC��MקݷSw(����.���$��t�0�~��V����f(�:H��(��vqt��8y~�a�R���e��l�M-<	9G��0�
��8�o��\C��u��"e)�y��S���|pi�y�q6�ܫ��<���홗��%�Q�J XTN 8�3�e#��*�eӟO��Ⱦz�#��4��2�LEw�*�37��ux}tn�����h����!R5�Hx���`�-sё�ڿB�{C��T����n7��������%�8Ag�D#<bI���4ٕ/λ(��P�.�>Y��M�͡������[�Hp*:u�<�ؚGP���%m:9�2荙�	R<�?t�xuP��;��{FM�]uvFy���K���P<��Y�V���A+Aĭ��[���;� aJ���#pV��W]>���N�a&��\gmu�]�V"��S�C�r�w]Ѭ��+c�U���R�0�S�0{�I�wA�ћ��  �:�mN$�fo���(�����M�Ax�8�ر
2!L�8fpW}�[�����֎)����k�rY�|�*QVF��w���>�XmT�,�ɣm��灝��Fa��)��*�����J�7����!�^ �����{n+�Zh.���'w�>>rPܨ:t)3����.�Ȓk!���q<���{
�>�@j�{hՎ�`ݜ�f.�`��ʟ`�p�X�\�>4�d�{8��F���㵕qQ��l�N�>r,$+�nW��:ՄT=wh����ṅx�н��nFCeF[�d.sQ�s^}��r�Ler=�����jq^��dMf����,��&�
"�4�aQ�����U�/�v(��"�K�%Y��f���X�@w������~�x�7� 4cK���Y5�S̾w^q��nO��B�b���U˘(!Y}Wy,j���VC�`'a��S�\�	�ו����\C/�9L����ce�U��S������s<,�(���l�;FT@�E�mW]3��R��r*&�;q�aʋ~�4 �C�j����%����e�U��D5Jv2f���ۮ����=�^9��qx�b�_v�ͳ�wt��C�l�ycY��w݄0#+:v7x���t�K8��jw��1Ϭ���2m4eݼU�(�8���V6R��L�Z�	�%״r�	�k��B��4�[��mkf�l�λJ�1��;�y�����rP�θeS�qW\�e�L��(������S����WU�>4eΓ�;]j�(v�쩋tm������7�E��XÏ��9��S�Z�χ,�ʳIC���LՉ�k�m���dN88��v.�숽���.r9>�]�l�6���('r��WI��_p�+;K��j"
ķ�v���7�۽���r�����7��Ȳ���q��%y���K�-I�f�2f�7��KY}�"uvC��y.\2i;�yvH�n�Սx�����b;O�������t+b�E��o�wj֩����G�����c�����ʲ�������u��w�=k�V��¾������� /#�u��k��z�d��Ě�i�7�*�����a��6R��mρf>�\J�WG���}�xZC���[w��ᄻ���z�u����j�{`~|���Z�@f��{��%��U�c�e���aq;1)��.͍v^G�K�<��|(e'/�
Fg<���� ����/v��0�J�<�8�L�e�D�wQ�|����v9c�s��ͅMKV����`��n��9jgf��JY��'�i������l�}�H��s)G:�m^ 2�p׺�t�u�u�w�s�#uw�c�Y`v��b��`��`����I.������^^�ת&�:�;<�- ���q���R}�N�&Il�D[O.�Z��.De�.VjȬ&a 5��=�_Xs�f�r�L�
ֵP���߁�t:���"jٻ��m��ff乢��j��Clj��a��Y]��a�q���a����z�,nG�n���:)�p����X�����[�Y��#u�hUҙ����M�!��9��7\Z��v��d�+	b��7�]0� .Ņ�E�i�a+[�{���Ee������wZx�՝���	�]a�Q9�۱�O.������S���Ρtnֆ7��YM� �MN�J�n��2��`���uݙ�6�A�Y��T|T���e�:�3�8�B���۠��vM8�C����L�FMd�aS#O5S����M��n�����ɨ�tޔ���K{A�lu,���~{�ͩ�����j�P����R���QyM��1�4t�dk3:0�:��AL��}�y�d3�T79��vYI�v+�v(�iw�#s�%o�Gj������ݮ�`鮷@�g&���}�<ۜ�޻�Co:�E����W�d��d)S;&I4K.���l�II�\�U���M9b��"�9�F7ݴ��\�E�uFf�1���&$��\݈�w]����ͅ�w:	�뉅��v�I9�4��u���C3 �M�s�D�]�4)9u%�ؘ��4�"9�2E
#f�tr���1�����)s��1$��1s�� )�H�P`�w].r�3ws�	�
d����b$	H���7X�':�3fr�L)3��D����!���"���c�t!΂"l�t��H$�����)�`��"	�Eݐ��d(�;�Ā�wWF�
 X�pɗ7I�w.F$%d�\�N����q�hU� û����'73��]d�ˈ�0���$�ݻ��v�!���
3���bF9�HS2�5Ҕu\�]ݲU�wwt\�g��P��RFP&����u��ۛ��x���L|@ (���{�l���3r���%r��H�i�Hש;F�Eъ���k�X�Y7����VJ�w��36�OXެ�fWdr�����k�����l��_�rf�!��V]K���3��'�R��;#�����ïV��ǵ晻�q�VB��4F�cۑ�pׂ�A]P��c���\�xL�o�X�BV�N�N���yQ�T1xՊ�Jv:,t��y`�{ب��\�$y= ?xUjǏ����n%�"�|$��3��^|��[�^�N�0��l�����C7 ���:s�|߁�>��^q�
���=+����)��f��[�~	��-��%�����[�n;���Qέ�C�hqE*ޔ5�kʼp��53Wa�.ta۞��+Úvh��ܗYy{=���p��he)xd�Y=^��h�D� ʫ|�����l�p'a��9WL~d��=هU��ڨz\B��'. �f���x�/�^']U��?��b�^���W@Wg��T��u����Yv|'��@�����"���Ș�k�����|a�uњ��_ubMIz����|ҭ"�)L�ҧ�a꙰�4ls�?]`��*":��l�4m!�����Z�\�Q�,��"J�f�w'��K<4�Cv��֚T�)��{bT�=f�B!���X��@���Nԥ�>���N�N��<FF�/b��EA5�#�՗\�$�_�]Keq�^�µ��9��Ё�X�=x{��k�)�+���ʻ�����b���i���?Ӑ�&t詞d��; M�V*�e��*k�{���10�y��C�a5���|�eqxM�bg�>��ڧgc 4�� 츅zh8�S̸8�l���UN�r@�d3�=�����e֟|�A[H]
�]������4|)��8���S߮�#���}�)N�=9k���r=��t>�\F�ʔlYd�3 �R�Y��bC�oX{�u��}�S��uF�(��{�Hq�1�B�N�����p�x��*�|B
�2�jb9NY��̟��gڏf���_l��T���22_��{5��������Z��������w2�FǪ9O�L��Z�WZ�?~�W��b�e�q�\��33�;B�◆�g_$^���I��F�+��(���-ע��e@�!F�]S��`����# T���q� }qn�1N��yT��)��ğ!���O>��ʃ��#.=���(<���	��س2��y}�x�/�w��x)R&�J'A#�=dhv������P��9���f�DB�����ٳ����thn�]X��͹�T5���ϲ:�>���޺�f
8x����3K�V2��5 �.wi>��ɵ7j�֋H���{��#�{v�4ֿb��-�{�'ک���bw�q�3W��*(�������L<a�/�������IΗ'���#EMK��\Ox��@T����<N0P�2����Py���`�@�c���O�������=�Utl�bPn\F������$t�z��i�>���
��~n�OA2'1��2=�+����]0Ⴑ��s��uPc�]͇Xz�Y��7�x��iW�w+.op�b������w֌;����oӳ+�E�sṷj�O*���3kS�5t���i��CPpx��kG��ՎFѪ:|L��J#q�uJÁs�3Y��yR�X�/}�MȪj��yk����pυ{O
� <* �*�j���s�����_+�[�l��Y�lm^[Xd<O��
��\�x4[�6�Mo���H,9��w+j�[�7�[&([�nyܸ�va����c.���23�a�OI����	�O�[R6O�s:�]��qt��8yx�6C�^����5ԑ΀���k�}yP��U��&�r���uL��Aeü�O��=��������sM�������vv�b���0Nڽ��U������p{_��D���x1u�u瘝֩4�N�	v���Fֳ�8���9��Ɖ��Ֆ�Rum	A�U��oX=B��^��p�}����氌���{| ��ak&g`hK���M��,_ft�r��x t�ɸ�w���� �4��Q �":y��2���UZ�n�4h�_j�]�
H�!{����T���#�?g�A�pz*J4�@�12B�o^d�cu}��y�e�[�D��8�:,s3��y��sѸ�wa�:n%�(�� w?��iR�=f=U��J��h�YMM�^b��U<6�(D\?$ը��
�N��[a�4Adu>HƓ�g֮r>� ���Fx��G��$T���@|��ZT�	��-ĸ���B���W"�j�~�m��:/)��O1��f�VY��b���Q��ޕ��O�ͩ�S&���#� ����f���ո�{�z:d�|�q�ͬ�p��[g�o�8�!i]WAjN��O��(V�]w���2��gX>�� �1����Y�D��^!�ȡ֫I��P����_P��t��OEN8ˣ����eu�~�u����k*⢹�N��N��A�!_�C�@� �̚b�{(Ut��:�8u�TD?f:-�gQ��Ys���u��Sѡ%j�s%]e��?���|��	����s���tWԵ�m��+�y36q���hC�^Cߒ���x1��ə�g7G�-������|R���.��tͫ��GvR���d������m��%�׽/�-v�5����.s6�>�[*s�h{��L+x6;�n��rD��� ���I�[��k���e�+ �"/�w1�\�ɷ>ų~櫠X띊��E
(�[�!�+�'�Il�]����,�i�Q�� $cK���Y5�y����5�nۡ��ז9�;n��y�c�=Rr���D��TL�;��S��`��ϹF�pl��^	�e.]�nqo��lqy}>��g�
>+ă���>��7���ݵ�tUQ:�8�o��Lc��Ł�侵�6�c;��j���g��x�OQ�"w��J�����yp���E{Rm���V���J���YM�\��#��J��B#ŏ��p�	�^���h!���ʱs������k�~��tC�zo{�F�+ب�u��'�N��8аx�sK�k,G��{P��7�X?!���}��^[�^�rt��9�����~m�yX��x8��7ٸg^gtn"zQx����s���ɝ���nX��=�~	��4�c:������Y���"`2�$,P��)Wz}��a��^\(�#w�i\��Nz*H�p�w�::\�/g�ϼ�hs����=�nj�4�;�Xc���;���i���Ձ�̓���(#6S��4�CX�da�*�V5��T��\;R��\�^m&�2���l���o��d�:�V���4�����wU�ot��m�X�y`¹�?{����[坵�c���G� kq"�l�2OB'�FO���"�+�d^R����(�%��alP��5,ʝ�,��t=�wQa��i�q��9�yS�Y<0���}R�0�K����u�e)�����g(���ذ0�9U8��k�и:\5�L
�n9�q���[�8�o{71�Н:�6*dd�:[7�j�dz�m:�F�����/c� ��E�^}Ӻ2�~�}Pp��*�x��wYU��S-��/���Us,�E���]_m��c�"T��-F��=pև[�ٸ����_k�����r�9.!^�S̸&����cVUt����������t��PR���������G�+>�g1Ǭg�����kX/3y����C�
��g�������dK�C@V#�x���������ܜ�hWot���>��UE���bC��u�ӿ=6��p�x�"JF}S�X����fw����ڂ�P냳U�,�S������a���!a���cmUyPh�	W]:���b�9�}�1�Z����ϯ���Ȇ;�y/9\�8��#�2�'���Q���"z�+M���]kI�;���J�s��%��k�c�Sz�T��Uo�{׮*3���,݄t��v��5I�Ѱl>��s*}�L|{��������k�����h����k|z_83M��Jr�\w�q�s��@��`���Y�}�����ubB�TZ3D���].�L�^�L�T�x�ޮ��)�d` ��<�=p�q�bmt:vsR��W�+�o��=�U��C	����ˇa�G�.ɗ�lt,�V��e��q��/9�>N'�x��s�I��r����[f�#�Ⱥqv�m!��[��h��Y7�UoF1�����9�d�fX�EX��Zx��a���b�m�4�2j�O4���E�܅7�a��.{n06�����8�7.#K�#�q~���Ϧx	g��w��L*hgǦx��hl'�u�gK��������:���������u���� ̂�b=j��Oׇp/0�\+E`�Q��`���^�����9��L��~��C�/��s+h�NL�O��g�=�Ǳ%X��l�t9�d�+��>��,���Q����5;Rʳĳ#��y�]u�{���f�{Z�M_�XxP\8W��n'd.@x9��Oz���aӨ�Eis���o����5�������5ʺ_��}�v�����w���mʬ�����0ec��V�mt����%(�1:�E}�\���ѝ���]J���5:h��|VnTgE>�p��+�Y:#lnwA��	n*�������T�lK�������ӿC�l�
U�Ҭ�?�[�8q�uޭ�Id��Xt*���.���5"��} �Y���������+|���Q��r4.T\I�$�%W1r7:�X¬���3��R���U�Y��Ӟ��,c��T�ɇ]ɱi�<tm���l�.f�
�h6	U3��;�D8��Af�qQ:�=;�C��p}��D�P_���M;�.l�<L���� pTOZw�]a]���UZ�;u���ț�j�U���&�{�l�-H��ƞ�g׮B��EIG��<��k���-�,��Eq/5x�H��5]!\�嬍�:���;�q���<�؝6"Y􀈄dq�H$\�;�Ϟ7�<x]gS|b:g�ʖ׮m/�X�ȮMZ�nQ!y�p��6�b-�0/¢�w(��+񋘜�h�����N��7�)����)���%5:{�������p��u��������b�ss����a���[9��4v��J�i>�6�Lr�L�6n�9��#k�η=q�[�D��[#� y�W+Ez�5s��71�y杤M��L�{P����謧�:jtU���S.�lނ�"�3'j���g}���<���G�PY�8XKUL\_[<1c�
��,Un��޻:�����܇����.�(���mN���w��_}U_<��+tܗw]���Fg�q�r\
�
�{�Vӊ�^XXN7)��e{�Zs��|q��<fK��D�!�tw3�9](R�
�
���`Q��οp7��0�#�=�H7/��EJ�=��,}^;YW9�N�Nf���Bʐ���wXk(W'��d���VF����[����:��	�2,s��Ӄv}>�j�s%]e�&l�B�ճk�������9~<EÙ����Hq7�<��U�+���S}�EO�,b�je�� ���3��Y$�����+zV�H�ې6v\(�Y<������`�#u�ط�kټ��]�;(�e�����I�%ïD��ڙu#Er�$PZ���]86��<���:��&�d\�DV�/8?ol�<7�.��� |+���?�Ks���V�?x�E�:�q�՘��t{�)�\B;A5a�xͲ��+O�:��;�Hi5�{�z�_yY�Y��%��	�췎*,J��yM���0�#��*T��F�x>�d(��V�Y�M1�*׌S�/jP��el�L6{z�s�Ύ�z+ k���+�j�#uK���S��[A��^T��SZ��V� ����"Vޝ� ���;���+��Q���jQ�ʅ�|��n�W�n�4;,[f�,��|�t�4Z�r�E	N�
��������t�ýR��i>��1����[^���.���N�8�d�uJ&��*T%n�FIo��A�و�}1�Ε�L�+v'�ƀ[�^���Gs�8��7���	8R�G��Py��9��Q�H��$��" �	��BzW��)��c�>�E2:��1&��YQ����e���uG�fW�i���)�31Ad̎vudC��ʎ�/zV�s�{�Bt�u$��f�ǣ7)*����9٣a9]�hel�2M(�}����E�������s��UQl^]�a�UQ��i�q�9��kʘ:Y=�2B�����}�t}����˸�lz�ΰ���d!����2�,sְ�\4Ș�S0/
'+v=���	�la�ڒ�<�&�h���)�$��q�:S7�j���g�u��,~�؂f*�&���r֣�7ְ4����Gm�4�ģ��|��U\�$LZ9�v�s�垫Nj^�Ƿ7�y8�@VFErp剕	�^�;;iT58v\B�4 ��GV:�����=�'n��2�*���ժ%h�\�9����:�ڻ��m�R
����=�g[L�47�k�&ڼ ��Z���ԡ�F�cӺ�4�k��f>��ɻW��+����;U��-�y>.�*+�N!6?�_jצ���b&q�݀s'
PšI��{6�ɨ�L���u�{9@%�iG�Bi6��^Վ��t�=�p�oNQ����m��k��ެ{B%�x�y�/�I�R�2��I,��2L��0�S�t�)]�������OUY�g�.��gޑ�0�z2�Ĵ�[1܊�T��f�#|��������x��;��*_B��s�N���y�,ow����H�dwTI�Q�3i�d��fV}�%l�5��c:�%���\�:�{��н��������m��`A�e����0��->K�T�b�P�H��ۼB�+$|5#,V,�ٍ�xe�L����i,R���ax:��ے�N���vv�VܭM�sK�;EXtư�m�;�qb��'e��=K�ް�7%n��k`��B��������n���V�;2��M_X�ֵ�`!���X���6�ȓ�r��������[�i��ؽ�S�Ln���.<��R����[��C$�6�R�����_tޏ��Xc���s�3����b��^I���s�+��
�M��)۵��z��GӔL ��6Ka�;�ue�[ 6�L��*�E�6RJGt�7Wc5��T.q��vr�0�8)է1LZ�o09�l������5Z��FM_<}[>�5ϡ58��f�,�jf�A��&��F��k�6L˥�l�J'�J�-�t���H��p�僨ס+U��*�z��w�q.3)�y�'/!�UrZ7fRڨ^R9�<	Æ/���3#�+�κ��A��w���{]�%Nۂ�BP5i�@h�뵝5:��.,��,���K;VЎ�@�]>̈��7F���<��/2<Xi�i1'GG{�[5>uoi3�����7�ћɩc���b�.�1�i�N����*!v�B��wM���EZt[I��u#8ü��c7s�]�0���7��q�B.���\_t�n�h}<��Lu";SXE��<�ɍv��4i�I�J���)����m@r�+`��gl�c\]J$�M��Z��9i5o��՝��\�usy��щ������mX��FS`�Em�z��V�M�ެ��GH<�dި�f��'�o��`99l3BxGpU��eK'	�Tn>�2��y�Wd�D y ��Ž����lm=����{5Wܧ+��W[�:����IG'��1�A��G+h�˕�o-�:��up�9eЇ�+�ӼI����Su��ՈE�)�frm��.���P�ݰ0L�+<�80X�.�YGs��Q�+��;� }H��-�ss�Q�U��L��?
�(&3b"H�d�$�����q�a�.n�;���t��(RdLQ�t��9�y;) 
R��R&����'v�jdB��1��*�H�L�a��q7��H���)�	]�59�"`�7wQ��i\�s��r�1�N�R��$s��q/�6d I�:.��:]�d�H���� DbYr�.��I4���wt�F�3��F:)	���Bd�u<�K��vn0�D)A"I"K�a����;�Is�n���9�%)H,r��d!�] ����9˴���%�t�"	�F�,u�)Hd�Ͳ���#Lf]�W70f9�d����f5�uwpbDwnbd@I1F�nAN\Ȥ�Bb[�ƍ��@���t�ι4BL�4�XK�А�9$Û���H;���nQ(�Ww]��WWam���r.*�����}�w��k�94�2I��'�
���;�b�t�0�|mdu�L�����w��p,����U}U�U�>�w�'�����VG�;t^���4�~�^�+��p�O�g�9�<
���e�B-��b�(��Ɨ^��l:p/��g����P�t9�Wt���bg_�R��[�;}�0�U��]�:�wpqn�3X�����w���X6�:tq'�wX�p�w�B�4��s[>��F�ˮe���f�S�� R����F[��³fc����S<s1��Z�;�t�6��똈Γ�P��zU�4�t�Jq/�>.C�Ӊ�@��(��f�٥8�+׾��/P�}i�N� E/��Ӯ�2J�2��3Of�ơ)�dU_1}v�w_F��U��vtۚ�=Ń�2&�NXm����r��1��jbS�u���׭8Hob�pfۚ�c��mG����C�-�,��Jq>*C��#���P�~���H2�p����z{~�d^���J��,C�W5L��ˁ�@T�Έ����
�mΉY�^�C��'��JJ�L�'U-;D8���
.{nSTTc1(7.#K�v�,C��؂�Juߦ�ޫLYZrd:�5��=d�/,ֆe�R���T��j�ݨ���Y�)�v��F��IȜ�靷}z�¯�ny字�i�k��$��=��ܥՎ����|�&V��̶7�Fʮ�8XsM��Q�ݒ�k9%��J�5K/���=�Enb7�9�6M������;��:��{���e�uN�,v���X`���O�=�wԯ0���0z�bW>�^�Q���k�1xK�c�'D��=��^C�G,b<ǽ剤u�	��j<��؞���kȋ�f��FP!CUBՎ�[?:�->&�n>U�7���HR]Kz-��7:6ꮰ�c��{pn޼�N�ma�\h�UpB�����V�
�l�ZKt�op�n�$3�"��N��.�w���{��/���b\J�Q����6A�C�X3�v���z*MV��k#��z�Ɋ�<��������/��ط��2� ��P��Z5۴���
�Y'K���FU{d�'=

4�]�����4����;�n�8ۚ��y�����;!ܽ�X V|ð�λ��+�]R!�y\�ˇ�ԭ��sz�ܛ���@���Ť���όf��Q3�@`:]m< �[��Wq�b��qۯJ�Z�a4o6�m4^wq�UF�Cn�H�9�=g�Pr@EIE�7]2��a!�%���n�����&;wM����ab�[&�uA#���y0l��-�A��u��Q����	y���ĳ��[3�n��T�x2��V��`�_Zp!s���m9���,�Y�oSs��L��j������a}�B�j8��܀��b�f�"fL��uLF������<�zgq'��L�
�=�W��;�q��wo]��q,�Q��1	��&���t�Oe�9�X�6�:�u����ը��"E�E�%�9���Y�%
u��7y��+is���e��8�Ѱ:�Ճ���y�~J��I��/4�#b�
2 n^����m����^�\O��Y��{9��s;Gx�<}~mH�Vy�E�����u���'9�����ڧ]��a�v��L�zh�qP�T�PKm�f�s4�v󷖺�5��z���K:!^�>�G���x�c0U��!uČ�@��"��U����L�k9������9-�}�s��9>��a	���ʬ<Nd+�P�5Ջ�kў<GzM��]F;���J�<4��@	�-Pqh�:�瓮d_9��9�>�n�b�t���ru���aJ����v�)����dd`3̞Ȑ�"�'s�l�}�f�5]��G���]n;wM��זf�(�;~��4ghu����� 4{�e²Yd�)�_;�8� 9���qÕ�l�v/����8C��q:,U�����=L�u<$��b�i�z۔�j���3j�\��4o<<�S�b澕Nas2ۊu(�e	+{�X���;H:��bNw<Z�zn�F9���H!��__Bd��]����σ��eGU��_xx{�k����"�족zjM���4��,+#~j��`�u��������6x���Ӓ�c���������CS
ӂ��ă���pu��~
�[�3�^8��l/B�S_�-��y��zƠ�F`.!����<f�`u��< �:�Չ=�wUM��L���� �8��h�Y��o�m���*>��V׮��_��["I�]K��Ek�U�0*��5��{�����-����|w|�tq6�1�R���2�

�j�<��}�]T�R��"0�c�Z��cL�/tD�x�����E9�~*���|7n#�B��X������}j�Z�=�#��@Wx訵v��RdoA�i�/E�Ո*��m[���c=w���z�)���^ �NI0�J���ՑR�8��,��"��i�m�y�IUm���.ɓg�d�N���#C+�/E{�'��nAvE+�du���ۇe��챮�֧z��4�C�}U�wuqf�ܸ�hs��k��9��u�-Wm��-��<�y��[CӴ��C��kb{�ΩS�k��Ҧ�We�"9�fERf��t템�g���qo�s2���z�Y�KAJ����m)����V�5�5�k�Y`qo���Ԗf�/-�=��B�[����]�K=�ul)�U�L/mL��{��}�}U�z�|��Ex��>�Y�r]z)��F���UN�k�f� t.�dLk��ɳY���9�{��#��@Xw 4ژ��&�WJ��L�ه֯0y�b�S��K�};:����f��z{�oG���j�6i�Џ��g���[��8��VyUs,�c�2��0��r\�Yj�Ǚ�1�_��sM@vFEs�f�\-���Xߡ��{��^�g��<R�m���.�*yfҺ�X�u�n{��zk3��P0a�\+�����<)�\ ���3N����r���ߴ�*aע([��g]N��f����@���q�F����w�������\��S�.ϝ*Wp{�w��X��,c����>����Dt��;�s�kz8�N�b�so�*�D�`ρ�n��m�2�U�,�Og�J��0��s��{�1�V��+�r�8�=ǧp쮫��W��oHyb>U�X+���|��7]=ҙ.;��8�;���C�^T�y�y��1�(�n���XsL�3�:T{�����_Æi�͝;�z��m$�vY���z'Ebj^��m��c�"%�.�x¼�n��E�桺�P��`������*��uT���qvv-X�d���ʖƮ�]�;{]P��vh��;6��j;jђH��f���b��F��]�;�Cf��\J�=�/�x{յ�[��[��gl��M���"�hmМ�T��)���k�D$wژ�y׆W/<5Θ��jz�s�r������Mu�Q�����bq=>��r�Jj�q�J��-�V��W��lC��{fF+K�����/�p���ԲZf\F��"$'@��qD�G.��QH�Mc�Σ,²�ܠuN�ѷ!����=�ګ�q��8�7.#O��8�`��ǹ^���</����y�m����{[^t��)_��ruXys��JTR�(sU�گ���Yv>��r	��+��V�F.>���P�@ _I��~���Kq�Y��yn��6Z���C�uȭj�OX��4"�٭(��
�2r�S�}^����%`Z�Լ���Z�.��]��T�8N#�����-��"#2Q`@|xR�z(���~�z��Y��流�È�|�31�
ӿE����*��Vv77*t�"Z�t��伜��qڭUok}0��
�TT��k���G;���dų�λ�\��q�9^�31���,���M���o{����.�?����Vp=�7�69��x���V��ہ�th4�`���4��_�pʌ�ؒ:�(���pn��Bv��̸I��v�f3��j�9���5��b�r��F�m); �L�O.����X�`L��P���~���xY׻r��;�*c~��K4��U�ڐ�Ѝ�U�Y��Ӛ|����w��I��e�SW�"��Tkt�JZ<	9ip
���M����יqQ:�='$�Z-5�V�ZY���a�)�>q�u���7�xp1"85o���w�����+Ёole��
�5e�v�߲�	f��~=��=��!3�d(b��\GuF��5-���.�gt���K�Y=}��k��[�Y�q�ý��:�%�8x�}(�G�N.�[n���E�5�B���OyK���FP���5��Soy�5�-�d6W��'�-E�wC�m[�T#�lޏ>N�(�	s�	��~e�c:p]Nx��<��J)U�b���1�enMz�˜�t��{�33�<�fm��5w��Eݮ�b����V�1>�-n�	�Ŝ����CM\�'I���~K|�!M�Wٝ8��մ#[��xn��LZ����(��eD1�<��Y�T�p��Q�W9�Q\)���Kh0�s��V:T)�@F�\�h�;�0����ޔ�_R��aҥ1�\���>�CDz7�ਓ�`ھ�#������m�:�ڑUhp<�W;�_!��'��]ݹ��w����Rr{:�(�џ{9;ٷ��퀵�k�;C.fx���+���X�y=��*�\��!i�ݡ%�e��'�-�aL�G��f���> ���> Vz�]����O9e�s�\�nr���F!"�&mW7�X���2z�
}ʍ9��]k��b��W�B�.��˙�m ՏF������1l��{Ӌ�{`k��^����!g�ڪ<�j��.juU宖7�#�!.�7O��+�ω�~������{���"g]�C�_�<<�F=�՞��ƀ�&�=�+����Lz���������4��5QQ��#�C'h�`�(��nWN��ZsN��5�]y�ل������(��ݷ��n��B����V��}2�h�qZy��Bޠ��׋}����'��"�e�1�y�T��
�$.Gxz����3���e��U�E�\�W���TfX�/���p��؎D/��?c���k��
���Сla�+/�4�@�i$�æ�*�/���	-�&��ʷ(�K�u�����'O��Q��9�\��V,
�&1��h�ұ���+m����[������Sc%W��;{�=��E��uk�<��EZ����\
Aۡޙ���r���-�g=^ɝ��3nƧ��c-��/}}��>�
�8�o@���g�����굙��hO�rw9���^8��M{�q4lk�p/�=�	�Ǣ;���b������N�Z��5�cu�yub��M�9����p{^�l ���w�uOm*G3i��u/3���׈^�;�/l-a�_����w/w um��/��q�)��LZ����{6�����O�+�����}�l�㙅�{��NN�=�����h��Fe ]��`��1�Gh�B|/�y���"°�WΞní�3���u��I�h2z���,9�}���W���oDx�R��=�.��j��7[�
�t�q�Yw��hqʰ� <��v�M�B|�9y�4��9�����qV�ya6�ľ{f�Gm��QÆM�����az�)�ZC�ix�k�Y�s�gMuj"�S�����Y�ܯd�Z�Ӂuj�w��E�d8V�2�K ��0�X�+ �[ɛg��]�6�EӜ�Ni�B1��P�v�ͤ.�擾�x�D퉠p�d֞�g5\���P�\��u���UU�Uz�]V��n������.]��JT���X���0�~��f�>;[©Z�W^�yY��P
���;��RKԪ ���I�0�!�-B�=m�9k�%c5N�PR�������=�r;����ޅ��)n�P����Պf��q�l�$��A�9NQ��#�&U]�;w����z$���(�xl�d�\�.�/�0!޵��"�geD-����'�Qm���s�����Ɲ��ލ�Ϛ�o��6�8��R=�z��Y��g)�T;���9ܦ	��-\��6�gy��c��:0%[��v��!ߦ���Z�q¯}c�n�4����[@.z��J��m�q1U#��E��^��j�����}�$q�"�����[�����xc��u�Ԕ�.�0��%Ѹ�t)ǝq��Uxn��-v��X|�s��o��R�����.\��CQ���On�.#םINwǀ�bY�#w��`�	r���Z%��wД-!-U�$�8�'R� ��u��'�^��y0	\�����挘 ��ڻV�oLnj�ź0��I˚��j��(���{DE5�q.�|��1q^o8�u�e;�Oz����t��O.�k�Uok/Z�.���Kc�s�"[�{!˙��H���@�x�Ul��chŸ�u��m��:2_n�U��4�a�5��J�-�p�֬��ɉ�@ǥ���r"邖
 mnbFM����iv��mU����m8';cF/t�,�:"� 9\��>K6�pL�\8鴣7��{�,� E�90���
Vk		�O�hFڔ6	s7Y�,Jh�����Z9��-J�A-`���؆��U@Iw�`���ҳ�_.�x��8f�ܮQ�JD�tba��ι49S��n�4�e��w���Pϳ)ݱR�Z��vԬ)��N!
�V�iv'R�>7�:���i�����G�3/����LK|��X�殐N)ҭm7�r>c�.�l+�4��\�.�u�GJ�k=QskC�^��ε���s�mRcM�T�bsDٻg:�����JP�de@d*�-݁!]$(vm���,���6˳�53��b�7�o�����1���j��ő�gg-ݑ�1[O�lN�XL���9r�<�	�5}������e�"��PWO��6&�O�ɜ	�&��&f�)
�۠�YWu
[:�N����{�������n��CVsSsh��fY�Z���,���o�n%����W��W�iʹ��wg�<�mn��C+�os<�,�e��|E�4{�M�=[}H���Jܸ3�s�#�ا� �w���7n;��@��zrm��I��侶兝�c�k@2�pu�{��.j!��8㬕y��
,��a[��-E-]��u��1��:e\��9ƻzѕ���c;X2	��d,����gNt��#|�\���`wC���������� �6��j��
�ZN.���E�ɩ��k���_�}���ކ�,�{6��Z���z���v�f&1�WN,B�%���n;���.є)	���I�<\��f�τ�3�f��A���#o����n�:��"�:����]��U��*��f_-�20�!xh>a��kۭ���Y�y� p�Cy��Պ���64�]�u4Vi}�:�X��8��駴�5�5�Š�;*�&��+��B*�o��2_T�rp]����[1�͞�C�e�ձ�a�z�E{�j������bx	�����M�����:��(�tc�޺�˻����EA�aY�Բ�8(u��;*��&f�+8Y2�('��
ڽЮ��lAX]�[aEK~+�2�u��(����_`�u��tA�2��R�e�v z�Ų�+;��	
f�n8ﲃN���ݻO��AI��@��u6��%��q� �����]0�N������5͙r�	)�ELc��)�+�(P4 �4lDW9�r����	��!$TQ%�Mv�2;��& �ݺ%7w�,;�D�9tJ6$Ɋ)(�c��ΤI�r�$�1,�dI���ܘ�2�c�(�r$MO;�!���1�Ƽ�0�����I��M$���fh�d(�6�$a#H���,!�H�ӝ���0�wqE@�i���)h��b�,�4b�!��&���n� a��b)ݹ$P�tk�"0E�B9�B��$b.�d�hK��Ĕ�"��p�\�.�9���� ����Q�Le�n)DF!2�wvIRI�2�u�X�Q�A!���7*u������I3J77,V""�WWUQot��G��Z�=_uy������5���Gx��x/i������c2��s7gdu^�R;K��)]���=���U�|�)�,F{�N/꥙���Sܫ�C�VOv�ZW�V�ma�
��V��'jǓ�ﳸ�=�H;Ժ����W��5�kl����ZW�'9�]��W��T�a�sӔ$�����$ͪ��ǝ7�%v���r��)BP�_T������:�m:���	X�t�qB�7����{J{5쭌��.�tWs=e���� �*�Թ�:�*Z�l7}�7�)7H���,l����^K�+Z�'xLw{�F�@�|�mJO�.�:�}1Ǻ����T�mӞ�s5��.ǌsگ)���������O�wY@���=����y��[��ovoý�r�v{X͠3��B*�����3��(d{���L�8�	~��W�o?FG��j��Ov)�9NY�#b6�9\��ɪ�9K��[��u9�'_-
�yoFW�4�}v��x#Jd�������]=��xL�٬u
��sy���n�ѡ8X9�B���:�|nM��;&��yy�)�A�v��㡡M�K��CWx�񤷔<[�@�2�)�� 17u�֫W$�&�D�@ۃ���
�㗋p��v18��Q�7��P�7�m���K�=�������ɣ�ʯAJ�`��h��67���1.s�7��A�R2�o=�ns\ogZ�W�Ү:�U���u�[�B���ym.z��g�hOr�ɔ��N��^�8�M�v�V�1�7�_=�ڬ�mR�~���s=��hS���]n�Zs�R�@7�Z��{����]�P��)V�|{�X��o�����F��N��c�R���9�}Gk�s΋�|.���q���ǙR9�M�.:�M��I쌼�$e��)���|�9I�N�/�ܧ&$3x�]ѝ�Ţd�a�4l�q���_$ͅ\�[�[�I��;�"��TC���k�|����Y�W�\�;մ�ki�5�^��Uk���v{ދ��y�~jy`|���Y�ߌ�,�9��kɬ�]Z;'=M�3v�����)S��z�o/�4�姷�/*2&���Ͼ��`^���ə�@�ƍvJ�9T����y��]$��s:z���)]�f:k.Eյj}7Un%WcPf���� sİ�('�#�N8���7v��}�>�|��:���M���.��Iαیi����"��}�o@��)��њ�w�kV/?���������V��=7����u5����5����c4И��GTq�\�^3�/��6�/����
��wƤ��u�Of�O,sƻ��O8�)J��s�FZ�(�T��9f�� �����[�寧h{���j���_8��Ӳ��':%�=���b�O����}��<���9kjw���$m��.2pç!�n�ލ̊M�;eD.��؄�nyv�)�����W9�hv��Q�n%4}�8|�	T��r���겵�Rr:z�ݕ�7�o���nvO�PIlF�B7��������O(�kp�x��:6����S�XR�Z�ln��Պ�N����4���yU�R��3z;bq�̘��*��(]ſE���BVe�����^�;�-������}��N�#y;��Z�?S�7R�u�ٺ�&/��F�W��N��'je�3(���c0A��~���%_R�@�*�,���wi{0k�\��,�3%��@���TY�u�Fo`�ʯ:uh�P�޸�)���R�R�6�O���me��Y}�������I��]�W.�yg �N��Mk�8�5z���{��Y���ip��]{pi���|c��D?_?�V��6�ќny�BΫ|z�KQ�����W������O�[�����U�{�^˨��SG'x�۴��i�0��[�\�/M퀫�Uv��9B�>�U�z뼻�|U;�xsvN˝A��t�an*�o/ɷ����}�g�(z^���1ر���WQ���=��h벨*T�{�ycn��^쟹r�*�,�5}r���b5�[fX�T\��t�>U�),�P�:{4Ryc�k[7��[��x�s1�n��ù��̟z`�}޷}�)v�~���jB�[ո��b���U[�FZ���m<gG�>��q	lo���鳣eK�IU�1=�s�����s4;�Ư�Z�5�r�� #�K#cf��f�]�z�j���;/ӽ�s̷A�F׹�A���f�+�8'�R=��Qr�>�U�4߭3�Egk�( �郅�98njL���~��^�˕��vћ���r��<��3�07��f�3v�~����������srɽ���-�8��sJ���x�і���[�j��F�j�q�]plϜr������S�[)�'a_�2��O��o'O�:�}SC�p�2�5 B=Mt��F�i��9�a:/e�UXoj���H���Ặ�=w��J���R�.iƾ��E\��e-�'��w���Vy�Z3k<���输�x`ʿn�9��Ό�%���aO^;�n�<7C\t�-u�F������M{�K���Sa��yҹ+o��N��'_Y*�
&ov��AwZ�i�����і���πS<�c�]c���O>>!oӭ,�iv%��%u�E+J��8�F�d�X�bo�fǕsq~o��U�s'LK!����}5�\,�|�5W���U�SS�%q������o�k�އ��/��g���+��Y���̆��@���u�y:Y�9�.uV}�CQgE7
���p�.�ر����/5�5}�����ƻ�tgԮ�6k���>N����A��v<r\�q��j�����Ʊ��:��,�"�"qڍ��"X�0ԞV�V0���er�	2����:��0>��Yt��m^Β���0tǵ�k2:�}G.<Y˫y��OY�:%�siGw;����꯫e+Eg��R���Ou��{[@<��&:��>����ZS�T-�눃|j�o+�����Z�*}4o���v�T���o������O�p^�)G�SD�p�0idPí�[�_gҸw�s�6�����x?8f�%���4�쏻wD'��[4'W=�X��z3�IC}ǧ�w���+��3�d>���2Szpa������u.��M>Q��������U�����K��߾BR�*��7� {��vZ��إf� ��:�����q��u�ʾ�����lk��Uk�9GH�[B����}6�㗔���'Z��J��c}X�$�o�XsB�����_�g�z*����7}W
k��^D$�/������n�m�K�Z�5���Q�vn6�ƭ�c���}IM�g0
���&��VFg!�m;
e�)��ηCL���u>��=�cr0'ډ�o�CEJwu���eܢ.v�Q(�+MԽ֊�&pO��r�(3[�N�Y���i��G{���8��^o�WN�uwZ�˺]��.J�2S������+U��=��Ȏ.j��s|�.�ep������5(X+��s��^Y���z�*��0�p�8_$��*��ud`��n&���˕�"�z�����z��q�nө���CX@�>�E+�����㝱���~��5��C�g�~1�B�뷔'���{�ʜ�o�H���]�8c}�V�ϊu���⭆��O�Z{~7��g��F�� ���:��%^�tˬw�;d��v]*U457��5����i�K[���1���np��G�f�̀��/�����.����N�sƻ��^y�%��˚�6N�����1ݶ�1SQr;��%�Zy��z���׋}��i�bR�;��Km��t�/�����n��Uq��L8 �6;5 ��'�t�`���r��Y\5n*��q���C̊�ol�#��s�ǽ�������5;�GYJ�Zκ�sJ��ck��M�;f�53����1P;�Cg�7���K�u��}���٭�q����xƣgB�����>}1y[�Xh'b~�I���5��l�e��D,����^�ֹ|±P��kns�벳B\e+r��c�p���3���9¹,E�Ħ�Y]X��n$�T���p�ـ�e��(I�
.���T�"��ڝ����޷�8t�T�4�i65�G���r��4`g�ut1�1��ݝIC�g(>H�-�<#um.�Vu+s�6�ms��ȕY�ŞU��O�����F��=�Lʻ��ɼ�$�Շީ��~���Aܲ��>w�ū���c��~�E�˽*�ޫ\����h��ַ���3�O-'9���v-����Ƨ����S�=d���p!��ݏ7Z��#�sc�u��'�������Hj������a��2n՞��ب�o6�0�8�c�q\���M��Wnھ�^�����Nâ���{��U�������N���+�ⅰ�Zm��|��7��uy"�	��J=űG�r#{�W}�:g�'��1�]�J�+���0�^0���ڣA��]��Q.�٥�y�t�W�+R��U����I�, �B����f3=����:�f�Bba7%��{�1ϡX,G]��s�块J�軄[��^�L��f�uw�)4�ބ�
u��1vEgtuT����Q`z�Z���Ơ:]]�
�`-�U�yՃ>��U攕u�j�`.�(T�":�8���-��(7;����H��y�P�mN櫗�(�{s'ޘ:��z��t]�(U�S6o���g���-܋T�eT�m&>�1�A�9_yq\G*߷Q�'��:�5u*>υ֜>���JR��U�FG{����r����9NY�#�%%-�d܌�����U��,���7�-מ�ms���C�ͨV8'ʑU�;-LbV�ڜ��l���m�k�k��y:����i�p��΃CyޡܡK�wO����������5~89�V�<?7�~����v�<����[��y����g�ωaMn�M��׆$s����e�K�8��T��c�N6�;��$%��$�7�ϟ��׎�h���޸�KxFb�M�����G�/�V�Q��gE+�S�:��y�{Z����fs�u�3(�q�o���P �=�<�: >��Z1�#��]�=�U�}{��i�hY���.�ը�^���_�td�=�sU�9��u����7(I�t�]�_<p=K3�܊`O�:��y@%l&�q�X���Z9�Z�xx��Y��L_k�7aWWV�L�3H}����ծ���u$��bޚxu�M�3���&�[��4��f���z�I���k� �����;����as�&�*GW���gw�c�_gr�Wll��%���ޫS�l^��P�K���u'PK�o!��g�s¸,�y���=�s��!Z�+��m����W�N#dr �sBuT�Q�ok0�gl��;]\��	[��t��5�QQ�9Dl!P�Pڞ�ibY�����u�쨋�T|�\������9m�J�=��P��n2���7�KZS�{��;�l�r�X-�_,k�Xͧ��9J�T+�f�*�竃ž���g(�毡o-}���W�5]��|��|.׻m�x��w���8����e���������Z���5V�C�+oڤ]�{��j�<��EZ�ôd"�P��؅�zWd��(�$��eU�1������K.�X����B�!O�2���Qo�/}B�H��h�}�8`�ʜSf�h.i��o�z#b�$���u�Ƶ��7�^ՠ�3�G[Xm�8�,��u�ֹ����]n!i>��5�I]𧁛�r�ƾj�[�+sy�=��*&[��]��ֽ[�ЭB
9�إ�$E ,�]�9:���	��Q]Fn���m�Y�nҷ �˴�G#�7�(���t7�`���h���(���Zz�i���B������o-6���fi��n��Y��'c	PG�[��,�Z0��^��G�h�tV����W
])Sn.����/l�*�5�#��$�e�!Zv�e����"`��ސ���i���G��p��gt�[W��	��"��7-e�W�9����f����z�Y�RT��8t�� �P��OI.��[7�5J{ƨJux�T��y���?p�c��L�3~��t�Ƥ��ՙ6ŠI*%@j�j.J"v�A�c��)��7>w8Ä���"E��.�óQ��Q�+���Q�I�I�<TodZv��˰��c8��;.�@XY�>Iݖ7+!�chVBT1�
�Y���U�l�F>���GgR��6��)��9�tgP���98�J]�(��@X���u( �-n%d�/��"ė*um�جڽ�)gM�WwP+@����^9Zy�
C�fZ�+��Ȳ��k3�fڻ��G���સ�� �|:�d�\�v�RY��F�R�f�=UՈv�4_a%��k�ki��n��5�ۙ��x)["���`o8�r<�xb�^4(f�"�2�<��װ��ۙA՜�8�(���%k�
,`:��8��!��*��"��Z�u������F����/k�f 6���B�h�S�6�B7.Q��H�qu�!
ǉ%�����l� �T�QHd�s�n�g��@n�t�����'$d���7o1�sv{�̘��F��;we�FP���ʼ�%1aJ��l��'��k��J��d�]E���a�m�'n64n�H3���k|5e�ϵ*���ΙV�M��6,g)��I�.��;��o*+#�w�A��2���o�]�l�����U<.K��ޡ�n��k��O�����7a^8'��S{q�OJA[3�O���y��%��Q��{��\ԧ�Ѽ��Roo�kzvq����{§c{`hFV�״F�����:�K�V�eaY%���6Қ7�%�+v�@�;ܡ�:e�w��ݘ���f'I�7�f�o����q�̝��";�^���i�/��<�Mo���֭��h�Q��es\�`�+Qw\!�2���RVX�V:��,��]�Z�.�Gr����k�&�J�-��b�F���f	�{�;�Lҏ�����u��q��s��8�Hf\��kf,ܮj��%;�6���Ϝs�����z�qW��9n�D�,e���;R0�Rwz��\�wi*T�td����v���U�[ʦi��M�vGx��䯎��"�e3٦�n<�u���� E| ���b
$��VD�Q#�����4c��%�$�L��"M�,A&�`
�r�E`��r�74���(�X� ��JwW]�4m&s��rљ����4E�زLBNtcb�Q�	6!'tt�E$����hрӻ�ȲQ�Q!	i1�Nn34e1�)��,�ѦP�
B�	wr��wX���@E�(L�2��œE%w\�	��nhɹ�1\�G����Db�^vv�K�LΥ�K���s�2I4�d�]��ĔBhJyݘ�M\�HPR�#EId���%Q�r0h���2F�滮3#ǯ����\��A˅��̓��X�xv��EwpmгX��資�}V�3	���q����j��X4 =E:�y)؃�����w�����1���f�]1?u����{E��[�{x��6�f��I��w-��:�9�״��XI�ߖ��m��s^�q�R���wI�K3e�7K��[�u;ٷ����5������ux�w���N㈷�W���]i_��{6����2�����/OW])�ON>�U]j�z��]�q��6��b��������ԏxlԾ��&5��6�]<�Oc�y�P��-mn����Vu��mZ�=��W��s��S|Ӭ|��MF�m�z�R�v��h䨌�j���Ȧ$u��W���g'���9�����ⅰ�Zi�i�{�G��F�ǆ����b5.�kd8��R��QZ�SAs{z�Yc{A4����{���(0�8�~^g,{M۷[W%�wv���٠Ryc�5���TC��S�3�LÅk�|���ރ5$ۭ�DӰ�K]X;m9(�����mh�;�rQ�;/�2���{�z�a�oe���l��4�9���jWki~c�1't��n���5|��CXΠzI�(v�-x0D٠0�B�e*�7�[{,�9�v�j�| �h��;;�X�fj�!U�s�B*���	lW��Y�Bޥ���-�v[�Y�}�N�S�lo[3K���o�r��aO��L8 �(i\��f�Si.D�=S�Sޥ�WB�_r�w��<ȯ6�W�� #�D�Q�|W�k|XQ�b�=�n'ފ�f��Sތ�Ϝד}ٷ�8$*Q<�d<�)���&���_3�,�,˦�ֽ��is�A���iĦ�>�8']����×4Jª��t�p���M�S�[��%ve�����umՊ�N��0����eP#��T���*]��u�|�-������K_w<W����^�p:m�\�X�������b�����iu��3ԗ<>��V��y+ׁ��s�~�������� E~����kk����~�����P�����f5��S�r��6�Aا��'��;S<�c�]i���^ۣ�9�eb����Ǣ]>4t6��^!4�wq�s5m��*͉&�ٞ��F�5��ޕ#�nm�멕�5[9[X�0���ٛ�o��x���N��ݳ�-hŘ�lܚOvM�N:���
f�q=C�� ,��ÙH�Q�s:�V�v�1�[9 W��t=^�V�Q_�nt����)�ll����B�5�ő;��w�<P�}A������`}]���J�ⅰ�&ޗ����vFF������p�k!mk�x=��	�0I+��2�X��1��E�o��{yO,,~�նkz���s��+ϕ�JK*�N��}X��i5��4ip��3X�Z���y�)JBc���JqZRPq!��o7�۾����M S��bb�__(��uo۱��o��=��G��z�י�{��m�Ҹw�w��+��p���^";�8T�Č��<w��dy9�<��{ȷ@=�������P���dDͱ����V��M,��A�^��뚛]�{�����T��7��q����鷫n�W(�������c�ߎUi��<-�ޞ~|`�񞺕����!�y7_�.9���&��Y����v��2�p8��L�{q�J�n��*7kVF�Z����EM�Wj��}��i�h��7 v�ZjtH��s��U�vw�xE�W�*\l�=lh�t	du�n���qa�b���
�Ή����޻ͮ�������zքr�k�9�O��Ќ��K̩ů�h����Ԥq�|�G8WN�����i��u��ǜ5|'k�]�OЇ� |o1mmYݹ�{��O>S/o��>���d�����~>3}��Ckk"8���ܸ�F�dN���N[�jg���]a��~i�~�c�ϸ.����d�z�йT��IA��7��3j���M��i/Th[9Ӆ<qMlU;�VQ�����=���ή�1k��v^�y��g��b��ND>~�gC��d�iDl��DU�.juD�O)�N��x���\�iSS�� �^6��'�kxLw(���>SVr�U<�a�s�m����[�FZ�ۢ�N��Ԟߵ���r�6����� ��NBV2��8a���b;�װ�kg:}0�^������O�r��Q��s�*��6��M��N�`�:�
c�
�t��ɺ}R��p_1�䲔W������Q�غ��KQ:��Ϸ�$�e� 2cӘ]	3zB�J��>jf�����prq,����9��z����=K�g�y��k���̎¾+n�Cg�#����؎a|{^�ZR���߾_)�����fBޥ���iX�z�<��
���4�]:z�)�6�x�B��R#`��f���:�{4\�ywfSK�/�I�����i�wG?F_E ��A�2g�$64�s^�]���MVUe
��&��]����m�;�,c�!`�)D��>��뒷'�ES��8��ws�W.��Z����mL�X�M6ƻκ1z�f/�v�sG]��G����;�xn��V+�N�ְ歡��k�d*�ǩ�.��
���I7Y�mT�v�}�����3���c�;�CK�g�Źe1+�L��u�n��̯s���В�2󐑖ӵ2�yo��p�)�Լ���v�~��}S��[������梷H���ԯ&^�wtB��3�[�������^��nT/(�u��r�9�}�>����킊�l�:.�m��18V���e��r��-֚�\GqR�'���GPm���m�,ٶ�([��
��O�<��~�����}��J�tc-:*L�����$���3[���Z9��dy���A=��f�0��P*��ps�gf*.�1����R�}Uk�7�-�{�7��}�o:E휡J#c�3=��m]+G#�@�cڂ~��3q������P��4���odv��ףE�9)��	ގ�`_���3}��vu�T�T�o;Xk1���{�0�_V��:6gks�^�{}{nK�C�I{HIOQt=�)<�x�l#&A�rz�^�V'�R�k��amvwV_�ޗ�w;W=}W�o��0}Q>��=c|ƙ<�SV��G��m�qර Ϯ��}c�;�$�Q����m/o�۰�s���d]��x!�E�
�2�.���=�3��N�C��6E���K�}��󖶇>sA7��S����6ᡵ/HZ)G gw�����>������ޏY˜:�M{�q)���9�=N�si��0�����N���V[ھ9T=5��͍մV+'S^XÖC��B�Ƽ�3���[����5j��e*���p����
�Aj��7Go.�Ι�@�,�����j�#ح�V�#���h�¶�u��
tN�.U�G�RL M��"�TS.�hu³��������	�����Ԯ��~���ۚ��o*ֳ������}g�ե�U����<��^��'�:R���Δˇ��>o��/{�O�]j��p�W�����V�A'W:��O2��]�W�{��Ʈ5:����T|�9�Tbu������,;nJ�V#�i��������,�BU=i6v�u>=�]ڸe8s��'v�g\��,%b1��n4r��æ����o�����n_Y�J��څٶ�����@8�
���wW�)���[���WЖ88b���3Dr�'k8u-ɛ`��]z�F�)ȃʽ�=;2{=������S��k/����w�y�V=е���Q�9Dt�P>�ʽ�),�P�ӍSS�
D��Ք�d=��*����kq���PR����>��pj���Lp�Q���9=���mk�O��}��v�S��e�0��ݩh�4T��iUef��©
���9 z*S\D���l��_gV׃M�6�i��NT�N���֯��^� ��,0+ov�&�˚x�(��o��f�ek�iZ�KT�E������{Wʅ�v��k}uN�9�S9s��Z�S�n,c�L�V�����/�P�W@a��,�ov�)�b�A�ƶ�Pk�p�q=��_�dy=�����`4Z���q��z6��V!��a�P�>�{���܅7�V>�Ut�GcN�o�r
�4&�mX�M������.P\��+���1��F�a�;tbyC���G4��煾e߁��xZYy=�nU����0�cZ��׆9�`���*�szԛ�W��0��wj�t��=��ΰ9:�Xsnbڹ�f��GL�������/�׼�|�.�g�׾v���'�x)��9��c�;@e�voc +&aXm�����wJH�NXU���/1���xD�c��ϔ�7qo7[�jR�A�,]_��%���d�=>��"l�J���ʦ�+�P|1
�̰����U���N�Ļ�{f�7�u5ĎS^���ȷ���g�9��G:��bۮ/�#�kK`In�[6$�_�����5���X��(�1�}N���f�oE���\��y�C�����y�5���>s���rw3ٙ�SJBP���s*�X�vj �IP� �U}�����`,d�����������e-l�� ���ov5$\�S��l��}�=<�|ʌ��J#gǘ�W�.V��:����Eo���]��.�N�4��1��z�'�iͫۙS��P�,��C��Oq��}�sX�T�%R_N��'��a���-���ͤ&9������@�H��}��1!�����_�ֻt�a���,k�b������
)o����|��~�$@ilW��Y���-}�iX�z��1Wx���=9�u�y�~���8ep�ʩ�u;�<�q��W˶��Z���Z��48��z��Zw���9ñ�W�x)�2,�)P��
�4:�l�̕�2�f����+[�WV��o���e�w�D�� AN�p��;�]8��K���_S������6�ibq4���F/To81����X�Y���Q��q���^ee=s���V+I�ߖ�歡M�9쫨C�_�H�I:���T�`\�xq�(��K(�;Õ�����r��@���'}��r�y�g�N �|s�@�$J�2��v��^��D`��xM����$P&L�ė.��J�GH�N�jS�X\�S��\Sf�Ǚr�YJ=��Co��Xe�uj�</�č�n�@�;�����-��ɿZ]��s��{�/W��{~Z�5X��m�\';�Zw�l��0��U�Rw�--�;-.߫������V#���hoB�؇#��X~^+!�ۓ���i��~�i_mzp�e`�\d_�.㻢&��{�62N���&K���g������d-�����,9�g_o��l��ݻ���}�HL�U�?[�v����^v�\�ݰ��9*#_]Xcv�U��Qf�A��~��YR�X�^]-��j�m��i��k�!�q��œ=}p����Q���X֯J�>|��s{cXk/{'J��k���2�UR���m�ͨ�r9Dt�������N�&{�~�����X�E�����^�{��6�q�
R��S���	lP��`Y/D�>�-ݍ�U�x�zx������+}���<f��*!X�%0��R�~�k�Iw��8kf��-�Փ<��9��;y��A���.�^�X`���7v;�ꖟIJ��8H��</a�2s����q&�2���|��AEQ��B�84ug�Y��{���;��kO+FJ���Z�Av%�#U�L�7��}[�G�r����]\]4��%�&R�z]�F����wL��(}�;�J픟`W����鰨�b�c���o/Jƴ�yien�蜉X��E�	��x�F�h4�X;���:H�=� Ց��Vj�O�����ep������b���f�7�5�ն�=�u�F�����Pa#����e�uB4���Ժ
�+9ʢ�����ϐpQ��8� M��z�p�z���Z�7iA�)(Yޚ������uё�š\��������i��X	�;69�)g+��é��}��\(id:�;4��E��� B�Q�m���Fϧ+���,��&[�=��V.S�mN��X�V�C����j�tE+���T�7��\w+�8�Gz���jm-<�2�V��=��t���O���6T���7��xԃ5;U�M�;l|1�띭k]<7��o8>s�����I��z���I��N0miP��i�d\��T�ş:ЬR���A=�$@��彩�P�����e��t��0
�]��wjV���0g<-��yਚ]�x�����t��]q��,t���+rn��]�r�����e5;���l��j�\���N�n�ثLگyS�0Y엤�@&�i�+�[�3�o]��p�K�d��J��Oz�i��ZVCm��3�Z�/�ǝ/&e���y�/z�����|���>p�پ����zbu"���̓3E#��]p̥ز	��'Y�����j��x#J�8S��l��w��;�4?tc���Ϳ�Tٴ8Y��+�yfb��~
��s+Ԯӛl�s�Wp=\.���z�B��L�孧�
i�$�7� N�ܡOš�b�)�L}"y>sj&�Y�[�$��ئ��Ro;�	H�3w�ۮ��^d�E�Lm��7WMA�m��olf�M��q#;��R���P�;n���"K�K���J���3.=��ot7��b�3j6+�AZE��-�������;�8�y�\�f�8�2Ɣ�e���'�բɍ2�����-]�޵��؜�&�E�E��.��^\�(oh�`&��ߴ��a�4�=���`��U�f�L�l�+<6��7[٪�QX�e\��wU�i#o!���J.��9�1�}kc��}�Z�ul�ot�������+q
Imr�������������ٻ��t�!1dY���h�ٜ��'�t�I'uׅYYM����DB��e�7v��,�w�����F�^,��+1S�a��]��He�����>ɩ���k���WJqov��l��=���Y��y�k���]Pv>�qj���2�p�u�:�^Q���&h�f�tEݸ�P@ "�
����ݔ��N�1����@�d��JJ�X�q�f	~u��[�n\b��c"�Ta/:��"/���IJ��&P��*	@�r��ܮy�M�Ay�1:m��)�wtT`�$�x�$�����I.�a%�n����rx�ʝ\��%��.v�Is�(�wvH�K��M��幼y+-sSιyݑ ���󸄍���bwW#cE%wW�h��Ν�,X�*M@���45v�M��·ݾ��]����>����|o4���2iRN�@�p��iJ��ˎ�Z�ʕQk�ۑi�Pn;NS����t�!_���3�%ubA]�����.�"R��T�像.u-�Zb3�_�����y�Fs�<}>���Vv�Ւ��"��M�G��rb��o"�k(F�v����7���� �T��M��MӚE�Bc�)�j���;^�m�V|��GD�����s�:��ۓ.k�E��i�--�r�>8��*6��U{^�k����fu	y�<��s�qyWq�Мy�>�I~�o9����y��z,�.}|-P���S�x�ڹI��w���s���;��[�=��f��C��+���7\�2���ΩN}ìS�\�+�f�*r���!��;
g�����t��x|B�"�V��5��'���X�w��o�(41��0���O}�~퍝�|v¢WoO]t�h:���[g�Gv��DU�.h	��v⭆�-b�9�K�P^����](-1;�ڷ3���(Bݝ<������uv����A����9Ou����������6�Wjз�+sf�,��n���c�* G�K�pu�q5gF��Ú�L
���U}p�Qh���S��ԧoW.軔:�?Orح�v���
s���mQ��lٛ7�~S)�K�'_{�{�^���z¼߃����G��ob=���NdHy�&��+ۉ�b�)�y��9����9JR}���	�j���й֎�[�z���yK��[��gy1���(�F]�\�s��G�[��бo�X5�(�)��yovp)�kHC̊m�Bq�vQ�u$�/a<���^\ᨊ`t�W�`�]5<�� �t�ms�C}�����=|�_-�Ug�\�[ÂB�3�(�z:���Z����N��_��K�%N�~�~Q�o���ۺ��9ð��B�!:1<�f
��J��\�{-�u���U�$�.�2u����{���M,a�6Ƶ9�s��E����B�NPR� ���S׋����ϳ��h^�u�N�kU����V�5�Tr���D�A�n�1*-ϦM�s{�v�m�5k��6:`e]�S<b�-�֞�B���������
���fЛ�\Uԏk��7JݎUh�(^��X=dWZQh�P�ۅ���y�cנr�� ���!�B@J`�����*v���c3%rS)�a�ߦ�[�o�lw�2��͎k�;���Dsܤ�z��qC~8tO.����>��p�ڼ��Q�k�u(n�p�����(��UW���t6���z*�(��=^�/�}S{����Ѵ���w퓖��8��iy^Ƚ������F��ө�:�Y�L��J�*���=�/bF�T�vZ���W��5�����|'����ʋ�WT��O�<Q���s:�t��a����:Ol�����(��s��wd@�|Ɵ�Gv�T�x�u�N��5'�5���0���?�E�(k�^�nq�g�N3�3�V���k�RVֻt�h�,rƻ���1��p�F�趡N�hs�c2���Dy%���_[Ե��m)��gi�c�)]޾q�l�.M��<f�y�2����U�y�ΞU�J󬬋�ͻ���nR�y$�汧����о�X9y�����!]�N�f�&v�j��:�4벬��5�J��8K�.@��e��/Gra�/�h-9v�I*���p�CeeoYy�r"��$T�� �:}o�WT� ��W��v�Juк%�Z{&i2�N,���wx߽/����A�2g�
U�`j���b�csT�K�ol��o�ey.sA7��0}*�VWg�����{4H�u�\h1ʆ^u��^�G{�jqdf��V*�����A�5߂3#]�p�FSˇ4�Nbn��)��������z��[Aub�����9�[B7��;����J�s�r�����\ʳ�Is�%3��T�{~/W�N�;3�k�Hw�Y<�.z���MQ̞ �˭+�_Z]�|��N�7z��g��e�=9i��ς�������Zy��gZ[��^����C�H�����ş{�Xw�z�T{�{1�Y�Q�����E�����~hq'�Tu�[���:��ck�ki��5���rֱ���9�ٯ)�B����Evسxd���]yQ���w�.juK\���a�������o��W*gd���QF����i�E�o�Պ�۠;Z���6�Koػ�&���&.b��hg,s�V*R<9�7��;y��ľ2n���t�=ÎV�i��)@nj��#S��[0]J�����6ॡ�|�u]Nh�1Ƒ`_��)���Y�:S�m�}�����l�s����Xk1��4n2�������{ac�շ�I	��q �wEa���E�����aw"�'���تk[�v�y��E!0���ЅB[�<�ǒ��������<��;Ħ�O�:}�݊��r���|~�we����+{�ў�C�)�����n�ދ�M+�z�y�^��_p���$�h��q���ѻ3��yv�G&���s�5��C�͸v��dv6Z����9)�97�)y�/\ܮ��X��ï7�49�'	�3�Z�/�r�|�����yS���=���+{�7�zj�N�O�~N�'�ݬ��3]���~�aMy6#k�V�1�� E��Jny-�����=�P���y���y����t��ܽ�����oj�sޘ=bo����c�&
����֎r�7�~������#�9l���Ѻ3VEp:��0gػz�b���+QOS��(�fb��,�-qVe"���^˷�`�7�5���^gj�I�ӣ
�5F�j�Mt�պ��J��V�f@��r�7��
-�Й�3'q�]x���Iڙ{c�����(}y#�1�I�="�b�I�ǫ������9��W���b�|ӵ3�ÜZ�c�͙��y�Q��N��ȭ�'im���8
�c���.n-�z�Eʾ�s��^B��ܳ�g��'=p�f7�pk���NhN����d7 ��K���5�ou�izr/�N1ϗ���:��V�{��{rzWg���-��ﳟ>���6�1�)� ݡ�ji�Noz*:}��� ���V�K�h���R
?k�O���k��y�^
��|�Snd��4�"��e���S�8Y�g[��Z�S���;}����r�N����O�y�g'8��_.�{�y��ǥ؎ͮ��	��޻O2)��ιt�B�q5L��V��9A}�Ou;�<�q�{�BS�b�Sj<����\��F��;Pʱ۽��)�p(ɝm�K���B���%���M�KX�eN4"� �N�pd*gv�t�>V���O��F�ƭr���T���h�p��V�h�{{O6�
<ZA;��*�-�6��Jݫ��b�T���fRP��Y�ʝ7t�э�I���d�o]�������;^�΄i��O.�Ѽ��6CF1卫��}��SM'�c��LA��;���T{,�໋�S2����]�X�K���׊�]SC�9m�|�Uxb})�س׭��G3��C��3�����P���7^뵓z���mkj��]P�ZF��{{�\x������4���wҲ3167)�/4sc��>��e�^�0厛��Ws=+(ԙ~���� YQ<�,v�9o����0¸��q�P ���\�6��نI�՚$��7-��~�)5�0�7.�v����7���~�.z6x�,�����ڰ���ە��LoM�
{�Gd��r�����Q�R��/������B�F�	�%<������P=�x�<��oGj�z[�l7w���)�NwTu��"J~W�nY�%G�ܒ����=�����r�}�ѥj��q�n<}&�H̏6ƨ�F���ݻtn��Q]޳= y��	y[�K�:%rYy�q<���ڝ�ݦ.��X��uB�qCnU�)�7ioQR�R�}�6��׵�ڹe�S�Ћ�J3���ݻW��s��=Ǫ���T��{z�U�ae7�dԹ^X�PM����V��T&1�Ô?w3�JJ�Ӡ��)<����QYRb(��oz�3�V��\�J�Q��}���毽|��?Mܦd�ݛ���c�.+���,�`<g�c�}��Q�LL�����-�Zsmy��'�I.'�s�B?'��g��Fˍ�.�^m� �3�	�>1�a"&����\�WzU��iz'f7��L���r�rk���,ۈc`b�Q'�;lcpS7Jvq�6����NoI��O����3"��^�ޅ���ϛ}3'��ɒ�n��#�b�������k4ʿ�̓��C����T�͊��L���K��!~I�z�X�9�co�"�8�꼚^��Ho�ׂ�w6<�\����(y\�}����c:��Gg2�\3{�j��gH̞Sr���u�G��f�at`s��[�NO���q�r���v�w��\x��X|�5�(�^X�{9,Z���D��;
���1t�0�GTi��m;�����l�x|��ȴ)��ڒ�c]M� =`�pF��wuX�}]\����h|S�UL�]��|`%��TQ���ʷ�=Zv��۷R�dM����>�M���讲�?��S�e��'>��Χ�_fV��rN_��:v�2�׏��Ҙ�����w�H������b��r�����y�Ns��y7a%7ǆ'"�9?���Cƴ��zjNt��p�kD���ʕG��!(��VL���,_�Cgo�[^�Q|}���Κ����o��8�聨����C��N���4���~r�Zr��~�{��΃wN2K�z��-��>ܨ�d"N�;���^ڙ�q{��Ы�J�yssb���p����^e�muߞ�o۲�n�zn*<�EI�C�$�!��@mJEg���C;�[�_�w�]������ދ�~�[=e��c���/|�PU�4L{�@b`���`��^��-*�D�;hln�n���4��>�V��OCu�C4�aL��玠e{�%�(�Q�{�Gt�`�B)D?)�ܪj�M�C�R��X��Q�k�z}���|��w��ݓ�mײ��ف��2cO8~���O�'�:�]S%�s����12_�ʹ�����Y��}Lz�}E�q�I���� �A�:&��Ѵg����o>-�����J�({�oWk"��3��wzר����O�p����*�nn���+sX��&��*&�r�[�/�e�W}�%Z�١W�*�sՍn�8ĬT!a�归ɾ�]�h1ژkO,�Oz��O�9Ǹa��[/�>s�J�Nt��:�U��,�al�5u�+ٳ�.rC�UH���;�;v'�{���UZ����p��k�!�u0Qd�!���};�Fܯ�Vw_�O�gd��[na��5]M>�%Z��遦����q �=?ai�����;�?�^����T��e?ٺ�zהּ�i�+���V�/M���z/��s��yt+��d�� tɸ���8y��w����2��	�.tOѰ�7��l��*�1/O��s�G�ت�r���3ţb���2Y?���+���☳��7��y鋓���(��ݐ����(�t�N�Q����n�z��5�&�wz9fl�u�~�R��Nd[�*:����4�#�d�/��F��L���3�y)^���r���w$O�n��d��B���P���}F�D7����޲��M֬���M^z�MM�6�q�ܰ��.�1�:'�ۘ%p�f|cg�^ډrLc��
��b[�~4f�ϱ�/2wn}�y�q�M�B� �*���%�w�l��1���5�i��;�]�*���dTY[�pZ�k#v�זph�j+d+,J�T�W�m��ث+(h{�v]TJ�Z�O�͔���#8t�v�gM_H��*�'k�u6X�1n��M=��HŘ�1`��U�&���ʕ�\:�����j)5uoJ=\fs"^Fhn�㜺��/�[]+5T��/YՋ��1ⲫ/�Fno]�d�v�9����]'�xYt}������JU��"�]%܆���9�M�wwK�^�[,�w-�֦��z�3%;p��3�;�c��ƛ6FSYO~z���,���an�v>x�fN��a̽ͩ�����\־YS�³�]�AW>�mEfP��Ɗ�u�k#� ��X��HM�X굵��A#G�`������V������@w���F�� ��� ��0xa/��z���K�y�x4c|��@9L+&�Ӝ���2�^m>Wx���r���������Х� ��=8Sٱ,|_c<��N���[!��2ծ����T�(�N���a���I���З�ˑ���u}E�nZ����T��i��@�x�^���,!��cն���&ą�l�c��f�ܙ Xj�cu���o#s&�&��!�˷WP�v�d�ש��c�Ӣre�hZ�<6���4�u���rʲPL�;@U3����e)�7{x��ހJM$ܮ&i�/{�q��Y�* �l��/C�,�.��re�7	N����s�@٫�
�x��j�i䕨���+�Ɉ���x��ɋ&�l��z��XGx�`����A}֘5�C�\ź����5Y�a8�]�{������:|+9gB��b9L]=���\Y�%7@���RV����¢���;WQ��և��i�i�xw|"J<���c��(^G��(u���/���]2�vM{���x���N�G�'��u״ᱵ�7��5��y-B�� �(tS�,�s�Dn�<F�f�!��i֭�p�$��R)��U��rWo2X��FP��5Cuǩ�H�tM#p�/Y}� �H�)��/K�t+gH=�d��l>}����؂��<$z���T1���S{�T�X)ۊ����>��l�M���+��s0䭑ٻ܍�蓑��Y;��V�jØ��	@��O�v�(�C֘�B`ڸ�q5�^�l�++�C�L���ư@gC#�םF�.;df�&>��τ�v��د�s�E�%�� �!���p֘�nu+x�)n��N&Ǝ6mrS_�
��mJ�1���|&%Ȝ�H|�oU�N|3^�ojv��,��X��>�j����AnU!C�v���;ҜB�h�Y:����m�ɴٴ$�9Ry��c�w3���]D��"kM�34P��Ʀvb��Q�$v��1S�ٽbe=
�^��7���;�gn����ꋦuujɑԆ���>�9D�;u�]�yv[��u=|u ��w�]�#��1�64>�{������@k�vy���&�Z�2Wwx������.�;nx�T��-��s�0�x�N�t$,׎�e�щ�\�I����6��Ii
1csk��s�`ѳλ��#Źwq�W3$1�Qb��ww\W�ux��E�ݮcG��h�sb^u��7q�����r�	��3Nx�1<�Ӻ�b���M�˅�G��!� �����>�{�}g]b�����\���b��Qۻ���PX����n�љ1��'[��)��өf�[�N��J�q6���ص��l�8_j7����S;ІR�,�Μ�'ڕ<7�8�7�p�y��(�U@��S��Ö֍���sE����P/k</:�Q��9�5���n�JdY���F+c%M����%US�v�����2.���x��|\�AK`�؇�����k�
jP�P�vgj�g'�fuMV�(����'M�N�י�ʀށĉ���~����>S�͢,>�P�/'>��72���U�=�K%ߙ���q�O�*�O��6���׎ǣ�\����kr�j���a3{j泔��Yw�O���5�Kߙ� �8�L�cc��>1�'�7���dz��]���n���|�0���M.{^w�j�J�Òڀ1p���\A~�G���(;�uCJOS���[�^�A?�0���{,v�,+f������Z�.Mz�xd�WF�����ŐQ���g��`�.��/�Q=?�l���©��
��N���(:ܪ���{~��s���\��fkm�Q������͏G�44�w`���#}7?i�J����q@m������F1$���o���$��[h:;�4gK&��b�����"$w6[�j�񫋡;�"��!ܩu�{����^�֞e<�..���4��k��s����::���DP��]w;�vuo����b���r�Z&(�c�[�I�;��8	�����eos��r9?z�ú���U�q�=�eL(d��C�@��uM�᯦!��zl\�d>���7P�@��p�n��Y~�ӣm\蟯c$틖O�@�f���\(�s
���Z�mw����#<#O���Nq�=��y���}^�w:'ݱppW�A'qM���9�2:Q��H#dP$g�ʪ��_�~�*kݮh+��,W��eٴ���J����8ۚʟ}Tk3/���yn���ג`�1�@+����1uT�*TH���4_���n97���z.ڒ#bs�x��������[(D�s�+� {�$&�����μ�։�I��${�bd��ڼ�r�"�E?�Hõ��fT����Pxϴ��c�ҝ'I�U�S��%v�Jؼ&y�J��u]J�6�1~*峹�s�I�~���_����#���ܝQ��U�Ew����]� ��{r�ښZ���������_-�>���:Hߋ���w(���`��O�A:=�{�J�~:��4��=��Ӆ����T�t_���{�}��\��p��m�1��FpeD@����&���4�i������k3=n�t�'�����q�G][޺N�V��p�ܤ� nq8eu�m%�l�:�
�|_t�h�-��ֻ��UgH�����Mq�_L�[���fl.�^Px�ms���J��1M�l�+c�Gz�2�n��v���7#G�`a�q�*�s���q[�ފ{_�U���.Y��o���oJҹǟ7�R}\ӣ&��?u�]�"U��3_�;k��U??It`�Ng�ǞЇg�sb���l��!��.���Ng�^Ʌ��<A"�z2�F0�_. �~�O��4i�O:�{`Y����9������i�<f:�\�\檞��2���!���B0Ӹ�<�`]{!��>�E�yg�7/O0�5�uT.Eڳ8r����I���j�Q�Dw��sQ�c�u1��]ЁÕ�B��]����G��-���We���LٯLBd�ò�P����x+��cn�Js�6M��W�Yt݈�3E��n�tQFθ�"#Cه'��!���`r��S̱~u��[^��0��oN�����ݮ�wζ�8��@ݓ94���ƨ�yk�
���*ߜ���1�r%U=c���(J<O���{k����oѭ�	?zqg�N,u�*�p,���ˁ�`�
�ɢ����<ιSS���߾�1u�����M�U�<k�Y'��B#�"��p~q�=�B�����j%1��Wf�vM��"��uҊ��m3Gr�[[�&M�v,��QSqt<�v�t����Z2�}pLi�|����zt:Y��_oW_hu�'R��yQ���ڞ��I������^��%s2q��i��59����D/.�*��r��8h�����Θ_)���� �6��~�w
��|k@�j���=�_`��O��|��zj���{|�`���sM34�j��#	=��R>��Q�Ԙ�:���2�.7a�#a��M��w��ݒ۟\�ENOW�!�J�Vv�������#|�Qj���B��Poy�;������{�S�&��=#�v�{T�wm�b�;�6�ϳ�OG��Q;�}��(���'�u�+����\�V��B���C5�ܧ�Uw��,�ˈ��66!�u0p)d�!�~�/�t�ە��u�S3#���f�f㒽A���h��Ԛ��9�7L5�&�kɀx�{<����c���\}����J�]E����q|{��Y7>���i����z/��|v�o.�qyu�x�55��{:��KD�с�ܱ���ZN���&kr�y��b^�_���V}���k���Ą?���������z�\lq��~X<����,���e9m_��)�v�s����1�@��B`:�Lʺ�Y�f4��
��qe���L�'r�)��o��vbC!�C0>s�ڧ^}<��Y��gi�3<J��y>�1:,:R���<���0`�e����Xв�v�I�!`�i�Ȗ����Z���*q�oFu�Z������z�=�w:@��m����#M�����
��Y5��eHX�`_9�`�+Ê��~���޹<�?�L���wy=3��M�,�����6|�i�I�N� ��>��S�K�/����:"���nyܰ���6��b�eLmܲO��4���>��������Z_I~ʌ�v��-��8��c�7�~t���EN�����B��f8��[�=��'����<��p�z�If�9�5�J�������Gi�W�ًEM�.@���N��:^[�`����:9��R(wتu�t焖煍玗��wo�rP3�¼^*ߣ>ʭ#�E�f�1	QtbD��LX2�q��GR�\4\6��P�F냯Φz�֬;\fq�Kc0��ף9s�@�x ��|y�ɹ�\^��O�R�K��h�n�L�����0?n%L_Ź�]��XD�� �n��Gx�H�B�ri
��ECw1x��{�i�ד5��'ؗK�ɹ�[���N>S*qD���~;��b�@��iU�YC'�aNA���(�]wX�\d��u{;��+Mi�Q՚ݮ��P_{����)>��"�3G C ��8����z�aGEcܾ˺X�EV���اBWE�k���[{m�N�iV*��j{��mo}7���Lnպ�Pp�w1��Ɏ�^mdot�8��P���u��oB�_.{^m��*�2d�y� k��ʡ��Aph\Fo}��jyȋ��"���
(c:a��X��vV��s�$�����\�e�w��˕wN6����w��Y�/��J��+6����;
��;�.>cr��__�ҳ��meþȷ��c���U�����QA}�8v9��!}B't�W�r�ѕ8^u U��7��n������Of�5Dl�m�2��sCt�۳�Y�T�"���!Ꮤ����L�:����N[y"�"�}�f���i3����N�_�G7�z�F�Sï�s�ob��}P�c+�e�Ɋ���c:)�U�^ǵ�Rk��^;*���d�8�^���͞�}^ݿ<��ظ8*�sLɸ9�3	ɾ����N~KF:	h�+c����\H]�.X5nC/���J����2!����)��r�[�]�z�ٌ5[&Q�#�\uJ����*Y����X��4^�9C"���=n.����+*ﲘG��-���xT3�,����=� i)(�>�^t�D���~ҳ�2�����|�e��cևe�����P�:�u}Yz�Pt`��fV��>Of*jggk*�}8�If;��ۛ�a���<���Ȋ�(��c��l:)p�]�kv�u�4���q�އ�B��u}B7���:�8��7O Z,�L����7��=��/�M���A��%����Ti�m(�.\��rY���P2H)N�^؎ef���W����{=bn!�������^5^��'��:��99Ѥ��Sc�A̗*"!��~�^Aq�l?�v���F�vqZ���>�5�'�^��#~./Kg<^Nۛ|�ى�%q�{�6^���D��F�6�,���5=+������|�����Y_8�d��3�zo>�sT�Zh\�G��Ȉ޲��O�X�Y�dg������ZW8!�}U'��iѓ���7�8���~�=�]�%;��a�d�C���Y;"�ϯ�?a%����u���W{7/2�.��"]'Q��3���������}���j`����0��������]P��ҠW�O���ww���Rٕ�ŵ2�ߖ��[ڱi�H������D煎gd�Jn�׀Q^��^Tuf�����.b���	���*b��3/TF'>�����}�X'\\�l p��u��z�ݖzs�i�8�=zngLF�xߎB������Q4�;m��u�Ӛc�r�~������y�t��۹2�Q�!{��]XU���%0�6�Q�|��w�˹��j��I�3E�s�*
�kY�����1b�a9�����]��!b�vӫjvN�{�V�
�ޤDܟK������4�[1N�;��圮��t��|/!�����_q����X�Y���Ip���c������+8���.�5�y����Ք7�_��!��};x]���^}�Dg\Κ�K���J1NΩ�k����#Sy�'�]a�kQYf�U߱�����zpx��R��ˈ� ��N/��WҮ�а�@�y=7�+<���JC��1:�x���r�N�zL����D��^_O��2>��8S}Wݾ��v�g����BT��8F�{-yL�v �*����N�9�u��N7�ݯ$�,6�)N^���3�z^ϝ}�q����9�'�s��%�;����c�<a�uYKTˀQ�g������A�S(_�oG�N�>�{M.0���!��]����]��5��g�	S'�>YF'�y����g.ޣ���B�����<,��/��+W�]���l�"~ύ^v�M)d�D�_X�� ��&��Ȟ����\=�W���]~̫<�m�#��URP�k�a��ѯ`�wP����0����Oжs	p�Y�o���4{���,9?%��j�\�>t��W>�|��[�pW7Cit�씦x*[}E�0_\�F-���ym7�v�c�?j]���:�.@L1��U�U�/���j�!|��� zU���/-=��:oR�F�}b�"/�5;x��X3*Ʋz�9���h���x���{��[^�5��i��L���9�7L.��rhk��s������[���e�lD�hO�!����~�_o��y ���t-5��e{�9�=�@sю������������y��9��<�ã_�#�ܱ���ZN���&k۔���S����g�Ϫ���+7�L]ּ�ezRѱ߿V/J����Y)/�1`�j��>k��9}������_�g��n�9W�`�pb�xَͺ���Yo��١�lޟ[��<7|c��C�}ՓZlʐ�����%�G�����P*��K�0��R�Kgo��Gq��z(geN����Y���3����"�q�4����[��؝ƺ�0.�jd{_�[�+�[�n5�0�K�m�.tv�@̨D�3����?f��6��:�Va�����k�P�3^Z����\�7�py�|���Δ��cGo��<�ՙP<;ε�����@���wO�}�2�1��K5�4&�*zo\V��v���d^uQ�]ha�s���OU�F�$/�@��:9��i���b��mӞPݨ����m����{^���}�CjM�Y�%?v'#�=�9j������r�\W;K��%��\X�A��y@ڽ�����zu]6:��dZ��]��:E���Ѱ͒���3�6�vVW� 2�k�11�c��c\N�H���G>��{���̶)�C���^�#J�й	��9�w8u%�_���fW��Y�
��xݟ$����f:�宸h���hh���+�on1e�U�<�N�m��4�ףy˟D��g�@J~��#�욝�������|�e�+�0������j���v�XD�� t��ĸ��#����;�ީ+	�f�iڭu����w��^Lן!>�K�ɤ��.ٖ ���PWr�:/n���ke
���~�,~��r,O�����gd��-5�.{^vڪ�^�d&L�m����P��[~�wC,,���D>��ƍ��¯�;ŵ�Z��j�����|F�
���tO�r�;�s�,�^��h����xb�{J%Td��F�ñS����\O`�v�`c}�\{�ff��"�u�����r9B�5W�6�*�3g�N��wHz++�4eN��b�2hvW�L
���*o�� ?]��-̺�c�es��,��w02Բw`�g�Pb�n����-��Yf�˷
WY}e�b��%�'��;�*�I�>��W�z9,���rv�'�� >ºI��n��&������Uij:5K��ҫ@��dC�t�͗��/ ��_ZzȷmN,Σ�.��y��l� 1)S���m&��l�����8Rv����53�qv]�F���2Q�<-��ͮ�:��G2X�hS���pG�t	w��3�A涇VbF�J�5:��%.7Xn�n�n�yW��-�29��2��:u����MV�e�Q��u(�n�=�i�Uݵݢ��I�[z�-�S�/��3�kX�s�"�0�� ��n�uӋy�:��c[3d�����L��k���v��}J��$���b]�UK�[�;�hus���X����37���ᯥج�ps�on�0Q���;O��h���w�/n
�m����j�h:�%J�Eݭ�J�+QX�����7OE��؏�Ʊ֒�!{�סq��:r��dJ�l�����$�5��n8)w;C�C���랛]2��u���qv�E3[5�O���`���ז8������q�:/�j66(g>ǹc*qA�r�J��sK�F����uk��%-r�8�Q�<�KR����3{�gV\73���]u"�	A����w4���e�Z]���5���*�k��G:�=�YWb���ku_U�v	��ۓE�B�CD�t;��ut���W�-0�Xc�
�3��|/o�Z�^kQRq5�t�t�6M�݄��xp�X��BU�u���}�����W�P�!m��}�ƪU��6���_�	�g9��Uu)+*�tܼ���@����2zk�P���E��{���G���_
9L>C.�-��Y�����L�U̫2y��>V�����DuF�Ɍ*Ֆ�ܻ�ݫ��[��y�Nf����VLGa1����B$]�1���S���r����NJW^"c�joI��k�����B�Z�:�^
6ة{/B:$�#gTW��.�rq������J��M�spO�K  5.>[c�9D����.m��7]}}�+rJ�(͎���k	뚃�ُ��.�"%�w �3G	z,ah�D��(=��`��X����K�7�si�g	��<�֋�B죟zmR�����v��A����!z�Y�p[��|�N7�x 5Np߲����z2,����l�ˣ�NL�՚�\�
B�d�]P����(n�;��J����o".g3���L�1a�b{�]=ִDn[4�Ż�ϡZ��.RQ�?����o���<��׺wk�l�̠��]a��u�"(p".�˅#Si8Ұ�(kL-�����v!�N��Q)c'WP��l%��̖���r2GN���xpZ6��Ʋ>�:�P=y�D\�f�]�N\�$�:opE��o��
(5�����umZ@��c��|).��z��+zPU�k"���9�ǑA���n�޴��v{!���uu���2�9���i�y�^N�
���ڋ};{sK���+�(2�H}DQm2�nRh5�kŞu��[��(��"*�/:���W����W.s���M�r���\(ۜ����wv�x�Y6y�s\�'w�^<ٜ��μ]'u��Ir�s�+��C��wrF���[�
ws�����؉K��5y�c�rr��7^v�<ve6%ݷ	�pwbNb�q.����[�-�ۜ�x�75ҹ�Q]܉���7Fع���4��yܣwq�\�\��@f!p��sr�q.nn)��*�|(��f��XF���]P��6�|����� B�ڻ2���=ǹ���2�f �m����/z�}�p�P���vJ�q2�\��4P��*�R��_�G�;*��^���S�Ω}^�w<��v��^_*�y��gꓑ�K�L�u����꾩+�As_-sA^�,���6�6z$L%S>î��W�eM�����#>�a����ڞ�f��s�Q"s�N��-��T���,������{���5^{f-�*�<g�,��a����BJ/�j}Ud\�*�*�<�,fK�T$?�Ҭ�Z=�k��k��0�Q��%��G��1�Q��Q��J����}���o_�O��Z��5��r��y9Ѥ�����̡�����\��/1�o�yu����!�)N��.�)��-�>��ܝ$C5��ł�۬�ql�y��'�/l�����T˂U��$8�<&��qѹ�Й��'�ϥ�L�%�l��W���,�USPo^]��O��NI��:�J���At�̋��w�Ҵ׼����>�k]�g�y3C����y��x�����o��O�d�E��}����K[{ۯ��wS�ؖ����	�oי}V}|9�t��-��t�C��ʇ�Ge.�֜(�&`�G+�k!�a��ꜧT.����Pۢ+f4/��[��[!{�2��Ϩ�rƈ�	�N$�\���
z�M]�Ր�emd?oe����,�\�:$��j��#j���Y=׵�[S�/3��U��3!���+�nk��
ד ��'����k���2�W�蟬��ν�ϥm+�m#Z�S+ە����e�-r��=����7�HK��q���|n�.�����x���]�~O��t��<'�Cf��J��)�z�19�5�u>9Yu�}�.�?u����m��o��;��)�6u�+3��M�ᯉh�5�p�'��W��L�,�&��mW���!����DU��X�z1�?Rfu������j��ʡ��KUFT���r^���9���a M�u�j�6t幧�vϳ�������e��e�P�<\_]W�n��2�}4PĲZ�(���ȫ�_9�x}�R�_���_������ڈ㞢�;&<��(W��3��gp�K�7ߣ��lC�Y�誕R=���`��ٵ�r�N�zn.z��F��$���e[��U�oê��U���Μ6���S�U���Śt��5�%O��m����Θ^S(*��+�MQF-#��@��5�m�� ��H� gK��ʼSCxߕ>�MCu�o����)�g��t�4U)����=���h�"���+��]��y��(�n����Θ���!�����1����b��t;u���֋��OƏ
�u5�ZyU��B�U:]H�n�y��9�Nn�Nv���5��x�Gs������-�X��}�%�����n�8ޮG�xe��4�����A�i���F�-���N�>�{M����r�e�l�ׅ�V��o�2�I]��U�Dz>�<���
t���ݓ�.���^�+���NV]N�]-�tY�h���CD:r'�x�"{�}_Q�+�'�V���G��I���/za�x����E{��K�a���F��O��@<Q;��M}��}�yOjVz�e�f<.�n�7����q~�h���y�\�X�6�����曦�~G&�{^L=��w8�;��������*��*J����Yذ�\���=/�wB�W���ruZo�-r���s��]�J7.�F��YQ��j��r�K7u{�#�znX��ZN݄���Pa�����ey>�����@����U�E��[���YhŞ�^������v*r��Ԫ�N�]N"����b{ͅv�
<�,ܜ�Y��#Z�O2��j7xugC>ʝ6d��2TOȸ��j��4�#���<��̽Uv��1N�w}\�<��8�U<7J��onc}�(���Vd�ϑe����+�l;R���Q#��~ԦR��������� 8t�{�fx*
���
J��a���T]}9�e�;Zcy� �/-ŷ- ���ӧ�����<�mq��pP���6�ǁ�����M�و���WRmnp>�ֳ=���ڿ�s�҄��f�JP�
�Jc��Uk{w�ʮ~&��7$w��7��a��]pco���Q3�I�=�G[�؎>�ְ)�rA��<��&��B4�Uyhp��8��>oa:Rƙ���r�뚇q�#o�u�gZ�rLI�I��G���{je(c=J��N�НJ^�����p�و��u��y
���VJ]�f�������x��L  ts1Za"��N�n����-><��1��GT;���i�i�>��i�FW��>^�Q���K�#�R�"���sQ�h�y���qKx_N�joҒ��c�J���i�N3	玽\8�b0Q� %>��'ǜl�y}Ϥ��]w৹�Wom��w=��MoY+�rj����-�A�6�@�n���:������7'��L����VC!�)�59	����e>B}��S�^M���e�1߂�Tʃ������;T�	�8�_Q���QO	����4.�	�����o�д׼��y�j�M,�ɓ^m��\`�#��	3�Y{9[=�z�^g�"�WN���k���a�)�~�ݕ�t��o�uZ|O�̾�-�f�fu�.ɹwW���/�U2Qn!�N�_\H����_e2�=�; ��{5w(��p�e���EQ�X��gDW��{�h�9�W��V,�x#/fn�|�U��IYܝ�E�K��16p�]n +X"�u�"�Wi���S]�bS���+�8�gh���R_޾�k��Q�-�B_�:Z��z�Ʒ?0���� �M���*��f�	�Ѧ��77�MS���۲�}�T/���ʮ'��k"��_eNY;���9�|��r�ѝ�������:��������m0徦-L��c<��*�ɹB\_��'���Tb���}��������p��&O_�%�&�'p-Tsp\ǭds�ѫ�uΉ�����x�>���ư�f�M�qf}�=�3'=;��ga�_ar��y����͞�}^�]ah�*�c]��0\Ȏ���v��l�-I'�L�z�U�H�+�As^Z悿{K�[�����ɽ�@Ƽ�ɳȬ�?����0ע�a�xD3�?�Y��>��./����̩f����)�5w�E��W�L��T���TKЃ����x�#���y혶|�T<'���q�!%y%�Us�6�C����K=0�"����;���k��k�'�a�*|�Tx����	�z`��^��U=�_����x)�񥯫�P�_.����s�Ix���eD�n��u�][7�|���S57һ7�F�gtB��_W6)wTBt7P����pǩ�
v,��{,A���f�ҧ|{�7-���r�<��(�ؙ�S�'5n�U�wD�W�ã�T	K{Ƭa���Pѕ+;L��-��s��G�C�ֹ�����������!�Y��S��KxO��:Hߋ�����pm� _����	fc��]㝶zm͘~��o���^;GМ𚞕�F��L��{�}��}NM'�g����r^qk2�����;�kb(9�31H����zdW���E��K�g�S�a������$���үf��y���>ns�%2�1�46�O�d��z�$>�������0�/L��v�Y��s˿e�,����ʬ/�:�0�@�V$=y0������������(F9�i�m�'����t���.?�>�4W�+)��)�����fy�Ќ.��]��d"q��n�"KqO*�v6�=��^���	XM��t&w%K�e�N=��}Χ�+.�T�8c�,-�ΪQ����ヿS�a�s?!�?c�b�g=�y�ƍ��_5^w�3̲o�Q��(S�Ԋj"�*��,�~���]����#�%R^�Z;Z�΍/�~�/�u{���ڈ}鎓���^ܼ�Ӛ�\2��O#�����u���vT�,���q��cJ�&�:�"��[�;�I���<u�M�\5���{6�뫀ʍ�����U�����Z�W\2�fT��٨¶mHU���/������^e���N�5������C-�����3Z�`�+c�hM�R���Z��
��	\��A�=��<��k6%��Ҏ�']�5�y�6�oN���e_b;~r�_���_���1z}=�1ƾ��;&<��
{U���օ�ݜ��,����s�}.�y{������{������7�GJ/��<�O5~io"�W�.�2��D�����\Ƣ��|Q~t��%)vw�p��c��y�B���ȝ�&<�z\��3;����_� ^���CAH�葚z^ϥ��q����)�g>�h�vEu����a���:*��&���@�*��1"[��|e�\hg8�ޞ~�����ӾTSq����gqn�~Mף)̳|�
��%Cd�����S�y�������-^��ݾ��p&׳9fK#���}E��g/=�)ۡ4<�������Ez˓~�=gn#�gy���A���[�ؗ�(:|����sR�v�01ߑ�`��>�D�i���\:
��~�Uy�v�Ύ��Yٽ���_.{L[jjMyc�׼�04�.$f���vss�;�kg⎝��
��� 갯���pʜ�^������Zj�����N�J� 9�_�Ps��Gj�Ԓ��
�+��M�<4���V1=Lb���elX�8F%D[G���U0Kڼi�v��zl�jR��ו*����gX�Lwʅ#�pQꗴ��^I8>,�=!��k�G�i�V�������L/��wF��6{����睜���o�a�����3�p�P���nX���Ҵ�;�2�)W��LK��� ��싢��vٷ�o�ٟF~�����F,�r2��c��ᑁ]NQرR��:�\CL��%���TE}Y��x��?`{3��8�uN$fdVm���h�wl!�D���
���<�9|��٣�N�wz��4�Km:�`_�s��Υ����a�,���(�_Q�+1��Ό�gMM��4zgk�ͿfN��s�@jƺ�偹#��7�w,>�z]pco�s���k��<�[�{��ͽ%Wh�D�?	=���C�?Q��q,���vqr��8���כ�r����k�J/y��������M��h$�K�*���zVɔ���RY�NhN�/2�9Ug���hPyz�Rr��\ϯ�~]z*�����A�."@�+�68�e�w\ͺs�hyrV�DB�����ص3/B����p0�y�FW�s(�W �?w����)l��Qf$�S��n�.�>ȼ���:��V��˧����cs���4�ף��	G�����}~��7p����?m��;��5#�iT��&������U*�R���'+�0>�3&![s��h���V֎be�(����nC�>��t68��Wt��Pf��uB��Jﮢ�V3{<�� oe`[Ɲu��a^\Ÿ񩼣�~� �57d<xM�c������U�޲0W�5HYnx�34۝�v��*!�r�v��^��Qs�_I�B��A�b�&����ͯ&SB=z�S�I��]��`w����/+ʸ2�"�.)�(�<���'��׏E��=�s�I߷�i�.{^v�e�Y	�'vx��$ã��7<�뙬`^6r�R/"��̩�.;D}9�V���k��/;��j���ħ+\�{(�k��{(�W]��>{�Ҥ�(nnJ���1f���޳��ᓁT�Â�ԧI��t��ɩ����gM�-
^U`bڗ����#�,}4#k&Ďu3ga�gx�_�C�Jz2gu�ճ5�5�_QfT�9x��'��s��y9�U����-�@��B'3Ѩzӆ�&�NS�JN?e��鹜51��,>�I��Tspm����������_g��"��L8�g诣?�3���%� �ն��ح�!��p��w��wO�;7qo�����^��;=��oٕ���pJ��:�.t��[��Jz��h+��,����c&�9�T�*�A�3x�����lm
9/����}M�5�ֻ����״����v,Kr�'k^�r�-_���@�(u�#����z�R�<�k<���7CvQ88��n�L�<8�ш�V�^J�m\�`ٹ��x�1��v	X\��Y�{,��]��i{����U���<v��+��A�Ex@���>��?ǤK�cP��p�YWdU��hܴ%�ي��~��(e��v�U�b��
��x�O��{�@����U�4�X�Gm��.�[��~��O��ʝ�Rsc}�%�����=`}��t�r�YA�bV�y'���8�6��iN_}���
}�k寫�^���_�ܾ;�Nti/@������ZQ:'ND_8꺙��s2ਰ ���� ������Ɩ�g')����/'�;���j��ѽ��u�����`?\Z1Ē����h���ק�qѸ:4���+�}NMߧj��M+���x���ۻ������N��D_��'�QJ"�GbLG�ׇM���#.�����Zk^��;��]Y�*έ�ds��T�W�N��N��F}����<;�[_v|Wdؾ�hs�H��wK]W���2��X�}U�I�H��C������x(V��}���Y���1ҝu�hC�޼[x�>�!˞ôw
��Lh���b��e�C3���F�d�W}�1��,�8�uJ�#ルLܤ��A�}��7z��S�C:@��(�9�w4Wh��6�����-sk�Px(�w/���j�-.�V9V�W%��|�	�E���*�vEzy\98��ك)U���5�oFb�,Y���Ԩ��W;��r��rP�y��і�b[������p=َ���R[r���I�����պ���Ҩ�����^٧\ѭt.�Gn�k�e�t6,�����n7 U:��1
����mC��q�2���kB����Z��.i��G�����om*K�Sr3�s�Ǻ;t�8����yGM8/���Y�jǋS�Q�"�t-��|�ý�+����v$f_���M`Ի��CȄ�a���;�1���*����t���5b�5m���"A�8�qmqw2M��՘�Fu.�Rx���|�*/�Jζ�)�x�68j��hW�h�0)�[d]�������,�	�G�6�����D��ՙ����L���t�u`\�#�ˮ�)������t�M�]WЪ|�0���,��klY�wX\�=�N����K&��e�]l!SXG�n�}W��[���#3xh��6e��zC���/�_{#���X�Skخ�R��g� �Pƫ,�&T�j�)����R�g�"��u�\���º����l�W���
��H�9{%\ج�T�3ή���(�ǅ�â�܋�Z�%\��Hg'���m�:W%��WDm�C�za�|�)��I�wYUҿ�S��V�3��ݍ+�Œ�6�������b�����X�Za�|����q�e�Sk���{���rN�n���� ��21C�nV��&d��,lXUv\[���n�Rۙ\�[���y���*5��c&限b���Y�+��{�
�)Ւ�J�ӗ� �ٚ���Eow۵o�J������	�&Vu���L͇�M��A�8���v{�X�e���򒉛+ۏ�����wT��?N�y*F6L�Ό
��KF��p�W����;C�շroم����=e�bN�v����l����]�O��`uđ�k�yV�|�B-��ݮu4VXWuxũDoX�]����u.�:�Ir��ь��ˀ��\�]�1�.bucUH�����ɳmH
��D��38�=��%׫�ta�N���A:����o��KӺ+����nQjT����]ϑ�p@������*��o�>��;ϓ�rd�_!��w�n����Z�����@����Δ�lۂ�<i]b��ʕ�1���I�ǫW.m�!�}\p��kq:]J���d�r4Q�7�1D�Hc�worv��i�NN�n��<���[��i��'_eC����fm�1���=�s�t���u��Q�>�3+�58/bk�lSnG���S*P��m;b}�cY�$$پ]���ǹ���{nڗY�
WYz�| ��mo�+%%z�a�#�ڪ��E}IZ�a�X�l���1���k���r0:Evv�[���Ml���D��1���]y˓An]��î�guȣ�^/	F���.��<t��I3%�v��듺�;�غt��a6���˻�(�wn�׎��[��:\�ݸ�1����y<]wu�\��;��ۼ��s���w3�<�5��Gw�㍯�r���ʻw�b��+��Lgv����Mr�w3�͌b�%ή���]�j�ss�/�Dl�vq�ĺ��a,��F��K�;��u]݋��T�w\�;�B������wwW5�w<I������˦�]�]�˦��wr��H��5�wu�N뛤G7;�n�ێ��v�,xN[���78K�\��Mӫ���u����󫑹�\��M�&;���(��N�r�\�p�]�r�|.�����e>��>Ra�vP[�{�)��!-���v�	�a��������r�bV�H��=�R�k�͍����FRDww��_�X��ok�Օ�7S/IӃT����w�`���3�Ϲ��u>98bN�T�1Y���+��`Pz�
������un�ks;�x�'���Ds,����Nh=۳}u��t�������3�.�0W��Ä�^'GnԺ:/�*CQ~9���UV�݋�1��H�޹�����P7�:��ܥc��Dg\Ν���X\eA�.,��&T!���[��&�fwu�b�?�9���.X"���~�r��u<�:}��2'pǓ5p:�/��P�uѽvo�ͮ�S=*/�w>��T�.͇�~��^9my:A鸨���Px�ڋ�6n�����OK�L���{1̥�U^,ם=�Mz���F/c���Θ[�i
�1�����/C�UvЦ��8�$�"���l�]\r.�T(��w�#�g_��AH�Nۛ��Su}��4�z�S�f �~�Ǧ���A���(f|o�oO��b��ҽ��̜������<��q�M{ͺ�ey̳1A̖��jCwF$I_)���|w`g�����>��«2�[$��y�H�S�۹����F���\0�)ˁf�[���G��;D���oU���Mz%:߯*"����&fZQ�<��蓖�4��k�Vv���]��r�#o<0����p�3{�P�0�@�(7��{Aހ2��f�koj{ze�O׎���]L!e��͸�D�#�ኔ�'��D숏s�xF���O��m�K~r���\^��;���(:�����E}�K%߼�03���+߮ ]W/��lSv�T<,K��۝q޶GQQ���9������ז��s�b�SRk����04�G&������W���`.�\���z|���kc�����B�r�~&�� 9��[y^: tQ���c)H�~3�^��+��+��x���b����5��n�f�)W�/J��1�{f�)l��J._Y���\�)�ϣ;���?��5\Y�?��Jj��>k��8x�������]Yy7��a��)��]�_�q邾u:�_�������۹�5��^1�~/�#oU�\:�bd�䜼���}e��gd�d�/��0;ʹ��u-��ζį<��-��?rF>W����N'�����f6|�T̘� .^ꇕ�tE���:�c�\�i�V��WfVM��]�P1�Q��g�R3�>u�&��B4�Uyhp����e��y��;����_?l��U�����^�������/��ǩ�:;:���B�^��p;9���7�f,���=�Y*����Co�������F�K��y/{!���.�V�E�':�|�Y�h������e��:���͌U�p���Ȑ�3MK�}7���j)�4�ֹ���:��\�0Iو@@}>U�����If��4&��S�=�.A���kn�]!�"�`3��ί-����H��."D)_��[.3]ֳ��lW�b�^OlR�Sr�I��X�q�p0�<u�����>^�Q������"=�)lm�dh�Av��9��[k}o6�}�k]p�~�6�.������t���^�4�ϢQ���*�q�P8�θwu�V��Z��n��������Ɵ,1��ɪB��nx����m� �O�=���;b�μx���~��Z��
�Q�B���\����j�ޯ&_!�K��M���� c�C��t�@_���#�kX��t޺�&h�'��f_�ʜ��v+F]/�Q�+.{^w��T�~{k���T%:��E:���/�� k�r�hwx���Ck�Ņ���Ŵ�_�ei���lG��To1����=�U�����ո@�y��:�������.�F�+��->���lN�+���W���r�8'{U���){~����c�Y6$O��Ś̯�{������H�}3X�Ύ}�`A.��2}��v�pZU���ln݃�-����W�;/��gR��ҝo���#u��|�OU�62#��/�<���F]�a�[�o^�?)ɳ۳�� t��wvʝO`M^!��J��ySIT�,����Y+�jH3Z�X̽'7:�V�S*Dш�_�
�������&��徦/�2�Q��Y��9��o�nF��sתj#�!\bqc��wz���z�c�̕��Ss8k�l���J O��w�G7��}�b��O��{�i�D�٫���c����G<�������ʡuRcJ�h��a�^��\�{7]�R����T��d!'�g�����W�����T��:�K���鱿�T��`�{\HU-޹���s�j��_{��C�v�q�/��g���y���/L��َ5�PA�0����^���K'��
�l9�ɗ�#�Dv5��qE���	�Θѯ���9�j|�g܅A���{ $VS��ₘ��o8��9���Gr��ڟC�:w�AI͍����\�;^y<#)S�B#��+���Ax��F�E���}���Q^�9҉���V`S��K_W���7��˹|u8�������w<C�������Ԥ!��� tg��#Д�:
���x�����"�-�ݧl���4���J{�qUTa�5jl��J�%q��Kf��1"_Ԣ�
T�����o�QChFr3%���5*��
��m�����y��#Ně�QK��A�{h�[J:������Ѐ�F���^����C�m;��D�]ƺ²F;E�`���q6�Po1��;3u8f�w=�je#q�⤧��5]*�c5՛Iv��wlf_Q!R4��Æ�I��1�����t�N��J-�[%�yE(��v$�]��@|w�c�y��y|7B��Qq�h�x�2��Y�PF���>�sN��N��<�����4�'�FH}q?a��蓜n��so8oVuuj���+L�챫�l!�:��C������x(W���3�Oz�M�4�*�M*[,ݿmx�'.suC��=��cE{r������!����X�5�q"鍿r�=fE�������p��''��F�d�����&�}�	��R���=���7-�Ŋw�[�{���T�?wt�F���0p�|U�.0(��91��0���U�\�tB�4�����
sz��KڌGS�ޮy���i`�ߑÒ���KGO�d�:/�T���(*#f�N���z7X�@K���q̰W�KgnWW�mNq��{sd"_i�/��A����	�wu��t���u�+��Nd�U�k�
�`���,e�-��S��3���ۘ�^��;�a��Z�f�mi�CS��X:1��:+�S.\_��}
��]+��`��ٵ�9l����MҋG'�%W�]}�ܵ��j��n���<i�u�36e��������}��If��8+�ٴ���[��������P}�����ztK��p�(�]�׃�7�����E�H�P7:��ڐqN2')�ⅇ�g1wǆ�d�{�H���XZ�L����0~! to��=�jR*���Ś�����Е<7�Q��@Z^#}v_���C/;�������wc��.}� ]	K��E_��ho���Cu�k�4;s��tf�0�E��;^x�3�|�F{�q�$�A�S(Z
7�nO���}���V�WN�?F*L�:�h���ͺ�e9�`O� ��3J�6H����ˊ��`QoMb��b'�&/w��.Ӟ��7�Des�a �Ie8�D�f}���	�,��!}|��S��a���u�>~�r��WP������ϕ�y���^楒�`c�#^�'��@9|<���j�MXM?�����O�l��T4vov���y,sjjJ� 9nPWR�6��}�=[�]T�ֲ`�������9:e��r��>�����rs:^��|�z�mE���ӝ��S���s��yt+�^D]l0xύ�C#�M�_OJ�t��cU~��ъ�F{b�����뚇�dĭ>���)�ϣ;ߦ����Y��X��6�1rpq��ϛ�vkey���V_	��Q4�_,��Ֆ#�n��2ep�v��A3�t@�X��W����Z��}~;��h׼(>{���]p��lG%/jkCoD�d]]&.oE�oV �_jހ�.�K�M�^�I�6��r�P��2�f���3�_�5�[���/Iǻ,	�[��
#�0S��z����ح>�[��<7y�+�_g�O���C��Y/��Y��p�p��d�/��09W:`۩l�ʞ�Yѷ�1�'ɯa;[�HU�i�l�v���:�Ӫ����]P�-��q���a��]pcv}5�b3��h��b��NT@��$韠�g�:|��Q.Mzv(��UW�����x�2�M�lr�[s��=up���d>��6�GxI=~�`�����[S)C�U%�t愺�/6���[f_��x��lV�d#��^Z"��h3����@G�G3
Eɼ*WΜ�y庭�0�dC�/+�	�N�`�x�q�k��i�FP�����,�@�%G�1�4`���dY����{p�u�GANb��اF�B˽�7>NwI�<u���ǣ�����95���e�o#
߄a>��.Li|^w�O�R޲0W�5H_�sĻ����m���K�Uf§�;�x�K�Q*#��/�;G�eɯ{����y3O��e|�S�I��^�=S�Y9Otda�B;�(?����;��VM|9�d��ζ��n��u�Q�K1�|S�����_	0_�^g��L�*}{���e&�T�{FM���]�3���B�.��i�aD��M���6�tz��uB5�E[���IU�{�oVI�Fw������1����)����e/~0�>���nc��;�M.{^sS����<���nX���J�{%��ɒ��1��ʂ}��$_*���������z|�a�)綘�.�-*����w����e�VW���V�_��K�V���u�kK�k�Y=�>]������>1�b_�K �.�t?���;�5{U���/oֵ��8ϱ�a��j���s'�>W��������~�b:Ϝ\=":,ﳩ 2�K�)�Z�bs̫�47M�F�87��]J�Z��ۗ=qr�s�#�̣vC���M�᯦!2z�J O��;���pW�u>ű��^���;�?E5�����.	�����G�PʈVA��_�_������¬.Y.��v�ј��1Fc��;�k�q�nT�x����n������R�N��؈�w�E��P\�Բ:���<�w�oD�rЧ�*X5nC/�����8��;f8שAg��/�:�~l?Td��fk,es�Y�6n�!�4&����~r�c��sj���b��
�ǯ����������*�M�T@y��n���lFk�-��#�(>�ں�����݄J�g�N�y]����e���s��%v�+O��Ime�ʣ�l�A�t�����zJ�h_ hԎ���P�\�x4<M���3F+��D��*Y�c|q����vw]���r_j� ��{� a<�w���yӽ*u���{\9�<����*|� .�+��Y������<3�ǸAnt���s+3��Ƽ��zk��_�w/��0��>OZ�T;W�zs;����s8"v �� �|\��5���x��xO����Ed�p����U���]i�/�rp�7Xyų�J�Fa#G`���׽=+���0����jg�_t	�������)-�Ĳ�q�hE��(�}����:6'�Q�ȹ@]�����=�{�s s��_5f_l�+�����O��td�_�>F}��ó�D�x\yo�����Q��TE]i�|u�?F�X/+e�ݖ6����N�Eyc��)�`�{�࡮���1y(AV�j�8��a6�{^�}��S�k�����cF�ܱ�r�|mk�����X�*6�'0����urꕒ�>�*c,t�Nנ�/���ATܾ51	�yЙ��T��L��;k>�N���z��~~;A��.��p�Nߋ�>?NñYU���_�ib7�}y	bl<��h�߸�L�E�H�(߻���(�����;�Q�\�^�f+�	ƈ���(a�1��T�;�oe�!n��)��|���7]e�#g&+�ŃA8�ɚ�*˩��F�P�z��i@��ڔ+e�L��*,U-4Fd7�Y�pOg-oT"u����Ԟc����Gm�^�t��0s&���\�Dh�ڗGFH���	r�T���]���&�Y@s��]0k��,��KgnWW�o�s���ۘ�TQ/��kA1O����auWM�á���2��$u�K����z�O�����4�]�Lv�j�=��]æ�q�����ڙr���s�T�]+��`�c�6r��@[I�L~��n�M?[˒�s��g�����c�T�G�Cڗ�����u��n����`z��d��-Ϋ����V~�.���S�~�d�
b#�5%���9�0�W�)��mS�����J߇ӎ&ҽ���P���wN7��P2��Q�Q ���g��(�oL&P�T4�xթ�U��Z����x��N�>�{M.3	�6�ю!��
�1�l�.w�.���ۙ��bC���u��Oz��}, �-�Y4�]�g��>�>��Cc�{1�g�uK�^��^q��"���F�定�r��*0㛪��j�/���|?�������[j����[j�����ڵ���Vڵ��[j�����խ��-m�[o�um�[o���V���Z�V���j�V���j�V���ն�m�j�V�ݫmZ�~V�խ���m�[o���V���ն�m��j֪���j�V��ն�m���m�mm�[o��PVI��@���PZ���@���y�d���Vg���U�HB��B�m@l��h�k6�)h-�J*�l��!kKˎ�$�2*�c[3&Jj��Slb�V�ѻ)L��sZE��m��Ѡmi"үJ�jzhr�$��X���6f��Ͷ���v76���٦�RkV� �me�U*��9=V����$��K��0�.�u���*��]wN)V�\�1P��Rl����� o
����Z2��G����  r�  ��  c  b����Uȇ0ԥ:��ֳ�  ����(Q��P�q��ՊP������.v� �p��)P�avY�5�hm�o  [���ea�*��&,�)�҂a�T��ڔ���@W5R����͌V���^ ��N�͐ݚE�{s�Mc�h:;�惷v��WE����4nv�-�vֶ�����vj-��ɛm-���/AV���5�79ө5W;�UR�r�[�&v-���we�f�����wr���km������!Tx{�P��ےs�S��[�]1�۶]:ls�dleڀ�N�Zsj��MGFˮm����b�l�3w�AG�`�X���h3��룮[��mM�S�����Tqa�ۖ�kV�v�l�C�z�c K�P@�B�]�#���n� "(v�:�9�m�%3i���^ݹ��:�a!��4���u��@��pi:�����H<      ��JRD i�0� � LOhaJT�� L�i��i�&���%IQLC@��M2dh T�A��I�z��C� bbh ���di��     $҈bT&�bd4�j��mSh'��f���C��S�.L.P�ɏ<N!7��cT@*bZd� @5����$$��}G��P��$���$	 $3����
&$�HH@F����?�?�?�g����t=ł@�BB@Qp���RC`��e��
� ��C��]�7޺0O��>��'�Ԓ��I���@��%�G�C�I��k�����T�%  (��uH`�&��o�l}dfŖʒ�jr�J�j���1h�e��A�1n�/pB��y�&b߶̦�f�l�hy�=9�X���[%Z����0�w�SЪ��M�і1#�d�;ڕ�K��@����<9pDV� ҹzT�l��֎k�brçu�T��r�^�ALEe�!�!X���d	�\��Z�t�����f��e�d���kv���e\���n�+ZCNFEZ�������A�$��d�V:�r��l��O[DXu�SEB�avk�r�;ŗ��Q^jYvfJp�ʿ���S�XSR{H�,.f1�s'RYb��Z�0��F����D�ٖ5��/[�{��6�H.��(�Q:���`1a+�J��k��.<+�b(�	�kS9��')c��V+�MZu%튒�h���W&��wx5L0��v]��Pm�4C�-Vc�^�r�B���vq�L�Z����-��fI��܁U�w��������a)1)�=l2��s2��W��
���I���
Ҥ%�fl�C�F+&e���_�	���A[�T[pU��VN\!�/i�7����Ytq_�\�E��c#����!���#�ʉA8s	�	�-G\(S��)A�dS.L���2$m�	�;�;�b��̵H" �e�9p[uK72dy���8�Xf�L��5�oJL��zq:[�+W5���^�t-� ��]\!�u��E0n�˘�[#�ճ�t,y�f0\�m�Ѝ��V�L��J^�dHc������V�o*-�/"q��E���zŻu*=�V��4�	��nM�El�F�D�aGu�R��̫�/�Ե�4�Ϲ�8%&���1��8 ��h��e7k%�u�eK1lR'���2��+U�uB�sh(�2=8\R�[a��$ᗸ���x���[m�0J��J�zHi��Q��a�3a�̐e�&���J�y���2Ob�$H.�*���^07Coc���Y�$�.�]Z��3؆.%H�z+.��M1L���`Ԇ����l
XN�-ʆ�rn��,Ojhh*?��U�Q_9-�(�IV1(��V�r�k�����m'HsM�����&:(F�POV���a��l��0�?X�XW��Tޘ�Wh�m��XL�N¼ض�3,�!WFʷh�	�Y�n�T�+U���/,�.�m��.��W��G���c�S'�=�*7�l�4�+Ga���İ�09qlhe�d��u�n�7$τW
��%\���wab�#�tB��Q������)�Q"朽)���W�3t�J��V�6	��W�����q����ڃ��o˽�XvVŢJ9��ƪ7��le/��#�J��D�n�*^�(��%����*�)+GCj�)����,���ۓ+2�tZcqh�c��v+ >�b^m�tA�[9�Q��t��J}�(v���+4*����#E�X}��R��W�-7�Qi��q�Bn�U��י�(ܭ��A2���d$�K-�ՆL, �ӭ�V��swn���r2j�n}2J"�.��F�L"J���oPk��-�~u ��0Z����b�q٫�t���Ѣ�l��[ ��G�d�ܗ���;�XX�3��R�2!�[ iXPWg(S��M�2}��:/]fVLfA���̀�ʭ
G�$�I녕KA�
�c6ŚXq^�cU�`�R�mF����,�PHe3����7l�wYxCעHwT��ĉ-�!�~׌�{���;�X�e�۬vR�tQo��WI�p��z-24��#6��X�h�Kѳe���ν�tn)�JnH��i-us^͠ʃ��ڎ��kohS��,R��f^�˘,�Ԅ�q��C7��t\pK���#u��0CX޺9
`����1lA���h!u=��- դ�6pC(�Q(i]i3��kBX���HU���̣�جp@��(��T"�ʭ���M�[�n�r;X(PS+n�	��� �(�n�pP�3~2�K4Tj�ʼ'�ße�]���x٫�֑�+7)�dB�J<��6]Z6��\ݻN�!5Xd�԰�t��bf�sU�DK�J����Ʈ�/�hp/��z���n�_ Z1Z��d�(�p\M�9��2�8v���K;	-)y���Z��+f��f�Y�:zug��ݣ�S�L���+G�����e�|dM�$r� ��
˗�%��
ʵ��7n�VM�YDD�hj�c�����������.a�L��nbZ��k\��z7�,	��&ɹfM�ת��1��Zx�ZAg0cH]GLU�r�TF��+-��b��ߦ	5�f�n��8	7d�S��'k�Aѳ�
۹%H��j���!J�+haAfb����9Nη�'n��A�ugtX�7�B�K37���ed���M"އ���9��
[V3w
��mh��J�,n���wp�*��/\�	�d�����j��4�^�Ac"n´4V�>���@�e��u��#�������w7��nMRK�VZߞ}�l�rQ�-n��KO])����6-E��AZ� �ϖ`�ۚ۳5��-�pA5,�us(�֪��!f����2�{be�,�k���SIV��;��]�ME�ͽZ��4&�_)��� EZ5�:Y��-v&�3RKF�k.�L��N���^���Zc�g،q����iE�YO��տ��QyHX;q�d�3b�Z��m��ˬ,gۑ�ɻ�Hh��2T0ִ���[4D�.ͺ�$e,�2�L�kЬ�I��p��`V8�V<�m��Y���1�#�k	s:�ʎ&���2��dk����naUVa��+]83u�����+6�v���c��cY�g6� ��Λn��%w,?��"Vf|A�zs.��8H��U�d�m�#�b�Yuȼ�p� M[�m���7f�I�D�� ��EQ6][��&;��wNY���1�T\M���"�㼶J�Ĝ�R�E�ɤ��٧�R���L!�8q�я�0f.��8�B7�1�n� 3��J6X-c�}e�T��Q�Y���S����I8.�_j���3jj�1-l�L��X0�׎%[���,�l�++�h�l�F�%|��X�M�������[f��L8&�5�ѷ�w(Y�!�*ٻkn,e���;��yn2��,�
��l{�lF����U�ϓ��y�Tm�������3����p�9w֑}�{�څv��km0:�{�l����EQ��i�1h0H�Z
��0rè����2UՌ�W[3�2�iEs&�3s�"�ɹ�5D<
�.Y�)���L�ۉ��-�[�]���I6�0e�hb�����~{4#���q��Ŋ��ʽh�c�n��`�2P�1v�\�ۤ�����$'[����N�Ih��ߖ��d�VLV�^�Ce�M�cD�P��O,�s&�L�b	��氧�C)駈$�vG8��e�/(S���]�P��]��V�w��!�l�b�ޡ|�\r�J�cn�m�2v㊂�J��ZK:�f@�ϥ�̣'��l��5n�ǇeL��7&*�g;�^W�`Zᖮ7��z'aT���,+NVĶ�ٸ��l���-�����P������la���hsp0��u�5(o�a��!#+�.�����J�=�ۙ��J��F1k2m�J;��c�2���aS�F�ͣX�[.f�j��6��yr���l��р-��T�^���Ԥ30ʴ��MؖZ���F�Ũ��`���-��Sm]e�u1g+cԍ^�T�]˕�bё����`l+T�Vi�)U{b1*A6�{���tbZ��5��5`��u��Լ�ui�l�K�މK6�5RYQ�ڨ��+�->ԗ=��ͦ�H�X�����n-��3OD��т]��,S3(J'i�a���ܖ!kv:/2��\s�i�(��fB��
ں��S��M�� �䥰[��H�қ���˶H�E��T^��R��n��[ۣˣ��3���I�?������R�����]K<�Fb}�}��|=Q �[�i������q�?��=Ml�.�[��\�=�\ر�@���7���[�<��Vu]oet��
�(Aj���r�
�;aTѺ�s������k�"[�;b��3�ꝺ7���憯�2rxɘ�]nv}�i�-;��X�]�2g��~��U��w�ɭ��gZC$����se����mJ��� 	��aBH�:����sq���#�	]u�e�'}�RF�Ts�$H��i�tG���qU�J���~�����)976J#(��f�%l�	g}�)����b��[�#�a��u|������壞�M�35m�%�����p�p�Z��F�9�I�G-�3Da�szye��B����ΫC���isxb�fe�K��Pl{l:�V�fÌQ��>|q�2d/j>om7�]������So>��T�ꌋ�G]��٦�IY�g�^|��h(���pÒe[Sd�r�w2�g�;iW��7nm.㕡o9ݸ�o�-������Ypn֡
�t�,�aD��Q�M�#F��{�vp!j���e�>�{��4Mp�ªZQ��U�y@�Z����,{Z9ky��GAd̼�S7�:X�&�M���OFu^�*��{��t1�\R#���J����w�iqP@�c��;`�b�U��� ��m�x�f)1S˙��gf�����z{�e��B�4�,W]%A�gm.��k>��+��K�
���wrʲ(M�fW��l�Vҙ*�ʱ�
]���A{�q����8��Z����0�V�p�0UY�Gh��;���S���;��q�X���/�G �rulT�w�-��f����G��ȭ�*����VG���Ғ��y�D���Ω=��*��ùD��pl޽���e�������P�ڡi���[����.��!��7KR[�n�8��������M��K\��/�o�h���{�5��A1[\ �A+�j�9/S2�@��*vW�VSRu۳�ߧ�76Y��YdZy&�f�`mGΜ³�s�8ݱ�O��]&y�oE��p�`�Y4��JS
��ż�*������\31���b��IN�����v����B�q�u���&a��J��],�F�nu!�
�gf���Z"WQ9��]��(d�:�]�D����Bo*�.P	uB��e��R沧��ڹ�a�B#�\ʆ�5�7pd�J*3�Z���]�׷�%�γ����$;����L��af=�n����{ �O����cx�[�Y�b�s++��yr��:;Wk�$��S��o] �m*'	��8�=�0���{���Gz2yfKp��ح}(��Y�2�#��������2XF�I�� [y[�^Ӌ��ê�W>+E�E�Eg��X�M,��y���T�����=6|酜��ع��ō.%����.��
��%���Y��k[���.��)q-�d�j�7�e�#sj1�4��즆�����k-q�~d�9���'��)aY{��5.����u
!oV�R�s�_s�[�!9��@��]}��4�������y;+.��pWXo蘳9oN�����p�ɼ�# ��(��%Vs�
��Awc'�OR0�K�n5��k0dͺ���D�I%�Vu)`��a���0<��y�&'F�F\�����Zʔ��g��dЬ(�N;��Mm�+�h�Bbtw���P"���F�[擋!u�wM|��!�M�T��[n��9Y�Q��4ê-��&��f�&�{,k���4ocK7P��41Eq+;�=o̠{ލc9S:�)ڻ�C����1@l�y|q3��K�S�c�i{�em5*�Yt���:��6�,���s��L��} �/��y�JE���fA�u�:���4�^X�b�xR�$�
� E%rۜ;]���	���KGeq��D0S�(WV�U���TE�G`��Q��{ ��Y��"��rq_0�;��9���)�^����{���r�;�o�1��Z+ ���^��GX���a ����kj���d�.��]� ��һ(3�;�*�@BG>���Ė�[��(.�ȸ���̧P��ٕ^����-++�(XnM��lI�'�)��ܩ�~#Ocʄ|s8����:3t�c�֩����X׋fW\JM���o/�W��WXz�SqM�K%xz�}�%��Q�=�v|���fI�쮽R�	[�佛�F�٬�2o2��9�m܋�:��\�*���-^Lڑֲ�|�*�r��L�c��Wu�B�j�5c\	��oM�'U,r�G��� �m��t�<%>�c�h����Z�=�:Yi�f�8$�Y	L��L#������^�U%�)@� �n:���r7Sb����
B[նMg+r�H=����}���
R�lwS%�'0���u���M��,�w��jq���ʵ�Ԫw���O�4mTH>)��KyW�g\p��.�֮�)`ba�$_�ǖ��u�I@qH\�Nfڧh�er�$`�h*f���r����3F���+���0Y�ٔ2D��عr�ۡpffΝ�4�:�/6��Fۏz�n��@d���/���V®��Q��Z�Kuر�X�iab���
��;�����)��c�n.;����l~L]��!I��0z�SJ��Xy|��Gn��u�A�s��˂T`V�z��0S��v
Y�h����] ޕ��4�˲\�-�����O
`n�!^�4ʷ~L E*p�f��+݃���ݜ��uO�컶m���B���:�tE<�0��mue!���x�#��vT��6j��@m���S:,��t"���Gs�J��:<V3����CH�krc��ݯߥ�]��:Ź�.�W6�n�����M���$�ܭ|1�O����:��p�nZ��I������;����uqQ��X����p�6Z������[i�ۣ
�m��s������8t�,�r�F�;뉸�����T�]wQ��AC�#�5���L!��T371��\�	���y�6�;�Ԣ�p$if���Y�g��h��L����P��\�0��`��v���U�b�P�I�E1����o5�m,�j�K��} �}3[u&w-k
��n���\TnD��q�uȃU��{|#޺������N�楥T]�Ai�A��b{��ֳ�T�y��ڶ�n�;�Zч�W-����1�
7U�I��®����s�u&c�֛-�K�]b�l��)-cu>�J�`���"�S�ثʾ{Ϻ��#�6�U�vr��[��!�QY��ޙx@\�+�.�Fm���pX�['s�j�,���\�K����+E�6�rCkv��Q*��G�J�U�
Q�U����̖�p3b�Y7fpy�X�����Ew���j�ii���~��[ݡ+��ٖ[#�j��&^sC&V�)d����w�9�V��oG���[��Q]k�Ҋ�\�L�Y�s+�X�?&����	�^��q����Ds��� �Yf�LZ��',NC�0��9N,ߍV]*�������E8;<��M<`��wtQ��(�r\��S|��Q��� <ݻ�|0�1��H�����y*]J$|h��]�i8���I$�I$�I$�I$�I$�I$�I$�A��b�{q�� ;�'�bK7���+�%��ݽǋ���i����/^�ә�V���l��][z"��u�1m��8Eے[��ik�0���N���7�ݻ��-����U4�r[���E�5��bk�5�
��z�
��;0��*^��\���l����ɍD͢�Dn�1j�z��ދ诜�L�OsOeKTN`��$;���Y��@�a��P�Ml!��s�ܠ��T�au\{/:��iJ#��Z���cL�&T�6�o��銒�����Pʗ��[1��N�;Uy̷���{��m����{�'/J�d\Y8��"��X��n���vT���ulJ\9�z�gK4���)�NY�EF�����w$��,�5<��ʘ��]:�I��ce�ۆ��7Q�eE>�QQ�F�I8���&ޞ�����z���p�|��.�<o`ˍ��EԦ
u��ǆs{�����>�������|��^|X� 	$$�	�q��@�����C��+T�?a&BB@>���߭�ϖqs��X�=|���X$�HS��mf\��TN��*���6�� c�@.cl.�G6-v��MvT$����|�*�^�B
	�m�(���᳍B��"�e�&�����Kh�G�(����{{���6e��*�nm�
��M�8;�N�m\���
�\����V�5�hǹ�6C{
�(�s')�{cC�ͫXJmi��B�-7v�����P�9Ty��c[�L,�GB:�Y��[c�B���X�=���/��d]�3��o^b35m�.���wT��j2()k��A�s/0�Aς�A<5kie�Xw�k����rzC �uj�N�%�a]��X-�>۲9_�KW��U��z�ǘ�W+!�qf�z�!�G-�;�Qz�{���5W�1�q[v������ �uE?�N������)�J!+�D��T��٨�/���Q��.�c�����$���9�s��Mp�F_
7���L�uځ�[sUe�w��Y[B�6n-�ئ,Y5bF��o���K/5֭�5�u1��MK�ڹt�7���&��|n�r�s�Mz�g,�O��ξV4�[h�1�˕h&ZB])u�y�fV7!]�sJ�j5l�|�.;|Q��dSu�o�:�г���#��@vS;��}�K���P�9�ٝ���d�F�,�B�w��5���xFȭ����)�j�"LhD�^֮�6帪0/�2$��q��TO,�#�2a���R8��zl��	3Z��q+��F�h4^b�e����&����a[U��SugP���=tU�j���O���1�%�7Gm3�T�ʆ�o*����F��V��Y�3Xv=�w4�-�R��f쮡X�-ˆI�Z�)��-�h+1n0AYD�T(�}���!����T
��5̋a%���X�W(������Z%W����D�ڬ�I*X/����Tfq�%�˦��2����Bɏ$ŷG`|�q���<6�'\VS$��7iգ:\�(S���'�v*�v�w��Љ0�Ew�G�@Φ]���޺�W�ՠ#֗-ٔ�}bSO�9�q��Z8�B�Շ�����*�3"�|*e.w�����m K�0�+�|�	ܢ�K��]ۈ_uwk5��1�Y䤱�sK���ϝ��*��L�{��Si�LT��t#7M޳�iǎ�T:����=��$�K	f�h��n�f9�z���❹gk��N֊Z���
b���L��'BmR=Ϊb=�U�/���ѻfbG�@]�|n�k3*�!�RTn�9o���rp:rźB�_cC��e�Y]��L�ڒQ N�Sf�jSo+� ��T)=��.�wmch��a�o���70&�1B>T��6��"!��ɽ����T~#�3�Bƴ8f��RR��s��EVm��:�¤��\�֚%em���9�ŅE��(�/9^�3����-\���o��3��h���	��H��r����b�:�MM�o�`��?]^�Qu�Cm�A;�)Vu뛽����B q��V���棓8)ϋf�\̈́͞�2a�\��MV�e�MB/�j9k�I��lQL�]勖�\�n�n:��o�ө��7z�n�)`u�]�u�4�6��Ĳ�\�M�@+ͷmٌ�6�A�f�j����37A;���}#�xT�(^���0ٸ��Skmj��X����җ�Fk)�X�leR�9O�y>N��F���̔۴�y�G"�HӒ�/�7ǜ�N��(��Irؤ͗�9al'Z+5()�)xNj�j!N0A1؝36\/�*���6���R���b45�I7י�x�^��Z�-���\6��U���,����Y�dB�%�c�o"�L.'�����v.6�ޫ�p�@�>�ˤ���QYjY��]^$��M����+n���-�[[��������Ո�ڰ��O2$ޝ�K�5�Z Qy���:��� �e����޽��� ���g��M�
#e&��5t�y�����e%�R�hS�tq�w�.[�*(��Xp���,b#{v�U-��o�ZAEh*i'X~�U�O�2�6�7RL핊�+^�ʛ��r��Tʷ�:�j��e,;`�j�����j�uu���]<af�)o,��5"�VXWy�fݔ4��f�WI�THB4*�^����$r�T�R%����xp����@~��#	�Bc,�yr��B���B���=��[��Z�3z��˻�¸t7�C�6�-���MH����μj�Сc�)�$wq��ͪ�^�r[t�V]h��<�1�3�i�[x-�hsS�>��9�/��Kq*��Y.e�
�RQjپ�'l6u�7S�ʸš��(J]��I�Fȳ琌�o1��^1��n%2�f'J��6�rt7�ųs�j[��FU�V�X:֭�<(� ��*Ρ�] X������Y�r�@ۼ{4�BE7$�Q]�B�������8������\�kB���Q�}\&�N�\��٬���|В��qt_r銰�����=��PV�n�駋\�jai9�*r�B�B��j��
H�[F�P�3�S�;\���zY�{�K������hYuj��Fl�I�E�u$���UG��"���ٛ(9h2H��grޣҐt2	�J�Tz��Yx͢Q�ht�΍G\�t&���ӛD>O��̩u���:Zw1�a�Ü���\;��M=fE��f<5��O�r��6-�"L�g�qTk�X�(ݘK5y��c3$l�1�-�"�CY*4��;���Z�>J�,Lж��[5��6jZEIiY���q+߲�kv���1I�W�{-�th�K�v��1G&��8�'����ۢN#	 �ʣ��tM�a>v][=��fpڼ5�b�F�\0.YA:����8�޷N;��љ��i墴,���	�_A��"�UԐ�ՙ����4�8��R�_W�f�H!�ܪ�g�G�cz������u�:�/3��O��-0Y0ć�,�@����K��`�\���f=Z.�]|�J��r�N�󷺅r��v ��Z��F�毖���7wp/�Ѳ�h�Cݶ�IB�e���n�vE���ۉr���yG�go!�l�J$5۽��Fm���̌-�h0��U���C;�پ8,��I��˼Ko͒*4L�TNM9Z~�N�V�����mixqL�*Z�ٓ:F�4�N��Wa�(A
��n�Ѓ)��%Յ��v� S�ٮ�]볍mr���;:;F&�
׻�a��G�X���y���v�l�R��+[7a�ó3)��Y��p���F��8��w��z˷��Q�yLÃ&ue.�vT\�|U��.��E����y!aͨ�7Qʉ�O�oۇ�|�X�)&�Q����!#�2VDsE�j�.��!,V�;�oB�(ؖU�k��ME�@�P�ӯv�}�R�1�n�.I�NV�ߏYu����)�Ȼ�Q'�Ka'{���N��Iw������0��[	�CL�I̬�J��jJ�jn�u']���
�S&����T�u3s6ު�P[��X$;���6���r�K[K����VV�2e�!�]؄�v�����k����F��aB�u-��7Qϳ�	.��dg.A`��+f'M� �T'��ӯ��D�e=�uݖ�V71���o���TY��}L�n���Q�ګ1�쌆��*tW�&k3
W�[�a����ewܫ�ֻ.�a6�v�fs뾮퇸��X�u#��"s��x���o/�,��A](���@�7ʻv�J�w T�������gQ�2_<vR�mQF�����N,3�]�]2*�R���w����bқ��")�زpjX'H���7�l����7Yx�  U��U�J�9).�D!Uٻ��N�#o40[�B����6õ���7om�t���Q��bx&}yg�7�*V��"�����z�k̼"�ƹ;�qA�傶]�$C<� f�Y�lr�����9o�[w���q�z�b���� �)"���B���o�,}�_|*���{��kGY�N�=��%n��;�S��r%��\!�%��A/�����)����L���诱�X]�V��*bB���w�v�O~w/ɓ-*�����U�V���;RIEw��oS�ZnoM��9�"G<��]F�S�"�8e��oc'���e���_nE�R`vT���0�m���ƶ��}��o
��4i��� �E̊G�#����g�́���%L�ϰ"95�����lޥ+l�Nr|���{5�J6ek�����Ů�Ρ����s��aޠ��_>A#H�ʄΥ�io/��Z�}���-���;�p����=�����V!an��A7�oZ�)=������-֮X���kzr(bJʢ�گ�t�,E
�)/.�gV��&�;}���'����7k������~�@
 
�"*����F%��Yh���UA���=��E+�Pp6�m��TډT�T+Q[Ymj�qK���4�V��ѝ8�Kl��ѵ*4�:acmK�p�\\+�-��kkJ"��1����iD*Q��ڪZ[K-�Dm�Z�-JZ�\8��qij��EF���eԶ֖�
�T�j9��h��նV��Ң�[Z�6��E�E�j�[�Y�UU���3�-#,T+mmTP��l��[���^���7c�]t~��v�>v6.�EoI������G
v{ؑO���{�J?�����x�ǳܬ����s�}_���<��!������ByN�]ojtE�׽��Z�p�[v�
���3�r��׶3�Q{��0F�s�z���`q�.A�fd�2TNb���/G;XjnP��C1��V�
�ə�b����Sޤ<�L;�x��c3���R߆����/�2ט�E�SY`R��t	5��\��b��(�M�WwZ/����Vz�%[̼���#`�9�'u.�j�3nɝ=!�܃}�cC9�#�̝?��ɾ���/���Cz�r�x�,��z�Vm6v�aV�x�fk�i�z���`g� ;K�ҁ+d<]"j�==KzH��I�b�B*�i@�JH$3����uA�wZ�5o�1�ɞ���(��&�۬�9�%e�����Nj�|�ma;��S�,�]*OjЀ�p�t���-����ĎFGѻ@W;t��m_�]��/�w�zk���[g�r�2�+�{�fo��<�흠.G�mD��y�_���C7��+lg���Me�C�t�<����0ܿ�5��j���"x`{d�pk�B�~�����5�z�@��>y���:l�G�b�ʭG�B�rO����'֔+�2x;� �0c&��"\U 6f]x�=7{�{4�,������f�b��ې�Z*%�m��&P̠�|+R�Y܌�C&���(�]���f-Ǉug��y����c6T�V_w�\��#�����ԅ6�N#^����cZxO^���5����)
͸5<��їC��M,h���^�=�g�zM���K��5������owaB1>|(ŅN�i
����F�rþ��"5izd�ǽe<���}��}�&ƙKj�x�����qi}i�`R�V�^oE:��Wz�\��F�է�#+ZJA���%���+.��'�}�W���y��n�w��z��ҷˢ�-+G��V5�v�^>��J������5]qb�˸�Y�4G�)j�����q{{:��"����juW�JҐ�2N�ӥ�F!z�z~����o�}�u�d���D=ƲRN�����6)O]��M��fD��q�XT�&(�]^��i�o�;z �^��v�Ά4�!���o���N�y^��랗,cܫ^|"���N͹�46�����OIY	�z�X��e��z�;"c�v�^�튞�y��V�m����x�/9Z��8֗��K�gF�HZ���c��苞|�g���^#�ZN��������6[���:Q�qN�Ӝ~5���	��{�B�N���ܐ������z57�.W�ނuykM��BVoNz�\�\iͧե�Tɀ�@N����}9��������~�3���1l����/vi2ߧ�,����N��FG���t��y��~|�@����߸`�����#2������anv��k�^�P��r�pA������o|���gi�G�����׮$ž5/;�_VlW:��W,���mzsq��ԁ�瞀[À�e�®7e?q|�3��T1(!�|�>��g9���i{Kٝ�ϩ�����+8�ܷ��!D]���o�I�W����a���,yS���P���v�c�tZ��t��n��t����;���r d�%o�{ͨs�-E0�$M�M.�e8s��E_*�A����2��� �r��]��H^u�r[�kc��߻	��\�Ș�V�{3߿h��%�Ӈv����7���6R�ޥ�e�>�^.��#�S���:Z�<v���%�lQ�x�v��Ǟ���zTat�w��᣼�ƭj߸��spz�-�̈́O�tZׅ���Պ�Y���P$qB��OK�׶���f{x�=�4IY��y>\��J��s�b�lQJߦ&�U�ӨÂ<}�x݈ۡd��Q�O�P/���JW��N��Զ|���ݬN4�0���=:�JS�������(굤�����̫�7�'PZ�h`�t�j[��$uhɶs%)t�r=8�SOǣ�f�YfJ>���zC~]��]�˲�頗����ƣL�95��j�	�z����Eշ�6|�I�����YX�k�����x�m�v��Z����B"��;ҳ��&��μ��\����r�W��y��q����E�Z}Yf�ƺ��8��¯�X�dm��C<����h����9x�R�o�w3��u랣�s��s$�b#}2�L���e��<�.�y���*�H�&ϟA`d���~��1�4�|���ب4Mv�M�'�&8�k�󷷷w�x�
े:K
�Zx���Ĺ��e��ܨ�uZ�V���r���7OY"7��S�X�Sr�t!�LĹL�(�����x��U�L1S�f�eWg�'/�\E�f���xg��*o��}�����J���aN�է|��)wkIB�*��U��q�2�u�db���tZ(�=�)�E����y;(1^oI�R��oV�Es��!�h�=s}����LT�6F�#����3�WϚ̮X;��O�xwg�rv*�JƯ��K�Ԩ�ٕζ;0f�jg��P.�GF�V�yY��'��Y����<U�kR��� ����w���ׄ�Yu�� q���P
�Ύ�	m�DN��vSM�	����|�����+��E�ݰ����m�qk)F����6�t�����Ynv�M�M6�G���	��8Pw��;�]�e;U��ޖ}�f�������zan16V	=���E	���ӹߍ�ߗ>rBUb�\�OZ��2j�e?^6�i� {ӧX��fҕ�,�}x5nk�ߧj֘Z�i���4�:�`p�4��g7L~�����[:��W��L�Y��=ν�{\���`���=�+�ﳐ�{��۞Rw����b���H���V�$�xw�S���֛8s;&����Y��-T����U��q�����9��;�q:�fY��%���PomN3��J��;n��&��=ܱj9$z4Sz�␹}�'5mב�=��V�^�,I��L(WrA���G���|冣��^��iJBJa*9\�gƦ��E�g�%�Q�8�a� �B��Ux����E����)�]���=�-�j��RYĤ����~�z��7x8�����0��ص��j�^���tV>�>#5��'E����{Z����:T�:<��e��ZoJLo����h��Z��[��7}1���$Y݆{ر��������!��O�gVh�	2����q��o)iعH�&�-��\�\y{�1.�����+�4� smAbmK9ښ0(Qv�)�{��.��q�f�\�P�9Aj�zQe�k%��4I�������j�i��f���ǃ�!h���˾��Z)��V�M�Q�q0k��بv�,��z��xg9W��L'�l
:H��Y�PYP=�z6�������3�-f^cT��f�������t�fkY�!u���}Ϟ�[v����֪毢��S��̻m[b�殸a����k���<B	�Ft�]4ڡj�m�y`{�$����MԐޗ���=Y&�{��E7tv�f[�.����94��K���kOKc'��c�u/��{�ᬌ�y>���+��ww�7q��,���U�����9�p�d�Z�ʎ�5�gW�w�-n�Q��% ��o=�Ėo�^7����x,~�_}����Wq�����c?os�Tˮ3P�fE��>��n�{+��-��+�|B������o�*�����f��>Pd���ʵ��t���
�WI���������mJ|J��|v���<��8���t]�v{���K��3�!���aV��^�u9�=/c�N�v��cS:�Kݡ5.�VS���`�O��Hu�+�t�*]�)X�yX �d��Jū=w�(JC�$&n�`ޚ"A�:�zQ�xѩs)
�u%�F:��<\��u�/��6���]��l�t�-P4B�٩NR�W��"�v���yZ#���q�IF�aJK�*�v���.s����mR�	�:�=q�u��Y��)�N��֮�;M�kzujW�n��o��T��r�l_!��B�o�,�om���-�C�L�����˞�wV1�ZXV�+F����Ŵ�V�V�hVET���e���#[VPr�0��m�W+J-[|�1j�m��Z�6,��-ԭ�T�D���(�J�����Z���V*���Z�J�ѭ��֔�B؋G-0+

єk\\b�ѵ����h��a�l��[jR���-��F�Z�����-����U�U�D*5-B������Em
6���b��h��FڲѨ#J�ZZ-�V"��[��+F�\�`qmhTJR����D)Z�c�%��UeF�(�[֪�\V��iZV�Ÿ�KҋcPVԣf1p5��,�֪�V[j�kj���)\Q�*�����1 ��E�K8V{��Ѹ�������ޙW�,vh�Kh/Bptrm4�S�p`��r.����vxVg.�|A$�kc��m�.����������䶣����p��6=\:P�`�����t��m�/l�j���S�\/z}1����u���������(�u!��ג�e��L���D\	�Σ�;d
��;<�zw![ysޟ.�j��x$Q����.ǌ{늒=
�N˕Dd1�B��Hґ��o���v���Sc؞O4�y
�PP��4�s�g�������h�ȴw���r�j�+�G`��g����\,��Yw��^vaVH�!ǴomS����뽰C���t�w�h�B�V.i�De޾��Mh�1��p��F��9U�0��㒀�Փ�j�k_�1�7��B�&��Pv5��ٿ7���;y/��a������Qn��{bx!�󥏁��iVM[u�oI��sȼ��^���W!<M�p���O�׸���'q�)�ݷ/.����\g��+��U]�ӣ��Т�H���W�6\��~ޢ��8�Ԧ��d{�(.�m�5O%�5��(&U���>=}
����Ms��$�9x��,�wS�w��ι��=\�I+v�u��;��*�K�$�_�"��f��g3���lK<L�B������3eq~F�%�{�~���\���
:"�\�1��qks�٢�II���n���F�b�l'eU�������2����L�����W��j�y��̘��5Q�+؏Z~��{�1c<�%��⢏�ӨXp�ýk&ˡ�[H!}F0�w�^bEK8��[�h�������8��1l1����W���m�����Rs�նƓ1���[�cx���Q���ꧻJQ\����b����.��`��9����yT�;#*��N����Vݡ�����5Y��i�Wn�;q�h���g5��C��kh�!˵�=���qr�ɬ�m��3^���*�}M��\�t��y�]��w����=?*�l�b5�KS�+B�Vy%��v\�!��yF�O�4vSO)𥆕'Z���R�]�c��1�w�4��Z�Uhi��6f�i���-����W5��i����1ɧ[P	�v�٧�F���k']��GON��>�x��ײ�e�¯��]�ۥ��a�c�`X1|w<閫;�s�³~�{�ս��lt���]j�~���Pw�$Y=���C���L�&he� \s���������C���AL�OY�3�!���
M�m$:ݒ�d��z�ܶI2��j��1yֵ�N7a���02�Bu�$�P�)6�1<��!��I��8ɧ�&�<H��^��5���{��'OlB�q�v̞�Be;f]�2s�$�P�e�yM0&�d�N�d���P�q��#��~�2��:;�����un��=�&'0u�}�V���)�V�/:��R�I�t|^��E�ڷ�+mf30���v���(�7 ��)#��C�Rx�����m�������6d4��'hq	�@��Xa�e��d�$�:u�y}�]��y�M2a��,$���I�MRz�I�'I��$=d������:�Л`)��	�N0�ɽ��{��M�B&Y6��T�$�&Y4�z�bHvȡ<C�C)��:Ci���&P�@gG����w����	�N0�t����&�y5`q$�q퓸��$��!;Hf�� ��&�
i�i�]u�4^��7�}����Cl��O6�L��4�Ô�� gVo�&C�`l��I��'��d4×��Ƴ�u�=ǽ����0=��&7d�$�P�'�L��=d��2C��$�&|�m�	��I�q	���i�1�9�֜�qߺ߼��C�,�
�m�m$�JI�M�}��@��z�P�I�$8�v��8b��o�uמy�;��Ni4��C��	�,��i��(C��jI�e��	� ���!��k����x���a6���i�a*�N��$�<�	yM0��)'4���'����xf�/L�6�����s���=0�i��C�4�il
�m�2Cl����v�v�d�ݲi�l��d��O��^w_��Np���_�������`�I�}5�c�#�픉{��������������_fLܔ5v��T�Qbh��k����ٶ��q�R}޽<ܪ�}�����
��t�)�rɶI���Ƭ6�m�� �L2��$�VJ�t�,��@��μ�2s�s�����i&ӞP�2͙zH<�6�e�$�Xtj��6��C�l$�� ��B���u���1��^�I\��v�m��!�)�'��y��	�=�:fY�w�&�%LN��!�he���o^{�����=�M�c�bJ��<a2����� �g�$.)�z�m'��d5��	:C�=d�y�Wx�;��9�xzv�Yr�Xm��N�2q����C��I��,'�� v��~Ra1�${d�2�u���G�>�y����݆L��T�'�&f�Y=zI�`t�y�I���8�)'���d�%OY!��ٷ�y����P�!��B{�	�OPϖH�t�'�O]$��j$�o�q��E��;͐�`ry���Xӏ{��8p!�2��I��6�:I�0y� q3L�L;�d��	׶I��	� ��{�u�1�Ͻ��vzJ�v�MRL00Zv�m3��B�,4�XI�2i���2qY�!�L��6�"s�y�^s|�:Mr����IN�P�6�d�d�'�a�OY2z��! ��>���g��?RۿU~��Μ^����YP{4Z���$�%��m���R��>����7偿����c��] {iL����<cQn�X(I��2D���y�������I>:�L0�$�1�q$1ݜB�4�%���1l���L�ɄC���H(m$����Z�]x{���u������x�XM>��3,�A�X��N٤*����0�6���$�<��<�Ƴn7�}ִp0ɗi a�f,��{d�8�m�Y:�I�1<�$�<�,��@�2i7�]s�u�����[8IY2������23�I��+$:�M�2�a<Bi�v������ֳ�<��·���|�x��x�XN2t�=3a8��VI8�wH/hLR�`���Iؕ�3��6� dϞw�~�<1��[߰��,��VE���Ⓣ&ٝRCW)&��!�ή�Jʆ=�C��!����u�s�޹�6r
�� ���Ԭ!�vJ�5�x�d��BzOY2a�@�,��L�^0��y�\߽���m$��Ӧǖ��!�d��N�7�/T>XN�2L<N2B�I�I=�=��n9��瞜	�!��e�)6�x�X!��I�M�t�8�MܲM�i�I6����6������η���^�G�:a8�):�v���wH���0�ٶ�w<�8�ǉ&RO7d����Z���O?�B*i~+[�C�Cz�ޖ��^Gf&W���w7��H]��.�3u���*.3�����S��츥K��m�Ԭ7m��o����|`A�7���8|!:`(a$�*|NY!qC�Cl�=�v���{��0��������&�L�O4�Ǵ$����W�=��ךֵ��"�\Y�i�6��,$���� d��i��3a;a���0��8���'�۝s]�|u�����d�~9�C�v�	�C')&��6���L��``͇�8ɤ;Ha��{��7�z�߾{��n�&�{7`m���I�Ēw����)Pr��`fݲ8���3a���O:�\�x�n{����6��2!9�q�0y@��	�WL�l&�N�޳�!�E��!�6��[$톙�y��g�{�p�@d�!�2xɧ�;IqN��M2u3`m$Ƭ'i�L����N�HT�������]����0�z�,�� L�Xm���� v�n��>s}�����oĘ�ʝ�Җ���c[Xʝp����6J�&��_΁s�W�.�},��J��%���"��4oQ�yu~��9�1xx���Z��a]���c��o�N�<[{X8w?��JtzU���e�,��2�;�ʺ�PT8hr���݇՗Ϛ������4�?���{�j�Gܭa����A���D����Ǆ!h���	^���7���k��g&<L�7���v׹�0�Y�Զ�#!�9��]���nܵ��xWl�+��nӲ�<n�Ǆ����~r�Uߦ�o��7A�]m�M��� ������K�%�g��ާ1�/�Eu72��s� 5���<KuF#������W���j�^V6�n!���-�&p�s��^yC�n���b����P���<�'0����2�O����WQ:���&�dݏ���6���KثaI%�R�}�Ս��⟍pN��=� �|���)�.e�s�.�}w�V�F�NO��y�>���[b��l�m��R�@a�qd�P�G�
��_���Q�W�B��o�w״�BS?�ϿX�ߧ�\�����u��I�<m^����wr
��O�i��*]Po+Fc�1;I��>��T�LY\���D��s�{�w�!��9����z2Oa"z{��e.&�E������.�J�^j�1������˙����;���r�8�	�<2��:wF������hP#��sj䵯]�%�����_����o���~f���V���/P@�f�i$��w1R�Ut˄)Pr��Z�t��)*4d�"��V+��p5'|��7�EWۗm;Q�WVf-[O�[�8Y������_T+m��c�F�2�TLƷ�m&&����(L.Z�{�.��/:����(
�T��@�]ppו�o nF=gT�/E��|O��v��ʛ6J��Pf]�䀶^���VY�u��+0���L\���47���˫�8�AM̬�++��+�cR���J��'�Cgp�cxd���[��+rK��W�P��;�NWX|�M����%E1 ��mEK� ���{�sn�-��V�/o���\�s3r�u<��Y��J�Mn�m�U��H E��g+;���%f7Q2zl/QpD4s.���T*!��fe_^��Ԗu�k�th��j5����Pemč�^��K@ˈ��ؽ�X�悡�J�]ձ����Y*�����W�r�Ή볓1w�UX���=��M(.<��ԛ��5��f����O�J��(i�@��W�7\%�1�y�m��D�t*u�"	�݋vVm��N�Ow�J�nvJ}���F�^6�D�3�h�o-τ,Aw��8�K4Ru�o�N��kWʏ#Ħ�U���ggC���$K�N��ɸ�׽���eW4E��q�o-��@V�����Tu#L+y����s��R++:^H8�}�Ja�����h[��u�*�6AŚ�6�2�2нofT̓^n ����+�}���]��#{����`�$r�(s��_kC�m�>g�C�Mr��������������fWi��£�5LT��b�F�E���$������]�s� �+�;���(tCv)�ӥ��W����8�u�BKUS��	����z-`�[-DaX#[l)ZV-b�թE�J-�U6VaEV��ҵ�R�֭m��+R�8QEŭE%�a�+ �DT)�X.-�,��)J�UP[mA��EF���+j��mQ����B�b1��b8
�D���j��+���1(��*��5����	�-��J�B�1e[�a+�
�b��V�\Z3֪a.[Pl�1G�1�T0�p�b��*U���0����T�mL��Kl�Ve*�R�
���ʬZ�Rѵ�,jUe+TkJ&���4*)Z*[`��)R�ci�#J�b��E
��B�Z-�֊�A)lB��m-��-f1�PPGZYKF؂
�*���*TYeE���r�Tͣm*��Z��S�e�	�D$�	�����?N�B!�{s-��il˫t���J9��:���'Ž�����Ǻ�S�@��]���������Y
�{�z�l�G��f���Y�</�q�О/8L�Vg�zǝ�22Ua��K���hI�y��J�;��ށW�����zc��F���vc����7�0u�i�t�ZOmO��:2�R���gP����u��^�^��1��-v������sohm��C� �,�7��ծ���?R�iR���dvߌ��U�g����h���ۯx���ρ�]ɺ9���@�����w榾���!&4V�A0�Y�Z}};��z2=^{r竜�z����~G��h��~�n��2�q�T 6F�.�a��9���^�eLF������}�Y9$���|A�5١�{���!T���ȧN��9A0�w�z���56+�mB���wi� �k��Y	���k���s��˱ڦ��ߵsn�1������i��O�ki���cx��Fqxiu�WK���)���xG�T+�Q�~~�Ӯ��s�U�� �c��ҽ�t����0��-=C��Y����:�Z����f���I\���}E[;�,˝Xd.�7ޥ��fop�n+�z�+��랑`7�e!�d;�Xгۚm�5�oR�-C*F�M����ph>Op:��6'�T���{�%r��M\bK`F�^��fɩ,S�ʖ�c'�O���������խ)��	��^9�;�\ҿ;����-.;�J2�}��z�,�ڼe,�PI�͊���y����-�ǳiV�S��s��<ԫr��8�%�ޣ��]�r��;�NC�F{f����w��7�e�	ZO$��2�; �+�!��媼d�"q�9�4���K̕�v;.�#[�y��ݿ��J��C3q۱��c��q�a#�o#PV�s�^�ݧ�K�O���]�}]qM��Q@��VL{�Yu뀃���/��k��*�������AA K#pm,����#N�����kh�'~��1�3�j̰Z�1��+4��˻���SiT�Yn���W�xo�_�/������P|7��M̾}�6�NeAh�|/'�qa�Ƿ��ʵKk;}{޲�tA:]�z,�(la7'X;�Weo{��.��P>���N��Յ���չ�&3�
{v�`S#Գ�������'}���^���R�]��/�Cpkp��K���[q��z�臫��#���O��!zr����ӯ.�;��k�ט������8P��<���oj ���=�t���+EM��2���zTwi/:�W=�y�@vm�>p���p5o��wsR��˜�#�Z�cW�~����s��XcR _r��a�-J��[#�:��x~�k�3��m��|����h�}��.�^�jٗ��R=G�%Yi�v����X�v����Q��v��l-7 �%�LE�V�������yE�C�J�\�v5�-��7cz�F��Ǥ�n�����r��m�1�y��!~'R�o�̸(�/���q"����������r�T�V;ޢV���roqV���e
�vn�7B��M_��X��`�����
&�C:�Y��D�^�2�����R����٧�p]w������:aW�v@thѱK�t�� ���&� 7��l�:Clr�#F�7&o!s3a3�t�H�t�É^�XI�f�S[����k���f��� �_D����d]�����f�6]p������U{�h����W������r.�և��l�d��נ<�k�=;,tj�{�N/�SS��.�'�z�=�����U(nl�G}�jՆ�D���F�V�����<eAy�4���(��Yc�����q	�5�N�È��:V�����\��6S�A{+=���d�vOC���Ox��}1mFv���ɮ��5�і+��[�rz����V�t�c�gڨg:�n���}ǰ@�z+Ӱ�t�e���YǇs�<�-��V��W��[�>\� �<6G�Tტ�f��Jr�7a��t��r����~���|ا4��ŇvQ��]sÖ7hY���^�F���x�wܺ�)��~^���f� pF<y=^g�{d�Z}|2�y���M�nnm'��Ed휺��Ө嵄c��M�tvP�
�1
ᯜ�2l]���G�F�w���o��s�[���Ώ*�h����Rh�#�e����3��V��JX��2I%�z��H����G����^va%���/��pr�1ޝ���hyg��`�]/��q������ �L<���G��r�V4�������ׄuo#�,�[j�U[�O{Y��I��V1� �O����v�e�y8 ��Ѐ����� �fE�9�mԯ���y�.g�l\{q���nt�M68WL��-���Y�z&z׼=��-êA�%<�gn�sEd�>�5��>�x�C Qz쨌�~:캼�����_��y�9�&��Μw���{����,5��}�q�NΖ����=&=ܣ�e�nx꽑���p½��L�&N;�V�XK~���5ő��D|(�{�>���^�zr�[�Q�/rs�ke z��|�Qiܻ�W	u�&���c���9ƽ�q�j��V�Ѣo@J��Ѐ9:��4�r�ƹo�0�8nYv�Ȓ�ᤌM���*�
������ԭ_YL�e�Ek&�-��x>e�O���}ݭ�<�(�?�7~Ig.4# 
t'^� ��c<3���2���U�h3qҘ�P*�+g_����7�!+K�uR]קq���э��e�O��'C��Ng�K\o7LB���6��ܽ^����2�˷�������m���Ǻ�^h��{"��a]uݪtC6���ū��>g��dw��鹅9+!㼶�y��-��dc�iV�+]0{��o,s�9ukmc���=���v8f�=�L>�*���§S匜5�t��^�H�eeY���Z��<�B�oz�{��w��n�(�C�Z�{ҜQ1p�XSل]\����fȬ��\�0������d�����J߼(����<������My!�=���\s.;��!;�Ot�Srz����&�Eu�i�V�����'H��\8�է-+G3��|��n�E�4bt6]h�֗��~�9�RMTϷs;�����:g����/1Y����ؙ���`E�(�:6)�yfD�ۏ.޹o�������D�,�x��c�2�͸�@�5__y�y}�Zq�L'Nia�&����Y�����A�͍ʯr��h�}+%up�Hn~0���f�]�N����1�]�6�'���%�2���f��)\R���/���TZ쩼�U�:v^���N��j �k�Y�B��Lr�u�1�W�,J�h�{!�0��G2��!
�7�d]:'u���©�v뢎����G����WZ;�k��V�R�D-u-���ڱͼ}���{@u��Y�������m�8��]3@�3F��d,u�ɒb���R)��;����>ʖ�Jm'�m#ݪ�m�0O�#]x���5�;�:���B"����k��V���U�?"z�r�l:W)v�D29o`�Zݺ���tvo`�ˉ8�\�򹴄��rw5�x�����l�q-���	n�m֑)�<��emJ�j&\�!�t4Bv�퇧���U�di����9�ܥ�	Y�	�I���d�Avv�-I��0��GHY�	�	^nv��riqG#ЃZ���|ݸ�Ղx����wN����x��ʘ㛕��H��҂�J`"`櫔��yJ�C�K�.��%J��Q��fD�Y�t49T/�0t��
@7���!9����;�
�kw4q��̊��0�K���f�Q�}7��.v������i`�#tp� EN#�Qfwl������7Õ���1}�d�Դr1�n�ҡG��ÍfFy.Ͳ��P�:�Lև�ێ���,����gF�*�7A�yY[9E��\��л.d�z�f�:�pB�P��ʈ��IJVt�.�kܻ��]Z�j֌��r�>=q�=\�X�������eܡ����ƃd���prg��$�L�0�Ͱ�}�Y+��B�K�%���Wecl��=�/
@�E�}��I���@p@����������qA�+U��R�J�6�V����`�E��Z�b/��L�r����[E�b���qB�����)F�Ь�[PF,�J�P���Z�V�m�JŢJ�Z�V�"[��#m�++k[H��U��Ap�eeIX��X)TJ�ֵ*b�E%V�T�
�l�3�*%�
YPYD��X#J��&SK�d
Ȩ�,���e�DaXm���E�kX�8l�J�	*a��V)R,�)+�fV����*�k)l*� �
��-"�2����`���` �A?>)�T{���,H�6�ee�/����%�3U:|X.�2�@
%��_� e�E�<O��o@>�v߀�?y��Z�.Tз}��Jm�(��y�Y����m����&p��=n��k>�3�k�&��8�m_9���3��#�ﯝ��7h?ndҊ����2i�J��u�z�Xn�X���>r�y�z�����Ms�ۊ1�ͪCȹ#c�X��9�)-�}�q���KFn��i�]��޿O{1�UPr��t�U�7~��O��e�a� ��{��m	k��ў2��D/��Zb�P�K�|NmG�A垤���'l<0.��OR��{s����V�nQ��E)å�w�i�I�]:�k����-��lq��>��{���>��K�D��T���A�V��E�@�_N���n�N�%̾�'��IG+�r�DmxT�@���4S�wu��T�T�C�͇�߁�\C�#���M�ٝ*��fz���#��a;��s�{�B�"��^Ï��.��.~�o����T~~˸f;��.p|/ƪ�Ij��`�/�X[����{�����]�n�owR��ӄ�gN;�G�'B�٣�5٤j���M��rxZ�"�I��걞��sc+�t��JT�׆�ShK[	aߕ����ʁZ��ގT��}P�fp��)|uAI&!p����%[�q�]�Sw��wc��|M��7�| ��m�2B
��ި^_Y�0�;��n4߻wI���3�P@�v{�Ϣs7���M��O��tX}��?b,���ɂe�3��Ω����]�VL�L�pLH^����k�z�"�l����<f��u���x^�oCFy�N��l�LD�����E��8C����	\��ݱ{�jju���tV�~�r�V;�i�ɚ��0����mi��db���9Dr�0���	]Mg�.;�ef�4� ��	��\6����c�SU�6�ӷ�s��X��
���L�8p}��M�D9jVݪ�����4�|� ��ݲ��'tSe�eDd������V2��]�� wB�)c[�}˳�3��64�'fE���+O���-~�,l-I��d5J�ӥr��6��Vw���r�����Yն�`̛5AL��z��;��^�j��-���_�ho'z�
��ڴ��]̤�C�I|e�s��*G�p-�#�;�����3`ܔy2���ޟ\V_&�}���'/4��A�;�r�r���L�r��K_�҅���)�}�;����iΑOv8~������ּ�v�Y�ר�e�rM>ݛסL��T�=�%�/&X7�K�鶈�J��*$VМ�|��t��N��[7��D���3+$�NbF9�����0� ��~9�xq�t߼�dHn���vfԼ}�
B�B�\F�tg^�����Y}���*�z?Z"$V�bǩ���׃�q"�<����{�xl�@�+ܫ;&�wO??u�QA�T����kބ7�"y�r�x?p"V����CsC���Y��������b�n�aLVl�V.S����fc�㏜�<�������]�F�cA�'��ЇG���o.��DǓu�[�β�m�%�������6{�5؟`��)��t��<��1��Sĺ�X�-�*��hۭr�q,ùoJ�&|o*hY;���>���`�SܓS��zӭFp��O�G\=��^(�͍���N~�ﾠ/ȓA��~�<��u�{d�K��:��{.>���O�:#1w�N�+^�ఛw�z���Dda�x��n L�uc��K�!����a�[���۔�&Ӗ�;�!�4�+�d�����<���~�=���I�q��¬6�d����޳p���ػ������X�(s��&|�'�"��H+�Ιv���<EJ��I�s���m϶	���uK̞�;.��F{�d�{{	��*R�eҗ���gZ��
V�S���R�-��Ǻs.n���X���en�9%C�K��[J�y�܏L䣙�8���H�8��<�Z��ƌ��\:2D���W�}��#���U��	[�iS���_!����c%��ll&);�tR�z�-���-���ac�9���}:��{+{��Q����v)K[�l��{�w��8u%v6���D�v�l��d�=��P|�۳�Hp�~?Y��$�'<�:�e�5�ܡ�_��gx���j멗0W����+[��a����~� �ި�u�=�n/O�,�t6;�����VR����ì��*���{�,��X��6G�S�a��H�dP�A�%�5iF) o�P��V(:�kUo�|j
��_=���_���̠6њєà�c����������v=D��pܩک=W7���#�P��{��ï�z\��p���&с)���}_
�����?'�'5#���BG^��,�^<w��L���\�	"�>$�z��(��>4]�dx��[�G�� �xGGMj��OX(\K���Đ��]C(,�k�2�z7��پW��U��jUy^��¡��Z\(�˳2 ��~�����Xo��/��Nm8t!�B�[ gN�Oz{����Ml+��Hx��ӿy�G��<z���ە/g�NE�:CQ�^B���,y�kOh4��.���17Zn);���
M��5T�!9Cb��/\&���i��΂A����c�juG��/M:�˪�3uO���W�֛�2��-��c�Y�Rü~y��B4h���
�W�撃��Y��\d�.N��&4���SX;��}��H�����Iޔ�p�C;B��6���I���Re"�c���_����sou.㬧�� ��'"~����}x����j�<a��0ܰѩ
�v{�*u^(C�Y:8AN�ʆ�}"Ղ9��O����}�h���A����S���H鱑�<��^��2�D��og�fsI'����o��m�E�wʃB�p}�J�ٰcR#"z��a���Uqv�x�8�2���nOp�98
!�\z��CJ�xZ���F�;�w�wl�:~z�]���0:I��IVϭ����:;nV�d7���5�.*�~`���byUh��BM�C��f�
�����^P�y�%��b���?�Y/ʹBք�r$���y�>�.���w�պ5凌��sb�؍��q4��q�uY*Ǟ�q�*�e����T�����Ok����6c+�*���ͭw+�;���֬���UL��o��G�����[R��������~"_ʼ+�z�������B��V��F5^F l!�y���]��K�����g���3nW�0��͚�~-����N<G�X`�Jk9n �;*�u؇o��j]t|��v]��x�G'�66��>�-B��?�Ͻ�X��L�G&b-<��>���x�Xe|9�H�=���V�ͱ�Oomt�#�o�}Z�8y!c����%�{�C+��6���adF4;�Wo�S�F��w$X$��Z��y(J�QUY2��5��f�ab��@�e���ʇq�
��R�y~�3N�:L�=Pa�6�k��^#B���!憝���Vg��1ztR�D�3��XՇrNu���:�s��W#���Ci�3�<۝Q�<#S�]p�μ ��ے����VLq1)��_K.1"�Ô�5Syoq��S���KP<��Z,s�뺑(-q����`e�y�s�Q�(�}z��N���'u����d�-����ҧ]ۣ4͈�1Z��b�k�LcS8(|����Gd�y̤��ۮ�Q���0�E���ں�i�p}k.�>!^Q��ݰ��23���֑�*z[V9Z8�9����*��HH��J�d�.7[P�0r�"벁�{�1Yf�9�fq��b3��O �2�
���!W̜f�9�#ӶհX���ӧv��Sn�Ѱ`�-T�]{|u
�Lhǌ��B�1�'��>��In�,�C)͎�P�����θY�@��œ8HI!Kq>�%:�,WwK�RT����MbN��Eß9o оA��,�c]��q��W��2�#���g�[OH �,"�ղ����^=X{)�Eq���]0�$;E˸
{�T!^fZ��S�}وJ*�@��YXJ;G��i�V×o�7�1.���;\�Sf�ח�"F\�,�[C-)�q�t1�W:�?A��כ��]�y#gV�[+!`��`���T�|Ml|�n��<Q6\#�
ʾ�D��o|ր�d���p��u�Bv��Δ���GhRE�87���R�ٷ����Rǖ��`h*��v�Å�e�s)e��33mI}c���A�k�[���f��6�\�ƚ�ٍ廛SN��Յo`����OuT8���J��ކ���W��rc���rYYB;}h����J]�K笕�D��.�=��H`2�:�c��	�v'9lv���r�ߊ�Ί�4�3�ff�٪���1������-i
[S�+���B�V�E�Xa
�ATP�ʀ��+#i+
�Ң��Y*V6�J0�
�,U����`�@*���a�RڰTdX���P
��H*�@Qm*����,�������V(����H�0�P�j "(
9��1�e(
�J��Њ��B��E
��Q�0@˔U��X,"�L$�0��"��T
��PDYXE
&\!)Z�3�9@qa�T�0�����Ra0�j6�����a��N���s�r���z�+��5T+�0hBWI�)��ؐ�$Q�����5�'��Y���E;��^4A���'�DC��^UK�7�&��$3��a���\�G���u�;�OO�gpsk����܏��,֩u��q.b�}a/42��fmNΪ/��t�a��d<��hg�댐������C��"�Ɍ[��QC{�����Eh�T����<8�~��p�J6���RB�]���`�<�F���G�]����P^��uS=�^	Y%��|a8�嚆?<�ĥB=���4�͈�U�ok+<�����x�Z`5k�{�L_�+̮��b�$��i!Z�k^�hkP�ˣoB��et95��hԺ�V�/�?_ā�������cA���L~*(�ʷn^Vj�`u��(�
�F�a�]Y����6�(�iT�l������}JN �ꁬ�5�p�9�d�U8�[��U}�x��$���:�2�у.���0�XKK!r��^��]��m��=Dw.���~#}�g�x�,/��$��Տw�l�#^!
;
��b)8C�!�֬4!b(}^�W��F^�{��j"@�_�>�� �g�Rꝺ��F�b=���Џ���W?#�|C��"��>Bţɏ.4�}�^�ސn�H�b(IY��x�(�E�QL�x(��v���˽݈��_���'�(/�5�M^$��z�������=��Q�/�����>�	?a$��С��eyD��gP"z��m����c��>+��Yђ� c�K���I��� �o��&��MN,V�u���T/�\z׌����f
C��M]_Z�-���q��&��s�e#�=f�h�[��~�޻X>D���<�ΧRj�X���P(K�߲Hs�k��|t{\�ynk����xt����4�xN��BIi,a�ﺥ|�>> iMU*HNP�\F޸I;'p�\۩Ӽ'�пk��8֭JQ����F��������'W��1{�%�"Y��!�y�!��j���[(BAx�J�ު�=�3h�`�H�^��Z��Z}�raq����sݩ���I�(c(a�H��ZP���2c�����X�}��>�5J~�0^|C�^�D)�n +yW�iȂ�<3s��y ��Q���e��I�^3��	M
"���e���rM����Lz�6C������iġ�o����[����^�@J^��<l���jӰ!X�#�����&��:_����X��xH4��Ϸυ�d�^K'�ɘU�|�.mԊ�%�F���3 �}L��(���K���#*O�W�3a��o�ԇ�e���<4m ��@�=�e7�<��p�q�.:^���@�o0�z�"t��}u�ݓi�Q�,.-�<ĉ���r��^���3��R��3]�����pЈ�0��M!�
���ok�ܶEB��=��;��N��]�3�rwy�K�����E�.�k��t�����
�aÞ�6^!�{���[�A���K�e��gt���lQ�z�P�4'��^C��9_1�X�~��{3�@h�(�㤕�Y��0���u�zU���T�U�+9�2MHçO���CZ��}ʭB��0Ʈļvr㙲z�!��$���Ia���	!�����?���!JI�zʑbL����<��;ψҺ�)!dK���`ړ/ǂ٭�[�OW:�N��y�%��Xu��)89���Y4y�i�|$�YLb�?e���ؐԑ��	O_�=V�E�����+�<�����?��o=B]6~�C_X �]���hr����0zz��a0�q�0�mi����Z80�柷sg������|��mW/�����ǰ!44���m�Oo�I��t�T�_7T.��."�0�O�\\�nI�i����њ����ǥ�J����Ib��zψ���QR������-�tY6v᧮�?2|0(�� ���nd0=�%�*�5��ʔ��Ю�zy���~P��^[7:}M��g1gb&�CE��R���{�_����i>��]+�=3�k.]����<)�<<����dyt<�=��ti�P������4����}kP4�
j��G\>�\H�<�T���'S�Nw��S�x�Q�C�{p�3ϋ�iN�Q��ꪤ0�'=�歈�$؈'�CC�$���5���<E{E���E�&U�+�w䬲N�<��KƎ��!��rrr�vw�>�j�C$YiRC��ե,�o-UU�^�/oR�P\����7u���"t��*Hk�Γ���q�l��gyqh{����4���k`B!���~�AN��{�.���1Q�V��V?��1�兑���u��j_e�֊�j��:��%`�Vm���'x�/�i"!�u�(�}y����6"������^
��pp^5.�_�T�E}�����G"��;,dh�1x���EcY�O,����|�%���<���b$C�HfkD`>iD=��L׺�K�d�u=�vK}W9�y���xo���Q����B���^���sеz����^:�*A�����\Z�8ie�8�b��|���S]v�N�e�'���R}�p*�z��\a'���!,k�iF�3[��M��� �#�\UJ���
7�3��'�#M٦i�����\��կ%�__��q�L���Y���ӇmY�|*�U�w�2y��S~�aC@���B4D�cK�b�><�:�Ju���Hժ?i��%�C��ey���/�1�ŭ-N�哬�`�����4����m Jj�RB>p���<�n��}�yq>��rx���W����ei�B)k:�/�o�_MD�Xw���ccVZ�/�cb+��|�v�n���,��+�,��U�_��W��Q[��6��c�!��b�:���xz\~�U(�E�w��}�У[��������|lL��pcd]�X�r�}{
aQ��j֛u(�I�KU��A�qn;$�R�A�Ô~&>W2O������7W�9��kF0�~���#?)�3}��h�Y(Ggs��0 ^3ʷ=g���7Q$�/�AlȣC�!%:OwsW4,D%�l��ȉ�aԡ�U����qn���k,�1xC��D=
_k�;�zֻ�/h]q��g�.�5O�Ư��J�W�0�$�H���}W�鳤�a"{��tk��7�*�~`�7�Y�&O7x�k��� �|+�X�����j��H�)Q������~F�)��ᬘ\^>��]OƄD�_u�G�ޚ���u:@�>��w騞hPK��Z,ϼ��y�K������o�.���I�3��5�OTl�E�=�<ܡ[U��Ssد5�c,�������ݍV].�+6d�~�6�-�BV�ՒhW�u�r�:M��s>�uqݠ�ܸjb}gy\<��0a�m���r��x�T��?tS�m��xm}m���pr�����RQ���|�F\���w�L:3��H�o��a%�嶇z�<"�w�{N<wk6I�O+>Z�x�|O!䆵��>�V��!㓱E��Wg��k���ŒwJ��A,3�$�#�g��Xׯ��H�b�O�8�(F��b�m�������왓�dBH���������l��	�'�"�A�gɼ�ӥ�K�|�&�v3tj
�=F��Wʇ�h���β䁯
4�nf]��U���e����C�z��97c�"|x�-&rS�H*wC9x�/yK�j�K�d��xiJ����D�j$2яK��
�~B��M�xU���Wa[�VB�b6���E�U�8�t{�����mEXs�����=_Ǣ�K��]]�o��;�do���{�d�X���_>���Ƕ����������F0����F&�J-uYu�tz�3�|0x��ds�V��F�i��?S�4|T�RR#��<�T�����.��.����m��+l�vئ(�1����d�~�lL�{'oW@j��i����Q�4k�Mz>"�}�:�C7�"�F�5c+O��UJ
�¿[���Et j-'p�=��S���.� 2z�@:W��A�]����,���gVE�CJ)�L ��9Bֽ1��BL���U�6�;| ��E�+{l�0V�h�J/���[#^�Q�9��]�C�C�����1�:rs�C�"�ݭo;;�ϾA	���>s��"r���������������/�<*�����ou��x�2���{��=j!2�AB�������P1s�=�QNUԋd���θ�2��ov�.��r�z���=G�k�m
ɼ��;������F��8�&Yۓk����۴�!���U�<�3B�ŋA��r�;h4t��q��D��Z�����;]IJ�d��1bb�S[����p�k����%	�mcD�a��Ƞ��Vue
�.�t����W���P\t�� .��ų�o�8zʉn��L��2��ǵ�1W�S� sK�W�0�Sm�@ŇE܌��@٫�<�V�2#��^�_�|�Q5��N.Yb��ǻ�v��K3��++k�n\�0%�u���[M���JP�R��$�[�:���NѺ����t������W9�x��|��E%��W�i
jM�D��&-�rn@�r��7�d
9m��K���Y����:���\a��خ }*wa�4�%:v�1��S��\\R�G;��U�s!��r�<2�U����Ⱥ0���l���4����*E�W\wB�8���/cA�ڳ�̎��O~�&oyđ�Ρ�J	aW2�؍0�h����@���ަ���i���j<���_h�}#�4�8���s�n)o՞�o+�����w�Wz��O����$	4`�,�u<.V[%ڣ�m�2�"�Hr�b���2�Q���^6��Ja�.�T�s�������t�X}l���|*�HV�m+}�#�:�6��e���B���-���S����sFrRX�멒�3#�]ۻ��6��t��i�2�&K�+zD��.M�̙H�C٫�۬p9��Ge���7��*�>�v�y|�����E}@U
�ZM�������ed��a+JإaPX-x�(.-�Q`)�RELPÁ�+"�@R,�B�&RVV
�Be��*���*E6
V,(-aQ"�d��a	m��b"�SU��U@RV�%�E[H��T�V6QX�`T� *$Pb��C�E����YDY�UQD""�����_7ˮ�/݇�:lr�2���y#xw^{�a��OB�R��v/y�i��%�ic�,K�㺅e'c��-�G�Z�]�'�P����=�c��h����ͳ���z�Y��,�wSP�DϪ1�_o"n$pꏈu�a(��Ct-�rY�q�[ly�h
�wRջ`Q·�W4+�K~A?��0����qAƊ�[㦹qq�.%�N\�M������E
��P��{3�v(Q�|��	���bo�W�����z�h�+���ܾU��u3*ؿ +5��C�ׄÛ��{=���dxZ'�ל�!���P�lx�����>Q���,��(}��<h�WHx����,z��-Į��}��-�px�E���#b��J|p���j��GVM��/=�a9x�߉��A��ʾj�.Ǡ�h�����Yw��l�v\���X�K�jk�oN�\��Z�G.쵡M���M��ɴ�D�����\�zA_�����������3��`����Z�|T�n ��z��[7)w�y�(�b��"��wS��Q��6"�'��_eR��zX��Q��<�B���'\�Z��v�h{#Gh����.���.��tw�Z�
����־�H�H�ç�/�k��2C�6�Ф�*Ǚ��g�l=Sˋ(��9��j��W)m۩�b��	y}�P�V���%6C��VFH�(^�}x�Ş��纰�ÃB�^
�A�q�!�l]q�X�zOw����-��j����	W��\��Lu����{�<���^�r�!ڱ奊��_�3���*:��"�{}��%pA��/�]weY�n�y��P�$��V��u,g&^��V�^i1}���	֧�9V��R�g�άvqN��;��Mu��c��������ۿ�ZF��VV����y�$C,�1->T�M�w	���,b�!F'>5��:����5�pZ64?|�.����+�b�?�����9
4���-t��߯��F:}1�ç�#e�@й�__���X���|�()ރ��hx��hY�Z��p�9
>"�,=Fu$���jI������UC$�t������A�I1֯J�}�y �aR	Ἶ��=4�\P��\ǒb���ܬț
�3��M�	B�����la'%P84�#>&�����?z-�ڎL`pUt9�#���[GHq�PX;�����=ٵ��Dӵ|.����10Sg��N֍���!^���b�]��%Y�V���l��&0�eQڻ�ׅVޘ'ݖ�I\��歴�E�Z��`xuG�3Pk�-rz<�ۮ$���Wؗ����[��m:������aF�Ze(B�=�����ޢ6��Vm��s���G�\F����y(���s~т�z@�� 0NWd];���ŋ@�~��U9e�w�n�	ӂ��m�����,|������ѨL��^��p���
�<||I����7�t�ˮ�[w��=9t�ڻ=Q�4fs���,z���⾞c�h��^/��.�c�����2iS:<�:鍈��B��_g�P��{��X~�	"�y\C����Qij,3��Z�w �3�Ӹ��lz�����t|h�bP���Onh��=/���M�1W�]0��� ��xX����=<�r��1M�'�7x36�^u�)���t%�Wc�}yB���Es���D��C����훬F:s�զa�v%*�\7mu���fe�"i���}������5j�
P�L�`M*Ӣ�^�E�î��t�+�����5C{��Zᯈ�I�N�F�R�����p�}m�4��^"�c	�:k'P�3�0�o��X^t�����x"0���.xm|���O�o��_�7����{�F����G��=��5�O��J��"]��<��ƹ���i{{'��~��W�)LZ�Ǟ�mq�fz�~:Q��{���MĎ��(�׃֒=����Z����c$�lj��1����֔C���DB�_I���ӥ�a~H���7�ň��i�<k_�1Nyy������jү(*��m�P�������h/��t��UR�Џ�ɌU�y�1u�c7���2��Z6�V1c��v��p���WWGr��r��<��(��F�Μ0���X4�����y�mqSdi��V��~�/��V'�_�ߗn|L S����=7�FX�X�X� ��	�����/�U'�B�>� ��Y|g*#.�$��*����*G���4C��N^ ��ƈr���[X���A�wU/��:�Z�^�����j39�mx�+�֟���
�r�����(�S;D�/��@aBC�P�z���o�����PA�
�.�v\�sΣ�t.y�^�������-ˌ.S��E� ��+Jj�������}������[^ �֋�h��ݨB/��L�U<z��AC5y��x�Q��v���W��uDj��wuY�걙�4�B;wv��K�u�np�;2������i\��,�Kf��4��
b��qm_Yvw���o�����+�֓���JA�U�#���9	c�!�P�C#$1�]:�t�¼��nm��c��k8�;�u�^�R�|�4w.��(�X��-SSWXo��T<~q���<ap.:�V+�.�3�N�$FFճ��Ձ�*0�W�_�'y�;_��_^fo���R���0�8E��i�W�'��.6C���{�U��%!�0�_p��|4��G	�[����t�'��QÆ�1�A��F�{��qNB�%�x����&�Of�˺#C�A�U�uc�	�/l��{�L4�Wt;���Z�T���C�ŋZM,3�:w���y)E�$zb���5#�C�a�	)��V��z��j^a��V:���40_R۟~�<|�y3=Q��9�t��}Z[�E�by����D������P�w]]�ɆC�	�o^��o�cq(7������W��m9C�ycci@l�ܽ{9����ܺ����R0!��$p��W�SJ�WȞ�dB)p�����v�#NE������Fg�9����پǧָ�8��P�3����l�5c��o{������dѼ^	j�q�-x����6p��kLzx�w:�=:i�!��p���T&��0�#j��ǈ�Wb��pʏcJ����P���U�����h�j���b�WѠ��w�2�9�5��x�$�ϲ4ek$Qg�X���PKw�>�o�î���cP*؅��	:L_]�QKǉ��X�k��mw���=5��ի>�^!�S�4|T�Y�W�sI9�k�wޜ�E��������W�}���g���:l�tHb9|�9{Np�>΂t��l��vμ�H6�S�í!�;q7'������Z�\�~ZX"���G�B�ET��Ub��Ǉe�)sR6�}>f�L���/EY:>\P��� ���Զ�gz����Z�(e+�L$ߐO���-|`�6kOzyЩ[� 䲞�u��ZA:ǝ�$��.2��r��h�l{�u����q�|"�;�L�\p��1E�i!'V0�1*��tw(I��!��s�lP"�+\?]�p��'Jkxܾ/I���y!n6x���/V�4p�9�Fn�>[z�x��'��z�t�(v(j��\��O��(X0�ϯҚw<���q���Zw�B����M�~#�ℬ~3P����<.�{$!趕44��a���y}��"�4���T<|v����ۛ�Vj)�kӷ���7�d|�x�8#��0v�	�%�6�
����!������&���*��Qx��j���O����ĺT�o�o�y3�yiy�����J>!�͎��~�Ԯ��w�e�4������h��
�b��Q�/�Ak�+o;�զ��c��*�(�Pq������:"'���^�:�����E?T���Vn��գX/�"�����҆��3������!w��P� ���y��ώjf3K�P���ܰ���z���px!��+��F���P��J�]�[Ar������C�t�0�^�Ǐ<�#��eW�����r
�t����u�����<�ȼx�����[^��cu��JˋH�P�_{����{�Zt�����ˁ�N{�X��8@���`w��ҳx��+�i=�@a�W�T\�uqLVt�=3��� ��D�#8���������"�������ɷ�̇��2�u�O*5����=�u�v�,�e)��5�z��ڙ��ji��H�ѩ	�˗d�9ݶ��y]&̩�	MÂ���$"�>���Q0˱��A��-]�Q�
�|xѧ����ow�����*G�7�Jwe�+j+�����7bw����s#'@�]0r���Zs�2�<�6�l`>jb�:`쬭��maĲ�E����\AyH�h�[�s��Ѡ�g>��b�l���R��v)�5&�UP2���j����ii|���)m3�Mgڲ$"TCŽ�Pձ��r�{l���Ƅ�{�5g+�gv����lZ�Ӣ��b��wIMdyS��i�u�.�-��ؖ`�0^Q��q��ԣE�Ш�9CxV����{(;Fd]YY'�g.͹W�ˡ�
�^b����)��(��ʦ��ޗ�Ra�%IP�5�Wp���;�3p9����sj�c��[k���.n��{ˑ��l��g�3H�өn���c:�`�i��F
w�C9��&�Z�7A�|���ޫb�q�f.��X�IPU�W5�7y��4�.�7ev����»���{�`Y�İ���e)�2ۚFZ��{��ɜ	�צ�n0�:Su>�������r���D��M���y����S�ӕ��͘�VںȨ��Ŗ{-�o�/�ن���S�2��*�wYu���0��S�1�ꡕ���F�Yp��V�m'�+$����~֘�nYӼ(/$�E��o���n��G�d�o��!��o��56���:N�{�_fMi�/pTFf:;n���⥣�:T��#]]l�
��v�]w�*"+*�E2¢$�
���"�*�E��H�[E�dPFBa�v�� ��"�.p �,EX�,X����ea1�X$
�Qb��P�*�R�ɔ�k$Qr�`�0�I
���E��
,��!Łm
��RE
�,
��L��Y��En�<5�s��o�Ůt܍1;Q��͗�&���/uQh��,���� �9�Z�F�c���ؼC0�Xm�����v�q����U�꧞�OpZ��
/i�3�2�a�!.~�a)���~��A�ݗZY�ykA���Z,yi����bZ����;��q�B�#��y�����t�c��A�$���k�n�_'*�o}��@���E�p�*g�O$F�D"�Tb��֙�u�T�Y����S�GZ#��L�4(ek��ԙ��o{{�!��a��T׵u��M�C��%��<aS<�o&/	u�ٽ�G�G��Da$KG)�//�q~^�	�۱O�y~�`����q��B�*�Zk���N�`���*�'���Q\a��'��x�ύDO5�Z$yo_�vi�b����W�xdEDTڕkj
���Ju�tD��<��q��N��n}K�s�V �Щ�U�+��=Gn+9�W;��oous\[�����<�����ӇL��������.7�v�.9��w^G[�wR���i�Tl��z_����4.u���1���f2�C�0�5��B=BΓ���(a���v[1T�Ӥ/�+6��Y��y"H�0{�fY�TG?���};'	��j!1}�禂���yC�yg͍�ye���=��މ�	��N���Uc�,gz��4���Ys�0��UTM��*�b�#NEđ���E龤�=M�>m���0����Cx�g]lWc�A����{ʀ�J �Тk<|O׋�<�m���Ǝqf�Vw�=;�!�4�>yT&��1DڱQ��Ƨ���´�}`T=�)a6��m���pa�6ғ���|��'ˎ�,C�Di�|��n�U��ܷ(R[Ҳ��KR�����aJ�=� .:��m�����nqi���y�����׳l
� �9^#F��Q��-j��?5��� ��9�K�����q'M���͟�c� �}�����g�pn��+�."x��؅򄗨���QM�<U�5t�%�^�o��c7����Yn�Z��9��q2଩^R�;�2�;-aFN~��ϫ��|E���h[���,���D>U�n����7�^��;���U�j�KL_+#q"�
]����:��/����?m�47���	>#�!�<�ށg1����n�0�E��w^�mU�x�`;=|+��K֧gU�������5�5x(iB��M1��J�"]榲≱��̰sΪ����Z�[J눭A��~͟?:��f���8�a��v	���k3��5/g#�ܵV;����>oJΫ5��z_-a��rJN-ҹLˋ@c�ٓ��vU��2}z�M����J�U �
�H����)�R��yR���r�?#�'wG��o�aZ^-/����~C���Ja�4)��i�%�X(����|�����Fd!�,K��P�2�Vã��g�6F�5�0�cc&ǟ�~��*��sk��R�N�1�>>(�>�w�w�,dh�1qbA�g�ɞ�������;G���x؄��u!�6����Ai>y7��fD�套Hx��E=`�p�.0�����r����)���Vn׶]Ql*�b��^V���Τ��?`�$
��3(������̞m���΀RD��p����Z'b�"E�h�$�fZ^�4l�h�%��OY��[X�t�9���*��\�]��R�[��J_��|���I|�^�]j��z�5����A���?����;�LwP_���j�e~�ų�8��x,LTF>��;m���X��թ������x��>�����z�b= �ު��a�C�U|>�,�B���Ð�W�0��O��ϋ�@�P^cz����'ڸ�Z{�Y���c^��T���PjXUB��@Ӡ���v[�)�{n���Tdd�,/J��r����LdH�(s(a��K��w��^!�G��)3�I����G\���e/����Z<tÈ/��@�]��sw�A�IL��#�!ȡe�9�mbwcʻ%S�V+��:m �����ySB�<į6C�p��M����1�������Y#��4|D��uyQ���W^<9�1ܽ��������&�홰��,�����4k�,���<Wm��+m䕠�S��\�iG��ܶvG���J�{�vaM����Y�y��}�v� ����G�_���ng�{��{�O�A	kY���W����6�:X�H�G��hYb�O�q�+�|������@`����
��Ɗ��]u��Fa}�G�z���e��Z�;�^y�ʹG����D�)f/1K2��P��Y޺���ڙ,i�4'n�
���ޯ+0��p�tk�_W1uƊ:nc�X�z٪�0��}��;ŢOu���b������(�h�C~P�oOj�aj��Uz���Їݬz����}���;�I#�����j%�:�W��!0�����	��İ�`��)���\��;��,(r�L� 0���N����3���Ot�_�7=�Um��ń�Q�S�X�z�-8�����,���TdK�ۻr���5����=ʷ��&w�e;{�&����6$�Mĝ*�WfY��)�������S���r�"B�ƾ�R�{�����-��C��F�cָ��_7Ξ�:y�(9��I?PB��ƅ
�<Q�^���O<$5���������fU�{w�
<��ӆ��3R�����DC/O�/��{����eY��Ǳ}���0����v)Hm�Oy�W�:��ᦗ����<l?#˨F8���H�$"4�h���RbeuM���#��XC�$�"���B#��z��_Ev_����	!?1���C��д=�c�O��x��ץ��/s}���C�+�AG��������G��݌
�����{w�M1�=��P�x�Mg�j�ȮR��7�����ۮ�ן+�yo7E�� o%���yV��ֻ�Y�vdq�/ev��5"c^N{{-��+D5y�C$C r�����{6�G�q�Qx�,��Ƹ�)x��~A�p{���%����R��ylL�:�ǹ(�R콬����Ԉ��i��;��L��	�
�Y2��
P��0��ώ�{k'xt>�y�ƅ���5�`�z*�+�/x�,a�J�y�v� {b���M���~zk��U�pR�8')�[4��s-=���@�m�Һ�-./��u2��V��b��?/lӺ���\�,�谿/�F�D���~"�b^�Z�v��%��i^#�b�yg��a�"�bI9������+%�u[��ha�ּ}������'*��&�4aw}#�oûr{�2�IY�|��B�<o~-�Iި~�VE���v��+ ·���w1*d��AM�y������V��n�&�[�	�B�d�SrdUd��c�9e��)Dԕ�7͡pξ��q��κ${��A�:�4�C�+|µ��q�x�O�Uurxs�(+��0>��wJ�Q���� �p�3�ʞxe��%�q'H�q�CU��/�z�h"����*�rm�xh����BS��E�tj&1�H�+�m�G�< |c���Sҷ7GP��B�$��ܧ־�#��1㝸_��<�����E{����ܳj۱]�c����;j�m�=����S�7��χ��ť�h�	t��;X�]���i���u]nH4����^�ƈE$2s�0Td��ۥ��,m*�{d!��/Q�k��RiYa�B�qDc�M�q�	Du��zA���ӽ���ur����{Ja$E�t	7���d{�������/��=�ah�4�zen\12���=)�(�� �w�����3�_w*��ڶ�9[����ډ�f����R;�3�����
d��d_�Cǈ��f?{=�b�5�Q-�,ц瘍o.7I�D�����E;�F�&���f��45u�34��Z�p`��z��f!����Y#ǻ>��ů�6��ǩ8�L��m�#�����s��C�pCAӉ#�3>�m��ﲅ<�W<RE���_Ui����t�D��}N�^-.��+�Α{�̼�	V�c�@�/���I���!�=�CV�e�vt�����j��4�b�M9��\@C����ϼ�jw��������W�yY�����X�Р��ua������eD�G�O��·�����/��.�N�
߿�p�L��hyĭ���0v�e3���[I8�)v]`�6�UX���M��zХ�W�CD�3�t[;�X�ݦ����E�5��R���.ƐY���p[�hb�H�k�-34Ԉ.�y{��T
5���^-�qa��dh��ܪ�{����#g���0C}��AYf���4�2�n�|ff�+y7#���+��WF(��P�¶FV�^T���r,�eݍ/������>���Ն�&����E�_��^PZIGz�!���F�vY�����.��a�8^ۜ�?f�&垑�r��N*���r]ى��+r�[�rD+{��=̬��jo�����đLXͫ��P>��*�D�i�Q��.5�ͦ�.u���B�U-|�VʴZ1�G�"�q�W `�j:��o"X�>
�5�O_�㓳9��
is�*9��m���x�w0�Pn��d�SR��fS�����c�Ǖ�n��fA?�������t���T�N�1�m�ݫ��G��.�`ܻJ`Fk/����e�]�n&��rIwg4�GS�F�:�9��8�l8a�6��L�ǦA���ǯ��N�e]H����{`��ՉͩΩJz0�8�v936��h����wvŮ��$����ŵ`�X�����.d����_�
��c�H(��-#�Ӕ{]�F�t%a���3�e&��-��!�v�$(��v�`��%<+o�T��@��oNlWë�FS���[A�)˂�ۦ5�ΐ�sw���w<h���ޑG��:�h�[�u�aHL���u���vp���;qu�WT�tcxt+~�" DJ��P�,���
�B#"A@^!Ra$�[!�C"d0�"�A�J�S,�!�X�d*+Zf� a�H�qJ²T�@��R��B�
�X��J������Z��d�m3q�H*��*T�A+�V\Y�\�Ud�Pֳ�-�y�l{�S�x�%du�v�nfӼ��b��}|(�ʯ��:I%%�gߑʗ�ŇJ��F@+��(M�=�W퉙��mn��wHd5�o��҅c��Q5([W�Y���B��cC#�Ec��n�/h{b���<GQ��/u�Vd�=��0��-�ݬlY���#ST�05:��>~�ޢ� R���/������lmc��;�G!��S��ݝ=�Cؼ�4����^"��z�־�����ڽ~ݞE�r0HX\�U �8�.6|l�z�(�������e���a�Y�ǎ�bj~�"�=|��=�w�.�m�\lrBk㑒4�6���wHKq{Z~W~t�����F|��y{�_�؄��qiiؑ���ͳ����߄��<�ovv;��p��`N�U�ӭ��\_ݴ*,j��6�2J��[I�%�Y��˅��L��kySw�l�����@
JN�s2H��KV[�,�Jj�������"��,��l�}��I��C䃪cş>��C�B�q�|��=T%Tɒ<>#o��=��W����룃oi���Q�s�`ުo,x�z�e����Q!�����\�p/6p�I�Ę,&��+W+�������Д6���A�ʽ���>?OM'��/�u���_� m�,_NL^B�ؘ��/��ڬ�LVӮ�@�}�Ej�5/�=i3�~�ox=Jφ�Z�]0����ƚ�����F�NT����}���x��D���r1�:w��M/V�g�x��wy��E�q�U|��4��H����<���=�f��'�0"�\%`�;b�����3.�AJ�$��G��0��#��<v��56�zN�';��N�k�:Dfb��V�-wI�ޑ�$s�t��ư?���¦�I�Pg´/e�{���-���^�!YI�~�,��D&�J�iG�f�������A�V]�3��|���gH��ry�)=76t�;�$p��/��4�Fл^><p$!$C�z�z���~s=��'��Q!���>c�0�t��<UF�~aZ��mӽ�{�F|�׍(`}j�~p�~⼠<A=�)�ړ�uufO
>�a��&�Cp�l�KMw?�<�*W��k�o�b����T:z�����-Q���L|�#��^�L�VOfq���޶<_��$���r�,�Q)���Yy�@�
��Q�t��ƾŦB�r���Ծ{T�q�TD5�L��Y-�4O���U�a����xuۧ���1ui���H;L��lik�Gd.��mS#��T'�62nW�Ħ��&x�7꿪��U�/�ҫP�Oc����,Ê�u�#sd��>6ms�0�~$�s�#�2kW��M�O]�˛��:t�㚾؆E�ЇZ/ð�TeY��9�1=��c%��تF:���a�&YCܢ0���ߟ��u�2Z����
�]����1Ԑđy��ܘ{%U��y��!��HY����.,��_(0f�g�zN�G�Q$�->��:`���bϚ�O-hki<DG���3H���ŒƮ>m��2#j�#��]vl�z�m��J
�1`�5T��]���l�oX����1�Dڠ��*��d��#���VE!�ey1En㥐���N�ڨ�m9�m�7J�^���QJ�:����y�^C>yh��a�cw�k6�\�Qbh��S��;��/�*rri���2��W<���@���DBN�j/��!�շ��I=����ڃ�;U4(���x�D�<S���u�s-'T�����0uX��C��G��^����3j�'���a���T���_i��&� F3���٥�+O���=Ws�XDm��~n!Ƨ�~F lW��&_8Cj��u��:�dNA�hw����Ձ�m]Ѻ�W,Ǝ��:r�����s����և�a��J�/��}�WU�=��}�y���e�p�U�ؼ����IHG���lff� ���P�l�C�w��i�r�(4���?5�I'S�� ����@ߠv~GGn��
�~�YmLI%�+�\�>��M`{�%�z�h���C0X��[a(��`�V7��rך���J�R�w��P�#X��$�LEѸ�D�{S���B�U�B��, �b?%ƭx��L�ɴ��Wl��Y���hF0��#5 kˎ�bj��a{��~�׻�K���1}c�{P��_��t�$鞦�m�gl��Hf#��>^�1�
���qa-/cG�6	ޕO7{�,��+��r��I8�VƟ"�ڌ[�w-���}W��o����������ԙ�;*�U���Y���l
�#����v���X�G��������vzgnv������4���˯���D���CK�E�>���!�]e�i�u��۠fKT�]Z>N�O7�|OL�m]b5p�<�6��W�ǩ}�:��I0l�(<X�w�Ʒ���ZZ�{d����zU�k"��a޻�a�I[�h̭F&���ilճ��c�/�b7��a�k8fćA�e7-��,��l���(y�+.b�|)aϰ�ğ�[��t���rVaD�i�L&�'چ��� �
���w�7�(/zQ���o�*\Ġ�:k��Myx���oW{�]��.;�ǈ�FyT��҄�{}L�ޏ�p�yQ̺p�P]�:����Ξs�G�#E�F-�Q��gM��rJ�.�]}��&JϢ�
��T��z�T϶X�ء�����M���;�}s�m�~�X֡���{�%�6��.i��!�yc�ٯz�=��#@�U~2�
��
F��ח�><߀���rǬ+����ɫ>���cM��a��4�W��.J2��%�R5�R�7dI\�mc���S�{qk�R0y�ɢ���*�3�p�23��x�!����&
¹U��C�T���%��(6�S��9��~kCŋH^gI��[�	���/.�T�oچ�m!7�~lg������_9����S��~c:
�}��s/G��7����p�9~T{;�N�A�Jj��['�+����mQ���-/ާ����Mkov):�}^&KC�F
���o-I��`4�;�1��坝����.�8��F�ﱮk�Սk�0�4�(_�!WF%�]�b���,�A��;KT��	��gT95���	9+�{Y�D��gr��]ڣ�ւF���b,���Yw��ۊ�"��]JM�ؖ��0$�M�|ۢ�wսyܥ�&��=CZ��Fb���������V�&�V�A�#J�nV_n���@6'��=E��ܸ꩟�6�7��|/�Z�xv���G����[��>賬d#"�V���=�ɝcC��C���2Xk��-�z�ߣ�#=�MI��B��^��7�����ᅊ�.xk�ݧq�������M/����Ȓ`�a`��N����C��ԳP�5��-��.���ukG<�
�T{ ��ZxN5Z�w�1x� Z�Wo��it ٘�ߒ��a���*V�ϙ���U�_NI�r��8<�[%�iJ���Ε�ѹ����K�v��R]�|��h>�R���+<W;�`c�!NzF��ڍ1n�P����6�Y9�r+:�n�o���t|��D�mgi@�v��5��,:�Ԯ��jgm��RƵ��;QcS��;g8���2iY��[jbRe	D3HC�XS:�}��a���{�������i�ҝ��\���)���a�K�|��|BZ
�u͋9Ul���}EC/ْZ�#F#q�[ٌb��J+�uX�,]��f�]�|���Z�/�`�丅���{� )8�a*��;�E���jy��Lu�y��^��(����9'uX��]L����r�/���]��,8jog3e�Q��c��!g�Y�d5�2ӷˑ���]݇�۰QZ�Д�kJy�@s��� ��3oS��Q�t��pk4���	Εe�u�B���z��ݲ�X)�o]��.�BYv�z\� ���Z�v���3:n^�toX-�!u܏ˤv�b�x�Au��&9z�Tgs�/D�w��}��cC(�	)kd�Y2R�ƙ��W+M�W-�v%]r��)�Z�R��W�>[2���/Y$T���Oٵv�/��鰊��۫���Wn�E����w����hE�7��:*�g.�8z&i�ڥ,�A,�����G$e*w�0����͜�׼)Pv2E����bX���t:�;��uB��{�N����:�v�%�	�i��$+�*`��S^���1����Ս�rp���3���Y�c6�G̍X��/\HW_�;�I�%�U�5vl���G�v���x]���s0lk)^l=�s){��{i{.�"���y=�`� ���x����۾qL�_e�S�R���8�g���bG��\��ٸ� 1]#Vc���o�T�ʸ����C��Y�����Մ�V�wۜ�5����j8��FZ�:7I.Ma��y�螱���K!�y*>�	�~�r��A�g��bp�u�(���� (Y�s16�;k�6��uN�B5������bM���}�&�%i.(�Z�Y���w�vK��)¾�����V��iݎ��1���to�'��7
�ʭ@�*Ad�J������[TqB���ڱ`�j���F�U*AUVAeB�J��+R���H�J9lf��TlX0�0����%E�b��`��V�Vņ��-�����TP-*VZ�0�*�
a�eC)�b�F�$�?}�u�7|��w��̸�dt�n�1�t��9B����j�7#~e����a'c���y�E���EԪ�	0�y/J����E�V�$�ʭ�8ʪ������T�˳W����mI��d͗�����BR�u�s�"����m�k�Wvj^����Ij��=���󈱋̛��&ths�^G�	3�u`�V}~"s'K�;�;=�wɶ)�ٟm&�
@�Ww�\s*��y����3�����F���M��ާ��Όz�;plӖ����^i���׺M�k������Q;=9�䳔g:y/PFҡ�j��:��j�e8T����N|��=�;���Gq�Uw�&U��Ŕ��YaCK"��v@Ի�����Ze�r�?��v}�G�`sIIU���yK�W����Ԥ���9}�p�Lq�z^Ȭ!������}Q�{�����֑4L�{�q�UA��_���FHX`;�kvh�^�}<�W룦"���j}����U�h>�O˅�c�Ѹ�]���#�#�[X�bń*�sh�'vH�������.泛'�P����}���\���-��y]��>�������9a���E��n&G�`�<�j�����ìÏ��3+�s���Z�{fzP�%��_����S�#ލ/`�(3�v�כ��h�W����x,����H�<S�^�w)��|Re\��N�u�L��Ӗ�Nr
m*�Kiɻ��;�'��/sP�~,��QU����*�2�.������^���+���ҕ�y�H�[ү݌R1����9���Ƿ*wf�Ok]�8؅d�3�j{�i���w$���s���3OmҼ��Z�s�M\Q,ѻ�_ξ��Ƈ�O�k&�^Ҿ��q���a>m�����z_���)2�%��e�X߆�e:�1g��5�<��lh�)���4��J���tdZ7w�z'�y�3�Dpun��g������y�K�pw�y����6Կ�V��jӡy!q�Mv�;XR2��o!n�p�sRX0ɯ���	<���q�,�_Z�+e�&ڶ֔�4�
2�8���nܼh�a=�D4%�[��m�VK}~75��'������<с5�T�d�]��ג�}:uu�������>�3�]^w�(/W{ڵ�'M6�����Xg�퍪;k��=�<�j*���1Pqf����\sS�xF���~�����#���F
��>���Ξ�Z�u��ܚ��)�"͹aK��<�/x�ۏ���9Ƹ_ӏ����f,��Ǖ��Cv<��\h`���UxЗ�]gx�P����V�й�Geܙ�������M��b�5�w�J)�%��>rV��1=Ǖu����Z�x�ܚԾ�d��qrQ�'W��X��o}QX�e=@b/OUҶu�мDM�=�~�x����=�T�Z��xh��M�;�'	Z*o�*_
��d�L�圽^����2�Ise�L
���O�Ֆ�Ao��K�UP�m����y�Af��Zwt�d˼>�癅H/i�j��װ�ż�n�#���>�4�y�r�����e��v��m��؆���y}3��;��way]���3�'K�\]��iAj���q�w����H�7��!Ž}뷝M�B��(M=ɹ�^�p�۱N�g��U�k��٦��p2�[�:��X6r��p���I�8�i��RC�I�YF��
j��Ϭ8dµ4Ə��쾴�w�M�4�Q���uo�5K��ϖ�l��V9[Ow���5aA8ԡ��Bk+K���+�� ��>�IY���!�Κ<�J��FVu5)B�wT�J$����Έs��E�o�������v��FaD�u#D�,���8�����=�I�o�Ǉ���5����4u⥶j_lO��!Jƈ���e��Y�f]m����)��`����_�6�B���9������J�^�ךۻ��Hĝ�q��`��
��z�8�uֲ��O%u�'���/��ޑ�/�tԱr�D��a��b\dٟa����/JoŜ<SBk�.��u��΁�fd}�oO�Iܞ����}�/t�F�cn���i�B�7�k���B1�ej����OӖ9��4`���u���>lxV��ݑ��uk��e��r묦\�nu��r|X��m�Tx}5gq9�t�ԻTT�T�C�(�YO�4f���Ӷ����;��7�8�ܫfP�h��7+qf�oҷ�g�^Ƞ�9~��^��izR�����ګ-�)����Ej�U�~�|���u��n�e��H ?��I�>��xTl�߫j�,�rf�ө���|އ����kF�j�`ڷz~cC����u�RM�mF�r�;a��+�G�,
��]3DZ>��X�j42q��JC��6�=��GI�>h��ʽٌ��j��C�bd��J��vuӅ���^'A��};/-l\�4F�`����
$h�,Rv"������7�g�c���_{����=Y/O��i�L�����cLZk�;�-˫ɠQ���B�
�H�Μz;S���f�EnziA6Wl�j���$F[Ƕ�M��z\���L�)p��}�>xM�'Y�|�<�/�����9%�.�}�W�����c7:�<�%[���~Eاs����������f��MG�r�b鲏]L�}�hD��zN7s�Dfȣ�g`��F+�y�Na��jNf���O[���aP>�H�>V�O[Z�����Ab��v�͝��k��?"�6�]�+�/���\��Y�ޖ(���_S'n��3��}[�c����Ԧ�wy���v�d���
E�]}xl�8��
����Lp���?Q\W��9�����w7[pD�B�4�3^��\72��F����bP띞������\�^oeU��7/�{aճ�*�=}7Sҩ�a�4���o�/ٰV�kѬ��gi���(��]�K��cU�+�nA�c�G�Hb` L.wr�!a��Hji�GQ�@%W�J�'K\��
)I���i���܌�)3'�M#�-�٪���'� 򺱒��]Z�PÇ8�X�ꪹ���w��ya5�w�(I�d�Ԍ�K�}�]OW����,�Q�=2�Ў=V��}���
;Տ{�'o]�Z�9b�٧��_rjRƅ��<~�N�'�Č�@�Z�夻���5+�93�ͷ�w���hi��o>��8zV%!S�O�q�<�J�y���SD.�ס�СE8y���b�D�p��߾G�c}�����,�ٜ,r�i`��w����b"��jEdU�K����JgoK͚�j����ǙukE�F��iȐ{��G�q
/V����Yf��Vwsm3ȫ���0:^q���W���(Ň-.�h^���ß=�nF�!VhvS�h�y�;&͂��i��^�e;�[L�|�Նv��	�▯b�]I�6*�n�V����U|��'��n��ъ%��fe�ku���»��ެ�=FIܔ��\���V-7��7i^.�oD��u��gD9`�4�m��W4��Qq1�mX��Ԯ���-�@R�8f�@K:^���f�0�/�.���˺���)ew�^䇑�{���:�rb�-��^���T�l�F�1�Ļ�u읦koF!��r/�\��}u����m�ŦŬjg���f�s0���Wf���P�쓶^hB��v�[w�lM�Q��[�LSpL[op+.#��[V�i��K� _t�x ݈�6�`�݁��f�F	سbk:��5�V�1a�������Z�FR3��vVNStw[W������6�nI`�����v֥-�0V�2ޣ�w,��t�&�H^U�7"tü���*p����g�W:��RZ=�Z	�vЕ��f`�:�^Q9Zͪ�)`��I&S��LA朏���n�T���~L,�2�q�`�c��IW�\��iXr곬���e���U3�D�<�C�A��y}e�S�ܣ81���/d̏tMne��)&�f��>���"�_2�W�}֡�2�r�\T��R�՛�=x&N$K7cB�x���zrԦT��/\��'k����Y��`h6�X��������Wo�!��$�'ꞈ�LZ)
���*�M�r�L�UU�Eci*(�U+b.)H��Z��G-�*�jE��D*�rҴF.�(�-�1lÉZ�,Æa����Z�Q���
�ª����R�����(��Tb��qp\��DX��Z��X�{��Z'�>�����u�uX�{K�R��	��>���m����nҎ@g�U�K��t��I=⊶�w��B��*�"���v�|=y9�s��}��I����v+�<�&��z��69��p����rP����]����loc�hƉ�!�9���y��k��2�ٛ�8wgi0Vl���r��_y����"��g01^��@�>=�~:��\4o�����4��<��������e��&���s^�R�+ҳr��k�����[�T�a���EDTC�8��dy��U�yīZk��x6�0޵�`�mM�����ZO%���Dc�������vu��fYT�"Hf�:�0��9����"r�X��I�d ���4M&Hz����M��
���٧���^$�&0��S{6.�T�]ʧ/77z��߼i�o��^��v��J<�rA�3�|�#�oK*�? �vc�3��z���|*�n�L�����{L��Xm����9�g��� ���&�,�.Fc�P0���0]��/��C�`�Sȕ�e��<*^M�7�w��E���N|�@�hXT�#"��D^ݍgɯ^�𾅭��&x��Ջ�;��o��M-gOv����gs[:F�M�F��.���ڇ��R���WNU�&qW��']�&�N���z�Q�|/]���BL�`��A;��/�9�*[�I������͇*)9l2�پ� z<�s�Ph�Ky���w6�/E�kdv�u����R��|F���a����y�)!,mM@����CgFru(]�%u��>�er�Q�(��}��c���C�\^�:Q��f5|���_��ь�B>��CN���7éYVN0U����_c�R���״sb�������﹞�p:�ߟa���f��5)�)�T�#m��<Q�q�
;��dO<�i��Yb�S�	�b�{��0�U����!)��`���b����f�[�-uœ'��$r���a7D�*٢�M�eHG"wd��Ũ�,���}�G�B���w��ƫ��6GS�ts�1}���AxUa�s�����#:�t̨��!y�r��-�v��h3��Xw���Y�
�����?W|��^Ӻ'9s��^�JG�97R�	�f�y��ay]^Ś�L���l��U���4�{�@hV�E�S3o�a�*��k���x�t$�����ڵ_w���X���Q�gq�1�dA����S��lPi�5����d1�����ﭫ/�? ��zh�e�>�1X2������٤���>��\��Ċ����y�<K(Y���m��U&��j�u��_2S):�WZ�p��������mG�Nk:��pv�1�ڙ��2����NZK���.q�׼T��Nt�߮��y�ݷ��c�=��'GL�����}P�J\�Y�f{V���3SLrb$7��2Ӷg&�zAU����1��u� M>���l����ǌ�e{;3|��!wl�UOq�?�T0�X�1,=���2f��'��~6��Z��XQ�|����k" �b��k�ڱ��򒋗�|^��?������˚���-vLެ��ilh%;2���+s�kL�>+=f�8/����c�1�ߕ^��u�}�H�v�J)Cͺ��y��5�z��>Sx��-]e�\e�[U�2rG�p�sH(��J�q��U�^�Qj�7:�;3TPM�}z�\Ν�~^ݮ�첁�����,N�M����9��'�9������%$�(�1g�e����P�=�&�f�QZKO_�d ӫާ�"3tu{4ۯ�N���lR8+z�z���ܱ��g}[C�4T�i�Ƴ�J/Wk~��^)L���m�cѭ����]�k��ƁS�㇃|}h����n�},9��{ѻ;��}oع8��+&�YVО���!j1!�NI��u��蜏p�y�%нǪ�$�߅r��P��Ú&d�v+�.��eV�X�X�-��*=<T�?\d�;fn� �6RR�\�vhō��ݍ����8�n+r݀�X�<�K�Ng?P�,�$���M46���(�^�^�oϧ��[�M��g��KX��)�^���{�&�u]A;ɧ\�M�Z�&�һ��p^���:}el���g{f�����!otv�̛bz��2!4X�Oo-�xgK��o'BY5�a���d����j�n_o��Q�~��oF7p,\���#�7�ٰ^���ϓw��P��@����������I��������|Lv��v�����ȓͷ�ߺ �LS�7+g탅sC�om��\�Y�z�\���Cw݌��l7mV���S=�	��T)�
ڧ�-w�N�o6f>͕�t�+=��v��g\M�-*��n��sy��x�Ca�*/�l���QI�}�FL9C�Q�U,g�7i�L��v�\\J�cګ�N��	�8���x�
+�ƴOg����[�=������*� �$�^��H����k��0�zTcǯ�`r�6? �����f�ٛ�\���cc7�!T�8�.� N�t��89���f�O^�[��NA��f:R�J�����Y����U�s�mL�h�ɰ�mG�=�E��c�Z��/9ea�\Q=.Dd�tu	�$���:����ז�د,ڗ�%c�T�%�6fSTZ�d�F�)Z�/d���y�����!i��5Vw�	��7�Ur�U?4%֓���W�=NfץBǃ�٩ۜ{l���Ц��z���{��k�Lcg������{�+���l+���.a����;"��K�_t�k���6e{�xi�Le^t����5�z��uv��_�p��J?E�r���#l9x^�R2�PUΩC���h�=��צ��2��>�d٢�H��q�e��<�u�������U�C"A�{to�f�C/������0�,�k��58`6��Υ�`����c�
��|���8/�_V*k��m���tǧo�:�Zm�pv$3A�\�l�������^ݔ
�y(��X9��j��v����׼�G�%x�)�*!�b�l��7�mr��zP�jۚ�~�(��y���o'�����f��6&��R�� :�^�N�"���F{F���k�al��63�M|�n�Z�[r�ru�a�Y��5ɫ���u{+lyM��<�*;�zȎ<^��ά3kT:Q��b�p@�������f�X���]�f�,��]��著<�~`η��?i��$���S�j
(*����$$$ŧ��$�����HRl��3a��gp���0��0���������d�vg�q6��$��&,���T$��,�HH!���B1ׇ�;G���v���
C��X|#3ܯƄ:'D�_l?�}�I		 ��E��0������^�]z�C�L0C���1;����!��0�K��?�מ%��b_L�);��o�y�%�����<�ɐ�����9����c��d�� I��$��� xI$��܇�H,,�>�}_�9�H|
P�I����r۩O��`5���?A���Ρ���4�l������\C��dDH{Ԇ���	���ҙL���?@p'LA܇���$/�s�[���Hï��?>�~a�����!�{�w.���褐����賑��;L?�>�$���d���1 7*��%�(t�d.��my2C�?/|�����?\���*�O�v��'���|ξ!>���:�����7'A��$���'^��?�P��G������������Ο���	! ~�3�}!�����BO�������
�|���0N�B��/��������ԟ9:��p�����>!�����A�~�����?HHH��:��w�D~���é4jCA�� P9���jB��&~0@&!�d�����O�B	�z?�	�4��L���%�I5��4tJ>'P̓��$��vфA`�N�����h�� I �d�tO d��>��N�g��̧0��(�>HNw�bI�r��&-!��td����!�'`B@90�������C���!! A�ϼ�Pd���>P�2c��$��||ρ�' �I���'�C ��!���3H��}����}���9�������>�����������I!! Y�ϟ_A�~d��B����?�!�?��d��|L�؇�a�C�����I��O�ć���rC���a��A����"��������������>v�������~_��!�6p3��~�|{$���c�~�O������L}_Q����0П��Q>A�|~p�#Շ�><�ߧGD3 P��u$>�I�0��$$�a�b~d0���m �[�����9����r����������d>�>߶��u�{�$�Hu�?^ ~�c���,DC�"�d����!=��'���H�
�7n�