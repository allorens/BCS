BZh91AY&SY����߀@qc���"� ����bE�          ��j��-�R
B�-��AI���h�V�%AVM�ѵ��
P�֨�IE*�D�ZbHH"�E&�$�� �^��1[U�h�IKV��kc*6F�F�͵!Md�j�T6�cl
�6�Im�R�Z0kkZ�j6��6Ec�f�r	�f�+e�����f�ֶ�F����Z�Z�WcekX֛6��cf�[B�ЩhV�mSh��YX*��h�(�BE�MD��MB���� ���F�0  �ƀj�t��:���Z���eUD� 	�GC���Z��5v[�K�ځ������N��Zf�u�[Z��iiS4�j� �RM�})E �w�G�R�R�˫��iK�� [սz���m(*�w��AJ�W�ڕЭ����A�Z/v����
l�=��z�uw���T�����[ie����+>}$�� à��ƨ&�7�;� �/8y�Q��}�}�j��w=��|����{Uy����F<�x5�i�l����
�^W��z zq�w�M <wmEmmfhڦj�2�dM��( ��!� Q��}��Рm}q�y@�4����҄� ��z��kA�h��y���@�]=�{�Uջ�ʀ)ǯ7<��ݛ%)�a�f�h�-�&�>|�R�9'�ր�����z�^g�!��r���7������v�3�k�AR�9�4꤯]�}��U�'�U��A�Su�UK�9�Ɣ�%+[,Z&ko>����Р6���j���7Uvpt�(st��J �[ui@5�[��bR���� )n�]@ qۋZ�PS����S��í��ٶZ�Ra�V�([W������4v� ����F�T�r�x製qnt �[� ��: �=�v �۫m��$X�x��Ym��jQaf��@�歹 o>�Wۦ����ہ�C�t=���� p ��e� �mP�����ӷ��: ��h�i2f�k5*+A�>�T� 0�/|�N�:n%���jd��^(t��e  �=� �� 롴�۽� ��� P'N��k�,t�Ŧ�Dj���J� �w��v��  N/N@=�`���� �wp �Om���� 9� ����� P	R�UC
*� j`�R��  h  SƌR��G�i�1CL��4�~FBR� �  O5JT�db0&����)MUL�0��2`b�j3JI&S�j2h��L�M�4��_��������E^������r	�Zxh���ay�9p�y�ʽ�҂ ��b"�APS� *�����#B��A?��C���~�*�� ���$�O�
 
�``EO� 
/����_���`��3��#ضĶ-�-�la��)�[�6Ķ-�m�0-�lL[`�ؖĶ��-�l`[�6���#-�l`��6�������SLbi�lKb[ؖĶ%6�[LKb[�Ķ%�-�cl
`��6��%�-�l4�ؔĶ�m�lK`�ؖ�bF�-�lKb[ؖĶ6�1-�lKb[ؖ���l`��6���-�l[b[��Ķ�-�lKb[ؖĶi�lJb[ؖ�����-��1�-�Lm�lK`[ؖ��e�m�l`�ؖ���-�n�`SؖĶ%�-�lKb[-����%�-�lKb[ؖ�Ķ�m�lb[����lKb[�Ŷ%�t�@S �lRؖ�����6Ķ�-�lb[�Ķ[Ķ%�-�l`[���e�-�lb[����-�l4�ؔ��%�-��-�lK`[�e�-�l`[�Ķ�m�2��L`[����-�la[��ؖ�����-�lm�c��������-�l``��
�b#lU-��T� 6�1V؀� `�lm��A�6�R�i��b�lAm����(6�R� �4�B�
SKb�l m����(6�F� �`l)�[b����
�`�lA-��P�
6��R�"[ [b�l@m������(�b�l-�b�lU-����(6��*[[`�l m��� ��4�ؠ�Kbl m����*��H�b�lE-���� ��؀�[`��B1A�6�F� �`�lE-��B�+�[K`�l-�%�T� 6�Rآ[K`�lU4��*�؀�K`#lm�-��(6�F؈�i�6�Vب送l b [[blP#-�-��6���`�lm��`[`�lm��H�V؈�b+lcb#lm���E� ��F��`l )�� � ���`�lTm���E�(�`�lAt���b�l@m�-��(6� �
:`�lEm���P-�lAc [`�lTm�-�A�(��"b�li�	l`�lm�-�A�
6�F���m���E�*6�ت�m�l�$`��6�-�lش�Kl]0-�lb[ؖ�albi�lK`[ؖ��%�-��1-�lb[`������i��)�lKclKclK`[b[`[4�����-��-���%�-�lf�[�[�6Ķ%�-��-�lcm%��%���-�lK`��clJ`��6���m�l2���%�-�l`[���%�-�l`�������ؖ���Ķ6Ŷ%�-�����m�l`[ؔ�KlM0m�l`[�6Ħ[�:`��6Ķ%�m���6��ؖ��%�m�lt�[�6��%���m��1-�c���%���-�lb[)��-��%�-�lK`[���[0-�lb��6���������-�l�����߹���@�_������n�H�6�WuJ���۔��r��D`fa���.J�UJ�U�G76�VNk�`�UsZ��S�47X�����Ec̒��[Wt�d݋^Z:�b�ں/-�b9H�̙�>�g4�i�M;ɯ!����u�f�ݴv4ʺ�j?�h�M��&�0��B�I�pл۰6� p�u�b�QwJ�8��'a�dk�H�[K^���k��Xb�Ĺ�e��]��n*�$�&D(ێ�M�u��f2�:!M����٤��/9�s�X��Ӊ�c//^Zou����1ʡ�K;V�,�T�R*�؎aw�f�Q�,Q��h���0S�ҋ��uP������.6�nVn�Q�`z%�8tR�F5J\�2'���/Ky5�6����-S�j��2���	����x��!��+�)3�E���N��v`"ALo�FV�+T���RMu쾭d���\�U\����D�h���U�A��,I�N�B�r1x,6]Db%AF��=r ��X�з�ءx"�/�5�L���^&+Vi�T���{�5�fe�M���͙I�Z�:oA���$\#����J�-{S+3I�b-��,�d�W5ۦ-��Vaz���*˽�Ж�=h��g�ugZ��,�GE��52�� �aRT<e��K.��S���Y2�nZ��q��vÙ��\�y�te6^	7�aÒk�4���ޝ�)=heŬ6����P%R�̡���tcw�IP��	���n������N��KS ��v��L/3oD�k���dպ�	�fQ��Gr��H�`�O'WT�J���I�d�!�zL�A���i��٤v�8�~NV�tȬBj`�z4��R�]!2���Ķ�D�m\ͤ!j�weB�#�L�$lj�U�Y�i5Gk.��cY8.������հ�e��^f���&�zh9����Q6f�֡w�k��+��u�rͶ�0aO�^��h8mS�Y�7�6��{S6����O"�F�������@����f^j9G*��i��X֣Gl4Y��LWZ�u�M�V�����R`�6a׷B���P_��%4ft,H�%�j��в�bx&Kb�Uo�L���w�����N=í�k��L�����aœF�V���>�ֈ�R�cY��Uǃ7qǴ�*Le*�c��U1�7���;If�Uo��6����J�M�{w(:�(P�]ef�xZ�t]*�G��R�O|e�B���o2�^TՋ�R:%oPf��W.*�9(��%�sY��GM�tUn�RE�Z:f�\V42Ӭ�^����z����һx4.�4��o��x���y��x2p�Kt��ER�J�j������ͩ��5`JQMn7O{NmÇr��n޴
�n?4޲L�X� �^b�U��Y�k%+���dj�e��:�Tt�<'G5��e�x����A�ʿ���Ƽ�˱���I�J �1��x}H�k6:3r�4�fǕ(����j�&:�~��^Ñ��0�U�%���
�����aMV��W'n2l7�-r�"�D���k�c��vTc.�S"�UK"��yO!�c�̑ح���jj�G*���G�ӭ�հ0�d��h��K���i��og��a�IS�	�ה�)YaPدr�א�uJmn�͠�I%�[�!�z�vN�ӤA�+yV]�ղ��*�,V�-�x�@꓊���B)��n����n�c	QM-��0�����D&hJ��YN���*Cz͞�x��I��p�òU),4'jY�B5%��74fJ���팉��/[�c������ݶA�GBe|��'�8�)5�ʙ6Mv��AM���4�s"0�9-Myl��0�A�J��V�thEjI��dïrګuy�i��	်�V���[ ��ҹN�ՍٙP����1�[����׺L�Öj�Ma�PF�,8�j��9���-L]�&]+�1���b4ݶ����T���M=�:�:�+Y�Դ�������*�5&�6��Z��B�3�#乛�hu��vμT��	f��<�[��N�dVة��oo5P{� e�̓bOR�%����O�t�e7�q-�ù�E!�n��Ӑ�V��˲1��Miq[��C�ƪX��-��-����j��n3[�t�E����U6�x�7v��Xn���f�� F�
�kIR3R�U݈���1�*lb:Z���Jr��m�!�U�MR��i�p#�54$�̹�[Y�V5�F���m��NśY����E�Ŵ�4��m�MV����M�_<�m^������T��5��ve�)�Z:����G��t�[�S�Gx���÷��1*��#X�-���J\����+F�y�;հ��&��VwՉ�M7[�*�^��gr��u+�Fm̱ǹ�O^���*V8-�%��Gi�f�ڀ�w�0Ō��CD���S5kUU�%7��v�mQ��[̄��Gd��)ި�����Fnа�Fh��S.�[�/H������aop�X�Aз6ٔd��/p�]7b{W�K�%���w���L��O2"����d�~��U�T�!J�1#�uuE�����.�i���G��geav�ʘ�d�(�j��K�UѸ�1ofV�Q��ݵmZ1�S��L��bNd��q��۩M�ғ�XB`����Y)H�:��iU4.�ˊ=ɠ���4���������P;���4���1���2��]&��tgډ��o��'ɕm�MsUZ�ꓭ�
����#�5F�ޜ��=ǻ���D���o��$���[u4`��bI�U&k��r�ՏNR;CK*��i�]<��Ĉ|��Y��\��,�RC{�g��o\�OUTe��j�r֡�6K�r�m��r�9��I�c��P����A7��E�����G3M�)o`7�w
�c`P-p�&��
��d�X/�7e�5���h�2��-��*3 "���VII�h�w�f�#p楐�̭SFɅ�nL�FJ��dcr
�k"�S2��AΒ�w&-S�.�#�~iwwn:�ϫ
n%t�5
�
�!&=��ͧ��NiNf�HJ:M+o6,
�(/���yxŲKp5UY�o^�+f�M��7��i����4=��c��(Ք1�ǮAbj�*lAQ���v�A�X�at�J�tkB%��N;AC�M�%"D�ʣ��+Y�"ƅH��W)㯰��ŗ�2�h<��Gg_�Q�ފ�t��s4(��HNܫ�oL�fY�/7pJ���Q˼�/ l�f%���)����f��܆i�j6��B�ͽyp�Xш�������[�f�n�{���DR��MM�
;Zr���\�u����T�9���t�Mb��HuO;'V(��"7:���Vf�Ш1�`�mnE��*�l�M�ܗaT.fV�YS\.��x�l�M���ޗv��^�Y�ҫ��5l�sf82ꚤ3Mdסcw��d�����gF��BӅR�	�31�����Y%�kK�{���1�&e�K'���5ތz��5��Â�槲�Z�יa�O*�����ޛ��ڽ#qF*^�I���eܳ��v�f�Y�%m�)ɢ�f���6��0LL]�b�.�"�X�z&��f[R;�[��wBq�Oo2��/3 O-�e�T�T2�׉���h�[
�u(ZD�`oܽ�V�h��[��1zZ��ܵL��ᵛ}͞��EƂĆ�.fM�Q�Mb�cEI�Uͩ��ʭ�� )�hê�GI5)��˳bl�v��̂��Iz��.L�rV7���䣘�[Z�2Х+MӺ���4D����뽱Q��u�M�{�m�.F�W���V^��x��
ɪi@�i361�\P#%<̕��ÏvfX%�r��+p$Mz�-ۄ�JP�%�l�1xoB���uGfQ���**F��X����bVL+%j�nm<��s*�ѢL���IW�R�%��IѓX����W�t�^y�i�
��
jSb��pDwT�wU��Kn�,�T���2썖ҿ[�R��iC��H&*��7�4�b�U��d�����*����]SW
5�^���H�D�sV;Z�;�jJ�Yje919��45����"�֍����Юn�$9���$���mWڕA[2m�]�T�̄�21(X6]��X����9�Ei�r��d���u-��)eƃt�-D9��[*��	��RXFƸر�����V"�Ǎ
u^749�hŴ5;~.n�m
�4�M�JȚFX�4�unK܆��sV�^�c5I-�m�fTʒ�#1
6�S$� ��)�S`�"x�ZYJ
(�pk�Ȭ�\r�Q��'Z�\�m���%8C^X,�,�M�v�HIvc�6O��(LW�Zd�M[>���)7.�l��Ej�L"�d6�cڛ���a�����Q�lB�LhPW{&�"a��[Y1=G-^�+%��ȋڕY�{RLY4�/u�+�yg�k0a����!˻S�R��^�d��c�����p�1m0���G�!��df[z����f a�ܐ�'�Z��UO��OFݽ�Ob����u`�F������&��9=&���#v�R�=^i9�t�i1S�!�E�,�rک�`qT�z���(P�%ժ�E]ɎT�앎���jᰖ�X�j`�qk���7Ff1fT�^2�r�9�ԹM]	,Uʷ%���ͻ����L�[�CV���J�J�y䤰r�3��'r�iZ/r��!l{k5 �DN���35��Ru��fɱ��GZ���[Xh�K��w�E]:42IWj�R��Q�oI��9�l]a�1�kn�#sMS�efm=y�W�[�{l�AD�`U�-�ˬ���Ú���ɐ��X��9��
���� �r�� i�Z�:��0��x�Ӵ�1�ׁ��57(�͹��i�u3C��+sX��H���@�ڔ���"�^i%��f,�ΏJ�cM��q��`̭��E�ڵ�XZ�S��aK�`��v�9�L���e�@�n����Aoi��*V�-�0V���ޜ��t�,A��`��[�4�ݠq���+D���f�QP"���iO6F�«ՙ�Ei�6�c�5�ia��D͒n���w�,/eSl۽��f�HIwoN�XW�O��� �Cq���J�S�h_�%�ث�w��[$�!5j�]V�ǡF�ݺ����*��	�]�Z��%�۴����0�݅#Y���j9��{�h�wR[HQ�NM_,Ѹ1nԷdI%M���3L;�����E�Γe��e�-܉d/,���tޅU�A���F�u�b�;9&���#�X5%�A�v��b�,XAy[ba~ؚ4����+�(-�2aj�`ȶ�
u�*�ʼ���f2%��0��iB� �NJ�(���!!N;՚U�FUvo��=9j�{v/z����	b�B�S���J�)�*�:#B�����)]���'J��=��5b��U����l�ۖ!cX8�7��ƩU槆��oÛJM�:��U3!���e���Uz�PW2e"����V�qH���7*�97 jٶ��B;�̖�-���طt�8P���k��VɰtnKٕH�ݷ/i���j�BE]A�nh�[:^Pt��{bS��Ÿ�<sr'$�b�[W��_Z���&�;Utl�#JK��Ѷ4\�s2����[8������z�G�x�4��jHE'N�׹)�K8խ��ئ�#���73�Y�r�Qi����@۶�s5)����˼��
���M�[^rZ��m�Z�y�YQJ�*�v�E���^���Z�*���$�u�'y�T�J4E<��9��n��q�ł�+�ȫN-�a{��1�;��1)7�>���x$q�.ɺ�[	�՜N���9x܎����vA�u�&����uʷj˱����V;94�tJb���`��
�-�pd�b�s��,%LQ�횉��d��Zf���QL�n�����m"�
�R�o!i�{a`8�3�E�䦃K㲰�M�:6�.}�Ws+��y����p�MI�w����X��ܦ+�@�G����W�Q>�U�4���RirF�jZ�,�5p&,KyV��e'�u�=�f&YA:�7&gb���K"�Rե�� ��5���o9�Z@�[�һE$�ijبJ��,�w�v%��)�d^(��ܓX�qu)��x��K�|�U���KTJ��KUEx��/�@�#JD�vŭ�Jf*����ȵ�U��y�Ti5i�'���k\�O�˳sW4y6�Fւ�Tӈ�}�	)cf�������դ�%�KO�c�N��u=I�������b��sU���%��TT�Xz�Lhڤ�-��T�"֥m6�JD�w$%��mj�rF�&i/��$�)k"ĒE���U�uV�ȃ8�O��R�Zxi3�b�TT���v�Lk�a|���a{%v�'Z`�
���%����,�|�,���ڵ\�*��KQj��o�Z�O��m�������WũsǮ�c[��q��mNV�v�Q�J��D�Q��1GTk��5���r-��ƴ�Z@���j⤫��\��Y�e�����+u*֥�e�[�u{���Y��7�ڨ�<J�@�Z��]}�qMV�qS>ٻ�뺦��];I{�UZ�R��;k9h=����mLR$�K��Ы�$�.y1 �hTX�����n@�rF���,R��ZƮ��[IꨤSf���%�f��hĈdM,��.U���+��i�ƒ֕%��v����Qĭ4�Wj�1$�KVjI4��!�\�Oy[վ\�j���U�8��qn��j�ى��R���w�]ir�<"4��^�i\OR�"�'=|����]�TT�-�Z����r��һn�&�r�o#i5Z�TĚX�I�j�K�$�0i��b<�'��T�K�E��,��=L����e�K�WkR�:6ڍ^'j�v��b1[J�	Ʊ'���J��HI���&�R1dZ�/6��ɼ�.�dm+K1LZ���,Iji7�wUSO*�-I&��Mwl��KR��v�<ڵ�7�:�fu�'yku$�UH�9F�iEH�Mk�e�5T�x���It��6�,�5�UJ�X�;O�����=��~����$�G�~�?S�I���o�"�3�3ĴP��T��a0���d�k����.�dvf�L��W:w��t���oeU'7vq8aҏ�u�x�����1+E�cDSV�a�)*=1�}�ٹ��n�.Э��r����Om�a��wY!k���<�}N�7}�%^<tݨ��5��
}wZQ����zgwZ3:}-�6a$����ts���TO�e��f���?[������(V�o2b4���f<a�.�sc��]���j(��f��6c}p�+7�iu�T=�zvPV��C%8{*nɷ¹Zڜ�-l_:<J݌�]'�Q
�H�u��;�E�Ĝ��\��o�S���U�<��b&��-�����tj���j�צ��xSl�{ZN�!�[]�}!'#oM���>v�/*zi9�
��t�w�kp���Y!6+]9���>NaR��UN�)ޭ��4Nd��f�@�L���oN�v�4\z��+y�B���x])H��wѱG8�5z,5���y��.I������E3v���<�b�k�N�DI@��ġ�}P̴v��_n����.�K+:gt����,-�ǈw"�C5�q�כ.��I�u�M-�T�/y�d:��um�Q����g��:��ƯDi洋�T3T��=f�uY�o���w����	�L3��;W���n�T=��)���oOH+���ɗOyNw��m�MZ�;θ����Y�"��˩����i"F��D����˱k
���kw������-GɈ�-�|^�~��Q/.�Ap��\�)26���nJڠ�sՊT���iU�������,�Cs�u#������RLZ^iH�{7�o4 ��Qv�d�U�B����<u�1w�1�AQ�/�V�&�qðR��$�V��y�*�bX�����Ɔj��8����G�mp��eW
�Ɯ�����o̾�M]��b�k������K�般�9y��גK�Z�O��:�j���:˝���Ms.��]��o홲�jrHcUå0��NM�nm_k�#�>�ϩ㭺W0��MD�]u)+��,�ՎUZ3�.�=�n�Ȣ39��E����K%X�(T��-ኮ��}��᮪�L�ӢWN��b�.G�C��:�;�湈�����ٛjw�0����u����m���Ĥ˝x37���{�.ܷ�����vX�T�E�ku�'�m���l�Tц�vK��)͎eg�Z�YCv�&�Me��)��&V���{������ʉ���*ۼ:1��{Cz+���[�5k�[VӶ�)�2ii�F�f�^�Κ�����IM�D���i�^��3{���s���q��oa���`��mM��
q+��/f��ە�on�Vt�	��`�!STp���Uw,����6��ד4�XnJ̈́�#{h��dI;7�������#VRTR�D�\�B�SnV�f�w%ͪ>�x	�b�cKv�Cr����z�UFd]�G3�k2Yئ�:v_u��#�'Y����Z�Цp�K�ϘŌ�vz�tȊ��������[�^#���J-�^��0���r�j�r�kʪo(�Y�z!X�%J�rd<��K��̳c�; �4����g-�19������C��mq㯺�8��m'}�R\�R��qmfH�κǯP�n�:o(�v�8x_<��7���^kh6�����a�Y=������Q"ƾ���D\����LM�*k3!{o����v/7S��&{�w͆�菣}cV��f;�Ѭ�LH��/�P`�u!��λ�����;U"��S��T(��kz���S95��N��E��b'o�W]�q��j�9W��ZV��.�G�~�F;�޼�*̳x�����u�Ok�v]�̒d��l��y��Y�V���5ة��ʁ̤����i��t.��g��?s\���bY|3
d*M�v�l���T��i7Ҿ�����!�_X&��ǹ׵ĻJt��]q�OV9��ԯ��2�n�!*c75�a��Ćܕ)�f�N��6̼
��]ՓAK�>p.+0�ێ�I}���%����x�����NH>�۳\�rsC2�_
:#�_&\��:��u���,Δ2��s�5�1�ݑ|$�v�#�B6��m`�vK���D�8:5-O��58�UI��+t���%
�J����5��zge�N�C���.S��b8�z��!������@��.�q�ofSgl��́E��5���ą�j�ԧV��88����bZAy�ֈڔtT�U�uWv+��,:{)��B[C�].��j��C��"�L�:�6�fq�[c�i��3�`�Dr�(���7&�6k0>�Q۪*Yؔ�%�6�}�L
�t�1պaR*��h��oI��V���UW�U�j:�#�u����6*Zݫ�s�[?C�,�i	���H�B��r:�JT�\5D��w��6���ngԎ�zn��M|��Kvt�"ðL5���ș�V�"	�Z8&#���m⺈!���-Y�tKw�n�󁤝�S���;%�S�񬖙�7��hU��9',��.���WXWPD�R�̐�1N��jL�tU�<rheXU.�9���sT�[QҔ��*�t�ȅ�;��L���W�u�|��}v�����TW	��{e8���Igi��{e�1�`��se=��\-�&�P��%rX.�Sw%�UH^=��:N鋡�|�n�����k`q��[�]N�j�u>&XTp����.sAy���e4i��E�T�|{[��J]R���_<ʜ��8c�p���R�&�����?��gX|L����%$vV&�B�u��a�4�gRi ��k�^BL<�u6.�P�t�m��Y�)?�8��핻gp�5*�����hӝ��i_z\��Nn���F�Gb�-�0&�����W̤�G��:���E��b�s��r�#�U��Q&�ٛ�>*L���0R��j��$EU��\&��[����t�ﯦ��q��N�;A�vVpb>#���5����Y��!���b�,B�9 ދ�j����lxqW*����L�-�v��1��ޙګݬ��b����x�����r�m]߁��2�c��̅�f�Vt��q0ʷ�k���qV�o)<��u����J-�G�5��-<��-�7c\�����K�=XaF�ߒ�]ɴB;ÿ=�d*���'ڟY�53*�s�l��,r�/O�;�|"�r]nv�a.y���v-sa�.QַEZcEv��D�,u>����ِT�G�ݎU�`����(����z�7�t�:-�l��t׃�]u����4�P���'@X���NB��wgF����L�5Qf�严���8)+GC�o�"W�x���8����n�T(˗�����$-,�,U��a�ј;��=>J�	;O�J��%�*erFS��3{Gv=:�eg-�*�Y�Uǖ�fゟ2y�����eC1�=�k��s8#F��R1E2jO�f�����wyC�k���}/�a��U����M杖v�PË��=תZ����KΩ ��-��Psڎ;�_X�����i	�;���vyv3��5�N���3�yx�S���q�XBP=�%wj�gVlR���N5��U�-�ɜ�W�4����e�z.�ι�����9�Rz�t��k�cexZ�FyD�����7�I)p�gm��Mb��+��WEe�ZX��7�CA+eY��k��#���y�R�t�1�R��x�t�}�Ͱ�
''/��̍����M�oz�z����u#��yx�m�o7(��5tm�qt:��jJ�a:܋���h��K�9��-OY�g�"�V5f��m����gs�^��N�(h�j����}(`�a�Bb��6t�
]�(ug*�*������i;��)�o���ࠥ�Q�E���2pu�'D�#[��<Q|:�{�%�D�m�h͵O]D��`�e�y(0�'����Ze45�]�;M��AƜK"�w����w�>��켵��^I�\����0"�:htb��u8�D�IΜ��;p);x㎲a�+21*�/ Z�t%�˓��议�g'�1Vʱ)�e3�#�����:ݐgnװǝ�.E�bv�΄;"�w}HҜss+5N�n�eh`k���j�ݣ��v	��qs]�y�����CD�I�t^��9,B�k��Ug�oOJ��ݵ��9u����ǷY��r�z����ʠ��m4E��4jl�9�H���%ПU�������3�}�	5ń��t��҈'�୉쩑�;BJRƅHq冝�킶�N�fh3�UX"�t>�_�o(J�.���=U�M쩖k<�=�I,9�:�Fqc�!|�z/d/�8�6�顺�-���.AT�*H�����k ��6�N츮��F�X�X�=:�1��qu�T��Z����J����K�B.�.�p�癝�����4�Z��N�J���7���Ժ�LM̕-�u��Ό�I ��;]�mp��vS)Jǵ��o��b�lj�X�R��ճ�]Jq��k���Xb�� �1��m��v�[�bݤ��P5�k��N���pg�R*����U��!�-��Gjbtyuʱ������ϵ�3�=Q�d���c��n�z�&��c�����p�:C��5wF�u�T�/��VB�4A��:M��?���G��C��f�U���ٝU��=�؄tm��Z��yWq���Ɏ�wwG�9�>�;-e:�]����ò�^�u��V����7\�%�m��JQ��v����ˮ��q졗�f�%�J+z�*�;nSvu��t�����u����*�
/sl�~��T�E�]jl��CkB/,۫��C�Yi���[���םۓ�Mٛ7��Dr�X���*�l�j�F��ed눇�n���וV���Q��;�2���U-WsJV�MϝO{t� {u����M{ڒ�:�4���*�W���õ>��7�Q�.j*�ֹɭ�|�N�*fhڜ�__>E=X9�y�@���å� ��XT��c��z�\��N�k��{"��'�t]6}�86�l��ڨ�Y�������=z��6���1i���YeyfQ�~�9��w�͏��x.�zc4�t�#y��)ݽ:k�¡��q�ܹU�аF�{:��GmTDz���//�Ӭ��NCe<&���D�W������l�Z=E��z�.�ʻҌ�׃j��,�7��ʜ53K��2d�]�U�
�b��J���զf�%Ӻ�\��t�Z�/4ۛ0pc{l\)�Ӗ�6Ϊ��^TEj�尥}BẔ{'�n����v=��;�JCfReKڭ�2y�*W�^o.V-&�l�X�ƒPc#��K��Nu��,%�G�9���GeN������F�P;��D�ʱꥯ2*�N��w����s)��y2�A��k�=x`g4޴�9�v�x��o;��y���u6��|ET�$�Ho������h�gl�:v:�$��5fv۰�\%��E5F�7��wc6���JfT���l�N�Ԕ��h:���뻶8Y��3&& �8�:;�U�V3)�}�s�QUr�g����+�-�i�eh�f�C����bF�J���*��e
�a�"Y���!�c�ΣN�Z�}3l0�|Y�k:�=C&��cTf��WAO5(6�֜3hr�����3�;���5��$D����Uz;$�hN��N[8���`|n��*�mgY�t���V�$�!��E�(�g�Z.�˝Q軡��ݱ��KMQ��_Rq2��Vs��Ur� ������v�3f�u��c���Y�uٹ��o]�0i��^.Q�6�;_]��o�7_Ҷ����_2����ܔ��xY�/��n���۝�$ØI7���@vPa��JJ�,���lX��똰JuNڲ��8����\��2�2��y�yq]G��2��u!�;p����ыaP��r�CF����`Sq�ys8����e�/�M�MϞI�����c����m�fǲ9r-;�˻÷�7���֟N�:�W�d:� ՚�AOg�� \�n��|�=���td�"d�sg8z�'�(�\<�˻| �恘6��z�g;N�/xm�]eX�!,�AxxEA�u�H���A��r簯k�P%�}�Z��\�r��$ȞO`̀jj���j/|)�hRD��A�5+)n	�S �	U@��r��C٪�rn\�{�CY�D�P����dU�zHq"π� �V���DS�{�����0� �OpX9��g�>���ԅ�|��W.�Z�H��^�Ob�y�Ӻ�M�8@9�{A=�{�H� ��?�_�`�(���8ϟo�b�����~���"(#������>ߗ�}����������K���]Y��O�Xlf_�ZI�<�[b�ۆ�M�+�2цR�T#��Pwj	ͧR�k��m$��˾˼�"�c��inW�_\�����3���\7�G��F:;�y�d�Ѫ�o�ykm�9���w1:˴��`��V�]�Db��d|��
,�����6)�O�N<)*O&���,ZJ��|����C�]b�/V���LT�Ơ�θ��ّ;�l�[]�d��VTt"��n֪���@�������h�sY���'MMGN�t��vn��w�M�;Hq���ӘTj���r"7I�`�i3��/��O��H���3�^}�Ş�À�S֡��f�_�nu���ҁ|F,�{�\	����ogV��0�n��d��[K3M)���u����Z���9��gj)r2�	jI��W�2d|���d��J��C��F�N�S���e;m�;7d����B���ʛ��Jg��ᏼev�î�V5pH�x��%s�=��[R��MO���h6��Z)�5:�H8E�`��Z{j�� Θ�e*��lؤ)Ѧwg�����O{��U�T��[�)G{K+	���L�e��S����7�o���rn�����o}x�8�8�q�q�x�q�n8ӎ;qƜq�q��q�q�q�q��q�q۷nݾ�}q�q��q��q�|q�t�8㏮>8�|q�v��8�8��q�q�v�8�8�;qƜq�q��qӎ8�>8�7��}>�?�峝�'E����B��3��s6Qt��BI�r��/t���l8J�q+�Jy�����pق�n���9�Xj��S�ݞ������風�ͤ�,���v2؁�]�찬���$�Q�g���c���z���n�+�w̵�fj�&
�P�VW����)���);���N�Υ���/�)WgT
4����l�d�,�WI�S��,�#,3�u��*�3�XH&h��N�5�S��f�N����D�ڹ�[�\�u��;��Z"�;T��0��A�b��"^�7U[$bc1g���y�u��i�h��r��h$0��2�f����CO �Υ�'3y��Sy�Zr���y&rLU=�'5W�*k��*�D��gg\���WPײ�w\�q��7α��a�U:N0Z�p��7U�)��%bq�M�X(m�2��ֺ�T��)��m�D�~�i�"�j����Q�In�΍"���q���X��DN(l��pm*F�ι���;wn���z�Q;p��t8��M��${X���ރ��۾��W}�A�/p�ڡ���M�[��Rs3U�'�ΰ���������;	n�]D_b�O���b0��2{��̧��A+ޜx�����ʅkB*B�+�j�۪}|t����q�8�8��1�q�qノ8�8�88�8�;qƜq�q�v�8��8�ݻv�۷n8��:q�q�\q�N8�8��8��q��q�|q�8�8�<pq�q�q�q�q�q�q�x�q�q���N8�׾����~��9Ƨ���aQ�ە-� ����^�D�5Ե��5��pS�Y����L��S:��e�ǜ��k��e�m�$�c?v�;�r��v7]��_>.�ѻ+���W��m��O��]a{Vr�+e����`��MQ����z���|�/����Ss��1�٨��v�[�;�N�bJ�^�a�T/[�*�*ŧ��j��A!��u;�]��pv(i�0"Fa�1]󀣌�n�swG^�-픩�f�=�(��v>�P>�*PWė��Q�[7)��Qu�T�r�ŔkbY�i��8�G9!�UXF�T:�QS�.4x˙���F��'V�Ei�ꕇD��V�|M�۫V���J�D�s�*��h���=-2�fѕ�[ N�Ӻ�����"Bm.jJֻ�5X6ِWP�&��Zx��S�|5R�6�%Z�w{f�PP��&n�.�v&�f^�Y��-Ge�M9�|���u�ޗ��J���z�����v;H�sD��YFQN�b���o�ml�9�uH�aH�	������Zg�C�8*�gA�.���vj�ckjӫ�
���HՖ�F�B������D�Q�v�uX�����n��_)���U�Y[w�w��������x�8��8�n8㎜q�q��i�q�v�4�8�;pq�q�q�q�q�nݎݻv��q�q�q�8�q�q�8�q�q��t�8��q�\q�8�8�q�8�8��8ӎ8�8���q�q�=^���{���ܴ�t��ʮ.���!⪰۟*�f�pЗ*��ܫZp�tÙ��vL���yp]�\5�o���~}�Y�6V�FG,�U�b0_���q:[m1�F�V�n�/(�"���DC�v]+E�J{W�U8h�������d��	l��h�%�,V��Iv�2ww:+��'#{K��͜�ۘ�}��1Zfαӯr��vp��T�÷)w&6�eo�y+Ϣ�:��uu��6��{P����'��.Ԍ˙��1rUe��9x�8�Y�;x�nӱ��,�ϯI��D�UzbCp���*y�+���mT�U�TM���a�G:��>���pF���C�t��1Z=�~�3�͹���V-�%ñ<㷹KjҊ�HoE��V\�nvҮ�����J���˓�4Y;��lAZ���ɹ��
���m޾ܹUȍu:���gRcoD�Z-.t3G�j�I�xr��9�˧����^b�_ 4�Y�<��M*i�s6��n����qW�I����D�oA=#"����{z�yu���m{�� ��P�a��.��靫�os�Rr�Q���,���T�%�V����'R-�|(h��[(m>v�$���Y��kb��Q7����һ.�\T��,�PAF	�d�hgN���7��Ft����%��D�ܬţ{��}׷n��pc&gs��,����u����ރ;��W������8��8�n�q�q�q��t�8㏎8㍸�:q�q��q�q�qێ8ӎ8�<x���v��q�8ӎ8�8���q�q�q�q�x�q�q��q�q�q�q��q�q�q�q�q�qƜq�q�n8�l�j3�$��^�ò��ձ��A(֊��t9��C�|��Pn�Ib��(�u ۾N�J}�$�pd����V��[΋p�K1k���@evj��ҭ<����6��>����w�6)��5J�0�G��l�v�,�,�9Yy�/.�<r��6ڪީ��ch�'(נ��W���f)��$�t�> h�����<��n)�Խ����ıwִ��3賦Sa�0�C�����{rV+
B� {�����D����cKRʋ0k;���p��a��ܾܱx�jv��e�8�Y���ZZ�p�����Y�2,�f��U�[гz+z�2l���+D��yx� m.ܗ��Y�	ҽ�1� �2�3�W�;\z�d�ێ�4�K���b��E��'g�V`���҉QfR���W&�\��x-�*�\_���j��7-�n��ҷ{�_/c�#��XG]5&��|7OL�r��uW��N� ���B��#�on˝���s!ʆH�aO�ѻ�2I7f��.]0U�]k��>��e9Z.VcM����6Gz�h��hz\��^B��a[�������cAH�v>8̥�[D�y��5�,8oώ45q���|�@�*��,^�nk��L�s*bZ��:�f'0�BS���9De����Τ�������WQf�\�n�Cs7�oq��F�<m�:����rck��檡%ҵ7��"� 2,�\{����N�u�2��9;��I�#�㹷S��kF��|��d�,,�FOK����mjYZj\
���m��(Mvp�n1ͥ�Fnm+|N�F��y� ���d��:��[z��7����kU�ӭ��,0%����%EOno\� ;.vo���!	�k\ȐX�[*�fPܴ�ʮF\z��`晼g:�Zz�Fp�tɜ�b�� _f˔�������M�-�ͻI�PZ�phY��v�f�w����� ۜlzD�j���UQ�w4�i�cṅ#�Kk(�K1)�֨��ƺ�p�X]�V��pz��l}2�>r	��&���
k�Y�U���mk���":��n�9�i�k��5Ff����5}���Q�,7��{���g"#��*��o�VgA�I	��MՊ�;*���+����EN��SY܋v�(�
K�iI l��eAX1�yYOv��V�q��^鄛k\���˪�g-���Z:S�UĆ�n ���#�s�#���+�0-����2��EC�,���u]	��Z���o��I�X�K�Lr���p�l�]vS۲^�#��#��f���F�1:i�Lc��/X�@����;p�S�zR�pڱ1a�wt+5�+AD��VjU	γ�YnKp���H��f���=�9u�5����U�Z;&C�����t;����ε�U�����ת=�(c�u=�Y�'���FiZ��h�P>V� \j��UE�j�_h������z�\о���{@�T��"Uwg5�ɘ.J9徍̆l�-�ԓ����鵖�oM�j�^�ʴ�Iu'Y}�y̱tM
r�M��p� V��j��,:k���}�E�v���� e��.���O2I���n�9��qd�K�7��a�j_K:wp�O{��q�8�7�18VJiW��9�-��%���cWQM��GP�gpA�;�n�ol�m4�i���y�N7��D�[����[Ŗge�����o�U�i�r�;+��;t/��ڰ�������Sk�as�wC7K����z�an-U�[O0��o$7ƖU�V�L��V�:�q�[(��ԧN"�\h�N6��� �ٝj����>���U^H���JG�VI׉=�/EY7�je˒�
3�mb�p�е�ayUcf\�����&ﵶ�R�y]���\a�{1��&;v��:mΩIip���9ɘ���L�q�2�ӣ�J�Uy�$n���z����34A�uϳo��V�QY�2��n���+��R�*g!�ջe�r��u�p�u���G;R��ؓN|f�kvi�tV�N��]c\��}�d������ڥN��z��ud|���-�Y;+�i��2%}�-�d�̓j)�5N�p�On�NRO4�)�A/X%��mmV��P;�I���]�TfYw�̯�eB�F�(!�7Q�W9ڷ+�������3܏�;�;1�w0.�yN:h��7-+1*���'�jH�v��&+�^e28��6s��.�,�RT$Ȓ�nB��cf/B7AԷ#�Vu���$�bH��O,��hu���e��+�Y��-��f#�vA�REw�jb�ӭ̧Gs&���N���$���ܛf��?�q}�z���#�Rp�s:�mAڕ}20��yc{t��x���(��RGU��+��x��!��(�cF,X;\�\u��Α����U��CT�ZC{��F�t�u���uGc܇t�&����,'5�z	u!�jI�B���]�Bkf���}��
�ǨK���Z� ԩ�m��b�x	��e國�~��}��ZcYw��h�W�ӛ��E��'$���i��}|�k7��,&J�f<W9�_^�ժ�LW��S�����'Z3��¡���;��mV��([+�!����rs�n��YfB�d;ʙI�.:,p�yWW\C``�4@�̹Pud�m.��x���r�g=ڱC5�ZwRoBO�8P�`᪦7���t����e9�?]�$��ݍ=z�U��K�mڇ���wV�b�:�SJ_gI��"�:�m����V��jp�
���9���55Æ��aǊ��[YP�Poj�9ϡ��W.�Ty5;�8�m��[���Xk���������"�X���uj�_#�]�N{\�4s�I}��[͡<Ӫ���`��5����+.�,�ɺѬ��G;d �'�Ν�!q�o&�h�VE�#v���Ƥ��-ne7��;L^n��`����帽[8K�J얖7�Sg)��<뼟5�X��l��VE4J�m^�2���`�=�4Myx�C^5)2�cID�c^�ynM�}�쇟jʢ�Wf桮�r�|��;g(�N\Qm7lc�B�n��r[��v��������ݚ�ln-�h��=���ᾨʵ���1[�ЮI�k����P����Z먟,n����sul�A��:��d�}�{�>�g�Oj�6���;,PK���݊�7�t0��6CV-�d��k�]1kfv�����K��jC;y�q[}���&^5&^G%���ۦ̝5��J�{|o�����}��2ʽ�r�$�}TRj�8��kg��͸�k���I���F�Ea�[�c$�2X��lm�B39�3�����&�*sh���(#�9jax����e�)�ɜ����l�Z�Ub�8��qD��icM�ĵ�g��� �:��Ř�>��G����n�[ ���{X���a#z�]%;޲���Eksv�]Ε�+��l��Ŝ��WW�'sh�&:��/�0�j�b
���]E��N<��Y]�	#���U�i��yxԂu�<27Gw� 4�Hw���P�H���³_
2�w��[z�'�Qu���q]�m�
��H�@:v��׻eM��Krl��vr4�ۺ�>;U�ݜ���0�rG��i�@���Ϊ�,�F�=5u�u7:&�x�J�tf�m5ZS�0�(�
��Ց܄�mp�jL�Tl}%T:c�U�:n^��uW-]�b�1J�9����.��/�,�cz��#}0�\��Ǝ㈃�1_���kiKcfU�`�4�Gp�\�b���٫��&PL��k����iU<�cL�+ɘCi<;[��V�v�ڨ���Yo_�-�k���㢱�r�vV阴�mJiP5"�/�?��� �����/��������������~>I��y*rM~w#��%�$� ��!1�dM��q�4C�e8��6bq�!	��-l(����R�S���L�E�Z(��,�.�
L��LF	�4�H���A0�����T������H�q�R�4$�̑�UHTb��P�W� �?�Ç�xm�~&b9 0ʦHA�F�`�Y!���P4|�p"�Q(YP�g�A�5	!Zf8�26r���v���6b^q8��e3t- ��L2b$�i(�D��i�&�t~%5�O�7�\<'t�,�wk�*���iI�vj�8��5Q��j�g�Q�cyy�DV8NT���#؋��T��]�h�ܻ�o^!���,TA����N��Y�Ҷ���V�u�N9G���/��&a��j�;�)�m�+�G��q�(�pB���!糗pr��&儱֮�OCDa(2���f˭��)
��J�U��C9��ՙ��&�w{�#�i�z�)�Yͼ��UFC�v@���-A�ڒ�IW>�r���Li5������K��Xbx����NNo��0���dEn�R��y��9�Pws��mHUVgy�����F�8�{7���3�f���v���<���
x��|�-4/z/�x/�zV��E�ꨗq���]XY��׎����¾]zkp[Q�]Op��Os5��}%>���"	����H�ܦ2��H�Z´�]�v>{RoGC��s���JZVH�{܉�EZs.�զ�2�L��j��[��T4NO��8qt�ɔ��1��.<�<^m=�D�4k�J�V/w�khR�+����j����)c.Ƽ��!M�}�>�s�$4�����Z9�j�ݡ����5
��E�w�m#��5D���+2t	R!�l4�E&+>� ��*
�?aA�ׁ'ѣG�(	H�I�J��1Q�ۄ�G��A�0"\ Be�FZ�[r!���M�8�j�4��)cNKQ"�e� +�)��fD8��jH�F$�D?|�q�ߗ�0��n�m@`i��L��!d2�F�~��T�L��F	⌍FJ�H�*�� ��n� ��"SJ@�n�l��-�Aq�[@9�4��AO4TP@�ID�	0Th&�o��A���� �^^���hF�%"[��H`�Ҏ!��!H?Ca8Ir	$�b��FJa��E0`hDQqG,B�d/8�&�1�	���jNr�i$Z!����C~15�@�i����*Q�� +�)����A�Ӆ �i�J�h�cr)"�E��0Be�%$H6�`H ����A0�� �i8` ��h���
��P���F9�"�"���-@�i��I���TL���eC"����z�]s�a�y�7J����������w�� ��g];�"S��^;v�۷nݸ��ԕ{���78:^���]���r���{�E�٢_�_>t��B�I$*�i�n8�nݻ{��{�}�����;�p�
��6}�y��E�v��\:r�(f�]��w_�<�]�n�z�۷nݻv���ǙRT
�J�R��-�W� Bd$�	�i4�C��6�ν��w+qݝ���yޝZ�^�u֮�w���nt������[^��w�gum�N��M�z���nݻv��ף�E�/�����&�����8�[c�Nt󭨓wm���t���cs��=ݹ�Ow�:�V�k�ow�Ѝ�{�{�{{���]3�v��ݗ�9�yv�9{j�q���-^���t��������W�{�q�ݪ��gw.���z�u�a��	$<�i�H��M���'���O]�������y����L�l�Q	#�	�Ke��6�	W���w��gOz�޽�$>�r�2.��ݽ{���]9��=���N](��Țk��~엝�v/��۝�ۢ']tHf��D)��]:7n�s��J`�B\���<ܝ�qt����qB~���=���]0̗��rM�1~�;J(��1RP���G7�x3=�~I3�P�RA��h�*��B
�D \�W�rD�P�F�nDI������uM�S����Ea��S�B�p9�<�N��t���$�TJ#�Dcv�4�2wF��U"���ΐm�!dH�1��"� .
 �Ce�a�.�"0�l�	H���[�9#R2d�̐C���!�������$$�����R	N	Q@���zwZ�Zz<sd��G�n�4DZѥv�-L��OM�����b?�w��=K���~՚߶�f�R�=[��������ɉ�#������>�\��o1�nlH���c��2G��U^���,�=�A&�߆ϳ`�I/�D��5���n+���{Ϗo���U���A�o�Kg��y=�ڳ�˖��l��wI�k3�6�)�O��96j"����Xˋ�?-���}�Qg��Snα�ޖO�q�"��Y�ތ�6�!>�b��9��(�����kj�D�~��'<:������>%���0��l��lc����a��O=��g�`5I{����-OL�)l	�ϻ>��u��K9B�����OݜCG��1��{l�)�d�m���cޓN�� �^zki�(�=��g�������T+��A�fE� ׵9ƼԞ��
�SƇ3ۻw�$]v�9���Rv�����ׂa*��t�\�p��ɹ8�E�2t�]U�6>�"���E4J8Vi��R0��zBפL��.V�I�;����h�3�ʎ��#����GZ��)��m7גu�d }'a���9˾>���E<aY�]�=ھ�+�9̆��{#�R�۷<ty��0<2;�@��t��׆�=�������&5j9��B�g��o�{��TϤ���Qg��С���¹^��r���{�F�g�o�������;jH`�[�6�����f�4�TU�p���4sa{��^і��_�������EG����i/];��_��Q�{�7B��܏owH��3C4�|��͌���v�1w�����>H�(/	�/�mk�u��ܸ��{��%PI�]{n�X�Q[͸�{��}���^׳�``��Fz�/��7qV0�WJ�{�������>���o��^�;�:������� �Y�6�{�`�웮汻$�c��^L�v0e���"�:y�W/C�ף�[]W���p�Ŋ���	"`H4���oN�>}I�e��
㙕����4���Xԭ�Vo���R������̭���<�͋c(3u�f�t�?��/6q�?�g��[���SAV��m����B��"�8 
�]���e	�T�;����S�}��;�ަ��)�۰�X���VG�}=������KF�K�;E{�{�{�_��t��X���yk��Oz3��Q������uY뻼��5���\��I�Y;�OQ���#�S*}�/���4�ޒ�P}~�m+���Y���\؛��{����@��\w�3Qs����ċ�}eЗC�E�7�k^��j���]�]���y�`�{�G��Ǒ���A�*�hiJW��c��d��ĉ�z���Q�õ����>r�h��=~�+=�����3��}�A�*�XV�����	?��xg�����>v����˒�Lܠ�p�"��,W�'����h��,��O�N�ıssj��"^����1�������)�����u}��n��~�~x����
��NZ�+�3�����so���-��@��݇8�LU�Ȋ0�i<�Z�y�����������Y���BqCX��N�o�K�����E�t*��r��_�a\f� �sZ�����ls��B�R�.�O���#ݒzuE4��<<V����5��?b��UI�{%3����b��}����7��`xK�f��͚�N熿'~��z���getm����	�n��v}���8m�ޅ�zI^.�m��0��|��}�'~�u�By����֓r�U�[��z�C?}]׏���\��g�:Տ���&��P�aߒ%zR�T\���\!�Ƞ��F��o�y�����m��*��ۛ�]�kx�*i�U ����r�|=��M��W�>??�W�ت�q����u�T-����}u�T	="���F�d�ةg�/2�,m���U��K�����Q�ߔ��zC3�,]��x�@�����r}Y.�Cu��a� a�Rza/�ݵT�qq�3q�s�	 ��k̽���RM�\�
�5^��um�Ϗ\�C�C�k/��'d"�˷y]>R�]����z$w��J�v�����OX���؍���邙��m��+���T�ZG�F�'g!���,=��Y�1_|%	%��>�r�ٹ�1q�PjM:���:���':Hl����T��v�y��I0�2|����:���j��d�}�JPS7;μ/���!}�_�ʃ��y�![�1>ݯ�б�.��|�� �
��?GsG��t�x�l�����j*��#;M�Y����ē732� ���&�=�\��C=f�^,L�&�0{�E�7�sۓ�Ľ��x	����cǣ����'X�3������(`��?R!�� )�;7č|&Ep�:�K[�h5]��N"��d�ھ�#�2Z�ll�9G�=�i�h�mɋ���
�qo�s\�=�n�)��}=�b�o4��-����������.��t+�߯x>be{����٫�jt�xI�͜��̑��G�^�[��y�!t�KG{|��X:�
k:��2�x�no/X�5=���:�h�#�C��Ǉ�T	h�V"��
]���T^�[t��c:=:��xVf�)9�V�:-D���s!������c��9Ȯ�[�f���SӒ籮�8�6��Qӷt^�!xb��k[�y�5]|��򩣒p��Z��{lou�Y#�j }W۸�.~S���+~ ;��3���<�l�.*A�9gH���pO�~�&}v��p�&��za����;��{�����&�6M��e�1���b�f(Fg��&��~�}&�y]q��^�4����l�0;��?��!^��u{}k=����D:��p�<dA.��<��G"�|���xze��`�h�~2��x+p�$��{����̜�3s炶ưP��$6���J����(�]��u��VF��h��a2)
�>�y���Iy CqY�{*���g��Ou�>�z`y�N��Z:����#��M��k{��:��,�mO,�Q�u=���b\��U�^�lNz����l�]<{��5�a:�gt�p�4.7��nCP���N�����z1����H��	���Qo�*�;�2�[��XV�OupRb��qù�|�ޙ�k�^�F���-�GJ�ݮ�:�<�m��|M�ZZ*Q[q٭�z��GF�f�,��u�u��ᩔnu_K�pe��T�,z����2�_Mxf�2.s�֣���-���	�:��q�;��[�:v�F��c���������o�.�zZ�ҹ�qN����?O>�����z�8lc�Fy;zm���WY���s%�>�G��v����SO4�7�Nv��;9�ola8��w�`�^�f���Ӏ������������=ce���`�:]�a=ދ��xp���<�d�6��7��s:l�Şl��1�f���v��-¤_�˿"1�W�
��<~{s�r���o�F��Y��Mf����}���t�f&Fb�I�P�Pu�{�5����M�7;�\~��C�V����
�>�����A����J�yH���e
�u֮�x]�v�_2n?��s�E,}I�
�x�tI��q�I�&�������FH�_�	=�Es�+����C�����k��z�3�J�2���F�|��T\��K�5j-����Ŏ�kJ�/M��J�WZ;>S�k�\:l��k�{��5�N�V��u��^D���Н�Q��SV�컹C`_a�2��G
=r��6w���jVی�����铬α@=}cv�����*B�y��o��}��dM7�E{�[Oe�}G�+�*�cw��]ﰰۊ�\�J�u?�6������!�ߎ	�$��ΝP�^}�9fE}X��7;�9Z|��tH����mz�̄I�o�z��u]�y�6�a��f�U�p���x��y�8$�d"z*1�n�m|=�FM���Xv2�L��x׾޾�	��}��9��μ6�;U�m��-�h��ë7��f��Uo���"��]���k�5ę8�y)�>]����`zS�G'�K^0�=��ǧ4@{�I�s��:�vcbmϲhY}���'��a�rW�4t����߰�Y��VZ��6-#ݑ*�}��W��މ�B�-�?P@�~c���y�#�t�[�u�^��{�Ũ_����)��:��{��Za����e����c#���Q)(�d��V��1m��:r�tff�z���;b���6�z�C2�w�,�Mʪ\�[�=�-wi(Ⴕ��������!�`���y���5s�پ�0t��Ւ�N�̪vo4�t�Z��֝q�Vv�E\�^UZ?x�;�D��^z��}]�R�U��z�T���;�L���$��OC�ng�]��N����$W�:������A��_W�'�g<�Y��E�����<��X�=�2�j ����li9t_�{9���K��1Y�w����ߴ��g�s�贈�K~\�o�M�QH`�P8���6����fV�D'F7�+���=��}��K5;�c�Zڡ�~��g|��mVc�ؾ�h+>�zrR��৬`��N�Y�G
�xl��yM�/g7��V`�Ml֛�Zk�Y�M�'������U����-���(>���B��R_�n�`��k��}�k	�MM)��kru.[�n���ڶ�S����5������6���n�Y�e�&�u��G�\��߫�^~"�6�U�I�T�Y��\�:���׼�:˾�����<qv����W%�Pm�sI�c�[��qT\�gw��M��s��l�:�S��WF���\+�����<2��t4�y�7�>
�[�b�[��>7V�V��PT?q�BMϧ�6v���U^���wR�X���V�5_����(���!���B�^�E�@����]Z���ل|ۉ��vbPg�q�Xi�N���J�Aǳ�q{Å�<U���HQ���%!2{�VFg���}<���&ϻk��8i�w���p"<������1����c:�c��3�I�[="���츫e��CV]ڧ�����%���u�_j�}�s� ;�.{�Ipl��2���8�st���\E��a�9�",Ȉ8-&C~���%�����5���q/|�y�}L;����>"��(�^@���W_<�u{�����2�S�)g�y��� ��]����[H�J9T�T�#٭�����#c�ٟ�Xn����|����|m[�$�
�[�$���-�n�AW^[.��5G�MĒe�K�h.�&y���p�)�f�Y�-Y[�:PP�J^����i��#k,.��:��O��E�8^�3,em���\�Oj�2�!����:��̬���b�B��&������z��e�Z�h�x�p��Z��[����v�"[�a�m�i��K�C5N�K�ÃQ^5���W��^>������|3/�2 ��B�t��n�cEPx��q�\�N�P�	��܁sp�n�]͑��r�� BQ!:�6]�a�7r��5v�C�Ō�s8s=�͊�)1d�h��5|4�ܓ\k=�z�;�ص�ѝr�E)TJ�T;:�$wm��31��r��N�Q�˪M�H��E��sǹ�*�MY�]�VNm�)J<��,ݮ�����{ԣRs�̝Tgv=1]7\�]*��:��j��Q笍`�J�K�qX�v�e:]]F��L�'��W��pǯU���[�/4��v.X�l੐G\�JJ
���6��I�w�R��kWc;f�a����9'��=��?v��=������ev�A�K�-=(b|�����};�c8�)�2m�w���!)ٶ�f5�N�pBiR9���J�V�h���ss��T�aP���e�bN=4�mb��Gi6����H��U�N/2����6�ڊN����UP�r.�Y�/'���U:�/Cz����]Ǩ����30u�A��v2v�즳u���!(�;Gp-�Y�o�EX�'�fqz�]�T��;R��>g#ٽ66�7�5�o;KT]m�֚.�b
e�;���hT�r�����O���1��_f����*��ڧ۹�Ȩ2Q1�jd�6�r6�Q�F&-��9S[O�&k��8�]qਝ��5ЅW�nb�|ݧ81J�e�u��:t��B�P���B��b�{չdk�2e;�3�]÷Lq�ɷ�j��y+k��'u1����n���_b��hI9M�(�\�2"7�����5|Y����^%T\�%�MȻ,�N����,'�GSUR��IA�3�6��x��Ӫ��h��CWе���̡��tu[�ZT���)9�al"^���p�Fa����^=�����[Ub�M���L�>�7�R���`���w�7鹘�4J��6M��\Iʥ,�_.�q�n1���v�{oиw�[�����יf�;��i��S]��v�����.t�x�Ntf���<���ܥ��Um�����N�W[�=]�9��|F�4�v�y[7����g��J��;�P��u�A��;n�+�����<�n��<��*E50�_t(K�ܢΌ-�2����O���@(��$H �8n뻮��)�J�]۲e���y{�S}o����nݻx��Ǐ^�^��I	"$��ہu�P(ˤ"����@�뢔�=q�v�۷nݽx���쌿:�H�"i�g�\��F-ݺ\�J!e#F!$`S�޽q۷nݻv�}�~o���@dID̙
�?��S�M�ӻ��{����N\Ĝ��	R�m�ׯ^�x�۷nݻz�q�f��i۱�.q�D �Ȧ\�
L�$PD�ID�H	&!s������뒂/wau�dF4�I.p���1&E�ĐRb���%��)D.D��b��Fdd拎�s���b � ���:A��W������II��4I�$1hB�F�4�B���t�
h�wt�"H'���w�y7������H����q�Ǭ���,N��x�ұ�iۤ2�u���-�]*��[��:rI�ϩ�c���N�\�{�up��֠d��d���V�ӻ���f�ܾ����R�]�mYg�/R���/1��s���@{�n��C�[�ץz/���=W]"lf�o	�7 �=$�xVlf;8��M=\in\�^f�����v19k��4tKS����~dw����T��>ԫ�ʂSl=h������@�rx/��{��aJ�u�7(!�ߝ���	�5s��b!0j������)��-�%�ôT��x.ԧO�ܪ�H�h�%�cc��u�� $$e�^�y�d\�\7�IżZ
��+�K$�X*�3+ThU����쿕R��X���'�x^1y�b!��q����Txh�Q��i1	�x������R)�4
4���mτ����{-��ݪ�1C6U7Td�t�.Cޱ�3�΀W�z,������}9!=�F�|1 &*��R�Ø��>�0�U�|5��6[^��~g���c�ǘZ�O�E����R�����@/ߢ��I���oU<Lƒ�Cd��7u�1-��&C�:�e�#�(okȇ!���~�� ����r���>�x>���=_�K�~�A��ٗ{�&�8�;Ӿ�.f7}3�WX�ə�TӸ4�ef���/-;�º7�{��4��g��sto�P�2��9�yoa(��a��C���D�)財2�K�����[�3h}���>> ��F٘${ݮ-�� $�_�`�F_��dA1�o�ܭ�����j�������fKlW���+Du��3:9����~��V������ �@DApXE���÷9j��*������>��X7���R)S����e��q���Ʊ�X�#��AGe~�>�#�r�Z����$0پt%������ ��9�3V����s�o
�"3�o,~�-F��Bۆ���|%{��μ4A`�A���x�r޹p�,�����.;�$�v�����-��j���E����� ���+W��"O�� 1��O�a'��9��<����5��%�a�	���������{Iۨ����:b��e���9���xJlL���nW�a��~e�����E+u({ۏ��y hd�VIE�i��5����A��mL���"�@B%�8T5�kS�cN��p��k�x��;����� y�|mЃy2��AF��_�R^9n�,�׬�3���D���%���}��  6��.��[͞��}#&t7c�l X�R%7�U��f�?S�܀���o���ks~�C�h�2-���ȗ-��[�^���C����/m�Zmt�g7H��[���X{t�Er	+r��i�ܔ+B�L���M����y�F���9��� ��4Ɩ���,�ͷL���X��۝aR���1��{�\�oW�{z��w*�g��+�����87�DW
L�iw�!W��Z2�n-U�� ���zg�XxG������TG� a���+�7��|2��,fJΚ}�nX��ʾ�;lz����X!���*S����9�p�C ��[�N�H� &E�&%��!���\9�����b���6��a]A��w�xa��6 �Y�
O��#=э�`!���jץV;��Cnי8�?A�1M���9ק�5z7�F�^�9j@�+�
0|��_���YǪ756݂�+/��)S�w�x����
�m�	��-F�s��Ɨ��N��������:l�Õ��*=�&��.�F�+����/%����rq[�U XU��c6���^�Z@���0iS�x��~��R�ܤ��^�C�5�����6��]H�Sj|)7Go6���2׿��)�s3R�[\�9a�]9����=�mw�* �y��,ᱼ���様&�)�c�X�_�V�בXr��"]���{�����~c��@���+ʆ���1��|����f)�Y� ��Sp��{��6���h� xn�N����(� I�ǜS;x�k˼ c�Ca{�<��TT[#yl}�|�b��=�*��ۋ)@�u�+�w&����d��Q�'�q���<�7@�P�Q��̇A�V[�qʷ���b��/�m�|����N��\�g�����t��Ы쉓CH\��ek{�]�ё�*�x�}�1�Iw^p��g~9^�Mj'Ѹ�';����$8�?qg�D��&�Y��Z��A�»]K��'�߾�b�E_/z�_�^x�T47= �B�0yN�
鋇�ygoF�j����K�r��vX$r��}�W>�T_�o�D0߳_
�Z~���b�&z��t�kf���\�9R��=r�y���.� [O�t&D8�t��%�d�?�xIkR�z�2o�CĬ��]^;*֒��v�����u5�^ |3�X��@3t��������,�_\�x�aex?�6nWk���d��� xg?k��������ϒ��rvf����R���@|����������E=�UA<�qVu�A��x��ϐ[�I�[���[��C0�Wx�a`.w�
K�y��-���ϧ����_uR1֦5�j��pܽ�#l�o;gtRt��(�2.��)�.�/��������}oۺ)�kzgc:q�:�#������ς5���O���B�����g���b��������q-yn��r��g�?xxf ��X��1�J~:T[!���k�dV�)�E�
���0T=�������f",�*������[zv�,��V*�i��B�d�X�?"��곖=��sr�4�*%i�&�U,읚7�a^��������Z��\���s��ٕ26,������si,B:_j�vUW9٦F��$y�{��u�^����Ʃ���� O���w����{�e!��j�{��>H��1惭~�L-��3�,����0��+\
C�vwr0��V�Y��Vw��/:�N���Sc/XF����A�9?�ߌh��<���+�
cv�TKauxr��`��w�dZl����O��Q��~�	S9D�#�+gM|�h3P�oE��6���������d��NFy���.��#y��n����f��]a���&��. W��/�O~+��������> zޝ�<<����)�	|`W�Cd�������C�@3�MC �30}\4�<a��3�r͵��&��k�^��u�<!���8Ƚ	z��7��{E�zڼ&�d�F���==:{X�ʻm�����ߏ�T�̴)�q!��`|�18
�=����G�R�B�y�Y��#�7� �=j�s7R ��E����{HY^����+�R@?XB�.��B.���x�^z���[�L�܇�=7mϚ]���o:!������cx�Et�xQ�t濽x��Ƃ�n���\�,.}����ɹ�Y�L�w�/ �����:�B
bY'���L�Vxػ
;j��gO4�[��Rp�)R�Dۉ��*��j61b����y�M�7r��\g\�FK�z�gk�}�f��p��s< �[��$�H��L�اH��T\��W;Zi@�u��O�̺��t6�Q53m=��ƺY�*H����mB��\�fp���@?��5M1�AB�wޟ9��_:�������؈��:oc�:���O��Q
ʑm��+�5��G�ȸu�w����tg/z&�/|�p��L�0��5����3�ԩ7�a�LU�υ*_3y��n�j8�������n~>%���8�-���9m��������Z����R�	�-?-�=�Q�o+���n�"s��O���,���&e����`k������s�w�A1�G��D�)�i��{��� ���9�0�p����%��&�b�^h|}�n؀�t�hL�N�&],쨐�:��A��X������Ky0�Z���b��A������Ƅ�揉�@`[���ֲg�}(�NV��.J tC;;���z8���+���(7��u�_9�o����Z����C��n�q5�(�����D���@C��z�n|�2�Rq�Ǧ��	:�q�������؉h}������gy���o�����;�|��Y*��,/h�����u+}�;W���e��XW� ��E���B���������9�F�_����W]B|H�G���κ�ݺc��7�?3*J�҃���Q�7�_Zr����X�4��Q��~�~��9_Lɍ��o�n��~j���B����%ٷi��ڪ��K|E�ӣ#f�et����ݶb�����l^�řu���\̰���dϏ�4�5M5�L��~gk��|=�}�g��o��(*)|�g��.�H��4˯{�]&bC=D?�lxw�9��_��g��I`�B��E*�P\����5��XB���B�ok/]E��!�pK$�(�3UĲ�l�珢��@�a�s���o2:rΨ���|=���A���ʹГ�X΄�qt�Z�_��\�C�p�~�A��?�
�m��%�{�%š�&!OG����������]�̱;I·�Zɪ,)�x��6�^X�`�ݬ쮢�*5����@c�3��o'0+&y�:llwM��:"S�*	UWUGE5Q���zj�\o<u����6D�v_WL>����%y����~�����ڑ#�U&R9�gE���S8���C���?{��[O�� �TE�B1���?C�9�[�e��D����n� 7:��I��)�u��~/JK��;=�g�p����	��E�mh�O��.�1gg�/`��ЍH�B�}����^ʂƼ�	��P�kHjg���!���8}����<{�Dc�B^u�(]>�IU�-tseN'"��kH�|����5
�	��v��Kj�fr�u�#��pZ���;��Jm4P�i0�3����v�a\���.���c��]�8"e�V��d{+����3��z`�!Se�ڛ}2�%:o���.�p��umv�O�)�׆�#}��I�|zԦ44Ѕ4�	"!79lQ�)x[~���o���� ������\Jn�.	=+^ʂ^����Ns==��8r9V��îX/k�c!�n�A�B����5>���ߒ$�wS����z��Ǧ��-�r|1-c�_R�k������~�{:?o1��W�:W�~ah_�)c]�D�򸉘'����C�fo䶺χ�L[3"S�P������c����<�������)�R�K���g/��^�y��j�f*�$^H�z�!��Â-��^� 3:�:��Ց�,t�S�AG�����lqz�aoMmM4��-���%�iff��C���M�S�0��g9?[�rS͵WF��l^����PK�;/��V���AR[�u��uH��~x����'\?4�#h�9{]�������0�f*(�x�����`$C��}L4[&��>�	MvHL���[�Ox��W������!꘡���e���ύ��`
��c�����cVK�lT��-�Kvd��^��#nD�H��e�P��l�9�|��Ei8���O�<���jr�s�W�0~����y�E�Z���,�4���VF[�[��:b��w�o���E�1b������3LcF9�5�7�o3Q����3p�ӌm�])e3�3k��n�e��4�{����o	�;n��� ���{[���jWp��	7�L/�|�������iR�i�hA��5���\T/e�񊊦i��:��z��s��,S��~�c>���o%�=��z�4�`d{P�v7wr�ꮙ���v��C����ü`Y76���]7�)���+�e�b�F:ܵ;����1��ޜY�T�Ű\2=w�.�����C���'q=�z\���~b���)N��JT���Ϳ-M�	x{�s/R��?�y��ƘB ֘ຩ�m���=��⺍�a����k�mBxUm��l��\]���ʒ�AW��t#��ڹ�o��Pڻl���,�튯���)P���|��s�T�R�522�Ű���`Γ H���v�֝�f�s6Ӆ�H���m1�4�܄^�y�y�j|�L�q���Ku����G��Y��M_�~���F�f�St�c�l����K�~��`�!��%�^gxט�Ͷ5���q��4^�w��9Gp�-K�0�}( '�!��e�!��LNM�z,;�#�{ta�a���t�OC�@2I�i�7��j'7��1��y�S�c\�}�n� �~��=������t���dzjvD�d��#r��Ϫ��>�7�;��[��>w4�)�kt��DTg�����������ڭ���N]��1=�9�%�c�ftcs�}�i(ʪ�{dQ��y1<`�v8h�q�sh�N��l3Q�sa�l�`�/���Õ���{��{M ��@��I 4� ��a�{�ژ�S�e��|�r��y�g*�a�cO������^\���v~���}���1�C����g5O =���ۄx��{XL۟��_D~c�4�-��{E(����׷-�3u�r�a`���ս1dD�+�h=�B�Z��=��H��a�+"��OM��Sjb�^�r��y�d6g[]�N4�2N�S@2�_�/���3�Gk���=On����7�Z:C>V�0����k�pa����MGc˘LK��.�"�QF�[X��^c�֛����B�A�8�P�s��S0P�G)o3�2��VG;��R��c��t9�Rh��2�K�T��!�Q@y��b!��Xs!j4� �~{aC�>����ڏ��A~V.������ٲZ�?T�����ǝ���k��3o���ϼ��"r��!�D���~�D9��/~���\�ܿ@��U�f�m"�/m����D�u!7C�=���>$��Lb��c_r�|{�!�/�
h*�	��܆��X�U�w��:�F
y^���9���5��c0i>�o���q����C>����a��Ŝ�c���i�p�7��6䩵��Z�VN�Zd'�+#&�vj�7������i��.���޳�v��-9M��.��:�mV�PSO����i@\���\����QH"1F�Z�mq�h�7�.�U���GCќr;�Սp��'H�7U+sU��E��6�]�����킔�]N�+i�tU��AЌp��dP�J�Nf��3��g�v�V Ük-�5���]ux����fIaέ�!�+���5"�֩�ݭ�[y���?]����-�?�7yz��2��W5 �*�V�)�+���OZ�Aa�}��f],\�%�{*��z�ck[��v��+��h��i�Y��v� �DN��q���ܮS�d�#UEf�ת��R��3=�3b��H*�<ֹ�������	h���'"�xŤ����͓T��im��.��x�;�16�CRBu��5��c�oe'�[�4\����Sc��*�r��Zź�Z+���F!��Y��s�V1�iT.2љ�:��f��;-��\oN;
�J��N�J�K�Zq�I�)=л� �ZZ[WO�˙z��6�S�
�r��aOw'3݅^�c3Y�*Õc1V(�eV\�33k0#�B��l�����Ѽ{���\`��2��=�]�bp�T�;�n�[�Ԗ����3F8(�%��z�G�,�E3�5��7/�9���n�
W���7_D��;|7
��v�l�hul)�����@�ĭ���|�z��Gc�,Um>0H1�9��c5z`z�du��(,8�>�	�ٻ%,�s-)�\K)c)�*P�Υ��L����d�{5��$��T��nı���B�3��n�)N�c���]�E�)��7m�p���N��D�e^鰃�V(�SCE�8k7]^�͗�v�3!�O��v97@�!y+N��г�?g��T��=j���!\�ս3J���u����8jm�ɪ�W��R���1u&Ҥo�#����ǹ�����O=.j����'XG���\�K7m`��I#��ٻ�B�ɒ3Ya}���r�YE�Xg���H%m�S ��+�xE�o�V�&ᨲ1��mܹ�۸m��&�:�i=;�b��C4�-K�d �]�	�T'm#���$��n��i9��"��{5���ѩ��=�,��d���i9��ܴ�ˣ�]6T��+p��9��BB���
$8`�6�̝�u7CdtǢ�{ICF��y7xܳ��ݍ�%I���M'�C%���f9:��@��2�SǢȻ5��_`Cf��D�]�D�ȉ�<��|����K��`C� �W4L��QB�M3�w��yt�I�뫒Y��f52Lh��w;�1~B�3R�	;}x��׏<v����{��u���O�"��؏u���i��\�R� B1��i�q�׏<x�㷯G"HI	#�*2�*$L�h��l�5�W#c��J��b$�N8�=x��Ǐ<z�q�!�'�u��U��ݒ4�7C��(K����T���d$d�8�8��Ǐ<x��׬bdBD���!	"�b1�d� [��2,� Tw� ��(ɲd�vAE��U��*SB�ԝ�F��d%;6"CH$�@��q��ѷ�_�Wih��I �`Ţ�2�If(�o6蟥��{����ܼ�("	(�"��$
d̎�F*M��3$��CC$M"HFf1cE�#;�D�۬%�;��|�>|�((�I�Yi�aa�/Ĕ`i!E"�%�Y�"d� ��M6|��B����Np���7�K����Gc�i���鮮�EIpsOA���уQ�����gN)5��9C%��'o*h$i��6��F6��h��! JqƉl�b���ٞ���\� v�Q2)� �DH�˂�i��!�D<C`�)P(�D�$ �(@�R?���y4��$�SM %4РSM�B��H(H���>e�^����Q��Y��!#��6I���Ζ%�l<��X�W:��>�1F���*i��#}S%*�~���y��x�"Z������l�GT˗AwfA�L��[;_��>�]����zY8�Ǧ�U�$vس~�l�W/��MZ캵u>�����&W�qG�0&���x|~���|޳#���aMM"�)f�s�z���+Z!�_�T5Y]=�D��e����1�/-i��z�w�{�l�}�ohT�;cFkŗ\� Ș� ��'�sͼ!���A텇��E�?Ji����l&�O�\Sm�'u�!����FCH��S���l��z�'�K�t=c�QA�]D>��~p{'����c�\�B�)���Cr(ֳ��qP�^�ݖ%"��k5��l��d0t>��&����+��1lmk�>�/��n�cx��+U��]��~�����`QkL�������J�i�_?���`}�Z?��o�ͤ�_d5��+x)��:�/��� ��R��3�Zõ�W��oG�=�d�;�j5�SS�=k���$�[Nus˻��A��8�v� ��<i�㬣w" [%u;o���~��f�����j5^����[�H��8���{��%�Exȶe��T�ʝ�f���N0����O=ל�+[���H���
i�@��U
i�	d �{�2�w��]��\���d�y��W�<��� a�����i�I���^r;��2a�b�8��nb�a�ijJ{F)�x��h�x���{m�a uRL�߂���߹�w�G���!�-3����u��\�+�m��_:	Ac^\jJxw���Ȯ�oF����o��P�	��9�zNz��Դ��N1+��Z��3`+�a ���_u�-g�/U0{�B�1��D�`˃�`�t�sM�����'�k�PK�6�R#��r��W^��:ϡ��=��N@����5�x�;�2�ަ�8MC%*,�:j'�!�j7bd;�>�n"�J�4��I^�
�d38�<p�a}3�����D��ۛ�|^�932�����vm�<`�6:3��p%�ↇ��j�HU���o-��
�S)�fo6U�4Nd��H�!�1�[W�۞�ǖ��CCN<ʨ�K�c������29>��=5[�V輶�	=%����4���M� »B�͘�`?5��ٚ������>�.�e]�����B�����YK+��k��2?vc��aԦ����sm�8l�H�� ǖ��lT88hU�.F�-��j�9��H��S���U/-sHtXx�D�����=�6um��e��@~�4���@�M4�2M4"�B(H�� W}����*-l/�/�<��~aA��D]�?L	lZ�[^ǣ���{�{6�%�ש��GM7v��p�b�T ���ν��
"+�'���%����)�x�ͫX�~����?�~_����ϱ�98��T�3
3ó�&ǐ��c�X����+�rBh���ԋ891���� LJuc��	�JT.�&���{gO"���0���\b���`lລq�q���2ͩ�tGo�b� #=^R�lli0���S0li���7"���_Z�ݜ�T5Q��m�HW�]��K��!ʥ\�,�l�&:ܳV�{��L|F�v��ρ��������
��qu�^���L�Uf��v�}$���⠱����эM5c�os5�Ŏ�8������b�����Fz$��LSl�F��Ra�+c���`�Ʌݮ���.�@�?*I� ��-#�{�~ ��:��� �\;�+%�U<&���۲ҳF�)aVc�׊�^��83/F���G@!���v�M��t�1h���\#�߲۾��.�b{c�6�0�*�t�]q�Tg d"�Z�6roˣj��7Z��������r[��������i!��S&r�6ȗ�bn�3Ĭ|��v��ʉ��UQN�m���M�0�գ^�$��nU|j�M"�4ЊSM�kv��Պ�cj*��X�ތ�ۜ&��%�*&��R+[�S��{��d�s�#nk�T�h���+.��Lk�;L
僔x�Y�v��k�Y;�y�?)�Xܠ7�ۡ3��Xh�9'����݄�C'~��sQ��HQ����Cs}N$D������2T2Cd��7`��Š�bj:v��&#R��ퟕ��D�Y��
c��%��z�!�$�/V�r=5="o �5ʮ^r��6Ѽ�
�ǧ�	���r����N�>�A@�����Ϟ��#�)�W<���n��!���(��v��f��w��h2)�i�X�����NiKbF�n[��6����>�S�6|��Oy>r���dIzt�
=�Bޭ�[ߝ� �����C�����788�[�C�;����y������_���L��Q,�T�U(�|j���ⓄȪp���3}ڝ�c�;���/O0�^��"��ߪ��b']��L��*ƶ��7I\�U*nt��7/����ti��L?U~�`�c���T��1	��W�a����-����g6� ׻��{��܄��kylш�>��s:������3pL���a=n�R-PW�[���.��+!? H�D�j�z��17�X+h�בm�"�4�Z&]�Zu{me�c��c��d֊�m�J|�I'8���|>�G��F@@��	
i��ݻv�F�F�jm���@�d�����V���k�O/9�'�]�9Ի�ͬf�i��j�/%��e%�6�J�f�%�#�!|;~�X&���6^��y�b� ���"l?�p��;5�g9�}r�Z�&�d[e�L�~��dJ!~�C���6�}�B.n��Q�>�C��_h�c�`�n�H�<�/dH6yB̄��;�6;�/�=����7̹�*��h
���B}���Z�dI~����Mv;���8��R�O��&FW�-�@�`םfж	B�woW���w�aa��vO��<����=��C��>{Q�3��v�.�R1 �{����G�lQ/��
.��e왽��S�dC�|>.Z���E�]�����I�[�l�X����ut2W�8�.O$��?�����a!�ߕ_�+��=�@��V�c�	�����h[�L�n����9Ky�ۓx���݋/���\�j��XiW�X�F.)��.Q�sR�>� �������~`8������T&���=���J&a��c[�y���V�f|�B-�����6�%6?DU�9{��)mǊD���\����&�Hj7�L��[:y��u�����4�dk���\�T�#�x��]i�1I�L��ƣr�+۠���\q���e0�Tm�N̽�/_Un��m�/�@$�$:� �l}�Ǳ�������=�jcYq塛��(��A'�|�F2�AkpX�:�\�֮<vŤrmo9��M��^�9�{��P~�hU)��R�i@i��F@E�@	 \��I�
��pk��Cݸ\?�m\�@�t ��@�%�}:�UcY�O�mXj޼�܅Ӑ�s��#�\؉N����&�Ʊ93��>v�ciH�)�gi+i�ǭ+�a�p�ve�5���k��Tl�����<��ƾՖ��U���^��{���I�.����T]��j�x�d�Jqo�L3�-�WN7�C�Bt����X���r��[��ֿ��z=�����ǂd��E'��m����}w�xa n@�:1�C��s�)�3�;������ö*&��r�'�O�� ps�L��ӳ\������
g��h
\F.��F�C��RL����E`�*�\W���
�Τ«��yj���R/�౥ơ���q��V�Nn���j���69l�5�=K�x�Q��tї`�E���c$+�`��hQ����ʮ������u����P �pZv��?��遌�Y�J���@�zW>�6;���]��:��z5����W�=���5��i�3 �c�&I^i�ֈv3򳙗����'����et��	���ǹ���0���P�ɴ֎!{���,W"%4��ێ��/�#�n3�:��t��7�l�&[�����I��
+��e�`�����6�f�7m1�&ɽ����J��+W{X9�/�x��� �@A$D�4��J҄}��a�-Ž�Н\��p�hg�m�u\=�`NPhsI�t��%�3���@h04�	L1�7�tmc��z��Q:��>&i/�ͪ���yྒྷݏ^`o�[ ��yw� c|��l�ϽG��lړD��>ؾjb�B����	
��	sِ~�H�!��0�k�%��:�O�{��}Y������`t.�!b�w&-U�5[�U���� ��B5�T�I��V�1̕�m�\��/�/�!Izo�=jj�W���?�}����b �T���������m��v����\�ԯ_������6Yxa�������%�L��
L8�OE��(�p�=�O���ww5�.w</w�1H�L�݊�'���y�ֱ8�Tm�Q��z���Y�*��r�sDJ�U�������e}�&\I��%:�Ҙ&��*k	�c>�� ��OwdP�9�/F}+��[���ް�����>Y��`y�	g�3fQs��b���ģ)� ��)ﲥ;�#�4[0��]Fm�M����1�gbZ�o2����.����eX#�i�����8�ڼ0O��{Jg�K��Tk�����p�:��%hN�^_0�rV�ǉ�J-mj�w�m�M�=�<�PܹGi�S��}�� #�_%?�sY}���,�,���Yq���dvwd�$�w|��د��pr�n���J9r͗هV���n���ТS��*SM*�4�*SM("TP�L����;ٕ�>j=��p���zhC��C��6Ⱦ�&��;���ភ%�TsF�}�w��/�k�ؐ�3���%ܵ����=�3��֡#Y�˫��0֟^�B�6�C{J�F3Gm?f��z���w=ydi��E�k	����Џ��-�?sM3����'��"�,EP�\8�b����.�)���Хǽ�#w�l���C���}ߩ�j\��7p�m�C�b��������N� 
n�F�M����Lz1ξ���c���XE!5m��OQy��3��߰/��hw��B��-Y�@6�d%��tz_�>�h�3UoW�ݢ%���kTAŴ�;v;9\������lgwD>0�yïKE���K�Cd_U��Kww�ۙ`w6��γ%L�.Ŕou�0w�T2�B��2 ��>V6i���,\q�k��ʽZ�אyz��#'y-��#׽�ɢ�ً![r=4^E��y�fP�a�rG��J�_�?>T�����1\'����Z�]]��C�m�j(��O�ъ���J�B�~?xˆ����\0�Y B������o�1{�b'}PvFǲ�	s)<���4�j˨#�rbfN�,��{�d�:˾���*��z����oF���%+�wR�r�&�_6��|��tP>�}(e�������Y�E�NMur����3tr5>���BM4���@M4"AE	�D��5��y��C�ݩ��wt{z�j;��*�6����GsM;�Z�}��
���"S]�2�&�Y0^��N��X&7^���1홯o-�xa�$�'��!���T@�s�ju�lA��d��SL�ʷ����j;[&�-�^��VnQ����~kw�n?8�����4H�8�Bb^�E�h�*���g@{�3V�\q�ōL��r'�.����Tg�C*}a�{=���j��s�݇�bw�_ՙ��z?F��/���J�5�9��W�ň�>�b�@AG�Ȅ�Bc�l��A{���c�ڌ��M�&�}p2��2ɂ�/Dŧ�O;��QhٳL'ú�{��p�ۡ�.3ʸq��6��Jv6̞
��&���hWd.�CQ�HM��\w:lwþ5�����?u�C��gJ!�F�s��v�ȝsS�1�\�c�Jq@Z�'�ʨ�x�H��)�P�N7-|Mw���_����>~L={T;V��}l�V}p�D�u�\�ό��F~��Oķ�-�Zc\2b����t����Ի'ɳ#'ײ���1�;��b�e��)�[�<�V��k�C�j���:~θ{|i��$M�%1��6sϽ~��bU���mӫ��dQȂ$=8.e-�it��9_c*��
o0�N�R���m�Z��D�Q�~�V��՜"us�����d�z����U���O��x��T**���j(1���e ��H����3{���)n�f���!�����9����$�V�.(��)}k�F>?}C&�}y6`�An�4w���Az� ���!�]���uʼ5Y]�4���8-��&
>��/�á�D���Rnx#67����<B9���@ǯk$M��Qz	@A�"f�{^��yǌ�׀��%���i/qo�|��
��>ķ�7��E4u���~Y+��2o&�W����mO�8U�W=��?t�G偩��]��H�\ۊk��I�gB	��l������Y�_�Q��o�r�&��K���z^�`�?�fXs�������>T-au�����c«f��Oz��{�ơ��%��&��E��=��Xo�B�#+i��z�:lgv��m��L�QҜ����\َ����$�*S%8���ȶ7"�F7�56�8�r�(��g
�Mۓ߇�d��"{�U�,.ހ�+��-ފ&�>�sӽ���1�(f;�ޓ�;/�K��9�V���*�y����[�!��(�1L���J��6��sם�k�}�x ��2�G���&i�(3/꾇ptGu������[؃�����%4���1��)C���H�ΒNħՕ�v��-z2��0��`��+�K����̜��˃"�u�U��F�J7U�eN���TL�X5ۤ�u��;V:��%�v�J�Fq̑�-�
W�����������R�P6N�s�n�u��ᦔI���Ƣe��u���F�wc�Z�i<:�-L�|~�]�E�=e��֮�k/:|��y�=����L�.$�*��.�q�*
�-v���lJwC��k���9��v�e=��MR��:<J[�-�����7Yx��Am%���s����D�J��,R�I(�x�;Oz�7��ҕ)�j�5��a�1{�=��T�V��d��C���{�+��[_)S323g�ŋ9�]�c�v���>'�tovCno#�jlA��f�d�Q��]cŗJ�WSN=Ĥn͑s�����0[�Z�;Z��UXtU�=�k��b�1��T�㛁ɰ���JS�)зP[�ޛ\��yqL�VnУ	�Ǧ��&'�<�Ŋ@�)e��ӿCL�.lk�\����sk^��Ġ���ï�w��N�34s;(�q]:`?5J��L��E�D����a)��;�+&l�+�������ѱ�nT�{�/7�(��2��ۊG}��nr��N$��$čD!�k$Y��/ToiU��/C�$�`�wFE�D�<S"EQAN�D#�[�R�@��f��J��^�l8���f��wSd��$��%��K�3]4�d�nְ]V�a8VV��h���DJ�dT��wU��N����Լ��y��3B�����V�%��tV�<�L�l�|q$r<������Q{�W�{Q��^tB�3*�����wM�gr�P\�37]r�sv!�~��%������ޓz����3�[]�ur�q��jmg��K���+����3DQ��e��e���53J�U�a �n�B)�A��sVHvN��r��s7j�Q��{Y[�Q�K/d���BI�Q+�#"��˾n@�7բV̵{&��4�s��i�,�k�6�p�|��9�O䵒�гd�����|�2-e�e�CQ�����$2բ�K8u�*���uEI_%o�#�dI�37����A.��u�w���'��p��w�R&+��*��/��K:'Rpd�	�������N�=J�
e���xʗ�C�}��K�pv.�9]��[�';\�	j�f��%��Wn��Ĺ>�"�5ݥ)�u�hz���-Tťa���Hbwn��O:�׵Ⱦ]F[Pa[+3e���Ƀ��57U[%��� �!�������lYլP���(��b����&͖4P_����t�`�i4&�>��I"�B,���i��n=x�Ǐ<x��ׯCHd)���DY$�Ys|��T���u�	�wlF!�|���}�x��Ǐ<x���2HI	$ H�"3
@э&I"�D�]7���BI4ӧq�=x��Ǐ=z�1&�W59��td���Kv�#r�B�st�#	!lt��8��׏<x����7��t�Qˆ�sq�Ζ	�L�o��4d�DD^��*P��`ѿY�^\�!���[�B����sf"W�Dٔ��wk��cwuwmWC4����wWa��;��{����)��˕=�/*��戌A��M�k��cF"���۠�ؐ�A�{�\�L����툈#˓��zL��Ё%FI�p�wRK�۞��fi�p���3��݂���w~�MHcD#��}}��_�*�y|U�����kM)[�'�Ia<�v�odtZ�'A:*��ϠަE�ǡ�-�:��j��Z? 
o <���< SM#DREH�J-4�FEP$�Td�޳���{�~s�̪����kG��c�B_���D��M�T;$��-^�r����C
�k�u��ڛz��ΧW;�or�����l���y�^K��mB&�x�� �E���c&p�h])�>�fp;�g�F�?���؁�f�)^���Ŀ�44����P�@.�.)S����c�م�������(�s��|���"<��69��yɆe����<)M�Z#�;���Ϝs,�4�]5����н��9� Li/A��H.��`<�j�ظ���j�8��}SĽ�5ΩL8oD��a����â%�z�H�r��.�4�1����5�_!o�C��� KkЇ�{aB*-���`�qM3$w=x�4�fN��9��7�uL�YGguM�׆��fh�(E�	=z^��[�E\yj�K�{��/QR�0qz�]j��s-������R�Cc���S�H�����57&�ߥ�eG��-R-��M��x���:��j@^�g��3[~��l.a�tS<!涰������./�[ؙ��Ӛ%߿	C����L��6���=%���o]c�M~��z���r	��i>$�r�[OEX�G�(�k��5�W5J�3��:��o��@�)~;8Ƽ�ⵦ�U�p��{���oj4�U_d{�b}%�+�c	!_�|�+���kT��Z�T֖ٻv����5RA	B@@r���5�眽���:�}�
N�俘�տcռ4�S�l�{d��ruR$Qw1Oh�Cz��Wxε�&ڻ�K�J`����]�M�׶=�xOT��wW�M�/>�ݜM'�[
=�O�Ƈ~Y��>���̢�<,Sި�%L:�f��z5EL��{��������r�Ÿ�}al���Wo�,���}�Sz(�a|�Qu���$U��3���6N�f�t+^���6g��������g����_?W���g��wޘ����͕��m�̈́�V�N���c�m���cP����Չ�a�	_DwK�/���U�p��x1�<�yC�)Cе�(��3W���-B^��:�8K0�� �ֿ`�x�n�ʾ7���Z��dK� �0�P��%���(��X��;���W�dI���b��'|#��t!�=�Z��f�� 
u�"yX�cϖL�q�Od�=4�DUԍN;����~�V_1;�b����~#	��#�9g�?,���G$^͗��?O���_�nXޠ�j8���sP�%S3v�,�ϬTa��.�^��)�UGog���ܛ�(p�re��Tr��X�,>�Oq�%����Z��"�l�]��XNG��غ�9����������(�������"]!�z�CZ9uܥӥ���H���O��?���RA$�2��H4��F4҈�	 ����l��;�y|�����kL͝v��W��������$Q��j��X��.T/6�v)�?�M�;Aݾ/�~a��DJ�/b_*��}V�F���OJDN4.�\{�!�?Fs��Z��ݵ����/�|c_2O�X�T�}�n�G��F�y	��Еy:�}��z:h�e�m�c�<�-$(�����=�=Ѵ';�O��[�@<U�A�QL9��Hu�6��^����v��amV��z-�n�F��7W"�4�4C�wx`��GG��0Ţ�ι	L���H2jY]�a��f=z���'��e�n�Ti�u7��2�����as
y��o1�ju��l/J	ńbZ��)M2R�Mr�k��\�i9Y������:/�����툑A@��f�N6P-v=�٤K#�n�?�o��S������Q���|�<d�uc����Խ�W5���/��}5�~^c�c�}��Mp?R�
��G�#͸��U�����˵�؎d���)QU�9�Ǻl��G�Ű���4̈́�\�.���3��1�����̬�<܇C/��|r�%�=�NV��ni�.iv%�w@~��&ְ̆:��-��~J���A-���
�7wJ���qA\���Hy=����پ/��ֻ��g�*u~S��i}_�'��!�����mh��N�i�����>h�cQ�
� ��ި�&G*�=��	�Q��k��.46�+yq����r,~�U)��i�B�hjH!"�@ 2"2
����~\()�ʆ8�y�NķU�T;$�͘	�:O��'�q/�����oPw�)m�	��P�5Ө�Bm�dN���-��<��~�^P#'^U@�x�H���Z�.����H�Fw;��u�z��pla(9/"���%�������K,��o��O�5nY������G��~��s�\г�.<�������4?r{<�#��>�$�-,�����Lc��?_�c��Du���C�9j�;�׆x�������C��P��lr�+R�xrL���r�	���;k����^�y�A`|e�����S�����s��xrΈ�6�r&fCD� 2�C�-u���[���	@A�cš����|��>O�����T���l����G/��c�{��aM-5����W6�d4�M2"i���2�q��#Y�Ő.� q`�,?'u��za�}���n/��:�(�@�;�k6ҟ�Ư3��K�v��}��Bz�1����а�� �O�+?�X_����G��zH��>�\�$��b(N9N�ݽ�z+���E���z��8���ۃ"��sXj�9�s�!��S���k1u���d��f�z;Y�}��^&D�XU&�5A&/բ�p++����<+�O6_�~Oy�	�+P?V�hD���2*F�UZ���fʯWbu�flC2潭�	��Q`��x_Sr՘T���w�����{a³w�+y�@[b����ZTG6��M'X�T�p�Jqo�L0>�ɶ��m�M��q���"_O-��.�j$g."��!�����H�oJ��u��_<�/Eq��W�b�=v��K��OB�7oܛV6�����=^*o�8��vS���'�b�\�pK�ӱ<��d9{�'P�|�'ِ�t���i���R�*���=b���lv_��e�KEz1�;[<c��Ⱦt.��8�rz�� ��&�{dr&�C|x���yT�EV�l�N-%�]�T����"7�an:ƩC.�k`5���q�pC�h���80��	���'��X�:z����Ywx�G���]�����K���=��y�zhO�]S��N�����3?���@|O�x�A�<m`m-/���Z�Aa�Gz|5n��%�^�49��{�@���F5�E���v���m} �l�bs{@K3�mٮ=[ԘV�Iz&�����%�tg/�X���Gq�������qV���ӿ֩�2*�ܙ��S��o�p%����}�6�Z���duL�������M�����sl�<a{bf֕e%���WC�_k�wΌ?�s�UOe���ʵw��r]o�2:y�Slr;W�~�9��e��@��F�hR�iV����,�"����������/}�`>�?�п|�}�t���d�Jk䈒}
�������x�/
s�PC��K/vܙ�r��踚xn��p��ğ��\/� Uj�Z��[\�KV��d;ph�i�R�1�j�xfhC)W�E�S��z���,��g�t�tb;� 3���G���-��~K��ݴ����jLY�cC*Y�:���Y�m~j{�K����,��q�g=�;�`�S=�vk���۶�˸�Mg�<ɑw�bө��������b�ᩭ����O9I���Ͳ���F4��vG\3�pk/�� �֠;�S�J`������2o��?ql���L���"��l<*�37��"]��B�W�e����=>͈E�y�X��QW�6Q�Ll~�,D��&��3̎8Ow0����tw,1����S��J���^�5	���"�ZeݫbF�F�a�^"�|d�nMk`�M����p����O���*{��h1K�_-ry���r�t�����9cCT�~`)8����d4_�t���KO�h�gg.���z��\��X��j;����WtX;X�abc�:W�Cg�[Vd�]�ѿY�ܝK��܌l�;>Σ��L8~�æ�x~>�#�Dy�O\��를��9��mL�Ԭ����hͥy�V ��S���u��ˀ�#B]������C�|���O�*V?f�B+"1���)i�i����)"2߯k�*jM]���g��L������r�:8��\�P����92��D�Z��ȍ?���v���*5�QQ��aTCs9zw�v@xV��4��?�H<�ODc�Ƽl}Q��M�BbX�o������7�v���l)PK�=ҁ ���ض�6�.y��ȮO<��PXȇd����ou~3ln)P�n�O��gӏ@q�i���G&0�:3RPæ�ֆv��g�`�Cϐ�o"[��O[۬�~Z�~�����������;}��H֌g����4�aݠbi>����o՟����8�wϨe(w˼��U��ؼ�a�v��u�H$�4��q�Ց,��d-��t�<Sս�=�7e�{:̆����vwwC<�Q�%��G�E���q>��*��-2U�Ŝ��g`�W߅$�q��[>���kߩ��|�#�D#��W� Xw�t ʖM�,Q���i�{gS�)�n�U��^��|EĄ�ke��b��^�.�vff�A�"Sr�A�RȚ�K��Q0��>�J\FD��mQ�Ù[Նy�.����v]�� ,�������#q@��)D��z\��4�my�|M�V̯?ˮ׵��K'��lv�x3#�[�y��3ϻ:_^�\�C�LNY�}�- �'����RK��U��r�INl�zJ]���R�vK�N>�)4[30�uZˑ�	�b��/�ȭWwlW�^v���뮧4�+�A�Ѕ4д�%4�V`�t���j1v``��
������|w�##�x..��a�4O�{"�Bb����T���.E#�}���T�BX����c`�|�q�ltzqmP�����j5���F�*]���B��kc<ti�ͨU���Cy9W��E*W0�LYz�<�=�l#�(�C�}uP熄�7W��:��y���ܻn:e/��;�^OK�Z�J�wgu9�i��r����Sζb�ԝ�����G.d!�w�
��4������vB�E�����J;]R�חzy*������g�P�䓇2��y��#������T��_A��!�n�5�BO�Kcy�y\�����^�߫`��3�}7u�����RO���v�?����!$���.9����n�{؞�~���l�6�n�^،�i��ya��f������5��*�O_�c���mM�!v��؎���mŋȖ�P�}��}y�|׏�	�EV��q"<�4��$�1��MN��"X�!,ql�ʧ�����@_��H��"(v
|��+�����w����k���E�\���"��g]vɕ�/V�~��-{Ɩ�O�*�B��;��G/]GJYKb�oh�lֈ���ς��Tڃ�ᛧi�sY�e��R���gS�k0M�aUL��{��.+zI�%���{�ѓEo^s3�?L�H�@�M)PH�J�*Io�~w���|�ᬞB��7�1�ݥ�:܏?��M{vQt� ��Dy���ҟ[�9'�"�[�#n�7j��G�̴\	���$��� cW=���<��hW����%�CW�2x9j���Z�H��ɾ��i��cn)���a8�a�wk�� ��z��I����lKx��j����<���P�[�OJ��}�� ^��_��~!ua�S����A��ܯ�Yߔ������.��}�ى�f���c*��RS%��mK<:�5)YO��?��.�|�Ur��luŖO��9`�9���azS?=��_�T�)�o�&�Mk�iV:t�H{j0MW���ڬ:�p���\����&��<�X�j.W���t��.h9"j��+~��ԂdsH�� y��`!ol��K��ʞO~&)��[�������i��[���U7&/����:��7�o��C�h�2�	r�6dOU�&�5�A��f�nL����E��_Zy���7ןY��?S"{�K��ǯ]y!0]�D'�^�m��	yOp���)��P9f��唣&vG�³cZ�fb�i�a�-�M�����E�ݷ9,��:t4�.A��q��Y�tW������O9����/����4g*cX�Bj���xE�dx,�kac�+�T��ә:-�4)�	b��뎫k����򏳸1�4%4��V4�54�PHA�o���ٞ��9�7��>���=(�~�t��J�
��a�����80��`c,�n~��,�k;iE���B�Tf8^�z��M�6��ң��lƜ�it�@p�@���P����~e���>�l����`Y�^_&�h��*ad�hu��Mc�&5�lq�ZFt�^�9���U�~0�U|�=��CD[W�E]y��D��q{��ʼ��D�'�=��@ȊcST󏲮�x��W6�g���u� �k�^���TT[#c��������`�V��؇�������=5���p̸(����DdB؏I�^=��|hq���3��2
e��Y-��g5��g�-�^��(k�o��vz�E���q>��M�fU�YwZ�}��[��_7G��Uȶ��� ��y��{S)� t�y���T?
���y��z�@�+4�]\v�t3]S�ެ�?�P��g�&T�P��NH��x�^zw��Ol�ʅ>�C�����m|JD+d�K���>��J1��O5wB�3�oaN)7�h����2/6{������4�&&��G�� �.f�U����L8%ol�p�!�Jfc�5����x\��ǉ\#I�^�4E6�uj���L�#ޙ27�4�Q՞ۥÜΎ�m݉��wY��֪r�2R:�%��U��_
��+�j3���\^���񇵕p���-d�_9�*���T��'�lÖeq�ΌN�]W�7xm4p��è�n{�9{2r���ݾ
�u2��ø��H�w�2c���P8�H�f�%�U�j�0D����,�!|s,A"�ʆ����L��-eq;��(��As�Q�s^\����U9+�)ӻ���-ܖF�l�׽nRdm8D�HE,��7<��v.��ӰbЅ�/t���VU0��Mq�뺩Kǖ�0��J�w{%���X�k���9�,�� ø{���mm���<�T �FF��p�v���ʾJ�]b�x�b�B�{�)�=6�
y3�,җ#�͜C��69�*U�z�_sg3��)�����E���2�2�b�W*��Y�0"=]<�&dg-I�tN���L0r���Y/���ٕ�v���Aڕ��ڤ�o��9��{J�%�|�z���f�D;����N���ͫ��
�y�#aN��Z�.ܜ���Cd��"�a#��3�K5[��霺����0�g��\*�b7!F]��sf��.�a���SԹ�i��sg�hKϝ߇t�Ϥ�j�6QZ��*�;45�>�q�q���D�s�V��G%�:���`����H���փ���nro�̓5��E�k�n��T�:�=�y���X:�5���:iQ�0k-7��\��.����!����	`���`�wr����-���ܔ�Z�Wkd�'xۜ����UU��M�5��/8�&�ي.Υ��z!�v�f�ա��x�vG��\��$&�J�fK�n����>v�a&6ș��oo���k۩�%�Ƹ��1��k[]��>L��(�ol�p�YFѱ2�bd^֖0+���m���f	D�Ǹ�4���[+5��{
����T�Y��{K��N0Uo%��V�$F��6�[Sk.��}��&�N���Sӹ�U���(w
��Ք[��5h���㽣�\BVeՔ�Z�b�g�z�˒�2:�ON�Q:��T�����6�n'O$�hvv^�����:Vz��U�H�Q_���(H�u(�)�%ԍ%�g>��&����M�븽���E��w�΢{��ٲ(h��3[�ʗ0�-^��W<��tp�\z�-�*[P-l��ʾ���d����v�.�H�4-�^az4���TU[�Xy�[�rS�S�˫�����v愻�l)�����4�n;3P�B�%q��l3E���\(E1oc��nqEV�k�'̃4I���3��M]����I%��8i,("P��@�2���m�o��8�����Ǐ=z�;$��HBBC#P���Yn�҄�(�BFLFH����|�ݒ�p>8a]ܣC{{}������n=x��Ǐ�z$��"BHB!o��k��}rL`�؂�n�@�.mҌW.�[����Ǐ=x��Ǐ�z'L��B,�u�	+��C:h	MC����B&���GN�q�x��׏<x�����2\���p��v��$r7RS2b)���1���[��#G|�1b�A�c~�$�r���[�*��ɻ�}:�e|nRo�̘�X��#TEIlh�(���ܠ��]q��C^h�\��󮴖�uSW$�E��E��\,��D��[���E&j#�ܾz���|�=��(D�A�N/2�pBCQ@LB8�26Kf	
!4����܁&a�B�,�eX�ѻz���X�]�Hm*��5���V��CkgV+M��ʪ��Οu�Tyii<���`�m�U��A�'��$BQ(E �ȊhH�����d	�"�A$|L�-�"!�#��m��F�)EM#fD�eE	Q(S�`�@�Q�"I�SM����Z���C����� 1��TI�H��J��@�EI�邏�|��}��)�v�pc�!ژP���Y���-�#�V/�>Z�!e��YQ��?+�?�>�ٔ\�=�i�p0
QLz��*����ۼA�	�Ōu]��=^���$D&��C�)�]�(�k`&��f(�lQ/ُ�:��<�CP��,�^�� ���!6ԯHf�>70I����K��.��f3���G3��{�8�Z�)Ĵx��-���ӟv�翹a�������x�ш���L�-j�v	*� �^\k��w:��=C�d�!æ,���i�H���>��u0�m��ƣv��q���A/t�Jx���]8õR��V����!��_uw
ÐK�A�/`��g�%۠,��f�y�MM��V��5>_��N=q�j����]�����؂����G～������kN~U��%�M�B;�m�=,C��LΪ�^3WoHv�}I��_~s��ZO��z{ɩ�禪i�x��{��bT͘�7��K`6�C-����;-cy���!�\bz	4/���㢗�[����1=#?|g������P�v�!��Ȳ�˘A��z��yV�d����q����T<�:�6��'�o�+%��A,y�i}7K�=����\"�f���n�6�wj9e��$�鋪�ts��h���"��U����T�����7w�jd��D }��^���j�1����#��5�w�w�,�=�>f�]m	��,#s,A��qBeO.4�1YP.4lx{G�ݜ�����=���0���n`w�Sм�e�ǤQ|�	6�5"v��6��ϥ���,�72����C�8b.]{C����<�ǧ��Q��\D��0�&V�΂\Ӭq��������{Q�V�B�<���L2D@6�q�Z�lw � �K$��/q2"k,4#�J.�kqkb�4)�lX_(W���e&-���k��:O�^�(\�̛�S��;ۯ�u�f.l[숝ua)ʇ�4���nc�:��O��ȋ?}k�:�yT7E�}�史�{���M�f�v5��J�|1�<�PW4[R��9��=^1a���Za�	�%e;L�����+VD>�ACL>��7$O=_v�r�_xŧ�ר�ꑧbXw<��y�K�ʟ׷wt�M�r������PE��dZ�{��P�Nt�,�y�g��ǒ�I/a=;�\�V��7������A�\�_�v����<æ�Cj�Fz��ST��s]�JN*�Kq�4�%l�����@qn�?�v��pil�L�8��I��畻����aTX�¹ʺ=�S%o^C���v?�̠�򦁺ԟ������l�etK���v�9���ʥ�Ql�t�d"\��¶�qnf�[��>�� �＼������ �|��� ��m�������׾���w9�0}a!��a�:/S^���0*���"�v��h<��E��YaS�[��������:�;t��KC�	�?ޙ�`����>�7�D�y��oԁ^˝.��l����P�}��ǭx��!Z���EqF�E�~5-ͯ��X̋{�'EiX\Ș�a~���,S{����Ky�q�n3�4C��V�+��"UY�O���1�������~�f��O��]������oMiՌ�8�������|��i�|l�yͽ��M���ƼUC���k�A�����t^&��5Ю	�7#�J����a����s��I̱��A�Ķ!�!Y�S��K�@�m��L�R���*���I�4�b76b��2͋\�zpG���,h��g�c��'�~��s{�����
a�B4�O����K���ӯ�^jb�w�(N���.	��"W*^����� 4�x/[x��� �M����I� T;�Ƿ�h������S�Ƭ�2�tD�V
T$%2SϚ�rq���e�C���<�4�^_�Fc6�|�=�eZ	�3p>*M�7W�M�
c\��Bٳ������
���o�.��>�(�c�ό&��x����g����m�ыM��Jiµ2k�7ڍ�ܽ�v�g$��y���~z�s7�3�5�Wѧ馂�Li� @�����mb� ����D>����ύ�&S.g	�^�E�4�j}����t�vv�E�I5���hb���P9焢|y��r�ş�wR3r�|���L��g	���!�#�7o�6Op��`��&�s��ɥE��B��p?r�Q�L��s�+�:������cʍ7U�+�_�1e���.3������><����a	��o=K�uBT��aƕ��,�im�G2��U&����fV����(t��ҡ�W�öBZ�!W��K5۳̼�(��̈́Sr*EO�EƎ= .{td�����q����P/n�|`0~�hs�j�C��yL��tD;�k-�u���C�e�N0-7�U7;��%�^�49������,��X�q����kNw���Ex`��~�$O�@���=q����Uع�ߧ��Ǎ�z��+��s�/����W���}&�-k�T
g�^甘�~a���P2��Ȏ����2_ޖ�[�K�;�N��g�W�Xe�����ٚ��8@��0O��C���|`o�>�X��Q�0����,�y����},�^��u���?{����Y�4���P3�k�Y4r˸�꒙ebO`�V�)HT;u�q�ٿ��=�a�W\|=[�����E[��\((Ƿ�m�"��\3A!Wp�Uz�Wt����vd�/l��Z������
����Vۮ�Φ��������R4�P?��^讳צJǀ���t�*�NV4������r�\������e�t�/����j��>{�}���e\��)M��2��\k��ܮ]�Ù�Z�x�H�=�V.&z�P�_�i��!������E�����d����o�gi�E���F?,��
��%��2G��ߕ��^=�m4���.�_e��4�q�:��,	���Z�D��I�5�<����倪��MJR�hy=p�L������������Ô(Հ�Tt�z�,{���A�>��r	xkՋ�ZX�1.�m��%�aU�)�"���OC\<��0hL!��_��ȿ*o����/��l��R�W���e���E�������6�zh(��!6�K	�����������p�O���C�+ە��Bž���Qj���,lj�����K@;捠��0t�r��wW\1����Dlq���wf�`��x/����|�S[��Ta�Z�cH�~	�4$��.|����q;�ؐ���+Gd�<0��#��ֹ��œ"X�����*\�n��y� �@��� ;apv�J�+򴙲��_~j�0��t��F��N�1��r�FA�!�{�t��k��8��B�`���u'{��7��/[;C�^}ܷ�u�͑�,�j�N�Q���s4�\�G�\��\b|3���>݋�y��j�r�����W�� �o7�I.DRX��˘o��8� ���Y�~,R ��a�3�[�����&}�ͭ<L*5�x�����!Ƥk?�[�utP��c�~Q�9�W�G��&�!Y�����������u@lȆ���aٍ�k���殱�cü ��"T�{��J9�02��2ċX��b��XW��;�E�Y���P����/kt�V8S��/�o��>�z��(ax�1D*1Խ'�Y0��u�&�^K ��E���Ȳ��謏D�,�;�䣰��`��AcsW�#�6>[�c��4��R���2J-�b�Hs�ٴ���[pz��denf>�jᷓ1P�5��S����Ņܣ��=��?�c��! վ�(2j�Ȓ�ծ��L�SD�~�wp�C��ϞOhzңnr�R(p���"�c� ��~�>���f��S��wv���#owE:�E��
��V~���_=�����J�}�D�AC�	�Й��	���%^I���L��Sg��#ޘA�y������eG�2>�F�U�m��ȸu]x��R.%:i�A��J��n�>�3k�ɗ�rr�՘��D�7f�F��=�4�aX#����p�շ��ޢ<0�\� ��_u2�'��ek-���v�V���%ъ�5=��p�Uns��fRs����=w�|���<����sy��3�U�X��?0�7
Ą�`���0��7遛|��s��"�9�R�Usc}dC�������nV���r=��C= ϧ�=�t�+L�;�̥�Z�G$�9�yH����N�x�*�r�S� ςߋ�|X��^k� �(���GQ÷�D���4,�La�%ϗX9�S�r��%��ZC�i��YE��ώ�r��n �ȝ�N&��n�5�@	8�R~Q�XC3�T�Ƴ��iL%~^uﻖ���������!X�@�����Rf�E�K�d�2)n=mG8��&�(3�aJ�9��<��� 'Y�>S�v�Mn��X�����4���׿�����s$�Kbis�+R���=4C��;;��~��_�	7J�h�(ȧ
�3]9,�N��[�dR
�D�t�^���};�ߩI���]��S�ˡ�1�^׶~���Чy�;�d"��Z1��u�!�h�LÔ�Ma9��U�H��%�J(��i֐�q�_n���آ6;�1�7��x䗨;h."�y�z���?�@.���3_�{�n.���̫��jŏ�WN�N�C!���*u���}[̥�8/��s"M�ʑ	f���J�V������R�p��sw�m[Ţ�pd$���HDW�!�����_���7u~�ޱ�NL�X��ULe�ỵ��v�@���儒���@��k�0�^�7��^Yѻ�T���l�Y9��|||||}�<�l�3*W��7��C^D��:���ʒv??,/�P5v���~�?u��K���D�i�{]݁�;�����v��!�������g�b�θf��%Ć�/��M�0/��4��^��˜�	*neo�]�2��vH	�*�.)�[����R������gy����������B���>�>"�[��w{�t?DJue*
�UR����l�Bb4{��bo�w�7�������2����/�@�i1��t��E�hs��sM�:U�^��t��%��vD��:1��ʘsȷʷ��nc��<��2��Ƕ`�ԞI�}�M��ف�"��a���{����U_S6��<�|�LM�>j7ᆓ
���o��9���O.lf��,��s�����R�p�o��,f������v�c�����dSs�	���2|��qvR���k���|�="���c�J��>�t�62�[.ۮ3FE�f�O��U�S �O�ey�Xs&�W��a(%�T�y�.������|P�G�/ֽ~w��A��˸%J��J����e_-��0WD�6My�6��ij�%7����V����f깝6)��W.��Ǜ@*���Z��{���өE��k!���R��gqJ/fq�*��
�kB�y�Cp �(� ق�9�9�`��?��|~?$L�`]�0�.fI���o?��ٛ��	�)�Fi	ئ׵��͎�ڸ+2�a'���xP6}�v�T�?/T*>c!����r���3I����wƝ�,��dn%SkC>������&&��\e/�NϼIZ�o����$�-�0���7��)�Y������ ��"X�+嚢O����g�S���,Kx~�"���Y�(x�J��N�pr��r�:��� Ę��tD[�<S�z`�l^<%�q�p��M��Tʔ��f.F&l���p�S�V8����
�<��H@�>m�~=IҀj��ObH�������Fbr�Il�c�P�V�@�qP)�E�J�b�+��%�Og���A�9�s��3�>��%q�w1!Ϝd!m���ג���>o	Mg�&@�P�� v��f"�����ׂgc���V#�M��E�]|����i���B`I�U��E��'���S�J`�U=o$�tLnl�{�o��eU
��½{��r��R[���I�_@"E��f̢�y��q��g+�Kv���t3o�l�*񿈰������IPm|�����x *x4��
��c�۲�c<�AcMF���b�N+k2���%���O1�B�}|�*Ha3I��f�#z�c��n��,ᛳ��Ԭ�� A���U}��J�~���^J�y�J>�'$��Gx~e��㴅��r-{�K����-f�S@���u{݃�0��W���yy�o;�����0��R��Z����U���J.���L�أ�C��c��;���47�C��ڤ�;��;Q�e�k(��oq>8������T45o�C�Rq,u��{��+Ҥ�1*��0�lV��A�w�t����S	����T/�YF^���0T�#�Z�/N�[�z��*�or΅X��}a�01���uBb[L�d��0�ܥk��S�Q/�n֤�q��V��[��-��`0d9	��������v�s�����\���+oaɖ2�4h�'uz��Bɂ�wL0{F�J���?���GM�L����M���5��,n�Q�~�p3�����K?D
�o*�i�P�6/׎%?�#�k�*l��m/��LlZ�1��5�e����~g21V0h|�%��- �$��h���]��c�C�4ſ��g�������j�S���r�+>C{f��9,%�E��o4�0���O6��=#��;̪�Ռ�h�ii��~���ϗ�<t@����W�_A��`[J;K��3?b����eM�%�u+�[�r�sj�Ӧ"��v{1�g����:�cÅt�3qX�4�b)�K*�s�#3�˾5���Krus�9�ki��Jfd-�ǝw�煗�2�y��GB�Lܼ�s1"��v3�'N>tu*�T]��jd�w��sEJ�c�6����,�8�5
�gx���Iu6k�T��kP݌���7����2�mAt٬�8Q|�V��'�Ϳ�Z���1�r������$@�ټf�~�/�����z"&u*6���T������D�����&u�Gf娥��\��k�yeҘPV�*�������Q�"�ٹC0�Ʉ�bÊ�]����n����r�dC!S�C��>��uz��X��0n)w�#w�%۾-w[���e��rӯ�%�����y�O~{5]�R׳�p{J��������[����	w�wb
�AܙOp�R���S�SԳF��ի��{6	ъ�7)]j7gM�Y�a�\$�˻j��5�`�2����g7�$�,jݓpL��U��ص+��k��=�:�m��r�!�R��(o�ãb��y9k�7��Z�:˲w�5��S�[��P�/�쁍U���F��7���q�C6��ܓqaz�ZowoM5έ���N�4b�5�7Z�����D�H�{d���t��4�> ��]�����w�/l1����Q8�:�C�	�Sa˚W�}��hV
}�o�K�Dm���,�l��_u�V�%���7����X.:���
���r��?��T[`��<�96K��׷FuZ
�q�Q%)�b��-�8�d"ƹ�� �@g[�60v5�徎�uGV����.���7�=������\*�t{��]U΀��\�u�
s�ݖ�
&2��j�'��ާ2f��|L�,-øٽD6��U����lF^X�t�=g�=�YǛ���ҹ*ct_b�E���"����d��KI��AS�]���aKp��'q'���jKfZ��uR�Ś�g�زZa���/��x_�--�yu��Jd�y�Ȏ��i�w���,�dXTy�UE}��=�1��St��Tʾ�nTQ��us���L�-8༭w��Ɉ��v�w��"�s�ۅ�56�D����n7έ�ۆ��w;��'��n��/)�� Ӻe٬����輲�6�=�`�R:��t���]���0�|wGA{�;�\�=���/�Aܒ�}7K��Y�z�>.����R�[ei{�= ;�O��p�ݏbڞ��j�ٹ��5�{i�T��Sib��C��;�T��9�+��ڱiΎ�(��G��]�����#܌q�f�$�F�v�;%�Lr���1���WZ7,�GUe�,E/
͐_�^��������X�(���(�j1���|߽�߽��;q�Ǐ=z��	TIRAd�hѪMIF3~oo����8��ǯ<x��רt� 2	$�����$�HIӧq�<x��Ǐ=z�����@`�Q�"�*��~m8�8���o^<x��׬� Z4��3��y��6��h�E T���`��-�Xō&�ZK$kEm&ɌX��TT 5���`���tX4����$B�MQ�LQ]���W*�����v }�SQv��s�9ۈ��o;(NGo{9_aL�n�6��-|�mt}�av\�!ȵ=E��۴��d�nO�d�Ɗ���i�
gf|���>/����ݺ�w~~_�[>U��X�V!��ν���T[n�q���eT�EᵷV�PU��mL�v�V�ݦu�{�2cV�۟(-�1pXp�H~�c�g��:�l��;�\�Skn�V�:�w5��?�܉mO~IM2R�<Ӫ7ڇ=����{�`B�D���&�����r������@�q��\�/��$�g�
���}4�YO��n�lW���Ś��?9�յܗ���N�q�P­!�1�
��'rT8�) ��0P�J��a�^1�9�w9Y��w_BFx���or�"2<�>�����7�j�i�Ⱦ�Nm4e�\�7'4,R$�V�a׫���O��-Q y��h�1���A�\<2ש����Vv�oKI���}�Wh���Ϭ=�0ni9�?8�^HW*J�C>�,u��?s�k�9���=Ϻ����5�e=I����}�fG!�����|j1��;hA�����'���g������ǯ����5n��t�r#R�(FPz=x���z�s�Ԥo�F]7z��A�¿9~>R/˓B�72'��,V��������_�×b�Tӯ��%.X�!�	�;48�E�O3{p��ru���D�N��z�L��]ʯ,��2i��wv�V�[S�]q����r��Y��o3���T�B���7r��r:湬���O�c�3���jw3���x����D����s��fs���3���C�OxP���>7���_���HqEI�K����j�j�C;h�<A�˘��F��/���x/�ݵ���}=�n����	�א�&���U0����%݋2����Q�o��F?U�A/۲K�	@A�+��5+V�6�։��ITP���T5KO�`�'��C���n�/����V���2b��=�k.k���52��ID��.�i��l��sӽ��$������;ٳ��Hf�
��oG-�Tg>5�A�,�,h�Z�F:�H���:��P-�6K�]�*�ċ�h�Χ*I���K�t��o����;O���?~a���}8�}n��u)3
ti�u9S�@u[|���B��A��|��-�#"w=�D�VR��)�QO��ʡ���?�_����D�����.= �����|��������_:��&8^2W�"��I�
]��xV�m��=ݙd �+����3���2p1m"'��ｚ��F��֙��?G���:
T�#m�{�C����Q��9}E+��8��lvJ�\-0��V�C�Q���j����Q�r�WJ1v������c*��f+�������uȁ�I���}8���9��r�㵸M:9��QG}���������#s��{sƓھ�uR�����m�t��6�3�x�ic97k2�_�b��z������I�Mf��-�[B~��v2'���d�70��ծ���\�P��^Z�F#=��RfZ�w�����0t��o;�W}�c6|�T�3�Źn={���P5�3Eט��QaB�L�9��Z�|T:lriV�s����{�e���<;���ls]Ln�}"�tqq����iA/m	��ي�?|�Dq�l��)I���{��]��C��_h��an����t=s�^%#��GMc�&<'(q��}��]�f���o���1��2��zC2�:����AUY]�>��"e=��CyĿ��I#�L��2s
�+N�f��Thp�C���)�%���? �+"�m�3N286Y�5�x��ˋ�Y��hB�F'�TI3����^�n�'�����Bo���O-ĢG��ͬ�7�>��&��Z��WޖO-[����d�+Ț�M�S���9/C^Y�s���M�]�������p��<��~�He^��Ņ6��c��P��'\>�z�sr���=]ya��x����VM������rG~ӭ�q��{��J�*YG��U�����[���4v'iE���Kp�M��>d�U����J��k�1/f��!г�&=8m��m�Y�^rE.�ʔҕ�N��U1��b��sV]�����c���[�{����L�D����OX�!Ҍ�8� ���� ��z�eyX���G�J�aMo=��3[5w��y��:�^�ᩭ��ń5��Tx�&�'��y��҄�P%�K�-�"��e�FRu�׊�gs����I���_삾���Er�T������B`$�}�"�L���Y��f�̨�y���ᴺ�ģ)�cθ绝>w� ��.�#����j���<Eh+_�sp�Ws��(�oS��yb�u/��;�ׇ�C4 ���`��i���U�Ɉ����]o�۳�8t���]Ď�^���Lb}k+=%���S�jזf:���u���5�sUj֛ގ`����S9�����cp�&��*��Q�b�T;��@�E�_j��񱖛`ήw������è~�1-�7�%��M0�w)Z��^��iz�鈉3ac'әv��Q�a�:r:'�Ct��3k��!�����Ln5P��n�!��j�p�5z���ǣ��^=R9�3�k�l�f>$B/0��^��:}���l~���$f�~I�>�zn��Cn[0z�e+���w��&E��̬5��/ ���8N�]� ���g����cml��(��n�IYyA:+"��Aׯu�G{+��\0��V�p����1�#�En��U�h��Xx�������o��É^,C3;;8C?��e�羍	�����ޯv���Xh�M/��+������)TN���oFB�u�r�VHl�}V�u�}Z�MC_���Q{�m5;�%��V��j����@��i�r���l�v���n\���%�5 �==Z�c)�,�O�_$Yj��X��V�^S�Lp|a��y]���?>SԨ�>�kZ�T-M�-���4�X�*�������ľ����e�@7��UW�Pm^��9��`w=����!5�+$؉��sn�:�X�ؒ�ǧXP=Y���'+��?U��2�1����� *����!��ȫ�����ffR��� LI�r�,��o�ųw�(�}j/l��Sۼ	
g4=���ñڙK��."��UP4H��y�L��DIu`�ʁMa�M��+&��;#!��N�����]۳�ɶ��;�,�dL>��X)���GuI˺b�C�|)QK�X�c���v�2�gF^jm�嘼�������h�ˬS�vc��W���=q�O���a�{��T�ֺ151��c�c����TnTYY����+�-*i�,k/]�D���J��Uh�u{�	9��^����jv�n]�c����F�D�TQ�\��O!�*>�Д��58��`�-�5�e�������y���wx6O��ASL'��s<]����������uz�z�T(v8��E]l��������·��p���ڡ׳!'�_�����B�,s�&�dN���{`�x�����+4n볳Ǟ"9;���M�OI����cj$0��&<B��S�t|�x-�镋��YN�;oC�ة��*E�ԛá�Y[���� δ��?�hC���8k0�+U�U̵�`�f�����]���Ȍk�)�[�`Hqף�sI���j�=�,j-c��j�kޯ���y�g,��XQ�.����6���f�K���N���u�����c�뵿u+�`����jҲ0�1�A��"a7�P��{Ng#�*���'v	v�-�b�s�6�]��0_���2��U�KO�l�`������//�Y��Sz�YZ������QyR���b�qx��K$��Q��y4˜S:~iw��,/�Q��DI��-�ʹ�/��{�~���̇r6�z	�l�����Zs(ֳю�shlw���#��/͢���r��1�$�7v.���)��i~�;Җ*�k&dG�u�^����ioWg�7/X�~����`�+Z��1���ʼ�.�jS���ˁKX����Ю�*T�駴�)ʾ�[�iL���LF+�"Vvٻ�`��1gva �}����� ��Y���7��t�e�Ŭ��'��框"2�	FB˦M��V$C8�J�U��?PU���m���C��l&5iP�aU��q�^�X�yA[#��Hھ�NΆ��dd����n8S���tݯ��"�	L�N/��ن��P�')��{6ߧX�.m�S���n��%8vA�_X�6`Fl�,s��Y&i��7q�J����@۠0���O�]^����c��h�I���#�m�2��v�]�0_(�ɘƻ��3�5Ɠ����\�w�����vk��6�lE��Z}��.����v�ŉg���q�q˝a)d�yjnQr�<\�UE�^�;������M�N����U�We�#zא�����\�2;FT�qvJ�,1Ls�8� ^�Z{=:�����q����t,�ĽЩ�0|a���<�����ԊM��Ɠ~�Q^�J	|k�����.8;��ś_���v>�5���Z��
��0z�-0�;2�<�4ޥ]�kW�^�%tt��<�AI��N�zs��q���8e��	������5ԉ���2��~"����*߅~�>�;.YɍΩ�!KA��]���Z
�fSY����-�ãV�� ��+[xFU7l�8��m��6m��ڏo��M��f�#w��M	����#�sj���H�B듽�J��_���%ثݔ
������y�ޓf�[A�Y����3,z&��<�_?+�7�χ��-�<
|����dZb9N� ܳb��0�
����\�����	�Sk<�7^@f@��B,�*4͛�V��2ӏ5�//b5cS;4�S�᭩�
�]�Mq���Y!
��M�7��P鋇�ygJZ�S�m�?Y���>�X!��=�e,���O�`[P�C2�P�'\>lS	����8!#;���.�(�3�-�X�L�� ��{d�d�0��D�-�ej�
O3���Ǧ'O6���rB�`�5�<�o-ML���4y���@F|��5'ƿd<ڮ�Y��������Y��S����?yL>-2XkR��U�M��P���}���"��.<�� �-�5���s�27ܼ��N9�^%�}O,x�I���o8k���5����g�< ���2�l��:ډ�7!�/��l�w��P�9U)(|�eX��P1���6��,��z��nM�u��C��F�����k`d:���7݆z\
�&-?5����	ߛ��k#d��wJ�������ٹ�G]wh+�)���h����v*Βޘ�5h1No_q��,TV�Ϫ
�����cuT�G�����bz�L��Ӣ?ITy�$�ᨳ� Xj��fT�p�����|"��,޳����ǯ�S7�k7k��)����������`=d�>3�a������#Za�:�UN���FEp��ը�+�j(w;�D9��3Iκ#}�mN����"}�-��c��/�uG}BA�=��(w}>��m����}i~r��������M$-썚�Ù�c��D���	�*�WE1�mnؤ�x{|��z#��g!J�7VX�~���w��{�T`(���4s�Q�!�������;�<�dY=�g؈�m�p�Ul�P�:=-=��oW��E�,t����?-���z{=�3v�u���\!��ؕ��F��m�6��c��4=`{����D_="���qi4�ɨ��Mio�3���6逸~d^m��|�u�&�d�F�X�ɇ՛��5�-�K�+��E<2�<��t��'���o��w�p/R�B�e�+���BR_���>�7Q��x��,a̻Q���s��^��IaR��a�y&��ɐ�G��>�j=��w;�� mC:x2iX�$����
ј��O�����<0��=.�x�}0���ߺY1���pѼz"t�6�����$Fy�'i�f�S��T�K]���݀��x-\o�$��˨�{��$�G���՘�jp��@���9J��S��Mi��n&�	����%�
����8��V�7f��l�����7�7^{%`|bF1�`���5���^r:�5�D�Q�I�>SMR�I���8Ξi��= ��h����,zV3�5��c�S�R��EBǐ�7��=��q4]b�ʊ4���O7����B�*L92��*r�D�M��S�d ܉��ƯѬ�9=��	���Bb��J�]�q�/�i�@��J�7[\�:���}����_���G���+~�Ϳ2/�
��?%���9f4�����x�2���L'��-��u�%��!�=xND�ީ;9�=]�5s2!l-��c���������'�p���Ⲉc�P5�����P�_a7��t=�d��e1�"�����k��bq��UV���Ϟ#4��W,�����_����>U�#���m�z%�-w���}��cv5������^c2���"��G�n���Q�Ԯ�o�F��x�V�uޠN���;T�)�0>�0/gU� rJ�eu�t ��}�UE���4ń���}����[P�qH&���m��"@�Y�J��c!޸,g;K��2���F+yG;�W���H1ҋ%`:��e�䵪�T��}��t|�<U�W
��3��;��E��k���:sM4�M����V;�+��-{U{�5�M_�X��]1q��2ʶ#ɣ���T��&�<a�����K坛J'XYӒ�'Ue9#��ZR���M3�`���Q��c:p�u�t�+���Ϊ�ۍ2�o۔�6e-KF�cm��l0e+���W2!�f.�V���6�\{�eg!ɒ��N�Z����r�:�\�BCn!ҶeJ�v@k�}���-��AEU��i�9h��*�V0�r�¤-�]�=!IB��9H�a��y��'v�-A4i[܏�ܣ��
�0��͘�$Fd��l=M���e�}1Ѧ�㑲D.�{�����wr�t��w(���_HvB�Ŷ6�Z�û�}�=���%L���̔��t臵�>)Pw���oܴ�w	s:��ԝ�a��[�ӛ�����؜��4���as����sf���4�0�<�YJ�n,Ǉ�$�r4l�̏]Z���:�/�#�N���P~��Ƈ1e�����^֒�NW��R��r�`+3���A|u��'EN҆S-w5ŗ�����Gͱ����f�s����/Ho�s��L�aΪ��qvP�M�`0�dؒ�.�MT��ۿ/Z��t�����TD�������J۶��a�.��5�$Z���T�P��x]l�,*�q�I�5jy�A��v�e^�*��8(�m��ӷ������uò���5l�\�����FY����K$:�˫�k��ys��u��i˭`��Op���%�����i=6�k��Ӑ.�i�{3hl�����_MAױ���{��M[mR�L��ô��s�)���ի 2�gV-&1���k*�O';T]e[ƚ1}	�2��o�۫�F��Xܙ�j�W�_b��tʠN��:��Z��-i��5rKK���7��<��y9иF��7�!���{ի%U�1��Ѕ��j�:��@���fU��Y�Q��mG�q^I�H-���4��Z��zK� �l[ٛ]̝u��n�r�>���b����߳��*i��u����.y+{��ʈͥD���5k�ܧOv��Y]���bl����.�#=Q\ͼ�.� ��x�6�oW��*��0D�����ʘP;�Lۢ�mӬQ�C-�p�3�f��Vċ�Q�bZ*Fo�2.�|Z��-(��Y֠nr���8�9��ٛ�������٨��u�ȷ9ل>��-j�y(�p��+n�Ox���&���n
��*����]n�nZޱ΂/b���ٶ�to�-qv��VL-ό��R��Y��ˑB�in�f�_=�N������q$�$daBI7���$ 22�o�x��ǎߧ�<z���$P��#!#%bSR����?�ыz��8��Ǐ^<x��׽H�J?J�$�u�D�!!!$�E$Y���qǏ<z��Ǐ^��FE��A�HI5AQ*��c�M��<x��׏<z�ΒH���$I9�����ە��h��ͮLI#�W#L�b��[�1�5|�ےT	���v�h�]1P�u�ޓ��6H���{_�J,;�5w]��Ov���=�s\��3Q>����AW-;�E��V�L�q&�m&ㄔ~��&4P/C#AIa���`��n4d~$C�� �#FB���̃v���A$6zdT�\t���K�F��-�L�2�T�.�݁^��� �͚Fu�_a�hēH�#FB�/�#D�!�)$dm�Y�&aM�am"��1��*$|R��m�����PDƚ����aƐPF[	�!D�p�E?6��7�� �e�t(�\���4���]�13e�\m�ږдlKy�Bֲ��ϣH*b��c;�6��##cD��4���1�u�k;n�����"���z�Dn{c=,����f0!&ݢ�p/�)��C��gtv��vR�3���`����U���q`�I�&�Jq�n����j�/A�ty*��	���'�=Q.p�j�2j����ygw&��n�����K�6?V�/1� &�w�׭)T�����Q)�-���:�c+j�Q7�����2�6!(�'��q�&��*).�;�{��ě��ǳ2K�.�~�̉�nB��[��o:K�D���7j����&9����qJ�g���2��@t���a2tx��U?~^�3O	ѻ���SiwoZ�ݽ��Z�b-��{)��7p]�H�cY/�)�=q�ܧo�ʽ�f�+u-�R��)�94C[f0Rى�[��k��_k�b��E���d���M�$e{z��K�9���<�?c����W�bWo ��ԍUrr�0N�-�=�����1��ŰqUN=;V��nS���K�v5��a�0��{��뗗&V��}��y�o7�����#���B������Mw.T�z��z����=9U_ukn�)4�X����*c�Y��ܤ���Ou+��10�N����3ySa�7�Z�q�^5��=���� <A�q�uD�+Ի���p���O3__nޑ[��FC7��Y�.g����P����f�;�]��u$3%JC�}Ǽ����&������>��{�}zML�@E�\�-�#T�̭�	U��f�I�6'u��1�>y��bU�	���ך�0���a��3�h�ܛ}yK�^�k]��b���J0g��ϙ5B�L��b7B��x�˩{��J~�����#>T���|6i��P�S��?�-��
k8���;
cOV�ս��˲2{7f���u5l�]�'1�Ǖ�K8�ˮ7�����ǧ��9��/b"�*ΡXo&�b�슍�aT�J�32�J=K��V������꘷��Go�4�A�Oe�N�L��|7�v�˩աyCp�M�&��$隡�y�+F�b�a�N81nc�S�^�H���}����~?���k=�|�خU	h������8���e\m2�=�y�Ė8�L�d�6��&9�Ժ
;=Uڞ�<U={o��/���^@(��<��l)��w�p�Z!F+�@�ԗ*V�<������Ŷ���WM�1T��E�p��v���b:��_��'˜��5�邓�����I�Ut�iB�	� �_���5���k14#�f�ѫ&��غ�}��9���X�b�Kw�9����T|�g���1�!6gu�2������Ps[�}���ʔ�do��r8Ì]02���4�w�X<WT�B_�W�׻@��{��A鎐� g3���L���\����F�܇��K0G�ߩf�碤'$�XXq��f�U@������T��{��{C���~�QHȱn+k�wI�,`�*��w�?�|�����e-���k#w.gV�qL#,l�z�f�uq���[O{>�딁]�'gҭ�]yovtw�tƻ������}+�+O�)j��X��d6sj=n<��n�x��e^_V�O�;]�*a>���8;ǽs������c#��/y3}��u�y�O��U��4��
��M[MOD��l��I��fL����On��Y�.�0�X3>!Xv����g�>�Z�wn�6�T.��n�66óXi�\�'ZFm)�e��( -��i�Օv����@�ϡ��\����\���<�(`��2�:x�#�y��U��a�]X�����!`^�݆���͚g6vF9���(1��\��,�Z�l��
���S����/�ȋm�#
�"�#�Q���ʇM�QS޷�O2n>�Oȶ�m}�����Y=A_=�p�
a� �!D�v���]��ւ�vXͽ6i�^n`|��!�r��2ُ��h=ÿ�[@GxlS�����?�}�O�JgY�R��ܖ����D�;!����C"7�!l���)�TLls���6bs�y����� ���^�0�R]һ�����͆�q���LkLgv�����9��]��7ꤣ�.Ơ.�u���D�,�i���F���{Q�\3!�t����HMFﮖ{pC�=/��ӎW�J�U�qu�ʉn�ߋ/�^��U㋭<R٣o�W��S��8i|��9�sL�z5d�8U�S��W�� ~?���Q���F����n=ٚ�|g�O<eܔ�y=i8��{�Q����m��;��M-z�UY;L�<�p�k�ջ/��[u��.����3������r��lؖ�"�ȥ��'�B��䋥���ab�0U��`���[F���my�d�/ݚ8�B�V�wV^B�:�Ԯ�L��xC�E�S��#������>�Y�����t4��@n��>+�^��i��C��<W���F��Vʵ.�N]�+��W�������-Wo� �ြ!��I�K�,E>������ղ�]>�-�h��+�@�#ג�r9>�g�l53҇Yk���/�*�ʟ]B�WxGH�3���I꧇7��']Qݗg"{�	֎Q�`u��l����5C���ƞ�3� ��ჭ��[����[��x�b9Q�n��U�r��~'WV�٬�r�ߦS��,Z�k�U��+�Y�dx�����Ob��.=��˲��l�.��;%.[u C��4�Y����fu������v��K��x�,p%���k�����5,�s�����M��߳�|~?7���'v�/�/@��@l����d�[��$]�Ϡ���Et����Ͱʛ%�7�ۖ�I\�d�2�;!���Z/�c��j&��i�q�\\�Gjk�g~\W�&ۍ�=+�륈������=Q�d?7,�燼"�ڸ�-"< 7��4�^����sַĤ�9�(g�l�3M��L��q���aar�/iق���2�U�y]�*V齛i5S���������Ȕ���a�>P7ݾ`VlWd��%7q|=����(.0T�O���;C-7�F���������a��L��S�p^���_�m`�ӑ��ޫڽg��y.��&��5�f�.ǌ�� �i�a�l���v�oe\XCp��S|��&A#��{<�#�ӝv�/�����g�#��Q��20��,�|��OY��"H�K��P��E_2��'n�ddNi��ٺu�z��WW�$�3]KDw�V�O5�a��ǃt�H�骶�ȸϡ���++I���wT���I�$��,���Je:��5���,�yX/8VW�{�\h���p�9j-v&c�s=�|���1�c
�9����{��A����`Z^*���
��D��5� �KH��]s�(H����+}}v\;�a���?G�]b7{��7\;HL�I��/uD���H#����oa��Ո5�#�ҭ)��
e�jܮ��㗽�������ɯ���*i�ճ�^�
&��VE��lu�ڻ:9��9�V���"*9�d3�9�����=\JEJ�k�Ѵ�i�u$o]rz�������_)�9�G�Q�s�U�K�hVS�t�ӭ�zMӺf}���n�:F;R�t���di5���y�xޥs��m��71�'s1�؜@6/5`#f�i��8+�GY��'"j#o�g&h�s��J�C]`r��b�;�}z�W�(���Jɍ4��g.��酹R欞�b^�
����hHވ}�{�o�	����SE}��u�j��1�(�e�t��+Bg�)�����cP��,�0XӃ�ތ�Q�-���ل�:���������A��Y\}�K�ɤ7uݕRj�\�j�qav�
�G�6q�\������9�Wu\��92��f��|��!j�Lc�y�ûZzZNfww��v|Q54����[#c���8����0����r���x�K`�ލ>�&5���;^��z`t���:8�\{N�.���x{�8*f���E\_�/�#�]�j�������q����53�=�Ж[�=4س��lFV
g4�����`Ƚ�_M�di�9%�ᛣf˱�,��Ѽ��%�o�E>�3� ���Y��Vy\�J�c	���Z�`�~0����s��Ѽ�ե��m�n^:  ����S�:�hֶR���N�9n7�{A������^�i/e3�}a/@�f��-��0�������tz�s�h��8���m���֨����ߏ�(���Q���Iު�?ҟG^�j\�ޯU���ffὓ�r�S�JT,���n�:E,���	sY���f X����cTVh����k?.�%UHԯ�o���n��������q9��ݭ��f-
�މy��3�:�f��7���y�7M97C����k���؏s�j�lع_pG&�ܸ�� ����7㎃��Q��;�6��#��gVǯ_VL����x��_W��}S��t�缥<�^L��A#Gwb�Tq����YX���T��&�����
�W�(��ns�t��s�1}�g�1;����Q�*��#1�m�
ۼB���N�u�>Eִ�e<c��Q1٨���_��i�{G'���Cc�C�����l<-c���e�ɳl���_ ��]ܻ�嵁f�D��y�~���q�7�=�x��]Xv]� B� 9�Uܼ�E-ފ4�ƫ/i��Ӫ�1�?X�ף=�2�0�r�qJT��sms��8�uD��ȘNǹ���
܊��ۓ�����f���ϛ|�;��#^E�KGd�ty�8������7kK����;��=A�t6��z��
���~v���3?~�'�U�q�PN2ELK4Ne�5��?�/�c���/��_@x*C�#/JdO��vu�#[a��$aLNdN�yĈ��Yk�
s��z�,�R�"��4E<D���e��hqE�X���I_��k;�l���!�����(=��S�g��y��\I�xhC� ~�����L��7��'3�O�ٻ�1CO�;����$�s5[�^h-bی�{�ݶs����o337����1�ts���goZ��"��ǩZ���+"|W��:����M�LE�Wk�Wuf��46|G�z�Okt�Ʀ����-���H=KDS���:�2�j��s�ql�ͳ��9p,B�=�:U�7��:k��Fo73<�si�M�ֽ��Z�^OM>z���@
ϡ(�?�\K�7�ywq8�h^�y���z���^�6�_�Qr�ۖ�s(w�<��׈Y���y\�ᵝ���ǚx�}�:�%�A\FF�j�9���u��	��Z�aoozf�s��Auy���������� zW���E�}�=!�͐�w��UJ�o��wN�.$#��6�q�R��Z�W�DѤJ��w�'i�쨛�Tn^��]�j��lj�?�%�u;�<�`���T�ʭw�+u�X�X̫�/fq&��7@�lL'�3��Ϙ#���j�2�����?
�b�γe��ݗ��U���+1>ၱ� Έ�w��7B(��q͕�m��c��̙�;�yK�f��(��Y���\��lo��\8��8>�+?R����梯.��(�p�1#����(���J�ܜ�NdW��7Ǜ��F%;�j��Y�; ��fB�l�'/��iD+95W�e-�ՠ�n����飳Υ����I�m'c�Bs���K�O"�ȯ����j�|xۭP�=�;6u2�iLAܥw(��}��c5��٬u�p�V�2�c-^E�O�j���D<���U���ʫoU���;���	�݂�իט��5#Fgb�!u���i.����Ζ�]w��Z�7�S�omPؙ�j-U��w��H�&����d�Z�q�Fi��ɰ�q���!�����]�\�..���x���A�#���}(�qD��[�	���Ew�182���u�zNq&�]��FFj��g���^��kW���z����/�޵�!R�k��Y]��+�,��ݪ̋�PLar�u]�^�s�E�N+��JY�Ƅ<
�Չ}�V��8 ѕ*��AH���*�uݍ�qV)�e6wH�յ�q)�dgJj�+�b����e�EU�jc���}%u���[8��U����4<n��Գ��mGd�)�AܝUR|wu�9��'q���=��L���a�u�5����^��z%�6�J�ʣ-��4�`��4���u91��e��f�yֺ��h�p�olVZD�I" �d�$ES|�<E`u=Se$/��~ʧ�.W�F��'w`Ǔ]�W�j.��pUk�c6;/Gs'���\C5iZ3�:�n���;sM�j�Z�*n��7���7��a:�UG���U�?������vT'�+�ʮHj���Z ^�ު
U`1v��㛹���> ᕓ��h�e�i]�=���+���`7aD��55;��{7*(PiL���k�_LU�(�Z/v7�[��W���y.\Ν�* n=��N޵�rܭ�n�}Kh��*�;r�7ӷ+kN�o����!)�w>"U��ǖ�5.;�S�	|���������;}n�(���t�e�oR�;/-�+klwo�=�#��܃��}QD�g|s�.��n�I�n�����8�ܻ��v�t!Qjfu^^�S��h�N��x8ď/���)jR�);�*��e������v���b$С��G;r�u�צV7a�d�C�va�94�.�J��Bܳ�eި2P=чG;��:�Y+f���(c̟�2]��K�)�v�ŧ��Kа%egh�Z��)ge��8��,����3vjݥ��#R3t(�6^�Z;���_ƞ�?6����A�s;U��t=149\�k����ƺr����οa��g���%�56AԤ������	���ƃ}V����65���S�@Tc׍�v�Ǐ<q�Ǐ�z�1�X�[I�u�2J�T��n8�<x��Ǐ�zN��.k�cͮ��ȝI��5
�����q�Ǐ=x��ס���UEUUP2THI�r��qEsr���3H� G�^�8�<x��Ǐ�ߛ�4�͊�n�h�1���nk����o������s����5ʍuw���7.U�iݹ�'�k�}�w���h�s\�wWu���.�#����;�(���W7$�n�"Jw/�[�r�r+���\�w[��rشh�(�������;Oq�H�a�;�G���r�����i�u�A�M��.�䡸��JT�z�0�곚�wa��}���y��o7��q��u���w�w������Y��m�О�w�T��ɫs�IK�{�y�Q����uQ�&�����=�A��=����Px���G'�Nj�Y/�9����5�=ܫ��gķ��x�`��6�Fץ��2d��ϖ��0.�/�xEY����0�y�`Is`����}?[1Ȫ���2�,V~���P��"OH��]f^z�lO����ۅ��$S�To��0I7lL���7��=�J��ɨ�W��iբ�����-o��6l�<��בS�lE�)4�O�Ь��0��+�%X����$wvN���w����rX�r���x��ʷ˟c�9f��4���\UGF-z�O۽���N�ɐ��	W�OJJ�|���_��X� �!�:P5'z:�/�,���y:"J�-�M��X���ơ/f�e/���5���Y���j���.c;8�^g9k�Y�R�C)�٣���w�%�r�.ʗ�긦[�U޽�0��[�#��b{���.�9�/&a�6tJ���v�*yZ�9��Ẋ���X��ΨV��İa��OVk�g8�J޼��{��xrD��1�c�o}����;�EdorNDyP\��ݰR�T��9�H��4v6�>N-�}-���a6�ԇK�Dj��rn�����>\�\�&�z��z��I���Ot�S;��4�ASkl5t09�Y���z��෇���Ǟu��	�;�pk[:$�����7My��}�,;#���b�EiL:q����\�$����1j+=����35+����Go�b��݁�kYr�x&a���q6�?���|�V~Hy��t�3_�}�f
z�g���mr���5�D@g�c�K�n)5��GGt7�w�����=�a}K�yu��&��1탕	��f���%V&��,n�<X�H����^t���!��>�%cy�;pmB��O7/<�u�8�e���f�Ӊ��,�ZB�Ȑs���>�9,�: ���h��P��P�,�60��M�L��2��{��y�KST$dq7B�U���X�9��̗���B�U|r �m:���\kT���QPe3�vØkW*�9�n6�j��q�ޤ.k<KOdB�#yԮ�{Ϩ�������g�7�<�%��Wx'&N�ӵV�f=a#G#:��{)+$_��xzɤk�l�Y�Q��(���yW�8���M;,kz����W�=�APY����Fl��u5�n��nꢩ�۟7�E!�LoWW~�~��-�i%)A��^�
�̦'�6SS=�Õ��1s�S!�G.�E�#�5�qT����to�=﷾�~�ޥ�GN�"˪�w�7�������R���S��p����d���Ӥr���f�\���F��C1���%�]"��M9��b�4��ǯy�Y��h��(�\�>�Y�������-�հr�YJ������;���"㫺�9�z$U�b��بy�~����.Y����;�y��!��6��Y"#y�m�����q>[y�ޣ6�U����GP��͖��W���y���J�F�ٕ�{Ӵ9�e{�uP����5~����1���mF��3�Z.YM�����2V⭹W��-e�ц��Ң3�7rlMp��u]^�ƹ k�Wž��$�����$Ǚ(-K�!��M�v8֊�LY&��Bi»ʫ��^Dޱ�Iy:�E������1��Us��N���3\���O���7��5�9e�V��ݲ\�f�M��B���8�=g5�g77��"|�t1��#e�`u|�R9^l�D�swY�+��x�c;�f��8n�=^Mя�p�7=`����d������ܭÉ��L���F�^���E��k����f�'�^�q6���y�������2BVF{�P��=L
�;�VDmmv�V&�¾��L�u��^��~{�ʋ�t�r��#��w�w�L����<�jg*�=�	�p�A!}]��ŷ�����"&n��+oe�À��Q�v����6c�<����~t�<W�;�#?l{��րA���BQ��*��4o=��T��lΞx5��>�YPI)0�S��ї[���E�J܅,u�8�P)��dȜ�;�G|Ei��q���J�<�J�^��t�7 k�W~���IOa�.lʛ�f���G���Ü�����	k��l�r��1�v�5Ӯa9Z��t��t���L�K]�����r��-)�[v���`9���=��2jL4�;x�l��e����r�H�S��׹���>> Z��q�xh�g�O#cأ����q���\pp�4�-��O�ae��"�6�gww�螳�Ta�Q�Ge���|=F�+���ӹ03꥜���[��u����1vP��Q9��UܹZ�0�6.��&M�T3�F{���(�o03�^6����Ώ0�aˤGb�fT��5/��f��X�
`��[�SCU�y��3�\��Ӳ:���ヱ��P*:.hL,~m���H�\���Pe�g����I�<$y�Ds���}kF�̲{�B���/-�R��>�$u`���;M9�l2�h��Qnٌ�3�E�:��E����dE��wo�~� ��゛�x���%N%7�t{=�rb)��M�?��B���*:��qVz$m����n��u����2ݻ��ι_g�)v��ܚ��.��2�U���E�l���y�%!����n�4��e�5�qۋ��jV�V�q�S��ز���WT3{�H]�%k�2�}��?��43"�����w/���ʼ��:��d;i�̺��B����f���ӅM}*��W��p�{|6]���1�ge羛�j�{bf�wvڮJ4�vY�A��ZA�ub��O�P�e�wS/2�Q$,R��{#O\�K��Z��M0��&lI�g�/�u�pm��-X�K#B����`�J��)��W[<M4���\TA���|�A:g<k�}1\�O��ts�U�L��������b���[k;�Ɩ|�z��>-�F]�Yf[v9O�*\P�ӊ���j�E��pl�ٙ���殖�'u�B]�-�����8��@�;M�v��&���1��`ˌ�e�	m�:�t�0��WC��{��W�
~���aTS�P*���kwY���^(�<�ݑ�q-����O\�k��HP�;h̒ݔ������KR&g�t����"��nK׫!s��=�>�R7#��d?�5�Z�x��+�6���`�u�?va�d}4.��5>.�3���!DQ՚�b��z[Яo���"E�8b7�*�`aR��֩�ӀY�	��J[c�"�&�����B�c۴rd�ﺙ�X�y�a,�t�E����N��byϥ ���%tKi5�{��Ők�x�������ʳ�f�1�Z4�������N�M��]3���rgd��u�A�{c��We'��&k0�"l~��~�0��߲=ϣ�d޹�l��twF᷽�y�ޓ�N�W��[��ȷdegr��³QiX�����bkj���N�Q�Nu�����f	X���c�^EuEz�׽l��b��<�9�pj�O��^=Otsb���,�2 ��T�LM�����BsMck�d܅��+=w��MF�;~|�W,����;2[��R;��؁�_ώ{
�^#�Q�
�����ˉs{Mt�]������}`��![�~����?���)g����<�9�W���1e�[g_��9T��%�P�`Vh��,�n׎@p������;os��?Cû��4�T森�϶�d�J Cz��U���xb�v���b��+D���������:��:�����x�t�׈[QÏ��k�����>��#@�t3i:�˖^�-�Sv��Ƅ�t�f-؋��n��.F�wc&���S�UI�y���Ou#�,�&��ń�d��*��*c,l���x�����!�J�7E۱%ދ�{�(^0j�C3�ދ|=�'��c��=�y���)�g�{֏u�SAJ�E�k��d�'��Z��>�c�U�BB~I��B�7Do�fHq|�P�S={�5����Ի^ .϶׸�3�~~5�������[�T��v_������wcXpj�M-ފ4!����ӗ"P�(oWF�(�/8�$w[����z���v��e=�"+��S3b��h�@oJ��`�0~�x�a��eo�	t��bD��ۥO��ݲ���I���9�%���$14g���8wU�#�V�'#N+�ge]l��"�w��6O;0w����<�ctƼ��;%���,�#��'{�<�µ%����zf׫��]�4��q�٬�I$@�m7&�ſh��`�.Ԅ�A����s�щ>g*���T� �S�����e\�nf�k�ww�j�7���FX�7�X�S�z���uxC�������y*д����}�t!�$Y�ύ��wMan>������m��Oy�2�{:�Z�[���}��Җu�N�
�3���.�ʣ^ȡ������K���P�V�ۗ�u.��d�j=�ǵ�a.$��-U���Mo��e�j��c�3���w���w5W��,�)��qQ,�:��+�b	�R��i����u�X]i%�K��Iy=]<��y�OsL�����plw�&���0#9��<2����Iޒ�JF�u�(RJ�̲��5h�������4�Ub�U���c�L���h6V��Y��Z^�!B��v��wGcr�nݗ��&(��h��H��m�(=+���x�*W���t�xҡ�#��{�����lP�ad���I}�Z�Wa�4���*���:�kIf�&�t���(6�a��z�T�3��P�㞻�%Qʋ�0�����o91ۏsl���,��`�f�vt�;�I��y�;��������cN6~���\3���bU�����!�\q������`�>����n������ɠ�3��3'��}�2bnN�c.�@_E��T3�`ۏ"�Ƭ�&�)�.T�r�S=�x��v̚��M�6ӈ���WF�}���
�a�*Ly�K�ȫ���J�y�;�����3J�εD�s�b�њc�#ǻ�+1f�^�Mh�u��@����>>oD����	�Q�N#P0��O9�����x�>���#��ۇEE��Ve�D�������ş�ֲo	��V�q#u)�H�Iu��������t��������q�^_55��g�م���S�.�Wy��Yg;��.��[��@�C_~�Ï���ED�5�A&�앞�0&d�l�|��G����cy�������^Oe�9�j��PF��!��m�5T@���k�p�n�5�EkyN(��}ו뛿CMX� ��M�!��n�����+����w����_��1���K�"����j��!j����nI����c�cײ�������D߹�Q�8�R�C,}�3\Ү����S�]���yr�-{��_*E[��je�lF#M�Im�s��F��g�̀`4T��7x,�F���3\�{��5�|pC��2�Ü�Im���zaW����2<�6�޼7��ᚬ�Lu�Zs�T�9���pRf@^�|�u��IECW۬�ɖ3V\�9]��7gs٧�jH�̛/�l��M-�:�E.�v�8٘3bܜ���*1��Z�6�qؼ۠�(˨X��W�_���֎5����J]6�iؑT՛&��k���7��hr��qJ��9!2�N���Th�":߲muLd��,��u%�c��xz����ncV�͊.��Q�k�6�lg\�.ȷt�t=���8�T�::2�B�1z��8����iw�m���u#�U,������zs���=[�U���O�K �/�-Ӻ���D����D��һ����	a>Y5�ׄh�Kdц��HW'K>M�V����]:����eLR7bsg�ucdj%}[B-k��*ۤ�>AGS�Uyn�B:��&�����Y���wwݫN<͛[�B0U�LM�-����[6�����o�������ø�'u�`��N[�Z�.�2Q�Q��_XSb�%e���a��J����'[�WK���3z�|{�VD,��i�C��o^5��ùie�Va�Y<V���;u�[�V�T\Ɵ6r��l�LZ���,�FZr��K��n�}�ɕ.���Q'w�@�#��j������=J�1�v�%w����L��V�V{;���opn�r�i�:����G)��Q �`�-���"�9��V�(n��	 ���H֪EYe��sc_m�Fh8�ٙR����8���]g���:[�eN�ں���q���j���Y^j�v^q���b���j��;�بn$�Ջ!O�2k#s���2f��������w7gq��w�˜čc��5<�R��ӘQFtqJ�򪘛&9��v���;x~�f��	�R�޸`�h�U+x��NgX��]7[�٤=L����ė<�ӷ���yIhs���sW'Ò��RGa����k����_N�>��t#T�̂���"��r�tb�k	cf����-Y��>�t�3���y�j�9����7A�UH%��y.Z]�g����p6�Ǘ�mWJ�̇D�ʍ��0�ۺ��p�F��$w��ek�oGF��$�����M��&JN�5>��j�酳]V�*�g3/J�c�n���uR�(0vI��7yKX��B�N<�d�ɗ�����j�`v˔#�gzq�7�s�ek�|u�&�Mg#;�U7���'x��n�:��!J=)[���fB��[.����51�s��"�j��nr���l�F�����E=)SI���'Vo;50�m�2^<�%bu��\�ܨ���W��e�]�u�x&�;'Y��o�&�>4�˨FF����22^���$Ҩm;R��|Q)|���|A%�ۗs�]ͼ�k��o޴uA)�n�8�۷n߳�oǯZz�ɯ9K��\�.mt��\Sd��1n��W�n�z��ݻv��o^�{�2�0K�t�.j��s&�ܭ卸�UP%JjB2��N��|q�nݻv���ׯ^��b�J�QMUS%QV5�s�͹�\9�A��IUI"��ׯ�;v�۷o]�z��#ڦ@�UUHU!P�UJ]v���"+��j�sr���/-�v�Wws��(��Q����6���H�ѮWwE�~+�y��t]M�+�˓W+�']r#c���ݷu�w[�s�Rs\�sQ˖�:��]���U���,�!]v�@E��û���y��n˝-ΑΗ:�@�����2�	�g0�5$û�Մ����Ȁ2jD�.F��P�*MA�Z	����. �0�Kb�	0^hح���<�0�R�es�6��n��p�;"�����.��U!����Hй3������m����+Q"�#q��*X%�#U��h&IJ2n2�A"�a�PB�i�L�H$ ���,�Q�q�(�1�-)��2FI8�.&
E�ATD + ������~?�w<V;���.o��{�a�m^�F#����"J0�88c���g��Qo­�ݏ����:�t��Ƨe�`5-b;C��Qs9�7h]s��;^����aID�[���n�]����:ހ�{;7��C����������͘Wⷽi%sSo�b�e-����l7u��1��玉6�˅�"\z���5���7��= �b�3Z^.w%�kF��K[��{�g#�d
�o��j��+�L��K��}��#��G�_^;�wn-��F��ہ��������-_8�7�<t5ۖ�`�yREc�m�X�����Aż�	�����&�5��{}A�^q5w��n�E缓}���@l�� �,!� ��X�2�y̝"�Zd3���t�2��>�!/PJ�׊:�3iM�L�e��[��{�5�
�]��r��*�"�]xAHW�zw���U~�Y�H�Ϸ85��W��������c�>��nmn��[�՛�U�t�#����|q���(��=��O�alʭ��u�5s��7WZ]��D_R}�3�IX�`z����y-���i^<��nV�s6�e��|||||@���'��k�Cx��v����+߆��$גR���Vv6�|��m��٘t�Ϋ~�V����Vh�=�[�K����I�5�ڪ\��6����w�uISl�]:���t���Nj��fC�0���l��8>�=��������c�:��v��[�ۀ��r�lDck�B��1U���{�]"�h��(q���}�,���fz�z����ĩ�R�Ubbv�:[zF���i�B���Am�]�:�RR~��@V������ ��S��b�X�a��/x^�5H�<ۦ{��j7��K+��j�r�u�vzϣ�e����f���#"�$\�mӻϫ2t_�>�Q��ύ�n�?����w��X��q�Kǟ��>Yg,�F��`�R�MZ�y9)���l��qOj��Ey�t~B��?���{��V��u�=��b&M��Ӻj�'�.#��wL)�Чո�1���/�uo+kϬ�ݙ=���^�-���1�H�2 ��-㹆�L�ZNN�Wj�n��3�L�[�
�R�dJkz5����#�1L�fn��}�����~o7�+w�I�-�;;�5���CwO�Og����n�it({�r;S����^/��*ϔ^Y���*�^ �>R�\Ӛ�kS��q's�U���9��� �{��ʫ�V�׷2�� ��4����ǥ��xڷ� �=���/t�އ����N�	?":�k�rO�\����5�2�CM�y�z��]N�:
�X� ;�H��z1���h�mj��+b�u߫4^�����yU�藋�g�3
2�)�s)q�54޾����&;����Eu�����Q�U^{�;��}��ɡcB�p�3�)�~�~M���6��
O{����,��|�(�f=�v����jQ����z(�M�<���^/(* wѳ�dV�@�TzW�>M���6͒���Ss�~�`�
���X�>��v��H�٧Q=Uv��Mk��T�a�}�Z6��<ި�Ѵ!��s���z���ߕQ�藵.ܷ7J����ס�O�@P�G�I)�3Ư�z^�_
l���:���Wh����q��:/D9�g5�H�K�M���ݕ7[J.�������~?���N�!�3*��λ/vW�&]�{����<�u׺�}�u�SX�u���F��=o۽i|�E	U�۲����Fo�X�v'�oU!3
g�顝�ڐ�J7xI��>�ԇ�?-�����hP��9���J�<2�{����~��O<k���4�q�w؞}z�!�+���$��c�.��w���dU�3Ov�b0/[@x7����H�N�<wǞ��������|U�]����y�p�8c�,��/4�����ft�$��n�	���M�:z�7�#��ys"�?�}i�P��f?:���]����Ϲ���.�r��A��o)H见�����F���EM=��p��v��0��WB�u�ǀƼ��l)��5!N(#�k�Ȅ�z٧����E�jw���Y�"�J��=�@�䊚{�n�rm��8�}�'�C5:<�b�ƥ%骦�9|��+v��ސ�X�O?Te��wb
.�8R^���k�F�Ա���l�F�x�	_)P3=:�|'��e� yF�(�5�Ui�h5r�K���ʻ%��̴3K�ʾ���eG��J`YgO�C�c�d�|k2g�����Y�y�����H^Z��x�ǫ����_.`���cv��g!�T�i�.�F9'�Еq)7�)*�&����zj�Y�*I���}�� +Zs!>�p�I���qVN�j�L�b��ݞ]����K�~��l5�p�DL�\h0�G��t�T�4��D�V͜�,�e�feYǓ>�ݑ�\�m��>���起�J��î�.e�sp`<���5�Y�Y��fs���N��(ϴ� ��G��P*�>�e9p����w��ݗ�K���TJ1"�s�'t����L��f[�C.c�Z��ǫ)S6p&$�z�#9ܶgwⶊ&��)���ݻhj��Cʈ��Mg�	��`���\�}Y5��;�d�f��Q�D>��3�{���sw���A��Ӎ�w~?���}�0�����.�12+9�!�nXt�̺�f���/UmyN�r����t�
�z0�5�׫5͈[��H��j��9F�"v_K/N�jް�0]�oe;u���̍�]mlYΧxf�x$l��/��O��d���v�wCG3S�o'���s7(�IEh��6��p���&]��*zs����}}�ٸ/dG�����y��9��6���0�^)�I�z&0��$��>��g;�+�\��ڨ]�U�w��o�
���5�|x���|�s��^x�M�N�8����X�9W|-�%�Nw?WS8h��m�@GH�p��i@&��Q֜�W,���P��p�2�yY�z�c{�1h��e_�ڵ��5Y����=�ojD?d9F�u�m���#&�&��!\��Y�W��:��I������W o��mn\���;5sDj�2*�Lf��� Q��a�G�H�A��qS���x�����Ït	K��=�>�9N��[_�>r���y[x]�7nx���E���9U$X�:�d:���2ُ�@ ��Q�ZM�[��
����U�Y�:���K�mг_'�T�s�Y$��Q�ng��Z�K����b��*L��=}�<WA;�˱��-�JUq��뉍���j�lQ2�m�{�7&B:׉���!v�d��x�P�Q�ߍb',�&����0�}��b��W��$MS��z����?V?���:�h�7��7��P(��W��R�>f��"�V��d��S��I٘u�:^j�̿y5U^��1��r��gk+�r���<�@`z�.������Wwy*��1�\r�2��i����*�Ǎ�H܂7�����eH}Ӽd�C�hkܻ�L+޾��~�1���m�h�5{��ڶ�,�1O���}�{����7Y����->� ��A`��>g�5Q���vɲ�vm�.pɩ�w�aU�(ѱ�}�4�8#��M�2ٌ��nK6�dv�E���-ᚃ��y��_ ⮺$n������Yi�:�n
��4Kg*�|y"�z�l�k�m���+'hn��VD��̪�O�h�s,wr�������g�w����>d�@����r�h�iޡ�������,Q�RI8�Tz�\����r`ճ�6��.����Kme�-���y������w�@�d�3ʨ���U�j�����:��33����S������8�n�L�<���"?r�}s���Y�J�V��x���x��y֜;EF�)��);��k7�&r�V��9�yU���V9��Vl�v��e�4�o%�w^��芫v�����D��������y����n���6�!=qn��g+�JLq�qt�)�vc_J]ȴ쾷n�n4������5� ��Q�t��Xg�q���Jvb�;�A=�[��ng`��	,�A���^�p��UŰu�TJ�c]#5�Y�3�'V��;٘�t�?�e�
�v�*�`�sZ����W��粹Y���ʣ��d�:���|��l��i�T�G�����T�8Q̭�7����P4�Y�����̀o��+U�����\���xR���ܒ0S�� �W;�.�d��V%tӳվ��p����� �T߭o�Z��_��;�,)���-�uK��W~�����7I�A��oeu���O�M��M��5'���"�8�D�����V�n�bƝ�'�-�eR���g@�h��]�U����T3;��p��M�g��,�i��W/�K�(�x���{:
;�z�YܬYN��*�-ʺ�<E>�� ��u�����Hx{w���dޜ�BK޺7�Jo`N�S�+N�Љ�J��+�tM�:_LgF�m=�7i�6���|�ߌc�0<�*���}��;7��}����@�����9˱i�osv˔6�]!�n�A���>#������/��`b��)�`|�G��c�z�߲�%��~���N:7��ܷ�L����x;������rw3���=�*�*M���G?o���<}��Tyo����Ю��Y�Jm�z�-�7H�$w{O���U�#f�=���EM9[O�
�"u����^��j��R޵��ȏR�b:�*��)X�*����c<�^ܫ4��7vK�����@[�+^�=������<����M�:��uG]���Β���<*]o���]B�}�(ųEC�մv\���/7{R��_��Z����[D�a8,��|wB�T�^���n0�8;�l�ԕ����w��߼O�h��/Y��?8�W��vc�S@����ݘ��.������k��8�`�Pv�nc&����p�|��֎���bU?YG���^�)�v��a���5���V�ɱ��D��2������d��]�L���H;���&R�=��=��&�;w��H�U���҇D-A���B!�خ��Π����y������f���-0LXq�Tj��ل�q[E�Nf,�B�&��m@�F��j{H�8c6SW���i{� r�wFSi���u�gI��p�U���D���&���DDw�z��c�hM  ���˄}}��3���,���0!�O���7�=j�`Wǽ͂8l��1����<+5���
�o^��8��3�Q��0y��bL��p6FC8A��o��s�ikz�B�ȍS��E)T���v3;���殌��~��b��)?Oa���J��+|8@�����N�ZB&W"�ߞ��k-�U�$�g9���ɚ��:Y�+�5C�̫&j�q
��
B����`���;Ͼ�x �h�59���`�K���s4�T��i�b�p��ۇ{�DY�ɛQ�V��g:�s{�F�d׌���z��
�q ��sS�F+4{�م�>�-�La5��́������I�p�v��C�죞��W�{�gk/N��%P/��?vB�yHbE_Tɭo�);7\��խ|r�L�T�����,�)�˾��H�{|�S�5�ۜ�]�^�9-huI��R�gC��p�ۨ��5�X�QZ�Cd�$���&�p������ST�R��^<wn�jtNb��j�5�T�3x�BG�����k��{�+�U����l��,HzUk���cꂪ%+�cCI���@����uG
uw��n�5�i{�u��gHe8�`��:�!6N�lа����|�9���m	d��K5��q�v��rT��ε���>�pmnt}�.q�w%�Ӥ7K��)E�Ƙ��5�*S���<�,�΄2ż��6��C����X���%G�Z+������{4�|�VGq�+)�͜��L�/^�E�ǎLg�}YJT�~��e�X�#%݋��,�lM�n�,XVwMm�(�)���sk\��ti�.�0��{5�x�>��.��3o�7b�]�+�y�'f�g^+wPp8��X���-�	S�;2�wPU�M�_f*7���!�[���`���h[�*��V�Yx2�Qy�t��}��R�06eq�[t#��2�����z�3��]�K�ˈ.k䒭�7]Yqss�q޼�u�.�2Y��5�K+=�P$���)5�˩�Hb�*@A!�T��mcάb���8j���bg@���� �1�
��07�������b{�LS]t50�%���`�f�_	��缄L��Z��K�xg(b�N��"�G��O3|d�H�`��ĳso�I�Q���UC�I���L<L�k�v�]��W3\�S٪N2<趞��^�&�a�O�72����2/"]��O-lhe����ׯ�I��}�mj�9s!��=ƞr7X����7ZuV��El��z���
Q}f��{����jU���٪�L�>Kr�|n��K.�lMP�y����m�?_���V-�<m�q�j��Y#�b鰱�^M7YT��{��lk-��Iq6X�9%�u��]�:r<µ���v+����᮵�ݏ2.b���Y��q#Ҹ�.W�V�MuTղ[�q�͓*K)���'+�T�8�7�k,��f�u�JQ��r
㻮��Y�>�����5ҥ���8�gF�Z<B�伶���!�ob�ܻ�R�3�4Y��{tvK��q�3�k+�����`�DV�m�s���ul�E�ƾ�b2�U��w���\���;��\8�8MHZ��s�N��V��̣��k�N㾚ܡÖ�+-ط�W;�-e�����t���6���|��Қ��A��WL� ��b$���Kpe���(���i Z�]���W�{	s��J����D	|���v�߭��[�}�v�۷o�o^�{��
��(�F�n����@(�N��IP�
�F�m����v�۷ׯ^�{ؑ��%5TJ�HU6���wu~wk��e��:D��sG-���ߛ�}o���v�۷ׯ^�z2,�IP�Uzd�r�� �w~w��W$�U*�QR2����t��׮ݻv�۷o\z�;;I;�I$��TֻiR��ە��N��wtӻu���;��nwqNu�]~���]��Lw-�u���wI���E��.뻘ȗ���䛻��v�rN����]:L+��^����# #��<n�4��{��8t�{�z��}m���wJt������:��뻸|]��E�w�r�yt��Q��7|��W��3�ݤ���z{���(�_=�dL�����w;�뛹�_>y]��E�Z5�CpJ[�j�I���5����
���%ͭ��>;��*Y�y|�}�>w�a��/�o��1��7�oGp2��}�#o��MqT�~*���Ս0�}��%�c�Q÷��`����/�RWθ�ד�W�n@ۨ³��<Op[lOI�n��)�N�b��r�S>\�j�&�>�SE[2=wMv��fY�kMnq�5;�~}�V��m�����s_B��N��M��s�'�DK3ߚ��g�m����x��A��3�����'���ܿ<Op�l��{�7J6�$m6{�m��
3tO�?VLUO>EJ���:c9�J~��q�zC>�.Ew�{�y�H�.��E�ខ��{:�2-��%b�U�7m-݌;�xߴ�Pc�D1>����J����s�>���]�-��Y�\�{7Ͱ=}gK��4�k8'�[���ε�	�%�N/c���h�yŵe^8�=�HH���{Y�.p��y�l�r��c�j���̹��N�>YS�i:��u<Vs6����h*ߦ_c����A��y��s���O�3�,�r,����}ٲ�9\���Z���]ۜf�8��э%ö&�Wc�;5eJs���4�xʶ���3���y��o7��u����:i��a:�~{�^n/©Փ��\�$o��*T)���v{����l�>C��7�m®��e�%/5=Qg��"b���\�������ov��ӌ��n����6�S�M���@��3�,�� �#�:e�w*����U�}W����L�B����U�y�/Bi�|[�h�"[J�Ù�_ss��xa����òm�&�^++�<j��J{.}���L�WA�ι�fo�t��\i�~�xWU�%׮J\�tƑ�5����ڌ�*��4tϘ��2�~[�sʼzW��3Mzxݝm�n��K�ɫƇmt��ipF��s��1}�Ft3��k�T������c�콪�/��н�-��\0Y��ޱ�*;��	�iG��q����>�̪�yU��+v|oxil1���W�b�_�x��^㔐���=V�������<ޏzM��-Z��y�c	~�g;'Ŀ�ߍ8rᳮmpX H|�p���	o�f{��=������Ε��Sr��I�ŖWwqnU�Uqm�c�|,T�y����6f��L�s37�ײ{��]y�|c�1�w��;3�|=�9cU����ݙԯN��T;�O}���8wb�j�;�_r���Y~&���]���;}�1荍Yue���Й`��q�+�^��Ǧ��f���GE��(fr���Hm����|��(�5��IWI oa_]Uܣu�kD\L�����{����,�]��}*��Y�3<��t�g[��x������r]�_�%��ݡ�s'U��ז
��y~�k����C=%15&n$_Kӧ�/h��/�J�z���������H�Ḥ\�*/a�X����j�6����������gșpp��/x)���Ƽ>��^��@t�4E�v��Yy��2+S'��y��c�l%�C�zyP�Rp��[���(��wez/C35C�[pۥ�r�²"�c�3�*JE�zq@k�Ɉ�҅�Q�̲�}x�E��j���&;�=\DOO���-\�+����pq�����W��םL�^K-��)�+�xĽʦ^�U ��<)��M/h��]
F܁�j;��%�8m�ѽ2�ٿ\C6�Me�j�F1ޣ��55Cc�}q�����6���ʅp�Ω�Կ�v�ugz6��||||||})�_���c��ܯ�$�Ny>������85���o˳��J��sln�\���e��=d�)yV�w��|���!��	ۂŐ6���<���s��D;��u�
��KQZ��>�Z�*�"ڼ����m�C�<9��c�B��ڤn��!���"
ٽ&��bi_�����]&�C<�>ef����Ռ}����n��Fߗ	���׏*��(�u%X�{"Zz)�ګo/p�iݞ��"�#�s����g�]�t�}Y���S�����h'H ���!�c��^9�fCtn���tm��T��ǹ��iu�_�{�\��Mѿ�N��c_��D���wF/
ˉ��잩LU�$k[�ا7G���;��~'���"�/�7=o>�D�{��ޓ.Xi5�`�6g8�6$l��W��v�c��;�nQ�${�S�ڭw{���E�&��Jߝ3Cݟ�����Y�$�Ş�"�X�Z��5�8|/��?<�5i�F�l�f	U���l�em���E�yCN���g2����w1���m�3�v���ʏ�9_m%��]��$z�a�;�ל���}_�y��͹� ���o�����UnЎ�uk�V���z��J:�x���Y���}�������z�0�g˽~�/a
� �oLݻ�i��%�N^�4o{{��niԁW�t�~�L,��Y���;�N�?qw5�-!�:�%)A�9W>�>�T.��ƪ�gh⚸�KK5�h}���F-�����+p^��>���QR�=�N�H��e&WB�!]���ɢ�F�IFw��R�uƃ��7�:���쎖l�M���I>Mj�C���C5T�=4�}&�2�Yި�Ɨ$���-��7Na���tn�x :��H���>������p8�B���u�>���|VǛ�����/]Ȟ������(���^K�}~E����y���~]�c�N�K�!�N�2{S�+����z׫N�2|�f��Z� o��oP!�Ň-�F�����t�a�:���5vf��3�c�IL����n�����==�g���O8������&r6��&���qo:��gD����rp+����{ULzR���T�B�u�U����.$I&�ۮ�m�%�6�57̫��������1��.o{���e��J�_Vq������9�lo�y�8.}��:Ű�x��Y�7Um���#�Ǧ��_'L{����j�y[B����jG��33�	!���B�ih���R4�5HY����C�h��;�s�M֢*z=��c��)�W]���䈎�/�z/������xff@Գhl[�CXP�v�ڇ��N��-& w���������?��|3WA'*�Ϋu=���`/�	@z�5ݍ	)��j�`�����U>���v�:���\ә��?�0e��UWc<��!mь�/xg�Z�熼U�*�yUx�����&����ڣvs�s����^��`��>����	���8M{�S�ά؆�^��]�3��ψv��M\�}*�'�^B]�JZ����-p�ؗד��^sT����.��6��DZ6��
��*dN8�".p�ILeu0�4��[��X�|�ݟQ�z �B	��{U���&�����̧0�{�Y��U���j��*<WǍdq��RU�^\���힣�����頗�������~?�B����9r_���M/��j�tN�v����t�i�{{�2���P{�����a�d#
�����*�2��e�����J�rr]��_��z���vzCp��*!�Ƨ�,�g1i��t���>�쁗�o;at���.�&W�3�����y�-,����u͛�C�/^��v�wUk��+v|n=�:���8#7��[XĻf%T�d ;0�a�s
�E�����++��R�N�N��7N���gvA/L��z5���ȓ�7�e�U���f�k��X2�;u[�5��m\!���z��P��G���
꣓����J�[B0��ѡm��C���z�U�E�6/�;9e�O<!���6���eo\��bW��m�h$��
�y~��o8B
�t���!s+Y�,z��U�5�$f���n��gâ�6��}b���1�
{�l7E]ͷ\Jr{Y��Ckoj��1�k\�O�j#n�l�����i����-
����&������v"��)�o�	[)������ԙ���t��r������º�h�!���Xfq�D���f35yy��o7���s�K��כ�p���P����~�}��-�v׼�;��N�zͥ�Hܱ��Dx�4�����T������%S�]m�s=8�;ͺ�mH1m뗯����~�����eaM��'~��գN����T�L�Ml�D���70��)�D��l\,�Q�[u�fS��۳oh��<W�kG]:�`��y�mwn@��5�q[Nt���Z�0�o��(���7�t��yx�à��]�W�jn�N�f��˅<���$�o��E�A���\孍S�Ϋ���\�{��Hpɇ#��wl��2/��� ��6��<q��I�w��[aN��̖q�`0��M�F)�P�wP�H���x�*+j6�v7>�ý%X�6�!����^e�n��*C��j0Զ���`B����ª�d��W���J�����y��vGI]<�́5�����;�*�P��>��v�n���Q"������z�l��n��wx����Q̙����"^�6wKΘ�Jj�tӮ���0��nbbY�����ʺ�/�?��=��f��x����2�ȯl���g�7�p�0K沾��B�����7�g��rF�ǻg�CV;:�����Cm
ˋ��o��ѓ����/���F�3źq�$��m�n�TRn�`����:+�xd��E�k�V��jz+0��A�{��qD杮|����ek�`aP@��UB6&%a3X�B����W[�Y�iY<`�ܠp�NSn�M����i�g��rV��,4���ۛ�E��9��$VGOwb���*����aTP��畡�n���Lp�m~�c�|�wR��z{f��~9��	��6�]3�{7;���kw�R� Q��m{_�)YV��M�{t�y�r��SU�i�w/g(�G_C�cbq-��r��Dּ�:��r+�:���������=�f���������Hԣ΂�;�d��w���Wh]܆\Z�8�
��h�9�]�����[_�ڊ6l&�y�:h�:�s��s�������꧌�f�o&��v�I�z�쭷m3W�R�{ѹ�;��x�=&��m�0��q��N؉��[��M���^irL|����T1��c6�8���y��L�#]�� �!=ߺ���H6��k��]���Yx+>���f��])Ĥ�h�e��`�oLANt�:.Κw_��E�^�啽�0��j��w
��GS8��/ ��3P�ݢ��ɲx�%Ov��q�;���kϦ�}�je�Uy�.#\�����H�e��uר�z��WPc�k��z�t�6����\�j��^_6lkۼ3>zzG �(6N�V-�Q��[�ٮ'�=���q�q�^���v�E���0�wf��9	����[�^%``WOzJ��τN�Z=n�����1d�ק����+LŪ�=WU�����fgX\)�� ��5xg��:"`٦�� �����'��_ľU#�( 
�����?��S_�A��AF��D�=���|�AQ 0��[Jʴ���ibͫ1�6�VV������[Ljj��Y�M[1���f՘����Vj2�M�j[l���Q��5U�ŕT���%�m��m++jdŕYX�,�fL�K5Y�&VҲզ,�kJ��ei�6�X�֘���X�U�c&�VjZ�m�ԙm�1��Ve��3j�U�2Y�R�Ֆ,�ib�m+*�������Ͷ����d��Ki
D���Y��56���l�gJ�V[f���Yb�l����ڲ��+5eeT�6�����YYm�,����Y����Y[,���X��+5��VVkee�����ef�Vj�f�U���[+5eel�Օ�YY����S�)5�����@J
�@|�
"�@b(�U�V[UJ�V�Y�� 0D�A�PU ��کY[U+6�R��T���J�V�YkU+6�W��(�@`*�@b)R�m���کYkU+5 �� H4
m��e��VZ�J�Z�Ym����R��U+*�J�[k��[�iY�Jʴ��Ҳ�+6�VmiYm�`)�R(���`)5YY��fڕ�����0��SZ��HU 0VmiY��f�+-iY�J�jVmk���iY[Jʬ����e��������D��!#O����y�{>���ADRH@�
�7����}#��~oӿ��O��_��o��g�?���D{����'�����AW���?w���QUD_8�V�������?H��O��s���_��������|�@+�=�	�����~�����J$��"*��P��JU�֥�if֓Z�f�M��KZY��U���KR�%�-5i+i��R�Zm�Zf�5�Zl��F*���$")�J�ZjV��-iSV�jmieZT��k5i�ږ�V����kM�6��kJ��֥���������-��֛SkF�E��ٵ�[im-ZkMY��*ƶmMYMk3[-�lU����lmcV5��*VƬ��b�YBE@ EQQ@$�� D ��V���%���I�Q����`	 )z?0����������V��cj��U���QJ>ÀW��>��� g���`�����A U��(?��A��C��{�z�������?��x~���p� ���Ɵ�ӧ�r* 
�x� ���~���  ���~C�B* 
�� ����A�����l#����7��G�a�,@g܇�~���� 
��m$��������? �`~��`>�'������W��?�~�� �*��}��hXK)?���4~ JO��S����|��D�} 
�'�$����?�(�?V�xx���3�O��
�����������?�������~�����d�Mg�M��f�A@��̟\���|�����(P���Di�*��@HEDRQi�UP����J*����"*	QT��RUDQ�H��if��kiVڙ��Tikh��[�ҕ6�VKM�0�-�[M�6�b́�kBa�e�U����l�)J�el[
X[cm53kehk2FY�����[Z��Z�H��i5�+L�fZ�´�4d͵ZJ�M��mj6�iZ�lY�l�l�Se�bҴ֔+M)�ȶ)��ٵ1lѶ�Vִ�Vը�4��  b�K�]ݶ�w;\�n�ݭ]���]-S���Xܻ��ѱ�7p3�5���ŷ5-.��M�McV[��wQٝv�eR�\�n��F۷5��:V�t�N�٣M4ɵ�[-��)*o   !"�
�*�l*���X�z��ȑ"FؑCu��U"�B�
��n���]�g9�Ww.�MU��;��v�v�n��Z���wv�\8�s��ŷGGf�Jnl��v��m�ԧ[���Z.jk[Me��lRͱV���W� w{�umR�l������Yl�-�۸��wN�i����*�nҚ�ܩ+����u��;m�em�7Y���w]ٗ����u�F�[v�i�6�-��i�m��h���&�mB��� �盶wq���ݝ��\�6�հ]ݍ�T-hm��먫Fͺ�Ʃ�wWu�ӭ�E�+����Gw1\Uv��m����eҨ���KVV�XJm�am^  sȋ�k8ɛ��u�,�v��wT��[��mU���.ũ�ų������\3X��n.�����]A��m��i[���sv�Lm���֡��6���� 6��WsIDݵ܅j�c���6�֕4�f�Gn��u���GR�΍���M���:ڮݶᅢ5DV�EK[�[�V0b����ڶ���5��2J[iU� �  ���  ���  ���  mp ���  c�: m�0� �u.  �X  	�r��э,֕kJ�����x  a�@�fF( �+ ( f��  	ˮ 
 ��  k��(�R��\ s����n  �魳U��#K-�)�me��  �  މ���� (6;n  ��@ .v8  .\   ��X(�Gwkr� ��֪�[D�ի[X�&�m�  ۼ �Z�� w� (s  � `R` �;�@8ƀ ��  ۝�  5���&d�J� ���$�����x�@ �JR�`  ����UP0@��)6UR  �J�eq8
@,B�E��抠�F�Q�ob%t����.��N�6/� ����}��g�|�ҭ�km��UU���kZ�߶�m[�j��j��Vֵ�[UT>�Ῐ�����RC�_��Vj��n���+�x�U��*������"S�����Po�]]���Kj
.Sx�7w�(5��Jن�S�T 7l�;�0�ģ{2�y��7)(#r���9Wd'F�4�M8U���&�K~	V���ov*2���$r���.���fڡkTF��5��Q��w)��Z��S���bq�\nm��%oP�r**��xq����w�����AGA�;�b찶�c2=Ƕ���=n��^�I��=u�:H�ܹOM]X���g�03ah�iA{EE;@ԔW
Fm�meGqeඳT
Q�Q�Y��*�.��M*���T���X���1*�m�{�M�Jyv�~1����;kK;���D�����A��-H�I%�Y�����Vp^%2�S(��ݪ-�*ы;�<�����_Qf�B�EJSp�5��r4u���,޻ԃEt��u�-�����p,J�nHu-z�6�G��â�Ӕ6ާ�Z� ԭ[9��|��Z�wI[������l�D�t�x�#q}i���֬��M�1�TkAJ�G�t(�z"��}�*��e���0P�q(�nչ,�N6��K����\���1(��� ��Hb�F�6�j.�R�6�0&1������)��L{��0�x2��Ti�U��a�вchwaV�5Q�@�9�Kk(�Z�iTr���:"�����wp�d
�FR�n[�֒�k5aY,�m���-�d��H��Fݽ�e�F5p�fظ��p�X�nJ�v5.]ս!��t���1M�
��ʷy٥��ni�����٢�SY�ˏtʑK��Գb�����wT6i���%F:c�e��)=C.�2X鍅iՁl�зmqF6K0��e�ŴU+��%��ѕ�L����w��כVB�Badֹ�
܊D7v�� ]��U�eB[�F�Z&�"-���2jY� 1E��&	q��,�;�0�w�¡�F�)M��C1�2E��fQJ��ͤ
x"�!��$,�cp\%PxB�w\LIEa�yW+�#kt����`���X��;����$���{VK ���
�Cj�Kyi�w�[�9���dN�u]�Z�BT�0]]-u*�{�+����R�-�13��t�ڂ����۹���Qh�e�\�TlE�飃qU�z�ZW5DJz%��A�2�b���TW
x^TZ�F�+NMõXLONc�%m'Hʂ�Ւ'�fm����z�X&�:��6�v^���}6���XU�B����C���vе�<x�ժ�u.���Qv��+o/F;��VM����:]1�^;��b1�1D�f�[���-�W����ƒR6T��hf�	�� ��j��l���L;�Ǻ~�0k&#L21�r8 p��5��,,�]6�����v��*��K1c��ۋh4(����q��L�
/t�U���Y.�>�}{�-��VS ����]��`t0���_�LMF�V�Dn�.��jʹ�̆���nQ:��{�cqV^I�Z�X)��B�m�;;SVA.��Ũʗ�cAI��J�V4�ݎ�haI�amcR�q��Im�����Km�Oe[���ݺ��ټ�)�1VҤ��e�h�e�kX��J�浅�WV/v�[J��b�Q//0�Qb��i���K;[f��.��kI`��uQ`��\�0淸���w+H�c�Ҳ���3\�w��#��Jh��$�fe��^X�e̕��<�yB`�������"F�N��n�*����X^˺ҫ^��ax�f#x��db9��5�WKh��͌����:9ݶ�zm9CD�y�.]�{j=����LE�������
�V��-�(�y�۫�\��ٻxR�"]�D[��iՑH��X��H��;bu$ `.�fU��kJ�0�Ԭ�N�2�
�t��oB�L��+6��qݟ�[�q`�j�Թ[LJ�{��q�8�:ܗYF�f��&u�3�/���R5h�a�FT,g+v���P�V���L���!��I
�y�Z!뷴�07"!��f�cH�]��v,�,z4���:x�[Lk�mն/��
��w3!�c��EV��x��:ZV\n�%���M�v��ik�ld�u��%�@C�&R[��m��XP�1jmU�ڧQ�׵��h^h���YN��C:�"�y��n�p^ޖmX0QX���I�� �xj�����S&7H
��o5R*�е�U��I��
X��.�vF*�Y��I�����Kv�I�/��(Vڤ��z��Z��E�0ևa#(�d{$�G��]�Pa:8eZ��Z^�(�N�k�xP���	ж7+t��4Z�·a�p���|[�!��E�i
���6B#t�n�� R���6�;F�D[��Po�EַQ��"�[�v�ݼ��Y�ڼ� q0�3�����3^��� w`�́"�M�jY���a,+��GlV��,*m��LLO7m��KJ��[�b�R�^�jSh�԰}��t^�j���B�x�m�u� 2M�Z�ZK%��h��C��\*,,�k^�b�8M��F��&*B�*|X���x�csO+X  ��%�bѺf���IF���Z[��
�$]hy6�jV�Ge�ݒE��h`S4��Ƕ�ͬkq։3�]��x�nŗKK��_4u�b������F�ǌ;�j7/i(���d����:/]♢,A�2b�6�Y�����9o��X�;�w6��0�X�*j��A��[��`�[�JT�7.ѽ6�P�{e��"6}�b7�6���3\�����{�$����E�#T�����e��.*M%��b��g���W�w":m!�r�ON��.Fh�5��l��j'�V�K����8����_,���K*�P6-&��{f9���t��#7�QV¬��b��=v"f�扱J���6ٺ��eXe��У��e�wnvak1fE�n��i|��ǋh��e��z���5��[�W�TNa0F[u�Ȝ����J� 1(A5*;w�\/\AQ��!��=�V1��ԱY $���]�ٖN,��M��b�a2���O౩m�ס�9F�bTK�q*���ܬ'!&@��Vt�/iS�,�U��f���٢��j:���CU��EK�f�Y���6$�͈����E����)
KwBiǊJӬwk	�q�EGx�h�l*U�T�%�Yy����I�Y	�,=��P�r�a����WLl:wE�,��y[w1J����u�kUI��.G9z��ti�G%��+4՜j��)�U ���wgU��;l�]���Ck!nQ�--Gqb�Pǡ|��=�(̰hD��ʳ�*�Ji,��͸D�E�R�]m���c.�[@�Y[�Q\�ùp�ĩ"����B�r0�HVV\"�;=����u�Mc$e�w�n4E�#U$�f�Z�ǫX;*b��)SÅ��Z�<�k,ڣO*H>�I���gcP��z��y+�J��W���<�HfTObkr:4��=�� `�ٍ��,�70d�Ņ���
�w��(������8Gj�Vf%�[�����r�bYt�˵�AR�G�`Ǖ�
��&U�n������ �hԡ���2�7튊C`d@���,�sB�0�l
YOh#5l����6�d�1�l�)4\߬��xm8�Qq齅c�Ap�j�p�cf�yC>f�A�)�7n��ƹ�i
�GF)�v���G+�ɰ3�����q�W�iau�Y���sZkrL 37ɡ�RZ�[���l�2m�)�u�,�ͣ����*��ݎ�h�h-U�^D����Ʊ�C�՗��A#1�0��T�Ӫ��1�R�]:�b�+ �V̽�vvLv���)��5#DA�]2e4�aF�ش�[9����(�SvE;�E
˱�����kY,��@�U����g���)nн��N�yj��6�$-�D0[�Rhda���¹�nl;t�%�Hڐ�+L51�����p��ʦ�"F�`���-ɹ��)�Ԋ9*��.���ibb�F��y#����Kn�M�Ӱ�q�LB*oFJ�$�bE�1]]	YekX.|�2jEp��T�XݥET�R�R���Rְ�q\�%!D�1�XU����B����)�乥S�K�lL�B�]��j�`���:���iۥ�j^�0����%���Px)�i�Xp��AG�@�l�e�bڵ��{v�BUۻ�)��0N�͍wY�T�Gd�m8ٰCڴL1V+7�k�ц�%��a��toω�&%�� ̏(���)e�E��,,��A��Gbp+Vo��')�h�qu;���B��y�6�*�f�Ss.'g�śN�_c$�X�t#���j�4۸v�mY��y$c-#)�?`�r�;Z��*�`�p�IU�T	y%m6ޓ61"j��t4�n�/�E����+��Gm����wY[�Z�Q8V��md�*�f��Voh	K1I5�r�S;�-O�}����n�cR�X�1�bCO�%�\�-L n����e�����%���lk���2/�4�Vb�f�hn����.dd�B\b��z�'tmm�U���#����w��!.;����)Jh��-�)LnV��ڻ�&�B۬x��+5<��n��pj�b6f�5P]���L��ݝ�@7D�ȥ<0���GF�&7x^�j�,TY��A��ët�<��V�;*�q�3���;��f�q���d+0Y-�2f�
��[�մ�a�!t!�y�MИjM��l�M��W���Ha8S�W�/ J�r�՜ӻX��6Jjm�P��ak*�l�#)Ċ$��I�:����d��F��߳J6��2,��v�t�2(t���B�� !��t/"��&�@�R���U&�l���&��ff��u#���Z���Z)��7.�#-dA`�A����j*m�!WA<�Z�5(5މthi.�͑O*���
ޘ>D���Q1W�[qPәv���5.�/$G./����SI�U���4�ǵ��Xn��5ʚL
�*����s�U�,S��Cl��@R^��aE[���w^V��oi�c��0̨cYd���� ���8%�w�B"�-={Y2;��ig(�e(�!���nnZ)��*�0]�� 0��P\��{H4�r�dA�,�ɹ�M�ȩ�j򓅝n�{�Њ���ʹ�S�K�����jle	�
Z����KQ���ǻdS��b��3\Waå7����fҋ%�5.��H�@��l�;<)�[��KAK �K�>�+i p����R�x֛�5
��Ez��ڒ�2�����h��H�i��f�@c��h�CL��#eJs7�=.B�\T��x6��SV���, &2�ݚF�ʅl7P��j�UWV�ͺxn1�@���ȪXN����j�Y�K�?fl��̬�D͗m�� Uؚ+)�5�1�H[۱.���b�2�"�R���zպ9�H��f|Zf*��KԱ���ϲ�x2TA���9�J�(�Ӓ�_�8݃L�A��#q��kw n�K� 4!!�0!����1�,������z���m4n|���H0�2ӘhCv�`�ţ��wW�K	�
�1V�,�5o\��X̺=�2*�ޮ��9M3����i\�-k�E�N�@�L6����l�T̫�b&홉 ^S�B&i��ᬢЬ�fh���n*�ա���kf�T���t�ݯ�Uu�i3K�����h��"�n�R���Č����ajQ�DWx���io&��a׻W���;�p���<y�F�{�̷�V�QJ��īm���f�ս{xZ{F�Qb�V�wdիn��HV�����	uk�J[����m��L0��[Cbu5���z0:u-�77�څ�9�[t��eEY������Y�YR�z�i�%A(QO[.V�S�-���nC/3�s�vUK�����mҙ�P*֧CX��"�C(b�˴�4�K��j*F�X�gFn��Id*;B��ax�T��kvƬ���h5g�av1�Ј�O+6���Ӯ��
k�o��
��9���'Pf�B�����匢�n��N�W�� �j��7��n��+-���u��n�h�.�%AEc�����T���؛*X�zu�`�S�QYw+Ix��j�Reg�jԭ�]-Zw�i̴��%�m@#�d�3�	��.U�*,C��8�w�`��C.����H㥎P�ܡ���3˧f;zs$mV�T����D�6�{�A<Q���q�(�����RҨ�,�ܱ��+�lj�'��+��n�6��6�7Jb[F���a�M7x"׻56�E1�LT�!yZ��͜pT��ڗ-�����%b��7CZ�'�ڗ��ȥ#V�-F�(#b�^Vn��/	�R͉Ԑ\�����[�5i�L� �i�n�&K�5f�JںV
���V+�YM{*KH!�Zf�U{����I�&*a��ƀ�Y�{�ܨ��S��A0�x�oVR��8�$ܴM��*aӸBGi��L�7W�eM,��H�P[�$�M+x���+^�V�Z^���^�02H6)�R�r�U��ҤS�y��m\iGQZ�`R�{06�y��a���{��>�4bcrQ5�5�����ٺZ���2T2���J�t��,�J��I�f�<6��3��O�YV����sQ�K�t>#��(�����إ&���Ռ��y��CDB*+�5�=�ٴ�ކ��|��ULj�T�e�s`�ʰ�hTf�1B��UX��%4���[m�a!�aN�~�7Xm]Q�wW�k�M�'���!�jlƙrp[�Mø���դuuj��H�c�0��t���N��A\���$�-�.�>U׵���U��]H���s��;6�x�l)b6y������l;;�h��Lb��/��HTց��j��/�Q�M�:.�Ww7r��(�ŗ*�Ң`��0k��%x�\�*N�Y��Q���gN��a�Kv�˥ɮ�����Q�Gb��WX ����豠�Z�6�W iJ�'-�]���yS.�aQ���e��](䖒l�
�;��`;�W����+gV��*8�a�.���,�ԻF�Ԕ�ӂ�0iWZ�)���ۅV�ޥ�+}���5��"$.����i�������{H"���I5�����h��E�2ۂ�Sm�F�)���`������֠�7Ş��i��j���p2�=ά��
��\Į���l�ecz5nQ���h�K������`�}|�M�j�A����l��w6Y�wx�+�80���$8��y�S굶�d���K/'3iśp�[�2�����w��㶊���wc�3��t٩J�f��-[�@*��o(^�᭍߯tͮ�f�T6�uv�g3��l��|1V<�M �z"����gsz�<ے�塤̡{�s�}m��p�u�#�<nb���jaŘ���9
鏛#7[��A�`�/E���n�Q*n��.`+T?e�+z���j]�,�W	����ڬ#u5M�BHo�v�S&m;��r��.�Y��=r�[t�C왲5��$��@Z���«{���kw��$�)�|4,�.Z#��V���O	��~�S0��z�i68v���'e�]�lUŹ/�f�Y�X8���;�Za���W=��K��p�48a�F��J ��F+{�jnfk-���.�\խ¯�owg#������<�u��\�������R�����xV� e�;���3w���ӊ�z�'�ZL�m8ka�]��������#)��Bvv�.Z���.;�U�=�(�_!�̅|u����)X7Z����i� �=�|�y,����V ��͎�βbʬ���hn���n�Q��XA���z�^�*�@H���Q�'�l��çN�Xܢ*����]	��Nw����OP��O��H�`��ZA��+�D@�Z��-z�&NBF�{�W)Ұ��x�p�N}���J��isg��iDeꥑ��幺�u	���SOg,�,�b�9L�sV�|�<h[(LXl]�Zȭ�oPұO�4�X%�źt���	aG�wt��e�sGDzC\�<�R�Wj΋)v-��󢈔q�7��������;&;�5t��
p�YV����؎CB�g�a�'ǎ��G(A�59�*��j�7]E*H�lr:W�s��C���րq�F٫�����OZ�}.��Σ�{�wV.�V�m����\��u���U��<�|�miW\hªP�{�����E���@�詊�4҆ �9 ���8�fʵ��J,z�s����}��[6�y�I#*%�B	ٰ���k�1R���gX���h_RՈ����2}��A��ޖ;�4���M�s8i:�n�Һ��Jt�^o'3��.�UL1n��7��֙�R�%c��,V\���ޥ�kR��2�\�x�y|T���zȼ�>S�ɠ�����m=G;�흡������IF��2���s](w'I�uH��b�S�-,�I�Ҩj�qI�/���`�i������\��6�-]�E1d�@s��q�\�]��/����������I�I�������ݏ���;;��L[�z��9�	�����:V��.�U �z�p
a�|�:��e�-ٴ�e�K�H/��U(Z8 ��
4e\���p�YB�<��^�t����T�xY�i�p��R*,�u;�����"bt)M��y��M�X��uuo[y2�Hk��ދu
������`b!�B��ر�r�g�@p�M���x76ŽT@�Q'���Y�N�9���W�K�~]��Ɠ#�C\)i�
Uԕ]�1R��/��7&���y���>��]�c830+'�Sgu8�5�F �����r�t�ju=es����������J�;<�!�m_W]j�,͙��m]����N�,�rgr�i��צ��m�OjWHoQ58���d%m�b����|�I�!�*��՗X�����b�M�"7R;Mc�0�����F�U�V�\���Ի�<��-O=6�I���ݺ�ne���#��̒�B�_n(��h#:]�M�y�4�ﺞeҼ��T��Z��,�r��7���1&ƚP ��zgG+zZB�T���u�
��^�	y(؉��g]ʹz���m]Vv�p�6я*���ǁ:��x.��N=�N�xʠ��O���缃�,���&�����u�+2 6qU�/�U���.T��k3��q	C-U+�s���[Dɦ9���ݨ�]��ϖ5R�[���xn8%U���x��%X�Y3�[	y�s��ӹ�a?n��&fj�w"NB+0:G	&���#CI��
|�X˯�8E�W7{&,��{"4�m^�N*Ah�(���QY�+����:oq�Lt��:��K�:�f2�oi���sZ��(�@՚U��'m�8����	����֢5˹, ^TU�uʧ,���v�^=T�M83u�n|s@�k��̊:��7.s(I3Fک���^�U�KZ�W����	-�l9��v*�M.�
�iWL�b5�-�6T!b�ڢ.�x��dо�@�D�4�XRn�ө1�u��hM�(������y G(�h�4��o���@�^bt���I3w4v�^��#i��x\ckw��9E`�R�@�txZ�3�jA]�1���+��;�Q�B��A�T>����vr�ӑ��\�M���')@��>7׽�{&c��{ҩ���Ղ#�eӥ�����:�\Qr���XM��V#����>[�j�

Y�����8/�"��v�
޷�g�u�Җjn���YE���4���%�7���v�*�',f�ڷ2�+��z������ṟC�-ZU���U�Y�� �)ZW���7mu�+;OP̻QӸ1�(;���&rܜ)_d��:�(jcܫ��
P\%�B�c8�f�2вôtc�n�����&kM�wu�t�5��CP���b����k�^S��W8F����$��@҄��m�bx�߻����a5ͫ#[�z��b�j��%2Crv����m���dT���Rݐ�t+�Q��b��;
t�1������mk�Ѩ�!�n�ݒڠ��t��w�o}��fK@h�nv��r�^!]��}�{��t���p�c#�����ƍޕ�-P��33��L�8,� ߹Z�VKPl�U�FnbY$x&��1 �s9MBW\u�,��{z
1�:�^4�W|7�u�z�S���:K�_!�����5��ױ�:��t{[��=dg_>�;l���=�e"��SF¢9*g�8`�Cϩ�6۲�kF隊wr�ۻv�)�[.��s�r��1�fcC���5J�}&C��'�i�U�^��nU�]orU�_�r�d�'�|���dN̢�c���#��4M`�0�`#h��3-!���5��h,�^f���g9ݚ�j���ᣎ6m�E�h:����*a$i[����v��:V���ͮ��RthJ3�.d�Qx^-@9r욖� ��t�h�!}���u�8H�(tE��$���n�0keZcw@�7"�(q��LGgo8�e�c�>��9k%�k1h���Ҳ�@�Q<�bM���*:�߻p�U��HG�̇��]tAgMٖ���jX�����s,�KAlp�s�>��B�p)U�+(9�C�f��^���m���|R���ɜ��6���eH0l�Hw�'_h�wzUs��GS}]�p�{v��us����dHk�{-;�i�s��r/�9|7�%�3En�؝�S왝��;��p*�s��!C+X�pl�,m��t�B��Ly� �R�S���]���X��G&{]�ܼ7wE�l˭�]RI�e;��&�;8o}�X0n����;NC�>�g�C��r3���v�B�v1yq��c0[��pd;�ܑ'V;�Iv<w���и���C/�/��Wb�7lݍ�������������l����ZowZ�]b%�J<���i�76�W���v��6^�Uyz�W:��e�17�J�
\�˛vo�t�R//��)V-'{9Y��F���ᢣp�.[ȋӲ[�bge������m�[�y�ܐ]��'ʳ��S�Gֺ3Cc�i+,(xi���>=&訨e���Pg�`�î�A�툯b��Zd�R�1³�K%*"�]�d�@�X��{W]B�aW�ʊ# r�>����7i��h�޻�x�t���Gwk�ݡ��$B;5H�seCN��H53<N^���U�r��(��p�:�O���_'��q��]��j�!r�д��9��ZkNNQbֶ��s��J$Ѱ��k���刪�8h}M���l�{O+����4$�V���\�^m�u9��eaa��[�j[�-
#^v�{�2�Z�&P�M��@ہ�{[.���^WKv�Br ��A�c�Wc��T�l���wE%r���A����p�,�\'�ՋuG��B�Ke-�BwV�Oi�}�Z��}w`��ұ�$����&N��Q�D���٣���܊�*ޭ9
�������]�5Pl�ٖk�U,4
9M��:-��J(�.R�w�n����b��m:
tŮ��z��b�\�	�4}�}��bTe�����j��z�\ټYѺ�uL1HW��]Q:�о"�������'�]�]�4$��ض��{t���Z�X��Oj�;�Ry�zPݻ�;�	������eyp��%�:�G���;zk��]�R�]�.:��&33�F��4M$S֧b���S2�a�G�F]qio�Ev.�:eZ/�l�C��!�z�d�i�G/09��{W+Gq��"����ݡW$�E��L����̷��L�[gN����
��u�W�rS����B�������Z,[�!��o(N�,͆�a�ΙN�k
t�B�7��s{�� �M�Y����J@#����Sv��.�K�b���;,t�aeKYt�]g����DQZ�3�/R2�Y��[[[� 4Q�e�Yę���mPK#���
T9��NX��+[i�$�x�\*�� �˗ �����ۺ�� ��=(��2M����%�	���/z�;%vVeC`v=�k;�h�Kr��jmN�S���-���b�Sް�Fy=��P��Ô+��&:r����,,%ݕ�eo.ֹ�g�{ȓ�y��3sh�.p�^�[�Y���$�\p
U�ظ.��E/�&7��OZ$���h�0��z��y������Ew��1we�L��:�nn&�'n�RBj�4*j��l��3��Fw9���6��x�T�eK:��E�.�wJt�jC�o�<�'�-e�D��]�,�-��vĬ쌤��}o�k�]�GV����ʪ��U!�,�&[�ÿ�f>�Թ�66�m��fQN�L#�#�u���7%7U�!3ع[���wT�Fb�E8Q��Q9LY��t���Ӻr�6:nA�{�b��.t��Pg/��ϋ���:�GkAh3d�R�>sp����D��
]�z`��-�'p���Oaջ���Y]x�]IyxM̮e��K�hk �Q]���&Ǝ�NڼZ�NA�T����s>:M:02���#.�V�٦�R�*�g���)������z�����N\���xT�Zoqr���3u���亘���6�Xb��,B$3�ݷ�+����r����V�c��GM��L�9�3l�Qf��n]��V��b��v,=���Ӄ��4p�*Q���+���qd-0���ݕ8�����Z�����lv���YJ�-��3�Ϻ�-�@�J t���E�C��qpa�:w�̗��^zruh��[N�\����J����]���gJ��^)��V��T�q��;4��G�����d��83׼�S]����:����R+�yu,��z�͠!�P��wA��v���%#ڕ �__AI}saA�4���-\L�;��܊��=��wRN�f#��(���;���q\ͩC�}Żtk&�<�&�B�A�:����()�P&R͉���ns���zP�᫄Q����|l:���Ȝ���]�>�K��N'(R�	���rr`�BZ��D���+�fc5��2���e�|#�J�=�I|�N7�^oD��uQ�Ԏ�>��mi�5We@���`�G�u�T�-71^��[v��ֺ�ݮ��d�-��x]�M�`0���x��#([MM��9�:��ɰv���-}�:�`y���Λ�کX2�����Q�n��9�'a@�4��t����G`ŵٚ7S�e�X�jg���fVn��wp�\�6�m3i�Jm�f\�c��oec1�rX�u����ͅ��>��x�|V�r�㋋C�_S��pkHW<�FgC@�+}��B4����t=�''s��*��^���\$^Z��r>v��i��`x�TrY�x&�Ң�c޶��:��.�V����K���d�"�m옶�N�$���T:��g��OGy�R��*ܡ}��L�t�сw�'��+���(��X��w�V%�(s�z�H F�n��?��Z�8Q��x�z:�0�>�.9ܸ:�r���׺D��^Q�M(y���S���w%gD]�^�݄�0�f���0c�Дå������;��-Q��)j%��m��#6k��.�4��od�	�^�+P��\�h��:r%v$+���38��e�m^9*sɚl#�,�ڜ�R��c���]�-���䨔�GuI�ޓ��   }����������s�#R�x�R��z��
�H�'��KT��:�� Û�x����wm�0�I�'v7���k�e�"��m^�P��?<��E�cdBN�z:�9��VS4�c���rk��\�
�;Q��<(�i�/�,ѷ�y��B�G]���u7�I�4d	ҟ<oovJ`��r�����E���Z�(v-wC)��unGW�s��:����L,ÍaQ�O!�sw W�l�L�w���ɶ��X-)�}	8��x6|��Ǜ�"G^�r�]8�y3���s����	��+;���	�w�r�O�i��M�#�Ì�����hۜۙ�����v��f��d���|E@h���&���h��_C+`U�����y՛n�S���I�2��&.Ɣ������31%>i������JԬ���~�ء����΁p;�<t�S2�LA]�]ٕ�en��tl�ۺg�m�S����ۂ��L ��n;����v���e�{ӫ�ꎬVg=z0q�nޢu5�y�F�Cͣ�M�f�u|2-�X�X)��{���se,�[����sQ#��_�]k�?Z�e:�8��ǘ�J`ց]{���jΦ^(��Sr�$���D�IB�s��x�.�=Y��ުu۶�]9A�*�͈m�6��Z��k�2��S\o!T�^���}�sK��i��ͺ��-Ylp������B����$�i�M
�ݼ���w|�N7V�\����� *>����Sn���f��oz.7�Յb��#3J�dsf���7�P���"��ܺ�xI:�ڵ��L!��5�b�����T����없�Wh�i��Mŷ8���c����#�.�qj
=+1�I�C����S��8�4���{�G��Z�^CA̧w��lp\!�Hl�D�m}�A�s�J=�'"̑��R�7��.��7 )-��̬�Z�̶��C`D�:�v��i�����0�1>��FR�Ι�[��C�IW��ժ*�s�[v����=��bl�]�L}6k�[ҭ�T.�)�A#��,;���WM�Ӛ𲔣�T-�*8�]i%/[��!̣%����%���ҝ��S��⏝`!͗�w*p��:=n'��s�j���[p�G5��f�Q�(�wd��u��ǰ���`��;짝��#�w�(�ӓ����]ZUZ�vm�Ya	Gq�]�M�.^h�]����zI�N��d�Q�� ��J���S{���&�*�UM-l6[�(\i L�GL:i���DdMm�<�/�7������;fs���*�n�'xҁ=+�3��=�JIoh�@�����2�k��sZFW0)\�-Eic�,XT1���
8X��q��&�1Uo[�շOxhZ�+2%� qo<�B��(��*](�u��e��tN�t��+���s���-��'Z�L�2믗KFʗ���<���9K��N��2�dR�YBˋ�̘���s����+U�y�;��mQ
�����m�o����ۙ�cK�f1�e���d�G��0t)���xl�lSr�O��)�������ni\���Ya⚼r����lӧa?t���/KV��X/v��BqD^]ɢ�<�x�trf*K��[���r�Mv��(<Y4 X�B�^��Z��3��5�Q;Z�gو\�����֓K"[��2���=���w�9�F��]9 ��PW(�r����d��$��u���O�h�G0�B���&����4��eb5(iz0@�a�*2ݻ���8*�!r�(9��a]y�� ��6(n�Qx8�����x�'�S�o2���ҦZ� �G�Jx1�×ϭ�i���둬,�LXp+;5}�6�I:�n���F�v=�˭a�t�&V��Rg190t��c�2�}�WiB��`��M��t	+���f>=H27T��#4���}��������A���r��C*K	Syo`u7�D��u�yY�J�4U[�[���;�kJ�db�}���m:|�R�#��3IeY�ؗ3q�h��9zB@�Dar<�v�V����KY�n�Z	Bi���.� N��+���v᫭k�cF�@.�
?#���*¬!H��tv.u�:x����ų^�#��ۥk�ܔ�}`�ԉ&�ɼ�Ba
�'⣺v�V?��pv���wi�EC�o)=�ƣ/��R�(���Z�h�#&���e=gK)�zޚ�3mv��(
0T3~c�p,)�\:�ر�:kM=�Yl=t���aǩ��x�E�V��j�K�y��cw ��
�b��.����`[l�w���s�pt���Y�:�r�sU�(:	��e�2tck1����5`�����t��+�pu���@�(S�8s������.�Cs!�+�bw��x{L�,�� դ���I��ޛ�%�9�m�1�+m!Y�Z(�w�Mŗ�N��J�̹�{�ee�y�Q廾V�!�U���n:J����V�[.�R��gaã�)]���D�'=2���ɐ�W]��>y�4�Vu��kClf��Yb�����$����HF�Ne5��܂�/�ćf�Ν��a�aA�7V��ݏ2�7����>�ڕ��S������r�)�[ut=���wN֗� '�B����Ֆ�ΙT�U��A���ɠټ1�]@H��ü���γ*�m
VcUe̬*�vFT�8j��P�gL諻���eX֏ n�fk*)�t^�e
�;FN��R�����}�J��L+%�9:�W��mH��VHI8��t(*�P��)������P���)����Bxnm&�.�gY�n�b��A�q9;K֎))-���
���b�]W�/Ѫ�Ӌ�T}�U�<!\&��}+\b�)ě���#�`'����h���^��M��n
�Q�8�XHfP���˲&+�ط&������˝	/�v��B���\$@�/Vk�`��vu%��Ι�����%��n�☪Mu��� �*�����"�9Ϡ(L2þ��H앱o-W��&�|�O���V���Nۈ�W�欵�,�sz�M�|�p({���mZ�j]]�v#(u�������cYw:��Uוme�3[�����K[Y�"]S%*T�D�Ӂ������n��;�|�`u��@��mE{u��^�nj;i����h�����.�s,�g������=���9d�T�*2�V�f��yG7���=�X��f��gd9.����00�.����G/��m7��վ}�F�wPb^n�Y�bK�,��6�Z5�>܍�2�u*4�J��B���[op��+��m��S�k���urb�Ŝ!�����y;;�\a�T�
�%���Q�8']N�����Nw�]-�0��WL�|8Cۉ��qS
����������P]bm��fE��[�C�p���Q��-���e+Hd!q�Q��k���n`.��k��+�ӛ�ۀ��/�k����p�ER�������^eњ�OtR�[��G`��I�fb�����B���C+W�k^UƔh2N�7�fNc�^21P��=V�M��yB��hl���üŏ-�I�[x�9�õjq\1'ݘ�1���*DS�7�]�r����:��Xk]����2�� �f=��PΣ����k9-H���
x��Хg�*͜�e����I�4jՓX�_���wI��SNY瓙Sn�ٚo��oZ�pfU���{��N(_i�h�X�H�9V$ �U�+)�ӌ�!]�;�ԗA����*�YE���b�d�jҝzؾ�,ΝN�mp��<����u�KsX&�'��t�5���G��f ����qڳ�UE>���8�8��z:Vb.ȥcXc�̡�*�W/-m�fs�O_S>�DT
�ȓ����_���V-:4Mt]�V[��Ѹn�Tyc9l�����0;�ƕ�D���fdd3G�ئ-���2��!uj�E��)�Y�sXz����綈���Gz@*O��6̕e���[�7K:("�!B�g6Q�D�V�6o�	���O���\2՟��F�w�YJ�ڟ5y����F�-B]_.�
�q}(�&�G�-���YᲤx��K�ZM��l��n����%��i��<�s���9R�e��tcg0�����ζ��h��3�J�0�����FWg5>��>Z��ՂyZЩ��x�cAN윷���*���P�n�������A��%�ҫd����]�X�+n�,�p��K�`���!��qo�1�̨�DE�y�N�ˢ�ZbK���{��j�ᵋslX���㙉7I�r����~�q��!���k�����j���eq�N�d4.��R��A!��EA\f
���9�=XkoR, ��挦��RvRz�����GF�����v,U�NyM	�����d�&qQ�&�N�#�n��%!�|x�v�d���|��W��FT�ޱ��̳�Y�����׵Ġ�Yy�n��3��5o����i�'QͷBT����r�h%˺�e��	��u������܄
Ƶ7nc���9�J�[!��Wb�mۍ��݃����]7C���ܗX��M��^p3u�e�6WA�U�T���D�Ǘi��NY�n �ioԁ��L�ƒ�Ԏ�=�ƴWK�4t<�ـ��w���H���5:���mG�fe�C���C�X6�qN�/o�U���ƛBaFL�A���g:4�K=��,t(�ku���㿷a�O%�N��qꂻ:ңB��[�)r�t7�u�)Kn�t���)�}�4JP�&��P�G���%f�*��e�r7�mG�ŅM�v���Vu���2�w�8���B�����_a�wX�c�Q��nRX9n��j]XS��]��t�����2�n�7�ө3X�Gg
)�rR�)�m��z�`V�="n�L�*�/i@��F�G��]��`��m��S�àŸ��
��KF��2д2��1��N�zMa�r�%=�p���h�YDj=V�W],{0�rNF�7�kJ���u��⡸��%F��;L��մs��8EO�E��1����wNO�;{��Oz o��
�+"��#�+�(�	������9�j�A�R�/3��f�Veub��ʲ��3&N�EL�b�V�ں�^�Ʃ]�R5w�{đ�5x�@4P��p�W�h��wx]ZY�G���1i[S��d�}���4��{(�Ԧ�T��:֝n��g@m��ݸH:�
HG6��R�'��(����[�(4�����U��9�g�|*ξŢ�¶����Gըn��Ϙ�7�Z&���X&�8,:�����؋k�`����c�`���r|,�oq�2�
�q`�X�}t�-�۱2���QpKsy��7L&��U�B5�3��xV��4EO�X�+�P�4k��n���h���w�/����8&��ý G��>�.�AF�azr5(�+)�o�l���d���x��iQx�5����V�*�9i�"�';���P�fK�������q����}
�e*6�F>О4M�
wZIz0��U�^K u)Q{O�1xz�#N��6L.���GFotq�-�=���7CD�(]��K)��wn2�}��N/!]1k���L�ܵ����8�[��sw�öo�P0LO�ճmM�d�X�v�,���+�U�F���G/�w*=��z�Wq��ӱ�C�ڏj �3���t4�QX�r�dL����G�G�"�Y�_m��Um�g�,e�b^�z�B�����\�7h=R��z�Qڌᜎ[�u�<�='gX��ӧ	�:��h��a���j�!x�q附�Y LE3;��M�K7���5���]$^7Ck��d;�Pm��_b�����9A5���^S�KR�K�o�쮘WR7w�2}N�"�7\���t�6)���C�A�qӮˍ�u���h+lK�1��/���]J.h�}�0Q6��^��R�7�-���1)����'1Z�*&��sQp�7o�w��վ�7��w�JU�M��W���e�Z7��|~�n�`w�r��V��CW�J�s�}�52�}v"�{���6u�L�Kwf�������2��s��l��Ǘ&����6��:�.Y#T�b��¥w�ḪUv𺂖`sPC �#7���=�r}����ĩR��	s!=K'"L��i�{��u�k`:E��\lجaܶr�\3�EL<�=�c��n���7{�lV)V����DvY���5[R�8R�kqQǓv�V�&��|�O�Pٽ%��C��m4RW�hpL�'CH���#u/�n��k��U}[fA6ۑ�[N����8z�c��Tt�&Mݪ��]@����#�1Uٚ�YRL�F���}ϴZ�b���x M5*Y�ͷf�ʎ<���0�12�isQ<)R)wZ��S�fJ��EˮY}�Aݣ��wˤ#P�n)���X{q�:6�X���VR�Mi��Q`.N;��I��a1�t�;���ch}ׁ�y5�m�R�ܵ|�JRnZ�Hit��z6ԷὍ�X�<��u�,��Ȏ<�",�����Wu ;n�]�a˵g�|%E'�ۋ����ہ+4�5�:�AN=���R�J!���܉0����� Q�_+7�PU�:F�w�@�m���㹌��Vm��WZC+Y=>C9�u�yn'�Ie��I&���w%�J=���7c$=�ą�%n�5��"i�T��>��m��k.+�)"����.�:)�����a3^��n6m	�M`φ�t��}�خl�.���zWB�|��iau2ٺ�[إث�)��N�4�HMG����)�%;�]v��4
J��r�4�s�SӪ"i^Aa��'{��8-�[�q�]@]�ԯ�y-��f��㴄1Z��=M�i���@ح�BĵVnt�wS�W����l�n^t��X�� ����}�����Lg��T�{g�n?���elFd��O��bEf��{o�Ǣ�s'�__l��D��]ܾhU����A�x����V����0�A�]{ʸ��3q</jj���O��K�b��Y�m��XW`��l���o�wBXr���]+���s
�\|�M&�����h
�-��g%3R���D�@mmh
�j�/�B��t8*�4V��!�#SM�|H��@eخ0m����*��me�|١�xH]j$.epѷ�r#�	$.�/����:2�-�mh����c:��.�P����"0l��[�
��b��n4�h ��w���uǩ�,:������+{�j�ˋng@��n+��{61'4��_�Ȧ�T�Ջw@p�p�4�<30�֗-��z|� ��АX�*v�܎�E����Q��H���'Oj��Y�w]�\ �`���ꥩe:�nI�.�$�[�c���m�q�Tʚ�����д�m�a�2�3:��7��&�Y-GT��ڴ^�rB�=8����Q�S��}���aC!F^k���%��kJˏ	Ļ�f�O�-� m;ۛ�02Aj��R�	��)�<8���\�
L��ï�>������+��y��l��Jb��`�{1T��1��hO���P8�D�]�ޫ{���[ըs�ѡ~�|�����LLj�ޡ+��2�;!�����+�T
��wi�ws��q�����6$����1���wN�L���\&���$wt�`��d�%���s�1H�s�#���sc��26"�4�J.�됻�4Ȇcnr�4��w]PI��v���I������wK������;�DF(�9����ED�%�\�TE`+�$�.0�������9c���
�	�s�(��f�.k��N��7.:i.s7w1���"��ni2h�뎺+��D&1�ӛ�v��q��˹ � c[�.[���)�p� ٥2�2f��j�ۻ�ܤ��E���wutƋl�Ѭ��'w6�&
f��QY"Is�
"ƌY4�L-��h4�ݻ��h�H����r�rk����m��5��[+)�Zy.��W��󵞚A��1���ec�L㘭�#76��{ŧ�]�\��c���[+������#�����q+mAа;��ϛj�aw�.�����ؼ�軰�MN�%�����ըCCyW���ig�=y�S=���#�u���Tj�����W��Υ�kS��Ϩ_+w��F$��^��l�k�>V%��NY�e��j�)���m1����^b�?V�5����D�����2	��0����!�qZ��77Λ�x'v5%r�~�l��*�=�%;���|���޵�'�zD�oN# {Эbv<�!�bsnB�Hj�EC��N�~\vx��A��]%S����c�{��
���ӡZ
g��[��;^�Ͼä��o�'�y|��@)u^�C�_.�y？��v�Pw剛B��u8ܮ��ɵg��3��-ې�$���!@�_!dy��)Շ�z��~� 27"ǟ��J�x7�4D�y���f,(�]2�8∋�D�N�uy�3�wLS�|7�\�'u��VRpru���fZܵ�Д�^F��M\1q
f�~�.2��B��Pՠ�Ag���m۝�~�,ſB12O����S4��	���/?Ym{����U*nkv��ӫW:����V��.bX�N�h¥X�øxz���f_c�����j	$��1u�£�xX������=�k \���B�ie�˷��7n3���N|�@�yxq�P���o���W��Y�t��j!Jx[X�#�k��\i���uC�u,�����e��󭴭�L������@�{������ĥݳ��:3���7����H���$g���ў�{�~���jCS�p�D�@�5�Lx5	���p���V���NxdMOS�k)�Z��3���o�fR4P��0��y�1�әa}�����$CĮ�,뛱��:���}j�@u�A�1`Jwl�U�3 �Zh��fr�+>gQ�3�ב�s�yp}����+�mA�S&���~���i�7�=Vb���-���):��a*����}]M��}^�cjB�r��pR�������T�cT|@�?�����N`2�-�g�3�0oR��XW��υ�l��n�m��w�?Z���Ҟ�[�z���叞��y߹�;�3���^��{K��`������p�+�����}-P�&�^��T�
���+�M���(��<`6FW��y�Ô�\d�D� �{l3
�뷯@Ͻ1�^y�����j_�q���BC)K��$$%6z����>��(��#{P8�l�զ[w<����5H���L�a�'����FI��!Skf�7�=�uD�F�t��D��7��Y4�m�c/l+�yt��2�_e��mFxFx1:\T�%��׻��^X�WY ٙ�e���|���W���{P G���;Q���ӱ��{���*���R�f7Q�{U���Z:hPKJi{U7KrG�K�St{D<qW���u����6��W�����"Y�� �cc�k���PÓ�8ʙ�>���b�y�����Ѕq��yÖ,04��j�ﾅ:�|m�]~!�e�9bW�W�A��W�`�f|�Ǣ*f$�֭_��X�h�[!8,h>2�V�Y�/װ��v��2K��BxW�[9�|�lp�ET���s�w����`Y�Ɂ�}/����1=��ڴ�������SA����j��_��UIb�����Ո��ϟ5�P�wx����	&=�{1]{����U��#'����T����ڡ Q���[X9�Z���د
^
\��w[Ƌ�$mD%���9��Ys�J�5�+���йuPF�B��eX71�ۖ&S�ׂp]]	[�et>|ѯg�2��BI�g�\�c�j.): V�S��={��mr�^@���/s�"C�_v7w��<��K-@��w`�H�^�9�X[���ݫI9���E\�������Ԫ�@���k�5w��>���\�f���ҍ���<y�6�/hh%�ۖS8�1>��RV�}�0�t�CO�k����;��RD,ez��J�{q��dBJ�&C���#���T�Qy������:0*�\���C�]��
�O���p��J��+����U�=8��e]�������*�� N�`��st�o�e3V*�BxmY����_��J�K�#�/Z�!��:�'<�}���$Z<�����֭�h��c����zt.S�u5Tc{S�3g�ڼ�^�{w�Wk�^�N�,#�ֶ������������)���D�FǞ��R�������N�K�����i��8'M���dHY����L�ڥaV'�&��u�B*%Hglzh=����u�#��3<�׺�MS�Q����C]�ʉ�x}X��Ҩ�|%4��>@W:�l �1����D�������=Ba�ꆺ�nkv&����+-�օ�lk�Y%�o�~�D�2'�Ⴒ�׍�x�.E�߲v��Zb�ׅ�������m���Յ�����:�t|����m^��Њs�����)1yR�O�m��%����ۘ��/�9h]�v�
����U��nS��
Й���^jpec��C�N���z�֖qX{ ��=y�.,���L:ls���hq���`ڽ���/zP4�{q��`˃��O�f�h�2���w�sCW���L�~6��O����E�S�EC6$B�0�@�	T�z�ni�Dj�rN����(�
N�3��Ν�~��u9�m�ϩݳ"�UT�p���Zݍi�g�I��ΕLT̵^Y0Ǡ!����Q	;AC����c̚M��P��o�}W�nX�����0�T�;sQ��#�|����N�p��sl�-g���-,g֮b@�sq:�w���P}]��G����0�t�k�g�ׅ�n�R��\�u��3�y��8緷"�����z	]b3��g=����![�^G�?{K��J���(v3b�ϖ�Z^��}��z�R�I]Oq8n�|��3��
��l\�k6� V��딇��ڭecW�G�Ɗ��=K���������F�����c/fX�Q8$O��X�q�L^cIڬ�fC~xV��r�Q�~��dܪ���m���v>�N�������ǘ��CW,���ۓO���;�v��*�����q;3�����*���~��[���z��>�ƅ����oOZ��-U��rWD:�U[��u-��"�XD��K<%�|[�~{�f��5:3e��X�X\ELZ���@�&�t�,��\�[ĚΨ�סc�4J3�j�u4 v���K�%�@��V�X̣`�w���6sf-zR>V�owtZ���Ir�3.ǻۑ��	�¾�Q8+_�|�� �2X2�cuV�4�~�5��)��קv��n������5�C}:Ie}fB�6�Ƈ��B
p��z��̠���<�9��v�� � !7p�	�3�/Wh���#��3�]Y=U���wN��,�Ѥ�l��ܨ�a\j���kq[��,�~cUl6Ϯ�b��ʮ�A�5y �vm���c�7�s�. ��\T�k7�_J(1c�i�r0��?^7P�;u,�M-Y~����H� T`.��t]g�{]���\�����@
��-�{���jBYʻ�k}Yi���*>/�"�U@�?�
&<�7�  ��MZs��c��4�����V���_�e`�s��J�ᢀ�9�#
��z̦{Ov�W���ޤ'o�Y�zx�A�z��Ѥ���L|#Q�S�`�J�9��@�����9z�+�<��X�f����9�X���|���[PEDj�ɢې1���V����}刨,[a7l(u�6+殛ѶE�x����z;C�^?{|����X��|m�-mKNX�P�6&lO_��+�"_�{�����Z�:�vz$,E��h���t�}V9�}}"�v��b�P:����c)��-�t�h��#H]��j6����<��mWm��]���� ͸��"�Z}������fY����=~}�5t2�> Ti�uy��Z�F �Ύ����~�����i|����V��C�����]gy�C���Y;Ҟ�;�J{u����C}��Z-�}�@�_m�]�W�������du�W�Wj��Q��׶�����b'�W���ڰ��k������QU������z�����pU�N����>����J�;����ӓ��}ˑ!�v�>sJ�� �/%� y��q]��7�+/eӋ܁�	��n*�B��؅>�=�\��3��Z:hPK8@�����g���Տ�r�Z��ݡ]qէP+eˣi�eyڿ��(^��,�j �?TJ��*�����X��|
a�˭U+\���+�鏮<���ŀ�)��~�������m��(w<�R�q��$�p��b�a
�ftk����(\*�<-�-���3�/Pq��ᾲ�w���v�!﫼a�+�s���9|UeG���>]�4����t�wJ�o9�jGFd��&`{����$�w@��/s�k�P�(�)������oSYi4�o'A�I�m; Wm�.y�a�������c^��@ 2��|/��1Uj"��6մ�����C�򭩊�s|�Tt�39�]8!M��ssU���\���ƛX&���=X���U�L7���3�=������� 8*`4{�Cx뿨*�4�Y� M	���t�hy����3�Ax���#%z8):�H�Z=� *P�A��C}WISY}/xN�K��AR@���h��ƈb��%16sl������";W��~�����ܦ��u�+�iL�O�50ʲ�Oa����B�<�MT�}�N��jo#v��6�s5�y/��9:]��J���j�0��7������	��v!�`)�3�J��[�I�UX߳��غ�K}fNτU��?5�vP�^���Å��n���Z���K���l�F��M�PS���Y��Ч�@�t�c��߰�j�xTG����8&�ቫp�Cţ�b�$�^7��ǜ���~�1"��l���������-/o�-����M�{���Q��/'`���8j����7�J�Ǟ2��٬�lܯ��sʕ��l�"�.{ǎ�u���g|�j��3ʴ}G]k0<��e���Cw�b�1���Լ9�-��V�i����K,���x��8���+'�b��`�j|$����mX�;�,�ى����fޫ���WB�t�D5hv�XJ�5�ٱ5vU�w<ځgV.��Vd�Mn�-ƞ
	�R�5��D1�j�RA�7W��_+�v�X9w��f�`����@�:%?&)�!�eP�Ƕ�gJ���X�;�����C���zW�H�s+Ml���wDz{�:0����~�6�!$�9J@�P�� �1����D������\�p�:��>����Kg�l�wj�F(�P��Z��dK�!�w��b��ڰ5��3���Û�-�,��7ʪq�;���s�*��.���,�����T��ۧq_�
�����;3��\Q,m�Ja��ю@���r<�i�H�
Ҫd�����M?cV�b�#,��:��ݶc��K��5b���:6�ߊ�6����[=�W������j�xQ�WG_�V ��V��t�|��h!�-Yg�LyI��6��r�cU��yk]]�ω�#��}Y�ف�j@j�V׬���-m����������<<Uڻ���ٛo��j����Gޣ��ZQ>��Mv�f3^�[��3�8Z���z�
^��WE�2蠂j(���0&!��J��ig�^a��a�:w��2 D��|c�/��|h̟]�g,%��IF��0��FyT�8DV��\�֜ʎ:3!w�c�t�U�w�x����2��GSS��>bq�hZ��8n��3��O�gW�X�M{gw��즪�Å��n�w���T��6E$��z��=Nq���Խ��Ͻ�������eU� V?�͋��m(< �b�Z���c�����}����~^���/r�)�p�,���L�1G��_��M�^��[�����w7��<��"v��Pw�Z5��/+&�ּ�l�ͻNN��F9�ucV���d�k�0VfP������)�W��U�
��N'fS��E��o��%-�z�]y���O�;��W��ϰ�]���Q�]���Yt�����~bU�������|1�L_g�ωv�p7u�q����z�L�W��	�I�Wzj�<�*�2�%�,�Q��@Ye
S�"�&�zh��&`�Z�m��MX�@G�0��w	��J��|���X�k:	:��P����x�-y�Tc	��^�k$C���ϡc���Ie��a������M��������A��Kx�-�߽/�yfp�S��9�b�f5�J~��R��X�#��F=���n��v�T��f<��b�R��h�Q,>��k��x ��-����g��X(\���Ώku�H���2W^*�tV=�ȆE�چ칵�D�%��y�8#8����k���V!ϑ�&�o�э��j�f����;Kx�v.-�W��c�4�6(wY��py���jjk&WKB_T{z���C��u&#u��,j�Ϧ%�yk1GCn�2/�p<�o(����b�M*g�T�&��9xxօ �n����!I��2r������[ҕ=U�=8'T�-�E�����"[�K�)�3�4���
f\B��".w�+���6[�tT0՘~�VG+&o�Ԧ��(]g (����N��a�l�d)��)#YB�f<�+��K�y�Mɫ����ib*��<�l��>}N��L晩#�'%s�&
0Wk�Z������.[4k��)��gKAA�$fV���WS�wS
�i|܊6�qPͮ[�u1̎�Y�RWw�6��x��AҢU����̳}�]��j�e���࿍+ѡ�$t�=�)v$���cX��/��pX���U���
�
����.�ZrL�G�#�續��Ǉm�zp�u+����]'��ۉ�<�Rя���	f��_f���W#�(�2�)��������x��Pt�������P��\Ю�δMct>&e������|���M% ˸˽Zb�����Ε��a��ݛ�Γ�*!�˪NA/n(��7;Wh�ʦ� !u�KjY������iQ�:��mh���\4>ץ����<�V|%ǀX^��Q�:8)�M�x��hlae*sy%��1ԤobG��t)�73���>�/iYtw�5�`ԙ֣�9urK�����sz���qi��LZ������vʬFS���=}79��+�1HsV��qc-����pj��M*�-"a=gV���y��e�Ujׇ�N�A�7�jm]uv�+��V&	P.�#��e��Լ��)ȵ�X裂�[�1�8����	��m���$��`�uo�=3i��kC��aZ��k��b�U��n��ܖ��mK���;o� ��h�p�1��,������Z�䭴�ڽc9����7�aJndr�f.��7w|�)]����wf��R��I��M��3��Y��YC�4݋�9��RQ�J��j[�r|��Jn��0��7���ņ��ۺ��b
o�B�-)v�^ެ�w�$�:Oi���,B��t������ۥ�Lx2^�Oei�C�TZZ1m֬�B�^�n�蚻_)��76� ��-	6�\��[{R�[��ui��1g;7ׂ��w���
�F����}����F�ĵ9�m�V��E���:5#������#k%$�+��]�pDMF:ޠ�#�g�%E�YDk�n�V��� ��j�h�:M��r7�Y����P]Yv�3�v����p{{m�*	��ܐ�Љ�����%�Y�Ǻ�qr����&�w�B��}ż|�qɅ����e񆷖���Sco/a������`�*��\�����<����߭��
4�H�"D�0�F��D"D��w\�˅��#�(g:�nQ����e��6ɩ�@@fBQQAI��h�h�DmF��cW74lXɬ]�`&I���wF�m#T$h�EF6�e]�i��Q���F�%�b��)$*L� f�-I4r�;�4�hȖJ1jM$��@�F4$�Zf��k%	�W5�usa,�ld�4�b��d�a���%2]�@�K	���bM4f"E�4Y�3	���1ݮX��h�+�!2le1E2����1���I��r钙H����*��N�!�q�[Bv)�w���f���5} 9|�3tn���\	���o�
{j�ILb��nE}ar�쏺����j�ӎ1��&���P�U}u�uy�-�׶�/���}�^�^/��owί;�77��{�ץ\��������Ү\��:���}�|�uzZ|�������ѹ�*��{��}����|m�����'�L�#)A�����b��� ����D}� �}"&�>��,}��?z:�#ϫ�h���^i���ʿ�
��|������^wj�<o^|��׵����ߞ��o����o��h7չ�����LTW��1u�z�@���DF�1�uc�񷍽�����w����ޕ~�o�����|�ʋ~+�7��|���޵��=|�{_�}zzZM͸m�����:�5�j5�����ھ��������ǩ����F�7T[�h���"GG^7�������r�������{[�sW��瞾u�����o���6����r�}~���{U��\���y����sz����_�w����z_�w�oJ���{����).����u\��Ԫk��������]��~v߭����^[�}{[�]����|�}�GЕ��b>�>c���������J����_W�x�>��|�����9�G�DX�>�Dz9͏��H�� ���#���ũ{&|���^� }�f/���->u����z��*��ח_[~�o�ܽ�}o��������kŘ�#�\N]D���G�}��BW}��A��>������_|�B��[����uodlw�8�q��yY�#�~��#�M�_���W�����zn^5��(�W�A�����?Z�W�O�~W��,}_ͼW��_7�n��[ү�����^܃�+�
�*�7��}D|�?�̚�k��kA��rwח��gg���xcү���ۆ޿�y��~z���cQ�����_��^��޷�o�x�+�_��<�-�[ǿ:���{Z��W�~����uy������/\U�sD}G����[�s�˝�m����1��U��_w���[��r���z��n���!������A��s�h���}���߾o�����oϝx��x�o�w�~o]��|[��{������7羾�o���"G��H>�*k�C.�u�5Ų �_��^>���������w�|�or�ޯ�ﾷ����x����~{Z�n�1�S� �������b< ���#�3��k�����m�����������[¨�F����ΡK��X(&�-�.����tu��^㾷��pY0�"���#��,�,֌�o��ւw�Ǯ���L�����M/�mΛ��7]���-p����7@����8�z�����nQ(P����b�(�u��hf����G�&n���͚�oq��·:�7����׮���^��K�o;������_|��_��]󪂾�O�R����ּ_V��~_>���|_Z�|_�<���h��~y���ƿ��WϽ�ήX�����>��o�bf)��u�qW�w�1��>�m��}��Xܪ��w�x����}v~P�ԡ��m�}�ӫ��ޠ {��/�|[�/�h��߫��_ͷ�~��M�ޯZ�X�Zq�����}X)
����|��x��r����x����oJ�˚����o|\�}��oO�\׿]�^���w��?>y~7�nU�rw5��>#�|G��?A\~���G�334�`}O=����tB�X�xGD��f5��߯���+�ţ}~���~�mzo�ſ.�*"������KO�ln^�{U˕���[�|��x���ޑB>�>�����돸DxG�,�փ��yG�{ܡ�Ý�� }�����EC�5����ڮ\�6������ץ�\�^���^�|�\ޛ���������*���x�ۻ����Wv�W����:��8������G�D!X����d�����F�7c��������H���U!Z+�}�ޟ��|���z��叫�o;�~�M�ۼ����[~*�s�����{��\����^���<�ֹ����oK�|�>��~�G�}� }F=a�%�r������1#���GQ�1"DG��{��W��_���ޫ��F��wϟ޷�}k������K+���]�����^/������s\������__|�UAF��U}U��jc����E�\�.��#DD�����O�"��|DW�������szm�{�o���o����m���Ž�������Z�������^5�/�wϞ_������-�Q Dh��3������YW�-�M���c�V.{G�xG�" �"9��>������x�Z7��ݼ�u���߯���oc~�������/��^7���h����o���/kE����>z��~{�\ߕwί��~���sL�ʻ��z}*-�H��_��ۻ�����zZ5~�����]���i�^��k���/Mx�����^���5�w�/�߫Ţ�z��ޟ�~�ƿ/}�>ur���k��׵_7�n�~tX��*���5�#�o����j��/ӆ���8*�\���@��)g)�,�}��C�+'�
.WgV�qe��ч��G�c�R.ѪF��.��fi��67�˕��a2����{�9�2E:�e��R�xD&�r�aK+RŶ�ۢ���yᖙU����Nm_����������Drn�,\���}W�}��om�}[������xޛp���S�mzk�����^����_�{���s}W�x���^�������om������~���W�}����B�}���8��}�"Dvw�����}y�ֹ}~��W�Ͼ^��q��Ay�X���>4tFq�4G��>��������6��߭~u�W��v߭����R#�!" ��8c�#�>���<�����r�1�����GDY��C#�������^�>���i�������W.�=y����{o�߾[����~|�y���x���w�_��h���s"�H��>̝ޞ�!���
����ݼU�s�_wu��E���]�������s�{�������~_�'�ԡG� WM�x�H�������Wּ_[�{���\�o��/�{{X#�"D}�iԢ�暡؁P�`��M��}��?:�c������W���׾��]�ͼU�s����]�F����.m���Y���zm������=~-�s����[}�ƾ��~���-�o��H�c�U7�}8�W��_X��k3�Vc\����=xW⿗�E���ϊ�7�{k�x׶�k��?��ŧη��痧�oj�.o��צ�/���5�{��zW-��������oj�|[�s��͸E��>���ףh�_��ޅW�ૠo}^�߭���o�|�j�.��/��矃Qo��x�������u�o�ۼ�_�k���m��o���x��~w��؋˺������k���||[�_��yz}��>L����<�����,�	q"$Z��}�����o��o������_[x7������ڮ\�6�<~~���m�W������{�}���O�ޗ�;WǍͻ�o���^����wW��x�\�|���Ωp9���린_CGΌD���~z����~��x�u�����ѽ�ʩ��D!`��nb�p��c�B"sz��b��B/���""���ޘ������LP�G�$D@�pB/�x�5���[�N`_�]@�1�"�<3�X����^Bs-��rꙐKk�,P�N;K���ls�Y(gZT�m�����j\���ٷ����)w�*�Z�2n�j��]h�5��$.ޝm���פ�ol�v���w�	{$�GH%Zs�ʧ�=Ǣj뱊���8B�m;ƝYt�Z�%k3��n��G��_woC��5��K�>�l 2�דB�L1�n�����=_����O�bB�����~{�����^�})�^O��Ԉ�Q��py�3�E�6�y�J�!~?m�l���^�W�.���T�r��
��2��}�Q����x��պ�J@j�ᆴҍ~P/ޫ�j���9`a~
hz܋0�d������a��x❜r�g޵QN?�+m{����xf5[{���}�`y�VxX�ؿj1'��#D��7&S�Ԣ��|�okk���a�h��04�xie��^b�W?S������`Aw�@��a���:��Q���@��[���r|��*|O�P�蕢$���<�����δ��tC�c�;�{�f_n��!P���o⫂�x(U�����Vx[}4w��C�{�u �{�x�����4�]��bE��E��@s#>7�T�X�oeߡ�L�����ZeI�w[x�\��ݭNiܱ�pxy���y��GI:v,�Q��B��3�٭��/*�]����.]�^�hl���r�-z�P��:X�U궳���^�J��$�L�I�>*�In-���c7��!h�JU������Z'2�V�n���\��_��+�a����{��e�
�9�}�ߢ����Y�
e������i:^��Y� ����h�� E�C[N�3�1��sq�GD`E�%�w�]�L2.������}�;�d�P5)���m;����,�>��P��b੶_�N	F{�,j�-�3 �w��d��|Nb�cYT��E,8k�u��=;_k��� D��oON�يj3$۔#����΁ � O�'^�zB&�u*υ���K�֍�r��<"�Ψ�+q�'/*�K����"Y��'0Y�D@j�HR�\	���  Q�>X�� >xoaq*S��o�7o�����xY)��[�U�Ą+L ��0�Ǽ��L��ȴU�z��d,Y}�i���Ԇg��
���5��_�:��S��x�y*�Wi~A�|S�w���5���J�gQ��7�_ h�r�fW����y��_0o�z����P Ż��B9��ŉ�%����'Uxj���\�w��G�>������k�v�H��=԰o{N�"��v5^?Uh�<��+�� m}��1ֶ�-�̛�>�݋�PK��oq"�+�o/�c�z�O����.7�{�M3r����P�v�fgvq�x@H§y�mS�7)�9�ǲ�2�C��`@�G=e���^'�ʹkV�n�\��)F����O�uL{)A�11�xTV7��V�Mb�u�)ᴜU��
-\:�}_U��Pܓ�������������o�'���n�t���X�`۷���2:�߇�)@�ݍ~�;��Ud�6��Rښ8[Y��$vҩ��W���V�O58�h�V�����+;�8uUxNo%h���V	cձ���rt3�NN�}ˑ:M��Iu�Ec���'3�RF��݉�<�|]���@�~�u��*��ܗ��=���EȺXK"^��ꗾ���Wa����M/yT~@htmW���P,�:��W���.
������e5�0bM���J�����h�7�l+����6����1]0��}*����W�+7˹�����T��r����/#7��,�P��P8���q3TVfK�_W.N��nzջ~�pN�����3��G�
�Cv�����F�*���@C��g�/�u�ߥ��1��Ad�NuRz��<�K��{��WC���u���ͯ)\@�`?�@X��{/m^W>[�#�¬t(No>�)�E�b*��6��2�Ո��1$�A�1ޙ:���o&U���b�\Zb�n߁�
�C��^{��%��带nCIdtUG[�l9�y>��ƙm#��r���E���1Wө�eT�s���͡d�T�ֵq˩NѢ;3$k���t��X�S�y�r�q�(��GT���;�r�S7qC�'+G}���sEw����jg5�2� �hЂ-/�zc�,���>s1��M�S�u�h8^}����8�[@�@�G�R������B�UҩOHCL�|��`�U����x_�R��d��΢���qs��y�����5K�W��.�hQ�!}s��0�
�zb7��J��02acyWמ����f>���iz�ˀ(r�ïh�����������C���Z:���Oz�ѧ�)�cJb���9Q�T=;ʼVz¯,S������B����0{L��땯Xî��@uZP���L�[B��=���:���%������t����)��9V��ߌ������=�׫Sxe3�'
��=�����@��s�{�������֐�k�����/*����<6Q�2Ǩd�ɹ>�!���P�Z>�:�Y��N�/*lFe�)�Qy�ܨ>��r���,ÈNpK6"�nі.��Њ�!������� ���4��}ճӏ30��^�=61���bgFT��6m�Xߙϔ��Ӓ�R�z3���L�����|�o�ǩ�5����
Y[k⍺Lɥ������.���Xj�����N�rn�86���<�	+ٔ�OU�)[�}#OZ�gd#:�ǽ�I/6�h����}�}u5�,�v���(�:�����Xwrˮ�ֿ�}��}Ty��3'W��z�c�z�ΐ{�w<6��B�@���K@�^dK�!UT��g�R�^+5���5��^,\���Sg�d�q�@,2���mםϽ>�=9 7�G@|�J�4��>�kغ_޽�����\����e�Ja����ڋn����Ex9�#��%���U������ ����m@�	��!a���ݶc��g�_w���{h/gz�
�^T0{&0[�z���C�m��@�@������|��\��F��jv��-Yf���	���V��x�g��/��>�zv|�����ӓ�����#F&B�����aA q�:�J*O�{\-=���t�P���C�Uӓzd�����T����^��ZQ��A�Yޑ��i�z��<ҫ�x��	���M2(��U��M���mj$IӔ��S��ё�U��.��n��>Z�FU� Vw�ڌI� +��Ok8]�����w=k>�Yڭ�0,O��(�d��y���*����_c���e�ᗾ�S�PWs;�Uͤ1z5Vd��G�g{ܮ��t�Z����,����pd6���sG�N����5��?:�Ks���ge��jRQ��Bu�r_]7it�g(R lz��tO;�TA4:�`@����7�wu�81�tq7E��S7��������P^��kV�@���yj٭�Z��ߏ���dܵ�'~ۮ\۱������['�e�����{ޫ�G��^��(�	@��\
����>g�g�U��A���WC����n'~�YX�ey��/޿�����5(Ua/`7�U���,N�� =-l���~m�Fyd{�V�������cuV�5���+uZ0cV���dcn-$�#��Z���3�^)�*}g)���Y��𡢺�)S@��T�hJ����g�^��sq��h��	;��^9�tֻ|��賽Y�(��*dh�����g;x|Ԗ^1���T�.м��J������p�����A�-���Q�[�:s�)r�[^����\fZ�m�񔼷�q�?+�y��h�p2�Q�Ut��-��t
_m��bR���+��ԂϬ�6��_�j9Sմ��g���]�B�(�?Rs����JT\^W;Y�����9NYG��ٜz]�V44Ӵ=}Z�x1���n�uo�W3pu���,��w�������s�,v+�PdZL��_��"��Sy�|��R[���D����i��BGC˄�eT�_.������-kR�n���܎ȭ�j4zZ7:9�D/�	wh�W]a� �s�f�{�.h�-�h<w���{o-L$��.��w:��p��Ƙk}U��}�Ǵ��o���d����w��*�Pɨ��h/�X"ы~N�Tۙ�Xq?V;���īn}3o7<����[P?5�8̬>��|�ڈ�R�4nt�s`f��?n%#o´؆�fz���n|�F/�1-���w��*�an˕׽��U�_y�^���.��	�b]f�����C?�Z�d�*��׬�o�����ٶ`�7_���;V	a�w���N�C�ޱ*��/O��Z_����b�H��it8X7k��_ޝD���/�
��2���b�G��ک�54"p��<���M#��@$�erC�~+^�D5��i��e�e�>1�
�� �UT0/�0ǖ���u=�e�,Z+��lϳ9���8�F�+�r�����xd�3�-I�D��p4@��u��3��X��n�5>�.�����M{�`lJ��;�4A^���I[1����UJ�G~NS+����H�B��X��YU�2Wy`��=Dexk
��K^�M�j�fD-�鏮Ly��7Su>q~��k����
���Y�Q�L��1S)k���C�Wy��;i��僶9���d�R'�,-�ٻ�:($���%�e'�Z�/�'�yڔ�5f2�̤���x�{c+��b�����/����0)�"V�t⭡�,�Cyh��t�yI��'�]v��q�J���p��9���f&�e7��\��ѽ��R��FE��/`�����2������v��]�sl����Lk�:��Cq���Ve{W��������[Q�J<e�h�ؕmsww|�j.�E]�J���5(�,K|��-v:��2���8�2u����D��9��Uj:y7�^.�$�ՙ#ᢖ![-�J�<tA�+q�o2�`�����	`7�<�˽��7S�݊����^uf����\^�q.�	�Ũ��q.PQVJu�.9��t�W�cs0��@�2�m�p򅠩�YǱ(��(.niğ�Wfa����PmA��/Q�t�vq�͵�g5���fYG��u)U��0f2�Ѯ؆(��g,fS�rtH�{��D�Ù�e��>}�n��V͉,�#XZ�P>B9��6a4���F���؏�L9�^�)�Yrb���)��s�B�,pX1�=&#y+��_r���GE~�N���0:�U��N���	�u�P:�4���R�fJx�jm6��#Q&�S�.��w^��[��₮^lαj1������j����_@X�.v��So\����+&h8eF�_aǠ���`�{09�TP`���O3G�h޹+Q�����*K���GY�֩��$�&����֍ս:"����z*y6���5�:��e��C�x8��9W��3�E �>�]�M�+�L�4BW�4�$�U�)�r�����@G9@þV��]��7�>�ٵ����P�w���b��4��]�v۴޻��+���[M�Ց·���ov��'�Sj��Ԛ,gt��e�i1�f
�uu��`�l\/����ڕг��d9��+q��q�dWd�a�ه1��;��MTu��C��	���Ĺ[n�:nY���H�tLAo�w-$i�xD���X���}�W��'ό��%H���U����Y���vsE�}�sx��(i66���( �Db�&�2���db��l�(�f�}�S����%ɣ���>�m��.>�����b�B� �e#T)��fu(Z*����b��t,V���;zƮ��(���J�aw��
�x"G%h<p.�����M�sv���&��Ś����t��3[t�~����՗R�|4���`F(	�_G���1��C�s��ڷ�����]�!�^;L�y�Sj3ʂd<M��������&���Y4���j�Z��K�Xi)HU�RqCwn< �l�;��\�[p�K]]�ݭ��C�o�Z�|Ȓ�������kW����><�ש_Y� �RŹ,=�$�vkut>44a0�#D��T�)�(��wL�-s�@��2Q��eF̎T��ƹ]#lcRX����1�@ŰEF�$FƄ��0���-�F
�5##�� ��*f��aDX�b��\��cPU!�)Ki#JF�F�6�Yb�Qō�TTL���(�����cA��1��0�I�ABA�ݪ7,�QF���Ɛ��f��h�Z*L���FD�Q,���f�Q�h�$�5�c��4Tb�m����?��y��ׯ�������k��1�t�l�T��mI&�k�K}�g%M��R��t��h�XZ�\��N*�;/cĹ�ꯪ���{~e��Z�'@�_��[�S^G끖a!d���U�G�ʲD�K��6oR���~q�=J'ҳv�̱A�BS1q�!��ƃ��:��}R��>�Rf2��
.T7�x^ �C8>n�ιϲ���`��
n����F�� �9���3.q �`��W����+&g�8��L��PaaB����)�G�g�>/+��n���I�O
U�-��
�.y{�y��~ ��k��gV�2�oQ��,��2m���*�9�w`^;ok���tx�1Z�W��K��F:�o�&�A���$�7Ʉ�vY{P�Ed��r^�խ�g�C��5I�^G%��}G��:�Q��SJ���xz�����s>y���z�\���$C������9}a״GA���G`��e�?W���7Exv��P��
�Hn�7J1X��4Pp�Ո���5nb�����PA�b��޺%���<{���I�R��y�vb׽���e
�PA�}R�N�!��ڝ\G�S���}��}�=q
x��N��v����z�;Td�E֠�c�$�X3��W΄�+�F�ܙl�"it���ܽ�i���2�h�G렪�Ϟ�7o1��,�/��ts�6q�yC��X1��˻g�L+(R.����E`��;]�t[�ʖmXo7$h��O
Z}r���}U_DG�V�8���ͣ�nt+��U��N@7��@jӆ��c�K��˼kG>��i-�O���o�~��̖����7'�Q'~�x�f�;l���qR�u�o=�W`�l#�0ESn��6�n��F
��x�G��-1�:!U�d���\�y��L.���L�S��1Xa&��O���~Zd�ҫ'��Rꄭ������I��⪹b�8]�y�c��H=�����UօQ�Wy�l}�D��@ƫ��Z������ӣ�S(&}�?O׻K��Y�u���e�_�;�zP�������9k�b�ߺ^o�`�=@ت��n�^)�|���Cl�S-8��ݑ�SH�r}�{"��O=�q�*s�p��$�s>�cY�!a���ݶ~��\����S:�.J��{�lٹ0�^��	���>� V��(o�1o�x\�P����N�AL8r��������|��Xx��čd���� ��k�Y&��?�����Fq�W��f���.ו|�U���x�Nu:���sS�^њ�Q�ˋt�]c��Y���_!M��a1�n��-�n�]�L���� <����� ��o�{�n2�r ��6ڒ�V��*�e���_.�FZ'wiQ��u�o��}���;K\{����͹�ZX�DX����s^F�J'�a����Z��7Ģ�"��<�#�oS��Z�{k�Y�?#��J�M���	��4<ȣ����~�>���bIS�����i���2��'�֩V�ΐnr��
�[͇،K�9��[��2�v0ptg�Z���q�a8ea�S%Ϯ7f��+�=�b�O����[�/�Js��vo��y�~�,
W]qZ�}�x��\�'s�*�o��Z"Kk����/���,|cP�5�;�ps��)Y ߾�@Hʮ�^����vW2����N�o����M�oW��Ғ~��To��y|�����zjP�:L�?*���bt��/Ƽu�WZ�F�� ]��� Ex��n�����W�:�3�e����r  ��p�n����V�̽�x���\����_p5YT���@W��%OO!<G�ܭ��>�K�"�w���mf���N�����3z|�"�����X����Ig����=Q�ep�/ī/�\q�)]��{yn�R��N�Z_dݾaZ�Hn+�j3�;��E��!nl�
�g�JS���]���J��������}Ԋ�-�,�c��ߡ�����㕺.Ǚ�U�M�	YS��걌My�tw|�4�W�}�}_V�y}<=������~���D��Z�ʣJ��}ӟʢ�ǅ��;HęsO0s3<�E����nt}��P�8ʙg!AUA�~ a׳X
1�u���]<O>X���R8*Uy6p����!�E��u�M������?&`�����@�0IJ�����Ӓl�acp,�=8l��7�w�U:s�J�ϫY��'u�\:�諉���F�id�>a�]r���asF��T�ˢ��xO�Lo�T+��-��Z�:��E���7*��c5��U }�y�,����~5�8���_۾置��S&���~���h�5���_�<��E���<A�
� K�l�>]�w����Q�S�N
�{����;��sk�i�Ag�ތd��l���6Ū�V;>5�6ϕ�Ԭ<-�m�8\���c�A^]�Q��(�GZ�	�E?H�_`����~�ŧ@~�'���@Q�5Ѫ��8X6�	VUG�o��U�,{�!��`�ک�54"p�<�����������_�}��i��r�ߋ��x�Л:k9&.	k6@V��t����Ej��:��y%�<�g{���Ʒ%�����=�u6�қ�8�Z����=C�-#\��}Wp�N��9� ����V�2���+Յo����X:�u;�V�a���ﾯ����^8x��C�V���� �{lz%UC��^��'���tjy�K�^�<
ձ��.����S�����*��ɥ� FP�4L5Vߓ�})�������,�b��I�lw�Ig�z�šߊG:'�0��/j����TmW��}P+eˣi�ey��h�DU�]烆׷
��/Je�v"�H;FXڀdB�-z#k�����<�>�xVuO�Z�
�c�`�����g+����)�#����>:I�V �i�U���o��o��Yj;���{,w�
݆=�X������!�h6q�w�7�(��5�)P�l�;��`?UM�m�2�|�Ԫ/�i}���ޔ�.�Z'(��;����@]9�����K�� Ba����s*y��?[ux�R����ڱS�ϰ�#�3���n!7de��?>WA��mk��c	��I[ 5�_IXX��zj�Im4Y1�ng̕x�ㆈ>;���P���W~��w�@8^wŉK��R#�p5ʼc�٧U�x���c*��e��2C��yT�\3�*��4*X�{�c}m$Y�/8f�������<��>�����yJ>9T�S5$�'Zٙ�@�EZ��ˏ�xp�Z�w��c�[68-�ޒS��1�J��.S���c-�ɟv[Y��t3Jv�`}�)�^��o5��p����UW�US�?{��O�{\�?��y
�U���^G�����g]Y��6���;Z� 9�������B�{��Íj�&C�ߛ� wO��]U��#5g+����� �o����]勯��c7�> L�|���<\�<�N�b�o�4)�yu����V=B6���&�~Wq�Bǣ�3Q~��<~:��lG�S����`��Q#މ��}1���\w�<Eh�xW��hX������,U>f�`��ﾼ�~��ߛq���R�;�w�d��?��ٯ	�����t<���%�*������Z>����`3����E�Bng�����b#9���g�������ʡPV�+��p𿟓�!�j�r���-�����Nį?ej�9w 6�����߽�ם�'�beP�}�t�|#K�P��nYO^Y��[�)����h�@����0Ũ������ʮ�(
8��v��ѱ���`��f{�|�ngN7�i ]�4�7��G��ݦϞ�f2�΀Xo�i�_��dܕw�*i(��W�E�5Ե]���Ɲ�
]�w�]0�� [��/	0_U���
N���^y��vo�ߚV�����A:��V��^䷩Z�Ky�Z4"�s�*}�Ǔxnf�dX�KT.�4��ͭ���`�s�T��-��[�K�����v��T����ݯ�H�(X��<;��L�=�W_d�).fw*��7Y�k��"�JqBI��S�/ݫ��7�i����4�Wu\$�.�gD\Xw�p=�����^�o%Jow|��� �]�mzrp3!C�K�P�A��ħʼ.P<5֬v�?DNDjr���l۱��s(�&<���w�S�wr����fHJ�Ht��.�g�ҧc��PV�/W>]m[�������Y-g�m֒��5���yx}tz?#+J'�e���X7$W�̗�#��l���R�m-�u��Z�J�MǊI��SC��f�Pɛ8r�:��^��pK����/+�5�e�=�S�#�uƤ�,*����Hp2���/S#��e���e��L�i�_����Q��e_x�X���g+��,_kv=�`����r`�&�{Vy*�f���a�pAo*�q��	�tk�)}��|�;�,�^���H�=��*������w�U��6�Y�c�gV{�a�Xnʳ+�vʮW��P�+��>�F���d�}N�3<e�ߵvgn�� ��P4��u�D�t�I-e�B��h�J��|y��4DV�`�����Gl.�k���h��v��9u^�Q��q�#pl��i�8w4�dR��B�� �ْ�:c�U�
�qޅ�M=Y�����v�����ە���u'�f-��n��6�V�Y����Cd�J�����;�^t��(^�J��۾:���|��> S�ŀ'��Z�ӹb5D:�3��_�k.���,�u{��{&ޯQ��W��e��W�C��
�K*�^�����'s�'�χ�^�3�i[
�xwbS{�eK���xr��k��$�K C��#DzK����,v��!�,�>��}ᾦ3,1q5R5��V�nT �.o��'�p��D�N06t�ZSLk*��uW.��Hf�5>�0t��W�6�<Zr0��ӣ�W��12�Y�P@�Qh
��8�ڝ�X;�vD���5å��W�9�����Kk�{d �xЂ��?Rs����~����:��݈d�d́��kg���;T�畠�γ�KM�p�ߢ�阐�i�}�ŕް�{+C�'ͱl��꣌�xO�Lo�T+�*�M|ۭß�F,�&Dd�v���,Eg������ӥ��B2�_���X���9�q{����D=��%�{�����)m=Y�K�F�vKr�A��ǎ�5+@�����r�Y�`�{)�����s7m�����52��[*g�|鹱XN⇼�ӥN*Lډ�4���_C�9�^}������OZ�{)�u��K7L���P{CwVG�x,{��f���_k�PBu}_UW�T��٬�����򼾀*�8<�|+> T�m��.�nqmb��̲3��m~)��3������h�|����oF2W�� =?����U��0.3Ʒ����y�+גD}B��̮���`�ڷ%z�|�C�k׉��k��:��{,�ZϦ�HW`�i�[�3a�ۢ�p��ӿ5�.=@�-ք*���2���T�ϡ�����Wɓ�e}1�١��z�WY�0�/'���t�z�EV#�Nϕx7��2�7^�?vW�t�^��t~�{,������b�+�æw����K�{�|m�1y.9� y�4�Ma��ߓ�})�PoT^�S&�V�A>��)�ۜ�h���t��t��^�R� 45�B�
N�"��R���M�s�ni�Fۿ�!Zr�"Y��d��XڈD �K^��������s��U����V����8���=�����|Ul?ev�*S$����3+>Ws����yTY)�.1��k�լ�gyu���*-��Ct݌��!}�~9�b���x�-�U�P���
��0Tg� fbzy���ٽ)��5�����9t�����V����0K�um
��*'.�~����2ǝ>�������ݨ��W;�AMe�\��6�"�Ηj�2*�ڊ�릥�N�1D��������}싽�7}�~)w+/P�=h��C�}�Ok���{3�w�x��!�=�'�'�{������߂��f+)��cJ�ض=��w��K�Ϝ_�K�2^� F�d�w�����
�-i���n���[�^-,Ǟ~(��������2�]T}\������ힿ��P�瞔�|)���H����3,��l+��cB�8�ߚ�jM�g(sH�w�������)2����+�~k�������y��O���@�,��W�^��4�c{M�I�k*<�������[�s��
[�9�Nr�Ś�usw�h����6<����&�[/���5�š�jq���r���?fC���[z����7���z��~t��-��l��.}�=l�i�9b���u}���H��y��䱚�i_i���BY�躑�,WѾ�����Yp*X��R��#$�����s׮���l�/�):]�Y�͋�NFh�lO�e+y�b.eL�]�0.b{�Q������ܰI)]_X#�&5;3,��vk[n�g�q�Ǵ�W�fXr�Y�[F�Jڅ
��&��Y-֧B�!c�v[	��e�\��#��P�PU����$���M�Y�%��f1ӵ
D;�sY�c���so�h�XT4�����$�m,�ѱ��a=��U��c"�1��%5/.�jr��1m�wo�[��A�
Y��U�a�!c�xLyyn�m^|�N�"�A��&�T�Zُ��R�幊�ٴe���q�����
�|���EG��Y�*�����Ԋ�Q��u�1}�`#��h\��������*ִ�j'�{�{����-�˨�P�e�Ӝ�㼸W��6�vnR2�W���b�K�����,B&.�X��+�=��_[�UÏM9�/n3/ ���m[�棝A� KX��,�X&�Wn���sj�G��'z���%v^
����a�4tMȍo�U�ej�ڥ:��;iV��&'#�	��芶]���S*E+]�Y˚ʝY��>[���8�gS�%��Fy�N��*��tCx��A�^�⾷H���d�꿴�b��������s�( �@�Z�`�mR�jeN�%S>k��wvwN�Xޱzc�CMt�e�d���bZ��c-��T.	c����J�1uD��=�����\d�F/"����.�<�KsX.DŇ�[�V:U�3��e97M��J�x�vP�.��MvtȜ���X�u��[fU���Ӝ�fϻ-��r�����-Sq������e�G��vO�1��>���zos���֒������`Ԝ��l��U��Ca�%�����h�J��-�x�U;��yY}��=w��
��kg\f\0,U����E�4V�V���sqCv�z,�qB�im��^Ѻ!�[ĳq�݆�<]����-��nٶ� ����,.3y9e�q�lY/t�%km-��}�RJJv\�};��wm�6j'*������v��eF�=+W�.�rx�8e�\�
�@���Hx��gi�ǣ�qj��	.�.PI�h*嗗L�Oo}o���6�Ĥ��ZPM��Wݶ�����垩1n܄��8���B^Ou�j!��]��\���J싥wq����<�X`�J�=��ӅI��@fp��P5�gIWhV����Y�h|j�;���R]���1:m>|�u���%�t���R-�4�6�h��^5z5S <jV��`�R.�:G�j�ڴ�c��
��K�q7J�jt��W-�⻲`g�����r&`��>*j���o(]pUjV3���G��J)�:��'����.���)�ͤ��V ��B����N�t�9�Z0��;E^Tu�r��ر��۰�L���thNn�Xgk{��}���d����E�ҡ*"���M4�	�RD���&����"M��أF��Q�-r�lm�`$��ѱ&������b6,h�шԘ�Y1���\)��V2E����+\��Q��lA�Dc)lF5�dm��E�ɰ��A���"61mE!�Q��V-�"5\�Dh,��n�ƹp�,Ti)6���RV�%$X�%i1b��QA���-��F�W�}_������Zf�z\?,����W��a�.�����g��G�Z��aW=os s��@-��F��<U�om��6�j��������o�g����S-�bݓ{��u�YM����C���3�"�U�u��X���C�X^��"w�[�;M[�ye^�k'g@�+f��ݳ��sX�X)q>�U�)X����y^�C��3�g�Go���+�,��l��fZ�pͯPR��ߚ=��_M��!�k.#�TE�Y9�����^�Ė[�S� ��x?�.����;Ǐ,��ws��Se�8�%�ᘋ��G�����_�{LB|�U ���bs�o�F���9���� )�Kk�3�N���n	�^K�iL�[���kɩX�qh;>����d�O��H�q�[V���M[/C�hbo�Ni�,�F����c��3���I����pg�'��:����z7{�7��3�!�h�,yky���s�ٳ|Y��Y�����'b�`�Bn1�4�T)ٝ����p�*r�׀��آ[�⤳���*�vɄ�v�=9v$�m���lC��f*�s:�5��;�r��Ac�b�L�9<�q�4U�ve\��hk��++��GYR�Ұ,j;�qbԍ1] ���ue�8 t��ݿ��}��}���Dy_{��^�����D����ߩr�������^���qx��]��m@=���Z��V���3�En�~�B����|�dl�A��}���Z���jB���NT嬙L���]L�K��y�֮���ۛ��~6u�'��Pk��3���O���-��}�z!�梱��^m�k"���f�5�8lt�~~%�|�{[���}2ݪ쨟��K4��5�˺�}LEq.�@󍯼TO۫[�;m[�̿��������&2��6��O���=����/j\j��KV1���I�i�ä�4�{7D���è3�~��L�m�w��:��>z�$��L�J����`[v=�iq��mX˷3-��m`K��Ӱ����LQ�K ��үH��߳�o�/ר7��E�.��Xe���O}��oE�7M���ڦ ��Lײ��>��g��½J󌢫��cF}��)ϊʫkA��O��L��MS��eo��6�hp��Zd�j�%�*�]�G��77�iC�l
�X�I��(qT�5�K��J�r��Q"Om��e_J[Pl��!yi��L��Ix���*b-�5۹��\ˬ�)M[�������f�OӍ�����)��6�=�
��Q.������d@�ڕi��>���7�ĩ���a�凓�
�SJ�f�@y�P��T9�5HV��V�[�1�g��N6��E�NJ˼�	���	-g[z;a��)���F�WK=��܇}Gv_�����3�k���[6��Q8�rz���\�����w�OZ���{���(�N>�/υvX=ܹ�6m�,��}�g"��!�7~N���R�5��������~��V��U�۞Ks��U��N-y��[��Q����^^�Ǧy�����^[�}���XK�Zʳ�iww����'C��Daɏgu>$���񙜬�����=�������b���sE�t��9뇫16屾q�׬#�5K��7��~�(��L>ຉl�f���W�I���:^�W����/�ߟ�.v��i��q���u)D5�K�kt�`����p�/`/~A=�p�|��+���hi��.򯰥^��|6oz :��!��7l���>�ش}����}�qnЏh����hϥ��\i�������}���|��,��ۇm<��_ >7�T����䟱������E�Q腟5�#U�炶
+}~�fs���x'f�Zi�זU�|��w�����.!e�w�l�N�^C��5y)�k�Wp�7���x�~
�c�v}T�
��{z�o�#rc(]�۷��{^<�h�u��l)Ջ����>p}�ynN^��sWO��Y�B��9OZ���C�}�xk�z�����Vk4�D�b��*|q���&0���Of�ɨ�m�}��lo���Пi-u��^�=��ә;_F��F������ʊG�����5�r�:��f��pX�P��m�p�9�R�ik�S�X�o���䷤=W30m��4Z��)�[F�$Æ��
��\KV�i{C.`����i_��������a���9���U5�1�z���}�����+9�{���ΛӋɵ\p��4�T�C+�,v��EX?��F=�gj�v�L��6A[>���:Vc��(�(a��놵
g�P�.�8��X-�
&��&�vQr�j��)q�{��AR3|��$9[h�V]�-1����/��Jn�H�s�P�ԇ��o�ﾏ�&�����ѥ+������t�VL��.�;���^����aB�e���f�N"�Z��'�8��{ȟ�eҞ�կ�;��W����R�tr��U���5���ٝ��t������j������>�N��	�&�P�Na��vt�I^�{1�ߗ��yZ[��_��������6�y��u��~^A��Qj[k�K������Y;5r1ƭ��Ad*R��7�5�ٯ�(�n��Q?F��r�=Q��z��m:�f>x��f�i�X����9q&�\'K%+��<��<_:O.ޫeZl˦��<��o<�Lݶ�
pn��u%:���\+�7�����\y��>����V�>>����Cڛ}]���xSuu��\�L�h����ܫI��lX-�g{�>��=�~�%�p��_j�(���l,����:�,#�Dx=/m��C�]rF����G�²� PM��]�g`��(c��2:?3�<;�chE����5B���IV�B��v����˭܉�-��Z�Bۣ�kz��Ƿ�bc�VU3'��^h�v��E�]�Io5U}���^�,�'�0�����	�
�lx�gЦJߖ��05��J��ʠ��OE�wύ���Ɛ�o��M+e�p��7�f\�
�k�"4(Kz��X!�7ȷ�<�
K�}oޟjϷ4*�Z�6�;�;���Nؠ��2�v�� ��e>
�o�R������f�F�&|��vٰ�C.�p�lƼ���iV��C���������"C���Y_G��I�|�^�X�2�)E|o��w`����u�!Y�����>�z	7�'��._p�/>Nkm�W�����ˇ�0�ܣ��ZZ=2�������$��g�A�-��^y9��q庯�~	<j#��zE�/%���}��;�$'{�w��{8��L����Ml�t����/��{�ܯvk��Z���Bŵ'`��}�Z �������o�_i������y>��.�w�v�6�9N[ӫ2���˖�;AJT:�=&�۳��/b�]���j(�^�zes0`T��f����/v�Y��>�Z���s}N�0��MJ��i�]]���I6_D��F���%۸�ʻH!�2�Y�Z�IJ�+�m7s��{c�ce���U}Zkg��d�z�ۓ�^$��qT��*5R�j�8�����w���/*^�K<|�mFUw��F�����{~'T�
��h]�̙r�ӛ�|�&Dy˵X�b22����R\
��М<�m<
�ў*�h
~9膗��m#Hg����>O<�'=.����5���ڋz=M�w,�_j��A	C��B/Y�~�wN����mE�9/��0��k���������H�K_=�:l.���qXE�U���3�{�,V���,��`U����x߾<*~���90��v��Lߨp��gpcr���j%g�a9��Ik-�@~a�{3Z�Ԯ�#�n���m�Oc���|�F:B�;��^^��j�?8i�S��Vؤ=B\&�6Ѹ�qq1���{_�+}�ͫw�{C��3�J��������@Ox^��y��
v+g![�_�A�V"�;���e��e����r�h��qT���6�e"fN�-���7ij4���k�<Sa�+:�-�v��V^܋�];�(u�pQZ���eN-�;�C��m�!!���N�ݳ����A�M;#�݃�p�|EZ�I���m��ղ�����}�������n�!/W���v^Z�_�ϓ>Q��%��g�}L��_��X�����{
c��ޕ�_���ӽ=�=�Uy���y���o�W��i�oà����p��7�+^5�S�/�/�}�unL�sV��j#z��}�6}�x�����Xsj�z���1�0ߟ��nu����k���O�b>'�����K��f܌qʰ�k��Bځ�z�!߱�F/���)���ZS�M=��k�*��Y.���~V�	-b�{`㬨}�=�T���
9Gv<�s�߯��|�yjoU��,�������^D+��;��~��q^+^��R����_�p���7M�QC`���Z�Gje�/;������C�ԕ�� ��h���q�l{�ض�o<!nz[�k�q욗ܗ[���B_b{8o��SJ�ƒ�"=
�V�'Σ1zT�C4������IwP�*���Q��XX�\f3�*�CA�Q����zZ6P�4:���,�ﬀ�m���Z�ޜ �Mu����Ŏ*+Uf�v�t�Z�-]Zܦ�����*������v���v8(��nn�x(�j#�_W�U�o���X�b��b~��>H�C��C}��zW���������Ry�{t{%I8Ai'�[
��	��'nh�f��!m@ʒ��J�K�����1��Y5��jC}��kd��&�w�ħ[:��R�J[�#b/�an_������Y�,��֒����yF�=���Oޜ��1>O�{������s�Kڬ�nE�_,�V��s텎�K�&|������6��׽��j��9暈u�����y�B�֡�٫_��)ޥ�Y�z�
x��{�uR#}���z�+�w�o��P��J+t��Z��a�钱:�w��w �s�{����I�\߶���~�i_i�Nڬ8�����;�I����4��{!���E�=Y�ٯyͥ�y�nM�q���51��]P�s�:[�g�}[q�·��{�.���^\{_&�v��rb���s;s���Åע��׀�5����+�V
oP-�t������ݥ���pte���7�~�ҖP�'�h���ay�.�l? �R��}.���#m�nPr�c����*�C�&���~���Q�<ҩ[�}�������N\z����F�Y)\n��o�i�t�#Z������'�h��~��5>8�`?��z�JU%�W&~��ކ���P�HͿ9?%Ml���߷77��Yu��T��07D���F�E2�2=�7a:v���eg�Yɵ�<�k]��\������)���p� +5��Xs!�+e��T�P������Zi����=�V��DK�iL��-�F�� ��s-ߣ�AFS�]Z��}V�+����L���	�E9�5K5Bӧ�*��dEvnU��{�Õz�'��K�?nhU�j�k�އ��p�1ZT0j�,<�~��9z\2���+=5)�|�ُ��Ԩ�LM�=5!�b%3���)��o3ӎ���)�@�u��r�����2���Ol�aCo����/P�+�)�V�W��6�@�� .�^�Hc;�R�u{���-�ɪ�`�[����.����7V@�ύ:��q) �
�����6��mݫ�(V��:��Υ�aG�3�ړ�㼣����S�;�VF�Z���Fӡq�;�)^-L����y��_6���'NB�C�ހ�;���<<�x�]Z�ua���eA�eCZ컘�TPݓ{W|��&GoG&D����U�f`�W����s����ׄ���luV��o��U��/mJ5��l�`?Nn��<j%h�������2���#��w3���4�8��pʳpD�IX���[]�o�S��8�L(�����պ��%-9S:𩚫	n
�uƞ�^�v��T���v8
u��}�%+�ã��%ʅQ� ڷCV�q����Wܒ��j��{�
�q�Y�����!�X��f�ɲs�l+ʾ����rr�B�	��؃x�ʦ�[�a;GU�B�����"���E�_A��v� x�R��{T�5rVo��%S��k-���DW�%�TH�1Ԇ��sn+��\p��.)�0�����2���+��*�>�����Ճ9R3b���*]����f����Sᣛ�<���K�#q2���۰�)'�`/d��#��x�Ezh���թE\�Z/쪊���փW��u\�_>��|c��v)��+;e�%�*�]湋��*��w�>�B���	��ob8Sմ�CJ�0�uV�p��Q	9��fsw���Z��r�6�丅!š�YR�Jt��I�)A�/������4�VtU����nt����ïLoAv�u����[(�.��k��1��DgR�T-���|����r$��̽D-��2I�6u]ټ��{�e%w;R%N�LXsSFb�Z535oL���L@���Av�(����s^$�-)��5�en-������!](AQ�e��O��C9�Kn��������D=�!��<"�������]iXbY间�y��j�HN�Q�E��sDe0e@tjqvf�(i�7G;��%)or(욨s2���c���;쳮��/z�u�x��q��w5����^�&T�\G��t���䋺�kDPZɴ�+�n�Ƞ{�.�xBZꍲ]�׺��a��\Vs�ӛz;��B�R���56�Ȟ��u�CB���E��Q�}���	�����]��}��e�O�̰J���샋�3˅�ʺ��-#�7+V[����4k%N���Y�YS!B�/(�8�.M�g1f]>�"��/3T�8X����PR������K��lk(��fݮ�*Cp���Ċ�M�ɨڍ	[�ƾ���ޓ%��2�{j%��ic�����ժ��QJ�u�p�_V8ụ{#X��Y��6��������H�!�Z���9j�z�m��i��j�xSAң�\P�o���Z�W���-�'�Q�#y���q���S�n��q�wy�8?��ܹ�L���l��#���A\��,D��$QQss�(����\�X�h�N�cQcIh�CѐЅ��F69�(�F�E���X�Gwj-2�Q�m c@�&cXؓr���m1X�wVK������';d4�j1j5�nW,o�b�"�W7Mx���h���wr�r����5sn2�x��ܮE�nh֋!X�p�h��W5%���I4�(�.�[��\4r�Ar*�`�us_�
����MK�ky��1žX�r�i��[�5�j+b\<�������.żWW'I�.�Z�T��٩9x5:�l�����/Q�c}\�V�_�����c�v�\�Ð�ܬp.���=��x�K���j��376\e.�k��r��?u?g��fR�X��*�Nt(ʒ�+���徣ȍ9l�3��==F�<����)�dhi������r��l���}.v���q�*7V�*���[�Mmɉ:�!F-	Mfe4�%]h0^�8�Kڕ��c�^	;^�Ұ��T2ןs8�S���8�qgM�s^qYm�9����g�[cH����g��4�ǜ<����+���K@CуtHiG�ME�n�&oX�q�o���7��}��?R�G�׽���|��9`𶫫,�o8o���{τ]^��Z�?_<��4wHxF��ޟ1�t�d�6�2��V}2أ����W��(��D��w�Y;�
�4��o�xUw�tl�e��~x�#��I���e�E̯e�k��v:��3J��|4�j�Nգ���Y.��X��3E"�-̛�#�8�BT��i� ��(W<�,��0�=p��zL�,�N���+� n_)�r��=�MiUh�z��@c���T��ྙ��w�`�ү�c�#������U��)��p�!���V{�9�}�RZ�CoC��1�d*ggϐk�}���}��8z�q��/��ڝ�>yy2�T�4npJ�8�Ww���Fe���5	�ƅG��ƺs�/6]�Egyf|�8#�^�4�}�Vw�u{����w��EyÔ�8j}_C�q������m)^l����~�w��O�{���z�_۲��c�5�Nr�9�ws^�p�n�E�,���X�{�+[�g˽��񙜮w���b�'�����o���5�WX�����Emo��R3�ƨvOQ���~y����<�{��yw����홷���Fe����\k�;����y�OV]���x��\8s�T�{>oʾ�5��Cw>*�b!�D�[v�������˟1�e@��1��[�M=��Z�ʽ��K��6`���w,Wx��>ہ݅9�j�g�OOn9c�����)?L���pr�/[�r�b`��n�ɖt�}`�@kr�g^�<��;C�5 �v��LrL$��w:�;�Zx	��s0��mw�R��gN6F �;L���N�]�66�w�p��_vq��r�1�����I�n3O�=3���[�x�����?�ƭ��].��7�9����{Q�xf�~���Q%k�V�(�m���ޏSt����z0	ʙ���8��{�������O���+3z�����^z熽����E'ټ2o�eo��Z�d��p����za�q7�w��u�+�Qݔ�<X�^��o��p���4(q��.�\��lb=���2 ��)������k��������Y����AR�ii��ض��X�,c���Qag��o4,�[F����4*'[5��<�ۦ��s��gf�����gyf�����i*��N���c����\H��x�ȟ=Ֆ-xj�x�-��U�◓|��i�R{Y���پ[�b'6�������Un9˵w��b�����ΩO[]b�^�;yҾ:�dXsm�X�e��O�J�Ҳc]M��m�V�1|�kl�>��F�Z��b{��Z�m]��o��3P�޾�dA��f"HA�!R�2����&^���2���J���|�Ӧ�nͽ�H+�@�*y�"t'T���+�kH��.��4���;�[
*��w��ﾌC�e�5nB���D7(��z�[�k�{÷��FϽ;���K[C��N���8��5�ݙ:�vy��	r^�^K����5�ʰ�yqy���]����޻��<gGH�?}�3�K��9�/sɛr_n`�YԶ*X�O,S��d��yz��4+o�+`{�s�==o���=6�I��颩��Q���`S��� ���^�K�K
Q����߯�8k��`��4 ͜@�q�}jg��6c���7AQ	zKԨ�^�oC^���^�9y_�ˣ�%��kw���~Sm��*�ڧ�~�`4�$�v�zB�X����UM�'���{�z'�S|�D�J�;-}�G�>	D�׳p�����{��30��df ��b���͸)�l�<O<)�o�t�B�*�ߖȌ�kf�W����n��y87]߅�}�+��ި���>e�w�~A7q�i�,�DdMi��z���K�2y"H��B���hN���5=՗qs86��N��]j�eۊ";en�.n�"Z��l�4zujnz瘡��M(�g�M�a>;�;A?mٓoU�70s}�:V��\�m��	�+b1ޱ$8QF3�%:3sOj���+//�"�D}�0)1�:�T/� }m9�Y鯣��hZ������؄n���Z֎�%���hO�(���� �"+vٞ�ѳo��1Ȋ$���g����f��~�5���=�z����L����ou\�Zf��=�m�/=Nw�*�i��%U��(sP���Bs緣?U̳�m.EVr��U���ۜJ�k�X�p��S�;6�&�S�6`�r�']��{fi�1�Q�j>q���5�D���W��Z����L�md�~��y�O�j�X�r����oFK���^{��j*��nZ^Q�Z=�׮/�/�[��k$�}�unF��ˆusQc��m��x��q.v�T=�q��cuks�v�w������O-N�����_y�������(�@Y�W�A�r{�����Wp�.�ӃC��~s�<�� 3��䧠j9D{y�;�佼��[^�:��Y�S�o�ir���5ݬb�që���Ęz��nY��Ҥ_fԹ��0�{�IK��WR�k�Y+1d*���@�(�W]�p�]����\]n��X�(�"��I���8R��S�H(�|��ꬊ��D��s�s�dngV�Q2��pE���T�[�;��?H��CV��T6�Y^n����E�{��k:��T��S�Y%��/�L����k}�=��z���(�_j�
�z��L�tǱ�؟W��eY^��<�/<�ݻh���'�*-�ꈗHο �nI����9��V9	O�/��0�q0�������f�@y�Y5�y)�,�c��CsNh�Q#��F��D�������H�R�{{��i�VƯ7O1�������F�S�* �f������ϥ���iJ���D����
ͥ�=6�jLM|یw�N8���v�o�Ohe����$��^Ng�Lt��<;�ߚ���W�����5�nT5>����p7�,>�h	BD��k�m^�7���痍f�<d�3�����b}�{��X{nP��r�U�N4Nd,�@N cځ�:����]���Ť�����˜ˬХ�� %�,4���d:�>|e�+��6�ӝb)���E·�����ㆉ��[��:
s�x6��J�>S,�S�|�a��Y����8(:�G��Ҙ�/S5�f�Ru2�;ѩ�>gs�.�>�tT�Zu��oZ2H�Y�G��woe���}��>������o�Wy,G�-9W˷�8�잹�����=ED��Y}3�_E�$0A=.$��-���9�ku�G��^��46 ��ʇ�gy����9��{�j�G��p`�x"�v}�lC}:�|�����=�Ϙ���V3]��r��,���ծ������=s��U�|��w�l��y.�%W��Yx^�-���eL���W)F7O��^�O.ޫ�e�u��&�ѷ����C�� ��u����;���J)�4��r�Z�F�B����ڗ���ai��x�AW�_Y��{֌��^�o,�~n�Jn����E{��mW%�Bzϐ�9C�H,WO;Ϫu���f��J�;6�p�Q��0���m5�<b��T�L�[!m@�05앎�͛n~*Nؽ�Đ̷Hm%�[/C���	��Og�~)��W&u��~A|(�|ORzu�i��%<25�ϲ��R���ggKB\�Tl��I�9u-Q�����RE���*<6�т�V�Yurm�P���뾫-�'{�rl/ �Y1M�z��W��r5;+���
TЫ��̍�f	i��kA���]��S+f�KfY��o N]�_�m}��:��|L;��c�F�8��jف+$J���QN�
�@��-��;����ۏ��U5i�5	��aMଉ�rE�z�)��~�.�R��:�{���7P7݀tY�O���?W��~��}�v;�{^ܞ�Fj˷�z���
c<�V�B��g�޹��P17P2��Pr��ƅ*8����c��r���T>�.�w���{����xzdS�9��@:X|����?��q���~��������߶���yZ[�9^s����OQ�<��t̋ζ��46E���\"��.�-����d��X���GJ�V�xXy��yy�*{�9�/�+��
���[��޽�OL�������RZ��a�/��[��`y�^�@:�KңVB�J�cv�7k�=E�U��f�ąW�����1[sz�Yt���~Q�H�ztEM�xe�%BI�C�q{iYZ�IJ��ۮq^���ߋ$L����Y�i�;,�f�J�����\�b^�8u*��v�>�*�eI�%��B0���_0��_�H"` ��J�"jm�0�(�x���5Yw[��we�m�")>V�k�XoV���kV\9��e�K�C"��*�N�z�=����Ϩ�m�Ş���{��*�q�~f�]%e���@K�x��O��Q�:Z�g����S�m%�<�'�*���Lҙ*�ߖ�˵+%[;r#s�4��Y»���7뀶w����^�a�
�M�)�9�:�0$y���ߩ�;�^���
;ח;m}����N6i������=�t��i��5~^̼�\�ѩد���)��sY��嚹ew{c���R��e�3,y��'J�W��9�/<��=s/4+��[�3\ڽb���bbk�\-����֫8w>��yO^��XWxS�dhV�W��z꒣x�Q����f�<j��3K�c���ׅ:��8n �v�
�VF�͙<����y��ͭ_o���Lwsk��~NS�Z�V&��{1���$c\ u`�+��gjF�A�	���stOf`t�z(�kW������)�Pֳi����ف�[�p�L�=�P���w�5%�R\ldj�����ma���̽$�������_)�<���)�6]eh�pe�J�M���6�������E�X��T����ƥ�e�+_����穡��]/D�����U^�`�����7rv�OU,��3�6ϫ��x鸶��Xpx=�����L�~�����|2�bm<R瘓����o��^����_J�����V���{�x�b�+��43�g��;p�h&�O:O/�*��nJ��4dT�Ym�������o�ǣ��y�'gq;�z�ǜ<��O��x�Z8s75��v�ũ��羽��>�������Z�������ޏ7-�����q�f��-$T9��)���+xX�O;ς��|�h���=���*��^�y'a0.����oL^�����?}C���^j���`U�V��uC�Y�Ǣ��a����$����Դe�N�5�5<���O}����5�.n�4�{��4�W�~a�#q)�U�ZB�RS�mg��Uw�q��4�;�P�������l�3�K%]̺G����G6]H��r�h�؃�������.����ӭ��D��C�7�X����^�v��w����k�멕zY��hب���n�W��ϸ#Rdv�فb�*�Ʃ�qT3F�Z���85j�li�Oƅ.����c�$!p��!K�W���SQj�eѣ��V�X�1]M�;+0ueH�Õb�.&���X<4|�@�:�1�.W
�l���_6�%`$��7]��ao0�Aݮ�b�}Z��n ��EQ�[w"�xEh�A��c�Gp�絊f����-�U�Kk�`m�t
m��^r�kC�Y:�xl�EuX���jb�z����%�7��%�Qd������~�[��>f����h�b����z�R�nr	��x��=� ���د	t'o �֤�G�F�}o���e�j�-N{�xͭj�.�����N�\-�q� �{�^�yL#h�Xy+�o�4�l�zS�jso���u��߷FW"�4�+Z�ܯ8IB��:�M��\�@],n� �;ѵ�l����;�uΝ�6AW���&���?`g_eަ���Jh��*޽��pm�]Wb�eB�l��3���3-�ށ}�L��(�+�DkPr�V��&�����a�3�����[XtK(�4[:���#Fn�kGH��k/3.�K�.��]``ⳇd�;��6��F$mU�foX��+���B��XR5�3��(O�כwN�B-�C ^
�������(t��u�2Fr<� '��Ա��a�Ղ�\Hm3jْc��fw\�Sa�JWU*ד/^j��~�B�B-%W"{AZm�-�0a-�㋌�+��.���z�縮=V;����ИZ��w�G��x��ǵ��țw1�R�$+�:\ �ttK�F2��C�+:���M��\/g]i��F�2N��^^.�-\n��l>ѳDN�R������h� �ΊS�/&�hG�f}'|���Лx�2�3w���Q��W���7��2G��3��A��(��\g*�n��zF�]�ҼGKV����4��#Aj��*ɽ����ɛ���ɗ;�ם�R��d���`�$�t>Pӊ��Ut;]M�Wĸ���5d���'
�3��;e-�/L� ���1eyԭ���x�s�X�V�s�u�r�җf���-m���6Br��u��eC$Eh�r;"mr�3o3Z���ǓS1C�x���x�5m̷�tP�n�7�-U�]\X:��xI��B�cu�=�t��E):���ݛ.�8�5�X6�ʪ*[r��#��V��[SzV����Ga��5�JI��'�z��dȌ-�{�%�ԩ��3Lub뫐�RbԳT^Z:���Jڽ��>��e�@�[hN�Vk�lh�v��C�b����tGq��ug=��V<v����i�s�啴�i��!���o�_������^�?���k�ь�b�QF�Rm*��H�EF���-s\Ѱ��j#cwv�C'��l�FMQ�RlHX�h����mcX�h��sa4V/��ɣE��1�#E��X���-�"�.k����E�Y��(��/;Wyں	���Ɋ�6�F6$��;Q�����Ur*+���/�b��H���W9�ر�j��񹊌V/��O�EQW��,�$�y�9��X޺П\y�K���z'�漶��@��±�Opd�6Z�����SJ����d�Թ��q�/u�~�M4�`�6��#q8��]9���s�v}bӷ^����ǆl��.M��oϖ;��EyÝ�����EG���Wf���j���|���VF�n�s}�:j�Q���8sO��-9��/7�瘶�!=��;��֭��	��b��%�y;�Ʀg+����gd�&_��w��Lx��^��kg%��V��9~]�����]G^�M��r����4���W���R�����WÍ[������&�%�S�"�3�ac��*����T}=H��T�-�/5�١��U�@8�R�5�Όik�V�Q�q�Jہ��E�M<�>^f����w��N�ȱ��9���{S+]¹J�cwo~�x&��ެE4�F���VHr�Z>8� �E|����jצ���^^p�߲0�?'�^%n��Y��Wp�Y~�cw�Vc��(�}��l���a�>�W����*��;����#2���g7����Kۮ�	�r�p5�*gX�.���'i�f	��PP����Pɇ��oa4��ԋ���]�z^>�G�<Y����ȣ{v��+Z�a{����kك�:���}�N|��,�J�e?Z26�!՝��+�Zkڣ\5��Ok잭^JZ�|��9dq�]<�,�{JǪ��)ormS�*�\����j�gɱ���9D���hF�g~�xbe'>��+��������z;a1P�N��,��B�Ճ*�O=t��6�/{+V_����l��΢ƍ|�a�q��' :���w}ٓOO���`�x{�����9�Y��d~�IL�Zp�Bn1�ҝ�˪�v��y5��{�k�؊�y��Y�9y����Ց�^�Pyv�(-r�W8pߧ������F�w�;��U���Z��<�K��+�]zs����\��v�\��^>�\.��T����n}+ڭp�q�&n�5�.2������gTZ������kҗ��yZ[C��8�!���I����k��U�83-�ܥ��}��o"�2�1���u��z���aD�z���F3�TE�-,U�W����;+�Vf{c;���r"gֶ���է�.�R��|,ݲ����\G�v�/���-)A(�ռ@��1k�Bt��)���^�6�(�[��M^��_J��qZ�o�^�E��׼��5�ڙ�	a�U�g����"\�������6|^߄hVߞ}[��޽��y?sMm8�s[c����fS��%]h?�5\��*5,)ln��}c}��hn�LGr���}�d�^8��gS���r�*�̋�g�g�,�X�-zz�u^���p�0��h'�p���e���(�_o`t.Kϯ�ݥ�'ag��W�J^��V�צ�{��/5���~g�.��캅�GO%}S�7j�y̅���^T���i\3x�<��lz��5�)���f�e/d�(�1,��|���=���������2�;�T&���T�܋�M��8���Ǯ���ah@�9�%ގ_:�<7���"�[�<G^Ò�Z^��#{U�w�HTl�F��m�k6���ir������«Nozn��'���U���y��b���g�zK�b���]�[�R��5UN���{q��&Mk���os\%E��]A�sl�S��u�ǭ)"�B�f��M�]��v�;�{v�0����\��_b�p�]�����G�P�>ȩ2�(s�a\��:�����)7���q:�ʸ�Ohe���J���޳xvC��M���:�q��Z�i��z�:��Ldz+vuC��ɂ��S��R�x\��������w�϶xw��{!����~�괫v��΍�6=�ڌ��n�M����z��ͼW�+�������{�d�'���
j��7Z�+�^mn��u��yz�z�` =�Tz�o�lc޺a=��{*�w�&�����X(�W�h\hV�44��=w����lu�����)�S:�=�������ӭ�N��1�����py�4�]1Aa����'xz�2�T;)}�w	��S��{K7%\V��"�=Ws�7Κ�!�xG��Ƿ���f7��s�~X߯硯\G�<�m<���e���!	�f��YW��~�jqCb`{΢$�w
צ�����kq����z����fBy"M�I
�hT��7�b�Ɠ�u����V-���r����f %�3��/$|wz�N�QX�4C���Ŝ�NNz7�ڞ'<��2�~�.`��[���[F2̴��ѓ~˗�C"a@+�%�*߮dQ��m�#��r�F��ӷ�ZSl�wo:w`}/��������|����u��5j�n��I�*Sy�ڝ�m���y�}�y�����P^j�,��Q�OK�i8�h܅��� c�Q1�W�<�O�Ni�D-!f�#Of�g�q={��o�8o0)�HX��f�z�~a�#p�1�3�3Q�� �����U���eS�)B���m�~X­[E$�ߛq�
�c�K}<�P~ո�QAv]�{ݝ�����\������Z��SV�3Pہ���k����{���ٳ�}�}��m.EVr�4�f�<d�3����-�3���ϴbO7���˵w����b����}[��4.mj=kWL ��R�'��}d�q���������f����K6J�Ƽ�aŹ=siu:2ֹ%a����>򷫗����g�E^��8���im9@�5Y�:����tr�y��:�� ���1��{�rz{8U�4��1��6pmy��@��߯���.�S�K�f�G����A���,.i
%\�:M�x�7^�ѿ/ Q��m��IʖN)+����m�9D�5�-�����\V�+#��\d��p��g{��63<u�Xo���E����-��x�n�W�V�-�-�Ǯ�n�%��˓~�p�<^���&#|�si��u�~*��Y.4�W���gήp��n�����P7�H�\�Ԩ�n�<��~�M<�9��V�9_	ʑ�EJ�^̽a�U���~UIJ�N뿕�M)O��1K���9�rv.�2q��u����ev>r�uH�sG�������}���U���ecS;�v�l�������;���+�w��E]��2���0�=7κ/o�m�ҿ��k���lz��9�2UG�!k�V1F�(h��d�{�ļ�~�T;g��P��2�;�?0�!��N��,�H�v˯Mg�8_�-�
��*\���m����AƊ�z��W�;�!ϴ]:��n?ml�ee�$Z}��
�;w�m��m���$�����=p���C$c�V�Q��rȔ:�B�������:an�c��)���S�cU�#����C��+,T�u�s��Q��vv�Fl$B֗o[;�ˡ�{��C��	Ś�5���c�q���K�1�7��*��Au/1a�%���v��4�R�~��Q�P>�S�{�d��߯�v��S��U{�mEg/3��7����Q$�T�
�>�^��g6%�ڽ}��ʷ�g�j���:S��]b�"���mzAu{J^��}�N`.�����s��=_>�Z��Dف�/{��E���-��=�LjJ�s�\u���{��:�g����l�5�䱚�i���)n�(m�~�C^w���s���[^�V��^��׮/�-��w�ߴ7�vl����=Z�X��Qc��oG�[��Mή�k=Zꋧ����{��+�f����(k��;�/�s�m��S��2ϙ���ƭ��l�.��l�}S��s�ܼ^&�ۤ��ި�+�� ����Γ}x��[�\#����{Z3=��^���ִ5��*ެ�6�e�Ġ�n���wsMf_���5):�K��^�N�>)o���F8��3y��J����m�e�O�k�i�[E�^����̹�I����n
��t���Юfu��-�h!�lw��Vu�t�9iu[�+c��_9me"aw�e̳����E�e�n����
ڍg\��Z�i(�Y`^Pg\���o� R��+������f�S����� <��<a����<�'�+�lx�f�ʛ�y���u�CS�?�Ȍ?y5���-���F���2�;�? �g�����G'f�M�QW-��<�KG�♯?�N�����Cg�:�w��g{1e\\�)�=��Br�����,	��@��A��xgm�s�k�]��
�7X�6ȥ��_�m�F����8F��E�����j��j��mdJ��]�V�NK~n����e�q�>��^�ʽ���˅������'>z(�8��Է�(I�����i��5v�����u饺_�\y?�K����nw��gĈ�i����ھ�|<����a���kWP���fr�]ޞ4��q��_��ӎ�Ŧ߫�V#MZZ=�9�^^�����T��5<�b�߮�udi{�Hxp��I{�yHk��^��z��y��\j�������o2���c<ܖM�b��eov�t���ޮɈ2.�����(��L�p�̓*%� ����h�&����u0q�[����Rc�&�E��&��5\l����>U;/*�0���S�ʛU�g��*m�L�+ۣs�틱��:\�=�uE�oUsnv{�{�{cgܻ~^��S�c�G���=e��ӵO��5�l�&�m�'v��W�M4�C����'>�n���<�hb�j���N�y絎|�_�}�-5EN,o���׮<��D6�Y^n���*��2����2}ka_��7xCO�w]�^�R��!�k}�=�g�n��ߜ�D�r�xr�����/�������R���[�u�do9��]���������Z�"s޿֏Wҩ��9-|��J(/5ad�����W��Nͫ{s�O�C{��k��oz׭u��P�*yڹ۲�~J���.r��fxjC3׺3wm�����`Og�3�3Q���uv���K�G_�7��N]�\�lwz�����Sn1���N8��v�v��q[gA�Ɯ�+�êI��'��p{�	����=�>)�4ہ��S�z5����.����B�7r��������u�}^���&�t����׌Ǣ=�\�@/i�r��ٔ�Z�i.ǻlO�Ve*ea�f�O��[��S��2P�Wu�r�)V
X����'#��̵$x��غ�lF�5jf��!���Y;HxO
���+v!su\�wL��/.8r���y^��t����'����%���V�ϥ%Ϋ��r���1��)��)�U0ku�GXz�7�إy��]�����ߗ�'���{0���ӡ~E�N��2���q}�]��5<���+KG�����t�M��o_5d9﯄k`v+|,��0Kq�^�χ��o�[���~-}��T_L;s��������4���_��[����^[���s
^C�H��L*ܝq�2K��_�T�Fd�M�HaFs��'���;eev��������;C��R��7�(���l	<��l�(.;��ˊ�tﰈ��ÛjM�Xp�
�^d4&��M����y�#/��zϤ�r NH�/��@�-��!�~�yw+�;5�ߏ�yV��o�+���9�qZ_�=�de�ճW��<\ �ߦ@��}��������ʞӪB��w˘�.�<���Aػ;q˵�z'�J��ƶ�c�.�Q����oCe.��fF�:�A�k�[y4����X�W�jԢ��}���8��;��}��sz���v�;�6�x�q�b#��C�PR�v�Z0�]�j$޼����Eh��Zn����!kMŊmv�H� ��-kn����c��k8j�LAy
����6�e튭6ֹ�,�c��b��Z
U�u 5�p�w��0t���mnp������vp��7&�ɏ�#��4�mf����7�t���
����������Ծ"Z�CN�\´T���;�e�6��W99�����j�7��P����M��z�<�6]5}+�����Zt���uJ�|v��bK�Av)|���5��R�F��nwwOXZ�2�u>w���4Ekp����W9]4S�ufI+��Ww��i��"�썭׉Y����Wh�b�6*����J���C����G���~}ޝ��E�U�n*s/י�� +��1��ަ�w���T�wS��i�g3��C�mV�y�6m���6c�b�qGV�^������M�V�b	�u�G��Γ���f]$�X]CP�j7:�Տ���,�1*�(#xj�P�x^$������^����77F�DL��+�B���6'���z�˖fJܢ+s8���{�Ʌ�fr��{Fv�$�P`ԥt%���fv��Ў�]�U�1�ڱT�ȃ�F!�5
lb�`�ݦ��n����%UA��%��lj��{i�o#����~����*��P�S���.������Y�L���ʊ>�>�*� �u�7:�]�j;p[J�ǚ5���5I�u�p��M�h̺]v�n��-n�s�!�n���v��^>�"TDڗk�Be�t.�s�C{3W3��Dm�F����n7%�'	#��8����[rl��CК���j�S.��W0�2��挛��Mj����y"R���;YN����R�w���S��t�<
�	�k1_WD:);״����9���]��g8�Y�a�1v�:�u<���d�5�(R�K�������u��"
�#���(���cV��0^���𧝓���,Db<����:��V�o��t�y��E"Oq��7��T��r���Ҡ���Ie��ʭ��<�]�X��v8�{���r�u(+�f�U�j*�����<���!�;tb���3j�P�(�' �o�u�#Hw8ry��lm�{��J��Y��ʖ�ە�qC\�uд� ���)����tMN]ȷtv�©��	����,lҡVx��}o�� %����40!��j�3Q�WY�.�
u�����,�D������n=ܤ;z�Qց r�\�Vp<��bWR*�n�B��R3%2��>�t��Hb|Դ��rKW��q�M�[�j�{��T	c�E�D���4YN��w]���Z�fub���L���a�j�T)�������0?�k����\M�t��E�Fܴh�sW��/:��p�(�˞-��.\�F�M�9k��h��9�k��;���#FW4\�����!��ƈ،X���Ɲ�
�Qt�h�68m]*-�c�#QQҸm�ɚ����#sr�j�;��D��*#�E���9;����M�N��s�[��G]us���k�N��5�wG(��
v����xOz�����<�i�a��t摨��!�|�J5e	t��ɗ��{�6+S�ܶ�M&��Le�N�]�yB��=��_���mh~��ُGO����ӸM���\G]�����T��X5ِ}��9:�I��Vp��zh\Ed���/e�6����g��Nq/�ƣ�+��늩^s�P���7�E�)=�t�X��/k���j�%����a5U#[u���t�ؽy�/:l^��VW�,�q�'P<�dr6w�������\eC�_B�����]���^�Q^ȩ0T5�kU�\O.���懮9\�feda�9>�0�x{➻�WtQ|r��̉���ݵ��G�����{�Q���[��CWH���ޠ
#ǂ�8�xz��*U�gӷ|�l�{�$��e3Qy{qޕ4��}�_mW
�}߯p���s�a��􃓗3�(�������v֕�,��I�>��E{��ǡU'�u׼_�+�c��UaʱX��`6z�nh��Y��]c�_@�G�צ��WH�)���2%r�@�Ϋ���M��rE_��ރ���T߳�C�ۮ>�ωJ��x��v��WU#t��eP� �����' Q�9>;ދ��&U�huunmMO�'i��Y��Sr��n7F���j]��W%j��TL���hG�(�g���|�j]���š̾�����2�;�7�8�0'�w)}�ᘗ)3�Cil��4[[�X`B�Z5w��yeܕ� ��\ښ�p��a�޴�}	�~���#�_=��\�J5%�FUC�3��3p������}JEz�v��~�������}n�o�z�~>���IU�΁#�C����.aQ
g��a�ǥ�kW�F�hM}���9I���3�q��+����q��	f��:�5���S5��o��7��>\��o�1qS<�]���h�m�[G#zFq�q9W]��;�<UoD�
�sG����`-�2�@9�
�=/�נ6�Yף���������ZMǻ���^�_�L�˪�7��.3Ӯ'����Ƒ�4�h�Qz{=�j�o�b��l{�����8��:&��N;iEN�P�-d�Uo�E�����|H�{]F�9WP���*V{�|�����I�F4�����ϫ�~\ ��u�Up9���L���O)��͊�^�
���(���ML����C���V�������g<��G7w&��&���7��uC�ʏ�������炱�����&����W��ɚU>�
/��ISy=��߮;�%�zc�����ap'5����G�l�oH%f���P��.�Y���q��=����{x���%�ԧ5��5��b�^�ͽN�#���¼���R���u����u�_��:ت��=F��P��A9Q'갞o��͖�3Z��+t���j�h�Y�Ų�bѓn mRC^�iݬ�u�-@�U���6�+�X������=L+����WN���T^]�0��\,}Cz}�l�^��⇲����"��P���>�}^<�A9��Ys;�Wi��s������{���w����M8�Ü����ܘ�Y(��d�C�X1ߪ���>�0�<��^��t_�2�acVGwG��6��e^���s����::���9�vR����s�*�������/}]T���Pƹ8c�9�[*Ty��t��dw�;��GZ����ag:�(z-I%��	��_� F�`�5<	�kz*�O9�����i�\gL��,�>����G[����ב�{+M3�Ix81��܁���N%�&χT�!2Z�����{��܇S��v��v�����8u�����d�o#�=�%ѝ"E����������xw=�eg��0���{U�O�����_q���h8y�����T�pȀ�A���n������J�eE9my���;��=�}�΂��QQ�����Fi��T���鿙 s��F�-�
����j'v����S��2��4&�`v�i�Ƴox+�.(�-v�<s�5�4Fc�򭁈��1dh(��T������<Qh�)}�wr���'|j
�C��]b�8�¤���B6|umܬ�|SNpk��]�8�Vh���ԧv�Ǻ4�����[����X�]��<M��.m`7����5��b�T���$�҅rG�]	��s{�Q�������{�Gf���m_I��D�}��`8��{�/��mL��&}���e�q;�8sv�RSy�;>�B��=����n��URc~m��7�t��&.3z���\�)�ӎ��}aX�ʾT_��bw�*Z���s�j�Xʅ�~z!.��~}C�{� r���7��Y�5K<r�7����ع��r�J����s;�������L`��/�ǡ*�ҍ�R~�H+*�[��F��]�í�'46�vg�{ѽ@�����ʇq��n��p�a||��;���Q�~�/�P3��D������ܪ�V�;w�z}G��o�/ƏNq^�Ý�`�|/�\䮷�6T{�I��\	��q��\���uՌ��˄��4���N��||�X���T�f�\I�KՊ-?������(�P<�Z��S�_�7{���H��Ǥ��x+&"�k
�����$�tA���g��L�n"�C*�49xc�c=\)>��z:�ޭ�W����|�=�V�!�������|,�M��
�ن?���Wъ�t-�c�Gk��s4mث޲ܦ[;f�8&�)Ý�*k��\��C��K�d�]��<�wbY�n�=E
�Yѭ�v�!��h �t�~W�r�)�u��
��j��5���3JF�����;5�B+��R44�����U1$�s盛�~~�?�Dv��8�_��.O��O-��n���"�ZO�z�~���f�Itf6�U⌶d�����r���O�����/�޳�s��w��i��*#/��xl�Kd ���t	�
��٭�s��T��o�N\,{�3��㶽Q]����&��/������F\uճV��O�����7�v�GU�;���S�w7�p7�<+� �4�kC�:�lǣ�6���<K�>﫮�ȸuU,��b**ꎇ��N�*��$H:�и�;�<_,�!�Cj�1�yY��Nq/�:��.D��q�e����ǹf��E�.�螚�7��2CPv�z^�Q����W,u-VC	����Z���[�}^�ЋcS�V����>�q�+�Q�_C~��h�<�ژ/g�;E�ʼ�xk彗�R�>@.��{nt-��K������6��=�L\���]��K�0{L���O��(<=�����T޹wК��x{:�q�k�����o��kꑛ������ �Q��F�l��-�ի��Mocsb��tՊ�Sn�yo����l)A�"=�K9p��Ы�>����� ��d6Wt���e�Fp����'Sثp_>��;}i&z��V�C���U��v�I��
Җ}e��J��*�q�Wq�\�O��t��w���s�ΌNE�EKd�=Ƣ���g�a>��z;j�V��^����k�� �}�� u�[���c�)�7�������'0�^��0�S�	�^��Ϧ����p���'�{}��`M�E�F*m���'0W�<��Ma�r,�B�hq+�z��s�{�QE+���"��h>i�t�h�=ݵ�����Y�)Y�~ ���}]T��Q��P�@-zo�c:c/�Q�#��<�lms��wz���Hp��?��۠��J;%�
�r#!��{Zd��v`�f�{et�'�g@[O��<{�3�)�[�]����@���`r�q���w��1��S�v���S�U&}��_�\=w�y����w�\=�t׸��l�K7	��2\N�O:J��zs�����S<�|��\Kv�7�m��U�u���W]���HV܈潜N,��t� f��@�q��SP�Yף��'����m�܎�ZMG��ʀ�<����0�
�[���������o�jQ�DU@�0WVѐ���L5P�|C	��.�{s�b�z1��7�@�����8cͣ�R���Km���T�s�*�!�C+��p �����gi<f�p���{3����(�ң�w�v9GX�g�ZU	�0T�T�˺��r�U�bx��������sao\}BE:���@��W	���wU���%�t���-�$i�����zr�2�����L�u��5+o�-P=��twu�7�H������ ���9���Wrڣ���ngy�#��Y�
��{�NQa��gz�\F�w%a�&�}���:���F.��>�7<��Rd���z+*�oٝ�SK�97����\*�^�m���.��{�]F�X���]��G�l��&��\4��f��
��\	|�W2�;��8.�p���:����a)�X����;f���b9^�gW�z',��E���e׏��Ne��a��9�׫��8�2�b��l{�T�?|��oS��[;:}u�쾰w��_����+^ӻj� #+���سz|6� #{o�J5nEj����ad��wRdy�p�S��ѫ�{h\g:�*����vv�B��E�Y�Q*=ٞ��7�����}K
��K�q����q~�W��c��((�$�S,&=F�zw��6�w)���3옺�	ͽ���7�Cι��_�\G[���^F���L�����~8����[*Ac�.�i��������r�u+�j>�x)U��`��"��Ц�f�چ�O�Q�.�혘���}��v
�Zz��q&��G/fv]i)�7$���%e���U���T�����<��+��Z:�q�v�̛��n��?�x_�=H]T����A�������c=�8������ϫ+���O��1Hy㳴�3�L>��S��Itg@��H�Pz[2J����O�<�gvǭ2#��<�}�Q�wo۱���_
7ϩ��;���Od@N�3`�@T��W��ҳ���:.�*h_��u��Ç��wO���ӣ	Q��#.+�؛}U=6���#Hn`\����.E]����Sw��=���gC�ﳘ�W�[g��>��p��q�����7���X�U%��$��{U�jK��;j�%�+�����@)��f��q��7�<���Nq=�f�>�q"�_�����#0-�<{��EX�n�ȹ��=/�����#%᯷z�w	��0��2TwO@��5�d?H'�&n��ݛz�\�d�r�t��p'|b�Z����a��c*��0�UP_y��u�j�aI��f3���\k�p��� Wwz+�=P*5�̕p.a���x��l��?E��[�,��z|��"�ں����{ۻ�]G�M��W�eX���顷�=C�ޠNP>�̘{��e3�':�k�~=u�Y����{^+Z^��I�ǈe�H�Q̜�}�@��?sc��՛��k}h�1�q���B�`��)X��GH;4�Yӊ�:��VE��lv+��z��5�A�G&\��6sf��.tP�Ik�e��m\D����n�g(�1i춊������VǢ%Uv�N�oG*���~�+(�>��2�k�Ӂ��31�B@u>c�`9�ѫ-�CO�����.�*�ߢ\����3�;��/B��^s�S���NCئ=��_y�^�[�7�}f�I�8%�+P�p�\`9�L�������`� �i���dѾ��*�f��OY�;���gKS<�Ӑʱ�C��c�c=\)D>��ܩ�Mk�2G^�6^��Û����}eU�F��b�R7U<���A����w��Ft��s~��
O�^��;o���i�C�R6�Y�Q%���0yT;�-�%��)�WQ�D�e?o��}��ն����w��i��ʈ���Ϥ��r NjN�!��4^��`5���;�ΏQ�q�C�e��"����ӏ�aW��#.#����}T'����\�`qi;�����KT��@�:xT�Vmh~u�ُGNm�9�p�}�'���݁6u�=qʻ�%9ӧ������r�Nw�z�!f��\GO+<Gq,?p{n��^�4�Z�U����OXx��mµ�e�q�f>Cs(l�|�r��p���k�iw�?��ˊ������G��\"�2k9[�Wf"6_<�O���ԥ��⤸̅J�U5�b{C"���S���Wk�4&���+�\ɧVZq����մ:[���zk��B�#���1R�����5���W�U���j�GUм�[6*�?si3~�E{[	U�*��\:X��x
}��}&�'��;u/k0��/�U�T<!���& �q���P/�~��Ѹ����_���sC܅�]^3*�����q]Y�%Σu�V,����=��ݲn�Ǿ��\?}������{*X�ߟ]��=3{�G`�x(� �Lӹ�F����%y�kiv�����K�p���쩮���+x�;j�V���c�Nq�?���~�����R*�{�f�������C'���Q�R�'0�2���cʩ?@���}5�'t8p�.�f�~��9������w�ˮ(x�{>�1ިȱ>3�")��)���dJ�ށ|Zƨd~�Q�cВӾ~y9.lf��B�]#�>%+3Ƣ�C��n���d�ཞ\f��r�v��[�'/���k#�Ls�8b�_���n���$�RZ5UC�yS��9��� ߹G�������T���]���<{=�u��>�����Z�g$����S:��{U���WQ^�9�8���4��u�P�Ǉ�Zi_�P�:4���r�����;���Wh��Ã$�{�vʹ�Q�pQR�ǤI��=�+&����lVR�:�$+9�!���uokqq�Wv��y�C38�̰�GE]��fI��x3&X��6�u�@X���������<�)]��\�u�VA����3�<�[�5O��2:M��Ʌa�t���J��Ih0�+��H��e����]GT�ړ��i^]L���w�nb����E��iM`'Oy
-l�O{+�1�P�;�����z@MN��E��k|5nء5�f���u�"w{J����e]�ah��K˳3�j��t�+it�|�=��6�/����dcEc�*�;��:��Qm���0G�X�7� ��R��7fȄ:����r��(p�sL��,oF�_T,���@N������G'
�pu��)���4V�L��a��ǫ
blY}��!H;v��&�K�ki	q�;��/+QY��Β_tCs}z�y�&�S)JG�Sl���6n�kAM�[�+i��d�͊·�/fH�	��Bq)�.����W�����W�j�J�u��m��M���hF�|-<�+|siǄU�х�;gE�[��<R��ȿ�͚���F��Q|��MgT9b��%�;��͛	��mV��C�zÏU���ӫrMA�iw�"3�A`M�����2�[�c�����N�j��a���h�Bu6f�1H=�V.=�:Qt��jI.e�WR3>�\�SS����r鳩VA3^q���Q���4t��>ln=��θb��Y���fn�D����ԯNr�U*q����B��\�(X�u�xY��	�޼�R��/e�Y�R��U8�f��D&�k������h�^o
>����`j��^��L�d��m�tM�)�a�fV�s&1W�m�]�۪�B�ث9\0S�˽v���]�B��G[�1K6/Mq�k~*W
C&���7� ������F�d�q�@��(Q��b�R߮rW�v����G$Ҥʶ2e���������,�ñ0�lܓwi�)A\�#���Ʀ��@-�d���5�.�#��Ȩ��MJn��E�ۦ�ua��6Z��mv_�I��qk��̝�@`��f�fY�Fk]f[v��aP��s����Ag'Z�Z�7g*CY�>����ή8����5�i��Z�c�-���)X��L��Ӽ�F��}�e�p%*�;��ѡ��7����Oe,�R�f��=�}
p��-�t����=���m�MU�.u0i�ڀ'%][�]apa v	���Rޜ,sk�z2��2ev��2��v��š��(Uqv�t{0e.Uu\�qq+Mk��-��Vv�����7�*@�*U��y��4�s��Z�ٗ�pϻC;����Ox��+�mr�g��;���޿߿��W����u�ݔF�c�wk��c��]�sn��7]�ÑN�4����ۛ���-ź;��\ӻ�qr�˕J4r��wvNwqK�ƌ�ۘ�wn���uэ]4n\�9b�+��1�p���nj�v黺帑�\��\ӧQ���.TL��wX�c�N륹��H�D].�E ��܉�\�I��X����j��3cf�u�ED���ٜ���]����e	��;�$r�77+��s�.�˴M�,�:��cs�s�D��wqɅ@d�䛗ݹ.�q��$|E� �W�}B�y�Q�5ו��ԲE����+��Գi�呎<�n���� �C!�a<N�Z��	�puw
�#����m>�M�RC�E~��}�zW~�f���>�Rx�>��v��+��������M�g�\:l.�E��<Iγ_���C�U\�ch}1u2�O��`��n���o:�9�#
�θ���H�5�x{�i��޸��x��ީ�p���|d�[ TA�\��1��X8tOs�=>��g�P뵃񜾙m�#+���z9���t��Mé�f�� h��������a�Y�!�}X���Y�r�6�{�w�=\K���ɿ�u`5��.��n�Z >�����Qzr����3�����g�x&�tn��B�����?�W 7�׀��|˯t�"O)؃�al�NԹٓ�u�5YԢ�u
�G(��V����T�⸚=��7��^�K�é��F�=P�i7?W��wZ����:���6ܱ]�������]w�<�����K�:��{��&]}5�6V�2|͙��} ���+I�>Np���:�/.��U����3���'�Be����
���&�'|�e׏�zA9���P'0ú�v��s���0�{��&���^�%��ͭz�P��ʓ�c[Rk.�@�2�$��7J{Wd-���K�,O�u�ybsݣ6�����h��J�	�b�~�*饷yR;rG_ZY���.���x��a�̝�]���x�r�F��Õ!l]��Mw�_sj�rEn�k���	O��n.��/;+�t�~�SC�NF����e��9�s�g�yT;��U���V�]P��.F�ۛ>q��[�GN�\G�W�=ޝ��{h^s��ʎ :����ɵ���<�~=�v�
Nh����K��0�P��ǫ#�q�_R���y�.3�m)J(y��Q3#���N�	���詞SNB�{5�����y�<z�����w�ͣ�=���[�Kk�J'5�8�S�M#�y$@�y.*U!2y9؇���_�u1�Ρ�m��4��3/϶�����·���{Lw��O�Q%��&H�_�̒����-���u�=.��B���^{!O{ק���U��H7�}qѷ3Ł[�1�$�@+��J5](RqjIF�W��^[��]���qC�CI�wQq]v����`�w�F���@U~�/,>���7^��R���yE.�;\&1���*����tϴ���X��� ��3p�K�-M��SO}2W�;;9������9��� �+4L=�����Ȟ,���f��$�L�&?8^�S�����T�����CV�)+z�J�>�t�N�;7�g���i}	�ںGh��-U,��)��*[��I����k/��jc�֧&5j��g\XaQ��Pb�-h�7x��n���%3n�V#��`��_&9�bS��T���G�Rz:d��mX�s�hO�Y�K�Q��C��ܘ�m��7�=z.�g�Ǔ��o,���<���NE�;���W��r���TKYx=N{\d������%�t'r������N����\*�=�9`���V���@����*�0���a�uf����ﶘ�nq�D�]�cT�Z7�z��V{�8�d�����CW{�B�z�9@�r#2a�W��������顊q^�ݕ�h�̦o+k��*��>����ܪ�V���٪��C]���yY�a��Q�����zy,�i�{��Ua��(��>\�;�gx���3���Kк��:}�:;p�T�Y�f܃�,��Ga��tL�z�΅'�����h�p*�\`{�]o�ο\n�\��Iq��M�Y�M�;l�>ݺ���R�3�� Ζ$�FYꁓC��;�+���KV��ڭх��U��+�V�~>�ۮ��5�b��ˮ>���J�3�A�L_�S)�������0��o�N��윉K<��˾��s��;h������\ܠ��T�p�$�c`\U�(�dtb�';e�t�3�ˇi�hq���8.�<<*���y�^�R%G��5��\TF�M���S��]@3�>5��ژW�v��m)^��z:������-��l)s�[}D���Q!�C�0��OD5�cHwT�/4����E�-�2��esݼuħ�9^"�8A��^���YqV��a�s��w��i�r�3���(>���9��:��a(~���kRܟy8�t�Q�/O�{��%�H����Ӑ�F��#��l;�Ě;/�%��zK���h�pEtځ�J��_,���뭳��6���<N�냜�[��эׇ;�k4�F{�fe��jH�p$�SSB��;�=�<͢{\�yY���vd�̗�Ӈ]�F��W�}�zBV�*�\�ID���v�W�����E����X��j�~�-=��Y�}�=c�������Ŀ�{��x
���\�}&ђy;u�猇��1Q/�7�\�s٘��7g<�\����}@t���4��9��B��3�H�a�Hf�0�zM��u)pQk��}E"�����\w�W]������q�t�o�]]"�kz@:z�{�lЋ�F�}�{��=�΍�ST���5���=��Eoٞ����ׅ��ߴ���w�s?�����^)�}>�AP���}'E)�r�%�?W�}zR~��8Ͻ����Y��̤1�����Sj��O�޹8i9��p4	i��`e�:�ʨ��B�r>{�VVMۙǺ�G�u���`��v��39Q�;�w*�`����q^l\.�Ǧ\=����>���:`jr%c^v�:55�aڬY�,4⭝0Qj�ךWPS��7����1x�.���'0w�aW���S�9^Sc�d>��<���~����|�#)_@s)9]�WW���>�B�9��>�>%+�0�Aه=2��9��s�Λǵ=�ё��BR�@�!඀���t�w��}T�R�h_Ϟ��IF��ѣ*���ȼ���w��ը��E���Bڦ���>��O�}�p�O�:�p�D�Z�6rK���IZ��Yqs�}��g�0����K�3��Q�Nt�DT�\}���5o]�G)<^�gH��W}�^���J�su�S��7Wd�*C�N�p@�Ft⁸����e>�n|+];Cy���hG���>�\�a���R^�%���uޘ~�ީf����� \A�\��K:�p=Θ��{&�����8͢���c�T{k�{��i>}Pp�WTKu5,�" 5_	D�WVѐ����[�q���mw.ށ���ϭ�t�"{ç&�}Հt�\VK��FIh�4���k8R��I����N�����j�퓕�uGq�Bc���=wu {�� oz�O����f1L�R���
%�[���0�SnVt��2���U<d���oX���Q����8�����,��t\�=�h��֯�S\���=���*��W��p�~�ۓE1�1�^�N���B�����{�1ګa�i��k�ݴjͣ`M�m2���f���f���ر)S[�:"wՂ���(��[���&��/����P��z��x�wفz�y�w��".����߫�9�s�����+�S��W����o��%�za�D��.�g�;&i@�[�ES�������cz;��͞D����p2�;��ÂY�}�(u}yw�Ǣ��E4�����v
�=���V�\/'���4��N�}�u�﷤�r�9�׫��9�r��`	�Y��B����"�Q��=<�GC�w���]<��͕����;�t3�p�˃0�k�ʡ�W�����O�ސ��[�y/-��ʏu�>�T��Y+�q�U�9N}ݔ�甇�O��'G��/��v����@��:�[�sqE�辯Ua���#@[]P��ǫ#�q�_R����b�9��BTu�%o�Sȝ��wx����2�I-LdWHNm�����x�<�_��w�%R��w� ��$\�����};���H+`΁?@<�*�������Aս�p���:����9E*�齛�{ۓ�,�B�z��r���Q%ѝAH�G��q2��C��
o�<�{�!1�����mGt7����{���zt+��]<��nfܦ쥱[5L��WM�m��=������nD �*XVT�-��/T!{�0wm���g-��p�3��n"lH(����.�G����%�5aK���pP4��I�kIoui�Xq���������ⷤx�u p�u��xo�x� '�c`L�
;+��v8�B�Ez9ڋ��oFt;=�n*���s��w!�!�߻�����؛��S�q�9�A#K��<��קz?ok�w��;�s�z��i՚*}M�3�=�>=��������ê�,
/'+{�H�=��®>��$H�\*K���_Y�������D������5]�A๽?�b��������l���!�١�;Ƅ�^5�d�5��C�M]ɋm��7��!C	V�{ҒS�^;��>�j=	H��?WQ^�s��![�{�w����<���J�\���N���^���]C��C�{� sy�+�!�Q��2U�.a�����0�x{,���M�~>��ܑ�oC��;:�lz��/zG}�c�e��=C��	���#q2��x�u<��2

���o(��g��N���j����J�xO����*�ݻ��*��'g�~z�>
�	.�g�4�����9�����ܡ�^��#��v0�	��q��L�-S�eg��p������i������±&^�c�@�u�w����S�/lT}WP�7~��PF���]�w��&wC,���d�޹��-���Nn ����V�}���1� ���Y���޵2��ʉKfj6]ÝMu* �=6��X��6N6䰕����j�_&o:��OV�F^��}�WWd�����ȗ�l%�������M��8
<��V��eCG�Ots�}�-y���΋����F7�HвR�2Ǩ����#t�2� d��� W�d��Ta��Z�{|�9FFٮ�\�����9�#��\h 1�TT��S)�����QS�;]ՆjJ�oi�@OH����zq��;_S��΄�����Q%ј���HX!ݞ�1�k2n��i�=�L������Ӿ��ry��:��>�${{��w�l�Kd ���nf/��O�����_�9���
��tg�i�_z���ݤ}g�V��x��Q��g'���f��7j���y�=�t�t��遀��B��/MBͭκ�1�so�ϏN��|"��;���r���lY�~���F�O�x�>�mU��h��@����o��ﲈX����܉@x"U
�A��Lm�x��%x:�@}]QE��+�2CWv�T���!�MfKʽ�ݙ�s����m�&N,p=�"�sWrs����o1Q`>��
9��M�$�7�ۨ/g,�n��	]3��Q�(&0��21��H^JPW�{<�� ���^-ǏZ�9I��}�=[挨!��Z��&;���.�i]a�FӸ�I���w�>�����Լ*Dd1gΉaS��mgj���(̇���P���T,zV���vL��*u���k�nOn<9z���T��Z�J=�'+���K{/��ut|�@�_C��4�����C�tٙX�����W��ڼ�Ѥ�>�Va���a�:��_��uޟCޠ:���t�o�]���=3u<�a�uB��Lм���`z�c'�Og�=�����ח��*k�Ǿ��+x���[|_�������q[��ߖ���k�"�ߦC'��Q�R����+ݷj�O��=��޹��n������Ϧ�K>j�\gf]i�3��B������;O~@~��K���E�h�]\����?	�st���zW>����|�i��H�ωJ��0�Aه讪Fv����'��:�/7��F���{�Paz:�u.鮹c���C���~�<�	E�$�_Ih�K��}���+��-���Q����a�oWx��Ǽ�:��Du��� ����\K��K�^�3w��M�π��Q�S/�.*z�>~�f����Rx�>�Α�}ʡ���� Xޑ٣�R�gn���	� �8�(�y�����}ΰUçj�����?]=����S��˲1t�q�1�{�`x��gv7Uh�}��-����A��7�5��IR�)�)Ǵ�w�#��n�v�H�������^�q�O����],�:�t�b���Ռl�J57e��f�Q��VC����p5���CKy��t��h+������}������O�������k���G�G�Bw�n/w`�+'q����;�;�Դ��w\7��n��������J��7E��og�
��:����oFt?tFs�_��==H��@��ɸ}Հ_U����u]3#$�l���x5��<������U���P���T4�t��:����}׀}U��K�t��a�޼��S��F6�_���b����W/�Q��r#w�����ܛ��&���{�T=6fƈ�9p�+�cv�kz��#��xml��7<��u+��y\*�%ᯖ߮�����p�����;�1N˨��t2ң�6w�%l@��V2�;���ว8N\d���^]�1��=�(���ފtqU�$�c��ٮ4�����Ug7��r�9��W���S����R�󛹍���n�8��F4��*����.�G)�ڧ7��_��ˡ��8Ne���G�C��z����V���Ǩ�J�`�g+"�WR�<�g)�����m�>��\��2�萳��?EI��h���!^�C�w���!��{v0�*+s�B��S6�nÖ2�;)��n�X�G�;Y�2��g/��%�_Ve#�Z9���1nNL��tL���|��\W`�3�9`@>ƸB7��V��R�S�t�Fz��𣂮��}����"��-�ܝ�5��}�뗷J0���ǻ.���ɒ���2�Nь��`0��/ڹ�Nv(�t�N�V�\�%/!���Ok�ŴI�ȸSqqgom6��hV�U�2��L�tqY�返�:�E�K��:������dZ+�|�YϠ��r�6}�V��<6���cY+z�A�X-�����+)
A��Hޕi���L�Wom��t��`�.�HH1�Y�
(���:+^��<���cp��ZW7V���\3@lB��<�m��,I}�ŭR���$;��Wl��@��	��ap�vpɖ��m9�>0�T�DݻC3+:嫼��3�ۺ�c�5-��9��6�^̕S��W<�u���;R��A��BY���m��v��',��v��S"�jR�:�fK Y�N���%�@��e�[Q���Gwb�#O����bgr:a]cE�%���5�t�x�!掋�7��c�Q+�P���f�R����ro8�j渺�	r3Ԡ@��
�C��y<l4v��w�\Ei���Or-��W��\oMr��3uU��èVu��%@ܬcPA9���nk[%i��lvЮ�8�z6�K���m�u6|��G��so�'�&�A#L�Y��ܨ:X��37R�np�k6���1WG�ƴ�rJ�Xݿ���wM���0�6T�w��\4*�A�לw,$������0���&�(���<�Ŏ��5u�W��y�%(�Mn*.�����K�[�`���k�2�	0�;S3����4)c����`䰐��a�]�}��Tw:8u[�gv�GPo�bs��b���j�i�mu�%���i�kp��=���c=H�����ޘW<�T�l)|�[���-Q�b�WLǶ�F7rw��.�a�WΪ2�܊?q����N+ݸ0Vn����g�c3y0T������/��KV#�'(�.ԕhe�O,�h��ѯ�\#"
�+U$X�eX���o1��D����s%��tY��qV� Y�K�с˰`p��WʰL�t�V�T�.���,�}O�;�0r��D��c��k�+��ŹUe+#���v�7s�����1C�e>,�cn�iΫɈ�7�aG�fM�5 �+��\���fn��W\tc�xa�hK��#oF��r�dgeL��ukn� ��H�5!�cR0�d��uθ�Y9�U�����`e\��S�m���4��B�M�I\5�U!�Djq�ϝK��;� �E�]�2�;U�p�ԁ���*�Cڎ��x���;�P�S<�^9o'`�9:=]4���!Ou�������r�����1;�����L�#��.u���܍�h0�w���;��s�N�ܻ�e���uـ����J�BF#���-��.��$��8ͺ��wqwwpP�ی	S(��;����t�'w]�E��6Y��ԝuӻ�w$��B�Ӛ����D�"W+���&��q���(vs�)s����RI9a��".L��\2�swti�t��s���d�w];�\������g7wpI%w:��H�뛻�s��uݸ���ܓ��77v;#9qr�wn��H�]�:�Ҕ;�'ґ�sp�������P�\��0��4�F�9��&��|E (P���ku�@p
d敖qL�I�b'%ڔ��s���w3�.Kr��VV���	:��a�Z9�ߍ����V�`b����t��O����u�[U�C�������+�.=Y�z㸿u���s�1��'�bko�%�g�j���죣���N��{�3��T�)��r��x��ި�<�=G��_]��&�C�5nGZ��Խ�����������RA@�96�R�T�r��u�{�0;�l�Fo9`��3���»s�v�;�����!�RͲ�.�� �H��ْP]]�o������B���n��v
ծ�y��edoP¯�u p�WTr�o�x�̈	��c`Oź �L������NZ��������1���ۊ�my9�r;��&���F\W]�/�g�Y s��޲n����z��v��cHW0"ϙu�&��&����oOq��_ux��PǖG�)C�6��t܅��'C�V���B�/N����4T;��}'��'����Փ���
�]w��z��ߺ��W�"�]%C[j�D��4.+�a��xwzHz���9~������=��̫hT/W=��p511q�"�	w���|.c��'|b�����=��2X�v���l0��I�i<��`�K:�]��V���*��x��K/a�f�����
Kw;\�-Am�R�����5����ir�R� �꾽DK�z^����ɍ��=��:�'j� qk7�"O49{���R��^"�V�;uZD]�]Ioui�p�Z�`������������C���#�9^��[�[�nsK�7^M�����c^_���*����q���u���hm���{���|�"�	�ޝ[�=F���
��6���Vi�/	Á����`���u:�}ʫ�o�w�/��YG'@zf�]��&�:7[�5�3�5g��Ua���k�g:�ߥ�. z!�VqY�v\$����a^���yWN{;|S7�:I×<=BgB��pdE9����U��K�q��W����F��Y�ma�_<9�~���7x�_��c�u��>+����Ji~�>~CǠɡ˷8��/y*����+iD��mj�9} 5�S�����;Y�F6<��貉*�3�DT���F�vʡ�f����7u~g��E{n� �����D��m����.nt'}R��������Wd�&���b�|�����M�L�\}�.*�[���ry��:�zo�r�2�}wý���/Eo�^+�=�O>���&��Ǹ�=&���f�
/���Ӱ��qW-�G�g�V���*�;:�dz��**g�ì(tsK�0�`aϡը���w[צ%�=�,8����wӸ���eT���f#���V�3���vd��Q��}Iz_�-�����`��SJ%Ѭ{g�&�,�K��J�/�职uը���S+-�U��i룙]=N؋[3O=�*��k�u��:�?8W��^;@i�Ԑ!��_J��K6�?C���{�6���r*>ܫ&m�q9Y�xKYP}��ِ�fY�RCW$�W)�qNw�z�m���^0/Ժ�O���i�`��=�Y�ǧ8��Q���늹s]&�S$5bv�TD���qZɧ>��K��v,	!��:3�������n����y��!�z�W��}&�'��;uYm2�Fѹ�]KX�E���G�ʼ�Xioe��n�����o����h{������fUV�t���P�i��dO�q<�B��O��*�7Ea�>�/^_��uޟ=���v]1[�}t5!��w^����:wu^��xD���8\:PŃҝ��%5�'�=Ư/n�%Mv�'�[����z�nn���'���&�m����V?՞?���k��O��uC#h��|�����;��L��=��5���ٻ�ow�U��w�|�k�Y�p�w�U�Y�s.��	�X���Xn)��x�]8�h��i����@��k�����鱘vm!q�.��d�;* ��:�4zc�շ��?�W(�K34�R�m��̮fŊp�=7/2@�Sju]Jf����Z[^a���z�Cf��SkR��:�ڥ��q��
��R�>��g�D�	���8i��u�����u��e��L�RP�Q�@S��&[h{۴s&���9s�v�����M������?ǈlT^��+�i�ަ9�:��~�.=��(��#ހ�VǠ
�e��w�qG���d���p�((Ηe�,�tFu��>�:�p�}/փ�p����_,�lNo)
q�S�'z�$�:��P�*e�����ϡ�i��z��'���q�B�/�S=Ҋ�����󾎚���6'������&�nc>���}ΰU�v����Qw�k�M�=^�lt�}����C�U��''����;�<n�2�-���k`7_��d:���/@��t��c�GO��nGu-&�=�pt�WTN:��m�� h�+�h��vj��I���6��y�vI��	�u�<�ŧ����=H���:p2nu`�}��zg�Z5�tW�*��j˛��eg=z�F���r�a�Y�a�M_I��GO 3��׀�}w��✠O� .왗~����w��tt��7f�D��T�9F�5��p����o%�4nu��=F
���7=�MV_<�u�}C�WܫéϠ��W���늕����W�K�_-�\?j�4�X���׮��݄r�-�"7�J�q;���+4G�C�i�j�Ef�\�T%���!�{��]R���m�;k��jѺ�2\k�;��_.˷arG�+�r3q��*��w9��:S;��
��F��ëZ���AȬ���owٱ�Pҡ&&�C�'�v}��YP'9;����͝�	[�\��*{��8N^J�i��EdN�F���w���=�z1���v�q��Q8w�ٗ^>���_�c�D	�0�+��v��L �4�Oz�{�6Tz��]���y���ʩ�����SC�Nom`οUd9�s. ey:�	ԕ�Ŗ������|����]^��QL�y\ �XՑr���u\3��vR��п��e���i����<�BΒX���x�U
���F�@�o���@W�:\z��q�_��W��ʲ�Ό��5G-eM{3�'��X�$�Q3�T	�I�1�NBsp�k���O:�Q�^yN�%5Y�3���xky���m\v� ��/J�L�RA@�9$�Ъ���?M[�������'U�l?���:��8���9�1��K6�$��:��"�Kff�s�Sogz
��P�O��U�o��P�O���s+7�aW�@��˙��:��l�=7ҽ]��w<�ݜ��:����	���v�UĶ������}Hi>�=�W]�6��zz;���w��ts��$kJdg��G���k�OU�7.۶�9�oD��5?uΠ��Li
�[�v:��NOׄ4Py��hݍw=y��*�Ӷ��x�}�� }�,Y��2nM��V������hfvEP�U�<�Qna�a�.��9��� ܗ�!��X)��I�h	u.�'�s?de6��t�=^�0����O���ޞ����o��P�ц&~������k�=�l�GUT��ԞSpH#����*^��_Y���������<v� =Y�/�]��Ai�ʼJ������x
�^d�����6�Hj�Պ�;ƅ�t�5q����Q�g3=��T�P�-cH��I���'�O@��3Q请�x��稭�1��N��D��������"���jby���7�g}�w�����ǟP���x��?Ea�C�z��Y�؜���
���~��-�[*1t�﨤^�k�
�����J����P�]�C�'~��Co�ٞ��oP'���o���� w��\oH�=ʡ_��h�Q�'�|j//m��_�Nxc=��W	�}۾�hX�����W�3Y*r�z���p8N���zpuת���Q��p'��;�.iqκ����&OZ�^>�$�'3������n#�*t?�쉖=QgB���8/�r9N؁��e�;�kL�{ʽ�IB�;\�`tu;|^u��w�׌�sʤW�|J@�~�gKS<�����'i��+��K'�ov���o���)����O�[�(�ԇ|ɤ�F� e�ކ������j��P�^v�yвx�kF;g�1��U���ae��ʪ���E�Wh�!T��O���^�����%Ϯ����qu�3h��� ���v9Օ6�F�=B�B��-��c=|+����(v'5�a��WeUA��hʦ$���a3z&ޥ����=U85�z�0�{�ô���Dv��c��ש����e^���Ut�uQ8�ֽ)3�
�FH9�"�X\|���[���ry��3��ܤ�k��^� ���vI���G�N������`_å� ���/v\U�v����>}#
�����Я{�=��?y9��zf�}T%� "�d���@�u��^�^���Z���cqrhY-L�Ϩ8�JfWy���'�.��UR�©!��\����|��y���\U1~���[@z�������}�����_��������3�t���0��uz�fD�B�̛�V��E�������ڬ�.Wr.!�\O{���oz�����������<��rwb�l1��^<jT��G}����/�U�Ga�[�|sTW�}@t���4����.�95�!��~��ů^��2��Ѹ9>�0����#K�Qy~�z��
��@u���ٷ����t���
a,��ַ{���y6�Fx3˵���뾑��#��u�i�՗�=��E'C��q��Z�)Յ%:�Ʊ��o�!��*[�C�x���	,Ew�s�]oZW|�FV��{RIB.�x3�I;zS�x�����EU�h��ȕ���߬o�}C�7|��|},+���ϧ����W���~�S]�7.(�#�L/mH�>�Vm�
j:�2�g?׸o��9ư���rr�p97'�"��'.2X�.|�m�)�yz����Ω?@�κ���MqK9^ዏ��.���s,�?W�y.�5����@��h[8�gfʏ�ʘ��"�r�@����+��t�m!q�.��d��a�����u79�W_����(�}�W���t�Ռ���
�c��5�ަ9���ᾗ�B�|��(�蝂�{\u��yl�I�5g*:��7zf��0�7��}�l�=����}����3U��EM�3v�Vf?�:rO\)@��g@�ʡ�T�szS;�L���}��<[
�]�[��R]���lY���	�i���k�{��	f��3�HR��y�����}ΰS+ �E��fǳ�*�b�XgxX�z�Ϸ�aW����lÎ��. �@-���iY���W]�f2��ہ�э���z����ok�/��i7��������nMK(h�4z>�;����J˻���֗oҋ��4^ٝY��90XN޳%	�}�m���+�2A;��%�&jfI��%�~��=`7i=�]z�ْX/�2�������x:�i�\�oa�ov�2�2�M�����d-S�eCY.�S�=r���V8����R�o���a��	�U7�1p�;c�J'�����V�]qY.��no}J�p=Qz�����'�@x�qE�O��hT;�5}'�������^а�#���6k�D���_��U5#��:�t��\T�9F�;�ꇩU2�&��L��9_�0;��+���U^�!9���~7<����+�S��X_�ʺ�Ѧ���j�~�065{¹���6�M�O@����C/��{�	U���W��Oa�|O����ұ�G�#��J3�3���=�U���c�����K��qZm�e׏���c�	�w�S7���WU�g��Ujq���E9@��0{���T��7\�}��j����y�ˡ���#�TEx�Wlɗ�~랥���[_���7�d��� X�����U�9NDwe ��m��~���lx�u����I�T@`�|%U�T�ޙL�V}C]�@Tn�L˩��Ǣ�n�dZ��.r�d�E�Gv{��cu�P��B(��:�S<�%��,��@9���E/r§���$a�z��Y���;���+rH�J��G|q5h�z��ov������~�E��q�Q�^�㙀ˆH7~�ː֋�w���I�����X�A��\3�B��}�Y$n�M�$+�i�[�vV��MX��t�=����dm��;G��|W��;/���+2��$Fcf�X��H\UO'>1=m!��A%�h~�w��ԏz���K�\3��8��Qؠ���p3�(�#��_A�#��"8���Ώmcڪ��:=S(kw��C]>��s��:���uuCᾩ���!��JC�n��gw7������@W�Ӝn(�þ}Q[-� ��#��F#q��#.:�ت��<7�8�c2�᤯����� 2H�7���\z�a鯖mC�O����i�p��ڱ�f���/۾�س����]����t��CI����6GN�����@|uf��pھ�{Vt˩� ��W�W�*7��G�N"W�f�>�q���]%CZ6�w���3^�ƺ�/Mg�x>��4yc�~�-�����"���oz!��E>��B�WQ�c�|'l�D���gкO;.��������I��7��U��UPQ��:f��o�w������fJ�0�{�L�r��ڍ$��h�bDM�x�����c^_�7z{
��P�W�V:�|�hj����,�P��,����,��Z��n^�B�E����I��X�C�|�eԠ�X����v��ҩδ6tv����G; 䮷p�CM��r�-g	�&�|Zg��Oq��7Z�1z�
;׺�OsP���-�|]����
`f���G�s3vh�����(M]��.3ڳ���T���f��Ñ�w�1��XUȜމ��Ԏ2[2�(���:"���(V
P�ʳS_3,i��mE/���S�s1�v\ku�s1�W���bܳt�I\u��'�p��M�0ut�OL��k`gEI�^�N^N�-L�W��^�,�����q�Z�Vm�Ly�e�6+9N��k�Xh;Nڢ�I��[��d���Y�X&z���&���������U@�y���Nc�"ͤ����
����L�mo6�76Lf�	"�B�
�[S�8��y��ixs��1N�`ЁV�f����k��}[}0��Q��\�E ��M�h������h:�D��;�Bi	]���iL[���̀ԡ�7�J����2X��ɦL��o�$���jb�WƗ���]:(��r����w�ܺA�UIx�,gDy=V�!vPL�Q���B�{�,����[{��\�b�j�鬥gp˷y�!�^pT#��R'��2����	�pP����6:���:�p���mjΎ�v������;�	�;7�A�]���wlH;{[��+9�s`X;�j���ԭ�@m�=V#�L�o��'�%v̧C��-I��(N�\$f`�5�6dǫ�k�)��PF�pq�^dOY�	[���JM�˙I�-��i]��N�]ZPii��ֲ��� �3��4����GK��"��*.�My4E��znB��[C\Q�r(�q�9���XT��uu��w�&�9V%M*�l�� QL�z�U�V��|%MkS��RVd��|��F�B,��
�Y�f���#&���ۜ�vc�2AB`�/x�Ii��qo8}N�A��= c�*��G:�VdRv≭�=}��)�*�$kvJ��ޫ��i��MN�����gHmQ"�����0!|ԛ�_q]D7Vʡ�)�E,Gw,���Ţ��(#��܂<�#\���uE�q[A���*�訜5-9P�3n��EVy��b�\5Bt��$݌a�B��tYX�9���N��mE�EB���i�`�����7t��`�`��֘�i�)�/&�vS�ai`��{w�3C.��s��lW!F��B0��-W%�cyD��T/[��YY�5�����V��uZ��ǻJl�����x�9��'��@n)�]�v�D�Z�[����Wf=۬2���
���ʶ3;�a8J�9�tcX��=n��a����w�BGKg�FI�IOR˒!f6�*і�o������"�[+�e,�؈}9T�V[�Њ��}BP"�Mˠ�$��s��%����i"R���wr�JD�Nv2W.FE	���II K(�$B�s+���F���t��@EFb4J,6QL���쑅���.L��0����͍"�]��"�F�$��"�.념�B2QC2MQ��pB*M�H%&0��错I�!�$dL�$��#&PR�3 F��r*�,Idb	1��L�K h�Ԉ4�(�Si&Y ��ۻ�;�9vJ�,"�wt���]�F
dX���g]�r��Qfr�E	FJ�%2`#�K���wp������\�Gv���0�w*d�&M�\����ź$2�Qcwn� >B�5B� >�Ю���2��V��XV:��{��gCւ�ۂ��\���h1m�J}�6 �oF�KB��ܳ`- n�'&�d�xe]휕�����F��T;�W
���'��<W��CeUv'<7��Ϊ�;�R�+�wkf���3�efgh�}��sЦ��i�8ת��Q\H�p=�ۇ�4�b���?
��"k����:\KɏxS��~��OrZ��p���\��
�z����SxX�xw?{�/ʶ�@�[�W��s��+L�s����_�7{��6=�.��"ωݿ���gLT��#/��0,��k�F���a�C������SA�Dw R���/��O�����0���H�Nl��jo�*���ᱻw[zy%>[�:*g�n(�}=�8�갻D��v�v��c��:� �7�,�럯�������(V���Nz����73�q�?L�%}�����u �4�v�((���H�����~��l�m���NIv� ��I�&�:R7Ft�*���-��s�+Nc�{"ymFf_��q/��g:m��s\s���<m��@ۀ�@�x�a����=�^�����uΕ����i���|=�p��P}��|d\:��n!��]�C~�;�%(�?�z_�b<Y��۝C�f�C�w��L���m�`�,�2�$Ձ��ά����a].�gG�=��F`{��q��z[c(�Gn�fD�a��Y�8b���h�OU���>�M9V�HT�Ʊ��n��������h�i�&�]���u�SV�v=��q}欍���c�*<\A��&��G�T>����\�I���A�M1���z.٭΅Z����G�&�2P媈��[�"�m��ǀ�L�x
}�Q���z��s/m�u]ǡz;cs\.�+OA��T�V�����n�[��WF��M���4��9��[**�N,���X/���lW@���9p�g'����0�Qxx`vr_��uޟ=�������Et�O��
�n������e�雿�z�(��DO����u/	Áqؼ���37���㝺�*:��Ƶ��ݵ\+{�F�~��\}􃓗3�*����M�8%��v,K�k��x����(��:1��aL�@O��}5�.U�0�;0��@%b�U��:�2���8m��N��mh���oe0u FJ�ށ�U�W���t����.��E��3�!7hFU�X��ՉF�xϪ:�+j��r+�Q�X�@RN�t�w��~�:��wH��\~�w븮����^���\�'MI�j�:�=�������z����Y|���ɛ�nj�~�e��3��z�Ys�?z��<�-�kV��>��ZO3sROj[����"/)�+}�UZ�aL��ĺ�֭���\�Tr�t5qN�4#�т�1��(���f*洪bsf4�e�V)�8ͣ���d+ttG]2/66T)P}�j;n�	���Ǻ'�h=>��P$���$r�w�L�=Z������]��ۮ��x��<s�^�TO�����G�����3|y|6|%��@L��I+��#ON�ǚ�+^
莭�<���w������u�0��S��=��l�d�Vz�ӱ|��֬������p:��z"�-�C�C�u��߻����+��(_�վ�Bf����]���)��Y�h��EA9ǔ{��|C�|�'x�87������*�V"q�}����w�������0�⺺����0��Y���j�M�wR��8og�@L^���v��׷�=���ރs�I�<dgҲ�U�/�Q��r7z��j�O��2\���i�W�-�&�|���G�#z���lu)ߍ�cg°D���o��<����Q�\���*��GR�P=�t{�����]&���	��#ܤم� �P2a팬���Á�_�'��q��[�r��|k����˿�����}C��d��C��p�2����	ʀc��`���7?e��F�EiXE!.�N�yE���i�ũ�p�
�FvV�ొ���=GcrS��1������e+�u�Z��F��;��F��hu���mnt�f�]�!�qI�YX�AWD-�v�Vf �[Uk\�+3d���� 7@�
�Hss��b>�`���^��t�ˌ��?W�m�|���>N�t�2;
���}�~�ބ6+�=��lb���K�a��L:���񐸝��@.Ut��Wjs�).�,Q�{'O�f}c�㶜�fw�f侅>%���3�
⺨W�\���o��%Ը���wnz�lx`ˎ��Շu�������g9�(+!S,*:�S<�%��,��{�sh��5�-_j� �sW,�>��uLw� ��6�V�f� ��1� �,\T�C�=�ٰ��5�a�EΚ��o���Z����{�Ρ�o����ׄ;���F��J����"k��?_�^U�f���F:n}������𡮟^s�g}�8�t�|v;��;�}R=[�������^�~K����T�;����xk}�qWKk�3s����F#��#��v9�>"qE���d�O�]�^OX����zn #?0����\z�&��0��l��}��ΤY��s�/�+[q�Y��G=��3L�C��,Z�-M��çD�J�� >;���Fq|-t��y�̽m��a���v���)�WAZ&TynS� Tі@�*�&j��J�$�����p�x���(��=GR�H`�6��}�mؼ��jbW&vzR���!8B���p�W\te찥��]g&6��[�t�d t��:en���7���{�*�~��>�Ć��v�s�K>�ӜK�6>�q�/��mL���ڱQ�xп����1ށ�}�����h��=�莾j�L_;�/���ކj=�x����#�Nٍn�����<�}4���=c���5�/}�c��UPq��:f����u㜇�B�Y��[����^�:݃��)���'�6�U{�������^���ޮ��{�8�d�����C_XH�(�&��.][S鮑�}@���"3&�^�?f��y{hzUWa�'<7�G����^�X5g�T����Sv�Nwv���<g/�6=���X=)�zg���CC�yQ~����3j�?�Ʀ���j?�D�u�}����q�T�Ւp��3t/EOQ�t�r��y�PWV�_���v&p�V�6��@�֮�K���y���Gu��r�V�Nf�C� Θ��T*=���Q����q;�G�$3�&�^��p���TC�|_����fm|�T$�;~��f�����Q��3��T�#!��n���Gh�㞌����������$��\[��m��paU��6fQ��pK3c�\�H�z�ؚ/���r�)x�+\�֝�)o6��'kJ��3ӎ��mPHN q��mu�̮�HF�̇�
�dV�L�
�:�=s4�xyf�ҜO"��vV2T�i�]Z�ۂ*�r�8�ɳ�̼55�T���)�N�0���@�=�⌤n�x.>��䫸�s��w��ӓ�'Ł��d���TTf�{q�tGw�Gxl䞸r Nj$����JF�Ε�_z��u���� ���95C�Y���\{����H­�\���gO��pB.�d��
x�	��\NLwVa�#���*�Br��9��ϧp�}�.+��ȷUR� 5�@�v��<c���?Iy���E{�����v�_=<����zs����P���%�t��2CCp�8�:H�q&w���W��)�}�Stz�<���c�j�"�սr/��q=�<�����p.��X�9�[/g}�r�S��OG'�S����������z�mMQqsæ�}|�|(��>�J�������Y�������IW �znO����7^�a~5/�WUaȾ�c�cT��2�.��v��e`e�],N��F2o�-)>����F�k�t�ሼ'�0�!>�z�v���UD��?8Ό��,0�D��\+}�~���7Ƹ��O��5@��_I��W��>ʣ��k�-���#߱����wZ3EM{���U�����NU���i]^��r�)5Fc�+��+���	w�"����!��12k���G>�{V�[���5Fm��V	BeW���j ,
�2���Uu��q�ԛ���dƎT��Y��+����y�u>�g����Vx�ˡpω���?s8j���}[��>Qm��W���a�O �;@��˽�:���uxn�>�B��yt��;�#�yCΒT�<eT+�+���t���Q�X�@T$�wMu���DzC��y��.(Mʰ*7�j��α��v�?\�J$r>�30�L��
������ޠ*Ie�<�R��^��z5x{q,3�ޞ��Lo�_��r�����V���u���U)�ϼo֟��B�P�j�}U����~��(�Α�n;��f��a�,�����!@<���e�2%w�������髞�*�W�|0{���r7�aW��r��w��7	��l���}�;G7w��x��k�����:�P��[V������ZMǻ����wo������P��o{�5�o	�� \�_xL=��o�b��lz:}[ǲN�&�u`z�uS�7�.��ъ�7}��}�]�=TzoM��#L�{�Q���9���[W�n;��=T�.��(�̻F�}[�^I�\���x�,8�S�\pb<�fWlz���\歮:�1�d���*�HQ�1dm��gV5�y���=��޶���z�%i��=��cyL��N��t5t+�%��5�I�=���:��:`�j�DsWŞG��+V=����w�NE�r��3
d�7f�D��u<�Q��w8L<������U)j�fw��.��h�>�{�׀���Y��:����WU���������ⱊ������F�c]��|�]ɋ�讓o��N�s�G*> V�U�{����6����Y�Ж��'�M���s�xeE�߃J�}�GL�ɾ5�����f]x�O�]3�x��Ű5]��ލ=]�#
��SFx�>��c�}y{lzS�Нr��)�ճ��r+�\����RT�P�s��\|f7Ơ�Tu�z��ī�� �.W����(u\1�3h�Q]1S�?��?~o�eǳ�~��o����;��82�e�ѝ�W]U����r8����oǙ�����o6)p����::��w��޶�ζ��IE\��:��)���!�ez}+�c��3틎~��̨Ӈ8=���sǨ�K�֮;|]y}/Mq�� ��<D(��wu�[��X���(���w\���ގ�����=�A���㵙�a���e�IsL}=f�X��bw֎��o�|�C{k�l+N��V{�z�Z��ˠ���	U�,Y��YzZ�J6�>���� ���ͷ�5
���O��e�N����O�3f�JV^e��@Dhɝ�ΰ.�<�W#[RU����R�F���eay�QL�6�\Ved;���UIz�o=��s�&τ��z*e�އ��/�O���'��gP����8o���V053"��]'�CS}8z5Q��t�pz[7S0���u�\Kk�yϫ��}@b=3�z<݃s���E�"���.#;��E\>��7�����P(l�*��	���n�?D������d/3۠e�Pcz���=���'�F_]_s3%�$����Ru/O���y��ߡ��Q�?�m�����'�<\A��%��x�|hd���p�Hj�Պ�\���wzcҰ���~���/:p�}��j;U�5w&/��Y����7��z*P���ޮ�p�c��e��-����<�U5Όt��z����P��6��_�P���g(��r�p�vJ�z��W]����^�%��j�NxÞ��Ϩ�=��c}��c�B]W��H�N;*�V�G�n�7 ��~�薵�g�����ȶ��XzQ̨w^��t^��7���S=��zzN����V��[������bw�w�/��YG=��×������m�3߉�>��_9��z�t�v��E����:9;�9���׏^����8�T���ѿJ�	}���cQ���f]�djrM�u�͊�GaS��d��mH���k`Czފ��U#�'8�h�R땭#���\l�����p�*-��Ռ=h��N�[:�Z��;j'<�3�� Ǿu՜}�Q�����7�$�ˉ�=P:PwS�8��W1ݓލL�]�[�Q��ޞE�>ֽ�WZ��미���\n�����{t�%-����9�Y�b��ͯeע��؛3�,�w�d���� ��w�VGz��C��漌\>yt�{/"U|�~޼k�6�U��$�1��9\$�G"�����?�Gh�㞌�c���ӎ���ٷV�'��+��U�ٝ���=�J6�U���	��ꨚ�%}Ǒ<�2�)�=���]y~j�hW�l���1M��Ϥ�@	���&U���ٸ������\Q~C{"$ߗo�J���� �]��^�Dx�}��#.������<\ �ِ6Cu��҅wM9��ӛ�?-��g:н��1���8�V�����"�UK7
T	n5<Θ��gV�y⩡,��@c{�d;o��=���A��%�Tz�_\U˚�1�O�K��c]l:���7��=���=���Osh�25:"�m֒��5LP�#��������km���Zֶ��U��m�mkZ��[Z����mk[o�vֵ���U��m���kZ�����m��Vֵ���[Z����ֵ��km�U��m��Vֵ��������*�ֶ���kZ��[Z���ڶ����[Z�����e5��T�P��!�?���}������s��BIQT UPPJ�P %J��� �@IH�
�B%UT%U%JP�)T�J�˞��
$����@�DT�  B@�U�Ww�� tt�
�6e
�H�66ee�&f-j��j5hX%)��)p 'J.��Eֹ��  9   H  wqu�-`�:j*��aiUe��� �t�흫Q��!6��+Sm��Ҧ��*ͫ�P���l����@�
42hPe��h [4�Am�  ;`j@(�\��X�@m�m݁@�EPel�Et�� *B��"ɪBp4�jC@��  (�V� @�� s
 I\�8w̄�6����m��0L��33kE5��@���R����k)��0Җ���j�%X��h�%��l�*Y��� ��bҕm�hl�f�d�l�)��ћb6*�I�!F���4V�E��������m�*�*�@�� ��*H�
� )���U*���hb2��4i�0LE? �)I*4��@ �
� ���H�Q��4���d�S�&��$�0&d L!�09�&L�0�&&��!�0# �IFM�Q�2=4�d���������z�w�����8cٞz��e|�m���	3���9�I�/Β�0I!"#�	.F�>J�/ !&)�F/��O�W��l�xC��aQT�*$c!$TYCB4�D!&ʈ�T%U�!&T�>|��f8�
~�|����-�	4�I�%�K�{���`�F�Y/:�OS�im�F8,�RUm����0��e���=Vw?��m�2E�!�wPÃ$��om8.�E�u{{z�T(����J������T:�S���w(n�U��1��	�j�z���tR�ŕ[�[�X��|�Ƌ�.!��i2����$�{�,�[��m��/v��(�b��Ҍi孳E@6������3r^%�[be*����"�)s&I�I���z�v��l�ͫ���������;�O쭙 ߞ��JQ6����ٽ//��a�v�; 0^�CX�I3e5�F��R��E�(����9K(�U�وd�С�	yd0>��or�c��ӚZ�ȵg��Y��
vj�ZX�ZN�ւ�c&芫b�ˢ���OsD�%�|��$dn�e�ϛ�rQ;)(a���+�Z�]����1Y5˗�5G:�+[���م�p���5��ݓc,`G^V�}i�ݨ�NM��n�6fU��.𬐨ɐJJ�f6dչ���`���̭��u��nAf�?dI�bI�s���U��ȃ́ضA;f��;����T�KR�h��y�b޼X �1��%�z��z��v�OJ�Ywi'��f&�v��m��׍���Zd���1S,�[EV��i)ov:WFm���T�����JY!G�t.��(#>���
�Di�V�.hTÒ��l��۷��B�m�Ia׻���O@�{Y��j��TD�%hܫ�/f�l<�i�U��ǄVf�V�5�=��ox.��qЪi�T���38Qae�6��wk�����1Q���uq=Sv��0S��+�7ku(vv��F�Ij�2��X�R�[��
��ãD�&ئ^屷�R��4f�o�c�Z��F�$��������ƍ^֍Υ�4&�j�8��k����b�Y�E�e�Hl�4�E����2��C]�{�O��$��.���k�m������s��p.�z��*M��9v��1���$0X,^]���2�u�7R�V^2��I5�Ra��=C���)=�0g۷����\ǡ�c�im��
�� i�7%^����ӥ7���JD�6�t�6��h�b���FP2M�A�t�_Y�Or�0�aZ�9]k/ ��YxȎFa�҅^i���y���V 6��K]�T�{P�cR죴�'G(�͔"rb%�+t�X�т��)���cB�k#��MJ���6ʀG+p�:J�6Q��@��B�����U�v��kWk$�C��b�[F�EXKx($6����[�=7�㷬lv�}v��թv� ���cK��5j觙���KF�)�����9�mj"mǳV�$Ĭ�tCI�K�k$䘘f�ѫUbqe�@w�Ej�$�jm`��M�(��姐�/]
��k�<�#t�6���q�*	EC����6%���OT	B�
O&�f�m�R�=�t(�97Hբv��X����R��yGkt�pg��z�e[�ì�Wy��Wa��m�d�iu�7x�YE�m`#��a�pXEh'l����|�ǅ	���c��ɒ]�kr�G��X�I�@���g
H�Q[4���yYN�b����:���0ꡳU���-���*��љx@.�̓p�����)���a2��tr�ؗ���؃E��1Fv����dc6�^�+8���ggvҾ*�·R����d������
J���OQQ[j�$�s6�K�48U�(��x����X�4pSM��:{�7o4;H±H#�,�gT�d�D@*eo`�Ҫ\Up��W�>���p��L�,(��=�6���N�]�Ǒ �bj�̲��35
��VL�E�.ՌSmX��s��F���"���u�����,���Tnm������w�c�:�,�L�d����4�G2��]���R���&r�ժ�L`^�����T�d��(� )Õ�a;�U��*Ҕ�S����j�A����
̰��2DWA;*ћP��#0�����Ǆm��hYh��Ň��w�G¦�9�F�Y��iSX�e�3�����e����Qբ�^Ѥ�k ݺպ�%˞��-���f+4��^Q3K�3V(3h�iػ�)e���R+SV
�tQRfkW��*e�W���႘��f��Kƭa���Y�)j�%S�l���"#a�K�i��.hb l������Mo:AX�}��Ƒ.�:$(�<Gn�fS�U�כ�!�ٰ;,r6��5yV����-��MU�czN�ݧ�d�Uw��ug0o�X�бn��T(h۴�@��v�,X�ə��-��Y�0W�B��E^1fjݦ�ڽ&�im)l��4VM�LR�ݡV5�;���6*��fLTī�.��H*87E儒v2�
r�e�w��\���r���iw7H�65)^�(o�į5�����4C�f�$�G]'��^c�����J�
���Y:�Y�`�Yf��5���:ؽ��&�"��D�j��v�l��W�5(�&ˢ���������$V��QԙR̡��`�I4^Y-�b̼�(-��E�;�1Tݔ�T$���Ŕ�U5��l�����+w54��B:ܫCw�m�[V��4o7ㄫ���S�gMj���+��� ��v�:�^^��M�ڽ��e�+�ゴh[��ͣ�b�i�p<�9�U�F����oC�B�c5�#�HT��ū�ۺ�ӵ�Y�	}��o+SO��sf�S�5*4�8l�,��t]U�!h�5]�VSb�	�W\�q�0`�0��}�-s`��I�z-b�K+{�Y�;6��������%�5�{y��a��D��Ƨ���6�֦iʗh�v�ʻ�����&SǈfZ������Q<��9�8ns;�e0X����ԉVB�pV�$�����u�ݽ�Z�y��n�C����N��N�k)��쾫�3�J���qp�{��T���l��������_��l��Q����k@�                                                                   ��                                                                                                           	$�L��If��.u�n�b�+�;^����zr��Q�����z��h��7����X���Y�rJv�����e�-76�m�ŉ�KC�W
�/x8�T��Y8;�R;��WOdܒ�'�P�1uL��:�h̜s��������l�!F%�n�[\�Z5Wq2��~}��z�w���y���M�=3�*�<6��7��(Z�͸*�o�ڻ`mZ=twJ�T��^6��e��@�����=$HN�6z�=Ǯ�%W_�n�������rTY��Ίw`��'i��k�9kS��/� κ�Y#�(���m��{�f^s�tӍ�#�<�_%����ЙB���*���Fď�ĳT�w�e�5٧b��ņ�ݥ�7�R��`���3+6����#Q�w�gbNcf!�ؽ� 
���qE���N�z��a����x2�>^	�Yt�U�262���Kz�+9ۓK5ZϬӗY�Q����&�|�k�#��W�S�:�)a3�^�M���*^�t�z���w�����˾��N�U��&��ݱ���ۇ�4b Y�.�mC]ոI�[�A岜���)=��d4�rՕeA��(��r�H	�]{N�/j:�9;@�Ƕ`��N����kS�8�������+s΂��w]v&���r#��;	�^.ZIl�mf���LnY�������g9y2��ܹ�J�P��ə]��-(S�:����lҫ��|�c�֕�@wd,s�:�58r՘�@3���	Y���[�*W�;��(��$�\sI�r�����3MY��t��w1�U�x�i����X���uҡ����ڡfEGV7|���m7��S�*Ȳ��O��)YP��p����*&S�o$�}Y0);�1*X�ZK�QɅ���i	�����qՊ��'_N̘s� ��{z,
���2�LZZ�f���������H=�⇖�[��7��e�C������_�����ܣJ��������Cʳ��E�cF�kZi<�yL��Aƨ-�^ͥ�2̮81)����6}ԃy�w]_h^�\�a�^s�aHp�_t�1�Z�ul��ެsd둇�������+]�{�g�h�f�k]�3d�Z���շ�*��b]���Fd�in*�0Z�|�!/M���9�Vn�̢k��(��qs-�XyB�]� �n��N�O֩R��˷�=�07�*}��R�ƅ�G�o0�Nd{�cX��.讫������i`K{|���x�K-r��&�r�v���a��Ƭ	�ڳJ�l|��,�ha���Y�k�"�3~4�J���p�:���-������f�������`r�ѽ�#C���S�۲[[]��m({���*9F���iT�ITrnp��d�fQu.���)��c�k�S�2ف�ux�Z�r��&�XuՔ�97�{1�Ew}�h�v�P��E�ϗKX�f�؊�Eu4�S;i��0eњY�ԑ�����k&���&�_Pfd�P�`�"������n�T�����Om�x��٭�^�m��CR\�#��Uv軽{�{u�v]�%2�WOt2�!�%,��}
Y3�a�Z��w![��:��m��k��%�c���Չ0g0ag#��֍�y����d��2>���$l]�U���Jzn[�+�w�ޖ�"�2�S��6�p%R��۴�;OYGx�Y$t������G��}�Lk�l�/9(�_:k���Z^�L�Z䑔/*+��2m�%��&ҡA��:�g�>��e��z��K�ܑ� `T��5u��Y��WkWs��g �힡�{�(d���i�P
L�v�M���/Gde;C�Ѥ�m,Z�G	W�0yi�&��Lg-�G���J�*PH뮏�L�Y���y
"�m�����vA(�C�u�. )����` �De����΋��^-�\�����m���t���d��!�m�m�J�QTMT��˷c `���OpH��PS�YׄD+4k�z�I�lܹώR�ѭaE��[}�/�5���ۆ�.�ht=}����-���(��v��y+0d렁A"������5#���ـw=�W�'�9uN
WY��(ˤ�lj��4Tb�FU�b�n-��K�(�D/���m�9Y�L(��1�I ,���/H�S��Q�ަ1�
�/C��ݭܘ���C.� Պ�Qr"�����!�k��-�I�2t�]�5y�}�mvl��{�Q�a⮿�N�E�J����j�`��#��H�������t̰qWFI�e�Y�0,�P�;�g-dNA�T�O]h���sT��~u2T�;���Z箞^�i�*�镩��*j�@=�ީ����C�n��r�_,*���Nfo'Փ)Cs�2�78>�\F��7�	&���2����V�����>�R�ޜ�U: e��<�θ���R�q5V�JT��r_V��֕�3���[V������H�a|~�R�;43�񮲮�k�=�w¶��)K��1155%�VY���8��f��֕��u[�%�u���j��Â�k�+*�Bi\��R\q��l:F�6���"	��o4��}R���e��gtډ�OPpG��7�It�Em�I�'pn6Cb
o	Z(%�:kj4�+6�s߆�]e2��"+����Q%�_=�r.V���n:���I'ZhCoq͸Y���O�{P�Y[� y/A��j���0�l}�&W6���y�:oyM �2u��W�[��ذ��ۼU����(�V���ׯ�tx�J�HA�6A��,�w�0����J� �
�"�9�鍬�$Q&�@�ڎ�I�qL�q	V̻�)պ{�y�%Mΰ��ԍ3����;���w�����   �M4�M4�Ï����=��}��o�uM��I$_lS,o�1D���t�;�M�Z��0BI ��g�����t緾���}tw�Z�N�����nr���6�8�0�v���^t��
�8���_b�\��$M]`855��U�&TĤ�Q�/Yw��v�a�]+Ȥ$�p�"�=�C$٫V�ޠ�����r<�#no ��'8uBnՌ -M;��-�� ��Ֆf�s5
�5�[��Y��Y �Ҽ�j٬5�I�g0�%!�ѧ�*m����Or@�>؈�ڌ03
�x,,P��vP��B"W�ž�ݮ-3���Ɋa�y;U����+��v�x��{�$1˾ 2,�e�|i�𭗂��\�F̐�v���X�eL1ms������>z���-\x�c����銭�;m�e&;Y"�]bk&n���U�L�R����*�p��a��w�������%�VM�$�s�Um�l�:]�zH��^M��Rb���-i9B�K���;گM��+0&r�b"�Me��3q�љf� eiB����P������J"溋.�ٕa�s`dQ}�6�w��f�v��ѹZ׭*�۱�I��U�j�\h4VݴJ�̡cn�A�Gu�b�p�Q�[hb�-^�VkS=�;'VB���%�mY�ɮ���>�=w����
�p�]��.����Bzuʝs (<��v6f[�J��y�P���n�WR',�iSS)7���u���ʠ(���h��*�Kl�	FpY�2p���t7�ST��f��L�մ)u��Uuf/�A�ǣF��%Q+��ٻ�o�5Y���S sƪU����!� ��Y�{��o`�<��T���dWV�Q0k1�_��F^�?1�x8+��c7St�Z�x@U��ƫ�7x��5U݂��ܮ����C�� ��I���"�YםV�- 3�}M�#l9O�6�[��Րwr�pZ5g��k�9J��2a6U0����mڽ�m�2۰6uC[���j�����ma�Ct�@�o�7��&츪;ݴ ���tɅ�s��:������4m�jE-�^�n�n��>ݣ�� ��Em����4��Y�E�]&Z��;(�EV��aݭU�S˗u����8����A,��r�𮦆����C��.j�N�َ�%�;H�ڼb�Wy�Շn�R�F��[C੯�ŉ7jru�!��H��Ǥ�L��]�uU��FA�p�%���"�F��8���㱬�`V���aL�dv�:��#Cr��u�:h������%�XKW��;����{��YtXnV�O.Y��=ksiz�Bn��jy�V�%�y0�8��[k����M囫����_���*�oƹ�,�4T�%�>%E��n�
�g-H�y!�V!���Y�g��L8;�4MաGgR6R&:B�m4+�ov �ۄ_!׆�nM��岋O1$��PV��GK
u��֓/0aK��R��2��}��O��,��]d�Pw!��wq��iQB�m�a���6tn�4�b6�F���tD�օ:j����f�B�o3nSs:�\��x��Y���.6ʕ6��khV��M8!\�(%����jt[Q+8ŻK�"2���J�Zs{No8e��1R�<�ت-a#>w�W`1+0�o�/��鯫�嬌���8�oZ��p(.{�2���-�+r�,��ݭ0e�6�4Y�3	�(����6�u�f�#�����IΫ.�Ű�|��z��5��V[*��T�e���Awk�0��ש.��2�f�i�rN�mj��5��*^V�' ��/�[4N��,��ғ�..��f�9�R�cY��5�YP$`'���*��,T�׳�6�4-D�afc���շ;��ߤM��ެ�8e��e%�Վ.��u	��iwD�����'*�S�.'���\�f��.��]Y5t��aN��buݓD�H��o���͌'�t!���a��9�`�pe�l�f�hL�(V��KP��/��.:t;M�OX�'kl��7�E2Y����)f��wl���Lo]�@���9ۗ�A"�)R�F��f��CI�W��K|16�pi��60l4%w��"�W]�5m�YZ��CTi�4Z�;lF����h���AP'H�iٲ���ɼD��.�R� �˾��(�Ϗ9i� J���npy�p�ǺkWvؙ���X� 5v��0.
��8$˽C:p���nk����(
]�:ŏ��q���kv�v�ך�ڝ�����f���S"I�3��s#���m���9ɠEb�\���R��5[,���L*i���\����v�C���REfu���uѡN�BΜm�g�L �}Ղ�C��X���\'vk�yWd�#V e�h��'D��ʼc^e���0�
V�1��A�(��,��WEf:�Z��ڗN����q���1�۝�ǣ��!���kq�ez�tS�:�]@ŧX�Mt׭f^�4��a�{O��;[u�@b�o��!!BR�۷�ۮ��/v�V���{w��X�+u9=�:4(Z�wr)-�%�oh�7'Na�Wu��G� Z.��2�׉��uY�+��(�2��[���U������
����x�f��"�� ���;�|qF�Cf��b��O��o��i#L�|{(Jn���uvivC�z%�g9�� �!���Ĥ�e��Dɚ�K��u&����1�Y�ܦ��oE,KB���^0�S�f����� ��LG�6)٫U���=!�u�\|�����̟��+,]YbS�2�Cxݰ�c窶��l]�;�Yw���rA�5��-'Z�h��(�U�vkz�����)��b��QEHҠ���@��|UJZ�e5�h�����P�������	,�<�*�%��7��9Ʉ�M�s�I�{]��Dz�IV0�Y���(��~5�W6Wڛ�$�J)U��$]
TW\��B0�`bYyֿ?9��9�p              2�ԃ7�yי��D�f	f�Y��YAc=.���-����Ʋ��yf	E�lߓ7�۸���kr�+�-I�B�p݅��E	��n�E-�[� -�&�i������N,i-byG4�-�i)�S]�����gy��XX�>ыF�Y���e.B�Ps���;��9�M�k���%��XE;S�OV֊[�e)�{���[��3��)L����p=�&^�9ǐ��؄�r�Yv�<������#��1��ٶY&�z��U%vWf^
�MM��L��Ĺjk��閻�b躉�'r���9�7����j�R�[K++p��B�&5%Lq�m2�i��bQR��Q�*E�CYҳ+1��Ze\�h��q�ch6��`�E�Ҵ�bZX��E�U�1i���m�S.8ȉ-�lY��P�*Ar�ci�0HE�UC�ҡDQUAb���jE�\�cR��D���Q���2�J��-�@���-�E�.YRE����d��U��ȱ�� �ed�d*%k`���������c�v���ܫo.�f���nF.�(s�Id���lMc�������[Q�yե}�I~��s�����u�鰅��J���i��j͆� �<��gϟ���kV�7l�'��Z)�cC��S{���-v�����������J�G�5������iȶ���y����p:�ee&j�(ϟe�.��I�k�4�/=��1:s��{w��mo*�I��Tl=��뾲���1�C��N��mN_�z�TA���5l,�S5VhC3�o_�l<�uK-o:�}yY�%�Fa�8�@�g8�AK�T�$�5�sq�ےTFּ�[�/^�]퍼�㴱v�RΨ�D��OE{Uɻ�v"t�����Q�bg<�gޯe:
XYη�٪���ܼow�NPRs�L����^��X�1��/�^��Tͻ����j��^T6'u�G��*^����W_����)mb��mw�v�o\!Tz��>����D��y�q>u⩚�M�Z>�^��u��Y��PݠLo��h}�fK�3A]�!�g_cSZ"Q�������:�\xC��9��ٲ�^�zSU�*�:T�rv���b�I�8�6�ڻ��ʼg(>[�SH��6S��p�F���gE�����t��d�[}N�z��'�f�Z.t�
p?%���N�<���(�*���f��=�.
<��
���؏�χ:��7弍bx��ã��J>����QM�]���ד�M@FV�6.zwϲ�g˥����\������r"D�L�k^���u���z��Äiv��X$�t���@�÷n�ϥ�噭ө�y�O�|GN:%V�Q]�@;;j,H�%�N��sDz�2��ZT�`(���s�yQ���sd��;�́������P2MN�b�Z��+G��Cޅ�Z�L�d�+g�K�l�զr	�y岮������ў��'���z;u��R��yf�u:�-��� ,�[�i5���]综�P᏶�yxC�gWjr�]N��wW���zjܴu�K�������P��lq6�WlySU���Wbg��Ȧ���49��+������gr����t����1�2�tF���.pԺ��,��r�gR���1��lWpm-����}�p�����:]j���gq�˙y���#رfʨ���1Q���5���FT���ۼ�Q:w���}�b2i�`��^NKf�'
��P��#�5.�����*ρ��qAτ�n�Hʎb�}�{`�~�]�O.{��}q"[����IsNao�K�ZZ�u&���w�w%U����U2��Y��{揬�R��js3-�!��L�Lq�7��Ėxd]ǎc��XIҤ�&-7��I;br�m�����~�	�ޞ��ʕ�f�c����j����*�v��z�wׂݚb�����f��X�/�gd��NXЮ[�L�|Mk���6�;�z�]����/m����խ�0�	�d]�e��������X��$�^�96=߆�;3��5�'�&;xŞv�%ײ�S&���=�U��@����V[�K�|&��\aZ痞�����-^��;�7N�j�Z����G�Sn��Qo�};�{V�~;N7�J�' �o)Mu.�*�*������Gi�t3f 58�[�5�r�\�	]�<�
��y��ɲ�_���u��wf�m�Յ�L��s(J~�:�{Z֫�nټ��΀z����T�}ΛhT���������@�>t�����ܰ;���Nf�P���R�-�'5�U*�f��y�����R��M��SS��q�S֯i�p�n��� �1X�����O:�u��EoO��Nx�tQ�sr�hnZ�3��p�l�:Q�s5�دY3ƥ��|����d*:��n��I'B���ŋd��J�|��t���X���C5��^U���5��N ��u�P�lm�1�_�y�>�O�^�R�v�ƶ���K�Ǒ��3G�ɵ��^�Ś��f�^#�W���-�aWw�۶�nG�l����&&���*/� ��޾�cͻ�:��Q�������fCu�O\�ݳ_�`�
��v��E��W2��lU���^�:�{&:�=��q`��ANT�v�a��F�"���ڞՆ�A��Xe�)�"/�|fօ��c<���G`sUD��(�]��_K������s��}��&�y4�LI�To�+0N���l\i��/��P���|��������>���<E@��v7�V�e��I�u�>ՙ��	��̭�=��/�5l8�s���O��5��Xg@؛�{�'₂:sܫز�z6W����V:���GUT��4��������v����P�c�7ٴ���\��)&��p��������}��i�>��3F�ءH�W��^m�nR\�w���e�j������l��s�RT���t�Z_7�uyj�C��hy@�h�/���cs���,z��Ӱ�{�^�#ۉ(A�ަ�=�V�s�:z�-\���uŴű�L��\o�S�����U4�}K����U��Lj�Ǆ�{�Dy[d�~[�ԯ�3����6G��S�3�ni��r����	�z�Qzc�\+[P�u=�{��`�4�V�y�ݳZ�lkY(�Y�������Le����>���O���o�=n��7ݔ��A�!Bmg��Kp䶶������ˈԵ�7�^wL�c%�}���:��A����E�.���%e�v���u�X�ٴ%���HM��܇7fe����G:{B-�s���dTo5�#EСz���к�>��p������FVe,�e���A�gQQ��>˺�tvŀ)*@�[Td\$�t�sz��������2��9AB�v�M	�2Tkm�	��/Gr��)�=�+C�/�`:���>.�&�'1Q��JT�d�>�P|4�U������q���&
&! ��[������(e��J�KQ�q�����4�ſ��              ⚱K1��:���]u5����a];L���5K{��r�Δj�1��kB�ٲ^�� �ƅZ��p	�{D#W�6�͹�[S���k�K(����E>nR}�@B3Ul�P���\QIW�����u3R[��dS;f_V���s��V����ӡz�F��ot�s�wv6m»�*1�ŨA��=v#6mR�h��A�S�;/���(i��8�8�e�If͋�Wm���i��#1uC�Z�����:2�%,iw���T�W��	�ْ�l(�ǢB�s�Әg3��l�+Iț���������+�DZQEi{ˍ��-�QU��hŕ*�R�XT���P�11)a�T(�,E��DTV���d(�e-f""#�-�*��J����:f0R/L��H)bX�IXEP(�ʂ��Y���6���Jъ�,̲�Ҳ�ʀ����c
���Х[*B��X��-q���F*Ł���
�mQ�-)�U�m`�(�il�-��X��eDb�Y1�$1��*�J�R�:'����ߨ�fo���(�f�����]Y o�Z������|��V�3��x�-5�::��X{5���j�RU��~
��'�<�nw��t���5��e~j���ц��-�ç$�^b�/��a��Bڭ勔W�}ؘ�R�mm6��]M�2V�����ܯA�G��j{��j�����[�Sb�~����S�S,g���3^)��R�ߑ-�~?�������ߕb���'o���IMK{�����W�d��ć�s�"2!��Z��7*ž�/}�W���	�'*���VAg�Q��`}�k��V������2vɫs�T�j⥋�<+Vю����{��ö��?���G���ܿz�C&��4�����gn�r4��P[����p�n��WD�o~z_��綿E��䴐(A�yw�?V
�i�Z����]�O���{_횴��S�i���'e�$%������[�ۄ��Y�k������s��}��rktE.�ͬZ_~V����}U[M��t���:Q�O�Xjɮ������j��vk�S��єn�'E3C��)-�w���_��6�4�\dE�G��;�W\�)빬���������Z��������^�It��:Q�����%��\^���D�ĪjӚx/s�(O��wC���٫T���F��M�����OԖ������I꡸
�D�׾mf֭#�[[[1��&�%�;�9�,����#i^��k�Ou��3KF/gq�a޷ؽ}4`�/=d�W�{�x��}T����xs���Հ�LRb��i ��HvÉĒv��|d�C��Hu�`,��q�����z��ՇSm��v��
�N�R�2~
ه���Ղ~��%Sܷĉ-R����(&*�r�U��>�FnC�C���m>B�|I���`M� �Hm��4�VI��~\3�{��y
�4�t��$P���L�=I�I�$�&$�o��!��6�i�I&�����_nI��)!�;d��P��hN��y�;a��'��	�bM�d�^Y�痻�z�^I�Hz���;g�C���$YRbN�`x�g�|�0Փ��IP$޺�~w�p>d�C��I���	�Hi��v
@�>H��!��!�OP� u�n���z�^@�$��Hx��RB���I��a'HI�\��Ψx��0��=a�ֶ}��k_k�4�:J�9��3��M{`0yd�L�d�xɦ0��:d{�ۮu���̇ۼd��Ւ�������)'>J�<�d�����s_o������淯dCL8�99`t�Bu� m���$����>`q����O"��,�d�k�~����<�0āRC��!6�L�BbI�|�̐�4�P�{gI8�m ��<}17�|�fy/�$���S+l
VNc�('�ɭQ?�V֥��gr2�#\uԀ-q���u�syq�k�<�$:B�<I�$�$4�� g�M��!�I�>B�5O�C�Z�7w����޹1'L�4��,���� ē�f�&�SHT>d4��(OY��M���y����}�C��T�<M2x�m�z�$�08ɴ�N�I�u����(|�:��������'
}�@��w�<d����'6�;Ւ�'Ht�T���^���\�u������i=I�C����2��!��8��CϹ��0 ��u�y����=N2əI��́�Y2q�<a���q'i'g���Ն�'���u��y���o�I�M2�Ȓv��q<d������2m��wHa��$�FXa9]t�~}��d�$=�C�'L�I�V�8��m�0���CV�q�ΩNw�Y�u�>ߟg�Cm�!<}:��� qr�M0M�m'lB&�,2ô����6�5��놘$�E$;OXN |j�ē9d<C��e2s �0� �$�l�l�g���}���\ﷷ����Z���]������wʿ��tQŧ���7���2��~���)\��à>l�{bZ�sη�8�~�&�ߞ��Cl>IP�$�t��I��~�d8�$׶�L��
I�4�k���3=�nE�L!Y�t�4�}П2@����;�ԇ�P�$�(g�b���{����N�8�`t��!uI偌�!��� ��)��!�0�ߝ�=��u�R|��H|s�Đ��04�������&�m���gT��>a�O�']��s�B�0�$��l�{d��l��&�bI=N���LM3��̆��~o��g$
�L��}�8�Y��I<`c&�=Ib�x$��I�{׿}�{�_k���T��2|���j�>C7a�;��!�] z�ĝ�@8ɟRN��1���Y�yν��lg� ��$Y�5�	��!�$4��q����l�`x����C�w���ϼ'l&��$�	�;g�I1��i��O;�!��z�<a��:`q&2}��͗7�7�rHs]�N2N2�N�N�N2�XC�i��8�x��VCl�a�Ԑ�s��yOՔ�Ã?oǝ�#qT��
w�_�sXo\[�/���c�D{R�r������x-��R�〈\�Ƀ����
�z��w�_�'{�d�m?�rHc'�$��i��m/,��e�ā����qt����5�|/�o�Ou$p�ư���}\r74m\��n�/Y��[����Dv3G}�W}�^��)ӻ(��J�k3�|E�[�����<���o+�켳��У��'qQ�M��KJv\���=t[ص[{U�1�qH[�ᕼ��y��9��]ٸ�]ٱ��\�:���sU݊�d�zN�J�-�~d�$dw[u��o)ު4��j�r��=\��
E�sE�ҡ���2�op�5�~���	td��Nr�%N�u�r�v\],�����__UU��Mo�����禟3�~%��o;�6��e��_
jLޗ����o��Ky��?<���;��nR��ϸ(ww)$tn��:���9g�i�85��tżM:JC<�����/L~�D�Y��oV{z�1z���鎖m�e��\���ze>�L�z����O>򊺯]�P.#�1y{�����g�尲��7��2�����nVZ��s��5��p��[`����D��Z��eĹ�u���p���2W�Tó��j)Wy���9t0�꾪����P )!<����9�ߎ}ٿ/����������Z��{��v |2+�*��M�R���Na�g���X��y�u�Yyќ�zd/#J�����f��:�����M>���x'�W���+�w}��9�F
j�.�y'�3�ŋh�J����>7R���.'��NA1�5Ny�a]�=6P�⣑V%��!��8V��.�%4���Sn�+��<н�6���<P*PN�_q3~˸�2n9�f�2f)��]?.�1���A4�ww�p"��s����s��;�s�k/��"����"���, ��,�H�,V"��!u�y�s�_:����s�Wl~^�G,���a��׹�t��**r�uy���:{G���D]����b궒�@~����������vˇfV�t�jOxs^���Z9�`�7t�����A�iSu�{*�}�f��������[����W��-�(�1���ѩ�E��mʁ���W�]okjJY)�{�z2]g�*=[{M�uT�lJ{*���?}����>���W4�}��:����뮭ݼ����f��Apb�
j+���b���*Z��{9�!�ԁ�?�=�Y��ݧ�5G�T���M�b�֜��]J��+c�흹(���P�; �47���Q�0s�{	�3n� �p9��`S�V�)Z�H����u ��[�Vz_>YְCW���>�*;޺�a��˛�(9��6��#��4zP�/k�����Yn��:�ٔ9�wXg
���@����,���w7�	�v�e�e�9�9�؋���U�'�wn��zD6�X}ac�����{8�nt�-'S0�뼦_�~��7&�c�               +�++o:f�"v�c����U�ڝ��d-h��+23������x=��C:)Wev�&��;&�;�F�se4I��C�gJCay%��w6�I�V���v��mVv��r�ĳ�#.\��������J����ʛ,���w�`�)\�೉�V"f˂�1K!�}�uzp��*�S��[�.�����W&v�2����(^r��Kf��7����_;�V��OL��.��^�W�M;�C�\�qVm��G�ec��ܣtl�u��"��u�7|���R<9yNCýo�y�o���9�y�=��������
�T+Y#j�P��ē
�()�U���*�B"PXE���L����V����( �X�RVG��H�"�M�@R( ��@�TA`�AAH(
���J�aP&"�, �a��	����5�����*�($U"�
�XA[�U�}_W�syO�����m<�^�ԭ!�n�^kj�^�r��-��UW�}US^�/����={��'�Wz'?f>:=���=*���|��H+�\�m�y���7�h~�ǭ��gx��J?Y6�Tjho�p�uv��:Oj�\��S1f�-zc0��<���˝U~�Vlޯ@g��{��*����+���2N��V��S�w~���ebo�sU�e�E�5mzJ�sr#ϣ��;`��`Koہ׻uG�=�q���25\���E�^k>���ygL��νFs�~O��b���'{x�˜+�_iP��s�� ��}���L=�}}to������������.�4|�ζ�l�f́G}���Y��I�e��^��^���붩�T�Uu��A�\�S��N~����MU����Yj�_k��v�}����a���E�9�J����'[D�27~�������թ�=��˧���*Nl��}�izǼ=��n݉���~Qtڴk���g��{՞��}��j�nf�2�W5������#�l���C\�A�+�*ֹ�6=���ɳ�A�z�s�.���������^���_����s)�������$��,��u�ޞ�Dz�d\R���f��J+6�zD�c��ژ��9�ʏq���p�`y�w�{*�O|�gZֳC�g�wJY}� �"�EO�6y�^YH�#�܂�:)�Y�m�pc���j���(�S.���v���V��.��l�i�N͊�v~��zr�����f�v�=��c�B�aK� ���Oi� ӆ����U�K�z��<;��.[iZu�N�L��6��]EΜӖ��U}�R�n-�E��u��G������R�8*J^:��"^����9k	r#�����L8����B��8��/mf�H(�39��On��D�Y��Ù�y�D`��g�8+�i��sc�܆��ҏQsr�M�Lt�L����k9f�n�������h!�K�zw���7�M�{���Ů�;�+,Po�:�(����W��jz²��9h�$��g|e*�V���#a(�Ժ�W�6o�E3��q���=�M�~��ﾯ�b�=?q;���j_��S�a[m&{�.�Oɯ_�u=�<"���'��g�����d�Ǽ�?S%�mE�ͅ�(R��wuݧb=[G��;w�ѼT;�?.����v��6Z�v�ː�qnC��購��ݠ�dc*���`��ͪ���z�;_��C:�9��[��ݺ���0�;���ݢt�׾��$�ʧ��W�H=�ݳ^�Ge�][�~ޡ��u�� �����;L�s(=r]���ݙu�%g<�J�)X�M)�C����W�;qO���X�W�m5�k�l��P���eAk'�eW�>Οk�:��Xo5����ƽ͟8���g�/sIn2��ٴ������M��\a�w��F�e֣�7K=��WM}�ʎ���*��NL��9�{�w��}����I�*�U�b�x3үtQ�G����LM�%�)�w�f�z&f:�SՍo!Ll9Ӊ�#�i�ͣ��n)�2�v�!���3F��:��p��ʐ��[���d��cw�ݭWԓ�E뮢38�Z����
T]�/E&�>����>�����1��n���=�t�0M��my�e-s����~�j}}i���x�VM�4�V�����_e3u6K��;�jU����Tի���an0�wF�s�ԇ�ݝ9f�&qO}�J����Q�,�a��Շj���
�:�Qtk� Vy���~%�tGm6���E�R#<̭����cjA��T���y��vw�g�����2+�S���^dj�pߵ����e� �K�:�5�7g$�v�{5Φt�;T�mn)��j��7"ղc�4~���v{����d��>���_`{`<���Um�~q����=4���n�3ގX��s3ɭ~�x�����u|wu#fy����oD^WҢ+��]��z86.[{�V'���<����=gb�.L���1��-�!���]{���cn�v-@=��tߣ{X��zM<y�#|M㹾��m��Q\�HDݞ��=:d����8HqDYmj��|N���8��ǳ���˒g)��P��(Q�Ǽ�76:-)<v�x�T�ӥW�J�������������7�*�~���j��y���`{��˞�6Z�Y<�I�'e����b�*v�J`�g�%`�6��徶����Y��H�@ϝw��|���Q�w!#֫Gi�g�oLu���u�'^�2���`����j�x���y�q�_S�4���W���w�}���t��bWN�{:WJh���n5�3W����!���ϗ�C�|�F���(Y�t���L�͗���Ů��~^/��y�!9v�(N���ĝr��y�3[|���qP�+y�|xn�|u�<�?B�����6�;��_��o�C�Py�7][%�R7�ͻ/+�4��}.��ϩ<�XDn�x��^�<��+�X|i�<��l,u���<���~�*u������b���N�-���p~Z#s��f�uQ�̥`���a��쥾�\�8W
ѣ��`,<*� W}=t��5�.�i���H��殮�_�4h���՚#^���*���^(���3�=w�k8�Oa��)��!;7�h���~�
P��&�Q���Ѐ�^�dl���W���c��
�Xa�Uˀ�6h�̚M�xZa����k*W_a�j��x�ho�<Wa[A�T���+p�9s�	�:��h>޳:����R�$�:\���4e[��>�ҷ
�:S�!���C�`r��ɀ'� F֬}Y�Y�J�����wR�'l�5q��(����z»�ZUj���=����]2��oaP��Q7qe���;�%c�YMH����V,�aE>�pT�#�;l,
��/�gs�x�����k�ӽK[�����I�s���P��~�@;�+�āUϻy��:r�r�.�ƺbz6��ʥ��
V�%5��:ĥ�Ͼ�pg��o#U�Y�㼴 `               ���3,��t����Tz�Fi�m	հ�Y;U8�5�$=��#�1��[D�P��p(�S��'e�XwW8��`�I�F=΃�t=�c]F�ۖ��
r2�4x6}���s:sV�%a�=n�պ9�j1gN*��u��{>�m;�pǙ�Uzڼ׽��U�6uwM;�pK���m�C�A�ë��kT�fAt�O��Sr��t�/]���;�Sv丨u+ll�zE�`�z&���`��Z�:�)臕�栧_wo��%��ٳ�PF�Ќεy�D��T�h�Zp��s~����`���EXDE�
E ����Ub�`��E
�PD� X(,�+Y"Ȥ�TY�Dr�R))���T!P
�# �%dQID���,�,��dYd+ �aX��@X\�߿~v�o��z�Z�2<�j��fn�*ș=\�K������:_x��+���r�ϳ�(.�.���r��I?AR� ���L,8#�H:��ך��!Q���޻�lة�ôҿ���%�/U���dUX�:)z�u����>'����^-�)�ī>�	~y.]pc�GS��{fG��v���(r5��h��0��Z=~f�w�Sǁ<���>���Ñ�Z�X��H���*��[�.Bd��c��a���f�K�^o��z��n�+��8Wx�x=5��ǚ^�˹R���q8i
�YC����PV�yK��i����t���l*�,e�;740�،ĝfŌ]���[Yf%�M먢���Ml�_@���W�U��܃��>�"�&j@�t8�һ
���{�Ү,`��τ}�;��8}�+4���zGWJWS��1{�Lc5�5~���$Ii�e�XB��'°Wx�Hyz��=o|�~�\�����
�e�h�"���H��^�Y����(M<��ث�E���l^�,�.w��{ݟx1v�|~����^�w^�t(Rd���ˣ��qҺhՎf�&T�xT������9흏ʸU���V��k!�i�Ѫ�lWw�Od�H�IR�^+c4ӡx|,}�-)5uފ_�2��g��L����d��u-��'{f�i���	�gk�1ö�.�5X��"��%�����}Cn9=+�ӂ��	VP�+��Ӓ�hW
3*��O]���,P��*\/Ƽ xPZ�Œ��\W��>�RŻ��J�Y�+F]^�*�3f�=��8Um����P�h0�|+�Si�d�J?g�X��PV
�Dx!G e�Q�n����Ռ<+б+��
p��.���-i�먮��<u�co������ݖ����k拾ԸA*����
�XΊ���(T �z�:Ȇ��Y'�H�� B�������Ơ>>^�nE���٦@�C������U�~��u+޾�}���k3�<�̾���� �քD�����c�n��Tg�x:�d����6��1I�_UWѭ~\=c�3c_�
=.��5��Bi:���Gΐ��;�8�k�<|Lv��{�4��Χ��z>�D{Ơ"�Dx(X��O����@}S;��Mމxh�Ua��h�����;-=o���4+B�WgƸؠ>���%գ�}�E��~͢������o�{)_O���z�S�zw��z�F�u����+ƸV�zi�����;%�>�٭o�(�B�_�3�Ƽ)�٥�uC�ev\��t!HxU��Dp��pZ�U��,�lQ�Y�z)
CG�:Ί���&��N�귚y�Ofg�B�NR9�hS'V��/w�-�k$@,�.�.��]�,������v�.��zŽ��ʕ��?}D�}߾��kT�,�t��oUN���YQq�{>���y�Ƈ
�x/ ��5>��҅1����nb{��Z(/V�J��
^$p�CQ�W����N5р�]XC���}�} 1�\��bR�'�w�^������d�����;�\~�xԳGO�^+oC�tiB�׹�����_�C^(|+��T�႕ߛ�������F_���1��>��9��g����Qv���iA
w��
0�?V��k׭h��j̄f�0��x|]+�^f����4l�A���w�%�����^�XԢ#�m4{�s��d�B�\���4�� ��>YH��:��:���~�B7���gO�wO�u�2�84�X���5���!O�}�I�_)�*Z�u3@�@��ɕM�MdyOt�bA����lw�wV<+��ƈ�.��P7����b��#�],�}�·!W\~�8M+wHgKkƮʿZ���Pу¼��p��.�:��t �y�!����(kڮ�|�Cc���yX>8��)�']����̸M�Pk5����D1���+�w[�}�C����T/2�xW"I^5���*�o��)�ǉ��{Ǉ���[˃E{�[J�{s@�mO^�^�2�xPg´SF���˥`{6Ｏh%~¶Җ�m�	y�l|�诞��ekG�f��r̈́�q�ܕ��iN�vA�C
�S����y�|߽w�����ϺɆ���zV�^)�����ê��^�y$8�h̺���e�ý1����;��������V/w�ot�+G�;c��N����e��h�^�vәt��	������G�ɗ��k��C��y+Л���}�F�Mp���5:�o�~�L�/�~F�׬[��;�to�iJ�9z�K��J�:0U{�h�U:�hc(}�w��)&�wy� ���� ��,U�5����^,S��ε�� x}Y(�����p���
pޫ�շ��'�w���
z4�[ޝ�����dK.B|��3'��v��V3,W]�z�ȟ. �/��?�}�}�V����Q_�����]�j��Ђ�wFw
����ݞ��]�yOOj�j�{C��='��g;����iEyy�G�Ǡnj8��G�W
�f��>^]rA���f�@r�(�����8!٦��T9-���ٱ����+�k�`B�P�)�=�۪>nY�v�fgyO^ӧj���o.���@���SÅ`������7W��3�v�~~��6"(Z8*�,7Ɓ4���//�,��{ܷ�aa�2���3;><lPB���
���~�r�l�u��F��a��v�a�h�+�ӻ�p��ync�T��b
v����1Fq�W`���3Yb�4�7���˙��vUE��Ɠ��6Xո-� �ﾪاyl�^�4!�
1\*��4��1�kh1���8��>��Ej��X�ఱ|k-�T:	�G:��+A'E!X)"h��M�D��ª����K�<�yK���g����
�N��~�x?��y����6��?z�3�D
�Z2����S���f�`���U���X���Q�,(Sb㣅*�A�{ �
�TX�4�!'�5dNM���І����J]l�5�ʡP �Y~�-R�8�=B���|)���}������̻�3"�|����R��^�Ǵ���y��\���~ڶx}W@/a�
�T��/�[/M ��r�Z�)若�K�wW���T��h�C�Jn�?��}T2M���_�?]p�t1F��.�]��~��<_��Q�݌�Ug�s�X������G�^�+��JG�����*��ܠ*�FwM6^uQ����,�P\(r5��v�E_��!ᵳ��|���Yn������P�f|k�+>��{t��˯Z����U�&+���D#��;��`�h׉��tV���Y�.��S�e��KMc�v���<�`�+8��p�^4���&�ׯ�A�
��A�i����B�y��R8�g�G:��ʼX�#����T:� �嚙#��w�S��J]Ցob.��*:8Θd'empx%5���+4r��,���2Pe@�u�Y����\����iL�6`���Ǒ� |l��Q�ee����sc�@��o��@E��w;�:���!��5���p@E�|�j�Sx�:�m4T���>ţ����.��,̓�C&�-�{\��,,�>�u��/�����n���|~;`�$!�s�ofj�_e�o#@3i���;�Z�՛�"��k���=�*í�C[�[Z���ߛS�0�����-�|��|n��X�4l��޴j`�q[�Ջ�,v��M�z�6    ����        g���W�1�
����������[*o�X�^S�9�v&���ɂ�nS]&�R��9�íc���sD��щ��79^���"���4[�B��|��32�c�B�u�ֵ��u{c
J���|�i�V��sZ,ܝx#�ot��[Y	w�Ԉ�udl侸V�K�D�<�}�`��P=1�Gq���$�#ӳ��Q��[v�V��{�КʚU^S�t�8���}Q�;�(����]�+���854cc��Xr��"IR�"u�ޜR]9B�i�,o8��#�+��B��P����
`
æ��+P=�"��R� c
+5��B
La
�@m%H��B��H
�a:B���P+%b�FЪ���X�*TXQU�XUeUVE��~浿x�z޺sڛ��v�h������{c5N��[�w�@#�s�zd�I���_a����>wߘg�ul�c5�jϞ���@����;���Z�'°W���t�b�>wub
wTxQ��p�S�ᵦ�=�\�{��g�h���hpU�(�]��q�%��ƋOڈ
�Ӎ;�ϸS�+���_��s��
�}�t��`��`��c�h̺���}������
��(Uo&��xp�*t�������0AP���K*U��W�ϗ��r�5�_�h�F�ƍ��Eh~5�P⿰SJ�`�׹z��¸U���4�b���Ŋ�M!�_ƿP���]�la\�6�V�-�߭)GPn�y��p�u{�9_`V�$��{��$t��5��Id��}_W��x|/��O��r��0l�_���п����Z��C��eͳu^�h!�#�5Bݠ�/�K��5�+�
�W�ı���5��������!9AȢc� X�
]F��<`�Ey�����$�]��ui�]2��CG�2ix�ZPN)帙����}� ��@�q�4Ud68}�Gm������=C�������pWW�9�;��I𮛗�����v����[��N>V����}�E�~��c�}��I�U� �jr�\}ײvD��6+@e�1�v]ACX�n�z��{C�9���Ӟ("U��b])l][yr����j�0�VX���s=�#Gk9�b
Zpͱ�N����jO-��5V ������c�E7�7R\�f�b�,D`�WAa�C��X��ޭ`��0p���k��;��AEt��!Gk;�:{E��д���`�c?1\?U莼1林�+���1�aA�h����t��]mY�M����a�CƘ�P�ń4W�i��Lؽ�I��O��h�EhEAX*#d֋��{���.?I�8��Kc��5L��2�.��*�ʝ/k�|���7�2��}&Qٓ�����NN��ޑz�����X�L�L�lB~�r��V��S�,K�4�qO�dIu!/ ��1��%�{�S)Z�F����G�l��j�y�X��u�ޮj���%�aN0?}_�S�\?#
��g�V�A��H��4���Mم�b��e��.;�/�ho���@���O]N��b�WY���^ᬭ?y��g������F@:~��B���h���~v�/g��Dm
����j��]K7T�������\��"4���5[�1�F��Xx~��\h/`X�����z4 ����z\^�a���>(Ւ2����Ο�a��gx�5����~�W����o��^���j��¡�F3��(i��Ws�7�5ܭ
�>�;��l�q�S7wUon�?-�q{\�:���>�{²�Հ�N����b�G-���o�r�l�8Grď����K~�{o���Ƙ�yM��1��I���<I����ξ�߯���A���Je�X)
��Dv�&���߲�^Yu�������c»����~0@��_��$�i&}(��Kƻ�����㉷�̈w{7ߙ�~��:]0�5�t�
Bi� y�M�&���~��4�]���]3�s}Mkym�<�ⷛ��V,1H>���S+�|F��0U���F��2���U��l�wp�*�{ݻ&Gդؔ����QY��rg�)�X|������(lU�T��5!���N������:�#7˩xU�����Mx�ô�OC0=�����љ��3����f��!Ԛ��ȺM{'��}B,O�Ϙ���J�κ��S��B1��O\Jx�}�����ǉ��{��_^�cί��3���=9���J�W
H��80Z$5�Y@��������4}�*���a�h�%���6�N��BFjr���y����������SpKٟV����Av�M��IY0׼x`����!��b
�������)P��R�=��X�
��vh�;+t�}��ꡢ�`>�^�5vp1�a���é\��j%��e��-(u��,������Mi�p�&�������W\iY�c���潲�Tgwp��S�^K�W�=
�J�q�� k���_w�6'��މ���S�wi�J��'���J	3�8o�5�ߞ�G�ګ�w�n��/�O)�>�8~���
�/ֺ )�F��i
�@g�x 9X��'u�o0�l�,<��y���~4�o�/e�����ޝ����{N<�8�:sY��֎���c�W0�[�]�V+,�B��V�<�Wy�z:�ɣ#�Y��ȥ0��f�����Ã�Vr��4�T'4�l�����½Ǝ��Y
T+�����t"��y��y�W�˧�C�/�+�\��R�.�+�&���\��xR��8/�X3���>5�q�J]J ��� � xX�4R�\2��~�Vd9anj�8y�T�{ڜ�%�6S�F6N����*o�7�����0B���f����Oy�F�~ۺ�P�F���B�6Mh�<s˽��r���)��RK���4?�F@VxQv�7�{˽�0�W�Nu�4Gњ��뤬
є8i77|.I;g�P:���
0�b+���Yƽy�,�6/A�0������Ɨ�n�{�y1���8�b
��`c��P�Z�A������4+��p���x�w�p�i��������9+��E]�ۮ�?beez�#53�x�c��~���
�rS��+�w��f�:=�Z�H����ׯ�c4�o�e
^5a=��l�N�g���(添l훎]�w��*Q59Y�e]��Ӕ�ob�3�mff,�鸆e�ܮó`-3���&C�J�UQY�����z����({��0o���f�+��'���V��n�Pn��xU��0�L�����a�}~O��Sv�4V���D*1Dc>F�3}.K������4��8B/�\]��j�ųp����Mn�� �k޻�8���잏���+�G�Ɣ.���uƈ�:��[�<�
���zj�A�JL�7�+o/���)
�2��5c�P�"
A�OJ�ח�݄>���G ���S+�((x
�v���Wk~(Y�4��x��hb���əW�¯���=�h߬|�`L�os���h�g\{�OQ�|+$������Y�ĕ���܇!�w��c��������
o�Ӷ�T8W��0���1°|I�k�gW�K�?-��A���޿
��
�|h�N��w��+�,eCc,^�=˿�Sʃ�~wS�W..D}+�{�¬���4{6��5c;�V�*^�%�}�6׽�+4ԡ��8����~>I�-Ϙ���2���ǂ�]+7��c>��XnU�����z�����P���YA������� w"b�ݟ{�.WU���/;c=(W��ԧ#ӽ��(jWm�����ܪ`�	{3�к�`/�	B�]L�B�N��5^x1տW��?���_~���NOx�b�kćmc��]�$���Rw�4���OY�G"��w9�D�F��'ù�]�Lm�9�2�`��-|�h���ʏ5Y�^�>Y]�ۍ[yE�pfeN�ܔ��P]]�7�K)�j94G\��7
����[����k�y��ά�HB�����wf���M�h�A�Vz���F�0�٤��ێ��h=߃�T6�Y�0M�n��q�G�A�t��ջO�J�wVէ�o��p3����:]X�)�Z/8l\]+q����k�S�Cv4�Kʴ��U��s��"5ټ���k�YPP�2ZSiG��U���9�ԙ2Ń�u������DI_���lm�              ����V���J���in1����mt��p�(�� J�֗a�l]��e#����;��Gȸ�f�f����ذ��/0������Gkl=J� ����32� �l�P���XN�5׺n���9��๫x[��f�n�Z/0$NY-]�:G�b�܇����֦�ή�j��7�$��n��n�]�	�&�v$��c�.d��)�S��{Ѽ�Pv���}N\�,\gL۫�F1�q总��p�^���.�{@��*��+��ʘ�����8����p���8�rE����D�%h����V���
$�a���UPTV8ؠ��,UQA}�VV���#ٍQdR�"�e��̴��\Lf$b,���,Qm�YR-VTPqr����c0����je+�Հ*�^]�W�ׅ{���>���;��.�`x!�eҗ�%.NT�ϮN�?��_U
ۊOG����0�u�C�+|kC���w�;�~e<y���tΓz)�/O���&�t����S����Df�_��˦��]�,����4yf�q����8�]�>���;M=!ߛ��o����]�xW L�]h�c]-���t��#�|/��ouV�4R�(i�-����?�l��/On}���?b���غ�Y![޺����^\75�xMVE��t+���o�+��.� ��瘌�Ș �¶�
�V��Z �&5�_��]�O{Ǟ�VJX(.*�L���,}]gEi�f�X��OZ`n�ibޝ;N&��<�1��BV��z�mǻGl�+��n:5��:�qG	��RM��d�Hh�/�~�c5hv�><lP���?w��Z� ��κ�|0W����N��L���V�{�o&��}N�Ee큨���ưy�˝���~�������׶mSe�9w���k|�����Zj#��m�_�hEA\)�h�^&��h>\��+{( �S�L���7���inɸE1Yd
�u����Y���'$@Ѣvvr��9�J�ʕ�EX�4���A^N�lL���WWXs���Кc�����������^1L6_�7��_n���<82j�?X��\ܫ����t����z+=��pVr�������9���S�3�H�����Wd��7M�W�eoa�]\�����7+�;0~�zy�h��@�h��`�E�+��
�ƻ�,�֚����_�qu+�DD�����YGo�]w\�^�>WH:��ut�CPS�վ���.(�ޞ^���O���5^��5aa�P��M�:��P���U�b��=��L��%��G!�M��X��Y޿��7��H(P�j8XƮf%�ߢ,V�^{�ZBY��:�w�͞���4���W���0Hh��#I��F�ӕ���v_��i50�4��{�Dxp�\=2\Rb�Uō]���ig޷�
�HV�5w�t]����ȳ+!I#/��6������jf�g^A�'��Ց-,�\������X�S��ֺ�Z�k1Ec�C-G�@��!���>4��� �i�0A�w��~߶���.�m��3[��x��6��4ȣ]Z?M���B�O��]�h�+�����=!����u�@3V40��NeՏ
u�ݘ��gL���V�+Ȇn]Ն)�P	S�o_N��R��զ�����K�P�`��0Wq�}�t��yU:�|4�p6~�V��q��	۪Q�v���|o�^ P�sB�����Cs��^��E�C���yut0��ؠMh�`��;�t�j�',mb0p�>6+Eh��^.غ�~)��*��|�t��WpGCH�c��F��qws �Ah5�br�]�!{�/$�S��Wۜ�G�@��3��#��o������b�t4z�ݩL�4��`��uZ)_[҅FP�>Xn�������k��n��|&����m�0F�뿜�g�y����we<�B����Y�B���^c�m;v����7KO/+�*Y-� ��xS�2i�o���*������it�z)^�];��^j��Y�Mzl�V;C��OǮ]8i�>�Æ�?G)Zծ�oɮD��ŋ҄�wL|Ƣ��ҿ��+�!��V�ϼ���c�
C��`�aЂS5<8~�S_{�&�cM���w<�;F���t{v��Roʜ���ƚ��U�V�=�#j[Ow���cZ�Z��+6��2�ս���TwINF)!�3z���zG=��kގ�'βν�m�^Ω״�w�pp���sS��Ѣ�/8Tg�2�p�5���Ơ����y���!YS/�3DU�+h�Q�O�/2�>��<<4R�k��P����U,7Ƅ�G����5�|)�@a�[H���8W���o���=���ڰ��hW@�X�++¸R�̔+�4��<���`�a�>�\.��y����:?q���8��������I�Xc���儊�
q�b��^�Ӗvy[�b��9��֓YL���4V�Tѕ�X���]A8��vP1�PشiߦA��8}$fr5ޝ}�M?%�f��w�<�z̫Y]5K%��K�7����2����]�����K/p�i�`{�j�Ӑ��w� ">��J�j]>.��Gt��"��E���o��xH~�V;ƽ��h
��b�&]���}�ſG�U8��><4�zخQTX{s+u﹧u4��Q?����~ܬo��Lк���m*S����
�4�xRg����o��z�)��]�=Kצ���@�"���u�+����F?6��t��7��w�u�.����f��u�M�}R�Dkx�vlU�ph���f���2�/��3��x�2���>���8{�ϥ���c~��5�J��ύxՄOՕ:�ǅ;�f� ��fL����t���C�8m�'���J����Y
86&�4����|/Į0�Ȼ��{$��-�ߺ�����ݙ��i����>:y����(�}6���{ض��t�j��
q�
�`����ǯW���{�
�K5�f��X�wW.����͓y�������������Mo�����v�u����+|j�L|hpb�`�^��h�Ƒ����
��x�|i��`�W�Y��u���}���������c��(�
��_)��5d��8�j���x|�wZ�|z���D���Z)�f
�D3�~b�Q���^%x���G�+(`���\�(k0AA�*B�l-��ul��� .^%]��%���s�X�K���v� �SO���8�8A��rb6��at�:��nO_��������X��)�Mfy�k�}8ҳ0�
$�w���u��h1oܧ�K�1[2��Hq?X9�,}�M�Ӥ��{��F�O��*�68p�>�,[>�l���J�Y�Y��U�W\>hۨ����O�^���]��+߶by�x���E�r��K���#M�5��:ex^��}}>B\(|�
�lc��Į�!q��z�AX>ǫ,PF��*�{-��˼��|j���!B�WP�<)\��b�(C~~�(��Y�=�ņ>��mu]X����Y0/5N�Z��36���z(U��Wv�h�և/4�[�H���t�7WJΥ��Ŧ1��NC�q]�$�Nr�a�w�y�=��4{���q�pӄ�NL�WCB��/��U�v����d��������:�b
T���z���v�u8U F�4 ��!�F*o�Ԕ
��S�O��pX�Bk�nB���W�u��wn��_����.��Y�С������½�'y ]�+���#���P�o�+)��fu�J�x7d��"�[0 ~��VxATBF�V���<e���;���4W���ﮯ�[�0|ë��������<��5�3P �py��C��E�|(��c�5h�*�S���
8�U�<}���;d�q���+r3+�U�-v<H�V����������m���C�\;��K�n]q8Hn�WG�	w87�/��HN��a��7-^�af��_oS�0��'㦥c�ע�;�t=!4�x9!J���d�E��yͣkn:g6����@cҷ��)g[����X%1��Δ��Ǐs��
��e����U&R�����ZL����/��:�pWB��h��w�v�+�!۫���tv�o��xc���&�1���x��"������^S��AI�LM����5_)����qXOq�H��ѵ�u�<�z��� �Ol\[3R�                #=\e{z�M��MvاN�ހq��X��!oK���&�p��քtp}�5B�;D��&�v�t2�ubB��
�k,��r ��1��⫳]�d�Qe'λ�mf��x��"\}Ѝ|��£���}�யM޲9<]�?�w�Y9��ep]k�)>GMl�;���u�h��.=bp<�ڧۦR�J��K��t6!���YZ}w�țKD繲c�q�3V뿔�B�>�p诔RƣN��sD�R�-ͅ�v�N�0i[���uU�������T�T�V�p��rD��I$�ٿ����
��u:K�1{�%nQ�@��[g-�T+,��8�E�(-F#hX�*��Jڶ�bʉJV�
cf	Q�)UU"��R�(�V�Tih���,U��)Z�֫"��rD���:]�l�ʔ]�լ����JK����'Y��r{+�0S����Y{`0��?
�Y�KS�u�4Fq��\=�1�� i��X;�-��m��a�²�i�٬&��/�ZQ:+��y�hi�X�=�^'���h���)�L��$�sّJZ@�Q
꽘s+'�B�9Dg��+f}s5X"��7�|;�x�����Je�oz�u����F�xoת�û�r*(��Jɇ�'��(O[��'nǹ��V9Q���� Uj=B�V��r���t���ג���C՝�g��!���i<(V:���]r�F���g�N�	�&�}���0}@`�a��M����u����@���Q����Y�Rޛ�����z�j�:�����
�\x	��9���*s���p��ж7�uDq�^�z'�͊��5oջQ��@��a��i��a|ʓ0i!��l��ɛ����P~��t�c�9���5�$���~��:ڌ��Ώǎ���O�z�T��M{��$Lޖ��a�0o�2�e���ׇaD��T��v��eN�NƳ+۪sTh�g���m�oSzN����8���Q���bf�?�W[{(p|t�r�)�:1:��摉ͭ���d�*�R(uvo^��n��J�c��{�"X��AuʍwӁ�'�x߽��:eO'�mߩ���|����;52v:\���_"��y��Nڪ{x�Ҏ̔P��_�����u�Q�	���L�Xw;OzU:��O!cs���a�z�?x�ʵ���Y�3�l~�:�(y7����u̓վ��1�r�p��Y�U^�̻k����n95a7��T��i.����|�W��T>k��Y~Iѽ$����#qf�v(��R�56�q�Ί�\Ɂr�v��N.Ģ4���=0g�6�+Z��@9�K��V`ɿ^����Ɋ�L�lJ�?��dp���MG�כ�㧏\��>�W�$����"��v|E{���v��a�.��<�M~��c��yh'ͧ�T�p����m��^��*Wl����7g�E��XK{
�R��]��� Rܚ�6| <א�����{}~���ۧMc�帨���K~��� ؔw֡ge�뒯(�ʗ�,�$���[����X��Bn]ŗ����?�����Z�������h6��f�{w����K]��]�`��󽺺ĕv�n����ϵu�:vRǼ2���I��u�����'{Z�)�8�n%��e����)/ʤ[�OH{C�4�w�'~�j��>K���y��;����w\b�Hj�yH7r�[�i�c�^���s�$b�[\�o�s�������o�\"�zŏUTϞ�[�uؔfNEʉK4�u�pL�B���JU�%L�嬊�Z�ԺW��7*;LH;��0T�s�k�Tt<�^Wb��!�ԧDC�����f
�^�t'\��x*���Ԝ�9�#�32�����ߟ���[�����[�6`n��]������S�1+�V����~�Z�J���v�E��ޜ�2}G�Q�a~}���t~�<�%j�VvFUէ6!���^�8�js�$ڤ�j����l�|��V���YC+$~��'	p}��wָLu¡ǡ�V�M��9�T���潇n勭�|^k�X6	)0��C����^_�s��,�:u~H�SX�3w۳�Zٜjo�/���匿J�xWA[�nm��|x��c*�nN��

�Y�+������m߶Zu��:,g_V���w���U~T�5����طIŠK}u�Ԡ��3�H��r�����V�ž�r�'z�'�x�ދl��Z��!yu���y�f�Tg�|�Ƿ�٬�*ϽZ�>��U��j�
5��Vjl� �7_����vW-u�2��kur%�����ܳ�2+��S���2�q�K=��n�-���S�ֵ�����x?=Vd�.K׎��OMlC�՚�M���v#6��c�ݔ�3��r��=�O!�g�į�^b#UE9n�).㝧3n�HQu��^[���q��|�-��i��n*�y��9����˛�f�S�g^^1ySެ啉������,���.w���(���C�wI�\������1=�,��p5��*�`⫛����4{鹉ήa-z����\_r8�ͭ0�ގ�u�|i���w�2/����*�T[��.3�o�ƾCy�7Zv�g�J{
/��L��ק��&�����Wz3���.��yVL�Ή�l�#B�V����q����+��l��G����;{�V���և�cc��TMgWz3���{=>����YދlT��䷙��4������tӆ��T���S�,�3fyyc�b��pK�:��ᘸ��s{�FP�PM�9h�r���"`�"\�剾�)����kiժJ����+'G	]�y��K�{(n)���}�O~:�Q���M�CPr�WK kϻ}^ge9�
��:���Fr����C����]�<'-�#�P�uKqX�/M��PUAqd����]a;\dc�-Y��d<�b���\R��'c��n�e���l��W���6�>lMa������GX'���Ǔzb���_�,����ϡ�����ߕ~�~"�?�
mګ�����7�]56i������.�i�����s��t�����3A�@O����u�fmgA���B��T��$����|-��ĕ���o#�f�B�mw�R��q7YqD}+C�̗5�5��r�ppY{Yȍa�j���=�VP�Y����ms�J�9$7eܔPashE2l˔����0#@u�졥�{��i�SbX���/���;�xցĎ�;J���μRſ�&�Z&�����B��˂E\Y�XI�HֻӬ4�=c^P�e���\��q��񉹁�зA�Wϩ�[ZH��	淯���*�!#rZ�⪵��L��Hr�V�               ���#��W�B]5�U]�o4����ha��c)�!/pt��[�
�b��¶�/N�v�F�Zghʺҷp���A�p=�z!�K�,y���y��Y�F�]�9�*�sW3�d�wZ�Lh��©*i}ҳ�M)J3{rV��RBڴ�bf^��q�����bZA­������ꥁ�;\Ѕ��@;����k��!R��Q��*s����SӬ.��L�k�9�yr����ԩ���m�n+�����;����%�՗#r��F�m�vb�k�Ӈ ��J�q)z�'rH���xU�.� ��#�%E-��1�J���J�QAeIm�Q�e`���)�Z�m%�m��,��U,-m�,���֤�%�J��*s*(�*maF��KJ""5�T��W.d��@|&�t�W^WT�[+g-�;5�����/�+${0T���Nw�˖�\� �r�;A�9��b�z����G�8�{��W��W����X��w����w����y�MLcgk\�?=��SJs�����p�1�ppCLR��R�$�h���9i�nfG�4����3K�����&�K^=�⮽}A��7]X�w�p����b�J���u���I�����T�)ԧ��\�P�Ǎ�^���$�Z�O�o�H��J�o�1��G5�A��Dk3c6��XEd�J�k�z�$"#�2�~�;��c�K���mO֪��*O���yG�e=��J������9U���8�,Ϫ�5�u3n��L����KS3ɨ��S��ψ3��tu� j�E~���U��e��3���|ZULv����q��p��Ǭ9gL�1�Z�ׯ6J�<��.}L�ݓ��z������<k�;��;�P{���4W�5����אr���6��-a�0�h8(�m���1�f�T�s����u�����{��fїk�+��Ӡ63y��"��u͏A�Ew�;L����i&��P�FE�S/e�|Y3׉\zu�p>ܖ�i��ݭ][�7Mx'�*i�k�O�t�ם���:U4�v���d�'-��'��g^^���&��3۫���R�PAط���k��P��ZFV�9]=OM=�����&������Nlb��kn������Oe�
~�k�g�M�:�m9xl{��QM,�3hmù����~�Ժz4�<W�#�ؔ�w|���N ^
M�Gh}�J�[�oWqKGs�trF�eW�m׺�V�[�2��mKӯ�[v��#����,>����"���a
�x� ����[��D��i��� S��W���eg�M#XW�{ʳ�.�1V�>�Us}oGS=�=���Zv�^����R������ܦ�{��P��E�վǽ�?B�����Y6�y�I�y�NI��
�Z��<ޘ=E.��b���{-Z�Ⳍu8M�lk
ڒom䨫4�n��t>�L?�6��!�]G�HG�_'��s���VML�����n2��y��X�n��:������L��¹�q|�����6��ݜ���p����1�D����s�z��!&�Uv�o��y�l�1tZ6���>P)(�L$��oe\s������x��v�)�CeaPr'V�>]���ӕ�7�W�&�a�}/TJ��a�=�y� �����3[����}��KG~=w��h�6GeCùw"βu}�T�Ѻr�7�����邎�{����:����+�90T��]۰���}�|�Lt�ʥ��z����aEg(�������Ƶ�&�O��U���%y�wj�K��yfx©�O�ݫ����ϗ��n'w���>�ڞ�����(ֈo����{k�DR�ǾF�ﶮ3��>�h&=ɶ�>So�qW>>� _�E���4��ѫ�"ghz������t��Ae7g�)<���m���G��ٺ}:���ݬ�ݬ����f۹|~�:Q�O�@��Rևk����J���*7B�QS
o��?��[[
)��71�C�u��麌K��;�����N�B퍥�r��I(pd�����A���]��������M��=R�MUF����:�i���٤(���ߥ�絼��to�ףzO����^e���q��q�=�IP>l�\�Ռ5#�՗�����1ν��5H��c�ײn{6Gӵ/�Sh�๪M{���U������8�%d���w�5�$�Bn�K0m-D�d�q���F�^�u��]!���W���Һ�A���kM�o;�|�.�.Z�᥌���DL��sU}�Y��e3Ly]ܶG �G�/b�ncOǏe�I�>��}�m��-=y���w!�.��yLa�M��+�����~�1�)�U�i���p��{k�&'�ّ;jB�l�[��ѯ���ř�q����ٺ�V�q���v����Ğ:x{��l�hg��~]�0��7D���r�z�.]3k��j�o���k��y[X��r�&o�w%]�l���,<���3��g�ŕ���6�]1���xK*.�*�}ݻ@��,�}|�W$�ה�sge�L�^��z�3L)�ͮ{�u���V�#}�G��Ot�56��h�ls��[Kޯ=��U
��C��.�*7�k��W7��F%m]q��Q/�gv]N8�w���}j�\VC�٫��'�v�d8mU���؆����.�Omrݘ��c���C�U���i�F⩞�B{/�:�d6q��Y���Q�O_L���c��\����JT/��ݤ�4tM���,6���;���έ���.���}x�Z�75�j!V���U�V��+E6�� ���г��u�k�{�C�!��w=��=��ݟ{UE��=����'�{7R5�F�O�Zk�[�弫&wu��T,k���Ǎ-��q��MU�%������O1xZ������L�s��Zs͗��ڣ�S\��EŔ󴆭�/G�p�w��t;�c�6n�c�ٶ�m��` b���$s[�m��Q��˱غ�*!�g`��'
ͧ�T���{���n��_�9��NP{]\���pJ���W-)Y�+�>�[��ŋ8��<�w�Ժ�����d�=�`��,Y��7�86⤯�u�gn�CӸ�<�f�1����fg9Fm��=���	��n]J��,Z�A�7v4T��
��Y{B���t�)K��Qx�[�C.���tȬ��f]-�;�Y�rd�V&̥�]VO�!���>϶죈�>�kw@��]{ӝ%[��7�V��Y��ﶴ�]X��Hm:Je��tM����E�|Ϳ�p5r���\s!C��QW��                FT��Q�r�ʬ�>�eJ�t5�]���FG��3X2�y�>5��C�P���mW8S`�/��D_E|��[��@�����u�a�V�E-�WT\��g+G �M*.�>79q��+c��r�h��k���>��e۽�5ISʈ#�i(2��`�]�0�`�V�]ֻo�y���tp�]�I�Z0�郛\0ګ���/�4^�X�a��Z�p�p;q�W'[[�w9����z�u�����֛0�.��G��:��>�C7P{pLp�XB�����{7�7ɯ��)��=�nI�7$\P	@� h�YQKm��Z�/V���EPm�5�(��҅J�-��(WĢ�J,b�)U�bem�Qb*[m+qɊ*��FT+Ls%���U[b�KP����ՕiJ��kiT[il�9B�\���.e�r䶹kZ�*/�N[kE�h�i�c[+D[�e�&��.3ThQ�({"~���W�W��E:ĭJ^ w����5do�)�2`��I,��R�ѯ){�5y7I&k�{0�&.b�
�8!C���yr�雂u8��{O�tH-�wX�
a↢a�(�v�,Mx��d����iv���C��_+`�}���|(�u�ŀɧ"�-{�*��YC�'�5�l�$'�����M�"�}�*���.k�̫s�{R�2���4w���z4;r^���X�bh��������������:c��Oc�z��yeś9Ș����7;qd����^�;�Vx�����LtކV����&�t+=�Qæo��w����09����2g�w���y#��3�iJ�ܨnZ��;��y	�$��R���j��k��-�td�u��ӽC�r���ze.����Oe�z���)��򝕩X�61v��Z7-�CN�H��^~�Oְ���m{̑��є�(�z�Q7�9�o�_T���4R{19�"�r�ǽ�$�-	�v:�ڍ�Z�Y��%Ez{�)����ˎ���_�1����ӝlewr��3�j����z}�G,'�i�o�������auz��{�"t�5>O���c������yd��}'��c�E+o��!��}%����^5�օ-5MW]^��ƕ�?w=��c��v_���W��a|_~�B%\;�6p͔�̡Z�=z�ӳ��$,�L�#R���(���底��JUq)?t�-�n=��_�ٹ�����6r捏;,w�h��W�c�|�1�&��8v�h��7i�n�CUuJ`<���M��.4Mi�3Rӆ��e�����ư���k�}���XH߹>@S������g��\�\T�_�Z�X/=#ԡwy[M�z;Md�m�*2�;�Ӗ���<]a���G�K�4P=�7�
��tc�:w�;�z_���S�(:cΆX�x�~�7���+�睝����1�f��I-e����jTs�^��/3���B�e"woӞ���#�m�5�Wy��Wx�=�C��#ĒO��3r��F��}ֳr��\;ogq�g_si9�]��]Εo.,Y&�ԡCs������/�vyS��T�GX�W�<qfԛ0m�d�ceu�@<S������9dN�i�>w.-�9+�[�t���f����E�'�z�O�4���k����Z+U~�gӟhc�^Oܸ-Sկ�;���S��-�o��s[��{4�մ�)\�y+{����޽����m[����؇�w��/�G�{oh�p����<��K���^�`=%��xS��9i��;�M^�gk��	}��]�P�ǽrm/֐�#�� �}����iz���Wnf���kRΩ+ǯ�|�k�OW�X��]-����^;7-W��Me���:�<���B�/[[g��5�g���?~��~�Nx��5�6|SU��:-V���3ؖc�K�A`�uת'�����Wr)�C�V.~f��J��N����<�C:&�}m����=EãL�ؽ�>�2n9g�����CxZ����o������m���N���HY[�T���r*i-6f��J����%-9��rWr�����b�'976v��W�_���Z��s�5[��V�h�U�^��=�Ԫ5��}���+�Z���n-+��#�?=35tr��k�Fk���=���^�K�j�9���F��̔��1�&�����ǽ�Iy�]�0�>��v�A�/fa:G5��'�oVM����Kv��E�P�bcf�J�ۇ�Q�^�"(d�v�zyS�_���/�1Y��_j��J���K���;|�6.h�Z�G%:��.�[Z��sz8O�_7��dY����.<��c<��ʮ����n�#S�&v9,�렷�,-e��&���ڊ�]g���K��>��^P���=���F�q�j�ժ��N-6�y���/��P!���*1[����3�2���ޗ�w�Z�^������*���4V{y��������l��g	�Ǵ�¨O/'��V���D�#���"��+�)�wNԨ��BZ(vS�l�
�;G]ȫ *s*$6��=Z#���N��b��V����TNgJ(�'w���x�7Eowh��+�+���[�E�ɑy�$v���-Z��.�A��K��yOw����>����wMe^;��r�W��._�<�g�p��*�/{o�1��5J~�Py4tk��ouy)QvL�K��}#⩻*���}�'�RT�d���Ϸ��^��8��Ǐ�o�dB�#�vm�"񰯕��OMm]=��0ܯ{��k��=���9�/��a�'�g@o������:uK���ڧ�`�@��ld�suǓn���۱�J(����S�(NC,�8���jw��qśK5��=���4+9C${���Hk����D4c���[�vz��^�Uz�R�A;^��<y(�h���ڇ��-'��������޻�i�~�s2�yL��5n۫t-��s{���4`n���hƪ��>r���{�����U�n_����m>�b�t��,��V�*Uŝ���k��2Φ	��/V�>�ݢ�5�,ק���4��D~��^�]�#~�����ę΢�i}u�)B��.�+�����ZZ�ܼ��ġ�������Ƨ��	;�i,�]iX^��ަf��������W�qB�{b���c�
5Ն�X��7�5���1�d�u��ֱk��6��]��[%d����/F�8(3�e�نq�����f�KK��ɒ^�T��/fX��ⶑp���DoQk:є/lokC��/�ew=%m�b���ֳ32ғ��VF��]��m��<}�4��ng�3]�t3����F���.��62�S.-���pg2RM;�:r��-W#��W0uD5"�r~��Kg���{�               �>�8^�iRq���^Bx�gz��3&l<Q�1jK/2w�8B�t��y�[�n�
�G)Q��2B9n�n԰�!W����
vJwҥ�_gn�0'�w`;XR���ݫ{òo¸��cx�%�3S���Mq9�;[�P�V#��A熬�ud����֌�ب��%�������,�=v�d��품�wʘӫ���w�3ִ<+��Vnl��pP+�m5���Q����m��8'�Z\nC���ͬ�VM9�}]�e2����1Z�.,�-��ܯ��Ev������l��J=��������㘹�8a�i���U��B�ch�mi�¦"ais�bًp���e�q��p�E��\j���ګ�Q���1��2e1�e3.fca�bf�)\H��Z"-i��q�-(,�R���h㈸�)H,*��Ʃ2�Q��T[E
�P�D��PX�f�����Aj4��B�Vm�"bT���b�4���d�LIQDa�<ε��� �n���������i�_ ��]19tlU�O}9�mJE�6�w���ζ5�=|�K7�Q�[�\��VR�V�BU2����{0���:���-��PjU7�ۧ�ۢ4+��C�&�޳&e{��`M�k0�"���J!ֹ��X���5�ڍ̌��X�}˚�����R�:�ٰ��/g37WW ����o��r1U�;z���5�����V��S;}��&{��d��m���Gn��T2�~ⷵPZs۽(Ǉ�z�W1��yޮlg[Rᳯ�4T�qA�9)br���rt�Xy��I���Ϝ���;6�����G�7F�����!�gg�jjw��es���q��CU�n#a�3�������B���y	���G��M��в�xS\�����T�l*�Mx����NM�J����p� ��^���y,?EOG�%쥠�����y��꘰fH���:��5��ߵ[��@�x�ȗW�oc��ѵ�ݩ�!)�PԵ@o ���Ak ���IiM�:�{�D;�	��{1#+]�r��6f/��b��n{��y�U�G�#:�p�{�T��9ˆƪr�N��=�ӓA�B�]3o����]���k(q�0���K���:�.{��Z��u-�q��]ì�b������HN�?*n~��F��S�|��6g�ǳ*���z��>�����7��|��h����R~�m=����}��g��K�Q���X���X�lW�J�ي~w(�������.=�s�o)�2rҲÙ�J̕�t�_.����[�k^��54����]J5AU����+�90WK�EY5�z�JPp������O��5<�N�l�s���P�%c����I:h.c��ָ���)=���玗�>�sӭ]��r�^�j���ޭ}�w_ChS�K�n1˩ΉGTu�.����rM��H�/f��K8�zve�[��^*��Z��x%������bԽ��pj��6�b�c������3�bO���{��eE�o�F#-�O�}E�wJ��!N�elhym�Ͼ¸UЭ�뼡u�E�68��V��A�WֳgȲ.QG�e�ԁ��H�q��G>��L
�f�A5��Y�<�]�X�����y˦�l�}��ڂnP��9+�.?uHD>)��(q�=��U��G�2�#�Ӡ�X�zi��U��v�X%�g��L�j�3 ��;>��W�g���Z���o�U:��*oW�X5\���}�t�ڳ �[P�az^7���=x>>b� ��O�^Y!�:����oB�汁F0O�o��m\��u�=�1^�P�i�Du��.�Sșý7	�Y�ؿiյ˯���W�6m��Eh�(UY��;ջ ��Z��8ĉ'�B�U��=^}$|8�N�X��C�':Tt_��<��'�QB{��=���S!�5mt���..)v7��S��9�$vB2���V�i�י�n���ppf���,�+��Bx�J��CY �e��v3�K��yZ�W�i�j����s�Ǽ�ǳG�.���Yf�#�����,�V�_�ݬ6$�k���gfʞ���j��R���{1J�����^�>'��;��°���/]��ѵS�r�t�9t�_̊jL���Ir)��n�Vn���}�^+jOb�I�;v�9.i���bޝ�L�}��B��`n�ʶ���u�5v�=�w�~t5��]�;����uw���]ʺ�ˮ�驕ez� O)���+[���^�|�_�k��N���s��Z�gp�zW'�	7�,F�S�T����y ��Oyr�i·�*�QQ^�.�]}�K����dꡰ��î�*����=�=�X���v���tS�l���b�ۘ�n��<��Xx�7v�e���x�{Rû���Cqi���6g`�h�bI�v�3�6��7x� ܅Ki�3΃�{�ͨ�7�H�Rf������붜���oiQۯ'���}��������d(�wg�bz��Kx�� ��7�N��-.Z�_]me�^Հ�o�QSϡM�¸���2-��1�A}��ES.�'|#��tŶ�#��o��.��'Om��+��j|WO�.�6ۓ��td��]c�׎6���צ<ѭb��g^Ů�'�y�_�yN�c�C,Ȯ�d:wc��y�yQɼ�1fIR��s����]�**cw���ӗ��'�R��&����Z���?/v�3���¤�d�����1�aZ����Z��L�-�h���d2+�޹B���K���o"��Ix�ekȝ��=�r��SuZ������7��:TZF�ylL��YY=�]�U�u��ߛ��}ά���KU�zk����Z��_K�*Ye3T�gvz3��o���gJ
?'��z�q@ߗ��u���<��Z[���t߫יni��NT;Iں�C���t���64��M�O2���\Z��ڴ�����9r/��ܥhu+d�-wM5e'��˵*���'c��59�7�f�UW�T�ۧ�	�[�S�ʲQjTՊ�u�^�Ц��v19�㯲�9���my�M�����I^\uO�ĿO%	t������:�8z�qe�����A���עc�%M�q�En�Tg�mt���48���=����ҩ��ɕӹo��4�=W�Q���A��h�����]����~�����S�T�UV,���Є�Iz���� ���&�HgI$��v�#6�
t3��/���_��t��w��D�N%BI*�"A�D��X�$TBF�3��g{0;�;td,P�?$M�[m��=����KV�HeŤ��G�8U�BH$�RUn��V������l���>C��"dԝ����C'��tP�������(oA�?<
Rjs廓>aW\ٮ13�9���$�O�~�-���ɥ��JI�u	$~�I�����:b*��]�?��捫'�'�"z��g���v?i�bv�D�go�� �Q��o�Σ�IJPٌ����H�H���S#9rY��]�1Eh�j�W��~a�z�I(ǣ���*�����"�K^��I�b���IMM��{w̸v�����HH~� p��d�p�H�aC��)�\��7�Vl��7lOكk�D�I�L���URYő�	��I����Z��__}������q��c�:'��͌^Û�{?��?I��f��i"H$ǒZJ�ׇ�F�N�|Q���wd����.]5��,fG��o?g6]]�l��8I�>�ߨz����9̼N�S�f�r��	7��IEj��u�zOSn)����]J{ņ�A٩T��a�"��\�$}�Ԟ�)�X��'*���8�0��KpI�Ȧ�1bF�!䌛�@���X ��2`��IGɩ7J��BKEI��b��H�~�ԝ���p���5��(����"C$�Գ��I�-!ɰ;���`U|�`}��$�Mr����lH��!$Vy;�~�$�p���\��>���Z�6����������9��2mad����]\���wM|�=q�D��tH���lj�>߹i	 ���pǡ¸����Y/����A%���e�V�w�}!���s��M��8	v�z<3֌��gK�=\�^)E�z�ɹCHs�Ѷ����kQ�����������g;��7e!$_��(�0��zb�n�nX�5)�̲���	�eTuTYFՙ�en:��,z�����D�$�O�$�B�Ǌ4�GUyO'	�[���A't�N���&�(��dc���$�*�E���e#tUJQDwE>$s�ډ����w$S�	��հ