BZh91AY&SY
c��߀py����߰����aM~_p    }        l t�  M+���N�^���64�rP�m��+[[�����Gvrհ=� A& .��У�1�`i0 p                  ��   ԳkZ��_g����:�딽v���Jl(5#Z��ll۾���>�G����
����J�@V���/M����M�gim��$��;��vǶ�(gw�gvVZvzL�����  �W!��3g��Tn���{{���|c�{�:��p��S�t[��l�PQ�u������x�f�}����W{��P�uyt=v�k�m��we۶涝����H��vIn�m��n�+��RE��G�   C��{��tn�������y�;0��ӤӶ�s�4O<�gvx�ר�;��Z[��n�u�^)^{.�r9��v<�ݥo1��κ��tK�. )�  ���z�h�:7-�ӝ׊x;�X�n��I���fw���[{k���
��m�w{��n;��{x޹��2ٴv��9�ؗ�^{��s��NZ�f�=뢂;   N���{���䍷A� n�ر6�c������̳�_ ��Uwy�}yw�Ϣ�K��۴�j���;�e�4����O`      B� �@       � �              �~�Fz�T�L	�� L� a)����(`#	� 4�  �R	�J�FC �1 � &F`��HUMC `  F  H���4&M���3$�d��@�jR�Q� �L` F# #�?0?D�7?U�P~��~Ԡ��T ދ�!2O��'�  T�Q �*�_�P�A+��/����?����������I�,�?���B(`�P "�����J�P�$��ѕmU~����k�e6�� �CQe� �;�}��'����g�/������^o�[��6���i$y=��� &��}�v��<$���V�e��MM�������'����y3�'�D�rL���~���'�nD�D��C�2'�p�&���N>+�K"u�ԡ4Hݞ�ǳ�����0��ȉ�5]8?&�U�JؔG�51��DOw�bX�ʳ�89	]�X&T��Rh�e|����DO2DGd�D(~DN��1�'G���;8]}F�'0s%|��x�)�J͕��jU���"y�H�r�p��ϒ����ea�7����a҈�-�G"P����ԤN7)nM�ӂ/%x��Ҿ~rR'3��%���k)<__W��D㒑=��8k�ӣ̕��ʮ���D��H�ܭ8<�}�5)��D��D^Jӣ�J�6;+�s9+�[�H��Z��/�����"q�H��V5�i�NO���ʭ,�����)�xn%vRa�eP���)ݕ�;�1$�r����ܪ/�}�ݕ�3�<_Y^;!�G��$NԳ����͉�ep�`x��� �p~r��}߫*�����>���H�Du���Zz�l�MI��N�7��lGbw�2N�N�y�V	�j�h�*�����4Z��E�a�~ì�S�dF��ȗc�4岫2��1�(jA飕T�g$��nA�=��{�vAϧ��3=�[�.G����~/�.	�w�&��x�B�	��W*UȜ�=���V;;�fy���^��W{UFvA�ӥ�*ݕ����p������F�G��N>��em�y+�/g99��g&�fGc�������󒝞:���\�+�r7)�yUy:�Wv'1��	Hv��T�7r�A2�z3^�����ջ�$=����e��LM�&Yg�d�C���$�:�LD��$߷I!;���������Kâu�=�<�=î����i�GM�%�E��¢K�K�MGR`����ӝ����|Q�����I\-+�:�I�H��&��}�1/��N"t��=��'>J��v	�yC(��R{��$�
nA/���g䚚+$߽�N�YO��&p�d��L�᧸���'��2o��&�=�ߋ2}�
2$J�:Q�r}��-!� b��,����8'8�5<P���J�!i�h�7�	4MHoɩ	�%"jX�l�?'�(�H��ȚS�)>�M�H��~ϓL;Γ0N�������8A<�tH䉂s/N��搿�t�M��i"&�D�����ƶO�2��N���K�H���G~xO��2�$8>�M&�ç['��DNa��"{�&%�!0�Ğ�ӥ�=i�R��N���҇!�i���P��N�D�O�6QA<�I4��&��y�x鍓�f��
�DJ�DՒ��
����Dt:P��,DNq"`��rH?%��S��$M<�&ĝ87	�'�O|���t���"'��7xl�!>��}��)��%��4�a���#���� ��"#��i�='D�
.&�%%��ϊ�'Q;}"jh��|G����L��jaʐ~3�Ȓ���Eژ{bxO'����NY�X�OP��ǧ�xy8xN��Oe��W�q�D���/D�Ӽ�z�KA؏ܜ�F�g��Dt�5����987>���Q,�Y��}��Mك�0�U,�YW87ҥ�gl�y!���v��
�ԫ�ȍ�a�tK'��*D�j#�V莥$�<C���;���F���ڟ�?'z���~?z�~��;0���=��T����S	���WnG�2N�a]}�4|�K/�a*���N˝�NOM�L�T�I��̨��1�)�Y㜈��'N3�=� ��D�l�Dg�_DE��=>������ȋ ��S�yUv�#"{��S>�"/*'����j$1<q�J�Dt�<S!_#9Q��"Zԡ!�jY��E�K�&�����wdNBJ<]�">$DRM:W"#�TD\��Zԡ=�H;>OyR��<�N�j"_�A��G��B"�J�M�����FUM:7ڈ�z�&>���J����r�"�D�֥	�5:A��	��T�ڈ�ͨ�|jQO�;���KeJ�Q������d�8p���G2�w�"�:{'L9mO	�jt�{,v|�{�B�r����rQ�!_2|x>G��'P��=Bo��!���b9��D�v���+Lz�rG>��<ڝ�gji���jY6 �u>�Bd9���}BO�ݚ�*���F��K-�vG��ǡ�G���]�]p����E�3�?a�l��L="50F��L#��vښg"tε0NƧ����aòQI�G�ʟ>�=Y��P��a�z�y����ˇڳ�'�����=�q���z��l�*�qu;���r�-��ڝ�T�I.�|���}u;�����u��O	�4�0�YV#��v�����OjVɞ�]$zI9F�Q˨��rg��MOSS�65*���[��fw*T�J��Q*���Կ��R����⯦\�'K�K�w+����r;�L�>��2G��̞Ƨy���Ϲ����u.�/�>�T}$�b{gOT��v�i|�M��ʏ�U��jdjp�'fT��Nq�d�;>vL��s��rN��z�>���Զ�%gj94�jeOF�j'�*w������+ە:���)��$��l����O��jz�cS�T�j_�;/�Bچ�4�!��M�%֐�T�rSۥ�F�=����_g��5ƣ�bi3�⾱�ʲ��	NJD霞�JMl����Ӄȉ�#$N�,����"uex��:<䯑ؔq�&�DN�����%�J�DG6W��R�K-�LnRh�+�
�����ea��N�9�����J ��[�H�ġ�����H�nR'��Dy4�����H�K�J�w��)0�2������ȉ�Y���y+��Ӈ�'^JD��i��Г���H�nR'��"�V�zW��JD�rWD�ґ-e'��+���H�rR&�L8h��},rg
D�ep�gݒt�H��']���U��Jwen���ۘr����ܪ/�}:'D���q����pjt�Գ�����v��/̮�$0���J�"�}߸�}_o��ܔ�4M�Q'�\Dweiݜɩ6z���>��%lG�='F�x��I�5��=�O�"h�U&�0� ���jx����v`��Uy��2D�~�e�n���i���{d���샟M�ݜ܊�vg2?d��~'d�����OC�a��z���<�n+<>�o܎����Gޜߣ��s�w���_n/��9��u�V��I8iYR�ܕO%S�V�S��J��~˩U�l��ٝ����w��jL�V�!�I��������E�/����w�w'��NG��^�e���MIs���;C�<�Ü����Q�#X��jJ���4�����n���3�i]�N��ѩ��J�֙��p�7F��ɝk���;���T+������9O�O��5��O���ُѕ,?,`b?�I�x*�I��%I�#���nff~�Sp�ox{��=><?Q�o}u�t����y2nV�9(�ROI;$��~��Y!V�;��E�g��S_*��z'�L_.,�.'�5��Yŕa��.������Ȱ������թ)����<��k=���o��?.�;�K��k��eI7;31�CZ�����_�5797ũS3s�R�92}�OO��w��rL�J�U���&�5Iyf��ɤ��������������;7=7.2�@e�\����s=}�~92dgf���2V�2[��GM���ύq�1�7�p{{5��8�8���W˫UM%�dYS�Q���������w\㧆��_^t���>�:�����맗�����\q���{z]���w��Ǳ�����\{=��<�	��7N��΃�<�=��۝�|c{����ӏ>.���ϸ2!�\MU��g%MbDA�S���6�鑟_J��6'*OaL�'�U�W�Wˊ.(���G�qu]\Mqu.9����s�#����#�}�fFl�g4�O���$�����ϳJ�����z�ˌ:K���S�ܪuv˞|q����6��ǡ��^y����c����ޘ�y�Oc�On<��ȏ �����|�����V��|^MU�U^YVgW�Sy�K�*��+~\^�[99s'�Ez|˛�62����wJ��v\�W��4ӗ6�٥T�=>>�8�;}n6�ç=�����7�g4z�d�������ꪮ�Uj���������&���Y�̪$�Z\UD��s��RQ4�Muo�ϑ��q����..(�eџ�-�:�>�/�S]Y�05=>�w&j>�'e���U§�3�TL֔Mg�=F׫�rE����7G�U�tv�Nz|��g�g��*�����ӌmǾ��x:v8���|xs�Ύo[�,x�RW�D�W��՟�8�~�//|�����dY�[��_���.��wuy���Y��f�y����-�Qdq��B㘺��Q�s���+j.㽔���Iȗ�s��=��
�q�sGQ��j��F�7\1�J��qw�����j8�����.�GQw��a�W��evzz�U4?@�!�[�ҽcG%\�����@9�@5,��
��Q�{�I��&(�	㘗9��e&vW��eGtj\,��s�+�Gc��wԬ��]F��zUw\u�7�����8���Qu����J�.�w���9�˝����/�Z)7��ʑ�蘝�Zgc���� T91��������Q�M���R5���)��q�vUF��ț�Ej�K���CQ�Y��FG1Ɗ�\YUUQN&!�R����w�}�=Ä�İ՝Y�B��eG�D�[��n<�IL�Rf<��sem�7.2V��J��(~k��y��W�u���/��y����e�p��qvVl��UǱ{��=� v5G0^��]��v:���=��D��y���x�Ƣ�j�G�I�f=��tQQ��29�9N4UGq�sr��]�p=���ެ�W��-�*Ƴ�>Y����ýeoc��(�W�0��eN�:ղ;��|+|*2QUG1�j<oM��cxoyo-xq��Íӌ��J��q1��ǓQ��s�\���Z�X�`�qcMg���"k*�"�3��sb�$y.=�M�Ǔ1ܑ��uyg�����������7��*k<�,�,�,j~�}I6�-YV5�� ��Y�,\_b���ӄK��3�R���j:��GY͵$y9H�&�/�E�qg�Gk�gG��Mg����{}oN��l[�u��>����ĸ��t)F���5�����nr71Wm�UJ��qe<���o��ޝ�O�-���F����ǆz嗚�y7ET�n\n}@�.:���SVU՞\YW|?�VT�=]�uU���T]0a%}>��oѕɭ�g!�?xwZ9=+S!��n+�r���I)�GӲ�=+�]I��9��%0$���H:��%G���,K�*�:����$_�Z&Vj]U�����qqg�uyg�Q��$��x�Y���U�oG�#�JnM���y7]��H�gVT���*���,�,i�Jh���,�̜]YWzBU�U�U�.�z�c]�ҵ]�k��:/��0I�}9eo��ݙ�b7*#��ȸ�3ME�u9����wE��ʍLƌSS1��/|o��1鼺n;n����<�/��T���A��7)��M�}'
�\y���8��єƨ�{�B�M�d�Gq��+���d5�u�R�+҉y��N�%zT��;�:�,�kʘ���GՊ,��"/8+Y�t�����V���8�h�B�M��w ���~d���U�FD�+:�.?QR5l�ǴV##��G��G�؛�6V��#Q�q�u0�v�@�u�F�Q��u�S��#�H͕�͕q��{��Gqt����G�w���T$�M�Z��Ån7���F�wZ.���\y�R��V��J�G:7
���{�%v9fY��pWaNZ�nK*�q���:������B�U�1�/��6FG1�C��7eFjG��{sE�� ����^a9�{F7M�yn7���Zt�������ĳ��!o�d7t8��F��:�c��70����V�L�uY]�_GP/k�C�ԩ+|J�x/���m>���S�%gGZز�c�}����=
��J�Fh���4oX!1��uG��s��mg8>��B�*ƱpueX�#Q�LC8�;l�ƸT������j��r�%�ck9G�tu�v:�!�u��W�+�e})�UG�$5�n�����f���~�1���@�2��Y\����<��Y*��sƣ��7Gq��eH�� ]Q��?Gq�w�G��~�I� �5��;g��nʑ��9���>�!��7�l�એ�+0�3�TwGq��dq�X�P�)��Q�u኷��dJ�@2L�s
��tV��<�Gq�M��S��q�{�#���<��Aq���8�G�)�;�0J�\�G���ŕ��27�19*J>������\GиjvH�3�����zS(��Y���ɩ�W�,��?N͙2\�ﳼ����lc;;�'�G��*���լ~���o�g��H�+�O�V9���^�G}�Ͼ8�?i��4�]rc���<Yx��w�s^���˭E9�c�O�K��|�Թ��F��H��=9���v��ᒨ��$uE��M�����]����yv��O�wy��k���˼�F����w�#��Yfs�����{\p�ɨ��ݱn˺m/6N���ٕ3d9Ʊ�"�b��e�MV��`��|��{�撍�L�t����Y׾�^�W���F���F�z����;�K��;�{=.���劕�%��sޥz���������}�/=�������<q���ͯ�t�,��^v^��#�{ǧ�\�G�prrwo�r��$��'U[�j�)�9�g�Kچr�U�Y��z'�s�є׼rÏ�w_&J8^i�3�Q�97]���s���ܞ�l}��Y�%=�kF��������{�+��/k�Y�[:�vs��v��7Zg%�*��E����y��hI9}�QΝ��/q�{��NE{w��[�n��{9�՟s~^���ۼ'�]g��쥊������5����7�3nK�v�+���k.�'�|�ߏ]�S��T��%Vʕ�����2d}���R#U~]����ys��>v�m�W�[��u.l�%��7�T��^j'����!��d�!��~0tǍ��q$]�*�
��bT@.!7G��	�{t��M@1���G�`��q�N@GpsԸ��+�W�E�D��P��j�ő@D�K������l��ů٠�3�����Mr����\CUI���	�Pj<�Y�@;���7H���73j�5��5���Qk�����QI��H��REj+3M���ˈ���8�Y��a���Q�� �� ��wf�Dh$�z�|���1bxD���Q��e�ƞ���E%�%�ܲʂ��]�5IX�#y�Fmx8��ʁT�A�;&�՘]�-,�La*3
�DUa��wOϰʄ�
�U�BY�9ǈ�1,�%��Vl�D�<k+������H���3Q�b���i`/�퇬CFU�ʤ�7���6�3�5 v�3V���@}C��Djq(�3X�&���5�T�g���a��ٴ��>CUcXr����Z���fj�������/lHL֦ .54B��9��sV��3\m8(ߩZ��{@�����2h��]�[oO�|]+zW�U|iD�n;�b��I�~ f%f��Q���&�_Ԡ�'&�f&��1�S���N�0�R���\D����n'�P>�W�7��/j��ں[��7�yv1�{뷾��O�~��#�_ꤽ_t�
�ϫЙ�F�G����!?�|��������?�����R��P�*�	 �dP�	�����|W����s�����/��^*�UmW��yU�W��U_"���UUU�������U_+�V�^��U|�UUb���^*��x����j�U[Uz��U򴪮"��-*���U|���n�qZUWU�UUťU\ZUUťU\]@��ҋZij��\�5�-[�JmUƮ+L֢֨�ME��Q�T��V��%DF@@�THADʾ���u�������J��^*�UmZ]b������U򴪮"���UW��Uz�j�U_"���UUTUQ]b��W������U�V�^�UU�UUTUUu���w�^���x���������������{��Ȍ��(H����E�m���Rljƫ3j����ۃm�	>�6|��$��V�WV*��*��*��*��үWʼU_*�Uo��W�Ҫ��UUb��-*�UmZUWUUV*��*��*��*��-8��[U��ZUW�Uq[��ťUUEUUX���UuZUW�U}��|kcW�r�k��*��lEY*����N�u5�b����~����U_,UU�iU\X������⪾W����U_+�V�^��U\������-*���W���V�^�J�⴪�,UU�UUťU�b��W����V��n�QUUU�UqU�W����U^�ګj�w����>
�O�������lkV6�qm�"�HTV��F`��bQڮ6��Uq��W֍Z-6�Q�h���V�ۑ���~����r��$�dL��������O���?i���`��K4��2�� ���Rt��B"tD�DM���O�A��$8'������&	�a�	�i�'���0M4��t�"P�'J:""'L ���pD�4Hh��'D�,K8'�$:X��bx�D�:"A4E��ibY�8C�P�A,�� �x�$,D���X�(�ƚi�&'JDJ�&�"h�tN�P�X�DA A �%�>6�?������}��6ʤ+j+mU,��$�EQ,�ġr�j���R7K�	B�<�5$��Gbj�r��%U�T�
6�UD�!�77^\�T��",��T�M�)%�ˌI�H&GJ�d�Wd�V��A���P�Z��X����Dݵ�H4��E�������1�D&KG�q&���I���,#�u�b�%cI	#J\YS�]�����Y"�*R)A6�UP�"�X�LJU]���]"�D�R��Jլ�K%�4HMtZ�Ǒh�"(܅��^8ݩT�m�Un9�i	Qآ�8!�uђ�db�	�� �LDuE��,�8�J��vڨ�chR�I1�S$nbM���uiDT;��ڛ��µI;�m!:GJ�E�$�8��40�X�%�KK%V���"w���)�U�j�j+OP�mrؔH���IU	Z'��[�1�,�.,N&��JDRI+�ѩl�VWfQ�#$ʙyP�D9��Tl ��+U�B���T+#ʋ �R���#l�dnK!`�DDx��<��\�D!1��Ċ�L�ȭ�����(W���׊�Ś�Dq��b�j,�"�Q�%��)e�#)$ġ\��L�GJ�\r�*�a뱭`�{h��qA0tNZ�"�O!�dN�F��t�
�D��"�@��	CV��c8kKRVG���ў�ZQ�ڌ����e+�52T⮸8X[J�S�$�B�2֓J��9J��LDo"���LPXژ����pec_Y�tp�Q�IR��V�E#"���]g"hx��7�FQ�!�m�FFƆ�]y�^;:�0�)FV&Yq�R���m!�e,i\�V\���Q�CvT�X��o.6�E�S(1�J2⤰#�Ą��-"1<�t��1˕Q�R����e-(ҡP�"By-�)��hi�Lb,B�A�T)��(��bǖ1�iZ�2�bj)P�Q���%���(ɑbt����c��<Q#Y$X���ʘ�Q%i�*�b��Y#$j"�,,�R̍�R(�cě����T���la11���an7D�j����H�OCTYSu���̱�%Ƌli&TZ"E%�y2�e�X�G2b�Rd�ْ��J��)�LMn֒�r��t����!f$�jZj"㱑eBB"%����+�*$F���LhP�V��'��Ea2�1��)�
�82�1�iīc���5k(��7�K���Ŭ�fH�ie�aX�$
��Kk7sn	�G�&�J�&*�ǐ��c�)q1�&BB���dƄ�rR�Q��c�Y�)	��PEedu6�X���������EECf'h܉�\l�TO��QD� ��QU��VQ�ڭ�*�ˍ�nRW���A��+9��X�Ȥ�ph��"�&,UH��)(��cQ+~Vi��[ą�,Y+l�YPR̤��FH*��r��#-(�����Z%I�hPD#�$�D:X6B�YKq<�i�Q�"!2�Y(��M��l��Zʜv�6TE�
a!hJ*�n��ARd��[,�9iFWD!Q�%$��e5�0ѲA�`���8&6A���R��QP�X��B2,�5��A����ЋE2eo.b(��(��P�X閡<te�u@cCDT���li�boYX��1R��KU�N
�q	�"�Ȋ�F*��
ˋ�b7X������+Gj1��E��+ЩK\��)2�'n'UH�=��Z���# ��G�B}�638b8݃8�q��T��"XKkU*�n�h���dL�b��FYmb��8�"u�k���TЛ�E[��A�T�I[v��ȣU�YI�H������D���\��B���#Q�h��`Ɲ�CepTJ9F�KZ%�JUc��bOU%�lnW�`����cIA2�]v���uYeiX�Uq�$qC�D���bDty)Kd�"T�N�I	e+����j�Sy-�J��ڭ�!;QH�Uv��j7�Ԓі�Ume�Q	�ڭ2X�R+Q��(Y�֥UYZTJ��d�*��v$�I�9X�"Pm%in*�N�ثRcUTU�JET�D�(��*���cuWb%C�J�Eq�;F([kJ���q�t�To)�أ�T��"Q�TDu؇S����(	5�
7Yq��UIQ�D�E��RDQ�UH�4��pM�e�I�EDHX�N9R���#V��䘜���뉑��kq+�7c$��e�"�N��pK(�n��8�r�:H�-�mQB��KH�R�)#M��Y,X�v��:��̍
�kQZ���"VdBQ�Uܬm��D���b)X�k)+i�+jye���$lC�e�$;RD��`�X�ݭ���euKj*�'$�)j���YIkMĩ[I��qE+�-m�Y\��"���+F�+c��D�[e"���d��4R5$�:D�J�Q�Z��d�ED�)A[*�UK�薦�4ִ������%Ln�js�eKcI;`��x��J�ė��D��*��_6�چ�K�U�W"��ښn� �5���Edlm4�UJ4��D���;H+\j�`��i�W[�&�d�bh,m��d��֢O�NHň�Gd�]�H�+^H�bd����ڱJ1[UN�`9�K&1�U��;k�Q�$�X�4(��Z0�cn�Yeo��c�����!Z�E"^�)%�V�D�-q�V�VF'$��P�b���&$���'T��H݉� ��
WI�*���u��U��2ܰJ�D袑��E�8�r�F�_�Z2��ej7$MȚ�N�R��R��,NUm��CI��m�%+��7EqV�i��;S�YZ&V�n�B"V���;�ڿ�j*��*�wv������Uj*��*�wv������x���b����wwn�������*��*�wv������������V��Z�m�u�_<�̺�8C�_g����o�톫G]�kYJ�T!:G-`�e�x��Pj'T�n�\��hi׊�

L�1W�8H�*%V�X�����Z�iGZN�.ZǑ��\�LE�FK��HTKi[��q� �$�k&%-N�ѹF� ��*����B�ێ�TIrJ; �����c�YcEp�U�R��YcIA�F��q2�Cc����R� �r:E+tl �L�"�u�U�<��D�bde�HJA�C�bʓ6CJ4�h��NdYE��D!b����� Є7�#*e�Hu̙"�:VQ�+W!-d!쌋1�Y%nA�;	�lƈHA�2I���H�7]�n��ܕ�Ӱ�u�:�L���EP�[d��I[�*�(�*�q�%�C,#��EW�P��&��Y1�H��F�J��R�j�T"�)U�G#r���J8I��vF�dm����)#�I.V+F��V&�v�*)m�޸���G�$nēme+��y*���̍��iT�]���X����hQ2��mI$�`c;����՛~�J��p�n�#Ӭ�Κpp].�y�C����xw��~�y�2S��O�J˽��o=�y���孴���*���S�����d�٣�2{ܐҮ���r����?^��}r�Ã���[���JO��2��Lk��GG��'$���!�����A��^@�7{����ۂ�t4�;
r��&ɿ����m��a����eѤ,r�Ys~�����d��r3V�!{���#�MK��[>�"%?�m��̺˭?���o<�:��e�Q��MF�P�b�Z�I!�ˁ���nGF���v��"�{\_�:�x�AU&]c�$����ͮ+�+��56�i��`�t�g4I&G2�֎�9�U��Ϯ�>�4wK�������?0���ˈ�g%�ӕʲ^0��7���ct�gJ��G�����>2�4�/�[F��ǄD�4O%i<p�O]��8H�dX4��!	�8>$�HL���(�*�����I�<���[�c��8�2�t���ɫ%	���2��]��w���pp�1'��6��6DԶWm��~�Y
A��DH:��GJ���6��aᦛ� Ӽɘp�5`h���Wq'Čxi�
l頳[S�W+�V�:�/2�N:��y�D�<`�i�0�åmv��^՝In]��I$#o�!*�<�x�����&`?��o=`�� ����4RF3}����SkE�X.-	��f`4�ɡٷ�Ӂ�˜� p�QE�*�1��v:`���d�P����ll��/�Y$n1bz<�Y����|h�e�:~�"h�'��4�8r�%i�$�Q���M4��2�ō$]ۑ(r��4�I$�K�L�o'��p�ǅ���U��V5�J���G�e��gG�s�9����ϾE�oun�=����4���_Z�Dk����vqz�{w[�v��_m.pk��ҽ���W����A/<{|��p�ήW�uνp읝���(�+��vp�g��o{�}���}��)�y��8�ްt�v�0�29Ö������?�C��!8��z8�$t�������̘�!#���ތU�rhi��2�Ӛt0�Ǧ�$iu�B\Ywk�����bXQ�GG�68r�9
���4�2�+e�um��μ�͸��ӄ<s�15��#I�R�W��<��|��,��x��d�[�i���������o~4I�[\j�_]���0X�hz������|�84:��o��#!4;��ۡ���� jĿ��LD&H3�=I����#����56&��AC������p��0v����"�?q�{�������Y
4D)!��D���&��	4�8QS��U!J��DXZX�NA,1��mI$����Lv���o�F�|0�;�	?��>ú���DP���l�@���Dj���6Xт@�N�Ò�:�p}Lŋ�1�m��GM"tzs�ۜ�3Z�d�l�8��<�S,rt9�MS��3�2�P�4���4ہc��SP�����LLB�6��!�|atX�/W�l��N��D�0�!��t�����ΐs�� ����I&��7�Fdc���l)Ð������B���YN]��Iɤ�>�{=���M�6�Y��N*��>!4QM;�͸)Άޚ(0����;F݊�So�4�T��V�+r������i�&��u��E7D%Ipy��Y<pӆ"~<"&��`�i� �yđJ�!�g˧�5�!�y�Y@^F��6p�i$�C�t�~d�����uQs�z��uϸ���v����>��;;��sux����tg����#���r�3�C�m��9Z��K��ᲤS�|=F�f��}���:���?���ӻ�MsMv�ݻm���<ka�Ņ�S�މw���y�鳛
����O�RNq��8��ɧ8�U'�h3���
%�|� '̊}�Ԯ����`���4p24e�<�	8b'o	��! A<�c����g]��,���f\�8�824R}���w*�`������xB�x�����im�����l�Ƣve�)����e�CI	煋�hB�!�8S���"h�&	�����:z����q(��G�*I$�s9��t˜���g�#%��Y.}ܰ`����Q����{%e���w�ᨲ�Y��(�a0i^|�U���u�#8#.�7���<j	y^���y�mb���[�$�l��Κ+G^#eP��N>$���'�F��>�A�W�t�����c��8O�L'	��MI�y�	��&2��/	���2`�	���i��i��KG���an�M����&1�Ld���'�~~$!�x�ǪK%��0C�
(���K~f�&ӟ��<�������y�b�����ao1�ȴ�Zx��x��>'I��&	��8pS�a0��D�CL!fD�a6L�!�O�t��!�0tL%a4K�D��T�a=r>[���KK[m�%����Vp�pp��������0vC㌚�Se�#r`�J�["L%L�d�{��w$�&�%�%ػ��Z-2�O�зei][%������<OgO����$0p�X��Ⴤ��L'����X|����y��]�q;	w�N��E�Q�4��e�����&��g�����t����{=7Z���[nz�9����m��)繳=�{MF�����ԥڈ��n�D�	;;/YW_I�0�W��a[��ӫ���<�տ"��r�*�MJ��}��zwɤ�y٨��˛8w��q-�=a��;�Un���ӋV���O�s~^=���~���l�8�%W�w��.�����>]��O3��ގY��Z����}��?�Y�}�����9��?o�o�-�{o���W���<��]�?���~������8�ڣ��v�ws~�ߧ�߿*�*���`�{�������]��߻��g9ϯ�G{�w���������-�{��s���묺˭:����:�8��>,�
��mEEEhH6TJψBB��YC�
`6�E��&X=X���B�&��
ܕ�}mҨ�b�Y^���%&��Ĕ��x`�l��@�C��G��A� R������.�.2�o��u��&k&�@���JS�^)�O�E	�F���!�&�3���taCdȯ ��"f��*0�i��U���P�l)<0����^�5R|d�QR��869O�<Z�J\��wf��H���> r���D��t4�@�(��m��~~m�\u�[u��xG�tA_�lf��).��Z���s����	
"V�¿Q( V��Z줣!��0����A	&fp@�3�^^�$��7�OI��9
��ƥU�9àn#�>�R�� H;٩%�X�-F	�GpR���J�L�"%�@�S�2�c �����(h�0Q��@��}���$!؊(�q��h�6ۂ��$���M�W���P�`S�8�L��)�w2�)����XU����QǆD�)1$+,櫥����cB��w��`|Ñ~vQ���F"Z]��<6CK�Y���D�4LCO�Q��v���(�̷	d^�2g,3�������sl��ݬ{�"���1���M�;�O���^��U�f}O.?maޞ��0�Ǜ֏�oK��Kw���owK��޷��x�}y~�};ڮپ:٩�4�Z���ٕä:�[�(�w�:W��Xx�p��W��O��I{��W��b�X^=�}y���$|ٔ9��|�f�)�>�狶�W�{7��w*e��:���r��~��J���3�;��h�=Ýq.�w���W�F��m-��c�q�[�'��+�uQVB�V�9QUچO�G�V���p��[�48 >aC���#gV�1��� 8堃���ޏFUZ��9BB��4%�l�i9	@�`|e�6�8h��,��� � .���� .�qG� `��.�n���0a �T;EV"��Y6���f�j���'�Q�P��	|��aCF3��|p�"I
b��b�yf��Y�b[�30�.�ύ��L00��@�P?,��40{m�`�MB��L�E�69b���U4�u��y��6��&��hi�J4�Ϭ;�W���/�U��!D�T	 �cF����# ����B�雙�D�73 �F_�ۣn�mҎ�V��fw<ό�:,���(`Y����4��H�L0�c�!+�Wb�PCQ��D#Þ*����(LA(�t������xR<a����h���b$t����J4�r��݊�����x�|�Q�#�*Yi�!c|HJ�\�=�ʫuc0`�Dݐ��\>`�b����$�aK��鳶"�)��� pb:#�.K�M��t4��į��y�y��ߛy�y��O���x������6�I6{Ȩ��	
/D�4E��.F�y��i�x�BJ��+���ۑ��A��!d�h5�ilL8h*� d�0sK���*�UVS���D\0wԛ݉LY�L ��$
A��cM`�0����2���d,a��.��LϤb�ts�I�)V�DY�ɤ�H�� �,�@��5�G Pŭ��.�*
8��@��h�1U|�uQM+�iP=�ى�a�ãC��)AE!��) ��ղ�p���t<H�YT�f".3q�9����E�7\.�ذ������Q�#��fI(a�H�G�Q��6?2t�ş�'����O:��8�]~a�V�'%\c8T�IrpZ'c�5$j5o	�}�EEhHQ?�WMQ!dS5���S��G����|A�����#A(1!h&�៥߸?���;|�Gӧ2ػ�M罔����atN�8a��kei����~�R��ç�����I����j|�Y.�P��$������J�h!-!��	]u_SG �eE}�w/���V��F�ᑁ�:��0L�(���u���3�-��t���2��q�Q
�Յ��*�+_2n��z<tl2�6C�Wߖ�#cL7R���1�I5J2�ھ#h�ˏϟ��x��"`�iƘQ��t�Qt_��M/���!���[�fQ �ua�.�g�.ML��clm�����s��x�_x}	�\VE��r���m8�n������\���w��ἳ{%��N�\�7���pR�&�A<.�}8|NA���\��7f�����D^M���mQ"׷���ͯ�W���a�o���G��ET��=����������O��{��v
��t�J���)�Z4��]G��akՄ��]ꏊ�S&cp�I+B�������^��]�:6D�����!���D��h�p[ O�)�K��H@ns"hՑB��f���E^��K]��^77Z�,tR�xm�a�EE�`W4��N\��丹��r�U���F��0�9Y�&A�l$�� ���(��
C���C�՛�4�&�7����-��%3�y����n��I^��w���w!(`�m�4� ���A���eP:�m7�|�<�+HdÈ��.����?6��:��8�]E�����U{,Ȏ��� %OHX~,sHX�j�acE6I3��g6��}d�A�ɃmUq�=��KÛ���+9�]����x|P�7,�k�Ţ��C��P�aц�9�(``�C�1¥6�I��c���2��xs���	���m�I:��R�h�D�+�}�؆q��%�)�n�X�v�sdx�7�;	����!$���C��͍s���Z�6$\1�e�'M�.D���a��ƌ�;�F�� ��D@���3c�U�wF+�Z��ɆQ󬭕�>[�o<�<�:u�qn!��)��Җ	�R!$�Si*݉��Eclm���|^�_n�=r6���"��8e�n�`L�6��4xs�pSc��hh�z@<49�˽lp��$�E�2�za�h �:�)1���^�K�A���%16@����{���m��d�K��f9̬b��f��8���Ǆq�c��ۜ4@8�hz(x���B�P��h�,+.j@��6@�(˒�����1�&r��4J�A/����|l���%��>T-�e_7��#��!�[t&@� ��G����0�6�/2���~m�u�:x�>>!����inYp���CU-Һ>��1�`$�����Y,-9��#����� �#!�պe�y�,M�8lpA0@��C�n~�G�O]�����oa��A�f��u���3����D2��	�#�����@��5c���,>Л -���i��Ji^>i_!�|�j��db��h�(:U��`׺�Q�Ґ6@��bcn j2�
"��}	�pZİN~h����v��l�t@�:����0x����5N�R�(�2i&�1C"dn�;�-�e��`r��\!��?d�NI�x�	G�=+���0�l˘8hp�On�^6�ey�Ŧ�b��Ė�KKy��mlm&R�"Ⱥ�]I*�%].�vf�]�N���r��q/�h�-[Jݦ8�N���b����h���b�-��~N���+G���bӫc���؈���Vͥ�ť�Ŷť����ZZa8B�	�lp���~>�?òZa������Ԓ��Z|�KM%a�l[,[Kf��ӫb�[+L��	�0��Y��Ã��0�1�&��ӃZ0M	���0tL:ẻ�]nvrN�;�'q.�]�K軜����]�3����KJ���Zm>O&d�{�u�-,�0��p���af\�L'&d��Z[�-�[J�2��,��w��%�.��s�����~#������N�Z����w������w�Ӛ����9�E]��[�WN��=�9xw�]�ս�VL=��)z��e'����s��|	s��l%��iD3� ���I�gf4o<�pO��`x��FŦ�#S��8��l�m�t�� 5FO�w4���i¾c��+�fs��wI�w��Ox�J�w�x��a����O��Goؚ�!"�S�}<Ez}7�����ߢ"/�R�:���ߛ]~G=���hJN|鳯���r�����gۢ�ڋ�m�W�Ԏ(!dX�������A��ԧ��W`�R:Gdl���[u��ۓn���&�-�L�ߨ�ڡ_����+K���߿o����9�?�������V�_߿o������s��������Ҫ��������9��>�������iU\Y�����9��)Q�Q�Yu�]|����:��><<#��1�ӵ8�tI�Ț��*��Z �'D�yI]���ƭp��hr��VJ�ʣ��Ҕ�5\��(Ӣ�<QR�����"�B�!GJ�*ljVY:ՊHd��Hn8�(� �:��E-̱Q	�9I�T'H�i�pIB�a]i��М�2�Q��%u���a]����TՐBH����X��bm$Œ�@������\M�cX˒��T)ji�Lq2Ң��W%p��$�-��&HIldD��lL��I�crʁ̰tV!K��ed�$G�"a#�Q�-�c�`���q\���!(Em�R,��@��h� �UI�DXªA5aJ�[�v�E#*%��b(�H!a�b&B��,���"Y�$�z�V$ҊiS��)dr9%�ղ(��b�YRmXXV�BTe�ʔKI��ʭb!R������$p��	Z�jM�e��H�mq
ڵɦ􋤸F٥�m���y������i�"!ʛ�������bn5�QUc��X�i��5c� ���6�l��h�#N!9RQ)duH�24�-J�7D��+��Z��t��APn��%j�e�mRT�H���Ili�K�MZ�n���1�`$�̝ߍ+^�/t�n/��G^}����p��=9]�J�͗�pݞ�r�fo�+9m	c�7t��OT�ew����h�1����m,u
���i]���g;�������=��ܞ]�Z���Tr�k�^���o�o�_���Ѣ!Z'e ��VlR�BFCXQ��� �.��*�n�,�-��&H`y�a�����oN�J6GD1t6Ī(,���o�IƍG���ч2�9�4��3'�(!Z��:�Hqs��zt0l��t`��A��t|�ڲ1�h�CA����X��Z�{6�_�$������B�	�Xl��P�c�a��ƕ0V���&��V�97��d����Q���ᘌ���C����t`��2wy��s���AÆ���!dp��
P�|�$�h��1��m��]y�ߛ[�:��8�]G�vq�l��}��f�|9�S�*�i��h�)C�H�(`�	��a006@��x�KWĪ��+BB!M@�
� 0ď���r`Q��!����P� �!����R�F�=����6�_4hh0�a�E;�_����5�ɀ101�����|0� ���ĥt����FY�j��;a���( BB���>7lbۢ�jm���է�$��i��� ������� ����1�/I�2̫s.P`!�,BPo@�mx£6���	���C �y���	����Sd8�d�t�,B���R�l��2���嶷�u�q�N��-��CqJa�������m�"�(�.8�8�J��y�U��#NZ>a�	@paA����8�n������l�щ����$	A�jP��Ev��QJ@� �C8�^���˳b�a��y��������Ig�P�|5�ڶ����m�"x�2�^��&k����ꑛf���>-��_�<e��vU�!�bX�@�D�y�P��&�aO�9fA�X�4]��Ӣ7L��K���xgDǁ0�?��O�:&���C6��l�&JxŢ��w�>��s�����rU���cfhiJS�:Y�[ y=�a���$��)�G�c�����E�0��/̺��6��u�q�N��N��W�{����?i�
B�#�M5��ܚ�c�@�
�~>�ƆB���t11(�Δ� M�6;m�d�c]�X�Pd����M�R�����_�m�]5ڮü���n��ޛ*�	��Kxll�Q���CM�9Orf�B�#�7ھ�&�vZ0�Lz?1�F��Řc��:�(�B��v�A)�봓�&Ur��+��]�W~7�.�z��W�Q0�Ռ�4`x���B<I\e3�����$�����4868�������qW0v���DI�m�r||ʅ� �F�cq��d�G����+��a	!�e��a[�%`�̰�m-�_�-����<�:u�q��9�N���)�F�>�]8\�T)M~�7-�4�(�!���w�-M4ӌ`$��zrOcgهvk��|k��ǆ�ч8w�{��f��l�M^�޼�9Yto���e������{�3>�P���6�{g�����L��;��������osۨ�_9��{{߹�wJ�_E�o�4od��]�K�y9HQF��}������^��o�S��R��?�P��(.���R��v3���p�
���.
 �),4T��<��P��
�k1˶��:�Z;�X`pPb,H��p�s!�tb��,4��m�IT�l�!"�C�T��u^o4Z��D�K�>�!��Mm��zƣ ��ii�4�,�p�p�T
��I&�`bA�i��((�G��Ԑk,r07
���@���҉9Cϩ��CawE��`ڭ:�?1,�8>���d�E��)�2cɧD���3���=P����Y*�e�»�!�����ï4�+y���ky�^y�t��kW���U��11$i��eUe��P����i��h�cX1YE=�,L(�uG�ѱ�Cc���=N��ʘ7D�D7Z�E�EYv�\��1H�ht�F�=v�K)�$6����c��umm�C��uP���a���h�!� �����I7��`�2A3��8���k���ez�����Nq�k?��
f�P�b��;}�*;b@0@#�T�y��t�Y{Q�(�p`�F#<������Ƃ��c(r@��:1$�<hКH��E`t�:x�l���~mkyמyǝ:�8�J�S��]vr1�c	 ʹ!?%[�#�4XA��W��aL��23�`�fXDR�4��*��]���CІF� �a���a�шd2|�I&���&"d��n	�����>����4Z! ��jG��E��I�5[)>�(�T���Fh+�|�aV��(�P��!?eX���s����4�a��AD��$���A�F�n3@����,O��S �nF��5��+"*��C�;�,n�nQ����C�
�HI�
����&��5B@�(����°�=�V��E���i����mkyמyǝ:�8�j��c�L�x�:8��$�v�2]9�M9R�@�Ѷ��=� ӡ���d'Z� � S��,r0 ��i�;��a�M�5�HE��}���.�����񰯊>k�;u&����+�����6����7A�E��ƴa�Z����2I��j��t:����R�p�ۖ
$�#��a�|(y�L�M�#� &�#�E2�ȳ���I\�ɷ&gq��T�A-��� Y��1�M)�� a�N(l �s�-2�Xpp>��9섘�<���!�!u�)�V06P��c�C!���<��6����<�ΝuYƟ}�e��8h�+�N[������u���nMj-�}���1�`$0޹�|A)WHTC��s�T\����c����f���L}u3��Y�{�ǻ!��>���s�|ث=�)�,ೡ>$�9��Ӑd97��x�Ϗ{�s\%U%�K�A�k��ĞɮO�]�����K]��A=[7��{�O|��#��(��^�v��v����"�N�I&�����Sl��{� 	b���!�b��r��Sb�����]�n�>=�&S~�I�}��PHS�D��� Y�c�>�]�������@�~Ǫ��6:Qе�;V*��g���P�#&���Ik���cō�5��C��6_B���b�"H�at&�E!�IOrRj��8�рrD���4@��#�I�90��pm����$_PQ4J�e�	r�_���:p�v���q��RqY����?���F��?3D�0a4�:��~ioϖ����<�:u�qf���s#bϖ
QL���!�E�@�&�Sq�c�H��H7���+���w���Bj�ã�H|�eV��]�
�E&��͗MB� fM"��[V�vVʾ+�+����	�~wf<O�C�� ��M����0J q���)�$�8`�{�zV̄ X�p}	H4��3�x�Aѩ�	�טW�P���H�UQ�G��,�ӇCN�CY7�*�SesBR4��=�o�'2������P�n��ƝXၢ���l{p2LI�w�cȤ�O���t���FOd�'�Zxa�p�[0˘&�p�y�l��H`ጳ�a0��a�c'����gdk�l�L�1�+d��M�.�ve�ݎN���am1Y[J�-+V�Z-8�n�Դyl<���-��y�G�m���[L[l~E�1�8��|�M?O��`�`�0��0�8L>�E��	�-�-�%���b��[,�$��a-9%���|�O���X����I�KM4�m---���6)0���a,��a��a<L&I8`��NɃ�p�����5�~%��Ig��?!�ѫ���$&I����q.�%�]�N�ܺ%��iV�i�B�a����y�O=��<O��	����I���>0���a�c'����gH�0xCĺ��2�Ļ��N�E�IlD��2�$���G�??S��IEӟ�E'*�y"�M���s�~��{�v}9�/7�m��suo~|s*�_l�_{�*8V�����g/�2���=�5U��1����N.|w�y�ֹ��.����M�ƾ��ZS��}9�C�8q��TWG���������\�՗���|�Ǝ�K��Ҋ�V������$�]�?"�yǕ�����窽��8\�L����{i�|�{�X�wP���;�[�O�'=����g��U|�_ݻ�������ߺ��U򴿻ۿ������ߺ��U򴿻ۿ�������֫�U����g�4�i֝i�_-m�o:��8�]GPM�F1�V���ܚ�]$� \��%�֙	40�P�Gý�bp�@�������M�$ d=��{U*��vA��m��6A��g<����s2d��l4� h�0Y��/sʰVҙ�YV�S�TdR�t��f��B��çF��C��	4h2?0,��#�Z�ct�R�j!D�с')���c�~h0���$�{<0d��
 ����i�A�	�R~t��Ӂ�~h,���ÃvW���2��h�O�u���oͬ�&���hi�0�Yɴq����kB_#M�&����QQZ���3��I4���?n\����D�ݎ���6�FG�`Bz�D��}��CN"�9ŰIn���ɒ���^:����;H<&�F$01� ��	4�p9 Q^L��Z8tR��([̔	ೋ����������n��\�`h>#8����c4��޲:�
�#$��r��BQ��|�����5�Ud�%��rtht��80�(�����^m��ֵ���8�]G=�fJ������vǛ6wc�:&�;F�4��V�iy%:��\��EEhH>�+�l����k����g�<-�gI�k�y�g;�o�&���#:�/���;ϼ狣ٸ�><w\����t���g͚s3�߽����޻�~��g��E��H���of�������Nur��w�����:u���rէM��6y�}�[v���}�ߡ�M>&r����g5�i&�i���	�~ąG�9B��'H\�=�d)�P���%j��	I�!螼֭�Y�|4<3I��nD��h��laL�n��Ģy�r�U�*���;�ƀ�[�!���p� >c��F>3�t!����b���d��$O��<��) ���8t�S����t���?.x])yU�y7F�.\ʁ.���WQ[��I�SH�jmYV�F�[�#��0v�w�h�`�:ˬ���o��-kuo<�Νu0�I��MµA�Qq�z���T�@2�|>���<��,�V,���බ��Қ��Q�?�������{y�IR%�7:ӡ�Ў�2B[��uWf�-�u�]�(dv��(l��O&��0h�sH?����"�?A�nq�]��{���5�oS|,CrN���+������M�0}�䪅��/rB-4|Wt~��m��_~�c�+��u�D#����.2������Z���x�����?�Ň���2��i�n�QQZ_s!�&�;	w��8�c���ӑ��6!=$L�!nH�:Ü�bY��}�\{����j�1��c_)��a��V��S�|=�p�ij�������F{;��t!{&+m�w6�e�V9��(�}��:&`I���sP�� �:f��&|_����ٜ*Ua[+���]M_�N��-!Y�GC��Kl����l�g<h�o�qk[�y�t��޿a[e�5uJ�	!{��o\��TTV���!��Ύ���W���!~���j͸�.hQ�����pm�;H�^���.��H�
�*�]�yΨ��"1V0����}VQ��!d.�]~�s'��<�4�1�X�s�Ih6ǌ!�n�1�!��D)�Y�I�e�ܒ\��G�3U'"�,��P�����rB׬	��c�'�`l��D8�tB�pXlv�ѐ���8�O2�km��ŭo-�yӮ�針f���v��4wAcJJ�h�^�*��*�v�v<���EEhHKͩ߷��|�����a�i5�I��{;�w5)�g8�L���]��Y��K����!�N��<��:xK,�i�&��{��F֜���w5lo���9�z����ϝS}Ϸ��zdwWR��g+����o��}ι��Ft�[�n���!����	��J�ɫS�烃�����Nt�:��ca��Ц�i$�4!᱁�S�����a��C��Jl�c�kZ�P����-��̆\��X�Ҙ�Hl���O��!hP��~�^����Ÿ�N6ht˕���56�S�$���>ˀ����K�J~�=BK��-9��1��?y�iC��k�u��H�SJt��ͭ�ŭo-�yӮ��{�B��z�bm�W�IU����yJ!|���x29)��$7��G��^J��8�U}�G��k���)F(�N��C%��C�HK�gp�r{�p,�C�n8�s,ޱ��L�^CD-�g!�u�ǃD8x��_�9�?�N�ѩN���q�n��d��	;T�K����Q!,�g�u�h�O�M���8�!6�P��B'�>�ry�U���Bf�e2���;��!���!�p�8[�Z�[�8�]G�i���S�J���АY*C��zX���GBf���la��h�����B�/
��Xh�4C
���T�d����Xh���2��k��-�����>��â8,l��DWc��YsLm�	$k�CƊ�uS��.q(9�l��A ��e���Z�G"�z��9ߕ�NF���O ���Ig��.~͙ćnM6d�#��0�t0Á��d��XZ�u���qk[�[�8q�mk_���9;xjfW��;+�i�^0�h*EhFVÜK��m��А�5�j��k��t�h:C8H>l�m4�L����WW�LnM`cR�A�vC.}�<=� Q2�[��&Cn��(� Q<�����h��D��]O����clؙy?w=�f��&N��k٪]�9�u �چ���3�f�C|�\c�U��3�$�9��{�DG/���]���n���?xwXv]o��u���������Oؑ��y!�p�^\p�&��φ�L&	�0p��0�tː�x��0�L<��crq��|�K"ȲUԑiId�H�%E��e�.0��VV���ZU�ah��ZW����4�J��ul-�-<�G��Qkb�a�����[�u8�K%��K�8L'	�����I��KM%���h�[�ZZ<�<�F��[,rKa��m->F��ϙ���~����?�~0|`��&��F�!���;#���!���;&h�0�՘:��/D�ƙ���&		��`���D��|'r�x�˓�y����4`��������0���xO���c'�у	��2�&�ra<`���#�0xCd�`J�]����q.�w�]�x�F�J x�G�{�&�ϻ̣{��y��y|-7��#޾�C�:G��#��'�.��Q����Ok)QN���!��l�����D��ti'G9�K�*.��ϩ�t�7U�Ks��_�=~�<���?�Ox�F=:pt���	����JɈ�	�Ü�͕���>���D�=����~�'o�>�����:mw���o5�J�o=^�{�__�f?���Wo�=�ֳ�$�o���_�]K�u��>���;�r�2�����!Xӧ)�1�ֵ$F��V��x���,�S�zwT�����U��Z[�;w��ww{�������W���o�����n��j���U����{�������[Uz����o�64ӆu�Yu�Z�Z����q�'�ɑ�և�c������!�U��r�Y2EZ��h�"���)%�)T�Ic�e�n�Y"J��ƛP�r�V�]C�i$���H&Y%�"��1LM�mK6C��\Y`��d�Kk$��I	I˕�؊���Ҋ��n�!�*R���;%�TJ�HE�$��c	\U���)J2TF!�գ���J�r�+���hd�l�&��Ѷ"X��l���&����ErW����ۨ�*�R�D�L������uQ2��d����q����KQe�mAHA��o&*8�Q��T1QFA5S���I���!,	�x�Fe�&�(<�2�y^*"�9D�JQ� �,)HE�T�T�V�IKi,V��I-u��q��*J*���,*�X����bI5cE��l%�RF��Kh8���pj()[BP�M�D���o#b�V�1�µrF�
(��V(�,VD7�@����R�64����#����HeNQ��JH�Ci��<�1��W1�ݸ���j&��<M&A��mAQ��kJ��n���7�"����$�DPj	�j��VT�,��EEEhHkY�a�X��6C�Fޛ;���Noo������G���Y���忳�O������A�����8"^S�FoN��������<n��N|n�G:����Ț���o	y�ogx]��x�=ͭ�ټ�^f��J�eP����O�4�BT.�?�t�?�+6C8v>rਕ2G�I�&�2Cc�t���}�b��6�G+v�i*���;B��B~9͞���s��^s��<x1�)�a�a���^�{�xz-͎���8ѾԪ�S����pv8ˮ��eh�����F�<0,8X$4QP�^i�7P��
*�4�2z,�}<���.ݙ���`Q��i�;~i60C&6`��F���ַ���p��޻��M��w�9(�Â;NA'�Xt���lm�TURQ������&N;0�w��9�	��~?�w�[$QK�\8y������ �gL�8!��:�e�B�v[M|BM��p�l(���9��B�t�`��	�8l�����os����q�Vmݥǳ��f֭ԫ��i��v�e���;�S�ef��~�j�na_R��%7�]v��n6�MEŝ����iW<�W��|��Th�(�N4��y�ߖ�ַ���p�����>�c�hI#w�7ޢ���$/�!5��T���*��4!�;0�j���d4�cl��'x<�i6f��ɒ����0��b|��]��ˊ7E�'&��Тu�j�ֳ�I�o\>�
�}R���4y�����&�D4D�$$��h!-�l���aC��<08C����lpC���#)���Q&��!���O���܌�d>��d�dy�!�c�cfG�6��~u����ַ���N�N��R��7�GL4]��D�e�t���А�H�?U2Q0d}�"Xl���S�8��!�������٦���b�Bͼ���lrq�!��k׷D����d��@��N��GEu]�h�8�3\.���_=�U�Dǳ��@�L��:�p~�LJZ��HGlz�t8�9�������p!ిv�#]����]Yustv$��29�f�;y�%�&��`��iכm�n-kyky�8����3�S\Dul9Q�6޶�o�h�#P�$���k�T��;��m��А�4o��7�����|����\�$�\�pn��;U�|w�]r����4ޞ����~�~D�{)��g8]z~4���8�����o��QE��'n;-�S�����>��MU	rw�s��O�S�CO;;�]�O��n�EP�ET�Ï�ȡa�Ä=3��o��2��~6�@�5�넯�i�����WȵeQ��������_tq��?��8�h���=��@�4�cd��AD#/Č�p�ç$6\��P0�O ��^�O�!m�)�?�g������HT
�h6B�� �MA�)pc������ �_8���8��:��o?8���x����0�f�,g��l�kz��EEEhHj�V��u�,8BIw	��Tl��c��!��WE��rP���Kn`x;c�XB�i�G.O��C�>��Y�n��.�7�d�
!��c,�d�À�&�`�\���%�p��B���ZZ��]�#���ez#�π<`�ƒX�K!���7FKx��D�փ� ����������|a�y��-���?8��ַ���::#�����8UC�j.�z���/�TTV��v}�,�&��7UAT��*��t�0�����8Pb&?Q,Kt�e̐L�G������\d'8hMŞ{������D8	Z��|Q��n��"IY�c�ڗ�x;����m/�tw���c[��S
˷`��̹�&C|&��Q�ht{rX�9$���7�|-zWò��!��� ��]sg�	�U���#�U�`�"h ��*��L������3��0t(�q��y�֜~qk[�[�8q�l�U�VS%ˀ�.u�EEE�������i���x8: ���D��N?�UY�Vmۻ�>�B��gC�̞8���CCh�ܑ�i�Z�D4�a���	�}1��ʓA�g#A�B᣾j�]J������j��h���Z}P���ռ�$n��k�XF1\y�u؉%��8ѧL�"�e�<��m�ŭo-o8����ϼ��=[.��!�$]��:�M��h���	a�8s=�F���W�������F���'E�||Ϲr�F�Å~�&z8��ۨkf�e�_e��`�,��W��wh�ʢT4\��oN�����<5�s}7HT��_+�ϸr�����$鷮o���F㏪ꦝ(�J�.�sǧk������l�f���S:��X�:[�־r�x`�$��|�D��6�9�L��1�Y
|4L`��,���?��^��1�q�AGt�?�$�����G�`|��&ä;���Y�2|���:���Pe��xi�pk�GI-�Yxˇ޺���<`���D�?����7���l-��v�R�bi'���e3�CC�K|�P���&�jF�T��|��~a�y����kqk[�[�N�!�8x����Br��$TIC+p�*����	7��TTV�!`��:�3%�(,���?8t��v����Ņ���j�J���3\��""I+ݼ��3�WE��C���۳[f�$1����&���2���!��h�a|SA��D/��Vؑ
�ʺ�$��k&�MV����~>!���0O`��0C�?X9��&HZ����C�y���C��6t��X�p�C���0DÂB�DK�&���tD��(AAA(���pD��<&�CD�4MD�4MD�4L0��h��<�4��4J(N�"&�&�:"t��'D�� �,DD�Â�D�:"&	���y�O	Ӆ��(L��/2���x�ǋx�H���[K[ki�^e�.�ˮ��Z�8~���K�&���!�t��AAO�!E0L?~������{d��.Y�5ۅߧޜ�����*��+�	5zl��{�2+,�ӛ�xp~��1j��%Ua=���N��w�m��+2۟_n�u�v���$>�sM�>=�j:��Đ��_{�l���)���ϥ��>�D��K߽ɾ�$���n"v�:����.k+��i+�7'"�ۗ�lz��fRW6�$��k���Y�,�no����{lk�]�y���ʧ5_?��}޽t��E���C6e���>F^��ҨWwU�j�Ux��������o��UmU��ݿ�����o��U^�ګww���www}��qUz�j�������CHiF�p饝un6������#�6�����/�EEEhHY�9wu��z-֬u�Lxvq��C�a`��׍����+�Q�1�n5�NÈ�hMzI0�1�;*F?nHBBX���8C�9���+L$� ���k.���$��N�/��/B�Ͼ�"y�#��n��QNU�cƉ�:Dv?:˔���a��v�Q�tt���2]�$6��X�0Q�a��|�N�<�o�-kyky�#�8|s��<�X���k�����EEEhHz���e2�	�J3[�������&Ma�(v!�HMy�aI�9�o�Ѱ�
2�c^�f�O�^C}���Wc��^��|��D>o9��J��t��d49��L�:eɚc9�p�h,����s�1��;⚁d/g8��U]P�=����Nm�h���(�qYWUs	"r�5���9V�!�o�6�G�w�������Q�������~[��ŭo-o8�:3�ŧ�aÿ�#�J(k$� p�e&p�pb;���;���)5�!s|���!������޽��>;,�>����������_���O��u���:x0zo��/2��9]��ͳ��v���f��Ǵ_����W�
��3�]��{�>����z%�Mr2��r�rw����3���'���c�������[�Ӫ#��a���$��uON\���B�Ȟ�6��vzy�I���!�#х���#!��a�� ���Z��HI�4��W=Y3���fA��썾���넊�.GL~M�!�I2:����:Jp��C�<\v�]Ja*Q��?��:�M!�6:��:�V��#)��L[�$��0>�,�ꕧ��9\mF�u�_6����~qŭo-o8������fz�]�J�/s����	I_�Q��GR�V��@�Y�(yr%��"YC��4LO�鱣!��ƞ�,~|�Q�:�:d#�[��$�/]���Y�ý6t����Ė��!	,�ᙹ��C�M��?��4s5ũ:C^-��������O�������;����)-��N�)�����ǹ��밠+�[���w��~����q��4���[�-f0��N�!�9E�7�ޅ�듒�U�75W����q�<]nDE=���CF6�gA�硘�"�o>���᠆<����و�P�K1!�f6����%��o�hڧd�ڸ-;t��T�3�}������C��c"`���
�*s.}'@':�!���od�񢪨������v���O�gD�ωC×��U7]ɥ�L>|���q帷Z����8�0ۊ{���b1����#���6V�W+��.��]	�!G"�W�`ɀ�5N���|�3á���2BJ��1���������7�ZgL�b4�������t��m�)�h�E::�M���ϗy$po�z��:�2O]�B��9��vd4z��Cd�HRv#���uӖ�M̻B��C�m�ʹ�����Z�Z�q��9���NnX3�d�z�4��k:ѥ����~�clm���w��G]\�F^Z��9��O���;���+�紪#M=]���wva����缘={W|�=�r���*��y��~�44_}���a��ҟ{�Ç�:T��k�{9lw��.M��sz�ߠ����{�����T9��y���g9��2����r��R��w�t^���&ֈ�� [l+f�]񛟌Y�*����1+j��U"ߘt��Xh�%���}?u��UL?HɄL�!u\3��p�$��~�2��[k��I���:p��dh����2�Ây>*��Q�.�pt�Bo�/�0�2e3�S�(#�����6����ΎN�^�&%��J�$vm�y��ˍ�����n-kyk<t���a���jZML�����	*�� ����S�!,��or>��:T�-V��M5�Mlt:��������4�A�[ć�,}��8|e��i��D�į�e��CK�/��,VD�մ���yn���#�1tFt)��M�f��3{+�IR������Qܺ6+�x�eݔ�r5�ru��x�H����i��~mŭoa�N����k�ɳRĻv���**+Bk!�[�z��u�A0h,�pj�ߋ�xpvノ4~��6l:fC<p`i��Ӑ�H! �QqԽ��Ҍ���څ�uF��{=o���2�2d\��5�%����։�u�U�D��j��|=��Ȟt�$��u构��:|~��␒�I`�h�n\H˓>�$��HJ�i�83sw�Sn*ma�Ym��u�Ŷ�ַ���q�q��\}�D�%Ma�!	���LԦѽZ�o5�TTj�����0����(���a�X����L�[\��-V�3�4Iq���7N)����|ũZi��Q��0>�	�����x>�çSe�aonݸ�ΏCOC�~ܝ()���h�2�E�W�q�t��%���r����_�<LJ�O�!xgu���3s��spѣǓ��6�v4<xGz!q��u��5�4��Ke<��2��"h�P�$�D��h����tN�(AA<"%p���8"tD��0L4M�4DD�	F8"CK4DL0��&�E	��D�N��&t��x�ӄ�h�b"&�pC�$��D�:B�2%�'��p�� �` �����孵��Xi�\e�[μ���ֶ�������<���tN�(AAO��?�ᤞ������wy���ʞ#�GV>O�y��rq	^�����uO7��J��{��fd�^O���N�N����)��B�IOSN���"��}���ZǇ�6F��H}�'�E�;���d}~�sP���J�����DS�௸}�P��<�L����������to��sy�8�>	��ӽ/h��0KW���wކp7�*:�����`z�������^�w�����O,�\���A�ϻ~ӿ���T{��v���d�v���/�̭��"�_<W;^���f��i�ů����(�KQ>iE%���o�杷�ݑ����ض����!"���r�f_������Y��q^*�UmU���;��wwws��U^�ګww���wwww?~�U|�[����n�����Ԫ���ww�M���Q��4�f�~qm�����qa�i�}9�̊��P�&;�;eh�< �Gr6&)jpd�r[AڑfBY"e�,b��%(�q��d� hP��)U��S��1��$r+%-��]�HB���bMJ�DǎH%^U$@�R
Z*�TY[,j�	��+i`��+E�X��WkU���$U��$8�"�C��U �"!���q��4���$,� ��ى��T�델KK�;���R2	eQҍ
V�-`Ԥ%���i�+G��C@�QZFT11���)r"\Pl�1��V)
!��#������!

�
ȊQ��-I��'A4�5^U*��X��.4�"�fm6�VZHL���
S��N,+!l�$7TJ�T����pu)k���e�HM�j��I$yY�1(�6��U*r�"Acl��G	f*��j�RE�
��mD��'`���M����%HQX�ХJ��q7,��H�"��Udq�Pq*줲�l�D�N7-�<��6���;�+FG#���n��a2�J�$��QRFԗ,u�VBKh�U(RE*A�Q��j�*eb��6Tʬ�n/�����	�r������sGr���rs���y�HЅ���&��K�p�N�����糾ţ�'S��<^�����%��[�Jzt3��{�|�Ҏf`|�Xs��wS�k��|�=#�����Kϸ�n�����>w�j�:O�9{��N�'�ĺ�_��^<����y�I�J���8��m���?�b��vN��rN�����+)3�����H�h�|`,��ѩ#�G�f��84���ɀ��9	.K*�
�`~r��l��@r9y�8��w�N�q44�����}��s&�*9y����Y�d��]�>��i�u��ݼ����f�__�<�g���#[�,,��Mm1%4;�,�<�n2��N?<��_d����ۆ�l�GpJ�d��S�����tY%+OJ;lch������4��a�a��eQ�$�|??eɏ������(��ɓ>�ƯF��kF��WWF�M�u)���$%�$�����M���t`C/�>�?/j��;]4�9[4�T�ێ0��ws��=�.{�d3|�kzq3��<o�~vczMNx�t���� �0w�`k����4vQ����4$w_+��U�6�O�[-�����\Z�Z�q��o�I[��7�#�M��v�Z�������֪J�!<=r�|L�ϪN9`p�TԔf��r�!F$%�wtԭ<��!Aߛ�A�~H�g:�4gX�N�#�y�aIDԼѪ��b^kC��9z`iۦ�����p����_�a������0��0��̈́8=髫Z�e��?~��8x'⬰��m�qX�TW9_�i��2�-���~[�-o-o8�����Ƙ%Jh��h򢢢�#��	"A�����08|l��>��8g��BK,���Ȅ&om\�0����D���/\�ʪ�����>�dl�Q�HF��6=�4x��UQ����ff��ӄ�ᰣ��d�j6l�A��i�f^��<�£PXF ��<�!����Seh4mP�?I	�3!1�vǡ�ޓx���_�!�����e[4�4��e�[qל~[�-o-o8������8Ύs�QA�芃K��5��s��s��u��**+BY���K�}�9���ѽ|r��ַ��5��g'y9b���;�e=ߘz����f�O{	�2�|va�p�{��]���8��Q���|����;et���z�W4�)*������i^͈s���ث��/�U�{�7���ַu�{N�g0Ӊ�^��3����{N��v��w�+�����K<Q�wۚ�ܭj�g9+{�χ��y��:8��rn;��Iυ��af�Ptpt:�(4d���$��K���ˇZ�7Im<I	F>{�����6d48��൰�L�RY�����������������^:1ӌ4�닩,��v�3��Iˊ�i*�Ԩ�M.ͯ�VT���^�r�p�h�[-����qkun���ua�0�?c�I�!�QD�j�6؊���r��5���5A��\$'B�߲�W��O$�"���;¶X'�o��vd�)�z~�^�Wkd�Z@�yK$�cAS�Z�m�Y�O��N��JϊIZ�IƬ����B���σ��{��G'?[%�tڮ*�O����١�f�����!��i���]��~;[V�?wW��.��l'C��x0C�e�^qלZ�[�yky�]Gl»(�9w�z���О���x��&�H��gB��uI��ri��e�0�#���� L8�k;�,�%���$�4Yߜ��g�A`��ף^E}J,�V�GU����"�%��g�w:���X���
!�2Hi���w�+afXd{�Rx��A�X�J��A���`�����H���'(��|UЏ��S��Q��[>|�0물��y�ŭո����u�q�����#�1eC���clm���2�-\p�i��_�ھ0G�R������JE9�jխ�ײHT�2�[f�5���#�)"T�5bG�Q�x!����Z~�ϲ�H�4�}��g�CA�b��h����d-y�^�����|�+Je��:�`2����<4:���8�����+�/��E���^e��帵����󎺎0ێ[Ef�N�!>!*,B�z
rR8�t(��#�I�o�A��96>ܷ[�j�QQZ��]���k����$۾��K�κI���ہϥ�g=g��+�t|*Y��s�>��hg4���駡�O,Q-�JqD�+vI(Ԑ��wi��/v�_G�x�*�o۽ꇽ����Vz�CM�9�E�8��8f�=220>Ԗdǈ;v8G��~��8��b�M�G~>2���'�d��t:���h��'C&BFB#���H�`d����h��!��h厌/Ca��$�����W��id���!�b�&�gLE�L�l�`�ȡ������r馑�y�Y~qo8��V�^[���Ǆxg	Ó�~[����k�C*(H��D�'_Ȩ��	���JÆ�>c*���I6��a<�|�p�BdY��p��U�+k��?���Q�"���`���J�)�WD$�l�:�;�:l{�`��g˭+�����ܽ\�L�6��	�A�H�̤�Խi=P��!���ZJ�B�91ke$��Y���PY�>�z�l6;vɃ��%_��u\��]q��i�agV�<KD ��"'�M�a�<'Nx� � �i�p�Â'����xL4MD�4MD�L<t�,���"a��!�8"tDL4O	bX�tN�� ��"";"aB�D�:'���k'���:!g9�(J�%���Ay��<������[�2î4a���0�H"%���?�-k[���l>Fx��Ǐ�&���9�ݞ�����IUa�U��>9+�-����>����\W���q�.{��܇�,���� ���G�t}��1���ֆ�p{9���w�u�{f{��v�{��6b~�2��.Y��.9e��~�Ϲ�I'3�>C���U�W����v�'�N�T���e0�Vo���;_��[Tq��}�������ػ��UW��U���ߦ������U�Un���黻���EU\ZUn���n������UW�[��;�:î��.���Z�Z�yf:||C�8<��TTV��f��B�K*+2���t�g�Ë����ѡ��2={�3O���O��u{O���߿h���#.Y��+S:*����8���� |r�oô0:��A�g�=I���WY��]9�b���%��H�#C��za=�l�H�Q���:�c�UQ~��ͼ��gϵ��q�e�][�q�n�n0��O��|<&��ܐ���Y�yz���ʾI|]��fy�)?MI
�h@���0�C�j$�y|�����y��,�/+�N-�l�b�B&Z�\���o�c�BH���C�u��H�EDd]&"Tjdt=#��ÆʹUɀ�h>��UQMUU{��Fg��`Pc�t���}N�+T���$����u��#li<��O�ο8��V�Z�t����x�'��NpA%��8K��(���94�����������{�y$I�_{Y=Mk�{
��o��^ߍ�tS��}�z��9��j7��/`��7��D\�>!����i���:jiAJ�:��.��9��u�i�z��]o{"��r1�-,�GdE�{��r���\��N�KY�R�cI$O8d|��~5G>���:򪤌��ގX1�d�L�'_FJ�������'�ٛ�8�w����Cca���MK!!���0{��y���c�^Jg����y&��Y��^%CTĘ�����7�Si�Y�v��I)�Cc�?�=�r�.�uT�ʕ�2�<��̿4���?-խǖ��u�u������ʒBJ�ج,��EEJ�J�HHa���c6�|�?f��!�1f@�M��M4�K�9�w��lv�J�u�qg�_I����J�X7k���$p4p�#"o�`b\��"���
�.�d�8L#Hb����#տi_6�ԭ9�xŤA�g3&���X$$y�׉�>��5��8BIR�����U�e��[.�㮿8�����������<>	4G���X��R��+clm��~���$ڞ>3�Ύ��䑰���5����ѳ�y;I�iR��}o�u�k�����	*�D�X�����Xi�o]k!��I���%��Te6:~���:c�	�'ǎ�v�̪r]�\,�bF�95ԕ�X]?��Y�x6�0�W�eci���yո��Xa��x�������Zl[�Ih�I���:�����$	}**��4�v_`����px����a���s����Ù���l��Q�çe]�n�Y�7"~S<��ظa���Hty�����"���i��u�h���� J
ӱ2bI���A>,<����z��<>��ݹT���R|��~~pu�Cm�6�-����~u�������[�:�:���Dml��}$��[�T�{pBé�Y�Iw\=cJX;.˅֝5�3��TTV��f׃f~���鳲�{�����6��p��/��w���o2���)Ɗ]��ߏ�����~菢�e���j���g�;���e���?��W�9�2{�s�'����(�{�<r�wy��ꡚ4_c9���������Ù��߫�y���b�g7����7<�x�_y;��}��<�m;�SuRH��p��]�z|8v��a��I���'�*�9�u5"�2�~hÁ8p�����yC��(o�%��Dݵ�oC���
_�}%qB��ς�͎�, �Sl�ↈJ�-�,a���P�2�a�(4Q!�z�ʦ�u�t�.�M�8u	z!b��h��1�}X��ꮚuc��^i�]yŭխǖ��u�u���EK��V���**+G��9 �;u���<�ꪨ�č��x5���&(��j�W�����@Q冹��
ز�4<
�C�fC$�^Y�� �[��h��� _ߍ#�O�X�s6�8VQl�V�\��W��Bj�W�=]�H(��zm������!$�C�������+���0�4�ɶV�ߞy�庵���󎺎�������Z�F�����\Sj�%'�X��:V�Kle�w�BI?@�W�m�c�z�,4d~r���h�R�X���!��bħ��U�z����������ʄ��K-�d�d�I T!
�w�YWW:Go�[�>p��x͉=�ɞbB�'�)$F3�4.�ܿ�ow}��Dӎ��n�noR�qhϳ�f��u��U��#�m6��[��8������󎺎������-h��u`���W��6�����xLϖ���=z;��a�\���^!U��r�܍jU��D1f��%��pn��$�����C�����!�q]���+��I'j�J���%0�J�%Qϵ۸��Ĳ)��7�`:�u�(r���U���nFI6q�|�I0�6��Ɵ�̫�>c��N?8�������:""h�(A�b"&	�"'�����e �AA<%��%�pD��<&	�i�M�0M4�0�Bo����gDDDL(A(�,DO�h��'��,K�%�!�숈�'�D�"X�'�MD�Ĳ4NP�%���� ��J�A!��~:~�
M:i���x�H"%���.���-����e�Ye�x���VE��]k^o��&{�e�m=Ϲ������l����p�9��7�Z��Nk���=���Β}�����_sw�?v�����8&�^�;��!C5e�x�S�����ɇ�t���s��s�u���S��>WH$_�G=z���L��8o9E~�)솴sF)M�gۛ���p��_uw>}���.1���N��S,��	�x���]�^�dΜ������O�����=���j^����i��]��|��%�~]�G��o����������u����==Kw�rUzz.r�o=�[���u(�IU��x� �tIB�8JG��:.���:uO��w�}�{�ߟª�-*�wv������Ȫ��J��ݿ�����ߑUW�[�������"���Un���l���묺˭:��qkukyŭ�t�!���]��qX�mP�ej��䊉�2�ڣ-�����K!AiRe)[��q�2hR�l+�ʤ��bdm+n"$������ۗ,C(�U�\��-�z�7U��E
��`�<u2Mu�[!Z��W-�4�UrY�i)��P�(&��n!��<p�X�%$x�[DB-pq�	E���RB�X2���B,VH"8R����4(JZ�9Kr�pE2�U������[]�(!R4�ƄTZ��1b��$D�ˤ(���IJPaf	V&�(Ԣb���Y&LqR.!�m!b(���W��i�ю�У� ��ZȮ!Qچ"*2A��#*N�"�f1B�b����b 1'�c2�����fQ�E*�U��%]�H8�M2$H����Z;*��#��*�;c��L���,�J6D�e������bq�b��(�[\(�����%J��[u�c�B��ĝ�X%U-�$	Uf�X�U����D�qK�T�`Ъ�����A+kn�ئ7�L�ѹIJ��*ұ6�I%MR��n�RL�Me��h��2�$�k�&�"r�4��ā5��**+E���G${�j���sN���s�z����gN�E���un�z?��wʜv|27|��;e{�w���g�=����ڽ੼ٖ���5�N��f��o��}y��������N}Yh���F��w�ڠ��V�-�){ξv�g��^U>X�Wk����i�����+|���,�����'�h�X��.L��C�Ǧ��$�Xt~j��F,����nIݾ-ˊ=�ϟ�9�p7�H1�}TUW�G��l�˧A����������%M�^p�Q^>%*�gO��=�>�fM*�%��I�+����y��u��~[�[�-o8��h$�3H���k�2�h]B������_n1���|UՙY�F�
��vj�O�k��F~�-�9��*��vUJ�Xǟ��r�h7�<�U�9������m%t7[)V!(*�O�VC�Q�R�Vn��HTL�!��$�TW�]đ$���ϰ$�}�>h��H��$��OrK�w�������tjLV%%}t��J�a6�̭�矛y�n�o-ż㮣�2��1$�cED����_�!!!,:o�t�t����+p>�����3��ݽr4|04`C.�6Uܫ�<<x�B,�>r��ǝ�/���f�Q���l����҇%Ծ�����M���܎�Ttc����P�:I8��Y��9Z�Kd$2�d$����a2�v�哯Gi�ɀ8(�q�~um�-n�o-��㮣� Ƴќ\�,y��J�5�3w�BB���̚r�� �wd�:�����_��O�5.�tR��)�OjY�3���{�ʹU�f���X�������g�q���5�����_�t��&��껅�YWr�˿�=p���zl7w.ҏ��88I$�B�r����!�=;p?:w�����^;\�˨묺ˍ:��kZ�Z�[ky�]G\e����M��k��z�)���-@��ĳ�ipBp�?T$$%��7�dQӽ9x��O5&۳���/�o]�/r}:��s���7�{E��b҇;�{=��>s�=;�.���uH���=�D=����4\�G�7���Ӏ���z�:�I:������N8ټ�!�Ҷ�x��wcK���t��Io$<��[��~�t���9-�Q.eB����&R;��)�?��?�深�mH��s�2N�|6̎��`|��*��K��od�'J�_J:_芳 ����u��<ÒD�W��u�z����`�J�VC �ű�pqf��&�������(B�l".��;gx�RDq[�9�t��ucG��u�+��$o�����~e��~y��n�o-��㮣�2��h��6[���l���HHK�F����2L�v>�u�Tn��UZ��T�;r:9pd8��?dk�B��G@np<PN; ������}�������������J56wX��$��m�J%�$�9����.I�c������X�z�x�w�`f��5���!��~v��­[2�>~e�[i�_�~Z�Z�[ky�]G\eF����,�7e%�s��oo^>�DF�{LQ-��i�{&�Q[�! �|�6�6J΋̄�&�!��.]U�ܘt0v�l8;��<���(4d����:K��#!k��6+�ٳ�l�kZI�w�\,����Y]+���l>�aD`�D���ÚM]���f���2 �Xl���/C�f�qc����i�q|-���Q��m��y�Z�����[�:�:�/�T�`���bD�)�4��BG^�baZCu�Jؓꁧ��?_���6f�^�Hr�U{�x\��2c3f��m�?7F~�[���6�ľˇAԒY�jW4�\�]{�������6̚\�R�5�~�?$�����Ό�U,*�G�"��Ѡ�4SPjH�͋�렆B�%X��|�.2��ym�kukym�㧏����<��ʮ,�e#]#AHRU�&���k�]-�{�HHK>Gy����rG�/>]�囨�?S��M*}�zM5��W�_��p]y�9|"��b7���4����i�^I�p��N�����x�p��r.��^����t����y����n���}M���{����ƣ�"MV��o���v��n�~9��F�����l޳�w;��m(�)G������O�������	��	xX���8�|88g���<���[��RQ�o�lLc��HxuގCNoHxv:a_��,�㘅��s��fsj��s鵂F-$����+b���\ڗ١��Ǐ��b��X:�<����O�-��խ嶷�u�u�]��R�S�X�27��_�BBBX{�|&�"@�������!d ���aÂ��~m���#�������+բ�W�r�	�����!bϬ[a6�]J-Ɂ�`�A�r����ڊ��+�w/�ţE�9�-�z���Á�Ǖ(����g�2t�g�pJ?A�"&���D艂&��&�'�8pAAHtN	Â%�N��'�0��4��&��4MDDM0L:P��8%	Ӣ""i�D�'
��h��'D�,K8��(��$(DN���'�DjDG� �Ț&	�:%�d8"r���A,�� �xD�����pN��i�M?��"%��M4L:'D�����,��,�f�al3�t��zx�3{��8�����>%����w0��n��<=\��J=���������8[�G���+�6�&]fx���e^#�:�ν�>�Mpۼ�7����o���v�d��*m��i}�/��z>{\|���-�7�6^����y����T��.NW۷����۹��/��L�����5�劳���[���jl���_GX��%�sk�r卵"����Z�^�]����_d;أ[/4����/޺���w�?Ky�^��϶���U�wy�7�q�^u��"���Un���n���������U����www~�*���V����l����߿
�����ݿ�4�i�NY�����ukyo�󎺎��,$���$HIE�2ZE��jô�t����q�b�P�x�����AA�T=!�7�y��g��kZi��"h���qj��K	N�fx�s�K��|x>=����������f�E���UM�6�HN&��p~��I���v�U1�<U��Hj�v����E �I�2���Y��~i���ߞ[�[�|��u�v�uw{��s.wu����:\�h�W����%�W���m�8�qV�լB���J�j=��?�y��Y���8q'!	b/���B粳C����i�k�Z�j���=F�U��f�Hh=���WkE~:��ɤ��u�|�Xi�dz:�����(68��m�n'o>��c������6���̸ӎ���[�[�|��u�u�Vɽ�m8�(�������F5���[�}���H'��>}g�<�9ᝏW�4[<#oG\��=�Y��L3�4�Ix��^�{���t��"���}���n�~]]�j���F���]��U�YIyh�M#u�9�uq�N?l���\������TUc>�T%���Nr��UV�wy�G�n�W�-&�[f�jH�>��X��l<]9�Ī4�#�!d�A��V��<`N�O���0�#��=BB�%$!�?���B������A�C��=\�uy����I �zsc���*�wߏ��}���1]�o
H�ӟw��k=3~�{�����s�4�Yt�~��m�+Յ���Ym��[�ͭ庵���㎟��e΀����.���*A!��BJ+�jI$���q��1��}�=]����²����V�{�Õ�Hd#�L�S�]~�IQ^�eo	�%v�*j�x8W]_��X��n�h=�A��<t<ѵ�_�pG��hޕ���>�L�d�Л�4��`¹]>������:lv7�= ���0!��=
��|U3�W�����m�u����-o-o>q�Q�l��T5ޤ�H_�i$����[m���zr�8���qa�����0Ӹ)��)��`i
3=������5�����w�S9f�^���8�����|>M4�q^��BYD0E~7��ٰ��ӆCƏ��לp3R�!~���U�w%����I�8��*�(��q��Z�mo8�����O� ����\CA���d�9�$�O��M=:H�;�I|3���?ň�������6s�"�����W3���C�=��r�G��r�y�%�|�-�y�o�fD[���şH�$���t�RN�J�>4{}>��<(��Ɋ�k8u�t�hxԓ�Aǥ[����l�,2�U*:�.�t�v%5vT� }+J��y_2m�i��Ym�_�m��yo-ۓN��6ˮ"q�1]������>st�o$@M��1{RI$Boﺿ%m.6�m����:O_�����p�zJ���t�t�wk�#�,˳�Q�(�w�g��O�:�R
l�xx�á�E�"t=��Ab�W��5oc��_+�M�㫨~���z��>~-\M^�_����j5ӻϷ�jH��j�?z����[b���\��p�է���ǋ1��e�CnS&�2��u�VA���䪯�Ͷ���'�	)���4��<֘�]o�*���}�a���y<dp��Á�|92�&�$l�ha����k
��h˓ d��/%�jE],vT�i?%�̟��h~3٧j�גb�_�m�\eƖ����y強VӮ#���a�}�McHQvU^ĒI����q����#�o�W�x��]pϿ*�T�>�rt#v���Fݛ!�#���%��HNdt���M�7m�0|Cd55�:�뉵�ʩH�x/b3���6h0d{o�(�(tpvm��ret�J�a�2H���d6!�/̼�ο6��<����u�q�=���1���j������Ȣ0�UD�H���=��Ù��Iz�i��4��$!���M��1�C�D�#�0:��M���Bc�Xh��}������Y`�!u�֯Y����vI���Ą	ѳ�d����8L�B����|��$&����=����P���cW������m&�5���"�������#m2�����6���[�x�SǄt���bx4�i(��I$��0�.b���e��p�IB����t�C˖��!���ٮ6��m��w��O��O�d��0xH�20��.�p�nHT'ǉ[��I���\�}R4]�HIW�����_:m�!��P����4d�Ό�]z�l6����;����dM� �����(��������0�렓�����')�� �� �!�����ZSl���Sh��
DQ�Aϻ�^)JR��)T�)K&JRʥ$�JL�5&L�d���K)I*��"d��)J[$�&R�&L��e,�Y,�d��)�L�JL�U2d�I�%�L�Y$�&I,�K5t�rK$�$�iK*��(�-E2̲�e�M$�JL�%�Il�Id��%I%Ie�d�l�4�Y$�KeI$�rܔ�I$�Ke���I%I&JK-�IRId�I���e&I$ԒI�J�s�[]I&I4�I$�R�d��$�Rd�T��Y$�$�$�),��Y$�RT�Y),��VJJ���������IRIRIRT��J[,��JMIRRY),�RY)*J�J����l���JK%%I���J[*I*J���&I,�����d��Id��-�%�Id�$�RʦY�ɲ�ٓ%&��&L�%Kf�ɤ�I�d���e$�2RI�%�[2i,��I�$Ԓ�d�Y4�M&M%I��%�L�K$�-L�JeL��k�d��RJe�L�d�&�ɤ�٤�i-&��i,�ٓ%$����*�)$ɓ%&�ʥ�Jd�RiK-�Y4�&JRL�l��)��L�[)%5,�L�ʙk���)2̙T��,��Z�Rɔ��U),�YK)�ʥ�L�K,��ifR�,�,����Z�L�D�e,��̖Ye,��K,�Ye��-�ZY��2��e�fU2̦Ye��e�U2�)�%�ʥ��)�ʦR�e,�)eR�K)K,�R�R���U,�%�Ke\V����Ҳ�VV���el����YYjVke\��U��ee��Օ���U+6�Y���YYU ��KU��`0V �����Ҳ�+6��եG����R�L���[\����Y��f�+5��ڕ����Ҳ���m*䤡HE 1P��ml��ef�VZ��U)b���(��X f�e���J�Ԭ�J٪����k++ee�Vm���+6�YmJ�jV�YYk+6�Y���ee���Ԭ�J�l��el�J�jVm�Y����ͭ+-YY��ͭ+*��ZҲ�+-YY�ҳZ���VUR����m��l���+*ҳU��T�֕��VVҳU+-YYU��֚������*%V�6��j�-eYjT�*[eJ��iSk*kJ�YSk*[f�M�EY��J*	JAQQ�*m�M�����e���e������ͬ��Y��V�Ҵ��Yk,֖j�*�+K6��YeT��������\�\��%�Y��.[�-��e���%�,�K,���,�VY,�d�YR�f[JYe�ʖK%�Y,��m*Y,�e��YK)e�Ki,�d�,�J�,�T��ͥ�ʖK*Y,�id�ZʖK*Y,�d���eK*[Id��)f�T�YR�eKi,��,��,�e,�f�T��ʖT��Ye,��Ye�-��[,��YK*Y,�o��eKi,�eK*YR�eK*Y,�m)eK*Y,�e,�eK)e�ҖYe,�eK%�,�e��YfYK2�,�e�,�Ym%�f�Yf�Yd�K,�El��+)Y����̳,��Ye�̳,���e�if��,��e)IZe2���S)JJjS+K))e%,���T���i�K)�,�����M+J��iKJJe4���fVeE%2�))���JeJRV�SJJeIL����^9WR�Қ�ҖSJYM)e4����S)J�S)��%i�2���T�R�V�VYM)�ʚ�e�ҖSJe2��2��R��L�eL�V���e)L�V̬��+b�*YYeYe2��,�f�����T����RRʲ��*YK*YVYR��*el����T�����,�S)eK*�+,�����e��T��V�*ZVYS+fVeL��ٕ�S+,����l�̬ʩ�JS*eYJ̦T�[2�+2������J��L�Jٕ)Y�fT��R��eL�)Y�)Y���2���Ve2�VecWJ��ۙYJ�R�fS)J̨�2�R�2��L�S)J�*-L�)���YT�2��L���)Je2R��l�,���)KR����� '����>�~�~hSM	�����~�(��H
*��!�1�?+�����M��?��_�=����m�s�]Y������'�?�� �ߵ��/�F���i�>�+JNW����F?��,'�5�?��������G�����A�'�[��o�{�*��T �������o��?ʃ���O�G����B(���P?���'�?�0s��?����@������0��a���O�����CO���8��͟�P '�S������H?� T2���bX�6h�1��G��-�������������"�H��ֹ�N��T���:���2��arH����׎�<oT �Yh�ڋ�����(*
4 �,"�� �>*!QUY����9Zf���
��]��)���'���VS���������C�> � 
T��moj��5��S*em��Z��T�m�EI
�/������'� T?w�b��N)��y���� *z�Ԟ�����?A�r
)?���D�� 	����v���с@
O������k���������?����!������k�L�����'���8���!�������A�^�������?�@T �+���Fu���G��+�?q��޻z�Ѡ"��qT �?k�@�~�� _�?���O�)�?���t������)�����.��lF�	���hQ9Z��B��^B?���"�!H��գ��e�C�ҫI)(����S�~��^�EC�i�(�,l���k���.G��	����v�* PA����RC�߯����?o��Ҁ��?�eO�b3��o�����,��?���o�����o��d��v���#����]O�?П������������EO�(�$�����?���ø�* ~g� ��( ��u��~e��1�clQE�h�1��F�(�Q�bب�QF�ch�Qb�bѪ1F�cEŢű�h�F��F����j*�E�F�QlQ�E�F�Q��m�5�F�Q��5���F�Q��j5�F�Q��j5�F�Q��V5�ƣQ��j6�b,j6+��F��������"�*"�-h؋F�4Q�����Qh����(�F�,E(�EDTEF�Q�F�F���QQQ6ţF�4h�Q��lh�4h�cF�4hѢ4Th�4h�Q��m�TTEF�X�F4hээ�lh�ъ�hƋ1����lb�E����1���,Tk**-Db�Ѣэ64Tlh�ƣ6,hьhѣ4h�4hэcF4cF�hѣ1�ѣ(ƍ,b�(��61�F4j4h�F�FƊ4cc�ƣ��F64Q��#Ѣъ���Q����1���m�F�Q��Q��j-�5�Eb�X�m�QQj��5�F�Q�QcF�ƍF�Q���mF���mE�QQQ��[����صZ1EFэ��E�4j4Q�[�E�m��*(Ʊ�m��XѣEEQlTh�*4m�Z*�EF��c�c��(Ōh�(�cb��1�V-�,Q�m����F��ō�b��X�*��EQ��4X�XڍF��j5Q��U5��X���lQ��5F�ƣQ��5�F�QX�j5�Tj5�F�Q��h�j5�FѨ�j5�F�Q���+6-h���X��(��F�4X�c�Ƣ��4QhŊ4cQh�Qb�Q�Fьh�Q�Q"�,h�1c�رb���Ŋ�,h������-Q�1�ѣF64hѣFƍ64h�Q�EF�1F�1bƍ*4h�F�4TQ�FѣF�(�QE�TQ�-�b�Ţ��h���EEE�ѴTTZ(Ѣ�E���Q�Z*-�Z*-F�5��ѱ�b�c[j5�EQ�F���j*�Q�*�F�5��Q��cQ��U�F�Q��V5�F�Q��j5�F�Q�cQ��j5�F�Q��V,Z��V6-h�����-�#E(�EDTF���Q�E��h��E��klF�F�4Q��Z#E�����4lF(�h؊����Ѣ�XѢ�F�4h�ѣF�4h�ѣF�4hѣF�4hѢ�F�m�bƌE�b1b,lh��E�,F-,cX�1EF�4bƌFƌj,lb)8�?���?���� � T3�?�O���'����A�q�f �Z�"�H2��C�s�80A��0Q�bȭ�?!���� �Ki�O����/�_;�;�)��������MP "��+����d�S��7������<������?���^�������5��ِ� �:������O�������@Q�����x�dG���ߡ�~o��(
?�?JJ����O�kSm'�?s��#�������RڕJT�~i����H�
Lc~�