BZh91AY&SY�K��;_�py����������  `����@  =   ��TU*���0����   P(( �@�����&x @ �hx� Q@  
 �E�=� �vi&�ێ3�[i�6���{x���\w��MU+��v(���l�]4wc� >�Ǣ��|  |+�t݀�A�t4�Gv�g�we>�9|w���o��V���e�s���.�˦ ���_ �ӥ:ѷׇ����&�78��ܖ�>7%w�<[�kN�]69rtիf��� ��� =�ӭ�n.]���av�����z��O��ޛ�6���}���k�ڷ�N�a�q�{�=� >�}ͦl��½�������w� ����_F�.5�Z��������]��     P    @P) @S���Ҫ�2b`&&�0`��C=	�EA����A�� & L@�ȩ&)Rh @ 1 dd 0�� �J�0 �  dh �	R��h#MLMM��OSe=���@TI)U"1��L!��0 �d���󒚄d�*���~���J?�� �#�������H��� �D?j���"���B������\:��^�*��2��I$��j���S��e�p��: H�H���[I$�I$��PPD;���O�W��o��m~�l�rh�?��Emߦ�}`��R�{�u`u,]k=�WJ�/ܩG,�k�nF"�E+��D)�~��L^G�H�9i�U�x�J�p[�W1!n�����b�\.��.
Ҩ�&UQ<�Y$��o�pw�-X�:�w�	�t�)w�qb�:�z��HDѶr�/d9le��/�U�J�*�s
�7H�~�\�9gKx+��;�O7�螱���>�9���]�=�A��\b��U�B�*B���u�;��k��=��I��Yp���;�v�8c�E��z�}�a�u�\���7�c�M��GG*ppq	�hj���Cw�;�;��|��R�0X�1v��q5þ38y����>�;@pp��*g��:��;��u��P�9�h�H��W����ZH��p��aư0(�.�FJ�P��5G����o���o�<���A��B��\a��)_��Y�avm�v�]��Ӹ0��5bprpE��;�w��q+��Xl3��;��Wj�7�u+zG��c�_1�����out�;��.f���yͻ�8�oS}��dì
�Z1We�ôY����g�G[�:�y�mʵTi�Z�\�r3���[�7�g>'I¨�&�"���t�F�xG{��,g�Pg7��˫���q�V�n[y�d{ ME��r��#���qү�Vʦ��Y檨聽;y����q�`=<0���WY�gX�7��hv��񜩓��G���p��TTA�>�Uv8�-O��n�����Y�]�:�o��"��J�;�h�;@�
���yV9��X�Vr�u���W2�t`�6 ���4,)Sr=�i�J�/�Y��vU�>�V��L88�!�O���Ŝ΀]���@�	Gh����iyC��ݒ�����s  840(�.��=�w��o���Pr�;[�q��m0�X#�+���Ӹ�|_���0�5f��n����9;58189�����-�N\.��j�2;�\Σ��1v�0޶��{�|��=e�gQ�c��3���m�6����ͼ��'��P���gK}�;�*�TWD��ð]���Ώ���T[���N]�!\�������u����I���]g�J��V�����\��\��QDq)�w�{�{CQ����ʎ)4.�Ah�+\�\�[�����M��Ck�zyW�tk|�J�O���8��Y4�i�q+�Ŋ��|J���������,\��W�.S�(#ቦ?%�k-�|�ڮ�V�x�9b� v�ڡc.кS�ݲ���Pr��*Y*YK���]V�'c]��[��Nt'�R�����.�#�iU]E1xڮ��:Պ񊱴,�U�\�NQ�S�3�/̤�(��.�T��V�/��Y|8S"3�嫃��X�-u[wx�t�>-Gw����d��G���]G)]d��.�]�GX{��,嫰���P�VK��׃��[���.{��KaR:O��5:OX��U��˨��cwj�ŧ������t���Tt:\�t?w�/ῼ�SCt�����Gؙ���b�5u��E�� �+�+�+Q�(���!'ǎZ;��r��J�1b�2�r�@ˈ�v���F��!WV�q4+�E�Z��m��Ʊ#)(S
�D%��g%���rk���k�j��.|ş`��F։��7�b}�|��-]�[�X�\�R�9QҏM����p"���r�ॼ�vHwm:Z����~\�B�Y�x*:��V�\��T�U�.S�(���5,��%!��b��V���q�1�u�5�i]��K�KK�����M�(���>X���o���Cb�j��#�BBV���|����.Sg:\�܉�ӭ���W
W
<���m5�G��r��Np�e�y�:Z�1���i���s*��WVbhZ���-^�"բբ�+�
W

��K9,�#���hOֵs�\Cv�j�k��-LBz6��L]X/-�}�ﺸ����B�B�c=�+uM���|WL�ou�s���Gq���.��G��m
����|*��&$/1:Gg�7Myb^[�3��\\ԅlN��1{����=���ؽHT.����L^Q�B��5�J��P��'h�Z�B�w�W,�T#w�N���ѝ�p���r�&�g��+W�W���X����Y��a<�Sav���.�d�>��GRT�T�WG#��iZw|��wÿ�~`��t��M�o{���o!o-�Y'�!�\pfu�_j%�r�rٴd!D,��U\��OVV�A*�n��¥�K�G��U櫕�#9��w,�����]��n|�Z.�W7[ƏX��B�r�	�9ND�ퟖ�~��<�}������7l������<�8��I���^�7�)H��"{���7�iA��!凼���/�E�=ޥ�/s�=ǠJ�4�Mӌ8�`��F���ld�]x,/3+�"%�sB5�D��[z�_��E������m�d���k\#���I_Ϣ�	�i��c���.�0�T\gu���]o.Cj#E�(���ʕr�\]f��3TM�����&t�j8����I�y�y-eD��>뫁��ߧ�z�z�YA 1�o��y��ݮ�{���sÑ���z�n.�$ �����;b�4�0��eL��ڞ�`�d�2�e�)��K��7�J��e���gL'�u��0�&�+�&�q4��4|=,���Ș`�Ƅ�@�y9\3&�8�2�{aP�"�J���
 �	܍ވ�f�o�"!�O�z �e��+�dfأ�Kuph�.&������$�E���s�U�xn�ei�ؙ����@S~O���8�@��1Qf�C���Y��QW=�rǱ1���i]~��8��ĖE�yq�\�DLQ���C>ȋ4�(��ŖF�FF���q�Qo!�o?~�Q� ͪ�'2>$����:�\�*z�,��}	 I�[PQ�Y aF}I��X��	0dA�Q�-]=V+m��e�gs;=�Edn�)�	���YJl��[9QlN\f�o�(�OL��e���a\�4�� �U�c4���׵�VC��tnP�1@΂rt��#`t�)��I�0"�0ʸ��ͬ��VS��ŷu�$�H$��$�Aߪ7�5WU��fe�m��0K׳���h�R�eZ��;"1�9Ȳv��SS�T��,���gׇZl�&eL�Z� �0��C\�:�J����_Dif�@�ȌS��87:�d<^��^؝x��=���I=�;��zwBɃFQYTF�Q�qf�T@U��mz(ȸ�V�Y�IYqeA�,���ț�d�> �rt��َ���8�0����=�G�~�$�O���=jp����?�4s7ʬڣM=\��2� ��Q��L��Q�!ʆY���;�w5u��~J(�����t����c) ��~��΋c��N�H�㷱�vI��e��=1n��5	��|mn)�O�;����W�+&/"� U��E� A��$��Glon���署���b���ҙ����=�4���ltY����Q�<�8+-T�q��X��Ut����۪�O��X�uSUa��!���\�N�.d���^߷�}�4��� �0�.L	�lP�	ڈ$���U��f
.�Ty���i Zn�"��c匽�4�
���q��� �q��|Q�c���<�k�(Iu;8��0�O
��,��F���	��vʘ�ė8vta F�p�ӀἎ9S�&㌭�(�HR��	�2��<�G�V�tic0� $��8d�Ie��K�\��\DIF�a��,��#J<�E�%Q�Y�`��I�Y=�Ǘ�4�KG��I q�F:;���Y�,�Ȁ�Q�%�u�ʐd���H��h)�Jc�1r�vpN$��)�eQ��`yWDt:$���2��,�f�0��4��=��Ҏ:z4�8Ê�Q���f���[QNt q� �-8(�j���$��H���Eie���'����p���\ @�,fDc� <���(� (�p�4�I�$i�<��4�����UX�$�6�,D� �K8�n�4�0��aG��d�>� q�}�|h��!��d�qC8É0�M6��D���Α�� ��/� �;��2�i%�d~ؖ~�\մ�,�$&����4��4��QM/��8gM�|A
3%��z��Ɲ�_�\�yz w�@�8`=�.���&Q�3Q��ꎪ�1yI&��'�ADN՞JOf��X�c�9��rgJ�g|tc/$ ��e��i
]]��<�
��+0����� �~�Y/��6�Zv�v�톔}��8��?/'��#h��4���>�%��nʧ�8i��J�Y��}�ǘ����f�bҵm�1/�ov,W�װi���%�bb��6/+�����FnB])�dnq`V�q�ڪK�+{��jYk�_�g�����^��{��L�/a&{�[Z��R/r�}j��z1E��)b�	N��̃�X���_��	���(�~���~]6$?S)��?��r~���c��?R�?"�bQ�����q\�o���(~�D
�E索j ����bb�Z�"�Ԩ�Q]��>���r��?tX��X72bb�����2	���J����=S蚀Hv-Ź&����ǂ$�jK$���9S^q�6�b�R��RkEB��?k��_7��BB\�mŋ��q��b�P2*JTUĢ�h��� f�%��ʛ[�)ʞ�X�����ӱ��z$�3�3�`۵0\y�f-D���Ӝj��,�����{\M1�Z����kI���f���.�m�T�[F��,�,��|[��ZSǋ]ш��,W�'��$��lQ,�S�P25�K4�5�QD�ǥ�-�^�+X�s,]�{��L]2ǨLK�g�7lġ�G��3R�`�kZk9��h���Q�x�8K��Y^�~>o�Tg�͟l����o-n�+� �ty�-�_I�W�ͤ���*Q�\p�L���|��L"��=sE�̘��s��BK���c��6���OgK��V+ǭog�&*��X#��/ ��[I����l��E��O��sb^���> �@36��� f3$��Ś���U�_��A���Y��hT����H~?=�����h���O�����������FA}�������_�~^  ��  @ 
 @�� , � � : �  tӂ, 	�p 4@ 
 /������ 0 t32��x`�$4�_|��K�\|�``p 4 �    <1�p 0� 0��� �@ {�t`@ `���{��`� �fe�X ��$�^$��K]p@�` �@ t � �  �P `� `  � � j `� � ���/{�@� 33/� �{�{�vH��NY<�k��9�
 @�` p�h D  �  �@� X k , �  � p 4��=�w�~��< X���� ��|�C�%�|�@ ` 
 @�`  �  � =� � Р � `�`  � ,
���ޯx�`��ú �/���}���M$;� �  �� : �� � @� : �   <��  t)@ t@ h �{��{�� c.��v�8 ���i������*!����UD�	 ���������G� |�p�/�?@������$?p~��_1�/t�n�m���m��m���6i�m�O�÷�۶�v�o6�[m�o^6ҶlٵV�V!
ЅhX��.�]B��j��hCom���;m�o^6�mi�+f͛6�ݴ�v۶�i�+m�fͶ��i��m��ǆ�|�7ӟt�*0���j�=�(�M�h74����l����pv)�u�����U�,j)3bkr�b��뼱���ڻF% �$�1�c������b�7h�]e�3���	(����3�Xh�D��R�3k�]-K�F��Fb�\@�eb՘����OъiC��-ָ&%+�s@v��01k6#V˪�GB����tmmF]�]|���F�#�e�E� ���_�6�j0�83]�%��e��ket���:�L]��e��s2�VD�jMBe��.��9|�GI�ǲ�&��X���bj6Q�������lm<5���Y��gf:8�Wg:��bf��lK]l�uX[?���jݎ���,�Ci�B�ac�utٴ��5$)������f��Ҝ�[c]�6�����a{[��v���,p,cy,z�4����P��K�%�.�Yv�Svs�nZ�ZD��WV�iv�J%��a,�8k�g��ǈP��e	Pź�0��k˘Z��$�
��ݓ������I���V� �������"�f����aduk,�4�%�-ˢ�v#���@<��\Q�ï1�DEk�y0y��%FYlL�v���aй��0���h7k	��L�HA��%s�],�LW��˶�F�cmL�ue#.���w���3f&�CZ�X!�nw2�%/��)�]�̪����7lz]�屡S���iv��k)+��ia�ݡ{(�l6k�˕MK!�JZ6[2�Lk��,j�\b�+y�.��,u.�
����Љ(��Fk��cPf�ٙqvT�֒�fօ{uhlΟ���ާ1[��\He�ݥ�fBVȪpj����R���S��ĵ�M���V�V;j�V��`$���ږ�6��h��RY��-��B�@�jKq�]�J,شF
]f��PҥF�5fI�����f@v��Rh,��b`<A`S̫m��/��L���m.`M6�륺���Ev��̚����-B
��Q4�Q

��uF(�hSYZS��m���ֹ�`R�&m��|�O<ko�h�t�쬙��E�5E	k{j�j83.y2�)I���։�U*�\[Y+A��M*-u�WYY���F`�M���7�p�(����H�����š�@��������Қ����0[J.ֺ�
�]��y���K5�3�l��`ڴ�4:��ml#�v�-�-S�0��š*��b*�H��!�G��D���A��#�=kq,֕��bX��/h�]�e�I���14 f�-�,��-fd�Q�m�- ⥘5d��hשf!y|��c}���yQ��{��1�{�ޒ�
)�I%���9�}�_}�K����7J$�_(��]�fE�����|�rI�w�|}�[���#a�8��G�1C���U�}+p+��3Q���4�K cq��]t�P�*�IIhS�VE��RQ�\�ǭ��X��r^%�h�`a�\)���k�rB���Lv�"2���$3Wr�'1��U����]5����1�IQ�h�hb��4�";�҅��H3R�S0*�����<�h�ŷL豚"B�s�SF��Y����j��L���	��,�̽.#uK��Z�D!չ��ƶ5q��RR�6�����i�΋�S3H���.��Z��f��v�7ȱ׋�-�N�t�y�-�RAU��Ae�R��HӔ� )�(F�o!c%�	�*����Y?�v236���ZB�񬟇��R9v�P�ˇ2{�S�	�6�u���3�a�4�Mrj�E�˦&�DUAKŋ�<�/�T�Z��vm��U_1��.g3.e�@�T�Q0UQ%�a2�qN��&n!����g	��b̛1-��pat�b�8��<�q�d��anM���S&�-�(((�Cf�(���N�-�V,L�4��m�U�I���΀b�n-� y�W�w�J�Xr�V�Q�bC�����N�ħ7]ᡲÙ��6M&\0�u���U˳E<�$����a�*�׭1�{��Z�j秈@�y��y��.w{�$r�Ĕ�ˉ%uh��$jA�8�HB�,���u�R�K��r*C!�ˍt�I#��ْ?����4�);�̶�|��k[G��a�=UB��D�MoQ����v)a�G͆��mH�$�U�f�hc8��gJ�m�İŻK��f�&��cL�[Y��UI%N4�7�@;
)4&Y�ԺԐ��guJ�e�%Q���g2J��i3�IC���OQB^���nIqɝ\KLS���lm�τ݅��eIw�b�w<��<T�u<a�;UWoZc�7[��t��Un�����}�Z����d��K)M�I�v�Ґ��a�`�T���3�EAX`�jD(�RA8T�9��u!,�G��|��ø�H�wN��l0Ǌ����;�ˤ�$�4�z���� �0�,1fdo���^�L��YL�;�q�s�w˕�� +ehU�J�q<F|���
n�︻1|�� N1�0�G���X�wsŶ��r{;�&JSl0Ǆ.-QEQoW��;Q��Y����n{ <ɏ;��GD��!�H F��®��2_�춛�d�v�Úp�#�fz���HOm3����w���R��N����F����9O߹�.o�I��2���i��}����PW^�f�Mo8����5Ӊ��Yo�:�<�B�X�MŃ�`B�;�i�]�1ler��G3g^H�������I�|-��d�nze:m5�@e�lӻ��I ��+vC����w�i5���@k9�[ڋlU�VEnH�U�F�H�j1-�,�y�g\_/%cˈ�>a�8WOi��y�2���IH	ԓљ47t��=�I�:��rf��)#:�e��R���&9j�g$�ĥg���_j�2�����+@��t@�� ��3��쾘2��B�iv@d�o��*������/~mW�3~,�j���[g�������jx���Ǭⸯ������~W���X�Z�+�W�U��x�])�׬����*��U�1���x�YǬ�\_���m�8������M/�����k�_��ҿ/�v����8�r���m~q����gO�ߝ����qzث�*��D��	����7�*���9�58阼/���X�/Oǹo�3���N1Ҹ�1x^-vg
�x�c�x�^�~k�.���e�\U}�՝8ʧ
����z�v�~_	ǅ"��=�ƋU�.U��{��͛,Xѵ�Bq6��S�d�5����-d�ʹ�$g�͋��x�T�g��C���m�α���TU\v�]���֥�z�{��Z��Z�kU�+j�gT���]�OZ７�=kE�����.�O��~��7�>_�f"�������7V܎I2��u�F�ۑ�&]���H�8ڑ�&]���%W8ڑ�&]����Sr9$˻��#u|҉E�Ě��o�qƚi����d��Z�jհ``�0�USh��#& �$�������8��a���i ��g&R	��Z ���E�Ev�����IZSs6�G��4� ��]>H�����r�"EKH\I���q-�|A�L6������E�i@H���d:�&L��,�e�Qdo	�l��,��,�}�<���|/-�U�nc� @����?ԏ�2�@51,Ԅ(x�����p���j���.x�K�7s����]\\�W��O#�l0[�"���$��5"TF�*��_�e�a'rm��d,��JU뒀��[؛�.��NzB��E~bex��������c�Z�R�P"bx�����)K�%#��jGG�ʘ�Ě`���Q��`�(�gI�MIAamɰ���,��2ng�/���˴�_��-���X�*�u9D�Tz�$ @�<�a�,���1o�k�TY]��Ɛ�JU�@���W��Z4�:��ibb�GWC95ᮌXFѣ�Ѧ�&*��6E-��=��I�[n�x���Q�FK�j"�|�w֑���>�  �D�"�pRo ���,F��H&�R0�0ǉM d��G���G�I��^�Vj=ȉ3�1b\S���0�Z��7�qrcfYN�hO��.2���W�?P~j�*T*����a�D���ɠ���,��29��/P�u�9D A�\2�ئ&��1i��rq8НtV��dF}xє������ʗEU�Ɉp�Ɵ.+2BV@��i�Kߊ��zt��x�4>)F+kR5����x��h����%F�L��B�8�ސ�J�X�%'s$���b�-+1Zc�<|�M4ӳ���?+�g*իV�G���Dx�Ob�	�0DÒ?!T�`1����i6se�@q��ކ�ѐ>�f$��)�]�$����|B[�6h�0!�r���*2�v�0P���8_Ğ3[�Yt�~m���'Ŷ���Wj][m4QˮL>��ɷ�`Q�(��h(���,�̆*E�R����>bf ��Lxca� A��i�\%Z�6O�e���o�WWm��)�T-�X�İO��׬�#0�#��&��>u�i�������i��(�'\Sn�$�@�S����r�x�h���-@4�<�8Z��b�%��˴тYYP�{ζ�������M4�N�?+��eߑ{ơ]��ǩ�	�+�� �\9Z{g\wz�9W�b�����R@(��/�73����R�6YV1�Ԇ�٭�Z҉\V0 �4
��z�f��F�]�H������G릋?��.L�K�0Yyr��:sڢ���T�s/\q> ��:�$��v\��×yi���i���;9۹��!��wvJ������p F;L%� o��.�(���R�We2�Z�ƭ��d�m�.$�o����ѓl��g���LV�Ꮫi��iٝ�b�֬LsU��+��
�Ra�/n^i�L�
Nn3X�]$�L��J� G=6ф6ҡG�΄�웪�(��<��8�]i�dhp��<b�Wj�y�P�)m���b��/W���t�Ax�M��e�䌗i t��ӂ��.���On�'?>��kGNՆ��1ٍ�1�i��(z5 �X'��ɚ�<L�D���),�h�{b�2mHӟ���������I!^$ɝ�
�>h�O�[.�h��ˮ��il��Rz�|��۞��ɤ�Lĕ|��VxJ��b��-�)�����y,�2Ra�䢀�P�i*&���b��a�!4�4��)�YTqXi������cN�߼�޳���y��b���s�O�&��&Xۑ��2�pV^ �;�+ݾ�d���.T]�&%�wyi�7�*����p��)��J�Jƥ4y�$2�*���8Iy���2�`Qo���a+���+R����v�@g�7�Ny0މG���'+�*��qx��ū����ǋ��~W�L��?1W���ϙ�_���?+k���׎�1x�xW����*�U_UK��OXǪ�8�^�3���:W���mx�,�x�^-^z�x�x�W�{~g����-��/����������QU��ys�Uu>��"��/D�&'�ی��q�q����x�xΗ���Lc��ی���\zǫ��q�[��x��s��L�i��*�j��+��M8�K����'��e���X,`�|�CG�@�@�f���d��t���;j�/ۯad_��ZP�ﲯ�����2NnK..���\_\KB��]�JB&8Do'9�_�7������c�6m>��ttd�+�h��b{}P�p�vJ����:i�9VT�l\\u;�S�d�H�R�ٕ�on�waB!�G;j����*�B��EQg~�w:Z#Z���Y1^�Vl�����}]4�D☐"��
�"��Ю���N�8���k[E2&J&�5ٺ<zH\z~�-E�
��ę5i�%�t�y��˾�����NI3.�(Ju�s�Mۻ��F�.Mܻ��IRl�̸�)�ڒT�ws2(Jt6Ҋ&�&���R�E��4�Q\^^��
Ȉ:)b�M�\�m��,�	4`�;:�lA[�-�mP-q�i.�t*$ˢ���n�e�*��.��Q1q��1t �յpW]@���Y�4���Z�F���]���ɖ���YN.+���Mf�M&��UMti���hfck���,���]qv�rͧ�`|�h���Z-�05���a���R��;92�f6..��Y����դau��[0̛[.1�]"��nļ�!�i���Qae4�+H�-���λ7n�%�a7z�����c<
ȅ5�nV:��fg[&׬��@�ݰ;)]Xn�I��-�F��e��5������5%�ϓ��m�����xI}�F\gM����\$�q�b[�9K�)����(�z�,L3����u����>��r�'�-b����Go�%֋�C�xek�m����;�I�8٣>bm�I1��K�9�ݫ
�Lc�O�1�iџmr�.]�\&,����ZD}�wN���5��	$�з�(�Rmҕd�|�Fm˨��ɤXtեH�%��Ky
 ��O�����F��̀CFv��������x���N��1�	v�L>=�������]�x�[���Ie�v|`��x��tWj¼i�~4��cN���^c'�g��dB@��{uc��oP�̙(I��[����!�7�-��;@�SE��~��8�0��Y����[n������n�nSuR	U,�TUm���I�zP�6�<�;���yǌ�Di/[�ـ+݅IUU0\�Q��]�ݜy�����2��	ο��$���a���	kه+
�1�OϘ�4������/][��}���$�0`�H�S"��K�\�/8x&<<c?IHY.YLI
L�Pу#Hb�7�W!�7R�Eb�w��mo���e1T6�ڄ����k��:0����ùԪ�Xѥ#Tiӓ��N@鳍)��4�O�a�i�y)��»i�l���ctzdz=>�=�pfQ^5J 01�2�1{>Kj2[G��$�A;x W��3�&c�qpc&/E�b[��T�)vb�w
XkS�!*��4��fw}zH==��i��&O�F���:0���������e�:ϝ�٤��lh�IAzw�$7|��q)�}m0{�V�*�W]�M��j�LɝZ�g�~ʒ��z�A�6�[�d���J�1~Hl4��Z|`�7��M&���"�9߮����ό4�(�+��f���ӣ�u���N��X�8��w�i�S�--N��#��|�3�<�.%�N��WUV]�Ɗ.宀�LB޼p�L�f��q�ph�O]T�U�&��4p�6�X���GS�[�I��+��=A����)���I3]��TK���S�t��M� �30�Çϩh�
`���%��I�%i?X�u� �H�g�ㆠ�:!i���<�Y[���%&Mi��q�dxN��+ٌ�!FNeg��t˴��d����&~��*�5�!�%%Ҋ~�;�:G:Zeu�ZNOX��$%ߎZuKN�b�À���ºi�zi�V�to�9f�0���j�غtf�mV�K�h~��2#o�K,��I��'�]]6څ2�y�"�o���y��^)�$e�Zt����a�M��ͻ-��&T�gJ�ۑ�P�Ř/���0U13������	����p4���F1XV+��O�\iўw����(O���5��q٪���)��¶��� 
fh����t����M�rt\���-%�͗�W֍��*��0����0�ckv��k��,-m�(["��,&#�ĖRf��`ݬ�RҸ�E�ܟa�.b���|����N�D��Kkd��X0�����:�M�vI�5���:e�����)yt��-�(�>�('�ì�mGJ< ԕ�gm�;i<BKSD)4|N�U9J2�aX�~U|ӣ�(w^�t$�I\��*�0��K���3Į~ ��+�����������l�M�&�2��
c)ϡuF�)��`o�&������uI,v"V�@ܔ�(z�$	8�<f�\0�F\��2���5�@u��M���m�U��)/f+�!�	�LG� M�U���z��q{WK�v�i�=g�q�qgo���|\~�j�U_�~Z����?/�U��}d���i^��Vqz^/����g���mx�/��s-�ū¼Z�-^+KŜ^���e�_Y�q�8��^6�/���6�/�{m�W��~m�/����x�q��3o�k�oK���:^.���1x�x_��x���W��x�<��x�8Η��q�c��¸^��1�3��x�Y��mqx�x��Wj��Ut�*�o?%�q���:b�WO���MDU��6%q��VƤ*�>檉�&:YR�=Oom�5�{�I_����l簝����teڹZ��ӎ�m���P)���L��Tf=U����m�����oW�.�k����ȿ	�S��'$���E	N�$�����%:�rN��dRJ��rL��dRJ��NI��̊IU^(��+���Uq�G~[n��������Pm�o��xɐ6��:���Dxm.D�0Ff*��tT.�������mO5��5I#4���׋@��7�T:w��\�wue�%4�N�?0��N� S���-���m�c��8�|���+M
����B⊥���1H��c*���R�A0��=�:�!����C���� �C������f��Ɠ����܄O1H!�_:]}6ӵ!
�O��FL���`y�IZ&*���y�3M3�Oa Y�aX�6���W�:3?oY��g:�)�kp���\����m���z�@�y�X4�'J�x�KR�Ķ�7��M��9MpL�b0♈ݴ�M�k�6�@�H��Yt�qvĥAW,�A�U�T 0tz�� �ɜ�!��Qr����`���Л6�m(�e����U5(�`�������}�� CFe��)�o�9SI�- ʚ���9Ǭu=z���w���e��HY*�Y$���L�^޸S�7�k�[}�X�z�gdö+
�iT!E�Bꊥ}ܲ	��b�<xḅ����8����ك�23�m�f�BT:@�e��/�I�M#ķ��ӄ�>��1˘��.�x.\��NchF^�X�C��e,���mˮo.D�r��L#�̘L��;}=��/Q�ÿ�����
�x�U���:9��ϪOլ�[:��qtL�kR�OzBGf�|���)O�pHwve�Z�U!\6�:Ǿ�$�O��~Ul�9eB|��L�tm!ƇN@0�!�����f��1�1.Z|X�N�ɡJ���u/�p��aX��*��U�}�[�e��}>W2Օ��*@2��8�>��+MBB��*��&�YD�!�~�|���9C�c�W����l�rDf'(*��ӡ�H�����G��쪔]��0JO���o��x��8D��n�SGo�±_����\t~�����[����q����!����Qn��%�x�J�5l���:ծ��+"K�+��z��5��A�5����k(�Lʕ6a�q�f��!�����Z�io��ʉ�,�w;�~�������q5����5��;��8���u�2�a۔>^G�0�]����~}�:bu�~��U%'�4̘!�Z���q�xcN��1�k����ptzҰ�W�ʭ;U~h�����K�]J��.���	��؆'N�ą�`ۛ�Ul��o^=1@|R^���0d�r�ap�,����<BCΎ�`���9�nf;UTU]��$�a��٪�O��$�)�Ex㳤��=��{�~�V�ۤ!E�B�u�;;6ڈ��-_���!� sQd`f%Zg�%�F�l�	$<� e�>�*}SЕ��d��!\^�U��Ƨ����@x
K(���ڎ�bt�L~m߱?5����3��&�8�+�j�1_�<�~���u�k�N��x=`^
��v�MRA��F�'ÇU`AN��:�p q�����4J�*x�餴�䖐��2^�8��D~z�&B���ˮ�������iu���+|Z^�0�����y�m{�LU�j���M�_-�v��[6�~_W���x���N=�ۍ8�7��qgϲ�k�e��qj�m��W������̪�m�e��*��t���U�zW�����8�.����8����q�^e�x�y-�-^*�qzW�ǌ�̾����q�|�m��y~g����3����D*��F��T(�N/*ꊵ������:^.���1�?1��~/���.O���������ȴJ����B>Zc��\/��5��k���g�U��~c�3k*��[Z����/��˺�*T�ul��j!H��"26��eEN]R�w��Q��T���T��[J�R�[soi�&K-�PKp��s>�v��sU���&��MlI��fj2"��̞�"����&�E�-��軵�zבr��rײ-׏SuIl����Ū8'H�����n��P�\D����M_QP��ڨ�f��fD'�9W_�P�E��Z��<�N�ȝQ��U�[,�K�=1���2�vJ� �)�M
���)�=���?��I*��I9&ww2)%Uy�$���܊IU^rI.gww"��~rI.gww"��~rI.fww"��}(�j�j��U
&�M��z���n�B�{�/f5+z�j�4��u�ƶ�YJ�Lci����k�[q���-�9KFl�Z���%�-���ۂhD�!Lh��u�ط%��5�X���F�l�Rl�\U2�^�F�;6:m�����Z���=Ẉ�Rg˱Mh̍���h�ol��L��u��!�]Wl���m�څs`A�d�$f��qP�0[3ړS"� ��M��Y�6�Ķ&ż\�GaсKt����L̗J�O$�J�J*N%�ͪF-
��+k�s�W���k[+���źIs*$Ɩ5�+��c9�aX˥�!Yi	��+*�W�����+�E=��@���N aϜo�TJ���`U��--�����}$�/tJ���p�,�ǻ*�\�h��/��%�wmM_��.�1>z�8&^�lN�h�䑝��iXV+�����|��N}�j|P���k'C�͂dv`���A������9�\���<(���o�N{^�N�	� ����ր�Ԭe޻�.���%��-V�_'�P�}�_*Lhks�P�1����4���9�����$�8mO�N�3���V�U�wVq��qo\`4`���z���4�^���ɼ����۳7I���;��0tӧ���Ne,x֘3ي����I�;���ؘ
�\$P�Y_���jI-��Q��d�O�����B���p��t:��\�ːvjC�}�l�А�L�>4V x����|�1�G���-F[r�;2!���no`lx-��C���x'$���+q���q��n�eb���!�D:��Q���I9�;a��֞��!�$��I&袪���礚cm���`�iLi����,���X�Z�͞�0�*$�W�&��z�?�n���|�u˝"�h��^�]Ü�=��a��\�lf���mi��%���y,m��함˥�al��`�kqJ��Wm4��3D�q3iK@1ʭ���U��l�͜fݳ�Ci���ݻM�F��):q�	��&�@�M����fBg�S��$(0D��BƾJCɯ;I��Jc��v��i�))�|��!�|�����'��T���Mi���~:v����Ѡ���0޷�Q]��C)$l������9H���D��I(tv�&h+�1�%���P��+۰��($�t�6�_,H��fX����ߓ�u>i,�A����X��z��~WO���:a�WS_����ɥ�/Ƽ2�a]�r�K8�M��B���C$�� �\�7�_bk�cY�n�n��n�h*UJ�>��<[�g߱���g5$�UUO��c�`T70��>�W��'��$�����_&@��;��4�1ZUc�ج~a���n��$�dؔ|�Xa!Qu���w��{HN��Ӵc�W�d�zp��M���NjI3��L�l�S��H�x�;��R�
�;O�'����y1�z�SZ�'����������g[��l1���b�z�U4 ߼Qϗ�nj٦�=wS٬��J�ͭq��U�q�Y\��~I!/�YO9�4���"]]�lKD�ZD2����A�a�e�m�$m����Y��m�>b���U|��3��C����#��a0�F�4��|�J3�&Gp�(i���>k2BL'��I�O�>�T�`1w;%�\�U�K�6�GΘ���u���G�������N���i��u=<m�1^!	�V��k����{dٮW~�oRFL����'X�)�L������&N1�&jVʘ�i]@�%m���萃/�/�~1zä�XR�*�(ꨂm�k��W�|UdK-D^��4ܒHB��2���s�'����vg��+��~Z�.�U��ڪ�_��������N/�1��x�q�,�|^�b���eW�W�z��W�U���e_U��������q�/��⸭���j�x�.9���k��j����qg��q�y���̷�\j&'��D��yWVS�J.�quP�8�B��ۉ�*�ʺ��N-��>/E��x�1�U�\Z�/��L�x����=f<�]8Η��q�c���x�xq�\qƪ��q����*�U�v��Y�����qo�߳zknY�PڧwS����SZ�����&n�h������A�E���I.&Q��w\�l�j�}�j�|W[��@tQ��7��������ب�Q���-;E(S�]M9�>b�n2���}�D�q��4E;i�
�#�a��\��=��Tvںȩ���u˾>g\�K���Ȥr�\�K���Ȥr�\�I���ؤr�\�I���ؤr�RI&w�~�����a�WX⫳��W3TL [���UTo�%U,M$�-��2W㉆@$M���p�����P�QP�k	��M'���>pjHdu2��)��lr��i�4�iq�A��Q�X⫳�9����5��[z��9ʄ7�!�&`m���4��(�a��C�*)P���jbi���6����Ve�|ڽY4۾;��ݿ=U���2�:{n~��b�ffc8�<鴇rBRbh�$��u�o%'�N�+��iU�*�8����bYV_�\2j��5��ud[�Yx���2ڈ��I-MP؂=��墰fҬ,�)mb�Y���m(��e�IV��JK�ⅰ4�k�]34v6�5k��e�y8���én�U��(�7���>>Jp`ʝ0=|��O��p`<��@�6y���M�U��e�C�.$�	��}��K�KZ�`WcLVȁ*���W��]�%��:S��GS��c�V6��6@��;!��S#%�D6g9��-'rs�N���d��q"i Y���Β����ű0��]1I�yan&���6F��O>I��0�:&|��
�C��$���HYӴ�T���i'�v��*�򫷊�x��*檳Y���H�w$��d�����a�d,�I��!,m*2�D�������&� ҿ*ד�<���)����s�aRa#A�$5�f�*T�����D���翭�V�����m�񆔭��V:Ux�SO9�s�M_.j���:��f��^��a c9*-U�OSRH�*��q�I�x���d�ߩ86�<�d�5�	y	�&�^��%�>M�O�h�20��qU��\x/盾_zF�^��-�EƖ��L��m�Lh3LbpUI	�>[��$�h$��.V��l���P�UHInne�G`L�P�ulμ�k�D�S3Sl�[l�)-�Z��e��
���m�k�w<��f�p�0oŇ<v:#�ܖd��>�	�^�CE��wXr+I����~M����nw3Կ`�Kq4�o�kNFRB��ecP���nE�"�Iś�8���>�}:SjV��V8�����XL�#�Ln��QLY3��m��Gظ��}苊��
���Z;cӣA)�RL����r�	�,&�wݡ�V9-#�6�@��sK6�}�a��X@"t�Ak��u�5�_|j}��ҕھUc�W�.Bj�]�d�|}a8JC�y�s��c�g#׮w��*��،�w����&�&/ڀ��b�g�U�-���X�G] ђ���2CҤ�V�$���ǋR:!�$��o.x�yf?OO�W�ګU|�o�l�w�&9�b��4�O��'�E�e�m�rƜz��WF��w��l�v���H�J��g�Y��nHp�Ùn�1|�[g�����e��F��#���%�F݆O���N��}��C�Ғ��!�W�]1Ů�6��1W��2���z_V��n1���N+���|�/k�e�x�x�zq��[oz��ϙU��}b��z̿���;g�����8�>c����M����x�8�^*�2�-^-��8��c�ǌ���[Ǭ��qU����z|�]���ܵǬ��p�m�]�k����=q�/e�8Ε���ΗU�U�x�\/��L�x����g�oN1��t�i��*�-^g8���8�i���mU�[Wj���.@���g��K����L�\y��:�%�ȸj������rΟ���9;�8���Sȣk��Uo�G0�^2�n�XveFCw[}��\,d9�Jn܈�{9�������M����>�����F��<�5�]
��۩��N����S�S�!15��O[�Dߞ�=��Yo6����%C*/�l���I����iu������g���ꭍ����ft�\�e;륨/�� ]�ɔ�I��Z���V���8��㩦�j�����+���hֆk��;}�����D�<sa>u��N�y}9UU_�����L����#s\�I���ؤnk�Iww�"���$�]��6)��]��N9�y�)\WX⫏�����1��f�"���L�c2�2���Y�Ф�\�;W�XXf�g�K�@	��x��-{[��r��]����uѱx�Mn3VYf�Ԙѹ�F��X����nV�h����Mn��-l��*b���ah��b�[F���r�+Z:��*ǭ�i�ŭ�eԠ�c]��c���i�f�e��`���Ֆ��&�L�C%�0�a�����������v%�����M\n՚��S�Uc��N�kvQ�RUٚ;j]^��b�]r�v*��\6`Ֆ�̑�Y�������лL��=R�E�K�WG\i�F��t�7��9e.;h��`����4�wD�:
`d�M'D���Κ-/�U�a
�A���u���or�m��c�&	��Ƴ(��n�BT�Pa�:�p�xm�M���!
<B4L����2V1W��qO+�wS�]z���c�[y<�Ɔ�!M�B�0z�P�7EUIR�y���G�p��c�ܒ���S�J����Bm{�ϑ�)���_rw�I��gS�]{j[�0���BޟO���W�ګ*��_l[�PzA��$d����ɧ�N���sV�
�p���&r�����(�:s5[��S	$�ݹ���'M��OBOa�@�Ѳ?��=��b&�ʨ�_�j��"x3y�aDh��	�B��5n�PlR��=@��l8G�M�J=�NU]7eYd��mݘ�]�)��%�)�Ou�c�x��g�>��7�(�B�6h�t��8�=ߣ&}r��vb�b�P�-<�h�4a�R��2t�&L�(�)�c��Y�Ϛk,˦cZ�UL	�E]j�4j̷wl�r��i�� �u���i�05�팚:�:�����u�v�mö�2��\�rV�\�ݪ����<��9����_w�׆#����S̝q)3ͽ%Ԧ�i�.��LJ�d�C	<QN��kh�k�bc��m�f/�����ն����+�=c�1�^�=1:z� �9�>N�;iG��^��UToo���f��&'�컫�Uu�nhө���ȝ�~3�s�^$���V�Щ�e��/�L�S�8����N�<v�J��?(� �����
R_�?Y���)�>c����ٛ��b���܋lI��T��=���pP��ԉ�t�Ry�� ʭF�BIR�QD�T�D�ev�GO'�)���������C{��);�Ӏi�ؐ����GLjo��;1J�N�퉦�\K�K�U��uF��v=�����k0,x�� �NR�x��x��qs=�1��b")[#B|TH��y#KI�f�~��T&x�y����nIQ4u;��ٷ�I�!׍�7\�����Z�7:w(��+�-Mq4�_.'��#��E>P�R_�y�n�lL�m,�	�A@(ǅ[1�ɗɢ/3`g�0��f�P�(:I�kn��,qՔ��8H]6�XͣpA"��b9�UMu��no"X�G$��k�^�Z������K���!�;)��u�$&�����>0�!���iΝ�4�>J��pt�ɤ��?}z��6��\n���g69�l�U8�5D0d�"�.��	`���ԯ����>x�߼�W����װ�&�h�K����Dâ��ьaW�}L[1�Uw��&N#7=?_�S�����L+(Ҡ����M�/�aԏ�I%/CO ���ސ�Q��G%����`�`���|m�q�Ot��y��o6�;lҶlٷJٷ���+�Ǌ�8��n8���o��;m��l٣i�m���v���x��m�m��1Z�!P��/*B�������i��b�mҶl�^<i�o6��ڶ�lٳfͶ�m�.B�-J�Եj��jqdN�I3?7f�1j��I��(]鹘2FA�:"����ErkI癔�������ʌ}pV(��mk��â6�C�]8�N����q.�je��˥r�[y!e�b��${��9�����u8���.��|FMj�&�c�j�ݼ�����_�nc�Iww{"���I%���F�9$�ww�)��]��Ȥnc�I�]uל㜷��%8�qN1�1�<_�%+�MzX�J{���f�Ͻ!=��e�~�Y�*�z���[e�/�N"�Q��ed�cӝ�s�4e?��:�Z���^L�l�U��j��J�U\c���y�)�4���}�K8��Q�OK�ξ4�Td�r ����%�tӋ'5!0`�E&��a��9�;7��\��R��Y�}�8��^'9![��!6��$��iZl�����+J���6��u�Z�o4o]�ͫ�C8fp�2T��ؠ$�ꦇ�����5�l3lvGa��ˍ���ح�31��8�rWvlJ�J�7u���#���-l�є�&N�FF�--�����w�����>I7£l2�,�J�Z#N���%����gv�ɷ͹J�L��S{%��7�ӎߡVd�r�H��mllk�9,X���;�?+��G�U񎇧�WJ��X�3���=����wx�L,:�I-8o6PY��Ԙ��Dre!�8N���̥�ҏ+,��&��.�v�Բ躪}��+�zv��Ό�n�!zi<1�n�I	$%Ӡ~"���ש���?�b�5 =/��<Ӈi��������. 6�y|z�3�ks2�DIi-^�vs�M�����6F�K[m�6�l�$r٧�"Y�!���8on�����Um�}�	��k�ҭ��\�n���W�y6���R�����1�oi�2�u��ω׌�tyKqU��O��_�!�T�	�er�*�Q��?i���O;$�S)��i�tvZ�x���UML�CV~��qU�ƾ��ѻU]��q(����Uv�lco<�ֿ^��kY8ڦ�3IV��ܵԝR"J��d�Vx�`�(5�im��\�ˉ�[�!�	ez��=nel�j��4xRɍ�is�gd�4BP�O���}��Io��[}&��*�aMt���k5U�BC��o�2��!��&̜�ä��(�a��5UG�������J�ߍ'�Rwn�I׿�[]ȝ�j���ʪ�ǌcW�����-�:ԑ��g�D�3�:(�8z�pt�q�oӽ���G6hң���t�шfy�:5l&
B�uUP���8t���0ON|�nq��>��>��+C�V)^����&�k��Z�l���L���
���t�NrW�����%��i�~L��_chi�"�����x�X�-:ƭ&�>����.�HI��$
>NS�j�&�:&��͔�q��|�qU_1��cm���5�u�ޯ�3�������&ߖ��1�MQH�mB��좮��Б�LrC���s�q��9Kk�v�8�~�xlL�>'�>i/�73�*�M5�g��N���8ڸ��m�m��z�m�|��+��8t������x�8�-��8ǭ��o��Ҷ�[0�m�m��v۶�6����!y
��X�b��.�!y�X��;z��n�m�ح�6l�<x��޼m��m6Ѷ+f͛76�m��m��U|x|||��#W����^�"�k���n��Qb"߂���\6�E;&-MVҪlB�{�K}.T�s��y�7�OH���aʓ~��~X���3����n�_%���J���]�9loVY$v��j�f^f^|�N�g�\W����N �[F�IUE2OK�|h}�/�̍���3r���j/������Y��V(K,��3�Mn���柳���VU�m>aE^8�WL@��*��]+G\涮Ȣ�6(��-�j�� �S"�����Y����k)���5g�щ�3s�_�����!�#�9$�ww�)��]��Ȥnc�Iww{"���I%���F�&��]��H�n�k�j&�qU\c�cux��u��[�KYc�Ƙ�Ě�)��m�c6��t4�4�a�h\^@6 G3k��Ck��\UrSsu�8���������1J�^M-X��IfL������6�t�"p$��
�C�5l��;�5�ǘڹ3�4�Qm�i�s�V�I/�))�e*�:�A�we�0Jͦ!Bj[K��np��n��43�4�4����-d�h�fT{X��B;K�e�3t$&nq����6�f&\\Пd���V�ڔ��#
˞����΄P��hB�)[,�dM� �UZۇjV���3K	&#)��4�>8��~&�%��'9�������c<}�LkN�%1�"l$��)+ѥ��BK�M��'S)�ӒC�i�C�a�E즃 MQ�.W����O�{��v>U|�iU]�����y��:̢�U��{��̩�R�!B� ۚ�����@�|�p�`�ᑤ�6�Ϫ��S��N1�����W�x�4��d�%U LM�%�{m����r��1~Ms��<��v��&�y��mɸ��M*�R�����c�8��m��=�F=�r�wu}zh�bbt�N:v}�%�Bea�S�s֦C���Ny`��Lm1���5U	$�d&�ǋ���M����e1���Ho�B�D"����e�w/��vt�W�7=G�OU��c�1�4��W5�6�7�u�<Χ�O�~</Z�o$�� �Ƥ��+mU��៌[L;d���Ym7���g>��03�3Y��C���U��j�ss��*��#�x��F:�q��V��*��=c����n��5k�eV�(�#�������s��w���v���
6�6���3G�!6�"qͻ\���fͬ�2�([����*-p�i��d3*v��ׯHA�.����fe�&�4�吰ٽ�u$�UL8
zy�ޯ�6�᳸%&�p��$�n��^̦Nw��2�o.,L'��]J��0J����Q$��ϓk��}d�/�-<h,!?Q��Є&���}��&"�;lM���ψ��N�2�0�BJ���Rՠ�ן���`v%�jE��릇}��Ct%%�;$��J��ps�4^4��_�ͪ�ct���q�b�[��Z��h�$�,������غn�ؖ&�_�H�-�B���c�BzA�Kh�e��}��Jw�z���UTJ��yOs)@zYrt����Wd�l� 壹�:i
|©2x|���1Ҫ�c�1�e�e����0�2;�ų1�Km�U�qc��`��'����� �&����8b��"r.�m�b�	s՜ܫ�x<;�n�O��$�N�я����?Me�R���ׁ�}u~��`���ʪ����c�UzǬc�_��^3�ݫ�^H���ڭ,��D�,���Sx��k<���.��+kiR�l-�fV���PΎmpf�iN5�s�
+	R����s���.�bm�n�YF*�i{���/�}������vO���_�a3�	nHe��h��;�ɢ���!�Ŗ�%���5/�B�-���b��շ����L0Ǌ����6��;�*��!�p��$�^:�*�xΉ\�A��%a�2�2)����߸J�"��s>�7���-RT|�L�"�*�Ж��{�利���5��HBB�m��|��$>N&Nx4t�Ϗ���i�n��t���m��m���1�f�m�====;x�qӎ:���z㍶��m+g͔ٶ���t�o��޼z�o�c�m:m���m��6��;m��ݫn��M�[6lٵv�맍�z۷��m�lV͛6m�m��m��p��|||�:��oy=׸�_g�G��jZ�"u��p(݇Y�&6��~��W}��{��:�rx�kp�L�z i���i�ù�U\b������T�j���k���0�q�;��{۴�jŕ�UH�����< ���S�k(S�g{�z�z���7K����.}$����e8��$����e8��$����e8�Ϥ�]������]�����J*0�U�8�1��4��<��;Ӵ�!���=��RUQ�{X���eM�"Bm;������s��ܙU��Pi�sL6y;��[;ELw��xa71�i;����y;)�0�j���
(���۳�O&���1Sƾ�B��X�hP��F��w���ͼ|I!9�I2k)i<`���a�����THW�ɧ	��	�>h�lr=t ]g���&����xۑ��0�ʪ鏘�=w��S�;֗^p��5$��D�ǭ�2�	[�)%�,4�ѫ]aH<#s)
ld��.2�
�auG8����,ܤ��wYf���Csv�"��t��+ݰ��2�b,��d��v��1�v]K�^^>m��}�j�;L��x��ٹ�Tda�+ڄ��2��oyB��2ƙ��ğaJQg�M#5�r�5Cdn˺���M&�JK0�9��SAE⪻c�1��w��x��Z�*Y�ٙ=٭�N�d2�Zp��e;�8ި���0e2����Ϳ�=O���'�%��Uj�&��e�}��֞y<e�yM<MRn����ff�����a�:UW�v�QS�U�&!�j&���b�țH�\��K��s71����D
8G?3-v���r��Me$�;�ͥtD'��]���a��	
��w��S�w�ߜ[��a���-Mri��9{��5���PP;P��Y�7n*��S���g6 "��U�n��##P��A�.�=�w;N=�k.�:L�^��y��+�B�9�J�u�)����}��a0 e��ە��ٶc�Um�X�5�W�R6�y��7��j눴Ó���޴�W5\���Sy*q����E���n:ڥ�jȍΚ��S$��`��;.��]).�yl�-�)Hl�+�J�L�ƆMO_`��]Y�2��t��}L�;0<H��g�BA��5G8y	��|���_/~@\S�>Ǌ|�,�+�D�$�\�˪�u�:k{v�=S��a��Z���M>�%ı��y�78����S��"�vrHB`����^��I]�Wisت��*%�F.��X߸PD���ϿFϝN���}�d��p�Zk��5��e�A���0��U|��<~��n�'+8�YE_���=�
��G	�'�M��/�N�y�s�~o<O������4�C�c��ܔ����ć�ܦ���KJ��Y3�Ӽ���~�x�̾6RqO�0�*��=c��]}�<��f��lz�V^n�}��vѹĦ&�O}�o��k�E�4�$#��ș*��˄�y��keǆ6��~;�T�D˳NUUIR f|�si�p���\0��-03��Zc�I[??����$HD��I$�I$"��QG�����?��p��hi����$!�
���ЩD@$29���o	l3�R빋V���Y(��RH�Y!�"�
EI��R�H�X�H����(Ңa"��*JD�,D�(�����(�H��(��R2!E�Qd%H�TIE��Y$Qd�E�Y�kԆ\E�.`Ȣ�T`��(�X��H�,Qb�(�QE��,��1H�E�X��*Qe(��YF��j(���T��b�(��(��*FEQQE���T��,k�(��Z,Qh�E�*(�a�#�(���F�����YE�X;��ұ�j������Qe(��QEJ,QeXeHȢ�,QeJ)E�,��,���X��QEQb�(�E��bQb�(��R�X��RJ�QE�,T�EX��(��T��Qd�Ģ�,Qe(��T��QR��YE�,��)%�X��QR�(�E�X��IR��YE�,��(��TRK(��(��YE�,��X\�F%QeQR�(�X��X��Qe(���,��Qb�)%J,��TQe(��QI*Qe(���Qb�(�EE$�E�,Qb��,QeQe)%J,��,��,T����T�Q,�b����bA�0bA$��,Qb�YE�,��ZB�QR�Z(�бI-�(�E��,P�Z$�YB�%�U)%(�,�h�"�K*%T�����eJ��Rʖ,R�,R�,��R���E,��K�R�,��R��b�JX���)d��Y)R�J%�U,��R�,��JJX��%�X�)b�JT���)b�(�JX���JY)b��K�Q*�)b����JQK�H�KE)b�JX�)b�J%�Y�Y)E,��TR�,Q,��K%,��K%,R��)b�d��Y)b��E,��K�D�R�,��J)T�K%,R�D�K%*)d��X���)d��%�Y)e,��KE��D���R�R���*�)R�d��Y)b�JU,R�))d�X��X���)d���)R�JH�K%,R�K�,R��)b�b�JY)b�)E,R�*�J%�Y)QK%,U��U��U��d�*�Y*�R��d�Z�V*ʱUV*ʲ�T�%T�Ub�4�,U���X�%X�b��UJ�U��QVJ�R�V*��U��H���b�U���EX�%X�J�UV$R-"ĊER*$�TIH��Q%B��,B���D��$dD�RIH�JE�
E�%"�"�Q�#q��*@H�@K)I�D�TE"� $U����E�=��G }��1r��(M�c������QAH�QT!I	�>���'����_5��7���������A���1�g����w��������Ϸ�,��C���)B������$��C��?���2�������sa�����
�? ��O�������UD������������C�b��� �?�I"?�*URY����$~C���������!��1(R���O�����~ç�C�R�@����� ?����*��������儐2����|҇�B��8�/�
�'����II��o��i�k����Ѹ���?a�������b�����\���LE�-qTM4b?�F�?%!1@	@[ـ� �-i��W �t�����lr�/�?����<@# -HB�T	h�ByBL���D�UHH�u���f��?���3�6/_������;���$�L�x?���Ą��?�\��~ԃUQ)?s@n�k�?�C������a����Gd�/�3��&�!�����~�������&C�12?�H�?0����~���?����6����UQ?A�H	�_��5��W�g�?��M�?���/�?�@�?q�*�����b���������U���(t���р��M$�(X��B��e���$!$��6���	o�� � @`XV��6	�rt���J!�Ԧ��t	�89w�?����-���t�Q���q> H�ɿ�*�������j�DUQ?����b)?�?c�
~WB�?���=�������R~��OQ�.�����)?`������zDO�(�������`����L"��~e ���?�0 ���B�EU`��!�g�����������蟑�������t�2Fp��!�#,�hg��7_�����|/�~ <�!�w"Y��M~��ߨdEUI�������F)�
��S�?01��c�;�<��o����Nq"��![сȥ��x����'��s�柬@���S����~��o��:O��ࠠ�~�������K�������?s��)�/�+��X̃QIb9������qw$S�	
��(0