BZh91AY&SY'�c�_�pyc����߰����  a6�U�    ����   �  ��-IU  4�             �      �AR:�A�V6`�8���Z�`b�x>�P��8u�H�����o{��W}��o�����W�wY�n������>�<����ϵ��6ׁ���ت�c�=��}>�*�_]vVmN�ɽ�	}�@�=>��"���o^��f����}�\�`>叀  ި�<z�<�ezꪢ��W��K���w�֯l����;ݮ{���{p0tw|E������{�G[�3�`�zE���}�J>��	���Z�f��r�������}�O�]��,�X]w5��:\"�A�π� �zׂ��[Y�۳ӎj�i�J�.��j��=�Aݻ�������^fۮSgw��;ך���x����Q���5QYn��<�<���շ]���m�JM� {�  ��.=�
�׾��_Z}�r�����������U�wW�W�nK�� ܼ�c
> �� F��]/�׬y�||��2���]M�,F{���t�jS{�����S���  {�4��W���ʯk����os/|��U�k}�Wv9W}�;kw�G���te�� *� 4*�+k�x�����I3k��o]/��}_���_v�f�          B��     @ P� � ��Mꔪ��#``   S�BR�!4h�  �M�����쒔�RA�ɠi��F	�&@ 4	OD�%J�A����`Lb�D�	��4	�M2jz4���h� aOLP�M�T���CL0��4&&&?A�?W럫��#Mb�.b7�?s��~��gO�* P��̀ �Z�����D�������P�UW�aT ���?�詎���?������r�)����F2�I�by$� *:Q����[�.��y�UQ@�#��0�UQ�[j�'�do�B"D����w��a���������������u��?�g��L��U=�8�"�H�ǉ0�R)����d�xi1'���>����&ӸY���6W
��o�D�	��ī��i�Q�9F��ZZs�S]�	4h������ ��p��&͚l�BFɣ�q1�M��d�_&���hm7>�&kRM��E�bl���܉�GY%�ɭ�8Yh��:S¸YdM�W�&�:����O��6Ch��١���uXl��D~��Q�%""sK��U�w	Oe?'jlM]I�R�L��hu8��Y��D��ᣯ�6:ԯ��D���5rW����jR"q;���T�@ܤN�E�*�${)}et����%l�0�D~���R%��%}>�5:%;���舺���\����H��lKy)�V�J7w+��%=��β�h���]����٣O�n�"`ܫ0�����R������舺���\����H��lKy)���N��+���)Oe"s]4`��s�f�>r$e�Ϸ$�L��#��򫌝�*��Z�\��9�:�/S����U�G�8;�[�j�p���nK�jD�	|7؎N�bwl��	�%CO��IDZ����TBT�}�K��E��1�+qds%oFɽ�I��&���ZvD��9&Ʀ�8򫬘�V��ԇ�=�ʕ��t� ��l�Sf�F�ç$MdL5�Uq���2H9�~�Ԯ���~ì��fHfHs�rA�ӽ���e9;���d���s����pNh��<�rAbAbA2��O�'���6�ݩm�+CПD��4OjSܓ��~��jH�����#Կd��p�]wU�2�$�.i�����97M&ɾE{�����*јZ�"aϛ�引�Us"u��}ʪ���UEx)_MOx���{�'�g�[�!|$����SUF��J���P�C�sF��_CTV��5I8�LD\$��Q+�I�8��{�t�e�M�I��&�&�m�s�bAH�a6eaZ*p�����H��Vkӄ�1�;c����~7��A%��	�Nď	�P��'Ru2�bedְ�g���oh��MC]�/��ʒ�7rkE7 ��rq:�LL(s$�0��IgH�D�d�Hu�sbUFJ8��Nh�9�}d��J�h�|_ņ�>�m�d�%vC�\�>փHZ	�qCΆ�f�}\�MZ�4&��19R<�~�IԔ��	��	0G�����Bq�̶J�i�B2E��G�S�?"L�$Y�f}ߓMlN�0�&���8=���$N|�G�S����enJ!6Y���n$D�H��X�aC�4HP�I9ĉ��%�|���H�BtHLI�ͶO����\"&ӗ�"b'I:K:V�"R"8l�Q"'-"#�N�k�	�DGd�"GD�	ؑ47�M��7�0�L'�s�/A�7["'8�
N'&:�>Fa6h�$A+�)I�E}�8��8p��H'RDG�N��0��$6P��$D�d��٢��:$�I��~�7��ݤE:S�Yn�М�,�����H�L1�B�}���F�"D��'���%t�t�ԛ1�,��d��3�5B\H�I�	���&�p�RQ�V	��FC��?\G���D�t���]N����D�U(Ϭ��j#�1��hoUˠnlNlE�J��$D�f�'ɶY�4YUO	�����q��
�CVbe	l��'{'r#��z�I�O�ʟp�QR|��M'p��h�4U�weU�NX�Q_o��'��&��}CuQY\�
�nG!�?1�j�J4���c,��}Ϝ�:�<�8n�S�<{s��ו/�H�֣���t�L��ڝ:VD���D�ћ���QIۑ;MM�/MM�r�_79�!�5>E�L�S�7��Բ�ltH��".�a���jhJ'�"����jQc��.�a3�#*�#ؐM-J0���ULd����#ƧHs������Q�M�ϓ��",M�gլ�ĭj�#��L-jP��K6P�"kwR�g*"6�Å$�#	'��"#�DFN�:�"A�D^�N�7��޵:Ag��N�P��Q�TN����d�4=�DKyR�fTDN�l���&j�7���yQ�u,�����uQ�j&yQ�jl�ϬN��u8#���/MI�F�O�7�TD��(N�DNi��l�D�Pѯ���V�_d���}�D�N��S�&ra�jw	)��d�t�Z_HzM�0��ӿHzOv4���5MJ,��iD�N�+":(����K�v]���b�ݍ==4a���Ttu��2�Q��V	�eJ9�cQ;�:m�H&�U��!��	�54NΧQ4RI�vC�p�i+vYzjX�Ԥ�N�f�ԲTА��;�#���K5�ɣ]��5,F�Q���GYQ9������8��v��\J�������;#2���e2�
[���j�ny��E���ʚ�Tѹ+�K�F��ڟ=�9>X�4�pI;����L��S�������#{��l:�w�c�Ǽ�y3���$����FUK��yʏe;Qr�9Sf�3(戸(�����+u��>:�ږ�'�GRZpd{����v766P��4o����T��{OT�⇸�8&�d2����}���H�ڈ�>�U��R;��c��"�u�$���.;��Q,uڋ#ʘi�5R�#R����;�G�ǃ>D$]4��-�Zh�4X�X�*=���Y1�oR��i���+j;���x��7�G4�����Q���rw�����N��Ħ}2N�*坉H�'Ow�����p]8φ*	9�U���a���>���Xa��*��';$��Md�d��"mep���67r�Gq(��L��9+�~D�5*�G���r�N���m�D�r��p�W#�H��+���DG�+d��ᢟ�%�R�ġ�����H�nR'�"�VrW��e"k���-�L܍JN�W��r�4�R'1��F?L6:쯟�V�~��u)���_@�:��i�H�~���Xlu�_ �"Wu*ķ��-e'4�+���{)�������|�N�+D���rJ)�#q(ے��vʡ�*��Tr�fM�N���a�d��w*�}��N�9��������rXԳR#R�r#���'vʛ�i�`��!��P���'^�VJ%����Jw)-���Kb�WMn"w2Vɮ�I��kS[�n#��r#�NI���8�c�]��T��8%�uNH�d��M�M���7"9:&��W�ԇN2�P�L�Ra����Y��H9%O��9 ��������2v�}�ݛ����/�.	�'!���L���|����^�?T��O�W�}�E�I�
��
��ؔ�!�H{� �	cBĒ�/�D��ǰ�M��}��K��a�)�S��>��7M&Z4�SP�!Xo��_��;�DԮ���f��~
g�B��XW���W�1�����둇�?�}O���g��ĕaЇ����&��l�o���Mfs+��)���҇;u�O6M%a����qz�g���^�K�;���K�����N��ID���W^�m�8��a�T��CXWv��}��pJ���a#���������i�����k�	�>�ińl�t��9!UE��Tg�R���E#��Qh{�JHZ[RSM���n	͎� ���M�m��^y��1jD��~d���4Ï6nYV�w�L{Q�z�4�����=�sī�l\s�.��s��0�y�xp+��J��%��cxa6v=��R�ͷ%��<����:<x�������[0�R�\I�91��.aOu���'/n�\h.�>�Nmt�K���Ǻ{�x���4����i�q�"D���۞�a=�����Y��<D����������!yfy�ܳ.�gf����-FW�QeA{�r��eh(s���W�9-]�B�M��'q�aD�s�U�������N�L,���l�#��Y��Y-5Lsd�:~�8�R�j�n�O�o+s�m��z��6NZUP��(е��0����ix�Pܗ����N�Օ��haes�*��x�x��d(�۴,ϴ$s!dM�=05��Y;1��<���]��l.�����`���{���q�[�.��� �xD�-��p�V���g�<x�#�ݧW���br����3����z{|}˵O�G䞉�٨E���g~���_)�r5����$��~�[c��|��l+��a���1�_]��D������+��v��ӱnh{��Q�9���Vg~���T�8{��҂E���2���&8���� T��,�nn�솕)$�P��:�8q|�4���g
�B�D�]"��gf�Os�y�Oe|Q,nB�|��a��Q�Z�}�1��[3QYq,�a��8���{џa$�QU�>�KO$�J�_�3��+�mp�	$�9������@��BM(��/��ܺ$�M$�I5�PQ��(�$�c�&��_y@ָd�X��kZ`d�ޜ	[��Iy�ni�$}����
��C��?ڊ�k��;�l�5�W|i�,�gp��xFeٳ�;�㓋�R�q��x�2扷�4qا>|T����a��'�g��7�����N�1�ō7+Ĕ`V�|����������v�t�F��fsٚ�,a���t:Iް���NX:k�3��sx#c��GP��s�:���"��v=�TIc��=��ku��X�8�9J�vMjn.ދ��1���^d�Km�/���2�`Tq-����SX
�Xp���J��Ynz7pcq�v��,]o>Nn��6�t}ƛF��Ìqǎ<�OQnQ�*K(�AM�G<�_���Vj���:�&s�m{s.{TYύ�|��R��E\FJp�Z2��ۯZ�=˔B���7=�?`��f��������S�2��D����ڣ�����6fi`�����!ф�G�(��?UQ$�339���O���r+$����Gy'������]��d��6��e�%�7�C�f	hy�N�`ŋS��iK��M3�!QU��dK{�CBx��y�Ӄ�8�y
vR�N��#�64TgWD�0FL�K��DcOI�%=����Er��v3f��)��-a]+���|����r�E��[�nm�e�{>�6V�Y�`�&+��ǃE�M�ՇQoyfS�Y�if��e��û���af�y^]�����Y9��3T���zIqoyN�x�x;�͚��l�+h.�I�������3�|��ys��ޮ�����[�H��SN.�~�^;�o9�W٣0�G�V�ך1�[��T�����!0����o��#�ۏ�K�����!�����0f8�����e;�;�yy{T��繌r���ל�aL@��~ۘ�_d����yw����a���G'��E�[���8s�I�ypF:f~˺����W��?C�.SB��lg1sm�Z�n>t�B���׻_�i�GQO[��Ṷ�A��$.�[S%�{���yȵfP��n����6#ȏ�\a��P6�c��a;��%��a���5$Y�_o�u���z8�w=��Y�*�![���3�*�vnC�l"�9�o37�K�]΍����»��=9s0�zm�}\[��E�r��T����t���,l��8l^���K���S5��6�U_y�'G��z?��2���T�	&N���]���D���a;:�e=~{��1�ǟ"�^�^����]�S�$v��[3�
w��F�2�_2����g�v��;���(gn@a�E`�R�g:�OF�m�eo�K���̌��¥a�W�o�zpl�\d3��y��w}Q����D�i2(ѵ��a0�>Xw�^c�'�~}�{g����3�ᨢIF�Ȥ_v���^^��^�V]~4o{îkEn�����s��B�Y��z۬�F�%���XꫬV<WZm�N���t�fz��s_�S�8���'�҅Zai�b)�1_]3=��{˞�ExȮF��rB}�dщ��f;�I{�%�2�c�ޓ;���1vg��}ԙ����%�c��	�p���=�o	0�3���Kܽ>����,^��BҜ�b+�ھ^�sf�O�)ʕ9O�.�uͷ!�������x$���9�k'�^k9��L1u5�k��F��,�~:^?aS[�5���m!}�⯄Lm���D�Yݺ������rD?~�#�Y?�����r���r1+=�v�$=O7��K�|iq�w��o����!�٫��1��5����*'N�k�
�{���x��֢C�F�8M?��Ǚ�߂�����h�nC=��^�5���h/i����q$|�+�jy����+Ө�m�̺M@�w�^�{7��۩��,���N��^p�̴����5J�g�	:�x�xϼ���z=�R�\+��{���=�i��w)�͕v�����bO�^�ڇ7�[�M��w�sOqU���4'ц�I�W��o7�>�ť7N�!�����c��*�%7�,��d�Et�f�i�5�����ϣjs'
0�J�}�t������8�9�v��Ε����;�n2;�#Պ���_w��V98�(�my$[i�t��v#���ϦFI. ���ՓB=�\x�zf���y껙
3'�΃�TϵB���Vw<���:�ENa�2�zw[�}�qEqG�L�9:T��vx��Ϝ�\h���!��.�_�D�}�oR��N��ß{�3�[�r>�T��y�����2�Ԝ-��uٯ�d��?,�+�t�p���ez�=��'mo|{#*�do�1d��G.q�RmP�ٙ#g�h�2sʹY�:�V|������o�@�%ٟ���ó}��$������[��U6�1f��g"�~{W=&��wmY��eu�\��zgӧ��u��\�J;q�6�G��rW\Z���M�̙�����Zߧ�dgן�%�������.��m�>0��}�Wz������>�^�N"u�)nO9=YxO�.^n=P:����b��rn�n'���9��5 �nkeHp���#�tGi������e;z����~�����=�j���m������N�0Љ$�\����oo�e��b��QQ�';pk(b?˻���$/�����2K��+u��?#��2�-Å�+g1�ҤF��s�]Ƴ&7��w*kW���k3���#��1)���ESp�.ID��ƽ�|��R?��8O�~�a82���� ��	��?�O��_���g�f��םk��@��6��t��2�"���A���-f5[i?d$�d/0cIkn�&A�-�ֶ�\�M�f����L�jպ�٬�+T�hD0d��m����fWE�Mt�.��](n���i�RX:3X�%�-���F��D.:�#��7�*p9|Cl��FE<�d�-:�xe�tw>RD�i�6D�f�P1b4�AD@J���"�h����Ķ#oc����坩/1��/-�
�7�L�2�}Ҷ����)�gT�����lX6ߎ�u�쐖���[�Ͷh��EZl%��ݱT_�O�����~pr�Y�s,ˈ�34�l��k�D�	�[k�#����;��r�#��)5,��,���
�/�M�(r8�&2�D����+����ț>�d��{4 �$��W�^$q��Í]�Л�:�E&rTK]��	R��AJ#�o�wVFRN2Jne �3����&�ΨŐ���]�D��f��ᅂmpA�6	�P�j/����7Dj������}|>5��6��"L閲I¢���#O��݋�:㮮�ͶR�LiVoW�8 5le�A�~�~=�a�YV���>�����vf�Τ�a�v�����M3|K���V���ͨ7�١3eRm]��|���Q��76wa���.�͎��L-f`�6ޮ"�te�D�[3k�cf�	]�E�e�SBWH�w+�dV�1����8���Fi���-���yf� Œe��V�"�7�4�3W8�D����m�d5}��\ :�K��*~������%2y�yܭ �eO��U�zC�$��&�"H'��p�R�<E8�_MtR�b�B�n}ŴWɅ��E����L$�e2�ڦ�?����>����d�M�e!̴~?�+r��Y#l1� zEc�3� ���x�}��:�nV�Y�9��DZ����H�NZ�֥W"���߮�u��Q=v�n&�a����j�����Tp�H1#���6�@�
�D�����}��B�����/���L�H������q�m�皈$!9$�%�Q�'�ff	�Y`���4c�9.���F]m���ݛ���[P�0���d�c���
	cT�*����CH,s��4!���VQ���T���B�}~�O�;-i8B*�t�(�� $�/�OL�e�
vHb�#�SV͔�-�	�Pإ
��#�YrX��P�j�?�H��fAm_
3�҉$�1�0NT�AQ6�մp?3q�ap�bC����6��ͬ��u9�H�4��d �����@iXE���ϵ�o&Z^�w�Ӂ�P�Bv�ws���i��-�o|��g�;�ٮﰟ����C�5�H��Y@ O���}	����"��џ�U$�D?�sI���<?��O�^�$~����~����g��9�%z���ҫ����[Uv��U⴪�QUU�*��*��t��U��U\X��]"���UW��WJ��]*�*���U\X�����եU�Ҫ�WJ���V�U�+UJ����UU�UUTUUTU]|����I! �@���}$[��V"j���jHB
��P�.A�E$��kVQQ�U��Y��	>����qU�UUq���ZUW��U^+ZUm�X��������եUڭ����ZUW�Ҫ�EUVcW8��Wj��ګ�]*�t��X�����եUW��1��[Uv�uT���W����UҪ�ZUW�Ү����I��!���-��[D���M%B�@R�hb �,���%��	l�i"Ő-����) H+!p**H)������z��Uz������1UU�*��t��U��n�]�J��Uz���U�Uڭ��Ux�*��UUq���Zx����Uv�j��[UҪ�ZUW�������Wj��=���Uv�j��]*��t�ګ����;a�DU\*
�b�T��*�V"Զ"Ԓ����UZ:�,E���c�{�����yڭ����ZUW�Ҫ�X������Wj���ҫj��*�W����U^�*��t�ګ�iU^�UU�UUq���1U�z��Wj��ګ�V�]�J��Uz���k]ZUUq���1UU�*��iUt��I�}_O��>ql2��E�qq�� �3T[$nú��BԚ��j�SVj�-H���uIت��u�Y�BU��d���˗v�`�� �D"f����T� H)R���5��������UE  Đ�A���������� ~ '����(�G�?i��2d��M�>,�CgH""'Dě �"P��:"`�����8YBЂ �	�,M�8'N��a�â&	�`�F"&Μd�K�	E��6"&��,�M��%�6%��"C�"l؈��8P�$܈�҄�(L�ن�,��	�(J��2|�!�>D��JbAgN�:p��l��B"lD艂&	�bl��!A8p��:X��]�?�d{�7�Y�N�u�b��j?��s���sspjˁ�[��a}lu؛D��mդ�MqXd䅢�.��K�����n�����.�v.#��щ��:�������9ң����L�~U����3������7�15H6k��&��YZ���M6�k��ـh�˦�F՚��4Y��0��;E���i[M�����W�-���bY�1�TH����t����l�5&�ٲf���·`ҩ�U�Pۆ	�d��D�ؓh�w����M#�o׷o�m~���N�h����bh��cCH7�M[�u�vש����u����V�,���LJ�D�]c�b,`���F}=溺�� g�f�+L�Y��W#Cc�����;M4�)�]_&m��pƆv��
����Kl�Ѝ���`���L��R����޸��_Ǚ�V�/�S���p�@S�(��5#R��LJ�Ϗa������si���0��S�J�>��e�q����#^�S�wZg���ݥՃ��\�{�	��ٲ5P�Xl.������b�|�.�厔�Yv���f�n�Ѵ`�ͥ.Ժ��R��֊V�0��q��QUU�*�wv������UU�*�wv����>X���U\b�wwo�>��*��EUW�������1��:c�;cz�}jY�Q�0�8h����/�%5sR����j�0=�ݓ��7l��ř��3�z�wM�k���&n@�E\�B٩JMX�ӴX�<��źx�@(z����%����WRڭ���>|�ۺCN���oMuොUZ	���q����K[KY.AE-K-j�A�����CN��p��(��J���
-�x�Lr�m�Z����^#6l�����d��o[L;�U+a�9Fp�A���L&����Y�(��y�S܇���������h6�ȕ��l�LdE|���cq�s�L���*}�~���_������������Lt����\q�ĳ��a�:p����֢jKִ^vI$����r��|�����:����h뗩�e<��*�J(�I�4۵���	�K��[%Pe�H;M����:m�\Tѭt��(�%���Y��][�^6��N�Kč�a���CH�rA�g�w�����jD��T�P�g��G�95R�*� ����K:�5xӮ���Wlt���"pDL������C�|;5نڵ���%F�6x%���d�o��$��y���G�x&LC�ߔD!'^�=�n9ㇸM)ã���bN�U5�QvY%�%����ЄTI��n}����m��6#��eNo1���BK�%J�Rp贳&Pw8Q�Er�M�5L�c�H��y�9�w���Ld��R��&�p�Nu$�9��+%�a!��6h�f��CG�h���%)�2L��R$��d���I2d۠֍��<M����������I,�D�����Z�v$"G^^��B�i���N$x@>8|�pHAޫR��.������Dg���i����r�����2��;��z2�EY1)s07.a8d�nD�z�jJ��}��Y�E	�J�x�^:n;=v��:x��8��L������G2j*o[��C�OQ�1"
9�Z����52�	�aF%a8M�|�*P�9SU�'$ȧ�q�<��L";T�݂����$^,��?b�5G��n�]�̺�o;�Xhu�N��܌������X$E $4���:Fb!
��UU-�ۛ��5��;`�&��e[J[�s����w�����t��4Ww��ĉM*p����$�ts��vSQT�!�.M�يL8�]�優���_�?':�!n0a�)Y{�T�LbK�x�������̸f�a��Y9�Y��7�ciի��]�LC)Ӎ�O�>Ha�U�.�됝v��:qӎ�|Ǯ8��`�����Fӛ��Au���@�5R]}UT��ON�y����Õ�UUu�cnNc�H|��
�]ɢd���J�&��Eˣe
a:�8��1��]�$�2�������,�ݜ�_h�3l��gJٮ�d�x�
i���4|�����(�Wiz��<��T�s��\R��pOJvqEU\�TL=��s����;W��>t�ۏ�z��0ND�t�%eW*��s��Ri:�_;UT���=�����Ue����E�ݜ�h��h���q�_Ã�x4����OK��l4�tf;�mB�]�j���#&\���:�.(xy���M<�' �!�w����fA�)�S��TD؎f�9��S��\�x�x�L%l��s�	
6Y[rIAl�����	�Řa�"`�&�Ç4`c�s��l{ uW�2#*���t��U<�oy��s��9�y_FWͱ�����_ln}f��������%����ѧ�[_�	�5�G�3�ϳ�
O�>%�o��U���}{�ݵ6��O-չaCo
�,��S�@��'����6LL��9�m���:KeT�C�-�pQ�vw�l�R�)l�	�BhK<pDL�tL0�Fn�	s���adE��F��ccɬ���(�$Z�govQ0��;�SMN�]����ż��eSsDjC2�~�v��}��f-}���R���)0�m:�Ż�ە�7g\Ii7�����U&I�9�n��ؔ%6��$��fL�L4�A���}����A��9iU�������bn�l��TC6Y�@��:;�D�
nS<GP�[jʢ��ɴ�y$�ɖ��1���z�I�;1U]r�f��0�i�y�:�[Vl��&��WZ.��wM��W+$��4�p�:���]����2i4,�Lp�,��"`�'�a�:p��=
�úK��<��Ρ��ܭDs�y�t`����*�8�!M��.��������ɝ�\����ќC�UE�����F�	�M�	,�4��a��@�e&
pGU��|a�j|��yS\e�-
��7I����p�F���%�a��n�9A;$t���ʁû�Zm�Vw��n�̔�7��J�q�;������v_���4����],�+4�����vN��xzB��b�'�'Ë���b��z֮5W5���\<W���O!�xJ<eI����v'����)�*9�Q���(����🄃؟�G?B��~Wk�go�?+ܷF.��4�ư�$4%��(�x�O	G�%���:ƚ�x�.��֗���5�Z�b���q���\\i�\^���mb��z�+k-�������cmL_�xƼY��b�鶸����u�����o]t�\\\t�L\z�..8�/k�4��k5�q���1�O�4�ƻ\^���?F�~�G��UH8�dS�>?�!�j��옞+�	�XL�*"k��x�*���k5��ƽcX�3V⸸��O�"�|N���~"}O�E�̖��ۖ��f�����R���y/����'?^W���N�@�wK��~���\Gn�CŰ�,=[�R�㾞&9��>���K��6l�	^��_o��2*1k�ϯn��}��)����fTO8����S�İ\�A����N*��;y���`�IOlk�����7�ݔ���;fo:K�[���9���T����O���k���ߟUU�*�Z��>��&fg3=�ǽ�*�*�Z����������ǽ�{ʨ��kO���̬��������{�QWZ֟}���h��<x���&	ä<xDO;��]ҝ�$���]�(z�S�ih�eI�T5��	)v�8Ah�m��`� �@��w|�q��ޒ�� H�LK�E�m�}u�ّ���Q��Jc�'�xQ{�->z�0�]�3��1�u*)�XUV�Dc�2fZ�MGd7rIW��[���YgfN����y7�]���1�2��!�A� y!��@�\�Ulٶ#���>�Q���Q����g�i#�BR���Dz괎��nV����p�a"�'C׭ S����;�1qd$�t�>ҬS�0�s�ԫ���06Y4pЖ'�0æ0N�O�pcA�ã±�Y��ͫ+��C�����*�(�i"�Ĵ�
:B4�L�Xu�6I	$���EL�:B�/���H����F!	p��m�]v:id�X.EE�D����rR��@�I(~D��!�p{�����&�0�v�礒��d.ZN`%�I�BB���4E��&��:��a�%�__2�He4�< z�$��/F�[;y.*諤�i `�j�e'��Ӥ[��Z�p��3ګC@3ʎE2��[SR>Y6�>Tm�s�>{mu����eX�)������BY���D�0N���#���j ��!h�}�dD�=0�ç��[)Cq]̅v-�e��)��_��BH�̈b�)�^ر��l՗��4�_����q��L8id��?Hc�3<q�ͷ[��~m�8��knu���S;j��>��HhY#�ŝ��#�-+q���i��!$$�� ��-�6i�#u�YZ�aCm&ˍɃ��`;�{�ZK��ŴR1"�@�V�!%�h��Ejr��"�+���?t���r��	D0��V�Ze)LSC�	�!�����d��$B��RH��L8ñ�R@��g"�)�,N��,r�åf���!H�F)�wmJ��&K,G'�]�,�u����雍���8CdF:x�L�%���]仳rH:����bݔ�p���5'Q���iM&�e:��8�o?2M�Â\�!�Q4���F"x���&	Ӡ�xJ0�ؒ�;e�\�[f�t,�9	!$$��*B4�hv��l�0�#���~pȟ{�dd�e>�8y�Z�57�����>*U:ޓ�\1H�2�܄!0q S ���ȁ�V��ۢ�J^ʭA��#o&��|:��z��>��="��)0R� ��f0OH@�C�rm<wK~�o\�^o*]�l�#ռ;2�p\&
�dX�3�����WR,z�M�e����nH�rzJ��x�J�:f�l�f)�d��O����#��X��%��> �b%U����a��p��F~6h�h������0DN���xvS�s��e��RÜ���!$$�����a��R�n�����}���ֺ5)���ŏ��ŇJv�jJ'�dX|���)�̔�ͱ; a"�ؔ��ThL$,��3�G0�j#���0�� w�l�w%)M����tY�
A%�h[t%ڮ��dpU�U��i�ăK4C)`�K��i>��+ՉӚ;�m����mN��.��M˕u�ޕ���i �4] w����l��/˓�+�$ F)�"� c�>A�X�!�q Sԥ���_Q0i�H��E2G	�d�tԝY����֍,?�c�W���8�??=q�8㍶qÇ�6Y��s$�R���B���6r�������F�]���0F��;B��^�����$$�� �$ ��CR��Hʱ�Ɠ,
!����E��;$$�1�YJ��x�D��1AɇBL6�jub&(�l�����%��p3�&y��!�� h���',�Nx�_�;{KKΥCD*�廆Wc �I���HQ�C�/�b�4S���fAþ�ym��u6jL�a�)�.؎�1 Q$ΒӰ/�m,�Cd6	�-.�H��'�QS2��'i
b�p�D�`ۂ���Q�Sit:�&B`�C�=�*�>Hg�IP�@ʚ�HҚHh�
Y���$���᧪��OΟ��8���|DN�a�:aY�u��I�\��z��G��k�U��Wf3��������CrE�����%a�Q,H�:����3���m�V��X��ڬ55ڵ2���A�m5�\Ռ�ֱ�kJ��f.ۧ�@ 2���mH��,"�_ѫ40kԉWv�4����J�d%9�䃲pܨz`~4�	�u��d��w>��t�ڏ��S�����S+o!f��U2ry�����Ut��+�=�jSز�Q]�r��w,7+�*:�2��t[�$D��RwKZR�y�,�ʆ�0&�"��!.IO`~=N�5�4�)�:�⦲{Ԟ���1aܖMt����O��	�q�0F�#	J��@�x�;w%]$���ӏ23�EK0��)vT��FB�!�@�\���f����8u��N~{��n��dV�f����燡0��4N�4a��?���"t��pѧ�~�4�j*��gԉPv5;8i�=�BHI(���X����U�ѵ��~�8�k�w�����[� 9�:��gY����gt�
 }qۚ0f'�ѡ�)��������4Dkx�N'Si�QM�	e�%���'�w����L=2C��H���j�n��ᔎ�b �u��V<F�K~�v�SV��K#�����Fzs���n�7>��@ش�@��� i_�e�\`�%�i7�ʒ�>�m"p��#��Io}�L	� A���H����i5��D�Æ|S��`�d�,�тl�~8"&�ӢC<Q�Osi�k5�L��t'!Nh$�H$�������M�8�IM�O���I�ɂ�%���0��ny�&�HH%��i��@�L&0��X����8t��16ZB�&O'����e�r짗mE��¡X:�W4��IT�$%�Oǳ��L'�M4��rPt��dN�'O��/�`���r�6��'����7YX�ӳ�qO�}g��{��)�n�Ӳ�8Dk?�vIvV��J6�>p�|p��R��L�F�GI9�w��	���37�l�"��L�f��(!&Pe�%�{N�Iy��Y�ǎՎ:z��Ǐ��\q��ӢC!��N�kZ֦���>��<�M��UO���ρTj7dB(Y�}�0�.��)儐�@�~�p�Nu�:t#��O:1��ϒR�ь��t�Ii�Ёnө�������p�a}U�X&�L�����Z���S��M:x�>�Us�V�p�����J�)�i�jbf�W���\�aƉ0��ͦ�y��a��X)rjH�Z`�Cm=H�0�p�KE0D�S)nz�0�yia�&�R⎖�0�O[2B�d
):�Z��WM��ȵm�֥�Fr5}*��~�z�E<Qgzb�<��;0��I��B�D�E=!d6G�4����8|C�h�<!���ω��G�|?/��������|)�>��[�b�Ʊq�[������OW�����-Wed���Z�+���s� ���>4���,�#��!��d<Cg�8F1�Y�M1Ƙ�Lq�/��c�X�����������Nߚ��q~t�X���\\V/kK��i��zcU�<cX�_X�-��cL]庘�kk�Zz��]��iⴿ-cX���c���c汦��Z\..1���.=k���v�0�xJ8O	]"t��p�(�x�O���>):����"?���UH'̋>���I�	�4C�J���sS
�*t��5�Y<��UcX��\k�5��j�^.+i����z��Ū²[r[}\Z���XV-W��g�(*���~H��\������hG]y����ِ�� �9*{�ff��b\-�5���q��pO��?��*�-�w��͞�0���������wu�	�4%]t�XD��`�G����W�sZ�k���c�ۂ��I���O��t���u��s��&J6��Ս��ㄚk]�\>X,��vh.�F����Z�yAI"vȍ�̈%�'P�nd�a�	m���i	N�8W�y'��W�^$��
vT���XA�r`@�!�G,�)���[!cP���%���	q��wa�&PE/��'��Q��#њ�<"�$��o��	��e�������<�j;�2��0��	�s�LB�6-���v1�,�X��J���X�t05?7�܍�H���W�1<��ȏ�&�هşn����ʏƦ
Aޛj�yj�����7��t�2\BH�O]���\Γ=�da��]͏�yuQ���3ۆ�*}��x��`t�	JF�[E�!F��5]s8�ǨD�n�Y�E����<D%ݓ�%�	��o��k{������I2�>��	fM75�@\,�`��4�ˈ�8�k��C�w�9)��2���}ۜ(Ԣa��*�P\�ٷ��᯵|d��5�҅�l�Z}�O8�0��Ւnٹ��tW��e!������,�r;���K�5 �M6\��.��m������؛2m M�筽К��4 ��n
b�f�\�q��s�j�k���9��m�)���5%��L�3l2����i
��8�P��b]H�>.�O� �F��.��e*;�d�nl$��(�H1-�D�"-��K�?���X?3�FU�y#^]�}MSUpj����O���{�V{����y�kO������{����y��yֵ���Y���ub��{Ϗ{�ֵ�{�33Y���*�9��fg]u�n#�����Ο>x�=D��!���k�_���q�fC2hۦ=�����{�0a)ػSJb�f�Z�қ"Ɔ��Im��ƚ[OXK[r��n��^�Ea?6e�a-�ϗMں�m��t�kk6�|h�m-�Td&�V�뮃�����]�^��BI��E�ml����;�7zzԺRJl���37Rl��O�2@� �JB<̓i���SQ����^�!�I(3����p|�9���F
\- h���IR�*T�%10�t�
u����ɧ]&��,��-�9��d���Zh���O�|J2��ۭ��e)���� x��pӄ�n�%J�UXL�ku�c�O6�&����:����\D:����ģ��6�
���dd��e-56<M��M��9�۩ɻ��ב�OF���ȓa�3\����,i��f��=)�4x��6'�"`��:$0�;>;>���>>�Ѭ]ﮢ��1�b@��M�`x�EP�=@�t���P�"��_F�����%<"|v�Ҕ�$1	_[����jp�H�������>4x�n�!@y����0@=����WG����J�P��~����p ��!Āi�Cm��-�� �ݙ�b�l����QSn�<SQa�nԧlt�,�����M���,��7��u�����x�I�I
 CDh]�:\$�Lm�[�S��Hץ������ۜ��CV�s9�.�5��cr�Ui�c�����1����"'N�0�O,�O�J��w5Ϲ��FI�,NL�f�;��e��c�!�ܘ���pӨz��)3��a*�K�D�%<L:0�H�����a���ԧ�9����L���:���s��ILa���&㔮�Q ������*B�Ŗ|�Zٸ�NNsd�۵6�v�0�G�xs<8�P�O#&�jz��u4>����C�*&��@(�$t���u5�騻��>�F�ӥ6�W���FB߈�<{�A��8i闧��ݴ��i/t�4e��+N�c��V6�z��t�Xۦ:x�?<"`��:$0�<t�<|��"�H뷦�}c�1�B#��:��%Q
�J���O��Cd<�0��M8n�j�1'�l���	��.q=qC�|/��dH:V.�6s���I �g'A�M����+�,Ɋ]6S�B��0ǊL>J4GL�<Za�Hh��#�e/�à�/�dJv.̌"6������a��Ķ�s���a�C�
SJ}��4|��,}�o��֚tۿU*�T�w�o-��7	,��҈d�A���$��8n�<�5����\)�hpEn	�$��QIT䰺M��&!N
XQ��4x��6x�p���"t�������-I-=w��Il���ZWݵ5�1<�b���nk��|[/5&&���	����d0Y[�x�Zޑ�û�W�&eP[�,,�Zd�HsK�Kp�J_%.�w����F�c\)%C�o�S���1�B�~8~���-mO�[��e:6l�\��:�S��Z��~>>Ë�ڷ�O%�'�E1p�*`!ၚi*$��=N�WvU\�0�c� ��C'�M����7�/R:Qҝ�tu>56���Q8��N�qUV��&#�~9֋�9�r(�[��rHG̡��Dl%��it�٦фn;䒏2oD�f�t�{���������\�!�ɹ�W	�0����|8����=EHN܃`�s�r��J۷!��PE�n|i�2�F�]�<����'G�e#Dv���n;��#m*��2*����ԟ*|~i�O_�>t�ǎ?=aD��!��������ꦒ��d�Lc�!���c���`�0RC�&�9�����`���3KʔM�S��!k�08@���-$u�,ۄKC��n�IdK��3�����a=��!g�$$8 ��rRՔQԤ�-��� F%ĢH'��ū^�@Ԗ�kDx���c����������>7�h��3VfF��v�a8r;l��ɞa���I��kR{�ԝ)���`�^W˾?~��&������(��Rff�FX������RS�Zq�7Z�Hry$���e#��e�p�gx�����&�ӢC!�pwغ+L����1�)I�(�1 wa��T��N/�	�r�h����B��e-!�p�C��2;0��Y,C))0C^�K��a�>
~��= ox���^����2c��W�P��	��x���E�,�~y��A��3x{��HZp)�$xC�������k������\'9$����t�K#~4��<��Ws�;��x�h@��4�u�fL����}�N�-�>��Y��t�,�����0֙#�0�H'���M�2�>S��L�wI��U�#����Řh���㇄L�D�C�����̷n�fD�m�7:޷�uz;t�c� ���;�Ƀ���U�.��s3����~�K�K̆�s��H��O�B��YP�m�S�)-uIT���l;�Ӈ뇠!�f�)H��0@����"�D��i�S� Q�A��������댔�a�'��DE1�EB�����#L�Q�@:b�Z.$����NI4[��H|@��30S��:u�s��d�8��X��L`ݝ-);�w�Ur[E\?�,hܞlǱ��MFA	7E�6�.&J�n�q�ڴ�Y�t�?�0��6~?<xL�D���vxw���gYi�J�2i��ٛ	�@,�GmR4vޭg����~ӻ�7��f7��/����^b��H��8-��v��,"���i�D���[�F�e4%MnK6�d��3kE��ߣ��1�As�I�$�j2m����j�W>�]+�ig�'[s̒`����->!�=)��Zk�,2@�|E���eD�R4t#�c��d�d!Mۆio�y$��[�4�(�Ln����>S���p��2BSyh0@���{�>�>�����sXe~`t��BC�US��J�:��#��&�%�=�)�~��\�U��<d�d�,�����)���������ZQj�3�l�T����xgۉ�����p"u7�L)>�&]�}4�4�??N㺘t�v�o��c��㇏	�"t��tu5d�E^�w���Y}�n_KjMZ4��Ι�Bt��,�'h��-J�*T
 T=�rM�Q�ִ[` e�A�G�UJ+N�IG��m�y7�I!!����I�d�����'ƞ �~�ި0>��N�TvS�Ѥ�1p@�|m,�d/s�F�T4�>u���R� t~J4i�p�a�HY��h�; {O�_�1��Ѵ�7R���������Lf���LP�x�2�gB�.=O���1Hl��<h���!]�3U�U��W��p�KB�`i=I�x0��C$OeZv����OFY���q4@�T�h��^�0s�	��4}�������c��p~,~>���~���z��֗��f�Lu����bxjz�I�xJ=�+�+�6MǈV��ar�U�VaX�qj�V,��{V;jv��xҮ+�]LV.Ջ��_�q��N4���������	^"C�O���Bx�<[��]�O�������X����V6֗�5��;cLz׌k-��W�4��Ʀ+jc箍�x�&����F��C�x�,�~'ˋ�[�c\Z��.�/Lk��x���p��	]'��xvL��8CO��|4O���HE���>X#���"?/DU �,+LY��i{\Y�ұv���\��ºN�W���f��6U+Ǫh���8x��S�"O�W��p��	���/��>�Q>O��_�}'�Q?
%'�G��տA�|?h�ȶ�"Or��/|'A؝�Ռ�y`\�,�k����D2���_�B>(�ލg�|�7.��Ʉ�c�B��NԷ�����#w�����z���a�;���ܫ�U�%�Z�3n�{��O�&{��P���y�\D�O�|xp�����{~⴪�S����k^��ff�3=�+J����޵�������{�Ҫ�X��w~ٙ�����եUz�_n����00�Y��Y�<x���`��:$0�5p��WЩ�.T�c�;�s�d�ʢ�\�<SWs�,joV��ۯ�8�l�|��f_�a�NBaѧW����3,8���0��m'q�G�m~v�&C<��~zl����&��XIt[]�;����2���rJNe�Y0!i�L[a������!d0�h������1RH��b���EG�2�p���|�*����'#R>SqU]K9�>ه}8����9n��:���ٺ?�I����t�I�,!��1jCf�l���,����<&�ӣ���F��Y����QES�w��pN�?!׿�u!��l��W�)��K�0x�/�!EOD��.�!lE��QC�桿�%�v����m��F�`�%#����TnX\`��]�I,�L�6k��&8@�[8���KJ=~��]]���m�H���	��A�D�n'f����s	דǝ�1�a��]�(�2a;��'[H9!��ȟ�i�%�$:%�����JH��<�G�Xz "i�fo�_2Ќ6h����H� B�$"q1D��Z����RD�$^�������)�Hyh�I�QM$tk��獫ՉN�+�o�v���㇏	�"t��toy�Ϲ��>�,,�朽����z:���4�*;�zAcY�Sq@�i��b��
�21&�f}VQjrQ\������F�ze��̫R�b?�FYZ�I&V��ee�L�8�hd՚��4���Ha-�܎���\&m�,�M�v��ff�4ŋ��)��z��	!$�	uN������s*\͵�V �/ޟ$�괺���V,l�O�d��iTv@�\f2P;#�4U!i��;!�N��E�ɓ�7�q�)JJ��I��AD<���U$�*�
"���CLC�"p�I5�pY�	����o�0�0D����$h���"p�Y
=��+ G��`8��ֲ��A�̶�z�bu���.i)���#�a"V���A9�y2�-���fլ�.͖M��"Jp�8~ØL�'Q�\8!��d*�5THH��Q�����D?~~U�BLG��L�0���n*xv�]�t��=~~m�c�=;;=��;9Ы�a~����L4��M�+��=S��Ά�Hd�>qP�޺��b��:�'�M��G�M�&ԫ&�u�w)�i���)����4B$O���i��hci$<�B�(��5*T��]6s�^�!
(!&�`�YAI�����N4��|Q�nJ�b�Yvb���v&�d��@��iL�����j8��Ӥ�_�!�>�>�+Vx|��<��=������>h�ō����bگ�%|M��y��	LH44C���ba�?<x�"t��4M ���g�� W"��[�_3���6h���p�BI�����7?)d8�)��d��b��a�HX�a���d7Ny�EcS�[���l����C>>��q��뱔s��t�l�>�x�����&�E��/�qX�q��FI$�S��E�J/��e<��ayq��94'2��䪨�CI�x�C�-8`lrY�=�T�!��)�MS�Ed��ӝ��nf��d�������wv�[����i�|���bo
b>�<{I�Z�N��r�"���Ǌ��ӎ��?=q��1��㍶�|���;����3���{��_{�$���a1>>Rh���6CA`ѣ�;4��L����ߵ��ÁI������+	�mn�;�GK$K�#��å��:�e��I���[m��HH�!�ѓ�p�4Cc���`�7���%��Ĳ���	�%-��I�#����pZu����O%��`��<�C��Evi����N�i"e9hQar�	��>�UZy7�ơUbƣ��r;�nGQ�SN�I:���ڱ�Ξ1Ç���ǏxD��!��w2��j���A�2P���_a��#Ac@ܷ�R߻�rkf�|{w���y�Wn̬�Ӊ�mЫ-ă&$A1(M�םBp�m�hX��̕pl��پ�l�R�#�ܿ�� �zΟ3��`݌$cb��M6i��n�D��a�:;��w����Pl��y�Φ*�9*��vQ��N����I�7_Ii�����p�w�5
h�%(��<tL��p�=��{uQ#�!$���CD�@�4��2}���E����p�~L``��ѸnI�oQ�~[�w=W�W�v<�Os� s4���M�|].�*�]�k�ш��B`�&n@BĒ.Ch�Nd��_0Ӭ'æ�^i�rx�(�Ǐ����##�r+��oc�x|�֟��O���?6�1�q��Wϕ��<��Z���m'(NE�(����V�m��k���BHI0�~s��SI�ނ����=)�Dd*�!nR��W��-��Ub���:W��jq]���'7�*Hx˒Hm�v���mi6�6�(!&׉��t������ESg���h�<ZG�GEV���?E��8Y��Jۅ���4��ܔ�-�2���\RB	a�� �	���=s��6�OjL�N������!�y7�e�M�4ٷ��8������A!�����E�9I�!�4x�Ɵ�:|��z�c��=;;=��;!*Ԉ���l$�����O�
a0�1F8p��h�����D�f����T$��.��{�Ɇ��d�Id���RSE��!��r�
cӰJSD%`���ɧ�y������߷��ۻ%��f�n�14��T<�J���
ɲ��al�(ڴ�T���GX~ܘ+?4�Ө������*�Û���P-���q-8gL��!��O&�������%Q	��؛K��rv+���Y�Z����8i'kEԛ�+�9xZ`�������;~t��1����|�m���N�O: N�=�\��䭅S�!m�y3\
[n�-�k��������L ��n�w��#,���EJeJ�ĉ�
!�'�&4F��q=�Ze)����TfHJK��l㳮�l�l�u8��!%8!��l�_zKt�re��q�M��	���Zl�'~�u*�N���:=vt��<|����OcSi��2KKi�AM�h��4��h�ق��\�.;�w��~��!=��iZ���j�u:���:n?Jb!�:<��YYI��̇�<��w�(�i�=�Gg���d>'^*�}�����`��GD��~&p~��?E4|)>��?��u�����j�Ӷ5W����Ʊ�X��6έ�q�1��4�ۯmƽY���V�d��j���
'�|'�I�.���3~�	�~+�Ř�\Y�5>cS�b�}\q�/Li����~c_+�jq�xJ�
�6O
�Ⰶ�J�8p�.../����cM~~i��_����������M~W��58������;cO����|\^է�mkc��cX������x��.�5����ǭ�Ř�X��k��m�m�v'G�z��ӄ4��?��⟍!��L��"?�W��*���4�Ú|H<��h��ا�wY�{���G�i��~!��+���<O+�K<Rx�ǪO	Ft���i�^�
°�[mb�aY-�1�Vҿ-_��knk���<Ck#?N�B���n�۹v(}��c:s����(E$
H&_�Bu�m��P�\B����2d��J��8̮&$�4��\-8�4����w*K��x��#�)�����Ƨ۬gzK���akF�
U%6�b�HIH��$e�7rc�T��r6�[!7��GI��\�Vs��2�P��pU�)k�x����֮�O)Da@^�P@����=���|Zi��$��1s��G��m\9.�y�nw~��ĉv���v��I��ۅ��-K\h�����ڬ%��=�2z���z�MT8\B!���G��N��2R��v��u��P���}��t�V$�2y�<�
㨩���+疻0%
9�0%a�����빻�)#���%[�q��<BѸA� ��S&������ �(Y(i�v��p�7(�툔[�1�qƱҤ�kE��{t�����TGy��!ɻ��ky�5I���L m��t�ǒ�ʽW
��i�(�3IO��I8J.�D&��m,����q�,L��hTl���c��W��٭R��st1� K�3Gi�[4\�����[�k[eh\�z۩n�Ԧ��.�ױo\׌�o�{��)믬��׀��]�4�$.`L�l@��o�u������"��+�H�z��wxwI�����b��2�\k�%��sk:�)�ۍCJC�"&�)��T$���GN!��k�a���|m����i���7W
�����_\���*�Պ����fe�g��]*�+~��Y�������t��V����^fff�=�UҪ�Z[���a��0�pÇ�<x�:t:t�p�8QR}r��j�-��K��HF�5(+p�fns��SZX�D�����)b�l.�4����+�'fZzֻz\1�7l�fn�q|x��F�3��M���m6��Nw��BI����[�!���6�s�����5�d��"͂mj��u��4���ýT���'Y��}�<E9�>έt���vn�4��p���v�`�0�Ã	�PY�̕)��׋[v�59�;x�^~�1�ji4i��wup��AD"Zi�Ӆ�"fT���C��)�y�S��d:�Sq�:V��v�Z�^ås��Ĳt��d�9�B��)��i%�������m8i�d���(��ȝ{��zQ�˺�}����,�g]�tǯ�\clcc�6ٶ���������73 ��˧e_�A$B���th�0[�>��h��pY�K�pz�<���U�cN�ƴ�D�S�"o�`[�~a�	�C�'�UT:��}�J��j}�th�F��4Rt�Q�=�G���f%�*��*�v�ʠ�LbH���	É�)�~��T��!��x2p���d�۳ǒ��2���~�}r1k����l��:���ucG��|�7c�F���O�������q�8�f�W���ۭC�a��+;r9�6�7y�w��΀�:G��t_���BI�	�?y�c�Ϫ��lpBz�H�8t�яL4?*���q�B=����&��6B�f�QgL�a:�!�N󣬁�E�$�k}Sv��asms�m�,O��ҍ1��(���QT�h�'�O�H�&>;9-M���~��L�Cd�q����F�'
��7	a�<8g�G���;Q��;G0�y�C�N�2~G0H!㦟��m�o_=q��1�1�l�؝�U䵷�$Y�rBHI�|��f說�*[���$�8j>)�d���$����L�������B{�Ύ�lѥwq7m+�,)��i�M!��a�ü��'���_��!y3��+�O�8~K�UU$Mu|�pY���:���'D�㆓����d�(�u��WWip�|l ���$�>�;�DO�)�@��&�
Lh"rnS�:Û�}>���d�*�;Nd���C�m��X�C��ת���o]�����c�q�Ͷ�]M�y5��Y�Z;�M�;��(�$ٍ�-�X��s�~������5�.�:�ŗ�w�!iYW��jBcSje�w����-�1+�X�����P��+���Ս��UUv�uۦ��fl��{	!$$�A8uθ� ��`웰da>4q���fLu	a�1-5�=7�Z�j�_GSlX��$��]�2h�l�aD�,�UU�]=>�Y��}�)�W�'�3�q�uV�ᐄ(�l�פ�`!6RkfH(���1�)ףD2�}�#=�h�s A?^D��ݵ�%��V�4�%���%���� �d<�������[-��U�UwKS�U]�ROb��4�i�f�xp�t����㍶m�zԎ�ձ�u��>����L �����}�8u��D�|a�*��?8t'���!���rޥi7�ދ*�N�[(6CG�&/$>M�a���G����'�H�6!OK��e�R�k�4��X좆�M%�m�Z�͛B� �,�4���:Ù��e2F�tٽ:N�.���Hu2n4m_�Z�I���~z��tz��w�<t��N��⼎<e��O[V;q��<|��6�1�8�m�m^�����1�3�B��TA$_K�`���$�8��ܔZo��B��L'�g��B�'J,�T�]5r�
O��(���`���>h�ϒ�<�
'f�>�b��Yl��g�:Hk�l�M��6IR��J�*��ᤢ�'R���H[�l�)F��&�	��Xd��&d��1�NJ
!��jMD<	h���i4l�`�&���sk�i�IAD4�Ae��h��g��aA�d>0d��8��m�c�c��m�z�T�"j�lT�>IЩ�%�Lc?n �
�����gɸI4�M���ϳ|:b2y�G��?pG���t5�8L�C��]�������k���յ$��\���ؕ�Tq=�<)��1X!�e��I!�I����{�mGm�Ǝ��Ӟ�ֵ�Y�����,ti_�i��ۭx��t�;����U���Q��8L!��$�^��R9�YP��Ha����>������g˔��C��۷��v����ߛc�����A��D�"cp��(�Z%��6��T�m�Ka�z�nB������70�T*�^�)�64�{$���ǖ�3�(r�0#,��ce�gm}ܩ��pa�bx��e��6���k�!��BHI0�p:yq�¸A+�B��3c"�UW{Hm��'��%vO';C��7��X������pNa�y�r��!�ɱ����p���eJ�柞���gWQD�<2�I�ʹ�I*<�t�Q:�Q���}W74��}o���[���?~�k��=z99���j��Q�zOѹ;4O'�W��5-����k�a7ib�$fg	���T^�;�1��
z��a���Ti����)��%�U���tӷo����������������N�t(<�Yܙ�I-��K��>ץ��6l|V��ͰM�Y&�fs��$���a��&�W��p e6OJ�2i<��a6�!J�eq"S �Ri4x�iA���������)=dJ�Q����bQq����a6y6�L�He*�/S���htB�k;1xŖ\5S[u��M��p6��b������K����p�Yߘta��B����}���P��)õ<�=��yh�coє�=S�v#i������Y0���rC⌛4~4~,�Y��G�DD4""tD�H"%��pD��p؛,�� ��Ed�bhK	��tN��0L,�0K�0D�0�Å�"Y�,M	Ĉ�4 �M	blD�N�&	�6%�bY��	�B�DD艆�>FH�܈����x���p����%�f�ДP��"B	��A���J��<t�ӧx��G��b"pD�8"&6lM�(AA: �x����g�������*ǻI����v��g^=�Zi��a|=_�z�OL��f�r��\N��]��D}�����p���	%/uȩB��7�2}ȗ[asv0{����<7q}NG�W:��b�Q�`�f�M�k>G�N��B���^����N2����>\��
}�Q.7�?�yj�z�u���Ѿ���{?�G�����0W�4�q�r�^�뿲���j�U^+Kw�k333y����Ux�-߮������{֪ګ�in�w�fffo3޵V�]�������aF;|��Ϙ��6�1�1��m[h����S�	!$$�AC���u���'M�+���r:w=�+����>ɽ�r�&
�� ���� Q���L����.��>�����`�Z� F��c�����f\�>�{a��0���Th�f�C.�&�䆝XCƋ<�&:��"p��(�bRe�M]:O�C�)d5���I1�QSL�Y��n��Lq�;q�Ͷ��Ǆ�Ӥ:Q�W7RH5ʗ*�]�z���!$$��'��2�(�(��8��7rl��N��u"c�9���v&�a�h��߿2�vC[.�c��������B�m�֭�b�����p�Ög	�g�hv�}������!�$��'�4�F�h�Ip2C>�n��N&�h4B2h�LI9!�{��)�ZJ~Ҽ�j:k���jt�u=*��|s��1��ֽ]����Wm=|���n8��~m�c�c��ڶ��_����^i){Vr��/��nQA"�o[�pW�mS�Xll����+Tĭ1�ƛ̓�'۾];abU���t%��5���d�R�5M�:�8�[7�~Жm~�7U-�L�.�&r[��B�6�8����+�j'�����O�$
!�$�;�Y�c����hҼy���ܷ��l~N��u����UR���Sү^q�"�]CSϖ��ն���u���R���1v�8�y�V�;��UU��S����S<�L�'M��y%WJ)��l�rq,�S�Gښ̟\,���� 	uFvR[F�	�[�UtUs��|�7�񇑠чIק�$�2a��I��e�Cf�l���:v��oͱ�q�q��V�z�j�N��rBHI0��\s�����o������|ƟVU���^���t�z<8���F�֥W$��Rq(S3�&�� ��n
@�u�t�ޕ\Ne#g������`���FȐ!��/+�ꭉQv�sSvl��+�n�5I��)i7O��?|�ᾟ=>&�������y�O[d�e�I&G�6@��G��i��+C���~Y"�p��ό7�i��	���x��������8�8�m�m=}��R8G2�C\#�����)a�ܒ�/�a$$��M|�a�uU�x�!IF��CZ"{x�i/���9֧�S�U)��2{	k�)�6D�E�1�4{����wb��Tn�\�lr@���Q[4�C���,6s���&��d��&!	$ڦ��<j�ۄ�i<��o�'�Ag���$)��E;:���8{����OѾ�:�w1f�4X<��KHRS�ʱΞ����i�<z�������8�8�m�m=d>��ՙ�t֨�����H[�O��p6g�n��7
�=���xe�8=�l������Q�"���d���V��!�tY�OqRO<��r&�2���M���	'	6��5��� 8$K5�)��O��R���=bm/ne6b�%�L�EU89��l��|���GC��n��	�)����L6>��Y;)5����j�O�<|���ͽclccm���`+|�F�M2�&"��5��ܵ�AT�J*�[j4����"\��I&�WE�^�,&s�y8�oyÖo"(�4W�;sm�بgim��*š��e9�K��Y�m�,r�>u#IM$�%�l�z��BI�'NǫnA"JŎKJt������Dk�2EM��������1�;Y��ƃF[L��4��U�UQY��C�m0Z[x���2cg=e+�Hv*?���Nλ�d��0��y/;�
�E=�RU++i����i�z�s��NuԌ��pܧ�*.�H&���5�:�Ha��SRu9��ƻd���V�k����UU>O�$�I�ϼVIA�4�x�7�|M������d��e6�(����O��1���lccm�bvC����Qp����5�s���7w3����?y�$���a
`�:�L�h9\���(�８�b����88p�8����ݦͮFx�~:y#���K,��CF7���<�e������tm��KN��#����!����EϜ5'����^<��E���dl���.+��䒖�໦�y/'8sw]H�Ę��a�~�u8�<��:�d̒'d����*���S�~O*�Qߑ�}�'�{\��<9.T�R�wL�p�|�;�`>>!�Lz���㍿6���m��	/we����T���	�rT����$���a!U<ɇg��<����CD�8�l�k�DxD㗊��wuWU��~S��p�3F���8�~N�p��bJ�FT�-�h�J=^Y��y��FM^L�q���X�>~�r_�ZcJ�۩֍̶����V���}瓇��_y.Ǭ�=N�78l�`��r$���Y�|�by�������vOی��jtgD�>m���ߘ�ߛm�c�c��ڶC���0^�]GXc�"I0�L��+V;b��e�0Y\U݋�i�'�rBHI0��O���X��l%K2d����y<'2�'�So��(t�C���~|'�*EKD��U�R��,��d��
{�g���
e8�ѣ��PC���(�$�8��PQ�W���Oٰ���↜�?aЧ�I��wT�8_�W�g���$��BXR�D�̚0`ф��=��V������ v(|��8�����U]4��O�?;���Yg�AB""`�(D�"X��0M����l�E � �"%tKBX�F�N	�0N��D�Lf	B`�""a�:l��X�"tD�H"hD�3	���%�bY�4%4"&�艆��$8&�K8"`��ӧ��6Y���<Q�x���p�a(,!B&�6$��8l��b&	�!�ǋ<xN�'D��M��E � �	��v��G^����ej	y	0��4t��5����*���Խ=��*��]/�+M9��n5��b��aX/9t���1C-�$�p�gɈ�h�ѩ*ߋ����D%��M�K��oЋ�(�<i�L1�b�����+/P�̃� ���͒kA&��f-˟m�t�C�+b��w
@�N�X�H�-4$q��dɉ��'\�o�ģ��F�����
���5�����ՙғhL��F�a��lubn�ꪍ}�P�\u+ ��B[m��L:3�Iܨ�T^60����:~Y�ؔ���[���5(�Ć�<~�f����4��X2|׊�L�6�'�6�Q���|�fE��pM�1���������)nX���I{}���ך�o��A��1b��ct��I1CB�1��&!�3�F��Ce��\�K��=~"Ąn����f`��ӭ�s���O04D���E����o�ƣĤo�,.�MW`6l��e�=kw���νڇW�µ5��w��az)��{�1Һh�u��]f��g4�Z��]`��^�
�-�J�#�GI#c%8Ȑ�����Y�3(�֫K�ƴM�ЗDyA-4��:	���LՄ��{{b��^��dާ�غ��q����������H&�a�k�#P�1	
!�͵�GK�d�Si!,AN�H@.wg����p��Wo8�<�J���U�w~�Vfffs=�*���WM���Y�������ګ�]7w��fffg3�Ҫ�V�t�߯5>W�>|���o�1�6�������N�ts���n��f��[5�Ve�"C���=������˽��j��Mmi�P��f���� Mn�53�͠mX JQ6�6�P�h�6�\��;�f��[f �m\�#�M7���s[&��	!$$��}�a*dM��2m�V�������I�@~<9r��8m�D��p�wE6L'�_���fL�I'|d��0l����cl�a>�GS>3>���ທEcgS���;��T�q��p[Pd�6�#����J2�p�9�!|g���}���w1tǛ��^����S��$8i>L���htp�}�Ŏؕk]ң���#���ǮF6�������꼫�>���S�ڿ �C㲜?zx'O�N�<xO�N��G��ʭZ{��I~�hI{���A$_�-6oӡ�a���d�RD��I��cgϑ�mZ���Eu�k�#��I3�1����a�ϓF�'L:(!p��yэ��1�����)��(���BtS�Np�h8��ز��Rʛ%b���L�,��f+r��94�N��}��-��n��Km'��r�8�=a��|�a�!:�O���`�P�ۂ>�zIÁ���2&�8��I&B �l�bY�'O�Ox�<'�І	� b�om4RȆ�!��)��BHI	&�x)�{��2I$(�4x�h�Ԏ=�LQ<�zt��Li�`�g�![;��#����������9�E7:y�_xH_���e���/v16ŭ������e�v���vM�������N�˞+�t<Å���[}3R�*H5�����n����nϧ�����ǖ�ٳcf�5"Sw��2VN�8n�%_Nt��G��mW'S���ƞ������ߛc�1�1ǭ�����:��kΚ�,��Oe���L!Ç�׬�y�qu�W�SE(�6u�M�h0}�LY�l���*3���I	R�{�;��<j1�l�r�}�%J���h����z)��vzp��<v���5܇N|r�Lzʹx��\�:�}��fO��-��a$�$�Lo��
:�)-,Np����5WY���w�$�!���M:��������_����G)ӵ|�n:m��?6�������ڶ�׼�ެ��
���"%,��Q1R�QfZ�ZH��qm�j��l�i�a�jÔ�&�6/������n�p\,9V[1�In@�`���iӋĎVn�sve�,�fM�L���%��h��h平��bh�6�i�?���	 ��"���;�c�im����T����+	2K1����~?+���>xG!�˳�:�$���Y�����\�.�m�!������S�jBI	(��<��#�	̥�$���Q���Q�����0h������Ǿ$8O����]s��l�%<΍:�d�4�F�FW*F�H��m��Y���O>آ��~��{�9H���UUt0XM�����o��Z�>xV����:m���c�>ccz�j�OZ�����iݒ�^�u���q�P��@ @�|򦒂���?>���ɿ�eI ��Ъ���3���}���??
��������<�<)�����eUH*�0�4S&B6���!�>(x_�����-���n�6��T	1����p����4m0��W.p��~����kIܵ����>>��<�E�2n�i*I8�0\�UU�)���C�r~ُU�O[t���0����Ǆ�Ӥ:Q�O����f�6�r�����L!����4�y2q�Q�q����%�|�h��=8Qk$L�SC��N�Ç0�ҜCi�6�a4�>�Y���,1��h���&�p��d��I��IR�Id�r�.*�?�.W���>��L���@��FY�rB�j��6��:)��L�G�������g0�y�6���I���/
v&�gH�G=~����i�=z��6�>|�8�8��ն����κ�eg�l-�KJ��6��~�� �@=	Hz ����˙(�|gag��*'Ɵۓ>�pp���>���.�	�Ո��1�Y!ad��|s=>�H|Rr�h��@��m�e]�޹8n����f��UL�t���$v�RxCЅ�y̇������ї��[���nGY-Z�����Gǎg3U�?g�}�m�vik����;:��=OM1���[V��6�^��>z��m���1�1�6��m������*	�KTOYI�
��"��.���6�{Q:f6�-e�u>�;$�xN���<t�n>�C��wF1���.B�bk��̰1��RٚmQYn0R�@#f��b�kmQ��i|b2�]t�sn��vlv�ƷS����N�>�]�n���3M���f�!eq)��w��T����q��>��׋K����S�L��Fy������K)o����i�y�,�\;��ã�D��ecd��Տ��ɸ�-�o��d�v��	����Y�o���Cf���O&C�<J�`|`�NB��c1��;<E��������c��-|�)�.�QRY�K�UG������?|�o�UR�<���~��I��4�]4��=cm�|�������W�:l쪵M�v6k�C��*#�����-n���	}��I	!$���p�fC&����S��֯��Sa�G��8h�1��v]��'DH�-1� �Yf�2e�}�n����G֚t5��V�d>ѓd0?~�����r�f��vIix(�*-UHV}�8�p�g_�$�ہ4j&���9��	�=�[ɓ{	���ݗW,�G-����tr��Ce	�G�?,K,���D�0N� �M��:pL:a�8h٢�A��6i�4&�M�bpN��a�	�`�&�:$N���D鲄H"	b"A:"tЂ$0M�"'DJ0M&���%�f�4A�"X�����	B"X�$8"`���g=q�n;u�zq�1�cJɖ�	�h(!B&��BP�:l�Â&	҄ ����<t��<"`�pѱ6h�A<���?z/��HY��9�`����!������2�����C7KO��ıZ���%11���W>.�ò�&^�i㞝��CnM=���|1t�l���;6���4���ܭ'��;����S34x�]
�Z�M"G�y{�˾��J3ۖd�Y�o�t��C�8j	Sq�=��3������Ì�o��sU^*lQr��+9/y�=9MQ�LƧ����r��/2�9�ś��/�H��u�pd�f�?a�����р��y�c���e���V��݉�����g�{J��[U�wz��fffg}�U]�ګww~������J��[Un��ޙ������Uv�j�����0�S�Ο:z��c6�8�8��ղ��HI	&d��s��tt{�D�TB���'I���l��%�p~7Q���/l8�h7^����H�@}T�X`[�駾�[tQ��}�O�ӃŘsEHT��^=���=>�8w*���q�oƿf�&*H`<��<���ᇢ�,�
oy�I$�L�:<=�Ԫr���2d8p���:c��>q��>m�q�q�͂4!�`���g�]��R�b�s���BHI0��î�t犩�b\&�$6S��ii�+��u0t6�e���_��7e���>v�[z�H�>6M7l���b]6l��-���dm���F�p�s�Д�2�I����}�&��R��㩨a}�[�U^����6����08|cy8�����p;�U.m'�N<l�Y�Z>~�8�?>^��s��vl&��sؾ�N�g�U�_[󧮞�c~a�OǄ�Ht�H_.YZ��*��Gi56���ӆ�s�ݖqJ��"�P��,�Qat@~)Ę,��2\c-�WK�����Y�!4`a$�ȈBM���&@�iGi�9��-���Q�u�gݵ�y�}��m���b�m�%%)��u�M�����Z-��{a ���i�[�Y�Е��M�F�o�$�e ]5���7�}~�:���ڬ�9[=�nC�O&xN?:�|x۬�4�~�J�&�sp��Y�(+��q�{�1!*��R=v�ެ��͇�����p}�!�cd�=�����8M�t�MA~�����j���U͗Ve��]a0v�6����l��C����ҹO��8���g�~�\��7>�kL+j�[�Θ���1�8�?8�a?�z���vL�>������"ҿ~H$�H$�x��>ϗ�c�g�=�B0��i�;�r��������$����N_��bl0a�l�0�2��|�@Xa+D̔B�9ï^�
T_L��8p����W���}��qYe�ww7K������x�S���8�0BI��\��F�5�iv�'�u�����N�kRUJ��Y����3Cӱ):_
tS����lc�6��|�[k�|�V�]BaiKX�a$$��d,at7�+WW�Ý���M����֩9jz{=j��Fy-c�V�!�'>%�Q�{�̫��֨��֍ۦ޷e�97 ��nEW�>ɖ=N�(1��;���٣@N�L�:��8��m��fV����f��Mh��x��$)v�k]È�M��ݷ��><�O)]+ֹn:m�c�lc�6��|�[k�ze�R֠}3EUTURl��::v��a��g��V~�:�||�x�Hj�M��Q�d�ȍeby�.Nx$>��Г9�����d�,�ݙ�ps�'�6�a��0<o6����T���S,
L�~˓�1!URX�;�4�y���CI]m��ѷN1'Sq��{*�s��=�ƕ����N:q�1�1�c�c��|���wL�o�o����'JJ�����f�o&Τ�9u�N�la��ciCP��"��T8n�˽u�N�	���k��a��
4D�C�*�бϭ��b��6-�5f��j�;[�WR�h,�i���Uh�r	 �	/�~�F-?8Q�)xf���N���2�v�Sh|�����_�Xk���8o2�B�����)�¼M۲ҍ��􌎤��6u8����Q*�fʛ|`�N�ǁ�Y��^"|����l�*|I8� a2\d6[�L�5$0�`&�;�+�(���Ya�%j7Wt�Ē�
�EU�HL'\�N��S���XH�0�.��n��J�*9�����m������ߘ��X��o�	�:Zzq���sCX�m,>�	!$$��37Ӵ�p�)�^{3E	<���.ꨔ8=��q�VYM6����:�H�Ȳ��K�w�:��i��98��\ܕ
��R��L��k�)5�K>41��׈��K���,�I�ٔ�h��=�<�0�)$&v;�⪇=HW��a(쳀�(���rC&���0,�
Ĝ:~tۏ�m�����1�6��׶�%�q
aY�dD QF�Z��8��眄��L<�0�7?=��{ٮ��|��`��֓��&�`�$-䓏;�T*���O�%�Ź4�g*Y?k-�9���Зu�њ�R����r����{�fw�܃��(ɉ����Q�`�����$���'h�K���U*D�z���%��d�繤7=�<ƞ~�?'2H��sri����#��|��l���uӎߜ|����m�1��>W�zOZ7N��#���ί1]廋�D�z�
"��yx�n���ѐ��抪*�����?M:i0[��Z����dy�M�貛nV%�Ē�Ļ�-��]�ĶK���z���G���Z>��ֆ�x��)!�����J�!C��p�d㣁��!��4�a ���;3.\=<
\��[	e,A�/�_N�N�q�>$y�C����t��U#؟p���&͖C��/Ĵ�l�g��x0H""lDD�8P�$�DC�`���blM��AALE4"X�6"l��æ	�DL�	�&�Dât�B"P�b"'4DDHtM�"'DDK0�4&ĶK�4ADЖ"""a҄ ��"!���������n�t�N4�:\�d�f!xHP��6&�::t�Â&	 ��""t_1�cz��<t�8p�Á�<??OQ#����Ó:�2䁠�ܞ�zwË^�孵�N�/��k��:p��-�d���Ÿ��Ba��D�UI�%����R�O�}1,��O�,7�(~�d.�,�e��|�.�f����xa|��p�G�K��$���\�B�;��g��3Rq�g�>n��3���*�	�m
���P�Bù��s-�RLV�ϚT�Į<̣b��@��)4��P�HI ����W�hpʓ�(�$4$�u�p����xyP������m�5L%�$@Rlsb�u�K�(<f)dg��[�8��0��h�^-�������~�\j��/�[�j2�ln�[*M�ٿ�4�n19���B�*	�%�&�E�Nx�1#�P�M �&%�v��5H@\B�G1:@Dr�}��H����S��1b�z��ߛ���=�ۏbgKê�0*��̨FޤH���q�9h�8��i�c�B����z'0��9��!!K:f�=7�ļn�Ql�uÏ4��g���0ݮ��ϴ7\��ȭ��[�����Y�i�z3f��?N/v����ov+8rm���(y�k�?+�uX��]�{ ˰�ZYPpi�f@����Z:R̐�n�Fg���W�������"a�J�}��i��FUZX���$�J��\��*�u�ճ�6�Ma�V�{�җJ���@'ml��_%]���]���ֿ���gz}�{��*��t�����333=����]*�wv������z*��t�����333=����]*�wv���a��4afa㧏1���8������Lw�Vk�^�y�ַ�^�)��r9o��[��Yi�y��*��jT5�jLM
�v�c.��� N�qs�k�[�&���[;�����tn��/�+P��qc�8�x�G�U�kf�S~��HH@=:o�цm�Sj��їu��ul���"�$�2��:�05�i2��~+��c�BRo��8~&��nBt��Ój�tÛ7T�f��%]�Ag�Ii�"g�d:R�^��4M-���Y�yHx�wBM%�z�}�F�^���R3����T�/��&��)��K|��W��Q4�>���p댾���ɒ4Y�Θ<x��ǌ<x�<'L0�4r� ]��L��y��Â=쯽=1\/�{ɣ���yك�95*T���6�ӽO�m4p5�UU��)���'O�����̽��;˝��}�~A��˴��@�6��+���o�\<�<�Yi	m��7h��H.B��ʇs%_v�J�t:�}���/�֗L{��GmM8��E�G�`\:L����qdq��A4OƝ8�lq�6�>c��8�������@��Z/ڀ���F���B�.�G�QNg��3�9��Y�6& a2^����M��꫕R]\���a���'�>#��i���{�p7��q���;0F�Z	�/dqO �2a�n�{���$�#P���ri#%��Y����gF��=����g��G��d�#�z���������*������$����`���|oB���&�4��|��یc����x��<'L0�4n��;uz�]��r��$7ʊ(�C��C�F?��A��i�p^�9��a�����8�ſ��{2��)��hu�ܦ�2NH�Jm�&mZ��;�~3��݋mvz�?K=t��n=��NA�eICE���tp-���ᦓ�t���!�O�ʠ���̞��$b�s:�I����������R6��-�Ԥm�S���FN�3i!%�߲W��3���!��G,�:x��~8p#���7�f�`��L���.4��F�B���"g�$̗����V��Vf`_�a]J4r�U�)��u�R!��]��Ef��ɫX�I\��e�ws1B�j��1p4�I��%�
�̶���M���G]��߸�(�^�xst�]-`�5#�2�3j�֒iZM.�Yq��?{�˝a��g��p�)4VC���r��
z�9R2F���!a���&���m�4>jI��[�u�o,!&��t�oAg��S2��%P��z�aOG��P2��ʞk�{��x���YF�K!ʭ�����is;��"%�:j�q��$"�[	0����;8xh����i���rU��r��u�f�ێ��z�8�lc�1�c��p#�7�n]9���gK�~DZ�=�b���ϣ��'��L{���ª��9�^8O&�4���N'�>V����=��d|�g1�+U�Zt�}�$�&��.�gG<`�P��6O��4^��Ir�<ɑڳ"Qf����wI�p����g�LP0������i���v!��u$�q���2�!m�3$6�2��,��uIl^���g�+⶯]�x��m���ߘ��z��o�8`c��i�./����?i�&�bI$$x�M:i3��E��%��G"E;=Kp��Hʕ'���$��tˤ���O��0��p���[m�M��i���FmmǗf�vF�Zŝ���������i0x�'yUTO�;�HH<|�N�ao[#Vʸs<7qp�:s�h�p�ʕ�l,�I{{�*���O9W���>W�:m��l~c�x�Ǎ���t�a�Gyʝ��T.��5�Bf��爢�����/S�/���9��c���Կa�%ѶV(�l��ڍ��Ԋ��֔�Z�h�54���p'OD��^��_��֦���#_[e����?_$&Ӊ�C�!�i:��k*c����ain{�����pޖ!ټ<6�zHeԸV�ᧁ��I�8�k6|�]���O�����c�1�<xN�a8h�J*wr�	+{�5w5�+�/r�s[tp�2��7�̸ʵ�")��ٍ3
�q���e}>�o��4_Kv�r�,v��Vj��[�.�1+�b� z� ��iqD��K7I=�Qp�����E��YT��f�65��2���/zn~��z9��n\>5S�c$��~:=��֫�*l��y����,8����a�79����Y�Z��ER�d����G�>�u��&~��o3�$��-�׭_�N���q�W�O��n݇8p�ʲ����J�cL�U���;JME�����6�i:�.�B�L'�눅'��^�Wɬ����|A:x����|���1���1��>'�GY��9 w�ݝ<8Nb"ZQUfghq���}QE{TUr�慨�^y���K�L���~J:>��'�z�U]d4Q������Ӵ�24��>JK����	�����3����#�7j���ξ�T6.��K.�iq�	$�a���xM����9!Gd�«J2��'���d�d���m��[c���u���n��F�b͞6l�p�4C�tH""lDD�8P�"P��: �"`�6&�٢� � ����h�"X�6"pN�d�0ق`�&	�`��&�D��:l�(D�6tЂA(ؚb#�"'M	�M�bX�h���D��DDD� ��"'"aDL8&�؅�f�Д%	Dd�����x<h�#�LcLx�qۍ��m���8p�D�6"tD���=V=i�a�q8��Y�ֻK�{r�7$�t���u��e�ur�i�s�w����[Y<akW+ع��s�!��'����g��=�S=��~���+קu�[&���e��䋀�v�:}\ƾ�z�^��w�|��Ÿt���b��$��r�^���dΈ��ܷ���9�3�|o_p�閷�����nt8����?'��'��(�n�Ź���<�ܧ8'�G���;{��r�����z����]]�Fw���)l��Ó��2�𕖯7wݜ=�uRvv�}X�;#��o{��C�+�$sT��n���q]^���77q�s�:�J�%�^o��b�Y
p�/S�!N�^�NJ�vxi^������*����Olk/���f�o��2$||��nT�y�o�����'�_]���|V	����W�y�4�h�.;������P��Fk�ڳ
��7�k`��5��i��a~�瑩)��{�=�����}%����w�:�B���}�z*��iU����fffg��UW�J��ݾ3333=����ZUn��񙙙��"��V�[��|}��h�ϟ1���c��|�_=t�����	�K�N�UUdzݛ>㶦u�����#�-�h�gGxtS��p�p}��?�e,~��6�I6�*Tu�8(���-<�&^50� pٓe��1UTɐ��xT���!�N�|���n���я�~�knOr�m_����σj�'_��0C6t����=~c1�1�m��|ۧ�݄��ݖ��*�g���֧˻s\����B�z�g���i�z��>5�����n�m+�m�6�X�
tD�IԿ��G�2<i�:�I	,:�ԝ�������q8�$!'�>�*�h%�!�ЁLv֟�p'������4ܖL`�HIj6�:���W�47y;��UiQ;��jv]{8/9m����Q�}�'G�9}7յ<=v���z��n>c�1�����6��m����5���?Rj����qeD�i��x�p�h�W�h���I�E8@݄T��۵
2���h�� a{U�JII>~!y��Ɣ�V4�)�Yvɱ���AD��h�%�؎ý��1���P�z��8����#b�h�ԎKIq�mn���̓@�w����/x$_Cς�H�a���&�wx�Lv�UJ��C�b��t��}'����c��굫>��0�h燘~3��>;C��Sp�9��x}�h2��p�a���{W�s�tp�<��Jj��þ�;d{eI$��)���vY��&��!��{�����������>5�aq>8?I��g����;��,�W��<t۶ߜz��>cc�8���<;)p�@�O��f������.�V��q$�@�T4���'�y�$��� ��p&�c�* ��{wmI�/rF�޺!Dl67�|���v/�x����㑟?�-�
�J�F�셻I7vH���*�.m�@O3������&�lz�SSu*�*GE&t�p�h����v᠊}D5
�����rq���&�v�O1ۏ���c�1�=c��V޺}54��j��ٲ�v���?�sOz�'�{é�N�l�o9�P�%J(�)�蓎����*P;��/��^�q;#׾X�K��tI�ٷf'����m�Ki�ӱ��?)���������1e��ep!�%?Cꕗe4e�}N���%�:�On�p��[���*�gR%v��Ү�u-�{�z����4C�:[�m�c�1�����>m[z���?qg~�O��i��Í��I$��5��M��Ԇ�l�
H�>p��5S2�RC�dl-��dTU<�������Q����y���{��V�8|i#�ӕS[�LW�Cӷ'Rͬ^[�G�ѳ$���8�0���SI�:q6n�vz�gZ�UT!*B'6S��-����n;�G�N��n�:p�	��0��<l�t�N3���OEiT��)�W10�Ŋ��|>;WS��\b�Ժ_�R��e��3������/K�/��8]��k0m7ٳL4ݞ���4]�sd�gF��VP/�jVlj�Z.�X�b]����k5��G��}UT���ޒile6�i�����#�jKL�Jh�M����Z������<9�)�0{Ɠ����'A���1�a���L�Pi�uѯx�����cP�4�=��ze2�I��MMЄ���fI$�p��zI<4�q�q0�h�a��v�k[��U��\M:6�>x�=�0��/s=�,Csk���v��fW�e�
˳�?~g��a#��,�$O}�IڕPt�4l���q��o�~z�q�q��1�j��͵C��>c��f�K>e��&n��$�C��`��&��ل|p��>��W,��N�M�v��~��x�]��g5s0�-x|���t6� ��ܒ�M�&��Dg�W$��-�|Ng����wuݕّ�D�XI���.ݸh��bBrc�А6�'�~~6Ų��{��D*�D�Qٜ՜8ںc�Ξ�q�=c���8�O���m��_�V2�+�^���-�ڮ�G��nh��-�6�4���8�	��X��p�0�8'��I��ī9�/�?��Ο�e�T�F�R[��I�-��Z��R8�!0�0�������&��FҜ%��� .&\�eÞ�	��/O�I!��a��zi���-˄������.n�M�����:�@���m�n�v�8��6�q�>c����''�\�H	5e�l�7#�(�aF�Ŧ�Ҫ���5T�M��q2�+M8IM�BQ�;)z=��uv���n���1wa�J��&L��)o�:�I���L=N��U?y��V�}�3ɻ4^03rW���|����2t>q�L��v�4Y�;�i"V_��	�Z/�VFJ�a$�6u>��|[�c���������A��I?L��I$��s�_�ا�����XG���Yd:�F� �U�"d&k���J`�e��@� ���7���"w*ZUX�UeK*���SE�,�b���)eK)UU%�,��eYBʖRʖT�K)eKK*K)e,������YK-B�YRʲ��;�jUR�YK*�ʖRʅ�UeYK*YP��TYP�,���BʖR�YP��RʖR�T�R�X�YUK�UB�*����X�huD�)eU,R��)Ue,��*�K*�X��)UeUIb��V)UeUIb�U�Ue*���,T���*��V*�ʖ*ʪ������U*�*�UT�UU�R��-B�R��-��&��))Ub����UeY*J�J����U*ʪ���T�%T�UUb�RX���*��U��UU�����UVU*�UY*��KJ����UUd��%U�eR�UUU��J�����UUeUUIb����UER�UUQ�HԕUeR�UU����T��J�UVJ���U��ʥX�U����T�%UU���U*�UUY*J�%UQT�Ud�U�����UUY*��UY*J�%UU,UUUJ��UY*���UY*��RUUX�U����T�%U��UU���UUU��'zib�V*��*���,��*��ʪ�UV*KeR�U)b����,T�K*YURYK����R�IUeUYT���X�T�*�ʪYUVU�UU����VP�X���J�P�T�eUX�R�GU#EX�%X�*ʥX��eR�URʥ(�*���-
����������U�iUeU*�ʪYT����b�V)d�JX�)V)UeU,��eU,���YVT�VUR�F��BRXJK%�RTRQIIId���K	F��$RY%%���RR)*E%
J�%�IIF��B��'���%�RX�J�),�RP��i����t��R�J:�w�h�),E%�Ib)*�B��RX��"��B��RX��"��IH���
J�IH�T�%B��Id�K$��RX�K"��RX(�#RIIbJJ�IQ)*IIQ),E%IID��(�#PRY"��%%%"����),���%%!F��D)(),�RT�%��!IR��J�RT��R5$���%"�Ȕ�B��)*�B����H��E%�))�"��RX�J�IH��)%"E���QR(�T�,��,�D�QD��E���QD��XJ*IQd��u��R��R�EJ)%�DQaQTE�$�DT�
�R��HT�"�R��I(��a,�T�*AT�`�X0VP�`�U�0 �� �`�X0 � �H) `�H1D� �`���JEH�T��,,J�R@� �H11R
H�,�J�J�J�R�*T*P�H�d*E�R�KJEJ�K!R�K$T�*TH) �0RF)R�I*Y
�
�*R*E�R�A�������b�b���X�U�P�&��T��uZJ�b�*X�U*T��U,�*���R¥T��T�T�R�X�U*���R�X�R�R�,�eJ�b�T��*E*Y*���T��J�Rʔ�*R���R�X�J�*UK%H��*Y*UK)RʕR�R�ET�T��*UJ�d�U,T�H�R��J�R�JT�R�R�H��J�R�X�J�*UK%J�Ց��U,T�K*���T��J�I,T��J�R��$�`AH�ab���)T�R�JE��,R�d�R�d�R�"�d���R�T�R�b�D��K)T��E�U"�U,��,R�e)K�Qb�K)T�E�X�YIeE��%��R��J������"�e)K�R�)K�%��YJ��U,�Q,�Qe*�QTX�YJ���,RX�)b�T�J�X�)b�R�"��J��U,R�e,R*�QJX��e�����Iib�QT��K)%�Qe*�QT��U$ҖQJX�(�J��H�,Qb�(�,R��R�e*�)T���YER�UR���J,Qb�J,�R�%)b���R�)T�)TYER�UR*�R�UR�eD�B�KI,�b��ZuR��eQhYAb���X��,RX��E�Ib�),R��I,Qb��*�b��(�I,��X��Ib�X��%��X�zh�B�%��X�(�Ib��]�JX��E�K(�),RX�YIeRT�YIe%�*YRʖT,��"�YR�YB�eK)gr�!e,�UE*��e*��eK �b2)�O��F���'�����BҚ
S�?�~P?c	$EP�$�0z5�����W��_�9�������' �4'� ~�������~��������������X��~����������_�?���8���ៈ�~�����h��kI���O�X9O�(?G���~���XY�@�T���������ؿ�@���>G��*�����I@����`�\����A�D?�$4�)�?_��p��O�������Ň�Q?y��TP������4��?��AȔ�����"���(�?�ڎH�-�������RRjl�I��SH��ֶq;�������dW��fl�#��������Ra�I�V�@']<�^�B5�$D�J��U#J"�H�\ _��pBD X�― T�ܟЃւ���Յ6�S��X���W?��~���0 �@!D�Z*��"@�ā�RH&���D�����Ah�I	z!��g�$���?	���s_�?���#������`|�tCH?����'�� G���V����P )?h�0�h~O�#�ƍ���W_�������Ð����Z����w����?Ha?�L� ���~����@���$?�����6X~��5TP�C�������,��x�����=:����@?�?fԠ!��B�a��������R+��V��b��)�j~��(|{��a�U���\8cJ4��j�T���\�_��"G�[3��Kl @ԅ%�����N��D��ͭ	IC��HR���-iC�e����dn&S_��28 �c&��?�;D (�?~S�H��A���miU �`��W�ث���������?a�s�_��~��������E��S��"~��'����������_���E�ܖ��A�[�����_�?�TP�?	��Q������U �?��~כ?�?����/�䟈�?C��1�	�������A�TbBC�g�a"E���n�� ��C	 ������=��L��"[���^fA��~�i�TPC�b~�%���4��C���� �y`�V?����!���8�O�F���������H���?�D� (�������K�Sg(�'�����px��?�4����x0����~�6�?�����2�������F�J
A�),I���������"�(H�ұ�