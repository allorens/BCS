BZh91AY&SY�=���߀`q���#� ����bH>�       ^��jD�"E���ւTٚklЄ*��HP�h5���&�*�m���3ZUV���X�K�h�(�
Dlp

����
4e��b���U��������#Ufi*�b�3�a%�e+e��6�Ll֭V��6J��m�J����6�iU
���n�5�fl�kkX�4�d��%�ؖm�5F���ֵ�j��lh-����*��Z-E�+l6[hm)d��M��ƣSk(��#kZ�K["��07*���[` p  ��oQl̶� �1��j�R���(�k��֥S:��d�����M�2J
4�5����x�����X�j�M��E�   <��i����`4 ٧w ���4 �c�hPSM��>����. 	R�4( n�sCA�]��x G�=��FJ�Y�[`�Vɳ4N    .#o �hз���] �)�r��@(�/Ҕ ��Ƿ�M%M�<q� \0 t�{�t�K�k��Q����v/�� 7��e6�PmZ��d�S-Di��  �ৡ�i80*�CA�ӡ� {��ى�# u��ʝK�ƀY�� Q�d1�: �s�@е;��h>�*����+,���Q6e��   �}�!�U�z��z�3��7�p)osv[��� ��
z w��(Q����� uK�G:����W\v����{F�ljk6�R�4�3c�  f�= )��/\;�t
W`tr�΀�i���Mh��1�Ƃ����: �ӷ�����h4#��(_w��"/-�m���V6�՜  ��/@ w�+�R�7\ ;��s��@ GWt 6�� p� w.9  mи
R� 
�SlV�l�I��[j�F�m&� �z��U�`A쑀�ng@�N  n9�)և:�� Pc(P� j�OC�}{ԗ��ٶ�kLB%32�1�o  wu��t��� �  چ �܎( u  �vv���G;���Pq�W�
�9�B����fZ�fȵ5�6�6j�V�  x�{I�h�� �p��gN(J��� ;�:��h#
V�1�(�t� �        � ʒ����F  � �=��))UM	���4Ɉ��BR��      5< T�Q       �����"�P�    JR4��$�M54ѣJx�OQ���4�i�����x��<��45;?��P�=�/	�lŹw�m�ɸ���J3#�ˎ���M�qO�����?�Up ���@U�o�T@i��G������s���_���|����'�@p������"�*�/�>�'�!�>IDD������7�'�d�a�"����YG�d_���� �P�d:½eN��Y�z�=a�YS����� ��z�=d��!��#�Q�(��z����X�+��eN��XS���T� ��:��e:ʝaN��T�
u�:�=e�X哬��Q� ��~���� ��z�|2�a^��X���E�e^��E�����`^���"��z¾���ṖY �"��z�=d^�XG���=d�z��e�/Y�#�A�(��>�z��d^0�XG���� ��z�=eOlu�z�=eOL�T�*u�z�=a�YlYG�����=`C�#��*u�z����eN��X��0�X���A� ���`��YG���A�(���X���A��A� `^���@:Ƚd_l��z�=a^��X���"��>�:�=a2/Y��A�(��z�=a���d�X� ��z�=d��Y�'�
u�z�=a��� ��z�=a^�ze�X���A�*u�=��YS��S��XS��T�"u�z�=aO�A���:��P�*u�z�=a^��XG���Y&T�*��z�X�(a^��X逘���x��d^�/XG����"�����a���E�ʽ`^�/XG� u��dzʽd^�/YW���½`^��c�#��"��z�=e��Y �z�0!�:�Xx�"�U� u�U�
��0=`z�"�����Q���Y ^� �dzʨ��� �`T:� `z�
��P:ª�� :�*���z�0/Y��Q�"��z�=a��X �*u�����(��zȽd^��YG���̣�U�"��z��`^��XO���4��߃��<���2�@g�k7|��fw��=0�34Vb��k JY���%nHJ{sԆ�7,�LM�.-�P!�F^%v0ژ�kz�E�e����C���a��UJmS�擔��xh�eT����
�(�rV@��i�LN�avFn��M^7���w��k �5"ba��E ���U����W�hYM��\�N��SX8,Z�XaC5b���̗2mո�M#m<���vJ"-y���[���F��tB��&YV9�l�Y��e�{�Y���@�$�wW�b��L��T�l�[�*oЈ6�`:IJ˒S{��LԁVL��z楻�(3��˅ҸEa��Ԭ��DiG��tK���i�37�Q��!:�� �50J����z�@<6CZ��;5�V���y���\ʱ5@6��ەaV�5^�wy�5x�g�}IY1"���Dl�nɛf杭�dP�Ӻp�yZ�Fb�Yi[�/�����uv�Ѧ��2�j�\%���/)Y0�fث���c,��#��ј!ە.�)��%��m���dxWPk����X��g(sN �,�y��DB�u��Dnúӄ��t��˺"m��59��p�Vb�h�cZ��n3rx� t���]3��5�F`!�l*"T�n���m"���Y�n�vS�(�'+Zs1-�u
�L����*ZQ�vM�ù�J,ٯF#�f�(m��T�yU���A�u�W{���I⠸�k�y�l�62��Q�U�ě�j����14(��w�x�
7,T�w6^P�Θ(MZ�%���J��f�Zv*"�;�N�7���{�y�3�
SGE�f��E�w,ffMY#�"m�^v�y��e��慾��b��˘����Gf	B�ZՏqZ�yB�ljG�����{C~EG��gnm���Ӛ�F0�o���4�vHR֤��3HRѽ�03�q��wrS`�6�IڽJUr݊U���2���׊�Vq��ҍ\�Qf�Kme`J�\���]�Ƿ���9<t�p����������Ze
�a9X��1�`�F[v�5�X29��5�-)��jX�l�J���Rm����]a���z���eB�g	2GM��")e��Fm������sM�i�%�DXz�{�:ا�����7�m7%�vC���S �gh��.��Ù9�]��S��n�7*Hҥ0�	ചF���0m�Tx���fY�ј��y��M���ɻcF�\�ԃ)�*�5�,ʓ�A�j-��IJ1��ٰ��4���3���n��f,�V�E�x*m��Tai���WQ�Ǭ�YKm�.�:�mËc�r0��j�ZI8��.�a�0�ݵ�G���H���`��4drO��{b�9&�%�m�!ซ�Qa��Q$LDY�6%)���H�|��Vvwc�&����,q�< �f1r=��I�S��,7{�0�9y�RkjQ�4�w�(�ǁ���� �b�&k���8�VCf�)A8&���	�10X:^:������"�����	a����h����,�M�S�rc��ى9U�`��i��%��7���t�z@!�f�*��!w��	�T[ֹ[V�酮��0wwj�y.�2�3�v��K��fn���~RMh���/]ս�6���WA�C����q�i7oA
�0�:��5�8��|�ɹ�H���E[	DXW7� �z�Lٺ���ȌxecXʦ>@��^��w�	�VVcY6�1��p+/lǶ4���R��D02�r�R9vۻotV��v�bB5�Ƴ0�mȰ�4�5���3�oC����ʁ)h�S��hٚ4HR�OF�*=A����9L����(a��u0B2i�i��1H��E͒a
V(���5[�]�����5�� �g�(��鬒��wi�t���^����;���Z�'�p���mb��5h]����8�jY�2�B�X�S�ld�5��kU�]]b���.�fч�r'1�n�c��(��*��i��nU����V�[�f3�n�C ���[�`�ţ��1+6��k0�H�'|��U���Έ��g0 ���/��qZY#b�h�0�I/i�`c{2[�̻��ͲO\o�),����&�I�P8#̾v9�Sh�ս����$�vC�ʶ����E��wbU���I�0T��KM��Cu;��mŕ�p�qp�V���5���&+�rM�h��-��2�je��mÕ�ҽ�ԥe�ɐ����/Q��a]1��6�9��ܽcoCZj��t����\�F����-q�l�����h2,h���t�ov�����;�*iD�Չ)�EQŎ�
�CK8�����tN�1�Z����˗$�bJiӏ%neAV춦&����4�7��8c��^/o�����]��ǣ#i�2�o�҈3I"�^�gcQi*D6��yo(l�gv���y�����R���L��.k&d����6I�X�`��Y�t]�	�7Mн�z�f˵֥V�S��f�x�B0�r�a.Cm�鉒�U��%�&Y�Y��&,Yf���`��I)��*�"yr�� V��X��H̻��Yכ{y@�2���R�;���3�N��[���3pB�%�Q�U���p�����Od��5C&�Cf��ٚ���nc��pWJh�)�E,�%޼��
:�wIU1/!g��b�d��N왴�e�ȭc�ˡ���Wm�V����w:�Ԫ�b���1�"�U�Z�ٶM�xu0�Pb�2赃2�S��c��H��К�[G W&	$���D�
Oc_P�7R45vn�]��Lf�
��5��hQ��7 ���7��OU%�E[[E��lچU,� E�-m7�m0�)�!��) å3I�S˥�49Y�mU+O癸J�Wa�q��'�l���"� �Eq��{p�o%�Ô7 ei�W+V��b5�
׹{�7c�|^-8`zN4-a�tȽR�=��2٫�8���x�4ʭ"���R�f�h;׆��-kR�o0�E�w,��v��-R+�������F� �8�0�i��E�XjB1-׷.��[ؤ��HcbSX���L(�<ۘq��Uvtco`ys5�rE�$-�)L8~`@�2���jcwje�N,[Yʫ�T��bD�ms��Q9W�mc� Tv�%p8�LSr�,e�X3L���S��.���O��y�ÒncuYCwL�BZ��-�^e��R^-`���N�;�u�/Un�+�3ګ��'+fȌ̕����@އ�]���z�0�F����\�7c�{ʉ�7��J�V�Y'cTn,�Z	�	K������`�����}t�Ɏa91�vV�8p�oh�Z�������[WV���̺Dд���f�1صQ���5'��w#��-��[��wu�"&Q1�(�ŰV�9�P�~�`eQ�3l@��]ŏ.\IYŵ+%�ـʨGmkӎ�)���ɗw��l�NP��r*��c��̬�RB��H\1��	w���3%�zpj�[��F.E�[|u^5�.մ�ehXᄑVܻ1�t=���1(a/
��0�]��Q���r�2���-��)ҘXpK�hN��J�Y�M��9&GROA7F��F�0��������J�.)j#*�!�7l�T��n�������x�c�cɟ]����������&�L���1��"�<[��M˻͉"P�["���Yȵ��R��˩c3TgZN	`E᩻��L��%������B�\�Ȋ�s6ǖ�����O]m�kr��
��[i�� �ǚf8�i<���A	TtI��NB.��mcF�M��yK*!Y�m�/>���Y/!�Lze]k�A���\;�T��$b��YI3��Z4���h6��b5�u��67��X�����ų��U5��[�o�մކ��ki)�[=Y����Q6v�=�6�#Ti����Ҩwa-�>��K�5��t/)d��o�AQ���f��k{f�h�׎A0Iz]f]�EP[��均I�ڎ�X���x	�r�6�ۋ+6�=n�b���`V�%�1+I��^�^फ़ӯ+ �@��z�\5����uaAIn����s����2X��,"����v�r8��D=aT�5�۶	�R�^f�C^J��m��@\a�c1BꮧTUF��قh,��"��2�]\Wv-�S`��\�,[ISҖǲT@Ƥ-Τˬ��ů;��k��[H����VG>�׆��+wT��ffj�ҺKn��i̬�%�[�(�����b�f�n�F)���w&ٖ&!���S,;w�1-toT�t���:�4��0��0Ԧ+BXv���9ux������[A=�5��F$�(� �.6֦�6�\���ń̏CH�ŨKŶMV
�5f(���Pv]^�s�@x���sx��z�5�T��2�+�'C-)A���S�R��!V��]HDb+';d9ٶP�3n�V���Xw3B��`�--��"2��,P.�U�nV[�B��X\��@)�Ә����7lǔ�
�9�j�h�QMa2�����El�NƱ�y2�k(�@[R�e4,���qvs�޶�f�Lf�D�4�=Z2n!z�#.��8�]=�Hz�`-�ʷ2�ۻ����U��R�X���LD�"A2)Nihڀ�)�t��xּ�ж�9oB�)���ණ6M7��N��#��P]:�	�lޠ���V�����Swj�e�)n���e���0)�;>���-�
ڷw0K�:+.�-D�v0ehwL����u�.]�J0��$*�. �����������n��E�F��Q*y2�Q�v)X��\�l�������v/2哏Yx�IFAmOfU,\��J����~��9A�`�n��{�	��84�b��57K{�4�#��L��S{`%eb�Wl�y�%���2(cx
Ʉ*��X@�&��Y��[�h�XE�ERi؉V6����T��F������LJ���^����'i�k�V,s�-�xp�Ƿ�2�٢�ꙙB�+6�&�I��ղ�B�����3]a���ѫ�x�a��ű�S�h�j����!�gwvݲTGl�t]Pz�J��*e%�e޿�c����r��@0����j�2�<
��C�����]�Rf�%�n��Z��ow7+Ҥ�ˡ�*'��RG,5�պuY��vmK8�+Ufł�U��ٲ�챦0eދUJ�O��W��&�>�yj�
��Bc*"�1rZ�7xg�ă�ƞ,��]n-���,6�,�W�X s�{G@�Hpk]+*j'+(����ilő��]�6��L{3[BbP�)�	��z�VD���ͺ-�Y�]�º�Z���T��R��)w�fn�:*+���7-fM�TB�	f�VǈC���9�b�	������-���&���P�N�J�Q��x�XL�qfi��b� ��%PM�r��i�e�B��d.R��2�lFɫw��{�g7f�	�ŵ�w��nE���S�A$�ɲ�ɹ��*�	m-�&k~�ͨj�LH2��Xwe�NT��.F�S�e@V��&���
�oM=b��<���:�留�_S.Ĳ��a�p�8���@j*/7N2i<��kMf��<�`�yn���k3،C���3m,��7.a����`��A�W��`�1)Z��zO�,�[w��D ��<�A[Չ`-���I����ϥ���5����B<�dY�޹+m���C�L��PK�mɛ�qM:S��e��9R�ꌖ�
uW�7�IG�#T�m��m���д�In���Bm�Z�2�W�B�;��/aT��7��ȞI�������J�*����G�y��m��c�&5�sit<0#4���\�ׂ�8iS�os	E�5�JQ����L��<��o(+�R�˲���a��5�e;�Hh`d�6Q�ٍq�۴ X�vm�5�`�YA\S6�Ě�û5�&^lɡ����1$�ʄ-��D�	WX��n^c*�Ov����:e�[�l��,�kF]����L�[R۶�VV^�Ů&+S-[ӊ=�rػ8�+ �t��7o3���B� ���H�V̭�Ǵ�z�J�C.��"�w7.���0r��M�Ұ[����F��@�he\��f���'r�`�r�-hE֜�Ͱf�D���,�"c59w{Y���V2�4l�ث�$ɔ�2��&:�Z���WmͲ��+�-xڙL�Rlܷ�!�+4n�ӟQdeSM�x�;'#6�,-f����� R5�>�$�1��U��0���"W�^���٫/3u^n؎�1���P�{��p�VY5�o7��m�V�V��;"I
,�I���U��M��m����P���L��w��U�qV�k
dxŋ�)
ɗ���4<�rnn�
�3F�������t4[B��(QVL8��eY���kr�Nb�Gw0�f�(��d�KQohl�K��g��+D���C��X��+,���E�eQ�V@$` �Ǵ�\���<��M879��v�aaA0e����jÕ�0:�"ŦH��H���5E����~fpHżu���X:2	����Ć%haA��X`-  �����6�	���.�)`K� 꽫_5�=���Vvf�$,�yh>¤�#��E�&$�Xh<DH3ܜp��(,�+E��,��2��R<�Ԝ-�hh�`Yd��Y�*J�kJ��p�K��fbe�vR9a�I�h�mg�'ô4:��*�^�0p�c��!�èFΤ�>�ϲ �)���3�tv��DaA|4���4b� 1�#D�q�a;B��0�=�y���pf��ٰD�BE���Q����V�-���g��!� �,AD����i�N e@HiH=� ��"��	�um�\�#J	՚�YH�`����'��i����Vv�}�� �����xO�?����$��o��4d�sW7Ga��V��T�W�ũs��r����j��[�΋�6V��*��u���3ˣ���v�$�A���k��wI\�f�XoJ�!�:�v��%R�uЭ]�vn8�[e>J]ԕE�w����d��d@�T��ŖCX�pb��QP�KzU�*(\_kc1f�\��I��l��XݗF��|�y#z��a�&���tA#ѵ���p�����ە
:g�ӳ�z��P�
8���a����2�^�	P�FJ�8�Ձu��i��iі]*�9b�������\�Z�(lm��Qމ�wX�2|�f�U6u=���N�+�s�}��u�Y���"�ޱ������j1,��Ur@rC]�U�Ʌ1�D�t�[����yÜ��s��sQA���9!t��ֵ�YȬ(o#K��jn�`�@�
�D+��I(�uck�S�+�1���o�����M��6�X��0��5��Z��*�W�b?��[7��l G�����d��;MB'����K�JU<FX��;�F��p��-��gnLG Zk��I���t�<�݂�T�35 o��:-N޾�[w�'hĹ�'K�r�g�8�4M�:���uJ3]\͔��lk�O6�Q֢��ꕍ5��Ѭ7��8�>���b�[wuy�d���zz�e��;�)�i[ 4���no	�v�2U>Oj�,-�q���R��*���Y�KI�2kn���0���9eiUV*n��d�����Q�ҥ�ߩ��_e�u[чF��=�B��UUI�|���e<��iˉ� j��BIu+�y��t��q�q4fP��]����U�xv�@�ۇ�f�M��N��BՍ:�Q�p���m��8O�PS)�q����U0L]��|j�G[6��Q��3�I���c�e}��9�P���%�t�fVJ#ב+[���S��w���͎㜻8��Z����j*�����U�N��س�:e�a>�w�Bo=O{�4
��yP�#��n�{ύ�!p<�;�l;���+�d�͚��uڮ�j�^(ƴ�7�*�f���]�(M�~.>�P���PG
(�ߋf=L�hz�ru���X.Wn��}ew8iw;�Y��8��"pB �9[�l��6�IB��Ś�f	p2騢�U�m�߫$}�,ݙ����I7ws֋"{B�a�t��me!sf��/p^��i�ٌ!�V��Z�xn��ykNbu!��*�N&�#�c��\��WJ�<2�:�4[�h;�(���L�cq�����o�k��(ȍ���WS;U]<v)sR��ۖ�R�r�nKYF���)�{Ϫ;6�c�f���Ɛ)���}]��?����m 0;��D]�ԅ���X��%ɼ�\��ջ��SS%J��Z��k�����U@.�Y<��w��V��Q�i�{+��"�|�f�,�xf"��ͪ�'s�r�kVW9�w
U���u�����)���Y][���1����u���f;���-��g0�h;���	��y�a���s�u�K/y�w�i�Z�S4�kr2Q�o.�a�>��uJ�,=T��Oy���,�v��h�Y���H};S�p�n�B�7�+f����|ɲ;2����ZON��
R�b5vC�ol�,� ��3 �3y�l�TL����Q�8>Dܻ�����S���� ��y�y	��dh9G�,�Jf̳G�n�$;���-֣yӐY_��{pGu���K&�	�1��}�!�]K�PK���������ͬ{ʗvl��*{u��� ���F�W�*˒��H��'j�P��n�b]��R/b�fi-7�A%���v����u'�Gi_ �R����P��ֹ]ު֡��p�ӾzE�DX�z�\یPfP�O���>R�E���%^�ټ��9O�'9�8N�h̡Z/9�v�AV��,���qk��]#�o@�pp�n�|�k��O�)w+3��������7��HX@d�R�K��ȳ�WG��Y*s�$̠/]C����ՈÍ>�)R�{N�m��0�D�y������9�cD�*f�x/Nh�K�R�p�Rk6fE�ɻ'7hB��:d�o�i�ݽʳ+3D.������.�d+��Os�i�uc�,��	O�b��m�.	��H��no"���dj�ngj�3E8��V5�+���N�vV���9�S6��m���n�Ѧ�ke�o�=�UֻXH��a햺♳r�5g����U��
�%ID��ѳ]��i�O[��m���9rЩ��}�f��c���C�4�=(ՇyV{�CP�zr���|����GۛuB&b����E졺����p�u�S]�%cr��Wf'-����Z�=o&.�/�/	g2��/��S�ltK�(�e���L�#�q`�3D-��u2Kq�����^��Kv�i�;A��Q�ά��!ѭ{��6tPJs�s �Mv#�aU?�X���V��Oӈ�˃�N���M95�B��y.WUo6�z<�xN��yE+��dԮf��n�gd��%Z;�a۴�ȧ4��uZ�a淚����K冲��s\�,�6���:��3���T$�I��h��}-�n[#g�y�gkM^b;��˳w���h(ZiaD�*k�g�ނ�ݶ�g��j�1.C.�;P���k�R�a��`f�^��b�G�ɬ��;�}K�M}o�ѻ�(^�nP�E�.ӳS�KY��x����%]�uR�,[L��8���E��2�c��ݾ��a����m�#���Lr�c�f�ef���N٫X�t���q��K9�p|�*�T��*�	
�N�Ǡ��5Ip+���kj�.#%�f86�Ϊ��ԗm����gs�se	l�Tg� z��c+�f룑TٕSv�{֥�Å��R�AUt���>�]v�9���J��5g`�ؾӳ���-ֺo������f�4P;׃,����q�����֑5��l,�.鈢��ǝ[K
��_:�N���3۪335wlO�N�Qtz�����Lp/7"��
���И��(Z�nL�jg]��λ��{�`��<�*� AA��x��cR�U��k+N��ݚ���]B����Xt�3�S��	DЃ��6���'��%�f�U��D*T�/Y˓w�V;��+���k,sOC�/��4tf����a�Ҽ�D]H��"���S�/��g,�BB�7ِ�y�+r�i`*dzr�ks9��j=\Yy���$%]/9�v2C89�觷f�_t�6���5��V�Xn���p)�z���9�29�|��A|xLڙk���1��ǅL��P쬝p�c��5�S,2-�wC;�����z�e*d㲠��ג�p�'��c��C9���#/1��C;��Lν��(���a��V����Ŝ#�nE}�_ț�
8�,�-�l^���t�Hs5#�ݍ|_f�n˶fd�7:60m��q�F�\B����͔��\DS��7j�[-�f�y�f�m�J�ۛ�*��1�2���{��d�	�emu�ʡ�L+J�p1P.��ڢ^�T35���w�P<���#Yb��ҎM�b������%
��&4C�v�tU�U=�A%��̚��Ό�.���Ks�{N����M6x��f<z���6Fg����Hrj�y��S�¥	��.MH�/��F�{&(�#WU�wJ�d�0��kSynu��噘+B���S�6
��ls�kG��j���{�d��Ӭ��J+����WjS�27�{�-Q$dVCv�"k�=$��<�1e�_9���9��I�8�
}��{���Ҁ�7fe��oG$��ҕ�β�^�}isE��S����B1b�'C���x$��Yj�[ձ��4\����6	J���y��C�{O,ڡ�78��mT��b�K�<�s޳SBB5��ֳ��:1������#iQ�ri�/*-s냃i+�Y�r��r)�A;��K�����L�0�hQ�i(-:F��ܷ��s������Y�Phl�R�n��2�:y�H���ī�D���^��ӍR���r�TxM�D�����1s�O1�٣k�����L)5�W��)�ƃ/P���dՍT9�+u������ǃ{a��T7o]�g)�96��-�6�]��R��f��达�وs�����jʡ�z�^��mع���r%yp'n`;�uSL�N7��5�j�ฦJ���=�>쨢�҉{�ǵCN���om#�T3���u�[{�̫r�� ��B(���oTOicԤY�"t(�,v�G�J� �@�vߚ� �9�5ftà�|�3�;t-E����7�Zds���vPdc훭�l$�Gf-�KH�n>Cw�؜�9��j��/��N�-����mndn���Xk�9r���j���B��{��ƫ,��j�dSsV̇�T#��U݋B�{�<�.WT� �s#����&�r�tH8��o,r��󲡛���nqw;���L5ԎwsՉ.e;��־��m���3��VS�zKQ�#\зqCH��[6�̘��G"�\�9-���h���wŧ�*F=�5�J�x��^݀;�x���U�B�a4�]�)x��ڎ�yc��\6�$z�A��"�����M�q��U�f�kh9.�Crw|*V����B���R�ך%��#Lr�	8%��5u*��˯MǗC��Nf�0�]u:�-�3y�K5ay���*��KD��؅������7���������T���L-fb�u�yHl��p���FF��r���k%+ ��[�l��h��&�I���w���K����,����Ʌ<���E�s�x��U��Nrz{ۼvTW�Em����|C���Ȯ81�̀�ւV��N�X���t�@��Ѽ�9|����{j��/�Q�˙po��_���n���j���<*3M�%�y�-A&<+ZO
|Z}""��b�ׄ�i-��qi�a�{��X�5�V;U�
&���;�;k�%e�
�vDw���*ۦŲ�*ݽ1m�sa��tM�z�dYA8�<�	pw��v� ��MUw� ��]����gʽ8����U�ۣ���8:�e��-����\�V��%�}��}z��*:ӵ����]b�5S�ѓ[�qH��w��g�th���a����)�U)օ���}����R��s�b���tv�+�SǛ����;�Kü�a��Qr�..�����X9�O6��g�
{y��N
^7����I4DV�p���a��$�}���xH.X�ˊ�Է�ɥ�)=����E�f�a����nݳ+^�j�z�ѭ<C���\ˌ�x:4u��X1�L�ISQ�R��[{�n�l�)�jb���:80:]�X��֥ԫpm��9bO�E�e,����T"�GG4�m��/i���U#Yw��C���5���0>�$`�Wk��;����I����Wm\U�$���2�1Ѣmm����xʎ�1�v3�iKah��v�C@��Z�����-6��̺-c��[\�w.R��Q����Kn,�2�<e��lR�N]�)�
Jr�Tj�&i�}��:��K���Ѯd��[�
Ԯ��&�\*,\��e]�P�1��7up������nvCX��.��Վ�g�;�#���[kv�sff�c�m�.�ɣs#SM��Rp	���t�=zs͵'Z����t�8c�nP�;j�?H���I̋;[�[D��sHr�������(�%v×*�an�;�T�b��gI�����rq�f��pe^��}L^��d� 3k]Q��1^;��̚]kU�Gд�7�C0vUN�TQ�iMN��r�j�q��J�a�8@!�����9Ԣr�CF��Iq�E曷���n��^{�Kj��3Ք�u�q��U�/������������;Y�Ít�YN�A��T�b�G騄�nI!�u���6�WwC*��w�O�u�&	�A^�eI4+za/-��.��{Rq��dꛂ���n��S
Mh������7M��rsYȕY㰴]��pR�3��H0Y�},pܗ��3�v�n9Y��Z�n*��aZ������,ty4��t�L��^Ȼ�s����o%�4���pۧ�y79�� kgn[�*]��K�37DU��v��;���/̩�Xʅ���>F���ӵ#%��.m���d�U1>��;��6�l�>wj0=��Ӝ�B:+���|a㷜�v�7��_:���Y�$_Y��Vp�Q�}>��w���L�z���̼�o�4H!s������T�;��6���L���z1�:��Gptko����k�-�2̹[�	��Y�Rv�.�7L�����=O%�X��9-��!�	���q��ƧF�s�=Yֳ`�W[=t��A�7�8�2��݆��ȼ5Һ��G��i���8�v�1e�����;��W)�����oEt�MU�//TVUr�+�뤌`F�'���R�H��:�W_i�go'��&��rHy��Urd���5�&h�g�8�>�q�KMe���M'$�I�|���]��>d��O���>��/ϼ�̯d;�B�z��@П2��=�q즟�>a�����}��0���&������H�Q��|Ȕ?2�C�1�� 4��c�F��p�%�yz�>a�>{��Q T����^�@Q��������O��#��tU�S�o��g�������ߎ��_����{�����>~=��^�3Q1��sw��5�t�N��i��cE�[����Y�ֲ�TX�G���r:��u���'��۫��c/&���Q4��t]"��("��ne��w��H�b��,p��g[=�!L�L:���[����;.J4��l�:Wo'geY���;����\�lnLj`�V�ع���%µN�%}g`z�T.���Vl����kQ�H��b�U��fu��v�U�|�����dR����blf�L���yx��Uh��9�vU�:N�66���)��ိ�+��x''}a\:�`��P�q��$�����<f¼�\#��x����p⅖q)������9��XꚪGX�\��ԚV�������8�;Ԩ����:�_��v�v�2+ѯ3y�f�c6S�ݨ���HgX��`�;�{pm:Y4h6�Vڌ��]�����C��G�(өX>�n�
9��K.k�B��R��B`�/��R�յҗEϡED7���Qb�Ii�`VX-\4����W�Pm=G2�FN<'j:u�0�����P��Z�V��+
��j��;x�Ei�r]��m�w$��_jW����r%�Y2�
ut�h�Ӌ���,@����|�o2GuS�7K��:8�ݝ%�;V��U�dG�R�Zg�2�:�u���������n�����6=.ʘ���s�#UZ�>�(Δ�ҫT�Z�^9���c�KJ.�G>�S�=���oQN���6�fo"��ğRj��HȇsDjvMk�][k����V�C���3"��0����L�u\��[����m=o��}[��D��Ik)��^F7��N4�����4���՜��j3��RP���;2Ѹ!�x=���Z:�>R����P���Qi�X���@���\�I�Ux���u뗄�qN�i�}�n�F��'T4b.��N����q���� ��B��;n>&��r�v����bBGu���ݠN7Ʒ��8�Xg@�����˷ql�%�a��#��ɼX�K���ffL8RxI욥e�:�*L9g����;Q��WQgFĻCskM���XLUuÕ�W���7��a.�ɸo2o���2q���7+��ڞ/�鏸8`�Ixif��*v���ܻh�o`N��a,X�	�V��D�j�u��POh��}�G����W��I��F��U�[�fE����gMVo�y��%@�������R����xJ���9�� }F씬]�7���k�
��:bk:����%�O�|F}y���C����`㊚�4��R�k=�mZ'��Ruj��A�J���t���^N!�'0[/b� m\�R`ܝP��
�sY�.����V�.58�J�.�:�r��]ǂ�DTs���\��<u��.�:�S�y��M6oFL ��賖%���Τ��'H�&j7u����ao�˱�
NoM;ǯY�*6l	�n5�tcw���f�9�E�x�l^�5��r�T����%m�;
�$4���-��<�ᦇp�;�]ښ�
��©�gr���AZ��
���U��%�ƑΡ���Zt;L,�9��)�5/���׉�A�3$C=K���][����Q�^�Ż�V\�Uմ��e����$��.u�Tۣk� k)ι�>����X��s�f�1��`���R�Q���0��G��r/�����V�W|#!�y@��H�0E����(�k-r�'M�I=z8�;�F��I�o�
6�f*��;�}���XM�=&�����rH[ŏK�o5>xpTቤ#��(`��]�̒�j�>��_nT�T��8�2�Z�k|
�Ey�Xɛ��݋a�mh0�������neK��jÒ��\ݤ�)����N�T!��uK3�r/Z�.�|�Y�c9�p¯���Sk�i�h�/¢�Nۇ�Y���g㻜��K#������l�68��tm�0eJ���"ȡ�|�u�@�S�q��t��[�Y�����e/]Ǻ��x��KI�-zw�Ht����PtV��aM���_���T宅�\!fj��h�3�3��h`�J�2����������PD��؆��.��nXW��֘k풷l�U:22�ˣ~�̧�ʫ!^؋��N\��X��7xk�� ����U<йv���a[���U ��|Fj*��>��&ػW�,!,-Óe6*�%��_\�s_Z�R�d཮ʤBv���_�CW	���p;�M�GJ�%��q��AB-�3�CַؽuX�n��o�uSEr���$̉Puיa�ҳ$���k��k���Y�W(��1M�VER�sX�v�����`�i1y�y!K���:42��]X��8nؤ�w�����ݢ��WZٮ�w5�@737��t�U�X�6�mL����Ӽ�(���r���o�x�oF���E�p�4ZE*�
f��-�x$MP��@�@�bqV+B��_!ף�n�*�<�[�tUԯe�P�޲�t�z�cWK�ŞL����B�f���nq�;��2��w�X#f��W(��|��(��<��u�f�',,p��ua���uWWt���F-7V���GFŹ�l�Fj��.+n��y�u�r�kG�LB�m���t�d��M�
�_�k�]h��#IQ��bV��:�����!D6���oVS���ck�
!�>S(��
ɴ�̛L�'ep�]p�^$���va�T��T�.9�&�|�l�f9��;QD A�n�[P���R��{_�.���`S,�)R[yz{]�oP�ΰ�\Y,�.;�	�8T�۾�M��ִnn8�YRv+J��;�{�I��s�H81�Ώ�NQ7���tV����:�t��{��ֽ5Ս�I'/��Q�Ypɘ.�atE��k��Î��Q�
ꂩ/���cK
.�󺮯-��eZ齶+�ݹ��%5� ��v�ܝ�{4�W�IܛkM�� >��C��ެ�B�5.���g���2�=j3y�X���+���l�D#��,+����sʝs�×_%V�c��ɠ�f�[*���%Ih��9�MĹ���b��`lh6�|��"�Ws�n��h�V�r���F�$`.[��ܗ�I�YL�gVNn��F)cu>�&��x����*��p�*���i;��ʸA�8:�`f�ZIT�
D��]s%�0�n`0�J����8r��c���ia�&�HĨ�	;m����f���uҩ$_hWzƼ��Nլ'�p�e�W�<��E�0Mu��ZX���{��"򜰼ŧ���s�5w
�����O=�<�+LpS�IJz�'SU�»m@Qש���}�\٣oC�6N�^X�{Y�؆��1�M�G.���r�ЂnT�Y]�>]N�J㫶�����l,z�U�)�>�.�T�q����e�l�cw9����vā�{�Y��f3R����5 �\���1�Ge�I���T/K�\�B`!���^n�O�:�z��E�}�1V9mE��$��R�����f��{�b�IY16>��t�s��tk{�ಔ
���x�l�	�GL�{*1�����3�S�I$#XD.�`�g]��q-�+�TPӽt����4`�,ﯯ��k�q��NcL8E؊ξ�y�Nd����U��Ek�+Mߛ��ن�%��c�գ�5��f�"��Ήgc�7)�/�H�*��v΁ޘ2֭]��ؠnIo�oNH�+��L�׮�os)�L�CM��(,�B�#HMԀ��4(m���*�^�Em8z�(ɥ��6vVx��S�2�b)��*EM}M��Z�S�L[��
'(L��c2�e��t��F��g��=�
G9�Z�Xxz��#��9�4��ȼ�q�S}��
	�s�Z�ksd8�B֋xd�3#T&V�u�u�O7�΁�!3��mE$\�}G��dj���u��i�ѴF�$����H\ogkҨ�����a��hޘȨ�N���6+�	��_6���^,�%�G^%u}.fYP�������:kR���:Sǵ��yz�Qb�:U3ln���`CiD.4��}�;r�n��͠�7������sAffjb>u���Ԉ�P#�����P\�Ҁ;���T����`'v��Y5z:������ErCr����ƁZ�J����	�Ա��d�;�v�JTe�J!��͜�����qw���7F<f8��9(.;��������t[QY�v��܃��=��m3��(�5��8�X���f��:���ɤ�����rī�zr�(��q�����[�ݽK����h���uN�Yv�co6y�
�߾�{�t	��8+_{�;���flj�nu�s϶�T]�R���-�Td�΋����̩@<���In��e=���+�x�:�
�C�u��aފ<�����9Gkh�Ĝ�j�F���NN���=�RT�4b�.-�D�'+}�g(��&ȥ�����,ԅ^L�We�xƽ��suSh�)e1�u�e��Dy��^��$�iŌ5-��
�l-��i:�ʫ`
+}�T>��dZ�=m���}t�5`F��'C��<�����fV�j*4q�"���9�70`�yX�:@�j,K����H��F�b�p�Ybz�:\�t�ra�-v����R1�.�WrÆ��.�U)X�ʄU9��o�c���{l���(:�彈�P�Bw�X�Nʠ�k �|nvK�]uQ';\Ǐ�8���E���;:cu���t�A݂�I���D��PCM>�x銣�ك��#��5q��P�!;�9N>N�� ��_-�g�[�!LY���.P���Ս�|�ˮ5X,ۋpv3�ዣ3����K��{��o��Ta������ �iV�պj"�B�eX��cHr�X��j��;Zn�J�l�j�������RA�����Q��!ѥY���f�Am^!5*�].���E����?sH�Dn�5-g���h���B1����7��6r���s����B<��v-N��e�ұ)��QUm���o�&�؜92�d;\�����B��wXJRQᆫ6�*�,���!��#�bg{B�L�o��D����>�J��|�'��i��L#�� ��E
�m=]/"I��\K��覼 X\n7
]��V�4VQ�J��9�g9R����i��&-I[x��b$ͫ)Iݯ��ؾ�������e`�1���dv3s/���9���$�¶���Lf(�<�ʗdN��ӝf�q,(:�9jYKbX����Y\9�f�-�z��,[a|4U��CY�g�ę)$��UO�CC�8��;g�25�]&]Z��e��r,�)�np��H5 :�&
�.�G»�MZ�r��M��2��Bo��0���YTŕ�^��b���b�/�4hN�(e��u
aqw��z6�Ǘ�׍�/��X�o�U]�]hL��K�؄����<�5��Bbac����+�����rX��7oԙΰ��4Lȅs0ԍo*"�y�ʲ����n͟n�ja���E�)f$��N�!6R(�cy�*!G�������+�0�:���ʈ����I��j��.�Ӓ0r��lqf�l��/9+��0Iv�V�a��7���	�*-�f*�g-ۡ��˃���LLѪΛ��]USo��q���;��/,�J6d'�_mi���:Y�S�y�2�I�_�}�Y�0�5�T�3$jVʮ�ld[6�(Ķ1\Ŝz��� �-Xzh�"l��x��y��s}]�-�DB�m�ob�8U�5�!��d�%m����o��;	)3х��YS��5�Utdso�<q.	4T�WAN�y�j��5����Z��$���E����L�7�WN����k�w]�i��@ͺ��p�y;A��;Oaͺj���Eт��ݎb2�Sm�7z��	�7J��Ʋ��f-�	��t����{�խZ˗�%��#�=ZFù��1��GՙL��\�j�B�J0����t����d��>��ܧd�1�:�q����ܰ%}���\ ��q�FG�3zNn�mf(���rT�x^��JC�`�����S/"Tގ��'&N�'�9��:��X��˪̥�	7_k=�rz_*�gV>N�[����XجGSQ) ����a�B�3��]yΌ��[�m Sz0;�ِ̛}@�v�-<��O	p�p�Ȇ��E���z�6��]fَa@%�]����E����3�"���EuI��=������nv5�t���t���
��u
ֆ�Z��}�/���c6W����(!�Q?��ťZ"A�7:��Ɓ�Ŷ�SӰ�0�N��,��e٬n��5�A]!���9�]g8��_���u�=��ڐ$;(r�ʣ��BB�X��XHw�Q��i��)��U�|Sg&j��8gS�Ո�*�$�k��e�W㌞w�6o�[I7����27e�����k!�tr<�����h�]���X�r�+2ˬ����c�����2dy}$�l,T���u��7y�j+L��Wڍ�`���MUr:46�/8�[�Ln$(]�B��Y�|��o4�-�[�e>#��s�LlUGcIv��;![�c]Mc)�;ˮ��t���r�ւ�
�`�ݾ�ֱ��u7��~�Ņf5]�Û
�T�����]�{8��uP6��̴��.t�i��q[����\�t����r[ܑ�/����=dR�/��"�j"��K�]��r�O���2��YΆ�ܮ��gS����㽁�_wl��y6�B�5��W���{�\�o.o���������������������?!��������G�|||��|||||}>�O�����~i���`�c��ߏ��I�D�i��
d� ��^L��2 �I5��J&Z`��E��JE�\H"J!0 ap�
�1!��v�d*��e���$��ѱL��Z(�bЦ�w�=M\p��`G#�IH!fw�lC>���{)��w���T4
ܭ8X!v�ܣG�E#u�u�h�s�GI�ʔ���h�*6.��m:���9=�c\��q<s��+9�FVo	V�_�p����E�w� �/4Vl5q�
���SӓhJ�j8�s�ۨT͖�lj�Zw����=%��E�˧!.��F6o�u��<�dOw���6ZU���__�v�j:>�:����Q��趣�7RY*Xѥ�$4�D�`�c1N������f�
Ӄ`�����{Э3>�\��͙�bNP��q}Q�����f_Л���FM�^�$���;+�!��ΐՖ&T*�wn�Q��kc.b�S�fH'J຺��O�e�i�c�&�=����<ټ���B�:�5�ゎ���ͩ�U&1��ګ�U��W����oa}ͻ�u��A� Nǻ9��e묳H�`ݾp��ԛ��A��8n�pd�p�E�V���)]k��*����O2�8M��:�r�P�؆V�/B��!����}�3|�Q[���w�`�xQ���:aY��i*cZ=����*q죳�TҜ�X�1oX��R��H�R��}��:�������%�Bt����y�(e��j�@�=�$x����>(1n�
���K%��7��@�Ow��"�-(\�p��0[�4=U���ne�mp���ڤ�I�H2H!G�PM�،�$B&!(�J,��A��qċD�	��4L�%y�a�8J7#q�I	���Sʔ��l�a�4�r2`��E@�
~4��J$�@#�	�A#`��h)
e7j �D�J�m�!J2�EXm�!(��~������Ё6 ����O����h��1��i�	m�!�Ē2�f@�02��
q!��IBP�D�!HT)��5P��A ��x�H4�0�a��
$�s$�PIy�D�+�	��A�4cj��j֊�`�i+K���c4�m��Ky�%\ب�lE�)�F�%�ō�-�m��>}s����Ѧ"��j1V�Q�kh���ōk�4���UAF�-�6ƹs�L�TZ���F�D��hˣkj�b�(�٠����kQ�h��h�b�6խ����譢���u��X�h���*.N���6��'��s�$�Ί��s*+s��&*1����h����r�cLF�n\�&�F�j��m�im�f�1�m��l�T�[�lZ�VËk�+E�I��j�[:�lVs�b��I�Ź�5D4ID\��Zt�D`"�T[TZ�TT3Li�i�m5Q13i�%[܌W,SG1���F1f��Ê&��&�!�X�:�QMTܜ�͹���M{ü��)>�H!z�$ ,��j�5���8����X���!��M�.^��gױ�+�Y-a4�9��d����[W�5�6��c�Y���ފX�����L�Ry�X��`�pG�Ԉ��d�h@C���!�(�m��W�.���Zz�<ʭ�^����d�����*{�ʟ9�����f������D�O=�}~��v�iOH���Nm�F�i�I2(��z�neĽ�|�]���o�?{9W?F��}K�>��_�3�w[tQ�ŉ3m�Vd�w\ue��#U�A�s>�g)�x���`m����I��$�ɶ�4��,kM��8��б��X��������_�>�@��"�!^+*����e�������<F��Y���%�A��Z8�&+���=�z�:Ǎ��t��k�񳷂v���O?�z�J�hyfv��7����u$�/tT2�������=۾O�=�M�t��AxG��n��6M��%�����-�]h�����U�/?9qH����<=���V���3y��7_d�������T.��l�_gq��^��pN�Ş�w���/B�aD�}����NQC���K����Xy���餞��m�Z�S���і�[��n��萙��w*��m%P�N��U�e+c5`�`�F`�˙%6�m����%�����Y�Z+��=�i\�r���[����E<\��p9U�!���M��`w����TH]�s#wؓ�Ļg��,z]�ُ��c5�P�`߶h9{Ԯ����<�S<�]^��nJ{���	ʗNJ�g'����	w��E�ePKrw���\׺I�{�ٯT|�]�r`�~�[�4��B���(�28=b?$��v-̸�}z��x-<=�|����:�Ǿ���&P�Rn���ws�<����gm����<��O`�L�(賓�{�������6����3��=��2�
�5O����OT"x^]�7'I���\F&��M�V6��5,���#��66ۆ�������>�Ws+{�F����;$�e��RΡ]L�Cެ��Ҏ��ķs=�$�O|9W�B�_3���*g��
y��<N�]J�s��﫟z:�E,,;gu_6Z��H��JfP@��'^�Q��u���˺qܥ$�P�:b;���:�k���kx9c��Ϳ���GHN���|����^u�*h�l<3"�=/���Ec��^��u^؊Ic32_0vC��KB���(��������s��R�+n���tye��[�g�C��a�^Ď�:l=�w�c���ӷ�o���o�qU/
�Cް`v@1fN�����H7�	�f�l�e�:�����:>
���Pn�#����;��}�Ճ��PV̳�{}�����ك�-��/�0��{>��_�0.Jg���uI����~�ɢ:y��==����S�M}� ���`��g��}���>��wuL_���/e>�Kx"��4f�?3H:�*�wnͻ���r7U�3�D������[I�`	a�V"3�zf;Y�>���W�M��"�b�4zY��Y}�r���Һ׵v��:���N{��s�s�\�X�\O�o��k_ِ���K�ޮ5{�ו�=�y�o�ϣc��,5˞Tw���롕������U>��ۊ�ᤂ-�9�&����uM���`˒q���԰ѭ�0Ȥ9���m�r���3Y��i�%��|nI��*|��J��[�-g:]�3]:�Kڎ�iz��uY+kX����&���|���6�jo��"�i$R~���H����kC[ �����{ӫ`wgf��h���;.�ii�\��6
��/&���y!��g�����j	�;w>�G����&'�y����iK	�w�U�;gOC�g`�,Y�B[p�����^n�k��Qx$�>�{n���ַ���棺��X�o=�
W���[Lr�l6/��*��h����%������{��#�ye�<z�.���^᳹G^<{E����&�yץ��E6񝔶^�q{}j����N���>���:=���}w���̛�~�J̴6v�=nٽ�g��{|�=�{v춸ay��5�4a&��ى<Y��:�L�gt�[���H7���)�����N�&�7��/�{�w����w�};����Oa~~���^�BǢ����yG�,�V�
/ey�}�X#��������x�Z�Y%��w��Rw���-���u�mRo%u]e�yt"�H���6E��,rB]�؎���5Y��6����W�wl3��U,���6ȴE+Ҝ{[~E��Y$	`������A՝N�N��|���|�h��p���'l��Y�تfwv�U$���|�Fn��l��s����tn�:�)%vëW�E6k���Z����}ʕ���5R�� �j����͜&+������\�6��c���t�~���F�4��V�tњ�o������?1o�*�澽��k+��?{�'�z�ɗ���{��ߚ��o=B�m�0Oo�?C�j�3������h����WG�	WUOzڸ��f������踩�c�^� ȣS�	�2�f���ɟ:�~x���f9���i�Dl;؋7�Cё�x��f�I�={��2���l�.Q���S�&q�tBc�:�A#o��x��KtD�ͽ��o���~�����O݁�3��l���o*},7~����KN����n�p�_\V���$������<N���w��b2N��r�Q�$�iȮ�4zO�t<�>g�"��W�<�<�]��8��7�{��^�:���*�q�����e2c�ze����=�5q���K;a�ah�^�]6��`��u.���H��@.f��{u��hj5�PM�/���9zK)���t�SX ��s�c2�Z�w�URq��r�jm��X"�'t�s{z8�t�����v4����{��}��W�����:�{/Zs�ך~G�-��LE�����o��K���L��=�i�I�Ryř�lQ�gz����TM�GOx铲Ov�=�5�Zӑ�2NG�T�nz0�s���ϴ�����B�����w�w��o��6��G�\��X��qE�����!�4T��hzQ]�n��<V���5�>���O}��*)|"3��Q�?!ҏ�r�%U�������\�4�_�r*䨆j8^u���y����������Ao��K?g5���g�\�=�ҫ;<���Ԯ:�ॺ�y�k�zwʼ��.E��6)k0����Y�ެO����ngfvE�V)��o�zy�~Ʊ�<�1�¨i����&�"7x��Ao,��i9}i�O��O��2��J�܇X�/&�s�D+w`�+�^_�MnL����յ
�à`�	���>� *C�-�]��(-���Gx�2���d��:�sS����C��U0��DI�Nҳ���Ծl�׸3o7��݅\g^!��9%l{su�\]�}�x��/����wp'��r�o�V�>��ԏ�}��uW�6y�KA='=�I�ꮖ1-������&|s��K���TO'I+�8�rN�A'`��%��Z�ΰ�/���:���=gK���'��Q���[��>�q:���&A�����d�0���6��yzr�Y7@�y��X�o�������w&y�
����{�c�4/3~��2��9�2,^�_��C��}�2g�_�w�;Qcz_�z����[ZG���.����C~��r瀊�40.���oۮ�{y�Z��ӱ����x�u�SkLwv\ܐ0驠j���䰟e������X]��~�=�*b�Ol�Cb�,��W��Ә���;_PA�z�y^,"3�v�^gT���N.9<,E~�R���������0MC5���37��m���n[�R�K�n�Lxr�t|�	̃&-��,�1:`t0m.�ۣ>y�w1�k�s��꼛CR�^nu95�Β'��ݣv�+N�����|��jf͔u�whcM�xf�����[+^*�tؾ���QT�P�.��b�nA��.�����t�.�>� � �䨆J�HU�ڶ{����zM}�a� � xo����眶sdwl�`��,
p���<���K�Υ�M\>Rr�ǰ��W��:���M-Ɩ��:ez�	��&�-����'����:�.���Vh��ޭ�'$�[c�W'fz��oi����>��r�� �s��ՀG�>Y��h��*��8_�V{�y%X�(�5�w���=��_x���n��_i�Q����"�LyS�V��������&y�t�>0j#�>�і��}:�I���'�נ�M�uM�69�5��&	���p'5�Qx7^�m��ݒM�4�'��³l���mלMG�x�v�� ����\�_���ϲO��]�MSwb�}^�#�D���)`�
t��yT��7r���;��68�)��}*�b�ɽ���5o�����_6��ժ�w.�i��t�������K Y<�9]��,ǃx��o�@L���M3�r2��މ]�]��˗��p�$x�`K�+U��R�j֌�]$-��}�=�Z�]���l���H	_;���u��t�YQ�,�����lR����f�zOD{���j��A;<���qB��!7���j~\q�y����{�otɜ���n����3p�o!9_!/t^[�ּ��C"�����D������J��г碜5����m��j%��|��ݾ� ��bu��,��zo�/�*�Io;E�wB����ѹ�6{��0�%��;wDxz�?QZ�Y���o*V�L\
����o�׺=�����W�`k���?�J7��zrvm�O��^���^\�5ȢxO�#O5�
3�O����+����z-ʣZ�y<Qw��������&Oo�?Az���O�<��	��^�H���Oٽ=q�&�(���v-��Sޛ;���ן��k6e�/=�v����)#t��Z�c:w�Qj��{��g����xW�&�4��(����֬�W|�W�.���oa�Q����y�⫡C�.�v�(��w��2� s�w*�k{`�v�*JFM��ʨR�4d-�'V��r�l^f>�"4��C>�N��z'*�Ƶ��WD�a�R�O����:����o��?@����D��ggͤM�H�����6����۝<�m-�K�ޮ4�ި�W�_V��]5�.�rOn�;�=70#u�G�`��3�I���j�9��uW��00��aV�K���u&�}�ƺ5��nI=��dY���t����z���~�t�v9M�����ϳ�d�;����I�
��?Y��3���iP����q���o���2s�2(�d����߳�ߵ_�8{1�E%9{���T�P��'�ߨx�<��bɾ�qd�?=���i���Pq��[s�o�o)'�}��ږ�ã����k�k�{>�����^�b�aNO<�D�{=�Io#�3力��Ĥ=(���Z�9rB��}Oɞ��瓖���T^:F�vw=��WO�}A�}������ X���7��{���w���ϏG���������������Ǐ>=O���.;`;�_ٓl��<U'�Y?f����J�	G���u�z�ܸ������n��EB4Y�$��T��DY\�@�AğR�����0ƶ���<��uz�@���u�,�2jE�;[��xA�maM�kU��2�Qݡ���1�e��68�цLu��0%�+`E��nIwOA�2)z��K�s&�*͜���gX���;�Ծ.�����wa�0s4�*99Ʌ�#{|͊mܷ:o7����W�Mf�7LԵ,q�����v�E�CS�ʼ�}z��Pk�a�fj���
 ���X^XK���dSUy�-�{��T���W�gT����'c&f�vsfS2�̬)Fn�:��V�N0!�n-?v���_ta�������sG�f6Oma��4�]�k榤��M��t+5Ӗj��L1U�I����l�	N�;^��=b�յ��d��yt�m�a}�_��B:�f�N���-S�D�]E���_wr�iu]@�b�<��gYH|�K��ZNe�9웼��=)5���v-ul�q�W�᭔�|��*w�����Q�}Wm%��X���ݎ�4�9�k�z��d}��d얰nI��R僨�OR��sh�hR��Ե)�Fu�K�����3A|v�ۼx]�b����X�el�z��a\j5+0b5�r.�����!���Y��ӷ�Kwsk$�i��3%i��
5�Yٻc,S�	IƑ�0\�� �p��c��H�!��쌺�t�7�HTR��,����2���b������=]=��7<w.fum�vol�0-=��dVq���_jgt)�cc��v�l�JWR�#A�Y�|{A�`�Ý�Z�䇚�D����f�N�²ҲspvJx֪�ij�'������spu���P��ew� A*<�'y�D��'��Z�G��eep"*Cru��8ӑ�v�I;�k�b�T��ZAl{��P�5��n]���h�5#G��evdS]L�V�IZ��g*�[�h�L?T	_u��}�ǿ9���X8��u��G&>��D�؜O�3�z,b<^^�f��
ܝq�4jŐj/a�B�dgse�gz���F��ظ5\ȃm��O3�wa�y�[UO�Y���]4v+v:�'��5�& �H�����}<�y�D®A|���{�l}��������Uvi���q����h�u-d�5�d{F�mVt�ؗa�vq��r�]�;� ���*��Ǵ���ET��}����&�
%��;@_f�h�K��ה��ҹ�K��N���Isa!�E�PLr����W��ZWs�uXj�+5�id���&Z4��a�	y�XKx�%�{����Va5%�}����b]�ۅ���
w�e	����`�vu[�Œ:r2��u���X��Q�Vc��WQ���A ���ڮ�D����H"I>$�H?2c�v5A�AA3\��Mm�X*c��Ab�lne�\�H�Z���)�F#\�A���kn:�3�m�EU-PSU͚*�b�xE;���Gpz�"�Z�V嚹��S�Am<�8�UL[b&�Ѣ�Z���*�A̺6qE3\��Zu���'�Ƥ�m%sh�]PE3��(�2r�F�傠(��.lEEbng4�uQEPD�@j�9W6
�b��j����.m\ê!��AMG,�r1EDU3�J�0j���h5�#�c4�D�͂""���M�[� ���X�c�j+C�����"�͈���5� �*�'mDէmj(�꒒�j�kƊ
j�e����F��5����m5USUQ��
�mAQD�b�Ӣ�Elh���Ţ(�mQ1kE4�lj�"�"l�[m�N�]�jb"���;g@j��!��o��rw0�"��B ���������k\�.Z1�T�N�'���|X�yx����t��c�jCZÕ��v��HK����r���ƃܙR�I9Մ]��:<�7_6:�����T6E�4���snbp�9���#�KS�5��ph1��X��Gt�8#GԌ��Z�kt�V8Q�uƊ�k�Sl6-š�\kH��<�:���g��k��Y��>J�!C��p���p9c��ZB�oO�+�Q7W�ܦ���������
b������W��.ܒ�IS6�Slzv�^$���<���Q?�{{��@�K��s�0i6!��}.�������W;��"Sc{|��a��ξg���]]�1��ū	�.��N5?��/���80����E]E�5�@ղo9�t;���<�js�w�����!�Y�'���)��T��#�����[���c#)D�f��+�񕶚�-���{����N���>�N��~�O�p1��Y:��E2�������j�p�yƬ�[��d�e�Wg|4bf�}P�a�c����&H�_7�c���g��R���j&0�w��ܠ�Ϯt�Td��C���"��a?�j>f��|�j�cn�e����s��M����y��5|�m���3L98~�l��p�s���_g�[��W5�0�� 8�y�8؏�v�ة���]�؊�B�D'�h[)�kMZ遫����qP=H�G5*�Q[`����\o��ň��k��?OcM�X�,�m�U�̅����(�v��;�_c�f�x�}\�9[��������|�Y{dQ��5:�Xj��`6��T�z=
�:�������t��v�61�v���`������ȝu�[���J����'RO1nM��B����4�v}sw*��h�c��A~ഇ�o(����oqj{��}�����}�[�+
�����/�����^5����}]`�sH/�������Cs;z9c��2�ӗ֕mn���Yژ���;k�Π��%8%9�a\Z<׉���1�W��w�~�nI����)�n��8Έ�gh������N:���oH~~;��P�]���1i`��1I�L�G<]�-H�{���6��`��l���>u��d��#��	w���Gf�U���;����N(��Z��v��-n�#.��}k/@��¡��jw�0>B1�=Ű��G��v������y�^sR��E���\+P��r�W�3���l��3��zw�`ǆ`t�!����W�.o)mZ��7�����#'ְ0�	�Z�,��H�3�1���/M�c���'���V]���k#5��݁Iq����L�|sϠ?B����.�,�
�R��YS�w����O���d<	�5i����:���1�>�3[Df�iٳm��i�����X�e��V����hݹS*e�{=0g�k�W|�U�k0p���k�/<s^��ko[p&�49U/�E�v6�RZ���îV���EY�c�O\�ׇJR�3n����m0��nZ��Ôf����(]��Q˧=�r�����7{�"�b��̦��L�K'�/�9���f���Iڇl�''[���$�Xs�ZF��R��oe�Gs	#_��U�rm�ݷ+X!�-�V�7��cO��&�[p�����T�g��LS�O�Q��Tǃ(�̞y]{���C�{�ɂ�3����o$N;j��"9�v����#�Gd	e�f	K�`b�z���9�{vL���<�1�͈���\��~g�/�
}�����i����c׿�6�ȫLI�����C7zK	]�����)=XJKva�4'�vm�|{|ɺ��8uf�[�b �ퟧ���H,F��� ĝqv	T[�gG2�ְ��o��NX0`+
�
��vڙ�t����
Sֶp��^v�05�wo+d뎲�+�҂^�¨��F�p�:�gN�������a���w�!�Z`>�ja�d�qz�k=j���=�Z����_˹�*ٙF�Ot��s�c�Yu@�U��_@?A|?0�/�����]b2~N�a�wݹE�e��zD�7��۶��-Rͺ�˱���=�-���yw�xL�?(�,"�\���=��CO.�-����]{+SӉ�o�����ѓnⱋ7�7�q=���A��7f�Lv@vd��#�̌4/��HV:�'�������U"K�V���{���^��Γ���o�������G����q+���7���l��uMJܒfh@��g�i?7��ˊ���,��1����)����H:"�s؛�c[π��B,���2�4bE�W��2j�UE��X;ُ�<6�_Aʨr����`=0t�ê���%���h��w��ݚ��`���q1w5�uQ�F1�0��L�|�1B�Хa*-�`��8��D�y�6�<�Q��tS<h���0L���#�%bv�����׾&|+FD��-Ԛz��1����7��G�Gm�S�;A
-�8��S!#���i�y���żf2�dM��.�Y����6�R�&�!%B�F�c�m�'�|w��-�$�f̘'�ƀCz�:*�f\��^�_j̭���,̔�ĲS�X n�d��e�>�\S��c�k`�a�$D&�\�+ܹ�im��0��;{��)sZra׻"���J.�<��ӷW�r��\��l����r.'3b�vxZf�B0Bn�Ln��B��P�xU�� �R~k	Ai��T8ԜK�+��讕Κc^�wv���0�W�2j�#YTħU�,P:v��&|����ds��R�;��|�N��>ω�A]��Y�ћr��Z�lr�`�_�y>�(0��X��ܐVbR�!��Q}�qp��G��>�gY���e�����+��\��bKX�X�(�,oiЬ��C��v�Ժ�y���W&���Cv��a^�XuЙ�]��w'��5�@�4F}�}ġ�{8�o��8x���4	B5�O�\z:��[�-l��=+��w�V��ۺ)n^*���&�4��q�!]�6��!0P� ?J��i���j�872m�{
�:��l���2�y����KX�xT�a���3<�d��hņv2d8~a=�D�+�75O��ڗ�u<�<!_n�+�����w�P9%?X/��W�v�LW��fmL[ ��d�wA�xWSf�a��:p�-�z�pλ/D���:�5��^dn�0v�wA!�@"x��g����5���D[��ꋟ[ǚ{��:F���PX	����:����;�i�(_I`i+��R]÷�`�=��o�n#�c���x���p%�=b9��a4�22��T�y�ۓ6�5%L�cǐtޠ�y�B�s:�'�f=�9��q� o����9P�V��O]�E����*��7;-��B�z�62�մ
�[۸�j�%y��l�YFi=�W�P߽�LH�:���M��,Y�:���$8��nD�ݎ͚�UZ���

0�f.�q���I�1,��������{+�)i8?1�yz����w:o^���5�	��}��^]�T8�x�J�]�>���;F?+) ���\x�E��A�z��K_z�p;���N}���7���}�jF�Xn�rƦ��./R��R����n��R�]�FT�ò�8����w�8HX�]J�jNQc;zW���RZ��.���Xg�,i>f�'���S��^���,P	*Mm~������-�����ާ��ʷ���>C��1i��̪c��d�#�L8��F�v.�)7H�^[E�0�f�a�>]�DoތakqםG�g��h�yЂ�S'ry����w�Bn��LZ~O���23��(�l�Do^o!�Z�:�3L �vG�G�L�k��ߘ��U����U�m��O4'M�W(׃���� ���1���X�:A�wh�;C`t ;�h��~l=_Nq����n�u�3UWgqچI�k]?1��&ޯ����U,�[�f��`�p1��_��9��i?i��z��|�s6❺"d蝠��4-�Ë>2�����5\ź����A��F�yÀ�����/k��
�����!��Ϲ�Ļ��A��i'1�a�Z�&(��1��%Ҏڔ�Wt-����_s��z&U��������8��ԍd�z����4!�K�v�e��[�mU�a\j�֨���V�������)��c��/��3�?�_X�v����^�ȖG���]���� .���7%�(f1��G�馇~��j��H�ndUL,����콠msТR� s��N�6!�&�MpEx��;��d�WV`Gq���dM�]|�����1����mP�v��4�9n��*�����r�z����`�A�|���cr~�C��<�{6��:a?.g��JF����~򍡩.��ԟ9��l�w��B1���E��U\���F��o	���&oq���l��8�r��PjHγ׳gV@�t���V���߳Qc,v��a��݊i��H�~���c�r�1G���#6�_m�^���	;����j����Of���t��1�/K�'�C���W2l���?B�오�}���W��L)�\[ �+��v�ң�����_�4�O����A�k�I��pr�`�����$��1)�FE'��r�D��R�{;��o>�F0G^�~�~��mw����n#��tCgu*L��uq}���S�o���;���`0'�I�pgם��N�AƑB~�0�v@�M��{�$�'�F&Wf�e�m(m��uI�ћd]`cܠϿ6�q��D�\�����ڑ�r���L��W=���v���Al��+Ee��a<rT{�ځːzJ�v��&�/q�D:}�S������ƮN�;�p,iwǞ5��B̀bN���*�
X|h��������n��?�WS����l���5��G�KA��ygV��zT��SV�ww
�T}��^�wX�/6ƺ��\�\�����f�h��.��ZrX�{�l��i�x;������*o��w��Usi��N�$TނWj�Dj�L�`��������7�w[�\�������,6���������4-��̝q�_�s�PK�)~o<DN���+R�n������;�����`69��s̳ ܢ�Xԥ�ħ�p������
n�a^Nj���
��[���az/a��2%�=��B���M�h��_vlGO�Y���n�R������,�m��b�'���c��&e�@:"�׺���>�����28F��<����v�E	+.��}ś݋[�i�a0��ޮ����r2�'DY���-3�P'���U���U�r����ۅҵ�^����H<�\��/^*�p�dy�\m�j�L\:o@�}�qU.�n�r�xN�f`���*Dc����&.���Q�]~��`-�J�����]
V������p��mM�vL�)R377�����
��z�lP��scO�L|�!�s��b�`�;R����%6i2kx�=_
�8�.y�֬Vww��BN�]���oMl�`�ҜI|����;(x���<�84�d�"��3�.sq^������(��Ғ�5BJ�ߣg1�_q�P���C�h�t��	���޿_�x{x��S˜���������.ea�Ш��ߑT�Ò����vi��c�3s�r7swcq��SP��z�&�i���	�ʽ:���Ʀ�����9՗P�q��d�	�ؖ�q!ޫ&�x������97���R����\��j���x��x{� y�37��9�B�������ƽ)L�u�bY'Y��;Ռ�+�L+˝����P��,A����Ꝡ��^#���'a����fı�J��0��Ȣ酄jQu�n�eX�;u4������3�5P�N��]��ͭ0�s i�n��hQ�v�8�8���='���:?L�fP<��ZsץMc�i���9�LC]���aP��kL?�6�TħU�%�j��u�/<�2�Gs�d�:{f�2�î��x�}�	.���-.�@p��������l[2Z�h2k[�E�򇅹U���m���e��|/��y[��铼|���:
���~�+_Vf�� ��V����q���')7���t�,l'���&}:��c��f��,ƌXgc=�8��p#�ۦ�m�fMb�^EV*��g��3۸ֆ��~���/�ŞA�&+���� /����pk�P�6ƃ�����V�C��xQe�j3\���a�������qhq2��[�Lq�c�hx�O��g\���X��n�= C>�05g�EX���P֝�4�/��5䮂<�@�z(S)j�{��|_oU���x�Q�j��N�[���r�K����:����8�դV�]I盳���hhu�/�]��WW^�7vNv�X�5���p"��.�K�*��1���nCW��n���䣬w6���ڶ'5Y��jy���>����i� �R~9�<JM���i�>\W?Þm�k�<X��KI
>>K�U>�z܋i��lo=	�� ��}M�
�9⭻�k���b�������{ڜO�4�<%�p8��Xt]��bUc�רz�v�;]�{�t����+$Jl&d�Z3I��^�通x/Mn�˙����%�7���Y��av�wmJ���A�uzd!^��淘!8�LK$�3L�ҕ&����^�ΞE=���Y��hީ0��sb�N����lJveB`�=� ��:���'��%:o.q,�2Z���X�a�K�T_UTT��n��R��P�o��$(��q�i���n�`��������-p1�Rp
�ԟ�ٽ��\<��5��Y��Z�� z3��#ϡ�x�#��Bm�1��F��Q{:�W�� ����S����bG��^�1F�X04����:�3LǠ?c�C�!��!�{Z���M�ꑨ�pW�As{��3}q�6օG���^���@�����xQ����B��h���i#�Q�5���'c7�]f��"�v`Kd�5�t��i�oV�}5R2���}z>�鼉��ӟ�����������z��ׯ^�=<x���x����y�u���.��wZ��ǫ��n��a������v������6��,��B,���Mκ=,�	p�h_sF��o���pXK��!��e^��{�BI�o�w+%�TG�ۚhFP����vv#\�!����1.�9
ҫAZX��R���p\�yuo;�d��j0�2Y�X���+].[�1���5�(2�X������{�5i0m�)z�U�[���9�y(ff<U1��OD\�o��#��e�R����B�t=�j��0d�6���껖���y�m�&輰Q��u�V�\'g^f� u�[v���T�mgkɱe�(�x*�Wf=F��;U\a"��^q�y��w*��)�k3.bvg0�m��}��*7ShS�֮��&(��]۶��g�y��;eon�oaQ�jZ�u��U2{U	����aH`���0�
hYv���ns�C2�l��#y�v���dv�����T��,х���H��b�);uF�`��9#5V�I.�)
���+T�'��/8���6��ʺ�b�Sz]uށE��-ݽŮ�B��ཀ�=VdK{.>1�iY���]�/I&>����X/xk�3SYT
	L���*d�a����}g�a��<vչ���ng�6)h�\f�����γ>�*ٳ8q�����[���	yB�	u6L#-��&��-���!��c�j��Q��7��+�Dt�`��rvK��vw u��=����&s}�!j�N�D�'��[\������uˤtĕ?
Y�`<ykG~ӆ���U����J��W9n�s�{p��L�a�V3M�Ɛ��V�F<��I6!�úQ��_d����a�Do6Y7f��:$�Rvp��cr��:�O(��Z�կ���S�OI���x�����%�-�	^d�s��nѹQ��l6��P�ۤ��֝�S(uU_g1Vj�Z5����6���b�zM֥4�ߝ�X{�Tǧ�2�I��G�]h���ܼpm�z�n�Cp���G[�xH�a�ݱF�Σ������b:5�s���(��S�&ҽט�+���o�F/yPn�%�j��[z:�����p�OEI;�.$��9��S�M)[ǎ6��a��R���y��ܓ*�W=�N�-�-�}�(`�.e)r�m��=�{+:1�*S���
�UxT�iNf���V��a��9���%P���Fd�o{���R�C3��	����%s*Ӆ&�j�/��Dy~�Y�fR{\wr���:��
�nL㧲����
u�����p�${]����ec1]��a&�[2޽��)�Y �jD��ܤw}��Ӡ����:��7'ùn�/ Hby*�{8w-�kM寛t;&s��쫉�qq����� kY�i�r���>uxhX�G/\\�C����t�����s�ùX����]�c���U�B ����͉9����"v�lf�r[��QT�����s8+��K�O6&('s�%�jl�-�g������NEb̜���-1s���cm4\���\��9<���*���������*�:�q�"c�71���)�,�ѹ�cL�q�l1���4ہ�Q`�p��c���Ztr�sY�\�ݏA��mR6koX��ĶW3�9�b�BI���Fw�	�PV�h�ϩ�r��n/ �#s<���b�12�Ŧ���6��1S�M�c�yrZ�b�Q�湓��69�D�&��9r��NTUQ��G��Z�\��[��T��Y#�ç��f$�L�':��Ep#Ss��A9�

0X��m9��j�lD��s�P\�Új���s��I��\�Ʈs�Ö��y�n<��X�i�lQZ�Csk��Ll�jy`��8ڢ&�1�F�
 ��'�SK���Vح�bTl�i���P�cj�#���Q�˦�(���9�UDZ4Th����<و�����������1[:J��b�����7�����()��U0I@G,U�7�b��`����|����B1Re���IQ2@]5{.��ޞ�
�P�O�����n��<בtI�=s�w�,Vи����3~Y����s!l��LY��٧�A�⼝))��0�H��T'͉8�Q(�eT)��� P����3���>m�����>��>F�ZEV�
Tg�]���|���?-[��nr/���heQ�����-�{��oއd�=	vO�z�Y��,:���̹�%���
��|_�?��C�7�v;sg
�KY�����q����40�s0����rڞ��>H�T{d���i�ps|LW0	-��\b�Ф֪~��Z5���v5�<�&v����h�X���#Y+���tP=��i�.��蛸�nR�١�������YQ��
���S���xT6DI��A�4[�|��uM��k��=a�
>�V,�{����̆���6��l�Q&]����/����H�|�PB1�=Ų.x�hP�V1�؝�=�w{5{���cbt���l�Z�W(5$gh�x��ǁQ�tx�6����ΊZy�^4����݁Yp9/L".��r�-mZa��0�J��ʂF���F;��[�S���(�1������������89�cOQ�oM ~4��ʂ�����b��FD�*�
`%����.,j���=6�t�/UE��g����"�a'�nK�	�d���L��s�7��8�Ȧ%VK*]��haRkS��GN0�Od���� ��ƀ���~�6�<�.�߫������MM��,7��[��DR/�����W���/J��n�'�"�;����-2^Q�Nb��DbSl3�['����vʾ��Dw4_M�\�x�W���Z�}F�M��o%��y���.��gQ���Ϟy�<<����EB�X� V� "P
Be��|}sF!Mn�l�n?x7H��&���3��|���4�r<#�!�BsS �p9B�V���_Z�z���%�k��v�"�BZ��5>Y~�I옦I�09���\>�N���
��!��_�������Ʋ"w��o�X��^K�e�5#��M���-@��OW�Ƒچ��nC���l�̶
�o;Qt���:6�>�H�	�=	y�5�B͘��.�TaK:y�_���P/���p+�=LU�syɜ�{�[wͦۻV8z`���,�0r�y�'�905�pυ-$���<�����'��5c́���]|f�;�`���r���9��Wᯈ�,�~h����ڕ���j��e�L��$�ce�������Tן��@��3�����h��#m���t޸�(��OW2�޶�]��f�=:�bK�&��f]�l��l��k˼ `L�����L�����x��*���۫���?�"��tC�Q��O#.�tE��tM�V�H#Һ��jY��_Q�~�ϴr�p��&3$�ت�Ƕ�{m̀|��U�B��^7�������y�����z�O1�r����Uu4U�jF���#���*�p�v�F#�e�q�������w�BV�;%������.������GHF~R���zQYB�U<K�{Z(�	s=b���@�)��g�:��L;��Mq�6��],����@�營;�܀
E(& 
Ji�B�hT�(ThA� �Za�!�o37���v�R��0�9���Dk��E�Ÿ���TcWX��kmJ��0�+U"S��eh|�(�sR�U{��ٽ�U��=>�D�Ӧ���E?p_3��i�9�أ+��nj��M��o9i�r���p�
��{nȦ�	�%�z{���,�VQ��ѯz�x��o�cϣ�#��aO��U>��Xw��;�S7{���%8
�RX&t���#g1����	���C�h:A�ŗ7ok�����v�5l+���_�[MH8k���)�1,���m��%I�s�8��s��_Xe���K�GdmZ�XpZf��xb�cO���>�.�Z5(���X��y��S� �a{�彈6:��aC2g/�nn���
7㴡�S��&�ɹ�}b�1Ԥ6��]Ma]���s��>���������1��6t�Oo�ė]0X�;B��ˀ�gYq~l�x
k��{�v�Ǳ��H��di	���^�1�z_�y~h/�uz8s��~>�=?LĨ���t�L��ҶbR��r^�ʸ�A��m�t[�����?�v�L��>�*#�3V6F�\ٽGn;+����T���ML<KV�2WZ�^9�4�\���{�8�B�;i殬����.+�ZJ�Ē�dT遽m��z��y�o]�j&���&e�VC�7*���n� �����kT�s���9o��>9�����}�`B�I�D)I�eD�%D�E&B�e�J J���RHT�ZPg��߾���x�*��e?ۙ6���I����l���׉�i=r�k�,3����぀��Í�Z*){�i�w;wB�s�銗X��v���d�loN�$�`�zK׸������-]b�x�������n�Q�{��uݙd�!�Z��I�O~ڌ�K4��W��5�C���Ӱ�y��dο����w�ޛ�`�'���T1��3�2L=�OC��9��|Mi��u3�X����{��4�	�q�&0��Z)��U�ZfP��	�ѯP��`yNo�R=<�7"���	��ƪ����z���ru3j�(2�Z�`��H���ϖI��D�<�� >���>^��w�2ڮ$�V�l�]�Ϗ�.�
�qBLW�Z"y��FPd��Y�V�E��z3�lz�Kϭ���o]h�;-SXo]VwwXR�ע��4�vAk���≉d�� �2�J�]�����P�Ӏ���Z�WYX�joOv�t8(
A�.��ۨ�G` ���A�%:O�bS��S&��������'�V�q�nV,dEê@P-�
�m�Lpe=��
�$É�i'��)������>%l�뺥�����t�v������y�V���I� ��D4@ɴ�J�g��[�Tԏ|�n0d���@�ā���XuB����<Fư�升��AO��yں]Mė�@����U�R�*.V��Mq�l	���ܽ�Rń��J��>>O_t� R(A �*C#@�1@E�(H- @�H)$ҠL 0G�<>������C�_����o^�[2ݷ��_e�H;_rB�أ���ǽC�W�����}�4[��=Ȅ�Bc�l��=/E�S.tNnU�\D_��=�a��u�-? ����Z�f�I��E�2�F��G8���\)�8$Z�Sy���vwJ����3�w岋��4�}��U�$:~y�l�zQC|{��m�qܤE�;����-�iS>��`K,=X�~��2m�ǕύLO�,;D�<��[b��+��g�^bƪ�3S>�=�K~�vlp9>K��^��Ė@�k-{����W4���I��h79R���PY����K�<k0Я���}^���e��W���=�Rpl'3L8����9�\T/��6j�ɝ�N���,"�@��?��rP�4kr�߶�k �P~ypІ�a��=�X��]v�.�j�mi�w���\���Xi|D�o�q����:��-�r^��e$zbg���>WܨE�]�)���˵�5'��6�v��&`�UH�o�ww1�T����i�+���T�n�UȖ�mcbr���l�Y*�R3���l� [:y�p����l#��Q�hg�XCSk�V'��W�����e���U��ۃ�f}i��3BX�6���L��;�MΘ��A�������1���Ywc���t���`�uj��ߺȯt
*�F���Ŝ�m�|�ڬ�aʬ�e�}�Nu	c��/��VF�YaQ��(I(&)@�
 ��JI��o{��`���Q�S��+�q�K�>c�
7#��2"�<4�	��� �ӈe��z���孕C)֣��Σ�Ҳ�9�V���a��e����i��_r�?B���^#B����|S��r�`{��K��dv8VÙ���z�4�ςD&��Ⱥ�I�}�.�$vJnj~��8�7�ҙ
.3)�u����Sk��R�j�*�qvt�	�d[CyP���`O�[%�!�e;r�����YS�P�W�Q}J���3{mC+4i2�0:�K�G��^��[�	܀��bϙG7��*�v�����-ww! �c�b���ʒ���d\��摈����>���3�ˇ�\޲�~3���W�j�������/<�]J�i0����)=X	Ic^GjJxw����dmEd����L�]8|k��L@-���^u�u�`��.�%P�,��Ua]kx+���Z�Mf��zѷ�Ƨ��3�֯u0�ni�a6C�ka�L��y�X�W8 _�����
�^*��]�[e�]bi�V�@���(~��0����'월[�X�z=�*��1M � :i��]:��cEx��O����aڣU�:GB���R�L��*��?���	9�ܫ'�}�UP��꫸��R����fR���=������'VpFb�[{QwLͽ���n�!<۽��q���������9�G��������� �Z�D(X�Z� !R�!�B��Y����~o��}�����[E���������њMKsP�az/a�ό�w��0"��x����`�93���Ukgf�g&`/}���f�:�e&�bK�&�� L˴�ly�3��yw���-���a<�Q��Ż�[�F9`���j�a�2}6�lwH$8�P�<���c>��:'=�,[�\�ģ"-c�y�fK�N� ́g���Qw�S���U�m���o�<1���*�!C��������d��y�{�_Tlc��L\9�{��S�w4^���j�ɟK�jP�΄7�qqs>ͨ�cҷjֽ�,��^˕v�z^^7�,H��{X�3����0��~x~���<@���
�_�·9����Un�\�f�9oY0&�J9B�׺�_Zm�S�;�� b�|�J}���9�=f�&fz�d�gwPd+���	LAp!:�%%�gJ<�S�]��}Ǆ�o��!Ű�B0���sp�Z7��#�0�n[3�gU��L�!'
�wL$�C�K#���)��&��q,U(��{�i7a����73���;�}�Ja��K���"Q�P�h�.�#0���,l��kz���	ʋrn��;-�,�Vgî�Y�ol�Ѕ��+��ǵ�U#����w|f��n�t�'��=fE�V���9�S�)�n��?20�yu���5x.�,�uH)�t�2
w]f�v�N�"�{����5��ٶʖ�a妷�MYy�X�)��}�ZE&A%h@$�� $!R	D�"JTb
Q)�'��׾���������[��;���K��p͍1�u	���vl�)��t��i����MmF�W�5>������~�k\k�!c�����d$��^�ݳ]P5:ü^�Nׅ��E��:�&�Eu[�5wWc�C32�t9/JwU~��r��1��*��?|���#���|С�%�?��c��u��*��໦�;�6��G����zW=����W.G�N�;!t� ���~@}0�k�ٝ�ᢢ��՗O/�Ͷ�ِ-���Lm<u>��}���|z��ы�g���j����봰�(:���	�(a��S��
��g��w�}�;=V��g��,C	����Ea��Pk��9�7�6�ý�	��bL�e�^��>&�ݬ`�#�zRe4����>�K�ݣ��{���N��)��6"��8�΃�rC�w�'�Q����m�R���qm�R��b��P�v���#B��) ����R��eX\O��|?|D&c#)��z9���ќ���G'Ǭ��ӵ=ܭ���S6X�C��ԑ��z͙�b�O��4��,X_~@_�����.lޯc�����܄�ʾC���cJ�������f�x����s�u��xez����'�I:��/#,QZ�q�y�D����L�6
�צ���۶�0Q#2�WPk1�+2�7�S�W6۾v�9��_kw�J�_�|?r"f�H�ZQ�d�f��I�~�k����ˤZ�G&Y�5��ٝ�����N�pO�}&���دH<����2�&�h�'�F@�z3���׭����]��T��]#9������,���5l�(F*��A8�bY'���)��R�>{�:��ئѳ�f���T�&��˚)�=����yٲ�=� �7d�v��d��ħV�˗<���Y���K������\Y+J������m>���js���d;x,�$wQ��T�]M��:�w��\�:��Q���j����GPh���C� siW�Z��xN3]������m��2��ŧ匤�5&��İ����A'�KP����r�{��O�i=\��7�}{�4��WM2������]ॻi���nv7I�`����f�6V�.,Sv�h9%�������%Ї�ѡ2'���E7WOV5���2m�¹�x�H���ٴf6�"����W�����<E~��<�Y�g��4�H���$��u��e����z��QjQ���.����E����[B�}��� ��Ŧ[Ի'�p�}픟����7�������1"��Y�S`�e=o�w~�M��ۓ��Є�lwG����ƺ�T�	�5�k�d��1	��J2���\9v�v������"�˟�|�/���ѯ� �	u��u�˲�wx�^����f����������x~
�H�H�0�RH*�R$J	0	A� �_Q�J���;�V��1�W��H?uy��>(��~6����O�f�����_Sa�^/V���u�8�!jk���b����tE��sͼ�ȗt��O��
�uvvD"�U�����ӭ�����e���K�QM�A�B2�m�I�a���dS��"[��nw*����A�9�=�o��q{��#$U�A�_�,��J@�|ض� [:u���gXB{-�_vwa�u� ϴB�C�=0����U�{T�Z��'��hH�3�j
5�KU=M0�
y��]�Ъ=��;jy�Ӷ��'��U�B��#�4�h<sW�� �ɊN�X���u��5v��ޥ�lu&��5�8��g�.q����(2.� \�#r]�vBndzw�]!6��r��ӵ���7���Ө��ci�ҩ'~��a��г���1�C�;�o#�Ir�0��~������~ڃ}\f|�*L��`&*ۤRz"h������}�����Tb����6�8ǴǇy��ʻCH�)蘦E�c�}����zk���3�����=��/w���_��������|z�^�z��ǏY�-@�0�����;׭a8�w$zU���;#4���^�7��|����o~�eY�TS0�x��6Kw�F�/hRӈ+�
?O;Q�ǜ�l˦-�q�sk��Xh���IitC+���)���l.�v��[�Qn��:އ�3q���Z������L�o����v�A��<��;\	^avG&�$�!1�3��u\�ݬ�
UG.�gI����/z�����o7��
ic���eb��{�u�nf�7������.���n�ӍZ>v988��x/9µB�Q�]�.=lG��(� T7WZ���D�hj_pdo]u7������� 
��S/��Z��#-pE�2�fj;SUL��x㛸�Rc��"櫌��ɥ��[�rk���0 �!e7��;rb�*���鼾c.�|N.H���sѵ����n��(c�\��s�Y��q����j�v�S����X-2Uvb��
͕:c�U����J��h��ˋ�U�jAw�u=#J|�x��'���M����b�u���\������&�e��*�{D��o����y\|3)s|U�QN���Tz���Sb�orP{��3{q��zh�a��r�C_���b�f^�@t�&��)f-�Z�Y��ZF:�0\l0��3�챡�Ǵ6CX��-{%�*�gMm(u �Lc��PsKv��:�V��d��4�^�n#']Z��8���b�5��C�p&�ӛ7��n�Z{lⷋ���n�I�¨M=$��
��zC�Gl	9c���{]�$��������F�Xk	P��q�7Z���@s�	V"����HQ����h)*u�V�����*�F���(|*����;[�`i��x�H�s#�xV�a�=ζ}�z�jv�LEºuw;ah�1�*J�(QY�a.���|���A>�z�hێ�ȍG�#SOn��:�����l����:}]�K��RI3�`l^��D����b�.f�ᨓG�7�JgW#yK,O��*�l��Tr��^����+�*��v���G�e�M�4἗�W!=/7{����ŋ2�x9�+t��M>�U\7Ù�9j.t��`;���N��Q�q&a�s���d`ʤ�<75���9,�44��tnR��U���Y�
����Uq�RiG���_}}�_�Pٕj��6Kq�vJ�)��Zܶ�����n;R��z�VaN����H�Vޭ�:�}�,E�����ڱem��6_nth#h�C�p��,�Q�}���1uƾ���(܂��G�$J�crHҲpN�����y�/u�/o�*�k�3T˕��dOGo���5ɲ0��nƚZ3J�پ[W�nSj.Xop�۰I�C�	�s�Ւ�Vd�v���,p9�_�U,��kܼ��P�5
�%����^��x�+�n�Ղ��i7Ũ����;y�8ܨi�u����*�7���ͳ�@���;�W�G?\޾~=�s��t�i)���+���R��bu��-��)�j
((4j�"���cˉAM�t�MDS��C�i"��I�(�c��j���J@�������j4bY��P��)��&
j���ܱE0LDI�530QAO1��b����
""�)$��l�SDMTـ�
j��lSZ5TULm��"��EDTW�瑉��eđS���T��%��"����H��I3z�T�SPSIEEUQ�t:i*��J�����h֨"	���&�
����h-f�!�����)���$��*�"�#m�芩��*���Sl��)4��Z�h��"Z���1DU4Um��* �J�
�"��M�Qƪ�lTVڙ�t�b�SQ4�0cY��U%$DQQUSUSh�R��i0|\㤊#k��h��h#X)-�%Q��h6�z}3�.���������:g�44�2��L�	=Y�43�-Z��;R�ޙ:�:��G�Ti9|�W�N�7j������1�B#���|?�����=�x]f�	�&�wfu-���טpm/R�_�L�:�aTrW<��I����4��0�SR��ի���v-w���ÖO�:n�qz����4,ߌI�`�E�ΎeAM��cJa�מ�s#�8�s>�� ��m�B�>���Jp]1�Ll��hZ/v��=ws���?u�j��YN��9=��Ts	 ��Z�XK�3�Fy�I/Ý|�dd����Wu��=�0c��o�;2�˩ӿMkϸð��71�\���L߁p�4Ba���(���CX����ھ�3�P�f\��3n�ܢ�	�/G���{�_{h���RǂЀ5�29�k�.�ƻr���!�^�<��6nq�g����'v0�Y�	EG�<��O���A����'���s�է1��ͣ\My	�q1�)=�@�mcv1�����G9*�!�w����)W��q��rw7C����;k���?��,:N$��/uQ�]~��]65�JB�ɵO�\5[nn�U�V�1Z���4u�׷�	q�_�B��g@��A�������������ߓ���pV���=+��hX�ڒ��ݜ��QMn��2��.�}	=Ȏ&)�B�_c�
������h�5��T��B�
��h�y���S����S��1��\�rwCp�.n�t}��sB�.�&�x�'��:i�1��V]�6�Oc]��_��{��{��0` ���8�:����X��� ���&BeBѮ�i�R[Bь��z���{gh3��3�ƴ�K�^t�(��S�O�+c<��;׽܄�myY^3͡�ϙ�+�yՄ��y�X���GNc�m�s�[���E�=�[|}/[���xu:^�~s�v k��	:��%�t9��*�8�ph���W���t�;_�K�`���X|�!�{D��a�K��jQu��)�z�s��f�pD��g�7�s;�# u?/=�p���{d�k_����7O�
6҇Gtza�SR�AT��z�h�wvb5�/b�eK�C�>B$�X[<~���|�i�_g����n6��o���{�]�]u$U��.�Gs��t9�̟���8~�B�:CC0�����;4���(՘��WUc[+o�����(����O~W�|��Nl�{�h�F�z��f罹o1Q�;��f����;3m:fn���M&)���I��עc��C1�����c���o�\�wj˄�x�|!�|Ob]���O�6nB/�Ǥ�- �<|�9�<��O�7!���q4u���o��"�u���4{"�]�콰ƴ���s�5Z�����u���ʫ��/���q��,Ɓ�6+wvǤ���NJ6��U��]C^�g[�;C���nv��Έaw; �;W[@5H�q�^�&���{X��#����| ��R�����-������-�p"&��F���؇nO���x@��\H*l����t��h9�n�0v�;��񳫲(��et�!�f;[|��kX�^P|�Idz�`V=C�m��>�D�����g=�CY��9�۝sx����S��ܝLЅ�Lt��K�{cR~h���1a�|>��/�F�慯�
quƜ���^���LI2�ha�cC֦�&�����@ǫxU�)��V��C1�0k�����������R��(ן`�"Se�eMV�z�>Wz�ۼ*�f�h��Nk��q�'�z�On�w�\rD����4��w�N(��I�$f�X�&�&�0��=��4u��F�U�L�Ǣ��=��6I�.͔#ŅW�̘Tu��$vI���>y�Ju�'s�Lc�`�9ݙ-��syb����I`��= ��t��vc�.�vo2��0�����{ģ����5�Rw��~��^�.�a�@׌�v����a#��~�!�_?^�5q�,�s}���g�����LZ~XH%�ړH�Fi�������C�����}���Lk����y��JU�o���&�̥���y�Ŭ0���mT��Ï��Dw)w
.��v�i��fo��l`�8���^��Y�*�f ��d����T����VZt�]je�ٻE�c܎���pu��Y���%�e5�2����NC\2.C��� '����l��)ó����W�k�;��H�R�
��M��Ļ�����4��u�ۺ*/Z;�ht5y��<����s�E77�t��_t$��-2m�T{T�M�p�����ڹv�-������viC!�8��'�v�E�	vokd��B���è�e�h�����61"�.�w_B;*����*�~��VX^�� �AA�7��#����AZ�x� ���ۼ��}
���ȗo�脤8�x�r��,C��<4@~g��Р��&9ف��l _j.韓+�����Uf� ��	�@���D�1i`��D_x�F����P���X
��[��E��f���ߓ��Q�7D��
��7�}_*�vO����$�QSl�r0��֟�h���"����:�;��h�#�h~a�-�=����m>�	�P��W(5��={6q���X�0<;��w7֨��w!l�}��To`eϐ��L+�7!r*�=~�$'����qz����3�G�rg���v�U�}ذ�
�3�Q�v���v�S������X�7����1���阬h�;j5l;k=��*�鞹0�sk*�/g�޳j�@�d���f-�.�sSc�Kc�k�8f6��P5�W
Ȭ|,m��[gVt:��R]��Pmf외3��ADj���JHେ�n�J�nٝE�}p��ur�Sa⩌�'���> �j��WI��q�;��*�Ja,��ۇT\:�q�牡�
�\���nK��l�m��]�u��Z�0Y'�1)Մ�W*�qw8�{"��oD��!�2�����Dd�Bz�YW�}���.�0�a�wQ����g��Rz	@����Ob\n8�W�h<���pవ�>��} ��.!�v��)�I�`u�`sN"�4�O?D�љ)n�_���﷦��MO�-,`C�<re���4(ߎ�aTrW<�x�[$�iIc�����oㅥ~[�t������,/�0f�ק�|ŋ����ю�Q�f�I�`�@��D�q�ۻZq� 6눟���C����(�i�B��0�צ�LO�W�I5���Umm^��v��n��훷�(u+��PK�Z��O~�Mr��N�L�b@�J�)񁄿$���<��oa��\ͷӴdB�;FfN7�2:Ui�k^�v��j[���t�/e�3�"D���`9a��?_Q��)�ǥ��~/��3~o �y��(^�3�v:�$��j���\S9p;����;���~�(~t�t�+sMpj��;la�HD�7�βV��׽6�9�
�.�ftQ=��\��@! ��!�`��X�s���l���8�*�޾���Ւ��-��y+���S9�0�wv��|\�5��
�<�W�����xi������"�������P��ݿ�����6!�%����19�L�dYx�H~@A�vI��y�.��'S�a 9�<[�e�lVb@?���O�@X�w�ׇ͍1{�������M{�T=�}w�t����~~���\^�R�����`!~�bä�sE�1��NT��Uh:yaV�/��|zo�m�]nR��(A�[�kT���a��*PئxB�8&IxXQ�wt{C$��~O}���\��Zd��)��	�.�%ԣ�.�N��=[�M=���[^c�;�]��񛮫��#����zw�a�j~BS���%�L����F�c׵��`�����wZN��N�s/s�*`p/#���g��	9@1�d�`��oS��%����nᲷ:�ۀQ�p�G��={gѭ4z�G��R���@��&�dQt��5(�P� �'ۛ�r���7��د#��6���W��^� ��}!7P�	�Ga�F��P⪰�7\��᫺�m��Ku�K�Qi�s�PX�]* \k�!cݬ-��@B���zz�Itޟ/?�[\�bf���q�n�swz�B�Ƭ�gx�l�`��|��Q��a����k�oA�c�jC�=�!�)Գuvet�.����8�j}\+�u�4�!���{m��c��keޡ ������k�EX��&�՝�7M=Vf�,ӫ�_E*��C�xxZ&�r�u��uWf�ѿ[��H� ��L�D[}4v��EQ��,��Ua]��s�`[H�����_	�%��燘�^yVu�{+V���^Pٔg��2���	�\��^��+�<�w,��L�d0`;fh(�̌D�5w����Zϝ�C���#m���H�f�y�Xm���Ll'���cя������1�4�3-X�̞��ί���c�_Uv�P�p��xA.��_%�>�d�l��E��Ǥ�- �}[-p��T��\MN_K�D����Aݵt.�r�Cap���f�X��η�����+�t���{�����~�@.l��S���n=����ωل<��k�����/͂�{��r��\�wl�w*f��,%t�R]x)��..�65(������|r\Ͽ�����d/�Owj�؟����{i��C3�V`���QLo�1�"3`򡊭?����fM,��}�²���t�W�{��b��/T�����^��%6_��5Z3I�J2 Fc���lg1{�]����ǂ�s�x$)����!Ő��ju��!*��=�#4ɼ�^o�Wُ��{b�3w.��a�NC�*v�E9�O;��z6Yb�GS�
��+���]ի6\(�~�������W�1�^�Q��צ��Ih�.�GV�,�<�*��vwjsEJl��s�٦�j۹��ִ�Ȇ<tU��җ>y}l�
j�3���>�G&�OA��쟵��7�휼�{w�
J�.͐��v4�'ݒy��%=.�R�W%�`��+o�ɾ�6�	nIO�&��d�Ac���9�1��~P	�Нk��7%�'�����S ۧ:�i�;�e�ʣI>1I�S���J`Z��jz����E��pB=Ȅۜi����d�j�=�ʽ!��T����L4�rt���Px�"�4�K@~�y��I�%��ݱ����2���L<6��Қn�v��;(����@r�����8�;�f�n���t�8�Rvv�@�'���P����N$St��k�wJNZ֙6�a\�3Ř�uA�,��778oG6�f�)lc�7k�jA���]ٵ�|��k��BՀbK�^5��D[�k֑Bn���*j���^���Zɺ���;�c�m��tŝ���˲|�n^h���97h����oު��zࡎ��½ɠQ3<����-E�;��x��сAi���G���yy�-{���F6��Rx*ovC�hEd
.�L�Zx�w���9����{A�4�����9٧_B)�`�=�/sɌy��egӌ�szsX�]�^�V%u�"���"�ZtFv뷕ȡRf:�N����SwS���4.sTr5��3Y�ئ��1Sgq�B[I��1�S�����2�}-%�r���k]^�߸��t��+��������J����������͆ff��1������u��Fe�C�@%ڼT� ��F]����9���b�Q��i��w��w�!�C�[o=�\���kFH?�z� ũ+��Fu��MB��sY.����ޝ��b�@�h+Ʊe~�3�t�U�E����@5A	��?�6���N�_k�b��B�V��g���C*.U�fA8�"Kϼ�/<�^�X�#!s�sh=�Q/%i�ε���Q���塣�r���FD�RXK �'����q��"z Pd\:NKK�eI���u�+7��PU�Y59��=�1)Մ�V�IŽ{��`�hUӍ�񣱜����1x��yu���C�Cd��dw:a���&X�LU�H�>���w��,6����qᄮؠ��Y(�U/3��x������B�8@��r<%��a�i�)蘦E��I����-j���5Sw<S	�A�7�{3��N��?;3����������=�hQ���Q�s����JON2�B{ۉ��RUV�x&�yC
چ<���=�����t����ץ�]WQ�w�h���w�������g��w���v��s��HJ��r`H��w��RD��ǎQ�k�24&q�A���i�N[/��}�gEՀ�z�b��N��Ņnqc/��zb���}v�H!�������Mm���=Cl��I�d��.�
�_���[��+�%���WJcV�XH/v��=�x��}n�ks_�U�2�Z\��jS5�������#u{bN��Oҹ�(%�ʮP��n�<+�S%�
5�̯5�k8u�R��Ko8�;[fgONaٺ�YI��v�@��}�ӴMKsq�b�g&;�ʆI�$��W�ک�?v�	!���![�;7s��Ͳ;r�^���L3z̻O���2:�͞�v[/���T��rϮ�<���HF'�����NN�Y�S�q��;���m�k����f{���I7ƿ��~�y�����3>P{.23%'�z��h݌i�d�)LD��5��N:��1�2�]�)^in��=S��Y�X@�踟���}]�c���K��v��ߺ|��� �f�2�Z���Q�[ӌ}�{g����ҩ>����,�L�j��'V�p9uy�\�Ks���D���L�ѡI�J9B���{��
{glI�s�[�;%����Ǎ㽂ֶ���	�H$Q����ٞU�`<�)��1)Մ��MBT.�l�:��g�����=|~����������������O_^����p�gK�p(��Qg����c� ����c����£�t5��:��E;�B���A1t����a��h�-�n��49�^N�cxG3���-�S6�r�o)gXu�2��&Y:�Y�������ڪƽR̰D���tVAю��Gj� �]�V�������w�ڸ�}�q9T�pz��-C
5��~%�3�����'Sia�&Gl�;�yL3A������F���r,gt����L�3�NYÔ�ȃ���T��Y�e��*�]���3�f� ̶��x̭�\�k;�����!w&.��ٱ[��UtjvY��iA���Xl�jB$!d�*�MO�2�}n����.T���ԏ�W���*�T��-���f@�\6�,��p��m:-���aH-�wx�����'��sE��/(wK����9I)	p��-Eq�ڋ8�
m�f�/�Mֶ&f��y[Ů��Du�Kw`�SՇN��@O��8���k3ӵY)�Ӈkx(\[L��E�(QN��o	N�)�{
f�ˊ�r���!���p+#�l���$�f�#lp��Zsj���������w}(������Y{Ǝ:���V�fK4nc��U�6���ȧ,�grҺ���n#G��9�DYs����f8�>�sm��p {����L�"� �w3����$/F��k�65���s�6�u��Z�@l˴D�����G�f�{o��Rn�v���Y�����69H/A���}��0��:�R���t��^h&�<_��c�u{��p��q��h�;:���<W"�u]�t�/��o*�-��UX��}���3i+�x ]�>�����t�/:s���fO�=����/G��3.ߙ���1�ڗɩ���p<`Z7�s������lg4T�Y��
Z�!�*��]�sSj�m���i��1:房��K�#�m�gjy�qa��S���Vd�7P����;Z&�[��±	K��L�vF������0�ydL��]}c�r79 bGv��6�W]���-޹sNq��wl�t�ۻkGoF�jɼW&3��U�[c[4���"fb��x��@e���dD~�����N,�щ���tΩ���zOL���6'/n�tɷ(��;�t�x1���V�
%��.�;��"��an,P�x8��XGjs�4j��;�l�gWR��<�`��Ɖ�|�iQ�ԝW�c[�U�T�}�w�ͷ���PsѲؤ.b��p�9�b.�∾B�RoZo�J�vb�L��)fn��/*l 7�w^�|��^jlia��q�y׬>]�Ǉ|�^��Q�3M��5�{Y�J�8���<cicՁ�:�sX�)4�{:�f��zwZ���Ny��YY/2��ft�룝���՜]�t����b�jd��tz��1���Z6$.!�Y%_3���1�9�||3TEAE�4;cTj��)"t��8������	��
)��LT���)IAN�QEKDIE5Z�إ���}N�hJ��e�h��F���ccZ5T!�h�EV�b5���,T�kZ�E1U6�
����t��I�t�SQLU)ST���uDM%$�$US5LAA�CA��*��kQb��m��������"b��"�ƹ������"���4�1T��B�
��F�"�(nYh�%��)5�h(���&m8�
�(���+C���(��-�MTA}mAL�`�gjMR�SUM5QPTE4kA�T֜N�mM4��UT�EUV�b-h�*h����� )t�#AcQESUUA:�P�M3DQI5-44�m�b)*��X�~���\���#3	
8�d"\a���Q�� ��NG��߯��k�S(�n��'[�KNi�n�,!e%rP�����x�z'}q�u*E�E��;Q.��7�bx	ck\!�"4\E�R�6���lG���0SF)2QFҁ�$�"L�J!4��  p�f�_UK���W.{�ԔB� g��Q�����SƝ�*��@�hv�wL��<ĲN�<��M�=��Iߌ���J�.����e��.�CT�]���w�LV��o��W�t�,��]r���.WV?fg.��W�i�S*Zj�4�Ϡ?<�{d-ٱ�GM�逛��Т��t������;��{خ}0Y4��='���4J�����-�������==���{��U�lC�n��b������5?.�,Rմ.�*��ydw:�
�w=,��>/NqÊB5�f���L*kh���Ň�`��>'4&�4Ǧg���Z�����z���>� ��6���|˦g�j�-n�V�~��#	���R'�h��_K?X*�	��ɟN�/�Sk��c�t�c.����{������s�Q���0��4]�5��.���d3n������]P�혣�f����8�k�8t�y3	��F[ }�!��z��������f�X8�rl�9B�l5mz��n;�VڦʔŜ���i/��ӱ�2%����c��{d�����tΥ%�i��#��p�e9%ԙ]��D6��
���K�8q�׼���O���6��о7�������q[����t>�ӕ̼����YV6mS0�.ll�[j���4�gpe�k`�x�7	���i6����u[͍NT9�X�����I��9���^�u�~�CZw@�L�W�X+��r���)>sͼ4�^Y�?45=u��V}�Nƞ���P`���O�_q�iJ�� ƔS���{Ȳ���%�\�����i뻰����8-íy�\zT�	p���q�Ʉ��f�ߥ�Xe35�y?��˧nS�M<k�|w����ߢ!�V�"�b�j�� ���;!ϛ6O!%���d�6���z�𻈪�Q�ڷ{�%D�f�t�gcH"{$��60樈Ӭ����X��ڛ}�A�Jsat��w�T����_"��?��m"�m����e+k{���n��ѭ7�C3)as��� �u$���

����a����={'ѡ񅠄zL9��˾��[�}����\>���-I��c����LZ~Y�R	z�
���0����b3V}���i_]��1O�{Gȍ��k��r!�^��M7_j�k��/5�5���@'�q٪�b���������m��k�}q�;��}>`�sȇb�bk���M��Ս}Г��ɷ��y��&��_�S�O�P��9ؕd65�k��~����_zV��3�>v��w��	�=�%26��o��q�Q�Z�Y-o*�ۋ/����'6���lM�]2��S�]RnH�����:�&���\ۥW����U��ȶEX�w ���m��� ��)=��o(���T����0M��c#��pna ���ͮ���_'צ��1%��i�[DdN�N=�����l�@j������~]az��鬃��S���[�2w��)���qM�9�o;��ŽH�7���0�- ��[��m/`�p�b�����^��o.o~�(�ҷ��N9[Rcz����5>i�f˵,���0]ĝe�s͟D�l�wa��Y�W��G>��u"c#�����L?�u�N6����xfY���%ب�A�t;[�Zw�g�|\����k�wN�ǎ��2�a y�-�{W>���Ƒ�*� Ũ%r�3�"k�m�g%_o�$�u��U�Fѿ��x��� B�~9����&�9m��O�v�_Ubs�	�D���4v�X/��7/"k��;�������("�Iq�����S�����j蓹�/3����o,�A���LRuc�J�ڻ'�Ầ���g�Xz�"�#�W�U3]j4��q�I�Y���d�s79d���%:��P�'��� �v_����y{/�ݨ9��Z2�%��[*��ڵZ��qhm»�[ѵr�YtN���#���Ogr�bQ{Ph�j���hl�!s�Îܸ��w$�G�n����ݜp^��q���M�t,���ڔ����;�ȹv˺���9
��6�*�Z]�9U�w(��?h�o�� 60���l_ɾ���>���.�FgL4�Q>�ρ��_��Rt���&�s�Yl��	4�1���]�u��l_�w�֟C�\И9�v@�]�a��T�z@��E�1���γ��jY���b�8wv�y�J	M�;�?<���@A�בCw=K�x(�F�i0����IܗK�ZL7v�N�vc�/K>�~���D�ɤ�X��X���=	��	y�U�B�VyH�Ѧ��TR��[j��Y2X/,��s�ŕ�%=��P/h&5
�-=$=<i��������2������Uz���ٔ,ߌI�`�J�%����`z�ksPw��p�3&uY���qzJ������զre��?Y�X=�n]SX�Aֈ�������f���<E�u<�����k<xJ��P��n�y�N��wj�T�bx�n�L3$�v�@�>�v�bK�&��x��j�d=tV��=o~����*����K��QJQ'���=����a���`�u� /�	�*jV�M�����82�˴�G�N1�bqᲽ���(=�d��uN�Y�n�4<����G�_�v}��$W��#Tr����ˠ�ݕ�{��s+<ȍAv+�lv���Y�-�;p�^���d�"��+amv�qִC�匦�s�ɉ�S�r$9�r�k�N�-睔ש��f�ݵ�cb]t�T�B��|���������d���kS�f'��IOZ�*��}�{*�!E�^��7C�:ז~��zúP E��t#Wn;l��{�ƃ�cv���!�m�Ɇ�I $-{aUj�R��p��l3�1LkbY�M��j�o��2Z�̭1��ݖ�%BG<�q��s�-��~BV�!2�Z4)=�9B���ƚxf�[q���نSMW݊Y6��s�&�>!�v)��~B�^� �I`��	*����g�.)��R{�=�/ڇ�G�T� �;xw�F�ux[]>ѻ2K���,x���	Z��Լѣ-��{���z�
~���s���H0͎���r�ݍ"U{��=�=#"6�+s[2*�� ��x�>0T�S+m�c@�T2�@�NZ��mx�Ђ�lg��&�ҥ�����uy�U��t�Y{=%,U��r-?2NX�J���w�������M���������v�fm���mjbK�*�Ú���w�o��=����]o����di�zp��xl��=��+[����M�Qvѻ�B��ly�.u��)���&u��zV��`��{
�\�Kz<�idv��5h�5�j9�a��1�v/]Ƣ��b��!:�Y(��סXśu���8��v+��{K�k�W]	.nW�&���+��ګ�5�[�L���ɻ25�щ�Zr���=�Y�q�l�۪����<}Pm�wٽ%n^�p����P��7�����~�\���>2"P�^a�4�vm��e��.�)��x�}&=���3��-R�'o0ꚼ�E���9�3E��+�1��h�^D<��{�dfHf�ܔ_�xŔ�ք�{��[����恻H�z|tE�j��y�ސr�=���`9�)����T�?,��\�l+L{��{�+�J�2�z�xO{z���',ȯ�!���,o�Ժ)��ED��׽�a����^���Cl�h��,��9I��WI�Q��Yްsuث!���|����B-��,��O�1�O��nEK5ل���	�7!�ٳ��۸F0��b&r�]ej�`�^J2)�88���ȋ�OB�`�N�zGq�/����h�'�YiF�zqgtgn�J��� Y�^<��>��
H��� "V�1#sS� �Y����H��X�ܵ==�fZˠ5)�W�J�n�om��ΞE=��.2��K�e	��H�iL�}gx��ɇ��5]����-�^s]'�9�N�ˤg����f��zyc���~L~b��:|��^�GM�:��r����Nvs�	��Aݑ�D��ͱ̫���Cjü���`D�K��(��v���[נ�����v�c�L�^Z�+v!ΪD��\�Ʃ:�|�%�j�V�c�X'��W���h�XM�o_"�[��8l�������=�٧A��na�?ާ`��L8��4�㘤�`n�J��,��Lg���}C�N�M�z�������p^O�uLpn��ME��i �&�r^��
s��H�bXV��[�0_����6��g�e>h�D��&v#�X��}z��������/ R��\��xy[j��_�����2�D�R���-&����C`t������L��TjE1�t�c]�INX��FX�g�Q�������X^���T�y���ٻ]�w�?0!����C�u�M=�9΄dq�䚨z������m[��2׿#���4�������GP�n��8k���Bd��؝���bS�Ѧ�����g;<�_s2C��v�N��v������[�>���H�>��0^Q�Ʃ�vꮎX򣻬��=��kə���f�krސ��w��f��0ͅ�q�����E<GSk-���Y-���!���C�h��	������u����e�^�]��dyv����*Tg>��)�6�]sͼe{o�.F�3�9���s�Uȯ3v��Zt��fb�w�����b�3.���9�ΰw��F����#�ޯ9�{��]WZ9�B��;�o�\������&�z�E�����yMVր.��k���r����QЎ���u	���e�ճ8�Bq���]M��[�x��iɸ�]���N�)5��O\N	a�� �p�gOov����ӥVl��{X���T���1z`�}�l�u�b�i��b�d"���з�ރ�s��}d1B	�Z�,�$j=�c��*.Ձ��
�x.29�b+��6�ۉ��63��gv�jd# �[�A����W:�F�+�0���'��ޘW�g�"-�5�pgD/1�׹
�t����L.v�r]���-�^~�ʼ���%:���j��GN0��Э�����1Ӷӻۦ��{��i�D8�����v���Θi�I�0~�mi���y�vsKC��4����Z�p�V�°���b�����^jg�3��%=Y3l���Њ~{���g�ڳ�������E�Z1%�~g�l����¤3~2a������7�M���4=@�˭�؊V7T�� 9\�=ZRXבچ>M ��Aö_���~U��|�Z^}��GMvwJ���◑TXP�:q���]i~WkMr��A���Ї��{2Z�")�c<�7�réiS^�����lI�bu.|J	{e/�?m��XK��>�//^bU��$��3�~���g�h�­ś��Xm�+]�Z���4���ó�s/2u�/QA8�r��2���7�5_d�Q2��]���U���ǖv:�����P��f��M�&mK�9[��y���T-m޶[X/��K1@��[�u���c��vq��=Ey���.�C��������ˇ�}��c���kojT
n����фR�NǠaw�0�3q�h�&:����T���?X��~7���*v��?|�n���lv�&LIz��^�ߺP%��Ϲ��wW������Y\��L��3���S�
78��u3̋/Si�F�v�k��Ԝ�v�|`pi�v��-�<S����^B0�����3�'8�yN=��_�߷SGtĻ:�^q�<5z�4��@�A�,�fc�kجt�f.�{�L ���+AFj�`�v��ٕX�/�%NT���2��Z��4�	Q�]ӌ&�*�'?����v�����~����b>(�����{ӧ�LY��M{�d&T-���vzw]�my�tŖ\��[u���V<2��v�-�/�0�^!�v)��%1�1)Մ��M��}S�S�����΁P�����r:e�oǾ≱�T,UAt��	�By�hO�{�!'S�v�Z�D�q�������2�_(��IRaA~w�
򻏕ZX~d�o�>�TI��$7H�"S�<|��<�<�7SH�ƌ�=�x{nW�U��9�=lb�����2{s�2X#�*��8*M��B�奊�Ʋ\����Y0.s�r-�+�n�(�]���smMk5!'oYU�a_�bR:՗&�eR�2�M��'�����b��^�]p6#G��<���oa��߮�1E�ft���PZj���HDу��'��������^Wj7�yb��hR����Q�].q�?7%�.��^N%�/�Cǟܖ�r��z'{agn�,��/LO?P�����w�Uz#��Z�α�6����˟<@�ܖ�|�ަA����0Q���|�^��S�UE���8�������Oj㙯�M�l[���ti����(k�A�~���}�@:�1�v���V:U&6�:�r�CX/)�3�ni��>:�όg�����ۗ@f�\>�E�u��K�}�fHf���3��,�L�õ�7��;�1���Ŝ�LT�o�-�P��g�]�,46
)yC��2��E�_}=m���gw�_��	��}�X�۹������ӱm��y���Ah�1P�r�͛҉���������*�׽۸��*�K�HCyIw7�i����%�"�R��sM��z����1��`Q�1���b�}<��M�JT͘a&�����������z����O���O���������O����׏=�'n��GCz�PbۗWa�xr����R����:AU"�����v>�C�y&����\GT�׷��#o�i�CZ2���!ֱ��Yg�Q�Fl�\��B�qb�绕�L��%چAg3�6�&�/�I�%,��l��Y���vI�jw�@��+�f�|�g.N���%[�ڋ��P1�a� ����)�w�`b�t9��"�T��+ဃ������n>{z+�AN	�m��rέs3�u�gv�j^�l�h���a��c#��o��W�'�[P:�frO(�`r��Fs�d�j�#w�x�ѿ��fs�]��Ȝ�ɖ��Wʵ��6��k�ztdji�;�d��9�-�M�,]�g�m�e=G&�l'ՏGFP'-mFwq�F�$2�7mR˷��4��p�,�15�P3э�KAv@���Ќ&�ӭ�r��g��<k��S�?8�ľ�,���ǻ�`�:�FJ���U5�a[�t����|�
��ۻp���Vi,�&v�B����Vm<�V,rQ,��qbo�*�]���]�Vq�[r�J�>�zx��n��*�ճ��K2�۶�Y{It��J��1�{{�d�X��*�G)�n�Y�r.�#�پyP�LagvU�Nl�s�)f˖��:Y�1w#P��{9��{��δ*��K6�e6Vu��$��n�Ѩ�dUl�˕�'Mea�o,���7b�(#Pf��,��vhmK�p[��unػ;��^�)�w�2�����E���P�r7Y�N˪]��*���"� ߷?a-"eZ�4��K&>��t.�z�+�gy�Շ�ޢ,�nL����WY����a�]�N������k����M�p#%jչ4b��B�3�1h���iHRŬ[��0�+�Ƙ#3�J7td��:df4���Pْ$�:1r��le�O��,�iK�LeXS�<�_Xs�(4\�]���m�ZǗ$E<���ga���I<"�sCРç-�����.��0���Kk),��+ǻITt^oG�� �XCO��6��}Z%f(� ���q��$���S(:��v�Ià�P�(�J=ꌎ�۫�j�ڸ�!U�$�IG-���|Q�.���ʍr4|�O���v]j�b�9�z�N�_Z�U�HvD	�ª�]n�d����2��{W/�iV,�g&��:\�t��jP<�V۷�v``�+J���l�o�V�ɀ��s���<B��K����֯���!�s�c��wj�g[�N_�J��r���M^��T���SU���Q����Muρ�sY��YB�0l�A]����)Y�5�[X�����f�_`2n��*U:ƊԮN�p���yٜpoFR�X��=#��+>#��#��MtR-3z�ෝ#]{�ިs9��[�i�!�J��on%�'@�$�p"� ����|���>z,}�o�3�i""��4�EU-T�DARr�T�	�+��7*j�B��.K�������g���2�(9[QEhEEBPD�UT�V�R�em�B��( ��i��D�&`�(�$��RkCh���i��䦋mQEU4�hĒT&�ր�خgj�R���)4�"�h�AE2T�U�RS��j&��i(�� �ص�ƈ4����hld�bj�����������d��`��s�Km�*
*���m�44�Tm��"ӧC��"%Ţ�M.��#gRU.�8��d�)"&�((�@m��h�bMCA	Z}sQ�lD�h�����A����mESM��"�"�$���DE����|>-�M�^��� v��Yb��D�fޓw�P=�������	��ݽئ.V����k��Lz������C�����x�X:��i��aK����x5�)�08��������U��N�zGq�,�A�`����vPۋ+Z�Y�ީ�uG�XR1��oV����/K�	:�A��\���V"��4S�ۏ�Uz�69��Y���(JSW�����Z`|�րğ��2�����G�z�cD�%�ZX����d(*�)ؼ'I�9�N�@�\J�[\vO5>Eê���l�s	�\?M>E�z��٧4���C���8�wQ����r�t�T�a�^�gK�}�?O��O��#[�(���p�v���:�a�6���Q{:��6���Q�@e#֤�8l&�~���/!�N�Τ��KX^:h���
X�p�qb=.��k���T�W�^h,����	���cn
ճ�o;�E��t����xQC���'�߰	���(�>��%��;��.ՙ��1V=2�ҭ�¹� j�e{b�ٶv3��@?pM���������ݶ���l�f����KF��z}\fy��a��۵�6h~g�	����G��4��O��%6�~��SuN�
�%Y)pcW{,��ṹ�ҳ����nS�7['y�m㡖�݈�E(�]tw%íu���8ZZO�������R���}g1��0��)�[�,�;�2hW��d���=t���꿾� �Ea��r�����ϟHb���%8E��aZ�^y��r�k�bO<3�N��]��Z�7-��S;/`�Ɵ�X��[�l��'pЊ�j�1i��H�ї��#�?/*M�Y������Gq_[�['�O��e����q��}}S���=wFDn�s�(�!�^l��$wZyNDn���[7;����Ʋ��6��߰((F0���E��W>�ݛm� �K2Uk��U�l茊鵳�����A��Ju��ٳ���3��z��!~8,�v��vz�������׹ٝ�>ڞ�Ō��	�� �ӈd�M����C'�7.r=�<��S�%�(e��C5�|	�n�;�����M�Q�y�?A��yN�#B�)L%��8������(��h��4odż#�p,o-�#<�:]�r]�vAnm~��=�1)�FE#?���8��$^4
r��AM�~Ĥ��͢�Io@��D:!���[p�����T�``Bt�@��9�;��^(D�9�(���.�����t#����~~�0��˰�6�ʒ�����Z��{��</���^Zvn�������n�!R�,X_t�(�)w�5�S��KVK�]OO9H�Z��V�IZ�����\�)�C��37�{�A˝:���ê�qPwx�ݏ]�T�#8�}J�J�,Ӹy�]�񵘓0K45���Rb��[v��y��&��܏+�U�\�[ؚə�q�5ߘ�ƜE�m��p��=4 �7���2��	t�=���M���:�y���zͰ���Jzk򻔞��4�T0���#ې��8�2m�D���F��ϓKk7r�Na�~@u	l,qD��,�9�ʺ��l�n�p�3��۵V�1�S{4�gv�l�\&��m�8hY�u�zW=���K�X��(`�Ꭵn�w9v�"������j;��� ��k	��1��h�f9#r��nԤ�����`N�0��ǐ�T�q����w+������A�P�΂��4B ����'����s���B����/�'�c������gV�'c�f  tE���l��]�.+C�}�LR|a^7:˰wS0�fc��UTa�1�/mS<����ɇca鱞^'��23�P{�"�'�o�B�L���˜쳻\1ݘ�<����[1���	z*�!\�y��m�P鋇��,�����z���'��N����A3Z�*�N��K[iP?{ ��z�-�Rq��l���rޏg���*��6�/��*�Ajh�B�KV�V��xg�a�'gz�x�+~K+6ح{��4]ʏʷ��՚�K�ݾ��ڝ���DVB��&'K�*m-#�-swm�0+g� w��NW�b;P�T��%n��JUS��ޱX����H�$�(�]�u��������4�/z?�G��Â�g`��c%0�#ú<E&�`&Z-/+bQ�{4�������_�òu�����w��k
,|9ٞ�!�耈���Cv(���%1/	��%.�^�A��ܖ���0v^���؍�ǭ{g�Y��z1���������3�X22z4�|�]5;�o^�(�E�tS*�J�
��_8���O�/�3\���kЗ���2�b¿*�Ƽ3][��T�t:�QI��]`n�eAi��͹mH54��>D�㰌�YD�:֮���w�k,k�؁�B����ă�z^�LZ~d��+�Dz9�	k��y`��ķ�m�S��f�������<;5��ݧdQ��F^�F��J�s�V%T���}��s�&��R?2���y����AÝ�CTĶ*��
e��l0w)\��^�����9���7��c��������5����0�ߔ�G]0͑��>5�����M?#B���=�j��3�עc�O\�sHgn���h�������5�?*����O������Z��=�A=z�_�෪����j\����[�ڇ@w��g=���Y�Y�؀�M��<}q��q��3���[�[�d��u-��GV��4�I�w�tf^��­Vk��j�;��L�9b��Ǆc	�[�F����{R�j��j���{�<OL�����a�������^w:��hvx�����s��;�Ț]���kN�e�.��И����;X��OA!������7C~d嘍��b���G?S�K�AP!�5���>{�/����4��X	](r��/�ԭ�V��v�yn�S߻������
~���>0ջ��H��`܋mIK6�0���&����A�Wu��8����x�t#�fLM�����x���L�Sl	�y��!5�z��EZQ]G�{�^�MD�0�c1�ޭ�[�8A@�����x<�[!kcWf�{b�j���8����W��d����er�
����s�:y�=��.9�!��r�:xk�w��׽��֐��<���v/	����ɼ�����$ȸu]�KH]#�n,�Er�fahk>fB�d�֗a�7'���Q�Q��&*�$R�%E���D�`�5�T��ة�՝������������ڏ���˯��r�9/I��G3x�z���3���»+G�a�噕�\�}�6a�^�m���q#�c�\(�͗��c�uY������:\�F*��k2��,!i��Ur��ш�V#ݖr�j�����j쾪`���@�b�I7�ºV���ݤ�j��,Wӛj��B�v'�o_Y��m�{]�Q�a����� ���!�72׽��n�ڨU��8Ce�=O�^Y���k���G�1c.q���]�lA�4���c�F�=��,;�>���J7i5FU�u)ݱ��^TW�����z�s��FW�-ݚ'!�@!����>�]E���ˇ��<񧪭4�޽X�Yr+�$��/�^����M3ܶ��h4v{Yh@�`�Ьt�cZ��Y]Kw���Ɩ^��X�.��>��]�S�i�i�qhIy���s>z/���:1�qx�����V����G�D��
y�:��T�Ɔl�ב��;�9�+�������E;���q�cU��-�-���j>�~zWF��x���&
z1m��t{�̳B;��h�mw��.�Di;]Hɽ��82Ų�_ϭ\��yǃ���	A텀�Ƚ����+�}5�߈ұ_����O�}�z*�_\��k��&�PH�i�l�tg�NT�������5v���B�+��E~3{7Պ���!��L���[��(�L�#X�LXGc���s�lgAE���}����̱�?�^e�R0Ou�u�������v3f�O<R�3U�Oro���J�p��W��B�㒪Hg[��uњN�Gʖ��s�by��e|�ί��
i]Sˑ�Oze|�v�Ŗ�Y�U�u��M+KԘ��<�PW&�X��z�wl��WW{�y^p��p����l���<��2ǿ	�zѡJ����6�:�!��l�:�ޤ�)��w�Q_{����Ϡ��}���8A�><��2.��:K�0K���Du���w�w4_mܝ`�������M��&�S�v�۝��#�'�LoN��Vɉ�{���C�*���y����2>5ä�B`�=�%�v��`B��4�s#v��<���(� ��1Lw�Pn��zk���mxp�Ѓ�� C�e���kk138Jl=U}�(V^ǧ�R
�s�S$��4*�ø��|r�����{u�͵����ς2/�ξP5��u��*�
�ΞeJ�Xi{:x�A�~�J�!}-����h0ڃ�(�T&7H�T-Y�:��\�PK�XU�A����N:�S��+Q�\����^�@`�Dy�����/B�\�����ڕa8k^�8��J�*v�" n�x����Y{�k��Τ�8>h��&癙��^na�S�;6`�T[�����7vv�1eC/mY���+���v .u�/X�C5׌�,��=�f8��L8���Or�ՠ��x���F�{#%�v��u���]3�W4�]B�M֜��ĜR&�j��i�����%P�x]-ᶎ�Ԭ��"�!���򃷲9.5�������tE���_�� `G�>�C�{aY78ȵTD�L�����s.5Y�ɘW>���5���%�>΃��[H׊xn���P{.9ҫ�7B7�ǫf��r��	U�^�~�gx[X;^�j0Hxk���VHB��M�ۦ���yזu�|��
��w���B,�h��W��P'�nT��{yHZ�]DZ�
���p��8�6�C�n�<G���ʔ{��d9^�Dh���<0����\�K	�"Se�!2�dJxMс'��T�fE��;w�iǻ>����w�<Qѣ���n7�?�^�~~��y�?!)��Zhޗ����u���U�q� 2�r�)L5�BJ�؍�ǭ�E�'�o��!Ŵ���@I��Z�D;�4(ݺGVeov//Y�)���I���z�X)V0��q^�̨O~� d3\���k�
�N��V�l^v�-��P�47��I���]0�jQu���,�i��r��^�c����#32-b�e�'�	�svn*o�iC���=/^�1i��(,WB��L!��W���p��M]Ӷ�|?ay���B�vó"'��5�v-���%vҶ����p뻹r���i��P7��{��ي��k�%���I�Fᙄe�y��[-;��
g5e�:qT:�ɦ+YP7x2q�wȂ�r3�j�^)mVH�N�6���&}�tWc����Lq;�-��o�a�2g!������j�d�'�_���J�s�{���U*.�i�x�]��r�^�������ZG_����_j����S.�m��+�g:��Dݽ+��g�����{2��W�
#>�3�-_^H�Y\����g����.��0���y����D1�'�c���%鏏\�O=�M^a�����kN~]��٭š�]d��l����s���$3q�)��^��r�������ڕ4J�,~P�����R[�u��ۧw�.�
'ek�}nG����cn�$9!�&��1�#�*���U��NB�Ou��4pp� �0C�����g;�_�̳F�,%t�R]�,c�xTnG5n������疙��
~���?��"ǟ+�U}��~]�{�nԩ����Fx��6���槽ӛ��� 2, o��׳��=���.�,8{w���τ)�ߧ"�ӊ��l�4UY�oU� �j��(2j���Fp���y��U��W��W��.zÄ\l~���g��|OjDU�(�v��J�.���+�!��b���~��l[�����{���*[�թ;�j�{{�2�d�^^�9W��J������6��WTo�ޟT�/|U�C/������o�ܰ��L�����R�<g��ݷ�m��a����5D�v�¾��S�A8�LK$�3L�R�I���9�<�ۼ�,KWL!�
/��t�(�f�&�,iOd�z~��=�1)�P6�$�57@fk��싇J�"2�^�� ފ��i�u�]�/h��u*��}Cl��vr:`�I>0���)PJ��y�ᚂ��(.1K��x�}B<��{��=7S��F�/C�L4ۖI����FN>���[�y�Abq�j]4ù�� �-�x��G8���k����P������=��wG�^;7L���]%�A>;��ݠ�ga��:��7/�t6lSA�2r޶�7oMvP�nwD���k�#<�P9w���>/H��0���Ǩm���X�<�.���fZ��M2�K�d�4-_�Ia�������3:��A�chC���`���0�i�^��w�˄kSO��w=K�>H���l���~�a\Z�&+���9h0Y�c�&��{�U�G,�M���=(��~� ��]cjO�߳��N�^&$�ň�z�>�_�����������������������������z������)w_=LOx*}8�Ҳ�Lؑ�r�}�T��u�&v�A�T�E�`Ҽt������d��ͼV�d}�1)˹)��)�A;���t��uv4�	��x�o[Yf��'��Beh�gR��i�tҎu�3_�ǙXa��oo��O��.,}�U���/��G4}+c˾�r#��Yѧ�����v�X]�5��'�q=���W7w�Ѐ��Zؼ�6^if��;]�0=�c�]��3*+���{;��%IN�J󶯨������Buh�eA���c������sgX5͍�3���/������Amv4�GT�f��n���g`�F��ٚ��L��^K�|L�������iX�n�v��k�����w�,���.(�1s}�&%�	2��,��X�Ŗ�=1<W��;}��=�.L4��% �/ZCt�;eb�ҙ8U:kVM�n��5]W��J�9=�5_�^�iq�M�)]D#6�3�s`�w��6fi��zJ��O�%��73kc<w�	�v����| YoT{\
�L\�l�ƦPv���w�'���S����+�ft�(��6&��r�(]��h�w���sY�A��%١���c/��U���ub�Y���LXW)�f��u���zx�H�X��lUfY¨����3�kR#>�1��4���E��Ms�ىᩗ���K�z�)!b.�Gv��b!�6N��iK�M�E��$��mL�ԣ�ʱp��U�.U8�ha�ǽb�^��E�u�M�Jr$�z�������)]-�Ok�ke���e�T�j ���F��N�A�mn�XX���Il��o����M�׏�H�u�L�;Qc�S6�%�� h�Pl���n-f�᝷�k��QS�F�e�}/�#12]�U��h>��e	[ux�+�:Bt�g^�*�x����p�U8���a*X�Wj,$�u��A�y�.܌�s�"rp�	;1���Z�-]s�q�Xq#"@��2bܵ�^��57SI��7t�ve�pi��}k�㆏����]�.�n�P�s5��z\��KV����n<��%J����3*��+�,u��+/pTV��*��39*;�$�2�^��t��ɤ�[vfh1��n�����o���AJ�ˑ�Q�p�/0�FaۓN.=l�MDC��҈�R)��2�M�*�PbZl�ɋ��R�2���M�w^ʏ9��s�9�:�$䭮YeP8�˂��{�V7O��͝��d����3�vΩ�g9'P��91��i�\�Q�V
�4��V�a�:���\P���QH���e,�R���!��Y��8�A�l"7l͇j���.��첳>o��A�<�s$�A���Ev��;c`��DbB��j���.v�jgP܈Y�x�&x�����Ll5�6�jc����|_^�s�.b�`��%U1�1DPl����h�ch�N�:1SE1SM-	�i��i�����SK�ICN�k��U2D������R[&�Mh��ӥ�#gZ4�I	S�i䘒�vٗF#A�X��A�i׮rt�e�[�+HnI����X��Xhb��� �F�15TP���K��OEƈ��ck�Z0it����Ǒ$MSd,`��� �]:*"�DQ�69�s�C�6Γ@U�V�N�F�̕�֊(�"�E9��Km4��JRMP�ΣgUA��p��"��5���1Ȩ����ln\�䘐�����F���<��s���ܓN����EU^�$E�j"-�H���IK�SU�j�֨y:�s��(��Y�>�9���X�Nz@��e��d��>-��@�=ʓi㬃�{���WIA�30��D�yJ���{��1�+=̌\��޳ɖ]����d��J(�����'g:�td�� ������)�������D)��3$��m�S�4�~���$8Y�;[��\�Oݟ�y�_S�0"���2=�$?�����^����`�|F�����Qϗ��c2�P�����}��ٙ�q��z�[��>��i�G�L�I}kO��sd38	�"�C�["�Us�\G'���%n�nOv�j��+�!�PJ�����y6ʺ��i!M���S��zcu�`�jq��Le�ս�f�� &zG+r*ڵAO�xaL"��ʂF���Gc���s~���X�]P��w5Y�sZ{��� 3�!+�D����3g�FA��2ǿ	�F�+U�{'c4c�OV�х�M�7�+!�[�S $�;�8H����	�{���H�Bsz����|��z���Ro{;낽8�Gd[A��oLk��F5�H8vA���.�4��D��T�B���;�t,������"۱ �E�H�s�>;ݼ0������	�G<������]&��gfm���,�UIN��"��4�-#OD��mx�<���0�s��-�Qu8v���(4)Xi0���\��r�'����}L�>M ��X�A>^�/l?��S�|���d��i��]�I�y�k����w�͡w]�V���ueͪ.#�������=ޗM/pY��A0N����FX��'k�^��Oz��;Xu3H��^�1�t�Ě�bk��u�3��l��?������g*z�&�����Q���:\���Y9�Q���?��W�r%H:vN��_�K1�ci]c	��1��EH'����B7���X`���z�l�Θ@qѬhLc;���$�'�s�PK�X
��lD�8�>9��y�[����}��.��"0
|�_��1���!ٕ�ˮ`Z�@J������bC�dN�91�gV�v��cqg�|��%~0�����Z댟�S1���8�4daׄ���vnZ�ە�,�k�0�u虑'D[���<�ǐ046v���;oT����{�"Mզ;��V�r��f��;�;�����&]��[N�S�u{ 3 \@�n�h��ĭ�=�X���^��^=���c���JA�a�3���r3��k�����~�=�/9v��a�ֵ�p�a��\L]�sت�=Cr����ˠ�WAP	I�7,/��kyn����5�?��:���qMC��v��c%~��a�D&�&Be1j�}3#r�ƥ�ww��BNײŀ�7^�iᮞ��$�0���Z��#Uz�C��Sl������Ca���r���[�;����u��	X��7�EmV�ܭ���Q-�p�8���xl��&�7sj��)X���	��ڤ���g��FZ�%��g����«J|�Z6�&��;Zۣږ�5^B�-�Ui�zEuww3����7zN=����Q)ͥ%�gH�P�çu������0[�N�{�	=��j˘"ߪ.��l+��B��5�bu��K$�Y$d�A�/�S��'��L����d�z��(�(a��K��+B�;$��v�l�`�ŗC^X�-4:�r�����k6�3�/k�c�8u;.� t#X������l�(�}&-?5�����T?3@��*k�E�ɣ��w[�[�4@g!�d�z���4����P���T����~%Q�����sǻ��]���)�7��At@�H'���=#�#���]Qßl�?/��>r�9�Oy�3<3.����a}/T� ���+b�>�D?���^@��=	�K�n=�B��;3叧��;��j�4:�Ƨ��3�עc��C5��(���JG<�s߃��r��T����
ƶ	���%ؿs
����_���0oǏgr����5�/SH�;c�f�S�k�{��-���]�^�nY]A�A����H}�x�v-��{}��CI�1�s1{�֧�����֎zӛ\|��{�xm�E,��e�!�!�(l� �Y��*+�O���۽ӄ�.�y�ۏ{,
lG�3(�V���;��
���Q�i��pR��n6�^�2V�:���&�g8fW�K7�z��ͮW�*rk9'�Sk�Z����e!�����Jړ��=&������X����i��L��X79������i�(wI`R�Unz曄<���X��nwr�p��Yz�k�-C^��:hd5�=ŧ7U>�z�m�)�;�6W�7{�.߬�������2�Խ�m�jIe��8��=���)&,!e���`��,��;Ɵ��n��ޥ8�y���O�s[�ӓ�ּ��%6X&Pd֞�	���馞�3j
ȱ��/�����ټ[���C�����U��\��'1,��Fi��T*���Ʈ{gO;l#!瘂q��|8�>�n�
A{^�*än4��'���&I��Ju`%"�RJ�[X���5�?q����=���a��8��[H���0��ۗ`�#��{���I;󀘬�)j�ّ��ٷswZ�m��j��ǣ9�>G�^�QG�Ȅ�SgrD���0�; ��]%<����Xw�O�۝ݘc_���ZF��:��#��c�?�3��$C�-z]4�C(��5�d��s;uL�]!^�����	�� �w=|� ���8��>�r���������Y_��I%:��D��|S0ֵ��-6
HW��)̦�p헓�i�Zi!����|����ِv�"<��JZ[���:�wU�L��l�l5of��#�T��!;m���+5�M��{���z��QWs�N7%�jm���up�K1����o'ڜV6�.����]���*l�H����}���N�Ws�
p�t�z�-���@�����8h!��&�]�w4���]�\:�ku�^����"�x,4����fn�E��0Z��m��`��`����|�ﻵ0mP���ͩ�w����M����~O�L+�@;^&+��h(Y�1��2�[��ս�d_��Ń�g�!��4(��~ɀ�"7�?<���n�F\*^CZ�gͦ�����Yb�HA�|����I�e�`��5���b�ω΁]>˴�X���HΥWz����N�a�z�6��d�Zz�o�6C6�{`��Ƚ+��f-Kk^�*�,��٫�y��`�⯠�-I\����m��gO�.�,p�>��8v�������s�y�y��9mZa'ּ0�z��ʒ5��c����C�"�v��z�Ѳ�SsC;v��2Р��$CƻO��լZ�a�1��=��L��	TXS-�9u���w�O`��m���Ol�?7�(R.'l�8H����2/a�Jt��w��K��<�����_rv��4hlj(��1����oY��4B��h����2�'��]#�F��.?s���/|/g�U�Oգ�ݶ�cm���R��o{��s�&*,qGS��$
H�D����ي�E�4o8{�e�jTW�e��L��6�~2��o��an;/���O��W�P|����~ۇn�s�W�c Lָ�V�o�#�wj���u!2��l��:{H�
��_=;ݼ0�qh�!����L�\�]�c�������ڥ[Z9�02�r��\HmJF"� ���1f9��i9�۷�ʬ�a]�;��gq5�9U��@7IPJ��^2]HPϸgKYaېg�K�-������;�]��$��ʠ;�*Y��Uj��+�܌��Wn�<X�n����T0.��O��H�� `䞏j�'����m�άSf�^Z�Q�y�����r4�6@�0�f�Ou@q�*��Z;R2Y/='`�3h5��OOf]\������`����_8K%D��ƨ�]���l��o
�^~a��� qm�^��+�M���t�]nޮ;/<{oN��+���;���mw�HD�<KA�Q�/�|�y���?�B�~ /6-�e�Ķ� �jyM):��i��nCҺ�t�4�^�z�۳y+u�Dş�v[0Ĳ�7[9�x-U�/[�S;NmG辂�w4�S^�Z�q�X���o�m��h�w�><��A�l&�Z�±�٭�:�طT��PU����A9T'F�R�&�.���;#����V��sg���:y5�!�l*!���t�園�K���d3��Z�	��˯H���Jk�m�;,�g���;7�i�e��}�l�Tn~�hժ�2 a
�3z#��=ў���͊�=���0_��۹4�@�g@�ȻrDxj�0��"ڋ��]ˮ�;��A�q�k��U�	*�۹�ei�@�vHJ�u����zb�{T{��E��Ot���a*[$�W?_O����W'��[Q�ӷz��=�����ݵ�yI�<O���{srS>Tm]���
|Y:I��؛��~��y�Ε@�x��t�\'p��
��eu֮ÝZ��2��]J�n�`09�c��NOwW�V߮�(�43�«W}(���A��&�o�0^���do0���g�6O�����	?s�F����W�4ڭ3�D��	
Od��,�y�l�/gc#gҮ�o�^�r��bo����?t�h�{S��gi���+�P�()´t	W<'
s��-��dꮺ*Дv�y��6��5�Gr����Ǘ�(!��ycUn�����ʤ�N��۪��ؒ�H��U��au��g|�#��]�b.��V�VO����)Y��c�˻f�q��yI�L{����J!�UW^���n�=��z����\��rD�i�}�W����wF���ƨ٧�X�T���NFi��mB�1�m�^�īi���n���"�d���a�&;E�m��m�K���!�"����W'p���y���,4��!]OL�e�i�����t� ��*�dlS��g:!᪑�����"���ו\uoSٺ}���D��I6��%����R.�Cl�P7b��>d�掹�HTK��[[&�ot^��R�	 �?O\�=�q.o��*�T���q�e⼊�=�!Z��:d=��D�$�=�Hj�B_��5ƹe5S�ҷ���`��������p�g�R4��T�����yy�W!�q>{���\Oc�%I�;�H���P۶|xƞ�[V����;=;m��%�+W���z^F��9�huJ��F���~��.ɚ�����47sp+�a՝�E����t4˕H�]�e����U���OsWE�V�\����'�C^fH�¢�Z3�H�����7"ڏ��4�_�N�0����f�B������ϝҒ�E��sT�a"��K�����Q������!p�-���m>N��<�֛���u�{uFJ�K��[��{e=������^#{"L'��5����U�t͐/zM������.���ס���'t?C����.5���'�l��Ρy���)+���wG���t�Pj�v�����{��c�8�ɜ���� 8\�n�b�C��T�q�oȹ5�����:,n��{���c�4����_tu���W����Zb�,�6�H�K��ʯqc��
��̸�qڿ��������`z+�ˣ�����V7��YZ�r��4N�m��s���q</�$�眸���UY#���B|���g��/��M�����ꆈ����9��<�O$�4�_-�C���,�!D���j��l~�jh�}�Ϲ~��z�.��!��|�7�C+�R������xc�X{8�e�C΃��J4|�U��]��n��H�QG�\�1�eU֕o�񆸁���̘��fuKUp��1�[�u:��oc���q*|��ҝ$Y��4��e�#���	R�����`�i��Wg"2&�bw�����h݀�R�f��FEo%u�q��RGO\>����h�75�'�u�
���f�3�
��!Xw���b�n!]x�f�I��9����?l3_Uw����\��OM<z@��<�����mn �iIJ��]��yB�+ʎ���^�L�$� �jF��̑x�$1��v5A�3���V�Y���:��[��(��R�2kd�s�^����P{Ll�l��b���e���;� d�Tk�뒨���R�E�|OKg�D
^ה2��s�WϢ�����e�b:�u��*�qtO��I.�K�P�z�3¥���9v��a'�ϝU脧��;*�r�Agr�;��q`x�����wu���`}I��Fo�|����w*0rOj�^�o�����=��/?����{�ޯw��������w�����|}>>:�W���\due�S�XR��)�wm�l�$/!l�,�X��,�q뵦8q��^b�2`#���)�r9{)�/^E���(�N�Qb�FsS�$�uVgI5�.Q.�Η'l۾;Q�������jt��NYj���8�)���]�����o�
�N�ML�QU��6�P��f]�Z��b^��vS(��]Mk��X�76��˘4;��/%ϧ��.�su��k��k�V�920^�;:77G��t���!��#V}kBSS��c��040�Ok�nK�J�n�\�!�B�I���yR�rWy�b�tjjc����#
�p@��R�g1�HA�]Y��: �[9�٬���}|R��g#�A�w�{����f.y�AWV����)bN���om��KDs.��7\F4�ڄ�3�H�m��XEj�&7�x�5�5�������텨)qU��)aT4Se��}��R^t��I�Q�����yI�6�0��P\Y�Gw4����!������F���#�����+����ů��Ӻ��^�q�H���`ч��:3Ii���:y�0]%={��ۜ{XZ���ɜ����,���eJ:�"+�N�V`O{}�u�S�n�m��k��Ն�)�h+�܌]�V�yg(�����1Y%�i��A�a�k��2�(ovg6�f]m�쬵ˠ��sI�Y�x�G�
V�/�ei0u��.�4L��͔Bz�-���oS��c�.L�Tn��
�[�����$L�`v��@����`p}>�������w.��+*bH��u��{�ڻ�45ò�ktZ��x�c�t���hl5m�q�Y'X���9��#53�RV�Į�-#oM�l�|y��-��\+�b��$m�'Nn�U\%��I��p�Z�hH�7���.p�-N���%�N&`�ݶʭ�ѓ��E��1ؒPeT�����3�fe��nΕ����wu,�v۳�"���W���٦�-Y���4�Ε&�c�e*��z�ؙǶJQ��R��_<p��Ρ��mV��ٹ��̮�XD�ن��<	����.#Z�uf[��=�6�6��㮻!��MHsEa���:dF������q.��}w\���Ľ�V�ٍ���Fk�Ԩ��~�ޢX�ۧ[���󉮤RŢn�u�X(����zT��YBWfU��̜r�N�Q�&F�1���IMږM���GcNʬS�hݳn�����;�\P�7K�.�蠑m�w��U�#�"sFf6�.Η2"O��C�d���N��m��y �h�{�btq-��U�7�7g��S��kD���2�[�V�/����j�;M�ޘ�|~��(,+��=È�F��⼃V��P0ʥu��	�F����BO�JL�t�̗J��]�I��NTE�k�/wj�λ�Z/����L?�e}�|<A�ҼH5,�QA5G#UIQRS�~��͊��[Q:\������Q֍%QTD�D��吪b��h���+s��
Z�� 䚶�M��� (��!*�9b))*��,M;8��y&"j��P�-QU���EE��:")����bvuS1I$�SQCE�QD�3Nۑ�-����)"��)��b���&����Iͱ�E�c����&�cY��n\Nf���v6�clSZ*�lܢ ���i��&�9c�j6�ma�L[f�Q�(�$�ߟ����7���m^\�s�s��Hs�AF��M^���4��OSAJ
�:ys��&�V,ղ�k:F֝[��*�s����y�k�r��#�j~��#�׆�4ݾ�Ά�L߮����E%�:���뤒�m���>ţ��Io>���p�0-1����}3��HyY7��zs8�o_�ɑŎI1�'�M���K�ҁP��wq���f�%��W�M�]û2�=��	$o�pT`��q�/u�]���3o1�~��vۼ�v{ol��_�
g���?O�	R�<�	4�w�z7'x�S�z�j��<�rb�.+5�}��(��S�,�|����{�����4��Z��u����0��/���Z��i�$����n��F�n�H�6RUhʡR�Q��4�E[:�峌pSB.��t�1��/�m����A
§�PRz�O%P��ګ�ei�X�;i���M�M�r�
؟?g;z���Ot��].['}@S���Ӭ�z<��K`�K�=���t����Uh��v��s��vo��y��R�6I8-d����s��u�u�$�R��Ռٌ!U���v��0N���]C���{��z�0�Dt��t�a��Q�m^m�(2�-��ʹXƎ71�����j����S{��;��|�r�<u��/cvy+�*�t�go6�}xy�}9� �m켢5ǚ�����ƭ�nt����mlH�n��1j%L����l��Gu��z8�>�S���!��#��c���V�{��̭ti��r$U͑;VA֎�ظ>�v$���+���7������ޑ��q�k�TB��5�ݙO���&�y�~��{��U�O��o��G���&-��!3��y׺r��P; ٥C������t�;#�Hm�e4�����������F��	*r��?����3��_[�v���҄��P~����vf9����1@x6v1.�m�;,��w'Ăތ[�m�ϯY+p��gwS�)N�9����C0�"��%���~�[Q�3~��~�wy+(�ݻEy�(��WJv)̌�S���A;U-��\>������{��WGʒ��ep�4G�:�f���{��U�y-���8j�!��ƴ.pf,k�oUz,���$%�G��:x�J�`�����c{��7�w�|r�ɽ���M޹���=Q�"��.�L5�i�����N�ǽ-m�Cn�d������#Y)+�z�+�$�os� V�Sc>�&I$q�fڛ�Q��ՄXtW�l��9uy9��{��[��B-����J
E(2	�T{2�\�w�^]���n*���t��8B��w��{[!����#)ь�۳�m����F��,y^����*@�%n7�p�n	%I���;&�r�5w�ү{c���܏m����p!~
2�T�sǻ�%�c����׳y�ۙ[d3ǹwp�f>�y.<�-�ᱷ��6���뉛�����{�O:��\�2���l���	N;��0�
Y���z���qj�^
:�8Ν����3�t��8|�i�{��H�H���c�o��e���y���6Y�7�bN~[�����[[�wt�]ä��*Ui@5Y;L$��Zp��.�TKh�\w���-XZø����4���մ�uQ��?���}��r���O7v�N�#|�_g�޶.U~U�znm*�$��Y|^;��
M�Z��y�D�O�+"��k�`�sW�W�ɾ��!�	�������f�j�$K"�k�7cH��������r��*ՙ�eG΍�����V���f��+ƈ�H���q]���;{a-��������F���rGdy.��+w�"���A��KTg�����tk�o��]�A�o��ρU�s�+�n38�����{U����m�Q�;�)�%�du1���1��a�dU%R�h��4j������1�s{�7O��e���H���<���iC���+���?G��q��ó?/{\�`ğ�e	��̬RB�����|�y8�ڹ�+u��.���^q	�g,��b4U���R�f��2+JV��/v������U�P��V�%���oN�z�_H��7 �p�Z�hF.B����*Z�;��M��Y�G��w���b�|s4����y9��������-��i�:�-�#�2����+�A�#A"��8-nS��ȑn�0B�B��A���������a^��#7���7|�R&Z����ngq��~oo��UZ��g1���荽OO|Qӊ�H#��T�V�6���Oי33�;��:�E�0��++�wL��9��Sp��W��[�&��<=���8�J�E�⽷��j�d9]�α�g}�.����]����n���v��<3�!���b�s���w�x�������rU��j]�����2�̿'�^2$�5[�CvC���_Y��ؕQ��&�*�]��U�ս���i������8��<[I���o;��$���r����M0"�чŗp�	��t�^G�X?��9��+�W?j�ΥFcD1��]��j��mΙ�˫�0��Rx#Cdn��a���އ�£��w{u��am�u�CyA?NQ���p�6��3�,�B0�n�.ܜ�/���خ>�v=v.2��TLzMqc�LA�]>���k�x��4�Gǎ�B��}�G���lw�3/|�{����!E&���y=��rZ��x�\���.��ϣaGZ�5u׻�3	"��)#�bf���>�������nY��k�zJ�fR�L���;��o������{���S�me���|�.h�؊!��+[���$,������er�*m�&I��S��Y�
�SX��[��s�� h�N���Q1��]O.�˻�ɳw՜&���L�cT���a�ivm����ո�)A;�OjA�@H�]�SI�{�'�^ٟzN��߮%͍�t)�#�طڑ9�eΊ�ޛ=�79Cx��껜$�bS��ڮ�^�0k�7��W ��9g�ꗀ��j�����|�O��V#!�y���:Ju��}��&��~��w��1�N�K�"	��"=�ƽ]Ԓ�6BT�L�IM���EH�	�O-��3�Mv�<�pEH~]�<[+�/vy+�[:
���O����I�j4�%sϫ�;�?|A���ڷ=��hOZ؀Otp�7=�3���׽ݘ��\er~�f ��3Ћ�����	~�}���*_o꭯�SU�wzf��Y�o��6�|o��=�_��A��"���n%�;���'؜V�ǣ�Wq\�3<�#��N�|��0 ��tg4:������=��)ˊ0>n�� Q��د���$�Ρ�6�����-B�z����o:3�c��-�O�5>a�y%������Rr��Jٿb�r�.�(�4e)�7O��g�[l����O����O��d#������!:Vnc�F9oI$�F��������*�� TZ��c6�Q�ER�U��LPENS⭾܈L�ٲ�$�u�i�UU��7Y���Q���9�.���Dye��=^/�>�n��N��/3��cݻ�/$5�p�a�Y�į6��p�a����N��gI�����q��R��Ng��!�
���K��N��.��;�wB�N����{9���υ�)š\�Ee)�E9�d��c�<�o5R0�N�(�v�N_N������f�y$���:I��$o��jE�(,����xV�w]J�gww`�A�L����\f��+�M(2=j�{2ni�΍�_����vS�ޙ�ܤn}^����☽�2��[P*�2���F0I�0o]�湻	g�rmS�궁����"�q�v.�ԍy�	^�A��D
x��r)^d���Gry�4�0e%q�T��s:_��B��e6�������K�;�[��ջS�X�#k�s���l���m��Ӑ�c����{|�y�4M��J�1�4�<�\���Lݟ��P{��$�]F���3fx����|o�*�v�b���2Ve7k���?�����j���/��7�n;�\���w�B8��85��F7�! ����,�҂�s�2�gV�]�m�Nw"��{��ݡ{�ԧUݯ ��������6�
tZA2ζH[*{����r�D3멈����l!!�>3һoZ؞���J=�K��mna��"�mY9����i��_��������J�һ��ʡܔ�m���J<V'��a����/��ۻm��y��)
F�o,��tq��}[@�[Yz͂ˊ�/wYz�����d1����b_�����y`���r�yf��+]��K[�&veդ6�c��=A�\���ϡ;:��rJL���iS;��a�peGf�U{��3������{���KA�W u1�i��E�C@��3;��r�N�KR��B�AOAa@_��]�,��jγ7�c�����a�xJk��SwY��GP� �T���*�E��ݝכy���i��nP�lva�Aty�6��dT�K*��4T���<�Yb��Nn5�QNm�<�Q��4��٦]R���-`d����M�x�l�tUs};n�T{xs{m��H�ݝOO���#��ƚ�؆Mݓ��#�Q�u|�ۮU��7����T��/��	�M�\t�z�XiƚUE:��tE�W�l���}7����9�4�,ʁQ/s� �8+�`;�h�b��*�v�B��Sob��=�\p�4w*�{2zi�M3�w��b�߿R����7Ǜ&b�1����zG��$7"�.���9&����[��fD�[���f�O��f�֨���q��":�7c��䒶�R�2�[>j�3�Ŗ��X�1hb�d_a�`�0��: �Rk��uɿ+=H�ڔ�-�z{&�K'��q4��lf���g��e����wH��f;bUGA�KR�����yXGggvk�a�d��; �>���AS�L��˕^�x�UR���u�q��v��nq#{������a�|k�uOj��ޫZ3�1���۽3{uDY'h��Vt������G1�-T�,�����ax�޾*�Ѡ�Q�'���q��L�쳦�|�w����L;�9汔nn�j������D��!��E�q�]��`���Q�=W�o���j�wL�K�L�y57��i����/��[thY�����Hkx�~��V��s;7�N[;�׏�T�z������h�'��Һ����2�cZ��{v�|��iH���-e�v.2�4	�#�2A1�WN�sJ�B�����Aǻm��/��`Y��^M�7�:e���!0�[g��۲����O�)���l�#�s֙��S0��
��]u�ǳ0��+��bJ��;�:�����5ѝ��zө�k�t���Pc����5w?P��n��+�Ϣ�_[]>�^u?eS��]�ڐ3�T��.��yj�^V}#e�!T�?�ѹ|��2�=<f��{b���xu�Z2�B7'n榜�l�a�0@��j��\�L����x��w���/�]ӂ�a��#θ�y*���}�����]�Ns+����ݖ#B<�͎$k6��t��1���d�$����،����=�Ye�9�c8"��-���l�u��n�<��iĭ���n�0���7����w��:�d�)�o�8nt�8�@8~��ׯ��}�=s����������������{�>�O�������۽�����kp������51ˉ}�Ʊ�rUزʓ{T����A��Vc�秲D0j{ݵ���k%�L��}��ۺ���:��^����Mz1DA�!)��6Հ�*�
��;��;�`��w��!������*a_6*����p"3C�O7:�t�..���"��=w�0[���ӄ���鞢�r��5���Q�/���O�
���<Ƚ*��֘ǧ;n��m�N\VN���*s����qWT���֪�3��ID�p�±�:$�B#X1%����l�'[�j���z��nJ��3Q�B_N�B�u\�n�ݶ�w��f�.}���A����홪��������2�G�n�]����a��rNJb��f*�*��|q	)Փ��hө\��6/t��I��;]��X��u+�X)n^�҈T+�{�7$U8��Z���E���JLm	g��q�N2�+V���$�[~����PV᥏(�F�'�6M��ʵSHS���}�/YiH�nf�n��rv�]X�ԣ0��e�է����o`��}k�)�>�L��{v�Jt��D�{X����t-x�w6eMX�����Jw҈���'	ѢKZ`�ں�F��sP��.�@�n��s�����*�wT�]�H��[�ٴ�6�k:�7D�:Y���^O��D�zk�����x�\JW2�\�
�9���bK����S��j��T{Ϡmwl�����\���I��
�����֢�o�3t�n.j�b<�G�V�M}�yJeJM��E��J�YnZ�+zsbe�J����\��^��
��雽�WFf�Ϲ�][��ە*��x�^�-u����o]O��v]�x�M�rp�Z��u�7[��O0�s7�EjKk��n]���^���y(w(�ES�8H0e`�<��.���;��-�t)�0�Gh�1��0�Y��ƺ`���͌��2�"�w���C�7k �ޜ6�a��f�O�Ne��6��dB����o�}�7]ү>#�u4Em�WWm@�ǡ���u��I6���N�f*0�>})��!���Y�bo;Xūɇ�ؼ��;�r���t�D�v�����G�Vj���p22n��ĩ��_�T�zm��/�1�
&�b{�ԇ?�3�=������x{E���-�;��8U�d8]��i�{��6�)�IUAV�-60K,����c�+�O��Ģ����s���x��I]�B�vż������v�t2G��6��F�J;�ZY�9��%��*��z��[tV�3%G�#)�rɒc�$��Qc�}N��r�V�)�Tu4�֯*Ի��pqs�2�[����`+�UQ�����h��͏"�*�C/��'*M���W�S�W��|�2����1ڳۥVZ��d�J�GA+2�"�T{���N;��qө��iV�X8���u����7��@i��uy��þPAE��Q�9���3[QK�cQi�u��s�lc`Ӷ�q��TZ�h����ӵ��Zئ1a�kkִ͋lтt�m�֫4X�,�Th�E�AkUQ�q���0m�c�F�4n\�TU���V�N����kQ��Ή

4�ӈh����Q�VɊ�4ӧs9[kEڪ �i*(�j"��Q�$�A���c��E���*���
�U���.Z"+�ݱ%Q3ATD�[MU5U��K�~����m�
���ѡ�R-�i��P��uT�T[��ү/�wV�cD�t�{���-}��P��bBhu�#�nz��3'lF�v����7:�-������)� �Ai��I�B)�KAP(�6\M�JM�ʑ��6D�A�I׋IS)�n>ٽ������7y�X�'��@�
{[3l��&��z���i+K��]��
�������^]d�ݙ�;�ˍWgt�C8�PE�+�	�6�A�[��fy�! 0�ad�v��a]�w������T�d��ڡܗ$L�*~���s|�1����-�S�&|:t9ѕpuL�d���[͊��߱���h���P�}y��7/�%���wTpM�e�O�8%�ۥ����l�K��L�7bW*#9*�Ǫ�9����u��V������;��xVkg�m��/k#OQ�J4K�y4kz;�nx!��{�:�)����Ю�>)���!mK�3*�έ�������ݧ�+�	�[=7��}��Z�<�SI�^>W+���=�34Dʁ)�\E	�o!�M�A#����v�a�JV���3s'�1Q��~����a�T!g���w��R�>'�P=�^>og�hAٝk0����v�ZM7t�O	n�4{��1��[$۷y\��nM�U�F7�ǵ:�����cב�;z��t�{�nOa��]������N�����0n+��A��2����WƻZ,���ǰ���qen�Ѭ�5¶�L9S�X����8�|���E���4���|ځTL�IP��5�ǲd��s}��:Geުs�����-槯"�ۇv.�Ԏ	̸�w�9=�C��÷��n\�aTh$�S��]:����H@~
2�V]�<���UG���"�x�ǈ�8	��	�3u��:`�#�B׵0J��Z��`D�Wv��ws�>̃=|�h��irwֹ�Gl����YRWF.؈�|'v_`�>@� n���W_j��D��Ji.���r����OO��{OO}ݽL�q�	G��aw�]&��ʡܕ����ѫ ��]q�~YHS�����g�j�`��# \7��,үtq� ��\sŹe�TuEQƦ/M�/�}�ߦ�0.E;��C�l�?b5f�ƺ.SsX�Ӻ���2󷪧�e�s*�&; ��s�1�mׁ8gU���z�;͌�X)M�C�0���ٺ�|�ﺌ�әM���s�����2���Ul�t��gE��03t�{��5�o�s�Z�V��������/�uZW�3�u�D�ı̥U�=�g,���U�����1��!eq�l�>N�s���9<-�tS�z�.}�%F�H�G�����8z8w:Ic�M�1�����\�3�]Ε�o;w�e�2:*���̴�Ă�gk[j�E�+D��#1��l�ӽ@踊C��Й�����GP��k�]��2xȷܽ�Y�6��N��j�3��S��Ũz�꙯Y�׬��_g�fQj�f��aɣe���*�9lv�D��,�+�X�� z�:�t ��MjS��{On<���7o����PyU {2GM<M3�y9�		�1*��9���=����9�rH��I-�E����kr��̐޻fͅ7���c*�O[�*�d�b#o����r��L��JH��ef�Ӛ�y�O��vf�q-@?;�i�
�)�66����O7+kǥq�ڔ�E���tIz�����ͽ���,%�G'���]�Y��Ī�.�7Iw����Jc�)T*�U���LY�m�T6�6���z�vv�h��W�6FH��C�m��#�����+�;
��Rq�z��ɒ�:�$����̎�|x���|�7�hI��*p�h�Rf��u4�U��kk(U�vN�Ō��:�gp˸������=<���tZl����>�ɂ�\�s�`1��m��{�uM���ȴ�5r2�wA��t�|�͆⺣�5���dw8n���i3]�Әr;i�we%G��`u7F�G4���:B�/�z�{,<0�>��J)�-ђtl�ӄ�bF�w"����mᎻ{����F�x��;����D�G9>&#�W\�R�w-���v�Ot��P����1�F�M�=î��������?��=]]!�Y�;F���i��Q�`=����ծ�D���3�tc�����3Z�-���4�	=ɦ�ۊ�-㡟�3�J=~��53�Ѯ
���v4��ӹ������u� �
T�%�ה�\ә��z�Bal��׋���k����[ݪ
�UFDxv���ܒ�hʡ܃�sSNdU�z|�C�A�rk�F5� �Woά���Mn<����q�$�Eq�>F��V�f,<0�̠��f�9m���e�j�o��Mە��7�f�9�C����{���9�i��zG�rMrb�r�[�ӣS�|9�J��	r�����u�H+2n<��j7P��y6ǟ��t�
9��e;m3�]��cN�3e���ՈO�HnAH=�<�BP�����E����by�����]��s��+K�d�����Gt��1��l�F���.O�/������v���"�䭠'��:�G�����U�7u0��h,��s�^owf=hC�;g��C&�􌌀���#���J��n�k�f}�W;}ڲ���"0��'���:��>\������+��C���S:���99��g�a�ȝ#g��-Z��Q�Y�@�֐mt�`����6!4��̛5�s�2s���i8�gѾ���L��m�{������O�"�e'��r��k�2m��uo_�R��7T�ˁ���W��y�e�;@��q��f}����cӹ�����L�&��.�Yl��z�~���p�FCٕr��8z����R�]!�k��;�/����%��m>o7��c���3��c��ͯ�:AE���5�J#����ߙ�����c����\�$;��ZwB����rVFf�d2�gqu�B�s��O��:y�
y�u��G{��h��ZT:�����:�뭔��iS�6�zN):�ދ_g��O�A�8�����S�p��B��J~5�Z�9�_�~������&���`8�F�V���h���b��KX����N�Yܪ�V��#:{�γ2�kۗ�!��C��J�:ٴ��.�����l�';���#>�����Y5�#Q+Ġ�9�OZ�w���v�nnV	���ӷ$d���9B�.�c��m@�a&.��4F;�]X�[=|Զ���V���̠#�:�l����O�;���#�pݫ�X��O.r�e�n8����U*	%T�p]:�i� �:�~
������=��6ۻ��w�R�׾/a)ĭ��6yuy��l���A��:�.mLB���f�[������ǆ�yWF�+e�k�8�t�[����#Wn��U�G<�ӡ�ї��"#�vzz�ئz��ZJx%ܻ��oZi��3;�OI�������i��yh�ҝ�{Y���q�򒏸���9~3`��`��j<�]ޕ8�G�ڰ���uA^{X'h�F���F��L��L��0$�cM����ǜ
Yz�5�U �����4�k�x�WM�!�
v_f�6�3^�lT��u��џ��vkp���4g����K�F)d�ϸtY������GK7G��y���.���a����|��~�܁�iW��VvV�C��ͧ�SݗW+�uU�=	��Lo���=��C�~Gr#��ꍎ��볚{��\X�/�������2��(rfç��)���`a�.N��l��������/�.�=.	���^c=2��It&.p�� �o:-����z�S�c2���$IDi��»-F�>v5���:�j�z绫n�2 �MvN	���˴H� � �C
�h�睌�{���KogwH>ˮ�O���`����y�g�2*F�^X�w;�c���%퍍�B�E�;��է�=Q.gG� �C���fJ��8!�2����79�r���'����=�=4�4�=
׏��0� m1��7:cW��չ��[;r\��M�۴�C��ǳ�>�l�����[J<��rRf��6�ҥ�_5��mq�O�x�(�f�r�2bK�v�Uz��6l�?��}��z�U�H̬)yA�)�9l̲I罗mp�m��X/`����ոU� �|�jd��^=���߽$�\䚠-Hܷ]��!�����15�����!Lp�m�m���Dq�d�t�"Fο����a�9Qsxz���=u#�� :]0F�Y�^:��=+��ԕ2c1ٯ�.��3Sb;�;����)�I�~��@fz�bUC���\��~����x�Kd�#�b�~�P�Cq�k��d>�� �$�1N�3̺�����멚��w)�V�&�&P!u���A��7:��~dsO�?�o{0U�u=�֏j�'����=Cz[��%l��_�ߞ�p��թ�I ���i��*=u��ݥ�~�����c������	�ŵ��g���J�|6�7���с�&}��b�\{-^&L�c�	���b�=��e9���`V�:��� �E��£U���p���7{� 7���Z�3�ů�  cT�d�-OdV4��ecu
ԉ���]���9F��K�e[�u�K��	բ�������͚ie�)�.�Ԡ{�]d�lL(��\�3*���J���z�!�̫Մ�����U'\�.q��o�칚8��l��E�ǎ��;l꛲����[�yb��8��f�r{x��/�xs�C�l���L{T_H�9�����u�:٪��ܫ�6Ժi��-57�{������<�}{jGE<{a��t �y����'��K��Ne웾���"�*A%-¼����o-M�9��΅&�3^��	�޾��]�#��F�/�ё�+䌝�>��!m���<8v9h����d��J�}�n��G�}���#�p����� �#D�T!%]DͦS
���mP��z�r����8���2@S^u=�Dvc��Gɸ1��nc3����c��������ؚ��:���\R�ü��:Ki��>�e�g6���ވ�;���8�WFv�-��� ��d�պ TY3�iIv�^���N���*�׺�b{�x� �~�7�����
�s���m�~��{�����r=��PÓܺ4�N�mt�a������W�)w���yX+��:�5[����w�m���i�vzKDF�FLT�뫃:맪�nuo���u�J�΋�\���t�����L��9���R�|5-�W�W��H9˪t|�gWF��h��l��kǇ4c���	���nU��P_�?O�.�Ǚ�w��ܗPH��T�E��DR��ƙ�ZOwq����O_�X.&b2 e�_R���O��eܧZ'sA�f�|�����+77T���8�bHc���5G�lȀ�Yl�n#�-�fc#����f��iO������Kx#3额U��"ߞ�8�����Tͣ7u�5[��f��Ϗ'ă���<t]N�?H�g��!]M�:�Y�A���Z���}Zwn臟n�4�9���ݚs9,�̝�̠d��Y����b/1�\3?g����r��J�:ӛj���D���o7/+�{����%��¸��{���E��Q
��(R�<a��<Ș���r�0��m=�t��f����ݸ����}B:�A�թ���|ЁS������U�Ӵ��������W_tq�W�����e����dy90��n7 @=��O��������f||||||||}�>9�������}>�O�ۉ����zQ�
����!�o4��0U��:�p�Xy>�p��U^�dM��nu6�j˧[���cb��U�N��F[�r#Oh�z���YVhR�*i`��v+�(��=�pZk��j��[��ew`��{�:!��Ө���o.j�"LVͩ������ԇo�M����_�A�x���\��K��7�eC(}���,��)��x�����@���%�ḷ4s��K���*�p�A�h��6F^ڣ�M�b�^���/.�X�Z����x��R�eI,(��݅�ڶ�cGqu���� N	}�U�)P�Åe�ӱ�IR�z��Ek(�U��M�p�F�C���������{�O�k�T�ڥǻz��S�*�Ɵ`��\�J�ý��K��/$���.�sf�����v������D�ڵ��-6aŔ��u�is�6L\�Ӝ��Ʌ��}�t_-[�f���������T���:��dYJ�λ�<v
ׂ�m�b��Ƅѩ㝈։�IL�2n���T�n:.��5��5�]��ګ�ëާ�-hs�%B�*YT]��Dr���%u������J�Ɍ���wFKr�v�2^vKmGj�!-��B�J��}�A�N�s%wj9b觛�i���.�E:�c��.Ƨ�6Q��F�ל.�Y�L�yp�̓�H�����`7���ש�c�x�ݲ��Er�m��D����Gג�Xr�ޒ�JІi�,����q׷W�U�1����؅>�6r���8J/�:��zvR��S`��ZT{.�r�dd��9Ǆ�ۧ��]*,�q��l���F�s�*n�fk��"�"69͕Cu:�R�o)�>;�p�n�D��P��9�y�8d�[��k�����5㖝N�ȫ����㶞@i��nI}!�T��9EU��ԯ���4��a�G�9�y���nf���{�5��Պ�}n���-b��;au�&$X��{�n:�_Y�M���m>�h��[�:��x��*�~�d�hnϜ�X��`s(��^Bnv�T'V�w��$6̥�C ��cf�!0�C"�2�#�ˬSx��3e�C
��BIueN6�ʥ�X�9���XcKm���,gN=N�^fa��%����\�םM�o5�ʲ���
絗�yE�Svg�k�2AN"��i)j�Xi���Q&c��%ηf�"����3E|��ջf��Z��l%�QO%Vc#�̧צ3�ei���75�.��z��{���|:���6*Wgs,}4��SVF�F����t�u2�P]R)LN7�<���5���"�!g� �_������#F��r�j=����gIvn��Nu,����|Э�2�)��q߮m���᝭��Y.�ӌ�0�I�bL��s�y�kD�Z����8�65�SLrMZ�)�ADƛkY��$��D�hƫ�9z�S��F,l�I��6MU4�֨�CI��E�ĺ�jlF�EZ�X���V�ZG�F�S������֊Nl��4F�"�j�E4��Ō�#l��6��6�6�c%DPR�h���h�.6��,s5;5Mli1fM!��-8��T�M"�ڃcRh�E-Z�QF��AcUY5Kmh+DY�A��-`�����g�#���kc&ؘ����Kf�h��&Mb-��XٶN\���mlQ�F�[llZ�v��UPQZMQE
 ~�����+b������s���u4�����qd޽Gr�JƔ�r�.�����3�y�f�n֬\�;׭��s-�{k��'�7q#��'�T�U@?\uө_��t�B��rE!��}ՙ�o����JA���%+n\h6ɐO.&���m�.߸a���z��,�ö���e��gT�+��-sd��W�Kő�5ڻ�n5������ao��V"��Ov(�Y�%4�sd)3v3U5�
>kޣ]�����������k��t0�q��R6Mu�ʯw%z�S�c����ݏ�M��_�s寨/�k��
3pY���^h�nܽ{��/{t��Ki�;��]a�,8>`D�y�l�+j�^Ix�ݧNپf��Gg�_eW����1�v��1���F���ӘI���]��c��T-�C5������É%��=LwVf��E\LgL�K��<E�Y�k��t�̲���D���<��ֱ�!�>�3����x4�����nmU����%v9]hwm��N�n�)��Ҋ(��C��;y��\��ަC��޹�g%�3{�;FIy`bn�5�5��o#��2@�u�[�*���KULP`��̩�o�J�������n*�L�8��_�?���=�4X�E�G�]Veǭ:��*�[�k�����w��Fǟ���k��[���`���ꧨL���B�%R�j���Øm���}m�Q υ)#m�����3�,�&�ŉ0���D�6�w����]��)F,PW^%zK�K}ي�0i;�ݜ�;�x;6�l,�;Zz����|#o�[RF��T)�3����:m֮�j�!L�4���Hp.9s��2;D���H�c�I��$K5�oX���;�/,��:����sǈ��Va}rUx��4*.�:x?0~�f6cM��(%�ˣ�0�Ify���\��jI§�^������k�:���_Oa�O�����ʚz[a�;�}[��i��&�;��J�Í�f�;�ϯ{*�T��M*ݓ{��F[#7�~iT�M��ay�zuw�aP(��v��[S�ͭ�T��s�uXk��v]��
�}kW*Z��Q�C{J�n��!���<�����+7(�u�y��9@��p��ݫu��A�j��u�n�o��5>@��tExݥ�+ޓ��A|�eu	d�*7�X��{{&���"�dT]@��u]��0p���Ou+�������TP��_sY�t�L�8mC���P��]��x�6W����7��+Z0����UWv�}���1���_T���Z&�5�5Ŏ�=��O�a�;6��V�wQ���\�V�#��24YgTld�?���;v���x�n�(�Z����g`����D�a- ^_��� jXJa�)٫�k��ƅ����ui���5�C�ot�4F�MYK^_���$����Cô��\%k�ff� L��y�<���6�%ּ���74�vX�^��bئ���4�F�?yN�եP2 �
��䕣��v�'/��J����������b� �$8���;&�������G�u��#ʄ<�sg���'4�]��tM4tDd�Q��m���e���w��u�U�x�d��ڃK�I(���(m�*����S�d�j\���i�2ƫ�.�p#D*�&�lq�P��"��q�-qم��8��[?���ͯk�n�%��/�<2Z��*PSj�+�%0���T�'p]p�j\�.��FӚeA5��{�lz��ӟ��e��ğ�?_K]:�k�*]�<�QU����ٺ��}����WO`#H�n�!gl�_K�jp��� �쭶F��y�o�nv����gTwz
�����wQ�a"d.OҌǻ[a�w�
��4�ڃ[����z<��ݠ6J4���)D��	��mq�S��Ϧn���_d�޺~����;�!��q>�.�ll�����r\���/�TR띳�^2�	����=5щ>��`�Ɯb.2�e�.u�֬z���h�˫ɭ�������u[u!�9�g���!T�3\��ל�XK��	�U�˴�N�gS(CK_���pv����]����<+&���2x�QN��V,l���y�V�t�Ϝ�F�>c:y�D�w���}��ϭ3�I�:���������]j���v���w�J���5%lS�3ȧ������
�N3K;�OTթ��[��lItG8��ƽn�z����@��#ua{��pR��>�����8N���7�V�V�/q��K�f�^�/ ap5d��Sq��Q+Z�h��-����7Է[<����d��v�<��|x_��$sw�|�D{p�z#���Ґ�W!�	���dM�mj[��u7�O"oN���N��n��PW���dB�^�3�Q	A>?3���	�W�=֗�T^m�|�y�m�*� �����T���y!�S�UϹ-S�x�v<�U�JԣA#*��v�}��H�g����Ewy���T��|͞�~��/y��&۠�*W�������u#Li�	�m��s[�����{��[�O��WK#�����`7.4{�\��}�/`���6���ͯ֝�����3�F!�}���#�ʚ��`2olzԤ&�D:���3`��S�>�9O���^���-�����ئ}ֶ:�S���:}�:��y��?/r�^����6E�^�7P?���~Ǟ��ǚ`��6�N�H�u�v��5Y#i�瘌�7�z6���n"�U{����U;4֕b
�8TRh��dC�C��b��"�N5�v^a�4Y��mf��E��V�S^�5|�(�h8����c6��(u7v�2��i�B>�pʼ�5��Q��V-�_�0�n��E�/s�|��fo$������,����lRb_���7����L�=��б�_���� �p^#nj1��;��Qq�h�hº�}�\X�Lq�8Pc����qh�K:�������75��s�����%�w�{ǘ�Z^��5�[�v�i7����WSa����C�P��^m�3,����%r�.�Y�G+��mx/˽�_���
-T����ee�G2o)c/fZf��J������'�Ee�����X4�=T�zf�X��:�ȭ�;ػj:;�c/��_h�Z8�z�����qbo�fX�q����<�{���r{:��W^'���o��4�@"� f�=4�<�f��{��[fL�ç�턟�X|#l추����"�$�>ZQ��oL�x������z�cNrlo35H����m�G��7a"9$�t��{`��V�6�*���g��O�
W�[攪6v�f�o� p���gL�7�}a�N�3�t"M�v��r*���tV�Tǋ�U%Gw:�TSk���`�;S�W'7z:N�-�sp���i�9�Jf���c{�fk�����b�
�?M��^>�"�$����-ݝ���$5S��3!�a�366������~��V������q�Ť��H����==>a���M��@���g�<����?\u�n���(Y*�Z�t���ʔ����9�����c'9Sb}]��/����z$��>y=��[_;��_��)S������y����8X�!��|_~Y68��B���/C��"����=�h��V����:����կz��m��q��`L�(,a�A�T��@v�i?J�KY%����m��kfy5Rco����w	A6i�/�Qv/-��=����q���q,9n���~|MvS�[���K����i�Q��x���u<�)��!K�ntr�9M����xN��������@_3�<��RW��<�V��~=�:v�7�sR���$<���)#N�"��S�O�;��Ɔ��*�*����G<��u�����m߽v"�i�;וi��9'_v��qLg8�J�8�>7_�I+�^���*���i"��I�»I����P��* �ZG�o"=�t��URv��ڝ_K�{f��2f�����WJ\��{Ƀ3})�%�wv�݋31��#8���+�O�R���o-H��9Z��
ډt�q/}���Y��یts� :�8r����v�����Uhʡ��s�1m���)�ռ[�t[�96�E[!�@�ܺ"5aث�M�)�0���Q*�M5�f�mWt�m���"�T�Uci��@�#'З[{|O�Z�|Xqy^��ݲ�����j�o�z�7��J���k�R5�.��������_�ۑ�5��1���ܒ4���R��Gu��m���!��OUe��fDr���V���l�2����Ď�:�$L���Q��mǲ#.�*�n�y;�B�nG����#'��յ@�HW�$� ��P:�����v���Þꑪ��|8����w�cfT����w%�56������"�爹����>[���?�A`k�h��q�iWA���6���K/'��Ev>��ɍ��A��b9�̾�����)�;��i��N��{{TS��gps{��i��,�qRsv�GW�ᄟ ��;]}[,%Ky��2�z�+y�wx�q"�Y��mf�DPL��[yyv��Pe3Y�w���*T�9*�GW�[��ȯ�+�w�G�����	0SR�1��?z��`���:��'�*g3o6`��'濆�W�Ӽ�y�>��4Qf��XC���$��^˾��M��+N^���n�����;��g�y���,��Ռ�Ȗ&���²�n���d`ۇH�{��n�wD<��Rȵ\��́w���ݲ�i':�Ow]:Ce�`Ȁ��5�93sչq�I	�C���i��f���Z�E#��$ͯ�.��m7u4���=��+&�\d�!c�F��$.�m@�;��yC��{v� �d�ә�ATz�u��cEE	:��{N�Q������Q'ԝ#�#'j�U��WQ����o���rۋ�9��T^�d#0�ҍx7A4J��S����N�;	��r&��إۂ��FW�S.��x��dˉ������	����y
���rMCx$r����N������:2�4e�S뫔o�d9��<3`�9��u��qTʪ}�:��u
�Ñ�#�/���5a�Gz�\�K��7K��ζB�����Z����q�#���V�[���*�ʈ���Ȝ����_�h0M�G�ucm<m���\��ҵ���"���7е��:^�?d�G���i��}p�}���;�Z�-�`UF�Gg�O6��N�v���2�{VR�r�'�mp���\wн:�k���<�`��r2��/כ�5�3+�I�o��je�ݦ�b3`���:���JP��Z�w�3�gۙ]C#�W�}ZOt��;A����	�x&���Y]����ີ�ۙ��=�u�UŎ�&:A�3��ogd�����S��݌aO�)��?�z#l�QJ��������Ow3Q(�����s{6���n5n��ͱ�}���(���V��;�cٖ^}�H[�����ƣ�h����l�G-���s:,�!FݣS5u�\ �&��i�syy�7s���$q2Fxpk��`(s� ���N�����o��=� xWz*�����I��
/�B"����<��9�BQ�dY�f�`Y�fE�FB�V`Y�f�FdY�fQ�B�eY�fQ�V`Y�fE�dY�fE�V`Y�fE�FdY�d Y�f�eY�fQ�VeY�d Y�f�``Y�f�`YFe�f�VdY�f�FdXi�fQ�dY�fU�`Y�fA�fQ�`Y�fE�aY�fE�Ff�`Y�f�VaY�f�G����80̋2���"�0,ʳ"̣2,23�0,ȳ�2��3
�(O��aY�f�eY�f��dY�fE�`Y�f &�FA�F``Y�f�F`Y�f��e�fE�F`Y�fU�dXaF`�fE�d�f� �eaRdY�f�dY�fQ�VdY�a�&E�@DBVR B��0���(�(�(ʈ�(ȃ��_\s�*���0 0��� � � Ȫ�*���<�  C
� *�0 2��� ʪ�*���>�����  C*�*�2��ʁ����"���(�"��
��!�,0,0p���0Ȱ������ʰ�2,��̃2,��(�0������������ ��
��
̟����~Ϸ���A�_���S��>#��c����g��?��������O����{���@� �������������� ���?�?Q�G�p��I���I�p�_��@{��p�i��rC������?��@�B}z~���~6+����B��** L��,�� �H�2*(H�#�B��2*(Ȉ��J��� �J��(��H��RUE���"�����~I�� �-
�H�_�~������~?�(>����|���*���?o��z������=��	�_��g�O��O�� ���C�C����y���Q@~���C�!�?x~��=���zD~p~��Q@|'��)�����x��`���o��z��'�����8A��8��*�s���������>=* 
��}?#�����~��������Cם���$����c�2T@|>�������_����{��h|�&__�c�`����~���_@u>��O��Q U�O���o��L�������K�ry��A_�>�0}ߏJ �����>��~�������e5��NI U�� ?�s2}p$S�<z!B� U��@U��AUU�h�
IP��
AI*
BQJ���QUP"��@�"����%���Qe�����	UT�Mm�%F���5�XU֩P���1EM��T�ƚҍ�%��fc�K�R�9MR)j���Cjզ��
T*�*�	���% kD�H�M��E2��U�mHR[2�V�k[4�Q�c�T�**�ka+Z�	���Q2Y���  n�ﮅ{�l�:��s�Z�/kn�����*iY[gu*�ڪ�Z�ӥ��v�kN��:{r�{e:��[[�Ӧ���M�U(Q��hR�M�ٕ*m�V�W�  �ǡBC衡C�c��WE
(P�G��9(P��D�
�_p�(t5=�VO���������=mu�w�ܽn�SJ�hK��wv�+�tn�w��(�R����aE
�յ�Jem��  �����޺�CJ�r�����N����֚��v�F�R��4w;ow{m�:��YM`mf����j�v�i�U5�������vu�'����Rh����I�-_   l�T}ҝ ��s�i�ە8j��mT/���^�pzS��m�{��tگn�hV�� i����T �s�'�sU(�1�=a��kT(�cBT���   ;<J��1����ʰU�1��m�ڪ�v�uF�mP M��vƚӸ����VĩS������S�  �a���h؃+�S�m��j��'Gv�0jV�YO�"�X�����vw (��KUU�V��+`�"�IMhѡ����|   Ǻ�I�۔U ��F���4b�!UbX���  lw v��v �@� �r0  �ET%$�lSZ
���+�  �| >��0�:w(� ���{ <5w JwRn�����+  SK�@�f`@���N�.��j�M�M�[56m�m���  <  5A� 9, s�p  ��P(5Р(�n��ҕt�  �`@t'W� J�䪶ҕ6҂T(kE	�>   ��� y�mp� s�  ���[z����{{� =:-�
t �ը:�gy8��z3��
@*c� : > E? 2��@4@��a%%R4#Mh5O�x�UI��� a)� ����`4�M� �T ` &T�3*�  b~���~�������؏��Z,�Q�F�V�,�1�iD]~ٟ'���{W�N	�� ����N���?�cm�`����`�� �����m�`6��������T?���д�t�á�Ӳ�R`	��Hm���ZJV�j5�)�N
�i�zS9R���4���K�( o)W�Z�7
T]M[h<8�� �z�9Z��l��J^p�&Ԭ˕b�N� d�+-(ؙE��ϋ22�&�PYz�d��F���-�D���ފ�X�N��\����} oV����dt]���,6QSjlm-��\�o[������Ynn6���m%��ܴ�Yyw"���22]�sv=�����$H=5wf�a�IX��1K3�0�"�tN��i�g]
[����[ͣ�/l�t��AM��� B���$H�ǔ�����iw,H�a9N=m]�B�d�m
��w���	�ճ0oƥ;�U�i�5��¬H��Pɔ���T�r9O��ۚ��KNR�����������OE!��̺WX�E�"�Y��j�ֶ5E0j����Y����cDA	�w~ ���J�A����J�Y���-J5�)%Ap�bV�@QZ]5�1��7S`�����%��nSQHE�8lҌɉl�n���^�/r	&]�
8%, ^(��B����N�\hm��P�̩5Lf��48UcRlj�sd��W��٢Y��m�P�x��%�]4����rR;�h�e���x�NY��^ �n���H��\Y���u��cr�)K)\�����Qk��Nh�yM�#�T�6c�K^"D
���e'�[�{t��nM�v�f�L��PפӅ�l�Xe=��)��V�i[���K���頕k��ҬC*��@��K�*��)CzF�˷ki�8�t�/)̀����n�P�kh�̠�&���f���n�9����{��GBs=�C�Hc�ï���%cB�}V���̘*�E%*��Z��2]��H�Řu�����Ji�B5��r���2ͷ�a��cQ�UZ2vbVv�@�L�Tp-Y2EA|oY��ʕa\֔�w�{�Rn�Z6�ع��lR�
�~ ^Y		��J��K�t���Łϐ�6|wd[y��ҭ0S켲VnAYJ�9Y�<�2QˊҖ�Z�Suj1���Ac�FK�y4����r���[3\U��V�-�����w�B�ـ}����B�D�\�7lG��7@��(t�7p)��i�b9N��(���En:X����
b8����� �4ަ>a�d╻vm�T K�^tŭ%(L`�J�<V�C6�*
 (��f�H�6�^'7��ʃ$�Yv���YgF�܎�V��Pa�U޽�2
�����;p�N�gVY���Q%[�.�N#�b*9b��G姌S��i|�t�Ȅ��bn������Ы�IwN�����c`A��k!KU=�P3�A��&D�Hhą^찚A�#2��WK��Mˉ�^�B��JU�sS�m5���s3�j�G{��N^�U�Yo4řYc*�ڴcɬӵ	6��1c;��3
��b���1Rf�{�5%�%[�U�jIJ��oa�WiYkc��X0�ue�-+�'a�7�&�lbzvZ(�)m��b����2�d��S��;�+�H5
cg�^\�FԂ`�����Ջ�E�3i�ۻ�E��=�`Bڦ�[W��n�s�6-�@�$9�3nf̫�N���V�j��V���׏F����`��:hXAֺr
�r��
�lb�DvK9n�Lh֕��F�0��-�)RYH1e�n�@ۦ�,�����ŕp2�ӊ�X�d×Yk^�E��jA���lH�ۻ*ֽl�s[[#��2��MS\�~�EJ�Lm2��b�wYb���ck6�V�2�8��t����� ൖȔ>�H�ؾ�V�G5%m	2Z�z+hD�~f�i�Ô�
<�T @;we6V�zLxQ�	cf�0x�ӡ�/� 9���'��S���dTS�l�G��C�� -4^�e�˼�4\���@�(I���D'>ݐFՅ��֬�2rK�#�<��u����@��N�Vm�R8y� �G�0ȻDh(i'0bk(�U�@�́Q<_:|pL���5�\���Ф���jF�-ص���ɉ=�9*蛏CҖŎ戱���u�\��%Su�꧶Eb�L��͹6�w0��r�!�U�ld �U�Xӥ��&�a��u�ڟMvQۨ��ܷCYw@��Z1^m:V�kMh�Z�֮���Eŕ�2�H:B�^+�o*�V(c��n��Z����0�Ⱦ��B��唴�����+���sbya�1=�>/)֋���4�'�`XbZU�h&��:���6��qP�iX�7]��&�{�ů�K��eC0L,�<ۥo�K�(Z�*�;b����Xj���+T_���Q�+)�t��mJ�(��Wa`u����X���5�enL�Gr事nGE�Y���ޒ^�� eK�43�b�,�w9�Q��Nދ
����| J�UC���z)
����aV�F2�em�X$[V�Kf�)nR���̻��nKf�X��=��Lw���2���t�p�@mҺ�h���A��r�3JU�ZH�4 ܇5�I*��1��f$�;vʽ�Q`-a�`�n�Z��jЧ���X��A	g,LC
��nf�	,���i�Ҟ��`���ŀ�m=`�Lf����K��dZ��w�M�/0"v	�k`��6��Tҹ��$�:Z�^`$F֢N��R
.ѧw��4`Y��?2��dAs&���9Q	j��I;��h�T�Uy�wh�]���R7/P���k3r������ � f����3�8,�!��a���g)��[2kEm��ꩱVE����T��
�	����-��H�d�b`���#�KR:M,��>�kژ�H��ݣ����Ly���J�r�{n�	u�UƮ�E>pmZ۱���4�c��X1d�DnX�K�yM��L�ͨ)�p}���W����DTL#x�p+]f�c�l�l����Yf��{z!YG
��.k 
!��X; ���N�n��Ni*S���ۥ`��0��4v�('[�^k��L�,� ��v����.��E�a��A�Gl�VH�ug[�~X)�I�n��б�.�@&X�h^����h,����1�o-���C)�y��(3&e&�J�ЇY���2�9*a���J�7Cq��uR|�� �m����p���̭��n2ЗZ���Y-�o)��VmmՕ@kҘbܰ�(���L7R�Ȳ�4 Xȭ���̼8֩�-a��1���R�Dj���NN�	��L�n�)�Z&:lU�l��$S+��T��F����1k�(�3)-ݲ���1����T):�����3w%K6U�4��-����iR�C�f���+1D��[�i�m=�-��%T�R���齔U���H�жP����B'{z�2����vkV�.�:�%���@�Ût�ܤ�4��zn�m[m������2U�A23i`����7(&�9B��V�eM1k�#2W� ;n�,4�d����޶�-n��P�Q�Ȭ�#rXˍT;`��@����U�oV
Isv�ۭ��f��<�QV�(��d�R���J��	VY�(���n݊-�Nd�P�8��n��gJ>D'���#q����7�nϤofKl�u�n��6��U:��I��)�䭦�F��JU��cZs�]6�C\8���@P�w�n*?�b(�i���9�&�2I�
3�`���giҢ�])�2�EXUո[�t�;B�l�]�:GZ����;����fQ8�M����h*���7�Nj[�(�Լ�N���p�6+q��	��F��"���bw��0J{3f1��/
#*;�ʻʸ��2Lj5���-��%J��,`jB�h��(��f0D ݑ��U��q�s4�^۲��dZp��I��h=
�٨�oc�5��ܣH50�x�8�"�lV�Z��^�.�#0F�*����A�1�H5��+�j�p��l�1�K¥n�8�ix��ݟ��ilMUn֧��zK-T� ���-����2�Ɉ��wX����EdT4��K�Y�L���Ah�r5��֪�
k,J���:��r��Xa=!Z��v�a�2[1�̍����CJ!nJ�Z��Q���%F�5�o��v�t[R�LM�1m6��wXӎ9��e#M��+C���r[ڸ�4� J�'P���&�%4l�u��R=2+��\L|6������$��ؼ[������Y[�a*ڑ�@-u�F� k��dG,�z�CyKVJ�(SA޳��T�D��PԬ�^��	�cᥚ�ɪ�9@0�m�ȍ�Mj�-�]7 �h�Â
v ��KF_�nL���ATY��F90�L͜������ �ٛ�.V���{����Ⱦ�b�ql9e6���
K[Xb9�)R�V͐Vc8�� ĵ+	��i��B�
c]����.�m ^t%M��^���I�S5�X)�OPj�[K*����+%��L%v�]e�8ݤ��n�	A�P"��X�`�׭!1S%�¸[9!ڐ�X��H����U��Y�U���Z���`��1�7#��J�ܵ,�Ȣ��T!J[z��NV:i��#��"��=��(Ep=�Dem^�ia��9���J^���W.�P#V��V�-n�\-�G5�K,�fM���xm��h�Xا ��0	D�x2�: D��n�*�*44���ƍ2���VM�����V�Q�F���F2Kb���m�Ļ��թ��A:�
nc3��_l.vp����ܬ�ۨ�:"�	��j��k"˳��O>AY,l��$CHRշ7*-����*-�yL�w�^lm�E�-*�Ov��M��tw���*���tv2�iaM3%(�v��۔3+2$VA%V��ˌ�5c�+A6~uH���T��S,�,��.���CR(c�s�p����6��X�MsGťL3Kϒ�&�rMYz�z�n
N6^���3P'M��X��h��p�ŻH*u�b�f�u(�w�*h1`z�'����Z�r��Q�f"�����SYL��-q��8�pi1�T��u��������.L�5��q��^4�b��Wi;S&����-��/rI�ۉ��4�.hw%9����Ɇ�qI>,'[Co���-&w
bG�p��:]�T�*f������RJ�]*���
�X���Q�&��*�M(R8�:��ؘq
3v%&\�Լ�S�/F�E�ӫM�ж%y�0��yr师��P�P]+KZ@�4��Zj����J�/m���M�w5V���N���F�+��q^� �lԫ�2�-QlKf3'��Y9��FQ�uy6ث�b�f��KH�tt/]�`>@���	Ct`��Ƙͫ���sZ��Bb5�y)^��e#[ʃjM�U;dV���m��^�7,ɻ�fK��1�B�۫��m��RY������9z�YY��6E4a/#�f���	p�*e-h���V�Ы{�Ĩ�r�K9�
����J�n�v"`SVm'X��-Y��VJ�R��a�M�n;��ӈӭ5�R8r`ڕ��1�
[2�H��1JXko3e��c/h��ro4hw�4�f��X��b��l9��kMnQÆ+��`8�Xg��Y���t`6�ݘ�9AH�t5KQFj�Ǹ,�q�u����X�ɷ6Y�5��6��SD�6��[z(��nR%"R��݈*.h�opM6�,��wɟc���X����4�uwGU�%LdYt3#o(lu��7�e��(
oD��v���-[y���W���x���VC)�9Z������,۬�E���6�V*�m�cZu����]�Pm�E�����q�`詴�I��ѻVki�4p��mb�V���KHt�$�J�[�y ´�w"*tq��D�t�[l"�dPhW$�tM4��聂0 Էhޅ��v��k%�{�l��*ӻJ� 3@�#��wt�ԳF�8n�d�/TqaN��C�<}�d1K�5��D#�f'b\>��#�L[P���D֦򦉢�~)�z�ɸ$q�	�-�62j�+B��R�(�U,�ʵ�p�E�� ���Y�EW�ѡ+S(`d�8C����G*�u��N����	L�������%"�0�B	�{2�J`��[n�n���Xf�_ncZ#��*T��d�T�����5<����j �2�pP�`���q�v7�$$��kZPuALד	=��A+���m1y*8�2%EW1}��۵�̙1á'fYv~8�^��'Z�wJi�,1J�^IP�sb�S�EX�䂈�@�;��j�3o�VisDiPMj�4MZ�3kl���A�XÅ��Ĳ�ͻQ)��KY�ґ��nm�5�v�W��M�&�r�M�m�q�%���̐=so^JY�eucr�c�©L|N�^R��w���+s&+$D2�^�.�8�##�����{�V�&6S Enb�nc�&�kQ&%X�j�S6�`g�:�z13�1�àC�ʽ�5e``S�{j��|��Sc��R�R����� ~n�"��X�0�'���ˡ1�A��]�u�W��7jT&^g7q;�κ�`�ӒB�Ѷ��ѭk��WwgEI���2*Ҡ����!+���m�q��[�����"vM�۸`��У��{���^h�{R�q�+�V_^�^��I��.IR�S8-�K��eq��Z���Z��B�*ڱ7niL�i��d���x4�t���y�yF4�_��9�ج�݌��Pj���T����t��*3D+mS�[M�T.M���{O�F�F���y���G���[R	�s-'z�;R!Rn;�c?���!f���%tX�uq����}�[� P3�u��ƥ!��������;KyT�oR�ܞN����[���
೦>J.�9\e.S�L�0�;�M̪)i0���YH�i��YK'}�S7W�)2�I����r�m�KG|@b����Y�e:d {x�DP)N�).��MN��ak��K��JK�n]�l�]��P׹JreTI�q�c�
�̿��i]j�oQ�ֵ�2�]ַ{y=7����pV.����͌
&Ysz�,ɺ(�O�4�7a��v�fM�m�K̛�v@�{Y��ZZe\�2���bo���E�Wol��l.�x�l��I|��WmvG�[��ˍ��^�\	=uҜ:g12&�w*/�e���w�8:�^eN��A�F^�cgG�*٫k$�l��,٠�Ƴ�]�#���5�sbd+q��ą�Ȳ��=��ө��9�H
���h���M���=���v4��(��������Ǌ�;
iY��v�Ϣ&&�,����|�eȸ�멏��&L��R;yݾ6f�w�>�
�pl�p��� ¦�9T��¬E:-q��6@n��p8-�(	K��%t�R���X�V�}�z>�eG��K�'H�۽��pYYhgS<�J��dc.�����h��\���0��X-3ǯ1� �޾��|tl��Y{:qȭ�4��
+w#�m��5�o��2��V�]�d��z�U�:'}�1>�Mc=@h7�R.I��:f�W>�3E�0��'N�$<��g\�Z��aS�ܹك�ɫ�ר�T,��c��}�Ȋ�c��u��e�ՃT9yɬl��t��BbU�N�r����]̮�_uZ�Q}��vW]D���3�����'����_�H>S\x  ήw��Z�^��.t6�����d\��y�\u���*�:������n�Z4�g1��xI���te-٧�)GkE[r�[�����m[�B;��3f�X�z�Ek=�%@��et������k���V#W{ͯ�fL�d��/V��ln!"�EN�ֳwi�|/R��"�|�w��ye �K�cݬ6%���ۋrmѼ k��knf_k�2r����/��oj9MQ[N��K�?`P��1��d�P�c�\�����%�r��is��m$s�u�E��EV�=}�`9-<�S�4i��i
׭Wp)��5�۷�%�J-���!���{-ۖ��.�t�\�BcO
�-47���|��xLd\6��]j��M��(:�[��Gpŕu��Қ�ŻKPÉ�]�F�cV*�F�i���t�:��ba¢���i@�����wS�k�����Up��k��坖"�+1"2������(a�LJK��кth,��!�S �u��[�ktc�,A���Y�� w���<�N�k�u�݃�ˬ^�wS����*ܙ�>�����"\��R���Z%�|�p���yE�
8��tK�9����Y�Ax�����V*�!�k�ם�a�|��`���,�[��1]��\}�O�_3r�͇[���p������ޞ�K&�#I�X�,���噜j�t�����=���Z�V�48�C�c�jL�r�.�Z2����|Q��1����w���;���K��l*�*�=��Yê�G���]D���F�ֈE��T>
��{�U�"��d0d�,1YN�P&�9�Go��u3㊸�ҍ�*뮉�8y:	l$4#81Ї�%]�)�/<�4���<����Y�Sh<�w����ŕ�b�t2'%��]C(^b��6���q���}qQ3�W#�m��;������y��(I�o)b&,��L��]������ၧr�~x�
��gP��
s�;�J�ʮ�Mn��z�X�����Ѡ2�$2'tp�q�
N��޵�T�ӕ2�R��)�7�.'�Ws�װbp�-������9X�cV�
��ƫ��f_G�,� Nskr�C��y&���8�eZ��V������x��Sm6p�F�0��[�萮ڇ ��6�<�d�YA�r�f��cK�����S��r�:˥Ī��J��y��=���e����bS�js��:�x^rU4Ӿݓ�3�����n�8Z�C�|�!�v{�L�n����P��"����.���ԺoЗܭF�D��\ͣ�u2�쇬Va#��ST�c-�`��oq�'d���m�,_Gs�/5Y��u2Z�����h��]n�k���(�{���-�Y��c��kmf�k.�c�oڹ��6*S=A46-�o���p�U�`4HgG��iA�q�l���&�s�"�^��*!ʚ?c}c{"=��u���L����V�Y��+ ��-�([��tn'�;���&�N�����,Asz�"&D��>�rg�JW���*���r����/j6e��8Q����v�[��0�\q�o^c}¢�e������FUq���+1�<�,�xk�i�>�5�"
\�zh=fc89o<���=cnV1_8�=��u�М����D��R*�!�-�4��^�s�Cq���� 0+��|DW������(�	��m�xFU+�7�}	 ���q]���ܱz�g�>z'�#
�:��GR����XV]���],Q�T����
�v�;Rs6墸9^,����Ҿ�L �PUQoZb���Lpq~��"r��稽#eB�Q�@zk�b5���CZѷ�Y����+b��S���-��=�ECa^�N��c{��4��' 4T�Nu�p�S.�[�uC��c��|:���+կ��_�`{SV�y�Y�wGwK��5ol�Hԋ����e�N�dV/���X�� J��P���OX]��U�#^_+F��6��Z��+��#���̼�N�:�e�
�|e��8[��]�ֻ�O��n�����)y`����sc霞f%D���2jz��U�ス��,�Yj�,��*��Nk1���-�PoodwsqR���gQ�����z��/+�̍5`���I#!�(�P�S����A�|:��jlH(Q�%uk�u�ow^-��!Io&3>QR���o02�V��w3�
��ұ�]�mڐ�[N���G����У��r[y��C&����;��u����,C�I�ǅ�N�em��p���3��sNIc�ۇ����,�'8'��CK�u�م�1�.�:T.���&c0�
=?*����K�(R�ӡ�y���MgT�qn@�aW.�C��f�h�x36n(b�#���L+\0�FQ'�+x��Eȋ.���sk�Q��\�e��{]�7�D�޻��V<
�붓��lO"��_H1���wTs^���NkYլ2,�ޤ��E%N����[�bsv�w��G�J��G�B����������H�	�^�=����P늮��>|�T�D��[�31�[�r�����amnrD�O\
� W��},�Z&�,hT��ٕ�:�lJNi�[��c����6�z'��[F�*�Y�$:���ܫ����s��مS�,��4̥��C�(��AM��Si*[qaӽC� �w\�o<k1�9gI�l���Cp���swz�k���R��OM�uQ�u�q_n}d�'N���E��̄YtF#�Le�]q����}�� ��F#��/xDk8�={�wƝW'��Φ�^ڧp,.s�I�z���vJt��e�Y��'�Zj�)7�,F*������o�~��Z%���Ol�|�37�W%=�o��+�;-��yX�-�5�T��!�d�+���R��+����,e-��M��-�+q-a�Ϳ=y|���N�kp�֌$��	)=�$Wc���N��Je$7�"B:QR��`�l�7�	GB���1ܳu>�=����z���v 	gx1�&��Xyu`�qs�4N\oU��ژg�G� !�N�C���eQ{���i�Qy�߹M���3���{�i����8�����mhg#8�C]7MϷ�ZI�6�q��ʐQ�n��[�R��DQ�ڙW=��osԛu��l���}d�XM1g�f�S��2sU1F��WucE8��9��뜞��a����m��mP��Jnu<{�K��W�yņh.��-�[��p�).�*m�:v��:�%�]����)R���k���n*��$o{�`!մ���f��hn�.�#CP�<��)�8���/GAG�{e�����ì|�Kv<+7�q���W`�'#݊#f�cffQ[b�Q�g Q�g�&�4A*a���w,���ۣ�g'۴hre�*Q�Mf��[�j��^�'�t����%�nD���d��]�n�\��
�z��ә���Z�\`
��7�~�E���ڷ�e�i�v�z�b����0����zT�v�U��/�X�q^�0VZ:�@Ӏ����Q�>�h�hrk;6��[M�l<�*:Mb)8u�����p��Y�]�*�k��R�4u6U����ϕ�-V�V�n�ev���d��&��YM�w��[�:�Õ��E��2���N�*��5�]/T]o6���N��i�.м(Ζ�p�T�8����3{��Q���{����Zܨ�͏x�S�V���KXV�	xo�@�a�i�Z'�M��m[��|�8m��ܺ1���m)V��=���6��^'�V)��AY%�u�8k�\(z�9{mڜ@�"��?	\@��8A�9be�Z3��w|	�1���eN״�Bz��}rq~|w+P�u�Ϊ\Ul㲧L��Ӭ��v%�N;g]a�[���v�3-uv�������A,�쓶{0��Xf_�hpB�VvPQk�Hbe�lb!atk�7�)���ovd�c�Mt)�=�/w�F�t�SN�*�"��n���F�v��mD>v�,f�,���]�;M�"��?������D3s�u��XdH���<�m+��W`��+��ĭ7�x6�<�^@��(��a�VQ�������ݗy.���[�*"��e��i�;n��ܫ�`����q~�c����y=]"��;������pж�'m�jv��/x΢Yά��7�F�:n��ih�wE?g������N��vf�#w�s�4u4����5ղ�:�7d�`�W.]�nbu��/�;Rk�ko�������B�Q���A�X+{C/t��1n3bN��=r��6�kx-�&�)�h�j���<����ٌ��ݐ���u8���Nn=��m� 7���ӠGs�)C6���䃘дoPz�B�_n=y���8o��A��n��d���qU�h'���ű�}g�Z�i���@`E��#�+��̊΁|�P�#�Feխ�)b��p��:6�Ր9�,vV���t\ؾy*����Rܘ�+P��{�@�<=����]�wx�2�$ �{x�ծL=h��
m�L�����x�|�Zdr_d��m=%��y;��ɚӼ��~
��l]�)��l���\����N!A�0�#'��'v���S��=�ڇ-t��	,A��w70���b�<לb�r��>��7i'o�&]�ǈ�X9��R�gcĩ�U�Y��B��ۚ�\I���',n����v�n�@��60g�>L�Bo��A���	���|�N1����W�3�kI?C�F��,��z�h����D��nV9)�t�k����F�vL�b.;1��%9�:�s�pR���G�X�\��x�.�&ޘp�F�3mc���W.�6e5K�r��c�J[��Y�m��(eL�tx��z���+��T�W-�f���U�"�ʟ\+{$�S���rN�����{�J����a{8W_����!r��D=��	�6�!t�R�;;탺�������4�� ��q֥J�;ݒ�\u�(�w<iŦ��tu\���i-wvP{�5��F�$]�-uo����������&-�:%��mCH!/8,-����vZr��ʶ�R�>/Y<�=��d���k���0(S�Ѥ��nm�	v-�d��X�%��v�:�v{��L�jR�[���e�����w`:.�N{{�P�]�q]�W��ɨ�`>L�r�If�nb���xW\{����,��S$�f;���M��,!�^��Z�+�J$�����{h�|\��v�3Y�KtXC/GP�Vz����Ҩ�ɻ�m�&�"�(a#�Q쓴=�Dt�w�:���Qnֶ�]�����/iaMC�FȠ����voI��[��e����>����D�eq�NY��ˬ�Wz^�`Ȣ�{�յ��<�(�ΜO����%�+v�}��#E~����&|n���b�>�{b/I�tVGo7@/�ΐ�(��+�맆��1�a��Gt����8�\M����I�J��c���K�}dTө�9s�������k맂�}ձ�6s�X~FgK:2������AR��SF�mUh���vN*�M�=�AWpy��z�[m�6r��
L�	��9�N�G*�vs��}�����IfU�V2���`jV���w�+��!��N[L���"�ŝ=l�I��na\��[�c��:=i;��jܩ�e�u�e\�T¹�[����YëQ�o	�*T���7���]�xwQG���z�h<N���K�{!'�[�7צV����NJ�Ǯ!(N���^]��,���5yY�@lq̻�����]��0;̴��)7��5d7.�r���DS�_�>3�goy�W7h�r��r���V:��{��EnN�C3�M�����:�D�EgksU)�=���o�'zȁ�����T�zg��e9y8��%����̘�w��8��Mv�"�!Wl��0���k�x��gR��O��*��=�.�	ۆ�P>�mlCG�ʽ�Ds��9ۍta7_�=;l�c���mu�뺑�wk��gt�W�޷��� >��|?_| W���)�],bi�e��"N��:�gt�y;7�	t��ŉ$�v�rTwyXp�Xܬ�5܊α]��k�6E3���%Ӯ�Vˑ˥ZO{X]�msU/,Ty�W ��?��������:�0��vФ�a��k)��\��>����r�3�ξ��k��Dh�d\�:3-�h���L�"�9͓����˫�����;o4��x*c�k��RCq_1��L]j����z���7�̕f�c��Z=N�<��Zn��ܭ�U��;m��/�讎��s����%����a�c��J��aki%Y�B��:ˎm�`�ڜVn�/eD4g�͌喵Ѧ�*��#;ِӬO�zS&��ܼյ�Q�%qv����l��7�W��]#&���:q�~S�,b`��*���$e9Íu�����<y<)=���9�-��6�`[Y�b�dwHn����2J]Lѫܷ6���S��Y�!�4���v.�B�_us�a�a�g������R�Oqa sU��5�,�B�õ�hҼ�C"�����e�q����I��h��{;Rɶ�Q^�Χ;J�W�-��/.]~G-b�N	7uI_��.���
�PB��_Qk�{#����=�P�m�����:P2FZ��G-}7m�8r���թ�݆�Չ"���t�#{�OV�M�Ra���o5sE��1�-�Mǂ�w�e ���Z&\j:δ��_I�o�S�՚h�Y���N��G���/Da��M��'WT�U���t�{��BW)����s7�EZ��8f�3���D����{�ɝ���U�:a��	\�������w���m���ʥ=�kp1�%˲��R�OE��`D-^��Q\q*���u|.n�i��%�JZsmղ隴�S�e+*�MT~�j��\\F.�wg_n�U���ȵ_;lV�����򻮓�g��L�[�b�ܾ;N�[�.&4�����U"�[�n���@j�q��(�]��|�\0ή���v�X��/J��B�a\`���ڮ�մ�����)���8�K�AӚŽe�hUL�ܸ��YR��]^L�Q�6���Ԫ/�ۊ�wfӻ��q!��4�
�����>A�P��A�V��6om��M��ְ��皨*���Y=)q��Fa���v���:�qh���rSf]��md\�.���{q� ,u�	<��j���G��py���{8sN����U��UF�,e�3t
a�����'ݍ��<,���z�N�a��ɘt���=J�o����Ewm���V�)i��:1���{]�s��oz�V/�A��G��%�����=�б6H�*V��p�(\6���ǲdʚ㧁'F�� %�ũE�Pn�Z��,K����M;@d�G�0Φ.�zm���ʕ}���12�1۲
��>z\yC	����C,�;y,YP���̣�Ժ���0]�aRN��%hW>�"�u�q˺RŴ��Y�u��y�n^�Skl��Woiv9�=G�t��v7�G݈Zή},r.�r��t�n��4����e=�Ms��(�ܺx�k[a��|��pWr�S��oD�Zy���̶���C��i�ƱWi�m̘���|�Y��6�GP��P�T�&(����+	�Uw2�1��P��gm]���Ϻ�,Č�xW:O�!�ކ��oXAf^���R*����p48�xp��5s/t�h_)������b{Ɋ��y����՛���+6���
��8+�}e��嬋���#@O*g�n��i��vd�ֆ��(h�v^���"9�����:�Q*�!}��Y��Шl5� �q%�K�a����%�f�J:����wm�җ��R��'V� (5]S�]7���wc���+^��\pNdQ����c���3��LVn���؝(_$�|���::���"C�	����]hΤ�yH�lz���&��M�8��0X�B��q {���*Q}�����J�DxW]����ĥK��8gS܈]�v��h���Elg���*�S��Ѣ�7�%s�5��*4o���HfҾ���3���$C���ܚ��v��N��*`�*��c�ޣ[1/��9BTi-�G&�p&�Ls��81�r��R��w�D��oyi�
i�t��\�Ѥ�&YWI�t��u�K͗/�v�L��k7��[>5������_����p�1ۂ���nc�}o�h�FЙ���%ŐP�ej�q�P��y3V�x��b�"�t����e��_h˚�j�΅�pƛb;���/��h�d;�#�Bwp�5�l�7Uލ=����-��nUؓg���'cMZ�1x ��>��&dR���`�J�5��4����G�u`�9�m�M�}�ݝ�1,��	���X��0�"�m�	���RN�i<��j�0ʉ�q�c��ʤ`\���;+)aĔ8��ZE?�z*X���=��SV�=��w)��2� �0V��wsf�rٺ�6��r��z����U.&������rX�����l��=ʸV^��t�C�����R�F�-f^E���9��&�6\C5%ǩ��.]'1:�'
[��|����t�5�Y���7�2k��}6��JAY�f��#��HS��5�s�#d�n�|��n���(!�
��p��=N��/�K7��Yڿ��+jDa������l�km����� ��{�*�έռڹ��h�b���e�2���� ��y4�Zj��ma&�\\��t] _*l$�j��
=p}74�Z�sFɽ�3שD6�&�`��̉�_[�
�n��g�.���^���8Wס?�<o�a�f�	X:>Y$�����Y'K��;��j�oPp��P�!f�9E]v���H�x��4�&NUl͡��Q�U���ם��t�ї-���NN�l����n�C-�uY�r����%�ͅ�.W��*�{{�J�T�
���][��c�k6��*7��^�e��픎��Tө�������gvY�Ni�+����Qե�tm0nYv�iޜ��ۜR����i">I����Q��Q",��6�*�iW1�7f��%\���ܜf]n]G�lU/+T��$F�X�7���::4�G�����Y�h:���`Vet�����.EXq�`�:&4ZOâm1gpm'L�)�R`5m�00��/s05k����2	҉�㝅G])��(}�u-���8�"�4�f�����|(1��;q�Q����4qڃ{l=��)A�GRu	]]��>�o�:�OM�/��B����\��1�Y`��\�w/E0p�$]A���,�P���ע<����V;��u�u�V��
�Z%b�H��]+aD���ec�R�vjGaÜ�.o`�VQ('-����Q��Ħt�FlW 3y��Rp��e�^��'6��5�a������)w ���&�m͑V9xw)�'�R)�YΠ������۩K�xmR�:�
(t�eX�ݤG*wd���s��c�r.P̍��N���5���Y��(��v�)(1l2v�S,c�%ܥJ��bF��u�ݎ[t���ٯ��.�FʖPAbkS�F���]�roW36�:�5����*��ܤ�Fst��ʎ֚i54XYRcN�����[�6�ѷ(wK�+Z��SXDtX��Hx
q��݆����8U��e�n��PnG�`'#��U�y`��V��<~`�+��H�*x����9V���o����]� �<�3qD��Yy�κ|�;v�v[�C�l5]�?�&U���7��X资�f�kz��s�{���O\��%���Rm��Z��,-��ʻ��9�4��9a���ۛb��7�]��'Y�Pc(��[ųlv� �l#OS%��M�T�����qzi���A�U���j�u� <l�\�6��!�ͦ�����nt5f�.�S,�9�9�Y�������SS�Hؕ
�ܗS��R4�Yֶ�L�;X��/��BU����١�/fU�v8B\ w6ࣅ���rݣ������u��f7P�{O;n���=�Q�nBLմ�F��u��)0�v��v,#3�B9�ѧZ���`�k&r\c{L�[���க�2�,B�dw����ٕv&�L�]��#� 	)wM�F����΂'E�Fd/��9{ׅh�vəԍ\�w:3���w(�<ᄝ�w��+'���&�sG���ʋ��sbJ>݅�77��t�AE����ݵ�V�]	�Π�2��ܬɘ��RR��2 �-o맫�k1�R�ˮ9�jS/ܠ�[��Y��՘����A6r��kh�RKZe��.�1@��Ȓ�x�� �ؙF�'�Q�{g;1րR�RD��$��c�dI�'w�z����K ��r��G���e�p��R�;���f�+l�1�Wu#�wE��=���&��Ea�,��T�}�Rp����_#+T�'��Z�%�+õlCZ��1۰C��:�)����S��"ˮ� �굤��q�L���#���HE�7��r�ǛrT�5��Eœӌf���_)Sf����E����0�MM�S��(v>��hBE���B�s;����r8y�e+�#��#H����k���VA-zv0�:�Ú�z���˽Ws$���o���5;Y&'��Z��PnŘqށ��h�wY:R_
s2Ph�^`����]=��[����z�#a鴬(�߮t�%b�(M~���s�l�`�>F�Q���FdA9E
uی�Wb�#yj.3㇫Z�H��0�](�8�}�f��yع}/'-�|=�||c�|�MO*��^E+wp�Y�r��1�-,\8p2�'k6C��A�뢶� C�}�HD���s�s�qdN��(i�e	7Y����kѺV�����͡����N������-��LO���ݲ���QYr{޷�3=���#Z�zY/QI�A��{p>&�w�w�Fظt_��=�J��Ogv;z�<�k���_`�Y` ��}m����y>t��n��z!�r���z֠�o�'��BVzјԬ�y+��Z]:F��t�<���FvIQJ�hfݏ�k����X"���%*]q�f��U�5���*�@-�I����s4pd>a2�f��c�i����uh�'�i��t�g]�Ֆ�#�����M�W'Ի;
+a�ǝQ@ƍ�@�QG/~.2r�y9��K�pb�dChAY�L�C-�Wd�ա,��31�7C�.�<�k�R{n¶]t�bù:�u��l/vt�*�d��j�c��d�]���@댏�Α�YpQ�RW�m�N�e�[igb=6up
��(���^��3���e��r9��$a�q�3 �uz�+`)��g��5��,���iN�՘���p�ɷ��Or-�n�X�$�`�G���6�,���3��çowHP��Kv���N��Z����rov/ۅ��Ի�_)�0��N�TMF�5�o�4��u#9ϻP�>����ϻ�f�κ������2�ۜU�x ��å�yAԷu����z�E���y�l�)���^�&]9�Ӄs[G�����Èq9Uؑ�w(d�{w۷�=z��}Ѹ�'_)۔��v1Ѣ�LQ���P���l��R(��ES2�m;MsƲ�*v�t����Ӻ|�YX��0@��k^�B�I�cznb&���AM���s��{c��8���3���V3pWF*���bR|��[�>^��c�KC��QE��׹���QN�#]g�O�����f.��']tk����g$X/��<��k�u�Ӝ,Q����b��턛�$ �#-�RY��M�1WdN
ՠUm,eL��Zh��G��-�W=�n;�\KxLKihzs1p��,�L�Y u�j�y���8N��= �֓�{8}�릔
�wx��ΙD)�9�VA����Z�s%�ݝu�����r�q#1�'koL�v��%��!q��8�lr���,iɮ�#V�xә=&�(!��V*E�Ȼ]�\|�v�ea\�{u��޳�b�*�U��k��x��g� m�9�$��y������<^���(��gޖ��v��������9����o��EZ*R����v���% *(�{�ڻ�W�l0�Nׂ�ǘg]�_Aw����ڗ۬m�Ľݍ����mE�s���[)������텢���-=����@p�R��Fu��%u5u�hU�p�;��9�T�B�N�Q
r����A�kY��uk�n�V���9h�Ar�Vk4�b=�n���*�e�ז��t{I�Y(WZ�v��^�fq�cw��X*L��o���¹.Ʉw](�1٧��gk��h��V�|J�2�~ '�װ%x".��+�iV�Ϸ&���\�,;y��x�e�K���mv�t�f�}�n ����mJ�Y6�v�z����p:����5�"ή.eu�2�YcƮ��-��*���bl��H3����,H����}�V�o,�m�h��ͽB7�����:oxWmi��6��q�z㝼�P]Yr�]��h�uG@xH�����櫷}N�h\�WiP�˃�ݮN\�j�La���\[a��v(�Zd����,��Q�V ��V�#ֺW�����ͮ\����\�w�ǂ�/E�����T[@��C������:3��N��Hc�\�c��E�`ЧG��5�*XTa��yt듵����ŕ}�T��b{v��m�������N������e	0�,���^�i*�ն�u닩]-�a\�Bw��/	u�+�_J��ol��.�øk}����CH=wH��gvB&��z��7��Wޑgw������,��K�y��T���2ޑ���8 ��㖋�P�׹�@��x���|���� |>���}�v-�M�u�^��ے�\�y@H��A��oq^�!�l���Y�JW�Ii�zUu�L;�=������nJ�`	v�q��r2+vg]���&������c���4�#��Y"��5%�cq:�΢TC�o���+��i{���-g	*R*��xcz�����Kp�2��)��;v|JC���td`�����zigU`�ܣ�>F��G0��#�oe��Mh���}�Jo�
)쫇M�s�xxL{
�p�;J�ml���.��8�T��iц1�W������,����.U���p��u��w��Dc�47'��3�"���[�m�uˆ:��o�wui�����j$�|!=�t!��,�}u+����>��su/)�P�D�7�/1�:n�/��l�W��BAN��p8������N���_>�;	���!�h�������ǈ����:yP����LC{NQ���	�5V!eӧ��ܚe�R�
ȸ�<n���zm-�JUէg��Z�J��5�Ĺ����{
d����*�_% ���g�֌��k���	���t���/^O��ZZ��kf���k�޾� ��;��̼��6����>Ǣ�c4>��o������wpEgt�`��<��>�r�V��(��:��u�}G/�%}��{Ed�����B`y�t��{�W��9}�FJ-�����w����P��G3���w(��\�.�.Q�f�V��E<x��+*��(��]:]P�"�PY�(���a��Y���"��E��$�P�ͮ@N\<�u���+��""+E�t�0��\")-)E�*�U�VQp���U�S.bШ���Y'(#�F�'i4�ʠ��BB�QUM�$9PQ�*���Em<�TDQTr�(�u0-�E���Q̚p���Mĝ���%��C�)R��(�RVY			QQ�U0���J�Bs�Qr�)BʦG�.���I�t�w�q�J�E�UGr�Ȉ���9A��Ӹ��5���S�ED��$�Z�3ȅES"�p�Uǈ'���	� ���{od�Y{��.vFf|�҇r�׋�'�VF�3:��F�I��9+#w�IRxj���o3���w�5�z��ӧ�}���w��A!����L_gxxe�&E���c��ya_p�h�{��o������Ѩq�4!Q�_�,����Prlt�t[\�ô��E)vñ��ę�	�����{�F��q��M��,F���i�%r�xV���_sQ�\����!�0�:����DWc����W�f��I�h���V�^�"���iD�W�r2p.p1�l�2`�Ȥ��ݳ�QG�'C'.���K!��J�ϥ�3�]�n��ꬖ�\h�RMI|M7�s�����yѣ�⃫��qS���n���,�~�̜��6yl�₲L�콮|S[���,7����v�,O�TX:�1���[<��9b4:"��+��}՞���G����2�#�� [�Cvck8�Y�۞|t��z��G)�n�#��������]�P���1���+I�GA'je �{]t��Ƽ5�<i3��:��Y�|Gr�Kw����Z\CRY|cD1�o����y �(�( px��g�.]D���7���8zs��ޞ�r:ǭL��ޢj'֞vר�����w��jH�^���4&w@��{[t�9g`�W��T��{����eN$�X���6�W�����b��(�4hӉ��D�¯�����s�N�'(����n>����q��Y���7_����C�8`���i�����ܺ�!D��Dt7��f�s�M���W���� N��EA-��q�"���_(�U��M��5�,a,θ�C���y��U;��=�\2 %���j���Q�/�5	.�'��<L8f0"V����ƺ�k�؝x��n���� q����H�[N��\v���;��Tm�d�7ű=��z��Zko8p�ǠƠ��^�'��q|��;|X�`ɝz=�����/E3�r9�9����4nt<�j�_La'�#ӐrP�Xu�Oa��-�Y�ɹY��gX�����˯.'U����O%��n���<�!.�㪳��8�~�m�z/�y�G�c8*�V��ó�l1o����a��k���������	i��&���n�Į���1��T����rp�3μ+��+��jWjc0�Ox�����v��������BJ���J*�ˣ��t���x��\ ����u��Vvb�w% ZZ�Tz;�6���Ƿ*�Pc�޴���n�1�w ��G;#�)6P�ˋ����Fqb�G�/��3�����!�k�ϸi�8�m2]�%�s�T����c��e�xrTtb���$�K�ڞ�lY���[�!|"�.�F���Y���>��I���9l���V��\K����y.;OUW��>��s��T�,�{{��u8N�X�D�픊퇗�
�c����k�V*E�XS?0[�3B��7i
��Twۇ�ym�&�_+��n`2�S<�ۿ��ơQ�x�8�+�37�ӳ~ŵ���5:��]dE*��wS�xă��������0�M\>«��!	��9Pr�nЗ��ѲM�3�H-�0��]�K�����R��ki�ȳ����z�m�e��N��A�+A�=gW�k�3��I�y���}±>���Ӹ�jr��e�)v���;��O)�Ӂ�TF?7�:�'Z@~����ʫǒ�u�ms��:Ko��ٛG<�����gn3�9�;X����؃*d�+�R7�&xAM�����|ܜ��xu��u��mDs�rn��i���+�6�
�9�v:�SZ���I�;N�sעy[�0R��W��1G�V��Έw�|jLrN���#]�QqZ�����*VU��MriƷ)+�1��4ݘBY��1r�.�j�U�ZN�t����v����΃��C@V�u��6�gH�0�ڜ���;71�x���]aV
�ÖqǄ[ᦱ6��\����5���1%9��t��:yv�q�/I�L��qǵܕ���eEl&
�������XDV�wm+5���a��!q��ȴXf�9`I�s�㏷t��	D&��Nw嗋,yc��WH;���T��!��1�}�����щ�fo���Unl����Y���>X"���*a����7B�st���M`��l�n#6հ^9����Vj����Pш��1j�'����p�`���~�:���Jv�N�'��ۡ�l�
�M����C�W�p�\�2���K��q��P��)^�`A�U^gҸ��6�$)z����&x9`+�mCQO2��t�Xk�f�'z�aXc�]H������9n�gjZ��jC�
��)��O���11������T�_��g��pk��&�\U���v6i��o����B ��?4f�!qS=��Qb�Wbn�d>e����7֤��6������R��u�G�֘�������/�S,���l�6�����>1�M�f�Ӻ�PÆ)��@v���F�Cw;�h��zw�(	�
c�[Uu�&Ŧ�p_u0��6%x����XJ�ؠ�t꺻�"5�[��ˢF�R��f���Г�Y�;<��&K�,ۅ:C;��ޭ���Ș��-�վ�6�2��Xn�<�-��R����˛[���m=rl�'����Qk�}�]K�y��}q����i���s㯵���rsee�:W�+�l���܌�uh���A=i� ���Y�ѓЪh" ���\�|o���p�s8�xo*vٌ��H��f0E|��9+����<y+��'��ڵF[��5�9=�h])�qe�q
x}�˭�2j�9LZ%1?FB�Q+j�C5<�Z2��{T:�P�]L�N�%tY��E�"�4�n��ބxOg�JY-,{�c"� ��Y�6��f��L}z�Uǉ�T
�Q�t�k�7�Ɇ6�6��\����\��[��8�D3���]-�M{��i�����&1p\9�
R�-d��n��jkq&&�n��ek�K�g�Gt���%���@97(��U��ٜ�0�p�7.�!�:�;�D]g��f�^�ru��6V�E�[��0������SUQ=��!F�T�KhW_�r�p�f�딎n��9���$�d��v��Z�c"^�]/�ؼ"���q}<_
,��7��#���f;���m�T�l�� �!"��G�T,p��-ޟ	_s{�/��͈t<é�{�>G�_-껵��pz��޺�t8�:'w}9�A�G���/;_J�sp�;�A<��_�r�'���Vj;�)콝�1�a:��BC�e��igv����ot��|��IB��L�4��L���w}��cp&:��Ζ������R��й���&��oc^2�
�_����Zq�(ِ�/�7$R���3��e��t3�������V���n�\���C%E��-f�ʯ���>�0�ij����i�X{b^��wp��]�r�c� ���&b�Ҧ7>U��@�c>GA'je�T�0ķ��􌐝�܊噤>[@�E�Ƅ�F�o�5%��"�cj�\!eͲ��piA�
\Nh��kk�|�^��?T%T�ϩ���9c����GZ�������u{����a��ڲ���h����� %�{�B+��_1xxc�븛��<sp*���9�ջ/PY���&m�2Ճ� �1������� h��ա���&'l�>s�b��7v�������_����8l�=�G�C����\KfO��5�P�T�*�^�4G���.�n����+� ЄP
e�(���Bdi����W�ѷ'�!E���zZl8����_�V�֚�"�Jd�M�ؙ�,��a����Pb�S��2��",�vXto.,�kѼUD+@��)�ؕ�$R�'&.��3����T4ݻ�k�U�L�vz�J�p���K�i�x��7�%٧S�[[sIk���j7��YU�r�cQ��e�/��m3+�������4��vN�+$�xv��??�c�+ �Zj^\,�N�dk��5%����l��p�����#�=e,�٬�KQ�O�1�h�Â��i1�Pk�l1p�>��\�q��>���.�ZY� ���ZL����\i�wA���
L=:
8v� t^��.�8�F4��$5'�5��ǯ��aH�}�����Ƅ����B�����:�Xi.�;tpm�B6g�.��&Gn�Ll�w����M�ϗL5��Fyl��Ո�'D���+l����z���H��m��}k��-��<��:�K�9�_k���nxF�UtgNI�w�I��x:�3�B"�<sS�܂o{kι}w=s�b�Z��p5���e��q��=>�5����ihr�]�
3�}?e�9�O3')�wh�b�]p���f�(�폭�t�d9���j��X��/W��S���L��L���J���*�����6GK��^�%s^-���k"�����57��F,�F��s��O(�<�k��mgLnŃ�q��#_p��>���N�;v��ET���MFܻ�^�#jR�@k
l�^��u�
n�V�\8�Rniek�a�C�}u�&Tg0�{��<
�5�OP|�y�>���
�\:�n���;n_F�(�"��vnVn�$��=��+�>����aÓ6�����M���&{����<�i #��A���RD.#^�7�	\VU���\g5��~k4q���C���74	���Q� PC�tWb��y�.g&;sF43�f�ٔ�o�%���М�`3L�Ѝ`��"��4fc��N���E��r���d�3Ӂ���*,�Zb�^�\�e�1\��FṊ~5�hּ� 5'�s2>�^ө�ޞ�/je���C9�4,�jr�u�i��]��'U#��Xf�9`I��}qҰV��XٹŴ�|�eH5x����N���\���Bdo[.0Ֆ-*� ��|.�Rr�E{r����'�P��;�S�ƅ;:M�`����^҉�*���W[�&�W�n� �[c:�F�.�!����O\{ۜ"��1�@vUQ��tv����u�/c"�׶eNѳ�+V�����y*k�d�Q�g���������1���Ä�x�JE�=��d]�y'X����?/f-�v\�(<�l��5<�\�yD��	ޣ��a�s���{�������k�=6�9�hq�&��Uw�hL�������샻���kTr�>ڸ �s��rLn�}g��)��ܫ�zn��	�ڌE���f
�1�F�k���ss����(Gu�L��9���P���+�s����t��X�V#��a�K�Gy9/nr���+�?�XxJih�U����6hu��_]�Ri�g��u����q��&ޑ������"�]�q�E]��?r2g�	'��,B����"�z1�U�|��+firv���e�H��vf�ۓ�V�c�3�4�0�	��6�@�LɈe�z��<=LcCU�D,��8|�7��IF6��M�������p$��@�RP�1!#�3M���Ÿ����o��ME��q ��yL��!�Z�~�\����$�[Da֐r�XEr`�`ܭ�O����w���F��Ô�l���H㙌I���ꙑ]�8�x�V�7�q����>} WHq'��Na���,+S��]l!��e�&-�����Cw#a�rR�ڍ��Kեj>�*�٦�"��v�Su����z�ܔ�\k������'R�Z[�"�����(���������טn�*��>��»}������Y��w�Vt�� h�PS�f�Dg�{Þ��|�GE�>k��v��}J�ɑ+���{��yq�<j��Nl���vZ/*XK��0� h8C{B��/_�h}�߰Rj;B�~�2�U��o,)�
�.�o�� ���nXd�:wJ�\8K�sP�!��Rͣ�'�
��h>��XW^��T�u�
.���s�=6�N��"�K�Wd؍��;�9�jt�p2���P��f�b8,tY�N����)�����j=����s'�F��n3����0������V�w�6�4�1`٭(�š�q)�.A�}o��]��vU���t��g�RP�s�Pz�C��WFK�g����8Î���%�λ���3Ǆv��+��P�(��j�po�%-ޟ3��M܅�'N�-�5�]}�{�X�ѻ�i����W�*'s>K����>��-
��mt�|k-�ְV�.z�V������]s�]����XI��f�������P
2��8Uq֥8'������۱�j��4C���1p럆_��掰a4��N4�C�떽��1=�׫VmK��<XLК\��ϡ�,�9D1�o��.��������K]c����T�5 �?S��DSu�e�6�i����ߏ�םp����^��jy���iF�p@H:�����y��q�"����M_��iCs�븑���t����s�M����`	�T��V�m��q�n�0:<����y�r:���79ɵ�y�:�մ�RQu���=ޡ#�x���X�����N[�-<��e�v�t�H�vq�0������Jf0sK�����
]zޠ5��-Jŵ��C�6�c�V����m���mLu�7�12��82�F�����=oo>xu�zt���[\c��ӳӨ�����󭶷���՚QA���Nj��q�O�m��c�X�k �]�.3���0��)��k���oF�ɝ%8]��cX�7n��݉>J���Ԫ�������N��#��te]�N��3�c�7�V	�h�JZ	��>ɍ
�b��`�!U�\��"(_�P���@�/3%m[^��Q�݅ʡZrdp���CkU�s"��b�n��&=]�y�6Z�˹Y�B����ݻ��1$�^�v'l�{6�I���U��^&E��ǱWv�*uI�sp��2�:=�&�J<�����8���U���e��%J*�e�+; ���lz'n��f������x�K�u�[ċ�[���� L|o`Lk�PP��j��)�D*��tV��6��_v�ԃ�[|�_ܫ���i��52jY��؃��ԔXS390���Y��xe��+麙���ޭ�+��Z��.v����O��y���*��R=�ާ��G���M	�k��H[�������5qƠ���i�J����c*�-dSs����yw���Z7Zr4d��R��\�݅�|u�8/�u�A^>p�ڃz��o��8���#M1�b��t�ݔ��Z��k"T�/u󗲷�j�ڡyC�w�j�ub�U�i%��E��+��7�u�n�;T������ʇΩt�w8fs6{^R��r���gys�2�eN[opWrz����>��Ұ6V�B����Ӱ�R`^��-����|2Zɷ�3'h�b���^e��@:�G��Rl
B�\'���/Of&����YǨ �rlXx�뭖kz�<�����_]�P̹�&����2W-F�����BVBΰl�{�2�X#齰�5U6t��FY�xcoK��Xs;�Y-��<6̓���<:�}s������8��Ե����4�0���4�O1�u�W�L\���r+3 �*��������LP��.`��Z��<�0��Vn����*���NǼ���CAڛ2�fIl�/Il-���gN�������[�P�ά�+j�Jns}0ŹE���+@ٝ�Uh4pp�S5V>UݐS(c�h:cj��&��y��Z�ђQ�[�Д�ۜ�n�i=�j,���\T=�SMn6#�r�jA�f��R��N��x*�Ыo�i�qP����;d��x�+��{��&ﰤ�[+�]�}�֞8�W^#'�G\z�@.��ICW! bSs���=:_4_�;��`:��xRXT^���
/k#�x�s7�RBZ�妪j���ϖ�
()8㹔yF��#K�S��Z9!�U�f�g
�yi�,�5��m��!�\����Qy����r�H;��y����p.]�J��*%B�2�N�%�1@e\#��Rt!"�"9��n:vdr��3�� 9�p$$�s�$�+��j�$��
���TQd�9x���Er�r���S*�)6AUW���4eP\(�'4J� �T\�#%�AW
.D�,"�E.s�r��I$��W)&��"��6'8���B���$�B9�Sdfr��Jʈ��&C(+s��S�D�BYE�MH�ʸP�q�y�9��x��I�o����s�1e�����6�c���s��y|�xdŔ���3�y�����-7w����E�!7z�91Q�X�����.-�B�'��#ߐs���<G���yc��'�8��l�w��Q��ۉ���u����n��;��O�ױ���i�������ΗN��"/�O���`���""x2������ٝ]������x�v�qSz}�2��	���������[�|}O���'g,<���.��G����8��ۜ�N�ל>��=M�q7���O�8�P��>JpG� xG�3�/��V�
�[��������$?�p~��_��v�y�=N����M�{��z����O��8��N��;{�1;�v~�H<x�p���&�=N:O�8�����p�#�f"<���*W��� l���9����H�B"�H�yO�>b��y�[�
����΃��Bpvy�μ��N=�q����z���I�����7i�BC�������M�u��0�q��t�����@�!��:���?�
~i�z���o��o�����z,�������o���M���ͧx���~��v�]㏻���|q�����޺�ES�qݞ�sn��];��|����N��ͮ?���P7�ٓ�z���9r̿��?~}��y�}C���=q�w��;8G�����'_�����N*w��c��!>�|���9�1;�k�w�޿��0������to������� G��/���*�^�w��Ž�|w�k���~�����7�q������O�}�s��aWz�g���L>G�q�e�>�q˜��v�o�>c��o��Bt�w����Sz�����
�AH��q�z�}wJ2��=��Ϗ.����۴��}N}��8�\���O��&�F�~��z��>������C��{܏]��w{���I���vs�^F�'�}�Qh
��>�>�)<|7�^]~[�8�+c<�n�|�}" ��}IT}`3��M��޹���z��:�y�[�n�?$'���1�����q���!��n��v��8��q�o�_�ëN�7��vr:w��W��>b�
c�c©���z��{�_�1�g�Z]� }�C�D�D��^;.���p����}�~�۞��刺���U=v��y�$��������o��q>;t��]��8o�t��;'whG�����?��{��v��s��2��
��*��B�ޫ�jX�ݩ�k��0��z�-Al��f�^>f��s��� �]�p�5��ըNް�> �-LJ��t`/�j8wMWeݻ�Հ�'�Wr��u+X���@V
g1Tٵ�����hтWK{�:[�E�O�̾�z��):{��N�ǧq�V�>�I��{��Ѻx�ݞ}���L)�������k���qt���z��8�탎�=q���{�|L(}w������8�����$ȑ}�}\�gv��v�Yy�}��}7������벙w��w�v��q����m��n���:q��������1'��&����������b#Dd�pd�8C�*�������k�{��;�&���o�Hu�n}��8�}C�r� z���E����M�$��z���o����C��������ߝ���z���}|���~?|��#�~��|)�b�Ǯ���5Uu����4�&��ȿF'q7Ǐ��x�|L.��(>'N8��w@�(��?;�]&-�I����ݿ]��C�#q߽�瑿�+t�]����{ٿ��
1*�"p�٭�V�ݏ_�H��ڮ��8��\���~v���\}=��i�B;q9�߽�7���{c�������um�����8�ڣx�ʧ��aC�G�A۾�\���O�$G�}���ڏ	����ӏ�菠�C�z{�����0���}�ݾ8�;{�s�	2���s��]�;w���y�=v�����{c���7��t�;q瑉�?Gn� x���9p�v�u��vQ7Lb�g�o{��"$}>�>��W~O�&���9�;�<w�_tq0���<����]�py��ߐ�z��n{�:��8�}O�9�v����;��'��n&��v������.�Ӕ��}�G%j���
(Dz+'n�v�;�_xt;~t��9��[}w����t��}x�矽�;�bw�����;wI����<q�v�hqǾ�� (��=~s�����O�~�t�P3�s�U-y�'�}"�}"��H�O��r۟�{_�t�]��s���a�u�G�n���Ӿu��x����^;�o�s
o������G��'���ޗi����y}������Y5�Wrǈη�x���>c�1�	������{c��;wN� ���z�q�������'�qu��P�aN�Q�n���q����c� �/��������Rw�k��w����ޡ;Ü�Ξ��&���%w�|�,"��5zmM��1�l)^s,yKo���P;�{jos\ͩG�\)v������A��
�z��aZ�K��cG�r]�^�c����O���2��ɏu7��/y9��WY[�Bz�"��ˡ��l�e�zr]p��"p�k��	�.wwO�v��8ޞ{�A�N�<��p]۴�������Nv�!���>'n:q+��$ߓ��>8�+�#�!㸒}C�t�]���;�z��þ�� }"��DP�7���)�;��`Wb���7L|�D�[r��X�� ���5X���ۉ��<�hz�_m�No|���0�~O\|N���M�����t�;�&������	7���G�Ei������^��'}*.}{����}~���?;�����N�ǩ�}C�}��(�����!�0�m�םu�w���}v�s�0�����=�x��©�>��;��� (��q]����P�}�G�wQ!לH�������k�䛤'���t�7�﫧�nӟщ��۪���t�����z�Q�~_{�.��T��&��w��#�;��v��O���7��aw�}O��y�'��D���N���	�ϞC����7�y;����ճ��|OS��:@�'|q�G:��n&�	�w;u�8w��������#k��v� ~~k�λp�];O���<N�x�W|�鏨G�G�H�C���Ϧ\�˼�+�\��>�����4�� q#
{��!���ӽC�>|��q!&��r�a�7�s��:;v��N�w8�??����.��C���m�Ϟt|M� ��;�_}�>���}s��QY9i����/s�>� ����>#�>��LE��B���|��|W��}x�:�������N8���:w�N8�㾜�L*좜���8�|��N���#�}�Bܨ�@W��Iz��C�������/�%,��}b"D} ��W�_�}��y��G��W}q����I'��^?�x~v�7������\
oD'�n'<�x�ӵ[?�����A�G�N]봩���׷��ι������V*��u��p��y^\}}����w����]�|��ޱ����8���+�M?�}C���z1� �/����޶���N�wÿx����M�|�:wN�)���(I;}y���sϿy¾�}:͉;u�n6�%��|G�z��=�\.�w\M�<N8��W���M�~N!����щ�P��~��!��	[�]Ӽw�q<��Ҹ�Bqߞ��;L<��>oc���ۈ%��ܩ^�H +�O۷I� �\�++l�X��#|�\«�h���aId���9ʴڼXU�w�o�*L<�]n+�M�K
��Ĵw�Py�ލ�%0L�U�-���W_f+�5�r@b���ֳ�����V �%�(����Ķ�q��P��Vm��_͎��������v�Hq4�X���n! q/o�'N���v�'C�����߹�t��/-�o:�֕�����y����B�1%��o�qާz�0���8��߹�~�������>��} ��@���|C��ջ�A�t��I��Aw����c�G_�!����8}v���w>sn����Wtp;@�$�����:��;I�B~��[v�W�����(ݚ����=�S�����4}�v���Ӽv�o���|�]�ڣ����w�C�7������[�F'x�\s����N��:����>��}��w����i������$����s�
&#JC�]�ۓ�;��uU�B����zۿ��ۉ�_��t�{H{q7�I;<���9��v�!�Pz�x�p�C���M�q8��+�M�>���&��bw��w��>��8����W�ʸ�=7*m���j#��>���1��9���F:WP��ϼ��0������`�"v9������|#o�۱|}�9f�nX칕��Qw�y�Ϋ�N"r����w�x�\Fu��ʘxb�'���k"�(w�(�#Y�I��ȸ�w�$&8G�d�w�NQ������@u�Yd�WF:�g���n�؀34$�����0��f ̣0Ĉ|P�q;1�`xK5�-���w��H�9��	��{{fo�>H{ܶY���d�pg��مE��:��U!�'wdr����a�]c*H}����t�t�7��muϝv�C'�a'�wŕ��!�}7a9�d��ȸ�LwG�	��9��Q�PjR�|��9Cn��u%#��6�J��.=������$6T��u�6�hV#w�[�{#�a܁B�M���o!M*��y7:�q/��6���AZ(�yfM��N���!��w|�<�="dA��ya��
�x���]�WBйm���U�*zr h�\c�L���S���(Ld#����&�l0t��F{f��am�u3�8Z����	�\��Ƥ����D1�o����e����vλ@U�[�D��l���TP �!���Z��9M�ƾr�	k���ԝ*�8��@W��S!q9��N��U�&�dI8_Р����-$_���̎2�TbuÃ����l!���@ �fq�|g���z��KO�q��3��;>�:�d�:2���J�u�.S^r
Z�1p�k�x���}=H�b,"u7Z�;w
c���� �9����E&֪�ֺݙ����9E�X3�|&1��C&�7\�,���UR�Q1 &F���6!�vl�Z�<���L��v���BOo����M�7@s�j�_�1���zv�G��VK;�Q�O�B�c**{�/i��:��ח���\�ɯ�K�;m�ٚ]Ag�;CX��) Zs5��ɞSv0��cu��`ӛ(;�ѰŵO�1s��pz��M�F:��b��Ud�2Q�IҒ��]�d��:�Oe"B#$�c�٨��P���T��������Oo��8�؉�z9����|M[I��skkC7��h��ǋ�J�ߞI�AH�ȴ4l�;Ky�����}֏�CO�i�]��7��eY��w I�3��	
�[������m��c��&��;4�'�*��i֣�hn�յ�FUԋ�bл�mڼA/L%��S�Y�s�U\���f8 �_u�S�l���}7��tjyl�Jc�[��KG3�яjM�mf^�}͖��a�ۄg
���s� ��h�/]��ss�7m��*#:rN�E���.�X�J>�yJ-�M�/��!8<��Sj���Z��t���0xn��t��V�!� v
�j�͏�^�:V`x
��עVH֛����>�|!���#h*8�Fㅦ��_��H��ڸ|l߯��"����C��]�l���Ϻ�!��Ai��b[9�g��������B�&Z|s�G�����8�?��	��1��OK�������y�[u��vgrޥ�ӸB��>;��M��#k�T��)�������ĥZ
������������\o�j+���-�_T$�"����k��w�\9�JR����'D\�S��n���ڪ?%gэۋF�]׼�X�6*O�%�җ���}�Po4���z:�p+�����RZ��,�����ĝ��О���3��S��\����-m�����Aa�o���:c���"���|�2�=Ѷ��8�֪��B�W�;�R��`wB�����6��rS1��\�%�6��H2��s���S��/ս#Tx���]҇;������pԭ��go���Z4�'f��s��4���)��5l�T=YB�C!�z���M/Lʶ:ɦk�Ciu��\rwr]T��]z��,�w�`r^�-h�r�����^'X�]����{�D���婻^ٮ!]����8L����fY��%1B�t�]o�@Y���ok�g�I�J�v�MӌQ��)F��7�j� �d�BT�4s殢y�h�W0E�`ٌ%Y@�Q)Ɯy�]�FVbJ���ɞ.*g�(�1����S\�'b�c=p����9�q�h�YR�<m�*\�>���;'�8�c(L�Ĺ8$�g��_�j�jy�S���/0�S;׎9ʥs��w���8X(��w�\:P�X���AXP��_?�u�9�[��Q��j(;����Ol�8㮸5�b���F��~�TV��[�|>�� �Ι���ڞ��A�؍��`J�ׯ���:��*�^Ò�n�$�[���j�`�{�W�P)S�9�c�=kڶ.��l�E	S�V^�r����4��ذ�i�v������	ݬ�r,]o��{�
��&��g"��MKm6N��BkY�]�>�膛["y�Wh��=�&ˈ�@=�N�zo�W\��#Ĕ�PYc�Kp��'��;���'BwCy+8:<��T�;If6� ��c�#o�����Y<� 3S�x ��Sf�;a9t�s\LH�/����Rj�l�=��L���#��q�ћ�2��Rv���5��{{V�8�@�s�����]<7�;l��)�3)7Pv�Ahi.ܖ��n�7E����=Z����+k	�LO�*����Ӗ����a ڢ�ڋ�r�f�[ˎD�z��.��Q��\�����(hfE�"nW������-�`�Ce��.9�J�#��ٓ��X�(��'����(��BӅ�ED��ӑ[0��DƧ����D�V!�/�&������9`ih��LGK'j���49�P�(F�G��~6�p�=��{Gn�ZN�N� 91rP�p�݋�/fr�1&$�Pg��Y3K��:�*��@��j&錿���<r7�3�N���I�k+a���{Q�CLX0�F���6�;n��n�����w.�3]( t&]Bx�����8�b���:�0`�ݼ2[�u��$�2Vhπ�5�y)���]�fX�Aj�r��=���������c&t�k���@�Z��o�4�˯���@�d3ˏo򪾪ۧ��"��(pi1�1æN'$��'�'.#��z�C.�������N.�[kJ�9c��z�_�yS���U��i�n'fS\��k�_m��Gp8^��ʅ��Nr�V:���ꦏ*^�/���yp��87\�;��ls�!������F���V_�j1=��"��'$S����1
�W;"V_���hd�,$�#�.���,�!&�!�y��ķnWY���p
4����Ξ�!����3�LnB���ba�|����s��T��N;ԯP^�;��c���jF���o�CRY|ph�6�T �R�#���b�.Ϊ9�\�b� �j$�B�J~ߺ�9M�ƾr���H�5'Ja݌2s7V���}2���=�4x�� f���S�0��>�ߣ������C����M�b�{�э�x����%�|�d ��0c�ShϢ���X�ie��@�_�j�횩��W|�&�: �]ʸ?��D�a��÷q4`���ҼZym�@T��؟�]nŞ��L��E��;�~ў���N܉��6P�=���K5��"ɵڲ�eU��~���w��kp��Rmp���_rp��.�͢��-��"ŭ���2".\H�� Y[Y��pWpXD��ƻR���ىU���/.Oz>��׎偱��z����B�*6�T2k��p/� ЄP�@�M���	�o'q�`1V����q���Ϝ�B���v��K����MQ
d�MH������0���e��\���Z���z��$�q���PRz���S��c~���;��J����=W�i��p����I3s�h�/��8X�;~�s���\�I�͔��6���F�ˇrf43�9��*�MR�?�u|�*͞+q� ��g�Ϭ$+�V�y��Q�r���x9�E,YuZ�-u���vl��1�M���ɩ�W�O�l�C+�����.���>�pV�l��a��a* �]d\O:���?c��v;�S�e�1���%�U��`�Z9�	77�+2��}�j��b=��p�,2i��_l<��V�n�5p�}�+�2V��4�/ϝ.�qQ��@��P&t+����T$��?.��]���2�ۿ������w@L��qh��a��<(�o�p��Z�ckϼ���T�t�qw���TvÏ|xZ�w:�ӣo��[b���3n3+#g�{h��W5��x��+k��~�#/���ն�T��r��ft��j��׶���ǉt�z.>�	������1]�c�iB:Ԓ����V �N�HKCi�%����x�����,z��k��w��GH/"�����cE�Ռ�"�W��NH���껼���ץT^�H�{�����(z� �5�'�k��G3M!F��8o
Q�����3\Ue�G^���}�E�d�u��*l2����-D���l��r��%����Z�n�����u����@�9[j�`w��:�rN���L�t��A�5�bM�9��k�,ow{7ȹ��	S�=+H����\�<��cA�#UX�yo#�0d�נc;�骘ǍaMf��wQXt�'U�N�v��S��:�=��\ݑ����vE>� ��Vb��U��6Œ�eL��(j
/8�-v�ƪ��wqwP=*�CW6q0}kR�粷�L�a曰3C��܋G΁�lC�:ƻ���u��4Mo*+��h�ݞ̆XuG�_Q��gZ����gSۖ��p&��%8�9�*��"V7 ��}6ܴ��v�ܧݫ�:�m��̺�#�%�!��49l�V�y��ʽ�23]��]*3|�GѓP�z��a8��' 2,aν��G��R��Ȟv}rx��d��X��t�k�*��HW�]L}��'�+�rn�w�S "�;Y՞4����Z� �o����|`Yծ�z��G�f�®du��۱[�yhԹPC]�:Ev�#�8��
��ir�N1ۂ�@�_ro���`��=���x*]�ܳ��;�7�&�q����U�mw`Jt<%$�fnՅv�(��GGV�K��gv��;��%k鸰W|9`|Nd%�gjg���L�g5$V����`B��dd:@�M�we�t�ݍ�mAg�y��BL.�J����,�z�>�!�`V^���	�%���H�s�tAm�h�u�}����u"�pB�ǅL�טgS�Z����z��tq�������K3c=�pђ����ٻOXO"ԡ���ƨ/^d�0wl�a���^�
�nJP,�*X}�qqe��p�����bv]�CO4�N��-��q��<�԰��8�f���M�ci����D��Wz�D��S����]� ��/�,5�^���U�C76�����qEI妧�^n8���(an����q�����Ia�n��#$i��4c���Y���+4�N_�O�ȓ�b�uU�k����|�ʑ^�������묾�Xа�q���vNp��*J2���LlF������=��Wb�� ^>��t��u���8���l�,�RLu�oDC�n��7�[��pЮ�<Ji{��)�=�j���6�5���3AIsR>�ڒ����9�>X�>��zh���S9�^�xmRu���4���'��I�A$�~�O�/��Up�D�)$�F�F���,$!*��r�U]JZIEI2�8�	[6�J��:r̋�r��f�g(�+DV����tʇ9s�		jPY"��C8
��0*����(�$� 9
��Y\�6���J�!�E9�JI��G�BI˧H$W9qp�(�;�q2�Цm��qA3�!h��q2
4����]-v\�2�򇉬õ$��Jk�&D���.P�ft�W.S4H�6q!3$�TU�"���M	�v��REQr���r�����L��BI�jhX&�����2
�p��D�M+�&Ds2�:�f���8�2��)K��A#q9����j�EY�b�.币Ū�i4��FȠ�P�
�K(K#�K�x�T &�0��#�f˰��+���ǀ]l4���DFDj��|ˮ�0�x~�%�|����Ě���a�w�#���޼�I���n?��p�)�~�b�GI<
q 3J�K˺hBx���}�x�l�[�1gYc��M۸x.K5��7�0R�&��V��s�����b�c�)����X�%���p��NS��!��ق5כ��$y= 4���Vˁ\u��݃s�5�'�#ٟI���xW�9H�3�9v��M�nlA�S$����s���w�K_3�ɀG�W�%�����L��6�K�ɸNc�16�x�`9�cr���N6�p��`�pfc��X0Č�,v���Zms��|jLTrN������gMs\F�a-���42<��p�t��!��+��2�Wv����X-���"\�.IX��@t�',	5�p}Q�*A�y�&�k+����۞ā�s���?6z��|���d��h�Ӫb19�j���=�L?�ƅX�e�x��]<�)u���9�W�r��٨��]L����3y���<%)b*!�������計�W�l���58�p��4�ɠt�{D�3���@�hW0��U-U�0��&�J���U��q@�/&�F�)�T퍅Q���'(�.��{�:%��u�5m�tWN�[պ9.݊n[����0J�9�_Ȑ_{
%�.��C�#���Oۈ��)u�����ڏ��$��T��|kV�s;��b;�}*k�dċgzW�\s����s����isy�D�������%�3�%I��*��P	�b<�S��.w~��vja<�94�wbQݢ�ƿWt�5>�`���n�����4�)�*���A����$IY�v��i'��H�C�)l�;�a��0��Q� FlA�2JOq�E�C/�#�]�o3�&�r����o;ё�&ˌt��9�Y,�cZCKm0�{�m��酗Z��v��o�J�����%��O5%��r�я���n��`�*��7��b�����V���
�6c�Tl�vU��"�Wpe��p�a�ӐܑN������+���F��g�C�Az�@�W ���F.���f���G�`�_w]�ʾ����2Ҳ���G�戮D*G}��T�a���,+S��]l!��z�V���2n�'�mA�NO�[��Z�`l�u�42-����#_�����3�2(���I���]R�Q����y3�g%pLYS�70]
0lɑL�	�[ߺ�kR��8W�RЩ;h�7@^J�q\ڦ��Wپ�4��Vz���(Ƶ�'SJo�����B)M��K��
�7�����n�='��w�y�G�G�D4��5Q�m^*!�ʣ�Bj�/���"�����(���d&��ڬ�����ny:f(���J:�Ϯ���-��Ԕ1��健����<�3�l�7�����a^�DVR��U��#�؉ͭ��6�Iۣb3� ��	FW�U
�Z�;��0�pڮR�58�����1����/>�����)��n����xb�qZ��j�%9k��7[�YZ㏹=n�Sl���V�h�-X�ճ�<L���:����\1�e�*F�{hS���w��wy�����L�S��N4��+�x?���%Ho�a�sj^à�U���Q�R�<9���:��u?fo+�����d�ݖ��[��9��W]<�:�.f��Ĳ+,��ꠄ_��)��s�n��p�1�]}���m�Βt�����{��P�o�{5��W��-��F��Э�ѨZ��dt���ˈ�p���J�3�z;�Mz7J�
�םչ��{mP�I�p�wS(�F
;#Bir��u^�|pU��2vJ��i�ή�s=!��^��!^�w}V��MYX*f�Mol�.�m-��K�{�<T8aƯ�d��ؖQ��x ��kM��ħϫ���O�]����k����ѻRέ-(��-�An��yf�x,e�`t�9��)ú�U �q�}}�WM�s����+���<\ 8a,	<ҟ�:�9�7_r��Z�"3��Svj��$<��X沛���2���.�V*J= �2�����&zbPg]oԻ�.YK'��Q�v*�a?Z��Ge��ӈ�����'�:z�����(w:���T��YB�z;T���c.��ޜ]���� hi�A�<L8�c%78÷q4`�_�Di"%�>꒝�펴ct����8=?t��\��o*�M&�x0��b��U�6a�ϔ�_Eux�9�??Aj#���$$r���+�O+�MTP�S&�n@֙�\476 ��nVt<�I��T<�\)�skl��W�<%�pv�.rw|c"5�̔#%��^>��V�\���T	N^ٿ�zg��\�����Er�&/��A��A����涫D��ᤨv+��a>��tc� ��w�}��7f�U5^���`�)&ܰ\�V�j� '�Y� u��r�NNlvrn�=ٞ���5D�y���w4Uu�}�����#�Ʋ�[5�8�]Z�`�;�f��X�� ���Hk���7��<�Y���fݙ��|7a��g��e͙4<��V�qJw�����XM��N�{���1F��R�5&%��Z�2�v_vp�x���u8���q,�)�j�I���������;ޝv:��g�+ L0�.�.'�Cd������p����Ν��Oй��4n��[�=�W�p(�.��S��u�Ѹ;.��'~jy��/����\ ��v��A�%��wZ8ޥ�#c�<�4���%��KڪV�aWc���5���=	�e	雴:3��N�V���aߨh�.�����A�
�ף^|��ʘ=�~n�c�V���&���U�Z�H�9��Gi�p� ��~�!	GI<
q 3J뺉s���\�Y�/U5䥛�bCU,`���1��;ŎCv�Q,����&�u�v,,��,N�Ū�ܞY]��8�8f�B����t�8Z���[�J{0F?����'���cig�����nZQ��:�@��٢~i:H�9���;X��؃�k��BŹE��mHK�����3�����3�2���mB]nJf8C��Kآ�/:OEMR���яNPf���	��V�1#>��i���Zms���pP{�fe1�-~T��H`���QԞ�ZuF�F���nt&ԡ��M���]j�R���N�Kx�V[�P\� ��;��J��jS��-|;^�{��+��w+�ߞ��]ϔzM��*�/+�⭝%YY���j0��gǻ�/D6̾Äu����]�>��%_^���6l���Lד�4�z�P�*m���[�t�Vqv���u��'r̻ro aE�:�D_*�ߴ?���0�����g*G���pe��6䳫�����|fZ��\������R�ʺ����тh����:͹�vn��Z�B��&�A�/����]�w�쭗S7y�t�q�ْcX�-��m�c	�J���U1;��ۜ-����:��N(�C-n�]$3A��U���VUi����G�D�cW�<�%��Zj���ܙ�w]�����#5?zeޮ�?Mc�T�Z���K������������0�kS̰ON<����ͣ��*}yz_�U�lލ6S�C;s�dxZ�qX��S,EFҠ��4Tve�Ď��A��%u��z9��_ �h��	�ί����1|b�eJ4 ܃�d�$��yV��'
JK�B5�]Rs��w��n�G`��FDk��2� ��;�鸕��h�u\t�Ί���@�e�H��Zo���7}���4���;Ѻ\u����J����m���zq����w;�Nw)J�>M�')R�����x������.�twW���_�LI�-i��JNɝ�-jY=-���\��*����&-uR��ѽL��)�4�<�[7�bcJ1ۤmf���c{%�kAspӗ�< 4�Q�S�T���-+����j�Н�@��c�"�$��Y՘"��%?���>���;�H�ծ�2}t	
a��$z���.9���Y�=�;N7$GT<w#��Rs�L�h�]�U[sfp�D?���D����)�|aq��up�T�l�`�>QU��A����g*΄!��A���3!QRH��1���#�^+J��\�}�4e[��J�;kt��O.�Kw�x�����>t�G0%[�٦�#�4����Cy��ú-��hKU���Q��*d��偮@�!:�#�'`����dU�j^W�_i�Lw��H{}0���m�_.ylgɪ�7��@b�����{�x~,����ǚ��`a]��N�p��ƃ���=���{E�V��Ӛ� ��Ib1��	L�;�C����K��3ۇ�2��V+��Z6��إ1�Ҹ�=�)���w�F�I��=�t��]�E�U����f5j��M��F#L�Xx��k���c�V�Α��nn>�_�W�p��%�yrwm���z����nE��|(��?p���W_އ�����0< ;B���K3���S�Kr�����r�eg:�QP����!���e�ɇ'�Tν��K\4�N�k�H���բEB7�AcM��o��
��dX�$��Xv����[�/[�5S��Ҹ+l���|9��q�c��q�ʷC]Y�����%�������B���]s9���"�%4�Ꭹ2��}�m���Sƃ%.�?XEs�ެ*IX��~x�\z0�������X:�1�)��s���3�r��ދrކ cG�ڭ����ޑ%���t�O�$��:gV��Q�^D0�Bf�Ln*��k��W��n蝽:���a�<	.���$>�W�L�_�s���4�[�Ie��
�&b��o��$1m�f,8=7�`85�	�Pǁ�ZS�T�f[���r�~h�݊b!�+#Uto�7����,�f+�Ty�Ck��+�ý�	ߙ�l }7��P�O�q8��L^�z-%��b�T��q�7!��&��<n���0���	T@�&9�4��rL�F���C�����ᚎv��ɫC>r��`D�n�N�v �f:��3����7��Ϸ�����e3�8�V���.B�yL2{��p/� �hŀ�P0��PS=��z�6��_��Gv�U���wJ�p����5PE,��f}��}�����ew
�Ħ��X�g�//�L	X(��^.z���ED`�ij���v�Z����K�++����,��Py��mwi�ưy.��N����l�}��OWl�J��7��ҝ�IZ�W1��.
Y�07y��*jJ�B˰�t@�"i#ۄ�&�ߨ�b�����}DG�زSA��mj�La%�g� �N��mm�����.������I��Ü���N����9����/rz����>¬��@j�E]���
��-�=&3J���y�`�&�d�5��=��F��]���0��|v��x,Z���zQ��{+�	
���y��Gm>�)�
��J5C��H�6�{h_^��.�8����U~����?��Г�^'0�m+�s�)���kb֥'�
�Ջ*^�3 � ob�"�y�6N|��}6��q򥚥1���#*{s��W]!�)���̼4gj:��T��LCF�ˀ�0�h�+[���p�n��B�{yrT�[=�O��Pz����*b$�=X:4����BLR�_+���7`2���n�p����k�g���>?3���p�C�0A�+�T�p'V�����|i��TS�|�;R�+�+�j���
��s�oa������K!����f�0��$2�W����mu����)�1"�U,`���h�F�x1��n�Bb�_�z`�(	>g�f�f6�9��+����G��{gOY^�
�sǻaE�Xr�R/|�;�sru�v�J��omuD���2���I�J���h�d�]�7{�nϦ2�G�a\�s�`!�R8�e^��H^��Zp����9��
����:x��Vuh7��{x}�337�x��S�=�A�^�T���+寮*�;�ܾ9��!��ق5̡(��ْ�ν+���� �b����/K̉"��+䜤W�gD6q��&��௯o��tV��J2�D$�!T�� ��_D��h)���6�.�&Ә�&{h -���p
�I�_"uƚ�)M�EB�����s�����$U�;L\wJ�p��������=;�JW��T8�kuY�{ɚ�]455��a����s�h[�.'=7��$���o��h��j�XO����܋����&�����9��'�d���N����\�9R�����������ٽhh�5e�J����3=��1�W����4*�;뾻�˽�{��µ�3��z��P��}��e+�/�S9���xM|�1�bw����Xǜ�Ρ��3�/3�N6p1PNك?LTE�ЖpiE�d�]��L�Fq��3�L5(�D���,�o\r�g~~�w�8j��#f�\.��eR^f�k���8��xR��ǛmJ�#p���x��t��<ʲxu�6�ho�GPЗg���K/5�{�����rՙ�-
�y�іN�J�R�ɗ���������w�a}Q�*JA�}��)�T�h��Ⱥ]
t�m2Q�|�M���/�0��2�n>v!���X�m=Pv��Ƕ�f�;zOǺ�jސ��0*�&km3�2R��/zWs��ғ�ݝ�c��+U'j���~ӏu���]J��L��q�rWmka�9�*γ����g��+bb=ϯ	hd<n/�r�l�95���YP����C��Į�3o��i�C�C5�_.ay(`�!�l���|���'[��%�m��8`�-"�V�j���K�N:qD�K�JtOI��ڋ���(.�e��ӷ�������fV�w[(뎗V���d���I��W� \f�8�,]B���5�[�;�#������F�9������3ԅuf��vb�]"���:������h�X��;�.�Sp�Ī�==J�W���o���EwF&ͬ��&D�#Mi�|l��P{}9(#���`���;MY.�jr��A���"���5:c�8q��q9x&�:@\��!j&�.�8B�,�Y@׷��E�Ѕ���s`�6���
��;�:�B3/>�_-#8i���̤�k^ضC��d�h��(��U�7.�����&5;y�#M6���ZqE��g���|6)P�5��v�9�p��!��1.�GӪ�t�:���l�K�K��dd��wm�%�ԩ�ƎP�l �X�Gc �Ԧ#�S��|\=��_��6��
;n�p���TV�i��7z/g^q��J��k�%ƞ��$�Z:���P�C_0{�k;��dq�����{ۆ-���[�uػ�\��3���K� �d��y*l6nes]^+��XM���K-8�O*f����$8�����yk9�!jL}C���t�/&7Wu�M�Μ�]�Jб7)6�E��8���j���7h��PS�r���D5�g�q:3���E�"��4x�Ԭ��=�nL2B!�*��T�7�Cn*�3���d4�y�����^�1�,ۇ���Yd>o�����Cэ����N�����3�/v\���m�YKQ�Ts�WL��a���l�5n�]����OVt�Q.6� �k%k%B�,��=Ņ�b�����"��۳��[C�:N�Z�c]Z�6Y�]�wb��\��]D�XA�u��;׻�jNɇo6�ͣx�M�N�!K�vԇa[���+Ae4�]����vo<��noZ���7Kt��t�2�����8�3+P��;�
�y`�$���H~n<��0���J�%���=��H��O�r �Vv5k�g�ޥ�N�>�H��MRk��	��53��Y����I�v�����ܝE��]�wi��z�����&N|��AvY��������}u���"�Ҥ�UNE��q8�m�H�Sf��q2Ԃ�	'2��LUK��"ANZU�����W��l�9aċ���4N�%$����
D�<I9Rb3(8�E$P�2���1��PdjI8�A�*�Њ�G-JBN��ӥns�Wn:Ȼ)��$RE*&re�����q;$7+,H�U3����DuZ�,�2�&��(
�)�n!<J��&��B�"c(q�q��r��������D�
ɬ�2;�hs�Qs���Z"�L��fy���\�r�V�hdDTr�f���AVt�8�^:E��$�͐ND�fȪEf1&����	9W1 ���U�#��\�Z�����Q&uF*4��Q���J�1e�T2Q�Qn	��wG�E䫥��h�;0�˾��4j�m-v�$�)T��rߚ}SSj�'��ݝWM�����/Hk�Y���菾.�띥���v̓���h��5�3m;�cE��~�w�@:xg�/
��q��{���Q������1hI�� �9b<��u��*���qb����x�+_�V�b'���6��X_�*��:��kw�5��q�����ܫ�IF��J�bȜs����OV�r���ê3��6T�.'���5t�ڎ듿Q����U�˵����V�K�iޮ�'x�;d��0�TH�}�VMTJ2�q�3v�nH��V��]��g)n;��"��}�+h;i�ܾ��Z!q���z]$`������7+�mP͞�u+p�bMNѝ���\'�ԍ#a
4�I��B��Sg�O�*��r9k�Fm�ht��8}.�[gŵe��4�l�mZ�NQr�6s#S"ߑ��-��iC}��wq�>���Y[=G�JY-,yDX�A<Qle�/eٱ��O��-3%-s�FM�-3���ۆ"�\��MMI_d)9`ix�����sxJ
���-��9��:��٪i:�} �h�{Kp�rV�uܝ��7�6m��=^E
�����W<0ұ	��d��耓@�� \�4wۑw��XM�%�Ei �u7��T����wMn��6���=@l�Y��f!��h�V+��jV�w���>��-Vj�t�����C�)V��/��c�ٱ	'U��S�����~3�ݛox����^�#��Ϗ�����ltJ�ƣ�B�kl,ּ[�T>?�^C�B243��Yqy�c+{ͺ{�}]�R鎯�5�����tk��͎����Ԏ�s��|������9�Ћ]c;cC��p�c��{���|j�JΊN�*�}�<.�N���OL���1V�5h��+8`L,V��<�c�L��u��n�nL��,��������步�y��-6#E������T����g��߭���pc�3��z-�u�+�z��%�j�� !�-2��ƴÀQ�Z��dt���<���&b��J��E����@�q�O^#�Ƞ�|&�`$��*��U4���0Q���+�=<Ԗ_z��n3W��Um^�B��p�F�} �(҂ ����?\u�&r������Y��s�0���9M����ή�ڒ͖+�T2�mv�A�3��`��y�� �T>�qE����J��.�k2�\�V��[���CPΡ���R�����iAm��df�^�jW.��:���i^��j�d����a�#��	��������G��o�Z�ZWgA-6iC�b*�+����K����m�C�����q�hM��_W��UWxv�oK}}ah�Y(h�*j��g4���w��N�,����:L�welFwU��͍O�̢����5\.�G&�T�0ٌ���h�D���h���\����S����| ����O{A���q�1P�
��U���-DLvk��Wx���E��̅A�hΧ�-��)��>�b���x�x�3�!'���j���d�Mr�-��N��g$��`,�2-��$�L#�PrP��1aɈ|-��W�G�js��U���3Y4��M+z�r?q-���w�o�/J�*���E]����z͇_=��Q�槎b�=�l��ظ��z��o�9{qй��	��s��x,Z���q���3�g��x�ҩ2d����9&&ȍF�������)s��r��){�n@�~{��̽3<|ըeZ�~&/�V�w35���E)���� K�z0v.�.y�6NC�����Dk��w*1l�o V%F���vmɇG	C	Vp��+�UH�WLCF��
�a�P����������i�vC���t�F���;�HsƯ�po�<��&�n�$xFCj�h
�g9M����k[W]�q��)���	&dS���gӕ�m�[Z�	:1��o���!R��՝e��,�Hr�P���fV0�9P�v��]j�f�C��������Kg�m�,V?�o�Z�pI��H��X:4���C�x+y�~�o����9�E2��R]=��h�i�[+>v���G�.�"�P�������w9�q���gHZ�Ѡ�������P�.�e�(ؾ=>yv�ZX-wL�`]���H��^;1�������vr��pV���{��u}��ǖ���_���з�����pV�qIۧ�L(��@WĶy�5�
���mӸ�����!��ق6�R�M����`[[��g�[�nZ bG��A�V��$B⻧�I�G>s:!��v��ɚ�yY�����W�?m��<o�U�(��������g��ؼ�)���m%���[=���I��6�<}FA�ɾ'��T�$>��E*�J�5ʼ��l���/ ޝ��ΘES��Ts��ĈL��	�f�f#e��'�l��+���2�=��s���:���`>�W^�ˮ�B�9;���',	<͏��y�c^x	HWN	�C���ݏ���
��͚�l
� �w6��(�RG5R|�*�ͪ������KEZ���@��Ξ�^�ә/��/54�n�z�v�`��je��1m��]�7��owB����{�	�Ŀ1�0t��p�/:�N��g׫E=�f>�Ě��t���_}�}_}��z�TM��.~Ş@ùBf����a)�!�t��s���Хx
C]1ܢ��r��t��XV����[��WJ���
fX���s�i^�e�*�/˽e���Oe�B��-������ʭ7Ig��1i�ev�q��85���Y	�sX�o>�M�GZ�u��b*�`��3*
�:�%�TIP��b�2L���2�֞Q���j\/�|�O^'|��{��6�������L;��̗����ohl$�-X��B��_��|��|��߫@И�\��ή�s�f����q�rS�uJUµJ��\c����ڄ��S|�P]�A�lZ�n'-9�}��
�uR돺��RҊw��km�z꧴ZK/O(}�t�������3=T�����%;�����S����Gj��B��V^N6���Ru�c�ŧ�P>�9�
��w]������#�+���[8�]M�H�uҌ)�J���POo�rb�R֣ڂW;�5��/)��wŞ�Ʌ-�U~���s�A��x]ԙO��A��m^��	�l�se������su��:8�=�H0��'�* ���x�=Luj>������гWS��q��Ӌ�a61��D)�	F�ϧ�����L9
sp�>���X15�5�iD2�;��l�)G�9�:�y��&nT��QŃR�9*yd�I���I�I0�q�Ѹ��&9|�[��<,o	��?@��$k[Y�:<v��_B�k�Mƴ3���$�.�6w;Z�T��Nʷ�K��2����{V�s��#�4'�:ъ���I%����T��;`[��[o-����},N�p�YZ%چ�T"��'<���v�w�֖��e�ۇ��0+�v�ꪎ���'�Y�j���<����S���:�*�rxU�|��m�b�6&_7����]�NK��c�Ć��͌�&�v��7�Y�vX1��P_Xɥ�Jis��U���d߱���y�41�Oy�ϩ��s�*�D������ІG�+n��[���Ŋ�kHzH.�r�Q���y,�R%L|��}��		Ik��:�7[�R�$�Si�ҥǦ<o��8Cטŋѕ^պ��f�Lc�N@��,���%j�k2����Z
��c���;���(�|�-�D}G�F����F���s�!��yTI}Q���Z�\o-�o.1����`�ځ[�c\�'Z�ޡ�i��z�Pr�����ʤ�Q�'���\���Vr��đ�Jla[�t��O8vվ[e�w���A��&K�����Mb#-�B��b9k8�oQjy�������P�.R�����-5u!�V����=�����p�*��-+g5n7�*>x�Ӗg�B���b�ؚ�6�ݘ����m�5������%�3y� �$/��7�N��u
���Bw�oK�%�)B��SR�'w�B�6�s5	��wJ���gU����C���\�j��Y�`�ɹO'�b�����E�[����eg�'�o<ԧ�v�����u���ʜZ��5oj���O1�b�.Dv*=���-(E�<pv����׆�<5|'m]�/]��oq��YU����ʴ�qL��_'/�F�Iͭ���4�r�|+aw*]����+B���厰n��.��o�����wu�s=
ݽ�̪MVf^�A(9����G&��3fv��=΄�,'���˾ަu�{ǥq�'���������v��{�:`�C�W�Ob���ƻ{'*-eWQK&�hk��]v�,暉YM��b6��O`ˎ��>���OZ�j��^k���=E���f��fvoG�0n��A��*�:1F�ظQ�͌�X��]��Tz~��')�ţ���{w��9�}.z��P�k��lTC\�gk�}����5ܗo��^�5^�ڢk@���U%�m()i��	�Y��)j:k[+�e�;����'�U�D.§@УC�_I�m�*�[z�Ur�y{��~��;+�MQ��������[���m=�+�����a����J6u%5Y]Z။�ʤ�����k�\g[�z�7p(:������:���s�u�Ϯ��09�P뿸���>,��Gn7�3���{�30�\�u7ΎQ��_wO� $�PZ�������I���b]��ĝö�se�K\&7oȰ�R�8�M����4ӗ�W��PC���s���S偳�u�`f�#3pRuEOs&�9������B�;�١qHqQ8+��Qj�2�֛\�n�˧g8�tϊ�X����s�w$�_m��}}��jR�v�:�Cݻ�_:e ��%_�)��ҷ2�Juxj�I^F&���c�Ĉ�;�Øvôn%RSx=�=SM~ͣ����y���ΜL�[J�wgp�Q�䘚��kB�]��l�����v��>3�����Ϩ�8��k5�ٮ\�X��&��s��vD�1��cJ�y��z���O�'�jVe}Ե�o=��i��i�9ۆ��^[���۬ݗ#���h�|�2*��jm�J�����s�	=i�� ���#'�s�cV�I��i�5�]���Sx���(�H�޿om�<���tj�+9�q��j�~��I<d�ZB��P�V�ď��2]],�U�Sr�2��Zc6�6V�qI~ΝlL�yv҈=�\���cP�e�ƺ���ε�u��p��V6Z�إ��m=_:��U��*p�����g.�&t�i�ڍ�j�͔�kz���^<=��^Ԍ�6Q��aC!��(f�y`meN����_���`��c�G�6�;g%�c@v�gS�����ι�TgWR�,V<RҬ�u�iU;.��ܘy�Ռ�E/zJ�֌��͘��������G�,[ϼB�:�K��{
�+�\c���=�M=�S|��.�q&U
�[]oP��و;�Q%.��躔�Ҕ����=�?n{�E����bd��y�E窣��(9����%�k].��>5��1w�ψ�S�g}�l�|婾^zQϑ��ό2�P��:n)�(����Nq|�oU8R���sRc,&�#�]�.OU�'��9�(�T���o3
��Foke:��6��52�;�<A\3q*�����@����:�X�������ճ}��>A�}E$Æ�w��mh�U;!�*N���3�$d�"`�Cv��yW���ӈMQ�X��n��P�2����v�J\v���}�s>�<��߳�,���^�5��|�%��:�,�$f��];5�\�ޱ�-�@�U�M���Z6����>�qAe؞��9 �uŻ:�FU؅�c���dI��t��S�#;��Y�hڱq���5�u��ҖR���o/�����ϭ�El���-����ϛf��ի׷�N뱞xrT6�գ�u	�V�ԁ�%;Y[���n�::"R'n��|e5ʱ�@�h���$���@f�WR�`渪E����F��W�� ,г�fa�@r�Fc���n읺�����5Æ��=H�������0�x�c��1�zXWu��U
K��y0���]d�tnbc��]*�b6scwd�#�G��$;�=tY�2/aiN
�����3����;1�u��v�;E, u���+<�㶹[�����;�--�J���'�Ft��0+rs�a�fG�-65�+��z�LP�׆�嚊��tZ�tK�X�9];GKJ��.�s%dT������k���k��<f+�f�sF�}�j�-w]svk��)c�5�p�A9�"��y�Vehq�Qv1���<����;G���2p�٧7tu�z��n�mwE��_K��'�][����#.|jw�*a׹�DL�r�4I��p���)n��r�_\R���=(4V솯5D�����J����|��K->] U�;5�]�|�=L^�7s/W2�[I�&!ή,)0�m��]=�Jy{�d�ݍ:���l�2��S1�-�Jb{l��ӕ!+����+/G���vJ�r1e�h�{"�6d'js��5λaZ��*��ǁ����c��|��3y���
IڭL�,w;䑣0�o7(����.y�lӟu�D�
rzb�w���A��Y���&��W�Of�\Opg	�)���x�Y�e�U;�IvvC#tiEO���շ%[��f���mw/�I�*�(*��G�+V�1/��kR��58���+22mu�/"Uգ-w#j��W���i�V^�Oۂ2��&�ɞ�};C���E� Xc}wl�(�ٝK7��$�歮�S��^bŒ���芔��Y���2hO��O|	��{ݏ�r�9���;8�w�r��Xڝ�xr�Y�.�9'|���:�aںg�h:ƺ��RuZ�`n���	N3C�]kQՈ#�`�Aѭ͆�E00-%�avm����XE�It�eI�y�+L���7 Nmdg����9�1�#�zz�q��Vŀ+��oB���] �Az9��w��W
jj�;p'NbY�5K�(�$�8���5�iп���X�x�.��{�=O�!�'jE���V.�4����b�F�t�E�@M�;l�k	{\ѽ�;Pj����1a]�m��P�#�cݝ'P�$�Ռ����=gT0�9�-]�0��u��b�l��y�µ�b��78���O3u��}���c�ˮ��w�h�諌���ג�.��qђ�P�R�b�[z{N>�2�j��H��[��ε37A:j�9��OWr��W�Z�3�a�Mq��<��ʄ���q�ӯ��s�y�_N��w?������URt9(�9Z�%Q�QC��.Y�:Eh�+��Ig@����(�"%��Vd�-ȐU6r+��%Dո��4�#�h\���%*B����Z,��J��:T�ӚPPV��9�Y�����2�("�.� D@QȦ\�Z	%�E0�ӥR�ĥ�0#D:r�9Չ�ĴZ��W��!�R�*eȋ(�ȃSeEEr&r3�D%�J�$'%�
��AHBTYi�r�ʠ�s��#6Q�6��,�T�J����d"9UP�"H��MD �ȢU$�#�ʢ��8�d�TU���NX!��D$�Fk4�eE� T�W*��9Z���UEU��E�ed\����G.P�#�TU�9Bu��S9R�TJl�6
��i'd\��dfQQQ\�ʪ*".ʊ(�4@�Z��yi��>"��^eu	|B�_:�e�����ڴ�α�؍6M�u�����ڏx$����ք��pel�59���I���",�s?G��}5)�[��Ƭ�g��q�>���6�Y��P̨)��Us�[� e�T/��v�kb�=Q5�;+'��vs�&�M�i
u�}�s�ݞ}�Hf���ׯ$��z�d�#��VD��<�����îݸo:��÷��-��,}�d3��,w��U��Wu���cb��7�M5p�PX��v��役X�Veմ���7
p9�v��J�n��Cy�ng���_::�����ec��=�7�$,��l�_>WR���=SݣeQ�]��*m���â��老��yO{��w�}�%A�~.\%�9��g"��8R�X�Ej.�ı�P�g<f�]%b����ޘ0���f���ԉ*��t��8Ƹ�᝷"���r�b�c{���r�M�!��@$��v=[�,�%5���J�����a�l_�ذ��g+�f�{�J����כ�.�0���a3y����ӓ��p�:�G":��p�LQ꾡y�{<r��^���e6��N�^I���:E��	�[{Bt4dלbzШ�dM>�7nLə�6�,�q]���.��IW9��oe�u�O͍Wz"">�/��S���Q��:P��	z�nN�>�r\���Ծ���9ˊ�q�l��v�
�i�R��3��)�U�8���9�O/5w[l���Ô'&[��ҡ�Z�Bjq�ћ�xG!��<���ۑ ��C��͖;���=��q�e^�s��Ú�ヴ�Uk�z�E-ዌ郟8��������K|�����q�lg���Q�~�j^��\k���ʋYUDR�$P�x}�iZ��OU���B�}�+}�R�\rz�S���K��:�Q��FOzp?p�sGy�KC9s�M�ALv��ظT|�soLV�b��r���˺>��ro�/m(���\[�r�K���F�Qm���0�s��^��ga���w����l������퉚�.�Q�Z��P�ʰ�k����<�ìk�eՊ�;{=��/X����O���V����1��3�
؀�.+��fII�-(����fɺ�6���{�͓iQ[n�pN�u�`X����	���Z���L�4�s��;��ni�wPc�wa����N��G��N����N��ʆVQfƚ�
�b�b6/��qbS����Z�V�`D�MN�=��~�����궚ךm��:�*�:4�������{_6��X݋
ah�}C&���vU�.̗W�V	���T�����Jx�5�5�u�ܴ�E�59��v�����WO��l�vkE|9�����/��Gn7�	᎐�&j�����u�[�Nqs����/�Z!c��u-�4��[Zz����M�u����X�����T:fQ
zBT4)����"�x��⎐8�Rb�{�����f�|�l;���R(�@<�\��w*�����L��L%�C8�Η��.a�'�y&'�q�Ѹ�vD��yVy�9�z|i��:�.$IH��X�ZÚ��3V�˪��'F�8sI�/g��E�Rkq <Q�] �8%�'޴��VeGS�ټ��i�R��8f�yNu���"r?f�N1���zik��}v�@�Uo�$�qڝE�'eK�:륻r`�G��[Ƽ5��DE��̫�t6k�sφQ�LQ�g��^�� �o za��d�X5��ٲ�)z3��NLj��b��(�V����~̜ɾ�uMd�wy*�Z���}$��R�Gt�y�^��̉���,�#~�[��">7:�GM,�y*=_�m:F�3+��`{D��D��끊*��
24ua��t�P�.��n�H~r����i
z�C�[�=�/�e�^��MpqK#wToh�]���P��!q+�\*�ۄ�Tga�c�`�n�w9[YV�fV4��8�ξT�(��[a�����CU힆���W�Ƚ��Ot����U}�瀰�N$�V�)j��[ˌp�cyɧ�&�eS�h-Q����rk��$[Z
[��I�w�]R�\��4ѽT�}R���n��^�o�)�nŅ?/���#��7r��;���Zf/�u��z�:�X�q���ؽ��K�J��﷤�0�A�cj�����˷����'����������Y�D)�:�'ڔ_S�6��̭�k��s�r�G��Fo&�2�8v��w�Ui��מ�|����[I����1C�E��n��[5�]'����p�\OKfd�T2r��%Z[��<�Ǔqe�i�xG\r�"k4���w7&H�цr�y��b����'�{�e� �0C6�9k�ˆdp"6��k3df[
p;�ҜM�X�-�T_�U�}Pf��謕���#5I{s��Ρr�Y�����k�nç9�m�8�ug1�a���+k�`��|��յ�;��X��c�ﹹ���+������С[�3t�?v��]���y�����[V����6&j��w����YM*���.3��U}�ֱ�/d]�n�'�����7�}W�)a .~�!�e�e�o(�u.�����gݚ5u��@K�MX����۶��uH���-q5�;���r��ؓ��m-#'Y/�+����GS��^���kq?�7Q78F���c� 9�a�?w�f��=�IH�/oO�i^�C�q�U0*�S��F��lS\��O�p="��bWl�|ݣ��ވ=�v�f�5x:�c�f�=v���e	��̂���*�ƶ��y�o��T�f
���UiW�ʐ-�L.��*l�t�g6I�/f���S���1�&��腮���\b@)��՛� ��uE��b7z#�r��H�;�e��[{�*5�� u�;����DW��I�7�7Wu���8]gU�<6:r�n��8KӖ�CWY���V۟n��}_UW��8��%������|�xR|�˶�]�S�u�������G����C�=��*����Jy%�s�{�<1�W�ﷆ�g�G{�x�;t���u����-�z�e�\B8��7�*!�;_9��Z�-�UKG_=�M��pn���8�[�694�����woD�e����槟�]�Z�s����(�	��{-�o�vh�]���&��X�c��mv>��';:ᛅ(_R;@���?�7)����u��1���Ѭ\j��st�R����i��MƻF�]�1�l�[���ިK�N�I��{�����o�9�t���ruK9M�͈o*�׆u��Z�H���#*��7Z�I�<�y�y��^ջj^�p��6��}�f�T�����3�/$��nm!�1�`]�M������s�;������j����9���C���r���$���V�e"��m��䮞������S"%[�n_�O���`��u�g��*��*Y6�]��B�Eɶ���]�fd�,f��b*��W����dmJ5�{Yq�oƋY)��p;z�kh�(Vc�{�2g	��J��_W�}�m���sɣ���p��.��w*-F�d�{Ko�[�lImu���W��b�̔��k\�����6�z�߇�g�>����w�ia�&�̛�|��R�A���Ozni��˶�A��yB{*����A٣5�'�ۇ�ym�p�z�_!]�,m=N��Ȏ�=:���Ž�u��PSR�a|�]?���T�������5���������B�.��T��<�*�{]`�9�tZ]}t]JZiJyp�[x����0.��tcƱ�ƫ���/��pGs9�v.��>4��_������(/����ӽ̦�V<�;NQ�D)�����P9��+��MH9�R��u��,�-b�7-������,�"���zf'��20��N�ͧ�bX15�mG>t���;a[7�O�Ԏ�<�m��wNaf�;1�:�.3���߫��~ؓ�G��z[��}8<�%��̊��)Y��q
�/��9���+3^`w��&>;産I]h��<�_3T�=f��|L��H�q��Eœ�W�9�z���o�uCMee+��޿}�}N�lQo��r|��Z�����DrLSn1�#q?'dMT�x׫7�5��0s���R�<$H�.�ͽ��v��N�B�i7_s�uy1�^��>���A�9	����<|��7�Oy�]��2�k���6���%�\�VN��T�T�?N������;S����qH�X��[뀑P�=Z���n'�kQ�޽�H�GE��^�����+h�����MZC}K���_io��j���<��x��<ڈ�{Q�g+��3(р��\�U�B�'%+��}���'%�q�׫"�Ϻ>�?gN��bg���������q��..��*��|Sf}Q�����j�cb����j��>�*�&��;�b�v�Y�k����] �TI}_m2�媔kw�Ἷ�ْ��;�����v�3�i�ޫ�A�B�=����.������&FH���\1>�;=�
m�g�<��^u�u����m�.7R���C~�x�.�57 	*c�t�\�2��I]��JXa�,'J͓�uV���-����u�u:�HL�ֲ�h�:o���db
ĉ��8gr����Z�~��g�|>�\������gڈ��Q	�w_oLA�X�唶�	��w�n1i�ޢ�Ju�x�q��OʗJ�1�oI�BZ��յX��m��|{v!��9�Z�������I��Y�D)�K+`��T��qF=7<�p�����|zc�FTF�i��þ	Tt��ؼ����x���S2��v�/(��Jv��[���o�r�RL5�n5���j�����uԥ�%�ME�5�&�
���&yi��Ow���&��w�F���){��ϵ�b�*�Q/2�7����6���T�Q�~h���9[q��/�o*�^�c������[���z��5o8������v
=�Q{N���	8֟I�Ǔ
h�b�y�Z��T
-	Y���v�q���U&o�D�c;TJ����vz�o';[|d�ZC�z���޿x&"q$wE��]���A<���.P�͞:W�/˚��.���ՑP��Z&0nhk�����Y�k����3�i���<�Bs �s�	�ӭ1d����2ԍ�a�X�S�+����x��=]�dQ���0z�nr��Ung{��L5y�<��Gw��������DIO��;�61��O�M���(�oY�Q�����轻�#����c��:���N�5j1�ֵ���{���7�o/M�k�f�����pr#+��}��MX�qQ};�C��.є�Gu�i��On�T*	h��Q'�e���l�9�]��h�K�:��|�x'�8�n�XJ7��T��_�=F�#�
Y�5�(��E�/WZ�A-(�nֻꇂ�J$(�1کr9x�L�i�׫>�pp�hT��8������q�[���x���Lj�o���ԑq�wR�mh�1o>����	�V��⺾[�i&����W�P�2�\X��ƫ9�n�T:fQ4I�Z�'��Y�ks��[�{=OQ�R�4�Cq<H���;upƅB�;�u��C����>�/}����Y�r=�iAa<��W�H(�]Ӡ.h�I�va�f�^�&��H-;#׮�ݽ7w$�̬)Rv��j���ltKk�M���,W0�l-|6Y��m����c�a?ko$�X����[J��%�Ĉ��Ս��௥p���pɒ�''b�Vܦ(�+k�u�"_L����Fl��������a�DP׏�,�um��^�7�ľ{g*f؏-��1��
� XD��"����ݦ���hF[nps�t�_t����u�ܫ�D�`���婹�m#���,&s1��0��G��T�RU�VpW)E���yT��y��|�"�j�<��W�.�ٶv�La�E�䫶h�QN�]^l���3T�+���s�|�l׸������:��ٴ/��f �@^\�A �c��2���9���������q*N	�f��[Y�2���r'2�s�a������.=z�jEn��,�\���nf��(�҄���#��o!��\u�̻����b���M��lM�R�n�E��ó�
�U]7�aZS��lF�T���]oR�4L5�q웛V掺�i��[��D���ӎ�<T'�jS}���\ݺ���IF��V,f��V�8�skb�6���}G�iUгt�u�YM��^Zq�ۜM'��$����Gp1{s��mn���̮� "�e�����y���0f�5;���Y����5gl��A�fw�#�yH�k=r���aV�����<�;�{,kZ2�hM��,|5��-Ӏ�oK�Vt��'�4�ܨ��܏5��w���#�h�|d���dLل���E��v�B$�م%�S´q�`�Zqd��ʝV �Y��8>�ϱ���W
o���`�gQ�������G��+IϯR=�^�⏦�qf�Ր�}��`������HS�����Hh+E*Y���XWoT#R:����qV����.�-
�2-���ݰ�q(y5�`ՖW��p0�����ۺD��\U�$�Kt�x%c˴�˩���V�"��Kz{�<�o�sw��g
cnK�<�TQ��^��Sڻ)��Tx�L'���L)�ϑ6Z��}���	vw^��"���E�X�z,�&��ge�QS���@���A����t7C��]��#{Y���E�J�̷-;k���gV�f@�ۊ����ȹ��}�B��TG��Bl�vٹ�wE�#��7Uh�ȕ`�]�xè��M���K�z@妮ˏ�]a�]ټ�;�xDUǹ�j�m�&P��E�{8�:ҋ�ݓ�8�ҫ��j����wN�i�uqv�͕f�
���ۏ�Q/N��_s�i�Wvڲe.pWrȺO������R�z�;���Zq�䶭��n�ڽ�ӆ�i�50j�ˬ�L����Wf�7��p��nt��2us�:�P�'op��n�r���׬	=��z�7�hݔ),_.�m�R�*��A�("
�TAA�*.Ub,�,�D��*���	$Ӓ!3����)aR�r#P����DZeȢ�8U�ʸDr���HAL���&�S:��WMF�$��ee�QV�@A���J�E�K2�P\-If[��U��eE4�����
�IСD��h��*!Rr�#�N�PMX�(�Q�����4 ��eG2BI9UR�&rq��Qv]�0D�**��
*����M�ȸT��I�a��

"�L**�����"��AT�g.p��eUG#�$�\"�G5��eA�q:vQF��DETfP\�ȕr�9W��#�t�"(PĪTEL��
�TT��s��H��f�\����ɗ��u@U�G%(��* 0 � A& �2c/��A������{��/(\����m�h*4�����# :6;n�
�ј�2s���b�B����|/��|ֲ�"�V7�B���'�j9&&�7���dr���wՀ,ZdSGg[��/�������{_.�W��B�i7j!��~C�_�
=f����^�ӽe�����{q��}{V�����xMd%���Fz�#~wp+�tzp�3G'f����Q6����2�]cO�
���=h��<���ͩ��A���K�q�}�g����o��P�/�Q��(^��o�����nL0��������U��]��-�=l��,9�V{2����p�-SZ������_1I�w�KO��[�i�ȃݦ��U��:�4���΄M�	i����Yp�|���z��;p�|�����H�N�j7��V�=ӽA��_TF�t��J�ky=e�i�����l�xq�͞�t�iZ��1�����B�����%-5
S�i����ߔ�Q`��E��+���i�]��]@���/�<<�stjʦDV/��C�Rw)V󥸖�M��q�Lu�w�TL	������V8�v5q�\�Εϡ˷��wT��XU���z�I����B����S�������f"��rk������W�'���.N���M�]�6����/Ϳ!�xgQ(4�r�;��ϔ���{���}�)���݂�7w�Ң�Fav븗 f�6�z\,M\3��ca7��e�e�m�<ǚ�H��ɮn����k�7��)��Is��|:a1P�)��\9��(:���E�b[]=E���|�����a��n�s�>�\�یw�MWx�h��62�R��tjg��{��n��N7��{����ѯ�8r���n��s�QM������c��sE���Y�j���u�?ENs����&R�:����k���)�V[Փݍ�U_��V�ne	�я�/��� 4��� E�����bo(��z���j!�7Q�fQ~�������Ⳳ2�������ob�X��$���G���sy��;&�f���p���g�0�k�5er���wS���r_3��.��*8�Wu��zy`T�.ۙ�)qWMN7��)������7�W.��]][۔���j,�һy���H��@&�?�����OZQC�;4���@S�s�[Ԝs?��{�%bĻ���زo�:���K�u��ll���az)�sR���zH�Q�qxx��7j%OV҄������-��)���>��鉑�-;X����iauZ���y�6�P�R��������N�7�W.��l�qԞ�)�W���l�_>W{�63����W$��;�j���w��zվ[m�	}��A�*�v��n���f*�u�����<�j�ı�O�u<g*]%@����xC�nb�T��b�C��/s�= 7��w������-+�sV��)��!�(_T�s-�9y�d�~�Y��wf���-��&���8v�n�@vR/�)��yv�=+BU��v��s�ͦ�\�o.f�|�^ҥ�ws�'V�Z*|n&1?s0
unJܚ��qܶ����DŞtZ�xq#�̪�սI^voMO �AL/%b/�U޵�À�(}��۟��zs�o-]�߫�:�����]Ѩn��<=�)v0���u>�KsOK�
f��XS7����|w�S��
�|�@l5����&�پ�@�oM�DF��|�JԦ���.�%7�4���!�-m@v�UG�6��j�!n����`�����e^�'[x�2���o*�^��c������eX��s"������j#���6���W�nڗ��kY��F<�Uf��C0[u("����"��W.g{/i���/����ڽ޾6�.���~|�3\�#*f�:�f��pfTAۘ��̉)����;y�c"c��f��U<�9?����h���BY��;T�ep7�\�N�j�k�ؾ�1�&�r����}�ޞ�{�{cf�ܻ~Q���󁨇����(Õ��p%2ø�Y���s�7��}p�=�S}Q���m�~�8���o��{O��q1�4B�Q��F����YC��4�*۱aJ�9��������׵�ծAC�`.}}tYKN��<�kZ�|3��r�m��XW��U�X�sIE�әhT�m�q���lE�X8��[��}�K_u ��܂���퀵G��J�9�dn�m�)n^/q;�t~�
����uۥZ0�w@oR+G���}G�˼�Y�*�f^;���(R�OT�w�I+�E�QÇv�@3?����[��������;5�9�o��'Ɯ��Gk{������ӈ��,D\�.�c}T��������KE����+����&����@SW�n��b��R+q�pW���GΙ�o��wo��|;�2US�eS)(ѵ}X�cg
J�Y��o���h�Ms�����6/�g����bc���m�LgY��-�\ï�>�_rLM6�]�q:쉈�6-j��xu���*Q})5�b^��#U���I�ޚx�;�6�8s_&��;��xE���[�S�Y�Sڸ�HpQ���J̩篷�/����R���sO(�T.�U�ь�_'�qm�q�fދυ�C1TD�ꈒ�e��{)�K��uM�+���y[���nl�}����*��4o>�u�1B��B'`�P�kKx��3���I�X��5�q�:��6�|.�Ǣ5���?-�ݪc��{T{򗶼�xogj/���T�k�ܕ����U���
w��L�c(�y�)�+~l$O���J=�#�mz��h��^��x=ݗ�2�HNJ|�P<�W�E&˻���&%��&��,R�����\�<�ud�g��D'H����n��=�B}�7�Cz->��K�\*������Z{���N���c����D��fym��c����%:t�+�l�|-!�����\�ʾ�]�U��5́��5�Gkޚ}l��+d���ڧ*���\o��C���Oum՗p&{��u5��1h �!�)u�]R���)���kJɭ��\5m��m��Ut��,p��t������F�I�K��j���3��{D�ۦ��J����*�k��/8�[�\7tzG{s���ޒ���"�;�k�]��Ϯ���sR�gp&�l9e �����X����2�j\Mˉ�"�B�P�5a�÷||vp0pqh�=�2L��k#����NoME���M�=��a����SH8p�������V�W�Dchv0�K�ˏ�9�f������p�\��v�hr�ne�Ԣ�i���Mɔ ��Q�k�б}���A9}L�̩8A�yf��T�ܰ-�ָ;�糧�7Y��Z���U��E�k.������@��;��n�e�*b/W��,5�]��B��_-/�ߣ讜J'z�KB�����"c�فq�Z3s�,�����duϑ���Hm*���.S����9��:b����m�DO-ϋzv�l:mH�����mΧ�Ĝc���~��F��c2���3�}'v�C�I^j�j��]�N"N��\OՉ;����K�֝f�kΥ�-�֗[�~�F�&�魔���U��np������bB�jAO-�U۷	�de
W�n��$(�tچo�6�'_r��f҄�l���[��DSMvf�c��o�	C:z-}O��^��3k��@���yTD��*
�Z�_�[�R�%�T�����*):P������oy���

ah?AP`>D$�:謉��]��1���얷{K�o=�������[��}	}��AP~�(bεkfaؐ�����u=��j��>,���-k���:�x�W��(��;��O�ެ�@��b!K�,���E��z0��p�����&�푷|����@d���O9�N�q��Q��,^l��.����X�D�ʷ�o7݃��n�Ȭ+}g���^��h�a^������Ni��\���K3Z�'�o���'w��U�.����.����չ����Ʋ�ml�k'�h�=j��s7�d[�������DJחR��7�I2�8v�lӋͪ�*�]d�U�q�Zv��ᘄQ�g�A+\�Jܚ��P���̺.1����:��v�ɩ��J���3[7�&9�:snMDM�ڸ��n7z��T��U��"�T��Β��bjq��Fn�^1�t�-m|��s3�H����;��q���/Vv�w����Nv��o*�^�;E���=��>�ާH�1�����բ��f����'�>�Տ*�Y��i��ҽ��UUʍwrwI�N37>�{R^�Q6��*^�X��V�h�s������˖9<v�����P��_{/��2����9�`v�צ���;cc�]�\$��_r�=�}qm9��7=�kW���urE�)V�c���y�_q��i����)fj�I݃s�����֕'�
�QӒ���^n�����k��v���oS�=�������s��\c���u��:y�¥ݹW4��nC8�h_�go'��,ѱ�B���Ck�nv�h��lǪ;R[��W�v�Y�wk@���UD���l�E[j��b�(�ɓ�Ѻ=��yZ�p51P�7��}n��S}K���wo(ut*�A�N��79Rt�����Q��OuM�����!4��n�XX���4Ɛ������$iwT��JZiJypֵυ�<ㇱl=Ҩ5�1ݥύWE�(l���PKE|9��Չ񯜾����҇՗:�E���˛���u�v��r���S�R4;�����_I\忰ڢ]�9Fr��9."�ޜ\���Q	��,�ȅ�,�h%zf�4��߫���[:�[=���WbI�)�l;F�~T��#�8�5nS3�3Μ}��Ɏ�г���Ut�0�>�Q�14ۍw�N�"yQ�im�}��wܼ+�.�ON��F��Ȝkj��[P��_ܝ���n����$!Z�g��(���)m��������"Y�M:?;�l���鹚���As�n��s��X
��|�N����9S�����-�s��N#���D�b�^J�KG�sQ8�J�S3s�1X�W�ŷZ1��귉[�=q'P�]y�N;Au3�Ok�ce����~��쪳�j���Kk'?D��٧�5/n18eM�{�R�=Ux��yq���o�F�-Q�D���/����]'��hh��6fj���P�A�oZƨ�F<څVn�X�
��l�	�;���SȾ��y�z����5}�˞lc�}��ߋ�-�����q�����{�zC��y���u���K��c�������r��]�'��;����]<˦1gV4m�:̮�K�`믤���k�l�@��v��O�s����N���k���C�r�u��8/� U'�f\���F�|�5��=���v��TYb�k�k6�Q9O㹪Ň?-�
�*�J]q�E�JZQN��t�� ��k��X]����yN;c���ʆ黁AL/���I�ޚ�2o���C޳;��=UҚb�g63��9_9E ���-E,�(�;�3��_��F`��{&?�*���ɯ:���B�)��ݫ�}u/�t�ާw�,f��;a�0��T�N 1s�>�W��1u`���8���tZ�쓮�����r�۽lXľI[���:Z��jV�X�x�	����h��Է.qWu�ïy���*��P�t�Vh����lv����y�D�V7׫c�C�c�h]wd-�1���g�o�����jm`��0s����r��_f5M�z#흖�D��>�G��>�h�~��=���I�X �,����n�}�ӓ�碎�I���Q�xr'V��;Wó!7�k������n��j��c�=9�I��G+����M����앷t�j���;ϴ�E�es�5j�J����Ytzh�9�sr�lo�@��|���;"�WN��d�u���ӱJ���Z5N �ޫAo)�Ä�x��P	�v��A�"ˮ�8�6�&w>�BZ�&33K����isf�v��U����*��]�	�L��<{Id52>�t��ȨV�9&�՝Օl�O��Ilfq{�{Wґ�07�.0�;7��
�8�z��f�n���e��y���j�yl�؍/E7��I]�wq�鎥�0k�[A%�œ��s.Y�|_�S0Vk�<ܦ&��{q;�8�ҡKh!k~G��N}6��j�05
%�W["�)����`͓�2B�j�U�\�YE��_��j��Un�wܥ���|�P�\':1�א݂�I	���zLmm'�2м}�2����s������xQq>/);c/�kgk ���Ҭ� ��2�x �4�]�+4t6�*��5a��L�Q	q���
�{7lT��tj�K��Ϝ��-�;N=7b�`ݐV�LN�^W=F�<��rc�rK���8�W4�p2��Qlr�cN�^�Xͺ��\v��ٱ�r�N��-0�y-n���Y`T�B��K-���15Oh^�%� I���w:
-Z��+�����i�
���Y��5���(�2��p�a:���\Q���M���v�gfuj/�8N����X�6���K���5�G��ڕ��MD��S��T[GK̤�A����{1��t{�[��C����+0I�`�o[Z��i��X]W�`T��m��y4�,
Y�#�<��@/���p&��2�;[J��V�z�_u.�����Ċ�MWzw;�˃KxA���9 t�W)u����N�7���&3��}�h$oim6��>1��U�8Tc��Gf$�Bs��B X�sZ$��l��s�
�w�큷u�[��s�X�<�v�"^C�5Ir���ך��R�S�"q!�ME�]�W۝�{�]n'�X�ѧ�iR�ym����:�/~8!���M����A���B�������Mٍ��M�W�s�7��7��;"�CG�y��7�W]͹��}�BP�{�v��6�_WnJG�p�F����/����B���S�YEeˑ\猊VȎUPQ\��Ґ(��%.��9M��n$*��"�<�8�g+:�#���E4H��:�ӄܠp��#�RZQR�s�N���sA#�q'"�ex�$ʈ*�&\��R��%�'T*"�ȑQ��<l�	�dW@�0����EDED�t�2�"��Q:�T�-�J$©�TE��`��Q[\�eU9H���Tx�
���f�(����zl���Ud�q�,�H���r��t�.T�s���OC���W
L4R�]M ��^q�9N7Q**�t���;�L���'�5��'#��̎W*
<e:����(��q����G$�kA2dEf���7)Ȫ�MBP�"q%+w�T��0!*)
���18S-q�9ENA�(��"�M������������$��gs3�8�)^��wW�ձ�b�B�ӈ1��˺���6>͹��v���n�I\��������q����5~�wZ���9�c;��ci��r�;���e�Rq������Z��<���U��P�5p������(��ZM��kf�c+3c���@)PW'�ME����:��:O��L8j-Bm��ǵѵ�n-�܍q��jgY��l*��2�9�f�������ԥ=�ӄ�P��>����8k�1����tc_Z3s�j�~�rڞLgs���t^:ѹMn�����7��s���s�u�t[�[6����L1.9:���b�
p��^�az��k>}G�=�ڇH�G1��ub�=��M������z�R�9*�N���:+al(���:͸םQVs%KnÚ�[�,J���pU��M�W�Uz]Y�]ע>�=��퍜}8�o��5ȭX��̩q�����*�U.z�iBWe�د��zn/�:E�۱���yt��Y��/_P:����ik
�c-���xvz�)M͋���ݸ!����;c9�8�p�
W���w\Nr��i����|3��א�%8e�q�Ϙ0�p[ϱ�t�o�W��d�E���]⧵r;�M�w���Ì���vОʱ;pzk�-R����lf�H���.Ѵ�oBYq��I�5ˢ0��*�v����V��n.��e�E��rs��/�ִ�������m�v����}�0TV=j؍�}��Mm"5.�䥲ޗ_e�Z�c�P񜨗I_b����p/P�.DG�??��P�S�w�⺢1>���J�g5n7�*-������.u���.񵡏T2��)���f�V��)-��V���\�]JOˍ�W��k/��˅H�Y�	d
�5��ɭ�k��@���M �4.��Cy�#������]�q*���6AN�m��9|��7|^b�m�Q3�.Y��y+�ŝq	�5I��#7���7���;|Ip�R�9{�v�{C�cu����5j���<N���yU��'�9���k��Wo�����M�x7Ev c���c��K�h��{�g5/IXp]�xy�\)�C�;q�H_�C/�فyb��I"�fe��h�c�_Yx�;� �%�;mCwǌ�N����&�13���4��#�j��c��X!Λ8j�Yo���ŜV\�s��Y�VeO=y���[�����Ƶ���W��v���+ێ��=����r��e�ۇ�k+F>���{�~�Vjr騇�������PN�2lg�h��O�qʡ��J+h��υ�m���ڜ����{�ת{����1���!��SiD�����,8<"���6]��P�n�
��/�t����Z�O�܈v���]�ծ�û���P�����Y�b��m��D�>���8)k��[yp�}p�=�Rf�Ўڭwo����(��ɉy,Z�q�
�Q%�F�Q=�j#�{o�YoC��4�*o��,���25��l��i�.��p0v�bK����KJ)޵�E�j`��=�|�y������\p��k�HK��*�P��q�ub|Y}�LkNa�EO�q�J���
�����_<gk�(��w�H`�R�]p[{q}���w���Gb�R����_i=�'��1�,ۛgh1e��ttj��=�֖�s�X�-����9]��
� ��&B9B���学ޠc��:q���u`Z��1�^�E-Rj��[��o>u���*1]y�����B��m��s㫡��!)wsR��˽Ƽ3[�w&�+�L�ȅ1Ҕh��KjQ�Iu
[Q�3/n��3�7��)��	s5�&�8t��n�qԎ���`M�S=+O�2{�yԱ�^l�|��'�F'�j9&%��������W�L���9�þ�b?B/�Um�ߎ	5����[_.�\��n���7Ԭ�Wf�K�a�x^{���ߪ�=���+���y��ƽ��,��u��ٿg�/xn�5�zT􃴥����%�|������� ~j�6�UoR���;=�ᷭcTv���ʬ�F��E\���nq��:���#<¨��/�;[A`O�&#�s�aD:�ɭވ���ݜ�����߸�a��ˉ֥�OW�d�R]]_LS\�-=�]�p�*�ð�a�xpz�/.�=����ưI�����nz��;W��}n���|�k��0�4M5{�k|�� ��+������yeR�u�s<8�.�fn9��	�3�V�^�r�E���n�A�OxY�ա�1�5���'�ve���k��g;/uH	�(�7cK,�n�WN�WQ�u�ѼM.�T��(T�x��m.��#��b��������w.�CX<���W[U|�B��=����
b��A�DIK�#��������wt
����]c�>��㇝o�T7Mą���*I��%�1[����:�h���+����B��h����uC�q�P���k�7�(RZkY6)Nz o��=~�t��g���}ʡ��I���D(�y��X{k��_E�|A��<�Խy|Z��6��|:atC7=�+{bnz��+oR/�������
�{�j�sQK�o��N�|��O��L9���ݹ\A�|�
��J��7>�V�sne�9�j�V�玩mfa�����fՔ�V��J:jq��*~"���yVc�Fmg�ڥ��1o.��tCǼQ�ǆ��ݕ{��tbp��s���G<7_k"�Fb�0��F����$�m��
�Wu���'9[J�03l�#F��Q����:ԗ*F�� 5�&���t��u��VI��̤� *�v֎3�u��n�W��T����ލ�'k;�(P�)4�cl�����uL�3R�W!�g�4��F�q#&I�;��o�Y��f�y�״��T��IƵ����z�Q�fM/W��)���r0��o6s35��b�T��I\3�GV4� ���v�����ϻר��8������{C�{��U��r���'v�3�%���;�K�<����Z�
�L�2�<9T�9н�Ǎ�v���g��x^���v|J@ó�z��W����@7�:�x<�o�d)�ЦzJ���-���^y�C�dD��ɑ�<I�RW�*a�>G����T`������o1ށ��s���/U�9��G��7��r=n�;"e��%�9�I�X<�*ft3׏Ws�5�����˞�eԳqO�X�����}�'�����'ǯ��}�Vx� �p@�[���O^o�յv�0=�A��</�t�r��Bo��CF7޶���'J���r}T�/%}���eT_]ʻ��>ƶ|l������I�)̄e��ԇ��3ӽlv�Ը��^��S^���Y�9O1�A���ډ`�r!ΠO+��n����F��|��	��>�q��| X �x!�E_z�gRG��V�م��;�ER�Ú�%B}LC3�R=\l�{�eg�Y����ԕ��ʉմ��$��z|���W�@��۝:��Z]��,yB�UG���YC_+d�	�&�3�E^Ɲ��sܗ��{�'}�ZY�'�}̟��>�ogEU�����΄M����.#��d�eo��l�$��*(�;W����1S�v7ٽ3�ޫ���r}���@����|�`���Y<(̿��௥�h��ѳJ$�|i��8�zU�i���w	��7�����?z��c5C/�lɥ0ʚ��׾��VM���o�l[c7R����gE�+>ާ��ˇ����ƿD�K�τ��׶o�>�8L��%X�y�L�ڜ|�ć�/æ�mh�/N����z���u��vFk�����Ҷ����
}+{��=�Xc�+ʜ7����wL;����u��.� ����^������^���#=3j�Q����\iS�/~��r���	��mP���T�1���k�;���.���s�lbT�w�;������o��C�/m�>�X�ȿ�%%�.��]>�����-�z��FU9��q���l����u�n<�x���e��~�Q��{�\#�xWOl��Ý\bl�n�eT�����T������	r��A���7�>>ӏ��VG��{��"³,��!����a���Sq.͒�����,�[��X)q�r�m�S"�0�����f�(�}��H�"�wеBYH��=���ޔ�����z<�@e���=�ˤXH�jEs��´V�We���V)]	Ydj�iÏ �m��i���376������y���ٮ��;����|$�Cz��J�M�z�8g��1����Σڶo�,� �����=S]cӆ�d�4�}Pg�L@)(�[S�.�}t�p����w�W�[~�~l�k+ʪ��wю��+��!r|i��A�p$�\H�Z�/uD�V�d��H�=G����������h���RM�}R:�T�ә.P 7#Ď�n��_`�'J߽3�L`��^Ӌ�z5�}�B���m��}��=Z�z��ߌә%�U-������T	�SѾ�]�Q����O�W�S:7!�l�>B��!�~�o��O����5�T5<H�|�3y+���P>��=�~�mn>>�^�e`���F��n�ĩ�k�G���L{�߬����o���C]��VG��_k+i|@�梃���7d��P���oFDV���ަ:᫼gП��\=�T���J�sP��^`���%��	koG�� �t��C&_�wL+��n����>[�Å�u��t������N^�G4�s�Sr�G��N����\G^T�҉̀p&n�C��+��/I��=�I�\��3�.�z�@�E�φ\�M�������M�K�ӠF�Q�*�;�v��� ���ɉ��A�
�lj�5���"�!ܫ',B�u:"�r﷨��\m'LHi�+�;u	���^�c�Ds��>}|0As�j���k��ES/!�kgM�N�ظ�.+��DO����'^�>u1:�ۜ.�IS�_9eϒ� �[�Gb���)�5��{Ӿ��ύJ�,���
Z�ǳ�sK���w�g���%7�Ǯg�zN�9S���/��:g��n��>��3��>��~��S�g�+���y���9^��*��~�f-���gܬ�ۇ�[�7�uzp�,�/��p;��7��2㌅�1�\-�܏z���p�K�vfVQ|�����`��U�ŵ�>48����PeSJGc
ym�q��`}i�|��
�=��. {0�G:!��1�*%� �d�j�J�3�*�Q��ŗq>6�D>K��D˫�w�R���J�����'�{7�����Dmǽw���l�9N�I`O���:*�0k|b���a�����֟[+�Ua3�E?+��W�"���{�t�o�Fc|����X}6j߱�F'Mź��~����y��� �P��h�F�H'>��x��E��Jn���^2�=!�ʮ�n���������I��1'�M��=㸌�;|���m_�}�g� �sĽ�꽶ctY��6bE����a�YMM�ڇ������ɥWc-Ws>�i����)[j�LkV���Jl�H�k�-̡��1X��4�/�f`���F�D�ƥY��\��O��C"EM�KBVZ�`���9�c�Ф�Pme_<gw��.c�m_�[X�R{D�{���/��o�k���=q��~Wr&�(E����5��^-����^�_�l�5g�7?e�5�OW��|G�c%�n�Ҽv����s��	������[��S���������P����0do{*A�������
�պW�7�z���k�ތ��X}R��u��ϛ���~�=&���xWg��e�G�3���Q�9>��ళ2�;�J:�/�����V׆�W�q<sz}�q�n��.k�c!�Ew���������36GF5����ȿ5��m$w9%t��.W�e�P����:.���܈]L
����.W�����o�ϟ����=Ǡ_C��|/w�~��j��c�;ʟ����;�Ǯ�aEd֛��@y`�`T-v��J�l�z�z�ɽ��܂������*�[;�WHw�=�/V��>%+�0���+�H�u��T<ӓ0}�~)f��R��W��>����������%��L���O�U���>�k���Hs��͎�=�%��;Ý{N��c�\?)�9���-��.��OTL�}�tzl/C"���.�J���[|f�ެ�u7����}��g*�cA��HڹM�j<��N����s�]G�ڦ��l����A>g��y��p*n�kA]��)P��[n�w�n^��D'Ǌ
���m��n�Y��K �;_+��y�xS�0Ԃ�J�cPb�1�a���� �'i-(�p:�i�؛>hK�E�1��żeEO�Yˍ �E�@����jnfq�%t �l1+n#]L�i��7�jZ���Z	��[�P��VO�vk���5C��m9��=��yɲ	��/�ٵvU�����!Y��x� �R�n�f���Ҳ�#�F��T���{v��DP��G9�Y�]�|nZp�(}}��Wq�5�wP����L����м���]�Xe�\Ti���]��3]�4�f'»@�h�
.�A#�;5^��F�'���%��h��wӂۋ�b&�ϩe!P�9�f`�Z�Zr��Pći�I�U���3M�o��r�9+C��{�5��Lp�2�{��g���v�C�r�m��2� ǻ��Z�Xe3ɑ��ǝ;w�#d�E�����1l��n�h�6���s�Lg�7���n�+f�B��OcJ���HYKn�J\.�Dڑ�d��cᣝ��{��x{���Ňh����v��)%�,���:WZ�=V+�-.ĉ�'v�.�����>7�Nu��}�L��;)��퓒�y�9����oy	"j>̥iPO��35O�������(s~�΀u�Y��S&!��L6Ե�8���Y� jK���H�i��w�ka
�S�뺍����Qo<{�$(dJҸ�*Z�uumn��N��+J�oTB	X��X4Y7[���
}�S[k�a�æ����9Mn+j^�\x��n!�a�쥗��CP��ՙ��#cU��Z�
�j(���v
�[�ʙ����z�3�(P��g5��1݊/f�rA��R�t��mk�e��G����ѵMb�+0����b�L;)u��rw���m���
\��틔4�bZ2U�w�!6(�A��f��V��+�'���9��;����P���}D�!�o��I��Y�K���ݵƳ8�	��$��U���̪�[���9]Je�u�����ܥ���d�A��jS*�u��#���DʭW���L���f�~f�{��d�o2�����B�"�9�3�/���\୧�:����Fd�уJޝ]b����q�qY�Y%+Hf��:���޺�,�N��������͹B����F_RC{�G<:^6���ޔ��i^�厝�zr�ۨo?]JX��am�ݻ�M�&�#*j��+�Q?�c��k^���LX�!w�ځ�uj�ᨹ�f�`BLs�C����+=��������9T�c���q�s/��������h	wZ��N,}N���o�v�co-1ǡ��E���-V��j��?W��~p����X��)�J�2��e�U ��Bs�x6��+�㦎'(8�9T\s�2%J�9���\\���7��A*q"`]Č�.DUsVSq�(��VWQb`h�2���EM'QN#�x�Z�7TQAZU0�
 ���JV�Ps�$f��q��ǚBI9�QT�sq��i�4rAy�ӕb!&x˧#Dʬ�,�ҩ�˔fp��/$�r�+J*Q+�r����dE$9�W�*�HN]6QE�K�XQ�k���FIA$�����p��#�J*��PL��/�E�M����d�Je�A+�3���*��9�'�HX���^M
��4��/'�8����eEFBjQuYgMˊ���,I�
��%Q��H �AfYb=�|���üC�����:1����/��,�F���+,G!�^f#����Ԅʹ::h�ѥQ[5:��(grn�������io�yu,�E7V&�w�>D��>�Y�Dg���>�����ñ4t��ޜp��u����:���	�_��<'�������>>�p����ѵ#��
s�>�5��'�f7���p@��7�GA+�s�ƿZdz�팏N����S�8.� >�#wo��2|���z�i�,�"t'���^��t_j���릗���5��}Z{غ��������ɿ��ՠ_��_9�L�Cdq#"_W���_�>����ez'�����,�Eb�M���@����{��x�sN{�|K����2R�\��n,��<���W�����j_����~wrn!�F���y��{��5�Ry�����Qy�Vg�&���u+N�����Y��>6���Ȅ�w�3_��������;e�n�e;sV4���p~��,�4�>��W6�z�}�E�u��DoSΪ����^��5��z]y�n[i]����;�עǪ�l�iD�	��wL;�����Z�� _^�߀����t���-�̎��k��I6d:�t�̃+)�Y�Pb:_;T�2�~Lf(�P�X6{�����_�Ni��ud3� ҏ��f���ܖbN���8J�-	�]�ml���z��l��s�]4d��
�P\t!4
�U��'yV�>�x�o��M�z�\��m~`��YYU���i���'0vG�a:ʭ7S/ī��~�7��{:;�{���VE�/Խ�;�z�7�q���нS�z�|Js/=0�+�7dQ�,yֻN�V}�����3��}�+�ݱˇ��=j�<���N��w�I���%�7^ϻ����C��돪g�b�P�K�M�w�����>>Ӑ�/�z�G�9�G��:2E��a�v�5�Q�S������>�>dk����R��~<���q�����>���Y�C)o�[��,�2�M��|j�J�,	�R$TKjU������t�z3��	��#=�J;�gZ��ӛ�p���������'�Y9Q�p$�\M�+�b�����]��A~����O���1���#��!��}27�,K�2\� �x�r�p*o�߲��F������]���o����m���;��;���o��_q�?�9���N'�h	���j�ϟ8�}WHU�S��܈�>�!Q������|������&��6�[���r��������b����!n��Zų&XuY�z�]�a��;+q�X*!��c�gtooB����HI���w�|�޵�M��yv�����Z�C�Z��wP�=;Q[�WV����tY�`t8kXr�ٜ5��l�6�KR�ɴ��/8t��^@���<�:]<���R�x�>-zH�~Wrb�~�F����;�~�s�v}�Og�`յ��t�2MC,��0�b�1R�ތ�u�7�,k�8O�r+�I}K�x�zx�'3^��v�z�<�E��mH5>%W�2a��
}9�x�>�}��8o
�zo�U�a��xr��G��uS��P�lМ;�7�b��f�No��L�ݨwY^Fy�u�����^��up���oI���Jg:�x3�'�Bu��s��u����ɼ������e��g�Ui�v����T���յL٩�����\{"L��'!���g���,^�F�4�L�����ym1Y`ǧ77��þ(�X�	�
��t\T�S�vX
ƻ�>r�|��?��\o~]=�����*�=xc����ݟ��g�*�,\Tϑ�rjMt������@�s�}��+�zժw��w�x=	N�v�.!��	���\�	n�왏��7t!���-�s�jD�+�my�$%���#��L{J�^RIf��J�0�(�ey��\x=3y�^ӕ;�2��y��t(9�P{C2����nh�$7�#�L�y ���Җ��wu�Q��i�0%������{-�V�N��oh��df��w�����b˂��zE�T�i�%!-�{o���^��b�	���*���<�DU�7Wb����}�yz�o�N��<���do�q��6��dd�� RC�{�Lկc�į�&�X���`>Q���X�9��&���H�s�i^��+�ꑝ�fj�,���w��`]�N���Տc��W��p�C1h޵H'>��?c���fF��Ƅo�=1�*�y��yӮ�z��	�5�5��doj���Y�yσ����m_�}�gơ-/*U0-_�*}���Koɓ�&.�~������3�{TK���˖�k>J����<4�ow#�jj��R=���R;=#Ϻ�.<|yC7�ԃ�Y=P��ϲ���n�����<��y���G�k�X�&V,�	��>���=V�~����{*A�>'��p.#M���^��'�V���>�C������;��Ϋ�|߮��k��7ۯ
�{n�#�ˈ��(���#����Q���g>�̭OW�?�q���*��7���u��g�潦3���/|��q��.�t�_��at��5�Q&�C�3�̳��Nzet{jr����^'WKE�G�r�~�^��[oT�Ƴ�m�vԻ�]u0�V�!8*|3��Cf���{DN�P6�췅7���f��wZ,����M�B(�&�[���w�����'e`���(�bov�tB�MSx�;�@��^�Gy�V1x뻺��y�1`֏���'LQWz5�#�e�*e��B�n��ѐQ]K�������4��Y,�|r&�u����!�\6����y)�
�x�'
�i`���u�V;�;�C��jڞ7gĤ;9g���z���@6�(W�Z�[�:30���Y~Ђ���"�ҽ�������hx,����mH�<I�W�A�P��^j�^w�n_Y����}�x;��9�>��\?)�[�ϝe���]9�I��lv���>T�s'�s����{Q멕�A]L��sBW*��yI�|r=�|z�<�M��g
��mÓ���z���ސx����$9@���x\G;��E{Ԅ߫ֆ�o�m�w����ُ>�����+�w;蛝����J��Ao��%yN XJ5��C��L)Ll��w��S3�kѕ�P���t������/�+�F�����-�2	����Ba�\u�����}P���cJ�Ec~�3��D� zt2n!�ՠ_��e��[l�~���d}�f��y|�1v�vvxgG���}�q�i���M_���ޤ����|���5
Y</��LJ-;߮��f��G�-Nq".��],�UJ��������n�Su�=k��t$���݊�fmD ��v�*5��_9|񜧕��YW�J��%�r��[u��[{���6�g+a���T�,�7�e�:�,B�h��ԃ��-�Y�s�?R����;G�)����{>~wrm�E�����y�}i�~m6V}S.���s�EϠ��v=8�JӢ�o�~�oS�5yp���w�3_��&��>�=KlNӢ��J�-k8��l�zg�%pɆ��Z�O�踤��ަ=y�x<2<�ݑz�4,*m���[cӷ��Ux')t�����6~�[����]�j��Z��d��qm0�p��
�!���R�	u��h�OR�#ޭecUc���C*�E�K��Y��Dl7KEDY��oK>T�%5w�=7���\�+ωq���=��R��ﮣ|�!��!{mG$�}s�Pۙx{�Xê�
�c_r���]�7��ɖ}N}������x�����e��y�W�{�\F��<=���[�srkbU���;qOx���g��<T�SND��ޫ w���{h��NC����w�����t�_I7}Yyh�b~�>�����9�.Ah�u*��뺔o�J�M�/z�8g�C�����eeX�N�|+ʏ^�]uU���g<��{����|2K4�U|e� �HuG���]W\t�J~��A\z	�>M�O�L{�Ƃ�Y̲w���]WjӥT{ܫ�b�V�:o��(Z�C���W4�'b�!���`e{��z��`f�}���s(u����j̫hST{C"ٯ9���=�� �����Z�Sdu��ܜO[B���;Z��]cm�些+{�4�l�8{޿\{>'ƙ9T� 7<ND�VE�y�j�[�{��z5�G{�q7���;^G�#ޤ8�o�F�z����2\� ��H4 6E���F��Om��ލ�ļ���f���ϐ��o���������z�~�����f��,��r�Ey/T�>�n�ev�>�}$��ޤ*��tnq��p�
��m_��C���<o��C5�z���o �޹Vqer��:H�u�˛�3	\X*}=�B�Ը�%O���#�ʪLt&�f���������N(;��h���Ǿr��4�'�d���O��DK[z2�׸�oSp��'tV@��������+����So��'�{4X��ԃ]>%T@ɇ�wL.��n��/������'#����{���>���[y~�U�9���~*~��>���>�m���c�aݨ~�[Cl��]�͔4�Ϯq.��d{��L��ӟ>��N�K����ׇyϝMc���g�f~��RL\w�����{Y�o��D��*�٩h�rˁ_-��D��NC���~u�z����{�"���H���n���s����uݓ�itDi��Y�.Wd�T!d�{�h�ƥ��r:m�� �I����6��=r�i�^��ƙ��V1MR��j�%���f�������A�ɹh�s�9mԝ���K��s	����:���k6��tK��j8r%�n�\Ժ:.���;,c]�9^>�z�����Ų4��j}���.�
���1�&x�Yd���$�#��2�頮:`�9��$NU�M{��� K���u���C݅�#�Գvx������4������W�+Z����ƙg��[���5z�g�O����D{���q.�K(i'���ʡء�#�����{�}۪��uO����%��.����O��F����*#o�z��� �.�r �7(�����yW�}�����y��e lx��A���uG�>��'<{Kd��D{}r6���3弣�+=��U�=mk�l���� ��p7�/�@�q�����ٌ�N��w�L���B
�30G�{��s�|o?A���#�!�L��ch�9�g����[�F�J�a��~�3*EC�s#�u��y�*�蕞,��"W��C=<�:⼎ςUߠ[f����ʸ�餥�y�%�����J�2���ȸ~u�}���7���Q�r)d�!�>ʊ�}[��[.c*mr�gmT*�Uk�F	������Ⴘ�5�IY��S��H�B,�C,��7c�9�O2�� ?.P��R�U��>���=�e���nĻ:�Zh�Y�B�]aB���=���G1]�6�U������Ѡ��9��)�R;������X�±_G(΃�ҭ�Bҹ�1�~urn!�U���>`���eH(��߁����F���~�~ћ�N{B�m=7�+�GyK�qח!�]�����n=�^����}�9��V۬V�n����9ć�,�����������*|O��\g[��K���ϛ�Wx��T�ｓv�J=�il�jڬ_��g�6���Ggne�P����*�����w�z�9Q�J��j���]G�Y���L������i��Vk�W�7T3:�Ny�Qb9;�FK݇;[�����Dy_���J�`� G���z�2�J������mO�>% a��=P�T��S���3��;�#�k{C|q�!����s��Sy�<}/-���G�<w�+�5��O[�c�Sw�'5{�z/�F_�Ǯ\	f�|����W��o�x�s����[�ϝe��Q/��M��9�{��k{�W�t��=�I-χ|��Y����7�N��>��������p�c��T�d��{�Y���=����>�
P4
G�z����z��O��}�h�b/�{E���{�<��=�7k����|���R���J��:p���\�&aVsK�U���S�ע��볬ծv��tm0�l����f�091�oa{5������.��]���H���L�]f+���)�]3���+���F��;XŚ󦲹V�������a�@�,�( r�2�7�F��3�FXW�ւn���]B��c�*�����u���.&k樓'�G��8G�;?s,���'�_lw�c��w"ӿG��.������#�ǟ����D����d��ޭ�~�����l����1�݆��#�?`B�x:�o.����G+Ϯ71Q֚�I��R�=^ o��԰T)d�X1S`df?�a����}��+���w�l�����P���=��h��ޠ;�^��QEPۣ����i]_�~�}1��A�c����V�o�²>ާŪ���'�1�k�W���/{̟;��������-P%���x�L�>%FkFևu>Ӣ⓮'�#z��uU�V�S�C/t�g��\%Z���T;���z�9{UbU���Xus6sK'v��/T	�0�'�d��s2.�W�h��mI�{� �%~���9	ֲ����r;�zޜ�+�� �^CG����-YC�)�w���W�:�y3�^%��k�
Zݑq+Խ�>���J~t���5��s�U���������Pe�����ѺeŦ��뭦�M���(�ak����}	�]���K��ah�x�����n�tk��=�t�.x��q�A���gX�������.�0O��HsVm+4cz��xٸK�z8���Ӥͣ�-�-s��Ff�hN��Q�ם%A�������n�����^��6�,�AcWO����TO3+z���)?L�>���[�n�X��vc�Jѻa��Ej���!]�n@u�@�^��g��,K|�9�O}I3m�]��,��]2C�Źyy��>��Y<�"�aO8���+6*���G�iss3�g9h�b�gV�d:);�h������-yNvQ��#�ַ�TV%F��+{~���:����:�Vm�2nV=<~g�����R��(n�ǌ���U���vf���֋�o*j%��oD�\�n+�eh��^��t5�#�j<&����=��묫A���m��6� Z+t�;6�Cu}X�����I�#��;l��F�G���-h�˶7���-P��w]�e�� :P��Sc�n �y�۳q��m=�P˫����I��Bвi'.��9ϔ�Y}��\�֒2�ŵsT�˔�]]m�����GR���/��7@G�5�.���l\���T�2�s�����m��QZ�*F�j�'jf��Z�q�b��Ы3��d++� S=�E���J���-/%cL�u�ɮ�`.�T� A��������@�Q��z8��x�]�-����|�<�օ��%`.S�㤨nm��,\��{��ݷ@��f��06��R��sV�
�f��)��ǋz�6g`ب��r�90e;��ف��U��S�д �	܈������F�w�G
�i�ԫP�M֙�u��l�L���n��S��[q���v��z��D<A}جp�ٽ��b�j��N�.����.��Z,�x�}�ݮ�v<�zC[��b�ޞ�\u'����Ћ�/aKE.�LU��������GQ�0�1�;z�7K8"�ZT�t��t�'�w0V�Y8�(^(����͛��Ss�$,�~��
�@�*�v�w��L
�SX�x-�{����|�-�+[t׈T�W%�+Gf2E8��3��֒�<v.�V��wK:h�h��9��c%���j+�[ݓVX���T���k8�ٵPf&K�9�]��)^����V�'2��4�m�]�h�ܳBx`235Ԏ��c��N4��U����=Z/;���2pb��8�9����>ʍ��~������ת�O^�B����N�gc�N�o]�l�FIY�G4��]&�uM�^:�;�ï�T�K��W��ؖ�g9�}1��y�9�}zK�G���a�)5�ڲ�5�{�`�t�b�#�y�9.Z��:����YO��]��)e�A�o0���ŗ;x\Bew�����%L�[gL�C�v���u^�\�9��>��s��DAʯJ�+�NR��\`j��a�JR��YETAL�����"�T��

;��]��#���*)D)�s�r��s�uq�q�i��G;�q�r!�TDUG��U*��E@r��r�9%d'K��(���s#�Qv��$�)
�%�"�Ȝ�TPE
���ND���NW8AY�%�h���.h�"(����G*(� ���Fr��y�n��㎞0�Ȝ�E�����AU`S�aD\�Tʉ���v�*EDPy0Bs��"G�G(r*����N�Ur^<��DQp�(��it"��Ge)Ȳ���� �#��'�"�B
�x�9\��QVUN��E��v� r$Q9�F��r��^ZA�*2Y&Dp�*�\������+��DEA(��).�U�G��8Ut9I��\��|���W.���Ö<B�Xd�Sz;����,���7��ɬG�Ʋ�o;�v�年�lf���;Y"��[k��\�w2n�Vv��.���˨��^�F�T3�z}��}^'̯k�\?�G�\wg�{�)����zFogxq���\��rI�,<�L�wS>Sn��}���xl�a_?K�T<��iaS��EOkܼ�᷾}|f��Xg���H<��,IR�UL��*�+ޯ7�Me�x���������E��~w���c� d�X�J؃,	"EA���>Yu�q:UM���S��Փ�ޱ#λף"���߻�4���HN��z�q��\�@Á��́����e�����)�]:}h���Bf�5�\Mǫ�g'����&���q�&��sP��ޅ������!7�]Q�<�w��J�@�)���4_!1���9��w��|vp����x׌�Y]�3'��ԝ�q�'�K�{�'�Rٲ䉉n���|tnG^6�
�mW��~�"|p�s���j�J�O�zR���>�=7���ʞ�L{�`��=�B�=K��/J��Dzߕܘ���m+��p����Ω�f�U��XT�&.4�2O�OT�}p'�`���~�u�7��Ʊ�o���r�[Gh}{��:��V[��~�v�K`Ȁ�jf���Kr�"�r�
���l�ow��e"n�HX�k��<��O����7��9�avv���lB$��f�e;�k>a�oV/�z�ԏo�_ħ�Gd+Je�v��)��%�J}�p��D�UT�{}C�7�?O�����b��RF���j����5ҟ�Z^�qo�\]]�ѝۥg����g^_�G�W���~ڱ:[ɡ�yR2���N���L�yNhv�<���>�]��o:��?V׼n�V��O�n3�߆D��i9	ׇy���D�����n�$�:�n��X����Ip(���Q�����TE����I)s<6��-�D����v#�;���p�ӽ^v#��7��H��:e�粏����zN���c(L�W�O�躗C�r�X�~�W���מ˾>���5��3���l�Z���;�b�յ<nωJ��@�."�|����4�|l��\�,��a���]c=`�C��z���J����kjY�<I�0�j�b�R-�&��,�ٸ:��@��O�_�X����X{���ȏu�~�=�K�AŒγĕPf�+��|�@ssU��|��_���+!��K7�7�n��NG��9��P�q�TF��^�D��r�z���L��>�J=�$f��~ fO�N�0��`�U���4r)�\M��is;�����*����k�ҟ�s�zF�7]m/��W�e���b�(҆V�S�a����=r{힚`��7y�K�<=�E�f��4z����ׂ=��鉷G4��;�1���P�-V'Z.v���&Vvˬ�6�=Dʈ�i��!B�q"i�������=x}�C�(��0��X�unsV����H4��>������ih�R�'^��dzw����BIل��:��x:���Y���˺�����E9��*���2J��x�#>�+#�T�޺�j�h*���x�����쳇Ӟ%�x�dNa]q^G`J���-�N���f}q{�2޿��×��ۛ�����/C�d!q��E�ɺ�>����*,~ːj�z����\�������Ֆ��Z�˨������^F���p׶�2�\�{��o��8��#�s �S�{'U�p�zP����sa3�N�;�v���;�񿳯.7�9�@zMǶ�»�۠��1=���-�_x<��~��|h䠣N�Օ�J��7���g[��}.k�a�D�i���A�����U��1�V'�9��{�q���8P���|?/�·u9GE�J���B�`T^��x
��TتΘ��MzuĭT����ֲ����Gz���ʝ6�'v��<��X��ɭ2\��
�B���2t�˚�o�8����+@����.�3�ƾa�R��ۅ��O�vD�DxYО�ҿ_���-.����x�á�y���3��"�����ۅ��_r�k�]W�dJ4��bS�'�ϱ��	�/[^
�&!�G)�"!�I`��{��iޮ��q�{a˱:KmN��彙�X���wVy�(����q+$�Q�=c�i��nMP����՝s�f��<{;�Z�:�~VG��x:�x<����o�{��~�<�=v���yh[[R:�x�ƾ�g��~����d�{y_��A����F|��uʁ>/�T8�O��7�<}���~S��u��n�P~�������[�޲y���& yTz�e��ϡeԳqMՉ�i߸�G���#�'Ǯ�O��=V��g��>��X��`�� jFX�G�Gz���{Ԅ�z�hh眰
�����5��m�b�ۇx�<��Nz+�l�υ�f�A� z}$t��1a{�!�P�z��^@���{�,z?[��c�#ޥ��Pt���Q�f��<LLD�WQF��u.�E-����=�Wz#ơz�|��	���R'�=:6���/�_�&���e_��l��}�T�ۗX�1���w��D�ңqu����x�4�GZj�&��ԁ�|=^ o��k ��t���3^�T<���X�,�$��3��8t�˯x������{�ܛ��F���{��_���Z����^ט�|��ɯ�1⦎O�\N_�+N��}~����WP���Lx�<Q��.-��b��Z`fl<��v�syioz��$0@�Y�;���bOr�T�"��Y��4�fWv�`3Oe�0ҿ��ӹE��ՠ� ����(�:X��1�n�E��=�-�uvu^-�M��b�.�a�&���;�55S&�4���t�Wht���`aHm�	w����<꼇�� ����d�W����*}�E��q=�,y4�ȼt}<���[c}�G��*}���P�K����AU��q���/o�wL9����ѳ�r�Ր�:��/h9�u�^�~�נ�'Z��j�w�{HV��g�l��!����2���<��~^��F��ڤn�y��m0B�싉^��I�]F�NC�/m�z�d����Mlg�G^^5�����%���z�_��n+���8z}��W����x��u�?�֮;���+8d߫V(��t�$rK����c����*g�b��	sp��a��W���G���,��6*�*ѷ�f���;;_���q��sX����,���A�,E���H\G]ԣ)M	~���3�Ċ&��d��+�o�1䃦7>�Q��~w��<c���,�<I@�,�ŵ:���fz�G��(<�X���yg��T�z<�|�8�Pү�HN������r|k�DTf
����Roo@��_L�g��}���G���:��%G��ȇ;^G��z��o�o�G_����̗9J�����T�#��=B�J��/��8��g�s`Ε��aIT��0��↊Y2ڭ��ٻ�A�G�
��T��F��<��ܾ��cwư���ɺ���%�c�f�)��Jh��La8s���ZBz�)���yق�S3��� �B��]&���������X/%:`������h��*9�Se������h7޾�vG�b�ߣ$=��R��X/� ׎��O��9��^�S�{�|�G6��W���O������f83��2o�k ��߉�}=6faz¬��Y�\o!*|m�Q�y9��ޣq'��ٕ���*�Lzs�Fߧ�;��54{� �i���ݓ�_P�˶�ޢ����v��(�ʇ���"{U�`~�m�	��E��P�K���٢������*0��9���W�����Z�~Y�#�q����b9[/�μ��#Ϋ�r5����{j����\u�H��D�/j�~�1]k8��o���df�o�+��L�IӋ���g[��}���ׇy�ǝ�J���Zꇽ���$��m�}(�)�+�%�G�V�KVUi�W�F�K�P����.ix������\�l�s���;D˅~�j����y3��^��ne��3�]O�踩t<�i`%]�u�wo�}��r��k��^ed;W�Ռ��V��>%+2�W��$�#�n�-��hϜ�����[�����@��p;ą'�"2�@3b�aHDe]���|�?o�D걞�5`{Ҳ�ŕ)Yܳ�á��9Rg4h��v(	�>)���5�)�X��:A$
ʕ���]r�j��{M]N���mV�_Z4&�܀m�)��JX9f{Gzux�9c{��v��ƿ�GEh���\O��2M�-�=���\��f�]G���t�:~����FG�O�܏u�~�=�"^R,�X�J�ٖ�j���w������Y0�FW��Yw�S}q6�ߴ�y����P�y�Do�U���:����/iw�WzI�}@���{��l�[4*����}I���cޓ�^EǅFu941Vo�˺�+�<�Q���s����l2N�ܰ�H�F�Z��Sf2��>���w^�W-����~h��S=��/z���|d2K)T�ݎ�&J�N{�r�9�7^mL�s>��ӝ)^s"�m0����ώNx���Q�*���F\����/@�R�M��-�ZrƊ���+�j�9M{ʼ=~N��~UR;��x�d@���C7D?e�5�OW��|fn�3�P��~�`�K_~	~��9�k��
p�����1��ɿ����_���8��#�s ��~����g�5��4.{��K�(/��\5���g?A���vz4�zW���~�=&���xWr���$P�&M�nH[=� ���5��Ϣ|ȨlV+���C�-ز(�7�-xR�UҒ{]]g�Whvj�����q6����æl�Y��so�C��@vû���ᥭ�[ewZ���Y��yh�w��N�5���U����}BA.���8܈b�w���9~�
5'�F�����ۊT��9�/��:�ǲ%�{L?w	đ�詙�U��^RUUL��Q=�޽��L͔<rp�ވ:�NQ�qR��;����p\�	��sˤi�Kgoa�]c;р�hs������Gz���ʝ6�'tw�|�Y5��O*�iY~��([�����@����lJ�lR����9����jxݟ���xg�����^�{"�+7���w�j�mߨ�G�C}�"�J����Ǘ��1�]p�C[R9iF�yż�7]
{�*����p��>f�3�_�e#�}Y����{No�x�s��\?)Ͻn�:�P|�C��[�ok������l��s���2��T9%��腗R̷4'~�����>/I�G0�d����u7�{��y��au�>�`����&������ȯz���v�]����Nz�dw���BK��w�):U���\N�z�qD����ʌ��[�"�%yNE;�+h��]v�����������C"y��޶;}�\M�{��ǫ��,�"t'���"Y5"s��6���6*�9K3� v��s�V�ԁr��&6�E�11�d��%��-�D�p�Ԁ�*��,h+g��m
��kzf`�e��/}ܯ
וb�Cuۜ]�`\H�E�p5S.���w�:m�4��ݹj���*8����3���٫]�ޑ�X���Ը��G�Q�{r��|��	�R���D� zt2n�Zǯ���ʵܟ	F�5ys}謧��"Q��&w�Ѹ��[���b��U�+��R�=^ o�!��Y�s�DRWS������X�6O�t�,W�e��>��W�]/��zT5��CU^7��~&��|��r���d=�v�=�T1��'aL2��9,u�N]Jӣi�xR��|m�ˇ��H�����|vj���7�V9�1�߶}z���7}��p�6<����[�z�[�F�`g��w�-����Ev+/�-����^����{UbU�E�W3g4������gՙS�{}:�ٵ���Q�d�s�>� *���ȗ^�>N����X�9�i���p�����^W�]�pԤ����s3[�F��7�\VUi���%Fπ[�
��zK��o���B���!u�J��GG���y&��G?}-�\P��U\n�T.4�
�c�M�R����Be\�{�"�g�_�V�|�r�C�ї�W���S�x]��x�	��g�b��	r��A��|X�Ȝ��zv3[o	�dD'k���8�fYv�Z�N��t�,�d�ql{��`	�ڱ���?gW�-L5k�4�C)�-7�+J���o�ŝ�mcCvO���V�f.G)��	;��#/��bKx��b:��<]�vb����"Ysg`�����l��x����=�]b6��,�_I��A�,_�*��뺔Lc{�{~��'��dg{%-��	���_��!�c}�|uC��dY���Yc�+`�`��4b�u�8z�o^߫�}+��˨�/��GC��ё���WzF^�Bt�{��`�>,�{,���Z����rAYH�=�	������o��c��#��!��}27��LM�C��`��]fe�U���F��x��*H��θ��؄�E|�
��o���������z�z�ut�.'��yW��~�G7���ٽ2�%�S��Č�_�
��|tnq��q���m_������:���R�tux�Z_N��x`��I��}��񡱗�\k!*|CK���ށ0�۸iRWi���{�ܘ~~�E{���&.61}BӃ!��7cH�˶��[�0�f]M����^��5�F��Lu�w����w"����m�|��f��{jA��V�2a�硋sr(���vŸ���O��~�����K���+��yח��U�9��<f���`��M���i����{�QVW�,�����-��QW;*fZ&%;*�,�x�~��y��h����ǒ��#1;�R�W|��h�퐿��o�jƉ�srIՌ���·��C�w�s�k�c �IsB�.�κ�q*��,�h[�)*��e��:����l�I$�7�h�jq=Ys��w���M��.�̥ƥms��\�\r���8sF�+5�u��w�V��,��fgs�a�F�n���{ԫ5f����ivф<yh�۱�g\�ǡL�����КۑT��_Q��oW-����βs��]ʻW�¦��
M�[7�9���2�|]*8*���z��w��8�%�s����ZD�xwH������7���J}����k{��Ż��h�}ٚ��E����/"��~�����}iWN�X�����7٦���7�Q��0�u�V��Q�:�}��+��kzs~I�lz%ɶ����>��8/w6.�Ru
Q�x-�T{$5���[�ތ��i������\�ef�F�leg7�4��$�x1W^��x�&�iC���tY@��=�J��9tcRǯ��O^g���齎�_f\�wh
jΝ-�ڭ�~Y���ᵻ�����/�,׽�8H�ӯ�`%� @��qnƉ׫��r�ÆH�Y"*A�ҙ�%��ge)�+��姹S��L��Pb�褺�'{|-����U+� *�u��a�.�0�^Ժ����t�05�`Dk
���-Wi�g]�R ۀ�ܭ��E�7G�&�.�>�X^j�z��_6)-�k�.e��t]�)���i�(�`+W��+�L}t�H��A�^+���[��V
��
ŸB��G�j<1;�E��s�,'��.��e��ǧ�Es�q��N��)�ӷR�(�C��.�a �.Z\�V;C܀@�i,[s�R=�ʶZ�Y���8`�L���*���+EH饙�]�_ ��BNr9|v�7W�:�D��@�_V�Wk:B
��z\kg	�i����=w�c��5M<(%n�;����su�b+�r� �����+;�<=�]5�)�+F��+%���3b�'H]@j�ɘ¡�8{�����av�0�M�6a��.�(�<ʕ<h?�|�*�a�[v�?u~�=|�0˗Ne�.T�v1Z��l�N��g,w.wa�ާ���/��&�8�:�|�Q�Ne'�m�9Z�2��9s����ib�7[��Cy.<V�DXx^�Ā��u���C��4���)���#˺ܾ� �	��F���aoL\��Y�0S� I�i^����qPޖ[j��tý�m�W?u��R[��.��̫�O*�,��tƝ�@�����L��]�x�ŽQ�Ρx��y�6tK�Gm��p��<��Րi@Ic����y 3u����\�]C��bd��".�v1Lc�lYAf��}�����"�3� �ۀ��r�+����+�D�^���$�P�Z���V���*#�**��TQʎ_����Q���*#�DT\�QS�*��R��vPs�Dr�E"��("�(�(rq!W"�g�+��J�RBȨ��*(�PUȠ���Er"5�jeːAgH��"�Q"	��&�kH#8����H��'9"�QE��D0�YYbWB(�jUA.!&�B"�J�£2�f�ZU�D2ƕPmm���JT�*3�9���f�gJ�D�TrT�E��s��f�q�q�����U�("C�T���Z�l���J�(R%E�E�vA«#͒J�Qe�ȓ� �s""��dES���eI�%�PQEG
��DU�"
�I�YW#�P�F"dVID��(��<��ܭD�fE�L*+�$A�(8QE��T*��QQ�H��r9k""U�I�$��=ĵ3����o>�mnbv��{(�&mK��ճt�l�"w����8($:�S:Ճ�A̪2��Ό���Is�������)ć�/��x�Aݨ��h��T��t�.��N����n�;�|�by�p7�M
}����U+w/�=�q�9E_��x�oʒ��[�iE�g��+�dK�^>'~��t'��-���]}�Yb��]�&{�;�I�"��L�^'l�Bg���Q�u.���,�"���U9rz���K�g��H�}�~+�����a}�jx�E����2��,I>G�L1��=�M*���yma��4��Lp�:csާ�=t��>.�>�\L�C	��g�:j�n��|Gڪ��N���c�2�o�t�<���8�z�{A�9��Q����q�yH<��Y�J��1u��}��p���Tz�(�ed,��񿩾��t��|���HM��3�gH�U'}yNk���7ƫ���w��ڇ ���|����-��h4U?+���z�9g|W��3�]Q��ΦsՓ���o�;���#o��[3ndT�l�<�p6�C-}<9�tz
�����s勈�n�N�L�{I~�A�L��qd�P�Hn�QW�кs�;^o����8��yl�N�ʞ�ҧ!���/.�Z˸�zPڏ�<�N�s	)��T�ك�&�a5�\�g�Q䡜�x]����xwe(�m�D�٢�)
U�[s���e�9��J�ǩ�4��v�FbUe�H� �����麳�n��Py77�xjy��V��6r�Wt�hk:��/+�c������y�Q�*��@�=���l��r�W+Gnފ<�j]%�}��ϼ���N��~Wr-7^'��O��c7�ԃ�)d�P�8w�ii5�(�(����G�w*
S�w��l��T=)�m�c�=�긇��}���Ŵޕ1NQ���%���(7�9O�Ij�����\���/6_��ˆߪ��~�='��^�=�P@f�t���+�Wz�~>ٜ���(���V6t;���6��O��_��:�Ƿ�2���&�f��؟<�����c�{ފ��Wq*�������l�<rp��᳡�NQ�u*���W�%��yfr#������ҽ~�z��c�X�ϻר���N�E��fa�}|��<gj=.��u�N�3%�	z׀���"�W;`���:������jx��)W��G<Q0=�mz�޵މd�~�U#Ԥ5�����Y�W�=^�<�U���D��;�8�.����6��|�W�g�Y'ƢKd0���Y���}�^ӑ��������� {�����0��MT���ۺ��Ɋ'r'�!fI	6��!T��5��f�{����owR}��+���dmF��`̇H��yL7����ėM��x����v����5�%G�8 ��.L�� ��"H�un�gn�k	^��*�ה:f�ԶTmpC�>��<	<K�yT;��n|2]K2�Н������ɟW�[ۦ1dwN��H�ö}����W�����,v9Q�"��R</����ًa+�f�%m_a��K7�bT�1����h�yIҮ=�����]�>%��Td@o��Y�/Ǣ��U{t��k=��S��������Θq�޶;}�\M�g�px߫�L�f��E�c�9���أ}�皏"c�Oe*7E2�!��+#GD'�lgޟR'��:/ޝ����c}��˓3�xa^�/z5��d̿|���rDĮ�FC㕽���b�����M�z�>χ����*�<��9)G�F�>�=��`5Q<(̦l��/�Ele���9��7{n=���M������ݓ��pO��|�>��@rϼj�q�L�S���KcӃ�V����+7��OܳQ���׽��� �~�ꟾ�8�)|�~�����>�=~����3���\2a��mhw>ӡ1��ڱ_c�*�3|lO=&����s�Q��;�����z�P;�TM�s�6���%ݳ��fdKWԙ*>���鵅��r܌Q}���ٗ8u1s��:rs�c{3�*Ka&��y8۰&��֜�'˔��X���8v�k�������c[/se3 [I��D��L}Н^)�y��.�����gS��ooRq���5�YM���}[^�Aͅ��{�~ϫ��YY�{�܂yg_U2�-v�֏X��H���e$=ĥ�0�����Ν����Yi�)kvEįR��ﮣ|�!����S�u�Vw7=T�2�';'�|J�/�u�n+���9��o�����sW���b��/*n�u+������=�&r�tJ��:����KG�K�*�l���}��W�cb�%��ސ�}�Fz��ǰ�ޗ���=��#2��7�A�X�>E���Hx�r:�h�x�l{��>�}�V'���B�!�c}�|u�T=�q_�3�8�q�l��-f�:6H�x�'�U�jv���${��N<��w�7�$[��ё���V��iW�'M���`�>>�o�w�>���·���A��zY9�-���4o�~W~�,C�y߽�C���o�G^#�w>����/}�C(����OK �K�s��@/���h�>B����s�;��:����m���_�������;�B���ߌә%�U-���D�/ԅ]K�s�2�n!Qν�͸�vF��F��RQp)�BY��3h��ȡ�>�y`�5�#��m�
�Ѱ��d�2n�[�R��cЬ.3o7Xrim������j|Ф��{x��Wc�Ĩ�湜Qe�s��>kx�e|!���w��qtc3�h��n2�u���bё�jQ�˸[�0~���)��|WN�ܧ��W,N�ЫK���Zkq�K̕��� 3+�Φ\ZJǹ>tB��w&~�EG�>��bb�z}�I�Y=C&X�a�V���g�'�`��������h�W����z�:�j�	��E���=Sp�>z�{4X���R��z�\�^7�+'��?@��S��(�>��Å�u��g�u^��C�o�V'M��c"kqp���з�a��zC���	�0�������t�.��N���i8�xw��~��:����}�畃��.�b�s�r�|����<t<�����L����[�q���ʕ�GnO���w)EgyX�.:O�β���r�^�F�M�΅�p�̱�����.�����0yŲ&��5��o�S@/|1_���^>>�S�Y���|�3Ʀv5����i^�Z|,����~Z�<��u���_�2�t�Q�X#�ht��C�?��C��F-��f�� Q5'��y�$�X�?ߏ��=x��#��
�7t!��^��	�;��=��Ǵ��� ΁ak��d]P��mH ʜױ��a\��g�,�PI�2H�e�m����@^бX�oi�0;�`*�xx�XI�t���� j���/c���M1�m󱐖j���"�FmS;L]naS.��ZeqRY˨I[����)�ո�P�Oj������+IK��wKN`#9��R7�9��鿃��D�:�j��El�Yw�t�\K�^��y��Ϸ���~���{����ŗ�Y��]v��l�2 �;X����-�kj�G)�\M��i��싹Cۄ������~(4?N�����y�7��Ae@V�2�7\��P�FZ%B�:1-+�lS���If��_�;�1���|[|�XO}����G�~�@����!yM���R�5�ǑK�-G:1�;�cϕ���c"�����}9�^x�d
�n�irz�0��V���D�Wlґ+{�(��!�=7����sϦ��8�vG���p����z|���)�.A�N|uxE�����ޮ��E��I~F��\�Oun���x��o\>-{+�C�o}@z��~���1��Zw�|��$Ν[^cОT�^�'����
�պon_#���Ϋ�}��;�Ǐyc��;�b���e��s9� ����
�=���g/���0�-:��fҧ���/�U@�=$P&�����Ƨ�饦1��]����yG�׼n<m��p����L�~����T�x�?���j?'�w7�޳J�+��^>�)+�k�5fގ�l� ����MᎳ�z��U���=��̳_P�W5m�1�%aMVm��"-�k׬.�4%[�۵YC�NǘF�Y�����B�d�ĵΦ��1S���P��[�1�[mL��l�j3s��=���P��o#�>�K��gӞ<�~����k�[���zk��qg�t^���s;�^�:=�H�EK�������"�s�;���wHw~�CVL�g=�,�A��5���:�ϸ���1�5UGK�Gc������}�!>��Ol_��?U!���9>G�`�s]��΂�.����H���G���l7'>��W3�'��[�ϟW����VN��H��ټ�7�m^����n�9��d��s��İ/��P�*e���Yu,�sBj*�Mݘ�4�ԝ����BRY|s�'ǯ<�M��D����`�`)@����j��颽�0��U��
Z��g�^U�.}H`�o�m�):U�}q;u�a�,�������O	�z��JU�V}��!��^��(��A�y��޶;}�\M�px߫��,��:�����\u�]�v-{� ��8L�ё�>��7o��?:aǧԉ����~��$h�=4k�I�U�Z��9����ı.�q>�&!��#�'�/���w\/i��MW��~� },����V����E''�U�Y=��^Jo2a�wg,��;KՕ������S5�W�C�)y��Rg�P0(����"��^�`��r���H�9]p�T=�b��[��DI[��Mz�e�XYܮn�J2H{QtvU���׀r�H�ʀZ_��VE�D��KG�ߡ�*ׁ�S�xT��8�ȗբ��^=G!)|m�mǱ��T��ޟ�I��vg6�y%A{���dѿ��@w����2R�eMA�c��Ƕ*V�O��fq�P��DVn���b��G���}�~����^�~��	���l��}�p��|J��X����b������%���f�����^��=�ԇ�:��G�{�3_�w��yU�W���X�yS�C'3����ߵ靈��s�O�}x��uo�;��a��`
���^�"�ecUc���C��Q�2]����VoS���9����J��VUi��e���� ���d\J�/zN���){+c��sٟ�%ڣ�*!���?�Vr�vE����V��O�|c�p<�A��c}^%*^���rK���6��)nrXa��yq���qݑ{�j8����:�����z4�r�~Ayz��'ׅI���`�f��/|5W��������|��k�����^:+In6��`9��s�E���MP�xS����iu�G��Q��+ޯ���7"=�|z���{���E���<I\�������遴�A/ao�֓t��A^K��(^[(M����D3������'�3�V���8Ҍּ����YVc��ؾH�Ncx�����ݢ�:�S�����00������7E��9R��j������\�����gLj'�y����g!���$Qr��]LO�"��/�Oף#ϫ̭��*���鸏z�q�=�z�ٴ;�XT^_\�׹֮>6}���@�>u���Vb5��q>�+AC��#~��pYH�i����.9��g6�1��Bk�s%� 9�>�'�n����!0�P�
���m�q�S�	�sݞ����݊�mP��h���}޾Ƽga̒�H��B�*_��W�����o6��҆�8y�����~�o���c�_��E;ǹO�l�X�~�:�.{ƀ�d��j=`d��;|�y��+ڍz<��Dz��ܘM��x�И��O��4�'�L>DQ�Ą��ތ��n���+�;���l����1�'���=Sp�>z�^�.;�R
�q�Х��}Uz�KQ�%Ƙ��;�:\���>��r�ח��3�*#_�x�Ƕ�N�r=��s�>��3�ۦǕ�H��/�]�t�*>�a.������:<�꽤�\K��<�[yY5�\ھ�wL2�k�yn�H���\��#�o�訌&߃G��齵�C,jc��X�פ��/8/�(�[�jE�:��1�-AR��1��l�AT��3I���<Y՜�=�����ʅ7F���Bo��nVR���F�����ӱ��u� ��ch;���]��3y$k��s���;��u�
0�	wcT�sjV��*�[�*[c;чL���+Ӿ)��o%��n4�L��:v�X�<�S�:���G��Q���-��Ϣ����� ���>r�|��O�:U�׬Ƭ���Y�)Y�2�$��p��߱��m���DT����/Mc0E�����~+�({���涥���'�3����K��S�$�3F�3��e#�S�O����<�w�z=����H}����3ӭ�5z<͵�5�+��'L7��o��l7K@��rzY|.�X�ߴ真9��%�MEA��7I]M��<�箈�^���d�����I`Cs�pʸ[V2��'ў\'||7�xmK�C��{ۇ�3��;��+�ꑓ�eÙ��qU �u��~(\�44N�]�V��>�]c�Ϣ3�^>u�l�zw�����%��{�^2)̖j!T�ݎ�l��Rꊙ�F��g&�����r!�a�ϕ����c ��ώA��y5Ә�Q��Wz}7������͡s�}��s�]F�.Z�J��TC�Qz���^W�9��~���� co���01��� 1��`cm�� �6��`cm�� co�01���1����m���m�co��1�����01���m�� ���p�m�� ����m�� �����m���m��b��L��t�Mll�� � ���fO� ĒwǼPGmT� JR$IHEH�EJ�H"��V��RJ� �PkQQP�%J���VJJT�[`3c}DBu�U*�!"mf�XU�)Zi����u���Eq����km�[P�UY[`��bk5k���Y�N2XT�zjv�K0*��B��ԕ�I��[j��ڶ�f�km�lƚ�a[m���3Q�[*��5m��V�5I�ka�[&la���-��s6����� �aIeZ6֬�M�����k&�  �D�mܪ[^��Z�G��c�s�\]3�u���To;�׭PڳW�/x�j�ڕ�y�;��p�j��6�����m��n��RRzz��EXZ�cmQ�3j�1m��  f�U���5Z�D�R�;�a�{�t}���PE=h�X�EѣGF����    =���   �c�( ����h��8�h����4Q�ϔ����eV�֖���J�  �ào}��岗h�Twv_^-�{ݎ����W�+��3ډ�2���X��mU�חz�֎��ݫ6��W`n����^V�J�ifl뫳%@Z�    l��ͬ��wz�wtZVwg24mh�=��P�t�������9�î:�6Z{o^�ͳ�S��gU��`��v����ڠ�筽{SMӹ��z#j�SaM��n��GQ|    ��m���ͽ��:�Ws�p��喋���{+���s���a�m����SE;�Վ���鋳�����ז�iMv�ׇ=Q�v�wOU�5,��n�%U�4��:�dQ��L��g�   ���W�N�����kCfvv��{�R]+q����j�;s�n��Mnݞ�޺�WY�sޏ5��.�:�F�wz�\��+�y�/^ݭ[4��׭ռ��:����#&m�k��2
2���  �{嶧�imw.��R�$�cV���Q��V���ty(:M�����L(mWu^nڕ)9w����Uv�-����r�W��v5T��n��v�v�v�ǵ�ͯv�V֩l�[3#V�|   ����tSZ��06�Zԋ�����wt�o;Ç�lR�;���y�����hs^����h�vb�m�Wyٝe��'�4v������9����@��n�vU�z�ڡ��E�,��  ;C�o�EM�!�۹M��;���»�ղ�R�{�������U�x��N�]��c�v��ݪ�Թs�j�*�'w��lP�yp݀���T��E7���g{L�f�f�Vedim���J�  w�'/[�v�գ�6��.�'SaZ� ��u�뮕�؛w]��n����ۮJ���O{۸4�
�M���6��3�y������`���J�*�����fU)P  "�ф��! B)�a'��C&� )� ��z�  ���U*   i*z��C F������������w?����F��;)���
�Z�ߵu���5���$����$�I���BH@�����$��$�	"I��������+k��4�O���~��m!)ѱ��uk6⣸A7�ʳHefU1��m�Ci��6"s))���u��@ZKH�@J�؉{.��*���W�@�3X�+"�b*����+(m$��A�u�˚������Lea�k���`�d�k�E��i�bf�����LĜ.�Z�S:ZȬ��׶�m�C2n�x�J�4&)B�˶ڴ+j<��q[�f�Ԧ!�SN훭��V�o�%fK×n��u�f]0�CktSt!�ڛG�N����	�ȱ��m����92��K N0�L86�s"�bP, B{�{V��ŋ��yLY�Vs*)[�0]�-�.8�CTs�ܣd��VV��7�jZ4�tҴ$x����J���n��0�rZ�4�1����aU42�K2nU��^J��nn�9.��)�FU�{0�7WWX�&�: �����t%*&�]F�f$��r���S�2�㰋�{�I�խ7D�Һ��̹�LRѪ��賃H,�cypJ��ئ.�j�6��Y�t���wre�iH�Qf��Q�|g���K�;�E��zb:x��;��$���l��DY�;l�o�Zd-:p:����-X��ۦ�00��?Jn���挘1lJ�tԼ�?eL�@[[���8�K��S��v�$�e�a�Z�lM��U.Beam���HU��k���v�n1���e
˭t�ܺ#p�(�\ǁ��FH8�Ӕ��"����n�L1ٴ+u�aR2�(*�ak&�*#Y�d��e-�uu�l���+olVMہ�B�Hn,��inf�50$�+i��Ȳݲ�ӭd��l[L��,�A�$4.��>#Uh��wSAy��FiB��3sh�WN�v��a`�
i5f���Kp�C��)!�"n��;1����4"���@�y����P0�6�+q���5�i��XJKQP�k���fۇ(�e�{z�nŪV)H����b7��uky��@���%D܍`ݽĉ�R��pJ�S�0qc�-�7F��Wq(&n�����@����@P��}�n4�cܨ7�4��5�2#�'�MS>Sv�V-�Q��ϭ�tht�֮�=N��E-�YJ��0���+ƥC)�F���	�c^�/�7�)Pͨ��bd�ݑ�R	W	%��Q���
)fR	��41A�1h˔�iz��,�v#ܡj�8���2DR�e�Ҳ�m-�Y�+�jʭ�H�U�GU�eӂ��f�}�.ҕ�����WM;��\x7�+�������@Ab�D�ߊ���QS6�m�aڤֳ�ŵ��遴�:5e��T��n�j�Ef�d�[e�
�eJ;�h�&���`�K`R�7u�Q��KelC(�ٗ��P�Pj�Me�KɎ
�ӥ�أ��r��q�&nA�SRu�ee
qe^�h�^2���,�Wk]�1Fr�����3[�eJj����cqV��i⻅(�9f�@��5�[�"���h�����[шm��ݻ�Du�Z-�U$6���i��b�ϣWX���-v&ԭ�n����WzR�Z�U�Ö�/S����3dF�.�����W�K��.�c2�a���IL���o7C2:�̙�S�j�[�w5Z��V�=����G^���x��e�ͺ,�����Hv��F�)8hd�Z
�f���Y���V��l��176X���&T����$���b�tm����׎��\�F�n�hӼV`����*8�c�Q�j��P��ŵ�a�5�-�r w@����k��S�Yo3t������ǨzN������"����+>����Q��l(P��!0�S'�JM����bFqYG ��]��I:L�4;�ݥB �ӳ����`]:�.�on��8Y�q�&=;���$}�TtU��sJ-®�I+�G�2�Q�Ekt60 �:�wrB��ևίd	�g1\Ks�ߝ����;V��M�*�+��fVj%i�,�m�l-ִ:ͱw#q:�Oq�lӳ4n�k�.Z�2U�]Y��R�`�SZĩ7�tM�R-,1�3[���J�v�%J�3�NK�I������*S�sUbv ���`K��Oc���ث͠5Í�,���0�$�R����`ۉ��1�i��jÎ��(���4v�a�����Dڐ�P��c�Lɍ�o|P�N=p�[�)�7d����֝0
0����������8[ꭚkL��J�au7%]6Edx4Xڸ*\^&Э�p�Uy�T.n@SOS�2'�oj���̬���,�0Pȡwj����&�$\��*%���d�rb�כ؀�0��X!����㼒v�[�*�4�Ȣ�E<L]�B�KMVBp�9m'��W<����7%V��e��cH���+)�Q7�v4��`Ee��gomM�A�y��az,l١|�ee��h����.A��9x�+��������ٛ�L�kc�A� ӱPR'մ��ӭ�lQ˽���҇*u]DK�{���R�cQd�
&�B��ͼ��n�o5�,f��gM�ȄAӿ;c�	,�J�ɳY
��M���N��e��8���M��U��IF�oe(���űi�����Ƅ�t�	�.�xXW�2�Q6\���:v�5vU��̫L$1ɕ��E7(@\d��f�L�U"q�H�Z�㔀�t��H2FlJ���I^g8���f�&w�-���"�;#�q�Gu^Bf��f�	��/i��[J�WW��V��W��u+t�nX/
�H����p
�Z�vK������t�}r���e(��L���h�q\�
�e��ˬ7Z� �;{WkZ�)��Z�[+h���E���f0Y�RGt(E2�`��^�4}�(�-������|���|S]�W�)�2k�[�'1j9f�Bt�Z@�W[-��9F�u��2�Л�6���(IYW���Eƙ��PY"���"�@�E����R��d��1��CqU�;{t-Xo]�FE�o˨�uy�,���a�Q9h�f	�~n[xmTɬ�PJ��ײe'��/� ��x��e@�� �� ��p�{���� �1��hz��$��D���݅�t4��7�<��1m։���4�d;XհG���V���]`5��Q��ڦq������ݓa��b&�S�L��V[��%��R"��5E���ud@2˖6����Hi�Z��L�w5�����
Ů;��An,�Ѻ�n�m�����b5w���l�.��8��ZE�v��I��Fd�߮�^���Mf��)�����dπ��ȫU0��p �����eY�i1I24�n� ����]U�N�#�5�Q�ֺJ�R����8���"�c�Oh+�u�F��m���Y��r��
�j�՛A�*�B�ؔ�=H���z�[��2]���4�����&3�X��je�іk5S�����شE+�53e4�z��LF�p�� ���%���,�	��CR�UD�[ڑ˛��JIJ׈��ȴ����7-Z�HC��vcb=�7Y�&��^��Hd��M�\U���We�pKWP��*�z&�n1�.��5�t�k����L�+U�t�k3k�II�k;k(:�f���I�T�Ej�iwt�r�	`�]j@���N�D�0مU[&��\�q\lҏ\�!P�5�9pU�xh&����S	�w���[Q�1�7�S#A[���8��( {�Gv$��\e^Dv��P��(���R��S��R��+
e�j�JR�A�P���W$Y1Ĩk��R2�N�X2�rX�4�Cs*�z�A�0j��.Kz���+{��݆�-^3��1�8Y��h�
�C21۽D����:�y�YP��0�GVV5�9-n�T�ZKTա�M�����G�Hb��HRqP���������9��f��U����VHr�Æ�ɪ��q�7�ST�a�N�d�GEI2�e���8��X�t��ԓ����ŵq3wr-l蹚lS��0�m"�-���`h.�A��L��V�6d�ś5������KY��B��;m�_�Cn�Z)�2��FEv�m���r��9x���Bl���!�H���7+ �L�M�kqƀ*ɹ�9ow��6�V���۲�<
��aP��t^�{C][Nm[�N�wpm�Z��@�f�D�I���%�ū6$#˛tҺ�t�z�҂�쭺V"�C6�/�E] ���m:������Gn�Sr�8��dh��m�G%yj�O�h���� ư9L��Z([T��x�U�n�㈣�gx<��T��P)85I�9x�����Ҙ��i�mV��2ø^��b�74�4��ꚵN�-SE�xY�max�RK�'��S͸Yv
{eҎ���';;� ט�
q!�na������i�X�f�/id����z#Z4���6�[4�`\:���0��b�l���O	���A�]�j̧����GmdH"��[�eBjRYZ�5CSC���^`�p���Nn�a):��-@(h�6+�MCdu�N�5F�n�ѻ1D�a7�or���b���X��N��eH����1�.�&%�	�ǥM�L�ZR���<Wb5[�#���q�3���f	<L�*v4 d�����R��El�vp��z��У-�wmڨr�.�4�m�%e��6|+�{sR^k�N��%����˼ ��U��� �q�5��a�rQ�pR��U��O(3�2�(��tFR��l���v[!'G`���5vfS;��Am9��cnX���1T �ߠ�U��L̽X�B����MjӤ��ǗR#T���7F�����@�^�LWhY1��� c�C��z8ť�ݔZ��Y�����U5k���d�X�͖7i�ED���_B�n[�5id՛�0ͫ��e��FtR���Ú� ���PT@�X�nhqX��n��W��W�:
�ֻ��F��un�[�F�U?���k	��<�v��,�" O��wr�2�oT�VP��1��Y&�\jGb�^�"��{���h1+r��j� �� ��,5eb6ɴwV�\�&췮���֕Qi�3J�HÌ���)l�� l��IڄT5�a��[�5l��d�V�0�K�Sj5�[�;��I��6h�[�x� Z$6���z%����Qm${Y%@ՓJE��n�h��Tݑakn��)�dS�@K���Ֆ��ŃAY çS��m�X��Gè;@k��3-��)BZ�ټz71M��B��V�H�a��[��]e�1���ӻ�J�hb:�ٕL5i)j�����B�]��d;C�(=c	w������^Jg0�KO;�/oi��04�1�7[�-���oX�h�i�VX���)hb�ˠw�P�9F�,N�p1�Yt��x6��OqU�B�Z��bVn�)���v5a�w��Q�=�bx����ǹ})Q�6���Dݻ
%lFeY�Ӣ���#r#M���m*ɕ%��&:V����:0"�L�#LxN'x��F,��;�&��ِ'�
QJ����W���+
��)vuC*J���ۡ�w ���6�ںS%t&��z�O�;��HoB�d�Fa� z����V���Sa��M.� ΅Q�F�YRfV��Ј�Xp�v�;z�M�!��?���Z�vDơ�A�gr�#l"6�Z���I���oh��!���{����u)��Ɩ��x�A��5�Ѓ�s\�g�<qdL� ��ywe6�=ŁуRf�w$8��9b�,�nC�ܖ�.�\*@�Q�P�N���b�e�UTqV���
˅��<�[+2�T����Fc�#4M��L�B��kiV���v ���7j�k{�z~:B5�t���ĥ�e=;F�!�ౠ�q�YN Ўo��ܸo�f��(mZl��CLӺl��N7��&��Qɏr�#�zP�T�6�R�2�ذ&*��:�ћG�hVSj��(�2�h�#	W���J8�Yݵ�TP�X�JQ7�!��1��l棩�ݧ�i��XC!�����ˢ̴��*ͼ���Tl��n��P�����d���Ҹ�#y��s�1��Ā����"��XU;�dI�+%�e��p4��L	�f����x��T�F]H�8�t;-��eGNm���UxV ւ��#n�4t����D��5h̗�m�*)P���� �;���FV��'�Xx�l�S9E�2��2�a������սى5����$Osi���-h@4dI݃35-��GM�3^�W��@Vc�&���@��jeJ��ʸ���(-��ډ�z!
�n=��#V��Q�B���چѹ��ַ6,�'t"�j�]˃)�Ç1Ө ƚ�f�h͹�2D+o��#�3D��̭��X*[n�+�Z�֍x�)�A��h�r܆�t�+�`�'I�:Ba�B!trQ���X�A5D�N��l�+/iVm�V^�3Q&���ߥ=�f��Ym� $J9��d�q�G�V��W�`Е�����i<�l�/;��r�64�+	�`�专@&VǑ��s-��17u()Se��5�*Լ�,ja�X�Uh��emf���v�5���٨N��(c�BlF��"���u�as3#�';YZ�1��Iq�fMg1�]ғAf���A*��u2`�Q3��B��V���,��H�ijz��3V�Z.��Szh�BX���c�bպ;��)
Ko�KQ��
&�J�6�O4�A��|b }�.q�rC|�T��Fc����u�{���7�FoWb��&e��cS�,��Y��?�n��UqR�ˎ;���mwp�����!��ޮ��ڃB�$���/D۹K�L�gcjNv\O�w|�}��ÕN�K����%U�-�A�mΤ�v���]�z+Y6�򴎛�gi���T����9Cˣ�Q"�8)�Y՛��K�x�.	���D���۠os�"S9r�e帡5�5T��p�M��H���=;s�'��.S�ۣO��w��	�/'~92iNs����yg,L=�$�3n{^�Eg���ۗ������5�S��`�;r��9��<�E���P@S�(j���[n�}�,ǹ8�C���[�W*�5kx�N<�7�5�u�K\_ʰ�Ч��&�,��/t
�fx��|�|����w���!�L��K ��+_<OG]�?�k��{OS��50y����C�J(ͮ��4�������`ݽ����ﬤ�ρN�wSo][I�!���'�,���0om��^h�̡�-�0���y1�No)�Fxp�,J{3�dq���W�_n�߳ay�o�8.CM���]�qK��+�;�kOQ{k�ނvN�o`X��o74;v����7EN���-��13z��9�cBԵ�eb��ˁ�0Y���Um�D���in2�'UY= ǹ7�n�N�>2Ln����c���5��Z;*�kU�ٚi�B�ͬ�x+2����5��{:<j9�Ts�m�G�%tfm���mvT�����WQP17�\;�9u��j��f�*��ͦk�����ċ�h�;@s4�.�ⳖOHV�6wk�7��Y�A�������U�n�Ť���4[�H�|�~�MR�wܮ�m-U�d]K����Os�1Մ��F�Vݞh���^S�����}��\.{L��R�(c,�Uw4���8�*l�eӮl�>�_D6r+�ap�b�R8�l�]�͢�r��j�8>��Y��x����J,n�����?`IN���u1]e�32�I@����/{���5%��.��ބi�4�jj�+*}����wNfC����̫�9�k`ɬ��}�h�n�km�ǔ�D��!�S.�Vq�n��W�'����_`ozM�3=؆S}]mZ@s�/��j�;�U�I ���cF�w�;zD�f��4���[�R��)2h U.e���s�-�9�uzeB�w��erD�Ս�шa�T���N�t��/ �莎�ͤ�ҏ99�]96[��V�oNga�Ғ�`-P\W4&�/̫�J(����kJ�呩n��e�c�\�O���-�f����s�X>��51��SX�U("��.��{�b�f6�\b��y� {}����*\�.8
Q]<u�9)╻�m�������WMv�Uzz�^G�Q�R�soA9ᆲ��PP�n֫���^���o�]��洔-�����q�dr��WϹ��qųG,�����l��������F6!پ&˸H����Z��ܘ�� ;({hgg\����(=�Q1\Ke!ݫN��(l��{vJ�B�wW�h�[Qȷ6�vM����Vr��ce��5M�H���(�j�L���1��<�mYZ�Τ���6p,u�=}J�	�w�L���ee���}�O^�{�n�����VR=W"7�}���,�":��vR5̼�H�\��Uc��]�7XR$r�BZ��]l�G���Rw���+���(4��W߻/�{��jS��KK�e��0д�]zxS��^�m���״�n��Mh	�����Q ��ᴪm�9Z��m-��G\Nw>x��y��G3`��w4�}�]���ﬃE����YlIS6F�s��T(�w��*$�w��7 ̗}��!ղ�=��w��[x�)�kY���m��HT�og�y1n�����ݗx�1�:PƬ>e�m�v�7w��1'�)���\��.X"w�gѲN��2�b��I���/J�0Eue:��Ga��N����T8ȫ�+o���o�y��Y,8Z���@i��u�+���s� Be�}��ˡ���#��Z����͏\����0x#�X�51x���O(µT�C6�й�Cn���=:g��24��Z���u�9��7��zr�9�z8Fs��}���m�B
q�pS���%�kn�g�NG�z�C/��sJ��f�Є|
1��E¶DWih�h�3m��
���c� �e�X���YpQФ�9u�A��ݲ*Y��΁4:�֢V7������:���!>6ޔ��:�n�����'Ō;�P�{0���k��!h�6���z%m0"U̫��f�W8�/w���)�^�Wǚ`{
�Ȓ��63�$�^�a"��oI��ݯ��e��+�n�������y2�I�.�k���6���cq1t�K�1��ʧ���-^�p�����l*��DLYD3���[�	=n{٫�A�����g����r���?Tif�=����	ԽᎤ4�[ޖzN:_/Wps�=�k7}0�\h泭t'xWyz�o}��[Т	��Y[�g�Pܫ�R�����3`u��hb�V;m�_H�V^S���c�^Y��1���C�j+N�������5��X:�U��cg���}�pqy�SX{M������G�n��"pK��S4����f
Ƒ�0�4뎉N��c���J���j�}-�̍KwX_Cf}{x�V��gg�}�����MhsU�{m@6������!=r��u_��"r�*�%3fo=�Ϛ4@\�0RY4 m��%%:�켣X7���ډw��G�Z��ʲ�w�nY�@�i�=�x�b̡�hQ�� 완���2!]�6�w�c�+�ݽ�+�6��3etFZ[��yQu�+18!�&�M�P���ŗ���Fj-�44��ۨC��̍��C6�n:�̏���Q'�b��iw�}�D�F�un�s�,�WuK�Us�cB�h��+��0q"��s�i��&�*h��cxtVCq��]��>�^g��jvGF5���}�t[��n��v0q�� �~8i��ʆ݋�#��潡w��m��uG.�n���hJ+v���!��w�o-w����<�KQ �a�ٷB&ōql![�s������(��ᛕ�6�]k���nQxU�]*�ԭ��qmЕ��5,B��s�:4���x�w㵿o\l�ծ��X�%i�S�5��ٓ.QZ��P�2�&h����9��A(,��GSX��9����:���q�7�{��Ҏhc�m�b��y����>ӏw��p��R�Zy��A�*G�sBQ����%F��ŤǕ��,�\�>�����>����(U�Ǽr���M#ݮ���T]�4Y���V�����,�4�m��L��{	[H��Yo]���L�ъ�;ME+e��f7a��/\ *վ�Vm,�i����.V��j��`J�K��Xe�v(&�s5���'E���;��y)G�>�u��I�%�''ͮcv�B�I�9�vվ�I�}��ʔ+6>�jě����+�
z����{�Z@d��"`Y��e��lX�SA�r�z���;�*�{���R*c~g�*�fd��h�����O�^Dmc��w�^͐�a�n^�z�����	7�rG��!�Џy{=Df/o\s�m'��v3�i��ln-T�$�����j��O(� ��ȸ6���Z�x+���AXP"-�NRt��T>a&���p�6��p��mDobn\V�4y��b�Oz�����
�M�m-e��Jr��i't٭��;����U�z{�O^�3���D��񇼋Ʈ8�d��\U�%�(jao\��؆�gqSI:�B�fn:�
��Qs����>��z����x�N��T�-��X󐎛�ʓeKO���ztΞ����kE���. �r ����B���D�Ղ�;�mTyq��W΢�j_d�r�*M���sx�Y���ψocL;��������Du?��0R9�+)����PNƱ�=�"�d��U�����.tb)Q�{f;�{�M��N�$ė��5�b6v�P9O<�|B������S����[�i�ݶr�B�q�L[32M��I���у���Нk�m)ԗ�%�WNlW��1ء}��b5l[ՖU�V�
|�@�F1뷝�q�wwa챏F�����Pɢ�k0)��"zen2��{wf&��{�n��tӬ�#��m;���V>���~�Wv�˕�j�s��.CK0�
j��OKѫ�d��5|��yd'N�S\���SMu�j���Q��݊�8�ElS� �=n�9���U�*���E���V�q���OE�άMX����[߸.������l�L%[j<ɽʯc`��M���9u5�F��`�݀�_U�`K3��-���T��$��L��;f ���%��=yn�r����Lu��|Քq�˰�o	z��SΏ�zLT���x�p�����L�J�.+��Mk+{i�/+ucw�l�$�Z�r��Cy�n�6�zd<��[OL=�X�ၭ$��s�;T�8+\�4�s(+|0���r>q<��Y�\��u�9��U����S��f�[�>��/����u�"��'4]
��^���������]��YF�^�
�EW[m��;�KJ�q�^����ؕ�E�뙓30D��t�2V����%��/b��E�D��1���\w1V��<D�*�1�{c�����H������q�n:�yUWL\�5%Tý��CZ�/Y�>~糸�p�% m�Lnaf�E�E� ���������:t�y!(�9Z�}�%3�7�2vv��[٪lp�WN�i�[��>��!�^����֝g;�M�eow�f� �I�>�ٚ�gv0�uK�q�Xk���wsG�Ay{A]v�>��噚� 	Gه�d�67��jl�XK�İ�I�o0�`���Qݦ���p�6Ù:��#�J�=��P!�=��"��g삮QJ`�,e��^h�Z:EJ81v����,��Xd��n�R�K�eN��M�@[Yq�,�����u���|N."�p+=��=���9p�>y�P畑���
F5��7JvZ�%���p�f`�&E��l����t�j��ޢ5��+Jr��EdJI�F�-EKo[x�]��nU�[.סu�K�1�Gi��N
�B�����fŤ��&֜ 5[��ҵ-P+���hÙÉ��b	���uy�fE�ABw�u�W��b
���7ULq^��-�U)%��K�i�zg���Ӹ�S�;���D��P�wx�Fw�^Дj�w`��n;�j�;ڏ��cZ�p��:�xp�P;��ɶ�`�r���FMPn؛[F��� ��V��^>h(+��t��S�&�}m��ε�:�E�ݴ`ᇬ`u&����rN�v��ʭ���8�xC�_[�l�ogq/'��;�H%s���\�[2�$c b����S���7ƞ�(�8�䲣���Wh���Y9�V«O���Qc��ݥ�ϯ�c��9�Z�����������nWm�p(�Jl�݂����X���+>C;tq��=6�GH]�:�v�F���m���6�a_WE�:k�4�z��΢/2�*6��Ηr����t*�Km�yA<�*����a���=��`����p�(R�4��X���]\�4�H�n�$��V�}�Y*�5H��<0�G���A�A���$u_'��<�hы����{��]{z�|h����>9ڍ�-��1:z��V��6�^�� �z�����|%lS�N�H�^���Lk���T�o�+�-�rӧx�s�!#M�~���ȷ��m�×m2]��yp�h[yυ���I��N���{�T�Mx%r��է���ݫ�	S{����VN�
���7�^�i�%���l��� �W���1����k4��)�����ǽ�|ۭ���$�'2l6��1���hծ��f�����u�1��.�ͲȢӮOi²ƞV��zK�
�wn��Nl������@�=N��u�msT	QZ'�,��5���=p��q}����,-�띴R��k'r�yԫk_p|XHfj熱��.rrf����)V\���j����]J�
wT���p�Z_eۚ�[�噚fCb��Iv��g��a��T�1R�P���b�����/,�;u�K��Xjy�{��띁WS��G��,J�ޝx��Z��z�;����]��{@84l�3�$���F��]w ��q{9G������S�F����[i��f�9�%;7��q�"5/=�dC�VE��N�g�Svo�}�D���4��(#@�lEh�مR�t̷�˭{���b�{{=�#˫� �><�H��q��m��O�8/�ߟ(��Vk����Q�@b�Uyyխʂm>�7���X�B"{����\���杫�i��l;*YRu+ ��+h��H�;��ٴ��n l�)+��C��8M�s.��u@(�P��h��0�l汹�)w�1��zf�6ܘ�3)�Q�7�j$_[}�82�����"�T����u�(���0徖����:�7��=����ʱ�ʊ:�Y��s�l��a�{����l6���~6n�����Җ��9٢�Z�2�����K�φ�}���p4�4�����܂m_i�cNE"�u%ю�Vv��#l6m� �VM�
��
��x��\4uK�B얦�f�w��U��/� �KiS�>�	.��p'�}����Z�&^�r��'�/v}�s2�ku�J0�l��hQF7�]��7�h>�����`��޾=z���������nPX&t���6=�R%���^7�~�v�85/|�����>��I���BH@�y�~fp��)P®�*�s/��y�rgK*���t��5E]���5gO�=�e	���3o-������`>	���Mb/�{t�^ʲƥ��\qG��Wq(�4;��1u�#����^�&W�X�5=sć��-kle3�!<.�vT��[P�������3�t�72���چ���wq�����u��<�#̐�˵���i��h���%��� �ܭŸ�Է��ns.�����骱�^�|�T�ʁ���߻D6�:VǚLFOL/Rj��|�;����fF�Ax��LXQ]��<������j�wZ/S0GC��k�x�o#�q���7v�K@:w����*��@��|��n�7ፗD�>
+�5���+��1b��,��j7D��X�sF�jC,�{��D���f�����r�Ycq�V BDڙ6�fu�5P*Z�,���̗��=�c'J���I��sg�|1j/u��n\�x�tF9��Ὣ�EԶ�����5������6��[������sXdǼ ��C�Y�m���ٙ��_�Fq�7d�7/j*j��җ``#	[1>،��J�j�տ�:vۇ�|�����XSr�?v�Q�{ݞAǈ��2^�<��=��;N��d9�ӕ�
@tQ#�kT@ޔkWY,�>V)�@�ԈLN�Ӎ}����#+
U
��Y�����I�˾�]���3D���5�ݡ@�)CkWksR���]�\�lxf�C��-C�.�2��
��T|��� f-zmi���0]5s3��>��Ӄ�ӳ�!�d�ƳU�%�4§n�.�'z�v��6��N6k&m��$�v�E�DL��_ ��c�p�F��Q��w�P��� �'��J!�L�z���,j��#U�IG�+v���N=feG|mq-x ]��U���^�|~I�l�e�T�/ˮ��"��vS��:�D�V���7\y����l�>�L�4��Ҵ�vV�Z��TѨ��t�:�F+#��d��o(����bS��Ld�o!�Q+CFQj񣻋M̴'9�`��<֧n����y9#2��ɖBv��(n�+#�LC8�](6��7S�m�a�<�Y-#�n� ᘎ�d>�f�*��+qO��N���kE+�d�G��iw��w�t��]m�B_uwgjՑeں�h����)�FLX�#����+Gtޝ�n�eA�,�z�}m�O��rC����c�LЋY5R�<"��j��r�{�M��︴�+% A[��vʹ���ܗ�SLZlѭ|��d���>:e���(J��ܒ��J����b�Y�|X�V�<���7�jL����I-<L���A}���v�TċW���гf@�h�;�{��q��|A5�>�R��ةoI���R�P����L:�dR��EB����#����Ί�޽�\���9j9k,˭f�r�E�K�0>Gm�X�b*��֚�d�;��TD�fU���5:qQ�b�nְ�g]K�܂�a��LV:RO8E'��D�q��Z�н�m6V��*.�1�F�ųZ4��)V��;d�[����������֜�J��JS�Y�mq�3o�ަ�[���M�E~
KVm����\�س�1Z��u���P��3A�c��І��%/a��i�}&ۘԛ�����yb���kQ�2��Y/8h��Q��wZS���|��`��a�3�f�d��5g�e��N~O&^YV��b�nZe�=�/x��Łn�&�VTɭAxq����͠9��y:���|2���.*}���������
y�ya�	`b��qq�Ä�}�X�u�wx���CX������6��ٚ1�d�b���9�oI��Xؤ�ľ�QȀ���&�e��B���M|�Ѡ�тR�.�t��7,�K%�Ϯ�ٮ9���ZiF�('v�bTmRr*ƈO����փM5�]�ẹa7ڂ��N_��թQ]�&�����y�����A/�Ö8�m]� 1�R�]hUweu#P�V�})\]�r�L�j��v�J���>*��6Λ�mqX���j�&��i^��<��we�;b�!̽%i6�f�c/+�MZĲ}��b�^Ü�]�]�5����8�3���Nɯ��Y�����~ܞK�`���WC�j�f�Q���(�cfa�7W
R%^2{��ө�r���a{��Zh��ME�����=��JcpPI�B)V:�vM�5��iۀ`X���I+M�8vx�d拘���wp{r$B�C��4l�"�r��$nĒG�.[����AOp}�i~g���z�ZI��S�C��9`����R\�����i��5i^m<��Y�7c��E��C��V�o�[�|O^佶��w�!����eጽ �7^�(ú�y���b��]���C��X�<����މ�|�=�S��ڍ�� �v#�V�������fqc�u:���&`�������ݵ�*K�����5�T�(q��S�R��u�� ��7�r��O���[O!����^�E����λ쥷(�a=��+Y&���*%Ĝ'Ӗ)ulo�C����z�e�+��ww��Z�j�G�;nR�TT��ty��F�o` ��&9&�볊h.ɂd �W3��x�+M�tv*�������iG�'MO�RH>ćt�������"Gn\�cxN��yj�V&]��&��r��X�.��S��y!]��)Ι%t��E�V��ņ�f��r�|�<[%��|��b�,����V�EX��u!�<���pLg�����MJ��x�U4��3ќ!���:h�)��1PsO%�e�ر��H3S��S퀉%iocvj��<�ɕ��f��7X�������q�\�����ap�H�/3M�}��W�!ܦ���e�[����9����Ƕ�U���v�O���'i#}�`ΪC���qX5um�����ٜZl��~���Q��7( �\��Kv�`ӣS�A�+.l�5s �Ɖ୘�U+�ʚ����e��:�;2�a�=��y��=j".Ɋ1�2��}�x��(a����D|��W]���U�Xw�JE�N�̘��2�\�g!�I�lⒶ��=�5K��+�{%�.��k4���TS$gjhb�q�Ñ�sl��6\�[m�Wwp����O	�t-&�����^����N�vNq$�i_0TgjreΤ<�pɽ�U	;
��x-1^G����{��6�J<��vP.R�FVPH8V�^o���V�=�o����fˉ�b=U��� �uJ�:�&��-����c��Z�9�V<�`,�)}�SZ�pa���(>�h�k�����j�i�]��
�aۮ5Ԟia�-��>�R��/�@��b�d�3 )�{{\q���%�{Z���ѳ�b��Ų���8�;;S�=@'e��'b˃ƈ�ա)uw�mk�\Lxgu���b^����Ĭ�kMJM���e&�JU��'k����z#$:�YA@)�zr�5F��X��z�*W���;
���6�����;���9+�e]���7	�o��O2�9�f2{(Hd*�ǘ���{�eŁ�Ʋ�;׻�gb<����q�|w�wm�xr�ī�F`�#��VRW���$l�q,�nB�[،X�ʗg��k6���i��\�LP�����mnC��K�:��j��`S8n�9ՙD�P��
0n*�d��˯�au�)�1s\���fj4�g��%�1P<9Oc���"œz��PC��c)/#ɕ&j��������!}��z}}O�+շ.%�擧Ax��lλ�>�:��ػ���Sڳ�9�G+N�=�N�L��ӻ	(�=ۢAa�qW�{�Ǵ_�
�s���8����n�獊Qp[�w*Q����4x��Jo5��zy��j���X�u4T�@�;����n&egܽ��=�y�✫�V��"�eq��bCi�;��)N�(�ʴ���n��cL�_� �שzh��Y����y�<��C�}X�s��zsnZH��L�4:p�~�F�OuU��<c�
���yN�9kh�cv���y٨'�VNk�GW4�=y�6�nnjRLY���)�]�9��v^�{�#6_S��#�/�x��mf�on�j�&֓}qD.��b������]R�c4m¥��6��cX�1lAL�G�-�K�) �U��#�Vq
�h�V�!ŭѦ��h"e�����i{�S��r$u����^�f���|�)@�ę��K���r�������
�^�56�-�ͳ�㹥0K��H|:�Ү��i�3e�C�)Ř��b���7*�y������!Gp]�Fh ��*9�6�`L=�}@-z�������{�.<�tD�Xf�+�n7u����}�>�d ��^s����ŋ!NFim�����"q�D	9'������^�zs��U��S$�PK����j�d���
��L�<\��ԮC�s�]��%�	���NC;:��Z��D'�gn)�g�K�r��������\Z��7"���}�4<��[2J��(���c���z���?^�vHL�X�(u;֜7����Q(њS�k�J�2t��.�ȶ��3^�ڜ$X���UׁkD��	�-��Զ.���s#��"�5Gi.Hi�r�B+.JP���� ��񓗻,���q5�+�O;ZEs86��v�U?�s�P�y�ӦAt�)�tE���*WQ�t��!��.�e��]��.Ѭ);0%X�z*�B��幺4M�y|mmD�X�#�i�[=/]�6�D�y2��2���8c����vK�|�fj��M3	:�cR�߂sd8S�)�&�cm�BB�u�^��q�����O&.yD��}$"�Y!�֟s%�<w0F�J��i\%�3M �厵eLɔ��n>hw�:�'c:R\�vt�K8�苳ɼ��Ǵn��*5*c�d`�8k+ugI
�;6�����F#��b�N�ۻy
��f�[�pʺ����7��:t���� K�v���Y�v�bu�Y1'}#�*3h�+�Z5��S̵���r�'�5ٵ98"�_ax�P�]md�V�4.���Y���d4��{c�r�def�4*�:l �ΐj;*J� �#�ϧnP�Č�75���o�;P�����NA�:�5M�!̺&�+����5��v-�-;%s�:�#~ަb�a�䯳΅�0�;�Vrw��U�*�f�y��%c9����p��jW3y`�1ƪ]\�٘6�1��U��n.Ao	����c]��N���;�gVپ<����yL��+���>��N�Uiu�q\�?��mH>|�wS<�)����0�V �-ù, ��.&��fJi-i�1&�|8��O���xk���S��5�N�v�<ʄӢ
��Z9��#!�9�š[}�y���yr]��7]��G�5�nZH<=�s�2�'K	�k�R�2�v�a�Im�Gw7�1E��qJE*ꖁ哏5���9�7dZ;LL, ���i�O5�YA��?��]{E���:��C�r�P�t���ۧ�X0����ZXn�y�Y�b�(Y�Yk�0��087(n\3�n��r�	���Z�xa�p��m�oSL�hjGn ��TX�ڤ�`�c�� �1���*Ξ���]b��qJ_(z���'�ьhn�L9*��H��d�ڱ��o:c��I����*�[�3]��dF��c��Õ���'�<v_`�\�&I�x��Ӣ'u��K5vx�_-	O� �Y���A�R#.��em���Gw[%�Kb��"yB�d_���}գ,�L���;4:q�8�jW�-�b���@��\��7WkWh�1���-�[�M��T�W�hQ�i��ı9��TӼ�bx��r\i!>Z��]o,ߞr�)�Z2���<,uX�vwl�,V���Zl�L�
�vR��J��fΕX�%��#)�3���8�M7���(��k$��%�k�Nd�Ջ��j5�q��ø�=}5FD��V&+�H��U'YY�<b�`L���@0(�A�H}���v��yeWT��G`���h�N�a�D]kƽ�-p�K� �S����5G��`�ג�a�s��jܙCV)�<� 0y����[_W;9���m��A�2�I`���R���u��r�7�:'p��	�j��|7^��^R6!���d�m�N��l�X��Xa�Lepn���t5���ٸ�Zշr��D���%GP�`�ۅ݇�"���&��&��û �tx5��,嚕��}` �T���v�

	$H[�I�C��۹[�P��ISV��c��!z������>�c�Oa�{��ڨ�J$�	���嚜�׏~F�r��(-�G�d�اE������Ȅ�W���)5��Z�:�Qk��j�rȞ3��g�q-���{}H�;���47"-�_��ߢ�w,�-��fWO�S7F^5,'Y�ʝ��ڦQ�Z,Rm��VҺ9(f���T��;�q,�G���j�vod�2�%څ�N#���ذ����I��,Z�\�j	�Rh	��Fm'j���E����C-�Y׿N�]V��̡���Q��Y��-�b�Ӥ8���7Ӽªv}<�����d9�6�p#2h�0;3h��gze�8o������D�4��1E9,H�>8p?v(��}�O]�B�%=׷=�{b�(��K-
}���n�D�.������C�]~��}�;�>�V�44v��qKE,�xCZiMG�5n�����2pX�	�_W�}_U}���׾Hq�2V����*�Ðr
5N�����rH�{���J\^����R�f��c��u��s�=��p-K��b�;:�6A���������8�<�p38���忞�R��0��d����6�d����n/4{��Fxc�vTX+0�2���ؗ��曽JO���6���ؒa�-�E�="�-�nٵ�R:��ԫ��o��E����5�a��`'3j'��U�e3b�cf��`B&=��!�[K��ܥ��a�L6\���n���PJ���3�u��u��q	DWJ���ސ'�X؂Hպ�wu���/f}8]oTd�q<�;��PMfL��*4��Ff	����ݑA��G��O�j���w!b���RPHꬦ �z�d�w��.�<(��/��ݫ¤!�6ș�왖����kq�Z�qs�nЫ�7R��M�8��6��v�W�,e;����s�;F��2�z�%�
�9�R	܅[�%m��Q����a�Um]��yy�*T+��8wϊ�R�F�5q��%aP��=�1t��GeC�w#�@/87�+���� `���E��f0ǈ"��Xeh����p�jj]򚃅cgP��v���v)��=ǯ�'F��&S��cM˃��"-�ǳ�ӊt��������wJTF�`jwopm�{R՜��+a[��"L�F��l���%�x��M�j�
���l�TA���(��墖����[b(���b�(!ZV��V1��j,P���DDVګ��E��X3(6�[�Ub#�++m%�*Ym���JR��R(�E����[QmB�keUA�ҥI\d�6
)��D)jDZ%P��J��)aU[kK+e`�F��ij"�c�F2 ȅ�B�[U�b#SL��li`��j-V*[**�����ʌE�%U���V-���-h��Ҳ�TF�UPR�b�����[e*R���Gh�E�TmDR������"��UQB��(*�J��\�8���,Q�`��kF1Em)j[��o�-7�ѡ�c�Ѧ�C����nj���T�������h�����}�x��R�i��I�A���)�J��f4�}�Sb����j�4t�ct��r�i�0�*�[��5�Ot���7]�x��r�uW$X	v�,� ;�5Wϫ����j�������4��4�7i R�'t�}����摦�Z�u��y�JR��O�9!}��b���I��o^3�nIU�ZO@09iy�F����_�^�ToPkò�(`��
���^^�W���ټt�����uzC�ET#j�l?Z�,g���+I�^vq\�� ��մ�%��zE�^n�OFR��(������>oЪ�5A�0V�#���|�<���m(�9�u���n�E$�2��Eu��m8�x��� ���;�^����#](�-�K��O�>{T��Z͂��=3۽<�y�-�Ţg�$+q��"�.⾏��M��tR/��}�Q5�N�"��ܰU��sK�I����Bu[�HzWEOMM�7nac�Ө�U�Ɓ� �/V�ˏgV��sL�ѡƙ�ӡF�j)C�E�^�b*�����U�z4��
��z����b��	��(���4���eF-7E9wP�WR�WOXfv<��9�y;&X7�Mx����
�2K��1����/��;�hWs��k��Gmr \!��|�i������tӽ_��Y��֤�*���t{��5�S���ώ@�������yDP�,>o�3	^v!�j"fq��rZ��5��H�낫wP�����|x��ֵ$$���\��62�����	�l9�w�y/�GT7%3\�j��\)Uk�����du/���4��_-ś�Vą��*fs]�mTB�8ｷ��'��ՍF|���*H��/�uw_M��,텣':�s݈���5ou��0Nw�G�L�	Kh�Ц�wB��a]�΍�h��9�/Ù$�V�����%w7�hޞ֥U���R�$N��OC��>����yj�7�t������� ��U��,�J�^�l*γ�2��U�R^CO��Ұz��ܼ[q���{�ht4h�x��)�Yµ��<3�Jg���u�ό����ņ����BΓ��<���g���݃�	6rW�}�թZ�X<v����Y��5N��셎����z�5l���қOE\�,��,�p�[V�d� yY[�`�ݴ�j\[�޼��}ϯ� 5
��_:�w Q�k']�ɽ#�˽�F�u�w�tT�]<㩓k�e]��2iF73�Xq�1����ޚ��v�u���Ԩ�0z��9�a��ew��vJ�k��N߉����u��{�0��9�[2��Z�o}Q�X�;g�}nD�{eI�uV��J~V��o%�nj>w<}/��r�6x����WÆ�!��BS�Ţg��CF=�Ϧ�����y�D��W�����8�_��_�y���=�:t�Pg���+0r��*�l�~�EY��3�E�9��zv�U���a~<�53��ĽP0���8V���8`�דh�oj��/"��]~䏻����M>�7�=�nU��.�(�t[$���]F =��d2�\G��Tz�/rq^'p��yC&�8�֮*σ�[�i	�6�1����w�(d���̻킻���}ܑ�J[��L�6åj�W��T6Y��	������2Fq��q�~���_�[�~�d�Xʷ��<��z� "ɹ̡��8��
��h�,����s��S�P�(p�B�%�캺�r,e�����.�+��� ���o=�}�	�������t��>�v)l]|�4�ԍ����_w�*�ng�����蛹������m�Z��ʜ-$�طWm�h���ɛѥ��2�D��A�t���i�*��$9k��������c�2������{<�Ѽ(��b�3y���+�,�ճ� �8%F�3�Hv���*@���jN�6��w{{�����t=�ю��+����b��@�KG���w\w۶�x�q��>y��-O�]�T���_�UI5ER�\;C��~�閖���Fp͏��I���r�/�����#τ�JAޥ��Tյ�`j%C\���[#vg�z]���.����ݳ3z�Q�t��T��/�va$V�v��i����g���YՊ��k=1��5MsGk�-�pU'��[�ޙGug�rܲc�.�r�}]��%�bw��(�u�u��}�V��*��N幼���պ�����s��(?�[��Z�vۭ���+}"̝��z�ß<��W��Y5;�k��mWٮ6�+������npܡW7v��f�=U�\�A��T�)��w�I;}2y
�[T}r8����1���g��G+�L�,n&���:�V|$���u
�Z�]�4��� 4��6I�NrŔvs��|��������l9n^:C���GX�u%gN��$�΂;_<�=7��eV�s���{�r�);�6��&��{Ȁ��Ξ���:�gX�h���Hv����#y��u��4.��Tɨ�p�(�D�UV��ͅ^u'�ҥғ'��2�HP�^o7w+mU��r�ĺm]��_*<�_y㛲�y9�Dy��K�O����שޤ��u��N������#\�������x�ǻPK͆�1�{��:e�S�;=2�侦��v(�.�>�Ը0w:{����y8���m��Ҩ>ǕE�U�L�)�R�/��uM
:��ӯ-`�/�'k6�7Ӧ�j)h�[�{(���I���'��J�F��E����+3x��;��o=�FqOo%'��]�:����;bIt[�T�vg�ݻ���U�c������T��q�A���|߉s���c��tob���ݸ�zx�Ӹ��k����r
z��Ykrv�&?}��f���;��R/���Vf�&���p�u���1�/NA?ug��3�o�,��
�=h� I	��k3=�ҥז��y�ʺ7B����zqW��ߑB�:Zg���;��0K�у޿'���*��/0�i��M�r�8�ˇ{��E��ܗ���7�x�\�������"q����eǆ�.P&���^#8�����m��o�Q�#�y������OORu��~F+~�z��~E��9z�L�In����a����yl�Y��t�q�a}=&�n�k|���:�\����m�b��[��ُh\'ɻ]V�Vv�2�8�w�d{�d��}2y�c=�q�8<�%��˽|·2��j�p�(�Ԕ�Φ��q;�1����j�}#V��sU�S7��u�3����Ny�.�_>p*���m�^$��3��g�J�-�ld�%wP^:�㓉η߄��՜�7����k���2�O�/�;J齙��v�x9��m_�\F���uZz��4�<�{	+ө3nC����ճm=��9�y#[�,Q�cjvx����#,��IxL^]�3.�d���z���x����r_��NI�z�����y����}<��
��
�����vg9�(ŝ��H������4}�gK��]=���j���y�ݼ�u��R/�U��U�	�`	�5s�t�]�@�5����;&yl��S�'}�.�t�jXڝ���is�v.޽m��+@S���%���y=uu�5�b�S���m��u�+��.ӫ�G����9�b�����w���_y�k4hG���]��X�O�W�yԕ9_G����zV9W�4��
�kJ�)�����k�����x�=l�8{R���v�{=����ۜө��ǝ��fW���./{��{d.Q!s���F�<��TϷ��Q��ғ�Dc7����izE���X�|�N�w�&���׏O�E����n�������	1�G�:ճ֜�C3��9�{�1���ȑ�j�E�rym�j�]"���aOy��{v�Rc���:V�S�%-r)���/�փ����n�v�Y��;���DG���=�����Rz5��l׍�J�*]g�(<��h�k�ne�[*w���u�S�͞�Sɰ��{�q}���9�wm|}mU�[�I�ħ����]�t����졘f���F6M�9N�����رգ�i|>�3]�ռ�*e��^�/�l�hs\���W[�^s�$+��}��9�'��N=�c�ք'N���ck�n�L��o��'�7i�P�G�	6a-%/���-�>��k���I�y]���uw5�8n ��h/$���m���7&��7vǘ���yz��}�͆�IZ.�����ګ�3"��w�,-��t��)=�p$uO�����U��=��3�T��7��)�p��r�C�^0M�<�mo O�?P�fX�4m]�5��[U������\�OӎO_��ǭ{��x��SI�
�JQ�ݕ��qlJ��4+xA��#N.�J�k^���DhfWNf��~�w��A��Sqm�)���t��=:ս��ˣ�B���kzs@=��̣=:�{t$.Ē���9��3�ׂ��<����B��2��J՞��K�ޓ��c�!�ַ���f���K�ca��5�;]-M^���Y��?9�y\�C>��W�|m��N@������-[/�s0cU+�tb�o�=1��5L�s�ހ���R&���c(��q�NӹUy�rϾZ��g�V!��G{J�t�f�<>g!~o1���m�
�V�`n�H�|*<]gE����LyX0xf>%���|�=�<��Q��C��b�L�cg�6׳�L��\S�h�8�r����}�ۧ:�o��u�SU����Cy�R���}�5`�Ѵ9.�wJ��G�U���_��kޓjk��(?k=a?r{��fb~��\I���˲�m��h��裭�O}.L��������]t�hr�c^���{8E�f'�ӵT������N*w�3��$���<���Gyˌ]^&�z��E9�[��~���j0�����w:c1�+�="s&�.V=i�s7�{��6t��F[TN���8/��pM��d��oh�;x��ٲ/tj�[O�!��q[�Yo�~v�G�
����Q���9���O��k�xt���T$�(﹐��9�t�7�T'���"r��h=5��9ٚʟl��M�o��|�4ӱF��y�]Kƅ�֌��=y�<�:.wG�9�e�V�3|�[y�)�����������g�)�͝7{]�ұ�uK���fm|�Ө�	'�PK�^l�t�O^��$�}y#��Y�C�ʂ��)�V@��KvJ<��{&�6�唝w]3Z�_���Z*�'�j����{�V�+\۬�y�N,_U���ޮ��X�e9�ؐ�Cd0��+cଔv�BIyԵ��/�T�[}oWʛ����g�{57:E�]�m��wb�<�G���W��⏾�*�w�e�/qK���}�������U�V��~��2��c����̀���OZ��Ί�J����������S.�X����'&�iǖ�XyW�鳽���I~��^}J���;>�X�zm�)E{j��Қ��ܻ�<�}��/�왪VV���J{\���b�y.��ڊ�+Kݿ�YΕnݠ����s��3[�R��WS�WH���������&��]6�7�6@�����]V�;\��]��?7����-u��{��.�"��������^ԕ��l*�q��g+z|=Mƽ��U=�u�����y��2�k/�N�n�s�H4W]\��n�����[qu���9|���ԛ��^[�Grw�Y�q��p�=.�zJ��,YV���v�#@.Y��:�0�5���R�2 !�u.�۩�uU�d���o�Uռh���u�B��r���W7]R���&%�g�[�fg6������z���H�`�����E�%��=�!.
�/����/da�׽��8������=��zwn"r�ð�Hzv��IƧE��uyA�I�WQl/ �`�5��;Cڑ�z���鸌�ŗHi	Y�*��^�*��7��Z�������s�|,��w�XQk)i:�ڔ��[rn=�;�9�48u���e"�*rX�	��0�cH*,�]ؓ�Sr��U�7��4ٱ������,-(J�|K�`bڸ9p�����gAƲ�����'���Q�A�l�4~<��W���<C���=
S��/s��qz���M���p��%׮��-Y���})��]|�w#}��MWl�X1�u�I�=Z��L�{ ��Y�}�82
�Ѭ-�f84�� �����*�.�)AR�v�U������o�o*�s-eI:	���	���M5��>v��k%���
�;R���..T�K��*V�sfU��������n)���sN%�ύ8^���H`��|�ۭo�ade������'�3��2�0hs�2g�?_*���ǚ�g���:��+/g���c�=�y�D¦1��a`R�������֖�T�e���+�72��V�K��7p�=���P=��^��I�o�\���9gA�N�Cy8�}�IRh�Lzv���':�|/��w���`�~�8�1��u>"�������jͬ����(�ʓ�{}\�P��m��G2��#	�f�9�R��3qw=ۻ1Tݽ�6j�,�.���d�a�}D��<Խޮ�%�`U�y᳎":�t��b�|U֦(�SeL����T�\i?$��rqk*�F:����1���ݠ��. �4]mL��'k���+n�"����K�.��]�&�.�F4��K�T=�L�ۜ�sr
baN�ҥg�x,w�=�ʰ��3�x�ݔ�׹` �J�FCJۻ*J]ث���}�����>�2�!ŝC#����t�8��SA�ҹB����pI�Pwѝ>��r���ǹ�)�seֻ�]��|5N�[M�W���/��(N41�����k'迅��iW-�}F�FK�;��T{7�z�dϊ&��c"����f�������Tj�oa������ay�}�f�L/��S�tG&Yp�9�ľx�	l{�wn�u�W��L�֖;|h�g�<ՙo����Z3��-Ҥ7m��w}��*���g^���f��w}᜛����!;�r���fI%j�i�B����ڢ �mo�#�V7hzƝ�ɭ��_h��(��0�DYZ���L�7ϋ�D}����-�*őcZ���5�ZZ[EDIm��eX���J���Kk�+m��
ՈҔ�b�����԰-�-��ت�B�ZQJ5���H��(�Ը�\U�1m,U�#lmr����Tb,r�ċ*�m� �U�\�؊�+Z6ՊJ��"�[e�E
�"�6��
B��*Z%DDej�q�֋P[kaKV�X(QYm����V,��QX�Tii[YZ����"�4�%��hQm�V6��eel�FT��mh�J6�j�JR�e���(
5���jPkV�kB�Xe*�h��k)[B�+U�m���E����%m����X�kR�-ZV�օJ"ʅeTkj�U��Ѡ�J�*TJZ��PR�W2��K��R�����\�wG3�tu���N�
�RV��<�Q��u,�tԵ��Ю�w����Ff���x����\y�"=�/;�R쾚��V���q������F7��	]Q�k�̎�cjꆹIL�p���&�r��R�]��t͠��l�R{�v�+�iV�K�v ��w9��@�y�쑵>F��\%�������x����r_���0�Ľ=��ɛٶ�vl���bc�)�i@�q��漣u9y�;ǌ�G��3�=�ד�^�u/�ɪn�Z� ����W5�Ĝ��38���睍̔%�cb�JI��+���,��������4]y��'�-�l�>���K_8�*��F1�}]�ڙe�{B�3�t����i�����a�Q�s��S�F�GJO=Q�z�ϻ=��˙������W��S��/h��+�/�{�i��O����I�#��z#��+ǳm�O��=D�[����G�9l{�*fo���U�-Ǳ��6�����=�gl�`6��jZ5J[P��`ь{�z�����:����u8��3B���l!g�S���u+�W^v�}�}�s�ep�1���~^���h\O˯B)Xw��[c��/Ktu=���l{qj����e����C����Nxf�����֥y�����o�+egV���y�?Shx��6��pj�U���3ywH���Βlq�s�+[(}���6�Ys��р�w�^�k`�p��U.)��uԒfܫ�_/{���V��d����T������I��O��hU�N�����;ҳ��1���XѮ)<�ڶܭ����w�{Z�Bg*�m�:���i�*�8M.�=~7����nf��Wr��+��yW��W���~σ�=�.�M�f��Z��n�:Φ��~F)�y�m[dV}�m]q�k����=��������q�y)���{X>�8v���e�|�5N���Y����v���7��avH_�8�v���Pś�ײ��o�]?4�8]�jޫ��^��f�E�v�^g����s/k�Q��=�c�L�Nd���p]"t՟	�k/H7�5�\�\>��V�u���]r�ú��yv�Dd=�~�ŖvT�yi~���������YmgV_�B��m�{��7EԳ��1{vG;����q�c�rE�Fa��t���ιs�+��N��3�]�j���ֵ�k��ԙ's���gvS�N�����'Q�����Hm���^1�X.Ռ1�Uy:��ZK��S�wU�󺤼�}^홛Ї����t��_�.�̷w�����SW���k�e�M;Y�ۚ������
��qn�tT9�XLs�uf��k���K����H���N�Y�����;˜7S�Y�ʰ��t�g���|��uʯ%U�I�S_���(���y��JB��b�^����o��5�VjqS���#�{��s'Aj���To��y��·��㗲��=��ÕK�t����S��S>�;���v�d�a+�����jy\��θk�q�u{NgSc��|c�Yy�s��3�̞��$��G�aBT��-s�,��oq���	��d,��8 �{�y�ڿ�RRw�Ԟ�?��s*�۫���`s0�Q����6��%i��S��Zeq`!��k�h����[8����Y�!�`ǳ�-��=�h�H���E�f3a�1Z��e���+�%����Ը���hu����܇Y�'H���#D����`�z�G�oy0G>�^�5z$.�Y�F�B�+[Z�:]re�˪�NI�u�d������cjꆸ�5�q}��d���Uّ�wQ{���$����C��ݷ��t��ȝ:�.�s�C�ȧ.��zy�~���y��Gi���y%����EN�hW�X���k3$}n��wZ�ݺ���ٜ漣x%��O`�%����fֲ;�w���ȴzM~Zs��/��|���������4���N0��xB�d�=�'LN�����N��|��~d�����3濾�מ^��>�=�|��{�	��w���$�<�*V��vE�~X����2z�u���!���i�l;��u��WN�_�}�B��R�u�鿿#�����9���&�O��{��8���9��q�Ԭ5�a
��O�5��I�ߙ%|d���H�w��8�4��݆�8�~�j���_X��+��'�W�*�������m���M��y�a6¡���PY%O���m����z��>eC��T��~����N�k~d��s[��.���ѬW믾V�哿S��k۱�\����t<a�'}�f�>aԟj��?2u���O��9�:��|���d�T&��ORm'̨y���>d���䓨=�!댟2q)�o^t��s�z�u���܄�M�r�l'S�k�I�'�o��N�@��d�!�N��k	=C�h�ru4�>g�>ì�J���s�d��Nj����Oo���}��{�;_|~|;,<:|�m�9�^&��8�(�b{���o,k���:��0�̀�cU�))�
i�\X)�w��_lk��Uw���O+���*�NL|w�Y�N�;׺U<�y#�?g�P�]^�ab1�
׎�����<�������0�`w�N�'�N&�,���&�Yg'�Y�:��Of���8�ɯ7�|�:��}�	ĝC�gS�$�w�q����֌>���3�Ͻ��������'=��2N2O]g쒲i���&ړ�N3YBz��:��8�m�Oڡ�I��Y:����)8���?
��u����Js���%������O|���6ÿfd��	��0�'|퓺�$�I빚�+��C�VO�qe��?2q5��I�LC�,&���q��X��ߞ�w|���<��sm��$��;7�HVN0����i'Xy���xɶOO�d���MC���N0�O&k$�6���̬�1I���u��D}��*��j��F��y���޳3}�һSl���>��&Ұ4���w������5�m��ğM� |�'��Oxd&��&����VI��?d�&�PATG�p����ˇ�b�~;j;�o?}��iم�x����'�I��8��|^`x��N�C߻�>I?k��O?2y5���x�����'L���ߨ_������.ٕ�Y��F��]9O�*
���,;-�6�l��i8��Xn�'���6���C��8��h{3�:��	��so<a�'�_~A��>�߸����^�����q���d�!�氕	���%d�VJ���I�zaa8��~���RN3����~d�7�:�>x��ܚd�}_w���'��%���"W���~�}������?2zŝ��	�=d��$���IR��}N0��J���N u������'���Z�m��$+�M2���*�Ύ~����8��W�}���om�oǘ~d�OP;�
�2x�ϧ{�C�MwX~d�I�Y*T�����o�2��O�;���d8�}9��Uܿ2+*�F��c�w�6���X��m^�n�>R|&�I�Pn�ep�T�k^���20)��hv�/�x]�m38���C�:3�l�M�lwZI��@[WP��zɵ��O�"��r뇳�~�	xq���2���m�\��<���cj���',�)>���n��̜C��rB�I��x�1+��:ì'��;�I8���;܅C����S��'�?�O�'h7�I|�N:>��T������c��Y��������}<I��v~��'Y�Vi��L:�����'��βLJ��ϰ�$�����8������'>J���a
�ԟ�"�����A��M��������}�x�x��Ȱ��'FXm�x���Xi����y���Oq���2��'�}�$���7�PY&'���M�d5����x}��#�7w_��1��~�5V���ۺ��>�?t�q����M�y�%t�|�0�|I���a>gS��q��[���'Ru'ڲm̝A��x�Xw}é�I��}�������9����sݚ��'�Y{C�d��'ý�M�h޾�	�Ԟ��8����O��Y�I�T�5a�a?ِ���(<�I��>��9���mo�=;�������W�����4�z���Ì���xw�:��M�$���O�|�w̒�z��OZɌ8��d=g�N�����ԩ�jÍP�ҽ0f<	"�럽J�9y�c�V
� �w|�):�Ԭ��0'us�f�N��y�Y6��y��P:��l�����:�>o�%d����+'�f��}Z>C�4���޿b�^|����xوi$��qC�N�`jy�"ì�J�s(C�����N��Y8��x{�$�>��{��8�q�C5�V���E?{e�Յ��p˚�����t/��q�2��̜ML�$�C���O̓n�y2q+G��,:���<=�H,�C����5��;d���'߇
���l��v�@��y�9=�_��N�~�+��M��>Aa��!�N&��0�I��6�I6�f�d�C���N2u�~�H,�a�]ϝ��z��n��b�+|-����6l�=R*sPն����{�|n���
�WZ��i�r��$�&vvv(�U��(��t�u�f�Y�[+���9�/FI��u���VB�
�LWF�mc���������R�H����
�%Sl/���7_It���}����s�~�� c�'~O����&����VI��9�$�(L7g�>AI��M��'SXY&�q?j�����.�m����0<@�]���ۙy~�ߟ��|�u�}�W��6�t�3�<d���s$�q�ğ�w!6�2s��$��Y%ABd�͡Y:���P6Ì�Maa8�����$�7�h�y���;�ַ���|����x��ԃ�>d�v�s�i����8�����I��'�?>��d����~�J�$���Jɴ�����d���u�3���ݞy��۾���o�7���&�6�0հ�a�oW�M!�~��IǨy��I:�9��̛a��w��䞠�S���C�M��u'�k	YXNf�]�í���3^�^f~�]������%d���R|��N?�A��m�i��Y8��>�xB�d����LeC����:�9�{��N �5;܅Ci=Af��!Rz��߹纼�}���Ͼ�k\��~�������ԝ��%ea9��"ɷ��I��x��?P�'ڡ��M2q=�@�:����I1���'X�LO��d�
A�ߎ{�|����~��f��}��Z�*2q*7���=d��c	�7�I|�Nh>�O_?e��&�]��N2�y���'�8��X��N���3�&Шezw���8�_�^{ۯ}涼����;�p���P��2z���%a��0�a�'�u��N�hߙ%��q�Bi���Vd�z�(i'O��0�4��I�o5���g7�}�w�w�=��od�$��u����N����3G>�Ԝed5�rz�l�}d���6ɶMoY�$�&�|�z�'̝J���'��e�d����x}7�=��u���o����a�0���q4��'�� �������I����SL��y���N2��u���?$���0��d����i=k'�N%������9Ō/�`�d��7C26V�O��/E{��2�*�0S��DΖd�c'L�Y֪(^ˤN����cѻ�Q6hg�2���p������d�eIVK}RvŒÝ��d�K�5��Yug[	N��`��]�獝�m�Ow��W��q�6����ԅp���T<I8ʚa�,�>(q��,��o �2u*}��q�Xl��:�a:���d�&����:��O�Rs�d�d���y��y�{�s�f{�ݾ�����C�VO�=B��2m��f�M�S� ������J����
N2q*y�	�a̧_�'w��Y9���ݧ��Z��M����o�y�����|�����~�����IRm!��+'�8���6��N3Yq�|�S_�:��m��8�����d�d�<��$N���~w�~����������7���I��0�N�d�O�T���M�w�Ь�l���%a���a�VO�X)��N3ܸ�m'_�:��&ۻ$�+��ww��2x�����_e��s�y��4��'����A@���|퓌��<w ��'�<�qa8�2k����$�59�$�XM��� �R!�N��M��:wz�}��~������k�sy�k��ӡ�|�~e��l���v��N�m�a�2�'��0��O?2y5�'�O~Oܰ�O̟sXJ�q���T'ɴ+'R�>~����9�?~����{�|�$�iFI���k$�t��d��C���O���a�OM}�:�'�>@�]�:�d�����rC�4�]��8�wY��>�����}�>�	�n�T�eI�(��&�SS���'�����q?k��c�'P��2u$���a�Iöc&�x����M2|�����N�:Ӿs^}�������}�����M�ĝ�ka=I�wY%J�d>�IRm����'̝>���@�?yf�Y:���Wl�CS߲q��+����X+�¾��b����w?t��L��Hw��*d��9�	�>d�u��I��%J�u�7dY7��)8��'���d<5C��M2m��~�>gY<C8?k�\��;�۞���?kZ���x6�ޥ�ZZ�2�ď��.��'��֭էf6	;#mf:�f�Fs���6ǲVl�Q��i܍7(B��ֻ�1�+:��i0����x�<Z���e^p	W�U�Y[[9���3���HQ_#0�����s����|�߷�?�Y&%a��z����d�]�B��OR��y�*OY?sX~d�a�Y+�I�~�N�`~2�&�tk��o�}W����&=�~�9��v�~�c�N$�'M� m4��<�y�l*��u�T��p�&�X�q'��w��I�'u��'Y7�%t�9�7�)<}d�g4��>���������y��{�rI1�:n��|�~5��L�aĞ�y�>M2q�}�$���o���!ϩ�N%Bl�=I��2�����>d��ϒN�o]���g�w�������������'���a�ǌ�ML����6����Ou�>f�8���d�!�N��}�$����'SL��yϰ�'������U~}�k�'~�����������N2t;��	�^�zԟ�6��!�8ɤ��8�=J��T:��Mn�c'Y=�y'�q��Y����I�'���>��j�ymg�⹨�����3~�󧌟<a;���'Y7�'��$�$��3�IY4��n�mI�'P��2u=�8�m�Oڡ�I��0:��O�������������3ؿ*����߿���'t���m���:����{�8��l�י'RO]��IXm�P����B�&2q*VI�M���O��!wn�d,z���{��1�4���X>�IԝeMN{���?�v�u�����xɶO~�O_�5�|�'N'�����AC�VO��X*��������_���wg��Z>��m1��&���d�V���d��=�� �u��M�0���}�;I�'���M��O���d�O�?d�&�9���������j���w���7���Aa�`i�q4Y'Rq?�6��&ۺd��!�/0<d�'}���r�'��3�l�2~d��]��O���$�i��\i+%z��;Zy�>ق4f�	�b~��oL��V����[bU
��C���;�3_r�	�'t�u�!��*쀤M�����*j����Wݧ5�C�[����8˓G�Np���$Ø(H[�ۋ�������޼qf�����W�S��><_�'aXM��RT'�vϐ�� ��ZRq&٬)&�u?�ݲN3����N�2(i��<v��:��	�w6���W��x�򧗌��߷�J͜7�|��'~{5�u4ɨwX$���%ABg׉+'R�~�m'm�a8��{��$�?Mo!�����;}�]W�;��/Ъh��G�����'�'�a�M$�Ü�u�d��<?wuY4wX$�����a3�q�d�VO�I��o�4~��d�?YZ��b�~����;~������;�kdo��x��<�a1�a��u�sǸ~d�OP<��B����w�C�z����IԛՒ�I9��
ɷ�L?}���>��4������x?_��>��o�������Ι4ɴ<7���i��~�2LJ��o�u�XOɮw&�q!��!P�'�,��a
�ԟ����'޺��,����}���o��΄�������d۴��N$��<?Xq��������$��y�i��y����ϰ�$����N �5���'������c������z��R!��{�U���Ϲ>a?2kVJ�$���>�q52ì���זd�!�)�u�I8�s�2��'�O���!��:��2�}��������f�o�w�d.S_�>�|�Ĭ:sx�2k�}�I�M{�I_N��M>���L���u5冘q����~d�N����&��'P~���+��TZ*���ct�|�2s�_�W[d�C�S�N%d9�m��ԝ�r�6ɭ��О�=I�Y1����4�e�d��OƬ:Ì&�XbN ���  rZ���q~���|�T|�P��O�m��f�OP��p�'>��N��Y:ɷ��́�'�>|�%d�������!��C�~d�h�8�=J����߫�N��kBk忶_S���b�����jn��򘤢bxh1C%IV�Z�;�#�Q���
�f�5t�M>�U8x�{��r�!������,��Mu}�|�H�i��`m���н�/c�0�J)�{rfL�׌�n�_l��n.a��u�oko!=q�à��]�Y�m8S��s>=��J�>��lA7&���<}�%��ׁ�q�ٙ�W$�IݙA�UԋU�x�K�����D7��?<3������#�^i����C�\K������vw&��R�<<2ʲ�/��ݥ�����#���F�x��:�1m�;���̩@���֭�6c�s�]�'�9�}
ٕȌa��twXF<P��њvU_���|Ãh�,˻�9�U�r�n����9SX��6vo\ʓ2�E���M��� �G�9ϻ�qlL��vo�&�$f
��-�"k#Cv`�Dx[�<9���-�I.��A�z���q
��Y�A-��6뷮���(��.[�Lڭ��qV��:iSX훅���wV%�v��X8(T��d!�${J`�Š	�^%QinB�#}}���d�7ۘ�M�ޫ}��o3�-�uFPƲV_T&��w����^�NrQ���J�4�����9�<n����̫L���N�+]d��i�Ʈ"���v��pzMK0�K����f��F§�W7k]�_���R��z��ު�c��H%��T��L���U�}Y"�)jͨ���O3�Խul1�e0�-U�����\����p��$���:k ����J�H5��b�.:�wY�gY3k�f�U��ݾX>�n>�-VV3AsMC����F����z�7D,]9�J�ɻ�p9�͈B��G�Vl�I_/\������w�!�1{�nu���o�fe���]-f
��5�t�0��yܐ�!�SG(���R��Y^k�|��XU�S\�j���R�S�������W�����q��"�5��GiS�or�=�6�}w�:��53]�弜�N7�9����f�ms8h>�8��ՁB����3�ӈl'��g%e]�6�97q�7�^���<Z��w����������ܒ��C��Q1ƏU^ٔ=A�o���j|m�6�%ڽ���f�Z�7LZ����g�t�s	��R�k(�G�n�?7����O�.j	:y�K��ux�O�Q�}Z��B;�����)�٥��*�����a�U��R�e��Z��q ��D�tf��k�Te��+����밫,��ǅ6n��Dy����L��B�e.;*���#}#�ks<K ��L*͎�|�wM�H���[Gx0��\3��B���:f�SJ�TL�W`����^�=�k�Ǜ��!�b��%�*��1D�Mm9�ի�meF/+�����Vio���C�Pc�77�d�f$�MjbL��z���OcjO� 3�[%KiR��P��Q�H�l����
��B��0be��eYZ�Z�����b ��6P�������ҥTf�m\�-��(�J�6���iR�F�E`���e��VJ�ڍeA�Ub�J�E�B�ѣm��B�[eQ
ԬkLsmamZ��Ҡ��U(�4���ԫR�J�4F�JR��R��Z��V��*����*ѨUm�*�Kh֖��Tcmi*,��AVZQ*�����e-���je2eQ�V�H�m����kS-�U�����ZQWh��TU�����j�Z��)J%�m��j-kl-(֋Z�����J-*�Z���dm*��Z�+m)j�X6�в�eE���c[TZZ�Ej�k5\��u��	��2�+��:ڵ��}y����e�Pv����~5<iu��� ��K]�w2��u�z��`e�S7�������|ۿ<�=���������ء�� �h�y':����q'P���u�a:��y�Y6��y;��X|�Ӿ{�N�O�&k$��0?Ct>J��'�:�\�d��i[�f����ﾡ;��/��3��AI0��(u��Xn�a�N%f��
P�l�쓬9i�M�0�=�ORk����a8ϯ��sz���3߿s��|�7}앆2�=J�Ԟ��:�2q=�bI�f��O̓n�o!�N%`h��E�Y:�������©����~����]�z�S�֭����\s�N�<��U�uO���m]�Q<��|�u��J�$Q����{JQ�)^�B��I��4�xrv(�W�q�.��t��Ͻ�٪5���r�F=T�<�R<�S��~hV��(���(Η���<p�3���+���='���a�v�M�l�m�(��@�c�?|��i�d+&��{��r�K�c���}�n	s�Ƿ_H]�$�Ĕ��S2j�n���?p���[v��^/I���{YU�NpϤ;b��K��BM�ڻ�.zcQ��+�d�Kܛ�Ҫ�=&o�U]�(�L�`�u��f�-�u��or��XeE6l�X�,�!J�CIZ)��_X����S�L���x�
�'��Gݯ֪Doȃ�lUvC�CS��̯u��2�����7�ˠ�FίI��a{H�Ҁ4;��9s��X*)n���c�XA���43(㳥G�������%�s�����&���Z���sʸ��ϕ8�yU2��b�M�x/k.����{���I~��^}K��+~�X�{a���B�~|�>l����7oA�;qaI߭�;Ι}���u�ǭק�c
{ݻꓹrة�+Bu��|v�^T�W���X���Ӌ�G�t�T�^�OS���t�*��w�7w>��Ӻ�P���,Z�mW��6T`���ϏxZ�7�gk�֧�7�3�$�m���{Ȓ��!�:���}��ɔ�/�[E�N�Ӂm>�����u��=e&��'��I>���[���46�}z5�=m���R���Τ�^ۣc�e�~z���u<��?p�蟩=~78\�k�F��a�f\�am��w��oshlZ��h�M��N)�����Jz�`��\���E1�GW`�ۧ�⹋���t��F�|:v�u�ϳb��b��[���� �����w����[��V��;��b�bt��ԋv�뭠�l���t�+�mnl	 kd��.3{�|�����8�X�`ر>���l!nWK۰A�c��k#b��%w�ݾq�����{���pd�;���w9�[�W�$Q��Q~������B�w��o�s��K��7��E��"�)�)�F�Y��{�-<��}[>�(�F4]Q��[۬��㳩�r���g�Ur�#�P�33�7���)A&*<��-���V��L|9'=��KR!a�s��y�	ʨ|=�vĒ�O9�&XѱQ�֟��Ql��-ܸ��{�]���"��k��R�W�歮��mC���.�~����yM�Ob��|�ù���>��N6��=�ѮOҀn��xnTX�뷞�P־����Y�߫sS��ױ>����b{;�d�3�o�"0m��)s73��W3��s�?M�>N�TW������]������۾�ifw�\ޥ�Zԯ=�{t?���t�����ϥ��>�k(+w�~ޔSӦ�M���2y|l+����ic�x$<��a�<�y�>��cJ�߷��C[����Q����[�}d��o�뒡7sA�α�By����1�K����3� �ff���tn�ӵ�ި|vĔ���uSN�Ԗ:4�Jj��(��cFV�.�r�"��1](���\��+��M���_}��}]io�L{5�?}��.tϩ���ߵ�L�ܢ�V�c������U-�e�x'7ݭ��&��uH�*�N�N{�OԞ���ۡ�V��b�u�~E��t��:9\���aW�I��R�N��͋�7�p�Z5���b�M���;�X��+�.�G���{�6�O{.��c �w3֫w%t����̣��[gM=���6O3���/����(c0�V[Z���bP���Sս���Mڮ���(��AuG�#On��qٶN�W��g��3��go<��Y�^ʒ-�����������Y{����M�x��^g�gGo��e�����_�I65;��q�]%�"�w�H�y}����^-z%���i��T���ꦭ��䰻�ٵy͎kۼ���'�S��Ѻ}׹�Y���1�p��ʎ��'Qv�ﲤ9"�#��7�����7{v�rD�:|֑�˼����]�S��w���c��g��u�G4:�WPf�X�}Y��[�tN��1[�=T�2��������혀��/U��D�cN���u�e����"�t@t���ɼ�~���ꪜw�l����;�5��ו/G;���9~�u�Vw�S�G=C�/b����it���U��|�c{��[�c_vy*/b�Mvܝ[��7H�ZΪ�����ӏ=����U乹��#���?n�W��>q+ֳ�H������r�.�S��E�{����;*d���w���v_y[��t����j����{�z���*���Y� ��q;�f��BI3g�Yg�bokѓR��fV�Q(�]:�2�2*�F����N�����y�W�g����Z�*+u{Nؼ�(�!a�o#������cΤίJ�=&'R�n�BL���wmXۀgQ�gYぃ��a�ӳ���j�]r����Jw��f�zh�ow;����ƶ`�b�1�c�F���j��w����X:�-풺����J��zx��sW�)^)�ST݊[���������g���~�LY��_�ѫ�ʥ%}�l�{L�>xrso����|�f�@x���4>�? @�	��IϝH�]m�ׄ�"w��oZ�����q{g�۹���4��XV�p!���V<|m���t����ˏ�_}UUT�Wv	��{�:����϶F��?n��m{����R%QS��'�ۖ�ӵ�=�n�0/v�׻y�Z�����~ȏ�x�k��[/c;s�}ѵ�4��Y6��	�ḏk�o���p䪽���#�-�L���}m'�c~���^ё���u�2�/s�W�����ḽ�.�(T��8�37���<���W���:�p��5�NyW�\~|��N��O��6}�[�'7ݱ�o��D�d�oӂ�<�eF=���`����/!QEyWw���-����~�+�-���z�O�J��;�1'��&�~Z��r�u�	.o��c�r�v�Y�VV����t�*��w�<��U�;ڽ�U+}l���M�C��[Gڕ�jQ���Vv�3S���S8���j5 )�o����(��vO*6h/�}q|_�:5{N�u6c~������̇]v��(V��@�dV���,��Еn��ës�Df)d�VP:���/�B!����-���Qu�oA˪.ft.�Gdn���8[�#\�ևܘ�������U�ࡌ�-u�p�Ckl�/�������-o+��(�t󿪾�꯾�<{Z���������<��0�գ_�[_�}W+�s`*�-����h�^o'2�}|#��d�7��̞;���>86�lj�碧��bp�>�Yy�ϥ{���>�&^A=3y�mP�vd���B���q�u�u��H�/y�g�QyU����j���������}���vu�ü�&�T:m��ܾ�3z�����ʍs��������������m�U�I<�q�9�=��6��ζ2O�p�g�Z�{�?}Kx���5��ǷP�=%oW��������ku؁��ľ�8hG�ɮ�U��F����]���|��������3L��σ�JAީ'��'�N�A�^�_yi�n�টrޒYY��,y���7�c�/����^�j� ��J�dMs8�Ȏf����px��e��Z��~���=飵�T�:��W�p��W��L�p���g;sʠ������F$�v�8�b��ib�:ֲL1�������-Gf^oM�Y�{�䭍���l0�(»'��"������Ѻ�Z�ヽ0�z����خ���sNҼ��*�|3�v��]&
�=����U�}�}��B=�Nw˃�յ����X����?nju��gl�4ʬ��#^q+�*B:��c9׮R�*(�W��{*�y/��_bwK�:���u=^��k9M��
{�@���W��6����m%yֽ�r��-��[F>���zQ�'~ќ���	��ɼ���;}Rz�A��B�gôk�w�\��h�͢�g�MU��lO7��L�c�W�{��46�[�և�÷�a�F,8��wU��b}�R�J��tbs�[+ګf7���[Kۋ ^�����((��}n�|y����IJv��M���¡�v=��]��^{r�ҙ�����k�\�0��{f�{�k({4Q���s1���-g8/'��Fz2�8;�jyl�͓��P�)��7��v�x�����sH����'�R��T݊U�@;��C��C�l��;����-Ǘ��_j��k�<�+�8K�O%��*~Bbԟ=�ΉFW���H��d�~���3}$B�H�Z�p*���z�J��g�X��+��zVqΘ��q���]�
;��nM]&tS���'o�7�Z4K�r�|_:K/h)Bj;�����}Ue,���-���	k�8��E��\��O��pʢ�_��U�i�l{�۽���W`w�&<���L�(��B�x	&xO9��N!_b�yn�V�e{7d�>�|ݗ��Ǣ%^�E�9-8�)�(ǳ��k�7��{���]ļ���T8:k=�ռ~Q��x^s�Od��{9����y�۫j�8�;��[�~��k��}�|w��+Ǔ/z�/w��w?i�5 -���P����<����[<�~�� �n't�T�Z�Z��{�oӞ�3�u�m�O/j�-Ϟ�'���7_-���;��5Y�UhT�3{;���^�p;� ��{�(�d��nX��~񴕎�5�vh���~^BOP�/�������u��2���w���z,��kr'N�i� Ʀc����`�,��V���Φ��R������P�{ΕY	˱^!�tVU7
���w|P���Ӵ�i���Z����O����{yʥ-֯"�~̧ә�{w�\B}�+a{�\��t��Y���N����xk_+�P�A�'\�۔��*��!��{6s�p�WO��,�ۛ���������9I<�}�W��U�/���׫i���,mxy�����k�k�
��Og�Ckz�_0��;��݀���]h�%�3�+�G�TN���n�ۥj���y�۱��=+eKSy�)��N=[<9;y��Y���c�]][��	�_���68=�5�~����_9�/>R<��nۦ��oE�l7�ߐd���k{\���U�W�_�vmt\�����I�U)���5�u<͐��6��6�_��A�
�_�s¡N�O��Jzu|c۩���Z�/j�<s&�K�׺����^��:���e�+�:���x^���!�ʵ��3֧��������~���U�����5�=ٺw�o��Qj�YI��z���W�O�i��l��(ǝ����z�_ǖ*���k�O%��w���k7|�X�+�����P����O=Q�_�^�����z��WB;\�ߜ��ݺ�Y��+�uۗ�w!��@�W@��^�E�
N+\�:�R77�Ͳ����T
�he��[�hź��7%�f-��BR�O�Uv{u�����C�D���	��W����I�R\>��o;�L�wm�K	{wODl3x�\�y#%�1%��.���a�N�S�h2��<�$�;��1v3M���+vj45���Y��Vf�)�FZ��G�|lfO(�N�.���Of��b�="����U���欂^��Ĭ�G��V��QWk���æ�U�'m��|�tZ�k�,�z����2��V�j 1�T�+��eLіjeb7�4=o�$GM�G��+(ūV���Eۺ&��
�u��H�C
�D��s����c+Z3�,����4���Ԑ	\�c*3b7m9�G�����f�]v���xm
s�G�aH�ؽ��.|��ZqVB�4�/h�Ù�w��}2T���	�x�uEa��_LV�er�`y��֜b�e;@��v{���U����mb������46c�d��[HK;	�=�L���f*jpjus30�c�pV���0�/SȖL��j� ��L�jpi�!�x:	��I;2	ͫ�VXkX7�X���@
��o*�ƞUv��\�ok&��ĺh(ufu��3��r��`*0�fG���_>����ʈ?���+���Er�Όp���l���*azfuu�|EEt��>����IKTw�v��VQQ��U�ǂ��As�-��z$�����ٓ����)�S��j6���f�^����7A��bj�{����C�qRU�;,Y��S=�N�L=����o4*A��_q�� + ��k7P|��n�G��-�,۠d� �E��n�u���b���>\I��)hS����mr�yk[ኵ�]-|�g6��x�;E�1x\��o�ݧ�9��X��/m�rFJ)������a��=���.\�)G[Sܪ��,Z��;�3�_!ڴ7�"��F�EV�����s���,4FX�����q�E1�n�u��'q�&vs/��X�]gӕ ?\f)#q&	�Ͷ4�p��ٹ�[je�D�8�Ϸ��J���4���C(c�X�'X� ˆ�3�A�0�OVt-a<\Ͳ{9M�Г,�;���X�t�h�o{�i�<p���l�\��ͷ�
��p܃	nI��I�d�S�W_�_����T@�Wu����»[6��s.�̘�&^&��9�$�l�^Q짤~�Va���ʕ�ǧ�5e�z�#�_�1V]X�ƲK	�p@���՛��W�n��#�����heCR[|�g�S8���\O����x�6ЫU����P�0r�t,Xp�y�0^�+�묻�t��1�-yb��耪������5`�V6<y;�tn;���Uv'(�F�V��[�F�nX(�:�Oַ�-^<���x�6(9W|x���c�Q�5vJ��4����2������Z�P��%VTV���h�R�[U�����U�Q�Z���F4Z�ҩLI�Z�*��(�-�¶ҋ[Y*j֪Yb�mDV,X�V�h*�PQh�H�F�m+F�ڑZ2��+j��h�U��)F�U��J���֊�-����J�X[Dfe0H�˖�R�(�[h����F[UR���F�TR1�V��EX�PE��X�E���dX�Z�jZ�QV1��i[J�)TeU`�h�T���X����"6¨�iiJ%U���-�QJ�DER�Q[eim�6�H��V*
�R6QR,DZ�PJťJ��*F���ƶb)V1KTlR,J4+"%em(�%j���Q�iEF*�������1���m�X�Җ�X����ZYX�ҕm* ֪�E��b8�DT�*���KJ+ƫ��մ)@J�V���fX�"���D�h�m��V([Kkm[j��֊�QF5�e�l��Ŷ�"�m���J���ѕU�eh�A"+TB�j���b��U����S\�Q���-�D-3.%�2��i�7/w���*D���C�<���)�{�'|6t�핝'=�8R��ԫ�({� ;ӱ�D/��PNj��y�m�2�k�]��UW�}T�c]�羓	��ܵg�?"�ן����=�*��nT��~�
�:�� Ɓ��'=PLx�����<�u�VV��^z�F����@ĤW���O\t�Ϣu�/W�ܑ����GK��pejq;�{�{��9�Y��s6RO���k�����@�G{(���]�6�7�s�Θ�lǳk���Ϥ��,j3���&��ud	{]�f�j:U뾀ǹ{�a�8I�\#&J�7���Oi�ͮۙ��u����w<p��%�����&�-^��{�V����s}[*)��9��%=U�*v{���{�wvQm<|�Z|�/'qH���o�0=3*ߡ5W�_>y��ü�o��k�� =��N�u+k#Ӳ�L8�3��lc��������\��ҳL��X<<�o�x5���r�]Ӻ}b����ӑz��[ ~����Y�+�;BS�xp_21��1�K��N�-��}IN]�#{�3t����� �w�ԪI�V����hN���c�M�>��V��s���b��M�z��i�=��l���y�){{�:�>V���kCZ�Lü�T
;dL��+t"��֞�����U}����Tu���x_�M~�n-��<�����8ml���U�WҲn,ÂZw{���N�{+��򄶾�w�UI5Eq|��|�����r�)]�RY��'<�W�.����E�s�ӉҐ?*�^����D鮢H����^0��߻���_���ꮮ��8�����MK�4'd9@0,�A֦�֏'��n޽�V{�y��#kz�n�^�O�[��4Ju�[Y���%��W6�8�~�8G/m�y�~�<>F���;�}h٣$Z��5s���$g�ڮֵ+��̡�)ޥ�}������yC/��&���m��O����d쯦I�	T�>{��-p��[��C7to�&�k�*��m/�����S�q��U#{ޙ�P5�5��b7��Qv<�����U\�oI��u6�>���3�R͓5�/ L�Df#�H1�o�mp�H+�#P:�:����r��>G]_�ᣬ{�������f��]Sv��������\�JOo��6dP�gOZ]d��x�!bn'��8�nR��҇����X�	���ol��e.��c�I��bN�z^���U}��T����o�gA���*k�:�\�Ty���ޕ.O~�pN^s�Q�Oi�����ڼ�æg��Fq��w�{^����=].�ȰY����w��#�҅�.|�L����0+w���oEF�]R滦e |F,�RՓ�i��wy�!�\��{x�%�5Mإ���j�S���f��ȹ\(����9��6�Ϲ�<1g`�{*��r�O(��@�c�{k޹��]-k�sO���3-��8m�����}"�>�/���I=�[�Z�{�o�&{ݼ��<���o�����z"^�E�9��} �R���zvc�e��{���:AƯ"���}q��y*����oB.��4Z��~vUǮ��ꩽa�p�����	β�ʏ9'=�U2��vZ
�g���9���5��$�z2�?_��vj�<���oj��Hl�6���It��@�	���6E�B�h���5�z�t=��)����5�X����AF��*}�-<
b쾈�7F�8rkZ\0�2�s��nqg����"����[@��5���������}�����8T�������Y'�y{\����3���^��^�&f��ꓹr۬���^V�q�?4%�X������[�PX� ��OWg���o�^�J����m{�z�@�����(#���}Q��p*�qS����}�檣���ڕ��72<��/P��C�'a�nL�g��9��Y��7�.�"r��d��WRO��T��,m�r��ʉ֮u���u&0�<����o�mMm�꺞����]^o�q�t+�~�|N���o7�5C�w�<�Z�O{]KSy����=[<9;j���o�g^���iI1i�V���՛����Og����5�j�H��NNߩ�[OS��:��3շ�\(�M�]�b|S�i����ܪ󰵋[^�_���"�q��Ƕ��gk�Z��ףB1��k��B�Ի��Jzu|c�W��xU��i2�����7�iW���]�urq���)mVv�s��Qc��������SՔ�m:%:��yh�$`���S2ђ4f��|���<{���з$�Io����;l�H��v�']VT=c`y�n�{6���I��� ]��;O�UW�U|s�M�OwZ�:���_5Q�
����Yz�#�p��"�������I_o�g��s)���c�JO[�j� w�2��#����zWo�xv@��Fs�f��J�d\�o�u x61�j�P]�����hgft잾����rN3}Nyv}�k�;�r���{1�ō9��2��l��:���/�yJ���1���tqnc�r���nd{�	C6^�] ���W%_Ly�M��n�L6�WR��6�sD���m���`�j�U��mVD�á22��D�{��Q˱Y����B^�G�<����ż�!�4<�����"ל4=����ְ�J�W�AӃq��^�KW풂�%l��5�$��r�7��F������bCASPT�"�1�&��~�1�>�=��eW�1Jq���*�{��샽��#����Sl���"���'<�������48�V%z�S~��a��1CC��l�J��)2��K<o:�LZ���iҼ��`��=�Ӭ|SP��zr�U߇��7�,�jԷ��+	�L��G���~���ו��U�;4�:��
VD3��Y �e.{ϒ�&>�}J)��;	�{3T������D;G>W�^��qt����U���Y��6l./���}_UU}[*옹I��oW�lo�dj��V5�b���S�jx�81�A����9iv�2��-vM����"�"R�`�r��cH#ʶ�c�b��}�,;��DP2�p�g%�U�_^���D�z�b�C����S�s�,�\���}+
��w�ywUN�v���^̐nΙ]�Z}b��>��F�`�ץđط>o�҉C�ݹ'���l�s��������>�46��r�fE�F�=P�He�B��$t1jT��c.��Ũ�G��Ng�َY�3�s*§/!��c>�[Y�Se?"�ڎ���{5��.�y��o�Bk^���v�˯k���JD�X�q.�<}*�@hS�E(qv�0������y�� �S.��݀�ν̋}u���oD�r�N*��/��6_R�k.](�;v��i���d��tX<�go�@^tyT����~��z�_L�~ߺx����|���Ɣ`�}:�0R�|����=]��f�А�W�*Ы
�p�`ϫ٪	Zq�"�ޫ�]�Z��(l��+���V���0{��H�R�ϴ&z>�ĭ�,�uQ}��ٴ�	�479�:���j=J�����?-9}��9uwC�E�i�O���^�����]&�
��K>=��nm`6T���6�b��$�E��E����꯫���z��v���4� �-_���F��.�lxr�V�ØS=�7���Gj]yވN���tg��S������q13�á����A[�a߼o�c/�f=|8���p�'�Rp�$Π���±��W�����ֹ�qq�r�B12�#N�,�mnL^���N���p�*�q�`{\$����U_3��ġ�{��������qU�;�G��ټm��4�]І�&�Q��2��yJ$U�!#a���,�$�V(s2��-d��gc�9�U{���a��/��G�k����KR�IȦ7��V�c>���<��;��;0^gV=�{\�:������<���"����E]Ni��J��=)�<��O.em�O8���E�A�LU������>+��DU� ��|h�e�Å�=���˛01ئ�c}ON��(gXS�hu���9K,zz5U2��!�b�w1��tڙ�:��J�Ԙ#���<+<�U|1�0�J�:���R5�bF&$�l�oM�#��z����@��8�yf��b��+�>L��ǿ=&����e2E�هiv1N�U��B�(==�hY[}�<sԨ�&;��]�C/��������/�֊�cݰ��r�>��YD���ϣ��G���X�h<f�8`��f�)������/.�O������p��Fً��D�B����^3��7�'�����n�[^]�"Os�����^��T�6_�u�V�#��B|tLϛ�	�q}�{�S�ܱ�����>�-=o�����k 6X2Bo-T쳆��U���g��+O�o�=�+ȸp�ƙY(m��g�v0Jg�ǆ�U�J'��`�K>���h���{~o���j�+��gK=�#���^��&�i��z��^�Y�R�oNg1�"W����}c�2Ҧ����[=>�����p,iJ^w¥ejT�Ϛ���2'���<�ˇ{Eڲ+Z�1ꋵ�tw��:)���x�Y��B2��@�&5T�1=>����|���~�H�e�V_�3e��KK�m�O���Pc�D���J���V%WN��gy�����������* �\|���\>�{��u�>J�,2q�۷=V�ʂ7�mzM���r̊�R�;��W�s�D<�$C��ω�M+x����5
9����3�c�;����ik�k¯��e62�ᄠ��X�����y�{λw�ﷸ��R�5�7�Z�~QlEz!B���L��<�#�sz�םኳ�"ܼb��J9��ș��AE]��I�刞����ľk��nW rB(\�s���������x��ҽʗ��3�8 ���Y9�X�Q�۾���#�g�%��j=��'e���y�.�뾾��bxߖ�'��S���.65LC�7�����S��CiW�M�k���ӳ�c�~�hJ]f��������T4�<"gZ�Vq�g�:�^�x��(��PvdK|�G���>�WN+#+���,���Pr��@_���/���<w�ɪ�z=*Lz�yN�Y�`��{�"0��$��/O���S~���\%�;��Wl�����z�{��2|{O��2} ��d���l�>�%��-#ڳ��N�;d-�E�o3����ٔ��Ϸ�U�� g�ȸ
�JsF�x�0���2��R�tV����V��>�gE��r�}��f����r�Of1S;�V�!n�
�]��=	���=|)����xoG��e��Ԡ���	C>�z)t��q��N}6��aw~�o:���f�c5������ޞ|&Z�ke��с���-��W�h��v*��q!^���/�)�)���� M�V��+���w��08٥�V�*"Yٰ\~��ha�;yCzZ�[���&z�9;ĭqp=ˡ:��M�("�.��I�gw�b�-ݘ�M�)�%���u֩�d�z�.�GxI�#�;�һ�UW�UWy�;���y;[�lq����V�����"�p�8x��I3����"��ur|������Ox�3��k�"�׵=pnZD`_:7
��i}G���Ƃ�9��v�6��N�����bw�)�;��2m��ɪw��Q���m�_G��]x��UW{rs�B�Cb�Q+�b�s����b���o!y��U,����2w����E��j��`*��m�3��J�����#1z�z5B!����È��.�K���{fZ������^H���dwÃ�n�T�ê:�a�Gc�b�0>�p:�B���y�3�����^Z�Zj# =�Hн<L��򮭈��d�X���D�fi�ʱN\ƽ^���wp˩&i�t���F� X#X�+��^kb���
q(x�yFy�/6c���7^����l���l��fW`w��!ZF(���b��`
����ŭ������Z�NOo�sf1���o9P�j�Δ�>�c+����5TĄ��6������bFi���o�+�����S�d���ڗ�8�p�"�7���{slǽ����T�W:&1{ݴӒ��>�y�����d{�fKF�^>��q�E�	0�����'��O{iY�"o0d����=+Q/j@�����7+Ь��B�w�G�8H0�%��_�����&;��<��m��Gf�'j�]�؍C��ס��L�:{B_[7c����l#v��H+"V�n%+d��ONgˊ5�o7{�ͫq[e�;[=���=��H"��qyg�h�VL���+o�c��p\�d�k7t")m� >a��<6��}��X�B/T'}m��"�1�٤�8D��ϳ1u٩�GV�SV�p�kp������m�k��+%���	�d��ٯ�>��3��zlZ��/5
d�Y����h�{�l<(�I�^p����Vox}�q��v���R�T6���$`+�Ί���F�q.\�GۏB�����#g�sZ�J�ʘ�n����`���aV�m%��$��*��4�ɛ��'_gQ�ݧ�nL�O�|{z� �B���@T��7��isG��d%
^6�V�����1�ps� �����)=�v�3V��8@!Ȋ��Nn���}�����Gb��,:�e�Ų���]	�QaPƷ�Z�C�Z��ǽK�� >;J��ѷ��~��s����B۔�E|q��L}~��5X+$N���B}~4YW���#�v%��!^��|ri����h��Ce�pwL7ܵ��9h��n��փ��ʏ��c�����߰,˸<�=FNr{�� 	<�žh�^!=�s�E��7��MD�y'��Z
@62���Tk���%�/;w��[}ҍ�o,��l��[�-<M�<N!m��{����uy���ͫO�9̍�0\\AƯO=�g%�:�f,���R�m᣷"�Dm�{��	��ޟ=5ӝ�씍0m�����]%b���y]�Β7q�x�
	�l߷i[X����o&)٧��
�p}��{%!y]a�V��s�]�\w�)�s�ʴ���M�ʗ)���]�h��yT�p�:�4i6޺/���wA�ƴ�S9���.�"���y5�����X��^X2�9��1�we�BmY�k$O���<��k{�P�5��5%v4c*�H��g���k�)С�G`�8�Ց ���̫L�G�:�¥Ӱ�,n�1D�1��PZ���kzҧ>�}�Eǘ�5�6���j.ú�N-����O��;�5 �h��n�>鲹���ξcT$1���:�n/�M��ŏ�r���~��ɔ���Lh�����go�����7d�bf�]-5o���ӄ���!�B�	8s������'f�w�-�z���r,��f���9�wf񐟮�Ҳ�}0����Q|�ڵ�������ג}JA��w��ȩ��8����\$s���o������eJ��J�h��Z����ōYlF�
���J4�h��h�kb�ب��keE����31R�F�ecceZ�Z�X�VܹQF
"�Q�ʊ�B��h��B�im��.8"孭�V"��DEKj�2ىUE����XP�(�+E�6ڭ��Eb��+kQ�U���ADED���������h���ER��-�F)�*��*����,b"���",*�b�%b+Qb��X�P��+QUڌ�Z�VE
�B��(%l�(�RR�jV�-����R�Ĺj"��TQ*�ѵ��QPJ�f[qb(�F�UDT�TY�2�%��am��T�h[kTA���)U
��Ԫ1TkH��1�LnKE����P`��`bcEq���,[J1�mV�lm�UiPQ�QJ"2�QQm�#iU���e���ZR��(����E����U���*٘)-(��iE�ܸ���pDq�"��kD`�Z�Z�,��,A`(�TV,b�3�EPZ�Lj�e�ƨ�1D*#amX"*"F"	���*��)*PVE��3.8�8�EQL�[h�L��w�����;�� ���b<�Z�v�O���:N	����y���V��[:���s��t�V^��z{_�U}_}�I�cQ���~�?�+�p藔un	����d�rثNf:�Ie�s.ըs\��ӯ��f#�E��I`C��+ЭG�����ƶ��`Mr���ԫ��`�b�4�<}��H1��}����p}�ҵxi��R�Ɋ5k���r�G���NK6s��o<Z�Q�!֡�Yw~~�wu�ܶ;
��uץe�7�#,�Kΰ@��ь�Z~U��OL�س8��0m1�7�ʗ(vN�jckb�yմ0��/ǫ���Z"�b��L�[!'ӫ���owzǈ�~�Z<��4������A[�m$x�+��6�����T��Յ�evN��թQ%�A�C�V3�*��SQA����,1���+}��d���;=��l�;݋	X�X�� m��� :����;�u��bc��g�]u-�%˹��<<3�r`�a,KB�����$U�!#>��S�+����Wy��n>���r�{*��ίB�^]��'h��t7Ym�U����\|7k�S�3Z��K�Ҳ���u�E�z��b(�*>�K�;��Q����s	��|o_M�y/M��k����bX�=�j���umiƖF����oI�C�c;6��s�1s�����	H�.�%��-'��ۀ��n�;ȝf8R�zջ��:���!Ϸe���}_U}CW%��\ߺ��K���>fp�GӪϭC�^�~G��0t���,0�Ƈ�[�@_X�}��/{�XC۾}��=n{F*�K�9���R'�{"c2�  S�u� �	P�&$��w?z�yϐc�xW'�=8z����)�:��/�K�wԢ�DT`zly���
?d]������7�(jL�m���}Y劫���T�������+T����ܩ~�ə������)���G�P=!���&j.�j/�m.��0�w2��Q�z�4i9-y�7���0_4*�w�F��l�h�K�E��u���φ��Z�4;��=������X3`��� HX2BuO-T�� �q�V;�綊4��V�Ƶ�C��׾K&�Ļ��Ϧ^�,h��jP!=�f�� ����b����mq����_^$��>�sqƻ��Wf�Z[&��3��֫�C�BC�=���u1�.�h��E�:\�����V��ī��o�%��V4��+5*p�53+|d,)��]�f�=���,��GX�]o:9�s�M|��&�IG2M��cUh��L�{�微�<�[����|/:P�g�Q9U�R�ǡ�^��u�ݘ���(��d:���w���PC�=�WR@��[��+աǬ�̛~�)"�uv���cټ����}_}sh��dY�S�Ὺ�aU�-:&�>\�9���ȍ�I�\g8�:�(�ù�Ox�U�y�Y�X`�P�u�k�aW��)M����>��D��fX#M�4�Vˬ͘N���`rs���K:=Z8hX5��b:�Yқ�ў!���7��SZ���=O�=~k���*�]''����=2�}Q"F��_��z�{A�"~��杽��b��|�uҖ��`�����OoJB?,�^�-���C�B��������R�R^�͜����P���3�cBy䩊��|�ީ�xtޫ�Q�)��X�ٴݝ��'�c͗�ш�u�$�#;J��������4�utv'�x;4)���e�Q�h�s�l㺳��C�=Y��t�<D_��J�wX��@����Y����0k׎�h�Y�Y8��$���X�%�J*���$��k�}E�����z�M0����rY��>�ĺ>d����dD\0<��H-��V6G�(u�r׀k�d�9)��V���k-L�LY�]��v���X����">�n�u���j��=��x�7�.�A��iM�s���+y(��u���Jkݾ��ђ�\��v�ˍ��L�m.���g�ͦ{�a�5�/q}���׬/��5Ǖ��[�i�+�C����}{6�������=�zg>��{*�<��gE/kUe�܂�AUH-�9�h�TP�W�#]�M��=y�`9K��d�ǹ�֚�_J||\�Ec9��qW��R�{'�s����hF{��c�ۼ�����$ �X.�nQ�<�}�g�2	�w����]%e(�` {� �K�5��0�%����v�fZ�k��i]R0zyp�p>"UǢB=�b���������菖�C�+b�M�n�U=}�&r�9��%BF�C�C�7�U6�C.λ�[�䡊X��^O;[��E3��*z�	��u�����F�qN$m���Ե[�^t�,�g����:�;ڶ!��LEM)�S���*kOOo�ݐmҌ������Ś��u��*s���O��z�v�V�4�#�4�Q*�b�L�a�5C�<�/�s�|xկ\�ըNM�������m��֢>C��;�����6Pc!�}����#숯
���t�vs*3䧫k�n�M��r$x�.��_�×E��ƐyV�u�K��1�0����#\����2���nQc\p��zB�p�9;���/��\OY
���M�2�P�����ʖd�I{h޽�zU���
�Mq�h�p��W[f�r��ݙԻ�z�yɞEH��쨉S�)]3�K�k:�7�_ku���se�m���������	���[m�G���E}�������uœ��[V[&*Ɲӳ�fR�>�s����:����n#��V�o:8o꒫O�����G48�<��p��\�M#�>�1t���;�Y��L���qV���A�ã�	
�1E�����������ԕ�����%���6W���;<s9̫
������I���Ck>0A�i	U^y3w��\.vߵ�ɂ��b�nGBn86�P���JD��������u~�|�(�#�/;]��!���to���gf�*C�a���K��;:둃+z+%V�J�'��u�{L7��w���j�^.�[���X�@^iݦ8'-���o\�&�y.��KW�mŹ�n�:Vo`�S V�^���W�$��ք'��`����XS>���'~53g��w�d�;ų>ʹf�g��CFS������O��|!�a�e�;5�<u����LǙ�r�׌j�U��JPʡ�a������>�NM�
�LZ7O�����51OY�45�X�����IVJ�B�ü^������d�o�]�����.
.�W�)����.�w�V�a�(���u䯉/�u�.
s��%�]�)۴�.;�t<�C]!�:u0wo����W�&&m1�%�B�ɫ;_� �/�d��`G���nyu7��pa��tgXf�)©����'��o�Rӗ��hє�V�ێ��+e��HM��w�C�]�	�(���U�q����5�d^�� �Uu=�z�Dw����*�9��53�n��v���dTH<�ڐ��[*�x�h��^�nK�֟.�۸��Y�neug�?O+�yF�p�%��;Ϭ�e�`/E:�xr6>�v�ͼ�i�_��V�Y79�=Y9��+g���
�PwN�*��=(�|�p���8�zs�N{�ȱ�Vښ}FyA�~1V�T�?yVH���}�1�U1������I��������n�K��)��F�f�4*��Z3�J֧���1�Z��r�z��P��8���'n��<=�n�Z�ɬ�-�����֥k^��9P��Y励= ����_�iZ��������&&.�f-�\d��ccG�S�H~�����0A�>s� ��Gfꢦ"�f��2�����
K>-]��yXU�g���n�L!~V�3��I��my۷�E)c���S��Uk�1����o]�>��܋U�b�
���e��$)2�:�Q8U��;���
�yY�A�,�T�����y�D�|���غ�0M«L`��<��r�b�����C+s��pl����\�/hkx�򪪪�/t+˦����ͫT�ZwQ���2F4n�w���w�QRr�XW�������9�ky{�G��yJ�
�pgd�F�V{���"-[^�������v�ո��Y���'��%�V��S&��3�������Qо{'=51ݿEZ8K�`�W��S��^ɰ�%f5p�sJߪ�%d�1�R�V��YZ�8q��Z$,��.��f��̈t`�w�{��qP7J�ץ%c��\�S�	�/x�W�G��؍_L�7��W��>m�Oi����PHw�g��*�+�[*ϑ�������C�_��^ͭx�\��v�.zB_';���!<���ז��]0��Z�u�m$K���S9�s}��K(X��%{�����h����}*��WO"}!�G������D{*�Z�9g�o���EL-�u��猝1=ճ �Ud�c��_�Ğ:/�o�؆������R���0�B�?�MU�Ǥ3��M{�}^S�Ox+keЂ�R"�̤��#.��wp��3�i��1oa}�iO��W��/c�{m�[h���gc�z�;pv�x��Z����3��{5�.���N�?u>'��f������ދ�����3Y�S��Y3��q�� D�]��VN�x���磌�"�>]{A�� ]�ü�/cQ/7�r@���D�����P*�:��^2�Iwq�o|���+�#V"w0��*駈оvC%[�ϒ��޺��WY�S�\����˽��f�g���[��Xz8Da	uy$qz���z7��,/�*�(%�gN"K���4ħ,���lV&��� *�[�2�b�����b{C�Ud��z�`�8��y���x�8i{5c;�E.�zeYOr2�P��
����o��X��^�֔����<�A��~�5����ag�3�����ފ��})U���t3�<X�Oh�n�;"�o��o��.!����*��¼/���:��x{b�e��R})V�R�������k�ޝ[���1��*�a����Y��டQ�[Mr��WP�|D���C�cy�F�û�]��f���d\��(L�n��tɜ�Ni�T9Ug�%E�񺤤/�Ã&��w�X����Wh���[���L��.��?�lS��z����#`�;gQ��Z~�Ҟ��E.��!�;6�&?V�qo.��v�`V���qp.R�t7�q���vp���⧴��G�f����Sl�F�9��N���T}[�oD�Z�� �u�O�J��;����<�3������X���!׶\���Rz�nГ�ݱ�W�R�;��IwxIDUe���J�02�SSJq���*����샽W����";��E�s'7CMi乮�1���Q/�b��R*fq�����5�W����nQ^�o"�Y�-�4g΋�ĵ+OEM�2����|�>��C4��X�VG��#D��g��f���W��r���
Z�*즑�#����h16��[T�k��<�/TXM٧��a�W�+��]�Ou`R��g��N�}���.��P�<����>JR1���'��.�0�SѴ�xO��<fۙ�>����3����σ�\�P�G8/�Gx��B�O��Wl���e͘/N����]��7��~�3<;�s�|$+H�QA�S*\��m�r��[���/t�g�u��*|U{E�s���X�/!�R����T0A�j���*��ٜ�l<�xO��Ȧ+�ʲ��x���}f��U���*�IЫ��4�t<|����{�N�S����Ġ��>3:���#��^�I�|�eM�N{pb��{֞1�U�uxy�e���b.�;bz�F�\a�[���5�M����XRZ�u��Wv�~�w|���S�O��\&ҽ�K�o�cRq�����W�_�1�n5���ܩ����9ysU����{M�xBԥ]� �KБ����%���L��}�٩s���:�[C�����ħ%kFW���Jɼ@3K���ag�a`Ʌ a�;�9�����+�^'L�� �O'��;�&̯JkB�U`LY�y��n���K��3��ݽ1e��P����u���b�3�׶���g��6'��>�v[���%h;FRj��m������=�-���
��RR���q11�0�b��OB2yٻA���g��-��{v,>�\S6����8�@��C��g�T��6�|O�L���AFf;��+|�tSU穑c;��+°������,�Ii�2l{C��
�OqW��u��z���W~j�`>�6�=�����U����s�-LtEh������$�J�eX���umw�;'0V(.2g��6�0��j�E������r)�`�|�?ggʝ�MX�pIO�A@l9��*���؀�&�2��'<�^�E筑��lФ8VP���Vxa��ax���h2'�+)=;�=c�<�[�}�b����!�?�&3&  ���+Ϣ�D�i�V���紴?`ޠ��5�l �\��4�Y�(L��+rk��8�N�ǉ5��+�o"�SyXӽv�Q0A��˳��q�W�R̜�8�Sx(:�w`oP�2��,+[�T����$�t�fc[ݒ�j$���ML9/��W�q���O���v��7P�+� %N�ݙV���Ff�m�Zm�^��왽L���[c)��j�#�Z����������-73����*X�v,�2���dbM��0杝y�1`\G|'����[k�����e�-;;F�i3@3�j�	ݷ��њi>=I�G��2�/<o]:n�^ܨՆ�����,m�3L]�zv��$@i��+��QW/k@�O(��{񘣓U���p��=e+4]gD���ՙ�������t�
<(X*"gpj�Ȉ�/�m6e�)Ń��W��;\���5l�L�b��}�ø����$����<�0\�Qm�Ts�Bi��E��e/���m��;J���lWr�V1�#��Îܽ�܃ۍdzv�} Pw����yr���8�TV�ʾ�_Yl�:�j�%��'o�����E7�A\k��.��{]�#D����uy���XЙ�A�]i�1�]��n�c���v{.'T\h�\����-�;N{oiTr�oZ�����x��8�[]/skHqv�ͷ����Ƿlv�}�P���g� dH���܌��0N�r`���"Ś�zr0���H�{ȯDy{w����LOvV������w}v#�O�ۨA�ɷ����!��s�f�Z�vҠ�ò�f�c�mrφ��/;�e��P����2�����B�u��-������C�����/l��L���cl>Yz�P�-R���ӖF��'O]�S��ul,}����!�ֳk7R��' h���-Ô)�������cj��֜���:s�o��d��Y�0˥��$��
�懋��Ó����ԽmAb�x��;��rѢ�[7Q�1�R�j;Ӽk+5wq��PC��������X窮>(�k(�N��ZچZ2�̩�t�pw����i�9�F.�MV�s4��E���,��ҵ5;���[�|�i�5Ԏ�:�\�o��*�G�g�����>�W}�XP9�+��(�%�dB�n�Y�$)���4�G���Er���t���Wc}��V�(���;{9g�{7����3H�Yp�l�[�^�p�b���x~s�Vu����/���P>��eq�JV2�VF�ԭ^Pg��ʞ���m�e�]�1e�,r�dM�w��t������\̌mw<G�Q6�����ZjJ��A1P�hy]6*ˮ�ב�b�]ҭm\��w��i:Ouj��/z2����L��WG%��C�N�������>f�v�ml���Z��fj��5:Tδ�u�pN��K�5�]3G=$��z����EQXŊ*�E_�|��X���@r�30E�"*�

�J�V+QbV���$PPcE���V,A��DR(����D��*�8����2�p�\�X�V����VE��
�D���*�(���*�����U�YQT��
¥(����A�"��m����TDAEƢ�V�QER*�Af5EP�P11q*�J�dmm��b��Lq������V*�D����QZ�,�j8��Tb�
�@X����DU��Q1��9�8�Ub���ت�
.4��*��AF�"����U؃�UQUr�b*�(��b����VQEr�\�DX�ETU�`��%h��X�UEES0�E��2�*��T`��Qƨ���[UE�[b ����Z�-,QDc���UQUEV0+A ��QTTERڪ��.&.PX*"�EK����~�ov����q]AN�	�&��=��<Px!k�����Kٝ�܆�iٵyO�/�����c�)���������+�7����ϓ� ���F�>�M}ONb�J֧���1�U#��׀��g��1�y��3o oO2���(�^�,�WlWY���V@���t�m���(s��a�u��RV6���jƙ|ו��&-Pp�SI=��N=!��;�=ʯr<pZ�Nr�5N��\ow�z��,:v��{��"��5k����m�x=��.����n�>X��xN���Vd�t^>v�KÕ�Ղ�}0N�2�Al �;#ʞZ���|i�WU]�t����B������n��|i�T��#иxZԠB���P�='#DUח�@_�Y��kK��Hm��F�\��~����-qZ|(��]r��GRg�"g;'�+���A^�GfU�Ʈ��-�<0�C��W狯��P�Ī(r�j�7��1��h�T3PGV�|D�8\%�f>�CR�m�}�l�T�Y��JJǡ���0�^��� 	����z�_{:��w�{������綇喤��6�u�k�!rF��K�AquM���&[N��K&������i_#p��E��b�]ۉe0A�������;�xP&��ȵy�		ҏt�)�[3����͋)��W�y��C�>ʼ[#���QJ����xd�Xy��RFAS��Mǫk���zn��fr rԾ��J+SC6��}�	���t�1#���\p�S<:rs���Byq���P����u���'7�|y�Y��n���Δ��1��'|����EZ ʧs����W�s�D<�$Cu����24Z;�[=��>ДN
h�R�U����NV�M�l� Y9�X�w����_�Β�$��jl��G�X ='H�5���i���6ñp��������x��Ks�n���N�-ʘr��5f��	_]�0��iC�-;1�˜7�e�i�I�B�ݲ���kz���sJf#V9K�b�Oi�49�%�t���@8���������x��9�r��]��˘�~&7�K���ϔ�)TUu<D���� Y�/�fr��G��}���s�K�]Zk�m;�ٜ�P1��4$/��C��Fȇ�D�/��ڐ����7ZTV|ά��5嶡����U��2����AoIΈ|yC�k.���y�E��"��y���f���]ʸ�o>�(f�J�l�vJ�B�J��nZ�;���������Hb�;��% �s=�J���(���m������s�L�Skl����������ׄ�A{��V*�k��yMڸ�jyR�n=vɝhUt-�'w6cU7:�X�oq𺗖�}���x��J��c��ܿy�����.G8v�x�g��#BُD��:�!�B�/��.^I��P����~~��˽�ހ�ХV��L��t��4�_nj�p�|~�+V��eW�0���Z�7m﵎|��{B[����7��"B���9��lO�f��`o��.�G]!�@yӷ4���b~|�<�xʧ�hu�@e{����9cg�b���(m6�����\����d��>�s��x�9u
��(��N�}�a��T�UM)�;��2kOOmOvAڣK9{Ɠ�K7�7Ӷ�͋<��V\9@7�[M1�x��3	�D0�"�����ԫ
j>��;<��ݻ��z����(���ZdTzcH����*��b����B=�ܱ�����)^�w�� �$9������v4�]�Ծ��*����sc�˝u�r�j��.X:�L��]��wj�=tǄ�7��{��)��EQ#B��v�=l<��b#}�k��Z��g4��b���x�%�.c�qOڷ3�	��h�d���Ȟ��S�#�8���x�����h��r��CH�v���n%{�;AgDO0�v�����Y*6����7r%?�ȧ���Է�9�T�vۛE��kyq����j	^ln��xy�{M�{�T;M���诽{��֮�����R��ٳ��sps�q^�����d��K�����_|'r���zy��w�Vz�}�Ƀ��]�*�"X;����G���i�ʩ�.N�{ix�V�'�N�?0e��ʲ�k)*�W�\�<��̮�A�tu�3��V$/��`.ޠ�1iSo*�{.p��k�6e��7�~j��1�^X��0�oL�%S�\�G.�:5�Kk��۝(��'��v����߄��>��
�ϟ����ٕ4z�fw��W�J��C�NB,�J�*��tI~gI�Tvt��Ġ��>3:�����9��q^�pcC+�sּ��|�.�gD��Y�]h���-�� �%�����V�X�MRȹ��O9Cc"�+���-a�Kf�����PѨ�w:Д���N�CC��麫t��ÍC;�vS��
�>ѣ��\�up4a>�_*ҫ1WK�'C(p�eeV�bcJa��f�l�+�T�5p/+߄����{�j�Yx|3��y�+��ļ*��8Z�(��h�U!�?1vj��������b�mˡȘp=�Y��X��-��Oix �:�l�Ґ���-��c�bō��;���tQ�<��=���� V����"���t'�y��	�Ӭ[�����5�����^��R��k$�]����S�lo����FȎX��`7/��w�?g����}x��ks�_r0�*�͏c��꯾��[�=(`���t��f'���R���5�IPҪ��s�|�1��V��͎��W��М�P�����$k�Oq��6à��Th_5P�gÊ#M��%��va��]{��������{ì���4���� "����
sX04ve���HЮ�4Vs�Vg��\�)���"��'����E���-�4��(5銴R��~�
KxS���������ۜ�Ǜ/�&`�&� ��c��(vSӘ���3�৪��t�*{���c�5��W��Z\�!*`p�J-�rW�|F��Gb���
�-9�tÇ�v�� ^�3jL����W>{��w5�b���(8|%4����U�Hiq��x�P���'�<��z5L��%�c�>�8��<�t2K"�AW�Y�T�*y]�Ic�L&xʸ��6��S������cmh���g��X)��-S�����
;#�&%��Z�t��N7�������W;���L�E����=���Z=(w���ZԠB{��='*�DR��2�f�籮����_ν��m^'�E��m����BR�ѩ4�_�+o�o~z�`�>����0C3QX �y�S����K�cX�4���W{q���h܋�p7��R:��T{�����K���/+g�)m��������,��y�i�U��2R\/���R�q������Ȩ X}�=�6{�]2��)�ۜ��6�=��h��a}u~x�U���TP��@k<�(v�w���	�O	Z����Vx��^\�;�:��v�TE���^}A�3U[�}�t��B��?r���v�s��ֶl`� O���ȢʌK~,A"�R�xf���ׁC���)N{J����e��ɸ|���f��y�F�R����߹͡/�Nv1y�Byq�)�P����>!�+��e�쮒-�=$���R*���48xi7�xL�`s�s���{���h�Xw�󖓨+{�����`Z�>(F�F���������Q�2�Q0�
�����m�ݖ�4D5�Yn8��~�D�{����9��@x@����M_Lz|]���x�4�]�����c��\�}ڊ�ϓ��8�[
��B띘J��ɠ�z����au��{��ȧ7�����ԧ�W��z֊�Rף���(1��4V�#�.^�~�N!	8����A\��T�uږ�$�b�����������Y��^� /f�o,�}��V_�_=%q���{m8ͭ?SG6�i�uk~��ָ.YjX�xzu�t�c#;��������Tk��\�Z�6;�l5->��g�������$�^^g�C��m��Pp�9��P?��Q��\���Ւk5�@<�evL���G�{$�۝/�ԔW�4��{/+�Չ�a��6�!}���1x��,��b�~��1>�ҕ�s�Y��Ĝ4�٫!���*�z�]���DkA�!}�ȶ]�ݻ�Z�s�z�@�D5��������ߊ^+�p�+���� ��յ�֔�W�+�����t�7rI���W�hp��ȱ�1�AAεoЯ�>��*�nd��C���':�6wd����W^NVӏ������+������XѮ����r��W��\����/�ۮyh�"SŢB=شL��_=Q�Y��3��O_q���v��*�}�{v}����s6="���Z�+���!/q13�`�WEOMeTاu�T��aH�.,����u��#<>淳�z���w��Z�/8��=��.�1��S���k��Z�t3;k�l^bJ�`\����>P�=_7�Q4�|� ��K������a߹MP��s�[r�X�~�5��Ľ�aY�
��\Wh����2��VQ�o�aH�m����F��2ejb���<�G��:e�]`�C�so9��]��:���H���#��Wp�r��t{V�t��z����C|zZV{<m�����hn�ip������=�����%�ƿ��*��������:����bK��v+�_&�σӍp~�yv��ͼ��Q�nJ�W�UY��ō�����:��ß]"�i�1� ZW�ZHʍ�U��}��l�ֻ�{��o{<w�\4��@��4.��v�����8eTH{�"ѓ�s���mV4�h�/����Sz��fp^ȝ* �܁�=�U�ᕶ��W��q��J5\��p
|�5�ޡ���:Ԭ��s��߈�Pi-M�^�	ta�?^Kɰ���P@
5�U��,J�/��T/��T7�}��C�o�l�g�mjv��?=������hu��B	�p���<3�Fx(����ό��(4�����W�}��q��0��\�t%�WS��@�3j���A���Q@������#��@�%��*���(>Ze�y��F4�G|�/}�+q(1�ό�i������D�wm��T������$�r7�{�/�E7!�>��z���OA��[uo���a�a��=}�����5uڭl�Av���]�~��D�2�+T���a)����ŝ���/c�uB�=�V��
N\�^�w��q��h�w��Qe+k��w|'@޾q��2R����1Q�)�(��w���c����gVo�Vr,���}�Վ�B�.5���v�+�]��e�v�|{��ʠ_aP�5�ܰJ�~�������7U6Od�j����է��=F>]u�)��7�����LqC|��"����Ƿ|C�\=|�\ُ �V&c\��{_�<��62�c��c>�xa3�E�hc��g�T�����o�������>�tLJ��4��S�PV堠�%İ>2�%�ҟ�h�0߮{�4Ō�3���k`�;A��b$��>������ uZX�E_=~=Vo��ܟN�H��=�|�ޜ�
_)������&z���P�4/������]>(V�O��o��}mrtm]���߻d�~�d)\E��qM>�3�
��؀�&�2���s��04Ul�#���g���;e�W�ש'�H���V��]s_b�X-���3�b]xWS���=Y"~*�� ��tyݏ�~�從�W����@-� B�v�4��]M
��Y|7L��[�Z�b�fz�
/\�d}��c)��b�A|��z�uCF������[�x��
�_¸b���LgŃV\�-���ͣ!�Sϵ�{��XUo]ZS>@E�E3H�˝�n��3��S���e>8��R��Ȁ�<Sʻ{̔܀�gm�Ȑ��6ޛ]P���ӷ�2��x��+ɋ�}��&[8�j�-��.��ڴ���(���4�9�I�h�h�CE}�JϽ�B�^�U}(8|%4����T����z®�6#�J�xƅ�I����������9���0��p4�`�F�w�cm�x?���������mwz_��,��RU�+�|<;LÛ�X/����d��TvG�<�P3�:Ńm�?7ޝ��8R�����-���V�Oh�_2򔰺-+9�Qχd�F���bI��K�W�#,!~j��u��ږ|�mC����|�i�)�]i��u&v������wn�~F�wy�[��wPm�\ܮu�CӃ�ݥ��I^).K�����d����R��:�W�Qm�w{�����<�MP�8����>Se�@��o>��K:�@U�py�i՞��^՞��R��9���ؘ��	�>���"�V%䡶��׈�/3�e�2.w���8�į1?{#g��Ϲ�/�č_"T.z��m	`rs����e.2�yjV'3Y�/)w������8u1e�A�~I�ర�^upM؀�"�e;���J>�W��T"�>�.��=5��$���&�m����d��Y�2%۩���Ę&���f�����mM�Lr�r�	�Р�+3�J��Y��4`٢�V�2���䢨�*�n^���e̱��素Ӡ�N���=.y�鳪��9�H����M���Ę�#K}k9υ��Z����y���]���'��o����WU�V�Y�p��)���{��Z��TG��hmu�7�;�[��A�m��e�̻�r!�`�tT�9���̆mYcIK��]�I��U��n��ûWr��� u���k8��s lPX[w��.��P�V��Do:+$���Мŵ�m&�oL���h`r.��"�J�շA����Bh=����3�L�f�m[��糪�SgG\T�1��*��7wKȿax�y�7�RYu�.��l	�"Ë���T���R���)���l�I�/�^�����yM���A�y�c�Ж<��y�4�T����o��� ��y��fm�Y��Yjpp��;��,�__Kv�&�jV^������v}���U�[���]x������]NM��	3��Xn�Y3�"�9��0�3*����p��>:P'{=rǸV(:��X\�dɺ�h����x�Gg���N�bݘsj��n�5'RuZ�V`�\롛�+B�{�@��[+@��Aމ��l7K�F���)d�iOVv��in���:C�u�����7�jmA�;1�z4�Lt�(������@ab[���f�F�
�&�r��eG���'� ��`����m�4���"g��]�����4(;�^�Frk�DB�7�ʵ�]���	%)�W�j1����]�_iņo;��Դ��<o�y.����)�o�S��>S�#d�[�+$���>�߰� ��DZAA�jJS7�s�h�*0Vܣ�gӇr�`��Lv��j�\��B��JkS�ISS��N��4��ɼ�H]iyK;v�8h�6�&6B���y��\x7��5F���<ЯC�;{��^I�v�������p�$���7�{��g!�RO��ܥ�����_6���2;����ғ�0Vm���Jt�C3fc�"�v-�vj��
���͋5�r9���{�,�յ�]d\�֔R2cO��r����3w �Iņ��;(����DY'��Oj^k闁0 Ne�
�ʗ�Đ9M�[�He�nc!�^�*�g:@�pR��u�ⓓ�kH���f]�i:��CR ۩��֢�a6��g��d��7�ʍrk,)�XV������0r�����[Y�{g5�Y�ғi��.�L[f]+���PL��l,k��;ڼ�BL.-�9qZ;�ٺ%�[LN�hc-d���꛷�'v�ѡt1}̼�8�w����;��	3~���Ŏ�J�S��P�Ju��zR�92���pY�MZ|=�W�eL���&�����1`�b�h�T@Q
�ҥDcZ
��������Җ�Q(ѣ"�AAF(� ����X��E�*�V�(ŋ"-�YPQ�*��Z��Z�(8�Q-,Q��1Leb�ؠ�EmU�S�*�D�
�U�1X�EU`���bTc+PE�6�X�b��J�	[F%���YQV*��"�&Z�"��(Ŭ���2�����%DH��j
�����"�m��E��P��J*���U����D��(�"�b(,b*��K���-h�PU?5b�,b�PU����?~���X�����0A�PEQ���Ԩ�\qA[h*���d��*��j��
ŌPb��R"R��+�ĉUb�*�Q5*�b�*(�)�����#�`��imTT��*�1QV�Em��R(���[i,ET�V
"�PDb�Ū"1q�f>����u������ʣ���m7@�[9��ΛX뫰ܝ@�-�\6.��6Y>�Ȼdݭq�-�f޷�=�����	��p���H��§Q"���U�U|�j��e�a��7�2D�aכ�#.��Y�}����9��p��H�z%��Z _5���i��O�.����}ptٔ�˙��j����\��S��Џg��������_i��KC|g*aq�]<�����5=6�r=^�_���@c��=7�w�2/Z�����*��S�hs$2K04W����f��}��p�4�ˬ�>d�p>&7�K��P���*�4I�����45�WjZZ�?L�v8n��n˛K�*`�-j��0��KL�� ��eK�7�����Fc����pT��
����!�մ�����;�����eꌡ�B"�z��kr@���{���q�`��g4?�x:�!�<C֚<%�[.�/���"��S��:����A�p-��^����'����*<#F��)
A�X������s�Jd���7[���y`�w떃x���\��W%1_,K~3���X�p��V�X���4�MO3��2�ݫ:���K��GW�k��9���|��iZ�l�Z���/{I^�0�o����C9�e�x_�}~6Z�����a�������^���|p�1�i���e��.Vr�ܢ]~D�}8�P��)Q|NG{�3�I<�Biai^ŢB=]�Dʧ���:��?x��H�3q��|9��ksk�y�����1�X��pS6�egU��ex�p����wߺ*zk*lS������#�a��9��rx4/��כ�h_�k�����=�zU�"��8��qW�ε��{��?F��׿�R��3��ېw����xM��Fk�{�uu��0��bf� �gX^���%��j�@}kL��!c b��wǍ�E��Z֢�|��Dm��qJ��Y˲QlӼ���ڞ~�zsO��eVG��5��V�T�lB붩�x�.��@�=0���O�<G1.zc�UW$�=-�~4�=| �i�g��V5�>�w�DH�'��cW%��A���QȵxhG�S�i\�V+�p�κW�;�=�ng�9�
D�%/���\o������^���su�u
>H\%Y�˫��\&�6��es������b>$^�T]��orU[��ՙ�y�=>�@@� Q޳����ye%O�����_5����:::�q��mY�)��o7X�ce�硩
�h�9�w1�������׼-9�Z�����T+�॰X��a�oSx6��wRz�r,�����x	.��kj�Վ�:ߴiu����e�Z���e>��<^������ʘ��Q�����`�'P%A�b���,A�bB��dS��Ycb��.�y`~��0���y��U߇���^oy���H~�oUp5�r�ё�LJ~��8�Hz���J(���6����ѬE���A�n
x:�畒��)QN*t��t�UGgJ�q(2�`C��i������>�K��]#�*��ք��.�cj�ܱ���U>��� ����1����ʥջ
�YDp�w��ѱ�ȳ�3�>�]pڬ*8j2,�~0p��C�>8hvN�f[kZ�*���%��o�{ե�v�ҿ|���·2�*�S.���p�ef�b;�͏`Yb ��u���r3��pg��U�^Ø�Yx|a~=@7�R���~���k<���E��[�o�l뗳�����i�}��b(aͱ.�#/�+��/>�Й$�J &��{#��]��k��� � 6q�{t�1==�`��T"��HV�%�S����#�G �x��帲��/��ҩy ��8H����&{�l:
�F��sV�,v�B�;���w�n�=]�h2�gU�9�g�Y�i{,ƒFM���I��9��V�¹
���z���1Ux"�������}��o�Ω[)��?��ߟ2���/yKlck;:�����ͷo���b�ӳ����Hd@�(�D�{��,f*���8u���[�i�Q�PW��d��PS���D*]B;����3c��;�g�#C�� lί�����ȱ�[ji�Pk�h��?y��(�����pf�]�)z�R�bS�̐P�HC����z���-���#�(o��b��Y]Yy%��б�:S��Y�OC�L�� HΖY*��(Sy���u3�t�x�l���u�-99������R�Y��R5�b��Pp�SI=��r�U��@p��v�Ow_s���i~vx��o5d�fK�Cd�+��Y�jȒ��M�%�� �5�g����V>2���w���+��;LßoE`�� �N�2�[ (�=�ݾ�Ųg"1O���Z�5�Ƈd���,���t����3�\<
֥��<"�;!B���9�G÷3F�#�u�jY��mx��������V�L��L�#�|���3��ax)�C�^qt��@h&k��R�=�v1g��>^W��V�vƒ�\fJ(�+�e`b�!�հ�dj�ǹN�YN��aRB�K�����<�
Ykc��<6��\;�� �Ҧ	��k��F��Wcw:+[��WW8��`u��9v�̽��Aڝ��x����*�&�ן�շ�����w,��(����u�JK+#z���
��>��`�+�W��f\J��d,�=�~��z6�0U�f�]��b倓�`�����s�A���潠I�o�� �U�(w��K��b��q_��P�u�k����Ǒ�YM��XKO<�	S��@s������ȕ��{�shK����_��T��W�����~���j�3�١�k�,�k�R�XXd�����ꭘYh����5ٺ���>.�b����l�W�ϫ�Ȏ��$C𾠨��+�T�U�W�:b{�f�A��I�_x�
W��3�k����gOadB��,�/����4��ǥ��\k��*纤^���3�2���J�'<�*)_)��Z�j�d�}v�g.��+��=��]8;u��/���&u�q�r��AQ�A��R�A��W�,o4y'�f����-����̓�Mw���_��eY�ǭg-��Yʃ��xF���'��O�Y^/R�3�·��3���)�
�q/�<:�7���\%^��K�hzQ�`y�$�V�~^3���s�*������&�V� G)`e���jnr�ц;�x�QqoXq�x�h|�WXg��7����E��_
s����#��Ηo�����#l�U�cI���R��'ίkF�܇�`o')�^�\�f��]2��3	4-r�5���u��.�r��`�jB�?@s�Y߰z���H�>�2]T����#(4��v�=�_r޲��tQ��8[�s�hEp��&Y,:���x8&���`��������N� �9�+��e�8�u#�=��<{F�J� �7����:$/޳����uI��~͏/��S˰���ҕkؙ.�b�:M�=����&Z�k���ޭoO1��s�]2�x�;�x`���^�!��9v+��ɲgq�wOT�W�%]��������Uj|�#�H��%Ь���n&&53�����˛�)�������ے����H�=
|�5�C�s���=��.�U1��ya{�j�jnM�[��|&e���^��-�/*�������ı��1�{����yD���1EI-�[��v��&1����p�z�.�/쁋��wǍ�/�Ե+L��oL����۰q�y�.���3}���� d3O��b��E�5��l�LRفWg�#�du*��U}2M���OxP!Q��1�kB�0������Ҫ/q��L��]�
��^z#���u�9������s����8Ч�}�x��yb)��;�5w��h��m�{�;�LL���w�:��H�M�����Fj����N�$��-��l�92㸳�+�]��E��H<�U<h5nz������|�����`TQ#@�����Eź��|ۻ����upE�ɋ�i�ѕE_a�_L��x4{$���D�pNo�Y�C�����R�=d� �8�K�H��s�q(k��CF��κ%\U��x�h��ئ:m���yI��k".\5����u��UYp��J��!�'�﫜ʱ�N$��l.w/ۡ��=�ƽ>)��H-�0A�bC�}�p����<�/��ԟ�F�iJ���ؓ�(��^s*�U%�V���C*K,�c�
bPe?Y�U�ʾ�Bꯙ����{���G����F���=i�`�WNʕ{�v(����?C���-F���|�ٙ�9�Wo�z��(�Y��J�G\�)����N���`��
U'��}Q�q^��e��v��g�q�����QZ��곶����p�d>�r�+�شL��hǱ��m��c�-{}���-�1�.as3C{Ps�W�xq�=��ӑJ��LJ/W����;�����j��Y	���c��G��Ծ��;��W�s�}U����j�8��u�V� �v1s�����E�l=�etMEݦ^Q�j�R{�t�Oa�2Jm�dLl�"�[���^�f�U�%[��h
�$�t��<�]:�c8&�NM�
�ULZ7L�|7tZy�(|�8�@��C	���З�t�bY}�y��$q�*ا
�fA� ����ʂ�>��l���	�O�93ʲ"�/u��0�7����$ھ *�L�P�f/ d�%r��[�1x��!�̫�>��%f簖�I����{�&�>�pvR��VԄ��WS�=,��6�0���9�e;ܑ��SVc�VuT����#X���q������Q�PW�XO-ℬ���Ip��َ�E�gMEy)՗�8-L�W^�A[B�'���s��ȱ�m���yA�h�Z(�u>���O;z=�
k��Иڞ+��L@@�� �W��ӅVp�k/�鏇m�-�M��f�s;y��z���1�U#���*T4hJ^��|��.���p˧�?*p��X�Iro��;=�N���]~�C��5�+11h�>��S�_�:�K��^g�/�B�6��'
���X�/}���������$�eIdW�*�ϊx�4�`��˔���4�q��޾�Ч9kW*PI_,"�͈��Tś�M��tDN>���4�G��΀���;�,�^�s�/.��A�Wns\:y9��6��iIOgz�����B;�rxӂ*=��;4B�N,�
	����2�Oa�8&{�N�9M} o�*��vu��Lj+�lz�v��>ފ�}��2�[ *���>M��˜���N��|�S���+�T�hq��m&ii𭢞��r��p�*��@�'κ+_\ә����1���NY�6;	�Ws"��n�xl+���?fu�,�
e2k�S9���'���e#F��掻����LW(hX}��'+�S�QV�������sJګ�4��K�{˥rHF�O�3v?-�t{��m��zU��\����Z:��6��V�l�Ғ��y���߻3�9=�Y���/�Kj��| ��؎媜�OO����\U�1g���謄���׳���k2�Fe�U�~��$h��J��B<9�%�s�׫e_��}k�h��@����<6^%�?jR�1���R��x_�l�"ȫDw���{Yݭy�u>;�.�o,Я/��m8���i���̥�ϯ�2r��bmgeo���]77�恠1>��U��;����lv}��1�OD�i��4��hp�s�g:��(U{$�Ӳ�?`�)p�q�C�Sں�O/uz�y���VS��J��X�=�����4��v���
��W�T���'u!p)cD����p�
��b~:���X>f���2�$�<,�����+���p*xzq���3(i��s���G��)�r[���m��SSP�M�+���zev�cZ�B�ل��#=������5ឋ��ߝ'u����s��;?Z�c��q��d���e)sTi��hz�xNΑ�}��f8���ɕy|9g�p���]ga���\���$������"{�Ȫ��\�u��9hڑ�Mz��i/��\o�_֦�/Qس�Չ�a����ݢ�7y��j}N�זk95�9���X��G�_��.���פVox5pv��+G��篷�f�z�'�"�/��oIΈ���!��=��Y�x9<��)24�kj�;<v@Q�X{yL�S�*��c��	�Ɯ������(�l�!x���+�*��ee-~����r�cKCܽE��tT})V�=��ʛ{�I�Á�L~��#]Q�sR�&[��Q|��}}pnW�@��P��-�a�"��҇L��VK{��'��g�6E�6�c�qƗY�/�GE6xU�ԅ}�V���x�p��LL��`�WEOMm|=u���{��6���|�3����1`
̲�*��˪�������A(���@3Fܾ����n��X�A��	!�ȼ�[�˧o�xO�;���.���b��b_Y�{���W�ͷ��=��͡[�88�kN����]TE�pS���G�klV܇c�k`N�eJ+D���:����K{���S�=���}��#�{��:�	x̽�z)ԣ�T콛��_I;���yՔ�x>�0ͺ3I�����X�/���fJc��V�����w�g���Z������'�l���
���}�A/!Ѽy��h:(ws��XB5�*��xaT�`��/;��CY���%D�Z(�R:F�kx�vg�:��`i��P�#)��	_U�=�G˻�:붹����+z�J*�����P_����W:Jg�D{�ZQ��{t�kI�7\1����³_h	�n#yw6�gX��k���0���6"=�
�J�޽�S-��ӣ˜����gt��75�1xűRN���B���͆M�))��ô���9e,%F�47�'QdЉ�L�q�7��JT��0��I��gN��I�}���^���T�ul�k�У]D�ٴ�W6�9��h�3h���NV���Pt��j�Y�&�f�M�ư&{N�RY�1l��g	Ѯ�30R�&E(�!U���&����g^�{֤2���fa��VV@'(��h�\]�C��)h��[��d�u�$�ׄ臫�u<�n�s(���H;��}{�+[K���\��EFz.͜�����SR��8,Ps���b�+��*�Ly�kjԾXшuÇOt�-��SW�0��v<���\�>"0}�,�π��=�0����0Si���cr��Ӭ���[)2�T�	b�ܡ�uD��b�ǻw\�#�+(l��0Mʄ�'y�>��@֌���g{%&:)��ɍn�z���ؕq�+���:gPB�N�.�����	��bN��FQ�	h;i��a�n";m�J�,Fw��[�l��m�.�%�|���"y�A��ӕ�o��K���o7=��O~�"�:o��j�Y�Ԍ\�f�"�6��Zc�`K6^��B�����JH�����Gx��]m{3$��t�9�W�W܈ۢ�R�	r��=��=�`��Y9�J��k�Q�ƟL<�h����v�P�R�����8��:4����nRF��Y��2�=0��0){Aد�-���(�;�wGZ�Z�P���ta46'�,�w\��<����+7!u��a�B���N�kocIvVi+��x�I���P��X��t.j�e�,A~����p�� �K��nT����e6�����b� R�s��]X�m���#eX:��:x�K
"\�F�d'w,2h<���l%���@����<��4�f����X��J��G�%�S�sm�>C7� �՞��a1�H֪����F�RZ�Re�[Kb�Z*b�e���#i����F,[lX���Q�PQ��fEUm�-�%X�
�����r�9j�bҊ*.4B�2U�YYV��J9F�(��l�*�(����EDV[F�U��#��d�����b[,A`����)m�Ŗ�QV9ZX��((����.fB����m�V(ň�~KdEV1T���?�fY�`�PX�AE+*�f\J+Z�E`��X,bȈ*�-� +��*"�AAX��ڬQc�T�+.e1Tb�#DDDXVTUY"�h��V�qc�E��\�c�f
"�
�ȷ�1�Ym�ȣZ�**,X�I��A"���ZV��3$�b
,�0ET`�"1 �Q�6�UH�J����D_7s�}��F̽|�gW�����j��_JL'�}L�ug%2�|z,��{�Tz���Zʅ�m��:�@+3�Z��om�]�Y��[)������Y�Z��B��C�ʾ�3kӮ����Y��yY��CsO	]mW�W�OOL��:yize|�)A�4�����Q#[�P�j��C�/`Ws�;�c�G�ST49�o!c쁋̕\x���ֵ�E@6���;��v��ؗJ�jU?>��s���2��,B�>Ȍ̯J��^h]l��x�쎮ޏ�(Řa��}��y��A젮̾u���QS�z �t��x/}�F|��h��`T[��t˘��9������B"ɔ��Ϯ����d�v�xm���qht';������ד�罴�Zr�z�t~�����U���*�СKx[%}g�쫫c�\&���Y\�~������
�o��Z���'��V��������}��
� Q�vx��,���^�r�v	��5�\|�����N�_�3<OO���|`�TĄ�,�WaU���p֎�#y5��-�yzR~�Xq�a�ޙVK�
�s1�Ϥ���8����o�WZ6}+PG������Ηh���Ӑh�wn����V���r�V�14�Ew�b�r���QT��4p��Wj�kÜx�D�Ϲʒ��N���2��v�Agq�K����Js��}9���ܾ/���X��1lwGqr�T.{��f��1I��N�.�g�j���޺�X�謝r����А�>'j;:WۉA���s�G_��=д��n�w�>�`zTz�<l1�Sō�r�G��>��� ��<��eg5h�<2i�9�J����O����>��9�pU�2�p�d;�hJuشI���MO���^�{���>��M�u��R�i����\54�}+2xWi˦+˩'C�RО�d��g^\���=o|3�ޣ�8���ؠ��Ň1X�^��z�y��ʁ���l�x�e��꼝�07��*>#�T�̃�u���ي��KA`]�QyY�����*�GN�ۑI�}��Z�p�������UgX��D=𓮣��݃�5TU�W���g7G�n�������̜6�6��*ڐ�� bZ����(8�5Q�|��������J����Dȅ��,�����yJ�,e[�i�PW��M�e�Z��p
��ŋ���-��L)��_V�";*�F�]Pb����]]sY���A�zb�/��R�wi�Mһ.�7�����-W^j�j�w�Eb��%�c�d������K1v���۫�R�Wn'x�b��=+��G��uʒ�%%n��[�R��:\O��i3�s����6T8����o3e�˨�B��jv�/s\��S}|�0��g>-�{I=�ӝʗ^���m�=��W�Ș̘�� @�H�Y��
�O%�V�����~�����WV��:�c֨	���R��<9���b{�fu��i��ozG��Q�9Ը�X��o�*�!�9R�أ�Hו�*�r�U�$�����6�߬��{�[�>'O
�tl(y����y�%S0@�I�Ϥ�+��Y����_l^�o�L~S�/���|�,)E���_o��.��qp����� w����^� wQ��hf?{�M���I��hʊ�Ѕu-J����W���R���-ѷ��A!��p����1�����g��E/�ۯ	U�-�MW�JK��>��iV{s)��0�f��ۭ��˩[���9G�^���MLwlU���: w-�>���0�H��Mk<�x�~Ɋn��x�Mo3�j<*SԩÍL��Q�<K�_���νz6�bŔ��i�\řQz�aJ�����f_��Ȁ��u\�g�� Z����YS�L����}�P��o]��.7����X%\F�|Ϛ�4RC����Nxfic���Ȭ8`��V�}�5ϝ6��Ӽ��+F*�Y�-�R��^��v���F�c�V��;:�*��]q!`@�gwf����o�f1�E��#��N�olk�b���Sm��29F�O�7{mF�1�����N��E�M�4����H�"U9͡/���yM��[v,vߍNۗsِxVr��(e:��<8�5��Ldn�.<����e�����Eͩ/�z���QW��г�}[}2q�G�ve�ҢD0�𾠾'�5D��R�We��M=
��>��_��2j�_c�l4g����U�R��~�����H�'�%�ѭG��0� ��gtJ9�����܉~��LV~��y�Bb�zw�3�*��<���pV^)��Z���@���H-}]���y\k�&d뷆�O�VC��:v[��ԻΎ��AQ�A����U���V�7޾��zn���v��~zhM�"t������@7����E`�Yʜ�C�7��F'�몮S��fnd���o�A���/w�,�����4Ǹ�W�wb��J~����>owx'�D����!���@y�-���8���e�s��5h�\��'w�5ﯧ���UfVvo04] ���t@j(Xc�F���־��x�C�o�c��'�d���Kpt�7:�7��p�Z<(����pV�����������G��U݆��G�F��L-�뭖/]�M��}�eA���5���]�og�K-QӬ�v��GqSS7�^A�F�Gh�3��x�[����!�st�\�m�չ�Ot`�g�:�-;^��+M��n��G5�[�Y[�W��*��c��x��*��4-�P`�X�}+�(��7W�Xrվ׳5�>y||*��~�P���<2�%rTǜ�+3�8F�"���U�����k����Ӛ,V6U����X�����L��OT`�M�;�&,��Q5�Ϙ���z=���Ik-;��IL�Y�I+�Ґ����t8Nn&&53�.砠�z�Y��/�8]�� ��MןKp�m���E_5�C�.cW�O��jP��3�+�k\q�Q���F�fg,3�s���}k;�/*^h�ť��y�)�4��]��7u�n�s.lŋ�g3U�H��MP�9��,����wǍ�E��Z�|
�"���]a74��Q}�/�â��^���
��D3#���s>�J����wg�RF\���B�w8�(���8#9t`���}mS���Nm�I�g��5�0SiJ�!r�ݞ��R����F���,E����4X�Yl���+F|^'��T��E{y1`Z�I�����⼞�A���	1;qm�����}j�꺘-r���-ӱ��d���GГ�:����l���9�)����/�}cw*3f�9*�r	§w
�s��a_{I!�[�W�͙����޻};7�����77���V���{�/ՍL8
��
5Z��H�{~��9e�`Xھ5��{���^���ۭ�E�����y+H��1 �� vxV\<�*|W�\�p�w��m�����Nm�Ş��*©/!��z} �6�����1�YA�B��nu�۬��Z�}���M�F�G�	��ч3��d�`��s1��,����B��@�33�ӮSlg���Fg��k��
�(hxwL,��<��#��'�\�ES��R_��c'�{ʣ��pD����^yn���l�����v�����<3�s���X<�}.�y��b�rL�]��|��$��	e��t��f��!<�綥����{�54ߩ}��^��K�n�$��7(`����ɺ�t��_����`LtK|d�y�Q�
Oi��*C~zo��7N�n{�����l�J�."S�=���=���1_������{*�Q����w���/
�����z�]�V��%�tZ;ҪQ���so�\�
�I��q{U���y�
������� �]���������A�Rr���-�\��(L�d;j4l�] �݉4��T������;D=��0�j�̓�%���V�Χб���Y�'�\���[n�7+��y�Ϸ��,�=�r��i����'��-���]�r�}�Ƚ?����J~`*{K��`���UP���3��ҕo�!������k57�����&Q:L�ʹh<���y��mHH�F��K*��/���29��v��f�[Rp�w �����tL'h*'a�f�<�[E���&\���W����M��rL9H��P�����3�z]4V�";)�hU�+`%��0���{|���-	R����k�ź�S׼���3ҌU��9��C�d����S�jy�J,�7�$�������J�29K϶��r��p]?j��3��V�Q�<i���^9%�:�P!�L��LGBY-e���l�s֧&�����C���}Y励=*P�dI�$�Pp��[n�c���vI{}{�M�_>|C�n�^7�=�����Ւ�� yB$�eIdW�e�%?���uq)�������#U夝CП���e�\,nC3|�/��\��r=#�Վ���Y��4�h< ��_<�S��{�{�2�E^�f�S���x*g��.�C�|ڬ0�s	�B�y$���B��4;��ЄG2�k��tkX)���.�?r�2V���v��N��^�3s�;,�J��F�mSs�}���3s��z@*��/����%�=*։��A���͝����r�<���v�������5��:7˘�X�E��^���f�� ���ۯ	�ط]�ayIp�KsƟnѼǥ<���ֵ���#��r�_3��τ�t=���MLwo�h૎�<�w�o��*<�UvߨΣjG�7R��u��u�>�ڨ���A�������"�}~^�z���0U���>|�gW*7�VG7�1�]��9n�X�K��#>�\ >�lGf���P�C�o2��b��\>5!�1����^V��(�5~R���K����F��*=���P�c�O�1�7
�/�^���f�x�yq��b����K��27�Xd�:�&��=�n�c{��ջ�΂��8c������.�y��o�iz	:GXH������5���hews�;$�귈��[^ܸ��7}e���v��ђ���� _�F�����m_=��6}9R�o�@]L�$>��_��3�,����%�Yx�Waǂ���`J	n���Nz���W9f!�F���"Ǵ�������a�z�R*�b���4=�Fu���B����r){�7VvI/�ï�W�c=~
���Lj�*������d�R5�V�����͈��5�����EcI[jh�Y��Na���OR>�/)����许��u:ܚE��ޑ ��;�^3��G��}����F�^�}�i��g�V�BGdq*�\]����]ga�p�9s�"Li{������<&��c�u����E�]�U�j���U��|����c+�8S����?�D�=���>�cN�Zd�l[�!�=��T�]E�}⬾:�)*�j�N��t�bL�=�I�l�zy̫*��eAT�]�Ϸ��V�s����<%����ץ� ���$�!�}��epu=�e}�q9U�R����B�<v<#B��Pg�``�j+ҧ'w��j[�����\���A;/Q�K�J�JU�bd��z��4���U�j#��돪UL�=�0]����?|�ٕ�L*á23شHG��h�]���Q�L���K��b�gȳ;�ŧ��ǺkXf%������VS~�}6�B�	{��;9z��}{�W�n��2V�SMeM�w^�\�ZD`UM�P�F���^p!��2�H+�ȷ�y��+�z�5�8�*b*�N0{�wxg�OOL�]�!���w�̫7\+�2��J�r��ĥ�
��{��,�����CF��y��嶻�L�γdny�����͝Z����O�dU���o۳G���E�$�1�J=��i�E�'i���Ʉ�����M�;��N4~�Ք"]1�o�߼��_��r��f	�G:�J�L {�CM� UL�0g���k�l��n��w��Tz�#��v��qu�{�fY�P6���dw��N*�<j)����+���">���͔��_l�����>�ط	W�����&sg�߻�̣�D��0s9tX�A�OƳ��9��I�g�Q���^�}�}皼�ir�YY�����4.��v�=l3E��&:Ƙ�^'��ng ���������=En�@��h��C����B�r�B���x����>;�q(}�wy�
7V�[��F��3R]<c�p�i��+�x�k������rb��-vxV\<����������^)IO��p�s�X�^CO�"OO���U خ�#C�G� ���J��wyر��#������0�oL�%U9pU���t2����S��A�%�R��׫q���k]�şN�+�B	�ؚ�V{۞z둃z]���*.]:%��%�t��{G?dJ�f��OWF�J�Z6v}��C�;���Y�[z�u��y�� ���C��ێ�z�t����lL��U�����8n����m��R#zl��	�:�lˆ�:�������u�����˾��֜>/ؑ�p���K�ۈs�E͗��h��_.U��ɓ2�6��@�$<v�g���V��u�q�S�הO�X��_�N nr����L�9�F�;X�eh���ۗ�}Wܘ%�g2RD��]��������o:�G�^�+o(�`����ω�/���#G^��f�z�J$F���㉄y�3%���(u�ٛB��*Yȅ��8�GR�u�1X�1�ָL�T:2i�2�Uf���b�rҹ@h�E˩�ඹ�GG̫w"�k�}�C���a�D�u��Eu"�Ut��B�iI<m1L�����A��|�`�8yyzVo�g��*�K�]gY�qm
cZ���^p��ۜ�K=aT*yw���|.��͹t��}x�t�[���\�����`Z��L���^sXv�v��&8�l��2�i�N�p��r�30i� �+�./�]±È���-�f��N��Ą�9��0�ׇ�QC�~�fU��-�8����[X�!G���fOFy�.�t��*��B�Z���j݁ 㺹R�
��ۘ4+R�-��X�L.�۽�R���ɜ�m3m�Z��>��Gtu髳!4`ƨ6;C�BO�uZs����Ql�ѷx7)��&i����e�˂��;�z��2�p� ��։_T�r�M;��ЩY��ئZt�*��U�U��j�'%1]t��[�LubHCH�*'��'�9��ve���\�B�����YS��q
,�y�.��%�b�Ҹ܊�;��2�oW_��I�$�B���GB������ �V�x;:V�/\Q�;ܜ�`ޥJ6��ܜ�_u=mf|�|p6̛�zbO�X�����S&P�ۻLo:w�>m��(�Re���7KB�$b���H\������"�L�[��r,����R����>r/j�Xs��Bo�����fbBgt~IP�{d�9�����0V�:��@B��\��ę6d��{_9<���&g+���nw��c���_ �uRۨ�{N�l�B�Y�:*�'�N*������3g����2��%���0����T���+:'U�V��������WJ�v\Y�{��`��|4�3���v��!Z�܏�4kZ��&a�C�wτI6���Xol��a#�ǚ�A�}T�r�wt�M�օ�˒��IB���:���=�f6�t���I��ͽ 	loZ2zN�+پ�9�AAJAύ�EW ��� �?���%��W�X�����qo�G��r��[�����YAܠ���{aV���D�F���o,碱���K+h����M���������Śzw԰��M��|�U֌��*��g��
�U�͞O�uvG��[]�+(����ľ��M�q���
 4j�(�EDb,q�*
�#mV"Z	-(� �,DP��+�UG)UEA\n%b��iX����r،D�j� �*�Pb������̥QEU`�2�-�"1m��TUb��F1�T��*&R�YR+YH��������S)E����LE�(�h(̴PA�UKFʂ"�+�\D-R���D��Qa���-�	hZ�-
�1�Kj�����A��"�,b����\5U-X��V!Z��Fj"cV-j���0O̢"��h�PAL���,T��1̅X �kE�"����E(�ŭ��?~
��AU`�*�Z"���fZ��Ec#�DY�DT~}�`��"<:%i✢Z�+�G!���O�q���.p�%*��i�{;`���X���g���C�!(�V�n;:��;s��q�Մ��~-o;��!�^4ք'��`���R��rޏx*ji�R ��v|��NU9{�ϗ1���%��m�����ޮ��џn�A�Э����S�s�]�F���7d��Y���LL��ã��N}6()���m�
�7y��<������U���̜��ҝa��@|+Y�*|GB���q��\0A���+r���d�^��f+�ݔ���bٕwpL�D�.���`�y؅	:�e3��ҕos>��Z���=0���J]І��a;�/�A��D�.�$u}����댙�l1X)���g��U�o�ࢱi�qM�>_&F���)@4��\���+R����e�-�o�M�r��p�꬜��z]4V�"v��y�0w�A�<k�WX��lfvT����C˼g�_�4�Z)�y�ud���-��1�,�v@�
��(If{6J�����1�Ԝ�+�f�d��1u��P�1���1�Z����R��R���Qh���̙�7�<��A������컘=0�e�����il{+ywO��aVrn��էvm�Ӭ�oSw5���Ѵ���fͶ�:�����P'�vuE�9΄Mŗ��3��a[���	�vE����v;�bsu+����J�+��#X��9���rE��M�n��L�hp m������2�EY���ۦ9s&S��xd�Q�eOmz"7�P9�a�>~�����`��Y�W�v�*(z��x�Ϸ��S0@��t<���g���R-������~�*P�Y��}�Ҫ��'�hz^Z/-���[�j� Ӟܱ���u����
��@^l�o�v��&wę��&&��+C����g�*��yd5�ۤ�rY�CD(&lg�8�ٺ�%3о<
إ��Y�J�y���Ѧ;��Iq�g[���.�9�l��~9f�z<ʃۗ�e{��[	(�T�&O�����*�Æ�[�En1�γI�].��tIi����g�ى{���v�@o)�cc����|=��y{=m�/��ŋNn��A���ŏs�pc�[�d1r�]O0=���;� �[*��*1-�ځ�r��%rh�]/l!�2�i��6��]c*ϑ�_�n��.7�:�	�E٣q>s�+�]���9AyӜmͺ��;�FR�+�^Z����5��Ld�7� �ĺ^���<7)�:;1m�׾�>��nz���
�J�3�N�*�Gr��f���.;�;uE('=��\=\��$��m����de�C��ڑ���>6m�z��k��;�:0���r^rrҍ�R�5�/�w��th�!:�I7[YVTF���&������5z=�^EZ �w;�}���!�H�� �O�̓��o�^k~%����ܩK�Ni��l� ��U��K�����t�C��� r�0Qڌi���W�y~�ͱc�h�������=>.��Ӽg��b=�K����Gm�����~2�'�ɉ��C�z���rP7ǹPaq�X��f:�7��}^��E�[�G)k���Ͳ�=)��w�װ;�P��O4�G����k*�����v�u���:�U�P5|���r8Uw����g)�[��L�ԝ�R���<D�����U��RPr�����P	���L��:��;�y.�I�j-��k��܉��F��C�6D>��Qu_x���:�)L�ʬy��pe�f�Y��,y6c�³7�U��#(��H_b[6YG��;��e�4���L��|o�G��}L笣4���oeoE\Nk������<Xӕ�V�-�IU��9�$��
vP�XvP���h�O��-�z�Od�}*��Of2r�޳���Bٔ��i�j*��q���-�����H+׿XX1!Z�WG�g�bvG�J{�yP���;R� �zA})���7�}�{��ޤ`��]^����{"��z���eT�X'�}�K��a(�����ܙ})\���K*�	��w&��O:�C2�u<<=���}���G�m5�c��a}�Bde}�Z$#�شL�����v3#������W�º�Y��� ��T��jͤ�G{��-1�H�+C��i}�6�s�'�[���jپ�=�}�S�YU6)�{S��֑b�9VuE�qWN�*��u��X�A���̡o���}�g�{�T69�4ƞ�����D08~��b�=j_�.ǈ障�r���=�px]���|�0�r���s��X�������jE>�i��篻�GH�0{������W���3�l�
���#���I�������-a3�oo��K���Q�#��×E��A���?��9��4'��,�S��}�j�/�;7]y^���Q����$h_�Y;AU���E�cLV�/���Wz��[D̓:Ӟ�I���vp��x4z�̚�>�Pt+�r�B�p^%��v*\7Nx^��󲝃P�)��V�N�3�N�V���A�ã�	
�.\و@
:��*ˇ�/�����+�Y�e�����J�	Xc9j>Kˆ�cFA��[�]X��n�ЯE�6{������VL��z������텮CU-]Zxv��¤f2&c�/�P�U�|��74��lE�o�iñX�o�`��Rc�3Q��a7�C�}Ne��6�;�A�ݽ�����g̞+��2�8T4�D��H-���$ ��dL��˴���+����no���H�u�4z;pO>FϷ�U���*ә��Ie���8g]k�U����]y�mٗmZ�2Ex�+qÕw�g�j6y�ﳠ�^<8=[evƊ�\���I�����&IgJ�I�����Ң����Y��:�U`�W��)k���)���<�3@�[ )7��G}Ǘ14e�Zد�Ps�M�Μ�_�q��7�-�K����R��ʗ|��/���6�K�����n�o�d�'=�ǫi�y�����N���[t�f*��VV�be4�@�\ؠ��Tţt�x^�[��y+;N8��wr��g��o��;�q.u*U��U��P��
p��d����0A�1T�x�7�^�k^�I����w�~S��� �ܰ%.���`6W��jN���1=�w�3��$���K;������.�qI�}������$U[R0dKT.2e���'�Z���W�����t t2���=ًGV�5�gnoq�D�$�ۍ��#�Xv5�y8q�]R䈎��w�p���Dd��^�TG_VK��H]ƺ��9�νOq���I�������d-E��9��8��l���O���;^_vP���E^=vv�U�E_oWA��EF��sU�|:�#K�Y;AQ; �{J�,e[�i��kT���g��d��l�+�b/�ns()�`P�Y��ȎƑ���0�f58t�{
Ͻ�I^����!����ъ�R�9��z�$O�)l.���}0 �Ȁ)_=Br�7���6�v0�O�c�{�������.�҆u����~�K��T�0��d�0g�2����ځ}ٳ=9��۝|m�Z������
���t�V�0�Ϯd�~�*�Ϥ���!��#8�6f�q�V|=c��D����1yh��K��/��zΘ&o4K@�s��v��I���EvО戰{���lvSIq�e(zo/�xq��u��ǈ�Q�0uy�d»�{���ްf>�-}�M�$�#$c�媙�{B�V4<~�m&V�
o������{���n�4����y{�x�x�J'��g�|�>�X�mz�V���LLpE��cc��Ǿs�r���K=��Ƿ/���n*�jJ>���驎튴p\v�yv�	�o���Y=X��A\6^Z��02�������N��/��V���n�v����\���$�ɴثj\�gk��9���=��zӳ_���cg�$��"��G�L>�9�G
��� �]�t���q���N
���)n�Щ�#�]�3��Pc�k'��UM�ļ+�>�U������E]�T2ԋ��9�P\�e�5�.^�O��5��\랠n��C2,�|A�z
�h�u\�g�� ��bg�E��ή��Ov`��-�{׬�:�r�P�u�k��!�Fڊ=+E>���F��r%L���g6�3߷���f�'l��e�[�@�)q��jG��Z�:�Y�ߨh�������u��:��sӣI�Qa�}� �"�39=;(�L��D<�$C����'�;��e�1N���G�o�={��b����D��Tx̱���¦�\Y����;:{c"z�H���/WNs�T�
�	C�;^��V��.Śg_d�EC+��QW�H�v�����N���{�h�^�t��^�>Tx�����iَ�����4�b��<��9��	�u�5b���<��՚��d��p5�A�4�-]ga����sA�<ܳ���(t���'��7�]tє1K��Uu�I��X�%}n�OW��;��!�8�S�c4�c1E~��a�V����}��N����~U)�oF��C>I�u�H�!P���
����=�w���q]�pm�{�{�{ʕ(��~���O;�qӤp�n5M�&���n�٧	uf�N��^sG��2��[C[ד�Jg\o[�O�ە�Չ�a����*AoH��9�l�|:�b{C�H���~D)8�f{��^���$��+O�%�?9�VW��#(e�� /��D����������N�<aE�yǖ�vG�&[�!�yu�q9_k����
�X��ʹv��}yj=O�=��&=�*~B�Ep�6���x{+m�2��_
O�*�{1�{��d�7�`�o�w@f���=m�o^K5�z�՘�r��q�p�|D��{�kV<�KԦ��{�|�t3�)[@k&ɝ�j�����9^�Ӥ�r�𤨱^7�R�V��r3<�ϛ�:zc{ܼ�=l=��Ȧ`�WEOMdاu����i�6-C�U�F���q)�v�\��:�z����;y�I�}�н�Txq�����U�����܃�x�aQ�|&�iB�"'�r�۵^��խ�1��7�b��;�5|��2��{*�۳1�6�'�w�������g�,J;e���X�I<&һʯ�`�c!�}��9(�������@��"���b�/��Tͽ��ċ���]K�7:�����F���k6��C�T{��
��+qAG�W;��Q�_MIv�V?yu����>��Rs'UY�4s��6o������v���w���ɝ���ހ�7;ͅCޒ�q�j��N���*t�O�p*ܪ�*��:�<&�kA�[T�h5nz���6h[�l�"7����@�x%���d4��@��#B��v�=l<��ؘY3~Ƙ�+r�.�쓳už��vb0�����;�G�&�O>�Pb�r�B�Vp^%�;�b�c��=�=��Z�Ş��P�7�Y�*�"X;�;�txHV�r���L@0� vx�7ʯ�gIZ�);���Z��6W��q���3�s*����i�D��H-��؀�����\��J|�y��")�Ue���1�����#eoL�%|��V�s1��,���'.�_KU�wo��J��WF�J��gf�*
��n�~~�w��f��|&o�%}�*/��W=w	`��\oZ*��K���,J��ky�lu�jj&�N�=�V�T��x��wZdw�M��̯:P��w�[͵V3�f���uK�=�n�V�ת��0�ç�`t��@+}1��1ɝ�}�جn��-R����{n�s�f���aUOd�~�v[����ǧ=2���U�}s*�<��ǔ�b�����#��T;�`�"����_S�֧��"�*V�Gr�2�����=.�c���=�+y�C}K�M��b�6k��`>�Y1�[��r.t]�G�p�e�ߕ���ɢ��=r�uD0�m�M�;3AÓ2%삐�U­m%(e����wq�`zhL��e���`K/9�Si�Usg+ef�����nyu|�K���=����a�b�.�Pmu����~�Y�����\��Bۮ��Γ�+gւ�����Ϫ�B���m(����p�@l��3��X�d\E���W���ӵ�{��g�)V���!��t8�:Nß_Z����Ԅ��ja���l��>kf�k�����z��U����6iug�5=a�O����D珢+GF�����$u}�0.s/gQ��P.�B.�w��&�2����<�]4V�";)�h|�h5�[�`!�~���:{U��0h����X�mM>3�{F*�I�~���^���Ϧ  _Ls5�y�k���5�w���7���@� �Q��}Y|3�J֧���1�R)�~ڕ��쫸���f>�ߑ�� �̂���Su�*j�QӚi���L���xeh��3[в(�{�r�{��,\&o�ꮠ����{=j�zC�o��&/����0J��}w"����m��?7}�\�Q�ģG{rݵf���[D��Ĳ�0:�[�M������[�L+���!��@R~p����<Z�#��%�9nu�<N��b+EݐxR��k�C�<K]]�h	ָ��r��h]n[u�D޺�7��x4ۘc�F�+�]\�9��o��g^\'2wL�k������]YL���\�Y��c7�x\���lĝ�Ս�uf�K\�T�>n�;ض@q�/+	��n�z�Ƞw��H���I��l+�I<.�*a��6p.�ܭvE[LgJ�e>Lm<Z��҅��}�D@�h�9����S�+�J�-3�}j#��]��+�)�:�BN�O-w�<u3C�=rq�y1Q��y��N���5R:
�����H���7�)�̶��u�V�]��KN��ϋ���Ү�l�yytܚ5��au�k��q���~���Ε��:�{!GP{tf̸`PZ�|^,�ހczjf���AJ�q��g][]�k�/�zi�pp���Êzޞ9�h��Y��y�{'�}�+d[���5w��	�ĹR�AQ��)�o^��+�q��[h�����7u�V�)�7}B�
�v-I�x��v�\�g�z���ۇ������+ـ��d�t����M{���| �g(���9�3 k6R��2�
�T=Z�M��� ���h�E嵖�~Z���3n��(v[6֎yP6�X�-l�%>����5n��x_���g�w�5mXF`�;�c�)������{t�ev?�u[��X�.�l�l|�\��&�0`���Ԏ��[�:&ҜmSt��lb��u-y2M	�7����rn>�Q9�R� ��y�ZU"7�g"'�R|�%o��'t� qեk��#���ed�G�tH�_c$�����+�`v�K�hk4'b����~��+U-�\���70Ve��mp\F�fwcNFao�˒�oyN�Ǔ+�����*��ոe�2%��%�l`�Ϝ,=ڣ����"�{��j��x��m�ų��!�-�eY�?,�
�o-F�1�
���eD�8���C�R��a�~�� *lf�����f�v�5�����;�I���	�}B�L3.�۪�w�v�zcb�x�k��X��=(,�4Py^�=�sF,w��,��[�S�A��x3� Nt�䞅4�d�^tFޝ�ֹ/�h�֕05��oz^VaQo��V�N�U�fg8I�,l���a=/Z�2;�|v�e	NL\��]s�����6:�qz��J.���c�� _��A�!��wgsQ'|���hp���{z2�+�0��@\���tu�,�
�4��TM����&e�TF
��SU_&:��ST�,P"�͙,X�G�7`L����/N�U��p��u�ԖJ%z�u����棭!�S���g�X��QP��  PB�����ZFZ�1�����&Z�1Tb1��V��b���,X��)Q�J���b*�����2QJ���PQb���*̵AU`,DQX��*Ď$̔QF+��TX���
�P�J��(��,Aq�#�b*�TXʔb1Eb�DEUU1����++F*��������Ab"��D`�b��bbV8�rՂ���QDq*9s%UX�1QV(��U���ʔjµPV*e*��T1�Ȋ1Q�UDD`����cDbF�UJ����Z��%��j���*1AH������ƥX�[r�b�Ѫ�l�ˊ�!o��ܭ)]s���bof��s� Y!�pFS]���{�A=���,kռ\���-���թ謨�>]��[7�s�o����~��FL
K>)�T�Ȓ��3�U���6����[/p6�l��nw�Z���W��%�s�>ę��:���j���{��g��"����^�V����r5+�*�}������UkR�	�xFT>@>�X�mz᳕զNT��<Qh9�I�8OUfKL�<(��]q��u*gi�������=驎튴pq���W�]����z��� ޥ�	�_�.K�yA���;���R��J�9ML��&�^�ؘ�ur�W퓌�<�N7|ǹM�TE���^r�ve*|�
��
Dp5� 3U�9ͨ�{]��3�<��GA=�8�4���꞊�*�8P�l���.zV
|�.���s��[��s';�)��B<#�B_ܜ�b�x����Q�4��U��+Q�H��9�u�^�y}�����y��'���U{������c���gJ��<�yQ"P�}�=���=ߧ��X+��gɥ]�_<d�A�'<���z�N�y}}{�J�{8`�	�C+�pu��d1���N��.A�X��gx�f,;���CZ/�$�Ͻ�N��Q�f�޹���]�Y˧��n�z��hvC^I=Z����n��a
��IJa��]�,t���Ѵ�|M"�4�3ݥ���;������=r��k�Tz�5}1��/���V��y˺�OgACJ���JӬ���F.SՂ�� |%5f���	WlFM+Ը]4xw�C����.��øo	A'�zS����t���v�Ջf#�*駈оvC$�[�Pr��@4x�CYW��s+�M�\�w<XmV�p�Pi1��Q�C��#K^I�+|��7�ՄXCu0+{Wx����Y�LJr��Ͻ�X�#�-2T�ޑ�.��.�@��,Oh{h_&����j������W��~^<�PU���8�:)v�ʲ��e�tH-�9]��a��,8v���ifם��{4q��C֝#�Y��q��w*���ԅ��g@���+��e�4���+��� �ݓ��K�bTȘ6n���s����G:��O��-�z�T�K�����˨[��g�i����`�s��Ġ�y�R�ذ�ße�hu���˕�[\2����Uq����(]�9������}����d^[�(A2J�X%��BV�X��Gvk�ru)oџ�x�1Qp5�%��wo��ަv�J�/�G�O��E{��[�~�Q�z#�\P�%]�]� �������N|�T�͞��]��G�)�ua���ts �j�g��u�[������8�{���[ݏ*N�D^1{/�a����e3{/3eķ9�Er����	���Ʀ`ޗOƜاu�����֑͋P��i0���oŽ�냶{/*��6-�I'��zB�8yP�3�4�=N�Go�\��U��X}w���n�^��O���)_4�#����o(��1E�L�a�5C�s��]?VRqw�~��q߫�o��:�*�ʼ ��88]�����60��>�C2>���MV��y�:����Q�綕AJ��U��<UdwÃ�n�V4�ϭ�~5��Ͱ��^ֽ����}�.���
�Tf��}�]�i�.�ʢF��œ�ǭ��WV�Yl�=؋��=�P}.��[�K��;dY����ϛ��(Nw�G�L��ÁP�;�B���߰N`L�<��fr�s��!�x.�59�Z�Ffxu3���e(�ܘ�a|�h���[���Nf�c��^�`ʳ���IS��γ�3y�X��i����ZX`�ug��-��TǷ�r��y��7�Ȧ+�Ϭ��]�=���>F�ޙVJ�˂�|�OU������NU�n��ȔV�Ⱦ7-���.ƈO���_\}�Z��j��5C��v��@9�OV�c+��͌E@.��Mأ1�Ӷ��K��Z������(f����Wv���$�7:�q���8_JQWzb�ȥ�\�Y�`���7�qιӜBp�{5���^֍�M@T�6�އ�U�U��1�o#iTq�4y�^-r̼U��	������w;�_ӚŞn��LDա���L��K\b��s��%�e��
��M���t�-S� ���z����ʦo��Ҷ�*�1zi�:�Y��rӃ�����S�,��شL��h�{�uV��K�����Y���׳(�����OR�{��l���V*��u%(`����LGw��f�&�o�-���b�cz�Bu_�w��:�Z�w���cJ�c��}Z�(�>#���U돰��t�#������ȱ���
�&n5��x}ʀm�2^�	:+Y=�.��-�3������VT�y�3�����HD�W�@z�y��z$w!#NVK���C6l� �-ױ�0V)|ɞ�6åj�W��[(�ڙX	rX�K"�������	5�:o��;�_��*����_��}�M���b��Y��;�%4w�@��X!ݕMl��{z͸���T��Y���4���+�*S-J˽�H׽��w�¢���I+W��y�5�`���M�a6�݁(6�q��W>CG.�x��[�� =v��Һ)S�`᝘ܖ��vI��[�:Lk��>?m��{z��ɱۗ��]�D�ee'��m���g���Z)|�?y}�'⽑1�1��z��nTi���s���r �{���s�Fa�y����/��x{B�7��m�Z�8M���`oO�X{�#7���5�8���gJݺa×2e;����	�F̕7:�i=��jƙ|ו��𚧂����Ȏ���N�ᮋ����:`�!F���S����śdϰ���A���#DX>��^���m4�RQa��%Ly�a5_nCy���x���M/o5`�� �j2Ԃ�TvG��UE�
�+�ni�U�)o��r>ŵ�9d4�=���GȾ.kR�	�xFC����^�]A�VGڧ9޳碞�2_m?L\�5�¶�d�[�4p��H���{��s=�u1��Nk�}�����N�p�x�p�ia����J���}�({r�T��ԩÍL��F���'[��g��>&f�c��u�Ѷ`�,�֕�C)r�]N`'�ȍ}}�0��S���݌k������,,� �]�+F�:�{8>�бk��n��9[��k����^�"~�}���ce3��w%��=�֓]Gsq�9�u�0"!�ԃ�5�t��!�؂��p���q�vlűX�u�u�M̫�a�y`�gUÉ���~���{��Ujk)�-���p�yU�ɳ�V
\H�}k����z\��l�7��m˼��bFo"T.z�o�����&�V�K��^Z��i����,�C���o_��g)���gO���:0Oz $ȫDN�c�*��L�}!��>�ͳʅ�
?s��t B�M�I�]�|�V*<fX�D��*oPeśN@��S�N�5��,�:�|�=Gt��a �ڏ�/���Q�4��ǧ�]���~��g�o8V�����;xA�q�x�^�)ܥ�S@��՚Ʉ�����ic����(k�G�_���˽:�/$�wt��^�+�����*�՚��d�`k~J^�謫�?:���{��7���[5�|���b���I���Xz8Da	c�� ���^��9"�;k�}k�߻^��ç^x�W�m:��fPR�=@��Dԅ�#Q�qK�P*x�^��V��6Ϗfz=iP||���>oE/��<n�ڴT��)U�<�B"�*�[�s�N_S���CLY}�#N�i�7��&,��}oC���Z^���4zG�i�Q�q�R����
5̒b�����7�Q�[�~!$�*&�_��q��'ۯ�T���c��Pץ�e��c�4�<U��O |o̞j,�b�����$6�<y���l�l�L9�i<cG���KV����eś�PժO��]ʸ���ԅf�K:=��0�"r�t�;�㡞�G���c�?�oҊ�2��/��m������N��[+<44zdڈ����*�0���[�k
�������'���t&@��t�p�q���.�{[|D�š��$+r������gqڞ��L�F�p���b�F���b�75��t���a�chO�؜�����ӛ�7*�#�Ũt��罒�_[��f��"�"B)��p5}V�9����8��qW�}^�==�=�:�r��w�VOv�]������!|-�K�1�{����yD�/��*�H@��`�w3Xv�8;3q+��}陜<,gN�xۢ��KQ���"�ޘ�#l=�qC����#]Py���w�vV>�=��M�>�\)}Z�*�i*��:�<&�kA�[T�hi�/Y̱�,OW��3j�=r�A������qP�E}�����\Y;A�S�
�O;7z
�R�����N��ݻ�ת#��ȹ���׹/��bG�k紩�ڭ��Uz�n��|��5�,s�Z�[Ds�R$.T	��_)J,K�z�u ���ޣ"�1����\`
]I�Lγ�r:vn�YR�AڜM��q��][���V�Y̏��+�����^U�;*���';��H�z=����0Ag��M��nM����Uհ�`߱�|k9��R���ǜ��̋؋��%x�9�I֝�>�۷��
��xH�q*�}���gYӛ�U�
f�|"OO���]Oupgp5��Z��ue��S;����/�»	lW���/,ϑ�7�-!����f�r��6����x/v/���9+ކ��jԡ��Dq�+_o�׵E&U�SG���bAy�G�6U�Rd\����Y3��V��tI~gR��b�7��թCY7�yst�x���Q��	���KI�Nݘ�;�yM>�Y���K���$�)�����6��f�1�iͤܘ��!N��4���|����PѨ�}��W+��4=�h�����aOd�j����~�N�C�)o}��
*�Y���V����]I:C��+>���ϚS� ~3�دV�̜D�x>��-�^�>�^}�_����PnK a�hc��լ��:�~��U��,|6j�AU�ߟD��s���t7)����41#=�ƺ�̖�X)
xs4��Y����п{
�ZzJ�s�0gί�Z���+x�ܻ:rIM�X�U���^�&��^�*��y���i���������*J��y͵p�u�=������n���9rE��,A��ʂ�>�U�e�z9I-^@]=�������q����� ؽ�怇;��1-��Q��C�ӉP҉�s�Z���+G/$;/��`T-�#_k���w=/x�:U��ʯ;!Rm�J�F��j�6Y��	���Kh�ͽ}OޓdÏZ��y�xt�_�c*�SO�򂽲��&�2��s��M�ȎƑ�W�:�uK�����H��d�[@�Mnb�`�mM>�<�|Ƕ���ޜ�ڣ�o!��z��Qr��%b���f����`�&� �P>F����s�Fa�w�^�Nݡʝ���׀�#����>����Ԭy�Tʸ"��e���b�������gJݺa��1�8�������76�J�)�11A(8|%4��cG�S�Hiq�QC����(v���cƜ�b�9�e�5��R(a���{��"��]��/��\��=�Ӭi�=��������tޤ&��lz�v��7��WϦl�d�
�O}9�}�Ľ�+C���w�WwHp��Gi�cKb���[, E�����L���+f�]�fԕ���i�n��b�z��Ug'c3F�J�%9]��;1%�,�&�h2����PP�ju7q'�y�-�I���dəw�F�|k�s���X�Uv�쇠͐�4��XᛇRqz �j�ݧ�*�j�gQ�3��x�J*���`�'܈�<�Yާmo_c�6󖽦$){�bc@�>?S��ZS&����#��R���t=���r�8�)��qɶ��:LX;=ΰhу�\����+�"\0�=p,}�({r�T�ԩ��>Ȥ���=y�kt1��}Fq����/6�o|pW��e��%c��\����>�S|��n���[60wÀgC�ET�3bȲԮb�k��>H�R�{J���9����7Wrf�@���$h^��*�8C�P��S��,M.�P0񉵪����k͡���-5�	��$�^|��x���JPaV*�����dC49ͮհ+��/��x���-���+���"ģ��Lȑ\�˱�����Tx̰2Q0�Tޠˋ6�y\�og=�Nv�S+���N���ީD,�,�
��4k�M?_Lz|[�]�M��ꐭ9�v�j��
��zj��Z�{���AV���|����p���~gHIO���$���$��BH@�RB���$�܄��$��B���$��!$ I?섐�$��B����$�!$ I)	!I�BH@�bB���$�؄��$��$�	'�!$ I?�B��B���(+$�k;�����0
 ��d��Io|w��DE*I%%BB�)(�Q%TQBIT�*�J��!HD��T��IQ%J�*����$
%
�������T���[����**�ъIIQDU!�*��J�-�M��*
����UP�*���HU@��hJ@J�$�	IBD��U*�*-���DU("��I��
���)%��l�%ElR*T�R
����i(QD��  tx ,0 �l�Ҷ���H�MA��6�R�Ul
�4MZ�h �f�i�AK)*@��"R���J^   w^j��ͳll�`YVű��l�Ҕ��,��@,-�MY�*� -`U�m���
��M�3E���]&�"�E ��B;�  ��t4(P�E��B�P�hP�C�;���
P�BΦ�@  P�C�.��СB��
�w
(P�C@ �W8P�(P�C��*�R�]����`���X,�k
�5Tld�UZ�S�  ����Ц��akP�m�e���ea�X�H�1m�Ɔ�P��4ʁ���+T���1�P�6F-`6���Z���("����  �^l�V�j	�4hқ$�+CY���P�3Z��R�ؙ�4��5F�4�,��-���� ֭�� m�Sa)J�*����+l��  �ƀU�Ki�M�ki+jضU
Z��5M(�a� �&�hi��hձl)0l�-�؛T�Th�b���CJ�I"
���IET�=�  w�6�(�f`��Tm*�kESB���`Sl�m[m�m �-�iCD�i�f�YYm�4��0���̫m��-��Ғ�֨��J�U	�  r�S[0Z�ZVC �i0���@�Z5Fj, fKP��a�Z +$! �D�"�Q.  �E 1� U[m��6)�P �cZР�0 �0 �	�F�U��-���Ī����EEAI
�  � V�� j`��E *�a�h����
�1TR�l �b� 3� jcA�%J�� E=�	)J�  ~���  O��Dh  ��R� �L�	5�U)� ��[�0���Ez�N�y��La̠P���nY��?o��\�v���IO�ܟȄ��$�$ �	!I����$��$�	#!���s�y�~_��0��UCx��@�Iٹ��ul�KBr��i���b�Yc	T��d����g0�n���\�q[�r��f�I�B*��|��i�9�ŧ�"�R�H�b�l�Cm]���&��Ґ��`��K��F@t^�m�[��ՙnZ��(���ś�r��6̷f��b1 �r���%i�%�W5c�<v;�!m�ڰ�A���5/Ml�$h�-n�߮E�$ئ\���M�ƪ� dS��ۻ��-��i�K�����#3ka��M�ݎ���B����5e�;9�*7�xp�У���%fG���2�j�0�v�Ц5Kn�ђ�`3-S:�P,�`P�J�{mۛ����Ъzq��Csn�w�W��jf<[����wό0AN��ָ�.kt�˻�D��fVæVTщ���mB���u'�cD��Z/te��"�G c�[l;n�������Zqf#�kN���c��T�7��T��ʹ�*��YP��Ɏ�.���-�6(r�
�z2md �	�hYx����6�5��ƕ�m��b`C4=M ���^���ً�R�f��e�L�(��^!`��n6�V2�LP�E�.�)��.S[+N*E�@2�(���押�%��ˢǘ�`-")ɨ������ó��m�.�,V�����|)Ȓ�a��7��5  pE��k2,����53_l�a�s4[�{P�w�X��Z��](ДJk!NV�Oaj"Y�&\�(7[X2��&����`Vm�T��b9��	��е�n��D6� �*�;���b���N񝺼�����H"�6�����������.�>�q��O�w���2�k�N��XDK�j[n`�wWX���[��M�*Jr�� Z�l�z.jx�mV�X�Vlz
/B��N�p�Gh�{@)�F�V76{�&!hka��S6헥�1�Ma�sr�[�h���u��7���[ji:��%ܩt]0������ɲ����z.�+U��R5s��X��A�5g�XoQ
��B�ʧn�����dͬmZ�5���n��I�j�^yYbX{b���j����P�4I1X���X���`e���1<�(��ki��)S#!��}�dlʥqܦ��%滇q0@�S���I=�i�<�a�R,���wSM��ݺʆD�_&�K	&U�ym��sM0�� H�w��v�P՚�0*�����v�к�����b��b��(I�V��U/ ��/!�@�	�61���������O):�m�ᗪ$�v�<�G
�@���Q2�`�h��{���X��޲��B�/^:"�t̡�A�Qy��(�W�����)�� �-%��cѕ�meZO$H��J�gw>�2�e���6�� �T���бF�J��W���	�hz��QL���g�V!DdF�D@)�LG�G�R�1�<�R-�qQ�����MXM�����L)},����>յ*37m�;��(:�=�7EZ��1�[,�tV͑@��-��\�F8v��9m�L�7�!Zȹ���$u7ve4�����fV���h�5�t-������
�+Xy�G
�Q�"1�m�<t+qY`m�v��\4� n���0�3d�h�|�����b����ՁOq+�eb)�m��y.n��WB��2��
u4 ��X�cZ� ���$���ۺ��Iq3,% �Iiu��;WrfJ�kd��N��R�v�ύ_pm�r���ڡ ����(��)W�;��t�H�{1�31��dۗy���Զѵ5a�'#�	XqW�h�3,�!OҦ�w3�P�S]fV��r�3�c�dR�-�<�*�S*eF�h[Ҭ��{��%� a,4��7�jaks6��	m�����̽��
b�Q#Q��굓2m�HfX�ђä0�LBƙ7KKI���-�K�ڔb�9�0a�"K�E�h������Ḱ�!Uva&��#H��mE�ԚF�na�xMs�EY�����K��Pm���g4(�E����N��i�R�{��Cx1^"^��q3r<�70fMr�Ci�P0�Զ���Lr�Ur9xŅZ��V��ɍ0l������L�&�)[36��˼1��"�,�Wr����6��x˺N]jOr���i����R�7t.� ����z��v��L��*z�奈�ڻR��"8����[�ע���bA��ϯC	�wi�VIi�#��B���I���׮��6��0�W抺pݐ�ԩE��[��RM�t�:zo��wV����i���C�KKJM�h�52���)SѠ������k�F]'v3���e�ݰ�f^�ՂSX-\d9�c��8%˼kr1�H"��GB�m��Ԩ"����P*׍��j��"Z̺�c-���d�̼����8�EP(�d��vQ��RfůE#��ɺ�H���e�y�VCB�	ɳaV��T����1q�
�^��y���vf�4��  ��C{6��39o��4ꕸ.}7A{�*L?nEc0��*��1]v�+�us�-*m�74e�_K���L��u#h��Nb$���(�Z(<�6�pU����-�xv�DtڷE���Kͨ,�Ús]�fKv�P�v�V� �VցWa�%��bXFn����L�e��7���e��B�����B�V8lٛ2�Xl��b"�*Vt���+���ZԖ���h��T��-�q*�d�����z��3bڍKB�46��J��"�)���Qb�d����P�E�Y�fnJ4�;o)ݦ�u�ŃM�4���w5�R��5���߃ʳ
4 j�,�7R<
^�I��Lj�	�u�.J�YKfc�[�Q{���CAmӗX�%lݲ2}qQ�&�
�D���V��m�#2
іST�V�ʁ�,�# �^�,��em��]����/(�!�3y�e:&��r!X��1��9�e����L A'�ǊŪ���j�ڊl!���gG�yA�Xr��`.��Q�]�Y�ݼY)5ej�S@r�^m�p˰�'�%�'x�4��vA�ٵ��bkm�3�j&�\���wEB����4��)V�V�+g> ���P����ћ�p�&�ئ��� ˦2PV�l+`�~WK�3\m��;	�%�44�P��Щ��OD⸊F�+SA1R�ѳ�"�;E�k�	�v,�e2Q�M�2�
�	�;F�Nh�FkȪ���!FVe�x�wOq�r�GR5� ��-bK)�� ��>Y����Db���⫗���9[l8Da*0]�Jګ���f5�mGj��ub�U���)VТ�Q0� t�f)�hd��	���ȥ=��iF2�#p-#D��
�Ui<����n����_ւ�$l7�x@���%nD��V�ܰ�G3,d{n�\Z�U%��7
��b\�*��s��B�Y�e��Y��
qQ��8��*��E呟4�����@M��fX�@��ݣ�E��*-:�%�v�ǵ�K�gB7+f��wb�\��E�% U��]���1]�`��Ր�p5��*Ɇ�u��F��- ^*��恚A`\�N�V�@n[ ��%n����D&�-BRx�懐��5�MY�3U�N�KM�u��$����pkaݡ*Vu1�B�`�@�KoVՉ{`�*����ME�����Ӛƌ������ܫY�z� J�!kǰ17�����1���[ӗ�^�t�&�j�z�ٹ4R����+lq�8�P��^kY�2��9l�j<DL�gZ�Y�A���[h��ƀ���e�v���XF@� 7����U�J��BP���Y*�R��yKoL�z����n�֦7@�[� ��q �(.��V��[���Z�Kv�D45��D�vs)bP<7 :��xwR҅������[����1R���6�7���2)��Vm*�����ضT��b�ء.8�c�V�ɗy�F+P[��D&�j�q�R�˫��vq�hp�p�@ɳCn�|���ND1�{�j��Pl�+%�ŪBT �B�	W&
�$�53R�oV�%F�F[���jf�K Ф����nPiPZp�,ثZ�zu=1��O��
�n@�4dr��V/LA�	��/(��3��U�-�I�,!R�n��kYi#T���sg�Ihlk3���A�����a�&ő!�b�+E�Z>_+�9nri�A��'�Mʛ�d.H��T�j�m�A�r�ƛԩ�+&�\˫�I��4���b�7ҥ�W��n�5���z�T�c�E(��{�m�1��-�oq�j�c�s��ܘ�m�%�n�)�z��*Mh���Z���D"�wH��C�6-���P
h�n�\LjtjmI%�f�<I�on��2�اY)�i��Fˁ�`��X�M�x��Y �ܙ�i�+n�(*),␱��T�h��V�32�=��R��%�8�t�V��50P֊L,� ٶ[��h˱�Tܬ-fSr����F^�"X���*��6�) ��c̩31�tf�i���R�kn'��Ke�ȪҎRTv��dV�ݤr��#�d6�c�Ӥ�7�N�S�+&e	%����
Ub�҃��E����DL�"�!�x��˽�R�ĥ؆�j�q�_B�k��n�cM#���6��0�X�
!mOlvӭ�L�ŪR��L5Ck��{%갩�%5B��E���B�'Y��jM�E�n(Q �r�۵@�*P���IU�)V��ܗ�j��j�Xi
N�Tܻ��u��S��@hu�1�[�E�Me�,�,�fJ����Eѫ&ۘ�Ia֢���S��퉻$��5Ϟi8����*�[�����j�+�H���E`���&-��5�)V����^*�X��E8�Ĳ,Wb�a�ӤT�. )�n�� �ډ���#P�0�f��t�yy�[��E����545RQ�c ��Ya�7~��Ĭ�*���a!�X*{hfK�����%��Y�ފչ��Z1H��b�ʒ���a�J��9�h2�#�����aޔ&��˫�u�6�@A,.����NU�* �ImՏ��/Mz��>8��N�]���#���J��B���F�e0�����ɡ,���w���՜so�0ҍM�ͺ���	W!��c��^�����bv���z�[�)�@e+r'�6�Inn\�wLցX�0�oV�V^�B03��m���J��Hf�?9cN���`,�&JZ�,�@3�=�`H�U��L��bJ�J�m p+t��X�Q%����F�V7u�8��o�R���R]��x1^�B@´e�{���#�ؗN�7M�����S.�Փ)�)�-�T�n�Melh�ch-C\�$َX1
7�)L�fwu��R�5�;{S�d�0�e%���5yn�]c���\�wf�Cr�m��TY��1	���6���O���=c`Ò��m4�G`�[��N�v]GY�uu����#D�����$��`l̓Vի�gM	��բ`�|v
�0��LemX���V���Iw�S�.m�%��A�F�OoF�&�,#Jn4N`�(:	݄�-sESgZ�V9�+�&��$	'��Bf^+S[p�ԩG)�:��{vá[rعwn���+I7��J٩Xq�6e�����,b^�a�yjU'	b�Om�9�z�s	J�9w��۷H=�4�b������S�a���]��r�8n�5��Ͱ���X-�[��X]��J�Y�Vv�d5t@�+%���V!&}���
�Ur `D�q\��Źp�v�L�-���&^��-3yVV�l�η���r��j����l��(|����nUз�U��!%M�ۣ�'Z�e-��5P`�.�S�fX�k��	zksn�u�/ ���
�V6���Y���^�y��9�,VL�7e"'zZ$`�5h4f&ӻ��ڳ)
�wZ*Ե)�����/0nD�k#�ѕ�v�/Mi�*)�j���Y�7I��W���Z�W�9����E%�u�ں�y�0�6��v����֤j0��.����Y���V`*�̊�}���>8e+8j����V�' ISJ)���n:w�Sv�F����4Z k)#b;-��1��P�1��m�xVJCi� �:�ɮl�u;���V`�5k+��ee�r�Bf��,�Qnan%)�l̊��5aT�6��j@��̤��m�Ab�#�)�O؍*����,S�0ƪ0� ]�I-B?��Yz�,	�@AX�9l`��kJLF�ӮG����*�����ք�5�&����yL��w���k+J!m��E�
���Q����B�A<�R��[l�`�3r�5+���*Ф@5n=O(�)+IV11��J�1J
/$i;�W�C�w�'���&��5e��Z�!@ZB���sU�7b�������B�HuVi[{B�:�E��O悼NXs1�lK$�w3qb�Q��v0��vJH�lg�޳EOc*�j�ɿB�cJ��P�:�1:צL��!Zn��r�nmB��L�E�r�")���Y,��3rTX(]��Qw��'ORx5Xgi,�QP6�X����6Z�7�����D�zc9u���p��1�U^�V�<�*�+ϡ�X�'{��(��]g\��Sa�c"9L�Ur�֭5.��Q)"��ф������j
����,q�An9ut��v��^�Ң��)Pяp�Z`��̴�J��;��R�Bun�+[ځ�q�۔,L�!�y#�Ge�t[�و\�+0�_9�%LJ/�������gP��/V��k��w�q�wA��b�^�u�ת�6���X�$��s�n%�� ��k�,[Y%\�&�1�K��yu�o�J�X�0�����[��K�cLL�i
�4W�Ss��t-ʱht8�i5!�����u����p���j��k�6qu�_&
�u���i�Εv�CYżr���Ǹ�4(؛e�냡�;t��\6p�,q��q�Ә��d���gL�޸����W�_BUv��gE%فµ+�F+ND���//�<���lmoi��8rb��Zm�����F��5��,��¨a\�AWb�]ӕ�R�%�[}|�oO�M�ٌFtK�n��ɟvU�=oq��*V	�E W3Zܦs{KY�=�A���'�o3c[�jy�ٝ�@S��%r��(�^(+qv�k�U�i�:��!�7�_r�
w�2K���<��R��!�6ᆥ�V����=��n!���q�F�|�PT�*uc����gQ=V�h����/���ʎ'�]�\�� �f��g	�5�/��o�����w:tb����[�֩:��&�Yc�\x�Mõ��om)��ƹ5 �;��򵈇]�e�����;8�vU��N����Z:����<-u>�%�+�8��X���`U�3gBV�}��{v��c�w��4� ��Nok�m��&q����<���X��7B����L��f�6���
���L>�G;��MT4�����q+�Ծ�uǤ�x;'�A@F��#4c�o/L�ؖ	�hıg,��koh���ΐ�`4fM�'�7�}�-������y;Jy�d<760	���s��Z�]δ��{�ӡ��t�hR�]ri��Q��p�t��#�z�S�'-�6Um�}�̕�s�*Å����ZZA7X�6����.���w�h����ht[�K��;��X/�䝍��C�&�.�ڐnWAk[��E��OM�Z/&i!=r��B�:Ccb\�=,�5�6�����B�kN\��6v�����a0�s����U���;��3u�.(��Y�)D���Z"$�m۽���M~�SF�K��{\Η��K���X��k��&�xu�vc��D��-5�*d���7:��:�c �0t趕��zmp�u)6��huǒ�>>8f�n\��S"�c�
؍fw>����+GQO��S�b�ƺVے$�4�ٺˠ
q�!.��6U��ؠ��-�IKv���]m������L�:f�6U���wFq��w.V#��V�Gh����w�.5n�f�[�jiu	v�ٱ�y������rC���x��d�3�+3f
ބp`@�Ճ�*���&��MpH4[fS����&��}+*ɴ���ǣ��6]��;�y�ª6��aV�����L�Ȩ���Re�mP������N��U0VV��|��U��F:K���c�TQ5{{����\�ȚD"j×��)ϭ[e/]��o�&�u�ǚ
��͌x2����J�v��f��zhǙ�*�NU{��Ҏ5Y.��b�K
Se���|��'����l��b�P���1R�y}w��s��V�U|�W����v
�[�{�Қ� �vq��t/i!eЕ�F�c�u��}
e]��%w0��L�Ű���nw�%��U�oV�ϧX���W!{�st��2�*�� .XMա&=�jvb���|�U�+E�$��3�hV����(�J��sHU�;(�9�	M�xv�o+uvu�)P�̪1Ņ��ok�Z��vT��P,�Mp�f]`��W�8f�B�b`��=顖�]��d!w���ې;��5��x0���-�wKvb�Γ�<��5/5s����H�.�w����G,���G��X��6���muSc}]V�Ϝ:J�b��w�vk�tN��ڏm�1��Ŵ��ҹJk��N�of���4�.�c�Á�$|U�A�n'�����5�-&<���ta�˩g�V.�	`�U�ዤ�>��|��}:mZG���n�:�>�����N�cC���r��gA������md�"���V-�R�nwg^pwmȋ{���H�7v�����J�ɩLš'{h���>sBem����I�i.�1q[�Ҿ�7)�U��a�R��90*�r���e�u���&̮�F���fv�PpZ�'VQ���Өɫr�ج���
�Q�T�nT��سJQ�� }���#=�A�ڠ�k�h�a)g������u�n����mi��I�u��!��{��p��M�3��k5n���:���[һ��&�J+��n���d��z)���\�}���9�UЃ���y��r�X�:;3��	t�j�\�]�lȳp�Ԯ�k�]# �%wn�c�f�܂g�����\w���׸�V'w��@�3,�3s+������P�ڗ��(wi|���%,\)	mݪ�Rq����^������[4��e52��ܚ(VD\�Fp��놻�֊R@j��yi�n�>���a�gK��T��ʕ��}utm��&K���α�T��jn�G��W$2��Rm�h�R��uv�K�T����2�ٙ��_J�1�wK��/Q9x��'v*�����kL�"�2�_����4m4������Np�;9E�fV�� �7s[#N�p�V	��;О�K��V�X�W+U�� �-�yw� �3UͨtN�z+�4'ق�F7v��w������`	s�;c4Ǻ�x>�V5�F�������q1��J9�����{C��f��S	U�o3�*Zdq��x�q�-ݫa�
P�6��̳�9�%q!���}�tp�9Jx��n�h�E�a}���}�6�=]�x2�u`9g�!�R��s�j��N�7�ah}�_
�u��m�c�Ʒ,$;�V���V���R�"��E��z�RΝۺ.�1�\d)��dD+���L��=udT���j����՝��n�՝���2���i���S��un���bo1��W��g����m�gz��`�
n�E����B�3�ɲ��X�O
��|7��iU��)��J�-�_�uvxX�]�
��C;@�{|VP�aݩ�]�����p0��ؙYu�º����Jy���γ)>���v1�m��P�8���֜6����e	(<��{I۾�<��>\��]t��3+�ܙb�('�����x�(��Z���vV����Xy�EE1�X��X(�G�f�v��Xh�6�w`.�'G}]�œ6��i�b���4�k�MyD��f��;bek���WAs��9wJ�ԃ�{]����3����
�;���}�
J��A]��ۅ�t����v���TŖ�)K�m����Ӻ�sqҕ��_,;�]�	]�&�n��B�О�G��α��i
��o<C���).|�3\q��>�`�,�+MNāJ�_'��Eu�,�p�v��:�'���F��r�Ϋ&�O�;�`Oj����c=jk;S�+�*��B�C{ �jG%tޫՋ��n�%��'J��NI|�%�ij:5�l�\�����Iy��^���ݒV]fҨ�(�T�L8��Wڊ�V����q���O���gӇHl:Z�.'	�d�U��.��f.0�}K��E�֦�������-�D����:���sM-��*�.p.,�ǖmW���2��'�#{Z�����ne�Dc��Wn��ճ�8��,}K1p��+�#�UKfn�[���tY�Y\�L�o42�\+c�:��:U�
��늈Ӗ1�i��ݳ�ĝ�>Ἇ0���f���}[ŕO�����C
�a��eV:ut��ܝ@!�޽*���(�GH��A����.�]�N-5�:��t�����ގ"_	˺�Sk�B�ٶ%쇷6�=�b�8'7�$`t�p��E`|
�������Wha `5}54�-%�A˵���[��=Z{r�9�(����R�.��3�E)�-�"�g/l��*%Gm���\���%g1�el�m�k�1���E���n��-�c����]Ի:�N殧aYHޑ4tY�C�k*AKx�|�����S�k��6�J�����m �w�	�z��u��yq���=�T���^m�������(d��Y�@wQ�eÝ�X�ֺ�u�]|�ĵсd�r�q<���ՙ9�'η�{��������mq(ѝ���g��C,\��J�`W6��͆�v0�RR�1Ss��{d�W��<R��ů�[c9�Cc
��u���ms�<��U�s�iK�C�^��Cba!�͊.�2�eB��"E'YA��X���c�ح����w�a�M��UaN�a�/n���Y/!hƖ���)���f���r�UɎ��s���t;�T�L�W�%褺L�p�*Vr��-�+���c�-�s
��ax��Y���7Av��@٦1i�6�cX)ek�	�;tV�M���j��yy�OB���֊=fל�,-^��8�oy\�b�r��^yc�>h�����Դ��:�<�\6]U��[�0<������Z������:Tp���chocsa�����0��n�C��DZК��G%�M��+B���W^�Q�W�����G�q�|�V���F���R䡄Ԩ�F^n�oW1}�F��1>�j�'��L�wzea�ɡ �2�]��}�]X����͕wY;x���J��i+6�x��+�w]3c���K���8d%��>r��e/5�o*�u@T�n�N3�m�ŉRWV�*���i�i����I�@�}�G(NL�,�<�RoMͩ(j���i��[u,�Y(q�MD�T��8�1��F�U�k^I�ۘk���ٙ��i	Z��t�$�!jD�Ϋ��7Z�����Z��3
y\&c8�]jr�����Rc�����K6�R�o@�:#:�Wm�!��ӛ	��k���]E��^
��um�1]�Z(�oYR�Y-�[�+(��*��Z�ث�>��D9�gq(�2�.��fa���E�d�.C�t���;�<�V�Q���=Lo��v�iK�����m��Q���b�#Ӷ��3Є�r�4�v�V"����U��a���>��nv+������e�`�����T������V���B����%�6�{L�����}��q�`A�����$0�x���͗rR���W�kqN��K�b\i.���lx�����Pj��\���j�� �c7�0}˗K��;�JS/3M�=�sy���̦��cƕ��4qw�P=J|W.q���3r c����rjl�U�;{�Z�@KV^�j�*���K��B��9m��<�ׂ6�$�Ƥį��s}�VqԷ�xk;��tX�� E����k��a�)�T����+��rjȵ�vf�>[|��>�Vs"�������@:Ane]Jѻ�!�.�X��4�Xn��ս�'g86�n��n����6tR8�+7�28	Y˺�[B�8{��eIF�sz+v�z6,3���*,�,�z�_[]�:�c�dܛpIy��l
�w��3Վ�g�L�[��d���[�1ø�cUb=F��7��_L��:I�O��oNµ(�#w9,���=8Ԟk�ggj�+�����w^���B��Lǽx��Y`d%Ҕ�� �}sF��3���:��q����hml�FC\��k��{R7����']L���H�Ӷ�f���2=�"�b��zN3MaÉp����o����Hn�\V�cOh^��y�N�#��k���E�%l���n����]��F�Nl��^֨��΢��g#強rE��ee���@��aވ\CE�]��1�n�Q[��Zk.�8��W���=j��F��������Ƀ!�E@qeFC�*_E��)��F�]��^8�k���NM̓GCu��m��Qo�ZoD.����u���(��.>��3Pf.ɯR�7.K�>�|�r7K&�*-�BC��J��0��x��R�WMR�U��vlZ�a�j+�U*����v����j�3Gv�E�{23����*�-9���N�f�Ȉ3�iڱc�����u�ѫˠp4h�ᕋ:1�`
��� ]Qs�Q�`�8��XV���Ä�&���òw�Z�i����u͢聏2�6%�܈&�Vq��P��mZ)�x�q�V	<�U��"�E��s��1q�M􆔷fn:��}W� "�B�3�u�D��+^m��.�\�4Km"&K'��]8��R��ᬮ���%���N9g*��#�����>�u��r�8��{ֻR�R���
�|s{����{mD9�3���-0�ૻ8�}o:l'ӱtI�60��FV�@����qe�f���F8�6�d}�)��A�N��IbL�n����[	��q[��><�Ң�<Oo���G,�O8����N"�=WY���F�ҏ(�5ǕfY����j�S� ��D�;/��I�x��V�e���݄�x7����]IWi$CfL��᎕�5.��κ�6�ǜ�,����G��[�JW&F��&扐k�Z�+��o��.��K�vp�g,
��
�U�2�hk�qW&�vGN՚�7,�"��nH����sޙuHYZj�Kur-��S��&x�w��5g��MXyESS+&Uԝ��9�Zy4";�5�B�9����X�gK���}��<�)mH3�Ya.��G�3�П��w`��9'-����'|6���o9!f�`'����:�����VK��<;j!�*����Z����
7�6Z��R�[K����h��������Gyvޥ��C5C�Xtv��9kx`�{S�e��b�guu+ޗ9�P�G�]uo)�Dvc����k�y�*���dS�2����;���,��LN��ɡTsRI$��Z��ŉ��<< ���?x{��{�c��E�+��;鹊ʞ=Ct�UFfCh �6�6�@�79i3pSN6�K�!)#�ݱ}��f�좟9l>�W�'�Z��0�H*�@0DnL��	�_.GF]�cN��܆���ٺ4.�mmN�YA�UcE�ɧ�#�Z/p����VS�64+}�i��M�W]>��X��0���et'��j�(i@,gZZ#�W ������gVͭ�[a*���V���]P��su����
�)c]����'�.����NA����S� �v���v��Zh�cu>�T�j��&k�@SG+���;9q��.Fଆ�m2�!}w���y�83Q�;"�۶Ս�����0��V�%���j��]�q��4�e;�,Y�p������v�@�F·j^
N�3�v�&&5R��:�]��o��7o��sl7�U�e4[q��إ�x��4�rլ��n,����f�:�̷T�>Y)h�Ӯ�v-
�e]躖o75���o1�P�1
�ꑬĭ�Z-���[�ὶ�sh��H��.#:��ne�s}���,���K�v�U��5Y�rY/�:��Sy�nS��zũ����
�V���`3[�u�v����i���a�oIP���1�$��H�I��|
���7�ˉ�U���˔�d����tp��p�T�]!=� ۢ�eE{��=7�M��D�ue�)�d q��8����'&��!�R벌8�wD=	�p�&_1�G��Z��(�Uo��Y��C�3��]a3��<�u�Y69����`;���b� W�����8Q�ȝ����5������xo{T�JM��q�>���i����c��n|�����&'�a��!YRCR ��9�,��`�B`0]�V9��V5����0^����59v�ޮh��BE� ^�%<o�]n��ú7��O���je�n ��Tͮ)��ĭ��w�%;j�"Wڄ74Dwqo
5��-��a���gui�BXoTʦ��t�.���Y��gS]�������초=�*E��?��!Vh�ӆK���籏�[h��jJz�i��&nh�p�n�h��B�+`�P��ǀ̚�e�roV<�HYC���E�"u-0��R��]l�1C�;�n�,��u'��Z�G%���A��z�J�N�Er�RSn�sb*����)MD/V�)
�Wm�1GD[젤hXx�	��)NPD��<�i;�|z�h�a��e����m�Ϋ0Q2Ю��+m����FS��62�E���]/�6����!�rcZ���n����dW��Hv�y=�r
b���[,\��I3]N�D�|f���&�o)s���Pۼ�uL'.*�;r�����pb�#r�+�^;s��J����Ь��#k,�Ib���8^Ӯ��wcvnV`댂:�8�Q���hic&�T�k��]����6᳓������U�H�5ǊQΡ�jաwE�)e�V�6��}3�}�ȽM�k��⮛ׯ�*k{^����X�����2Ea�����5vF���h�;&��xSGI�<�b�.Ո)���F���v)�vSw)��6��Fr��f��l첮:J����7Eԧ���:�+Żð�*1��Pn�x���`����ξ�ʥ.�}��m �dC���i˺תq|p������9#���퀶S{}��}�ob�Z_vV�E(`W��7v7	m\�r���ò�s����2��B��2Bf�k��mf�ާ�3�ګ#-NZs�c-����1],T��$R�\�R��2L�Q���[+r��k\Fp\�^|YK�J��y[V�2�l����f�7g[i�J�V]�-��䮘�F5�-d������sqv+�*�\����ST�H��X���S2�]LrV�3y��5�+����݄>��:iL�w��C�[���P�v�8�cvD��=Y�<��oV0�sT�ݬ��R��tˤ��� ]�5�P�(Ӎ��j��2�;V{��>�=ʝ[ʾ�1�93�56qZ�z�u��f����!Ju�l�}8�=���&Q����0
t���Yѐ���U�?7ך�!�szir>��{�6��'$�}a�X������;�7�T��E}K���R�!|��鳺e�Dw��ܟf�p���]�m�s��3v�e���Z5� �����5�����Y���3H���KoW�<
FP�`uv��ۼH��R1n�*�㗢�`s��[�(�j�S-��pV5w�gz��$���.�R7�EM�6ЗgVH�>#���ѝ�)5�ޕ�naD:�.�v�SM���tLR��M���(l�r\j�p����%��:��᥹�G���b���C���\�Q8��n;{n�����	V��D*���)BwM�"sB�d��p$�9yץ
Wz�dgw`��9�B���^��1�L�5�v�c��t#�]Ã_U��M�p��Iƛt�M\���/s���A�>��d�@x��@O��nr�.�"ٍ�9�@y�_h�i�IV2<�V��|�Rѓ,��%��2�9����(�O��Pg�"y%�%��6����1�޼��q,�[�c��P�V�j�a�juF�lU�����n��j��z>8�����p�w4[�E�G��������2��50'�9�(*���;�K$V9`��g�՘�S��ٺщn�n�eA@��@�� ����}���y=�y�������sz�{�lsE��n�")��Q�<��;J��T/���T;���]sZڱ���Oq������mS|З�j�y�q����=9SQ��X�Y.��M�A)me<ʐ�v���w��91����X������
�e�K0�̊,�L˷n
�|kMf����)@��LB�[Y��9�{\q�PxE.۷��}�
��H��$�e3:D�S��'gaavƴ6�Y��˵�4�r�x�6<U�6xb�Ơ�R��礜�{��G$D�[�wju�Hҕ��XZ	c�GHӯj��@�~�(�Euѽ�`�V��޻�K-qN�3�}5�'���\�	n�b���;�U��g}�%�N���������Ԟ� L�9կ:���̅!R�V]�Pe�y��A�J���ᑣZ�n��x��ܧD:��"����`Ӻ{�cӸ��k�B��T�����;�(�d��Ω��]u;�U���VBP-�?wu�J�]uuJ��:qJ�G��:P�u���3ೕ��&���t��;>\�7��dp֢Fw�ݪ�,;ƏS�{�y�&���6���iկ��ɽ��ivnr�E���J]��Qy6���
���MZ͡�.0ڏ)�cXœ���R��*�1Ćξ�{�;�}��@n��}lN�-�� r�[�`�����7����汵��<0:�o�mg�MTLɁD�kh�[�7��x�)`�pAff�@�f�7���S�o�
2L�U;�wiIn����o��������=H��3�����#���<l�l�w�m��]f�id�еfY���<��A��|S��Y%iM�:��R�Ӹ�����)@���ut�ZGU+��F*�Q�!E9}7�fBsCF���#�9R�EpC*V����k;R�	����#�&֬�q�=��´G��2p�Q*�LY���ق��Q>ȸ��#�\x�~kC��:@f�5�+9��#�k]�'���`�N�t2�5�V�i�F�[��fH�@b�*9ʎf`T��5�,�{��sQ]�p]�)6{[X���V*sm]�T{�%<�v��'7�3��|R(Zsyݣ1���mrۣ��余.��\�poR�Um���[Y�����K�,�{�]=�;��;J�wr̫h1k@��c*&;�q}�)�&�ƴ��j���Wv���0�/�^���S�Z�V��XD��5��m�5Y�.ڦeE��YBX���	LjZ��Ā�bc�Un�F�[�{�&�}yWpjF:V���O�\��%�F��+52􍵏;w�)l��25+5һw@`�:m�&��i�����O�7�.�ۂ�K�K��Z�yJ캘k�ǯ�YdN]�b�wi �<�
��n����π8(�3P���}��܄�X��(r�8^rWSp�e�T![In��ώ��{���Yb��̀8�� 흹C�/tA.3z8���MԘ��=�3:&�}���k�X���O3!�����|/I�� ��3z�7��su� /&|z��f��G ڻ��{$g��ϝ*��4��|Wbu�Iz̛;�����U�Y�9�W]�%���^�L�Φ�k΁�yu�����h�+��5t�o�M�GB���)�Cf�D�{b�M���C�t����h�mb�/M�9ҟ@�Z!�x��{h�cf��9Y�d���	ڹŤ]�Y# l�Z���W=� ҔM5,�V\خ��u>"ި����/�Z���q����MJݶ��Sr�^�+_-�׹�e-yԻCx�yW�E��� �*�Wá%���B�h�6J��qs�^�?J5tE�ec���ӥc*��UYQ�ޣZ�[b6q�7��&	׺����V�3kq�za=�1�k2X�Мk��o7�_B�Z�>�dC��9Q��u&oD�{�&K*�c�z�X�s`92ᇄ���q�.�K�ub�����8�0���S4�;A6>�&���6�����o��X����K*,�dɣRO�R�k��З�'e�Z�ޔ1a�A4��(�M1Y7�����V�(��6��]p�ׇ�1�R��jJ)�^��졽ͷt��ն�לq��ѕ����]�/T����E���j�yy˲oU�><��Q������3��r"��&�Xx��,�넭�#�I+�p��]M�ϳ��Gr˕҄�䝽t����I�7��:��Y���-������V��S���@b9Cmc��I��Oc�7C]���B���-Y��V�l;/�c7)ܤ���+Ƕ�rV���N<�q�m��Cx6� ʺ��'�kh[�V� }�.�m��m�[�)ҋ|�p5��g-$���I���x����.�D���Z��2�H�f8����y�ɑr�{�Z�� 7���󦌉�U�u�r�T�ts(<����c�	��;�ͩ��:,����v,���.}��/���Y[r>:%�n�>$w �E9q9gb0u�m���̫����3�)S�W�8v��2�����evȐL8�%b]�@T#v����	I�3�(�Q��N��؆uv]��f+��x,���b�r{���
Z|
���2P/rF�o=YR�9b3�r��t�[�\�*L��|�b��Q����v�k�:�h��ty�>i��
�H5�k��ռ=�����Թ U����9��S���m�������[�X*��T��3��XgP�4A��R�.��.Hӊ��^i����ܷu|���c�����Uʈ@�;CP�lн�ɷ�Fm�Ů�5���E̔�X5�q�?7�8�|���]N-ݨ@;��@��ca.��X��̎�i���Nֻ�PM��P6)��h�q�L����V,�)ʹ���k�i�÷%ݪl�/v�w:P�}���9�jC��
�:���b�(�W�������Q���Rf�5h:kΪ='e:=�z�u��t����4L�|�ԓ���C��v�>�����i��U���n�vB/v�����\�hו�2�V���9�	R�"�N�X�FLD��]/b����	yoD��O�qmf`z�q:W�eJ�K;�Rv���i�òK�g���RCW��&��ͼ��jQ�֪�;��:i}dR��=��V��gMr4HӐ��GM�R�giUf�@�1����%)�t�Lǌ�]w��D霞\k-)���\	��������I�l�fV��TC���5��R��S�wB}3+	���A�F(����hA�_R[�%^�v��ĩ�g�k��.X��l���:w}|k�I����,M����J����朗Z#dW��bs갫n�m���ҍW��|��.�zf���S��!S8O
�ȵ�[&Lgm\2��p3-Z���<�Rv��v�-㧹/�&�2���S[��p�"=q�6^����C�����${%u^氳�jneH.�$S4���=W��ӝ]od�]]�g"ѶR�%����kq�k1^%��}N���h����������[y�&T�u/H���'��@���D��V�K�J���p�cgr�v1��9�)*
���[lY�h$4��s�xnc�Ѻ���f�Y+8��پ[ O � j	���%2:ڽ�R��t)q�y�I��vt��y2�%L�ёm��8L�pA4Rq�t��2����&Eri�8���Ӛ�b��a�����Nϴ����[ulb�/�;��Xi��ݽ��Clev�}OE+��1		Dp�<��7��I�:�$4�F᝽���!Ôo���{;G;�9om$y�J�VC�=�Zᝁ�I�t����zj!�o�o�1n,
2`|f�b���y���н������g!6�_�7�P:�Ɵb���,<�gZ��d�ڣ�x�ZS��f#�+�}++��j�9�`�̊��=����}z�oo-Y��*�n���lZ�N=���2�OBW�+�W1�Ҝֶ+۫]�)j40p	�NʣZ�l%�W�M��y�)���%�\cA��Ŧ�a�Vp�Kk�5�ƍ6Y\L4���S%��L��ʐ��8ή#)椃�]
�eI���V�����' q��trݬ�&�j��]	X���N���v�a�c�t{7Fr@.V����w,Y45N ��g��E��3EDhڇ^���$���D]��z�A��xx{�
]	TZ��,0v7i���cs��y�����ҏ�v(*��9;#��:�\�S�c]ˑ0Bj'{ofM��y��1i��P$�Ȗ�тiM�����듥˸Zt�=!C�T�B�$5�9.0
ܛZ^�P��ױn.J[XX�n�3�]�gY�ݜ���lH!�I_e�.ӭ�X�st�UMl^F�;����4�z�^�zɾ�s���h{�i)~�|Ūc�]ۚA�T];h�љok6��ϯ���V�!m�_8�f2o8� �H�s��̀��:�GՂEF\ڌֆN��Q���w�u�Bb���blv	�%n���nc�4>�J�;�e�v�h]�ޖt�v����,kqU�n�w���6+�1���zon@��T%�|�%e\��"(�V0�,˫�G�+V �,kޘ�][[O(�ϣg��{Z��O��M�;�t��A8>޳o�yȵS �&=�2��䇈kgufؠě�7�.+�rI�݃{/��]�h�����ಆ�B������N��GhC��*�s���h$���Z�@�q�X����V���'!�Yc�8q�����,k۶��%H�����-*����/��u��$Jm��w]e�M�;�!:6P�哋'�u�s��H��aU�&*��۳�q�mIe�)�[�D�6p�=���I֚1���k.�o˗cF�k��~���DDc�����Zi)�&-��p��R��mm�[l��Ng5�֐����Y�m�M��ڱ$�ؒBY��3mkl��!;[$ֶ�f�ql���Ͳ��m��ţ�L�!����NYgcpض�[���nKkGH��6�ĚVIm��q9&XP��,��k2	$#���1H"pF�gXgk[nÜ�Y��M��A9�&ئՂ�m��٭+n��!;0��vkc2Z�m`gf��Fv�g"��-�
Ӝ塱�p�6�4Y���8���m�-��N .&gD��8 �ۭ ۛgY)!Νَf�:�Dr6���s��e�,�6�R���R�tde��:9N��jmJ+9��p-f�8�.\$�S-�'m�@t$9'B㑝gi��f��h���)U��A�����M�.1����1�qE1xK�N�+�,��%�U�gp��h�� ��m�;��=
��:��u�5|r��&�6^��T�Vd�^�����o������ڟ�3�e��_%���"b�����UmKD��+�����=Q����s�V�U����嫻����J���U#Z>��"v_+�Յ�M�i�#J�Xط���?d�__XL�=i��!�č�h3�\\L�yqR�y�O�ΨU�p�Zh�h[��-�Ump?e{ȭ�X��v#⽨ݤ�ΝW�^��V��+v8����h6�;d�u<�zՄ�s7:okfrk�����k]^Uۚ�ѱ�[�pm�y挢��^�ȆD�:�#[���,hʡ�:��'b�*�a��ct�[{�mmD\^
�	���������3�E��f�s
�{v��|P}������\2�᝛�1����0�q���k��>��(�N2���ƛ�HQ�'��*W�#^v��d�ofŃU �Yذ(��0��kvKh*��wu�8�r_M�W�)v�y�/X�;���`$'	�|huH����x{,��&ʣ:���E	�-yU�i����[�G9Eh�YYC���W2-��ib���bt�<��U��!U{�V���oYv���f�9Z�lH��R�9M�7:֬��.��H+��$��5`&��e3;7���3bhnGiA��F���w9��z���g�>��$b-�4Ս`��j�w�}��S�t�W�YWV���֑��^��zP���;�|S��m_���Gj��e�a�c�3�t=�wNF}W���c�N�K�]�R�;�H���H������[D�+���b�c_C>��%�e��^ޡ,$}U�%�c{�Fm�[s7g��T�g-��S9*�ܞ_7�(�FA�
B��CH��]����Ak��K}6��������sJ��|ϥ���pQ���
%P�uS�q��j���J�:�{&ߨiN�7R�Q�uC�O��j÷6&�fP���c��bJ�<��p�vКX�:��J��e����q!�-��cn���%o�Y���*��r�dË#��o*�p&�7�cO�iB�}�d���@�u�n�ѳszg\�!�&��8+T���u�3�SV�i%�dQ'spކ���NvK�N�9�/,�r�T�j��	l�؊�:��X�֯� �5�qNm�N>����x��r�n��K�Z�.���j��T��b�(nk��ѽ�ݎqLF9;O&�j4��[��.W,�RUu�g�:��7b�(]�>�v��7y�y��cR�<1�����4��u�[�0)"�t'0��c�9�C�W5�r��כ�z��Z��3مZk�|V�j��^
]���W��ވ���2�=�o#չ��uzX��/v�!�[ٮ���@��w��/#x�ep�v+�OR���i��%�f���.�)�;7�d��.o'��j�;y0�T����:�ӟ�gs��Cf����<�QRB1Fko+��GV�'�=�ˢF^�� R
�u����ۈ�
+���,�����7�����j���b68o\��X�R��<��12$�ܽ��Τ����[�g=n�Ȱ�k�28u�u6<�7R�tN�z��P
��`��#���f��}��۬�f�tW�8�&�3�3^f��i�o���:(�����6�n4�������F+q�^o���׶R�u��=O},��[τ�"���F�@���F:�{eM�7�G]�}�'��̩x�z\�������zS�c�P��dE�wr�[L��q$zӴ�g�mʁN{��;����Ձp��O�:�2����,���#�B<�twHm�(K������=
0r�mN��%7��r��:�i��^׼ӫA��Π�(��E��^yc�toā������P�j�÷�"�㭹
	{�f:��q�&j&�c;�V�����:��(���4�l
f�qa"йQ0{i�
E;d�T���kP�s��������R�搛�bU �|�.����qt���Qe���b�ޙ��9e��j�X,�a"��������'(d�"��k�N��(�nth���痭��{�xe�W���۶�0s�C�C�;9s�U�U�p`P�.D�~�;۔��q����,�a���q_o�q�f�>?I3���;Ze��k��n:��v�BQ+=Yj�I�Mwh�`W�.8BS0.)h' ۧ3�p�">�Ź�|z.�WVl���2l!Z�j噽ӰMA�s/��g��+^�M��?�^:'֗W��r�1,S��g��Ό^�.��� 4m��K���I��u*�dj�ڡ����߹R�Ea��u&g$�m��s�������|� �L��P6�5:���͉<!ف�/7j�ػSt �19Ų G\�=|7��˺�bS��qw�1`���;�����O;n/η�c�&s�����$G���AE}t�{���u҉����3�b�g��VܐyV{�9�E�ˡ�*�mN��yֺƐ��_�u
��M������K��jQ�U
]E���V�����cX"ֲ%�eF9�T6%_��&�¶6��⍎xh�Y��eWw�a��%�DƩQPx��P�X�炠:�L����Sn�ئ�K�v��_,J�0:TLX��h�"�(��n3�[��_�:Y����ڝ�.���M��f��\ն��n��Y�a��[sK=
Eyzz	�r���t�*.,OWB�R�B\(W%yI��Q�,��[7�����Q��y�x*�qt���ѡ�}N�Ԙ|�k�[n�\Kf]��Vn�Qf;%l��Μ(2��v�3z$������)�پ:��j�/�~x����c����9��V}����O���uC�(�]�PY>P'�0��fd�F�"/��x�'Qk�!vLeLl�iF�^G���aŎu&^�vjO��#c�&�Y�*,����U�$3X}��Ո)���t���;{�K�7n��(Q玗H[Ux�kxb�Ϳ
�V������,4aV�".&�M�����#�=ZOJ�ܥg�Y0ˠ�c.6�ܮ&^�}S��N�6�%����*gcʳ�4n����`�[�a	�:VW��~��q�6�)EA�jŮF܋�:�b�.*{���n������>s���g�3��	222����9Ir���6��L����3I�{��dnd��kx�E��E⣲KD\��}����*rV�.��%<.f�zMffN��ְ�%��2X{�㓡��}Ad�k9�Õj�kʱ�e&(��6�iDD���
��}Ko/r�6_U!
5ȧ-:pe^F�>#c�5�ڞ�؝S�>ꂲ��x�o�9>ݚ���q�^�p��`�g��&a�nl�.V&}n�!9��4�N���O~���#Ќ ���{u�H��PT�T���(_PQ0@�n�8��)`�V��������v�dq+R�s`Qc
��mz�O=~4�h�L�D����g�� �ث�T�{���W�otX����p�G�XJ��CK�z��/K��L�Z��mK͡�u;=.�S�/5;�z)�=
��p�{*���qu 8�����P���|~W���#�rS�x����䣖�ݚ�����ȯ[��&w�lXm�ϋ���]r�S໶�!�oʞ�c�to�~W�.�t5��a�V��,4��qg���jv螪����԰��ܝ�e=ܬC��WB{Z�oVt��#�*[ʏ6:�R��[w�T�WF�ڑP�/�B%�w���rj��a	QPª�r�k\b:s�<f�Z�\��;s;t�r*��}9Δ�g�ˬ��L�lBr$R�T��4�:(�kE�D�k�@0�{:p��7��Dl7!xj�7�T�a2���ˇ8�E+����͵���r�[�z|g�:D�p���42 ��K�����Q�t�2����Sa:��u]=Ξۮu>Wb�բ$�A�>B}U��I��IAa�����s���<|W�+����暝��"3�$�A�^Ȣ���x�;^4��`�.ϼq���9�$)�і��iN�ydrT���=ψu>��!z��No�؊j��
}t���l���v �Cۮw{o�d���:�Z%)����3���'k�ÐVQ�ǄTQ��H)�W[r�}7�U��gw5�L\�:U����E�~�ɦ!�j�!�8�a��x��^����E3F�����6�>�Q*cg�&�H���a���eոQ�U�bi���qnr
t-��O�d)�bH6�����gq5N��ܭ)Щ|�Cp�wÍ�J|�����2�=�̾b�c�}����w�^��>]��h�M]���ư�,ʜ�����ts{�]h�Sg���l����r�V��>�ջ\W��P�c�Ѹ{
&�b��g�N��u�d~�A�E��`L!.��J�gQ.�Ɍ������vXKu�<��:۽'՝���q��J*��+�X*ҥ��WP���ઞzr;2��Ɇ��k7NW8U��:$��z�y��c�&VK:2�p�ؚ�{�!;1�b�-�v緒+Y�����-U��9j�Ȱ��])�nvKJ�Jb'�h/WB��y\�̭��E���U���egc�w�)fܨ��Q�v:N�eE�|r��P1"T/�!��I�v*���Q�φ�=�
\P����^���pLo��X���\����t9M��\ɬ�k�F�j�/�a��h�i��DHn�=N)�T��t��(�\>��	�÷��z��\�9���Ķoz����L[�����I	 �	�+`DN�,�s^�Q1@��ץ����3������R�Tv?=���ؙqv&���b\�ԑ�Tu����wKCyPN+�\"N{��$�x�~�E�T�܇aں��6X�0`f��׸S��r7ӗ����*tc..S4شQ�Ń{�|ڙ:��z{���C[k�k���R>�cFh,.�>���-j�bs�^y9��-!�Z��!�˷e�k�	
�XV��S�t�Ju���<�;
���h�J�o�^��w�|���p]]�×��3�H̯a�V�Ks�Xb�.
yGg.Z��A�@k^R�"fǎ��׏�%u�/�^��G`7�/vi3��wR�i�B�e�=Y��B��o{x�s���/�v���%�E@���o�e��q@�����&qFfqռ�'�o�fzD����ú�2�DR>��t~\U+^�|GdK�D���㣗�o'w;`՞bڕմ�#Q�*�?2���8]��{T�1 ��)B��U���M�\B��N�����.R��ۀ��)�x6H-V{�9�Eŉt;%FyW��U�4G�UC�t�i�]+6B�V��n��v�1ڢ�oz�K��)�Z����(W�eF9�Pؕ~�ؔ�vu.s����eu�p��Pb�m��z�Lk�/�_�6�@%����jN�+�i:Z���ϑ��^�ځ��Ԡ��цj��P;��g�<���_K+���Ne�û����9��������}sK ��"���DC���t�YB�G��^�)��h��s�J��	��]���$��>��j��W������S�E�ᗙYaʛwz=K��rފ�"v��6�x���w�����ͼ�1	Pu_E|����sܾ�>���]G+u������$���M����w��U���)�r�c��՜�(k�]�[�:.��zv:��n�z�|��<W|s��F��)�:�������OU��<�Wbၮ)�S��(���A���&oD��d���A
�DUFΩsc.�u�UUx�"��gz"&w'���i�r��vuD�;�'~&\!r��.�L�ʌQ�9��0�W�:��^-���R�%�6o[[��ZdQ�ב��p��Re�y�5%�b6�VMk�w�jI�B�B�u�3I�u����=�#]gȱwv� ���멪������qQ��u��b&��F�܈�2����f�O�PQ^����dU�92K��M�-�*Þ����D�u��몜�\Z�Y��0n�"�tG��
nMN@*���※d�ܖ�����1�iY��� ��a�Xdt�N泛&������`T�9
1*��./Z�L�p�2�Tt�ʤ!E�T��Ӏ]�k6�ᮆІ�c������~!tK{xx/<�Ě�C#*����/�*���Cr��):�h2�8��䊊[�R0�5޺���y=;��� 	b�̒��m9W��ד1�'g5n�:���>u��[D99���dcE0-WH��Ԋ���ȴ�P_p��*R�i��+,D�b.�nA�dqx���X{��P!��鬝�Z�#�_L)Z�1Щ:�"5b8��3 Ļrܤ��V�]^�I�Ř�XTw�/6��7f�2���\�P���C�&�$�6�}�P
`��1�r���;B IC8�����4�{ħ�7��.zV�W8��|�T;�cj�M���W2h�����z�ۄ�6Q��c(���1�hm�哖����%f�"s�=b��vmQy.�7������m�N�v�n�2b��}6f( yܩ=��約��v5�J�Iuv�6y��Z�iog1��_s��o ��J;#V����;����Z�ϒ�,H�����u:x8�s�����7��-�J��jj�ңp�G�S�	�|��ihX�Ig���:�4.��	f��T*M�5:Wf�j���W"��z]L��^��df�R�c�*��.؋=Sn-]�Ꝺ�H�o��5'Z�y/Z[�H��<k�Uʼ�4�.WJ�0��3�C>��׽��e����7K������ FR�%��L�د/ME�[��/P�mZ2�5�K�\�(���U.C9�J��Ȗn&�ō�{��٫�Y]  �J��$ӛ�S����Fv�y´=
�u޳9��,V@�����t�T]w)'�9 u�Izx	��͓\Gu�\�j�;8V=Iތsb`�	���/U�j��_o��\�@�x����[:���NJ-:�L��ѵ������$(��h�=p�O:�Px��|��(wj�"�_GG�i#�q6/VaꝛL7�h���c.P��gm�mou��r��.��-�bK� J�ra1^�Ά�H���CF;�-&�������o��,��]��: b��b��u�n�4ٺ6�*�\;�i���=㽴ˆ���̨M�\�m�m��b�_1�1x�oYlդ�؉�5�K�n7�xg�l�v� �G�2e���q9��Yy٬��{�ܗqRd�]N�mɵ�wnB��X%�5��� ڹ�/wn]�v�e:���`m�w��zS=�:�\z��O9�s�m��XC��$&S���-0z�Hwk\�1r�W�L�vL�|]���ZL��X�%qkm�������m��k�q�t�e
�]�5%J�쇙7W�̰�����s�J�i���(;1rM⁋̡OH�]nq畅<:�K������U���K%-�rJ�J���M��8�Q�x���48-�֓A��@����yU�
vSo�^P�n�&���Y��հ�!9x�IPW���9�z^"�AN��b�Җ��|��[kNm�QF�����w�Լ<�>�����^�5�w�̰s����uՄС@h�D�G��B���[V#���ē��rA��DL���::G8p��\m�嵈�e��G� pp%$����$"�Ŗ�	�'(%[�㍬�i��"�Sm!�m���'8II�	5�Bq	H]f���'Km�tR�qC�$E�qɕ�p�B�9f�NN)�N'ke�f3N:A$K+.�8�Y�p�S�[�ֶ�6.,I:�S������S�p9H�m�����HY�䎈8�:&�Q�JL�kD�:�L�(�M�$�Q�m�[�!$J$���� 3@s��)#��"cd�q�ۭN�N( �!(c�e�J����78��H
HB���R\�E��AK2F"-4FU5@�����s6b���v�Ƈ\XWw��5^"�Y�AmX�h4Y��aʿ"�<��49�j�U�u�x-n��������d�6�7:�O��~u
\C�`��beʁ��Lb�n���+X�ReG�U�/81b��.W�$�O���=]��蘠FנC{<h!V�D��1���sV5�r��.D��!����o�]�C�>w���x���p�C���<6c�=R�( T�r}I7�����^�wv�ᙜ�"S ���	�
Ľ��#쪰�8��~��W�%�ѺzP�ҭS��o�,��o��r����p�85�9��,�X	����N�����8`��̘�-]�FҦI����ųG��dX�JU=/�:P.��������d�3~��Hѻo)�����p뉹�<�Y���)ň�nGQ��j�r7�d+���rU���+��/G���DE�T�h�Z���X�j�i��BnG� ^^�u0Tû���!��j�E��a�@�,�Z"O�jJ��8�=R\�uW����ϊMZ庪���ͮ䉺�eMt�:%�Ѩ '^Ȣ���ci�� pt
�0L�Ks�����mv�֧Cj�;:,�~����Op�r�A=�y���r�)�ww�L�6d҈���%�nX�:����db[��9� �o�����"�N�v`]}X0��BgX����b�b��P-� �{��K�R�����ڝ|gs�sn��x�����q�	M��Fs�h0�8�xk`϶��U���~)���~�=(/�=}*г.�ф���}C�/�v��2�-������_��v�.������.È�	E1�\YN���$YWHC��E�w8�aٗ�׼��6c�X^��q��a7=�f�^�AUZ���Y^.����k�e�Q�>P�l�r�2�ܑ��eE��ع����ʄG %=�\��h:�<$�5"��g�+Υj3����3�᭘-�S\$�='��zǻݾ��p]�t�S���V
��{�l��)��.�z�t�P!γ��;7��4}z��{*���Q�O�}s~L���$tm*������]W�&;/j$�X�<�|�{c�j߷�EӅ ��<d��#��X�T�8���7R�D��=�u�
�ib9݅v�<�}�ȷ�:	s`R�E�_)�nT.������lʋ��L�{Qt(�x�^&�ƞ�r�tHcEtWL�P��mK���=
0r�mN܄���]R��0mU19U|c!@���nH�|�e�X�=����4�ݹ�%�@�ޱ�5[,*��7� q
}i<ZQ��Nx��7��
�Z־ 7����wt�Xi1�nQ�Q�L<��|��J��-�ޙ;�e�9h����{�u�5*�zU�3]v�D��u��U��pr�z.NN���]OW�+E��hV� >F��Fyt������C=��83�Q�G�Ю���ٵ��-�]����B�}O��9"'.$A:A
�&k��t<W�� n���9C��vf�a�W*�.\8
�f)N�e�ġ&à U�M�x����ゆ!�b�'7.���F�|\�4G2��m?9�k�	�86��9C%�{]zhp�z����������=�Uo��B�)N g6Ne{/8� ���s9��/���x1�B�݆f=,��z���vk���u�Y�a��=�wҰO�'��t;���!~L��<����6o�޽|��Z��KD\ϔd_�Ks02)`' �e���Z�o� 1��Ep�Jg7�9����;�=�l�]���pQc/~"����?.*��	�#�藎����#���[��e^�p)Kh�@X��W���v�s��͞��>��AG�e�}e&�Q�d޴{5�\-<�V�au�E9o6H-Vsg :T〗C�Tb�3]����m}�Z��a�����b��#��Tuj�bJ�8ؔ��)et���Lp4�n*;H�˕}�s�����Z-%�>�&�>�a[7�y�3ˍ\[�O���*u�l�ժ�27�S{jƤ69l�Y�[�3;5�u�Veϒ���[��R1��P�Iy͙��Op������P��UM�U�p3�*��-X�aB�eF9�Pؔ䐵Sf�z�.��c�>�&ġ.X�A��nU�D��**���9ʱ�����jdwE'$Tb�OdU��k�,��,JӰV�D���A�K
z�f�(��e�����࿎t�t���1�uuh�9֋�,][��}~�vJ!�[
�q��h�D�����A��У�k�r��eq=�����r�*q�v:ɻga_����OA�Nr�4:��qh�>�ha�QWp�h�Ӕ��ˉ��:C����:
-`�A���&oD��� PB\J����
��~֓�7��ky��U���gvҜ�`�Q.�N�L�B��ˬ<���EC�\�y�nqo]�Z�pB4�+��",�N�I��c�+7Ҽ&�k�;���W�t=���Q�R�ɝ�8[+�v魥��V8*F�gѨ-����y�ۑ~�[9ێ{{s�_p�7U�_��z{i�3�L.j��XÐO�PQ^����}�^�G"�K���q��-Ů�sǇ.��"T!l���C3��]G);�+�U��ZI�묕��#PT���{��]��H��q])]��P�e�xhtWdk��rJl�^����^��!'R���Wb�,Տ){�d�0m:]Z�	��I�3���Zwzc���x���]EkQ����l�X{}{�Y��ms5�}��{����|jǄԫ(.�����noY�w�{İ���^A�eх���|�����sd���s5����4Q�u������1��Е�:N��GN��LB��@�n\
h;Y�`'�ltf�Sו��=����j�']�j���нQ�����SЍ�&a�nlmQr�&}n�!9���ʜ�L�����{u�6_fw.��������],O������`�n��9Z��<�e�v��ru�%�8�:nUt
��LQ^�"S��h!B��7̉�}A9���W3��q�ŋ�]�wH�K���򤠛��~�2f����5<!��Hq^)2��s�p6si�:�
�T1��u�Ҝ�s��c��]V���ԋ�{�ER�i#OV��œ���C�X��P)����"��|z�w� &v��PE�n�ߐ��n�K��h7��;�p��l�;��$E�T�b����:P.���WL�O�2p�o����_�ҵ�����l��+6t�թ][}��n�1(��LZ��~�s�@�`<l;ˉ��a�����H[�OW�;
�����r�}ټ�r�b<��,�j�}��gׯ4���OI0��ɝ {1u�Y�;�3qØy����-�	T�J��#�x{�)��J��4�5tl@���qH�*�Z$����������W=�^�y�H�GS}X�\x�E6}
aț�*�C!_�'H�;����˪�ޣK���d�]��;yT�d���@�0�N�������r��t��%���P�9s�{|�b�Y���j^B"��F�����ѹ7��ԟpt	B�	����3���|�v��rºi�Z�`�٨nW��Xt�b�Y��3�=&f�P��|�.Q��ʋ�y��y�N�K�4�Qh�&I��>:��������g�=�Ŀ[����U���yh��˻���C��5��V�7L���5����]���P�F�Q��8�o���s��m��'�����I��[_���(�6��*.Q�ɉ5��i�ێ�Uv#��\t��{�؝�^����IRjEC#��@W��V���;�a<����9u�-�j'�������*��7��-҅N �U���T���#�c��b�:�O�!�#:�ڙMx�>:�*6l��Shd�Kz�jKy3�+og���@�P�N����#�;�Xk�
"uOT^`���q���g+/ɜ���[e���=ݢ*5���Q���/�WDo;Ж��SI+���KTp�1�>����1kV�UK��]M�[t��j�(�k又��S�J�L�M½5�a�Ֆ�^=K9���"�3\"�P��P��Q�65V9��(W����zh��.;'M���}��]��wm(1,�(dU ��\׫��H��JFlە�u��ӱ�Bu�*!9N���ڧ�J��EmuK�J����"���U�p*�4�to[/���3��o8]Ь�������t���n��q6ȕ}�F����7��#<�S@S���A�e�r�]�>p��bo�[����h�
	��Cub$���D	�+`Dlb�H�7�����%+����RH%�ba��+�=
�F#0��ˋ�BL=�@DWML��=X)�z��]�_b����&�.+Ţ(���Rox��=C-��)�/H���]zjv�S�#��c�xzv�!��Ү�Жo٨�5�����
���0s�_�ú���kA��)�-�q�'{�a-�oaiz��+hp�ZE�F)ǭ�uwҰJ���O�P����Մ�w�����^0Q�g�8�5C\qY���o%�7�o�Mw T‥��	�e�	�=j��|7,�gUgH�쬈�ѕU��\�gi�Z����rYzo�2����[�A���9�Z{R��7rԥ�����qU\ZC.��\��M~���#��������u�{�l�#+>��`��`\Tɇ�ˍ��q��5�2�1�'5�Ur\�a�����a���9U��4��><e+^�������4�&wj-��3��)�6�_��|�"5=���	��*sg�H�%
�������e��~q��g�W@``֐�c��^�p��Z�	��-�\쨅�6`���*h�[�-<ut6�N��V�O�e���T��Z� �����P��Q�K�7�Wۃ���ޚ;����c)��+c`��N�AT"�8碠��[3�m�aP3�r���l�c�¾[��"��&�G�x��4�:5�;)�<�*��y���YPri�}�;���7JŹ�WM�V���IxD����x"�H��=�\%T+s�ʋ�lU�}:�	љOWU�Wqp��jntr�v�¿'ہ��C�Nr�A}�t*ߍ�h��XDmtbkiT{�EC�vw�B������:
.�.:�ב���� �!"8�*a����Y�#B�"nv�T�*:�"��"-F^L� ԍ�7�뗃�*�[���]���'<�	��eM��eWS,d�ꅷ"��a�·�5mlMa��͒�&x�U���ƕ��r��ꊳ� ��9�J0�.vy�4⳧G���ή�ӭ���}�}��Pd�֊�k����'�l�5{^��[�yO��m�z|���|%+�_N8Zlh�KO����]ݫ^����4��#��)�-�(�]y�7�/]I���Sӗ�1Ni�`���Z�
�ldM�)���b�p_#^��#�|K����E��t��c���`�k�S��ՃH��>���	��^�j�xPQP�_���N^2�[�-Rxq���=YJ̨/͛�+g�d�����I63^�>�X�������յ���u�x{�b���|E�R�����ن�`L��PY7��$���s5�����륂�J���q>K� 9�����-�0ʴ�C��U��
^�M����Z�짂W]�P�}$���M�1[|�P"���u!Q�.;=3BS�4�w�>e�N}.���n��ϲ&r��]'��r*)f�D���������t�@ _PP�]�q.T��mݧ�'0�.�u�]hh8�+���jl	K,����wZ���AS|�dj8_�ߠ�E�Xz)�6S��wP�̤8����8R��S��aU^%<|W� ��d#=������d�Y�v{|J1yZ���/�VY���s���QS��G/��t^�[�>���X3y,�֕9N]C4�]̩w:���@Y�V�59K�Oa�٧x|<���[Hr�����m_J�qT�1������8�ؤ|�e��%_�kz�E�v��i��5��A+2D�g]C������M�:P�Z��>�{*��qu>;ӑ��̸��i�Mի�n��� �H;&�z���9�U�EE�ǡ�~��V�vMA��{�
Nn.q&2��υ\8DDd���k�b9��5WC��t�]YwЬg���7^��Ǌ��|w�b��wkţ׮�E�/�\9jq��v�.���ۜ�8nE�Q��X�NO\M�T;�ձoajW�f.\+%���ʙ��l�(*�"hp �F�B���&(��GM�k� ����jo�R���a�L�	ש����������/���]��ࡽyZ#7��.饻��1i�7��/�bKh�'^�-ѹ��pjH�������Z�/C�uf{�҃�9�\b�r7f�9C�×���7�gۃjݐ	qі���罍x�V�J��1�&*8�{v��N��B���2�l9��x{���^�8A�xѳ�R]��rN���!J.��\TV��/'1ω����؀��"�=�������+���A�ʭ�CU�޶�=�Vo!&MVjp�A�G�^��4�Õ"gm�S���N���>ī��ǂ��3D��"y�f呠a�N�e�R����(a�+�#��mД���s �0�ۜ��[�f���M�d	��Y.�NF����^�����,�!hk�yLL����j��-���f%E�Gp�ON͏��!�����勓��o��ڷ�i�*�(,�����)ڋ�V���gaS玭���������W���b�}�2r�W��n��ٖNnT�.[�rP� tW�J=�ۑ���5��|༳Z���#7crƍM�؛5�Ql,����]F�m�����U�܏N�0�[�B�.ʉ�pKgW]��mU&B�@��m�7���2@�َ�0Κ.h|�BGNP̨����r�a�W�W���>�v�9��X���Xn���|�-�JF�F�k��xs�F�a�t���Y�6�Ų$�n��lt�8��쨞w3��K�9cG����w�!-�s1���.V]�5�[���K�Ye.�|�_��c�V��-r*�k���:lKV�ĴvLޣ�ݬN�k5m�vјk�ؓ�h�F�v�m�׽��vi�.�#�*��=�����������z�YZt�V���;���,\+v������dTFd��_6_DUI��yS���;��YQ_U���Q;�ʭ'bJ+��u�@厂��W|��K]���Fmr����M{f����d�)�7U�P�`�Kg����SŶ�:,v�|��;g%��NO4�h^�쀁��M.��R�{�d����u�%ˣ�f@3J�իF��S���1i�n�o�=iDYol��l��o���z�S�G:�
ٻ�ؑ3rT�I�L�õH�b�t�L��'�v,��JQ���b�^��C3�!�qL�˼�2\�Q�>�UԲ�5��o���\a��2��J����Yt"�x"xp*<.�uҽe���w�\�����R��E�9�����8`��ö
�+2�^4^u�Z�]Zr����:�Otdޭ� �S��-��Of[��2r���(U�0�����@������!�T4$׎�X[�X� ΎD��C���c�6��с��^���9*�R���/6ު���[�n2��v�L�O��:�j8{a<F�Aڝ�Z^4�H�X�6�T̢��Oض����׋'*s�ss��8�(R]g�j|֛e��I�9��v���4��nrz�5g��4Q�^dG�r��c��߭�:�� �g��wn��[�Ԕl��T%n�hV�s�����Ϋ;��u�����K$�ʤ��t�nv�XA��ofi��S�B�x��}�@�$�u	�]����w;y�+7M�:�"·�6���۾JJ6hv�]�ܮ����r��ϫ���{�ؤE#Mj����mv�#��p�qҜ&�G"'#��%$
*t��w-�H�N����Y�B�J)���&m�\�m�.qH����n����s-m��Qf���ӎ 蓒!�7rqCkt��rp��N�Qp�9s�9����L��d��6�N�\#�9�	�C�):IgZ��	�!����$�� �(�).")�m���"!L�Y�g!s�����D��$JB"\t�H��q��Йi�;�
'"��%��H"w9�E$�#�NgaȔ�hr�K�8m�q��:�N�݀�#�AB��q�ڷ�]�8�T�ՂQ�$9:��f����u�|>
��Ĉ6mcܙSyޱûk5M�����8ק��,�Y��Uΐ�-w7��7�Jè���d]�y#J�F�J��&�~��xV>�3o�SF�E\�?����ʌ��V�$.�@��!�f��;��^M�Dm�]7�'�/����1m��ȭ��D׶�ϰD�����5����xp�K�v�1��r���K�β�啳��qnpAN��`cu�=e�%Y�Ӏ��r�t[�K���N!I�[�n��<�������	/�s�����R�,2�|�H��}���̝M��AI�;th;�Y�Q
aU�×D�u-�E�i6�L%#��!l
i�U��uD�(S=����L=��,����{��1�g���%;�Ih�<g��2���Mr�5S���C�o�x@�RC�F�K%�(�Y��Xq�AI�]�̧Y6ߨ�EC�)���互ٶJm��s���_oҭY9�n�o��\��� �L��6��8��Y�@����p�e �ٝc�
g�R,���XRq!n�ہ��ah���Xa�Hu��L=Kd���ׄ8��0);��䲡�㏗�K�J���
 1������
e���Q��S<�w@*�:�1dRS<��B�D)����x4���ZA~�٦KC�R,ǪKd�)�9;��*JN����ѿ�f�������y@�� t	�s��f�RZ>��a���'h\$����]P�m�aI��"����gS&*@Qvɋ���Ra��6���}�Y�j���ZK�λ�b�-�4��#y0"<�{b�{ I��#��O{AnP���v�)��BҐ��l�i �Շ[i��H)�v�%�0��qD���Ob���ja��x^�yǽ0 �N���l�o�9���k{�+���p�X{��C	�N7��z̰�
|�����Udu���Lz��P����ʲ��>�����S�а�a ��v�3l)�.��m�'�u�ִs�Ү����Ms������ � s�dc�/qmN���ۼX�N�b�G�
YSuUh,�:�Ȏ]�b����Z��f����eպ��Q+�٧���96�Q�u�R%ܺ$����vP<��c�m��*��[�C�@}��b��rsSiޮ��� �[�i�{��@����aH��3���z�d�O�v�:���2O��Цy���>;�,<����Q�&��y���aUIHVYI�[l��X_(�0������5��k4�t��@����P �1��8�"�b�['̤13�<�R*Mse<��2��/)<�3�T��I^�R,0�Ͻa�I0�2d�c�,�m��}VXJt�H��{_o��;��b��τRk{��� "��يa ��c�8�4���8��f���[>3R[>I��}��A`c>�0^�I5�ԙL��������I�Vj�r�2R,
�=�_�Y���c5�~�����P��{v5Sl��A�B�0���n�u:�H
br�O�H,���M2y��>�C>aO�3�����ͲS���{T)����q�>��쟢��ㄩ���Lwr`g�B�|���,�%�R�fY�0ϘR(}�%���&ó�2�uP�0b�Y���RbP����Ka�T�P�%9I�0�HS<ə�gƾ�T��_�~�������S����k��9�u
g���eUI��>�)&Y��N�Ì3�!Hj{צy4�l�ZM���a��0�9�ZAd�R_(S�a ꂘ�e�X[&���`{�c��ޒ~�v�Un������_�Qa���\�m&Ц�p�hY:�3�v̠i)�%#���<ɔɠ�nM$�;��9��l�P���r�N��n�[8��@��*@����}r��l��wf��3�E��)��T�@a-�9P��qd�e ����0L�d�Y4n�(y%>a�5��9��N⏎��e��n�O2R��0)�O�H<퓈��󞙓q[о��{�;�s��<
m�Q�H,�Ki�wB�_]@��VR��%n�S���a�a��ܫfY�-�aH��v��):̛��e ���}sH��)�����f+j�	ڵ�r�`dL(�D���0�IN�چm
e��(q�!L6��a�qD���7&T���a ��b��-�V(�95�3��fR��h��0�Ze���%��RR(������[>��]��ݫ1kkӑ�Ԝ��o���WQ����)��FF�Π\�@TN�C
�˧YI��#��-���Q_e��Ůgu��m:כ@ŏ���!�+�@r��e�s���9W9x�+���^գee�q�g?�W�\�;]��W=���~>����i�k޸e�4�al4�L�����ꩄ�r�M���S4b��вu�ћ�2���&1bβRAp�}�d�E�{b���S�TGG��Ojj���k�8 ���=7#�f���L��e ��<��p��PƽpۖhS&Ov�;@i-�;A�U���KH)�ҩ-��`������\3	6�a&3����g�3���1�ַ����i�a_\�gP����q���m���|�����o�u�7P�&��
���
M��U�{#ã�c�#n�c[�yH��C�Tzb|��,��,��l)0g�C)Un��ey� k}l�IO�����`��Jt�/�%$��38��5���g���4�h�(S�Q�J`*�Vu���4q���Xߏk���AIY���l+U���
gR�u�KML��a�1��0�Y0g{��O!i���ĔřM����d��O!L�(���i ��2_���&�I�+F�sw�3;��p?R��k��DG�QQ�ty�2��"�8�H7E��Ĵ�ຆ�jM2�A��)����z�&R0�3]�4��) ��˓�X/��7�%������֏�Ӷ�Ɵ���._{ l�ﴙ�IN�ǵ%!���z�*a�P�����2��S���d��'ͤ�(-&P��&u��h�0��1~�����l�dV��p���)=�U��?sw�f��1�N8��ߪZAI�O����Q
N��3�Ka���a�fжeNT�AaL7tRB�*g�,0�:`��%!�J~��xeȸ lL_�r��U��|��g}�Gj����tt1ﺑ���C�c��A�e�Q�'���^Y�J`*��!����F�aZ�9�\�3�l2̽p�Y����Ii��}0�>�*=�pTLUk�.�����K=������)�0P%$����I���:�q�Y<�N&Ø�H>�d�o>�� e)�o��eq��gܰ��O���ׄ�C�2�������6�N��ӓF��9��Lu�k�&+��n�6����ja��f��V^n(�b 었���2uz�ׂ����Ѻ����qd�CO8X���ӻS#���H�C.L�W,�nn�2��w����-��3;y��ѧl�Ԭ���Y|�9W��ɹ8�ݮa��=�=�	�܆�8��� (
�G��}B�&R�Hb��u��)31@^����c��0��ih]�*J|�Iɾ�<��&���B�jy�=�}P�
@�=�`�CuS���i��C�j�k=�	ӻ�#���"�x�@d�i8�%������2r��&}F
g�L9d�С�Q- ����C�+�C���B��KM�`a�g��u>�e�����[׳Z�3��ګ����)�:��^��y��f�S>��L�Ԕ�:͡�)�4���B�������>�m��F�1�3����5�aI�) �O�a�y�0�Pw|+\����ֻ^������[6��I���L�i�G}���R
d�\8�CI�-���n��,�m�9FP8��Ч4;�0���K�ai�O6�����A�&5��0�Jw�gd������Ø��E��Hx>�|�ԶM���������uTB�e�n��zÉI���&�}a�I>JE�Ez�0>i��ʻ �@Z[0������Ka�b�l⤧̕�{W���O⾣}&��=ϥ��L�.�>��<�R��k�ĝ����Gݳ��C�S	5��PS̜m��\$��M�[�!L8���2��Q����<�N�1t)�T�X5�E�Վ��sֽ���}�*̡����ة�T)�a���l�̳�[/�E �����e8�P���f>�y���0�Y����IOS?�$��L���]�)'Y륜d���S�w?v߷�0�1׳�&�}p�v)_��q�T���
�2S&*�T�B�wd�q�a\���-���S	�a¹�C�R)o�Ĝe!��Ϲ��)�4�tg�@�RN�^�Y��Q���g�~�vo�|6=�}�@���@��̙mW���n���a��n!��L��:�I���.�<��1D�����us��L5
�8'��i4o�I8�&��a\���Ng�?E���������#�dLxDd��fRh%���9�CII<�Ͻ��ڤ�2{�e��!�ц�yH7X�'٨u�!�L$>��e �(��>3��AIhRP}گkkq}��h��eeӁAm���;;��5��_>�@�:
bf�-���V���)�� ��[o���\ޏ����n�1¡���;�����O:빣V�lK�8�9*ʩ�q�%WB���+�`E���h[���]o;���1�L������x�V�7���W*���H�?����=�����2�)�'n�}�R
`��:��I^�>�[�
e���Af�/����R.n����uI�P^jah��/d�2lK;��<� �\���]�7_�n�2Z���pL�`RL��n�Y�O_��qk
aL�#tf{�C,�%0�Z�M!L�{�0�,�l0�[ǰB�e�KfyB�&2����&�ר9�Y��u�g8ޫ|�ވ
 �Q@��M2��mp��ԔŞ֬��|��E}��]�-tow�aI�O6��������:�aL��פ˶JE�I����(�d�\y�
�u���h�S=�o| p=����B���L��qD�y-!�]ͤ�i4��4b���a����ITf��a�T-)'�¹p)�T��2s�QH(u3�Xe��l748��
<bg돫����_Fϲ=�g�,)���O�)UL9�
)L/�	&�Ʊe2z�r��O�a�&�F}���l��&��dR
C&����C�+�>��ɖT)�gsu���a��6����Wj�t
���P>��4Ͱ�R������mC�d�T>ah�uA����7Xi<�h
)����Hb]C�'��'�ja��S2é������S:�W\4o�w��l���'��w��wwu�P���$�6�3�����S3�ng�	��}�q4�ФR}z��e!i�ъ��IL[��O0��Hd�
�����1E��o�_������
ҕ�����|�u�ZN�I4{��$�aH|sL�d�Y�>���@Q|���o��&����T:�z�S�b�'�Դ��$�i0��'l��)�(� ��<uzo�r�;D��'o���<��xS�>�BҒuÄ��*J|k�&H(g}�a�!l���1��d�*C}�����7�Y-E:�z�nR
M���̧Y6ߨ�EC�)�=���v�|iJq�f+}1ܹ/��c%6���qB�P,��VRI[��juP�`�.L�[2k�S<`g\�0�
N!�-Ѿ�}P�E5;�Xa�Hu�߮e�!��UP�~;���+�C�;��*,u�o�]��9C�p��fT��ei�l���0�ĩ%Tp��y.�*1���a�״���k3�x݂8��:�G���,�w/x�[1g.��o+�s\d22�]��9�4OY�M���q����)�f������)!=X��_��=OX��rÈe�d��������
e��F�B��O��UI�)�
���6�����ٝ}�a�u- �Mݚa�:�"�z��M���@mMOs��W����K��d�������[@�S��nC,�%��h-aIl6v��N�L��M�Ì)2b���d�YԶ���R�e$�C}��M��D*=�D����f&q�}�8fv�+����D�|��ڻ�I��i+Y�$Z{�r�$Po���i�٨ZR�v�&�-Xfv��%"�R�B�ߘuC&(�U6��T:�e�RR<�R1�C�x>����"��ן{#ޘ �����:� ���n��m����s�e�XS�O�F7��:�NS!�\9���>��iYHZ=�3�!L-P�=�a��Ae���C�
�=��
�٧�=� �Q���00���5��U0�Ʈ�R�!����e�u���"�RS���Цy���>;�,<����Q�&��y���aUIHV9d-&mG��O��k�on��1��G��-��)�f��31E�,<��Ф]b�['̤0g�u�T��.,�u��eܛ��'��}���d�Xa�'��Pu�L!L��c�,�m������O�w�;�6�w>V� l	��z�g���0���b��RZm�2����a��<�Kg�jKg�6�L�}fH,�׆�) ��.M&�{�JO�zÉ���+>�k���)Qe�}C����Y��WU~?�q%?0��9���Lb���2�ɶ5S̔���vS'ͤ`��C	�O7ڇ�ja�
|ɓﻃI�d�S��{T)�1�{�������_}������ZN+)��݆wD)�����aĴ��fY�0ϘR(h��L0�
L!�'*e �h`�(��)���)-�y��d�KE�S���I�)�dp�.o�����o�r��u��zB�m�3����sD��3�{a�U'�$��e ��:��Pq�7D)Oz��&�m�KI�˰Y�KCS�����L���
y$Pf�,Y��d�oZ�u糃����!�.<=��f|)ފ��@M�p�����m����/))���N�C{� uv��c�=�do���p��wVe��I>꺾ZW`x� �{��.���rc���h\�g4�t�<	b�ev%z�ٻ���E~� z2ݴ��;�>p2�1�S�~��Qa���oؓͤ���_�Y:����@�S�JGG���L�(�M�é����݇3R|��þ�,>aˢe:��L�Km���
~*U�û�Z��@P"�@��dŶ�)�������B�S8�m2�Y�_s&_2R,���P�J|��n�dT�'qG;�a���{⧙)�v)�M6�tc9���{��1���K{�&=����1[>���1��a��(�Af�fb�4�ۡH-0)'U���%n�S�5�`2�0�[[��g��y�"�r���Ru��(a �ԭ�}ε�������ߧgXR��>��)�8�l���0�IN�v���B�l8���S���P��8�y
gqRZ��S=��AIL���[0�Q
r݆G�����}{S��=j��8O��/����8�ih|�Ũ�N�>��%�ith�b�'X[
�O&|�3>�䪘@QaL9tS&�I�)��I}�d�l9���a)�%܈�8�� #��ӟ[;����M���3�2�$m�C��6��=��0��8�|wפ��$�n�w�"�P��\6��ɟv�;@i-�;@����i7�U%�d�Xb]B��zaǃ����~����s>��j)lzq �=|�!����j�rw5<�L5���)�N�������Rq���k�,6�����i ���XS�O����]�$�������<& �ӗAr,��]u��舀{c� S'�R�L�ΰ���0���C	5���E�aH�E�Ĕ�8�}{ a:��&���I8�3��Ǭ9���0�>���f�m�e��l)q0�լ���ݥ���� T<r�H)*Ϯ.i�z�g�ϒ�y�KL S)�R��[��)�;��!�����W%1f���풓	<�3\�㾸iE�������{�h/�
'�.�.�B�ܜm'P�w!��Y0�2v�0�R�0�t(�����7e��䴂ຆ�jM2�A�&S]^�Ʉ��$��y�$�)���I��& �ee����dUG��MǮ��FVD]�|�M�ʙ4�
f�w`=���z��$q�ϡ�U�o�k���i�(L3d���*����RՈ�W�n�k�K{��X��x�g`8]�X��X9�)w9�b�j��ʉ�,����#���(�Kw�U_}�|���m��y~�����ݑ��{ \-!���'�%;d�X���4��C�א�A�L0�(sP�
@�R�>��d�}1P�S̟6�3�(Ri��>�r<&<xLo�H����ӿ�yY��s>�=���>=�&]2v�Y5�\�AI�Oz��RV(�&����nk՝&¯D���A�!�FFG͈ݼ%85M}Ӷ������Xo~#�K��z|%�g�d�o"�f�IT��ڲg�Z�y'��X:�a��j(]��ķ=���Of��2:HV�����{�I�T6I����:B@�O}Ԙ�N�����C������^ç ��͌�"�\�����Ϲ�c՜�C`������+ƈ���}q}W��3|:<e��ك�EE�e�0�Z�nH��xFC	"��ףj�.(ht���(M�t��
;o���ڸ{����8Y�����V5�-XN� �J����Ǣb�^�"[���*\\��:��>zy�<��D�k��"��\�*DWK��ٸ!�@F$dʯ��8�L�An���o��vPc�֊�oRʋ��U���Jr�)jf;ؖ{��#F2����c���R�Zh�&9@�L�k#��W=���6\\������{[@����ö��$hݽ]e�ښA>�Ȑm�NTV�3��P�wҲ��u���c��������Wc'+�1�G�;y�W�F�S�F�rrF��.�:��j�=ڒ7~T �����C��mw��J�3b� �"�x�W)�6�T?ǡ�ܝl"w��U|_^	w��DoMC�6����30磯ƎI�q̨��}8:P.���=֩�R�+��y*���r'��J����p_��"0���n|�.�'-��TWoTV�QG�0��N�3��.��[>�UD��Q�Q��~�T�h�ˣ��^�w �n�����0t�"�\�R�N�M�nzh������>���a�{K�s�3�SFE�U\tJ|oh��f��ķ�P��{ ��75��Gg�!����2��[Vj�WK�"`�(1RNv �Ʀbc�s�ŀ��� ���'П�=Mޗ����jn*e�����I�ݛ�`T�0����s;C>�>Xjq&��y�d�m'�~����Euz$`U�<���*����]C�s(B�n�]Q[q܋��.��Esw}!����i8��!�򫢂1{����ȉ��b̞�>�չ}�V�Ca��}���X:���V�
��<�_L[Y���V�c�٭�Es^�T7q����F�����YK�f�*]IE���Y2.�Cm][� ̰�엇��wnM�����W( �t�O �����;D�w������ =�vV2Ӟh��YU�cY�-�8.Er��.�`����Ҷ��)W����|Z肑���U���5(t_3'`;�N�gQ.�3�q���^Ƿ�h૳$tk�N���Sm��[WJ��pN��1B��ʠ�e�y�*��uZt�)���b���P��d�/��J�h���FFѦ=2�tO�Ď�4�P����
�QS�uM�s�'R�9�Y�&���p�����S���鞩y螉��]� ���NhR�{Źlە[Xȼt%N�I�\����/����?/MXe_*`��Rૈ�:*>Β��d9뷆x�"C�/b2o�v��C�ړ)0�t5M�:�
�]ᘿbv$�#���Tƺ\l˽��s�$u�މ�}�q�#�R�Q<�L�x��Q]O��~l���N$F�BpNj�9����|�\���{���{�-��_"X��[-�
�����g�..�4��;�: S�gs��~wn�����W�K��_U?y�u5���k�����7��9�'�Q����h
o+zerȝ	�2��{�����K��րp0U}�U �D�&��}���W�,62+j�I�#���hayN�����F����
���e�����/��1��z�Q)74���C]�L�QY��v�éH,2g.�7j�!�]\A�I����u��p�0]�1��@�����J^���T�KF�C�a�s���y8�D��N�k�D�Q���֚C�&K�)�lo`y�l���z��
!��eelF*b�^D
�4��%D-!�%0�极<˖�������)u��g@�r`���It\�����=J�k��$�^��-�`TwBsԯx�>��r��A�b䯯�#���֨5�q�ڝ$3gb���O\ޮ((�л�=a��v��QSk
�u��y� {�z�-��l�x�֤t���E.鳤b]��ʮ�Q�v��A�ϫ����)X�E7� _'^<55fJwS&ߊGa��FN����6!ׁLw���4��`jZ��I�q�Ot��R5z��,�tq����s4C���2��m�|��|�j�jD��1@_��R��oG��,c��VW.��=��YJ]n�uwW*z��2�����+E�I��#9�5Ձ��(53{`mnL��-U��tw�p�7�rkߝ���)s� �V�T�4�̔EHX��gh�u> '�=zR���m!�nP�K%��ɭQr�`�:����w]�Z�����Ӂ��v���XdK��e�����Gb�5���^�v��2�m�ٰ`������Sw�Rg0΢� 8ܡ��<�Ik�ս��z�l��>�:�G�;�W9֛‱ُ;guvka� ۋs�;��\ŽxQT�"NrR.WW���>��y]�g���w=�����#�31�:���ki+�zw23�#3v`��\��h#�F�V殕.��:g��e��u�H��Cn�21��N�7���>%�պ�r�x��7@��O7�(����i�*��wI5�*�G�߹9�]��:��%�i܉�mrR��We�o�\�����M`|t�T2F�6�죚����5�CLa�𾐳ܟYF��;�]�]���ʛm�u��+��Ku��ׅ�����07�N���U�1'�p�U�c�Wj�{�
s�[Q�*X��@N�JMi� !C��w���i�1�Ƙyxkc��"L����sT؍v�6�Cu��a�0󡗥����
��W�Z)�d��CZi�A��"�@}yk)ڷ'qe}\��͏:l�*bZg&uΕml�;�mv7mgY�l6�i��	$�fI��6�����d)]�+m��5���/ �J�U�n "�j�(]f��I�A�ƀ�.�N��62�,Q��ۏd�}��:f����I؄k����1E�R�,w`
��u3�������S��I�U�0��;KW��ȕq�2F+f����ѳ��]T���������r S��9Ŗ���kN�u��E�؊�N���s�6�@��IY�;���Ds�C�t$f�Q8e�f�'@��R��wgiB\uq�$�e;kve'6̶��t!��rR��\�ӄ�q�t��g`�d莇�����9B�@����$�Rӈs�YdAP�QD�Y�5ݵ�� "��#�8� pw%�jVۜE�F��R��̎�"m�f��vv��N�I)'��	��H��s�[`N$���@��A'h'���� ���	�PvY��#�$q� �R[j�N.A#�9"��-�I'gaH)��<��{h��t¨  �@Pwk^�tka��o�sS9�# r�N��R;�&3ԓ��er�m���pl�������e�].PW�ksٽ��..xxx����!��b�:W�"EE�)צ�²Qg\��>̯I�B�wz����Ms���Vؾ��S���RCC�@�vV��6�^%(x1K(�R�"�J����j�:��[z�j���˛M�6]��wVR��X���C���V��x����yFE{�'�# �"�����������ea\�kK���l[��H��aȵ8E	��zf�조�%}��W	{+�tp�<�'r�ǫ33�yrPw)fz�v{��p,=g��W��#�˙Β��;%1(Tfj|З���L��] ��d�S���gQp/�!�ob�5I��2��r컶v��k�ؙ<���OC��z�h*�k�i�]A����Un\�S�HL����ge�ӽԵ��	oU��2�Ñ�Y�G�h��ؐ��Z%WD�:�EDm5b����{���a�el�J��㾙i�na����|��t4z�좇��,c���
����0��1�ۊ�,~x�A�g>�q�a���c�F>�0[�sOT9��t����"��^�'i4��>��5����;�	��aD�v���n��Kּ������8���`�օ��fP�+9�{�w���������Eu6��:侩ʭqxMѦt>��7_L��V�bp���ݚl�s7%�{Xf$�ܽH�ю���D~� {Ӯ�6�&q�;�'⛧���:�p�ʽ�C�x�}�����!/P���gX���*1�ߠT�1�a�J�>���T��5�����QcTWCS��WN:�����hM�99��{�]f	0�\LK��+!��nl�4/kā���5T�;:�]��bRm��>��Ng����}shK��t���a?��(�<
�c��*o�&z4�<�x����2��ۀ��ג���I��;5%�b6�`��B��>WְW��j��{�䨣-��N�(��QP�>ǂ��r5��	WECM�l��M�z���A<((�]�g���}[I-��2��s����^�'�ၒ�\�(KI���f������9��&� ̴\�NY�Z�})|��;��u�E�g��Ķ'���9�0�&GA�+���ӣ'`]iέ��@�v�Ň�P��5��e&(	�\-e�^�reqڨ1�t��1��h��6�n^t�K<���S��qX�=mS���,OƧ���~ ��}��n��u'd�`b���<.�08��~�'W��Ծ<U-����u�F<~���^�6�$l;��S�*�ߤQ(s��lZW|o�w�b����QpC�;�Π����/�Y�����T0�n�1��]3aU4�.t#��N�;�����{-�Y�ʲ_r��ϟl��/:��6��X4�&���N�!8)ҁ��T���W�ۗ+�K��ݡ����^xu�ZL��CάR�zꭉ��6�R%�<�W5*�*��+2���	lP!�w��/��	���V�g��ARq�֛��~����6+-W#�(�I�+g������5��t\���*��h�U���1J�jf8�=�Y��mMek��ٍ�X�����NÙB�H.H�^��yN)�"��ǡ�~�J�r�<�͸��zgXt�A�7Bo�J����*x;&�"�*P;U_K���~r:쒲Hx9��{a���kC֙8D��H�)D�UP�k�S7y\&=9�"K�<��q��z�gLS�\�,,�sb�e×3b+Cg�)T9����nR�LԷ���	��S��� 	ܣ_%n01����
�	�P�Rc�<��{�M]G��
�{�A�<o����5 �B���6���ٯ7��p���P��$��AN���C�sO޸ͤ<n���~�S���&���%����N	�h>�I���f�T�|�k��Ӣ�u���R��^�V��^�i�]դnT���s��4ͷ��}-E�J9����G5_eh<��r�M().�
H��e�2��_D0Y��պ�N����Gb�J�:u���3	]�#��{����RB)'�}S�6�<+`P���� 3�.�\g�ڑcv�6'>!ۧW�9�?|v~��߹�d�3�!����|��.��#<\<*���F�����'�Y#{K'�����^�|���Oq1*�� ����\-�hx�8�ehw�Tw��}1��4����H�ؕ\ض�O�
]���껛�o����eB�`�霔e��R�g4R�����a�zd�t9�(�#nVx..-Ȥ�C�9��k�
����#Dt0lP<����w���	��d�
���E���炚�W�v����E��J
��j�}/j'hdܸtWlI��\�;y�)� (�V��_�Ez�y�M*��)����u����~�:��g"~���t��
�ݬ�Ȗ8W���!�!�	��
�T��X�dB�5��]̬������2��E��鞩b:'W��L���Fx`�E��
D�	�*�J�d����2�0r�O	�Py�̨�|r�����PRฌ:
�K�l���y��i�U����>x6S��!�*�L�m�[��J1����-���S��5Nc8�&"j	�l�����B(�F+V��p��R��������VN��w��l�%�zc��n�K����:�Z&�U�U&��<'t`���������籖9Y���7
����:.BSqNF�Nn?�xf,bv$�#�ъZ���鮛/.�/�r�Iƅ�][���ǈ��ƨ�s�ɗ
+�>�u���-#/�촯�o+��hc�t%஁^$q�%C�c�~�+���t#���..��p樌Z�fZ:ts��K1��]��9U8�}�tYK|_Ⱦ8*R"�l�7�Z��N-ʇ��,���8r��;5�8���9��)	��n���M��p���Y�8��̯Mv�W���btJ���نu�,K��V��7ίMX��tFJ��xy}���(w�$���kG�%�@�ۻ##4����B���b��}"�OV@�c��OP3���"�	nE%Q婥6�R풒20NB9��b�u�n�@g݇"��ECE���:E��r�Z	%/j�(֢�XqÈ����]J/��1P���T���F��z��U�'��מ��(k/��
��G�7�ivX��O��
+�2�����Qp/�!�ob�5]����uV��ʾ��m�h[�n�!]bh��p;�LY:��0�c<�%+z<2'r᧽H�̚��v���T�����Yo��£q�U�GQ��+Ժl��Uv6_s]
ݭJ
ڻ�D
W��1d�w�֦i,#9:���UU_Wǳ#Sy���Q��vU�<���4�X�?*����ᣜ������-!F���=��k��򾓨0}��u�a��aJ-�K��[a��[PB�*�,��D��z��Bo�k��V��zݣ89�9x��w�#��2/�y�~���C(�#��U���_fo=/#O\��Ko#�=E5u�������
v=�X�nY�}FMW�3bta��'\��}�#S��S�'��E�T��q��M�g��>�^_	z�F1��o��r��7{��ȸI���Qѿ�GQ��+�p��h���E����),�Z������c\��9��z$��Q6�d"*�e��f��x��-����{����N�����[/wyA��~n�L�V%į%t��AY��`<%'��]4<T�:���Z�#bcvk&�RW*���P�Q~�Rerf�y�b6�`��d>�T�B�!�Fi����{�����Ed;OEA�b�x9r9��eB�l�yL.V���<i%��q7�͢z�bDf��Eu��B�WJ�4�#(Q|�:���bW;����iT:���A�۽"��q�ɬn�W�䩫���e* �4ڕ#�V�*d�0�W�hZ�#L��L��-�:�Q�:0��X8��Y�����]S^�.$W�s7��.�6�8���x�_$�U�ڽc���	U{#.���F\��6��L� Cl����x9��&���O����oE��o����}T8RREN@.�C!�v�����:�ÞˣS#���U	3b�RK�?S��Q��G�����v1ײ��Fzf܅N�GN�R�T�!�[o/$:�K�8R�V�\��lXO�`�u�U������:�*t�?���F���j�A�b_��Lyw��9��#=3Y:�>.��NA�l6���c��6�Mx?�'�@��1Z���Gw;�]p�������h�p�f)ʽ`�V���X�W@��#�1Dm{�!;��=uV��=ތ�)���@Z.&�"b�Br��r�\D8�(w&� \8퐮�Zq��]m��ݎV� ̰��s1�:3¤1R"H��=������w�K��{��c� �~�Lw�𦸬Ϊ~]]R/����c�X���\�U�w����"���Ј���T��gNg}�����2�C�j��Л�����UT+���6Eߣ�QGɪZ):�iuK�-���(��J`S%�vwVD�l���;]\ �ܫ7�9�k�@����$&�D�ǟvX�Y;/�����Y=4����1r\`t���vK��O7����K�f;��x/*�HV�k����ΰi���T��ApJ�"L��9Q�\�z�r�����zq�bP��k���l�/�@���K�����8D��H�)D��
 �+�D ;���O���힩Гk�XW�Q�}|n�r�W7O���:�G͟@����o��ig%JŽٞ|^���)b@� ���k��1��u0T�!FחS������4U��V��o��.Jì.�"v劒�;���	O���ڛ���^B"��F�9��fz�2����zծݚck`Ԑ��P���5r���
�G"��ԋݣ��s��4��'������;z�L2��~H�jO�򈼣���K<_��*#<_�
�m���
�CF�����t�k�|����g�=���*Ai�m��o�<|�̷x8�׮��� ��No�Z^�ȱu1�� ����l�͝�a��V���+���WW�>�ƞN�ч�J�������p���^Q�5r��qns�S�D����_MvW�(�S�{�Y�)��kY|;=T��Pՙ=�J*6j��k�^�q�p;E���N) ��{�n0OEt�m[�5ۨ���T�̓Hq�-Tj�K
`���FD칺�w��r�����i6#Y���|�0�ܑ�����z]*\�f;]\99�� ��;ChԲY:��w=Y;�M��"�Fv-�K=}�������U1��X��<3q�4�׮�n�@��=3^��2D��$!��/����)�aM\5��ִ�-�X&3�޸W�{s��c���1r�N��_Z�]C�_�uS�чÅd���5m�\�m����u<{|��C�t+�T�{=O:g�}`�=��֕Wf��\��?K�^�bh�W+�}y!�ە˫�G���k	�/���H�K��"��j��w�l�W�A�z�6o���;	�ʇ�X��r����6����xf12$pU�"m�I��]t�{����*w�QNR��ԣTO9�.:�r86����wAv�wa$�=�^=�o hz�^TV��H���St<T<y��;W�]z��/�EU��Yff�/Z^j�q����NAu�8J����R���1�@Ȣ/��&���s�7��Ԫns8���Yk��w(�*���6}P4����ipoiX�W�x�3xn�Ӫžе���U�u\�'���������Ls��
yZ#߹�����h��c%A�ec�Y�q1C�P�a�4N���T�����W7#�u�Prǹ�hc�;= ��.�mŽϺ�l��a�]"R�l��8�2${��ie�76��/���Pu��#gT�;AZ�*\�o�l���V�i�������{Q��X��7�ξk���gJ������� {z�3/�FEm�fڿ�,C�Yse��� X�Gd��.h
�
flq��n*�%oF%��gK����,����g[�%@7�r-�d���(���2Y�.m��핏�v�` �dzT߫+��W�0lOE�R
{9��5�U�t�oGWS�ճYs�7ܦҎ~�t�9��$G��PQBT�6�!gM8���l�Z�J���3O���t=�X�_�vTA�������S�u���]A����;�h���T�N�	��A��`�I��/S*1�	t6+m��+c`�B�*���U���˝:�o��5�&7%EC�nٞsn[T�1�L����峰X�FuF��"����{���cj�n2]w�e9�UT:=^:��X�;Pr�ϥXnTl{�X�!�w4�!�Nbr�Mq�a��r�����g>�]<ty��i��~�U�(xh�-�`��]����ޓM�x��m�)�U����q x��ia+�S�p��{��p�}��ʥ�" ݧ�*��R��ɩ��6F�5쳜�7yc�}���V`F�@���bjw3+@��p@�R���U���6:��w�L�vk���͗]3��zζ�ӮQ>z!�ӏ�vjk)���6��0�smm\N��)�]R�m#5���U�˴8�WO�\Κ2�%`!}���̚J�h�w
�Ӳ�1�&XaF���-��d���R�U�;n���.����umQIeE��I̝Pf��q��˷"�)�e�j�(]
2vN�4��ɬ�%�U0���d��� 8,	k�
6��rp�l��'H4�Bv�V{<�zoZ�T7��S����3b�����pp}��ǳLɸ�k�����m���m7Y���Q��8ŝ�)$L���ow
�I��=ZwQ�f�]j�u{/QފƙQtI��܏���dv�W��=��
Z�g+Dp'/�;�cC���P �K)-�	��][���n�P����z�l��Gu�;7��ն��;% ���gQ�]�v�8�A����a�+�[�|�3�s��#���{;$Ӓ�۞���VJ��e�ʽF+Q��6�Ԥ��jRc�V���:�k�섶�YS{�q��a<��RAo<�ř�D�ܺ\>])m��eG	Co�v��hFh�]`;A��k�.��غj��Z��o|V3��8.q'�+�Yi�\�pt�dY�z"��vçm�hq;L����XlU�o*kUm�Ԣ�Ι���=Ǎ��ua�zG�Iv^�{��
�U���J�K�I��"�)��]�)ԗ@.�t�w��ݲ��}NӬp�G�<��9ȑe���*)�}�b�=��-B9�+���D���r\)��e;���!z��M���7�+����!�+�w)9z�w`�Kr3[��fv�����21b@��V鼼���B�j�ھ��w�Gi�z��7z��8�+��H_Q\���e�4nr�3]!��A6 �h��n�)p�]0�,u��V�f��`S�}pV4yj�#k57�2�S~Y7��2Ni��=Ӫ�+17a͚Mͫ=���z>y�:6ۙյi��'����C�t���mb��s���*�A�{ʔLҤ˛��v���dVv�P��m�z����)n���.��-��H�vr��6WE�V�~]����g��,f=;,��%����!�Rw+q!u�;����[�4�_�3��u�%}��+���(M�S6Z��h�i��暂�ǜ8�B����}��H���}�v`콙�:��-v�Aer|�*�ؖ�ES�Ns=�go'2�iu��,3������Qm+���W-U�ب9���ym�]��>��4�(@���m,	�}}q[�#��jB\i��YtR�h�M���pd	�B�L��
��L��ZN�l������[7S��o��h��6k'5�N�u�檱�p�͢�*�b1X�s�7Y�	��$G8 $�c��W���ԗ(�v�(�N��$y��s��3q�\!*]!qA�6��J*N)9	(8��;4����iX/1
vv��6�(�$�����Y8:e�q�jE���(�8��E��p�v���9罓��.!89� Vi`��(�N�����ډN�y[��q�9�Qw�dB"qy�R)6�p�*Nf�;:�R��f���,�9֎V�D��Y��ol=���#�Y!��W����C:.���m�=�zmI�w����+N���,����=�x�NNH{g�r�ז��D!���z��ۼ�2�^��2�����m�����E{n<�∦�QEeT�Pm����ɑK8n7������ja��*M�ý�Zb�w�nߜ��ݸ�dGݜ��fwp8��/�I�r;��g�_| ����j�z��T_�M^Gg#z$�C�4!*&��+!��nj!I��o�n�����V��/�s��^F�v�G��:�]��gå	���E��a?��(��x�i�������Ȱ�ݩC��s��ݹ�)�����T-u&W`N�Kr�d�N�\)EG�:0����d(24a��o�3הtVṫ��/J�ʊ�v�|�a��QPS@�N�d�W�fS�gZ7�{��3��Z��)�UZ�}��ߔP�G"�]˃ct��3��PC�ق\��:Sr�^w�l�߫BW�G�B�r���JEÍ��>7Ķ'�uy�&%���_o��__�Z�b�=�����^����xXsT'+�fQB���5�U#l��CL�K�x{��K�1jJ����J\�h�aӀU��fŷ�ltk��+j+m/�*��'�Q�����Of���)#�ٙ�&a�Noj���L����C�##[EE,}UrN3��V�
��=Zg�;��R� �t(�����3�k
���:�J���#�1��&���D���5˧&%'�NDL`�m��۾�ݦ��P���<���V�YWI3�=����m����� ��8۝M�%��fYx�QoU�%�6ݲ��n�%q�BʝE?�z��|H>��1y�;�����Qt��V�*��� <:��r��H���P�=�ȉ���	���V�C��S���	���]�4�6qd��Z���ć3CF�)"�q0�)$^�ʋ�,#��|�l&)B8���u�콞ښ���g>�^��|�{��pQ�v*|�T�%`�\�U�w������"��y�1ͺ��tu�	ks��.��ų�<<5�rj���«������׼Ū5��`���}8�<�Z�H³p1IS�%O@4˾�~�w'��Y�#��J򨀢��(�oO&d���o���]��5�W��b�j�\��曢�'�r��W2��9�K�$6}�C�;^಺VM	9{�a�-!wp���ː�=��]���"���SJrs��r���G�%�y���[���H���4N)�*J��U\dn}F�ڛ�o��ʄE1%�j3\�R��^��ꥐ��G�:��W��.��S�8*��m�"���sjE�цę�Z��/�����!��Q1^쳰���jO��ԟh�{(?i�u��o�u��z��ű\[d�];R��m���k�׼c�i��;����{"�Ԝ֬J��
����7n�	��ݜ��8�^o\�x���$���.��� Y�q[}� ��0Q{ɻw� B�f��N��/s{Ӹ,��p]0�YZ���;�-#��nMu���{��V�}���-�}jaO�p�3�|�t�w�A�1�GW�F
Q�*���*�M�ܙ�*��]�VîGo�cB.�bq�.���<�#y!��f�vaϹv��}t+(��ӥ��v/,�`WV\�5�U�ըQ�گ(���x���8 �@�^u����ꌷ����]�Bk���]�=3a�����Z�����^j�یs�v��g8���fN\౮ONcD#�L�]�`eP��:�HB([�3}ET�uZt�I��q�QO���t��ԅz��)U�)�3J�6'8W���!�i�i���z�9	W�b�[;Op񶧯�!o��bT,u�!���jp:g�^�w�G:J���K�WPӂ. p'K�fV"�Vr�_v�r3�6�@�]^�)��\��C��*o�@�
 l�0�����W4�5Zɜ]����l(ء�]
,vԘ	I�]Sa:�
����&D�]X4���i��$e�n��oÐڬ;%�j H)@��b��<�.:ې���h~rb��
X&���LQ�٣�v���X�ȥ�gvQ�ys>��3�M�����g��8]֨D��V�庮
u��Z9N��q-x��{�^�k��s����S��e�Spi�sn�T'���͖ႏ٣>�
Ժ���J4��ڋ��3f$���K|�:]�k3W޼.$AaP�B�Dl��hx�x��?x�
����qb|�nŭ�a�>]Q���C���ԟp�CE7'�%N��T�Mx�E�-I�ֆ�n���Mmf�3}Β0�\l
���uu:Ce�EE�>�^��J	�Y
&�?�1\�:����g>|�G��s���v��s�C����3�NBm�:��-��aśQji?k��z�k!���l^m��P�β����-PV}~Oz�����>#��w[���Șv%)��NGf�h[��$@dv�S���ڷ{�b-L��s팆���z��$F��1r�h�gԦ�)Ŭ�>��e�=2�=��ÁoY�OSUʕg�lV���zFU�}���;'������2���k�V3�����{����I�S(>�='Ƴ����(��#�r7ܑU+=��4G�0��')0�r�UI�=a(�����cڪܸ�)ʽ`�V��K���ح�#�4���A
p�
b�p�7bos��:���s�u����xb�L�ŧck*��;�Q�q� ތ�E*�Q�삝:fC��l{�ky�X T߷�������uݾZ�n�zJ�}�)M��C`�Y��;Y�݁��5���l���S���irg�����Mbk12��ؓ<�EA���fy͹} V�w�#��\�u�S�K����y��/�Ol�!�cԎV����J�|��s����jg>�s��ͅ;�|D -��{�8��./g'?U^_
�S(BV	H�T\_��t(�T���x�e�^�o  gk��}'WZ�&�S�����<|s�Dx�h����>�d(��+���z�1:J��=Xg�V��⭱����E[���m�>�(KR�����/�ӵ�Y�,Eh�'ng_��4���S �޸�����˅b\Xi]#�PWG�p�j���u���78�[��zT��EZw��ބC��Rerf�[�# 8q�&��h�**�Ô2�瞣�]����F��ʦ��z\TgZ���ۑ|�a��QP|�L��)��E8;�|�#=|�ޡ�;7~'��4�ҭX�ޕM�aT����=����[ $��Ǖi�N��1ij�w}���I*���h�UX�䊜�T������P�gޯ��	�$y��N{�����6xl��t��p�E���8��v.�λ�ǄX�8ᷜ�����x�t��n���CI���s���7��f@��� ,I��8K�(�c3x�;#�݉K��L<�
���Ю�RA�Ԑ3�ݦ6
=�WV��՗�1��r����dt>��N�9���ɺ���(T�g�p"Ѱ��4�2����b^-�	�����
us�^�X.þ͆��F�t6���Ț�N4�ATm#o�j��b�Ovw q��Ɗ���!)[T\�L��d' �y�61�TR�4�*a�@�{��s��Ӥ���ݻ{�hz���N��5W���\�5�-&\{��V)�U�'��νY�7�Tv���a�^��'�P�z&�dL_HN^ė<��ARq��$��;�����0�ӑ�u��W�L���A�bR�)'׼��a~>�Xn��ZIGJ�β����1/�a���U[t��E��z6:�R�P�2�ѧz�KyO�AkvV��^�}Hfs�\���qP�[�ru�+��\�ZF��x!U�W�xd}�9Gw��M��9a(hܥ����ҁue�B�gr}~L�"lBr$R�h*�
2J$,���mj�N�@eI`�lڗJ�R/ڣ������X!\ا�n2���/�
x�^��	�6Ma�o�Q0�n^dN8*�`�i��L���V��
�����l�MKQ���睹���Vd�`q��D5
�8׿�G��1eS��3�R��hu��K,
Ͳp��b��N��S\+.t��G��]�7�i�rc����w;�:��"pul~hd;�.*��یS��s1Jx'AA�ÎN{���
뻵Z$D��A� p�D�RjK���� 7>��jo7��x�LJ��W����^8�ry~�>ϕ�}�F�JO"�![�3W-�x�@�.���xV"rm֚�6�+ۛ�~��.:}�!~t�b�Y����jH�WR}�\8V�"�vn��sHL�me>x�t�ҾZ�����{�mOF��B�>@�V�U�Oq1~��YZ��p�hx�g$E)t�|�m�������vU�3�q˸��8�~w}>l�͝��E]`7�ؠ�P4��_G|�@����ŭJ���W�V�FmW�v�.Z�qnpAN�����eC��M�:hGz�S�5�½�'�:�	.O�ECvd�yԭGMS��'Ϟ�q�_,�/k��t�i�}��5s_93��P�p����;�pSs��A�n���Sy�i�̓19V8���n��[�:�Wŕ���W��>�
ןa��4b�(�m/�Q����ܨ�nAQ��X5�z0՝z���r�>&h��W������v�*o��yh�W��]��	y����G��p�����l�WA��zc�ȪT�fj����gF\��,���:�u ���=�Y.�yz.����VAc��+�Ĭ��p��������´}����ٝH+��oQr���"�1J�YDӯb�8ߗ���|pw%U�N��n$r֮�}
��ۙ�Q,Zv���ٷ*�W��'aA�[2��>9S~�@įJ��k|���5���a��$á=�U�BT8&7�B�V��w!)���j�N��=	Z��u����{�o���^x����^��i�����}Y�o�`L�x�}r�qUD���ܝz��b���k������l���:A
����C��Q1@��=
�����Y75Џob����c6q�ˋ�*���bU ���E�e/x�E��S�E������U�����bV�q˺�`�'��_K����]AN��xH��]zhp���:����8�T�f1^�^~�I�G@;�v����1`K��Vжw��YC��YG�*��ܖK�^ah�[�>}Bȗ���Õn+z�vS>>7�҄;�3�Ŷ_H��Ր1�d��zz���3��-��.�/�싊%)>��92�dnu�n����R������ǟ�_=*�h�8j
z��!���Z�Y�)fZ.^ެo�=�� �ʾ��u/�X���;�+����q�
�ŝ�b�K���X���^��nX�;��<��+��+���Qp��[Թ��ތR�C��z��u-��Wf�S���M����M_+���Y��?}��4�_myU��Jׄ��A|Ϙ���AN�#p�01`5.k4�>�k�j�08��'��v�����zf����K�l��z�p�u���p/H������Y��l�J�t������à��W�$<~Tmu��e�b����M.SP��������ˁ���k
���
����<�D��������"x�cWj���& N$��**��l�u�^yP�;���.x	l�0��JWmwu��1�G��B�����4a̅�������s�E�Cr��{���7�����o��g	���5�z^��S,BV	H�T\2_Y}��G�\�n	ҽ�p]���NF1�n��rA�J$A	QKӪO�<#KWΤ��p*�,�>��q�m�7\����GA�)�C���ɹ�X�|*�u}Ԭs��x�G{�p�,@�S���z�C�/U��}���ߵE8�����.�qa�`�#��?p�XG�vz�d{,�?
΁-���l.�9��sfY��N�ie�.�m�cud�V��A�X���5�e4��Mݠe"u�U���u:*�7%t21���a�ך���a�a'KU��r��V�}(=�����/z�T�w)���S2���wuf���ʣ����j�_<C,�ϼj:m*��^G����q�f�o�b��##�,D��A��Ч'�SLܢ�>q��(ؠ*B�w�W��T�V-r6�_:�`��QPBh2�_!��l��.�kk'2K��M{�)�p��dd7U덻G"�]˃{�З���6�es��]9�#6-l�۷��C���ؼl�I63�=&�7&� ~����>>�%�<A�]�tj}9�O%��2_��7��:�PY._��a��	���LR&x����Yx�b�\���&>��Qh�LΫ��!�h:p��l[|F�Fk��4E�D׸S�#j
�XB�o��ͭ�a�od�ꞆE�.:"��mQr�&|]��NA���EE,O�5v��3�W@�Z�܆��Z1ңOC�E��*�PP����fb��b�\���U���<��ܵ��Z�Ŕ%�Q1Dmz�O1=R�G�`�2&���Ir���*UD<=���Hn�K4}�⮍��X�3C��A(C���RT$�;�X����{tљ&2�FŊ�;-(�Dk`��2�g(���ɝ�F/Y��R�`�H`���8��M<�.!�X7{Oe>��F�<�e�\�� 9q��s5��m0��]	6�3��2AV{;"�h���]�PK�Wv�_��v�+{/��P�46�R��&s��+�-Y��3�	�m;�E�U���b>�*�y���E(�v$t�ɬkt���e��:��.��VkLzl������9�oj4���x��XY:D�}{{t�v��j;���pT��Mvw;9�Z��!Հ��]�P�g�h�$�n�9{a�um�L���&Ź͗�(ۓ^�9T�P&�s��oA�wUf�E���Px*�q��r��M��=o}!;�P�J�0Y\\�W0�e�I��[��n^�5��AR���ʗ2ꬬ�����N#U���oyb�z/v�ĺh��,=ݲ��(�������ǅ�}Ҵ����}SG��؄a7�wQ�bR�����f���p7Rj�B�����q�W���޳���e� 
�T�.jyqR�V�ӽ��m]Т�#{�T:����U�����i:CV��-l"�C��a� �{ա�Q��g����U
fet�V�6u���.�[ޭ,ř�];;ض;��H��:̻.L�Aǳ�Y�K����S�Av��ӧ��/S�ֱv@���
'��Eϯ��Z�7�xm�*����0S����Zv���y	��
qo[��i�mA��ھ;��>���SE�}���ky�7R���[\&ۭ���1��^�ʜ.�V1)��:\}�dQp�0�ו�^.�I���.��0i�����}�G��⮂�I�i�[��9���3��D�뻦�2oS�V�I	5M�p�ƔL�p�
��bYt1Mb�����짗L��F��
7�ǶM�g� ��M�����l�6�d��U����1\)�[���e���8�Wպ�r�;�뛼Q�u���/%�/3�����@y]x�>�c��gww7�P���R� ڧuݲ��!�l�ST'��3]��n�K�;�,�-��r�;�G����T0��7��Њ�V;�c��fֳ��S�x���WO��nە:#�R�k;;oj
�{7$��|ө�\1 �
�<N�Ӳ��.V�Ρ�0˫��8k���73��a�V�7{��j��VX����9�f*�e�حv�U'ۘ��9@�ݫ�{f�F���x����m�͵j��r�FY����czK갆L�6�:MW{(�ZԦqT����^���eݫB���CƎ�;�䬥®��{O.el�1�9��֬�H�У��d����Q#,B��;HW�:��n�k��?G�{,���,��%�A��sy�&91t�[�h���V ����k�C��:��v�7K8u:���s�lC�6��ǐ�AM�qɒ��[W�I��\�����h�&�
b9�-���U���h���O{��������Ƕ6�,�y]�����J"98�#�r��m6���������ȓ-�o^O[ll��NY�y��G�Z�י��%�{ol\�����p��9�=�K���佛^�8;3�f�`�V���D��H+ۻ9�H@8��M�9���l�m���I�Cɳ�Vpv#�nm�'8㶳mbZNqΙk4�dR6�H�ť��+N��";j�fd�H3E9mn�lq$t�e�ά�kdq�۰�Y�mY�İ\)0�p��Y`���V]�XZ౎���H�"�:�8��3N9�,�YQq�vY�v؛b��5����3e�cC���.knYŝ�ͰI��]��6:N̴�2q �?Q E
����t-�ұNt���_C����|d��ՃE}2��8��$����!����ю�S����uܠ��r�7Q�\�����O�t+��c��{*�7N.�X��>�N�
�!+ �\�R�A���Qw#nn��)R�a]�5�9_�p[�q	��WG�aA���x}X6RCǇɍ?�PN���;r�]�X�J{U_K��n���B�[s�L�"lBr$!*$R�޻��[�z���1 �����ύC����(�#���p5O9�d+�}e�K�'u�%U��Ǔ�I�oz}�:D���(���;J*.�]���!W��
�:

[Z㼖b+^�-�F�+�z������	�H�X�b��ZPXt=��s�.�_����B}]���Ѫ�����"3����>�z!ѹ�X�;^4���
D�}�t͊��ە�/�8�U8�5�����Rn�r�h0��l�g�R}ή����k�S�7cOqKh�I��k����+��/	];C#���d�F/���� uz0J��1|i��&<S���Bb�a�U���b��U�/�ňp�w!�9�����7����*���Cy U��]�uewĥ���@����{�.���^Y9]?	䞫,�7��K��\��}����Y;|�N�rD��k)�����#1�g>*�}�Ap*v�
��J�5�)��9^U���'u֡}؍Lv��{�u�9Fˉ��ۣ��0����l�=�5����x(ٟ(��m�����9:MEE�5�.�b�/�;�R��0��g��e{�T�R*������:�p���v��Sz��e�f1�X�iT��轖:��(��|o��J+����*^���!n���R�o���V�}�-ˮp�1V55p_���8��,�V��L�FҨ����HBq4�l�y�;7q�g����/�!@6���85V91J�eOشN7�����A]������օf�p�;I�v+2���a?H���]z�r2��JNODt?s��Qc������ݳ@�S2]��h^G�E^�|�Қ�a�����i}���ף��_����CTߓ���wY\�l>Y�<]�$w8����G�/N)51���QA�Q���^��r���c�rjYJ�r���X���L[��|��- �	�+`T�l�H�4.TLP;�����C=f��?�>};pF�u�\<�ƙ�..e0��\�ԟp�C){Ţ��H�={�������v�\b�'SޗӨ�,���Z��|��K
�,$��t�����%]#)�u^B4-��r�+6b��s8ER�K������].�jc�6�.�|hn��o9X�?$A;���kf�.��[�Ȃ�&���n�q�i�f�^	�!�l��U��{��Gw76�̭C|���9�p*�&�|�!��$T\5צ���lp��nݕ~��ӓx)sO����^�6�8��ۜ�>!����1�[�1�C���ۆ>�e�E�Y{=)+�!|�b�ðn��e3���oP�|���}"�z��os�{tN��t�$��RK�.g�2/�H�*�9�f�㻨�E�6�]+���=��1��}d=�!R�K���ᩅ2v�j�ǎ+^���L��tK�AO@�;E���L�c�u��#Q�*�0ʽ�O��-�s�������A*���z����x�ѝ�{V�r�[�p�Bv������.,K��87�j;شN��4���̃$<���Ȟұ-\g����
6�E�ު�.�NV�@�;�*1�K��[a��Ñr���Ky6ŕָuJ�~4���$N�QPo�[3�s�r�ʅ=v�ƶw�O��ހ%&���O4�����؟CQ�T���0Ȫ
=@�;��[*
�ϥXnA��	�z.�2x�բ��v4�׆��j͝M�;Ech�[.��g�����t��1Ч�� ���9�9�	�~��|�_��hu
�]Y���A�u�)��*5�K�8��GK�v>�����l^�{��S���K��X�|�ԏ-oS���j���D��;��Sϥ����v&���i��p(��&X���t�eE�t�(᪃S[x�B���{yU�Y��_*�Qї%�ӱ��nr4Z�����}��@��t�,-_:�|L㽮}ȥ]Ȫ��TwK�(��]��I��&,d�����)��nQ��ǎ���1�q1�r���y��\��:�`VOj�q}�;�2�X�f�N{�����X��R&{���w+@߳^�kr�ׯ�E���oC��{]I����券0D��sn�v����]�b�����B�pT�u��An���r���_#nE��L0|�QQ�j6��_Q;7�%r�Dgz��M�תkL)��#���aI�ī>���'�|���x��X�����:{U����v^���J�fP�>���rV(d8��}՞�y�M��y�Ve�<�y$va�I�`�j����Ya�j����*ǔ��L�
.[�AN^�wq��p�2�"�R��Bp�A�v��-���o����k��f�V%[��xҢj�L���ӈSu���������c�j��t�z��
w�߰��V)�
{�1^*���rNu�I���M�-�,���\��Au���3����r�[�7�� 7[�,���+c���PF���㙂B��e��C�yz��V��'r]J�ez���H�T�q��=�0�%6�+>-�NG	y�606��B.���E�J��ow�Td�!�]�LL�P8_PP���.�=f)ʽ`�I������ߴo�^��{[�-v}�A	�/�Ə�GQ����7ʈzk�{|v����]#+)�&�;��w`��w��tjv�B����}R�8"�1R"oy�E	��V�ʊV�t��r��(�p�)�&)B��c�{�n\��6;ѱ�T�%T)�RR��R�e���t���+��=ܴ���"��|z,��&ve\�뚃i�6� ��GU��wn��hll�]Ml�L���T�����\�����t�����8D؄�HT���Bnr���/J�ǩe�+��Un\Vp���p�L�5�ʹ����P�qn��E^�i`�7^��6D��
�F�B�$'J��/�ی
buc]L'3T��ѧ�r�$��or�,���Ct������w�$n����R�.�~5�䠰Ǽ~Nc�eUx�w�����*�T����a�F���w�%z�V꿯��]��Z�.�O�3X��U���\�]p�`����%D�Z[9d���\]oB��󩕢�I�T�p�۩��O���m�˭��!)W60.
���֠[p�K�6W�VL���]ܫ�XU�Gqno7ܩMt��Ep��5'^��<�*}����������*x�6)������k���}��A�W�;�	��t�b�Y��3�<��H%�>+|Ws|.R>M�Ts5������Sjn:༻Nz6:�Ga�͕�nA�1���uz&Ⱥq
Mmc�o'�\�1�\[[}U������;;��ӎAv��<Ce^l���q5
)<5�X����LVu~Ϧ\e*�qg���
��V�F{j���Q�/ |\[���p�@�O+�+��Mvn�PS��J�
�~�\ yE�t�!܂�n�-�.�6�)TJ�7��i@��Ւ���m��ָ*������̐eѮ��wJ�
nz���P�^n0��w%me�ov����r�j^u[T�I�[�@Z��y�el�1Ѵ��3�5½��C�o5�(3؍�W��]��#5P��
������X�_��P�YS ���R��Ե�$�/���W�����C�䬁T��U)��w�m�͛r�Yu{(�vs��Q`c�-�;�a�6p�Cz.=�Q�FS9��*&�|��J�"���r@�vqˀ�FIZ�GI�h�{�;lwUÆ���_��jC��i��N���2N������yIm�s�q��7֕Mk�'��)u�s��g.�-����]�ݒ����m���&ʺw9D�K�{�tݾ=��ߨRд���Е*���PH��У9c��nBSv~�e>���<;ٳY{p���yO>��?=��61"$Dyz1M��5ҰD	��Q�#_R�Q<穅38��[�,��{�v/v��pH���N�Em��D�*+�`�H�}��i�.�˖��Il�+�{�.u��g{�2��P�҇�P
��E�e/x�_�u��^SQ�����r�z�9�����s�E�
���]AN��y*.��^�Jɂ��-��V�yd(~����9�s+�o�P�]�89�\�p+�Z�<5nl*�Mޣ[ȯz��r+��lR�,�j���0f]���z|��(C���0�=�O%@��}}t�ͷ���t���65^Q�X%�5# �'!���c8�\r	���*\l��z�^�R��t.��*,5n��}�/f��L��ו[������	�|E�>�/T9���ܓۚ�ʽ�(�R�|nY�t�F��_B���IS�=2Dz�
�}�Q��H�!�����4���y	K/�i9��^�S���\wB��_]��Kv!ZD睙�m��<���O��2͋٧oWP��in�&	'ZĩH�oQƍ�(��,�=���q��kYdU��{=��c�����iJ	+��۝�،���҂ݶ���#�k���!�� �X�9���<ka�����Š��k� �����Ȅ�:g^�=�"�me4p�SS�gڪܸ�)ʽ`�V��
��%�ئ�����}�wbPw/�N�_�$��'\���(�=α�����N*��R�z'j�|��\�JӰVEz'�4OA,)��2*��Q�wQ,v��W��r l]G�e�bX�ퟶz<�>�0|�;�y�P��*e�J�Vå �/�7�7yzl�74�s�JJy����]������OA��(�!*)zuI��*&�e��f0�N�:���c���_N����t59΂��㡚yy�3z$����^B�a�7�6ő���n�]]lb��������9Op>7�>l�t��<��;�
2��9��D��J����\.c�`��9��DU�7�oC!ōu&Wg����b2�w�"43��m��v��]�Μ�GMm,X�#^�Ѩ/8��yذ^r6�X�STGK#�؎��ŉ��e:n�R;fE��9)�W�TG���72H��G��fty��L���fg-�i����*�H�m����]�\;�عx�8Ľ��&�x��od3m�K"G[��m�*p�����Gu<7�wj�V�v[]�V.Tb��h3~	U잟L�r	�,X��X��y��ϭX��e��<5�F�N7Ǡ�٨!���^��-�u	YG�R���F�>��x]9�}x�/vB�=����Vn���-	���9=�ny2:}Ad��l�7�s9N����m�Jv��1��p�PS�d�)WE̡�Pb�pg�#[�6:3]�����le;������8�m�z���>5��4�4�;�V�+g��d' �y�64p]�Y�cx<qI��W����x{����k����b�(����6��D�S�cX"��*�����O��m����N���E�X���	��L��؞�A
���{hY���Т����w��<9�F�:�K�q�DAS���&��bv�V"F�����!��b/��D�k�Yfz��{g2�#��Wj���U�ϟJbP��$m�lK=���B���֗P�ܫ�#��{vl��il!�,WW��v��r*)�lq(�ZgfU�q�5֑��8R�R����ff\�t��^DSyW'����׭"�ڮ�ǝ�u���D����!R���s�&d� ��Jj\l-Y٥x=Myѳ���/|�^cW�wn��Yp���Б�x��Nͳ��R⯬[�̌ɚ:���	�#�{��X:�Ήm$�Kw��Vk��3�{
\ĿUF�C�E��qȨ�����P.���ܟZd�;���e%���P�S�v��Y��K>���yJ.�K�r/ڣ���<�r��g�l�9<D�q�[���-W�C�X"Hl�*�"hp ѡ��@rt��&?Z�w����1����+����7w�LfJ�
xQ��:�|9�jP�E�e+�B�J����+}4�K*�s\�F�땙�6�/%�LI�PS�d;�:75ci��<���2����]a���I��\����f�p0Q�v�6'=ψbç���7��jyɩ��\�c�_SwEj�GV�U캞�Nz�a��nz6:��^C[+f܃�F,c�*(]3A�]��kp���7PK�v|=��GZ��,���p7S��sJ㳸���rd�yG�����M:��ކ%>�|�l���)�����}t�z#�v�SÅ�b_p���|�$�#q���[�	v#��\t����³~_`�^66�����^��W������>�b����-�{wW`5����Bv'��7x,R�8�,<�a�cw鐀�Kփ����a�5���E�{6��&��r�<�]�w8+�4�뜞U���䚲~j����M�`�B�Ѵ�WKX�l��3Ek��1Bd����i��x�u4r�)ű�Q�X٫}���=�e`F���d�2�$�ֆ虆]|jnB#������_���m��ǲE}�mWrЯ0���r}��s����j4k����Է珜ڄa��
y՚RUuq������+�\��a�D�@o'g�/���G�GȌ��<
t�]������Ia�k'
	�ۼڈ[y��֮1Dk��ר㒞f��v^�'Z��Z�2�Ϥ�j�+]X]n��E�{	&R\ɬZ��N���2 �n��v��眝p��w{}�C�lw��째`�j��@e;�/��m��u2�V:���:}Ԗ�D���W�=�':�����ջ�p��� *K���6�f�cG3��7�}�m��{ܬ�pq�#/0�D+G���R�vHݡ���qǗ�Q-f�xOʅ��a^�cZ[��\���� ��b���ֳJ� N��5ʙL@kx�uأˋ�v�w��U��t1��:��$t.��]D�z��9\�o"8�Yǹ&K�1w߮�i[�)��h̙!q�	��+����!�Ec��>���t� ��9q����gy�&�Sa����a3�ޓO>j�%�6�{w ���;A�3�G�wb�p�2�pD�[5(rc0���e�!�fﴺ�9.�ǲu��v�9�.���u�����)��#k�LY�ii|�����ˤi`5ݳp��lfύc:�b����|����zJ�AI�1y�p5��f�U�4^������Q%�S�����]/n�]<��?�{��"�[��/ΰ9�!ެ����[�^N�Z�q�b�Y����dθ�n� ��,�T��V�^��[�ӥm�٭�V�������
s͹��^a�s�T!���1�w�r����[ޔi�������2S=������8:�a�*���rg`��I�@��6h��R�	P�jX�r�;��5�����owl�g��ӎR(�M���$�]B��ս�tj�!���s�����V��:Ş�|��G�*���S�bg-XLYT4WX5����^���:����Op�,��V�˧�]��m��6��]�}1mfk�{�S�el?d��x�M+�7�r�6a4.�\���v�OQ�]ħ^5 �� ;ʛg��';$b��"j%|Z��C]�S�Ac�Woe�Ņ���SkF��HB���\";:rI�ǧ!5y@d�Ye���g����,���=��O'�I�]���;�n�J޼�6N�*V�����ӇmK|i�%����X9o�:�c�`�P��X�n���O�+��S:��7��k�)u�1��Wj�Ƃe݌Z�(�Xtݬ�k7�)P�\GƩ����[��f;C�`�S�ܯ���cʡJ�T�AR�f�M!�5��mm�t$�DtF�H[%�6m��rBsn��m�ܴ�Yjsj�e��2��*H�:�K�)mv��Ig��N�3H!�Vu�ͫ�4�������M���-���Љ�Be�nNm�[2n���`NҶ�����鑸���+f�68k6��n�۶i��9��@Q6��ved�Y�+JͶ�E��m��k6�� �bj$����&۹83krZ6��fZ������e�q�Ls��u�fݶf�i;-���-��N;n��1�i�6��9��R�3,�3M�J�:NlI�|(�
Z�N�JfƘ�ʾJ�^cz���c��:{>��)���f��;�V=Kj��]�3+�I��B*�LF*��ɍ�k\�9�qi��ǝ���N4�</��9�zg���(T����R��=`E��==�&�^�7nQ�T�{f�K�:��ꚸ
/X�"1��R�d��#F.S�p[K��®�O�e�6��V���]w{T*�VЗ�
��<gTې�1J�S!����鞩x��)��*��B�iA��OBu@(DH�5J�I���ʀ���E2.u�*/2���bO3���~T�;��L���=(Rชá�>Ω/���У �ڝ�	M��񫍼"l�z'��uҬ�q�����z� +��3`bdHD���$��h
4�p������`vwo��Ύ��Ti����x�nB�@�����h�� �J�.f6qUsM�p˅Q25c�v��0�a������
�s��o��$����ʨ��I�*&�Sr�U�u��������h_s�32L	������߷��s����rj7��/"EE�>�^���щ�J�zZ�vi����>y�	�*�4�
�o]�89�C�^V��<��Y�~��z�5�@��G8aҶ���ŵP�@(��!�l	�w/+Lǌ�@��OVq̀)V��B�Z2./,������K\�J�)��Ú(�t	�����	z���*�\�q�w�1��mc�� 7��g]����`�C�3l�;;�Զ�B���<)i|��/dnb##}�n�wik��b3����62��]�Uu��=!���኎�=@�
��	nH# ��23��օ�J�ŝ����˜>or\�a�Ⱦ��MV�zw�"�j�A�[^Uc��R��:鿐w�;�v��m��\r�,N���s7�g��*�/�򾅣�Β�=��$G��PP����ۇ�Y]�VA�.�鬐�M(�!�n�� �I��	�\\����WT���`�k��3>~���U��7��W	��GJ�(�g��UN�.\�)ʱ�jӰ�K��Q�M	}��6���_���'cc=C�8W�@=buʊ�e�=α����y�.ʮV�޻,Ho�s�G��`4=�w�����[� Ԡ��0Ȫ
=Gy�E������E�qu>ع�Ϡ;�jp����zm��;�x"�
^���%��t�YQpU�'&�!);{3m�yR�aY����SW.:9I.�;�O��=$Z�#P��n�<&z����:�-U��`2��B��67.\����`��݄��d\ (;�f�N��uܕ����襅���"�&�C�9��K��<D�E]ל3�M�ٍ�S�|�ؐ��,�����\�����w�]9`v'{Z�`4Y���]�!�8ݕ2}g�s��l�)蝺����Et5<�(4�8�f�^Gbf�I��p!*&�3����r�Mni��~{�h�����g̎*b�����y��;65E8�����p�K�uX*HHab�"���n.^�ܓ�����]
�/��WVB�P毙}k�#��oC!��2��w����{��ow��J+�C#Jt*�p.
(T���Ʈ0�qP}yذ^F܈���=l����F�jɌ"���@�N�d�W�kL9��\=��XRs��~����o����N��VeAm��+g�f�׮d�.��ins�J�?%R��H�K��Y�Y�b`n��a���;�JB{z�Òf��2:}Ad��3�&���:�S�V�/bR��mI=˾j��e\�S�O��WE�S��5Pb�Ӏ]�}������r2��d�e�ǡ����h����D��la��[EȺ��l�q��%+�T\����!9	P5{{�W�]`2��@e;�d��{��fQ���~�J�(��]�{阧+)RĮ�A��^�K���W?U��:�,9��|LOn���rH1p������A�f�}zA4�Uo�s�9�bk9���������$]�<R��g�u�ki��5�E��'lgQ�WV�93�؝�y�mt�Q��d�����IVWZ0��x�:�N*�vs�C�?O�z�ʦ��Nz��D�3˰��N1jU9���ʏ�`�R� �8��ٸ!�l�`D���]�(C�R�Jq�v2�.�b8ل����Օ1ae>�LR�L�p�eU���ԋ���ލ����Z�+c@�;j)��fqp�K� �U�;ǔ��X�TS��En��3�*q������׍p~�E�����Xo��Z���@�ȻȨ�����e�B�gr}<�l2��6[�/xV{��4|/ƍ/�K��@W��<y�CJ�Z�%�\��曧�xTi��d;Gί���vb�²_����U�$�Ϡ)�"o�0� Q���@s�t��>��n.�������r[�MD罜ћ�������H����d��D��H�.B�Uq���_\;nqA�ׯw1J�in����{7��VK�B"���5'^�a�X|;[^T�u,9��i	���DrA����C:ސ`�7^���f��Gv�6'��a:q1O,�~�}�<�Ԟ�[����CR�w:��kh(],l�z����vՠ��*�u��ݓ$$Bg��f,��r�۴p�=��2������n������ZӔ�ǒG�J� ����l�K��8K����+
>Ω6�����D�Q�;vݾ�����v��L���i��u��~�ݛ�~��&���yv��h��!�v ����6�wW;��{j� ���}H/}k�k)x[�4�:X�r�p7S��7�q��X�bq�/&��Ҫ�1�����;��}�)�W�,Vi�b��Ҡ��k�����<8]b_p�<�n`�79QEv1���m5�+g��܊N�z^u�����l	�� �Ԋ����	�#r���	G-��{����y�e��竀��Kt�\0����R��v��J�����<�G����9�[W��#j���gU�MD�
���#Z��y�Y#F.S�'�O,������b�|��!Fb*��&�}}EO�6�k��k*d��-L���A����t�E;��K��qĸ���f�dS��D��nB6�@���Q��(�g�`�S�=;�9j���~��T��@ī)B�=B\3�
+cx�(���=jd�q[�,3��w�웊���n�����&D�Dyz1L�k���@vx|7�3�>k&���T��W�S���u��,[�K�����{F�RyV]��l6�?z�ij������r�/o���O&���g�!��-<Nt��)����7G^k�,
T�n���N�z�q
��XY�]]LW\�7Ժ�S��]���d����~���I�h�
�>�L��"�q"AК�X)0�xŇ�H����&�m���QS��n&(E}8!@PwQ�fw�e�إ� ���T���E�g�xVq9ڂ�a�U��辙����1�G�|/��&���s��T=��]A	�/"EEǻ7.oYN�U�ܻ�}/�)A>B�M*�:g6s'Ӏ۰��m�=������AZD�����[�ז%@�t�J�YX��5��f+��w�{�a	� �ݵ��Ԣ;�y�/��ܭu
�_p�t=�h�AVNC9���|� ��RS���wo�� �� 3�r-N�P�g6xt�����V�ˊ�k�w�Ku���n>�¸T>�Bz/*�SܨÀ�W��9��ίd����4�Z̻���Ǘ�����w�L8S�7�,�zC��d��`M��`2���vN��ɂ*��ڵ�+�C�=��wP�zZ�~a�c��9LA�8�W�J��."����a;���7ZJ�5Ì^_=]�^�B*E��R �\1'�mp#E��B^��;��lEI�ĶV�����^_*y�o�N�����w1T�>B���v�-�b���*��q� �s�Nk5�XM)�a�����ENkE�@gf�s^ np�YD����Nd�Bإx�;��n���b�+�4S�1�TTp��s��c���,��14o9g*�[�P��&Bm�na�X~оP�:�Om%\>O7������Q��tm*C39~n���ӎQ����Fǻ�>�0Ct�i�p4/O@�P��5�Z�8�z+��d�N$e����]���G)([=i��y��9 �T�D����9.�]f���T�6И�0�R+fS�v�;��t]X�^����2\ �q�+�Q�B� ��ˉc(�U
S�aM������S �����w�}.�p�	�{wH�j�fl�C��Q_�U��DO��hq�H��S���(�sl]z�R�x��:�WN"��V��\�V�[��!��C�����/o��;�=��4殽�H��E]t��1��ʊ��L�N�d�W�hi� ����ހO�:ç7Ǳ��S�Qۏwtdq���G��= 6�C��ؼ�o��D\�h�U�nj �J�8l��ua���ݧ�|���|q�i�0�~�O2M�f�8�����d�2��罗�����/�1F���ǽ3ǣ��]d��\H��mG�XW �GqwJ�m;ʲ3eXWD��W�v٢�#IbCx��e���[h��6�j�
���vQ䁘��d(�w���������9>��p���Ϫ�4����?L i�!Os��`n�Ӗ�϶�i{��*&q���X[�}i!/ڨ1�8�wٰ�P�ؾ�qxg)�M$�>�5����v��3�rXʕ��^Tp�"����$u�+~=νL5���*��ȡm�Ļ��Ԉ8��a�TR�4�&���ӂ+h�2�@�/�(Qch�p�*{7����IY��b+��a��:�0��_�~S]ձ0�FתD�'��B�-��.�TY��wxK�AY:�R�tչY."
��������`C��
�F����R�8Ӂ�$��;��g��3���"m5u1ae>��b�+��q�eU���ԋ��b̪��s�q�����vu�񸹜���)ע�w��������G-߸�veX�j4��#��7���sٔ<�KϮ��|,4vH�Ȼ�E@�'��n���BA
�]���T �sy�V5�;��>'���H��(�UW�{\�j:e���|k8jc��7p�Qu{av8�S"�Yۍ=��}ss��M�]��*7f������[�ɣڂ�St����F�:�z��������N:.�Z�'G��M��y��v��wC��7M]���������a���g pk.�^N�v��Q%�M�>��rתM����;h�)O�P�ӊ�p�7��-H�Y
��>�qlD�^����ᔣ(��V$ �QPe�b�"���|�{�ʻWLC*�]L7��(!����DI�A�(O�}��I���L��cF��s������f���W���P��%�U	Ϯ�F�i�� py[]�egyp`s�/�ܷ�};讼!:p9���Ftڑ�5�״n�LW����?Oo��Wp��-.�ܜ�{�P�������>�诊'��\�!����+e��������ͧ���Ta��*(��O�R�#*�"���a��E��7�q����:}QɈ*�'VBG��%
Wj��W{>L�͐��V�����&ϙ�|�Ү)����͍Ď���"�ׇ/���z`�龳��AN�^u�����l	�Y"��	��U��p�� ����Q2�ӷ�K���5�k�����s��#u802��үt�ed����J�J3m-=��2���W�ב��S`gU�OT��QcX�"1��R�d�3J�J����uK�ɚG'��R��F��ީ�.�����O=2�j�;r%����{��yn��� #Ū��,�����̺�o�d��Gl�OV���*���T��NN���.��q�Nw�-sw�d[�/�e�껻�rv*s�aʻy'K�b�[���G �o^R[q?+�R0F�HEH�"�h��C�|)������+��dI�E�.�6�;���:ϫ�^��A]��� t	st�D�{�܌ٷ*���Q��v%鱚X̋��#���|i�� w����H߅.
��à�𮴾���Kse��������zM\�RQp���=�r9M������d��3iА��#ҽ8��ƺVDg.w��d�w�K��c����N5��I�o�B�E>�u�3�(�.$AAД'`]��:��ɮ)�G^�G�!ѳZ�":h\����R��A�Fa���e��Rp�@r��I����އ�T�����W+�Cԋ��Qe>�I�5���W���xR�������w���D]�r�Xۥ�zuXb�Wkⶖ�������&���6�Pq-���5v���9��:v��n�^>P`2�a�������k/*�V�.4��&|~�n�l��s��d���Z�<#�ӱ��l��q�U���𷪙�_p����Z5a�V=UC�<Lx���{�$��n����99<������8�8��j�/+�q�
D���v�&��Z�y�Cݤ�
��n#P�7��>Ty�n�/IΛ2�˟oǃm	ܻ���j�o��W�z�|��U�jɹkhBv ���h�ouF�5lN`<�����Jx��{��5M������˴)p�K��-�tw*��ë*޻�q膅�v��X&�s��u '+6�t��$YK��!D��[r�繰�5�˜<|p�[d{.��.��)>�Q��T���b�NY	_#��ձ��q d8�t1>��4� �%j�Jz���օ�p�f�4ﷳ ��R��H��4����p�|�W�7��f�YKn�}�PsZ_br�i���\��:��6q�-�������T{gv��}�:�P_`������,+��Ov��,lub��2�u�"��8���]�gk�[5##N�so�X�.۸˭O�*�<-w0:����N�j}��.jVDm��LY��l�뜩������w�����kV��U�<:�Ʀ�Ƴ��yTf���i��]=���f��v�9âr�D��	Hd���U�ih�5�B����]��|0]�ہ>B��r\�W�;��ի�퇧.����:�t��h`�V�V�a
vr����y��/�wF�u�U�.�tu?�1o�d{��P���ϱ[
�N��,��EV�BR�̌��D�����t�>A���H><ir�PIε2���Vhtpy�\>+=ڞ]f�]�u��Fc���bⷘ賉�wkr��4�gd��.a%3�7��XmԥX+68�Ɠy�ȩ�Z�u�'�+��7���a��Z��<��Oi�ϭu��c&����eeՆ����h�k�Ԧ� 7Nˬ���x\,� �-��>��m��Y���˥���NAx�9�-wr݊�E����O�	g9!�b�|M�=}y���� �\�i�]�ʪWZ�cP\�Θ��w��7]�٣X9�2
��MRoL�
�Wg��y�nF���f���E���W�M��v�I�p]�����.��%�
�l[e'+��7
�-l�#�.wau9�(T�ڶpճ$�-�In��TZZB��m<��-O�.��ܠ���y	Zso ��t���<�GF���T���Ot���e��u�9��X
�و+/&nP�|�o��j�usq��]�9Xt/�v��eԙ�������C����ʱ���K�_.�D'Tg*]U�B�{q��շ9wZ����N[E%��֐�e�W	Rnb2�]���1�}��3zbl��R>�)[C�u��)V��q7fu���Y�6��Kn����Y�9��F�� ��P��Xo{*���}6@&����W��1�� \��]O;uv`���[6LX�O_I�1M=���y��7��`*"�C�u�[m��r�{׈={Iͽ]F��MB�+�����V��m�ZĪ���i����j����nѴwm��Off�kN���m4٭��[��-Dm�:-���[m�;[�ٳ5e�lٴB�[,۲Ӷi�s�-�L������Mn0�I�m�m�z^���m�fI�3��� ��n�d��Ckm��I"��7h5�ۋq����-m����ٓh�ٷ-��խ�id6�ck{j/n�q�@�#5dn6�f�ZQ�v�B�ӱbͳk6��g1�ĝ���I��m�r�&;dӬ�[ޱ�X���e�ݶI�0�Xe+90�ۚյ���8�v�۰��޼��HmY�6��kn�̷%�i�d۶֝��2[gC[3bN�mh�@P�Nu�y'ŕ�rqdb#o7�A1��{�����N�|�Om+�7��;��J.6Y��tt�ݔĊ�Vk��y��-��=���H��*�К*,5n��@��P}b���쥣�ࢥ�<_�}#�6y¾��L3-��2��=ʌ8�Y��v�uޜe��Po�w��E.�4�]���X��ޖ,P��L��=A�.�!���&��*�P��읍�ؠ�ZG��}Z^��_j7�����Yi?)�B��B��U;�Un\��X��g[�'�c{Γ<[��䮲p�F����s�].�u/�U�-��M|��:u��Ln�ޞ[��'tDc��i�na��/�W�}�'�Ԡ��jU�a�0N�듽Ew�u��~��s�G��S��8����t�i�S�AzzC��l��P�T�c�[:����˥/U��K��Ro��GZ}�OA�֩D�!	Qd]�F�:��r��Yr�c�A����{
��Q;��t]]8�r��rtpI��2��FJƹi���� z'bk�+#���)��L_7C1����ʬ��_g��E��w��lN�P�5yr.�s7:�l��ڊ|����M��X�9�,��So�ǨE|%�2�iV�U��.זz�]�]y�W�c'�rj^�/;%�}R!\�+V1Ӈ&�3����@Q�V��p������w��g��ч暃���o�(��Ϡ�ΫI��1Q�b��G�B�P��=4���/�^�%�A�QmG�dk���yL��0��W��# _���t*��>���5�=>j�/�3���]w"rj�<��r��`6mH�s���@�N�d��g�r	((��q�quB��3b�o�g��8�d#=��%�L� ۪��y{{���[����?/BmE���G�}�Wr�^��~�PX����Ǫ��u�fa5ϩYю��c��;tVcYH#˺�����VUo�d���0��[�͘�z�������<�j�W��^�ȑ��{*���U�>����Mm����c��%=�a����dC����R�f��=NR�m�%�(�j�z�b�s;uG��1[k��X)4���.~��*���^�A�3vt8/ڞ�nQ�T��v�"�m�KW�}����}/��S�)�V[�f�[}�� �-�)D���詙�8,닅Lep��'9��Z/���D��;�d�'����s7����@.�7���m5י���Q���-F���oSڛ�4�N,j����L��F��=]���Kk,�PCq;�V�WeX�I��d��;�d�}Ԧ���*�XL$F����f[�"�O�ҭp��G}���U:�(�r�b���}ʬ����Y��.˽g�&�aBs
m�/wL�S���ҙ�[&7�_�_>�ҺUt6�ͬ/�z����~s��Mna��ǽu��P�R5�(t�Dƾ}Zn���srej����TWZ���ŢD��������U��t�X��E�#w�\�K���n��P����j���C��lpQ#�1A�T�B���F�X�5���Қ7���/\J�)�l93�]N�_A�\Tj�4�Un��|7,v15iI�U��ot�,s�ni��<z��D�\������t��Gյ�ھTn�O�����w �f w��9 k��s��d��h�X~�{U��(`n�9�]eP-��j�j�#:L���3UR0p_q4ZYRf�����e�ˤ����=N���n^�Cv�ЂĘ%6|�g1�.�s�S�mK	�z�h�P�/B��:��������h���y?�z$�G#��}?�Ϯ�Rz
�]���E�"������ڔ�����9���>g��Vnk��7�<`�s����u�L�;��ٝkzy��r�a�5��=e�e3�9٭���ؚ+�,�K9c1��V�f�[�����:ͺkb[kf����N�_�\�H!�c�7^A�a�V�N��:��Ju�bA�D_R��Sx:KW���R�2�>}���:�����],�,C��'��B�J(jM�]W�ھa+f�8�F��ܾ��+章���[���6;��(.5N�)Ex��ح�f+����C+8k=�s��L>�|9�,|gm#+�{;�!�@�����O/�/7O*Ԍ+�c]��i]X/R{k��N	/b�#Z[y��Do{7M�Om�_u��˽�9�i��ľ���M�
A���.Ma�
rׅ�K��#;':h�c�#��g�4a�}�J{���̝F�^��wDEQ�H'~=�hn�bT�ꛛ'��4����zi8���g݊]s���_�V&�W�0Bue��&�|��c3(*��K��Hk����W��:�m��Af��K�6x��3�M�h7�b���7
�����']3/+����F䗙:L��n��ȸR[�����<}|��u'Mee�Sٷ���a��Y������8:��	����ԛe�-���:�drv+�N7�R��jhvh�#��>�f��T8b���U���[���Dn�{�'ue+(��"9�,����v��P��NaU1�mGb�䙇��}�-R{��2;0�Mw�t��LI�Fmz��/-��,�Ɩ������سZ�*���ג���v��l�OVo{]�vIdf;�T����b_k�P�˦+c%��W��CdJ曷l���p���Y�Mȼ���<���{��^lO�nW�7�>GeJ�o:i��f�i����T���
��S�k}���$P܀�����^:��MZq`�:2�d%8�F���p��0��sݏ��E�����Ď:�(.>�v�r|^�����Γ��-��O=ýJ�����gWDf�j��}���
%9ٿ���r�G6��7�4'���8O�v��S:�_T�屷�;m�8D�����V�SL�Q��A�DM��}Ӟ
]X;��}(�S�t�*�*�T�Vf�n)?;j����4�����Kl˱W���ٶ��������.	��%i1���[U~�*�_q	�'�u���I�f;#���9fe��C�79���#WU���v.���i]Y|ϥ��2TNG1�&�(%��}w����x�S$!��#�]�m�Ϯb]~��Ih�]�A�W�#*f.So�Յ�D��hpQ����Rk���N�"r���w���˂���+�Ӊ�h[�x"�5��઼4b�4�]^V��*6�ܶVo����
�Kw��[|uRhs�+��5��eg(멭�bYo[�Q���l�vv{���[����r��:ʮ�2n^��nx��y�mj��I��-�X�	��7ި���=�U���+�ީՙgA���&o�$mU1f'�7+�)T�*rj[�%ژh<e��kۮ�����**(i�]��=�L���&�:��Š�����s�AP�ײ�\�A�畜� S��]gw����!h敖�S��.v��R�8�wm�b��p|�Ղ��J�t\��uwa5�wz]���ʽ�TV�mՁ�t�T��8��'q���Nfk4S�v�'��5ڳ<U��y*(���+��K�0�wZ�i�-VL=��\�m���I�{x�iJ�f��yC�:����]���)�a�n|�;�l�ObZZ�GɦD<�J;gV¡�^���w���q�v��0���"�%'��7�%�b�c��V�C�`F�",8k\�V�u�}o�.tvB|yE�$_Z�_w�a"5��|gݾ����)^�T���χ{]J	L��Q@�V1[UO�R �㝜^���)���z㳖��v�ɴ̂����􆑪���Lor������׫ғbHK�VkY;�r�s�����P"ӁAb�$kF�O�#��[� ����\���FU�~����kh�}l2#N/�*��P&��6�Ը��y��ˡꌍ�ޓ��ƛ�]i�r�wP�S\W�����W���h��cbw`����o��;W�t��I��M�fM՛��dL@���Q��5{��/�'G*7�Y�"ղ!��T}\�di�\Y���[�=ْИ�u��;���E�����U�X�\F	�ŔW�-�=ޮ�*�(VRyͩ���>�+(��,���\�-����b\�؎���������^Oy��=��2�����;��\��r�UZ���Qr������v�l�huC�:�¤��YyM�w �1��x�Y��a��2����[�-=�ʭbp,��NaV+*�o-U���؟�7t�X-��l�{����X��g�����5��y��`�@N2�w.������g.@�+�Q|iu��_���Yw��e�vkg'xfĊ}Z7N.�D�a���)���CY)�J�i��f��nݲ��<�J;gs޶^λy��w�F�oBr�H���B}Z�>אmS��i��_V�ryV(%�����J�i������8nC�RR��N����E���mѻ����KV�Ǌ��cWB!�Z�9{,l`�oT���:��<�y.a�:n��ۆ�+;�YGrT�ۭ�k�yM�i���^;��L^��)�s�)�U�K�#IĞX��/8�L ��4sj����zD����^q�m�Ʋ���'=�)�^��	�H\�#v�Ы�c�څZ���0�W��S%%���ڭuXM#�a��m*�䗷�4��\��R������x���x���8�OYkP-+�/R{k��i�AX^ő�<H�yݽ{��q�a/�4�[�����Z$K��<^)Ǐ
Qq�*�p���v.m����u����z�h�@��&��������v�C�SAT�N��E�xelg��珧�y%�!�j©CQ�u����%�C�d�����+��JZ���|4k��ޝ\p�ꮸ֊���x&�h�<�Q�f���ኧ1�8�¨]�8�6�;��n�^1�Z;�5�>ii���o�ڣ�1�e�m�V����$t�iy[�'�g�b���|P}���}مZk��s]�Qa��ڐzn�ڴÈ�$O9�zrp�c�%�ᨷ`=e�Y�'��늞��FP{�y�X���z�i�����hy�
�~�i�N���1�����q��r�!�۲�;�$�$eY����v2�=���rMA�)W��v�\*�xp�I&�zr��۽7p�w_Viхw	2wG�^��o�'��3]�����-RW�7s2Jy��ެy� P�	�nym�5c���f������R��B���u�*/�d����:�m)W�؟
���!e�"�p]�������5n��1��'}�MX��؇�[atH��R|@�
��V�;�3U�cr��N+yL���X�m_0x��⚷b�v#c���J��ݥ�tu���}��[�qE5?"�S?m4�>�8�\��2��Fm���-{Nb.�nu������eܦF�.���_r��'��>9V�ow�b��7}�����V��#_,Q�_��ue��ː�R��Yzm��{��ろ�����CH�ȡ�\n�cTq�];+���&��a���ǻ�[m�jÿ9�5ʦ��D�CT&���랜���H����8�'\������8�зp�Ek��pUZ1W��)�]f"���-CQxVF�Wg�8|�9�~7�i��.롟9eh���T�[���
 ��1�ZM�ZT�T���w��2<�!%�\N���}�-u7�sh��]D�(�P.SZ�.��.]%�����qu�o�9,�N���MyVV\��c���,/�wY��Z�`�fQ�ۙ����!��H��=n%o069l��oI�`���,��\�*��񮇤�J�v7��(Ğ�\m��U�g0���k��LZ�^��N[X�nr1X�J���@w8���u!���ce���o�̱�H$Θ���Qˮ]hN�ղ�Ö́�5�\�z�]����^2;�LTv+�H�0+�)��ϩ@�
!X�L��s$�]�c����A��qD��1�\4y����o��0&2X��f�SjY��|��l<r�-֫M[\�Y��,�[��-l��V�v�P���Q�杠��μ�&�ya��F��9��!o�C���wS9>\����W�m�4oE�grhmQv���F�q���s.�ιX r�4FZM[Gf���u;�v��nط҃�D<�f�XV�O]�\J��m`u��fɺ��g�s�H��q�y]�S�'u�P7��x�i?1��Ff�>>Ը��--3PI�l�&�ӻ��Á]4FgP�ލ�����a�j���h��uuˮ1�J�ˈ*id��+f���y���gj���f�&Q7�A����j��0�T�F���Wc�i�Ck3�X�e+�q%��2�z��ü�w)����үC�F&���h�ϸ���'Of���;l�� ���"GK���ab��8��)4Ӻ:YWm�6ћ3�X�:y'&)R���^�:�+��J�KM����:�������bA.5u�������Y�;�����wv��FVKr΍�7��:�Yq�!/����,��81}s��$aQ6&�[I"{)���VT���*K�9�Ik����u�+u��cv��(�.K�8���ٷ/��v���EGof%�Y��Ƒt���7�N0�Gh܆Ћ����9�l�j먢�k��&j:ԉ�S:�P���zϋ����w�w��� 1���Z���M�s�)u7�e���X«G�R���h�ۤ!�N\�1O��w�e9���׶�9)��>��*�Iӗ�~*�^g�1����!�՛4Q�|�̨�[9}S_Z���D�u��`q�u��{T=��\�|
ͭq=��#�kʫ��4�P֒ci�}�x�W��<WW UyEf��+j�1ZTQ(�uz�e���
+����Y��2<�ۢ�ɳ�4�\�)���;η]An�B��n����3�e0U�i�|F>��˳��G�9m�˺9B%Q��]v�!õt�����D���$T��޼RR�Q��c����1L��ҳ���t���>�o�]���&�4���u�v���f�f6ֳ۬���g7��l��3{��v�ݶ�1[k,�ƶ�YXݭ�k+y�e��d��ml&��ƙ4v Scie�8E�ǖl�f���t��[�f$���sa���;L6jٱ,���ս�:D����e��ibv��M��ll���q���w�a���.��$�-��h�ܤm۝�kmgn���"q��n���e��a���S�'%��n�Z��q���dv���j,\Y��El٘�͸Faݤf�n�m�k�ͳNB34�����N�+pxk���2W�zۋN�m6٦l���e����ۦ��ͤ۶�Zf���^������w��P�X�>"� $��Z��oI�Vk^�[T��C�Q�p�իWgn�$8�Rb�����2��\� -$U���ӭv��2>9��>�.wB-g�=�wx���ښO�Q�r������4���ɈUm֕�:��^�r�+�����/�{��mKxw:ʫ'{/81p�k�I@;�ͷDzWvU���^'��5��;�g�
��DϜ���;P�=|��c�Q�1>��R�t���ƛ���'��[s{fu�9]�W4wHOV�{]�Q��`�br��Fe�+5��&#U����qJ��D�&�t�w��ͥ*�lHW
u9He߯FLq9��=<�Qki��m�K�5��i�yؔvέ�Cr>]Ü�v�Ň��A?W	)�ԧo�o:KV5�����&��>�R{GI��Ц{{!��0�N�q�$����]VU���GZ����5���X��iu��an�W����BXJe؞Pw�Z/����C[ùo���7�N�݂��ʲ����$�%,��d�������u,�e`W.�j��B��"q��k�;�q���ۑ�[�f��5�.�%c�S���G~zA���]����3R�Rv"T=�^�ԇr�_N�u;}wF�o.�7bJ=r�v�#�]rm# ��^޹"*��-�ۓ�ݽp��xL��=�.QQ�wo,��O��"^_XL���
'�b�ԎYw�f"�P�ʦ[��������G�h�}n�;A��q��7����]ofw2���7k]��׏kv9B.��.MpP.���5̐� �wg�9��&Zh>�;*ic�W�-)�om�ݎqLښ	����/]Ɗ٫�I`른���y�48:��jۿU�]�>�v��6�7Vz^����Ms��o��;�*��Fhhu�	�*��]�7��J�E�p%H�F7���.��Z|��~�{T}�$`YCu9�NO`��nQ��Џ��|R&'��>����=�͕��k����`�� �_?f� ��Z�������d�i��W��5��YvM�u�����͊��;��z���{+:�,]����;�8�d/�藍����:o �����K���������F����w�RWAzM�W�a��`�x1ӽ�:4�
�\6x��҂�4ӂw"��8m��,T�
�WE`��)
������Ʒ����
Z�T�"����M�٦���rbv,2�s"oqs�:���Kvm�D�ܡ#�@�y}JH�)��i`�7�f�/���df��rq��=q���A��!>)E�M�.��kt*NM�b��6��.��GZ�{�8y)������eߥ(�&��j��\���+���UZi9�#�}r}iW�W|�
�rkb������=y��T�&�궻i]Yz��\�i��GJ�e�e�����;���X7��'�\�Q�X敪j�K��O��v�7�x3��^���{5q��7u���u�F&��s��荷N;�%��ʗ��Dr~�b)uO47ؤ]7<m�{����n�fM)�ܧ�yFf0�M6�0��=���*��	��'���jm�z�,+"��l΀�X�]����?��K�s��k-rU�>_�xhc��Ĝ��e�V�|H�d�}�Йݪ�]�9���.;��惍=4��;' ݸ�Br88���Ba��D�n^��#��K�3�v朎�G�I��w��|��ۗ�.�s9G�����b��lՊ�W5r�����2����\ln��<`���==��3�Dq�z!eJ�ܴ���O�r������w�}L=�a��)>~y
����Ԩ�� sޓgOI��WHR��*rj[�d���޺h2��2�>:�o\�"�ϋ�~N���-�ʅ�5`t��ĵ�j�.6XOas8��3	u�:ƝFvnrJVlm���q
/���)�������C]��(Y�ښ�R��W-c�C��'�7(HA��!Y�"9Y�>)��F�v�-����ڱ�#G��b�v#bxh�E���v���k%Wp�I�u	}R��}T��_�=��}rClˎ5�̧1ꫴ3zN%���ק靹H�F�+�mU�ܪ�}�=�����en=�ˋCk�SPio�+*�����%B��y6���JC.��)�:��2 �f��z�4-M����=�^����ў{���.ϩF�ku)�0�S�)�{{�����7�0n�=)i�6�,�Xp�|��2;��I�	wp�{|�;������b�H|�v��'ѯ��QϬsJ�B\�V�U׷eOf��ռ�ܵ}ʬV�N �|�(�eAZ�i�z�nɫ��z�f�,I�t�ɺ�Eu�������ؚ�hpQ h|�����hz�Z"뻖W{�v�f���~��ӆ�/!��s<൰w�W���7��ua��0���}��n�����|2�3�u�����׭cY\�m����c����ڼ�v͍҃��X!�4��u�S�/�,ٺ�7�je�IYUOOU�c�9�N2U�>�E'��U�j/�l��wgo� Gu���Yx�j�����	�U�Uo��(>���B2H5}��H��J�R�zʰ�kz�xk�����*���V&+b.�33�ĥ٧�\�$v�/X�a;��5a6[��vkk��͊,p��|�hа���©��fJ"ej�{�#�1,H�Uw��;������bS��X�i����d�e�s���>�;+�T��wv�R�CAV��D>�q��ܱ�2���P���N�q�ku�15y���u��1nwTE�Wv���)]b9�����{4���M^�QM3;)�9��9�SĮ���u��I�	4ă�u)������RᏣ�M[� ���mDE��G����EÉ5B���J+y�_Z겭��&�DV]�Cު*�^�;嫠�n�̱����F�ОQ^;ܬb��G
#r+�H�)�;x1ǹ˴����{��i>^ީ)��ꆃ���a�X��U�Ww���<ZWT�t����P6�!kdkJ#4�Ѱ!�5�U���]��m�����G����-�������<�b�\�GiFi��.�HYbk;$,zOk|9B.Ƹ�ɧ)�b�\'�t��q��}�2�(��M,V*�4��o����`����3:�ޝ�ќ�j#��m\���ْ�X>�+>'��^=��E�n�G���b�� =H��j�e>]� �{h��S3<i�7�.��P��c���&wh�U ����6=CR>7�xb4�{h��q	�1��^ TS���F������;v��r��T���]�yT?\T���oV�M��ǥ�Y�U�W�g���W��oK��;�Gh�3CC��t'0�n�\[�:�:zn��S�����6�#� 6������{Tx��YCt'0�O ;��ɡ��q�p4�i�k�e�g�����w�W����ȃ}Yo2�N��cm,^�bv�X��>�]�2X]~�[����)��;7=��g�V�r�@�w6��=ڻ�?1�A�Ꜧ�9o��+4�ؖ��m�o���,��2Z�ˤ�����[(nW�����/��S{I��ZA�����#�>z���W*󳓖���=�0me���t��p�=�۶�V'�f�WKܜ�
�����a#�G�j�}��`?o٫�=]�/�����:i^��XJ����x�]��\�\�U+�+��1pH�輭�b��^�����fq�V��ܯU���4�^�{���m8���E���p�����`��ǢT;�?3L�/�q����&�l�l�u��܁���y��3{�<eI�t �Y$��X�6Q���\C+z�;j�#��><�h ��E�Oj���#��f�����;�.厈'È��Ua��	���ڷy]��w�#WCdD�W�9�ҵ��D����8�x�[���W��X�m���D��F���;��(GoT3�|�,��7����M�hZ�b(s��pQ:���b�H���h��*�A���uv�f��*�Y��e���~�X�R�2�.��^�G�WN<��3�i�۽'��z�v9��4�FQ�3���4:��<��1p�.�o}G�Da��W}�ׅ3cu}�!��k��<IֱǺ�fc~+MĜ�r̷};FK��=9�v��gs�aV��˥���b�<P��M&g�7��%��ѹX)T�*�*���X�Au�-�t�s�1���E�������c��W��J��7b�U�5c����E�O@�̽�Q�QA��:N��ǽ��W�_N�S���R�8�x�G����e��wr��]pKi���h�뗅rOC�k��D��wSֻ��r�ۦI��E aW�K����ĺ�2��>8��Y�R���T�QSJh�
nbzY�B��Zv1�uc5�!K�N����]��\�p��S@�{h��t�o���}1��+��\�;����M5~�
)����0�+7ˢ@��BB�p^��k�����~�ȯJM�N����n�][V�C{N������DN��������p �:;�U<���j����V�G���|g� �Up�&	�Mjl½X�oN�g1(%3�%�c{���/I�~�I�+\���\���3qO>�0��i�A/Z�����W�����9��ec�G���(V�<��gWB��8(�pQaT�nGY�K�����)O��X�We�p�ߵ�=a4H��;lMr��
45~��Y4\�G����v]�@��ݒ���RZ��'���u5�S�z�J��L2n�����q[8�r�=��ktf�5���I1|��.�-���L�T8gT�'~��k�ot�[ss�؝�/����۔��r��8�5kw���=QWZ���h�'��� �v͍��iA��NK{q�����3\�d�$N6]'�Fku�9%k�\�e��G�[[�j����zYfs��5�����˶!��}v-˃X�7�u9�ϭ���{�Cz���ޓ_��|��+΄�8��a��lvw0�(�MS�(�L^j�+�%���R���j����
T&�WYTi�IV����+���ss+���D<e�g��Y��w�D^D�y�U��o�ѱ�FP2�M�HE!Gf{_J	X٦�t�r~����ͥ*�lH�ַM^Gݵ�.�Ogz5>"�u�;��J��6�f��`�L��ģ�w����w�eqZ��k\a�9T���Ԅ��@�R|/�o:KW�q�tmc�S�@�W$�'%a����꾏8۱)̡����	�J(�&��U"�+62�i=p,[��Wv����h^b�L}rCl˱�޹A"*�r��;ܷ�[�)�{θfs�J�U�u?�S�G\�U!���BCJgv]�rO6��:���2�+'�����SH�=�Vu�r��
�
$1H�w-m/V*z�f��:�uwc�h5��y�uo]�/���&�ߐz�Ƅ�W�νZ/�-"H�Jԩ��r5���$"u�g'�i�eW�񞔶V{�
T�ӑ��h/N��ٰ�E3�ry��W%��1��g_5�oo�j�Js��GE�w|^_rj�5�os_��+jΓ�'�/7\����8������V�{�b="*��LE*G�?�q���x��R�/�[���|F�����\�%��ƶAOP�6<9�xr=N�`E}*]L�R�d�-�ޮ˝�����?�Ӛq�7w���K9#�	��P@�F	0��)%��jcZ�{K���R`%��,�ٔp�����[�_:p��1�ޜ{N���v�`�N����,vB�
n��L�&�3��^�1#^ۣ�3�
��j�G1����*�����:�jПMںۧ������g2��&	�'Ѯ�뷷u�I���o�ԡg*,���#�=�=���;�Mv�'��F�61+Vv�GC6�>G&ޒ^�ƺ��8ٝ��Kob���R��9��wEI�k�B�\9�����"a�!Yi���er�w]�hp"��J��\"Ur�+����C�3�\��`��zr�n�a�M�7	���]�jV�v��#��T��xXv�)^x5������Az�r��3t\�4�fr{!�C�̀�ܔ�}R�oEъ�v���죵f޾B��|�����8dR��QT�C�ǒ��&h�˨}εd��Xs+/�f����[�u�X5j%�o�\O��T���P5��k�am������^Z��v,�ق�L�Ot Ӽ;����6�mg[�4N�TewL|�J��N��`��K���o-�
ۄ����+���w�V��\�L�����5N
�a�X�MN;M��0���
9}y(���vw34A�:q���{���C��맚�(�^#�͙z(2���������iW*�ۙe�i�oY܆f�S;2o�G3����8�=�Z��t8>V�y}���ֱ�)����h��]I�BG��󴓏m+�9�M���C���H��m$��Хˎ���=ţA�ƻs�62�2�@+bF��,V�30�]s��S��<Vc�E��`۷���)�{�t7#��9!yǨ#Ó*)�e(,�;3�*�4	6�V��N��TMgv;+Ck���<�Y;с<�Avw�=�]�l�L������D޻�uM��eڈ�]S;���r[}��N]u$���Kv^�l����|G(��&msQ�i����*;;{�q�Ļ/,�frA(�:���ɷb�u�Y�P�E��3/[��w�`�n<�A��xA��X�s��Y7��P�������Jμ���.�#�v��K�����u� ��L�8�f��� ��ۦ�ճr�4�\97Z�\v6�Ǧl_������b(�b�s����w���]�r|LgJ��zJU��D�B�e��z��j(ѡ� Q� P��	Yv��������fmͺ3FܜZD���m�bӴm	Y�Q$֨�5�;6��Q-m��9Vvv��ֳZnڲ,7:vl�[ma�K(�;��-Nv�8P��T�h�6(��4"�&jf;&͵�6[m�m�����ұ�kmM����E�kh29�l[l�,�t�f�,�nL�f�l��r��m��Mږ֑��VV�M��#c�2��-�$����n�MMa4��nE�؊m�mn�3��6b�'�d����Z�ɷg6��,[�����]�m�h�d�)�b�\]�n��m#�K	[k�����t�E�5�7e�ܓm;j�f�:6��[lض�@? ~�*�� �m�������r��ށ��$�q�mZ�:�;dHl�J/E3f�ϥ�vųp��[�]4Ԧ�>�v�-��������G��#>2cW+��v�s���L��p�Ey��%���ލԎ̤Փ��|.��^�X�=�������E��yU�)Mdv�[�u�ڭP�3,p�ъ���uy^��7���-s�aӯDL�����-(�\�Yhb�UruT�\1dշ'3�k��n\喲#iX��Ƶ�{���Bni��69��34�T8c��*�Vݨ�6��[�-7��^���Ů����mi���q������7t}5�f�j�V�H��{`����YTWa�(>���c-�f���pk��7�����8u�M���Xs���ŊT'��������J�Qn޲�Sq�y-�M񸩋zģ���ެy�C��zr��T�>���f�x�5z�}8�ΧJŤ�eo���k�'z����=�ֶ&���P���J��MR:z�3/��(�,Oq�l͵�2H��a����K?iL���qnpxv���X8'Z�^*��<��{��n����@�����@���R�f�r��]Y�è��Ӕ�mi��e��uY�U�ّ̼O��
_=j�<u��}�|�����)\�Q׳��n��|
#%~���s�*�bGʐ��H�����_ď-t�3�f_��U����%�G<��Jq��ް%�M�]%uR5F��s�'��le��SOj�w��&�簎>�"�2�@SFg�X�\�ݽ�s�yw���o3�BS$F�-E�@��������*����Ϻ�]<�/V�R]�z`0,n{��������X��4�S������N ��V5�;[g[P( �V$n"'����#����5sƯ��7��/wyE�6�����b+�MpQ hn������W�/�q�Vo��r]r��~��_��=��[B�ì�5�׸*��^6�a�Q<O �Z�c���c���<wx�`s�s�4eg(�fhhu7��/;J�6_e�WkW���rWW�w�of��A�=a����u�G�UNģ��Hqw�f�f�Ͳ�����grkc�',�Vg��B��Z-�%���WڦQC���c�}ß>6��rn�-*N�a���������̂!Dc��[���s_wV֒�2���],.����}�����Bʵ���^ĕ;�֫Zɼ�W�3f��k�����C~�H��	k��B��(>���¯ɮ�"k
�Ⱦ��#*}��b�5^�Y�0J�N2�&���v���i��ܘ��v���3���Z���t��of���͉�u	�ny��q�h�cVDj�{KN�:voq���
ky6Z�)�yٹ��)Y��PܩМ�8�1��\nZZ��ҔJ-m98�o=�M_��Q	��Z�j���?}��SM)��j��̮�/BQ��
N�H-�jo�:�ھ`�>�O�	e,Z���X{��cFrԮ:��U:R�y�+j����&���챔C��봋BwsE_Kn�Ab��,$j���c{��U�V_r���{@�{���;�r�~ƱZ�m# ���S;~�D���m��B��V�˼̈́/;T��������g���:�Z-8�!�čl��]p�3�lu��X���VEӬ����	��ڇ���`U��NΤ�r3ʇ�O�n���˂����c�����P���{�.[7��wD�4Վ���t�c�e�H���m>����ɒ�K�:�5Pޙ�\u; ��-�I9��}Z�V��X4��R�y�iEV��.��7X�vƨg�&�Z��9�<�o��m��Ou34)�d;�&o:r�g���{�Ǽ���v5�.���x"�����$��\Oq�g\.�;��;yV��7����s�`��4C+m���mF�O9ˢ[���{�XH�ْ��/xiuD�Ҽ|ln��z�[�_T9�IN��s��2�Y�6�ڢ8Č��t�8��a�-�}�7��k�t����k�a��6��+㽪#�N�0R�t�VP�vw��4槁��b�çw�[y{����׭����� 7�{�ڣy�(`�q�|�*�d@U21*��xa�R���S"�>�a,�|�e�e3�yٸJU��ŧ���̕Y��Z�C����A��@���l�obZZ�E4ϡ�bt���K���#���=3��]yMS�Qސu�����Ս`������k�>Ő������'Z���<^M�\�Yіj\�N�gM��+bS��[t�R>��>䯙��u�̓��8�o���~*�UMe�В�07��M�[���[�Γ�;F�8M��Rڷ�ݺ�y�}oG0M��ޭ�3RVvcsz����gq�_9/}^^0��<�v�S���$���}k�T��p'sGix��--��F�����.����J	L���Ee���/�u,e�E*\�+7����UO�<���OuH~AH��!�F�0��Jgo���]��~�����+�|�J���e���r��PP�a�s_t6��
��K��#y�vq��(�ū���e���b��Ko�ۈ�I�''K{��Cю���]'T׏kw�z�V�M���`펭���wqV�k��vNg����U4�_��4�?9����c]zwQ^�B�M~���u�]�:�Z~�W']Mpu�5mث�k!rU�N6"I�Y;�)YE��!|��sO��Y[�fkC��3)�y#�u�K�ޭ�d��ç#m�w�%տw�����{Tx��Y�:ӡ�<	�Pk�f�{e�hLC��6��g[�K���o&X={����\Z�Y�K|"o\�ۛ�E{V,�e���y���2�l�⻹�;���������R�aΆ	x
�rk���[*T�ԤݘH�ҵ�X���ڑްL5t['�;�-^�~�e]eW��"���=���t�n&���k��l�	.�U��.��r�ºS��X+)4��J�j-��[��M�P��^+�1*���7ۜr��6'�W
U9M�r�_RV6i��٦�f��i��vK��Ȅ��T��]k��:��gg.y�SDW�6��o��Ƶ8���5r��k���1[Ry^�Q�(j�9�68e�A��,�4_wH����#S���ը���%�Gp{֭��w����-�0gE6�RK��;2����u�K�:��V�S:��H��G\�i[�g^�U��֡�P�.�y:1�[	U���cڭ��ZWV^���⼇o�i����'����H�S��b�#Z46N"v_+����+]������<�gl�k����U�S�A�1T��E'���V�1�����m�y�j�t]�@�s�
6F�Ƃ�f���%�<�o3`-:�p�B�I�+j��\�,e�9��qt^}����ehpoFEEf4���Şߞ�1ӭ��'��.�l<��s�����u.�T���7�ܪ,؅��g�z�{uJ��oc�Zh�-v!؊�S\H�	��#6�`�i����W��n����Å�V�s�{m�׃hc7�Ci�T���R�y�;�[0s�ftU�uj��SFճ~�-��R�h�<����C��V��1�����<}(�*�s�����^���s�oHz{��o�X���t�7��eU1�$pyC*�U�����/���{w\2�c�c��'��o�_?��nW"�N2�
ʠi�ג��p�#�0�*`�N��K��U�2���{Y��͊��gZ򬜘�S����Cѝo��9�a���v6i�7n�)�;7<9%*�N��Mg½釷�>�xF;2���FG�}+�Gb~�NO���jưQM5bZ�~��[atPzM�z�f�wf�5��b�������L�u)>�)Ձ�ڱ�#G&��G��͸�x�K+(��¥��E���z�ͮ�/���.F"�f��9�An�sY��T9��+���W����@��u�Z�G�Y��U���}�Ħ�n��iP���|F>f��)tC"ĭ�Nk��ئ�fi�K.�W ���y{�&�թ�!FĠ���ԥ��ڪg�����I]]P��V�9����?[w%����!{z�����j�ѽ�Qj�e�j�W�B"�X��J��e�;�|��>9DZFAA/j�)��N#5ve��X�jm��j�#
�޸k��WT�����ub�ӁAb�#[]]
U���Y傫Nf'{,�@��d�$�Tq���j�Z��͉�3�A�Vh�J���촅��쐰�Oiy��qK�8���=��6�sɛ�����gGKኦ�+yBۚ�ѽ�ݎqL���D��m��Y�r#��g(�S�M��s�W�.�^2�҃&E�G_��(N�;�����k���#�G�NU���b����^��"���gwk�{�����͠ϻ0�Ms�Vw���L�J���Y�}���{s�&�(\վ�?�<_g�i��������{��xf���a��M���`�}��www1���@k�s�R/r�K���#'�C�HN��S����t�F�*�W�	ۘ�
�#�������[/�����EҰ��wִ���¸پ璂�L42���f��ڢ/"G��`P�b.ֺ]���^�s��u��Sݹ(%cf���v�a�^7�<��r�e�芜��>��ޥ2�Փ(*`��E�%{4��l�W�@M8�1,N�}|�u�:t�6m��2���"�+���7ԛ]%�w=��euU����](U��a�V��28pޠ%�S
QGy�P8�&tU���ަ/s�.*��J�a#�G1���.�c��r�DU>����^.�=�������߱�UO�R�'��\�U#|����I��Ěh��lp/o6�Xװ�*��2Dj�cU��i@�P���r���t�W�Y�36I)sA���|0,,�#�P���Lk�cڣ�ޮv�����$K`Èڒ�6k0]�+V!�n:'�*��WA�:���n�B.��.�5�2��+*���#+oU�(`#%!�mm.́5�1/��R.ӣH���l\�e��1�]-h�r�hDM-Q�v93ǂ�4V.�ծsu�&��	ZSb���l��a�:�_���Π2�ADDa���Q5�z�C;8��D;[�������7u�E�\�NݝG��W�;@�tb�&�+�ʶ�ޔH��oGtk��I�7ܩWbȝɩ�&�;�:�:�hpuC�*�շ~�ͭ��]߬h�3j�����wV����1`s�m���9�gh�3�́�B��4�٢w��g�OI�.��xS��A��@�֐��c�WTF���;ĩ�9�p�#��a�����A�k��)Wf�&Vj�Hl�K�Ԭ#���s3�FX�QeR�Q��ܭi���X�[���I��=�q�u���r���C�}�X�v2��Vu	�n�y_RW�m�W{ݻ��K�ެ�ܧm�=v�2����Gl��T7(Ho��$�*(�R��Rͭ�]�!�e��E4��V>I	k��63�7(	>�.7mNv͗�6�x��Pw�+��RE�]W�W�j�b�����V�>!$ I?�	!I��B����$�H@�~�$�	'�H@��B���$ I?�	!I��IO�H@�~�$�	'`IJ�$ I4@�$����$�`IO�H@�~�$�	'�H@�~P$�	'�$�	'�1AY&SY�dJ'E�Y�pP��3'� bJ��w          � �� �F�    �           4   "�4�v덟m;6�mX�U^��XF3l�a���L�5�ֲ�!������u�ڱn�]M���֝۵6h��v���e1���Ńi1[c����;�[4���Z��m�Y����j�]rWY�e��"�Sf�ͳk1-fƖ��͕E=n٫+�vL�ۮT֕�cZ��uܵ��ѕ�&��֎%N�'֞�+�.�F  �=��i���W�׳;��un�׳׽�ֻk���z�{iWB���[m
a۷���n���jn��ޕJT�������6ڒ��C�W�6ۦ�{x��w:ٚ[z�=5��[n�ւZ��/wr/w�  {{���ݻNmn�{�zҫy�={J����]ݵv7mJ��W�[g\��r���:�^�p�D��C��ǽ���ې����z�l��jZ��UJյu�\u�6!�������U�K{�  =Ͻ���l:ݭ���ޭ5��:�oyLWz���V�s�U��3��D�ڧ��{+���d�ivm��ۖ��mg��/� ����({���(P
�����n�}
(P�o^��U�ɷ�8ҩݕT�6��|  u�
 
  /�˼B�
(3�xP�C�hP�B���B�(P P�����t�x�e�m�Q���J���=w�awUK�6s]��=��U*���{����u�v�U睕����C6m5CV���3�  �l}���X(P=�N 6��h���f�ҁӽ�\*�M��p���{ݼSA��L
݀����{WG�u�Z�ݬ-�d��f�s�Vڶ�|   �hP��� ��C��z��r{��q�=u�:X��ˀ4��\��1Z(Μ�A�{�G�su��v�L��2ʋme�|   {��Z�Oz.��r�@����p�w={U�*���<:5��3��=�����F�mP�d�:)@f�m.SS��h�[3-S*v���  �����z� :��hoO+�kݡ[�/]�ۗ\�j����ٺ��+�y=�ڴ�[^z��eWmK����=N�;�^�8��eK��nY�⻭J�U������le--Sfl��eg�  o}i��3v;|y�׬�J��wz��ޚu=[Mww��-��n����T�n�v�ov�Պ�m����z�m��=S�{oZv�ʺ��zUUjZ����y����v���[e=Sk��tZF�75�m[Ukz�  p���]�R�=��#m�f�]�u�V��.�v��ַ�Um��՞���f�j��׽�{�٩Uڷ{ٷR�V�۶���c�Z��OgOomv��]�/=��m�mv��S��$����4O�1JU&� h�)���@  S�%*�=   j����U&� �I�U%�2h<S�?����?����n�����bK���q�B��*Hh� �Z}���6N�:���ꯤ��S����$� ���$�HB��@�$�� H%���"���������7��j���4.L��Y�M�r,���t�v�����dS�����ޕ�x���7,��h��>��K�3�a����w&+�[d�t����W�"]������"���^=�aU�T��İ�2j\Y=��T5�F�9�N`�uh�x��=�*7��Pָ${˧y�G��v�#*U��tS���N�'X�[�-����^B�u<:ݷ��H�s ���*��M6�M۲��Wo�n%0�j�t����)P��w{I��njۗ��JsZ��wp,���#l�rѯ7��`�<$��g<��0���;��'��,�k���-X���Iᛗw�SiK�7��"��Q�a��縚��C<���yh��:ny��,г���Ƀ�����t��X�x���8 6��u��C����Zy���梴襘$oW	�7���=ہمqq�3ai���Wr���ƛ>+rWI�p��P�m�uf�Gk�ۧ[�;��Wn���4�;u�N��ΐ6���b`Z��x�R�n
����1�%�)@ ���M�9`�q-ƣ�=�[q�\��[�Zzn���3��3��4M�h5��GQ��gG���1�s ���K��a�V��L�t�۱�rqh+�	���a��X\���ي�nL�4v>4,�r������`����l?WK<�����sFCs�i[;�ԍ}F��m�n<���r���c9Zuu�q��ӥ,U�l8=xoFp͂k#�=�;�r�אBE�愅[�سAy�*-�;pi�d7�!�l�rҴ�]�w''���u��n&^�o��`S��ǭK7D��I���R��a���SB9�7���Y����Z�(��aN(���ľ{'��3��O(W���T�$���Қ6���]���Ň��.w��}�nq�fk�� h� ��Vy�Dy�IRu��q�W������\���pgR��hV��@-�xJu �/ \7;�t���z�����hhɍ�DU{�����ˤ�sWmڵ���{c_}��:6eB�\V]CssvRV}βȸu�yiQ<�^�k����ΰi&8j���4dwP�vu;�Ĺ3pq��r���_L�.��ͯ;���뇣��Q�H��-ͽ��3�%�工�*Pн�2�D5�Tw�.sJ!�"�X7����3`�:�UK�W�&�]��0����lhvu&Mf4T]��]k��fm�D&,Q�^��#SN��3�M]�ڭ]p���[z�d��7��ݬ+_m�m�s��w�r��oSV�u�3Pĥm��N�O:1,C��O4^�����_�dò�7O�n=-��>A*��|�f��y�&m�&6(z,\6��ojK����У&�V�Be�ږ�.l��Ԣ;sR�2g	�(=�NwoDM����,�B�me����S�U��.��oN��ok��I>�`��R1e�%oT��ov?�t��[�u�5p�B��`xOn����b��7�0�f�J^׽1�њ���;�<{*�7m
���`���
(�3��'sN�0,��gG�puӔ�ϗ2������NA�p����)��j�\4��:��N�=���Js5{D�:�����=����h.�;]���q�Ӗ[IМf���.0w+��q\�z|wu�q���ܒ���qTvR�O:c�)"�SIfn�뷬 ��jc�(�ĕ{�kL�u@+�JsO�������D�kW���/+R'�=ۯ�灺���\ƕ���s\�tݴ����p޺ ᓫqp��p��3i�g;��-RmKN�q�b�@���Y]��#侏n�+ �>�tM��q3��Jv捪1�M�m���^�i\U/��0�{��n���B�9|`4Y�VSEZxN+|3�ؖ<� �s���M%E ���U<Nu�;��̔p�U�s���x������7��8�Vva��,a�S㪺����`���4u �il]�>,��T��K���5&��ֱ��y7;�pݪz!����>C���r�%7yOBe{|��)�w�t����}Wq�vv��qvN�Ն	J��z,%#�:>�c�T8u`�0Cھt%b�Ypvu�U�Y�/�#tD@�����`(����p�d�x$���{�",b�-F�\ח^�0��x��F��������
��󁳰���ۀ6u.�G>*|ٜ�)�oص��	V��P��n�u[��c�y���$�Kب�O@�#j�i2p�S��.�<"=ݴ�lZE�@��ؓ�������GE�.����e�\��V;yw���M��lkU����v0f�eW���xαEƫ�.MwvRx4%n�J�.�9�ju٭x� w2T�#W��,Oh�x.�s^�x��ׇ�+�����Շ]�����T�7]A��I�\7z9�7�l��SD�I������ui9�%ؖ�.�o�PN�oM8�\b����CJڳ�������+��{5��v�T�a�!�4���_�]��e{b��᩵O�����>��>��Ku�a$�ɛ���.;a��޹!ދ�I�3Nٍ��,��ιۣ���L�2�:q��p��#Kx��Tՙ�;4��J���.�7��ږ&�Ǟ��VI���l�k9�(ڄc���>���ٍ��Żr
Ć%�#�3�)�tmk:H#a��NY%(e��i���2���UU%y�����NqT��((_4����C�Խ*�n��G2�/]�)����y���Y���mXe�Q;띡��$`wtՁsa�b,��:��(�͛����S�<�rɸ�,k��r)AΫҖ��iyI��nɩ�˻p��P�5y/�P�ަ���IΧ;F.����]gK�.o���T�L�b�ܘZ��W�bZ��シ���w{Th<Y}�j�z�X�G�lVL����-^'��4�هS�.��s�F�tl�xP�)���[�sx�p%�sg������EѮZ�j8�)к����|$�������gYK��U��!0�)p�{~�����lޑ� tYlEY�W78Y���xq�9F�l�YZ��.��]k	�O ��x��jV�݆ɃB���r�m]��Eb�O�/�wR~��Y����B��M�]��,��e�F-7�:6[�k�{7���r�J�o��8^;�Z��5�Q�$�w%��G���y��خ[B��R���I:n�ۗ>wIq����ݒrD��c�������`b�,�t�޹Bn%���hP'��᰼�&GB<ksE�D{{5��F��s�vE��z��]�{��gP��;�����"By�±j�3���c%\����
ł�^��KGZ{[���T�Hb/>��F�6���b�P l|�X4��!���v��5dg�
�9v�L3F�����'f�o�46�M�N�����2L��ʶr����ר7Nq��D��")C"qw7�S������gT�(�V���0wU�������(�\J`��&�P�D�Ȁ�Dٛ�.�@�f��v̡P%=�k�77n�pl�C���T���,�:�xI�OQ\q7Q\^V{v��Ӈ�.R� WV�ݗ���K�+�{�m<0決��߃�vh�y�>�/*s�C���5�%��W�����74��&�����v�)��S�T�w�'^p���P�j��5c :X������Ж 'n���5����x��6/`b�k��{$2��Gj}kش��P&�rC���ٛÞY%���LI�.;T\g^sj���{��VK�B�k_bc�C��B+��mwٕ�9n&�)�[��)����#�H�XM�ڳ��l(�^�;�tS��~�-��äd�V�]8�sI}:��q���
C4�c�3{��62r�S�Q2��f���J�qG�fh�uT%≽5����o\�V �WW\:�=��������]�'��ni9����V���ա����x���9�z�eYD��̽^����7zh�/t�kT��"���Su�l@pu���^Zay����Z���X��Pl뫈�!s�39�T|-�����9 2I��wY�x�a�H L�[�LGݍ���m���H�3p����뢵N�u�p��ƚcۜ�p��	V<5 JМ�x����6Mzs���k��eyK�~\#�~�Z*��.�I�J� �B0��"iW{�aX:q�6bqq���񨀱n��N�6goA\3����@��8B��ȕу����P(`��5���7p':�/M	�l'��uh|lz0׶Z���:9��/^�.�N8��Y�lm��4W��p�O{�4����;!��@jC~�V�]��"��1���jН�LU.���כ�%sOjE;�q�oCaen���f��I���B潵�<�X߶���XL��F{C��*�gNuۯY��(�%j��Dx����]�ZE�٨K�hyN��v��?5����@�ͥå���T��᛺$ï������1s��Pǡ0���u@�_��rk�ycX�H��{nUz'��,��rv�geD�a�h;��5��{��˛*�o�j&��\Ƅ���,��-�E���Z:f�,:��2�f�4+���F�����A-\��.�z7/=�18�U��TŌ�b=���tQ��;^��N�U�s~\�7n#�td�;���5<�Fu[".�3�(JZ���oHp7��o'��6�9�	
���Xz�ȣ��yn&0-��U�C���\{���ye���"���2]6\�ٕc$2�Ei�goiL$�
(��ˢ��ۦ<\7v-q�$�
���-C�,���yH.�.�jgW>�.�Ҧ�`]�{j-uևCctv���Yp|q;FAo3v�Ӗ��$s93)��7:
�ɧ%;V-�����>�L��'?vⱽ��2�#7\�)��W{4��C�4�7r񠋤6v�23^�L�~G
�0�C���q\�oK�2��J`�b[���V�>�qy۲<[m�sol��4����!�x=}34 @FL9��p��sὺ�ñX�'^������u��hwov�};�3�QZݹ���qh�.Á��ԓkս�����yf�"�w5����nq[v�)�c%@@�%Niv`�rvT6U�)��wa��c��WW�q�k����vm�#��,kHb��>,]o�����ŇiK�!��&LvH�����ӂ�s�^1"�ns�:1��5��%�h�D��4%�"��!�nM��c3��ٹ02�#y�f�U�d״����Х[0�ҍ��7f�S)�go*�a�v�Ml�-$R���k�L=�;7�ֻ]9Af���!���4p��QJ>�6	����$x=WD��<�:�u.=/�X�v�%�˳�0K��W�;.��=�Wmv\ܸ�K8.8�pW��̭�+����b(о��z��I'��6�ءط��F�;��<��ӫ2:W���6G������m��uݐ
C��V�c!<��D>�@�4��bN���<=T�<nZ��JpG�*�$�F9�bqn�S����0�`�N�!̧n��l܏8l����S�M�F)�0}��읯w5i��("�y1�ù(��-��oDnd|����23�}���xfێ=FL�v����9�6��_jD�or@��������Om<��V��­�S[F��u��:b��\8{������pj�`��)ӡgp�>_sYۧ.N����w.��T8��3��V>l�Wm�6�K������=-�nE�"�l(���9ۂ��/Z�P%�]��Ut�;+���8��lD����t�Ax�S�8!�L"��D)��^��������� ^7,]�˙B�v��/v,(�֘cZ|��M��� ���)�i\���j�M��{q�Ӽ��HW&W&���>2���՚�'��R��j�i���l�a4v�4�v$���8t�w���3GW3p!�w�ઘ��{V�����>Ǻy�:n�j����I���Z�y��{x���InwM��A����iͦ�;.��Zn0�W���Sޑ�۪�+2sU���
�z,Z����
ǋE����F%2����4��jC��O�-]t�e*q>闶ػ	k ���� �}�]�D�Ա+@4s{�^[�^��Y�5�m����2^Њʌ8&��
K��U�y&�+�qLv����՛�ۈ>�j4ͧf�^�[�c�t苸8��Pǹ�}��j��$�D[q��B7��6�9��6�L�3���h$M�Tf� �2KIm)���ի��wb}sw��D�&�s��ÕHy���w@Y��o����T��Z�ݿwq����H�,C���!�r�v�����k׌�y=i'[��R �rk\ؑ�3,�#�`8�ۄb+{"	a�b��rū.��wx�cf��p�����qt����4[�4��2�\��)<��P���9�JS:0��H�x��.��]���+ˠ�q��s�s��h�7\��T��I�f�и��^��e�P����F��a�{�<oq@X�ڀ�`�twu�� �Y���ūZ�K��Dh�O�u���l�b��B-\e�OZyu�����w�]��yX�����(���R���I���i�[���+wӅ���պ�7n�Ϻ�!n��F��7g��O5�m��h�e7ԃ2���i�a/5康wNoj�3�C����(�S��F����O<�=f-4q/rhc�^�FI*��`�j�BЬVV1P	U���n����f:`־�i�T����*�ղ���i�F11��<Y�{�Ԏ<���D�\�=���F	c.���Iz�*wX���ֽW��Om폮^-�f���axu]��jzf�;�t��yN�U�������]�gʗi59e��{S�%M�ۢ�Ks�9�'7��Mz�$�wDKU���k)����ȶh�����cY˭!��T�39R��c��CK��X��P{}h	ZV��V��(��ﻕ ���/WR~Ǘ;+\ڷ90�������sٮk��������TGG�VD/pc��ܱ�r��Յ$7;��aNn��Zt�aͧ���N�Ob�F�ް��TOm���Aj�2�mU��*�^��]!pU�j��.R�Y�8�]x����%\L���1�u�e�Y�Y1�Ш���g�ҷ�����X���K[y���*�8�K�ޤ��b�+mV�j�u:S[�՗viKζ�p[1,�*t������w��:�:��ɥ��+-�Q�د.�r�]f��@�S�g:U�Sܘ��N�ZÚ���Z�z�*�{�o[}1t�S�h���;g��i�I�A���t06v+�j��]�.9�������a�*ݍ���$�I�h��;�%��c�[�5���i��^rght��4D{m�͘2S��s���ʲ��RGF�E��~P��?{g!��k�1�;9tQ�©�ɓ}<�y.cɋ�Gr�ݡ�jU��{\�R����^����.��G[z�%&ml�B�:^��w:t�r�=�OT/�*�\�וy\S2B��+������[���w��_a*'i��Љ�.�0gPs8
���X�޹[��&�v!i�����Z[������C \��w���9�]�VAG_@{j��g-��n�9cN�U���,N�����j^���2�mR��Mw����(�b�k������ۏ^'��S�1].�O��-1�4V83.���|2�Z1�
a�5�	׀w�h)�Oh^�CCdl��ro��/p���e����9せrB���f�ϰo��Z�<��U:a5�S��^I����(��
�+V�K�qLѢ;�ں��J=I�Lso��V���3�q��B$S	����)�5�"j]��n�뭈}����+�[�!�D������͐�w`�{��yw4�����%-�����9�����/Hq��G&z�#W�s�LQ��X\ɭ�H���9h�ƚ�W��_��q��uD���r��H�4v�����^wBv���ʻ��kUi��؎sVszxV�ѭoJ#�7��f`r���ܡ����%u$��X��[2�
������K��Ae&�ʈow�k�!�@�3ف�Z�e�]x�i��H��2g>��s�0t�Y1zrڏ��7�C�>���/sb{Wg��7;]<��A��J�s�\2��"gB�L�,��u)|����wT$N���I%�%�
�m��2\h���K���w�ӭ��AFt�q����K�`]׮Q��d����d�9i�˥n'���'1<����R\���X\)�r�T�e$rӐv��-�7s��}x�U�"xB��tߥ�&���u՝p����,��J�ބ�x/���twH(F�H��j묻M(�eG�t��ZC(V9�f�dY��Fjun�Q�3Ap�:��W9fm=+��-�#�,?�e�lSv�}�Z����
g��E��]�}9隡���������c�m���.���y��4ʞ��z��n��-����(evk�J�g�x�r�mb��31����(������R�q�:șD@֢o��ݩQޝK��f�/md�Ռ��co��ʓ�&�+�r<�V6\�X�p�{�q%ͤ�n���klZO���.�;�J���L:��:7:yf��RKe�^�6��d�^3��˜8����@S�<yZgE-��
�,4�sO��O�3�_S�ĭ��F�_-P�1�B��z���YH>���ýt�u;��ޡ���S�g'hz5�T���k&���� �VJ�o�������jy��?QLDw4_����h[�`#�&GY��S��o]>�+�Iw�e�g��`�>�2�Q/��+��[�1�ҭ�G+�
"�

�b��-$�R�My�hU ��e<�-8�7�.��r�h#@�疩U�u°h��3�;���Q<��C�n��M��B���:��$��i\�^V
��`cCF����ip��qw�v���9�aF)n�]��]�ȟq�F�C�ua���]�nݛtˡw��Y;�c:3y}M2y�l�i�ۿ��R�`�Y�;(D�U��f��ܭꢏp�8�b��2��v&j�X�7�̲��ӡۏ��lQ�{[�&���o(��ئ]��;���a'
k�Vu��+�uѦ�V����@LFN�Y��˥�>B�ܥ&s�Ms͓-�so���.Yؗ{~�^r���!|
���<�|e���g(W^�w�I�����b��P��<����Z+x��??=���x�M��rr��Mj �չn&�e����}���7�W��^�jjO�H����ʺ蒪F���Ĵ]e�?,tK7��*�h	�,=�~�8&S�SO��	��W���PG"���bo�	�Q�����j�n��E��7(��)��Y��Pkr���y̤��~�9��|7W�v~�1��ihQ_Pu�R�OrV��}7�A9�`���Q>Y�Q�1�3�0����|����=J��hf8_�ɋu�õԖ<&�0jR�0��żq�mî�COf��sT]���\ںv�[�hL�zMF���\\�rCL�F1��]�<a���֢��yݓO7��Y\ީ;�;��A�B&JFoO�������՟#��������]S&�e��d2��o/�E��e�R�$����q�5���6�����i�D&W����S�[�s����y'��11>�+rmv��ֲ�~��]�63gf���!�گ)��ӛ+Z��9�eRW}]R�i�yx��ptq���K!e�v]�i>�Y�|�R��ʽu.>v�d��Z�X�LA<�'-�!�x�S��f�5F�%�Ot��В�l|Z'0$��	�3T#8�u�qV�iQ��D��R���c�����K�9M&�lv.M����΢2Eh�2E�W�#�<�fÏ�%Y]�6�4�ҙ'Q�T7"�.�Ǣ^�W�y��c�i�ܼl��o!�t�2������|��X?1�2���S��u�Yy_��:ٰ����x�����ف� �i�F���y	�W9�Gz̊o��oV�G�r�dL�;�bV� .�֌��*�G*.IE+�K����ɋk+�Б;�º�aߜ.U�B�4��,[�����׼�s��*e]�������ᶳ{Wb$�ŋm�&����*Σv���bx\��Ucv��"��7P0�嶩en�p216���",�4����ja�|,�D�4���*��!���7	 d�;umt`lʹK�i�/�๪DC���u3x�����i�dꕛ@�eu�o�L��&�A��8�Sy���d�UH����y��`�Z��3�n�lp����3Fko��xH��Ru�~������kN��P��'6�%��2��&�Y�ޣ��_5z��n�bA�wj�'bh���7l��1��UsݻH��$,W{)B��[SD�m��v��R��/8;���r���yώ�� �ӵX�bl��:�s�>��J��ì���9��p��B��Z���ؑt��RM��ym��c��X�r����U�e��ɽTڬ����W�;&F6vgg)&}�V&�ߣ�|����z*7M�ج"���}��,�Y��X ��G�B��{��e�ك;n�77�����qn�k�]F��_y��#���`��;Vݾ�ٷ2�N˸�����<��2�S�������]՘;H����*�Ϣ�r4�,4$���[�u\-����t��
s4���;),�2�eXŲ��-l0�hM=s+9Fuɺ.��<��̆W\�(��3َ^��*{�s�����]��"��Ի����5A\���S��˯���dGv���X0M!���Weq�}.7C'e��]y�85���Ǝ3�`���_G.s��f�A�6�Y��)g=qP횓LM�Br��l�؎K�>�,i&4��-���r{n�� ��[��������w&%��:��9����njQ׮��sB�9��9o�+��"cp�ڀY�;s,W-���w��R]17swu��{�,����QZ<�b�;s7����Mi��w��i)�^A��ہ����;�(v^Gn��G%��a�\�}0�iIr�Y/�-�qa��xsk�kY��Y�kUAd˩�s��[��MűL�/�zr��4i?0�kޖ����v+e�}h��c[����P��x9W'�+M�"|�&A�@�`�M�:����k=*�4E)X�{$GU;,us&��+m�)�g�p�sm��@��E����yR���"x=�;��r��[�\Ky<I"#�I>��ڠ�y�%cM�(]�\o لЂ-e������2`����n�����7��lz�9Z$�����X�9�j�b;�^)�Ɓ����-8P.�+$���9]�5Z��;u.�;R�+�{sv��W5FX�f�F���l'&��pw����,`8�o-r����Ruu�9{��)F��R�E�1TBTpu���d��PGf�Ya�G�ݖWaƦ���gP����o[�ٻy�q�%���ZN�+,�Yծ���n���Yu��^m�����j�F�L,��ڔ������{?��F�h�gb�ѝh��]�^���u��÷ ���{\�R�I*u.�x�����!c�^c��]�2�LZ��f�g�"^���QpW*7��^�2�ʃ�aQE�q5sL��L����L�sX�k�m��m�'aml�3��D��ˎ�u���ب�[�����E�����ג��5Kof'{�+�c`�0�$��O���z��fe�i4u�')6�K�
�M����ș�*۟$�9��	[}�ٖ��L���K/F�q��`ۥ�f�ғ�u���v�S���U�RB΄���yQU������{�m�Ys����qˋ����^���>�#Ӝ�;s��[*p���L ��/�\b�Eow.�a���X�Bb��M��41L[��T�']>�;��,���T��Ύ�oQ�5�;�x�0i�vsr��ٰ�t5��Ys��fB�,�{hw��Y[I�;��J���;t�G���x�_rt��*u��rEƋ5<�*�91�v�h����*ܷ��q�˸�E�|��L�:�(L5)���c�[��\ڐ�}r����z�慠���Kh�}�1��_��b�GB��~��c����6���v��Õ�	i���u��Go�sx�!�U�w��i�>�] ǫFH��ٸ�xX3\����hk��3v��)�+��v���_5;��������r��}�� 
��ǔTɵT:k��4��7��|VUǍ����MYɸ����'n�.�g�g=Y0r�5���0���x�1Vk��Q��$����!gm�n�\��Zk���Co��V�ۚ���[�n@L��Q>���L�$��K;���$�ξv����F���n2�/eJ}q�Oo#�������L�ݗ��B�V�C:���J�r�W+�>R2_�;�y�,��ɜ��k��o��z�'W\7L���;{ƣ�XH����)��Fu�����+�Jo.D�t��|���F��k`���d�mK_���N��7\؆&M-�i��WY�ޚɘ�AݮF��Q�Ӹ�z��!7�:��c#H�����ڞU��K$T���-���Bi�30\m�Tݛ�{][|5���7��h0�	?f��}��v����ߖx����ǀ����U��u�
���,d��B��a�R�L��QE\�u���bV۶.�ɝ����A���AP��j�.}��uk�앵t\Ws!�����.�軻��*�6� �H�-k�Ƌ���i_-�Ppk��t��,ٮ�:�bnd8��j��4����8)sEřًk]��[p�:��3�O:�n��M���U�(��%��T��|����=�w�~�y�j�Lڎ��<[c!�X6��&^�i���*�Kafj.��Qy��a�n{��T��6j��7�4^�\�ڵ',��d{z�
7y8������B{wԙ��ٶ<[��"	���]�w��BL{o�-��� ���{:<�W��N���'4��|�u��-�x����m�9D��ݘ��눷S�c&��{X���y�D�4LǏcj֒K��=��;J�O�s���F{q�x�eD�r[~<咀|_���7�Q3;f�T}����Iɹg#�q�>�I�"�̧��4�˽�w`v�/V���,����"��_Q���$�Rδt"8���"�YA��v�si&��#�̡;@�7o����k��[�
����+W�*��6���x�͕�)E��5�X�%��9���T�^�2�t\~����\g9"\4�GY5�*L��m���Ղ�m�:�3X͙Luh�ᳺ�����Fb�B���*��3������<< ���?��=��{��~��ٚ�؋׿FJ]�z"�n��f�p�홯V�52!�����kg��h&L�K����k����ڻ�A��)�
�<<�p[.��Ƴ���_A�f�W)��$�z�AA����>���5�:t&J���*fT�Ll�|&9��ךҍ}�p��w{�f�>�+�w�Μ�B�	��z�`���&������s�j�j��sM&��X2�[�
M��G$�A�U�;����1p��� �]zi蜻m|�&�^gc� ��K�1�#KfZ�D��S6]KgJ�g����f�[�2�J��噬�C*�q�l�ϧo��]b^�֬5��p�3�R��NHdsk�:�do��I�s�[��[�-�^9�p��<��9��/o�+1��a�q�1�4��2�y��t\�̺��7=�ڲ�-���4sk�w��ح/fLз.��T���e9�j\b����=2ę���b�h=d�u e'�}y���m�7���׫Go��:'��-�`���{u\�u�P*�+��	S�Y��m<�Ҧ>�݄"v�퓀�v)q�S�bNcN�5�c�t���R{ݸ�*�`���]U�='r^$)_X���"wp�SĦ��||B�˳}�+ݻ{�T�3�q�ͺ{!�2��X��Ǵ2�\&pd$����^��j0��k}�&f`��u!����w�Ǽ�?iF=V�N)ZD���c'�a�M�h��ț�u�����(Vs
r�]�k�cr��V���� ��+��.%Һ�Q� ��ѭ��1ޚ����r�&��&�jM��md�vP��T����}����9D�J���{�N�&�0��w�����	O�,J�ΪJ�i _Aov�Ѻ)�hhMgA{xR^�P��ž}��Y�{XQ�^W��۫5�Bn>0W�&�/@��ez��߬۷� �<��G@R�gwi�4������Ӛ�4���K0bї�lf�/븇9ԞS����)���e�۳/`��G���٣\��*rGA�E�U���}y�VKw�=�˺)#9�:�!�8h�`[���x�/�H��B���h^>�>����j�����8*�tpGI��ܹ��:��;���2e�z�Toi���b�G\ı�,������@��h��V�d�8b�'l��w�R;݂g,�c�uʘg�X�� zs����}����I�P/���DW=#>{LL�P�R�Za۷N���{��q>�i٫��4R�<.�Yl�RF����,�®����V�V�s��mcf�l*�!@)�[���LM;鯺��Nh!u
2�n����TW�y֥�}b���)���oR���vT~1�Q{�!�}ɽ�pK`&��.��EI<L+�O+���P��q:��W�J���mm��c#�i�;�CG��*ej�Pa8u��Y�F�!���\����w.�wb��_&D�rwxgx�c�og�%09Ɯ����3����H}��{xts��9��u� �[=<_��xm�V�܈t��.��yK��k�4n�PP��kw�1��զ��bӥ��n���:��>�G��1T)�5�ࢷ9FI(5`���,Y�m.�B�5��&�∢�C��DYgſY^�E� �Ι�ǷK���%Fv�^	O���8���j��������j��e\K�6�Y�f�\ݞbe���e.6¬��*��G);Z)F#��9�%\6�h_�r:#Bү,��Qժs��ᨑ�bfdإ�PǼ�]��X�JX����=���W��)�8Dǡ 3:��)d�v��w��5��`z���#v-�(��#
�S%ao^�ګ0c�w��z���=e7��5�R���T�C�:��kK�'���;Л��"*DErOV�����-լ�.�V��`^*����}H��5P�� ��+��e�FFb��#é"ݜ�c�>�Kwyə�� ���v��Qr������a���v�\]�F����n���op��������r��r�7��1�����OMC��l*��%$�m����dƮޚ�ZPخkw^�{[^���io���H~O���8��y��6�l�] ��l�zNQ�	�I�+�ݲ�O�cT��3y9��M����i4s��ִƬ�[��ZK"�W���#�s��4�s+/3�������汸���ڭ+n�w�x;�`��Ó�S�)%�.��V��/^}ضVA��'����RwInd�2�T�����W�N��X���a��\&q#�4���7Om��8^�z�xV
[O��/A�����h��T*�%-��7�-�w Qq:.U�����t��I���FD�ln�]�6��&ԓ*^�"����9e��yޛ�vtʧR�m-b�-1k�N�1"�J�"�/r>f>��L/Ǟ�HﳝԶ?-�^���j�&�}q�{�p�;��lc��V�:����C��ع�\*�\.^�-�P���*�2������=�1g��w'��4v{NH��e.���{������f�_LΚGx������yj�j��ۀ����ў|Sp��W�X��]i�#g`���v���'nJ[ӝ��ZfR��I�/-[��`�p�ӎR��#t�{2��۱"B��(��,��v��W�|4zX�����=$�i�%M�=P֡�����
�hOZ�m1�8����G���`��ⱒ��Qܾ�&��	��x���:��'p�r�M�jc���۹#gX?*��Nѧ�T�]�w$�)�Uy��`�$�OoR�/wX��ڕI�)6�$@y��|%�W&tK� !"mY������\��V�U#�>5p��{����\[Ձ��5��lv���F�B�k@�we���k��U@e���QO㵽3�bW�N��n�����A���ܦ�Q �od̎�m�eZ�����[�=U!� ÞG�yI� r�a�e�o����RrpSN���Q$#*,��Py���y%TJ�J=���XZ	�7�0���1+�W8%z�xF�W7y�)qa�r�l���4��N��Z}cpB�SN�U��U���ҩؽ4�4�RU/7{;;�fm�z�=ah�Ht�BŌC:��Q�iN�n,�0���a�͹�)���6�W��կ]У����߆�o\�;�t�[�^��;u��n?}Xj����;���b�}�Co1�Kv�.͆BR�-&�z�'/�^r�Tv]_,�ڰi��u��VkG]�R�$�x׀�g��Nw
�Uk	�Z�La��b��м3�ډ���\��!�6�*R̄�t�K˸���gc�M��0�E�KC�����a�2u��l���تPw$�z�d{�h\���8钜�����#��KOs�����~�Ֆ�#
?}�zf�<6�n���È|$|i���*�B���ћvlI�VU�컷�o�v�\S4�N��usnᨅư�'��+m��V.�"9�,�R��J���ö�0Rд��nǹ�ٚ�fio�F�k�ӶNt]\�@��X0əy���&�]<\�1���ΝD�eb�˅�'�s��%#_��Z�y�%P|�{��#�,b�%�ǣWotWs(0FO��6]��)�y�u���OsI�J�H�C��� �Q
���6�p�����,07���Q�7R�n�հ����y��Y�x���Wfw#]��Ǘ�����邂*w�WakPKOk�;}V��i�k<�Ɣ^3�՗����Įۂ�w �5�>#	�Ȳ�N��+��`�@@ٮO�I��hV�x��c'70���������lZ6eĢZ�I{���4.�yw3�V;�]2�ˊMx�b]In�jjN��"�a��
���^�������F}�N==,����fL�u��0i�H���)���?�b�c�ܭ���%��^�d.k���L��aFxfk9I���;�gozt͝K1�L�[�FM7lm0��+�c��kS������sF@��u-��5e�>���G����TX6FЯ,z��(�YwK�:��u`+�;��[��X�*��%[ivR�5���_c��+l�|q"1cM(��J�ޔM�A]��VNQ���|��H�}��i�m� �{���\���k)����Թh�5Q�[���F33�w7*�������R⥌fWv��&�7�Tޛ�:�Gf�Xj[�_����&�1T�O�� �a4T��Xf�Oj᥆�1��7�)\��a��lr۝�ƥ�a�'2w���I68+[ӅnZ
�^<B���7[��<�g�ȗU�����*]������y�;eS���:��:�sc�����۾(O��LR����.�i��k�t�gn��+��9W�f)c�0�܉�L� ÷2˖�t�Uq+�.�S�/6���[���Q`��:�+'�ъ����X�#֙��O�JG�r�)"ɛ��OH�^�h��?Q��~S7����������c{ 5��^�b4�U,��F�*�)�2�~$栰�׻%�p)��uf��]F)6pkYU}C	܅�j�fۖEÊ�Gkd�i,�Ӓt�n�[���t�>�WG��q�Wم�y��XL,����%���b��Y�ܻ�ٝ��}㝥�qcWkd.�`����Qp}f�n�4)=�s���e��om��_oEJ����9�9��қ.���}�$�5)�n�w�Զ��:͗��h��1^�;a���s�P³r�}�G��ʎ7��2�t�RZ�::RD�\�����j�I���]������l_\�T���c�o� |U~��q^������S<�����\ts3G�s�ݚ��hd5*K͡��wXm�0n��w�Y�;�=Ԗѝ3���q|���G;&�))�kuYX2�l��T
�g#k�	�ueF���9�i�u�T�y�6�D�L���������N�nRlR��*�:e4xm���<�U�ϙq|{�61�<�ɺ_i[����Z�2{�Z��4�oA$9����ڴ0���B 
23���Ē�lv��
�'4�d���gq�k&y-f���n�P��!J�c{��<vD�Y�^�x[n�*�4K4a���;04�x��� �@o\�$��ۻ���X�i0�z��;�M�f��s��qS��J5Ֆڴ��.��<��p��.��n���5U����|�D`Ԍ�j��g5��v�[Y,�k��c�V4
�sL���o��W��M�]��Wm�H�n3�6OA������҆�95&S
��}wv9mrc���ءX��j7�v�����F�ZM@��9�Y�Uw:�U٫V \�*G�o9M�y.F>0�.�N�m�2��ҢgI\:����Ea����FX�RwE
�� "l·(���W�A����ZH�h�m�n�q�W���[��m,����C��Ok2�lkS����[�a�����O��j	ʯ�W�ܩ�ku�X@��bˍ1�*�yv8V��1c�,*LN4*��B�<=���E0�!&�G��"��1I�Ta������f2f�
wwı"�f��Gi��FgE&>�Z��%�&�^ z��}���ܠ٭�����u�6��c�D��r���uʱH	˶�zӎ�l�����ȱFK���UcP�g������/Pz�PrQ�;��n��@%wk>��o^t;pՕV�㡸ЖZ;kL]��G�^�ڤk�bC-��-c�ST^�Rp�{����\��j��l���[[�>|՘��F�����r-I)Yq顃��-L��H���L���p�SYM!�Y5t�^��X�k7`/U�v/��Z�:͔6�+��,cR��������֠������Z��s��O�x4��K��W)��7hl[�Σ 1MQff��f�wI�^qZ�7�*Pn����}�B�y ���f=S/h�=�+�g��v�+�x������T�Dt9���y$]�b�������<�5wC`����{L�3s�Ȍ:�Q��5W�HP�MԮ�����I�Dz�4��xa��ƙ�fk�/xU��Р[q�2ë���g�n�Q�W����Hh����ƣ��m�9�\���>��ᷲ�[���'f��w7�� �a�e�f�]��\�	sQkxPv�Q�r�^���:�E�ܻ��ﾛh����̰^��Y�
�2B�k��#-�_N�%#WtM%b�1Ph���s�zy�>L��ш��9�'���V1 �ys���G� �g)�R���m`�u�*�jĕz���o�� �L�ukm�J��jwt�$�r�c�d���W2���x��8�4�<�Jy�T:�ۯ2c�i[܍�$�z퇘��#0<�:x��W������if��lKQ���L�����*8��ʷ+�	7�Jk����[W,�B�!2ucx>!�����.Z��ٗ�>f������H2W���ڻ;rw��N�F����Zv����t9��|e������ARO������!s��5�XYت�u�!���z)��c,g��ϲ#^�wϵu�_!.��gw��+���{�$��.:������C�~Ջx1��ז��4��o0����9���j�f ����I�2mJ��Q\��p�]�� �����de�5v���s$T�U�
��Yk�ĝ���1��]o���@���d�'�K�zV�7�dڱZ���6�sάoM霶��o���%i�TcotIrPVW5���6��t��	�� �t�:5�l!�R-���;8�X��8�L�Ǹa�V�%O0�I���ڊV����`�a��C	=7E�G�ܷ{�h�5�ê��Ę�[3��{�� ID�{n���l�_��w�]7ܫ�K2�2�b�)s�rZ�ǥ��w��:�K�ɚ5��E;����'X�0�e(�X����;S�k#ަ��{hf]��b�Gd��W.G6�Ǐ���#}r��s}@ٵS�b��G��M�j��̬���*��Yl��^�����{|v����v���8�{zB�Ëh#jk��&*��y6m�[,���u*l"<�&Q:(��nv���x�ӗ��![y�=���E��)����4M�%{V8���:!����8�'��sv��`Ņ�s:��҉���(K\Nw�}˰��{�0�W9�l�����Bu1� �r��ي��*Ϸ�Pu�ŏݞ���S7L��itM�lҺ�b�|�Lzq].��Z�������@�f5��0ekc�^�~;Fʤg�q�<��h��C銁�G���P��~������r����2�� 6���csv���pף}�x9vЦ"K���=Fg������F{�u����Ὠ�\_K��t�e��
�ٻ�c�t^�0f��<`=%���Ѽ������ �SK�����:������q����b5�.�.[d�E�H٭����3NU�ժ;�_-��k!ǜ� ._5�:�b���ݜ�sp�u)xyb���^P�ȅ\WWh�[q�>�W�M�=��~��q��~�C�1T��������Z5��b1b¡U��*��[k
��m��Tb�`T*��U�*(���R�E��e�+*�R�ň�"��X�%Kj*�dPY`���E��P��e(�LDET@XbQ�Pm�("��QA��m*�D��Z�b��Ȫ*4l���AVbKl+�V�*�,,�
ֵ�b���ۉ+-KB�b��h�QjV��"�b%�RULLq"�eET*�J��0���.0QL��DP���Q�ыQX�IX*�U�fC
�kV�dJȱ`��Em%Zж �`�,l1�ŵ���
�TY�h"���5�a��０귮�7z-�x�)��w�-tFR��iP]>޲�6�Q[���O�xګ�:답�u�}����Ӈ���|�15��?��Ϸj�k�ޓն�$3Oh*�D~t�W��i�Ż�᳖���ij�'D0���O��_A����TlR��:�Q�X٦	x��7k18��K�櫗_��������ttT�e{��b2Q(��d�d��v�^������'�d1F��.������+��a�]��r1I�ɛ>���Lí��܉ln����ɤ���&42��'�s�b0�����{Cv:ެqp��7�t�z����E7�w;C����E	C���b$8v6���u�T'� ���Zk�x�����l|X�Gc�|W"D��2:�"q�y�uOqu�d��=61B����'o��޵��qE�b�K��Eg���,7��~����^�⬽]d~f�:��=�ҦOZ�ݦGn��ls�79�4'CC/�#��;=K5,���~�u�W=�u���j�טk�sv��;�e+y7���j���0szZ� N�:���Y� 
<ɜF�H�z��B�VOM,�e.
Vw�O�>����J�=�^\5���ۧQ-��9�9��W����?�4i���̴�=I�K��޺Е�x����.x{_��6��ӽ<
�Uh|U�n���
]dރ��%�˩?���Ұ����-<U;�F�Ｘ:�� M�)�ֈ�٠�6i�f���u\�/�=J�7��y
�8�UwCx浕�w���_����ş�˚�hI��{\g������5��[¶��`�8�=�(t�v|�H�gNRzBYAoh�e���E���R���t�u�8�kV���1f���Gn5��ֳ?qƎ�Q�>C\��v� xv�c3oyy�DC��_w_�����ג�7D�=���6:�_������qB�I�f�laA��E��@"�2�|*�U�$�����{�)���[Yc=��4o"f4d�#�������:��yГ8@�k�Ѻ� ��U�IY3I�aዒ@�Kr�]&4ӪP^��i�p็���v��M�+���D��lW�8�üŲf��@iPŬy��i�u�R����B�;��/�W$�^	鷪�E��E��9�]c�$�@���@�Y�,S'q?c�r�����`�BD �4��wf�����w��Owvj�ż)\��n��jG���+%c��zL�50���]�nIT��^Iێɔ��sӝR�����ݾ��� A��	��y7��랡���򭦕��&��d:#w[S���b	W<�ʝw�n���w�k9�є`��?	u�cu�9����a�**��(H@��c�s�a.Y�{�����3����}R���<Mㅾ�@�q�������u��E�UL%���uhjv��K��>6Y�3<��q�ݶkP�LԒ�.�ܘoCC���XA1�3j�.�ەݜ�y˺\&D)�W��*4D��{/�@������罞 e1y�����b�z����tާ�v�ڗĬ�Z.3�>��
�S����WQoy!C�˝}��c�H���R�!]:Y9�n����4X_{<5�]!Lg���^�t�<o;��:�������fx\�yw�>q�7���tA�9�f^1�Β�Ϩ;`��M�����䳜Òk�H�S����֟�D�d^���:b��	��shm�����I��C�gcQ�jW^@�Tb��<��S��V��CE+��C��m�ΌWI�J�L%:#S.�Y(������U���"����,vm���N�=\���&��g=+��VK�����.�T�i�L�z�IlL��o苬vN��L�KVs�#��������xzϹ���]/{p�p���YKd��U�)M���U�Ɔ��M�Yإ��"7���8���}"�hўV��.4���9's$s� j,��m�h1^g>M���^�����<o�u
�d��YtYw�����s9�I\��ҞyFK]�5HĶ���z~�ORzQ\�VA�*s�;���d0���*�e�P�_�Е)�А��"�axV�ҁ�SzK(i���.����N76��{�4�����͙q�Pq�+���xhV��1N�:�H��11�{Ul����A�ϳ�H�kzE�w���]�R�A�_��C`�]��Sd�O���"p��ݢ���y
	q�B&S�_J��Q��."27���r���cm��kk����j�Ų��u��9�>�4��,��{xЖ��#����(�W�;�Nݢ���Q1�`���`UZ���Z�|�ѯ��q�������g1,�n����wy����==~$�B�Լ�oW��?��vi����Oyq��~�F�#��R9^x�`��g֬�ö]�)_!wJ&�v��g�:XX�� ���fk��Ϋ.�ß8K��B���{�8R�'�Ǯ	DhIjg,��;���Uɥ��{�ɴ��nC�@�s٫3��l�Zg��}m\O�bU��
�}�W@7�en��{0v-(����黒	ӸE��ζ��[Œ�C� ��R�v��:�Z-\�Z�ґH��ì��W�2�]���v�bg
�~�Q;���X�BˇiR����st�:Fӹ��7�Z
ؑ�XB�E_P��_^�clxȇb�ή�}�!���JN����d��MY9�X'��C��+��;#}�ّ�Ӵ�E;�r�˪5c��cG�⤛�>��O=C�y兿K�eK��(�{<<�h4<��o4S�F�{)3[П$�efK��ہ��}����,+��2�Q,R�^g�A��wn��vB�d��֚݇�<v傁����os��^w���(�¹Q14 �����M^��Kf�
���zT+����;�.;D�	�a�T4eN�Ģ�$�f��j2�R�y��纳r F���fs�U�Z[��S���0t3r���	�U�[�:2-�Ol�;�6d'<��{�c�����dB�ψ;[��yv,��Y��fk�����ٵ��G�������r�D>T�@8�@��m3�:�N�ۑ�=y��s�3�w�"��/)��%��������Jv����S�4tө{6�v��Y�5p޶b���处ٍeGY/q<���`��m��⾄����c��KS慵I�>��ma�Qd�Q���`*�6���*I�)�>Z�=����Ԥ� �-Sw$e9��!��:��,�q�y%�G_$J��B�-���X�2K�$Yϸ��^�s6*��噖�scT��Fń�����e���W�(�gr���mg��0�w�O�vGԽ2�gѼ�U'3	�Bj,vy�@؋.��!�h�P�=���>�ԗf�;��W,���6��΅�J�M��� 7LE���)Z�Zt\^������0O��d�� dWi���>ŧ���B��ק�?`{��;�.�ԗy[�7�fOU��(���!A�8��JJ��6;r��뿌���O��3�ʕt���s{2��'5���y�_�,N+���)�h�$~���">O�dҋ�u'��[���0��5�"�s1���LX�⼩y��y�ֹ���/���T��OH�h��\�gDdFqx\�'DC`��2�w_��yU��ג�F�=f�l.v�����K�v_�N�Ff�؟-B�a9QD7m�
n�����V=�� �R\N����h��Qj�B�^&�%Jޗj�^E�9���
��:��UK��G�ñx�&:ߝ;����yӑN��O-8�p��4h�-�Y(,�"Is&H+@W�TL�3b�KK�+��q�,t9�"U��!mEN��S��F�)M���'bC�7��ŲM�"K��=��l�)-��.2X.��G׳��5;�tSj�7��7[OYp�ەuS��n�eei��ӄi�Q$��1���|w�._�{j����=�[�)TD��E��X*��h�3ħ=�g����/R��?�	�庳�L�4��*��&*�Wv�A�-$�U�o�fwP^S�(3\��W��u�̒DhFJ�+9eŖcw;��^�}����B�~}֠b�iNˮ��<�n�v�=R싋ĕDL�)gly�C����׺�&����گ�a}k����p��`8s6e���'5�Au��B�}�s��=���Ỻ�����,�!���I��G9������@��X�a��q"a���iKX����˱�㚁(��(9��|��f��ｗ�C$uJ�oW�94EqZʞSʱE綸ze�������;_���>�W��Hc�%x�E�L����s�VN��vG����B���3�>lV.+hg1@�w��Y�Y� &�g;Cø�Q�ŋ��5c6zf��/=E�Zw�_������@�^c�|��Dfm,�n�U���[]��t�9����	���}ę#12�����]�p��O�x
�N04V㒲�1��e��]�.3�:Z��.M��h��۫yI��y����J���~]�zMK�JX��R�b\A�vY��r���㴧b��ݼ6�cَ$:�S���;ꬶ+j���&X�ӄh��ȼ;�Sҳ��㘾��{�9�������~�&���􌯛�X��[�lc��JE}���Ut=���{���]��[|�;�g �=�G0Pʢߐ뮪"��{o�*^�1Cc��}\��"|���(�e�v{7y߽0��$ʣ�-�B:D�A6"2�v���Ì��ҡ���%7��1p��5�(#Ϡ�!ꆑ/%�M����BU'��i��W�������d�5�a�k���ʡȷ�%M���<>=+��^���b�zK(i�c�굻x�P]nJ�I]A�Vt�{�2�t�	�����ث	�b�N��#�&GU.9=����쪕�C1+�����^����C��{N_���f��9#mj��%�6�h׋�GNPw L<`"{~{��}�=�}��D�'a}��[��Jm�ά�eշ�J�Y��z#2��z��^���ٻ:�R����,{_IF��o����a��H���-h83�u��nbr�ʴ��&��3��ׂ�W<���ܜ��Q�V���99�wY�M�>��G���Qy.�p��jg[�#X֏�.���}Ya�V�	X��U�1
��N��Ƅ�5q$����*���s.�d�M��_fD��'p��BuP�"W��jej��:4���A���P�X��eU'Ӎf�J�X�M��w�5�s�N�,gǵ/!�����g��m��aҿ�&�g���t��Q�B�}�~"^�]�����!wJ&�v��g�:_��uo�㋴�����y>�W̰�
㪶�L�ZLU��;P��+���D�s��Yq,��LUWoI1{�_
�.�SS�H�k"wh>�xaF�wc��˭�:�q�Q��i���W�=���a��@; ��4�#uU�b��F���{]�X�i�raə�S��.�{�*�$���^4�|��������?��3>
єJ�ER�>�6�Z�pN�q5��-�)"b!��L�PQӁ�K}����h����/�ސ��SEݾP���בr��{��ܚ�cX6"�ה�7��X|��;��^�EE�Q^���y�1�������%w���U��iY�À�j���2i��K��o���i=�N������~�hВ"��Ø�T�6W����Juc�ER
�Z���� �%^��b|us(��I��޵I��dh�ha{71��]�����2M��r�܊���ċ՗da����Y���_xgQ��<��W�	t�UGe��X�@�ɾޭ]A��*{5${䰖Vr��c�o��,�B�Nvu�ɛ�6#�y1}��s����.t�y0���E��/�0 ��}���b��b3�;-q'����}*��P�͗/i�N.T"��`�8��C�`O^{k�V����;G)�i(��/�k����llX��/�{����"D�����$NX]���|��z熭�9!�
����ۦf^�69N�l_���;઺���Vu��lyW.�k�;�p�|hz�걛)�Bn�f��9#`N|N��_6G��vz��̷��/S�p���ʰxh�ug���^�2��x���*3�������lU������W���R�?Z��'Y�;,�?	�U�3�����k�˄�X�@�T⎡orf�-�K;S���e,�.���J+�m|W��8�"RWB�o���y�}�P��)o���u����)E.��4%���Յ�n=���h��o�����_S�X)���7�,��CQ��hS'x��.��t�90�|o���)���(�b1u�җ/l�Gu�4��-=6���wB��j�J��w^����!OyO	��0>}�%,9{:�J�P��c�f�p��4��L����B�s�ӎn����OV�D%�⋘��v=j�0z{��)����{Ir�\tz�f������3'n����oMqdE��2���{%�D��H�G��W};s0��S��n�=|2��N�A�]i��E9��C\���ۭ��4�*�E�[�O��3�S�>nE�#A���n�HD��n�A�Y�WOKg�Wp�k)v�Kp�,c7W�8�D���Xڊ9س.�fs�[y}�'V ��*�er��'�<�=W����8ؐ�V�5���|��<�?�����e�c���Okr��˂,��,�%k��g���+%�x�:�cRX���=�$��wĪO^v������ ��v��y�t*	D�qN�=MYt�;�����a7 �yy0� �����?^�K��u� ����w:qA��f��	�=q���A��4n>~/���st��d7c1�tBu�*V\j<8e�Y+��}�fq����U�MY}%\N��P����+��.�V#����iPA�t��:���ƅ�տ\&�R��LѠ�<#n�J�P�U�j {#I���G�TLQS������uܥ��p<�,U:�}�Kau��F��R�$��Kѯ;152��W�H��8C�(��s��8��P�<sT����;;]@��Q>g_!���w��6<g��Pd>�~�%��:�*�f�j�"��j��ќ��!Z�*��U��ږ��T3C����.�AGڼ��Yx^',�m�����1P��k��;�`v=��j��)�b���]׏����	"�2�{�t���a�@����D��Y�U>�ҧc�/dN�]�@��ج��÷Q/Z�W �����3�/V�Q>���q���u� S�ˑoIt��3����I����jҝs49v�&r�|6QL�I�S�y�]��x/B��l�;rfcL�S&�}�n���젭�%�з��|𭤈ȫHۭ��9�y�������~�֪�����6�Q8N��9��1����c�h�=�7͙�C�x,)V������t(L�GZ���Xl��L7�37l���[v�܆g"�8�G�ak���Q��aW	�0�(-�(�g[��������Ug) ���B��1�k$�v�:�	���+\$��.�Ѥu�t��T���)ښ��U�x��P7;skK�N3�B�2Ӷ�A�͌(OX�â`�g�2����Bݹ2�&#��4|&�9�%�[b��AEV�*"���E�G��V(�������J�V�[aVڶ��J�E�bԊ��F���+jڰ��)m��PD�Vڊ�Z���[E+(���Kej����(�--eB�6����VҲ��iB�iZR�m��*,KJ�B�[-"��D**U�J�%�ERԨ��Zօ"5� �E�[�mU�(��YP�2�,Q����aPX�PU-�m��(TTAV԰R�QF%�-b-��ҡb[T[eE�[J��R*,�E"��KJVֈ��գkb�#(�5����EUV�DQ�EF�R��,�EkQ`��ڕ%Kh*5�Z�,DQE����jQEU��Em��(������VD�T���%��������:忮,�@|�N1�U��V4M��zybX�\���g)ǽ�k���o}&�,z�4.���)<�yM���e��P�'�/���G}��ks�����t�ڝ�fĺ�YC��Is&�e����ZnZԒ��k3pv�ua�B�q�u��7�~-���`���*��ι�|��R����M,�R0��ꗎ}�а�DW�̩�
�C�ͼ��t�og@�d�\��T�����\��*3eC�Q �O��\�NTV7m̷J�����sq��l���ed
��k�Lcr�-�6�U�)q��]�0�x���AD����Y�֤��������b� �1�P�M�5�.������b�U8/qg�i�p��1T���\=�k�L��~�r��JY�>e�@Nܾ>��R��B�KX/�y��m8����7�v�+�cՔ9e��`H��3>WzPg��滹�HU����cC�9��717;�-�RU�6�uLߵ+03�S��D��
3��eO/*�^Ȑ�P��*�@=���Y��z{V���B��L��(]i�0o��9��KwCy:�r�1�c�^[��.�V�nV{���B6/�*"����,��ޜm-�T��~[{kq�^��ˮ_��U�j�y�PǇ��ƨ����M�t�-��f;b�nSu��L}эx�@\�vVf�ܬ�s��$��vJ+D�{�mXm6!�{:��.jF�B�>�m���.�Zag���!��۶�}�g&hI+��*��}P�5��B�7��xz���ҟ>�b���0�Eu�@�WG�}�ФP�v7�G�M�.m(������M
.�JHx�d�&�P'��7@��~K(�;�|Xʳ��U�
�;���ѕǥ�p9�y+�_�4��/1RM�"�u�o��1�4,,t���a��.��
��<��[2�յ֮��=�(aI�ݺ��v+��?\������e�c����pC�R�]���G�՞Ð�L��Ľ����3i�"�|�.����Ǉ�G�y�E������\Y�-��g���A�5���8O�G��e��R�juʌ��ΰ����}��n��=��H��VE��%P-����������ʇP�ш����c���>z�R�|�D֘��r�`�&�\�P$ �5RlJi�+���׏O�y�5b�HH�7W5�A��j!����ֺ_�lI����Ў���{P��b=7�����n�C�Gxǰ]l;��T������nm��v�µAA���n�{�Vϛ8"^�4��E���E�aPg�E�{�Fܾ���Ue��6ʉ�hg�{.=u4�dwM<X]�5���$��Z�Dc��c'Wl[�\�KF+���[S�r=3�=��H��*�9�9�%M������1[�-�ef]��omGӥ����t�s����b����8�P8&Y��^�]�!:�3�xBS{��2�����M��Lk �b4
�Mv~�׽xlG*I�P�@��7�dtn쫣gsw����v��J[D(�yJ01o��l��s����N+�[�[�N+et��`���߹�S:R[�`�1q�R��x����5�-�����%_7��*��v�^�͇n�LlX	݇��u�S+Q�͇�\j��8����Dq83�S�;X�A������Ne�P\���E��/����Xߝ��:n.�r�$���k�ZC��܌'u�Oѝ�6/Ml��#�b�y�B��_3sӂ<�ő�����=og[�	��4����h8糨ð;s6q�̌������C��;6�<�F�^Y�b�-"�����r���E�z�íǆhWv:1*��{9�ہ���]w1���w�^uկ�8�z�t��W)�é%G��H�b!a͎���W-��Ju���T��S�pޏՂ���k���ݴ��x��η��e�>K1����l��o�*9��r��a��,���嵝W,�|�|��g]��n��t�����.:����C@�"7U^L�$s�Ib��P��A�WU�Os] ^$�t��ɪ������/y���I��B� �>>/�0ɔ���}�3d��P�K�6\�PQbQ�[G=�W\��f���[��K��j�{�;ɋ���.#tV:�9�;ck���72�Ϡ�ޗ޹Se96y:��[���k�ǌWxr�!DI afWޝ|}�u\s����X�ǉ��~C�n�t��!J%���$XK	u|䜺����X�r��o�v`�R�4�7�i����K�m�hد}�� �����A1����O-��k9������ulJ��6��T��%b�<�̞T5���4l�����ʇ"`�|���Hp��
�Q�1ت3w��5{�C5�~(�s�]q�FG���G�����0G��D�<𺭙�L���
�o�K��EUͰD���a`*Ën�K�9PȬ�!�S����7��YG�'3�bbI>�â��s�H����a���N������*Sbv��us;w�|��}��d���G��/��.5�ɩ��}�,�/nx�?l��i�c�e������%������^`�Y��%�z<*Xv�t�tpm͍�)�h�uw0NR��TA���Iי��mk��ܷ7��Sv�469����X���Z�YDP}k�OV��\����a��t4`#����~eSwO�hZ������R|�10�k��xA�f�ͰxnK^@�`�g�e���v��g�i���#YO}�ÁB�Σ�4
�8��Ūt�c�C�J��	������k��F�^��h)+�7��u�[�fu�ѽm¾�.?]�-��~}�`��F��盅��bqgע��]hT�2�NF�=j����ճ1��l��N�5�"�lf�����ș,E�����\�	o��^�W��f�C<.���] ���^��	�x\�WFE���oF�]7�YL����b�����E$X8���.˲¬�<��y��DIӋX��Mڀ�Q�#����YӗmL�-����<V)jHj�"!��jq'�2 �g��p}yil����>x78"[�$�\Ϯ{4�Ҵ��p�k�Hj��B]&!��o���tCC}�+�4�&��u[�����վ ~O�o���h{�<Q1�e�sF��3-�\C�׎�φR�b�;suʅq�$l���=�0�7��"U^�����f��W���<ڏK�ԍ���[c[������4��D�5�h=f��V�WR�IJ[FD�}�dL>e�6����Ƀ�Q�TwGG�B�{�1����ѯ�EYJ��N^,N��A��ތ3���S��]��$��@f�C�J��뽜�k����({�bV��u���c�iL9�d��pkǂ�;Y�1N�Acq-�O΋��F�@�� @�{G�r�f-XQ�6u�<y�#���8ǀ����vu<e��ךzGx(3B6��Y+<Y�&y��{>��,��g���ܽR�JJ=�=˽u�6Z�8M���펳�^��Ԯ&D��бK�T_�S��N@[c{s�jn5����+nL(S4����؈�s1����˾_��>;<*��^�g�+c9���<PF�]���Vd:��IL�d�s͊��hVc(�CܷV��xQ~[�p�Η�P~�b����Wut!Ļ�|�~�.��@���&Һ���]�k	�2r�G苼p��U���8�k�w*�:�]�Ni�C�W-�����B�Z밐�6�\<E�A�i�R��PC2rܒ�:3-�T��{j_*����A������q��u�S��cZA�p�j{��E7��&�3�P&A꒔������}�-4��T{�.�:�f���A3{Y|���;��;�l�ɨ�C^K���
�Q~YQ�[`c��JE}���r��=���ޮ�����^m<0cyч��#||Ļ-�b���2{|\'>�ш����nN�<��L�+B��uG�������8a��ݷG}l:D�I��4��(@N����Yi�H�YkL�ظeq5�A��Ե�q��a�C�K��)?��=�L��Z�oe����ĺF�3�9�C�Zj��	������AE�%���^�%B��u�[� +BF�'�ܖ���HW�R�b���c�+��E���q�S��xN��c�%�ڍ����O��&Q��	�,�F��{]��8�z�؎������0�-��s�oS�-�I�zmm���TBL�܈#����$���&S�_J+������D"�[0cF*��I��g�$!�ٞ/[�!b?
q\T���\u��1
'<V�-�D��/1����B����1/\�C�:��ش�Á��]��R;Z�ӛ\j�����K��d�M��e�Yh�[F���g{��z�.��nm�%O�ن7D�J�Dx��^t�:�b�rx�+Zf���o2>R��7��*�ZM1F5���s����մŮ��%袥��Jʼ):�Vd���=o9A��瓆�Eמ����0V��f�M+���4D�\��g$js�MoCXl�/#[��=�_q׈$*]h�u�rՙ�.�:�}R���CcL�y�ܠ���s�r�Z��^xQ��}Y1o�NG6��x��׶U-���Z��4��n��̌\Ż�sjh����O�7����ik-@���¡�Մ+݂�$F|(À�p=˾�]��Z�9#)Z��]�I%�jҿ}��z����^�W] 隃�&U�bgy#f2��6ɭ)U���zK���NB��e��߹ko|c=͜�����h���Z2�B�F�v�B�@Sى*��mt���J��`O�\�+���O�k}�[�s�2�$�ɥ�x��k!k����R3f�p�f���紅b6|����:0J�ΧMM�Y�v�]������$֝��[����M���C�vafz�7��yq������I�|��:��nze`ػ�ֱ-V"�"��X+�Cb��r�]%��W)�Ɩ�9�C���j�ߌզ2��^�^e���ՐL�|�-@0���k�)�g~ǝ�~(��g׺h��;<�jI�'��C��T�ن?����ï�an����k�{�liEa�y�d�Lf��+�HN.��g�M�h�>�WH�K'K�kY�9c�������گƊ����'=����c㔵\D(&40P���Ȯ��ή�E���&�5�Nt=2�H\�ܕ��Ԏw�q�����.Uȃ%��R����㘗�u�k������II0��p+x��\eF�#cb��<�^�K��,�S*_�K�$�y�e�����[�1�a��1K�H��qP�(t\���↙a��ذ�޹�]q���̼�p�F	1���BUq�˦g�k��Fș�369�r�7�Н����iz�-�w���޶�2lW �y�R���@��jg����+�p�޽���y7���RN΂�疚�����]6��ܨ*�t���F	���&_ń*��l���Z`l���N{0��޽5�|RQ��!���
�����kDE�A�.�3�X���Y�˯2�TD�5U��Zk+-VP���c�<�]�g[�����zHƻ}�����4�z硩�:+5�ͧ�ü�_�=�����2Z�����N�6k�E�꡶������[��{|��F;�w�2�� d0�1,ޘ�Go5+g��W�/�p�����:��r&e3I�9hxm�]���{���	��;��X���=�SBM�R�b9%��w6�,�[60���˱�+yfL��P����)mb��C���EfB<(��8�U�R��� }x��|���F|#��˭�9L�^Pvk
��^�󎈆�o1����v�' I�z�o7���b��c'ep#MX)�������$m�����	:qk��'�Gb܎k�ͥn������g,�}ψx�����&�-�|��N"dܗDP��?�=��N�2n�e֫)��T�7ӏ�7MZ���i����4Њ$�����,Rb�$��̬���y8���^����,�1}�Av�0�]�||;Kԥ���C>-��(��f�����Rv�aI9�.�(�i`�X�lh*��=�OK�A������u�$�^f����*f>*�Y�)�	���nTC3�рC�R#��O-�y�Ǻ�ñ�.�z���-e���q�&=�o\��Ͼ� O`�#����WপXQ�:���G��+eЅ��˙W��,�4��6�n�dCÞ
�Ѵd��'<Y����^��ޓ�<�5.�dY�C�ZJ�����(Ā�j,n��ȝ
�����BÙA�g+�VD�����L�t�f��1cס���.#y�oe���&6���K�Qh�w��	O���]_sx�aof[w']	�v�@5���y�̘]ˎ���K�R�F)�f�ɇ��b��lwA�V�rKu�:�%�wδ5�>�,�ɝ�'��6�B���{�U�vy>@����e�s�8x-�Q8�LK/����ɪeʽ{�dh�DΦ�=��B:���Ɗ�ĔhZ�#�'c��ᓷ�^�r�k��'yd�H�#�x('�a|s�N9Nv���0��2�2g�c\��|�F��q�n�W���ݴ0YZVM���)Lqf�z�$d����Yհ\�|�}6��cn��s��T�u&�e.}m�e�,}�cb���Ә���7!�d|Q"t��*`xTI�D���#����3I�v�o&љ��V��Yy��LS��ޥ���WvW9�%����^��+�����u�������{���K�����kzxwW�V��ߓG|�we�������5�ڲy!��MTk�8u�bW���4ӽ�QM�+o	y�����-=8�`:r⯴;�!�Vz��)
�<����	eeb-�s�Ҵz��ym�X1��LӼ50���'3$D����c1����`t��IG�l�II��;2>��~�j�����Q�F��bo�܋��Uݨ�w���ͭ�� u�-��*��-�;�+��{�&����[ה�g+N��7R!Z4��82J[��B�z�}��v͑�c��N��P|�;�jCA��]/��U���nY�fp�.�1�O�s93I���(s��尖�}�P�l��ީ	�ɘ�J�#tLn���5�^ҋ�aC�� �Ό�Ӊ�"�݈rF&+�/w
*s�r�c�|�6H{�h)u�m��mV*��/Z&�(2lū/t˟�P]��]6�4��8��\%��M-�D�M'{�9��ޚ�c��&�� {gAĖ�U��f�uӤwu�����·kx@�x7&�N�㦀�\N�]>=�n���hXm%�aM���)9\���5�ͨqV���1|D���n��s�z/�n�EŮ����lև\D�d0f��n�rUD��	Y�O:af������8��y#Յ9�Zq��n��o��J}�v��1�nҩ8���O^�u.�<��}$Ϳ��M6�.<��z+�ڈXV!ՅR���S��X.<����ղ܂,���`|ڜ��{����,��u�R����֧������;�KE���;t"t.��q�Y����3��t�S��+�C��KZ�<�z5Pr����/[T��J1����޾܍��<��t�C�����t/�d��
jt[�g���H�R�����?kl�pt�����N���Ɖ��Np�������� IR��1'O��fd�rb�s�!��D�;-ћ���m�,�p@^e�Q��
��j�YbJ�hd"�[���}n��5���ś�mj*�5������[A�b�$Q�X�b1��[�
[
��D�D����*E� T�XV-EUb����ʕil�keB� ��V+�"�mP�QAH�e�"�
Um`VE���6¤XEb(���Q�*�6�T*#���5*���Z�jҥ+AVڪ,J4Pm(1�Q���֬Rڨ��4�b����*PETU��R��-h�6�����Z����X�mF,F4�U#��Z)R���b�0E�V�Ҡ(�X���hQPEڶ1��X�����cE��
�ъ�(֊��c-(�b����EV2�"ձ��b�QX"
��DX��iA�R�E���90�B9��d��oT+YU��Gir��uy�����>֔9ٝ��%�OM�����[��V�E��I
;m!�x{6��Y�ڼځq�$n�X�O$뺸��	���>�o_�{e!9|/������ϻ�z�f�=*�����yL]�=^b^�]�s:���S�@�^�wX��ttFm��{��R箒����@V�՗HSL�8�j��}�~�|�`{����%���1�qڄr��8�J�a��&�{_�_B��3� ]=���ё�SnK��:�
�7ڼ9^^��k1�M��P���P�/W��w��&7f�8�-юǥ"�S.��ۣP\m�����3/sk����<��ttb�}p�
���$[��`R��s�6�#�I��i����M%�f*bJ�.��t��v��9Q��l��]�
�Q�ʋ����������7����-����¸��Qlw��Re�jKp��/Hic���R�-\�S�Cf���z�����䊌2�9�0�c�J��i`z!�02��Z�^�t^V���1�E��K���,���a���\�����C���A�8.�-LȞ��,�U��ZOL�7.��'fn�8m=�%h�{���'�2�k�m�f��V|[����I��<4��i�f�~�E�e����saE|+szf����dxNEL�N5�!ok��;�۳cw��Օ��34MRī�K|$�kh���}˩�y��R3�U&f�1	XO	`���y��w�xlGr��=��W>���D�A���JH�`�0	[w𝢟+�A�'R"I���Q�g�S���yL�|�9[�zJ�x��~�˰�Wu��+�2?
q\T������_R����=U������ZR�4u��� �.��f%��x%�GƧU"�o�N�2�gU�u�T��ۭS���C=�\;;r���P�I�UKA�rF�>$�B�G$�ޯ��&�v�,v�K}c7T�9'��O/\c�z���-�Z:��
�߷p��_�+���
����Y�E�
�FjJb�o |Ə|v�ڃϮ��2��%���i1Kz��iT�V{�����u��߳���'��'�{�,��b�6GnUl����{^g�f��Fm;[�5�$�����>up���:8ߓ7�`�?�����!(U�b�Ky#�k=t�$����d��`z<z`L�NtS��-m�s}{����S�:#`1I�;��&~�j,��L�?��h�Yow]J˦P��B�bE�����v�^-o�yk��G�@��Vp4lP��x��w�ٿm[�L�u���R�7D���;�҅�B��(ѬS*mD[[�sa�i]�J���ޜ�4�SzGE�9�IU7w;GU]y����{�kwf���c2~��� 8����9�7a�	F��6���f�elI���8��e1Iq�r5=Ӧ�E��9�A3�4�T �y�x��)рГ7���%<tbT;��jlZ���f|�(�ק,�%6��A�7]�t��T��!����ovk���9����o;ǣF�x��1�ZlEE���
�2�����\+��`^�k ���/�'��p���
�r0ɀ�Pp�G\꿢 �I���I��Eb���x��Z�������FI�����[/���G+�/� ���9��W܈2PLFF^kA��1o���n�Q|41�~Ճ�,V�)�K�2�C���m�ˌvqx:R��q��}i��{�t}�<�mT&�����ꗌ����,l��_7ڻܘȯ�ʈ��D���ˉ���[h�Em�˖Lx���KȪ��Xlg��6F����9.^�.�ew���e�{��]��C�������=�W]׆5�ή_�M���0��y7.ṽ�DNgt���'`Xk#��Z�Y��M������4�z���讒��(F�Ҿ��s�����}����v�rř�ۙ+���͓Y��m��k)�ڌ��N���o��X��!Q�s��ז1�bU�3�p0�h�gOlY�'�о4w��§,�P����{�~����؛-d􀾗@u�����O���U�9xd��B�e�tM���'f�sj.�^;�mh�-F���4�U�D�q;�/Ԩ=�-��{�j������Ճӝtq����|�����.=6�������9�����|�\2[{�ɍ-N�=sp�AŊ�fv|�]=��7V!�c\r/ꡳ���)��#�w��<]{�&aN�1�<�ۓ��f���vk_V���f�N�es!m]>}�KYH���i��;2lB��K�����$o���/D�ii���p��)�vm��u��۴�˜�Y�U�|C�b���:����D4Ꙝ�Q	g,���p��'ҒPz+k�$)9�t���C�J�(����Q$��0vЗI�J��q/��9�W����ٱ���5�q�s�}B�2��Za�ۗ�ô�J_��#L`#�����h[Y���>���J����ƕ\��X'���b���FB�x^��>g��}OI�\��7�v�YG��x
	����8�}%�X�9G'��b��J����w%�An�M�~��Mڮm���|��[%���8C�iڴ�D":0�I+�9�W�[hJT�增S�w%Znsn��sE�W5��Ļ�y���㑻#}�� ��ɖKsȘ��~���"��Q�eD#6�fNҘs��n���x(]2)��htf<esUf��N�W*2Qd�F�1A�s��5W�D²�(Z�0mH�v/�o)�l��=6b[��.X���!��
Ѝ�%�J�h3·���n�3�t�� �eg:��-����N��q p-E��γ�^��Ԯ&D��Я���S��W0]���[��k���k"���8�IWJ<���\N����>�o_�{eY�qN6*�9橊�,Ȝw]��c}�ttq�럠+�ܱ��A���� b�q��$�wK&�s͊��k��U��xV�O$���Fl�.�KUѵ"�dp�.o۹��5,�{U1�{]ۊ�KS���b����]�db�F����M@�u��o�8|�X���=��jW-r7Bǃ<�c�r���UT+�!Fy0�V-	p��M٬N.Kw%�X0-n��s�ڜ2Z�C�������*�����A�קO�s��YF��%�-���<�'�Ɉ,m��ʹ�h�~�%�5��$F_ߺp���mI�z�q�S�g�ywd��G��;�wq������N�u��V.��m��H�ZM<9ã7
�����oi����*�U��Y��g���3}CK��b��H�5i]���LF��_&��xo��ϳﾗx�W&��'j �F�G�PM��t�V�?�p!������
5A������)�ns=�R�jh���>�=B�t�3ڃ���QtR�y�J]�5J�R�nR<Y����:��G�U�^�Ѯ�I�WJ��Q���r�s<��Qwa8j�m��3Gt���VTE(��\R[M�,4�#)��~��(�����W�qu�*qt����w�r�6K��gMږ5&f���Jļ%�"4W����;޼1T�a�O�S��N�0���S���Sˮ��|C����!�h�ˉvN?��_$�ń$.%X��7��\:"J�G�k^ �tϓ�VL��:�._L�Fߛ�q����S��T����q֯a��s�a'~��^��Jhv�;*��-#.��Ľs}����N�8V���v!	�½Y5k3�]�r�t���@���p4o9��Ȝ˜�	�ń�h�k�iy����5w�����y��ۛo���>BR8wì�Ǉi�����K̹���+�C7i���9�����,��@�+;	�B�O:L*�C	�-�=�$˧/���V2ҭ����*6'��#2�H���9e����/���y�W�3A�LKD���t~�4�2��+�;jd��o.E��WI�u���Iz�,��1��c�4�I]F��E|=�� R�ԩe�:�!Q�Gn����/̱p��p,�ۼ)3^G�9�U�@����I$X�z�lw�����P�ⱋ����
�{����TU�z��W(�p��;�4�Ѿ�_M��~7v:3�Pe��J���h�L�[]t������ř�����������ͥw��|���σ�v�˪��{�͜��wB����v��SwQ�w��2�&z�|�ʩh3le�Iy�[�F�&c�=͵��n��D]%���Dv����{���zG��g�v�u�M�*Pl�]��HV"�ל��ns���p���<s�k�j�(d�\E[��Iߡ��a��c_�ޙt�i��1
3�����.\r�퇛���v3b:�+���g���v+(�`�� �3�܇~U��,r��xt�E@���m5��T�Va�e����[�w�2RcC(BK\�YB�`H�i��y����
nف�������n�:ޫ�F��p�ӟ˕D
�%8!�p%*�}��5�;dgu�˷�.}�g\�ڴ�����u׷��P�o Ue��|�~F��.z�-����Ί��:̉S�vn{(�KUy1u��;�]u�6�>��뷓�������4�j]��$��NW>���\]7jM��T�����xx{��DYFY]\D|"FGZ^��
�%:%�Q�F�ņ���;9�4����]eC���I$K�J���]�����߲�ϑ��������=Ci�}̛bΰ�c'��&���f3�xw7��!�۬*= ����53�Aϭ��)R�վC����=�0�%~݁�LB��^r�-����Me8����c6�I�O���+�{�@�N3�!�)�4�PS�}��li+s4�0�cgSw׻�������s=�����{߷�o�E*���P�A}I�浩P|��>�O̬�옟$�Ă�*r[m'�*%x�����XI�Og�<�4�į�=��M��0=�z��f>���ڕ��{/�H��2x��^ϻ�I����s�M3���l�9�M�>�3i3��Z�R�S�}l�4�Y��b)6� �Ԙ�a�g���}����|G~̭���7�f��/<��,�����hJ�0���wg�L@�W�S�����Y�>��6����?wh)�Lv�5�Aed���y�/���l+�~��I:����ُ�
����L��!��$y�;��ޯ��_�k�|�w�{P��=a�c��~a�f3�g�m �a���6�H�q+=���l6���La����&Щ+����6�HT��w������g;a�5�&ٌ��O�i��d�9�>��}�|�w�ƭI#|]Eǀ���EGީ�0Pw���Lz��f��q�c<qR�E*y?o��~H/���m����c'YY�,�������s�d�ZN�R~�����z���y�<����{߷�>��1��&� ���1ĩ��8��8���C������x|d�c��wH)��ɉ�(�26���N?&��7����'ݡ��f�8�Nsϰ�W���{�����;}�˺�|�����xD{`}���5��@��p��|�������bL~M�q"�Ĭ���C5g�����xi�d�_����J�U��ZLAH�P���/��'/�|?�Ì�寛:�6��6P����h`q7Wjw��:��9\smܚquor��Î���2��������-�a�^e\�]��a^�L9h��q7�\y����{8��[�pf�p�|��@3�N�c��\��(��u��H�^;+w���x *jɢU�����\d��0����`I�u1�w�o���jb!�bC�;�N�X�L=LM W��3�~CI�����IR(K�Y0�u���vM!RW�����n������Oy�ṷ5�P=�� |��3�(��C�d�k�N3�ܤP:��&w�~`T�gK�ki>B�`T��Xz�>J�|��q�&0�տ&��"�s0:�!���>/v^���z�ߴup_�� ǜG�<>������Ͼ��)�%H/��~ѶN�N�Y��4׬��AO�}��%N2l���g̕�[߲OoX��?2bcğ��"2q����xw��OT��a���U%�s��#��L����Q�m ����$��1��vc�AN�w��|��� ���~���I�Vs!��u&?0�;�m ��c��d�EIYӹ����=��~��|������߼��S���2�����%B�d���̀��S��hq㴂ʆ����i�!�린*N'ɉ�)Ԛ~`T�ì�C���gri��X��=L�w�!����������lV�F��)Q/� l���;`��"���y���*c�Lw�"��I^r͒�i%B��Z�l���Xl��%���bx����P��fOY\`T�~�:�'�͏w����;��*�K��P&�X���0�w���������F��:�$;�z�f�uIY��&�1����R�~��%d���l��'����0��P�<�m��a�v����l�_���>����{�_�>Lt�����u�2bc�xw0�AH�����M�x���u����Ă��9����N�0��t��)��i��Oɉ,�z�H��L{�Ў���忺ki/����ȇs�H/Y�<���R(J��0�&�Y�LC�3��&e�M��6��T��wX��PR)�}�W�ʞ���'5M0�Wl
���.kψ�@6g�L��}T�|DU��6>���1��g�Y�n�H/~C/�m�!���?}�N��?%H���i�aS��p�r�q*%sS���~IP�l=�E�Y4�A~T;�*j����y��7��Հ�K��$�@�����f��>Ci�D��cS"7Շ� Ess ��B/yC���7�+�<�vs4�?���H����P�+	vԙNn�y��;ݗt ƃ�����l6�=*s����6�f������J�e�w���v���Ē�~�����ys�%@�\�|��tϙ*�̧�,=f�X�<g$�
���vi��Y�]�ag�:�͞y��x���/�bbOP���z�eA�%yܓi�N��Yώ���`���ֺ��e,���P ��3@\l	dդ�?r� �q��MeH�u*|���L�l��i񓩏�M�$��_P1"0ީ���A�  ��y>��xEF����}۽�w5}�=��oqN$���3�s$ӶAM����ԝL@{J���E'䯳�>3c�7%��i �g���4��"��f������Y14����&e��{I��B�a����_x����y��F��3Nd��UT}�ٙI'�$�]2i�'���v�!_�
����hz���/O{��>eCHz���ȳ��>f�<M$�?'��L�=C�鼇P�m*E3Z��ir��ş��b��{~`(���3h�B�����ĕ
���i"�N��|����w�O����z��9'��?v�봛B�����H,+X,�~¤q�ɝQ�+ΟZ��z>߱����l�!@�,14������c�E��6y�6����eO9��&�*T<�&5+'֓�N�A����'��5�"�ԩ�9�I���2Vs2q+�&�$��k{�]�o~�#>��ſ{ y@���Ͱ*
Df����Ă�S{��Y>~L@�n���$�(c����f��٤�8���<=��S�1�?���H.3�1�{�C�~H1�{~ͪ�@�W�ޢ�;&SG�u���
=R,�{jc<d�g�:r��Y�����P4��*V(U~`TnاRq㤃���&��>�4�?s0����ffӉ�u%|d���:ʇ��Q5�������&�RT�G��gO��C���]��s�h?3�:�0<;�i�!��R.�dSV8�ٔ�@�*�+�X������~���(�P8��}�Y�����Vn����8�O��s�m������yD��\'��=B���;�m��a���N�H,����?0��&$��$SHi:�!ԕ�TS�� T����q��*Tٔx��� @�*�F}�\n�d��U�oC�56�M.YלDr�f,k��.a�e���LpR��M/�2�2����P{��Y�e���`�H�F��3��a2/U&}�r��}e��NAu���%�n�b��:L����x��b{@��$�	+�����c�>��V�];[�2��G�ѭW\���`P��Ee`�a�V��� ��]ո!��4�}�_W[l�g>1�LV3Y`��R�n4�g�)}�~��s�؟Zȝ��\�z��&�,���WI���z+�p#��b�c������\8JZ&����`TD�KvK��_ȣ#?(���4��>�5�ѕ��H���9�.8��v���9�u"^���(�
P�c��L����Xv��\e�sq>���3��υ6��+ņb4�ʰ�2t��w(ʨ;N�x��)�R�n;�LÈ��F�ƣq�5�[�k}{�JgBLG�"F�́�Ǡr���i>K��hQ�2c��\��Zi�{S8�r�^��Ǎ�BIj�4�!Z%�v�����ySN����ŋn�� [�9�|��1+�/'�/z?yU����ČN���N"+)�s1�a�-����W݄�vo$���*ˌ�;�g.�E�s��2R.�i���&\l���e�G�!$ʻ���r0�ۉ
3�<:���W5���z{/3��sz�0�-��h�P�O;�CTzpyH�Փ0�Ci,Bn"tѨ)�W ^��eMA�<�-�[c{(��zdz�TBV��A��/�����*�.�2R�,dձ��3c�a��τw�\̧����q�A�co+�D�ow�]��yM��2��a &��5��U��t��ֳ3l7�I�i�%M�rvCz����x+v�M@ɱ�1h<n+���9qǯ�;�$�J=gU��}N�����L�)"9n�]����N�N��� ��f�/�]�9�IIv�����#����O�n;̧�9Pm�Q6�v�2+�8g���ź{���R��ҹQN���]gj����Ӽ�ǜ����e�������k�!ϟ��9�Z�������Q�����r�tl�7�[s��,ә�!�nˀ��4�4��M�Y�F��o��:z�s)_v9�.d��W"�Cf�{WX���;�I���n��Z&(t¦�:�L�(v�-��Q����cy�l��=R�96V��>$Y$�th=wJS}��$C\jͫs"��`%�"E�Z��]l��(�2�+S�w��*b]������Kcλ��^.���:�PYJ�~�ǵ&k�p���C����6����2ڗ�u��m�u�{�ƍ=8׼�����x7�������w���Y�:�|&Ec���E2��u$ѓ9�M��[�x#��1�6�X
�ԁQj̭Wu��	���Q�����[�~���ṴXnV���~	 K���X���
�%�AU�UU��b�����*-eUTmm�(Ե�(�+,B�Q(�[F%�-+QDE�1���%�EPUUX1��Qm�
�Q(��-�mD��1V"+[X�E�F�1Kj"Ƌl�cl����Th5��m���F���m�#m�Z�J�+Db����E�����U��F�T�6��Yj�e�����iQH���QQ�#����
���1VYiF6ʢ���c��"
�"��m�֖���,cPQH�
�F*��Pm+��m[(4IX�Qm*��PeF�F1TX��"�[b��EX��*R����V(�[e�EX�X"(�V��icZ(�Z"հiU[j  D|@\����9�e�j�)��U`�������*���s�X�ӸEt6CV�_[���6h��$�dͱ����j��� ��G3�oZR�@|�^;a��AH�z�9���'g*xwXOo̝Lz��fB��
�ɹ��������jO�$~�ך�ݓO~�v��$�)���xDLx	��N���ۛ��|Q\����4��wI��x�l�bA}g�7�����HbAz��$Ǭ�6w�M��K�u��h�gY?gwu�
��*ns�ԛW�
�����=�d\ 7�N��,����e|_}�|�\d��5�20���Y��8�&��J����>eC�6~�i�B�vy�a������!�m�C}y�^0�����;�@�V�O�̬�@�*3�^�k��������~�1�X��<�&�R/5d�~��R(K����J����}�'����n�I�uĞ�_Ǿd ����c?%H,�=��:��~f���sOY�q6�?h������-=����}���v�H���{�l�@�Y6}ϵ6��Ɉ�eRԬ�Zk(z����~����R,����u���%�����'S���&�q
��x�{`ltx	�" 3�rn��� ��RϿ~׺���}0d۴Ă��Ì��v��ǝ�4�@�5���¤�k���S�4����lgSb�?%H/Y�6[4���1�����LzɁ職#�Ƕ=��@w�{_��-|��~��>��@Ĭ��?~��*O��ލ�m_X����E:�箘x{܆��J��^w�?0��|`W���x���W�p�ɤVT<E<LH,�?Z��<LH/��+���:���׹�y߽�z��<C��&<a����2�|��a���_Y1�S��ᴛy�y5��AH�����{����}�u'��<d��{܇���&�_�xr��z�q'����{����~y�y��~��?���2�3�R=veR��=LI�+�"����۴��"ʏ����*��d�6ϻd�O5��m �J�y��N�R����Rq�"�k��/��G�������}�{���x�dی�ÿ������x�ĜB���a������P���Ɉ�Y�F�>~L|� u�?}G�4�Z��5���P��N���?$u:��>�y�o�fzͿ��hs���	���P�J*(h�w	�h]v?1�̭�N���U}a�Y��d��Ao-*��wS�yQ�a�,��%L���hm�J��і��Nⷖ��T5�ʓ����gL}�X��Y���l�԰4{'P�Y��򾯫�=շ����o/��`xD8��X�A���O'{�OYĘ�'�y�q+1��4[�&�:��'��kW�I����L�_�ެĊu':g�̒�L�����������}�_���}�;�=��y��v����%vL�Tu�w��q?$u��g�&09��x�3��'(�!��]e� z��E�:�ɈK��4�O9`c4�CR/ݡ�<�G��Ӹ��+*�)t��'�?z� z �����c<d������2�'�~�6��n��A��
��a����Yԩ�w�+Sl1�&!�r�ȥC�Ƴ�E?Kq����*�W]V�s.��s�
K��ly���ݚM$�Pٮ���8�H?��<d��"�̇���O\g���r@į��;�4~z��6�]{�6�x���s���ɏSl�edm��8�_�\l��z���+�r����̰��H-f��b
x�O�l�����'�7�ߴ�Rǚ�Rm�!�8gr}g�1�*sĬ�����&�6���jO߯XQ�A�Q��0�?o\�ު�D}� h�v{M �R���s,ed��Դ;�m��+����N'Ɉu����
�ϙS���M$q��i�:���N�Y4���c1�C���A}`�
���8�V/~�(��9�4z��`z �>�Y'��L@�<�HT�����b"��[Sh)�8�퓬�m���'�d���{�@�N3�!��a�6�PSg>��5c�^��������a돍������<2a��1;��=dR��w�*H/�?wZԨ>RT
���Ԟ2���b|�ԩ�[m'�*%x������8�N�x�?�d�@�X1�cT^v,�.m��皫�y�x	�~gN�6��c��&�#'&!���i�dm�}�5������5�&{C_�(AJ�O��g����'��٤�R��u&>0�g˞���+��]d�R���ýJ���qq6���0�%g�<���ɈJ�=��~�~`Vs�:���UtÓ�p6��N$�}�5�Aed���椾�������M$�bbf�f>0*>L����g��s������O��ƫ�ט����%ESo�OXs]�9�s���`�+���Uv�ګۼާR�SX&ӷR)�$n�[U�O9~�)^����^�?s���8�r<kъ�U�jO)X�����C\
9��<TX;��  ��-I��o� d��?��!�,񇉌?[���1���Y���Èf�����H�q+>La���&0��2u6�I_�d���M!PR.|w�nOS��?�@��>�G�=��Mm}���G�k�����2��v�z��=g\kP��A���g�Y1��0�cg� �2)S�������o3h<���5�:��yd�;� d���X�����s__f3�����m
����_Y6�ܦ x�1���<d�R�3�������c�&��4�
Dd��b}��F���'�Iě�xu���Ш3*��ؾ��u}����2~�� )�
�����Ag���{�~@�*��᧌�&;a��B���1�=-Ċ��.Y�& s��u�y~`WL8�%d���O3	��u�s����A�""�J[�"/��
��*K��O}��q�v�~���N�!�w	��
�ǟd�?!�bC�;�N�X�L=LO�����bjߐ�Ax���-4�J�@�]��i��}
=�kɸq��t�69q���àT������I�*
�i��u4��|�L퓌�~y;�"���Y75�jm���</9���
�S����`��7�gbcM[�i<"{�u}�#��d���?�R��_|��<H/��7C�)+��I�OYY�퇟����H.�����v�u
���k�O] ���p4��S���ߵ����q+�;���?=`T;�*=�P�{��s;�������W���_yؠ�FO_�̺H,����Xz�6�\Cr���N��2~ݘ�PS�]�_h�'S�Ag����? x���s!��u&?0�=;�?$�Lw�w�����d+��aM��ϻw������d�Y�&$���*i��f^�~��J�J�U�d"��Zx� ���f>�}�i��x~�k��|��<�I��A{��4��c<���ǌ1�8�0)%�G�{�up{v�~��~��0�g{�ڝC�At����A�?%H�~'3��aS2c�Y�*J�n�i%B��KA~������ľ�:�O��q>�fOY\`T�hIu��پf����V���ї_��H�矙��/_�����u�E�=^�g�sU�f,(x1}�c|�I{%p��Msz!���0��u��Y7U�Mkd�0����rW^qe�Ke��R-����D�,Q���BJ8���(�n����_�ԉ�)����f�����O�_^�?x <<Vf�Ͷ�C��ǉ=B�`]�jZ�gR���4�q1�����S�A~d�֍��uH>N�^�Y�4��g,4�d�Vs�~- T��x����HW���=��\De��tn���|=��Sh}�;f�*�y�_�:��Sa��u�2bc�x�&�ɩ�y��H,��;��O^�$o$������?��L
���i��O�P<"�B�8�f���Vac��w��<
�������c��~����!��p��P8��)�MnͲbs0>Jβf]$�l�N�R�zwzZ��5=��%|$T�}a��Nj�|	��|��9�͗���߀Q�{ j(xɴ%C�&��'P$���y	�����g�I�n{�N$�I���"��I>9`|�d��ے(�u��nT}����t	�Q��b�χ�%Ͻp.=;<�=K�O�v韙*S�a�1��X{5xλI��&������R�0�c>�y��x���/�bbOP�ܦ=H��ĕ{���gn��ע>�gi{$����P{�=1���ܘ�R������+&�'�ۤ���O;�`bR�ɲ�x�2VM�^&�:�����q
�ɉ�������ï�� ��=ߛ�=���v��ʼ\~آ�J;�R�{#`T��d 8�O�C�l��Ro�`i<I����+<OXb�^0+�������4�^3��hi��q�j韙.����N&��L��=��o<�k�O�y�s�=��sﵮ���*Vn�W��:{�h�'�]$�]2i�'���rw;�W�I�~=�t~C���|����m!�c?ȳ��>f�<M$�?"��g�bA~�~��s<��w���>>���>C����P��aXT��?y�@�*��]7�$�T��ċ�l�M!�}�i�{d���S�>d����I�+�Oǝ��>$��G�G��������Kz���[wx���+;�H,���Άd4Φ��~�����Pğ�C�YP�r�@�VN�����6�R��)1�Y>�����m �z�{��A@�T��$������H��VVLX?*�V�R"�i!׌`�r���guox����%<5z����mM��Oŭ5,<�s�h@�`aH4&��M��5�)F.`#�n�dU���za#c�'�����+F��P��3�[R]ǹ��9ij�Zv#�U�*3��Oh����=9Z1"���?�.�ܸ��)ǃ2>��d���R�"��NO��9��%K���
��d�tIG��r��Oc��L��	`mQCHdt�P��y��6�E���o�����)���1�\,S�6/���k�,H�����O	eH�|W������*�h����E��[<�Y؃�������
�g1H�Ⱥs���P���'ٕbr<Q����U)$�	�]>VU�*�-��F�v��W��7�)"�}�����{�{�$K^gP��Y�Ϻ�{��Y��g�wsҺʰ�摳��C����Y\�v?M]��7��y�|12�;Z��sm���1�t��'2�=
���2�q^��4O��dr�L��a1\IɆ������YH�Gh�Nz3ݴ6,i����.rL:4�m��8�gA7$�6��]���������^F��t�Bk����A�K~<����x�i+6�<��ej~#��7P����=��v8AoP��\��������.ခf��'1��%����b�����p�Be	z`�L1D�
�ˆ5w�*�`RإX��,�n�[��dy{XRV��r7[���ˬ�]���/(�v�9��WX��i��Gv�}+3&�|�n��^��"l(�WԎR��=���p�5m��ȕ���6=ۘaƅwc�Tu�j!�鎇�Q���AFӉ!S&�պ��U���ל{��¶��3R9���k�q����.�ڛY�6s�y�˃��Mm�3���7;�)�-�Wf��C
����T�c� Z~���3*�Ǟ��]Z�^6R#Q�rm�>�z{�Ae-|}`��W���uZO��h���u��W���e5y�/�$���eu�5Y��s�إ
(j�-3E6F����^Ђ��	�}�׫S	��|��>!PO7�)��}�K;P�H���7컐�As;��a�c�t�v�4�����}��Nr8�;�n\ߣ5i;hq��j�JLh�}�.�&"����$[H�.����t�R�f#��e��u1��V8��EuҌN�.U�cF׳{|�7�օ���2r`�s6P�(@����%�]r#�ڡ�#cb�Ǘ���+��9.6!�o"�+���~<W�#�|�8�ޭ5S��#N^�61�A���̿�y:�d�X6����_�J�Un���G�*e��#m;�.g:N�Ŋ�F_4�)���V�h����{��ymҔ�z���n�͸�z3��|�w2zwr��K�G�s<�t�>�bwH��~�W:�/q����:':5��I�5�W
սEu}���'����$���z~򛁱ceW�z<�z��~������X�5a˔��]@��m�ޗ����{��A��neκ�!75��Ȃw��p��@��S<����':�\}*�w1��vſp��ݼ���ʦ�n��j*
��� o��:�12�.�!f��A��!�XԺ:x�Fd�>�ch^K�^a��.�^;�mh�-F�řr\�iw�'�38k~�l<�A� ��٧J�������.s���2�PI�A{�p|s�t]�K��>vqw�{ں+Nal���a�c�)�h5����u�bx�
0B�q�T��42�voXq{9�����+=X��qo.�B�g��~�˩=��(E(О#x��.�Y7��E)��b�\!C�w�}���L�	�xkS�#¿ 3�ҼL��ȣ��xJX�懲H�bT$���uw+]P��Ƚ�r��8�ߎ�6�b��-��r�w|�b��#w�����S"�=��MW�p}*<0�p�$�z?kks�>�k�n����V��8��I#Ǔ��\y	�Фr�mb!�s�C�^�R(�Xo��MT��v�f�*��ܹc/e�:9t΄r��lok�*ǃmg�Ԅݎ��#RRc#Ȏk�2#�jb*3���=�x �Z�xNu�#�F�TH'���.��=�\x�9��,v4g-&K=�/���	������T�|�!5�o|��1���AR&QVgP���67�W9%����{nH���~��{k,3�C\��G2I�1(@�.�*!�jv`c�iKГR���f��"g�@&XN��5��X��,E�J���(HDoc�9��f��^�wA�������'�za�uZ�<�<C��r4:�b��2M�P�d���֭�C��ͽ�������@�|59^�e�7�=��.��б~�g �+/�_�2%^v	عy����Z�3^����}f3�t���()+˜Ra����q]��P�cpE�C�Y��]4��;k��W�u\�NGJ0 ��l�>�k*2�v;����Q���`���V\:�αTO6�D-�����u�d0��Ft�C.{�Yt�1���6�����q=S]��`��Y��iޒc�Y���������Mx:�ê����8��R������AXd`2�]or߈H��Qf���YCWLPT[|�ؿE3�+gV~ c�m�~�@��W��'ؤ�|�����j�8�ٷ��S�T�z�]�`D����RQ%�ў���`+7���lÅɼ����(d�v�s��w��4>�� 7݆�Z��_IѝS]�>
m�x�Rf���x=,(Y/(;�п
�Whf�6�xʎubIt���g)�����Tˡ*��
29�x`Ǝtb�}p�AbxF���x��UĘ�hS��猝�ʡ4=�b&��':n�<v��k�
3[9pS�nymV��楘��dD:nh�칢g=r���w�q��<�o ���!��Ȳv�YZy�O���:��˃R���I����B2�W�W)�����s����#��no4n+��rW"rx���J�/��+o�P��ZH#H�#.��Z1+�ܧ'ggU����E!ʤƮ���Xf�<'�9�w�ԙ�+�&B��*Dh��������[�:�Q��II�Y�b�0b#�k����:[w���X�A	8Ea&�b�)L���w��@�0!��DZ?y9mJ�9E�`L�F�y�=�uZ�b�JH�[]�쇡�Tܱ�@��gK�>�j�.�^N��Ƅ���"���ҽ�8���	�}Ǽ�,z��3V�bPo<����6l�_z����(:^�n�I<%u��q#�x��T�Z�­m��E��/����x�v��.ъ��l��ת�nLQ���-ͻ�f�z�{b����F�=�{�!���Q\�"u�f[�s�|V}e7f������ ۽k8�KWV!�?{��]b��J��k"�#n/.����a@�����NeȆrGݫ���ު��j�й�%�d���1��k��������v�;4���.x����W;�SE"���{̳�/��&�ɼ�a�BN9@iTF����
��,���}uF_�a���/�)��?k̷y��̜e�/��߈��v�cӅsW�w��^�.+��?���q;���3uu��]L��z=(��m�=�fwc��˭�:�u�kzB����tge���:N+)F���*��M?V,�+���`K��|����N�ܴ6��9�����zk.x�DM��ߦꌹ�7�+D�
єJ�>�V(m�� ,Iy�[��Uuݬ>7���2N����%���ki��kvnzՕ���Ž!ڼ�@y��c��)-�Ү/,���f��=Q��,o+}�:̕��'>����B�g_�]�c,פ���@:	�~S�M��te����G���Β�{��b'�e�0�,���`��p�S��2���^�m��	��Y֛�jY|�rQ��a��s�'����k�:D��a��=}�V����9�/���4 ��ĺ�W5��4ưˬo��ӂ����x(�|�c6""]��*`r<g-7vwG�E)о�:w����v%�0�o-���_y�غݩ��6LZ����s9#ݘ"�w,׋��bo5Z"�a�N�����34WM��ux!�@�·�qB���&���n�,��I�����W��/��m���`.�sw�
�u�4��.�5�����ўM����=^�Fn������m/-:A��%��G�ܾK�<j�2�c�n���#�G5-�(��p�(�D��zߖ���"ZXCK��$�v+ɍ�L��o<����͘�u��=m�q�p6�d�b�;:d�0��7x-��΂]�ۚA�h�9�&��|V�2�M�W�n
ǣ�g������ƶb�y�b���!�N��+mL���{Qv�ӕ|s5=X2�n��M��)�&�vf˴���*��m-�
������`~��-us��	�%���>}�L�e��c/��=G9�[���\�̽3+v@�lýoQ�ɻ�ӯ��;�#-�y, M��H/���_s�FM��eF1��rU�t�4*�U���3ˎED�K�1��I�w}�L�YD�w�D5ٯ4e/^g�BX(dW�s��:f@��y��Y�`��3g,M����L��ڊ�m�5xÆ�	7��P�����I+�;wS7���&_گ&n�����c�a��Ϥ�R�oG��GҮ��4�z��Tb�D�S����䱧AH�E��kO]FWc��D��<��X�(蛗��}�Viڍ�����VM5�q7����[LX٬u��u�k���^�35ڡQ��0��!WɆ-u]sSp��)n�ْ�֯��Z�S��MI����At���{q��+�A��!�u`�k�PMb<�J;�%C����JgsD��
F�k�M�ٵ*����n un�l��'��x���Y�XN�%Mk�;-
8-F�ЭWe);{���$��u|���!�L{��d8�[�\5����㕘G������Ć�h�1w�>�	������}�@K���z��'��8j��ه�`��J��%�[VG�Ν�"��;V��M�{-�5{	;��vlI�{é��Ml�v$,�躥[Ǐu��{�c�JbS�hK�	2�v�+Զ�a�e�:]妣�Br�e��u�	�P{�w0X��p��b�y�$EGD��!���L#�Ka��-.'�=#�IŢDu��>`��j���B��N:�����A��ˀ���[pF'<�p����	��?c�Yjc�;���[MK)�Z�%�:P�����^�7����u廌�{��K��I1n[f���
wF#S4:>���q^���������b�Z�"(PQTV[UV(����[eARڕ��(���m`�Uk�b"5,Db��Kj"����-A�kb�AD�V[EDV��TDQ+(���",-�F���Tb""��4���Ub(� ���D��P�F�[F6�(�b,*�#�A��"���TEH!iD������""���TF,Db
$APF�X�-��UH´Q�*����������DH��1Kh#$�PDUDDQEmb1EQ"DVdVDTb[Z���U[J,F#QTV����*"�")Db
�E��((�KeUEb�b�DT`�EJՋPKje���Kj��"��DH+Q�Db�EX�lR�
��b�%lTQQR"ZX�(�H���T�T*��  ]��+��}5�R��r�Ӗv�R�(FI���wc�v3u�9����h6�}.^^ ��r�{��'ێ+��һ��l�K�������*xMXL����my-��^.Ⱦ�浪K0���ֵԽ�\�T�0��o����պ�Bb�L+��ɚ� ��zpM{���/��4�J��%M�]���%yl���K��[�g��0�tQ�9MR���U	\�,Պ\�3�J(�כf�(үi���vZ]}pXuߓ��N�����Wt%s��ݩ�6�6+�jWJUYv/�)*�}&]XI8x��f�Q��ta���u��x�p��=����pI+�g��y���Z¦��4�9�������	�1כJ�k�,ם�+�UqM[��oz���:�c�6���mSu����X.H-?M�nX�sb(��S�]c͋���S��?J��]^�{����m+��N.�wk	�q��n����.6ơ#-�3%M�N�^t�y~����OV
���O\�*��.R�X�=K�.�5��q_E�|�QD�p;ܷ����j�v^��p��9Lˬ�j��#t�O/��^l��.�t׍Q�Ģ�����4���<Ē���$ܔ�n�Uݜ��ǫ��Z����m�ޥu57/�T��Ut_4���|
����}��#4Ձ�²����b7	-��ݽ�c/�.�0­G%RY�E�6�f�k�^A�+.'��t`��nﻸ�GUN6t�	���0E{M֋mۤXK	M���?"�\C��U����6Fo��M��Po5���NZO%�tl9��w���pݦRŦ!�o���������a���0��B/	E�	�7 �[�����<��6��Ox��iX�NI}Bd|�y'��z�c�Z��l=��rK�MS���N:�%�^���Յ�v��=VS���RJ'���������͇Fڌ�y*�����1~�\�q����δ��M��[M,r�<s��ݾ���S�҈K�Cv:3o�3���{�Nc��7�&Z%���Q����lG�o�>�Yw���W�<[�H�^�R<���;�����cS�կ�x�v�SR&kj��vN�H��JO�-S�]c��N7�m�+/3 ǊIW˭�˩ڏ���;s:��H��U��3c�jh�&�֯�.��=�j��j�B���vDثuX�T$e��UU}��l�&��!v֊+oqm�>X�����[lQj#���/`�ƞ��+][e����!�ͥ������z��g \èQR�Ɋ0���/���̡Eګ��F�v���������ܼU���$�������袒�����/\�+Ү���qo���a����!�]�<���Mm��i*�fog�S�J�|�mx�kF1���ӎQ�v�|��;$b�f:;Ƒ#1`�/�S�m��͞�����J6q->�KV�����+�J��B��!\Rn��v�wK�G7�AY�/��R{�Lګ���H�[�oԂW����b��T�^��|X|�wr_wr+/h�+��ҥ�xT2�T�2ҥ'���j����#�i�{�F
�z��i<�<}@"�����=&Yo��F�ǫ2m�
�vd,�!��*bm��%o!���M������-��C��ֳcss�3��>�7�e���Þ�7�]���&6�$��V�o����e�k#Ra?skU:$����3�˷��#`e۔�J=�8c���I����=�_}���{��J;,ѝ�G_v����cxM_�9��{�H��Jze��r���:M�a�T�.�a*�H����u��NM.O��~n[�r4�K�F�ie�v)�	��7�P�Ҭ�����{[��V�t�Z�f�y}��K\il�:�T`@�qF�
]��:�Ҭ]Xm�y�:˫�z�QV�#�`���3���d�SL�O��랯����mOY��kf'k3n����c����ΣE����́�%������bVŃ[�{NW>2�����aM�؊i
�B����i�<��ߖ�5��-;�L�j�v�ܼx8�9��6;Sm�@��Y�s��L\�;-��7Z'Z���_bb�Fߵ=���5K�+e�ӛz�p7�Z��,�L\_I��(���.��i���.j�,�
��R�6�����Lʳ!�G{i��4gP<@Dݓ�aR�F,��~)9&>��,^ӵpْ��M�ʧ-C��XvBD��-y̱�df6�`HE%�4���4.�QFҥ>�p!�;�L�B�t��	kF-��(Jz��8���%snX�0=At�0oE}� Q�h*�Z�]%�]���VX��.{}H3z���+�/���
�5��Gvm�.�q��~��bl�ٮ�^A^D�e{f��{G�H�/x<\�]$P<5s	�a.9�٧J#@~y@��[��3(�ދ������X﫯XO3��[��W�I�p���R�\'����1�D��F�Cy����ѹ^zM�o����T�Fį)œb=΃`�#��u���$��f��J�V�sv!Z'ak������n�B��D̴��<�U���)x�	�p=�¦NB�J���r;��c���/�����j�*7��*���J�F�kJ���$f�K]��e$�0��x�Su9_H�9��d�r��~o�s�TԼ���g=�K
���l���I�p��m:��Yp]n��&g"����v�Sm�4���e�n��.za�[mo>�:��u�k\�%X�bX�Ջx�H�r���(��"��X�����]+"�_
���=��a�o.���l�t�T�u�
���.읽l�hV��N�6̎嗫�_}�5��(���ܧ�>�t�g�+���6�4�(s1��\0�bc��t]��c�+P'���,�=���>�uh�����V���hvI�j8G'Yz:5]�W�m�.��K
u6�1y���ʧ޺ǚ���c�W�`嘕:�����)+,�}5�n�����?u7�_x<r�nyN��s)|��-�{/��������[B5e�*rzP}a�Rs�zS=�V��M>j��~9��^J�މk;<�=�Ѯ��4���\��l�Ťh��b1��b�{4l!�)7H[n���Ӊ�]�b��]���1�#�k/97|s��Om��W�A+�J��7��a���ܴ�B\`��q�/:��ƯٽY�Þ��33z�RS]%�R��l��}��Нum"��V�n�$����s�GA^K���CJ��)�Y�d}s�����Q�ά��*b�^���f�,��>����}��vj:��SQ�t��J��y�2�7�..I��~V��YE��p�G��r�ln��OSZ$76�9=�;|�Ot:Hs��Z=ړT4鷹w��۩jS}Mv�\���2,�Ho�{�
��VBO�d���un��q�߉BG��s�B;��x�a�i>�k��h�&����7�F;sn��S�U�%^���/�.q\F��܊�tʉ�њ�A�]+�ig���&���֣������9cMuwNa�Wv��j�l{q��eZ%�l�NX��m�'Z�3x�s]�(�Έ����|��[J��f9؎�=�-��oy�ĕ���lTYBs�l|qL]gm��2z��p:Ϣ��7(yY�6�/cQ�>�	u�[�{{�Z&n�1Tm%=C)�b)49�ʮq�1�������Fޗ�`慝8��nOS�\+3��{�\�x�s~�E�)g��Ѝdn·�V��-w��U�N��6g	����^��#�hs�u��y��lmՃ2�[��{�x�I��ti�#��Q�4��*�&ި����v��b��j�_>����a@�}�Ɛ[8e�CD�/��jm���N����-�A^;=��5nF#��%Ǜ���x�h8<���Y�U*IZ���6�5��A�w�Űu�vHF�J����Hb����o`�;op����n;��>]{-��JWJ��a����!
�u�۰#��b5����Kk�~I��>�ȎS�A+�ޠ�b�紧}��Gf�|���]��;9�����k�.F�Q ��S�U4��%܆�ufF&t�r�)!ʸ�6nЩ��׼��c*��[���"�����l�6�����p�=����3A�5i�y�����*�,*�̗p��U�����$�����o`�z���V��_v����9�H'�Zۂ��(����4��.Ln��=v��zU�SK�?:�מ�{n��	��;��,}��"q⛱�R�'��3V)vߴ'��qEՆه���SSz��if��VI�
��V���׌�2�����>{ݳ�x��s{�U�\uB΍��#�i��Rlp-F�:�����Gd#�)�7������k�H�o��z� _3��]=�� a\�P�}]�]���"k���Y��A��ӡh�('yp���V��n�Txh�m�\Y/�0��W|�3\�8䕤K;�V�K���i,��#_Y�VV��;��*���'مw����1Ҭ|�F���xʺ�baM�؊i
�`������i�wO6"i�1i�Gqb�`絹x�q�pja��-��-f�g8���d,+'�� ��]��b
�+�S����冩rT��,=}�åP�����֜�Q-y���r�N�^�ϭ�65	���T^J�Ɂ1�v�n䧳�Ŏ-�Z���чNb{*�צW�\�C|`O�^�qFPTߣ��2H�Ur�"����[5�/ נ���V*Y��@�W��=�5�{)�#�bP�cm��x%�f�Z��,�)e��n�~\v0��['ު�iJ��A~}
��L#����`%�	#IH�Y�RM����v�Ծ�RJ���+Ot���ϡS�j���)��Rv�������'N�}�����3�SS�>y�@StK{����ds��t8)�E��sI�̼��('��.]�3}���b�H�P6�p�a��YJ�3{;_&�R{w�>�n�$��_"����*D�J�DQ:��ʤv���-��{U�ی=�.�{ܻS^Z��Lqe���릣h�i>\�FcV�[�!T��� =ة�.	f�Q�K�K��GL$(G&s�V�SJ�Q�GD��CGM]��ΚFyYMN�t�x蔦�"5b�;C:4C2{]��ŲN��A*���%�r�<s��w~N���j2P(��ً�������7S�����fZ&��N�8�i�h�^��,�]�{��±b|_n�,	'�=H��=���IU,`��S3�ʏA��)]ͺ�;v'+)gY(��ګ���Z�(������x���v=�w����\t��e��(ګJ�o��1y��<�޼y�w��n�$w��o���)%�C3L������un5��V�;�-��w?ql��^Z�]ƽ)_I����*�-�Z��^�j��#V_��u���%�ұ�څ�d��V��8ɋ�x%SoD�����5�]��j�}���<��׿b��Ŗ܎y� �KNC���H����.9��H_�7:V
nX��+r �t�A]�룄���UnhEWV]Aג.�Lq88W����!���h��9��`3:�t���#Jm�;3^�NL��^���6K4F�����v��|��{.3�FC����ϻyL��/>�Sn_j����寭��p�L�:�ҧ�N�]q�h���y>��bxi�w�vشĘ(U{�^n�C4��u��ⴭ�y2�ƦQ����-��l�Y9�_
!�:���:�{���<�Q*�T^�u�{���d��]k�w8�,�-*�8�����*���re��T�Q�\3s�ROv87É�q��{��{�Ӯ�=�V�<�pn;�z��ͥe�ϕgD"�+�Ȋ��󕻭�\-��H7m�?��cU�-������gb�ڙَ�Dҧ�^C"A��xO*gG�0�o���������RN����n��V��8K�i0��T⯈�W�����0.���;�R��b�&��Sr��v�׏��b��֦J۷fB�&�����b���bz$ݚ��d`*9b�5i�A�u��g���i5k#�j[�X��n�`���v	�1o%J;E��k�}ȵ=܆;�%\Q�(r�����ں��mǗ��i�?J�Ku�>�#�R�05�r�C�-��	\=�Z7F�)���΁Z{���Fc��ځ`�,'�*û���t8v��hN�u�;^4̻������b}��bse��,����A�Enf9�5�B��S«s�؊�73��1F�\�%�s�k�J�F��_��@����V9Ϯ15=����z
��%d8!�|;v�a�jg�ȷ��Vس���˕�}�4�ݵ��4m� ����wr��2��^���E�7=�=�_�PF�_�ҽ�&]v�gze~��[ZV�3-�;�u��[�e.�ϞW�tY3mZJ)��<�~�Sm+���� ���.,ܹt3BcVt��������f	�������Ш��\S:O?ཷ�P� 8	g�4���t��Ӎ*G�MCz��b�y:�f���X٢\�h��R]����JK���HXr��v���%�3��9\��ؼeL"�}��=��c�]Ae�8�z�.Jޤ6U�1�WA�P:�}�1�H�^T��t�t��k%�9Y���X���\j���U��i�͠]B]�C'2�-�|���6�*(���͒��Vٲm|���w���.9�<�?O;ɔw�N����Y�ޤGDu(��W�ͱhJ�W�4���!��M���n��J���R8N�K�XtI\�q�X�K�+jZ�2��Sf���`���ǯ�Nݓ	Q�nlZ%y���^)�;m�W6���ôi�1ܜ��:�'h�Y:�ʹ.}6���bSOr-u,����ta��j<D� �]�T��+�$�kC�X��r���M�r����>������EXƥb���jUD�j�DQDT"
��"����*��
��"h�Ԩ*��DX�Eb���(��"Ԫ�QbVR*
QX֢����YUb�Ȩ�F[UE�Ŋ�b��E1D(*�DQ"*1��0PR(����DEDE��X)U-�-���E`�P��X�EEE���Kj0TQX��D���ATm��Db1������DX�,Db�+Pm��-lUE��X*��"DA�*-h(�!YXԩR*�,X�����("��mV �	Z%�R##QF"����
�`��*"(�hU�b
�"De��c*Q`�"�"��-�AUX�R�
��UTATF((ň���*���Q��"��� ��TDR҂�bAb��U""�
�*���@3]��4'd�M�� ��]K�p�:-=���1#��q�v�7DQ�c��0�g.)���F��W|VT�Ǝ�9=�����5�+�66iXB0��Sm:E���ٮ��Q7��J��|���P>YUe��j�cPo5��>n��DwVfm4v*�}p[=(�:����1�m��xX�U���¥������#s�h���׼�Ʊ��1��,�y�GA���O	�=!z��� M`A��M%n�0�y��
��y��Ƽ.��ZN6~J�t�B��/s��eeE]jg�3�攐�f.j�Yys{�v�ão<�`/%BNF;�yu��B��O�Wu1KM�F��`���a��۷�gyN�B�����;��$��~ ʥ�e�F�*�.�ͳ�@��l�td̊,z�V&���z�j1�ܼ�zeˣ5�U�7�-�I������K��b�監Q��D�M�=��Ȱ{n��v�\�<���q�$6��X=X^�D<�e1����^�X��l���y�C��!g���XxS��Һ��(�F�R�ܔ��0x8����yb��._Q|�=�<�PU�,�26��W=:�n���,��*��㱜��m8�I�UӺR����ćފ��']�iFN_��XƄShP�cj���Dn�=�W�F9ʱ;��};r��إ��꼰!�s˘/5ӛ�E�)s����~��k^�h��J;rz�3C�\��.�����3����ͬ�6p�6vkX��ں�Νh�p��`G>�Y]b��cP���i�
^��s�6{o�R��Ъ2��2J{�Lګ~��Q��9˒ill�CB�����>�9�z�x�Y�[O�kf������S�H%`j�cPa<S;:'b�7�C�T୷����ȑ=�;� ��_��e������]�w_^OrM��%��`���A���M�؍{~�<�`l\�ͺ�X�z�u1�Ve����b�	�KB��|��3��ͷѰ��F�slN�sWӏG5�J՜��(F>Ya�a}b�v���H{n�Ѵ�w,؅uQ�5�̴�6�2����ߗ^�L��m��(iZ��=H����(�*t�]m��8q�I��=��R�:b�V^�u�4�V$,�#g�9���Ik�ʋrR[G+��Y��л��\7��x(�rˎp�^޽fΖ����[r�����(�O#.�w�xR�{��U*-h�4�_6��ۡ�Q��T�c�\�#׵�#~�l)��(�;]9��[�%8�yq��]+����W�9"Ł��vw��8� f��+�X�v���}��r���q�k��&i��V
N*�`���4���f㲄��b�UbęK�kM+�`���Y�]�&�؆��f0s��ˮ��@κ��zD�K5���sj⚫c�k[��_9��v��B�Y�Xv�v���S���D��Mw�wF)��<s��l�c�3���9r/�;N��m�K�\���a.�Ց�#^\=W���. }���UE�M�����U,3vIh���ⳛ,�k���4j��O�]t�7�Y���k�j����%��H~+I�T�	E� �+�זY��;.��A��T������D	�.�`��Y�6y|�Eǲ�j�d
:��5���Ubs��4��	Û�N�t�MK)�^�:�Zs��0��x���z<�=-�t�'f��3� �G���_y�I�z�Z��|^��Y��FR!N�ʸ��-̤�V�	[y�Y��죧�M���"��j����Z,%�5Ԙ�"#�(u�|���`���0���q,T�ت��J�A����&��GN��V�FhQ��K��mi�,O	�ةn`�Ib����TQl��FaY����Y����=���Q��!!^�����+��V�����los;Ij�Um�)Tk)��]o�.��T$t�HW��8��ZP�Ee�*�u�\�i�H
~�Sz��n�94�N�Ja.����\�	�
�nD�\fszҔ6�[����a�������^yN�W�0�����:�}|��g���{��[�d��e_�7VN�1��:�^���N�]hƺrۂN	&�������Q[cqn���%uak
�c�iLm��ʇ|x"�%k�a7��|6�J{���xr���j��=��똔���#��#y�}n�s/l��h�G��j�<z�u.j]ΒN�=	t��pڲQN�#b�)U��K�����lG���x��Z�>��c��ϵ�8�ZCǮ݌)�|v>��GPY����JW����*3�>�	����e�=�ɷ��݄J;S���
Q�V9���n7kұ�
Y���o����z/�i<7I��M_����u���ڞ�aq�F�q����O��6s,�]�z/'a��$�5��]v^zU>Z�u�\�������/����ޛ���s���=��;�'0e�eSn�!�{�k����n�8�����ç���z\�x�ӿaV���r�0��{g4+�ʄmV�6���f�](� �b$��f� ��cPo5����B��Lg;���������W�p�}!+�����Ib�w��ۀ�*T��C����w��+{L'��k��y�DU���s���ت��F��B�3�G_v�K�,����T��P�hb���n��WUVk��E��K���k�������ӎܹ4�)�*��K�:�Nt��'�-���>+����z�&�2mdΚ�:��PI�*�)�0L�A�'�w�sƻ=������w{��5W�{7 �	brm�ٌ"nT-\v��2b�n��::;qi�s��9�{�0�,m��C(ֻ���3_M=�3%D���%$]CIG|������b����zQM$������Cu������)�E�0]��<��v��L��V�0�1ܗ>��,^�؞(=f�=f]Zc<�]X3X���Ԟ��[{ϖ$���c�Df��&NZ�)I)=qOܘ��Es1����E�:�Y��X�ūb<hӜ�e���m�2�����PUh�'S�ۃ}AN���[�kTq�U�X���K<�Z���]�����e>��CES�x_A�:<6�'����o�5��1�[�^z�Fޱ#-��j�`J�|�����׽Z�ch��v)���o'�utr�%~���RpoP�(Śe�����k������uĵ�铥��m��v^A�՗��є�0�7�M�B����.�ŋ��D��(�5��k��o��`D�R̠�,��1��yD.�Ŷ��}�c'�VV�)������\A%wP>�y�y[륄��O�tcI�qvl<P�(S�4�i���]څ�K.Sй�k�&�ۗ)�l��c[s/��"��Q驇�k�jsi,4 pEs'w6�+1j9��d���+�5�7{�Ġ�"9�M�i2%�#K-DH�¡�u$�l��y7��v���`�|�8{{X��5�{����Ш�y���:��	�ݱ�-�r��r�1��S������Щ<�_2Y�>xMXL��>��c6�Y���O6&��d�J���4\rG=au��T�0��k}����7�#Y�:&�]j,�g5V��Ǆ���@鄅B�j���3:zO�xz���2�h9m��WI�U��*�x�aT%p8&jWf�L]�.�9���D˞��g7Ke;L�<q�j�l'Z� U���%b:�ҹՁL�j0̨�[;�Ė����T�N*�lP-F߹�h����n;� �a>�Bڎ�Wgq��>�m�M��	wV10��b(��s1���ۅ$�����Z�<���������U��3�So���;"��kݜ�ا��O	[	��7�G���8����\·��"nmp�o�	��{A]ԩ_Y}�co	���io�n�ž�:h�ǌ+W����W6ּ)!EN������@���$��h�c�Ue�e�[�:Y︦��|�f8��ͣ|��ٽ��#/`}Y�f���ƌG}�+�K#oSܮ\R�	[.G]��y��SY����Rʝ��k�
��v6�j��]eu�.�j0��M�#L0uN�[ۦ�/J:rܪ\�ޜ�,�k���6������X��課��ں�̒G�,fn����(���Z�V��4��(p�O�̍�R�X�JG��`�'p�+
��<�v%��ZO�f�Z��Wq�15�+�t�U�"�u�`���S).��V5� ��ЈM'��N,�j�k��LV�i�\�s��'��%ߪR��^Kn����,���,����v��#��uQ�Ills�W����++o�ͅH��V�A��괹�`����yF7�պ�X|%��T$t����������=j]j4�V ��¢^{�k��n�94��tJS	{{�5�Jn���;x�hz���<�A�p�$Ӳ�ќd:-�F��Ll,
O]��qJ#�1ȋ���O1Q�H3��yQD"�ȸ�ٌ֤�W|Ʀ�
W[�1��{��if�to��V��p�Jo��M<��i$n���2WFQ/	{���	�3F!�m��<��W#7~a�c�W�X��V��ߓ�x�u`�%v��7N�N2�]�n��tN��n��V��I8n`�~N�E��P{�a�-?)�:�_�0-v�{^��_4�QZ¦ر��C��¸u]׼G���>���r�Vg�W�lm]���P�7Xv�Z*ٽ�4�������Т�mU�Q���V��Y~��$�U]<`��z�Um�N�6���`o�~�o����ڞ�g^�dn���_n�#�ߦ$����'�'�H��un5�j��*�-�Z�����lmՑM\�l�rz�.Z�J�ʞ���ߵ�(ƚe�m薳�6�k][�nr�%����bI�"��;p�/�SyU���ZB�&�m�a�/(P醋tVZ�oSt�r[<SE��0Y�UԳb�JƪZ�w�3�7^Ea��������[<�WS�C-�w�Z��Kl��ȯ6��n�������:jv�RY�\RuMнHyۧ~}���'.��O���{��߃�-/:��Y�nQ]��I@�݄�q�Z8�IL�VS�S�mL5۩�W��븁#�!�1�Ҝ���7�Ou5$��9Σ�� ���+}R����UL]�!�Tw��F�y�9Q(���B�����y�}��F���G���WA$\���ĝ��H�'V;���h������î��l3���:�ELrc;��u��TWg ���
玚Yyv��x�˓O���%�9y9L�]�D��YbLn�_����e4�9f:��������5y�1-���N<Q���밦��\��.��ߴ�W�K��a�Eq�c��rn.�Vն�����ҧr�u`�5b:��WmX��mf�>\�;��J/5B���)���n)68�\�h��K"ٱ�������6�͌��-G+r�&�����Vp.a��^m
�cj�s�^�F�n����;��۽Y��#���,Q����Ŝi�\�y�t����N�q�=�q.�L��J��]׭,�����9�8+�e�����`�Z�M����rh�^K�w�����о��.�nu\b��8�-�1�{m����	��O��j�θ.�&Ns��q���T����H��\�;�"eB���7�u���y���U��:-#�e�%����u�&�� nÎ��O��(���9��D���>�Y£��Zt�+���wE�`��!U����%�f��cu��'$��{_�leJT���,��Q#An��.ӫ���g�XS�xAM\����$�]��9])X��N� �$�5=�T����*M��78��a�֠�2V�f��8�T�-�\���Wu6m=R
���m���Y]�o"�U���L�qЦ&Ir��.�O�|�-W�jOw������cn"$�P�xo|��8C��9� �s����F����O�TH=���u;�Ss-�*�c:�i�V�u>ʅM�m�����D��p�W	GI�L��A�h�FUlb%O3�[q��``��!9�O�󫒢6��x��pE�n՞�F��;��m+�~�p�I��x����fGQh�x�6������9�3C{��Ǚ�L����s���ag�eJ��b�)<2|����3$9X�8cΌ ��c�R:���8�A�;��0o@�>'�۵J4'K�����i�4�9�/��Zw�[AS���	`V6T���f4݊DɉM�ď[��|�xih�N't-�|Յ�S��>���7���Z�^C�o`(iS�~c+$m�T73�̑m�o�#�Js���<�]$LꙖ��VȦ��.�h��U��Y+;�mp�׀�[��>�^�����+���7�av޼"���nr:tV�1�� '��s
��ڣ�:4�\B�V\)����΀�{��|�"��S��&��V�K~�2a�1������ڼ�)o��9)rb�<L�l��3�%�0̅�q���3-��}�ݫ�����b�_;�K(_��=K�g��ƚ�w;��ʑ�Q�����Xz��sk�p���쓭��D�V��i}�p��+C�:��s�z����X.e�a�vX���?F�e�[œ,�F�Vt��>ˍD��8��ۓ/!ٔW�ɠcma�n������)7z��h��%�^"��ر��I��Y��t�[H���Z�'`�N��-�Ѹ���q���̅�cBr��wOc��ߜ�n�])s�j�9�8�[�:�A���4��|�n�5��]�=�/n���m����J�t]�6Z��7:�Ò�c3[W�	{�süa��tkeefૠ��̬Z��1�e�Ѧ^���X ���{��i;� +�.�@Y����w/��n���!͹����&��Jnom�j�R�-�2�6���oa�')�,�'0��a�w�Z����YE}}��&]��c�<�����y PD�~$B4��Q�������TEU��,UTj$QQ��R��mA`��V�,�Q�kE� ��Em�h�څ,�""� ��ѵ��AH�"�l�Z�T��$Eb�`� �
�6��UQDE�D`������#X�"��
�
��*�X�j,R1�ƲVڱB��V�UTEE���(*�2�5�1�E�#"(��JmYPQ�Y*�##��T����E��,�XV�"�*�ڍaUU��
�m**"�R*�бF ��dT�Qb�X�l�PF1b+Pb��U�%*��"%�`�Tb�"�5�E`�V�ȱDb�E�TX6�U+X�+�"�F
(�����QD�H�F
D`V�UR#"�jő��%�#*(#�VE��X�@��A�T��_�y��ߵ��dcaЫ4p���rW7%���͍U/O.Vl���s$�RY�Đf;����I�}4��2�Wsk#�"�'+�X��h��Gs�m;���-��_-l�\"�4j(��gUkckލX|++�Rplj0�i�
^������A�D��%;�g�Yz��4�`֍u\�.'������(aPd��$�m6��Jrn�����:�Վ+�V0�Y�2���H��t��iU���=��4<A��k��x!.+�R�;B��QP���h���r���-�f���W��a�=��)�<����R1>�N���O�e��g�-Y^�v�xF>�%u��!Z{��'Y�xMrf��9=���g�`s�r�8�/U/���K�Y����wе�k}�v�ȸg+*�ӾjF�S
�����!k�]CJ��H�n_t�%���rQ�$z�����Ox:�j0L�̔F/��je؜��c�<�t�:�=���׭)&�K+2����w�ޔHl3�{A;U�U�m���Y��r�1!b.<�Dx����VF���'T������4�<Y�:�LxF}����3ZX�-��ҍ�M����ȑ��������դ.��di�!+���&�6�<s������+皌�r����hSI���{�y�Vpm+��Y��0�������Q�9�h���ȶf�;�j��I�f�����Gv�a�]ΩL)�؊!\�`p����j�|ʚ7Qô��)n�<}�����q�sژs`c�3|���9��s�L�Yh0�f�bQ�#��ыܪ���Y�}�sep�z���"�'e��$�6��������r���(���*�&�op�Mǆ�6L�����aK�|�Ӂ�{=������j��3�f�
9<�0ۛ�J�q��W�j���^J����8�V�� �T6��K��mR�=R-��;���o���!XT5M����ZS]HQ�#����h�{=�OC�I-:b�1��I���T�j�kn �6�}yz�L��:�wC�I�y�T�I�a�z���[�x^ԋ���&��������ԴS��:��F�M�U��#K�&C�%��19]�%a�Mu��4&�W�fץ`s�g���ǵcN>܍����Mrk��	���<����6tUͬ��A3��#}'?&y^�K*��Iީ%�-�V��,>��a^��"��Y��ҼO*�O������t^J��	y��+n��}���U�+�cuII Ur`Gk��7O�=K�|%�~J�#�	*{�Vx%�df�.>�f�����ԱSK!�$�3�ݺ�F�)�)L%�@Ẍ�l�:���Hf�.��`R�z	�a�w�X!�<�u�ּS���N�U9�Kp^$�$�s�p�V�L����Eu`$�<r�j0�:&�L�m���iq2�.���UjY�W����yMG���URL��R����z�#8�Ĺ֨�����!�6�������<ګ�ګc�kr�����֛⒌��$*c��6�j2��q��So����;�G��{h_[��w�Z�R��`a���������?I�z�q>��.6�͈�P������J"�~�� V*�ܺ��^V*xZ�ku��G�Qh(=��&0����
��MŅ�Ĳ�!=������q��}�J%��[IE ��u�3kf+N��hfڻM������պzf�E�d�مR�;���=M\�l!X gN�!��=se��č�j�)����r�ȢuEd�|��Xu�5�Wg���we�����m&���������!���F�̪m쵝��{֌����Sm��3j��C�'.'���@���<!(�L[m=�.T�'q���ե�ܝf�
��f�,�H��ĕ`T�(%کj���Of��4ݔ��*pV��]�i<�l��!#pP�SRPk�D� �����-�륒���M�;�A�g�B���͡��89�p�!�۷��6z�/t[�-t��s��i��V���K1��u~u֓��C�OY��F�0�*�-��f�0 �c�������i({˛�>�no΍�ڌQa6�;#k�#$N��~��U�\�#�zU��X�y�:���_f��E�u��Z��Y�ªң���.u+�-24�V�u���|7�bU��>�p����E�"fx<#i�neR�_V���罃j��e�֢e�/���b�=�����ʭ�҉ad�*=���7p'O�Ν��J;�K��f�=���#H�����*��J��YO՛QT��rL!u.��oG7��bwSR����
���,�b�S��k�8끘huB����k�s����̮�}�b/=']Z��6��+���K[7��Z�J�O�����mg1$���M�7z����XІ��s1�W�F#�kT��1b��靋�x��ڷ���Jܫ[�4��9�6�?'yHlf�`Y�f�q-��UA~��n��9�Yz����<j�%O��3u�k�5nf�a��R�]l��s�ckѯ.WY])��B}�2�HE�����2�_�/�L�^���g��k�אj5`�2����A�;1G���i-�(q��L[nè�k�)�w��n0P*窄�ܺ{3a��N���z�ư� �-�r�y'W&@)���e�)\��S�C1z�W7��J�c{����ЛI���{F���#�-�D��:M�7�okԱ��vz^ȡ��.��4vY�7 �MŽ�t�L���8�������4��I�q}�n*
H�ޡ�a�PڱwC`UKrCU ��R�$��Κ2V魉�Ùwm�c��F�q�Oz+��@���?^{��@����3E>�V��N,���*��a��7�K�i�z��f5�4��G�Ln�Չ,�ݧ��v��p�!/qg��Յ���v����[��X�VW�����]L*6�>�����	
���0��d�;Ǜ��XG��Wq�+}�IP�z��ۍ��v�<굨�+�BW�Й�]�ɺ�F��akJP�S[��Eզ�<s��W:��
�шK�{���r���}2'՞�jE�Y��}ڻ9C2�7WⓊ��Z��ΣE������7Fİk�z��c�V}�����j<}�/]�&�6�4�W�F^KZ���ڰ�5*�V��5��v�=ܥ��r��͉�'U���J��@���\�x�Y�a�+�,۬�kь؍ڕ��dm�t7/���*�{�n�I(٫`h����}����s�cF��z�
��.�/%�����#���\ʸ�wl>lv�Ko�8�c3��A�L����#rE��εd��	���]e���"�LҼ�!ި��0+����{�k«e��f�]t�����Sn�d�P-��%f�-�z�Ȼ.��:#N�����W�ym�9���i������ZRUr����M>zzp2�f���_F��Ŕ�T�)���0䩾G�`�zD�qe�*��^��+�k��:�6b﫹��RX^�:{�K۩�t�7�N��+�T5XmܴXKMQ���FYҽ9r�eh�ȼ��\�DHI�D�u$�SK=j��A��a��ЁH[:�v绸��w2����\pL8v��������RW�n����eN�c�=-�t�)�ߦO	��V��&-�6���6	�P�=	
��������|�1�W&�^mC��KeP�7�yWʷʺ��P^&�l�$q	Z��z.��p�o:-R]Yl�.劚A�$����v�ão���I�-�v�ZØ��o����VR�ܶ��Ŧ�~��<s����ߓ�qA� �}��03[m$������/�C��E�eѸ��)wU N9a(��!��P|�>�T�S��V�+��V�կ�We�e����JA��tx	�y�Ł�S�J��iو���nw�x�G�A�v͸c�����ס���}y��[�-r���p(72n���*f�*U�Iڕ�������c�qe�n�ޫd�K��a��+Y����|�-�1n���ߴ�xWO*�Uuv���Ƕ��E[II���1A�1C��97�(5���=����9�Y�p9uzY��z��aՌv��B�Q�W��lF�zV=Iޗ=�Ȅ��۫K��\&�����~������^ğunB5�Ӳ�4+6Y�~��5�~��~ϩ�cr�,5EB����u�\�_uwG	�z���y8�ň?v�Re��gPх�i��U6���pn4��CM,�˻������R6�F�/ Ђ�G-�FP'�i�YE��"�
�(��0f�1��(�:�4�XS][]�~%X,ؤ�T�"痱�E���6҂&���ͩi<�����|�D�<*Wꔻ#*���ޜV����}T1�o�{��*��PgY����T��̝	bK���z�Y}��~Ʀ\X�Ӆr�Idfʻ����q�$�Yn�f���;��F�*��:◃1�Y	¤i�n��Ӽ�v\�"1_��w�ru�� c�8ޤ*�+Bۆ�Y����]Mt�\�Y���'c�s$��t8&E��0o��˝�?�$'���ٍ����
��s%�����T_O=��k1Y�لƧ�G�~4��Q�V�4����k}�1۞
u28֕�$����N�d��
D?+�)s��zU��Y�9f{�xVp(�i�5���N�Uk�)����V\�Wg�����Q����94�YI;O�7�ҝ�'Z�k��j�mm'��A.�a�=Ü��K�,���?ww<+����6��E�Ƌ/],�f���7����4���-��j��?W��s���%����W�hE6�s1�V9��j�nA��jRz�<�%R��O#oK��Ŝi��s�*mp�V���5;7�N?,رK\������7�j�F�2�,�v��a�Q%½�k����=�+/&��|��qJf�=�*���I��7�
0#N=u����݉rb�f5�]E-*fkV�|i����k9�䤷\��u	��h{�](~C�1��ҡ7fG��QP1�{�S��MKKn+�6'�/����\{:�ji�E�]RԾ��c���U�$]פ��J;×�r�������QӖ�R�7�9���h�U������ѺA�u�&.��x��)%jL����h�݇H�4�k}Z}f"Dl�m��b�L��e��2%�״�}��@�A�p�N�r4�Z��LkWQP7ae��g��=�=��=�S��T��T�j��y�ۏ�Si0���nyD�7\Y���p�^YTh6,zL�ۤ��Z{��d�f7�N���m�[h�]]T�+y����?%.�xX]C_�	���k��+o3�c�J��*a,��m��:6���a����	
����9J�uY�����t�'�79��s�m���ׁN�VBW�f�\��H:g��s�H�S>���_�.�6a���\�Z�k� �$���Jk�)sL��7w�ݴ�#�7��r�5\RqV�Q�:� ����G�3r6%[�g+$������F�W�	
}7��*9���O]�ۊ�J�6�td�:��3q���M^E[�Śc�[���LT:�5�k��%�q�	s3�.����,f��>�H!�B�V#Yb|�=N�={-��*�'Q[g�Pa��91����Բ�9:i+�S��EگL�9�6DP������ݾ��t̬�U�[�֩vfc�Z���#I(��꾈�9��Av�.�Sp$%��M-$���V�.����1s�P��Oa��Ω�S�\˯Ӷ}�"د"�ҩ��[��wi�"��4��� ����Mجw��=��|��%��!Ǔ	x��P���+¹����k���юƵ�@��	Ϻ$���u���;y���=��{aܭ�$�s��ay�ۇZ����O8{�G�*{X�gs 3F+�E
F{B�|�4�<�gRrs��wFR����iѓ��-3���x޴�^�|P�vU�[Tz'f���S:v^�.����ŀ�xn���/����0��n���3�rG�r-����]fV�S�>>
=6��)�)����Pi����
*:��p;ӊi��.;%Y����l�U��NVq,�ԫ����_3Ԯ2믜�b��n���؀��9�T�×���n�ktCKZ��%�0@XW@a��y��9\���G�p�VL_S6l�H��紩�k3{Q�Z�vC���x�*����).;2K����
�$�����Z�l��C!%4�Q��掭�����v7[�R������b�����ԓ�c��f-�S>D�[yj�V
��k:�M��ײ�b���gL�	�z:^�L�ſ0}��/F�������gE������ۆ୛�V��8nw=3#Q���q��Hrj���X�]%�vj������E�L�{]�$)KV�xȄ�œ*��ޝ�j�'6](�8aM���{��Q�͗v 2)�p5w��VQ*nWu#k)����J��(M�D,
��+4��E���ƨ"b��V��-��n. ��WL�Z��Ľ4`'�n�`焸:�(bɜ%�1�+}춝`����̣qwӖ;���_ @Y��w^��L=p�s���'L�eS���W%�m;GAǁ��,ι�`�F��̌�4���ʀ�.�L��Wձgr���T�1a��q�T�uo�T�HV���������)ݫ��+��{R�Z ��^]nƮ�>
�wAO��f�z/.�͉�ށm��efr��u��Ú�4nTz*�"�p�P��Ы�,}����mIm����Kkw6�l>�K�̮S3B���8��e�a�씥oӊ�����v�H!ɃOl���T��.�"��7�B�
��tw�p�3�^���-�mbC�[�c�я'�����~npvw���K���D�ZrƢ�E���(��Y'!Wt����E[KV"�"��Q���b�Ȋ(�E�1`�A`��EEPV$b��,�������b�,P�P��P��UTEUADb�Z��b�QQ�r`�XbE��d�H�(1*TX���"���q����E��P+��"A��X�%�T��Z���b#���QX屌�**�`�dY��R�j*��+��YQH1F+`�Z�*��\�b�ĭ����X�TQD1#����X���E@Eb�!�AU��,���A��\j�+�Xe((��J�UX��
�,PYR�QTX��DA�ł��B��R���ƈ��Uq��\�Ke�,P[U���QZ�F�P�
��Er��b��U-�����`6��U�,�.5D�>O=��5���%�-R$aѦN�{)�b�a�� �A3a���n�j�(lE��	��{;_bYX��x��t#x��G�R�7[�/���I;�)��Ŷ4ެ%�Z�6�㬌Ȅ�x�h��&����iA���v̕oX���Ş�L�<%�M����K	�I.�/�����˭�F3�7jV3�������y}<ʥ��5׭�W�m����C�9�c}�ޭ���=W���԰�[������(��Ⱦ���K����T�o���V�x���F9�4Ç4��};[�z­J��~�N�:��C�,ʤ�J/��V�հ"�k�>���ֹ$o`��ˉ=~�&�of��aP�cmܴZ��V�s2{����%�X-D�T�:*�Yj��Po5����JY(�lݑz9�}��SG�{Po�D*���S	uI.��B��r�j���M�!�R�����B6ɛL۾Çj}#�`_=$��v��ThxoK��pM0�~�-���0�cٗ�U&��x���K��
ae�l���F�y}к|6�ʜRVw3f"e%��ڜ��^���<��q�ker���(�谤��tp�cT��E�kp�,�D�Qj���{Ii��{�'��T�V�t�;D�k���h<.�κ�'�]��*��VӚ�y�#+�XE�U���
Ӟ������SK!�%�s�~Nܹ4�N�U�*2q2�Ξ�=ȸD�ap�Ʈ�;�a�E�6a�V��Ξ��C�{�^Vc+�^6�j�ì��)��V	\�Q���w��D�pI8s�SN�nھ��Y8*6�U,�Ճ,؎�)u��)�����p\�q�ؽ1T��e�I��.(O'9�9҂??�����~��ʳ6����.7g.T�� y�sog;�|P�����lwl�#D΢z�>4at;��Cy���bⶾ��V<<�{�7L�^ٚU��;+��1��_��@��fo/l"�S�N7_F����v�']�4�VX�>��"�b�p����2&2���.�%�U�{UG]��?�ߊ��6)Θ�}��/����^��25��ZY/��|/�x�/K�cǴ�5���]�vۭ�WH��M��<��B�:}�-������K�kj�j��nR��X�i	�k#�Iئ�i��Ѽ����4����\�l7Z�6����$2�b�]�g��=Ŏ�a����,�ԍ�r	C���_E�@/s9���b��g.����o����juj�ӓs��Okr��h���PwSt]�Ssق� 6��ms��Zc
)g)�EhUy���+OB���;����l�H����Ж)>��I��R��M�E�^矦Zrs*p��+zz��;�t���=Za'�d�8Re��d+��w������sPr��Ғ�F]'�"�w�Or�G��젢��ݱ=�j�}�'<�"����q�8�Nk��x�Y�7"H����L��%}&mI��U�γS�v/���:�S�ޫ�R2�����,�^T@��`+)�,�G�uay��;p�#6Lk���EP"ߛ�_�Z��{�����D�ӏ8�DAr��YJ�(x��Bm=��
��G!�m����5Z�9�Is�ZZI�;��|~�������YJK,��<�3�޶'��������U�Wf\�$��М�V���J�.�l�T8�����Etz�5�Xk��������z걆ұq]t]�I]ҳ㼑��Ěކ���j^Gy��h5��{�q���{im�܅<`��t���n��L�%ҙ��V7�P��5��TW~��;sԡ��l�z�[�:�Znw�շܦ'Z T�;sS���jO<�}��#���'U��٭�"C�I�����Kׅ����Ϻ��N"i8.�g:>Of��`��˜dgm��[`��;�i�w9��^m`��Ϣ^�,o�n��6��i��>�2�,:�l�[|=��&)}�u�!s�P����qY3h����f��AC�M�B�P�~b���m��1�
W-�� �^\ s3+C(gn����d}y��M�V��K��{�84:���j] ��CDv�(U�b�JrF��&����F>姝�#�Z�T�a�}mL��jmg�y{�P�^�p>�o��@�Z2��)�dq��j�kܝf�6�u�T9J�WH1C����x9T`g4��[����|	7��ct�3��g�T~�Rk�)��f���M�Unpr�l�Ad7����J��	�EF�.� s��pN}$���Ep4�8���diDt���~կ\w����Pm,dM�Ò3׫|[�tX����YچE�(n�O)SoX�<jr������� �k��LaW��E_OK��Ohq;R�r �A1��!%�=�0PQ��@�kh�0�hv�t26����hѩRe;����ڵX��i9�u�C��q.:a7�yK�q�dY�wG6v������M^i�6B�m��ά]Qp����-�1���^�-�,��R%V*"�j�u��O��%���Nr\��}�����;e$�	Q@nJ���<�1������ˉ�>,MI@�<xP��M_9��8/�/�+RRDM�	��jB��o���g���:�f� T��2:H�)7��q�.�=]�u|2�ٳ=���S���2F�/qP��C��ϵ.��ƹ�W#bӻ�3�����'���!�C��m��{�>�-3��CW\��.��M��Rs7)�|��o+ޟn@w�E��dد�@5^����+������+��U7pn�c��<�i�Y2W��B5HU{�{g;�@�:Z���u��L��!�g/y^ς��u��!y2x�c睓�d��~M�@�u�=�ֈ��k{r/@4�z����)Pf|�g1lVK�/�=Ҳ��e	�gr�F5�<�[���?*���w[�+���+���շm��L�)�ේ=�!���/=^"'�Y��MK�R��x�F��>�
2''ny:w��RS�iZ/�����N6��-�L�_y@_�D@��o-:"�"�v6�(�]�Ռ��J*j���0��@����.ﱮK�e~��I6j��]_:�������~Z2��J�	����}r��Ɗ����uj�3�o>���CY;G���s���8�u9�ܝh����}�NT�
�i���Tt�����1��\�"���w�0����6���כn8�l�Ú}��'�T�t
x��M���$n}�������t��7m�1	��7�s[d��7��G���B\)D�X�["m�t�-ŗT�u�K6*��B��]g�QC���B�)�A�PA
b����_˶��I�i��{0-�Y�ۻ=k�ۻF�TV�:���u�VD��t�;j��iz���0���y-j��6���ZQ�뚀�ZV!Z��(��3>P�J�ܰ�V'e��2I!�8Uj�w��*�� ���{�Ε�8㝜)T�d��^����v��	��X�fG�=Ϻ$A���ė�Z\\Ť���e4gYd�Gv�MC��j�,(�6�� y�#��n�*
��޴o�*h��A0�_)�\,TY��K=-SP�g��<�=^ݶe��L�\>���mN�첺�\�1 4�X�N�b�����#h��|�P�Fr�
ȏ��H�jJ�쩃z��)�r�1;��o.T8�4[�e؈�f7`��r�'!z�>��>rb��4�N�*���4�lcӷA���·�����3��ml\��G����r޺�����0���q����ٯl�t+�+P����-��g+��m}|����`h}��4��#R�n�j�9������D�eNj��S�+�ɩ��J�@�[7��ٝD�X�]�,��60�[��<e�v��{]�Rw젋u��X�s�cjE��{%M��`Z'ꟺ[���>��+�(�	�EF�V�xn��[%���U�_��c���-�՗���ڪ:7VT��s�Kup$���2in|���u�"�6�s�b/%�>c�`�J٬N#�tp�F4�o��}��)�k���<Z&g��1R�#�&����F+��dkX��&
�D��Q�*;�P60\�csKIt�����K�Mq�:�����ݕG6�$#�MEk���3�Xd0<�Q&��=����qѬ*y(s����7����0J]�}8�� �?��jt|��Vח������A���D���䊊h�s��g���W۴$=+��^��:�g�3�;Mf�eO2N-���C�do:uE:�bWѓ6���*ÂgY��O�ai�ԏ���'����ܜ}],�"��&J�2p�W�����8�z��>�<y/b�>Q�m{��c���v�-x��� �Ӭ]PVӭ*­�G�1�eso�Gc�����L�رs��۾�[w��b���ƥ4�O.=R�)sx73����]�[#iI���Ӻ#��ڨ8-bys%񢹼�)홹V�r.;o�,�㌺��H�
����"�n-����p�]a����}�陚ܵ{l�{�,��$�F���%8$|e�w��߹�WR�JK,�a晘�\N�v�}���f�Ǝ��I2�Xmىz��hs������jetgU����B�r8�l��k�������ܱ�,j�'2�#a9����E���$�O���%Y/��D�b���)�>cfZb���k��72Ő?�r�<K��>F��s��
��u�cRg.�7Ѭ�KV\��~�t�NPdm{eS���U�=�a�ۙ�0q�̌��,���*&���ۅ�c��E�'��'���f�_V��uf3�F+�,�hQ�
�"t�5��\�1�^\hU�W�GL&S63� �+�*i��w�Ⴒcl�������{d��`z<zL`6�9�U�D6��3�9����2�ePB� �6�//n)�=���lj>õ�M��F�*ӗ}��t���#��������Ekmi�*U�ܲ�ŗ;�� �U���U���W����-eZ��#7�-�Ob�4NNL�wz�\�b�+F�p�Ԭ��)N��^�O�[O����KDٸ�n';��v�c�%.�-Wp��-.aR�,��ZT�F:���Am��U1*�2�P��E5�(o�]�Q�xW�%7���r�^ה���;����L�7���P�\0�8id��F{�?\�E?��	��zz�4�C�bfz{��?X�C��*	��Ox�{s_���o�r���%��"�K	`�ԍ.��.���-��W)��K��M����h6�Q�W�N����L�p�Թr �A1��!$��[���v��������FI���d��=էlv]��	��ʇ"u'�j��]��'aZ2Ie��ݡ�`+�O���.5��ذ�<����<,�S%�$�W�z�ݵb�S�=]�	���k�d�X��B_�(sU9�����P�i��{1���3�G�38�ߝ���7�?g�g��v����(-3g�u���PT�3rBt�v�� ������c�&����v+��3���u�Z09_�W/̯��5V�Z#�<�ƅ�Y�į]�U�y���"���쏁]ҁϷ�� oX'F!3���3���R��*�!�b;����^����A���a��謃�鎓c�|��-Pc� ���rhj��'�h1�~w���Q8�fSj��RQ�T#�޹`�� ��vQ���C(�;9��v4/�ƶ�f���ږ��[ȥ.�RU�%��ӗ�z	�S�pʳ�7���7�w�-�Z�܋�Ng�'`�6�eR�]c�s�v��>��.e?+��nXq�jN������^�_o��p�פ�P:#;�^.]*�BeΫ=sp�AŊ�fNz��af�d�C�����ݖ'�ׇƮ>�`�L�,(��y+ȗ�� Y�[D�ye�-�L�_(��o^��q���]�5����ۻ�o铥��B�T�^]��%��4
�2���H��uY_�J,n�݋w$ؾޖ�p�/�&��Rv��N�)ӁNj̃!�L�i���\d�r��r1{±s�/{�4��VטHRs�Rڥ�	Y�}�Äi��J0]�%�b�Z��Ys��Yq���͎�H�t�#�[=�X�h��if�m�}�^�,/���*�p�8�E?F#\����G~�`x�y%�*PӡG�Y��ab��zPf�!��u�>wI�u��n�&�t~*6	#{���������[&j�鵤_��HG�!��l����[���9�G2A���ezn`J�o:k&^Hf�݁��𽑛�	��[[�'�M>�ۣ?y�Ȱ��S����oѣ��r����"l��~���I�ʛ��U�p͝��[�8h��O�1槾�!��.�1�̗d�m2n�=x����]�T0��\�*M��p�wiX��,-�xU�%+h��X�́
4�h�&�X��]�w\|c�ˑ���n�$��H��<���B7��Q�ȕx:�u��le�,ͺwJ�2C������<n�b=��r[0'�H���;j�s�|9�p��̞�J��*�M��=�f���;�z�H��)7��Q���F;Y�8[4��5�&mc �\&%��Mk�gp 8��r�ǳ��ỳ�s��ҳ�^ȶof�X'�w�Ʈ�����g;�9�t�<��3y3>��2��B��|���`����o�Bo]rS�v�6�k�Dm P��Q͒J��iN�O��3��j�1yT��_��LAn@�%�o���j�=�����"�n�Ѩ���t*V/��w���4&e�-��S'>+w��fN>�+�I���7�q[B����w�Ș�w)��ظZ'�k;�iu�#K���:�p+���7t�r��\�7.ŗ=ʴ�J_B�U�𧈔��RNS��{�F[2<�;,��f�æ�D�HLC�c(��\�k�S���!�X��GfU�S���B��ż��g��`N���A���*˙&�|��#��$�����`d��,�'7!��#���mK�׷v��V����L�,;r=,IF�h��.�jЅkX�1�2�<�M���Ah���k�)ҲЧ2�N�IU%�p4��2��>�>�����߂^k��Yr��n0�{���Lۨ��Q����2��=�y�W��6�׾��\�3{����.�V����"����y�	]�������ȩ>�=��x�����Õϱ���5�}Pu��{�{}�3��Q��;�~�	��m���2��t uj�D�����Alz��8����O*��X��=�#� �zqZ��h����GqT��czgYM�@�2:-Кɽ{jU�kZ/;*^� �E±��$�������l��M*:[J��N�u�A�K���|՞[�2ۻ�f[���Iw��v����\C��nJ׫�;�kT�蒣�Ac|�+r��<�MviWܶovglݿC���Vo:=Үh�w�����J���gu�;�'�/��#�*9�{l�]�>rڷoy�KN���#�hpx��^���3ʒ�#�N~-�0ڊ5t=.�ŏ�׎�U�� �4J{3q[�2�E���a���m��K��j����i�b��AxV���y 5���u����cnPb:F䂗ftȵ�i����T�)�^sB�ۂwt���V9�h	=1U�@��f�r�G�ߦ/���~u\���H��((��%�0.aT`�E"�+q��q�(�
,�"�ɉS1-AƤU�F��es3(�es���e2�T�-��D�e1���1��m�PDW-��	-,Q��U�����U��RUcl��2U�KB��D����\�P��EUEA2ªcr�Kh��V1UR"�!11$J�XUq�Ui1�J�ZE�9B�EEQE��Q�����4j���@QTb�DD1��e��VҨ��U��e�.%)�+�*�YX��"�*�Z�#�Ɔ%T�e%QUX�V*DLK��F,T`�DX���#&5[V(�D�"fY���Q�4�R"�F1Bc(�+�����"�)e+r¨�)I��TLedP\h�(�E2�P���(#EKJ$P�UEJ�!U�������̓Z�+e��q=�W�2����a�E(��Ruw')�p罕7�!jڏ"��f���hC��'��*����:���$�9�''/��W�X 򮦌�,��b�P�+�v���m�@C�`82><o���]2vsh����9s�A��ђ�yj���?NV�A廖'|c��(�߽'WQ�flq)Ó�CC�9�����Ԭ�Ee�Nejr�U��}W�	ʜ��ra���vt���x)q
j�ݰ1�(�y��N��oA��-qsV���zF����j2k�f�V�X��&s'� �х��N��x��O�pe3�!���ӂ��`���v�t2ō���nv��O�8�| }7뿢�Ҏپ��Wi����ޖ�ι�ig8k���>~=`S�,�zy,�����,O�[�O�E����j�p~�}p��ߦ�دWI�$i4�PwQ�~	B���cǖ�����=}C���$��{���g�����Ǝ�>��:}���_Q5	Z[�%�U�'u�Vx�g9��{�;ozK�oƸpf"�PM��n�<��
l��@S�§7�Q�Lm��*m�N�"]T�9��>��yg���ov��Z�^l�*��[��8|�;�)9����*�{�q;��s�:;ˍ>�O�6k��:4���]
|�Ob��Na�S��.cm9���d�d�ol�˜ѽC�‡���,� ���Ti!���񓹽>�.�vU9� T�{<��Y0��(wX���/O�'ءKL�dB�{�m�y�=W�U{�Ѯ�|�RqH�����ܴg3�e��
*�ݰ�U�'�����U�������xQ��V��$�Դ�(i�1B����d�7�r;���l�W��@颏D�bW����!o��c����EJ 7�'�H�����q�޼=<o�ON�US3m�`�H��r`�����N����=
q_�De�����J�N;N�F�V"�3�q�k�|�^b�(�)��U�����!q�WR��iIe�PՇ�㯭�;��t���!���P}��HJI��vb^��a҉>5:�q�S�L�����{�5*��b9$�O�]�����ܰ�X�����"XPc�H���]�0���%��W�����tK�eͷ�_{�!2���F�7��ˌ�m��[`%�Ѝ1
�jP�^J��y�gx=�^pC;�s�Yg0��G�����Ϭ��,<������߈��;P���@����&oR�m�b.ʫ��Z�늤������d�����dX�_L#�e�j�
�s�c�HɭQ��fˍ���;yѥLnk���n��b��ֲr��)/�Ϩu���H;�qo\=q�7�]��2V7u57q���B�e�v�\��= �b��$4���/�U��υ/�Z����ޕ)Vy�#}o��}6c#��l4�2�y��;�ꎍ�2�&�`�����<޷M��Y��cg��i��U�0�3��ə�6�9�w~孽�o�`�K.���W螁��-U���ߢwy����Ы��d��s�6���#x�N]��8��Y��Z;���z�DO4��j�,�kQ��Ғ���-���� 2*�u������(/���P1�H�ӊ��9�p/��]�����5�Tn�(��&�<���k����afW���s>ޣ��s�6{d��7��N�Sb�hN,�Eñ�KT1$p���[�\�VO�ʲN��ɯ`��Sq�JeC�����M�)0/�3a���:��{�J	��$��=幀�����=W���JH����03�������룏�f8�ȣt�=�����lH��:%�A"�L���s�-��ӡ�kB�WK��pL`��N�U�\8ǝ癫 Tm*������h{A��nE�~>��̢����U�V���+����'܁=l2�I�%�1W.{Z�|���!�G���-A��;�r/i�<�.K	K9����a� ��k:܏��|��[��2�P�⮥����9�.e��;ڏ$��_W�@v"�j����d�,^�/ej���R�r��5,֌�t^���z��Ί�4J�������Ag�e���x/�\GS�X��ՅN\�8b�udͷ�s�c.�P�6Ku`�톆D��}�^=KE!�-���W/̴`{[�h��ik�	��	���I!�[7�ʥ�鈛,`�k��:�12�c�39{ək��>̊j���"���t*��\�`W��wގ���z��]~'p+��Ӷ�6���S�����U���='�l36;rg��[��������}���X{�v�U�1%]��f�Rm���i�H�a�4R%����{�c���CS�;���1ѽN�X�E-�5>�Kg�.�ZX,�t&.�yV_��ˡڼ`>D@�޽��M ����un��meꡯ�<
5�齛���萍��<R�7�M�d�����W�X8}��բ�4�um;��T��YI��J�VuB,"�V��>WJ$��;l��ͽ�b�񒷇�^K�1�7�Ǒ�+Q�K��~��<��dZ����T�;טḮ�YNd�Fg����E,h5��.n�M���w� ����"j_4r@*�x����b�j�y:sp�I�t)r��:��w�݅%Y�,��-��<��N��^n�w��^��^��]������p�hER�c�Bge!�Q�x{�c��b�dx6��ԩ�5K�>>y��,v4eڴ�;j��iz����(��N����o[t�a�0C��@�fx\���ʑ�*�̷��eg�ʱ�:2��y݉K���`�o��EO0j" uz@�d�h���&j߽6����E�������3L~}���i��o�\�/��݇ҥ��%E�Jh�e�#{X��^;]G��@��Ǿ�ꃽbc��Cz��f
#N%Qt�42���9x(3_}��%�^ZF,���u�!��S�N�����[p�d��aP뚋	+s/|���X��b����W#A�B�ܦ6���Q��i���I�*%3`(i+˕!M7n ��9�����oA�K��a���)���.8�Z}�t�1�k��%���9��0��M�����1f>��l�n�0��������v��냖]h��\߳s�-~���u���o�_En,87���k�:
���^�����=Ԫ'C��:zW�א-�1d�d<�@Fa��D��C���q-��nsֵ�TG6dӧ�t��z�E�Mܵf�"��$2�tzpn;|����L]���;i����{!�rt�U���QV��\#S�%�ǝ�:B��\$xY�B+xv���)��5���u>�}�i����6/cgwg�uY�RFNҙ�^�1x��H��C�����n�b�����	���v�:٣/���V��0UZ��+��p�Q���קO�s��}Do��.�o�]TFS�D�[K�����6��3}P����LE�U�
r��a��%F��	��V���KڽNR��!_�`���
[	w��oN\�ޫ�Q�����̘}}�;�t���=Zt�ĶHr��霹������җD��Iȯ�O���Z�z��/g3�gc
*��:s�;��ܭ��J|�Wgi���+
۔I�W��/←����7���L@��Nex6wT�v\��y�~�#�#���ue�/	�jDp$ɟ&F���FP?w���ۯ�yh�2��R��;Z_ZO�@u<OC���3}~!P[w�E��Z" ��'[�)_Ԕ8����:��;���sJ֔�B���Ώ��}Ϫ%ě3u����!q�WR�"iI`�Nw2�N�s��ט<`S 3��2.�pp�b_�V@ǹ�����I���'y��}r�^ʗ2�RƆ�������LO"��2ӧ�w����]q���4r���Ú�	�')�Ɲ�`I��]"|�_�A�-��1�Fn�K���Sq��+>�8�Wm�{\�ٯil�۳�͸�t�cbӻyUk��Y%��.�t>���v�οz3������eAO|�I�F{��}ރ]^����n	6+�a�y���/��#�"������q���Ł���K�3�F��r�HWU�Q�zc�x���*�
5;7}����~�*���ڭ���Q�c�3`t��!�&ٻ��;��E�l����,���unk5�s\^� ψ��^jyq㲻�pK ���'�Ӹ�ާ�`)��Ъ�l4�2�}ή�sz��GN��z���|�?v�˓�5�:���˅��l>${��מd�y�=U~��M���΍�\�V̪t��DFF>A�8�µi��L�s�Jn�g 鰄^�QC������t���-��Esс2*̷�������W9r�K�p��"�hv�����r���E�yAy��7.8ta�*�ږ�����{�)�9�f3�}���0zؖH��zKB)���Wxu6:���Ѯja�a�%��}�*��	X��Sz��卖⫵�R܏S�tz�8�wRy��L�gٵ��s{������c�Ţ�{��7%��Z^3$�=w�e�S�n�^ m�������MUӝi;;|�;1���I\N5�Ɉ�A�0���@�yS�]/�bZ�(�/䰐wR6�Ț_oc����=8������AaH��~�"�K�H��q�r�+�2P	�P %`7iV���o��/<-�$��5}<��o�t������َ.,��79��P�A��Ѳs���ʾrnG��0�����Ѩ�=�*c�������L!��/-����4ڽ���pO�;��w���Xs�1��H��	��kg>Ի�r��G����/�+��w��3L{�9��1a�>�PY��x�e��5u�S�اQ���T�oZo�8����5e�]]s7/ܫ��ŏjDY9��R�HC����?���*��62�N�/�vE������wT�G�}���@t�oK^@ްOV���]1WBx�W�٠[�ʸ�:��k�޵h���jz6�м��6���w'yOֈ�-onE�s:}��T���0Sْ��[�o!��(}�x���
0�B��%���Ҁ��}�����	�;=�A���꿕�T;��m32��!d���3��5��N��.?�[u�S��)OZ��6��Վr�h|t�CRǤN�{Q��� � �o�Bf�1�@JiI�|��<_3m+y��9X+׻�����]�e6eN�Í^m1��^8�E��K�>��h�ha��o%��������hj�|��
Қ|'{n��i�ê�Jqt\>�1�x�*�/8}`��l
}KlS�W�P��/7�y7X'qy�,��v����DɨT97aB�L���;2h!����]7�K�����w{x!�4S��,|�]$QĘ��qy���O��^ճ��X�	gX�	�{��9�5���j\t��v^�@c]Bu���^�����P��x��:u%�P��`��1tX��5�p�i��t�,�ow��s���o3���4e.e�<�|<�DĪ]�����b�Sޏ���~�����qȮ�#�w:L�!��){�G��L�-�=iuD��/yȚ�������,�z����hI@����f���kH���^\����J
c�m�vSϢ��ᄭ`�Vrȱ�Ĕ_��;�d��'O���a��`��Rm��졉��7��IP���xsw�Y���Y�xs�A�I��,��cG���_��ϯ\��8�H�gi[��k���XG[e�Λ	�c�bIw��R�)vf+u)pWBJ{v�tCt�wͬ�ʑ[e5�H}�A8��jC��C��U��Ѱ5�p)��Hܡ�ݒ�9������,P+���专�WV���Ǔ�{3}'7*mp�ݖ$4��m�&z��oCCӓ^@���}J�L����C������KW_pQ1�9��N83�+˜����ۈ�]��W��ܡ���n�[���k��"\��B��M��?��Y��_a�^չQ�W�Q����u�`>4au�t�n;�/�&�f���d�1�1��XV�.��ac§��]��{%����D�S�n�>���]����班zN-�m�������boܳ񉓟�<A���������U�F[�
m󠭮���a�I(�=�N,��9�������0؋�z���_+���+��-�(��e�����A[���%QD��C��o��|������b��Z)�wSt]�P>]�A��R�e��t�ٶ4{�l���綏"}��J�ǬuK��*Oyf��
�×ڕ���\SV�Z�.�X/���S�/��g�o�	�}a����q�R�1�b�@ԕVla$����+=5�����x
NEb��"�w�Or��g���W�`�8����V��:��iL�9�g�ͺ{�ؒ�#Jd ;3g{�7ۢ�W�JV�R��L��ɪ����Ϊ�x�ȭ�4U �p�:�ܛ�<�ZU�=u�Jw� ߝ�4#{�m^-*��i�+�ԓ�����)_/N����3l��G�cE�O�cI�Xİ�5l�����Ag0=F�;�U��pTݻ)^6���)MM���p�<��T���������|��RT[���oZ!mIݴ�\�������������_;�'���+���~8e�Rgh<���� /:�㭠��	�,7���,r��Ǫ	'���=F�4���/d��Uz��:���{)V�g4v��F2��	��e��}�ś1ww^`�՞��F����l��G��ߌ�C���[��q��*8�7�	���h4��|y�M��#�u�li�ծT�D9�yCs�esu���M;�ӛ�m#�B�v��#��Ui���c$fu�z�H��b��~���7Pd�����qG3N%7�3�_��F]�]ٱ�wkd(5�>���r�\wI���py���X��w
锯l1)JHtk�쥵���Νe�o��{�P����*u�F���w����\�yl��9�Z6o��"/�2��g;�^�F�����Y���Gw]��ޕª]������������զ'�s#�ԄhUՊ��k-��zӽ;�Dڔ,N�N]r��r�м���2�b��8w���̳J����.[#�ĭ&j<\4.r\ƬYV��|i�.�H�`�e`ѝ���8���A�;�9^���8\��'��i�t�s��:�ꇥ��2h�r	���G�ym�O{.����H�%��Nt9�{��9 )
~~L(3և��ح�c�3�.�c\�oF��#�W6��H�.�Y���2�S��ӭ�s7����S5xj";ؗI�:�pi��x9�`�]{�R��۹X�@L.� �m�Fv�*��s��n�VWJ�u]�X�%��E�����?t�2���p��^�dС�T��Zα�˰�=/ob��/dG�x��g~��o/1�BIWqz�f���6�uY�y��mjt�E��{�X���yD2���eӓ�oTg�v�|�A�,��y8�`I���绫vT�RffѱՊ�w��X��F���N�ɑlo85Z�a7A��ۣ4�cOV��������ur�٘B�3������s�^�M�L�{ !aqz�
�M��;��W0�;Buonj
 �\��Ԛe�ͦdkj�k�D+�uXMQf� 66un�݊�3��%Rkā��һ�i!�S����S����� #d@r�J���<ڬeu,�RIZ�a��vhnȺe�ѳ���Θ�fn<��Ɨ6��G���.�Dy���Ḷ���z�M +���m�[4(�ɤM�1�y�Ф�솝pΎ�Y�;�Dd������\�gwH��e�����λ���_@P_|}@}�V,R
J��ej������Q��PUUH��(�)��"��,T2�QQR)�E"*((�1b���(�m�QEEEF���V�QUdj6�UX��aX���*�Q\B��fa��PX�bV�U*R��1����
�(��ȸ����`�kUb����b1c ��"�jc��(��",EVTRVܹ1 �0U"��(1EEĬb
���-eAc����QVRRҪ�iPUb�`�T�hW"ŋX"����!F("1PTATYH�q�A�PUDX?c�;+�Vb�Yy$�$�!�%��MuŒ�{-ڢNlw�Ff'�Ĳګ���5�<'lE�����u
�c���b4�r�\�N_
���(����
@���s��%d`6�ƍu���G�+a��������ޱW՗qNK#x"d��'�Jb�O�5������d���(l�v6q���+L<�(s�wP�Wψ\����
q\D���唥=��z�^4�^�Pd�6Y�Fg9��CetP�s�q&���?rW�d~ԯ�Rf�[̘��3��<��Π=���R5��tޛ5!)&\���ۈ�J&6-;��-\A���[��=�{:�ܿ#`�^��C.vh�5��YPV=���H��=����u��Ķ�w���o�X�'��K�ԕ�9`��v�;4ma�S�\W��ϟ[w���ѣ`{���ߛ�=+��6��]�p"td�c^UZ�㥫bm�}_0��/T~K/��_�,(t����.���ʠL��W9�5�= �:���\��E�ʾOK��������ʾ�um��Ȕ�W�7q�]���%A�\��ި�߱{>��`�0��5�w�U.�hn�%�{�7f�\�&Rם(�q�Ɠ�K����2OmT��{6돴����'���/syrc���?s��>��d�C�m��
�CK]O�������{S���-MuhV�놖\ʘoU�R�iV}ƲU��#jA`�;�ZP56\-V髵w�d���s1�ݧ;N�ܛy�͜��ie��&�b�U:�����~KA�Q��/URbΛE��*ӗ|<�00���K���t��U��0�����134��[�(4;U�W��W�A�?��.�v*��h"��{�$ڂb�x��zW�zk�Q�P���&��X��IhAbw@�!�^G���"�h��v�TriAU}���&;g�(����[�cX���(�,%����H�˜��#��yq��I3u��՛����o�/.\��b�����g�G\��0!(�BU��A�WkK�LbmJ]�@=i�*��k�h�b��ϴ�z���]�`������J�������q���s�`�afP4P��12��XI�S�����9�<�Ü7E%ֻٞޛ"qb��P,�^���$�$�fui�欿��8��T%��N]�Y�K�l�k:B���Y5Y����HYᲫܔoǩ~� 9_?�yʯ�O�CW\Gi?e��G	Ŷ���S}9�A�>��ɾ�4�H�I�4���Y`�yR��.�a^y�aw�1���"/����r�ښ���31������l�}M�v��]#j�u�n���d�9b��P�S�4Y�Y2˱�h�2A}�4�*G�I��}�L]�|V���R Ί�]73s�N��	���T&��x�-�6����jo��.�*Vi��WF�U�}�kn-�{3��j�M��F����%�_oK^@ްN��0�"���|wjz�<�7�rt�K�Ͼ�=ō�|;:�4��絎S���KkG��"̹�k�P΁�8]�a���lB�bj��K���z�Q�jN%����ˏM�o��l[�bt�Z�;�Ts��i�-�'�p�D<+�;c�����zX�Jt8�5�"2���s�Q&�����c�O�Og
��w.�,C0*'Gw՗�<�˪��� �����ĥ�>��ç�dY7�.�\"�v6�(�/��NN̛�Bb���i�*2F�*��;-o\��X�����"ĨR�E�v��7jj�ψ|��I0u�Б���}�v�=,蹽�cQ��O̚�?��&����`�)��t!Mըz!+0�a)�!&m�[fb��&�M?{ZՐX<�(z�1��oN�}r�!j]q��G��yY�b�����p�\���ħ_jc!^U��� <m� $�I���6*�bo$�V�����i�[�t�v��7��W�aݳ�^8;7+��-hn�RDL�o3�{&E��v��;�V�m�-d(�]tf�l����n
1I._(σ��k]�F�������z�Ӥ�mG5� �K����	��9H��#ƞwX���cO�~��7�z_uk�&�j�UM�Q��P�P�+2�]c�$�@�J���iFO�00*v������Tk�*����6.����u���U�E�J��4d����b�j�~�Gz:fת��G_S|��1���&(����n��f�NO܆��A�I0��MC�P�v'#AZn��z+i!5T��㵚g��0I+��}ɀ�ކ��	Ζ 5�o��E3�3�/_^7k2��tR.ӗ6d1D��ʔgrr�ӎ��]�	q1:�&�ޠO�ᝧ��g������M9ff��T0'G���>�>䮥� �[�z쉜���'Y�Ɲ�4�:�Y��hF�R�M�+!��;z3�<6�`�=㍭U�q�����؁�Va�.[Iue�Wn*:/Z�9�g�5�^d�;���y�kK����o�:�;
��d���_Iьur!���xw:"��g/9�a����u�~2����M�wNö|A�v�M�p	S	z8�7��t8��Ső��+=��.G�zg`[����b��v9���ZRi�J��(furo���4zd��9�|����~�HЕ.����R�X.�h�V��PAgnm�GU��	ӕ�ҍ��[W;5��+
'�2.s�k�(k�`�]J��<5���Çs���Ȳ5�b_� �{�1���*��$ґ����� ���]��LEꠛ�����k=�J��	���e���'���ѷ[i֝i�	Y��}C.��V.J��0�����B����k<���=�̑��O"}��y�/=pE����jU'"�I�z�e�ק�{9�C
܄RzMgd�ؾ��8�+�9-&p �l��Vk$�԰�
Ct�U7��H�Sʰ�/����e!ʤƶl8&u�D1׽b�ue�^�֤EpD�A2q��#���s��Y�����������8;�o8�3�*;[��~�Nߝ��#|��ҜS����x_sm�t���[=r�T�����[R�@t�L�1���q��\���t�ۀ[1�w^��mO�"DC
zM�r�F܄��pԅ�L�vb^��~����(r������Vq�M˝1�#���)�L��ֻ4����1��MeAY��j��H��c�H�����x��[~+g�g��%-�֪����8�`"]�������zG�D<�����J�'@�m��N�tLv�/���Y��
�R��ى;�&��ƪ����6��:��]{�[����]�a����7&�\�*�t����mc�2�w�����27���pa���#)��~pGM�
f�;n�ˎ����ʇ:ޟvsպ��_&�d�d��!�ߐ���t�s��*��:Z�&�����K�,:���پ}C���f8�z���.VeE3ٛ F�20.b˞sNims\^� �>#�����=�k}Ǹ��d�6NGK꾴T�@���@�]���Tu��\3�ፄ=ӽ5�Dct��t̓��s$��M�p��P�s��m��.��{SR:��Q�W�;���^��tF�5:�Y�v��^�#6��)ZS��,��aAqz�R���*yIc6T��]C�G�<�~�%J�33�u�j�[;�[���F&f��J�ސ��^��z'�A�7'a��qC�#MY��=INz�m��\�wJY����Mr*6)B�`��hze�M�c,פ��c��=˯y�S���2)���1�T9��'�(��X�s��ga��(��b�|z9��&\2zZ]+��W��Z[��+��c@kz���Kqi;hq;R�|�2~^����^@M�Iawq�i�n'��_<x�I�r���z�T�Y���Ժ~��w$E�Q�-(�ļL��.q{�km2]��ٜۋH.m����	z�4M��X��K��(�[Q
�8[{��������f)/�n�̼�)\��e>2�������7^���CI-[�R�r��2���g�b��?-�-������FO_T�蜽;��� �##�(x�@����a*N���\x�6_��W����[מ�z�kr��`�x�S*_�K �զ�S���8��bf��K5�W�Aiޖ����ɒ��ƹ�dhN�y(ߏR�Q�A��r��V�<��aq��ra�7�'9��T���@'hT3�X���ƆX���5�^=K|m���1��*�7bw勑��#z��L̹gk��r��[���c��鈛iX5�-yk��&.좑���2\��b�ǽ�^TึV�L+�B�Tg������@��M�ֈ�.r�����~D�cQ�yY�_�*Plӫ�S�/T�ϵ��J�2���ǧ8���H�s2�*��YK�ީ;�h����:}hQ�Hw����!��B���X��\Y3]�j�4���#�W{�8h_?^�](X,�wTís[�����Eʵ��׷r�_�{��=�*園�r�<�ed��6�^&(�oȷ�;I��oW��<0�cnB3������Rm-.#x�r�ٸM��x;����z��J�X!���W�d�YTk���&�f3c�)��%��n*Wv� ��f.d9�3��KB[������gc���U��s%�&���٫��DC`��3��C|�*��k�m!�V)�o��;�R:}/���7ۖ��}}|6�:ys�����uB,ȳU�n9�.T���z4*��3�	[	q0:�͜u���ˁ~�P�{�MN�s&;�C�G�#N��;��v������jKy1���'�&8�m���˘�����{�Nƌ=�K9�Tk��ok]���0�*(̬��h`/�%9H��L�y�bԹcO�Q��B�<}�@��!��f����a�qp��Z��I"2��99�""3��+|� �ZW{坥m�=$�<��;�%v�����K�/�IQF��$ F��A�s�Y����7k��l3�II�,;ip�C�`8�w��42r~�7�
ֶ��e+�{[���d:�e-y.��v�l�v��m�b1���%r]�L�X��C~~[�*2w�k8g���*k�4X�)s(x�[�dOP���H�<N������~7#����\�7�Z+�3��X�|���6?A��d��R\3�g�_�ݓ R��ar���K�*��xÃ�̥�@��-��S��Ț��ե�V����+f��$r�D�{Y�p���R`k6���}%w��]s�Wi�3{}�I̓��&M�&P����*r�^�2σea�gX[#*�-��<��C��52{�\�-߳�fv��l��v�&����b�q]�C�U�;�{Yt�0�x�6�T���/OWu�aκ)��隹.H���w���>�YSע�U�^.��kò��%�e*�cĤq�S��M![t��t�U�fnЮ��*i�)���-U�L3��/%��OY|DMi��cw:b��vX��cv]�B��J"����2�o�]��aEƐ��7Ý��2+��Z���m_�b���q��tL5���	sO�w��1��n�ۧ�0�(�1��a���u$f��)��������H@���b2�V��@D�J�Q�j����D(��ؑT��+[z���$�����.-c��Kʗ,� 0{P�IȮ��"����Or���XC�t����i8[�Fl\�`r�.n�v���a�x��D�� ޒ�(i�*2S�g�E>ѧ�v��rWQ��s7�ѺU�Άj`Px^�}��~�֤E�%��
��)�������pe5("���2u�ខ���^�f�S�l���p���c|i¯Y|��#�ɲpɎS/���\[sP6/c�W=�חP74���ݍ)8x,�x�b.u�+h�Bx;�rT�"v�+y&um�&��]���[k����7K+^�YbwV&�}_����:�x����J����c8n�c��K�˅T"�@7�D���3:��=�Y.��qx}XPc�Tj����3����v�^���n�ǹ�k��s��l$�y��7����3\���y4��	Z�ƫ�r�V]���
	� �ݘ��͸���{۠FcMZ��垸ݦc�fS�~�v�WGak�_9������S�ϰ-ݩ&���x�S�tR�P͝���H���I��#_Լ�}�_s�k����_�4k��ς�wLcR����{r^���)^���z籠i�w9����C;ib���-[l��aG�^*��@8a��Kǲ?d��L������-�;P�3�o,��;XA��Yqa�3���K�I���]�sU��mK:��`�"wi�p�xaF�]����2�}ή<�{�T�#c�y���Z���׮,T���\>P�_f�#�g�����c�i�ӻ�-m��ҽ"í�}����T�Q���yan��_Å!Gp�:�к�L|�8o�U}��	'���$��@�$���$ I,	!I� IO�H@����$�$�	'��IO�@�$���$ I?�	!I�B���$��B��@�$����$���H@�xB��@�$��H@�{H@���d�Me�}���~�Ae�����v@�������� (*�JQP�R
A@P��� PDH�T JJ  ��T)I J<�A@�$��U"��QT�R ��UR)(P��"R�IA
�%P���r�UD�IQQU}�($��T����J�)����$%P��J����U�{qR   �"�*��՘օA[kYJ�R��"T�&�*�+)�kSFPY�ԥl���J�����(  k�JDV��FL�A[)�UA �-��2�*�acTPڍ�0��
J���Tb�TU)��TD8 �+�)a����Hh�Ѥ���P
�m����ґdcX���i[I�L��ҠUH��Qx  ۴U`��ZmQZ���q[5��Q�
)E��E
�qҊ(QJ7#�E�\s��E(@g, �A8���PJ��(�  ��P�[#ڨ�wFn��E�ZY�t3��[��mn�m;�j\���a���]Uݺq�5�t��[
U�l�������á*�P�RTA �  {�U�=u�\�������1��:j�4��uwv�:ڪ���f�\]��3��Q���lٵ���uL��t]�w(�5C]m�B*�UDP�  �{b���j�G[�,e�[�Wws�i��kE�j`l`)��j�;kU�L˺� ݪ壪֖(3�qJJ�B�%QJQx  �y�u�m&Xj�m����h(�mk��Ձ50�`��Qtԧ(��n�ka�mR��Tj�t]��]6��]j�U*)R�  y�z����ֵ̭�kw0��.n�ͪR�`�N���K�۪i�1�\Eڛ-ck�M&�û]��X�R�hԥA(RT*!�  pU���۰\-u��3UUKM`���u��uVk!GVr�U݊�U���ض�S��t:;�Қ�Ќ�R�xIQ�T"y�))��� M  �{C
R��2�&@0��2&I�Jx��hL� yL�C1B)� �EQ��@�4ɀ��j��	�UP �     i$j�H�S��ښz�T����H�׬ݦz@��t�Nt�'(��F1���i�uwV�)B//;5��~~�@������ H���IBM$� H!?�0 �0������4:��H�0�P 	%C�$�B ORK2��T%H	v���;����u4�������  D;��՗��̱���O�O��Ӱ�P�J"��ßO�5�����tw�e����r�A[Lj5��+5��h���G^6���Oq�1�70�	�d��ٽV���K��ʱ62A�`&;LV��*Ee*eՆ�T�e37S���6KB-ź��P��4�v�c)\W�-f԰�f���˰#&�u���ZlR�a�y����MM�m�n��\wIbldˎԫ�c2[�4�N*�'�
�N��حtjd�jݺB_L�J]c[X�jˍd���NnMR�X֨����Yb,���r�57iX�Z�h�Օ���e/�|�u�u�+G�	+���a�[���Z[�	@j��1�lˬ�r��{�K1Z�Ead��)�R�����&9��{{nBv��6`*X3(m�kh�;Pj	��i�l��{[RBԊ�h��Z�3����Y #I�t��˺���YotR�ۧ�*T�t&m�������T:OqM
-�����wj��� ����_؅�MU�s*4����oo*�P�s4��L���d��Bf��X?nIE�5|�̫9�(�h��� �؃���ũ{���xu��)Q�:�K��"���8u���o[�4�����#h��}ėF���Y&�u5�U��U�Q�$ ё`9b0a-Ls>or^Q;U��I�l`�p݄�mbo�@��5W>�.k�csi�e�ًl�jy[/��z��W	
=[7�E����u��M��sᨑ-�Sۘ����hͶ�6]�ҎhJЭn�{�呔��o�w�+5���yw��Ym*Mml��wa,�R�Z���iff!�2ʓf 	��f�:�Ĳ*x�����үj�h��*��l;Gl�!�7ԭj��Z1E!ڴrU���X.0�ʫ��(m�*�㬗X-��,���	�6�wv:[U���b��ħ�����;V��[����.��Dh�X��(Q���(�2���n�@=���:ӗ�m�K�`?	�b��<�8���nP�;�s� ��v���kڃ�|���w�9�.�=X�6)�Z��8�i��Ӡ���m�Zpi�Y�vN�K�7��ϖ�K\�1Y�n*�Qq[��FՍܬ$/g֒r�74mL�Iy��� �q�4�bR���h�ț���::���%�c+x���ѡ	��m��Hi8ګ"�e:x���i�a=�n�`-%�se��Alԫv�i�VM�%�5+@5PG�)��5�l��wX(�ںyY���]5���JMhӻ*�tj5�f�ܬ[)��z�tXԠj5n��kC�`va�C�]�T��}��h�g)@% (FfAgm��؏6���yCe5q�lc�J���ׂ�#sYb�;-�c
4,�(�1���$V(�z��ծ��+ ��*m���X/7��]撀x��b�{���wd�3�l]GAm[5
2�.^���b�x��e���Q碖Yk
ͧov�
XԨ�Zy��b�=�����{yb�ٙ4j�|1��
�;'E[�"���H>�	u��"����
T %��(�7CZ���&�R�PZ������S5�T��Z�(0L�R���J���%-K�=���.�b:�L�>N�V�����	U��,�me���q�D�i$��m3�Vkb�۹XHW �����ƩٺBe�%եV�eV۠��Yv��LH-:����7R�h]��#-%eGn�T�m[�
� ��J���q�@��uA�P�	����f^e���l(�ޜ�ET"�?���a���q���$�
�U���2�����R ���c�1�;5��M��iR�E�D6��0�L������P"���sk�tt��h��
�e&&��`E�nc�Zy@��&����F�`�(+ծd�����d�k�h&1���X�����,�i*w)�n^�f��u�;B$lG���2��Vv��ýJ��H�M[׉���@^�iM��nYR�W�o$|�PÚn��x%�OLt[ϣ5�A��Ô��J�){��7�Oh��*�WR�)R�~��t����u̃��{�޳��W��g�jO�k��.ƙJ��	�1���h�(�Y�Z�2���L�MhOQh��^�ʂ(��r̺���
w�v��K_h,�����Z��I��m^Z�Y�n�Ԥ(�,Srֆ�ۤY"�Wȅ:�� ��(@n^T;�.�1]��O�6#�����ٲ^���JkKz�u��_Z�X��\9��Ϸv���O�ǻV��d�1��dPc_�۠�gz�u����Hm!�D���rf@JiӚ�`�Z�}f��ð1j+u�h�6�*SQ���%�y���6���A�@��n�X&AY�Tw� *?�ъK2�cV{c9���v�Yj�8j��
�k7-�Q�0�x�,)�D�Z���y{�	�.�ރG�*��jg\����U���f2���2����%��ػ��Re��
|rlm,WL����n�135	�YB���5�'/^G�yD��1�*M͕���Hn���F�1�5���"����WV[�е��oS��yL�i\[l�*@�ou1�V�ǧt�[ڠ���'.�ͦe�uՁ2��h [�V�1�F���c&UȲ�JBr��=0�m������i�/V+�*�o]*Ouwc�`W�ea�hXZ�J-Q�{o3 Hn�r�G`4laG7M�4S�ZXi�ę���$�p�''��餲�+NaUƻ����°
��`�j� "k��1���j��&Vm��+V����Ė�inQƎl׺	�,jo.�ɫsa&x��@�l�	E1�Mыn*B��N��eZ2��k��+EhI�ł����V�V�k/J�X�ߍ��͔I��b2�ٳr��wQgNm�
�"�W
W6r�F�ß
ܼ�J�+a�Si)&Sg��N`y"Y��-�����KE��ih'���cE��4j��M�3`V��C*�(.���j�B\0,-����r�d�w-w��V37N�o+wBN�z�����Rx�nb��c�W//nӔ�O��`�<��cT�h�+n�a�@Ϋ�g�f�m�s��3	:5�ڹ4�nV���f�(�m�j���ӝ&K�[n�kQ��J�nVd4�h`elT�`ʲ��n]��n���� `�2��]�VӶj�`f�MaUK0���i`��%ݛ(ǎ�ٻ5��%4��L���u�+����n�4�5Kb]��a,�(�Ɲ����%e���	d��42��a���\��sE
7[�CP^X�@$m跕���Iu���|����}E��WOC4ղ�\�AYl*ݺm� ����Ih2鵧����MV��fҧ�\��6�h��ob#w�e��9��4Yx��UފSE�n���I
��J/�I��L��ȝ\r��@H˙-��M=��q�0E�8��x��!o�ú�̹�xx5aM��܋-�@l/R�3+,�q]�ue��Z�]�A�6"����KH�6�̀c;�t��&H�U�Ň���M��y#�����0F�7��Yd��RZE�V{���X�b��5��Po��Q���e2ي]B�T�7f�J�AIZr�j�����)�:�1��7�X%V�oM��@���jϱϮ�<]�{�ޛ���*ʳhY�R! ��e������l^1}��;iq+�1v0��Jʫ���2���V���e<hP�lU�����h�5�d����
��<�yu2kñ3�R��õ���e�un7���d���G7��FՆCP-�ξO�:�:J5�kh���|F0v�x�Y�m��+K�6qKB�of��nځ*�2�w6*��P[V%����K׭QLÐ�w;[�C���K��*V�'m;TQKvOm��wn��p�cF�8-�+^n�ù&�+)m�֒ͦ"!N�̲��7	ZJT�w�H��U]��8+�ek�A�䳳U��cm�d�
�[L)�` b�x.�ض�B�=l-�TG�i�k�-w��;,4��:�A�6k!��S��l�V�6��y*݁S2"��2�1fY���o4k��O��,V�OQ3�ucB�6V��J������͘v\2
�v���8E[�\;n
��n/�����uMd`�{u*�0Ӱ�7SR }Zx�ɹ��;	WfU�F�!fXkx{00vۦlB�LtVbg^SkbV��r[��9wy�R���G)��?r���1��b�ƎJJ�W��y�fV)���\r]9�7��ދ�9{�S�t�CdEڎW��!�8iCK�l�z�;;�]��lҙvTݕr*Q˹��5X��/vÛ�e%vh�UbԷx27Q��rզ���6��%Xx�5���x3^�Z���º0��t-�a^cۛX6��0���Yʺ�^;Ŧ���vJ��|�mY[o�{J�vRYݤ�VNZ����Q&�uaLsb�]�*�m,���l;��t,�9��hiS�onj�9���4F�2!�f
�6��٥*Lfm��&�U�3n��d9�֘p�e%��*�w�%8�T�YMM��G&�R��6t,��a�3n�%!+$���uӮG����"�U����Wf�M�ŧKM��e �+u^������h�Zw��̠Lf *mbZwb��
��ɔ�09������h�!Dˬ��s1��R�)%�,��E��%�!Mu���E��.�KY6��W
�q\A�^kY-��S�#P2cŒ��*�(���Ǜ����T�c��4��%�(��q^=�-��x�p�_QW���&="���2�B���oY�v�9�e`��U���Q��*��Ւ·JP���Q�4�6#�Lg]�T�oV��^���,�̀�XAkt�tƎ*��y�x��ů:���I#{V�O�X��^�u
m޵�����u5dS���ݠ�푚�Wiv�_-����1�ZW(s�k�#h�m�]�z�������E��S�L5��WK�a�f[Q=�@�+�,���{�[`�Y��1'o6����R�{1ݪMn���(�1T1Q"��ܽ`�f�v�Q!+�V6�X�bv�>��C��_�R.��4��hT���f]!.h�;	b��X�Y����ZsQf�5u�o��4oV�C��;9Y�z
֞,�*����+j�������
۫���G7(��a/�%]H0����J�C�(�#V�����6�̧dj���e��iO`���@<!U�Z0�Q0 (]
���TB��x�Չ$���
9�GhÊ���QM-�M����6�-�WX��]�l�O��ʰ��v$R(��P��1�nY6�,b�:ۻ_X$lQT95kN��S���VS床���A����m�t-�e�lt��60CK.�6��2�FdkB��4k@4�ʿ�h9iѰE�e!�w/
E��X�Lmm�m�5Ğ�-|�p|p��|S���ؑ,�ZU���XR�����P�;���ON Ϭ�t3`qMܣyA�	6��*[t��[QY�=�h͹�f��[0��b�X�y	Lh7���W3HgZ����_��¥l�$֔rţ`�j��Z��62̦N^�E��y�~f�"���ʷ+rj��DQW�Ѽ�R��o`���
�`�R5y��Z.���.��or�n��f��C��@j����UƳR��pY��b�ֲ��WN�Rk^+�;g���U�Lw���3p^�4ZH��q*yZ��pLb���At��oÅ텛d��̀h={�
��8'M�j��kµ�����䭇F��W:j�奧q-��k	Ư'�&���Շ2㱖>�xFm����������9#>��YRu�65,'��W�w#Y;���j��ܝJK!��096ĵ�,å$��2?�#	�r��v}���f�Э֥��ۘ�`��;$n�ݭ=Y�+��"���Jwf�|
�n�J����[�]�EC��n�j�ѓ/��[�/��bb8������%c(��>*��7e���滧��ung]ݦM��l�V{H#3D�f��ͪ�"1��x_vPMU�̡�3(�"
E��] �R�@���	�w���y+s� ���t�YE�&���=͌ԧ�M���]�k$nr���'G9C��գ&kF���*'Σ�N�v���t��x��1\MoEbY�tG]�B^��d��o39�r�eI�ԝzF�{���)�ښ��!�]7ó1��M.��p��R,�V1Z�����b
H�>&��[�c���f'��Z=ٸ�X,�����z�Ri\/���!c�:�e�N�A{B� �zUo*r�β��y�^�]�h^��ZXs�>���肎�9[�<�Nz�G}���"�6�[��^�T8��z�S�*��+&�J�����j���;����B�1��Yx�q�,s���*o:�Wa�����֖DZ��4�����@ouպ�:�P���Ű7|;���z��%<(����XC�+X@Zz����ܐ9�J�4\�7v�:ᔻt�&s=7IF��g��:�U�Li$�_]h:�_>�4���&����S�A[J��ֺXz�e����R�u�����7U�|�S���.���sNngE�YX�;�S�5P��N�\�������N����ʕ�+�s��}t��WIu^�����njW�z�H��Ƹ�>�E�lR�"]�5;Jpͳ��8n�e�3F�v�,Θ.���!dM� �F����\��I�v�Y7��[���3hS���fbI���rCO�[�@����=�)����5�;��z���;�gu2Ve8��	�u�F�(�4q�w�4(H�MT�U�-��x�^�p�A��˷��y�3	w��`��
�����]�dd8�
�N��Հ��{-�����f��L�ʗP�Y�=]��܁�`+�܆�����]2�J��4-R'��{�e4P�V�����wI��{�����ʻ�I������ڜLu��x�4kܗ"���@����-�7y9����3����Bҷ�(+�c4��t�f\�p-�2,�3�9A �K�v�5�.��Ck�[m-Uύb���q��}�)^�S���]rY{N�$
��/�h��}��:���W�J��k�V�Cv]�@Z��9)���J.�-Ѳ�xT$�|턷k!ݤˬ T�Ȍ2�4]��x�X��ʚe7϶V�V��d��}�&�m�J
q��he��vDS(濙���zX���u�Ћg/[��"mc`V��t�ސ��Nr�9��6�d��1�k�+��R�ܱ 6ɕ�p
e� `I�fV>"��0uB��h���������5�G�E��S��z�Ml'��~c�`x���G�Y����N�2�����rD_���'bs��ճ�X�N�x�h9Vx٘��+F�@����a
Y����ف�"���KQ���o��ǘ���:��!O&�0���I���Gk3MG!�V��U�n�8E;Q�t���!�)�}��Ш�,A-8
�h�8lFi���}���>qv�f�.�W�of2U��yn��#t�j8��v�˂��|�*�r��&�b7���i�uv;m�����Q���=�jZ뢬�*�fT)�{�{S>�}n{,�:�7������h�ɼn��Gq�be�uݵǓ_*@�����[w���wd,	,��v��u����Y��|פ��SfQ�؟m�������فq�ci�Ю6�>3��R���1�M��O��&.� �K�)�[��X�<<�e.U�|^c��d���A�Ц��ET�n�Ӯ�|(�3����� :X�k�F;�n���FU�|N�͊U��!R�	� �k�j�ǆ�t/c�!�������]הK=��A�KA.���\j��x���%Yz�,�J�5�%�����0;�o�2�n'*du�lfm+�r��w%�,�1qV��Y!7�/3��HŻ��W�ך�e�Z� "��K���J��c r̷����Y�#5�ǹw�&CVjn&GM�%�V���|�<��-�w,e�؜�T�k�\9�+�ŚuF�20Mj�md�zQv�Jۥn�;�q-Jimm���]w��ծIQ܏R8�acF#��E�Nd�PADQJY���7ҩq&m;�y��ӳrW[������3��g,q�wU+��im�a.5����#3��o�M^Y����A���Z"�Z�7�����O �]n��B��vb�/��6-È䦖�5l�Txt{]W�iy�����y��X���[Y�8��2�]N�7/�+-]q��WtC66��xD��Z�d6^�3n4%â�r9h���<��x��;�t�]��Ro��f��z�b��Z�hfY�DI�T`^v�J	]$8�5ǁ_��,�*r��0�۸��:Bp�Hߜ���Hm̱�>b�.\�tP-Չb�摶��^�$�.����RUI[0;ɼ�Ծ�ظ:�oa�`�R���H!/'��j�R�Tv��ͧG�C�Z�C�]�s(NJl]�6�!�2"���P���H�]\�Da���hՒMU�;���#����T��ҭ<��|v��u����*$�U�f\��fYu�^e�f��,���Y���г	�`\���ʀ��ȶWW$���˒��r[4��h��0��оP��x��˕��K�e��{E�\�	�~��f��������r��ۈ��m�6OkF�	i��+h�Bko$��n�i�OmJeZ�&l��cٻJ��{fY��m����4XD��e���f4�7ǂ���F��}�� z���5zE�t����o����(��7�u�s����D�Ә��v7��e�ϲ�H�%�GP�ӛ`���"�m8�k[���P�V:�j�[�W��m��O`�|�udL�s�7��C�Xa���ݻc6�&� 1���U�2{Z팉����I��Z捊z�ܹ`�gE���M��	.�*�Ų�*ʝظS��ɏV�Q�-�+_jz5ۄ��駕6�r�!p�(ve�����>�j�\�ؐ��Z��9˦к�4��"�`;y`�Nn��oy-�u��ˋ��!�.Jξ�5N�)���Q����Vu,}E\(�$E�2�����+���t���ۏ�֮�����6w�s`����$��dX��}S+��{2��,�%^�CBm�������
d���Eq�o,{{Q�a5�w5�L��;�H���3y}�:�A�H�R���w�0er������WD���t���L��lrXʸ2Z]Զ�����/j����b�;En����6���|��WR	3n����z�A�TLIFS��뻑n���J���=��O��}�{�1Cn�l�[�Q� 6J:Z.��W��pWi���p\�+�,��;��a;ݨ���YX�k�6sa����r��v�K��� 2�@%[�켙�,�N�N��mte>Y���:�
��s8�h�w�M��~�>�U��.sܢ-h
�����y��X�O��s"���h��v0q��B�i����"�;Řʥo7n�^抋a����Nf�f��QÛB���U��qV\�b���&�	}Y������wd��9�T�V:q�ZiM��p0�>�h�ˡ�6J�2b�z��Jy�m�WZ�Vu_#zi��8󺘏cY��Xr�J]�N.��Vخ:Ku���X6��쿻��๜��_-����WH�l[x�oA���Ew3��(fΛ!Eҧ��w�2�Ǝ9%^M%�Ƭ���.8����ǂt��Ș���V�D��e]�����+{uݲv;*�Zئ8n�1w��6�(Zh�u�z�����Ol�c�,ﰧ����x���s�U���MC�Bq���8�L�}/�j�snb���jã7�4$�\��?Z$��0�E���o7���x��-o�N.�VDIs,��衹n�wS-m��e[�h�u����֔�6k�t�-�Y ������Q�;t_\�v5����9���g˹d��>]�^<�ƝM�ŤK��B�Q���H-�ySkX�7s&�қM1�ef��ǦF�P���Ua��Ӳ�M7�F����n��޻�����aSsZ�iꖲM������g� <�V/Z�u -�-�N���^�e��5V�J©�r��a4��:�]�8h;�X\���:��vs�7�v�U��A�[���b���t��S��4�kh��__IP�rN,���_S� �ON0�UuJBk2�m��SxT���[>ݛh�m������[4�ݦ���_;�FC/����8]�J.�e��}/�&�+�\�)_�z��j��@+Î���"oPEN�n�s� ��G�n��r%hq��ok��(N&C˔�T�u��
�M^	.�c/�6\����1ڹu�Ǳ��s�LT_C�Dw��$JYWj�=�ݍgl��:��Ϯ�U�k];����ɒ]�<Ju��Z�
c���lJl������(J�ݵG/�o��V�4�봭��� 0���ɽ�U�g�eA(=���h��e>̪�����Ǻ��z�ڸq��5f�� ߍ͐��t���@^�;U���'�-��0��T���*��T��m���{=�$4�v�I�r�֧�N����:j��k��Nw�5�퉓&c�lp�{ʓ�-���ba��q*,�\J2�|�ïu6�}��ٴ/o	F�e4����-�Lbq�̺.\�nó��_]9�E���z+�͉�q>��w	Oo���ŵ�5�q]����{��nr
����4s��|�m���7B}Zݏ��z�ͣ��E��Pi�}k�9S�!�4#ن�K�u}Љ����b��;���`�J �ҭ�)�W*�/��#6�i��k5��)u�PjėwS e���5:4^� gJ=w��GZ:�"{3iue ���g'}E�^�+se�Ҁ�0�!�R�ǲ*���x��)��4�2�b�Z����_S/�PvS�X/K\)T���8ٴy��W�nYҐ�'*�j�x˗�K�0�i�E���۸�#�:0�7�`���w}rCm�jcn�����3�b�R4r���k.�77SO;NrA��޵��3��͜�'M�U�	3(wi�io-�w���d����mr�h���d�/4p�\��t�$��D�C�n�pfT�ᾛm��X�Լ%e፝��3�n�YV�X=*	[�e�-��s&
٦BT�W�D��
͏\�Vܽ��n�ڳԳ���N�٫����f��㡎TX2��؎9�+��L�(�%�e�6\�M�&M=���Z�tRqD�doW^&�U��7D~�I��y	<�;�x���b��j�+c�(��LݎJ�iw2��n�߂�
�TG\��C�(�ꑺ�+�>[.+W�@�)���St�>���+%v�Z6�;C��gX�}����{d��5��p���QR��Oqn*��:f2�J܇����;ϸ_j��%�V����IZ޴�M�nڰ;�5�qc��n�L�k��L�\���n�8�v�xf�!�7��b2�#����}x�'y(�,��P���!;8wp�F���@��_$�����t����wN��T�k��/��u���4���C'�����Jw�N���	-��oOOPٛ_�������j�ɟ����Đ �'����p�! O�ϰ$�&��� H���_���]u��=k�󼈣p~����-�"Qu�B�m�5}�n�ͱ׭\�ar_��cfq�9e�uI�Y��&V�'�����&�O#9�X?_Vޗr�P�m�*݋�t������T��7:��X6��V���I9{���5[�5$Cw��P�ā��fU�I��R׉��e�rf^|D�q��U�K7�4�Ga��9m%XN.�ܩg��Z�ڈ�SY�ݸn��Fc����i}�0"�������w�:X��Cs!n��Z> �^� � �����Z�����{��EsJ�'+��{�`�S �}����^�zS�V�����>�sEpf@�V�kv]�M!�������k�����;��]�a��¡!��q�@��L�k��2f�m�'�q��nK�`wn�Q�Q�#�tņ+e�w���-H�wx��SR�z����
���)����싪��]�V+�M��c�*�u��R�KJ��p۩�x�P蛡v7�g�m��u���X(	��q�F�<�� �#�r�@Us�S;�l�.�r��`��)�Ů�p��
����f\z�#�+�*��e<BTh:�w]>�r[�ŉ�w��Mcuz��6�;���l*�ǅu�:���8�ă���U��o.�q ��/���p.���ya\
�vd����QkI���W�p�,r�&@�g:�:���J�>&����;.)��Vҙ.���(��v(6-�
2ѥ����7���x�f�Y-��v�uԧ��>��LC�;�H�u���ᤙ�A[Ӯ��M!9�u��E�fỴIѨH8��W7��<U�$�;xc���WR��3q��� &8���#�_1|C�6�Vg#�R�Ү?;�Q�l6����P޽YV6[���|��b�����m��evu;��f�))�VK���,��&3[�o-Z����Z��oVuԴ�e���TI��)d�/��Z�7���&��������3���g��X{G%o���J����JW���7���
�"�jeu�fV���Z����⥺�؆r����o�)�"X���)e��je	��{@w*�ܻ�F �tx��Ӱou��1B�n�X�����J�jDк�IB;�&����"���ܢ��p-��!�An�dNm��̦�t+�p��pհ���R=}��v{�>n#��չ��|�ѷ֙F6��o	,i�^+��2�*�q�v^�x�V�fF����Ex�y��)ץ,�S�p��rb&������A�k��/��EM�6�,����#�k�X֢)f������*����}*��$b{�����7�Q-�<]��ŭ����
�Z��8*��ndr�G[c.�6���x #�ܘ���z����݆E]h=�� m���f�ܒu�R9�W;�ߓ����F�I@U�:d����6Me�B[��.����X�)P��|���$A�"%$n��1u�qc��^U� u��6'q�]�9��-a&uօ/�ⓣU*o��s���b �Y�ݝU	5V�㙵����ҏv�5�4��X�F���H2f��v8S�ENT��C0-:ţ���Ku�4H �;���31s��qhHU�����鎍�U��Qj�X^��ुER���j��Z�7�V֝��{kz�E�\U$�Mys�Ζ�L���g5�܎�
޴Q">,˥y�hĨ��K��~��}�5m]�붝+�V\�0�en�Z9��r�'g�X��R�:�B=;K����Bo#X��s8mu"N��;(������ǳ��eC�R�ݪ$��\�7��_uE��('�U�s7Z���)�"q}ʁƋ�l�9pAt�@�C;n�/6�2�Z���wz]m˽�zC����Ktqv�Z��H�9�]�-�|,S�ׁ���WZ�hYӔ�N�s����$fT�h���棣N�'lg���9B�>�6vS�6Q����T?:]�t�0_KΜ��x���Fj͠��0�`x��!�@]l+�m�4��n	���aN�7�9��'�8��6�;(�U�h��LBp7b[��Z�gM��8$�
���r��3�']�f�Z������ɺ黽	�p�3v��|��N��k�V�X��E�2�gv���q�-Ѡ�:�*�GN����Z3-���P����#M%�SP��\�P��e��ur�,�=���R���ҙ݋E�v�I��p�P�3�0��V5N�˝�*Z^s��( ��wu�	��F�rO�����  �N���wB�%�U�R᳦�Wΐ#vr��;y�n`��'��W�e�Z�Y�O7,�5�Yc�����hb�$�H�VZI�b�s��Y�b��Jx��x8Ԩ9N�ʶ^����&���d�M���2mp�L�/3��4[ٵA�빤�g4^���9�SrN���O��lq�A���p$�h	�Z�WW�&�B��S�>MZ�.�r�u���YN��ٝ�螹�J�Y��<8M��$u�.�ij��u�R��1'��&�j�Z��J]ŷ�5Ʃ6��e��
Ph�R�Q����V�[�>���C�3p�=��,&�����"AH�ݝ;�hu��岻4]&���|*�e����2��#s������A�Y5���Mo�S��e�EX}��r�N��e�-lWǦ�%Òki@�Q�����@)�8�o9.؂�3��c=]�ZuqѬb���&��
��p1�v�z�)�4��ͬsbA��5p1�Z��.:Fc;vst���h�7{Dv��*[�w6L���\ON}H����u���|��fe�[pe�5�bM(����Dr��q4kqSN��^���,j�e�p��ɥ�MB/>4�5^�=��1u*��=�k��l�$n�:b�OE����e�-Gv��h<N�5�+k5_��`H�
���	��f���m�:k!�Xԫ|5M�挽a�m���^�Z�닖Z�U����n�g���WB-Z�}q�������v��-�gq�]OCa�����LԒ,�Ǖ��{�)�U�uA��} ]Zpn�(�R뒘�&�U�v%R�!�#�:�]cC �!h�QbZmn�W.�Qm
��Sln���l[�x�2���Qyf�n����Yd�9lt��,&��Nb�-*坺��[&���n���ik���^u��Fh�,
ur��֜�5fp��T���V�&�f��f��S�WFV���ոb,���׏lb/�u����:�&=x�)���fr���pd�՘��T��ُ��;���V�UGC�Ӭǆ:b	S/��%�Vm`)a��ב�َC�K&��Yb_M��ֳ#N�m��V���X\����ݺ5�m-T�)�������y�;�H:{Z'p5i
��J7̮&Ѯ�AZ�w@	L;v�s9���&�4���,��;3o�R�Q ;ֽ�eE�HD3�!�����ᩂ�B�<wN	;aA�IثA5�ۑ�{��ۗ���kMOH��&r��5�_LB�����Ye�k�A��W>����+S��Yc3��TAly���U���S�ɑ���;�aƷ�@�a�}n���nWe[�ս#����ç�W�A��I�b7�(��)oٻ�t���t�q̂D�A%MCF�Eudeۥ�7ٮ����k��!�)ك��ʁK��UӰk,e�&(&b���L�T��H:Mɱ1���˺����t>�-vmc��.��׸#�w^�h0^3CC�7a1�od�<���2I%g4 �\n�TۢA�4L2��b���d��yrSܐY���ǛN����G$��#���Zel�>�5�P�呋�)<�H�W��8��>�Ұ��WJ2�L�;��Ѯ���a�Ώ�-�1cV2�8�A]D���M{ש�xVb{�w����{dě0�mt�.��Q���g�E�����r�2�;���o���6�@�x~�w�U�I<{�,���Y2T<�ѧ��pڷSc}�5j�i�,ӛw��=`�C&u�fժe3�݀6�B+�t/-�7�yf�Jɪd��)�������충mws�v�NNn�iɍk��ˈwG��&�M�B���fM�*����>Ng�-.w)�e��{��
ݡC���Pf\�h���lG��h�#Q���a���7��]m��T�W�Q�M����-e�G¶e�`��u�7G~�A9�7�������QČ�wt%uw��v��2^Y�Tx[#V;mӻ[���DMD��!�]�[��6��I������ᑚZn��.;�X�L��� �&�Z��do#Wr���ye�.
���=��:Ɲ�%)uPNζ��v������=������p�46��)�������T�6E9�f��I��4�W��]��T&��z��YηV�+��b�$dS��S�,�hcw�a�ܩ��"胓1��'�6�_]����SzDqv�
���,��Ŏ¯Iuh��J�1��v�ꀔ�r̷��6���}n�^R�LH���\�1�Y��B*Ձ�亜-����v�̘.�I���M�C�ʇO@+�u*N�9���mK���w&��@#�ۑ!�*9�����I(T�t��U�����bě5�n}����'U����2MEX;M�4�FHw��jN�b�Rw���9ۚޖ^�'����Z�cg5C�o]�7M��um�v� ��N����̨������e��=��lL3S8M�U��,q��I�,m��y{ç3;W�3v6�|)�	�sy��G�t���uyl훃Z0��\��-,be�{on�p�7G&�V���؞m4*�:�c%b�t�8�^2{J��!ٗwݭ���Ra�6�M�ZV�H���`��E��ֈ��N�miv�<����v�;ЈҪ�0�6湵�ǋ�n����TBYZ��ڝW|�o%�΀�mq�)ǎ=��e�:ߵ�O	e���Z ��lO�+)�X�Sj6][��`��mk�(m�������G�۝ϛ�avh<E]e �YA�:�늋�x�4��&���*Z�wQ��	�����c�jg�A�on�	�SSëO^T�l#���Tm��4�U�ott��<�'ƛ�ݼN���!��Ƴ�}��ݬU�ƺ,��Qtm��#D|�	�����gүW\�s��f\�
�V�N�[��b�3k{`�O�,r��,Y&[��v�$�L��ظ寇�6RgVY�4����5�  K*6tcYna�31���(�쫊L�Ev���B����iY[��e=��[0���TH�K����"*k�����|�^���p�����3[�)�19R���R.�c�%=�s��$�s�v*h�sR���6٧[ht�����R���=	a\g��i�.��y��f�s�����՝҈��hںY�wṻR��k�F�L��B��k�_��.9�>F��h��JJ{H�b默RBh�*v>�lZj-���f+��k��Za�m#Z{��ݱV(I5�������x�_A�b��\�s5���m; �͙�/
��W^O��ݬG&�
8��>����_Gԝ`r�˒��W�q�	�%pY����CK�˹�c�z���0 �'�R�V7r�,K�+����f�E\f@�թ)�
�ذ-��:^�d�#͊U��1b���$�xe���k�&�>�2V[#r3��E�G�;��x(�;�5I���&��Ջ��cS�,7ҩ�m�m���7�Z�H�U��'Xb��\q�+5ф��&Ŕ��S��;�����~  $��+��d�zLO�����3�����q9$���ОXϚ�є������[2�
Rq�����|'X��Y��.އK�*v������v��qor&�JU�4���=��N�ۆ�v��WD��Y���
޵W�έ�V���mZ ��p]�,����'�0�e�Q�yM�!]�v<�u]X�2���>#B��b�Ӕ-հ��	W�:�>X7���/���6o)J�v�f8��3�S6m^`<�n%Vq_`6�w���a˔W�c9�`%�&����T�(���Ⱦ�=�����Hi:'�"�*�t���.  ���Qw,7M"�U��o�ٙ����K���8.n�j�K�"�u�]ϻgX�P�jH�m9:͛l��V�+;+4�Գr�5�]n����Ih�G��B�^8�>B$0HO�����9��rc�����+r���Z/��/�0�e����ʱ��S������Myչm]h�(�Ye�iެ����������w6WV�7�^ۗ���Kʅ˛1�9�E7/C��б�;0�B�ͽ'�����q+ǰ�sP3H�rh6����1���w���1��pX��X� ,D�z��V�aR�i�5��b�X��t8���+�*(�X�̥-��6�)�28�k`����"����hTFZuiZ�լ�jb���b��b��2�E]%:pA*T�VM-�������+Eq������c�S-5IEkUE&$P��\n!H���DX�*\ːmjU�EQAD�Y���PU�\�QG��KU����5UV:J�Db2��S�M�6���
#[�Q�R�+R�(���U��8e0QKJŴ�V�n`�("V�����Dm�0Q�-Dc]Z�+�TE�+TR1����"�EUƦ�Q5j��s*��b�ZƗ,�UX��%n5C-Db�s(�R\B��f�i���5F��QT��4�B�LV
�V[�U]���� �%�϶�W�첇V $���f;�=�M��3�����ӾzAܫ���]!,و�ݽN�}�̿�P�������'A���H�����JR�s��)��P�v��,��ӮJ���1��o;��x�����s2ڗ�_2�l�<�4�c������^x�d�S>����S��v�2g6�v�����(�S���P^��96�?{�/&E�x[+|L:SθM�[j�h�;�P7��A�X{��c֟�,�C5����%G��j���GQ�q��}SV�����l��F4�N-�ۅ��+��2$�0����y�֠�ڗ�D���õ]����R�s�9����ՙ��V�s�s����a��\UV�����q��J��vtR����{7����k̊~�dE��ʯV���v�ۊX������r>�غ5�U��� i�����a�9H%�M���Z�6��d�xm"4��9��Tog*G)��{0���N&��nge�,��Bv�����bbfW���of�$�3��To�"�Qt��Φ[��U�����`���N�T��N�:r$]9�vr� s����p�*f��"�,��U�\!_o?n�+�p��H� �F�z;B]�O��v��io�x�Y}����Gb:�ɘ��l)E��L_�>�c�_S��Q�Iw&Sf+3�4Ncv3g�;]dI���Vw����<j��sSO�ρ�R�0vӼ�W������u�aa��jn-8�-S��|�Fi-<��i;���1O��\��ñp�ꪧ`I�i�m��.�ᦹ�<��յ�j!f��ɘa���"�1�;��+V��\��J��΂��
ι�"���ӊ��_kYsS����z&��D\�����[j`7L�e�n����7���)�]y�F�ٯ�["R�	�����e,W�D���r~�wQ�������ä�JJ+h�IF��Ɣ(����0Q]�a�x�<R�-HU�m%9��u�)����׸Nά��.IP���G8b6#���=/*�wo�o�i�O�댨�C�����V�C�t[:�ʿ,��7yoϪ?k(g�B��-q��z�ɛ�H�ڊ���h�iW������z|{0F�{�i,��B�Է�~��mDE:W��g-[�{�ć;uLtWm�o2��q;�}el'>��nij9�ܵo�G��.H�U�&?,�%IXu�1��b>���	Q]�iM*�l���S<7H�]��U$3}0:�����- mY��	BB�ơw���م��]�*�V�i�0�uQ{ts��ʚt���)EI�c���J���&k'���y�}�\ �ZUq���g��[����9.�=Ա�E����^�i��9�[g���{ҹV�T8(Nv4WJ�)Z�WI�fT�e�0� �E2��ͭ#;��Qa��lI��ᶽ���Z����9��ں���U�����5{�oJ�'5����c�j�ֹ�[!�à�n�29���2ILM륮,�WvO�!0����{��F^�/��e�^0s�����E���	��ͨ¦��z)�x��ON'������rj��7����=,o8�Nnuo���M[���H����o��f��jV)�%ePS׼���I�_�W�H�Ce��o g6&��)�R�`�F�tt��8�y����U��p�kO�l�2u\b��q�����2��Q�u����V+��^=y�I��{��&�J�M׽���k�؟!�SG$ �^]�]��a�L����{�.�W'0��LG1��	���yOXǭؠ|�igjӽ�+[���z�����W�@�}#�qf�3W:]��%�9W:��w|��G�ay*�p X�����Gd\��Z�����p�D+1�*p
 .̚4� ���X±_�v�k�Y^��v��{$�&�6uȲ�������V�kqR�Jlr�2P���}�H��bc�b�㷣���АZpv�)�"}�l-��N�u�p�-9Ŋۖ��Ž��R�7A8��+�~G�c�-������e����;2�OD�D#�*��.)�W<7�u��T�ʫ3��M:�����:��WX�Bpc%�������zj:�϶*�־�n��>b�2m�JNJ�r�כ����m�-w�ڂ�9�3�z�=-ɼE�T,�ۑ����߈��x�y���-ၧ�����@��^�G���V�9�,�^3����0�{�Z�z�,�T��{���w������s�5��Hde5��/km�*���U�Tcy���h�|!vAj$�Z�vS�|��5�X��]V�y�෭C�q�&�ƍ����EMJ�TSe*cydPkHc�A�Q��ܲ�&s%adR��$޾�]�ub����'kP�s/+o���cz��9S:�BL��a��]>����+�*Jk��uXU�E)c�c�Mf�qq��ez��o,�_9�tc���~q�ޅ}*U�8�^�֬�a�5#F̾��w��f������f�v�Oy%p��������r�U��[��������w}!�+|5�ru-�
+'o��kf�Eg�[�����b�~3�'ws:���'����5�{;����ʈ�CD���\N�����ܫJ�_I�v��0՟����ڙ�:�"��J��*��6�Z�\ʺ+�K������F%��s��_y�_2�.���1
4�wv��|����M��}O�Uf����Zc�1�C��Fb_nv=t�l��ٺz/j��(�u��51�6m�q�[~��)j�F�����/z�'�(�����	�S�7�L��]!d8j�{ǹ��7��t|/8q�/��JI[�[|+��,.��m�m�u�fux�,�Yo�~�H����4����vZ3\�:�}e%}(�u�d�S�AvV�j��G�۶alc1�9#/'{���=�.C<��w�Z�Uǣ�l�y�.�k͋a�I����T.y{yW���B����*Ċq�t��F��z�*��u�O�;����ok�u��w1��J*k�N��kSv��<�r�߻��R��+�{ޕ�#y���\���*�AvÅ�☘�T[먾يx���cl:&ruȉ����|�Kc V���Cb`-��{��}ws�ͻ���ҕn���Ns5�x�=ɘ^�YiW��y���#����v"{��~eB��hM7��H�Qt��߭[��ʵ&���i�N�Lc���[�j��m�5��9n���)u�c�8���:v�:˯W�nq�*W	QܳT��H�W��*�����gEue���f�D��d�bZa���`]v	�R�J�lw�T�J�I�3���1��$�\Vkțw).r��ܼ	�'E@�i	o)>a��V�؁�ãwl��a�@��\���z�p�pgb�H6:;�sTq͏��p�:�pwWd�秡�|xs��o��K{�"�,�Y^��4���B#M����׽O��ٳ;�d'tyټ�cfꨃj`��Й|�+�{��M�|��i�/�鍋�Y8�Mu��+3�[S�\W�x��)�[���}Xr�k�O&=�t�k{�}6ݛ�	��x��� ����I}��3���'���W�T�<MNKg�]ݧ��� �]�S����8�CZ����UF��cx�j�(��t��$�Μ��r��e8����Ts����m�pf:"�v�(q{��7a��"�`�F�tt��8�k��0�{�32}3ܧ�^�wb��p�&�����B���q��+�n��n�n�C���q&��%�˧BGچ�R�iI�t#Cr������+�ڐ�J�(�h!�����D�h0"�� dӼg�:�J����*e�{�w�tg��sz=����O�E)�܎�;��3��$�3Z�=]�;�c��S��mmC�a_T�z`�;Y2�'��H°k/�����;5TJOG�^�粡�\�d�t���a�y�s?A΍^�QX�'zks��ǩ
�]�6�o7�lΨ�n̤8�:�N�1:.}|��c`��)�[2��6i�T��\��/�,)��4D�Pـ�GԎ�v�1S2T�7��>G���K���BY1	�;G�c�-��%զ��K�����ŉ����8QJ�Ah�������}�#�uF��1�8y����<2�T�+�PrZ���q�Zy��P~_x�%c�O]�ʇ|�R�_���o1*��;J%T�Wr��V���w���v�1k���U�Y���pW5�!T�f+��	m���o�WT�W\�Jוb����v�n�~S���+��k'�L8����V��{�;�C��GGbg� 1�-�@s��,�J��vt�^CqY�(%����x�戓�+G޲�.AxV֧�k�^V^�y�;,׆.����d���Gq5b�A�y�y['��jC�w��W������s�0u���˽�j�Ǚ�9G{�\�oV'o��so���.X\|��嫬�����,�jڗ�?ty�x�-��6���n���o��!�H�U�W�ᑕ/�A��H}�����]1Je9�����VS5u͉�������"�w�l!������k���UJy�$q�7g��緸�whz�j��J��g��U�c�C��j֝˞���f?u�f�ޒ3=\��V�Bme)��~pp��9_���Ff�*�pov4����B�6Z�:	����-^��ov�^�N�^�9J��K�
m�8�d���Tw-Fe!dn�Ӊ��?g���z>��3����?�V�D�U�l3���1�ChG6g*�'`�T�Fsn}��;�^ű:��=b�*�"x�͒�o\)�|[@��b��%=F�R͙�wJ�.��;Dmrv�ßj)�> �]��Y�n����9���zm�O摖B�aZ�&����r�l�a]�4�Dr-��S�&����I�W�y��&ܡ��Ɯ�[[��	��y�G��]y#b%�Ik݉F|3��Y�{Tk���ɖ�<ُo\5 � �CMr�[2��7��
��hw�x�U���j������W���gtO<��u��
��������L�"�y%I���z�3�*�'�[��U�GP*5�J�w����kIw_%-�Ft�l��z����K��i����P�YZ8� f��W4K�_bX"MiM�ņq�օ�PI��]8��plv��W�&1�
�;nǬӇ��R��Z˼�[�ґ:f��\��mK��3�w��ώ�p����@!f��5�0�����l4���Y��ݨ�h@�Z;kZ�ï3���I��jK9�u9������kmX{�x�chnAɱ�y�]�ԺX'\@uݼ̩qX��fbm���h#4tG�kWf.ݍ�5��o��ii����nG�u��l/������,��bg#��L���T��	�ѵ%k����̊�GW]�:8��O[�6�W+֪�fn�rf�+;�MPP"@`7ݼ��v�e��$�#�U�'���Ȏ֮�ϗa���򠂵�9�5��y�y��zn
;�W05r���%ƨo6i<����81J�u��ihr6+�C@;5�h�ų@v^*��ژ���N��o�,�X��J����K\Ca7�P�Y&r�¦;*f���w*Υ�P���IŻ69fGY��i��B�j�������Ap�-�2�%�tT��@]�Ό�9��QN��E��˗f@м17N�1������ğ[*|���ɲ譵����nq�Ӂ� ���E�zR�,�.������):�>���q����
_\�,$vɇ[�,�ݬ�;&��@+7�1x���5@�%�ވ{^���L\�:;"���U���hBwie�P;�yBL���bq��f :����.�Kb�/ju���6���2,�͕�e��R;BSiM�rT�Us�"':��!ME�g5	@êMq�5��r�]��̴�E�5�1�g��2��&r�����{-����F�adr�b�TkV,�*cr�F�
ƩJ��"�R��\ƙmn���a�����+++hTƠ�m�2��j9B�Ѡ�-&4\�F��Eb�`i1՗��+(ر�6��Tu@���s	��Jq���V*i%�5J�����`��()���U5MX�5b+K
T�����m�IkA[j�0ӫ�P.WJ��EJ7\�1�q+Fe̠��"�[J������EYm���m+J�QMfJ�T�՘�T1̪����X�t��m,ZU1�Kj�V�WZ�-��r5���PY���KKi���mULe�f�(���0EL�ER��*��KTŦf�Z,Z�F
�h�TjɌR��6K10®���1��j[M[���(��*0Tb�F�]e�-�b��%������~3w3����r���1Tt��ͱ3pb�sDp(.#���`%`�=�����V�Q��Qƚ����s?����.>��r���Е.)�9fm���WU��Q78m�8+"�x�j�W4�~]M����s�7�>��{y�9CNc��u�/h}�˃�gʣngԭ��y�uu���ݥY�IC��.��~ov�]񬱨M�Y1�a��]�1��>�	��y���N#rr�1>V�\sݨN�osM>�Rz�nrwU�;�7^�����k��Lo�z����;Ɇ���f��ɐn���&K��ɜ�N��[z�{��wM�Վ�я����ò��ü�~���W���Bz�S{]����t�qgl�u-QںX��cI�=LvҸ5��&,rw��}������K��)����=�R����J�UCaǯ�֫*�ʿ,��w�Ϯ:�to^Y����;{��3����sXι<�E�y���[Lh��!8{lb#fT��w_їQv�n�J�� �E�N�ٹ��4�5��%3O'p�X8՞��7���٧�d��2��T��8S{�����g�ڬ�{��o�
�:�Fxn�8�Kޝ�����}��k�V�.R���խ��Z���}��{N+3ݞ틐@��Y���[��*���v����M�{v����_�����Ԥg��g4��1��b9.Qn,��mL���4�(�ǋd�/=-v�,��Ao>�_��}7�L��Qg�I��*Bѓ��J�:�Nx��9��wHv�*�%c�IGe��}Ɋ|.S�5�W������ژ8���Nv<��F�]Z�U^�aHt5��k'��OP�����m�s.��^�E���WT�LjA]7�3۫3�VU���ky�@��V^Y�w�������ES��3��k}��{^�-�ɡb��\+5n�:r��6�æ9dD�;	�����5�GK	���l.�W�>�x��Vnpث����eQA=���;���䫻�������Wf���a.\$oH�y��J	5g6y��-����Rts������3���*����cT��m��p��\�>MD�L_%E�B�z�3���C�2U���õFW����PN�{�fS��=���0R_j�
�������{���-��5��MӸ���Q����[����^�8���ы�+5TJ{����_L�sx3F_�?BI��-\���oC�Q��ʦTڔ�Au����R�YS1C��n�Oqz8��AZz�PN��>��5u r�̚p�����ݜ��uy��c��:�D�3:.��
�덮�}�\Ӷ�8��첚o�X�:�������S6i�|hc������8)3�	�R��2в7X�b�nn2\���� �5^XlО�EWdBi��K�W��kyo�ux�A��Η�2�V.��ֶ�u<4[�b�~>�C}�f����RgL�W�Xj��spq���J�VGl\�i'qӘ����u��2��N�����o�ޝ.��D��[��Gg>���:ļ�h��ՀUs���^����mLұ>Ό)[Xض�N;�j��6�=~��e1&�;�ճ*���Id;�&z�Cq��g��b���l��U�G����C��W��������艋��YE�.o����V�(��s��W�P���eV��d�
�o��B6(z��1gC���l���\�㷴W^(����^�m��^��z�"��W?=��o����������;3[�d��w����/�k�\�v��ٯ<��St�N����[�n�kVgp]�>�/��Z�T�{��-�2L˽q�ٷ���t������Cv{��=�����=�T�3��s�
��+4y��\�HB�ѭ�/q�S�E�|�#����[k��T�%�	U<���|�*�֎F����z�^��U�����:�_%�1�Ͱ���\��dAS˽�%p�̢�
ҡD.�LH�	�L��\o�Y9͕+���7��C����[Yn����ڵ��]<�o��;p�K���Zq-UDQ>ޥ^�&9l�r����{�k��2�]+u"��u�6��6Z���X�ϩKW�"��zϟ�OM�"T�}��c'փŐ2#�%���5J��لe���ۭ*�P,N1���-�t���d�Tv���̖�U)n-ɺ��)Vʴ���>cf���T���2�PO��������֘��3I�m	1�V�1��;c�6hOk�"z�='��׹���+Gu45�ڍw�(\j�������������&�ؽÎ�xT�7��	sQ<G�Χ�@���S�C��v:�S���gj�;�F��*������U�ʔ6h���˶K�FK;t�&������&�L�(���0��z#5!J�<
�֏�C�k�,M�s�گ�9�L����*\4��մ��p� �+k�5�T�R�Z)ˑ��$Q�v,�&P�QW��2y�rS��7�S��h��������e�پq�.U�>���ַ���O�m!ھ��sW� c>���T�7�Bt���f�%11�
�}u��M2�]�tEO8�}�9Vʞ����^�9�t1��fك�$s�pܣ
/�Z��U]��>��y��7�W���/_Q����B�`����_�$-	�>W<���~�M��DEg��_�k�b���4�$	@�6gY�����l����=��[ʋ8YN��{)YG���of��v8I��D�=,fbs�� �����$��t$�K4��_|�k�#~ك�},=��5�m��u����T9CLd�tг��U�G:K����2�,d�M��p)���i�o�a%�ݗ�%Rك��n�-�*α��_p���d�I�R"����̇����t'��-��-�Fy����>S��o2�o��ap��.F�[��%�]J��\Yg�M�tNdw�5��l�+�vs��+c���"��e��ͼ��;[��W"�lo%��#�W�.�}ꮟ'2y��X�j�i���V]����~Ԫw�U�J�ʨ̟�ͪO'R����u։;�s�	ʹ�q�զ�W�]�S�6�������_'���gu1Z\ٮ���:w��m3��YW�ʙ0/J����7��{_���'����/vs3Rn�ھ�sF3�P51��B�F�q�(d���{�ާ7���1C����R��)�����/&�y����g�[�5-2����Ǖ�8�N�CͿ>t���l��+f���35�Z�x�o�Oz�[OAW�3�w�/fB�z�y�3�~``ɉZN��mbs٪�'P]h��l1{�N�v}��[�KgPA��f�)*��\�{Cf7%�8-u'K�� ��(N]e@e[�ồU�������z��|
�yh�⛣!`�[��D��YQY�ظУp�2+�]�u����;�d$l�`���ܠ{�R�G��²��x�{Ei�ǐ�h]��(�pz��s��Eb��a��\��[�B�بk�����o��K��;9u�lh~�*yJ�\�)����d,P#�����촷Pj��)�v�\����K&�w��]AZr���\3cq�cl����Wt����R��R�	�s�N���[ݹ���Ԕ�T���,��d�E+х'��~hbb�;ӕ��4S�|���Z_��ʇr���?�PǓ��9I�����s}4���)jh�R|���3�/���yކk��j��vf�9������.q>�s��]NKg��#7�m���*�u;ɺ�Lm��I2�q��V?%3�j�.Or�t{eΨSJ�n	�6Z�W�-r�׻cj*;t����W�K��x���=Xs�D�o|.���iK�Zxc�u�����ޅ�����5Y\�ō"xg<��;m�]M��t�/�a��r۔�q�M!0�3w����r�V�VO>Z�Sʌo:�zu-��떁�+,X����'K�ru���B������{�޼P�n5���,xnm�[i�{9%S�AO�vÊ�������5Ls�������l���2�Ku�lo�-�6�{�=���/n�^�1��U��[nV#i�Z+�Õ�c���[Yn����'���ʰ'��o|�n?r��~�7hM�Of�Ec��YVЖ*��`�vN��S��N�x�4d5h䕎�6���JZ��~b�}��J_�����Q<2m�8��	�	Ew-FeP��:��0���,�HT�%^+�3H���EGhJ; U1j@����:wf�8�u�Y��C��ԛ�.��7�Q�a��ı��8'�m��v��J�ͬ�)6n�N�ye�����w�P�M�:�7:��~z�Y��΋w.R��A��N�_Y� P�{t�K2�e�,Y�;m�<�MrQ۸��J֌5�wO�G��[km���}�����;�vn��ڀ���r-����b��@i��R�u͊�����~oR���XR��������T:��k�+�ok;~�Y�O��Ԅ�o.9�]�xv"�3jV��7�օ�*~�S㳰��.85zs�\�>�^������HՋ��el�|R���;�G��}�u��v�<B�U����r�4v�-�B�:�|Ij&
bb���=����n��oU�qy�Ov��R�qF������­��zm��̖ۜ�Wn����oT6�^��xs���cb`-�����,Q�{ۭi����qYŜs]��T=\��c"`n���s�ɨʭQ3�o,�"{�}�~|�y2�7�m=������3����8�=!e`�;�	�̙��Z.�+i�[=K�lx�F�X�E[�����VE�dy��Ӏ`��;%�wX��8Ʒ�d�bV9���721^Yʵ�w)oT����2���	a�p��+k0ޣ��j��F��XV��ru�P��C�'zy"���X�����b�6�7m۝��g���v�ڋ���L�ƾv�C^P_Kx1g ��*�?mF%�9)���Լ8��晬�x��.-M��꒵�Mc�*K�+��?��܏O3I�ڥ��bVC�WZ�QX����,��5<��,j�#��!�c$��enc'mb���ѴH2V�\�e���)�*��I����;ay���6��K�y�[T��5�pܥ�P�d���:�c��,о}�Y{k������mmM�~���m�;�={D&�:�5�������p�(V��a���T�ev�OLl���&fC�۬kr
@-ҕ�����ㇵ�:��;��m�<[���@o�.6���v�<ݤ��"����A^��((:���i�j�I�v��{b"��f] �ąV:��U+L5�m��+�Y ����qa�FN��qCH.�'�7v"Rt�Y���Jᣣ��Mؽ2�?�^Y���~v���4�3�����|�q�p6^gkv���ot��dXiQ�ut���w��S2�5��Z��LkQ}�sV�N勦6R[� �h���6M\O/!��rfԌ澇!b�tY���W.͐��H�)���T���B�OxO�2�A�J�����>��V�Q���*,� +��YU��,F�  \[��S��#���	iT.u7]CD�uP�%�C���v�㰩����{ϰb%Vݛ��F���VP�� ��"I2�� 5u���.�E��z����cj���ܽ,tk'�Y��
��)+;��sn��]Z*݁7�+@�;�wJ�U�H��A���p�S�D�S�ϫ�1ƞ�H�S�B��ƌ�h�>��Dyլ�W�o̎�L���hJb���Ʀa�¸�l
�S��1񭺂�)(j}էyخ��<��rR��ݖ���7��Z� 	�Zq��7�3��َ�iU�|��ԠW]#w0Uޑ#���ir�����t� vU�Н�P���Π\���cz��n�I|E�٧���5�	��a�oN]�`))T����s�G��JVFN��@�)m��W�d�~���O��/�(\)TRҭkhx�Z�i�*Ub�l5j��Vj�Z���Q�KB�Z4�Qr���UR��*9[�Z1`�u�Lu��5���9f���TƹJ��a�PX�e�Q��&\.fS�-�( �e*4��-nj㖮%��[ie��E���J*����AT\�\-r�c�.Z���"�[���4�R�����Y��,DƵ
i(*e�JZ��˧J(��H厖�Z�GVV*��TAUM4u�fSYDEFj�c(�1�#�V*�ZƦakYZ1Tp�b�� �eL�eu�QD��D"�R��Ur�A`�~�>���mq+F��R�p�ok���d)�Q�&{1��p"W]�3\��F���r��q&;�q*�_}L-���&T�{�hS/��̌N����}�G5A:�sFA�+䷔�Ψ�TC��	8|6X>o���0u��]:zjx^-��n�2��'چ�����j�X{�@8�ѝrZo��>E���I��cXꨂ���9K\Q��s�	WN'V��)C��C�r���f����]Qs8L�k���~/��\�U9�'��k�c�=B��S��ծ�I@=b��{��ٓ�m�y��v��7ݜ:r.��r�7)V�۬/Ɏ{Wwo���[~½=kt�{8='�p^�g�ܖפ+�C+yS��K^�y;:�UH�t"��v�'�fS�YP�i˽��ˎ�W25�S�7a>���'��d
�d;�
(<׭��-��^a�M�a��X������v[���2=�RΉ���V�^�Z��r[l;��D��1+�`�1\�n -�汸^��}�zPӻ�}���5(δ��m�?�U}���{`m��1���k<���R�
�oã��{�u�ݽ�:��*-��]�O5-��6�ܿYBW���w�gr�/|�����cҠO5y��Fu#<�p��TVV��'$�����#HCg�=��u�mbs٪�)<�h��{"�[�@�)O�'/�[ϼxS���k-تA����� 7�B��S~�ޮe���s%�j9�Ӗ��5�)`��s"���v㮏s=ӵ��~�����m7��6�Zʸ����0L�������+~��Ӫ��	ED%��SB��c��e�C��O���i�_)pϠ��un}h"�QKG!P�dǓ�˖E�lKMㄨ\�|��cŭ�QJ��taJ�lO��X|��e��Í�<T(K&����B�{�tΑh=�&,�U����qx�Y����C����Fc��G�5T�򇺗�uuq��ok���1�zqw)<�x�.Z���Kw���Ž2�⑲�p�=s���[6l/�1�=�˪�v��?��Z��V���[kl���!�iR�Q�E�rK1�5ޚ�èVg��}0nz�4=�F�,ɞ�ob�o	�g5Ejq�mM���v���ĺ�*���s,=ά�'��C���>E[W�9�}�[����9���r�/_`�]#�fҳ�5mj�ϖ�N�+���+�`�Z��"�4��Dm{����PO����x�f��2�S��V��{ڋ���=�Vr��?Y�M^�9�cj�����-���+�y��*kb�S���֢|�cf{��{U����C �p&b��֭R�'�8����YF'����o3�OYX���g��)�f��*g{��>��6�WR{�F��x"G&^�-��X��#uĻύr/�U�����w��z��8��nؚ���<�ӟ#/|b�����nAZw��8���ƴ����.�es�4��*��Ow�.c}�E��f�Θ�G��nc�S��	j�W��ވ�I{/����.��Nv�<�J���TD=l�\�8FN�M]J@�k�m:�Ψ�2�y�r	�`J)��)A��t3ޘ�l��"�K8x��q.�]:@W+'�y\7�9ʫj�M2��W`��l}+������5Fh��[�>�Ph��;d�Oa5WOSAk��ȨK�v'���k�]"�L�3)����9�_'�+��9Sa��u��X?){����y���sw�'�	�O�إ�nr�!0���{�����������������v���59'%E<n�1�s;~^�as���=u�ٴ�O~j�oԋ~�V�������~�&QN�g3�Q.��`�mU�V�����rKOrڠ�q7�5�z��h�e��o��[�͜�����n�cz=x��u���F��?_a��=�������L*S�CW�.��4ghF�
��Yy�/;��\�{�ꌡ�M.n�.N�q�X �v;Fu�����%�(�c����Ep&g7��ꯩt�{��U��������R�cA�{0)�)���WvRͺY��9�y/W%��9�9z�W��o��1�!l�=��iU4�\���w�^tM�z۾�VMF�� bLt�5�s�I��AO�u�zu]ס>���PU`�oZ�cZDm]��Koué��y>)�L���N��1�ޮ���oF^�M4�ݜ�gj:�Y�	8`l�G���S1��'�9݋]�7��(���%�&��M*�l�R�\F��Ao>���.�;���l-���<�1��8ԆJwM9�Ux���ޠ斍`�y�����S��|y�ME>LS�r�Ѯxr������k�|v�yݻ�̊z��7�u�5�:�Z���]�ì""k:���˙`A}F�a.���5��N����/z��X����m����w��F��墑�m������n�Ḍ�ؚ�X��qˁ��B�ڥk������vm�bۙ�BY֝�����K��c?��慠�E�=�E�X-T6����a���T�N�'����c�a-d���@�3W����ګ�<���Ci���+k�8e�;%J�ԋ�&rSӊ�P��[��LҶ�y��n�:Y~}��:��2)�������swE�k��Ñ[�P��S^�\�9��8�}W*c{:��b�}͹��F	�R���8�f�&'��ak�-���~/�*'�B����}1�Lj[���޸)�p����4�b����a�%��[�����yZTܞO��q��o"���D��������iY�����[X��j��{J�Z��oy�Qx����ܶY��4Lف�����X�w������N�r^�!�;2�{����ښ�C�G��J�Y r5\�Lv֝�%|8I*!e�9R��W:�`9΃ΧՃ���3QX�k�YN��=�ĥYIt�P�j���s���b��4���W'�t�s�5Z�P�|D˛��M��Η;a�Q�s��B��P��ģ������{�w���u�aM����.c9s�w��uθ����;2������i#��w�q��\3h������+�'T�#+��q���g$��P6+��:����uv�]��4S[��lH����w����;}�>�fL��4�LgF�f/�.�i>֓&k2�?Gg�6� �9Uqu�q���y�q��3(�����k|y^>�;�KW��9��6�Y��\��*,{y��O�/W�ޣ�>~�J��:x���[l���TAQ�S�IӴ{���e6q�c��[V�'���ז���֍ꂶ��n	ܖ38������d�嫣S���yU#�������f��(����	���:��>~3i���ߞq�� !�+s|h�,u�k���6���k�[+����z��j�G;\}o�ʒԮ�V<'���XU�:Ojދw6'��U����˨������g�2�j�ƿ������p��Q9+����=���\��sbo?�;6`=����b7�W'j1po�o%Ҏp���i(k.�6�mC�U�W1��exd[�c�~Qk�zn;�w=nL�{WMf����Q�5�b����8tv�;�_nvMyH�nBB���|�����M�6��\"��k��gkk=^ӥ%��,R>��곔g��5��9QU��õ�OK��|��"�h~=�*�ίK>����(Y������,����}�6j��#c$u�U��-�b�����b�y	�{I�ٳ݁:�Z-Wz?J�f:����5Fj>~�Tⶉ� N�u����2Z�P�����u��^�J���3ui��R��n�f+/�8��*l(ov�]���ճ	H��Զ�\M��ِu�l�ֆn+���y��e�� 2� _F�n�!64>�k�}�OB"�f�ܩf�[�]�͉�ufQEL��G{�y�3+q|�-�������Ҧ��U҂Vy����*Q!|f5�������ғ��N�[S&rӨ�|�����|�'}��zm� i�|�LΦ�s�B�����|�v�C��哬�V�=�6�cw����^L�2��8�W�yײy�rP��B6�����W%��}IO��w����}�!ڨ��}G�n�Pi���o���{�f�Һ�C��mL���c^�
`�-V�q��ݕv�s]��;[v�i���(�0�s��lH[BЖ7�n6�kQ����s�݉���_7�SW8+�[�ںBJ���,}ʍ�dsj�{����'���m��u�Z��U��w�O#�fx���J�V�d���r����n�t�ۼ���v_��.鞨u�VD�$�i�g���O[�����z�>������g��������v:),
ֳ3֤bv}�d�%;:h�׳�5�l.��Kn�V�������=T][�1"TC�U����+��b0E�)���-�:�hܟ����̜�#�i�-�f(��_W�}��PΉ1���JBz)s�e!DljtVσ�;Wغ3� `����ˮ�	Հbы=0�5���^y:�Nx����E凲��o^gbA+�̪��@\j��[��>)��1�u�U���3*���)89���j��T�B���Wz��N�⡗ݻ���7B�����&�ْ��t���R��}3x�����)j��ѷ5��e/_:���v����Bx�1���`Oޞo��$�z�礸��5{L�u�����q����jx�u/)t�Dcy^m5p��A��s�j���.ubn����?Z�W.w���ڇz��
Ux`���j%�S��lIʖ:0k�-p��K��ob�y�D~�;��_��f��2�.W�r���u��坛Y%�'�'k͐ůsU�\{)Ϟ
���k��pXi�mo.J��YT�n���;�������T3[{B�Wa�����R��]����*f����I�WB��sE�o�}R�XQ�mQ����p���E��K���SR��t�,��Ʌ+uѠzwj�]���˱;���u�C0�Ek�}D�TC5�j�H�w�n,��d0;�{�J�t�m�ɺ�MV�r��3ke�C���e�,�R��W� ,�ٝ��'�q�)q�c8j&�u���Y,^��&%b�K���u�����3�p��eέ�*��'Y�ԇ�q����! >��8��PoA��B��Bk)��;;y"���<m�֒���*�����2�$�>�s��&ӡ��=7�e�)Ɖ���q�G�j�C@����-��ؙ�G],t/����v"�̄�s,�Lw%X��y��;���i������#��M�������o*��ą�GWWJnF�+�;���̵@$H��8�Jy���ob��q�#e����-A��o��̍�	�x�y�\/o�6���D�])�I܇S��,�m�+K�t���ha2;��2�z�rk,��1���W}�k^Ӗ6�Mi�W;�6�jf�3���"�����Mޞ4�*ͶhJ5�f�:�3��%�m�q[x�@*j��g�=�_�6:�Bn+!�\�s�_[�;nr�X�{�s���Z:�j!��ñ�\�L��#ה�+�%	����K�n);;).B��6t�*�Q��gM�q"-{�p�!��������8g5-���!κ�t��3D+R�6l�w
.���8���?�]v�B����X����׻{2����1�WRǚ1�ZjU�[˄�u�>��\��nۮK��h��k
���s�$�����:�VUD�=��^�s��>I9|��y�N1�}�T���[Sx8�e�S�Ð}��]e��	�;X�pq+��<�k+��3QoMN��w1ag5d�%�V� v�}��H�9�VNn�v�g��!֤,N�G&�(�G��˯S�L�/��r���L˕�6� �� :��r��[[sQ�:SoV[�a�2L���ΎU,ݪ)h��6KPt�r��<��6�1��N.7��p�W��M�W.m���v�@�˹�c�7���m�1)���R]�34��p<�Ό)^� Ӑ�)���s:����z��ﺙ�VX �0�kN�=ںj�����r��-��k��a�	���[�RꕹQk-Lʈ�e15t�V�e5�X�m1�&J(�J�D�t�ȣ�W*���5.�+&�TTJZ�+kkR�PVҋKS�e��2�n[�2\�V�QQF�m�)Q����҂����J�ʪk."�Uj墈���+����`�db�aR�	��[K�-��������"f\�T�"ņ2��b2�MTLJQU@PհDS-U��2�#��*�6,X�+5j2(��J��1nS�B��
jҤ��uj����!��i*���bb#Kb#r��1�Q��2��X
�
Ț��*k�{����޼��^ofJ���{��ͅ��]��5 F�Y�����.6xb�����:Ó���݋���DDC�乢�rJ����0d�.������+J������L~Ԟ���Ï8+s7�lH�cj{GW�w�b11�`Y�Sw�ہՉ��t]h�me�cD���P^��Ǖ����o;z�Q=��G���v�s�9n�E�[ِ���Vri-���J֌/��[�{�^Ǔi�neCPh�Rѵ軻�n4+!)��g��
����pٸF"Ѹ=>�	E%��S�;��38]co�Fnt��AX[�Sk=V�"�8E��h�+�4�7;M�Z�+�a<wT�֡�P_X���c:7�i<�}M�����,�j����N\]~�z���Ӧ�	9�#f��y�&R}����Wm����M\����B��ki!��܅��e���:�z��d������,�t]su��������i��o��Mv��:g	N�:{a�'L�O��ˣ������)���}L��bʭ��Q��z�t�詝�\�Rd��p�[��}_}UT������{DL^���>m�+ݨN򽗆}O6aK6�of�l\�rF-���2yW)�j���C��uX��3��yi*s;�rg�O�z&�W�W�y�-U�cw�kc�`��y�u�kT��NV�
�'�pj,�1|�z�Ls��Y�{n����J^wM8݇�~֛��F�{!{���/���c"����{wx���gO�[��סWOsl�h7h��ꮇ*񥍷�n��=~���f����\��YF9���I���Вt�7��H���S�YPyLF�u�J���ޥ��cKK��T�R��e C��U�Zcد�{�k�(����Gˀ�jj�5=3��"|��%�H�vı�h<W�_GC��_�[.�"�hEu֕!{E6�cCt��r46�7�k):�7�����_�p8�����=��ǔ�<@�o��t�O�����x���⬎������Lxz��v'#7�R�	b�Q8��u�G��G��y���
�.���c��}>�d,�cn=t�/�S1H	A���Y�y7����jܸb���1�g��G3U?rYۇ_�,�'K�5���5��r�T>��B�#��f�5���]|h^����K5����=�뙊�M�jb}����;�֬5�՛�{w����P��^��-uE��nr�!*�ˎ{���<���bMX��ȱ�f�en<���[��is˭k/Ӌ�z�3]ܛ&sj�*��^t(-��e�\��K���~�h����b�֟ok��..��\�c��W]B�ss!t��&�Lꬬw�ЧNݯs�ZWZ�W����8ѯ:�:M�]^R������.b����v�*�'��\d��vNR|�rI��Q�̩�������M��U��+F�k��=Ir6��w�GhТ۹Mрέ���5w���j*-���K�7�q�ɒu�����i�Tڴ+��ǈ�t�]��z�R+6�8�|��I���Dz#ވ�icL22��s�λ4��TO=v�!P����yg�C].Ja��GD�{!��K�Q:�V�}�;�������M�=��N_���T�����U�ܘN����o&:�k�׵3�jGu|1V���B���M��u>�e�#�`.Kѣ6�����t|��[�flڃ�▻hE��[e����]ZJ��	�u�Z�Y�Д$-'t�#)zޯc0"�Wo�n9{�g[�Uv����u:�ox?h���+�h��ˡ�8m�#���������Pb�9{�}�իZ�=�"�>t�{�b�x^C�hY쳻m7{c��Ʉ#o�����<�O[���8��Y�:��=�%qׇ�A{�kv׃�5Z6�����ۣ`.��7�:>Y�/<=hjw:�&ky�fM�ϊ�a��Uc���ۂ��Yڝp=JDҼ�/��C��d�sKb��]a��n�%����[���{̮��Q0odrd�X������N欺IC��z=b<�~GG&�'�[��N!>��>d��6w��zï��>$��z����ީ'i�&�&�Nٮk|����ϳv�N{��}�^{�o��6��� ���$�OY���OX|���c	�{��8��u�`|��O��a xì��I<d�M��;#ޱ=��]��GҦ�^���f���9�	�!Y�8ɴ��w@�N$���M�m�m:��i8��ty��<v�|��	����O�9�1���l��햳yY�~��"#�>��E2j�d�!���>d�2�a�&�Rtw@�N2}�;���M�GT8��4s�C�{њ��DG�=���9��vL����5���,���O��x�-	�x���x���$�T�V�6�����&�8�����l�ug��'�?��{�/ t��]
/�1�cޏ�� OXu��I>�y4��Cl8�d���@=I��J�=a�o$�+	���O�q��d��l�����]boY��{�=�y���|�����hu����!�s:d��a���q��d�&0Xa�+'�Xy���z�R�%B��==�%��!k����|��g���" x��'O�̡6�g�8�q&�� m:d.�O��<3xt��>N���l��m�VM��R$�w���{ߏ��}������I�Nk�'�2Mj�ĕ큮�6��O's)�L=���|�G��2tޤ�3��i����1+!Mk�ߗW�5�}w�>�Z��0��Ȱ4��'/��I�N�{���$�wՓ�+�������L��f$6��l��>A�� x���ϼ|>�"mL�	K�%}��:�KH����,���A�{+��N����00n���f1`f���r�E	R�h=83��l�B�E�Z0��;�V�:������p�ݝ3�w�=�G��yIos�ճ�1�����LƏzAYSh&��te��OY4_0�h�d�wI>M23����T��>��řG���N����T����~�[�y�*d�Vs�p%I�>��������L{a:=�*M����06���<�O�2��'��	��]Xǣ�"�ƾ����m��[��A}� $�=�C�O���xÌ�2�>�*N���;��1�P�0�N��
N�jZ���>d<2���7�G��q��O��EW_��1菢�m�t�ٴ=Aa;|���O��5�xN�q��;�2C�OP��t��c|�i<q$׿d
��ċv����5��ַ׺�����W��$92���u�!��m:<�2�8�d�w�C�M�`k}�m�8���������s�O�Ƙ��l�����Bn��K3{����9l=d�&�z�!������îX!�'��d�i>N�C�i ��2|����d�'P��0=a�OW�|׺�߽�޼ϻv�m'l��ɪI�i�E�����I�&��P�'w@��>OI6����>��>}q�!�{�=𭓿l�G�R{~�߂i'o�s���=aџf�П wl�J�v�� �E�&�yd�	���M�q+']�6Ì�'i'̛Oy��
�p��}7��ԠwލG�c�GL�h'�̇g�dXI���y�C��0�@촞��=f�hN!�&����K�'XMZz�l��d懽�o����{�|�}������,&�6��Xz�q�����s�,'����Y'��0�svB�����=g�����=MgFolUjي�������S���jm��w:xjwexAgWy\��ui�N�5�t�j���vgZ��N�0�#r&L�۶��"9֤��Zޙ�d�L��r�Sr�Zf��_k�S,>�1�a�3�_}_W����}Ͼ�}��=ea?ɶO��:�O�=I����!����x��|�}d8��Ι'�P��
�q=��:d����|"��G�^��*��=��ws���+d��%I>I��9�I�Y=d��I<I���P�@�z���I��E��\���#���{�a��zO�,}��vh����~�޵�p��R���Jɴ�4e!��<�2w��q$��ORW����I��w2��������>����c��鏖�4�7~��k}�{�'�zÆ{�H(=�I1�����VOR�є�=H��|ɞ�;I6�꓌��]�|�Vq4yOC�j}�1'���+��ݩ���p�D|y�P�'=}�qXu��I�$���ٓĘ��k�d��&���'�5y�0�`u5�'o�'��Մ��<�:�\������<���$�S����&kL� �u��C�N!��������������&wa=N2VM�$�a����pǼ�DV�L}s�m�ϒS��OhM��C�ć���)�XI3��q���7��'̜J��섬<a��a�Xo�����N2T������̎���6��ۭ
��������C-�i�	�:��v�05��$�'S�AI0���e`h��N�q��S�s$=@���a۶I�<��*~ٴ>w�{��ǜ��4{�z=�G���N����h<�|��Xx�@<Hv��6�{�$����M2OX|�c�z#�O�{��.�O'�N���g����|��'l�!��0��	�'~�Ğ��juv�6ɢ�|�;N���!S�1����2q:��6��h���_|n.�n{n����h�^˜��U�F^t8�%+
a�ct1���o121Sfl$]�'r���[�p��+$�9����&g�;��X+5�����4m�i���]��
%���C�����ݸ�J[:+#c����ꯛ��Sp�����ެ>�~{�b����"69�<CS�a���ĝϩ�O\Bz�wa<M2h��`�����3�� ��ԛd�}�{þ��μםy�<��I<a�6����,6�Ǵ�S���'z�ÝX`x���6��:�ɴ�'n�a;f�j���mg2O�P�}��5��Ҩ��WZ��*����c�G����=��޲������$�:s!�&���"��N����2�&��!8�ݲz�$�����y���s\����:�Ϡ�����I�T�}Iěed��&ޝ�I6��h�O�o�I��C��dY'�5�0
�3|ގ��@��ts�oG7����}��{�b�Y�Bq�5/� ����&�XE�O�7Ձ���l�{{<������$�C�[��OG�ތ����y�#��fY>��_|���
�9��i���I�+'�,դ6��Gt��l3�&�����N=�ui>d�N�S��>`q57C�ԁ��~���bJ���sܬ8�_z#X��蝘��	P�{�v�>O��l����t���T0�!�2>Ұ�@���N8�>묓�O<�����f�=7�^k��|�y�g�wמ{���d;E�Bm'7�@�t����'��xt�I>M�N�1*ɻ>IRm�e �%�4�6ɞS�	�!�~��#�r���?__���x8ua�$���	�X�!>I�o$�i���{�O�������:>�;d�VC�|��{�'�X2z���������s�IUL�#ޏ��XB=�({�Wl��IR����N�VC�O|�Vm�h/��%I���;N�'��1�ޑ��ad��e��rlFWgmuŹ��}K�-�A_�V'^��%�.��4@y2\ٵ���x��̅�x&r�D�����W�vt�ae��3����Y���wR��M�j�D~R�͋;��QH8.\�������UW��H���6�+&=��L�;d�'oFy��`jg0�> �':��IYS=�m�`w��>Ad��O�q�79�����UQ�%αu���ʶ~�#��=o�<I��'S��%d��d�l��a'�2���hm��1��Հt���0RN�5��O��9�=��g^h��|�~��s^p�$�'���i��o�Y&!�ݝ��l'�X'O��'̓��2�a�bhw<�<CL��]�{�"������~=�S8����у�����zʁ�}�;I�'���s�!�M��|÷l��<���8�z����'���I�y�i̲c!�>�g��7{�|������c�{�=��|#ܝ}a�i�x��>Bz}��>d��<��Y=a��ϟOY;��$��]X��Gz����`����ߦgN���UC�'&Y��q�]�ORm��Y$���׶M0�gA�q�������!�ΰ�<a����t��N��m�	�<��o��<��q��	;M2,��7�',����6��VN��m'�>g]�MOl6��6�Xm'���,$���9�8�Y����ν���]�<�a:@�O��:t}Bm2j�d�CY�I�I���|ɶT��m'>�<��2m�:�����$����K��?ER�}V� gu��������,���sGL'�x�Bq�2j����$�{�q*H�a�M�<���&�8���|ɶo���:��u�\3�y�5��y:{I>C�^d<I��C��'�7�p
�a�{��!��F�8�d���G�VI�5��Ԭ&ަY>IǴ���9w�[Ϟۡ�_t��w��f�Ѹ�9�R�˃uw�[���*S�
Wv�I=z7�4�5���Y�^�3��yq'�
��p�&�]˱faر�綂���k�+�v�\{��C[I���F�KJ��fv��ȭ���$&��������u��;d�i�<�>@��>�紓�g���!��gL�Ԭ:��q���;I��q
��VL�6�Ԛ��k�o���k���o���z�$�Y&�|���l8��N�S��'̇�q��N�� m:d:��L'�Vt�$�<7��c	�t>aY6ʇ|�[^s^k�k��Ͷ��&2p��ROY:׹'d�5d�%{`h���$��w���'��a>I��2{��I�<a�}�H,'�gC�;���sͼ�W������;aY6ɩl�zɫ�t�|�ѯp��$�N��q%}`h��gvC�'h��6����*3�D�|���z�>X�Ϳz#DG��ŏX��3�f2bVCA�>@�6���>d������@�s$�I�wՐ�`k�>d�*m���^����Z�����!�M0Y=��P�'�Y�hJ��9>�����S�Lza<��d�6���,�06���<�O��N0�3G�'I���/���.�*��7�诼���D，F RL���q����Oq����s�	Rx���N��La�S�L{a<7`):|I�@�ԝ��'̇��޺�|���{��w�8'l&���&04�2M3l��Aa<t�m��XwI�2p{�ﻫ��5xg����v*-e/��w��79^X�DaZ�^.|���N�$��9YJ[���X�rsq���E����P�:��Q�g�ե��DmfK�3��܁�,&�ʌ�[lcw{\9d���]�+e]?�����lm��i�9M���N���WNWE77ttTj��fq�uX�p�tT�+hI'7�j^Di�FA,��ɊEνe�wRn���˻�n����'�'��&��\�Fr�ͬ@fi ���h�XB��n5W���<���2���Ϙo�G-�q�(ͺ�gd��Ă���Tt��s��02���R�����3��.DN[�I;%;��,τxLVO�#p�zu�N��CS3)>�5wv�fU�׹j��D�U��<�Ԭ��B�jŢ|#�k�ڭ�6���UqVKCy���7sD��y(��`���p1�iGۀ�7�xN=�6�h:��¶�L�0vP;�E���ڰ�k��
��G3�,̻�ɔqMYr�R�l����s��A����f�@G&�ï���a+8�SU��hj��ᓲ�f�nҼ��Ć�bek������pyj�CA��aɝzH�X�JZ4�of�,��a\:�T�D���,nJ]���5�u��@���>�:O���ۦ�:��l�]���4��r�q�ޢu�B�c�F���;������n芷,u�m�]M����ݼ�2���\]�?��aw,WfRb�OM���t�#�����+���iz���Ŋ�^_iN�cH�c�uB��,�H��D:�Ce������a�OM*�_Voc�}��}e�@��_T��e���|�E+�*U� 5���ʀ��v�m}D�q�8nSf�彲6��L<�8��X����we��f^��[*T�U*��5�r&�P��vsv��b��9@vK��Ӥ��m�P@��Jq�gIөd�J��JQcPk��V�����))��������w�'\��k�z��mGF�GBz��v��2��wt��z����!;���F���VU�|��SQW,�q�s(�,��yA�'�sO�����H����8��-u˝Wm�4��㴟~�n�k�]<�t��1�n��2{e��Uu^u����۹ralS�.ɭ�#����8Zˎ���<K�����,t��<h�I\Dv�0��+.����+,uG��U���]�%;r݋xQ*� ��IV`P�Gl朴d��^��f8��6�YwB��ܢm��U��
�u�w+8(��<C�zNm���d=6�Z|�N������5��8�����֤�����KN�W9kNZt�v62+�G$t��3��{ٗi�B��"
��bc+
���EH��Dq���̥QV�ڂ	��E��
�X�*8�1��+�D˘��Jؕ*[ET@P1�A\��lq
��*J�11�S-��
V�-�8�q2��J�H�-Q��PY�[b��IR(�e,�E++L�*\�P����ٍDD�.q��X-ƆV���Y\f2[�V��@ƥZ�2��0�k
V9B��,�*���j��,�[Unci�f���h�jT���h�Z.0�B�ef%f7-�)���l*b-E2Ь��S����J�+� {�6F��Ι=t�lf��U���@8:�ŧ;37���@�2�-����2��;Ͼ�����۩���Nҏ�wx3�d�$3�IP���;�����T9���w\��^�Ej��釮q�cJ�4�&�{����8�P2zPd�F)�j�hN�y{�7:� -<:1D���s��L;I��hJ��<gz��:�:��ߟ�ZӰ���KgB�r9��!��D���#@�P�_�����M�d�����D�����&(��7�/6X��J
���Lq�U 1>Yu03\��	��J֥S(�J����p���3�)ʷ_g�0�*U��u ��/v�q+ڷ��ki(�8�AC���	�N˒��Iڍ���a�dSɷ�[ar'5m�qe��JT��	Ã~��r���o�ptf�x�F�1�u�'5N�1���Gq"4�C��BB�I���z$�4]�"��J�=�ƹ�]p���&v������t.�3�o��g��������>���t�0n���Ѯ��Û]	��[dL��ɬ�l�������q�+�{}b��tuM�P��Y�U�}6�wV^�!8��J�>[��|kFã�[tfvټ���kn9@��+���LJ�s>�v+��ď����Dc�K�em�J��*M�4���*��m�"&1͂+�Tၔ&zƸUf,m�eW6�ae��z|s���F-�Rɯr�e��Q�EbG�ؼ����.��eh"�ȑVı��J�CF�c�3�("q�#��f�H����1��9⾤)������bcjy`�Vtv#I]���3Ә�{ܐY�5��V�\���<�֔�y��X6��S�ph�PIj��t��o�x�<vP�LC-�A�6���c��v��+�*�j"�*��Q���S�Z���d8Q.,�*�*�w�Sҧ��,^(nآX����-Kʼ����]�kBN� �L������^��Mu�:[гK�*��#X��^�����~���_�<>�lՏ���y�r�[�dB�i]S�o��M1r����?n{�=��d�8*^��u���`��E�BDpY4;�(vșA���CЮ�P {g�����0vh6,ψ��v�X=
�
uJ��7K�u�����֭��V|S�z�����6����jl�|�̶�4D���1vd���SGN��/6��J8�VB�.��D{�;z񸮬Q��`��'y䮥�u	�o {��1Ƹ�`�O��wD�mس��u(O����:���?��o(����h��t8��[��*��h;0�����%�c.RyR���Y�g��rL�1Z�M��pk�
a]z�z���\�11j`�Q�@�q=R�������p�j����Xq]�V�&&�`�jHWpe�~��+үn.��VX$�)���N���<�a���o�)�yWU!��57`|��8|;�mCg.+�B���G"ֹ^��m�5� nY�>�Փm�,p�Yg�/��-�a����N�s�w<�J	�O�aO2E,�o�a�p�\��ufZT��٦8U�Z	�8<�5��l75�Ӄ�8vu�i�
���]O>��9�%�<����[��[��\#ml�or98P��24D�uW@�ɘ�Ԩ��ō��0��1����ݢlh~K�Ш����)��4?:��	��H�xGR#� ��1;�X�bR5�]��TwSx�~�grU�8�=��YTէW����iŢ`�X��e����BչJ��o
����S��a��>��c��K��*�_}U� �OzS3��u8p����"�2��j)�!�V|\^�����dZo6���\��IwX�g�pt��{I����t[ۊ����ݬ�#�̾u�S��5/v@zb��&&wla lzn ������Z�.����*�BO��E\hM:Ю�.SB��p8�eT�Ã���%N��תʭ���w��:�Ղ$2卸��f�*��.]�ek&�8	�t�����g;�"FC�;&:����׶e	�,1t���@�OU�Bf	_[�C�R�e����K��'ԗt::�Ox�tΛN�a�]e%�ަ:U�W�U��ƚǸW1�zG1�)JY����T��[����r�N�ac(	e�[�S�j�<�����@�+�E���-��\m�^yP1�6�5�,���*1I�3���*���|�B4���rG��܂��Z�Z��<}><�, ���6z:���
�@���r�����)�B�JL�*U���-��U�A�+�"�s��g�[�w��@�n���S7DC,��;����W/�FWҺ���O���|�,�ȅ���.���}L�����;6��L�oJ|�����މ*����ᱯZ����l�樍�ם�)�NL!Xx�;?<�j4d�NՕ����~K����98*�5��>��h��,�y����͍u�d^�ԋ��uuMk�֍܁	�Tp�ʦ/�1����Fˣ�Q*�X�p��h����:�8=5cN�T�<]�V��A��T�*�yX�O��w���П���L�k`F��IuY�ș͊��D+U�=�X����2�'�a�L`�9mT�E�*v��;�?E��o���H^�_�Fu-m�K��#ad�N�3҃%�`K�W3��.��wo�����i�1�Q޸����S,-���VR����E���Mgxa��~��J�P�ЅG'\�8g=�%gU�0���A<��)y}��wt�cr��Lz�A+�̍�=5�H\R�)���j�,c��	���o�\����DC�>��E��	�l���u��L�"�u������(֧nDR����G�k#�4NK!ٔ����� m�~��1r�s(�H
2#�8����ē;�`�����64���
�'R�������$�8�n,uq�I����>��+G��U}�}�Wm�]fL������0&9�h��,�	�؀HK�x�W�e�x"���ܣ:4�<��,e9zn%�T'S$�qd�5.xTA
��I`�Z�W>��K�����`[��r�[@]z�S{-uT蕵��N#(��'T�+��ϼUvvO�E�� �q�x�%��Z�����<�gg&.9�Y/y-!5uA����sz��.�� џ-�5J�8f�"1�F�s�U}�4�U����/ؤ�v
,�xc�YӔj��3a��E�|�e���b�sv�n�f��0�nY�X��x��C֭/de���YTC����U�uMr��Nfmf-^�I�|wtf��-ұXD�,�*�Q��&6�y`��@�%>��1��%L͹�Kv�L~Y]��'��r��BiE
W��b���.e�P�J����OiPgK
�j���qATd���j���^�ٞ�.F.K�n�a����5�m&�� ��X���!��yJ�s�Y�V�o:Bm��8�5�ã,;o��++��好����{[����z��¯[� ��dƟ+1S��%؏{��xAc��Mf�W�W�KRM�wgf�]~Ɍ��	~ʤ��TFʮ��y�n��]�o^>rgL�}���i(��L�***�n0�����[�b���#�]W��!�E�-�����$S�oG��#i�,u@>�#��'��Hs���6�ry˽�@�LJMu+�ɢ������f�8-K1�|�p�=kϧS�y����d�3���jw�!geC�)��u6�������6�1ƹ�OB����Y����u�,!�fxlІ���]o;@���h���\��k�ʑ+��N����È�� ��S�U�7��(Y�7�|�>m%uI#;$X�תz��Qd��TJ�� F�����EƟ��S}�Cu��7�j˜%��B��o�឴@F;�:��)+��������NR�u���q)�CO�%/�ۑ:�Xu�Dc�(p������bB��`,u1�1�h�&�7�kkwUCo�;!�u�_.�{�8ΎNCv�؝��\mm�ܿ��O��-��o��,o> 6�[����� F�Z���A�ZVDF��y!��}��+55N=��r��V.�=芥���hF��p��,�,+��Jm�e�8},��ʕO.gtK(n�������>{2��{D�Y��N�r�F��Ἑ��'PB3����	��&�Z�e���92�sOh<B�Go��L+�A��:;x�>{�� �7�@"t]�~�~�����0 �*���*(^���a'tƊ�Ȭ�ݻ�>�k�zH�}��Ыǀ4&�E\�0�mB��OK0�3��e�M�g6'׏U�U�N�zP��TJ.}'�q7c�Y7P��ܲ�i*\�Ψ|c5M����뉉�n�$�M��zY4T��7&���FWf�$:�����+C�/���w��}�R��bx�1b�wm9�9��y|�K0�ne����(JR��]���*y��i+�n6�G�A��
"�YJ�v���v��s�\5�p:��3���"Oj�rbB����l��kE=�a��YC
�G:_B��]v���%]z퇔�ҩ¶ݸ.6q$�
5�%N��+/-���x��@,M��ǘuv�\ˋs6��Cw�GOI-��c?�������MC����t��X�u0��3G�MA��ܺT�T^mŰ��.FQ������Y�ԲS�<�D�b�x`gѡu�Z:�==`38Xss��u����;^��(��nIg��F�f�øG*I�k�"�4<.\��84�
�gy��z'���`��@T-��I�^O.��'!�\����g�֬����oB�ٱ�ٺ5jpR�LmK���'�6�^vD�'[;1p���2����4*^�w�*�*h�u���zW��`o&M<��npfƺ�2)�f��Ofgv�ї�T�o��j��׃V��Ƕʮ���dT3}t��;X旆�{�/H�@�~����q`�x���V��VPYLp&H�EG*�ݺip}}�Z�E��Yzc�zq�Q]w�(�ɸ=<� �b:�����y�[��H��Іq�q����z��c:W\!d�6*8Ȓ�5�>����Nܛ��\�Az�SJ���6J��5i/\"���:���]C/SZCã\��z�=A�*c���='��4j���7]��=�`;�u`F�F�KEEa�Tm����L����t��J�7-Lˎ�	2����UW�JI?jX��9���oi琝@\A���9ϛ����:(���+]������ڙ���0κ�oإ��(u(�둇�D�����@Y8�kvc��׋�^���R����p�y+�'x�J|�=�M16��_[+ro��=i��mL'9�4���x�N�+d��Z��5:�bIK�j��$���2�Y��vr�h*�DitW�,^�4 �d�'�v��H�>+޴+�F��͜�_��u�JT�T�JXp`J�< ��h��1��ƀ�̭�⫯0>���bಊ�Ep��d�w�
.��`�T_��{����%�	�n놧|�9�F��'y�5�܀_z6=�V+U�t!���m�������Q�+�%%I)�N�j�cS�ǂ�5dGP�k]�>t�l�<yS��I�� ��l� �W9F���3a�����)%��2Vm�2{ފs�������wXޘre����;�"%�Qt��`{Tŋ)��Rr�|�(!��9Q2k���;�ׅ�fd��?��5���_LL�Q��:sd�KxU���w3�v��U��KI��	t���p��!�m:�ӗ�EKu�Τs�<U4�2���I�"j���T������]d��k{L�X�Gr0mc���e�V-n��Z����,�X��Trx�_mc��q�tT�m<���.r�8i�J�o!�wy���TH-h���m�s�Tx�Y>���]v�6��,�W)�&��'3��h�2n����|I��Wdv��i�Qsi���{�r��Q]#TU�qCW;���ȩ� �����ʗ6g%�6uHs�>4���!Wfu����mL��@�[:�d�N6v��'/x��Z*^^��]��J]��[�J�Ð�j���x7�7�X�����r�i�5r�8��ƪ"�mX�b�j�N�/Qxk!IaV����x�̱��=�@��H�B�J%��Z{ae7ady�fcI�"��.���K+m_�����;75w ;�wH�Vuӽ�V������}�̧h�'s�͙���ԬJ�9YH���Ή˘yeC��0.a��-f�̥ǎdG�����U����wQ�5�j�`�{���b�Z4©_*�/}��|�ǵ����I,�rV�bJ�0v`��e=ؒ�W+z�	W��٢TW��b�ٔ�z��;�d-f�������,��;8aln��Tm^5�ʚ�bI�5�u��M���]�5�r���Mn���K�X�c��{2��s@y���@�v,$p�vxi}�4����p�)��M�>��;��k���Gw��r�ѐ�t� s�ch|��&�r
R�;��*���B�dܸ.���x�m���
�:�r���H⬑�΍�*�a�|�Sq�J����U��gE���� k���Y�M�8�u��ߟmAx^�h���ѕ�{�Y{��9ړ`NVW%ozb#x����FB�'�� 8����6{}7�R� ����;��_|���[��FkU|]g$�˩�WsK6�L�ܱ�+Zw����	X�&���}a�����x��{n�ulGU�ٰ�Q�{�r>�LW}��ɽ3�AG4�Y�$�ˎ�V4�J�b�Y˄�$����al.<�U������;����?
W�|c�(�9T�̅�V�+EB9h���ز[`�Zȥh�D��Lk1UJ"����*���R��B�K�\(��[k+)RЪ"���a1m ��[J1��EF-Q"�cm�P�T��V��U��0��R�ic ���,̪,�"%�ڍ`)�f+l��%I��l���R#R�)���Xbb,ƹs+R��kle"QZ�ferŪ�"�FڅTQ��L)Q1%IEAh�-����ʸܸ��b4�ԩ��YZ�A�
���.Kq3���mJb\b��̥jVbL�V��E1��R�f\e�Z\�Aq���LnRbG*�,\���fe0 ������h�Pwr�|>⧳4��oo�p�چmư��cN:�����T;"� �Wg/�m��<2��q����z#�z�"skl����F�ޞV\�;ȉp.����Ba�Z�Bݼ�2N�*�Zy��
��3�����s��t=5`�k	T��C��q�bck�	�rp�S�ҫ�,!�X�J�e쵳�O,�
>����P�{�p:-��0�d2�[;�Ot�ؾBU��%�fK�L �2Pxm�O�Ή]��\&3pS�p#���r�*��pY*� ��L;���)�Tl�������X��֦���!
�"|�� �LLR3gϞ�/J�%*�u�4w4�]S�'1�@��\c�tD.uHirGx1� ���I��m�8o��5�^c���M�;Y�\���N���[yP��z&LȾ8-Jf<o��Ǹ+}Q�y�W��N{u�w�+YNe���qR�3.�I�j��{r*� i$vt.�t�/�<��%�v��Pc��B}�Xu�����o���4���p�&�L�.ҹf�����S�"�^�-�����˨�Wp>�G� )o���8k�R1[�ѱ-fپ`0��j�㊡9�jk.�*G}��"*��#F�ɵx�1]1��ڮ�ť4��4�fRu�6!��n1����UO�����=�t���T'��O��xpk�d=W�mB���N�ۼnr7^&��6C�GmO�Ѯ�G��l�]qx�S��>�Gl�TUL9Y��V��K,����+�Q
��!\2�ã)zd���|=`-���_�����~�ܫe-�T���r��w�Uu
������(�B�e���b��f:�禩��n+��� J���:�' !�c���e5/� �&Vw�Y����憼Ⓖ!�Jq<(u����}���!e�{<ܠ��M4��J�y5�p��
lP�n^{��KAA�7��
�ӗ�ɫ���)ڭ9�r�v�,v�G ���`%�gQ�X�Bq:�@����Ժ�/\�
��0�'��\����M�n�S�n)U`pܑ�8*�pa .����8'Qݯ^����o��v���u��a}�>�m�E]!d�7Q��
*%
�>�Ҹ����ٞ�����"�u�K��(0�H:�[{*���i>���ǲH��� \�U��Q��Mg�L��E��n�����cb���W�E���JZ�A�P�f���t��=�$���T�8S����K�n%.��o\S0���pay7v� n�1u�j�fQnhGS��e����k<�"�ل6nps�O��3MCX/*ݷ�1�^��oH
z��>�o�\�6T�:�X�\���A׌f�+ԕ1~�u��Bɂ Q�W��^��%���,�T�-F�T��#����!�OT�toSO��h����n�v�@��JRx�P�u]s5G�MaA��ؙA%uЁ����=h$������5.☸Su$�=�
(�o����m��١�7��l�S//���!�Lؤ���ẍ�Q�h�I5�rDX���9<5�qV�0T�F�Z����A��Q����=�9��O�����dvL�����B{�p%�G'E�&�N^�P'jX�W-���E����d�9C��ժ,н�'$�ĭa��|2��VT*������S���K%�ϛs�;y�"	��
�4HBi�E�+qa�b��(Q7�KR�o}�6��ׅ����aI�T��[�5d�I����m�;t��ܩ���+"/}�=��X��ˏݹal��^Vm��4{���$oH�ꮴ�~z"=�v�n��Z�#/fG��͐#3B9T���`�Q���_�R%�#]����l�ͭ�	T�����ܝ�<pn���j��Z��$V�W�/�Ԣo��&��B;�)�y���hG�nX��:�y�t�TmOo��.��ܸޅ��*X�+L*���o\��9�a����\�ب�"J���t����n�Z�r�S��x�ʢ����$-<.#Kޜ�>nf@:N���2k����B#&��AQ1>��ɀ��;�X�w�t!Q��#��Ci�\)�ssW2�rƹ�X�|�v���98	�y��+}ei[/�fz���е��*A��U�Л���Ns`ic�������Fuúz�*_����\�;�C%s�N��'���::������Y\>CG����Γ���u4���o_[�:E�I��;�g(�w��BսS�����O�V6u�1���[a(��w��R�vJ��R�iu4�0õn�R�;�x��W;���m^=kȱT��^�����sS�ЫXlR����4�m�̝�wL�\_E���I'+t��{$���f8L7�~����K��}��ؙ:����,Li�0�H�{��۩��P�p
uoEyR0�����痣�)���f��	B�>4N�6�V�"�t�����94��솷*�n�Q6��UzN�EcW/G\h�Ţ�.�(��S��l�M:Sf���e�g8�v���k�<�}��e�U�Á�)�
���pM[�p�7$��|x�=Y堇q���\0:�.b��v_Lfv�/g.�y�r�	�l�m��#j9��ΌVE�V+���Q�G{u�e�7���K������x�]w����g���,O,>9K}!4���+p�3���n����}��j�ת)�Ru��Pj6�������T��7~�#���u�8��^�E����^pa�Z�>�Mr�.�Ҫ���5�����D��h^�ᇊ|�������IX� ��b�r�&�
�c���V��m֬�[�����Y�u2�Q%K'�c���{��p˜���!����eۄ=j�qWkK��4���{{�@�U׍^c�ͦ��u��qjJ�-�C��k�P wW��S�zm�l
�2B73��#L�m��{���lVvk����z�x�7��4#v&1l��W �c�����D��}����%o��OV]�f땝�Tt��0��B
�����8pZ��x��'�*����f9���gs�5��AY�3�R��i�+���ͨ]�Ov���J';5��z�֠�C�*#ͮ��d+��>�Z���3���y���Z�{B����z5ݩ#�n�=G����{E�k��^-��`��Ia��~�R���
Q��ތ.Tx8m\��5|�9+Y�k&�%}Q�XQM�g�ˣ���`�$h���Z߃��/�fP�]ʢ5߂�v���R���9��"��Փ����z��� �=��
wU#�5�7AC��NR;,&ON p�rj�vU�t �؉��1�)���X���UҊY�<K��xz(��}F'�.)u��%Q����3�\9�N�D�Y��N�($k�la���_t��/�d5��zff
�r��ZW9%b�D�Y���t�laT���N'eS�`@��RE����s�WG�sv�n��,�w�[;�.�6�!-x�wt�WB�` ���}�gv��r
�K��}�ͧ�8'�M��)���^�!
�q�zg��R�����J������WR�?K��ռR��H!��a��4JFB3��ɘ�J���l#��\o>�*6ۀa[:׽�Ƌ���Б#:�T%� ��"�*��f�*�m�v6g(���zn5���WzxS��|%��X�0��.y}�F�����*��/ˏ���i�oa���[q^�zn1HL\k���SEګ�!r��i\��o�����p}�s�fL!���J��a��+	u��,��ER�t6y-a�!�&:zY+fP�T��(>1�P�J���u��!��!Y��y���m�#����E���=&���eϯn�>���Şu��r�s;���y��\�|>?S�:K��cp�|]!�����0�mC�̊}O�������d'��<4�S�+�h�8}���<��n/\�Q�}���ب�U|�&�
�F�V������V&u/���B/(��N-�tV�yk��I��)@�cn�DMwu.sm���������P��v3��#{8�Vf+Y/5k�	��V��j���ޓ�z'2+������":	��.����0l3Ta�r��)��`C�_Z:칯�d��>;��g����"��ֈ���.��uu@lp�C�20qߗ?"���s�,8��n�z��5힁;R������j��ם�15�/������tnwf�z���,���Z:�UN�~��~s<׉߽��(�x�\0R��M(\��i2׉�W�\��}~=�Uv&-f]˵y}���U�U1�WZ4Zv�d8��TڥTqV���w�Kz��F,w���t:��d�?f��p�wa���Ol�/����:�:�]C$�	�ܢ&:���O���.��|rO岞��\��9�WT!��6+��#�^��U,�"��]����=��1�n)�lt�*�O���9�Hn�g��u2�U��D]x!��rF�O�G�q8�}�:��B��#��CyJ�{�,��^�ɱ7�ua�����ʛ5��z����t��ٙwdv�U��W�[�u�U�]�f���傖���+gc��r��}�,k���o�;V"g�J�;/�ʳ{�4��Dk�fXP�o�UW��6���x��YC�# ��G�������߉\^dF����@뜱]Nʕz��E�2f]++%7�}1	�W�X��9��V��$�Ϊ'�������Z ��0���Оj����+���F�W�%8{H�!�����U�VJw:����F��,J/D����d��� ��sdGa�v�:�Ƹk]��k��wȏa�xPU؈��ɧ]�s ��dL��On��Z�v�8txW�|��\%[Lm	�
}��iS�8qS;�Xce-L�[+�'��;95>�r=j#[��R�u�3t8P8�R����T�-։���9%�x���w�ToD���#g`<:���~�W���6�\2�(��ӰEUٗK�=׾MTY��4�J�n��;^��^�ͥ엵�6��f׼��$�k��5�ȱ��5D�a���=�t��^Sб���xE�1v`潊�r���݃�(��s�A�]��6ؖ��}�T[Ɏ.!��x7�3��%��aC�X���-ސ�G&t���Z�������f譣fO;c��(�еQ����U}U�I �:0��m�x��w��z�z,����<���-�HM#B����[��뇵��A{�9
2#��N����\ε8kڈ�A�mK��3���Zk++�Gt��8�&0E�e�uD�P ���<��eRЇl��l�l�\���y�9�d^5րHc 쑡�� Be1QG�08�\'*1�����ɧټvk]��Wٲ�[1���������䎠Xꪱ�l���❋��0�mɏw:�v\q���ۇ*_�o*/A��ʩ;��G%	����u��H&�h�c���a��L��o\S0]N���T��@�a����
�>x���w JDn,C�S�־slז�}9����@-��L<��{�u�j�t��aq-�WG���b����^tk��J�M��D�:fENg.��r8k��{@���^_Ϫ~2}+d�X�aS�YUQf��ʙ
��M��Z��L�v>���k����Z}A�b��[@��d��Mn0��i�v���I4�LB���w��97M��(E� })S��JSjV�%��A��iݥ�`b*ֲwH��=��8�m��,T��|nA]%��_�RiN,�if�%U����������tT�oo4�\f�ۻ��mi���^^�[x/��t�f�aE@����h�!VkR9G�oy��+���n�gt�ѽ(�7 ��	琇6��S:Kw�C�s
���n�3���%yW �r��2�W�nH�X�Ӓ��]��)��j�-�)!eH;���R�YEA�g�+s�fAE��٦�FGk�2kL��i�2�m�"�,h{��)��m����u*�4�ƥ�3p�¹�v�Z�\k����J�V��,YjL�zn��*��H�?�S�q�@��n�H/t��� ҂��w[2�$�s*��`�X���62���Rie�'!{��!Ǝ�1�کN����h0�:VM�<���Jy�R�xl�����VN=xL��Yuղ��k��.�Um;R�[)��`��w�[��	�eBf�u� m�U0d�Wt��ˊ]*>���F�#OL�@�@��^�b����~L��Q�A�B�Xh�=t;�359w'gCr�8 ݬ�"���`8����	�6gɐ+mS��m�xE��q\׷e+C�fۂu�f\ْ�6��k ��5�f���%'�{b����˦�9�lP͟(��͕��
ڵ!7���)��l��O�N��m#x�u�֍���� -�W�K�����k//WX:~� _\3f	�[��X�����ݢN��62`��(akK+md�Άxt���r�[�|��]��2��#T�1!A;,Mx�mQ`.�8�e۔�`S�g0뮥n��Z/������o�U��ԩ��z�:>%jEI��)s�ɲ�i]&��Τ(2�8v�g�,m�f�x��۱�VLe�)��'V���ڬ��1�w�MM���X�X�y�W��+��p���2�_d�,NI��s���ꬵ{٧W�IWdi�؉�|&kr��n��Z����S�ك}$t9C;]]�|���U�4�J-н�T���6l�}J�W�����H$N�z������!x�5k��$Kw�ǣQ2E����8ƴ���.O�.72Rl=.��S�Ļ���R��MG���I��Fmt��`�L�S\�9���(����fV��\�*)�`��SL.\�T�q̦ZҘ�iR�1ˉ���R�1�j��
�4��ps
�ȬX��TTm(��V��
Ve�啈�.8�j�%@�.Z,(Q����,\aR����+PiT0��*�Vf\@�f!�\LLkZ�.f`��F0mP��Y�ZK+@�)Ps2�L�b�q�X�
������V��+1*\�-�2�U2�J��[K���.2JT�a�LE���ea�Ph���ffn�3�T��9�Ƴ-��s1Ɉ(a�[j���UJ��LLejQ`�b��*��ejZڙs%ZʌKZX�Ȏ[�am���mq��e�Tc��*��Ե�Ш��(�HV��f*��X�T��
ԖՊ��!Ed��!��e��#"���3%LkmDı }MuE�1�<Y�|p�z��w��>�z����^��D�Sz!�l��:�Ɓյ�)c1Y�a�*������k\�G�ܔ\ZtF�b谉�25�`��vvxT�ۉ���E�޽��m�q��u
6ru:x��=���3u֩{����a�z�t��{��M:�v�`�8(X����y���Y1�Ūʉۓe�=xip�����vgw�U�\8�(TI�*�gE
��8�ϲvR$,�og���s���TK�,׺���f��9%3�ه���U1RdpC]�x+�/B�K��e�U�*���&E�]�o��*�a(9�QZ�ө���gb�tsv+�\�i��۝��3A�ަ�czWe�Ĥ���8[('�-+�ޮ�Ƿ�щ�ԷڊNa~����⮐��ޔ$d(W�����z��rZ�Ꮳ^��h0�m\�(uE���0���HLk������+�H�b�+.ēg'���l��^�&�z}�����789E*|�1�Z^�.��F7&�me��������砸��B�˳���K4ӎ+��ܱyV�U�xr�7�ْVДz��alm����dt�E+�x��ڳtm������򍮆-F�8�}�*�B2� WT�͟�mx��d�F�q&K�q*Ȉ�{:z�iٞRL��%	:&6��q.�X�⧆�A��(W�*b�.��[��W���.��� |��5�=���S�aV�åϯn�:X`�'9��E����[��w��1��[��g��t��K�1��	O|]:gM�g���GV�˃��U��6H�(W�Mg�<%TJ
n��C����֡�w�E+�$ʴ�:�*]�f<k�t� �wJ�+��u-=0��!��Q�,ι���WE �\�=qX����<i�J�]���{I����]P	����nާ
�F��a�s�#�*OZ��xNԡ�k)�q�#Z�	mUv*n����������0+d6���d�dLEtū�G!�8Й��y��EH/
[�k�����+r��gG����,���FT�$.�3Y�sA���H��X��u�E�z�	��������ѩGh�W���~uY�Wd����T�w������{@v�&qoe�%D����<<�LoQj��o-��]e�td�WĹ��Ȇ��v�d�f݃�L�U��GS��_<X��I-��Gt���&��@��ԥ`���G��Kw5눠��M%U�aB9�<u�+��d"LR����ѥ�l#YXy��{�6{�z���*x;�ZaiO'��)�ckҺ�K���z.#�����w�9�Q�=ND�A�q�ʢ���zU����2���~�}p��ċ��dXpHSɚ�a'(ONFl�W�9�R�C��C}��#F��k��6����#+ y[�$��n>f�\�~S���d��m1�;)s�1YU�|���ls�ꕅ-��=��<�ic�v�{	J�<�8�T��)���r��n.���Cj�pt�t3����c���{ȍ.�K�>�r��N^Hh��i���`�Wc��}��@�k�t���9�N�YJ:���wROO�E��Y�D���&����xk��e	�2%l�
��CRi�-��� =��m燊�&�g���x[5,�+��up�i����4���:Elv���	���ܞ����
��+�IU����a*����i�4F`�z��?����!����T:�T��yQ���b��Y�'Y�2�G.4�иۛB�F9M�2"�N��þ�z���T����<��fqZ���Z"����pt�p��]0����~���9 :[��+v�_[�=�dD��#����M���k�q�.7&���Z:8f���H�������,��F��62䉍RE���4W��/53����Fܸ!֯��].��'5eL����9�0��v������EWŘ�ݛ��T�[~l��s����lG*��ZɎ��S��y1����B�z<l=�	00S�pz7��S(������(*�A�mS��dr�P2�
���͝��<�1{.L�1��@��,��<�ɔyLhCM�T��k����;��T�-���K�Ӷ bCvH�,D� Be1QPyWq���V6�� 2�N�j�b5�inc��q1�h��j�.H���}�G0,�����k
��ޙ�o�w.;��1՛P�ԩ��a��LJʩ9Y@����*���i�ɗ6L�z�P��}ys[�ZKȨ�<&��}�H���g��m̫�h���es�4�wvIi�:�������N��G[�Ү�u�	�[٥�'�E�
�p��X�V��i@�S� n�E�"���}��r$v��~0�\:��L��o\TJ��Cۈ;+�ʴ�j�.2��;4���Q ��Nq
���:0T���(l�#����5��!\I�}��ĳ������p\I%n�<~G��U_*�5���֏:(&�P����w�c���c�o��,���Z���=���u��iT�D��_� Q��_m����Ex��G�jw21�τ���Vy�Q\2̥�C�^�+ӌ�,����/s��6��
�R�1�j\4�]ȇf,k$g�ԧ(�zy����~s���q�@�ʞ@�q�J`�w�}�p���ݍe]e��o�	��!�8��ӢF�Nn}�)*e7�������E�G��)V��0���''��̪�A-�e\i�
Ժ;��.������Z�W��"sj�bp��u�n�p��.�7����C�*Y��%���y����C��{�C�����Ӿ+�3-f�����@x�|�R����I��ߙ�[�M����(7���z*���Yr#����5�cp�qҋ\��+7XM��L���S���[��s%j(f�>�Q[i�%�od���tƋ���ѐ���8*pa #`�f�zo�r��]�+�N2�4T5�
�����q>θN؊�WH��l�@"��LƼN���z�՝�*y�f�xP�{qQ���)��	��3ā�	u�v�.j"���xTOK&��p�x;�L!�YZ�|�����r*���ǯ����B���X�ղ��q2�X�*xm���iB�*aN��nNt�r�o35y�@�<#�L򓠴w:*^Z�t���a��`<;�٥p�Z}�5�\�zm߾�sF�N�a�m�_}p��� %�{�/�T������]5Yվݭ�0u' ��?a����t�w(�.��� �\,M3N5��VV���]�U�w(������L�K��|��[�&E����	���r)�Ybf�m,G{[P����Tة�.��7����Z����YKr'{�K�Og��odOT/^ƹ?
PK�O"�ކ�����X�+i�1����V����nG$r�-J �}5�+I�&���
N�&�lH�5 |�z�8���,'{8�ͳ�R�o%a<�5��-=�NE�g�<J�x���bd��i�]NV�5����߼N�Ɔ<�R]�<S}�ø\�/k$Ç)T�6���p�V��XPOUN���z\-\�|�8��%�ey�u�n5�q�{�R+�7�Q5j�θ:V�1W��:)�����&T'휣k��K1��u�Bw82��"��X6����;=xY�xB�s'��.P}s"9��*��U�#Qx[�^�+��b e�0�x:��l�ki��"����S��U�ʞ��
�e=��0�N3mD.�C" \h��ũ�+�0� n}�.Ыa՜X� X�}��ڥ����W΄+0<��f�|u�L��najx��=Bxp.F��R�����T\�Cg�o7&�ѫ]�S��ޚ9;O���q��&���5m�f�\�ܮ�&=G ����*��K,Dy�,�JXn�8��P��G2D`�!�{����]���җ�wi���:�a�F��B����S���;r��%�!Sw���0f�z��O��Y�㬂��Ж.)]��(N���r�����H��oWV��l&�Bf���l�ن�E9�0i�Q������%���Q�צZ;7x:\��:��]�#��Ơ�-۾��9�����R$xܝw(���gOzLl3�Uu�3ԥ�/Jt�'n	E��X���o����[���]�<|�ǽ�>�q��j�u.����u�:C����=[8��p'�{�:���"��b����48(�2���Q}{�ɛ��C��#)u�;��gվG�Dkc�n�5\.��� ��^�;�ʭ��Y�u]l,0�5dD�s��9�N������aGA�ѷ\v�|�U�\�#���5�'��Y�Q�Ek�e.5I�%pJs�m!Њ��YD�r��q�^��a[sQ�J��þ�=�t��h�t�6������՗���T�B΋��t�L�b;\��\l����J��O{�M� FL�z�U�}q�g
���$�\��S��}J�u��\ߎK��] ;�6mu�P<Kr���9�.�u�&#3!ӊ���z�7Nk]���[��,���nynۘ��ŗs!��c��3���qf���ݜ|*��mK{�na�Vd9��C��x�O�X�i�z7%t�8�o?��s�0�|B��z�Tn{�V����Mpr�WT���ƫ��o��(<��/K��K��D�b$ )���U���,ͪ]Sɶ��v��Q�ml���r7��P����5v�x�#�:����b�&]��hbm=j��ä�\���Ti��VmºT�����D�6UH�qd�Nq�c�nq�kh2:Ȑ�¢�1�4+�	C��L����E1J�ݨ�õ���/G�n�lqʛ�T 	�>�ς�oʈ�M`��	��6:c�mR�=��j�Wg3D?�e{]�k|�#�jUҞ?#�}8�<0��v�%���ϔW`��0	�^깿�:�#8���z?�Զ\[�Q����w�~�����3u�5z��NV����Nt�!�O��e��ţ��\�[��k�u�g
���'�N����5��yw"5x�|��3޶�/�V(��e�[dn[|��Vg�cޮ��#�y�1;���u{�e��&f#��Q���-<ѻQ6��%t�W#�3/k�g��E��Ӫ�u����E���Nm �F�(�Ǯ�.E�{����k��/������g -�n��<Y9��	�w�-�(��dA���yɖL>>�F�9pt���&�;+��Œ{P���nM�Ot�;��kR6a�{c��5�W��F�?�
�KD�4?��h�U�����Tjﮰ�6f׫��/Ƚ��v����ݖ����X�A(eA��L�������:���\;ދJvJ�,?6����+��$H���
�8L2���-���po�o�1jX����Խ���7�u/D�9:b����n�P��<��U���m���r��K�Dpj�aC�-��G[ӈ���F���Mݱ{Rgf��;�yٝ�#��,�{�O�U���=0�VN����b�h�OcUW$�Ut�_�F'�:�[����*G���k�����l�PZ}�xN�qI��r�m]3��F5���6��<�f8C=&E�=7ϯG��.C��e�;�Pw�j�����F���2Qtr�o��!�1�u�z�޵QW�d�6�uy����^��W�t��Ru�5hܒ�����/x��2�^T"�b�Kb�v�[��E)�����OH���JXL}�2�A��7�/Pޛ[]�	�:����͖��kL�/u4>� .$L��ͣ����s49!Iㆄ��[�F����{�z`�=�,��-�R|&T�ȌyC��8��t�d�r=:,��=9X7���pZ@C���3jԾ.�ǭ�b
��m�=�7��.���HZѮٸ���8JY|Z�������`e��J\�m�X�C��m�e�	J�n���r��i�"q���>(��2vő�ˉ�.w�+'0$��d�A��SuKc=�][��+xm;�WNNuzZ)mi�6���LA�	�˚������.�l*[��en@F���2��Mv��h.'����>�ŧn��
�N�8ޘ����++E6�BE�R���GH� �xo��K$��o`� N�]x;��X�
�9��]٩F�7u�v+��w6v@4P�p8�os��Ћh����*y���[��f&�Y�'S�r�4�=(
��ET2�ٺ�"3z�CV��Od�D�:k���3��͐ǻ��&l�V�`;�{��w[8�ӎ���fd����7e��i_]����tz���U7���	��6��6���n�:�Rl׻�۴�
8�)��RTC7����j��;c�}�İ$ojX��B֚����_�H��d����9h<�ۧ�uHa����h��Y�K�ð;�Ua�u�10�zc����x��*Ҋ��f<�ggyu��+:�փn��g빍62L���i�bU��tŋ�֠��Rv[�����*%�,�0���>5>���=2��^V�Y���X|]��&���P���\�<�s{`1��A���͎��fM�x
R��R��#�@��d�g
-�qS��kۗAZ��z������M��Y1d��t��h�����#�$��(bd�R�}���!� AO���dB�R^:�ɉwO �nS���X��ϻ"ي��q=�Q�Q�̥��f�Z�-M�5�B���=b���g��_^���ݫ�"k^��:dN�eIl��Yǲ��5ۼ�ȱ��A��oi>�m"�]|i��tS)��WOu�I�F=�de2��nP��A8�4;�ɭ8�Lo)�؜c�"�N��MA���<kAaJ���CNL35�{����76��A�EV���>�)Q@Q�2�j�媩R�J����Q�(�D`�KB���
	Z��2�Yl�pb��F"����Y��(,�U*�dŶQXV��ԹLm�A-��U�P�Pf1�+�Z�.31��S2�F1f51�+h"�`TPKeV�&��X���K�1�&\2bo3M�dD�8���is,(��˙m��D�r��rej�����k,Ȏ[1�m��q(�ڥ�KK
��m��X10B�b#�)�2���m�efW0��X��QL��m+�Z�a�\��r�s+���LC��ę��+��c`*V��`��\��qˋ�Y+[2ذLl*V��ԣYDm�%��Յi��Um(�F�8�,L�-V�ɖ�-U�"#Ү8�������&X�33Q�Q�6�������։����UJ���-�2�U��mBq �6�cM�u+}��\I���r�Y�����f���A���N2 zG+���ݲĘ{wjc�|������Q����r���\��oF�>�Y�l���Rx���^uO31ێ�k��m��⫰�R��z@b3be�z��GEu�K�>�Q�k��t��3�)�"��5l������Y���x�Q�r9R�nx�k�����z�:�Ė�UJ�b(`prxT��+"���a�h�@ߗI���.�+{2�y�R��j0X4[<Oa�S�f�H�pxc3��hX���c�C4R'�J'��L�x,�B�g}=����'�n\>�t`"��ި_�K���R�m_v4��a���5�^W��)����&Z�j���J������fql{_V���w���G�M�mC7�H��j��q`�mՉjïL@\j(���5z)]��O�2��m9�Z\�7�r/NC�^��g�'ܢ�2ߟ����˫g��puKW
u��2����­��o\��9��6ON�U�qJ]3�!�j\���4tk�g��5ԗ�뎷tQ����NG�Apb��7��C&�tgo1����L��|�w#��W��b��s!�f�V�3�+���\��!�z�[�ǹ�sjǨ�&\PGʵ������M�*��C���W���b��٫�sck6[S��a�:N��_*&$�d�U�߱K�P�]Ŝ�ko��nn�n�3��Cj1�:hy��460�k�h�>�;ۋ2����׻}�w'��f�JX���YS"�ɺ˧k-�o2{��|dv�$ k�'h
�aV��U�Թt'��/6:�0�`��GK�3�� ��f��=��b'ke�$F{a�:���,J/:���m�q�8�vk����b��Z< ��,k���|����P�$W.y��d�os��O�t$���>�[�T���%(6�GT�x��8���tVq�Fv�9{��p;
�����	܃�\V+U+|�Z�#[�\�u�S7G������������0��@�G�VDc4�sʜ:ɳ�

����_��ؘ�j�{=t�K�����+3s2��a��t�n������+Sl/��_ku&�l��m��f.��W3a�U�q�7E��\����k��)N����.umI�vVΚz�QA�w˺�p�G���[n�kyS�:*�Z[��{��t�v��1�}P	��$^8��+j�5���w����(!՞k����J�F�[QϬ�.��tEM�0�c�a]��)7��qY0�f3=uLT���S����r���L?�<��κ�{�&g��x �C'u�"�?Y�5�"P�:ʁ�Pkj���(+�P\�i�0�^g�}
/F������?
a[w�L`�&�T�T�P"�K&��"�[ٸ�h��j�k*�x'c�T����nCv�A,P`i##K! �����R��c���kZz�%��aq����f9pbߞ�1�]��\���ީ�z{l]k�动ϴ0��'e�ND�<��5�p��>1m�B%�1�$+����z呷�s�in�UxT¨�#C�(u�%ٵҥ3��@<���8��f��S����|��*߈J�{:���t�p�>)	��Ì���Uq�� n$d��Kt�7�e�L��2�ZX��2��aܺ�Yp���7R�l;>^��V�~�ۺ�&'zjk�ZIu ����_@���1N�iH�W����vܝ0��5������iToo�r�3���� k7��H�5*�x��(a�a��r���ڼ\��<;���a�spu�Fq9R<5��5��r�Y^dS�/3.�t�m�uN�	����T\%Dhb���f�rG]�Cp�g�����]�v�����]6Rv9LNS��pA���'�r,<1���&�S/SK9��UdK�s��N�jpP�B.5H�<��5:�' !����ס�������NY��:ڿ_��>T�.gf,M0v}���]Ĉc+�5�dp^�T�W�K�k���<�6i��Wih�������vtdv��	F{_>h!�q��	�}L=WZ7���3��EY�5JFBuʁ�$kp&�^���Z�4�����T�;\�԰�J��Б#:�T@1����(wV�v�� @������eT1�f)xqA��N؊����'I��n(}� �8V:��mhH	�"5BTj�V�z�*����� ̣���gN�un3H��y6|_.��M�eN~͊��߯��Cf9;mt[k1�yS9Qr�	i��Ze�w&��&�6t���i@��n	����$�u��LW��>����A�d�C��B�zoъ@zc\���1Qy��M���WXpH
|v���tT��h��G����1YZ�|�,�i�E���Ƙ�[�RBΙ�円'(1�b�S����G5NQ��p��)�w`�ռ�p:/
Պ���e�o��΂�*��GF@��i��58�(�C]��#Ks���"�<�� �!�z'��7���܉�I�U�ږ0�񹷇ͧ7��{C6��7�yZ���!����Ju�1���xj��=��'+�૤.�V��r�Ma��2	CWIe�s5��v':cZ�}����%�)",B2K¶������B�#�+zu]��c����]�%�ywX4s�Q=�������c.r�^-3r#u���׷�7�8��L����{q):�لl�,vY�C�Or�fz7�1�+8�^�zͮ�d�w����J��/)�J�s�̻ͰK�ؼ��lg�ȁǻZ�|хZ��Y׋oq�{F0M�R�a��[�|׻��
:�r�\�F��&J|�x�.�m��ډ�l	N�̯;�u�u�񑗓#�I+8
8}�.�e
I=����R��N;�Uҁ���
�2!��7�U<u_R8�w��טn>�}��G���/��L1�q��L��yL�{�6�r/K�>j���{fq�;x�9�@s���CJ��U�	����9l��z����,�TR�[�\�ؠ��pŒ����8�������ʫ��8�k��=R�NO,�.��Φ�]�8���h=ؗ�>YС>���,-�vj���Rf�q�X�p!��O$�s'�.�B~S��Cn�pΌt���ACj
��zM$[���������g���s6���m!t���c�¨�Yu"��H�+F+j��jeR�vK�m�aa�U��݊Q5�'��=�^�ˡ���l�]
p�}��\��O&V K3��`�yj>�x�z�]#G+ʼ곞�Qj�9Z4F�V����,�f�8��v&nm��<9S�G�NA��/ �ã0����k,,�Xb�NV�%�KmM�}cp�,�-<�:���u��i�o��hl*�
ۉ�r����νܬ!�2��w&� Y�;priG1b�Y^���j������&c���.�ɏ-T��)ʵr��r�dNl��Z6�U�$.d���9G������8t}���wg-�w��]�����eI���b7�II��x�옮rU�ɍ������������t�E�� �N��]*P.�}DU��:�[Vfy���Gve�����*=�_Tb7'=f-��Dך�e��^���#:�{;��v�$���"O�J�V�eVeD���:�xq3
凧<��)d�%�{˻��[+f/
�xX��*�q�y]|������g���ۼ�v�o���h�2p��V*Y���.��U�4sǨO��������v��̧ƚ��X��Vlu�	*a�^���{��H���@��&�b�m�sux�~�5��wil�6�N=��D���0�����E�B$p�{�rZX�>�a��5m�V��޴�J��r���UX��@l�(��p^p�F�.VW8F�e���/{��|��K�=:� ��3tF�f͊������+������2q���v�\yCc[q���pξ鏱(�E�%^��|�;Q��-��2�FVQش]c��$���+ŭFu���2D��\o
�tGueB�T�ť0��=���צD(	�}�''�E'|#���8C�������*"T�c :��lZd���%�d�5�����<ZF8P��&cϚ��n��9�w8д���Q�ps�L!B�*P�� ,��i�đ�n�S��i��wG8t6J���g��%�g
ك��a�d-�����,�Y��tOc��3٬�j��{�=�|�B�~k��9�`�q=R��`�H�_%D,�#f}�����y}���<�rR�	9B����Fv:�Y�3kKLVk��V�����A騎`��"�����,!*"}� d��Gd��Ls�G"�Ҽz��8{��.�a�T�4�˃�F�ي�OT��Y�siD�q_�]3�Z/n\e5��d;[7U^��g6�MCG�w�u���C���9�r/q�Ȥ�A[������s���S))���kt�����^")�14�;�<U�0M��<��tVF���_uuZ�H�-��yh�����Y��?�I�軷\#��3����`��a-B�r�2���}/=��;U�=�ծC+o�@;:2�욹c�=I{�2ҕ~�ꌪ�wJ�V9��RԱ��+����9[�z�<No3���s:T���Gƣ�y�~ڨb���-R��>��HC�*������oyY�8N���4�(�=�̑4��n+�-�R�aL-�}X��'���õ�hd�M�&���EE���"a��'3Z��QT�~k���l��7H�}�_us819ps�q����ɑo��b6f\�*��/0�#��(8n끸(.����:$2�F8Q�۾�]��ZZ��e���VT�>���Q�R��K�i6 �j����u�9IÎI�/e�"[Z 9�C�����ѯ�C�HƷĨ�R�f e����l��Wl��d��M�-'k7u����{�b}�l�3�ϡ�ԕ ����Qpa��4�/2�������
95l���떏w�v:���+���' �Kw�T*�{{��`���<X65�١Ⱑ1�3���R���ox�ҧo�WB�Vz`%hږ���61�tW��s|H<k�U�!y0�����ĩ���Xx�ꥮ�'�������v���S�3�]%��-�i:mM�R�~�n�̌u��E�yڵR���,�� �2ݭ�L���E9��=7��i<�;n�m��#l���M��1�/5��<y�Ŭ�q�˪��;@�eɋΞ%�,�#/�h�p�V���ZB3{�xd��2N��Q9P��68:�R�j�^�����r��eYB5�Y�a�{��y��}���� Zj�.��^KA��e��I���P�1)��sw��l�9c
��8VG�o�0:��2��J2r/��g��ǷW�]�o9@��6���P]��s��a��ct�5�R<�M3����ʯڗfQ]3^���s�����|�'Oa߃8�����w/���7�A�b����J�	�=V�V5Q,i�T�4�u4�s��ڐ^�ں �YOx+��;��J�`�{9���y���k�e�[y�F��]B��� /�na�P���-���iҰ{L*�oQ�d�c����F�/y�o6��u����݅el�
d��n�d��i���t������o�X�Uy|�n[zm�wN;��Ѻ껻{��fʅŅ+ùn��0FC1IMn�U�]�u%a2�PSu�,>�޶Z��ۑ���m��+}�H�d�.�3SU�$ⳓ�ݷ�L��s>g���3�"�U�ʂ[�H�@�N0�'�f�ԎP%�U�X3�yw�o5ƹ�5((-�]���ܸ��樝;(^��°b�:������q츙uj���-e�-����Frﯴ$Y��M�/�Ğ
wY9Zf��C.��]t�F���X�S��.�cV�=��J��KJ���1C0W|��.�mNc
��p)F��ݠ��<U�՚�0�ua>]#�>����������#.ͺ��X�\\�X�K�0����s�Iɸ���-:��v�ֵ����맱��ոI�:���cF�vdHr�(X�h{��_>��t;�v-�C�K/C���Hit�-��%��G���]�
�Weqy�.<��n^�G,X�SkcpV�1om��a�*�2�:�oh1�&u���pՀ��=�q.S��ۧ��ɻ+#��+w]�>��i��Z���E$����Nڐ�S'�ټ1�Dh�M˾4�OEZ�L	�od�7�/9�ռP-�ց[��V�ͺt����g[��#�E̬�Qt��r���0���}�&Q�gmh�9�ɒ�Ov���Yd�&������j=��>��=�nVfH��|	��0-������M\�B;���,�癛��`�!�����v^���N�\yn'%
䢹77�����Z�����d�}z��͗ה����p�΃J�x�������v���/O"2 -<�ͣW��*W��R�[��f曢�Ό'+0��� l�ݜ�ΧA�{�yYx�y��"V��{��>���.���Y�+(%�W�n�3m=�������Źtњ��a�"lM��f&�J��yE�/�d,��%Mb��2T�8X�9:��h0�;8���Ьb�|>/���h
��*���s
3-A�1j�PQb�ն�1AX�[Z�UVQ���i(*�6�h6�(��W,�P\s**3"��q�����q������G��TE�5��Uƶ�J+-"�p�0��*�c�V�մR�*e�*����Yp��e
�l�r�pTD������2�4�J�ȃZ*mTX�jc(�"8¥����[L�����hX��9KJ���5�V�s�������9����[��5�V��R���TC)fe���K��R��c*"��11*ۃr�䡉��s1�-�Ys&ZQ�2�E�\K�\��pb��L1
�QfZ"J�奠�VT��.5H��)�fZW���e2�W3r�eq��1�U��\�-�1c�UJ�D�.cE�0��EDQ�T�	s�=�{q{�����SY�sP��.'��=C��B�Ѐ�t��LN�O�S3&���q%&Elǝ�tn����΍��W'\�8t��}V<�h
�����:y��RW�q0ʗf�����T���pwGZyP�$39�}ٶ��{�/��#�H�8�7�oZ�[2\<�q����<�y��M����쎥r�;T*����8�ǪL�rU���(;��0v��=F%��s7��26��]�!r�ـ�80& �01�R��X�l����43m��Oծ���]K�2Y�T���0
ugA�H�0)�5����xj�������{3�	~���_�	b))#*!<��"�Y����zV:w�"^��)w}���~riB,F�]:P�����-�9Yޘ�W�<*��e]�M
���=^�8��NQ�1h����,�{�9�@f���G�o����ɹ����B���+���+LX�Wj�=��*��#j9���]���*:��Ł�ZZ�8�:w�6씱HM�ʻ3�N�w`�*:���U����ԽJ�ˑ����n�uq��wy9�pd���b���<��v`*
��!mC�#0̰����F�s��zj����Uf���*�Q��p1�::��P�T�e�fg@ު�R���^�,O0�)��E
(}�9b/��P�:ʁq�ו�y��]�^7�h�5��xn!�L<4ʞ��w�.H���@��cG+�[]���Y�ȗ�<�_��GL`�Y=L^(�3r�* �C��h�VxQ�:T�G;۽�$ ��K���'
�aiQoj9�6�ť�DrUHR�|�WO{j����� X,*�'�&J�xP瓞�5�p��>1m�-5���\
)�\�]u���Q-K����H��k���+�}*'՝�q��|vx���+���{kh��S	��Dc�*��<�1��S���i�N`>�ks�!�M�P�8P8s^FL���l�+5ƀ�[jnz4�V��]���m߹���է(�P���k�ȗ�-ukf~�+b��Ya�;8�y��-(w�%��'v�Hu�ڟ2����V$F��n`J���@i�w�š� ��(�x�+L|��a�1	%�rxd;O�4�qb���ƨ�2VI���:�������1�zw�"�)���|�Q��ɟ{=ϩ��YB}Q�Rcǖj��W'9��}�u�5V���d�]ܪiU6���=>�x�5�Tl�t���Iܤx��ff�p��t}���l��+1A��/%3^:��c�K�j�k�7�7N��B�E���@3S\�f��՜�'�iM��ѮT�,C�%���]�*���*�眐W�y7���fRG�5L5a�Uy�٧��O-4wJ�)��3��k|�_.����[S&��,��S羿%�<����W�"���(h�b�N�k4<��mڪ#�rTtueTr�u*1^�1b��A��0t��Ѐ�����A�w!V���;x)�80h�z,�+fa��-�W���g�ܝ�8Bx�]�t��M���|�B�C���?��޿.��b�y�q��,�\��Vk`�nXai���c	P5�#��:�K:���j��\7���=:�^| �.� �.Ϯ^	S���R�kZ�(j���I5;�ڲnj���rr�jV*�L%�V�ua��^�t�r���\%��&ᗫ���_6"z2���L��/${�h��w�������qc;Z��ʶM�p���
�y{Y2��819Am����7�C���3������y�T�`��:�c4�(���p7�9YP@�N�;NA�1�GZ��gi[�$����!����c�8p��Y:��c���?-�t�{Qnf��R"G7�ޤ	RD�1��Y���&��(gOXjU�E�e;���vɘ���oPF�v��ǺT|���(x��t�-�x�)�Q��g�ݞۢ�[�dȽ\z`%+R������|l���3v\�Ᾰ���i@�ؐGe��.����IS����v�G�0hH���ёb7W^����M�R��\�OCTF�g�Qw��U>�& 8l�+�;.���*���{b��C���R�F�)d�'����͍u�d\nI�M��ٌ�g
�Ls=�$���V��z{Ъ�\��^rD��b3�����V���P˒���j9��]�����v��K��ud��=�ǣޗ��x�An\\��h�ܾ�+;m�I�A��P��R+@ٙ1l�%*�4����Z:�"����u!Y)w]J7׺$�ƻ��:2J����	0f"�\��WnV���8>�yL�+
ȼ*.W��IYiv�ӫ�1���51th��S<*vX��:9������\e���ͧ}��E�ml��z�c:W_�&�GT�T�P*$�ɾ>�:�z������x'������.�P�t��L�V���++(L�йi�Oq�Y�S��cS]�����)ܡ�XCy:�r�1n��}V"��gzf,c�����>쟐J��/��i�-���j�T��=\t��p� ���pF��*�_b֚���+¬j���}��5��(�فWm�����P�,_��*I�=��x����'�7d"1�o�A��-ܫ�}��W�{�<gOxX��%�Ң�^�X���*�����:�J�ǆ����0����ɩ�j�K�I^�!�F@#����cT�BB�I��A�5�+Mx��0)��f[�uS��:��Ke�P8�μ��$��7I�Z���wM��s��aj$3e��z�J���i�vh�ԫ�˾-�H�Q���u	��52�<���f�tiQ�����LM}R�
 ���|�<)�"-��A��{�z)H�O)����SƑYFフu�'�! �����J�0�4�ȉ�NlQ�*p���Cn���ʮ"X,+>ÛP�:r�Y��Rz��4;J����=�Y&S���f��L]���ć<�+���Ba�d�	��q37�e��Zܶ�#
;jzcc�s��(��)�(�v뽓#�!�"���3��<.u��]�R��
ھc�8a�SӺ��QC�@��d�F����r��FS��E��P�T�R<:�Xx[R�ph1�����c�����ӊڷ7�nf{�92��z��&��*��P�0p���/K�ݰ���#�[��vW9��M�8hC���a{+�=5��z���,�T�Rc���c���(����i2�rJ� �4c�'�Q"bK�w+Luf�-�T��YW���#O�u��:6nOqTtfB'hF�=+]%�m:e��c%b��q��r�a�"�gpN��ت*��+6=�����ф����$��e� �Gt�ⰧL�'�|O��ʐ��+G�N�1�͆V!�/+<wr����+ps�pռ���N5㺸�ӱ�& �r��񨞬P�%3��;�:~��Br�n� �1Tt!�|���H�z��i��d���Q��(L"�u��0֮ζM�h���h�_n��`��<sٺ�n�k���yW��6B:jc���o����!�r8m�m�S�i(3օ?u����ã���t�L8v����UPX�,fK��*sH�i�LM��-I
�����t�R��/ꇁ%i�>�(`�ǚ~mBWy�=���<�{���Eu��e�q9H��BFٱ�R���ȗ�{S�R�z����}}�;X��&��ܡ^��z�bF��S<���W:������㨐�e6[:7�oLVĩ�r6i��硧�5m�Z��
Li��~�
�eF=��,��>{��P��Oi�k��_p(>���ʇ���r��F�Jh��%�T�O��O}�e(�T�:l� ��έ�Ss'������l��?7b�|+i��o�N��!ZŌԣ%�/F֥m��#��2m�S���ﬧ��r��T�����D�L�/��{�e�������;���Q��1b�.�;�4�X5��]�%����hѠ;�üU�T1\��j���\�;o|��2U�}���؜�S\eN��0*�7�;J6>�\�&����;y��u�N���JO�8Qy��R�d�/��&!7v��0����ɨ=>�|Pw�:Ĭ�wrO9�{��hO�psr�L&ai��D�븾816���ʜ�2��׍߶�s�sV�˖6�x*��
�,T7u��!�T󓦉�3��"��#�d�]��y�.����ʞ{��Eh���ƍf�=u�Մ!Y�;;��.�,�w��&R�$�L��)�#1�t����|j�˃���Йi��;�̽�rԳ�*sH�b�=	O�x�k�|B��B����^���q�5v[��f�q���!Z ���dT�ڒ
��v��S����G@��mu�{��W�F�fѶh�ñ�@��r�� �� Rl��(UٗS��I]�!ca��r3E��ǜm���J��dsr�Zt	W��o����y���kj��m�혣�gq6�y{+����~�;Q����'!�G�<4~U�l�oT?��oYqy0'��IC��)2Z�3�sssd�%��!+{<���j)*>bdMlūt�G"��O+͹���8ȿF�%8/w';�A��Tp.�B���J�ˢO�"<��!����Ր�;��ǋn�g��ܞ�l�h(`�00ƀ͆ߧ܆<��>��Pl��2R�_�p*�A�C��ݲX����24��ZԱxS�3�x:���t@�ל��"h�\�%0�NC0�Ԯ�W��lp #��@�(2J�wS���mf�f�{}�.tm)ZP���M�O�7S��bt�4TL/y��ǉ���zs��v��\8*:�8�RNj`ܫ��6�Ǜtj�7i�ʄ{n�o_6�)�0�Uzu�%qy�j��A%umT�U]=��������0sk���Y��R�:�ٻ�8�`�ݰy����:��{ �z8fD��:��+�*:�*Ģ�Z{���&���4�+if&��"1�iv��vm^�h�\WҎ�I-��c&����V��U�"��Cȍ�k�����O��~�k~��a���O��'�j�2`���s������8\��:7J�z$���}p��v��M���)���»����Nf i�� �":����݄e�Stu�Kq�:�Gq"�Hj��Z�T�[N�ᵂ!�ݴW����;��Of=�c¸=4K���&�\+��;ѱ�,���[�O�������+;�T`��u�H� �7J�!{Ϭ�L�!c�/3]�<�\�.1I�AX��x����6"��
�D�58�"@ˉ�ݻ���#����:�+�'��D�AxU�𿕦,X�ʉ:U{γ�=�y
9���[�EX�;�z��l_�����L�k����]W�l1�E���W�ٛs�n��¶���8a�[=	�hQC���hyYU��}����!����ޢ�v�����/id�����el�e��(f�޳��rėh��]�w���
��n���U8��Q'�lj�N�U�Kp�7�}}�V�l�l
��Ui��>!�w91����W|�Eu��lc@Nf=:��n�a���h�GU��ݡ�:����dglb��ɗ%�����-ܕإ+h�;��F�o0a�0e��,��3a���lV��S���]q�$�*RN���٧_�{;p ��A���*Ɍy	��G=�\3����X�y��M@���L�ն���=-��5����us&�*�7��Zan����g��:P�꽋�>z��s6�e*N��2й[����;R ��U��]���٦�j�3dM8v�xn��Uz�]�؏i �iTZ�ٯj�㗜�Qٝ��.4֡oE�)sU�_p�t�L:1�8��ryze�1��LF����$Ҷ��f�E7�Wd�t��XC"6�Y)G��Eգsndbey�x3x(*���o\���3���.�m|���f��F��9>�%Q����uZ����k�[�
''|1T �\�����7w�f�����YITi̡o���ՄA��! �ǎ<�{z�0�¹h�̝��d�Jͬ�S�(�9���w��d��#��f�v��� |l�{W`�0�&	��mT�%&tR��x,��(�$�T�yv4�`���,���jZ�L�p�-��y�xk�:���@,K��ڦ+���xq�`Q!ws�ڮ�;�M�B\�P�ym�\xvD�7wt4�R0ᤐ�G���w��μPξj�y{�(�f�άiYv�`�+An-Γ��S��#�ϣt'A��I��'��G8-X����?!s��^����֮���5Ma��zL���ʔ�Ӏ3��a砘�������V	TIǣ{��7mdٖ�8�T�D�������,p`�n�si�p���J&;��0�ٛ�]˲���w0��N|�vN��/iau!��r��W�)V<b޳7^�� ���k�޲먙&�Ӯ(����,m��N����:�c��{�dk�XЇg��1#*��ט��&�>��:�iYv�w/�K��uѳ����Ӵ-���u
}�ɹ�� �#,��Ը4p��֎�,j�5$��VL�o^]?�J�����r��w9khCq7#�U5!�P�b�I%�Mq�&��-��Yh�X��gl-�'K��.�g �S��ث�b[ec�r�-�%��*��Q�YZ�����0i��T*%i��2�KZfJ�2�FaB�Q�\�-ƪ���e�J�Q��\(�*�,W-�*�dV[D�
��%r�J&P��X��2!U�6�*
��؉��}u�V��ƹ�ƪ���4�V�5�(���j�ƺs4�
��q,f*�.4b(��(�f�QqmKi�K9��5h�FR�ڊ���	Yb��V�*��f+R���r�Ŷ��f`Զ�*�j�V(ۉUUq�!��c�Im1
%�1Ub�iW,RTd����*,SL�ʈ�b�,U��TQ�E5��V1��QH��i�X�J��%J��b�#���Ei��"((�X�T��1�:�R �$UbAE(�H,+Z��!��4˦�DAk�kE�N�TT��Me�QATrت� �����k`���,2 ���ن���5��W��g\j��u�ڳ�q��fn�Ր�sMꨩ�(�@�q��.:�&+���ք����ɞ���JjXbB�{s=�X�&�%�n�+z8��Ժ}˞T�F�c��牱̮ʨu��£���(,_7H2bBK,s��fV�����;�C��L !2�EzyWxXYyP�׭��s)1�VQ�.5�����}�׀\;[v��,l`��z_s�HS�+�e{`�o��2�¦��\fM]��6ض�!��1[�s�s"��u�%{X�uC]�����'���.�>�U�dj� ,��w<&0G���fک�X����aᡋ�xha��#<z�qʲLW!(���2a8�v!(���<�"WE9�������,g�ÃapZ�R�Gr��򢬝�\�ܗ�ލ�qD7���\����4����Th_j��2�yt�ސAM��I䚲��y`�{�9۔\c���*RW���*.U(ZJh@�˗���iڊ������ތwu$W�=٨��t�<'3ٌG��_ >É߷U�.%M@�)w��QdS��o,����r����|��-VʸUM��n�FS���O6g\Iᕆk��E��3Z$q�m��^]�~Vb��F��C�ߦ�<:�@ê�
g]�V��빽���Z�g��<|Mp�/�%)�͟�C�U�.gYڹ�ŻL<����WS��_Z��H��;^�ѳT�N̴���N���Hʪs'���ש�����e�ڀ�Պ�y��|�)��_��yۿ'X4m�܆����Փ�8'o(�'B�#��Ҁ���9_���s*!.�;�4Kͩ�f�'��5qJ�o���O�lUx�>g�Cf�"�j���
�S����Z�l͟^=V�R��
���sB.3�����F��>]O7�6](�2o�Co]X�z��:�r��{�����Y_�A��(��ۭ������=Vln����S��*|�2����H��w= ���s��*�̐{��=ĲP�T���A��(TR�*��l�VT�9:|�}�\⦒y^�6�A���ʽ�u�i �t~bp8��+��Ou�q��L��",�nJe����:��Fc��0댴�;��ՉLڵ���m���Z�C��Z�4�~���]ħu�|�M�.�[���ctR*h`�b�md��O��~ä�O]@�4�:yN�횥�ê���t�2��sW�o��0ڻ<=�|O��˃�LtX�0X�u�j��pF�q���I�=����,����C����*�׫5>�(쏣rK?C�c�5F2N )�h����K�Y늼<��}�`�J_kJ�Zg���f
��ym��\�]뒧X|NٕH���ݹά�s�68;7F�j`"��T�ꇶ���{���(���ժ��L\��R'�.z�
��� ό�P�D��!Ӂ�'���F��!��X��&v��h�8��(��WθJ�
�vL����=T��6���)f3����7����8z���L��������F���`��{җ��V�t}���^=��]IC�ͪ��Ls/N<�L5�x2&�FF��y-�/
p����{�Դ&E��v����-�݅)U��w9��6̰/�:$�Aα�z�����g::*�����uѼu�3�ɹ���iEuJ�n�n��XA�4xB��{��{Xx�R��~��S�͍9Uכ��������CsT�3mD��!���2$��.T����m���st"]��l���<���
�Q/6r�73�bcK��N9ښ�9k9�L�d8L3����"�"���W'\�P�
�<�[�pTK�&��>���z�����;�s8
Q��Pn�\�Ez]�k�{U'm1��G�S~��Rx�����yJ�h�5�v��k}jQ5׶ju���D�y�5X�v^,�..�7�0�Jbx�n�DcJ�:Q��m\��(;�YA��3��Ù��x�:a�R�u���W���)��H��O��G�#�x`c�nQ�]�
^�|U���a��� �I��3aU�+�9RLt��V���q���:�I��JPDN����3��28w�$H��]�����+{����'f��WOб�1��'��;1�U;:�5��졯zr���;�Y�^�gQ�0�A:F;)`���GCI�uZ��5��5����M�̝�/�i�ܬ��A���qީ�2�D�3��;=���NUڌ�Y�Kǽ�!�N���� ^���	�;\v�c%��j͖/�|w��7h!��~u��[.�X�zx�wR& �{|���+O=7�e�b�7T�ybP�e�ɡQ�m�(&86o$��խu͍'����7=�ýT�Ւ�ʴ3ʭ���6,o,k�&yQ+V�7.���챴�P��h�@�'��)o�КF�>���hy^������yI�t#~�c�|C��u�oԏ��mS �c+�ۙ��b��ٽ��<�4ĝ��ɋ�OY�VL��4vt�X�X���bFŌ�ź{v�et��RB"� p)�\O*�n����v�U�[N
LMB�M�#�:К�ԁ�ظ�������  ���'�Y"`��7�(s���r]����gRjU�'��bۘZm蘕�R82u[�9�9�[�B��.wr_��ԯ3w7Zw�+�e���pQL��]֓q�WJ��Bz۰�d��M)Z�H�ORy�`�5S"�n�K�^��Y	��3��
�[Sc�����ٞwX�uN�)�F�H���yZ�-vh���k�gU�^Ҕ�>Rr6�o���V\Kk �I.��Y��ݩr-ðE:�Pc����40�8P<P�� .�U�b��J'���sH�Sk/9���*�nz?H�[Z�KÃ�>�
��e*� �؛��1�a�҇�ރ	A��|\Ԭ�Q�����_�p��(��L\��цkvekoٺ�g��b}䨌�F�xX�8�5�r�3���X�sڗ&�+�����[)m]p����y<��3\��
.�r�!��6(<���w����W!�@�U<��S��p!�mD�(��M�=1��d�*u��Ǥ�ԫR/T�!<��1[6>���d�Y����_M�fZT곑��[�c`t���	/�hq&F1�ft�9��6:��{���u�X47Qw5�Ư�'1�gQ�X�G�:���f9oR��P�K��5p�8�&��ya���x�l�7hC�ᡳVy�0��ڄ�%���٪��):S���m��̋�$�b�t׎dtI��'���ȑj��ۋ�{s� t�T���n�@�R%�3X��L�P�6�8�Vu:u:􆾽N3��#��hna�#�)lد)W.�yU��
/uV���;�툢�u�a6!ّ�Tt}	�_i��\��U��o\W���7����P�����7p��ǨTdp\T�^Ўޤ�r���ܱٓt��\���g��<��]�&ݳ�){����|�\�5�:�@b$Ys��A��(J,g���o�r���	Ԅl��uBb����혍 ��{	-�4���x��ۢ�*�Ã��Ykc�K�/�hIT��u��(PpJRx��CjL!Q<�Ez�����'�2�Q^��=-�Hjﾊ���(FᨗqQ\�C���f��5�١�P��&kݹ�����Qt8�}��Γ"�u�P��8`�<*%��H3��	ݼy����N$b�V�u��J[�Y;ުZ�{����7'Ոb�<�h����H��8���7F�L	��Rǩ�Rd�TFּ�S�p��].��a�mn���GJ\f]�ٽ+!LP}���}vݠ�
Qb���huzV�
��2s�����me���M=�;�]�V�qٝcz:�؄Rj�.�g_���Nv��S�FMvh;����׺gq"�A�qr�|Lܳ/w׺��c�����MU��YpT�8<��P�W��Z6����F�U�<����#��Ӈ�(���ve��z�fc�rb�J$]p�h�k��D�c݊ŏ{���q�yV����Cj�
�����d������n�.|;3!�J�p�s/K��k�� Ɋ���%�𨝖#7gYq.bLe�uKt�<oB�򥎸(B�CsT�0ƕ��8�y�7��|;�(̞���'�(-�LZ�uD\�u����B-Aw���S0��'r�-j�NN�{����. (#X��E�[}��r{���&�M�|ogM�p�zmW�������,�}��Vq{�Gm���������<�C�z=	��fW/��Hm`�n��$WY.��7՞扵�ls�:6��U��xLF��4oS�W���Y�1K�41�<l�����E���w^����:3����ud�V���ed�����"�X���{�lHdΗ��N��t�뾬�L�7�}ѐ�^S&%ll�bs"�c[�\O��{���7�E��	����=�Iށ�Ot�ܨ�N��;�]����Y���?5rSp���`�j�48����Nr�T�ڷt�R �$l����!���g�E��3����q�M��AUAʘ6� �:�t�{nR��ɂ��z�L�4�WR�6�;����P�����j�a�����f�ۦ�F�.�ݹô:5
�
�\����\�K�4����M)m�jI[��j���*�ڨt_5�����iOls۽�v�:յ���޴�S��&��zv�^hwy�:m�]Ϛ98�c:�*Ә�׽��&��.�e]�t�\���R3�5�̎<�O�bk{��ם^�v��߇-�d��y&6 �^�����	�{,�wb�i !��v3 �*�Ё��U�Ց��hN֫�+M��yi���3�wu�M�lgl�L�vc�J������Nq��d����1ۛ�{��U��T��GGL�Ǘ
���[��|�+�����qo4��a�.��|;$,�:�s������f[t�T�N9�T���·����g� 1��d����n�D��ԕWe�a���}��A/h�m9;E7F�gZ�y�����K� +8���9^ߊ1������Ǫr����C�rX��u)�eק4�z�9�>,|h<�ɿ7����+ŷ=;IX�;�0�`*��{qL;�v���c��ԭsrf�J�qt��p�kB*懷�{�YPz�����M�\�!����ө�xn�X逺�ڒ���=�x����{�$ե�lJ�ǕI}3�N���X��g�?Y�����V��j���A� 	9i�� @���d�p 	p��^ß��t3+�%3����ц�3�Jz�i���g�E� H^P��
O��:�SC�{�$�4K������  �'�:l�}I���?����?�'������x���)e��X*�S�Zѕ'jN�/a���Ѱ��Sμ5�� �t���w�����!C�?y  O��$ $	�X�2 ���~m(� ��	%�I�Ng���?��$��:P 	��������*:&y�D~��&!ْ����'@5R󐛰�C{�&	ᐺ��f�.�>A��I���X �t톽��h�9;����|� H@�J�������0.g��S���?�tp�� �?�M�C>t�Zd`F��tt��2�N��`��G��ہ.A��_#��hI��P $zeXjX.H�~Ծ�����MT�b]�p�mֈ�J� �C��.K�>��}�C�  �-BѓW�`�����h��t��8'�w""��H���@ $	�W�̑?���$�O��5����4�=:�!?#�?����@���Պ��ɂ�������$$@�d�����Y��a���܉�U�b�܁���$�p3[���ֽ����R �>0?����|���  ����!��!H3ax������,2Gu��'���[&ϼd�Pgn����G`#��ߕ�Q���@ H������HO��xl @��O��%����K5Zz���.b�Ohq�R�LC��D����C	����� ����8����=����@����:� 	���-�|q=��9��_``#�s3!��������@?� n� � 	�L%���9т ɹ��k�x� �O�'�����ð�;��i;���蓯2��u�?)'��?�P�!�����]��BB���