BZh91AY&SY��UJ�i߀`q���#� ?���bD�|   || ���T>��j�Df ���BAYj����Y�T���lV�@b �T �2͒�HR�4jڊ��M�n�Ul��V�Ҷ��Ւ�6����R���F�J����S3VՒ�)���P*�lȓa��5[2%mF��M�V2ئ�Z)��5�w�{KQ1d�#j�m+iU���m�3��K&��ٳkll�2M��H56��J��Mm�+YjYi���ekZkZ�j�
�M�I��U(�4�m�  n��u����i��X�m��N��U���+V���B�]]tpà6���ժ��F�5�غ:�V����޴��a�mJ���l�Z�(��  ��RU�Vw�N{��̽��8y����2�m��x���R�^w�����QPyYĽ�"R���z[hK�Kܩ���4�y�nW���f�o<�1Z�5��ִ2�����Jֶ�[i�o�  ��έ�w]��Ϊ>���2U���������[���c�|����}΄��>9��^��*W�+���"�Y���J�K��>�ﾾ�[1J����J:���+���^��S���6cU�Zֲֶ������/�  sχ[m��wz�icm���r��{;�v�r�ǒ�i*�O����l4}�y���I����vm5RP����ǯ��*��}\�))�n�O}�_Jl�i�>�iUm��0�5�%RщS|   ;��U!EU[���z�[�������֞��{���z�d��f���C�ݫ���=�u��U�۽J��))��9�J��{�����5�W�;��Q{��/���kL�����d�jm|  ןU�d��מV�WMU^w�ꦴT��{�w���*j�n�R���y�.9�{��l�۽��lʶ�"w�=z���ǻʽX�[jx=a�=���Z�����f�j6f��٩J�P�   Z���WL�R[���ڒ�Oz����*�ֶu-��QN�n�lo=R��J�z�{m�+��ۭ�:Vڕ=vܸl�U*U��Uǣ��S�7�g=R{^w����Uj�ͥ�֭Cl��   8�QA��Κ4n����kG�y�ID�����b����ox�U��+�hm=�^�5�9�׽z��Z��]�E{�M*k)$�ڑT���k|   g^�V����*����^��zk���<��=���I��Th!�;@���=
=n�6��X���ު��=x���U+Ǽ�i�U���m��[f��g�  v=�RA��ڭ�w�����M��tjl�w��hw�:�������UR��ۊ Rݙު���QT>  4  ��̪R�#   �� ��M���@	��  L@�~JJUF�L &�	�0��	*� @Ѡ�����jm j��Om)��P  I��PiI�4�O@��h h���?b߯����rƿz�������ܳy�f���7rE������CHj6�Le� ����{�0lm���l}�m����7���m�lm�Q�����=���|��C� clm��2�l�o��p�v66�����G��o�Lp��hv��4!�84&484(�hq�!�;mmm	��B"�hCh@q�!�&�ƇcBdv���l�hv484;�6�c# �C���Ѐ�&��B���hv И�Cq���0B�B` ��`��c���@�"c	���� �� � �0B`0C��v�&0&�dq����C����l86�l1��0C��!`!�����m	��Blm�66Лhq�v��� ��B"�B C� B�BcmmƇcC��2&ChLhphq�&4;b�4;b�"�cBcBm��@v�m	��1c�����;�g����y���]-;eT �C\1�t�/����sf�d��)��Ж���r-)���������P�r�H�E��Ŧ�;*{�\���ᰥ;�=�P�YE*<&�'�/��n+|�Rv$(�'>���ض3�i �����j4,�X��^v0�k�h��&��A�r���q��kۍn5�4�݋&� nn2Awp�'{�P�ͽ���`��a��:�#O)
������i�GvճRw�|$ߞ��un����R�7w"r1˾��x����}G�$?<-����:�	�8�@��=�Af�6Sњ�1e@d�`�/�@���n#��F�2�V���-W@�k�A!{��焌�]z��T��#�N��Ld�Jyo�x��Ln�^bT���v�s	ƻ@�>�Z�+�:�0��=`�m"䜱�d����ϟm_pǒQ��u���^�7�}w�P�w�[�m���h�n���x���p4J;�=ݝv�n�Y���5���p�,hd;!�5*�Y�5��X��n��%`{��Q�e��c��oV+/E+���0b�uV���f�eG�Ee���d�9����n͵MPc͘nVt��ƞ<���yT"�Yww��0v�d[��Vh���n	��Aͪ�H�i9f�VGs��i�SWO
.u�� ^�O�B�a�F	E��
���A��S`w���)\ka���f�<�]W��i���<�գx��a]����q�jú���,.�]��qǪ�t� p/h��&OSV��7�����>zX<��h U�]^:�,�[o8īR��Ӷ��V�hc�̍�*q���`9Cty������Ӣ��r����6k���T��A�Y��ݹ�&w:���9�p!;:�pf��z�L�#���6���$s��9o\���=��g|k��	����s�c;-"��y���<3�N�B���?���f���Р�ݶ@'v�>J�V�� Jw�FF����z;����C��Q�8�Ff*�nR�W�-&w�׶��-V���f�! ��0�w� ��!�̰�>�+���\<X�;y��v���^�/d�#�wIŃB���B5�+"s���!*�7Z�l:�XP����܃��~Cx刬����ӛ1��#�X�S�j�z;C'GA�{!=�q���OK�/ά���� �s�z�:cڭ���<�)+�[�`�ik��e��-]����E8�ؚ����r�` �Wzow[���+3D��afb�Y�kj3�h�n���j��,�񱢎5r�ndN�,e^I6(�s��f�T��	nX9ųHZ�u]|V�ɀdɭ��Χ���}/��j�o
0�qͩF��Y��jG˻v���b�42޳��f޺���]�_e�*�C�ƹ%�J}���u:8tRu�d松F��v�Kn
g6�����{A��x�;��f����m��9u�z�X��>�g}5�8gL�r��y��u����n�Q|����al�����';9�op�F��HnΏ�r���ߓ��u�w��̤�1��ݝ�l�v�Y��w���=�ev���H�*}�o.��5�Ԕ���cǎq]��U�q-�Sv=�.ܺ��w�ݹǁd�lv�f��YA�h;y�;pMcjcx���D�ۍ<V2+|�=��t_�:ɋ-�ӱ��{{5 3���5h��o655��E+��Ӷl��ę��wO�X���۳h �˭<��Gx�>MX>�=�A�D�\�y7N�Ŕ��XJÊJ8u��������" {!�2���Z �eG\SNWl�Âȍ
����^�u�v���ު�x�Lؐ�o�ߑ�{sl��562[6�!ƭ>@=�B�ó�]	�	��>60)��oK�4؇9�r�e-�ɷymx���N�#�ŭ�U��h��Br
ZǗocx����Pv�#�h��Ry��q=��җ'0J�ǳ�!�mQ�f��� �WL�Ռn��_�xk��hw
�6����D�+�*�S��ע� �d4�y�U��lo�*,�E/s�/J0���Љ���(��8�j�u��s\��ap���1��<�g���l����K8o,c��;�w$I�9-�����h�/�;��|gS��T�9pٛ5 �Kz0�&�֝�Fh�ܑ��4����պܭ%IY+������y- ޥ70�̢^�;�Ԭ�+3p:	�GP���I���˯ ���U^/rY-U�`�:������'ڌ6�;�Zyi�˂�.�ܳ�u3Ni4Q�	��0�0���D��#p)"���!���0���86��Y�CGt䋙%r�GJ��,*���wpY�
ZqT��S��`�����0AB�#�y���v�
�c��m<�(j�\m7����wݽ��PI�4r���g���ۧ�N�$�P�x�7�҅���F�~Mdk5`��D�(6۪M���J�^z��Q ;�ߠ�j�l9�RÈ���z�9Y�U�[����[t�li�?��o��6N{�n�7-(���2MԻ�����^�q'��A��d�O����6�,�AY`�ż�.���0m�Ɇ�¾$C9��\�|����Jc�Qkw2Z���zwC��$�1Wut�<F'���E��m���#���������l�Ԍ��t�*W�ҷm�vL0=w���I�ݽ8�Ѫ�z�:�F�׸5�u�ң_i<{�"*��.�u���=;Q����V�{�'P�:w�u�z9N�n����\Τ��h����.9�0΅nn@�M�;]�5�!dq<Vj�]��n�sKj.nv��D�6wf��}D�]���6��tͮ¦HK3S�������5��H���cC��vMvEۻ[{N��Q�X(2�#�&S����nvt�@�����B`�γ�W[����b�ivh}�{�ROV�A�\[�[�u/�c�l���	� �Q����^v�O�^wl��ئE�`�tݯ]�w�:��4ly�윐ͻG+uJ����Med;��cU��� X�4Ex��-cK��&em����:��`zC�y�[�M��.�x�5���x(��L��n�`wɅ�j��[g{C�oC�0�;��[�K�HT]�DÝ�l�SE8-��<�2����F�1b,{r�K��]�w�� �Lt����hCwnS���,f������9ǝ iO��wN�0$��z75�5�r�V�e��	�S�0���M�����B8Ex�\��~�XK�;��/N�e��mt4Gô��8]���qa:��<�(n�&��Xr��D��`ںw�b"S�J!jI��C+M�Mf��S˱��R�<��N����c\a���'�c�h9���t� 7i�]|�:a�4��;Jz>��
��{��HD�
V<cv�֖��]��Dj�e[�I�7X�+x��2-h툩+�Ѱ+V]ړ���U��/��9�|Ҧ�f�7Y��Ș5M9/Cyi2r��ڟLt���Z�H;�Syv��l�˚ePy�v�&CsZ�n~�x�!֊Gz�����N��t���\U|�W@�����Ge4�`v�A������2��poT�z3��*�nYV�:��8�wkX`k�9K��Q#iq��!��9�ߏ`s�-��M��hn7a��(LI��4��Y�f�N�`ӥ�'uT�A�Jv$���$�yJ���\��0��䣻wD�JwͿH��e'�#E������6��O|n��u.����R6�
wNM}&C��u�� �n:ʝ{b�v���	{@���^�.W���<���Y����Nr�r3�=�n�J+xf�Y�-���*�v����^.�ه�L�j']�,,{�j�ĉNU���[x̬�[��gQ*�c��"܈j[�]��w�2���ͻ;xȴ^��e��	Ӧ��ڒ�&:7S.(�`Sؐ�4�6�y�n�D'�0?�&/�M7N��5a�ȲSgH�u�̺�
���͸��u�H��a�����Lo�o�7�G �'�8��
r�R�0Ey��K��aOt��X���rUwn�)�b���3,����&�t�Mh�m*CA�-v�u�v�b�6���X�)=.i��,"�R��"��t��s%:�.J��@O�������tkq��PpiG	L�P�{��ǆ�ʌ�V�-8 ;o��H�����6����w����H`Z�q�0h|�8���=����qp��Q9c��b;/d��4t��3涷�"�롕%������&-�G��Z�
9�z�4�QϺu�?
[|s�kd#���o5B�-BH鼕3�x��ˊ��]�8h7I����S�iK�ޙ6�ׂڊ��q/���q�qpٻgL�]6�oH���:Is]W38��I@sZ������@���sI���M,��2}p� ���*�F���#�Q�\Ed�������s{A�)���u�t���ȃ�{��	t�Z7���������L�E�9����0���[B�-V���7:�F�T��Y����w�@�uW�3Z3*�u��&��2���4ؙFKY-���㔳���޶m��b��㺇5�f��J��6dZSD.�<����p`���[��v$.��KN-�e�;��p�vGa��+�g>�hCWv24���zH�p��8�mn�Â�w��3s\�{��	9ni&�hho�W����zr�`d��p�R����N��]�np�㧎4�X��5&�ydY��]Z�E�_�r���,+[¤�lw�X�Y�9��V^䓈�"��9��!�*��G�X���Q	f6^�q�O_�)(�BX!��q8>W��eچ�ܮ>C�p�ٽ{y�]��7�:"��;D�Jgz\�9��Ec�ۉW5�q�뉘4L�U���7�fX��p_��sf\1���a��w;��9�o�a��^�*�����`}r�_㬓���ۼڡ�:ڼ�a7�6�{��U[�L��-(P��\s��e�X��UXw((cTi �\[C��=�Lp�'f���Y��F�bCE�n�.�v��j�v��	ۤ-9�L��
9�e���7O;�a��9�.�e�k��\���� ������6P
���:�=�TvY]�Lar��{����v�xͽ��ͨ���6E��v��2�ܟ&ˆ�ڷ�(cN�;sw�(��ϓWg�.���Z�fbT�p�}��:1ӛ���Acu�7P��#w��܊�ф<o�=�#{Ӎ^.��n��tnh��JD�4r����\Ft�ͱ=#��u�"�+��&I>y�4�Q�f����)0_lۦ�������빩�Of5embvudl-w�����"�-U��Ph�̋3m��Ъ�M]��u�N�^�1:^�1�\��2}@l�ԅ��O�J�4�B�����K�<�k3M�9�[l������H�ݱj�%j�֬u:����ᆤ�u�c�Z@���|`����;3��D80L��7t� B��sAh{�M����G4Sg5=�nc�^��M�ZP�Z5���:�X˭T��#hF�Į�#�[C�Fh|����\#XyÜy�J5Gy Y�XY�X�AUk9��u|G�:D��5�Ϙy{��8�&���Q����X�cY��'­_����]Ũ�@�,70����f����ot)��P�
�˺x5umC�gn�+tCt�X���zU�&��t�v���F�l���咁�t�>�.V�'.��N��܌Au�[�k�V�^Wf-̸dp>I:�7�2u��*�Wc&�u1K���G,!Љ2�#x^�'j������Y��\pa���&
7AJi��K��x��V��P���*-$-ksn�`3Nm=�'(��?�nϧB{�:��fG��Q� ֿ�qHD�9)����:@.HM	GW|���R�C�P��D�k���]ߵr��Ӡy�*���������G>G���h%]OE���
«9��wk���g՚s]&Mg�-�"�D�7������/�=�����sB��USMl�e�k�,��7BˆG��3 B7NQ����sV�C���׃&mݿm�
ѿmMBX�B,��Y�4�')�scr͏F��ƃ%f4���Wu�a��Z䳨�hn].��x�{�L����M%S�Z�MQJ����w՗kM��@/iR�T�"�9��V3d�s�K(=٨f��"㲙e��pT�l����k���޻�dfYf�ŏV���l�&���ܽ2��0n3ۗ,X��Y7�3ݦ�)S�!���ǣ�Vr	���#Z�O��`8���i��vwT��a�:�k�w�^3y��u�b���@\ �,�v�Ա�OT�'u���S���7�_��Jq����)E�y�y�bi�t����ٴ�Y����{��:1��1��z�I�����[|�Yw����(�pa6O0V�хX|�n�
��` ���� u^�́E,d��ZpmU�P��[��a��J����8��Ѻ�����2�V�4k%�rLN���w��U���e�+0n9
�et�����H/1q���U��_"��{��L'N����^��5L��e�����_k�yZӔն6���1˕s��M���ncv�5Lٻ4��d6���eK��ѥ�7��+��
�
w� ���_t���L�F) d^��.=������o�RԎ��,�ޫ�Z����a���Ǩ��ĉ�o��[fڋ4�[6���8��V8�9/s	�qV�t�nŭ��`�f,�6�I2�he"�u��ļ�;�P��8��h~{��	��{�D�?}?��w���9vx�QÜ�f�����U��K���x3�1��� ���|
�iռ6��f�S��:�yݤ��|��&5ٶ�.�_fƯ!ԲF>A�����*������*o^�����D
����@�׶�ny]��.�e8�I|閄�����;��o2���T<���81��i[���4���v�4�W'�8�(E�tes���*�;׀�����Je�"%�ט"��q���2c8�V3���
�#�A�i��L;�9�+h�b{�=}�]����(Y��->w�fv�gQx�T!���R�D��4zs�2�rylmI�Us�˘HN�	ftw9�v�w�on���X��hn�1�I�k5�7b; W����_�۳��o�M+���یؽ�qW�ax��$m�yul���-�5^AW4�7�7����ݮD;<��]94��:�J�XM	d֞`�O�b�`���TpH�y�KBC�(������Nӌ���ܴ�,1��2��������]?c��H��n�V�U��c�Wۉ'�9{�f����ؓ��+�x�7�<ՠx!tD;�j��l�t��=�XI��6�QwQnl&�V�w��*�^����yo1������e�+�-�g<Sh9������l��35�nE@Z�Zf%�9�kH�l�pW�F%�#+k��v�]��
�o-���mN%Y�Y�E�]s�Fm���,"�$Y�܆���IfЌ�O!�T�� IZ�{����������mQ�-�UwM�v���")������;ʹ�d�)�Q�h�F���݉W���n�M,������G�/��컔�����e4�{}�����[� +�rz��S��O�X��J��º�]��0zt��g<�<�»G7Bee��6z��ּ�)�磆���͙��䁬�af��Y��;m�q
�̄�s�Bge�L7�B)�����cu�f� �F_f�u�������?����Y�nG��d���pw����_���wd=P)zާD���G�J�[���R��I��ҕC}R� �U��Sj����3����s�/��I��iX4q�:ýLS���ny��K�+�����Szf-��#9BS{R�j�YL��V��!G�.'�q`�� Ս�b��9ǺU�ɛ�>�nM~/�d�����2�����N!�f�{�~�N���,pcF����B�˛'q\J(k+����v�_����r�2 �=�-~��Ae;ވ��s�[t{hއY�m�o�,����,��i�4���꧂���'������g�O�3�SlK����۴��>�@QL�b�}n�3e]1|�K:`��#Y�5#�}��LG3�#�i����G ��#"c�F,���G��h�V��̋~>��=}�L
�>܏�o�D��݆�����\�7���s�P)��pMQ�F�	}��k�B�
��u|��TZ�sZ�.�S���\`3�-�٨�ymL��s��zwC��X�+t7\���ׁz�\Į!��=�/=���Co��vA��<�H;�Y�Z��)[EFݾY�Q`0�r�:�<�Ѯ��H��,��W.��s����d��gK���ċ(bGK�nsh����"�t�|�����g��C��H��םy�\�yj̨�b���RI�bz�;|���G�Gۑ2�A��A�<�Ⳏ��C��\+JU��c�����+�Z+k��+��Z�U5̬�B��ë��|[��*'�q�^0:����䷝$���M]���;�*7]��m<N��Ի�p��ێ��h�� ����Ǘ�,�9�9�9C��6�f�+�P�Y�}eNzv�''�f/y�f	��¶��!�0qrǻ�\��92�T��2��ř��0���-с��ԙ�kΗ���͝�A� -�V}�a���b���T8t];r+�L�j�{˸+"�Q�u���g����XG@����=іbQ�>���˖�/=O�J��	ۗ��Tv.�l��*S�	�8�rԶ�]����6���T��z�=�I��#�e7/��'���g�C#f����	z4�y[����Yi��C+d7�}�;�%����	�k����zd�t�g�W�Y��:o}F 3ݳ�vCi�(�^�2� ��8���]J�R7Dز�9��ݿ�5�������|��M��Ws꼁�YCAKu/ɪ��qvEa2���23([Ƃ�2�GU�ˇʾ~�d�Ф��
�p���by�[Ņ�����<��L��1�a�{�����Fh��1��$�}*��E���F�;���|���h۵��;���7mA}�L��aEm��t՜�e�U���k���T���Si�7�[<�7k��FI�,읣��y�v�n�I�J����}u�w��w���^������,�ړR�˻��Z��E~���A����m�JK�����v\�U��t�`X�/���9�l���A�pG�d4�]��sX�s++/�Iȍ�R���}Z�[�8t��ej�M^no���`�Q�E�D�n,���_V�̓�Dw�3%��r��µn^x��es�$�|�.op�`O/hM9�q]⮈n���Bj֦��{��9�]�ri�T�Mc�FGn+��&�4k���kػ'x�����މ����tn��(�^Q���3�뾃�X�#���r���ǯ"]V6�t�Y��cAH+��Wf�t�|l�(�gV*����eH�3q��\N����qגp$�
�U"}�uI,��K���T:��qge�����F�V�ǽ����Y��v8�q]�w�����Zy�6�����[2��p� ���u!.�l\�ͺ[�c�G,Gn���v�{�O&Rسm��b1�}p�ig]D�K<����-`p�`[ָ��{��-�U�ψ��M��f�l�r
dE���n	S��=� 8���b��QSnl�;�4�3@��=Q��o���C7�ͪ����u���@]h���hS��	z�'����~![J۬[ܰ��r�֙�j����AT���y}�^����Mn���f��m��N�/�:�7f �n\��<E.��}�ӓ/�[m��7&E��;uD���Y[sL�}!L��G\>?� w�N4t��C�Һ�k�[{�����y2rr�=����z�s%՜����'u�r
-��T�ej�sS�b�:���7��8q�%���)S�G�;�y�'e;Z�u���+�G�����Z���UҲ^��:f��aFYd���:7��^g\����:��sGC@�E��t[)�O��ߕr��P����qC�dv��r����v�ŠOu����c˔jN�N��*,ե��E��	��
�%>ȣQI�����i�$�;���n� �OQ���_�Q�/-e������8�z��U�� �ݒ�m�̋�p���U�kM��$����&o����Z�^�Q[�g7`b�R�!��=�E�_�\pܙ�.)\�ˮɪ�J�o�0��䞘[�Ԑ�~&����ESU�d�*j�'R�����j&���{YW�1�.����⡩RU�� Ի8��M��"��F����c���4y���vԜ���+�C5�q����Q�w@���g9oUY���B�|�q�ǧ=wco��K��l&.��L��r�1�5���sy��������w�N����q��Z�؅��~o�ݽ^z�+��Ww�%�V��zKp���l\���M�{V^<���J���,�ߣ�=�=�Y%��������N{�d�5W�)�R��פ��U���. �<>K��OK|4��A�:���{��G�ݓW�&,�=���G{�d�^�ǻh�&������VB~�.&X}�+Ar��q���%Z��^=nL
J��"�����o��g!g��Lf�`s�)�d�C1�4�����ն&�h�Q�p�w4s	s&�:�p�3��P�6�����{�My�:A��#�>t�wp�z@�a�1����n� U�6�(K[�v���c.��w��N�blk?{;�UyϷ���靌ѽ���kmXn�ĩ�f	˖p���V�Y���jC�)�]?��꼼��.ޞ������6u�
JL�w�
�0b#����.�%XAV����ވ�۝;�!��Y;�Q!�u~���;mM:-�Ǹ��؋�ٵW]����Y̹�t�C~fe��31�y����a"���3�n�:y�{��q��&V-źs�-���L��Y������;�ç1��}�V�^d��@Tp�V� ���H�Z�����Y��v��Mc̉��w[x4��X4�V>+@�'2ӽ�˃_n��2y*C�Ց�ڶyǥ��-ዕE�W����[��������	�/��z�C�l���h��{2�1
P}H�0�׽��u�S+t����:dn$&^~9��L����ȗ��l�,�����S�n*�z�!���y����&�~�.!N����g�QV��5ow`�<�B2����~����az��(��0m����:5l���}�q�,,�Ԁ#ǔ�Fr�g�IM�Ll`�O�u8�����[�P,���"���"�zI�'Y����\a��м��:Q�=�����d��e�)sW75K{p�=ؖ��μn'�o��T��U�
���w��;e�<�"�'�z���<�,[�B�g;��><�Mg� �-��_�)�`�&xeї<8�W��m�;���Z�a�Ĥgv+�Hd����I�68H)��1�۽٧r������9�o��A��(�<
#c�V9�H���W�j��)��E� �칿{+Y��\�kgl��N��Y�{������[1��`ƨ�����]�k6������V�̨���M���1�T+{�konL0>��&�{
�y?c�>!����xL3O�{���PQm��;m}�9M���eɒ-u�.��^c
#�S)o�N�[�s��`�-]k��e>�nJ�.�D0W:�I)QK��-暈Q4�ك2�C���	�2�LM���(��dc�]��i� ��<}v<+��}��y�����Z�U8A�`�3��ޗ0 �T��pʻ�ݓ�,�b���%sR�4Γ�c���7D�N$�x6�Si'X�*u�-B�Y�A�T%wA���!w��0%NS�����ˤs��AK�`�跍:��k7P3��еۂ;���59<���Xe�ow�I��K�*s�� :��G��L��]i��_]:�j:��}xh�^������ݝr7�`
d�F]f&�[7J���a��ؘ�9�>p���"Ϋç���<�Rv���n�λ��V�=O��`G�;�u2����ۑL��
��������"^���0���趠U�B��.by�f9YjlO��	�y��oeV#Ӱ,�̢�3�ܸ�):�{'��N�ѕ3Ҝu��6�:���
�nŖ�ѭ&ad7���*YK]��G&�{����]F����,���@�)�4�7]���'��Xq��x��:�Eu�N�:��,䥃5˙����:�g���|���$ve�I�ՙ�
z��O�kH����u��iՉ#�&��̵�%��Q�������Z�Ż��f?=����^=�����wuk�,o6}>k�:�%h�b�]x$�M`l�� �rh�v4��;<4���!� S�v}�W{NӇ��}��	���q�����(�:��6����ɝ6r����t"缼0�;tv�R��2��͙LI�J�n��)���gt�c%�(ir�9�jƵ6��&p6�wSb:���l���
�6�s��V�	�[��<�x�n��l��dQjp�um�����qgw�����V�bI57�p4v���%16�3�8��r����A��t��=�ɧ7����ya<]͖�u7���Mo^k�������\g�^���C�০lpy5ڤ}��=���H�ۗ��W!��������d����m�/�ׇ��Q��Rȿ<�c�S~����B*��7tһU�F�uH_�tP�T�������+;,�4�D�	�X�a&���R���ڏsd���AK�5����SQ��%�"���x�PY�o6�uԛ�kBc��TY���Nae��]�_p���v^�>�_�eǹ	�Z[F"�L���I�,eUJ��N'J����:�l�=�]��Zd-;n-yIv����_�m�F��-h�۴����!{�!��޵��ׄ`�z�������@}xU,n�U��,�ёB�R��j7�,���%ǝ>�:��yv�;2�HK;Ԭ]���j�x�C�Y�@����k�w-�Ʈ�gA S�5?f��뫖�d��F�)כG�3߻�,�)	"�t���2��b��qh��L�$y���6�ǵt/B=����-�w/�\����xQ�{O�����������)Tݔy��JQy�w�P�HD�	o��\�Zy|/�'�	8K1.���!G��l�hw�/b�u�D:nG��(��pk7���JJ��S�$7{��ٝ��]y23��Ǭ��c�����w�Q��3M
;��i�s�*vŇ�b#{�I)�(X�nC�n]e˻i^�q��Fؒ^,����'6��b�G� {�}出vN�����̾���^m����=#a���9��lݾ%YnN���IM�4��YŮ�=C����2.	�.a:7�b312�Gf�Q,4�W��!2r�6�� ���s���MH�I%.��d-��\��y�Ů��䳲�u��^�˵�w���7�77���S`�-u:tuy�T�W<�ts���tfPwk�UXpj��v�.S6�r���$&��4��#?8�!ʡThCr:��]�e�lZf��F3A�qf"����j�"~̪���5qK)�)I���X� dd#��M r�]�8ʆT'��)����,��������������l �|��O����C����=�������_����vo޿��0j{�p�)��{}[�xf�%�~��䫆_),L�d�zp.�h%J�\w��m�6�Z<k�C-W#y|\��h��*��ܩ��+)�<H�@eϚ��D��,��@��}�.��3�c�����-C<K=��F��gt~��_�=�I��N��,��~�w���4�poc��o�3�˺��*ߗ.�]�O!������������$�bɕ�+ A
���ugY��'�S<�E�q�Z4v����h;1We�Ӻg]�W"�,�7z
B��n�v�3��w����}�/&H��8N|5w̋��~�����-X��~�_��G,���v[/�]�o5l\����3�N,Z���-��߻�Oo����y=ꢸ�|��c���YMt>��*I�]i��؅���c���h�<X4��\4��z�uq�T;%��-lՄڮ�� pޙO�d�,�a�:�EYc�SY1)7Zn���;!�ם��%q�~�."ZK���юg�52nn�-��S*Rźͽ9ܮ^HF�⥹�vJ�\��1���`7�띸r�	ɣr$f\|�U���c]٫�]�Q�`VL+9w8�b�e^��<�GDf���}�^���o������QfC�j,\¬�=��I�&�k�{5c������V��U6l�[H&ѧP1���4pc�8AÇ(p�Ã �8p�Ç8p��8p����Ç8X�Ã �Wt�(�����A���v(�22p:����oj���9pŻGw^WH��^4dY��-�^�{�dӪ�k�·�sb�h���0���(�a�����K�u�:�'���\�S&R���Ws��hu�ƅj�KyR�ظ��{!s䫜	_��l�d`ڕ���W؃��BN5G4�3Qg���*c*��P�!���V^����E�	-��2S���9X���������y�'���}�ل{_�ξ[��ۭ+�_}�4��|~�xܨ���(��\�ݲ�ą�C^cb����'s�#^iۮ��;Wf�N��tFɮyd��n���msN��Jjkk���[I
����C���y5�ĩ��W��_	=���aԛ�vo�	+]19@�ó�"�C�z��Ie{��z�I�ˑ�v�>�3��/�J�y�s@D��zIs )��%wsޢcc��o�x�]2o�����Ƭ�n�۾�k�T����Ɖ�Iq����Io_eԦ�ά�/�S�ǔ=n�ԭQ�˺�����N��ͦ�n����p�"�2����m|m�k^^TQ̄�.�~�ab�#��"M�h����k4�l\������@�0)r:yL��P����&�����lM�f	ݓ}�*M/�涷��]ux���jbޡp��=7<����s���Y}�7�x���n�����j�����4pᣀ�Ç8p�À�Ça��Ç8p�Á8p�Ç8p#�8p�)ԩ]$���[YKz�^�7GJ��;��;����0�؟\��٪�,SB)ŧ�t��t�[5�\F�R�̎{]p��n�t,�$~�M��wZ��Ui|�^�K�o���`$�����ln�J\���S��fj�ʭgo�����h�M�n�{��N��P�xLg�e>���w�Fk�X�p��O#�]~}k;�r5�_���k)��F�Ǣ�=�t�ԝ�|iaR���z�� U��T��H&Վ��d��q��ɓ�.�A8�nk�6$�Қ�;f�ݸ�Eu�M��Ӂ�ݰR�)���/�C<p��)^�-�6���{��E�8�漨t=��z{ݜ1��9�D{�-�b�O���H�\�12�Zd4鄞f�j���7�i���c�������k��o�$�tn�������yH;]��ۡ��m��to�0�>�M�2k �S�O��G�5���{�e��Or.��ʙ�8k:ks�Ŋ��O�hpl��^J�P=��X��g��؏�)#\^���=jy�x���ؚ>Q�Y��_��y��im�y4��|�%���4�k�1k�ΗgI�i��]�h��J��6�[�v����vX�@�p}3������^ۃ¸��ޓ*�U1����bNOg�}:�n��L���cݐ���sX)�G������/=n��'�qҸ�a�)X�&9��u����:���>94v�s ��RZVF�+��c���)=c�e��c�y��W��T��N@XةMY�:*x֌`��H�;��Ɨ�L��K��7=8�����,�ؔ*~�W�:6c����E��	8�fD5=f�*�ߢ���w/o���{m �7R��������]�������&�<L��z	"�-\ް8g⳨��u��ߛ}�Պ�͢�>��%�ͫq
�[�*�����X�՛�B��ok�p�"Nm��f�K�	ۯKѢݘ�u��I0��n(�[�D�6��,�AY����N��4�p[�B��l�s?�֛�so������J����P^j�CWR�;3b
�W!��V�6�,�4oo[���5�Q��?i#����8_wU&n���×�Nr���0�h��\�F��M��"�=Ӕl�Aݽ�u��Ӳ\�-��>�1�˷{��ev4VJ��!�)��'�&Ⱦ�ÛRK=�:&�UT��۹��
Z�edwsZE���� �y��ն��{I.��컠
6�=��+G=��k�^9�y�Q�c��Z�ʚFj{!Ԧ�̻έ�6[���v�dK'LׅY�P�rva]���h^H���
�޷�kl�,��3l����v�Ѳn̷�P�/Bc�j�޺Z	��{�zc7����C{��0���q�>����hYj��a�%W��Wke�%zi�f{n�Z㇇�(�����|)D�73�xA�j�r�ww�k�37$�������z�fqrJZ����x:}L�B��j4�?�	���r] ����яn�������ɳ-
<vK��B�t�:w1�n�;��<��Ȃm�X�X��m���|�#4��d������M�\s�	�]kYsn�( Yn�.��M����,��r�"�2m�R�#S�ePН���")w5��ԃPLŹG�/��~�x�F��(Ag;<3��	�؍��}xs�������:��K��;envι�ށ�xZ3�M��>�����H�����x�NRV_!��9Z�m�-�(��2\�	�7���8TQ��}�H:��8��:1`ыV$�;���4+���S��;0֯��AȮ���zsG����Q�E�%&��C�e.�ާ�O����٬ltv�f�ae��_7ݘ��_q������?�D�u%�i�{�|����f��ٲ�҄Ǫ��~������vk��'g�2��&ڝ|)/�۞������|���\]�(|h��Ѻ ��nNu6���_<F,�ą��A��6fӃ6 ���wF�B�0��y�\S�����QS�?8f�ZW4dqٷgz��`�-jnE��;2��t"��hֹ$ln{@��;�&�(����+���wsY�|����zWD~�yw�*k��f�9]�{������Ơ�e�0�ԩ2��0�W4qt����4�{\V+8�7uE��j����Ԗv����|Q�ex�f}� i>W_�|u���K5;,��U3g\�ݗ�ws�n������
��m�IY;ڪz�l�����1�-��z_F��;��A�xMo� �{Qg�/k��?n-!�Fq=uXOG)�e�)��3 ɉ��Q�b��2������n-�"[x�m�n��u�/2��f���=�w�'N_s:1��M����V���-���ΛCS� �}�+�1g����ssiT)�;sE���m�y�{�I�՚8P��c��[�8٭f��\�4ђ���.��hk�Z����Ux=��q6���3���%�ҵS�G�W��|�S+���;��g6��P}۬sU���Ƃ-�1K�{)�6uj9{ǹ��8t�=��ڑg%�^3��L�H��2�͵=����>2h����e���뷣��w6a��y�p �2b���l� �/����Fnu����i�������.�t�zc�ň�ۦ��O&�f����G<�"�$ y9;�v��V�y*���hÞ�m�gf�0R�L�+is�KMx�VG���Tb(���=@�g&�?�)ܝ���i��R�=�S��Ä�u{�*=}sw�\v���y�x�6.��9g@��o�ve]����`�z+Udӏ�<�k�۝=Uwc�&�Vx��I�+���wAYn������ʰ�v���n�����aU��oH�xJ}S��t�9J�n��ٵP74���(;W3zLѹ��+'�M���G^�!J��fd�+����!���qd��X�~��^�J�����[���C/���'[�b]JږV�����Z��1ob�tLEoH��"�K���=B����c��fx����)E&s;��c��\tp�ˑCe��S��O���F������@);]Hq�JD�bY�t�<�|^r�����,�n�_&궸"�3`vl#�=���_t�/����9ے�E�B��U��ze��
��&�����w6h�d��n���_1�x�E�o���̊�k{i�Bx$F�.}\����#c�loq�C��J�CJd����4�.�^Ͱ�2�Qjc����^]�S����ʔ��w�+c∃B/0�BY(p#k+OU\�W��G�[���=r�*%�݇��i�}r��˴�L, a�Kx\�n� �i����^1l��)Z��_�xQ��f9�ǵKk�)pt�[:Ύ#�7�Oix�ś|8�,��̗��wB+���&J�B�����kfL�L�q��b�W����C�wd������8�*�5�P;���7�K8�����n��C���J�=W.��o&�.cq�kS�cy����85ľ˦�(�%�(F�"��iv(��1����9ד��g�T��?{�/|�qVv#~�u��3�g���^:f�k���;�ds�̪����o���N,\����4Gp� 7��C��y�.e���Q�	�����m�D٠�+���W��06{�om�9� o��ƭ��U���N9����"0�vp��6�Iy�E_��gƣV�,��8��uC��/�B�*s�>�h0�fC��婮g0S��݉�zQ�2���EF�n��յ�����O�M��^���0�f����}[�7�By 7Nל����r�oR,îs�+V��"��9]�ѵ#r�ւ�+�ڻM����P�畖�M���5VE�j���r��g�~�	��z鐤��������yw/j��G#�Db8���N;-g(܋X��U�������voG�ep�l��1�	I��6#�����
eTh�ԋHg]�y?v��!�7��~�k܎�q��O|;��oiǪ;�$(AN,�:5�w��T#@��})�t���Vǝ��:��uܖ���޸���Y��9��X5�)a�$��{%맠��w�5�Yp�q���z��8�/�+C�}�+; gNR����� g�Q��{�ם} /gjs�`��2t�?b{���\nc٧v�h�t
����8$�f�${�,<�̻�b-�)$t��뽄Z�%�j�b�\с-���uXw{9�����~�RZ�ݰH�w��v��d�y�-�j{�L�y�/3[v�i�m��7|ڄ#��]�9�*���c�9�L����{ќ�%L����߮�ڐ����9�Hy\�!ͥ;[m( ��7k��9����r�d�v���@�=7��N��<�r�ڴ�"W(�,�[#ѪѴc�Oi���7��'�9���-a�� Õ�cu�ܸL��:�i"M�;vj�q{����^n�w$^bF�DLKC��	o^dYm���ٞ�/^���>�SUC��f��W������{�v����_����\�4t�������E�qK�ܯG^����@wΏTF��Ow:����;��c�l���n�>&�4%�`ߪ��~�s}�^���j��-3fMX񩓦�ӗ6�X���MUop�'��K�-Q՗T%d�7/zwRu��� � ��hcxo,�|ܳ�c_{ޝ��Ǉ���U{<����7��<;��K璻=:�GL���X?w�����,��<'z�s�Q��yD٭�<��:�6\�?7�oVpl��d\Fߟς����}�2Wi��vk�N�7��څ��\�2RH��β!��k("^V$�=�6.��|2��}*��	�&p�E�py
�{������W�gky�N��+�ɢRM^Ԕ- ������u���;���[>�@�]�eɁm��9�|[�W�R��S����u�g�\X�VC�M��P��T��{)���n��`��R�	�<�ƞ�N�w�m�au���&�Z@��pp[��*�d�К���..��iUx+ui]].�#����9ϒ�{Zn���a�[T���N���N��F�R# �R�[[�SH*�Q�0�4�t�b�.H�9 <��z^	���X׸I�@�3t,.}7R�\�\�z;1��7i�3��;��C�"�8���K�"/P�?o'��<��w�T�u���L.���4qt0K6ҟ��ݫ!��L���5��n":�4���4��&: Ֆ<s����]���rμ�ǏEuG�-2x�gӲ�#~�z3��P�|;�Oء#I���q���m�;�[@�Z�K�"�P��a]�^���v���2鍺��{��8����w���r�ί�p�0N]�N-P��NЄ7���i�*MI\����:8�Zc.�d�9wI����8}�O���σ�5^�O�yxh�H���w���/t�EV�/�m�~Ӈg-b��r#�z$�f�x��ʡr��wSw
��Ơ~:/-jr��;�D��פB�w�×��^��r�Ӕ-l�����ɪ��w�i�%�w����u���2^μW�����x{�������?_��?�����/�?o��?_��ǿ��l����~׍:cN^ddW��˙���^�Xc��ft;ٙV\���5��
��W���:�X�Dכ�r?xN�������=|m����/5c���.�+L'9����-zl(������C�E~7��p�ׇ�Yt/�eN*�j%\Ur����Z��6ڛX���5O�ʔ�X��q�\:z���j���gMs����=˅�E��Y�;��������*�p`#+69ۙޗ��� �w���6�@�z�w3��5n�6�t�7��|%�Ĥ�\�T�u���T]��yi����ů{_ݶ2�Z��D��.��.ǬR�\�)���["�a7�Y��e�F�96e�^)�9;,����b(�Ɋ��ZqXc\�-�5u�mK-��t��OGa��9�>��ӫ�X��z�oK��Ӿכ����b�]�*Ox<�AX��q��ef�18V�۝�)��TF{a�B�ʜ�,&sm��]O|�%�Z}������Te[;gy�/���U@�;̚�dΛ�{W4Xa�9{�Bw|N�s�&T؃���mOC���Za�-���'����T�Vh^�.��#�`y���4���v:-�sZ쭽<�\4,�P��wSƷnkq����؊^�Y-�hR���R�%Լ��9�bi���|0NS�D�N�Vo'ARQFɱ.���kd+ufV���yɤ��3��9�t��o�i�M-�\p�#	��܅�X���7�Z��粁�_�%�exer�������/]q �������G�=�Ȃ*��3;"��r��
i��mC"��L(����Pf=��g���U�)�K*�z��,�\�#�B��5iG���G�Ft�)�P��E�p���("���Pn�Us���+�F�q''u��"���",ȋ����&|8�Ur8Us2
U���y���Y�aS���xʩ�/S�EUTzє]u�/p/E��8S�ePT�ǜ�0�x��"�QQ/ ����r(*Qu9�9Fw]ܢ��ZUǝlx�(��E9ȭFU���I�2$�|���P��gǑr*�D��U�O)����Ը������U�ͷ�[�����F���������@�2D�f�t^37%2{��QT�	����/d{��ƯV��;����l����+�������{<���{C�7�ș��`���i1�Q?1p��f�{[�۞�<{�,�K�+�}���e�^ġ,3�0bxU�38�RH���V�w^{�_J�.�i�\��Ғ76�:Gl��f�{��7���S�gxQmYM��2���~Ku$�*�5�y{r���E�^�(��O��\�eJ��2̨Ey��w�n���6�sY��/D�/$_��l�דL�����kG�o���ުX]$�M�L����K��`��熶o����e��լ���g�(*��̠��~7Y�����E8��zf��d�kf����B�����\Y %䟅�k��]rV���V�ER��^�]Ʃ.Մi�7ԡn�%>屪���}�� xoP�坔���ٞ���+jL��Co"U��lw�A}�CVKర2���^�[����ܪ������(�/2�h �-���]b�\�wSRcц�b���=����eRP���c�*X=��-k���ˑt^5�w+%��q٭����(���Y���k�M����:�NN�pU����ߤ3��>��:�כ�?L�V�XU�M�k�򵕏��{�5z�5�#�2��^FL��V�j�V���,��]C%��#�-m�u�8���x
�O�{��B�X��C&�g�exsc��Y�w/�<��+���-V/�Y��V�<��P�t��h�z�d,��ԯ{��T*v�ݮ���y��]�^�Ԑ��AYE_.ȿ��i��fp�?_{w''��ԍ��[�������
�!�!��֣�]?OG���T�S��,�����6eX�P�K�4��qm�����/�ܺ����[՞�@{�Ѥ�3���� T��p���g�W���>�����e��ߺ��w!REm�	$Oӹ�.V!׼2y���G�i)�v�ng������m$d�y��kɳRt7ֿm>�{'��ξ��+�[�.f��s\}7�m*OU5�v3�q����%�d�s�C m�ک���a4�P|h�M' ۆ��wP�c��L�1��oz�.��>��x���@pr�Bb��H�n 0�ȕ�@��-���8��F6Y�6__��{�Y�n�=*��W+gV���F;�o�ŵ�`��kT��z��.�z�7N�1]��ׁ۬��V��,��n5My�^�7�����gX��8r˓Ce�m�^�n�yۧ7��x+�K� �����wCڻux=����1�N��s�]�9\��K�Ӧ=N]/N�i���ԉ��eh�a�P����p�az�io�,@�{O*޿�J�����ך������L���*w�ܭ�丅=h�P��Uִb��D��<6+��}~�B{5{Ӫ�߆>[P�F���TBE	Z�+��=m尡^]�6֞����C�����󙒛���S�w�%hj��3����$���9k�>���\0M�����I) �<�Scz؇�	��:J����埯z��ۙ`���$����}����w�z��q�J�*<bs��(��l��q)��A����Z�k��q���f5|��J��8���-��ڳT�=|edZ��C�,Fo��֯�rPޑ����L���� $׾���� 9pL	O��L�<"�@4���ཫ����\��=���)����ݗ3�xI�-�+T{�JW����ޡ��W����?E��l�7���&�������I';������IIp�֍%v�^ٔr2�yZ���6mE�E���s,o�B�P�������Q�H�������gr���c���UD����Z�%�����hAwz�S�m�Y�r�6����Əo�vUy	'+ՖTu�Ĥa��{�%p��+�W�3*D<��)��J��Z�T�-���>�f�����~��G�e��]t�;���}6�3b�������氧��D�竻\��� {�x��j���k���}�uuhV�J�.��C:/�f�N�Ls�Lkv{�|߲{VTݤ^�
R����&g�y��X6�u���צU�yQL�M�׳���OI���|��5s���`Q����+w{O�P����B������o���Od�>��쾺o|�)��:�
^����<;�����(2�zb�ӗy�AM���-�+���_�����7�ಜ�;R��X�$zvY����ޝL�%�%�/�1���ø�-�Зw��aR��o�t�TzNۂ�=>o�!f��:�fp�H���uk���e��
�2���QY[W{ۡ��t2d�*�u{wHkS��q��v�|+�z��ep��_0��~�W��&��>��䲒�J�Ee�IT��}��rc�W��]0��b;�z����M�=�����r���s7��%�D%�XI��md��#O�%��>�u��#;Gq J(�^�}�x� ��^��`fӧc2���Xr��=�ʩ�9���xQ�T����D
�mƠ��.+��v�|���Z��sp��B�7�=��~�Cƾ��RCs����5�GRE.I�#��4����b�jz7�w���UYLz�����M��o������]��;E��Gl��ڰ�^?~�{ޤ_U�*V�>�������"��5/}��ٕP������J̽Һ�,��a{g{�����kG��ýo?P5zP����G!�Lf�z�?��)W������y��q]ƹf��Hr�b[��<�X�\f�?ە��EEoLtV�R%��:��� �"�q��}GiE�OI��weF�}���L�i\хt]J�#yf��B���ƪmm)��}"{�&����ޥ���Ջ����xl�=����]�e][@�Y_����:w�j*��)'	�/��5[�x�;U�oٴ����6��EU^�̫���*�������/��"��z�Ȋ�(�K,wj�;�ng�,aw$<��z����o�6�1��6f>oT�*C���[ԗ���~�ʵ�Y�[yM�Mo{��M�x��T�԰��(b貼�+U���o�d��MXvl)��2O���{�9T��V�j�<���*�c�4��c{�b�X�wO�܈2}�k��{�rB�A
���E��P��u)�Ey���^����rV|{;V��Bl�VE]����^���U�Y�y���1{TG�x{�M�˺�ܣz�?g �W.1[傪M�&��d�ߵ��5�}��nnYu}�����DW��PY܂v��O�m�`�����Ð�~'N�@�y�z�w3P�P�Fa��˔Ĝ�i�i~�.-����H��ny�h�� :+��xn���2��;�3L[;=��5�du��v����p;�	^� ���yY���$�7� �prywy�۝'�������__t�����PrY�QȤ��h�[B>S7�ze����T囀�=�%֍$��̽0�1 P���I����p��w����Ƅ<q_Ј���X�\�I'sF\�#��O��lK�:͎��s[�՞��R5�w�y�Gy���^M���u�i��*=Gδ�ZJ�q(�t�5�u�}\�z�k�ڋ�'z��;��~�����4��o1qm뽛���O�x|�#���K3�3��^{�za�/��v{�A���Ƣkݣ7߷���j�g����z'L���Y?�M�ŧ�Ip{L{�Y[\uC݉��'���������d�[t���)�Jr�zu3MP5��ݶ�_M��}��g�&j�2��Lf=�F���U?�J��^�T^5��K��j� �~�i3A{�{�w ��r��	WZъ������#�Ix�&x��y#d�	ڱ��Tq>X}˟�"�g.ZUf߹���@!��x⹧g��]����]�-6Wu�}6Ҽ�+�zU��Ǩ�^q#
�y�C,�L��745Qm�I���6n�W��82ˢ󯴠�ĩ�*ӎe�;c���b� ���Rv�ߨx%Bkپ�wv���g*�CR	�]ʶS�s`���Hf֔�^��b��@�7kVm�O`ݜ��l��a"�����h�5:�f^�e_g�FW�B�������%ͭ�r��
��&"ʷ���\��=Z�Ѫru�>U]��P�bǽ�2{?I��nm�jz\롋�N�g��74/��J�.ȿ�NX˥�P��J��K�߈��S�k׳���ݢ�!o���A�ib�R�����m���j�yM�G��=m+v�~��\:�N!�{!��ԑ����\+	dny-�\��x>�2�'to���Vʻ���HT�{�·:k��X#�#kے�H��+h����q�����5}�pu���m���+�krұ��{��>J,������l��}����}���v��^{�Jl��g�j2nN��:	���}� /b�;�	����N,�q��=�Z]E}�wl����c��
��$�)� `���dv����[�6{�I^�t[)��D����_y��a���e���5�B-ZZ�l5�e
:��j@L�y�Wi�h
���X�v��"��/�w5����f��ޗH�"2����`/o~��p���d+*��ɜ(m��ܵn.�Y���=cL �*�*ڄQ��������^��xW�b4��x{�����7����Sٵ}�	h����Y�}��~�ީ*���F��~j8��<^�z�5S�L����ɵteމ�˾��e�h?3����
�{ƽ�7M����%v䬓-�Kٺ��v��� �t�˼
�1�=Q?!���M�����c�#�%�㝋�V%�B�$t���h�_�0uP@�]f%�|py`�����'*�IT�y-�_��Bo��$��~�p�'��z����Q��OoTE�]N����V��P���~�{�ŚcK��/�m9w�������𳦦���lG�꾭$����0��B��B���F�[F���ܕ��Ԯ7��dw{��?�S?GB[P�z6[Z��Ǌ�����l]\R��'}ΙZ;��H.��������͈���X2ZsF.�u�d��-�����p������]-'r��,G}N��Wp�cܼV�[iW1}�k�$�o�f2H��F���0�b>�^�:��*{���Hnp��[b5��IG/TA΋��A^o.��)Ťϳ/�����PR0�@�	^/�S�W1��'{��:�{֤ݳ��jY�ͫI+��&U�H��+���f��X��G����҇g�}����/�=4;-#��,��/l�uw���𹲽�{�K�����wH/ߝ���h�򛿻Ճ�i.�[�#o�p$o��wL���,�~)m��z�z���j�+��i����?w.�+uQ�3K}�˫�Ѕ����\e����411�@����"{l]�����e��[=!��^J�_�=����?�Q���hؠީT2����QIvꍗ�=��x��$T�����.�Jf����M����R¯L�o�k��d�y���:Qu����v{�J2TG�I�Ul9!������������`���;)�뼚>�l�K��n�a�xvȽc�o��o��\��Ɯ;�J ����օ��yb��wdWWb�����}v�L'�s�e^-u��������)@�U�Y���r�e�b��#��{�"{@st.�tr��t=Q/\��MaO�&�s(9,�jBn'�?(��Vr���I�ܮ�A��v��/-S�������Dv�Q��t�vؾa����Vql��+C��5�c
3��sY��Y�	�X���W4��li��M���}x1��c�0#�8�y��7l�{ҌY��F��l��V��a�/�S�U���Y��K���]Ը�I�̱�h�q�;Ք[�ϟ
��΂�<��Hp,H��/0a�4ꏦ/+=aq���)��$ϏVx��{�/Zȫ�ַr{�t��|��q}?+�'�l�.��*+��-���2m�[��n�r*�Z��N*f�9؟R�����q�\H�6Khb�p�1����9��I��${ȷ���������s�,]>�d2e�o{.U�o�@N�<�����װ;�w\ �v� ��z�V�c�%;��5������oKsB�7k� � �p��FV-��x�}�(9܇�e���ib,��� pԸ��f��D�(����-]��v���x9J�(�Eojy�J�$U�f����I3�s���:��w�Aԋ�I9i��q��Ķ3��RۂJ-oZ��7����w2Ե���Lږ�w��/����I��5j=%B0��9���`�?z�"u��:��7�N8O�ݵ-�JpQjB�k`y+u���s,�$������4�_oV��En���z����_�q�޴/���%wPO��k�2,g;��pRSu��F��ݪ̴��u�k�oVJ��&���'�};�񸶤9�U����93&���y��B�k�XsSy{�W��Ɇne=���9��X��^��a��"^�U��8�#Ք�u�cc��C��U�s�9j3%\�^�B��U<=�0�F[�7#^�?x	旞�o��hw��fuiήe�q���I�x�镆�I�������\�"���fw���:~��=c�����?9��Ο��N浛}����e$V��ܼ՛u�⋩n�s��2�7Q-���5A�)a��"�Уi:FqL��)fmvR��s=����՜3sc#FM`��T�x��S��;�������˾�:�g�͙/����gf�3�<ߟr�/�J�#�Ocz�c6���xs��T������e����Չ'p�Oj�_���yx�0��9�7��t��B�L��i��-�ь۩CT��0,L�*��k�;�:ͭq���K�u���k�J-u�мJ�����2�vzSV@H���];�;�S)VV�����3�)��GszH򔉝�;�{v��Z.���ɚnq�RQ,s|�� gRRm�����*�3��_�N�%���x�.AA��k4 ��3ּF'w�*�B�(Xю@m�� �i0+�ސ�P����*&}:\���>Pɘ����=��y"����=��.�W�!ԱJ�̼�#�DU\֎l9�t����竻YL�+��E��(��˗#�!ʮ���
��y�2"�۹A(!Er��K��y�Q�N��h*+1j<{2���&�C�[)�(�$P8X�)$��F	bl�=nwE�����\�Q�+t�ͅ�^��#�p�#���K�TYEU痴�#؁�B�/h9ܹC�		��P���p���.�.\�����y��$&��(�k(��t�����!" �dPA{��9!DG2�KͪUz&�B�BH$uX<�^�	p�HN�ף�5�=�h�n��R�D��&$�陸����ki��Km>��LZ7�˜iv���p��Ȝ������l��߾	
�O�R��'�b?h�Xt0��k�����U6d��E�|Qc�����#Cu�e{�5u��C�Y�"�+p�!�ժ�6i�Vz��Ǻ�j��H�ٷ:��a���Êk�͹뙏F�qڒ�o^�B��y�kI���@��Yu=ዔsn�a�3E��`I.�)��\b��Ӣ��vu�{��`����θ7z!+�[Vb6�b�f3�ᩐ�'Mz;��Okݚh��o�l����h��3᷐8%�qc�敺ɹ� ����BZ�O�H�o<2F�]�҄�NQ��4�jJ���� ��'2J+�J>�`�}���uw��=L)��g!\-2�"��<"���Z�����ƴ�zr�k��mFh��J&���G�,����C�q��Cж�^�R=�Yn|����P��{a���}G�)FXj�v�i��[��Ɠ��+��(�4���~��k��^�s>�zGU��qu���6�T,ò�������e�����������'��t�oo�����~���s��GC������k��k�{1e'�&5�>�Q�u��ϻ�m߼���{�[B�6�v��*��=0D�TPc��pZ(!>r�gj���ng*���88]!�lu�����U���gm���8&��W���.�ͷѓ9�جmbv���;.���7;f/����`s�Fɦ��[l>3��%�@�9dw�fD�U ���+����Y��.�}��D��^U�>_�y}�\�����041�u�xb�`p�lz�}�k���k�1��#3S]�ae5�^���]0�q|e��w|�������p���~C�>�N^��`�l��gEy�W��P��q�K5t��D��-.��ʳ�P{��P~GE���4	m��`v/�tK3�5km[��Y��M�U��n���:�[�9���8�Δ�̬�cʰ�E�v�r�Kߍo��R��B��:��0�V6c��G���5S���Ŭ_wA�u�ƬJv�������br����*����)'�������g�<s��?�uG���k��}�o�_^��[W��X�AGCsoK�e�]���[�b�i�^�8�#�s�e��Z�8Ф>/lg�껦8���Sv3�*a�9SG�$*�A�G�!�C oo�ǊHE���.⻽�V�1��!z����H��!�s䨹x<��̗|?����U�v{����zo{s`2����[�{�g�t�����{9m��WlrY{�?�r�5>V~m�ĖK�V\��������T9˾�KKOv�����cu���^�;�@�aL�h0=hKL��SB���47��BM6����m��גf�2vWS����9�4����F�WS�}C�n#����\��Q�D�8nrU[���)P�)U�V������՞35Y��
�	��}�t[y�ms�@�|~��0�h�+���\?T'���vk$'������݂��[iH�~��$�ax1���<��Gkf ��{C)Z�f�uj��ul����p���G^^̇���nq�ִ���	�:l�g���L>�ۦc^Q�zϔ4�qY�R��wP���=��}�q��sm�=�ｴȟ&�,n5� �� ���؈��$�%�x�ك��{zИ9/�4v{>#*��3e@8���{T�	Ɲ4Aa�4��t
`���3q/�w�kj`Scz[�)��l�nt�T[��z�N'INC�jG>�J�w:�Q�¦,�l���hZ	�.`>f�����+��C��T���9�;/��A��w$qM�����.�|�����)z=� ����19'l\�2En�6�[���;S~�NY�*z�ѽ��0m��_{�#?o�L>�1eb�ү��#���F�NEE�����ON����	��a�o׊eݻ�e������ ���~Ve���{Y2��v�z���{��o��e�a�t���VY�3�2�)*�Z���r�Ƀͫ�	����4��aa�!H��/�OvR�Ou�.�V�{'N>�'\=�	.�Cov�U�
`0��	�u��N�a�u��Y�^MB�
Ek�F�f��Ϗ5>ʼ.�+y(:���3fYyc�9� ]��RU�l�%6��*Ƽ�X����ݱ�����c�X�0�~���_ZS�;Kp�P΃*S(� �lS
5�o3	V����}{�����]C�\p��`���k]�7[uG1N1�a�Ƭ[���6:u���Yݪ��V��;�]cݕfH��h�LYƎzh��nCC���ϸ4m��?O1n�B�/�fz�q�]�X�䱻nit����gS:9F�G�Va�@܈(@@��g%��Z�U,�z��	uA��=�������{���~���T�P8��O�T:3��?�voY)��r=n���4�n��ߤ5�v�#:�9�m��p0s6ԿF{ƣ�ʑ�dF�-�+�����e�T�˪]����`R��T5�b�.�:�l/3�$b�sџ7J}j����\�UW+Z�3�#�E�./MWu�c�e0c��ֶ��N.^|�� PBդf�W'wK�xGA��C������-�O��;�t���s7��~��(���V;:�,����w��@�dP�����d�o&�t7{^n��Ӳ�y�����\R��i��\�K�m!oeʂ27[Bb�Ȏ,��&�yhc�t��w�pNY�l�5MDwn�u��#�����Z�;#�e�N��.�����G�k��+'��1������x��%��WS܊�,�xtgVdE�����V�e�ˍ��;!zz
�ØO�����:�3#'}$o��e���F�[{��Wٛn�ǟ���9�5_���+��
�D°�Cs��4�0�ϝQr��z���\t��bc�/[S��ք���$���=74����\��!��4۾\W���>�*�U��g�l�䈅y�l��t���p�����8F<�5J�	��od��k5�%�c�`������ns��f�/..:��b(����-Z��oT]%�lyk�4�O������h�ף�1�{��&c��~�]�ͳ��lC����y�5��.f�wwj0�W�~�g��+�ٚ>u;Iq`�g
���$�c�a���^0'q�:��Uv�]���T�%�.�a=�v}4f��6J���]�܆�	ҰMXc�;)�6��e���B��SI�A�]�:�U	Jj�}��i�LQ�4K�@�M��tN0��w�zi�:�l��'��R�r빡���3sS�BY�!�>QȖsS���G�pT[9T��a��S�
Ex�-�#s������ІV�9ʷ[)^f��۞��{"�6P˭���B��ʝ��C����c���M.�)�YjʳSz���@]_ar�u�ǌli��3�n���[��ݎ!� �����m�f�.X�5������Vm�qO�������w\B?_[�-����n�Z��r�m�lGX,����!M?G�yEn��l���Ə�����`�����x#�6��t��-�;@�t�}�����ɳkݮ�XÂ�{�`�����'���z���6�![?r�n�߫�c�+�ͱUoEթ���W%ת�cs��tm�y�}|b�#���,���q ����T%9ю���,�;m����ӑ�9S� �h�M�_xM�^%�/������ y�4��5�C�6F�9��Jbb��v��t�T�:����ut���b�🯘�u	O�"<+�Y6��غ��դ3�
q�T�{��s���D�Z[��ʳ�I�-���2mSF�����6�l_X$/Av/��q�nhx~����n���|����w�`�q1�V�q�zg�0UD��u$�|��F(��� �.N
}h���E_�ch���E�t�=.�t�ߍš�롿x!Dn3u�0�q�W�]l��$�}k����ݑ��{ƍ������q1T�p��k��jG6�!:�^0�c����$��������QKu���Ì��LĤ}��Z���yR ����۷<=�E��$V^(˪�y]�u";�Ub�G�?����/u:-
���qM����KSJ;�1E�@�M�!�6�X1QL���ǧe������~�-Tr�;ej>���W!#��*�yt[��e"�ScL����. ��ˈH�JTaq�Q��5��+ �
�Vw�r��Ý���t.MD������Z޸�ћmO�-�*���!sfm
B��8�^i��Wdl�����=LG�Ӂ*.^4Ay�%�0_e�+e��Y�Z��0�Wwkj�c�C^ؼ�������4:E��p[D{nk6��<���%�)iv�)6�=������6�
�e�E���a
ޙ�F�8ޏH���� DV���0�h�+��ŗ�f�=���d�eM��t�^,T^1�T��"
W�dt]�. ��C�����ǰ�����hi��	����"��e��O���\P�1���Z���k����-0�f�~�i,�Xt0cY���.�tyQ��������o���Ym��w�n]��0"�8�sf6��Ӕ�y�N��v�=��h؜�a#Z�t��T�>Ukdf$ʁ�������0N��Ɯ!����~�����OK(�n��ܧ.}K-̴���ԓ�����ž�N�Bkҫ�o��.����:�݄�Te�\��##�	�3��e�XfEA��f� �������j��-�Q�jsFY���=���_��+��)�$��o��K*L���zRTk�{���{8��
#���}������NJG��#��ĨV	�Qt6��c�H�Dc�����
z�N'INF3MH�r��(���{K�V��	�!���!����(�����T����X�켏N�wt�u���/����a��?>��T�� ����H.�Gh�fH�݆m��7{ܠ+�\����gW�ف�4�vO�P��B���,�(5D��x�aa���DΦ�幛 ���[y���ȿz�DwXHJr�+�������L��k�bz�����X�>����0B����u�8e�ʳَ�.�\�#>J�!>]��|��\˕���ڷ��6MTD���y;�L s��?��/s/�^�����{>R�2͋L%=�u��ۗmW}���_f������KӜ���涰�6���أ*��m�<Ÿ�|����Ȏ�D��/�I��f��+�}r*���l�hi�8��M��nZ(@HPܟpn���vWR#Ei�;S6���k(u�/5�"���&��)q�5�tv����B��R݈��p�������z��(�r,�o��ʝ!xn��at!r(A�5ie�mu�t�Vz�5��`��.�)��/�2>��Ə]UO�nH_�91��U�I�Y��f8�NJ/���llLe:`��	��ƚK6�ң�a~�}p�1��^�śz�ؾ�� Gйw^�g��\!���s���(qvL9�iyd�������C�>�q�;5�Nr
tn\'x���<X\��$��b����ýEˁ�����:���f˶Ϲ�O4���v�Y�l���I)ξ��~��'Lz�|���=�@���E�^g��)�=�(D>�S��ڐ���2ES\��c�K�B_��0%�Ŋ�[F�.Z��
5j�3e\�y �ץ�Z
{t����>MNU��j'��ϑ��8#���>`���<5��֘j��R�������5^��{w�c���AR��|��g�������k��>�"u|ldd�/���tWs�������t����Q�N�����~�9]�.5%)�	|�Dx)(��ʳ��?�ܦ��v/����9�+�]���@-�n���	!!AjSx��q0�U̚���/�Yxx��G7�� =ܡ�_���O/���~��t%M�!�A��hわ���'�͈����e7Gf��Ƴ�p�����?*;?|��S�W��q�Gv�&�+pf�ݓ��7e�"]�i�iw�7 {����3�R��5�@xwޯ�Bw�}�z0����<XP�kܮ��T�{�^�[�C[z�˨x�k:8�90%E��k+�	�=�������/h0�v�]:#�B����=����e��V�Y�����f>sD���J� �{f@JZgK*�����Uc�_H�?.�Y<�1��>�Ve����z�mY���Ȅ}F�������NM3��xH�P+�z��Ӣ�N0H=Sa�=lz���Up����	�� ɩs�:!t[�Tn�Շ�6�J��aႾj41n�9F����_q,a��a�^g��SBSPܥ����A�l�N�b�I�z����8�;���}�}f��D��>�0!;q�d��)<�����RX&�𥶠��v�B��G����ݱSy��fy�����Bf#�%�A����m�~��v��s����l	Xi��a�mˋ�/Sqprhͥ�S���5Ũ�ߌ����ġN4�7�8��~������q�1��z�{g}|�u�[r|�l%$kqc��C��t!��|����&�ܬ6<f:����W~�q���J1���5z�9�w>�Md�n{�Im8łG``wLy�#��n�(�	ڇ�b�+3h�O���~v�F`��G��f�������D�f p:���� bO%���LɄu�`��&���"߬ҙ#�G�+s�ں	���E[�S�Ǟz#;K���۪�C�EhmnL��kk,>S����z���;�*1�׮{f�+��+7N:�ʂ�3��{aڛƲ�h�{q�G�R�۸��\ȇ�yj��Mˣ�"y\��1�w�w������ͰB9v�v�3G���T/��W}u�V�S�+q.��켴d�{RGS�m�:��M�4Xo&K�;�в�N���7n5Y+R��jP��/-��S�Uշ�c.+; h���Ao3,�l&`�T�
�mzi����m%�l����{ϮeovOJ}��8ۧ4r��l9�#'p���OM7/��y��<S�{�a��[�����ϯv;�GU�?�^_�E�9Є��*8�e�ܭ�Y�m��g}�QG��i��p�v�`�%�w��*�r�4�FN�{w���+}{"���vc����n���R�IHf❯@+�(�!���{鱑�nC�����sk�$�&-��$�� T��.�ʋPC۝і|�/�	/�ͽ���zo�͞���j@$�<���3���l���z�����u�3�~�wO�{�\������`�.��2��m��Ѡ����xyg�5u{��zG�R��hns��b�.N1��+)���<���W�hD�3���P����a�D�q?'�m�-�S��1`�^����BA���Ѫ��n�M����O.Nz&K�q%K:+��N�Mǹ�,֮���7������';�eׯ��=�K���YS�6��VS�Mb_n�ڪ�֯1��H�w�s6ߗO%��U�q�.����n��>3�`��}�N�1?.�gT�x����<���س�z�F�����\�h�y"�o�O+<��/�;��{�O1O����~��~p�k�<�WY�^�xV�SWq�/r�!���x���Ҙ�v���G���4p�~@M������`��W]�h��KvݙUn��3|9��2����Rm9a�[.�s �n]��DqV0K=�=���W@�F�-Ve��)�3چgm:1�l�QuM�C۝u-Z��oz:�Uq�e��lx��i�}�Mo�0vv�Ϫ�EYGP�N���sط9��%�gJƲF�D��h��.��#��[��'����eܽ�F䉌Thۥ��#:v�����q�T�_t�wJH�m*ob���{)+�t�@�ͽ�e<(��inQ䞆���W�8:���7�>�����ss�N�V(AH1�г��fh�q".�^�w`ݡ���)���hl�cα��әQ^���ĳ��^"[�;��+'���-�p�jd��˧�'=���9n;�B��r��t�PD)������7af�����;Z��^	�FX���u�f�ni�m	;DK�3hN�],	:�2�/����Ո�t�zz�Q��5�������^K/�'sC�j9[Q��n?ć��g`25%&$��B�a�|�d��W�t�
�\�x�(���W��*��Pp(��oG���g��:Z	�]P9C�q�/��s�aE����zJ�F��/����:�>�G������]s��Ӑ�ydG��T�ζ���~*�<Ih%��G׮9�*��Wq��X�|y��$�I;�F��y�$�Гng*�'��Z��u�D�u�(��^t��Zj<�v�O�V9UꇣL��:b̙D�GD=����E�ZO:ǎb�����u��uւ���^�G��������W��]Kj�*��V��n��:�rnIK��3;r\�:�Q��:��&�s5�;���=��-"�;��7s��s\N}]��g�7q�r��2J��L�yg��Ϩ�*�eNc��9ʠ���p̪Ȣu5rp��w'4JU��(�"�!+�s��N�"��Pr#�l�CC�ܜ'��	�!�"n^l�r�w%���ۛ+�UP��2
,�!+��)Ā�@�I���R�~�F��ܦ>�a���p� M9yH
r6���}M��$��)tUt���A�%�����)����L��=<6硇k�̧�'������o ���<� R��'��ҙ�S�?�j��Dc�V�qS[e.��y=OxO��T�L%��I\���)]I��Hҗ�����
�}X����x��Αڈ�+Kr|�Y��'����WT^�1���g��4��9*a�hqv.=���X��O��C�d�`:�/��{μ��A��g����ST�vJf��8HC�=#��_�� A.����]��f����]�U!��>f�i.��2���۷]��a��!��4l�˹KOհRL`�ఋ
\������	/LQ1r�b�Υc�����_�+�M>J���]�}y�m��'c�d>�>�3�,�u���A�M���Ó,+���;��ལ�{��;RÒ�T&G�*x�G�k*W���V�vM�]���s���*ܨ�h���csO��B�@à���U]"U �pU庭�=���ڣI|v�L`Z��Onj������C5KC�ZF�,w��Az�78%U�zZ�My7�RCc��ֳ���{����A�쿫�L#����?8�)��~�3">vze��/&�����Sti�����?-A��z���=}�����Vya2aG::�c�]o�������:�f��q������v!7��=���H��廠�Gé�nD�Nu+iT1bs��\mkX�N�Je��VJ�5�ƥ�����-�!�i`�gRZ�/�۫
|���ȘP(�E��aM�  |�'\��>�Y{�l��o#�$'ȅ���&}�P/G�SW��Jx���
v]��V`i{�r}�����PQ��]Cx���<-^CR�
�DkZO�lN��}c�6�!i��^+���ݟDU	���^}�(O�S� �K�H^��pqe�7�7ji��� ���`C�b�k0eg�aF�(�����	p�U�rG=+��U����I�WC��ð-N`�����}/(��z��_�TV�^��MH�ȁ��~��AS�~�c�{U��ս��:�Gt�u��=}D�2ڳ�;{r�B��sHF�=�0�|��}hpm�d�C�;J��B��\E�j[�먻}��¨Fg�R�� �	���r����Y.4s��������\�2E&���ɣh-.4�9j�h{x��c��p�St3v�-�>g���ǌxa�P����EB)���S�������^Vgs��u�K�w�^�bDwXHJr�i]B�&��&���G��%#����Ӳ@p~DD�ܤlL�a���{$n�bj��-�kH�;r�@���W3��V&B�A[{�b�au�\H���Z���5u�:�t�bs!�jm��9�%�X3����qMU���Ǆc�oI�4v��E��ݼ�c:<�]X��Y�z�c�l��.���RX�ge�VĶLG�����T�s����A��p������ٟ���3�> ��PL()��L��0o3�o��Th�د�s�9���bh+�`��e{�8��e�b��q���Vw�΃)�D���cSSR����7��rC)�� ^]�Fщ��S�E���p�4��Q��FL6��B_�yh_K/r_��O'��ϫ,����E�w��b��X��/Ý���N(Ǧ�{C[�Pnd����l��j:�������LK��U>Eٟa�.�5�Ⴉ�lNv��r���UuE�~`��.��@V�ݮ����*Ɨ�RR�hy�V��t��~�����n�nfru�iȰ������\�1��a��������=�Q�R2�޽]eu���=�W������8<0p��1�|x�}`(D-�
ťԂ��{c���G�����2��ZS�om��!ݐ�"	�����y��L|�����B��Z��ęW3�}ݣ'Ew������x��B�ԍ�>V���h��A��;q��ں������߹b�6y��qg������J��>N�����ڂ�p�#���|4k��>�9l)��}]��Q��r���u7hr�K23	�!��9V��i�@��]k]�k����e
��y/�Ջ���C��h.��"�&U�^���r�%���{����\��kN�ǫX����w�9�������Tw����J��mx>��;������}�}�`��șC"l�M�(*�.28�8�Le�.������<�����}~2\F�w��9S�	u�u*��w��A�(츅j�DµB"~�K8U,�lo�g����(��N�����A�/���3B��ZS�'�Btr�HJ����PG`��/�M�{�ca�'ZiF�VJ�u��y�b��d��K�u�S�{��R���:����N%8���o���t����G���?�>�pTv~�_�5y%n:v�Db������T_�v:�߯��[����AV:��g�5B��������հ��G����&A���4L1���N+i��/nS5��7Ry`�=ˮA�Ȥm�K��K�"��`u�~{!de�a3{d�����跟Gr���Ѓ&�R�jE��׻>�3E��Y6N.�j|�w����^�,#SD�g� !/ju�J��츤�%��	�]�ʹ�(��T Z��=�v��W-�s3��FP��LF1N#�D���k������74%U�xX0�m�}s���;�X3H+w�o�0�o���9O�������i���[s����c�T�o��L����4�{��;��n��Fȥ�`���Ic���X�֣����ou�"5�hOJŧX���O��ʜ�p�z!m���F����,�HAW�Vir�w����t�(�s��3�n���"�8�U�ܱ�c']'oJ��˭s6�0�h58X�>�߫�f�d@P;
���a@�Q@S.˔�)��0����9�w|�]���}|������7��������:'����� ��!.74��;o�T�Z���F��v檲����۵m�f����t��4\���ݰ�`�ü��<4��촒�!ի��걨���9����sx�f��ĊP1��I�L�#d�l�y%�k���=�e�2�3톫���L�ޞ������n��~V�FwSsЇ���l����P��5�D��+�!��t30;�����_K�W�|r�0o�p8�kV��l���,=����t��� �>�k��>ͽ�My����X�����ºX��򓦡Ξ�D��nBAʳ�qa���+�o�xB����Y���P��(�sH$ 4�X��y��G�i���w+|�şD���{��P���z;�b�0�z�ZT�E��OM��;b	A�h>��t�͘��<i[�ݱY	��u^W;�������?DQ}mL�!�]�Q��d1E�A68����ˍsb�K���ϳW�'5i^����=��?ySbA��p[�b �>���e��Su��	s��Ŗὐ�üa�O�<�����{٠�ڦ�~�=�9��-k��z^5l�����vE*�0�f/�X�Zz*��K��'���?���Ю�PlH+���#/V����xG��.�6��}�n#
c��S��`�7e�!`򓨉o%��?�@�0�� .6\.2���#���ap|�}~|�?>>>��Ǳ�#�����4�X��HJ��M�PF�@�t�N!�.�c��F����ܵ�
�SsKֺ�ݻ+��8f ��4M���Ŷ�1������ef��QT-t�Sm���^rݖ�U^��׼E��ngc�x�H��/�;5)�r�7nkH:���_yw�Z�z�y���{r^�#�H����l�:צ�@���� D>?g�sB�<��f�W�����N���(�^sA�x#�-����I��M0���=�<Ӵ��fᕎ��ӹ�����u�,���#�K��:Fw�a��!P��1cJ�=6j�'�z�f��J�����pBv]J�'�j��� ���_�}7[sxv�֚�l�,�W�Tȇ��9�{��d�p��!���ABrG=+��U���e@8���xvᦳ�ذ�F�������q��D��F��mh��}��F��Q��ս�ا���ve�r�=���ިج�ڌ]Fڠ����ksH%yP�#�}!�������:n!��@����6>���Y��>i��|�nR�(�l��j�G.T�����G�7�,��mR����{����+XƂ��t�͹�?i���ݗ��/I�'!�RCV��|4���Q��.R��Ʌ./��t��K��B�J0G�}�*M�j�md�U;�wyE�g7g�����}����p)���`\�����7��Y�=v*�Un�_�N���J�'u
4>��T�����P��N�w�Ye?Nќ�A�S�O���%3n���-ɶ���s�m��r�����~���ne�0"������û�
5��7�����2C�
鸦[{���h_�M�		)�b,��Xh��~꼗nv�xPxr�Cҧ3y�y��X�>)��jx�͜��F�6&����rCya��H��Z#���;���$��}�!�٦YNr}�,\Xt��(FCL]��Y5�R�7���]���u[�5���Y�=��w����/�Vȝ�0=�yr��
jl��~h#KN(�J�f���6>��1Mg�ii�����W�1�\��3 ]{�G���Ș�c@DGr��!(�І��$���F���j��2��L܃��nxERQ��	�Ȼ3�,�2(�/ �d���y�p�|�8� ��0ʶp�ڏX�H���"���RJS	���wF�.L�v1[�G<\M�݀�����Q�}a�O�i�ElX��n�Gz��9�jX�m3������\��e5��ڿ�x����FԪ�D7.�:ٓK�[���$�}��M���$��o��;*g�!"g]�!x�L�~�f����:٥tjPi�],�����Ψd���1�c�>�BV��6�!Ĵ�8�V�{7a;�Ѣ��I~�`����o������0����6 �f��f�����F��)6�y�$7 �W�*��_ԅ8����
ťԂ��﫞��R�2��S�3qfl�m9�iW����ڂ����?���;=��KЍ���դem�{E�����N�-[��*`�.�4���F�+qz\O=_q��=��i�x��쌘��J��M���͸zA>҂�f.
��]Og�~�Ph*Q�!]�w�z`�����zy9���#	]�EQ�{ܐ�j���=���a�v���\gq+��$r��?.ˈEV�W�K����9K�9�^�d�@���φ��G*����=�8���g��,ГϠ,L�cE�<�Ӷ��h��v.�-HK�/�0q��_���z[_$D-��S�SbKb�������ll�.oT�f��VxQ�'yr����?42y�a�5������)��v�J>,��%��y�:s��s�kQ�1E���:��N�ͽ�ZM�}//����W#ms�evog��07܌F�S��y�5�$�o��8]k�&�`�g
�率�ݴ�1)�'U>J7�=�b����t�e
�Ti켩��+�v�u��ǽ�&�2^xŏΗ&ݴ%�w+K�T��퀟5iEt�y�e�rAaL���~q�	y�+vNV�vE�G�ɗ{�&�sG���z�{|�I9�}�}�����7�7��=�Ú:����p�k�C��p�/h�}�^3�+bj˚j�����њ/�E$˧/��!��t,�W2��\*�v�4@���$=�֐u�r���mY��[e�L�NFQ���i����󳪖�↚%�k�d�x��a�`�m�p���2u���xER��-f;�smV��ķ��]�ކ�-l�ܟX���f��Bv���؈Q�	ȏ�R�/��k��/6c&���;����QO@�)W��>��l@����P� �5�;��-`��oE��ț�˅�;x�e�;Mm�����tT���XG���u��"��ʉ�"Vz�_:�E���;������;o����U�\bi@�Nd$��Q�m�G<��6�&1��晻Y����ݬ�������e�S
z��T�T.�G#3�ە�]F)T{����,ٙ|rHl$��ot�m�Ӝ�8ŉP('�n�6y�j:w�X-�8�S[g���|��ؑq��\L[�/�j�V�����v@��A�(���8�� �9�nt���)܋����x��
I��*}׶��8�����P�[�)�ۡ���pܒkA�BF�津�Г:K�7�������+����w������NG�L���ᾳ׼7cr�F	B�v?	�}�@�B���q��k�C��΄{�.�d�4����߁����7��0���,��T�֫c
��-<�y6�)��C�K�|�Z�<�ʣ�-������n: o�Z�ߟ|���Y��eߏ���B{C�..���D�#�|c������'k0�,z�j6�l2��:�Ǟ>���%�4��-m�g�����I1��M�k�F�5�L����l˵�8�\�؍���J���m6� D�T�8-�5~�#�y�Pȗ9�tp�� ��L���Nx:�q��c!�0Q.�c�{�m���F��=˦�q�ǉ~��7���E����M���U�pT$eಥ���EL;ױ�>�S�"z���Ĩ�uD,��:|(�x[����6������Qm>�zs��{b�@~o;��hAH�e�mn�Yc�1�D� oq�Q�
F77�_��.}V�)����EP}�a�e�^ŷ���� E��B�MT�J�
<�����������9U�����)��<���Bϩ_��,�ȃF0����6��m_z�{�2��}NFM��c�d��pם�v]7%{z)�m�5�ִ�x������� �!�P��t��52pz��\��GX��� h����[b�(�5K��/����9�z��&/�d�P��cˬv��;���')��-K��ro���J�F˕�]��>ʌ�0i��c�Sm"(�IO���%׃���#h�x�F�*Pk�ɐÍ����㰎�i��a;�V6�Uо"����>~*��י�c��W����G�K�<��Ӯ���D�L�]��o�A��HJ�(�Ͱ�����vZ�GKíRG�Kр��ɸ��+��@�}��=�:�-�D�V��ڏ^:R�@U|s31��#�Ë�s^-܀����bbi���yh޲%��IϦ�zwQNf�
h��y�e5�ɹQ�ŋG����M�4�\�!��nWv5�d��jU��:�ܱK~Gg�����0v�/�Ɠ�妌��eix(}�_
X�#���b�Ƴ�hSh~��gb�O�Q\:�m�,��˺"Soy���ǫ���*��"���������>�۴�
nWN�95gH"}�ts�����ʣ�w'z%�I��im��변;�#A�\�b�^��[W%Vi͉�6�1�j����ѧ�S�x�ߣo���wn���.n�5����h��4@;F_j��;���Ex_Lѷ2�Wnc��%�6F��A��!^�F�E,��L���~vP��2��Ê5����{'pu�c
�mo�"��V��9��`XY	k����I/����q��i?j���/���x�j;{X��2�ٮvz��H�M�΃�+����|��9�G�=���"�}�dt��5s
Y����ә��oSBtr��<Rf���כ�+�t0a�o�Q����>y�o�#��Q�Z�N�ٛ����{�k�wkY4+���^�G�A�Z�u8[��-�F����.EBB�e����P+e���G#Tޝ�y==S��u� #��lu^�����r�*��D�e#�:�9(�bB�������^I(�ôz���]{�v�-����ӛw�=����Dt� �_�<��;�^�u����;<^�o}�;u�G-�PwU��k!�T;��%�;�C%:��L�(3�v�}�������:tP�oS��8UD�e�귐�C�P*�;�c ��Hs.u�'}sܻ_u����kR}{$O�������?~�K��{Z���~%ʒ��E%���Dd�s�>��gmut�`{s���&�K�ѻ�T<@��m��
���gi���5��M�
�/3)ތ�7Fk�( ������#��$|�ל��{�\�a?��v�V'Y�s��%���s�ӧ�	����,�R�ąf�Q�\ �r�����.�g��V���JEמ��f<��Y~��&	C݊PomH	�\b�����@d�[���V�~X������_Z:_ fI�n�}��&�ử��|Ľ�ەz��&T�����Rn�n�Գm�]�]����pdӻ��{Џ>��x�?�~�� pg�@
3z�]�!>I*��z�U�I%T\MDT��dT!Ю���z=��c�i*�SC+{�!/�9�1D#���!�QEEp�'pL�F���IeW.\�q��z<=��-i)��.4$�FV��"#�m5����T@�#J$�]!���8a�EAv�*H)R����ZQE]��]G���r����E�ӎr���
%A���@�RJY����g.<a<Cΰ�VQ��T1.f@Pd��8�j�`��H�+[�ʛ�$P$�e���D�SN*�ĊH-Rj�%�.�

U�3X�AUEV��J�L�-c��mU1�$�X`��bd��F����24-9IЙIS*擮N����UEQ��!�kZj[*�&d�nK�PQ�GN��M�uH��I+�̪�b`�HO#��Z��aȮω�Ij5B�ZDU�DQ$�D�yU�AX����{�o�9�s�3����؂����Ȩ��I�;�2L�fެ-I:4�h��i8`h��N�]�/��F�7���7�������{���i!S~{L9�ۦo��J͋Z��z�M�Ym��v���	�ic<��W���Uo�я�b��\��'�X�.:�PQ�O=/���V�FbL�_C��s^��3\Z����=���C��V��<��B��8]t:7���[�v�����Dbwc*��սVSofZ�+׏��(+��-�8�򰗠�/��W�_>^��a�䝲���N�&�x�#��@�}�R:�؜*҆ ��nlc�Fx�b�X��	��jW&�w��:.�uʢh��*�FS�G�*~	\B�������+�[$%w0�I�*of�n���m��>r��t��U�lȔ9o���7��F�p�1����#��BO�:E����Z+!�pJ�`¿���O��ٹJ�FkTᘎ� pz� L]�F���m¬�c��qA�U�ׄe�7�ޜ}(�wsT�5��L�=9�0����"���[U����L54��@X{]��^>�#A^�̬^3�h��VQ��El�;א/.�J;F&�b�z/��Y�)�"��]��h	�L^`�=Q^W�HG����~#X�v�-̸�D�<����� ��}o��Q�v��#��麵p�WӰi�2����Yӌ)=��޽�KO13)�j�Q�*v�Wߕ������B�Ս�����=��\^K'N� �`? ��l�ܨ9v�=�|�{��� yբ;�^&jc�'�^�n=�����^T[^#0.�ՆRf�+(�����~.�[ޢW��뫞���ı�3/�!b��<ŸX*�/�`�C��U �fp�FE'��nw��)��X�	�[�	r���rD��������!"�7<2EX����.���=�(���槻9of{�)|'b���#�T�>��BءMe��ɷ*�s6Կ}Fq�9RYR�TW\�����=�=��:�AQ���<%�p����AKmԋ��z���^�nM�2�����L?m(D>�S�\��5�������!3�~|�����G��5���K[7;��-���x��t�3I�J�07N�n/O4�kq��;�} ����r�R7n^D��[E;]�E���W�]o�>N�Jr�;P_�q~Ud/A�+�0����S�deO�C�w���#�,�4t;7Y���e^�R��;�%`>�UF��IV�A��5�I�PL����H��{�c�d�#�+�D�_zڞQ?R��PZBT~r���R�6Q_V���ę��{1� j�^�n�q0Y�e�/k[���r��5�'^��d��j3�66K��Vs-�7W?���G.���}Q�w��w)4Vm:J`��vR�eyׄ�l��m�rU���r�<�23�l�����p
5�srg-�;?�����o{�x{�<"�u���l-mo����ǂt70���4���z[@$D+t��)ShED�g��������Ӻ��,1�Fb��ϧ]��O�<1t47<�&�#�g$���b���i�t%d�b�Q�5�6�){n9��U!��A�Ȥu�K�a�.(>�4 �4<�]�r2g�Ԛ�D��%{�_��ySf#py[�р�Bk�I��/�CZP�)'�>��$����{��)2µ|vx/h�c��q�]2j\���]�Gkݙf��m�׏0D5Ly�vO�`*Y^�2�%VM6$��m�y��'�� �W�j��ˌP���**iWz��Ѥ�˧�����er�������n|����}���� ێ� ��)<���nx�޾\��iI��y����"2������G��;5�Iٶ�lpe=�X(p����\1�zi����#,���FɌ=ɶ�@�)W��>��nd
1_T�N4�6�����w�Y�澗�u���e��q�'���;	N�9�\
K�O	�A�}j���;��=v�S`���f�6gŇ�ѣ�[O�h�Eݠo^[�oե�{7&��X���)k�P��0,�8�.0�����N�ɝ�,�x�U�Mٜx*-�U�D���$�E�y���r�.i�\�ZU�L-�2�t��zQx�������ϳ>�0}���� <=���l���#�p�צ�MĲ���:�C��J2s)>�l�m�y%�_�U6���z�F?n(c��}�-�p%������}+mX0�Z9��nT`�V�o>yc����SQ{��7�;tQ�[��f�%�7��xÖ¸϶]��ΑIL7x��2�^���׽B���5�^̽>yt�N�O�"�(j �;�N/�O�A���m{�yo���T��U��?������م�b	<�O��e4�����xcX��aҋ���[t6�r�5�t��׼P�#H5թ�	E"�;2mGI����_�ÓA�`����Xa<��;k�b��N�س=�_?�U�i֔�	�C~�b�v1��=WD�f{��
���X7�}��2�>0qQM�ؙ��ڼ��:lH?c�!�f��	��I��t�,� �3�s,��^p�8P�$���. �?��|�L�����k�tơ�Є�C(��r��Ģ�/�E��Q�]�+1Z�F�n^���8f>МT
Se4��m��Lh�<u�ef:S����nm\~��I�}3���?!ۂʫK�� ��<:l���	�W G��ñ0���d��lPc���%���U�\�� 9�l�ȼ��Z7���p��f������p��G��C{�:�(ʨ�{��C;��@��c�U2P����~^xq���:��>^��la�l#�6J�ׇ|�#+ �_@��a�[Qm�i����~?��Л��#Cr#�޶��1A��A[��¦�i6م����E*�"*�}�am�O�-��8=�9HZ�f���dm�r2�'��CR�����X�:�4&:����|B�W�g��a�EE2�[6���͖�i>|�@uT��E����+��_�鄌��S.*ۜk@��h#�'LSݻ�MYQo:b�T6+���-C,�{�8�&�JM�=+�
ť�$/[�8��1IG7BˡV�gIUZk��3v�N�ji�%��B�F�Ǽ�G9}����M/H:�*W*��������:sչ��oude�|Ts�N�9"hl��lwѱ��
�"Gj#eǳ�ԙ6&�m����OY�zGluwK�)��	��C�g��'��4?��CX��RO��}3��u��]>^�e�w���`t����Y�^n��7
����+3_pT&�24\]�ta0��޾��15Oҝ�B�K��:�|T������-���Ņ��H1*W�2�n�����CaٍjN�tyY��N��-��<.l}	���M���y�������F��p+�dwb���+���{��yf�8oZ��g'c��r�̖ki�P�y�dC��(��ki�s+����o�ԡ[�O����w���o�L����߁���0���o����Z�=c\���0�6����.� W��bD.���t�i]G��v���&���r񵢴7rk�ɨҨDH�t.�B�H��Ź�5�9�Od��bj�L9�q�yV{�z�r�j�:ņ=���V�P~묩du���R"�測Q�]^��ji.pm�`��u�����]Ք�ٻ:��D��}^Յ�;�7�S��C����Á�(_Ly��gP�/>����3�~7
�a���Pp�r �����]{���i�)Y_G����@���[,���g��0�48���j5������^J9�b��&ި��Gb�k5�E�Y�o;X��P�GQ-x�q���8F�O�ݱ	a��*���N���i��`°�b��fj�,8VA��C���:�=U(��Ɛ�Vŋex���Qe0���Y!m�ȒG5e=�ˬ�؇�����PG�"6jD��Dz,W
q����b����t���H<�yl��9\�5��n�dv��5���-�s�(� �r����cK�|m�d��S��.h��i|kP�WCp��#���-гZ�������`_�i /Q�.=������p�p���j�.��o�Ds\�z��������Jd�Z���9����pp����+��T|�ą�9,⓲^[�3����&o����>G�O��~c�X�67�@ G� U>u]Vy)bb��c�ްl��s�T)��PV��� ���>����J�3�2�?�-J.'x�=;{���!�}.���:Jr�J>����&�+#tr���&��W�嫨b�ÖínY��W<��:���ɡ��'�%���w�]-��g�ݳE��^n<*Z�fA`h}F��^�vGd^@-���︿����;:]�{2������UD\���;�(���cYA�-.L�<�����Eq���)ZDB�����W����U[�s�J�%�;�sX���ys�o_�?42y����͜X��������B��Ȭ����#���� b��l1��U"lVE"D�ha��}hh�	�^(Q�5-���ۃ�sW�'Q�3�3�q�96c���b
�&�D��s�K�I�q*1���W5�v;L�h!,�� (���B6da	\K�0�wP��IF�M>�%\��kݗ�7�������IU�n��|(a�xoxXM�h�ؒ;�a^g�:Xr5*�ns�ڳ��$����J�͋6��<y�8
��Ӟ����W�>�9���9��u]z��}�>[�ny ���Ӧ����_�3�f�p҄����{*Y�rېL����)����l���@B�'v\^�"g�����y�o6{T�;��U>���O�`���8�m��rG.FN�j�;�i�Lt��D��Λ%�8�\��L�8�q�d��)y��&iYii�xOs��b�A��ڂJSSP�q8����c̛3���NЛ8��X(���Yڈ�(�`�����{"T�=�Ǻ|Qr����YzzA	W���L@�|x:l���ج3&j���)^�ۯHkB�-�����q�<�;	I������.�=q^��9�D�]_�8uV��`>��^���*��ߙ��m��>�caԐ�wI�6M��<��Es!���CK�͂��^��q0��Otة��g���`�T���u�*3�Zɶk��^{�FE�+3Ϸ��f���D�t'`�X ����Z�ƣ�Oݨ�y�p8�5��Kѵ��ƴ���E+ݨ�^�W/8ɲ��Ȑ�ۣ�`��
!�aE�Sѻ$i�s��<��=h��s��W�wr<�z���@Z��l�:,��4	4�X��O�xug�ak��ЂuW!�NV����j$6�/�4PJ)Iٓj:��^Z��y.� A/��cǸ��\�e����F�Lu�򼪵�C�u\��#�X�;ۊ�Ap�f�@����<i�~�7���||a4�ag8N�avl,�w��^n蹗o�Dw���i�m�����1��Fv� 	L��ٳ��P��P�L��ӷf�Mu�!����X��+ll�  �7��<�����T�k�fV�@������V�6����y�w]1�IL'F�5sϺo&�����T�W;��V�J�N"|`��!t�����}rؑ�14�jj��բ���
�c��O����`��C َ2K��qp,:F20�bg$%B1�A�Ý�TÚT�
�5\p���	tV��c��c�D�]��	������p�B	�E�q�A�,�h܂�ܬ4�l��F5ں:�����V��הz���^|�p>5��&���+�4,R��:WS�H���E����UQi�]�ܢ��[&�Ι"�]�.�I�$D��l#��P��x<5��˖�g�=٥�//�F�͆����4m�v�}��5_�#�-򰐥~Rf}�P(Wv/�2
��U�_���1�8!]*xl���
VȨk�!�6�VOܯ!�~�tXϸ��[��j;��'���oQ���>�1F���L9�ۦDk�=]5"V-.?/[�#[sv�ܼ��,k�n2���<o~���]�w��!��ps�\u���4z^#�1`Ukda��^$EFNf�Ͻ�F��2s���`?]K�J}t���q���W,��@W���\50�?;�7S��BH�</'.m�D
��@ZR-�0:R�-�%������@�Z����q�o3\|�o�}�R��"��]�8����juz��|��/_c }�lam��=�|���9>O}���l+�;����dM�<��-<`c���ꃎ����}Cv|t�~�nز�^�Gb��ӟ']ƙ�\B��Íz8`F��2u��C(�*1�������
ny�7�G�P:
փ����Y�^�A♸P_P�dq�ǣ�	۽ƻ�5юϕn_���i	c�8�{'���������J��iL%Q�A+���L*��ۻ�*�c&[5Fz���[�­B����I���y�q�2*"��vY�ٮ�n���6B���`݊���jS���zkG�f�숍�T.��X�0�z+Fex�5n:ØR�dm> s�c;�3r��h�c���h���`��)�̹V5��~aA�"��測�TkWbfeʤJ��f���~��,����g�X��Ǆ�&VȒ7��.:kڡW�3~5v�����RwI�G7\�	�}�P�^���<Ÿ�%a�8��[^#3�׻>�3Q��D�M�m�FT���˷E*d0��t9��ϐm����Bu7<"�~`����E;�]��O��d�N��Fu�����^WF^w���p�+����B�z�'��ټ����5�ko�bwz5v�Sqe�H��0now���n�5?{����V����'��լKµ9�IL�a��
�6�\��sK8�ӎ���d�7)��`�`��3Ee���2�ʵe=K%��(��f�X�3.@��uxA���u�$W�Q���й̯��?��hS��g�-t������������˳���k�����ͩyOR>��r�m�\,,hܨ��m�Y7��Zt
Y��"J]�놩����Jыpx�B5�v�sq���7�7�Z��;���ru�ڌc��	���B�6��v�a��C ��B��FȳS�b�[�4g��E��z7�c�i�Hݦ3F��cҐP��47�5(>t"6eu��0��*�=�u�.��<�I	��2�7�I�¸���e�i��GDwwn�s'[U8�R���n5{b��-Qu3�8�}���袧WhW��WQ�B�®9�ga�iRf-�i�֊�XOv^nr`b��C#4[�����p�� �yϟ6-ck�tBQ�iI�E�z���<4.���!�8ǽ\���Іɽ�m�0;;��>��~��۰X~��ɹ&�.�����wp���E8�>�o�֬��w��]�sd��^@ۃy :���Y�qa��h�]9*��#�4���Eخ�q㱕���6T���p����V��\�v]��:
:�ܮ��w��&�b(	o@X�tRmT�v����"z�Dn�kQ��f<��r�Z��G�vs�S�sS�pWGats��;���=���Q����Je)}N���1�y���m:���Nt�Jk�ek�����oT�L-T*�G.7��eٜ�Ic����5Q DDV�K2�&�1�H��'0�����'A�
��jz���'�6I�9�e�/o���:[���7���vJ^�!��06��d��?e�C����'��:✳���ܬ�
h�}3�Y,���(�+�����:ܗ�`��^���r�3tS�?Zx�su`LLn�۾�GZ�_��6v�-�[5�
��;��4���P����R|�vt~�Us7�:xSz՜N9I���p��W�L��$��Ff'J7�ڏ�h'y.��;��=�_�09����]�-�!,l����7�<�C�si�y���!*����O�\�^����qLuU��U��g|@�ޭn�&�w�M���c���`t��^o"�k����6)t���c9��6kf��[/J[Ϥ�ybF���c�v��[-�7W���j��Ej..ǝSL5og�Q9�a�&�\�y��S���]��7G����ND �j�����;��G�0N��x�}��ԺI��X�j"$��X�d���3�z�K��4���1�&�G��-hƊ�\uQ�{r���G2NN*S�q�$��kZ��#� b4��!�˳���J�r�CJ"3�J+55ek �Q3�%d�*U%EʹAr��g����=�!z��V���L.��R]!9DI� �J+!��)�G����3��%uUH��̨(���E���ӹ�6G#4䒳1�vӔ�L��-j���n^�!V��\(�Đ��<�9�IŕGdr�R��VeM�K5�Y��L
�+�B*f����	'E	�\��4�譜�G�˸e�Z\J��e�t�WC��"�ʖT%t��L�*�p�L�IM$�9AZ��j�k�qȤ9�VE���;+�刉2�X���H�9HUZ2$�v��e�S�P��s�ƄGIVfVb��Q@Y
�%ȥS��n�	)*F�*9����\����G!)�ȃ(ڭ2H�
�+1$I ���EęI�
.��Œ�re%Eˉ����ď��}�f�Y����#�e���v�֗t�/n��:�$,7}9� �<\��q���:B[�H��#)�{��/�а���P�u�MK���oxx��=�D�|\�z�q~?����
�9H��gm�p���k�E���lM�K�׹��T��c����D�U�}��<����#e�B+bŲ���ޢ���a��FH���M���غ�k͏-�6�}��y�Ć���&(0�#�uuuB� �����Z���۸����ojF?�x�������#���9֔D\n89 0o�64����]���O�-,�kx�[�y�֍���nd��w)�3I�J�07N�qzdq��J�8׍��UkS�yA5H<��_u�@��������Q��;g�K���M��A�J9���<ͼe���e}�C,;���/��u����9l:�óg�ϲ�)��B�'��>�������g�-Fu*��UYb�W�=Qx�<�V�v�3��+�1���K�;>��[#nQ?R�s�бܲ�,�vu����8ǐX�I����ϐ<�_O
+�i�l���U�阰K�<ӛŹ��p)�o�� ��K@わ�w�;#�9C���eG���nP̛���z��tx)���mj�|K�`Me�z�a��SpJO�:�����w��0���l�nf���C�����m��C7�h��a}͘� ��&Hu���0�}���xyI��/�U��nn��Caef8-���*>&?�~���7���<<=��ݡ�D���Vߒ�wk1F+p�v�D�ٷ�H�-3��_�>0ҥ��}-���Wf|��b{��U�}J_z� �m���%�zaL�9u�7�(�4]HME�c:�ۚ0�tLL�,�A�V� u�(B;��~��s���!�Ƭ��m_�(g��z�v�uޘ�T�������h�l�9�Ǭ<0W!���� �mF�=L9%W�wO�_�v�������;��_�4W�
��(y�y'�J�K���Vk=W�#�/�l�a4C&�E�S�U��,jͬSF�q�^`K$�&�E��[A��+O�8�f��J�Ddhe�J[#T3�O��{��E�\���0,�>UE�~��YO@�Jq`���x�郄���Z �Ʉ4$�I}ʠ3�o�4����-wQk��JU�y�C���N�՘au���CqZ��V��]w%n{Q���vN��cn�Nq����g��Sk�v6I���2��m��4�Zg�=Ϳ�e,m�i\K|.�D����lTDq ���EZ9��ܨ��d�B�c!M�y]Y]�1(W5-w�V��׷8]��$K�a�����ǰ՝���{�,�����U���h�bJj�=O�.4���zs����g�fJ����	�u�m��R,w܉�����ED����]�05eܷ����!49w��V�=7�� =�ox0`<=��7�ʔڥn����)�e��X8@�[
�>�g5]�=c>��Gs��Wg��ۜ�_f{�bԿo_Ǳ=N�O�8���9�t*~�Zsʶ��o��/���8Ɍ���kg)yQ|F�#�,rhd$��!SH�@����pb�a:�|����߃�=�`�NLe��*�Fy�05��n�m1�}+�(�Z|-C2h����{C�*��Z~�Fe<�{��2@�]��5�t�����lŶQ���y�w��Q֔�ta��j�,d�c���bY΃�L�)*4f�uΧ���P$��q��QL���G�kq���H�΃&)L}V����%����:,���{�z�ߤ=n��$�.1*��2��>�*��U�M#u�G���Ȋe�\J��w���МqB�ŉ;CUM����i����#(DHa��Z��h���l8DC�3<�-�=�q8{ڇñ��	�~y|�/>d�}��<k*Y�ez&�)G����w��a�2�]�!��n��_��@W	��Jd�qty�E'P���.��YןLW����ݝ��ˌw߸���-Ct�0I���vM�zc����^�|��v���Bݻ���y�A�k�-�u��g��Z���h�2�V1M�\f��ʹ�5�q,��{TwgF�G���0nӭ����ѳr�I�D�^n��Ÿ]���<�(�>Ͼ��f|7�� ]vc;�M�D>>R;�0�X�+���\?)��<���)@?E�3V�|쨷kE^-ܥ�]��! �mr�;>فÌ�8�]j�na�9����UQ�Z{��48��]����u���wk�Q.+Qρ��x�@���b8AX����o��5�=��'dr#`Z�~��K�U}�u��.�e��l�&�Bm�l��TMȮ������Yq)�U�z�z����ǚ*����g`Z�"v�9"k� B��08��qMӡ���¦j���Ѓsj��Z�$V�<,#hq�ZhO�i��5 ��}
�^T O
�#ƻ��Y.���hW�s����BZ�~f�����子��Y�^�A�7
��A+"^�lk.����x�ТU�p_�>�pj�%z�!�hw\GX[�%2)ThJ����ׯW���&�ذD���j؇1ej�ip�B�.j|��t�����D��ެBh��HK�<$���6�6_l��J·h�����,\3a8�������̽a����{�0���ʕ.T��k|���6)�DBP8)���{��r���a��2p�7�Cؑ���1��Y�O%�[��E^̕�ƚ�-)a���JY(LzR1	��
;��r�mD+���D�E]NԷ�.�w���w���.|��>>��S/��<��0a��f�yk�e��Q���r~o,0~i����.]eK�yb��������x�y���$A�W�y�����Yu7U�Δ!<xAx�["O�#� ��G��)��^�'�r�4G�-��u�F�t/fV�h^���<Ÿ�T5�4As�[^#1u���զ^��G~S�.a�s���#��~0i�ܴ8HmǸ6�|n��!7.�ԣ�&�:JE!�m�᳴�fV�=�xz�҄�3�_#��leg��N{:��}�����G�G٧^=����<��跭W)L'���5P��lgY���a�4�%�B���]IZc}[�&k,������v��0Y��0��#�y/~��%���Ȝ6��=S���1j,�Ӣ����0��3�$b�sщ?7-~s��9��0o�65NYf��^E�~������8 �uxl��#~��j���@eT��v��;��Ft� ��pF�Ǹ��/�g��T��0O����LKf�l�S*	�kaݮ��(%Xd�v���\Gf�ȭ�.3�n�6|����wg�\�Y~���u�/ΐ""�Z�����J��Y�co	��o�r,jX!��l��UMe� �5El�JY��r�m���j\�s�$�"+��ډ\��#�wz�ڛ�����`��bg����P�x���ZP���x����< ��洭���T��&��P4u|fFN�Ζ~�B��L�d�s����L̕��lj�s&�,�u�����8�X"a)�
���)��a�42]����6�q��Ǔ)We�*N�S�/�	cފH	Q��Z+�v���ׂPn�05��KEq�5�*��8����uu��>�q��;�uI� d$!�K@わ��s�o\�l�K=r^�1)K��Ԑ�H	���Q~��5�9�|\t�f"�S������Tq �<�`i�.ц��n���w그�g,=A�V5��<�]�3�;n��5�� _B��Sܺ���E�z�a�\76��T�o�|�J�E3���`\\ztP�8�*�>�n�	���d����?Fs�Uw��#R�vs$�I~*���Bqp,<0W-op�=��g��#:����B����٫���M,h��K*����ٶ����-D�N4�Z��
��EOg.l�Ңh*m����|�TW�<i�6S�*���|����n5��ӕ#_�8�f��J͑���ꦌ-�V�i��Z"��/<hm�p.Yef�P�a��A�;�0��
זD�J����VI&m�ciiچ�P��k���}�=S������Kj_�hO�P[�l��jj�1��O+��}=s����]��-�L�ɢ��(J�2�M/%k���_ʯ�����`�{�ٽ��F���jC_���t�_ˋ-ϕQr��u����:J��+Ux��{�T8���тgoV��J��7\%�ݷ�.qk��^�r��<�;	I��qY�K�y���"o�s5Z�t/0{a�ӍNti2��S�nz;Y�8�jl㱰�Ku�<nQ��Dvt����#3�~�ݟ$��Ý$_ϊ!�p�
�Ot�L9\x�z]*	R�wZG�ˉ/ĆW��&�F�v��T���y��a����K6a`�X_�;��Ll�'�GN���������{�Y�`b_[0�ձ���Kδ�9`�`�Z�#DtJ�D��)����&p�9u3eo�P����"x�-�Y�f��X|BO<Ҏ�)�q�H}��π�30yDdL��r��tW�`�p�\�zvѱ��w+|�ŷEL0��8�t�E��H1E��zw'u14��0M��M��,� �L\�'�f-��^�y�륙�vҘ!;�b5s5?k�a#��Å�M�U���� ��q��ze�&j=;^�y��Zt��\�2e� ��
���u����?���sS �F� �Gvx�eߙ�����3���t�{�j�O�@:�'E�r�94?3���-;��5j8H���p�ܒr��ŧR�4ޝ=-vB��c�������vm�ڱ�j)�ף�ha�2ww}��>�7���{��S�r�%@o�{�ldȦ��h&�V�nN�l����!����V�١��Z����of�}��A��B᦯$Lj��m"���H����1��Z���6��Q�n��O�Kk'��gǝVhw<��ֺD��C`[Qm#e�ʣlo����/T����&���S��g|[y� �f���󅧮!�鵰��#G�T�B�)G^�_�ޙ��@�܏M\�w]��_�������C��}���;�y]E�ŗD�	���-�67r�M��W[eL�Z�8VAD�a����0T���a$-�p׸3q�M�IϹ^CR�R�K��j]d�f����b�{i4���$;�0A�~-1�<zH���+�ص�ip(";<�7����vG]�ݬ��wQ�b��n]��3ȹ,^�o��ð�������*��/���~G׃(�z4��{�t�!e����6T
��q�]}ZD�MV��0x-=��������8��7	{�wcM��?Z���<+#k�v�4'�6Ί�5n�*pL�
����E]���/��|j*��9����AQ�V��(�G�;�ƛNK	�6�T��Q��C��q�]�o&Օ�pr*Zy$4]g�ڔd�~���e\�5׻C�8���D�'&�nx���/5Z��b�ȣNڽ'j�v�v[�=s-�V-c\�`����d����1:N�`>��ox0`=��+��,��o�'�!��Ɇe���L5�v&B���� �L�(} �D��U�N�wW�ؑ���j��JМ�"n�Gg�7����:���*�0BW�su����O1O��{,��U��_��N)�1�0K�ÜD|a�#�P�s���D����?q��{�`�=箦mB^m"�+����W�P���+��|�*fW�)j�]e���՜=9���v�� ��N�w�����o,0CH���i�u�T��bk
�-��QWS�j⒇׹�['V�UP��^���;g�1�xAi��﷯"��`�	3qc��ﲖ�	�o��dxT�n�U���{���b�f��8g�h����3>]{�6sQ3x�Wb�O��f���1�q�ܴ8HO���#��@�b�,�ܼn��J���`�'2w�l]�l�����]��E��%�:�9H��g�l��?Z���t|�Vv���a��+Q��mayn����y�/���tt65���]R��OB--�-��������e�?�rz{=Kp���	��>���D��i��دxwE݃�0������8L�0�HG&���3�h;��ё��-K_3�Z�R(oR��*A���|����#v�;���.�0J�B�*��.Ĭ������^�x ��� 
����it��[S��z�O@�Ѷ��:�3��5U"E(f��4�"͍^|�F7MW*�K���I��ģ�dy�{;��u �;��T��G��-�s�>DA����0n����|R�V}�c}|-ؔ�p�ｷ�
Z����*���w�|���P�^��D���U���'�3�n�P�����ݖ~�f5���FCϝ����O#�f
�}k�;Ak����
v�v��L�Al[�È0Ȗl)�\;6Y���L��Jn�O�sg]>1;�a�yՋ��z_�n����U�$�y�P����򁩫<�@��.���%�?��S	���̒��h�xg��o8���G�L(�`0�u\�|Ĩ�|�X�w�^�m��q����0~Κ�����6�9�)� ���Z<8��j�OU�����J�=)evƖ�T��`�p�]ts�rvJ���A��Y��+�0IL0j�$�H��]�U�w��L��^&��z�%�VEŀ�D��orU�}Juz� �m���+b:0h�� ��mlD@�Bw2�dA��ˍ������"t�9��c�u�3)�~ʓ����܁ &�v�}��z�p��!�w���lo��Ti�h���B�|�̗����1�sg����]��>�}���l�r5\��O���Z�v��1^x��+}l�}[�P�U��R�S�b]��Z���<,M0�]ݚ���o^Tח�Z�LCC�GgP�&���b���=����.�%���X��u�α�����y��9��e�w|z���->�'j��{\���sW��qe tv\���@��t�}]7v+.��3q�H��.U��LJ��4�#B�42v�op��=�z<�?�`WƁ�՜���?R2�Q;/T��C�(�u��*+�M����RؠlΘ ���ق��n�5�9��D��=~��a�]oE�
�� jj(�Sc���v��`W���Zo-�o��=�ǈ�`vء:��{���Hj9Ô��-xJ��N7z=6��j�}5�t�@�sY��Wʰ��:iڷ�g�� �ؠ�k���s�.�6�pFoj�bZ��}��5�D�5]:`������{E�=-������TQ�
r>w���C%)u�z���˥:㦁z�9����x���|;d�����w#�O��]����}Gs;�SL- I�Ka�%lT���x�Oa�4}���������X�t{j����qQ6���:�ĝ�m��T��i��p]�TzW������S{paܓ!�9��(�y��F�Bq׼��ŵ���Zwb ���r�E�q�'�Qs+4�Ub�ط2��cF��+w�m��Ɍ����v��ץf�R�&��"nM����v�o!�^w������k�=�8��W�r�5 ��zr�8��Ğ��m��]oX��yg7u(�^T��
����Y��'[�4,�E�if�N�akM� T��2eF��\y�cS��ݗ��0l��^�gNBT�0�7��۬��ñmF4l�%����{�#tii|��n�l<q
����îb��b�Fu�ر�mS\�/���3���uL�S:�G�T�-J�. q4����pA۬�|g�-7}�f���*ݒzM��r��W;�Y�XSq�6��gNm�#eF6�7���k� ����.����8��_Ky��[PŹ�a��k�{�G��قt9*
�ͥ��75���B��5{�����v-�}�
�y�O��#ݧ{�	��+zdx����K�l�i�o�;��\�;��?M��v��˼�H�_*a�o�kx�>�=<{��.ŧ���ov:o� �����gn���dٵ��m��1wD�� WL��)j���r�H��
�2Ws��g@�B�T� w�m+�ێ�]��$���Θ�Τ���R�}˻��@ˣ�s�S�k�P9I�[��3�ؾ;ۗ�E⇇��s�����ogC�o������$�R�(��A����]$���N�aҹeAApH
xx{>���쬈*�"��CZF�N��a�	�fE*"�.P��g����E2�e�d���e
��m:vb�Ӫ%�q�����R��s�ӔG
ɪ'#5l��vV�ZpitVˉ�h�J��Vd��Z�ĥ�9T%r̵�T'
t ��"�5N�
�������L�ĺȨ("�sIs�z	IR$�QT�ӧH��U6�p����jӑĒ�͔EAd$�(L�!�X,��Aq �(���$��+�
�ad&�L�*�
�^���dQB�t]��0��fˋ!.
�
d�!Y��$r�}�ғ}b���D]��8�/�H�\V6 �5�k��D�,*}{
�)E�6<�<�>$#�M� ��6� ��0`=�W�fT�rU���Ɗ/�d	%�L�q���N��)�	U�����[�7s<�D/b�������Q}ô�f�� Q�PGCe�P�� �:$������3Yd����L�N��u�!]�2F��D��JS]�ذ�++�)ZN?����9_��Z*�f��#�r1�6&T]^uK!�{*-E�H��U-�,�$�51�}lޜ�>#�4�fN�cV����+�ÞZ�B"~�,__�#�ۘ׭ԅ��ઋ���u��zzAJ����};ӹ׵]�2!EU-�
�-?��{n��6Ϸ"�x��P� QM��GPN7J�@�1qF��:&��n�/aŗBY�^��0O�xi쇆Zv)�=��Z�vBSg�v6M>�ۚ������g/nuIQFZ�����Ki�,$!�:<���s��<#&^}j��U���[���J�e���y-�땂c�\f�/��q#]�N� ׂ���H�_y`L�׆�<Eeg��xh�g��,�נk
ka��.�WZ��i����rۥ�H�u��)Ǵ��=B�x窎F�j<`\i�m��<�A~�nāֈw<���*_�7[��Qғ�'n��y�-f!3�s�������x�g@O��_���x�m���8�x���l�i��>n���g)U��J.��WH\�3-��n�Ds��?Ͼ�0g�ٟgkJ�i,M˘����l�}8'�[r�K\��'�d�(��4	���]E�w4d��t�Qս�rY���4
��J����JU�#����7x��C��JdZ�X�EP��[z��z٬9��c�|W	{;8�O�\�*�b�(��Ǯ롙�v;�O�EAA��o
�e������ngUF�5)�<�e3�uyI��<��<=E2�/���y��N�"��O7�]��w&�Kh����Օ{����S+"X�cL����.=a����[���'HoD>�v�Q4�ncv֘��9Y�W=,���G��z��e<�m��Wd��Y"!� ��V���a:��_�'~����s�E���a�t&1Ӂ*.^4Ay�d�ϲ��eK#+�3FM.W\"7M��^����������3hsh��.!qͬ�S$txE$����f
��:$�z��=�YRkX����ګ\����x=�9H��������.��ϣ�3xwY�up��Yy/&��5SL!�>E��r^h�
�!��"���?q������+̻F��FmI�x&��2�hh��".p�
���u�5cz�?+e]����0�������g���4�uɢ1.^x���Yڽw۾rVpx�wqE�K��Ǡ��h��f�q�VV�B��|��S��W����ը�K���,�v4^nV�%��K(}�=��(�V���/�r}���
/Ϣƕ�zl�tO �?�!i-��M��WMN���¨�sSov3��N]�ݶ�`g_)�#:�$m�st��.�.K3��p�d�m���.6��9I߻�7������q(��vK�Nm������I� ���w���ߍ�xOp����Zo_?�ރ��-�
�>�wx9���<Q��}��|²6�㰴�=�Y��!�#Z}Ɓ)�=�LQ��^j��>k����D�2�,P�l������ؠ(?{[!`s�vW�����B���3[pu��+��]�7SO����Ҁ�������Qۺ�nZ�1ַ�@����#2b��Wܱ�r�%3U��r�v�S�)�00�.1�2��%�aC"��u��0X�ֺ���O�߱b��"i�X�$��"�J�/墲꼚�FЈ�R*جR,L]�E��Z�'m(=�J�װ��a0�}]�F�6&���o,0~i��V�����s���x���X$kcE���d92Ԗ�r�f_F<�7���T�3�/el�;א2��W'J �D���?��+�S�`�������.k0��"�:�� ZP���ʞ�6����{��7�`���>%F�Ȣ.���nr!��8���n�kfp�<]O%���k�8=6�#Ϛ]=�~n+���v�v�ʵ��kw�����:���ʁ���>��V��^�����kG��M!�b�d�ѓ� ����8g ���"0��{�h�����vM'��e�P�4]��i�>�zh�!dE�l�x��_y�A�b� ���؁��c��2S��Ecd��ES�]�r��Q�`0Vk�R��\pGm��o���ї@��c6��6��j��&ǆH�c��R�P8��I��GcX���d�!�T�X!��c���Q�����7f[�~��R�>fڗ�!���
�i ��X4�y���=F��T�Q���.{9��f-߬z8��Ax�R
󽃢��j	?7O��9�a!8��q�̺AaUR�zݨg�ʽL%�/Z`SkG��[��˗�o��H�&U��wIfC�;��P�Lk��ZVꢒ�;�Ҹ��	��6�ra��LKk�|Td<�� �S���)˖�^�h[�ƛ�Js�HtY
ۆn����{�0b4k���4��p��g/^YoB���y�Yِ}���^�>埳������ś��b��3g�s��q�9�7Ʋ]��b�}O�^~�QyW9ڻ�������/�� �ջ��xr��z1�����Z��5���;���N�@b�R��I	��f��Jy"RT̠$5*r�X�L%N=�7�j"�w.b��\&c��ڕ�͌⬳��o	;�N�oeH"6�px�q�Q��}��1��z������$�QAiJ�ִVB���irPna���Q�OW�P*�%��>���eKk�[�	
��>��HJ�Cb�9�1jtd�{Tjx�U���N�-h������(p�Ma�5�Y���q���j!<!�9ڙ���=�.��<���Χ��&�i
ظ���G���M�}'�w�G6�F�SˣC����!����c���oP9�8i�K�Iq`�g�����|=l���?_s��܌ᰠҡ�z���Qn�zs�� ���Nd�$�~2(�(".���
�4@H��@��ٞ�$}�u����s8���ñ�>����%�BR��;�ii�0$��
��:�1(f��]�lo�u��w�*�S
Wm�p�ώ�"��y�Al	e>IJjj}�֟zr�k��df��in�7O�ܕ��C��b��#����C[S�^�R/�Ŗ�ʨ�O��!����d��6mCι�7r��\�r�x��
�
�+�BTn�p��o�`(Z�Ï"����a����ߧ�DC��y-�
�V�K�,K��X�$�_qe��VA�����1�Mg֦Z�﮻7���w�H0!�����;�}�2A�٣��R2�)�*e��!L�z�K2]�MԵ6d��m��຅-'����ץc�ֽ���������@7��[�j�����C~܉`��a��G4�A�͚o�7���u��d.0wS�n�`��.o�j�{e�
4�Z�_ybC��8�z��X���ܣG�ޠ:�W/�9���h�]Kǉ�5Xr�y�`�-A������m����j���'uk�qx.�D��Ȣ:�;)s��� G<�_m��mm��.�l��1=3�sۛ/|��ͬ ��W,x�Vӫ�)E)�/0��R㜻�s��Ȟ!inB�*����������p���u�w�7yQY0q�1/	�E4�c��z��}Cv���Y�g�u�t_O@�p��G���	��o9�,°��vq��Z"�q�F���0���;�)��	5�B��n ��%��_E�{��/'c�Q�^�S<ğ�8�Y��*�~��ݮ���7˴�HE���]]�֫�r^�~��A��E��]��eX�أ���P��77��n�@e��=���&�O��/��y�,_���=�Ý��"ʠ᦯"s��F�E�Ӟ�R8p�U�4u�����}rkp��D���l�üKy���fU�ٚߌ#��`�Mx�CN�~��`�D-��nWCEz�D�s�<�Ef$��luL��?`2��H·B�A�G�Z���4�&:�}�-*�ݷ{��N/h7ع���uv\�ƪH���M�c)���0�4T3��򀌑�4<ai���Cۭ2u�ef�s�*��Ax�p�/��&��oI�+��5Q������W��Ϟ�n���5��;'��>]2p���+R���E`j�����1�]̪ͳg��zS�>������_¥1"�ig�s�(A��/8�ᨐ�6�}i��|7	���WJY~��r�YU�H���_�a�Ƞ�ms�?q����*���D-���qU��t��K�=����ᕙڊF�,gݲ�PK��W�|�Tx��O��1`�;Js.��t���f�����	���MuBF)(���%�B.K3平l���սeI�L4CD�HG+͏ Z(�4v{��*��3L�_C����#�jAƝ4Aq�0i�Z3�^]5�d�g
3 ����y�M�-񔍘����R����8�-5���5z�"|���U��{���\$�<��$_�	�d@z+��u(O������)�
3�Ő��=gg����[�vAd���ī�ez��Q����N� �L���(�\�2EP͂��q���4�gs9(ʚW�ߥ�������_e�ye�^�i;���Wϒ�,n��+7Ļ�J�^O0�#[����݉�ʯ뭩�=��~�/rE���!��#Ճ�ڽ�{䳬�]u٩�h��T��n�C�w��ٷ?��0��a����!��~
�fXd��;�v�,x߰�.���hy��a�e�?z�<<V�����8�T]�ba����ނ���@\���"�l��VG�U��-��x*lV)69�7f���UNZ֜~�+�/Xi���7i�5��<�X`���,ei������My;�g�5i�H�0�zB~���s/�=QsM>Ԡ,5��A��-^~el�#z��!��n2Ghc�o79<bPw��*9����/i�v��q�g������nb�7^9��qm��ٝŪ�w���^�='&���}���Dp7!��Cn=����6 �В�{�=��a�q��27���_^Ӥ�UȻ8�Eі�r
�)s�dm��i�(����pk2i�2�b+�R�q2xd��/,�"�q�H�j�ќ8��@�f��`���Ҏ��S-H�=�5qW{J�Hk�gk�S����)�j6Կ}Fx�qR2� F�H�o�}�3��b�������F��zՅ��AX���W����z3��7-~s��� �4cg8�,U&ouՆ�ݽx6�;yu�0�į�
�����gTϵ?_���+s��V�����A�.ﳞ�ƙ���C�N�Ӽ���ޭ��F���sQ�7uǄځxVt�q��u�x����HG%�hɽ}X�� ~~�=�NZ�ֻ���{g����������+Yᎁ��?���m�>2��˗���H�&U��Y���)�l�
���v/�L��|a����iO�>��i�
òLKb����x�@%.,��[�<��[^����]f�]>4yUC6O���p��i�~�_����nt���
���zj�lDZܽ���Pؼ��6宇a_ݒq�u�}�@��`����sC��59j��+ʗ5.i.V�b}پ��
ue�azڞϔ�ք��(-Jo����S��O�J�cЉ���n����;Ϥ#'���]/xWw@n��`���PHPb�4f,:2~��5=y������a�N��ͬV�mt�0���|����lX��1�JL�CUtȞ9�pd�ұ����&x�NgW%Y�.݁B�/�;�����V�y��~���K496b7>�!�{ Ds�I��O��l��څ�!���f�+��Iuc`I.�*0CS�z�������P���L,�oY����3#�+�tR.��Z�fE���Y6�qv�W~h��4�~��?�)ct�����Y���s��m�wS�-m'�%���A\U��曦�	����=8S�U
<f��(�T�bT��{�n�bچkC��v�f�KU��үu�2(��Ԣ2�<����{�q��
sG%ូ��l�$i���(����nd#BtF��%f?U?z{v0���U�4���ǝD�<2F��D��BR����f�@�LQ�I�^8�3��v\1�.^��Ҍhrښ_m�8C ۅ���)<����%���51�}f�5.�s��u���߳��,A������o\GWSת`4�ԋ�qe��UE�~�/O@��G��WL�����y�{f��(���L��x:l�dƆ���*qk����).u9|�;a�}�����7���c��������.�=p����*?B��د��ݿN4�{|4%�;F��jV��e^����d�tϑ�F�<�1�c��0;��OBh�����&��N��^O-�G}؇m�Qm^����ӕ��V�m��]��v�;?k ���sC������=���[�QE�`ڼ�LLYC%�ϖt�T��q|e���=;]/:���,l[t�����R�Ҷt�=�V�!�K�N:&9���dr}������z%��rh�n������pwo��˽���o��;��g��O����~3�ؽ���k��#��[�E�93%q
;�G�߈����eb�Yg/3�;���U����p�F��t�����ҥXqP��Ud���!RfI������el��o/���P�i9�2�wk�:����t8w�l�'\Mq���:��.���ѢÏxJW=��}���k��c��ܲ�C�������d�"��AcÜ
�a���h���[�?��-�9r����/m2����:��Yw���
ν���6c�8�l�s�-d�mv>�\S8�����{nEK�u`>����}�ޑ��P=X^O�-����Y�=�4�,,�Z9W���v�d�n�
#l0����r��x��iɻ�u�	\1���p*�������"٢�<�j3b鐶.��l�C^���z�^id�L�|O��`7Û��1�z�X!��'zR	�y�����xh����X�����/w1+���9ݝ��V'4�����=F�C����B���b��=���'��7��[�%�`���UɌhGro@3$��goӳ� ��%gx�U�Y,gh���IŸm�6�,������N��u+�v-�C�n�2���H�6�]�yqδ�6f�i/�_M�r6��NOkC۾��H�ʣ��q�5/$�
���j!r�{�>�0tY���z�s]~��\��v(}��0��0%����,�=��]����=���A��x�T����a]�[Mβ��2���%t4�l���|'>�c�[�jk�ݺ���n�_�%k����*fa|n���{��a��g����`H�����޴�#�-���[�NU9�j_��x��ݒ�����(ޏ�Ȯp�I���yo��%A��z������z[�t�,��j��t�&���:���`��#"�感J3gr����+>V�[�����ީ���aa�N#���:��H�E0F�������3�����R��,^v�$��=�K*'�ځ-��zd�B�M
,7F�-�𦵥\����d��t;.��)&͉u��CzR��S�B��1�)�}=9�}wm�oػޘx���^r�s�JQ�A���r��"����VB�������Wҹ��̋�с�����짷U�or�:ʭ8{rK�YR·�ۻ��#;V��v�D��t��ؙ7���<=�[�W������=�𐜸���<҅��Ss,^�V����dNr1<�s�0��uz��D���<I�[b^9eH'N�v�Z��i-���i�9��%a��@�]yz�;�?����~��>����<|Ǽ�����݉����>��V���԰���u������P����x�֫P�Q=}g2�쫔��NW>K{�NJZ)��q�u��5T��pI����"�#L��������jݼ��JЯB�Wɣ����R!v6� ������X��s���x��p��h�{'�k	�~�zS��E������@�-Z�	����AO�E�%v�����@Jΐ!�Qh2��\��1}���=��qhg(���jM*�2���!�Ӱ�
b�� �I8�TI�h����{=����Sat���|{�#;i�Q8�$DȢ��'�3�͉�i���e@\��ӹ*0�¨)�F]�˕t���.��aT�NPS5���NY��
�
"��*�9�+���Zl*�J��;'��N���i
����.S.;������W9�r*%
�uz��\����EUW�ERa�J��.'.Wa�C�+�L�G�e	U�L(��k.ʸ���y��8PW��T(*��w8��EsKa���:d(� Ԩ���Q�"R	�ju.2+E���\����\�[59Ts�\���f��\�&h'3*�V������¢�"��y:����'c�e�	�9��p�hꬻ ηf�v�o��N�;�Mj�b�k\��#;�RWy�໩���u���t{�NTO%�Q"4���Qu9~2Ƌ|c������������FW���r)W�����������w����ʹKOհRX<���������G�x�g���x���SU���}\������� ���$�o!�A�s��qv
G��u��~}�osW����1�K!��r��yKV:�}�V6��8+չ�=��v�l��>?q	��Z�k�c�U�b����a��S鎖!��T\�5b�d���_��r#:�V��ь�O�Ub뢱�!�l^�{�;5W�"�n[FӦ��u�$h��*�]B�ů7��x8<]ܣ���?z!���e��-�m^r�"<�)�����WP�ݸurf��;�k�xc=�x�DR�\	�zp�|d���#�-ÄD��-4x�AIh\5�3�&5��s'����zq%��P���ՉVCR���i��j�<p�d��������mҰMb�,�hȜ����kZy6�ӄǥ�'��}7�Ym��n�"֚<�H��֨Zz����3�Q�~�������l=�dՁM�����f�n�s��8��&&k1![jӣ9�v�3{�4��*�v�՛�`h�g�z��)˅�e��慏U�raD�fc��͂������U��^n�G��Z�x�x�9ϣn��Ǳ�W�WA=�H���g��@ ��Y�����*�����H*�#�bϕZ��&T1��;�;�S�N����o�}
����l���-b?�J�b�P��C�ǏG��>uo�;����:Jr0[��;a��L;��{qx���TB�1��)�<���í@86��L3,���{^}���aC����}!<�ڏ4�iq������S�%Z�s<�#C�]���3$Uxf�m��36�v<N9>��l�/U�����BWs��XݤK8�N9�G�=����Q9:��������hXٽ���ސ/��ON����_�Ed>�3P��"<���ٶ��(�ʫ�=��a�Ww`sr�Өؙz�M^�u�s ]���d%p-#�@��NAu�-Z���"~���l��y�׸��� ��S��֛5�{��d9�g<��x͋{�el�ї�z�/�(l�>�9���{���@�? o.n��ڽb�È��3���T#&`�1n<���U� �mѼ�Ҳ�ww�&X�/��ޜ�3Qpbc~Ah�C�h-�m��o�]�\�z��1���7j��v�����Ƌ�5�[��_!�i�]D���aR���RnpY�Ǣ�}�#|��-Ά,��������m�W��Q�W�����g
�,1��F�Y��D+xX��i���bq�w	��iXq��z�����6>��*���p<�4����#0V߼q�����d��@�l���ٖ���U@XM;��>��s�p{�?[wm�`7y�*�k�)IJa'^��5P�����]��&�^y4/���K0�z
	�+�/a�{)r�Ƕ�QL5C�-�Q�C�5~T��3"6rzԋ�#�p��٫�n����51�U��8�Xp�[��-.���\�U�z�	 ��O5f4��2lj��J��4X�AR���K��¶8�6\���-ZF`	2�H�]�온�s��CGb�g���uIB(�*����F�/������0��٦�k��!�} �Q��ok߫8S.�ܸ���̥P���
�F�����s�΀��s	�>�_����ǴB�����^x�ǈ#�����c��;�+��Oܮ�
츄~U�&�8�q6���>���n����u�%K���F툍�SSܦ��$�QAi��~����:�Gܚ^�
wj6X�#~{�ć��-ȿ���nse$ 7Fd��}��K9���]%��ςϻhm|&Ao�ﮕ|���ݬ������Ƒ\
+jh��l�۷�H� �_)�a/|.�Ӗ���h���A���K���נ��oXO�H햲g��V�51a-�Ye�|�26!Y8-�U���k���x$A�����a�x���hz����eͧ��\/�l-��M��"�O����? `_6���=��V9��O\p����!�Q&r���IIq�WG�0��R��=j��cS��ʊ��=$��~����3cT)�|a��|p:ɖ������{�y�f#N�5wO�筈5g�܇�1`��א׈�m;�94��f��P+����E������f)�khqܳ�Y�p��ֈMt7�M4�%�.�a=�vz��x6(�.N.=aႽ;[�E�y�˵��D�H��+�=t��#�tK*�%)���ٶ֖(ߤ�9��f|�D��/3uh�![Ŗm���
v�(27#��^H��R��j?��}]�<��=�[۫:��9��8N�M�4>������G�eJG��y �V�Zg���tJ�|D�I8{.��;�꠳�f�� W���P�E���}}N ��E���d^��������`�1Ǿdj��l%$kqc��Y�K�O}9o�tL!º��7�5�i֌�S��v��0��7"�5+��b@�9��tϑ�F�rZ��(���ߏrD���c_=�[K��j���hp�c���ii2�/�[�ǅ,"��|�'��k���^��hy����<��d3�Ԭ���Y�H2�u�I�Z�A�:?@f�'�W7���3N���[��m�z�G���6d�-��<�	=������x�3_ǁv3{�d�ٹ�E��Vl�,���]�@}_�G�W.W�cotF����.5WY���ە�&���Aq;Y3�6�G�k�K�L�����c��;fB5
t��F74�w|��>{<������r��{d9m�$��M����>姃1���X��a
�l]Nǔ���Ξ�D��inB�*��Ňź*��b�/��������X�l��$?��X��c������[t6]�GM��"�Jʘ��8��g��cΰ�<w�ե�d?utȰ�V5\����"!?�����?�__lyT���(?)Q��mY���[��&O����0S�� ����;���y4�$�y� �<!�r��^W7�6���lƲ����������SbA�LC��(2�zc���d�{ [04�48�ѧv5>��0����Du]�@FJ�i�x�!��^��=�Ý���t.MfĐ�d��eN��fk�ٻ���d������n68<".Zi��^�l��b�)�-4Ax.��qX4��-�Mvm��e엧;>��/����Fd]70F��Q��z�79���-{=3g�ڳ�`�C��sWU�x����=�F����]��pE� ���o��:��3ݗ�s�׋���*��	-�[ޱ�\�!"�QY�Tɰv�1�rLf𰡖+�9a_wE�����r����?;�w�]n�m�hҔ�G!OPW_d7�mCe�;H���[m쿨t�����ƾ�!��vD|��?��*�&�?��l�����eKH��!	oH���_�7E�Fp�+�b�<G)�S�Gl��E�9�䰣w=u�m�Ϲ^CR��ϢƮ�ӄ�,�4�XL�en�WC�q�M��gs�n��/�}=� �Z\B�����,���P�kM@�®�#�g���a(mWF���a��]��Xؼ��V*�ƹ?q�ҕ傴V�F$�@/kO���8�}��a�Hw�u�_{���0b8l�0<��qM�6`kd�z�ǀ:���z�N'ING��n�:�z��Sf�.v�Dڙ!{6�sJ4	P9�4?����5��L3,��<�[�(
�Aݢkf���@�){j*o���t�_�+zAc��O���&��X��d���ݵuqEB���t�RڹLUja*�^�	]�_�Ed#�2%N�L���D�:����xT�⼡�KV�U�v.t�I��5�ݻ���^�4{�$%96j�-�=2��]������WΪf�ٟ�)׵_�}�W�,���؞���[�Uļ�9��pqY]��t�e�u��Ǔ��v ���;�����x��W�x,P��,hIĎD��}˃���ܑ{�`�A,B]�F�j-�q��-�(�mf:Վ�Ih�	;�j�57�a�q�m��F�W�2�����1w)�z�M[����t�x b����4��yZeǙ���^��PB�9����ָ�s�a�\�" =��q�8Ѻ"��Rp�ﯟ�2�R��L�^E׵��Q�����c�"wh�^�yr�c��魢�?5���أ*������gֽ^郱����8Y1+Y��	�bԻK�f|��d��95�LPa=4yl9	���ݢ�kmҁ'�24yj����u`����[�:�/����R*��fF��Ϩ�. �ǜ���]$�P������פ8Q�b0v+�C"^K��W����a��p�g�.�߲��7�0M���bʢ�,��"�R��$q�މݖ�llڕ ����^�a�����Q�;A�!��u�Tw�7�s�mh僬�?~|���x���AX�R	���).z87J�p����s��X�;2�j��!��"_����?�`�������<���G��ZF`�*��VM�V�M�;�}4��f���ѨC�R7L�[��<h���4:�:0e�r�6y��R�3����a�7D����?Rk�F=�U�PA�W#N��x�ZL�Z����@|�Z&��U���8���ۖv����a��b�i�E"wk�Nv�oj���o���.�p :*b���:*�qs�������i|�Dn*���k뼸u*�[9����_^ݏ��_��]@���9~�m~��7�0��5���)6����N��d.�tØO��������U����Y���O�}v���g�`�/��q�J����+��e�"�L%" �8*ƚ́&�G�dR%��z�'⃘`�8җdw1�6`ۅ�k��8I�PZBT~��VB��*a?��Lz/��TSdc6_��V��=��@�":)��{�u�ʛ`��ptAАp�{�3�2""*+�m]�f�����t��ڢ����:hny���4����l��w��Q�gZ���J��#tF�X8�v����q �<�i�.���h>�4������&cѦv�)���ÁVMFT���8�7-�c��3���^ ȼ�FE���v� �)��ƅ�G��K��1�V�l�-�p8���~���q�	[��sO� /�W�$d��F�ɰ�qr�%�X]��T3�+ހ��"�{D������A����Upܶ��w�)MT�m���0�w�V�+ck�UU�oo�_��=D��z�a��6��ׄR7���[YH	)MM��@�_�f/�d�.g��Y6��l�;8O[���n ���i���>CTh�_9����f��iV?�q75�㼞p�U��N �<��E�4;�ɻ�Ln��9xfGFU���s�pFgc~��~����y	d���#�>�(�$=�v۱���۲�0����{�v��L�o,>�j[�m����Y���C6H����p���l�H�0�+͙�T��Y7�J�鎳�܎���|��G�=0pA���t��Ce��֞5ء������fI+K)݃T����+l��޴�l�wĚϗD�x�v<��{����|�����~^��X�:~��z=�G>�=�B���c��RCu�%�$:8�z��k�y����WT�j��{�E�Dmf(LLԅ�B���S�WqnTxkV�o_�&�<~�ɘ� ��e����`�1���H��p���Ll�5:{\�d:w���ϸ�k�|����w�Y]p���t���k�`�s�n<� ,��l���!O[x�>��q�|Nz.��7w��q�7�ݗt��m�D:��'GG�Fi��b����x_ݛ�<c��EW���C�V�c�$��	�ד��v>C���Z�4�=y�՚���6}5�ov�z�c��M���2���4�dud�q#�3�9���l���5�k]��y���;د���M��?��e�8�xTl��Yٷ���ή�̤+5��=`���,�3
kS��ݣѺ-P�":�/Ypɚq�7��mk��^ �L��p޽�w��w;tS=�>2�j<f�|��/m�׎jPv����{9��ǐM�ŧ��.�侨˾�dz���X')��fc�U��J"�����r+x+)�!5����7�q.&�"���U�y�f����l8�ꡟϢ=j�H{[�x?bV�վ��mUZ�"�t]EU������0�%X��M�u!�"������g$��KX$�eP�^
�;�f�*�5y��d�N6�۸.�HT��~�,����>V�I�{��ǫ���6���]{цU�a�A����=���'�I�������!��W���E����<�6��덍��c��ɓV�8��9I.u�({o�V��Y�#��!y�m�{��-�P�5u��H�FO�|�j-@����u�3�(���ϽKu;��D�
}D�i�jجv��Y�bǖ���Q7����]�r-�վ9�O�vw*��Oa=+]��o����2������k5��v:[�sS�:aU�h�&u�]k6��ƨ��"�|YT����Hx��3�n��#ҡ
կ��c։N�9#Hm��;?I�ls�2�����e���a&1�Uc��8����Э�����S�F�䇳H���8�mY��.i�/�Ӳ�ڹ��4�����eb9����lS�%�w�.���D�ϭ��V����ۏcђ�cFq;T�
�X&F[9L��zёɻ��q��k41��}�(~��y��CB�Tv�8�\[�1�Y8yc�u�b�n�Y�ŚYn�'rҘn�k��4�'%vd��:��{F���d�`�z�น2�{f�7�y�R#۾E�*I��_�LM�BK���U�Mw�G��<����ز��%Y��/KḢ��-%��yk��	]CA\��e2���؂8`{1S��JV��qԑ�Qu]֔f\�Op�;dɆY�+���
���딻}�n��Ŏ�x���YK#��P)s�K��U�,~>�P��������ʬPBEP\�q�9�Y�����q�g��~d�;���䰶@��q����a����Ԣp,�}:���j��/��(�!��p�k���n��vZ혌��Y=�I���͋<0>C��5k�h�=�Z�H�����z�|A��|ٷ�#G�
o�u}���3ԇ~sq-�g���{��y�k���6����r)Q̡:G� ��ј]���7HPM�tq�騹�k7zP6�1���1�i����!~������ؾ~��te�t2��t��8���{g��n�}�V!X)B���nWt�V;����ߕ�j�3��\�ۺϣ'J��~�]�.�F4����]�b-ΖSˎ^��uͷxaIV��;*ЉԈ�Z�dB�gr�A�������WU,�ض{�7R��kf�ɵ5MK�6���c�5��RL,�CS~������$��a�n�@�MWBVV�Qvi����lu\]�ç���	:�˜��0B����"4�F�̬X��W&�Nh�M�Ȼ6ӧ����u��N�C˔0b��շr�"Q��I]���a���)�Y[/n7g �7��$���|�8���)ٓ��D<�׬�=P����L*h�Ny���!��ޕ����u��Z�kh�uU]�y���-7�=��$�� �,�}��,�%��aK���U�T,m�uũ&�}|�x���{����'Q�<Fɒ�_lYyN�6���<ߔ78���TlG�ҙ��i�#�bS��+;�]��Ċ"��b�XM���b�*Y��GP��RFj��#U��v��6��Ȼژb��\ ��9[޵V'���;�Xq�ǻd�;��g-dq�Gjɮ���..[p�R��neҕ�A�[���e&)���ҧ7N�])0#��}S���m*����ewC�N���mĲ�j��֋��S���{������{I!����;�M��:�srS�/�wm�ݾ�#� �EI�A �J���r��Y�IA�Я���9E�ʸ"�gۧ�<>����S�iT\e���(��J��E0��<��*�CK"x�/0�ǳ���{=�����*��DQT\>2"�6$D")�tIQ&P]��(����Tt��U��\�#��n@US�$��*�����Qs�n������H��
��(�5.��@PW8��f*|t��(����J�!'��T���"�ˇ>P������UW��i˕�U�2������.wt=aQ��Nr�:����"�3���>8�y;�s�\wv��EkN�k,".��Y��NRg�/#��1��ܜ�A�QQ{����|e�!�$%��{�q�ȫ����;���q��������,��ATr�S�.p�M�U��ϪEN{�1�(�x㔈��B��g�wRȌDx�����꼣zq��9���v�_+a	�=�"�$�Dp��w�H��!�QE��u�!�5&Ec�;�L��� 眈.QBIW�%D��ph|�h<�E>�~��vro{�CH�o�꺆�y��T��ڒ��k��A��~���d��{��Ŕ�������O7��Dk�Z�WC�������Hk����;�B�7�y����㯱W<���B<�}\Z\�+����V�Vqs6�k�@X!)��@�j��:��:U�؛έ��N�g��d.GP^�e+B��U��j�W�!�+�|�[}{��-�I����';�����'� �A��E �}FW�S���\�G*Oyw��-�t.�˳��;V��bl��P���m�Y���'/�:r�]8l�5�\`O{>��˿�J�^��߿~������7x���df۹6�Gu�%QIm=�M�5\%�*2�P=4�$bč��}�x���z_7l��}봔�\�x.��޼�*�Ȑ���C�M�0�;uF�v�����1�~�;��F:�!.l�m�;�`o�]���P�᛻ZLsX�<�3z��w<��U8=,�+ḝ��o!So>���O��θ�/f*ｷU�sMݯ���6�6�����oV7|h�pt
��e��	_��^S���}y۹�0��v(�ϻXy�l?��ިm�`��tpA����v�O#�7fne��u��I[�����)4ɣ;�M�m�;�r���}W*t�x��ܟ��tI/L�V��Uj�$��ᣁ����XW���N�X�r�z9��G[~��D�Z�NDۃ�7׽FͿy�s��Å���<��-4�yͬ{Z��]�:�`�9��g-v�"�m��v�;�]��;�O��>�a�{|��_���Wbߍ$�Epș�k��h����Տ9�C����	z��]�� �E�sPYy��u{8^��t�YX�$zƗ=}�p��?Y�,�5"࡬J2vk��gJ�{��u�
��o�s�?U�����0w腦y���T����"�}�z�׳}An��6��q�OZr�����N/g9�ptkژ���%��h]D�N�򩥋h��ѽ�btRl_͆�4G��ѫ%�ݽ���OբT�Tv���u%Cb�{���u��k�Q��!Ř�o<�t��O78$�<|]��eXq `�a��o0�}}���Ӧ����	�����E�NWS�/te���A�)����a�d=��8A���)&&��և�Y��V[�uہ�m�K��ơ�l�ޓk�F��2�Ix���B T���5oA��	�R�|p�pDy�}{;:,<�{%ξ�:�9}~2K�m��i�3k���Vh��o���&��.��2�n$`YX��*s��5>�WH�����~�x^���I�_R�K������*�9�Vl-bj��#tַOxXu{!���B��#XL�m�ճM"gs"J�UI��L�Fb���{+L?�nPT�X�i��	B��.��6�GW��������I⼩����q����цv��1�KclV�v;Н��4��x��W�ͫ���'���Qt�\��ų���vr<�S�2������i���u����si��$���P8ҳ�E��!�X}q��ism���Z��Ίa��s\�R��UZ�L�_�����;˪�z��o�=,�Zϩ�.�������y�a�K�׀�����\�*�篤c�4~E�$zƘ�Gk^)�[���Q�oo�
��5P��7�V��qd*O��z~��{�{�}A^Ĕ8z�q��ѱpز�4�Kq�w��}C�Q���{�->x�Y:zt���X �kz�u[��U�c7F�ho8.�6�N��el`�!�lZ��c٘�%������g]z}�R��R띒���®�����Ṽp
<�ݼ������*���z`N��5��*~��d�͝k�}ǭ��1\�x���Q��/�:�,U�h�c��C�4tX�j��/R����Z���سET�nJY�p������;-�>]�}�s�z�XUZ3�i�D]u����j�N^c]q~���aBX�HX	��YJF��i9�$<�����9UHp�{�ՂO{S�����cͰ��[�[-ur��Ӽ�l����ǉ��XZDV��7w)Da	tc�b
���AN�Mz2�ڛ�Lg��ݓ����ޯP�շ���w,<��5磌K
\%,(��v��d�	��;b*ڧsv����o����4S�0Kc�p�Ǳ�W��dEf]�̾8�7<�_��G���,Ҡ���q��d���aCc0V���UT^T+�V^3�r"�"v�6sE�J;����ʼ�
����Rz0Y�X�u�B�������x����������=ܧ����>97{�Q�]�D��T���jܛ��S^"+��7�z�����;C��fmゎ�룎�7����΁=�o���?L�p p�����D0Z�����u>s+�"Aoe�K�+Z=W0�]z�b��Q����ǩ�)�Z;N�gB��հ�NGll��n_Oy�Rf����۳\q$A_hoo�ѽu��V|`�����\
-�o��z\ײ7���G{�Oq��3`*P�@��i����B�)Oe�w>x��g����
�z�;77;�J���p���#y���4ϣS��������ۼGՒ�Z�E-<�n������-���y
�}�C�#�_�?mY;u��m�n>�A�iaAq����a��p�����V��*�H�~�9��ϻ�+߃�|t�;�1sNd}^����6�������Y��Ew��FW��#(Ǳ���������A壕	��v��`�C���rB��/��V�b=T���L�>Vc@�=m�9ձf�	Q(uR�s�������[`�")B�UN�T�cʐD�gwA��}aѕ{hw=���"�e��$�3ljhb��У��?�������	�h��V��&�׽C�+�o�G8M9 �m�,#'�L��?N?l�����߰��./f�v��Q˘ݎ=����B���p�Oi؜~��x�:���w�SG9�1�/�c˱I��"�,7;q1t��qp�ci;Ә�r�ڴ��"��=���2���}�
U����z�tC���zʆ|�7��W"��f���B+�/ݗq�=�b�V�/t0^�T�ث�;b��!v����j�����y�S'*�e�PC��xY���Q5�7�pf�plǂvC79_˭�����6���L�gv�T�W���]^f�^���H<����ފv���I�2�τu���j���{�Ν��vLέ�A��!=BXB6���ii���n����Q�;;z}$z����xW{��x�.�ۍ���,�6*�3׉c�r���f���<X������>�^0�W��n0>Cy�� ��=^�f�ِ�+�f�[S�w��z�2�>����~� �������â_rsus���8���w���BB�j���[ߕ5�)���w�r���+��+��ؕ�v��0��P��.�g���n��ΞU��;���r��bx ;�l�qt���A����9̎�i�;���/���]ZT�5�͓�:��}'�_kFT�Y��q���b�&���+��L1w�����\�6'��	�949Jc��73�d�����67���	���|��pE�6m����(!i�*1U����^��"	�os��/.��Dz�Th�F�*Oy����=�N�M��
�ktүN��p�;�H��{b����=邂���U6��iﺼ�g٘�B�[߂��DM�ധ��g6�cG5@�����q8:�0�^e�.��CރF6h�o)����e�l{9�����5�iw�Y�`m��Y����l�2��E߳|���W3»[U���?��}jW����2������C,��s�{���\)��[b�f��k	��_[dչi_2���~���$��wl{PǓ�#(,R�`�i�ބ(w�\m6��I��&j�iW��y�ۦ�+�^�L��Vw�q�C䯌W�vb ��z��@����D��^�Բ6կk◕��� 0�P�_2̩��O~��A���_a�6I�	5��S���c�#�f��P`̕�pC����4E����%j ����Mݷ7�|n>р>L.��Y��h-�
Gʳ7��:AnoI�fn���=f�C���_�Gϗ,��+k�md�N���E��G{��ټ2�;�mA�\�ta�{=:Z�ap/������}n�.���yTʝ]ETf,�;�	��J�[u����h���~�>�����u����V��~�O�I6'�'��侺����N�e�,'���u�]"G���eE;���-����G�5F��b�����Y
���zyw�)�z�����n#���gx�!�n2#�w�4t ������_c��zߗޒ���J#ٖ�ӏ����)��v8�w�THh��Q����6����}�;~��<��@+�*h-�7Bw�E-_Q�~�(s�
��.�GW69\�ZpS���ǝv��:��`op�G����@���o��/}:�au����RN�%�,���s۳������'B7�Q���yoۊ�I�F�W��2����a�6��S�����L�R���s[àO(O��I�:"���\�1�}����z�%8~m���YUI��fN��p��?7���[�̇�}y_:8L�ۈ�Gs��~*�X�.{W[�����{�-ʗ�ap	���!��D�u��P�������")w��I�
��٩[��Ldԯ2�7)���$Fvq38goޅ�r�̫.$py@`��g���H{Z5"y�D�ڇ�������V�'{�����w�Ƞ�����ō��?doE�
]&W|�z��yJ�~5��`�M��E�I;��e�f���1����7MF���.�`��=��ޖ�Λv��	��2�x��~�AԹ�c��]��<3��B�:z��n��V�y�l�r;c^�j���^@����j���(~�}�û�֑
���6J��=)<����C���͂�]O���IK�[[���ñ��z�6#W<�_���Fϧ��u�w�ۛ��ֈM�	n�q����m�����P7�Bj��o�[����R�G��ܿ�G���1����Qw�ڷ�u���C��4(�7��jʓ}qu;kG�w�DevU��ĺ|u��	
�)�-�_�*�FF��
#��;�|6�^m�d�'X�]�L��Vx�v�5"���0,��	C�"�������L���!���ڶ{{!�%Vڐc��|��h]V�R<ޝȅ'L�sՓRZ4%}�F[���/e�I��V�q�<��-��[�ʓ�.��F��ukjuD�k�ب��[�����*�h�lm�r?%hZAz�L��]7ֽ��ϧ�����.��d�� �JC�	��F�y,�_{؄���M� ���l�MX���ru����nqq>�ŗY���gǰv��lN�¨����7�ا�䆓����v���6ׇQ��`J������_ɢ٫���"��ϰ�o��Y��?�PvY�<����I��22�:�*��e�½�r	�����Z��������������U��r%��9�J�+Å�������"���y��>��?GSE.l�IL��YrQ��pС��D���C����[�5�>��avBs����B���V�O7{�ro����EW{��'٭l���;��CFP�o��^�h��i<�Zp�WM���H�|-]ui�K�a��4���d�适�AY��]c���� W�j��W��md��a�yc�e��?M�#ط��s�^��7�E;V?b;�4	����p�!ݺδݡVP\+�c����6J��ّ���!R�%=﹍��S��6�.�N��"�{���p-�k��zkr\.p���ײnO���n4����0��h�|���=��Mޒ��x�����7�V�S�وf��-����d��`������'�����:S�5���Řa|�)�ٺf������g�[Y�xd;�T�p��7�n�~�)�b�6�������*J�	��2�Wc����~ΧP��7�S`�ȭ�ob7��:���T��ܘ*�m�-+��vp��wBũ/k��Y�;2�D��`f>+��Q,��!��;�r]/�Y�{�&jU]x�9{ޤ-�g�9�'(2�:�[��x��i4�Y�;kQZ^�gL|T]�<�]��j�d/��E��+�$P(���v�,����V[gypn�1�IF���u�����Yγ�+7�$��mS���������#�U:��}�PgD\�����xs�������/��j�#����w�,m�Z6���W�[���Z���Ǳ]�6���ױ�G��o#+�ɔ�t��L;ӨXeg��+�[�w+<�� �S�rR�Wb9�ef�AƬGz6�fܡ�I×p�Э;`�S4�9�.w܄��C�T�Tn��m����k��W�s�}���#�x����;i���S����\�e�W��u� ��y)�A�����Y�H�gQ���!��ڥfGS������sf��oBܛJ]\��YRL��3I���)K��9�,Z��_Tn+d|�ЦhfK_5�1Y���� �v��@*��)-{�Dn��7�$%j�͍�KV��c�o�w�o�\H�~�����Q�c�l�88����n͇���Rwbj�4��q�DM�4��Ĺ����91�]��-�e�<�W��y��л c y����U�KW�*kS	��zD'0��O��g���d^ζ�>��&�,�hŗ�t��s��S	��A��w���NI�P���\�wќ�VBtW�ٷ��¤�{�w������I��1��L�<Z�=]hl��,)�9��e�H��}�;ͱ�O(�soC�XkD2R�L�4/h�`��oA��vJO��^�q��Q4\���}؏���_	�M���Z�v�^1�� &���z�z��O��/��/F�I���x� ^��l�W���3g*;�����6��a�F8m� |���ݎR�U�#{gJ\�+����*Vy��r�L��gzL�'wkD�r��6)ׯd�z�P+��W��ҫ�Y��<a�$�`�;��K�y'���o��k�uW�i��:�m�v�T[˕��Z.�M�Z&�φ��x��w^�Ptz=���{���ܕo�kQ�n5c���^I6T13	���ۉ���	 ��^ATU<��=bL��E�+���9ҧ3��<�e<�����"*rH�����Ï��=���O�y��"���5
{w2H�"�:�Nq
� ��;+����N�����g�؈��ZF �\�*rA%�CNʠ���*�@]4-4��P^Wp���A��\��Ur����-�y�(��*��� ��!���R�U=�
zv������s�䗨E�*�:Ȯ�]�Ӻ.��ʳ�Ȉ����
5�����r���C��\r��;��L��J�/"�����0��EQq�E�t��J���ʮeA�yo<BVt��Ι\9Pr�J�����Y]$9
�����p����E�p�:�]
�T�$�FPQsA+�N�.�Q�\��ۄ���_I�*�:ir�">G<*�9�UWH��,��w���,'q�H�.mܨ�t�~loE���F-c�Rù��7v��㷴	#g[�'d>;W\#,n��E��X����!}����uo���Iw,Ӊt�q�V�m�Ǚϸ���b�l�xWG�
|X�n�ͪ��Uwl��V@���/�*ΐaV�f�x^w��r�==��|�c!.|SH�gh$z����=^�Z8�kk�Ho?v�#a�z���~����E��E5�N߻����\B2A�{����ˍ4l��n�EwL��51��o�Q�滂���I�����ۣ��3K/٫.�C:�"}�	P��SO��|;�P��:
e��J�yK��>(ww�]�]���D���ϔZ�����%��WJ�꾗�J�-���>�'SM���E|p��h�ڃ���a��+L���:|e�&M�=���?�z�Yɱ��s
�E��F�Kʹx6�{{�ꝩ���n�X�F��F�R+նs�(;��Kq���(�7��6�ρ�]�s*_��o�Ie�ˆ��U{��I���U�	����s:ĹF~��ٸ����ſ��������쾻亵��սm��[5Z�*����$�V�{x�������o���y꾔y`>�}��ts�g�y�љ�d�7���]H �K�J}�Tׅ6=٨_ӏn5��	[d6���FdP��*nY��7��E/�qසnCȫb��
��;�}�
]�I�`�{*��׻Ug�׼�-�H�θ�.��!�
�ж����g ^����&��]������V��)yX�zw쐂��Xۄ�xQڴE��6�z�b�3/��<[�|���V7:6��u.��Q�%^lzо�g"���=���<��wJ���w��y�YO]��[gps��
Mubb��naӈ�f]��o�*��!s���~��UK	����������E�H�Ŗr/���o�S�p��0��?����l���������������%��(��Ӌ�'�&��Duwѣ������������Y�����&�4�b\s=U�gm���I�`�E�F���.��d�6�];f����'�e�|��,,@�C�-��qSj����͠v$��9�H����lrT�ޛKo Waػ���Ej��� �bi&w�����쫴Y�	����&e^q/[9��$J��*�\�@�u&��&�O�kQ�cOZ����I>����b�]|/����(����2�z�C
��r���U�*���P�h��ސ��.�Z����v�{����HZe]�E�2VJ�+|���=^UG9bل0������v|{m{Ͱ�ba�e�	�Gk��h�֞�6i�E�n���o���^~`�s�����ﯞ����6���Av{�c���DJ�C��>��N������Y�T`aӊ��=j�[w$�ݗ�4Blgl6����p_�+�b�D+L���fY����ϳ���賓����ya(��%��W�aK|�,�H�;���y��������W*�����7[�l?C;�m�����݆�q�w:�a��ұ>�E��_�͝^]`b���'G���c�퐼�e�gQ|�G>��;�Q7����9��e�ۍm�x%������?f���'���[�P7���UWF����ȄG��
^�78���sJ�~~zeX��k��c��ٵxhY�?t��Y6=ܛ����~���,#Y'�޷kܻ_����m���?K_6�m�{c{�wO��]���^�xs�Ψz���]&"J}ݹb��$�㫹���5�ڜ�O�o���u�Z���{o�X�z�w���
!Wx�Ty4;ʛ�Nx�����Ͼ���6�͟v��6X���3}�~r����0�{V��)���<�M�չ�=�+yw[Vڿ��_�
��1��S��5&�'���J��Z�c�/s⵴a���³{�v�Չ�*�*�=�1\�f�8���"�hN�׳��4��6��ȥh${������ԼaY�7��h�%�s���]��s��Z�U��k�hu���HXM���s*p��df���r�^q�T�*Y��>=�v��lI��h����[��b'Q�u���7�Ł�]�:�
dq��K�{�`�B�;���׸'ũ���)���j�'���$�>ؿ����e_�p�Â����lQ��돌ߎ.�,��ɲ+����;�g�^[^%w�e��9Czk����
lX���`{Cl����v�������s�3c���"w��ۭ'�L���ǿ�����j�(p��)��J�����;�/���o�E��剁�G5=����g8�[�`��`�� ^g$��륒gcGά�T7:��$rj�3 N˒:⇝�q�+X��1�}��4c����6�|r��X瞪�VN�ʫ�ګù-��^����A��+s����
�ciM�?+�vS��g���G�靖}Me1�Z|x��z)�s��I�q&brwm�ԣ*s6.�)5���Ñ�d��a$ ��:G�5t�\s�xq��_
��91#K]���J>��ׁ��)�j�Wloղ�ch�å��*�!��o����"��~��S��n�W���Ad	��������_W���WYK�xCH[��|�Ȳ,is��&�����H��.z�#k8^<2����N���?
w�],U��R#v��Q�*k���;���q0��ܛ-�Eaĺ/-"|�pQcCU5��������\T��kFU���կ˖Y��հqb�a��q�v��a<�t[���{�D}��O�s�7�L�8��������������=x�q236���b/��j�<�{&o�V���+n�z�.Ug=p�x��p�b��@��	]�K�������հr��{��nA�Os~��2(��
5�)R��*©�Ž��/��8����[x��B��#�A�1k>�Ĩ�v-ء��W9���W�6���M�s�]��w��#�o=l��sQp�FU�͎���M}���(��QE��U�~-��l��e�9�<~�am���iyW.���2����W�N��ق�9׫�,`����m����L>/�K��\l�Gz��9�ӹ��w�5m��G��oE64,޹Ƕ#XL���xĨvWU3������ݓ�P�72��9�� �V2�C������FᲛ,d�ֺE_���naB2�)2�m�'��a�j�A��{��3g�k��+|#�ƭ��F�����;m��|�m�	k◕���2Cf8#<����D�x�k�����z��)��۳Ⱦyk�c��n����]�w��F�Ȫ�����y��3õN�v+o����;���ǵ`�n�}�Aj½��h�5������w�p���MP�I1���ݱ,�:5h=E��գ�I��<�O�5�>���.���X�W�Tы�KΔ����]��IS� D��s���^r��o�o�����1��m1�Z=uߣ3U��+�,�j��xQ�TGGoo��?]��u%����	`��,۽g��Q
��sv^�7܆tX�m��˺�t�������4f��ڰ:����U'ۯ���s���$v]=��>�ޮY�d�k�n<Dw�} ��'���qF1`��m�ƹ�o/�ڎ�-�.?)�o������C����5����1e�5n�*��+��g��ށ}Gz��1�9{���Õ���AV8¡�By�v,$��91Kپ����'�8���b�;�(������z�s0�����װ�M\���߫�+����p.��cX.ω���l#�&��c�j����3�V�!�j����x���0"3����֧f������þ�N�@�^��r#�>wܖF�5�c��!N(?8�h�V���e�懴�1-�T��}x��,;�Xu�\�@]���NQC���~�b:��D�=��/��᭗[��~4L�@.�9"�NK��v��E��;�x��|�";C��K�.���߅y�~��$x_���9a'�^��+����D���'-�9|,�ũ�K2^�����ȗR5�eMf�V4�5��f�]��ѹ%8�J-N�j��F$�n���A{���X!Se��JHǋ��%�h��|�1ϱ�8=��4A�K�J��[��z���it6�=E�����Y:�Twu�p�v6�����Ղ�B�-�dpݾu���J�oSbV��g� J�^��p��@�'�]!WD�	\cϫ��cd���k�����||;.k�}2}�C���W�tխ���{��i����&��ٯnxu�oz���c}΍����ި @O��i�s�=b��wd�y�������^�]�嶯��:�0�wѡG5�U)�ED�iGr߬R���/��PJ �cq4������	W��u����A�mHplp�ȶG-�V�`��p����5�=�|�+B�H/XJ�}u�]t��v��l�>��P��&��c��+�����]�3@��1������-Bj]���ٖ6>��|���1�f�WIhwQ��_�{�gO#�K��˦[t���}ܦ����ܾ���Ql�ﵔ�������Q�j����9Z^b$��P>�9��염^�˫mM7�Dc����VʧX���{�X��a��n��% �7��Jw�5�T���)oƾ��-vnU��1��l��������|��V�&���c�Gq?'����Or�k��iv:��b�#���O��л�Ј�_Y�XuZí���������W��e���E��v2̫ۉ`����{��7��6���X�[N�.�ЯWk��m_���E.���e�fUL`���\��Q�=�]�`=_k��l_ݞB�ϬG0�u4�6�6ȁ;.�1��]Oc�����̅B�(gz0�����턕 �bE˴��f����2��_.3��W3=�Fw�����������_��������@ݹ��Rk5��v�۸�^@fN�A�+̏n��nc蠂6�qq�w�h7�uj;FDEڼ��y����x���[�����_@�v��8�%'�i7u �ۼ�`�n��6)+T�7V����w��6Xe��,<GsG��ۋ��7l�����_}&y���:p�iG8SR�^�G<��aS�htr��_97X�Ǫ3�p䀵���4=OE�_ʿ�}�d�s��{�=�NE]��dZ�G���9�����D��[�dIV�C9���~9���r��n`�J��' {a��I�=� /�$g�ޓ�=O�ַZ�H�f@뱜rt_�yr�i��AI.��6�����-t{ eǲ�T��d���n���ߜ�}�4w�����z�j�~1��}�s��tz�+��l�]���6�MЩ��y��&O��څ�+2�J�h+ä1��nͅ�]WO�-(Q&���98`�Uz���p�ӏ��ضï��w���3ޘ 12=Q�5zP�%�>���N��W���<��B{w�-�9��p�0z��`�3�r�� a�km��G�}v��g6ƞa%m��{tg�A�y�;�v-7r�K����۴*�����T��^��a�Lj{���;^�~5Wy:3ydo6;���2���4��E�#kx���C�x�S7�۷�~�lŁ�l纵
J�-̽y.�D�
C������c�/k{eaإh�]~<��԰إ�R�h���q��-M��zݳ@�<�ٌ-6L�aj���8�g��hCdz/l��f�4X'c��]Yk!{��m7s%}����@��2��4X�R���� ǪnQ���}�����<S=Ќ�{���΅;������\�+Xc��W�Q��-�,crQ��9�3��o{[z��L��2����/�Ѵ�fl�hZ��2��$g��8{z�f�w5�	=i��`���֞�S��j�9�����H/Ձ���Sm����e��V��{a��Gc��Mw�����~�{��U�Ǎ�mq�=�<~�m�)���y�k�{�T#{��f@���ѷ���c�g�X��d��O\N��򈳛[��7h]0���љRWQ�-����gHkeLn�6��t+gb��憦C�5��`��C�T7-Ԍ��Nk����=5J�>�m+A����ʺ�F�z{�l�M�k��[�flI���5��ͭ��p����{w˼h��,@�x�P��ޕ���~������x�xV���'�&xh"oZ�w�N�6�S�;A�v���V�Z}�O��諒����J���[���+{�C:۬P'�9<����$���G������������6�������7���|���J��gdʗl�����,�Fݍ;�~|��e��\�ʆCR57�6.+�+�/~����q�5��cJ�CnI��g��u��4ǡ�L�*�������M;�K�a� �:���Un�f~�ȱ�G�>�΂��ɧf���N��"�6��x�mF3U^v�pME������h�B��0q�Ur�[���A3.���$���M�`7�b�SM�ႷUgy�!Զ�V�t'LV����"h��w#yk�oS��f���#<����w^禽'�kTJ�eq�#�u6>s�i��׀�� V��?C�+����Z:7�i��}��J�=6�M�h�j	vni�|h�2�駒sOo�C�J���.�p��e$v�E�I��:ηK��}����6��;�h_R��] �V#Sk�թM�./VC����#��ur�7g�+.���{�cׇ%w7G?C��z©������c׷�:�3@�7�Me�	]:�\,n䐼iU�����A�oY�ܵK�=Z�Ci��v�(ka�.���S�ݶ,�|A�Z�.+՘4���#���Co*�f����ֻӗmrr��px{}����nzc���&m���$�r�=47�<����6N��M�77!'�:Z���o�8�]�g+e�zM�"4����������O�����I/{57vpe���*�d8xm��%�E��I{�y�BLxᾸ���$�h�{��Ln�� ,J�Q�]O��vd�����v2��9]u���A���Ҡ[����ˈh$�$��cD"��2��ğ%$o%�*������)ՒVD�"+Wɲ�.U 窥��������>ǳ��ϺDG.G9R@�������PQA+Zp���D�{=��g�U�.Q�\��9U��ws�E\�*DV��
"#�a&*}�쪽B�YD $��ZjTEQ��G(��PDTp��*��ȕ(��"�UF�TUDTvfU��)6���*�:�s$�"�
H4
"���r��G)���Q§t]wn&T�Ay�L����dr��';)$���)���j�^2��(�
�*�D��nnBTᗩ�\�M2�JH�D(�Brq�(��"�L͔R�TT�"�(#DQ�Z�[�E�p�B��Zd�i;��:˗�QDA��@ �g{���~�{E�;��Vv���6ܕ��	��˭A�`�S͍��c4sV��\�Y�aaSmՒ$�7UD�ﲺR�?���t+���=�~�"�[m�Oe�.ƪa��NK�h���v�����p&e��h��KGK�cmZZ�,Hwӻ<=�D���Y�Јh���0���Р�[H�RJ'Q|�����m�U�Qa"�]z3s˷|Z}+�2���흉��O�ic��I<��&[d<9&�(�h�O��oȔ0�!�2�=�u	|�n���QT�OsfA�7������kuv�i.�$z��}~���#�@�ی��B�NUP{켽���X��s'ڷg��=�C6m��n\�	�辉r];���$p�ڼ^�KSc�����ye(��v>���_�7J��8���w�A�dWl-]�7B�%�øj��_7��~=T��{AZ'�<�o셁�1�%=�)h���Bl䅄Р��os~=Qy�̸��}�_��??����t�z��������(G}8� �f�]�w:4�{��VU��KE+��������TiW���0Q0��skF��%&��u� N9�t+A���'0��hG�En�I>n�={\h븍-�)e��A�ę��v��_�ϟ�FT����k.ω�/_�aL5�l�� �K��g.ô��__k2��\N$7Bs0�֐����rb��l�L{3Vo��`�l���@�ʿ(��yX)VUp��ϫ)���L��w�n���&$���}V'=�WbKıC���9�3o�Jf����TP��VxX�B����5��6CiA��k�ytU[�z��<�<)�[�eX�F�Q�:��p}��v�iI-gX�� �=� ���{���0�׺>5��p�|%>���X�+k�tv[gU�V<��v޳��ׯ=�$����k�ϼDA?`���x4~[����{�Q�>��_u�ɾw�HR�K�{�\���H}٥,E=��!��ś`dG-Ԙ�ѻ�vd�|���P��W�y.hc�tE��\ބe���y�F�w}���)�q�q�sg����W��Ǖ�1P���/}dCc�qn׶r�kɻ�s�$:�ǫ*U���f�� ���碚&��z�p��q��0&�&<��m8a*� �Z.�p��rn�c�m�	����wӝ�ڳz�뭾dm�{����אח��C��z|-t����]��.���V��W;��z�3�w;;$&^C�[�E��S�WKWZ�L�i��oN��E7��DX�#�\ƣ>�]^��@h�f��}a;�=�����$�Yc9�\D��)K�,��eZ�8NGyQZZG�] �����պ5�.뉧y��rJ͝����3\��Z:�! $���Cg�Ά��X������g%ʫ�rk��y��s7��%J�(.��i�������6%j�NǞ.~Λût��<������x7�{�y|ðYi�������}�Z�n��ε�UZʹ[��4;`���ཪ���Ͳ5nZ>��+�֑0,�9�ў�g���ٷfʩn+�:�!W�=��st���vfԗ�k$mU����1���m���CV#:��C�Iu��w���>�x�9��l'% ��m�r��;ve-�W�t�[+�'�����6٬�=��LyH(_Pv��Iְ�(*�}��V�݉*���B9�bԵ%�������77g�.f^�+�bԤЌ��_R<�S&˝�{W\�m��)��OA�2��u^�W�{���}W�Z�I~3��e��5-=:x8�e&��^izѵ�=�-��� �i�u���w���F�,1"8?c�j&G���9(�=�C�_RH��|2��<���i[�=a����7���S�^D����W�w�_�y<=C��m������/�R�Տ�V@�H���#�� 3�%{n��H�0���� �'��(�������wP��z�v�U�G�ʏp�y��d@��u/p�jak��. ��Sβ4�]�W�1o�^7����k%U�n��k!�yN[�g���A��5�k��i���W}�Q�ګ�:O�p�)����F�S�`�x����7�<�x:��]�r�u�q�_'�ܐH+�-m�
�<��[���R�DC�hJ�:C?�u!Y��l�'w������mNχ�u�s����[�\g��J,$�p罌5>~�zݚFa������P�i�����9�r�����k����O1��c��>�"�y�����m\�.Ȏj���I,�tb٭k�+����"����}1�\m�Σ�W~^(�UEn⡵U!����]�w�/�m�<´�"Mz�����fn��I��[ن׌e�!���֩�� �V���?�F��h��Z��Γ�{���K�M����u�\.Ȁ�$O?{超��w�{�����(�]|�`��n�z-�ڶi����̿�A[���>ꋅqGy��^m����<1�V!$��:�I���&z����o��b�M~����'�;�lp7b�m7��6�v�J�ҷ�����w��m WO���HQ�����?w'��	��}n���E�RJ7�j�X�5�x�F�=l�X/չٲ��iД���5�a�J�i���7�w��cڳͺ{N���E�*�-��M�켾�$<�ue��{#,0v�>�/��޳�Z(�^3��&��EsU��r}���G=���"G�i�E��^?�#�k�nM�,��Nn��?æC�V�8�4��,�o���}��X���&e��0&~���:Л���ש�[��k	'wc|�;y}1����6���Z��%B�����:b�]��u�HB�t���~<��w%t�^�<���K�['��٩�5}Vg6���9��p���-y'������kd6��g��-�*�ә��ٌ�r�9]�.o�Xް����\�i����t�������PzM?�R�'��dD!p�u��M��5�V��_�ÒJ���S�J���E���Gr
��'C����;�h�X7h+��	�䅦������U8Ff^�NX�yɗ�p*`���k>�>'|�~m�<|�{W�`��>���x:����(Z�e�uČ
Hn���<�N�p�U����L:���N�������3�a��;�~	�E��ѫ�c��
�A�bv�>��L�^.�����7anrf��s�$Օ֊�d��Xt��G�5���)�[>*J����?�4�=ţSk�*l����$ϱ�1בn|QE���f�j��Oin��Kc,V��w�
�v*����:m�V����k�r6�۷R�Z�lɵ�*���pK��yr�bpv��w5}��B�lH�NE ךH;����L��t�y|�a�8a�@�S�J�r0�2rL���QUr<*b�*h4C������Í�"=gK�}ίy��mğ� =}���*_z����NW�[��	%F88[%�28n�:�u��P��L�(�	xq�59���Of�S�sZ���9퍀��a�r�ж���:�6����m�O�ow�̿�w*��d7�aoK�P[_�+�4)"�9伱�i򡊳�ݓ$��5��Gr�F>�E�Շ}�l8fлId��Gl>D��+�6�����V�:x�_��qt���r�]�{�f�N^K��&���%ڑ�@d��������Xյc+�߫c�,��]�؍[�Ү��d������~��#��}��xn>D%hUy�Iq0�7Ϸ�Q*��O	�p6��b���v(q1D��G��ȿG���0s�l��o
j�G�����P�t]1�;�\��n��u���N�'1v�[�����5*��]�/7��u��wp�q�O���͓����I6�x!,����#y���zGr��>F����n~�P�so,�2�`���*X�ϯ��Q���qb�U�re�[N(�m��hG]��3�h�CjP����@��K5�Ġ'�d�sˬB���SʽW��E[�S용Q<�sjϿ�>^to��65&���.�����+˱d߽�bF�^�/ݯf�5P�v�^�@�T
�a���8չhޕ��|z�,6r����&�NEi�����[� YK��DSb�<���a�u4w"�i ϲ����vO��^h��s6�`�(s�4=��V�$t�2V�Bj��z����ͳ��z�!m�$��::�a�l	�ݾW[\�p_ME����;�Ǘ�9<�'��O ��o۷ݝp�h@2�Zo;��uF�)\��ѧ���[+�k�j��km$9�j�cz�L�v,�
�f����Y�����<<}T��o;�k�Rj��6ݵ��}����f%�<��0����K�z��n��
.�z�u������	�k�M؝�s
I���۝��v9[��G�9T�5|�4Z���{>v���딚7]�x��pY�ٝ�.�oL�Np���թX���fqL�8��!��E�������M�^��z���3��N)�.�f!�x3%�H�I�;B�;��B�mv!�}�E-�<j���^���2oJ�p�o�@����ٸ�U�m�������=���]k���[�#GX�5G/��\1��(͚�y*6.0}�o毷<�~����-���h�|DHى�����;ꆶ�t�Ը�j��Z�c;�ݘ36�: $ذa���]�]��=~��Q�fֳ��pr.��Ԍ�y��iW�/'�l���$~o�9����H�p~������T��[��=>�u��%������}ͼ��j���^p ��uYFⷆ.�9��^,0�n$��z��$l�����g�USWs���Z14H�}]j�evz�Y�0�+��[B�5�5��^�:��,�%����Ù��Cj٦�i8��`�PW�F�g`w��&�����N�ʥ����ǛC�-I�@m�D�v\��W�瓽A�y C[yo��a礫����%^}|�yM���(�V�>!/'�����ݼ5|�Gk��^��5r�iW
�I�{���+=���E�//Ch��P���EG�X�Qt�+��N�oE�9c&ef���*ֻp5��Eɹ[�sQۥ�mK�f�3)SQ"N�%�Qf�
kY��<���ktA[���W��{�bLQ�Vh�w5)#O���H{Օ(-��ޕ��47v~�_<��ȸ���1��Ou��k-��OZ�ᅑ��}(j��m���;���a������v3��X�q��&�n�ޚLX��48B���ⷣ"1O�:{l�-�������^^G���.�+uQ�D�X`O��/�k\�L(�^��N��Q����R|�_�r�*�h[�lq��F�ų-?^[�v8ϡb��:���9	o�����^k�
v�������D'i��ے�ijfؑ%^T�
m�g�np����	�W�7F��M��kǥht��m���kk�b�!��n��5�uP��	�䁶3�~����|�2��t��ϫOVJ��0*`�Y�e��#|��t$%ѭK��7ٗ���g����7���%X�t�	P�oW����?���c��cmn1��m�����ll`�?��7A�=�` �m�@08n��؇1��d  ��n<�1�A  ����x� C�0`��Q� �� 8�(�  �ݶ�z�dp����;m�A��d�	��m�q���m�v�l����&�mw�h�m�@ v�l����8 �l�  �m�M���m��m��m�@ q��m��&�l�m��&�l�m��&�m�p���;m�A6�d��A  A�m�	�� �m�	��cP�D�� �0;l��hy����0���0l#�c����������?���������v_���_���?���������	�������=�������߿������1�6�S�6�������cz>�8� ���o��۶��6����}#��\	�7��x|��;�3��-���m�c��� )���Cm��m�Gm��m��d�m�a6�d�m��� l��gm�	��( ;m�@v1��� ?plcy~����~_�����P6�1�������2����0{7�~)�������~��[������筼��|�����'�8�o�cm�O��~��_]߀|݃cm��m���o�C���0clm�����pccm�ɭ��-�<��=�������_��x}����o�cm���6���� ���y���(��_����������ѿ��2���� m����� �o�o����e�o����8�&m���}0y�7��w��2?��cm�>K������7�-���G�}���7�������[��{�������������to����
�2��Al��������9�>�����"AJ"�%*�%)*��*�����J��P
�֤H��dTBP*�UElV��)J"�A6ͲlĢ�H��L�)�ě6Flն�M��{����%l�VԲl3Q+ZU��k%��)*ʥ[[*���-SVj��ZV��L�gj��˻]�^��'�ͩ��f�m-���`M�mlͭ��ʭ6�"�IMh���U�-�Zh�m�����6CJf��m�ͳ-l��b�6k[jR��������R�h����  ݾn_kv��;���ymj��׵�]��7g�[y��wn����w)��n�q�n{ͭ��c��ײ�������8��V�;�ݖ�+��emj�W��:=`un��m6e�����ʛJ4ھ  n����������|
>���B����@>�44(w��СB� -:�s\}K�����n]j�Җq\�WQi�ݶz���r��u�{׽�۴Vp������9�v�jcj��D��5�f��  o_�Qն����W-��٘uY�s��[���-q��񫻆ӭ��֭�+����,�����׮�)5��C��n]έ��wn���{�2����b��Ԩ6�Q�l�  w�N���F��}o/[�ڹ[F��w=T�k5d��t��܃�����]�u�wq��s�Zwm��s{V�m�ud���]��9�ݡ�ڊ������޴m��mR�bz�L�,�ֵ�o� ����	>�y�ʶkj��S����yo%F���vӺ�t=�wuݪ[����u�����Ruq]�N����㡠.��J[1Z6��5��֭6o� ���f�L����iogO{���4{g����ɻ��K����{��՝=�ysD�g���.�Z^���C�F��t�U�Gi�&ZdJ�c����"�5�� ��})B�W��@zWS޸9=k^5�����n��{�V�6��sڦ��YsM1Q��:��WC�D�-��:u�u�9��R�٦���2Qd�5�=�   ��׽ g^�� �盽 (z��� Sw�.�)��7�`C@���(� ^����h� o)��P��{e�RD�$)���%�o�  M���>����sqҝ�+��y�	/s��Pz
��P���� �P�x��@����(^�Ug@�Ѡ�UG��m���d�6֨VQ��  ���i@ýpz /{���Ұt�P��  w���AC+�pE(w�pz@��� U�;�� �S�)J�hF�4Њ{FR��   �7�FUT!�� )� ��� 4 56��*�� hhi"LʪM  ��~?���0g���`~���$���;`�!�}�W��7�yf�|J�=�4���$I<�Z����$��HHHhB@����$��! BH��$���ϻ����]�:�ɵ�2hj?��Yp�wr�QƔ�ZMlx�U�����yQ�A�r�#&f1��
ktn �e#j2`������!�L*�hu�Mc����%!�;d��d�ya�E�Z��un�IV톩c���`���*IB���b�%g���M,��)9F�ܕ���tBd2&Xlnٽ��%KܽL��p&��aDI��U�o2�qcl�X�.
���/r��b�͹�l����fhCp��J`w���aݐ5�i�E[��kjJ)�Ae�G��e��̲m�X˻�Tk���p8�p��J��~�7��I�.~�1D�w����*�r���H�W�^��O4eQ���+(�M�j�6��*f��n���.� �r)�4G��lm(�]�Ӄv�1�)d��-��j���Uή4�SH�^!B+CcL^�A�#.�C�n��qc��:#�B%�j��em�����U��0.Z �!�id�N
ˆ�I2S�$[JT��o.����|*�2ʩ44D����w�"�p�4eIvsK�1��
>�R��\�eխ�w�Q�j����c4���ʊ���-�D���a���u����\���х��e;H�h���$�ӗ��Y���w�i�pB�]�x2�+�U�Y�|	97 �!Q(02��ӽ�rĊi��*G�m�1m#9���&��N������Mז��X�'���h �)�M�fjU���]dLU��i�2�E�#��R��=�U��"�Ǣ�B�o;����\�.�}�q*:��`}wv/tc7($,�C%Y�cq�O`)Z��n�Xzٻ�u�)�F�y�c���J{��$M�V��h�����kN����Fb�6�N�ʻ���/!.�lR7����9t��6��=ITo&:��ZI.��r�#�X��wc5ն,U��Ђ�Ԁyy���5�{2�̆�2!��R�&�� x�m����T���[��c5�!�����92��J�V\{�iؤ!�x˶r�Q���~D�B�9�]h�@GV���,�{t4]l
�MkWԫvB��h+�7a�z3頉�5�R�l��uk
vEQ����S�*�c\�	�e�Ōt�
ܒ��f��MqX	콹k�0U���V��R+f���T/����a@T̻bџ�k��7�=���ڋ*5�K1-�tf��I���:aұ-����dѵwG%����;fE��jVR����.e�Ҁ����052QxT�Z�a���Zh�N��$q*�,ۭ87E�L�R���� ��6�V4K:f���"gH��%��˛�D7N�܃v��Ӕ[��l^�.���r������T�xwc5m6�Y����̓� �Os0a�RF��y��&�j����A#U������yqF��صd�f2�ck)��V�(����\���JSe�nYь�y��	�44㎍�.��v�ϭ�B*�T��*�`_�-�u[��Q��勊���{��,�i�``9{#���r�K$��̸�� �EZ��+e��1�bhA��V�E�Q��e�n��)Ik�V�����F�Д *�{,:�X��$���a����b�'�BsQ�[�N�+AQ,��'2
�l^<k8�ij�c�4աm[�]n�d�f��[a�t
+�͂D��\��V����RYN탬t�u�L�`]q�CҨx�.�!�Ep�A�e��a�30��P$�҉���L6���R�h.3��aCC�j�y��L�],z[8H�a���"B��6�^�a	�L$+6"��Fil�L!FGu#�G/�����R�Dӷ�c4����S�)<����"�L��X���u���f^��QK4^k�CKkc���l�p�m^��B�K�G�2��R-����?��'2�Y������%���a��}27��2�p� n��ܔ����@�\�F�%մ1�ߦ�4�j@H�Ṣ��a6�eXò�1��XXD�T��!�sjV�GU�BI�jM�|�H��5�0�
ڳV��J���NZ�x$�Yڭ߈v�A�ɺKt���k��ok%Z$6��m���N%G�IXU&���E�ih1֍5��w�B�c8w]&�vL��?�WQR�J­W��-@A�q�w[��m�bը����p���������+iÇV���ʳ�z*�0��!��LwϜD`����mÒ|e�*���k����ml&�ƢDl"���3V�-l3Xm�ɂ�g�qV�i+|ni�f��I��-9S�7dJ����LǕ�j�@�3 �F<,f��N��V�d6�J�5w)��
�r�Z��Z�7+(�.=���Ȟ*��TX@E�x!�ݥ�5��
f��ߕ�ɩ!O2H���Lm�R�oQ׈�W&�Յ��ɓs�Fjr-�P��>	;{v���"��kNk��u�*t��`&��cX2b�ٶP�l9�q��R�]�r7*f'bM�:�͵�S��  v����Mk��Z�CcLi��"��������$��i8�B�Vj��D��顿h@�5�/ܥ��$�n���S�i�Yz����!��j���1QۼKRiإX$�@6�T���v�����hi$����ox^�r#@����IB�ԌVñDl�̗kP��ޓ�)*X�q*�f��6��W[��B"��6J��f�M%������T��/m�g(d�ooY*���6������̤�4,˚I�	Y4��ь�(:7#�HK���X�q�`:�m���%�AU��Gә�h*Ʈd&Sa,Zf ��5pfؽ1L�=�R��#!��ڌBl����a�)����2ZHp��Q֭pZ�Ij컴io�eM	3��Kt�݆f�4�C˧J�?���xa�{sv���7�,��ɭ6&#��I�o.�K�7����N촫-��([�'�A�!t35�0i4"��x���U���-ԓ5J�J|E:���e=��`�����-������6m35����	i��fP��`�75�m9�S��fV���)l���A�T�̙���!�D�$`C6���KVn��ex���B�n��-���U�j��fe��A�\��bXx ����:v�&�70��Ǳ�:Ӊ�G��zs.��ŷ�v��*����
ʗ�b�Yh�L���թ�����$�#��"�r̂�Kw7,�+[Ʋ�:4~i�m�Ɉ��K p�h�bic�r�T��Y���M�ڌ�JTL�:8p5�(���f=��� �b^Y�����f±�!��q�2
���!��Oks�M[�-��y�F���7*�\4�mO���m/�qV+�-L1Eq&���Y�����v�kh�21��MJ$��fVjʔ����u�tb�ɀXw��� n��w�n�,�&Ħ�0���ַha�%�tj��`�N�& D��ĘZ�h5�޳�jY`�2� �m%Z���Z�Yl;A��YN3,��#���Ŏ��l;]���Ì���Uշuy�qͰ�^�Q̙p��I\���94�=kS��Pڸ++v&���ZW�\6�^�0ʄ�-:���j�K #쭛iR�[��ՍA�OYt,e0&�x�EԔ�$q��e�r�s/pY[Q'���;��HiWx�hJ�]�����?�{�SE��Qٌk����)̀7
51+��R�A�@7f�jj�*]bwn�hƾܬ 
ܵ#�Wiŕ�
��`�Z�J�@M��t�-�݈Ǒ^�cY�Y�2�^����NA��o1Ȯ�F�h�:OP{�NΉv*ٱt��NG/(��6�h04�e�i6v��j���&qQk51N�Qi��&ʪ���f�*:DSh������v�ۊ;f���ySb�ҥ�[k�)Z��e��A��"�,��l���Z�iy�@��i�pBn!��@C2��?��J��`V;ו��m+'�~Sc��=l�u��F��u�ld�>��W����]��Ο�m�����q�j�ڦ�
�ô�:��-�a顁'B�R�`'Q��`�.Yo����B�}��b�w�YJ�A��G[�̚&͸d�Iq���L�ZRT�{�صrEz~�ec%[��S��Mȷ	�C&-Tu(P�j�2n��:y�*��ի�oZ��ل^��k6�݂��p�Q��j�[(���tR[�@����Zӡ�E�+ͻU.�64L�j!7��y���A�'�6M�d�[,�I��*��ɻ1�x��"W���K�b��ՇyY(B �^V*���h4u�h�f�����bb�}�if^��� �cǏ6kIF�jTʷxE
B[zK���Fɢ*1��(Q���V];8����ƃt�Rn�WS2Tr��۔�����s(��@��l�����	K�@���Z$Ș���b�%]�٠mn,��v�F�Akz����xԳ��w���>�˻xen�pԤR����9�ɻc/]­єB���ί6+H���p�r�)�7����'r�k�D����YJ�=�VJ��r���Ұ��^*K(=�e��vPU�#QRaƄ��㦱U��L����hb����ZHoXz>SAҴ����dKD��F��א��S�����c�nʭf��Rf��ʹ���j���,��l�	9L����A���ѻLj�ރY���Q�E��tZ�k)�4�5SpTi�r�]^L4@̇(֣�e���A<�T�)���R�Ԭ�ށ�HpM��.���]�P���͸k��)nmn���Tr�����P���[u9/1���`�4X�n���ū<KX��x�u��0�j�bY	��Ū0�����&���b����S��C�@6ibj�F��ϔ��Fs0�Vn�):�$N?=Լ�~��R�����f`ɟC,'�c7��5�Ai�'���kJ�JB
� m�J�HT�&�ù�ʻ*'��,h�����f��j$�k��S��l���];dh��*��(%6����6�����1�:�E-P�y����:�!�6�=��H�%I{Ce�J%�7��l"s-�p��IGq@c�ͣ���7xD�uf�gl��'r(K��lں�w�ef���͠X������ó�1�xHmPe�0���λ��V�~�َ^�eJzH���:n�ޝ̚��j������6��I=�r���uO��4�����&Q�����kj��n�K9b��iY�@-kt���[y�j�2��n9�K�R���2[���,hݭe���D�8l٨�-�a�k��j�RAQ�Ii�k��� %G�su�2�^���e�4�c��J8��-�7��]^�3�֘�ՂNH�*����Y-P�bm��V0��w��m2���6@��Y��rT��M:T�iǐ#�$��Dř3eilKP�.䚔(ЛwH�v�P�W@�o��eF��SE��ҩB�	�F���Ԥ!5� \w��� U���Z�V�<7@n�ȶ(���Ge�*݈�:�TIlVd�ǐ��/	��õ�2�y�-�cX�];E��z4jt�I�X{6i�3�%�[�e�m�я^]O5�B�j�����S�Q�@\�I�-�XA��*bf8����Ԑ�˹	;XX�Rf؁�
��
����m���5e��ܬ߆�X;BCE��:zh`��Y��]�A��&�Fc�Sb���C�C0���F�S�b�C��A�1N"{/3V�KQ�P`�m7�m���n��rf%��ଛzӨ�-cz�A�{2���+�j'{��yi+w�U�ԱAT�k�eZ�*dX	"�tդN(�w��#���l�2X5�Ÿm	�e��fͳ[�J�Vt��1��J��r/��,a��FAF�5D1�4�x��"@��ԉneY5(;���e3iIPT��;�2��mb{�eL���u6Re1���Z�H����"�l\=�j*�۴[��A��*❑+
�,��8���29Gv�X��ma�L�0d�3s���cAH���&1�<���S�V9����3��w(�c�>��Y�l��/oـ! .v��φ��r-LԈn�A�D���F?���h!�g��9:zh֤��2(�˂ͅc0RƳ.lQ�a�Q֍2�[(*����*�����h-0���7#9�R���m)fSb���&��PƩɇ2�a�\2� z6^�t�]]D���H�`P�{�/P\�!��/{y��+m�&����"h�&�(̺�$qQ�-1� 5��ɷ[%��u�n���]P�R�tZ���qݷz�ͣ�����ue���Zm$��E&�4g]�P\͚�wF��[�]��I���v��M�E�h\M�U��# 
��Yl@P�fY!Ĳ�����BV�X�R�oA��a7�{.� )ef��X���8�ӓ,���%���Ň$��ܗ1�r�؅�4"�2��/U�� AA�Ypж�I��޻��fG2�R-5�����oqڼ�M�;�݂5K�8Qbiǰ�����E�)(J4�X���x)�\r���r��t��F�0ҷ>N��u0"�$�IyXC�V$�n�ԧ�%n�`�
Z�$]2�㭗em<b�dSF��(���Iec�: j4��2�P��z���4�����% ���D���晢�/��z��u3 ��p\p\b\�Ͷ���!A�����-�ߎ�׵'S��Q�����t�L������-kk�m�Eµ��en`�KEJG%˚�(D�r�33F�x���v��a5��Z.��э�X(��K	'\��C�!��hZe���,U�A��X�$��f(�S��w�g>��e�q�m�#vU�:Z��:rz�:�X�{�u�����G��TiF�$�幩v�<
�m�3@})&�����/�g�U��^��N�H�fQULz[^�z��c�&<'����<^�љF�E��C�ݘ��`6��*��z'
[�k�ev�b[ԅR�Ԩ�
[���b�qɏ.l�(�&o+�f�������=���l���Y�!��V��`��`�M�2l��9^hv�����Yz,=��+�t�ښq� U���Z>��Ƞ"��:�x��e��a:��~�6t��������vV�Ҕ-���B�/a�`t�̢�`�i���*V/�����Ŋ�w�n����V���l�j���wS��]>!�*�[�(��e8z�k9�d୕�q�s�\.�]ս��S3Kt�?-�����l:���5u����W�勾��6�|�i4~5�wQ���\�ñ:�I�Oj
���,&��V!������X���V^�&N&�rܳ���@ݎ���V��%{���2�mpVL�p�h�����nn`�xt�n{��;��}`)V��/f;�w�]%J�n�6����Q��D-�t���ӷ�p���\ �jA{�(4�jX5�s��@��O�h�F��e.b�NWz��jĚ�qd�ov��qʂ��gp˵�+�o5;*�`�Qخ���o/r}�Xֲ59oJ�Ȕ���C�w2�nf>�oa�C�j�}њ��hc�n���C183L<��JG�+Y�$v��m�#\w�zaf����*o�)�����\q����^.��Q�|RX�>���d����0a���v-G�+|�GDh˹J��-7M}׵n�k�H��z�E�7��,�Ζ�����<	�I��˚q�Y�Hu�Ɔv��؊ƭ��/�`ڑj�����T�d=Vf�n:��k���7��@gI��\Y2_es���J;�H���h�{�^Oׯ|/K���V�]>�]o��ag��a�Um.Я0*m4�� lÅ.\�h��EL��7��5�YoD|�� �W2*5�z+x��Q�u|8>I�ӈq�Q�A�������u�kMtb�ݻ/��	Qq�X�Ҋ/��jr�9���5�v���5S��&'Rs��kn�t����$�ݧx��o2E���VUszF�)��yΈj=[��9�^ZU*Ȃ�����>R\�gq��u�O2�<	ق�ӗ�5y��t��i�1e��X{m܁�W6��F�-0{IuL��ڷ�-/:gs�o�c��;^���W������[����r���Y�PTb��2Z�5�i�תZ���eLN�;�&l�df���s���AV�F�]�W�s���c�������������ܣ�� �F�������X���p�_�[�b���5���
n ��*u�8�g8lHJƮ�Ju/����-Sqj�N����=sH��p��؞�U�78vB�Oaw�ݓ9f����><�\�Z��؇=/{�3�k�����)TX�s����pu"�x�Q�Qe9�y���t�:㾎p
#���%\��>�g'�Q�	�8H8<�,�=�%�h�t"��G�_ ��>�h^qH�n��3�����.wu!���t��F>�-��%��2�)9���o��]N�pƥ�uh#|sy����;2�����=�=]	W��L3����`�:��P{�� �ÿ1�:u)`T2�8%��{�-��h��=Y�[w� ��|(l}b���"���pd�z	M1Кʹ{/eW���{�9|`Eu�9�p5�^�Z��qĢ]�+(�Â���$9plz%wZUl���ݼ���w��w�_pҚ�}Y\nŉ^2��G�GJ�Y�v��;�m���ĩ��K��uǶA�1ɕR�(���Iv1��߸k}�m
�lW�K%�Iǜ�R���r�_H��ӍM�4�<K:�&��r8�G0[�YkmU󕯐�(�
����ۛ�A���㹂�'���im���9����Vn�K��y���g\�gb�0Q��0��\#��5��Yپ���t�]��H~�ÿ��*�!ި��II*W��W��_kݫ� ����/j.{7@[z��8-�3^���ѥ[�s�T ��n�IgX��#��e4);�V��gK����^=�'4c�Wv�[Lbf����V�x��'�\x�o���g�D�sښ��2��Hf=��1��) ��pY�-M�/�|&�x�tfF:����+�"VM��b��6�<<DOH�=�kh�-]^�������pꭗ�5�gĆ��u���������]�,�9��^�cr�HZ���=&�%hp�7UՓ%ty�1�Ѯ]�H2���e�;��q��6���|���|We���mL<��P�.��q�ṛ(��xV��ݥ3u�p���M�#;�^Z�� ��}�Y�A��m^�_d��/[�Nn����8����M-xLu&k��m��څ�!vd�B���x������i��\�Y�U�x[��X�~���u>����P�2T��1��yl�]Ȅ�̸�ܥwL�o��;.��ȷs[��ըn��Y5���f����{�FZ��S;�3�
��v�u
����w��OOe�=��-My��*jy��u�44��;�q��znq���#��i��k���ʗӒᵚ��W�������I#�KS8�%4�7�J�����B�1n�,>�n�N�@`Q�$�%e�w=����T����4��:�}p�K�l�Ui�݉K���/h�d�rVE-8WU�9a�Y��E��� �ۡ�h$2��*^ٔ�h�ٓ�)kk�f_�לimf���eѕ�d�P[X,Ÿ���nh�)�U���J�7�ّ��hԹ�-񙄂-۫L3��o����}R�B/��Y����v�M���k�y�Q�Z�'��B�^�f����镣,ޏ�J�~�9�!����y����y���7f&��L�O�:��G)Ee�%�\�9I(R}�նUɯ��Um&d��7��m5M;獵��fTr��O��zM����w@�6�9�V���Q�����Y�l�*�6�5.��ق��F˺�eR�̵��M��}�_c\�(/_[���)��[�OmҊa��য�R�^�M�����X;K�u���ӱ�ik��w�5�;^�;G��u��Kr�`8�޽��4�ԗ�#PpҎt��X��h]��VdB��>\��7SUb�u�H<�̷���c�b@�iX<Ş���as��]B]�ģ;*�uj��Ѐ
���b����9��^0f���Y��sF>n�Ac�	ykU�Ӻ��&eƦ��o�On{<{F����o�bq��B����n�V�9�}ӭ������o���А�������$zZX�[����+��..5j|UVUG)�}y�G��y⾪U�!~L�mo��ɋ˗j�y��^հgV,��������"�ű=�K���\J��w&���s%�x��o0�_�,˛{��C����K�Pl��	ũe���t��o�{Df���
�oGrs%�Z���K�����v��x"x$D����qwKv"(%}�������KQA4�]�[���q?�ޥx��[�̝O��`W �Ρ�U����:<ԡ��ѮB$�Z��FÅtMf�n;��2�[p�Ukg��GϞms�#=�+A���P' �;������o��uY[�q_�+EC�ocgdӝt۳gf�U�W�hK�i�����R��q{�f��R����eV� f� 1�yj�>=��l�;;f��^6CX���K��O�j,��%޵�L�����z�7��jg�좯(��3j3������C�Z����uy��մoP�;ʊ�xi>�L�qI�Qq�T�R>FV�*};]���pa.�抡��7=o�w�q��Հ�)���T�Z�58Vm	v;� f�F��-5uӁ���L��Z���b�jltL�2�i����3�+�����#�֞��)a��v��X�[I|�(�����ӻ���CDScZɀ���X��+n�2��Īr���=v�xx���M��+�.��~�����]e�2��c��R�w��j��%d /��ھ xnoH��)��u�������'�c��:�+�H����[O��aV�F�,���#wf��*�Q�}�vFow�N\,=���8�Yƚ��?7�^�>3�/hݽ�Ӫ�F=���i���cՁ3/B�+#A��Lf�4i����f��=��9T��o��v��k;Oe�Z��^[�\@�top��b�P�J�پ]�"xV<�c�$DSs��b��\�(h��*��h^-�5����)��9�{^G�/�^o�7�,�0!��5�{vq:�ћ��9�gH�ãy��i=ٱ���[x�k�%〪�˺\ͭ�0-��z�+7N�T����_q�]�&��D�vf}6�v����Y:��o���6����vưj���-\|�7d�ӝO2�䝨�^;8�ϟ�\v�W$η�eqC��+#V�Y%k:�3��>�Fy��E�NɊ�z��[8t�Ѵ��$�__L���{�qq���Y��f_/a'��%^Pl5q��1c��J��B��+��b�������;�aܤn���΍�R8���YW���l�#f�zf]eʺ��#�I���.�@��#@Tw��X�I�̩:����':�2k��yQYx0-v�	s��s�Euf��_4Z��H��Pq�fS�S��nڦZ�W6�;�w=��a�B��:褔g<�c�N+�ͮ�z�H��O��1mk"�Q~ 	�:)j����=ǭ^&�0 �s���oT2�v����ƞ�+�81*Qs��bC6<������'��/���к����c�頤;3en�)۲`7agc�"��ǐ�T�b�����P��^�����t�)u���o ��.���ޣs�͍p�{�VTJi����qt�/�����O],��$�S��P�۹��w����W�"8�b�!��o]�����H�tg�b��P#��cZ�s-Ϳ����S�`x&���N'l�]9P�(~�Ť��7m��p��f@{���!��#]�]݄��ی�Ycr�#6������f���5��nCo:����1��v����NS{w�W�7z֚�X��^}���E0뷻��a����\����+�\Ӱk�}�K���j��o��֍���w��9l
���X.��"GʞW#'>S�*k,�����*p��HzIKj�b�7��8����L�52�;��K�+1�P��p��d:]��r�88D���=y��_����ͬsn��k�5g�i���5|�k.f4Lʕy!7'kU8;��N]��WMN��m�8@�+�ٖo:N4ZkYu
�g(�K���d����q57�₏:��V��2������t#�m��n
"S�{x��T��{n0�u�)������;I]R�2�*jM��Pgn�\-�2Mוy�����: �s�P�$�/Vt�o��LuƱ}36�I�DP� �`O3$°
�ɳ�@�d[np��%���osBf��o����T.�k��v��d�5�8��tUܚ+��=��s��L�u/o�F��a�aVñ�#���
��d�'�tN�����<:�3e�&"c_+���'XՊ^E}��Nx���|"�Y���ʟa�j���6��Zxw�A<�Z��^J��V��� U��7Mw�_u��H�����f����ϵJ�N�P��wkKdɢы�RAQ���>����1t��%K[��Q��&���傂�OO��G(�T~����v�N��-�Zq��y��X���e�IƩ�γ��g���ɭ��.ُ���ӏ��M�%�r�]��%����LU�:����+#�;��83s��b�j�	������u�T=����$���J���`�ev�|c�F�+��T��.s�|<�2S��ѳ��5�,m���pD���ۉ����e�~��Z��Aݗ��d���A���|�����b-�1��ɵ���.�H�L.�6���Z�xJ����tP̦�$����g��n!j�<��Nc%tA-�������M�_.RE��]{�n�*bbUv���k�>�렵�t�/M�**:*�-�W��T�)�����ض,���������щ�_Cc�S֍C�t=+7H��Կ.ճ7�=]�.5��3��E�i��@�����&N�j����jaS��^�qfx_u�w���X����`�<�u��y��͸��-��0�v_r���0��F6�b�K�c�O��U�P�*g:��ְt�*|�h_f��p�GjN#1R�n�^m��^m�A���{��S��f��.��b��p�)�v"�v�B�L� �vC�r��9��X�|&��	��i'M9p
�1}���5p*����b���n-�Jj���iv�u�/�B�o0>�[����B\��e]��2t|�t�h1cYF��;G�ݢG�s��gm�&�.�ٖ���b�L�w�Z���(�'��`�*�W��W��Rٕ����,�==�'���źUӷ�*�n��}�pH>=�;0�ԝݜ��왂�۝@7O�Dvxd��S��]�=��w^{%���L&а@}_.�]\�L��f�iY�1m[��������>yx��"�9Aq;�"3$�i���=r�w1|��SKwm�T����Y8K����C���Ư5g=꼍$��@k8N7ۜ�F�w���"�=}kV*���Yմ�홰�qͼ�͂ڰ��٘L��K�ܬ�W� ���L�t�Q[
5c^�|�F{z����vڽ.�½�yy�~���=��+�����[����II	�{�x{��+x���C�2sv����?���ӡ�Lw��'�*�+yV�!Ên;M^���35��:���{t��N��_$r�k:<�Ѳ��A�f���bc+�Q����Q�����S�?��n��ǖ��c�XDP ۏJ�;�>��a1q�>����2��^��0��w}�p+|&W����.1������D$_�a��a67zN�*!�K�V��n�ۄ.�J8dfeL�AȘ_a8@2>�V��S���|�O,G�۸w���^�6�e�!��7*:�De����>
��Ҧ���$���Vo���������L�!b����Dm]+wA�M���zWe&x� �c����"���Oӕ�/L�C��ټκ�R��Q;��u!}���@�_�PT�6�䦅�7�����`���/p��	E�fc%nX�
�J��*�,p��J#���v��Gkڳ]��8n먃mnd������|bYM�m�e�k�
���&�Jx���yl�H�T��ٙbѰ�E�O:��xS�(���R൝��PY�^8�uo��֖�.wl^? ��Sa�SL����0u2Ĭ������I=8��04K��DCM�愻�V��C�V��Z�Z�'���#1ey|��Ρa�����9mɞ��ND�Hj�{�`[4��|�Oe�M;�j���4��޴��J���\K�,{V��8`aQ��p�����f��z�Y�sɪ��l�]q���6�_,Z+���p&�j�J˸#��,'WL�$��q�=�*�]�u����*�v�j��5ئ[�3�j�A���d��� �7���f¢�S��j�@m#	�� ^.$ܱO��wZ�z��&MS�It���:��T�ɹ3�h��ǈ���y�A���S�[^b.7�M��s#�f\����u8��w�U�u
gucP�7�}B�2��i�9)�ufT��}uB�y�醝��'�}ot��,�<��^ݕ'���1�xǧ�K6��P)G��+�MX���h�#*Z�[�<�w:��C�ͷ)%{���:�4�~���tѶ\��ńWu20����K{8���}��tUr��P!<y�ed�G4�S�x5�|���L��sppҋDc�A��lJۙ��T�x�"�R�(��us�G��ߕ����ЙC�j��L�u��wW�s�V�C[V�}�X����{F�صU���@UY�}j�Ҋ7��k9�iP��O��s�8��nz��q.ӣr��:�sZ�������q��wV��ڳh���em���E�5"�U���S��nVe9kY�|G�x�׬Њ�=�k.vR��s�$ ��{{O>���gf.N��(d����%��"e��5�2C귭��G�.�,S5����G����=)Q�8v�չ��εX�qf������N�Q녋����o���ʹ�r��2Nw��P��tTw��6��P��y{z������[�=�� ]��-�S�͜��N���n� �3D�d�����S���=��+�8������ςA}�nkc����_�7�/��c5}ڏ�tyL���.����p;լ<�]-<b��
Ʃ����,L��s2S��.Z"X	��М�ږ�_nn��e}���G-��░��t�3>tq��3w�V(��_6���+U�޴����VSț�/@�r���{���:6 r�d�L��}tV�z��=3�=�^���Xse�+�pAʗ�h���|�qS����mfֽ�Q�]��`��������M޾��z��1^I6���o�|oG��2K��`��9���xp�z/&�yT�O�Jl+�V��]���v�9U���A%t6o[73 |Q*YO��'&^�Y��Ia��p멚&G���OZ�m%� &��I�̢lR��Vk��>�6ࢵ�vWҏqRw83Y�ܭ=tn�s�[A
�n�2��X��y��є;Q�%f��ެ6����Խh{�F��T6̜����-(3CŇ�+�`�Sdn��$�{9\��k��-�;��hGl�9|��1B�[MAt�?dJn�Wf����G�h���}�gPn�h�>c*~G�9?�`�w���F͹��#����xv�ķJ0S'[�Ԟ��Lt� P8hC�ꩆ�Y���뱥�pX۬�t���]��]oMW'�(����:�q�Ӫ��$���DR�MvF&'J��)k������+���"�S�1�{l� �C{:��Vs�U�NR�uc��2�d=���!S�H̨RZ��:����I�u��Iq������vS��������W���\Y�e����ggV ����/gI�#ܩ�_wjU�����x���Eu[��]C��o��� � �q��-<~���{�Zo�+�=(.���l���]|2e�S���j�m����K7�+Y7�D�k�;��ve�$V�t�Q���0��L|�l�����/%�ǔ˺}��Nekǁ�V��o{�5�Ġ�%ϑ�\3�@t��6�m�[an����3Jb��9{�c�Ԓ���Q����T}Y}:��*�s�GBܷ{����}n���n�C��5��o�L���,����Ŷ����^���	�]�e�)�w.������n�3c��Jэ���M�?�L��
5m��:�p����Cy��{6��/_9ūpehan&v��#חn��Zl�U��.�W���$��,�Y�o/��c��!<7��'��W�h�l:D��
��E֊|S�U�:�����y�ŏqZ����7�؆�1���3�w���@\:�;�ޡ.� ��NF�7
z��D� �N��:�:���=�l܈�e��R��ԻHsh��B���t�6�^��|B:�O1I��}q٨�n��7iv�LJVI�1��8�|+:�k���\�:K'�M,�b�m템+�Ӊ�6���VQ���V`�%��(��/�NG�u�u��-���3�*ׯ�ѵ� �Ķ���I^�S� �ۖ	�@TMh+�77+6ZyD���ՙ� %(f��v�$��ޝ��ˌ��W*�L�XGMAک슺��<LSnjsq�h�>���
���3�x��mCќ|�r��o��	
 �yJ���
���n�Xq��s̙&���M�i#F�H��xrTv��)̝��f���#z1\�\�ܠ4KMq�)K6hݪ�o���X$��I�ZN��
��	ԯy��a�7evF��i��2+�ݑ�x�E�z�pdh,�{�v��PQ�m^�k��(��I�RpzNz��궍�4MCa�y״λ�1us�1�kn��&���I�r6�qԢ.����m�3r��uû(������O��i��TA�*�N�'H�[����1]����Zq��� w��I���_vh�*ɼ�s-�T<�6_>76�o����"����so�m�u6�5I���s��c�Vl�ѳ�(�'v^ ��)Kᆴ�L�ԭǀ�82|�nY2i\3�J����s|��W�"2���*���yDς-I�IWu��մ
)�ZF���\�#*�r-?�Xzg"^��{���}ݺ���id���˷Wd/e��x�n���YZ3R�T�oi������� �Wh�q�u�b���ZH3a�Xo6�����ǓZ��9�&v뺔!!�X�s�\�"r����|�0��6�p���LV���,���_j&%.�S��ۧW��T�uU+�Ӝ�}�]W{�eu�����{;&���n��,�H�I&*��k����w��G]�h��=�l�Z����/�}��*7����wU�U����UoD��{�4��K�K��t>����(���1`���&��!^RXY�X�J�����}�Ƌ��xZDP1�.�'�||��#n����m�aY��2�wG�]H���X�� �����?eC�;��8�s�j�.:�7Y�|hҙ�e�^阝X���ȴ�l����=X�
�H�vcA�ۏ�.	�k k�=nQ��G��8E$�9mZU�ۗ��e�x���ޫ�0���'b] ���7w�Y��X�u�����w�:kR��3]��պ9�{�w<&�ż�:�ii�j�Sw�c���Wj�_V�S�j����ͽI�"����|�T���%��1��n��/��4JH9e�E���Qt>��q��hD�%�m��W^��<E>}��g5Eu�t���ΐ�q�=|�,�ݲ���Rm��0f�oaO%	E]Φ�Y��M�Ȝ���󡃝�S{i��^bIӡ�i���r�;Uw|����w9�gJQБ̘��1w�������؇[�^�d ލ�1ВVjCWAۜ�w�gE��Ge��rΘ$A�wN���KC*PkM�����>��) S�z.w�q���;n�{7`�<[�~X6��z�'r��z.m����:��qgi��pҷ��N�`^΁-�&��ט�{���V�+�h��\��
^b�?*���C耴$tlɝ�pC���w���1k�b�Y�V9��e=ǥ��.N/�[+z��9�->�j�*���4��C+myv�BT�݋�Y3�,���ڲ�s�8wC��i���\k}O�9��C��3�5��Ӂ����5����x��Jg=�[��-;Ek�ܷ��9nΊ�~��gP����>ǘ�ڧ5���X��<Տ�9�ᗖ��}כ��� ���I?��s�]l�Cp�����l�/f�Mg���vh�	�Q	����)^^ۦYt�)Ʒ�x���jVݶf;4�����i����b-gL�B>������@8��r����0]�E����޹�U^	�[��mBt_��o�bLQ�`���V�s��4�C��
�n��]��Y����B��|���}��z:3Ń5�z"�c-ؓ���t��m��/w��N#DIr��tT��U�.���4Tl]*�"6�)�^��$���C2���(,Ԉ�X,�š��]'���8���}��S+F��3���4Z�X�m��nd�"�	�^��@�����K� `�����v��+]�������JŽ��x�RU҂��*�4hޖ7���V��5"Iȱ�e뫾�c�z%n寓�����-M�eW-me΀�
��t�1���S^����U� �
�b�eǐ��.�f����A+�G�������^��w��of��gz�踊�W�����!Zi�"2�*��v�yCx��֟=����ڵ�v�GO`�&b��-9�r���U&<f���̭�m<Z�U�	}���_k}S���Q���f���뛳�f���S��K^b�F�/��DG����#*4�';ǅ<o�秏�����|�������������5��3�	�G�̽E՛F��R�'�T�mR�M[+���.?�mc��tD�B[�dy�`��Μ�VK>���B�6DUqʹ{fߜW�Ok[˰�(�x�A������K�y�j�}��(�qa{��L\ܠ;��m�|���v��;Zk��1m��)�s]��ou��)2c�;>�N�;���E�A��b#�r���ı<��.�t��i�P�55�5d89")$�羝��i������:��y�'p<I�c����A9j��os����U�cL���'�y4ܵ�w]���pf-NS����\A��M�ґ�4�a�`T�J<��	}La��nfT�S(�m'io�sQ�4��N���Q����ke�N�f7����&��"�7��b��c$Րi���GU��"�bNzw���U�f�|s���<������ѧ{�Ƀ&�L��`Rs7nb�"���7Yh��u�/�J�/QR/9����ݱu*�R�"hC�w��τH�@g�<ņ@�U����svl~E1��B�I����9�p��`��>v�)n�ћ͆��5cj�S�ޒ�n'ʋ�8��3)uj�qh�)cc�`�iP6Kù�C�t��B�Z�������6S֎��ى$��Wa�t�R�P��7p���V���!���n����wJ�B�Ņ�er	�b�si
 ���ͼ�]F���{�[gn��Dh��ws�=���K�/$��-L�pͭ�B�'�Zze�Eؙzu`���[�k��w*Rd�Ҷ�s�Gv�����;i{I��_�7x��ն�6��iv���\�5�	�75LMuwe�b��C�j�3���G����]i�ʉ�+DW`)b�I։],�o��*����Ն��@q�̰��5Nr�f�2���&A�vo-�۶H\g5r
�P�6���ے�P���%��/����g%j�%W����}��.��Ge�lN�$���f`%��d�*���κ�Fq�h,��Xt˃�)�����3�0m���sSM�D9���:,]��v�X�)#�kU���u�
���I�}�U��کлn��X�KH�u��䙮wvs�Q���]���o����[��&�ǃ�i:0>�7|��K���Ka]e=��T����GO\�n����˘��#�GL�	湫�S�Y+;d>���:�6h^w�m���I�x���ӆK皺�2R7�UvP]A�L�9����M�7�a�ie+���g%�s�]��←Iv�P�~*��\��p�:�u
�L�G���FDÒ�>�yW1y�)�o��A,��T�.;1��E������+���B�f���E7�\Ζ�=ô;jO� F�{Ԃ9�kfU�5�Pv@���&wn��w��%��<���;�>f����
U�w��s�c�>x4�NáS�u�������-�3�O.���>:ȃ V��l϶u6M[���F�e��J�^������m�uܼ�N�u}�VnUtڸ:��}���i���������y���*�>�
�e���r`�뻳;H#N������˅IwPW>B2b4�h�ɗ}���S�X�L<䈣O���gs$ݝ�]}��l��B�h�	�ī}�D����4Z9O��:H��	4	TH}$���+O�:�n��R����e�lɅo^�����t
o�~��ס�bo��>�;�62(0�T�o��r�5{Yz�>Z1l49\ıy��mb�;ZLo������-��j�zx;�<7�*F	����Yz���Kh+��{˹����&2�b6'p�� +���j�FS����]��B�H��:Y�ñ�g_ h�v_sUx�����|��X���n�ՏuE��<P�=���O9f����!��9wKnFu����ӷw��pl�s��2��O�z���PS�Em�ڱ:���?	l4i�ʍ�X�uu\��{A� 5f�Y���CWP��f�{��8¼�}�^X9zW��k~�|W1�+e^D�D���B�u�V��.�݅�kY[}Bd2�e��uu��{lgq�U8|��7s�G(�C��ϧ�q+��/��HV;�@N���=K�R�S$˲61���h���HZ;V��gX�,�-Z���i�m��F1�a�I$��O���E��s��4q���O�VmXR�m���p�WmKX�;_{6rm�F�//�YҨԤ��H�Ӟ��}w�<��f~��nؑE��+(�
��X+UQQDdQUb�,]!b�UUUX��V"�%eZ�㈊�dAEF
1���UV)U&!Ub�IZ*(��*����e�UQ���"1E�1�DUV*""ED��D��0TD���V#*ڪ �E�J�f%Eb*�����TEQeB�(���Ķ�QQ`�"��+1�`����%UdZ�UX�E�� �X�-�&Q����*��9Lrk2�(�#UUQ�Q�(���q�UV*1�*�(��e̘3)UE-,L��5*�#���TTTTTdU� �j�1*�Q���F�0I���+���� ��*V����#�*(����Lcj��E�X��X��Qb*,2�ĩ-��V�b"��b�TQTEG)TF �"�`�IQX�1YWA�*�+ܟ��z}s��7�����>S5W���Ǘ4{;6�e�Z���qn�Zߔ��i�s�]C'RЩYY�^sސ0��^����ݚK����x�<}�p�7�t�}�7X�*#ym�������MS�p��@ng$W@#k&��u���J'���9��g�A4wA��5a����6.�����^ܼ�?<��7N��{c�Ѱ��֕��^bᲅ����϶>� �97է�=�)��d=˹��9�^�y��E�U����<��!AG#��tk���Վ�xeqxm4��	s�g�z0�C���V[�/��z}��U�i��j��c��ɲߔ�8)�3"��ʵγ�" �!"�+ʽ2\�q�Y"@�k���+��B�ۮ�^��{�(XQr��S��s�)�m�;3�N@u��Ь��B�d��r��߭�Ӧh 0le�M,�f��Z3����dh[<IÈ�W?�5^��	O�ܮ|9�Ӥf�-_#�E�VX�z����6���Lu���1�N����������}�
�,k�((��om���2,Nf��ڒ��D1�o����U��ƺ뺂xg�-�Y�p֥%��7���D`�*��
�}2���Wg#�zѾ��ݽ���E���C$/t��V���J��U����1"�}s���vd}����$Z���|���c�/��f�����y�Fp�*�<��Q͡P:�z�٢v�<K��	�\me����J�@=��?z��7^�'�����i������9�!D��@���n��<hX������N͐Du�)�jwB����������7]��Ƅ�Q,��C.j'z\u�M^�`��4"#4$?N��+T����_h�j0W&��.�1p�`D�ų}�j�k���wo����Z�����
`��|vH�[N��H��W����U���X�.i)݌��凄��!�g \�"��'��Tu|�c���V��3:Wb��o(�0�û]�.rny|�:d����F�v�V��26GO�k�:s��p�.�ෂy�-;�e���ޫ���;����iiϙ=ndn��iXgƘ���3�򔶢��k+*9���zn�mi!{2Xw��_�ʟdgڝ!#]|:��P�wSf�쫎ȍ�M�OC[$�0�D]�܉���d���u Dn:�-gQ����٥��j	�rK{�՛lsp��;�X����;�횶�����Y���|���6L8������a��U����=�vT�z�A��c��K��%�G�>���r�D��K����s�.G��U�Kd��CF
U.T:6��-�y	�ǈ�ݜ1���s�j����J�u�P ��O�l&�LK��5� ��˛�L���s�l#����T��������;вnH�Qd���Y�g(j�Ң�[ >��ﲡQ�f��������((��_�s���^q��^ �lO�J�bND�TN�Q8;^j�\o9����\���+�3z�w��L`2��7)���O��V�t�|�8��%�{�,��{��M�[��ړ�U�Y���&&�Zq��w��g)�A�6�au���r�E_aLk��I�e�H�y�#���F+�.��"��,`���h��r��,!�2�pŞA��5wf�
N���."'Ǻ��	�]��{b��z�/:hl!�t���s�Bҗ$k��U��H�Kn`�s(NB�*j8��Hc�R�����D��V�Z�r�#�Pl9��H��ԃ��Z��k�((�H��Z�3�hT;�E?���WI·/���|�1Q���}c�Yq���S����a�l�� Q
iLȡ�F3#Z����!�=He;ygI�3#�i#��B�/
Φ=3$`��%7 cC�Datd�4�;�;��Ҝ��}+w���4J���}������9����[���wC�MJ��j�ݻ�	zs{����I�W����\�p�I��j�O��T�1����L$A�ӽV�(}����~u�Y�a��� �d3����#��cڔ�"��g����d�#j��To�;��Þ�:�鱡��U��'w"�&B�����6>J�(Iѣ�2���@�.'�Z��Ta��\���\)��Y�.����0�������D�[����J�`:_�ĉ��R"�&�
�e�C����ة��.��+�1+`>�%@���|�R��%j�i���TfW�7���6i�B��c�'r0����8)��x�S��&�x���<�%��7��ݛ��D\X�&͠�t�o�{.��<o���;�q��5��ٖi�#b��)�eI���A[Hm]uצ*oh_c�v�[��6�e���e*KS��+>�������r�6yt�Y��1@g���=;(��{�KDD�|�ό�t,U[NlT{�	�JX�md^1#��I�k���a\ܗ��s�J�2��X�9�),֖I�|==Cw��exQx}@�S��&���W��Wd��x�k����٩�o�t']j {UIBJ�b*4�E_�j���.-���f��B%�[����ƺ�-�Sy�{�L_��xM���1�&7��Y�����L�.�zk�<��t2M�����j�E��v���H/���k]ј:���\%��s��I�;��Y��uP�<T����f��7�:���3���0������*�MX��<_�C���03|��4�ҙD�Az��D��jnx�m�C3���N	u����F#Oz�v*i�,A����ȸ�ne��2{�������웶���2��v$�١qM�1�K�����a�-Yg�zW��ys@e̲�8G[Z6��.wgH�	�D�BNGI�R��Vl�>֮C�Q���L���9���{<�p��	��7���a
^��*���:cA����ok��>�>�]�ӀbƮ:� 'k'R�x�i��@%:��iECG�#e���>�4nTj��7�S�_]�N��)O��\������Dj�|�V��\��o��TiY3�a`YC���`����c:½��*�+I���W�/#��n��ԣ��uƠ0�<MX�|�l�fn�2�|�t/�8�j���'C'.3�Yo�8�n����\rۥ���E�3��MuM��n녹��3H�e��ʽ9*�b��c��fD���]&{+��ī3�k�ؠ��w�g��J�'a���+���v�������U��В�b���'F�,�Xn�:�#��<�w�2��#��7I�'\��vhTqA������]1�>v�,zOsYn�m띐��˒�T�oH�9y��vr��m�1���2�._@��婴�)Z.�CՕ,ݖKW~��W��&�U �Gv>���"��n{�X!M�ܾ�:����p)�r�iS�܍��8H��+�؍yá����^�J��܃ru�,nP�^r��&b�Z�;"r�u�d��@��2���� 5W@p�I˲O��g���z�;P(�:(MCN��e�p4CQo��_��t����x�gϳ[��|�e�-�e�f{O�ʬf�u�.6.K]�u�:U�g�0�*%�}
0Pȧ7�{oNK����G��$:�)��FxE-uÆ|�����t7]��7�Yc�y���o�L����}�~�48���	�K|����Z=�9ƫ]p
�MZ��&&�R�Gp[��K�p��K}8C�q4as�?$k��+iѾ�H�%_0��Q��q���W��!syln˛�$q/�{]�i�F���U��)����P#�_�u|;�t�k9F8��8>�D�����z����>�c|�u�%su�ô�`Q%{dq�P�XQ�7��{ۛ��ז���4�z�>{G[I}��D�7+6��+�j�_��I���'[}/ؠ<�_>�9�<�p��Z���-w-�|��y�~/����gnrI�up�λz��w���^8w�zfz�]���sT{r<�F�I��Z�ɝ�����W�WY�'\�d{$��S���B�r�w��,c�2yn�/:�5��͔0��*�3.�IRW&2w����p&u3�R�&:7e{401qʟdf�HB��_F׮�T[a!9�6�&S�;�h�������٪���CA��:��Cq�N���Q���3U���%T'G��鱡%j�s!U�Y�?����	�K�+$� �i܋�S���y{+����}W3Ig�.�A�V�^s�K&� Q�\Z��4�CSJ���D���.��F=\�=��5U�p�h7<���MyƯ�^9J�p��I"I�tNU�kmAC��P����U���@[u����"�)��z�M�jjaU�.�� �Œ\H�����B4R�wL�_eU�9�˝��a�E�r!����f����mL�����׽���N�
��
$��<����2;�ʁhSw�0����^}tь��p��8ut���Ɠwݩ%F��!pl�WC��I�=�`�DD���W�#�Y
~��E8t�8pc��3q�zu@UЫrjº����0V�^��P޶��л��SַO�5�2if�����5��"����.u�l|��s"�|_9\������tH�]t���xf	ܬ쿳�1����# ����ѽ�[�ܓz�ے�,�Ɵc���}[N�,Ȅ���� 4�`���T��J��?>	N�ceq�w�(�[�l��{�՘V����\[���s���8g�I�lԤl� �<!�EOl��}&�^�,���74��:H��v�%7#`8d�K�x��$�ha��te�ܒ����K^�bT���G!���+�Φ|fLl4��-��jh���')S���e�z^�ՙ >�g����[��:�鼃���W!rwr.d)����/)��)|��}>,>1_��aܱ��x"v}�G(����pŚ��oU1��;b���f�X�U���Fm�/Ɛ�i
�g��T�c���ƎT�h��3O*� Ɂ��t��}�Eڤ ���Zu�G�L���)}��V�~#�WƳQ,-��软HLt�oKԎ��8^́!7��X��e�tB�7�ڶoqC\�6OB3w4�3�.SP���Jٵ�����(dT�	N��Cf��jS,�t�RxE��*�1����;&����P0V�
��R�o%^ن�a��M�b��������r�.�X��L�kፎu�m���70��K�l�5)��K�����KN#�q�6P���BҀ0�u)^/�%��2`/\{�X�b��|gV�S}��d����ǰ�﫹V�S�b0W���Y�q����]||�:B.��K�����K���GN[b�"�u8R" d�w3�бUm9���q�[���bGE�Y7���Nl��T��\��"����zM��44�'�����ث���$*�b��QGҽ�^fF���"
�-��55����2�٭����;5 =�Ĕ&
�b+�0�@+"��d�8|�:��E���%x�;�t�q�[&k�D.y>)�r@�_m�]/2l*ŻNl����[�=�p.wJ���_-���]6a�l�r�`�����ꙑJd��PV�<����������y�G��ʡ��
Xv���S'-Yg�d�u�l�F��k�����J�ޭ� {踟?�U��4���]8�M9Y��C)�3�}O��-2R�ܵ}��*�NT�a#y�u���F���B���
���3�8�ј�@���8�p��ꙻ�˼ZW+���*N� �ۖ��ho���Z�N�����,n?<ûq����x��t�\�;����:��]~̾5��c��m���Lݭ>�7O	
m�JU�əm=0]�>�С�-N�VY��%���uӻ���3���]�8��k��[���8�:n���7�p������cD=��f�.8ku�q���Dđ����k��Ħ��7��Xo��u�͌*=����ɜ�1�nP�?-��z�T���R�hh�O���[/���eL=(cuZ�9�hqz���F�Lp��Sb��f�r�y��V�+�
PwU�~�<9�(�q��3�n��,�9�Ս쎭��{�	X�u�N�ꚫ���t�0�*�*�|�s�\��Y� ��22�w�.S;�2�V_A�m)o7�x���vX�nT頉��?XD->&qH�:����a��]Em�u9��y&O|f���l�\>Q��Z8 äwŕ��X�y�t x����{n�Z�\�;6�sc��ON@�,�{p���j�윭`�1�N��L*�͵��C�f�dv�T%�ڱf�jb���o�CRY|ph�6�T!��*��x� ��{=2zQJ�f�7�@p���g��l�3�;u�����H�N�l����A��sc��TիS���7 �z��0��[3�N�#<!k����f���0��ۓcu-
�P���g�8e��<�cV�Κ>G��yK�� 4�ɯ����˾#q��x-�\>�D�6�M�����Ev��+����.Ѫ�s�2�c��|��m��zoV�X�QN=���J��:�h�ۈ�[�A��H���\�Q���9;�$3�:�����ύ�]�Y�����uvr�w�"�tb�sN��L����\������G�hKV�E[�w��5M#�w6�'.��U{:���<��Ń9�w�^�Һ�L����j�q���Ṟ���۳��t�*�_60��}���U[���p�a�r-)W<���:c��E��W�0�{a�*w]$^��'��4���R&�x줏zZ4���=F��T�EK��� ��2���A�sE�%1ӧ*����WK!KT,Y���3ve� ���i|��J��r�Á��]��KGZ>��sso���M������vU�����_T�U.�z4�A��b��H��?o3��P�W��5k�pr�з|����_���X䃾���;9|Y�.���-��Yia��X�]��f�h3}�.A �of���'6�7͢��ܫ�#��y�e�(����h�ֱ�E�:-l��70��9�����U9���r���oM�8nF���3	U@���r�C�P=Y��)�J�i����-�y�rVo!l�R(i���,�v,ܮYעr�F�a�k(}�0�Y�����)(�wF��ʗ�n{<�7�)�#7#ɜ�Ѯv@.Nق�3�����{r?PR�od��$�b�Xw��z�4�_cC��^-����Ѓ�܅��x4�)c�m��k�S��;��_Gsq6��n�4�e�Vod��K�u�d�Jehf�ˮ���=�m��[�n�I^8ͼ[C3]���� ���h6���kO��ȆNm|{���Q�wf*;��������&fGj
C�u�H��u{V��[Yaְ��������`q�
U�ŝ톉x��0f�2���9������M�Nf�4�%�sW�s�����XvAQn��y�8�sg�M��ٝ�*TWk>�5�F=��쳗���I�++by?N�e:�oM��f��6���V�O��}�D!C�.����;��ب����J��3�#P���[Wo�mmm�+z �J^h4y�z�/�����ُMv�7S�N��+�=��i>wx�]��8��"�J+.ݽLE�u�B��� [�׼3x���J�9�z�<mY��(S&v-����2�BcB�d�{��"O]��3:'��~�f8�<�Vp��{��gm:�"�ba��M	7�hÓ8��t��T�1����{��c�sB�3@�vgo����o%�Wm�@��pv��k*�ɧ��m��3�ͺq$��d�y�0��ވ=��Yܭ��Uq�{
��!���kל8��y��xO3ǝ��{��z�K�ƿQw_���iU~�Qt�X"
("� X���"�@�)�V�QV0`��EUQF(�La��+*UX��*���*�����,e�+e(�B�m����5PX(2 �@����ZTV"���Ua����[T����T\L�1E��ŶIQH�PPUJ��U�E����Y*�jeF�Ԭ�Z�Ī1b�e�J��+��H�73"��A�8ʮZ�+"!r�UAdWPE`�Ҫ��fUAIB�H*2V��*AEk*6�2��c�TJ��h��"
-J�Ded�IiaDPU����DZ�R�8�\�b�X����S�%lR(�c*��D�EVQk�J-����s0�-Y(�LjH��(���J��Q-��)ULkR*�E�b��Q|��*
���{��׹>f1�q�c�E��6�\;z;]ՊY�wlǬ�Gl=k��]
������1��*������ޞ8{�/��Txd	� �i�H*��"�N!��6�ZB��ݦ�Y11 ���ݲo�M��}�LT����������'>�,��ĩ�>�u'�J�������<m�4��X����B#��� ��3��������g�����'��M̰Rq�Y�LV����̧���B�F���6�I�Ğ}����O��?9�$gRW�>kߺS�]JY[Y������	�6�Y�v�z�Ɍ�;��m�2\��;n�u
��}���I�
�����&��i��q��f2T�N�3fS�V�F^'��?$��~���<a=�	5�˜\t�����>��"��~� i�!�1�w�=CiX}9�h6���9����bc�L|�rN��V>z�;a��'�VM�Y��c>q ��'ɤ���&�8�aC����%<s�_rbc�<��0<��|�>���|5��|���_,�,�:��>9����Ă�0�}����bA{�jE:��<O'���!Y���hm�ɴ��g<�f�<C�s��3.��O!V��I	q@G�1&��@�q�����P8��Fd��?2T��0:�ߙ11P��rI�+�O�oE�HVu��9��N�'��Ǽ��O�Ŝg�{��`)/Կ~��Y��p�~qp��>�}�=����Vi�����I<LC�+>La����$gXh��?!������E�zɈxf`q+=d�g�<����N!YY.翻���B��3Z��{I�1�O=�����lm�,����[*�<��т"�"=���2T���g��1X:yg��m$�Ry�3�c1P��0�Ag��w2�g�AVo�����
��k\����'�fT�a_�>�m�hM�sՄ]7�:��ٿp�^�8���*A��'�װ�58ɴ������4�Y+P�,�f+'�tĜf8��_��Ձ�q'�����m ��y��u<a�1�9co�`��ξ^R��� >�#r��r�!Y�ٙ��bc&��ɦs�L�'����AT�%���>C��Ρ�g������i<dӌ��|<�q8ɉ��2ɉ>B�B���f�躉�>�21/���г�S]�P��q7`�+�C�&��.��~	�_��s�zt�߳�i�׻�q��>VO0a㾌v�q�㼦�yX1�"�r]�!݇/�=9�d�c�Վ)�{t6*��:Z|�v�"�������l�Vs���9xot��bj;��pY�x��#�Ƕ<>ː���
���0�&�i�Y����AI�{��:�r���eN���Oɏ{`c8�a��s}èx�P��e��P���=�R.'̘�	��o���{�ϼ�����&0���Ne��E&[? ����4��I>d�~��%~I���a15��Ԝ@6s܅N$�'�󔂇{ 6GG�� d:���WR.���)w�y��}���!�:�Щ?!P�i3���&?!Y�J°��?$뤚B����4񓉌<�����d��{��>d�K��'YY�%g���d �>�LQ��{�W7�g�CU�uw�>4�?$�~q&әG�!Y�<q�(m�M�q�<M0ǈbM�����S�k.�0-�*W�i���fa}�&r����ɴ�ϙ.��v=����C�}9ʅ9�w�U���jod�l��k'��u���{�6��W�LL�Cb����i�R�f�CZ�c����2�T�kE�Y*AC2����K���3��"DxG�&�	G��s��ǽ�r��#���N���CiϹ�oqd�wY5�
�z�d���4�.S��2m'�VT��yHT��>��L��ԝC)�M q㌩X,����8�2й����u%��z��/�����y��'��z��}/r��:�C�s�&$~C��&��i`|�i'�T�B�r��RuLz�a��XT��M�I�I4���! ���>��$�z~ңuJ9tZ��6�_�,�4�*u�:��2Wa�d:����1���i'�<��ꐬ�O���f���a�Oc�1�	�=N�f���O��6ln�l����ήJ�����p���116�Y�,����CI���fv��1 �����O��V~׹&Ӭ����aRu
�d�{�4x�Rq
���Mꐬ����d��Nk��^u���Y��WD!���">�Dz�x�R��}��L�(l�I�q1�'n�ɤ��'�<���=C
l3Xu&��?!�?}�C\�R/S���a�R��K��O1'P��l�gi�����lќe�������Jb�������&�=�v_ol�r�gg�
KE��AB���zxW����f��N��V$�p�x;�xk(�.M_V�|�+.����M(�d���7�ܵ�W{�%�[ػj����R;O�������>׻�W�{�X
N����d㚤�?k�Vx�P1��ghc�d�z�M��i�V��8����=�<�+>C���e=C��Ag[���3��ɬ���T�!s.���bG��З���o1L���p�d0>�N=<@�V���bu�'$�~�p�A^�8����'�m ��ɴ�?2T���SC&2���$�,�3�dI�x�:�~�+8�����͝�<�Z]��>�u~�������1���4�0�1�=C���4��(h����=`[d�k�6�=I�Y13��Y�,��<;�!�AT�<>���OP��=���@h��jb#�(D���#����^֍Z��<��w�>{'�>B�a��I�`):͜�m����i
����Y7l�x�C�gY*N>_u����P7�f�s�1�d�Mv��q:��sz��T����y�6���H>z�����?����u�.��8�����������dP���l� u+<a�i���LI�+��L��X6kܜCiY8�)=���6�P8�/���,VJ���N��q�V|w�M$�u1�o���]�ʽQy���ͺ�\�O��#�Ǻ �&�����6v���m�gP�ya�¡Rz�)��C-1��HJ�g�a�O������
�W�M���O���/�ԝO�%g׼�����*sp�Y��v|F��0G�q�������b�OS��s�`):�\|5a�����Xm�ϓ?}f3�11�<f̺H*Ȣ�i��x���~���8�&<d��<��Afvɛ�w�����Q�ezyo1]{3>��DH�� #��Ro���ğ�;��N�b��w�6��S�����p��i4�}g���ڰ��C�bg���VKl�~M&��2T5��,�%T����N�꿾�3ۢb����������,�>a���	��Af��r����Ӛ�JΤ��=C?�k(T��l���O4����hkvq�i8��d�k|�1+'�}A�~�躮�	�GW|� ��Ǽ`{�#!`��帓���aU�� �=O���h�������u<C�u1 �s'�=f��qO���a�
�}�u�Rz���oY1I}t�����^#���+�R%�6�sWlpvTp�J)��[���{=��Wvnc���-N����֩� �����m�N
ʾ�QxU��N��9��O]4�v�R�/����^������WJP���ߛn/3�Jj@��1�;{��H��������\��:gC,�H+�����bZ�}z��i�d���$�ld�+=�I:�����J�'�o��^$���O�u�I��Φ0m�g�:�Ȑ���L禰�7��{��G� |E`i>Cn�ٳ�M3�1���&�;�M}I�H.��z�{I�1�ߙ&�O�1Y�y��@�T�'���f�*N�_;�jM�+Cw�~�;ƫ��5I��GG�DC>�DO��^��>d�����x�S!�tŘ�U}a�9�1���ٚ�+8���0�Oɴ�͚�0�z��c��!�gRW�O=�(T�������ʚ��8h8S�����DCY�߻�7�dĞ~��++%��ĝB�d��o�,=Cl񒠡�n0X,�y��I���!��V���bT��7HV|��f��S7�~� �~����z]u~���"�G�>b"�{�V�Y�=���Ry�wA�x�Ɉ��tm�aS��u��� ��:��I4�I���&�L�'���eM|d�N!~��k�����>o��|��~�+>V��e8Ԟ�|�;�7��O�a��1>�����0����!�AVO&sZ:����{���=z�'ݰ�m �>�����OP���*x�r��1�/�'�}�GWp��|?y���.S1Y��H�u*q�Ι����<��o�O����!^2bg���m�d�ɳ����AgY/�wD�,�%W�]�4��P�z��܆��+=O�s<�����)��߿�~����|�$�bA�=O�6�C�c:�U�%|a塉�*�/S�L@�Wg�a��~Y�&!�zÈm�|3Lx	Y�~22)/_��`,��uhJ����9u�Az��Ƀ^X�3��� �A��0��*MEj���؂�fk��9��Z�zc%�MOS�#TK�t�����l�#�,�:ƫ��m�7ȈNr�Ϧ\ȑ��Jr:�f\��;��Tm���ɼ����;�K_)�o��}{�57��S�R
�5�{r���._.q��7�Wf�&�颇[��I���J��{罏W��q�����nʾ�5lg^�mu. ���-a����Ń��^7	�9�ӃD0��Bf��1�9Z:P$�(�L�'���*36�ЋV&�^]p�1��C,P�����e�q�e��	�<"�饺��.�ʭj'� 	����f�L�~��eV3a�^�ˍ��;�����<��}i��7�'�7V�\�gr�'����&$��E}�<��<"����>?z�������L�v��윑�@�)*�����G����0y�Q��#a���3�1q5�\�H��D�</e���%�;L��ȸ�k���Er�&!y�?$F�
�tz:�#�ڭo�쉙jq��{b;ToyC�(Z�A�A�\Ȇi�8\#�J�Rf����L���d�u'�*n4ْ�7QWƴS��7Nѽr��{_'�C���&Jn@֢{�c�v����c!V��7`0#�GPj��=����T;7�ZE�s�O+uPq ���7U'.	�����沴Ζ��B��D��S!ٸCR�&/vPw�C�>����-�x�#�~}S�\CzljA$ze̷r㍋�"k��g���B��ͺf�)\զ�va���!�Ԥ�`��9�>z|<���s�JԞ�m���	t�㖭qM�th�b-j텢��T5u�k�D]Ň����E�qR��9&�Q��:�c9H�����}o��oo����%(g��	
㛵��u��x[��� �Hز�R�������:��u��5�Fa�>��L%���A��_W�j�!	��O����T(%:(P�i�/p��nr��$K,E������t:��t��r�� �'uñ�=��R@ono�������ˠ�K,��s̽�לj����XjMŮ�H�ڔjcvp�=��'��i�ب�/�3�W*�R��`U�r���g��7)�������T�5���Hc�8�*R(��ϑ�X�
�k~9��g�3HN.v������0ك�Eb����]�׸�6���-���'�,����;�f�dw/��7{
z\\5*�"7B�H ݥ��������l�1��R��.J5>���AJ��#�KDu{bx�љ��Q�8�Zl]Z����8#r��n��n��ꐚ�2T�q���U���������N��@�Zs��|���b�^�u�o�g 6l9W}�x��V�N�ϋ]�k6��(�i���e�']�Q���u�%�0Zە6U�(K�r{�v�X�:��c��&VǪ���!챖7 �Y�*rԤz��О�ֲ?(p˥o��|p��[�����م�+H������p�W��7Ӣ��(7ɪ��`��W��zkqv�L����z��*�� x_P�S:7GJgG��[�q�pa�l�ʴ	�����1�~\ۭ�OVj�-{�m[>��oJ�n��j�?��k4���$9����}�)��Ugs-$j;���{6��� F�D��	�B����j�m��O
���+9/t 7�S�/4��te�mB����y�8��DL�Jt�G��U0h\�.�#��� ˫�~�=����Ȍj�Ȩn�h8s�kꘌNC3��f$N��XQ9@��n�B3���̚HÁS�\F�rn������<�1rp	.�g|�y��R�vg�V.�2z;��=��9��]ĨLMb\lTβx߲d	_'s�̲lQ�&�{t�9�.)S��2(4Ԩ������gFA?-�tpmJ���̰�l�MJe���2�*xFl�L$L���l�^�Ƚ�!�PY�ۆX�t�K�N��h%]|<޺�n"W�u��yȶE��H�����4�m�,P>������Cc�R���xL�f�d��#��骢��3��]pW�lV�\����ڸq���%9���x�3�e�Ҟ{���Eg��3�D���Ԡ\^'xw���<�5<3j�Z���ᙑѕ�����:�sW��q� ��Էs!��r:u+��.7����E����x��<�{xL!�d����������(����`>(
��H��;p���U�*j����6v�(�G4��n���!�ײB��fF%U�h��� >����VX��X�WO�=�=��]���F�h���<���!(�;��!���nH����eÚFQ ���Niq�E��Qy�R����iˢ'��ȡⷧ��*vٌ6Z8�c6�'ts�Y�z�Ε]D�ާ3�d8����?,$O�y�п��C�K�^����E���z����
����uՊ5T��g��^<��q8�U��٧H��-��iϳ_O���=8�d���u)ʹ(��:�+�<���~N`��(�`��a��t�^a�x��Byt�{���!;��)��M�T!5��MMIXX
�nXZɡ���OK'��~ZFr���@0�:��<�jsx�⸸IV	�Wg�ޓw�\����62��B�� �q��
�hTq���ËZ��:o۳̭���􇇢�n������c��s�Nv�.l�Ǖ+*��wDO�[vF&�bڼ���R��\C����jh��ԨB�+;e��y�ubIՅ@��_OR�=z �FՔ�^P���}�c�Rɥ����e�_��|�I��o9SV����	ʱO4\�9z?xU[�Rig���Xx��k�jǢn��#�����4��_���+�t����r��z���l+�ｮ
�\�5®ҳ\@��
���ӑR�0Cc��fB,�o����̅{�o�����˟�v�?���X^[Xd<O��k��$v�_m�t@�	��w�To�%�G�wd�1�Y0���8'N�K��bn�;��.T\I��G|Y\��\B�/ߦZC3p�����ppH(�7w
9�¾!���d)}N6�7Y"�OA'1����:@��B�to^�<D�F�C��^)��|�&�+|s椲���m��@	G�)��U�7n�!uYr��s�.6O���37e#����r��i�0%��IҨN�T�����_U�g���ˣ�����P*O� w$\�ZH��g���g�TB�\8d:j�.�s�!��]������7kt��:TK>�F= ��13κ���p{
c"��m`������&T܃g5�~r뉋�c&������C���AZ��N�u��M���Di<]7]��E���f�#g�66Z��
��^�Ke��-����ʋ-M�g���wW�ށ�����{D��|���)�f�D��֤��6��mZ���i�9]֓��^5R�;��ٳV��Qk27F ��D�G����n5,���*��^�1�hoPd�n���8����r+uq?/��]H����n���bT�#9���7�^��~C�������V��2Sr�.�q�$��U���l�]>q64�;�!C�1V����¼��׻U��7�ZE�2z���s7�<z�G����0z��1�@rW�PUc�U�6&�zMJ�\=1P�ťO�`�c�^T���Y�ī�J~���k��=�j�&���ݚ��{^`���#��*>�$ѫ;j(��d[֕�S�jxe�Fq:�c���r��� ��q9���/��?���<Q�׶b�wc\���q8� L[i䌥0�!����*��d���1QE�\��u�S�UH[M�LL�ˣ�_7�Tk�\�)�����K,����^�^q����Caa�7���	��\�Y��=���I�|L�%��#|�J��"+��k�9���m�ee7tX��z6.�痵�ZϪ��e�DuEh
�}�]t�}}�Q�s%s�>����}^����nN�\�Η*ܫMw9�g%gȦ��К(Ķ��dq��h��'�`��/9�&��ꦌ�Ȥ7[ӲY��"�xH�!�_L�"�c4���E$�:]���rP�����&��N�kv�V���kt��v�.��a�r*y�(�j�2XI|��=�����т�p���-��{p�꼄��tv�|���q,�v�X;}�8�Z*�*���m#[R#�`@P��>:�L��Q��Eb��P5�̞[��oGw+$��� ӛtg����e�����[��z��]�˙�aVkz�K}��b[�*�׎�ۙ뜷J�8�˔.{�5MΞ��<�}Q�����қ�$ζ_oʋ�@��w�+�|p-҅�+U�Ul7�q2�g�2���Zڲ!y�Sn��hHjRG.ĉ�g����dw��c��+��{RM}nn��U㝯8�ڮ�T=aF!<w�Y�;DR��%qtM�Z���*�k�	38E�Ehi�[�3ϼ��/pry�;�aV<��x�3�!F�Y˲��;�jiE�/$y6·I�#�\��i�Қ�ʝ6��<�h���v�!{6��"��0tǧ���*��S��}��uX�SC��X���+�n�lf�AS]�//��n�T�gBȤ�t�X�IRm��F���mϭݕ�?�(;��k-vp#�5�{�[��LNT�ک��W�wfnM�����T?A8=���C1p�É�%��ήg(d���ג0�$��WMj�%��i����-p��;�V��*q���]sl���^��G������
�3�Ӭ��j���nlL3��g�CD���]|ɱj�c�_Tʉ�:�mw4\;����=�H�~�5�3�v�}��5���Uu��	I�B���-��]��� �;��3�7�f"��*����F��5��_J]`�3�`�K:1D��:of�sTN�n���m`|�g9tq-���7w�����!LۻKe�x#�k����89MP7�i�I+J+t��C�;h�d��]�NRio���O��J�=jp�d�j��KY<%�VX��>�ͥ���@snQ����^�7V�	���c��ޝD��U�mӵ4HТ�ð!�i���z�T�utn�����c`�Vn��D�	��B���d�]ӛ�x+�_uN�qҬ�(!�{�>h\yA�n�
w��U���q�V�U�}�d�.�]���2�z���r>˳j(<�{˧{ϫͫ����2�Ok������CͰ3Z�s�XNzb�+,&]�7ڑq�\4������o����͙@$��2��:U���n���8�S��ུ�f��X��{1�J%Z.�V��0�qA����-ݺ����xϮ��­�__a[�&��1��f���s�g�|�vV���d��tls�\6�3zu&t:&1�N
b��rQ" ƫ"Ƞ�����X�"�LX�T�DQ���#Z��-��q*LJ�m�"�Uem��X�E,�UTQV##2�A��IR�UU�
��AQQb�E"��Um���iEjU$T`(�DX,Qa,�DX�������CT��
��,��ذ�,� �9b¢��RV(��L�ff���EX����)�QI�#l%�J" ���SH9H�RV�KV(%��H�ƴE �H�",��b�EU�R)R
T�[��Qa�X������b�,���Q�ڐQER#"��
T��*U@R���lIYRT��T��@ET� �,XT���TU$X�l�
ɌYm%EAE��bc!�~���]���O�ܼ��C������������t�e��	�
<��fv�yg(e�ţ��v^f���k�}����SϪ�ݞ��q-h`�F{r�o��?T
Ã$�D@L��E�L�GL��p��:/5R�M񪀉�ܵ|����C��h�D>����p8T���.J4>��P`�ZH<8�q��-�e�	=^����,��S��n��nv0�$���钦��!��c�p�і1��5���R�2{���O��o	�'=�Ù���s���84 �$�<k�e_"��T�WF;պY0o"�W��3cxuݩ�A��s6�}7��;�(ċ繱/��U��2(@D�u`�SH�(v����i��CP_��vd��¾Z�M$&�q8H��u5V��YD�<N������iվ�Xr���pxej��ۑD�n�B���=j�$���_�ԟ��i��WѠ]Z�|�Z��9��e�ٽS��Q��TXr&��Es��uL��a�,\7T�^'A��,/Ɛ_Vz4)��n��.�t�;��˹��7:l=��yUڋ���.��e����w�;��ώ��o=��E�A�[.�E�]ykI�8���@�h�:h��tR=�5��E-^��k4�]hǡ�[K/V3�Mms���2�&�[�^�Lrt|���h>g�78����x]n��-�wuu����[j����uAC	X!�����w��`�ّe=�7��!o��3��ʪ����w�c�d��zvV����x� d_5l�I�L��s[W�_Ni}w�:cQ�\�&�MR��hw��J)�3ѐO��6��ѕ*�S�2±�ECR�`�.�܌U�U�S��u��F��Sz����Y\#�V4|)��Z�Q�~e�� ��� nNԮ��t,m�y-��N�_�ޑ]�S�y�|~�Ek�-~[vA:�$�|�KU!_r�Gf�����z3��aO(�������!I�COz��=<�V��9"�]�O'�J��c;�UQz~��<9�3�HX{�R6�U|�'���0�<�n�N�W��XYƻ�L0nE��#��J3M���J2��P�a���"7�x�F[�F{#�%�F��w:,�R��T�8��c!}K|�
��qњ{6v3}��dXo%�d� �7ѥ�����g�z���u\f+�d��O�4�G>�ʡ����C�c]L �I˜�*e'ð<ĸ�Å�3IW^Q�\��q8�	V���W�#�ȷi�+u����/I�۞�"��5׾��i�&'PRR�F/�n�V���T�/��:l�L
�Rõ�r��渭���S��O�j
���|E������e���`�C�s��������9���Wt�n��Ӧ��;o����B�7EU�X#�')]��m����UA�T�,Λ������_4����X����f��(��d-6^TTD��c��>UO�VV9�ԭ�������h���a`+�健�ڱA��OK'������u��K=�R�^��]���=�dU�z��tè`�����@j�H};�
�ğ����CT����k�{�(D
�z\4"�΄ʎ�Z��:ovy�ḹy���[uX�f���ՑO0�	��z�c���B��6-�R�.�㐚�G�N�&н�����Ç.C�l*�yB�[K|Z��[���ۊk�N����@7tUp��x]l�0���0ƕ�gr�0�ӭ8*�2V����o����:�yma��}%�v��^�'K&����p�I3}�K�=��J<��LRs��ӗ:]l8�u���ܴj�p���;��=�.BwZ�mH]�qW�H�-a�_rC�Ѯ��Y=�L��T�d�h�Ɍ�,�T�����=��I�2��S�X�)��H�ʞ�IgD`�/b��p�x2�y�L�e��=+cNs,��H�mQ����PYn��/Zw�
i���ɤ{��������1�*/��ۯ����BҸ�����j�k9�5��l�}����3�-U�{��k��%ս��a�³���r��ʛ��{���מ�6�2�I�����������r{�6ܞ�_��������f��G�8˧?K�,p�p��H�����W\�bbܔ�s����頴�nǅs/h��ϙ	�$:ķܳ��R��e�7l�q3	��V����ɾ����Z:1�]���q<n�����&Io��6*��(��Nt[�Y��;=�6�n�_$ա�9t���c&�jpJ�D!ˊ����xsr6�7��w�����\z���-h�e�d�n���0G ��T��O®䵮H<��!��p=j��,������/T��QC6{J����Ϩ�.�d�^��#]��(��E��J��o�y9�׆to%XIF���Z)�9�{������0�g���o4���9�'�"�wY�������9�#���*̬4*Wl
�p����Qo:�~y���!�ʷ����R����s��5�ê2�P֦Q��n��|����� OFA�����dԃIwj캙�Q�ݠ�y�g8�9�Gk���c2}>	��Zx��2:���2�J�B��DxN#Μ�3ڣ��Sw�P�u���|X�p,|����9��XsF �e��]VRw�t>��%�BX6{����5��ړGx��˪�xS�R��\��C;�%�;O3kF R��7��.S�Η�������������g#���ο�_W��F�&�E>���ei,��ϝ�qJa�o��S�J�s�S��V�!��K�9J��Y�9#W��l˅�X3�������2]Dr%�Mk�e�&��P/H�N��lɜx��t�f�fj�j��8�$�'�]�t������
ʾ����?9���pܦP��u�9o6R�U�m}���tAf��$�![U�L֩<wÔ���֜y\W�F�n�<36��*���6�l���p�������;�HJԫ�ʾ����ypc��K2�s\�]��������'���^U��uϝt������Ep��{V-PZ��������q�����9u9�S��%=�#jR\��ʭz�D{��.p�7��c�`|/��qJe������'Is:!��M���h���ՎV�-��gz���� "z��R��`��xEGT�:7GJf7��Ki�p��b��2^p����)=�ۏԷ�`�����Q����Հ�HȲ�i��zV�Nd5}�tf>^�{��n�.���4g+wvx���}��(:�h��a+@�Vl���M��B�Sz~꽾m��roX'��z=h@M_�V���vS6�۩a�]YD�#��`��
�����L�iǋo�j�B���o7��)v�ż/��{�;I�-�r�AL���UVt�/B����P��P�5*����S¯��8�#�����S�u��8s����뻑a2�e�68��c:4�����nPY��Eyݔ��z6n�����F.�C�XX�ULE���fx�@��f$N��XQ9�2nWj��o���~�D��j��~�����d�{-���qރ:e�ϊ������	�_@-!�_}��� �Ĵ_���ܘn�]��Ī����ߗ>���x3^��r9[N�5n�*;�,�T~1�S�M�@L�^��nL�:6�Pjr6e�cf�jS,���(SbA8�"��ٵ�NYO�.��H����p�k��G@�<%��:Y�q�L{M�`t��v&�v���Gt������C�7)��u���9�*!vT����>>�d��B�*��3V�瓘p�����Ы���ʡ	���|!jч���	S��B����$� g¦��a�����M�ķ�N�U;��U��x}^=�����Q���fb�W7�?�d��Kֲ#e���
������g�0��Z�X�6�e�s������ݧ���Ǥ<U���e��@�m�Ov�ͳ��Abm-�a�\�TzgY���	��ã��mJ��q��5ÀJ�*���h��!p�`�F1�U�ޕ���^�87���ָ����"*g�Iq'$t�L�[V7�Rj�l�=���1�r�#��e+k��l:�N��I�v�q2� q�䍉J��S(F|�4���b�m��se��gEI٘ڣj�0ݥ�I��;�D��31^��(���/�<�h]r�cr�Þa��h���u}�%�f�ҎU��,5)�g�����s@=\N0�o��5uH��*�*qC�h��Л����-�;�����T�x�9�W�
sGUc/�#�h�+�?W�n�p�Spz�ޣ:cFS�ۆ"�S�cUro�, �|ܰ4�[V(;?	��d���;��(���;��:��?uƇ8w��z�E�p�Ɗ��pBI�a��*^�mC���zr�<C����Kh�1h�-}�(������L�ү�
�zP�굕��̓��O>��\�*��<�Vi���X|M[�\<��w��tx������Ʋ�
�fmk���B�N#�M���1Q�*t�0eD�$C⃭��y��j�ǷQYw~E��4��;��Y�<�v��S�݃����*պ�f�i�׵|.7 f)&��t�2���w��	,�Z������S=��oA'w�����U�=�b�t��w����:���.R���8	B{c{j(��D*��6}��G�tg.ni��6��i����g�)W٦�,�����Ҿ���|��pu����܎����O#��_�[$U�M��t�j�[6���7L]$�w%��X��o49�j�Kn��C���"AF�����CD0���&b�c�鷃uK�+G�'Fw+��^��&�R�C�q�HC�b��,P�ʞ���s���apL�ЏV�<�=�ׇ��0��k
��f�����(	���΂����k.��=�8`S�L�fq�O.�(�����1o	IҮ3�T9�!D���;��&L-$i<��D#<!�����eģ5wn'���R�P�W5���q��n��4'J,�x�� �w��+'�h�Wy�n@�;%y��� Ӯ��j�w`�MZ�Df0"Z6�Q<as�?$ut���0����x�Q�n�w)������}���0���p-�`X
!U)3h#8]���`�n�=��EY5@M>���Q�v#x����(o=^C�P1K�Y2P�����l����{<��	��2���]<%�
�_L�-ڥ���ى ���x�f�]�CZ�\n�X����wS�N�h�\]����,����%��%4TY�����`!��v��f�ʕ��}�TW�g,���2W�8*��������k���Ϯ/^����B$�r0�ѹ��ʝ��}��1��v���ovru���9�be��ˊ��|�~�l���T;���v�	��xlg�j����A�Ckj�r7"ʅ8.�>��N�����Օb���M�0�9��vG����h�H�����*�7���68�޴ �s Y�2�ֲ5����fO�&�ai�n�e����Q��#���������Ǯ�u��H`	����2"��d�b-l�CJ��Ŏ��X)�zz[Y[�בx9]6�JE�t9M**�@|p���%�Mk�e�y5�HWu����a���]�V�Ȑ�ܖ.Ԓb`�	�
�U:��z�
�u�^�t�"�&7�J_Q��u��ecy�m��u{`VpQ�ꟑ�p
����n��<g�r��/�K
ߋ���R���߷���D3�� ���g��4�Nў���̋��a#C:�������5ar��g+AO՛}K��O���l���85
�B�%C�2��fB\iٱ���9Y<^�-�y���k�d�O�ًaMV�}�%C���\�@zg+ks��������w�Rr^b�+�0���kf#����{�����6V/�dƺ�hq���7L{��=Z6=���m�����s���
83�N�� ��O&6[�3����������9u:�>;��M��#\�
�<���A�U��ivq��h�6�=�����V蟳�|��}_$�#�gD6q��p�h
��ꍧ{�w�s� �$�. ��7L Bg�TuJ�w�ҙ��b]NKf4B3�157�e���ZT�"m­~sJfE#L���w�}*a�P�1�VNd's ^*��qKc�WW$���޴d�@�Ң,�2Kx��Eϲ���uچE�9��ܚ�i�(�J�y�g��������XL�3_Cr�(}��A��jL.��~�M���@ŗ�.;�J��w�۞������XX�2�w؝g� ��c��12��v�`�:�vmu�><��Me�r*f4F�_nڶ3�C�2��y��R�Uqݪ�\�U��ؤ�������ŀ٦NB�+��Ɇ�[�x� b����e��D.8��X��ak�t�s�tE����hB�+�Rp����׍�Ms��wP�^���	��3�5�T��j�,bu�!���"R�喪q >W׷}Wϝtj�U�l+nZ��Y���J�9�1���;���e���H���Z �7F��j����;IJ�i.qӠ׹ӓ��m�&7&��0�!��I��U�W.һ�v���L����B��7���fcVy}�L��IJ�gʩgj���Hc�{R���B�O��Cx���BtEh��ej���+�bS�)^�TB�-�7�|ff��	Sr�{.��t0�m
.�;9Ӂ9}/ ��ˆ�6�G�b����q��m�"�s���	�nf�W(;��GE��v�T\�������h���x�]��WC��n�w�m��smf�r��(L�
P��y�M�{Qv1��-|͘�?b�H�3��Cw��{U��l�SŲ�ՙ�����c��E[o8PU�/U�޳��2�h�B3u[4���#��޺�C	MJ���=sCu@e�j�������Ji��%5ɛ׺�;<E����qܶd�ssU��b������Vc�
�;1�����$uϨ)���r��u,�6s��#M^��V�y���b���d����1�j�܆��ٽ0j��m����+���uT[o��V���ba�wGR'�w�"6�8E�������-�8���nۢ61�Z� �{�;�dQ̻��Z�ú,U�1Q7�kmG��
��m�[�.ݓ4�6M���Jm2m�� ��7W�Mw}�Hc�R����C�x��t�u��. E��K�ș�/�]k�&*N�0�������i��8fwr�B {V��-<Y�Ҭ��o��;�Mb�=���+z+h���n��y6�ɀ�
2�b$_�x����{M���`�n�R/���m�,�=��"�g(����5�Ϻ���u��}8�t4�s6�NJ��ᤗv����S�	�v5�;oJb��3=���0x�k���']�)�lt&�%�I�4��љ�{���T�{w��n[��ݤf�xy�yQ^�q��o$׮�OZN< �nz���b�^���dĒ��!a�6�P��v��VWb�#p�z�.�
.�����f!��NNn��ɘ:�����2�N�	6��a�-�Dk�n�vcs�Lа��5�!p$بe��!�w,S� 9Vı���]](�W�8�͊�.�ǜ~Q���Vf摝v��Ϯ�}�]��ݐW�0��3Sgve�+���Iv*���mks�9݃���m�M���F쓇h��("5܎���C�>[]y,��l8����1�����L5��m���j�HA�v��>޵�m��n�#��v]�AJ�w��ke����c+c�E�����ٽ���B�nhC�]��^>�����c�g8�x@[X��2�_�5���SQ/�mW�>�88�����U�n��]��N�U���gwל?������,�ṱwF3���s��py��{n�_�QUUE��ʶ��PU� ��
�b0U��eecZ�
���ֈ��*ł�DAUX�TEh.�Qk2�U`e��ImŬZ��%��b,D�IU��0R*"0��bAKs(�D�*��Q"�-�
!Q�3

DWb*�
�
��(,Ym�*�mR��Fڊ��DR*���T��mEk�A-�c(�%VB�@PYXUQ`�1"�*Ҫ���R�2F�,�2�a�1���U��X1 ���m**"�PR��)��Q*J��ĬX#*�*���G)(��B�m%B�X���UJ�Leb8�UImZ�r�b1b�J�(,PY*J���
A`T*g���>��W-�r����e���6���խرyV&P�����&�w58,y�LȬ.�o˻zR5��>����;WXe���Ν����=~���+H�Y�p�B�@:P߅Ib*'UR�XlH��u�ܻ����Uv�?ޯDPL:���3�N�X3zE۩�$��*���vnN"�^K�۾�$z�\�1Q�r�P:�kk!�НɎ���¥N����Q�U���Y.yjAw(�{-���8B��^F��,�z~	K���ar�qO2׻w�})%��:+��Sfy�d �ԞL1�)l��=\�	@�;��7�&�P
��&�iO����3�g_[m	�'�?$�U�G�TD�U�2�B0!�V��ޅN�#z�)@Y��S��;sV^L�Ә��T̊�2R�'�H#���W*�7 )a�g���Fʆ��o(�̩S��l!�Z��l����T�(�a*�@��:�py��/����f�v�K5{;�)�W�T����R�h9`sȯ�����B�fTa[ۧ7�FpͻM�����b�C��b'��Bj�N C�nX^BڱA��rs�2c��ز�F^=$k��%\΍�������*�z6 MsMS�ň#u7Z���1�D,vx�f��w��gj�/q�L�/{�����27օXac0�v�.�˩��L��d�m�լ��ܪ: D�7���f<�9�2x���{������ˮn'�6#���G 15�oT�Ǹ��&�r�&>���=��7�w�>�Ԓ��˱��r���3o�BnP�?"l1ss�J�3�g�Ƈey�����O D_F�E�}[��1� ye^�ha�j���c��w�h�2j�3�I}�Fmm�b�K�t<�A�R���F�S\�/-�W
�Kheu��:�+K9�o��s[);���ʻ;��8	��31u�נ�l�]^�(u�E�ÁK@�BXۑ1��"�.����r&L�LF��ҏ "ۓ��s��8�y���V��i䳕Lޤ*,��\�^�&'Q\�x�r=>�H7��v�k��� 8�O�B��o^���*��y1+o%�{50�T&�W�N4�	��]!^)��|�&�r�ŢYxm[N^c�x�c��K��sx(���n(b��e@�x�t�P���f��G�S8�;u��㫫[��b�Eg<V���#�����;�Rt�8���!EIF�����F�	�r��~kr�ۙ �X�=V5D�:p:8h�\-�v��xI
s����T�ҹ�:4f�n���C<s���)�4����,>Vqu�m�Կ�������ݻ����_!��t���1����/���w�6���t�M>���-�oL�0��u�&:�c�{������|7�^�� �+cb��/&o���t�4'J�K>�"8�U�'�LQg�`���S�2��[E�jFGe�圁��ϗE�.���c&�������!��5�R�y� ,�B��z�zLO�6�5Oq��_0�5�Q��*�Knx��`XЦ+^���!܆Z�r��O%&_�,�O���|�^U� j5���l����z�5PEE��L�JD�V��j�t��vXmeئb�3�L#�G%�Ņ�=��]l^F�=+�����`�[��s��<����'�:�v�e��6P�"�
Gj"�L�f�]���Oo��cԙ�sɜ�U�,ظp�n�ذ3�t�>��](����l�(�����a�3�Y�%��P�և!Զ�6�`6���c�FY�g!:�
3ٶ�M��|w,��%jc2?j���.Q2BS��VTh��e2Q�6�����W���yg�c�d+�ik&�Gŭ���,��C����鞳Fr�Z�TUl���2]DtC,��{N���)V�5Unn{-��w��j�.cJ�sHP%k��1\y6��^�y{	�T����v'��r柌yx=P�&�s�tC�g]�F��\}����Eۥ��Is+�]�&���C}\����hS����:'��p�q��{qf[��M轞�����  <���5ξ��k��:Ц(����$Ңts	`�U��T�+z�
�u�B1ӂ.cY��grrg\f�M��9��y-���٠��F��t�E) �(B�]t�E�QE�n���N�n�%I���S%������:C3�"��l�}B*č,��g�'�w|��e�,;�<�; >�[�Qű������XD�v
�x��d����[�n*Ugت8,�/aSY� Ϊ��A�g����lP�z� 顰������F��H1��U�4"��F�n�Rie�x������yփceq{�	�8���Rt�d��ʇ;XFm�s*Ყ��Y�˫t
4 ��<����7�g�TuJ�tt�n�1��[��׮��������k�	�a��i+!ր�>IUƆR�����\��'�R�WaI_�Yl�C��9b���ъi;2n��v� ��q�����h[�ކ���� �n�j�=�;r,�6�7]W�ruR#�2ۖ��c�}��j�Zގ��U�~�[Qմ<���9L��U��1ԕ���[!���e���rٛ�&T��@��w�̮�s�����r���%��x(��r��c6>�L�qp�Z�0��0<�n�����R����w�-\�\�-�=�;LuRGb��yg��<�������N�Q��]nw(B��c��ÎULE�t�ϢX�t��ču2 s#0�ӂR�lM��HI~��ʇq5���1�0g�em1��2�������vnh[[0\y�'w����ү�'�DuZ��uD�,�X�Iܘo��'��� J���X��e�Gz���bS5��싟r�A{����Lm]q�g� �D�Bg�ڧgFT�NF̰���eoe/��2�M�a^Ժ�'	c;'	�ܗK'��MX`ٿ�p�k+�`�<)�D���Һ��)��R,����[�HE�)��<#9�\�4 ̓�e�=zC��?Z}�=�꫍��`�P��uƶ�,�#���0�6��I�r������WG�ܯ<� g�}�|x�L�UPYb���)vw��cm����z�hwΛ�ީw�65�<����$� �!�SEi�����ct�>�<��P��p܎�n�p���T���yuo8TY�,7�bӚfht�:����|*4�e�o��p�aK�O�(�d����ݵft��xR8��,APjJ��g��r����g�hڣ`�lL�!6�q�R�#&�(��d����9'V}E��|up�Ql��j�j���<�u:���L��#�8+��1�ho1�UmhK!�
�)�__n�-��F��w��b�� xH�����������۝�a̋�^mМs,�q'�~ޡ����S�W��}t�Ȟ��x2*/R�X�C�eB}l!�9j�8�J�u�"�@��NЙ�v'��}صoK�uv�.�I}ŋx=�#��L;�Z�1�~K������E}`�0DpD�����5�.:úд����e!��@���8�ϩIB� !Pܰ4�[V5�kJo)�*0�=2g��S���[���}а�4���H�u)������ӟjt�7���)�e�y
r��p}�>WT*!������`��4��k��;�����m��H����ۚPGa�o���Ϊ-��HŃf�J&2� �d�V��~���~!��i[��]����[�aŇN�������Q�ck4�g1�\*�-]z����oc�@*i�C�d�fNH<0���v���I;�\�l���Y�n7���p��_j�x3���}a��A|C�%l�9��>�-(�nLW��nw N�R�aƔ��*ůa%�ƿ+���smm���8f+4�49�����Ur�vz�qyE#1P��3���l���1<3�kb[��]б�]��z�N�|JL��נ�i�9}`pԦ��a�4+b{Kw֌���9a�����tޘ�X�7����j�u�K�7���������n��Fz.Y'I2��J���J�t���,{P���)�L��:����7�k���&'�,v�P�B�!�F-�(J�OL�U�mb=s��3���
WR��ڗ�)p�Ǡ �<��)��UZ�*7��Z6\��ͼ)]Lץ��ۥ�|ԝ(c?^ØBI(�A��.���\��+����,7��|q�@s)r�cL�
llXt�y3x\e��t�n����Ҍz�.*����t:�YGi��L9�[F��0���q���ɫC!ˤL_��M58�Q3�I2���U:3:��/��B%���0�q;��V�|v����|h^�N��`�f��T�\���l���<��U]%?,'��#x�:�G��s����3���o����U]�k��(1����XW2Q��o�� �L�5WN���󊎼U�|��jp��ghT:T$��{���#hvG��e�oZZE�s�O!n�9+��xzʳ+����eV9�U�6;�u��;d�t|y���.­ɝ�D����n�X6ݝ�qM���d޼��	ZA��k=W/5��i��*�E�����s�'9�ĭ�At2��qN�g'�GS�Y|�3��GE���*����Qw����w�(��xG������ҭk��f��n��h`c����N���k��VU��<���'1���/r�C�I�%�æ����'���ր���e�Fr��S�- ����1�����m�<1��]���e��_WVTh$�J�!�'��Hȥ0�6X�[6Ү�k;�����m��y�ɪR)�1_Qd���8�Z�TW�l���d���	e�Z�}����23��+N>Z�iϰS��5y>��#bUO"M"ty���썺��RDlbu��x���y��4R�Y��3�Q�a��z�6��+��M�"2��pc{�8u
�=�FZ����I�7=8l��+�!�Ч����m=�6�H�`t��ӥ��:�M'���\\Y�W��-�ғˆ���|3�q�R��Kt�J�m��:�(k+�X,��a��:�@�{5�/uy�{���"���.I��Q#��fԌ<�T�u�dp㔆	KE\�Ψ��2�I���}c:fb^+�Gs!;X����FC�d�)����<�@٭����U�>7��^]�u���0Em
����0i'BW����u2 ���)�8��$��McT�V:��S�P�)+�&��)b`�oz6�ֻ��.�֣��e�]s���� Q��;��1�V�mǢ#?q�JU��~)�����ɽ�k�-�j��_�� ��v����G��o�W�8õ�T�g�Cf�P:�rmvU#9�K�����]Frn�T�u�O���&|��w �����6~��;;�t,ֶ��6��u�S��ڸ�[�m`�tW1�Cn3h�|�O������Sh�.�u�*v��n���Ci���)e[@oK�|�:�mFPjdE���P���K�]���.o֗h��~�v�N�Y=�)���|�g��.�zN��̥Ȫ85��$}�C\]ä#���V��ѨY�1��Nd�{�z�u���x.
�f�byv>��WN��k�� �6��b���b4��<�Tֻ�]óJ�
��|�)|�	�^�Քn�]h�};��:�]��^�0Z�&����=&�9=.�[q��րo��/^��@�Gg�0h���<n�i�8I�ί��|J��	����2�Ҡ����?R7�Mm�������Jz�Y�Ns/EDk֎j�F��ι�Z�l�ǋ���[�V�6,��e1�;j����3@��N���֪v�����w$�|�Mv����}���{��ek}�����-V���+`sx�5o��{f�������P��v5���a����|�6�W���Of�����[p�-�Bz���9��[橙��Vm��B���&+�)+[[�><��Uc�!N��Q�i����;�u|�e����,�^��d�;l;�WJ����8�˪�{)��sZ�wCl�9f~D.���CA���5ү3f��Eh��J����7�=��\��/a�3n9;�<D��#]�'�����2�j����G0k�h	\�[�����5�I��>�ZrG.njM�	��Z^�|��+5fz��ANZ�.������F�ӄk��kl���3�ubݷ�xym�F$�xne<�9����Œ����^S{��{ާE��&�w��~ރ<̬�c�_	��|Ҟ�Z�F�����;3qa�WK��E���ZjD��K�p���#g�QٯEޢg��CM6M�����A�t��L����fP�8����hm�.��d�ul��Hގ�y+�^+"ާ]�5s�*Ng[|����q6���������[���{�pGw,�����W�I�vI���9�\�6����T�y�q�@��ܕ�v���m�ݰ���p����C�Ѝ�8>ΨnT��}s�*7�.z��gpZ'*�F�sd۝�Q��t������<kؒ��l�5D��6�oA��ʦ��Gbk��u��wEH3~f�;{rˢ�g"�h.i��;�dQ�E�ɓB��]"���`��5gv�84�{jV����jH�Yb�:w�����J���)��Ӽ�[�㗆����|����S6�ِ�O����N�.�f�9��k54��vXCh�2���D�C�+r�0X�.eY��36���;%bZ
a�f�u���釓w����aL�b���5�d�m��q٫o��Go{^�#6U��lEJ^H�&��*!��kZ�ͤX{�`���G4^���ꙧ�T�I��V& ̃9�u1cMf�l���ڻ�è���]�$����p��tE,�u��K�a�t�y�wݳ�bͼ���<���<Ѽ|�^�(ݸ�p�9H��]<ǸeJ��������f#uX�HǬ��oT3�N�����R�N��x%k"=��Ӭ+Mfv��L_P�{QkSGM�D���q��jRQq�3�b}:���2�E�V�S�� ��է
�Y5[������ta�:e��j�Q���-c{��}���$#q9�!�����u�NeZ�+C�D����$$���*I�~m���l����!� �r���]���+��(���Ո�K���u�,#��]�S�6�3N��)H.��Yr�V�q'�	���ٰ�w/�2z`�t��E����{�щ��g���RM�3��+�[#3{X�8���v?B׳��E�Q���T�j;�/=�h����l3�_-�t��%[�V̥o�.2�x5�4�ũ��ܥ�M='Щĝ�7�7	��Z�n'}�jܱ���H9`��h�kE������
��-��V�A�ƹ�F�ݯMЫ��e���]����h�诼t-xM��t�Q�$Z�;��{i+Ema�-���R��ڋ��tϟpo�]t:�k���:�U�q�t��g��KXz��sY�&a u7l�6՚�<����[�?q}��5R��2�֢z��b�i۹�C�:n�\h�i��юo��23)l�x�$�8^۾�1��Yl��8D�"��omŏ�·�`V�p�_�+�_P���ЗyF�}j�K��v�"�Z���QRK�3����8�@=��6�g\��Cx3�]j���+v�#e�^W:��P����0߬�o�t��YO�!�{���g������O�"�TA@P�s�1�K-��d[-�2(
�X��Z1E,�
E��TQIiU���A`���kIX���ҭ��FcAq��HT�A�,���*J���"V*�,YYY+J�+ZȰ����X��T�&diPX6�dD�*(�T�EP�����B���Q���X#d�QB��2�@���E
�X*"�
�k!R�*�b0���+)
�1ҰP[m-�*�m�DPY"�
� �H,����UEĕEEU�J�Z�1EH�*���
�b�,YmQb�X3\q��Z�X�e`.!P
��Y�
��Y�H��I�0�`)QeI�\_W.DI�+� 3�rcCs~�g�.��68}�cȵ��Y	P(藧l���⩰�z�I�����a��=�3�?{�x{��ԛ��9�K��y��}~�Q�WcZ*��t9������V������G��{�'-�p�6.]�&�����7[�wG��Fm(Eq���Z֍ǕԮK��8�|˔��{ކ��g�ϋ!^ٓ7,p�dqd燃�ؔ�6�=YN��8w!��(��M�SO�_>Z����ٷi
��2_+.���nA�[R�_\�X�(����aK��������lmӉ�|+{E�����_>W��N�P�ԙ/%��@�x����{-4��;�^C�O!�{׾5�@EF���cu�{����fDm��vg�b��Ѽ��]k����R�AO}�?)p��al��]d��
��<�՘��D-}̴�9�q��m�e��ۥޙ�3�e�r��c]Eۈ=�j6����j���>�����߫ܫ�^�w~��z_҄ό�g��ˈ*r	MLWt��e���������z�ryd��l�̖F}�q���Cf��2F�/�c��x��T�=��r]�QW���Ҏ�}�j�$LO�5t��m��#f�������Ͻ(��r7�e����]���	�'_����J��_2����t9�ꌈ�r��ے���^���ok4��f-��SD>��ɥ�)�)\��p��L�0
t:�5���<s�}��̖i��PM>���rx�΂�͌kܪ@ƌHލ�B�C]�cg�}=�z�SH{�7��ed�]�L)���ru��2�����4�0-u@�B�Z�wg`��W�PI��oz6��W��eս��o���uB�δU_E��B�R�J�h�����XòF�OJљ�.���z�B|�9������'&���'�z����O��{*o�q�ˉ�i���.րkd����->���ӌ�d-�|��ƭ��ۛX���v�n�Q:���JX��_u;��[��^{+�� �;$��'Z���ݽ�z�q�6�s��y�y�y�z��z�����WDd���t�ؽ�V�3��-�Ir�!HL<`��^��i������D���`<�hx�uo�*��#~�MF����� A@��I�j��뗴�(��\�j`l�B�k���n\G�	H87nZ{|&z��������q�.�r���t�Yy�3�:����<��e�+[Be�QS���	˙\�7��zt6��j$w}�W�lU��=�+@2��Jx!��C[�T}-颓ˈk�|3�q��)I��f��jg61w^��bv-��t���ב@a��qٷ�N�{����ϛ���v�ev㩭��j��mQ������BP�|R�CW<����������wQ݆��'��juKb3�Z;�4�
i�:g���
}5K�r'a{iS��
3�K�r'.dS�L��4�0��|��n·\�V��0oU^g�Ŝ�u�z�gf���UI�����F����q��Y]<�ȵ�m_b�
��Q&�=~���Gxlh�~z[篪��F�1Ƽی�S"��|��6���}�/ie.B@��x�f*2�:W=]�(,�hoK�|�:���;�̽O�c�>��9=Ew�k*��ե�0�\IZ2�9:��N���h�ĺ�\�0U��~�����_Ś,��@z�S���`
Y�2�t%<͟{ʵ�y)<|�-O��u����]���ٜVW��T�Oy/?L�gv>.e�:����:�G(�T۵���`�oS����c�ݡ�o:RC&_L�uh�S�U�=�j��,���c���C������jD}}^2�פ�Ѫ�
��X�V	�{9��(%�!ol9k�7ٺ�<�7C�̨*�ꍧZ�hV�u=��i)Wg^�<�6+�b�Z}q�6�t�휪A�U4���& g�-�B��u�n��cT�ק��^�됋n(��^o��z�+/q�g}T:T�Z܆;d�B�uFԩW�u�R��9�����{(7�U��[w�2�b����՝w�/�C'��pQP(����*��٨)<�p�މ��\9۪��oo��r�v��R�D
�>~	1ZRV����N�!�(ǚ� ,�=	���_63���(�!O��t�`%��Jk;l�gyBȌ$�x�x�q���jZV�kX����r��!u	J�2
{W	�eI����Z�=..�{a������������"}�c����q3I�39��<�B������<�����3������<雌�s���B�ʘ�\Ff�1�Oӯk�B���=F�`�c�[>}�n��j���KY8s��E�9Ǭ���ZYG3�g4]ne]�e�Φ�"�3��]�I�޻�۝�?�=���\;XMe���󚉵�W�ru�I����q��N��	v�y}�y,#���^s���9�+�umjz�Tk�NU��MPK��p�L�3NT��%��khe�C�6j����ˋ��^��	�/d��Os�cyzڌ���r*���.�wۘ|�M�sk����E��Yꈤ�@3��u`�;Vٽs�5���p��	��|�8͌���V`Z-��IZ3O[���׍��,�Ѻ�wH�Y���������MNN�Ip�����4��M��m�]y�6�M5��J���[a;8q�V�U���i��ꄴ9\1�V�{�E4�ch�It�);X��ǣ�|��񘽐ۧ�b;��w�5��b*��Q��NK�ʜ�kcWa�2�bZ����C��0T�>[)>�A��6umJ�2	gF^#$��J�7�qB8�&&�,2�U�J�h{�Õ�F�Y꾷LK��ؽ�av�CPJM�%��)�]X��.���T�����V����(j[=�aSVs{�(Թ����<��
�vj�.!Dav��-T��� -��	� �p~�����[{����eO�3^'��y+�=�F��q�>�������LV
�O6����m����j�o��.ƻꇌ�9J����P��3�9N�C���o��׻����c���M��r�d�=�W�5�p�y�mACi��#A��f��=Ϣ�X��ri[/�b�3i���mmM���Ԟ��VC��/B�ʾß�f�x\�mS��:xl�{+���J��N%Ǆ����~R��Cd�lG�ӏ}�Vog34l���uwep��t��a�@.��͌k�O���!�ka���<�
Ӂ]/�4��3��Ln�W�ھ^�u���3���Pjg��������9=Gk�+h'E'񗶝n�,��eս��E��׎�k֦u���R�[�y�ynp���\A��_L@�Tf�`�|���p�^���QηU��WFA����.�+�q/�,�
VT�9���01sƀ��ŷ�i���R�]Z��5�uΆ:��~���R��y%�Ӧq��Tep��QބPh�+��vcp�ٸp{�.��P��q�p����c�y��)�R���bѼ���xx�ǯ�9y9R�h��J��";z���)<㕖$-|���t��.�m�4/�}�r��}�?8~��M�8wG��͡��hNp|�;(F��-crB/��u]p.����b�z�/o��9QH�U�Թ[|�:�u�J��Jn���wR���xˆ���ͣ1}���b�Օv�9�s�0Ou5AZV'E�컧aWʕM.on�އ��i��m�;MŠA�eʮ��� ���/8֔��*�[�_��{��/KS�4MK=��Y)r�=�������	h���Y��X�_n�3op���0iX���i���ӕQ�D)�J�)h���y������b�*�L�����͢z����qj06�)�2�]_	J4YO���n��;��z�o	����9]��>f����l>YJ&~�6`qԉ�d�mj�q�	���bӶ�5���\�hL�]��Ȯ?��� ٝ�M����w٨+Wq����X}"ݾ��+`:l8�B�}���K�w��.��c�j��]WR��	wu�OQ�>Q�`��T�+�j�lm��׬�}��h�݇����tV�#��>����Mha�6���%fecy�je��u���MƵq�k�9m��Z�6_��|o���_��8�=4�=j�rrz-8E�3c�g�&@��h+�ڤg����Y� ����]�z��^�;�/o�zVQfV�XԜ�����c���H[��]E�P2��=�j��e�;vjv���|n� �g��k���'���x]��*3u�w�D�E
�äHy�V��{-L�	����p��ؼ�f���Ѻ����S7�7=<��G���'���O�/� ca��/��]������{��b7+���g�9���\U�rq��]p��|�}h7�T�}f�ȓ9��Z�kl�����������w�JV�o��D=qW�.ܿ[Qk�վMv�:�fu!�� �Em$�1Pn^Δ�q���YiQ�m�����[��ִ^Nt�>Qi�B��r��4S��\[����Yj��w��퉧�r΋���t2�<�:�,;#2��S�.6[�%ِ.�7����n�{�o4Z�WHT���x� =��uz0���7lou���xN�<�㡡+��7(;�t:{���L`$�iIZ��f�)��2(�P��������2�Tѳ��3or�q�P�r��!w��X%-�������J	{z��P��o�RҶsZc,l6��9f~D.���Hl��R��	Vv^�7`3}�J�{�6���\ղ�;gW b�Uo�RW��T�Nbz�>�"�\�jA��%=�[���Iԓ�7��Ulмy�{V��Z�O>�;DO�H=���f��v��O&��㖙6��q��;\���/�g!�u8щ�feE��e<�';^�����e�RP���GM�W��b�3��/+�g2����Nڻ줧�Y5֭kc�y�$F��u'��ʗ��k#]���f�P̢��D�"&�:����jVT:�A�\F�{��~�iڔ�B]� �^b�tQ��cE�[��{"h��*.ή��H�6��Ꭱ�J���l� ���L��.^�HS /k/s�o��;]�Ӟ	m*uюr����gcBOT7���]����'���n��͛J�
��n�q#i�]]�4�\s��E������_|Y�<;q���7��)�cu�u�I��,-i�����+�UӀzޅ�e���x.ˍ�.X]�܃���MN�J��W���E��ʙF�-ގg:���,Ei̯R���3�6��G|�y�^]6#��J�uw�g[��BI�kvt׺�z�_���[�������ʾ�I�=�e��U[p�gU�k���s�)���4�z�5��{V�m�J�P����1������Y{w&�ƞwK�;���Ƅ���}��5��g<f��)T

0�Fn��T%�;���ꐃ���iMb�_s-%�opScݮ����x���u;ʻ����E}���琳�����p����M��5��F]Z�&�o�%�<���`�+\�u.ٽ���t1w :(���0��:|�ku9W%٨&[�u����ѓ��^=�4�^K����x��{h,&��=R����+�����W]�����]<���d���t�L$�Ւ�A�f4�L��D�f�Q��]�)�r	����w���EYٻ��˫r�ˆ��˨bn�s0�R��שׂN�{�EsB����P'Y���D{�֭���
�uq<�ҳ�,�}��|��v�S�[|Ƭ���4/JV��H!j��{(�i��]ms�� 3Vy���U�%;����K ��$wf*��(ua�ݮ���Uv��0�k$�V��QjDQ��,���}{ڎ�&�P�بm'ƭNq]c�8������XR����K�f�ّS������8���Lӵdb��T�7[�v�@S|9�9��J\�]��D���0���
'�9�&폟tЪ-$:�DR������AVxijg�X��)��7 k�S�U�-�S�rdX��<1Ǖ�ɧ�F��!��d[z�������U��3���٣u���3MO�ͱD2U8��Z�dv\�T�о��$f���ԣ���2v$t��8��&�ts۰�V�L���D�׼�*��m�X���r��Mh��Gb��C;`;�#�:���v��{�$��z�exY��Ӯzt��X�<Եs�eŝ�}֨}+L֧lB�C��X��G{��_$�I�i�o�:O^;��cG.�����M��/mY��@t��z�L�N�T��ګ5;2͐a���K�)k�b=H���m�w6o���@a��!��h�+j�h������;y�̻�XJ�ƪ�aCظ�lZ�l�l˳E�[3�8�Is;/0�K�f_N�$��Ч�;���Z�1J��^tr�vfm9�9Y-�L�i﫧�N�Ր��;v�S�}D����{`s�tq��8����d�ܾ��ڳ��S�9:ğwk�4�6���Hܳ��/i�kI,b�s�=̢���C-�9�z!	��q��ǀ�b~N\<�w�-i���i�v@,Ù9�!�=�ٶ#Nn�ڔ��z��^D���ܼǺ��ݳ:��o��� ��]���r*q*�u��
��{�q�\�_��g�����P޺�q+�X��)׵�NPE�kuw�e0���Қ�����ˊ��{R{f�7;W�f��կx)N�	��A�gbJ]��D���v�w�d}Wk���u3�9�;*��{��z����.	>EK���;A�X��@Q<�d�䛛W׼�x5�ud)�Hr�'i+�6�Z{����	{�㸗b4�J�8��������[qd7���<�*���:�WC�oXm����h V�s{�޺�y��ss��M�8��Yםq�`7u����Ȏ�/�ˈ�kmu�a1o�ep�H�,Mg]]#�!����-�4��?l��G�fuD�� �M+y�\����5��r��sc��vγ��Φ
�n��{��#]���W̱�a���&K�ȗ@�W��,����~&1Ea�<eC�(-k PQd�$D�3,	�E�+��b�R�*)Y%j0���,*
 ��m-���B�2�XT��4�R������I�%�$��1"��-�k��dPX(�c���c+�J�VVR�d�b� ��J��R�Ab��!Y*���X�V$Y
°��VHQ�R-�+*"���XAd����RQ��V�P�%�YXҐX
�� �*B�"�Y*@P��-d��}�TEiN�tw�� PK�󙝶M��)��Z�d;Ϭn�1w�o��-aq�n�D�4�07���Z����L�!+����lf�֔:���f<��Ϩ�]�xsc�*�1�ѷ	mh����gV��5D�����;����K1�ھCy�/_0�!nc)���K؃��4�k�f���ђ�w=,&�켞\6�S��+2����t:����}c2�Y3mz��B��w�1O �E�	���:e�����H�8�IO�W$Ͻ۶��^S>0��:��ƽ9MZ̔¼.&/�d'm�ӻ�3�o6�jН`���Zۆ���ٷ�s")�U��C)�М���D�z�x�F;¦�k��T&�ܦ�\�͸y��휔�p5j��ڞ��bo��Ԕ�2-��sz7<-�n����=^��W����;^����e�pݤ�sF���r�,�U.]�XtWT׻[ǰ�py+���O��ʐ;1��D�\��!��s��`>gBJԆ�%�4Rymc]�>ļ�󤦸�{�B�dc+U��ԢW�g�����Һu�Rh����3d�Y�8K���T|����X�F��iJkI���7q9�Nʱaߞ�@�u�j'�F���y�3��J۽ΐ���J������ݣ���5c�ִN�7n�}��x{��vg7
mm+7�s}QQ���*�TF�k0-�O�/�B܂`��gX��tx���O�I��^~�pϑ
~�Jb
Z*�y�v=ה�w���(�̩�˜3��C;�����@��h	�ͬu[��u�+9�x�Fw7�cw�=�	s4��ضB�EQ�l��g�%�ɵ�qշ�?�,���,���^��4�phlcC���-�=���pu__%����m��y8��U�����p�6ƥCdc�0�\�rO_,k;Z��F%���'�V���Tޞ��<��^3��XtU���=��/�6�~���މg����ȅ�]� e=R{"н��)d��)+ƸWVB]�\��6޾C]FW�r7�*��̨��G�s�ƞ,4�B\j�H=Tul[tJo�����~o�V�H	�u�qw@�e���LR��9c�U˺'0J*󠴣���f�	��2tx�#һ%�Du)\�4��"����%�J�� '�F���ovAk���^c���q}��DC:z��K6���u�g����rdqy�{�+؞:&�}E���}w��XKz��.�e�xP?ǽ�V[id���_�V�c�l��E�M��i��+�U�eJ��n	�ʪ}��5�P��g.w�*juBW�ҿ�cp�|�������5e#��6މ�[n�����UG��걭^�`�K����b�N'�0�F�U%ml�>F��ku����0:J�(��Ib���OeD� �hlgS�V�{s!v8z�<㔥*�P����`$�iI-)�V90# ����ji�V���_r�9��P�r��!O}�0X�ޅ4\v险-`�}tv9�v!�����:_r�ֱ��P�:�(�w(���{�M����s��'=+�pM��xeB\ղ�;gW�����m:����η�8�A���m�Z��쭎���h��>�P�a�\�f�\]USr�����u5mIS���j�� ��ϛ篼���V\8s����Y[+NgL��]�6z;��@ {�7;�{k���zZNr��H����k�\`I�u�amI�]$r睭�/`Z�ב�t�Y{�n&���'�|I�O��8�Z����].��H\ɼkfV0CV�Z󓻮��Bnv*R�V�軜���xX5okim\�8�a�ͱ�����q����[YO1zs��+0�=���X�Գng��nVo'9i�<�1�ڇs��^ �����Ie��Y�I��3x�s������3��Z���Xnq��uV�u��:.�)Մ��wb7�y��O�wy��w���*z�O7����eભ�W�k�*��N�j��x���3U�\�+o�*��b��nRl\��3�����6� fm�������4����9QH>
�U�ꚝP��t�cbd-�L�}�������#x�����z2�����@�:Ƽ�}[�z/PVYes��/ti������v�C�A�=^��P+6�1����$z���83O�E.�F]V���mN�M>O_�=j-��)h�����vb�z��}U�q��X㍯_V4%�4{i����^Ӷn����%�������Ҽ�;m���G�c+���X�;4�`��{yy�j閤6]������hC���WV��er�5:�������k2�����.��ѭ��9.e�����1�wM�y��.��;���T��P���l�ftr�w&(1��Y��%b���x
���=�N��%'@���Y��TB��nZL^������Fdv�y�Q�J��a���CSA��f��=��b�|�rD�z)�+K��q�u�˫�ȷ�4TCy�g�(��R���Z棩v��o'�b�x�9̝+)�)��Ӎ�f�|�ˍj��g����\��1�<���zԝ��s��Y��/���o}%ŭpkÛ�*���� B�0����;�G>�9+Z=�:}�Nv�f;��W�o:����[L��UG�{YY�e$��p���Pe�_�φ+2���k>�C�*��U
�c�V����y�h��軍w}^2�/D�E��i�fy�����Osd��-�Y���N��+yy>Z��軠)���s�'�r�Ƹ�F�wj1�թMl�RE�8�.֚�s��yTYw��hq�p��ચ�wR��<ͼ�3k��/���a��}��{x�r��q��w�jz
j���XȪQ\b�J��v"�h������	c`��&�fS4-	����6Wr@��(��eq����>���
��i��3�-�����W�`iTǭxfaYun�3�J���cd͓���B�_�%u-ƾn��z���A��X��tFI�Hz��GpQ�)o�y[u;�c3�Q���S���c[�5���%��of;l�A�[�G��ĳr���َގ�@���vOK���D*U4��|��c���3��:(�ΐi��4^JW�,P�h+���iI^*��5'��5�|�.4=&o�T�P+p�R�D

{��T���<�B��O����/,�sC�pM�F�����p�U��v���gU޵X���[��5W��ri[9���5�������P4U�Z�3by�J����;��S���n��ʈK��m�w��A�J&~�6��rehW�Vp\���)5�zSܥ���2����CI���|�;���..+�����g�1����anX۴�7��]�9�:�e��e�
��O����X�-�n7X�� /]�ݵ;�
u��ڬw�}�$�c��r���St-k�@��og�D=ޣb�j����%�������^Ƿ�c�c���7�uo�;�ҫ޺3����T���п�h�4�
Ŏ�y�:�8�퍊JD�B�������sd��i������zyT��,��Jh�$joOERy�ʷ�3��E�.��v�j�'���8�(�@Ɗ��~����OTOd[���g�L�
6�\�6s">/{ƽ���7�s�����#u�fQw?b��1�䄄]�}�e.��D���q��8�)7
Z�A��[y>M�k���j����(Z��Z�P��N�V֐ᮌ.:������`���Wf���B[Fdˁ���d�_ ��8�=�.�U�Թ:�,t'�\;So��Y0�:y*vkǵ5ܺ��e\��.�8��b7�ʝ��j���*V9�m�-��BhQ��3r��s_١ki�A��C��ϔo�I+�T����2�'��צf��w�'c������JU���邠�c2���{��j�gy�=�u�yY�Ξ�y�޸Gkb��6ܣ(�=�s� a4y<�������:R�7o�n-ݏ�J��[s6B���n�W����Y�+±�ь	��j햞�y����{�v��涄m��]��{��j]p�*Z��� m��������kp�5s��F�굼ve�R2�]+��o{o{��7���J�pq`�E7��[Է�n�ɛ��-F6�W��vnT�p�c5�{�/9j����O:�h0y��u.{�t��T%�[/��gY��j�+y�DNT�''<g�d���ul-s�6�j�������=��y<�X۩a���h�21����'$j�����9�j�Vִ;(="\��^��B��r �*��x���8�lc]u8щ�gл�_=�z�����h[�x?�a��~ΗS�ؼ�ڋ��I�Zp�<v5ѽVn�s��GqɀT3�����$J�~�ݍC1�˭h����>�uB��R�,� k�C����e�j357�{�н�"��g��^v���O�բ�%�p���ǌ擣�=ih�^��������%k�T�7�,��s�om�_F$��� �%b7B��<�vK�X����;�jAz�(�E'M�h��̻��{)[�h��KD7�ܩ>��}yvsN5�'�v�+����kxzp�Hg �?a��ʓ0��PB�Ǉo�2����+�\��o1�r��3�>��6-%�����xe���%��d�2����T
���Ņy��=��}އ==/>���H��`U�.QD�!sL���M��)^O1ݠ�Z��z���
͡��**WP�a<�j��e+�n{���t�k���m�jr�6�@�ܣj��ůj��Cam|K�����5�b�w-��e�X�c��6��u�k�����v���/5{��G�w`���%\����Ƽ��g\�>��J�*�&�4����2�]B�������j����!!�3j�6uKɡeS�<�b��k"~T���@�QA���GR���t�J�̌��#4B��1i�4���q�\b�O!�����0	�F'��i�j�2P����&���Bn5ں����V�J�,�Il s;B޴l���S��"u�״��\ru���+�;�g7i����[�k��w$z�ߤÓvGS��]9�L�t�l��){��aDN�
m�e��8���C4��k~X�ui��u�Ä\/������f�釅�ꌬ�O<
�^�F��TX��i�-˃�k�C��s�n5��*�a/�D(:��y�l�o]�
�����UNA=�E۠eݡ;����.S��^��5�*
ٓ�v���S��ӓmBW85����U[��:�.����D�E�{��׀�ڤSӽ�6�{8�9��5�bi�gY7���:b��z�'n����ɭTr�����7=Q[��\�q�m�{��[,���壎U�&x]�lx#�wˮz\�Bw\*�ب�ܦ��O�:,��o]���+F��gp��wQ�Qp�*�5����\lW��A�z���
�B�:����nQ�裮)�`�ʶ���PZ�T�˛��c��{cL��2�l*�i�bmq�X��*���#��Ғ��Pu����wy}�.��ۛ ׼���O�婾P�)J��>
4%�G5|�N�}f��`37"{W�]d�Q{)��q��}��3��D)��JC �����/*���!���0Y�j�[�֪{f�zh@cA}��Yy�jT���Q*�t>Kk�����&.k�S���1�4��v����-v4��[A<��'Uw5�+��d�V91.\np:�y�C]9�L�r����r�b�%�{o�%�����}͛�=����_E2L|-��:�^瓒��0�ygIT����r:/vIQ���#U��t�0����i\�gtR���8��>�n��U�)_'�)Y����ٕ�eZ��-�����6 ��r�+|k��x7���|0�ɴמ�מ#(��U�1��Be���=���^���,[�!r*�H���U�9+��H�s�6�Nc���ȮJ3uF�LS5DGv����(i��9PB�j���r=EW��}��+G�=���ΠƠ3��ƛ�Fꮋ��Ty��5N[��wam��{w��WK�Xw�\�9�uZ���K~�����&ī��+)\<��+6C[�8Pۤz@!�o�:w��}��:���V$5�ㄡ����.�Yx��O��ɂ�����',��mԤ�ͤ��6Ԛ�:�{�vs�ulC�:�ˁ��3>�YXyr������n��b�=f`r�n�N�['U��דC2�[�8д�,� ����
��IdR��I\Dt�`f�:e�x5�VQ/������/_n�����~s�{�8Q�y(��N޹2��D[݄��� ��
��L��	n�oa{]F,�P�
�N�H���������;���l�,ZR�<��Ď�}�h�yMva�l-��Z�
9Y#˵J��"t�ǩ�ː��g���S��Aufq2�wp��)��R���f��-�Aʙ�+p�o�����9�h��37W��q�w��P�"�u���Zi�3���J��֦VN��+)M�AR;�9��ϖ�IZ���Co:wH2��*�3�p���s��Wv��x�ވ4�٫ �d��j��gZ�9�٘ATu�R�L�ll���]n��(HT�ۖL��.c�l�8s�9��P��op���&��z�w��J5�A9�܋�w�uǻVrl��WYĮJfR��:�T%�WU�lѤ]�*���-�wE�]���:��	ʣ�I�N>���ey�uQ��[]yIp��m*M�՚t���',�r��q�ތ�z�,�G^*���r>0p���u�NR[�s&ܣ�oH�r��ۺL�(>,A�eG���;e%zOs�4���ywb`䬘S�Q`Q��
�d�,�]\�Ӝ*eN����i�R�������J{Kk�!�xѹr�&l"I�z�N1��3��^�z����Y����o{[�,7cz�ɽ�g@�聲r.�ːe�8��De�7�d�����J�^�PJv��S��B(tF��}�?^��]9��}dm^>sF(;�����&�LC-@�Kj��C]Z +��Z���yv�S�b��u.��Ӫ1���ӗ��I�I�� �iԫ��I�ͫ�\�N�i~aDJ�Qd�VTZ�T��VB�iYF����F�+�TR"l��E�H�,��ihU`(��R)Uc�a+�m	X�P�P%�[H���RT"�)hUk*,
�X�UX-TQdZ�T"$kJ�j���B�V`�V���+"�F1���aP�F��#kl�	�W
*
V"el
��"�1EEV)
��VT�b�TZ&!��
�ʒ�1�!&*��bCVT����+YQ`-J��*TbEY-��
´e`��	X�U�b�(Q*�U*�"��T R�Kk��@��q��"�6���9gH��ok��iE�h��FOY���᪸zf�{�c�TK����uX���i���Jo%�g+�#/�=�	4��mD3�)��P�����;����{���DD����Y�]I��&�{�*�[|��a�,��L��	���&�)��'�?��C.`�����W�o-��ˤ��CI�I�֊9*��SN��K��}prHV5��J��7�)fvW���xo::�="�&]�k{�v�&$��ӹ�Db���fp//�k��s*�l�!M�Ҍ��l&sh��y/��g����jqѥ�_E�.u1Q�}��+{t>.����t���-Բ�W��o��#7ד�F�#�]�-eӯ�qq]�Xփ��Sr�zN���|Ӏ�a}.ֶ�{�m��+�{�T��^�����s���}��HP�aq��lW�&�Ĵ���L�[���X�T�]ˎV]}L.�.�Y%��p�^��m�&^��ޤ��&W��F�e�±IpW�R�7#�0}wH��isn� ���kpNڎ�Z7� :sI��ڷ�(*ѫvÚ\����Im��DP��9C�ۛ7o�G��+�̗0�O��U:��*ӱX�7��uXԵ���i�$���/�!�.��W����K��+|#�T����^�`滟u^b;��{��e��9V���=��u�Ci��oz�P���0T����p��7VFΆ�gR�����鯋o9�X��X�zm��a�[��Q﷓;�*՜7�Y&��-�79���T�Y}܎>�lgT<g+�r��3�p����}v�u�.�ꐃ���i�>z��m�i_�浐�����ލ�Vk[���(���ʆ��M}Թ��C�\�����図�ux�UJ�	��Vc�G� �F'��6;�m��M.������g"�6�%{ct�)<_����61��䎎Cd��[�s�Tg��Ъ�#׉��s��k�MI�8F�mƴ:�q��6avTZ����u����['y�w>��{Y��N�ָr���w�������l?1o�ʕ�(`�Ukdu�T���,��pWz���dVxc��'��΋�)� v��ۉ����7YS���煮�w��o�b�5�Eox,틱�o^���Im%&3#i.C�پ�h��Z������H���iHWN!���ź�&o�g_��X�]��A\̱�n�^���N�r�ڙz��k5����ݠ���Q�j��͵�F^��7�c�7XG1{��r�h��R�qݳ�?(�nf��I^�����eDs�|�rt��|�+<"�0'v<3H���{U�/���?gD�ryE������V���nn>��N�r��2�$�ٺ���*�oe����og��TRf9�.frz�����!��ͱjOU�\�cv�C�A�=/�o��:��������R�ydoְC
����Ԩ:�N��y��5�C·���6�E\:V���[UBU��r���|���3Q�%�q��Ơ��mc]�>�h�����0���w�k0��{m^����`�`���O5��-}���٢��]f>��_hB�z�v,`n�E��Y�B����`�٨�\�Ո�>�{3 �)u楍O�X��$�n��}��+��Vlw�c��V�K���o/	B�5�ˠ�՟������*�Np*"�<���;^��la��/7��Vi��[-t'�u�E��7b��2�s����Kt�Ft��gAvL{���B:���0�ܧ˹D��H�����4ͱ_5�*��⋠R�k��D��7���O��ދM�go5K���c�{�ζ���{�:x�ѓ�r�-f���K{0k�h*׳{�kS�&�ծ`����D;���I"�p��K:-�ג�r��}�cۉ�ή7^��\���ᕌ�ev�����8���g���z���ߪ���d�m��SZ�j{=^��3"��u�D?.�+�y�nm#������ѮD]�)��OdZ��s|n�sWv֊��K���y��=|���C/�HoE۪=���]�ㇲD�����N�vv�Ԏ�ſa�!7̡=�������4m�F�WC��;Y0�B������6����뮩�N�-TalW4��SoT��N�V#~�暨�M�J��8wI��mL@-TmJ�����\l<_Ci�_=�sZ�{'�Ob�DeHl9�1po�F7��ji��Ehի���F�gS6֬e*epA|^��0��x`���80��	�ޔ��W�'��3w*�ɹϖ��R��ǻںp��s��j���#��i�ᐋ�J���/3+��0�r�)�x����s�s��,ڕF�@����z^�]aWʕMB����c]:�PiIA8�f���l
�ُO�ơ�#gǽ��{�}P�x, ���=+=]����� ��=�|3���)W����BZ+�<�a�Ƞj�'���E
���̅�L�������۟7�3���B�3)1�z�+�]��x?�}�-ᔓJ�������l�!p2V��i��|]�����O�J��A�f���j�{^�ʆ��m�v�0�C̞:9�ӥ^�=�[��WC� �P�j�{Е۔�r�L��J�@�m�	��Y����J��d�����/'[�ν��D�b�=-��}��}*���sP������m���b2�M������^���eݡ���h��ѽ�J�W������yums���2���G�ٺ�2E����s1j�߭*��<љ�̜ў�U`;�?�qzFk�u*U�ibV��CdT9�CR��2��֠��9X��mk���z����srݠb��.���ц.���Vf���{���̸gv0V�,񏪰<yr���zA�t��Aa�>ygu�|3�����^���یm�O>�2�o��t6�y1�F��G_���б��x��ޅd��ћ��;ѷ0-|�=���bo�V�r4/Bղ<�ejkۛ����p~�KK~�ƭ�˛�<!e���S�n�z��*��ܶ���O=�)嗝8�Z;��8��PR���]p���]��!��Ӷ�Sɩڜ|6����/^��F�=T��)�<�OKخ��,º�E׋z��S9���.!�k����oz��@t�P~��f��=���_�x�wY>��X�h*�Sٯ�O9�X��[P�T)J���f���*����ј:��b����kz�T�k�/����ؽ��[����+##u�>�d���v|4�EF��d�P��mKI�֓;� ���NA��ݎx���g�d.���C@��qԹ��C�_r�}B���.���mA�X��ϔ�ej��K`�%fL��aջ�n̮T�#˼\Ӡw�+r�hO���W%i��mt*�e䎮�s��&Ÿ0�yr=�!�ݱ�[��0*!ouE���#Z��6onj;J�e�v�G�b�f.�K��A�U;5��k4:�k�	y��T�w�p��xb�w�dG��ҝ��n���i��\ӕ�*�$'M�O�Q��L8n1�+��1�l� ��W�[���ɡx�vje��iF-m��N�4ί���7k*c]��v@���� ���W8�1�S�<��n�۝\�>�{Q�����������`�%�y#W��O:�s�^�$a7_�S6���|:�S���)���O��#E^=�]��U\��<u���A��Bv}iu��}�zѥ:��{������`J�U�;����c���𤖽�&溾��V���m�fV!�Z��!�)u�2�.'B�[|k:'Ų�[[��8����nN^ �������bM*���zz��1�Qm7���/�
۞�@g}�`f�]�_>1W�4�-��X+*NK�L�ĩX�����y�=@K��fע�Tȍ���MJ9F�γy;%�f����FNClWrĶ�Xk�&��e]���{[s���5��6M�ל{m�D��;�y;c9Rw��pY��`q��;U�7�o�t1I���uc%�pjT,�wUyBf,"�e5۰2Jf�:�isF;���}������ϩPt�������kn����z�
lr�!c4{�[��3�{j_ˤ�?�kJJ��Z��o�Ao��kPP����wW�-j��*!Ov×�c������V�k1ꏖ��&�q⺭��u�i��y�e�Ub���EE�6��(�=	F��gv�=�ɠ+{K�./����g�?�8g&�5�6m�����R3�#�dB��Hl��dd���{�9,*�ٸ��kG+�\�6�;eƻYJ&yk���V�N6l?oT�o���U���f�t�����O}%Ů`��+�''J���P�x�3�{1��k�e���ǞF�>��ߞ��W�{Y]���ϥ��Y�,N�E��A���3Ђ���g�%�g�9:[5M����^�Ώ=:r���a�es�k�K5�ꌹ��f�̨<�f*�a�5y���\j�]��������%��}ʛ� ���S�c0P����L�e�]r�C��Tݣ���˦��,;t�9�i/�T_�V�ԏY���o>!�� >����n3�!���\��e}��m�R�CعN� .^*��݋ZX^�W�	�8����LIZY5&��6s&׾���ٞ|w��{m<���r�T>F@�V�]*<�h�랢;x\M�L���ciou���ʤ@�	���]�W-�|%X)�*ښ�q���_P��P���m�z���PR�A�V뙤�cz��~�s��D��>�Pbt�ka�j�O����OM�[��V���X�{e�Sd�?ʣjz]�u�P�T�o��\��Fd�v�o8̮�Α��?^Ge��>���x�~$�x�b$�_I[2�v1��2yѿu\&�Ѽ�$+�&f�O���~ӑ�my���Dj7�R6�uL;˚D�5X�-�(rr�]�L�������F�7�Wz�i��;���:
���u�zi��25��#oh���������c�S������7��*6�[f<s��/���i7����Sŷכ�x��v���P*���^��D�*|�	NV�ॏ{��j�&/��㞙��1�d��&�ҍ����5��Az�$�I�D��25ml�9�jk�frő��7J}=��ǸP�K�gv��hS�c����gK��bF�3�[�����R�5�-��Gc�6P��=N5�Lf�:4i��d�+u�nb^�	.�:ҺÓU,p��zZ��X���FN��P�M�H��	��ߥ�i�k��w��fG*c���G�����9�ݴx1��̷����}Fg����#�&;�R)d������xK��7��[��!�oc���ۨ��d�̥aÜ[�=�Uɸ��Ͻ^ ���&�F���Y>��pwv��o��_����o�g)S;�gl�j:ϛ�q���o���iQ����}�ʃ���o�hܬ^6�~�_�����+H�Ϳ+�������rJ�x�ڧ�7��<�ϴ�>��W:�;��Y����߅gux��lvyhy�2s�3�gC���,��*6e�Q��#����/�V3����9c\�^Ϣ�0૥�p�-x%��_�D~ݺ��|��+gOB���K�<�i� �o����~��|�3mϫ/{Cw9�����Z���W��[�(����|��g>3��TϨ�s��>�܏}��K��Y��yZ�:%2=�|��{�ǔ����s���x���<j$��ʨw�4��}�샢H�*�����B�v}Ϣ���ǽ>£�'��{��q���j����UD)`�$0�(k����Y^�5��k��i����b��T���UwQ erD},�5c�h�3�������}ʖK��Ү��[��Lj��;r�G��o�;�Sn���
A/1ԑ!��%O����n�C��aj�)~�/��ZӬ��nlge�;�b�TK������X�+!c�2$s�߂o��x�a�+քQK�0Pb-*N7n���9�듯�V!��u��>�c�_R�8+�up��ސ��4���_rΓ3[��k�B�]ʆ�BF�/57a�f�yr��-ٞ��->��,�'�S�ow��\��d����4��%�U��"��;V�Q��w0�Vp)
���,�R�����]�Q���2��"�D�#��X��,t�!�ۖ{�)��ɧ)�z�3a�Ncx�k=��k�kx&7A�c+������9�Sb'��i���3����e�˻�.��3O=�Bp-�6]1�}�z�)_�15gb5�9���l٢�ϸ)D�f���-w���"�|��T���X�ޥ�]�s����Bn��0n��k�3n����_N�Z�Ӕ�hTz�����Έ���ZU��mKBŶT]4(�̤���Ϋ/��פ\�鉲 �%��"wDkht�j�Yi4������O�#�P^<��*����u*5���Y��1V%1Bkу�L�	S8)�Wzn��qɷSB�Ii[ü)�[b�Ig_;��o9�L�j�˟Q]e�L�/��|�i��ؒ�t��ug^���m�ץ���gs�[[�..��;���p��ff���b�f���Ż�KU�t����X��u��l٦|�X���C:�Pǟ;v�c#����;ܔp��g2��ہ�f�\2�bK�J�7[����Z��wMV9��Q<��]��(�g���7+��M�Ѱ`�gR�0%�K����^�. CCb^�8�S�R��|\s؞4ݎc��:�t�>H���,�I��t�Hz�L�L˧g6��8���r7]Fҫ4t �[�[�aRͦ�� �P�v��7.��`����A��캣���M-����¯k<�Ȩzp(�=�q^����]86��(C�Qj�'\|�.҆��� �P
�у�X�p�����ز��&*�g{���;{��W�ݸ�#�+��ҐC�z�w�퓱�Ֆ�:��	ѻ����3ziN���TY��q{FZ*�������n���n)n���ɞ��-�2��ҷi9v�4��.���R�wu��%�]�Wegn�Iv��2\]��N,�7�P/�.a�b�k^�YJ��zٸ��(�ۉH�<&�jX-��Yr��d���{)i�s�x}u��f�m��t���{��)�|���#o3��O��k�Bw=�d��ʆ�V��h�7�f�ɬ�&�(m��x-�.�;^3��\`�rs��Y�y*>�x�|��j.��*[�v����9ÏmZ���H�$�x@aR�,��aX,5*)�"�+m���
(�$Z�d+%aX�B�R(���T*Dk
�Y*[V
������H�1L��XJ���� ��"�V)���"(UAH-��%T�%bŖ�+Y*)QhʣUPS��Ղ%[J�h�Z�eQ�m���k(����kB�H%�(QE%@����EYX4�V(
��X�P�"ԣ+`�6�DX�,���1�d�,���� �V�Ķ�* �FV
��ł"5�����YD+R
+mB,��B��őB�@D}��6g�w5���Om���wPvLU��*өu��՝��#��hf��6{a�YW�r-��A��
�sf�w�T�PO�u\�P��IK���t�����>7��\U�w�8�#���t�{ڪFt9�]�6
;���
�vFc�3�2�
9mC��|��`�/Ņ��G����W�#���>�8yD{}q;���˟J���j��H�q��d�_z	TQ���H��u�wC�
��89�zw���R������M�����ՙ~�'։mTN�G��P̖U�����1�J�*7�+���~�={�����D��>̖g�{��>9F���)U�^xΆ\�`��MB�OT!x�ʊ����3���Y/;/;�:���`�e�@-�.�g�}5'�6��� z� �d:�'��O�3/��zv�Ïg�g��p9�W��Ͼ���Y��q����C󻓏����P���خ>ɓP�����^������sg�d#az=t��Ȯ�"����{p��V�_C�Ez��]A��=YF���uˇ�յuƳЕ�Fx��,�T�����F|��%gu1�������^/�١!�crn�<��CW>�W��q�+�����t���X�����z���3���������hX�V��X+���ɥ�f��f���쏴�M7�g��g�S�����1#��^F�Xѵ�l*C�P, �jV:d�
��7��TI1MV�ك(��λ,qrDv%���tx��B����=��V��=��w�	aZB1r���v��MF�ˊU��+�7qy�*u�{�c4����_�g,���!ٯ���ʭ=.���1Pw�6=���=�n{� �.~����.+���e���k�}�9'n.Y>F�K�Fz���Uct��q^9'�8P���Q�d��>���}^&���}��_��ȯ+�Y9\*NI�q�ޘ�{����5y���[b`��y�W�b��Rη4�����'�����+����kX��(�9�tqBU��c���@�,tWSy����X�'^=�Ҵ�%��H������{5zy	������g4Ê'�!Aʌ�$�28�����}�Z/����/�����ej�'sݪxk�=�Qү���q���;�rY�D��ĉ�i(l�|^`f����Ec��bBѝ���Fe�T�Ǻ����ӵ�=�G�Hq7������Nd�@��zH����;яQ鬟N�9���I[������o�r1y��f�?}]�`}7_AC�Y@9L�\���'�/x�ɹ���6�4��-���ǈ����{���3Q��j�'�>D������c��s2=;/�@��ݦ�o	������弩��sy �Ccuy�Jt��W��l�7�kt�c��>h]ܳ}�f��|]�<��\{������1,������w�N����2�R4�l���D��ѣiij�=�e�]}���$�t&���w��%Lp�ޓpƧP����3C�8*%Oi�yj���O�?mG���z̗���G�&}��Z�_>�#שּׁ2O��L>����Z��\�x�Guxu�Wzϓ��C-F�ߗ��m��p�8�&4_�L���#Ղ�������2a��a�ׯt�'H��<9yI���њ9�u�}�#��Az_zh+rhW��R2�6Y;���ߎ�C���q���^�[W롻V�B��/,���
��uU�s/��.��wd��iKN�D��2��C��b״o�=֮�ʙ^%�ٟ@��^�#�Q/�ϙ��w�����:l5#��Lw�7<�p��k�Ŝ��a/��c����y�tσ����+��}��~�x��+��^�e���%_k��KF{hǡ<��$�d<X����t�~�7��G�������3�S�z�u��Zօg݆��q�s�R�F��=�`	>T�Tʯ�B�Ziڊ���;�O�~#��[�֮9���ﻢ|�纈�{�Ǵ��T8�QCĔ��8)����l�t��������n /�X��hK���3�\��\q�3{;`�ۤM�R�Еީ.��w Ջ��J�)��.���-��K����`�V���j�eS���omv��B@�b����vx˃�[����зլ�#�L�S��p�g_�6g7�'��_���{^eyI�}�U#m�8k�Qs\b#�\;���:�Ĥ��9o(���+���Ƣ��\M��i����;����������2/QH9n�-�=^G��45TxnO��H��*�7�"���Σp�
���m����_�w�=��{޾�V�!�Y��q�J_##�s%�nL'$d��4.��Ƕ�=q�VF����Q�yY�}C,3�6���{�qB�k&��`OާS&�OP���*�dK������yʘ�~��f!=U�>����>�YW%zG�Z����z|{!��;�C����J�R�����������v�>o4�����������������_�=7&�F���e���gv�/�LN��w�Ul��z�q|{��{YLy��q�~�=.s��T	��Z��`E�1��"�>�����+���/����#T��UP�k�\��zW���=�oOJ~���m_\��(即4wIӷ<2�9���j�Ό�U�#fX��#�>��~>�V3�{Td�����+�ZL�K�o�����&,��s81�vV9�V,O���і\x�-U�w�������+��2���ud�<�ջ�:����+	%�����b�S:����������/��YF�4�Vޫ�{�����ܜ��R�PP{���m��r����,��w�A^�yS��N�,^<P������y��������Q�sn)�En�Y�͎�`:�>�^�YN��9�TVvT����0���b��Fy��N;��GK�=ܣ�vN�W�B��"�=�w=���ȯZ'+�D.ʔn,�O���j��#+��U.��&�	���u?:9�Yj7^��8^�a����{��q��yׇd�pV��K���'�|A�yYB��7�e,d��;�����t|o����qzG���%��uH��dWo%ev纴�5]ϫx)�O�`��@L��7e��>��s�~�*�=^��3���G�'JR3�s�QίMW`^B��]z'=���ȯL�iA*��"~��I�����s�[�hps�L
��S�[d=��Fh|�O�^'p�}���q��D�K+EL7bx����To�r��l^�݊�zǷ����g2��X�s�����"}�3��6>9>tК�K'hA��n�/k�31	c:������o}�����f��x?)�=�n�����C���AE�.|3=|��ӱ��hd]��L���NyR)�b�]޺�Ϳ{ ����]۳ܯ�X��qv�x�q�L��1��a�WT� '�7��5���Km�]�`ʐ&`<!%gS��n-�|��jx̞Z���:T�I�檅�[���OI�(�r�xo=wcಎ8�����{�������!
����uǳ��w&���rn#���yT7��d���X��Pr����,���?NG*��\�������n~��
z+�^F�.? ð��xJY��Y�5ߩYXgǏ�u������g<pj�H��,y��k#�W�"��xW�p���{}}�[��R��{*���;����Nb�3�'t�Me^��U�wU0ק��4.CȽ�{�eF��ڧ��;��W�4��z�-� ݊�~�,�=���*�:�ͩ^o�������H_g���2��zL�|=�SU��OΜ��Y>G�K��^e׼��2&���U�8��x7Ѿ�Wtn)Ϡ6r:}w7��Tg����/��g��~��ZnN
�*�g]^�����܍�Y%|����5��Ԅ5:�o[�;��+�'���t�>u��>��4�A�޶.5�ㇾVk��8}ă�� >,:�o<)ԟW��>TƏyS�g^x�)'�SJ�=��6�Uow8���uǻ�8�Q�*2��/L�������ZO�ٲ��lm�QTY���NW�������g#�j��*�mr�C.�ٝBkM;�����-X��5`�3(�.'�mM�-<�&{��,5�)V�1������x�16��CʱފhT�t�5�*�6na���5���',��xBWX�D\X�`2����Ã{������*:U����鸏S�w�,�Ȉ	Q��q7�+��q*�	RYG/��Ef�F�z�yם��zv�ǽ�᤬�����^���̗5� 6Gw��+F}+�6�jw�;��G�s�_G�5��>B�n��r�H�NW�����3_)�3�~�?L�D��>dfxZ��^�w��>>�&'�xU���Q�_��3Q������㞙��9�#w]S� �5w�o�VV��S2=e�H&��PYύFz�W�j��OJ���|�ܔ��>k�d����óF��}����p��ljl0��<;��O��F�m���^�����0�o}�N�1�LV�p�5sӒW����}����X(V��Y>���j�\~��[�9/�(�~����Ћ�U<z�m���`�Fu��{�>�_�x���X<o�4+��q����E��"/��3u�`D��vp�{T�Ȓ��>�K��~f}�eC�B��z�6�+Gxܛϔ�t��F�,�={��Ч�'��z�V]�ȩ��G>��p+��g�W�&Y�;�ݴ���}��`~βj�0��^�P�J���[J�d =�a:�h�=�zw:v�n�r-S�'�tЗ��O�y��hHs�e�ɨ�s�M�݀���ŉn|��{��
G��A��FgV��Ҭ�8Ifz�Ƿ����5��lt�ڒ������gx%1m��ԭ�tz7���̱�&xz��Y��y��'�`��r�c����j��0���g���W5t��9�=�S�������,uL���:�k�Xx7��A�d�o���̚�͆�Ӏw�w�ޯx����>*a��嵦C�k*�s𕱾�"�TX��3��#��K���ף#}��u����qȜ�Q$���=Pf�>��ڞ����pڝ���3�{u YU�ڄ�-������폶�>+�U#n!�0��g��!���z�;Gt{�B�7�#�u��3�/5�r7��_����r#�;�����W�{}r:���2���6����t[�콦����24�Sޭ��g�v�F�*��o�ٌ�N����L��ز8��݀.��I��j�F{'8�d�8fc��m?I`����r8��!�Y4���=(0�E��]�p�3�,��L���Tl	�ө�'��3�{��;Y=��7�O�?y��FX˺���9ٹ�<����s�W�>~��U0k�,��!��B^�ac3�I�h�-9,�k�e�e�x�e��,鶊/v0S�����D�A�ߊԁN��ƗGv����xuXj�%B�����P��B͠�|&���O�<
Q�S3K�Ίj�\8��m��s��&����63�(�W��Z,"�P2{n�it�Uz�ߒ��Q���������@9����q��B��H5,���n���xV}w9�O�X��s�\�Z;�S�7�{p���q�@r���tv~���	���M?w����X���S���.|=p6tz�ظU>�x�~7�|���k�.>��Ǟ��:��
koUVb�CV{��}��^��w��`Y���=Cӡ����b�W�o�1y�x(��~Z�N�:��󃵑��ŭbzul�o�����p�4�s��#�=�_R�~�u�a�o�)�阸�m{#uW�N
�z=����}O��)�Fi��D�b����'�@�,5�����;W��b㘠"=}���Jn�{�g{���4��E�z|��{���>�<9D�p��eH���:j$�����X�2dy*��}ޱ^���s]G���F�w�{N}���#�q�7������%k�g:k��"a�y��G��P$� z b�W�OŌ�t|o�_�&�iߴ���=�|z���f�F�L�lX��o�r�۟$k�����π���֙H����r!ߩ
��zЋo}k���Pe��fu~_��G�ؓ���8}x�����^�[*�f��:�cL��������Xv���7�`܄�Y�W�<�j��%$����y!N�l��'J�N�G�[b��l�E.��ն�x ���C�w��Rɴ�n�A�*���"WvF�Wn��㦽�+�ۏUx�;��|���Q%��8�#}�S��z��}�wުg"���S�̒�c�t�������q<n=^���d��Cz'���W���u�G�~��K�3��	j�	X�E�*"�M���_��t2|,*�{��d/�76��o��F]��n�����W��+�x�w��O��[S�_�k��D:�'�TA��N�L���A���3;�1+�����pTJU��'�;g#T�<��O��N3����@�臷a�[�B�������S7���/�R?�*������ذ+_/��g�)��:��-#!���E��u{�ܩ�H��r�Eq��:�5���8n4�U��8����[�OwK}�q�F��������_�L�����B�<��z�{X!z�hޖN홅���(ʯ�ة��N��_$�KC�s5/Kܩ���=}��2#�^�}�W2�顚{�xV{*B��a�؃�S{��h���P�P��>V}3��#MxX���2)����z��5Z;>{\+:rN�d��'�p8my�&$����'F��؁��^3{�1AR��6���N�Y��vD�yiII��4>�1��J��,���]N���k���Ӽ;Yu;S*46�ϝ�eʼ�uk�w"Q�K^�_cZ�����Ӯ�+c�Zy��`Dc[E���A�E%���X�V�{
V3x�l^c;��o<y��k��WV�'�3�ɏ@�g3v�<�|�P����ֻzw9�Jm�ux/��0np�Qb�	"�T��pM��%���;����]�q�+���m����^j�ΓV;8 ��B�!6,�-B^P��=fcOa|���v��V�n���ku�̊��L�^�4���_���=n��e;֕�Tk�O-�ۤ^YSB(+M��^[Ƨ_)���YLu;v*.�K�����T�@�fq��gn�A'i���V��h��84Ö�6*�]|{�aL��������lW}�>�:����#d��>DӪJ�e����������o�!�-uY�ڿ��C8y\��������ɝBY�`k�l���e��T�v� N'��#2�T�:����4��N�0a�j��)���8Jd�nn5[x/������F��ǜ�71�ƀ 3Q�p틵juJ8�s�݁�k�#Zs���bf�;Z�֊�!Ķ\���g�Y]�)��)���+mZM��z��.����fr�yPX^�x���۪�_6�f�p��H�ǎ�d�bT	yx���p��*=�n�w���qz<���yz�Ry��q �[��s+��^x�U��ޙ��R��R��5��=�}�{b���v���H�oM���A���66�b��n���(/����歝\��"
�y�<9��9�hU���V*$���qgOX"dE�������ܖ\��,s�+[�[Y4q�2 ���eN�׊���J�Bd����[�p��Ha��h��ѫ��W�y<������z`Y�]ovuCn�M�2��
��	K_4z�\4�]�o�g]^��H;�H36�J{K�	veN���Pj<o���uq����
�/�	��V�:r�l�0�K����^�^�����橊��/P���㩕���N�9|�d�<f���x;7�]�R<\�Č{g�����-H+2�_g9�V���;;���M�F���{NY7��0I�oep��ό=�$�X����[ٙi[�pj�Gr'!*�p�V��O�;�y,'&rAs+ϳ:��K����}}	v-�Y|qH\
�i������Kje>��^p��^w]��>>�/����;��n.�a�;���9GsSR65�=Nb>��+]-�o�;�^Vv�ia�*��}�WJ��3�����Y7���;��;ξP�/�.�ʒ�3C�
k����;�a;���v��99��/��f���y#8�A\�_l�x{��\ޙ����:b�-(�E�
ʂ���
E��i%Ve���X� ���X(E�E�@P���[i-��E���l��VJ�"��
�"�E�R,��-�X�TDT�	R�����(�d1�*��B�T�"�Uh������jU�+�VT�� ��(EU"�U�� 6�bVE�*-aUQAb+Y*�����+R�E�QEF��*�c2�U��b9�,B��U*���Qb0Qd���6�%�(Ƶ`�b*��֩R�i���(A����H,��UAE,[K*T����(���**�aP�DX�E���EAAn��+
 īlm�Q`�"ĨT�E������T��F�[@�m��U�j�X)�~�~u���۟�;����u^��;�|�k	�K�ڲet�����lA
�ܝ]�IWN�k�Ep5sn�X���Z�f�u�%}�~u�uU��@�9�O���x�^�������}�j���b��~�����_�l�ֱʏ�����v���UfDmUz�6��=��a��W�ǶO�Ñ�K�U�����O f�ꬦ�����7�{�9Ƽl�� �`H>E��U��J�;ub��~$�E���)ٟ�ff�{Up�͒�ߚ�|�(�T"�A����E�L��5�G�3�yXC�����w���$zy��d{�^elG�*��:U
��F�� yW�|"KuĻӋ=�>*�ZڭR�A=��7�47��~���Z�k�=��!��{�G_��ʙ*k� $D��5�r��ቻr%c�z']hr_��Q��>B�n��G�x�NW����@�sl΁|QoD�Eb�[��ڠy�C�fW��FDJu�V��<3����5گI���Y��|;�IR�雛���I��Ǵ����$���'E*�ib.Z��U�5�ʟ�~�����@I�P�	5i�Fc�-|d���y�}fI�E��2a��'�cg��N)�����n-^,`����m��}�'80N�h�2;R������r�_X}v�vׯ��pT�/l�'f׭W�+/D �^OM�p��5���Q�KsV�RI�!���]�7�7G8�*�f.�й�e ��S��3����Z�x�Q��~.��Ҟ�V8C4�@rV�SS{\��9f���z�1�G�W�>�Ղ�kʑ����\���a�n���F*Q�{�j�[#�t�~���ö��;�꼎k���OG�hR�T���d�^)q�{=�W�3=UX�s-��C�Mz�9�q:s�R��x/�U{����B���ܭޜ��y;+�9f���c|�s�c�p2s�2����ե��-���b0��.\������=�:�����4%7Z�^ѓ^�>�d�?�lφT|&x+������C�s��W}^ש��c�w���y��	?s��?F�~4��\*R�q�E��%W��.:�F�u�h8<n�qs����9��:'����7>������Q���v�O�(����>T�TʯK���*�[����\�����q��z27�>��t��Q�[�l��Rx�I�0�O<#z��#ƞ�X+�=�+��UA�Q^�\In����3��>�21̰�Q/n����Mv�~B�#�=� *d��}e���Q��k�O�"�3�+��ӡ_��#��[��&�w�g<����W��K_F:�]�V��aNK*��;������td�|n�cJ7�c��k0&0
8��J\E�̽�;�����߯�纜6��8�t�����}Y�t�5�-�kY}eȲ�C��;},E�&L�+�U���뛫��=�UU����)��?�dk�A�I)V�W�� �Q�ʣo��m��N������Ϭ��ku �ݨ�}h�{��e}�_���r�Z�z|5���Pt��x�"ǽ�Dd[#����}m�ҎU���ʊ>�����ꍁ0�Ԅ=�f�[f�����kp�h������q���F�wG�lsb��됃��n�O�|�|�0?T�6���!��������`�Y0ڦh�O�?Ob@��;}徸������{��8�вhW��,����3}4�pϹT�ߤ+!^�+�8�|��H�Kν��K��9����F�*�w-??ߘ��(�L����+�/��Kƾ9<����ꬿU/�㑪_��\���S_iq�����=H����Ł�R�J���Y��_���F��c�?N�q5YgFT��M�b����Ο\��y���=�U����X�g�F��f����T�����3?|��}~��.��pޯ�s$�K�z�t{����L�y��W��=~�]��劦��~�du� �T����(�0�*q�M൹�Y>9x,�uԟ��s��m~��gQTz��.PN���!�<#���M+����R�`�6YVR-�͛�q3��5��Y��߮��D9x�8,\!&h�l�������r��n��=�|Zч$�}ORm���Ag�0#s��3���������4��E�z|��}�W������s�B�E�t�ĔWh�~+3'��n�����A����aug���{ND{����uǸ������U�gH�z��خ�/Еy��P$��`{���$|5ԟW�'�ӿi^#��~�><n�#�7�_���M��ߣ=�.��|j<��!��PK���ץ
Q����S0���z��|���oBRt����ۈ�S1N䲠 ���C{$>��9�::�qn�D���J.���:����N��d{��M�{޸�>�LN�%�PC`�!O}[D��H��.�"��+�6��ė��G;ê����޶2=>�O��t2o�p	T�'�'���>�{[�Y����̥V�c��J���z_�^%q��3	�zKn|�%�5�h�1ccۉ�yR����n> ��(�����B��g��/J������Ғ�������tځJ��4�V�׻ه��B�\���"��=8�]{������>��V!���iP�z�L�O�����X���j����S.��H���a�$�aZ�����q�;�����%�or]*���Z�H6���	�y��MGϺ�]�v!2�C�b�@P緫.V��.��K7�QGh��x���+7h\���+݇6���EwH����Tk�6VO�"�mE�MW�tb�H���<���ß��3-���)�u�C���dy�{�8�U��l��J(ad� dw���+�U}�*�����7�y�w���G���V���~g��_G�\����i���{*E"�̸3��^�s��ϲv��oF�7�m��r*g���5�/?\����s��C�q�Gd=��9'me�#�X�E!O�MÛ_���X��7��:��ʮ���>�q���W��}�Ⲽ�:�,���Ks�7�ݙ�juh��F�H�w�L�z	�q�U꘸�U(ޯU���^�>/��N	Ѕ/Zر3�w=��j6=�nwjz�F�F����� y:������ό����?=I��eD�gN߯�0�!�����ǶO��ʡ�8�;%D*�,	��2.:e�6߶�z+��r*��p��sk��O��ў{^eo�Tt���4�T+�%�>�~{����U ����GW<��O�&W��Q���+��O����k�=�O%g�����+�H��a_�~�=S=�w��J�t���V�un(��t��(�2���k�yH�)`��a�j���t95N�{us5��}<囟A�v�k��宱�l���r~[��(z������ˢ�X�F��u�(50֭紬M��9cۚ��_u���}�AJ|2:�"�~����Tk~����x{�#ӕ�o�:�7uzc�Q��upxޥ/��$�<fy��Dħ^p��<29K���kj�%{��O��
���#�y���uJ�0���@��צdT"�H&=c��}*wƆR�i��T���ǟ�:���ށ�����5/]J��O���-^�%���͍�$��Y=C&A�������x5:۽cf�3Z�9=���3�O�r.1���n=��<���53FK'�d=Ȝ�9�ʦV��wR�v�����?շ?���}߾J�8_ݷ���y��2����<n=�C�s"�6Y:r�≛���9�
Ǳ�Z�g�U��e�'�N�R�{iW���W�̿Lw����;q�z���"���Q�9�5��v@L�.r>SV��=�<VL����(�O��ύ��4֚&�=<w+�{g1��D_��8�����i�ӷ,d�du׬�ȩt<�6g�^�W��g�z}*4�~��}}	Tg���^��j����q�g"����B�5U}E
�A��I���2R�0�:gnG�F�K��餅��ިܛ+qRݑN�	[0�ܑ���;W
��^ب��=���;�[-���n��^u��:�:�J['r��Y��-�Z��⏓WO�;��2�;�g�n%��^�Ǫ>�
A�ny-Jm	T��adl����vN�W�/U�G�zX��S�Y�C����(v�Od��d?�=N'9��?o�f����_H�]�̹�?:���e�.�~����FF�'�;�=�=�c�r''��rQA�V�����d]z����ǯv1nJY�0l�w]���w�����r<���dG��|n#ڪF۪aˤ�ps�;�o˽��FZ'=� nj$�+��o��^|��r9O��o��H���b=�:S��%(���.��u�]K��#8���AF�A��D灎/Ō�s�ޞ�׭���gB�{{�7~cP�ʷձw�Ä���!:��W�b�s%�a���D�^SB�:^=�χ�7ݧu�d]i���3�S�/ݮ��O����������ԁP���L/A�1���EO�`by�h˭�<�J��|�o�x/Gy܏�U#��x�`���C��/�R
,��C�['�w~~�]|���9�Ƒ��J��3�~8�{u��j�/��JM�� ����}�j�w��~�?<�W��oE�nRhO�9�|5�����~��r��)iy׷!�]�ȍ~�=.s��T�u����,�B�w;��v��� ���OL��3&Z�u���	�ٛl	���(�a۴AU�n�C%t�{�+XX�$�����C؁��Q�����JWk�8�nj�9}�@��� v��;7�IPDe��@���&�����&s�>�CӶ���k�z���YY3���,��%�cgC����܅t��7�����Φ����F9�K�
`���B�my_���^���M�c�͗�>;;q>�l�w5YgFEJ���}��<��$]�H�>����E��1�~����go�Fm���+����^���^2T	�,Z������q�N�&�V�%*����'�����ddS~��^���t��Ϟ���A��Pf�l�i dλ���/|�o�}�Z��t�@7��B�>��q���Ol_���+և�ϧ+���h
e:�>^޵��t�I6}'<k�.�_)�E�]U��m �F�_a�}�~/>��.+μ�XߏM�f?��ؐ팥�Vs�^�l���J���X<��u�g�#]���zhV���r;�<_u�y�G�γkn�}��G���^���e|ZT48<��B��7�l�����>����c`���A�Y��^�'�p�Gwz�>D������Ǫ��K8���|}DO�[�#�^s��=�t.�����lr�zE�7�|��޿�z�q����W�%�Y[�t'���!�lz��=z]���0��¯�f+��z����g,��%8`�^�DC�ܱd�Q��軫�� �G���,�Z�pO+��ݍ����{�G�{E	�j!�W�f9ԈԞ]�#汧Gh�i�c�;�zq�Jv��}��r�ʚ[�R�����\Ԥ4�t*7Gt��=Q����П�0�>�O�<gC&��@�����R��P�s1�b�+c=�~��t��&yW��)cj������j}^��{ԁ�}�^ w��u�H��{)���r�b�����+\�����' ̶B62"}բ����Y�R��s�\{>j��^&J��U{i��k�{���o�u�#�v*<^L�a�;%������w�����?��7��Y�rQ�������+�^ө�T�>h����o���M��/����D�j6t33�8B�H��g�jV^�*c}��8���̟���(K�֫ޯ,����^/{�`���*��Ɩ7l�/T@����,���.��ARU^�>�*}\�F���7<��W������x�顚w��eH�R�����x�x�{�kOB.&O��Q�[UǪe���k�
��쑑N_�&}1og�N���y�k�{�����4�m�IQ�I���e	��$:�&�+'�8X�#�E�d��S;��<��q�>\Uv�o��Ԩ�C���'W���*yu���%����j�:�K7�V|;��W������}���e�ێ��>��C0Wo����3jk2����y����^�,�`��D�O"ݝT�J����wnѷ�5ˎa]��kRP8���*tX���������:i��u���J#˞ƻ=�{N�s-�)j���W!�J�T�ԵOw��z}Ⲽ�<��:̣�nH=QX�bⶹO�����wy�"�Mh˥���5�'��ϰW�+��C��纏�_��=�g<a���|��(�22�e�\�ts�EO��+o��}�P\���GK~���V�QҮ=���r������Q&g(��Wg�i+d�:�I�3�/v��m���_ޯ,A��#�ޤ8�o�c4}T�V��[5`���}Tm�]��#�� s5���^��8�G�cQP�
�����r�x��cӵ����{]��=�3s�,��u~�=shω%2$�e�&%����t�����#Q����S����K+�\�	N�_�@C��َ �8��3!zw�3�V�x�߲�.5�r��8�=^U�m�{�n�=;7>����ɋ�~�&�ޟ@�d:�&:}fI�Y;B.C�~D^S�>A���6��>���g�M�䩎���}	��E�?P���{��z�V
�*A��O���)b��gD��fetS�zY�������E��+��}����ϸ���������<}fFG{*Fo�Բ��fvf���a-�J(�Œn)�f����[�1���;r��󝕋�h'-y��.m�|��=����{o���H^q1ڋ��C�;�`hs;�ɒgq���ou��,3}-��^�א���nD#�"޽�;Y��{u�{�7�rg������ۏ�}���Y��[t<�+&ܝCb�* �܂�%��N�c6gC��U9�9z�v�+7�5� Ѯ�jk!{b���������(2�VА�˂�}T37(W=9�G��z/����W8�M�AZ7jg.h�x�VVR�Q�|ԯ����q�c
;
n�z���Eƙ߂B�0 ���_j�Oj�e�,{w`v����,u������nC���QW�Ce\��hX/�DJr�)�lJĹZ���WP�w�r�o=)��z��U,�o)�-������:�G[�jE		΁:�ˢy��r=�]ru�gV��:�����[�/{���n�\�-9��{��Wr��#�����x��*�v�/�o;Ṝc��I]m�u4���%�Wg1x����㓓�$�z��t��Ir����no7u�����I�-x��,�@�x�@S���%�b�.�Tt��l�����,EWR��vum7E!ĝn6�uT��X�y��ݩ�Vj�f��N5��.�Sw��˷vDN�D��|�З�j�A��X�)L�WغhH���wO�a:�ͪ�2������ 1��9/(�#�z���c�Pkd�����c��wgo�$H��t'h$K�{HS�h0R�}��ɾ9��R�Y�彂��e��\5�JT9�O��mB�Uh�Gtk�q��c��
��[e˺:�`ە�뫏!��b�-�NK�Y|����K�
�H�$o�O��g)�6ŵX_MpO��r��^�)����CZ������o��� U�Vȕ��']�Pc��I�\�,�x�m	l)�}fG�C��m�F�쏳"�QV�������Y�]���g=Ԇx�k��}ڛ ��b���\�S��_�j5�j���n��YI@s���q�4��^Gzk��Q��{�P+��F�݅��V��%���7,�vI�w	J�<;I����͵�}Ƭ6P�BK��gDV��q�������ԝ�lv�Z�WM4�U7����q��42(�D�KW��y.̋{���N��2��{b�U[���٥%՝��\s�$��.�O[m�K�k�ѕx��3¦����5QOv�Ы��9U�v�թ@f�Wn�����!q�Y����P���;w���.�w��4\�N��CQ�M$sZ۝��ir«��i���J]��8�2SJ�E��%�L��6��p�}�Ү��8�ttf]ok��7��Β���)q��a������S�]y�}�Y�c����du���vg_1
˸&�h�I�zuV6��Z{ج�5f��}u�_���o�������~�}�U�+
�V�D"�"�*
�*�Q�U�@Q`�Z�U�
!DADb"*���R�IZ°EF�K�EX��`V)X�b[F�V�dbAb�E�d����b�DEY"*FՊ
(2�P+D+AH���c"�Y�Ī�(�*��EU��1�bb�T��(�b()XQ@dQZ�
��T�2�`�0(��e���\IE��*�YQEV,U`*�Q1E\��5��U�U�r�V8�DUT`��V�"1D�S̬Ub�R��T��*�ETDUE��*�AEL�-�EEE��V��V�b�$�
5(�+DQUE��6�DH�b,DPn\X�J�`�X0Y�"�j(�QH�U�
���()��Um�EQb#iEV"_u�����y�t^���g-hu4#�j�g����2�O��g�x��Z�j�n��U�F�X�Wyš�N:x��-��t�%B���&.>��s(|�5i�S���Q~;���e���B��:�y^U>gE��9�6j�{�W��X��t.t;�&��J8K�}�LK���t�ԕǨn\яz@�q����bzw�{��7�l���^���ˋ�;��^��"���ٟ�������n�UxR�xpW�>�=OŃ�^������:�"�n�
�,��qb�����eg���&���I)��La�qUa��|_{G��Ͻ�~+"+ԇ��1K����$�|f�WRJE-�w9�]u���˪���_���N�C��ё�x�G���_�l{�D��QD�8Ȭؚ�Hm��qt����$Ͼ3�1J>����A�_W��D�~Ӟr|��D>7�R72+�����g����{�z�v� ���u�o��[顨�~W~�ZG!����zZ�����Z���7����m�zk�î�}
EI-�c�����7�Rf���s(EzyurW�0��ǔ�3���n#����Ǫ�d2KK*�U�A���~���.�s�3f���W뢬�򛗮�mP�p:��ڗ�-�����hq�[�.ߙ�(�U��o��o��n�Oq��"Y��J)��|���b�wP/�*_���:�^��<��7g��7,���I{�xf�i��Ӧ�M>�q��j	�d�.�$�	\���x�;�fk�3����O���%�Tl	�ө�R���L����͖�,j��GY �
��O���%wM�z�=}�r<-�]ȿ7^'�=>��,l?]H5
Y<v���u���Q�{O�?]
�Y��d����=:�����ɼ~��{��8���>�ߏ���}�5�f\s��H4Q/��ql.�[�u�GȤ}��^�<o�|s_�K�ō� =��B�U�N_0��zz]
����^ρf�K
4�}U���h�{��ܮ��3�#as�T]�k\�:�������U��~H_����?��(q���>�l�fg(蒧�9t��;�|&;�k���˙�X��#�>�?_�ȯV3����ﺷ�V{*t�"����|��=��J��~���|u�K�|���h�5�����߯��W���r�i���ӶY>R�^���A���e��_T��r|e�z���tn���}��bF�z���N�����^�<D�p�eft٬����L��G����'MI�4eT;���Qy��f�[����^ӟ{����u�򓬨~�o����-ӃY��Z�m���9�Ӈv���V�4*�#��3��\ډ;</�����w��Z��Y�dC7-�M|/C�+)�-�V5[N}��^,�{���r����\��5Z�7��K����W���0M\��r�ޔ��t����NWp��|	<K��C��φ������U�N���poQ��d�/���?8���L&��~���6˰lT <��`)^3qe��C��ه�Kf��uj�-3yS>�[*������w�N���D�z��qD��( %_Q7�E�E��6�&nez�����y;�<�Ԇ������ίQ�.&����7��D���e\|����,Gb��Y�Gk�$��eR�?nC��C�h��팏O���ɸ��v�%`���^�==���[��k��f�����F�O��ϒ�~7�f��5~�~���� ;��T��:�f���o�X�]��UJLקI@�§}:*nW��\�����򪒞4�����7ihh��2Wl����}�&�L2��K@��w�].<2��������ܺ��$.��}�5�}�%�X�𤾡�{�rsK�8o�,�PɆ�gC����v6��]M���WMy��xz�n�xd'^Y�=��@��k
^ʜ7Y;�ay��N7��z|(PQ����5ei�wL��%OgD9���XD�fY����Z�	F'H�O�{ M��v�Q
�KG�b�X�xuڵr(G���"p���6N6e�������R���؟a��
����`���f����-	�`��gH"��n*j��i�Z��ʼQ�e�#�J��V���~�|��?R�x�V;�a�ўʑ�5����73f�гz�D�z��_�G�mW��x��| �^~����r�Q��<�p]9�eU����h�����פ{�nO�Oĸ�&~�Fv�-_%Ez�X����P�o�����uԕ$�Y.�j�N���Z\n��U��m��nN��I'��>�D��CUW�!N����P��	_���v++K��ݝ��,��g����3�i�(ݹ �`H>E���s�k�=�;��[���BnzY����W~��=LnG���\G��=�ߌ8�QP��*��qS������^Q�,gȲ{T㩂�^�p�q-��g�י[�GJ�mtN:RYܪ|�\��Gv�Z�x@��=��7�/�����W~�,A��#��z��n#��ڄ;����������\�SQ�f��H�n���-l9�E>B�[�6\A��x������2��)7��ʴ
��3Jd���͞�&_�
���G�B/���F�viS� ���z�{�8z��Ɔ������<yn�*���ھ�6Ҿ���ޮ��)k8[�H�]�$˷��F��<���\�un�_^��*l�)��gosb�W]�,k{O��DU��5�FR��nX贼	�f�VT�2�CsA�Hf�Yv�9W'�O��d����>��ց.i��A��30�
ldK��e�\i^_*wX��6��]�����V������T�����G���>���XQ�nd��}p'�a+V|W����#}�am)�1�n����j�C���\c�L����*�B�ו �d�3>ݚ�j;V�z���B�@����{�"ϑ�J�4>����꼎�H��U����	Uܺڼ�yQ;��U�f�{����@89;���������/����d:��9�~�^rҍH_a���=kҨ砯<�F�����A��w5�|r*ex�t��y߀1�d��v�=�J6�qW�����3�n�B���3�x�8�X�'�κ���K��==\����c'���f������NS,W���E5q���ι�4>�e��g�W
�æNz;�t=���:�>Ȏ>�7��B�h�1��?>�=�ޘ_.ʔn�$�{}����G����d��/z~�G�X�y���[T\C��!��{ף"7�>�܏u�c�M�	��%��5�Y�#o��xԴ+�Tֵ�m�4�Lfju��ҝ��[�.	�پ�r���>!�<��}k�3���s�G�5�������S�	u�j��(�H�u3DP�8-w4Y��h�Z�omWS���FN��t�y���1(�.�n�)K�Cx%���\/>��.�3
�*�R�k]�����n[�i��s�����	��Æ��S�7�k=#=���}P��$1e��7q����c�ȧ�q7���\�ﱺ�D���
=�����Ӽ}	Iҽ����f��,҂G�E�u����/��Gc;ޚ��OU�����z���ߙ��N�����i7�z�z�U�"��jo�S��"bJ����K��9�2�[�T���Y�|��=��ۏ5~x�Q�~���=Q�'�N�
�,��a{�(��qp/L�뭥�&Y	N��r��V9W��#��G���~n�O���w�E�~��w��v*���u7�Ơ�I�b>��QR��N}[)���|y�k�C�x�@9���i�^�=��s&�ߵ�{~C�Zʐj=>%���������=�/��pwO�P�X�o�2%b���M,�fg�M��Չ��*n}������l�|k�:EV_��+��G;��� n'ϐ\�r���)��:.ס�#jk�X��������q��M3���M�_���,�&���G�U����i���R�2�-��y��Y*펰���E%�����B{Ʊ��nЭZ�u����Jw�B�z�\�SֻY��v�3 s�]AG��s�^'�����r��37��$h�3q�^��ټf>���Ef�ۧ8&2]�Dz����2��sb�sPU=��K�G*`W۞y�W��M���ޫ�[�+=�:o�Y;�f{��zaP��9~����:=��ٓ����-��߯����~+)��>{<3�gHW�ª�fxy��z\.�"k=cpџT+����t|=T!����E�������R�f����{�^D�]���P�ByR=\�O��3�����`���Aߣ~����'��[r9��~ճ�܍�B˟}]��'+���U
|	=_L�$yT;��l�dk�>7�U�s�����iG���ҭ[9d��~�~/M��O�P�����@A�Q��<�`\+�o��X�=�Uw!� �л�i�U�F�R~�Z2�[G=�I���g�N!滋B��#������Iw����6rmG����RG�2es����z����2=;����������~�TMC2YS.=黐4B��V��5S3�|LL�^�u�E��G;���4Z~vǏ���:7s�Z��{�`����oz'�,�P29��=$LK��E������;��u�j�&�=�R�����~����of��n�ð�9�H���a����2`��l��Y[��c�0��"���o�vo��SjCgo4K�or�w�zZ�5ú�$�r�5�w`+��,�ĸ'4ͼ��GbN����d[J�E]�a��^���d�$��0B��?���wc���r>��ꭹl ���L�L��Y<+�3/��*pT��VR��9��~�>���HUv�D����;����'�g�L���@w�݊�>ɓP�SPrX���:�q�\��\��R��k]ߩ���.Y�'��}׈m�%�c�O�y��Pu{�5�ٛ+'�2a�ZhQ�c��!F�7�t�m�=��D�wW����G�Bu呯��)���[6$b�T�,��|��*�&'|����oB�D��/D�_��Ɲp;�j� ��+�s>�fTC�/�47Ov�B�X���ݛS5}��r+N���1�jU�{w�I~%��5�Db��Hȧ/ޓ�W�1�J�L��]v�t�j�_���X�{7'��~�Beك�:���TP��#�s�P7��D5C���� 4}�׻�F�Q]�q���q���B�:rN���$���=�yu^���2ʸ~�=ue_��S�8��O�(ޖ�,�>�z_�����3�i�(�[�TA��>E���3�#<�C�L��J����Qf�~�mz�8dyS�������9�(�r�%ct!�8�;|g#&2gR�@BRf"�FVR!�^X6���C�M�鿴n�1Tv�� ��f���&Y�O�r���5B���&�4��&��A��*�K���1 b� �b���լsWh��.�������Ӌ�2���K2�eg��i��q%�Ig������zu���{8H���z3�k��x}�p���]� ��c���!��/�3��R���J'�t�#��< ��\M��+��Q��>����3��u{ԇYP���`ͽ�{���sԺ��7�U�k�L�4�f����[��-l9�E�	�Kԑ�2��Qd��g!���Tw����Nփq�V�Nm�D��D��=$�B�]4xv�R�IÇ܄>�=^֤N��}���n=��'�"=3�'��:�&ә�Q�,��A��뀫K��j^8�`�s��������^J����G���w&<ߨ�_{�����=>�$�Ȳz�0����S�)w�v�+��u�g��^�y�uxu�Wzϓ�܋��zf���=*�B��H$F>�C���̯r�9�/D	�0�k׺U���~.;oo���:�#�y�㻚"{��ɓ�io�zx�۟!��ʑ��d��fL37^�Խ'�:_���}f~�3K3��GJ�^C��-��އ{>��uor�r7%X�pp�ٓ��55ii�T�|O2�ߢ���42+���d#J������YU�˗���4�f�^��uZ형�����5�f-���[��E���/*��q^�� �Ɔ>�)i��<fk�e��|Yܙ*�)١�d��*fʾ0��H�걙��:vq6����>Ug���Ωq<�%/����m�0=;L/���=��;�Y
��\΍�zN���2��}u�<+����}��5O��iJ�8�3��GL��}>�������z�O�Ͱ�8����("�����#�|⦤{ʆ�Z^�<=�]R�t�A����a��x��1G�O�dW�,3�au̢�1H��k��ww/tt>�I%}�"�5�.���Nl.��n�q�}z7�|�8�u�z��jΌ�F;��j�0u�j��+�@�:k�U|f	>T���'P|U{�q%����s�j&CfJ�]�[��J��P�G��T�s>�%W�@SRXρ��-��hj*��Ě��n{5���_)�x<��6�i��'J����m�i��2* ElD����[��K�cq�����;�u`�z���6}�f�!���ُ��/�=�����'�3�#a̖�I�㤏?J��<�[��M��n�r������|=>�r�6��W��z|���G�wļ�F��t�@������3�c�W �C���_�"yseєRٵʡֵr�ꈨiS%�,S�B@����$��$I?�! BIB$��B@����$I?�! BI�$I?�! BI��	O�H�P��	'$�! BI��!$��	O�! BI�$��! BI�$I?�B@���B@����PVI��uć�@A^���@���y�d/���:�� {�)!@*���P�R�  �(
�RP�(���WX P(�5u�%*�H�AJ�*R��TU(���sa`��U,��1m����mPi��R�v���8���A��  �  m`9f�T���UV� ���m,��l�]�j%*H�j���C�T$(�ۘ�ś��۸���gv�������ݷWs���ĕQR m��3[vd���.��i�軺M��s 3Mki�m���ՍJ��aҨQ��B��]�E��v���wa��r�sQ��������:�Z�I�T7w%V��m���tPviu]�M���c#��mE�5)IE�9�T����V�jɊ�U)�KFT
م�(�JG -�f�#k16��V��l0��ֆT4J����50b��%j��HZ�fֶ��б�\        E<2��P�  ��i� OhaJJ�h      �101��&5O��J����   4�4d���`F�b0L�`�Q&
(A3@���j~��5=FC�7�OOQ���}_��3���ٝ}�|�<�V�A$	$<�����P���H`�$��}r I$,!���4�E�I �C���	/��|?�?����?�/���|?�!���a�H"��	�I$$�J=/�=� �C�C���0$) P� $����������_�L�?��������ױUUUQUUQ{� SI)���BJ@$�� R�)�@�H $�$�! �!B�	 R"�I���R�R��*��*��*��*��*�����U���	/����|�1��믽�C�TK�n�?�C��,��I�h�,(�$^��~.oT��&��[�Ż{w+�A�B��.謳yvi�AQ��8P9t8��g,/5*=]�DR��F��6��J警2�ڒ���3���4��k�]/�-�lR	�(i;��&졢�V��7t�da�V��¡�gXr�j�
)�4Q*��z43��$aUsU�*"����uݮ���~cCN�N]:4x��֬�,J7�d��1C"̬�k�;I=wj�^V�С�f嘬�8���ȃyu]��aׇo?u��KU�w^�]��M���֛r��Ɗ��2���'�P�'-]XuN�j�ފ���BT�^�R�C��5�c�iY����H^�܊�Ů�k�Mnݺ�ͥ��T�I�`��\ڂ$.�,{��%J
�ѡօx��/��{dq[f��O��KK��"�eޡ���Q���B����{h��rUe�Yt1"*7��WX�/=T�����Y�U>Wc>�qi���'���F�mSk,-�&!kف\XfA��M�)��d���B7X��ɖ��f�v�[c6H�:�I�	�qVڭ���ceԻ��&S{��w&hŉ�Rh�윭5*�*�.�ҹt�|�{�-�2�|�}���t�QC��Ƽ��UML�l]1%�j-3V�|B���Y���i.��ٖ�YտD�a���I��fnK-�3�tQ�0݃L���y7V��&Y���95���⬺�y݁Ri5�om5��0���{Ȧn�������&��tw�y����غ���8�81+͍�g;��6UizF�#i[b��٫��)�YTk%�Ԕ�v2A���v���5*����۵�sUr���WU����TA�v���i�ꩇ�lŒ��U7�x�3�57v�ۣ�UM�?�
�����%1к���u�X��+�$Yyo^�M��@aj�ԭ�6���k-a�1�B	��RӧlRi�y0-�z���Q˪�Y5�h��qѥ������ѩ�X�Rk�-�Ô���m����;�*����q���:��]U�	�j4ĨыC����Ec�"��J<�O�V���+��Q
Ρ�֖FU��"��L�Ӳ�1uY��/l�m=�r7	5tie�լ�%�6i��� �%�w��$�3�I�t�J������.֨��fЄJ&�.Y��G��r�I.�l�\�+	r�Zܨoh�ٕPځ��Y.�1O��7X�+��h�O��K�q�9-8��H,ɹx���V[�H7[Kwqͦ��X�6kjQ��>fGX,��à��orU�i����X��z,��¤od�c+6�ō��2*��9�Q����Ve�w�UA��*�r��B�Z���ʁI;����sDV��Im�C5����������M��ָ�Ud�}Vkp��n�<��;%��!K.��s#ECn#�u:�ө�����Z�ӫf�ܪ{��6��$�W,\�${1om阷�R��S�`41����,Ҥ�k%��`�Wwo*�ZĮ]�qʼ�r�W�kNR���Z�;�Ռ�Z���el5IS/^'��n"uT����n��uF�0j�Bղi�0ʺ&�M��Z�G9��v��đ�lk�'�xAz7[�'���9�U�tu��E��Z6�\y@f](lj߮�8��$��`�,�Xf���MHIV�i�V�F�B�Vہz��DaQ�a1^[��]^d��3�r�I�Um���m�����@H��P��5�"�,��T�7���� �X:i
��f����*��e;�G�ET�F��퍺ݭh�az�*���f�ãU��j�j&��]n׫Cw[\�8^.��ƭ'gU�t#,!I7�%Ɇ-��k�\��� �1M�LҶͩ����T[J�6�Z5�P�U]n��(�޽n�V�����V�hS%m�#��jӪ��b��y��un#t�Z���0�yn�$2�2V=��5v�7/�c�0X�Dk��.<���픢�d�2�P���yGH�c�j���Ǻ[ֲ�e�*]�r��m��,u�������U-w2��{w*�yy����klͼ��kqԲ��Td�݋R��2*�RJ��+�,Vo&��%嬺7P�-�����uGSz��~��U-�Q��bF�K&���T^����b���I&��i96�][6DD�5V�ĨQ��A�A
���S�xX��cW�����l/!/B���/iԺ��[{B�bEl�J�9�d8�[Cf�t���	�ช�q�+s�[���(��֒��~��&�Xvf�`l�gIxVUQ�WGN�`�����<�ј�A�$M�l'F8-��	8��ٷu��+n�$\�h��-�i7p`�4B-�r�m�M��z�l���A�U��cd3L�a\�&v�j8Xe��9v-�牆E�YI1D2��<O*�WɫL�gcW���4�"VU]iR�ӫ��w���˪CN%F�6���Z*��WGN<.�R�N�m1���2M-�e�>W���Wy��5�RdϚ��Z �: �;��J[Qhn��]�Ա�`�P��m�kRܗNbrl��Ȉ��@���c2c�6�;�т��e���Ӛ�ɱGa���I���	�0���ӆ]�B�>M���1=�@�d��{�h���9n��O5ܑ�9��Z)!�	C#g�2v�F�(���	)�h��S��F���t����xk%������w��Q����!��Ͻ�}_�F:��?w���%���C_��࿏�)J���p}_���V}��?��2�J����mI9krA"ʹ �:%Vཚ���Nw{YP��_Sw�A]��E�n���v�InK��T��𐍹6-�&1�L���N#��g��Pv^�˛ñЉ�d�Jߔ��\����ke�R����6�U�d��q�֮�U\��{t�Kr�>�PmP-#HgAV-�+���25u�}�f՞D0p�y˹]m��Z�-�:b�71:������"�,�ވ��֛�ϮR.\�����\;\�3R9\��|�!�'�����u����4�.��@+N�Y���ŕ:��9Z�;���u>峆T�/h�Dc���u���t��8fc=}o���թt�t�ո#kq�:іa��l��Eӳ�㜤�s ��9y�gN,���X\�V]>�M�T,�6giھ뒤{�Q`

���\U���;OKh�Z�Iyµ:�}U�2�H�T"���S�E��/_�[ٲY�f����T7n=�Q�DǦG6hep����Oe�xMK5����7�*P�ӥ�}�kn\������f(%�u��E"�}�D���f���6�xw*��%#H]��f���Q�_#�#�ˎ��6j�՛3u�N큐&�+�gw[���]r��5�3Z�t�D�ǣj3��u^i�Za�
���F{4Ce윬c�K��k"�$���G�a߰nҘ�;'a]�k��'E�L�*�P(vv�'.��Q��g�G��Zl�wa��n-�E��ʛ�T9ѫ|�r���ҙGz���y0�TPt�R�]��ei!�ty����z���[�-��_u��`�
K'
*h��^(Ú]u^cޒ�"�e�+�z.o�}W��]�G�,�����6��e޵�Y��Gk�6����/M�N7��P��Q�53q^���L����9P�-��j�Wd7[2�p;l�I�tud���ixپ���Q��]�J�ϰ[�I���s:�c�P[�J�^�@�5�=�W*�BO'������8�&���������QdVr*U1�����SPa�^:�y���,RǳzGh�!�nJ;:iZ�; iu�ot7[�QV��_es{�y���˕}�A�3^�,�4���VMn��{��7� �ʷ������R�nwk��ʠ��-����D-�X�	G�i���s)9P�R���x2{�ee��}1�Egec�%`�°].�eB��Y�D;��oEF��N�0@���e�"�3���4�I�)�j�d��]^ul���+��Y+�6�q�N��u�kBu[(�q	8�z/1���:+��zj�3��=����NŬ�y|�tY��5��%nV�-Y���V9��]o���D�V�d+}�zx���#�zģ����P��rrE�W���$�,� ��u['i�RYD2�}�l�G�;a�*z��64c��]��T
�BkӺ����b����9��e0A㺊��K�8����{e���x�� ���)�k�Þ8����Nn&f�G��륧(��@����r�:�m΂����ٔN�#Oq������\��WW��9YZ_u��FTu�Ͳ��=�eR�Y�c�i����у�Re�.䮢:ѓ����qN�:����l�OӖ�dK�/�c��F�GK� �Si氁W]Q��c�x�����6ܺ�ַ��*�	��BM���gm�`Z�f�֛<��/ K$�ѝ������Db���9�ԍ����^��@��uk�m�F�QG�{�(��*�eiW(i�S.ZC](�Hr�A�x��wQN�
lIgs�Ng+;Z�7�]�Q�Q�'v �S�gf��H9X�b�-A
���%ݞ��*33k_�+gt7[R��%V	��^�Q���sM��6��ޔɬ�Ӻ,m����'�4imm�{�ۺ/�$��Ήol�x��)�}��(6�l��k�s�NZh�A�K�q\��2Ʈ�r�ͧ
j���Z����j"�0�=�;	�Ƥ�v���vr�S�;��HjB[�.:|��Q��*nLy\;��G�c�(����0��z��A=�j�ӯ����r�]ħ�eϯ����Y�1;�-�����K�^ܪڠsh�2Q�tQ���#NF��2��q�r��eO��;n]mN�7_;*��k���0Hf�%8���b�r�SХgT�n��V:���w3N�3K���wjl�K�ʉ2����&wEǷ��r��N�v�LaL�`t@�`Wu�JX�s:�ƛ���Y��2;�WIQ��Tsd����Y� ��"3�ɰG�����t�SjGӒI��GQ��m\�1VЕ{��r�B:t�!RZ%��N�Kz�(��a[�αD`��ʛy�I"�L�RT,��N��#�6@2qRglNI0������N9&l�18����$$̠�ҽb���MV<��+7��/����/y�S;{�
G��h����%��)��74�jM��̵$��r.�%�%��)��#��$�ˇ��|�ɰ��Խ�+)+��v\��u:v0��3���5����jX�}�G�r���#�	P����j�AKq��R��⬣ �vЛ;1����d�*�Sm�G���YE�.�K���4�G^m�n�[4&ۺ-��}�����b���k�|Z"Z�Ŗ�S�E3d^�&�����;���Ӝ�9��_����{=?"���|�>F�/��	$��pqҵ��<�$ H�~����	$�����R�?pL$����3��3�>���}H�3�Lf�vnK�,�ϵ�����u[�n���@�m�9�#�2�H%�uE��̭s�7n�*�Rj-�����+@PU�uΝn����PŴ�tt����釯{j�O�u!J���qv���*sklhcq�v�*1�ˍ�=��Ti=�f���FY�h�n��GH�m�K��]�Z����X��&�#�MliD��7pod]�x�����P;\{@"��'m�9�]e۫�ܭY���;��-#�	�J�71$�$�Ԓ����I ���I�����2i��ᡋMf^�o=�5i:�{[���L�w+���'���G��%U7j�7�]���ˌ��KoK�n}�nv��_P��N-i���gUd	-W����`�c���M��+���LN��D���6����*�v��Į��$���T�����!�MZ�z�Qq�~�U�n[Gb��H�<�k�u(����D�{�N�o���Z}'IȻƶ$�m�#eR�/6!Q��Ƀ-,vo>S�ݹ������T�I$���32K�I$r\�I#��I���9�b��L��8r����;�j�b�ۚٺ�k��F�ӎ�f�	������Q�����K��!�&�bL�ͮں+���&��dݥ�,xj����v��̗�'��=���J�&�.ͪH�m�S���cy���&����n��uN{d^��
�j�Wv�6QF�2;��Gz�W�ѱ�ef�jCX:8����ٳ)h������SkbJe�zq�9e��nQN�����Z�J"�%K�����gS��G6�t����68�.��H 뽁g�W<BR�y�:��7XU�q�;Ε�Kc�}4)�v�������]7�B�Vk�(��(^��]aX��F��W�Au:��9e%ݺX�=of��o�mVR��ik�����*�^݋�B���qJ����&.��Uw\�2� +��EQ)���u�9!B,��fb�k"��/�����C���mv�&�.���KLo���c�a�z�a{Kw2����z�Q��Kt�9���"���pJьM���h>�5�'�T�#�ИM�{]n]���j6
�`��lhQF��l5�;9��|�/��j��S��5gC��F��fS���x��R��;��ϳ
v�;�j�D��Kj_�BPZF��e�;��y��m4��3+)T��i����0�A��2Vmc��Mfe4hwrek!�+��[�5���%Tp�yTVR�j�oʱ\�i��ӑnd<,!R�K�m}��j�^l���tt�뢺�-�Vřp��wwB-T�y��k�Qmte7��2�[K@�!�G����LU]w4*�l��Yx��.j1��Ej���Ը�Mg0�P�IP��8&&n�5m]7Ku�j�I9�hs��3�nhB�}}����X{&h����In��%v�]4L���T�hڨ-:4�:�1��U�fѼ�ly�Q�]8<��Ѧk>;��X��mV^�i��t�C:�T���)7\�����u�|i[:����3rj��m�a=t]uX��M��
T�(����]��l�.��N3W|+l������%�h��7f��9��k'b*�<vs�Q��ӭ�b���N��y��V��I�Y�f3ŕy[M�妹^֜={�~�ңƄ����N���*�#�kK�2����8E�E,�1A��a��1�+0��q��Np+���1�N��i8M�.�I��*]WZR���n4�$�|����}ܲ�K@5m�{�����X�Ww�D�èd[F��	\�w�g��),tT\kI-��BZ�T��Yx�����G�I�Ur���n�Ζza��T0��nht/��s3k\`}����.�KҠ�.`���w�B;�@Y�{ v{,L�,���oj����a��K�dg��Z2^��6릴�6�*�UU���w�'i���>&���P7����*�֣����eѽ4ى��#eu(�k��Te��	-i��rl�qҺ��;;���J�c�z���Ч{�9�&�.Y�[���VU��;B�a���h�QTO9c.�c�#���\��b�E�2�X�8�
R���V&��㳙)���sh\Z.I���F8��׹tm���)��gV��=�������
.�eo7A�^���N$�=.��:��Ηz�ne�T���Ɂ��Y� $bظkn]:�e��N'k��{j#�I3��������WA%-N��-�/�ml���L����+���2�;����*��U
�0,�jE���uz�T-�ѿ���gdL=��9���뷷�\��p\��A�k�Q�)ԥ���r�L���y��^�/��&.�pP�h���e憻M�{&5'U��v`TP�5�7Yr
���$	��ZJWҨ�K;{G&!KN8�x����,�$9\ӷvvW"�cE �ܙm�&�ܽ�,�}b5+*%vt�PkYݏ{+�βIܖ��s�(��lBmn;�{xpߚx%p�6-fiSj�V��*�Z�O7�Y��Q'�1_dnw�Ͳm�Zv�ތ�z��n�G�z��(��ڥ{�N�0J��9;�LJ�u#�\;5TY�c��j271	�D��pi��
y�r�uo8k5�6sF�n��`�s�W�ި���<m��O�$�A���+��=HP|J7A_�~��=�T",���+�,��X�p���;�_��uӡ�2�^��K2�2;MP���/t�fn�3��������=�"�&��P�ݧ\�*�r��6��)�Z�v�GV��J�f��d�Xܗ�V�}�Q`"Y��l�q*�J��7���PLإvʰ{�m���JD����0Dp.X�z��~���ù�F�zu���u�~�&f��L��x��=�+y�I���$�|'Tp��1l����Ghs`�´q�V�Ff�R�'2ol��ۈ�$QI"q�$�sN9u���א�rWN�:�~��]N�Q�((������JSJ��c=�\���R]R�X��ⱜ�:�R�U�N����kʶ ��*�0U[B�#e�)iH�H�e���ڪ���%!mUV(�.��
��-��QmT*�i����*%�BCIT44�m��ڨ�-�wB�K���7u_�=w�s^c�q��T�%�j.��تY��P9�6�nu}d��?�����w�m{�'H��rW�/mpw)�@��v��[�r��p���r�ڇ��<O~�x�~�x�k'�t�A:RN���1��[���`e�����
i��2s�f��w�K���������&�:���'uIuE�LP�����bU���l�����{i�G}S��A�I��� 5u��|hG�	ݻ�b�l����ݝ�a���L]��ݣ6K�s��xΗ���i��YM��E'�ꮒ,�^�¶\�n�z�O;^�"1��>)���C�Ʈ�~�g{;�,&M�6&�]���/�.��C"H�f� x�WǁY�r4!;����̌/��+5�Z�W�L#��������"
N W:�����L
�"�}v��������2�?!��~���j��p]�
LQ�{��뤷ɇ�Q9�TۙƟtv��
R�����g�޿*G�-����w����ͅD�2�8�^T�<g5���wi�9�uR���^��Y����/�2U{�Uk�o=��3��߇�\��fPN��w�����Z���6d]C8oc�\y��8�z�+��g�o+߮�"8�1wO�"~S�ef���v[�C2\�F�;�~W6�xI�2�7
y����ψ];&N-��Yè��&:E���6�.�����իl���\OF�:����b���q%�����ds�F��p4��'���������GM�܅�q7x�z9,f��0#�1����)�Tu�M!b��.����[Ι�����lAǝ��U/{|����'�������]����V�ㇵ	ūM�2����9��Ճ�/Oc�� �|�r6)�S��5��
�t���SjX
�L�Uv5K��������A=�%k�)�a[9��4�܋m,Je{g ,��D���*���9���X����B%#�!h#}�b,+���h�s�kL�W�u2�8�fW`�9���+G���K��o@�0�ً\m�ٟ��M�V(=�	dB]ϕ��*q5}� L�k%�ହɭ<��<hVoS�F/F�A=1��/4��y8���S��i�Z���s[��&c�Kߍ-6�}�K�8Sۆ���/��J���+�s8��sI+J�N�Uӵld�'"�(��E<U{�xJ�8�*WWV�V�=�W�gvӶ(q�k&��6w�w��5w@���+/b'؀��d�ę���=�wZ�!Ԉ����Nn��{oh��\�vN��L��.R�0�p(�����quv:9	��`����]Ke�׺���YF�<�u�qMU�U۬�
5׬���ɚd.k��2��F;�we7#�(������NVU���\��W%m�5��ME��B��xAvᠴ�������L�3�HRt)��HΚ�z`{�c��tʬ�ҽ���ɰ"����7ӻ��Q����쯧r�ւm��J��W��jw&���R�֮�Ş[�uv(��a�;�*�=�Ю/w7d���Fuvf�3lb��W���,�:E���2�G-8x�>�(EM11R��SHI�(�sx��v'�����맣Z�-{Vf��Dߵ2mVH���k7�'���S��C>����� Æ/z4�Huj�&��p��˗u����L+Wͦ}S��9����L�g�<�=Vk^v�����_�G�i�]o�:�ΐ�h��=�������J���9Fj������d=�g���.'7<������"���Iꗯ�ھ�4�s��3��Y�f%Gg5̵c[��Ӿ9婼�rvVvsի�)te�E��qx���0__�z�T
�Χ�[%���ފ�k���x�9�]V�[*��u;9��hPj��"T�+/c��ƣe���΀�Lp�ѥՁ��/��="|��p�*+��8����4��=��#9�m7U�q��^aܝ����m����u�.�����DnW&:<вy��᧦r����}���#Ȓ��1����l�i_uE��p�1==�O�7bGv���4�f�F�\#/0�|���>��'�x�uH|i��̻�I�u�#�8� i[��\)v�v����A鯊ɨ�kP.fl�k�]��vU�y_�0x�6Q�Z.�g[�v�S�ڇ7�=�U����&j����m]�n����� <���#�;�V�~�y�g�s{�]�2�.��q-�]�K�vRZz�S�u)��@u�y�I]7�Q�kN�.��]�ي�8Ó���8��}�j�7_����ȥÙh���7,� QxNB�N�Ȋ�PK�X��a��k��-<��5��֬�wDn�-EY+Q��*����C}f:��c��IS�����t�-�Or ;v7�ZY����t�V%Z�,j��em�j�q�o}�LYz8�/u����tR6�:���)nX��GP�Upӻ�ݶ��`��`6;�-�XޓT�nn���Z�蟾B<��NV�E�td\YQo{����W��*��Ğ��*�P���v������:<LaWnM/Cad@tʱ�D#z/�-LS�*&k%DΛIc��4��M�9�ͼ��іTt��KZ�W��mv�sV����-��@̱��ɖ0й�;b�iZn앍`��<j�ضIķg5к�}�J:i��O����PcZ���"u�J�dv��C\q�F�p���O�p3x�;J����I�R��;:(���c�&��8ےH��9ubSx�w�R�X�q�6���t<�
��P�DX�hF��yϡ(���af�����o:�s���J��*����`Ŋ���*�QTXYue�]1i�D�(b�6�+uJ(R�P�i)ʢ��m%�)V�Ք�P��)X����k���E"��,RƌU7Ta��1u-�	$�J���������j�љG�p������s�B�6��(����7�:O����-���?yd��p�辻�6����j�+�\u{�������}��^���TH�?K���|�������3�XL^�.��~/��f���F;"�c�޹�ZÃ�<�J��q5������ne�'��d���n�{{�߱'}�]�s'�qP��WMՄ2�h[~/Ƀ$��_s�ƺ��MMۑqƫ��ޏFᛯ��Y$��㳖z;�u|��OSrH�=N~��7no��ב"�u��Z�g�fNB{�6�tn��ݛb��T���xE� /Q�C<��[^W�����9������![G�]�'3-���z��=䷅�]������g�����]7�5o�
�Q�pAfB���ϋ�K��I�;���3�jIE�wz8Φ��'��5�,&bݯ�0���GR�9oݸ�aŚ�I�7r�Z1��O;�{�=Zb��j��V�P�Jnz�����~�^����wv��r�Z��UB���
c��.�5�5,�L���:�o�@���6�q>�CP8�����_��V׏�ʔv�t��[/��e�������`vV㍑Z�9��=@��~���+��y���\�������|��-��1�˭PW�<ɀ|ia��f�W�o���g���ή#��]�j6�nM{[����[g�/&�L\�3�r0gm�ib�ֲ�s��rk�'��K���� ��C��o$>(���;����F���_�_8���]q����k� �~U�Z0}�>W�g����W)5�bX�c�۲�o���<�[){z=/�,3ɓL��S��xz��Յ���o�(�=s9���#���l�� e��+�n��;$8n��&�cU��ā�Ru�x�aL��`(Cl�d�I#��w�;x��-!�d������6�<d8�m�I�C��!F��BY��Đ��~k�W��
�/���uO��G��a��jǫs����z,ƕbi4�F�ׯ��U�f)=I��]}_W]UW�@�e�$2���:ɆBa ev�l��8���x7��=v��2�$���8�m	���P&Շ�Cl�C��!�I:�ў����\����2��i���� �a	���M i�ZH�����y��=$�N��a��d�Y&�%�O!�2̤��!�I�='���7���$9�L��'1RBm�d�B��2)�Q�H
w�yy��q���a2�6��Il�N.�l�|��u!HY0��l&�@Bm�/�湼��zBq22�Hx�)�T���:��ACi�$:�$1UhM5��5���=ϮZq��2J7D-�2�0��L�i:�4�d�X)��湬���߮aza0�q���$�ʒɦ�`,&X�`�V�\�;���e�a��Ȟ�M�z;P-$�Chq��!��xÉ$�&��!��{Ԣ�n�u��]��*'�qAr��C����~5�<����Q1@�T���N�%Z��\���t����=HCL���@�2q�z3RЅ�C��Ğ0��Q$��;���J��{�(\��sS�~�'Y<d���i!�u!���RN�6��-��4s�xoּ�Od�^$!�Wh'Y򃬚d8��8�x�=0��d���=!�8�Xoͯ|ִ�=3��l��$�H"@<M�&<řN0�I�B��0�q������~���Y!l8�M�u��S��e���!�+�!�) m�u�޻��=S��s���oU aZ����ہ�L��O$� �$��&XKM2B�9��~��nHul���3A4��cuH�:�n���i$��D�b,�������)���$��Hd=0Z@��2���0�I2a �$;~����N��gJ`R�gP%0�`m&�q	���=3�C�Hv�rM;I�����d���q���i��4����b���gjC�CT�ИI(L�[?P�t�W�U���o�"М����rFNE����ּ�^�Zժ�R�qn���v�u�'��ܑ*���M Bx�4��L$<I���$�&R�R[ �TH�� xh��/��ᔁ�֙&S�'���	6n�4��m 0�`Um=!3�W��w=�Be!ҪHVj�OI�u����d�@�I&X&<a�=Y��k��<�|�-4�H�$;�'Hyu$+��;�|���|���8��(1��{��m�@v����K��[��Щˋ<,�0^��zm�ȩЍ�0��@��R5,�̙ǅ�C�u�a�^H���M��3u�<n�L^��P�����mV(�a�g�5��u�5����,*7F��#��{d]��V$n���YAHm����w#�M����ϟ{���r���Y���u�é _�f��z'�������!�v�v͒n�{k?�;�İ�4Ã%�U6�IG�8���t8ξt���r��Y��;l�Vog=�)nP�˞;���ו�6$�%�S�2�}[t���B�&B��3�zQ�ƻ�@k-��a���`�?;0s�t�eR�<�g�z�VX��kV�`V�VT���֧xkqt�涚Q��mIa��9���67����{|D֓jdLb7�G��F�r:5�c�����X�x�o�GԨ���[�ܨ�����zuP�����N�)��z��V�����Tz����C�owj��7�2�zo� ��$3f����ut�N ޻v*�%CAہ�(���Js�c�50���^�Mֽw<�	��R�w� �u�t�m���s~���%��ӽѹ+��q��I��ĦD��N��_���o�I���<��Ӊr�=����&����˂�~��|=+$P�Y�#��������Cj	m�f����6�1�#�&�f)M��8�껕3Nc��m�
ݣVcwu��:u����a���S���ze���+׹�"ڽW7�#J���YDv��4���̗�_�}�DUG�����~���h�Cot��ZW@�U�*fS�e��z�H9֭��r�N�ԥ������P�����ϛ��C>�_���>v����B�-��Fi���a�;�t�B:�xN�8K��L���SDИ�ӯ�4�2��yь��Ի�q�˭"��s��%��w�D֕�ue�g���yK��h1�on�=��B�wAb1�ܼ��;xS%ūj�n��}+���$�h�i73��9�G�*���7���u6qmE|����xӮ]�k��9��1�j�T��B��n�������j{K�e4�uE�����G
�N�ƽs�ܩ�Qq=�D�AR�um>�jQ��Km���tB��f�X|v ��v`�9`	�*�N7\����f
.����z��3�J+����J޼�A�V�O)@��׮_<r�w8��g!��t�-�=�u�U��73�v�f�+2y�]qE��N�"������n�zsnSj���ٳ �ӆI��J���zm�nS���\�� ��FT�٢q�v���5(�:Nʕ��I��֣�&��8ےH�R9tW��O�4eIc	�������;�|���U�4R"�UQUw^�G+�s���Ky�b��F��)��WUH�y�9�L�UJ�����u-j�UYh�Q�]�(�jꮂ��Q(�i�Zh�D�(i�˦�I"p�Wv��M�EV4���).�A�iDb�Pb��U��iEDj��H�h�R�ꛦ��J��KjE�����uh՗�ŔRP�7uMUݶ��..�HXPx����o��r~���i��o��m�Ԣ��P�'��M���~�������TsfS��[eov��Xb�ٚ�S��/�tv���1֭ۜ�j
g�M���ENl_T5�M�L���}�sqf��c��Z2�$x�"����<�s��ȸd�'wI��Oo��u~꼤I�ϒ�9����1�\��y#`���Ĳn&�]�O�b�	��Ȅn��GH<�
Q�o���a���&-�B�vQ��xq�F�9�̓�{Z�)�rPE>���#޾�	�ܽ��6�[��W@��<7��T��%-�J��X��\���e2��X���T�t��a����6�	0���i��M�u�7�3u��rL�_�ߋ٥�5���� 1.����R��1X��������Ήx�m����v��L�}�/��z5OS�+۶6���^�W+W\EK�NQ� Y|�GE���)��}wҽ(J1�7;ot���asggF��~��:�5~�s�V���Z��{|Q���5"۟߮���k��5��Y���]q�N�VQ��	� ����@M_H�v�go!�v@E�G�/���aT��~9�k�O*֥F�Ga���o������4�A�ڡ���n�������WA�י�u�c�Y}5��Y��l�����CmN�ץ.&���zO%�:��)r�����l�.�Us�Z�^�֔��u��Ux�ö�N�W��:���3�[53������f%��SmG?�_�uU�q��=�7��-�yyO���X"�n0�ww�rT�:냘�V3����v�]6����6��sJ�0�C�e�k_��/,V� ;5x�E	D��]����6zC#��Ӿ��b�L��-�y�!@��_�>rx�ΛڵǞ��ʔ��Md���a����Ky
��/ojJWٗh鋚���4^19��A����\�z�xdNk��Z�u!k�wZ��nC��~��g�"�m�p_�÷+��-�Ӓ�<��gjL�5�	���Ś;:����fׅj�򦨦=��@gU�c��8��';c4�����(��o��}OkE8�j8��}ه.��X4*�Ǡ�R�N=M�Foǅ^�
v��p���%.�_��g7�m~����8X���yȥ���k}�#�-̩m�U�r{�>7j�U@z�MY�Tz*;:)�%�i��r��T�osn��o:�9쇶A`޹�o�Y�]�;��.�E�]`@�5�yđ�[.A�������# Co����mm���2Um�!T��GG8B1�����obկT���O����f�;�.t\�K���L��e�B�o}{�Ű��9�,�&r���#��=���x���@�Z���9�vU����45�ۣ�*�K�j�ez����W��hV�w�W��c�O[��VT6&M�e�f�����#���D~���~���I���������]b^)����[�1�8.���8�w�׾/,�[W�I��Ԧ������P9�Z�3�֯�����ޘD}3�����x�f�f�
��;�އ��\i^�w�:��ղyť=M���;�����x��^�A�*b�h�I波=�@�}bq�����=�n�^Cp���uƌ�e��|G8kۤ��J]�����ˡ������Cj�0����W��_L�G�$R� �_�]Y��[��b�$F��9��dSTa>��
j
*�|1Vm]������b|�.����)gU���ԗ�����@_Pl�<& �F��{|���ܐ���{_���I�yi�8�{S$*����#y�:{�^��z�b�O�'%��H�X��������[�xd�#��-=7Z{`��i̩��e�k��:{��_5����� 5n����JV��)������$B�Ǜ�=y�n{��9�c{߆��^g�tB�|������۷L�=��O��ON�M�&};9��Vu�������j���0/�V�?�~�7����}�e�2�K:)�7�2�,��J/d�s���5�������%�V���ƃ���9�><<]X��oZԘy������Wo�ʋ0��³\���-6[����ۯ�ђgOf{-���5cĬ�y�n�u�>si{_7���'��Y}	%��ߌ��r��!�;��X�*�y<>��j�z�Dv�Ԕ�C��y�m9�׉
�Ϝ{��'a�� �{����wm��.�Zg�lN�s�,甭��H�T����z�P���r�qvL�s���V�/���0^��"L-�U�ӗ���Ň����@�Ѥ
�ޑhY�
-! ��Љ�3��UGNn詏Ϊ�"�4H���u�(SW�k3�g�&h��o��]S���;ܵ�g=�IБf"M^�̲�`޷��*�k��&)�m�����HQ�����n���ǻ,���.dޥ8�(�4v�|Z��H�J �R������P�ⱳ,�mR,ޗ��$��*���&ty��h���zq>2�w5+G2u��X<�k��4���H��-�a�-5���ەwB���I>���΁�\��n0�9��\ǆ�D�u"����y�M*ͩ��s��C��+N%������Y�Q5��_u*fˮ��-��lݪ�Z��4��of��	m��2��I�KuَĻ�F���+
�}Z/�	cFq�p������[}�\�@�xp��6��9ǘ�.\�󊱝޷j�K��WkTr����'.�A���gt%Y�Q�<��܌$-��dM���R������86���+ɻ3RiA��� ��X��c٩���Q͕�Su�zڛ7bѝ�8�ZjLƁ&T��	�D7K�H��D�rI#�u m�7DD4�e�n����fw�=��wrզ�DX+�e��"C{6�5wL�e�D2�% � ��sWs��Yh�n��X��44RR���cU<���j�R������e�UCE5T�b�҅�P�-�ꩤ���B�*6��Q�Җ�PZ�KV��e �]�Ж�)�]�ˢ��RUSL�"ʪJ��H���h�J�Z�D��7h���m(Ř��Ԑ'�M~y��c���vV�ޔ�:�[�ޫY�wG
�3�o|�����O�)+IM��f����i#��Աz��x��+�U�i�G����*v̙[��re<@���GF�uY�_��L+��^~��]����ݩ��Ja����7׷���}oq�ue��uc��?�v�J��p���ț�d��\(΢:U�������n:�mp��%/uA0\ǯȞ8Ю5Kj�B<�{��P�h�_�wzC� ìsn��C���̒��x�+�����L�Dr�m,�w�z��q������w4���(m%���ގ�msЋ�p�5�c���8�Io�z�d�T�o��'/���u�c�k`��^�<�"����u���·fnZͬ��+\�Sٛ°0�_tK���5x�~k>���P��O��0�o{V���yU�K�M�ٯi���P� �#ٌ����d	+�g˭��R��2q�X4���P+Z�w�1f�H�I��c�xߜ����g��=�=��! ��o��x�����X�ؽ�f3��KP�3\��]ֻP��(����6�`�b4�Q�T!�����2��@(�;ޫ"H�So�젵B��j�V�פRwH�tyֹ�l��{$!6�Lw��N��L����-�)�$mξ큿�q�|+'���A�fZ�ӄ�cQ�I��ñ�^�f��nz
�yЗP���
���dQ�˓��q�������s���o|�=�{HE@�9�/fo�W^�
��\o���-�mJ���zV���v���4���"s�'�%����^4�	�P��4�2協z�=���<�׽A�5�����wN�x�����^>9�ky��GTw;|(LU�v��Žgo�LL�a���~~t��Vouy[�h�/D��O}�7d�DBͣ���SV�ӫX�Î8����+.Y<Kn�a+;�69ַ���=�"�M��ww�^c]���#�103��B'8�B%n9�s][=�߽�eq��LFC�F�y{^�E���� �ɒ��cx��Bj��j��د�M�GeGm� ���������.9�Ò�:�N���nޝI^�B�4�Z�&�87����)�56/]|8j�1��|3��~Gq�:�D�)a���?2�z��#v�g%t�p�s5���x5e�|�(�ܡ̖��A=� �I �9�s�{/ʼ�����x߬�7���Z���d�LV�7�%u�8&�
*�î��zҫ�=���l���yH�r��:��0���Ϧ|ėV�:�Y[ĎӬ�ԛ.���/�����ɮmTm�9S�4����s�eX��ʹb� �e���Y;}q����AAP��z����Q5��s�+�9��<�&����o&�������n$��H��riw��fL�9����Z���{H
��7���ӏ`���8��ב���nk�bŞ��~�;^�>[��h��5��U*N�2���ا����m�S̔pU[�CVy�V3-8Q-�h��I�y�������ȋ���4���F���W4����q굗���W���i'֋��l8�!č����w|�L��S��׳/�&�'|�hʻ�}[_+�)t�5�-)-6��ӭ��I�<S�)η�k|�@�����߷���h�xz��d�
�E��{����b�ݷW�xZс����bQ��=���v��q���޴}sLR(�
�y���w÷T�`�;ʰ�6"�u��̮B��ѩ�[���Q̵~g���x�E�,��EЄ���p����R���4j�ؾ����4Q�um|�	�7I�_�|}�3W���B͑�?C��v�z�܎����*/`8˗r%�ҡ�șV�W-�t��WE*�͹���(�6��kz�=�{`
@!�o���&����m�4�:w��	�!�����(/z�~�3��˘��t%��`�C��1�v@�N����j�m�p�9�8���5���o"v�zm��O/t��z��������<���{[?"���k�	6f���M�o[񭿹��׮["��)P�u���Ư}Ƶ��ުQ��Éᢶ�*Kx{ǧQ�~ߡ��:}\�8A��� I���,a�����Naڸ�s?>�s�x�C���Xɮ���C�?n!N>�U{6ẅi�(S�����;چ���E��V�;x�קg&gM˖�朘�~yy��y���u��{�'� �	s��y���\��L4���)���m��n�s�yӰKH�8��)A ^���L�Sp��y����	��T�iEn�����0��*#�#f�CO�G�A��۳y��!\�6�6�B4|E�[��R�v��~�:|t���H���.D�LŉR2Ͻ�Z;�\�Q3��|D9C�&�餂�$E�yc��Z���뭿���'�J��{��i�DK�q�v�:Mj�D��tc�Ϟw:2��N���u�e�*:��o��&�8f�t�_}��r]K�.F2����T%Y�"�]ރGX�M�Iw=�_A{�m�$��zsꇎ�wKȅ��Z[Tv��tr�G���f�<^�]6�*�+^�(J�/V�#!��tET8��}��r�g8���et��AɽsI�ٗF���n|Z�V��u)�����\����29:�T\n��9�۪�XŵM9����á�\YI7Y秺�Eo3��K"��F[y+a��b�����W[�z�_��x����
Py��5�Y�yg��׌;;Mt֩�̎y2�D�n��4m�	4�6���w��-x��wWZbj+�Mz��ۘ�vet�6��w����[M(��G���0�y���V��6��;����2��]x���J�����Y*�O:���
��
�C�&�彬R�I�yO��K��U;��r節{�K���n\)u��[�:�K1��&�%� ���{1W��8^Ǧ��tUN�b�=��ќ%v)����l5�!�j��Û�n��]�2��L�R	�����H[�D�rI��u4Ȑ�%܉��-7߈껮���U�4)i�xJ���i�T"�F|�	MK��qMSuK�T��<�|�!G�Ln�F+��1n���V�1Wmإ,QqUTT\%6U"��T+X��8GX���F�b�ZQT�Um,K��o1n�J�T�T�*�M�M���E���SJ����
Kpմ��a(���\qJ�	Wv�T�.]^1wKH4#wx�ī���bܦ]�[WU�(����k6�
�x,�ֱE�IEb�4Xa|�5�]��p�/=���.��MY��:�Γ���*P�Kn����]}�Bw��{�P��b�i�n��8��f����M�Q�����<D![�u���W���V���9����|"_�F5�	ʣ��o���t��x=v�2��Y�b��||f*2���2^�����ޮ�Η��#u�ȬN��A��Ǐ�Oi���~������W����,�8�����G��~'׹t��QÅ�=.����Z@�1�+:�������"��0�XI��!�D��7<�qR��4aDe~<���/�jʯ�_�<T�e�F\ڂ��[�B^0�wݭ�	�N��\Ŧp��uKjM���_Uzd�������8��)��2�*ʺ���֛i7g���>PW!YzL�b������͓4g�^	�!��C1�ۤ�3��*m4�;����̛:�P�&*6c�S��z��jT��V�c}_�iǎ�a�� ů�g��
�۫����}Ş"��qD#� q.{���e���y�f^=z����Pf�4��8=Www���f��W,\r�:\�X���.`=�{����/i�HV�?O �OO�`�
���bU&E�妒~˦<_�m˭��{���/V"�Ꭼ�6+i<��g73Lr�X�CK��@OE����u�gK���i��YM���U}�}�[�9���i����N�h�e���+��n�S��cH� �~����-�k���k�e^j��ج����h��IwU���G[�Z�Dw?8D�*"ȅ���������:Е�i��S��+oSi�I�&1��<u�G�ݕIC�X���+�߯�]&8�C��\�F��I����#����=�������t�h��o7F�_J��-0�*��<���S-�����
����$ٿ/��j7;9�i���ԾVݦ��+u<N���G���ڌN�.��e��I9��xo�PV9si���˷�_�*m�4_tn�M��gZ�=�l���&��s^��x��~�}�É��i��aZ�w��҆���sf޷�3T>r�i�Nt��3�r�"D���/�!��ݬ9�:Z�o�z�*q<v"�4���u�u�(�mۜ���Y��w;��hE0�%�b뉼�v�t�7OW1�5�d:l�D(R�����XVptGAב���a_�R�u��D���.�����j�,��?qg�g��7�c�����i��n��#��J��s1x�y�!Q���r\��T�r���|ǘ9Ǚ��͝ق��r�[�����c-c{)���I��9�
������<N����s�������� �w��֫�e��T,ו8�>:�]e�w��~�e����F(_�����u.��_܁�)IG�t��J���b���6F%�!� l���K}��#���z��h�x�t��Xl�����Z���bEEg�q�!؎��WOJC6F�?B+�P��"s�Nx}��6�i�ǫ�0M}?T])�9jV�.�)�q1C��?/���E����ſ{0U/�ְ�����"_/��|lM�{;���"�Q��ўC���4'�n��c�qW�k�ҧY�M�԰PP�2�i�uJ�arw`'���_Os�O5G
�y��|��Xs��;���xI�!�,��j�V��tcG�h�;��Ji�ӛ�6��۴1˼i0�9�,��Ho[և�w�,t�Yy�jz�^��f��T���P����B�x#O���d�ś>�a��{h"�?
#�=�0�أ�>����++G��ܵm�r���Z3]�Y�2�Dˤ�є�+I�x�/����1�ڂ4I���:GyqgKO����b� �
,?x���v�T9s�V����5P�}�rf���|��Є?&~Y7�x����}�:<r���+��Λ���̱D������۔�zy�f�R��M�J��)�7�D���@���s��J�4{�q��bpM!��+�_q�ּM3����3b�P�8M�������{������!��0�S������[���y}G-!�_e!�����J�{�yQ���e7�S^9�q���i�~�����"�Т���l;\Gg���{����ւ��4�4a�҅���E�z�iw����b�i���?��j�,�I���uY_sC
"��<Y�8��O�"g�[��shq�CO�I��+"�����M{�s����J�{������zw*٧�V�`�:��Z"�����A�!sqp����U�h�u���������"�I���v_+ؚJ�e�Vc����>�����}V���U�.X����t�;����}���e��y��rQ��Qb�$~hY��p�fm/z�i�ټ�	,נ�\����;�5t�����#q���e��%R�V٥G3�h��s]S�\�%�v�(w��YL�*V�uqd	���_$Bk��*���z��U�o�4�g��������^U��A��E�(��?S�����Q���H�_x�-?5K�g�Cղ^n��,�Ͷ%��&���Y�{R����%\z�͘NeAe�Gz&*Pس���{a��;޸ty����`�����@F�`o����'��?��y]�ŏŅ����wJ,.<�^�F��l�Ă0��j�W����w��)��˦G�u�,�3.��m�7����Y��9E��N;|u}����o{��p�A�����b�#�B/��
�ď��o*^h��N���_���]+�i/�uW��8�8n�֮u�;GOg��:j�����D���dB$�����w�7��U[Z�n�aL9�_)3��N�K���e����(z����R���2*������׻f�g��jV��O��SukZѤ7�%����o�|,!����(�j�N_l���5ZV?����\D��*vq�wP�\l����G�|�$Q�6-�gf]�?!J��~�y����u|+W�~��C��xC���W0G޸�ިR�u}�<{�󂕦��L�w[X(�!.��7Z��lm���U��������ϋ$��i~#�kչ�ϱ�k�C U 0�}z�8I�9����o�I�{�8��E,|�NW&�ۯ1z����z!�Vm�$�!���ܘf��e�cTy�نw�/9u���7��޾��x�=\h>�(z���y�]-]���}a�5u�9r�)��c�ג��d���۵WȽQ��rg=�Y�R�|FI(bJ���g�Vv�`<�n�^�5<�nԝ.8�+B :�JKXp��+p���UegVer�{!���E���3�eM/�u𭺛�oLX5��/tZ����n�R=�P���S��엇N�[�#��"�Q{i!K+q}t��͜��L��r�tV���=f�.�K�[/1���*�2����Qf>�u�m�Y͔�6���"r!o&̣Lm�	���H�}��s.�)|��H��[S�}��[���z�j?�{l�	W�*��"�dnԬZ�e��f��f^j��D[q���u�.�DC�F�n�[���J�4�9�D��Wi�;u`Υ�+�<�*s�8Ӻ��pڕ�¦z�,R�������KjI��^9�Y�6d�0n��/��H#�h�"�H֋�'yftr>������y�y�R���t�8�֎�0�Q�B��tfY��}��y��RӔ�o�2��r	��(��rIrH�H�>�9sE�\�2�C>�Ϝ�5��~'=kgj�lT)��bP�mSD4M��tR�E��r�)PB�c-��Jᦃ`�\U�U
�g�������U��GB���W�H2i�A�h_&Yc�U �,qWiU�QTeխR�*�j��H�T]$�M�*�/�hQd3��Z)��5mU]�t"]a�-�Ueʦ쫶���Qj45m�Ke"V)�[���*��	H]V.����T��wE��R���()Ta��4)�T����65AE�%n��`�KE�qe-��U�R�ݴU�����ED,��L4�T�*��TR�j�c��V����n�L��i�Vxf�ߜ4�5��[����s��o�Kg~)P&��yq^��&c}N�S0L9�SF��H�����C7vQ.�ng��ڙd{�#���t�_� �y�1��VܣgN$<~�0�-|�hB���kY�c>t���⾹F:x�,�3�Mby�pC����Q�P�	�B���>�Ľ����_?;5i�!�@~���zEX�n�4@Ә��Vi!Cɑ�<C7�f#��#Z(�G�c	�:��8�|Mr�����h�tN��7��=hnW��+*�S��z���n��2��R�F,�7���#:#j�۵��w3���� ��*�����Q���W��$�9�sׯ^&ݯ�\�ta�`�L>2�$��k���տ��~J�^"�߮�W�c:�Bˊ>�*���]Fb��]7K�C���6�9�=/P�5}G�Ⱦ�@]Z,�uV��){�g<���x|f쉁3?R���	���_��I��Np�~�c����D�mq��sg©"3�_�6~EZ�}X�á�ӿeCdth�`����n�ӿ�*��Nb����8k���;����F{�9뺨���77�2׋�`��=A�u^:�ze�e�&`��;�0�c�ú��䉍��)�2L��%�CJw���k|�9�'���/|�{ܖ�>��O�n����zf]eh�����K�}�t�W�W-0Q���,�G�0�x�˞)����ў�̽\�NQL!I}�<޳�g���\C��{�98h�D4F{�H?z���� W���"�Y����q�UMT"�n�#W�"���I�����!�FT�4&(K��|5{ ��aNJ��Ul��h�T{�z��maF,�Z�$yvz]W^]?")��V� �_q��b�^z:l�s��Z�~$~C ���U����FU�V�}J����͗�H�f��ۇx9E�/���PsrG��ξ���%�qA��?�>�$�H�9�v���Tz�6i�m5��O�çl�i6v�\�����"u��N�I�T�jh�x��/Z׏6Tڴ1L5�+����9n�|2���T��NN�
�I��j;��Na���p̙�0�ʘg52��0�!�/(��_�t�6�ᨇ�]r�5���qM2w���o��<�\��:/,����'�����U��a���t��DX��N��V�G�ӗ���%��/�l���h��=z�r�4t�����7�.��0����i���x�C��y�H�^�T"sA/F�l�Z�]u7����՜ej�I�%O7�q���rJD��J�_�?L}3G�6�ƅ�蟩ǏȆ��/��P��S̙(���d{�����e������u�����0�.=Q��ՈQD$�+|Q�}��d3�y��|��:_/k�,:�4����]m���vP����@��7w��α��9����T��@�e/���[U�^�`��
0��c���8���
l�f��$f*0�͇��,��Z�H�.���}�в��Fȟ>b8|z��FV!��J��u�Q����@o����u�9��~�������Ɣ]HǮў��4(>�����뾸)���[���oZ]��T���{�|e_&���������9�o�4���ǭܻ��4�[�1�7�~]e�V�t��4F�<��+�ӔvP�_��\���DaDaz�0��O.k���ֳ��ۤ�-�&_an�q���v�pv���3u�U�&-���a�k�u��̔~��f[�y���X��=����̳��x�ы1��8Gqi8�Nnv{F���!���#�8�<1Eo�o=�3z���"�4�Vq>og���L��]�����駨�_B?-q$m�K%�yZr��^��lE�C� f�d���/�Q��H:4��[*\	VL�i�Ғ�*6��YB�7����*kTy�wl2��Jǫ/[�=َ�����(:�7�S#�\�m�m�_cW��;,�8�r�8k�;�Cԭ�����n��l�JB�Ç��:��	�*<�}۷V6t�A����7��9�=I����~�_]!9/W�E� ����y���+a�0�!�#���z��a�5�M�ƻ��~Y��I}�Ƣ��?P"k�K̿gϨ��o�i��Z�/�<�hjM:�I�Od���_m$Q-}�#<�!��, ˤ5ѿ���k�e��!��� >��z_�0�Q�"�M�.Z=�0�=h�ξ���}�g菒I�pf2~�=���{r�̻-��4��J�9�]��������0�d_�3p��칬:E@+X7Jդ*����_���ǖ���R�2�*��.D�T.7��0��L���V�_,�x��ѡ,;]f��X�=�_<ט�q���*��K�_*j��}��/3�L�DQ�_D��Ċ+�CH�%���޹�Z�\�Q�폍��#�Z��!䇻������xD8��!�_+����)�SPa��7��p+۩*d�sj=*&�{���%NOJ;��<xMG[z���#+k���kqo���bĬ���;���Bc�N;�~�13M�e��֨�+nu꧚��*m)q�9��&O��5iU�#�o�d^Pn�zf�<�$q��MyD5k�U{��ݬ����e0�3���8`8|ƽ4x��-wY����+c���_xч��ެ�+=�.>$��! �p��u����0r���K�(_ݫ*���]2�|�^?K���c܃?V N�t\��g���dY��a�.S�>#�l��X������פ�qѺ)��R`JB��dO��~�V��ݰ�'6<	�����Y�^9,�/0���͉�[�Mr�{����#��?DGؗ6߮ruA�_�������.�ݬ̡�|�盭��!E���$/��Yҁ-@�mJf�k��F
#H�r��|p������;����x��L���fŬr�:\��q~w��q���;<Ve�h����> ����ܗ�to�zm!�Ս�GWVrzЦ�G"�A������0��D��ڙ���.!�P��0�� ������^r
�MB4�;L~��C�~��/���MO�ތ�EX��|)�/n����(VX�Rx���:�����6#7P.����=�N��Ēo(�v��]�j�m��ۭM��Ko�Sz��Hn�-�}�5h,4��s:�3��2����9]4��Q^-�زU��!�B�p9W��ΡX ���a��f;$�5Ȯ��X���x.��b#R(��x��"Gh+�A��_̦�Ef���M�4�r�ɜ{q�x���V��t6���:���u�b\���ѣ���T�*wW1��U����-���9>�D)/qR�b�kj�f�q��g10��W\Uڲ6�r-G�c���pCM�R�Ձ@h��q��i]3�OI>�Ͷ�7#�<5��x����G��T�M�+��4������W��]"��:�W^[�F���e�K�(��%�ۦ�ik�w�9�/�l�A֙�փ���?��YE�;+�mo��@�e_��3YW�|z���ljU��.]�	7Xqn�s�����l���^_*������.�XM-�k����O��gv�-�j�=1v��Ge:/�'��ʸ�n����4�$�I"S�qĵ�$��*���Y�4h��} ;�i��8�T���R�e(���RU1��}��q5l&�*-A+�UA
�����>g5T�P4њ��i���R��S(�V�����*��70�T[(�Ye��0X)2m�T�5B�m�d�j��e�����U�\1���AL�*m�X�-� 4�A_�D��)�1b�q���7T��iV��K�-��wn*�q�^1Cq����R�0X�.�J�]mW��&�"˶�Uw�`�-˺�ڻywAp�=�#Rs:�2u�a�ݗat��{��������i�����	~�qm
�b~�.����V�yn{�v�9:g�S����GTu�yy<�����ӧ,�oU:j�5YlL�U:�3�9�u�$��Y{��Oa���"4��=z"Q�H��An1u͑q�J�O5[3��q���L+���]���<G8FR�#r�}>�FR�K��e�_1)�S��+��:6؜�S
��?q�3����F�?lsq�)��
�?3�ӓ1s��r=���3��t*~1����@�g��l^]�L�I��JoNI�/��E!���Fd���ӕ�[I�9;�\�yƗtv��
)~�3?}˒�\�?�|g�Q��l�LQş�|\^���� b���=5�=v��9NgZ֜�8��&޴yB��lr�e	�W�T���\�����?\�ʩ�(~F?�39Aã'��n�m�����@���v�B�Y�^���N�t�ٺ|)�_���u�/��%j�%r���]ְ��>Cו��E Ey�D����G�#gI#����[��򠻫\�i3g|�C���y�4z}&]�j����y��OS)��NZ�YM�똡|���NG�{o�3�a�jd����
L�7d�)�\u��헽Ñ��F��� '���D~��g��M�wJ|G�����J?
+�B��D(�٧��Pf������"G8~�f;��m��X�xo���ש�i��gU2�gv�z�h/��<��Zl����G#6�éٷ��k�1E�,.�y}x����9~����R
G�B*���5�-ɼ_{�oZ�l��J��ĵ{�)����d�r���9R~��Q�ő�XmZ��^e#g�э?6��j��"�NaX�R����i'��k��P�� �
8S��}��e�˕��R�8+fX|k����O�*�����ס�̓�A=�%k�h%t,T������o��8zOo�U��Q��e��Yl�����)w}����T6ۖc���z�ڄ�C��T3�==�v�����Ņ�)3N�7G����מy��SL��T�e�tr�@�o5�v��g������;||Q�o&FGN:��7n�H��C㪘��H�}Y�R��7�C�e�7<�<��J�4���Ϭ?.���p��*����|�SQ'H{�^S��]�A�������^x2��ےa�$t&n��8�4��=�����.�`�;HBw1W+���r���g���ۤߞ��kP����\���s(ucٸ���P�+��Z�'Hӊ)u���Gd�˼x������H6��&�Q�&�}��4�7�=���K��rG7��v��R�.�6�����8{7<ǹkqx���ئԾ�[o���V�����1�YO6mB�Fv&!�}�t��o�����0pZ�ܫ��b��[���mn���T�2'5�]ڋ�HZEt�t�=ȥ�#����D}�y�����!.��_p��~Y2���P�^�iU�YĎK�t�i��X';��M�}���Y���s�4�7i��#r��<�64{�>�jF��s��yc����>n�z٭r�*��Wq�n���R�}�ZW
'6ۨ���{�ٚV�;��4�Nz��}}�I���o	����Wٌ��v��x��v��mf��� hַ3��2��z6*Vle9?����������6__��S�o�O�kF3n����L�?\R7��S����V���޹�
ȻB��G��=�u�*��RfBV�jx6,j$G���q��.�J]�1J���kȖSc�U�8Ϭ�� ���xL�#����P�*:��]T��5��9���u�Ω������[���=4�����
���=�e�K햬���ǂ�=�"�&�r�R�S6l]�*�vr	�,�Q,���1f�h��s��������#�iO�9[���끔�5M���Qٶ&rڶ���h��똷=��h�z���Gvb���O��v:��Ɋ�#�)���k��}�p�*7����皨щ�Ux��R�Ř��t��v�}D��g�/	��k��z�i�&�$̉ꗗv��'y�o���� bK��S�+�4*^m����x�+��mγi+���wF�הIp� r�W)����D,�N�D�ǽ�W(q��=�=�E$������_y}cm�~�}֎�P�lRI�z$�ܳ���ұ���Tv���3Ovbw ��g7�G�ڸK-�f�@�x;��!n��T:kq�B�V7vE�Fϰ�o}�m�-wI��q��P�!�,U�e��6#��������+�;�gk-��U�=�I��7:vZ��謶<.��2�˩����Q&��v��μ�EI�٬�� 4%Z�m(&����/��鈙��K���?�۱�R]��o��?6"��^E�%c�n����}\]W�o������;�5���ё��$Wj�g��cե��'v:�-�B1f�k����E�aVo�em���l���=a���z��OUE�4~Wy�u�0^�
�����ꏩ�
o;����n�3�W]�O�tIͣ�2�8r�3#<�vn�k4�T�	��&�o���Ȫn���tړ򧩷��5�˫�
����F�P!�����G,��v�����Qۧ��)�X���GWW>6�[Q��1����cz��쭂��y��j���mmԃN�B���^ͭ�*UN�E)�k/����H��\5�Ο�dnVv��S-�����������u�t<;���=��)G+�WZQ\^+͋��|�p���$�[Ln���g_W#�i�������]��)p�����	�˨ù��3bѵ�e�������u�/V��Q2�/1Ŗn�ӏj(ź��u:��Z�@��V엧Uv��+�R�������q���ڙAf�Ҭ�}�j�@R`N.6�>�U���q	�H��y>��qU�]����_��z�u��.���W�SB.mؚm����,���ÿr�Ä�S+;��H���WZ��L9'k��k�ֳ{�����Gm���w&Q�d,�bW[�Z]0�� H�nsg�K��P�f�NRNy�#�I��STR9V����,�V����`;�G�<S4�b�&�I��T�'�D��a$�UK�7�($m"�`0�Ոga���VUcϙ�i���v�4f�.�vն�WutU�]������T�Tj�2��&�2?&�n�Ì8n���)F�,h-��*�G	M�0�EQr�*�KE�����R�ե[q��s�ọ��v*�+*R�B�]�P�wuCcUv���,�J��*�AE���KM4�$�#T�A�UQg�UW̲���*��i�����B�ɊtJ�UI����	�ˠ�#Ha��m4E�����eWt���|O]�����/�t�I/�zfc�o�?|gG�}�,qJG��׼�QWw~��0=��|{Y�ە���ǠOk)@��6 �0lL	��t^]�3��[P9��0h�1}�݈�� eא�L�V�XDp��ڑQ�W1��.]��X�]M,�U�����S�����c�L.7�Xټ焓}�!��F8v �㼅�����ա��B�ެ��n�`�\�c��&[�y�έ&S�/[amܡ��ܿ�$�~6���o�ӽ2��Q�'�أm�6c��)[��CKވ�Xz ˸���yS�=��������=�X��baؙam��ߕ�/:F��qw�/7����N:
�Y��y�f9ȕv�����cc�q���g�4��sֻmm��A��=��:�6kv���Թ����xg{���הO���2p��H�i��3���V(R��ra��F�,S��R�e$�l������S�Q����Iw�V҅lrlJUbڙ��S)����{�xP}Y��q�i�����l�u
�3w��vf�"�0_�-�c:;5}��m���k��[Cޚ�Oŧ׶5�__uFL(#,��3/K�������X����V�
�\��	tݣpQ��¡�Y��u���Pes�J��NC��M&�h�Z���ʾL�&�^��ր�2*E�%�&{�1{��O�_H�zo��L��
�M�V3Ҍ�٫���'(������|N��Fh>�=ML`����M��^����fh/���Z�gj9�E��3�a,B�ug:j�Z�p�'��\X�Q�L��汻ޱ���Y����^�l�ؓ��3&i�cr�	�;y'R�HT��P*������I	,��bK��T��K����%ls��ڝ!3uzn��L�@��v{9P,uv�躈�y�[���<����TS��9/"�k<�+~���V7��Bh��;%P{mg�۹o��vO���G�vT�ұ�w��A>�������%�79��-cܶ7e�P�TgQ�c")��n�JちS/	�u;�ѷ�ܺ��':��b�F��m�D�H}��,�%�x�����c�Rq�Rm���U�+ve�G����f3��%f`��1�؉ҵ�p���` o��%JS��zoJ��ޮ���{����!�!�҂qw��u�^վ���q֭wv����ٰ�k�$[<S��2����ywE����<4�o�w���U{��q�HLoW��7Y!�s�y�����G�bޝ�t�.�,(7t���=�%�Vr5d����>ƌV�P�Kn$RO�����5z�t0fs%��
�G�>���z�@���j�݋cy�ؑ�?o����\��\b�Pb�Z�l����(]*G��0L��x^�M�:�PIr���:�)p�p�V����G���M�P�z��Z�A'�>74��>ܪӵ�Z�ݛ��!�U�|��鑷����k~U,Y	ۆx�S�����Wհ\�g"�w�G�9@�oD���g)��������/֓IGl���$���`��oA��עz"��X���~�p��;�^�a9��>�T(�-K�.FD�~9O�}��k������e	��oE����Z�wv;��3{��_�w�����\�~�[�#Q-�j�������MY�*7j��pA�&t�I�"�U�ɭ�}o��y��{�~,ٳ:/����˺�n���B�"�&bi�{ o�p���]Eaד[��q&W��e���IteYMD�H���޴`e���lr�-�ĺ`fŹ��[�g��]F�I�֒j�wg��}���c�L`y&s���S8s��M��bc8�U�� ��jݲ:�Z�����[s�Ϗ��ѕ�Y����Vˬ��ʑ}z�m�ܽH�G5��:���0+t�y7٣5�0:w''�r��}>Bo����͙&���/T��ߔ1�ϸ�C�I��o>�m��Zc��_
Q$�C�<hgѬ��u��Zw^����/b�]����;�t�0��n��UiT'!�k[�}��.�բ�9x�N�̢{*���8�.-��:����i�A�S��3� ��n9��3�%�ֳ,<�rq�m�h�w�;ec1�)UEV�����9'�S�`�OAV��u{�]AS�0;��wx���Ɍgٖx`
�1�{��s@��QY�~�z�����j�3y�oA�D]�v���@��Z�����Xp+Y`�m���+bN��Ծ��p��ӫi�]*�9]-�Y���9�C�u�L�p��;f]1Q��7�p�7`���V����p,(a�1�PJ�y�]r�yU������U�,f�\Ƚ���7���cf��u��\�ܕҩ���e�hp5�9y��R�ϻ�B7�z���}{��38\}\���!�c�n��9���P�;5k�n��l�[U��U$�f��Z����3L٩R�.T*[�w倷�;&=�1��E��pZ1�Čl@�l'�f*d �3�D�ܭ�};y�mI[Ҳzؤ��ҷ���J<{T����j�]�'Y�����1�wR$��^N�U�=�5E�e>�!��h��Z��"����#���s�����;4����J!��d�ص�y�r�c�[\lL٢�R���ޚ��9R����Q���Xb��q�`���L����䑙$��m�؜��Ao'�mΊ�d7��ZW��L��v��4KD��l4B%�Kd&�u_�,��#o殂eQ?Pl�(�j���)��)��Yj���3*yn[Q�)�U�RZX�E�Um�Wul���%�T*�Īn�e7R���tUb�i[���c�Z�1UUM�wwiV�+T�t�YE�]%�km�t����2�W�\�­�uM�Kl��Kh�.�m��%U5SB���ꨤ�l�VUU"��UB�]�ICE�8q�]+iJ*SiWB�V�VԩF(�eV��"5UTҔ�P%�wwq���]�XB�
	�����d?������9|��6�7�ɂZk��w=�9|��\Rq�i6�����Fq��L�8��v�8j�9���.V`�αj4���tc�����7�Հ��m��X��+�R��f�����E/��G��u�����"v5a1��Р����	��������zt���7��6�t�%i6sB�i�R(�9����|h��A��'$$n����kq����v�֕���+V,���d�-�6����uN�wQ)Z��u�Y���VsjI�JR�ք������=�h]����Z�-�`G��&iD���t"\�)��Yt3U[�g#�^9v{���Cw3�%[[MVƫz�Gtd#tXi�:^XF	� 3�l�,욻��G�f^X��\��VK��O<@�L/_N�&Y�:�.��类����ϕ0�8�|VX72h?,����ݬ�ʛ�^���/kJV��r�(']����JS��'B���=7*+`iM���ڍ��E�qf�͹׮����#R�+�eW�iLgx�����W�'^Lj�o&+Yg�ʉ����^��(����tʔ;�o��t�AQtȫI��/O�ѬƖoPU�:��'�xa�U�'8�'s�Ow����"��0�S/�S�����T����(����x�#*��+Pu��[���<�u��9���T�9��'O��b����Ao�`G=^[&�VE���[e�o0���Ք�N�k��0�0�y��1�m�a_�^!�9#Ԙ�Ar�����)mS�N+��ek�z��;nv
�ano�偍|�E�e�Rǳ��'Z��\�6�0%}U�Њ=zΑ�9i�N1.��C�!Q��\���(lP�T�>�-�V�����ſ�
�Ϣ��ژb�y��ڤ���17��S�B�m��q�w��u��;��&�T������*^���wln�/��:�k�;w+:B���Fw�W��\�!dk5y���0�Lq��kd���uT�j�gz��ν��p[�����4�Gq�UX���(�0MF3:��s������O;>=�Ǐ�#�>��*��8��w�63»���6ly{�L�V��BtA��S�ޥ�����hF�����,J���}qVb�Xq{�t��q~a�5B"�f�5�c�b��3-�&�/jle fs���҄��-��y���3-Gi��^��̻Ъ��l,�=�4=����^��o`YP���+-�kbx�D��;M��GfHO.ɘ"�27�(�'�t�e�\�����,��]�%Tq��6Ȫ�����zk#dD��S��8�d��î��5����=w�-Å�x��翽�a���f~�θ��]D�Z g̈�U/hug}�וJ�id׺b��'v=�g�̺y��u��4�ӉrG�wE�ŘR�xj�qV_�Rp�Dn?m�-��&o.J����9��`Hx���J�$>ņ�lk�j0��x��{��<B8{�]X�w]z�{i��}�c�ɺOP0����NN�Y�Hݭ�����nf�.:8;/�������9~���s����� / )��-@�O:��p��x9��1��+o���G��}ٜ5`���P̜k�Q�ʴ�A*(��\����8s��	}����u���-(�짶`�2���x4��d�Z��.��MPY�M�8�����\wp'�:�ⶺ���b������'�S!͂G�f��:�r� x�q�ո���\^��w�����_U���l�5{=.BL�OZ0v*��!�,h�#���Z��s���T`��ѕ��},a�v�[�[�@�(<��L�wX��nI%+��ӱ��d�.����n�;� _y�1�f�^�.�1��׽3��ٶ��_F$�4���ZK���p�w����*��b_[�=Q2;y�����S�w��zd�쉊z�rei�;ΣD�B��q��3ŮQ]fo���~�f�[��|�)vg��r,��Iƃ��=�5�WGq�%<#����=�H+H�1ݖ��X�����,�U�{ɧ�#*Q�m11R��Z�����OW��y<�T8�;,x����!�W�X��U�7�<T�݃����olUo��ݜ���A�Z��3��y[�_u��|��0^-�Q���m��[+�4&1W<E�g����]n�յ��O�:h �f���yF����w�+x]�X�f�#!`��=�f�ƹ����[b�H����莰�JZ^#�C���Z6{V>l�-�v����ռ�q��XMu�&QU��V��Z\d����N]�����!��V�J���,���}d�]��	V�
��Rˆ"���E�j�puX�U5,!T6�,�w%�}�1�M�v#�A��-Z4��,"��0��ͦb����V�k�d���*"�Jo�����Dp��� k���Z�F��''���Y�0gmJ繳��4����{]�v� �'��r���oz
Պ͜53�2�KX5�/o3�w7�:�%`�0���̕B�;����沝u8%��Qu��R}sf"���d!ʔ�mlʸ�l�<��&�h�s"u����L6؀�s�{X(N�4���j��7	�TU���Z�@��CGe��%�P����˧N�i9��+�g-�緐� @�m��{Wӝ�G�ɕ��s�Q�}�@*��Q���5�V@�ꛑ�g *&�jyg�,��
���^�ў����I��#rv�2I�H����=��J��\9޼`�G3oٯB��m��������B�0�uS^eby�����C�*b��j��U7W������G5B��n�wt6�m�N*�R�)K���j�,E%��+�1n��H⬼U�PXb�Y1�D�l��4�,DF�m����j��R�j��U*���PУTV�]�T�
Z��v�P�����We,L4�źh�"*���*��,i�G	m���8l�4@D�=^��l�B�&.糷.d�3v�J��kYj8�M ���Ʀ�ﯹ��Y�ש��Z�IQ�w#~�֤���/��c"\�in��8⋱WG�Ŕ���;W�p�ǰ�g����)�ۮGy��}2�fn��{�>9��콁!`�q89k�١��˨���r�v�+�U��[�v��u<{�����M��N��u���D��F:�ǧ��ef�W-�}�z���C�Jy��,�����iC�t��e�9C�"����.ʓ^��ZW�1������J��7��Q/n��܍���6�ϼi�9V��*.��NK�3�7�W�Ţ�J7��3�ͧb�E�\3�R
1tBJ�1`��-.�� N Oqo��6�!{s5�Nŋy�g�),��������S
�{K��}(H(���SЋ�xλc�әuIm��O����Ķ5���rv�x�����[	T5})%��qΠ��Jg�j�r�V�R<�.�"�	�t�a=<4��Q���ʭ��L�p&�&q�F�G\@c�Bo:ʚ�3b���'`n	2��n�͗�!��>ȱИO��*Zv�����XU���-����<�_�h��y1u��m�F_/5�r��n/�9��'��L�t��XuC�ν�=��!uՑG0�&��{&C=�aŸnw2�Y}�{`s.��Ii�b8{%9��N9m�X��|x@��nY�c�#�'�`��;X�e����I:Ծ�ti���[�\��B0�i��׻l��]b�T�Y]�7��{t7�X)9,7���ἰ�{�����b>�/*�/q<�`�U����K��bTf{4��q�F�(:����}�����.�[i�z�������΍�&#5ڗ0�W8�M����o4o%E)�G-i�-[zk��+w(r���Nil��u,�9�v};.j��m��4�C��g�*&Xo.T�6l&5����A��4Y�
���rE��\dZ����ټ�Xb%yu�Љ�ڭQo~���/g����:�=�������X+�m���]�v^u��lS���M"'.���7J�nJ ���]�{v��!2���sԱO}�8x��R�=�MJ�Ǎ_����x#�i�����<;Y:\�&�\��d�+��;j	NkZJ8Sm-��I��;��瘬���/I��O_c�/~W6fǰ��qW�ݧ��Tk�}W��iA3���/:c��	+K�OUO2np�=ꊬE�Ќ{�W� J�P��}c7����'翀mv��^���޳5
�m�z����+�-�ZQ�����#Q)��ʾ�_���NM�������5ʢ�ßC�f��)&t4XY�N�v�Q@eI���j�ת4���[T��{��ʲ����6��6����b�c<#�D�"�[�����M�zm��׫n�%���W��S����ޢ�1�c�ځM����ղX:ǣ�K���{̏T�����x�g���ܸ�]�/����Xrt��3��n�cuU�][<���xa��� ]���;x��Xi���{��=��,��C���N�z�k�r��ʚv[�Ĺ%JP�R�q�ʙ��q��EL����
Et�(v�3K��]�n�������Y��9ɿ{
����q�5kAľs�c����h����a%�i+�
W���_p��CM��##$�m��-󗮡�u�M^ѕۭ���������J]�>FpGg\�'��T�����ц��*�e�}����W�Ѣ��7�L�FY�:V���]��n ����3W9�2壼��K'r�x�JN7m�@祛��`�x�c��[�=e���S�����ٗ�眮�����D�{,.�B�ȸ*N׷]c����@�ط����P�f�ZI�&���c�5؊��uju@܅���`t#z����$�W���?jW5����;f̀���4��7h���#_���fӶ-g=S`�v���M�����/0:��7�#�ذ#i�}i�6�P�Kn$RUꠃ!��TkdT���:-���;��p��23��;�Z���$/�'�b��~J����5�T��4C�.Qk��*�uNXoo}�('�&H��ژ������	ÏNY���V��[ǕWJL�s�m*0P�'k��G6_rL���V��9�d�X�(�ֵ�ky<3�o��g?��?�?3�YA���>�AT��p� �A�(���@�BC�?�
'HHHt1P���̇��<�4\,�1���h|LK�WD�'���u,g��UB�* @(��HQ��$	� I$ %-
UQ_��V�c'�QG�e��
(�(*
(��P(��*��DQ"
(�ȣEQEQAEQ@T��ˁl�Щ܉��{�e���-|(=�%I�T�kP� �2�}��Y �R
|HG�o��W����u�:_�!P>��bO��hbY�<<��>��y��fcA�=s�(7��r���/iR�i��B�����g�Υp���C��~�ك�>�;O�	(�`2I	�� �$���(20*�����q���PX�'��@�H?��=��|������3��h��>�������$�HI��'�R���h~b���H`9?Pd5�$4}�L<���o�Ux��I���_D?���E�����Ud�P<����O�T4�����0Lʴ_�~�'�2QI	���S�a�K(�ķ�1�1(�$1��Ő\!�ݒ� R�]hb�!Z%K(<ed*¬<?#������@|}��O��́$���
��C"RD����h$dA,��C�����8}g�������y�u��� �>��ч�����C��O���r�|C���A����YF��g������� I!��I@3����_��d��Bw�!�?�̘
?��k�����X~�$?��~ߴ��O��8��O��?!!�!���t�� �� ��'���?�og�|�$����>!>��������aC��|� ���6"���~s��
UH/�� �A���HI�?� Ä|?�!��E�I``9?_Ԗ�Nx	���ԆO�� C$��h���'@�V|���6�d�	$*F¤���l	�Xl����{��`0�e	UDH��nI1��H��X�?����vj�0Q���7P�2 �QA�?
?�����O�?��I	!^�O����$�z�O��!��e��|�����'���|d>�O�� >��A1��H~���O���#�D,�"�=���6���	0~0�$��'��������I$����}^�O���G�!U(�~_����v�ĒHI
��9G�	�g��������{�~���"	�|H~�����c5 2�����`FF�,~���0|�c�����1��6~R�����b���i����%�0}1_���I$��|��C�!�A�'�Y�Q���|J�3A�08!��(G�>��#�a>G�I��Q,Bʆ��%Q���=����`����>$�XD��BC�!�?h���z���'���\�ߌ���I	�O����M�����}�L��G!@�rT��}���߆�>�POւ��?��|�$��&���ܑN$'u4�