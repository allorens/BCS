BZh91AY&SY��)��8߀rq����� ����bC�>  ���[+-����-5[j�P�A�BQ���$�JF�l@٭��kc*MZ��F���Z%TС\؁f*&��FZ$�kZʪ%m��k"�%�d��U��Ka���������6�I�-��F�[a)&Z�Y*�P��[�{�J��*�f6�Z�Z�6�-!�j��ְ&�k$���5�B�31&lى4��M���,KcZV�k@l�U��e2�km�XʴJiM�c��i[io   &�P�C/��G��Vl�â�j���֚on�ji{6�c��u���F�]�� ꎛjk=�W��QUW���tgwn�{ڱ��&�VT��D�Sm]�   �{�����ox��S�7wG��󞠩J���u�t4�J��Wr��������P�ޗ���=n�)���*��ԭ�K��J�=;�<�=h��-;�UJ�5$b�k	/�  k�R���A�x�ozz�S6�[���
P��G����*S�y.:^��y���{jkIR��]�i�=��(����[jU%^7[m-�������-h�*���RA.�   \�T����]^�x�R��[Ǯx�*V۞��=�յ�e��v@���:=���K۠��^�ަ���Κ��{��;j��w�]�̆���'r���uKʨ�R�l�J�#F%)��o�   ����Wm=���<V�gWa���2��6�S�o�z�TUe=���L��t�ǌ=OA��A�:k��z�us�
ҕv��ܶ�v��7J�
j�R�/l!TB�`�(h�   :���oZ*��Okޞ��:m�{���]��[h;�������z����[V�����)v׻iz���B�je�����t{wz���*�-'��x�^��&���IE�mV��Z�(��E�   {�}�Ҟ�t4�RgR�/k�#{ҶҪ�y�{��aлV�����{`�=y�U)@[�g���5�N���ڢy���z^u�Z{j������ozK�f�H��EJ�U��   c�>��1����/wp= ]���j��(罵�EU����=Eގ��
uۃ��h��G����z����*3b+lKZֵ�W�  ���T<;��=�X P^s]AOF���q@ �+::҂ܷ�( 9Ѩ �5�w^�� nQ/f�K�Z5J	T�|   ��}@�+ >�zy�g�=�6�(�Ն����<�� =ޖܠ��i�ʝ�5נv�Q� �*TJ���2�J�4Ɉi� �L&L�����ъR��2  42   "�����*0     ��
j�P �    &RJQ=Ri�Shb#��F��Ci�L*I&	���h�zML�4����(�?y?���?���7/1Yq���*|�yr+&��Jn��qG���33f������cm���	�m� m�l0 �ݿ2cclm��{w����������o�k������o�1�ccm�����UW�ݍ��6���?pq��j�c`��~?�����������_�����ɿ�;Y���rm���Փ~�6��y����Փ~� �d��; ~�����8�~���&0~����&���@1���Y�7�8��d ?2`�@������`?Y�m�ǲ���1���L8�l~�m�1��l���c���~��������L��߾v��� ~���d1�߬����ɶ ?Y���ɰ`?Y6��;~�o�L���m�Y�۲߬����~�m��!����d��Y �,�V����Ak���"H�y�'�0�ĵ�a�
&J2�)o)�esֵئK7W�ͮ�V���zή�F��op��d`���!�ɴyV�����.�ik�R-�W'^��3.] �Ct.�`�[��(�^�A�i�V�2�:�5kkn��E&���VX&�@����Of�ɱ��K�R�f�q�'�na��'n��6��A����[$�&�F�Y���L�*^��H�[2j]M����ދ� 0$*�d-�5�mԈ��[YPn3�2ܶ���������p���	5�4�p�x�B��z��TP�I��o�����*���C����Gg��q\��h�N�v$�m�����Ky�ZFL��J㽗�Xf�X��m
a=Aެn�)��w�o��P�v�Ù�^�lf������yq;{��ϊ�0�Y�5��G�M���V�GUZ9.�ix��*U���� .dŻ���Fi3�?m�,7���k[��S�E�-nTb�zD���t�*&�(n	r=�ǀ\���WS��4�M��i��r��X��W�̴�	ӁeV��Ù�%����ر`�\.��i����T��bf@X���-b�� T̥��kwl�2���+m��FY��5��V]�O�Rj��A*�Y4��(�I�SZ]d�>���X�[����RZZ�!1!�a)�GV):jm)��/7s	vn��R^ �nGz��!�e^��#5�j\{�hS��P�)�����-a�aH�aє���	�j�;v�����]&�E ���H�����j�13�� ���p����%K0^��u����pU��<+�P��]@�nM�D��
m1wf�t�Л)���*��(C�9���	B�kuV�R��nZt����:�:�N�uoeUT�f+v
N�,��	t��n���N��u�nm�P�݁]�Vs�9�����*@V���U12#�}/	�H�u�+6f�l1�iszs8�-�(�m5t�䶐˹dю��fL��ԡ���=�m9�P`ęۨ�m�Xԣ[A���t"���Xֈ�fH#s�8b�51z�um��N��n��zO.u�&����vc�\ͼ��Z[F���dTh��u���^a3Q��)�q��5��^�+��܆�vΰ�I[���rhܧ)�3����T�8n�3�c_;��NN�J�"��^3-��d�Ia�{��k-��ޙ%��F�X�*7�]�f��v�A��r�j�f���V݊���|���] ����3�V_g6��v#L���Rm�[d�	m<�N��hi�u&�F���Z� �n�3r���L�{�qO ?�V�%	F�ܽ�T��[�]mc�b��6ԉi��eKDM�m�m�h<Aw4b���+`Y.,�M�f֬��j�^�$�i��-8�Cf�h��Z�.7�!6\�T���Z�%�YHa�2�&T%�*x��+6���3ct Ү�"�#�^�YH�����T/'������qVj#^�a��قb�JJ�v*h�Y�u)�&X����NQ���}�Mf�����D�� `���f�+*a[��%bEg+(JrCy���ԫE�j�1X8.[MX��[U�v`?J7���-tvi��A�y4�.5�;�'Z�ua���Ɲ�7�����bْ����4�"�f�M�+e��ٚ.L����2�`Rn�dP'�LkH۫E餙Rh���H��� �o5% �#q(sU�o�l1n˧��l����,�-o�Ԇ��Zr�C�+"�f��P�r� �E �M�A�B��)�]�iݡ��Z�I�ջ�i�����shaNゎ��`�&`�0��H�vԭ,�a�yF��^Hf+��[w6�ڱ��!6k�BU��R	���KOQ�d!�ĕ[��hFXI��\�,j�L���8P-̨�A�+Xk*��VU^�d0rh�pCv�1�!o{@�4)�ٰ��;���*^I������ac55����Vca[�S�O��P�h ��6�<e�ԙ��r�d�E��	����Lj㽅&��,��(2��ǈlHh����1]=�/j�E���1�E�,�+5���V�2�K�T�ݼ�Ï5�(F���
mQ�2���3!�.Wf���,�(�Z�a���cm�Sd�r<Nw<�����7�r�{����{����6���2��O"Z�i5��K�xU�3n�ts3h����ܭ���5������f��,��4�N�j��pXt/�P�V��R"��jM�����#&�J;W�ka�ӛ�CnZ�pVv!���nY��8�����)��mv���t�Kk�]�
�}��{��*������svenV�v�W,V^�c�䐻��M�&��ʖV~�����a�a�#!j�)��lB�i����Ē4���f���2]��,�tjؑ,s-��S
*=�@�6�^�i�v�Q��zʒ��2�5�5���xRݼ�CA��[z��4��5L�P)� -ޅx����=�u+䧅D��kbT��F�֊�uuta�S^W���̷�c��Ԛ�nl��ƞ�ɵ6���ԇ?��O�s���+l����}��oj��S�=��K�{�JO�{h�dֻSb�E�y����$�RY��N�/�m��/+V�r		JF�,א! -;a։��]�oa���룪-�m醴O��6�V�[`�{��v�S,VݹQ�N�O�W���V��NV<�<�""0fRj�m6�v&
�ҕ2�	��-
U�LKu,�L;2=i����qְ����;R�?
צ��y7c$r��X��rH�u�����d]v���8��t�*�<䨽18���'(8�g��.nZʽbZ��cT�^R�q����`4��ۥ*���q��˃6�Y&�b�j�I2��)N���6^����I,=�i�XK���`�j��v�n�F� j�4��xDyb���ø��%��68h�5p�4�c%�**î6�P=�RcY�7N��6���2ۼ��֦K���{�AN]����:ǔҡ�8��L{��6�R/q�nm��.AT4�R��(㉄�Bn%t+q駵���iIb��=�Yiq�r֋�����'#������3k�w��Ȣ�+%����/v�dӣ()xv��Y��f�ED@Hl����F�voH[޳���n5ڳW���j�:.�#)n�Wx�g)t�����Kв���Ѣc��3`��9��
��ڢYE�*�a6֙x�l6�m�vi2�ȯr�2�ӌU�v�'�Ö��ʚ�?C�Q���A�oc����6g��K�!G�8e�%��u�`�������q��QB�iMUzQ8�r�h���k *2F0Ka�ڼ*�63��^�cU2Z���v��m��ɥ�s
��qV�s-u�ׁH�,m
�}�C�yCȕ�M9��U$�^�BX�,�1j��k^je����+J6�j��,i��m���r�c���}j��6m^���@�5�K[�/u� ��%�x�/t�nS�c�.�=Q֌QV�{�3�-n�Hբk��0�I�^j�Q����k(7�t�7Uݜ�w&֜�p��W�&k�0�8���^[#:čko/p�FD)�a++^���	��(���M|�oƓ�V���(V��sso&!z����Pcn�\YKpIF�3�-�B|n��wp�2�S%���,!�I��i�n�

�'�)� nL��Zolee�K��T�v���p��xY�Y�Gj�������P���n��*����b7�ښ��kr9��=.�Mu�+�{Z6*�JTi���oVctkf�2f
 ö:F��W2!R�ԗ25�ic�(����r��ec[�[�_���姦`����OB�gZ���-<ͭ�7��P߲�Ml)�-�+EӼ3D	,�4ܖ��xĒ�H����cJ�z�rv��-v���B�:k2'U1������G4fS����n�V�� ���<Ou�s"�L˭$j���p�)«du��X����Ƃ������Vwȝtܚ�!pl�ba��w���ل}����u�CÏUm�n�%�j&n�f�/��a� ��eZc)ڣ8V�;�M�rYǔ�iBJ��A��A+u�.�0��N`�s/�@��Ԏ�{Y��'l��efF�fVY��ˀ�n#��� �wyn�c�c@��@�5s-$�c"��l��%VGMn*�"wC	f�2�*����lm���9k�&��
�^!�`�wai3cn�I�z��YMd�@��L�c�#��]��j[�Uhi*xA·t,u�ҍɤ�,�"�\��S�A��pK�X�C��j���T5k��0L�-�y�[yh�]�ə%�L�zU���CZX�hثhQ5	Ѱ�Q͒�o�FS���.ay����bL�[�W%�(�nmn��-`�M�ʻ�%�Vv��M�ͩ�7�^�欪��.�2�4'��ăo6Q�17�jR�OT�vMN�3X�4�"(CwktRוD[r�@����e�̳G~��*��_6��1˞�Ÿ]ц�P�v+c���
f�h"�%͛��+/+2GL������lz��I�ĤoZ��#���$ ��e0'�k~�oe3
��7[[
�V����"2�����x�V	١Y�e�'m%�2�����i�˭*�jŻİl���0�M�����T3we�c!I�y�����h暶��+2�����QTB�U���줌J�y�s#1<r-��Wv&�w�6��%7-����14v�#�75M[uģ\2eԘ��F@̇jƠ�멍�� �H�,m^U�U%!�,�;K�<�)vci���t��G��ʪ^�#��+����T���V~cF�/��qw�H����FAg.-�V�Lx�,ⱃBE�E<��3c6�p��I0���c��|LK7��TL6�r�5��+����

%eɦ�,�%9�-b�ˡ>���o$�ɶ��ƅ'z�ձ��x�JҤU�8Fb�̦޽U�R;6�U�5�bm�࿮��+n�c
��E㩧e�Y�tI�j�p�wcP��xĶ��jSeLo6�a1t�1U�V��Aoc�$Vr¦݃����e
��m趴�큚/,QCq�c�hJ�jkAE�5��KoZjꞍĵ�l��ngY�r���;Y�R��&�f�1�ݺ�w�(X�C�)��A��&s1e�iZ�z��j��eֆ��(,sM�@զ���\��H�-��U�:��똲�
��:ZQ�oCs��f۲�&�ؽt��Gr�U�b�R��e$��,Ј���)Uc�I��K�X+0�Gv�+ZLk�z�6�*��bp�@aZ6�[`E1�7yu��d�F
1�)��u
Ⱖd,�i��n٭Yp'�L��2�?�պx���%̻��Q�n]�r*��{3V�7l�j�q-@��Чa��k+
�rم"�m0iM30�
,���(�w�+I�LF4�q�4���w��*�\��1ǵ6e�zmά[ 9c�7h��dn-����Y��V���b�Zdx�����M/�c�wu��Z�n��ѳi�r��5s[4eʼ�+�F��������3�l,�7��Y�zt��+P[P��6T�ZwI�0�w6�k���qS����;Z�.�%�%g%Y�զ��,����6�X����swS���:X�!Y#Y��;e���pm�ǐ|��Ûm�u�I�"��CU��ԁ�6Ϊ�%t�QoUe���է(=tLM�,^�3.�yB��0������N�{0$(C���[�����_O�n�V+1(�潨(�Tڛ2+y2��0ώ���[�zYa�@���S[���J�wub�i�%����B�fU���E["�n��B^��ZjÆъ7{�BO׺����i��Ǵ��M��/ek0d,�4r�{���:ʲ\��M�����ڍ�ؐ��v*�@�
]���1P�n^9��X�!��^�k$������֐� M3
�[�[	��6��*;�[��n����/w6����V��֙��oE7Kn�T�1<�s6��]0++�]!��+h�4eZ.~-%�j˽���#�F��?e'vkPyz\s$ݫm�,R�U0(i"���Q��!L�lL��i�w�ލ�:C5廴�[�8Z����6E91��lH6��;m8[R�񭵨kt���v������4-hӎ�k^����5���1���f��>�7M:5E<�LJ�)j4`�M�3`��kq�mS�X�)1�:�n�� ˫7oj\�Z<ɾUz˽Τ
Lm�آ���'�˔ƚ�kaZn��RO%e�4�IJ`��V�!UK��u�`�͖1��sϝw��]H&�o+�1E,Z؅݌ "dv�ِ�r����E�r��$�n����J�_�3]�.�V����X�56�o4�e�ճR�YM�*e�]̤)�UXa�қ̆��)�Ual&�ҡ��sF���t �{X���z�q�SqV�DКmaDf��u%���f�Hn��S�I����+B�mOѲ�d �	e���1��W���-�F��x�lX�V�6e�Z�&���1����KjSe^�gb}�Y�����ի��)h����.�61G�N�a����Zk:(�8Ȇ��T�@,�s�f���!MGQx��ֺ�r�V�7r�`�J���X����&h���o>g���cSAv�5�2��m�/m���7��ow�gt4�2;@��V�61a+r�&��f�%�̈�b�<�*�w5���/��]���-,�[��f�3hRQ]�d�F_�ҥ�]�2m[�pf֣a�~�] �h������gR4W�
�$�z8�OJ(�<F#�"?��>�?��^�&������8?�p$�{쾶g��w�^+�yc3�O��`s2Ħ���G4�>�]W��'r�׳����kS����	���gm�̝�rg�X�%c��hy	R.rI�WH��I(Э,�QF�r�K�t��@�b�f̢����\������I��X���Y�\��fP�w�+$�b�n�_k���N`cf�9z�F�9yJ��|����Nس�_+���Y�ݮX���Z�vED��Z���!���}�rQ������;�;���[$�[�}��ktҫ�r�YC�ǐBv�[�3��Y��e&�D9ZJ@&S��|�"�+�x������\]�ֳ�H��.�q�V��a�m���VXg	�tz��L�!�5���ïp1��zdl�<��un�S"�Q"	�c^=<`��֮<P�J>�u����̽Jn�Kk�kj���b'r�P�ݼ�%b�e��Ju˝1f}�D��웆ؾA�fG���b�̓�I"K�r7�"�P�w���K�_<f!y}�7C��jVb˂Ȱ*���d[�0��}�1�4l�:݂w��Q�b�&������J���K� VEG3+^M��㻵��g\���ޡ\Ǻ��R�A�w��
�Q9�b�`�r�9.v,��:�ء̖i�u�v���q�`����T����m��x��{CQ�k���u������wT�aJ�Z�Ƶۘ��v�g
���%xd�j�K���+h��:�限:����).°���.��C[�0:��4S](u��N�e�7���)kLk����]Y��q�%e�̌�v[�,^u��RGM��4�v��z��v�Xj�"$��˭ ���9G1����nv&��3��|��˝amB-)2�vov��nBT�S����ޕuH&�N^�F���'1/D�֒8:�8������*"�����Ԏ`�82��DFɸ��
��9`I,F�BQ�wky�;�ǃU`�x��^:S]9K��s^�ɷ��RDȄ��90���p�����j�[:��F�j��mյ��Z��y������͕�Q�Y)v>�'k����f3��|�j�1�v>�x[BGi��Xfv�5�{�:=P��<�vN�j�Wd��g��!��SѺ��ז��l˝��=Ps�}�,�4�tԬP���֘��2�1�#'N݂��A�)m6ze�cK�nT�s�k�+�L*��[G6v���ʴ�)G��vl�T�9dvggl��e$X��2��)��ؾ;{G��֛0��Zse&ҸyWֆ��Ǝ����X��H	W`���N;A�3�)�ޣ��S���Ar�WpnPSA#�P}J�t�E/��wR�m�i���Ḫ�슈aa��[{|7��\ѓ%�9(�i����ы]FE��(=�����;zr�7Z��C�]z4K��ou����9���a�y����`W��3z�gm�w@����II+�i�U��"��o2o_gZ&��c`G�Ҥ;��];8uDh]�p�S,�JZ+��)��9ϒ�uVJ�@v)P�;tl�@,h��X��iɭ�Nn|)�M>�4H�8��R=W�8.�RsN]�)$k��/��Z���EQ�֛�p_)�v�<�� Ju����
��z�pd�R�9�PL|��XB���*R�r���V���V<O�r�Wi��.n�{D���6��b����ɩ���h�T5�~1��j�:�z�ͤ;S}crnҺZz=7Dpz�ݓ5,=�ȫr9�f��r��F�*�3:U�k�MKO	4���ќ���SK�\1��
v��p��;��5�����r���:I��ʓE��I�ֲ��em���z>9��[ν�Jp��%#�]��"���z{[�u,܃z�WR+��局�I}��j�Κ/��"���bP�����aKi�;n�+yq�41�6W
�n�bP�O$�e�q�á�;k6�j*V��g ��K�+wm��Wy���`i��p�ǂۧ��)����[ZWb��1���`Ss�
[��me>�n�5%:��.;!�u��Ҵ�Kfl�A�R/�e�0����Q�}Kʓ���;h#��;����}��joE(Z���Ck;ɘU����i��	��e���P�Ҭ���B�D��� �g�z9�&�o��v����ޖn��f��dh��*q��=D��r��Vo{AzH�Cd��d+�p�nrJǁV���M��6-�9���}��
����򹲈6��]4�k��S�n�>-����o�{r�`����^m��u��q:q7k�&�w��
��G+�,vy]�W%�T��ގ�0��J�nE�֪o��b�k%�x�i���qRVq�`���^�ս�m#Y&R2�E��9]��p��������`Ka͵�uX2���\Gp��"���r����T����(%,��_ �k�z�7�.	
B��b\��fc[������'P�FBM���c���>�&Wdl�"r�k���_�7w
Y�qX�(������kB�s$���x�x�]�2J��VU�V����c@�yq��0y����u,�r@~�;�gn�ֱ�8�[9���y�]���@��,4P���FN�k��;G7k�S��lW�m��r��} C	0-i�D��7(aR���Z�ׄ7i��{�������xf4�j2e�95��s�h;yKmn-5r��6�KM��HaJ�7+^:�.&q�o�k�h)�W�]աn`�X�\��7q\�C��^�B�SmZ�+��ͩ�FSJj��B�Ag�����5�ԲY6�׫^[�!���
{�g��I����� �i��μ�5:j���<w$�M�0�u[%���7c�s*�F�3ӥ�q�yn�b���[�;���P��(g9��!���Hɽ�~��LD��1�e؛����S�����4l'���{N�_;�V(�EY�!¨n볩')�;��[�,�
�<�Q^r� t�)���B�����ѽ�ټM��b����kG"�Z:E�ܬ���]m@w����E�/#ڂ�)B����2��t�!�VU�l+���b�A�Q���
aK6����"V2�*|z!N��˩<.W�<���$%v���AEi���M�fث�z�䛜o47�96^�l�}6+ܥ��u�)U��`m<cN��x�T�d[�80r��e�$�)g�ڛ������Yqφ���N���]�.��d�,i���
2l�h���6���Y�a�]�Yݓ�3�&��{r�R�b��.��q��L�=U:w[7�� �`�W�A���1*W]ʱ�q,�\���V�ι���� ��^sZ�P������.ى=U���[�x�k.�RC��W��b�ӂ��2���;n��ݭGb�rnV����p0$�����P�ə��NR�҆���\i`T��oRuN���r=�4��xc_��w$��Z�(�r��q#W��k;H"��j.��]{��6��	U;��DW"��[3���ʟZ�S�e���M3ӵ�Zz9��%��؁d��+{)N-�2�i9¦�0qn�����.���R�40X��B+&]*8�ܻ.Δ2�5OP�(Kt�Vw2+l���<�f#r�e����z����n�1'�,댖�J0��)�/JEj��a�Y�Gs*�ڝ�����v�Y�g�Kga��!E��a NǶ֞w,c��G���DY'l�׶�����;8 �h���K=}S�ӆ�i�+� N=��,�Ӻ�1�4�ݱ�� A�������LP!��y�s}��<8��.�+�s�GYB�F�k�t]�wͧ۰r	Q/5����w%nEE��o Zq�]kR�]9�6vɕh�fN���+� �U�8���m[���N8��ls9���X���|,b��&Xܽ�&R*�V��ۿ�����^��lJNt�X��qc�X��c&�ے��V�b���A�EH���ڍ�ϐ��]�5�8rbH\j��� ,<=��gX����M���r.��y*кdTqK����ǘ�m�tJ$+7]ܰ�Y�έş ���ɺ|zjj���2���Ӑr��F�sM���V����+g[}	���w4iN�1��̗`v ��mgiW-�
Б��~�s��V�)f�i�6�Lgt�;����ɴx��Chp���h4 z�؇^�2>�
u��^��Y/p�wP�4�m�{�������XUkG�ˡ�l}1U�8)� �I��W�b���l��ǟ]<�1��u*�0Mٱ5���l\�L���ݥ����+�u��&���V�G9j��Ԅ���`R�b�GH�錾�$�ȱ��7qog\��$� N�k�k�V��p0�$�l������m�ud��j9���9����U�=�_�p�$˔F�B��%q�S�N�Ni����V�BD�&���M{h���B �}�Z`�f������^s��[��p��%,����h��$��78Z��r����:c�{v�,ʸ�]	�:�7�\�� X��g3R]x���(�KuKRh�ܳz���jp��cy��r�˅�R7��O�u�V-�����[h�=�S.�ц�Ι�!F�� ݑ4%;���_��+!w��i�b
6�'��fl�����T�ޡ�(�|�
N�ZR=�7%�H��L��d�ڬ{;K���J�1�喡��3��!B/6D�8���x-���EJ۴�z��n���&�b���4
���g%	VCt9�����9������W�;�0t��"Z��3�2��eg<i�nՎ l��y�TB���|��������-��ө��OdZ�,+�4��7�)�H�ň�}��U$��*gC��2�QX���3��������cؤ��o=�d;��8����81�򭭻��ݐ�咱�"��H�;H�;�kW�>�vW+T�L�Ա2ΙzUYW����`�kZ/��3'J|�<bŽG�iU]��A`�x�WUɷ���U��*��kR}�X'@����Q���r�D7(�R��I
]�$l���ѵ��R�bjӽ\�vJE�r���զ0��c���Z���p�:�P��1��}��f�k�"�H[Hk5d���mmG4YAjlPin��?�\c��r^ hpIa�ո�`��rr��s�߱&YO.��2v`.��,�E��qȆ^TY{�=�I+�F�E��b�N��Wl�	�VV:�N�d獈�;շg��a!I�se(�u��BEۄͬ�5£9�,����+;�:͊��7Lɚ띾�� z�k�y0�i�gN;�d[�7S`	M[%Y��@.��xRΊ\W��=Ƿ���n;��3�3���|[W�싆ĝ�Xd[����m�)n�5x*3��-0�u7��g���Gn���n��h��+5�[�g�}�N�IN^&��7�;b��u���t�ŕP�B���zю��fsjK��Si�n��zz*Ovs�R`w��-�����E�8��.ѯn�)�jBᗪ1�������,RY.�f'�Vt��b��wέ�s��y��Z(�\�]/��zɗF=��Mʂ	�p�:L�n�M,K`n��X���"�W�J\��N�f#�6���8=�́X��U  �'��]���'s��^�m��eť1G��DM�Z._!��+ D0jM!��3�W.P�"V×k5��c+4#�:�]K0wrH5�tۡ.�n�a<IV�j�����6����w��\���c�k�j����_Gs�7B��6 ����v˨�5M,�9Wt�͔��c-q��[(<��pg�x�$je��K��]��a��Pxyҷ]gk������Jxnz8�9&�N�6,��Ig�tJ���=��$�N���f�q��Ue|�%G��2wqՔ�WZMvC�)m,�|em w���6��z5�Z�8�`��*#��kn
Te�aw+l�u��w�q�%��U��W,��Hع��]��ð�>��!��RU�Vm`��|�%��c�w'�VJ�)np��\�ֺ�
L�1�05J�*ǝ��{r�V���C�=��S��%*�]�z|�t_;�1��8D����&�ڮޒs�)�چd�zp���.8��Ӿ�%�gQ���4+�U�����!8�n#�hԴ�'�0�7s5�����{��N�u�˵��t��0m`��u��/
y��j�5��t�(�<ֶ�<[5I}>X�#I�f��u>Yݡ,w��*"wv9��L[}c���܁�ɗ9�r�Ÿ��ط(^���ن�=�\B�.f�^�X{2a]|Q���}�5��٘�p�˟"���7��V���2_s�Yly�����s�^! [z���Vr�hP�l9\O:h�ɇ0"�LIoN��J.uϬ]�X��e���}l�#x��`�h>�&]IS^�&�Y9�kr�v���X���
Ntޜ��ގ�@�fK�A;gXM5���2�<���U�m�|.�l�\qӫ���h�^�,��K���u�;�*�x��M�a�[ls@����t���	=ܖ3�*u�e��=mU�b��CvLi�O�ćʧ}�o��<1S�*��z��X��J�K��yt��ʜ�����Vjl��v��N+���;�VhfS*�Y���)��m�Μb����l�������3���M�s�������	J�[�fJ����QJ�'a��X���eIz�6I%�dr���)kr
Wx�S�+q��ʒ��U�.P��nk�.��S�Z�]���|��c��v�k$�ntV�6�].�rl'�b�\��6��]Sua�tݢ��Z��l-��&���Ý���%�^�)�&	�g#�QI�;���Ů��$w+/U��;�������w���ǯ��b,�.�C�����噊m�9K�1B5���*'ΐ������޺�����"�Sg,�We*>8#��~��||p2$u��}����u���0�ϻ� 333|��#�9��Հ������ ����������ϡ�������������W�]X�S[��4��rUƬK֖�0��q� �8'wuw�Al�}*w%��w,�䷙�P�ݎ�Wr����kԐ���=VC����Xp���'Z��l��^��2��[գNe���g%+�G��r�fku�؏+h�4���?q�n#�5���wn��V�/���J��p�rb's3���cO�hڭ_|���r�H��X�w���m����&}6����nU���7R��}����n�nL&�a��\�w5������9�8§YW>%�k2 �y�Վ��D�	��A:Ͳ�q��w��h�j�k�ΥVje銡i����v�B�Z[�S��l�J����]OP���&hc����/6�ID�<�J&����w�̛։���^��,*p��)d���^��ЀR�{w�.�ή\�*e=���TԖ&�d���+%�^�!
��V����7�sF����&���c�2^���3Z�n�wn��mi�;�T�'xT���Q^�V��姌���u3L��\��;
�s:RR����8Nb��ov���tT���%�}{�!"�`�T�A��3�>��E�hU��UVֲAƶ�݉e��wb:0F3��vp9*�l�]&�V/`�UQ˼;�.�2m!MQ�:���bw,�(Lj�oi��P�%J�L�/Qj�%��V�JDC�9�'WLH�W�n+�J'5��܁��n�ցZ6=v���֙���AK��-�ĳ����¹VY��ֵ��C���lpm}�^���&���ٹv�R�'����W�s0`yc�v�U�a��{�k�shf����2�|���.�/^��E�vbW�d���u�:n)�K�7�hz:eN+'Cףy��,u�7d�-�������V�����[��`����\w�՞f�m�_9՘�U�����B��{1��Z7 ˙�L�x�L�*�dȺ���Qmh�V5$����)��sx��]��xd���wkx���pWa�6ﵳ�5ρ���L�6�E����uХ[+�c�
a�3���d���)��i&VXB���Z���eǼ�^3��H�v[[��ʝ��Î�]�[ׁ���(B*J��fu�ȺHM�4��4c��T"�ʽ�CXX�.�_���2�P�P}���-��j�<8C�f��}����3m���֌���a���;t7Q�]�i����S�Z�E�Y�bc�$x��A�4�O�έ\�)�h���Q'��MĨi��[�L�Ōfb c�JC��h�j�%��SŔ �4=�ʏ�o*$ә׹���+��țp,_[+���`�,-�(pt�N��`b7��ŋ����|h��=�a�R�;k�y�����)���fWd۽���-�Y�o'�]s�s���t��其����^��rv�G,q�U��[�-A`�ʚ�9�j������Ѯ�WC�$
�M�4�5�[G(K;Cbж����&�m��QY֝��W^�_
��b�l�:�y�K��=��mν �����<�Nw�ud 68�N�]p�=��~�cyE&�h^i�F�-l�.'"�Y��6I屙��x����1���A���|���M�������j�r�aL���G�L"�u�;���>�ڴpn��z�8�!�:M
Hn�R˧˷�t�Y����.���d+�P5��#}��<��#�RYD=U���:I�V�kP��y�qo^��uw);(�S��%:۩.n&����gUKi�Q�!z���O"�X<(TP+Y�u��W��^��lp�T��v��o\6��Mg�(k[2��t��ᲅ`Q�G(�󳉪-e;H�@r���L<�ٳK�k(��*��Z���ɧf��ѣ0'W�U�aΗ�u��9T���Ɉ�Zβ�<�)���2�Y
�v=��}�/v�(�ԡ׮�O1wh�7R}zX]pCV�bITɘ6d+4��w������e��B@��lN�k����=U��q��l2h��&!�:��F�;����	�]�h�Ԇ�.�0�T�j�����T\u3DO��X�0�s�x�>U��G/�Q�WQ[t���:x.J�UN�@�Ј����ϕvX��ۛ���Mx:p���J��Klfwu�zЊɴ��m�(�@r�L�D�HtTR���2��۰�V��T*���ѧ'o@��\�k9������n
�(�A#���UyV¡g�)��i�Н�=Bj����k.�.����X��c1�*.-u[G7N�Q�X��l�C��p��؀�:���4�c-���iX�[+�Q��ޫ;$p9RovmP+8h@�>��S�N�_�7��-�)�*�'��n+�0�r���s:�uP�.e��Q!��v��V{4�v������P�˥鏧XtnB��َM��K���Chkx��eO����S���a�HIP�ح��w2�E���pt�;Xq���;)<�뛎sg�Tb���.���gWw��	��'x�l���|�&��N�<"
۵��0�t���7��V@;�N��h-��l���&�WXƥMS,��{y�)B��Ϋ���g�����ʔǮq�y
;Yo��X
,�%E��/l�J'�=�C��y�Xd����ҕ��5�V�]J���2�Wd�Q�%�#��E�n�,�7z�()��h1�bە�T��XDޥڊ�%S)��T�k���Wn��}�g����Z��I�镆
��+ou��frh��u���C���1R�,v��d���hgvBYgI�En>�Ӳ�*��E��0�]�[�;1r�scb��|
��н6S؃n2��L��X]��)����(�
��c�I�;@�bRor�������o]N�ld�ЉiF��ݲ�/���A���n�DT��k��m�É�"�,�f�Q��������#ж�8��!}��j�"*�L��o+amof�Ҳ�ri���ۗm���[��5b��]�&�q�3s]���M��Z�̬[ .��}�V�A�s�hK���B�n�[��u���A�i�w1	a;}ӷ��J�awf��hn�U�� �y�R�d�[W�x�yR�YE�m�*<�T�oYRZ��c@=f��^-�E��W.ē`f�7lCkN�aF�'��]�wv�t4�޴�	d�,)*�9��@W"F)�U)���h؝�a�K���b"i��YFݺgK�-=��#��,�"9n*�5Q����|�D�ʻj.r��˅����<ĖQ"�E!N��Lѽ��K�w�.�Y1=c�'�}{�d��t7��!9q��Њ+���Zu-�*:�WI�K��հ)�Ѝ���vU���t#��
7�8%�������X8Aް�ߞ�a��G
�oi�:\,��˲���\7��\�<M�u�e��/�b�fcɁ��5w{��wMt�n�ͮK�o��QU�Z��N�E��gweKu����[D�!���}�`9H�h+��]z�NK�@��h�JW�u�E�:��<[�Qf
o�άuz��K�W�`t����=Tq�r�:
w��
1��l	/(;V��Y�2���E�\w���4��Eh1F�uj�}���oT�����b�s��gcҡP*J]�U���±&m&�<�q��N�ິ��m�S.� ��<W[z�g�#Ci���u���]��v�L2�"�F�*2��:����tf~��t#���cy�)��$%��S�ϲ�D�76T�.�-���Z��d7f��Y����꽶���O�GZ;t�P^����)�H;�7��.z�uJ
��\lB���$mՍ���d�q�z��̇-1x�Q;�TQ-+�l��Y���1�c��A�50���6U��f��e�b놔Ⱥe�x�{s+��O^"ުS{�v�k�m�t�mK�ܪ*-=3�J���ŒQ�42�^Sat5s�-Y��Ʒhҷ�\V�������1i��"��庘�����l紞��*���'uc�a���[[�&����t����l�ehbӏ_wrɰ��a���!5���	YzU]L����蹈��%ch��A�@�+A�v�0Ѕl6K��[���M��2&��Z����JӏF�S.bX╴谸���[�Wy6���
�w&����kd��ݧ:�7��#���%�hޗFM��y�v�&��A������uTSȟA���QѬz���Њ��C\���|>���9�GQ��;�X���ĖB`�ϴ>2��P&�jn٪�P��)�lsf�J��t�76�� ���T��*S���+��x276�����m��<t�ֺP�y-5�ca���S㒦�Ɩ5�1Ӧ�3m�VR�|LԈ
��:�[-��N�lb�\�
�ͭ'l�[�n��n�K�O������:o1'&�bg80�V���*g1�3y`
iq�r���� �%K<l�&=ʎ��؁ǡoZ˳]+C48�k�ӳgr^�F��V�`LP��ݑ�M%ܕG���7�ߕ��(&4\�s&pǃ�4(F�]��Pݽ� WA!Gwm��Q��y�2��ą�X�Лu�W�䤛=�d��d�!�
A�Uf��ZO^���[O��5ۓO.Z.
�,t+'@T2��`��f��/4<��M�S�P�	ʙ��gW.3Oa;df��V�-�aۘ�zV�U�9t�]�.�7P�Z���ޤ�*�f-���uvkxr��f�������-��<�;j��@�_1&�ӗ3qЦT�P-苧�{Z��[/#�}����4��x�n�ƪ뾕I��A����Ϛ6`�*_=�m���+k&l�D�w)p�s�j���[� ¦��:��w*���K�q��f�7�5���@��g�ȅ;����o�qOk��i>�$%Y��K캱��	ۼ�VDΖ�H�aʖ�a>j��Y�*��,��*���<��\�䥃5��8-�(�ԫx`$3�����՘Lz����(�kv�<O��[�O��MDzp�M^Z|]��ܳ3��l�^�*�vM�C��3/U�j�[�	�<�� M;���ӳ9����A*���Js7�%L}u��ˋ+�mCZ�\ɽ�a��$��4T͜k�p��T�o{�_���p�CZ��q���i�Φ��m�6���\�棻90\�:*
7gs�^�-�"�Ѓ�d��6��g>i�e�Q/ú�v���:R�,� E���=���cU-��	��<( �>�s7�n��'QЯkJC��O�H�=:mp ���<0�̗���t��	� �Ye�f�1f��vb*��ϗPF���ZCk&|���2�b'klwQ��6n�P�/n�Q��r
ڐ[0�Q��:���d޼eͥ`q���C��S�7ZJ�+T�˔"��)�N��ǐ�EIM�s���]j�oλ �����I�W+��[V�p��ذ��AB�K��GT�v;�+Ss4j�,T&����kOV�z�塒Yݛ�Rg1�c�Z�4�u�S�5�׃���z��y5�L�{z�h�D���<x
%�����|t:,�G�2>�S�F	��U�L7w�ǩ�C�̃	��Y�}u|&��K�(37Y'��S�)l�|�d�]��F�L���0��5r)�S�ur�Y�Bb�RD�F`�@iTi^�f�8������^0�^��J��nȔ����@��[�^����v�A���:4+�Xq��-��%�)ܥC6�a�YYS1��R������=�C3b�T�3J)�l�v�c��WL�r��o1J�kH��r���Ej>J|Sy=�D;G��l�<�S�yr�6+�<W!�ˮG�]츍���,�f78�����yoē] 
�-�����/�LRoݸ�أ
O(G�\0��2n.��u���B�j�2�gP�p�u��C��To�Fc	e�mحk#�z���΄��U�"G[�w*���oH�&�+s1��Tv�E�k'����J�~+"����!�Y��H��PW��7H��F��B��\��v�xڋ
���)w.�٬�N�g`��E��(�j��9$t�v���`峠�yvv�F��D�����7/��#XDu��9Ykz�vfe��ϸ�gRU��TkR��0���d��iSPU|����}���w�"���� ˺0.0�}�J��خ�Gl5E�G"�"�A�J�	�-�P̃O3df�0��=�Q�|�.�p$wv}�6�ޙ�⬤�m�s쭶ބe��A���D�X�.q.��Rͷ��m;�T�)�P���ä'	ۃ�T6���+VJ52f�Q���\��fݦDsj���v��47.R.ЍX��[j��]�F�Z԰��̰)�avj%�.�,L��d���ǵ_��'(���� tw��j�L�^�;,\�A�p9+�nc�V��Vi�c�2<锾B}�p;S@W��հ���&n+&�J�O\u�-��m)U��*���ި�vp�R����Y}���q�sG`̣�<R5H��/�;�w���O�����G ��]Fs��rj��x���LQ<�b�'k~&���:�pܩ6+p[[y��ӂ��4�}���ս�w�u>�S�M��e��]� jmt��f�!�&r�0cɐ}7euNy�x�Uk!p��{�x����w��p��>i�S��u˘��A�N��(AY�>].�:p������¡6��#�Gl��Χ^�V�'>E�cٙ>�����
�@
9�Bl�4���ם]}MP.����Z��iQg&�ky[����*����Z�\���1)t|�}cE�P{|nq�ÕbU�H�ϛ�������������w@u�x6�GPi��M�M��O�K���נ�)��M[ə�zu�^-�	��&b��ҪCt.�p+[�HF�W�;��"���JMw��7�s��#�ي��k\�.�.�ig%��ڰ,�QWoN|��6����Wh:2lO]l�^ƨ�I������ �30fbŋ??��_��?�����}��&�7�ߓ~��������ш~�^�%��fQo��H�C����C��c��BU�s�ٻ����gt��,�\f����{<s�@���rio����LJ�{��:z���������o}J�V�6i%;R���[��!-0����	k��9 ��5Vgl8r���:��6��3G|zIJ���8;�o8�:�ӵS��W=���V�GV��I�����R������+R�B�Z��d�{&"�wK���ШM3u�S�7#ƭT�+��Ֆ6�>��)`�	��[YT�V��.T���N���5��K�;V��ˮ3���'�Xa���J��pl}p��.J�K2h7ث�ğUQW��\�ĩ�pNb}�i}77{�p��d3+(�j鹑�$���6�A����.r�ؖ��z(�4�LCn (�h]*]�O58�\h�[,����-k�ޡ��9˚ �[l��2:�@�(v��;�Aؼ������z��q4�̈`�wFոXj���.�/Qy�;$��Oj�Cq�X� �u�J���\��YJ�`%W����X�һ7��u��5%S�Kd֍R��9�����a��yG[Q���t�j��w�hf��2�pE��o0޴W#��2+���Y�tf��X�0gV�}Z3&�)�r�9VE3���fq����j��c�0�=ռ%xxQ�Pd['1i턙��QϞ��RJ(���зPɸ�͏����}�Jx�����w�1(�s�#����q�s|�E*��9�Y*],̝ЦS�̴��jIE'���K
!(館��7�%rT�M��Q+y�yiYX�d�|�35d�WN,�����t����,����#R������P�X}w��}���.���'���e�~3�Uk����C�t2�+�?:yjV���-�>O+�$����څhR�(�*�:���o���}15+D�����D!�_{�v��{��>��%���S9y.���x�0�2���d<�34�Jy�Y4%\��E˙��#,.Qs!?{By`���r5�g׺r?'<����`fp���r���Ι���E~eNp��)����%rs��_%���$��w����5UXYN�NQ>c�rK�'D�DNyܵ�{�z���=��!��~��FU�V�����?�Ӿ��^`�-Kq��:��&� ��v��;vue�kb��x ��8j�3+:<�3��r���Uv��DT��/�?��{\�Nh��>G4��\�8�q��'��DY{77�L3�^�������_�}��^����;���k�8����::i�����'^̏������F��qZ���^���l�#˕�+�Z�@��FX��et g���م���3Wcr8P��ݤ�t�J�9�[/c/�<���+����_�*W�Y*(�<j�xV
U�w��2ƞ�}ѯT�-y���gƼ�f�3堈@h�N������-�C��ustP���Id�'����/T���u���y^�5��|��$�״�=�Ql��>�7����ů��
j��>835��gD�`u�f���]-F�)�3�����{G.�F��ٱ^J;}�T�V��ۓ�h_�tW��Br=�=�QIqR�ڧ13A�'h���r1��z�F"�j,`Q֚��E�ښf��#����(k"{�����i���'6���\����
5Ա�vh ��j���Y'\W�lB^�G{7Ҷ�uxz���t����lN�V��
Q�΅n�sl��	�Z�/&.�zg���,�@G���
���:T׳�����'ތ�����ļ���{`��Xח_��3*�������tχt�S���z��ˏƼǆ͹de/}G�ٛ�3N�����t��i"G���G�E<��{���q��Kz�g����&�.��,.郖��5ꌔ�|g�K��H�3�ѻ_�³�Vv�ԇ�!�凭.�_��]%��Q�R�U�Қ�,3��s�������	M���'��}����Ǭ�^��br��ˤ���G,3���N���K,�����'ݿW����Ɂm��dz���\��MK�^�6rK�<��?*�e��/��>�~��FS4O���=�;�@�xj���$B�Wˑ"t��W�����Cّ��7	�>|nv�(ܓ�R�����O=���{��k��3Rt7־��e`~���J�� �^�M�ڛ���c6��4Z�;5�|�Ab��3�Q4�+xn�j��z��;�q�J�x��p�?G��R+�q��\�)U�lk�N�ҫ3;t�b�
jN��;�IdW�^��Y��M���||�|ƍ���;�g�jԛ�N�xq���m����;�lv-�QZ�	+�T���!_�O�;ۆ�ɗ�8��>�ﮚ�M�x���=ؽ0��x����MV%qG�]�׷W/z���7(��v�-����}c���Ի13=Y�6���]z�k�A�k�p�m����%�L})̡K��4����J�����~ee�89`�u�q=����ߤe��1��i�[ڧ�y+��>��o���{o&�w����:����qS֏ܯ���O:>_Tڱ�;�v�Z�{wV��.�;s�y�6��ʊE�~�H2*��S��� �S��m��6_��N���<�籷]�(��-wOgt-�~3��*�I;��L�@ѝ�q#U5$��vow�|1$/��)��D���������w���I�S�ю[a�GR���,����&O�����1���C
\��'t��-r��:��ߝ&
�{��ۣ��0����� �5�e9��;�%���I�|��i,T���樭R����	׳����m�������wh�I���ϯ&6���{!Us@,H�bWn�9n�s������q蕮�kU?W�=Sƺ�6[=n�����e%���r��9����T:�T�O����a�Z#���ogG���2����6���ڟ��"��F����=4�.��R�cǾ}�ݭv�5��'��޿V/:�ܠ�b�^/�S��zz���l�ޒ"�\u�#:e&�����*�>�T=[Q^e�PŞ3�2�������{-g�e�-ȓ��r����BfмS���ڱ��<��+���2}�N��͏ǎ_*�����s/{��7�|�W�g�5�W�ѭ�*1
��oE�������4�K��y��n[�9��Ǝ��އ��~��+�ۡK�I�]'�X��Y���S���//w��_�y�f��:���&��[,/ �1���&Ê0���[�)6ЬvT�
�My��������s��{�K{.�l��C�����c�y=�%Y�؎�G�{Z�$��&s��V� �	�j�����-�__]��*����l**��O��iL��A�V>2�,��O����w#��o��j��Ia1�enp�(C�6�F�D����X�f�GcdȓnV������>�*ֽ�5�{[��ӡ�%���{nNٙ^^���Ghz�[��_���,J���>�Y�ө����2�R�Tw�W,��E(b���VS�d���L��
��W��'�>�x���/W�����+w���W�ۢl�
�-w
���?3b���k���s���@�&%�C��D���9�������^�>�z;5�G�e�1İf?pX=6z>��jϰVPU^��"+նj�J�u�]����p���<���۶�� ����J�"��·ٝAvd�D\�`��]7�p���qw�=�D����/�d=n����@��u�ul�[���>b��w ;g1%=��۾�T|~��6�7�<~T�eJ��3�2���=���i��â������9F}�P���C��}��s# ��F�J�ߞ3`�L]��Aԕl0��<�-��3� V�p��������!�}��t�[ͦ��sk.�;��S����7H�33HuJB�*�n�/1yL�x�Ev�j�:-F
�B��<!�����7;�/.�rfIvɳ۴&��EX�:i�)��y�t��!Ԋ�S��N�͇�����u������Q�.�UB��[J{En�*����z���=2Uo��i�f����n�c-Ox9�����7�Y�>��o��ߑo�!R��j�zM����`��~|l%��l��7sܜ�l���,���{]Q�@�\�-�<G��wk�����R]�O}��~�k��rS�}J�,.��5�R�Ky{9
7��Yٝ��q��ឣ�\E�ʊ�/j�k�ԫ�>�W��6U����S�^)���;����:���o����Ͻ Ϣ��@�k��P(H�e��,���s��ӧ��ps�Ux�ا�mz���F��؟w"�����P�l�zk>V��X�VZ����S`X̊�n#�6�MT~�.��J�l��]���'�E�ٝ<�P5�3�9|f��8�ee�9��mb��^�=Q�](Jh�1E�6�{�mg�v����W����ԣz*7}�/��N˔�vN(-�~S�Kz��N�̦l�z6V=�m!1��/7ޢZ�i)>���K#��Dkr���Wb��/�L����Ci7�UO���,v�׃]!�Y��b�M���w˧\���0uM�.?V_���vϯ����^��ޣ��(��;�0�yh��3;w�o�Iы��r�R��	�e�Vb�/`��A{�����/�o��K'z�.�ΚH�[ �)r'�ӣ.V��#��ٸ�z	K{��gS�o
��i���/�xeRg��T���:�lԝ
�f��o��ʇ�og}�܃�o�[��p�u#�T�</�������J���v�ʀ�~�!~ˮ�uU	O>Y�|Ȯ-�W��^�~�/�gmz�48�i��������}[/Y�j�8���%�j�'oa������Ӽ�]���Rng�
Զ�b��ST�.��S4�Þ�Wb����>��{7�]�����&3�3V��J������d'� �*lr�u��M������y==~f��:��V)�r��^�����^���q�ӎY׃�<�-�j���ΒG�s���G�9�u�}�f�۬��!:�=kr���m�t����]Vk�{/9d0э��T�l.�VE��c0�S}�3�m�$�s^0�`�g�븁c^����;k�g�����jM����_{�oR;�v;�ʈ�"����zA�l��^��w5�O6���/���{�5�)�]�(nJ/ފ�5~ݮ)�7nl�R�{��[F#�(��r�z��d�RJ�f��,bH��%�J�t��GUo�v���{�nU���p%@z��]�"{�/݉'���`GZs3�*]�z��S�Y���q�V׫�kk'�g�gL�G��[�ND�p�TT~����I��{���>&����޸�	m5n������d�W���p�����I����rz{v��������V�m�^�dԻ)�C'���ӻI-�r?�Kn�8���z���u0��3�����GӮ�f��H��(	�����Ի餯O#0��{W�#�������U�dL#yn�U�W�|%6~d�mC�g�ߜ��ecʴg��+U���P0�ȇ`5*�g\rp�f�LF�;�:ܷ+�4`y�v�m��L^n0img.m9ut�-�*⮚M�q!��Ii���yٙík��,>;6Ys�Ć�#���u�����e����Z)f��`��I�G{^>t �J��f�ELV�ٕKӓ����7<�Q	���A�m;-���T����u	\j�����ī�Or��~�G�&�E���}u)=y��^�9u�����77+O�)�E��߽�Oj�<�������G<b�(�,�f�h[��o�����eo�>��>�5��-G�'��t��_��O=e�[y��q�����x�H�PU�D�)���2�^�n�t� ���h�)VJ^�8ߥ���zv*>�{s){�@����� W��n�������m�7��rw)q�}Y��I�9�
��=�~��H��ĳ{%0H�	�_� 7����=�H��OP؂�|�Z��+j��/=y�][����#攓����Oۯ|�o�{��Z�h��l{N��#
����&ld�)�/�KثWfz�(���V�^�<��h�����S���'DߠY�͚A�z�&:mQ���<�!{��8>�X����7l< {:�d���y�1Y+ľ��{��Z�*쨼��v�!�zs9��Ry�%�L%	�~�u�ΔމΚ����5���C��2t��b�������*L�Kgj(�*Q#�v�u-Ͻ���y�Qu���nލ�lO�����Q���Y]�>�o�{͙%�C���*�GީtW�땏���GA���^����y�idm��_�6��*Ǉ��2����� +p(�U��u{����d�=��ٴ��c}j�22 #ȈCF�
3�s�۝�ϏRӍN�~��	�'
�;�}���?W��TV��+��͡s�d>�Ǌi��G�WZ�*��\�zE8�瞪+uQ�o�k�`� ���\nx]��o\h��+�b?@R /m���k�)X��k����,��[�##o��,�~�~u��u�X��^8C��Q�@�\�>�{�I,Qi|#}��Vcs�s�j{f���*�\e{���]{f�+�7ϣ�f��U;{�!sCמl�5�z;<7���2��nV�C²فdɾ54�64�b�~���^�uPo"�v8��`'���@����h8_j��n�ڿ����:�ld^�D>�WhL*�T�];ݣwaG���Ԝ$<�w���Uæ.�(�|�yI�7W�}F����,�W���g\��̠ȃv�N�!V�C�b݆�.<l�&2Ձ�3�Q|��7[LL��D;n�έ���J�j`�R��s��sa�3���ge��\l���7�6�:.�򂀼��3Ů%��(���	ޛ�����܏�]w3)�ɐa��ra���bZv�y=N�p��s`�R�z摼��_8i�q��v�H�k�Y�D�@蒕�Ƨm���'fsuF*=�������7�:
�ܬ87	y=��*p�	�0pP3tWi��� ��{�)fP������5�����Ի�c�)�{����s7�!a��ě�F4��s����4n��0"P�;��5��a6��%xMt� ELkD�Z��Q5R�ʹ���/��VooҠ����`���T�ZVɯ��]�cL��NTЖ��i?	�����FΡ-5�,ʌ�yC�Oia�B��ks� e�l�H�f�Z̓t���b�9A�c;
�G/�r�#v�ܼ�Sl�pp�f���m��K��҅0���"�Ǝ;%��e��o�$j�d�Q��p����JӸ��=�%��Ⳣ�fuC�##r������JyL���U._ia�yѓ��q��]{��W{$���֦�T
���;��YX���ۮ�"��m������5/{��2�6�}Evi�Mr����zKb9�f�4�״Y����7-e~���.���E�p����/A�]61���M<.��6��%q��x�+��P��z���8�4N²$e�m�҆�cK��Ur�ѝH7�1�9�/N���˽ӻ�.��gm�:v��0k��]��̅�����Ҝe�g3���:�jÍ;�BU��S��*��H�ty���L�h�l�{ϖCW��7:��yLAׇ�_��}�=aĳ�,0ꚋ�ט����Pr���(VJ;��:9�9q�"�p��z�ɓ�J���*��V7�k,F򶞖dٹ|��=P�_[7B+3�J6Kߵ3$�2����zS6���J����_Y�(ÝWYG����C:�9	�0_nDzje6�݋; g�m��)cm��{x��y�/3N�!�}�^�U��9�]�}+���4!���O{�@337�,뗑"a���v�vvp�DN��9ö�醺-h����JL����rl3��M�:�+-3�w{ŭ�J�<�,��c�>H����٭
;�����:t�%Q���9N9i��ݱWc������
s׭	8t����J�s"�4	[�:�.]X]��a6��U��0x�\+�WV-epȻQ�Ё��OCWһ����Yy��p�bW����/�es}dv�d����ζ+���N����mMav��nn)�`96.䢻,�nE
p��{��Fx�V��l��Q!"K=�(y�Ԉ℁���v�o$�B�G\p�
1(�|��$��|�tIr����}��J�w{��L��g��4�[��}ܿ:W֥h�縪$k5��Sq�wR�Kz=��T���������ӒW*�ʧ̹�
g��.��%W9��$��q�y25�2�#��y¯�V>�W��i9J��p�9��wE󋺺$�u.9SṴ�H)�e'�}[̂�DG.���U��f>{�gp���8�:�9��9���jM*y,����g���ﯓ�����.�"'T�Օ�iJ�{�yP}�.�z�z>}�}2���|:wtr��w&��������]I=ps���;���ȡ躂�%~)9*��C�ܴ�w]�z��rP�"�W�rs34B������s"t�;���=Q�	:�t����v�D25
/s�۞<���{�{���oV޴��&I��0�u��چ��E��]ÅA(� ��L�Ֆ�՟wu�Z�R���ц��/m�E����k��v�6�R�{xѻӜf3�Bt����_��H���N߾���@7����[�ؖϮ}�˺�w�yT�%M�?��.cU�M��)��0�ܿ�I�`�3;��t�=���zi�=�N�q{Qq�ݮ�+��n)�5J�N�;�����V�X�eC&^{oxO�&}J�af�ß���<9k쪟�*�Y�w�D큟O�c�>-?�����e��s=~�R�
u��yM'�l�)�Eju��4�~�#�b�Z ��|�y_=�/^	ʥ��Ge����>dFC��.p"��(}��U���Uk~c0&G���
���R����뭳E��`�H8c�'k��)U�s�&���h���Uo��Gܬ�)J�b����@�ߞz�����������Ű4�Pв�e�U�nT�9h>�a��.20
쾃>��}?C"c5SEdleV��G;���Aq�Q�7�[s����cx���T]}I������8��<�L;�,��}��y���#��o�9��!�C����&�t܁se��{}a���!Nk�,�7(���W{R��5՘o���6�P׎�
N���W�?��Lh�"���*��I�}8j��j}f���&��hyT͑��;y{��=V)7�pJUr�F�L�kٹ�Y3	�C���jA��|)�1�*��b�y�[��8�e{����\�i�t���F䩇�eJ�}-YT6��>��/�:4�U�{+�!CzwY]��u�����lq�x�w����f�,:�c�z7��L�����Rܼ��	�Q�l11C�ˣ�x�=/6/�g��zM��6o���݇Z��m��Q-;�d��z��AX���F֓�o�0]�eB�ד>��}ހm�N��Fv|��*ka��h��tj�	��C���AMaaW��I�؛�1?n�|R�ڰ��c�Hf�N��D�Kr9V`<N���	�|k˅��a!�Z���{]f���a����K"�&�q��kexq���u�����0�L(`5J�nœ�fd\3Ne�{pCs�5(���*^���i����ɏ���j��%���`��?<�B�r����/�hnz3?8'��^m�'+Ɠ�K/�K���Sy��>��ŕW��7j��B�`��k�<dwTp;��%���O�Q\�b��)ϼ)�ڝ�0�[��H\mꋨ�>I˖7���CT���)a�	��\�M�*�'�@�Y"#�O��S��s�do{[����W׹�^��r�S�"z���Jm�OQ�%�0�L`�zuŬ����ų���c�z��Ӑ���	�q�_I/Z��9��B�[7cjYc�]����Ɂh�w]��o4'j(ʌ�J���N\���w#�D�w��]Z86K͢��3�Â�o3��2d%�p�U�g@��Z�y���c�s/y47�A �I"�g?owGY~¾��� ��a�~�p@�Z���p��-5ղ�����d�,��&��s��}7���8O=���R���(C��\�`w��_qe��SA�y��7���oz�K���c5�R�)3>ɨ=#W��Ps�}��
J��3Q����5'���y.�K��;O����(����܉�	aX�^.��H�9��/<�g�/�\v^fØ��֣.���E@/��Aƭ��QM�w����&�*X��b��1	{��P�w��E�鬼ʎ�Fo�_��#|����0�P1�t8��!�T�fF*A8���t3��[��t��=�is<�*8PŇ=��_�[��z�N�)ȧ-H���d�\:��U[v��}�}�=a)�pF������"<�xۘzGiP:�a ��]���׸>�z^���}Z��=Wg�m�Ǜ��إ��t�!'����N�K)��	�]C2	���v����H(�=O�W��|����D�5[�֧6F`���g��,���Lx|ăCϔ�˟@�6����ry��{<5�nX��;�ݸ4��߄��X�5��
A��XS ��$��12JQNq��0U�j�2J�>��u+���)�;�`cw�ɷG�� ��=j�u4l�P4.��6��,b�}��f�1���f�>ۥ]A�Z�6��3g=���_���Ā��� �X�w�;�'�GƩ�xM��Ct��T,c�}W�PV�%��$�@����Ծ����t�+�n��oil��M��8��'����~�^2��YR�n'���(�;��U��۲Z;�b��4N��߼qJ&�ZM�A�vN}�LC/�Am�������=j�}~��뤪y��J�џ��}0u��u�Qѳ�[�g�Xp�� �+�S��dTu��׸�L�V��y�j�)3`R��_},�����1����oy�A�y�p��=��!i�q�s�V�%�^�ޟ?�m@p~����~����~RԼ�;ʝw�c4r��q�}k�xm��"X��Q�}��{ �2<�c޻�}ম���0�	��=G�̺s��c�M��=������B˦�z�j��5`����F���~�S��Eˁ�����:�2���eA��R$���X��z�ޞ�*�r�5�5���#����)G���Eo�)m��|��\����Br�!��U=ȹ�s�RQ��~��󼷮
8���|U�g�&'�l=�yz�_$ʹ#wH���&l�WV�utV�LiY&��Y������;P �87'&��Mj������W�~�y�����2`o�5;t6.D:��)��@.
gvP�+Ff�)_dL�f�u�9˰�Ύ����	���f�7 �lrq�_3;an����k��2����m<��$$̈́�����}�7�kD���4_ғ(/�w8C�6�_T����4ٍx8��v�.�әE���cd�W�O�k^������B�9�H[��(`�	��P�k� �tw~��g��|:�P�xeJƫenn/D^��+н�f�E�l،2ە�z65�85Aua�T:�^Ԫ��ܨ�w��#w.���������Dm�ZS��F��P�^k�F�y:deGa��'�^q=���`�`k�-���~2�|WO�f��4�B[��IJ��Hc�}�Q��g�L�N��x�N.a�c��-����éŃu����� �Qq�ݮ�+�[��xCR��f%�Rͳv�;"�l��i�+��R�Na�AN(>0�5����e]��ӹTc�|و�V�2�P"�9��x�yx=�+�Ef{h*͗ʱU��q	W�]�.���i�Q�dwSE���ޞn��;����^�Aн��pF5sʛ�c�N�ה�)����.�g��鋰ؒ�4-nUz��l8ʏq��T��4G�Wm��(99U�s�&�æ������Er�IT~�XX๘�B녚�Sy!H��U'}����"f+˽�C���}H��n�g5�4�nî�8S���.wb��F�kK�����ɩ���u8;Lw��=|]p���d���s��cXzK�Q���8��G`��:�n6���Z�,�1��;�v7��?�UW��vԑ��y�|�"c�}"��a���q?.��NS}`�!4\dev_A�}YR�pߴ��s��=�%|ǆTA�AܐxC��0�z�H޷m�|Qr���==��.�2&�,��u{0�]���[��C������ܵ�`9#.<gU0��s��P��w����!:o��`�z/}�W�J�^�g�$��p���?��#�Zap�{�D�����]�5�jɣ�C�W>��8���_t�ܱ�u%:���9�41��c��b�G�l�������FO�e�'��t���F����^���Zr�<լ��]�H��x�d�F�����|+�'������\$��8�li=�����휹��c͑��8�}�����F�ᑫ(&�	�rl���r��	y1[��:
��0i��k�:�[/�.[m�Iʳ��tT ~s�%Ü]^�M'x�u�v�wx�d;�����L ��Y�����C}�#��[�\[t\� ��8\��0��1�AuR-	>��-?k+�!���1o��S�^��SZ�r��'�H}�;�3�픡�k���3QK5P�[��0
5�n?�Ny[��?-�EG�9Rj��^VR�A�8ڶY�*Mև@�8\4�*0`�;�����t	˺ӒէWE�A[N�K�v��@��#:�)���sk:���u�ئ���|��2���x���}����o�ٞП������nØj^5�\���~�)'��$b;�}��Us�t��Ў92�m�sw�)�q���U�؇<� ��bO����s�s'�����Y[�V^Ϸ]���2)����_�����G,���{��;��0���\2�;UvO��ʔ~B#s�|���ʻ��ɯc���Բ��G�Pi��/G��S�3��?JSnZz�/ d�{��93�9B�p��دi̛��5���xY��	�0��ȿB8#=p�\{�k�t�	�1٩�o���M�ߟ��=J�G:�,7ʋ�=lnF���!!���#����fOO�Q�D�u���V��R��|�Yc �`�?r�Bϩ^)3>���CG�0��&s��)+h\?�T�6����f�a�W���$��0Q��9�{Wy���x�\�Dℰ�^/>�(Gt�a��Y/x�lM��wQ`fο{Ҡ���b4��'j���ȃɤK�b������,��}2����o#P�JH�EK�p�Y�[#1&T1��;�Y��"vNH�{QZ���cwk��r����)�c�xp,حJ���R�Y}J�2��-��u���Y/3����A$��)a����DCs.ڬVSM!G�1H���6���u�l�ټ�+�`����YZ����L��h]Y����0�g�"�f�ޭ%}vd̠V�����j��r5m��� �ðVtÌ}=#���=��y�{#�)�}8�%9n�B"/|7DVڅk��0X:�
T�m�  �ؕ�H�]����z���0����9�;-�0Gs�p�SN�!�\Ŧ�n:]_r����b�k��:%�,��z���d���"���!��:�wګn��f��	�B��UQ�V�qEj��	?r�"��R��G��]�r-Ǩ���#��T嗝��/^����bg��?wXHIn�m+���Y�^My��w�� �QH������j'��ݘ2����Mf�Gl�O�lMA�L9)�W�˗�YR��m�dە޻���a�m�?�������0-��z�J&�
_i7w;�<��x͋z+dO��.ߖX\fY�S�y_��0����%`\|||6އ���h'�Z.b:�b�{>	Xp��ik��z!�������67�p�.=r*�dzԳyM'0%QEƍz0!��8���m{���"���犩߹q]Rt?A}5���B4�4��2i����د��H����(׼����s��[��r���(���\������	
�坔�s����u`Cnv�]��P�iEG3�z��S�S��a9G���.z�f�-�vԳF���,a2��t�`�+�2��#wj�"v�ґ�+#��YV��3z���vI�/��N�P*f"��o�3 g�U	�f懇<,|��m]�/�M\7/��0�V�t��A]��Z� �������~�v|�s=�r��w��#��
Z�]M���p9�5,l�%�j��	�>j<�-�. �]�d�YC|y�<��|��d�㳻�
ťԂ��{c���:P��U=��?�Z�o
z.m.Z�-��5�%8��l�
����.^#~����i��s!������c�eb�j���;v(ެ�ZK�\ծ+�T�v�p����6�v�P�S�i��q*2|흁݊������f�vgo{�Z�K�����A~ˈ�ע�l
1�v���\W�7����~^�k���op�i��.5Ү�݆�Rٱw%��נQ����\Mh���yP9�yJo<L�6�w�K^�����Փw ��3�ڲ�S�hR3K�����h�
`��c��Wj�SE|�n�s��p���,S(�O��[�ߒ"���Е6$�i]G����_zR�� :;���VL�݆�:�f�JY�u����Y���Qq�Gv�G����|�2��x=��&@��8t�@�	����Mϋ[TA�� ���R�70r-�ݣ�|M�T,p�^ �$ۼ\H�������/�M�M]�����+�%['�aP���]&�kV3rP* j���b�4��|)V��]�7�n�|�ϟ<��T�}U�W�ܖ�ʟX�~;��4�W���˕��6�~0&=��i�hŞw����m^o��'�b���M�U���]^��7אݹ
}q\�bS�� JO��j�G������xjm�qEd�^ȕ�S��oM�s��p��g+b���ϙW�
��NE�,�k���2=f�#�:|�f����_���W��?OSA��{��=B;g�%t����Ie���O!׮`����ءHƱUjb�EҀ��E�,���'�ܷ>�*�r��������/���������+�.���[��q�M`��M��`=#n�N��x���*��?|#�������H��e]��n�=̍hz���>U�,l���Bc�q����=ջ}c|�r�;y{ي*���Z>[>��2�B�����?f���C�n@YC���9��u��X۫�Ӄ���P�+S�Y�ګ^���:�k�ս5`��R@�]�~s霎 k�G�GCl���<�k���P�3�򵰝�×*�޿��ŷ�=��a�̎妇�ciDs��b	���Dݢ����B[�-��k�}>4!�)	��?ÜX�^aޚ���)�d��&�ufERR���[�_�F3졷G,Grf���=r�n]M1,j�VsqX"�]�$�9��Nč�v�M���=[���:.����ݺuA.��Γ'ۨ�+x�)&`�v⽩�!�{����F_oo�3����(Io���Y����vս�]Т�����n]���oc���f��u�	�8��D��"���cc9���8޷��]�l^5Չmt�V���nƻΰ���ed�n ����ր�r�2�����b�u+�1O�����7��C����Y3i�X��k2rÃ:r�y��f�����n��TTv�ofG�jܙ�ܷzZZE�1�d\�%<��5�=���D�j�ڸ!b�n��},����q˘��0;q,2�Y+���V-m��)S�ý�����m��z�a<�54��6������y.���Q�c��v��E������F�y].��D�Ѫ��q�P^��\�#���y/Tk�%���ˍ趎cӶ@��ӭ�?�ESbճ.L�m�r��\��Ұ��ja~�3��[Slf���³��_��Z*F)sg��WD���{���(u��i��6!3�%ζg:����u��U����-����e;.�EX5�4�M�o�c�������fS�+��t�)*.nZ!�2����Xh��.us	�	ֆ�f��Z	��r�O�^Hz�̢�O65.��'�أ;k�����q�k)Z��
�H2�1��Y��[<��WI~�l1O �9P�:�}�ttW	ڝY�+ntoDZ��T�kv�5+8.�-N1�:Z65���7��������C��'��fź��t: ���ᇎ17��-|�	=�T��0�V�޼c
�Wy-�k�|I�D����F�yV^�95�D]]Ųe�Fw;��:���dB�C��ڋuvZM@�8��s/9��W��=B�jk/>u"U<���I�@J��An^ڼw����Awwn�$�h��AE�n��"F���Jt�|'4/��Ǌ�[ifm��w�d/euz���xʵ�!w�i� �a���fS�n����w���dַ��b�YFlm�϶.)=������o�
����29u��,h������47�˔�'}�-&˥9�fa��e^��� 
G�G�s�oM���ӽ{�9����%	��k-љ(����ڲV.�$�rv%D�g!$�i��uktШ5gPY�{�
G�V�����.m�:c�����0�^����JJ.�z�J͙G]o����2v��,�qVk�ư����EM��#{"���]��#���iTn,69"{�$Em�hԾݬ�J�
��G[&<�`Ng1�����E�ݕ��u�����ڲS��j��#_+SӬ�dPv^LM�|�k��{�@�7Z1��mV�)���tC���	��$pJ΄N�� �I:QQ*�i�g���i��KV��:�lZ�Y��w
.%��9�*etQE	"�Y!��=(�*'���K}�	�	�=��0�=G9E��MSP��8\�֩uKQ\�"?<z�K
�
�\�BQ5C2P:j2�"������*��{'9�&Tz�E�rEjf��J��B)�t�fAVm@�29Z�QR�I�E���E�*j�QQ}<�i��ʨ�54�­L�6G6�Z+�_2��Q��dQ""P�.�X�Ȏ�UE��(jR�W*�,2P���u�R�#e�B��a��D�qv�fV^���P̿G��=�ȟtgs5
�� Z���./+��X�J�Uiu�$ֽүS��+T�+���=����ܖjUY$��n��Z}B-{���F�$�h�i:dE�!D�0̜�}|���ts��!�eD��G�(!mjbj�EXe	$�jD/��X�[�g)�i/D���w-�*��������������Y��&�&w�,�q�t�=�s4����_��O���z���],����ة���1&Wd\�O�f S�)ؽ˽�R��[����r#V�q
ka��]�Tz�{l���{���xoGy�{3�h�:���OG�N��;ڬOpZ[��*����	�P��b���Ϣ�Q�g51��'�PH8���.��|��ko&Cy�Dt�[�\[t\��_ΟP�WX<���ޜE�=���GXz�8������2Ƌ|eJ������}��f^j��ʌ��T�]�y��[�"�׮`���0dv�9�KƹKb�O�.��<5�@��Cܳ�O�����D�uW��œ����Q��I�1��&�bH���8��@�'j��gG@�5�!]�o��`G���Ӑ;��sϯh��L9��*a��.M�!Wd��eJ�Nw��o��hG����CA�~���4\���pk��L�1Ӂ*.^|�^2\b�(�o+�~�>� �.���khxS>?�?�7F?y܈���q�!c��T���8W�Ã)f���vY���K^~�^�a��;�;-p4?�=�
���z�s��@��`=îX�Ԭ��wS��B3OG������}�E�L4\���oCٗ����c)]l��pͮ��k�����w3tP8u�,�I@kp�MUv��� �7x1�k�ƴ�YI�f��nҮ*�K� �aȞm0u�Vj�f��=���"(]sHmT���}�?���}_T�um��K�ח�c�6����|�X�V�	z��c�8p^4֎Y904j�g�Ϯ��(�O���}�T�1��<��X^6����5,)�4<�]g��z'���r��z��dk�����/�*{�b���o����-�ލ;�p�_'H�l�+�ળ/�3Ԫ}�����2�(�qgq>(ŻwUZ��&T�>��y�g`XS�N�1+z�j�(l�z_%�8�"]ȁĨV	Q�!K����F���{#�u=�N���ë��+�V��.͘6}�}6�$N�{<ܨ%������C���{��{s{m@�子�a~��d��j�L�k�ֲ�_)���7
}C�����A�|�cC�-��>��f��E�����Ss��'�w՛^"Gsƣ;�Nڜ؇06���lqEj�P�|¡w���㓵qƮh՟5�r�����Q��� P���#��BKt�i]E�
�g��jB#���T�*w�O�I�y�����	��"�7�s�5�9;i��lMA��'�����,}O�\m�-z��}��,�S�m1K�Z��n���)�\֙��fi���5�i;�nN/3���Kl��fi�>T��g�~�q׹�~pT|��{�j�1��A@�4�
U�勗���]�5�'�Y���b0^WV0�?��Q�ʾ��ݭ2��p[x��	u�����`>{s��m��ˬu����>
9W�eK�}��Ǉs��|��k[N!������g�{���˥"X�~"\t���tS��8`��dbr47�O���e�#��
�6�F�z��L���X~ͺ�\�I�a����U��aH��"�+ܱ�G;�^J�^f{��+]�½B��++pi��+��)kW����6�"��]�{���35�f��CF�ؑ���~�nZ��jPٸM4\=G�F�>�;��i���vnԲ8�u^��'�k�#�رl�S}�.\�m�~:�2��G�#*�y=^�|�Үsu{��0AQq�ܟ��8�� �Z]H+���.vN�+��Aezg7si�>���p�ǅ!'�p�v� �����r�K�ߠ(Z�`��O"�h����'R�9����'-�����T��!��t��P�f5�ڃý���Ńt�U<��=޺֠<{}Ӊ�@N\�n4�����B��0c����TF�(e,�>1����x�/�$�Qr�At9�հgkR��2T :}���c�/�b���� _���ڑt�z�������t���N�Tǌe��-�1	��:H�la��㷃�=�;�\�Y:���p�Jޠ��&��)����꯾�7�5�ߑ��c_���;e�����W���+��
�~�0O�\���韘�d��=����څΣ����VH��M�z;ViL�iC=x��m���FPtw)/VGY>��oP`,��}�{R搼G��D��VD�Km"!X��I	SbHN(1m#P��{{#.��V�fNZ	.�G�w��x��Q����k����CԢ���npq����E�Gv����n�E��/����_[�\��
ܞh(/%�Ô�ΖU�|<�j�L��
��r��,��=��a�+]�Vz�<�:�J���ߨ�Q�5�*��/����$�,��)�d���N��==د�*���ɝ��\�����k��4�����p_��8W�]Y�?Ui��;!�^B�}��|�v��n��(�v��02��v�?���^g��V��<����j�<���������0������I��]��zg�KF�6��M�]���޵�D�[���U[��>�a��.2*� ���[�潫��^a�(�9�ysӬ�9�8�&�>�r�1��ۢ�u!�Yn}�.S����~��������I4t.闔�uI-��۷�+C�щ��:@0�p�:pe�]����ͦ����@���)���2<��������ӽ��~�FZ��BqjDƛ�T�NJ=�j�E6nr?[��KL��_.J���:-Pݱye]��B�
���X�8�{�f`�b�dV��З����s�i��j��ep�=�Ã���?���r[.<gV�;�n��D�cf�]��]�m�m��͖��A@Rݚ���7dQ�x��#�:шCZs؞�s�~���%.p����>��ҟ�=��6F;���wI}3��U$_=(���}?���>70�nzg�ݯs]��OkH*{6"�����۔}��*5���l��kzH��rD/��6s����_;}�ir8PU��Ř��QӾ�`������;�]���=)���X�5Rzc�WY>׾`�s��!��B�(�S��'MC�=������!c�fN(=C�Q��VN����n�FV����A �br���Eǆ�ŏY���8��oq�-�./�{g�&���b��L=��8�ʕH��V)#�����$�x ������T����a�_j��U-J�5=���
����ш�������WQc'юOM��;`��)���y��n�L��x��"������y%�r��s�}ʛ1K�O-�!5{G���z�D���2�ޯZ)������(y��� �ukr+��7Fg�9E_V>�ޡ�����.��y�!�k��=�ڇ0ZȎ��͉:�s�;���uU�E����X��]�/W��Ǜ��Ic�Y�Nٵ��Jo���Z�jkP�4�ðoׇ'
zS���)�j/#�  $U�l�l=��h�ٿ�����:By{G �Sv0ySK��SGbHU�>��w�*j�*���1O]y��%xh�A��.�UA��pk�ԙ�b�)�-��Ϫs��I_'	��Ι~�E_Ѝ>�}��TS�ů�`��S��˄to�N��͘�ʪ�݊��{��M{zq��+�:w��{��z/��,�B�n��6��ۘ��J�
��f`ܬW��=��~�󨽿_�XSA�c�[�O�)^|�%��h����_.;���1K��{;�u�4l���\q����m�דڻ��a��@�܉�	aX�4|p�����Ѿ~��8��H`亝�%�=+�b�����Ym��v�ۗ#�H���C{�i���^�uٙ���q�ws�B�]{>�[Z�$�@/ka[���v���Qu�7ӂٟ{p�мz� ��XVrVpÍ~(�6:4����?��������t@M��SW5S.����!�NC��O��`�2�	l6�@A�bP�/�/r�h��z{J��ҙ�����%u�icR:w̤�eH⛋�)r>�oR��Fo���!�=����H�[�᣸�q<z��6�^�����r�gM1.u4+��Jƒsy����}m<��-��CsM��];bo �t��"1�yk�� q�S��}U��yr��:��/C�|�&�w:1y�0t�c��A[1����
[K���s��q~Gt��뺿-���*#��u�u��*J�LKn�;jFlC��Ge����I�k�ȏf�|Mґ�&l7��۞L�����ױ˺�z�	��		nB�WQk���'I����&YV��B�/F}��3�������L��
�z����\7_�2+_�)���챓qov�X	ʲ���4�9�ʟF'�z�)ȱ���){�e�bϴ����A��T�<f:��s3c�*�O�oDj�{��@޿@���^�tS�~8f�3#�����{�+�na��Jڬ��+ި:�s�t&4As���3�����Q`�D�0�"ÑhO�]�{��u_<t�j=�L�h�m�"R�(�r�;PKN�����-?.ߞ�(!�K�=�w�/��i	��]6H��(p��?X�n_���n_���M[��z�H#��4�����gY��&�����у& �����4�"ŋd/Sc�Eˁ��n:�7�u>�_����>5u<����0�gk%mض�,Ti�RP�`�S�-��2�i����n�'S`�ډjU�N��������GIs��z��#"��-=U/����ϋ��ꃚ�-���5�v�t�͔"�|9m+1�{T�S_0��;R��'$f��/�>:VNK��`���Nݍx���&~>�$���AIq�ܟj�J8�6"�V|�R	���)>u�T2^=��8j����F_p��.��s�<C��m¸b��\l�|g$\�R��@Q�j�2�9��c�:����&����Wt������T䉠;hH��t�O�!����<�yWG q���m-C|]�F��Ӱ.�Ӊ�S�8[�?e�qU�%* �Bh1\���'����h>�Z��w����F�;���>2�[.��ѝ���{<��5v\B*�DµB"{VOU"�t��x���Ȧ%�
�
�<��T�.ud��&�=�4�}
�K�����Mu��K3�jN���y��:�3W3_h��B|�z�ߔ��^�m+���R~J�BqA�����4����×[�x^g���J5��
c��xz�Y��nz��ڋ��;��sl�����������9��E{EfGu��\���)9�PS��7~0��R�L�N^�<���z�u}�yE;�|�u���h?^@PSZD��s�4���,�� 7ޮ�~���D��շ�����:�1b9anS4f��|���zˡ��~��ʻ��9~�9J�q���}sHbzt�W���,=���)Ttj��ގ[fg�+���3D�8nA�ܕ�jr�����F�;=&&u�y��]���,E:�.b��(���ճ�hm��0=�}�z��nx�>_,|h��1e����-Ǳ+b����ʽ�WVzNIɥ9��<��PLtX��w���B���W���{=A���A���9U�s��0��h�ɝ���d��l�cr����܎ұu*J-7�x�O����ދ�B~�Z�"z��s�Un^>�a�G�l���i~~�U'fw2������6;'�ч�nnc�Du��s�ynۘ�pD�l���7���e��`��0���Q�e~=�c�q�o�q���Ng����s6�/3;̼��P�U�ے9V9�PJP|����
��XX��m G>u�����룼�<�<�-�f7e�9f7�=���C��S��^J�j��c�Dp�7ے��]��-����AfK����$-]��Z>���nTg���x]�A����17�k���C�pD�̏.��?z�hW���yd#��"���#%�=��5�����yfmy�����`����g��<�p���s�U��>��>��̑r�.��m�	�U�Q���&VXDgwE�X�[��+8��[�{��"S�Ev`kQ��++���r Ge��7b<�v�̈��P�m�m��k�XѲ��RY�z�lӣׯA��So��'JS��.n���4��P�^��]qF+�Lr�M��u�kɳL@���i�@	�I/�����U{�{�;4f��F�w�p�,��j��|NU�������[�	�wS��޺�E��K�5�D�.���y�׎a��q�W�	���\]'��$ǂ��ӏ�M�1l@��l��:��F�ת�����fF�=�'���nØ��\�R}��"��0|�����W.P�8G���a���rじ�{g���^�>��M���;���?������+�z!	�{�(!�z��=N�_�Uz'�N�n�@~'Ho>���{��;<��/�*���ezd>��MX7).��,ϫ�zu��7��.yx�|�ɧ�b�-�������,ן���L�6�������(o���p�~�Ʋ������k�!�r8/Ў�㇃�/E�G8��·:�o�"��G�����^��t��OqD@�=�a��� hu���}�"��a��Һ�zK���`~����V�E�Q���C��u����QS���L��~	OI쭞��t�*+=ݹOç��:K����E���'�����u��N.�r'%�b�d������}=[�Z�OkK��B��3:�@!�ku���gSb���f��=yW�ܳ�ٖL��;ӷl��f�zv�T������M��v�F������ �� F�8o{�����lp��⴫�S9�4ָ�>�yW�vY�:��
ՙG$�d�Ù���;R{��ii�f,�A���8�w�:�;էq.&X����b��l7�\���rf�,�n�حv�Dy�1��E�0Uĭ={�ݽ���\�Wa�,6��-��M�Tt�=l�|%\�m��D��y�0M-=q᝸,.��v�S��5!A٠�b��0:��M4�^�|K�v�8�0!�L�nomP�~}p� �dx(al�(�X��{��vC�\ C2n[i�޾N]K�G�o�ǵώEvc��8��Mm�
5[�
�}��E�2�r�-�gv��v��|�ᦋ�w�y6��0��)8	+��MF����#51>�WBv�޶�1�',5��jv-��K�<�WKdV$h�ulb�����&]l�YZF7��Xb��=x�>*J�(-(�Vb��N��z:U�ǭVC���	�k��[w���8�*P�T�-���R�j�k-������z���b�����sp�J=��&ͶK˘���8�QY(�viE�wt�p湝,�K9Eb�@�2�2�7���W�0ǨfZ*�:wEGG]>V��e�ɜ��gckD�fkx�%�����sK]�⭸��YYy��aY��m�X��+Ν�S����1�VR�cU�ެ���$��u��c��r�^�Pۣeҡ�a��\�Yu�>T����%Z�Eq�K�騺�z�S�sc6Ƅ&$�KОr(�%��Ӷ_1t��0��!�0]+�9z��g��B!��g>	bz9��ޮf����zL�h�vw�wG7tP�ܠ�Tj��.G�8eG�騜�z/��ӣk3F:�<����m_i)��/7MQ�t�MY�z��
Bf�:��_�N�l�l:B�k�2���^Uj��m9rP�Ğ��eP̅v�g@�������PX}iԺx�h4��Io]o�V�_��ZӍ�و���6��кg�+�nkxX9՗nU��f�s������@Gp{�Ťy�:n�_kY���M�oiЫ��k��͍u�P��0��������ڕ�����"g�k|�vF	�g�G4w��orW�܍�Аꈂ��67˒��շ�S��V�93�is�vy䒏�,/�Q[{]:�;��,�%�S���A�ME�UK�V�n��Z�Z�r5���M�g�)�����X�"=�@�7�3V��.�u�G4�u��;YM��YL˾�*:vl�Y������x�h&є�]�<�C�_E���a�v�^kT�7��1V�z�䚚���h��O��b�u�@��j﫶kx��诋�&Lf�j���T�y���v͝
NiCI�E7������Y:/X+�n$y#�vw
8$�(^��H�a��quT�&�����UTT��t� ������"��^�CZ��=k� tU9r9�$Y�p����~���&G%^|������P������w��򾙋�w�z�f`jS�州�o#��qGu�yT}}�o����u����I��<��U�}�n���оC�n�~�rz*��~I��!�;�=s܇ʑעy!z/uˑ=]��g�� ����zm<ڎxTjU=Ǹ�U:�����ܾ��q{���(�^���{����e4�����uY�z.�u炽�ė�Y�F!b�TYyo{�޽�΅^�p����3,Z����ЯM�z�<ÞNl��'����p���׺=O9��Qc�*{��t#�G@�H9\����qϝ��{��9�W{Ǖ�3��>������EǓ�r"�{����6���GVU�����ϾN8�[��x��=o	"��w��{�#�OSwt�=�Pד��z����/{۹*�x��t��:���uJꕆ��ڨ7jP��QWx���4a5u)���_��x��Q��3KQ��9ϛ�O{F#md))���s'�f��̭��Ͳ����C�6*xBrG.R��kB�����Ym��N�"֚�#/}u}ssw	`묿u��$OF:����x�;�9�FK�Kϑ����$ʀ@����B�U�<s�RF]yf�$p�B�#� �Z�g ��C��L7��'��:�u�����%�L�ɫ��\��]k�,e��B9�P��B0鐖�pB��Jck��	��0�l�$?F�YQT�{x�p=g���9�;/����f�A}C����V���
���N�������kh�w���x.9w���?m�t������;jYf��06���Q�67>�R��y���R�����0�'ޗ�EO�f߯a���P�]�܆!���𬇉���뻩�Mﲤ�o{ox?>L� NA�pw��'���wߺ����wi�5�TÒ�i�^��f�ɫ�I��C��A��eO�C
�"�����k����q�{��Ҳ(������gWE��<|lZa"�D����.�J;F&���~J ���w�O��eř;z�u���ˬ�������I�J��xݕ�W)V��a|^pѶ�-bt�o���cL����:�乞��'gۢ[l��'n.=s+�k�\�>K�+�X3�σ���]E��U��n�=�H�;�cJG�:��}��s�t���US�������O�L��g�3`q����w�*�r=j|�����s�W����'�J��*�g��w'R[׌n�3��!�WF�1n|�����@q-;r�'vw�NNO�K��� �TQ݌I�o4M�g��`�tP��=�љܻڞ�~����.�zCT��7����==�{�Δ��@XU�PIiElX�B�}�䏖�s�9�j_�ubH�Bq��b��M������u�Zd$�AI}���>㓓���H)m��k�Λ�ғ^���fʣm����T{-����Xe�A8�p�v�b0ρ������ُ��ΓWz��U_{��Q�c_�r~�]��dwI~qX�U ��8��F���ֱL�2�����8�3;����{_�Q�Ν����p'IM}�9�n���8��
9��������Wk*_�w���X���)��zw�F ����7[��k5��ʂvu�v����Wtp*eJ�KǨM+Tة��t��P����q��Քڝ�B��.6�f����������Mu��IOFmV(3�ţ3Zq�On[Of-�⍖���Y��Z9`[%�RjcG^��a�r򘎅��A���M_
H�{m6f�[�a}��G�ZJys.�:�D��=ܝ�����=�͂;�������h�oY(I�',>fD�E� `��U{_�r�B�>i��:9^v���kڄ�|�Í{��|�������M��d�Fmh���O�*b��v3P�A��j�Ozj'�ǩE����͜^�<j�h��t5�rVT��_�w���/��`2��T�D���o&��������ç�_�WDgTpH���J|�>��d�3n���1�y[ߨ�Q�&����s�zNM>�s9�#!�=	��\Oe�Z��{��-���m��F}|v<�~��Ÿ���p~~V\�U����~�94�(�bȳ�8��K����6�ixZ�,<�1v9��m8W��?OSAJ��MY��[e�_���*�]�ٷ�*��1��:�U%I�Va���� �F�M5�n[�*�r�g{F�{<���\0���<�.�x�_�xѦ|��!y��■�5����NKd��6��7�΄TKb�2D��ʻy��� �KTz[���T���w_ڏ�+�!�8;��3��w}��/3��G<i���woE'�?},kWP�.:���;�~̈́��Sc��7 ,�_�l9��1n������=S71Щb:�X+ɉ�O/�񻶙򧀼6���o.��ͤ�Jp*ݢ^.��/jh�kr��2'~������ݫd]�U�mL�5l�u݋K5��W!���;�nj-d��!-g���%;(>��5�+�v,LΖܖUb�G���{�` *��]^�T|��>4��ޜ��Y���z3�jl�v6I	�t��g#�Tfb��&��J�9$�{�lȖ�@�Sb�6W$���0��}��ܴ׻cKQ��o6�A>��7~/R�Vp|쬽�U�H��A�഍uSF�j�2\�f����FH��z�7nCe3um����{����We�.����hm�豨���S���|�����P[_�JR���+��n��;V��2�N��\�fd�<�X)q���A�')�>X���*{W�:���T�y��@�V�jrww\\��ϵ��n�����8��*����R������X�o��|� �̚��,՝ם����޺��+v�~*ɹ̍�g�(�2ݻh��/0��d\
K=��އ�<���3k�Q���߸>!��(�k=��Ct���o��z�#��Z�lA��I��C��4*P��4�{No�f��Z�T��h���O�S8����!�ٳ��g�T×�LU���wuY����BT��sS�/B�W����0k��A�W�2���E�2�~�3��?H}9��5��X�'|g�����)��-�KV��	�T��˘ޥ��F�Μ�<��l|����]8AvÇ� ���U�/f@�]��;����K�Id䬆�<��mƬͲD�ak�\�2˚hP��Eǲl7�e��-lY,V8k��bϾ�ꯀ������[ߝ���X���%�0CܿE~N��xS��ǟЛ���nDx*�ں���Ϭ�_6��{��/�a���zT�9|�#|�NFg¶���dS u�>���+�0ؑ�\���٪v�A���q�c:�8E��u�Yp��p�}`�)�!J��Dϲj��Fo��x]k������s���ؘ�Ӎ���.^f���ۓ��!�~�C�����Y��O��_,�o>�e~��X_;Tk�wI�EIH��X����}7b�no>N�+����,�G����^{�F�:��S�K����^9,9�4�/97��Fj�^�u&T=t��D�Q�xw������ƠX|9Z	�@��O@!Y�;���	�k*ݲ��O���9�u����ӷ�)�Rb����`�:d%��,ġ��8^��:�6D
�y��5W��ua.c5�s�c�я��N:���'s�L�(} �ߔ��V�T�eȃo����Y�*��ߙ���j���3q	K��@)U���W�H�wQkEd":�D��@���)�v OM&sޘ���T:�����(�(�R}��e�E#p�Y&ʆ+\i��Q���ʩlc=r=�s�S/6�NVi�]��Uv��):�.��Nٵ&��䚟:@;x8���_'y�Y�+���LNA]�,�fa`���Y��窡o�1}}p}2��L��V����'��A���)zdͩ��^�^� W�X��u��t�+���S�ң�ۋ4��O+ٿ%H{�~�-3��	C�]��b�`߼[�Y�����O۴ؚ�RÒ��-���pr�t�g��u����yK������O��a{�L��/m��=�h0=�g/�եP����'����3����< �l��$o_�^][6�W�Ƈ�>�:��<���ݻ�Tz�}�q��7+�P��H[�bV3�\�+�f.�l�='&���LS
��K��e�{�!��{�ףּ�m��Z~?p��}y�p�)�r�;P��Fg�����列��kL�S�D��3���`~��z�Y�x:9e4`�l��]�/�M\7/�:� �M?w�.�H�}��u��b��~^��P�Z\���(��P��lX�~���]�\���RϗO�����ث��;�˄��c}.v@��Ze�Ӡ���O�>㓓a�+|AKmԋ�z�����J���o_\����q�҄��OC�R%�'n68!q��=��x�ŷ�+:d�Q�wzRh�����>���=�-�E].���ZyBW�f.��0j�.w����ߌ��x�`QDY^U�R6���=D�!���,��iV�X�e�!�r��Ssḁt��Ҝ\�w*��I��Y�'"���$��oV��=*#'"r@�� ����us��7"��ѝްu+��1�t��c�^H;)NH�nq���lM�/Wc�[���^�kf��a:u�s�K����,��=��:Jr�ŻPC�\G)0%{�bM{v�W�̟(�����H/��@���~x��I�yS�	9�3�W�����e�!�<s�����ޜ�eo{��&4 �����E�j��<�X]�&�g��f�ϡX�.6�'4�M���B��g�,�2�����B�𖃤N�~�ϔ�q�t���Hn�@u'.,���s��Y5{���m���Ǉ}�g゗��5��)�?�3��?�������꿢�U�4�^��!�(ܲs����&����?�l��H�#�5�P��R1E'0�)�
�a˄%�*s������q]ג��`^��Q�M�G������
kH���/ʱU����R]V�ֽ�2��1���Z1��D���������n�o�w1n=�+b�e�2�`�VzH���YtT���O����q�\z���������z�0�%5�|����=�	XO�y�Oj�̱�'B�P<)��5X��:n�G���QԚh9֎6%���k #@B��W}�gdb�m� ޻r����brV]=��^TzNz���g>9�gTW�tR�ԴB�5(-,w.��o��Z�H^��Y")n�{d1�se�
XЈ������3^�����wQ�~�im*?*+�)ZLA��?�9�?��0|'d���-�j�������1՗��mW���U����dϕd/=:�ML�\�0��F�������
��rHrd�_H��E��,�{R݇N��U)����p�;��X���QA�h~5b=�\N��5��5���wYz#^u�N �]B��������%'��lsUqY���]{˧�?��v�;9g����#���j��sVE<����T�qڢq��u%:���9@Tfc�k�z�
�&�{}}o�Q-�B�H�Y�l�s8�6"�F`��G��f�w�x�ؚ�����q+�~�:�\mB^���礉�����8гTF�j�G�^Ȯ��Ff��֊�;='LeHK�^#��f^֝���mYA4d�G c�U��?�>��r����.�n��<�Y���~��g��;6���U�L7�y�<�R�:�$�9N�
/�Ϧ�0�R�ԵG7��W���Y����=�GM���K����N�[T�E���OE��I��=_��G�[�y����W�+{�,�̆�D�؛��k�Kv2f��ź�Bw�eqk�{k�T+�KH���J������;�+7BQd?Gή��(����={3�Oh5�/��r�R*t�ncvMV��84i5p�wQ��HE]�X߫꯾�gKMs��*����N����*�%wW��b1Gu�0Cw����dz�����8si��=������T%�a�aQF�zf��+-��ڻ�Z�z�����eT,RK�!�. ߥ./C@�Q�e��ړ3X:��%9�ۭ����ལ�Gu0�c�Xs�A��H���G̹���x3۞�*�y��42����+��\�x�N�G��ǫ��a�uv��r��W���]R_��t�Ja� �� �{��<k*Y�+�٫"�|��F`��s�D!kW8|}Pt�y	4�43װ��%R��Lӗɢ1�3��S=��R_�2<Y�h�����,�mn�>�B4�\����,�~SA�y�u��ȅ���3욁�m�nAV]ѝ����bG���LM}::V�/���3Q}�m��F��o�:�6;����K�z�l)�ns�/nm��\� �_B�:�s��݊�l����}&-nnF��gi���n����L�l���%�μ��lt�}Tr�ƏKϑ��V�FG�j3�zɛ�����;6H:��ܸ��Y��ݶ����yRFu��֞C4�h�#�e�x��\hq�+��*��Ssu#ʀL;Md���Pݮ�ɩ>qVj�au��­Po� u̱��L�b�H=�ǻtK<,���\��gL��U}_W�%�&�)廏�.���2�#�ȽU!Y�T�v�+B�� �g

\/i�ѭ^���A�r�n��4s{�����{������S���5 �����[\�bxZ�U�{~�����w����Μb��;KҠt��=ge�;�<S7
H.w�8"U�2X�DL+)K��u_�~�Z�{��0��]~7�WuDw-�PJ�L��-�9]�-aeeD�����u-F���]���ԢOG��|yGN���ٓO���$0=��&�u����1�� �zH�g�w2�,VG��ɨghDO��v�b�^d����Q�����_�>���yp2�)\���s�&���7�a�$~���J��s����!�a{�L��/m��e��1�or�|�jk=黦�a�ޱ�>R�2͋M��D��~�ytjQF&������Ey��ގ�,�O�~��Sb�t����tG1N3BV21��k4�U�S��,���l�>|���Ku���ءJ� V�B�n��?!�w�D��g�jܼ�;Pi��^�zX�	���߷��O~K)b;����׸	Ĩ�9Γ.s<8��[���J�9گi\���}J��ޭ�k�r)Җ;t��;��1нOf�] ���]0=�E�ia�w��KO���*%����W��x�X�|>+0���K��Ԣ+Giv�ƍ�h})��eq���ʛ
�[��0b�)wX��ΐ������]>��ZV=���2B��i����ܰ�QTvI��g:⥁���0e�*����5Yn�I��|��nc6��pЛx�S9igf�;��#p୫��ң����k����*IHju���q��J�˶��I�@`��ؾ=	�4�%�+�#���H���:9\86�b�|��6'\���ދ�;ͩ�Z����33B�_7��LM�3C���2=�,t�RRT�O*�>[��f��5#�����x�M�u0��)Cʪ�E�Чs=����yw:�	��^�'�c�*�y�mb�6L�p�&��'Y�J��	���H�۵Y��2J��J�y��Շ�ҷ�	D�6�e�˯;U�o:���ɹ��Y��]s�C�@�cNh$2�+=\�7ب�he��]��cN�R�š���66á9��`u�Z��=�PZl���#֫_d�y�5m��APu:����o`��6�`
�
w�(M\�±�3D��wYT6���V�U�e��n+]��[ǳk&�{F�{�u�Ԫ=�U�6�b!3t'i,Vky��0Eȕ���6��2�|�F[r$�$P��\5li˥�Zn�zT���6��o8P����u��Hպm��;v,A�Y�]�li6mܹ������ʝl���Gِ�s��ma�o%����x��[e^υ�m��������m�/z��I1�[ԝ�����)��uSG����
��ު���^�S�b�Һ�8�v�]���yt�b��q�"��Q�W7�fgG�H3����'!�d2���[(B�K
�u�]V�}ܯ)^A���턧GJف\�ػ��֙�b���)f]�av�_	n���L�D�� $[zM[ס���V�j���*��W�AkfC��r]0��+(�6���@L皅rus]VR���T��k���7��hg��u7��#zW(��\%f��W0���
�l�7�9m��s�����vV��ϫQZ͡ϭ��Y9J�{�5�oB��7�+��޸J��x\��+�bђ֗��9�ѝ)rAv��4p:��M��Z|M��[HG�l�X��`ϹZ=��9p�m'�&m$��x���_B@��G������v�)N�yg�'4��-��{o DU�8)����3�t;�y|���#eD֌{zZR���o�o{�g�E���32��u�%���eq��1���=�`w j�Sn��դ ��!z#Z�qЬ��˚�"��p�;+d�[�cǤ&��Z3MF�}��
�z�w[�.S�c�[�jU��{P�͙�	}���⋬ɳ�o�{T}ј���])��gX?�昉�"���H�(���w=j��"�
��y�6�:|��E+���	��yt/</w��Z� q J)�&91�SL���&O{�>�����y��>�qt{ǻK��
yJ��9����w4����V|q���/W�l�o<�>������{����x|���˓��s�S7��>扨�$��袣��Tdi�������:��Q%���G��Y�e���������z�T}����ꜽ�ī��뻅��z���8�����|��_�e_�����t���q����癚�gZ���?$��u޼p��uL]CGT��{ǻ�I�s�7�{�'�qL�A��9���u"�9���ٕ��{����P���=uߞ�x�)�^�;����tB��G�#u�By򸒧���;��2�I��t�3ԯ�����<y|����y�0ry7�/��n��Nq�=f(�=�ȧ��﻽���D�]���ɾ��_r1V�]��]��H����;��^�N��#׻]w7׼O��9*�G��.t�w|z�n������H[�X�C��<��D�+��:K�H=�i	T��ůM�8�����;Z��}��]��]W1_�=r.�P�`���������W�$�����/Kq����!��-��ܻJ�jS�����x����^}Q;N�?��r�]�ʀд�2r�#ܫ���ŋex���ۗN�J+��1Jqޞ�7gj��^d㎣��Q�Uʍ�dF�)<9�A���Ɂ�dm�D�B��d���b�w�YE�H�ŧ�N*�=��vGdk�3�B	�ۅp !��/Դr�	I�L�}�z�N�owg'����i�&U��]��dwI�+��Ae����l:�!�d�]*�?n�_�#�y�&��}Ĩ�n�����S����U���qu_�J��O��]&�u�4%">���F�P�V?����$o���;Cc���r|�t7a��k�e��~g�x���iׯw�iw��T
�i��(`�	Ň�P�-{U\��w ���v����4%�g<V�����p^Ȉ���
0���t��-!�/)�,�O��K~		G�ob��q�9
��yf���}�/���%��Ɔ��GE/׭�]_�H�\�ta��0Tv}�Gﾓ�� y��ۡp�1�-�/&���;s�5ķP�޺��	��˽��6	��B����������e7��{T/::�];�wklM��:д�n���c��ruRd_�	3rl,Z��m�a�	�6�Y��F�U*!�ْÝUM��x��5�͛��� �:_����������s��8g2�Iyj��6@ީ$7lk����\�b�Nb���\v�Q�Tf�Z�9߻��p[�f��N�������xM��ϼ��o�`8К�$�o�IɧS�Jl�����[HT�8���Q��4�ٲ;��[�Cfp�>���c��8W��H����n%����K�r�);^�'��2~�១{ �a�$w��W��"z�rJ�/�9�Q;�Y]u�x�UqJ����x7���++�F�c��s�N�G����ֺjF6�:����}ܽ�X�r_U_K��4ո1��}O�*\���5FY������yzW^����̙���T]9��g^ԋ�Qn|Qr�� N��#�V����Q�G�ْ^��{9�o���\.s����ZӒ����N ��E��N:��s��\�%9���فV�����O{ڹ�:�O��^KfC�p=]S�H���]8Y��W�ym�6F;��]�\�g#���n.�q�o���r����?!�C���A��*a�.����lJ��w[r��_�}�����Ǎ޲X���-�U3��d��{��Vum��6��F����!��w�9���$6��@�@�{��6gދ��Q�Lc�chP�tj��x+K�t �Ob���/{�r�!*�Q��wӦ䷠�ვ\��V��k5Մ-'!����ջe]5���ٴ�R�����0^�r=���J>7�NO=$O@� ��aj����R2\��������k��w�v������9��9��YA4���69aaN4?��5�>U�i�-o�����ݝɆ�5LO�/�BQ�pN,.NmF���V�)�|Qc����;�t�}}�
����v�s�zl(O;�����.��;�qmR���=f���3�����p���{�Z�����W^�}u��R�����b1�IL7D�<;v�
^5�e�C!lz����Td�w�{�y�y�.
KF��,#w,�>'/���mA�ă������x"��R��mg��ll����}U���QX��)I�q�ܢ�����Z��A���s�"�����\nޕ�������~q�v<V��G+�u�@�7qQB��Ƌ�S�^Ä�n����T�s�����L��>���SnZQ�%�0^����?�E��������`K��9Ӛ��Qa-�x��^Eu�3n����g�c�nqU[��4F7v���V�@�ެ�g�¾��o�X��Ӥ�y���$ۡ2�X�ӆqn	���%'����/��1f�?���>��j���!3�[�U����ߢ[�v�̫��ҕ�8Z��o����O )�f}���3Hkq�Vu)��5�Ir[�u�[��
x会R�O��3U��߳؈q�ǜBE���z���+���Yp�����O�)^)�yP�1��w"/Ak�ť5�6�E�R��#����.^f���ۓ��!�~�C�[Pglv�cI]kʩ{�y�"��g�yJo��=1!��J�=snV���+>K�Hd�(s腔���^�u�}.�x�
��Sݳ���i�<�D���"�^=U��ƏK�|F,�43���U{�׶��_)ǟ �����v��:p�
��g����_��E>{aI��4�I���׷i�F��Dg9���)�|���uQ��ڄ�P�3��[��1.�ט���V���y�-��Y�(N�����-=�@�?-l��z���w0x�n��9PDJ�I�P��*�d�A�.$+�Ź�<5.�n��V{��.��qk|T�Uj`����y]�ul��B����9����(v��qEb��	>B�h�)�F��@���i}�bz�	�;����7���?D�`��:or�_������g�:L��X'�9��� 7����͜���pm#۲f����?�\��aV�8A��J]�0n�O}9�E��$+G¥1ֺ���}6�%�|�U��ؤ�����h�u���樭R�����O��ylC�/�kVҲ�6�}zh������)�@^I���z����&�5�r �k�݂�G�0����#�>�7�|����t�����,ex˃�]eK u�xR�X%����8��H�R|�#(����[Tv=&� ���ӀyS�Ǆ�6~��[P�z�Lx?.�����|{��~�嚷�������9�7O1n=�%a�Ƭ[�ex�����}'%���Td-��#���dm�<у#N��q|%���6{���#����˱;PM21�.Q��A&l�8b��ic�C��%
�R=�1е]^.�������6��B��P����ϽP�����/a�nz�Eιt�����8���-��{����>jMF��{a�M��L^�!�Y����Bϣj��5�FTD��"L0�#ѕw]�-����9������0�u�H�����sКӺݑ�L�i�!('�p��\�!q�"�N	����5Sy����5�6T�ߠ(?�Hĝ���vU�����~�Z	���+����<YY�O��ݩ���E;}j�\ě̈�'���Ȇ���TsM=Ѧ{��k�u��)۴�S�����IV�1���,.��W�V����yJ�٠��k]Na�bQ%�� ���`�%n��5�4���ת s�$��9ݽr��fJՓ���T��7��oC��"��\e�b��N����(7�S9�U��ү�}T�W�C�o�7<���?� ���������to�Z��G�c���'�W���Y^��qϳ[��ш���)B�<���)������c��C��z�%�,��}�J{�����"st՚���u��mt_���lז���t䄎�t���h�)=e�)��k�-��#�f�V��\����6����%8�ņ������kt�P�
�_k����)�UcC�:�^�>�y�������Y��1[��6j���+=x䎛ɨ��q=Q!��O`MFfaI���
���o��w_S��]���b7<��d?^@pSZD��rR1���(��]��\�����ySz=8*:l��a�љ�8��m�y��t���'��j��)�F�q�&�H�\��4��ڑK�`�=M��GzL@�$�����= =L9�S+3�*��x���/�ja�g�}{�1��`�������UZ��N=谅��q~�ʩKq�vE>�s�};��U�y��M�Q�W��v&�5ɢ���-����ق�m�{����7�u0+�ɥ���K2α�*������W�~�!E�V�j�Zq�or��N�8��Y\v��v��S�^��ӥY�fto3\�Uۭ���6�(����ܙ�����%�K�:nu��h��&A�#�I�;f*�iR1za�򪾪֦d������V��g\���U#�Ŗ��*��?}`����0��j�^vW=�O��Q�s��U�́A|���7�8�ߠ�Ů���\�ܫ��R��v8�՘��g����t�;�J7�Y�����)�C�:~#����"��up�s���`��b�jmc���HN��v���[ayΏ�3ނ{7�F�����R.��Q0c�c����92'`F��U�����ە���v�=x��Sg��̯p�f~�7����]���D��kr�h;��ѵڧ%�+���+��X��}�S3=f����g5'�[���5��YA6@H�r
�C�ҍ�x'j��.	Q�s��\��ٿ���]?mG�nBp��>	Ņ�'EAs�%�S�Pc�)����!ߴl<����e�� lߔ���О}�Dt�y[����0�L8��*�-�H鼚YӼAW�(W����rPS,"���q`پR��#��;���#G�Ҙ-�CZWP��&~�P�A��Þ}2UB�c&�k��fhx*a
�����A9��>��M���p�R�?e���\ԧÞ���'�3���c:��{{���M�tg[W�	�0��џo=eQ���ڗb���V6��"�Ӗ)�Z�&��P�dSmd��%'RK�����f���S���ȸ[.�:$7/��Fl;P��O_=�?c�8�}$A#��U}_p���{,?��g��C6Y��,���RLX����;S�&�t��f�I�C���X�q檼N/ P/��a�U��~�p�W�
���Kӭ�	���*(<j�t�^ua��Z����������:|׾T��}���V-�����Ʋ���D��)G�U��+�bh�����eD[t�`��s/�޵z�7*f����M����[y��VE7�Uê
K��>b��χ���pB�>�����fwW����cИ��@O�
�2�#sa\�ـc¶��{0�]����ND����Cه\1��񰂒���!y���m�Ϲ^CR�ڕ|ѥ���S�dz�x+����2���@��8�C����B� u��I�E�W�-j���ԑ�^�y�Fe�������i�M���uͧNi�t�|�(/c�sV0�y��c�sO�3�Y�s���=��U���M� �1�a蠧��"[W�+21R ƅg����},{`oi�Ik�[[�on�G��F<u~�Ď�������S���=BGe�:�%��\ [�sĺ�18�Wv֑ݸ�k�j�4�Y���:+[�-���yFj<���v.鉛RHw��W�����J�3�sO�k�֕ƅ�yӊAC5p	湷.�v��V���DP���j�f7ԇ;0����y���9�VN\��C��x�>.i��`Y�v��7e!�K�1l��;r;K�е�	9�;/�'s�f�A}C܇��K���-�K"u]��ۺ��r"g��1�V9CC�,���'�uۓz������~�]�1T���cy��l�؇p�.��X���S�S$ �^�|�*��3fM>�;���c��vQ�Ê+��Iڭ�p�cpK}A��J�-xVrt��5�p|�����@*fW���ޫ70�Ǎ�`�];��wC��+���R���X`��ѓ�묩}7���F�.E�:ɝ�C�����]y6�N��q�4����A���!�< ���$�_�^]��q8r��>�.
:��+(z�>#��Q��M?z�ڇ���4%a�Ƭ[�}�mg�z#Â�a(��Nzn�o�������ك�O�c����h�;�3�[��i�N��=�t94��˫�y��0j��b���\璉��y'���@u�����QCF��FdG9y�{.�{�㱵L浵X_G��GQ�SE�3�zA�˧:#|& ��#�S��H�HB[)��O�9�E��%�ݛJ���˙��v�^�]A{���R�+.����N`�j��\��v����[�=Y��
|���<@M�pi�.�S=c�,$'���+ˣ�`������XM덵�/�}2��Z�Fc�\c�Sump�Hڐ䩗7�m�-t�O]��-i��<�N��W-_ ��������z��Y�����O�TvvWMKGQ�G^K��}��Y m:
K�r|a�:nX�&�: KQ�����w�u�64�X�^��י���Wnz1:P�}j���"�'n��֣���lm��҆ѣ�a�'ujZ��
դf$ʹ?c��wn�t���3�A�4�FR恳z���J��wv�1!�]}��'�YlƼ�Q���;.����S�6�(8�#�3��O9p4�I��B�pA��>��H�\i���-�t}������Rۥ��kہvKOe;��2���F�rz��v\�p����E�ϖ�|�1�sS�����Kz2�z��\�n��=5��$7�T~��Q��T¾���Ĩ4O����|�z�e�gK~�����[D���������Q�t��J[�8���F�F�?`�鮡��x?�=�S��}/֖����ݘ0��t��Y��u��]��EV�2�-Z�����t�MG���X5��|D���������Z�L��`�ܕ�o�R~�q�}�'�#p+b��lom�I�Y�676�0��.}�B��l�5�sB�&�d�P^^�T�,�ɝtC�R�4�=w�H�eJe���T����ܮ�md�oy�4᱘z�H �u�ڪ����դ�ZaoF�h�y7f�c�l�2�X��L�܂�
�In���X���E�tn�M#��˦1w7:�-�K��h����-�Nl{�{}5���fq�ۮ>����11b�E�E)f9���.�N��QVs��G:���1V��D��^�ؘ��c{W��z�ˡI%i^�vz������_@�!���/���]�B��m΁���D�W@�y�~�,�c�\�DqR�C���������(�O5V��
���R��}e䔻"�rnԽ�?:�"����gd�j��oe��2��.��ٗ���8��)�)�z�������1km^	B�������k�u�C��zo����y0E0���K#�6MI��Ac#�r�K�[��=���_��ô83S�m�w<nՅ���vމ�*�]fY�{��r���^�c{E��2��h�TuCm�JD��B��CG{�t�hՃ+sM�ښXFG���h��	�5�I�$;Y�R����gpa� 8վ��(������堷�9'KgBtm���:�wf2��X���s����u�4ûV�|�D����R��	��ӗ`5z*`�bgr��X&Jc)�J��B�9rCݛо�:2Ƨ�ф#ӯ�Ki=�N�y`����V�GZg��G\��] ��)	'4��m[��49�wX���T}n�l����E�KKw�����Ź�݋��ќ�J��|c�����#�4�=�Ir�U*mq�v��5�lDu,3.�i�_g2�sE��3y���{`�wzqܺ�N�,�#:i��Ӹ�Zt�e�<��L�6��s�$�y-�}�b+r1Κꂶl����۾;��.����3�E�zn*Q��5��K�A5*�lwiދ��7�wtq	�0P8e'�Q	���=�oM	V���7,��oF"B7p�<t�q��>h�����{��a<Sߵ̷b�o���(�ڌ��̺+d7P��bPb�܏R�RZT� �2��EQ�xPd����E�Mp��U5�\��՝B��)�.1���S6����[s��|�Q�3Ki��s��7G@��I۝�
�+�8��iF�u-ڎ"]bA�ԯ\}��xb+f9w\e�ʱ��jpխYץ���t:2�S���[�j.ԥm9t�N�}/�#:tڷ�u�oj�M��snCsa�k\��f�KQb��e��K�0��P���M���v�˩�䴹���عyͫ�NG�P���j����ԟn��;\T30��w��\�amb���q%��;z���U:�H"��;��ʖ%�>%���s��G�%�ٺK��M.�#�9��3�'5�r�u�e㗤�	�y�_g���A����1�ݰ�q�2A9�k$������9t��qۧ�&(8|��w��������}��\KQ��������'dU�V��n��4���6{����9�=ܿ��|����n�:RD�H�H�\G���C��e㓮d~��{�S蹗̋δ���w��w�u"Q*�0����h����7t�t<�_x=�3�-B㫨*�/��׫�=Y<���|t�<��._��^���x�O�?�/�~wE�%W���FE-5C-y���NނS���L]�I��u��p�"3��w�䒢z/oOJ21p�r=����"����<J�t5�S���R�wwA�x�ܣ�}��|���{�[~3����璹9�L��p�(�9��3�E7�O�B.<�=��s��%�"u��P�xW�)㏝��7�C��wv��Z-$��u3?G{�vd�\�#�	ۮ�!Q��pu���Q��%^o'�zN��zĨ;����g�����n�T\1,���3�����x�9$�g�
t:�~{މ�'P|t��(ŤDYP���Z��硳ϺJ�ֳ�Ou�#�����K�*t�\�U�τ#���E�ND��*�z.���5����=��Ǽ�T�Om5n���}�:Tg��c>i����{ŝ�J�/f�A1GY`�p�\ȕ�Kܽq`��G���+���Wumw,�`�j['H�m�ʐ�%��W�w_�����z�;i}R�O�R(���z=8*:l��f��b�gu!
=�iLeJ{=0�%�,U�1���s�dKv=yM)���R�:��W���lI���A{�R*ІM7U�9�/�K������s�j����Ƹ7�������'��h7>D�L?�,̎ƍu�j��W���
\���^��4��S4�?�X0�m]���8�?�ܾ4���^Cu�t�������k�hG=���/[�7�-ϕT���9cKu��v�U�vWn�|D������^�!���N�P�m��~�����q�w�c�~�%$>Sc�Mz[��D�ٷ�j��{�=b[/�F��b��Sd�$���5�m��>�caԖ����zzՊ�}�<�~�\��G$s�E��F8�,Č9��b�Z�0�V��yPcw�o���}�������3l�������md�F�d>��(:���-r�{f�˷��k"��(�����K���ő�U��ݷh��y�#VPM�9C�`�P���F<�twG�.���(Wݐ�������'IWg[�0#�f��Y��`8�\+���7:�v�`k\�oOň�#�'�8(w[f9�c�z��{u/p���h�eQ���f��Ӫ��%��-�j���Vr�НR��n���m���_}�uGp�����_d�a����'���	9V`<�'��L��K��T؜�Tg�����0�į�����z]-��lt7��GM�yw�`��aņ�T�Eb��U��;�K.������
���߮���p���'/@�~��^��{��;�)���1\�ͯv��
��+�^���9I�^7��yKO�`��yC��Grϔ��r�=�v��y�bC=x���569�P�2=�[�7ί��5��^�Ox�Tl���1�1��\�*!�����vr�:Cct�ŋ�~�^��=Jjz���W7���ͮ��c�Xr���Bh�Im|��>v��[MN	\9�@�񫍍���ڝ�����yyu�ݘc:�t�ԺL�1Ӂ*.[�b��� =����^�o
E����7Cy���v�=�V��|�d_�=p�,~=�R~]�4F<d�#3����F�j�!���r��E&6�P��z,T�$Xۤ!�޹�"�y]E�\?|����P�>>�U隟�=��2���x?K�RYi� ь?�躔��������^wQ�w��$}����RHwQ���C�0��E[qD39�D��N9�&Y��eS�k9mq��ƓA{Mcڛ��;�i?q<��LPAB}yGr����ϙ�#n9�/l�HMt�EP��Q;����\ł[C��wC�ګ�����.�d���&'�B��_z�{=^�=F�P�4�8����±x �\p��n��8�r�#�
MlԬ��K�V���_@���M�Ŗ�� ��Dۗ"��K�y|n��� ;�9��h�(��8�0ے�?���9���~���Z���c��w���jp��#�$ĸ�+B����Әe[��=~��p�?�m(E�
4�;Q�:��;���	�S��[�j���}N	��S&����|'ޞ�fT�!�O�Ϧ+Œѷ0����Z�������Zf�Et7=��f���t�[���_�8"uФ�8N��p��P��=˳�ͿN��Ҙ��^��l�4o�.�v�jy��`u��؄�}N��$ㆸ�ڣ�^XE�ɧ�gu��gz�y��I��mm�n{zviw��α�Kr�+����zF<Rs�n	M�"�֡1�Or�\�S���#�7h绽9il��OzXݤ��V��	�i�'�.<]eK#�����UÎB�O6O������w���g�3o�l����ǚM�A��}9�LC c�ϛ+dI޿@��5*>�7R�(�oDH����~���&k|+������f�R`�<�a����ʩQfSO�@6�k�p�2c��y���O"0�X�خT]Ey�� ��m��2PcE3�4mһB ,��r�Pn���n����ʏ�+ޡΔ�t��2��g�`&�����So�W���xň���з0u^�y���3�[�bV3�\�+�f���S���.�0�~]2{qu)��U\Xǣ��8��?!;����(�r��.(�w����E<��]�y3[��X��!�H���h�tPѣ=��9w�:g��ښ7~}�����gϦ�9������.�z�H3�t�h����#�T�>��B/F�O��)"2�%�z�l�T]C��=Saz��3mK�ue��?'�ZI�&
OD�ڍC�7�(?�k���ny����<�
8��g�K����\�U�z1:P�}j���"im	�y�c;��s������9���G��l�Ұs��!D�ˈ��W'wK���$?PΙux�k-p��xE�9�z��K��"��؀��%���f5�K�h���"[w#�So>�P��^�К�b'{ن.����)!w�`�	ۃ�M�4��F����G�t���.N���_�3�ߩC�c}��z7*	�נQ�����ڡ�Z���{�%���~���R������讃�~6@;��ݬ��J���N�Hv�^r�Wvdt�)E5G2�-��fk6Fs���bF]�u�
ŨAۃ��e՞���Ad8Jܫ{1:5-��{� ��TAo��LJ7�f��j��J�$��`ɜ��π��?�o^oO�	�ПE�_+�v�4���ז�
�eGc$��1�g�-����%Qil=X���v5��ה����t��!*lJp���s��&�w�Y>x+�h>�x��գh�7s� ����p�Tv{������\\twk����S�!�U"lg��ɝڦ�׺Z��f��B�t�36S����ы�==J�0ъFz"����1�<��e����nvc�ɻ��ǚ7����V���)�� d	I��
th-�2~�=Zz��w���]��V��2
�/ǻc�k��;U���{ �՞Ve'��X������������>�>�S7�+#��	5R�W.���q:=!�=ʆ�Ğ����di����qQ\��US�5V�#�C�{~��uNI�U�ϒ�{^tX�a��I�n[�3NZ�����ƍ3�	�]����b�&�8�5�<����"8�<�[�Xt�ӷ���s�{Ŗ�ʨ�Lu]���:�W�ɴ�Wq*G�_[��F�y���S�C��сڄ�F��{o�T��u��\�U�{�z�,Ųay�%��J��ҩ��A��Q%Wq�[���es���.���V�'���^������)��V´�A:���xM�S6�	�c���Q�3�F����`��JW��@��n�P���TϳL�H���9����X��{�&����`�f�S��Wr�l����w_��$��� �� �|0h#�a�Y�r��fwn;Tt"��+PV������.��ϼ��)9�8͏e�G���,ĉ幑1v��u��)oN����Gy����xl��<?g�_��i�gm��}6��7܂�,!�B�P*ce��v���U/��XZ�j�:�r#;[��5��q.��������Htr1�6+jMY��|�w}>�ޫ�a����,�)��j"x��[��*��8��9��K���?}Dc���D�o�j��xh⋶�}0މ1��i�~o*�}!����x^�~�����p�SP��L�r�22�ɼ��A�8�������.�z7+u�!�{ղK�RS	yc�[�O�n�N��n�LS�"g�2��\���~�), ����w.�x*������|S��a���L��i(�}Z�>�!�U��؂W�'�m�3�,�(9RN���90?yM�uYu�MQ��F��3P���\���h��;<����2�;~U�>��eJ9B!xy�?���������ÌHL��ʶ�K����B�ٔ
���:����b���<�����n�B�z,�G���,��G��Gp�ڛDб9p�㋶v�%���[:��⹲��MGCxݴ���Ř�2#�#��s�)S��)�Ӗ++��b�{�WϪ���}�o6�����ͣ!��M�)�b����Ĩ�x�[�p.�dp�YR�c٤P��)Z����[w-�
���C�|rh���0w�1ýJ:4OS��>UV��M�>d�#
ߋ�u=�誌��^�`��'��䎏x�����z���tg��_ø�ᨐ�<30د���u12ǲX�6C�W�Lϲj��
a��]Jx񰂒��� /3Qlv1QZ��+����p�K��u�s��T:-�M�?.��r��V(Ax�pC�C:�s���#ݔ+{�LV]��1Y�k���	?���H~����w(�};��r9�:D���`B��ea{�!�'hͫ��\�Y�^L����JizAГ*�_C�,�St��h&5ݏ+*������)^�v̇PX�9(mtq�c�Ok#V�Gb��Ҝ�&)����U�������~��)�,%<%�pv%`���{�ȋ�z��a�Û}�=�<�7�l���T{�i���uc��%���D�>ah^"�omu�B}���L����p����:M_��c�2�	GN�ZTk]��OǰR�i��(EU�.O`�t.Q]Y�"G-*h����� 1D(}�4n潽������޺֑�����0V��K�{����z�fWVt�>��L	�E���0ɛ�yV$���V����dʙ\�E��~�����Pu�|�G�U�=k5�϶���lqEj��P����g�:�¿^M>�4\ƫH�Ԣ�$��]]��HyUA?��w �5�P��d2:�&���G��V�b��zM���m��W��;���jq�?d�۴ؚ��*aIO,0ZG豕�.:�Կu�=Y1~Y �h���N�������8�ne�c���d�a��K����D�V@ʸ����|)kN����z���`1�����o��z�ڸ�"y�q�JÆ@ƈ.\��Sb[��uOعDɭc���d�Iɨ1�1�:ȷ"ПA�Gx��w�tG1N;�pz�wyJ�K��T�͓�.�8/�F}u���B���Zv���X��bG�C��v^��~5��Nzo�@��~}w�=ম��FM �'��8[�aY���S;���Ug��h3ߦq�=����F�����{�n\�c�w�y= u����ZI�*�ʊ�����.��.9��-�d:�J<G���G� �Z]H$/3�'c��N�"dk�<C���p��J��(1;z��?���ȁ�|����~����N�4�NZ�A譊��lu�oF-��<u��xT~p����f���d_f���ٿ�KG1I{I � R{�v�X� ��{Qw�����ڗ�e����yT���}ͅ2�o���9ݽ�z�|b��V|`=�����.^o���#v�W��]�dwMO�8xR�jH�9��FK%��nB0>��� ��\<�3��P��K���G���OGY�9'6���h� ��P�}цF����ע�� ����~�@:�cƎ�Ζ}>=p�}A�[U1>��{�9�Or��6-Kf�a�7*	�נQ����\'�����S쒍��'��vw=뫷��Ք\d�α����=�k�BH���ʏ��0��
�V:�f��o�Uy�]:�sE{_�um�~2.�/�Xf�ҟ�H�W���RR�Ĕ��H�Z�?XڣSڽ�Pgaf1GP�;q����M�1Q�eC�!9�Ƴg����k1~�n?'�0Z�R%8������ک��#+��R�Nc��P|�^jT0k�&22���a��(��t�%��#+���n^wg�N+ksҕD�"��=��/�b�O��RO]�_�����b���U$c�����9ު���5�Z������U���ӑ)?�Zğ�1�#��@L���n"v�ׁ��YOs_A�k]��ܒ�хR��]�=|&��3�����>i��{�,�����)X�2�^�<Rz�M�;-�jY7se���F��A���Y��2��س;^�x,d��^-��вU�ّ/����i@���\]|���4�ޛ��T�యѧ�����\78��-��2�}>�ӑ.Ld�XT�n��&�UV�|&�x|��n.�/�c�z�N�U�n|U�xX0�h������г�~Z?/M��Kߒ��}�:�������ި��6�2��k��G��,�>UE�~��[���j�/��I���~��&l.s��b���т���
q�u�J��~��k���q�O*�<�Ӆ�~��oFjBe�2��m}^Đ��y��G>gZ1���rXY����F>�^�������n��n弾�(�@�Τo>b���Q��q�J!�c�B�Q���t�r�|��2|tC|�{��e��ֲ�{˼xOr�o�ϡ�f �H������a4,�h� W���Č��9���'�^�:^�1����d�{=j��CN>�æ�&̐��"O�oAPss�fUv�sx?��t��N��:~�dO<�r9V`4��N���.[�u==jq�޵���_�NS��⎍\|��幓u�{}�[��tW#,7�8\q�Ss;;[y���H� �r���rM���~�s��(f;D��:k{V�^�l�I�;W�P�
��2�&�᭘ڷ�>8(��6�vGeL3�%)}����鮳��.�<��Zxf|NI��VZQT'�/(��0�q++���$�ݥ�T��Y����gp�%p�BWWB��Q%�.��b�j��+��f�t���xz#-D2=����d<�e�u$�cy*��1�&kUn>���6��g�6(.�������`���M1f�bH+�4K8N� ��>�2����؉N��ʭٸu���.R����ֶ�r�`έK���:r%�x ͽ�������w�jVr��VJ	��VP��'ʳ�r^�颳�ϒ�lS��������@�ݧ���.Ն��]L�;��
�mN����k��Z����3��#��ۛ��:Q�i�ۊ������{�n�9Rr����n�;��\����y�F��2Ѩ�>�HnMD��n��w��Mq
�h�p��K'00;	ّ�v�M�xl�R�4�}�ą��f�ޝ&�u�n����k�Z���N$2[���D��@gfV�|�z�u��t]���]����f��c���MA�x����[`�J�G�R�����- ��7kr��ު��r��vfÕ��=�I^�ʇ)(�n��J�o�+��@Hj�t�*�Ĺ���;qI�&_\B\u���ܙ��.��LJ[c�Oh�C:B���m����8[fhK�W;U}�,$/X��O݂��k5ΐCL��g�rd�6>['vK��:�5H�	J�Z��v2�o�����=��n��Y�N^���GY�/Y�\���&�	P��
�xrܹ;r�[6�mv-K�ܼ5w�����PUn���Y��ԋ��rn'/Au��j�4	e�GB���;�e��B.ǳS���[�I�����sU�*KU ��3r���':#A;aM�\5�=�+)�,ڛ]���r������I7FenLzP�q5E�՝�J��8�g7���M�*��hk�̚��'͡ѓ2bk���,�uYWjR{ox&HR�`�+Y�K��y�����u*A�g2��/0��
�j�r�k�����ɫ�	F��!�T�K���(�+J�t�3�'��T������k\������c������e��.�%�uoEܱS�Q+FM�7��ۗ[Z��|�^�a*Zy-7�p�U��`N��:X��������+b]W���4C�vL/	�pSt��RFK`R�U*�P3}�u֊�=V�zs��:���`���9�̇��<�E&I����K�������&�5� z� SUׄ�Z�Xȥӎ�s[�����`P�Zc�e�Eu�9�V"�eԿ��i���9�z�#{w�#لM­���[۶
9[��P�����jB�;x�C�5dlKr�.���p���Q����N2l�{��u��5�}:�!�R%���y��9�&��EZ��B���#�����a�4�7t8[��w�y}�}�p��{��'t0%e	Rݻp��У�D��ۯE��nI[�*J]�w�=�QJ.���=��{�⺹:�B��㓺O��#y�:��s�-��:Vt�QE���Ĝ���w%ܜ�N�*��\��'=�&���yE�Y��5��^��������KB8d$�B*i�y�*�2�7���~{��s� �|�QP��
�Z~q<�w/T�9�d%G�#����FZb'�����FK}uZEϬ�nZgI���*gJBB�QB�/�"�x�J�J��D^nX�*"�}t�TЃ�Y/��H�j]?';�BI��z�(��Nq��[̈-^��o�9D!�1�g���3��.RXIeU',�k��s#X���tE�%�OK�r!E�s�]�%,�Y�o�o.\�c͕��͡QY* �O4�9��t��+(�04	w	�gDA �%=5ف�ѓ[W5����~�8Ȳ^�^�:.(�C:,d�[]��x�;i�����g:�F��`ʮŎ�[�:^Lދ�/����l�oۚ9.�G�+='���i6Ť�sb�i����ɏ�����V�/0S����V+U��	��1�Cﾌ��^Y�ZV�I1��$�����-O�9��t_��UU���/�j�RBA�pBylA	�ؓ��%χ*I�1���x���{�N.�gq��׽׎���,�X/h��L9�ϼ��$?P�d&�ĩ�95�+$D<�+�������}������W����i����>��bN���x�wn��q�zX������U�U:���M����	�0�������Yc��U�V妬��l�T�V�MZĺb|��w���'��P��|��c�w�a��WQ�n�;{���|vU��^c]�VX�$z��c�"R�Rf}�P/���1^��A�6R�EC�o�b����Y�WJ�5ٙ|�F����x{Wy���x�\�ȜQ ;�X��^.8H}3Gt�P�����a�wwQY��x�������o����no>N�#�Zj�(�b8l�����xl������#�2<d֛��|(�i=o}c��eͤ��U��j*�H�E������Rop�K�kާw�<Sɧd�X�iQ�c�y��H��:@Euc���^�&�����m���9�&����:	�fB�t{@ov�[�sC����]"��������V�ݨ��dg�U���EKϑ���V�FbL�c��w�v�����"e܏��@į/F/{��A�,:�Δ1(|~�Dc������OX�-;Ix�9�~$�q���y^[���i`�=J�W����m�P>�p�^\i���)���N�]���n}�f�CD�#�l�n8�R5P+a�$�5�{�PU�=먆���Ǔ�+a�z����oN�k0u[�!;�[$r������8��CZ��j"��T��^#�qfc��c5	ת�1o�e��[���&���!�U²꼚�FЈ�B�0zN�QbYn,�g3��02d]-���5�9�-���S
S4ߚG豕�.묩g��	G��C�^�|ǩ�I`?�'vG�޳҉���wPa}��>��!������$�z��P���{"�ɫ=��8�u��<��������|�>#W�,�SE�2��q�|��xw�����F���W����L[k�^�c�3VI��e���a��a�p�Ch6�� o�zy�w�$�FN�=�w%�3�#/���gq���li�,l��s5e�iu[��N�NΥ�{jR�۬�p{d>A��zਯ+R���{ë0&ŎD�����2��+Tnj�k�H��ᶍ���+{>Ey�c`=��ե;t*ʉؠ�Q����y�J-�R1�t���UMK2v��������X�==���=<k�b)a����,I���F�ಁ�|<�3���$+�����WPƋ�_�5v��)��厛��F�mE��T?+Ϡk���w�۞*��L�onR��xi��,Z^�S�6��|͵/��a���G)W*4	�>�u�����7Qӗ7�P�����OH�a�+|AX���O����).tt�t�P�O��}����Y�Qx���Sٛ����Qk�_Y6q
M��=����]Cf=B��BL����]��0��8.�^��˫W����µ�Kc�/ ��CB�6،vp��Yp�o��gM���d{�/-�C�ו�&�ng�{�Z�K�����L��A9�H[�(`�	�>jD��U��O^<���gG�6W40�yz���VB���E��gr��� ������N�j^T�Y/:��$���?v���˽.ud����v�����r3^Z�y:g(:;�OQ^�]X&�\V,�w��xO�!ի���{��$D-��S�%M�)�-�j-N������|}y�Y�Ơ*R��Y�|���G|�k��ݵS�K��r=��u��9��`�[>��>��|a=f�Ч�צ^Aj]nX�6Ѵ#�L�K�..kDϯ�붧f]��v1�H��oݼ
����Q��?`Lpk�����{��W,Zٹ���W�]�s�OՃ�{�S�Oa������.��+l��U�ܞ=wk1F+p	�e�>م�vftU��h3��.������Z����N,��%x_I�w��5�q��?E�UW��[�Yz#=�`(c��'�E��O��J�!d�X^�c��p�=ZG�|�`ȯO�A����L#'�}�Qv���p�԰ʽ�@]Y�#$�Ҝ�L�0�z�*�?x�0�Rf.#+�����޼ctK���}'�� �W�|��-��0Uo���b\��L��~I�R1�g��nYp�G|D�}#s����R�9s�Un[��m�]��΄K�x.4��o-�j�l�!LA�);��4�kj`=^�R,w[�*��?GX/ѵ�*����&v||i�r��wa�u�$O���!�ѡ��\n���F�Co���?�n�x'����-�=��z�s�����)�ū0*����|獵��5�}˥�{k����L��O���V��_z��ǝ��Ca��N�����Q��|{(�1��!f(�,��OR���T��Qے������\(a��0S<�ʑ�FE��R�ܵ����Z2�8%�yK97���T%u���Tm��d�z���K�v��C��6��6��N�X��v3����ƁJ orn�(��k$�7|U��vU�_��E�)��_ϫ�;mK��wn.����=�<l������ە������1�ԤM� ޅ��\F�'m`9�5�B��7�ۨ�xe��ce)w0�{��ji@މ�/K	u�{�=)�ђ�5]p���d���|����Ȗ�l(�S��4�)��j"x��,r��xqarsj6k����AFuY5�Y��Tz�����X~(�}7�6�W��c���w6<�����9���d������=��E�}��О���[R}����A�ا�/ܺ�&=�����[z���^����{��)���0[��!�U2��3Im�3^
���W�U�^CS�K`>�0��3�������l�C�ă��LC��bM^đ��%�E���`�~�jU`�+�~��>��������t�x/h��a���L9/�.�4v$��Ax�T����{I(����>���C��h;~���4\���pk��L�1Ӂ*.^ �[�p.#<�^��;�V��ɾ�oB��}t��`�����Mُ�F��G�z�tl�8npUn\|^e+��\઼?fdk,U��)���bi��c9[�W�C{$��U�Z溵��i���W��������D?_	���s�Τ,:��)d|���i������-��T�	�0��Ztg���)�d���N�ܦ�˱��>���M�ʪ��M�E�����u�E�rOq� ��}�2<Z��pB�A�l�#���/��W�Z�*>�v�Wz����y���oO�p&�F�}��,��t X��Z9fC���#̏b��\��M���=���/]''�})¡�ozli]g�Ȫ�D��b��T��Jk���Q�)<4T�kV� ��o����-���;Q��r��@�	�<�h�Ԗ��ĿR����[2A`@��26O��G�`G�b�V�Fg�2�}}���������ޱ���;��]��A�t����t8Dq�ѧ��F<��ϔ���	�S����T����.�zc��}�/�~C���@�A.������p��dF����P:9kd+�4�UR���M׹����\�Ϻ�'u
7��1ʂ"W����8*�\��nOg��7,ly�c]޻�����WoE�8�0}��-թ��!zyUT%��C"T�T�*cEyL�s�%�3G���q�3x��n[^�������q��X����!�U^��c�';-n	�0-U�*yg'"߳��G�<ez�@��EOm9�W���+B=��4)o.ș;4v�[��Yxj�QC�Y3�'���kyw��a����mw�����|^��0��U�uǺTm�2�f.��V哰������S}c&��ɼ\?ʯ��Z���M/�{�+#�������c�A���PF*aI	�ũ>�=[��'s�{.�:/�y�﩮k�B��C���E����){�e�bϴ�����>��!�6-����ĩ=ý���R�����R�_��Mn�U�3�#��V�h�q�y�q�#c��(elm�>�}�|��c7�.U��uu�d�NME�9�
�,9�����?!	�.���e��xwW�W������xS��Ѥq���P�y3j�O��%�=���ڔ����﫷�������4l��~G����SW�7�E�3�zA�s.�X6K0�AJ���󇈩�t�O�;�����p��E}��llڕ ����^��~��3S%�^ݷ��g��֡k�o�̰$NEpڈ�X��8���V�ԂB�=rqV9���
t����LB��^i�+��C��!'l�
�6�M���V�mթz����i��W:��q��Y�������80^���X�+$���81����s��ڻc�}�����6�NVp��}��3��-W�`^�`wA��{勏k�_\���Ӱָ���,�yg]�$����N��	b�n��䩘S���z��vI�k$v�#����f.�PŹt;r�o�ա�c�.��>������5Q3 q�S�^�Y���s<��]o�6>�y�UB��ӝ�sT��� ��c��x�l~�cS�h~{��h�y�[M��1�,g;��N�$���J���9]�N�A;-�@������\'��6�ʱ���Z��~�c��]8�B�#v�F�zެҙ�+���漴��t�����I6+�e�8N����-L�'�)��"Ǭ��>�^�o�$D+��I	SbJqA���oy����L:<�=^;ڢK����ˬ��V�G�L0�{�d�Z��ܞ8df_I/-[G9;��Oar���X����{�̽��<�P^K�C����
�>0����2e[�����*�Θ��C�\Ewֱ�o
Ң=�Z!1ׄq�����ǔ�~��)?�]�.�2~���}�K���o���R�ꁸ���>i
q�S��+.q�{ ��x�����Vq/!x�V��CR\H,�>/V��02�]��H~���z��ߒ���j�<�ˌ�ܜ���?��b�{½jɮC��W߳hT���XB�z�I�n[�3N[�	(}{uM����ҽ���������qo0bZ�^ʼ.���%�Gfi9|\rn��~���!Ɲ	6Q�B���ܶspv�[�9��	�ɚ>{jAf�1�GhDVCF֕�q�k+�1>O���&V��bݙ�ƃ���c���i�x��`�+:�\��5��4����&��ۄGF�9І̞-ʙ�)þIq��V ^A�`��L��>�#v��K/;+�=�c�q�X���_+���2�ې�:S�ϱq�U���/r�%�m��Vl��v�)��T!���C�>����Ð����W��s��ELe�ϣ�P��G�1�7���u�Ϙ�r�TrXk�G�D�q�D�I���$��ct�wvZ���6/�Xf��B�}�u�*0y�Y7����7q~y�]�.��o���U�~�?���^���"A�H�Wj�^��+��<q,���%���G��=�~��(��+3�/,φ��<%�(h\S��L�|��:j�j�=�E��0'C��8���w3��<���
Vdr��p19Ve�5�Ǣc�o�&�̐q{|������w^�}.����!T�L��#�5k���Z�b�O�p!'���-����Y���2U��~1����u:}5'����ts���-wM���@��v�FT��59�/P���K��)�s�n��/�z�Y]F�[�r.I`����=��h%r��۲�x$��]Zv�S۔�a��vӘ�5,���6N�RwX���*�d��o0�=���4�]�^�}�scr���".��������a��vN�ԇ�����^�hM�q0�2�}���w�3�S?u�D�FxE�8̽�[��i|�(zpf ��/�N�;7�����r
�X퐚ؿ�6D�����z����V�q����EqM�r��M��hX�j|�Ds
V��k��~ДdOvNj�;~��19OJ8ݙG#�!�"��7�56�����b�z�m?=�N"���"�"g���w�{��4x�
���:�sQ�}{�Η��5���-��G[��qǆ\���a�P�P}���޿�vy(����5��]��|=~u��M�mޫ|�s�{�ϡ�n�]v6w�W谼�I�淢��~�N���� +���w�Ϫ�-�O�~Y��&to��_R�{a���[�}fT�>���W���{�4>�G�{�Wz�z�dH��]}��
���Ѹ���7��s��{=#��r5_\,�����):��,��?7�ac�/����JJ��x�����>�f^�XqVuO�_W-��9	W]����y�T��.�}B�i��7[
ER�W��ۈ*JD����˨�0*-�[mn�7���T��@;[p]��	�����9����6AO�o�N���B�tt^@9���t�w<r�]wY����)m�q�9���__k\��V)���r�R��� ��8^EUm^���U��<3C���2��oC���1G�9Bw�S�Q;dV]-W7
�α{�y�S&���U������lz\�k]���'oKp�96=!e�D�w(�r��a}�Gia��/n���y��cYt@�3/�I;)�(F�E�$+�L������Gc��U�ξ��;�4���_P.�.�q�z.`���L�6̙}ér���uԑ#K�2*��@�P��0i�M�vH����n��l���߱.����ub��p�������9�:6O �:K���v�U�
@O@�}�WJ����2���(.E�ɕieX��dV�����"K3)���׃w�����cd��K��˒����n<ɝo#��-��_S�-J\q�V#����C��
��A�,�.�hڔ$��t�$�Ugs:=�<MS����a��wK��,�xE3NN�MmP�(5�uN�5:"U@X_l����F�"�ᒦac�gV��ַ�/+":�W(Q8���5wu�y<��5�M,�Č|+ 7s��7�#6$9.�v�p�Q}��Z�$��f}��R�j�������!��5 ��S�!o�]s�V��ӕ�����;��b4~��w}���&P�/.v�� �Vc�;n�B��m�@,�e�>G�f'��t74��R�eX{��[5�&{qeeFS��k���؞�6tC�`���F�6AK�.lBI�S����V�S������U�����tԛ�Rvt���j(ft�'r�]����Y����0:DF���\ܚ�Vg1�w��M��Qz��ff��4(��/��73�w�fU�(�O�+i��+v�d�G�6��������/(����1ĖХ��M��Y�fDs'Tw�a�mWj�������M���9��n���Y�r��
��N�-�`)����-�>F������f��w[��	��j�u��s����*�$��qmZk2��u�LjL�+M��R��K�Ř���Se�7��b�a{�ueC+�ޅ��=��b(ֳs_�{W�*��<�uB0h�5c��ĩ�Z�m�Y��+N̸�7��E�%Ǒ���L����zF��쾄��fF���&���#)E��t1�B��|��W\�d{
���]��j��u�º5^)=q�E^DcݰZ��Zg�;���i�%n���8e���ؠ�ݬʐ1���v%ӫl;,SS^U=�Rs��ٚ����G	����Ket+_)nbf=zqKBD��ڕ�W]�~���2��#���(��A�I6�Q�bUTa*Q\��c��B?w�'�ȏ��Z�D�H斝(�(�ʊ�����.N��7�뫭����xIk%I6#�S����I�n�冕"]�<����ܰ�W���%hmk���!��J��d�͘��P�r�٩s��$�+�z.d�j�U��^�*���ŗ9W�(�d�cݬ�zМ</����,%�͗�ԋa�*�r����s�I����D�T�"��ZЈ��\���K��/i�EG5��*!*$�YXrI�#]�sB#����&e�<�NV��F�"�z!yz��7
)4��D���j��L	��<�TG4n�ES�㺻�u)2�1*j,"�trp璊�!�H��TPr�a(�ܶ�We���"�)����Q�Edҭ_';�҈�B��rQB�Wg	H��D"	�Rg|c�[�!������h2T4nĵ�C,ޡ����/�E���4KB":B����;�`L��[�$Nb����N_!�A�/�����u�!P�B�7��5>��o���t�1�EX3�+9���{z�}~X�^��׌��*���T��p�����K��{�v��w��X�Y�k��s)Z��L���z�Ւ�`�Q��#L>���s�Zw��f�]è{���t���^�{�;�B��~���>��4o�Gw�X���{���bl�_���s����l��Č�VW�{�>����Сc|ŏ����	ҏ޺67[}�L:�� ��c:fc��6_?v�|��|/>Û^�r���J���k��z���r�dD�ꨓ�^�AўC9�F5l��a?-�X�2��K+��C�E6�L��gc�kЪ7O{UI���{]�H4GM4~�͚i�>��rנtE� �X����m��gz��;�v�	ш,��s�u6��i����r|'�X�2����%T� �U�E����^V�r[�#V1�Ν�%�L�?�H�_z?'�aE��s,p9����J�gI�[��;m�]�(��cV��\��'F�̨Z���/`�ne�}n�Л�A8D�]�h.��2�^z�ӏ���/s��-��O�PSzn!"��C��z�ʷ�&�A�Ƶ�B���_O�dqAX^�v��nZO��؎�o�;G��*�ge�9��A���8T ���nm�D-���4��#�k��\p�<�T��]�<��j�m�A�lۑX�О��ݧ�Ryz�5�wշ���{f�i��T@��kq Oö�ʀ�������Z��ܚg�oTF��!�4|���~�ϊi6�Z�6��V�â~c����ǆ=jA���������oȢ�������ޞU������U�5Od<.V~$O~����!�S���=c���c����G([r�Z-+��Ӟ��Nώ���u��*$x'A:��o�^kx;�{��o�6��T�=������E��A�_@�te���8:���_],o:�JZ��w�LU\Nm{���޸���{}�k��}�rS��v6��q?`ꯃ��aX.����+.�P�z�]�,]�Kݲ��Eȵq��À���o�f��z���`� �"�a��D�5�5z�L��	�[*JY�䃇��kGK�������Yn��:%Q82A�[9�$#/��b���sʺ˫װ=��m��6Rr��m�jj|'Wf���vj�ϻzl�=���g �al��/�^U�϶�p,��A��x6kЏ��d�{.�w�w^K����^�x�	��[U���=�r��bq��������D�����Wp���8��XM*o�M[���fJ��[�{��G���]�v��4S8��Z*���x��nC~kM$V���w+z�"I�w~~ި�Uj��b0�k�eKcoo���&���w[o���xa}S�]�[�*͒W��W�{]�^G���n0����ìw�ӥ��gz��P1�=�5����{(�U���+|����N��u`.��ʄ�%H�
�!��5��ϻ��ye��^�$��S�I�p}��*�vƱ�j�%���~�C����4*G����=l��x���#q�O���遪[��d�]�l��ڞ�[_*�5P9>���V�T��^���e����2A�q�耠*���˝��G����X@��\%PO�Wlk��K"r��y�ʰ�������s��5�R�Rl��.�o>l����vM�;"=m���7ld�9��M�V�6���RY��p��f^ˢ�7xVf�>�7�e�3a-����ܫ�+�@5��8�������]����[ےڲ^��Y9¦yU�憢W%�����<�uF���U�,�\�p�p �5s���>�U�{zvkl�4��'��4�U�V=P�#:�[l�T|�I��6�r�9{��k8P�����k�h�}&W��NM�}��b����{;Wfn��ګ����&�ቆ�����g��y.~'j.+�ؠ��;:�{�/�1W�=��z��u��m�a�������k��j�_�e��<��l�X.'�+7�hX��F���s
V���� r����[^�{|��n�|�:=�yAuk�hx�Ƚ��Cq뜙ɽ�=��؞ڭ�bG��x���SE�)r&}���.�{�aT�2�J񨑃_�N�K�ż)Th��m_5����i���x��Z=�1�l�HL���G{î"�r�Fͣ�z��[|Zu�S�����D��	��.X��V�'!諠!�SB?3[[s���2$o6�%���ʛ%��6�	ފ�v�=��Lo�`*^i'���W0aN�<�`���tC�����ս��i�԰�X�61�c��������������U�C^������F����ⶀ�0/Ӟy���lh��]�B��?w�$/>����ޗ��^dm��]������m�Y��w̅xx���{�2�U^��Ǯp���Wz�e(���(�����-�7�6��{�Qn^l�̻Ȝ�7�۔�;�*��ۙ�^�]���~�.�\��P�xW�Cݫǽ��&��U5W���j����ן<x�ϓ��	�XZ�|�'��{l�7n^���ޭ�nvv!�;Q�tmw��	Z�g��S�٫%l��O���<�]��/�hW/z.������ë��bw$,�j��#�m��҄��z*��W�ժ�<V��1PY���gǳ����bJc�r(+��*:g��xY��q��;�A���7=��'XϽ^�O��G�c�'��߿y��e�C�)T��w�h�.b!e����̊�9�z�|w�	dZ$Vvge�6�8-̟��t��²��h^��K�25�*+ԋ�NHQ��4Y�����z�躔�f�T�-��yWM��`�V�D�:�EB�ڛC2��	oNJ�,�;/�+��ͮ�ɉ�\!�}��|���#����U���yC*]|��G�?C^��'�����&k�Fh���#�G���e�VC��$`⧽�)xwM�;����x��������ˇ0ց�M\���d�]ƚ���]�p/-��>��jM�y_��� �E ��b��+���4��j�rdOs,��W�3�4�O{V�t�ѲX��mFGF�"m��5��I�~��}�~!�uT:�c	X���y��|`q� �AT�{��h[�Ey����f�>�m#Y=[}�tGd�;S|���屴 gT�<7��?u�]�!�/*��וOٝ�+�w��ŽV
�T~��ac�*��dCp�v"���̸́����n뺯���_?K̥ψM#G�k�,#ld�-��[�n�U��G^]�@�"��
q���J_j
v�W;�ʺ��Dw� �~��{´y��=O|���VG,�8˜#c��#�r�&����&uL���J� ��2@�Qp]u�����;��O��ǃ��tJ�u�qwMT���#2i��n;KW4��UO�K�w��1�wy\n��t�]lH�����R�a����k��)Nc�|�P�K��l�p;�yfd�ǚE��9�}�?z����Q�滔��~�lr�Z��ާt�)~��+Rdm݈�L/�'Z<�z��g^kx;�W����&�t���Y�=��>j����E�>_&>�^�k����AU1�����u敟-z#c���90���{3v;���w͟��Sm�ѕ{q?`�a��0��F����c�O{W������c�9�ke5�{Kʹ}L�������Y������|KqH����&t`��g��os5&���������e!���'0�}'��?`���)��xvj8�k	�V�j�i�@�z�+�U�Ag�߫Dg�����eH�
C.)�@�D��\~���t�S�Q;~��U����6����?	���]�S�2�����|zX����_N?]�J�3˽=y{�1�y��:݇�\�!�>ߠd��=϶�rk�_֭I���;W�H%�@�XP�ʑ�Ǡ���w8��j�tc7��ǈ�\��d���φm�z�v�Xz�8Dǖ�2f]�yT��4p��)c	�yÞ@{�|���D�;}��6��U-ہ+�A��.á��pe�B;V�e.ӆl:��7{�o\����頱��OP^��oN����9�#����3�Ea�7w}k4�D<�wjZl�7�� +������>� ��6��O�O���ۑJXѯ/�I=�j�=�u��~�e�/7�c�4E�As��o�j5��:���2�/�C�	d�k�w���>?)ק仏b�(8jKWuy�\\ܔQ��wѣ�Pj�o������c]��d��"��&�Y�EeN����:V�|D:���#���~[K[ؽ���I��[�E�^H�:��v�#���'m)���r�z�XUCFsr�hX�r]Z\w�[�]�Ŀol�M���Tw�ݾ�y�����g�D��v$n���s9�^[��^�6�#�,XO��x��]�G@���[ޕ��)��Ǿ��{�ߙ�n��W�y�|N�@7������$���}>��;mN�nz����^R�$���%	}΄�y��Ux[�a�(�C�n�n�:�H�I���\&�V|�!j=̧�ݛT����5`1�O9f䝃��B(�s��l��oizy(ʢ;-t�n�X8�!N�d���(N��,�m���ên��{���	�農��3���0R~?E�7<ѯ>����6f^ќ�t�R'�z����u���{���.�"E�����]�RTV=�7ʝ�����/o�}�}�4�M+���>񗣽��Kc�Fx�$�W_^7ởwtxÁ���v�[��x#��˺x��e^�)�W#՝�
�3u[�S �\�#ڨg�|y�X��n��_,�9���;au�{P��̊���	K���A�%�jh}����ꤼ��y����U�Z�rZG�G�~���&�w7�Iv��.�|�z��� vО\�]�*𢫼{�8�o�)�sUU�U��h�>&���,#o�	�@�7�����{QhGc������g[Ξ^���2}�?]��[}a�a
��B�cz�7_r�%��sV�x����:���@s��s����k��}�V>��{SXnӨ=As� n���k�5��e�m��dm{V�U�ݫ�������z��y�=n���
c�]���ԃǇs�]Z�i�Y���,,�	E��:�*�#F=�=�u7�H�t�@�,�c(�Vy�9L����ŧwL��og�e�Ώzgo�fo����F7�֮.�L�r!+B�B���Zъ���I�,ɍv��=�W.�Ѕ��5T�����b����!=˂�S��UK���a�ӟ�+��$H�Q�;`'<Pb�������{n�$��F����Jù�{��*�L�gQrݑK`�.���,��ڭ��#�C�����{�o�/^y����śe��X��ʹ[P�=������/*����Y��MN��ET�[�9s��W��ఎ��ƭ��aZs�fU�r%���')׳=} ��a�{�g��<�����stK[˛"���7+r��f"��n� k�M��Υ�����\Wc���W�u��M6���\�;� ��M���u_q��=J�C�CFP��₰��c����i���W�>��.�A�bg
��5au��m���uq������Ql3[�[�Y�tEc���B�0g��4��3pz8V�����G�.�[��
���^D��kڋ�.�Qb�t�'(U����4�Ùfa�c��6,LR��%y���l	�c�k4.	��B��T�Kl4�PcX�^ۺ�b,���`?�j�=2/��lS/o����Qpzz�ٝ�*mA�մۗ������w{����M��f�%Bٓ���w-�A��U/�n,Zi=��i�iӝV�}5b@��;�ʟ<F�J�--��c������\jR�u�!9�b���1.�8T�P�+&�p�&�o��j�j��:�U����$��&�>jY�����6L�pmep'���1ӳ�n�aF<Ci�=W-�,��4���c2�b�hŬͳ�&�4����e�J��
څܳ��3%a᳡�&#�B�� 8,�Og_(Z�w;aV��8`Ҭ垚uH۸�.<`q}e��6m����"�]��S�4D�42n
�]�̽�HNuʶ=W�o�����GK�BI5K;���&�GmJ9�hdl��5���BwiU��ܠ��ɰl7yOns����t�V�զm䕵�gE-���N�F��H��FSp�E`T�Ւ��s�WS�'/Om]�������hdkw5�=j��f�&��LqJmt��(�����z�F
�R܎�7	�w����6�f�i���I4�}�b���q=�p�D����������9Zͽ��������o�l�n7n�& ���e`��>�[�:��:>}�ƀ(�v�{Q���s�E|͡C&�5.���s�1T@���	�6�^�Ύ�Q�q�GA����6�A�%_W$op_7�Pz�S3,#�""b�N��o%@;��Z�k͔$��%]�M�oذI�k��9an��u�_A�1a2����bN[��,Ǘ\+VB*E
�X��U��yvʂ+�n��z�P̾*ue���I»x̏�S6=�YMy4�O�j�]�+ *N˼��oz�JY7��ǭ�;YY=Q
�/��yyuل��V+ �28��e޼�Ȭ2��;t]]q��驴��e˛.G��Hh�+�I�����N�9ǨR�:7���OKOo��:��	k��[:i-Z���x�W_������i�19Sn�m^��������㵘���������v�7�Wa<�Ίm�T3t�4�̠����LY��R��l�k��²s�2��✒�[�CE�66�h�W�,�a:���X�\R�q�o~N��(5&�o^eB�f�G��W�&�盗\���OH�53���Ǭ�%s$o_��n-�z��ge૬���(�S�ލղ�k�I:T�����.����v߼��!Ӹ\��fD#<0�%�����䉍R}6WV�������07�yV[�Ck�zsNPh�9n+9���$�f�-]�z��Z)�G��WZ�܄)]8����k�o��姺q��t�]E��>ȑE(*�����.J�2Ө�V"f��gZ�DM(�e��Fu���:�p����]�t��h�)[��Gu2�Q"�����WeQN�,�Q9в��/F�"�bS��\�V�E[M�s��z�e�<��i���I
")��<�t9^!W4(���Q�a-:Ô���E]H]#P,�o��܏Z�I�{��&Eq2��Ќ�UW�C���tH|ݘg��8��O��$(�r�4��t�;�9���V���֔��!a,ₘ|��1VZJ���USJ0�ʨ׻��_*CJ���U�MK*��=�ú�����hA�"&t(�
�+U"O�@�j2s�o�"���*��O�+�G2��db���B��AJ�2��NU�R����Z\ͅWKrB;�F躢7��Al"A�$������薻'popy�.sj��eb��]tm��� ���ʰY�'ٴw�8��A��J�fS6�\�F>ΙU��K\�v��������j�!lo���O�۴𿐪�7�$�=*t�]���w��mS�=w�1���Ւ�D&�,p�r/i\/Gs|��ct�v�w��w�!Z(�K̥ϊi"��7�\���P"����ͺ;�KfD�ԍ�b���e�MqS��;�9W.��6��R����ɍTon�^��n'�H�n"=aＣw�����~�m���w�Ǫ=~�{
`��2!WT ���U��y��Þe��ؖ�8I��x�1�W,�|��B�8;���Wה�c�F*�],����|}����&����O7����e<b�iLP8]�V6�F�a�����w[�'�e��,]y'�S�?��/�M�g0�al��=���e�F�f�^���
{+Q�W��=�>��𵩑^��a�÷�iWcл=�]�F#Ǭh6���m�����=֤�K"�6�@Tw׋]��gVĹ���1d�x��ju���9��:kng0�v�s���M�&��A�²�c]u�6�h��ͣ�鼅G`�%
�9�*n	X�	�rFK�Dko�|E���ɽxQ�X��O#I뗦�t��z��6���S^1m���/�Ƕ#XL������C���sW��ES����h+|M$퉱���B�]c��mz�&����V�{7
�2�i�;�q�]�T�-����	�b��VNl�Q�����uvE�]����K��wg����=�߰��BP{Sle�@=}�������U/k���������C������Z���oԽ[:|A���F���(O�;w|��wc���>�)�����8��!9�nt>�RKH�C#{��!s��oYh��⹽�}ƈ��'�#e��\�޻�~!<3�A}F�W�r��kV:�z��U'�5���~���7���*z�ݯ��2���rE��cc
��v��g�3�l�W��9�~ۊys�k���;7���[x���a�.��!���GG�De[�8���X[����Վ���NJ�19B��̜>��]JE���3�I�A�N��.:ke�C!�ҍ��*f�.��;���ݸF޽ѹ�ë�v�.uJl�\��4r�.p��ܓ��Eㇻ���ӧ]hۋ[�b4�Ca��*�[o6m�������f���:�ǉ�V��P�J|���ʱ���N��	Og.�W����;9ovxe�uy���4�n��g�
�ܐ�����ﺲS�͛�e��0؋Q��틈@�U��WY��.Ϗ`�_�a���	�Dwݛ=я;"aR�Ӝ\P/'֮$��?O�|��l��F��a��9�v{�˫�8'�^�܊�!���ط�/,˲�C+�R~.Ic��S�\��=5���}�d�v���T�c8�[�\�2F=��\�������2�0db���B��_j�5
���sM���4Y��������c�f��{��=Ռ>�7ٳ;V�^�6��G*x�igKi�����'�_цV������;w�Ƿ��<	��û>�,v[vF��ds�zuV38�1K^�ӳ~X�D�R���X���Ph�y|{͓��겋uzo�s~yn��:hA6Jt�.hZc&3���6�Y�8��j�	��1Mt��A9�چ"��V�'x�rM����U�Y��fY�*`\��\9���z+Q���}���;�Pɧ��,EXF[���bE���ͅY�7��� �cϙ��1�5��-��jJ�O�qK��@����=�m	�Ȏ��~W��m�r�����>]���Ӌw����D{����������P5W�W��V�wx4��y����}^��ho�!��q:���/����Bϻ�Т@cy{c#����x�{�A�7Ľϊ��s���q{�{�k�~X!PUw��'i���5��$�_��Y~���X�9���O+����4r����M�=�GsIf炵S��w�]����`�H�UC�*v�mf���3ޭ�37Gwpц���ЕB���P� ̫@�2��'���IoE����=���ɑ+7/ha��͚�z�u	���{�X���.��~��`o��~%P���õ<e�0c�9��k��&�Ͳ}��H��Y�mD|Xy�=�Ϟ��ڃ�sd��>=������x1�5�����ƭ�k	s�W+>9�v�2>b��+��n�ɇ� y��Q��գ�<�Ofɚ�2�5c%d�;�HV��!�A��	�J�+��C*�y{>�d��h<���r�t��8��BM=u�R�:RosL�&*�`:r�>�s��v��sNS�:�ص���8��t�Q��W�&�Ho�iH�=�z(
��Bq]ó�h�>��#�� r����$O�:��Vf����Ǘ^�^��ȑA�Cc�)}��nr��m���?~��ϯ)��p���5�Ķ��
��g�0�^�Pᐓ�PK�/�Ѓ��:������;Y~�cB��%}k���u�Í�Xc�<�s[��Zu��leW_�g*|w=�/(������Z�ɤ�O5R�ځ�B�xoM6-_��߯&�v.��'�Yx���JMW����,� v���/>��E���Y�ȳi{���s��E�W?y���i]p��e��*r�wHmmÍ�"��~���P���27��X�X��T�����w�r�k��f_�v����ڌ��K�<1|H�Rq<hh����s{q����
���x�
�{ދ�=uˇtE�v�m�.��,0�h�V���5�ý�_d��/��=��u�sq�!�]�u��%��>|����F��G�9G�ރ�E�rn������Wr��^G}X�ީ�Vb;&W5GmJ�;��Fw�3$`���;�oi'�a�f�3��W O^>�tiH{Y>K���5�u�w���.I���o�T��,7WϺ{����o�'�S�],mo����x̛���e�ٻ��&���O<'��*��k���YR~õ�"7G���p^����e۷ޓᩱ�3�V��Bkb���f\8
cgp�:s}�\cja}����x�K[B�[}�?��R���� ��EZto~bV����z��^�ߺ/�٨X�{F���+n����v;6��n��R��t��ʸ7֕�����2�SL��
��ِ������j����ꬭ��r�ɖ�wӹ��^��c�m{�f��ëvl��һ���^\�.���ǗMi��|�m�^��伮=��2Xc&c$�[Y�k�>��չX7�a{/��4;�?r/�}�zw~]n�tr��
=ㆽ��+�VČ+�����{v����夁�}VS�I�p�}�>u�s��dlQ��,C{T���ER0��(���m!>'4]�YO_���kk����EB�w3/4�T� QWiq{`$��!7�&��]g�[���j�[{omI@��I��F��ٴ�`�G#������/�;����²2^�X3��n^��#�����~:���>V+oY�E�x����78����a6h�����c׾ĩLSv�u�������U#Z��޿��U'Ͻ9�C8���禎�g�g��yf�=N{B�614��1��ã�����=x��"��Na���vxU5���F,�$����8]iҷ���!��Q h��hſ�ON�>�[�ä��yw�M��jm�>��1bvա��;iM-tܬ�F��G�l{|/�W���?��sμҳug�
�rA�C�.鯁~�9�14ߠ���6����;8���V�y��cYv|{>�_�aL4�c0�ሣ3����| ���������@�����z�������F��a�.[q^[EB�&��������1�l.��e�V
�`��D]�`ny���i�Rz�s�rf��њ=�oZD/u��2���2��M���đ1p�f�7�y]u�������\��틥�b�_v*fO{��5����?W��O;N���9Y\>������|+�L�!vWA���h9��&7��:��B$G��a+m��u7E��;[�� jX���i���?>�x�=����n�{zo=�͏
Y�5��M6Bh�]�����~5�#�oӾ;�b[��Oq�u�
BOn�+�c�Nn�K���u�	��'�G�Ϻ�g���n�Ko wS|:X�����C������e�dj/�����]�+yM�5�{z�j�o�i�*4�A���`!�~붕�����T<*�w��h�\�m�>b8&��r]�z��ޏTo�L���\�^(��W��Sx�r�\}���Q���kx��{�������	oT�	��l/�;�%GZ�����ݼ�޽n���:���/ �����5�q�}�*�uA�P�֭�V��(�_��|~Z�?9�����]k^2^�f��V���y�J�'�X�J�m@���Ko�ë��M*C�v!ʧ])y��+j2��jdu��z�E}�֋^���k5���_{؀2{՟U���R�r�t����	����I�n4��[��v�e)��Pg	�@m�˘^5�:���r�9I[6����xpŽ&Re�'&�T���N��`dΑ��C�͵4��o.�D�̩��:�/Ix�Y3WI�;��!�G��BW�����iR߁�FU�D�*c|0��x.�l�S�E{���o���rv�c������s��<_Mˎ�S�	P�n�^�LZ���FLz#�L^ӞK'.t��.��>�a�,�o�3��Y�cn'�zo��Q�Ef2}F~�J䟟m㟊�����<#�Eu%Zm��fT55�bw����x����F�k�<b����;Ϭ}�G�h�\��g�N}�׮��Y��
�maބ���r(>�&0JvB��Q�M�
i�Q�=
B��r7�����§��_цU��(!�%�Ǌ��������ג�X0������_��';��lw�\6dd1�n�gn<�`ꆸ��aV��αG#��ׄZ����Yo�'�9���x�vp6͹�G�{�2�w&v{�e��.�����������7�uc=��;bc���6�]���y�.hZ��o�53���W��(c�&4��Fn��ف���i�F���5~c�-�:��*��x"!
���總��Vk��8�.��ɇ5��[���Pj��jq;)lMVޝ�OЛ���s�1^)\B��n<��ɥ�s�JF�����K�	񩓼ۋ����a�G�d8��"�Ͻ��ٞ8�sܻ$���
@A*G��6�����ʧ������z^繟�Rح˘������䢈T!q::%�w�����Q�;�tD��1�\� ����������Z-o��"@�%CCt=V������z~4�H�NJ���r��_^y��	�}��w�w�ў������q�7�m��W���Տ;������\<ߘ-����FU��3�J��|m3>���4�ƶ�,{���s�۶{՗��`�
��[)��m��Z&����ݓV+u�|u�Wq#���z����z��wù��a�����#�&l�eT��
�9������<���Gh���Mvk�8��k	���$/��VO���>ӋG��V�׎^��`�H��9@؊i��p_vv��cky���b�jG��2��5o^�@�	�M#�Љs�>Mf�t�)�*�|7kt�z".>$�د�N���
Q!ۼ��5��ӆ����J5��b�.ϫo�-��7�[/VS��\�ފPtT%pT��4�^f-Tju�p'x�����g����� V��ӎTQP=Vk/0M�2���v:��ɶ�n�0S=;��;�=�^����ؾY�\k��Μ]ҡ�'0k��"=�EA/Z�x��Bv�݊�0��t�����A��32��*�Ql�����.�p��`�M��������!܅m	�*��+��'
5��!PJӴ�ﭬ�����F,s��:C�Ȳ�6��8e����{S��9&������]p(�R���v���xѻj���|���8��f�^8h�,�F~pT�p�
H^�P�.�<�{R�ؚ�˱�r[2�Б���t��MmD�,�_F)���
��g�w\jR�X��F�N��x:h��ލ��GM2�S��;�SU�����qnX�5�3u8#m;X#�}bn])X�Xi,��p٬ںp�;C�^~�G��S��Խj��{�����
 �xU��1H�s�NV�ʍ���/�̥x뫕�F>�� ���ci�݀���M7��>;u�P|�q:T6��z��G��ԖMwC);�6V�����y��3�%;}9���q\��f[zB�w���r[V,;{��1(�7l����dJ��+59��ٸ^��jP���0�\�w�2ﭮ76�\�O��RS�ߛU�$��œ|���jf=Yo�'�d�bf�g�wt���sz&(P]//��p�	��i�|�X/�CV�/^���[�n�9H9n�#�P��³�뾸�^��N\yOJ6�����$�b�����j�JM�R�E*�n&�M88��c�C����۴��j
����ɜWa,2�ZCu��=���]��7)*#��5[gRݽ�,�����9�S˾CP��V�:X���^��vFF��q�+����Gz�*�&���̸�+a����f�Z(��=0�Q:�:�g��!@A�V��u�}�>sl�Q�gz�0Dj�ۜ�Z�v�b@�EA��t��s�Ӳ���xJ�Y[ =��V���������� ��mQ,��2�-�(�8�q���7��^�)5i�+�"�r'�uy�������� ¼a��Y[x�b�]YMᠻ7����Q�b�q���F�Űn.�`����u�s�J���e�j�g&��o�ޑ�Y$�oCVF�rV�5#%!.�o������al��3K��j�(��{�+ι�x��Z�d��rk���͇���/,^��z�͙B���L�XS\�v�b�L�r�˶_VW^��'X�ɳ�U��vА<���2gG�����F�;�l���K����lG��s���c�B�㤈���T+O�
���e���`�+��T�(Q�Ɏcu5٘���N�������Oم�u�TݪJ����q4BԢ�E(���崪�1R��:̢	"�U��^�A��i���+G��">y^*��s�ww\�T��'���]�I���{��J�w��f=ǻ޽�Y�;uJUE�tD�\#a��P�T�-����#�z��T�����s�^�zUEE玹�t��q�jj��g��;����u���{�<4���
�J��qh�9-YdV*/�܇��'��������Nk�'>t�z��/%�#2=S�Q$�$��|W}ݸ��ɸ=�4$��Ϊ^)*��G�SZFeh��s�1O�D�U�{�y�}��JN瑎����5q����,#��R���ȝK޹z>[�Xj�p�(��o�s���+6�����fc�8�n��h�%!�}B�z�sY��q�V�g�rSP�Rکnc����<<m��b�g����+����N?�I��4��Z}Q�;�.8�jo#�����t��}���$��e������s�;"��#w��)h��Y�L�P�2�T�e	l1%��q�������xy|vX~S]��ΗȈ�V��!/+=顣!6'ރ�s<�
΅��G_z������#�|��{_?l��m�u���z���>w�5]�sE�J��Ջ�]�ח�w���{V6�>�|��v��wb�J	��5Աs(�<=�w\����+Z/���Q#|</w��:�u^�j�a3�֊�Ɂ�$y�z�H7��z�̩�v��#VNuJ�W�/]k�)z�7d>�����d\kd�Gc��n�9�芧U}����`����x�%ا��p�ӥoK���u����ӱ��s>���un���s��i<���%���oìj��%4�`q���
�0_U.]�I������XC��rٰ1��uP�b}�m
�wIYB�+�hV�����2Ϲ�7J�fnյ{�ou}%`����#�n�m�ʆ�FXXYw�.��Rgp�O�PqӬ��u����`,3����ٛMo3}\�$}�,Y�y+k4��֘�8�K՝�a:Y �mڬ��z���h��o��[��S{�Ŀ��}�����#�R�Ij���o��Ͱ���(�3O�˭[<�'l�|^���U�Č��Va��:�tn�ڷft_uV�������K��MlZ�@�ʿ(�y�Q�eW�ݪ`.��~��ʟ6+u�$�YԵ_2�@���Vf��:�A��n{�t!���=�}vE!�h��ۍm�SM��w��D��v7�/��$��XcJ���d��>>�^o��;�mp}�z�Y�M.��q���:k�q���l���vWw1�{߼2~C��J}{hwySX�}�m��[���T���QQe�Q�	�ЗOO�oc�#�] ��x>���{/���ٟj�����
k����������OH|��eЊ�BȀ�_N��iۯT����N\�r�P;�'�K����lq���z�������BSpg��Җ@�����S*���Xy���U�tƽt9߻�E�u��F��i���]��ت�f�w�ƕK�@ΰԽ�q�leŖ���v�����Rc|rGd��Ǵf[@Y�;(<���S����[�6%*�S����x6�������k�z�.��v���m[j�֌*�-��-�w�˲d8~���9�=��Z�?9���^�����I۫p[cn�'+�w�,q��4����]������ȥh0�?*��9��{�c���`�S�yΕ���h���U[@\z�i�?�Z��lx=z���ݗF������«�!�l_%4��O3��7��n>-���јK���z!uMU�=�.��y�	@�����^x��������N���w��������※�X*���}�y0��ȼ�;fV�,��=�y�Ex���a�Y!}�J��:�3�z����w6��ղ�e�9^.��#�F�<����>ػ� ��a4V��F�X�b�����ýT�.n����j.�s�L���/�c��Pk��=b��6{������y@_�\p�G��}Ns|�8X�$��.'aй]ZI��ֈ[���(X�ʥ`3k�y�lr��'h꣠��H[�D 6��1��[����z3��޽��$�n|�Cw{l�=A�-�4��ՉsDi�A�D��s}��le!���G���&7���=�ǘ����g�z{��P�^v6$ k�h�Oaz�Z
ϼtɻ1Gj��v{��M|����-<֟�t��r��bc��b���#LM�����^����~R��{x�i���~��A�����1���_��En����Uo�|~�zRj�����i�J���*��S/ʞ{��[j�z��]����ꁮ��׵Z��n���� &��/�>vg��`�[�k7��|%/n���R�>��(��i��o�����s��:+������Ҥ�������ϡ�n^����q_ް��Q���G�1��+>��ۭ�c%�n��u�_��1�G�^�~Q*��v:6�+���^~�=��݇�W��&���:}���m�LĹ�^y���W��0e�.���y�b��(N�%��S_.����͸y:�]I��YY�-m���$dC��!���o]�':�[�p��O3t:���곢M�qvq��X���tj�����q����cN�Sw�2�hwM��&%Z�Q��v�U��'Nq�~x���B4��`���ب�/�H�'۟]�_�՗��y���l��:���bm�d�b��3��.��c+�$�'Z6�qz�4~�V���P~!&H��xwP������7>�g�{� �2�3_\�D[B�f�q�藘#�7{Tx���:1������C�v�_J�0�)����2�o=c(K��I(�	-k`�x_��F�G�i.N߃i���P�2�`��+v�OFnF{f{��_�\=ad>�)���|�m���yx�C0*U�.��vL���){���'Bw��ޗ��n6��/�z���í�n�
c�����ig�����3��CU���y}�u��c�#9�Q�:��LX"�^��=�"n�-K��s��l@S�%�]���o�?�6����<�
;:�"�ܼMn���UI�l{n�h�Ƌ�old[e�hGo�h�;��\�D���c�ꧏ9v�C�����%�#��`���L�?+[6N��Yn�>�{�y�u�̙�,��(4�Y�0�YY�#�EY�e�*��4����$�.�����a\Fz�YG�|ߗjJ�s���(W8s	0nt��}��CY�IInj���/>^_ʞ��{���"�$|kd4v"�
^�t��5��j<�Z�/w���1�a�m�k�S��|�.NW�������Fz������-y��E�<=1<x���`�X�X]\,��%B�堧�쑙5#]����M���o����u<W�1P����>k7U�!V;��לI�=�w���;øA���)2����*���k��;���l.IkP�g2�[��*����^�p9K5�q�Y��_=��kpGB���R����w]��wH�AXX�������G����������׽ۗu��מ�@��kˇ0�O�:�W̐��4,��z �jqqB�m��B��pw�/q
�lF��4�i�ҹ���t���V*i3ޏw^�=��[�[{h;�B�7i�����:���B_�6������ѧ�m-����|_U��GW`7����Z͞��\����5��[��̄�7�;˶(Z�uˊ�I;LRt�k�P
�["��gk7�vEy��T�0�6���pճ�	�7"��g@� .�5���զ�ղ���,�B�r��:Vp�PE�S6��/��=~,����wҥ,�>�T�9�M뚏�
���6�}�$�\kv��l.�����bx>���{�5q���L�5흚�-��������Xz]�P$w��f�	׼�ߝi�V�(��I������^z׻ǹs/uS�o�z�o�x!��9�Βs��np�o�Q�~�ԭ�#�]?X����qym�|GZ0�"p�8ͱ�#������Aġ�_Hޡ9=�˖��s�������[�-VNr�TufbHA���k�<�5��Po@���n>IR�_7"�e�Ѱ}yg���N��Զ���*����~ֳ�t��py!�r��x�N�nJ;�lkJh/Cf糣U_1���E��#}�8�e��n�풒�9{�l+ˆ��
 ��͍��0���ly^hk���o��@��� ��~�7G
{�.�ē5���0�0E܏1�tR->8��+�;�ݮ��p4�z����'4�Z�u��wg_E��d<�����wG(�?Gί���5c�����;����6$��[C�qbQN������}(
t�v9Ǆ�8�*�b�a����oq�z���i�]�;7ڛ�<�w��g���,�W����T]WE����kRv�#�����[B�]�3����*|��[���Z�?h+�|w��_2�F}�e��	l{��_y�������f�^r��f�P��������$����f&�?\�<%����$���;s�`��?����Z��1���|jz{����2�c��Zzt�w��ݕ7�[꾧�k����.���z�=�O>��`?n��}��"�����{̥G	z���_jܼ���=����c���+Zi=����|�7�����efz�U��x���̆X3�t*�\��v��'䚢��yn�X����}ʋ(\݋�swz�2�(%Bu!�X۽d�}<W�s|SHרA���s6�`�\��/{��l��X��"��ǇHc�5�c}���S��{L�kI���+2����9|��1*���bS z�4e��u��Uކrߧ�
:1�vc�8�@Vd׻����w�2ͮ�01�Bn�λn>��Q3G[��CǺ��
�s��L���b���"V	���8�Ѳ�k��8�E\a��,铯�I���q����~�}6���׼V�+�����a��^;׈p�Q��v^���	��|��'e�N�j��*��"@ن;��]��x���_GWM��ŵ������ѽ�n�&ŧ�t���]��c3�dGB������;�0e�%5Ϩ�df&�y"xŴ��/<����wV}��'zv{Ϝ����M��C�T��WWoz���ذ0��o�W{��m��R��2��3���یj��`k}^�X-�dW�{�y�#&�qz�/-�����^�W��y��=t2�2D����hvk~������ک�>Z��mፎV��5l�j���5�9(+��t�,�՝$���ں��3w�z��XΎˆ��܇&Y�H���2�;���P�v�ч���ޘ<���{��vyM�m��|�m�K_,^L|/�ܜƿ����+%e��b�`eaZ��̂ �ff�	ff��ʗw}
pl��Z�uN�Z%��Ǔ�'q
J��ժ�t�|�uΧ2�G]՚�4Р�'K*P����; \U�J��Ӯe
]9�GF^��i�=2���+��9�c��ZG��ea[��մ��-����R�e	�k�{�J���n�܋���Զy���Sݩ�g�ζ�s���ǘ#3�:�(j��o��y|Gy�c���ػ��Y�5F�)Dp/>�vzk�07#�����S���h��b�j�3���n�W���j����-� ��Fӯ���`H��Cz���؎�y|�g�h����]�/��:~T�(��[��%�lo����h
l��2���n�X6���.��[c��ך�M�p�ӥa�w�CӃH��U��4L��v(dw��O�m7�t����X�/r	7mP���q�4Ϟ��#��<�D�u��dզF��\߳�z�Ԟ�Z���_�Ԩe��.�e�����L��V�Ƴ��w��|#E�D丘��{�4j��}��6{�%h{��#�W��QV�$���#� ����>�W�և����c���66�۟�h`o�o�?��v0�����8�_h/�~��� � ��1�s��0�� �6 s� 9� }���Y��g  ����[��l�6�;��m��m�� ��l���9�m�� ���w��m��m����r  �6�96�g!���6�96�g!�ۭݶ���g!���6�96�g  v�l��m���g;m�rm�609��g8�l�� �cm�� 9��v�l�6�9�m���l�����m�� !��ɶ�9��@ ��g;m�rc`��d6C���m�{�0��k���\{��O˻���� e6�l9� f.Pbņ� ~������?����o������&���d߸�����4�C�_� �������/������0cm������������66߇�	� 9� ���������G��� #���lo��?�p�~M�1`?��f���a�?���oϰ�bP��[G� _�?���a�p9�TĀ#������o����_�  ���[������`�a�� p� 0V�m�;gm��!�m��0x@�6��c 9 8�l�x���=��N�/��� cm��� )�� ~6~�� ����~��Ȑ��?1��}��A���������s����m��������7��Gw�M�h����?�}������� ��1��?�D���3f��鈟��`� ���������G���u 6��>���������1�3��o�y��f�37��?�Q��~����o���c����~��?����#�?`��<�����O��~�~�8?`?lm�������1��������3~����ɀ�Z�?��n>�������~M�������<o�?X���@�,����|����Scl����q�i������f����@<=������0 �������G� �X~.���/�Y�7�� ?و$�A��|3f�Y��X�@Ƀ�	p@n?��D��߹��L�>����!����}�߃ �0fo�5�~���~`m�0`�3�a0[�0�
S�Sw��}��n��(+$�k19�q@Jm�0
 ��d��H�{�U	��!JT����()I"J�� ��P�$��DEJ�);D��HQZ4��X���(���"� �%Q*�BUTU!
�P�(�(Q()I*�"B�R��)UT ���
�Q%���@vj�R%(��$PUR*��
D�
Au��R�*��
�R��EU*�	 B��*����%BT��B)v�*�A�   ��i��r0jF��:t
֝��446��r]@h*�h;�j��Wl���ha5Z�Y��t�tU���B
%��JR�H@^   ns��#֝�٭e��2���QBDH�m6f8��j�zӦ���W���֝�W��m66��6ն�5�ܫ�l�M5��ݺ�uJݬ��f��1MӡӦ��V˸dwk��0�r�k2���!T�*E
T���  �x�l�\�I�-�B�����T��k)��Rm�]-�q�����V
*�-m��ŕ���[e6�wA[�ɭL�!
R��D%QT�R;�  熁��ӭ��SF�[e���5�V�S�۷w.�:)�t4I̛A���j��歴�*�bV�ev�d6S I�PQ*$�HP�  �A@k� cSh�U�h1@ �7�m�+iV  e�J��Z�p�5U��
֕a� խ*UUR(�IJw�  �� �XV�-�ڍ@PR�cKa��⚔PTm �u6�@4F)L�X PTkd ��ERAT�B "���  �y��� Vj*�����Z�a��`1��*͈��h̫ ٌL�e�@ 6"��)Dzd�TU$�&�  �A@  j  �0  Q�  ��� &�t C�V �aL� LX  T*��@�:�!�  c� l��  &&@%	@ ��u�� ; ZH  	�� l hR�F U�2)t4TU@�)u�*���  J ��@hU�  �0  �  R�  �@ �` iA�0 �V��)���* @S�0��� �)�jzj5  S�A)R� dh a	�*S@� 	2�mU$  1#!�����0�����81�: �$�&�%���j�o�=�f��i�#-1��	 �O�ׯ����6߆��6?�`�1��v��cm�f�g�����y�_�������sE���[[�`��d)e�v���MŋH��Z�PdV����
��k Z�B~���$�m,@�5k.6���j�5�(�;@ly��ok�ʕ2L���H��%�$V�Ǣ�A��!!bS�f���r�B@�]
���jM��C���5B*Z�V�Zz��j�O�����L�1��%�SQK���S@ѷ[�˽�%��Ne��թPV�v\�	,Sdi�N���XN	�C��(5�-��+c�eko00>7�3HSn`0|U�5'��%��T�bq�F�8]��i�������EV.��XqmK���@M�әd�[!iۨr�4�59sE� ��ܩ�u��5�E�Iq�u17����B��4%{w�������R�dJ�-I3j�+ ��Z�3���'2��
���*hm-�&�&F�����l�����y[t�&�l;N�:�y:+���9��w��Z����ZH]̢����n�潥�H%�&S�U,ڳ�TwaX�k/Ke�&s���܉kH�v0�e
�	!5����)����v�m�K����|��);�&��毐�qe-��)�6�)h�r����X�iF�4���"���mW@��OF�̺P�6Gn�(�Z��{��S4Vm�h�H�_Ak�E��[iV�-Q�f21ue�ѷ���5�c\(�T�mV�ɛP7�<#u+Xq�wqK�\8�LL�\L�Q�+TbZ�f��������v�!`8��e��ܢ�(aEQY�D��iՒU4m�x��K��X�8[��lT�K�r��Z��ZbS8�aɺDY��3XiցLi�j�~Օj�wO�ؒ)e��Q@��l}��5	+&�Bÿ���V��X�V�k����v�>[)�d	1JMZ��
�qm��/�+i[1��P�1�&	�@�iDi��rĒ���n�
9ZfmK�B�կp:�Y�oBQ2�ϕӴ�8#,�J���:�.�2۬IE��B�P�*�N�$��I<;�[�V�E���ú4�T�i�ҡ޷�ch�����Yb���j-:U�2+�)�9��mp5Ot�偸p�Dp�p3W�l�`�v�7F��Kd��jք�h�[�Sw`�Ա��C��ݪ�4�`1U�B��L7G+8�7Mm��*��W�|�V]KF�z�i�T*]`��ڦ��̚I�	ԖJ���j;@�͎��̶2��WLY%���4��84f��x�<�ŧcuA��4�é4.f$�T�`����fV��*�'.$����Wj���R�owؔtИӪ�i�%cCd����/���1\hSߘ�ӗ8���I±�6u��Ƽ����n�a�����$�r-�0�uk%5���hG�.�qXu��5-E�sN�0�n-��#2��&͎%��U��.��Ĭ�*��5�(n�3N���(��Ō�2��m0�즶fB�L��R��1_:�<�w��U���u{H���%�5��u"qۉݍ`KM�ݲ*&��YKtKA=Y�m|����(���t_\�U\��ٺͩ���FXn�ײG ���49��1r���+^�"�
/b�x!��9&�&�Dc�v�\b�k�����..�mij���e�B�����CA��I��b���㲅;� +Pڽ��R�H$��P���*!/2� ������
T���B��e�Z�كN3�� � ����	�r�5gN�f������b��e�v�x�×LArk^7��ң�Ee�B�2f��<��Q�єB�y�Ի���E�m];�*��fY۬�Ś��:ki�IG�kpf��U��k(�"w�`�B�۩���4Y��r�eJݸ�CMF��I��I���N^�ɹ0��e*	`�E]K7w���"�UlX���id��d�˙"������a���"��i���1S#6Q��o.������9v�FiV��0c��؍n�l�j���ڒ��VP���BY��c�[u�&FQ��zASq������!̩�F�HUY:�nӬ���!,5��gu*�Kyb�#͖�1�n��0�$�iV�P�5)1j�IzhX@\i�(�8�3�l�#ܽ�aԩv�6�H*� fJʐ�p;5pf�D')�i�d�I$-A�2�X[������H�P+�-�Tr�PNk	�(���H�b�v�r:���6��{�/m�,���NG�˵�T�S�,Ԁ�^���߰,ڰ�.�O�@ŋT���3��4%�t�m1Z���KF��dѧO�"�S&���7{��H=��.���%L�cwh�����	l�3��SwnG)�r8�����P���n�����!xd��L�l�U��&�˩Q��m+-® C�[B�)6��l�ɩ+o3J��`y��!]f4���(^b%�_��vݒ�j]�����K�����ȩV3S�o4:j���u�����A��A�w������/C1����֯vY�>'T�:M��(j��h�VY.7nm�zr�sc:��'r��W5bX�sX7��B�:Rdn72e8^<��+d,
Gem�ཆ������:0�\J1K��+��*0C-�R�V���7,ʑ2F2���h䡧E��H�@�O���w�ei1m��Ȇ��X��aZ��t�o*+�DQv�J�[۶���kԆ<�����c

�����۹��,)5�R��jN��ZҶM�[w/�0��45��1R�1JƧ�{���'I����	^�e�.�`��`���]�G7FGR,T����u%e������i�5zi�y �b�=])��.��plV�:Z6��{��4"F���EG�!-��[*4����@875�Cj6���т�Ň(\��V���wi�uy�9�kl�9Qm!r="�TP��wX�6�G-�[��ܶi1meL��RS/1�s@Ϳ��̡FE&l����R��]��k� �E�7FLn������e�biGY�S�����r�o4�A|��P�LU��wAyj�J��.�����Y��i���0���
-���y�~�&���p���&&�`��*U�Ϊ��ѭ�h,�R��M�j�[��i��
Pl�R�)�jY������*�O,*����q�`�[F���.�V�v� 	A����1���zv�wkӦ�7cT:�ŵ
ׂ̼�.0n�є�X���.=��awa��[��K2[�og�9F��� �i�Tjh[F�b|��/�,Xj��WH'Jfr1}�u����� .���b�]]bƞ; ��eܔ��a�`��ay
jlZ&n#�m�)�-͎�ؕ��&�M�ʊ��Ҥ���jA]($u�����La��j]R��.U����Ԕ�*fZ�����ةfВ��S-f�O0�#�ލ���u�����6dZ͡�gn���z��5�Ɋ,(⺖����d���wn�Q#�{*ݍR�nE��a�aQf���+a��Z��ܸ3Sx�I��ӳ(�m!�,�����c�퉹/�	j�\�B���l��36�����-�*�D�+n�[�~��*�P�n�l��x�!�b��1d�`Nnݺ��B���dLڲv��S.��;0�ۍ�	-�l��e&���hÍCz�.�FU��OsC%	����
��raF����:��ksH!`�Å�"];Ax*Z2�l�r�ٸ(����7q�(�r�Ğb�z�)�2bmQ�MЫ:6K�CX�_�Q1��SPUu��=
�Mk�Wf�B	��$�"+F*�:`���Y��n�)^�Ъ�)�X�WGs�N�v<Y�����2T+b��9B#�?�d�&f����7AO�e�0��[���2�-Xv�y6�ƨ��"����f�zR��I�t�0`I��D5E��Y[ȲeZ��E�;Y��e�9Bm�nV�lQW6͂��5��l��[P���W��.ѳ�N��G�b�36�4{�Emɑ�[3Fn�b��QՅ�I^T0�����i�ҡ�؎����S���@���`U��5�yO��G ��
�qӦ�Q�ChܺF4N�� ��@֨(7PBP�yR**�&vַ���n�^�e��V�R��OM��P=!���wp����lf��3�Y�!c0R�HҹSu*w�<���^�#�e���2���*M�Hn������mL&U����w:n�o�>��WM-�aԄn=�v���v���jՇͱ�۽*�g�ES)d��=��At�Cg��
°FKv�kDT�*��-U�	Э�wx�ZQ�U�*���m*�۫܍<�i^�,3qZ�6Q�=��MڳY�&�^lV���k g*".�1�Q��an0\�*l�B@�5qd��`�]i�����>w\��έ	Rif�n�4��љ��·k�D��YL^E3\�d+������]Z�o^ Q:���
f���/��Ԡ*U���!�K:@nS7�u�1+L$��e��b�7{�8+0%�����o#��<���h-��/*��p��$T0U�>H]��pi��
��N`v��nݛx��]Ұ4��cY�X���(�w#�]dQ�6�]�Wjb��5h�S��*��!�*�5{�ʶkd2����@j��yM-��4�R��7+P��s.��z�7��N%���'%	{e�p@�'R�l�l�{�$����.�e�1����L�K[f�ɦrGH�ĳCM�$����Ŕ�&�6�cn�͈�Җ��Y�vf,$�t�EVքo*S�Ú
-�ii�gocU�0�t�"�:����O-���o!������⑸��2��T��u
��b�3_�7l�ŗy��8k)��XRM�,Ƙ�&R��D��mM��`�BdB
�]��aa�r���+5�Y8pj��%4j�i:A6�A�Ō�;R\ŉ�1���J[i�؆��(�{�]̺Uo)�[B
��u'��ldLCwd�Z�rRm4(�PE�5��-P&�,�A�Ke*���9%*�iRǛ��1^)�����!���X)�fF%8M۔=5sA��*�Ks�"ڹXkZj޽nw�[Y�����#$����ڤ�S |d�q�jFIj�u9�7e��JR��ȷFVTuf�<�i��5v�a�6>� m�(
�45Q��Ҡ�f�NMd���XI�k	0Y-r�qm��
8�����WP�۬���)�%@�5�@m+��6����J!�T��I��0-��e� #����4EL���1����95%X�L�op\�^j1����V�E[��[�~��Rn�;'��L�"(�Q�e���TJ�и�l�r��7SsF`�4�ԑ�3p@T��E��F\҈o�/
t\Ɍ���T��㕶N]GkJ�hJ��vH�O4���\YKoRA̖�)[�,-�7�52$(�U�d���Kq�N�yn .�ز^�j�3*�+h�ͬՁ�1���1�qC�b3r6��Ŵ�j��		Th�S3r�L���JV�_EI���-�o�*���v��CH[KU����d�h�V�K܂n[���4��[����v�*
leIq�X���@:�[��;w[��"ƿ�Zrb�m[Sl�p&�p����[B�R�s��x��:-vb��p=6Ѣ�6�ƁN�����SF�E�C)���n�v��د��&��h��6��+uf^�o���GiF�POn�*�qun�-��;��Ի�mm'%���_h�p�U�Om���Φ��j1�N�� ��ڷ/\G��] �<�]`�i��㣻�h!&��æ��m�r\�b:2� oF�����[�=�,mM%�4Ȋ��rZj�,XK������328�Fӫ$��tV��XL�w�p���)OB3����Z�7p�Q� �ϰ}�j)�[$ ]܋Vr p�¦�b���O�M�l�ڛJ�
����Tlb̇,���8�
�[���$��6�-��ÛQn�Ebu��+�G1}�^͊�JX#țǙ���̦E�a(�^��S��Av��g]0^�v6�ƕ7YX]n��f�����j�v��� 6�[+����sN캽��V��n��V�qۇ�E��Cl&�Ӵ��4jF3����(���ˌ���L�-���2��7�s_��dU��nIR��3fн�'{��
�(j�0@�Sœ+Y�qk�w[��-�[�y5�u��ФP�ˤV�dܲ��l�>�!�g(<"����M���l76�j3d��nA�f!rZЅX�	���VݝKf�X�� (V���'��$���l�:�6��;y	��tP/Juq����pZh13�C�5��dZ�ؗ�Z��XZ�^QFQn1lÁ\�t�1�Z`,7X�;8Ő��PF��k+����r˼2h�)k�S�B���{u�o���zU���Xڜo&�Ryp�cn� �ᗒ�^+����bT{i*m�h#P��KE�0Ǵ����9i��h+��tH
x;4tҥo�0�چ����bSU�Z,�0̤�;��L-�iQ��Ǵ�X&��R�N�gw-���aA�i;6e"T��m]�y�QA����/죬J�l�h�Aif]iJv�WR�K�W�
1ї���W�͇�B)�e�%�ԏ^�j�hr 
k5N��Z:5�]کa�0TYĀ�-��q�a���B��mR@�{2X�!�ҋH{�Z��0m�E��2*�]�Ol�ZWy��6�Cn��8�Ш����K)�_�)6�[������S9��\Ws��(����jⓆý����ԨJ*0xٛ��!Ny�LHj"Z��8�n��0���v��}�g�D�����{�gB�F'�L�5����o���#��z��f=���$�����@i�/4�.R[ӳA��-;4Wص.�o�r�O�V�j�4�ܫ�q�=��I'�Q��)o;�<���u��2Cbr ۬
�N�xY<Jպ���#C��9KZ�ix7ge�,�t�Y����-��nBz��/��D++ uϜ��OMbneY:��V�{r3ՔG"���[|xdg�8�F4Go{᛼�����]ݴ�#{+;����[Z_%r�ү�ۢZ���/p��k6nt��9�p�ΜZ�7���a��Q��]�s�[/ǋ��~w]k�5ӣC]�h�.��P&�E��4���+�[�H���]X��]ն�[�K,|S�x�h�
��6ݡ6-�:u̙�œ��Ƃ��8#�n&p��9G�g�+jQ̣[On�n3��1v��Nwvu�t�H#���
�G��(gFsq��(3�>��"[�W[�y}݁� ��n�ٵ1鏷E���]�Stt�	���]:��MX�6���i�������o�1W3f�v�I��R�c�t2��KvV��:�o:�ц�7��]�o1ӓB���uv����1�v�+�a�]w�I���O:�ewj*5M��Ru�U��N��:��zM�t�hܥ���%{Sm*�ЃV��`��ɐ�(��ׁV5���S��ŭ���x1�����bs��83U4�1�1;��Q]i�����4�My³u�ZN�u�V�����s���-�.��<��{���}��^H���z��ފSwnܸ�)� <���B��%��߬W��]9u��՗
LpW��v�z}���i_j����O��XY�í��ΫK^c�7]���@���L7CF�é�����2'w�|N��(�N�nf�ݸ�Mm.[}W�5]X��+��,�wyIe=0��ٲP՛�C)ݬ��g2�@�S�I�X]	YmV��s�2�w�hJ.�!i�v_}��Q�h<�m]l:�����+���]��ׇ��@ŕt�sa٣�gih	l�m��ò�F.׹w��h�؍�sj���B�Fp�U��w'ت�V"�J�),��Aŉ���oi֣�J4��j��,)c�R��8��{��T��זWR啮X%[;î�j*�K"��X�!��W;����H=�j�q�z�� ���\V>�Ԫ젙���5t�n�Mó.-+Ey���%j�E��-�E���sMǪ��H�q��L�3��g�.�Xݖ��9s��v�^8(vn�N�^�19	%�W=Nr;ɺ.pǭsG����Q`�XZ��u�ӽJ�L`�O4�k/B�h}�:�-g[,ڙ��U�TR�8�{oX�&٧^��T��ϖ�G���s�I��e��#�r�����ٖ@��Ք��1LP�t��o_	8�ӹ`j���^nq��]�݇&>=��q�j0�`�kUdǰ[��r�B��)Vh�A���z�ٛ1�{��l͘����f���Ѓ{�(�j�7N�ݜ�S3����Rokx�cF��4���4q+�ͻ�^�AӁ��[���gY�o:���́���d;�cjE�w3�yX��0��b��ݙ�X:�J�0�o	{�轨��
���i7�ce��]�>k�]桝v���=I��I��c�c.��9g�e=e����w[�ֳWmxJ���"c�Lw\�;.����J2���ؚ��XDft{l���ͥ�C/�f�9�kT1�v�Tu���k��W�ժ-�i�=y�`ɜ��Hu���Ƃ;��V��z�;4mob�g1�����Lu��`�r���{\�̃�PxЏ��d�h{�+l�IX)���֍�u'/s��
�xΥX7`�G�7���?�S��~�>����>t��ѣ�0�����g��n��_@�&�N�:�1]Z¤�Hq�qۥ<�v��gL3�T�H� )� �|��v`���y�Ǝ������*:]d��u�V%W��X�.Ӻ���4���ݥ0e�b�)��W���ڵГ!"�,-�����[��s)`��`�F�����*z�Ky757\��{im=GJJ������}Sow/jnrG;#�n]p�@J�R���L�w����.p�r�-�!oc(=��-9��։#�|�!]��OB�h�:�Z�W�>E�_U��NhU��F.w@�|�8�8엨r�j��_wNﲰ3l��r��x�CxA����7VvE���8�us�z��yZ(�����=.�ɉ򻅗�]��.��ޏ�����f��p8��p���ϴ���=���-�ѼO2xg_n���$7�7K2�:Ev��I�]ybݾ{���ce���.���5���o2����}��3�;7[|.�{U9��uaG/z0��{e�b��PQ�鵃Z�?u����}N��b`�[�-�r�+l����J��R\:�:�oU�%���+����=�a��	iњ�7�d�����*�e��,�O��AsП6Ùu�a�j;�y����K����t0��%�h*	���O���$btW����]M<�WV�p�)Hc�t���)-��iy�]�	���~�1V�����v|͜MP�h��` �%��-�[fѵ|��P�X��]���#�x!ʂ���*bH��[������d�zŅ�L�kbެ.Q�n����7�ϸ3XI�<Eb�[N�D�L�4l�8��>hՓ�^N��$�=@�Skw���c�y}`����#�U��-]�򲠊lxfpb��m�x���fK6�֞��LNkU�%�+M��z�+v-;��;�wJYMZ���Nj8�QÄi�ջ�
�Or���X�ہ$yR�IQ��^j�i��W�@������u4jY,��Ծ��_v[������dL�]�����W-�0D5��1�5&�|�Nv�k)�م"41�Ź]8ս��0�y����\�u{>+���c^��.V���z��V�:��\7-7��>�M��y��S[Q���z����[[�1�+s��t'�\d��MԺ��[�y�i�`Ӣ�	����ۗ��>W�c���['�}u����P]������V.o%�H���i����і�u�:��Y���1���ҕ[*ձ�+3�K��(�Z�2[m]f��T嘬Թ3��u����
�buw4��1"1�E�٧Ǧ�{����:�X�CP��.}�r2���/��]�a�s��b��T�ô�U�k�K�Q�].�*#5Sv��׶wk	�
o/\)�Y`!F�
�S-܀�����vK���Bt���i�*��\�$x�Y���+Q��XE�)��:�����0v�c_YHYUڪݲ�'\~9pZ���𻆝,�e��4b2�(ġ[h%��kZ��ݾ����B�Ҭ)gGfX���S�4�ۖ��W���M��j]eH������2���s�B�:�i%��2t͖�.C�A�
*.��jt�q�c�h��[W��*ʃw�v��yz��+N�IO�=ȡ�+�Z����$�w:����[�0:��K�Һ4�4�_yL�A
ެ���4⌼��KzK�N��` Jv�jh�`9��vf�@ͥO�䙛T�v��Ӻ�k1p4��}�yuь����s~�"�����+	�������,ĺ�Ҝ��3�S$MB�-����tj���᧚N%{���c�؍�Iۋ�JNۓ�M7M6@ Běg�s�y�M��W\��ɱ/��}�/No�g��t7K�EX�Q-�f�)�
�p!�"m��kf��i>c����Յ���j��]Տ���6�7�sn�n��.���p�C^� �޶j*�v�ݲ��l����w��vE�P���&���fsg�Q�ͤ1 �1.����14Nݝ��w�1�u��^���`��Vs�q����B�:�j��; 3���Y�D��Lu�+h�Ae����-��w�5�~�:�W[�)e�|�=��B�V8�=e?M[\7�] o��n�������E�S�JŜkb���C[/w�̗�q EС����SV{�Zu�mN!� Yk�.�x�|3�������͗��.orEj���^��&��)�#R�'5�����cY\��n�bL��/�X.v;�͂�ݚ���Z@����Qu���e�FuVQ�%��VfVj}h�ISa���B�b㘨ͧu4*�+fә�����%�AY$B�F[μXȶ&�J̳�Lz��:�Xyj�S��1��:k#ŢG[��}t�ˮ���!A��� A�����2��LҐt+B��ס0v�_�5f�����j�z��.�ܐ��.��/]��<�j�A�Yܶ>ަ,�D�ZD��\��[B�gd�w:���u����MӖ�լ.��Y��l��N�T�-wG�j��0Z���u����@j̻�#�xC��X=��+aU���m�4侣��˗lLk3:��]2-�}3�H��qY�{3�kj����ݗ��
ǽ��Q청��$+l폔_r�U`�A#���Cm���+�U����Ȱ	G���F��=z����;�V_g-��<��nP{�-r+��^�5�\3���Ӂu�g֊k������w�HY:%ЍՄ������eӴ��������u���k�B�<z�����vq���#WG�Of�@�ܦp/�6!v痈-���}r��J����N����1��=k�wia�����v�q�Z�y/qf\&�C@W[��Vh�����+�۶��I,f㥦�+�;�7A:�X�/�o�j��n}KQ3�P�³���vP��2�j�G��T��}A)�7M"/,�W��7M����M���OD�i2��[���>�z������ͬ8u �����f�F��k8�n����Y���i]ض��������`B^��u���W�q�.���t�E�[
`�X�*Gm���j��e��Ͳ�ZX��F�֍K#�8�p��1>��F�D�Gb�Uǲ�Sx:7LѮ�&�兲�Ԭ��r�r�'[�۹7*	,�ut[�6̸yf�6���&�a�5�BB9:�Z�s��ǳ/�l�G��o2�Ƙ�}�1 9 �Ǌ/���pk�}C[�i����7WM�rd�tx��	�WX_Z��N&�ν�,ư��p����<�aR[.:z�AS��I�=�s��_=�]�K��౧a�!Q�5�-F�$�k;.��l�v.zw]�.��q��(��:�T�oi��iI�V)rLe�33�1WS�x�zu[�{���H]�{��ɘ��}�9î��:Ҳ�kS)��Z�)���I���$4@n�>|�]����<]J��&R�O�ړ��wL��V0�����]�1:袅jn4L�n��K>x�mmBN�w��o-��0����]�p��u�5�͆��z(jhͱq:WO���B녭V#s��C��uk��,9|b�B̡�t([�ϵ\�d��k��&����j�Y��5'��6+n����0kfSQr�t��vs���],>'��]���4�[՚.�&�7�$��g@�g,ք�e�J�U��$ߍ:���qlps0Ꚗ�P�)�\$�Ʋ�����!an��ܡo]E�6I�۬�3I��m
Γ�Ӯ�<�iW��k;����1!a�4�A;�c��@�[n��,��^J汁�bqq�)^����m��]}�-;bX8�6�vχ|��!I����EN�աЭ��V-�P㺰��kR��$�+j��/;N��:G&,�Z��X�D��ؐ%.p��Γ�R�ns��8^�`�F�u䡱����e[�n� z_���ok�Z�.�^YE�0�ݜ�N�����+ L�9�v�J�E��\P�r�gS�d��Ѯ���0̦���؞���m�۬��{o��O'�w?�V�]�T;v];xy��0qX�S�� �5�2^�ce�5��v�V��wq�;	x��·j��J|��}��]M�2��uv�;YB#>H���Q��h!�Uu���j�3��4)�x3qJ;����c�T��w����=G9QK�r�ٴ�n�v'��U���:��x��C9��kL�;n�/S���4pS���w�]c���t��O�f5V�ݒfbR��+(��-k:��ԗ#L�P+E�ռ�Ѝ����J�g'*�+2(��un��{8l��k5�syV��+�M*g6���<9As�8�����8��x��P�{O���Ҫ�;S���>W�x�B�CI��Hq�����*����muw<�"��� �8Q(���Jo�1�}f����Ǚ��!�@��ؗd�;,�W�kGF�ϥ�cp�)5q�e���r���j�p㙠��+npz���>&���{A�.��(�ɇ����K%]�:3>.���r�+�Ţ{Om%O;�sc�M t�Ԓ�,�eF����a�3]�QvyY�ږ�t+z��y�.���8�,�s��Η1�WK�Re��
�\����]��������
	��0K�O.P�sw��}Xx	�e�m��7/9@�i�B�6�q}�����%t��Ć������ر�� �y�]��	�8;7ge\�D�3�hu�C�u4�G�ŲM# |��M`�{:s=M^�m���e�+D�u��5��g&��];�� �^�����T�a�Im�,����23kyM�A�z��!�뱙(�P�8z�p��]�Ӻi��-^�yƔ�MNo��koR���fN�����"����ai�ư�J�*Xx�f�q�&89����(m��t�5\�������eΫM�z�+�\z�-��}r�;,�I���R��r�U�dJFwm<�V��0�˸����@$�H�� �$�i�pF�uB�]Ek�*��6�,�V#��|�0���K�"���{Z��!��u��Sqη]��a�]�k�`�����SmU���j�n�0 F�g
쫥R������VQ�N�_j��k
���Vذ�TH�Un�A��x� 	�-�Mѽ���΃(p�^��*	��o[��������5ך�P9t�ֆ��7z�.��ll�;�;��8�6ޣ&�0=��}te�nXh�aK�
���u6 ���]�8c�]��yZh�5Zi��h�~�k�!B�5�u�Xs!Z�t�I�:E޳���t��0]v�B7k��g�S��a�a���\�Pb�v�B����`ǊA0h��'o�!]�Pw4f�(�F��ٺ3�4[�����֨
���푭��r���Eq�T7%wNr�[8K�f�n#W\�+� ^vDCi��t��`w����{�f��5�X�u�g(��ڠܫ�� �=d3��\��,u�2��&�r,�g�'n�%ϔu���X��+^M���pu Z({��)3����|��{q��0�e���򧰌�1�D�ki���s��S�o�׋~ԇl�5�r�	�xfPv3�J�}��a2���[�s�4�����ː�jʤź�:�X��1=�Ȕ�7V�ދKF��.���P��6�"t��,er�f_u�R\����
���i�Uݒ��4��a�q�]ˮ$whEmV�"�Ʋ���`�銹��݂��=�OÏRG�=�m�~�\��ŏ�Qj^Z�]up1�:un�2�20!8���a��2�.�!�e��x�4f��㾱ګ�Pa���ӫ�ah�2��'��Pծ[�8����S��@A��n�GjX��B�5�^T��z�'�+��:�:��Y����Av7�iC��T�ߖ��x����zS�EJ�mc�Gq�D��E��x�\�&E�fn3�L�+�gD�W��S�q�c�AR�w��7NLxgprz���MA�Όr�L9y����[ύ�.h�4OP��X�Z����p��f�k&�R���M;ۭ������I�\������v�����U�K��8��ƮB�XrC��#F=�Y�{�r����k1k��Zq��G�"��ٽC��V���]�����1]�G;���Ao
ݎ7�,3�s:��'�.���㒖�v��33M<�b�.f^��@��(�N2���g*���S���jy�h3�Z�웛N�ER�򗘛�ME�;o8_�:i�n�6�T�y�zS��=/.����� �Y=XZ�u���,�@U�.���ǳ^��Y	���"����V�[r�c�/������|���8�-&��Vnb������� ���A%X�n�;���.:��8��p�c��SW�0L.��`�ش'�	l1Q�K����J������5��/�;UH�E��H�8�a�RU�xj[y��M��S���KL�ܲ.�"���D�kɪ
tOJpĒ�2���_ט�}F�Rh�n��� ��HT$����A�����K�Z�9KM��:�R#�� �-ޛ��'eإi-kR��7d�y�ُn�8��gmi�<-n,dF��z��ޑ.��GJi�IP���0i݊�f�Ɏ�l+��'%`�;yp�<�3t�c[*��Z����,vA��`�h�{֎ZM��<��e8�WE�d�0��A����rൽ+mѮ���/�v+��'����^�V�6�k�k�Z�*;c;����%>MLX� �mP��&t��E��ݢX�Kk��wj�B�m��YpŬо}��]�	v�7�&=�N9����T��kNY�h��6N>�%��{p��}\�gO�Sqh�͛�������.=�r��J��t�)wewR����>�-����xmVeW���r�vSdo>��t7��>�\�c� "�<���A���)!�I9�1��L���֤U�Î�[;fB���e-U,r������4zm^��!�����u���F�z1��ܵw.n���"Q�*n:{�tt�r�T]����ݑ�)�L|( ��]y`�����;W��r^�Z6�ӥ9U�PRC��e�Z@����r��?�Q��S�ŋeu_ð́NZ�w��U���n�S,)������z�X��g�t]j��X��М7����:y'�c�S���/9[w�vGnXe���CC��.n��(ݦ(���Ԛ��W��D��QQ<����؞��I!��a!ݸ��Zn���� 5�� ��߅�Kg]@�ӭ���pO���u_]�i�,���/��x�,�V��yZ�j����PM��wj).�é1`Q�Ƿ)L�Cm�r��yWn��s���97��*���t���=�C������ ��]�5�L�=��۶�(���f���y]�D�E\�+�����칼�j��&�%���në/���J��ع���܇i�Ι%J�ڤ�	�5����Y��I.�4v�Z�����X���&�����3c�O7��(�_�y�l��G�9���b����]Ǵ��g�����f,m��g�i��ڥ��o�J��B�a49ot��1���#|K{(�*��fܮ�8bP]vt��L�d�ܮ���m��ηs�T!K�r����nYj���-EfQ]�Zܬ\����V���˕'�+Xo-�T��o TrB��s-��t��S3"�O�ZY|����e���m���-bui&�:]�9���F��Ί��J�:���K:�t��kX�yզ��&2�iDڹ��LU�l����|�n�y��짙]y��ܭQ-��]Vi�����*�NQ�2L3���3UDr{1)j��Z�{o_IV��LscK-1�pPx+�̹�l�j廫-.T�(�a�c�9�|����pf����)�<�� Χث!1��W�`Kİgun$*|�s�8����01&�Ah;����)�f3Ĩ�M4ΩW�.�V�7]��Mh�p�G�tH�׹7��eru��i4*c�O�Sw^���| �z��ʻ��fj9���q:���µ�e0��D��dI��fWi�uj�5|�����IH�K�Vr�)v��5���#�;� �G�k�Qs��ˎfZT�̻-Vܙ�r�8rXY��S:!�@�x��E��Ծ7�h9O@M��!z-֚�%O�̕3��t���)rQ�Jnةj�Յ��C(�N�#����M!�o:�]��vt�ZC�B�qs�&[�^�oa˔P=��)��O���H��Cw&���#�����4е���(8��V\������n����v�p��#g�:Ҟ�b�Geǵ��k\G����Ԭ�(�ՙO��s�O�m�� !rs����xga�5JXzi1���agΚtd=�����%���M]��b�����A�7�b�e6��}O��w�#�%�9H�f��}u�����ӆhvn2�Zʮ7����+eY�l9N�N��� �Z���,�XAZ7���W&��sU��3)��y�t��@��ˬݸ���Ƭ��l�8���1��Y�����|4G�j\�f^Jj�(tW&��X�Һz�4�wn�w��
6�n>��T���	�t��ݙH�s��Ծ���w���c9��m��Y����{N��\{�S�����-�|�R�ۻ���κ�\�t(�b���Tr��;�[�y}Oc�]ߑ����_uf��K��`�Ҹ��Uv�<� �^%�U����E�v�n�
��z�c�]�°�/gv��"�]65��Mc>��)e�x���*ɾ��ΖՋ�s�DDN�Q�W�!�t6�mWi�5W|	.gj�\�ܺ�З�٬K��O���Ԥ�T�aFkr��w���U��}�gM�S3�v�*��J���#5En�2��g��\C���M�e(P�C|s�h)��^���P��(�����枼�w��o�e5k� ��R`��p�I��U������9�pI���i��٩��L����������M"�C�9J����K?l].�圃:c�B�f�����˫��v�|��4V��i����ܺ�_ڒ�VI%��**,��K�h����=�.�U�"�FV�c�/'gs5��$uf��7ϖl���}��ClclJx��,��:���H����Gp���=6�t�G;(��7��ڭ2���mm�U����j󑃪��Dgm*C�c������H%�����i��o+l�2e[�5rZ������5/�)�'����ͦ������nىQ)i��[�ob�/w]�Fá��6�js���Ƴ�����2evu"S?eaJ_pW!5�t�I��-澬35���w'V3׽D :�'�1�\�;/t�ظ-�v�E&��ݏWt�(��!��]ҙ��ARR�³���s)��WxZ��f������X2I7��A}68��bH�w˝��(�7����n���$���l�Aq.�1�]�fE�7gfQ�0��kљ6U�V�+
AU��;���	r�
V�l��GC�GsU�Ǯ=�/!?�R� ��[�3P��u9[�1���t�zS�M���$�o�>��M�����h��e��0_b��JY�N���U�ʯ����hD�c���m�U�I-�5m�j����Dnt���2P+�>����!b*(�Z�(iZĪۚ��϶�W��0.����V��lW>��ܭf��H�P�qӕ�ia9�״C��Y�//��ۅ[׎��8k��d%oM8�!]��ܗ25ݘ�撽�n���6N2aC{)U�K*�n�ز���]�o��VD�h�d=+6�/��e�=�Br<��7�|�A #��12��a�<��I��S�gP�W�p�TN��^���ܛ��N�扢�^Ԡ�:��ec냶�[=lm�]mq"e����̣}�s�'���l%�:��fJ�{���wu*���Ƭs�	���a�tqf��du�
���)]���H�o
	E�>i�=KOZ�-����[}�9���Vۣէ)%j`S��J�K�I��L��|����GOv���󾃹�����ۆ��d��u�.��V5����oDwκ.�v��fJ��QF՗/��E��Z���Z�t���oPD�� 7C���w�����σJ;����]b,�T3��u����M+���ҸD��6��.m�B	V��i����0T�sif��T���Eʗ{�FI����X@��Ӓ�U�ao�������O/ńj�sn�Ƅ_��)۳��Ϯ�IyƖ*7g5޾�c�Uc\u]WL�*A=D��Ƕ̭{d��7t��Y���N4oY��r!��>@��"��K����\�9S`T;����Wr���:�VS�����j��[�pC���ٰ#f��x��؀�rt7�ԐR%f�9�����=��ۍ�kOӑ�.,�:�#�bM�tm��7�T�n�ȴ�X2J\(�S��6�𯃾��{���|7U�;�|����j���湟�ҡ�R�b�9)������i�&��}x)��)I��ltξHk��V���9��\k�O��U�q%��2ճ�B���սGR�]��XL),��p����ΊCvA�TIkv��ff����/�K��*r��u�nn��*>ڹյͥЛ��=�u�(��Z�=aY<"hogQ�;�Zv����Q����"݁L5�+�ҟ^�7i1���) +k�Xn�hqw�o��]X*^0�z*�i�[�*��B��u(�C�-j�������+q��C`O`b��Y��4��ݸ)u�Ǔ�2mp����ɚ�S=�{DV	/�n�3c��X�Dn���/�6��� �o�c|tl����/Q�a.�0�o,�b�S6x�e�}.�bW��&VX���\o��:1Go�c�t"��U��e#�Y[�S����s����Q/I\od]��fvEb󞻅m	�K������z;*Ӳܙs��ӺV��.z��h$�2��;NU���N�6��>j���aCۚ�-n�*�b�"�P��6�&^|Reڗ���o�R��ޤ����MV�T��^L��E��eq�F�w.]�B�o�s7N�h�]�.B���AD���"ɘfr�67�ڑ��d��*�>�G�L��I�#w�қ�����A�!M��v)BqP�˹�S9A�a=\_$/l�E������W7[X�ۮ&﶐9�MP����5mENɕ2���4�Vӣ\�Vq<�.Rѻ�F� )�Sz�����ͳز���'��F,�Y��'�{�*��i^Mq�4��:�#Y�A�Ϟ�y�,T�9�%��������*C�(JŁ�p�CE1����]�'GyY�νn�JgI�z��ռB��{h��DVۭp�)7���e�ra�$�wZ6m���]g:�Nd��W�|U��˔c��Č��W\sy�v�3b|۬� @P��7`��N���;_Y��1��k���S����Y��6�9!�L@/�v��=/Lg�NSVb�8��X��}�G�A��2��(#�:���J�T�g�4�� |�]	��/:��d��vXi���vُ0)�Ⱥ�WW�y�^#V�c�V�if<��S�1���j٣n��t�'-�Z2�����
/j]�tv�+��U�r�jh������-�f�cY���?AܹcyQw۸Z���b�.��=�3]J\�ʶ���Ʌ)zvӈ佫�eq�]�\!���TT�[�2�ғ�#�Z:͓�1O�][e���W�v뾫�e����:� �I]���n�����­tn��Tö4�_��pj�����yi�O�n
�]S��O���wg$E���$��jA��-�-WP�)
�~].ɘ/6�Y�6I�G`4o^H�t�Yǌ]L�yҥ���C2�V�j�$O�@ ���oz���4h���dɡWp�j���z�oz�<L14�|��KOu�%,��h��m�g\K/��6��]�,s��),��V\�٫q��ڴa��q����;1�s����k��Y�@��6	���L��^�-�a�-�Yu�{&)l0��yJ��i��&���j�k�X����5|:�ȕ��.[צ��X�\�Fި���Ã��S5�υ<sN��}��P�B�P���3��^�S���sY9�\���}'v�s�#s^5�Nvu9B�޽�����еa�{�'<JO�nc�i떌2���1��}y�7z��'3*ގr���\�e���+�Z�E�p��T��K����3�H6���E��SU&&4�݂K]�����#�����]����s�)`�m��y`/�e	�U��a��/'�䫭y��E=�E��ѕmf-:EoP��nL�)�;��E)]ԗ80�q�`F�ڡ����W��nюfgkUyM��]�*U�Ĥ��Ĥc�C�km�N�^�<K��-��F�!6��>�L����<�1">�9��g}�7h�ۘ�V��덌���Hb��3�ۂ�N�s ��7�e%{o9��7�왷�t���.}W�c�+V6�%�%�]��2���J����«0n
z�޽U�jV����ؑ�Mh�γvT�>t��lo�^,	4C�A��aSa4Ą"�-4�-;�蘙EA'���V)�r8U�d���u���2B����[��*ȒC	LE9j��\��(�,���XZ�W0��B!H)U�e�V�y���GD�5
�0�e$��+6G.7S�*�J�	�ȯK�zY����j����#�b7]��P���^Ij��(N�*�A,wr=LL�(5�l�S�RBL�Ee�EȊ4# 2I����̊�6�iUa������&UFʱ˧,%0�2��T!&JwĄ��D�XW"�rդt��iQ��emZAIZ�^D�r!3�3wv�438V��r��6QZ�����&QV���Vf�D,�*Z��F���
��$��3A9E%1	D9(�ҋ�UR,Ĺl.�	%M0��%i��,�j$�D��1:���<~��;'F�vj�B�μ�;\us��H�v�C�OGA�R�ӷR���b �v�q���e �+5<{<,�*߾��7v�;�_�U���Y�Bv<���R�`���7���������\��V�H��o}���3~�����8�z��C���q��H�u�9sb0\*��PY�N�yi�Wi�=�w�^V2��!0��p�
�TbᲨZ��7�*��+��޽��r�b����w��0�����{f��1`٨�(�ʃ9���^姅�vc˚w:�U>�K��:Y;�P�d0[�bͩ���f���ӫ����$r\[���ת�c��e
�YW�*���ߖ;�ddE$��p�=����7
�B�.���/�Bw��x�C� |F|o>�:��Ԛ��@%�wc�ܑK'���yLB���!`J{8�܅Z1��}1�S���n�<�!��v�7��!5�͘\9�ӽ�b��-���v�r� �n�����Y�*-d��؂1�m��jPo�k��7��f��P��<pR�=:Fޝn[ڹ�#D��}�!�,�:>c:�\ ���x�t�%#���L��|��
^=��Y4�82����� ��2﷧v,��\���QJW���	+'wS��2)`�έ�b����`^�u�t��Uy�ǍYB�)�Mk�¸t7Y�2��{�v�l�������ZMޝx�{��d�td�Ƈ�J3R���*��;u�Ӗ8`k.+��*�X�*��T�j#��ݝE)�)n�j4���c[+�"+I�|�t)�]pѐ����,n']��7PpЖ~�oa͈��f�=����S��LL�]F����� *�Z���$ա�]"b�1���Vb���{a`��8���D1��Di"�Vӣq])��>�~��}��Ĳ�s�қ5���B:���\ �������� �.�̻*�*x=��uL�8n���}u�k\�|��T_E�L�7�n��D���b:����ױ��d�2���^��tKռ�.V|%�6��0�>��эg�O'�Bv�e�+ῴ�`\������.�D���'�P�82-��&7K������B��W]{_��o��:���y��ޮ���3�����a�qUQ�@cA�� ��u\@R��N��h��$9:{pl>Fe����~�Dw,�����C�~���s2�+� L|���2��d�TC&�>��'xi��I�tH�
n�[�Y|l�RQ����� �����cԵ
o�-���do�.�Ⱦ9C1��[k���*Qۼ�hXs�1��"�t��n��ֵx!/�%n��f9.�J;J�:�p�����1���0�ac=q�;tssy��Q<�'��e��񛞞�.�C��-��!�j��ܛ똆�� '�˥`j�//3�;����KE����W�nۨ�7�rpR$��x8'Bϫj���;�ʽ��rS�\�YS"��5S��eḄ�y�WQ�bm��h<r'a�rjCu\���=:���p��F��t�y�(�+��+�1�C���0�M\>ό�?P�Z��̜)4�ؕ��YGk�|y��$jdY鄍�b����o8P�R�ki��Fp6fv%TO{-�h;��l�'�kȃ( �'"	�ef_p���*�;�ܾ9)�SI9q���W�G]>�$Kf ��S]2zi���1��[�8�}�$��4�����b�n̽�o��������Nzt������V_)�b:d�f�JF�a&��!"27��r'ohw
	{+%õ�z���qj����5��c�0��_���;�䐜haE*�J�_��嘺����t��L.���3�鋅Ҵ��D0�̘K�)�NX���7ꃀ�_�]�؛i.�����m'q��S�Zeƣe����U���=u�P���e�5�R��]��v�ړ.��C��Bڼ����#Np��;�b�r�*i}����ς��͙�;V��)��q�J��A�q����_�����ٛ�l)�)��@�0u*��7�Ǯ��9:hWx�K������q*4xK�]����{:����b�{`Y��Is�7OWk#z�тh������3*�]a�;g$��z)��H�KF$Lo]H��
%m�s�����G�ne;�f<�����V�t�u�N�J����Us.#]|�����ˏ�z*;�]GKPvd�p+��.��L��E�FN�uN(}%U��-��n!]��
�E�P�v�5l�T��W����ٹIp��K��z�=%/2m.g6gƝs�vXwf��2�P�+ �ݸU�b��`�C�䫷3H��Wwo����2�dh�����k�"��
X1üW���_P�*+$�����X����ztK���+ʨ��*���<oS�g�UZ9���b�:ꩡ%G�*nj�֯i��~L�5c)���OU�|P��\��%��Og�T�7$ױ]vV��ӷj� ��@X_غZ�ٓ���H�IvD�z���QV�_]���n��g5���A�:w�d�2w��������YQ����[u��&�#�X[9�A]R���]x�]`���Z�u���w`
�Qm�Am_#{�W<��ݙha��w�WmXt坮Ǉ�>�ŗ��] #���kQ���g�]��e��i��������R.�7���7�9:ۢ/\�2�E�q�tB���f7�}׭�Z���9ɕ��wtP�8g�<7�;l��-��0ECS�U##�<�MO�M�N�rN���r��v9RC�=}4.)*�7����k��j�/�c)�ъUHw}}7��k�k���	%?��%	X`�'*�q���A�U!��Q��T�y��)���^Zˊ��8^$~��t�8Y;_���kj�t2�̯[�I��[O���!5W&�Xz:��wpl��p��':��*�|���K'���96:��q��H�v9Lh�k=L�QΞivj�Z�m�]�ϵ�˘�?fú�ZVL��!�7(u�2~U3a��˗���0t�vǇΔr�R����gx��x�;�굕�]����iB(7��LeA�ZB����Kn^k�N���>?^A���R��ֲ�n���u6Χ47{��mR��c7.���;0F���-u��`��-:vU��4�,``O��22�w�uI��u���r���
~ǲ�݊��ڥ�S"�{�dI�Q��z�j�ug�����!�_*�%�*n`�������>�o�I�$cnC�T6�%k�>��C*5ݵrtZ'mv��Z+�ar:h5���
�D�H�_wn��w�ww��B�̋1���&��kzT�'@�u8wV��\����Tkc]
z��fU7hl��0�]l���VuP��7$TB��綜%4�ե���.��)��o��-�й�8H�+��E����'�H�ڡ�6��τ�79y��@R�.���&b�*c�&��Q	�c�ݷ�Y]�6�������qu�d^�R���n����B_*zy�>}����u�#V�^�t�9\���	�*p���Un��8�p��^�����c.��=Xၬt����ү%����!
�%���]9�7-0�n��F���� �H�4��:"���51zX��t����s8��q���`�o�]��0���1q<���Et��Tb�W`����2�D�r�<�u��M�����}�ڰ���:;�K�i��K����wh��Tm��g�=�riʒ�F���D��ySÖ �Ѝ�0�����Q1 &n���Q����|q�&}'��ܮL~��2+sK�ݷ�����Jdɴ���c4�$��WL��LxAˆ��w����ԤY/Җ
�M�8�\�U��ϖVIG.�M���C�_I}��b;鯅�fK��
��r0�������4�U	�����b�g$;kQ̠;�i���KGq�\XN�b���袜%�2��[���3-Hk��yB�p���<��gH���6��Zv��Mk��Y�ݣ��J���Bv��QЬa�*��{��rk��=�a��+;�	�FBÂ��q1{����p0����|�W]{_���a�u>2��ź�4��S�kE���LΗ�;��a��UP��(h;}���^��!6��u��S�)�Q��ۛS��;�@��v\<���Ȯ(��3j~���IL��a�&!cO$G<��Q��{
y:���)�S�}���S����S�M�'��]e�X�eS�H�����v�*�z�c�]�ҽ\(MP	��I��}�/�<*�<�B�b�؟ND�D���%��A\3t���uʍ�s&aR��ꯕ�t�l.}O ލ�]F鉷��ga�sJ�q��uoS�̖��o��6+][s�#�*Q�s&�;c������M\>�3l�訾U���sI�͉i�e�٤1p�M�Iq�@	�lB�@�~ـ�C��([�cY-_F�zh�VotI�Qw��ͮc���up.O�p(�R�&�&9��}¡k늿�;�t\F������� ���E	�_�m�G�`��UX�ow���Q��ӨN�������=P݈�̸�l��PEb�S��m5z����ɑ��wL�ZĚ��s4&D)���cc�M\Î���'/;vV��;����0A��{˞9@[3��õ�y7���1�u�Hq,@�ꐚ��=( �d>%*�cJ��I�FH���0����v'N��ꋑ�7�\�9��&�ߡ��+�PQU��3��q��;�E)/�mM��1���k(�WM�ٖ���6���&Ṏ�f�/�V ���@�	�b�Ë8�&�d����Qnܣ�Ľ�b����Ҵ��D;��Ԙ��$�ɿ���w�K�$�ڠ)��=���qO6	�Vs�b[�);U���
y^���o�9:�!L�rćò[|j��:������>�igI�P�]���??��7OW
�]Vl��,�|=�xQ=$�(��l�j��*{�:��zi�g�B�Y�m���9��|��q�iV
�+qw�4����+ξ�Kt���#o�_���j�'=u�c�0E�`ٌ���Nu��?�����d|<�� 1�*�%L�YDĊGɫ����B��Q=�k3�b�����Jg/��::�F��S�e�cf�Jy�C�L�����4�Y���R�C`}�I}�Y����c(!Uͯ�EH�D�\_g#`��*�vm��ݷ�%f�zM�P]󵝪lB�6���+� .a��9�\�
8�=X4��m�0��Z��C�o:�W@"���q<���)��D����8���Թ>���U�%. mv�J�d.�!`<)�<xH#�fҠ��sA!���LE�)�u<��ƈGP�X���*��Oh��ks��*�A�����!V�t��g�UQ��^W�yj��<B�U�Bl#��T�%+�7�vۇk,�P��>m�dJ�z�l�WB븖n=��E���o�ũ���۷<m�p�J1������W��� �RP�*a���"�g�;?fN��6;)ێr��[�q�;�U�QN��n�1�r�#�-�#/�sH�|�A�h�:יu�D�x�S�3޷����@s������z�v*vٌ6Z8\�h��UH��O9��Ӏ,����$���'�+�h]s�cqa����j�aZ�˂c)��nvQ��.��ǐ�ys�6N80���0F�'>���*㺐w�\�/�z����K��B�8!�hq���0�R��+�d�&N�2��c'_q�0�R�ێK�[	QmN.���ݎ]A"1\� �E�?�U���~�d�|�MAɱӮ�fwx,�X�����i�����j�T�e<����6���/{�Ф�Y��z㽖��\�z��_�`#ٌ%�K���x�����ͩ�;*�nKZ�f����`j/u-��v̅�\`��v�%�����9�.��<*%ud�Z�J�:�j�����Ws<�U�Nj��A1�ۛ��w�5:˜����i	��+��W��1pڳ�#��w������Gh���t�<w�e�Z��
�xXNg�]����B(=Q1�xy�˝g��}�}-mʘ���ᒛw�.<NJ�|�g���׹ׅJ�V��uc�#�8�X�U��ٵut���C��XP����ۘB��������������L�o��M���=�{������<=�S��Z�?X�tB��Ԛ�TQΨD[r@*��1Xvt�����J��[�B����b��˩��z۶�s�%���@����&stʩY���
;М�ZcD0�D=�L�åLvD�h�L_	:O({]qR���V��sw����k!�`�l�Bj+|q�,�9��6�-��	�/�P`麭����ѝ��d�{mm�r�(.sL�-�#V3��_MC�8`�k]�w�r4���>�sB���r��s�ܫ�e����PUD-$_�g��ЧD-s�C���g4���w>�>�FU���_P��Y�� $����1J�2V���{Chѡ}��p�TɾK2�ao22��Ƹ�ġ�����c�".�v����"v!�u�{��R+��u/W�A'8L�G�i�`ܱ/�T�5��N!���]1�ⰲ�:d伾�[1iHq�]�3-�6���b���"��ș�TF�$�М8��g@�]Cb�����č���R�!Ǧ�/��]���#��]O֙KH�X��y|���dst����BoY}|�K�f�:+�]�;x��R�K��F�nH��	��(p
�a'������t��%j��~CY��{�ԣ��1`���ѝ�-� �Bf�#���Alv-u��JXq_wRu�/C;I�vp�� 6uS,7�/����<�9�@ԭa����!���KU����Q#j��C B� Ѽ��/��.>��ʴ6c���:�R�U�w�S��(�c��xZጢp9��n����^�`#;����Uġ����-;�[�DL�b�Y\�d$�q Ms��̺�a
X+~�U:�9B����Y#���)
&ժ4�/y�|e��lLPk��nS���x��,q������h�4i��֣�G����J�f�����XSI'�d�u�oU7;Xz��g��P'�)[],�)m,��c��9�+��uҵ,ܭ��*�<�um � Ϯeeo�:Ue)ɭ:덊���I���k�����dh�Wp�j�7�؍m�\ŶKGw��Gø�	��e���\�x�s�/Q����H������V:�!��pu�u��'���2�6z��]i\�n�j��R��;�I�����M��MU��+f�ӵwQ7D���M�Ң�,�7� �X�ɕ�U<�%`#�:UyD�s�ڷa��t{{h�:���*Vۤ��-bIŻs[� �D����S)�Y�m��C�ڇ+�GNcNuoe-ER�ߙ�mn��"�Y��L�{��}��)'8C�� �kՀ������hsK:�������z�$�49�;3��n�oK�B�b�٥d��,�n��p�s�3H}����Y_wo���}\��Q{R�D�[i-�����	�|�b8p�6��V'���� ,5��e�A����7C6t��w�eh3(naw[1�`(���Ԩ
w7���˩T���Oe�뼡�o$���v�Be9����6ˢ��]ӵ����#��V��V�"�Zg-�����fۘ����҈��"Ş�qs-�:��0���}A�{Б�����]�n'HZ��u��J�u��V�*���=��N�X���$��tn�꼉���t�Vw^镭�.�y۱Z��̹�g�HQ�K-wa��u�z�����n�[@D����f���DZkk��|��хhm�3�a�\o��יs�}ڡYu��N� ݾT�sK�k{8�L@�E%@���
J�DZF�T��30��6+����$z�j�L0�(�:���f�hX�t�������а�G&RHQ��8TZZ�
��(� ��KjK�Ȍ��s�N]S4�Eh�Qbff��Uf�Xj�NU���g*�*YK*���Ȍ�iAt��NyD^�(��ir��s@N*[(��B�ͅ**ҋUC9�`��P����kU��U����-h)���$	K�����*��wJ��u�;��y���B��Sk5+�*Q���ኰ0wJ�,j�q�
͜T�(@��eY8PVK�NbG��Z�EAg.Jk
��ʨ�Ċ�T+wk�)Z�h�E�&�JB�#J����Z�g"�3���ueص9\(��.Q&E�		����hQ��j\�%@��)+YF�BQ���P{�����S���΅�0�HH �/jJEe�n�Uco/r\#apR3>]�<���^&�
��o=S�C t�]��^u�n��.������h�c�:��w�R��K���쿫�8q��90����"���s���Q��?P�Q��v������[V�i
�RCQ/�`J/1ȝ���a��hWw�O/#Ȗ����E֟���!�����H� G���t��	�v��x�;�[��`��O��ޓ��
o���8�G+�M��T!�D�0CFL�DR i@ΰ!C�� <����$���}s}�q-�%؁�o�y99;��O�4�B��eH)j��M����u័6��M��k���`97�$������ސ�zC��� }y���nv�}O����q�\�[�w��O�~��A[u禅$�n�ڕ�����=@|�U����C�s����zw�?�����=o�>&p��@�  P�D��!
Q0��v�'��?��,~?|Bv�����ۓ�s�o��a�s��zOa�㷤�C^�d����͎|9z/���1�p�恥�}���0� /	���� ���%��"(gޓhy<���yc��L/���׭�P�9~���޽@���C�
V��!+#�ɉ`�"+��Pzl�Mj�u�"����Dp'k�
~!ɇ�|q�һ��@�O}������~;I�o�P��;rr��J�|��eH�`��ȗ�2O��aw����[{M��]�߇�������=/㈙QX�ly���*p��>����y����zM��������Nq����ø=&w�=j�����~�����/����4S���u�����}Bt�{��{��Sx��/��m�1��D��B�I�d�]o{uOWzB�>�B R�����	F�-�byZ"U����x���_#|?����r�~�Ʌ�P��:<w�=�w�v�)����<��B�
�����>�>� ��@�7�˫���]0���7��oHHy��q�/��'&�β�?�6��ߤ�&�PadyGӏa��C�巧r�{����� ��YQ��F��G�H�>���>�"$}�{U<ᕤœ�6���қ���$JA %@B�7d�M�<���D���;��;�&>`�9�Ǔ
�������$����y�w����NOnޞw����O;rr�h���_  �P�t<���?�t7W��2��k��N�w�^�s*8��4oWs0n��hsڙҴ�f����F�ܾ��ε�T�]]���Ӛ��s��d��f��k;���"��حG}�ּ�n��(�c���g(�v��p�u�m�ճ�N�!���>��J�e�u�A`�)����}'������>�{M霻����������|=r�<q��o��������S��S���!�0����~��G�߰I���ۑ��=��JsꅿeZƬ}���:�h������L�����w���^M����Ϟ�еCj �0��A<����� i<�	țBw�j$���]��������Oڏ�� BA % �8������7!�ψ{:ސ>��p���@��(��l %r'��G��yH������H�u��~��I���Z>����d�0����h�sn^/�x�r'�s\3�	@�mB��>��ɿ}��}Oi��_���zq��97��@QC��t���Q�(C��X��!�#�2c�6��@���]��� B�ٿ��a����o�s�Z�|L���Z#�>�6����ǝ����7�����|��B~'�,{Oc�;��n��ԝ;I���O�ޏ�`���j>/ 	G��D!���&�c|:��sW�W�5�*�h��-|~ܐ�aC��z7�돨s��n��L�'��y�~'�|v�>��ޓ|Bt�lz��rz?��zv翣x�?:=�z@r����H�K@�|��Տ�
�W`��B�h�����>B�~�k;�<w!�~�z	90��~}���;�zC�yro�$�!'��8_��C���Hq'��zOo�ޔ�e ��!4N!ǭg��Ç��h�����2��*|���hR6�h@���E�H���9 ��h�:;`�F��ד}���F'x����ǧzNL/���>��>8������7�?X��~���O���iu��;0*�����=���hR��!���2cY	ZL.�C��Ѿ!ɇ����g��v"Z79r�ȜP����$��Y��y�x�}$�K4|_}'�'#�������x����H�D�봛�'���|v���������>o�ޝ�s�O�=��zL.���>g01�@��L��J���E��"y��)|�"/6��8�v�"aG�|�,h9�F���tF{fդg�ŗݰc��]�9����!,�:�$1��w�
�� %##��1y���!`�鞁��)��Σm���wuy�c�[T�>-�K6$��L�}|�*�;�&���{3�]��*WwWwW��[�4�m~�!�a��ACD_ﾫ���y��=����Q������;H����p�Ӵ��x��ӏN%q��M�99��]�1;��#��BG��>F��@B'�`�H�G�"	�^fV/V`�71m,]�d�m|~�Oȟ  �&&Hh|�7��ޓ�}�i�|����Ͼ��i�]�����Zq�����Z>DQ�zM�����&��!��=~@��#��z�ɑ�]u?f:��w�R����~�ӿ\x����7~��% ���@y|��nz#��>;rw�>���[w�}��{L*����=|��� (�ݹ]��~p�1H}�>Ž)����^���z�[���+zB~��I�\
o��z��߮��`��*"i�~\��.2�~D��dF]㴨�~����A�����<��{w���'�~��raw�~��zO�!">�|~�`]6�g.�q����#�$} �xj���L���=�c�ԝ�[�ۓ}B7��ӵ�8{߾�}AH4O(���@�|�h��y��!".�����'��ǎ%wϾq�&�����م���U�s4����3AZ���<��!�P�#(���>X�q!&�}u���7�w������ �>��H�CT�~R�T���OO@� -|Cߤ���8�h���{Kk*$�L+�a����P�5}�Ӿ;����i�o����\
o���)8�^l�)DB:�"k^�}q��9��g^�
�(�j<O�.D�YR<��6;}#������Yf�=:�稼��~^�qT?�臤©瞿=m��7��� ��Sh���R 4"qB�j&�0�k���ڸ�}�}�rw�����ӵ[x�'��	�]�>n���.�� Gկ��=S��,ښZ1�^����������￞�N�O���Ϟz7���]�>w�=c���9ΎWx��~!�G} �l�KP��A4��G���	�}v�ޓ����N�S�}��I��%����z��u�����O���H�M��~>�.I���zM�?��}Hi+} ��5@Q����:������90�v�C�ޝ㾡����Ҹ�Bq������Ѿ'������!ULQ��Y~,�~���y�ǒ ��FM�p���f�eJ�i���a���(w�t�K��{�WԹ�Z����N�+�{�F��Ea	!�G��]y�+�}JE�ӣ7��sF��ܓq���4�e>J]t��U/�6���C5�W��H�9��U�P��bN�Y��V!��}]���[u{��G��>b��[��
�X�Q�=&�$^����J4�ju��HD��F��@2�� �d�>�0� $#_vϐ? 0CBϞ���_�9�'8��8�9�?_��{g!�9����xa��>�} ��@�B��f��2��0�E�(J]�>z����&���v���F|ɎcQ0�4����h|��Ϻ|��Z�^�6I�!$@H	θ����NT�;���W)F��>�DJ?}������m���{����v���.�iP��c�}�9ߨ{�ޣ��뎣���aw|���i�������JH��k�� y�/v�� Гl�=�V�Eϡ�B"4A{���{�oNܛ��y�'Nה����7�I;~�����?����<~<�p�C�ܛ����~��S}O���!�@Ϙ!��xV@� 5�B&���Q�F�wH��w�*�=���}#�>����������h�˃� B������L �}"���J�)c'�90��w�|Oi��&�~��o�oI�߉�@�����:���7�/�"uB���^̬f�F*��|�DZ�f�@��v�z��T"!B̀�x���~|����]�w�^�h_"���H�����AC�����o�=�F�C�=��T��to�p��r7�1�-^�z�|���hď��ܾ�H�41-�R��Z�TR�o���S�^�<C��;�����<�m�@{>�B�!#�%؟�T�G�i_�{�=&�������c������v:�T��/=�t}3q�p��D�]��"�����o��q�=!�w��+������pzL>A!�|O�n@��UlDי�L .* )�6��	7�I;z>�y���o�zv����_P@��K����t�{9��+��k�����k�x�p?00�e�h��s���ޱ&Ȗ <�f�c�I�0*d��Zs����1���ۘ^�Q��ra�9.6L�����{�����fd�B�&b�EgrĬ)zpxe>�νA�vP�Q��4����.��n��Hݗ�j1���w�jL�]Vu�Ԇ��]��o^#����H�A���ć��Z�!]s7�b`�{�6��ָ�n�=X�,w6�k�ϻ��ӕ[+��}&�q��adTP2|�n�`�ON@�<�{p���J�쉺єBt؀1�m܈�JĨK{f��z�%u���P�c]:Bz`���Bk����e�q��6���M"�P<V���9�\N�x�hA8qh�iH��Uc.��,���k]�v#��*�2X�@�e�˭��V ��:�!8�T�v ��"~�0��4�S���k��_w�	�[���'��lׯ���=�}�r���ac�M-�E�td�
�s�1j�"���u	��]>�+����S&,1��MNJ����^@��F"�~f=]�dɞ�Ll}o��C"��0Lc��5��^|0-R����8��l�Mo5��Wmp���s�w���l�n�5��p�W�W�����)�&�7@sϞ]���Œf:a@�<��*���J�jޅ�����bz�R���:�ؼ����yp�:�1������N�β�@�MT,S!�}�7���:���	X�;�Å�~Tr�q�q�(;;G	S쌍N�Bֵ_p�S�#n���-�J�c�����oָ��'WΦ8��V��\3��t�۳�b�N�5���#M�(-/f����;�ڛ��\�qЭ}��F�R���,�s���z�(�T�ϖmb�:�BF�N	�d�S��t�wk�&r��������ŜU&�3�>Ub�FvT�(��pv
~�S2:���w�:�ʾ���U���tfQ������o�׸�Ӆj�F�MӶ~߭�H�(��3���"�f�3�n{�&��p�#�qH1`�d��0�6��{7sU�.:�C��t��q.��+i�[��S����b��Iq�#Y���V��)�_;���xF�è�?^���qjI1�k�-�n��V�g^[{[A12ºu]3�Z�P�����`��`2��r�X���f+J3.]w{ծ�e�7O�B�j|�%@��j�"�*9�TF�ڈ�+�1�D>�̂�ge�s2�r�Sqx+ٜ��Mqq\��ʱ�o$8Ԡ���E�鄍�+�.ݼ�B�K/�g�T�fn�S��N��4�a낇��*��P��DvAq�%�ߋc9ＶN%00�^�m��u�SqJr��7+N8N��g�����u> p�<>?��įCף���N~�����.��/~��t�ϜΈl����5X)�~�'����)1���;�J����+��o]��ˏ$�'��V8_�:_�����m��3����<�9En5�p��&��Z��of�n��\��]�먻�cC����ѽ��6V�r�ڠۇ�e5��wun'���^�|��#�w��W�UX9�q��ʀ<.��S�tn�l��x�����&ۘ��f�/�V*iL��ې�B�Ĭ�S|���8��]����W��P�,-0��<���5&+䓳&Ṉ�e���:��y[���hՀ��0�<ګY�߬qM�avy�zש����N�9z�:~��L緣*��s����	���� ��ʪ�4�%�Ʌ����L��9](CY�lhBͯ�TY�׹�x�A�4���ed:�M|�H�wR"�
' X�Fd�ꬶ�uD؝�p^s���7� �y3�֩=~J���q���*�*"<\��%Yh3'��M'U����q�qU�l�T�D�4�o��S̲\
��j�뎛�Q���шꍗd=�]�XX���%qg���:3�N�S�e��b*�e��C�L�5�7L�OodP�XmP�{�w9�F#`�_B;_�p����P�X��=t3����X1�Ԋ�1v����ي�ʎ�:��W�����qb�����+�+_�^V$?s��H+���9��ˇ*��i�)ɞ���ܼ7tHйS�a|�	����<��(�h[P�Hma��&�f�i!C:�[r���makhZ�Ypr�bd2��]��G�^>��E�^m�}��T��@!�2f�"e��*���%N�[}�+^��O���4	���$�S��}}.�]k�aUv<�L!��.��z����UCǋ[{`8!�ǠTV�E�)��r�w]�{�.��/�Y��9t���If6� ��>�6�Wʾ���Pښ<4K�Z�W��]�M���3�"5��V7�B��({�C��;NBru�D[2��S ��|4�Rb�dӂ��D�t�����P6Z(F@C8�-��ة�f0�h�bƾ��T�d�x�
w��I� t���8$˦�}ʡ��FXw�|~چ��C�e�юTM��*;S̙�����\��F�%9��
 gPQ�a�]>��\b�����\�v'6��K2N\5�Z#(��yS%�,y�W�
s�>�8�2��<���t2��kU�Tvjr�^��֫�j�����塐ګ�a`,/�YV*��Y=@����a�t��Oo��"w�\]�)��3���r��Q�u$���jt�86��N����b�W��a���V���d�\���#���7-��@ T�w������N�Y[�Wq={Y�xT�t+o��X������}9�r�y+aYh�֨���ĝ#���B+uz��E7��.�BL�f�64���r��e���?wo�R�,���׷�tޔ�f���ƻ4w�����wN��?��{V25�o��:����uk��Tۓ��\{���n��"�e7[�(BxP�b�DЦNqU�bNlv�����P�_Φ���x�75Y"��yjels�H�m�3�M� fQ�C�����%Hp������_n�"kM�آS��|8y��W7�;u���etX/"Xr'�(��Gp����P��b���{���kTP�\>ޒ+���lC�b��i��;n�eIӱ'��2���$nʦU]�%.:E�9�M}U�,�:zr�a�ڄ�(t��ɺ�� �11�N�9��5SvX�����Oh ʍ��S��-�,�ĉϟ+|q�,�9��6���Y4�ۘ�����3w՗6s0=@ �+Ni�6R?\b��qۯ����X�q\�h�^�H�J���m���x'/T�]I*a듁��!���mPw�kbЕ��h�t��B�D���gb�]r��R�Ә�tNf1��BKt;l\gN���캡ί��`ֹ���=���)�0���C�D��c&���*�IѮ�wq�c�7\m��}���w{(�����ٍڄU�)��{�L�L���	F7%I+^�͘Ǧr{���G2v��RA��q�Q�M�쭖s��q�ԙ_%K�ng�2%�r�w)����oRpq�Ĵ`�#���3KKt�ݶ���V�F�wF>_���>�:�j�RqN�͝�5!O��ێU���p/ :`��?*�&j:Q?H!3��a]LŅY\8t�Z�[�+~p^�yS�k�q������*ԦL��7@sϡ�خ1d��I��;����wNy���*_�'T����'_[4<8��9G'v�k?2y}j����R��5fOG[�5:\"��� t��]bc��!��q֫��ݔ��8J|�,��>�^N��W6�'W]�7G��/=�gTE;��ݦx*�6"y�z�7�ݰ����7��o:����sb��b��W��|j}�Lf����z4$��N�����U�D�V�+F�n]P}v���e��c@�<���&��og��c6��!��OR]e�ͪ�nm��ݹ�V�eF�{w&�w1	:��N�<�����¸s�7\�
�Rl�Q1.љ/=˥C6j�t��^�:��f����޵R"���X�L��^NS+��ZQ�P��V��*k�-�rt��GO�� 㢸
+�X�/�n�Q�s&�\폭�t�?�={"*��`�τ�=4����v�H�۵CfثZp�ެ�/�z5֪�p�h�v�C۳�5íF���8�RyK3���E��C-���J�K��oM37�s���[{I�4��R���t��t�.���t�����e�vj�3f�G��MGո�Ŋ���/�ˑ�9��QhQ�n���$Ὤj�������8.��o%t������>���#��n9�iά�3��Zv��S�*�/�l��+�h�po3�*۟H؋yN�v�O1'G�s �^�#e+s�7J�����KU��#��:_q�i�za��Ĩ�� ��b�e�� ��1De[�Q8vKq
n� �/3k^�;-�B�7@άOG�@jя�m50����:���$��#�/�^<q>��suk�j۰f`��bٗ5b�g��4L��Dd|8�@�4���s�|Ф˽�*�2?��n;f"�Q�{٘ہ�Ճ����u����ݡ�w�:��R�Y�Z�a�	m�컵ԧ�Y{y�:x�+`�R�H��4���?7��k^�t;`�5��*t�Їn.��([B�Y��!��d����T��Z���s ��-��~��d٧�z;{��t���P��*v����DsV�y&�X,V�}�3F���a*�+eJ�q�7�5�����W@����;m����9��4�S=��!��5x�hYS&���{H��:�n_]�=,V�	�xsn����m�&����7sG$w9n��@gs�������@].�Q�FK�:�/5	�)�صr�
5��f��Y�Pu#П,��k�^9*Y��MvM�b�*[��k'+9̲�� ��A�d��r����A�NʫkZ���Y�vw
��"X�J$]st�>Z��0�V�Ӛۣf���(�k�ް��+,57
��[aj�z͞��7N�DisޢAWKʦ����o{wn��B�{6�M(�����Ѵ� j��i	����n��)l�ST𑴾�;�.���k�w^ؽ�;��D���{�/d��ם�ˎǲ�9|VP����R�_�Y�3��ѡBu
Z�����sz~�JĲ�Y�K]:n����UA�i�uM��7��_��H��ZhW#K�֙�����T���-��N,�T�f��e(���+C1�䄶�H�&F4�3��'�����Wx	��@�>��kd���������=.6��'@_N��9���Gn���z���
��i'B�J��_W0��u��Git���Rm,F�������P�h�7x��ku�!��w���V��u0�)�Z��%���n�p��~�0�!�ұ��d�QS�֥�����c��7����S�[��\n�PDV��Ɗī)m�}a��F7Zs$z;����A�9��_r�$��§����̮��MR�d6m�ҖY,�x-�b%��$��Sc{rTYDe����5�t�JV>��CV�F�7�4��a�����f�
�m�(6�M��f(����u�E�Y�� �Vh��Y�KV����Z �QDT)g"�U[��DE\���g*HM30�]�	5b��"���AE�EҌ5QB��4�P���+I%5������UEr��R�S$���
���A�)�w#%E+����$�Ֆ�ŕTEd�����4TIL*�+B2*�gY���NJ�Zt:U�dH�ՕGT�:�J�ĢaP����L��H#QP#�d'-ifU]�I�E�U�g+H��RDT�^�QG9:��%���e�$���h��M5R$4J�"�g�ʜR���9�)��b�SIQC�V��U�!*(L���)%e�E�&agKVV�U**�(L��y��4�N�F��2SC�hs�C�kB�"��Q4j�ɖ�]�{��%��y��M����u=�&-"��3a1fJS�;�s�'��pF�{��X�VL������������������ꒅ��^�.�3h�B�p�,��e �9�8�F�L�v��}*�fؔine��R����k"��85�T+�rS���jJ��i絓�c�P;;V���Qr3�3j)J����>;�����3�$dCȒ5��A\�Y7h��
׶��|A���$��d�[�I�k�[¾�I�GΈl�{XS`j�x�y���g�8y-AT�fe>��+1�c���q���6/�'��s!���/`ݳ���,�w����a{�b�Hp�&�=C]��u�����-t�+����2a��vdC��z%ɐ�t2N~���k6��!��&�ZϞ�X���v�o�)�z�u_ 0Mn����������h�����i�bEq��⺐k%�.�;��=�����<��5	[yy|��2F�&��U1��fV:�M|�H�w�u�� �����/;o�'�v����E�T�1-�siS���'_4m����u�c�0E�t�pǧc�r)�](������(�r�7�EX�A��f�39��:���'9�����O�u�0�ws�f����YrC(�c���m�r;X����I��l�2os|�g�^v��N�3���"�E�����T���� L]XL޻��M�;:M��u)�˧��DDDA��V�-�s6���&n���O�#��}*��N
�?w��L,W��A\+����bj�'{҂4ǽ�ٹIh���叡�e��Xj l���X*�e'���4����.9�m?��L`�p���B�+	L��X�=�<�����9v�6p쎩�ӎ'u�ܧ����h����v�\eC@V#�x�+_�^QT~I1�����A���O��9�n�`Z!v��;�鹩��D��(�� �|���7��:��mW�5!�^�/Н�J6)��P�SÐԖco ��U�Y�}�'^��e��#�·�ŷ��Ԡ�=1�*���Ucx�j���{���c��ruE�dc2����/�iP��6�7צl
 Ï��"~���P6S(|���[�ñS����Z!���H�������X�jqA���"�d�"O�>$LI��ByL1��2����� ��+)#]�X�r���G��c4�y�\y j�q���l��E�����7����fq�b�vT��I޸�u�RL��i�_.�д-rUú�qY޿?MA���ں�w�Z*Pc���NR}�f����ќ0<.]ܱ�	ڛ} etU�֮���݌@rB�R��e��㜱f1�S���v�;N��E}	���Kɪ�1ki>��������:t�͊��?~��L��,y�}`�sGN�!i���qu�s}D(��*&��NG,��L`�o���鎄�\��, �',/U��Ë'���� �0xcg(UtՇ�[hu�Q*�a���O_ٮ�p�X�������]Pc�\�Vv$�͡�a<3T�"��t
)նcD 0�ȳ���2��q<w�e�gZ��
�xXNg�]���v��$���O�ћ:"����1�a�?�
⪲��x�v㶐�d1��C)�z��¢ɕo45&M��ҁ0Oi�/�w��_���@7\�i��ß�
����[Y<�-���q���:W72���]}�m\�ܩ�qe�?1(�Ψ�FN���a�6F%����)�j�àW8	]��brE,�n{a�1]+�����׹>��8H����\�7�j�[UK/����N����]r𨁢yp��3�S�u���l�Yy8�d,}��6�������&pNadEu!-0Ya��+|r�΋��eE����j4U*7rcD'���X�������=�Lc�VY]�t�+�$vvТ�ϣ���]��A�����j���cw�����κw��%�gM}��6+�s�n#���i�����5�ƪV�z�����^u��tݼ��4�}�<-NbE�������TA Fe���]�FT=��=vX�ޥ��������V3��}4�-�v��'1[��&���(q���쯜���P���d���cm�.�;b�lZ��-�Y�ȡ��y0;���=���_z�>W���n�����q�p����O�<����u��9��死njۋ�cqm@]\�H���KF�ϕ�%�C�&w\�pҐ��멷�f'r��\A�.��z����Lf�d�6�x0F��UJL�t�~N�����vVVGM�A���;�	;�3J�i=����AjS&M���9�<��od��9��-��p:��TY%��0�fׅ1�<{��K;g�����^z\����)x}�@�x�`��Ne�ً	���gsCx'�;e��*̬4*Wl��<62#�W���;G7E����݊-���"7u��o��㮭��G<��q��f~ra�30��(�;툲EE�V��x�H=��1����f��ƥ{����_O4����̅WYg��Ɓܷ��9�ы��\g΂(KV�&в||:��a���]�TMA8�	�*LҐӳ��oko�OY~�0e:�~�f��Ʋ����iJ��6��u��K;���VVw�1����"e��ܥZ	�R�h�+�j��=��MΕ��,L0��3�UUU}���|_t�C�3:�ya %cO�|��&W��إo���Ł�V�?��=j����_˄�q�&�<�3��{iJ�M�\�4F�p,2R<��/���n��W$ia8R�j�N�9Z�a�I�0o�%��<o�V�HW_���3��f.�')��1���b͋+���\��'�-�\��i�z��Rb�Y��ʔU�9��l}����p�[�T�V[�nq:ڨ{�f����(8����TS��A��C�R%�A���ۓ����%�ž�B�c��`o%�
5�������T+%�}�� �I�3�mV���jEF�\�*��=}qW�:w-�S�	�K9�kR:�³��^T��J�L�q�_b�>��n��nđƾ[¾��t��s:!���`-M��(�W)iVczk��/�^�Y6��Ԥo�`H����\to����?��rn��Ys��f7b�[{�[���c�r�
kfdVf�7p:�Wӊ��Xai�=�HN �KF�kU��BR�Qꆝ�:��Q3�Lb�ӽ��PV��Ѡ2\�]g��{`�̡W�+��pX\vMw�Џ��_{fsY08��q{7�I��[|�Qh�f�Pl�ɚ�yY��뮦�;��uH.u_aq��
�{��p����޵��>��!*����d 6h��]�U��pX�
%����-}��}5};X�|�b�j��}]��f�����YoD��?�u܋��j�$p���(�.��]��Y��Iyݘ��֎Y�����)�i�����Ֆ-��"��̬u��f$O��FM����k��qe�-a�Cj	\[��l��3#E��f�m[�3���j�'.?e读�\l����3E���Q�.��.pm�eޜ��L�r�D�ƭ����d�
Φ��S�q��$�q;�Z�K���Ǉ�½x>�6nR\-�K�t��� ]!�Ge��b*�e�+U��ng�:m"��ҧAtHۃZcuM�����B�*��(\Q��TFҠ����([��L�Y�����o[�`L�|:���NS=���k�j�F���2g�	O��^���R���o��g_�p�������A�-���z�|��MN�����Ox��/�x�c�׵�p	S�ymTJ,S���ʧ���n9�ڿk#%W7�PD폲���o�N��t7ڧ0�'$ؙuϓ76�X���Xg���U��ul:�ޏD�t����C=A8�2�򀭵]��[�M䙞��T}u���ږ2�q�c�,��qn��!x\&Y�H��Z^�C�֒�>|�)<7Y�վ���{9U�W�D�VRp�1`���tO�L!4$U�*��r�qWY�,�c��ruE�dd52�������M�U�&\C�D���$\JU��e��q�[�ò;l�|l�s/\�1�Em�,٪��D�Uڣ�҃�H�(Z���B����3�FXv_���cc6�riS�SiHɡ��ҝ�p��J�_B*d
�D�	��b{T�L�\b��>M)�Z��V�ț���}rc���*d�e��W����� �Zl���Po��|��x�j�)�_Jx�c��[�I��[]<��sUrn0�	�KϖU���c��ƻ�9Z��e�^.&��ko��wҋ�xm���@�fwx9�N��7P���`M:˜g�uCo2��0�����������������<�~�~�z��L�gZ������N�YA���\�g*�
}Ω�A������E��id�A�@���*�,�bx�w�P�d1�;�HG#�f)�u��
�5Sl�rc3k]��Kq�.�\�i��ۘl�`x{n���<_JV5Z�S+�LG�H7�b�k�]OK�4F��+z�>�C��W��|�՛.�ѩ��D��u�Mr �/cz�,q��#�V�w�]]�**� ��V*R��m��{n�w.��Eл�ݙ���<��J�2��f���.�UUU��7��H"�Wt���4��n�3����gE��%�>���J+���n�����k7�y��6zKv�y����7$,<��yLB�u\ܛ��;n�e��$�؂$�y��*o>Yה���. ��ǌi=�(�Z��`�ON@�<������\����k.TT}$ǜ��\���l�$��`H}P�+�b�l�f��(M|�[��,�/O�lS�mޡ��Ys��/1F��&���g� �������H�q����n��r��6ob�Sێ1��Ҿ��Z\'#J�G#�P�*a�,����6�R�Ov7��;�-�5h�ռߛ�c;ˌ�y]Qu�48�\��/K��u�M��A�EG3X�BinʋlDgNK<���v�m�������}P�I�C>r��c&���Z��0�9��xo$�1��)Tj���r�'.�e#�Е��C�*6��Pɦ�p.��(
�I�s�Ej燝t�:S�mJ���<��5��u�V��Ws�{�m��룭L�jS&M�n����6cVT�Y��Sr����n'F���g�
����p.p�S�;+z�RJ��X�"
�w�o�L՚,k̪1��V7�3n�_u*��oz��ʈ\�-˭�V8dg�9U��V���Ub;��lH2�B��� �W_r�ފCR�����>�ﾈ��z�2ߑ����N�g�K;��y�c�}eU~ci��\���xV��P�0�d]��'[7|R��Q���q�l,���xzʳ+�T"��X����
�=�
?7�~S�Lwۈ����X���2xPo��#S������.9�Vea�s!_yvk�n��9����JV�x�;�͂�%| ��U_�K�fS�f�MӟnO�n�E�J'tVqj�r�99Wb���ef�U� �e"T`o��R�l��?[��Dw\訽ł�9:h;`�e]y,ڷIߗZ�:��e�*���T��똆���@+�Xd��O2�b_�+�<#w�`"S�<dou������5h>	`��ә���T��Z��c]0n�e��y�1x�A�)����J��~^�Z�A�����8�cؼvD��ELJn2*6j&XSU�{j�@T������gŀ��&�d�~�B8O�Y'�
��䄪:���*w�t��֖�n���E�;��A�b��[M�r0�c����T+�rQ��>�2�ءL.L%7��Э�=0xbu��+7rƞg ��X�k��ɭ�!��Ί[y�Vz�5v����Z��i�KW >�_�۹��ϹV�M��ca�K)*��T!]�ΚA�Dָ�F�`DnT���C�u[�ܛ���诫��w�}���  ��9��N�oC����u�N��P���\:w.>s����t�l�}��'U�[�B��he_+�6�v�pC>������ E���'Is:!�����U�q�6r3d3q��d[ږ�{�͈(�V�jR7�6xA���2�OMu�-��f�,�U�|�8ˁI���Z�H�D�̀�әA�Ɔ_�}���'����=��\�c:�1=0Olf�)��Í[���t}Cf������f��S�.���}�`�3y�����g�<�R�@c�w��N�E��S5�rĊ�6>��u �J%�]�'t�_��쳏�[ָ���ե�NX��z��q���mU1�+��Π8]W� �=��7�z�A�a��_�t~y�8�ʻ�M��7�Lƈ�}���͵ld9���捵u���F�{2�f`��>�H���J����X"�#D�~5��aV�O�ت}�["Us,��L�G`\��a;�h�q���>�j���e��a/����:0Ҡԍ,56a����*���sv�,I����;|�s�ǹ�V>z��KH�rۖ+.酹Ռ��ǗZ�����f9�qRS����MUն��۵���zT�c&U�PK�ٽ�y\]V�U���[���ǳ�e��w*�����U�]	��_#�s�bu8�<�����}յ�p��� ��R�BT��.�[i��rh6 4v�������*�m� ��f㬳���rXܧL��)�&�R�w+w��u�m5y���{sxR�kh9��20[��w��w
���%������WG
c2��̑�/�6HQs}f�:=���M��������12��iIS{�y�Z�u:��*�|�v7u.#/�ӐN��qپ�{+0�tU�qD[Q��	Sf8lGj��w���;�)N���r람/�U9
Q�z�Z�1]�5e��]8�ұ��i�e�;��,�v�L�����Va�lѮ�\5��-�*�V)�&!4���#3�zBؘ��f���J�8��ŕ����l
�$�3�|�ˣu��6����G��B�X����[ä��s�i�YN㥘��i0����uxjʚ�n԰g}|�H��a���U���%mGC�>�b�`��e��;%�-��[��i�;v�\&�G\&p�tW�bY�8�,Bv�j��2E�N�j��GWë4S_6�7�(u�]��K;�>�j(U�x�탵:c�����/�Ձ��w�.��H�:^ػgR��Jɬ�.)n�d�@�{���m�b�M�����a�ٜ;{oF��]�p��];���u���Wd�0e����Q	�v��|���"�P;1�i]q���X��#��%�y��u��5�Vw�q�V9�M묔�=9��)�[�m�:�Ug
]t�̅!3jÐ#��t<�\�㾡6�w�1�k*��i�1Wo%���4����2h��E��K�T#x9�~�yԷ�d�ދ4C4U�i��`����Iw@����e�ȼwC�-+��я'�c��	�Gn��(Y��%�>b�\G%s�]��M�]�7"���t��ztҾ�_0/���K���0��l3s2�@�r�ܝ�,5��<����sn���̈́uH�>�M���XM�1m� 5ܶ��i����2�@!�8ww7�nN�+V�K4꠷%\�(�}�w�V��=)^ж�=�6��N���s�g=���p��2L�ݓ�V�.��8���j���sF�\�����TW̽��qq�j�ъ���s���n�d�c}W��w��S�YsίƑ��L��YlzL�]�C&o:��[��OX�]����z�s���z� ��.��`�1��{v���.:�5k������Q��X��\�O�N����宊�:������[5���wb��:�9w�%�4*P��:�`�A�v�>�p�Q���iH��̚��G��D�凚�ڮ��c8Sr��[�J�w>2�u*ɼ,�����i�{�å�.�[[����A�$�ĄVaJ��V��
5�aU�+	9]�*�%B+%����a��IJh��I3i�k-2CR"�Q��S#Tf��g
"N��,��j�ubp�H�r'2�wP�J*)3�uB����������\Dй$�$�PE��T���UjΖ%���d�Ҋ9UT.W
�4Em�"�^g"9NHs,,�t�!�g�����
�Q(��U������Q�-r�3L�,�r���,�r�r�2��Z�=�ݻ(�V��V�g%hN��E9.�Z(�aDUI�Z�ęC��T�ӦHeADDgB�J��Y�A�y�iEʣD������*����[���U�eDUTQU	�,�"=�r*�*������/Zr����Q\�ԏ��T�󚶄��ؾ�Xg�2����sS�V���+���9�޹+���qY��ǘvEposjV\tT�h�;���}M��)�+:��2���S|cp�8j!��p�2��#eHEQ���K��i�]z�mE
�Уv~XR�$yU:Za����>���T~�Ek�oƗa�s�s؊Q�9�*_�����؅�����0�c�rw��q5::�'�IJ��^�|���%��곀OJ����q,ا��9T��CRY��t�x��ۅU��s���א��eU�Ȁ3%�BK�b*����U��+j���m���>N@�3c�k;u��!EF6�9�Y�3xg�Ǚ-Dn�B���0-^Ƿ����N�0�)v"yF�j��:�\�@\�q����7`:���
ND<���mT>}4.+�C��zf.��8�
gv_W*��~��;dC���[%s��H����J��v#��lW~�̽W�}6�R��f)���W�\��?l$����_X)�;���]��VQp׻�L>�j�Y�Ϡu�+��LԺ���&��� a2���eX����'�Rh���Ń�(Ջ�0�7}��A�B�TXa!`3��H�rF�D{zn���Wt�yFۤuh�X���:��}D�
�v���}�b���8�l�Q��4%�yfh�)^	g�j�7j�꘶'���sEgY�jx��;Q�4*ML��+܏� ��ۑO���[z�?��|u� [3�=��vS�k�=�&��\�����}�S����fgK�-)3�Fħ�h�
�^V~��(<.Ul}���)�����0�6�:�Lm���i�)�*��;�����J@�Љ����tm�?@����������H������[�Y]ۛM�L
]O:�!ɦq9�����W��M���!q*����Y��Xmr����y�s� ���p�*�du$��q�3ʧ�ÿ+��3��%���c	�U�(k���k[yX�J�����P	d@�v>��������/
��z<2�n4����1�@��y�S��>"ې�ȋ���0��p�]������x��3	Ҧ9�K�̇��dU��36gڰ)lqǉ�m�T�T+����/����(K�OO5%��Z��Ŕ���;�NѴ>����\'�ν��'�K��z���₸�f��k�v���Z���d:�e4�bx�$P[���iW���NaU��8Y��Z�m����=�/�x�u��V�ĺq�ic}�63���6me��F�&��d�!$7:�OQ+�ުߗL;������Xx�%6�.={�J=x�;�����\��/VL�|w�����hl9�����}����#(�"��{s�.���0�M����6;5Ƕ�o��>����-��/d��{��FC���g4��	�q7�7PpЖ~������1.Ol>k)�wԨu�����9�;r *�K� ��5hg�]"b�1��P���\MA�!ೂ����:�3����=��n"�Z=y�W�����Pɦ�p/� �� +���ʨ�w/�Zn�j˪�-���|h��-�ګ.Vs�t7#q���[�!�5�����_[b�T�'S֪B�+_eب�)��k��~�BJ�Kfnr�w�<�]��Z�.l�أ�1ug��W4�$F�ه�~d��"s]e
���� 9�0��Ҿ�~AY��Q�ޛ�h�6�х#}��#�����O�3S�����ꌫ=��fa�s!_y|ٮ:wh�G�c�޹�ZytgE"�,���D^��!6̧:�?���7'�u2*�Q;�^.���K$��/��ye������+*4\̶J�1y#"��d۟����eѨq۴W��O����ǉ�^�t��,�u���FUlU^�y��d�u����:�"��R��.�(�q$���5�:��st�ʵ�N���<���~I�����^��+��M�2�j���K�☮�1wz0�^n�s;�O7�y�4��gY��>Ncc*`�V�o"��}������v��3�[���=�HT�}�w|{���>߁EF����;tF�s���*��D�D��A,7�l�>�?����� �j	��G����뺲�8uu��p1���N�8Ԡ�ʸ:X�/�n��ۮ�){ϳ��CcD��|>�������j��D�~���>m��'��	{w�?C�Θ��I�⬃�;A�<�����G�jg 1����뭕B"�������@���V7�yMmj 2�����zy�U�
���*�;�r�؄�&x�Uy�\��b�<߂̑g���0M:�<�� �E��6�����!V�s+�I�E��+���q���י�%�譺���ر]����� ������!3��h)�x��k�ɉ���z�<s3��ܭ]\� 2$F���)��`*�O�A�QJ�����_:�b@�V��Ҵ�� �p]�{��uZ�J�X��F3�jLWͧfKf#*�'e���z�?m����ut䰲����P��a�cF=w!��H�	��j���Z`�_F�uk���Z�������aT;��Dwm���om VJ@F�W�Qt5B��=Yx��^V�Q�\8���+ڴ9��үF�zOw�F.x�����6#��}�.⤾Ǹ!�����V����
�6�[{X���;�l�g7��A�w��2�BC���/����������%�=�]���~&�Y�xGw�z�тh��U1�e9��35�Ȅ&��;���s�xg��m�|��[����wN�;e3q���}&C�3��|Ѹj�'/��v��^V�;i��W�[0E�\�d����ҩ��
'ǎ*��հ
�e��4�0,�6��i�����}�횦+�Շ�F͓�XK�ki�ё��>;,4��Ou7��˞��+�i+�Q"�h�]Jg���
��:O�P�;$�JqoT&��5� *
���u��x.����dd�]Vu��:b-�L�C����1P�*Q����~L�n�:7��Oj�K;��=1T~�sw�!�b����ޟ{�M`�T":WL�����<���@�q��$�?A��@TV�Eb븖lS���.��RY��tӏ���z4K�;Q��co�\�ɃD�b g&���^�`�=/������^;�y*��3;��Ng]XX�WK�M�z�푖晔H": ��肔�.�eȀ�q��\;�+�8�3�V�(�J����o���GV��ϱׇ�{-Cf��]4=���+�;�kH稓o���$Fw	S��f��M����_|(qW�-�罗���㓴c.��]��t���.��cp��f�r��k�xV�N���q��W�W�Wދεgbsh����q�G��LS(�u��Z���BG}����x`P>Q֘{(&�ZsZ����l�?m}u��9j�9�2U��)U Tt�v�L�;�c�}!�|��컣y�A�2]9�b�S���z��	*d�X�����9�"~�Ӫ�[,d�s8�l��g��[[U���V̮���5.�x����xX��健�ʱ�g���"�Ӹ�P+y�]���6NW�����&¿�U���H�v9Lh�ܛ�:�=��\�U1�E^hB'i�4��R0�;S#�rҹ��U�l���Px\��I�T��
oo�rO�����A��{��%6`�������gV;�,���պ5��Z�ѷp���p���U��W�g�Z�Μx�H7�8{�!�Z�b�g5:���|c�1�N� ��0��|P��f�pV��g4�w���iN�oV;�de$���S;�+��M¹�Y��8�r�w�s|�D̋���l��E8)�[}@5�E�$u�Ju�~ҫ����Q�/�Y<�^{
�b1#���d4y,'JYy��t!�
9�LHڍ�����W7��T�"�۽3�57�^�G��Y��Y��4�[5���>�q���f�9�FN��
雎� ��^QǷ�RB�^���q�Fދq>����$Ǫ�C��6�^z�|I$�k��d}}�ѡ��?��/���*�*���j���t���ˇ�	�x�y��cc�S���Q�jpl
&ǩ�m�Td��9:�*;p9<�J�|����j���v��Y{�� 8��x��N\�\�{I�x�K�Z���o��1w���*���������Wr����-�.�i�r4�,}z��^�Y��Z�m���Su"lT��F�N)��}ENҞ:"���51zX΄븛n�ᯄ����TH$ix�b�;��_�7�}|�G�}T����U�TcRj�ȇ.�?1a���V��t�5P�Q���m�j��3�!0~\B$\��Q��H��_0���?�T2[s��0�bZ�QO97�H�=\ݢ�������_#;&	e���W��{_ɪ����;�m�������Q�w���������Z���mu�߬�o��1�}�����'��H�AĹÙֵ��z���+�c5�̔�dNl:�5�a�: aoD	�
����}��%]돳��ﳸX]+^�S�WfMD�3���Ț.�T!k.�:Wrצ�hϺ�*@���-�#�ut��oRp���̯�ݫ���a!�]�9r��>q<{�^_d`WV�ᗜ$n�����fW��0V�9��}��Y��zp�ظ,)�oS��{��3��v�z"#菢��c��2�	�G)�����T�##S��WǪ2�P��?1�6F}�<��:y>{�x�L/n�1N*�7 ��v�����1���_y�Orc0�e���hD���G+f6JQ؍c�#P��$���a������ʍ3)���0����2)L6K?S�u=�.����D2����Y^�w�J��[��v�F�<O��YtV:�O}"3d�4n�\�&�)�_;�wµp�����]os�j��+�)���
�����lJ��I�TN�:	`��%R�g4*���^��0��U���N]�u�h���X���=�:����;A�;;ep<+�X�/c�Q����#��{ij����*�H��H|��t�d;P��}��~�#�I���Ô���sA���Ww���&C��7������A�bƵ�ь�r0��85�:������r����W�n� ������A� IJ� BE_@U�
Z��;��)�݄�%���[*��In�8a��q ���>O)|8|;�>��Dg�[¡&��s[��oI.ˊ�їK���	]>��rQa�3W�%`(�r4�8m��h�2��|8m�#�v�T��R�$��Wd�t1n������9��뱖��8�4H�u�cT�7cF.�si
��`3���4p�Q�B��ՙ����`��U�����G�DDF��}5IkS ��f\K�3�r�)P�J}5˷r8�X���7 u�!׍����[7�ë��t��.%oT��ب��9J���0j̠��&u_U�V�hdM���M����q�Tk�;�فkh;镋�<]P�7"�tr���¹e8�5�}���tjӄSg7��Db��gl�Ĭ��//���۪uҜY�˚���m��8e=���^nOu����ljq ?UyZ��K��0�������^s��9	�B�v��:E�3.;��E�~�L}���9������Q3u�{ð(�Xӌ1��w)Is���+iCD*��U���ʨ^}G�-��K~r�Á����m��(�ֹ�mf�P4���_7͋�I��U��nPz૘Ujѭ�-�y��X�7�ç�᪕������i���\��=�R]¹�|�"��:��'��vj 1��nA�v���؞���΋#yO(��Nu�ICkgqXme屆V�������{����Z`�;�97:�ɝ:�ˮ�ʀz��}�gZ����锝�	Q������]��{��v�|�s�d�ͽ<�w�興��j�����Ԩ��:z�:��R�o.���=��Oo�[¶ΉU=�����������(�ԕ����ٯ����kq�̃vC{W$ޜ�ç�r�C�/hPs�>��I���7�
�K/�`T�R����t�[WN+Zq�Qm��r��������������Zn]�I�ڮy]Qu8�o!x���*0��#�@���y��.H�UY���Jwy��
h��e*�|u�i��B�9øE�Cg�y�r��bT�.�#kz/���r���v�����'�i$Æ�+)��38Y��s�M͵g�� �7�:��n���f���5'�8f�7�\��8s��3K�Z�δ��>��g�-����~^kL?w{b��5�����+���@�N���3��� ��k�f*����Ըu�WBfp�6נ]͞�Wr�z����C��WZ_Q�=K�gWYs�s�l�]��j�h���R����ً:����ri7]l$�x-B_Z{F���K��cjӨ�0�st�F{ ��+��7{����ؖ���PrԶovۭ�^9s��Wf0�Y��{S3�Q��T��rS-�N�t=�*,��I4p����]_GI���D֬=5Uv~��.�S�7�o��ōx�iX�&�R���ڰ�l�.�43kN�+T%	��ĩ>"�����w�
�%���I��.L����L�;��.H���q!H�Y��vS�k������P���|>�7�ΞAnN���u�wM�t�=;2�$*�ءzwY�ԟ#[ڳ7�dۣ���QT��w"����7�*F�ı���DfÔ�AZ�O�΃��]w`:XiΚx�����W&�-�]ǔ�nr���7�
һ����%�,��	i�N�_Z68�k�)	_s�%��k��N��\X�X\�q,��,����դ*�u�5��5��:m ���I�-Jx���c�·�h����b�1nG�4 yZ�Z�_Z�usHĭ4�OJ�V.�����諂�5`YV�6���Kh\`hyy}�"A��.X7u���eԫ����4cI�ް�|��ф̼ŧC���ݤCe.7m�V�W}OK�BT�����#��M�{��ml�o���0'���B�F���Wد��[R�M�5�j�!�;{x��Z�Vؙ�)4jrl턼t�{ymd� J֥r�M���u�)3��A����^����B���E.�[���C���3h�,��f#�;��ӳ�v�#�X�x܌]��u`��E��행�Er��T�.�j?A
�/a��ee�YV�}�x�d���0��F�S|�Jhu��ZOU�^	z�
V�����ӴPɪ*�wM
=�|�Ϸ9t�Dg��/��}���ƈ\��ۦQ��w��4��1lb�|z���՝J�c��5<o�Vܓ*u����φ,�$ჷbJ�t�}�����.�P��Ԕ�y�3ۃ[�c*[����[-%]>g�Mv��3�K[��gFlYt�� ����8�c	�{s"�Gx�Q�c5�_T+H�p]ݽun����!ݭ�̌�WD�<�V��ǽ�q���D"�Im�\��';��][Hi�0Iu������^��fܗ�c�Cvr�w���wI�l
gR"�eck��5ő_
�7:��5՜k��v/?�2�������oŎ3�vt)�k4�+s_�h�v�����O���1�>z�̫�8qH1�S����_Z@����\s%�5h�S
���<\�gc������w(�
2���au�������,M�����N�Ԟ�e�Vk5�R9�up<ϛߒ��yu.�Xޮ�m��0�6���L3S�Rt��3������:5{�'[����~�9Pb4�E"�Q��$�'R8G(�9Up�B=�rY�r�*�&p#�TIj�sD��ds�5YTEGL�e29b�;�Q\�B�L�IFJ`\$��Ge�H�d��B�����s��霨"��NT�.W ��(�qK�U�B(��2L��*��%��r�28I+�W�:$�H]p%B*j.�twe�A�Rԕ9Q)M�=��S�Jt��8RgHBI�B��R祚�Ar�9A�V�N����uP�#$T�'\�*�]*
�Tr��B�G
�!EԮUA]#<3����g�j.��3*�<�0�Ȯ���Tps�ʲE�ՐG��"9��N8f�!��**��ro@3hձ3�9�����/�T��[�b�.��.ۈ�t@��Ivu�Ջ�M�5���V�>TEr�{s6P��4��G�}Gt�r�N��*�|z{g'�v���.�
s3L�e�{�n��Zo�)�˰��tLV.wsb�[��'�/(���S�-��������_T�-��<r�\K�wz��b>d�l/���{cg�ϋ!+}�Ӎ*3�f��S��Xʸ��F��P���J�cb�s{��5n����kSaT�����L�l����<�GK+z䥪Wo-�o}�R���D���L�4�;�Q�B������P����A�N��mN���<���+�- ,��*p���{��	����E�[f��;�}�s45$�����vU�J�w,��q�/-í�/��k�\gTE�2��}��X���;�2ބ���b���r��˳"Ψ���ܴ��y�'�)�r���lN1���������� &0����b�[�*i\2�;��5�շ~cQ��@Wo�Z�i��p���Ӗ���������a��@��}V|��ø~�6�鋹������	� ��Q�o>\�6\�x���H;l��׉���p�h��ȻJMҗ[��=����[��ǪV�[&��e+f=DG��绀O5��T3� �P�`�sQ<�j�7�f�˙��U�(���K�b`�%�T���≮cd�s�y�Y<��]]<���ct�k+r(ƨ�FQz����k�WZ�C�� �T�n�N�t��M��'*[���w��u�A8��Z��v'��읧s1���F ����b���&Wn�>�֯��Ӟ�R���^���w	K������z�.f9ٺ�C0ku03z��u�{r��N뙽ۈ��m�ڢb��eK�S�ϧ1�����dK��Օbo��'�C2���#���V�IL+�c���4��+����"��D�3��s@���|=T����ʤQW �T�[J��P��K�x��31*rf�� �W�v����ʤ�p5,��+L>M��u�M�jݧ*u1���M>�t�����HG��o
�U����h�m�fU؛��+&�S���8ά3�"op����]�8��L������n�b��L��=]Wa�HW9��T�ۮ���ӆu�&c�.�2vs�;4�+f*��u�2kx�g�1���!�ot���xK��!�������>��:'(�+���T�˛�|ˌp��Ol�s�ƪ���<ԥ���/[��.��(p/4�|�Hn=��)嵭vk��|1����%��m8YIeX���=�Z#y�_�����_s�9>��-�\�|���\�9��<�]�R���b�w;���W9�]ޒ���]({
T���k��@T���%q*��#��F��5���;��S[B'z����7�fq�m�w���R��7"�P:����i�T㼌�ί8��oc��{���$�5�n5���ƺ"c���Z�w��^�'��ݾ�b<9�#�����O�i�J��N�Zp�Bl�u�������8WQ�l��V����4'��ʁ��켞|�F�ڽ�wK���U���[7�f�4�B��`&��N3FO�ۨ��}`��}��z�x��X�N��NNi�:�����pYYƬ��&��b�r�ot�j����?�K�f��D(�i��ݜ\����p�-����r�J�d?IS��Vu�wJqm��֡%��y��	���\�e��Iewe�ҕ�R� z��>�i�h�P�#�sln�sNiz�����5�zU7(�ժM�?^Oy��̯����M�d	����R`m]��m����5�_J�`Z�g[b�ս��u�/�[=i_i��9�c����kiYz���k#V�ܨbb���ä��v���9T��j�V��wM=w��䫷.QsДc��h5���m>��s�5��m�Y��_#�lY
b8+&j�g��벫�J��o-�o.1�ڄ���|)m��t*n�\��8� Ê�Wө+[E�C��NSˆ�[TsȾʾd�fjo�@���FT)J$w|�$b���g\*}.�I��-H�z��f�WH�3��|�gT[c)�3�?G}���Z*��i���bk�j�T��⌑��;�ZV�kY�
��s�f8�uR��8ΡV��خ��Y}]B�p�'�Jո��1�ֹ��
���;�f��;�pL����0���/��\2ؾ�� ���;]_J}��u{}1D�{�{~�ꗭ�K�o��7���u�Q˝H���b
�4���G�Ƥ3�MG�{���k�,o+�­<�;&�:EM�ToZ�jG="�[��Oκ�=��]��ep�ݟ�W�W�t�C�|S3+��OwMD����:��>���a�n5ڱ.O>���	<����Y�yc�n>m<s�M'�]<�~�v���3w�s�Д������u�u��Y�tVy�7�?c��_9��l��F�=�.�<q�p�T��2��ڇs1���؃�]��_L����p���ո�p����P�@ ��oB;�9]45�u��oY�%��Q�-�3b��T�3�1:ƽQ�X���sb�ս�N�n�yG�-�֕8�y�:�l}�	]�K��b�T�����j�8��>f�sb�'�bN��o=l*!�ݭ���d�^��WU\���Nʅ�k���s{��429F�ğQ��Pg���)]�[1�g%��� 򨝖U��%TBR�cY��z2
��{p��we��OC^��_�kz�P鏹�|�I�[E��Q=]�,����f[��j���:�n>�O%��3ae�W��GtR���VÒ�l�g�_AF��a{H��k����KC�C�MA;�@�w�)_WT�f�X7�11�����e^���m�rՁ��Ꙭ�V�ťKZ�A,|��Ed�ݧ�~������i�x��Y���w�������k�|�J[�LwϦ
���]��e�;0ޑ��MtcHt^�%Y�_O9}�ֵ��:���(����x�1�ޔ��^R[H2��@O�d�K_m�9i1z�=��sY���
+��q�׳�Zu})?�.��-l���b����I�p����2��iHP<��~�����d>�3�t�>Q���5˶�;���mG.fJB*;,����+uW9�� =�w��)D�r;b��lFW=���r�=	�ƙu;x�m���Ż%Ŵ���q���ƻ"y�kj�Q;۹��c�9\�%;����QO��}�Z���']x�2��v���+7Q�9���D�r��w]ץs�U�%Nf�9��۽�v����ֱ����vn��j/o��B��gBN��Q3}����o���;��x�Bzվy���ybu�x�bI�Yj��o����m�$!�p�'SZ��S.年畋��V��Ns�*��O[=�BO@J��Q���u+1�Mr�˵���k��P�vZ��_�deoe�x�v�pE5������Xn�x�Q���{8u%�;c��G�Cqy�H�}����ox]����\�{+nJaX�f��͊�13}�sļ|{/�7�=$5��[T��*��tk�X�
���s��˻˷�I�!���;M9��w״޻x'����xLW��(��4��L֤FQ��iX��C��\&�9O8��FD�޻yT:�Ax��Ncwl��/C��r��vUB�SK�ۇ���:^g���ۓ���k��x�Q��AT�� �>��RKd�t�YN�ֻ>��{E�� ���cG%��w����g���KDo5h,�Z�j��q���Z�:���
�rR�V)�������R=`w;ڷ��UpSy�s��ɝ�Z�.�[���qs��6��j�J7�Ώu�0=�N���K�tv��	C5W^)�h�][ǧj!�f�|�0�B:�f���t��4�t�ח¥���q����뎾�e��sh·�Nr=��&U�b�+i�W&P�OV)���G��]�f���+�Eӵx̢�K×tg�L喏WKY5v��'��^��䫹����ݔ ��Ӻ���C��.QVS�d�Y� �듫�G���Sf�A�d�W�^��\��0����I��6�]����#��k3+*Y�z�*Z
u��g�ES<����k��V���i�<�;]rr���.�|��'���Dp_�mQ�V�mfrF�t�'��=�j^�'���j̉�y�gb���"��D�a��]	���4��P]�&�u���3��^�I�[�rʆ���/^�ԛ��y1�F�̢�G�s��	�	ۋA.�W�J��� z���_���ս��5�q׳��9Q�eAW0�+������t��t��Z����Ui(���5͋t�\*��W��휪A�q�Kݸ�(S�}�ޫ��
���Sr�ca`n�O�������B��� T򻹮ܸ�G�ޝ&z�yP;�勋��*�R�p9�z������Ε�8��3Nf��d��:��[E�:{,�mv���9����.��ݧ��8j�۝)�TOet��=�n�>��yO�����$]K�}n�+�}����\�4�R�vl�9N��hnm�J��;9*>V���V�6��ڍ|9���8�xMs"vu-yq:�wN�;����H���=�_UP�=��ӄ +5B�}k�W�R�:~�ID$�I^*��{��m<�֧�WT]̿��gnBq�V�ʈr���S�wI`��0d������]�k��U+��{ݨ��3��@{��0��#��&��ʘ�H�����M���Ӛ���n>;MsV������R�]I���F���L�\R���eޠ{��9���ܛ�'�RL5�n5�Ѝ��q���x gv}]4^R���f��<�U�y�og.x�!5Fk9��-�/f֞��1��{��ƻ#�襛���{�:���<ܓ/�@0��y���v/!�����U��;P�gU��R���m����[�i���9\���}:v�^��g�w���MjU<A�֖���ES���RO�y����}�wƯ$�j>��O��͋�ս���ۍ��vq���hr+0V|<�e����w����oed��D�k������y7��h����w��Ҝn�pM�A�����wXx��W[�P��Ӝ��.����.q�R��(�к�,���\�f�cV���}�ǣ]��gD�1c&� t.S��>�n�F����	z\>��{+`�k�8����\ظt�\B����M8�|;Ej�u�B�U8�l��Aus��tkiBQ�WDlR�ohf/M���j�Oo�m��ݳ^��*�!o��ك�A�S���%o�U!8��
��řo�p����,z��t�Y��;��A�ԟ=Jn�Ѹ�ڶ�t�4��\C���k���Yƒ�wϦ
�;�Td�ޘ,e6#	�Iګ���$��^:�p���9}�cZ�����2�r�HY�]s��7�W�|�� ��jJ�^�Z�n!�I�ם	����̔)>�8�uh�o�]���%�4�d�琯�-�	4��_D�gn�.��wqnn�Sz�H<f\K�3ß�*�h%k��]�ܚ�������=Y�:�M(K�5#(��Æ�B�?)D�C�X���r������;�yp�K�M���
���F����#}2wh�T���7�����Y���5�Q�Y�>�ܐ�5����jV^��b�m�l��
&4)�r���b���ë،�r�3u0F)٢��r�m�]�NS�+�,�y�|~gz�_�9��q�6��P1��C@�e��n���Ǖn��륓h��}n�;v�O�(]M�O����|uR<��y��m��1�9�K+��ה�nkΊ�־�;`#�fڥ�@�HMѬV���6�cK��D5�����9�(��wW���ka����p@=@��2m�ޤDe�kj��7M͒P��̡yZHi��N��ih���7s��,�]ML�XE6r86��z��gSzK�a��weol�+�hD��*:�\�E�w\/8���9˪�-
Ū���4ed97:T�u�"���\U��G״/���d�^�����:��x�aI|���8�+�{��S��d���w��CW0pŸ�T��[uw�i�B��m���F�.n����'Z�W���%�6F�b��B���k���˯f��h��r�K*�޹�'iVQ娍��=�	KN�Z�H��:l9���A�T��F���;#�����E��\�@��/�AUc���0��b�ՠ��-��]�:d�2R����v���[��B��P6%KIft��\6ba�xH^k��Q�o@Z���\��)괰(�c��K�Xٰt���@=�� 2��#0v�C]h1�9�3�2�$9�咻.��C�펽+�r9�čIq�t�n���t)�IǷ��Z�������
���&��b�>ٛ	�Hb8�E��9�����[IT���f^�"c��޲�(u���rVq�Tm+�eoQ���g4�tR��¤j�{�uv�[��%�t^�T[b�.���6i��t��P���Ӿ:�el�sU���=C*�lfv(���yk�#��|�dW��뵊�r�j(�?��4Q��D�41��ntںS�q���m�����J�O4�f�W�_�"�����	twS���z�L�Kp�mΤ��s)X��v���dJ"�
���{qR���/R��lS�	�G�_ ����սM��K�T��9�,���^V_&Nvd��]�Ԇb����֧mf_S	����Vi=ǽb��XGcQqhS��颥CQ��n��T'=�5��2Xx��%��Ij�3&�MrJ��W��[�;���O^�:�FV�@�h$Cܝ�w��ro��<�����˗�M.hȲ,搫�ܭ����.�T�F\Ţ KwA�%� C�ݴY�;z�pЮ�\�
��:�\��oCfc��G\/�nT�����x4��H-�V4��3嗧�_THW;w���YF�ĥޅ���i�rإ�+����y���p�o{|�ɋ^�\8rSi�9!/-_wr7e�<g_�����./J�����=�>t*r�[S��m��@6A$r(�r��q�p��E��c �$�5L���8�w-B����N2�ЫP��NK"��	r��wi���z
���EQG+��C��hE�E��/G+�B�a�a\����DL�+D�QJ�3�ajܩ
)����Eȋ�TG�d���!�L �Ҡ��NC�z�\�4OADAtu��	��0T/2��waUQG.�y!ȎE,�z�q܍@�E֜�U;��B�S	WD��j:z^T��!Q�I�('gY*2�,�����E\���Մ���
β��Z�Z��"tQ
 ��YĽR\���\�72�VE�b�Q�B��K�mK�2���KC��r<P��'#�nN+��es�+D"��99�Bp���\����r��
��\������"�aA��	4b!n�չ7.�+4�<�����΃���g(��x=��u������/z�����gp�H.�+���ꔕ�s6q��}_-�}�[C"�?|�q[j�}��7�]Lk�'����;U�e[s�u�\eۑ}�9tn�8����5���bp�({'j��x�k&xn����nM[���WJ�TV뉕�O>q���[������Y��F\���Ux�K��8Y�ʤ�X.�ޑ��&m��Z6�D�cN�x�|����9OU	ƨ��3��Z]WRv��G!�_s�쭸�)�cL|��v@��mV�'�����
�?�[Ԗ��,���~Z8�6��F���)��xv��Vm�Z�4&�1���o�܇i�uۮ�ol�78���5l�Qj� ˮ�R��u��L��+�ا�����t������U 7�)�J�VGOZ}������J�=}vU*U4������p��Ol�X��ٌ����ϣ��X�@c*\�@ԕ�h�/ga�ypֵٮ3�+ ,'��Ej�N��7���<�d�mu�:��0^�����&n�a�V��N]٦��[����>�K�U�l���q� ���
����ư�ٽ��T�Q�g/+nu[_p9b��yZ5��J𻼁A��mr9
��	TjX�Z�Ԧ���IE�/Gľ��|�^�{_@���.�+�F�V�Υ����䅳[{	�%ͪ�j��ek��Cb�G@ޅ	C�۫}<���mM�rf`�ajE�T\�<�L^��=�P��¤g�#�	\��ԱJ��Lm�od�a��&^_��>;_5��;�v�Х?r��k�u�����jV8/q��5�k���D'�jL�c�pu��Ԩ[�V����;���z�{W�u��zk5�k�W�ѫNM��W�����Ū��Jg{���t�-m|3:�e�_�˚�s�h�>5^��zt�+$�����3������lJ�����Bo��)�-ڞ:���	�]�:�^'Kt��NOb8��mQ��y=�n��ʂ�=�>��U��ط���u�ْgr{"m��8�)6/�V��]�[N����el�A%A$a�Հgf�kY���&K�f�~���oMCBn�����5'��9�=�;�~��$�b�Ӕd9�4z_>�o�r{:�[��m��1�8R��1j7\����������k�ϯC�<�a���IwE7���fX���s�֥f���;�Е�ƣ�\ݟoz�cf���.R� ��؏��Ρq�v0B������_F҄�k�c�7��|瞅�����r������2��*�����+��.�벪!R���=枛F3w������ܨ�/_-�[�#�9��A��E}:��[E�{*������L��[���b(
�>	�ㇵ��JR��C����BLU�����K~���/x�9��,��b�p��1o����:�����
c��,E����QN��,��\�Ha��|�w�����|௚0��b�`,�bz]�.�v0J�
|�>E���Z�/����ø��6��+�"�vJ�c�8+�6�ěV�~ͪ��骓�C�B}F�L<���)��ѹ}��J�g�jU!D덳�DO���+h;�p�yoRq�t��oh3���"�j�j�(P�]��j!
�ip�ӷ��}�.�J�����V��Xo�����1�Ecb�ˡ��*�ޡ��zF�m/o9Ԁ�Hl��sf��� �K�u)ݲ�cc�4��i$��Wl�v���<�8��!Mr����I�t�K���/F�Һ�J�*uF���E���4ۍw��ds������{�W>a�HwC��ek��A8�ի��]q��*���^�Vt1���N�|�{��{��a{ki�7�>}��&:��N�k��T�X��O����Y��gz����֥9�ȹN���(�U�2nu'~�C��	����������4&˃vM�����Ӈ�0m\@�U=��%CQ�5c�o�\�r���F���j`������^�jol�R� ����_N�5J���Q��(\(x�Sj��8��7:�su�D���6���b;���ǧ��m�i�ﳦ��y�+*u1���7j#}:Oh���+ f�pC��f�fCwK61�wBj�U\��:'i?�Q�N��'�����c���`����P���ʤ�o+�҇�M@O�����:},�����ȍq�m��)te�W�g�X�FD� K��bz�"�i[6��;���.�MzU�Ní�I�,&�_S�RY���cwe	o��'f�t���x��+�������=���{#�OV௳�m�B�r����Q=��Or=���Ţ�j����3'�<[^W����,�3��r�y��%�%��w��+�6�k�rҸ��׸�h�h�`����e�
v�^��!��ɿ]{����7On@X�o�I�+���]/^gR��!�5��)+��H���9*����j�t{'{h�W��ra9O��w�M���m�v�j�!J&y�S��?[�Ѵ��e���X�\d�J������I�_&�]º����O�-l��7��
�j3���b>����q��׵��_ܝu�bpʸ{'j��wCe���;�S�S]vR��t&6�fuL�a��z3S�ڷmK�O(}G������3�<9�&�j��F�̯�s1Tͽ�+F�j����vΎ��T5�s�ʦ��]O�n�m:5�]��*�쭿�JaX�TI,����s*�����.'[b�ս�v��l�R*
�`~�*��?]���u{��h*V������9�˽���ó;���F>Rv���,����Ҳ����}�=W�9ŋ�b!yaQ᳞P��oQ�C6wR�̃�mpqS�$�}g�]��,�G�l\���Х�gi�Ld��&QZ*���r�պ��5X�(�Yb���U�\��;M\y�d�MUS!�T�_�Gq�T�sYw���_;�vQ��qT�ҍl;[M>�t�٭��Ϭ�+g5��A�X��A	�����:쪅J��7��5����Oo��:�ު��7��	�=5��w3CRV���t�i�ymk\�����]�g+s����5j;��K���)�T()��}%A	h��f@Y�_I�QY@涱��ޣ�T�G܅� ������e�W��m�����훶�"��ϴmCm+��o =��FD*Fx�t%*�h7y�a¨�z�м���=2V�Ƌu�c�s5�����(�CQ`��&1NK�n��+H̦.��wU�8�ծ[K�u�}F�I0[q��\U�=b沯"���*�m[Ϭ��\9�^����zS���<~��S�b⺵���S!��}K�U�] �E{n#��or�e}�vg9�v]Y��VoHZ��+��þ��Q�6��Y��;�?��\�yKV[�z�Z��q���������vԤfsx#9aY��G4�Idۼ��z��ӳ��\�Z��`Pƪ)U^��Aw�k8�!����ņ����ϻr�g�q�iz�,���<����}�����r\X9Z-�KȚ��a�D]S��Њ�{gj!��k�u�d��t3DL���jօ-6T��x�c� �W+Gh�OZ���z�g1�E���%S���M����A�H�ұ������X��)6.[�Mwun۳��f�Nr����ޫ�yE@T�*ۈ���Ƣ��l[���Wn�+��ƞ��;7t36�]���Y�\1QW �:Y�P�@�J�6�O��:�8�vy:�+��Wo�[1�e�Sf
r*���/���T�G7{2苇�d��/%]m��� )[�p�����D
<�邠���v�3�A_�!��mm"y1��8��sr���c���e)J�:c���U&.'u�����5|c���J����r���ې�gT[cE ���=��Xs@,�B�$t
a7���܂;�V�����N���f%����X����5�h������n��AzV5k����:I}�Jt�5n���;;�'�\�wԸ�O�,�Z�X�U����F�f���9���r����\�eǫ;v�G�˅v�6�<���/~	r��,ꅽ�p����K��CB��F�bcU!m��})*�����%�����Pmc��5p���<aU��c[����{7�|���N��6`�h-s�k��;�|��O��@Ct)	A�:�s�B$sc]ò�1�l����kw6'y�\f��,��:�Sm
t���o\���F��f�MƵS���:b�:[�V���0���7&�����c]��[[�|��{�U����C��F�s�	�N�ff�3��Z1֠�8��yp�K��{K������]�~�L
|����'�n�Y$5�]	
S|΄�݌�ș�����QX���4�����q��S��&S��Y�#���#�u��C�/ӫ�쭸����%c�nW6�qL���+���S�At����[��r��}PTTsY�quwm|3ϯ��^+�:�4�V1
�N�t�J�U+��Y�-�QC3x���m�Ͳ�jД�����$V��H%%Y�m��N�x�^�*eur�\2TC.�Y�T�`����ܭ�j��F��J���4�WD�6�ܸ���Ḻ<*_gRW�Hp����5n��َ�9T��<��Q;,��������E�릂Ȫ2��(��z��}p�=�[��܀܂�]�Y3ؕ��y{�vc��\C�.�t�j'��[x��}o�٤�G��-���2Wt8��񏻜��7RW��ۧ���ֵ������[
1T�=n�Z�Xƛ|��q���\�@�R�_��Z�:���׻d�j��Ĳ]��RD�k����9P��EA�S����b�[�-�0�`����kk]�x�\�)�p1P�ĪF~�A�)T��o�:=E�B���oo,>eo��{��U���6�湖��q�T"���6`���UV9�}�ȻM���ڦ�^����;MQ���5	�֪s]�1�t-�Y��t��-OZb�*yn�\����V������=���j;{���rr{����+�`VA�5��_�#���C���bTk����(�}Y1�p��x|�e�<�6a{t2�{H�����<�U+l_uM��W9�n��{p�	`���R��;5D0�d�5#|p�\/3#�[#�S]��ܚ�{_d��[<�h�V�Ϧ�^���F�t���N�j��R��ֶ�G
�7��#�^��$YZ��.h���B�S��+s�|�����ͭJ�p�Y��~�q�^�jڭݭ�vn��3*
�|�'���KQ��^�R٬Ź|��A�q1�͋uoo����������~y����L����V.G6�p�ƻ�j�C	sx����]����U 7iq!٢�}�ʲ��J�����k�Z�p��C��_К|�<�Z��\O3 ��*�s��*h�y���wvUB�SK��|��j�
�K���JS���Q�q�T
y��}���Ԓ�-��G����<�͎�X�ӷ��R���8Ψ�\1� PS�|�~*@KE�����R9U���t��.�Q��-n8O�6)�{��:T%T�?������ϐ8;���g:M|�o`�F[�.���M�X8*�l�paXI�(wUca�6�g8i�x�z�۸�{UA|fVwF��6,�(��M��j��9i�i�9�)ͫ�K#��2��-�]�R�4�JY�'�BsK�����cYIF� ��)e�0��t�S%�ΡK�~�]+Nf������F�q�LH�`-���$ll�V4�'t]r��+Cvl_Gu���V��1=�2�w���u�I�+{���
���(�8&Z���8ֳ�{����ns�9��J��meG5^u�TQ&������\��J�h��U����5���cp1ܦ���eM�?�p��[I"4i�z��e�����!�ݡ*)���2�,�Q���sљ�n�f����ӷO��ݗ��]��MS��b�E��]Rc�f��n��"���Z�'V%�}��ܾ���-���x���DN�)�-�.'���x��ٕ;�I��;��Ee�} z�A8�phE�k�.�����$֕^�ݾ+,9i��uO���wsT�������8��"�D��,���Y�D՛��;ye7x�x��p�<��du� ��ld4(	��f��p�f6v�9�E�Ӆ8�Y��k���M�)�+<����&.��݇�+([�Y���wW�Q���^�*u6�� �3�u�;'>b[��ۛ��L�ry���G%Kb��chm)��*�C%
U����5̿���w&>]������5� ��Ь�8�Ŭ7�1B]����%��Q��j���n�ض�Cz�WY�x�G^Pj	�l�>�f��K��Vu��<���w�h�u�X�wvQةk��-��|������a�V�vc���2E6�����;��e��k!w�w����5r�P��l����}�6�U�W��!�L![���ܦ{B���rI����ٹ��]ƭ^'{�+8��PL-X�e��Е����)��
W:��n#�XV����	�y,�.�ʅ�y��;�-r�3c��o*���m�J���K��w:��(c�Os1ӱǆ�t�,�	�gs�vQx��Ux�ٟFہ���ס񔫞���Đ�3E�OOb�r��魌���E��VމYWv'�+�t�d0D�Ä=!�yI�i��^��KBѿ!vC嬳�e޻��e��)E�R��Ù����V��+��d$��޹]p��
 �
`��X��|v[ZhU���ήD^�ʘ1�x�J�!ܭ�����u��]i�Fi6����{-Y�#���M��������G�|Z�E�~��Lܽ��ګF^���g:�uj&;�
nā�kܝ���>����&�N��'t2�с�ڝn��ڇ#꜋�L5"��u���6��L"%v�������c���ف<�VeJ��7{��F%]V��e�Ҩտ��@��V�ɹ�+�Yk:L�Y���f�q:k�)��v�oj @Ka 2�T��S��M�=j�8���Dr�%H�Q�Ȥ�!
�Բs�u�/V'wwJ9��i��䘤h��EZ9�9{�wq܇,��Ԯft�e�3RF�r��z��;���Q[q"*8AT���U�"���,�ID�MNP�JDQT�Xf�TDfuK�!]D��N�]@�IΙ�=	�g*�s�qe:�h��1P�Md�4T���9Q:����D#*����$�1�!�Q�xm�:��
�\4�T��H��Z�j�R���E�ҍ��Ԩ,�Qr�3����j�^�+ʝhys�W�*�1�s4��r�H�5IH�w
T=ܤܼ�в���Wn{�� ����9�����'+:EQg��Zw.^��a���rL���iUku�w]�a�đ�)�ݻ��.E�HYY'R]��q�zR�/�A�e3�
�j�%7���WC������5fW�N���_t�I-���i����s2a������&2�bc'�$�t�+wyK/���]��5����)���T���D�F1Ũ�q��J�tԮ���Ӎ�f�m�u���u�I#J��NR5{v�<��e ���
�n�t}8����u�}F�L�cU;*��cs�.�#��F�Hq�l�-m@W?A�ۧS�Q��\��䝝픉�P�f�ԋ�q���ON�\�k���=�қ�g�5����,gA�~Ac�4.�SO�s�7�zdg�^�xq�̆��C_T&���&{u�uҋ2�^���ыz�U��.U��s�*^3��MI��^w���3* �팋��*�c���y�9�h��f���aG[���������CP���͙�I즑�/4<@��� ��N�m��\5c�ll5͇)�*��QW�uu��a+ɡ�}�w*��[e�Ԃꂮ`U;,�҄�\�بX�����P3E�;/�uj����p`���Ĳ����h2��)����9�괭�}.�VW�c\�h��b�ő���!f6DŐ���ݎS��oF6V�{g�hވ�jb�G,���B�ޱ"�t�E3�/�t�::*D9�3xΆ%���D��� J�ʵp����06`�?ʧg���*�R��Ã�I���No{���떂����/=���5�_
<����0(��IN�j�P��S��ǯ���O�Y�P�<��[�S�iJU(t�|� !,��fZ�KK6��ps="v���u�����_u���!8Ψ�le9F~D-�̶��ګn��k:�����>9ov"���浐�hX��-�3�Er�&�7������
YA<�j'�=�����+湫e�cm�t�wr�=ɚoR��?��b����t6�s_M�ڸ�N� �;�b���mv�ɭ�H�R2��L;ƵI��!�
�ufֶ��<��ǭ/�3R��1Q!1w�/TdM�{��Rz"ӆSq��WS�ȞbeY綌���_��è���SҚ�q�ky�ܫ�I�\bpʿ���w3����۠��=�����ҹ����w���L�z�X��o��_'o���;W6؇VH�^Wu��_#r�ˡ�0.�Vw��u T�D�ס�A_
|z�\����Ӣ}����]ݓbK�����`�'c�AT�sV�ca�����ы�5;,=P���\��:Ҷ�7���0f�L�v�ޫ=ۘb57��o�^OO�g�*�c�/�4=E&�.�3��<+iG&,�r�'\=�w�f:�����m�ڢ����ź��3���!�k�&uB�DUR������̯����T�V�P�q+39���y�{|��R�A �G���퍞,�	o_��8վ5��5�RQ�npbG��]��&�1�s{�^=�>��hk��[�v��X�f���{n�>�,����*1�oCyx��)���;�k�U�f�ėm�5����ڔ�-�ܹ��=�|ۇ��}o��K^� i�.BǑ�}n�r��t0���+�U��>��/��kZ���~�S�	��ՊS0�	��L�������@%���Y�uB��nZR����L��S�r�����h��0��J��P�y����q�U�Y�|ܡ�`|u:kx_u�"h���FJ�8��ŋY��uø��MN� ����{�^Uc\��m��=ȡ�W �Z�arܒ�ƒ��a�++�.��q�wve��4��Ʋ�ݽٙV�x�v�·1�����][�ێA��hcõԹWa���ٽ�fQ�\S�e�v0�FB�f9 �.
�*�M��Y<������]�5o9=����<6!���q����(�Cs�9���)�ׂ��*3����Z��W���圹�MQ��)���WS��5d����+勫k�y�b�hu���ӯ�^<k�W��^'���'���E�D�l�+\��J����̫=6�.ڬ�$rt�~O���Ƽ���WZ�u�vҏ(@Mu�N�V\��~]io�{-.ڬ��/����!�͓�r۾�kt��L��"�>}9���f:�x]��|=��m��� ��j����U�e�O0]p;�^$�\�P���[����u��z���<���P�vk�yE�B\5¨�������v��]����m���o]5�BW`���,l���vx��*�k�q[���\Bi���������j�%u��d����S3��돳r���OZ�5}]Z˭�݌�]E�:�n&�;�j5��WB�eCG�:3����bv�o��B�;���/�T��
�$і��:�!�йҮn:c9b�z����.Z��vIX�p�n���۝��GlW�T��Q;<]�u�T�T����|�x/3�պu�����c%�շ��C��%}�͍I_�h�t�f{6��A�%�v�,�(
�q�>���o�"�H[��T	h��f˲okv��l6��Yz�$e?��K/���ڞ��l\�9Fc���BP��sB f���{fҍBzD,�/\-��M+������CW
��#��,}�8W.���̔��{�j'�n����k��m�v0�|z���Ѹ�gK}�י$�c& �sֺ��Kj�-��0��5�`��=�)�ʆ>��f_V?3B��y=o,�ڿ�.����z~����O3�똔eV�ˊ��n�De��4�;_G\��g����jқ�����G��3hb��;�v�N�����R����p���W�Y�c��M�w܈W�x���;�sUȠB�W��-��c���E]�+�W�jz��0I�}���5 ��T���q�.ʼO�����|W
y[2��#]7i�L�ӱ��3x��K.*��� G[z_@d����i��n��(�=��[�p�ͺ��$��p�,Lݭ�D��{�Εw�#o[���vT�e<|��9Q��������ff�G�H�\g%b��Jm8�Q7Y!݅D�|�$�N���&���23�"^WY[�c���"����5��"����P��|�6.'��T��n����=m�+�%]8�����TW�U��t���r����l
쮚���ۅ�� /-�\��s�5��z��@hN�N�y�$uj�v!3�=�Z�ڼE
�N�e��7��8{P�{pkz�:c�0T�����S2)��Uyƴ:+i>T{��v���ko=�|2�R�|(t�|�e�U�y�U�5қݼ�[I���x�:�S�/��}�	�u[cG��gu+�N}�lSnOǁ-h���:��m�i[9�C��`k06�W'<Oh��Ps��`�U!rm�m��jys�M�|r���E<B��4�`P���*Nͥ���v[2]�sQ�Y��v�P�ċ}��^�����MP���Т۽����@��m
��������޵�jl��h�6��Y��$x���	h�E�#�Y8ޢ������a�K|�m��	\/���n����t��i���5v>�{/��[�_��w��l�:��%k��]�}ɚ�����=���^c�/��зv�$�v�w
�BtD�!�
ڈ������~�����۝\ʕ��zs�Ƕt�|��Mƻ�u:��:`Zܮ�蕢�Lu�C9Ź�Ӊx��'W%��j7*��u؜3�흧s���#Lm�6��l������Jmf��7���{~/c����3�������o�f�m��^�����Cf�G܅�4���d��w������-!bv���FtV�ݢ���]���ϙ��K���km�G�_�u
��]�[5ܭ�r�����ظ�I��ll�e�K����j�~�~Cِ(u��خ��#O1�J����Y��;M[�z'r2�*�'�q0(������T��K�v��T�R�n��o/}>��d/5�6���,�T��9
�L�= |��9ze�&vY\V�h����ɀ�"l�w75�4{B�.�v�R��hk�ܟf�W�ڢ�uޗ�u�e�n�`��k���IZu�݂���͗1�Q7�,M�v�g\��CMܫ�KR���v�e�뫺�p�9��:���u�M|�=�|ۇ��[�x��sd��(���)��ӟk����fƤ�1V;t�k�/��ָ�#e�QyJ����V�t�[C)�T()ﻦ �~)h�毂�Z�۩9]=�RwV����6���-,'��=�r�	O�A<�j'W=�7{r3Ѹ�pT��8������i0�51_5p����@фȋD����+�k�>�钵e5���6�s5��7�\R��������jw�]f-t��fiEP����ͮ[K�;MQ��&|��w
����Y3�hZ�|�*�<����x8��������~��;�z� 2J��^h6��罞��ݲ�W�����闙D����f�Q{V�bL�+�e��WK�����˵,}G�치�A�]io�{>�K�>n����-~��ȗ~x���6�#�J:�x��Z�<��%	ôQ����*�l5�-�7���ݮ`(�d��i6�B4�^ދJ�%�5e{v?*�'_�H�84�3��������oPz�]�Pv`4Z������L���V<1��&ȹS/o�'Z�'Dy^3��ы�U����l����V���ͻ7\�eAW�I���ۆ/%Y���u�'1D�ƙ��sa�<�k���ol�R�����^��[8��w��c�)�.�"R�Q�����6).o]'��n۾���}7��U�A\���<n՛��S �:YͤUB�Jƶ*��4���aؗ��`��(�3Y?n�UH���������o%xfðNL�վ1d� ��ͧ�Z�:y��E�cR]�G��v̀��o�{T��h��W�4i�k�5�uD[�
R���>���я_�bB�\��qY�*����s:����/��}��h��0��:b$�*�̇T�eӌ�R�=\(%�1ꅼ6�&���pT5q0��ّy��������`�����꽊�>���W����N��e�\o����W�1~����'х�&gn-<��Y��.gg��r��qo�z��|�K�<~�x'�8�:�O�0� �0�O��p�ua	n%�Z�+��ڒoj��K*
(]�V'w˺�L����]Ū�Q�u��Quc���0�8N[�nPc�D�ڲ�wS����2[y)v�:�����us���������U�2px��1�X��*'_��k��ږ5C^�<�T���]�$�\F3^��B}Fg���w�׀	��u �)d�a��z�:u��;]/ǯ7�À�ò�M�%7�ז��(O{��Uro=���?_��M
ו �d�`A��?V����J��T��տ����-�ݷ��u^G>����#ݕ���zrN_�,5%8z7�٪���q��V�/1~���x����\}�{]Q�D��i���)������M#�����M�4��$Ҏ!x_2|Y~�gFTN����,��4��NF̰)�x�߯��z�<{!��$+f&S�L����e�lNǻ���Zc���S�pωݳ,e|�B�+�U�ȩt��p7��E��_��zB.�֜�nשP]͛�C���s犢���MŖO���xh�S�WUzOS�C�v!ť{5���z�R���v�	��G�z=v��ɺ��Q߬�O�*a�tғ��1�����ˀ;�^m� �*�Mz��'>£�'�ۛ��o��^jx.�%R�	S_I`/�;z��������ѽ�液��!�bc,]N�L���|z��n��E�J�1��9�i��"+�w+k�p��o"׋�b��bn�eڼ���c�����Բ��.�=�E����֗ה-�4�j�Y��)�m�m�7o�
��U��0�����$��A|�^JL�p�=|�sR霪�3mU�,����S����M�=�}����Ҕ�Q�I�5�.�Y�	D�#zk��t��՜��Tz��CF+����˕�29[N����w(
���we�aj��46��ϯ��.�h���=纖�(�Z+�ۙ�K�E%O�+�e�]Ǘf�_*�ke|�P�����$"�u�i����������U���A�E�H��)�����zHẺ��v��7�b�{3d�b�M�����I�n���;B���{�:Va��&�ˍJ�髢����˚�+2��jN�EK�Os7�L�l^l�e�L<�Gu��G+zs�1m�Avŝ�n��͉�WQ�.�+���+�MTt���Zf�IϹɃ���҅�왃3�v9���V�7��;�����֞��Ww�QɊ���Ѽ�6��P���x.��=�	��@��x9�ط��u!;�Rd��;�/q5(�V����"��Oo��Ţ�.
�W[]M"�N��Si{0��9��̎+��r��V+�Z�c��c�=�6FP�H-�ǩ�݋�fٚ��u� pY�ഀ.�!٢ �z�$��� �١t�N�mrrk�3C�٫o�L����C9w��y9���S<dyh�8�<t�{�t��`6{0#Wc9���d��:�Q-^*�]�-G9���֊�v�0���2�u+=���Id�H.@��zRh桌m#�SV\���R`��[h���oTF��YwpoH4vS�)b��7�����sQP
�絅[xE�`檏.�� Sԋq��*Q_-g,Q+ax�{VO◐��w15�2�?T���JǕ����mov�hz�'���a��Nv�A��s�iC�!�f�`�Hس����!����f�=3[����k�YM�Ǭ�d� wk�HiRWXv���O=3~�A-��e�SZ�0��T�E�IB��KX����E�S�Gsv#�7`{/(#{���A�˱sͣQ��#t�Ҷ*؟ft����&`Rf3�\��@��DS�����y����ӌB������gj�͡s��C��	^���8:����g.�P�SvJ���3�2hY�\�3��r����E=������+e's�������e��-�≗lo$k&�8���pG�� �!au�
U���sډ�+��mf�D�մ�O�����3��֤�P-�)59�%��Q�-��A�Y��v���A�e��٩}NlH4��vɰfv�RSk�����3e�O���@��΍�����;2��-|��
��ӷ�T�-}���QVاX-��|Ɨ>m�j�ޢ`ZN,$�l.hrt��:n�����s·p�N�!kf��'3 ��aD���s�F{��j�%�2�ꑄa$f���D��D�.�R�$;�r�Xl���s%�g\�r���h��$�QU�BJպ^�UQE��&dUX��YT���M֔C�D�3.DU��s��u[�QE�J�Q3���7v'�$I�GM0�jj��m]�+�wpk�!$�����ed��E�"%36�;�E3��ZYZ:.QPQ�(���P��'2ç"+�hE�*r�$���EY�N�ᗐ�%QdXP�&\�UTf�a�GNa�Z�9F�Ȉ�X�*`�9n㬹;���"�r=C���	ӕJ�٥��Z�U�s͕N�t���!��i�������{7mν����yO9��ViNm)�"�>턴\R�d8����V_M�`N��q�fI����{z�;����\3Q���/�w��z�,dG��|}^�����ei��G�^yYp�w �(�x����7��Ȝ��1/|gD�[���l���P�ԅ\G�֑��Ӿ��_�iW�����{ϼ�ݥEގ3w��?~H�.�����"d��E�yי�t+|��:�3ӽ~f��G��Q;�o��MR��2=H�n�>�18��]�
�n��12�J��JZ>��:������r�O�l/}^�5�Y[��iH��D)u�}�ӣ��x����/�;�v�5����{���umr�&z��m��{�dW����({�Uro��xG���u���A���x_�beVT�!�W�͑~Z��;���K��9Ҹ�^ۏ?:�+�I��P�yv*8�&J>����qs��(ws��m�n���d�ۥO�����<����˅�߮ь�~����츞�VQ��f.�����V��+޻�I�,a;聒��:�UVx�ȅn�+;��^u���u��6����=�����}��yo�#�&���+�T���wo�0�_	�,L�֝�ү˩���7P�F��]���L��q�}s��������xq�Ax�-V-��1+�ܙ�4$���Q7����l���@����yJ���K�3���X΢Wq)�3Һ�f��yv�_dZo�s=�N����s��Q�W'<�%*��L�}����t�]��+Sl�#�xTg��M�,��a�SR۾9R�;y�ب��}���ŏ{$X����^��Iȏ]1�r!ڮ�+�}�9'h�|�}%�3������\�l�y��7�'޹������x��x�\{.�ϣ֯ó��K�$踷$�˸�3� zR�:�r������A��G\R����=�Xx;��9���9��_�����vA��z&��َ�k�<��.��X(��$T��X����]O���B��߇�!�|s�'ǵFmA=��鎹�����(�*�f�a\���X����۝u8<�~�(_���r�����373�ʷ]}�J�g��CJ�����S�v.K5�	Q�-�8����U*�+)�}o��Eo��7��S��r�2=;]����!��ċ؏W�&�L�.�#�+��T�����u��*w�j;S��]���j5�܅G\7�l��P>,�k���u�S�fQd�i�lܿg�Ob_�'g�{�����b�)�G��%>�Ɋ���W�7�O�>8}���:�&ә�kb���[��l�2&� :<�5��g#��n�=V�'�>�r���cW�S#3�����5���0,ӽ�7�ك�Ֆ����j�d�zt���k2�])]F5'N�o��{���.V�rek�7�)Խ���k�����:!�d+��j�/�*��[J���0n�����9�]x�>�3�\8*"s���ͿW��|�>7{n=���L^7�2_��o����ʸe�^ݸʷ�g[G����2Mq�*�L{�O��<��w�Η���xu�z��~��	�xl�^����\���S7��3^T�,�PɆ��}U��9� VF���9��K����QJ�ڳU-�{�L��nu��hOF��^��y��ݸ�0�k�P�"�/�l��9�ޘ����sw���%�Cj�����%�{}2�1�R���gep��NI˅,;L�5����A{����9�h��w�+�w�$�K*Ϡ=�IQ{œq��=���,�U�s���]W�&����(�؁�e�&|2�L��]J�b��C�p��c}^�^>�{%������P���F�O /Gr�Lǡ�T��֤��Pt�b몽&�:�K/�4o���}��طL[sw׺�����o�+W��1�����OQ� R�EuR�ND,ʉw�X��y����������
�X|#�����c�r&�P�\�iUA�p$�^�	���[�$ŗ�֩Lki����B�����jx�ar�Je�̊P/ C��.��ꝵ�����s��t�`i</X�;���K��ԙ�C�W�=�/�GY�xw�c� њ��奧���d�pu��׮B����,�d�|9WP�.�7[���i)`�1�y�f��Y�#�]�=���n��7�>��\U��~���y��F��*#nS�.j yMDK��I1�ߗRWf��P>���V��F��ʢ�>�������/�:
����M35���a[O��X�.�=\{�Y��R��>G�X8�|�G\7�l�Gޝ�������q�X���}@zjk��}~�2=�>S�n�Q>�#B�):\{ac׾W#��_��ǽ�g�q�x�L��Kd+���rԪG���ꌁ>�S&��=_	�^��+e�>�Q��O��,k�QN-�a�C��}�v�Q�#+�=�׌����;�� w�d�,��0��\�֫t���~=}������m�'n�f�ȟH���屑��7�@9���7&�kʐke��;�
񣜰e^�#�UY#��r���i���~>gyO��m��g�W������=�Q=���9l�t�ϣh�����;���}]����RG����㋥��u��d��i���)�������6��t*����v�&��S4e��'N����G�g(��4��NF̰)�x [�x���=��SQ�=�3j���2�G/��e堤z@�Ч�
n҈S݂���w��7��}3�E �ɇ����-��$�	�@�9���ں��ݘ�gφ��]bz�p+7�i>ٛ���4�u�y�S��v�����]�@���;�\�\A���B\������b��eN�G������."��|d����xVot�'{�3�KA ����w��t�qǊ�:�t��Y>Vf��S�>������M�����=�����*��n��h�x�{�ǖ}�<D�p��eJ7e�x�D��PeT>>@u��S��{�x���/�<ˉ��uP�z}���>>��X�?:���&낰l�JX%N�@�6�x�׏o)-����3k��u�X�}u>>�uEz]{��O�㑾����yYqi�_{c��9�{#n��΍�o+�
. �2ğz���l���N�HUǫ֑��N���0�	}�����:k�����3��;�(��,�( %E�[�"�:�;��W�Z2y�U�)�^��Oj�iYP���D3�O�����t�&�(��T�wx����Tn)KGݡׇ�v������m5u�b�#G����J'�ztx����%ӹOo��^#�c"_W��K���̫Y^�G�go��pٸ�b�.�\���xg���{`~��n�xT�ƒ�4=fǳ�VOk.�E�j�Y"��JZ�m���=���V@8��[��h��U�y�"%f��t����Q,��J���V���o�4�N-��9��-w@^�C�jnT�-3,
%�(n��v�w��憽<H��m�����tt�&��/�g����3��Nb�m{n=���M�?P�qޠ;���Tq�L�7|�\�gk���M�%��Y����6p;��\xOyW��>���˅�߮ь��Iy츞��w_�=n:�OG��O|��8n8�U��⪳�B�(�ݖ=�ε��\�-����),����_ajQ�
�������1K�S���waU��s�Sv���������V���T�2����׊'`�t��z�<{>~�Ǭ�\��,��a�S{*��eO/C�woNN7w��5����T���d�e{�}R���v��c��YӒv�Y>F�>5�z�I��;ảw;}�33o+�W��W��M��@l���<���=���߽���_�g�u�q�:[Ľ0~꿨Ω�22;؇2N�e���q]T�|2UK/��hw��s�'��r7��V}�w�ʊ�W�8�+��˕;ex�����e� �X����]O���B��xh���>-��rC'P�[�W����wΚ׵|fهb�P����K�"����#]֏g�օ	�(q����~��-���u�՜E�%�1���������0��8�ͿU�IES^g��i�7k!��|���7fP����Ȼ����]�ֺ���S��}@*�G����Ϯ�y:	B�K,aɁj�Ʌه�bvYdT�ow��=�k�X����YI��q�3��[��{��>�l���4�����K�|.K4��� ���Ӎ�#~}pj��YU9�uR[�嗊.G�l����z|�����~�8��zH��z�j!L�.���29���}��K��7���>�������n!Q�߭���R�����_9�f��|2ǰ��	�"aM�̻��6��},��2�!WJ��Yĥ���LTu���oޟ"|G� o�ΰ���<}�ٜ��(O^{*fCr|f|#c'=]��m��Ʃ�k�Q������~�$�j7I[&��'�DJ]�T��Wze��'!J����O��W.��W��φ����$�Z7��s=���I�9a���^�o�L���U	��Ղ�����Y>�0����gոe9�y��[�z������yl�-}�H��m塑�U�9��Wx�����B���e�wA��3&NY�왽�t��������̟��W����;�.g���j}w\;;+�Dg�$�,9�zt���Em]ҿ:{�'�ȷ1���L��(�.��ߤ��d�;�x�B�IM�7�ye� T�XddW�gt�pq��g&ұ=Yb��	�u���;�ʏL�ܻ_�n���Xw�+��f٘-�_kD)������t�!\8j�=�/z��6�ԉ�Sr����� ����c���cw&>�'F���L���Z��,d�'������ȗa-���k������v7��m�^>�{%���Z���Ǣ��X��	AN:�X�VvT鿯�A�(:�g��^�u��nz�<��"�m��Q'��]��@|3Н/��w��*i��m��}���^ /��~���s�Q.��-����E�K]ouc�1S�=��|<��9�����q5��.J(x���0�IJ�&�}��<���6:+�e���_�����|�|�>���g���:�
.q���~�y���w�}�y]��d�>|���Q��uG�>������:����������2^H"��I���}\w�Y��>��$L��c���Σp�
���m��ίx���7�	�a_@9o~��X�߰ѪaA�GK��~��E����[�p�V�T�֕�0#�C��2���IW~������>��}�����ɤY=P&azĬ1Q/��g�7Е1Ρ���I�UBV�z���Y��F{��E�μfoޟ޿�, ���h�����G��g�n�7qu�^a~�ܞ�74�;���.bӣ[�Pܻ��T�#i��NyY���M��R}��MP����]����
�횖iΝD<�vkWWG,��Ѭ�c�G��㻙�R�ST��}c�ֱ�}�ܝ���,pw�ku�L�L��C��$[�*�*�W~���l{��屉��N?HW���<mdШו ��'�0>7^1��*5&OpO��8�^���Y~�>-���>�W^s>��~�=.sݕ�ˡQޜ��a�sp7bys
+��ϸ|zxu��
g)#���<rK�εq��������wq;:CQ=eX�W�-�Gv�߫O�gQ�)��6g�ʁ���g(����Q�,
{� d���.����[�yt����!tZ7Ϫ;������a�����W��V���4�5�����9��N����Vv�*�N��w��T�P��.��}��:h2|���]��j_��� �z���赫�4������]�y���"މ���Lyz�_M�
]�(�Yd�5���G=�y�<u�Ĳ���T�ў��Ӓ���eĳ;wp�/W��O��#}`{��:�숛�
��VճԬY��f&v��ǡ{���N�1��]M�TϏ��Q^�;��2|^��=y�dnv:�J���[�{c�:�>�.� ��e���x���c5�j.�(R�W�#���/�3�ŉ��cݬ]�������>~YCmX��\�b\�@,���hc{�m4,��V�#���xHNC�p����$��μ�����H�ʴ{�
42ue	�3t�	N�}�c��;�w���IwoL����7��g[W�թ�p�k��G��dT9��( %_Q���H��μ��s�[�hp���ݬ�>��ֽk7�D\�G����Oi>s�çQ5�G�������*7JZ>�6t���cx��5������\��lg�ԉ�N�9��0�܁P���^#�aڮ��'���������.�Ψ�<�ߚ�������\�mׁ�W��66!��A�,�WAL�{��_zV���Vٟ[>�����n���WKg����6׶��ΪJ����m��{>yv<��9e�^U
&������{2d��N��O�\@���+����_���>�v�\&�U��EzK�Q���tQך6_�15ݭT��MyVQ��f�}��� d��·uU�:1[�J��=gZ��/�O�U*)��~J�۔T$E�{�:�e�X����LR�T������Q3t�S�u��f�j�u,���v�^�=����O�^߫<y�hn�����Rd���a��]��ymNϪ� OV^�x�}��@�s>��쁴����#"��zO�c�{��\;W
���;w,�	����CƱ\bf���"�����h���z�m�@���C�W�h���)��݇w��ĵ�=�;���R��dcV�3r͙�0f]V��nn(�t�������IsD����U˓�Gb���6�Sr!�y.o;�ik��+�8�;g�qޮ�H�G4m�ڧ��oC/e=�t����g��v��D&�ƫ�[t��o�e$74��!.k��t�;�u]V'��
�zs"�sV*�dZVk�|�]�ac,v���Dd��ΰ-�ɠY��F94�}��R\u�'���;9�]���`��D��D�C�y�ug:؍i�nPʓ�9ڨ_���hS&���b��M09�s��;���]A�*��z(v��x��O���$��]k��K�B��r�O��5����ֺwFJ�E@��B�LhX�(�����U��;�xw����d`��}����9V��w,,<� S�L�gWpͧ�FM�&V.��(Z��^�[��nsfv��Ydj��sq��f>�uN�H����:E!s/v�ڼQr��i��t��t�.�R�n�B�k���]{�r9�ށeԶ3��q-�i�K�g)[Շ��Kt���\t����aWJ�����rW��'fr���3鵩{#v'.��&g;68�QR�T�:�BΊ������*}����s��j�Ѫ�n��jT'�YY��7a���Q�#W`〈�oa->z���J�������>]+��{6��mv�z�K�Y���l�R�<��m��B����X������np=��U-�Cs�l��Ki�,������N�;-%Խt��Ōp�+R�j�i�5��Ŗd��ܐ/�?+���&�F䫷�1����-e3��Kb�sW��M.K��
6��i��l��<��j���8?ZUH
Q����kh�C���K�ڬ���:^��!��j.����XW��Ϋ�eZS �}��[��~[)]���1=��t"����"�ד�;�H�I�w��}�_gu�jv�.�5�bu��-���ެ��m�X"I[�[*�o�l�qu���b�+�H�֤���{��w���5��'ACu�V^,	,
z�֛ܾ֨�CL6KiC�gM�Z��Ы�{.JR��vK�`����Y����qD�כo�Nm��ؙ�`J�,�w�"���hd�a3o��n��3�ڣ���H�ΰ��}٫�^�ݻ���'�Z��W�2���E9Q:\��bƱ��g7s�:ʇ�Ȅ*���-�*�i�꓃�GL6(�d��\��������l���{I���Ŏ���wn-�FeC];��p�j��k�ڠ��6�ZYԶ��U�0��K�����P�Jq������vG3����}s�h�u_WIk5Ը�7֫`<�g
V+t�"�ut�Ԇ%܀Fʑ�w�E����u�yeV�W˟w^�&�r�A�g��G��L"LP�e�%s6!NxE�d���IX'��\� ա���Z�#@�L�(�VY�Ie�wr��\��������%U��y�F�IH�{��3�I�]E[!D��s�ʒ(�d������0�+�C�W�L��3(䑩"���j���eu��YHTM(��bb�Bb̔��p�C5#L�Qf�����N*sD��@X^��UVN8�M��"fU�[9��
45TC6K1"�-R��T��E����),J�����&J��U#ݮ�s��Y�Ah�f)mF�-,�R��O'=P�	�e
��r=wKB�4�J���IP(H.h��UOv��24R2���tS$C-�&rj$�d��c��ҶH�4S��'�B��� �/������ɹ}}rb亭p�Փ`ܵ�Ը�i��Y�m<b$RQ�2=zt���=�!�$�rwmto����/6{���g��	�F\}M���*�P{�7��z����e��y�W~���_�3(�ߦ�u���쓃גIu(8&ٟL�ݕR��M�w���O����D�=Z&�TL��8�Ww�E�5��li9 �|e� �.�W�ڙg���Wz�8g��U;cgͯ[�N|ǣ�O��y���fهJ(��)zdY�mκ��ϰ
����W5�^�Kj�,�=����l��}�U�*al��q<�τOź�v?uQ�f�v�=�(��Z�u�ǻ�����hdzv����Hq7��$ez��L�� �퇽���Gu�ӌX�x��<
+��D3Q���*9�SeǦx{� �k��G�`�ٟNߺ\��|�rSu{�D���$LD�RqJ�<1)~7�*:���M���O����I�rq�X<�q>g{����OA��S��^cTNy�Fگq���Qz����L{X�0�v�1�w4�D :Y������=X'�>�$�R�C�1�]��}�����q�?j��ڰ۫���]fR�>�.5��<���@��^Y^���l������u+�\*��B������+�9-J�ɨn��b�,�pv	�+W�u}hu-�R@�(�xx�u��#DG�br>�þ\A,�6�/�m�M����u^I����`!~�cۮ��g�A̬���O\z�P���H��,�W��z�lW��[�����G���9V�o��`��n�b�:��2<��>�~���<o�4){*F^�'`B�=P ����`�o�����_����2��8�X��.���~��9ϼ�o���7&�9��4b�1�^��������鎩�ӐK�(��p)��d�^>'�o�_�Gv�F̵̺�Ɵ-�kO����i�6K	��l��Y�WW���:r7�C}^�n���y���Ʌr��*���|ٿC����X�g\Ν���2�����Ϥ�9ao���5�w��ӕ<z����I�0+�|:P�?S�Y��m��1�s<v,�OT�	>T��ʟN��hx*�;6�=��EdU�&��ܱ����p�x�o�u����970�T�5Y'� �(9Ͻ2˩�j���(�v{�ȯG�븟���+���{�|�do�#q�TF�:��d�?l�j�E�cSx�wb %>���&t��-����Q��y\Uǫ֑�9⴨~�
�ޢ3��1�v�qX��ܨn:��uvqo��~U��@teӅC/��j�W�Ӻ6��
D��/�g��U^��\���N�A����Y�w;����e���}d`�٧WTx��ǏM�^ef����˚���,��R��
�C�Xdδ\�J殕rp��������g����@�ARD�U���e3�΢�LoC~��g�z�̙y��6<�@1J�Z���Jd9D�7j2���2)L��I�㤎��2*+�w�j2ǯ|�G=̕zm�����êk�Fz�z9?Y�ȃ���=Q����>'XJ�����j��|�nSί��Fz�XOoד�i��{�B���w"�^&�ޟ�u`���K'�C��P�\�-{� �3^�|�;�[�������7�4k��	�jO���so����\ЭyRGK'�=��߭A�g��U*hS>91�)��ȥ-3���n3�..�{�������b��C������*X��i`_{]�����:jOp6t;����R��8�_��Z��D��i�~;�#.8��}�U���/�5�՟�q��F��X�|?N�qU�t	S���,
��Y�߱{�.��=S������>��g�cu�W�3�3�x�wA���P�����@y����ӝ�ױo\����p"������z���wHwy17�S��}�f6�Or�~M�bT�~�eL������^�"��W.����6�v�S�b�s�ton��	�d:B�q3T6���(���l٨��
,�ע�@�|u�]��!�O�Q���_��fn)]0�
vݹvp�-����K��s�������5�6l&�!�{�_F��T/���_��s��=�#��}���Ly�z��u�ǔ��:l��l`+	l�ɲ�~{�|?|1�C[�ك�W-��C�w /W�����g��?:�쉺ળD:� ԧRk�/r߯�J��&I`C�@dV�E���S�z�Q>N����O��#�r����,d��u���s��7xa�_�oǬƔ<��%O��)3�W[��HW�ԄN�z4�L�T=��e�p������U�pw�,���䲠 ��Q���H���s )�ŷ��=R�X�Ry]Qu�=��lgޝ���~��n<��N�j���Cpx��^���>V꼧�����3^�=��W��/��c"=>�O����:z�<O�!x�Z$�՚��v�3֥z=.��r���J��7�y1QQ	�zM�ۯ�� ;��Il�s}w�-��^��M���cĖ=g�*pWӋ��D���l�+Jk�q��U%F9�����P��B�8.��w����{G��j���2,
z}�GW5~�>�{�˅�߮щ���<-ϼ>��P�]�r��J�ʑ6�!7�*�����P�r�-�Ճ�韂���I�V���;?Ln�12#�&g�qۤ4����4��.\���.k���q��'ĴeDVlg�9����ͫ�5S���D�V��!x�R���$m5��W�橽3��tΩ`ǔ�N`�]�K�8n4�}P2c� d�S3���%g��Ǘ��5���=��U{t��E��h'3��}�V'�kJ�������3�wLT�״�y���mʪ�z�n�mjs�����@
����ϥ����g�c�X�=g�g��T"�̸3�}?~�)�Ӡ�ќJ/���O����(�����=��H�r��>��i�^UÝ��:rN��WJ��X�Ś���zIcĻ5�ۭ�7�.gz���W�l�k�e��y�W�}��c&�1S��[(��Ϙ�>���qjI=Q2��0���e쪔nz�<�ޯi>>�fo�v�M5���s���7�j��A��H�(�/I��'�|�\���mԲ��
���5�7[K�֊�bǾ�
�/�'�m�\>�6�;�\�k�D*�,	�R��[s}�jB軜^�[��q�_�����C��V=�#ގ�*�=P0ӥP��G#���F|!��B�=캧j�ߡ�;�'�O2�=1��}�qq�+C#ӵ�ߟ�&�ޒ2��Pf:d�����گ�w����Gh9�4�T!3[�����6�Q$P��P�U�r��Gq� ֶѼ�:�)�T�Ƒʿ�����Kqj�9HR��xﻄM����f[�_"���]>Y���!V�����Ino=Y��ֱ'm�p�h�3+9iO�lp��"�� �Eb �0�索B�z|��Y��n!�ߩ��3��9�^��:�*�y�3������}��۠5���FY@'���;$�²)SG�|���!Q���o�z|��A��( k����R�b��k�W'�u\L�_�K�矌J}��T��5�h��ꑔ!�c����-��Ƥ����>���X8z��p�'� d���1Q;�z2+U{�߭�B����m>W���Q�}#}�z�~��~��y9�;�X(TF�����s��[��4ӣcoէ��pm/~MB�է�~���z��g^_�G�W��k�x?tН=��hT/eH�,���#&���FT���]*q����qU��d������^�߆D��o�w�~��9ϼ�v�B�:�>�^V!�m+��}�����PTǪ{.�J"ˀ��߆}.W���\�z�B=	���q+z���E߽X�F'}�O��L��&x+���f/��󑾐��'��P���u�Ι]E�xx{�w=��]n�y���a`ٵEp��Z|#��#���gGx	��&�H����<���8��3.7{��4�3|�[*jUtH�ǴŴ�퇺_W�nz�7dK@<��8��G8(Iu�[s(�͍%Z��"��6mu��9Ö�]H>�k�RZ%:2l��	�n�����;J�-�QB���wR\G�z�5�_�z�z֘�ܩ�YD��1�0|���>����V��U�̫��D�\�eD��z�X���z�d{���s����qɹ�_
�ǃ$����F�; ���ݖ�m�%�������ȼ��q>7�u�\z��Nyϙ���*3ʈ�uL:�,{������r���� nMJ�$�L�t���5��Wq���r=3�+��N�q;�b����n�t��[�;�{�7�i������ �)V�p6W���s���Q���1�?Ǫ�Ċ���J��*>H��{Inb�ͳ"��^����v:��>�"��w� X��F�%����:�:����k�6��!�d�1p<�Ԋ�Y=���/��}�?z��O�{ՙ�gm(�gצ��L;����o��Cn|O�X�� K�Ԃ�'���G{�(�Y5j7=��V�=�����b+��׽Q��_���O�rn1��s?_��\Ш�yR@'Kʲ���ܛ-_�=ĸ/O��è�W�s�S�|��q�μ��k��9����G�쨞���Ҩ��΅�N��r�3���a�A��Vu�rx�Y+=�.Ľ��(�0燗���P�谯S��c*nM�'s�\�x{1` ܛ�z�_^_p��rB�1i9�+�����j�	׀�vҮ��N�E���6^����,�|���w�m��n���G:$��C�3d�l�<jO��l�wU��j��<rK�:�ǋ3�>ދ���u�~�V|��E@��~~����zP���"0�D����t;���:0ү��b���;�P}�>�:�ls���͔��'`O{��s�]g�c�Gq�X�_�� �F��kg�0e�=����`�.O(�Y���HS�^_�k��s�]?���.�o׷S��}�aa�#��vIe>\�ו�d��z}��߭P��؇�7޲/������<��&��\�$t5��FCX�D�>�/M|g��iI���U	��z��"=�|}��i_?:�U�Q*껅L��;;p25�����d�R�$Ԁ����}u>7��D��N��#�O����T��F��gxݾ�Mz7�q���w �(҂�,\>��E�W[��ԅq��e�^{��V߳m;���>�OJda�n��T�S�,��	Q�1%��,��|`_�w��\�r��#�/�{�����zw���������t�&�(���<Ld}���P����5���D��:��+GQtby�r8N�0�tn�z�b*�\a����vk�J�ϑ*�48�$wwiM[|71���Ǔ;��:�B��j�R�:�{��4�ⴖ�aU�����G4i�L���w�U|���p����P��Q������}r0[^���z}H�`���>*W Tt�}��x�U��;H�ώLLAJ�G�+{����W��6��� z� �c��w���׽V&� z���}�tQ��!���;+�l�>�����{!���>�Y��鞜k֗V���'w=�#�k�]�̔`qP�ӁOO�����>ޟi���¹�S
܅w��Q�H�wf=�Q^��=��#�tk�/������8�U{�B�(�/�H����Wi%��{n���^�c~~����V'�lE���3�d*���+�BG�u)����ߴ��gz����`
�/|��>���7?Vx����=�<3�2d�����QU>�J���\c>���ۊ{w�*e�<�mxO|��3�+ޓ���^Uñ�pq�R��|w޿ܸ�z�]7f��o�a�|mS��w&�nz�@�L��)L�D;�L��0�@�2ڡ��x�Ìs�J�u�ۜ^�G��D�t�0��Jz���YU,�ϽVD�x��3���>��8���#�TJ(#�ۭ������@�3FǗ9�zM� �������F��%��t���2
���|f$vj��ls&J�緘�u�̶�.c�Y:�ALݺI��Q�O�1��'\m��\�fE2������;���tn�=�W#�[�����x�S���3|k�{�[���|�Ԯ|U��3�<�ڽcw�s�k�Sf(��z=�hpϼ�����Q���q��a���H����,	/L����U������c����*�=���8P��Oף>���+{�4��RM�u�%��D)�������{u^]���ט�e"n�"�C��ny\W���^��#��Hq7�I_z��5�����9��s�꾏a�~�@h�rD�>u���h�w�j5��m��>'8���uh*��W��
�����f�X+W�?hSzf�d�������D��HU�R��@��B���5~���q�^j�ܧu�=w[ιH@{h�>>��}��bә��= �^AV
�u�62>g��5}��A��IwQ�ol�I3�g�2��{��L_����7��{"`>� o�<�+҇�*c�E/�s�ñ,��fz���o��Hu��b~��x�C�u׿6ϫ����h���t-W�����𿲷ڨ5ъq�6b�n�DW����ח�u^㑯�<e����ｓB��R3b#��6}X�ۆ��?]����Y֋�M;�2�+Ք�ޛ�O]�OgT�׼
�IðB[�S-x��Zp�ap�j�so�Xb&��]�"��@ǘn�ծZ^�y3�]��5���i�Y��$+EF(��95�����Ș�:j�����������]-��.B��S�9�R_
#�v����b�i��Jn��gf�l�]�*;�J���oWWWL6g^�UԎ��w%t	�����^],9��	����B�K�[5���G;v���Ͱ�v��Ǔ��&S�����k"ޭܹ���Ӷ�z�wBn���smV�e<��m¾b�-���œh\R��x�^�YNs�Pf��s#��9�˱:��gl�bĜ��#Ԕ�ꧢ��y��,h�a�@n�qԨ���O�`Yb󻀴m���8���ٵ��_Hʼ����u�9m�,k���rlY4p^�%^��u��'kxe=wӶ�3 ��Ԡ�2!�X��'U=Z�K,u_ۋ��Sp��O�n�����5ة�.Z��Ǯ͕ʺ-�Uܳh�>���+�t�e� UY�w|��@Pq�mr���b���ǵ�]YiLe���7)�&��ҷkzŧ�V��!���T�K�&�r�#�.�&���ࣩ��,�z�bΓo�H)�A(r�삛��XNw<�m"���WMT�
�����W�<�e�:K��7�4��|j�2_T
J=��^ǎ��i��dB>n�wq:�o���u�SNޖ����"�5`4a�`�x,�
Y�Y�\�I�"�{+���T�Rh�vO���³'��B8]�Ƙ��7N���]l�/�P*>̧�l��9�E��9YB���9֨.��j�Xz�:x���R�;����j^]8�p�aj=�r�Ӈ8T8������n���.���ֈ�pK���m�c�S�����R�U��1�&�l�*�gS]�v�ܡ{�u8w ��˥���a�W�=�#4�%݃f�ڲj�N-7���:U���}����J9���NY�5Ť�5�	�E���PɩQ����̛�4�u�AGv*#��e��4g~m��t}� ��&�7�Խ٣c�,��k`ÊR���K!}u�3���;�n�ܮ[��F�7�������+�O�٤.��٭�T�]*���[��4����l��PK��S*���{�9�+��r�ƀ#�x��0r[��x8��mڕ�؀��Ccw�}Z�K��(a��o녲U+e���o{��oN�ك%gvY�T
��pB�<� �	�F�� ԛ��k���y:���y�s�Er� �wAe=-�V2����'��C�G&U^��K�u�����M�����J-ۡ���A�ƙ���ξb���Tq�9�t�X�#4�n���/v�u@z�h2�L��6�eh9�˶!�6����:�.�i�%Xf��AO�U�,zw�ݩH���a4�M4�M�8
�!�Q:�p�в6:%N�(tO)����S̜Ȣ��]��U��G�UZX�E�"+u�(�K
Q�b�h`���ֳS�p�O3���3i�K���d�R����^N�a%��k2�8��NZ��aE�{�������窅��$�d{��DK��Q�rqfTF-E]Ƒ:R�誝HrH��(��w\���G�n�V'�����w
�R�4(K[*U��".ViY�T$������R(�'NI�6YhEe)���	'��!Ai�j����֎��t�=-V��'�G�WS�
2�9�JZrK�ۙ�����x*&B��{�zG��Rk6e)�ʢ��bt�K�O3
(�4Y)��H�2�B�µ�n����K�9�������Ҳ�LD�c�C�uAB��Ӛndo���X��v�u6mNQ]����y��2]�CA�]orͮ�,(�Y��r|u�tӢ\p�=��T�V���r�]wºm#�%��xw�0��-#�2��8�_��[��u^�L��Gy�G��N�)�a�1�W�����}��-���P8sO��t<��˾2J�(�.�*`z]/T�0^�$w�zv�H]�3}��uL?����J���ȗ��	h�����i�����/އ4B���>W�:�s�����@��*�>=t�V|�\wd7|i��Xd>'�J+����>R��� c-�oN��BY,Q~���<��������O�dz�p5�7�]�(�d��0�O��J�bI�glVUfZ���]���NT�*%���X���^��	�������L{J��ࢉG���9���dt.�"J��c`O�����y��|o�_��.����O��}��=��<����3�l��RW��+�פ?d����j%�[�[/��-ߕ�\z�i����=����T�����v��B��E@cM�;�dmǦ�e�9
ET��-�_����Hvo�cz ӵ�����V��"�Zc�w��>��|��fEB�+��n�u1%yM���x�?��&�4��jS�	^��ِvsx>��nz�ٮXR�]�2V<P6����>l\Gma;�)��.��.]�"��w�QA��+�v�y��KWu�W#a��z�8��5=r%�8ծk;���١�Y��oR��լ��)ԓ����f�,�Ȍ�ޜ�k���9r���1�z|�����y���H���&az����x߽�T�g���X]}T}�zW�o!����y܏��]ȶ�x�dO��g��??]H4���z�'�d������g�ʊ�n���Kg�#z�q�����W'�)��g�*��{��z���Fn��yv]zA�zp�����7g��w�r�Z>g����u��o�ZWѯ����ޭ�R��r;�{7,�)�J�g�_F��Oؼ�6�:X=>n���G�J9���εq�ƺ&D��t��������"�vp{��Us/|��z�Vi�g�3������gC���:0ү�������{�:ʽ�}�����{w؀>~����~��7�;=�:mN홇��"���x��s}���gvy3�z��`�`T=��ׯ�����t�q�y2��[�m�ݕ��NR�^���L�&:����S>�>�ˊn�M���z�C������zv�(5�]��&��Լv����n��v��2��Q���UxϤ��eP�_:�k�ޯi��I���G���H���ߙ�p����48�b�)Wuj��R�ݪ�2��J�:L%��T�er?mtƽ�Py8L17
�}��R�w}��`f�7��ŀ:��Žت%ǀ���_a�Mbu�:���pD�W[sym��y���R�a���Z��+�k�Q
G�eR�vy+�_`˕�8�
>�~�����6K�,x����Sg�!�����4+�״�w��꽧o'� �����=�T=Qm�p��|����7���k���ݾ�m/L�=ԶS�ꋯP�}���"=���{�a������Lÿ��f�A*>�&>��I�&O�4��Y~���W�����
�޴8g���2#ӽ~�Ը��ި8j#��@�\ ��b��kf��U��[إ�c�J�Te���F��Z�-�;c�҉����o�p
v�@+�]�.n�7�s��K�W��K�26\�{�Q�R��Į�Ǔi���{ҁ�� ;ֺ߰����#����L�����2���N>��V���-�C^ۏ?:�7�^�r���7�vu#�8*&J{ k�{.�}��2Q�T�,oDN=+������z����vG^(����=͟c�Ew�=�ь�}�Iy�=q��:������Ɇ�gC��a�n��iVA����)���#)�/����xg�׻<7ʫ�^��f;w�7U���]���}?F*� �5E�8���ܮ���^C�v��|Ry]��ftud4lWWDc�״+�za�)��:b������L�����L+�T7���~8"���
}97� ��Wzc�q��
��&7���\���,/�%ʶ�'�ޙȀJc�̦��]��J�w��$s�P�f/�U���4�����
/|��%ׯ|e�w�?���q���ʑ�;ޡ�&r�����}$��1�G���[w�I~%�O���$g��{�r#�Q��^så8��t-��\z+Vt���}�˧$�,�0�g�3�
�w'��e� �o�ĶW��)�=��ï�DέU����7��\w;�;:rN��I'�&P�@���+��2¹�g�z�?rf8_�BT����6�� )�>�*(�9����G��{����2�ےQ�"�}]J���=����ŗ�~Z�"m͟z��U�;���=Ln}�>=o��݆o��.J5���������:�*���i�ɐ����P}~�g
�~����V��iY�@��t���,�_��r	&�ͺ����v9燄�t%�d���݀�5}�qW���2=;^G����������2D�zO�ݭ��C��U~�>�����F��&%��lt�}��j7����M��[*w#q����MWv�R@�7k ��M�4�IL٩l��"e����M�~/�r�j���&~�K�O���N�".���U�Em�t��I���-�j����Cg7?]$��ֹ�[f`�A�)%2r�?,}Y|�v���57�+��:Q����;�ia9�j�3`�5һeZ��:�j�+�Otn��.��{c ��l��J����i)��R�O�A���\ә��=;�뀫N:����}��MfMk�Wz����wQ��Wrb�m�̛���;�l���&�d�a��}�1MF��ٛ������ϣkk�=^u�7����޻��|���c�3���OZ�+^T�Q���B��sN��o׳��u��E?@�F�;�9��缯Å�^_�}u^��<e?u��7ɡ�&��o9��`]�+���O�0r;v��V_��_��t�η~꽾����O��K�	�Q�i���h~��D<�
�9'/���C��}:�e����Q�;.�:����ϩ�[*#���s�=����Vq�>ɝ���;s,e	�
��xdt<���ۯ	�w�Zk7��� �7k��z����K����v:�c:�t�d��b�(M*��S��g�ԥ���C`ߺO����`�Vo���G��s��~+#�H{��]s(�Yd��#1� t���m�r��S>�;\.�WJ�w1-Ӻ��^��p�x�o�u���~�Y������5f�_����깛:X�ZѦ����d�ty1v��wt'�v����m{��>=�՞B[|V�rT+dX�J��y�wu�*���R���9��=�ʩ����ԇq�G�鶨�����#��Qm���}7h���e_Iw2��jKt�e!���7b�/�ߊ>��	=Pf	��0.��/]������u�>��=���=Ś�WEFw���,{!��_�j�:���) yMK�& �^�-���ƣ������H݋�﫢����VZwJ�/���iW�{�F�zi���24��UO���끸/ō߃�E\��M�fûݐ.���w�:���7ޮ��dzw���Oi7�Pr�S2+�2W����w���м`��z�^�ݺ��ͻ�
�����x����u����*>,�wļ�F@�N�Y=�f����;#���'�z.{��n|�Ǣw)ќ)l�%^��ʪG6��� z|{���A��q��*����s������<Ip�>����qu���x�����s�߆|������C��><4˨��
^��k�5�S>���,����vp+��_qϫ���w����^\,��]�߅_��w���t�@ ����Q=p��W�9l�|Fa���/�q]4J9��{�yK~#�ޘˤ�3}Ot����{
~����w���M3���h���>�l�wUYgF�"�s'�e
�F��k��lnI���uK�6��Y�Q;[�z��z Nn,:֫v�Y��>���;pr�Uƈ[�2���|�]1t2�T����c@�����6���;f1��M�0ǆ��'_B�gݓ��d�
ym#�\#JwhW�ʝ���S�)jS���%�:@U�Y�}-��Dz�<{!��wg�Y�7��n1��c+�Q�g�:�Vz8ߛ3��s秇���~9�@7�� �Լd*k��}R�y;�;�C��Y�S�נ��w]��g8
9b�^��<4eTu�r��}n�n;�B�o�d[�^��zX�~�C���=s��ʜ���g�-���(�Ą�U�k�Z��,�C�wz���O���[�*�&�3w���;��5s�V���7\���O�'�e�#ʘWSg��L�����W��u�gf+�.*����2��]�G��}�#}#ǯ<�d�]�6
5
UX��-�;�
T5�\����r�z�$_��=}HUǫֆ���[G~�Hҳި9�z��v.K5�C�@�N暙����lZ�}>�R@g�NC8;��և���lg�z�;~~��߽Pp׫�P��\���;�-�%l������/�p����Tn+������5޵�47�L8���>�'�� �,�h�M{k�+�_k˟H�=8N�!#����}^�qJZ=y�W��Ɋ����Mǽ�@������>�N���u4}׸�^���չx���6�u��`�>�u��+X�X^6��̴�qY�3H�q<��2sz���:-�����N�<f�ZB>M�Q�݇)��{8U�N���J�Y�kvjza�,�ˠ��"*퓱" �V3�>��� Wl�UNLҟ ̿���q�p�����q�|Z�T{/�����솽A"3�'YL�-�_�yv*8�&J0ʝ9,u�NEu.<2��𸡗�+ը��IX�kVW�uhӧ��ˇ���c#_��%纨O_�(�vf�id��L5p6�?Sѱt��{��'�|�����:t�{��u1�λ��7^�������V'�k뙳������>�ugJ��ە>�~h¸���9�p=�.� ��������w��:��s����nv�ǾT�؛^V'�����:�D�=qKn��EL�����?\�g����]F{�^�Ͻ�y"�m���������~���z�g������+]t���FG\�g ��p7��j��1S5.�ɗ�� <��z\/�z��vG�Ь��p?N�%��	h�������x�<����{�*_����G��r���S���3|P�2�ےT`L�X<��=DQ�U}��tNW��<ʞ>�4)�W��}�=Ln{������3~0�\�k�|ISއw~P�v�"�MĥduҘ(+o{f�?��귴۩{�y��2�O`�ƚ8SCB��*�rk�8;{ܦ�}.�+"X�9���hu9���ڱ�=�{Mu5ws��j]�&�ꦶR�N�P=e�'	��Y�w�񾭐s�JNOB�m�9�oa\��R[M��szd_�ϓ�u0|����C��X;ϫ̮�=~�t�Q��כ�3�n_{*�h�<Dڃ( <��=+��Q��>�O�����y��C�ʉs��_x���>�z<�'y����ʩ���.j����2�p1ţ�P�F��	���m��{1dj�V�1N���]�������+��3P�I^6j[6zH���B��T����#��(��TS���c�r�R�Y���׻]%���}Ӿ'��	��9���Pfaz¬���}� ������[VՌ��q���^�*||�$y?+�0��+ޟ@�9�7��d��Y=_�}�>E�-�b0�`�8��E�1�v�8O9zm�W�\w��0���(��JW�/�l�a����>��B~��f9����������
��G��8�~.3�/�>���~��/�V'O��C��	�.�hIQhy�T���'j���;�g+��L�'���_������g�M�x�Wf�ʤ����ϗ��wn�lw�$��7����ӡ�Ue�%x�_��|������0nOԆw<�L<�H�����(���]hyVeM�&0��<���(|�hP>���þ��2+Ѷ�y�B^���+J�*(���d:�\��ocy8^����q*�:�hw�����6[�կ��z���,�]��V�2 �i��g(=�9���R�8�g_�]0-z�;,&]g}��K!Vq��мN%�qg�����z�UO����E(��>�8�Q�X>��x��]?��\wc�F+;*tݖO���3focXi�~{o�+��Â\ʓ�Z�ˎ��ho���z=^��O�dz>�試�m���f^�l.d��/���r�"N���Q}L_��J}92�]÷�!�����'�;���o�Ǹ�5�̟(�nfǫ`(�r��
(�|�$��Ǡ)`dEu0�������*�N��<���;~��z�EZ��
�àx���u��w �*��<��s�cKe=ucQ�~W�^���"+w]�W��P�V�zg<}�_�iW����2��C�� "����n���X͉]Ygg�~xݮ���,{���C}���ٌ�N���>��oΠ�}��
d�M��n:Hݪb��=�~�ez���=*���ʼ�0|<�|�Gy��a�z|�����y��2��Ԁ������C����̣l=��]�)?��u���o!*�Z��bӪ"�IS%�-?O�G��6m��`�1����l����cm6m���cm���o��6m���cm������6��0l���`���`��0l�|��o�0l���`����6��`�1��S����06ߘ�o�����)��&*O��o�9,����������0���<�y -��4h(�`hJ4 �@4jlE���TDwP����jj�����&�m�i�klM�[U�0+5d�,,��֭k`Q��ݕ�ͭ���m�YmP�i�V�ɭ��lM�ȩ�Z�ѥ���ԳBT�'-T�Q��  ��n�n�N��wC!����q�����c �`���B(gz�*��#��>  �}J%��SM3��#]�p   {��   s   ���  z��S���L핃�i�W>  /�qlb�[w]�ֶ���ց�j��q����:9�Y�t\�i����LؙU
�� � '��h2�4�nT# N�hZ��mr�Nkv��	��<]Uj��P��[T��� {�U����	�j��ӝܪ:h6��AkU:���3*�Pv�vj���}���s��լSY,Xz�  [�V�mL�OY���of�un�d�])���m%\������uM���J͖��ҷYl��5��Sj��� G�����h�U&�s���K�F�r�E�n�:��ڮ�������p�gcZ��%M�sQjնحJ�P� go&���N�V0I�fУ���[���݅�Э�����J�]� �M.��p��m�mV��I�Vm� �^�7s��mpDZ�(�`)]�����5��΀��ܜ	�]խ��t8��< �ޝ��٠fj�n��]��n�i��A�]g V�fņ5��s��      L*RJ@d���L� ���0�IT�4 1 2h!�2hE=�&R�T�0     	�A�~%*U L &  �	S�JU&S(`�h�L	�@�h�CL$ �#"i�#"d�@�Q���mI�}�̷�옵�߷���ɍ�[��s���*ٜ1mn�Z�(!̿��(��AA��(4 \T~�PB��H��Q"��۟���?��
������u����	"�D"Q �hPT���H�q��-@
�(��`�g���^��������/��(!ϱ�Sl��o�~e0.rj��۫��b�AE$?w���叝���U�T�j������L�R-[�)aa��:E�.��de�X�T�^���L2	Tƭ؅|�ya�o3ZW�Op��S`�,��kS�չ���eH�ӕq!teQ�a�r�Q�]�V�uZ�}�Wr�����*��Wn�[��4�8p���)`Y��M��5�ء�T�o%-��lv-dffoZ�Z7t+Jz)�4�0��Q�u��]-ĳY̰�Y�o�r�%0�,�b�2�i+�FJ��e�X�� 1���ࢷHASJW�)'U��{z�m]�&`߆@X35h�f�s-nE 0TU�~�
�w�.�#ߖ�vF0���I�]A2�����Y���.�-�,����F0������/�a��c�mj*A�%��a�&ܫt�$Ck4)���F��+�vf�l��eP���-���U�W��VX����s0���V�.M�1��lhц�]mpΫ������!��f��}�l�!ϻxi۫4����� �v��ĵ���V1i�*-�Xʺ8��j��,Ed׸,�R�,�V�fP�W�Le�x��Z�G�^���טiv�h��=�;6�Z�o1Q��r�x�Ӡ�p�	��9�j_L�j��%�Z��lZԬ�1Gh� h�s�АV��F�F7.���w2c
`1k��k�rUGVrL���Ն��^�xE��mͤ��Cr)�h/��$�XOǖ�2���A�"�	{Yn$w%ừVVҔv��˙�NU���ђ��h(ݶ�#��J�
�y�qX�g�2���eX���݅˒��iz0\�V�Ǣ�db�vU�yw��B�b�2���aCn�\qo���/)��h�,П=d
�w�f��S{�u�{��R�-����*EASWAr7�,#1<@��3/�=
w���n�Ȅi	N4Ki��K����&S4�1�{��	�D���ǮP�P�E��ZU$�ǕN�,�/2-#�.�FEQo!��'UF���9�#�s�5'p(*fJ�(��ea��\D�aU^�^�"X�f�����J'6rΣ7nU�U7V�Fe\d��8ؽ�+]���2@T��+8�u���Ƶ���Ֆ���4���f�r=Pi0�9_=$��k����XE�����YP�925��a5�ܭsqV�u�61%�cF�x�F�khZ�g��2��[��_!��l�f����f1Q�Gs(䷅jߝ�#%�M�"�yywTf+�ȑ�S�U�;��DojMf����6溋S�5?�f��b�K��h]	*���:�Z�6l���Ɍ�Z��xwrKj�;;wZi���`��Es՜�j�L��)��:nf����7�M̧,e��vl�,m�$е��T*�N�ڗo�V^D1�6�ݕ7ICM�5���W��6����fg-���+l:�y}�z(�^R8�5[Co2BT/��1��v�u�M&R�u��v���ws�l�2U��u$��d�n���zi,f�y�5��9�	*�J{X�:�Ͱ���	i7�Ʒ��0I���5�a*� ����z�e�6���J`Sf����7���	×3ַ�����@ӷF��5�wZ�YT)�GV�f0o��t]����,h�V�`��=�Vrmn���q۷&�)#.ֽJm�+pv�F(e�sL�)�w[���1,��B]��kv5I�R��\j�b�Y�xL�ʵ�.p�:y���"��*��J��,=$rd��7iYڙx�:���&Λr}����,��2qa����a�ҡu>g"���˼!ED�AgB����+k]BX�a�رŸj�v���^��eϫ0��[y��������ZV=��ST*QR���wuZT7X3�yђ��:n��v�Ȇ�6�U�_�&�Ln��F�̪�(��;y�ʬ�̭�
^���8����-��y��lٚ��Em�rGN��0���!�i%f��]�ZA��4Ixq��vl�@�ʴ@uw��x"d^;�X�*˸u<��e���4	0Ce]f4N%f^�ba�q�}�w��|��}��H)U�����l��w��)��j��o!�jA���4s*�,Ǝ�h^���2Q��+�Y�[y!�*G��;�N�`"��43[7�L�cu������A���#`�R������ϝP�6�9bε���٪R�M! N$�������N���b���9��/��*��H��,Z�V�en�WB��ڦTa��*��37�V�y�Sg.<Y��\����w&[W��mu���V�+V�,І*����������y���ڦ�Z�r�ٶ�㖖^!A��+�`v1;'VI���/^[�ѹW(e��v���Tmϱ$pVQʯ�[z��*�$�	��)���
�4M�laFimh�JN�j
�G�Dn�j��j&	v"��䡧m��T�Y1�U�����=��sr*Z�œ�
�YF����.�'	-�bP�_k��&�	)ͭ���&�]�}�U�wYX4���U���H��N�7K��ܢ3��xu�ʮ��v�.��Zɘ
NJ�y7��Qj����MB�JS��ĦI�#*U�%��Zk(�!0�YtK�{6�e:6���"v��F6"��平LR�(Z`ݥ��6�F�ӻf�AĥK�!�¬�n��铆�����Y[.�̄ǔ�UQ)*�P�*r��2�'��v�m�ff2�:Q��D��X�\�d���q��I�b�@�5�cU�o׳tE�OI��0�e������T�Y��Q��v3s�ɉ���un,����Q}1ͷ���fټ0R�TN[&��3B�{Z\��1FqLˇj�Å&e��OE驃lkhɘ킮�l�ٰ�mл�N���H��̋Rp+l�AX��lV]��h�k.3+M�I=x�䪤�4f�ݲ���*6N���}{K7�����f8v]���XE�M�u���uW�Fږ�,�����uS-�%�2��L�E}Z�:�[�O�9���n�tɕL5cjԋ[&L7Btd�� ����"�Ê��Q�Sp��yO���m��hdج��@�I�	��A�e
.�풢ӎ�Ѻ3�$�n����0fSԕ�GrՖX��Y��D5��T��,}Ĥ*���/�7O�E*7cI�˶�/sDqZ�7h41)F�m�r���&34�HSz_Ք����O�Y�U#�N�x�mmgQ�/�C!&���w�%���!m8�Q�5T4k�c+Me�{��;�����~w��ƶ��F�e$kRv��5�b�^U�Y{��+��KE��o1@ټ��UZÏ�9pa/kl��E�)rkM�"�[��/+���a�'3[���S�
�!1]O�4FY�R�&�G�L�y)�,�<76.�Y�����;iV�ݫ72eZ� ���7��X*Ў��j����,��0㧔�hF��BS�kN�j�b�y�S�ܭ(5��`U���)ݻ���P���5;k��VY���ξ��Ea���YALQޣR��������x[�2�A�d�[V5�f�͘1��e�+pۓ�����U����`;O`�/"�����{�����T���(�e��0��k��Z;ڰ.e�� (�Y��r	��4��L�����<�[��.��}ULڪZ��
G��pj4ҼK��a�y"Fm˷X����ӫ!^�ݼd�w[J��곘t*H��Y����_ԙ�kKT�o	ոe�����N1�Z��#L�m��lS;b��8�&&�R&R++XF Udݥ,�ONL������&f�ĬHBZ�e��8��SqU�Tbt�T����w��\��w�5Z�c��:��#Va��?3��6*<Co%��ǚ���Ӓ*��i/r�M�˼�i1Z�;ٰ�h�B����Qqc˴m�f^e)Z������nWe5E��H@ۦ�R��UL�;�j�2�!C�bRKK ��4�-4]��5�uk4X.��0��B�d7v����yH��R����7>\ͪ?b-+[7�b�g �������%e��R\˪7a���ɡ�[��k����,];H%�*�!*�EyL��r������9Y5ϊN����j�,E���'K1*�{G���Q�Ѱ�a�!�i2#��;v�q7����pРj�y`�2�G�m��ϤԬc��sX�{q��%�����5f�/뗚�� �v���&��Q�d�$U�Vr���1���5��sxO����J�����_��i F����|�o�HD�Q���ި���/c�}!7�|�g�x��W�+|�����q��9^l��QVq#�\��o�m��B���k�2�[��EZ9�F����v!�	hM"V��2�k4v(��J�Z�:���2�z-��b`CE��8���P�bU˒k(F	�;��Y��m�`dt��i��>ihwqb�����87n^��+J�ӂ�q���j��@s�X\�2�Tz��o�+&�o���2,�L�%en�*��æR���+j��oC�����4���B�[ܪ @jO+N�%����Y�m�}�_8GV+�����b����b���I�u�FA/�J���B����wk�Lj�rJ�fs�=��r�푯3f�L�,dUܴ�n����3a.�7v���f�TF�������B[�S�n��}sg�Ubt�h�yo��9�m�̈۵B���h�l��<Mv0q�1@N��l��tF�/3d�&��\���x���pX�f�!�<��#q��D�y�n�Pӽ˱��Q��*���=k�}N�>NF/gn��I�ݱ����͏�Əb5���5-�	]9�v�e^E>�6�X�{�i �k��;q�(u!���2�C�8�ƪRk�����3�v�PB����>E�vBwb��"0U�h������k.�Zy��V/h�GJ]��
a���}�X�^��%��j���C ��)R�|6K�v�-f�pH��w0�Q)���Z�k/5S<L�-��ș��8{Ku���w��S���)��f��4�or���S�d=�,�J��0T�gڮ�Z]?s�_:��'1̂�:2�Ğ�>��vB8�YkN�c�ʖ�J����5rcC x2b�Qa��dz�GN����u���Ic�|wP�5cepӴ-|�%׽5(u�5��iӺ�җUk��:�[RJ8�J�;�U2�±9.���Rn=���/a�<-�|&g)x�u(E�KO��G����'�󒌇KV�qx�����}C����7�wU�]�2�yU����9̻'�4+Mtx�k$^��Y�i����/c���2�>ϟqX������{��*�`w�6r{�
�����֜�閁ͺ���u]-6q�,BM{�*g�Z��u��2��EQaK�Y����,��4��xNol�������['��Az�|�?��K	�}�;&�,X�(qk��2�c�n�>}0�ޥj�7��ê��xܖ�u(t��Ȳ��Z��;+�If�`�+h�3<k��ܔ0�Ք��t�v�S9Q��v���T��pPax̬��0�a\Z˜[�4-]�yb��+s��75��"0/N	�F�ne5Y.���u���b���)B�)��ǐ��w7�t���a�%+Ni�;a��⥔�ZԲ�ݭ��1<�$ݍ����6U�o��J�Z�e��6���f^L�]ͧ���Û��
h��k�u{$(�;ǧX`�nK̵V�Z�L;Pӧ,\!]x��+)�U�+�USO+����0��V򡉉W�^T��E��9s7{&3pS��'w�tٺ��2
v�*Z�����}nC�_֦3��'wmp�YF^�]�F����d=q��D�oU㰚�:<�T�;�� ~"��O��m�V0!�J�\���F��6�Ȣ�=ƏD��Hdɽ���t>�H����n���������3p�u;"�U�������)�d�\z�S�{+�K)�z$Y�a���[������ǈ����%�
��J��Z�+,�R��G��	��LəMV��^{���0�"��4��S��[�P�]V�)2�׽������Wi[󬣡��yY�ɮT`�ρF��T\욡��OW|nc�Piɂ멳m�V��d�+r��Jf�v�h��O�#0�z�P�������k��jX���Y�B��pfe�&�[�w��]�����F0�S��e�sn��+pͦh��;T{3Y4r�$�l�%��@�rUӴ䧵݌��q0��eky�Ve�oPr�;���X�M�ڞ�_"Xg��L�X�����U���0�8[��ت9�&���.��fPPi�����÷im�w���a�=6���]�$���]�Z;Ŷ��*C;ziՄB3�+�;2����0C��p��n;4:�P����( I9�->
�8NZJ��Ӵ�3{��+�p��8N-�X%�r�Mй6��¨l��^���h�x�Ѳ�*�s�зLɫ��F���2�����+\:	=䢫��`�}{�Oۘ6���[{!��6�{e3Uf��@b�D&�G��n,�.ŹW����k�)�{2��[�eE��<��v'G�pJ���lx��й3M�徏N�9nٽą�w�s:�<i7A�xv�k�{}���Wa�\��O��:`-�q�@�R��dK��tfA����Z�¥&ͦp��d�:$�wB��/_B��+�~ս
C*��ݥ#��kn�*�չ{��A�W-L&�zf0vbE1���l��;E�!�#v�`wd��qq��� �+�5!�Ch@@�|��x�q��|���h[��@���:��HN�wD��ZV_@��"K�L����p+��٪�[d�B{�Lԓ횵|Zl��3*����j�r0�a��IW<�}4ݒ#[�m�����"��9��Z1i��QY�J��C�<n�[�	]Y6�Ot6ڮ;�3��+�A\�T �4����lK��<s��sT��yc�a���ygw��m��T�I|����ի-ӄ]X��e=�Z�G�;����bGA���k�;il�ɮ�/�#�����۪�d�ޢ/�3I�V����b�ufA5����Z3�'�#{M#g�Q��q�w���[��Ff!ƶ�4�c�g�sG*Z�����3f���i$��mm�k�kb�3S�M�����޼V�j40�"�R�iV#�x�f�I��))]���3�aQP2U+i��d�܉��2��ެ�`�yj�ʅ\k�e��eDz�^:6i٬=��{L^:�ޣ2�m�J]:�$��V�1��rJP�Y\�q`֤�v����[fF^����]F��	Y�@\���b���î���5P�� ���y/y���hj��N�a�}���6wW[)i�`S.��t���aa����wfU����.�@ͤ*v��I^2znK}tkK��o*J�.v�!bp�]M�	d��J��j�y�zz�5�֞�k���l���&:�,�M�ެhC����*9�������1�R�+N��	jU؎����Iq����ՑZ�1����F�<�	Q�b߅	MF��\�����D��s�]Ń�Vwr�õ�+�i-���Sn6��e-rmcY��MXz)��)\��d�b`����u��0��-��H�]N#�%J[�;؆megW�]���]*hX�6a t�oOHh%��� �/;;��8�r!,�W#��u�	xٳ���RSR�u�J���9I��<Ƭ�y+(΂D{�I���|�a���I�yp��J����9G�� i����mmmF�;'E�1=��-uF�vb����n�Iw���2��]�h��+&Q�^��X=��i��kF���kO�6N���7�x�W��N�ʄ<��lA�JB6=3@� J����z_f���=��53�!vQ}��f�4哄�1�%����:��g,����\ʼ��sb�)Ո��S���_[w�]΅�Uԧ2�u�%'d�9n8Wj�xc�F�6^ܐ��͖L9�6e��P��H���	 �ƛ{�9(�j9��y�fԕ�
�pc6�,.˔�����)7b��ճn6nУ����l��6�pJ�6!�i�Ҍ��vJ�2V���1qNA��#�L�6*%9s�E�+=�,ŲK6�TZf�%�J0�Is�N]���ND1Z�I�u��ָ��t���Í�k���ZÆ���V�N3wP��+�VRk����&��ܲ���f�ݧx�V�g�^ln���j�@n�Li�A�:�=w��֍`��pe684[9$�Ӕ(#v:dV���ܖ7J���ɐ&�� NI�_L���������K���C$b�]���#���I�+����Ove�͓�'�m�y���㳔�u�C�IC;���^�)8lqRI$�I$�N�X�b�y.n�Ԥ��U9��{%�ZR�I2�IG.��3x���DtUf[j	1�e�*�=��2�ŷ�V��o��������r|W/��|����T��Ż| �"*�G�C|�!�C�G
 ���?B=>��p��{�7Yw�k��x��V��ȑO&fV�2K�����c�o�k&��}X�ݣb�������f}.wm���ö���Q�̠mʕ�Ƣ��#J�ц����Vd�1�@��v�<���6+YX͜B͹�|xp�Vuj��=[+jX��4^GX~2��By%��K�<�)����n"E ��,���9\t9UY2h��ʢ��>b���r�&��5����$S,��@�F2��m�'d�jU�+����L���T�r�s���GX�Y}�3]V�y��u#�¢
LJ��i:����ڷ���y��&��Bԥ�p��l5�aZ�Wp\�;
e �v"Eq��ԙ��wos6��B���9�̠n<��GÔ0�4<��E{iJ���u5h�m�QCȘ�qɚ;	݂�:�Q�d��%\�^���=x�ix��u�Ҁb��k{'�֝[b�
����\�
[�䊴v v�<���"
��fcu�����^gq���u�lvR��Ѽ�s��
��=�	#7����Hrb���"��Y��*�m�̸�sou���s(�]�M\N��MC"���1�p�>����S�Y܎�B^�b�����V�Ȱ�{&v!u\�=�U;����6�պj�T�ౙ��ޥ�����O#�>E�b�^�6,?��N��m�UHJc/)�Nu��,�P�9*�v��Ts�3
0�jg)et������N�5kնE�q�^X�֤8�B�T"p�6�7����*�42��˽f��Uv��S8��cWe^^�j���"�5��W%�}Tn�ݝO;z`ѣ�GNk����'��R��vgQ`�GJ�G�:���D[�\�7LY]�ޖ#��*�ǝ���J̗ԫnV$��wt�R;rV��㬹�/�vdO	��9�D���V�6�Zu ��K*���)Na������5d�+��Ml`ЭŻt��2%ڂ6U�6����wN�0a���+y5}�|Fe)S0��n�H�-#Q��Gv%fm12�*�\�;�p�Tk��$�0�gV:��%��ї[^ujY���r�$�\9�u�w]��������:�	��V6�nn�T��F��B��,%���^֎sa^�ٝ�\}yo"�k&ե\ 8��7w��"Dp��$�Yn�mU>O4���v��Yï��e�*��Y��'�s���Tr�R�Y��p�T��`�`v4��JY�q�NstD_Z6���S
�R B#����
���H���²^�UCy'"+/+ay��i���S�)u�*a�a�_e+�bf��Oa���6$�n�=B�*[����p�2n<�W\��)l�܊���*�P"�4��r�ݬ�V�b�ɓ&
��z�w�Zv�v��2�u�`Sn�=��5���#;
�+��[���qT�-S�n�T-�-�/`垲Fe18�J[�3���Ù��Y�$z��uش����0�p�?)A�1t ��/�:������5م�M��s413�GDN�����f��3,�xGa�LX\�0��!u6��M��s���d�%��ʌ��
�[�[�R^I�.���Wc���i�몡9��Xr�8�S{�������iH^�Ѽ��l�N�x*V�֘�ki��/�JY-����q���������f�޺J��dj�"`Ⱦ�ʶ;4��3�踓����p�1���$�LQՑ*�Jf�wyILśHmݻʱ�ѥ�W[eT�k�s�B��ᕗ��ȻN8�϶����U&9^ò�ZT��͉�od���/���,�z�ƒh��^U!�S;����]��9�yoX�j<{��v��[����t��U�\�Yv5ڷ��J�+dSi�.Z��{z�qNf���>��
��,�X�|�㔸WV>,4o)7/��K+�m춵���w�I ·��7"����Kf̸�٬�i����\��I:��x���t��u�M�q�ع\;�J90�������b��|�u��pj��l�5�: I�����nl��d��+�e	�+�7�_�^1f��0$Q�)f,��i҉�B����X~
9:f�A�\+C�z�`-q/S�s)�)��خ�X�u�"T���]�wF=���g"(\��ɹ\mҮn��OZ�aŤPݦ�2�E#}fVwU�vT˘�p�N�lnP,�QF(9p�̍�����%(,v��_m��o{-�N�o�.IYd/�����L	�g��y�7���u�:�EwHr��ٕ�j#W���1cs�J٬G�~X�J�A+B��K�ټa]��V���S�>'-���ڳ]C8R�y�E�d5�KF�a�7��H
u���vɭ�ʵՁ�CCb�IQ9z#�\��Q]f��k���n����Z�joE*җ�f.5:�ϋ#Cl,�3���JuvM3�]���4�^,�Y�"	�F���3H���̤��ڼLr�j���X�m�07kk:�X��������gY��qFo_\�]v��1X�hT�k�[۬���t�.�@zL�DuF"4(�a�8�mD��tN&�i�%���DE,��Z$���>�V	+0a,U�"��Ǔe 1�GP47���륓�:��m�ƶpi��_Ӯ�R����WL���MIٖ	-E�U�{�U�_.�cj�v^�'\,���[a�f���Qt�
1^�s%]�n[R�m�i�A^�
TK�K�VF��źӲegm�E�����嚻��n�o5��{tHʂ�%.�h9� j�PNu�}y��/)Q$��As�݊8j��h��m��#��r����YQ�t��e�A]v/s�$���>����gMK�ƣ�\��d�[q;�UȧTP���F5���%vP��&�Jn�RJ�L���+�l=�M֋؛��ْ�;A�r#�o:=�n˜�&�n�i��gtY�د�
�;�0\<�E�!�9�i��.9(k�(1O�Ĳ�AQ���tl2�Zμ+E�nP\��C���;�1�̻�_ӌZ�M�q�y��l{���U�0�S�����ҡ��ǫ5b9DѤ��Z�UG�֗E^i��"���I4Z����8E�zugdO\��jvhat��"6���ͭ���!��B*�v�>tn�VT� ٨^I�����c+��Y����q	]�f�2�X�����9>�Rn������r��|�L̶��\����mf�R�5�(�Y�9���꒹ۡ��*�[�����ٖU��X�|��T�E;��>[2�^C�����w��E��'AF�eWSssr����[��'p�����nB�Hj�䫴i�ou�\[�6��}���&e�mGwv�#8��Gj뀹����Zy���JI�+�ɝx�[}�p��o&�'R���e�ΈsL�b��,��y�����ـYǉجV�:��x������	Z��}��y;Y2��wCJ}]X�g!�F�y��浦���%i�gK��w0�/�����3��|�[7�U�R�A϶螑�އV���RԂ�wH��9����=
]f��"�����f‒p�I�۽�VU�bM���j���������PaV�R��3!�gk�S����YVn����z�u+���>!�'wj�8w2���Y��F�*���t�s�&�(�3k�;gd=�cF�t���Tśr����nK�����\\mv���WEv$͌�R��PA�V�w����>�zI*m=�6���]:�3�T��i��FX�R�T��*�tN��F���c:6����n����&�4��������t^)�w���#��Uy�+��]��w(�(抗������Cn�b�,��Դ=(�C���F��봮#.bvUX�E��)��($�"3�p��[f����HS�7J���R���%�n��0���ʬ0LB�+FU�hg�b�ܡI�ƫ!.�cl�#����'�Lz� #i��s��YK�1蠞C�c;���3��X	�5�|�`��-��aK`���jW%V!k�p��	���Rk����E��q�=�2� ��Mڑ�Q��{�j��.<�y�yNM=��W��0�K�q���(�jgܯ"v!!���t0�kA�QN�	w1��e�`َ�4P�X	1%e�=�1��l�kސؾ��i�c�"�*�\30�b�S�[�����5����:]����O�Y�Vmi	�~b���� (!$��2�B$�İ���Xh�HX�=�[X�s�[W�x�z���[%�ܨ�g3<��e�om�P�/�+0�|�=A�5�vB#Bւ�S�`�]j�22����.��r]��s��;�F=4?3�zxf/l�V,Hگp�#���O9=};l��L�^�h��� =z��IX��.oMB�sLy�]u��m�C�+��<޼5ݗ&�.�����)��}��Qw"��7Q�i�/��A2͚�\�KI����](f�D��h��8z��q�O���e=@�G��V[�7�S����i���CG2��E�'6��̛uq���6L�#:��feT���=��ʡ*Iaǉ�t+)��"��iK��O�����g| P�g��Nl�����ki�8ĭ]��!˕/�$ �Hr�0G�7���ͬؓ;R��[�.*V��)���q�u����+;�oᄵ�o��HIH�>�^g�)ZD�#$M�r�1Y�Ƴ����Z�md��L���iy�2��V�"��X�
�ϩ@e_R+S�`~�����i-aC#z��-�L��PP���k̿l���S-E�J�M��͟gf6�䡽���>��E/��I��Le�Q�l#fs3gy]V����(��٬��k^|��ێ�ϙ�.��8άi�ŬmJ��k;o��es#^ak�$��#X�>Y�T�m!i���PK�6g�u��@��+t�+$��}`���/��?i��*�xd��;BF�� O��َA�,&�q��n8�r`��Xw��w�*��T�D�)6����<��XM�~�g�^��f:u���]D"Grn��qF�X�4c,��MW�Eh���gBq�pԮ�ie��pmON��ث�ﵔ���}��D/|�=4`�3}&�q!VF�n�GC����եLu��*�
���p�+fV�"5vA{�KMluv$�qq�e�z��q��2-8�&���޹5h�V5e��r�5��]�R㓸�f+Q�c9o�rW���0�s���ƥ=�$_�YfE���u5tSR�;�\��;�B�{�3غ�s��Y�g1�Օ����wa<2>����xYA����'`�%�T{9#�l�ky���=r-���?>����ӭ"57Ǵ8�+Q���:���9,�q1}aζj���3}��&�_�u���}� �N�m�����fO��丑�*���3>�V��n�w�>��9<�����ݷ쮂�8#��8�f�eZ�����l#�~��V��ȧE	��!"n��ND]�|��η�pSA���[�}35�'�BWYx;��ƛ5�6�f�j���s����`�]��]�߷���˪q�3F3�y��ظf_�S޳C�^���R3[�7vL7Z��lg��)��,Ex�d�{CBɺ	��@s+�r�g-��9l���GM�<���4w:ђ�Ž\"\��Z�R�F�qR6���s���ʜ�&k������[���*q��zY}�
M�ؑ!�g�x�����@k�k��WT��N��P�l����bq�;�6�$d���ɆrO>��� c�
�ŝ�.�J9|�Le�z�&��zR^�78��;l��yл�3_+fx�X�F����(�N2�Uu��ng �f)[2$wBo24�:�3oi�m�!��z4b��w��FE�v%�勇3�̪�g��w:�|]�;Ͷ�_i�7U$�-�QyĜ�ٹƲ��[4VJޘ�8:Ҧ��q�qޮ+��u���#��(��v�}"׼�!/.e�0GqY�6����IN0�ɘ��esT�*�׳@�����z�^��9�"��N	� Y�@�d5&�l
����&��A$]�o=N�pC��'(�]`g����.�<u&�B#�Q�9[k��W�՚V�1Eq��ʛ9r^�`���g����tqMkv.����;X����u���i�XpAcv^���z�R#��I��݂�W�x�1۞6͝]�����]�|��yX7|����p"b�pUg�즛�d�̰,9��6�Ô�i��vD�D�fzdr��%��g9*"�WFyjۜ8�U([v��欿J*p�o�s���T�֌r.�GB�s�����;\ν�FQ����H(�.:�z�T_!�������֚��={�Y^�Q.YO�K!���t6�)P�ZnV���6��t
�q:�`ay�j�
s_pO�Z��J�����C9��+$�|�g{�9�j=&y�<:�;���6w4��I�%�仌���u����(hzom>��<�h�.����s��C��x�Lg-�.4T�Q�-�ȋ��/!cU�u�x�ED���*c)�w���;ج�p�nݘ��}�m��F��,��ՅL{�ۓ/ۓ����+��*���.��B���Yڲ��%d��YFr��KxLݺs�T)y��>ӈt��"K��^ɔ�=���0�+ȣ�������r���N8\ڗZ��J��זI����g��.��3뇜��_��#:��f�E�aŨ����}���Pa��W}��bF�u�jT��{�CL(Ɏ�L���k���QH�]l����U�unJ���8����E�c�v2q ��E�<���6�^��[�jo�a˥I�h�wۇ��m�k�V���B
�2qXq���F9������/�r�o+z�[S��No��a�z�Z�o��men���ݿ`�W�b��D��eV��Vbh�2���0b����S�&f���"qa�{�F�eG �_XR̰�i\}:���Ά�6�'4&LRܘ������辿-{Z����:�Iŗ����Μ��:�i	�]e��aaK���G?3b�=]}�Pa��`�92�t����ٙ��_���Z}����a�?���X%l�����9{R�S~�A����>�\f[�.�ǝB����;	��׀g���l<�u_�h��)m�6wKJ�Gm�����>􌛇>�A�$���q�Zx8
mA�>8��U�ܚFw��A��X5&�C�DΤA�<����ܞ2:���m`=ź�5tAՋ�*��{]��D��\�����,�82[qC�Y��-�&*��J�Yc�kr�ʝ,��N�ZC��h�#��x����W) ���ö�G�X�nz�9ڀP�z��S=�zෙ��к�Rq��a5w�}i�l�ь]ķ�%�n�3�zξNSʥ�4��
a��tU�L� ����S�{�!OP�h9��0ֱ�;�H}�je@)1EMZ��y[m���T��zi�)צ��#30�X&d�{�+2p��Ogz����[ �F�]����3�he��-n���kT�Њ�̖u�����!W�bM������D�!^���j���d=�>��l��F�8���WQ��0��Y�v�-G3"�+��2��.d�A�Mm��+S�mN���HCr>�މ��ST��ǌ���y���$�f+��eR�|i����Vd�u'g����%�9�
���s7<�CH��oeml�Y�᱁Ns�M��!�	��Y�����۪�V�Y��CW7��u9 ���Z*z2r7%�dX鶞曈���ۂg14˜�А�b��:.��b�����5W��t����i�u,�!�D��ul�ᯜ�2��G�`�.Y�q8'U�W�Z�OF�~}v@'t��*#V��|�g�:#^)�vY�p���2��t�!��r�U�/5Q�DN��2�\P��m�؋N�o˃�Gkb�m��q�Z^H�h��n�%w���tR�B2���V�N^�北���W3Pc�ҕ
���i:�=�5Z�h����;�!ý���WmۂyN�O��ؔ�kʮ2�&�"�0�o7a{Z�&��˗hi�:�/,ls�V0�:�[ha̗ok7��cW�H��q��t�k*�7��;�#��ơl��*���V����w��DT�E���q���E���Jsq�$���yq�Q����&1M�ń�X�3X��:'K��t�kwm���P�D�ȅw���s�n��EضS��;j�ˣ�֒��^wVq��B�s~i�s�ʭ5b�:i���r��,�v��T37}ư9�4��wΖ�6�3FNdK3PET�oJ8�b]��L���ɽ�\�Ky���'K���iG8Gt[qP#kkv�f�滯�4���wT����ڽNf!�ٻ�}q{����$���|�z��B+�
]G���ʴZ��;�.��M�c��lf*�mN2d!n�Ƃ<{��ī� ��w9��čb�F��ڽw�;/A�J9�� n^pyE�d+��g37����vP����n�k�`n����V�nSr KIHf���˖�������(��M�d:��B7����K���3�k�i��4���p�嗔�9Sq�ݢ[��j�j��*].��Zt�D]=�!�w�GV)d-g��r�3'-�we�DGk��8��yi�R�vv�o%>��5�0(�xDf�2��-�"�ؐ8z5b�_G�O�to�
��u�g�]����E��U���}N ��|��:��� ����!j�xC�[���r�I+��$���k�wV��BE8@��ԡ�8. ��Ԍ�TaVܗJĪ�yWj<��1VښE�5W�l�6�#˞
���i�����j�.Y�6 �E:�֡ڴIgu�s`�g�і;,�+�i��"��͠�ݓ6��n��ů��ь�����"�Va�u:����Ϙ�=��ٱǊ�X��C�M'd��L���U���݋ZT��7�iȪ��s_B3m�k�lS�k!-� �UG)u��ܴ������dHd�Ӹo��*�se�˙Z+�m���UcNe&<���t.�grʌ�+����C(�笗�pM�x�L�%�f��@���������f\|�n�eJ�᭧��P�3��<_'�~?�~sZ�H_�0�l�Ŵ�.}P�����kɉ)|��\�v�gm��l��jFL;�=���(����dγ���l�/�g.;ϼ���&cP��*�HN�B��M��ME����t;z|���X�NѮHU]%ID՘4�دh�DF�#*1M�rl�]OW���i/J2O���Ⱦ���C#t&d���!E��,/��gB�(�e^�UUEV�j3��(bV��&F��J�1*yER� �H/hɴoM��"�y�g˵	����	d̑�kY#j��ka7{^�c��+��[����r�:1{1�S�����$];8@���E8�t.8��w�ϫS�|��u�ד�F�C�����wE�)��v�>��������9|�`��H����ϥ��;{�V|��r�E��)��[���ֶ��щ�3�"CS��RV0	s���s�3��co�
\Y�އ=�V�t&:�X���]��<�ܭM�a7QYu�ЄN�����y�Y �<��*��]�Ȕ�4����wU�2y�E���Y*����s#q�N�����X��p!�R�Kv甼�Hv�5�����[��[�+�Gg:f��)�:�
�=��DAOh?W�wO���wC��˫��������a4��P�7cS"3��yQ���K�,���l�0w%:[��p��\'��a?�^N�_
���挈N63HaqsEF���m���6�����z������ɪ�/Xh��}�.�O�:��:���g#]2n9��D�������9Mp�*��\�����91����[����$E�R���|ӳ��n4N��Л3h�u�\1��l]�y�]��Ƀ*��z���Z8�]bu��
�9�R�*���Y��������q7*)���QX�����W����X��V�r��(�5h�P�Q���^,`�(���5���l�Y ���1}�Kr��U���º�S*g�J��)�6��8l��/f��a�rZ�d{�D�?+��\*��wXT�4K�5�7��۸jm��/��̻�n'*ԁr��z�
�~9w'��]^Y����Y��� 8�.�����T77��Q"���2Z�:��Z�Y���#�ۗQ�sշ�X��\1���sViI�Z^c��ר�E�@���&\u0��
��a�!�l::�x�y�W* �6���l��s7�j�g�k�N��3���
��;(joE( w^JT ��I�'�'!�mu�����[��p��˃��a �4��dћc.Vf���T����[�ȍ"������W�z��3���	��`�g��j��5��J�\s2e(S���%<<�so���1�/�@=:-;P���h%����f��C�5�Po��Z⋘ø�#�;�J�@���7��.�"[��a����к1�yg5�Y�B�]����
Ŋ;;2M+5�fXMp9���W�%����R�b'E��Lc�����	P��<KJ���ߜs�C��B�s|]�I�:+�]̓�0�z��>��d���y�<�R�ލ�E�o����q�.z��P�D�m�y��شc���������7��<�#���j�q]G�M�mF�COE76b��@��pj���*w��b��#Ｇ}��_�W��C�~6m�.U'���u�҈ck/Gr�
�n�E]�K���;���}�8x�dśԹ[�G^��]��y80w0�N���ȏMV��}_Q7|o=�K��S�t;��.v��B�B��|Л��%E7���o��G��V��;p_l�Og\ޭʾ}�rt�\��i�ͅ�B��y*+x!�B�����T�h;�\��y���P{\���{0�}��:�=<bx�����9F���Qw�ͯeKf�@u�LB�U f!~������}�w��sm���k�PmQ�{T!��Qɨ/"n!�-⽘����ʤq�Pb5 -�G�F⻁�_9���+�=�zxS��(1Ш��;��1Jr�zf(j!٘�� r-�P&a�R:�`�Y�MsW�l�^���k�<�`b!���N��^L��]�o�E�_f�:�KC0]������uŹ�I;}��I�c����>��SQ�
�r'���B�P���v&��oA辘�`�A}��;����D�jC�J��n����^��.a���(f���Tۥ�����;�,P'�f����o�S�����jq�*�o��_Z���阎 ���"�.`v+��,)�n%E�*-A{p��"��Q��$�R����n��g�����7B�����/�B�OF�N@�[�JZ�P�/f�T]D3T��Ⱦ��*~��[���vg��߲��۠ē��[7������V��!��g��DA�����Y�v�ó����=j:�Fy��NC|��!�|f�s�OIH��_UUU�����[��sJI���@�ct���57@�S�� ��6����-@r�E���oY�o��>�����QK��CPE5z�V�Q7$�)�pK����M���@K�׶�J��_x��_�SP]�n��B�P%��s���/A؎�z!x�)�!ؖuCȭB٣��-�{
��h��I7�v�Ϸ�Eݩ]E�Y-�G��!s��V��G�q�R�M�Ņ�Ŀ�Sɪ�M�צ-~�Y׻�r�b.aQN@�ME� �]�����,��=H�z!z��о�M�o���K��s9�٬�~�y�_����Zx;G"�#s��b�b+x.�B��P�T ��U;����!{���W/�o���P9�1M@}�PyP�m2j����G�p_E�AN�b��C�dGq��LF����}U��u��z��A9��1������M��*9����+���z^#�R���st���YRn�Ǧ���w�N��QG��m�Tf����Rn/�Q��OE�LE9�;�}��CP[n����w���߻�ȕځ�RE�^��5q�G"�!{R��{Rv.���)ؾ���4� 7������[�+u�[}Ϊ�Z�/+Mh��m�N;�'ݕ�Ng�e��#�N�<��)τ񽋓O3�,Z��4��l������Qr�~̄%����o�� ���s������~Gh1lz�EqZ�/�y���r�D$W0w=��o $���@��9�g���jϵ�{���7;5��5��G1�[j�3T�@l������n/����Z����3��m9|U�3���λ�W���AL���Am�7-�]C�L@
�F�9�ޕ0n�E�*-�@n'b���i�_]ק�^C�i3T!x�"�1Ob���QS$=�C~�-w�p�qBڽ��V�n��s��s�p���\D=T�b�Z�#腱I�/�r	&`9�z�@v+�7@��� �\쾫կLw����wg�3v���G�d\K�;jA}�L6���p9�X�Aj5��T�;�U~�����:� �^/�z��%�b�Q__V���K�B��7��==�=�+�@ױ��/�w>����-�r��Kz��^¢]�v'��|�bߘ��(��,I��硏R�Z������}�kym]ޯ]ϳ���m��1��y -�w�K��{�pE{��b+ȸ�,����f!"'�lg��ߕ�[Y�w�ַ:%D|f�B�B��3PM�&hC�-�P�sA�j)�t�b�fx.5�*^%Ay_x�=r��k��.��G�Nk��뺲5G'6Gf�<ݐ����\w���Bnv����e�[g�(�Ʊ+�Ԓd�]�1���:5Z�6��)W���Cq�\~#x��x.�P�T�Z�QMſ(���]�#���}��^\�=�ȍ�F྘��
vg~�U�^��=�c\����5@Z��3��@��iAm}X=/�Sq{
�":�ؚ����z/�H�F;�_|�k�.� �_n��^K���30��Aj!��@�����'"!h��غ��4!؜�3�Mw��7�vx��W�=�C��A}5�J7k�$��T ǨM��B�\���B���&��5�7=lZ��3��y��]R�u7E9�7=��1��y\��\���eKj�E7A7�	�Mǘ�9��{Z�u�rt9�U&"�)|PvɈsB��&b;��� ��#�r-��ȁZ����Ѹ 7��p��ڽ�|g~8."�E}1�(= =D�_b��C5�C�9������;�1 *���s7�sڴ�;�kfx�@|j�D$�=q}ځ;^����� >�g4�ɨ�-B���y ��u�}~��/��]�:`b ^({�����Ƣ�ԏ��Z^� �qA衸$��Z;��&�@v�}XŦo�{���`&��b>��"�t�����
��:1�OY����>���Z=&���Γ#N�F�Fr;�g���׻έ9|W~eVj��>ux�IS�k9�R�j��K[�â���U��;jKz\1��j�����R������P���ֲ�M��\ɫ�{OT9�(�ך�*��I�L�~>r�
��&��ϸ5�srt`��h�)çf��W��}xT�`�^ޡј�W7�t�{�;�A,;)a��%l��R9��ʭ�'�m�Y��4c�^8��f.d�7aH����s�i�������9ed�r�$�dܫ�'��W�B׍l�D}c�o[��%����T��6Q�a�{|���ځ}b��3׶r�8XȢ/K{ӀGeB��g�g�G��TYy�G<�����KDml�l�R�LP.�v��/^����5
�F)�q����
������fD8y��J��ZS��j+s�Ͱr3��@��h������j�Jo�%��I��U��%�j���;x
S�rШ���5�'�ۜ�R�ڴK?;>D|�~�&�T.e�7�ہ2h]|��pP�j9:��&8���Ef��P>9��cn\��G+�ӭSg�d��@��
���n�w�	ٙ�8E�@�Y��tveSM�g�I���b)��fz79Y��Ѯ�h,0���9h1�vCsl�����;غZNY6s�F:ӻk�y�x�.vKUFm�g����y�1[���I�����C�~���R������em~���ͮ�!�Oe���m[���ٖŽ��V�6HŃ���/�g}D����'����l��ٝ{�~iL��0�ۼ,�Wgf[\EK���2�gX��)����Fެ�+��i��h�b��X� �k�f��o	�F]U��(�~�z��O^�h��Z1[ݒq��S�3��@�A��Œ�d��E��Y�������M�h�@�R5YCq=4�u��ŋ.�n��9�������v�L�92l�f<T��u]JO6k]�р����<��N���tj�ԏ-S�;c��.��}�Mc�kNb��VRw
N�j�
�s!�B3�G�1�����e�ꦹ�J� �Y�9O�e�;���e�^]rK����hnjv�4̹�E������eՂ�Da��t�U!Dj�ulfa{ԣ��լ�	b�Y9�_4ͅQ���ٌӾ�j��aL@���ry�>�O`�+�[�Ћ5*�+l���9.�EC�����[��О6q��/O��&�f:!A�l��WJ'�N�h�x�+�l���+���-	�ޑsQȦ!2��M�\�/��]E�r�pU2f#7{t쫋*B�{�0C���  ���k��j�6�6Fĝk'�P6�tgw
.4~�=�'3BŹ���d��D�r
W�V�a�`����S�Ww�6:ڍ��;V���u̝т[�$�t*R�DH��!�z����vT����k���yKK|�ϸ������n�ؼ�v��q�Wy(��H���yqu̓�.�-�����PA%f�KIJ�=b�4].��&=Vw�������w�^�d���In��nc̗hP+i�T��f᳽'�AJs5�@E�Y�|�J�$\q��r��*KH�Vz����n=6�Y`j|(�q�0�B)bc�I�q~}��ܣ�~���5kFLKZ��dGy2gV�VG�Y&I2g.	s.��G;y�&m�CS0�z�X���(��l��~4�� �&���}W��"��6HZ�h_/�e
���R|��v6e$f�Yk�2
+�֢����i�J�c�[�Ť}f�*l�[6Z��5L�i�ڌ�vj\�e�ٕmE�7�u�7C�b�f+i9��R6D��#��U&>�B��2���H��Z���	��Mz�m�ѕUOI	.�:W>͓M�ժ8�z.�M\����c{zql��E�]��g)�h����1�;*6����IW��߉�����~o��\��4w�'��vN�<�V̆�JP���Xw@U�������40��^ӫ���q�-{�A��� �����ˬ�������~�
s]2yޕ�+�y������q��0��9a�����[7t�N"�Fz;�� ^��9Q��֞din��s�B3q���s���F/T�xtVN��=�L��p�Og�ܝzȄ5�~ڮ��"sσ�T,�}.y��f������[=1��mb�X&����w��W�PKe�f�jm���&
��)㞣��-�T&�Z�2��d��aSb��<�'�������!3A�3/;=��MH��՝>|���J�����gK�摙:���(��c�K�r���u��~���S�ʏMwj�t�mi4�|�/C��]��G�����d�Q^��	G����*��	���	d}r69��U�V�����e�|Q	����seP(��d
btgE��� Xuǘ1�PE*^�z�����DF�s
K�^&�U~�W�5[�;��o]�̉�^z�0�:�{;�E��{�*��Xv���
R1��OU����/4��qܮrf��ENn3��ݞsRQb��<�ن����8_���o\ӊ�0��b��uVm7��1�8_�]�4g$ˣ�WW:w�t��e'�/tRY�<C<k�#fwߥ��n��#2g+���}�d���a�jV�[�WСES)�D���ߴm���К��]�����峔��6�a�;����w�٬��&�2��V�)Ǻ����Dzn*~�P��	���VF�\���3��b�#ޒ�xܯ\qBM96���@��=�R_Mn�Hlݨ:����[�E�������C��թ׀3n:�!�Ⱥ�8�����%� �ƈ�U�^.�gj7�N���s���'�C�0���*��#��L�pF���F[u��ð/m-����:FV�.w�}�F+f&eĆ���ơy��<����9x�ns���9���q��d=W�ߧ�#7���Mh��5\5��r!΢���"T�TFh;g��2��rWi�&j�,;�:7aCDhY�;f��C��zn�:��%�2��PX�lu�"����qMz#�`�K�z=��!`pM�G���*������T,��:���v�I�#-Ŏ���k�6�*�ʽ�Y�͇D�..�#h;m3xk��.�N�v[l�&]Jj�I�G�9�F�"�6n����`���ʹ��Zy�]�5�0u��	�g@N{]r�ӵ*�2*E�7��.r͔�<۬��-�.��q"�	S(m�;t�sL���Ήf�R��L��#�H�
n:���ǂd:��j� �3��[I4����
�PuV�	�X��M>3d�]�W^�3u
C��8WLuµ������Q�X9_Qt�9�j*��9-�;ch���<�O��.��~��m������}��	�cK �_�;ڿ�{X���w;�V������b�q�b`P����M�
ܐ��{���g:��$�1��5z����6q��Q�v���)J��Qtp�`~5z�J�IX��卬!�$�I�w��X��gb^\�Z���[Ţ|tҔ>K¥��]3��(Lm`�bt������`�`5ډ-p*p��e��ʏ�9BOe�2V��{�=�g��]i���^�c b��WN�c�#�~�Zw�=�Q���w�6������Ya�Oֳd�N�V�j�ĝ(lCX�K�6Ҭ3�]���8s�w�2�kӰq;pN`��Io��	�QZf@�0�'�}U_}S���9o��[##R�zx�i��o��]b�o��g���[R���U��SI���.��J��3f6�5�4��s��Ε���zZ���s�^w��vw�J�6V�{�\�Y׋�1}
���JU��OE��Q��eMF��T�8�/���Є�LS5����w����S�qLF"=�8�\nE���˳�g���'�[lqf�Q��ÔJٽ�S�_��U���W���=?z��������9�\�^�˞�+��V�뮰F��)-�@�����)X��Y��F�yoڰjݛG}8�:	R���e6&a�/�!k����_B�g۞ZWN��	G�z"=]�����*6bU��ek i�k`��i���>��z��wT�ʽ����fF���\��-��i�[`�P.�ә��:پ-�݅�Tx^l�"�6"�p��t7/�W-���0�Ҷ�3.�!������{ֹ	{nM��{��g������U��+C�����#h�n�i/P	�wps[ޭ��1��_�c%��QQ�{���hy��aGl�0�QlCG3��Df��ؠE�,� B�{�n�z\[�*�ܷK`)+8lέ�Y��������3������e��X����G�w�re[bY������$C�Jkd*��<�$��(�1'�U}��Oo&�'G5*C#��0߾<��7��T�@�^6ND(=��3{Z��V�ڃwq��wXN�e��q�1Hn-�T�z��7X���A����"A)����w"���Y�{B\�|"�8��O1�]lrʵKF�2�'-f;�N1���u�nT��17&m��ry�!��ʞz���}��T�kl�I���cc�H.����Ҟ���MG�e�ֻ�`�2w�=�
N̗�2�%�;��YL�<�s���J�&ۓ4x×~Uwa��~��̓t��ƈ2�c��]�����%��eM��լvLŏ�����zXU�ƮT��$���.�H����G��u_b�Z�x�`K��;p_$�	M�����@k�罌Z%�uiY�YV{0��M��]uV�C�md��o�֍b�^�9*:��L]�Qff�La ��"���4���n����F���˿b�����-�����Ec݀��c#�qȽ�vy�/\	�n7��Y�5�x��ֽ~%)�h4�>�W�B�Y�>�L�=�5�zPqn'ߕo�I�|��v�Tխ�a�ʺ�����Tɾx�z�u<U�{��;2P�}br�,ֵE^e�G�/v��CEY�f)�W=�q�i'9��]y'=���(ļ��s�M�b	]܂��ޏ{���֛��1?{rE�����
m�r4�;B�i�m)Ĉ�.�ŗW^r��&�1�q|�G�^�1�{���Nr��딫[\��ӄ����?}�!��Z6ɽ�ْ%��n��}*����ٹ|s���(�Ro1"�{�L.9�)�S)��5��<��F��q#*�`��[�ڸ��\KUF����C{�wa^��v��#�c�OmDhX��v��mWL�G�B�j���U���j����{b�G9ȍH��*�F����d_����3�����FB(4]J����j�:�=7�ا�HHo��+�ܰ�T�q$�:�b������v��A{XF��WT1�ɫ�wgZ+EvD���M��n�t�����EZF�ްY�ޝ����򎻣 ��w�6"z鹔.��%��אk��w&F:��\0�Om�xӺU��Ӄ���[��h�W�h\6;j�M���m�*��a�=��Y��2�7�!�;V��&��4�����k.UA:�9׻v͔yl!��x�����>3�y���l�ot�*�DҪ��\�>AZ�g����(8�5\����V�e�u+pH*���>�w�h��&�iJ
�I��';jη݁���)^i�E�\{^s"�L��z��;�K����fv�{��e����b�ɁB5��/6�bA�
�F�
J	�:�;(��y�����3L��)Y���U�?�Y/4K3I��O�:�&x��;��U��}2�5�F�����&�h��"-C�ޣ&X( ��"�I��V�z���Ѭ�)۹#���U�p�i�Si]��9w����#��b��v���˺Ka�Mf����U�`����d��&���@��sj4�nn(ޓ�f#��q�řyl�s�y����H��$�ӥd֣r
E�x+�ݫ��O�B���x��Jvw������,�w���Ƃu]l՝3�bL����x49O��خv�]A�X���ꖨN[�oi2�hcQ�/w��)�Gd3{��&@��uԚִ���1�U�E��U�|p5�YՂkk+�{;��ܽ ܍'+'�����vd7X��5�bWJ̝��q�̽�)8y���G�\�ڼ� ��)]Y��L�	w�B�f�>bq��QDqn�i'�������.��1$��Lh�����sN�Mom�R�)b�&צ��Z�]^s�ѽ
,^��p���M��Q/^*՚6`�އ�C�F�M��ި�j}�қg�>�
{{�b��ٲ2E^��v�(�PCL
1{�n�LS3����)%/"��e�)'�����$�TB��E
��_TZb&�{٥&H��A@Nv�RF���Jn�L�:m�B����ĵ�mK�TY�:-d��u��!S�np�v:��lO����a�'�u-�E%���)��<T���u,�)�H��IO�N�_��u�UoAFپ�AgM�}�cq(�.���5��9�gZPJ#�K����腸5��t��kH�WI->�V���椒8�5�0s����5t;�"n[�2{�)�\+���T��يBޭ�3q(��h��m��Fը�j�S�X_n��o?�X� ����<�'�F(dB�HP����'5%�3�q�s�*�[c#�����5�x<zm�-� lƊЭ���tG"_��}_}e]�Y����F��1�Cv�P;�~-9�.`�n1���9�f��qG�EOm��k�j;����jN�����e#g.M-�����ظeYI��4�8�屧�o;�O�D�k+]��Z�p�Ȼ���z�eGv\�Sx���[�)ɮ�gwle����'��%/�z=�J��i��]_P�Eۀ�1�C-]��<����1}9e��+@�3J:�caY�y`�395�ud6�OA�Fc����:&�!��V!T7�d�
�����Q�͘:�� ���_��쥙G(�u=�	�ݜ���D����۽C-t�`UIԚ��q:�9xd'���E]�"�{/V��~ޢ�4��{�PS��s�E���#.0bB;9�p�k1�
kc��@�{Z����O7��W�NF����شt^L:�%Ȼ�;R���n��01M<�ۛOujTA��G3�P[��ʓmg 'J�ȩ&rv��.�'T�v�5sE�Z�FҜؓ����ރ�{�q�V�,,����7k���ɺ�}X��s6˨w�yȨNı�=�},��{�z�yqf�+�o�}�!
����FON��u{���G'x�u
LS�YsE\~j?[���p3�s���u�dMv�A�f0OQ�c+�R����ֻ�����2�TpW�x.�BkgD��l���{�l�#*m��hH��v�Vx�~�E�����*���󉻄m�u��Ǩ��|֠]�d�k�ӕ��Y�!��c��Ǿ�4�e���Kmk C6<԰�'+�˼�Ixi����'T�,�eVm��(�u	���w�1�������*�ga*֨�]�I~�{��D�iG�Y�An>vT�{M{��~f~��I�O���W���3�Rd�$�>�4��K�'<&+H/����䵇��±��{���:r�r���g|�W��:�ZQ%;c������h�sq�v9r���L���� �]Q`��DĢ�Q��w��]�\��V��U�&��*�eu葲Uy�w��}�r����|���h�G���f����B�Q�w�O�������ա�&T�Vr���b���;���x�q��Ӌo�+}�8cùr��8�HCdm��jg_g6M\kn2$5���}��üa�a��B���v�wښ��2\��x���X��
�#�E/���"Owqm�}θ�$Au�k1���Uu��S-ވ�[�P��;Uc��ƥ�y��&_��s0�k�F�W�$e��z4&�������l�)@(��SXWb�[�{�b����������CΫ���N1[���y���֡���"oiA�Xs�5bKprN�!oU���-܇t�	A��d!fB��Dҁ�(���皥cE��^�i�O_F*�g�Tq�:ګ%��w�ko���"��rr*w[:���5���H��9n�]�#��~�Y���e�*C��w�(����W!�'�(��b���Z�����ǋ0�ξޕ�1�(��6�,!�"�����UU}U7��n3 ��,t��r4�[�[p1�u�������P!A:R�b˵GF�Y�f���*q/8�&w�3�rW߰O#,º+^l�)�k�rw�>!���ԨV���%x]72,�k��$M�TM�����.K��f�뚒s�m,��s(_!���h�(�혺ǁVCKd�G�c���j�K�[�8��d�^���ف0�f6U���,�u��+��=.�!S�˸�7���ڷ��X�o�p�b�#_dȽ�Bc`(۞������PZdjv*�Ǳ��:��+��F�xX���&٩��9	��7ķ��e�"��QܭT���n		I�W�����U��-�"�hM�j�8���N1���KxX���Τh�Zy��oF.SV�#0�+��E��-ԭ���
�1r��^��*��걱wWiԤ����o )Z�)�9��Ap����ĩ�}aN�6n0��tNRJ���ӕ�.{�/� ��	c
xQ܉i$V3�����Ud܏i�0�`����^9޿��Dy�E�u���Nٻ�s�Or��=:���,�[X�̯�/w���ݽ�:�ջ��"���NG-]��d�.��cu�Μp�]�C{��{��ʯYK1!��u�����f��w��gN��ג��ϛ�\�9�v���i9i�����" ���	�������X��5[O�&�d݆���3�H��0�C�n�}Ffj����h>!)�m�/����˦�Ѷ'�Z���Ztm�z\Y�o>�7k�)V(Ξ��TV�T2޾
r#ktl	��w0��n@��꼱��N��P�	fF(:z%S/��+Q7+M�����iyEa�u��ZM4'=,�M��3s/��a�T�F=�&�h���z��H����md���^��F��5��e��c�
=�&���LJ�3��8+GX�x3�+��g�ѵ��[��-PO?K����+��5Pf=��8��]Һb�Y4���Y	)��r�NEd��S�*����ݥ�%�"��z#��Ws���C���+m�ˎZ�!�D�ƅ�֎�^i^�H![�lL9�N�.(��ت2�8퓢/��M1h-�de�=�Y�����㜐?+C����Xc�9qf�3s��!ք�Tb'RZ���ԁ4Ѕ��<�B��}�t�����X+�[!��_��!�axbZ|�����ǉ�w=0bȠ�	���&&�,E)yPh\	3Pb^W]xo����.G�t��z_v*���3�sd�57��-�`ͻ��g&�6$�C.\r�FqT�X�&w9���0F�KO�|s͇2�/�g/Jۣf����PP�6��/.��R�M)�N�b���g���<=Ȟk��C���Rf����C��'��T�'�*9r�*���n�ׁK�w�IX�k����� Ly�"����k��%vVq��0͝����:�˔\ ��ʎ?ϫ����i�缔����І��bK�� 4�PT	�"q���vX��i�O0Hd�N:�1k�}��\tA��-`�4��0���S��w%GH�Y}$ѓ.���Q��>b챜�fj͙����x��/���\(luÛo�I�8�%��v'��v������4|x�,c�_G�T#�ԥ-.{)\ ��@���4<�ϧʄ[��]�p�&��zC HaM~�_�j��~�a�`/}����0H�t�����e�řy�+i�d���F��αͤ�\��=-�\�*��fĆI%���ֱk�y.8	$߲�/^no�3-�&�����ø1�FbXU5����^o�yY����������^"��Ǘ�Lb����f���%���ߧ!m�N��u��p�l��΍v�c�2�s�;.���^��Y�����%�h(�p˵6�Y���ι�v����1�wD��K��ʷ���c�wn��F��Tچ.y`V�Zn�-�S�� �n�r��άW�L��,����WJ���+�����wI�);��]0��_<o�M�mvV�f�J�ӻ�F�G(�Zs�m��W&Cbl	+�eZ
��6��`�XX� R���0�:]ru�5KΙ���ۮ�̋kz�HJ���q����VY�Ew�Ը�]�>����������$�� ��6��)Q.]rݛwt\тq���m�]ٱ�>��󦝣����of����5��]�θ,���yI�J�T���jSb��\_aF�4�="v�D���C�5���Ũ2MDmM�7���,#K���Wx&��U��w�D=��0SJ�k�6j2%�CU[���4�r��~/V\��@{MhHE�3F��1M� ���v�͒�qI�wXv�5(�J$���ִ#��9��.�n�kɶ�[���	IY]��WE�sltk�d�7�,+X�b<	�����g`��"���\��s�]b�Up�v�Zu
.���v����?��2L��7��o�Fy�4���ζ��꽲hpU�c��]5dP���	w��ΫN�0=�����&�4��A�F�K,�ņ����vy���ɮ�%ݷE�IVL/j �yu�W0F	�³+jc�����C���pk��SePs��_JT������Kg;t�tw�kR�۳(ݺΊ���
�.A�Xx�je�f�ѝX��ي� �IB@ը��e��"���.�"�KEۊ�ަd�n�O�/�7$r�&����e
.8���mTQv-�1"˅�g쯯�����O��,�b��A��$��b�}eHrd�G��OlK��>k�Im�Em.q�][G��lrr�Y��3>��:!��� Z+9�'���UFS�%ݽ�e�97wm�Ԝ�-έ�s<���m���F\��7F���	��}��������1m����0����G5�<�}r&^������˭���>~�0��ݬ�
D���CF��xͅK2a6���||C-�o�N�7�:'_c�^����zee/\�o��_�0"���ȣ�k�����WW�Y� �C���(J����u��ԧ�mZ����Z�v�ڏ��=%)��"���K
�kM���=E/�""=�n��EO�[9k��A��������9&Gkr�ߪ��ۙ��$t|6�;Ȑ��V�=�!k'H0S_=w^)mly���	>;K�B�5��9��������+�
ٞ����*6G�G�P�]pu}��������KSC}�b�棨4Itny�쌃q�pʜ�P��&��s٦n�31�A��,����U�*��^j�þ��(��q�(zoC.��ە��}0��xlaӤ�__�⍎V���yvf���I�c�M�d;D��F���s���qa�*�x�}hN[Kp^\dwRAȌʃ0�6fr�O�ikWь�y#�4�Z}���9UT����U�����o�͒I����$7�������h��*$S��aiy,G���XK�%�����ke������̮�Խ�Y�)]�L�qK �H�A0���I�,X�j$�}j�X�ȥ?���G���	��Ɂ���}�4����7�H����A
�u��gP!�S���S�]Nc�NT�UlaƑ�N1}���v����3B�}8�Ը�Y�zE����N޽0����s�W�,�@`Lϥ�/k%�u���{�J����Qj-�>�'���ttJ��6��$p�^!�a<g�1H���}���$�˼���<5(��[bຈ��lP�t���)G�j�y�٘w��$�TШ�ԉ2�ʲ� eVTN��g��8�73}���H�X����G�Ɯ5J=��.��#���xo>�'����.;��j��1�����}�J��y!|�Ŧ$'*#e1��ㅌ\z�'���z�Vpfú��g�+v�`+�n=VT��̕���Y"�o�e��ʳ��PQ9�����H;��՚�l�wdڍ�9�R�R�;'�C�J0��>�����K����I��څ~��;�l���-2�gz��f]/���Cjx�@�]���+VK�� �x�
�o}���c<򐜻դ��/!��y�zZ�d*/x!����^@�V�*��9�fbc)��nD(E&Z��%$7���Z}V��ό��\G�s&��#�үw�S��2�=�$h�
x�h<�����g�<p�l;��?Uԧ�.x4���r��װ*��aw�;�[�w���� ��7#I����\}��%�,9�O�:ZoL.5�O�Ɗ��s1p�؜�'�q���1�W��Z��7�K^��f�&F�h!�Ì�4����A�T�^�x�٤�A.�tZ�jP�܌]o��T�lC�;�]{�v&�'oh�<J}���k�Gp*A+��P�5VJ�����G�f�a9�e]ç����?��Ŝ:t�%�FJJ7P����¦/���K�8�)�	�QZ�LUveJ#��b!M<a��r�p�X�(/���n�d8�{�b�׻ѵ�w6�.���Ŗ���W�H���Rf����C��jak/�3�`�Y���B�a��q�_#�Rb�g��%�*>���jg�w�8F��=��Q�n���ث
�]{ωm�+[PQ��>���\x�W�����ݖ3��M�s3|$�#�s�	1����6�b��:���tT���0Lmq��Gǎ��=���n�E���!X�И���t�{�``#���D����	Y�;���&�Eg� u�+���g�i�֍��	=��[��-�q�_j���sKȍ��q��.X'^>ʋ$<y��X�Y��Ո��Y�ĭ�`CCz(%��G���x6�F}bb�s��/��l�B�i�a��-=��E���u�u�"��[?D�^�w�� Lt�Dɡ�z�������{]��^>�����C-x��da�Ǥ0Y1�F�����nW��nӳ,���PK���T��*��؈�1M���d�I�FI��nAX���ARӤ�Or�L������!��&�m�Hf�?KX`���:�Q���L�ʫz�"�#e�3	Puᑨ�����T�G����m�����U�̕r�
�q�Ŭ��e�j셥��R����I�=��Oם�^���#ðkX���8�Y���҆g?�G-��������C��V�)��CW�L�?T��\U�{�g�S�g��v\�ºLcϸ/1<ǆ�kk4���%�s%�uD�>��[˦>ǹ�-�x�)�AG4�,��9;ñ:�˜��򫎸=�m �2��z#������G�k���x��hi�ZI��P�a��Ե��`�Ơ��db�«�S2��n�$��\Y�f�a]kşZI�y{�oe.ZjOKU�:bf2v"�*���,xu���#>CJ,�g�vm�5�`e!�1��a3e�N�j$g/5��<�հ�?�~�q]q/mZ���X�J���I������u~��+{%�5lV1�^#=l#���i�{]����~�aa配����6��(Z_�E���Y^*����wg�i�;ZԠo�,�/�	��`R���\*S�<�ӽ���s�;0����wU]�'W�69���y=(NӉ���{��ᭇ�H�ϊػ�C��KP���┆�s�h�/Ͷ�%M|i�q��T ˬ9t]ƾ���⡻�l\�t>8�x���bљ1;5�CL�,�K�1a�U�O��8�Nr��c���)}�G�4�u?{6�j���t�2�<���n/H9�
�Q�Oj��N�Z_)��W�c��%K�i�����Y~~���%R�����s; �+��%�q�Tx�ڡ�����=���x��gKHh�Dl���䃋��5�߽��k�#Ǐ��Rb!��:*y�k�ߘ񣇖'��Xv����}����� �[S��
-�	妦>?k��=L�Vno��i{�!���腍]�N���
À�R�3A�/U��'�������w�}S(�eR�hc �A~����~�y[�#ǈ��c#�g���\�'�>����2h�^̪���"�>�UG�.mX��X�n�.�P�2�7�ǰ��W�e�+���<�����yGĝ&-BMBq�e���r�{���u�ڷ�YO�U������%��uaޭ����t�;WN�2;ٰ݌�i�	��'�U}T�sJm�m}
���IUS�t$���P�3����H�,tt���*�)LL�q�6��O�Z�u.>�0J�z<�~�m��~�xѫH����?i��HpDؙ�*�Ԟ��nXX�3&n^ԅDe|�i�����_cq��нK�\����|�oI���;�^�QU�Y��㥍�8u�,�K^�NZ������.��)L^.k���	�AP�@��pi�A"�Ӓ/G�m��^�m�_�x�\B�1�5�!dA�c*��-]??/9˿}�VnX>;,�1w0}�`�)�r�3��OOze�Y~�ތe���p������a��.3�/��):���4��7׾�<��ό���͜#H��E�9�4�39uz�X�.(�oK.kVĒ�ײ�3:��c��ti�ݫ+���t�u����4I�k��'I,�ϲV�qs��@b|BUXjVu��RpK/�k���ư��	���A)a��L>�|x��g���&�Y+T���ɗ���$a�]��������^t��Vz�~�5<{@f��s��u7���P�e�5�/+$��q|���g,&��[O�\CU�$��I6w�l��!�~�N����`��u�q}1~5βT
�,ZԃZ}z})��3�;�֝d����XD$�k������I,[�a�z��}�oe'S�3���KƎ��L+^<a��õ�H`G\A}�w+}��ݕ�q���ְ�SW�x��[<z֞��)�_�|4a�B�`�E%���T��㔁��!V��ᶛO3s���K�B�ݘ.�=Ȑ���rM��;¹��*ع��x�t�1ѭ�v�_Z�N�켯����a�R��E?���.(C�9CN��NM��������V��{��ͭ��)�]��=�J���b<n6\���Iupň�[C���%S���䜷�^^����[�ц�������@��[z��)@���z�}����v���[A�V})���!�ވ�C�F�?��3;�)�e_L�h�x���8ޘEy1He�Y�lN3jcg�\V�XA��3,����r��K=����{[��9�[:�`�-�P��ەO{���h4��� �N�:0�t��7��$I3[.l�D&B7�s�Cua�!֡�	I�	�KX���11�ޚ{��H+������D+7�N�v6I'K5D�(;�r��{��g��?�>"��MQ�/zE�z�ľ`�QŴ��Nu��
AW��z�#�w�w]�ʝ��V%�F���h����͏_�_�Mӣ�\,M�v�9�t��S���Þ�}��t�;���uޱ�c`���s���:/V�͢��8�d��p�IgMvn-�n���|�f�t����ǣ��8&NQ��n.��r+��Y���AvS��`,��fA�/C2;'�
��|�5�Ā6R��A�
�%�L��a���ʌ,���h�7K �{̆l���������tљOCզ�����LU�&	��ٛ�Jꃹ�j�N$�zO�Vk��m�1:���"&/�p���.Y5�5��
�|��zl��E����T�Z`�V��֗^<5sӗ������$Q�Pt������*m�#*>y�ܛ��㧨J�l�_d��[ʇ�j!�ۿ
t��Oi���7�acR��X��s��b���gS!���yl"���R��y*/����ЍQb�3
����6�!/V�cJ��G��,�2�u<�ʳI�)���'�q��� ;䡋�v1��*VJ$͍�J$��u|�ŧ7�։�\�{b�kV���t��m�:�R�����>y�uR�S�;x�'��������Gsr㬑��qֆgi�#��^�=C���G'X�C8fKM��d#t���-U�[ܗ�3KwIP�ə�h�l��|�YR9g閕���WO�M!��љSVe��ّB��E(�˙���;u\p���gj�,n��{��쏍C{�ka�wJc��w)Ť�/k�CO��gQ7�Qrn���%j1�@G��Pܤ��)l�b�↖�,ݬטx��'�/���:�r�1�%�7��I�ɢ[���\���H*=Mwk��
h.-���I-��PHWYW�p�P��76��J����b�y�r(
�V����[-�ϳbB⏱L�yYy7���"m#�YM#�Q
�e�U���}c�v>��=2픳�>�F󩨹�S"𒚼�{�{mW��]��������G�g���R�1��u݇Y�'�ow[L}�rn��\���)�lC�qƪ�����,�>>�Q��^J�!ԫ��$]y��ɼ��|��(�]��vy V0��r�7՟�=Ҩ��+��~��'����Cl2�s��Y�a�N��p�Ɏ����v;��5<��=��/s�}��U���v�%�xxzGNJ6~ەh���K���T"�>y��ӟrd�۬����(�^J!P_'̾�F4�Ϝkj��w�I�!�1G��l���Ƕ���Q��1�}\cf�LE�u\j�gEx���5�	x)gHGK�#��7�7jrL��B_7~�������>8�^l3�[��N����P�C��y$�����b4����������=��ʪ��3qդbD��l�\C��DC���r�-}��z�{��Xl��j$x���.�0b]��iMT�y6���*��oR*cS�r�4��c �j��^=,F����,�~����N�ѿ_�U3Sq���YU[�B�Y��ϵC��Q.>���zq�L�+��M�zsd5��/x�N�ݫ�p�x���Q�P3�Q�u�j����Ӡ��a:��ea�UK�>,�&G��
�0�q�!�ݎ�7��yBxu\#Gi���7
��@4Ԉ����Dd� ��+�N�3��GL���m�]��ԫ��J�Q��Op��H��[/�ڸ��2殮���/Jb�btqSR����$�]zZ>1~��"[ &�xLq�j��_������Pj��M����+=����u�fw������NbӹoO���0�x��5��A�|�\on��x��.'f���ٽ^>���9��j�)�z�y�P1�,37;�<,�}���G,8ghv
���~�B�k]�P�y��s����F��)�{>8w����M 6���Ec�1�kz�q~tM9���
�dȳS34͹;v��D�P9�$�&�i�E������l���w!������=��u��4�Wo�34F��!��@�0:F�1�����[ɛ�+����k�}A�8��bk	?@8��{��L#?_��FFp甠hJ�T'Fìu��g�+��~M��Uxqګ�������WY��6�ő�aj��9 JL�qou�g�fR�Q83[L�>�wb�z�T��w����G$��w7��ɬ_etNe�LRܟ�@&��;�{�5-<w�似/,f�RεT_;��n�/+&�۪Jf�%�Av��ڦ.4|P��Ƶ��I:xw�^ǚ
�=��R�׾YN
�9Bo��hg0�\����z���������'k�g�2�$L��-�yp�n��]�<M���NdU��;�]��a1Y��zt�!�!x��'�=�OM���+��/�	!��a������P���"\婾�P�-7�4�3�x�z���H���B�=>ld[�X#��Q���<���i�e)��
N�Lg]�̛°�Y�y�H�6�GW]���NV <���G�+�4 ��l�B�����Ѣ0�U�*��o��bB�zF��_1��-E�O$A��ar��#�a��ǵm��]��Ir��R�H �|mSl�6��Aifc�y�Ͱh9��#��{���kQ���=�(����͹���䐈��~DDG�k拇[G�.�^[�s���TLe��˥b�_[��t��j���dU%�x5��c�W0ƣI�?."�l1�ǽ坰Wq�m�r�1:�D
<�jbS_y������Xnʽ����N��L�o�h��H�	�,I�NU���if�ٹ��'؁\ŗ��/㚳P��E�1ŮbU?� ��_t��kdzP��ͭ�)ȗ0q.uu�53{*�D��Y3'�2���l�)���3z#!ŖP���U=�+3�x��q�B�.i-4�'Hc��2������%�����%��5ȝ$�
�ÿyi-}|�׌Q�����z�=�]��C<ޑ���sʋ$��.<^0��*���z/7�׻��О'��9u;(Ы����9��{@�'�_!{�	��_& ��6k]�@l�M�g1+JD71f�&�B�Ň5���U�&��J'*r��'��_}U�����EO�c��P�7\u��CN�X��F1��Jn�N�7׾�bX���du��=3P���I�Nj�Ffd�����#�Z㚸�Hy�8e�A��%l)ߋ���Ј��%ń�&�R��1�^#=l#��ֆT�闛�<64_܉Di�1��^S#֪����;�t�pP���$�ix�(w>;��ג����0?0�UT%Hj���i��{P��e�J���`��c�����8��淧�З雛兡	��ϭ����i�l\����,����Zĵ�f�Mv�&X�ڌ��~H��)��.#Oo&0��5��w��Ad���D#ƹH���(�s^�p������G~q7���r8�F�1�k�uږ9�MZ��*�3�$')7q.�$2ʤ��]+�栺qʈ��`�nЕ�m"#h�w�s«�[�{��-4Z��b�U�˜�Vǧ(�Byi��2A^Q�W����7�F˵D1H��"Eyf-,D�6[t�=3p[���qX8᳧E�H/�.h�]��<(��n�@Ir�]�]=�(3�^97��԰�>?v���R(�=�f�["%�_����t`p��1O��A��$MO�l؞�!���-�\Ȩ��Α3m�� *�9��OeT��IG)_��n��R�fe!�V��_��t�����V����(<D����YC��;AcA�~�N�оξ�y����Y�����P��� ��Y�:���P�h̾������P�`7��yq���c�P=D�������KU{cʬ�vf��� �Z��U��%>�m��Ī��VV)��v벴�I�ڥ�VfmGieä�Z����W����	��㗨NRNR8�>��	���;6I�ѩd���T1�v��UM�x��H���~�{s;�����GO��vӤ<��O�Ӥmc}<�K����0.�Vzk�7&�?=A,��:Xиث�~��Og����P�8�.��$C�Z��C��ey�s�G��nWgyL"�@.<oˍ��Ƞp�,�+����t��r�����)t�W�̞/�M��WT�Z���R���<(ك]{���J_�9R�����Z3P]>
�YZ ���W��I�g����3�M��Zó���zע�G,�4�����:QH��^�^�*�TL���7���=:f�g�B�Z�s�A��9>~�ǵ"H�/��I,�,�c���k�g��@�i.uK'K�h;չ��C*Z|ɶ/L����e����ɺW6rQȊe��U�9�hM�3�spȴ�+�T+p1��Q��}_}UW5-�����!_�؜���te�R�uP6=¡}I;2��D-�{=�����c���Ѕ<�;D�8t�V�ސ̬u2U��n�`dxU;�G��P��x�Tt(,�xC�{��f�1��E=t4�*>�H��!N=,������]�L�O
6-̍?|���9���R�b��eş"�6���==�ᐏGZVU��,W�j4��o�T�ETm���%N���9�Pd��M����jbGP_/��B<55Z����yT�&��m+57��Ͼ?KXd��C�u��ʮ����ք�O�Hx��M���Xc#Qmc/��J�=w��$�ݺ~�{��F_��^��P�Lv"D�/ʔ�H���Jz���6�N)u���4ʼQb����-�<|��'���g��]7jf�ȳc��E�y�V��N0�|��jK�n)��l[�J�F֛)|z�_{�Cu�\V�}B���!T����y�9���8�q5/�IzV��+�;�}�]ր��0��fV�=o��{�e�����r����?҅�y���	�|t�}|�N��f���s�6v��TfE�GLȯ:0Ĭ��x�$I�u�^w�b/
���m��԰�	!E��H=ZZ�$�=b����Hsp�UK�Pg$���Z�"�3e�N�Z^5'��H� � �gu�뢅,��9��t��.�1�Eg�&>*OR_z��^ �ы�:yR�Ә��.��▲�k��vk��<�3Q(�9���(m�OŋCl�"z*�.�r����B}����:rN�Y7N�"��|g=nn���0�;絹%g})���"n���jIunR��<��W���/�cO_�l��<����9,�y�v�V.����c�TNw$����K��!}�s;==0 Q�ܙ��z��%�kG_�NP�n�󼆗�gb������Il텙KQ�u�:�"��ڙ�t�=�� iO�+4����Ń�����yk�����+C=��!M~!��<7F��,v,�Gێ (_����q�g�ݭ�0p�a�V���:��x��)ƺ���{/����u�d�t뭕=;1���x|��(�uӿx���1g���k�,��dQ��4��lFה���I8��X�!yݵq�{�y��z��G�ٮ3��Q|Y��Y�F04�
лIk.D��~�fc4Yu]_��d{E;�6�Ϟ+ZO3|
O��~'���BO�"f��oOO1da�Bc�L}�sf'��VÕ��`kdOA�h	ԡO-l˗̈́�Ql^�Q)V�l�q-ѹ{��[+
���y��]lI86��}\;n�Fܙ�	ά�h��h��q
{�Ϩ�4q,�=�Q�|Ժ���:��E�J� ��d���N����K���Uۧ�e�55>z��A�<�A��� ��i4+UF�����o!X�[�4�wPZ��=�^ h���ۗ���5w�b��M<�jۨp�c:	��JF,�]j�f\gQ	�fZw"u�ϊ�,���^.�,��.S�G�`^Z��V��:D�+TZ���8�%Z4���F��S���o�][Z�k7lan�~�<J�s��qȞ�nԬ����v�^i�hT��u�k 2�}��Y]��/�Ҍѥ��J�#�}���C��㳳�= �n�S9�ӝ�vѷG��]q�U���4���|�z��e�᪉��m-{�qaqV��R�q�p��A��\2Q2��K9ˬ('�[T_Y��P��N�{e�oE�D�)��utg����GA�C� �kxN��5���q-�)Z�{	�c��:��i�~�e^�;QÙ�I�%��]��#N�\���{��m;Ch�J+PE�uyD�ڒ�i��R�^-��Z�,�Ѐnt��kh��'��bt$k㚵+9(m���[ј�r�4i9���s{7����"�K�"�|9�� fTnc�4�__D"���CBO8S繕2o�J�hXh�OUr��]�����PY����ta����fwo"�L�Y��'g>̍�yI�"8���
�;Z�LIa.�^��K��q��V��T�s�	ܓnl�F�N_vƮI҄:hݥ��m��by
�(u��7��~��~����Щ3��@��"���Ğ_>��� �<��Nd_s
_^�y��>}�}�a��G�s�"/�~���>\J��I�es,�}�}�������|��~|�Wh]�=�����#�ourF�cm�E��!E|�|��Z>{��.���#�.��o���J.�L��
uqx�_m�y|�/�d��7�l[�3�n�þ��_-�A{��y���c�_�~�7Y�2��!}}�ն/!0����`�^��>}}U��/m��l^�Zhګ�^��(�/T�Z.ر��rqX}]��c�$1>d>��!�^�����瞽}�Y���:����aG�}����� A��'����j�8�!��_I�]�V��=Ȋ՘�l=���D��n��|�lc|�K����9!�C$�7*�;-gOҥ�ژ>�jU�yv��=��u�rǙ4q�/�:�E�6����߬e9ۘF}��h���n�Oݰ��}����I�h��|�?,C}�ەO:���uu3i�9�p��Aҝ�j
�r�w~c���ej��!eIv/z�%�<{�T|����gHB�q�#GB������]7�O�r7[0�*�����'�PGo1*5��q�G(wt�����oN��Ma'�� ��Oځ���6�3�#��:h�D{#��RD:\p��/�yj�������^�Y1i�ZC!�"X+��Xw�6��ue�u��R�<�׌����M�WT㤞?\D�[�D�EV*���-��b��X(F	�;�pM͙�b
�1t%��i�gW^��fS'8t�j3˓(l"�ʐ�͉F�p�������[��NEO��xx�ô�� �-��7�Ԅ7�l\�(R���;w����Ŭ#F϶ߌ���Vd�@�3S��O�ͪH�:�KQs��'~�R�\vv=:gڮ6v�ɛ���e~6>��m����t�~�͖C~�:If�e!ƻ��.��JJs�ɑ/��՞�7bgj�]s��E��"i�ƗrTk4��EO
�3鈴��n�7B�@Ţq��I6w�&��Cҷ6�N�x$8�'=�G�����u�6�
0^Q
���\�)�캊s����s31��f�%W��d���ϟX�y��]�4.�A�<u��.4|k�u�6׏l���k�vgw�,׹��y�)w ��y����>5�.���f���=%�
�s�C��G��=�EqyjY�Q����R�}�⮺ӫ�+WyhV_Q0���7&#w�=C��%egu��5jN׭,�C����`�z�������*{Ý+�_�cX���bXy�"��/���˾)�Y��ow&����I��J�]4rs$B��+xs�`�J��団����uk��w-��&p���I;I8��U^i(V��Zp�L�*==/����W\)���~�h�D5�˟�t�K�Jtzy�/7�3�R����8Ze$��Y��7	S���y��u�;�`<)/.Ě
�^ry�i�"y|FS���W�KI/�/���yl�9�janC���Ŕ�é�qmY��.=�<�I��Ό$�����*R��:�<�'�W�%�c��u�Vz��]uw[d����i<�xO8Z����=�#�igN��>#�1�P��f�֝�y�Of�r)@�T�+T�){R�j�g&�f�h��V�y�܅O{پ�w���B��l8ВNZњ���%��2��3�䍢i����O7����?���H�H����~"�j��R�0X~rC�9��N����to��B�}�O/E`.cּE��AէD��ٽ��Y�r}���LY�!/���y$�&y'~��Td{P���/�e<v�S`@ �[����^T�Mt���\Z��yg_�L� �yi%�Z8N�!����mV{����9�A��\�;��u�@�w���E}��x�!^������KN9��¸$u���]]��N�o���B�ӈ�a���P�ִ�>��
Y�t���[*Un�8�N;�92��utU	n�X�H𫓵�Ƚ
��X�7:�Y�G�*>.���]�D��LZ\lvK�n��G�lm�����zଋ4��_Ǉw;��q��k��m�`���I3Z��P��b��}��m�7"o)�}#2� Q�t�+ Ԋ_D{VL��y."�cؐ-8p��P�<x��TC�⢯m�p~���0z���CN
X}k�g��Q|~폍�0Ń\ʹu4Q��������FcU���r���
wv���#E�+�ҟ�����z�� �ظ�-=�(�4s�-�&m^��XGsc�Cǈ��RB�ϥ�>�s���G%�=�2���x��܉�����8gicA�~�ʅ�u]���Cg�b��E��IKASh�$hya�*/�������ܽ�/+�
z0
<��2��%�)L��)�IvfVQ��;�������,�e�Pn
ꂟ��6���*�����(�k�� M��.�3�m9R�z�j�G��׭u�e*�9���=qaC5Q�]\�3,hsVT\��\���/3��+�`Yg�M�Ti��,� 8����5��mtbb2�+Y�4q�@�K���v�Jo�������7"��J���Qw�g��a��w簨쑶�-c�Q�����D��-��hJPr�=P��n^���uh�[�ș~qV�D)�æ�i���B�Xg.!�Uv�G�Y���{�<5�P��a��O�H�:>8I��/��y�r啝�47���L٢%�CP�3�����o�f��Q������L�b�I���8v��;���Pf����.��<�n�eD���:�Pi!ߘ�XLVw�N��vF�����B"�Y�9>b챞H�0��a���<�J��ț�x#����uқ�q쮟-o	��yi���sn�*�=��2���>X�ַP4!X؂�8�å���|Ǘ��%S�].��/udxN�5ـ��0�Q��8�J�-�lk-%"�ZK�M���t�/�9�IAr[2ʄӼ��%�1I��������x�;��C HaW���Z�%�F�Р����n�3ʽ�q��L�� ��k��O�Q�
G���������
�jpDʎ����uws�b�S�S�Ny�!5�ʛ���q	5�h��>5��(��k
�i�li�B��j�߈,�G�չv�Mm��8��S�Ǐ�X����g�(%��LAؼFN2�T�����D^�1m��G��8��h��H�	��]��7��C��'ڪЮD��:p�F�<B�G=����W{��yk�ԕ�t����1q�ښ�8zv�mZg�ģ��r6�׹џ�!)q��:=�!�����ۂOe^{�|+�S�*����H�U�"%���F&�Y'e- ���S�S�#&t��w2o\j�@bv+��r
�"B�bo�.{1�I\�\2�ܙg0�|F 㣗���j}sju�R������]��rnT�B~�mLn�z`m��
nU��K��'li~��˿e缛$�Խ�ý~�^�<���r$�yц%g����9��g����0��+-x��Cf?ED)]���V;*�/5�zJ�ߩy�ʌt[��\Z]��h\Ǧjm���(�N_{�$���n"F�������~"�[��{�S��"K/��"Eډ\���ZXH"��>^��:���Ԧ�#���o֎װ+�l��F�asCK��?G��d������rbW���8�YiW�L�a�ֹ(��}B��%g�Н��٧N1SulWg%�FN�&էnQ�՝�F�h_���Fٽ��{E�!�a�B�'�..�IF��Ō��WuZ�Z�V߹��M��"ᮭ��i_RQ�TT��:��θ,��{��pJ��0k��4�ĳKgg\�;["U��PB��M�B%���pw&�*c`�_��:�JB��"��
��><ok���Wfz٬���j�������C�DP��|z�U{�|���-*��4����'����Ӎ
�3�yg���j��>j�me�[&mu�]�<^��:�Ӆ�V���4N�}�1�R.8^.=JG�y*;�1Ѻ�Ĳ�����\[�/�Û������l��70�ڜ���9ń}z�Qx��\��8���)��=ĉ���k4ɝ*�|�ۅi�As���c���zzy�!�Vb����TsZ�/|�<D��[lZ�gǏ�Tbz%�n�>MeTÃ�e�<���8ЭH�8gicB��_�#4��g� �}F�T<�����8(7Cn�Q"j��l����|s]V�
�
v���gLw���� o�Fe��I:���᭺��d��^��MfG�NA�H�
��
Mc�Z>wD�(�&���"K��`�)��2�>{�|���J5��1�9q�s��c�3������'�O�����,�aӜ�9�6C:E_l$&�
]�����c$>���<�N4|x��m?�ƨ�a�rHeS%��u��ɛ���F^A�U�a�u�7N���BNG��E�+,��ZY�#�����)q��A�}i"�	ѹ��j��>7�+�I���Zo��Ƞp�)�k��w�xz�$E�����KS��<UuN�L]�k�p+�ђU���^h�3���CN�/��.��d���*H��߼"j�ä"+���_z�8w7�8F��"���k���a���9��P#e�p&����(t�${�۽W�Q�!V7`>��W3u�t�nJ�!�F��y[<���~��[{���QK��6mֈf�N�͗��n6[�ݐ̺P�3Y��T� $ؽ��r�sd��0l}Э%,���׆�u�F�X�wos�
�;�Tz(�7P�eakX�ִ���`�M�z5��WJyw�'�h\-�M��0����ݢ��%��M�/`�X]�1f"Cr�N4��e���ko��=Ǯ�{����n���{,�}dMcBf�����sa��p�.*�peP���W!��9ݲPp�A�u�p�O���F �Q��(M�)�a�Wy�.��Ɍ�.wtH��mE�-"9�[&^���4�h�Γ&W+�4Mb8%^=x�4��d���Es�����RZ=YOLi��XQE,�ɢ�=��_pXZB�+I})�ԯE�Û����sd$�qu�7���gX]8�Mikt.gn���}Q��5a��#V��34�3bV�Au��&�j����%�t��%���x�E���;e��sc�]��J�������S.YcZ̚h�#r�}�3H�f�ЦJ>B*߷1
�(im�u��ef��h�	}���&73(���N�;�9g���L���0&�9n����;�f��������Z��b�Yt�읹ׁd�z�l�����f-�!�J�Za�q��q�D��w=ZBp�ΰe�m����k�4K�B;JuZ0�`��k(u�!.�ʋw	�--��C��|��/e�f�క�R�z�K�YF��ft���'�˳�ss��2��������i#r@�]���NF�z#[�*�L�*}�&i��7Y.M4�n�r�+m=G#��,�C�t�)G��-�~�B�'7��f���f3�$��p?^����:���r�zZ�J+�E�"=�uS���?(����;}�}��U� T��k[����C��!�&��9é�Ж�K�N���>K�b�뾷w�@�"=m���|�����
S�Im��
>��|?,�}Q�M4��L�-:��}cy��G����;x�K����I�}�o'9�:۟#6�Sm�;�n��7����ܯ�BQTU�
m��]�oe�N�ݜ'v+'6�'�wn�8��p���M�w[��۪{�yS��;�$M�X�ϡ-Tg��zUnzԧ��f�:enm��u���&)F&FJ/"�̭�L�"��RMz������wN�qM�}v���`�!��'�\:w�H�Vs�O��c9"H�/���3�tv<��F�]*������r#U�垣v&v�\�s*��C�b�������S�>#҂��<��ַP�H։��2�z��7B��n{�]�u�מ"��v��;����B�MYs��<y˾�t�b��兠������]zv�}n��ͧed��)��Vw0H�I|��$=b?%�
^.��e&%���W��_o�٣�Ŗp����!�5�#�ͱ�+�i4��l�$s�����b�6ƞ>:{ÿ����I��(��U��A�f������J�N㪸�>_q�oM�����V�:-cV�������<�*�}ePe̩AӼ<��B�չ�u�c��ڥ��W()ޯgX7�[���KA[��c�aMIy�/:�8�>����⤺�������-V�+�/P4��$�9�5������h�Z��8��J��K�t႕�zX��?G�+��"}}y�<c<9�Ք�^1��HJ\rS��y�8U�s���w��E�
W��)C�m|e�d��i
��!���H⻦��f^�ޜ3�kf�x`�~"�|r��3ȝ$��4�*����;=3>�[�9[�b���<�-�TY�=nfy7��|{�ݖ"�ҰZ�`���^7�!֡��W\ںx�~��h�"^��
X���N�C��P���D�=΍2�`$Mo��H����?V�0��T�+�����.^���x]�̪wZi,-+y���й�n�H����m |�a�Ƚ��\\���{t�1��T�X#ٕ�b�+�+v���.:����R�)���8��jյ��JU�I��iD��\%�)��c��u�~�#X}�ض0�����s A�,O5��M�)��Y�Ȣ���O�;C��Ƞ#M�ӱ�k�%��d�2�;|B=��ң�������&}�-"cd��eL�ge����d��|��ϐt���H^�F�t�|b��m���hlWmDG�/!���Hz������2&V0�b�����L	����{�!=�C/�E����_g�RrjY7�:���
�".���tU	x�׮��I��ĀJ����*##���G�)Q�f��D��H�-�������"��*"�H<\p��q�P�.Z��AC���F��B��L8��^0����短Q|YOWcU=,'�3�+}E��m*l]�ب�N.{���C$}srn�5��mۋv��^V�7#����^Ε�5R\�v	�*�7���k%�
Z�FҜؒ���%o#���#}�K�c���%_[�{X�^����p۸�>�wۣ�Ļ���{WH��g�I��O�qݷ��=f�n��G�aO>��36A�� ���4����ʻ�l�5C�Y~�"��qW���)�y�&�w�����:W:����KpU��<�Z�P�Z>wDB�Ƌ�h���C4��W_o~�����:!�2������,�Ɗ9�r�x����=��I�,>��}H�di�-u
�뻘�Y�:����d��;�*�c3��x�qt�x��ڢ=Hq��A3e�缺��а��ā��z*if��w�eϮ�\o�\�N��S���3��\F���d���$C���uC�Ӧ���ź��K4U(/��w����P<6���-e%;�[k$�R�1d���B^����4ӎ����H]�MIݬ��N�������Z�$*GwW^�-cԦ(+%��	�@��N0^=0�!bЭ�g�m�#z��A�A����P������9igG���դ$�/82Q�j�C�a�N9Y�lw�r�iBo��{.7�s�=zu��-:~�t�Oꁞ8}K�;���~v�*t�Ѻ�7O�W��Ҭ�VE;	�A>���+$U�wv���k��y�3�[Ǉ��O��se������[��{6���}G*^}!�kW�r�n��*h��񕞩T���;���6����!��Q�ڦ� �F��w���\\ι�.s�NYWs3FM~�G�ڃ(G�<W�+=�8w�{�����,r�A���Xvy��^"D���w���l��jT�����t��N슱�e��3���z�ܭ���-�:e ����!͉�ȋ�Wz����c�rr�SNc��(��`�:���J���u�|~�l�>7���;.{���fzΆZ�P���77�}�H���K
���li�Ct1cΟ�&eJ��P�����\-���=cX����),>i�]M�9T�{M�����ʽ�-.49/��Xj$rr��g����"���ɐq�Bj'H1:<��3Wd�,Պ%���xJ�k5>ZĪ�|p˧�����q۹[�.u��qc�o�r�u�:�g����i���Yu%�ajz]ԿT}��e��Uic'?��K�C�����}�ݞ�שzن
ǆ}��E�.7�����K#��t�������,$�~T/�.�Ǳ�F�@�i]�2<���Z��_ f2zׁf�+F�(��ܶ�T|��2DWQ��,EnL�Gp)VY��%Y{�%v��Nط���So.+���E0�'Mr��8N4|�������Ňt�>8}js�������`�=�n6:]S�<l�^xz�c{䏈�b-,_�GZb��7��e��N��w��=�!⍘�>-,�H�H�ϟ<>��%!�R�Z�����(�᷐�z�X���ZX_�!�<�Lb��
�0_r�l�W��_L>܂5ǠT]���F�`"�dA�3r�cw���j[�F�n�#%Ѻw�-��3\l�x��5N���כ#Z���	�_4��R��B�.>(������wr�ɾ���XM�GO,zC��Lwa�Z��ӸU�CŖ��m�Oި�z�^Cڸ�R��x�H�@�{��,_��v�0��gǏ1�pL���~,$��C>-�)٬)\Κ����-9�Ɛu��)��J����M%�G{�ƨ�{�mN�������]�[�Y;Kq�ǆ�����Ķ�h��U��R�[ʦ�mc��{�(�h���Cl_���O��w�2�����D��k�79���o�.�ݛ(ߩ����i�
��4D$��M�&�r��-cSSP8�3yw�[0�1��bE��ǩB(�����c-��}¼����{XN��c��������\�^xn���"����\LC�jDH�Z]�-g%K����厦�^Uz�}Ǯ!�-q�R���0�R�3jO�3p��9�ӥ��+-�ʝb�L_�qs�Wچ1�1.!�#Km�@^������n�I2���
��X��;P笚8Ж��
J��f_z�Jw�!,y��>9h+ۚj/�P���I{�S.b��OG@�����e�
}@z&��Q�.��<��K��t��CU��wk��=V���nC�ò#���2��\�w�Za��o������NNk1��D���Sbn�=���֤�Dќ�ȷsS��Q�N�����^;����	dB4�"`<��pVNλ�q0��:�$v����$��x񃑵Dx�����%e���Q�Q;�=�a�	c��T֟M&�Ӿw��#���%��S	>�Y��|Fե��2עD8��!Su�U���QS�0K��@4���Zl�!��3Tɾ��x`�+L��[��խ��P�����sj�so�8�V�J1��U'��)0��,.&hr��j�� ��P2m:��O�Izx�U__������dEu<p����w�"���w��;�T>�0���X#���_hA�(��F�=|�*��*�R��mѹ���c�&p�(���xy7��C0se���x��Z�R��2MWh�,���I��;;*{	�<� Yd鋊�b2�}�,�����ո!)�E��.EzI���e����T�yzg-ex�Jk-e���S�ڼk��s�u�&�=ܶ�z�H�;.)\��9DMy��1��o���yU��s؅f�h��Mrz���Q>`�:`J�OzBH��E�ⶠƴ��3۾��j/.m:��ZXAa���ҟ��H����٪���fo���}�� �H�ց"XD�W�)��8C�5��u�gT�p"��̋2��c���7�*�� ��sCXjM�;f�>��Ii@
������i(�WSm�����7�0(0�s���$lu���-c�34#	�f��W��6�l|˺�Rw ��ԓ�O}3A�e��'gk;q�zh�M�8��Fu��cV,�5�Q*���oX�l�W���}Y{e:r��C�y��_x���yhVv�N.{�9�s��\Z�Y���6�s:2,B�mJ�n���t�/��3��p^$���R����Vt�ruڃ�O��J+0�!kr�T��J8;�6�EA:v�T��o�8��"��ʃ��ҭ�3Wγ���A�����,i)�]����Ν�3�(���͊����u\����Ke�J��]�f���c	�+0+�,�;FT-�	���.әܨ]��o���L(���:��u4�24.�]�y��V*�%4�<�91���#y�6�ŀ�ͬ�2;]�m���-͚\w&����y�(��'[�Nvc��(nؕ���uVJ��g�//,YWfNg)�ڴ�`�o���Ksh.-&C�H�5>U��y�D��s\6tVN'�e��N�ksl����v���˚8�od/P��<h��n�.G�{r��}��v�֭�R�Q�DgM���;q�U��N�L�Ֆ�Ws�]<�=�]��y����Ւ3��We�&P[q��A�jFeY���N�,�d�H{3���]c8�(o��E���i��zb�7����C�u��a1d�o�4F�5���@�H�)P�d*.�X�1��z�wy;2���Ź��y!��A�C��Mm]�.�=��o�Jb�nƴ�J��֫V�=3�}�>���Y[�]4xI~��*s�œ�������˃o��o�#�r��fM��鳦h�-��g2�n�+�_%>��ZMLW��0�5m�rH3����ɇ�GQ�m�ŏ�H"���V;snu$�t��g�y����:zj���NG�$3�_���wWwWw��ݪ��;�tn�O��?��L��1>�[[�E�E������Z��o��S�`��2n��o��ײ<�wmm�3��/���$*��aO�e9VKkĜ�+������"jG�23)�J;8t���˖4ק��|�m����e9|����3�����0�W��̇��#!T��R'>�
'K�h|�J�<�R��p�v]v�u��w�>�kF��J��ԠﱗD�U:�uW�۱��Fז�/lS/�m����W�%KC>�q�}֪�0�e�d��IAGݹ/�����k�/�/+8���9;����U��'���'��f�46�>7�8q���vKkb��GP��/�Oy��r�g��9��E��u���̴��cY0��tE);���z����k2>�[wЎm9CS\
��{�}�b>�&^K�|�
�l+�&48uwR���rli��.T�Q�Ⱦ�
Yhj�G$�Y��R����
Ȕf{=K�O'�*�e����x�ܹ��]�MĚ���π���Mмs�~�Ǎ5��
Yb;�6Hy��>���_���Ã�f�c۴�g����Mef��B�Y�mz��
-޳nSA���'jY��~�1ܩ!��.p�Ƭ�=��W7�R�5$8��[+3]��v��.:�Zl>;�R7yڒ�=?z�vS�8c+S���#�oO��O��d���~��CZ[���ȒK؞g�?Lf}��:�p��!�5xq}�eD�W0K��5���o�l)��͌�)d�����<U9e��T�U�(�vf���e�����g6�B�q��̓mXp�`��t�Q���W�kY�ίH��(�즷�EH����	7��l��ϕƂr9&�wg�jnz�/X��yp#��W��ȪY%���14Cs������*�l��Um{k �Q� �ͤ=E����6��l��^
`뼣:�̙�Ҵ�M�u����G�NI�le��E�T�γuކ:�{V��A����J�v<b\�騺G7S{��F�Ҝ���$Q�Z��dRŗ�#�r,o�����a8�Sh�L��J�B����7�0�Q����wr�dIy�te�g��M
R&�sA+�kɇ0U�q��N�Qҧ�"z�t���+�s�Aq���ʼ�t�k��&g,� t�u�ƘU��J�����n��4�CO��i�O,:��pRH]䣹Axe#�6
��{�x�,k�
��D�	�����n�Ƽ��m5:s]ٸn1@3�5

��K�Ůۼ�ʌ�`տ)�C�YkLh�	�ҭ�3�c���JWu17�>Ԓ-s5�We���b�c����I�Y��}¤v�k;�v����h�e�ܜ��&0�[��ɾxܨ��k�4���;{o;xk:qD��dv�r��&�[::.��զ�Ѻ�=ͬ��܄���<��U�5x�LSVfUFp�o�M�Y�〰��₿U��,�1(K���.Rq�V"�	�m��a]�"'�*��W�ы�i��Yb������{˻�!a-esl�J�WtE��Ɵ���3ب�{m�B��|_7+Z�f�L�mx��t����I>z��^�]=�%�sP=0�	�NM
]#j�PZ n��C)�{��T���w�"�I[��,r�fP��1W,�FK]��2�vj|P�r�k������ŷ����]��i�=�4ey�'��Wj+�ɍȌRi��SO2iFbz�D��J�2̍�w)�%��	�ܦ��@�^�ml�	%����S�ł[qz.A��yªͫ=0��g�Ź�pr���y�M�BVȺ�@Wl��-������|��"/_m�w^�o��x�*�\nu���`�W�r��A�<����x�N(���2n�Fg�.�"����x�
Fnk�J;8�p�K9�qA#B�*ٛ�5\�ʍ<�E�q���̖��Of�y������V��)/k�Z�J*�ݫ��;��BU�ۊ�.xC��bz>�Vi �ɵQ�&�c���
.�2�\�}��i���]����Va��3f+<ԢQ;Y��)��i�]Pl\��������7*��x7W|Q|����~1���}o�R���&�J��n�\}�#����$���ת�{�G%̚m[�M6��J����OGH�w>/)ۓ�C�V�.TnBxμ��PÑq)��Y�`�ײ[������z7���ɚ�$ E�İ�l��� ������pg���f#O!�d�|��d��^^�6c���`��{�j�S&gN:�0S�f;n��6�F*�:W"}Z-��XR�o����Z3[�5描AkBXE^J��m��)�V�e�&wxh���rlܧ�
9z��؄�aR����^�{I�Nh�v�$���eU���a�c����{�l�X�O���lnX�yD��f�`���z�')�n2��:����F�|���q5'EV�/2U����4}�"�Ab�:�l������%Ї����|��+��b6QH؊�4q!�p	��O۬y�7[
yx��9r�b�T�q-�7q(fD���GEǭ�����Ĩ����Z�΅9�������->̤�����Xɡ�a�����zt3y���'\2���{���0���v�����b������tbE=�ig]� oj�E6l%���ZQp�.����ͱ��:$ 56^�������,C���dX�E�[��[�bsV�C)�FGڇ���}����R8�B�Q�^�*C��mg/I~ᚻ�̵�L#�A��dɕ�A������B�tBǊ��5Q+93�X�-�E���s�W�"�7�B�c,�5zo�r�g-ap ������3Ll�u�Z�r�"&���w��JٽA;B��6�ۍb���r,�}����wce3�ruq݀
����h����t��()����Q��Z��ч�$��Vb�|���b0��"�`d���fg�yK���2�,Y�æ����煩������dH�I�e7��U����ETF�����$;����U����Id����h-�3r�j�Ȇ����2�'0&LR܋wuI.�T�����ӡ:=L�w��4�aϘ�)��Dt��d�H����<��@#��{E�����$)�L�i<Z�:��X�\����2gG\�c�>��:��b�1�V��'+�@L�LZ݆Z��ݒ�yQ���!d,j���I뗖(���4md��{KAۼv�����y	'�˂eVk�!,�;'>�y����gȉ�r8Z��~��*[�]�=Յ�N��!v�~�>`�)��袥�=�1�;P�}�v|YZ�7M�x+iR>vWg*�a�Ӟ!f\����N<]�]��֡Y1�A�f	B�d{�G��ԡ��W�u9�G|���X��8�9%71H���*A~�rr��hU��ݍ�����Ʀ\9|�=�3��Q�w��%�:dl�]D��Cu{n^]΄vø�L�g��.dnܨ+�0�s���6kc'��r�Ýe�������d4�K��F�����3��
5��x��n��3�S1� h�yVǨ��>r�_h�����,Hk�(Q�%{q��u�B���y�5Ď�pu��]t�zp����X͛�Ǣg�]n��յ(��_#��s��כ��)�Z�;6���N}.h��/|���fl'�r�aeS��|6nN�=HUƀ�&tJ�횐L��cW�aG㔲+�ʬ1��> Yk�&��(�E��H;1�ifR�gb/1�ҷ�n��V��$�vK6ɉD���`�����ȪÄ,�
#z���g����B�a�͹r�l��W|XI�3b(v�M����m`������!�1\5��C��6YM��4E�i��(�?����SQ�;�ڦu͚��������6�#ۘ�L� �&mor�:���Rt��3�n��z.�k�;�dy�1+ޕ�U朣2t�c�qҳkTlty��$Sׅ�q���,M��D6N8��V1���
�P�U0�+��kd;�h��6��C��ܺ��k/�{�^<��h^��vڬmNoIon�D�e�&�87��s+�-|ᗍf���YY�Ph��7W�Yb����������1������u"�7��vÄ�a����ʼ�ʂs�,[E�<�ћ��u�0jw�v��J�Kh��3���q����X@�����bٺ�u��?�v��9*�K,�wXR���ұ�RjD���cW��6�:����|ol���F�n�-QƯ��HJ����5�.+g9�S$N��-٘��h��y��\�Au�s�`�Z��f����K���y��,��~'��AK�_'��ӛ��d�5��J�໣�e>�^�KhlB��q�^)��#�H��N��D��T�r�m�X�v7^����־���IөvIy��*����ѿ=Ux�:wF�̼:]�o,ɬ)a�2��#������9/:+�Φ�[]F��M�aە|m���Ax�G�2g2��Kz��RYj=��d1�7f�ue�)�T��QR���0ӕ���aǌ�J':C�Gշ��3eׅ�4"f���_wwQ�!G�M�My_E�H�Fv���R�M�>j�,�[ª�+����}/��Fe�yϬ�yB�_>]J���%1m��oc^^���U�ל�>��=-�37�S�3�j�E��13�KbD��UQ"��z}[J��XU���䜒�����%�%*�KLki�T����ή�U�ZY�3��C:*%�]��Ds/��e�VƢ�R�A��;2����;Ҫ��س^�v�>FR��v��of�B>y�|��Jt�r�����\��W�D6�Z��P���)�ޑ���`W��}�g(�ؕ�����ќ�Z��KN��l���w8��2�,'*\���r��ѹ��W���+
>1g��t9�F�i�1��gb�I�e�c �9��w�$���q6}��ă=/��z��]�y�x�O%�xec���Z�C�z
��y��*r�v2�:������_$Ue��6o38"�k�4��x�p
��do�T��L�+Tf�ZH)q]�����c��Am�������n�� �#y�4��J2h�b�*�ݕ9�AJ��a^f��6�����,UԦ��xK�RLn��o]٣�#��>�[�6�d��.]�j4�5V��L�)k8�2����(�%_����h�1{'۵�-��,ۖ�D��)�ڪAb��]�\��n[6�Zz�� f잒�� �&y�#��E_����Ճ2k��-'[�!�W�TX&誢\f�8H�q��N�7��պ�S��.���b�j��L��K&�.�2�m�h�;��]�8�nj�;�k�P3Z���к�3i�Mc�8-d���2�k6�δ�4RC���d87�'c��ۉN��n!�m�ʱ*�y�6�m�7���;�Jp�Thb�h[+�woω/;)V:�ee�����	���l;�Gj�d���κ�	VS|H{w3�]�lz8�x#�xqSR������D�K�h��ڲ!-@Ǿ�B�x�Y��.�b0��Z��N��b*;u�1���L(�Rvג��Pͭ�]j���W$-E���������˜��}be�J��cW�=�m똲�{��EJ�u��]� ����u;q6y�;�K��Ht.vbEN�;#�X.�n�U��z�8��=�Q \�\>�Fj��� sF�����F��_���T6��]j����\	�t��-���]sE�++�N9����W�9��uL�ހ�^N^���哦����[�Ubf:���R2���Y�j�i�K�f8^u9K9D-��5��}�y�.�f��2�M,�w���v��CQًN1�9F72�#:���:���$�>V�cGF��N~zK���ݥ�9�� �0;�/�����ʢ$�%��h���):7�����84����q%��� �g6�˻�ﳂ���C69�.:�;3.�����'v3�uzPΉ6sK<�^l���D߫4�\7�/3U�B�<]�� G3���������T��g�g:f�vb7{����s�Hǫ��ȹ�1�kM�=�D�Q��?G�NHC��*?Fw:Dȭ��曊�m��W�-���������b�"
����XQ�]P�sz�����M����s�g���L�`l�F����8���=%h.�L��P��{�.`94� y ���	F8�x�AV$��Qˍ%���������ċQӷ*alX��6$l��X�B��+y�ۅyk9ʝ��R�sPc0�8�)�Y� ���u��m�T3#��yj�M�ݥj�ڪ,2[u��L�uw\�yt9�f�� X�f��ƣɋ�F� A���㈘N���M;�$�c�E�M�9z��k	m����{��<����7���`�(�sO<�{�t�+�R�+�ϼ�k|��(���z7�|�m)�ٯx[7�N�ϲ���>4��cɇ�}g�kr��:�v	#O��82n��9z]����lt�j��nF���U�P�b"$9[���4L�APAZ0�t�� :�F�y�F�1V�B0�˕�C4�ӹ����I��������^^��o�yIrx��ub��zp:��N�5�<:�\������:oŽ��o�� v��������;Ӣ˸cp��٣�-e�8�lh�6�cQ�5�i�~��ys��b��ͦ��q��@<��=�\FS�[�rh�H,<%G�0��|�#�0��$L�W�X��fl`h�]�Q�[}�W��p$���7q�}[���H������¶��m�uK٥��#�A��K��/t��)[����
�08���>$.�D��cg=V��]�؉.+\��	wI4�Y��.���j��Is���Ӊ\��L��(]�8Z�+t������{�宇U�|E�g"��8���Du;pjԾ]�y�ɷ"]3���9���s�N�}�]���ۧn�bp���e�U�s�W%��9fG'S�W���پ�i�܇z�_:��W�ṱ�4z��X�v)���&3���|��T�$x0c�.4�N��N����{�#'�aXA.j�s[s�� ��E�-�7Q׷;��Jp�I��}q0 ���b/on.�0w���^�c}�籨�x
.�U�Źf��=�3���qw�Snr����| Fq�H��|�n��Եwz�b�/t���;�p�ȣnGzO&Л�]����5zHzGf�S��[�v�1C�#�(�N�j0d���cTZ��H��G����p��9�J�iTZ���E������l$�[�)�{e*�x0C�d*j'@�;�sV�n�Uں��nSAD���!��^sٯTeD����Xi�>y��/b]�b������2��Ud-܍�YS����.d������1ߔ�Sg���g�閭������q���#�)��,�M���k/��%�ۍV2�`�5�>��v�[3\�+���lWY���Qw�jׯ���no�������aN����O�t�"%���J#,��e�pl�nn�0��% j�8��Tq���RK��x8����dI�F�_0��N�IY� lZZ 
�ܞ�Pؾ�Q20wqn�������
����J+�Og2����v�&PS9�K_g�D�u�b�P�"K**uĪ���.ė{�F�7�5Q�	��*S*z̞4*O7ۖ�F�����$��۔��sQA�+��a��N�^^�z�\:�.��u�6$��5̀#�0�9��E^5��2�"���^K�o�w�4���˪1̻�F� A���<�9S]ux�u�����6���^	�� �E��ӻ�*_9Ԃ��f(��^E`\{S���M��MaIQ���Ź�Þ9:�r3�	��xf�C��͕�u2�ʐCZÌ�'�R���;fگp����,�̝ܱa@���Kї�p�\v���@��r�����z��c���5a�
�1,8�&皣oX��㑶d)��b&�@��gu�&�K�Q��	������n�Mr�g�Jr�8-���%DX��:5��;@�|mq1���4a��uE���wŌ�cV4Z�+�����yW��НC]���W�����=�[a�F�͝gp��_:�}��~��~B?��$�Ҋ�II$���(
KU��?�'A�?��{�%�X�f۬���5�a�?��/��!AAaQ@��P*�� �?���屢�0�L�JI�
�a��|P�!�7�S�BL%-z���D@PC� ��s5�O���������@>�`��<Т��������A��h?�oN�D5��o���*�e礭.�iC,X=��kn�(!������-��Z�,J�� ���]""�C���%-��>��e�!>
�����?�醏���o�Ad���������������@PCa�����>��Ȑ��
X6�Q�)�����&�F�|à�,Bq�(�h�_��ҫ�ʰ1��_h}c�B����l�!�ZOă�l(
CgՂ��1�U�B��_$!qQD��"�%��lP`>
5����7��e����σ���%ș#$�G��~(|��y�������P�U��������R�����\ �<`�!�O�V���3�����>_xƐAA~#K�C��O���C����$>�����G�C����
R�J����~������d���
�>�����[�_����?�4}g�
x�����'>�������`vl0���@{�?vТ5B_� B��A�?��B	���>�S%	�,�������A�J>F�H��XQ�d�Ё"@��,؟]�M�ɓJ���\�>��\�÷�P��T�4�	�����Zrm�N:.m�I���T8�G�}��?q�O��b (!.��z?���g��������!�w�����>���a����g��K�~�W��{���	�m��֥����M����"�A����>��>j$!'�QH���h�I�QA
_���m����C���������]���c�'����5�6��,�?��r�`m?]�|�?Oޯ�~|��� ~����>?O�7d����>W �e���#�#��>�����|����d?v��}A��|���H�lJ |��_M��P���τ��b�(!��b�ȱ�����C�D�S�?��>�>���(���1UAS�/�~#�H:��2���C����v�1�~�C�eO�$a(~ć����|�����]��BCa�@