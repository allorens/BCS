BZh91AY&SY�)4Lٳ߀@q���b� ����bF�|      �����dPلMEm� �-�VV�4�A@*�h*�2��6mi����[j� ٥*$��V��he+6ֳj�lvc����M�J�,mm��R�M5�ml�604�]�R���!mZ$m��՘��5m��lj�6���V��lj�0&��M���<��1j�:�h�J���s���Pd-�նa����ҭkY�6֚�mYl[+M�(�-��d�m�m����M��3��M0++Ms�\�B%) <   ;,�Ut�]+�J��Ӡӡ�u^�[nְn�dR%n�;=��յSP�k{��QG�mTmհ�`=uI�Z�k�=�jԶ��l�JU�#|2  �ϧ�JiJ�=�޷�*T�V���I
Y����V��R���z�$�mv۞�x�����-��eK<����!O]���U%DR�G��hhԭ����IL�l!YfŌL�-�O�  ,��Wգ�B��Z��
���p����v�S�z��Y+ݨt7�7�}T�����Ǽ%B�zug�q��v�=����h�s���[J�M�o<޼�Ql�S�^Ͱ�Z2ɲ�1��5���  ��}JU��Ӎ|{�ER��{��{T��;����*��Oy�t�R�w����
V������cMb��(Q�*��]�ٵ�l)�<���_Fا��\ڪ��KlѶ��P�   ����ƥ	R�����@+�K�*َ��K���kJ����R�s�ڥ+������6U-����U)
]m�i���@�/Y��Z��k;Ы�)(kU-kZ*!Yo�  ��7٣��^<X�V����yU&�Ke��W�U&�����V��m��޽cm��m�<�]䪕;;���HJ�o^מZ����=y��n��V��Ԣ��޻�"��fʊ �  ruo�iձ'�z�=)
���RU{j�{�w���5V�ޖW���n��U�-��@=ޕ��4�s{^ 6���� ��"�U�Mm�2��+CT��  }���� � Sۥ�  wA�@��{z��s���:P
ۧ�� :�� �W��@j�^��kMQ��vS�h5�e|( Ύ���{pP����t�c�	�ˀ�3� �����W:�=��[�-��wh������l�Q�mc	L��(  ��)�,���`v�%` ��{�i��t�� jt�t �{�  ��{� )g�w���47�ۀ�o�    �   j`�J��  � L "�Ѧ)JRP0i��	�0L�)�)*��hz�ɠ    ��$�J      �A0�*3IzF� �  %$�%F�)�M54z���jD���>��RC�tˡ�}��}�����jɺ{ّf��{ޣ7W�I�πff`�ߝT U�EPT��
������TUE0�	�=�_����?�������UW�pEU��J��AT}��?g�?[	�L0��̎e3	���09�09��e3!�L�fC0L9��&e3!�L�f2��c0���&a3fa3	�L�fC10���&a3	��f0��a̦a3	��fS2��̆e��&e3	�L�f0���`�3	�L�f2��̆d3	�2	�L�f0��̆a3)�C0���&a3!�L�f0��as!��f0�̆`3$�d3��fC2�̆a3!��!2�̆`3	�L�fC0�g0��̙�̆`3!��fC2�4�fC2��`A̪��2��D��@s eI�S0��ʃ�Ps
�`�9�G2(L��s e̪��S2�fȃ� s"aBaW2�f�)�Ps
d̢��S2�se� 9�0�� ��� s d	�2 ��� s e̠9�2��L�L�9�G2��P\��fA2"�P\������2��A\ȋ�Qs 3*�`E̊9�G2��@\�#�Ds�e	�G0��A�#�s .aQ̈`D� L d@3.a 3�As
.a��@d̂��2��\��f̢�*�e�*��S0
f2�̙�d3!��fC0���&ĕd3L�d3��fC2�̆d3&`�L�fC2�̆d3)���3�L�f2�̆e3	�L��f2��&a3!��f0L9�̦a3!�L�fS2�g2��̦d3	��f0��0L&d3�L�fC0��̆d3�a3!�L�fE1��?ł-S_�4?��@&�e���^c�{�����Q[�(\ؑ0�G��n������֪|�ȗ#�+���)�tPs)3+2��X��KMY��:�*�*�T٢@w��Hܵ��B��#�y=M}��d����k�C�z��Wz̖��/�뻝������j�W�\��o��d2gZ��nυ���0.0r��^:NX��������ب�w���%"�8����K�zF�F�ķHP�7��7Dk�f�n�ז�N���XK،R?���8���έ�2RvK�Nl'�uT`��ː�D.S�I���θ��u��rvS9f�ӨP�ci���!4V����\���|�p4��v(��+��<\#�����I^o.H�U��o9���5�#s�t���a�cF(zT�������n��:�.�k��=���H^]ڶL�vO�Q���޳ZVK���k,��za��{�)P��:�����E�Q�#�vł�{�Pv�R�S<�9,驆�9"l77��X��y2jWA���z���fn5������alB�m^mX�8R�/28������Ȏ�{������@R��wj��X������:��'ӎ��܇���`s�Ls8��ޝ.��*J�M�����79�Kq�ꦪ��w���Y�f�����h?,�,���q}������}�P`Άъ��⮌\�+ f[ڱ�qkkm��e`��|��D�z%��{s7I3��gv�C{t�^�p�k{������,W��� gL��`Pn,wn�W��=�׈0x�Ԋ�ɯh/e�h�s)̓��bnI+���D�u34m��m,1�Q ��[�]컏8�ḦM;2��Wh<ာGn�~��hU��>��,�fN�(.S6r��V�μM�Uߎ��)���@���S����ڜ[Tn�]P��0�kph�J��N�U�-�y���iS�Gpg`���J�av=�V�H|�����N�N��'��
��^Yݛ�2�v1UV4��T؞[}`��2�xl#�V�;�����f����kVtL��O�����ۋ�}���4b�����J�˲MՆ-ạ	ѧ(�ӷ!�,gaۼ�J��50�iC��s�Hs�^��\&���b��+�2�J�ק�wד�gv	X�5���f�f�����ֶ�V�Xc�
����V��@��ÁV5��n����iz��dԽ�M#4ۯ7��ï.���/K��ϵgF�3F����D�IF�f􉱜��<�Ku�a��ƤD�VnB�SB�y|��ռkiv��]=Ō�z��8�T������b�Z�-2ĕkZ�˻v�e��t	㧧cNk˼s9�FW�Q�I&��z2��pq<eـ�r'��z�0�'} {��Rs.���5x�5�5��!z�z=�P��3j�)��a����Ř�=�h/�/	F4�b���B*������A�L76�֖�l��]3�P��j���,J���pM�LV��_�U�ò*v�跞��>}u.��x�!{{�w�覜�����h;- �i���;��ی�����>�sLզ�@�Q��:���3�٩p\�b;���I�^�Lܽ�K������\�z�]KB�î#�R����o�k�%I�LIYx�^�6�>c��1���ˉ�vj��לf�+8�q��K�I;�k�<�j,o@�3�T<Śf\����:���p�������1|�>H�S�����m��4����\&k�֗.�؊��7�ٗ�����	~�+�NǛ��'��YY�&�*1�����9}NDL�}OU���5vts�DovK8��H ���Z��ܻ�:;��΍Y�S���e"���,"2��l;M���=��mwn�1�5l�7Z��P����;k�� �+�y%b�:��f�ڢ��0�M�4��^�����y��Ra	.e�+����-0d�;ҙQNH����V��e%g6�����s[P��5�ʶ4�o	@�aQmV�h�wX$��5�e�w���nڳ���e�q߫,�U��oB���^�)�����6r>H�].Ԛ'&>��)���}�Pz��GsY�I:\��{g%�Y�������~u�S<=(���6x'�-ܢ��C��	�-L��3P!/NB�'x��)����g���+�]F��YJ�h���m��N鳣V�g8r5����Y���ayf�|#��jN�����;NΙ�ƙrޔ�sZ���ͽ@���wKw�N�Ko.�v����^�9���o78�8�YzU=�S�X�j�\�1 7��ɛ�6���e(�RCt�E�t�	Ű�&�9��5��y����\9E�ZWf�S+];�R��ća��?�ɹ�`�l��*�׃{��w7�h�a;xRM.q5��]�ʑ@l�ϐ,eaxȼ���������hV�V�]��9�+Ԍ1�}��5��t��|��J�>�u��[G����Qպ��n�;:�5_��Ҿ\�>��ԝ`��^�&�˄�
^�|k����ܼs��/��Y�9��A"�þct*O�)�p��/N+�f��2�UZu��p�k諘�m8�ĳ-�u�C���JM�$�`�fV+�K��UƸ������`2�H{6��qk|G�Q�*�ąq7��E�@w�\�F\�.�ER�2k\%&D#޹7��=3PP ��G@�R.�A�֮��f��u��򳵹bjq=�MW���JK7z�Yh66�ŭu��[�����܄\6�܏������tX;�T�љ;N�fjܘ%��C&���D=�x����b���y��_sG�!�^��q@��d%a:�(^Y���I��]Ö�ZRy�٘�+\`�4��%����/M#�t�1}P����[k{F�����F�ݜq�����~�o�;��Ѡ�9��!�ݶ�b,�p�+��h������:Ӗ}�{�d+]�!!��\�܇/�~LIm��w�aJ�H��(��'c+	�Ƶ���j˝�b0�4rk&n'�o��-V�ǰ��U�i�rwM��Y�^�wi9�X�1��ߢ����}Kv�@�z���ν���vmܲ����l����[�|�OBB�os���	�(��N٫7��r1���~��e���Vd��G7eJ��q��v�%P�>2>z�p�a�"&�u�fս5�@���kތSI&S3�Z����^���Q��Zɖ=�6ɡ	��U�QuFsl�tظ�;c��#�9<,Vgn��Cl��w�ԦEqԃh�*���"o��9�A�U)���Ŧ�=��g80
�ِe��(��5���2���·W5k��;
���-/�TU5�t�������v5��wq��*x愵��ѯ9ŗ���^��e/�����-���XA�jnb�{�q�j5Nix *�i��(7��޸�	�T�e-hӬ�X�^^1j�	Mo����f�C�'4��K�D{�/�]�\�����)[Q��0�ᑱ��*X�ܵ������+�ݛv�df�Ю�YYr���c�3c"nR[�[n-���Bu}B9�8e��u��ee����0hT�LYi
�bqv4l�!�z��A�8D`���]6q�YvC����'�[�����4����"�ה�B��_U��[���D�f�W�(��a���:�(�-���wŞ)[�X���Ykmr�]+��z�ԴEMxɺw�4�v�nag6<�M{�Ù#��gY�w�L��3sn�iD~��َ��u6�c�t�J���eƇ����aK66q`�XWQ�x+nJ�Q���M:�j��:%=s�ha�RZ��Wa�eZ��8h�$�9�ս\���W%e�s��^N*d�ݦ�w�n����9�Bł���uU�7q�F,'-^��ynBbp��Z	=R�e���-���i�.��������5�n��x���3\;A���U0F�;��G&�Тl�J�/M|�W�t���=���bذp{OGѸ̅��{^jf����(��u���w�MiZ�r[�0NaL'��ۣ�biCY�h��m.ةP�m/;�͢�p���4�'#�FN���ڰ�N;�tb�r�)+��;.�_;�_+M}�V�(���(�J|&�XycciH1E��[�Z�~Q�b�������a��PW��iH3�#��׻��gS5���>a.h��z��;����ݡMA��̀�a�b}�N��t�N�{��ZI�go0�r��3�����N+Sy�sܙ"�pP��v0��fi4��vbZ���Q�[��{§�v;�so\����a�m���.�L��(���[Fk+�U5d"5�wn�܎ ����]�u5�9D�\�NNY�l��o;�[z�j����c.����]�[ԋ�y���ٜ��)S�T}���%��w�բ�`�,���߻��4���(fˡz{T޲􈖌��ƃD�̗y�:.����C2�&u�����s�c�)s���z�Ë������aX���$�����f�!�����.��[���s�O
�9���z&A�Y+�Kc���J�'}Ch�ش����ӗd����ḷ���jv��%ûU�8Q�-S:^�;nt.�ޗ�%�G)�$f7�l8�_!F���_q���=���l�v�ıUr�7��:S����aT|5q�x�kco�`��l7��O�ǎRva���kc��u�a�^�(10yoo%v;c��E �"�e+�E"�sbVf.JJ�/�����Gµ޹��-�T��7�D���(s����N�*t�7�����v�Ji�O�<&����JNE�U�8�z�-�:�0p�a�v�8���~r�V��́�F����4c�A"�X��dc\����6q䦂�ŘYŶð���1g3o�0�`���ԸF�r\�iw:ض��Z�AV`ޭM�H������.tJѪ�!�۔��
`(����"�7�˪$Hf�ȨVd�T�	�t
U`\]×Gc�2�Do�;FP��`QQj��h]��9Q�
����AY�J�ք��1������jc!<n��
�L-Ƕ�e��m��u���Z�^M��������l�tz,�rO�����ʛ��{�
�q����Q�xZ�a���$5e?d�aL�󛣓B$�up>�N���!f���7WE��mx��k�����2��/h��x�ݶTi�����$[!�����T3��#쭸ݻ:�����Mm�h�U�v��;�%
�Vpf�	эcD[�7�Z�mk��~�'G"�g
��fQ�+i��W�Y�R�R����%��U�Sх�&EJ��� �n��D�891t;7���u�z�d'��b�3mȆ�6��AG3^�M��^�C��pYhe�E`R1��`��4M�[�y\�ޔށ˸X�sw�]�[;�okN�b�ҵY�[�d4���4k�e�l�@�u͜���lkDk�7��Ǡ�GL��Q�y��ov�r���~�8��jy]OL�O�2-��֜6p�Ӵ���0*w"�����&`0=�u�Z�n����gr5/"�h���ymK�Sj��*Z���e��m� r�q�F��e60�-Z���m]d.F���Su]�����6PM�3$NcܬcL���v�Y�l��RN.Zz��[�tAw�`m���g��F��oS�ԍ����RjS�{Jg[l�#{V���,C>���]�KIg�{X����7q�w���^�3��4�\h�U�ɍ�o=��w��,M9n��-��sB�o��m,�-<W�T��8Z���	�A���g,�_h#W]ٴ����,�l��rN�SȲ:��/�9�,=�X�-B�̛��بh���CH�0X5oI�D><���J-�|
���:�9�l�VV�]����.
��j��-�t�	u��X��^�\���n4���[��kB�Z���r��9�Hl[��n��,�N���6-�k2��.��F$:>����:I��N��WT�9z�m����I�4G{�L/$/g�pgG���=G�As��BIx��*�_n��C8�!�� ���;
��o��V��Pr�Ģ6{M@��+Q�.�#v�Q��|���vJ�'uƊf�e�G.Sc����j�lG[@�e�&T�V�v�Ǻv�ʡXU�ūsp⽷��m[�Y���B�Kk!wdb�*mֆ")�9N|k�զ�F9�mPn�vr��w��㆛��� j7��a�ڴ
'c[��%T��E����䒻Č��g��X�[��Z/L�6��ѡ����%-6�H��S�q-Zā��i�����_d�����tߴ���$<�=7F�]b"0a���U-+�j{v�<e)�a��[�Y�iE"B�y>��X��v����V�񎳌eY@4�@ȋ��%���]���`D���[ٹ�+�ح$��m|8����(f�^3,i%@���:����(�~��h�]��D��oY�7��� ���Ta�&�`�+�u�X�ǚL������_�}�+=9�f=�`�QԵ� ��z�&p/�u�7�����HEZd�8�d\���N&�k,���aI��#Ik�g����{q_9C���	��vex�X-��S�kYM�&q���NJ���;����)�%�eV���-;~K���;ID�ؒ�O����/���y�:��Ot	C�2q�}�X����*{��Ɍ�N��+8#��&�wi�}���2�K�J���!:F 3i��T���}�␤�ȨX���������Ž� ����~ja�ɋ����=�o��sy��0�MꚊ[oe�Úe6��*n���i����I��N}�|�{��#�96՛�y��3�=�pN���,��1��p�9l>^G�dR����1i�'W�bjǆ��5jS&1�e���S�o s9L���w�{�~�ں�����<��>F|�}�퐗檼�xk����q�3e]��Kjsu���*�]�oB�&����f���ie|�g��!轗[B<���z�3'ӆ�*�E�Gu*��#92�}�<�t����M��/��E}Οcᱍ��1��_�'ה�9���q��Nr఼���G��g��&��X1J(l�*�ڴ����+��3������S:L��,��tvo*áe���v��]i�Ϭ�bLT9lthV�2�O{7E���j���E����R���<�E\�Ko�tF�V:N=��f����>�̙(%o�����6�ղ��}�{�/+��}2�wq<�W��X@�7ZՇ)��L�Iu�gW65�n�r�]p��'4�ǟ�����IE����z֙�����(�'[d��Yzq�J_�o7�9�k79׮3���j��آ�θor���.�|���ץvB=�97�7�^�T�+5̅.+�2����U��96�Y(,aT������J�`�D��%O�����%�q>�ٕʐz�8E�x���Fzf��.,��Dj��.j�_���%w,�2������Cu[����(�u�q�af����� �-v��y�'��S}ٮO[�9��	;zx�Q�����\;<�����)�w{jc�R��]��i�����{����ǧt��_/R��,Y�=��ؑ��]�8ɴT��}�V�ɕrڤ�@��v�;�k�U�ZM�K�0�/�2�V�1�+�M�}c(�ac	��+7��4�ڸz�i��o��pd4�>N�R�Z��Ϸ���e��uME�n:Q�ue��=�@g�gR�*���-�.A3L2��0��V+��雫A�]��W�x���i$p_�ȅl�q�;}��.Fޘ�_yTM�x��~sf��
�P���ؽ��gwzYW�i-OA��v��I8Ų77Yiȝ͆�+����B�,|�`-��"Z�5r�S{Nt�ѓ'V�ȫ$o3���q��J�{nc�ŵӬ]�I򢁽�βC��9'k��jL��*ko�z�\�IB�kϷb�i�B	Y]��*YN+�ڬ�GB��Ԑ�H�].s֎aĪ^�Jްh�����JY���u�4����N�/�%�oU��t��>+�0��U�����Q���;��6A�7��ݲv�2�_�x�u��w����d�� h>̗sq���4,�ޮ.(^'.]HN��f�v\�X��ڮB�0�#�RԻ�h�݇�K��6��_$�+�^������j�f�?/��l�Մ�����ڝ\�n��+�%�7��92�ה��ҳ�Z\�_[_�<���n����qE�������4U����ם�P���gG�t�y|�o�	��aE�j�䅟zTWGt,)a���dk�<{�1h����bo]ޭ���ό����r���{V����q��C�Z�uÓ������{U	��N��\���L2�W���r�Ǎ&Ԗ����
�Pp��;���9k4�Tm3
B�هdY3_C�z�է'R˰dt�;�S21ٱz�Ut��F�d���J���8G�I��on�9� �Ǌ�S��}4D��y��ˋ�O@%uG6���DC�u�3ni\�.���!��.�{5��+f��`����M��W�i}�k��  ;2n-�i�´�����?���z��Wp>K��%�+Ө�1���}�{�ڼ}I�X����4������Z��#���
�d���8�Y:wy����S��7����۽a��=e��A��p؈�؄���}�9��J3���V��s�y[ǩw h�V�	�Gi��pa�����b�,��W�^I��ZwXe���3km8��Q@v��G^n�N�����ö����R�/�/!��������&�x���}���5��u�z �O��6�}7��5�]����^��	�S�P�;y��庛���M5���Ԧ��mҨ�^<�pK'N�BM�%�X�__iA闵��xȴ!��6[�7��gD7�=9�*�پ=N������q*8�2� ���ti:�َ�αR�Ά���g?�Q�*&��E
֏<�}X֠����)ϧ\G����w�{��H��u�^`����l\����09�J�3�k���r��U��89���j���A���7��(�/U�@:kv�ȩF�ؚkyu'��=�"4%����^Z���d״�.��&����_u�z��BbJ�K�b�X�5��Iuiy��7������Gd���1P
���Px�������I���������t,�ܲ��f��5W�x��n�9l�u��#��>S�믾ܑ���󰱝����U}C�j?^w^���=M#!����kў}��c۴�Ӄ~c�n�_(�\�R�Of�3�yB|���}�eV��z�=7�ps�mA��C�ؼn��Y�ݯ͑�kc/͕菒�,���Mq�Y�a��l�R�AP�I��ьjЉ �h���{`�n��D(����=�6�E�������u�	�p�)@in�����ѥ^��֥���@ׄ͗���պ���xw]��!7��' �t�.��\�B۾����[1F���ڗ���e$�#�ye��5�u�� �t���������*=mtSZ�q�偩Ӊw�;�|zD�\�j���.պ��=��13x�I>qA7Ď��������C����v��=��4_Rf%�mi}������L���N����
�i���K�^A�u��7�t��uG
I�'c^d'�u:|O$����ᛚ�.V��_y_eޘ}�`�-뢯���{�����.��3��ΐޫx���R�̃�񗬽�הd����!˾�^�9�i\�ޘ�ڰ��!+�SE��og�Gq%a1�j�K])\�R�1��r�:�\h�����I�r�:�-�}���tr���e��m�5�2X{4$_�`:=JQs�� >=uט �q8^�`#؂+��V�^Gbէ�T���%��s�%�V�S*�o_rZ�7b��xɒ�nR����VW���n�V���%�ym7{<x^�"�J�[d!�Ra�ب>�sru�a�Mm��"+z]�:��ǰga��=����Y�@GN:5H�ɺ�=}�%f��/Zw���YF��_(����ɻ�Ϥ���x�����-�O�	\��Ӳ�W1�!g���0�蚓�jX�Xf���.���Vd�e���w�0:9�3q�W6W���ӹ�bW�G�?Z�\ժ�'�D�L���d��v���0r�I5�b�F��ps�9c-H�U��-e�a��ǱM�t�fd{DI�x��T{&��|�N��+/cX�䝩ß y��y�|z8�L_|<�$=�F�y���_T���Ե��Ch6���2�]Gsp��v�Rn�p�Ue[=���$�d4�F�=��)�g�`T��:�#���fɴ�Ǟ����t��~כ'����[�bO�_L2���N0����/�Fص�7���R�s3%u#QXpBj���eq�|�4�%sWT(:���(�M��b����ђŏo%8�{RA*wf�`*�h���^��h��+�ax�t�7l�5� ��+7h��ղ���9j�B3�+y͟ePioqb�c�r���K��_�,�e��h1�f5e�\��MP睽����+�MY1ܛ�y�)/��LIp����T"�ƬT�^]J��Jb���1��l��vƌ��,�5�K��w����5Ua���U�1&	�m�Mc�u�oS�R�A�l�0���*�M����ƻކC��/�k���C��߲�:ڔ�5��yۭ<�瑝�L|>WD��)�3���������b�wn.؁��S��Tv�� <�j��?���
�����Z;t��59�y�8�錜��nPW�U��k7NeiD��v����$��L��d\���/tpL���������� ���.�*�gG7+�'ub0dXOD�j�@Ȫ��N�[��K.����; ���i؈̖0=��T@�������v�����އS�À�����BS��*�M&�(2"Ws�v�w��G1����x;�S�F�$"��?1�_��?ggw���K4�Z☝�������.{��L7�Wv�Uo�)Htkk��3!w{	�Wq�ܚ����g8	6��h�fV���v�p�%D��C�D�˝���M̷ًJ:�-?;�ַ�Z��^���iN;3˲'/aF�ou;��EAo���ofە�2�a��TDh{u߻�V_�+6���N^��v�5E��e��OƦ�RQ@�m��`��XdjS��@�7k���E�8�s�h�q=���a���v�^'�-�)����j���]�v��ZVt��cͻ�j=��0�^
�xv}�q�-v�����x����Up�x�Ǯ��px2��,���pҫjf��jT�tr��t��H�E�ц���Y��w���<<��.q�k}�Ot�j�>�&Zއye�E��LQ̘�!1^��0I��._��{@٤ХU�7{,�����6/z����}�{�l���H�zŒ*ƾ|�_!�eY켫\y�n�����ٶ�8Vٗ���;�L0�g.�S��E��ǆt���\�I"��������zL�3��M�6�q�T�.��x�֜�(;��qTQ���sl�EIMs]�1���u�%�9�L�vn�& ��ɽ�h�Κ�ϝ����i��}`�݂��de����|�Ls�P��&�Vی�4ZRc�|���A��@�����H�d���CA������w�D4ށ�x���ψ3*��9u�h�o0��Y9����-�c��i۲K��:��<�<$\�kCA��w�[���k���$\��%�s��x��}�H}&v`Ǒ��ÌC���������p�3ê9ؐr��8��3k쇻�ت�$6�J� ��x��v8n�w�P�!�k���s:N���R��3�B�:z�1�;��EVPs���D�^�=Rp]p{���Ŵ4�\�_ש�o�p���˫C�qn���*����v��j�3+��6T�9�YOk�������z�+�Ib6[�A�3D�=�|�'���f�S8��z�ay�q��[����!(�ve����*�K7��k�Θ�y�j�c���6n+��E���*�<|��w����o.�'��6**�b!��n[�T��.ΦNێ,�ua]�n����w7�K5,�S�au�UK�͆��t���8�6��ã���A�_�זj�������Sv���2��aQr(i�Nk��}r䝙Sl�n�����n�M��p���,��X��5�j2�����*�+o*�|�Z������u�����������͜"�w2&�f(`�δ}�5l����waz_h�sa�yY#���I�]Du\�N�D��,
_Fh)w�-�d�������;?pQ�֗�ٝu�����pR��FP�4���2���<N����V�a<��;�`�y���if��Y�����]�}�r��a��"�����]�9��n�ȳ�v�c�X�oY|ƍ�������c�*:-�hS�5�^o\~�z����u���L>�����{��Ec�.�1}N����'��R�g��*�E,�h�G緅����V�5��*bLD�wz�K�@ζ5�L��jܾY�}�����k������"�l22��[�z���"O��޴�P4�jZE�_#G}�~�ӥ�t7R���U�*n����@��7d�D�H�l̭pL.K�ݛ�b:�qy�	|F�x4Q*,��"��H��L���)�.�^؝"0S���,�ef��b!��z��R�t*3���-�{��^׾@�+�O���7�����&�o��V�#�zN|1���͍��U��>� ��i�{�v�x�r��>��ʖ9��-@pS��T����nZ���2��ɧ�<�����q�2%&⭉6l�t2Wf���rWi�J�-ۖM��Ng	I���.���;Ȱ�q8�\��	���P^v<�ZoO�+꠪6K�v�HT�R���J٪����f:�;��ד��������I�����;���tYܮU���J��VX䮖��Ǚ%��7a��@�ϕ���w��H0��uO�_���R7b]�<6L־����'���u�q���h�B,�y�P�Kq��ޓ�[�{�?w�J
�4>^+s؛�>���t8�ѽҞJ���H���<��I,M��8�R;�SX��'��I�b�!�i�OƘ����08�@��p�L�E�8�d3zK�0)"ιuu!�ȭ����6�=,�3�?�`�)����٧��g���5E��z�)�^o8��`����� �ͭyw%9'Q�<��}s��xF�Ȓ��gIaE�Y�!%���>wk�r��	,��X 4@M�U�q#l��e,S�if�Mu~�#!0���2ES���0�i���ᇝ"��Y�V' 9V���8(U��;��q��y���∢ ����_�Ҡ� }��E����S���r�"������w��}��?�%?���~=m۪?�M�N�|�2k��BL�7�ͽx��y
ۊ�r��'&[T8���k�Ңϭ(�,���֏ݰ��뷭w.5ss�Х{*�A�S�{�L\v���J��s1�R�ꉍ����O{ny�h�����[�Zя2�I�fN9��[X��:�٭��6ˤ�g5k�Ztm
�ȭ���͠�V�R��!�X��aY�#�/����CQ����!.Ų^L����~{7��`&n����u�)ǰ���׷S�Jv#��rJ �v�4�i3CS��km�m���N�c��o,"_lO;����w#���Q.�V�Kt�+0��nY�
��G���Ɵ֫2��j�oM�rƢ��/��f�V]+�˖�m8������)*�_�<���$�>�z���\����|��x�O>�H(xVL���W��)�ic�L�����j��Krn�(ػbsR�Zt�Cg��v�d�<��nn�]���9�ڎ��s 6j\�ϴB�(,g_e�O�n�Q���3Fm��!�"�#��h"(@�*7Y�Ѓ�p���^�:�Rvb�[r�\ܮ�֘`
ݽǼ0���g]�D黜z�@��9o���Rг#�"e�e7�c<��X��G�W�z;�%~|����M;���g�a�DZF���Yj�����ַ�S9k�B�}�\���)�3̓����N|'z-�u���}�_�����{����������Ƿ�||||||||}�>9��������|||x�������||||z||||||}>>>>=>>>�����������������������������������������������ɱ����������[�[�[66666667�Yˏ]��̉�.��� J��j�]G� ��5hӧA�)Z�믦a4�{&7��9����]�&&v�]�u5��^���LSKQ51��/uՒcYgy��X�=<��b�v<	�%��7��vK�,I��0U��7HG�+[Ջv+��C�35�Gh�'ff\����[Ű���P�bޝX��Ef\w+tMwt4����if;�F-�i�.kY¾�c���i�q��AA�}j�
��]X��R!{n��:^bE�;\e��ftgE'��v76�g:��q�Z'0V�1�y�m�CF�@�2��>� zy^�)h�u��L󓑮;2P�}Iu��N�LM��C��NԾ=L��B��#�����f��KV�ҋv��x�9�7v���-P���J
��q�.`�;���������t���yM>�;��n���L�q8BX���k8`V/�ȗv��Y�X3�aԜb3g���#
7�͞���x��A�� �g�T,�y��=8MR��{O���Y��>+z����Κ���a��Ő��.�����Obc`b�Y��̭�qb�C ԥ�ٚ����=��:&�̹JZ.��:d�@�KAm�9�Y}1��].�T�M͂���zj�^Cң7]�,_���ijklklglllllhlll��-������������o������������>>>>>>>>>>>�������������s���||||}�>3���������������������Ϗ���������cccccccc��������������>>>>>>>>>=�1llllllllo662lc�1Og!�Nac�y������n�n�
C�Z3/)h2��t�۸܉�v�Y��hȟ__U��H���'V%�Ҁ���#�|�75�>^5�|a�N�>��d���ҽ���:��^I'=������<���o�L��y
ؔ������"t�^�->t�?r<zN�Jf'�1_U�z�s���d8��NR�߬��,z�%���w�1��T��s&�v�.�db!���{�Ų��}r�}��Ӡ u�z�S��See�D��0,+m(������dݽ�sk���.�-���41Ȳ�A�	�X;�ૻ��}���w*��ZE]�0�\=�܋2�J8���E�6�n�댩��
��s�����k����FB�5%Ut��ݖ{�K�ue����A��t�N#Cvz3b.+����M��9]��_�3$kr33`�i����vs��n�.Sc��k���婭��5q��!{���|:�M�q��)���{�x\�z�=0f�w����|v� �T�N2�Ҭꅧa����+<�m���s�7Ѷ+k��oQ��I�1%%"o���TFӬ��̆���vs��𪾥ٔ�wMw7�����j'��M3�f�&+�����0>+��oMcX��ܴ��\ǎ��<��K��&/��+���{���pW:ٷ:�SDƻwb�V+m�Ud�Y�-�U���jN��J�����1��%�(�.S�P;]�к�?�ѾhY{22�FZ�2�e8�=��gn#W[Fw�°��	�v����qnXZ�|-b�'�[ZM�hj�Q�D�w�K��Ek%�)����f=�س�[�s��aw����\$ǯ,���vʤ��cBP�.�ҶM�5|-~[:�'�.�/��2��7����BO�z`�B%^Ń"<��n���ͻ;��6'v[��\�e�uA�F��������X�w��C�z,f�ͮ뱜�JG�x�ib�T�)O1��g�1�sr+ɲ�&�1��>J����� �����⥩�/JO�I�o�F�/������hA�]�Y���E{P�S2v�||��:�Mu:4�U��h�StH��y�5M�Z�e�r�����0��9���|���o��啝Wb����|�<KޙA5��Fu��v�����ͪ�;����	K>��GR��:u����弝�q�$T�R���-̕oT�Q�0·+��|WHL�Dk2�V�v$�=��f�c0�-x��b�2�Y6����\��O%.����Vge��Ʋ�Hc�M�W!�Zn�����W�Ú��������B�К8��ۃ��r�C��δ�	��R�;�����FmȮX����^�s|�ttx��i��;$�,�H����:Y7X�,�\�/ui���L�z�U��vQӛpiCiՔ�^fZ�쓳BFc�?ђ��eQ89`vJ�W��c��ݠ\��O�L��d�yM�,�"z��y^T�2�3'��6��5�y����k"��_-\U�v��I7�/@Z�$��i�N�c����R�l�"�>黛��s� ��]�dĹ	Nj���D��m�J^�l��y�}_?a�m��@�#�������|R���,1�ݶ�waB�c4;o���돝յNyj~�!��>�a�6��m�lJ	�賺� �:b��@Y���md@(���n�V���2u.Pu���3j����[�������L�$�X^+ˑV&��tp��eAOt�ͭcK���Q0Y����L,��3-�i]��]^7���^�K�z�ֹ�\�I�m�9�o���[�$�;F,���)����no�7X�Z}��F[x�ĸdyъ��j��]T/K�)�`ņ�s�EHł뭲C|����V��y�@�ǖ����{x-^~�P���V�\$۽ᢲf9�m͊����V)XZ�p�Y�������tD����/ˢ�@B����¹��Y�)%
wJ��pV�2`%��PI:YL�ݍŎm/��I��c�K~���&k�ytU=�ϳ�x�_yL��2%���j9��T:�>�jfH�pk��6�ؚ
�{�Z#B��3�7P�ʼ���}�e���H������m�\k�e�l�m��Bqq0�Sn�=|�qOL��%�����v��[�:���E�X��Ŵ���Le�*8����x�]Z�K�L-
�ե��MV�ԡ�M���A�yQ��&��_��yf�87(b��'t��������S�l�w����n\.WP�6Do��������wF�QM�֕���/�*=J��'8o,r�b�M>i�dz%ưt{�D3����n�����v���d��e���7�ŧ�ۛ���7�-/��t�D��.w���YrǏh���ڱ/(e�yOv��*\��=�[�G�l���d�̅��f�dn�+����u��C	�c��:b �/��w}��/�K��&%��ޢ-�UÊ^p˶�]�"v��Bg.]���n��?�,��d�Ŏ�ɗɔ��9�]dH��㣥�t�qł�{O$I5���Ox�������@�\E둅@��AJ�D>���je>����r�x7f�|:C+�l��@q�mM�xA�.ۘTI��(�n�6��"��u�Ќ·ʲ'r<b��M�fo�FG5��J��b�� �UƄ���ܝ�Uw�gc��M��t!�c�=��yeR(ys���a,�Wt��=���k��u��y�����5ǝF�g��C� ���aZ��̮�4j��3�f�w�dF��S]���.�=�&�_w�,瑹�.�������^�W�^$M:"Z�i��@ƻ��v� **ۺ�U#7�I͂+1h���ld����R�$o6�]ry5e,��^J�i}T�c]� $e�f���K��b�Ns�����h%�)]������RZ2���el�|}�pg%��-�7#���nG-c�����-�0�x��׳hAh�{}�5�jѸv����y4m�
Ifd<���ʧ*l���A>"5�3�3�����I��� �u�8k����]�R&;���!��p�e�U��j;���"�� V^1wvF�\yg��	�*��x:^�F����kM�:�LU6������r�6���|xR�ӝaa��(եJC�dǋ�{�ݽ�^Q�'޴QUG���)b䊐ɮ�6�$k�f���1�wھ0�y��pM�{ץ��S���ŧ�}�ɇu��2a[�J��.�j��n�����+�H���U�����0���0_�xm8�����������V�ʪ�ye��1lM�'��6Z��-q�gs�7X6/ت��:@بo�Wi����&�L?ZW��S��Vu��N����jLU��r�ֶlNR1� P^է(i��)=<��t��:|�������;����K��Q�k��Vf�ttQw׮K�����J' �&��XI��m�Wti��'�۶�4}W�=&V��OK� �غy�w����ե�v��YB��:�Hf>0h�&��i�t�'g#�̝W�e��N���̹,�p�rڕ�smU���4��K��K�#�Ѹ�F�cJ�����mL��r˅+�/wQ���i�P�@i[�w[g���� wA���Щ��q��|�՘f��+M̳WP�u�D�[Va�5�w���Iv��}J= {N�s�9,�Xs�X�I�j
쵮��g�e#�dg(hQ}L_ZB*ݠ�}}w�r�����L�6a^O��W�w����<]�}A	X,���9�E��6�������[��nn3��r�j��F�Q��g;-��0�����%�`Ǎr�Z��J�����0]^�s
�7%��:C���'���D�\�+ �H����`֣j����e�}�0��J��zb9���<����W ���)�]�*��t7��+f�85�J�9/>�����®R��x�b�Ϸ�(�u��՛�x��[�����N���EX��^��z�y�D��c8�e��ǵo?zL9w�������븵V�2��q�k�1��n�G>��ۄuu7Xꒌ��� �Қ͋�=\���g,��n���ت�7�����<𕛵wx_��q��}�,^������SvUm�m��b/�@�,��K�e>P�MK����;� Y��ի�٫(�R�6A��]�������SE0bl��H�Ƚ/�k�무E�ʹ�C��K<���ܘ0�\g��1KF�����}u��,n�0�'瞆���%,�\�e�,Zt耶�a[)d���㔅��Zh4��f�R���e���F�;}��L�R<��x-_W�!�ǚ.��C|DE�5�#�̻��c.e�6���5��ά��Z�o�Rh='�C~[U���#����z��������S���﹗&��x���syi�P�to�&���nlyEJ��"�~
�U�;MqF�ZVu�AXxF�̥��J�|
�=�(sϺw���}��1����J��f�z_g��z��+��jPgq4e����p�;ہ��_-ʽҔs���e�sn
]�4�������$6e=&�������O�^�W5�[[��^Y�,��`Mm�[x4�_4��F�`��(����qEHzu2�|="�խ�>'S��ڦ_wwvf��3��6��״:���#*�\oz��t�s���c�����L�g4�y�h��W�,�[�����e����
�i�&�a��4�VNQ�:��է3m���.��9��R�CqD�}�����,q)�:�v�qO}p�|��f¶�!��{\Ӆ4��:`٫�֑��x]��ȏm�v�o�wػm�ϼ�-��}כ�x<_��f"�22��:H��j!��6,\����b�����b�c�|�^nc�{t�8h�]��VB�Ǻ�՗�yoy^̻g2�r�u�k<�f4���&0�#�g�������&�H��7.�u+�0�wgy*ӻ��Mf��;�{w]ys*;���/��P�}e������g.�x�.�
��՛�q<ƾ��ձT���vͲ�ח5Lj���2�q)�\2؝ǐ2�s�������Οr*��ˀhw��tͮ8^�'[E�3iG-jᶒ
];5BM�j��F�lf��]Ji܏�m�C���#]�[Kx(@�_#<^b�������MB^r�2G���v��ϼ���A��٨��4���Y�vd��X!n����X	�)����_ �U�|߹cd��%���c��U�ڶep�ZX��YFؠ��th�1/
�p��-)xb�)��ی�}�3��\�W�:�W�b�
����v+�o�]kKP��t���)�+�U�/j]�̯�`������Q:���U߬�'"�hLY���>����37�bG���������~P��7~a��>��9���*�B��j�8�0P22��e
�AAT�)�M6%1��!$(��
$%�fD�E�͠���!U"Aʪ�L`��R4�-�*aФ)�Ɏ@B�AIJ�q,��ܽ��U��4W��T���-�+'�<4kۙag3�o[��5WG�:{|w9�b,�D�|Yǆ���&�I�Y�G�U��^���]��lS_<��|�{Iu�x�4��l��.����[��ګR:v�SF��']�@�dww،s��Y�r��!ǎU�rc�sҺ�~�UZH�-��mޝ��}��G�^�8,=�dJX��c %�:�֓��KLin�	9V�7��&QX�z7]d�ΰH*t�]�̷5K(NA�{X��is�_ϲ��]W(�غr��c���d,:Bܳ��,�sw�?u{o�(T�^͛W#�\�$���`w�0������I��0+�fwy�4�/�xӷ���,���q5j�sGwB�WB��@Z�r�=P��Ǚ�n�]�rK&)��$s�fq�ukgE� ����m�\ճ�n�lK�\��(��|���2�y���g^����1�=�k{&Z�g�g���z �wq��ڮ���ҕ�\��5@�ܴC�c�4�uQ�'i<���Cl�L��L��{��ܙ��WR6Ե0kx�v��Vn�5qɊd��0�^�p���e��b�m���K�'"K�����Μ^�e��\���:�6�mH�t7A�5���b����Wq[��R^\�����,�jouc��bP����p" bHDE�$�D�"�E����$j~�q�
%8�~U#S)���2�!&�,�Ȇ)���	 ����\R&"(�YT��H�H�uQF��-�!�FD2D� �mE
D?΢ 6Sp�DA�mR	!DE�Ȇ$!F!a[hS-�f�N2�n@�~d?�Xt�aBhI�R����Z0��~jͤ	D3��-���Ө��V��q�&�ű���� ���b����lh�9���Z�4�O������}��o�����(|�V���QM�Z؍clMkEI�ƝU6&�j+E%iϏO��������}��oo���M��b�&bJ(�kh���8cl�cZ��EkF��X��[�R�G6y��j��6*��W��նŢ6�X��k\�͈���M�Vb��#z�
(���11&6Jڏ#s,�ލ��Z-lDZ6Ϊkb�Tmj/Q���$�.f�u��WX����Fl�(��v�Hb�\N\�1���s�1��60_v�͒ر��]�9�\���s�99�V,c����>�����j8F*(��s�r�O1�m9���	�s7r�0m�h��ns��9����:��*�s�A��c�5Z�G$�6����w9�T-�����:��N�'lhMh"ms���W:9��֣m[�Dryp��9�cFQ�:��F�-kG.g�Q\v�`�z��[c���1&63�Z �G9�p�<,[����@�$`rDˊS_�E��@�a��3�Ά��V5(I�xF�r^�tMi3/�ik�
�=Q:��5�ۮQ"�~\�;|Y��v�;l�</2�r8�$Dm�Dl��D�C��"D�����%$�`�fd4������OM� >�;%��{�T�_J��5�ަr�h���B�;�3����H�ȕs߽��O�nl�~(i&M�4�U��4�۷�'[F�F�;lq�C�����qo
)_�9Ld���+�<c�O�ד��au����WwW��/x�� ���g�VTpy������&ZHK�,G�1���E�����U9��8\x971�cգ<\����h�D���'%L`s�S����z�Of��}�b/:=���o(y�����f��ޞ�O^������g��8ײ��Zʺb�����N��Þ�zfhN�L��7�uCx�ȣ��Rwd��,+��*	����t��Di�g�ޫ�.�{Y��{���>������<���|��m~؊0l�ѫ2D���l���q��������y���z�zԺ����̃w���NZ�=}�_�[���1�I�쐶��wޗ�!�G".[��Ӣ[�"�шا��\�hç��nL��z7�JF>\*yo\����7��ٽ�f�k�8p됙�a�0��GQ,u�xrɻ}ri},�⑈���R�7�;�{n�]:�R¯NX�E[^xU�Q^�3W��֓��>��RUfR1�I�}����5�"�|[č�ܮ��5]���Rt����O�*xzPr�eH�TTo�Y��e�}S2�����t��=�E��y6�t�Q��wb��D��I6D��v��~ا��Xy�h�C��<�P��S�:r��ݛk.�2�a>7}<{E��||x����o���.�B�
T40���~�
[��r�����OԼw�қ�
�*ۢ�
�m3�Q*���lT̇�7����ߘ�z��֍ﯳ9%�{3�)���N������u1(���|.?y�]J������D��<�9�C=�t�|�o��Ć^��f�����ޤ��.�p�0y��y��'3`q�����͎'�<積����*��eY��*d7z0ߡaq��9��]�C6����űi��=x�vԬ,k��.�J:� ݠ���ĞH&r��s�m��n��D{�R���J=��,�gq�z)�����C,-�Єy��Wu^wx1��T�V֩��DT�Ծ�Vv�`6G|�C��j���I�}�-]Z���Վ�|T����5M{�[��36�\�����|��	�9[~��',��]�DJy@ymbz�s�'��2��S��^��ت��~���Gϗ��G.�v+Ԟ]7�
�/uc״$�'�4�����~Пz�{SQ�j]��Df~������1��gW���6?��st���v����W��|Ѩޣ�G�me=���}+�+�V;��f�_-�:,�B%�#�����a���M��ŅNΌ½�Q�����3�Q^��Y�mr�Ͻ�c�N\�Ϣ�5�>��+�ޝ��7��@���o=s��ǫ�����s�8M��[��_�w�׽۳�R�fخ�dA��P�MNм�	�F���f3����{����ߔy^�I_-j�߲�ݚ��\��|m`��+$�z�߯�L�f#���a��C9`J2eb���4k9��\���u�j�{L
�:��z����>�5^�Q��{����W�񦄨�bn�̻�b.{�f���*>#�~N�t�����fvvrBO7���b{��}��F]��,m�S{�RSF*��7��~������xz���n�76Y�簚����ݰ|�t���4�4pɣ=2r�Y�������Ե�u>�+<Ϗ�*�����qb��'G<�I�^3ƈ,m��{��zY%./=��>�^���C�3�E�o^3d�|���d��.-��{y���>Y�^��¥J��Ւ�Qy�.Yy=�����Mb��i
�yof���dsY#�Qkڷo.��W�U�S?>��n9������a�ۼ�O^�x\z'|ت?E�PǇ�M�}��=}�W\����N �._%'��a�y)�G%�wޙ����s3�Ux�ߙ��I����Cofz!�f7�ȩ� �='<�:��~�JxBs�<���3V��{�J�kh�t�Q�3]�������@�Óz}���7���{g(��b��q�Kc���Wg���w=&���Q����ޥ��E���D�������u�hp��Xs�7�l���i�� �Q�N�^��w5ۜ�^,�1�#ú��;y,�L���.��Ô��9b���!X�/��Ρ�xΰR��өC���t�wy���*(B�(p��^��]W>}5�2k��A����\������ޏG���ڨo��,�R�`U�S{�i�?r�Tx�E�O��Jޒ���<Tgk�rU�H�N��o�P�z�������H��z����r^�д�޾�#��׫���e\�ys~�g:�}�m�\+��a�W;ڝ;��~͛�1s��w�<A�=C�֜ڊ%�}�ۂ3u��E��Oθ�U�PW}8��[�i�^E����{|}� ��8n/Fa9W�o\y�e�9q��{�:� $Eo�;�$��h'�rhL�K_^��U��vM�ܗʹ�٫g�O�ċc������Qq1�yi����ѷ�~ǫ��|�{���MPT|��^�ګZ���s,@�p�����a���c	��;��'/ڷ�4����c�0���=�t��Ah��[
1{�<q5��
�m��W=����Y0epr���}�o����>L��Sm�bS?�������g|���2'd�����*��=����N�^�vB�uy����V�N��X�پ�pS]�9���s�i��y�:���[�=�6�\�Mn{ݞ��c���MY-3\u��Ǻ|��ݯm�������]{��㺘�^\��^{Y�mc�����7�>na�7��n�w��:�p�ۂ4Qn�`��~ރ �|����s�5�~���{����ɱy�_�5�hܟm}�v*S�B��R9�ψ~�5~{Ƶ����i��}�99WZ1��8�������c��z��Ж��g=�I��\ǵ%�ڧ3"���\���+���3��\��d�$�(=��� �l�|���p�;�g�=�W̳�*�yc]���)�=��Bb��PQ�d<_6�t�Eɾ��o��x�~xE�n�އ�sO��k��ȋZ�6����YgI�����w�'����<�C^��>��W�����:}����sS�&��{�V�0�Ƞ~��K�}���y�����{p�����`� 5&T����.�{c{�9��ߋ�	c��w��y1�}��j�
|D����u����5��'#�k�ً[��}�/zk�څ���׎Y��Z�b�ˬH���i�6ys@.X�aְp��?���ٙ
	�r��횱SA�ձ��"���	E��u�e����wz))��#.�x0��&�ת�����14�np��^�9-�ZL_c�1�vu⳻7G���x��6<��O Uy��\��kP/�f*�.�ޜ��}l
�|f�[68��}=��������Z�){��};7�v�c���!��<�댚�&y���	<�c���嘐�	����:�0�m�0���#i�����ӕ^����'�ݔ�u�?f��5]�W�����-l�Ba~+G�ȻvC]�$C�U����ff��o�a�������^=���E	1��x�L23��_��zD������C��>4mgz�8��D��P}�7����y��݋c�e��i���m*����i�E�W�Q�-�~�7� �;po=��WN��j>]�\��޻`�W7�`�::==M.'�����e�G�do̙�y�j��o��2-�&Q��	����<�ou���0�Ք;�kֹJ�KL�K���,�Z�R��W�3c��:Um5*�R��d� s-��������-�}s�SH����۝���X��[	��zr�Y��:�N\��6m=�V�X#���1)��b���R�Fe(�=ὑr�x������=겆�A^ne�S߫o��u?��+����~�y�٤Y}M?�j�&�\��f���=�'��O�v�>��]������럿#ke"�_v��Vor��7��s=\��y��d�w��ڹ4�4�6��s09�K�`��r�ō���=}�bW���$�0Ll�ؗ1�m�������CwDu��I��ʷ�y�IYEW�������I���wϵq���c����knp1y��g� �r��ק��ց�$��<Hמk"�{q�ւp6D��C�ûw����XVӝ��}Z�~瘇�Oӗ�;�}������fb������hx{�Rm���>�Yd�Ӭ�C�����7ퟛ�-�Nz��n'B�g^uH5�7���4,����v�bT�K�^p��/��|�>ܒh��,��y���vd�z�E�oUګ;L���d��(ɗ��c���%�3	f�_k���{�{pTi��u�܏��{Y�رܹ�V��3T��X#�(u���m��ؚ����3��ta�%�Q�Lٞ��/j !ti؊��U�:�&���t�{�\ݞ�#>"{�s�����˫ݳ�U:�����я���x�G|+�o��
g�!o���HNy���f��u�Ň{��p�yq�o���^W�
�b�u�?x}��}��9�x؅�
��Z���7�dd鬒_��T�J��ʼE��{���s�d�l"G*z��[��Ӟ�d�)�V��z��Fxs�_0��4�Wlw���/#7���$��9��"�(^X���Oь�>}����yN�Ƕ�]䗽�5��zDyʌ|6A6F��	�;�Ndl��c���=��������Q~�����]��s��^�m{�a���3��!��s�vt�Nf��b4��^w0Y5�>��sI=�6hٜ��6E���i��Q؀��}{Z���vߟ5�y��AZ�yd[Z�׮/�Xx�9��
&�߰�2�3����:��츭�Ѩ��2MEQ�Nt�2#��ܕ����sw3�_umH��:�F��,u#q���b�2��`�5�Q����ۉs4ϣh���D
�5�j��hs��t{G��������4��gC}���;�L�S����&l`��Ǽȋ�*��b����y���D���q^?OOm�tx疏�
��=�)ɓ��4<k4���y���h�#x�z��^�'��k�H9�����
�z�] ���{���+���3t����Ξ�fy���o�p=�e���>���U�F8w��s���z�w>���~�roG�]�P������m׹�G���s�7l�9NꐯVˣ]�]D�3�����I���3��<���K�޹���Z/�6��hkSh�t���z\�|h?z������'<�yy��3�9���~������F�(`�4�������45hl瓨�:S���f�c��7�rw�3���v�#������|�Kؾ�=��M�6>lb��V�ݽ��COp�R�}(�Ƅ�ջ�l	�f��|e;�
�Lr���O��L��L�@��]2�������!�u#��Sv̡i�k,87ۿc�d�M'�;WY�tl�er�;d	0���t�� ��HVݒ�^���D�y���Ff��<�/n;mi�vu�����凲����NJY���q�r9�����L�7p�9��ԛ�c6S�����q��w�d��e�
�=3�q�*Y����H��ë-���9��`P�n:�ř�q�?q���d���!��쒧͊'�$�����kz�:�Mԏ �S�{�j����]�x�J��F�pQ'BU�(���:�uଢ଼�7��[K���z=�0����5�:.�1H�ޮ�x��#*�d/���8�P�6Q�\9ge~�]�f�Ò;A7�k3��(U��e�oOD.����i��95i�%Вؑ^����=j��sr�E�n,�x�_$�,n���P��[��]�s���7�7�o�ɝ�T�����[���{9޷5�3NH��L�ڇc�6���͇<�}�g-�����p�*{8О8;h��qhb��ݼ�N��U�Et��b��w,<�(�&vh�Z@�z$�G_3b�'�<�i����Þ�VKڗ��xjގ��d��5­��v{��g��ލ��o�*��d�p���r���u��ڈ��۾��ۚV�[|J2�C.^9_
�x�ݏ�� ��mr����w�g`�*N�w'��Z}Kmf�� �;�*�2��eu��g�c�4��[^W>��WǺ��������.e=�9��L(cx݇s��ٗ�<�{���/<��%�u�Z{:a�C�B/�9r,b�Ƞx�(Gxm\ߺg*58���-B���>��?�u�Xvy��v��,�nZ�U�7*+8��Iw�Eh������n�H%�ut4)fT��U�j�H���ܳYmm��ɻ��܍������(���Q�1���Ր�@o���eKڲ��nu�B�
��Qf	3#�̽�Չ��*P�0--7Q�A9�V�Je�-6*�Z�D9�͙';�Yv���OYڌ��g�sP������ϗU�LIm�pk�߹.���N��H�����vl�)��|�Z0U�4b�]N�wj���G۔U	/ �����f��%`��- ^5�H�]�e�馅X��֏N�k�]�x�D��o����1��qT��d����>�{���[����cK��ݧ�8��}.�&�'/q�ڮ��]�l��w��LK�..�ܳ:9ۈ-�%:�1�Kp��fX;g>�:.��ea����Z�3/�6��M	i#Ns��]K��&�ߨ�\ͽö7 �%�������Yg��<Whi}�4��;�J���A+Z�N������{6Q���&⺕�﵁�~(�yƹ\�9��ͣ����[o�s��'5�q�lk�s�&���X(����$��5s��m���>�o�����}��o��������IE!A��)"�e��(����|��,4J�IT[ ��( [a���b9˜.F�E�<~?O������}��o����>=�V��N*����|�*�J�q�r�Ƣ ���6�A���1�1�E��U�2][�h��^W�Qup�4un��MQs/W&�m�c��g�(��4A��b�Z��6ıV�Z�L��DTu�p(������`�:32T[4b�(��E���:�]�f���:qIl���[�<��1�QQ�㘘�*����؊J�"&�����c��QR��SPsi-[}]%t�S=cUTMm�����DUMEUUIA<آ卵EUh�DZ9p"��s�*-�T����6z�9T�M0���<�Z�1I!�?H%&�6�<�y��e��orQ��mw�{x�wߞ�iDW�3�+L�N����]���q�c!��>^�Tc�?��>֧��~����ۍ싷�^˕~ޠ�#6��!�z	C�@"I�-��z�"���%�MG7���[�?_�u,�C�h:|{=�huGyLcמ�t�k�2�&�@,%t��o&��ͥf�6��eVK��#�ۮ2�)�xa����?<yK��?NT/^�*f�e5�1���s���֧��"Ob=�!����|i���"��7��Xt]�1s��UX�-����"Sn.�*J�iȷ��uX������g�{�t��0/�I�`��1������-!��]�|�{1��7qg{V���k!�� �t�-���+Ti5��=�_0�`ʅ�I��2��N(H�w��{>��k8!������ڞ��]'�)ͅ�)�Le0�#�y��.WG��t�}Z�޺۵����-<��c�1�����,.)C�2�Ӏ]�<s�"�j�a�G�ˁ4)5:�y1��h3N85�e�G����o�q�u�aR�e������-���T��dlE��F�N�!�8�5v��Uxτt��6�Q�[E��ǃy��U��Š��667S�c[7����#�6iW����Ϊ�Ou�(V��ێ+8��ι�0���m�5���K�`��h����]���_M�lEu�&�>	��4�\<"ɓ��c�v�#`���3�~�;q?s�Pe`�0�Q�X�mʺ�µ�ա�P�]�~�#��\H���D;p��1S:%��7TȜT�� ���gjS�~���ɭCٽ�� %���u<У<��=���z�3�?="x.�h��Y��C�Ҫ�J����gf��(vu����0�g����=������@��1ueЖ��<���q��h��g�w���������z� =�d�&��ę'6Y@�Vkό�X)�F�	=u���k�K�J��;x86�)��Q�	~ LL,u~��f�}}��^C��v�ŀ�c���AP�競���(5�=��yE'������j8S����7N��8��Qq43e'c���i�qY�Y�Q���z��<�y������E'�Rv�����������^��MWog���2�����\U�=��$8B��g�Z�#{b�
@����W)��� ����t�jc1�-��]�ʼ��&��v�X�M�	t ����A:��A]Z�9~��̨�sW���(��8��5�v�Z���=��|��6s���v\gX�FB���c�yN����
Jd������͑�P���^yBQ:N���*�eEn[��Xy�NƇ���;�W=�f�Ƿ2^s��{���h���8��)�.��?L�?H{F���:z�L^��S�w�(���K�w��5,�>����+�֝si6w����jݴŪ�u�/\���A�-@������#���muz����~�^������d-/�Hn���;{	�/�49��� /�ϑ�$�Z���)Ž�R��t��2��U�t�pl�:i�����p-�L-��3��n	�j�aF�:8�6�;�w��!ف*�3�-Z��86j	�M�7�"��NEv\0����`:��&h�}�u�eڰU7?59�0*�/Cd2V�f[�u�Q�]�}t a���'|�h�*���Zh9�Zr˾Z���J�j]W�&r�=P0��4�¨Z��j��F6�i�ۇ,,rt��yB�C��rt��om�^��(J�Z�W�;�zeSj�R�B��y̜��QaB�O6�4��ʥfqR
��A:���7����X���h��ǈr���Ϧ�еa̜�=+\�$�2��-�����
��x�'���2�6�z��fB��ve��Xcp�J��]5�|��r*��6{��~�̛�6P��e&�5�	���!,��a��^i����ْu�5z��N�	���)��8�FĪ�<y��gC���&fK�A���(�V].��Á�H�/A������a�_�|�|/T����YC��w�,U�ʚ$s�C��2��
�I���<�M#;�|e����!�O�@]U���#�x#�@v��h�
�s�I9;�����!2�Qgn^���gB<�˫=�ҟ��	�jKL���0k;-f���J���6b@�}�{�����L�C�.��ı���o ծ/N��E�=��{��צ���_�F�c#�yj�G=%��v�1O�\e��v()@@�X]x���N����5��H+���s�UNy})᭼��
<d.{;2�,�J�����Dc��X��B�Li�C�/���x����_h>P{^�׷`Cƹ�O��*�՗Ol*�q��C]�A�{���.�	�4�(��=�#VT����^!��R[��Le�ԛ�)a�g���ׅ]�s�絽)�R��Z�V�j�Y��ԀРc�}�YB1�/7�<u��l�/Ij���hYhy��@rN�{����{W{��Ӽ�6��UP���Y�r}�Gb���k�wA�b&:�i�����1��Z�w�}]0�0��9�Ai�cb���3�L-���Fq�j������b�:� ��L�oUxQ�4��YS��-o�9>���N�g4�-4%I�n�!��5Tg{28>��A_4��ه��v�%:�=%�P�r����Q��Q��lR�@�U���n}��W.�g�k6>���ș�݅�^����oPs�	�����	��B�PȦwF Z��������=d6���Vd��ئ7J8wWp���3�h7m� Z1p�Ne\�F�^��e�`�e���w��9vE��p~dŋzw<2���wC^�xyR
�%�8Xd���.�� <t�]�93l4q�Z�4n<n�����������U
<��ژ&�Kb�@ ��a1�}�'W��D�+:Y�����'���ڽ-y]�x�xŵ�0��a��@�p0�s���(�v���`<`~��C����8|�������u�a,��!�M���a�IR3K��j���kD43������5�5ѣs��l�Z�`��MIOr�^97�^�����7��Šh-�`j�I�(u�f�y�7{sy�r�6y.��`�P������N�ޡ͛�Y�@�������ԛ#�YJ�F^���l⇍=s���m�KW�IO!����q�?�mD��3���=��1�]�l��3if2�!�M�X�7>d�W��]m��M�����<3�E'�L(�=��Ӵd�����2�Y�/NP٨I�Z�5w�{G0"9�{�:g��%��Mӑdn)����}SH$���2~"�n~>��Od2���]ɯ�U��\����B4���bN+���P���g򗌾8W)�& ���/�{���O�����`���a08�����q8�V����jjݭ|��RH�7Kh3Wv��ں��㭑Q�nD����g����ܧw�q�,ۥ�U&3��\VC�,�S�V�����Y�4	��
�a�����Ju.
��,[�����\���4�4�H��V��${'�N;�n=��]��v@֤��8��Λ)a���뇇�ٰ_9y�Ͷ�#�_�p��Ƒ��j`�R/���O����56���"���xb�a͏ZX�ƿ��c�Q���ljMpc��w%�\��&�������p}6��*���󣕯�9����8���su���,ՄS�w!�/����8���1�2�6�!70h�!Ӟ�@M���Mѐ�w�Cu��Ww�9���4�R~aYͺ[HYͯ�����.��8c�c��ǁ%ά-�'�*��B�Yx�]O�!��jK�冽�J)���� x��T�7�rvഎKq��^��'}���5���әsY����j5t#��a]�u3�i5Y�V;%��#d0ڮBh��H�`�,��ε=验�ŭ�{s:�ŤC��z�b��� �})8���0�-�qO1m�s���=r:���fĳ���@]��\p<?Z�C�;=r�l�l��͉�g6�yp�9�.=�&/�,���P���^/6��I�z-�M}��#���c6~b��}����;���&�����A�织n��{|
�',�+��l;�_n]��{�<z��U�÷.L���x��Ӷf.b7��v*ךּ�����d[�'>5��������>����P}r�͸JpU��q�n�R�Y��Qn�)/Y�Y���1b����5���VtD.�ܼ�𗈖CĹ.�xvG�9�a�x�)�����5��!�#'�&�}Fo��@���TtK�gi�ָ��=����	w��,Ud���}͛eC [:y�^��\M������8X����W�r��]�LZ�8<�leE`��O��a�Cuk9Y*�������S�U�w�E�A!���/ENW�(=��Z����2,����A���N����,)��[
�Q�N57.��u����q��������[������U�8 VG8��>�N���js1�\>�<͘��-w��^�5�.<Dm���j��K:�z' �*��y=<zL��/�&���UH���=��5fy3��^��9@�Eyt��@�����Q|"�xr��B�mf�%Se�9�x�g�({xò���QC:(����c����R��wD ?:�:�ȽJiu�mu���>��5XI�3w�z�x>ە4hR�T�Uz̮Nd5w7�j��ӽ��#�'Hg��/s�.��&[7n�eOr���9h{CZt�YsԼ�5<�Y�2q��E�Z��3b��9T�21R���~�/�QViӼΕ�]�L���)[�Mפ��d��^��#�^8�Y���[ �tk��$�W�9U����5C{�m�z������N���8z���׃}�%Z�sD8ttQ=�$�0���_(���U}Z7��&:D)Sx�b��Ϗ���U|�ӪIf����y��3D�]y�&֟@P�*`ke�K|�N8�bek�-�^��G0��*q�5�wZs_���u،e�aܗObtZ� 8^�O�[�o�� �e�Xꨎ�nZ�Ek��]�rP�iC�^k����Y����Ҭ�`?�'�.������?���GL�U���k�9���+���i�נ	�nǠ8̹�
N�qEj��p�­�w1�[���׎�
ƺ���f�ut=1�z��^E�����%G��ʇD��`3`."ۍKN��s{e[�eQC���%�j/��cZ}yC�Wd�Id��-۲�)�+��=:��
�U��]t�������6�P]�@TN=��Ʈ���ƥ�B�vd��t(�U����	|�jv&�h�ݝ����|=����1P�Cs�m���������^�.U 75{��M�9HL�1eY"�_m9�g��y�p2ע�Ep���>SI�4�(��ҜI|�&Bo��5�fYU�ڞ��o4�wkuL�C�H�cl�Ϥ�K0,���]���Pո��U�1'A?���Da~��_%3Y�����=��j;���f-s~gUO���^��і$��}ĺ�*�7o�3:�G�b�D�3��r���%���v��.�u�-q���sJ��1�RY�(q�Ws���#1Kޕz���k��Q�{��Jp��U!>�Lk�1��Y2��A��[ �2d�3 ݙ���Z�C�����5��RtY�t�<SL(>�s���׵��A�lY.s���Cg\����C����Ժ�dH�B�������E�s�1������=nZ��s�\��;\���;'k�aӂ2V��zq��dN׶y!UeWC�zO���yt�~b��Ի���芺�ãvVW�-'���nr��<�H�n��$��N�`Z����+��ը�s)�c4���hJ�'۶rѶ�U�4z�@*A��COjP[��dd�΂�X�ϻ�:h�݊"n�<}�2pa���ݬ�e&�w�t4�/r򟘦0M[�3� p���M�(�r�o���e�CV]^l=��<z"X���PPi�N9O�ra��b�;��p�rafwu'�{����襘���-��-��}V��1��F�'6Y@�P�yh�'�Ga��.^F��hU2�z��΃<�A$a�
��FJ�Nf�q�����7���- ��CH/��m9��m����ڡמ����+ur���{0a�y����)a��[�Ɇ8d{kv��,	��: oGj�t�{;���Q��up��ļ�=+�w�����j�[���j����lvlŭ5{���`��w�f��d������;�Q��kq���8��#Y��&s�}1����Ȋ����a��P{�S �:�Q�_LC~~������ �8>0f��d��də� �^�T<w{�o,h/��ܼ\]&oT)�|a���3����Q1�/���>�J����
�LTm�Z��d��u�� ͜a�@q;A�fͷ�cM[<u�	Iǂ]�ڕ!&3�<Gt�t��Ҝ�;W�"$���|�����]  ɖ(����XP=�^�o��<����%��-�Ӯ�G�z-U���{�9�VI�j���(�E�%���}w_���4W�)Z[^_`�R����2o�!��P���B`�3|�i,.%.�.��)��Ǌ4���s���ϧVI��/c���h{��<���=:��d���·�䎝~H{!I.�E7���K	�����t�8Ы=�c1�$i����e�e�Q�H��?���0��3����.e����Uy��b�{YSx�����}׽^琵vm3��1$Fㅐz#`�{0�F! i��=�Ci`@��-�
T4�hYY�{���o�հ�ĊR1����b��n�a:G�9-������r6�a$ʾ��r7!v�dȦ�#�[]��)��M\T
S�[�u��qnA�p�ff�;7���4��G��l�m��]�mv45b`��c	f��b����?���^�e�Z#�-���ىkq�F;��C5W˯�;5�V3���u�j�]�3B�t2{��ǌ�qK�1�/�U�9Q�5/����]�N���u5uq=�@���oA���*-{�lO�bP__�b����xG�)o|U�w��zCp�%�����Q���mѲ��C���v��+���W}y�y}7���=w�'^�Ȝ�E��z��fB����Ou�B�����x�= ������/�A~�ʡF�#z�>NT��O-�X6��n��^i�����������&UN��6���l����̸�����	suD�[���ŗ�\�7��թ[�uԐT�;�$T�ǫ����k��M]y����{�m�!�d_e~o_}Vb�Zmݔ�Z8��;M�����Vu
H9X��',�ȹ��8Q��j��o��iW7�Zى���G�`"W�����x��=g�Wi�eo7`��y���o�\����}�R�j	'�w�S�=�}����Q�)cq+Г8�J�nT�D��S: �A�lK�{K��z�mB=��VQ�a���5g%o���<=BL�5�9ebz��*5k�OtL{u��u���̸�6�.ڧ�Y'v��ٹ ���3�g����S�#]��m�M�ᝲ����f��G3�)@��^��s.�J�^v���G�i�K�	�uh�I�牮B��^�zK$3�IN렔3�߯0�K�[|�{��h߃OfUQ;<���w�<���o��-vvI��룼���4⾾�y����2ބY�]dk�+tA�t���ٵi�j��Tw*�A[(��-<n�\�KslGN�.�x�
�����q��g��Q�B�����Ga9���˛qCp��ok�2/	�:p���p{�S��Ō� �H�ޫFL�k�*�6���3���~����`\����7���lu��v*��l5�N��c�@KZ*���A�8(;Q�kn�a2�vl����Iٳ��#�G��0ORk����G=�=���k��H�BK�wIBu����"Ř��֦����ׄ��(V	o�L�&�,t��/�����,U�_!V��s�Mu��1���4�Y���o�ͬ�~W$�h�2���o<�A�����*�U�nk����[�k9�2N��Ѝngy�V��]3�^N�P�%md	X�9�����I�ܣ��a�9��F��-u'rsא���}���ee��8��a���V�bu�X.q�Ca��w�4Z3�.�s��Y�(��q6���@�*ǀ�+�����3?j;z�쌳�Ƈ��3/+�{
�+Y�<�u�#�{����\�%���P�?p\���|{���:5�$5�w�����Kz��O%
�g�vn��E"���~b��vw;s5�����# ��^U^A�ꀒ�% HA�����"�Z��v|��m�
(��ƹ�U緧����{{{{{{{}�?��&H)����,Z�wfd9�T�SS[�9͊��`��(�������~=���������|���*�����"g�FűDOq��)����mQET�0U2Q�qULE��D����4�X35T��d�
)��vT�Q��QV��*�*65T���1-U^�<Ψ����H��4TI5���8��1UE�SM3UDELTF��1Q$T\�h����IMD^�S�bb"������(������DD�U',h�4S2Q���6�MD1\ڪ"�#�SD�QRELr�T�j
�I�6�L�.���5M��@m�*�(��f,`�51h�5��肶u$QY֚N)�8����L0f��=�b��޺}�~��ؼ���>��f#����Ś�+���C�2Ȩ)����c��d�r�<�/z��/�X��j�0�BQ��I���c`�Y��aFӍ*nM������ �A�id��&L�0f ������=ܺ���
���>z��h��*,��	㯤Yme�g��gd4�����&��<�!��=h��]�M͇;|A�BQ8��L.7���~쐻*������Gq�@��w[���D���q���0T�_P�'��$Zr�,(φ��x~��,����hE{��v�f���ڢf����Y�"������r����J�O��E�4���%�'�s�z}6S�����x��y�{3;�	Y��v��q�j0�M�5��x86E;ǰ>B2�g_�/x�&�ڱ��{�e����J	V��������A,��ϹqG�7�Q\��SC\z�gj{W]Ң�c�Z�e�g���$r���V�(�ñ�rƳ��z K+�����o�YQp��@/�EܸՊ۪�f^���2���-�0��e�|���U
V�,)��F�I=3siwN�����%��Ǌ������aS܌z�������Jr�94�`ވ/b-'%���w=���|�]�3l$�[B�Ӎ�cH�H ��������{�>ۿB��P�I�>�/uf���NE���ﬨꔶp��������R�W���K������g������6����.!� _���M���g,u:�>�S:��"ܮR�U�:�૓FQ\ao�X��4�+�hs�uֶ�^�߳-���" ��W�}_�v@0dɓ30fk��n�N����;�l�����"���A":l�6S����i�'�R�/�>�V���V��f�u_{�c�e�U)<߹M�.�8�Y�;��,0Ϗ(*.��)�9�}QJ�Ma�S-�a��	yO��G�b��L*�.x`8Z�E��RXבچ���||ڜb{
�e�M�h��Tژ=��@,y�]g��6�N8�o�X�/�1��XO�{���÷���VCa魜Ln��k�Ё{ć��!a҅.;�qg�W�+����cҵ�r^��o�M���* �>���<�seȎ3ʂ[�C�.��4���ИfY7�Xkg% ��Medꨒn�*��ENF]��ܔ��k��яK0�8@���L��\:V0k���vN�Kܸvy��&Ԩ)篦�k��n��K�<�:�4_��v?{L�4�Ge����	p�ly����t��ѐ�'�\M�R�{`���K��z/+z�@����JFa�,l�}O,s`3<6(M6�l<�F0Qٺ��C��@�'�V%;�f�o!8�����(k��sג�P��[�m�0V��"���1�*u�O־8�!��~��H}Y�ӇԐ�v�Ň�y>���Ce��Rߘ��UN֛�^���8V]W_�*�'�A)6ºO5��vr�0��������5��˲>�;�|�߷$�yt0�od���t�b�tU�+�f��ɘ0	� ��0�/���z�^ȷػ���z�/|�ܯ'�2�65.R9�A���/�b"���;���v}ڂ��Y\t׫]��!�à��׏v\�2��#��q׺g�ȟ߭_?Ԭ����дk�g!��kÝ��',�ǘ�����^��U�4Y��Z�:YW<J~��S���]�M�־��{lw�Hql� ��m�]�73��~~���Pw]��k��7�Jp ^%�>�N2��I� �ν}�b[�;v+ �x~�R�W�~�ߕ.%�;���XE`�Y��\G6t�.�s�1��P�@�S��K�����Uy�Ez����qC\�}�&q���F��wVUt=Qi��y�r��o�_Q>������6C�ݮ�!��M�"8g�[�z�K�0�&�G(_&�p������n�,b,�ty6���m�#��R�v�;p{# 㳠�ٖ;y�D�C�����xUt�v���f��
ʓ�iA��|��- +�f�,�tØO����_�x��������H����4 o YX~���d���)�e�ye�,���Y�&���9����2�����2�����}�s��W$����ȭ�F��2YGc�Wu�Yڎ<W��oo��T�F��}m�p`8�1�+�y�)��+������f2d� «*o�wV{�ľ��<���8�cl����O����v��ы��=� E�F{�lTz����{�T��ɻ}x�u8�=�vO�/$;d��J~�.-���K��ז�a�鑔�2ol��F/]��AE�N�,���	��2��/x�^����&]����$��n�؂�kjqb��)�3f�����W�����&@�o�����/^�49�73Od}�
�4?<�gI��}����7�#��u���A��T\��ц|>�"�J��*�xf
������7u�ݩ�P���������,2��AI<Y{���O�����oWD>b�]�gF����+�!)��H2jX���UӬ(�Ƕ�x/Mn�P2v��&9�Q��6�l�X�`t8�(d�殈A8�Q,��IW��[t���K�qQ\�����ܩ"�>^����t=�@��͐��Wp���C�%:O�"S��%��&�޹�N稪�6�U׷�Y��s���6*Y��82��f
o���ޣI>�NT�Ҟ� ��3r��y�C,DGE�w��k�t6�vӹ�-Τ݁\d�֞.Ź5��1{�_'F�DU��{}J?�t��-�Fg^�<S�9諁��J���6��!1��X�2�bU:�Y�A%P6	�WCo��t��M�i�BP��[�W�u�����x�|~�&s��=WY�7i\N��;u�?gFt�pq�7��۸��ϽUI�`(�Yz6}#�gh~70����3��Ύ<k�CZ�BO8ǲ���[��Qk�Xb��x��Z;5@�ǂ7W�=�`�{(���k�_Q�x�Ȕ�P|�앬o��yW0����+�Y�R�y�$2��"��~�!�Y���委v�y��o"4Ү^��W�H�T#���z}b1 d���Ct��Z���"��Գ,�4#�a�ك�P�#�®PΏ.�0��E_K
�`�4���g��gd4�4l�B��X��ګ���H�����7���	r
�iO���E�{m���������7s���i�{�@�+z^�'��ݓnj�l�o���	lNU���a����$k%{��A�T"K@�����T�PbaQ�d_��n��z�`�~�(
��$��X-�M}��?����v� �0�'����gS���^Y�k�hq����ǰ��}�1KƹkV��<�R����c�%�*,��a�kO5j��
��j=;}8�-���9��RY$5��=ٽ���(�{Θ��IS��v����}�ک��t{����yr\��3^��NJ=/i�VMc {��{Ww�ã���J�$�p��9}�R{w1"77���}#�kH�/�̲��AV��зf>����ْ×�x�p�M�C>ӷ6(�w��n�_L�����0�2d�0��ݹ§��8G�"4��c��M�]��m�����;'��%�x��g�c���z}�k�Od��W�<d�dW�˞p̸d�)�T���zu�d:���2ױ�):�-U�K��1;6M�U�[�=���Y���Y4�)��g��w#�'5dqơ�	�{�a��E�5�r��^:�9{�����3��P�D@��##Ĳd$ƿC�L9�V�1��1�`�s��WCGff�v^ԩ2����h_Id������K
�!��s�n5`n{�p�MM+]���H.����K����QL3��j�N0�x�\�v�8��/(p�Km������v;�����`�l:�>�X�/%�r�$��L*��\���W(����;P�3���)R'����ͫ���d���A|� B�����ץ�]T�f����6gV­t��U�*郤R��Y����n�ڜ: � �
�@!Y� tq�n��V�[u��Jד�s��"��V.�F�Fr�Rz-��m�fqPK1$
�1.8C񁅇���#'콞#O��w1���m�����&�b��'XHp9X{o9�jH��7C;�
;�x����� 56Y�wlj֟�<z`9��a��/LA�7)��)υhٛ��r'$����ZX�=��k�z�}�� �t��G�f�RVu�G�Dg��A�{���%�H���M��&L� ��/]�����z�x������F=9����-��[`BN�h��#m�.�s�:4�LM�'��+�S4���v(a�L8�����D&^�Gdc�+VJxk��833��pZ�������b�51x�t����F��|���C�Jy�L�M��e]ocS��i���<J�����k�@P��>dx��zm��"�-��7��,��"k�W)E@�~�/Ux��p�̎��
m����C��&a��@�̚/bj5�leT�5.R=���!�˷s�VV\{Ͽ<�&"��P�����n�~����PWƍ\q�|Q���\�\�5����]�l%b4�aUVxo8\�~A��ƻ�"yWN\������kS���(�z0�O�&B�7.F4��<q�I��^!��t�B.�S�J`�AS>`+g'-�_q�=z.1�EϬ՚n�BD���9]'2X,���1�b�h�D�eW�L�N��K"�9��F�?����!=S�䛕T]ng2�P͒B`SԺۜ�J�5���%��R���'3��{����;���ꀸ_⻶�k4W`�Z'�����;������kgn��S�Z8����@��U]拕�V7�L:���4�|`��}ұ��Wm��wSɨpU�:�2�^L؈�V�U���a��c)�ʒ��޸�Sn+�J���6`�"���	�2` dɐ��;ٻ�+f:����$�J�0͌�:n�0t��У`a��*���z���a6��\n1^�K��5������3�ue¸!���f�{9-%�t���WJ�UI��4ٖ��L��Öˡ�s7�T;��@���c�􎀎��ں��>�f.����&�y�\Wvib�r�1��ek���W�q���P��9��@A��(<#��el4�S6�F�S[�!̹�M���1�
:�/��q��6��K1�b�GӘ%	��a�1hX��^���}c~������f�|�y9/g���c�^���b�t<�j-�� ��h��V �Tvk�]a��j�D���� A���P��:�oP|�s>!���
��E,�*��M�=���l�d1�[�A��uC"Y��S��'�&/�oP��4�1vyiV��>�#k7~�*����zy�����R�3T*���&||�95>�}(�l���bN��D���VwK6#�CY8��v�׳f���o
�E;��a�z�m*�FC�h��������*�E�C;n���.����`�9������θE��W{�BG�,햛�b��=�ݔǎ�^匧[p�u;fh�<�,�� ���lR"�Y�9��g`�(�ږ/�,�ѢU�q^h��9lYs��UU}�>�&L�0 0��6���U��IYr��ECD`��^��Uoj+ӥ	M��LV)���]:��ս4��}��s��;b����ZSݵy�.��O	���1���!
%W7;��o�D�/i)�O��h�]J̕�G:ߺ����樂��>ʿ��]��q zy�70�GV�'mfDJt�������*�-�ۈ�:�r��Vm�w���|&����k�����u��VA#��5!��ܯ+�X7�Gv����g8[�{�m5�9��e闝��z!�`��C��n*��^�ւRٰ�Z��g���N�V�e^��;��ս���r�"H����UqA�
1�އ#�q"JB�'R�鈡�۵�q���+i�^����&i��.xV�k[�1g/$X�H�?�,���q��&�����<s�p+.���c}"y�	��B;�����O���5�1��9�S�ʙZ�"w��޽r��c~߫4��fjm���D?��P���H�mz*�Eu-�#��cYc����֮��14��2�Vf䧽Ν	�zC�юXJ�����ϵ�K�|�2o�'D���ޛ�������Ad��7�^�͒O�pG���p�t�,m~Oy~�i�)����C?5��S�O���//�xiڽ�>__D��'��΁��sm���2�yk�ۀ���V9&���3��/��4{3��5J���a@�'�U�p9��a�~�30��d ɓ 09��q�_���?+����Z�ו����cC����,���2T3k���t`���6�=Q���B�5��'��0�0�zՅ�Y�y�$�r�)��x~���A�Kus�M��-꾍�E��G�/�M��F{���M�揌��b�O�p%'�I�������U���<4g�0Ak��T�57@z���B7�í�)\�Q�g��6ʲ����qw�\se-ޛS������!v�ya~����`]'����9X�]Z�>݅�p����Wt�}��'�KӬ�L���xF.Xs�cO��>���)�ʇ7�?j�1I�˥�*�_�]��s<ځѼ�͈w#U�)�.�ƣQp�1�$AoG�M܍^4"��x�qÝ�wr=y���7�vf�r-����WH�|���]�6�{"�F7�H1�" �}C%�᭸��>�g�}�4�o��C� ��&Y����uKof���Z�%�vrDM�!y��l��k¯3�񭌨Wy�FaP�.��BS�9ά�F�cyFs��]�jq�^(;q8��±Xa�:�5b�����n(^դ2Rz8���%�8vU�1���xH��� ����{Z��9NN���0`��NCZ-�]�X��,k��,�j޽`����ڄ�E���*Z}�q��)��V#�����XE�M���ɬq�N��2�f��r��u�*5��^s�memҁ�D�հ.�a�}�j�G+��Q����@�Äȣ�G#hM�����v�4�+�>�p2��E��n���Ν���a{(�ŝ��Wd��\����A���IϸD�d�� G˽���N�M`-���S�g1ԉ�NQ�fU�(J7���2fq�VEm|Q��"Ģ/"��4��HXpt��j��qܫUri9��c��I3J���/f=�s�x]<�MN/+h�`�X�S��y#ӷi~��1G��mD-eL[.������T�x�^i��V^����X��|���,ɛ}��&[�I�֞���3�]jSڰ8:;'u�.6:d�8�*���O/�G���:��%�ܺn�HD*:�w�H�{�]�oC��=��t��
9����^�	���H]+f��E>�'L"������snC��>�n�Z�Y;5���_d34��1��p��`�栓C9l��Uڲ���`HD7��q�xVO�e�\.U�����H�X�	�h^d��`�=m�&^\�+�i��1�Ĳ;�Wq�ӹ;7�	׹dn�"Ϊ&vY��a�����Ku'��ΥB��f]�d
~fyu�����G�	����{béb{3ݗZ�0�X�k�c'3��}e^߼�1}jΰ+{˝�'�Z�`u��H��AN�l��MO�G1�t���C�(-}��N���[�}X�&�h;�N��(��%k�+0�3��05�m}SL���^\�Rl�ټ:+����=|�W/i�
�-��?��g$�P���2ھ=ؼ�8���n�h��qj�(��g��_���<�B?q.w��y5�����>�9A�ũ��R���QW��y/�����J}�r?]T-�}�a�¦�.01R�P�fj�3c�9� �g��9����#(vMnT�穚���[W��N�m�X��O��*�(��aH��/\�[��`L�u�<�@,���=���M�#Wm�`�u��()zd�h�,(/,��5�Qm��c]��"Õ���ۋ��r����t�c�N6k��9:�+e��T-o���g|�c���{ݗkZ�½YY_�t�di��)��԰�sk�(7`�%�kt'u��ʽ�S2�4�4�"p��}�b��yu�\dj�.�# ^���9_1���z=�;���{"�Vӝ�b���"}y�N8F�����,��P��ز������.o`2����qI뼼�>Ѓ�gz�-�xv��y��C4�B�;����5���r��������q</V*���"j��f*K�4�UQS4��l�g1�x��~>?�������ߏ���QERW�%U�{�QUDTU݈#�:��i�#l-�珏������~=���������UD�4LKDD�{LG��*
��b��
*
���T�M4�P�^l�-�UO�D�1�*((�������(��mIMQR�D�PS��TQE6��*���������(����	��(���"��8�f���j���R����
b� ��#��"�d�[:��Ӡ&/Y�EM50RT�]Z�Jj*B�
h���	��թ
*�(�"Bu�J���-��z؂�
��"'Z����&h֘�8F��Q�-�����i��
M�UPD�Ԛcj���A��E8���bb�Qf!y���ߙ��F�{z׼�~���=;����2�^yf�g����뜗���y�����*��!��P�������ϯ��[kE�qv��2O	����Ŝ��L*�Os�Z�E�T狛U�3oB�|^f6�v-X핕}iļ�i!��;�	�z��~�c"��2q��E�]<�����nx���]��˦�Gb�\g� ��d�!Y�㟎�}�Bչ����u䚥���f�1����\/_�Q���:�=�T�@�	���P>�hr{�̩=��?e�#�]Uj����R���]AXe�X���+�j[�8�R���lI��@|	�ݬ�zߋ[�	Χμ��o2�e��0̋�͈��^"��yW��G�w�g�;>��[9yחrI8;�++�vU`�1申���.�1G��r��*��wД|��i[+��8Z�@��V�3V\��x�?!��s��X�.&3%'�5�m~͍k�$<���#�+��⧞���w�i�������ty���P ��������5���ʪle�׌Q�٧wzԞ�V�.D�h�[�ȶ�^���c��8`��!r��k�����W<*"&�/�YE�㹽/��>�1=l�';2rV�n���A\[�zv�t��u �9�-���S����g1�:Np�a��`�8�ma}�JwIs`\�������mu��G[��.��r�-�����9�z��m��1�g�
�\ ��*��L���d�3�jn�4;����c~L!%��)	��>���������z��Mi�kс�F�C�+�TI*����ϻ�C��>!��k!�D�V^%9*t����K֯��H�䕗h�fͬ���jq�!�>��h/���!
�q���):,�ȺQ��i��O�0b��?b���%����Dv[�7��%�>�HP����n)���5`�"�u*���Θ���3�mm��.3qU��ٻ��a�a�r��@�p����O�>�!���ta��*����bΘ��c!Jǉ��g�Y��u��&4&���K����v�.6a�=�l�1:�c#H�{�K��N�jr�������=�j;��}rﱎ0z�;aA����� #��(~bk�����v�%6��[�f~����k[+ʱ�{�J�)�z�>6��	��n[�Y!�`�
���J�oL��7������\��i�D�(i�E���Ԏ�<�+՝S��,�m�J=ʁED���>�v;MQ��-�PfCF@{��r�*����@'�*�e1�h�9��z��+�a�4jJ�6�YA�DcA����퀏qv�rm>ȢSWK5�Z/��j��̽�`|�Ӷ���yV�Wѫ��ISB{QU��)W��:�ܻs|�f�y�{���]�x��ފy���7�m��b��Ng�41���|�Pzr�	��
���s>0jo��dɐ`�3u�SP=�=ރ/xaB)Xp�%8�.~���t�4��a^����+��}���6��`�~�_8o#�~�Y���œ��@W�P����EC��D���s;ĳ�uG�0���7�K=-\Z]b��8f����ݪ�ɚVd�#��8H�t5z*9��'6\���`�ABk�	ɚs������dp���u�l�/�(�\T�f���dXiGh><?���~�DW]|��l��?iP�����YΠǦ��7��[/>��%6�2�\�����f������yp˗Ut��l�m�]w@pP��an�{��E���
�D �P�Y���d��j��9��d�n�'�'�u+Ś����˄�J!�a��􊇚\G_�@� ^I���)�`3��ol5~4����1f5.��{Z�sg3��sƍ>Ta�^zu���Ƹ�������VA#��K�=hXE�7:�3�j���=<���DO.��<ƶ�$�8ۏZ�y�\�"!�"mzc�m���f�����]}�"Wgj���*]�Z����?"�-�Ը��]� =�|�l���k	����g��d�ͮR;=�
�OH΢$���l���2�5|9v�j9}�fa��j�)f��}��}��'�(��8�ğ�U���^I�x0�Z���1��a�Q�,����[��	q�丑��,r#�w��z�Vd���`=Oz�#�G�67�L�dɘ �6�{�j�ʱN>�˞���ʵ��EⅩuԍ��Rܼ��N��∎~���bzU��wu�鬾�<7��D�{�H&����)�������)?5�b2m��)򨁙Rˢ�A!��mF��������k̂������T:8��a^���]L��C���e�k��C�$�>�3��U>_�΋^��3�9�-nAV�a���x_=�k�e��͢\lР:]m40�.�/7]�ȰB�@�I�K��dCQ{��r�X|*ՎZ|��k��Ǎ���Ǹ�g���3��U��\�f�]�z��Y�Q��GN��C|�����\K���]���-9N�#~�&�Ȱ*��b!1��V�<6�_�F_H��I�jJq���݇7���m<�>Q��R5ӹ9�q����npj���{�b���ϕ�|�<����!�ڌ�=zsj�����*���#ˡ�N�c f����M�F�TV2�!>��A=,�,^�n����Z�[�hD]wn��uє�g����@�⡻��B�Cƣ�{<o�������Z�q/���B�G�.�}ޙ7`O2'�j�/wzbM\"�Dw�;��
�M�]��+>S1�	�5M��_��<oe��!	�3��̆nm�i��`�fmx����.��9	{}P�Uܥ��VUf�����o�1�9P=~qJ5f��|��|ffo7�L��d�3  ��͛��Y~���nwW�md��3���-�Q㐥�J�� >�����?�f"��(�j|�[��k3Qle�	�{���T-)��¸�ȝ����a��}�A��]�?3,�i�v��Nf�Wl� ֺ�oQ��x	��9�Qz+�b:l�y�-��@Ue'�m��|�9G�/�`����_� ��@�U|i��B�䧛��Y��9�o<��vk��"Q���˫sg��:� ��m�gZb�
9d�fȣ~�I�TY��b18�E� *u������;��&�ϏkϷ��GؚA��b��\r;�9���-u��ӯ��oE�g��jœ!��{ne^t-k�7<G�r�ؼ�v�(pX}+9���ʦ6Ǆ_+n���XE99��[nmg#�)y���a(%�ң�H[Bu�s�If;�0&&�h���_,�����?n�޾�n`]��5�VqT��{���lك�q	�z���!'5¼Ǻ�Ӈ�h����Umxu�&s�]Q-�����������9�C���]��=���!EyG5���P�^�,�$Tq�ʽ���A�����6@��������Sx�{�����2;[Є�ÎUp�_�M�y���\���X���k��#3cV�U���|���k���C<V˚W�a�u]ϴeҽ��'���.K��������络�u�}�B~�@L�(f`�^��ٲz�7[�A��x?r�u�¢�؛�m;�|�CzA!�(4��L2�­8�u��0R�l��1[o�g	��Yp�����^=��6+��# ��ݎG<�s�O��*�OU���(�R�B�!���g��v(*�N�NR�D]��^�j<6�[XI�QU|����,�C����2�/,�QG�T7��.:kڡW�3~1��g]k< ��]�ʱ�uk���校	M�9HL�e�X��^л�5��ռ4�{gh@ŷA��5T���sf��{�B�^!�_)殄%2��NJ�J`��J�b2s��C_q�9�`Ե��!M.ה��*��{a@�Q}�8s���<�� ��>�锝`�&�[n} [=i0���� ��J=lj���[N��yV�0y�߈���K�����K�E��QuwN��_:������ov��r�9d-7��―n�ه���S7_w�i;��`�㼭Y��������y\:��~k�PX����8��m¶M��b�yg$t������xo�㷑�����b߸��5��S�x���;��H�֏q�`y(���U�̉d�h3ի#�z��Z�oũ��wH�;�m�MAL�nm8�4�s�6m�?w�96��6���Q��"s�j������fLD��4��L2dɘ�Mh�Yގ
=�F�?����-��'˘[}���F�=��s'Ԩw=,c�T�������.j�1��[��O�z�i�
��	�d�J������q�\���U
����&�͏D,��Q+3f$��O�ٕ~���\�����d����7O���O�ϒ�Y����͈06�	�f�]��T���љU�;Fx
pJ9�qa���t�yX���1�s��ˬ0��]��l��FX�T^�d�MZ��xk|�?�ƣb�xwA�x`��\<(��/x�oH~�X���BaT�^DF���t^kHq�.cU�M�.�|�S�I"4ɐ8L�C�$��o'0�R�HK%-�R�;�������9���3J�Lx���B��S��3�_�KL��aqf��|�5�u�B/m1&�+���}9�6TS�S�糔H1�`d�t�������m���A^=R�)��# JQ�؛��)����5=2�(r:X��1�ڇ�3��R��Mu�҄���(2jb�OaWN��z/���=x��u-ރ�=�ju�/����7X4����yGd!Y&����yD�/~IM22�}���5�6����^�[�T]�x����E��7=��0y��t��n�o�??:����]�ⶵ�ʝ��R��&#u����
'T�r��\�X��^Dt�;ƯM�x�~I������o���)Q:��d�{ӂ���^O0~0�nd�&L�`ӫ\�k��mcS�S�|^�����(>Q%ٲ��`��+����N��޹��SV��(�<u��y�n��-�i5��ڍ2��t�vq�V�~w&�謂B�4׷o��3*���g��;k�a�Ԩ�:"�����fƪ,R1i��<�-�B=r!6�VT�����[#f��k��R�zKR{�e�˦�}���'�uOf�-�D6ㅐ���ؼ=�ҎZ7rN�Y}	ó�/~�i�9M��i�����*;��O��Ļ�L�-��v���iv�{��G3�^�d/�@���W��tz��7{��'��FM�ߩO�����:����޾���dL��	�H��r
�{��T3�k�H�mz^Ȯ��4���+���K2oLy]����+�Qs���F�KeG c�S`XS�~:`:��S��^�w�Jp�:���\.:�9qi��"{K���k�Ղ��2��qV#
:��D��BjNl+���ds{wYT�j�Q4<�8�M{��v�Ŵ$E��;<R�����A�	��^�C��Ano�7t��@̮���Ն�-��E;a�T��y��b��w;���$1S�8[�W2�u�H��y:!g;A!�V1R�Owayu�/w��![��:x��z�s�|�N��q�*G~�M��^�]��mX#�{&ѩ�����y��	̃3&L�`�ٞ���y���,o�c��[a���ޟfّ9�O;PJp�3ۻ0dyY�-/)�ץ���F��+�����׫@t�a�� �c4���|�m!l%���l�����Q�g�v����q��!cFi�X܁�l��^��(��"C�)�Ԑ��7jQ��}���(���lϽ�v.S��|�.���8#-�zu�)�(p�am����XܴcD�<c�<���u�6������:�o�5�!��ۊ.V���,)��[gT\:�q��"z<�Ⱥ�I��.�DS���ש+�u3�O6�x�&I�)��"�UE8���;���1����k�x�z�;=9��ڬb�ǚT��[�j��b�&X^b���(���7���P�1�],����I�ջOל� ��>�� ]\�@�ُ	eB��������6����s-ǁ���J&\T�4#[������%컄��*Y-)���Z�\sЗ��dI�4�UE���b�E癎鄊�t��������X�ٓxw��Q��[c��L�_d�P�X^��/���1���}�,�Mb~�}�M��ܫM��%��QM�ȶ*g\ɑ��[��ք�ɓ&�����s����ɉ�u+<�:�~��ӣޕ��q(��=��9��Νr�Y-_����_�u|J��}�q]�P�8�ժ{��=}k�~��v�� ��s���+
vF]^�-a|c��L��������qht9-=�(j�0��J��޳.o3�Wu��v���$���1�Z�y�U*9�	�db��C!���CE�rg8��zM$�]w]����k�f[ Z��Z�qT]o��;NP͘8e�V�2
�p�P�]'�^r�%mᨈV5\#XC�+|�f��e�g;+�Wy�*�4{w�f{C��1�X�I������.j��}uO.��@�B+;I}a�Ql��Ӱ�y^w�+Г���,��0�s`M�/u=}��P�pE��^)SB�kpJ5�GV����ܨD�b�y�M����3;��T�����>!u�j�}�����#Eq5��t������|��v��kQ�{3h��s��Φ�[��k^�]yl ʂ̡F��{�T7��.:kծ���`���9ؐ)�g.��Y�~������ �#`Vܷ5xt)��	�yb�I��H��0T�9�\��Y#�ɟ~31��Wi�I��!���}wR	���"ʞj�BS+�S��0LRU�ɼt�*/��Y�̓;�v:a�����b��Ț�pRk�Q|�4�ur+�(wN���Z'���k[�M���^Ӷ�x��OqLOA)�veڅĸv-}M�(i��l�����f����}A�x�qn��0f���n�ͽ�po}�/���x��7���z�{�]K�N$��W��%ȟiXX+C�H2h����v�Og��k<��u��q^��v���c��b����Ǣ�0�mȮ�K�~��!�E�����&R�̓��Y+�?i�!)[�u�������7��P��x����7yO����
B-1�	��	�Q�4��W�)����N��:��x�:P��ﰃҮ�w.�����r	��쪻��[��&1Ȓ����J�R��#}���fl�e�ן&�.�S�9uj5Y0Bs-<j �?��Y�g4@T�Wz����o08iҬ�Ō���p�ҖӥH��e�l�)>�ʧ�f"���囩�ޗK�Ǻ0��&8Fp�W���ƭވ�-���̴�,!���Ȋ�9������r�ˇ[�{�73���m:������4<��kmW{��zxq��;z��tN�[SF���5�l[r�-�+sY�t�����`��xO8��+�o7�Q��Q
�L��z�y��N�L��$��{���f��e����gwX�ypr]W�B<�_&��4,=5κ�os�!����ՙ�ϥ�[&m֛v�Z��IǞ��5��KN~O#%*a��ɧ4��w���R�K�7<��f�؉y�?YS]e7:�E&�sv���H'���
�bx��w�ܰt_{)���}��x���$[��V�Q�
B��kp��+� /��#^��=���3g-˵��i�*N�����^+�[��B����p���-D� ����>��Ь��"Y��ei'�jh�|���Ek�j�����>g	��8Ѱ)g:`�vv��]�K��_n:�ݰUnA��i��ų`L廮{�Ѽ���/q)�w+��)�0��	W}o�_Ҙ���9��nĥ�����<�¬
��ҳ4m��$h�-�cw6�lo8�1�Swk�e����f�]>�2�g�h�7����o,`Yu-ջv-�Ґ��V4��֙�aR��y���a ��WNg^��>�LGf�W�O9_ъ5c1g�&�E�F�Q�����L�������Y�b<�հt�;O?e�")��N�����w)�E�`^om �G�u�����fJu�5q��>z���[Y�J���%�z]�r����5�c�6�o���Lw��s��һ�f��2����Ȇ�..N�6�[�Kl��T�>qۭ�	W������ζ8�S&n�������r,.�t���jQ����WO>�`ڶ��
�;	��3����.O��t�k�4ĜB,�^��UEAAPL�x��]X&hi���&��(��*�+Y�gV��-9�����������oooooo������Z���Oq��&��H�&&ZJ����&zz||~���oǷ����������r)�4�UUEE�n4T4�I�0K3L���'�*X��*(J�*���� �����(*
���QEEEM7#5DA2U�tS͆*��������*�hj�������D�A-�D�TTEAL�SDTQU	N�5T�D�Q1U#�ETLQUA SS5ML��Q%�QDT�JP�]cPTTO1��*���"����J�&
"*h*����(������ ���*"���T\ƒ������rGVh�i*b�$�EERSDIW�T�RQD�Q�4SU1A�KT5TD�SA3EDDDEE4C�p����nP8�$pV��`8�%��_zl/{g/},U_6�-�x�3�����x��J��X6_HU�:ȠeaY��7����6"�J4���d&�B����0�M|]�<mDT�#UM)��(&/��nd��dɘa�L^d=�uS�������X^Ǥ=�,�Gv>�OW����(!��_h��/� �� |g�=�2���YY�ǇV�=M+ >��q�1۽0�p���jr��Xp��8��}�"�=��}}��ǝ,��z�Վ��Ge?��h�=���w�_by9;y.ru�V�d����93�r\��d8�՛"wx��t�+WY�˘]��tLe��٨��Csh���Ӊ8yy�n��:�"Є��[�pv�!&֟G���gE�cU�ЍNo+� �2X&�+(]�Ta�֣���e�祐8��y���G�D�1ޚ�{�{�ŕ�|����S��;\��ɛa�ac����{�(�W0͹�l�0kl4Mw2ٷ�yY��u�l������!z���2� �Lm�u>X�>�~/��|f�18�uw;~�3��:L�=�F8>d��\'lԡ�Z���y\7� �@��_�1�I|1�9/!I!��1��Y���
��������xI�-!�8^<��,�	{�J��?��s��{�T��a��hz�- �'�K������S�}0xyiFOr}3��z����g�y����z�D�9F*�btM�M���{�CoTһ&kuݓ��y4Uz*%�����]�����[�ѦbWR���+w�V2z�<f̖�mA
o�7n^QzN��}���*�v�����y�zT��SG,4��&T8��o���&L�aW�v�MdZa�i��=�CZFnu3Od�K(!Hɇ�/,���8�������huv�������}[J�Z�Bu?_��Ҟ��cH\�3m������9!�fͧ�z��[�T�0���8e�Z����\�"�ҩUc���H�"Sm�5,S~����\@g(@,\R@�>�"w��䬧\�o�}��r%�X��� Wl�2�h���Y�d���������}�h�����b�Y�ྡྷ8���a�g��6��`��3��y�`�}Ȏ��7�%��{8�}/����˗�[+���F��F�.��c�q�(�?ts��
/�Vվ���G{�������R�Ą�RO�1���(�a��Ϻl����A�@B�z�����fmt�mJa������K���&�~OI��	zyH��,0��*'q�L»�n���ބXr*1�C��L<1ס;�M��kZ���V�kr����>;��QA�G1�6���O�����	���@2�b�tw���LcJ�2����F��zUyG6J2����I�L^���nT�#%�f�.�1C�9�<�nl��ˋh�[�z�>��cc6����=��g����d���$�j*��Z�[G�^���[3:��|]��k��V�ٖ\����l��z)����ӽ�}�����G�)@���qq(Dx7�-�dɐf`��~�tꞠ�����s�ޒ'c��,!�,�ѵڦ��/MV�K�PIv}���Y��b�e沲�N�u�CM�u5a�Q!4���[� ��§C���z��V2י'����r苎��!�\�pA���mq�桫-2ڨ$����GÖ���)�*OCllx��λ3&�[�`g��cz��3��ƭ�W��ވ��˚���r��f�B]�8�ޑ8�"��q5|�L�H$�)<������m]�8�VK��%�(�A�0Ә��=p�ۍ-Q�J�-�r˜Y��E;ǰl	!��FN2/sW>�yխ!lt���!���w:�a&�f渣����z�Y]c�jc��9��	y�Ȱ�A�X@:ƥ�B~k��)�ӽTt,���z�5X��R��f��R5��_���pJ9�E���*by�WN�m�͈�on�۽�]�"��Q�Y�{����D�QaM^[s"�����O���?Ai�����5���V.~���۲�!Z�njY'.��IP�j����oM��R{�H�?��%���6���4��uV�)�qI]u�o�/����v������N
�b��}y|����~
*�i Q$�x�ݍ���O�o_u^��m��87���h����i�Vܘ�� ��B��"һ͵`����j� uzI����8�>x{��W���ɓ&@��ߟ�.������P���l'�`���i2��m�(�AN8�8���X��DF�dU�Z�pn�8���0C�{��gd�L9�_@�T/�;M�IO<��H���o��ˤ�;y���V��~x�g�u�b���v(u��)�(6(��<�xY���jۆEԐ�E��w����{P�<Ƃ;P�Sø��ͥa�`,�� u6>=�QL_P��[1<2g�M7�;uf�e�n�����$KWdaة�8�+vXeC�ht�csd	��kFd@�ZwFc�ٵ�K3��������X�d)%�Ҡ�[�#ꠖƸ!��G��"^ߎ��j�n��eL����f^�a�Y�P4{"|�������[,47\z���i�ȫfx��'�v�;P�t8l�`��<�
�ؘfI�l;n�e���0����30�b�멣�oU3u�L��hjY��%�S�2�ڑ~^"�^�mz��=9�V+�4�ZL���v3�s�?܌��hv{@�-3�� ,bJeĈ̔����7�<����l5��C�T����_�G� ���ɝ������+��ŝ���)����| �=s��eq��o[]��`h���89f�Q�}5�;����_l�1����w��1�����oj��`��ܫ:4ne�9���ށ7Ʋ���������A2d $�˾�̳͞Q5�W�҇�3�]y���3`���V"�ߚ�Fۦ�=��9�O�� �������<û��ī�:7�1)UKcW��!s�������P�`�<����L2�)��,�:mm�r�.&pʋc��Y����,�!!S�ut�Kss�	���,T):����5�cռ5Ҕ�%#oz6@	��=9��n2d�\I|���AC&}�!��T��%2,��R�&�)*��<�����_���u�"��^ŧ��`�i2$��B�����H��j��n�Ҝ��)6}UP�����:��]9��E��Ѻ�p|z�%z��N+09�w�;���"�H�@_Qw���i�ꞈLI� �?Յ��Ʒ!��G6�� c��wl�X�%�C�6i���ɗsI��V�-��Z��9��(aCM'qT-*�{OIa�Xsm�՝ �K<��1�Ǎ���s
��T�tgdWGw^�������1)�*KՄ��qTa�z�w9oL�έ�5��H'i�*w\�����3j@O��:����SA�ǡÒ�Bb[l��Z	�a>�ҵ�9/R�X��6ѯ71Ɗ�]�=*�G���>�lU��=~��ޭJ�R�|0�8v�v���-��y���s��'�$�y7Gk�>��?*Қ�+;���M\�ss��;�yF�|���S,�<]�����`j���ze<�>��"O����{�a8���|��,YXgnvF��OM����L)��p�p|ԩ����虥}�G�t&!>�ޘ�[�Ǳ�r)�ʍ��nOb�uM�נQ�����N,?j���8�+����	�{>����/�r4��h��17]]�����ng<��)�P���<$��,j���U7���y��u��M�Z����n���L!�tC�e�81����Sy(tZ�z �K�<�&�@���ʙ���ٛ���^K�E�1����{ ��	e��)?t��'6\���"�̜�������ÇAi���W5=���ZQ�L�vb�-�2(���6��Y�L��R�d��a�S� ���B��q@zvQ�6��r�y��%6�)A�R�4�;.�D�1���^�w�߻����g����m��S;���d��ar@$:�F��\��'T��없�Ts�:�8��u�yL��ӳ�
�w�^2'rW(iT����]�*a0W��̎a���4�-�s���:)�r�	�]"��(�kk���^zuӎ�8�a��	�rͭꉟe��.����`��eu3aԼ�R{{�CL������X�!Q�_kWiy�H��RL�'a7�y:��,R��n����4�w��)WE��wܯ!��:���E�!��H,�xw#Y9���5h�4��k���g�V��ԯ�.f����{�7��{eD�j��r���󸐸ںO�"����(�*����w�#ϡ�Z�=\�%�a)��nea��Z0,�g�3xi`V����z-?,O ��o)K��[��\�Z�2�s:��ן����b5��u��t�L^D��tx�{c�<��uԶ�1<�����q�����$��ᥖ��r{~Ć�n$_�Cc��F�˽R	�W��Suz;���zR~b5��6"%�S^o�e�c�{Ɲ�*�'!��b�\�M�[�Pఇm
�^@tqw''���"�
�f����i	ͻ���s}�K	���C%��bN�@M���nAM�A})æ-p��_��jq%�w��WWx��{;�[yP���Chؒ��2�Tx�+	�N_p<�f�����3�˶�Q���KYx�]Bz���Mf�}y;	]�^F�z"���4'�;�9KO�pjм��]{U�Q��z<��	hP (M10��b�)͍������'�k�� v�9Ͳ��Q9��g�]J��;:L���e����<��"�u���@T�Ϩ���!lP91k�W\��~��w�P\� �N]���Dt�H�u3xVBv���c	��nb%3*���:B[��x���'�K�٬�����y�0���Q���i˅cV/VD�m�]�U*�o�6�-$�'g<(r� PVa��pݴh�7��Ŝ��G';L�Y�:ϛ�k��wX�� �%�5�Ň�P{�H��r���e-3�4�ڶ���nz�l��g9����YX�ӌ�u�5xeE�٧�p���x�=0��U����
Y�]΍dv��,��\��X��S��"z�gH��/G!K��E8ZY��`.0���6����d�!hL.v�fG	қ�wL��"S�H�XzL���FͰ�Ǣ�"֍ʌ�j�z���W9naaQqIpq C�e[��H��*�,�&*ۤQzq�b�w23],����T�]u�&e9����1fYӴs�48ъc�0zZ�e�cyVs��]��|�F��	Y;��{c��q8�� ��m�jC��H��Vl����7.ȝm�կ�r��'q�!9��q��Q����N�fˑ rt��yה�!q�wo�(-���w[�9�z�����FT��@��X��"���k��̩���r���`!iu�0�V�R���J��E�՟9UYM�jÙ8���u�Ϻ��Q�� uȋ3��������|j>��� D	ݴ���ҝ�<���Zͽm��������J�Zqb��z��g�CّWL�x�����6�D���h��U���:a{�9jSбd��3C;#�e�ޗ�@��l]���]����sa94��o�<�x`V�zlݨQ�	���ň*���]���3OɮQ�bd�T�ո>�OX��;�7]����3��m�Mc��s���~y]�mEu�܃{|�?�ܿ:����'�PQ�����erw�y#龍"��s����6���Ӧ��ʽ1{g�8p������b��j,/j�u�%�^�m_��<��$R�N�mC�r��x����.�����l8"�F�S�u���@��ˌ �I�z/��y[ ٴآ�y��m�\�i�!��^�Y!@3�ی�M����b9� �8��[��2�3ne�u��ص\��P'��KcR��As��4�( �:���d@,�V��i�m���3�W��.�� ��Yq����Ym�;R�o���M|�&(,T)=��@�^<	`}�'0�]u/ϗڷޮ�Nl����="�DD����r��!<��%9��0M*Ӄ}�)�ʟ�uE�@l�1Kחj��D�I�\j����V��^��2���-K�-;��O�����~x7�ȷ^z�9��u�i0��\P{�}Sh �\��xnC�U��H���Mv"ׯ�X�4�#U���Ū���ү�~���~WU�����	C�7s����-q�͘����<����B���-s�rν�Ky�$�nNV9m�V���w��2����.���3w����=��cΧ���5@ܺT<�ŋ%uU��W�޽Թ�yq�����9ï$d�疙Hk,p	�!�a~�h���;����ν��w���;/4)_�RweOC�(���⠱��a��'�v���{��m.�f�WYRu�r���e��D&�C�sBvSj9e�qTa�Z�c
����4�a��i6Ƒv���5�s5vJ�Aa�(� ��]-�DI����&�>d�y�֨PKܽҁ���>�g�[��v�&lC���4/��O^Q���7�f*��m
9P�c������7�j�m��g����n`Sb�Q�kpJ���~O0��^��'�����r{�K��v��R�{���GTe������GXnY�X��t��w�y���ㄟmd��r���=�S�F��CMki�>Фf�\ln��bSP�yu�NU��=י��������:���l��e<�ͯ@���i��%�RYA
ɇ�y�o�F�+۶Js������C�ϡZ25*mYn�v�SV�1��$����z#N�zLϞ��&��!��hYw�Q�2�Y�ܡ:-N��i�v$š������<~^�J�²��o�	�[�v���0��]�׹xg)YJq�E�66�U�k��=�5�{���f�F�sx=�xln�������x⭠��֮۩l^P�Ю�2V������1<��p�}7 ��eR��<��qn��<��f�yVv]��b�}�w�j��绖��V{P�{1�����FY/'N�;�>V+ĕ�����MOL���I�}�B�X.�r.wv��okV&3{�b�K���^vF	zy�s�q=^��|�u��Yr����7�{��r�>�C��)�a[�P�J���r�W��ڥh���5��#�+!���%�E�i��H�X��6^���1��(-��C��I<�罒�񊝷�:��ehX��^/��}�sɻp�I�f-W�-��0�J�ʽ��}QET|���8��媁gYB�ڗ��������y��Vf?A/x�.I8��i�t2�ׁm��go�-���s�Y_�Sj����Viq������]{.��N;�z��o���x�U8wE𨲆�Ff�����A��
@�b�����u$��#BC�c���o����ܟmV]�*������w'h��I+�t��A{��֯}N�=y$�VnJ�������Ӳ{".��99-�r^�<�t���\Ӯ�\)j�������_G��E��z�p)s�ˣ��'w���O��G��s�#��T����U�WٷF�k�u�/~�:E">n{�r��Z�+d6k�e�'3�f�Z�SS7�2no>�'tq�0�kM9�h^p��9M�(�d*]�%Ӧaץ���m�	�G9��Ŝ�z��Z�s:jS4t�*���Z9Wd5�t��nW`8��ӯ]�����˂���K8@��.�E�{ �i�`c�ie�����T[Y4��{�nN�	G��5�}7����׼�jUyUֳZ;�E՚��Av*-XYg-�ɜ��������N�w]��$<˥kT����K�:��Kh;��e��^�6~gN3��UY���w�P�+��I;�g\[���<�?X�T|����.��f�VE����]_�b���m���m�+��f]1��/S�l��Rv��-�z&gV��+�hz�-(&*(�A�˲>���{+�^��z+ޥDK�{m��7N ��C��eW�wz�ѡ�JF"�u��x���8��ΏK�n�?mH��Nt���%�p
�*@tzvф�4w�OGmb(��3������'y]��t�(+	�Y��a��=�yWe�I|]դ�OޕA��WݘiH&�S��nH�aL\����QN��p{|
6x��������f��8�oA���mW^tw�o˝-1*�as�!k�s��ru���ID�.M����OD5p����Yy��ֽ����Jj���	 �@$�a�j"� ��$�"��Q3QU1EU�b��9�4��b�i���������������������~>|*���
�� ��j��)��I�(����ƪ)�c�T�L�MQT<�M4I?����>>=�������ߏ�����(��QU{�&5������c`�(���(��b���
(��/��b
i����z�G6*�������*Y�H��i��<$��:�MQDM-UDT�RTLQQAUT��OXMD4l��(*�*��5UQSQ$��:�*:�G��9��W3�*�j����)������-�EQ!QDU������Qu�N�UQLI��TUTT�-Pi�y&� bb���(���SQͦ�i6q��AAPIIM%mE4QA�
j"�ncR�RrUh�UDRMQN� ���"&��(+���EDAUT�S�&h ����I�0j�y9��fn*�0����˾�^]d+�잇fO�:'�=EL�y,u�F�.�KpE�8�����y��ڳ��y������dd�9�,/���U�@���\P[���3󼑻c���;����d͸�d�;TF�ī��Y�����4��;�B�Z����M��"�D��v�y�ʚh����{��1�����uL��Ds�-D�純�+ThUk�qQ\��RN k�.9>�i���Dy��r�h��_�Űu���W��?��4b$��b%9J���&��uȞȸu^��dcq��{�#�dά��],.��t�d��#!��y==�R�ؠQ�Usj=^��y�U�5���5]�B��Χ7���!����	�f�D��P�LY'\�����9�\�4"aڢP�HQ�gkin���6��O�����@C��=�>$��Xt�H�ؓ���[�)@M��f�z������2���Yo��";S�\z(�<���*`�l���ήL�S��5m`��e0��P�]�h�5{���x:RK̨�yT���/�ACB�hW���ڤB��~�^���sѻ+Q�{x9��IO��*�k,Y��b�^�� ��� ̈́
l�������^z���z�b�_~C�םW�"��E���΢6@�u?��y눭o#�\~��	ڒ���=�`ͬB�M6�����7v�u�ب�o��O�.�չD갹Ӂ
PZ�lG�Q��]�'12�	|\�OWP��/ބ֣{�������~s�����Џ-��J[ș"ǲ{����E��lל2���L��NP]y]��*nk��P�(�`��0�z�8��#�!k���B������q�����颒��&��Z;z,r5���֜Y>�`�`��~q�ʃTo���+�nt{'��� ��Mu>Δ��]�;}�fj�x�R����N ����,?y`�s�3'c�m��~Ɗ	�	�Y��{xw,��q��(�kȖY�-�<��N��0���5��+�q��{	�k՞��h�����t$��<�OK K�<U��!T�j���8�	���x�6ˈ����V�dn�0P���$�j0y��c��	�,T)XU\�v�����S�?t�����m�e�y�5�7�B������gAb�:!2N]�9�^S%8�ئ5�2�{:�n�q���slag���.�=�9�yw�Re�/1VØH��X5�֗e���Z�gn��>r���"f0�x<0�?T��0>1X`K*©���Nh�1�ڷ)
����A~NC�^�0�ʜ6� ����8�S�{.ۅȭ�f��g!�����R;�,\�>Ti�j���mT����Sj8�lUWp�ln�5���ٽj�ɪ�e��`���K����ɶ����;�
�h�ŋ|#��[�}8��.Y^V�^��(����?jc����׶W* m8A%�!�P��H�� 
͑FX��D�A�f�"��15�oQ`ؽyH�_��X��Pk�W�ø'�����`��7����ۡ'�����\�t�}�RUk���ҭa!*6p�
Z� ���3:+}Q��ٙʳx����Dʘ�"��Zc�q�X�Vb���Duȋ3���1�d��g�}���i�ń�����\Ή˚��	�g%@��@�{�r�Է5Pک0a�3%��B���l��k����Lp�o-z�_�?|�^4r^�,+�It�άs��Gr��)�8r�����A=������X9D���=<�R��<��7��#0U�Kb'�=Q��E�f��
[uƃw!��)4-<�9>pJ�%����{�I�?=c;y뾝��x��c�E�-]�K�Y!
,SCTzN��R����Wk�tj7/(�v�������r�LO����B�:� Ȭ��8��6m���M�ʞ;J�G-o#�0�Y�F���Эɇ���M��z�r�(^zLċ�)Mh��j���<�l��u{�na�yj�ж"��s*�
V�֍C8웡�h�H�k��
�iÈ���۳�/�WE4�/�Z�������u�s:.�7��ӓ1�'�����Q�H�*�G���/C�3�����{�E����;�H�U劅'�]�;bo#����pG�����O\�1I�(�яF�� O�l�O7:���%?.J C��K�uF]c�'��izc*E+y���eyAJ�`@��<��YN�'�Ƽ�H�vh�t�"���";�7�(x�%�QLJ2�p�\���'�>�ɨ�GZ��g�@��d��n�^˻{�H5}�+T�yJ):a~�R���'z�j�Xt$�JK���	S�����D͌�+�
ڔ�Mֺ{�G&S�9�n�T�eg4��-����[�~�\b<���U��t�־ �L��b9�N�0��7"���^�X�O���Tn�נb�	�/q�����N�u�%�Ƈ�}����]b8w�B������P���%�]��ݎ~���SU)��8e����B� �1÷���V�z���
Λeb9P��l���p�Ӳ�u���ņ}8��sH;R�<��-�)��p�.�L�ϵ9<�{���wn���'��)���m%��ժ�c�Yީd]�����w��Uys���<�,��? �Qf�����^��G�������3f���6z�҈�v�,�	�����}m������\��Ɇ��h��#���r��y?)ݑ��2��ҋ���=-��m`�u�v�G���`ji0>�cE�O,m���U]-�67ufee��d/R�]뀮�(�>��� n��bSW�"�� g���1�˻!����v3r�c��E��3�;�D)�;Cר�kٸe�tq�n��[a
dÉ�i��;�k�E�We�b߽�3���ߩB���1Ň���&=��l�J����)�<{��=�\4.��g�9��'j����7��[���P%'��jT��Ͱ&���q�fY��X�ǜY����r�����:�z1����ر�x�V�΂�r,D�� �y�B�5��v-��C{'-n}y���܎p�D�/~)D��:vD��P|ب�Pҩ'h���u��&��7"�Ԭ�Nv��%�@�#��}Y'�b%9���bQ���r$vEê��h���v�v(˩�ps�j��g���05��լ��^�HM�4��1��_<�4
�a�F�Ӆ�6u�38�7u����^|{`��#��G6��o®j�΄a�i�Y�ygh�	f{~���],�u�Kܙ}�ZS6c}�ułآJD֮��[��sf�3�=��;�Ԧ������D�i�T�"��s��Y��]�S	�F���2��qg���>$*�n�A�i4�F���K�ͦ|Q�+��˞�g��$a濿|>���}��.D�]��v�K�0�lJ�ZvKZ��'({:D�lv'��O�8�>�WK�����Rc<:��|q!�M"��D?�1���ǽ�	�
6lc�kN��;ڌ���8܀���(Gdf���n�q�R�>o"
���GWjǟ['F�_r&c���U�l��	�pѤX�i�;!�k��P[]�� � �'�"{��^3�&�mu]}�[S(|d���'��#tgIN���%�zs^pά��F�&i��8í�~�%��ù���hy
	�������mk�����{���0P�����aϞ���Jw"�2�ʊ�g�A�[0�樨Iݥ�:�7g|�}�����]�#�K��6i���Q����
����O����p\W���nDTy�^N��U%�ִ��+����ɧ}������b���$5���ף&�P�Ҍ�p)�4p�P]�U)!�o�ܕ=.���Yѹde��yt$���4�p�]Z�F:�H���:����{�"�A�qx�~=�"�f��mP\�4D����(�	�wy������oQ��SӚ��ǖ5�z>��z��74�&<S�F=�{VA� AI�^��ױC��ʕ�(�7�>���&*�;mWLܵ�iPWҎ_<�n
!�j�0Β�Y�8u[�w�ӻ~?����u�~��fg��tS"Z_r��*ƞ�٢��ba�}�q�PɅ���2��P�R�B���"L��I7S㐥�Mm!D�nN��f
S/��'}<�p��Y�>@�������}}%���2O�"S��J���N.u��-�^wZ��������qm��z�#%�x!,h=r	�5x�ב���o��&*���B�h1ꮼ��绵o��b�J�9�o@��=�|��y��	cB�ӳAb��3�uo9�!��z�)��ڠ�-�����n' ڦL��#��:���T�;��=D�dk�D�Z�0�4�UjW<5Z��[�N�vl�ܟ\�iZ�!��.<,�S2��s�\nm�N
#�З���-d߲qSl)lkt�J��kml��>�L���ɒa��ϫ7E�ȯ1�79����JӔ!ǏU�	�c|���:���Ru����g,���0�]�}���׊��,��u=NV�M�\0 >'�C�+��`�FrT��~N"�J|�K�gode�E��M,� _=��d�%�X\D�w�,�r{�y#�WӤk'���Ӝ2��8e!"�)7���Σa~"^P��E<b	C.��5��qAͮ���y�*�n~W%�Oߴf�aUF��-�E�!�%�uW,q�.���Xs�i>��9B�nt�X�O.�['���	���𔇡����x���*m�gOv^I��t(2k3��`�կ��_��vf���aD��Ӵ��:���B���1E�w(��y��g���$�>VC��#�3�K1�y����g3u;W���]y�p_ywl#�k�* �Q3��+��$~CV�?̵�^�Y��5g7w}��➋�%��"�8������B��h��t\��?43�7]�Ӊjj��^!�����O�z������� �*�v�����f�f@�jX�]�n�֨�&�!l9�u��M�n��=b`O<�cYu�ږ����P"*�^5���֞ގw��zB�ǪSI�	TQq���rj����|+:9�t!)�����d0���S9م� �H�G����%P��d�=k�:y�=��
.9v��� ��H��W��v����hYy����Ru��K"��)�x�<D�y�%U�m��g~#�Enץ��-Q[��J'2�z��B�s���\Ft?j�lO'g�$d�疙 m:R��7�Ce�����no�af>-�09�oM
W�������Qi���������kzd^y>�+?�Bh��Zތr��=��]H'�������vi�j�ҕr���զkAg�u��%2˝(f�����r���Z{�N�ĺG�b��r��}�����H�$�T1��r�[�-��;��8���#��1!Ve;߰FO����2` �w73�6��!�=� �ir�0�{0��G�V�0��W"�qTa�֣X��w=��Ԫ�Jۺ��nR�CYzp�Ł���#]� ��H��yfD���0�aw���5ka����h�^V6�A>�oD+�h!��Y� tmq�L������s���)q���޴����m�z3���#ڮ��KJR3_��p�(�pJ�������UtVQ���Nk<��GX��`�a^QNh�;⽒���υ��@�'�Ptl���ED����g��͆v��^z�D��%񉡛A�s�CHބC�gIꆖ�b�@�yu�і�r�g���;d��x�#�F7G�!��4���[W�$���%�RYA`Ä����q��6��gٔ)X�nGN.kQI�j��������/B�4L4b�@Q���3�~&�:^Y�P���OmWd�.a-y�!�l�>+�$�!e�_yGo��Id{�S�aei�^L�F��GM],��W�O-K"K�+�XP=�Bޭ����
H��c�Vf��7��o^s<۶�O�O!�-�
9(�aۼ�3��A|N-��B��?_�����O����}���kw7t�I�̛Ʃ�+Ol�y���"�A���[�ٶ#)<w'711B�n���q},�<�)�Ӊ�8^�u~z��H�nb���'����w9U�۸��3��Q'9D�/e)�JL��o��L��Sۼ	�?@�KC�5�����ٮ���B�����~1��X�Mm~���<��~��Q�
_��/��ߌ��#�%ǌ3�A(�=SpHڷć����,1	���"�\Ø+j�A=mz��gQɌ���\��;[�4&��~6���^��R�6�z���N�i&{��)��t���Dx���6g^R�ꧦ�jL����i�ׇ!L�����ם�
�闇핏��_���+L�����_H`�i��!�1����(���	�:��Avl�ھ|��4]I��K �Ƽ�)������J|� e��n�>y� ��Yb59��oq�+*��]�g��޹�r�hZ�2Xp5��c�#>��ӞYA~�m�� ���o�z�ۓ~��J!XA�=6��L�ᘾm��ғ�a�M�(u�y���^,k���^��vh�o]�j���Wx=\p��R���3h>�v�$�����M���l^ �c�rd�ɫa�[�*�,9x:�V/������W��|۷�ֿ]�eP��NM�}����iw�zʶs0֨������c�h�w�Z���y����=�����C�}�.P�x肷rVY�Y��;Zݰpj�&olv���Z[��eN(=��ŻkK���o�l�G�C"u�@�X{Ҧ.��WL��VJO9*@�>�R<�rIZ��֚��mG���+���E���_
�]��ev�z��ɍO_6�/S��g���u�p(�e����A���=E�����Y{T͉�J7Ho2M90vׯ[����E�D
r��H����Gl�i�x���Z�nv��/�fF{��s�ob"�u_iq+z����	sz[Ӿ�[V�V\Nw�p������#	Uߝrc6���5F�Z�)��O�,��o�z{�c�=7��p�a樨�'�;S��������NGҺ=���*˦�C�$>��VQX�=D;���#0]�@��O��F��G�����qx6��<�u���B�r�g��=y,��>4<��߽�
^z��78Ѥ���y��(�ړs9&�����T�,��=���u6�2��Z)�u��h�	*T�m��X�,��=�:a)����$�;��6��(��T�´:�Zm�ug�� �6U�n�fi�G�&�v8Μ~��:e�4\�<}�����f�L����m����-г=x�K%}(�=H@��M`���^]9�������G��/J!gng�ˮ����J��Ck��/��hj<�Ԭ*�8`�S޻�����2��	cw.��t�?ˈ́n'g���)���he6w���%h�,���;Qk���'f��z�����\<o���'A;pV�,��B���}ň5�!��]�?-[t���V�!�4�G�P�΢C�"Y֭ ��Z�P���K���=R�< oW|�sW��3ɗ�د�U<k�˸n]�Y���+��f��O4��땶j��c���#�J1���^I	�6ݜΚ��뗪�IVn>�'6DS���P8�7_������t5���l������P��eg������x�nX�6�V�Ǽ�_N����p�����t����6\�u��ַU}=�%��U�6�gN�E{� R���1�,�j�˧i�F�:����3n=���uc�]�Ѭ*���M�yދFs�kX֠,az��f�"����D�f�g�QY@ޕ�ӓ+"��i�Z HQ�r᝛���}#��fQ����
�F�ܶ/f�����eAuvz_W4���[��En-����F9FX�uy{�H�]�.�%�������~þڋ���:u�׍�96k:*(kB�a���X�wEgnh�r�(����8��!ٯ�k4Ei��Cd]�ּ��b�2��G,@��DLS�UU{Qkb����h"j�y:*j�(
h"��4��:M�X.cL�����~�����o������~?�D�IU@RDAS1EQ�h	�J�(�**��ݤ������>>=�������ߏ�ς�K�I�M�pyTlhj�(*��@Dyj�Z���[5�L�%E#ˈ��h�)�����QD4��QPRS2S��UBUW �1LM4R��k�i墭ji���zᓫTUST�,�L}np��TTPS�:��WV���������5��Q�SALDML1\ƪ��(�)ib�b��CUT5LT��AMTO[T�$T��ա��).�k�$��Q0h�RR7�������("*�cƠ���WX5L��UT�D�CO9�QP�LT�QMQIDEUW1�
B��t�>���r��˕�6�PȣpB��S(�%�ɪ�{�z{6WJ�!Ӡwd�y(/��:�u��Ib�|-A	iv��u�q�N��4�n=����tN-Q5{���I�s��iԌ@[T�m(H`��e�O��:	���FC�F	�}Ks"��@,}����Vy޼���A�	��!+�Hl
�}j���:ZF�)��x~��돲��CZ���?۱Z)q��TC2B��S��M����b�Ԝ�S��݀��B:��u��Z{~8�8�wg�fĝ��Ϳͫ_�8^9 ū�d���ƃVl�*�ΞyE��0>'u�o6S��l���u��n�צD�lʚ�\�>�;'�,�,J��r�N8��s[�Hǻc2�Z��5u�m����%�p�n	��ߤ�W����`��D�^�BeAb�J����5�Ʒ�'�]4��]������
�C��������2��|x�6�'��Nl$�%�hv��l�j�N��7~�߳��=�D��v_s��d�f]�u��	� ��X��zx��3�V,A��;��˨��~�7�3�֜q�4)�+������ @@�Ɵ\�O�&�Y�,�豜&p�W�M��+Վ
��A��3�����W�j��i�׊��N)K�Z�����P�A�Dd�`�͵M2�ΖSw���wH�fK	����j�����ơ����"y�Lc���w�����m�^������o��qi�u�	Ϙ�
/vj��=Lޛ�Ku�F�|Z�lF�<W�U�<�\�V������3U\���`@�^6������a���oH l�l=;3�ޛ$��=�����;��91��?x\�"����ͭݹ/�ٮS/:ާ�}�����v�3 ��^�Bŗ�[ȁ���K�sSʁ��N8�⨰���d�U�Y��PY�t�ɾ�UF�ߣ0���A�X���U01���Bչ��8�,w�T����Q�D�˺����?�=~)�ɲ*�9�T���`��"8;���� >�vf뜞`��rT]o�$XzY[}��k�3����ld���{�\"0����S'{��Op
�����$�y˲yz=
��p�Ey��ٴG׍R��G<�f��'gQZ��\55�!��Y���T'i���У��ffEd4�S��y�#6A���Ey��l6�ьO)��y�+���!�c�ٽ����eW8��/F�����{kݍk��[{ �J�!�^i�v:l
b��$$���Wj�����:#X@��Hw5�sP'�f�vyH\�d��*N�x,�]J�-lX�W�mU�a֨m�:a��L��h���C�矶1��;R�x�M|�&;ֺ��;Z���Mߵ��$������p��^��/<[&�b $yux��_)���ߠ4|���N.*�25��Uܲ����W���%-��Zp�jj�j�eeyy����.4I��6���n�	˯5�Q�b��MÑp���I<3��&|Ӕd��:x�[��՞�죳;�4Y \�����땁������Q��?�D2�rA�-�L�Aa��w�~LEt{�p<ߘ�S��])�eH��l�={gO"���0��'D>P�	>�uDA�)�y�Utwf<Vq�ЁZ����I�14�*�c���<D��8��N�_��V��X1�m|=��z�DR����W��*��u.�u� �Bw���)�]/sץ��.��5��Zd$��n9�SO	fE���'�Qd�j�a!Ђʽ0->���la��$YS��9E��UzK�Ö��6���I���77w�fJʫ"�m���p��y���мQZ���E��ޑU�Ӯ�R�c�{]�����df���6{P�u��C"���p�+#(��]k%����ʄwU�R׻�Y���ݝօ=Ww�r��qL(�6ɮkL�Cܵ� ���1��~h���N;eo|��ԧ>�j�;\�� �1���)���~c��=%��M� ��O�5ك�`GTk��v�9�������9!�$^�/��A�(\�*il��ᜦ��t��g7���kK����ɰ����v���9�pB�ύ됮�>!��Ϻ��(?��~92������$b����F\�}]J����R���yZ S(�81V"MX�Q3dxl�ܪۻ:��Q<44�⾗�;&��Y�r�V�#鄯D�W�F��aO��o˳M2V��Gc��k_t}t�no~�7���cD�(��~��2$��,H�̧��VC�����2%��b-�`�,�З�z9���nf�gXu%��׽��%ˇ�+�է��w�G?�ꮙ��M,L���/߳�`�������_*�%L�7�c1O�*1n�>���a���,��Cn��\{��K=�����4��z��L�3l4�T�ld�}x�q�q�����9��ՄG6/(2e����a_���Y���Z'��BÄ^�wY���s��r7gXw���:d,�%��N(r�d^�Ji��F�'�{��ό����Ij��k�ڌ5��sK��<'f�r��萅�}�D&I��Nl%"�׊4���u�jX_�d�[���zP1��(�A�L��v'*Q>��Ȍ���Z��M��)SK۳�̪d�h{9۫i���e��[��HZ��>uo~iO�J]��(s��kĩ�N"�W7+Y^��ګ�nv7cn(�l�
��d1���xr�~�SzQ���Y�n�i*.��6*��o��Qx�Rr���ܼ�~焎 �Q(y��"��(u�6�/���<��L 
����L�!3��O���g����|UCt��)����ƕ4X23}CVs/U�9W}x���'MJ`�t�vJ;Y<w�M-����p�}}��Qp��L�����7��o���@SQ`�4C��bž$�H#-_�]}C3�o19�;C�BD9x���KDJߍO+����8�"�#5E�BZT��zH�kD}a�b��m'5���uU�3tp+�^�ls�R��7�B�,;���e�k�ӐgX��A�=B����Q#WB;Y�8L��X@�\h�:㘦��k�ȹ�GrD���6��u��"�]d)�y-U�U��������\s�Va�	��e1�J�uל8����������K,��bp��'���d8�tE���l�vD$�r�
uݬ���]x�9~O>����c�˵ܞ��gw!(j���� {q��<���ݸ����Rd�<^�;]����SJ�U�mn��ދdr;B+�:g�Ѡ���5�؄��1JQ�mH2�p6�>f�J���z��
���^��݇�*�ʓ^+��M�K�t�\أ�W��'!�QD�cs�c1uܷil׹�Zq̚�UֶmMwFP�7��������>٧�j5Wp��[�=Z�X���#&�!5D�)��Q�Z�Qe��Bu'/7�s��'�㞻�;��X�g�+�d9��!���N�~�V�/���Me�ܭb�Ģ��RAzvgX���H�J�^��hfs�#X���i��'(f��O\'r�� ��</H�tJ��0,C2� �I>��W��M��%M����R��"���F���D�뮨�w+�7Yz�DA��ξ#]���d��������f8��H�"i���9gا�17����ٻV��WIZ�q>�FB�}����E Vo'i6�ޕ�*��ҙ����'�{c��J���4����:���v64`������i:0�0�����͞����W���%n�!^�l��/�XP]���sո��`�-{�˲;ޚLM`ӫ(q�������:�h�_���\��9B؋a�p�t=�����H��XԷo)w�|�܎��/7G7uֽx���GM�0op,���y�/�%�.z��(��'�����uQRr�z��Y�Ľ�� �p�,V�ש	Bh9�74�ee�y�(f��[����E��q���,�+3^K=/��V�����J�j�φ����P�̖�X�.�\ݾ�� i0=����eG����w"7������o�|M����������Θ�9EeI��a�݃y��In�����������S�燽�ޗc�\H�I�w3؄�Z������	� �"���o�5ߦ�7?�ѶԼV	�������=�D�����{_l�]I0ۺ�,�q�T7u��X̀AW��$
1�Y�������*�/5M���Տ�$��Mov�1ݤĹ�l"�#@?GO��T#"0�]��̖��͗��&g�)��ԧ�lC�v.ji�[Zv`@�Y5.H��E�Δ��Ih����q>l�0A��z���K�HW5'�J4��<Oe$�HT+x�U��ٯwA�\C��V^���x�~�'ў]��̃S�*6z�"�6Um��z��y�bv��4��������F����T�j��{�3x��o�8b7$F��^��)�QZ�d��Q8�鉙}�{��qQ��UB��w`�}�o�Y��Fwug,���S�4��׊��gؾ��7�d����/�!�;�-�o>�����	��y�C2��;�����tʗrE�uDd�U��a���~��-P(/O`�:��w'}s�v��˩���$w��v�/1�����
�� ��#���.~��L�s�=!��v�m@��z����\����ٚi7�*��U��b�&F��kFE������xtUU���9�u�����5�F\]{)>��1�a�G�OUɰ�Q���/�V�E�R�~E[�w���z ;#�6�s>�b0������깬��mӖ)�Z��q������ù/�5���9���El��0��(�M�wSv�2��V�<+U�P�m��1#J"x��{_WgV��ϫwx��9�l��%,�~��!�]~IP��7����}4�|m߷�Y��_��+�rC(�m���%��:  �s��y5�4/�uD�H�C����ƷU͛����� dp�4��v�a���Mp:Y�u��0F_2W!��e��Yѹ}��!rk�
B����|shd����yX�æg����ۛ�7�-R��3p�}���`��@�*���NUϵ[���S�#+��ۅu5�i�)��.)�T�F�7��_�t�x=D�%!��TD��M*yl���x͝|h��R��(mn\Y���MU�� ��H=2�D�5#����F�y~�߉X�[���q>�+����yA �ᓰ_,��N��q�w�.hU)ur�F�L�{g���n#rV�0�v�@n6�|U��~U�Q"�M!��ذ�3	�������>�fGY6Q�����������{9��b�`�i�]������7����u�n;gE�Nȧn��%��{��f���2��r�5�{1�"�jh��$�����w\͒�׺��k�����{%H��xao�Ñ�"!m��lE�T�+r������i��Ӝ}|o�VM<�) ����ϡ��M3c�y[��hd-lю�u�z�Y�Ui�A2\ǫi�$-ފ��FX�a�xeo��V-1fy[��	X(�	ۿV*U��<��]�PvH��k���%h�u������u���Zro����������c<��_�fM�H��c�2G2/�U�+Ð(���gwP��Ν����쾓wc9���Tkk�s���x:(��:�m`����&V���ש;5���7��ӑ<wż��=���xź��g�mt���J��p����f�U78�8�g��2�U���!�r!G�C:[k��]��L�MCs~������r�0�9Bz��@԰�Y��[���{"��tł�tc�.�h���{4�(��� �}.[(s�\��Lg.��&��� �u�������ux^���z�B&�Q̏,�:�25,� �*�N�u�a�n�y��R�%������P6�C�ⰏvM�:
�i����F�t@i���2�fOUdc��G]�X��t���+�Hɳ'�k�\emM<]�޳]��m�[���4�'�o'6��"�l�^�)-�lBv�Z�\r��g��^�Q��x�k^���n��#�E�H\�(�;"Hí����4��"�	7�t���%q��;-T�Fd� @��J��4dM�m�H�19�����n�h�
2��W����};���
�	�%��;v0���X[��&+��_%VW<�]�w�\��3yk�^�����^��5��0�dt�t�G>��U��Z�0D�ٜ�*2��DaQ�f�0Ve�����0���a�#�#�H�4����V?�z#�Dp��������z�l~ꠥ{����a�-��{�S���6�E����h�λ�"���f!��Y�����h5��pd&���MEysQZ��J�Wo'ʇ7.G3�6��w��I�0��|Pۻ��E{=��9=�v���]�n�}-�a}�q𶨽u-�%S�'�ze��]G�U����;?-�ӝ-���r�W����`�eI���׾;�kd{b���^���������IrV����ʶ�3V7�n�M�r��λ��3h 0:��ef�9|��긲phmX�;+��\�� �W��i9=��m,���W�]�����am�!�%�(�g]��h��B�������0��ƴ%��-�jol~�]�_��#��G��È���]�� ��{N��'d
�730�<�滖�$]�WD��G�HBv"�GQ�}u�E���͍���`k����j�kvg<|G��fKM�BS��k�^�A���oQ���4 ��J����Yՙe^@n��.l�AP[4�&��s����wn�D�-䡍L�Kj11�_�]�v������T�άj�_�I��>����� �쪱hY����q�W�������F�y�ܙ)z����q3z3��d�#m^��Fhˁ7|�Y"+<�^��7x�{p���],��QE*F�.J����zN�-�V��Pkd͉�ε*w�*��ޔ���W�9�rs|yi�}��Ǯ�LU8���*wd�l���n��=���G�6��C|�.IlN��ZvdZj����{���R�l�G64U��/�+�Ϊ�*��Wg3�J�s����*N�L��t{];�2�u�������~��=��龇�,����)��"<�簧uwW�޼���N}Y3��ƛ�SRH/��u��|yk�螢sѷ��n9��=���u�4�*Wy<�y �����~#�9�}1
���Z�� �\�o-w�7ǵ�S=�E��w�i�7xx��W�݂1����u���	V�9;x�S�VS�{��.�
�8Kl�s��_N���7ȷ5�t/.�1�+ʆ�O���Y�P�Go���!�u�|�O{O�`��v��^�Y���Oޝ&��Yֹ��ޖG��s�xv%t�IŞ=�����j�c�&ϤK��{-�s�W&n��vjB˂<�c�����o��}!��@�u�,���y���
�U!F��}�c8.9O����V8}�sgzgG�gV�B��@~���L-dj�ݚ��9�/��M�S�����ͱǓJ�EZDFZ�l����Nͻݮ�v4=�Y�OC�����AWtp`O[����bƳ7��@^�g�@���}R"M���9_�pX\��t-�^4lkC�������o�u7���k^��\�hX^�rT%VއN�;�s��?��D%P$DKTQ��D�TMID�RP��UDG�i('�����?�������ߏ���{�li�4�s	���"I��QPQ�l�(+��Ǐ�����������{{{~?�	&	
ZJ�C�LMsj�Q�MD4�,Qͨ��4DD�-5�d��
����)b���TSMIU3GDy&���E�AHD]n@:1�ڗ��&������"/X4Z�5PPQ�SI3KM-QE����UM5T�1'V�N�"��(�n���ъ�:j�.mP�LT��$m�����N�4P⍍�4�I�z�K�]F����%�T��14�z�Q�����C������j��5Ai��T�.�b]T�I\�ERr(J5T�[���cU��F����Z֪�C߀ҧ�}ϮuW�h>�J����W֪I3k��eB���X6���Oq\��\Nc,Eu1�{�%>Aph�,X��mm�^�#��7g����?H�6�gg@q�*���'����"H�bܫ�l�Y��H7���^"[62 ��l��PY���J����X��c2�5k2�T��cs���u�sy.2x�W��=����g�#�b��+��e:�f�M�v|ɪ��٭�/-�f��Iǚ�Q�/�gnr@�ͩ�'��X	�	׸LE�����z��}[�/#���"@=ɪ�S�Q3�M���2�}�^�ta�PY ����Љ��Y+Q]`�	�D�a�n�&��WFmR���7��7��%��>�� �+q*2"��ݏ?F�ӵ�æ��u��p�\ib�R�GWM_�i����nM˒���E�|�����_�����
uB�$�^R���������w���W?l��|��Q��#եN����h-���s�6��������/~���5W�!R���J.����vp��Π�	`{���h�m8ߝ`���d���x��z� 5�1_Z���Go��_R,��N�L��dB�Yp;YX��7�SK<޹vu�h뜞�DR���a�:����9@�A�����bb�3bu����� T+�I
�+�-���T��wv�t��G��u�Nv�S�c[ �M��C�k�ճ{�l��+^F�:�Sneb��P��|����[6����km��� ?�r�Fwvr�R��j�S���v&\��c��ן� ��4��c!�A���b#��XGu�,�}Sݏ��ҥ�kz���Q3)����O���G�8xr�@�Q���_\���tz�Qn[�n�� ⢸�!<��H~�6������^���ݓ/�5���s܀n+S�Ը�3y��z}^��g�Fu���a�Ea����WY��;=�a��{KE�d���$o07Jy6�4廉I辌�۞�>���:�d3��r+�?$�*�нQydC��f��i�:��F�f�*���x���觛�KX�(0�GDON��'6'���j��8���πΧ���ٟ���ua]Ƽ�{��������3grP�p�M3}���<u*����������)���������g +iȊ�;x'�������,�(NTu�@�Gu�0�AJX{7c;o4Q^ɩ��e��ŋ, ݄f׼���n��?v��Of����`�o�#���8�4Q֜�R.�F�P7aHECH���|xŧ^�sv�M8,h\�J��(�
������W�n���2Y�f`ܷY�}���!l���U���@��IJ�=3㴽�+y�L�����������Z�k<p��,�*�X�|�u�5���G�Q.1f��闻Ӻ��fQ�n_�rx
�ΐ���՛��),�e82N�ګ��~�}�sg��ڻ�Y��gc�B��B��p��l�1M<S����=,�g7��$��*Y�X~��� �����[����{}�/�3�RX�#��Χ��N��d�U�(�c�+�|�{bS�q������YҠ೓e���u|=Ay���c�aq."��EIJ�/i�Y�2���Z��f9���ԅ��YSu�V�=A���r�;�~ס}��g�̑�Fn�U��y3�-G�ڎ^��,ͫoy;`1�J��sN[�+.\�9�Ȋ�n��׃���t(j�p�`��&��@�;�
Ą��N��tn,��)�6�^˄ފ���(���x�-oBO��`�d���'/ >�V��i�ŃH[y���&G5��>`����#P@�&�.��eʩ�̅X���c����̎ܥ����q��c�9�(�G3�26lIV�f��f���[:�.bN�z9���Ftd�6��s�M���; ^�_3��5ɀ�}׈�U�n���گ/�z�t���99Y��nO2(��Z�_fM��ʣ���z�M]U�{ �����+"�*��9������^�.0��zGzs���=.`c�;�<_v����䷰����6G���0�*�f�^k]tcz�ľ���x�qb7HYh��]<���$�F�t�M���I�8Y��m��Z�v�GM<M3�G�t����Z����3d蘘Y;�O��m��9��~�IF8��[�ꅃ�$7��B�C_+&�M¦U2o��]����`�����a�L�=���Y#�I��J%�������Q�ǒ��y��s�A�^P�R�s}.8(ū����)��K����\���q�s�y���A��-`a��&��ђ��c�wU14�g�c�gJ���{���>:��;�֥����5�����j�gfQ�Ly�M��8�iFa�%��0Oq1����! H��-��RhYM]|�T��~2�샳�b����~V�q�ǉ���c{�pUs�A)�.��{r�����4����:x��}y���X�Noq�sdݒ��P�*c���9��SZ�01��a�b��lf�uɜƺ�l��".�Y$�\h1�qH��x�z��bejy�������p.��.;���\0�'/���h�t<��^s�&͌���|ٵ�㳵�B�r���{#�ǎ*4�r��`F��t-���#n�3'mgl�̯U� �U�ǫ*dϸ�r8�v	�M��k��~���є�$��4�`��6�ͧ�ù��yo��0Iǘ��2��0/<��_كM�Oe�^>Rg��>�>�/�9���݋ĄO]x�#�mC���ʚ��71$�m�[u��O^�l���BP�UD�H����fC�>L�\�k���f�MX;)�j����l��8�#��@�9��/f�5��}k;s�6�[}�=L�HZql�{��Pԋc���j���pg��NӘ�FD�Xu����`�g��>�Q�=2R�F����&��خ�WxNW��G<^\;hbŃz�'َV��m
W�����=yJni�쳎B��Q�0f�}���+��{���%J߸7Մn�ׄu�����J�'7f�%�U��md7��C�2DDN�Z-ϛ���bB@�zG>��\���%%N��϶�D�1�u93��&��k��M��Q�G!�� V�)+���8�U�.����!3�"�f��nVk^p1y��8 T9]��1�ࢸ�ޓ+}ʑW�$<�<�~^��3O�7�}�W��Y!A�57�}{�p�'�U�E	�����÷�w�__�3s(������|��:l0��0X��n�Li$��-=�(C�x/��r���s�QC�������}��-�B>/�5ȼt6�A���g��5�+�}���1�e���+
�^��3��s|GW�&��B��ػ��W��n�
���H:�Vu*����|�,��9��D��\�^+��v�o&B�F�!��W�NO�vI�C�y=�1�v��	�1��*�5����R{��H����6o���M�ElB2e�f^�~��2e��oB9������Qܖ4�|^\�~� �m���)כH��VQV�X�������uE�P<n����Fz��z�rtX�J���<G��`�թ���,���7��1�ޟ>�_F�!Zw.2���)�m
����vѪ�Y՛�J���H�n$m��O,�Mv�V�DT��/�hTo�22�wB��J��M{6�/i�C���[����7y��ҽ��%hj%��X�#�-��g��[�����=y����xIA,��	�Cd�F�:ٲ���l�����ҔF�F��3/�>ړ��/�g��\>.!b䂐�:}�qP=y74��L�;���T�����`t�B�r��Z}]B��	)T���)�:�v��o'�������J��*�O���B*oG��5�5���Ne�p��s������gsL���Zn�t������j��xC����j�g�R�w�מ��WP=df=�w�!���p�~�a\�&�3ϟ�����EuVu�W�3J�/��۔)����������u��l2��:�k䋠�dc\j�*|�E�n�g���ge�7.���>r��(!6*��x͉��ٛΦ������G���Q������c�bMy^eL@QN;�X����f�}��Yj�k���E�+M�s_��������+5�&���4�[n�Vl�	$D�;&�F��>���+�B�x.�6�ދ���K�]��U��g\����R�#Ve�3���ꮧ7��R��IQ�S��;
:�6#�e�ѭ���X�q����OdV�T�Pue]�M��;��{������������o�|���������i�nK��� ����9�^n���+-�)F{��� �l�!��9�`N:���y��~�U�s9������鍜�*|8���Fz���g���������+r�l^�]�e>�uZ��^�� ��Ϧ��ſH��]eʻl9F/�K�E��:5@{��/��cٙ������pC®閚��ݪ���{�ٍ=w������.��.�D�{d�d��k݄6�����C'��V���<��31���&�uvWs��z�|J�Y�*�>�J��Ժϵ{�_��Zk�v֯7����g��i+�<�o]K�볢��e�7��*K�SsP�1ʅez�_�M���p*�������Χ��U���/��^��F����^v�y7Uދu�FR�w�w��>�,?4�-�J��!e�esg^��_��u�(���{�UQ����=4΁��'&+��K�h��6���ɩ��/�7�ۤU��JK�1ƚ��e�'2 �n!e�m���4{9D�����8��$Z>3�%+�(�n�W�vCU9̰�_��7�je:��k��!���{F��R����P���	�]�:�[ϧc�(&����F�q3��
!��#�GvB�3��OY\�)R4WuKG6���v�顲c�P:ۇ{!��9�a��kv�`�)�ٳ�4��y&��a�ּ�Fte�Q&�*�
��zO��8CHa��q.��^�S��5�(w����[no�{�=�Ou+��[o���G4��-7:�u2�C��0w_^pn;ؕg7�4.��������h�pp�Z��|W�Xٚ��:�]"=Y�A�H�z�8����S��}��GL���q�%_U���a�o���ce��3(� �M�Y1���2��tC����z�WULy옳�W�uMW�D9G�tz�S���m�#�)��S�ƞ���x(��رb ���{gf��'J��n)3�>(�<Y���c���6���X��׊���R�5�X���y{�\�ˆU'#c vö���yЇ�hp�iUL��}x�@��y}�L���,�%q�]wb�;Ҹ���t�g�O6|ɋTy^�K�M�w<�E�S�&��{��;v�g��	���[{����ޕ��2S��>����ϊ�Ɇ��74�}����?�#��f���ąj_7Ork:73���H7ZRT�J�����߯�*�/��ڴ@c�Ј��n����7-۽sf�Rz��|��x,�_���V���ڹ�d[��7��s�����e�]z�K�#cFO��
�DV�)"����q�-��s�K�~�Qٜ��>��Y Hd�Y�r��@�W��<�)ED��پ��z��i+��̞��m��bM��Å�0uЈ#�Vq�k���$H]�3��F�f���'U���[f��@�N��n���.���_.�,�X��Cp�3	��,�����e�6g��"��c�K�9=%b%��,��Xrߊn��.��>��^�ڄn�ٳ�̹݇ }iލ������V�z��Tؠ��{��M�5{#�N�f��"\j���e_�u��.E���M��C�G���o�`�WZyQdó�8:ii���|��Qj\y��b���;y��t穃B��E둴mJ��}�'�g>2!}ת�3L����6q/�����F�`l�}���)e��.j������Ɲ������%�{��r��-�)�(=�n���}�?_4,��0Q\p],������r'���;�CMūu-�G��; �e�Bt��p�����زkGU�&Ⱥ%�O�]�˲܁��a�P�GV�Je^ǫq���G�z�����=�	��7�|��w��fa��u&����"��vu;;�,�݃5f�|���%^t�$�>�l5Y�0��v��%A��?Od�L���~�Je��Ԯ�W��e6�ܟ��T��W�un���3�_j�Z�pd�:��t�x��q�+~�R��t�*�w�A�SGM�V1l
s��ױ�����.ݰ�����m�ژ���w��y��f�>�vg�n�bW-Ş��a��swX�:m99�]E7.ԋ,��3�)��4j{7��`|��2��=�oU�D��q��,���6i���c�ld�3E�o���Ö�~��Z=���<�t;\ixp���7e��k�ac ע&Dp�֓p���v)RZ���B��s��t�w���i��%�fq
qU+N/�]�}P��8ݮ�X����Xƪ�q�ާxM���;N��P��@��n�n�9��<-j�1*�T{�iq�;H���d���Ѽ�ɝ�I��Ns��M<���cBpar��j�"�G��ݭ�^{(��C|�B*z�\;qn�ꟹͣ|�m�:�m1�21afɦ��D����m��D��ڪ���=���We�8Hk!���#l�zgD�>��mfԷz{��\B3G���7�:�ޭ;]Z�B�y^V���k5dW� T=��D��؅>�w��]�]bA+f�5�T���Fy�!}w,��ܓ�t$��7��v=;��u��:T�iR`�r��m���o}��HD�|h�K=�6-�*�^U�8s�hS�I�����_��(�|D�j@/I��M�0�H>0�h���|Nj����u���!p
��3��>��{�f�k[�C�3
k�����*�$�W�o)i���(�+�yx�,��'yu�0@W�}�M}u}1�x���w�
.��$�q���vi�J��SQ�Ьa#�i�mF�ѝ���o�j��wY���c��3��r����� R|�P�EΦ�k^#33b���D0%��� RAl���=���[hۜq/'H�i�o������}��o���}�s�?��-�7f4չǄ�r3V��6�A2Ӷ
K�DIhmhjjjlo7����y�����۳DQU��#Cs���j��kQr_$��ӡ��U14�Ej٧M	�������n��l�AQ%����I�11V'AF�ӫN��m�%�m��5��@l�6��h�
�UF�n��u���-�r�TTO-Uhj�k�)Ѫ��s�sa���SF���Yɶ�yb(z�4?=p�g��J8M����"��r��MQ���li�V�*�;b*���Nڕ��*�\#��W-���͈�\��5�TQ��T1���5g�mr�rޮ\sFՊ$�5ch.��
NN%��n\�HD$� �h6RHr�p-P, \5"LB�(%�,��뮳jy\L�R���R��uë�Y=(=�׭�f�$�{�r0l\D�Z��#�u�_��q�7JdeH�)H�P¿KF�jnE��,Cz}��0A5{w�u�z���K� �����=�����$"���:���`����t�U��x�y{�:+�%��'�z�s���jn�vo@a��d�<͎�3��kTȩ�L��۲�y-�Q5�Opj��k�ϻ�9U-T�0}�	v��`I�F pJq�t1Q�?-�7g,��9\z�*%7U4[�=V�;���p4Bd0tm�~�a|�z�W�ﺨt����ى�~��7�Wݲ����=v~��Ѝ�+5��6E��,���*�j�'��gm�"�<;�����?H�gA��WFG$�ro^٪ԫ��r�ﳙ�����\Nur[Q/�E��E9�j�Dy6S�`�ǫ����N�ثÌg��l刔'��M�@���+.�l3��r񫫳'�]���wR�M��|���]gJ߳�w�0K�~x�#]�i��ޱ�&�5������+9���,m�+�}�Щ� yam]6����J���#�|6��5�z�֥g3#��$�w����w��¬������w`�u��\�{��n���/��9�l�.l��ld�����ѥ��|�b:���!\�DGv��l�W(K����Ҏe�E�k�k���^��xg���M��9�Ⱥo^�|�Y#�V#K�{̓�_^:��ko8����T�(�n��S���:B���b���ԩa��,/&�ՒOA�����y�����H>?~	��9x�P��ٻٰ��]flcq��5g��%�i-�,���T����O��Tf�#����6��+ᛓۂ����؉S�/��rע��+�B�xڍv�e��u��n�7���\c0e���R�T�W��&iP~��*}Kw���z�~�7yY�3m�WmU�]0����z$_n�z�szpc�kF�
ɦ[]w�H�dgJ�#: $d�h6Ƿ|�È�:�?Z5�"��cn�(������G3��o/K �vH�'hϺ��/K����h���V��_Wn���v���e��(�۾y��K�͘H�Z}�Eu��oeq2N��g;E�lİ�A�2-�yi�)��v����ܶt����#$�5]���
R��YDw�U����J�/UO9�|�:Pz�� sn)ϫ�тLE71b�uU��Ƨ�M�N�ڽ1����#�y�d�8�>@�i�cVl��[�����!����*����'�Ǆ�$D��9e��26.3�e^<.�ܫ�2ݹ�td@�S]��MNy�^�r9*#
��7�є���d>�<��A�ń�MUq6{!��%��Ai��CK���Zd��^[s�d҆v�Iꊉu#8�
��w�Yh�~R=��=��o{�B��t�=�9Mz��I�&��UDm䎚y��'7`B@��m�{��S��w�ù s��gG�I�8�#r�H��4H��� �i���1����V�Ȫ	xA���3a#c�"���Ƽ�;>j�.���E�u�!����[���ff>�C��#ko�V��FuP����H���ő�.�ԋ<���&�2=g�<�!wB~j��_%UesҔl��X��M�!i�/Z���޴9s�g7��-
�I(R����1��-��ep�[�s�ə��ZEa��x�܈�J{�ABŤ�HvaxnBEGe˾��2��n�٥��k�\۝����u�����g�-�Ъ�Z.�b)h?���z9gH�2{z�{�H0�;=~���ި��8���4�;��UEu[��s{��aD�-�򽎖6�w��a�X���KK^{�_F��t�-�%��&q�W0۽���OTv?\��b�60��|�����ލCv򘞻�T@pv<'��rF�.��j�����QՊ���<էb`�ݗKz�#�k tZ��yP/ܤZ��������O\+�슲1����utQ޿q~��Z��� �Y��lЊ��3[f������!B���0�MUU��X�S����e���L?��,Ǟ}P����7�"K�B2�˼��̀��k2��n��q��,	%6l�{���?�w@A({�4"c�Ιm��ɛémY�h���[ץ*���
�%O���z�_��8B��#�lU˻gj�7UU�n�����'Ǽ��I,R�)�#f�TәmMa�Mp�줿>����ќ9��H�c�:8�1�_g����)�ކ��=*���(��q�g#��Q�_,�
V�+貳�]g��4�gޓ�9�#:N����K�ַc�����,�rg�ǾK���sz��r#Z�9�wj�i5��_������Nqj��e��tU���_-
���~٣]�e���AN�]@��)06��5���[r��:�o1�-�*A�^_8b&����IYxF��Qʊ���`d�/]7�a���n��}��)� �[A[��@�
 �-��F5H|O'p����wu���u�k���ư�ɶZ��k��ozn;,�s�V��Y�7���D��Q�%8%t��f����t �d?�����g[��0�� ��޸��P�U(���~+��eq��Ά��օM�m�Wm[�������l��~��v_0�+hME	F^����W>l��טV^�-�X� � ��.+:�y�l�b�ҧ+�7CǏl�W5����:z�T��L�4��:�Un �/�z�Pc�#�aŽE>U�*1eg3���>:)t��v���X�ј�/eְ��l�2���&�$�%q,���w��9���h������'���<Pђ�2{��>��+n���`k���P��sK`�w����HV�R����h* ���q�������6�/d�Vn��_�7qt�!�Vuk{<u�&^�|o>�=�/yy������/Tr�������%�x��v
3�O��@ �u���Ag��w��;���u�n�[�ٌ�]A,BQ/W*��9��X���Ԟ��4;���/ݵF1�X�=�"T��\P]hl�m(�Nm)�eN�+zb�^܄k��p�����:��d�j�2@\B��	[�q�Xj�ca��R���ޖE����� �PF�<!w)ku�+yJO��̻ݸ�+^�����793�ڽT�i��t�Њ�z8_.����T�{���=�9�9�y��VѢ�����N�i@7��\����W_�^���������=�b�Σ���=�Wp�ϛ1���!z��k%������E^v�&3�4WGMie龂��R�i�k��J������Ɩ11�r���G�n�9DA�;��3�� ��F(� .��/��j��}�_
��1)��_�7��m[�4v�j[��I}W�[��a �{E�;M��B��.qe���!��iwvuG����NF	S5�V�;Es��RH�33�upDk�
����ܪ.
{���j��7�ڹz�Q�P�W�>o7���r	�VGW���w�Ō��sR�[��K�Sx�݀W]c�W��)��wUE�j7]ڗd�S���oC��Qٞz�6W���Yޘh[�	��啛�n�[ݴs���d�`߬<n������"�f�Q0E
�͵�4wDMvqc��M�#�t���N_���9�	�Q�J����[�n���2j�'%Fkl�24�o6���<�
2� �ʛ��s�ok}�gV��m?��a�4���ח�#x�{b�Z:��]Ɏ������q��Y��@�����F"^��#�a#�ݑ�:�XEi���B��v��LN��su[�-`Ƞ��tw�:�l�[x�w:]���5�;y�OfТ/N�֟�0c�Y�W X���������O������,��r�f��P�>�L�2h�Tv�z�<7'����ߐDR���?O90c3M��v评��5�v��6y�}�W�� m��Ы��F�=P߷�mgv��`k���~�_�z�o�[�ˮ���㗳%j�Uy����	��>�Yg�F�ؽ��<��ɭ�}��jDe��ƾݴ�uY���~������OG/����"(�ϵ���"RE���ґ�q	�2C�5]Ա���i�r�vM���D>�^�EoFlE�:E���2uۗ��VL�Š�M�%��y��ށӬ���Fح2�_���ڥq�tf�3�ξ&V�޷���4���}��D.�1��U^����hS��͢3AI9���372�i�yԨg�1�|XZ�=Mr:v]�l����M���\��'����f�i3\/%��E�w������� �tB���Zoe��m��#���O�	ۉ�w ���?S�>���q˻8�J2�l������ܰWd�w�0U^	'Ι�<4o��q���p�43�!���3���7A��7`�	3��N�n�a�͂��@�
��x��U��?Oo���v�=��W�^�i�m
��V�z�)�8c�}mQ^W_�s�ঢ়� ^~"��3�dJ ��*���HU��A��-2��(�Ru��i�݄�%��E�2i+}�=�$�[���O�eў��0rŧ�v��<o{ӏݹ�ŋ�� �毷���56��%.�éXΠX%�k��ou@5�aE{���E'$��1��Π�O�gl����g��F�J-�`��=�=�j�+���[Jɞ��wͷ��ퟀ_��nF;O~RJ͍{�"Ori�J 觏i�	�	�1C��~��~���4�_oWWlnwn�Zu���E�)�3���*�dÁ5s�[����:��9ʽ��1c�F|lɣ=��rMD���Ͷq�*�����&�C��8��9@��_.�΂�P��0�����{ꑏUJ�D鼼�T�L��C2��DV��IYxDJ���^�^��sA���/g㓥-Md!�뷮D`���'4��DI�B�*��6K<A��δ�Q*�����v�H@m�jo�,�m[��$r!��jּY](c]��9�^�
�~������|�=��>~������nc�'�kGb5��}���'㻦�HKy�����}���k~�o�,�]jz�q�Q��]\�XG�<h}����v�'eg� էV�[�}{��(>�ea�XƣG��뻜s�H�b_E҃i9GU�&�.]���z��[�[z���ѐz��sa���3ڹ�Ώ)w��-�����f0I%�1b�q�^{�+|#�  �$	��F)�e�k���m���N�����-=+����k{��4��߫�N��ÍW02Ⳟ��ݰ�����R����2�΃��nNWk�iܠnCt:����#O�g��̽E��Ec��S��Y��]�f.Oj�+[n}�6Gh�&�_;8@�Ѧ<��1+�q�e扼T�n�;p�9�����J�"8�=��%$8�~����º����Hw�]�]x�o^n���"��N*�w��o�K�KǪ�N�9�m�S�@X�*�l�V�i7/�l��U�=sJ�:�H.�4�GJ:�m$��*�f2��WU��n#���'���
�=�ό��7/����9 �+q����f6^�eR�KAk-~�W�:��"��s\*%�
r�ON4��{;#]��V�馥3�GWgv��F�g�N��YV��c�ͺ�W�������!��r���7uv�Rc�J�9L�[dc�YJ��G,��b�M���gv�����Λ(������/gB�+;q���۽)��W�e	K�{O�(���l���C�"�-ξoԩ瓒ɾQ|}v�k2n��W������o�,�-m!q���1C6fgu8M��Z���45�ܧ��L�0��k`{�*x�w�L����܃;�3�G��T=%���I���X�.|q
;���*u4��� 2m���p�Zh}f�y��~�c�}G������ճ֔��vfAg3&@��Ngv3Hl%ft:内�k]��p����ܝ@��^e���N��w�$G��Pӯ�xw�G�,���[I�7��R�������۱�%�6E�\_j�]�qIw��VY�Sġ��e��ڭR��Zt���ۺ����]j)r�XCx�s�lX��Jc��l6ib>�.���	=�=�JJ�fh��#a��c�<�`�z߭����yS��v�\*�>�l5�����Wt3���.�������ȴ��m,����}P��E'���=���0>aOM�ub(�,���ݿ��LY�#����z{��r�3:ح�J�G�S�����v��ɛ�|��"+[Y)+��Z�	��"�4�Y��a��QV�fvq3��mP���C{2�����Ir�fѼ���x�Or3�Q�p��ƒ��9K���^/���L���J�#����"�v#q��슛Ԩ}u��-�·ua��,�2�/g��f��� b6����nK����K��>�ǝaǢ��$����c9�����#V�ʰ��+pU��'�GXrV��!r�O�Z��5���Ѽ����5�k�o�7�y�|:��ٹ�ޗK�֐�oEJ�J���<��<ߍ�O?U-|9ۍ��M�	5�w�=n�b��{�C\!��������a[�bֵ���ܯǷ��E缎Tr��ȴ��Pq��>}��b�T4N֚��k�t_�5��\�-���	���{�<B?�*�d�� ڴfK�F}ݸ���SI �r7�ѝ	�lreb�R�E:m�����"ȒC������ŷ#���=����r�q��3��6�V�aĜ�d�3r�)B��]���r]��>��o�,Q��V��ZY]Y��r�Ż��t�����{b��o��l���� ���m�5��
h�i�X�̏*��(��r.�e�\Δ�AB����	��J��4���A�Q.�&�z�![i;�0𕆒7��p���:"�kt6]��-r�J�������Q[��a�p�֊�_5�}u���p#o]�Fly9��!�(�N\���6��$v\�AW��������puv>@�oF�F�}&���=�,���{�6�.֣켂n|k23=4O�!�%$�$Ȼf��(+Y�kPU��U��V,س��+\�sf�������o7����sy����HdI�����8��峳�15��`9�1jZ�b4i�~>��������}��o������E�#F��h�j���8����nm�Eh�b���r8Vڤ�]n��i����,�nIl�)���O*�\�E\Éѵj

s�5�m�s�`+#V�3���:8lV�N��sU�5b�CT��4S��:�:�5�5���SV�#��'l�Z�Z��%����8�Ȯ���r���O7.F�<�yln\nk�j&��	"&y�*�ƨ��E�hz�3Il%:Ս�#m�-V"�[cHD��V��ts/Q�(�9ǬjNmW[EV֪�h�ű�WV9�U�j4�͍�QV��mT��Y�Z���4�kG�'#��UU&��p�3Zѱ����b�5�`�j���a� ��A��s�������om�p�d8�u�KZO��#�yu''7�r��8i}�n_n���tN�Ί�~$vz�VX߿}_�4���I9��=�0�����T�Q�N�K����]S5����9� ���[��c���������)	��hO����,���[
kc��I],5R�U���'�(�a�M��WW�m��C_�����m��������4�����1��~ɾ[}��ۺ3�c�v:ֆn��t\f!g�~0�$�\��m��[�e)�J�n�Ό��(������͏!���b6�Ն��\��3����7nV�-�7��U;�y6��������d��( ���zd�8l��A����糃vmq����eP�ݕ�1���d�n��h�I�̩Po��gQ���m��H��kl}j}�:w�L�<�㢋zGS9{���񭈱Y�왼��ݦ;�q�>���<%!��W��kכ��C��F����
�[h'�����ٞtu�t^=�޼�H �+�o+��ۣ�v	cQ,��o�x1�oc��=<�8�V��v��Nn�y
��g{���{�Ԛyz����<�k�֞/�6��Fk@�^���Xr��2J�wTŹ�;>ܺX�ټj��H���Ům����0,$t^�J���(a��0���k�Ū<��ٌ�ͭ�_N�X��X_0T���mP�n��Lo�V���u�9��=c�ۅF�]�L�D��,�+�b
󹈁��v�6�`�͜�&�;w9tI�Y\�6d�3�=e��{��	�׵6i���W+&꟰]����;ޮ��T��#@���T�JF�ꭹ7�#m�殖�ᐐ�����O�X���[��������K���U�B#3P��>�5\m���5�l�{�Tc�dy����ZbS��WIU�W;�Y�7s�9��#:��U�I��g���}����ir
��>]�WG���䦵��{�׾�c��z����Nnp�t-����8#��ߩ__;�@����;+���-�9�=Y��tj�]��(>WvM�?T�yP��b�wE�����C�R�e�"a��-i�&~��h{Λ��
��E�@�MD)}yǴ,�
�Ǉ]�؞��9nǖ�����,��d���ؽh�4�4���:Fԫʝk�o���ʇ��>S;�	yS�];��.�4d^�:N�=��ET�E��v��������MR�͞��M�ą^�^�Vg���h�4���:���R���F��Nds0i{�����z�G�<?XL��0%����FrF�t�j������G1配��wF��ښ��(���$5�g|��x�T
���Hc��;�v�b��7�l��v��N�w�B��A8�hȉ�4U�Y��yo����XC��'#z��\S��Ǜ�Q�y~�k@�,��R#j�zhK�SBٳVS9��ܼ�c����'{���S�O�9��J�O)7���kg"3�5������i1��`)i�	W|i�b��m��ә��;)�	�k�˧ox]��E�Q��G!�VF���U=�v�DE���S;��x_�.1��g:��r�]�H�]̂�j��	)e�cƧ�b���s������|�����g���3 �0���ޞ0RRSFf����v�״�S{�-�r�*&!�� �yᜨ���Ɋ��W�=�׾����S�
�0{���u�M>m���������'���*䙁�X�y�ؑ���rm�ܨ��KW���Z�V�1We��3�[���0�/�tK�0�`��D���ŋ_?��������۹���j����u:����~�����_��/a�d�/o3YYٛ�c�+�"��M���-�� �n+#3��/���麫�-w��J<eP�Z���4u_�&|��O��gϳ���2�r��kc��,���>���Ҏ�M�/(��>1Fv5���i�B{�s2՗9�i/я��l��`�5-�T�<������ʐ���V�[EQ^�qbXO�����[����t���0p���B/�喩��������W_||�1�ʧ�Oj�o(�/:H��ۏ�z��g#���WXwѺ黑9�1����zε����ܦO3��>���:�k4!���xX�c{�����gi����q�K(��#{�8����;ا��^�� �T�ܹ/e���7����-���Dz���m]u�f���CJ%�^='�Uu�Gs>a�_D,R�A�YO4v��T���W{�.
�{)<b����W�����ȝnmF�]{Y�+L��w,�,K�1V5o��S�geG�2�G����=I�KҪz̻oC��a���o]J����^�J���K[�NDF�w(����,p��Ϳ6���\�$ؚRk��(u!��ml�YI�cV��/Df��ݖ��4�%����ɸ|����9 ����d:ꉑ�dms�nߑ�5��gӗa9�*���d>R���/�W^s1Q9K��v���l��nQ���ג[�Q��7��unB�ƀe:�⥛e�̂�M����{tpXs'���ĩ=�QUA��uө\l��r�Zꉞ�G�"�6�3�l�q<�Is.;�0G@u z̶c�۞�Զq�v�w2����r((�i�ۭ���4ZJ��r�'՚����^nƷ~����"z��rq�B�t0�.��7�D-�F���"�k���BA�P�o9_p����<��>�\p̀�s.7�O�{b�'�?���)�l<�^S�aҡT䁴����L�����J�o���Յ�̔0Y�Bݽ�dyFHn�j�
NI��-Wc��u�f8��jD�S�(�7�͏KH���:w-����E�������G��g�ڛ��_e(-�#B�̝WFN�a7�/I)���$���[��s\�7kE�\����ъA}��'�d��,ug.�s����۾��p]�]����cG8�oM�e-�P�Q97�p;�m��:A�2:��bQ�X�PM�6�r�W�&h�Iu�x�;5!�;e�vȸ���i��m;�=�'��y��2��y殣I~�����^��_[�)y��63Lf��3�R!��E�i�k�Ǝ�<�3�ݶ�b��1m�N���Q�8�]^�������GL&n�Px�9f�N�Ъ���sp�*�Ϋu>�g�xz�����0��������W|e�{s{�;@�A�&�]�zl50��X@gq~���d�L�:���}�����ǯ����9�Y\��lɮ4㕮��4�馥Z�aCߚUd3�vv����]0H�+P��v)^�
JLq��U�q;U���x��ךB��v�ڈ�2�2}(�"��ٰ��t���<y�$PAý�m�ܭ��w�P��]0����e�V�?Z�16;Sһ �sv�i	7k/J5p�7�s_\f���&�G'����f����2%o3KWrθnm�;r���ta�J�f'��#M>Ğ��J{Ŷ���+�W�=��$�km�X�Y�OQ%Nm�aɲ�U&"Hx���1��3+��Ct����t� �:+�U_��(<�'lZ�j�N��ilv�{��XF��y�A��1�it
Ș�aua��Q�ɝ�����1Y׼�^��J�����S���L5�,mY�8^���2�F�7�8��3|ni��yP��b���`�m�pFm�:-��kUT^m�V,`�s���k�}�ym��r����n���{o'UΚݖ��	�HV�s77�s����v�oe���S�v*��\C�7���K�wH�WHe�P8 Z0"ϗ�(�k�F�tq�s����`5Dĥ+#VVs<�q3�(ͫu=�E�uE�њ�
.�.� 3f�ůTr�g<�"�{�W�QɑiE@�3e���Y���ՃӴ��ԬT�=Ou��޻���\��y�D����{�H��>P�@�3�ާ��=����vU��u&����`�o�&l�ۑE&���M˸�g�h�o�'�e�ޱ������� }����>;O�;��r�B��M]����;F�cu���جR��L�\���ޝy�^G�M�(�T8��0��71bљ�Y�;^D��~���7Pw�yn(�2Wc^J�sNr<�7aw(�V��M�p��4S	vl:�+� K%�g ��^Ғ��J�=��^
l�m���*�V�19�9��r�P�Eh�v�M�ǉQ���9�S�>i��F*ᫎ�t�s�zY�쁺�V���4ϵ{-�4�:���	@���3�T���9Q6�6Wo	�'3���g��v{����r�����<���lH��Å�^l�_n��ᄴd��(�h�-.�=ey��ڸ b��LN.ͣ=,,]:����ŧ�>t�Q3฿#[:�*FUa��5�z��+%�r���FwOg���,�㻠ڎLy�n�i��\4�(C�WU�y�	����
m���}�8���+(��E�r�����۽��n{��ƚ��z|�K4A�=!���02�O�zVqnl�ó��(Q�ufɷV��Im����ݭ���]j���co���6����_E�����]�{�C�w[��k�e��.%=�|�U������vl����@Y�����bv�wuf�+���������X�N]/+MǛ5�2�A�p��
�r�<Tē�LZ����2�f���ֳ��%�`P����9��[l�U{�;��+~]�ا{�u��\B����s� v���PmfC��y�,*Ό�ݯ�g�;�Kr$�����r�ϿbstCf�}�N��;�2)Km�H̈��x�խvSX(�ʀ�QW&�*�sI��X��K���[0'%��CO_k>�1�ג�K>� ��o�=={x�!ֆ�K��c��^�*�Q%�f��|�_��[Ut��g���6�s!N�6Lj(7c�u~���Y��)���D���sŮ5���r��EO�GnxZ�Ab�F�Du5��mY"��{��r���*��L��Ժ�E�o�8Z�����ro-?m�kEA�	3δ���J�EN�6:�ԁ��n!:������F6��%��c`N�9���R�9��vq�~���yݤ�.GV���,P�쪿f^��x*�/Sk����W]����n�u��q��uj[l�Z�#/��[��Zq_]�]��{�34s��⼼u�������s�H�عR����]�"6��ޫ���#D���#WQ������U.�WֹNcҽ����!p��"8mk������TP�K���T@��1�������ȣ��o��S�[�0�цz@�[ F��z�L��<�'u�0�ؙ���w1�y�*j���g�k��o�Pu�DF)�'�,��M�m�[��w.�o^�_�;�$�
�6Xg���C� �|��t�8���5�2�)�^�g��rx��]A����=�;9#$m�w�*c��qtg5V��`�!�$�f
ӓ��|��]5ɺ��t�v��aAˈ���god�p��;��>�Y���������J���/���g���J��¶�?� g�N�}H�ϦX�W�UӨaM�y�x޾y�s�����ۓ�3�s��x���ngo����S�]�Q5uB�;��fb�K�+:�5{��<6A5�6񋉩����L�F)��_��7�}���#� *���:""���_��"" ���p�S���
��}`p�0��C*�*�ʰ�0@�0��(C�2��C ʰ2! Cʰ��2 C
�
ʰ2�+(C*��2��C � C�0�C�0!�C
��2��C"�0�(C�� ���0�0�0�� � ���� ���0�0�0�0�0���0�0�0��00�20,0�202,0�0�������2��ϡ�� !� !�" a� !� !� !� !�@!� !�T̢q�����(��p C C
 C  C �C( C �C C( C" l�� �P �T � �A � �D �dePas�r`@d`P	��@!�Q���e ��U�fAff���0��0)4���Ȥ�
L
M2�s��0��4�7�@�(ʰ�2�2!�U�P!�a�a �!�eXaC�w��_Pc���TUEY�D 0,X������~���@�����W���@���>7���X����?��u����?�(���������?p(�+�TUEb�?�@������'�����8��+�O�������}q 7�_�Oa�_��'}�O��~+�aQU"A��B � * B�  D�2 B��  @B �  �( K" B� �2�(��H2��J�B�"��J� @B $�D+, L P P�H�\?@���o���R� �@(P�>����?������@��{��x
�+����o����~��؟��:��������~�ETW�~(R�~I�QUEETW���H�?C�*����<�*�+��_�0>���C�\�A�����?P��?s�p��QU�?����*����Ҁ��>��a�����z�����}�'����!�p
�+������ETW������)?5�~��t~`X<O������^����̞GҢ�+���!��d��{���^���'������>�0}��@��������~�����~i���e5�c��P/�ݘ ?�s2}p#��χ�JQ
�B� ��A@��!�����BUR"�J�RQ P�J����T�JJUT��BJ�I%P��.�J�6�!C٧@1�$��D�Yb�R���R��[2�m�	J��u��B�ųZ�P����U�N�U�
��ED�d*Z�J�GwsMI@��UD��P�k��%�4����"����D��DU-j��EE	B����$�!�  L�'�;gN�å���5˵�k��5��p��ų�� s���'C4�k�ڦtu5�C��B�ն��ʻ���iձ���]!N䤪�"P��"�T�   a��CFFF�P��+�]�dKR6��V�(z���aE��x��Cl^Ǹ����9:�k��e[�˝h4�Q���gr��Gq�V�Z�C9��E�@�wG[��[&����)��J�UE(��/   ǀP�k�n�wZ:u�vуr��k��m�4ӹ����S�a7v�뻷u�jWvn��)��wwD.�eWk-s*�J��9gX���k�Q	P��!iJXo   ��ZHҝ]���ͻ�v�Ѯ��J���e��)�N����*�F���)��wt@v�aY�jn�����ΦQ�[�Q%H$GX�)I-�x  �t݀p����9���R��]�����kh���:'w,K�uvl�ږ��6�v��� ��v�MV*��UP���  {��k���wA][�590X]����pª�l�i]��k�ݶe�wG�.��%�Pn�qu�D��mH	B���Rl�D� 7�R�V�ۂ�ATfW,�r���V�\�5���q�U	+r�m�t��+���
N�9)T�(�]�m��t锪�h)6¨�Ƶ�����蠥�j�T nJ㔤�ha�p��tY�) �͹B�R�� ��;��4��V�)@���%	]�+�jd�V�i�V�U-(�x �	QAr��(%(�v���4��������JET'k�ܪ��Ҋ���H��%u��u)PDc� ����6` � �x����RI보RE�WP�tM�Jk��J�A��̢���4�RR��mt��]�Tݪ� W-%u:��*)Ex)���R4#MhE=�	)*SM ��`!�&�O��E ��{M��i  OU"5U@  �O�������c��J���k����/��Z]��P�������g�A��> |>}���3��֫Z�m�m���ۭV���v�Z���5�ֶͶ���ׯן��_����jܯ��Ub���h�-�z��*]�lY��wp��\!�c���PXj�;�a�
a�u�[LZ����!�f�԰�2��j�[,M�;R������w46�{�U�̱��͹��Ơ���ɧN�2�V�<Nc!jĒ4"�4�,,�H�ovś�'�(�����Z����2�9����A.إW��6��U��;��؀ݑI2�
Qe�ˤV!WSf���R��0U��+�M���
���Sr��6J̦]nޒ1ܚt �J��ȥ�("��̶�`se�˭,��N�],�R������Ĉ�[c&S؈����t� ����!kW�xp1�ʔ������{����
��e�Z���P,Å#f��b�h�bU��ߦ`2�S
W�Y�E� ]�����LfH@Y
�M%���i�V�`0nqn\ܒ�cYX���.��!�%`����ۂ��x݈�=�ö�1ؼ��5AGX���܁@���#��)��0d���#�7�v�D��4�-n�[��
(Ys��,a��ҫڻYta�Y.�;��Ϯ�EK�r4.��Ƒ�+^�ºV�(en�s�ߕ+�L�q�j�*�f�Krkx�p���jڢ�ݛ����-�*�hʒ䛒�u����4��5�����#a���ϒ�mS[�婭LY2�ߓ�-L 1
	;�Ŗ�@,AA�iİZ��Niٶ
��w�B��)i�&�"�Ьjm2*i��u3U�#`,"����W�L$�Q4&f�լ��	��-iP96���)cmL��[Bœ�@mi�pb4ph�J��aj��Z`�w6���6?��9M�k�eڹV�)��-�)L����e�Yy�N�ܽ��G�j8�[��l����^�����$岫5��@n�.�X궶���
���i�4���6�JD⊕�-�l���`=
�+z� �(�XL����ʔ��Wyu(V��d�^=�ڈaR<@M
����Oܙ�WMnVˎ�?<�x�U�
�k@v��� �FGz2��x�YR�X��a�A�O�x5#X�#�r�Й#I�6�۬�a7%ܢ����)m��ܨ�f�a�:]i1�"��P�ZB�E兂EqR�u��r�� ܻ�c���-U�6���n���Y ����u$�,*�x�"�P��{�#�5Tú.�If���Ϙ2չJ�s
sf�kj�T����<ӥD݀UC�u�����j�m���Go���`�5�p�0�uZ�6�Ռ�d�l-t,�A^��v�Və�Iqkl]0���71�4��(��$T��ՖK�N��0�߳�*�S(�I���ԓoR��r�7�����ЩѷYm5�Q,6�a������d|��+HL1��	*RĘ@FL$b3KU��2��H5{Vi8��;��΁�jS;N�j�{D$��DH
��.�6Ml֫�>rV2rc����C)�u7[���B��D�̫�-c��r,iTn���wZ)f
���7Z�t�ݠ�-���Cv�k7*΅>�eE��MBNY���t�j�Ŕ�n�Ũ�q/F�h[0%�d�[BC�Fe'd/�J�خ�(���Q	�X��چ1�t74�
A�Z6�ګ�T�q����K׹U �Yr��J�'#�(.;w�-ZcI�-�b�CSoH6����fF�'�R����m�^1�	(-��Tj3c	8k+.V��F��Z��SZ��C\fȖsmm���Ǯ�ώհsI�v�EVɫU�h�&.KȰ��@�i���lZ������Էi uS �dsm���;FJ�ҕ�K�w���1L<�3/
�Tq�s:Z���s7J��F��UA+��K�YF�Z��$kd�H��wy� �mn^��i�T�R�on��YQ^6��t��e���Ǡ��vv����^�IY��8�I� җ��0%��l�n���z��XZR���Qj+H-w)Pݱ�%�Y��/k��(5^|0��5$�yK��1���אI��N��6-��t��6v��6�N���ܸB�{bm�Su8�-UXrЖt d��Cd��H�N]=r4�K0Ա%ѻ� :�,��0��qR��5�P�EH�ЪQot�H�/N�5����)�P:E]7��e⫠�a^R EYL<��F�;�
����fE�mj��H��[jL{yj��TQ�{��*鏞]_�}��K�[{ziC�NH44B������}�6�ʃ$�u*㊊M�B���8�V�@�%K��'�A;s-�iH�M���2[xE�M�,z�c]����l�:u�4ԖY��ƹK�J��y��ðF�dr��e�%�w4C
�`FigA��D�J"�DLB��B��4Xʚq�b��i�� U�����n�x���E�jGM'�ڇL�2�5�ĭ�\f�+Cͨ.�qg���n<S6�L�����G]u������1*��A�Ұ��V�l��B�������ъ��s�wlLR��ۄ��S	^�d%�f�XC�r��'�n��tU@p+���Q��L�/VYaot�.�K1T��ۼuj��i�A�m�{b�)VЈ��me�j�b��m*t݈ɶhĄ#���,Y�����Jr��G���9� �Àɱ�Ċ���;��6Ɉ`זK���Ś��;�����F�*�K9I�QIbZ�&�{heǮ��%Cb}l��4��sq���a)E����l���t��,Ҳ�K_E��ܧV �YW{�q��oB����{mL���3Q�R��iS3u9X����1T[a�7q�mbxͻ�x<�Z�#�o
A�0�qX�x�����>�ˡ��8�����ьk���v��-3��Zt`��p�bM�@��l��*XV��Q <�7$Bٽ��	�$��+^3]�),�vP0*f�V���U�ܦ3d�F��# fZ�����8�U����i�;�\��q��s%�ޡ�-�4��T��jڭq�r蜭�Ӕw*����QX4Vr��R��YFjY(f9�RU�^ �Tұf*3#lX�N�7zdzTeT���V��^��ʊ���h�@��d{�q�/%ݥ��s[t6!��a��6Z�3-8Q�ʈSX�V�ǲ�q�y�*N�<T񸴴R�su��r�̗W�T��t��$ҩ��37�v0J�f�r��ĸ�f���x"2ҩDȝe�6�5�u���R�څB�=7�R�B���e���8��W�u�2Z{�4�^b�+�
�JW	�m����� ��ޥ��sb�B��i��L�ndؕ]Ț��l�l3�U�.���[+v�%��T�]��0���:�Mi���1JS 5c2Xy��wf��R��l�o.���t�[ve���m�+5z.`�Mb�F1��Z�����6*�[�1�� EՋ)�¢�ɩ轧�O�z)
�wnȺZ�E���!"1M����w�*�����3.���%"ɰS"\��D�F��kU�m��f���6��A�m+n�P��r�wX^M�{uz习Ţ�+K%��Չ�[��j�2TF�ʹZ7-�@��I�a�8j��CY�B��W7ik�l-�{%U��طhk����d䔫A�����L��d/$Y���*2�d��5��S�̼P9V�{f��L�nFe�Z��q0�:N����P,����;���7��� �o/.]���XܗܭM��KV
L*���)�&V`p$[��!ue���.����SK0VR�ɢ�7�K��a�"u�E<���O.�E��ɭ�n@�EW�0̏>���{E����|�e�@��;�O�t8��Y��l`���c��/6����2�ZnV�D5�ۖ��-$�6彲�5h;;��N�9d*��JƑ�֤T���#2ڼk�#jjCf�A�WN�/sobm�%+��^�1����3l�Ȇ���)8S����AbӼ �e�u�f�4�2�7.�%"��V쫩J���!�����$�wp�	�,mjZ�Z���SF�+r�����/5`n��ܻh۸��6�lQ�5N�y)���Qr�	�U�a��iV*�,��Jg�w��b�f�E��ӣZ
�)J!,׏j��mBm�cF���KoAJ��sv����,EDD*��@\���&@V]"(t�a�����ʒa��5���eܖb�b���XAou`'�ڛ�In�k,��Y[��VD���T����F��e�e�N報�bm��ɕ1�Y0�"�ɐaӖ��!���E�m�n3��*ٯ�baC(U��:EG���HQ�*6m
-�f�Bhk��Y����.��D�G�yrj�čBّ�O!�Z�HV��Ju��K*l6�^f���9���c �TN����k��L�Z�Q���j!e,�L	{ME2�K]�[�쵇תu�mIM}��jK�2�pQ;V���k�F�nn����Qi� ��F��(�O+s�r�'X&��n�`nn�HՇiq�3D5Q��Fܥ�a�^��)h�R���=yV��pJ��:�qm�z�ٳ��nÁc�U�ǀVQƳuc��ոn;	�X�0���P���7�IT����m
݈+0��n�'B�PF载n�l�)�ތT&m��͋3>�vbK7(6��6��Li�4��KCN J�h�rW$�����97��ȲLH5���b�C%[.��E:�,��u��*m7l�*�#_��<Ǫ�R;W{�'�*\�l滼��bM-�L�����T5Uύ�Z�n��x�(�Y��
�8�'�o-�r�Q�AAb��Y�gE�x����
	+`�V&�6ΑOu���~)(�3\�y��OscC.��;�)7
��r���RM���b�.s"��%�6;�e�@�A`��ۻ?8�Sr�Yj�H�6u�'$���V��c�k�A�_����mSh,ʹ��5�hm�Gh�F�%<lU�XM^3�ȩkQZuiF���v����nQ�ܻ=�KK�㻢��$��[�P�]je�q�"i/v�w(D$����;t��sN�w��.2j��(���x�Վ��J9V�׺�5r1jM��n�����-t��ݩ�&9s`�� ]^^C�� �pܔM�AQ�"TB��T�%3o��v;-�ӫ�F;W2�s�H�%˽6*�!&dCFC
�s�SJ�pd����Vּ���+X:��h�cɐ�o1�©w	�\j�t�S�+�G6+�;b�`^�T� &;Ҧ=$����5vԷ&&��d)�o7\/i���6�n�4��dn���n��̊�w��ն-�ܶڥ��(��Du]��6�a����6��qM�c�[���$5�v쬭mcc�5sAA���4�[[V�1�ы4�e����f�Or]�!PoY)��#°iԈћ6n"�$�Nk�KUlá�@&�^bH��p�ܹ,-y)%ᳰ�6�/E� �20	75�8@�/3	*lF�(ՇKn'B)Ffc"�V�Ò#tM'�>��1�Y�
$�^!�� ��m��n<�c�M���7Z��X��й�������r=�Z����x^I�%��T��n��9�Զktf�*Cj6�*�ȝ�������!��@ӂ�e֬t��[��^��VD��c���qШF\�e���l�,�2Fmsb�M�r�c�N��M'��[f�e\2�H�ͱK"�Z��&�;33�0�@Sn��i�.�$�s4�@VR�A�6����>l��`�����&`B��0f�,���I�@�;W�L��hX�H�N2��h��ȭ�{���opV\s�e$jE9���Y��,�3U�,�m�i�4�]��nP���TrF�6�b� m�8���v޼2-���Գ
�T�i�F��]7ZՄE۽�&�,ֶ��	BGp:۶t�J��`ټ�),�/VUʷ��lᔷ�*ᡘdt(k����X&×�K5�M�Q�V!�5ƒ��5�+A'N�f�|.�,[�2)��
�0m$PGv,�M�[{�<�Xt�D�6.���B��2]m�vҵ�*<E<dQ�X6N�ֆ�Z�0��Jѡc6�f�m(�����IjOB�\�2�՜���r2�d��K��\×>�&�-�v�E2�E����TdM�*"���.%=t"a=��r��$�"�aۼR��Nd%�XS�i��aR�j��V�Պ��hT�EOu��v�����R�.X��T���q�	)�o��3q۫$�{�C�����Zr���Z�&��h�t 81Œ'�dl,�)��K{�a�0���[�w���c���rTKpv�Gv�,L.=���3�6�B���r��;*8Lװ��!����ڙ[
�2CJmX���gk#(�Ępڦ�(���G��2��Q��*��$]��>(��&�शMM�2�L��K��"P[�1��ɀ]�Ry����F���M&���EA�5Dܠ�K7��1��ѭЩOTx����`�3lq�kv�I�h�.�d��d�c �J���uz�G���a%ݨ�&��J�!�VmA�JaE����#]�,Rµ��y`:V��Cl�\z*�Ā��i��J������.�!uզ��w1�Ʃ'��I' ����V���L�Y���LW�����݇p��cKyL�r̆��8�@+b.�歽�kA��Sq+�Gs0�J���:vɩ�YD�I+XX�T,�(d{Xɭh1a
0Yv����3q$����V2�h�Hj}���V���	Ķ�XҘ��w�I�tc�n�)��I�l�hk�Z�؈X5�yh�X`�2ٵB���˘�5���f1jd�����*� r�&����7
�	R��S����ҍޥC9�)����B��K�*�W[34̈��]���4�vVb�|a��}�]gRVh@�:�®�J�[;�Ѯ�zw����/)�*��N�i�>�{8����o��=�"w9�5�KWb3q�R��*�]f2@�ݫR9����� GC��H��j���m�偒���V5�򜳖�V�R��Hک���F��8�߲�t�	w�'����re6\.��bk�ȑ��p�\aQ�{.����c.ʬbM��֥wNĵU��>��bG�53���]k_[�P�һw����I�2�i�c������W 7�e�qG��Ʒ��3�hl�A�����|4	\0<��7vn�\	b�S%h�j}ܨ-]W|IC��;v�� ^ap'S�8欝��G�&%Z���嵁m��k����x�nc�f讻=%�풩?�u5�n�W��h���m[�a&���g-T�R}�i4�R�����($���D5�kA��`�9�J/qSjd(9+.��e2�-�g*P����]�VA���S�is�'��&�w#�2�< ���u��V�\���J�_f@;����6=j�=\O&x5N�]u����s+ѷ���,/d���f����y�����݉՗�l͡��BŒ���~�;�%� dѮLLB�.9��Q��jK.\Vl��s���칊�ގ�E������0VV!�qR�o`'>귴�c�V��s2��6 �-v@iu�zK7�u�˥ãa�9�|�i���[砛Ư�2lg:9�^r�ȵ���ߴ�&�U���Hc�oD�Cˢ��6!��5�b���k��=O���x+{o:hJ� r�Ma��Z{v	�.��H���RDo`S!��[[[�tzu��ʕ�ۻ�+FVӖ�+�"����_u[�-*B��Jv�4�VÑ=�����=s��K���Xx���*b�xnY�aWpQj���z��Q:K�n�x�94:%鰞9��nL�T}��x��!U�%Rv�$�����#H�0 Q��w�����1 ��2+2�յ��#A�hmǃ�p�^-�4�yJ����P���޸V�3�����֙�D�;z�^��'Gtftų�]=Ԯ�8���ңx�k��cd�����U�cRޝ��M]N�O+f�9h3��y�&��mwP��Y=i]_e��n�{�;K��� �,��M�:��p�ڕqrִ������w
��T����V�&?i勳��lYd�
��{)m��u�f�c*����
���՞�R�eocb9������'��YF�� 'Wm�F�<��ͯ��yɂU4�k���Kָ��J�����v|>c;��\��޴(e�N�v�(����+��JLQ�,�Z �R�����Z,d�{P[]]q�����ح�l(\d|6g7��ݺ{V�P�����h�ۃ�q�-}׍��OpZ��v.S+�UXb����,ڙx*p�C	�S�X؊��f��6�ݚ%�P��9��βZ��me���\�-�\�2 %�C a�ӱ��o���ˍ]��vB�,
�c&��p��^���A�Z���at�2j	�@��
������y�խɌ��z�`���}j���0WV�N����Ѧ�� >���y[V��2�.�͍�C�E#>��n�|^r��ǚp��nը�ID�R��K�{�!��>�ރd�B���
(�v�ұ��M�m켄K���륩��z%9�畔�˗�i��䬧gt[�#m��q�Y��K�F/yV?3�~�|�`ܽp�\���b��-���OK�2آ)��� ޕzX��K�8���Ʋ;�;w��|�3�ŀM���5�K��dm.ۚve�p�ZW�W
��Y9�h��]vE��j,t�O �ܷ)k@V�6�m\�r{,l�uv�N
���u�-˚\�Oi.Qֳ-wr -:��%���+�zh�Q��7�m�t��Z�e&�.�9u|�{s%�JWrf�N"A�w��N��U�[`� ������BF llz�a���-gls�g#�]V#�]ŜDuıb����j)�ۉc�k����V^�/"���%�,Nu�×�鉻r�#�o^�ټ�ա�|���;�b�Ї_�5�Љ|���V ul�ʆqk��\P6s-k�y�s�Rܦ^'�}�Q)P}�1��]v>x]�PV8�[�g3��I�tբc�9���r�f�k�3�eL�v��5:1V��M�Un��ڵ΄�Kx8Y�bs%���9��Vvy�F8å�'eN��Tr�.�%b�4mwj��b�����WF5�eaה��i��V3�T�n�����_f�r�l��չ��>v���v�4;�
幕a��}L�R�R�$��ɞMZ��yl\�!w0��]���B%��v�댘��Vf�MsI��I�>.�]<χu1kc�y�CNf��z�_yTJ�w����Fg0L�x���5t�/k�LsVc����k��r6�f��(�Xq۝�Tjq���,��5PIH�g_��r�n���v�3���,���,=zI��5���2!�FҾܷBQ����,�7;oo	���ܝ�mF팵�/�m1D�(��v��f��Z7�PG�j�o^'����,�j������:^�:���� ��iO1ܛ��Tk-t����5���M�������.�]�T�C���˱�WM�e��^6���m��PW�9 �w`�8P���ɴ�U�I�Wt����xd��6$$FQ�GL�]��k,v���ҳF:W���j]�TJ�\�A�Y������[�<��U��(��Z�0I�����jm���OyX�]E��oGZY˦1�髻���V�.P�ʹ����;C���c�a�ďib<kX[hκg3^��]��iWe2x��ǪGjٽb��cq��Y�I��X�%�z�ٷ���SiQe�3h$���C��so���d��m���aӇA����퇻i�5��ռ.u���
҄��"+��廷�J�[P��NoO�"����*~2�yJ=���,{*�E� A�Hە��'r����_I���8C���i��P�ʱ>��Y�;F�>fQ5�N�K6�g-��9�T5��@ţ��� ����>��0^˕�Z�XOy����������o��{���N��X���T�C�Z�\H-��d[�/opl�: �-�f�;So%�Бdt���b�K�Wpma!V.��q���r�kx�pF�=�W}�6���ƟֻX�jT�]JY��:�Xp��wa�<xe���\3�q;.��0�!m��F�G'��Hp;�0h7����o��ۋ��vV&����+>t�p�*�n	�CVr�@���̹��$[�YI�yc)�F�ڛ��|��]��HXd�¾�:t̄�H���x �{F�����G\K���9{¥U����0�^��L���4Ȉ�Ȕaᮻ��wԷ�M�i8P3�Re�o����;���ǔ�L`��;�A˦��ӶU�#��O�S$���Վ5Ch��s,�e"�9����\�C�}��.U��z��U������� ���[hr��<]	w���L�rd�x�����tѼ�38$�_,%xS�^n8�K�b�Ϡ4
;qZ�S�uť��M��;tI�*Ա�ܼ"ɭ��ym{���\�y�y�^Na�pZ�������+�3j�T�{�hm+h5�c�i�7������V�y��$Ut�/�u`�Q��|6��'���W�S昳J�ʐ�%��u9�HF��$����M�l���[��GCϳ�8yZ��B�����ni�����#��˕u��Cr��(@��Kq6���w*��ilb[����u�"�x��3�YC�[�d3\��]�{�ǪX&����L���/��Oz��)P�r�[���BJ�W�E�_Q�6f�:2��ĸU�\7(gwr�����릡�t�"Ӈx-�m#W�р؇w��;F3�-�t5 �G�'�k�{���em�n��7�[�َ��Ҍm$.r��ٮ[|Ň��"��f�a�R�)=뛷\�G�
�X1�)x����[ԫ\��:�mjߦ�bc,<[3K-0�r�@T&�V����ݮ��ɋK��]�+)j]&B�Z�|�-$n껾�Eu�:;�3�:,�b�owV۫�����
���4)�^K��TY��U��t�U��&Y�7s�H���<��b'�T�b�o�a-�im3�S$�6�̲uWrg5ݘ�9i1�8��]-\v�xg=gF_D���`b�f����m�(<�_�gK*��0�W23F�d�,ѹ��{���w�84�]Z�z����ec���ʕ0-�Z@�Z;����B��;��м2g��b�Ә�}��g^^��L{��|���٠o\�������{s�NqBh�i�a�L����b�in��Rs�n{W��:-9ש's��!j嫺���\��;�%�'rׇL?^��z�b�#yX�n�v����P�9���)�b3F��u��&.��r�i*���-���\�\��_K�ls�wHK`P����~�ݔb��d�-2�)�╼#�}��)�;��au�˛/F3����@����έ�);���hK��WX��i�4��������9�Bgk����\s��r���8w;Z�1����|ef�)��.��Px��HJ[v�	�ّ���j^9'c��֧zr��.;����!Bg�À͗�d�(���ȂvA����N�O�)��Hr�p�ho]�oJ�}xe[�9��^T�%:�,P�y�<[���=��+sx�����3,c&���u7�.��)�Cv��"sB.Rb���蚲��v�h�������v��sE��ga@�
鑈�����J᠚7�m�B��(�w���)3���b�
���f�o 1�&�� Z����f��\�
R#fk.m�5ڻ%^5�)�;3^^sȞl��<S8sMJU��R�b�Ç5ܻ8���۝�
o�u�� gmc^�g���kj�Ռ���w'Wv��P���ie���U&������Q�-s�v]�K����U��P2�i;Z�w����J�zQ�5i�P�[r��y:�vd �gq�k�(�U�����u�ίhg1��]���+]n
MZ�w���ʦ�AZ�\��)գ�P�^��`����ٺ���� �PZJ�̱2�x�l|�U�j�M���cRr}��.�B�&�}������3�s~F�7:�y��;\�ƴ<\�M5#�ì<��y����s���M������+�v�0R���w�<�U�LR��B2�&U@g,�}\wQ=�;�+C��04���x�;�/z�A5Hk�M,�b-�43\��H几�.r���mw{-)v��x�WUԻ[��d�{8pΓ7x�W�chi�tAALVE��a��Lp�CX�1`�d˽��|�jOu�0��Q1�.�Љ�{��2Dn�WN<��}���K�sW.*��1�a���]XYS�jU�k
8�ЗV�ҿ����%o,R�Ƀ����t��FE�]�g_Yj�����޽0��2����2^r�_<8J��u�̬�A�{� ���m^C���������o�6�>����Y�������ϩ;[,��TZ��"`�@ii>��P�٧��nT����[w�n�9��w2c�̺P+=-��DT5�l���3�Y��x���-!�!ϕ�PL�����(�p���pY�x�
�2t��::ȲH��N�v�W��58���S��7l#��)�����q�Pe��٪7}���#� ��ysl���赇[�ͻ��ےW4m73E^,4/�on�h�8bs��LP�vE�]�L��ЈoJ�ߐx����fm��vM�-�����mhmǐ����&��xi`��\�L�1-��J� 㶤qC��>+U���6�>��Wl��Lq�� -�
����)�[;F����S��3���I�]��RU��o,{���^֋t���Y��p��Cj�l	R�Dw;��T�m�i�-� 2���
����o)4����I��DI`�]Ac5�X�]��)v��qGx��{��\l�V9�	Ω.R�kC.իH+��PE�F���@���:�pM�Ql��:A�/z���S���g��+c�)���<��q�;U�X��W8ԅɒ�.ۘ�ڴ�k��J�]�#�5���v@ɽ���ʆ�']f�i�^Z[�������*ʱ�Y�{\@�,�'Ӫ� \��
����i���i�-V�
}�=]�����::f!�p�n�n]���Y�T�ڬf�r��x(c�4
0y6��b�U5 ���FPǥn��%��v���R�xP��N��T�$i_���}�ǯ��xV�tG�ͦ��T�'�T��իg���(��Je�R�S�5�ύ9�R8��ķ+�wq���=�.�(w�)k`�|Z[:���r����Jj�#���s���[�HV��p�ν���.��tC����kU;Y�7l����5��2����Y#`�M�v�����1S�rȻ��ׯ�Wd�P/�/8nܜ�|�N� �&�<#F�t ǖ�e %�� �[o&|��L���Vd����Qz�͛-R��%)���p�֖��P��;��̖��\�Wj3��t6��i�ef��� ��l�\%V�5�5\��#ѽ �Ya\f'�hȷ���k��	-����e[�ʅ��E^���Jp��1����ok���o�
Y�S��8����i�W)�+k}c_N���rl����}N�ox�����α��`����\��U�D�3T���&�mg+�3{1M٬&��JP'�3�km����8�hy�:_�q�z��Y�V1�U��\�F��h�s�D�%W����s���c����x�<�_N�kcS����\<z�u��)��O��꯾����������͝=��_@�~��RV�6�q��ފ��7�졂�
�6�V���9%�^븴�ڬM�5(������y˩�cR�4�3K�� �,no�Q'66��;Ē5���:����-���
�poob���"��
Jңd`��T8'P�Xt+Y�+:��+�3^�r�@�"�V/7k <3F0�f��vwv���D�ƖM����wW��κ�@��ƺѫŘ��j�x�P��tt
Ķ�\�`o.kee�c2�毛�	K̝����y���v뺔2�@�����WY���K���2�%uc����/>᙭�X2�������U>�u���&��4 ��P��[x_�6�u�v��f�ͩjJ뺖�"��`ǆ�î5�dP]�>qP��;.���T��y��SE>2�(��'>9k^vӷ��v� ��	|d�uڸa�X�%[��*X�,�vBYoK���	S �nsȓ����x��$���x�h��R�"U�m�y�t[�*��R+�f�>�����[�\{T�z3��Վ[U:�z����u3��WSg`�8�B$�;�W�4<����b��.��WK�g1}ɺ��zT����B�����l��&:n���V��}�˝\�A��;�q{2��0���=���NĦ%�L���^^��$+4U�KU�%U�V_7SM��}�)�s��_e���kjd���v���u�0�'�iN�����*�!Lne���n�+��!З����m��k;���ZE��G.
��u�w�,��'O ��B��ޕ��ʍdK��S���
��E�M���=V���ɖ�X�rwv�I�x���p��:G�j�����]�t�Eo"bIs8>˦��S�\9�nҮ����E1�yb��;�[!�1�M�4M��N���WJ���uٯS�Si�5�����;)ԥ��`IX��e�(Sp��1I����U��华>O�Cռ�W>��<
�뜅o�p�1��(e7B�(��N��(Y�y}u(V�ʠV��>۰�5ܥDC��`7�#� n�8*X����k�0�y��%Em�ζb���Q�l4�1��8�gnb�r�]Bdܢ�Z���KlҽpD�nAF���,����(
N]^U�wQ�FdZr}�(&&t��-�ދ�C�\1`�k�͒�@��f��Vs�o[���U�I`ԍ�v�����Q�!P�f�6�C^��]Y]�Eme��]��i��#��bM?4�ڡE��!�m����U�]�[�0KvF��?)����7���g���0���smvR*�`�yҷ'sU�pIm�E�WVg����+��f��>s(�
�
��8V)��D¨a���-�Vl9�rr$)�XɈ��BͲ��2j)
珕	̤{mX��}`=�h�$F5�@cEa�/3OWl�"DE��%�FV_D\�^e�U٫�� 8b����!'�Q'%HD3�z��o*
jm�h��}[�W&�t�aϙ�����w����3�6�9�Dø�p���D,֞�լ��gGI֣�:{)g��uv��=���4�'����X���k,�I'���k1����ȳV���@ӕeb�(�����7:d��̽u:��ZH�qᖹ�_}n���l>9�T���N�v{���:|��&�Ǵ�Y7�pͬɳpQڽ��4��|p�u�\��iX�J���)-���ca��_U	���v���9�x��KKz+wt�y;T*Q�s�RY��Z�vus(�5��ȶ�
B���o;iP֖�Z��l'y.�.�8�n���LcZU���]�;�%��J�n'���5:��}u���a*r��Q����sMmoPъ�>�[�-F.4[f���f�g_3˓�e���7�#u����l�r]u��pٚ�t��]�4���҃{{��;�Ov��ԧR�D���a�)kh�m�t��"_nR�윁Σ���7d52��[�˸�J�+�: �v�j�`�	9�S4��������R�{G���xC�:��1��cF��������D����MAK]�w5+���qPu��-̵،\�H>�n�ZJ#�������Z��Z�����,a,�B�d�|&�����n�s]<&�
x
t^��E�EԘ���̾�����Z<uV����-*�C�d'k_I-�f��1r"=Odi�(��&օC6�q�'�{W�vbo]4�����t���W��#��:��?HԘc\`*R>'�����iqVqmǀS_i��{��9��j��â�Id9���J=Δ����*�pDc�������e^p�>�V����1C}��F��4yP��R���j�����!dC$����T�p;h7/��-������{��wsx�����S�X�s_�����X�+���e��P.�D`z�O#��L{'h���(�e�;d�2V��u�7]R��BR�i%�V��;�.�i�Π-���V�2�V�Kr��z�m�U��[�_`O*f���I69��[D!
O,�.�T�'�P�K��vHY�6���R�-"1Q��ݎg���p!��]v�+�%�0AG��2r��^pJ�X��΃����g}�8��Knm
#���{D�����,]�8�L*Z���+�,|7���c��n���+5�݌Z܈�)Nʛ��o-��a�B�21���K䲷��²Ԭ�Ō�Ę0+�h�6K��qՊ;�SYtˡeG�����Y/�#JE[l�Ŋ��2����{�P�k��@r�q)9��tn����t�/6�k[�p�Am�Q�z�-ю�0��JWYCcd�.�Ad�ݬ]P��NV�=T�����ۧ��e(�B���8�]��6���t�:�9䃫�{���a��[�b��P�/R7�jZP�O�ì�xE&v��-��:�*�V�;T	=�����P�=��M�ȼ������H�`O���C�1�:�@�a���]ZWi,��k�FR�6����Y[�5e�oZ�4������@���|�bPk�JXs�t��������~�K�v�8u5�Q�2�����R�n}��BZ/m�L��x̝H
|������y��y�ΣS4w{4�g�����Mh���ə+V#k���-����)�}�ck��E��]�25����p���%
9An��G7�[2Za�u���؍t��Q,Pq?`G�E��t�������d�
^���{)S���#�o`�kB��n�\l�%�Q������B�КR=�7u�NڛƵ�ôt,k#\W�b�ǚZ����d�����<5o�2������x6�*D`й<��_L
�aU���/.�^	�n�|��o%Jv��zF�n�p���֩��}3�7#��4��-��ֺ�
;DS&ڭ�uve#?��=�&�LV�Q��� 0���ԗ�ѯ"�t`9��klnu�՝H.�&���nM��dݬt-��Y�C5mV����w���ړu�B�y\����x����9:�]ɍ�u��;���>]�oI�`#����>)�-6~��u&b�t+HPvv����k�͈�]�zjb��,Ejb��vbb'F9z,U�
�_#�����<O�w58�M�J:!<w-����J
�u���"k1䒲����T����|6��1u�s���t���x�I:�����e�^������G� nV�e���Wz(�b�v��27��&�VD��\. ����V��}�4+�l�Ha�_!X-�u�ǌ�j��'��s�uf�uv�)B;櫳sw�Ju>Kr������H`�)�s���h�(���#I�2�;�{�*Q��BfY��7 Hfqj��v�V`��DnP�%^��H�*�Qt,�c�vRQ輺
�!R�ub���@"���r��C�qYW�p�`:VIfJ T�)SS�s�Mw,��}˵*�Q5��Ԓ�۾|���Q7\�+ô 7X�Q���L[Zکiję'�{���/��CD�EeJ���R��BY�]�� �ؼ�!������X�C�_R�sq�=�͋�Zөݱ魏��\�P_n0v],��{vv���P/���ʑ�pWAo�V�a'�����vqw�I�ҩn�DpVo1�q��5���L=61 �0�@Y�	�gP����wl�/����\��M�����<��}�?����Wo"����Z^�{oUm����W=�]��{NP���sL�/D%��z�*���kq����VlK�����(qG:4�U���Z=L�vf�4!V.VG����t|R;8��l0p����(k2��6d��v䊝�uo9t6��4宱�E�}q��M��jݫ6љ���S��j5+�u<E�xe���6�Ɨ ���j����:��W�Li,����d@�-N�B䷠�[LuֻڻO���f0p5��ɖqF4���p�t.S�{��\��nR��*N)�:�%��/��@��������U�}��Uُ�rՍ��#͊d�\�̬7�#W��Էi��L� 5��p���h\�н���D��#o�Lzͧ�hǗ�b�;�*�����}�K�w�*�$���n��W8H�3���b�t��'D�R�0e��#LFԂ�,m��O�A�Y[dn�v:�6���U;��[ϫ�L��P˹	��{8A�F��̾.�SEKn��uܖ�<���(	υK��׸�#�8�R����慐::5�'g�3�ff2��51�ڤ8�.E��V�\�]\��3!��-H4^7]�l��(�y�2�`&BR�Uٜ�X��V �_n3�R�.�s9�������?Z�\�����^]���ހZ�z�I��r#x;ӡN�#�a^�/[�-j[��mbTW��� g;�QY �j�k��F0���kQS��v�����ŷ�6(/�S����y�칼�f�R�p�y���,�(��)dl3F��+o�,5/�rR��j�6�LDZ9$��R�R9x�H���.�	c��Ɩ��b�]
֍Mp��IO+��c�d�8�I���;�3d���2��I.D�����$%0#Pk0�I��o�g� �R/+>Ι�[��y$Ggc:�k�lG�Sn�pM7�(G��4�Kr�.����$��,H�|�F���gE�ۥI�0^����Z嬎�\dT�3p�2��E�D�h[�K(���f�v�@��j7"�YVAԎPr�A�F���ET[È������Wٙ3SĮ5V��M���D8wY�ڻڵ�!�d�ɡX�&��3
x(ťt�^*���x�m�;;��R8���g:&�Uδ��s������1"~ź���O�n�.m��Z��2��?�u	4r|c���I�swI��)`ӧu�Y��&��&�B�;R����t�~F���ݬ��6����� 6�
fl�Й�T��� ������v=�g�^Jw�|x���00���K�P�oMO_B��ɷg�g:Zk�Ej(]���G�(�:��@㵴���[V9��Ҳ�ug$v´; ��h5���sOV��ٵ;I�@|3B;{����f���Ԛ̦�m
B+/�ʓy��8r=F�q�ɣF�Ȅ�Α�]��0P(	�����]uh�b�0��Y+�U6�,K��z�ʽ͖�3(;��jL�9�db%�-��vh�8�?(�ˬγ�p *]�7r�U3(L!����c���-�����EjT���[���������J�]c%�nН�FVKB�U=����ɂ�4�"�@���M΅�
��7�-�:(Wo5�uej�G��Pʼ�W��kv1��c��e�gTzwU�w"�"�3U\���&Ӳ�;j���e�`|�>��]ʏ9�h���fR\l��ɜ�ۂ<[�of��6��z&���]�)w^6��"���n��ӯ0q��0��e:#�&�Jl��1ד�����Ƞt����/~����5btQ���d]�yS�:��6d$�**Kd�Q�*(P�;`��2��+c%CP:ݏn����A:1}ٛ��F7zڹ���)a�U����.W�@�	�us�R#В��ww�l�-�Z`��q���j���}`P�ΰ�V����ii���/�v���C�n
U���ř+�F�9����@ԝ�V��I��º�s� ���m6^ tkZ�i�����i6*��.��F���%J�sw����hgk�7�2���@�����j$6+p� }YPp�)*�dZ�um�:8sT7��B�'���4�ʽ���̹®|{vG��mD2�J�)V�� �t�P&��`��j���v�W"�t�6��x�[��;��t�v<�}����Tx]�!��r���H��������"��z�XQ�䮘�ʽ-ȳY��5-��U�*��cb�R��P�s�����K���j�9|,J

�tr�W+a�k�'R�����I�L���|DA*H�.��:T4\�ہ��� 3���q��ckeꘙ��R�8���.�Gps�]^�1T2X��R9���ӯ�%:f�����;���n:�K }i_W$FSYw�#cBW����w�)hzyq\*,�3m�w�hSa�[��5�pM}�KV�7Ê\�i����ʅ�A9l
8�h�3�՗�;]b�vJ�`rniX��~;O��;���՚� `�b݃z2��׮Z�,`s�j�-
�Mwrd�e�NM�;\�ʈ(�����5�F�-�Ww�ŋ��.3J��W$t\U+�ޡ�T�7�wj���b�m�C8�س{ͲW	���1(�G���cm̹��N׿]s5d \Zy��ӊ�-��Lr�va�o�?��H�3�9���a_gM���<VWeĲ�˫�u�����u�ľ��1���gZ[�[�ܣ�8ۉO�C�sjc0B�8X�z nR_;�S��0l������}��}��u�;��2ۚ.�ߗ<l�aR�1t!��Ã�o2�d8͌E�Χ���-ggiG8M�) �vV	���"��`,�<-�g�x���z��dER�mm���*�������UΔ/����_p3��������8�J#ku����.��<[�޽�4SXy��x>[�t��&w��B���z`�4̆@��un��:�sf�8�7��.�Y��$M��4=��,��N��7]i��I�K�o/����j�PE��c�*D�dw8`ռ: �����*ŝ�}��Y�Y�Z���G�ǯCI�1�,��1�7KVa�&��S=`��V�ںѫ�w`�
��˦3���91q�|�t��� Y�=�	ie�Z��:=9,.�)颱r)_aXTI[p�ÛZ��p2թY����mBf���oG�vw.���%QWX�S!\p��N�nr-U�k�)��7�/`ch�ʆ�	\���F�������m�d՛����&�
�S��E���l:жpn VE�\���ռ֭���Fg!����y��f+�y$}gF�h
��N�cz�D�`ױ��3v�˜�ъ��N��P�%u�e�H>I�+/@���9���+2ه�!0�*KK�pd���{�֢J��8m�ƫ�����Q|NZI��d�ttr4�)��TNeK����e��B�FCGw����r2�n1i�A�q�HE ns�clj39ˊn��9r�ɠ��e!.8$؈��,�BDIc7�L�`j$R��D��`q"��!������ ��".r拜�q�s��BL�s��$�$ȒXؓ`��\�	5$'�S&cF0�4�a$��.F�qE�\ع�F8�\9���i�DF2I	)�)�E��&a	$�I%�)3#d!L�..(̉1�M����
H�����Ɠ&�B`bd�&P#1
��W��~����|�{c�C���+�cD� �����ew[��u��]�%�@�]��>�c��T��o�Z����㚺nhr���f�=�W�}Xl��Y�C�\6�p���C`/�]С�Q�L�8|q������r����ۑ�0響c!�?Z�N�~�.��:?<�2.��9Ƭ'j
��<���JӮWW����/u�p�wy��eg²}�d�G�)�k´#��k�t��O_i:l6�M��v�*�{./w=q����a��u�#���,����N�!xP��Ph�2EX!�7{�4�c`�ި�w��z�O��:Y9}��T^����hs4�7*31���V�DE�>��0��b�==��41�W5�N�o�a1د��<�dC�L��u��ok��w���QBK-̪i���49���'�tC�,O�TX:�1��nuE�b)d�f�d�Tn����z�ηs��~ک� ì�~2��H�(!�1#o]b7�a�P\�����s���FU�����	�&b����ϖ�I�GA'j&P�B�Q�5�:w+�FXR����͙�%���&�_qȆ�����m|����2� �(	�<5d�a��b��Mj85our�/xq�F��.�����z��Y�
/g�}��ˬoy*$�S�NǼw��#�b��a���5��׫8��.��ܩ��Y}�W �(�9ͳ�e����t1cL6��sTe�ԡ�M�Z�P�ցg�<|�CWJ+7U�ʾ����yS�uM��n��-�9c��s����?e}��p.J5�@޹n���Nv���iN��E�NgB)k�1�W��9���븛��8j��k�q����s���y*i��_�D�Q13κ����~�P�����V�nQ0����$E�@�����s��Sosג�b<��<D�?y��B]�̡�m�۳����O��x��l�+2qm���^W]P)�L��F,�7��S���#�]_/�c��5�8��zf����]\����s7w�>hAܾ%�1ϊQtȲN��̓r�(Xr{ݗ�.���ᝊw��{M��Z)�c���˅����s�%�p'6��/�a����g+��� �MpQ9�{V���W[����f�(�y��2��o�}*}�(מ|��مn!����E!�����>�M�~�0ú�zhp�� ��u\.p�T��4dn���1�v���S��+�����U)������P��jE������?_.�.y�6K'�錊&�'`��n�����pX�°�H-ٛVM���<0�!2T]����3�1�����)Xa����ā����Jh\�W9omCX;�藹%>2�[SӶ:��i��X1�t9��X���Ws�w��e�mRgp�W/���g����(�������lw;{9$/�<N�ЙvP3�m|�&h���rxCA ��%>�<he��5w��i���b_�+�<#v��!�jN���$��O ;幞�]��{�j-��X��awH%ɇ	��3��� ��pܦT�_b1zx`���� �<��B%ԭvɞ��P�����݂�'�VH��L'�����pt�d9���Bj��Sl��,B��=�|��{m�� '�+���,�=��wQ-R�:K/�{M�}'�8$]WF_a������y�ɨ�$�C�� ��k	�w��e}����PبS���>J�.+�֑��w9C��ф�"�TP�S%MG1?|"4�A�ǒ�]�.�~����i��ߏ7�nM�Sy{6�G.!\�.w�\:��rD�kG�@J㢝R=���A����-�֍�X�T��������М�b˛d�&��6�
��31��V�-���8UZX9e\H�Ň�7OY�7Z1�{J���Q��u2��2^'�'�Y��O�+��ܺ[B���DCl��J�G���}�Xѭ"h3�L��(H�4�4��|%]��߈�$&N�=N�̮�A'�Z���L���*3�&WZ�;4���tY��m.L戫[�r=0��j��ZƖ��JU��V9��R�P�+�Ź�����r�z�e�)�X�R����Q�w���ȴX']��u[�U��9۳Jo��Y�ďr)$�L��J'k��T���P�ٽlh�4XJe��R��$LI�k�[�Cr{]�b��ʘ��c�̠`�F����h�L��}����V��ұ�Rf`&-f<���\U������=콎DW��6B��?Mà�,4
��,�Hj2d�YX��̍�V>n��g�d�C�M_�|�8�4cs��.et�u��ZKj�@)�Xy�^�z{�q��=�%�:�1#vq�å��S�3)�c"���wMr�P�4�	�jJ���B�(�$���Pedi�`�X��pܦz\�|���9�%���y���Y6{4��t�0d��u8��wMH��Jܮ;�&�r�WD��\H���b����}�{�lm�Iet������l퍺�<hBy? k������U���u�Y�j�I��F�ޣC��� �UB���I@B1�q��VYT�3���<��Ԉ�wo6�:��X;�.�x�"T!:)V�Z���*�-�	n��(F����]$'ݣ�ƽ$�z��;]�o�ouS��1�N[}�C�͕��b2�q��E,m
�E�S��gE�]e�4�N��Et��Қkt�B�yvZQL��Ɇ;CrDuC�r2�wV�"A�GAx�%?�*4�R*4ޅ��M�H�|�L��l��z�v|��f3�se��\���u����(�*�#�6�зQ�cst��$�t�]��t�8e�����З[c�����J�k�R�':�e���G�`K
�[�3�ہ3o�/TI����&�i�Q(g���K%�(O*���v-�-Vy�/;�P2#��@Hg�� �m��r�fDt\�*�8�޺�|�I{��^�F�<y�$7�g=�1����@��uA��F��˖a�^��ƹ�G��x�s
�\��ƚ�Ӑ���d�#ʠ���g.1$ܱ��Y�ma�Z��đO4P��}]���M�gY�M}�#��_�^uBv�"��C$Z �a�*{�,e�H(b�zi�Y()7'�'O��L
����k=�j�fwi��8Qen1G�vw
���Q\��;� x��><**��A�@1�ʴu�uM��S��K�wVX%�B+w.��. ��Hs� +*�����Ad�n������ݡ����nIܝ�e�XԷ��q��j�!C��\a���ئ�<�\�!��	+5A����CT��9���wf�J+���r�>�� ��(��y���g����A��R�5;W^G0�vbs��7�{��<q�D*����TX:�1�*�7<U@D�Ƹ����R˔#zgGj��}���,$�uH�+���k�pWP<r��R�/�l�a����-���-��<�{p���Z�;>U��`6L!���T� �{]t��\~�n��������.����-�&�+|q�,�9��m<�-��/"�QP �A(�]��7|��5���W�����l�;u��Al��r�i�#OY�~�uP�+�%%V\ۑC#�9�f��Q o82�Ā����]p���e1�j�� �?�%'N��,gL�U�C��s��#�?8F(��:LO�ʵDdu�Hm���c�rd���A�C$B�y��&�^8�q��|��n�
5����D%���g�㛳�Y�X�
��M�ؽ6�l��V/�뺱D�� VL��2R����� ��A��Ax�/�"Q��C��X�	���nt����ڨ"�d�M���>e(�dY&F�ge��㗭�Ú2-�"Xk6��-�-݈�D�їYq�p,�k|���AB�wo�"�W�����b��������+~�X�d��<훺�au̱ΐvΣ�u��[l^���G��kb�p�.�n֥ڊřw���|1�:;����ݣ����^��j#���������[��ȍs�&�K�;7{f�O��3M�z:�r��O�m-[��=S�Lp�0�ஷZLf�١a����jt8���͵x,�����<�ri�8G�� ��vXHW`�0�pV���]C��yS�1�:��;�g��bM_w�͌=>�c�ոВ�q9�⫬��j��K�N��W �{a|$��lX������[����j�G<�����<NŒ��q��&u9�Ң�ˉ�\o*vVl.U�@LM}	O2��|�(s�7o���tܝ���pN�r !X��=�۴Y[�-��S�v�I�[?u@�H��Xm�L�����Z�}�]���qb���S ��md�w(�����G���Z�&��c�|!�`3���}�X��4d���v���i�bq��*��&|H�.aq����j�p�j����1����ͽu�3�B'"����JE�K�n��rYQ�͟��"�&�;�ݲ��U����=�-�g��[%�n	�Œ�W�.�x=yT���*�Q���ÈPCI֫C;[F���CJ+�m�����,M���@zz�ߨv�Kb�^]=LE�ƣ�r�Ue�1w�v��r���m�g�����l�]��0�[[(t��c\�1�m��9�*,�x3�ՊA����}�F��*"�3�>H�z@�md^�`=9:�40õa��9�;"�Z��?�u��s�9�yXn��U�%JRWH���3-�3J���ܛ��;�E���V���mD%��c�0�s6�hN �"B�EG��[��!^lf���l�Y�Dpܗ����c���T�����>�5�1q�l�2K6㫊�.c')c�w��~}��}5���\�e�U�ջ'�&�w"�`9���$�<غ������<��F�ӎ��V��?^6>��b@�(C��cE�,ZULD�6j9͑��suZMGu�4��Q\:B�94��Q�N�l;�Q�uҝ�q�4��X�����hnE���<o1Y8�J{[�C�L��o�T�4q����{s���"���CУ�X�N���(�G2Lį��9劲��8�8X����*k�d行���O�V�ޙT)�Vo��q.�]�㣛NK1z��f
�ٷ&*��������\����`fP}Xȡ��0��ڽ�+z����c,ԙ��W�O$+�1�fx���\��
�)��Vŗ��������WN��s*ۜu��[B�7�Tr��=Q[����9&���ʹ��
��q�0
��}HT�_a�XÕt�}ns�&��X��������n�;�d��5b�3b��,I<#"6�V�!�5��T-��nS=��Ad��BQ�11�V��W!�񎻙������UEk�)��g���]:t���g�0\>b��:5H���c�3�/a[�@^��vN���rYA�$�g�@��F[;m�K�P}����/�P���V���[V\BrQ���B�q���n��p�@��~��|+t�B�{�E=�[b�LeN'�]5���p�;����
f�8ܑ_<w#-�Z5jdiꉐ}[=gx(z⎂��-M���
��/�0���Ἡ�f2 �h�s�u�U�E|�K6�e)�=�&��kuD��.H��8�h_Ԧ��,$x}��[2�\@#)��'���7�N���i�M)�Q�z�b��^eN7����rj���(>�r��z�ܔ�^Wx�
�[��Z<�;]S�y��ޭF�[@N�N(3����0�#��
��"���TjM����.C�}:�K����Cr����e��Lt�z������R�p�m����0��}9J��zWt��ַ�ԋ�&VM�+����ۆ�f�4�J�w�
�a�y���R��Uˮ���b���Z�*�<V0l�������uќ��e����*��b����Z���b�օ��@�8��C���
����4���ltr��qj�M,��]�)ˍ9��U�k���,F�7�b����0�p������5A���[1;|2T7���r�'M���4/k����"��,���'��(2*H�ת���#}�%�(�2��6��V�8dY����D���不��������3������!j�3J(h8'�jo'�OX»O���(�`xK5�)��q<�φ:��xUf�2��V�
���w�O|����L�����tB���� �|:�1�&+�/mڹ�y��ζ�f���n��n�������R6�t���g���|sL(��[�3�f5�_7e^�ֻ�r5������G]����������4H��A'�. v�v�m�$����wx�^m7����u0x�&�%o�5%�� h�6��\!p�m���(�B�	��)ě7"&�3Yu�А"M��֧��L�;u��l��|��Gc��=g��$����쏺ڡr���Rh��m|d�I����(E|��Z��9��NwI}S�|V\R��>JԺ��=��{����v�����Mp�6��5��a�$�m�\E����+ul�ZeۅA²�_%V��v�hͬ�D�0�h�X$̓�ۜ��Z���W�Ǫ�I؛�7�2�r��Ƴғ�S���Xط�*q�d9��.�!N�+w�5�o��L}|2r�&���7o�>��V��h�U��p1��U2t}�V��Gu̇*;�ܣǖ{��lQ��V��5`�Y�� Gm�OZ4�*<��3%�qS�6Nr7�}�X��o!j���\7��n�e���4Z<��!h��}w�ͅʰ;U ���-?��1o-�EM��w�^��mQ�,t�
���n�vu%�V\خY����nAȌ�Q�p�̹I�ԭ�n��_6i��U�8A�;EoL�Μ���(j\����7DJ�^Ɇ�c��
y�Z=x��{J�;E�Im�+�Ӥ��ևj��j�Z��y�&zj1�h�`6W��U_mG��ys�w|���"��ʵXʰu�շ�#�"�D�sz��_LJ�gd�m�($u���q�1˱���G�:5+�i-�7�5��T^Vl8��4�v,Mw=6Fm��։��tő�i�5غJ ȈUt�:�K���a�e��ʕ��;�� շ�ʔ��@,\F]��`��phB��m��X�Y�b�	qp\t���F����Q�9����涘X!�o:�mu�#s�nu�"�ۮm�vT�����1Gp1j�� VyL������qt�v+Բ��]�1O�XX4�v�o����
n�N,����yK��8�!��<��ޤ;v9�u"%M2L����M���ɹ��T�ƅӖ�iZ�Z�'8(𻝅��_o.���յ��aoܶ�V&����M�gx����VX�:�;�)�Is��yW�v�vD	ɛ�5.E�4��4����s�R���w��ӭ��114ܧ@1-2�԰�ٗݚk9lҌ��4�+V�u�ǭ\�F�����b��g8Q�֝�`+��8
A�(��dU;N'���ȭ"����A�-��gu�R�� �}���a��� ��W�"!j]7�q�v�e������V�	��u���G�����+��ON�J�����Dse��j`�o[�+z��r����Kuc�5�U�R�`�L9Pd�B�PA�͙g8;�4��$]�4^�]�&�Z9�`���dG��f�ݷW�n�Ov��ز���H�NH#�B�nV�uEGJa�fk֏.��P��Hz�r�+{n+���A9��Vk���V���W;7]:���.G[s~�Tf-���I�}�Ju�ao�7�m�Q�u����H����(v�:wQ���F�����h�t[�{n�x�7�����1���3��噍w+7j�8l�jq긫9����y�(�
�Qq��52��bm�{t���ih���XN8Qv��s���9���*��q���d�ԪH���pFh�%�s���e?��3	�"1)"L����DƄ�܁�#
�.DR&h�Q)LٌI1�H��R`��I"L�e	&I@	H���H	��c$�a!�&Js�"a$C$�M3���3��8���J(㒉(�4�"��2RP�b�Y&A�IDq�.Y"8�%���s�2�8�bB	D&D(��0�d�$2P
 Is�Ll�p�
C$..@�"�1��I$�dI�rA����e	db�3`q�cd�$�e8�)F!�3s�Id�����%2������H�(�7 �$+��s�:�v�8S�{-<pne�@���ڌ1ݸ�v�[�s��Y;�����k#�LCx���c��ogr���`�����]��z~WkAz��Eq}WKw_y]s����^�˷�n�KG}���6�������r���<�{�y�zZ~���������U���~��{~{o͸��M-����r=�q0�т!�}"$o7�u�{W�t��~��^���9���Wǋ�ѻ^�\Ӯ[�LU��]E�~�t��/����\n������[��o~�]7�����7���^փx�|��9O'H�u.s~�*���|#H���ݏ˦�6��μ^��nu���7<���+������ʋzW�~�zz��\n���^����F��6�ߗ�����CQ�?/�ڽ��\��;���ν6IB�[9o����}0�c��]����7���|W����>�]�Ҹ����]��WK���=߼�o���׏��uoKzW��y�>sn�Kt�]-?s��Wk��v������~/ݹ�X����3:S�E�����`����7CS���������z���6�~[㦾߾��|^֍�����w{k��Z>o�;�b+�Һo[ϝmߜ��n��ߞ�.6>��L|����~�Qd02{{��ӹJ
br�������c�<��]�>r��t7��U����x���ۋ�}��~W��n�B��?��k~W6�w뻞�k��n~��{x�^֍���﬘�	g�鈠� G��-�p���מ������7�c�|x��G�f0_��[��^ＷM�t�K�_���Z�]�>5�]-?r�^�v���mҽs����6�\����[�ߕ��|k��UG�D� %�ޅ�|}0.��&xSM*����]#��}�h���4o/<��6��W������5�j7��ޗ��]��|��t�+��_����֍�_���^7�zZ�v��qo]w�w���].�V���*���A�Ǥ���^λ����J�Gz�<����+���ޭ��Ϳ.�����O������:ߛv��r_k�k��7��k��}W�۶�m���7N���{�˾j�-��z���/KF����^/Mz~Q#��݁�r�P���;˵�"�����^u�����o�z�_��6�t���n��ۯ9o��y�kAx۟�{�긴������:�c~m��WK�n�7�nz�+�M�]��m��UǊ��W���؝-�c�3�07��ܛ7hgK��+JB��X�����߻���ŝ8NA+|&���c�z%�@����A���w;���B��y�Np��+�"�����c���J�Z ���k���M�'L�v����j���J �I���}���������}�o�kG�\�6n������h����۝sW�_��q~k��o���sWM�x�K��羯�h����������u��Ŏ���&������Q�`�{1vz>����}�I�#ط[�ߕ_U�\�m��kz�z�ޯ�vp>t@�<��� C�~@�����G�C}�99�>��"8G���V�r}���5��\}p��D���wr�r�+���]sv��Ƹ�w:���ۥ�W��/�����_}sһZw�~����}m�^�=߽u��7G��B���"�~���G������E�K�C��o/�G�>�">B=��}�[㧭���x���^�Mt�]-���*"����v��͍���??-��ۥҽ��t�|��~�>o�u�- |��}돐��@���gGg��Cϫ(�W���� ���#��ީ�DX�>�æ�k��ίK~W[t��^wk��W ��	�>>Q�q#��@�q�9�~t���Wu�/߹^���:#�$	����`z��4ɟC7�|8x�y�2��~�����`xw����|
��:�o�~WM�]y����ŏ���^w�_��۝r���u�ok}W��箵��-qn׭��k��:��\z���6�#���I�@��G��1���A�>�Ll˭/c�x\	�������0>�`ks�<��]��~n�����닥�+���{����]5{��]��\[�q{�;����+�����]kү�Ƹ�7K��n��\��u^���o��yþ=���箖;Teng{s�`|!�<	� T}���W���]Ϳ7����}��ۦ�����[�:[���׮�k������Mzn�KG����5���OJ�^�yջTA�<1��b>��;�i%3���%����}"$G�b"G�O�J?E���h����n�彫����;���7��ow|�����M�{����ߕ���>� ��O�T
D|}�/�$���@P>����m�+L��j������-ۥ�}��kE�����|�M�nu����]5��k��|]���׽���������w�Ż|k�k�}�ֻ���ǋ�_7�ޯj�\o���|��������3x~��t�R(nݜ�X�:�Q��������bȭj�7�d��J� "��.��u��J��nQ���u�m�gEe���q��l9\z��4#�i�)��i�o����4���N�*����7�m)ě�K��([Ui󷣳z�rns�a���uck=��d��D�=�@T}� ��6��n������zm�z�����Mv��|�t����_9ߕ�t��+��hߝ���o���5� }X*���Ue����/`�����i�s���+#�&�ֺ>���|1JZ���Kt�����^-��m�u�y��{W��|�^�9���6�ޯܽ���7�^��]���6����WK~on�RG��|}������w}`�b�o�<���~]5yu����Mt������Uv6"������^֞so���zo���n�_�]Z�|�u�����U�^ւ���|�^�r�UҢw��n����b#�(D���#�u~���
���f������~��o�zW�]�E�n�~|�,5��*��П��8SX�W�}���-����Z
���뵿�r�o͹�/���W���5���7���W�����~�"��@��'x z�Հ��vs����{okq�_�鍟�\X��/.���x����s�]�6�o���n�����7�v��󯼷�r�n�qx�ו��;�ѣq����/m~k�?��(t@���C���^��/|,���3;��||���%L@ 8E��^۶�+��5��+�|u�Z~�W]����oJ�.7��.��}}m�^�z�ҺW�p�ͽ߽�����pG��=������#�+�(TI�}�a�c[[�D}�G�>q��� T��9����ν�E�o�Ow�׵z��\o�^�5�~]6����}k��]?7-�^���_U���5��tߟ��>�e�X�����EP�t�R�mhM쪯p�y�mx}������O���d}�]-���U�\�m���{�?��*�q~m�������oKv�?���W��j-��t�ۥ��j��s��ns�>�׫�U�~m�r��-��>s�;���"�il��������}���-����~wo��ѽ.u�Z�}W�t�������n>����y�v��ŏ������Wk���{�{��ۥ�/w�|��?�&��ؖ@�Wb�/���48��1��ϽX���",E��^=�4h�[��:[��t�ָC$>�����2>>p�/�+�x�Z|�u�+��o�_7^uWc_ƽ_���zZu�|^��}^׷�����z��BP-.VݭkE;%�p\v��6�\�,0b�K�S��3V��-�B����R��p���TWm����ޑe�d���ۣ�ık���k�7�"u��4Nt����me��h�q|�g/�wc^�E�;� {���E�#7�e����&u%nv�w��W
C�!���SHW�>s^�����+���_y�o���ۏ~�������|{��V�o��������5�o_�}���+��k���}x�綺o#��}����D�=����1tNyg�u��ϟ}�������U�+�Ӿo_y]7m���?�n�KF��5��]��+���w�W�ny�v��׮m��_[t7m���U�W���o����tۋx�=��� ��
���x�����mGL̍�uތ,}�~�����>����?>^��F�ۜ����������]-��WM��\��Z�~_��]^-�zZ7��u}k��W�k��7�q�ٳ#�� [byL��]i={¼�=[�7��� �c�}����g�}0>|��۞s����]�⸸��ל��u֮��n/��x��F⾷Kx�]5���Qo���~�Ż��\o�J��2W��v-v��	���������;��+*c�	z�N.t�p2���ؾ/fr���M�6��N�1�N�U*�ʔ���n����'ODoJf�6�����E}���/9�	���L��DT�Lؓu�T�}����C�\���t����u��B������N��S�w&3��w�� %���^����9թ�L������iq*�f�M@b���\؞i��vpZ��Ո3�X:�A��l!�����5��Yq�@~#ĥf~�0vaT'�Ґ��|�`Pt�^Ty�l
�u�$r=�uۦ!_Ϋ���;�?�cC%E��/�wŕ��H״Σу����m�ҷ�`�Iv�c0n%Zԏ3--���1��X܊ԫ�J��(d7���e�)��F+�f�g.�*��]CF�]���$a�ջ�o���U�K��3a�Z�8m\�G������� g��I�&��\��,�|\��� �m̜t��}bwnѠt����DT�ƈa�{p������S�ú���〓�.���[�k�(A�uV�RK?wؤV���m�i�RY|ph�6���[��^@6
7��u���j�c嵵�����0z���@)��㮩2���:,8��;�F��o��h[���)۴'�ntכ�V�`D��`1ј��<&'{f�2�R�\89j�b�w�5���hշ�����vOn��=?XdC3����$�h�~F��]]���Ri�����]���-�'�(2[s�8y�%x�~l��`��Fa�6����K��t�h��j�����F��T2Ss���L��F,	�UH�3�5�_Zsy�=�.��}'�Ͻ�k����7�t�6���5$t,�ɢې5�f�m��d��d3�p�$r�J�n�*kbz� p���AOY�Zy]
�C��R_%�8�?2^s~n��Q:zB�)���nӑ��u���l�dDh�;l�p�#���U����L�jT�#>��q���ZR��y*���U�WyX�Z�>aw��*de�!{�{�$�4�3�w�ΣcD�>�g��^�r�dw-�.f�9ͦ,�9��#f��� yǮn��؏'ǎ�Pwѧx������m=E@v�A��J-�H�Ӝr��X��Uq����s���C��;�e���upl�
�@����+	
�[��6���XW�hW�������M��{8�y�`��s��jhw�^��WR.�Y;�Uu�G��j+ ��;�6��\3rٛQ�Uƀ|����'����\ ���eLx+~�Z9����2��=��`=Q=C'��,�Eù�\F�p,2R<����a3�369�!�jN���O��]���^�T����&x+���/�BLTB���*@�A@"��S<���Q��a��G���4!��ڎ���U��z��(xW��$~|���T¥����Hf|�:�\l��2��F�3��@���6��XA$�|e0q!���6GK��hcy���J��2�l�{I��u��WiQɣ|��e��|2K1��� %:NA<��'���qul]����ϱ70�3��h.r��)��n��^�#4�(M|�J����~iV�#�uin�@����]2s��\k䜤T:!��9��nw�_��I�$O��Q���{���Qkp�Lo�DX|�:�la�սt0�9O��QP����6/��"�7I�ŃK�Coq-���^��T��9e���{1�L�*d���(�KKUc���i�Q	]��E����V��AX�Q���Z��iXŴ���뤬�Ո���З�<��Z�z��6pQ�	u�&loQ	u�6��-��%�#ZB�D�rwr��r
�oZ�:fae�`��0��v�+���q�1�:4z!9��x5���XgF8�z����g��)�'P���CDW���笫5����ozD�9��hȽOi����oH.�#�j����x�b�IA���b@�P�]z*p�ݙ^�މear\��-вzsØlr��k��\9�v[1#c��D`D�|��ݘ]YM�ɡht�'���1�sU���p�xB�_*b9�WQ;o/EB��.�X8B� ���Y��@�
S���4�����ĝd���#o��X�+x�"b������Cy^��p�t�B��W{wo�e���x[�%�4�͉�|ǵ.!�����\���]��`fFByw՞[P���
�H�+��6��Rm�0V�^��z�
c�t3��;�"����L��u�-���K�o,�;԰n��i��m��}���(�|#Kt���Ӥ�D'*A-۸:xk�{ʋ������wdF��JW�X�VR�`E"���:�m+�Xb�׮�~i)e���Rv�9N�p�����17�;�B��t��&Ev� ���	����������.;c�E�7�����;�����3���{��\2c*�%�V�Ԙԋ�^�N��ω�ٺ�6&��@=��礪��d�P�J�?A���gb2�Vk0H\�r�1�q��X����T��RY����M�ꑶ�Ͻ>�Y=���u[�V�r=�' ��E��8@�un����u΂�<wM9��i�nH�x�E���ѫ�2�v�]^����,�fާ�CO?�d��_�HzS�[a���,7���="�>�5������;#{���=ƃ�L�i4Ek�H�jbS�^4���G���0�9j�*��n��֣�U��G<�d�����J�.NF�;Dhr:JE���N9�F:6�j�o�Sw8��X���+,��t�Y�\�D'QQ8�����v��t�xZP\��y��N^vWʷbD4�-mUɱ���7,/!��^�Od|�H�AJ�i]��5SW[��ٲ�β���1��n�_�;�8�����,F��C�ɛ�dV	Γ5W5ų9��M�,�|&������7�/�������E���/>�&�/i1���:������
	䧔�U��7Y31�Ak.��6jn�$e_��i8�'�R͚�d� �80�����Wě���~��Xm�O�UD���jN}�y�W��+�f��^ec]]Q핔 ���Ð묒�+V�oﾏ����Nt&�TX4ti1�pR2p99& �d�}���ֲ�/��ҫ�|m�z(�c�y���eè�-N��p��{���5>�ma�@I\½��q;0�`xJ�5�*��A��"���O�4����+Ż�n��Y���m�p���qe��?Pa��mP	e�S�J;UG<�@,����dp��{�C�[�-Ϫy�WJ�z<6����lhd������-}�y^qH<l:h>�۹ֲ
(G@<Z�w:zph�=�L����[||���N�r���]NE����m��ۈ�"���x��H<j8�4������D!������}�3��O�xg���˩��n���	%!��?uL�[�_MAl��q�-v��r4��u�*f�+�:+2��Jp��_U1�Ǡ��d ��EDϧ3��]p���e�����L#��5urn+�-�i�P�4!.��"�(v�PXM/���1���iu��n+a�<��-,�C�ڴ0�H���ņM6�@�x�$@f.8��������h��r�u,e�8�U�iՙEg����L�׃^��n焮���J�WY�H����C��,�y�O���$á����w��b9,��O2/�hV�jS�B�����ᴺ�.J��8�����[[z�Y������F��.��X��x�=�bF1q@����2�� >��辇u���:Riy�}б��V�8���-L���b��T��Jg����2��7�0m.O.j�K����z����Z;F��qI�|�Id�Mm��H^j�$�Èq-�
�
��7^�]��0W��uMm���d�wGa�q�lrw|c#\�ɨy.���L��k{hF;�}l4=Ps����]�+��:Lnl��6hXa){p�Q:70g���L�k��c琱z���ɮ�
�@���C>�XHW�ܯ1�8+�Q�������$ޏ:cܵ�W+y{<��ɍ�u���V��>*���/�Eb���n-T
�0�m_`�-�%11�	��ȹ�P�9~��o����b��䐂<N�ЙvSֈ��Y�Y�O���*D�
5=�w�h����p�,2j�e����a_�xF�:�z�8-]E�M6�?RvO�������$��R3q�N�]1$?�Oڄ[L(V�nS+��{]A0����B�a%�d.!Q�$�,B3���n�ҕf$J�L|�Hc��T$�J�����rkV�B�@����q�\����0�ɲ��b��n��*���_�拥�enb�϶ԏ$y]��i�t��k���5�7u��SfXXT.���^t
�gN삚y�ւ���x�>��s\e��,W9N#S{M�6a�ON�:`�"�ͧ8r7�nl�JdX;�cѧ�_*0`��5��Q����B�QR���t���2�Ɔ���БD*JwMɕ��#}�])�v�x1\3�u�����ìVt{XqH�6�!YV*�l�8��#�*��ò�6�ŗs2�a�����������.��^����5��%j9{���
3�5��ڀ#ײ}�Q�����m���b�e��U�{����'G+'�Yͭr��ܢ�ӵ�؅���_�1��a�5�1��T��S��]kM@��7��ۧ��5��Y�.����2W=��s����)����l8h�T�`������ޣ�����ׄ��Kcl�����7�]k��W6���;j���n�b�c�r�@Һ��#O��Ara�R�V;�1���wn��R�tv�U�t1lR���wNo�u-�2�<�v�jDb�ݬi\��:Î�e�S�x2���:�s�s���G\�{;6��$um���Dw6˦�<����WVu��#Oq�v�9y��B�빀����Y��n�����J$�8d���wt�i]/�EW;��������A�9�+������ݫ�7p�nU�'h�S�J����׹X_�0��-yn�B���=��[����`�G���/Ov@\� 4ۀJ]8���#�eu�A.ͫSoN��5}��W!ä�J�Đ����GmS2�v�c�3����sܑU��x��ܘ��-���p!u�6�Ҷu�KJ�%.3<�����?bx���{��۽b0*YTh<0n�;X�ax�h�6��ivfV��٣-����ՠ���p�+�l�|7���k����jL�*T�xz�Co�@�7J��`�U��Z����U��J=Pw�����fT�f��Y�s*�[�	��EM�|鈵�If�ˍ�i���=��K�G��ز�Yw���$�tv�O���׸2K���������v?Z����~r>��@�*mh��@m)��R�3�5�����^n�6���^���i@uPnW�w5�S�Fsd�'m4�0{���Gs�G�L8�9S�ˑj�	�,�
�7�y}�nOIG��V����1�����L��8�/� �t���L���oM13r���C���]�´k�&Ħ1�]�xSZ�֧�Mܮ���l�*=�O�'v��[�n�iF����*eګ#��l�#{�R�x�b��K�ެv�esˇ��*�3�.��":��]>���P=34C����2��S�nձ-f p⽌W$\����xd9��C���\^���.|@����Uo�q�%�G�wcA����u�Ff�,�XE	�J��� #&�%,d1SE$�T@�a;m�$�9�a6�#�A1�!E$#�*E$��,���!�	HH�IA�8ۈJ0b�#)q�"1Mj4�㒃D�AL�8��DF��c�Bl��T3�`I�PPb�P��Cb�s��2AD!��#04�FjJ�(�У �lh&d�Q��ƍ��A�%0�
1&�N+� �%��4A1A	3%$�Q!&ɀ�&��"3WQ2�$DSLc%�9�e[��"TD�F�!���6 �A�#���h@�B���B�
��^�qt��Aء�|�>��-����ǉ[��]3Żq��0�ޗ�r�����\̽�
�)`EO�(��}7�������V��r�+yp(��I�>�*���X�&�O��{��.7�]�K����B5��l�0\�B��e�{\�gϤ��������<%��xP4�ZM�<��Y.X�}�s�IS{R�-ϴ6�\U�w/�9O����M��#j�BQ%NDq #K�b{�ud2˙�9���p�ْD>8���9�,���s���n�������_=�cL]�j�󼋓s�d�K& !���ؼ��)���j]NKf4B�D��uF@���ӽK'w����vg$1+�8A1���J�bE;W��+M�:!�|jLW$��(>Cb��5��/\v��-�(XA˳$�,�Qs�  ���Bℹ�*�C�Cv��qͳw1�v�aSs��8e �i9`I�s��A��N��6>�����a<U֯G^���\�9IV-5gE�T�-r�bB���P��c��@��0�:�ý�SG3wX��r�����'a�۔\EL�����H�ٶ���C�k�1��������;�b�Ϡ��LA~�ސN�ZE�iE���wp��E�n	Zc�y�H֢�Uv�<0����nح��FC�s��ۙ�(�^(:����LJhLxmq�&=�O��[Ci�\�ὃp�2�ECz{�7�U)[���Ζ�[F�Y�Vq�vZq�pWl��决�Zw�������b��M��"B���[ZD��G��D�����Ҧ��N��_˝}���=��^5<�$f�r��(��	IÄ�x&~d�83�J��ώ�F�R�������x�j�u�)�nd��p����`��GuB��(]L�J�+#L�k k���2�:a�};B�aV�!�<�d;����nef��_��QZ�Jin�H�W���׫h�sU8�{.wR쭡�J�d>e�c��'=%T�Qd��$�3����]֢�r�mj��~�.�?jX��$'O��~��U�-�b{D-7z�m�wz��\���+���/y�{�S��# 0�"D6v�5U���qW�{�&�=���ˇuhֈT/��H�d���l���;W��q����@S<"���-���
��~��ň쉩\��.3:.��ƃ��	<6�L���DV���H�1*�÷����u���a�����:fHZ�λ�(�~'g�_Ծ�|�=+�������:G�3�i?�_��[\���3��q�����o��n;�d'�������pm�u�K�C�6��E$U|��ή"W\�RĆ�z[�����������l���t_�4�������=��ҏP�b��ӗ՝Ia���fw2���A��{�,��>�����#�r����;uV����?W%L��E�������a٠z�_K�pd�ݨmgV�[;��y�1s���e�����2�r����e��H��u}���.���L�a�� �Y�\U�v�]0�+^�H&�090�Z��.�rM�h�oi�q��8���Y��Ppjxe���M���\O�����_�zG��}���ު]΢�����vBS�f����7���~8����<9�(����3�{Ʃ��;��z%]Oԇ��2����77y����4���
�{O
��a��P�:-�ݚ��zKU�����φ|�+"�}�[��ѽ�<n,�R�N�U���5����He����M���
�!��䊅���S�#�y�u��Ϋ�42TXI���Q?�5T��;T�v������e@��Ɛ}9�ӟ�ˇ�	������U��@d�Ԣ+��=z秳7�0g�(�����Y�}�AҀӰ�y��w��9!]KZy����T�`�ř���.7�u��45u�L�*��*yQ.5�Z�.ܾڱar`!�w[C�������݋��^.�/\�/1Qq���:]�W�ja���[:��'N��\X#�A�g+S��γ@w=:�ۢb��*n��T��Es���$2��ۆO�?��������,�j~�b$?갬A� `Wç��ZS�T�eӟ�����E�W�t����Cn:�+O����t;@�( k���T�P���ŭ��]vFД�����s����=w��U9�����W�X�Y=�A����w�g7g�4��p�ڤ�EN��@v�'~0Y���F��-�ؠ�����{+c�SH�GY�Cv�p���V�8��;�����@7���NK���K��x�i�߳ݚ��kἬ;k��2�Wq�����j�����4m�@s�f�nnUh�N5F��u�����}N�ݔ��nz�P��v��Zy]
�CںS��\�ɹ��ϻ�ø��Εի Or��ᗦp��;E�.�1�xlu)�c�e{4,0����ޣ�}�JA��׫��+�|�<U�5
�@��}ʬ$+�չ^b���W<�&_/T{]�&��Uu�	����o�>sԱ�s־�q�&��
��Ϲ�y���t��aecR:.�b�c;I���4��X^�+\��16���=M�j�/��k�z�0��1�g=v"���v�Z��	�����[5� �L �f��HOk,�k�i��K�%��b`�hL�S�Zgs�b�]�[M~���ﾉ�0�H�A5f��d�	� L_.�.y�6NAb1t�j�E�=��$��d���c�/��ȕի�YfUC�uH�u�CF�ˀ�a�P��/���s:#1�;�6e�Xf.���:���������&����ѥ�U6s��_k�pP�6ܦVU�h��Y��)�ˇ�[��e^��L_ ��[$�(C�vv0eR��ù
%}o��庾z�+5��'sl6�AV�0��Cނ���W�	:���H5�sdt���n9��]ї��e��т��F2IöX�p�Н���$�o
�R�%��ޛܹ�df�3|^�Il���|�C��p��p�S���s�I_=�#j���O+� �����97Sp�w���%pDk;[��@[Ҿ@7ɳlCeC���w�\��6��/�V#��Z�j|���/f�� ������̍2����j]NKf4B�2X�.{��1�gJ�3B�.W���M�"��
d>5%��QѶB���w����T���&c�E	����Ʊ��Εm����s�ٴ}��`���
�a=��&8��\x�{[2b��J���S=9�5��d�����(�n�t�&����,�9x:��҅rR�P%�x�`�k�!f6 �x(�v�<���/�`Em�ʹAg_Cbu]�R��}����I�N/!��u:Q��|�K�$�D�����ي��
.�nL!��`��Q3�X�ȌkZ7\kԦ83�y'�yx]o�R��Ѡ]Z�8Ūݔ1���D[�}p�؉����{���$�j��xj�	L�]j��;-���k�
vx�t�:^�2umA����I�pV�M)�p.(nK�x��D��u�tܬ^���K?x�9��~H���\�V6;Y���v�.n6�����ģ�f"{\<�T�2�߅g�������Qw�1�K~8���k�Dd!��f��,%��K�6!|ǵ<uuKug�-��wf{�����bVy�����|kp�8_¼+u��0V��O�j�+4��gY��7���k2�~�:����3Χ��b��R�4|�W���U�eH�LW絥�>��	���"�}v!g�S���-F:�u����e򵃆��߆}B���"�m��u|�9�"y�;m�	f�'���xq�,ƽ��21Cw;�C��|����Moj�2@�îh/�>�=���U��Hg�c��v��:�r�|+��z9�5�wm�O�x�V�[7����;A�Ncm����&�rfŭ��'9և���q��]у�ymlϴ3���sD�k[Qi��Sf^�tYW�!����G}��D}Xj��ST ΟI�#H���ƪ�����x�dtn�i�C��.�'1��
�=��i��DN�U}2��|(�����_-����*vٌ6Z1u"/�Y)����o�������oP7A�W�e�":4��D�}4.)L1�	f��.�vv5{�f(�Wy�n[��1����r�Ji\�J��o�[f���o�{M*v1J�Y�/{�h��j�dk�>��g��_G%L���\�'Q���(u�T}n��	Zb�"�;�ǽY�_�����ׅ�.V�{�s����8��~ 1M�K����^��K'���ӢQ�Fj�r�|��.͎�;�(�/��1��f�+��ޜ\�F�e#o���!lt��6��hi-ճ8�!$ܡƭgݵ�}h����3�
����^"��6Τ�*2��mN�r廢��U�q�/��tk���Վ�5l������@t^���M�ۨ�D`���'��⣪�{0�5]�nIڸW2�뫲P�C��	�6pҠ̴����8�x�o�;P���1����S��O���{��W8�`F�Nn�bx;�����ˈ}�{��t�!�'G�c��f;I�͏�g7���z�Ĺ��	�gi�E�t����s��p�Ce+��}/Q$�.wt��ֻ_J�ݜ*P���DD}��<�զgj{q�y���Iu��war�0��ű_f�4(�-�~�$�DD�Ra��aI`(���,T����g��طLB�[/�ݨ��s-�8�W"��o����1y��r{�U�3k�$�҆�(<Wp��Ξ�!��n1q-S���!4��3���β���䒲a�q�I�\EGj��?!�A҆��ͮ��O���hu-輳{�'�[�X� +v42���;�	%x�ZS���T�ȇn����b�yǝ���޾�Y��2wYj�&���i���?eC��!_��]�@p!i#`�}9�e��=z�ݝ喪,�ǮNN��T��=��g4���wo]��N~B9D�t�"w���1�����u�d��0��]p��&���"bً���dEu�	C�#O͐�����w<l�u6�z����#�P�6��ݟxgqU�ʡ�P���t�.�L�a�Y]�ߡ��Kz�ޘ����,�>_#��/�#Cv^��7�_P|�0�%����\e�Cgs9&%��_d���6�\:.����yD��D6�+TR	��r���o(=K7+el��Q��Qj)�y#C(q�x��ܢ�^C����*�=V���ۮ���}��e� R3���fgl3!8��ï&�s�6��p��t��F��V��"#��>���|/9=���,���0�M�"�1a��|�[���|��У\�x�+)_>���\s-N΢��Yu�~�\Cr�N��� ���%��vr�P�|�W�W�
�&/��A��D��3�gcm�d���w:]��jt8����Ub�u�N�<Ne���!�R;	3��&bu�j��ζ��� ��U\@R��/\��Tn�;��)������6��E;��:�K�V�;���*8��v�a /�Q�O:���,F.�������rH��xå�pFF�T�cu���e��;>�T��\�4l�
�a�P��/���
�s�7e�]i(�T��9�=�r�n��T�I�4z|��旵V�A��_kρ��Y��^ѶE��roTu5t��]_e9�ve|�H8����W��$~|��S���aZl+���[7�C�T�c��&�6��,Bi'��~�{��\r����ʎ��=!.�1<��g

K7��F3��p��X�p�N���,���ޓ!���?�8�^Iߎk-`���6d�wn���.5̭۵���r�+G@&L��e1��3R5��ukO�~�z�m���OZL+V+{�ur��΅^1���������u"ƞ:֥�|E�`�Ɨrm�%�Y���z���M+�
/-ebJ/e�� }����C-�S�U�|<˻����
�;��)��熒����'"�R��81�d��9�u��� a�����z^!q�\k䜤C8!"��9X�ܮ 8Ց�3�k4A)�X����� ���%i����L�|7�����rn��5��ǘ��A*w)]<�oz��{�^ �OWEG)V�|5�k�xH���a�Ұ��!�o���)$�[*UVj�c�_<VjH�;��F��:�e
'��+ᥓ�E�ؾ��B��\P�=eD�wc*/JOonĪ}6g�_1m����e�'~�s:���N�Ɏ��~�{ю��Ω���(N�[}6U��7��&��Sp��f��4ǖ)�*aָЧVx��Ea�~�LJ̙�Y�>�p��Ɔ��3�L��q�_�����R�4T5u�����7=��v�X�n��.���(773�
��Y�H6�hu˕�x��P�x@�1�t&-��9���i
ퟹ���P�X��K����O��t_1�;(����/�
?;s�4��%hj8���<qX���S���������
5,C1�S��B����O��ڝ��&\=�.�Q�!��[�!hiJ\�i+��E���8Ue��$j��Q�1u�XvV��i<ߎ�p���5�
�ڰ��'�c�oQ�On���Uc�Y(���V�����ͬ���]�г�����kw���#E��R�ë6�N��Np�㢏>�_U�c;f1�6	�z�n�-��oZ��g��JsM�rn掸�7�קK��d]cB&�:�Pf�2����_L�Ƙ���iq�u�T3�����
���ϵݺɵإrY������O�ry�h��r��ޕ�m�t�bL�M��G�`�W��n��:��T�W]�Ru�鱁̵�u`���1��f�9����T-��&fAz-vu���Y���Vi�/;s��n�lb}S��ѝ��,�!�xU&�����5V�|w�����U���;��]-�G�г)hC��u��	O�Vȶ�f��AJ��k���8������4V�Y�0k��._V-�*X�^X��x��r�n�v����ٺr���{S�2�u[NVj���`�ۦD��늍u�NH��^�:�W4�K�e�Hܫ��f�M��7��ځh�+�j1�_�P;uǴu�&a��a�-֪
�-=�pp��=�w&_rL:}�dF��5�.W�12��Q�`��\�]{Yb$'o-p�����t���8�÷��q]=�׳�����+يTV��:ݕΝ>9fQ����'���օ��������/���Ѯ�Ut���Z�����U�_k��Y��Q���i���DC.��M:Wn�ՙ��J��	�Xv����W/H�9���(&ZV8㬢�T�b�����{s�T���}}����Y�Z�tu��C��E-vԛ\�Kj��N��A)`��0r�:G���`Sg"ǀw0�9'�RN�v�WIkA2jȜ���0�u�%�����\�9�����H���)7���D�g��<���h��J]����(wK�g$�7���l�ܚC���k��N���.��3l%�h�j�K2�����\�2R�bܬ�ɕ		��ڸb�S�Mݥz���h�0���1���=F9ϬV>N9��qL��8o]�-��lqh���R�p���wImۆXbń]V-0�&��kW��^l��!��h�j	6�vEU�zмݘNDb�g�<�j�/T��/��O[S�٩v���H[&�m��5��v�\�ϳ�	�r�'�~��/y"V�][��.�#�;ei�E������\l��XO��,,N��E�c�Os�vݶ%����NT=��dTz���0���:���ڻ�"d\�ܞ �/�
wwp	a�9F�N�t
kc�}����H�f�6
����W��rhNB|��̹;`]G(#�G@="����׿�{�"f�#h��",CƤ�Q�d��"\\D�)�e�$�4`�.s�fh؊\�f���AJH�((�i$�4A�b�I(�q�Q	cF��$Ѱ��s4aD�`#hC&���1�"��s4Q�e$�H�M�)�.h�����㈪J(�Q$G�7+&������.s�&IY $���b(2m&�X,Ls����&�c!��
,2FHM�I(�b��qq%%��Pd�1FJ��TI�f�F��Ë��2�61%������A�d���#HF�\q� BcDT��%���&�Tm��cE&˜�(�Fb�@PU $��Y��rܛ���vق`��G]�U��V��ɲ]&f
�)��{(-���p`뾭�{���2q7a1cqFU���� | �hW]≶�:�g��<#vӽF/N��#�L�u�+	M/
x��<�[�#�`�����uH�p�_�T-��N[=�;������82Oό����r��xE�\v��)��(��QB�Wbn�d>f9�'=7*���Q�G�,e�J���i>�5\۟�VF���㷷T'�O'�mu���_v#�R6ۻ���Oj�"�[�+R]���l�1�I`B1#��k��B��*��=��S0�i���\	ۘx�w_Sȥ�s��V�������j@�[Da��@z������0���z�vB�m�M�-���f�\�í���\As"�:����I����"Ԏ�S���xt�x2嬹�ynħك�i�ArՖ`d�'���_q�'`��{TI���!�kݧzrI E��\^�����l�Z�d1p�Q��9*d��9`kϨ��'���:�|CU�C�}hx'SS�@�+�z�Ltݮ�h�+���]�ԕ��nXZFg�YF��z�9Z����{k 9���F:��x �jm^��%�t-Ғ�L�b=\8l7x�Ŗ�b����>Ӻ�]sREB��w�^�_U����l������<3I�Rf&!al�c�B�l�x��g����k/k�{����*��O�ᒽ��Tu�[�h�/��S*�lB�I��ϗ:ь��eK�˰N�6����	��7k�+R�F�V���`��5�ǯ��7�������yW���P�{�����c��Ҫ7��P;X��A�Ph�2EX!�H��
�*r��pd�}�Hk�@���<t*by�J�dگWfN�r*�_
4͵�W��>�<8���+�h�=YGo4�(��-*�F��O>��.���a��[3qN�Kz��J�n޿2���j�)�/B����f����A���������1
��pc�#��C�n����s�_
�p�!osZ�0�g������H�(a ��:��:zr h�\Cۄ�\KT�Ga�����kɽg:�s��.z�+)�`������]L��F���Qǅ	���-��;eh�D:�/Mf^�c�CNዂ��y �(�( pC����ZS�T�㣫��rЅ� op�͚��jj�P��=�h�G9z�8��N��J9�@�e�@�a ��|�v�k��s$��R{	ǖ��{����O37�ۓU�Ux�G�hg��yly���QSG���u�]BVLM�q��nn�(��kG���&)�[��k<FB�P�ݯ%hn���P�`J�9��:�x����*b�Η7%�i�N����`�ҿ >��
��s��^@����b�51zX��t���O�N~�����u|'I�ЧD5���i�`��3c�6�i���P�A����N,�H�������Z�ǑW`�F��_Tq��z��|��p�$9j����wW�b�1�9T2ju��r�9�
Gr��5���Z,8ڢ�jo&b hƟ��{��9�/M�+�|�0��dщ*�g1��{�V�Ul=����J2�r,�#d3�\���AN�����aд��˅/{f;r0��
i�p��5[��s�&�K�;p�����8kH�ي��p�:���k	�{0I��[�ʮw���9�cE��>���i��~h�Vl·w I���감��	�0˲���ƭ��<��z�1�v+��P�"����O��CSC�����EI���W�e��7�_ ����Ǩ??���:){I��*����|��&τb�mN����qm����^�Y�$�ܑ��7K�$v�$�mH�d�@V��)L�ߞ_�,���;�1�*l��]-ɒ� ��[���t��e��lS���u���i�b��̡�V�xNa�[�f���xvP�c	�U�Z����Χz��<���.Õ1Y#�H7�S�}�Ai]Y����"�9��������u��ݷ���Xc�}���Z�'y�
݁;������B�"M"ty��Қ^�R�s���}��*@�1�]T��o�Y`x\7<��=>�ʦ��E-� ���|�p'V���"m��l3�T&oc�s=�n�O���|�9B�C��|��}�Uc?\�W$�<�wI���ζ��Bd��a��,�ͽDi�yϴ��9l��4P��b���G����]�h��[��B8���Oq�l����Bzy
r���&���]&�܍�&�ݚ���7�<n^1" .u��/]�&Ҟ��7ɳ`���c���#8Fk�[�}M���]�8�X �)�xTGT�t� ���-6/4�f����P�����X������S~�5�\=������?�N$>��R������*�A���4��]�ں�3:�~�VK��F{1Aj���^��#A�{*����(/�z�BY:�d��A�!}/P�t�KW74hg	�"�ެ��kNJY���rryc�4����g]�1�l����|"Ƽ'�����4���:���K��؝���,�����r�Bo��k	�Y���-�����o�P!�X9*Y@����M�`�����ڱ8Y��Tf�Ѽ�B��ڠd����`9t���Lή�n��^�:���N���<���}U_|p�D��/Ք�]�o7�
�]A���J�]9C�*��m,6���1�&��:Z�8�C1�M�+�ju{\�.��z�|�՛Z.d���:���m��w|���xfT\����*��X����<ؚJ�c�p,PuY�ե|;�������h�`�s�}ctQ�ɛ�Z@o�ܻyD������E|ֽ�/s(>Ưl�p�uG��H�`��z�C�������1���xS�5��}n��Uڻ
XY�7xl���j�����^׫Ԏ��j�U��R������\c���{pU����uG(�����j[�p�p9��-u�]�l��'����[O8�&�̵e<ڮ(�-�y̴��(�ϳd�����=����H~�^�4N��Ns�5�=�ݱZ��UJi��ޓ����+�owK�ٓ*H��8��y��������
��HX�O8悓*���YS�h���A�,�vR�uz�ެzz��P����񴵷�rWi3���wy\�h��s�q��o2���J��Ժ�o�>�J7׃��&Qi�i�f���[Y�9
S��f�p	�\������ıD<o{ȳߪ�k>pT&�S�sH��.�����_JאU���k&�+΋�kt�mK�ahM�a[9
Q��@���e�kc.bVU�h���q:�ku�\��O��L5��h�L'q<��@�u��(�C�7���s������'$j��a\��'���'�c�5��h�{��wS�,j��E5˰�����}Q�2V��X�����n�9s� m�*�8���N���Xjs�׉��Ѳ"�T]�&�НyB����>�I���n���J��%�g:�o��kY���F<�Uf�P�	��Q79Q'��x��T�W�7����ݮ
�q�y9�٧�j�δ���N�����ND�ס��#�y�����:^Ѝ63�M��3[ޯ���}Lwt�nfr�����gU����U�����j�6����s�C���s[6!iqTv"ț�^�{�t�@;�Ox�T@#�n��fgٴ�,�f��Oi`]�}ۥ�Գ�(�A�uC�z6ŉ������w*R"L�h�9m%Fk�vek�oDں�R�
�I|pⲒ�|C��ga��|'d��_�������{E����ɠ/�S�ȇ۴��Z�\@��ކ���|�����[��9�c�y���\
	h�T�	dmIꎮ��i=W	�X2嬎Xe�FVu�J���-���C���Tw	�������)��e��!%�I��ܮ]���ۗ�<k�\f��r�uI_���zL3-f`m�����6�=jR��Ƌo_oD9i[9�r��uNi���t��Rk�ZVJZl��Y )�s���\���ГJ�ؤ6�)͹��K�/V�0'X�O�Wo�����[s����Ԏ�.e7���c�ٵ���=��!W7��c�}5�T�~�=�\89�߳��n<Cw��>h���!mIYu�Ў�������޸Fr���!�-mDo��[�؟#�`�Ֆ��J�L\��s1��n#�^89��V�7Q�t�]A.G)��|u4^�+*��ŉ�
��-;
�����v=�/^�8[Mu�t� EЬ1�u�kX�o���6<4�	�ʷ�"%����җ-��T��ı��������+I�\��nHs���A�c{dzn���4���)��4rfjꚆCȇ0���[^�}��o`��휴�;��z�Z�l�;�m�5��U{hj���va���c]���a���=�;\tV4� �x9<|����}�Vl �f�E���v��Jg�Bީ�ʁ)���(��¾<���/Zkz<�ٓ3�eVq����]V��ݳ�.��]L�'�V&9��x5���$����|m=юZ��yVuku59v�C�v��{>��k�Ρι��i��2�Z�RCy��y�}��Ν�9>�kW���Dd�X";Z��aG>��*��*�����Ne{�_T�{W��j�=SO���?���A��r�s�k��o>��pp)�꒔��<�V.׮3j�N[�a�3w[�+��Z_g
����A.��+�1>5��h����C^�ǣ~�w�Ɍ�f����_��;�ih�]����$Ҹ5�.Ƭ�d���:�u�]��I�k����;�7���6�&#��#��xS�U���5�Z�����St��(u6^	n��]֠�(��4/9Ρ�PFW�2����z���d���q�]a������
�Φ�.=�Z�l2:�9;������>�%��m#�GZ��Y�H]P4)���y�:[�d�[Rn\[N�^�t_<���6��q�q�O>_`���g�^�U�"�\����(��j��-	��k�����n5��l�[Aڜ�%q|��hS��a���N<�ŝ�MrtV8s�ہ��F�!U�a�\���\��Zyr[�{�#���z�X���^eGR�����٧�������9��9��ě�Y��:�	�q�-4WnŊ�O>��B]š��
Ž�FOZp��I�F���;����SY'_�b��n����=kbnrxv�Q=��#�@�:r^���Y�$�4U�n��[k���p���G��5��Au{k���,A�VTvc��<��������J���;c��2�c_^��F����EEG �9�c�va氦�BW��Kc���6�:�Wl.§@ڞ�3;�捑��*7p�m�M%vri`[�`Բ�Z��M��]�� ���@B.r��{�g�`�ZO��.0�l\&����+Q㖇���o}Ͳ{������� 9�kgN�ɗ�je����Ls:v�6Ӻm`K0������[vQ��F�ź4�.jo��l�J�W5������ڄ�ۂ������ ��	���w�*	��(!ꨓ�ﮋ�T���Zm�Bء��z�ج��;H��%��C����PGA�mo��<k��7�g��KN��S�s��6^�d��m|���T��aO}�&%�Ǟ��F��.��h������x�z=�p�rb��О௓c)�9�B����4{=��5��mn���l&1$M^�q٣*#�4���8�7�0��@<ȵOEp�r���W��w�5=:�Vc��1�Y��w��h�J��6���fB���Ư8S�Y��)��,���Tk��Cn5�ON�����-�zn��+0�P���:jz�Zy�/���Y�U,��7�y�Ռ��1r�u+��^�q՗�VL�Y9�O���pk.\Fpbm��;�{y�:�I�Z��KV�+��n`ݦ��fV���ڞ /n(]J4���k�Jբd�ӹ%W����ddJi�tMԥ��������9��@oG�R�h<�}b�L�y��.\j�Z:��&�T��Yk�t�No�7&,uv�G�����ir��F��W��'0��c��t.e��(2�r��gq��\��ݜ_�fC������*5�gV��Ǆ����h�N,���ڭ�#� g�{\Ƭ��J��ǖ�GWq��|���+G\�A�ْ��e�Gi�*5AVs`���6q7j�S٫��ú5�9�wYwv���������j�K���#mqU��q5Y{/b����ݶC�y��q�hvܧ�{����. 𧹒�������Үup���۬�7i��7W���G:�N�0d��2����Ǧ��R�$�}�@��A:�Rz2�^�P��^իL�U7��L�D�+U
kc޻�T����3�»�W}�p4X��=��W�F6�;a�g��}ؕ5\Z/����PQ�P԰,��t�K�jձ$��ҋ��w�ͽvm[�Ƹ���IX��.̳B��u�����n��-�j�Z�9̾#����h=.����x�k(RwX�*}�����,���
�8ǔR�*�r��t$=nH	�]�Gn-��#��z�;��#��\�Z�h�	�`Q�h]L�2q,�VS�#(�,����uu-����f�;'׭��Ĳ㊆Iv����N�7��/�̭�U��t��}���-+�A��q�h��/��Y��6�Ӝ�c�\k�r�!�	�6�)ɗ�ڜNVn<P.-<굹��\k4W;]m-¬��;6.�S:&���:�ޣ3pVjo7%���`p���
���!*��KC0]�B^1��
��َv���vqP�6u��	J���;7"��V��@ m[�<.���A����h�3V}c{�z��vj�o�`pA�>G�Y��Fc9�\+����L��+Sy{�ʭ��4�䝮͈	L�Y��>-t���~d�V��ׄ�)�
�[F!Lw!֭�TG����V���\���Q�j��A�ۺ�b��������t��t�.P�1����r�ݺ��J�v=r��{����w6����actЬ��/n�V��[��]Fէm����>E,Mf֋T���$r���ݳ4�mF�t�2/�^�����YȪɝ�x�X�pl _Lz�Y�J�G�HT��_��W1m�n�h�)3��p��:b�cr��`;�t�	�6�L�Z-Y�_1ݱZ7��o��@�Y�^p�(͔�ef�a�e9P�Ք�=LMn��;ţa��nl�v�U�'�t/Bn���Q���WH?�����tż��1z+A��]��'N�����Vd����O�1�]���5�,��ǎ��z�u*b�1^Z{\r>�2��7�+U�]i' ftW�uª����� �4�"CRDTh�	��M����L��iI ��P[&L���MH2lD�C,T\j��R6�A,h�F�
����lb�+���4hHF�Œ�(ش�$�A�Q��1��T�Q��F�IQ��%9��D`����j(�qqX�Elh��8ج��Qb�(�2�L,h6�F$�X�b�Ic!�Ѵ�&ش�AI�e�#2�h�F�5EIl�
,�,%�b�F��B�&��h�F�ƌb#P3B,�QAhe�F�1i1���Ԅ�D���&*@��
�
��z��Ԩ䭵���J�qڵ�H�(*�cfD�eو�4̮�EDv��y_]��K+�Y�O����vod�5�k�UU%�z����8�~_k��g(�/�~QH[���r]{�1���QJO���7t����m� \�C]<�7x;�-Q������xZ0��ʮ1�>��k��79P'��
���s�t���ݶ��;�WH��	u)1)sw���@庥�����P��D%��}M5n�N���jy�&���5;��iYU�l���T����Z��9:3�u�ugʲ�ԩ��aL�����|�,N�~��o��۾���U'���;3G���!�ד��^�tӄ�v�^��-����z`�?�.����֬��3}��q�<f\����MAI�+kV��x+>N����o�c�m��0�t�jnCu��_t2��!o[���v�Q����H�X�}�q�ך��q��M������oI�����)�����IWp�N�A^��A�vYp���Z�/Y�a5[2��m��qXU~�9��D-������$���z�)=x��q�Q�.Ú�jl�3꺾�k5r�wH"j�ĩOS����G����7��ԭ��[�wA�{}��%J�]��wc]j�r��+��|�vF�G^&�6|���c����V��;ZqB\�o� q����"�6��gC{J�p�p����v�����9�O&�V�s}�p�\��n�����K��mƻG'�vD�?[��g�\܄%6m��R�����M[S��:�p۪�ᚈM��o*�^�������!�C�l꼐z�;�ݴW����y�+����yú�V���4��c˙�ܢ��������=��_j��i��T��rz�CU����Ă�Bhe�����f�C2�;p����=mڕ�g�����Vyt1�z��`��@�[妅-�i㯲�O1�_AW0�K��%C�£�ቁf,rWz�f�+��1���ܳ�����н���;� �R=ut0��%g��}zR�ԟy�=~z*-CYm���WMomحg�����8��������}:��� nV���T�kW2���D&۷�k���f��u�+�|�Ɉ7zz��J�
���Ql+���k���;>�����|�j�т��0X�^��Oo*q"�^h,LՅ���;l�̔�dZ�����C�0\�Z����Wڏ������������t�W�[ǡ�QC�M=��P�������w
rկ�c[yg.�Ja������t�l��Sˎmn8y��e'M����m�敇��\:*�(s��]��e����vNH3./6��7f��s��Փxk'��_ޑ^�������ڄ�W�����B�:���U�8�3�)'��(��T@�`�'������/Sqn���󘞞��$����m�v�0�ȕJ~�G`s����㳮����ZQ��_Ϲ��'�k��ƅBNȞCam�8��]F�HG-Ҹ��w���g�aE|�5;�68s_Cn7���d	�T����O-5x�8y� ����z7���]w7�}^���cpjzb�<�!hb1c^]k1�X�Ѹ-�����?A�/�������ָᜄ^�Cw!�(�{_h;�r����&�J���0-��0�Ԃǂ`�|��˽x��Pb�HsX�h�����;��!���.ԌYW�}�[��1�e��l��u74vBW�+p�UEM��hЍJ�`�5Bw�!\���݁��[L�
��H������UW��Q�)	�i��Ctw��H�GEܕ��jjm��/��:;7��559������\�c!�>o3u��eYʏ����?f�^VE�����f��=��Gh�����k^Խ�}jѩ�JP��2���o�h�3��r����-��بZ�_ɶ��=�����t�e$EW�|!�׹+��Ybv��~z�Z�F7kV��M=N0D�:2'��e<������P�����~�ԣ��<���[�]�9:��� .ͻ7������}��A/��
���ܯ��5/����,��o�	�<�AR�T����ͨx�T:��,﷦2�d�ʝ���ިI�l�Kw[|�ܴ��}�{��c˜�B��HР��d�$oUM�sML��we����ܚ�e�v�x?z�s���.�y):PGr��We�����m�>���Óv��E`�V+��]ܫh8�T��e���o;�\�-͆%v0R�B����	S>�39����:�eޞ+�ذi�D�vxeۊS���(��0;��x�go
���]lѕ�˖���(�����
�2��SV{�f 4���Mn��Oܵ��v�w�^:yۧ�c��|��T>�� �P�{���Dv-���h�}�Jd����Q�KZΞܪ��A�1�'j㩩�-<��Z*g�iQ˛@s��Vմ�9�x��CyZ�:6@��U�'��ӯ#$}�� ��;����8�%t�}�S�K�}���.2e}n.��O¨�� 1��kr'�.��
ru��މ�ĝ�.*9Z��[��;V����lmc��2� �K�~�z�y�M�P�}qT_.y�Õ��cox�ܞ�4��
@���;�u�qLd�Ugw����Թ��i�c.V`j��(2n��u���!k]���"�Obփ�zZ�睰VZ/�t���Yк��\�Ĵ���)!h�Q��措�H�^e�~�JC��O"��t�m#�XF�8��=�Nr)��<ŹH����ჷ.hnb�NI��3���t��9%k��سz�h<�\V�&VN��&wt��TDwlLY�9Hp�9�J��p��G��ő��b�[�y�J�6J�Қ]�2��|Q�e'�n��XJ7�VД�i������e�s�����_5������X�dk�����-�aO}�v��'.3���!��ה�Rý>��k��q�opt[ck�TU��t�ͻ�J�m������0y�D���+��6�iXzݳl;c1��`�<szξ�۲�=6�q��,���Jܨ��A�� ���B
���H�΍�++�Ba��n'�Ht�� ��mI�s_Jy=�K���.��+���[�>��1=��#��Cr����Nݍ�!`ڈ�ӌe^9���^M����S�Ӵ�qA����uѲ!<�+��ВW��\����O��i���?s�y�я�ۭp�Q���@�M����B�@럅ۯ���IX2��u�>������j���c�#�4���Q�ח�n�C�=� .��p��w����C6��;=GG�Ec/ʘ�/���9	�]M�Oe����\��u�0�J�2%�Z�M$i{%a�־P���X��H�4e������4�a$3g[������Y�KB���N���u�+\�Iz��u����}�CpО��Ԭ�}P9�ct��OZ�Z��eByuX�mo_,��,d��U�;������0��q��tɲ�������Ms�]���u�.SC�I���������p��%'g��<s��	�3״ew#�6�\:y]5��zt�ˎيE�45�Y/�ճ�Iֆ%����y�Z;#�=:OB��
�9��o���uݭ��� �o�t[]�%�*[5
S����8{o����s�󘝪�ɛ���^���\3���s9�Dv.�Z�i��B�g3��3����)��糘{�z�9qҥD)����|9�໖�����u��{�STWa��^�pkL]�����8�S�W�@zj'��t�T!�ӭ�n�����X�N�m��s��p�0�x*ϻzg�Om��;{"E.�.�q=H���*-�}�Y)�� �wm�T������[�~{^*�O8���q�eg�պ��]^SE�"V��J,�X�>O�u1���u��ѱ昸���*l8ql���Q ��T
� �g����{h�|rн��E�Q����a�^�޷<ϫ/��w����I1M��h�LBvD�!�}���zC���6=�yB�s�rG',ߊXߏ��(;�һ�b�d�����蚮:�]�4�ȷ��Ο��������{WQ�ޭp���9�,���'qA�e.�;�Ş�@��̫>�Uip>+';e>���JH��L�C��P�u��3�Z��[��G�x�&ioE����.�Sj'|22	�vny�ʺ�j���ކ��ɥ�T�aͽ��v�5�VU���3(���y;�	
�ݼ��wޫΨͩQt�T#��:���8��IFK�"�:�&t��'6��P�|���G:�󿰶��;m9�U��=w�.�>�ƪ6��v��ʢ.A}"�'�}���9Q�ۇ���i�t/�ګc���ފX�gs���e_u�
V��|���뢪jW��`'�� �Fd�@�uB��,fl����#nequ43�'\}����b�i��9�ZY���Oo��"���GT\��}*K�m�lS�6tOR�9˹X�����n򱮤�b
���X�ҬK\��Ƥ���޼����PƓ��\��y�w1�2�%�S�amB�Zͷ����w������)?]�Gu�v��$��R��ˎx�c�P�T��
c�ޘ0�KGN�����
.��N�kcE�����r�b��|�h���:�(���홉��JEL#O,��Y�}���~��i&��P1Q���l�/o!�2�TMi�1�4�4�Y\�j%nMF�:��mr�j|7�H����6�r������Mw����g5�U��6>rx�w�B��[a�}�m�	k.��D�M���9���7����Sٙ+\�,�b��3Ω�����W<9��sYA�����q�HgY�3�f)�w�ȯY�_Z@
<����'��Y�狫m����}���ϕY�B�;��cw�d�k�u��M����2�]ej�x��������[|d�i�Y�=���wŋ]���H1�����gp�,�_E����]�/u�·����nL��yY�v�r���1�,�t7"5ԕ��
Ρu۝[v���_w$�*1�jB�k�d�O�^���wo��wI�c� �'��NǦ�������:Z���J��,��i��i��hZ.��+@�e\=웜�)��*&�p�<�cb��8���v㝛Z��c����1�_p7�\�m(j��P��}�=���r+4m�P��j��C܏k�ʾ]��s Y�ޘ8�v�&O9-�R�4)D���:ҳ"�@On�CLs�M>-<�9Ժʯ�@Т��_IU�cD��ɔ2�*��G����Ԟ�>e�8[I��[w����Q.*�y��lk{ ����-W��jO8T�BN���z�6�qʄ黁a닭�]��N+�2�y/���7���8��Z�Y}�[�p�h��
�PWGb��N�Y[���q�9���* ����w�u-��M+5����jTD+"�'qdݬ΄�.�;������9/WѐA}������\�Գ#^ �H����e�z�yye�ml;F�J(�q��+Zt���Iwpx`aM{=�eJ�]�`1.�M��8�g�a�{�O�Ӻ�E>�w9�2�k�l6�<�Q#���n���d4Y(EU1p�w!ѷu{�
�C�0-��g|{[�9(��Ҥ�gn��;������L2�j��\�Wz���QΗt��D�e={7x�2�PD�w��!�J�j�z]�	e䎬��s���L�,n�fԻB�\�ԩr�אz	�2%�K��;P
�6�b#bw�oR@��%�&��$J)�*���p��Rԡ�f�ʹRX�
,�PHd��@��Z��2r2.��]YӒ���v٠���
"���i�� �hf��k�^7�&nv���]}����Kꉶ��[Ds؂π<�.��j�}�M�>#6&\Iu:���}Xn�u�b�R������,���YӁcy�*ͻ2�wj˳��9B`�-^䁢�������J�w�F��3u�+�B�ު����6�%�6��",'��Z-
a��E�bsڒ��s/&�󖡫�ަs��woqs��Xu��\(m��s���,��7-���m�22\����Yϻ'�ڢg:���iV�A�b��ieع��p#�`�	)qaY3�����S
9җ�#���]�إ`;��+�e��-�WM��+�V�(��u�d��D�2諃X���;T�X���U��Z×i���b�uڶ��=�_T�kf�Hv��ӄ���m ��#F�̖��VE}��TgG\6V�AwQs���IRiB�gx]���Q}����lب�A�{�X��:��j,o$�]�aйc�:9>��<w�JNa.����dc�V=0�}��kИ�k̭����v
�F���L���7I<(Hyp�p��j�IpԘ:z٦��LJ��4�ċ�����KU �92�ɢ�,'���6:�	+k0��<�J��N�����&����N+�M����m��1upk��ݼn����QS{�C9	�WY��@�u�7xt�;��Y&��t���B
G��E
�;���)d�oyc�7�|UG���z�U���l��Q�9!�4u�:�Yv��Ĥ��$Q�LY��Q��4�ڮ��v��
H����Ɏ��.h!������T��o+�ul�y�!6�&�S������eG:����G�SKp�i�Ճ��'i�R\� �w+ON'��7��!��#��S��P�o�R�fa�)�uN��gy񾮰$V��jTb�S��Ո�}Ќ�*ws�(�*A�L��k��YV��LM����4���nV9ʦ�D6q�)Lщ�rVR<��AVK�X�5����;��e�}���'qQ��/�t�w��v�7����+�ovc2�0+SZeD�d��Qwv_��'ZX�EZ�XLt�$V����#[9�p�f������T�Z���:��L$Z�wJ[�u�A�!v���p�-\��@��R	̰-s/.ǔ)I�-�Y��O9�o�:��׷޺��=��=������\�T�Q�X(�4l&�B��&Q��XD$ؠ��1��SXKQ��FH�P�H��ɣX�JX؀1��06-�LmBƲX���EQF�Qd�e$��TE����F6�)F�J��m�m�������6"
��Qd�Qh��#b�W��X�A��D�X�Q� �L4Ehɨ�*(�ch�6"�%In.1�9[�E��m�cEF�����1�Y62lDlTF�X�B�hтИ1���_}�}����}���ims������`�BX۝B���Mcǽ��/�5}{�|����#*T�}�^\ӗ�c��;Y�B|}'~䘚�Mƴ.3]�1�lZ�:�R6��d
f���nc]����vM���S��u���޵�F/�돰�H�XmcV�^י�9�o��~��^^}Ե�Do=ܚ{	K�Z���7�eR�W\�;E}uUh��&��7b������!X���^�wT��'�L�Lb�a�f���0OO.ߦ�u���8��v�ŵy=p���3�ٻ�tG�sSUa>�⹻�<��~��6�����Kj�Dk�^V�.�jx��0Gyeo5�>��q��a�-j�v��Y�v���
�j��-eT!�싰�d����BV6z��+��K.O���S|��߫@�<�6�~��m[�ש�o������j�U�+T�[���o/��&��|�q��ͮM����e0�O[u�F���v����<�O%9}u���/�eh���kԌ\~�B�tx�*��U�-T�3f4�[�����Z�hcNn�Bsn�Rvf��d�]��]>T1sX �r�vQ6���"�LvbvdUdm��zB_wL���%[)�7��:Ҧ��Ǭ��M�����n*�:��t����I)�_*}W����EoP�Oi��_t��bw{oom�]KQw����Ա��t�"��oI��KE@O�����fq�8;a�0&�[&�-���/����3�*gj>�L�"�H]_��8�5F�T���M�l=jM^�N��K�a�j��9
��,⃼1�6/�9�bؼQگe��%r���{S��4�N�I��>�n%;"��(`��jĽ^V�u�K��T���G�0�s��k�����n5�����A�OUnnC����z��*q�Z���@Zyۚ��X��o�fa]�!1��9o��`��오Y����V}7�K���o�9�4�xW�dӬ�A���so�=9u��s�ڎ/z�ɚQ�f��f#g.8��N�m��s4��Υ�(gwC��s�*y��:���n�ѯz����u�}�zR�bQ�5K(dk}XX��k]����9�TuKk���:Λqj�3*�P�Y��Th�[s�0GB���{W�_T3��2	�&�7��#� ��
�S�iG$��Ft<�wQ"��oJ���βz2�k{Y����0f����E���Ш4^J�ծ���^Џ��l�{c}�'��v�B��i��ci3Օ�����uD���i�We�د����|��=�ܶRtE�������ݔyց�9�U_V҂�j�c[ǡ������6u�cG�n��u�ν�KW��XR�
+���޺*�*��jh���9��,����a=��mC�[p��	|�B�Kʹ�A%�}���.ldޏ�)ޗ��Vֽ�ѷ�+�aw��a���U]}{b͕���܆u�\��-+��׹�h�x�WΩ�B!d�&wi7��T�f�_��e�חR��o�I��h;b�y&�Kru�B'�]��m��6���� ��(Jܝ�kxb���o��H�$��t�]tލx���z+\d�/�*/.P����:����Jb��S;��j�vz�U�)�Y�,�f�l��8`�h��5�;�R47�����g�r̼����.��X�
�빥a�w�!��f�Nbwq�9cf�Yx+Fl6*��ܭutB�l�B��f.\�pgBe�+��m�	�w�Ğ�K��z���S�Ҷ�K���q��Fr���t�[�DOe�i�Nv�P"�����9[��KyUg7V�s��Ú���yU�ֱ�-u�6G_@�٣�16��OtӇZ��Fo4+u精��9�Lf��K�ҷn�!^w�D���L��*(��b�YUVj�z�xۜ�魟�)@x`��Wa��f��+�{k�"�B%���|�TA��s7.H�A����Y;��w�s ]h��9�ON�����k�؂�� �sZ�uw=��Y��5:����*γ�Z�w ꨒ�eAD}i֮��T�˖���uN������i��-=F�au�U�hQP-`��=S[�M��Ol�T{��RoC��\c��	��U�q�t��k�@nfL�w9�x�]�Ja��#Z�/U-�����5��6�qʄ����λ���)q��SGK����P���0lM����q��z6��6��/r�cR��@�3`���f��~u�k�2�Y忢�p�姎�BP^Cr�D=�)w]Yl�r�8����n�<��VK��J�$FFR��*����w�Q��+
�`�GI���T�3�W9���C|WW�_MC��p�>����\)>��Jw;��kgyr��k��s�vG|�C-k�⺖��I�������\mdq�A�vN'��C4�|�SҺ���O���F��뗎bu~.�˖���w��P����i7��v�B�!1Ԏ�Φ��?ab6�r����Y�	.�������4�N��14��w�N�#�k��Մ��Oq�-)C�[��ϩkܚ�x�z�־E|:P}��z�u��9���L�q9��W�S������ۛ��b�l��yå�nq���������;~�ؚ>�)zii�Ygޤ��މ+\v�{)�R�T���|��va).�n��tw�5�k��W1�?�V�|6ꑠ�U�=�_�o;Yr���c��u�Ψʳ��1�_��K��GE�酴D�W*|������50�K�t��^���Ct���K�d�A�j+"�����n<�ҳP�R�v�\�Ѩ���:��.u�ha|���	����fc7��D\'�j�����czy�����YZ%�'�*u�o>Л���7����',j��Օ���T� 淒/{���[�P�l[���U۷�x�:��1�PU������v��˾ג�Թ<�������%}���{)���Tf��w@�޸)ƧۯXୟ�J���Q�NR�*1�oCx�<�O\U���\���+5"�y���tϑ	j��.�T�w���OW��k.�&�S�j�i�>�[���j��aJ�zJ�b�	uvR�/��-W>�WX�(Sj���l�f��
�W~��*�����ΆK�P�nP���h+o3Z�^p��y�#��s6�Ժf�
c�.���L腐ZB�r����\�v\qJ�q�K��_q�	��(�G5F�����_	��o���yv��II}s�ڝ.A�'�k��7���E��J�]<�"�¯F�d��E����<��~i	㌮r;|��K9�1��7�cE��7oV�4���v45�F@Ӄ����V�ǹJ�E}�b�qαԂ�����Iv-�r�Z1���j,��C��8�B:�iʞ����y�^�S�'p7bX�l�n��!n¶��9Q���J�����5��w��ge��;�7�u\��,��9�9�4����E�[_Y�~���=v�<�3^VJky���*!'����Dl�֫j��R�S�����xn�X�=����uK{[n��' !�9���I�޸N�]�rq�d>����ish��ۋWn};*�rǺ�F�1����)��2��ފ��#��:���fƽ�9�]���Y6���/C����;+��8��jm���؝����n��new��q�P�3��{5��!��}i���:�%�V҄�4�Q��Z��v�3v�au�����woǛ�5���8�"2N��֤�����Ɲ�ys�%��.��!��	W|�O��{e_+�XR��=B�Ӆ�yã��{�B����'����5.ʙKw��ޅ����q��PS��*��˅qs*��#6��>���O����rƻ�x�S�J��?w�;.���E��>���Ed��V�T>��e��3����+:��7�;���8:�d�w!�:��а���$u�RܻI��yCWF��!0��ڳ�:}ζ�]\�<N��i�i���y�^ {+�`�Q�J�wq6cw4�Uҩ����^��l��r���9i\3����T���Gr�8�����`��<���٨�Z�\���M(o�A��fL��e��{;���K���2�A�2(�(K˕��r�Y��&D���;����	����\h�!�ʟ�˕;�+q�K7�
YC�@}֦s1���LO6�]�3��f$k��"�(��'n��g'�bP�76��z���7>���N��e�:P��;M�V�7�v�\��.ؘ�K6���wnZ�Z��Tuv��ME�[H���=���9E(��P�ٝ��ƻ\'�ػ��k��Vj�x���U9t5�[�1r��f͵v���_Ti�@�H\�&�*�;���p��6 �@�(ȹ�����u{��Hjs����r�f�'�P��:���䕻f������)V�e��OefĦwr E��p�v�$�HuƲ���܊w��%��&k[���;�������c�@"���}�;��o<�b��Շ)��±�F�'�l��}��G+�9p"!�9�5��w;E"� F-�3��թ��Wli��%t
�w�k��SM[�ͽ�j��/�Dd��"5��ң�ڳA|+��u���m���'Ԯ�*���sϲ����h,��,DO���ʁ$�S�9�����EW�]SI7��5��m|�{e[w�#ifp�yJG=�� ��#�����R�	;�o��ڇ�ru�Nm��D����jru���~�0\���տG�_O|��Z8�Jޚ��v����$��r��y���jR���O��-����uB���wv�EԾ�m���ӻ�N <֘���snP:WT ��R�03���P�gZ��Wi^�&��\�D&�;��#+�	��8��?��M�^�IR���>U��=U2S�����}��o�P�Oǂ���/*u�3x����sBo��X�S�y�*����}s���z�����ɸ;��]L��2`��Y�kEE���W��^mJ93)p7��\�X�����V]L=r��,>7yr�O���M���@��L��p�����_v�����g�v�1�c�9�L=��䥤S`���wsk;u��+u�dQ�8523b��-���g�4ww!rZ��g�k�JE}7��緳O~J^�p焩x'2��(�`�=�5 �9n� �YUfv�]�}7�+_ju�����[�N�:��=�uij��?�Z�5GkmD*�u�fW�\<Ys�y�<a����mb�*mƧW��{_�O61�>��]��sά�9�]�W{4u;�����4����R����GTLT$��:O�Wn�7����DSûZ���M�g�c�>�`�<�شs�:��n����ӽz��X�,�X:�vB�9t����TE�=� �#�>ڧ*ժW����n����L�$���9�9��Mf��M�_�ZO�|��w]P�l����Y�D`�s?)ո�[�:ڰRz6��{���;���!����OE��}����m�OF�o���=�p�>���D<g*%�5�#��9����s�_]d�W:��!�Y��4H��,���vΨ��3��4L���@J��-��]� ��-�5��8��ϋ������r�O�G��2����nF��� 9�\7���IV��ʮ�x�6C;Y�ʛ
�v�Q�p�iӳR�`�Z1\��e�Բ[���;�������#���Sk]�}C5@���œju,T��a$I!�sE��t����(�![l6�<�{)���m!]1��tEL�Ί`��=�v���rk�v]����H� �\���gu��$���z"��̧n�Yk�7�b���=���u�;5k�/�U�<tVws�WJ���!u:��_s%E��O�@�4�ed�t:�%�S�(CX��z1 �ҶX��3
�9ާ1jl^j��2�m�Y�Mĥ��
ݚ
��o���|�����H�fp1�Z��y�m�����.��%�{�o@;˫�m��[�{[��WJ�eg+M�ƹ�񌿲cǠ]�����(�]gjVj	�X�,�ΰWH�����W�zxu>�ٳj햡$��#j+�~���I����&n`:�|T�	����X7�u�R=ڦ�x�IV�����Ŭ�79r�{�1Q�p�r�+"�N��]$W��SH�_Vå��O��镣��K����δ�	�:z�*6�뼕h�cnas7�V�[CAU%�^wr��(�ӡW0v�N��Kt���4�Y�N'}��wv�j�� �,&�ߦZ���"F��xc.�0��H=��*3/l7���i�uÂ��C0��#t�k�FJDH;��Z�����+B�lbYr��;��1=y]�i	����b��I���"�
�܉���4})���V�t��7��r�"{E��x!j+�f�ǚ)�n��F�9�ͻ�+gwi	��3�������)ة�Me��S��fSG��L�9��ns�J�k�B[ԶuoY�٬A�MulХ*v�cZ{-��l�ut�x�EU�J<��D5�x�������d���N��hpjU��̢�%êX�[{�h5ļ���a�H��Ct���-�w[��P����ƙ[O]�n_+��Zz��y5a��	�$�������4^U���Kڜ��vp}�Xi�����Z��h>�_5N4��ąm��;���n������ )��ۑ�r�T�(:ܷӪ+�+x4���&ܮ���+B���g()�
��3�P��|[ocF��}6��.m[F�WA��Q�-؄Bb��T�˲S����iKc�]L��L9�B��0g}X0-|a��tA��|M�N�}��4L�ݢBA�w�o�$������r,��>�C�3VG���te��{�gkB�㯞�l-ԙ��ǳL��m�4N�in+�۬���ڡ6�8Dͷ���+�F�'e�. ޔ�g_"���ͼ&��9��-��d|FڐU�ӱy��:$�M�C=�V��7�����!`J�LX��T�+Ð�{].�E���w:�u���׿���F�d�Z4Z2�$$������e��b�Z"J(�M��5�cF�lT4b�b��AQj(�R�,m5b2&�Q�DhX�-��`,�F��cb�cTh�ţcTQ���Wl�(�#fkDE�QbM1Dh�	D�"���+Q��fX�m�5�Q����̖�����E�e h�)F�1Xȑ�Tm�5���8Ρ�^3��B�7����=��pZ���u�h��Ԉ�;X��v���
���۸e�'G�ҡ[���E���/����g���浐�`���2�
zB�r�¶m�B]����u�p<�P�{t ��ޛo6_Ű�Ș�H��7tT��kV�J� �Q�'�ʗ�(n>A�_ڊI0���k�sUW3�b���kv�s����an^}<�j�os�ɪ-&6�&�u	{�g��*x>c6��ΣO��ƭ�䶖��T�7dJ��l���L쪍�c������e|�Jk�o����xn��:~��f#n�@b��,��p��mf���+�O��y|�kO���ם,�誎�)B�ܽ&���kF�;K4nh�Gk��Ϡ���}��s������Mvw��z�&�ܮ�����_MM�÷[oc�n(��5��GF��P
���ؼ�k3-�v��;���UK����	_�e�����jonge��x���y�[�Ɛ89��[j�eS6��T�1�[�3��<�Q�܎��ҡZ��D��W��10���h�Ȇ��GL�&�]g=T{Sy͚=�uu^]���)�}�Ssb\�*m"5�V�;q���ؕc����ڌ�(�R}]/���B^i��T�����g:sZ���#$�u�'�b`�4�3�bGd��/���kn�k��n1�����M������*��m>�T��=p��Ӑ�j<�f\jOo�p��=	�NS�b��^�w�*��d�;5��R�ɂg��\!-wSw:}4[쿹c\�^s�r�RW�S�vi��Q�aZ��xD��gp��]wWT-}��l�Ops�r��!���HqO�7|�ޞ5��	�Q+^\qJ��ڈI�a�~�c�2=��j��n�+��[����.g��h%k���5��!�N�7��j>��qr��n�yGwK��G�H�L*C��:��%nI�r��e k+�q��2��Ӯ�VڣKM��q�V�"~�:E����	r�f�Q�V��ܘ޺+�W�4/;z����*�(u�8��!�f��Ѹ�	DK�i	���Fi����Kuդ��\�t�Ye�`����:ԱV�$bS�*�FИ�)�fn%�Z����:�m��҇{�+/�f4nKK�-Yf�����9���[�R��y����Y@�(`���ef��Jg{�g��0HH�WR��+R����:s~��*.�ʼ|�b�����|/��������N��!!n8m�r{�w;�+��]��Fb���%`���;*^�X�Ќ�׎&Yj�j��W8���;�o[V���eAW?ʦ�(Jc�W-�V/to>���W�t)��]��3��E1�PU�޸�=[J��r����+�p���"�i�^kX�#;΁���U��C"j���̔����Z�X��C��\&�\���]eWՠn�ӳ��T��#+sqN��:
�	=�bE��T�ɽ�����j!4�ʶ��j�r��u�|:굶�'`)�
��.����Kf����5���Ntu��V5���i�N��S�aO��邠�����ꅯ����y�=$�b;^�1Jqt+���Kp8X�WΩM"|� 0`���s�ү�z��M졍�R���d�4@�ѷ,��o)ϭ��U�;���1>�5߰��p��L�)�3�4驪:ݒ\��D�"blR���qVv·G;�s��Ņ��Q�ly�z�Ce5n@t�U=��S�$�}D=w�%��L���}��S�{��dܭM�����%�7��q���m�#JZ!Lt��	O���Ήc,;��=JMc�uxm%��&�8t��F�U!=H�|:�>-��2�1�B]����ӛ^2b�k&�V�w0��;�15	��#�?k��ˤ��v�:�o��{Y���$H��&�=����wå�
�����r]g��aA�ζ��r�t��y��{/;77��W6z�M�����s��yz��c��k��7����E�5��m��X3�8˭��9�ʐ��i畽���q��MIΌy���ֱ�C��79\��fEql[��Z�ԱeatO�;*y��������g+�̨�*�ۖ�w{WA+������Ph4=aQ����$���=���*γ�Y�̈́�w2�#R�������X$߶�%p6z�������O�繻-d��%5�<��p�����A��<���cM�Q ݋ԃ=�z.�nŭI�f�77��&�hZT(
JW�z/B.jegdq�Q�	fM�4el�=H�a�:9l�oÅ˾s����˟���9Y�S���O3����y��we�_בkвS�hO}ȅQZ�v*�=յNR�+����7��1�w�
��j�D���u��V�o�Z�P��F�����	-�<�ܢ�T+��Nt:�-M?��{q���o�Rt������F����]|:j��LH@��ꫴ5��d�M�����=�L�ng͌��ĺF�
~ﷄr��qUd��E��Bݧ�u-��Rҿ��k!��P�;N��"u&��R�`�On��*�q��`��Z�]����/�|�J�U�g��P�M�䧹A/A�O�V�`�sR�'�>�\����5	&w �P��=-���5�h[�hHn�H�ω�c�����=��s�~8�^P�4�W��ZUX�gә@�xz;������Uǽ~����_w����������^Y�������}E.ͦNB��3p]�S��>~���}�z��H���^��e�G�3�>���l�u�Z!;G����7��4�кzeVc�/K�� ��-��+�b�,�\�n�N�7�V�x�YN�]ǻ�''��!��0D�|�I/��5�RU�:��8����%��Ǹ����j�-�Ys�Z١6����{�_Syթ,+@ѕ��Y*s��{�c��ΧQ���z�Wx����'�~���x�3���k�R>�r+0v��_�c�!�<��\�sau0*��#�%��x�,�~�����k ���z҉u<4z��nk�gË'2���O3�r���r��φ�k��\탎�2�G��h@;���T�w4-4)|����ڞ7gĥfa���e�tyj��φ��F��O��j���NP�jg�l�����z�����v�5$�0�X2��ϙ�z����}2���>�s-c�u���mO���Oi>>��P�9���Ѷ9e8��u�'�`\@�k饡ʇng۔O����?w����G�|�Պ������#���t�z�ڮg���� �,� r���PUs��݆r빯PG�����K�lz��#�'g���98v���'<��:f���ǎp�v�N���y~6lD�L�I /)��e��ԇ����Ͻ;�����NJ�D���<����ƧS�>��*�%����A~�G~G��q����8\C~v���7�Y>}y�?-�(똑�����	��[chm9Q;b٬��w7m�F���I�:�U�Q����������z�Ԓ�]���䄧6g�}8n�4��P�w[����=����iZ�G{fJ����;a�������`ޝ]Br�{/;�L���4�i-D�#����@��؃&��h��Ĳ}2��G�����7G�=5!��&:S4rw���7������~V�������}��`�5�N�E/~2�����s�����w}����sحk~rq{��k�v��5Ryl����� o����2k�0ʚ���T�U���w#�����oc���q�Wm8V3Wi�9���}�"��߶|'����l����Bvq�"�6�_�7��q5�"�f��j�aȧ\����L{:�ǃs��F�P�K��X+���?(�Wu7��2��R�p>v��q[���q�~��a�e{�Ժ�uu0��;�.}X	��y���0�3��z/$t�/ه}���f���O���]d{UvS���*z6�\���̯W�3#�>{7�	�a-��x�D��^����js�y��нS�v�O�q���YFuAy&^�T.�oQf��_�Ӽ�}09DJƺ�6�_��y�~Z���e�S7�b�d��eǭ5��is�ʬ���t/)���T%����a�z|
�������y�y�{o�c5�fx�LCNuWVL���-�i���p�(�����l�ᄉ�[� *|���ު�A�t��z�f�A��V�du�����bUܩ,��}��N�����b���6������_+v�>��Z7���k��3Y�n�Yٳ�'PQ�|�a�p����n"`�=��jS,㦪�W�b��������q�{z�W��ڏ�2ڥY�)�م�'�G$�|�)�jz]D�ݼ�@���н��V�N5�s�7#����v*�=�N�'M�߮=�$�� r�0�L뉲W�������*
��9Wz_�O�.��ar�Z���8��o�ԇ{}R6��ݱW�9�� 55���?Ku��|}s�zu���8��BW�sM���>�����]�<oO�{��Őh{ޭ�������zjy�d�S�K�=�V�ߜQ��)���B�S������Ƹ���M�O�>#��O���`m�)\��ǲ_�/#Q�����D�V�f�ӕ��K�З��[��o�h���{�߷4�Ų|���ۛMk�$�8N���>���dX���+7�����1����=�T��^�]lG�焵�+�}�Oz�/���>%E�{�wL+��[��\�>\��Cμ��}Ό8�y�~��cZ���mHf�M	�1Ą������sz;��i{	ө�
`#J5i �<T#;�1&���1r��Ve�{1OЊ��������b�w�m�[��q���iG�
�	:����^�q�Z>��eE�r���Qf��B��X�(J{�����[�N�_9�*K�:D���Vu!ְ(�"s�GS9uw2Sk�w
�5n8z���h�W����v�D��i8�xw������}����䜸��:v�eᯏ�C\�ީR�.�m��Q��O�|K1��wڇ�=)���#~;�hn��MǪg# ~��^^��#�E�����ޱ�JK��ƺ���̰��~ӧ��r=t�{":���Y�3�.�z�gz�Qܢ��ۯOE�����S>G��e��A\@�Lb�Ln|�O�H��뭟gM�xYuM�g����dPn��GI:��~4eSJGb:�)�ǖ!��z�q�xD����Sz�����dzh����~�=�e ��rY�x���0�)��e���q>=w�'*/ �e�_g�'m�}��g=�������~��N�#�k�&1��߇��p�_9 r�����u�o|T�O�����6��#%��3�f�g޿+����l���z}�l��b��q�&�PG6,��0XW��Ʃ���s��]h0(_#-�ʐY�m��ί3�r����Bv��Ux����wj�{��O��s�W�$����Dĕ�4.����3�����ڿ3�O������Tw�̊�"�dp���L@�J���a��]��/��,�)��+��<�t{�����GYX��`�vfA�S}��OoR+=�� U���5��8�}q�R�����7c���i2�a�ݘV�\�V����ej������y��|�-�L�w��<�P����"dw�D퐥�z���j�u1�i���C}c��g۝π��[�^ݺ%�9�����]L�:��1�c�"�ڳ��3n���{�m�3��wl^h�ʎc���W&�{��~��>`��\�*�~'_���2�+>�a_�/P@�\��?/u,Z����>��=��������6�P����{�ţ��>���/Z����74�fvnۛ�}�c}Y^t�i:o6{ƅ�uX���"�x-��4����~��q�l��-�>�vg���}���F��e���·u9G@�>'7������R�{<��|V}�U��\��П{r}S����:�L*��<<Ng�1�+�>E��ɭ6i�Y�����0V�ib�;��EK:�:;��N7M�bqC)�_Q�-�GY��:גf��DwXR�GzFO-����>��'xk+k�z��Oz�&=T�ѽ4�o;S��t��2���]���~9�=��r�ŵ��(���<�s�i���q��~S�^u��r�p(��s��İDI�7����G˦v���F�egt�ڝ�M[��-�o5���`��Ŭ!�ɡh���t5�-=�P��U��8Ӝ�Fiͣ�h�F�;ɵ��ޟ�Z!۫�J��{WNi�Am;��*$
�1�*�r[�V�$���;݅T�{��G�B�;/@QNb�uе����K#i�:r��4���d�K^ތ<���t,V�RW�8`���ѯ^��Ư�v�(V�hq��ۊ[�V덄��д�i�4Ԯ� �>�R]<z/U�>ꭕ�G|����UcUd��L ��==Ig�k��H\S��;�md�}�y�UY5,L�&�FuKv�Yu|�j����ϳ�,^
P��۳};�b�q��W���Dre\F%���r�h�u9���\��iN������Dmqi�oS���m����b� N/�V�&�75�f�6omJ�Ll��t����־i.���]g ��&��J��@ť�5ݏ7; }j���������č��R��pU>�IT�u���C��������뮆�(U\�ZN��ׄt��&�h�N������ogYrH��<1c�ltL[���-��z��l�Y��o˛��f���۱6��GX/W��vM�lh1pW�c��;C_���vyڀ�k���T�jk�|8�G+V�s����0)�h�qmṀ��8��|;��-
�{�n-隴'�A�j��:�
��� W�PԜ�ڔ{�� �*m����ט6�f��ūuRnХ^��3�j�a����a',T��Gu�i�M,љii��eB�V�x�V���B%
Ozs�VH�|�un2:�uӱ|��N,l�@q�����|�8�J�s���0ȴ��|vs�*hw�-�
P�u7��5[�_t�r]]l�+�j��~Q[��ԥ�B�QٯeI(y��0�8(p���ӹk��ʹ�T�^�&�h�REQ.��Zf]��9[{>�'lm٭�N�f�2\$3npO1�GE��޴���9�\P��q��w�aJ��T00���*4ܼ���,3s�i���oC�"��f��vP�E�ݺ���-He����=�$'Z2\ʶ�ە�.+�Y��8��;ʼ��A�Ú�u��`j˕�8V�=���
�չ�����̕�P+m6b�t+��T[]ܭ\�n
黂�jڂ�5��x�j$�h���eZX4νh��Dr�k��Xsz�'$�w�5��$U�U�3��ao�(�]�X����Lb:U̢��,��n�E�.���k��i#�;m�r�r�%%{�j�{Ϛ�*��
�mm)!7�d�t�֙�C�^�����Ω)?�rG����CGh�Fʎ�v��i�����7�����1��:�TS,5�[J��x�>�mAsv��4t�(������]&�=yӹf���SCDJ�����9ATbo%��7/*�CYy2q����1 �n�!�2��(�z4�ې�\�.M��m�]Gψ�����uB���B�6Ʊ��`�hƠ��k�h�A���cF"���ɨ�llm�Q���MQi*4�E�lV(�q�\l`؍��Q�X�A��jqͨ�UpjM��DE�Rn.(э�؊���%n6�Fɱ�(�%�5F��Z�F9ƣn*�����>����5�v���{�ȖZG���y��X����Ŗ�O�_R7�ࡹV�<6�#�4�]#݃�A
��-��gA�Gi%�u76翢�EL�҆D,��]9�[���GzG���,�ǵ\>�Mo���l\�g>�U�Mx�o%P6�>��ީ~>�y8^�'��s9�'��z��^n�{χU�w֧{�}�c��g��@�F@��}$Y+�q�P�ւ�:a�w�ã�����4���wo�}���ۤ�W��ߨ*�'���>��D���h#�}��(s���)1��lz3_+��Ǡ�ԉy����7�z��z�jϦT:zH���z��|v�{��ו�Q�ۿr�;X�o�x��
�����K���=^ o������xQ�~7������Z!h��4���UyB���kv^��P���p�_��q�z��123z}�&��*nB槝Z}��f�o+�r����'��87+��
�Wi��z�H���4�|�ǽ{eTg��6��f�_��s@��>K|��=�Q���O��V���c��x<1��dk����i?Y=Orw�$ʕ<�KY~�{�`���N�>'v��uwL9����փ���`�:��f2���0�Ӗ�~����{|�Y�lu�ڭ�;{��:,�/
TF_nѬ�W9T'^��t��՜ܺT�����]dz�T��Y�1��t:���!bԛ
q0��\�Sa�bf�h�r���j<0qӕ%�;%����{Gw^F[
�-�Z��ʱ%�-�߮�վ+��>紅��H�R�ݳ0���ʡ�eV�5/ī���^�陷�g�����.%�^�����kS��B�[�f��>'b��0rF��j{E:�<��3�,rˢ�.>=.���6ܯj�����}��诱�Iد�d�����ɏY�;ccʗ.t3�	��g�b���B}7�Vw���$��>�~��+·���=~E�u��aM䅝�{��,Ւx��bJ�::��Z�kޯFŏ8����:+���T�������s��
�Gw���Qd����%Q���ڜ��Q>����B�^���3r�����s���/*��a�y���e	����d�����bÀ�$⯄��:���߰���aw-�xx���iz+ޥ؆zv��lC�!��{}R6�wlS$��@H�"�[�VBjl��+���Ng��y��h�u�߭�<s��\mh7�z��Ug�_�d�����Ŗ-�}�VԸ�a��u^#�wZ*���tnq��>B��W�/�ȟ����3X9�E�T����BU�u�+M��^J�n��6����f�/������S�+���A<G8�y۵oqX��!�����~�+�%��~I|
G�<��q<0T�}�$����'�2�az�����X۫�̆����D���<3,>G�f�nu���D�q���O����y\!=;�E/K©��4�1��ꤊ�z�5�z|#}�7��-�A�Ȼ�yU����$�x�C�=dT���6�{�f�1�]�a?UH����Ny��zUW���,	�o4X��ڦ
��-���C��i���<]xp��D�Vw�U3{V����啘�y���}�5����Վ�����86s�V��eգ��F���93���'G��u���u^�r!:��9�;���e��s�r�|���^VC��x�^#�p{l9��ъ�����,1'Y,�����hy�&wǉ��>�}�Cu��X�5s9
׽���.tˏ7�,��a-*���)͙`+���t�|G���c�q��N�ݒB���8�Ҽx�{����R���� �.*g��[�ˎ2|/�A��.��+�J��uDc�v=Of�����E:A��5���YR��g�<?2����R7�u�O<��Y��h3^$�xW��[u��&
g=��=��l{�:�A���L�%Q�p&�C�[*2�����kP���z+q�KL��OV��b��cҚ]��t�Ī���Y�:2�*�l_^�+)y);���k+8r�Uڐ�P�n�s�h�nk���$�u��a�����67��p�lf�>8��V�l����9ܕ��.YX蹁;KS
u�ɍ{����u�N���y�o�iQ�Dk�W��Y-� r��,	��}���,	��4�����J����)l�h���\W�ԑNg|W�=�:U�}r6��U�7���z}C׵5��u����zd���6�C1h��H,�^��gޝ��;��o��������� h\yo��>H�D�T�zQSSB����3������j����Y�v�^t}'M���u�͎[���Z�H�g�����B���iy*��i����G���h�M�m���[Y~����L����7�TX�RN�!i���s���v�<��s�]�W�7�s��O�)}�:�7��P����q�2�ɿ� _/��l{L��ǫ�W�S�^"�2��l�Nw&=�^�>���s�9�u��]�ϟz����u�]�m�C�3X}J/�sKB��rg�=I�_�4Y��|�te �����l��}{]C����a�~����w�����S��������8M,��>E���A������(�4���WD*�;���^�ޥ�,&S��?/q��O���y{�ޗ�����Q�)\��)�:�N�<w��Q]����:�-3�b�J��Y3x<Z�fq#�Q�8o�f�Nm��^R���d�g!J���S�����-�߱Wt��%wҺ�N�������C[ٖ�VC�͹Cq��m��u-NJ���myB~~��1T��9�du�"|�Er���r��4�Z�*�9\�w�3D+]��8W�=�}��?��G���c�:j��nvp�T;��R7�[���[�/׍��B����{����zu�{)�<���:�BᬩG�<w�+ƌ��Eo���ǳb��I������󻇐;��;�<}���}�^���x���I��ܤ)�Ix!�f�������u3�J
�g�Ӛ����/K�������J�%�}��_�,P�PyU+ɯ`,�`���2���@�>nPȅ�O�=~�+��CB}�h=Oy�G�N��^:�p��G��7;�;���h�Q�P@�PdL�I�)̈FXW��Zz|��q��*�f�p�+�YW=�~�zMvz���PT8�♁Љ�D���i��q#�Ep�ڦC�5���˳=��}�D� zpx���Z�=q5g�*���Hȗ��9<��o��ˈ��C��T��|���i����W�/ޔ�����N�P����2�w�y2w�zv<;^Q9U}�A��� ����4����Y:�����d3
��Ap���B����]Z�Q;5y#�tDhOee��ǂ�`O��7���˥YR���y$�r0kmb9�p���e;�u	Ů\�X)�,#�������$���XI�g�x��v�>g��{K~�<��U%�~&���@w����>ٓ����XN��2�R�W�8����V=8=u+N���mz��@s�����ZE���5���>�!{�M<����o�O�zg��%W�&�Z��N�Nx��ަ=q�w���vG�K�|
�qM��ޗR�u�|3'}�U�W�E�w�8t2s��9�;���4��A�k�#X.׶px����k"�li�eo{G�}]zCu����άr67؜W�V�.����GYG��ia�� `,�(͇\L窧W��K��� W�ڲ.W�{�w�Q�N{ΐX�օ꜓�*|K����G���W�3��U{�o�w�*�n:�@l�����-��{�����hfh�e�c7'a�^s�����+ە�w�M��^3��L�#W�%�C�U���^�'��_�g�������y;�oOF�B��sҏ��2��}$�>`�R����S�x��[�_���z���]��}�9�x�+U�Y�|߮=��u�1�%��x��`_��H�>�����!>�հ���DR�M��R�8�gMѳA���(|�PB�d�(Wp��,���
��6�x�a3���f��L�|��.��n�*�%����D�;�W9x2�.�Q��s/��
�nÒ���&��k�L'��}s?$zh��u� |:�����ڙ�s��Z�ٕeŖ����Q�{�{�8Ǳ8�4;��ȁ�|X9i�ps���VN|�Y�o�1�f1��ڞ��Ѽ}�'qW�,C>s��{a���o�ꑳ�'\�sP��@�LLҜ����CT��z�3^PDv�� �g9�����>���زG���=3~5�C�%�����Sg��wW�|gg�rH>r�eO��܎2�m�m���~�"|G���/��L{zB=^��s��3���G�w;;7f9\X=�C~�J�K���Dz��]Ʉߨ�}�8Ecv��}r��3PI_��&2<��k�Y=C&_�}�[X7m׸�F�1�]�`}�y4�d	��dw���v�#�·�o�~�=k٢�{&Aߺ|J����;��yf�i���b���;�y�T�j�#�����d7U�/�#ƽ�A�ϣ��j򐹋��ǿ���~���.7etE�]zrz;ۮY�L��Ӌ��q���%�{I��ü�c��'��|;�s�r�|��ѕ��vh{�'kع��|vx;���H��(����\{>�=��t}����%�/^��ꮊ&s��릞d��0�->��X-��U��G�[�2�w�~�us���:���agM�3v�$�w�c���\ʇ+ZKvQ��������f�-=��dN7cR2Iǵ:�T��)�W���Į��K-���P�����8���Vw��E#�d��9!ӻ�9��y�Ӥ�pOuO��N���,���4;�x����ՃY����L�6��O��c"�ڝ4>��[�g����Jg���n�/ t��φ���ϾE	*��#V{k��Tm�\`�?R�S�C���p�T�vx�0�AR�}S)���
b��ĆFz;�}+��u.�t!xy+я���r#}@{���qsr�_��IZf�0�1?6w}!�y^!8�t�׺���w��;}qW��~Ӑ�#�{#}@>7�Dm��߇�%�9 r����!7���FK��YI%���\��Bڰ�ϗ�W���}3�/N{�p��T�O�q�d3��|�����o=�l��:��C��p6�C1h��H,�^��dzw���ޙ�6">,;���+�ݟ����l���!jD~���B�w�A��3�,,]R3~I[��̙
��_�q�{�g]�,��;�V|�F�t�'�'����B���h#�%S���ۿ"�M�r�n���+��Ͳ0y�]ȸM׉�x�������A�,��C�g�QQ/�p���ѣ9�F@���7>DA]���2;\$�,︱�����-.�>Xx{�m��g�J��*	}d���9kln��8�*�4���∴��z���&J��+���j�A�-]3��W�yX]w��t�\�ly��Y]O�N���ī+[���܇a���^��u\���=K�z�g���eH:�Ī���^���ޏ.y<�%��:��Q~V�ۗ�#�r���:���7�8���߶�ж���E3왷95)u�c#TJ������g�%����YLm�J��7��oW!��}dx>�[��<����[���3&�Jg�/���� xpx��>�l�w9GE�U��],
�uǇ���xG��l��K��Y쳩��r�dVU��L���GZ��=�Xh�QY��72<�r m�Z�W��S ��y�� ���>���y�;����vL��wxe:�R�L�Ċ�3ː�g�~��)Ӽ�������_���}/ޞ�e1��<5C��-��G�<vJ�p�_DyO|����^��^F_E��:;�y�{No�x�w��/���[h<�gr}��]�Gg��^vn��s�8��C��n|1eԲ��
�n��#�#���ίj�}մ*J����uf��z��
O���ʌ�E`��C!e��������}�CBy�|M@U�W�-�&�~�n4��G:~} ���R��&:Gi
�3Xܧ�w��I����e8�2ݐ���Z���Kw���,����eu�p�F��^+�/�5��,�Ljf����G�,=��輸8ƅ��ǫF�7v���d��a��v�p��5q;;�f@�,҂ @��H{��#,+}�A�ح�����j%�����x�3�����z���^Ag<Pfs_D�"e�j3�ֲ�o��w��X��R{���D{��8\{�v�A����'������ә�ʰd6o�aP�!�j<�����䏾Gx�ڏ34�GZj�%�ҁ��z� �c5�TC�`�B�s<	&���u��sow���>98
s��*[;F�t�7�%��C�oe��7���}�61�1~^#n��y��ɓ��0�n}<j;�9�W�1��Mut:�}�"�w�����O���2;e��lN�R���	�'{e��h�|KB.G1����S�9떓�3W_�*�_Dzoᱽ��ӥ|�K�JA�W�~�|��w��M	��`���Tῴ�s(��ح{M|��A�u~�+Tߺ�2����U������^��w����Q��\?�U��g����Q�C�T{η{�,�i$N��ν<|
��.��� ��Ցr�Kޓ�z�5�����օ�9�;U>%� 8��}qT���{+jw��Up̮�+�}�7r�{pe�]�=�����g��x`����wH�ht�Ӓ�������̙ӂ�D*]�nT/t����"���ԾЂҍ-qm���}|C��.p P���|�tۊ�ݧy�X81��Pp`wouJ'���!K�l�Z&h:�ܜ����g�Em�Ɖ��riI�@J��Qw疨�L��H��\Qn`]E������Ť�jr��hP�ټb�s��442Td�-��#"���Ӳ�oM�]��6���S�ۂ�ճj�(fy�^��ᐠ���o]���� c�+�Ԙ�V_�x�n�m*"U���9�o6��1�h��N�Y�Lx� ���7[[,�dM��$Au;Lm��r�[zd� ���e˽�U��')�x�U{�u���Fj��b�]���o���{̄���o����fԏv����m� �
�4����
��{e����݃�ʆu<�wJ(=+��	O�s��Q��^�w�+�׶mlf����b*:��ɡ���B�к�;��GmN�^���2f��SF&9Tb���Qa��\n9-FqSE�pnZ�P��E�D��Q��.f�o6�RvD���;� d�`J��{�L7��
F�I�:� r�E����.1��z�Z���
���;4��+��ݻC{��\���RE�P�ķ�c2�����R�;�$��Ɲ,|�`��}]/ �-�X���y;5z ��T0� �ᒢ�@e�J�(�픯.�72�zc���
I4z-I�h$R�l��Ь�4б45��t�+1�B�����#�~Y>3#ލ����7N9n>��&�2�CL���/�+��W݊�!����z���(㕬����ۺT��0�Eٜ�U�G��1�.�PY����٪.<��67�l��w5\n�'�QU���:��x�N���n��Y�V��k��ρ��12r(��8�X�9��������(�'�Y\���RX�&������w��PX�!3g�|�F)@�����.���]G-�f^�1��ڼf��V��Hy�m4�Ժp����o��5���3�@x��_�,J�[�[��	woK/= ��ͣ���}ZPY.���Mh��
_��5��.E�eh<��N�\<��n��ts%���|�n&��v2ȱÓ[e�Yw4��`�X��F�ܫ:o��5�E�t_B�B7o4�st7v#.�3-�K:�;N�g.�0Ћ4�66�i�d�厽7׼O��ؚ꣍�n�J�殼ʨ��aq<l]?�m�"�+�Z��;��i��L�������A\mn��I�;�S1ɐ�6�����d�F�޼������������8s_�ε�� ��r�0�鼟;�HU"����Uჩ�E�?4��=��ǆ��e\�-����5Մ��2�ֹt�Z8$�"i�f�7�>�_�|.��_#X���5s��X���9r6��[��\\X�n.�&ŮJ���9Q\\�.r�Ƹָ��ۃ���s�+�8�"ė9��r��U�rs�9����js�%�ě�.#��9ȭ�qō�q,nis��m�si�s��579�U̸
�9L4Q����U�\�.s��ؤ���Nr�`�9�ƐqȊō�q��s\͸ۊ8����2h�ح����q���5ɭƸ��Ӝ�\��@U|Չ��fA�;�C�D��@���Pͣ����[��A��C:�I��٢����[�����hTCq�#��Ի.�cZs�GF�9���B�e{���L��r�y�=>����Kex�\{.�y43��5���"<����ث��mz���גIڙc�&x;��|�:��s��V�x�mi~/ǲnx��6��/x_V�.Q9�;����Vf賈�e� �."�Rw^�8�Պ�޿<ӯ,:��{=ay^���{�<z��ǻ>.��=���C<IUX �H�>�ԪR'�ᚦ}�d3��+�Y]�u��=��~��/ �(ô=����/!�D�����u���;�5S��o}�潒s<=�^�:
�����s�s�;O���u�&�s%�" jy��NϢ��,�1Ը�M��Y��09����Q���.�x��`�kA�{נ_��Ɣ��wh��HB�k_��Mǅ�/&���/҅dT�:7#��|�G\6��_��>#��.uW[w�Q8��Ȩ[���}�z!M�!QsӦf��K��>+o˩�Dy�UI�q��Bbp�w�fŗ�u]eύe���5}fI�Y=_�}b}d/��VF.�aO5to�j�P�Ѿ�^c����9�'�*R�վ��� �;���wY�r�t&���Sǳ�4��gZs%�A���6:��A�2)z����{�/�..��77bG��I�X��"�n��}����R���f���u3�}Q�Jot�[����-*��M<9��Y�Fh^[0ֻ7쌏w��E��P�M���	돗�E��mH5��P�;p��/,ó႖a��O�����V��O�������6/U/F�%�7�o�x�Ƕ�z�s�갪�E��'h���xo�<�f�\%��~�]�߆x+^f���p�{=�@^�W���^�m��o�s��'k=��]SrmUR�>J���]�W����(���vWǧ!Ҵ�����f�7<!<�P��J~>'=S�.��A�ƎTy��Fc�ݣ�{מ�>�o&x/�6e��3�]O�迍:S��c��n����Y=/��S%�|)a�[W�G|����W�jڞ4<J]X�x�$����e��{��z㪘��^�w�O2����
�c�]������J�Ev��Q�N���TĒ�O|����Y�3U���)��B����z5z�~�	������[���9���3Ĕ8f/|���Ҧ=��1Py���o��ϼ[���ާ�Kw�+�yθ�P��yQo�~ρ�^�r���GM�k�� �kk�S��7��Wj�EוE/W�#��s������{=S���k�{��6�g�.�]D�sUf��l�	�w�Sk��!19�ޒ�l7ZMn�3�i��@h.���o	{@`/��^F���[{���FA���^�"�:fż�gK缪���UH�n��[��ϗ�`���\7����:u('׏"�����?��>5�t������p0���F�*Ac�[f<s���C��g}E�ى����'ɫ��w~4-̖iT��t��W�и�=��3���j�vߝ}�=�ƷՈ^Fz-<��=�;,�s�����W!)��;_D�~��B�O��ї�Y����n�8�^�V-S��e��~VG����Bn|O����|��O�rB�OP2>ʇ���c[3�3"�o=Q�������x�í�W��ܪM���ޯ��㽷 �)�*���;�빷z:�T�y]-����
�[��n_#��_��ˇ�߮���P�{n�+�=��{��cۑB�ƶ��s��=��9`�PrXWgC���ۥO����o:ݏ\��a�'<X��pэ7J|��nU�D��V#��o�p�?���L�~�:���J����u0*��#���IF�,���O�a^?����o����7w�*��Y;�ü�>E��:tӠ<���TJ� K�fgj�g65=�p��[߯���2�O��Ojڞ4<J@ò��T?�S^�^���,�^J9; 
���)ek�J�S5�������>��!Y�J�Mɶ�z�JꃪnmNr�����Dcjc�j*+���}��	�U��9�V�e�d��|�̄c	����n�W�(ш������aG�}�~�d��5b��z+#a��˥ %�d ��?C�~�������]���� ��F���$����N+��Skca�H^G���Y�C��5�Աƀ���#|����H���o���yׇ9�A��6X��?{���n�K�K����`G��ȩ���]K.�Э�n��";�<_�Ig�F��,to�VO�5�˧u�~�?{5���lp@�@�>nPȅ�O�>�_�
��z��� C���|����̟m���������:�\�(F�����.	^S��
�C��5���w�fw��^az��3ӽ~�Ը�����q�\U�%���<LOҽ]Dp��H�˄(g�_��d��iCޡ����w{�����'�ƣ�����"�~�(}�>�u��)���iU�oՊ[���n�h�Gj���LLoD&��_�(8� 7�M���e�Ύ�Bn����f��|T͏��<ld��u/�h��|R�TyC���E{ޠ;��]�\�����{61kϖ���B��&��x����X���ԭ:/m��V��/��O�|c����ԏ����;SoDH�,�EXM��Kko�҂"T�7���B��Iȷbv��rЁd�E,]۽����N��*���6#ow#��}��z�쮼�{W;�`��Gv���3�U�E��m��33��ުQpԛC�ρ�ݚ&���;(�Ԧ��}S��m��2:
8;a�����'�����f���U|2a����*}�E�u��oS������z���F��s�4{��k#_�o�?*�*�}z,\;�6k�FC��#�+^�S��^���j�z�+���g��y� U�w�.�zs���uc���m!q��#-O�ݿ�����O���a����m�w�����O"V� ��ՑJ�/zN���jr=�H,�{�G$�	s�)�N1q�:n����IQ~����Ciy&k���q�>�3������χ��x����2q�/�w'ى�]y�f��xV�'Tˏt<��)��t%��>�Xqޟ���1�1yb����
W�ojr�;;��=�kQ�ea�k���& "�ԪB��/.���P�YlW��3�18�ǲ�}Bǡ�:���P��~w�������3ĕPe�0
D�>�Ԍӽ�6�K�,�F�m���j�J�޵�Pr�X9{�̮�;~�
�:��|j9T�<ϓ�Ne)C=�6˖��O�����}��AW�����^gpw��&��yLe|�I�y#�v�����eZ6,�]��N�5�װέ�3��T�Ê�[ױַ�)��p�}]��|���I0�<nQv{�T�^��My�Nl�ig���6�����U���P5���˼�Q��g 벙u9V��5qɲ]� m7���]��1�L�;��e�X]��뙝��b�f��P>��P�s����M���>���Y���@�{��\ٷ�y�K�[ԏ��y̓�_B�-M��'���
���͎2�m�_w:����'�ͻY�����V��^-�}��&���"�˞�L/B�K��QAz^OWio�c�m��(W�זd��Y��F������O��(2{bL>�>�-m�ͷ^�V�3Ҧ��d+�S�k�<�V��w����G��}C�7��'�{4X��mH5>%T�}p't��gE905�>��wYc�z��g�s���9_���:�����!��x��G�͏{UE ����<N=��ÞE�Փ��oR�otv����V��S>�p�˥������%�{I��ü�~���_
��f(�9�W��BԶ�I�9`�ۉ���������Y�nxBy�랔�|NT�2��1�4ͩQ�s�[;��nz)z�|tU����:v�X�'�ʟQ�%��%����1C�᢮��ސ4[T���]�����]w�ϝ�����a}�jxݟ��c(���ϑ��t~m~:q
��ۜ��t2f=�g���]H�*֚V;ΓV�v���x%�t�꼿�:��u���{���.�G|�C��qp��u��km�W��!*��h�1���F�*�Y6��Q���W����U1έ�b������Rd���+].u�ko9��N����[�Zo1XԷ�#W�yZ^��xn{��V}^�<��F9��f�x~ ��-Y�چ��rxSحžu���K��:�X����G�x�z@{�~�=�>u���%��x��ڼ��3v�6n��&��?#��#>�v�O�.��^�y�f��|o<���z��ư��1��lP���Gy�{	~� c�������8e\-�w�q^�RE|�w�q�����5V��\s^��ޘ��U�46f)�Q z���P�EC�H,�z��K�(��#׬ym\�8�zgp�ޡ;䗊��� Ԙ�_F�$�9QB����B3���]<���ɽ�j���#���c>��Y��L�~c�n�P.N�L��;d/���#n6�C�+�ݭqU�9���T��vG�����Zn�O�z|�����AP��� �|F �SEN���J�oܒ�5S�}�G�q^T{O|���2�\�{��q�_�����q�ېw��wW�|��lyW��w�d߁6�?�����L��?ps��
5�^����Ͻ@z���¶.���y��C���������*2�F��a7/�g�����6��N���t�b\T�:g���;�X��E��֑��W�q��z��_j��s����bj��2���XӄB���N��Sg�|{e�y"�T���^�3zJ�X�A�Y�rT�J��c�U��X��~��8�7>�0�v�^���i:o�����=b\״�Ry�x���l��;>�	Ui�f��w��{��m��h����3���l�u�G"�M~D凫�͍�aG���<�����G��s�A���=�Q�{��F*�Ì�9�du��z(r�����^��HTЙ���Wy�7��,lO�z�
�������Hw�{i�V���R�3��ؿvz�����3��X�)��G{�ʯ��Tyƨx<����p�_�=�~�<��hx,u���YR;'���Q���it��<��p�O��A�P���\��>wp�z��|G��Ǻ��L�χz��a�e�[��s�Y������.���'�g�CS*e��ϖ]K7�X�����{�x�>��d�X<n+Y��s<[~6{���ݑk|}���8 r�,	��@��C]?����^�mz�&��P�5�o��c�3��N���	�$���#$�_( r������.	^S��n`�.+��'g�-|;����y��޿~��W�����~��	e�<LdE���Ƣ�5��2�B�y�ίk��Ʒ�a�G��D���Zx��վ~��g�������Q��GOeۚ�5֘1���%` �:&��wWR�Lu��H��x�M�i�Uݚ��N��EA��Aڕ�Xs]N7�
����K�R�����Vw�)W4�ʽ�H�����[��y��p��팃�R'�����7�z�_�%��a+�4Ӿ�]~��~�:}�� �ˣ#��~ݸ^)�1��j�&�~� }��������;�*��cՕ�����t�L�Pg�4��'ڲ��p=��M�(z�������M�������]�~yǍPۈr�dҘeH��G��I�82�ׅ{z���������@׷E����d{�{����ϠO{Քx{���y�Ɇ�gC�hvx�`F?],3��]~��$·{�_�suV4{���#5��z^��V%o��ujl��z3+�!�|"o�0dg��iznrwD���[��d�s���n��V��\�����w�����p���߲�>���+1��|�bv]���>��������S�J�� �5d\�R����1���xw=�"1E��-z�*1��.��I�r��P�;0����*�.��M��:�|]%>�;�#I܀�)�%��E�◽��5�â�I=S(z�L�w3�1}n����z�<�ޯ��o��h'��m'���v�o%#Ւ�QM��M.�e����0���c��)B��u]wn�7�[:za�Mv9^��ϳ���o��'�Ӻ�M ��=�@����	(���*KA����VY��KC0_V�Gy�4+�)G9�H.�	9������q�fq:̳ZH:̰&�,]J�.:�N}Kq�y �ʵ�f{�k��yӍ���<�2��<u��{C���Y�g�*�2��R$/���2g��ۋk}�ز}�'�ul(�]�Ȱ���^4p��pp��W�z�d�d@�B�r�P�דW��w���#��֓D���9��o����/3�;�cI�����z��f��k��Seڣ~�Y�98 '�\�W�����b(s43�Chwz���Ni��|�d]W��ϐ��G�k�\���l��Ъ���2J
��Sg���_�B�"��ѹ�_���*:�W�6�˒���������}���%�DNx��3X4�
���L/8
�{Ɔץi�]O��dWP�^I�zKݧ3|b�;ΪH���(�z|#}c����%3��;A���+"'��U}�jЙ�31�Ů^r½�'C�U�E��܋{��~>w����c�� �t��C&yܶ�C٪��]�����k1���zUq|���p�μ��}�C�P���c�����&9Ą�����7�Vd��j�jq4{h��Z�ùx�ok�
3ji۷�C��A��j��_%w����3ˤu�FW$3T�v��v��1G`i;Ev�!X v�dD�wbb�k3�����.����J85�e���D�˖�}V�d�tq�n�c��l��
Z�9ǯ��	j8���oN�����nm�8K�3����02�:i���d�'v�v6ۊ�ͭ��)_Ô�u�ڰ:-��uua&��b�s�������F��)'5�v�;�]w`u#���j�����`z�׷Y�6�)��O���	��.=�S.�}��`tI��80��jv�Z���˲e��+��](�wEI xEͫZ�n��U�_Cm���B�ց`M��QU^�|^Zڎ��:�2��u=�$���8f�Xe0H͛�7k,>��N���ӧ4#Pep���‧yJ��v�_G�(<<�`n+��#C�Ju����XpHe�2f1��b���F�6��"z��j`W�/.�A= wZ��A>��oɁ{B��L��#o�e�S.Y�$V��P�a���\	��ugX�]u�`v�V\�mwVi�n�X�-�Iܱ��˹���V xskr R�cm�n
cXΣ�\��f�y�M�܃Ô�'�h`��1Yb�ܣ"�h�m��3|�4f��NTf1u�{e����"&����SOj��`]p�o��p��b��mՑ��oIä8��r��w*�FQ��G��Y�3"f��8����m�ȴ��4Y�v���-=WEˡ��PJC���X�{S���h�	�Q��[�E�n�	6)���f�s�h�F�\�9����D��ƎL�W�qR�i�n����8��uc��M�n[�ë=݈��b�� �p�w���x����V�pP vt�|�kc�vF�����vu��G2�W�M�G l��f@�\��r�e���w{���uΛـe�˦ur�����Gx�U�S����цjW��WC"C�3BX���Yu��܆�j)^A���e�J�=�Y&`i���m�2����.q���@��v}���T�ռZ^�D���7/�'�^7tn+ݩ�5$�`�)�>{M�����̔�n�"ks�W3
 땴����@`���hnu)�
���pro/ʖ��r�(�
ze�U�NrV���T��P�#Hyu���-c�q��7k���WGY�^	�ٛv(ƶ�7��{�)�ۥhb���D��AjT��e�PWb���z��D��ʓ��.i�1��|�<&��:��/�Ճ�4�;�rwl<xb��)Uٗx2�A�bj�����}�U�lQ9�_Q��\�Xo���w��	����v��ñU��{��eu��8;��H*�L`v]j�5�D��	&�]T�^�HV�lK���NǼ�Ѳ��Q<��0`�|�o�t0�Nm�O���W�����[�ց�Gq�E#J���鸵0�z�dw
L�rR���ٴj''Ǿ��X�����5qFs�c�6�qs��\\lW��I����NsW%n4h������\k���c�q�)�\[��),pU�r��6�s��I\�
����1I���ss��"�&ɍ+��Q��n8� �T�95s��%�Ѹ�\AƸ���	�9ȩ�W3\Tq��Mq�&��-��9�.s��k�n+�(�1b�D��W�؈s�W��Zqs!BS��Q� �b.4q��E��Z)5P%	qŊ\\����F �.7(#U�]�_�wU@C2'u���!y�6�kqW8r��z�V�;��I���
;�0�=��@��Wx�9��V�a)Jof��O�l�.���\�zx�a[�@�=_+\̓�M���x^�W�����'^�;�u�<,Ϛ;��Rj��o��g�y\䜾��o��!�+*��+ģ�v\�UQ.ix��hcL gZ�+��G:�]����K>N��y3�x�9�,e@�஧�tY�C�t��˭�#�4�6'ΉK/\細UO#�����~�f.5mO��R�2�@<X�|�n
�p��7|]������W�<f�x5߁������?>�=��q��T��I;�Gx�O�!8}�iy{z�j�!�L��wHS�x��8�z�{A�9�@{��c�q�R�e{��L b�7��گ:���K��E���C��^��O��}qW��~ӟ/H��HJ��*#w�E�,uu[>��c��E_�w��{����:u�H�zh4TC�+��W�#�g|W�~�u�k��;.�cC۷ㇽ	����:�e�;
�dCs���P̈FZ/���Wf��wrFſe�v����c1�N�����{I��Q9޻��K4�Hj�DL��4.����;�_�{�z�azV���;b�7��d\O~��:��v�kbbs�&^�����,�y��N	�ۓ1��v^��8N��HU�X,)������퉃K��vb�D`�m�*�b�Ug}%��n�X�^p䶀��,�k��;������K�)M�,����{���r:�W��G��ύ�g<O_�(`�]"l3='A!�"v���в��7�.Qj�m�j�#1�r�'���dx[�p�����ϙ��+��	���S���t{�yiNz�u�x�����%��6�㊅��M�+�`w�T�}@z�����q�347�>���Qb�Mr=�˳�
(��a�������ݹ||���_꺇���C�P����àd]������>�]��,\2�g8�zO���·9>�R�����~7�u��\�L��u����}�R����N���w߿Vq�fp�>;:O��Áɹ8:*�N�Y���P���\��N��iP���~�3\s~�U�7�YU��AN홇�|���y�62N���*3o���Y�t��H��#������.���y8�>�K�1�4��j�]n>�EVy��d����
�CԼ�� y��U�7޲.J�����1��<9|�-��}A����B�M�Z��W^��l���_�UA�=E��[�w w��w�x����KB�@;�M�݁��NP.�{�.e
����T��Tbu.d+g�����w����D>b#~���'-X�U�UmB�����̾1�B_0����qx�[��YL�S�k7���1���cH���Z �����Ӻ�!�K�����m�L;*n��q�5lY�9�Xs��{V��T�YY��+�z�]C����`L*�u3�"��R�MT*����&�C�5U�#�vedz�ly��	7g��Y�z�x�x�@64��ʌ�&�|��2]?�<���n���mmrᛕ�ٞb��|6,|���g��;^�P��UW�"��L9Q�=��1�er�4[`^�ּ����f|=q�����Θ�ͦ7�Ը��������AW�d�L��w�oR���s͊��u���H<���Gx�q#���#�~t�>�"}�x�~���������y�O#ٷF��ïv���L���Ϥ���W��|r���x����j�%�ҁ��DFxF�i~������	b�z�'�#�:z�S�h�.�a�a�k��5���>��և�4�����d�e@�7���9���w�����7����l�FS�%�����Zt^����|k���gު�uUp�c������uV���>��<�޽�|}�p��|J�0������Njުn�a���暴��md���{�_nUXc�זF}��;ӑ�׎�XUs$&8��+�wկm:�l���!��eZ���C��kC2����o�($���:��n�k�Z�+/���Rr��G�}�WU�M�Ⱦ��Ɍ_w`���B����*#��v��N���]�ΕԨ��7{dv���8)w����ܒC�r�ʤP�������Օ�7*��]~ ^�ׁs��}�o��ң4��؜W�V�.�״ץ�r���g/��o�4����t����Tl�F&���^��I߽u�����~%E�j�Ǌbݛ[���%;%_�>%'���B�L�<#�X;>�=>'{���Pw���R�3ugA�W���z��}��3����$�|��N�_�/ܪ}��'7���I�`Cٗ9���d�'���@�ޠ������P��9�F�Xe���Q���X��T�nq�}��t�:�K�:�>�b�>w��<�����~u�]g�z,�u�$�X�d�o�X����o�ɏS�9���ױB������2�ʎ���RM�_�=�$���6jqcсv�Vo�����f.��L������C����AP��Ӌ����Hq7��Hݻ�-nxq���]��	�K�B � *#��`�>�&8��k��m����>����aJ�r�⣞��9~��Oos�>�L�5�s$�J��6zH/҅g�/���_���Tq��]��n���v�9 ��=�a;�	^n��7���޸o��)���a=�b\���iS�X��և!7k�%}�v�J��76U�]�QV:�c�<.f�:^$��f��wɰ�n=�\�DN�
���y�:�����y��K���Sp�g�e��)e�O�ޟ2Y�>��>ϙ��d�E�N�fC�\)���/
��^�{�IPv�v�ڽ��N�|;��{ΪH}�Ez|#}|P���d��:,��}Dv��w���;>�A{k'�<��kz|5CWxϓ�܋����~�=p��B�֦
�'��w�<�i�JJeN��ѽ�9�:�[����弯Æu]xsi{M��G��J�,�{%G��}3ހ�Y^�'.�N,��ߤ_' X�Fd���2��9���g[��U�'��i�mn�"C��^�ω��sY<%��쾋�\���Û�xd�t;�����Qώˁ_-��i�o��י�"��syy�ǉ�z�|W��;���7��gE�IӤ��3��)�9�\��W�ێ�FW;CȊ;:�ؐ�X�y���^�W�^,�>.�\�n��q�x�J�ޙ���<X�o���z��ЧEh�̞k=,�R^�4���/�q�csާ���!�kQ��e��<I��&�f5*VhM�}z�q8A�C�3�n:�Cǖ!���F{���s����c�\ܠ����z�U�ٺA���J����)�:7ɴlQJqr����m<XE�Y����q&�]���'#Y6��JnWQ ���s��*7��ջ�:v]���AME��Isb�RpeoWWe�"�V=�S��g��յ�xa�\H�c^溋�olRYO[^<|4�'��G�|��g��I	��؂��a~1�~�!���t�'-n�0d{XY�)�#��߂ρ�}Q@���n�P)��Ts7��AW�^����rxu�;h�'�U��h�?IҮ��m��f� ����*�����9 �3>FZ-unZ��A�<�Ӿݝ���k�/}���c>��_��>��k��	���:d�MI�cdŉ/�hi޹8��{R�6s���Z�C�ף��>t|lzg<OX�C!��Jf\��0���q�&a�M�dyзY��z�Ǣs+h��j�Si�
�܋��x�d|=>}��`�P2{�Q'��%�H�J��u~dׄ��Gւ�f��ڼۇ���߃󚒾{��q�_���%������Ly.���o�ېi�%@��������n���||��)|n3�.~Kb=�^b���L=�|��DZ>�ޥ�]��e�G�3���Q��O�����O�o��i:lf�x��P��X}Y��K���������������Wq=�^�fl�?�,�~���,�ճ�f�g��r�w��47*�b z8�����*��<G{�e��Sꩻ�8\:��%��X�����:4Ԋ'y�I��݁�޺���={��=�Dxy�7�vv�na��4`}�������9t���|��W|�<���['V��ƶt#6�'��}Xw{9d��P���{���1N\��`^�q�%��@s6��7V;�9�#�U��A�'2���W�*6�8�@R�G�k��CՓZD�,�K]�E�J��x�]?��C��Ԇ���=0�ĒT�F^\��������#�W��Ciy&z� 6�uP�y}�"�J���/�ǟ�������Q��&�¼�R8|������I:W�{�-����G�O�H>�7��lg�<}�O<ǨWC0������v_�gO������%Ӟ���`L4:��t�IK-9P��z��'n&�_��;>>�{�G�ޘ��7��k�c��c�[��li��`O�J��ϸ�\��:-g޼�B�ٗ/q�Y����s�Z3����ߣ�N�����v��v�<'��h��s���D�x��e��YRG��S�}�A�W���zw��{ӸK�z��Uz��2x���J:7^YVW��;��"s�D�"D�MG�}�P���p���;c �ԉ����}�N��ܡ�^�=�W��xO�L��f1�����7E�ھ��p�i���~� A?~&�۠���LAXJ�XU��t̂�������-�WH\����i���Q�ۮ���ܠ�s[���k��U�C*]�PN8`̾{p+c������\���]��,���fhN�w$����ÈN��g8/w������*ӽ��l�9����"׉y�Y�������`�)�3���񿊛�����AOx�4�i���P�o�+�>������{[��h�>��P�f�gd�F�Q��c�zpzJӃ~�}~�豷t�08�.�,&�9�_?U���{�ZFw��O{'�'k�=��;�4pi�,Y���]I��~��.�ϣ��$������F�x;�ۼϺ�}��s�~�/����g��@��6g�/g����bk0����{���'4��������qu�E��>���w������v6�=v#���j@�ߣ}7��,��F�_hz����*{Ļ��!|��K�~���!��^���D{E��~X�_������_���z��ᄻ/�3�
��3_mO����<�L�����A�o]]ϗ8��^�Z���^�b�T�}$���=Qg��|�7�З>��y�7ݙGgr�g�o�w�w���r<^�K�S�Q�P�ea�n/���e� �/j��礑�F���/���1�]ӧ9X�ޯ�z���}CǮ�ǻ>.��=�$�L�%�E���>�� �;�#jb�������t���]Vb~�{.�p���OF�ړ�7V����l@�R�7�վD_5r��*�mɖ%0�'b>�(gAʡ<���;}�ʹ9V��D	l0��H�He�j:zo5:�ޜ�M�M��Áw֍�u�N7s�F�L�ɛ�����f^jqe�O���B�?^���2�<���'�z��X��st�mg�9�G<ۯ>���2�/���]heg��Ǘ����qy���q��^�$���W�y���W~q�%J �I Ǜ��|}�L4q����7Rw:���R��>��u]�����XG��Ư�2K
Ijt��2�HUԾ:78��~����n�z���^Gy�ۓp�>D�����C5�3L���\�a{B����׶�ק$���VxZ�{�¼<�����]ɋ�߬Ѹ~�@�11��?!�o6�ezcK�4v<tx�7V�珴I�&r�H�ؗk�oA�������'���=So��'�{"�G{*AWq��<��@�����M<�{�=į����}^�Ҩ���z�4<���ng�S�P�l��l��ΣԱ���1/a��l�{#έL]�'�q�9�u �y�S=���{Ưk��O%�%_D�2���ưY��GK��͟{�Q=q�s���rNq�8o =f<r:ե����Y�O߾ʊ�(Т�4}Jɯ�~
~��߳c�Ys^�p���B���(VP˵�����,HWVt���q���x�n�mNu�^�}R�����ީ�ұD����.��ޤ�%ԥ[X]>o��w]��aWu�f�Q��I�r�F�Q���gV�|�=PA��[�1�������~�?M1�v=s�+��Yרޛɝ�t�,^@���N�0�c�2/�Edy��y��s�L��w�*L�r�&V}���[�c��:(����US��\l_���8nf�v׮Z�3C�S+��Pe��f��o����=LnG�O�ez��Ϝ�dP�jxϪ��B=�g�o7=^�M������Je�Cj��u�����}�pǸO�w>�P��������I�f�d���;y�^�~�*O4�'�2<"~>ht��lu���t���u�<�jvy{���t�s#-gG_��E��~�6�z����� r�����7P ${{�a��ʢ�]��`)UL�sj�5��O}���8;��W�����ճL�Y�PGS z�~(f?i��N_����;>�����{ʜ;���E��ͯq���'��~Ix��d����t���k޹����W'�/ ת�hz�R;����9�^x��Ͻ3�%�Ld�n�ic���.Lx��f�ߵx"8Ki�1��`z�'��p�N��䩒�9`m�����D}G�}�>�V���ŭV�����Z�ۚ�k[o�V����k[o��U�m�εZ�����k[o�kU�m��V����k[o��k[nkU�m���k[o�֫Z��j����kU�m�ƵZ����U�m�٭V����V�����
�2���Lu@"r�������>������� ��(P �@( �(
E (��P(U@��$�
*R%$AI*AT "EJ���
R*��)U$�U	@P
Q$�*%��& �Z!f0ղ�X%bB���(��;��� �S��J��G �  	�  �mc%�*�J�R�B\ p�"��T���
�ZCLl��l2	� gH�eB�V�ɠ�2�jZ�t�͹'gwq��m
��EBT�� Ym�Qu�3�&�ԕnn�Wwwr��lt�7�s���WmV�7p(��)$�`gv�9��ۧB�����5��ݻYm�)mZkMf�Wu�t��4�**� `m��+���i'vnn��G.��fԢ�lJ#6�T����P(�.��6��Ba�3
��B�R�354(�U(W ;BS���lJȰbl�lcM��S��p�Q[5���iU	h�ͶKf)[1*�l���    Q�f
�RH�      ��0�)%2i�4 ѦM@2�#j2d      ���R�OS@ �L    �$A4	�0�Q�ij1�&� ��JR� '��! 0 0�̆Q�(�c�#c	&HZNP�� �� ԡY̒A���Y	$H�@��r0���R�"b�Xtb�J~R�'�g����
���QQ#	J�(hF���D�Q���*�Dʑ�їl��Oחo/?/��H"iғ^��K�{���`�Ek�^ugs�U*s�i�X��IT�����W�+���'3�����g.�g-�T��y62�֌Y[J�A{�:�n�)�CgE�ɛF�Ur� �Ѓ	{u��34����(=NՋ�IY�VQ���⡂�Yl ��v
vL���i������X�Ѵnܰt�ws2=��ncT���f�%�U�� ź%3)�w��a�A��,��Jk��:��e#�B�?Y�����(o&��=Vt�]�-U��Hd��BnR�ʹ[�:���y-�Zv�A/t�ub��V��G����:�M[Y[�l�g�
�.���Ku�ޜt�m�7�f�W��^�J�ή�m����s�f$�6��l��D
cO^��$�`/,E�h9V�7�<�t�\�m�vx<���5�#��nҷ
�,m�)��RIq���Y%9��l�V�jр��<�1��m���00���n�bJV;����#�Ue�a-6l��kī���mԦ�f�,d�6��-iZ�PI�)e]�R�t�1 �m<;*%� ֭ԏσǹ���"̷���Q��=B����}ǝe������%��X��C)�Q��m���MkiKh�e֬�o-��
���y�ZR�&ҕvmfD�v@[D�c���i�����.��U�v�-,B�vӥg���'P�V.�<����Ƙ�v��կ���۱�X4����R��۸��`&��@�����M�q���v<B+���ҬCŤmʺ�E�[�z�%h�h��m��-��7����8X@��!��ތQ&��̬�b5��T"�2�k�)���-ū*��Œ�-gB���ۿ�]�-�5���Bن�{-Y��ޠ���[��@��ܵ�;�i�Y&�N��l:S��Ue��,ohB�n�0�1e\t�iˈ��a�Q�U��{���H��׋5P[8f��XLz�s\E�gd�V��A��t��}�n���oh�+wk6���ni�YSF��j6�7�@<x�*�10sY�{f��8�m�;��$��pi+\;{���4e���S:9�H���I�����<1<�׬��+�����YwI[�k*��4�V��&��PSz�f`�%��hXu��P]J�[+si��k�(���b�6 /)��*[v����7�Y�V����VV�n��pkt�H5�[�ܳ�H���ɨ�ֲ]�Td�9;݂�T�u6Ei�6�+�^�~i���i�	�Yv�{f���&<�.��lq�,ec���ocý�ss�Ƅ��e��]]3��N���aO�R��k4��"=�c�XU�ɶX�n�z遺��f̥�V%�h���Ͳ�>F� \�X��h�΍t���6$�"�������Xղ�f�YYN�ӼU���@k�@]̗�eAۢ�ЈL�P��d�&Ι��v��M@���wS@��B�V��Mm��;W�<������&��"�5t3d�+�3� �qܫvԺ���A�z2^�&�y�h%�bųa�Iaol@$"�	�V.BkK�o	����V�<�m���\���1//*Z�iؤ��)[���l�1�l��ͬ(lی��� �S�wm��L��׶����]L�(����;1�x���U�[X���w`d �z��E��9��x�D�mJ:ν��81�@��X@�4a�{�R�b[۩��Jdp.e�4�6�dl���E�Q]��,��oXo���W�WW�a�Ckh\mqd^��ɳ�f�5�h�Ԃac�Y�k]=��+h�	#s_̽�4\(<I���B��U�+z(�Cm�J�Zg�e�#o�x@��U���5VD�֩e���sn&��
`�f��701/T�9���J�Roj����뗚�P�Z�E�z���7U�
f#�~���<��o+� {�J�����[<錣�El�z�/�#N<��u\�kQZ�%���{J��n��qV�"�2�~�#�����v(>YkK�Dn�8�내a�v����q����
�j�k�"���PM��8<Vn���d��к�6qrY�n�p�y�z��N��/��n�ˆ��YR7RW"ٗm��՚�@��K����������p�X���h�h�Tb�o6�ƭ�ͰbEZ3f��[�ݎ�^lג򐨤nXFC�YZS�T՝t��m��[/3/�TX���w��,
C.ek��Y1�
�z@ٷw��k�&�\F�WYrv���$e%��r;�4n����k���ϱ��wa=yp�)B&a��c@P�-m��]�d��6��6�)����7F��\�����v���5�Ң �w8�Gv������"�h��u�2��(`�.�مD�(�����1���pU�S�
i��WP�Wa�+{x��Ǐi��eh�s&��hIdM<������(h	�a3�aЗ�լ���Owr1����4+2��۽�3˶&h���JyxaЌ'�wS�i�?1�D���ʘ�E��\�j�ݕ��є�iM��f��l��"�	��a�x�Z�����P�.9�(\�sI�ە)���v�����MY�N��/�u�cv���U+�o\g!4Ľ ��1Y`�'�wa�F�N΁seKoE����ۣ�Gl�Z%c�����{�o(��t��B�T�
J�EE�9�[�{�[I��ky�\(�/�.��=�7A�h��zLW6���8Nk4r���b�[H�B�u}�[���aB�M_=��i]5d;t�;�Zَ�hj���i
(CuBLz�:��X��E�In�����ai�R݃r�ܭz�@��FV9XѲ&��I��<1��e�}�m��[m���n���m����Nc�("���ߞ-�4�C��(��u�E�YdF��mA����eք��
�~���i�(6֏����{�V���䧶Z�Cy6���f(�Ս6��t��	"��(��Ԗ��eXW7j#�J���5�&ν91�ug�ȍ����3R#���9���C}��o�s��k�o��?�?��ضS�"�����䦠��?������?�������R�����=�+�T��q��k{A�s� �C��"�����)�tXR�z�/�%ǣ��^��q>���P/Y���3締�)H�x��t���x�f�eo`P����]�Fq�T��%�F!�cOc�m�A�-��[�_\R����8*2qC��X�����R�@�{P.�����H�^h��:������tnȹ7t�v�����	�x�
�,���@R��c�he���r�!�.V37vcb;+gU�u�"*����n�݁�.�4sF�o����*�a�U�@C��n�h���nV�I�C�EXp���G�Ϻg^ ��Sz�kz�w[�(�:>��C8r?'�q�LCa+�K�+2:fr�Z4nݱ4����DU�ql�������q<��U ҧMd�Ĩ�Y�,�m�+�f7i��:r�0�t��{�ړ�͹�F5Ii���D�j��;7�0�-�����aףVu���K�����C)�!�y�;NiJ^h3,bvN��I��Y�����v�����/[�c�69s��Ą��#�V��Y�v\���^g�܎ޕV_��� ۙ�3ϯxi{77�IA�]p���#���g3�XQ(g[{G������3��U ��i�Y��6�8��n���p칸��/�z�FyK�-d��{o;���	�l`��_t7kB�H����2ں�R����pŇv�)��a�2���z�7YA�l�ldD饉��:��n�)���Ɗ�mҧ�=���A�V�zr��e_TK�e����,��+�%�7�C�\��@HV+��Wm�۝�y� &[�wg;���</OEB�ޚr�{��	b���)+�R�ô.B�0�D��u7#�m��;�Y��j�AQ�V�$u����F2,�I���v�V͡nZR�4>��	�N��w��ld��U��������4�u)WB��'GW�Ir|:ƘҔr��xi�S@g��At�ϧC��Y������-9[u�ZH�kq�iU�fMyR��ђ��{��E_��e�����l�R����\�nS�����fL-��+*+�R���[V�W[�sB�r�f`O���э&�����Ec��c��R�t�[�o'��X�4���nt�W�)Iir�UA^�6v;��eMV+b�X��m(u�&G�[�}Π�,�xD=:�e�ƄRl� t{�勻`�b�� ��]�n��ں�R�k��.��{��;�7Q�%vJ��u���ዢÕ:V�ۇ�fᐛ�GO1�p����]��q!Zz����CM�ݻrO�2e-�Le
*������.��Q����b���/���oy�S��@�yM{R[}����ćj�(�X3R U�(�W]��:���W�/�BEX\HU��V(p�@'}1�cof�o�27��M�g��0����W]@��HB�gK9[�Q}Q)�N���e��u���>%m��v8�^]ǳ䵺jh��TwD�y���n�����]1"d��],*��՜Do��VD&i�����umv����G}˪̂�n2ܕ�4FNfZ�K-Y��형�q�,�i+n�.��ܩ����k�ph�������,�o�/lR�a={��>;/g9��S�0{��RN<��P�1c��|9��c2`j��;i]Ie;ְ�r��n&����k�
�{pE#S[���|��9��c�
ūv��Ô�Y%G%�4��I�� ��*���>�������׊�.V��gs)�4R=u����n^w7����X�0u��J�z"NŵQZ6�mJ��9Ckl���)�F:��n�`G��Y.����Q�\ݗnU���N�J@�]����.oVn�)�^��a���NZ+ml��!On��͙����,�K�8�N�r=�j$V��I�C�Ù�K���!�Ԍ@^��_P�l�CV웏nh��YqZt�#J�Y��:p����ҧ���R}��+z��V7,�\{����Y&�;+q)u=��- �;��61�G.U�se�8K���W! �=����t�����.�#�
N��r�V�<�	��v ��f�ʲBĘ�*=A���/��{��]'���/~�ɘ��-Z5;�����[�T��$�N�BK;��N�v�*�,�=C2޽��R.�����ڝ�����ڎ��｢��fzmf*�KW�nÔJ���}Q�� �c��j�$z�YM��ۡ(r��͕�M��r����*N���9]�3�!�8��t����׏y����Q���֚t%�y%��n��#��V#e=�#�����+$����K]HUX�s.�v���ˆ��;:Ӭ��S悉�ҡ���.	��o���_�m�W]M��FE�v��K�0�	oX܂�qp���J����8vr��"&�qs��u�IZf :[�c��ͼ�SB��ͨ�4�O��vҤI�w2Lnk���aɒ)'��$�I$�I$�I$�I$�I$�I$�;r]oN:�1j:kWf�Ǚ�J�e���k]`��Gj7��nVF��&U�+l�@{�i�E1�,e��Eٶ�fup�ѽU�yC���R�u,��5q�����p S�hqlt�N���k�2�n�Z�]*�8��J��r�H�Y�::\-n�%�m�u��C��G����:d�&V:Mj�=z��*���R�M;����ɲ�B�f�]�2LvmJ&-Ǫ��F�MD�y�Nǹ���(.N�_X�6 rA\�Y��l]��l�9Yh]��N;�0�M>2Z*�	�h�ٴ�_)�N��˻|$`۫I��`��{�
�]Xf��e�c�s;����4��j㭱f);Uo���A�R���&����g:�w��ԗ��s,d��R�t�Z1<W1�y�oK��$,�D)�H��:�tK�:IٝR�;���J��+��)A�W�{OU-�nJ[4�" Υ�hh��+hoTp9�q�X�AtX�2B�i"tؖ��*���ů�ΪK@��P*� �A�"���c"n�K��֍zlR�;ф$�'�੣~z�گ�F{��V��b�V�H�h��v��պ�.Ym'��n�a�D�PJ����odNl����Tx7R�8��11�
�[��+zNG��eY�a��Y;��X�m�ÆӤI�N��`1^�H�1��A�ʭ7�	�t�i�CxĨ>�s�=Ֆ�W	�t�]��P�6'P��@V��c(�kE�J^�@ʷ(傕�IU�,���)�Z��9�������
���R�"K6��b��(����|���qV��S
��Xkfd�V����n!�	�\�r|�֞]�/����eM��xe�;ie-����򶑘��5Wc��EN�V����{���(Q��o�|r!N�xu[4�;���,^Ywf��F%��\���F�v�)����5�H1Xj.S�����	�0�����p�T�q8�b�(��e��U�آ�^����НE�#F���ZVVn���������pL*�	iL�%ol�q�[K6ȡ�p����бM�̊TAٗ�j$�*���hz��L�s�0��ẩ �|��
�vk�5�b��N5v�
f��ެv��k,a��x��Wv\N������%��8��oT�C��o������=�Ki�yj�]}��k`��3X���f����
��ᯨ�a�6h���Γo�ķVj�^>�lV�%Rp�.�`
�]�z0:M�ƅ��5��e��\�h=T�.of�c6��Au73���h��I�*������|��4�T)CS�go�۱�&��� �7ճ��砭��n�;n� ��	%Fjj:�	�
�`�h�J���.[��Mg.��%�k�Ӧ��H�e�I@}�����}�+��J��n���7�B��}�Y5�D��|+�x�M��dZ��1�*�b���b����ev��L�7����;lVo-*|;I����]2G-��|Gۛuw��B�1�M�K�7�@p��3+>j�*p�dR�QE�\�]�"z�r����2Iw�w%��g���R����%1St��Z+��B���Ik����0�t�i���s+��h<�����\��Äk��� JWS�f��H͒TF��0S8�p,�y�2Ýiq�&�Vp\1.���-���]	F;� ���d=#��;t�f��o_\�:�=�87'�]����u�<�냨�|9��0�W�o�� �(;�N�Ʋe.&��]"x���X&d��eh4Ws��q�+s`���:=�t�n1��5X�E+V������hλ�D��na������ur&u�%XE�Gl%X�q<q�gz�#�=��fR�ע,ƙ�g�d�P�5��;Ŗ�]�q�م���������:g��cj���H�`W}m�E�/I���c��Sm�<�)8*o^Ju���*,DNR�S�#b�\�]Y��3��ʷC�勰N���̽VE�:<"��]-��	�B�w����I�dawneJד�Yvu���L�;�r���f��ZOAZ��T:uk�h��J��h`�ʏ�x W���)qӏ���'$$���#�^��a]�\�*m�O(��Yi��l�d�F�wN��]ܒ㸄�VRĔ��ޠ°-1�,�2��u��;f%gV�(Z�nm	�f��#ߔЪu��g�<���KdVfs�RW,����(�B*pcM,Åʓl�E7�a]p��5�*U�&4��trU�)o���V��X�]-52�J�R���+�M"�,<l^G�ҟ(��H��qL;�:s.X�T�e���K"�fǽ*`i`���٫/-r�O����.e��HVR�#�9�/�N�(j�vXWп�]\�J-�5��Y2��F��&ᒙY��p�#��Yg`Ue��,(�B�O4#���ԬCk��b��$�E�[�W�6N���+�:�T��B��x�����M����5�U�s��T�UwZ ���F��PEls����t�m�d��Q5Id嘕j��IЭ��K��V��a�b�tþ\�B�d�G�bu+zֈF�[��蚮����V����g��WS.��ũ�u{u���S�Z��j�:��t� *މ�Mr�H�6o�f���*�:v�w�JX8�n���+��(;b�W;eM�/��I���������^�mr!;J^q���H��Q��ҋv0@Q�`����V�z溂�y&gI��V:f�Z9ϝ����h��^�(��\���@W����ǆ��� t��E)���8���yL�'W>�ˋ:��z��4� 9��@ۧ	�	����Yr>�Pժ��ܟ)�9�ΛԞ�tQ�l�jNeȬ@3V]�d8�QY�{UƊ�a���ulW�N�d���.�M��R�dѹ�j[�tѷ��孰i��5�Um8m)F�Ǧ�ݸ�sn�P,��b��)
��ǥ'I���8�e4^�"�N�ۍ�V����\#�k$�v�n�)�^�y��Ǝ,.����*�|�b��G.�����Mug�[&���tv;��A6bB
��kgS�V��T��It�}�7��-x�Qb��h�M�;�ڳ)<�\Z���	��YzV3�0�!]2slPɓ8R8jL6�6s����f��<�a!����}�V��8vjn�ѺI%Yn4�X�.��TJ��딛�& ��ݞuv�f��Oa۹ka+�P��lK��j���6��Y��M�P����T+��S.�ԫ���e���A]��j�a3q$�+:@��&�l�i{J��\�I�
r'j�����.4{P>�GN�e*k3Dy�a�&�{���K5�:�6�T
��\/�+w)�^�$p�NnD���=7�k����˦{���e���V�j9%88L��U	���t�<E��(h���R����n�#q��t@=����j��uB��wdX�o-��@�:j�����8�5Z���H�=����}j��o�x{����B ���@�C���d�?J2_��?}vr��~z=�.�����8��tb�o@��)�M�����ז{)�Y�2���-oU3t�p��)֭��zAci��>���0�
�%OI���w��S����j�s�=���S���r�[���ZeBM�	ҦM�)�.��Jv�|�"����t��Ƴ/uhP�wt���m���s�����7(!хE|�5א�D���)9��2�k��%��V �qw��qg<ɉ��	�c��{0+#Q��nb���8��8f_P�9�j�J���+��z��v�E�lZ����^�zÜ��5ޥ~˕2�֪.8�%m���\�b%���e��ĸ�r�ZP�q�����z_1�D���-��/���X�)AlAZ�9Qs��-�FU�iV�C1kH���ژ�,��L28�ۂ��r�(ц8���f-�&V��&�*�3#Kl̢�<�Tng���B��g���[m�ܢ�D�[�┴Q�<�L��1��*)�\���3ƴ�Z��k��מk�h�{�o��|���C�����3���b�.��$U�I���:q��~���r��g ���2��tg&6o���!۫���r��^g*�F�z/g/R��3�n ^ѩ�+F3�i'w��SkT�.]ⲎQ�=��}4���כ���V������IL���:+��gD�Z���$���vz�4P�U���^X�?r�]��ǳ�2�{�#\M�7]��?�N�.'}n�o�~��;�3ߖ~�a�SiV��"�g�e٘�<�^�w�q��fˑVIbs7[�iIv,�[�f"��[�<�x��[0�#�w���~��
�޽�Hv%�T[�z�#j���}Kw�	t�ٞ�b�g��9h���	=���J'5h�!���y�����J��g�v���y����k��S��������XTWU*�ʄ����b��Fg�:o�+LѴ�lG�L+��o�٥�F��|���}�ћ�����[ט.c�^�������[
n�jS}��P���C�d�d7}1a���t��J֣pc��lc��M�k~]~\�Y��œ�@�W�0;
F1�/��f��;H=�um��A�o#Ub���b;���[,�u�3�a2�Gܧ3��Ѽ�e�I�-9���֡�ᇾ6E#\�#���jٙ��R�'�b#�T���
/}�+��vZ���`@�q��3���P��
������ܧ�Q�f�}�PC�U��
��`Y��+��t��$����ķ��r���'c8�p'�E�Wʈ��b�;��8m��`+ԭX��bQ�ԁ�m]?z>�o�*��פg8�K��ә���_g95x���S��B� �/�`4�)���X�6��!p����rg�8:��[�w�;��w\����)Q�+_	�ҙG�/�]���s���N܀W_C�ߝ���L�^x����(��b]{�'�б�Y�kH�u�$8^l�x��=�cS��܇[6�ԥ�������น��jGqD��b�N�{�bDVY�Wl�]<�b���hwx���e��z2��kXt(���-_��ov��b(��.�L���y&�����<&�D�ʉ���uz`5����y�����N��aS����a�y�N4�5i�un]��q������es�ylh�iț���MP`�%"_���H��V�:��u��(ƽ�B�ڮ0�,���Yf������
��Y����V�p�g$]�7�ۧ
m���v�NoG��z���Ѥ��8��z��ԃδ=��[�=c��^YM�H�tx璮�UY.��i��8e�෽��j�[{s�f��sa���q��6K�}�+��ON�#�䇰O�3��]�:8�X����G��4�����j��d��L��b��+;�퉴l<�HgKc*H�'�'��,�N��{���Fp��u��+��3P	�;\0D����ھ3b���n���Ak	3�i�FCYI��rO>�.���|d6��y�P��'���ד�T�ty���M�tc%$W�u��0 �����]lY�:��2�櫴�:zF�y5�}6��)u>�"���5G���#ޢ���3�Ig^�_�ý^u���Y��S�ddQ���RF����r��[�=ia�����u���=�ǘ+%���%N����R�{A^p��;��N�f��B�J�p�^
8�_I��G�*��;$���E�����ٝJN����Q#�I���6��b� Qi"�������ۈ'~���t��	����{Z�7��C���2/�u5FqQ���R���D|��36'�XnH����%� ��V>^�.�/)��\EMR��m@ZX�ؕ0j$${4��c�5��f�����^zV:����8�Q������[I�{�Tb�8=`����lnvQ|kZ��D�%kV��L��Iט��v&�d����nX��� �kƯӇ<5��DE�\��>�Ai���K������Ezky��sD�]���� ֫�4hW�M���^��	9e�Fc���g�Ю��=���7�Crc��^�S9�3x;[�͑����t���LI��`�a���&���D�=��+�dH�WY��	�v�����HE�:t<��.�䊕>����r�mY��H8���<�ش�Bl/{�-�Գ*zZ�N64��'�@���Zv&�fkJV��v���bz���R�p�N!Sm!pw���3�z��HXi�r�h�oU<�d����ɇ\�Q�|��*i��Y��\ɜ>�b�9��F�i�~��tGu�Ep�GZ2�@�M��{��Of���Z����kcT7y�R�`e��i����-�����Hou�Ds<3�]1��87x'�FN�����t/���U��W�{�/�E��, :���;����U.��	z%�=D�M�S�ʙ�j�[���nT�j��hjwEw�i���%��]ʖY<��$ECx�Ma�r�q"��d�+�3;`����͛�A��.۹��Uyݶ�b��@#;bM�Iޅ�ita=Ԃ��+5��Kr�\���,ޣh���g��}P�������/�n����f�g��V886�0ys9�����[uJ�J.�D����k7sI�w��i�̐t˙vYy����mM� xB�N�9s�L�8�ut2S�@��֗���GĎ�������L�R��˫A�ڃS<C���q��
YW�j���2~���n��������������}��!"bԱ�Μ����ũ6�+r\�1�[�Y���t@�=���F�t�%��%�+I�]�d�Ii+C���ך�o{�rQ�j������mY,+�u�^G޺o�b������:v2h��]��%4f��L��G4[����5s�f��=����n�!�W
�j@r��=L>g �|:a��Ήp����:HM�t�2�y1�+XM�	v賗I��]�䇠�F,L)OtEND䵝nb�Ü^��C��r�6.�%s+��Z(��"��[��V�>��R��t1p&�z�}�7b����j���[�U�[m�Yh��fe�m|�#Iq�R�(�k1*�b��R�S��ZyJ�yA�
����D�T*�4h�elE��U[il��J�D�YR։DR��U+Z��R����ۘQ����2�iVҫ<s
V�TjE"��˔�h�T�\�r���Ĳ�U�m(�,DjPb�J6�KF���ƬZ�-+E�)m�iEQh��F��[Tr�1�V�kEm�Z��m�O�*ūVX����Q�%Ƃۙ11����e�YqU��nﾧ��_�u#ߍ#�r���׬��&�A}A&�]ir���v{������B^��u��=��E��_�9V�z�0�~3N�����k
}������=	��!�c���̱�&�N͹&����6�������p�@t���v���� ~Mӕ�=��i��Q�>�Y�u��87v�4��jl�>�U�Dq� �9�TU��{���#ӗ�`��K�W��>�b2��s@��o���A7���{��A���h��z����^mg��)f9M�Wے�i���8�6^o����yyȉ��T]ۗ����<-%O��g��i� �+����|M��F��=�+s�r��n��.6�+�Nx}���Ĝw%<CY�p��QB�v=�y�f�a�;伟������G7��{�g6��l�)tݨ7̉���4k y8��ڋVW,�*QK�5�IYi�{T
�6OZ�GF��E�y����v��&䚳�>�N�;u�ߢ�D�sȽJ3��pl[�.e��S9(��8�eI�C��c���\D�D���Y7�>?=Wt3�^
���<��~"'��ɮ�{�J2#�J�+z�1��3쵳z�J\>~ȧF�ק�+Oq{&q����z�%yv=�y�JAޕ��q}4���sD�n�S��06�+��9r�Ѩvx�i|2�8��V�@-!�w��e���)HP��+,U��z��?���(�:b.��p��^=�Z�3���E~k�kn���u"��3L��˩,f�%8�sS[��<F��%�ӣЫE���vi�T]v�PN���!A���[�|f#�'��>�y6��zP�m�l�^��U[I�3W�5��{�;d�z���>`,'�&�!R
l��q���Cn�����9��;������&��	?n�RJ��R|��Md�����d?2@��0�w��w�w���@�$�)�C9`�ē�l�%d�0�Y!FOY4��<-	�!�$\������=�s��:�|� (~��:�u��i��H)8�M�q�m��@7����o��~$<a�&�~݁�x����:��� �:���Ĝ`(m �'�d�@�$0�kw9���rL��I����r�f�̇���z��$=�6�P���&���K�������s��>����u��ܴ��*�Wz+C?��*_���z>.��L�pޜ�<.N�&�2�}������-�{�$��!��B|�g��!<aR��z�P�{HC;a���y�8��}��=��ہ�Onj�u�Ld���<I8��� ){d��`~d6��'�C^КI����/���{���!�����̜I:�z���1��1��!�6��I�~H��o��=��]�>I��5Ha���f���L@�'��L��>@4�~`T�$�����kg?k�������~`,��!��C�N��?2�!�� m�HCi�䆙*�������{��Xa�>�c$��(q�6�q��x�4��5��l'P2x�i�{������9��i��?0?	'�8�d�C�d>�6ɦC��$:��hM?sڟ�����k��'Y>d��2�ԟ09J�ui��a�@� �<���	�w������w�CI6ΰ� �'�6�:���d���T��
[	�&�IY!�sǾ_������u�� �C�?0�@���2Ci$�7`,��$�l�J�<g��Ϟ���;���?����'�BĽ����v˥0� ���R��o����*�g�n��&��ۦ,[�;@�d��V�B�T�_Q�=d�C��@�̟�'�Y�Cl8�q�n�q&0$�	=@������g����O$9��Bu���$�Xk�����H~`u$��'
�~��g;��}�Ǥ� z�͡>d9��01�d<H�i'%OS����a�}��m������'I�&�?2OBm ��v�M'�I>Ր�C<��!��Y!�������]���`,�}����r�m�;I��6�+����ć�&0���!���wN߻�~�{ b���N�O�P?$���&�<BJ�(�~B|�=J�d��y���o[����d4��hO�~C�Xb@ϩ������T��IY'������w����?~��?$�������fR���>O�a>�I�'��!˟�n�{��u����	�:�V@=C�g�Hc0�i�P���8�Y�!��4�j�1�O~󝿷�y�}�ߤ��'�d�$:�̇�V����;d8��<��m�l<���������9����˜�pO�8_��o��n���\���o�Ѽ0��]��Knv��N>x���������n�����'�Y1���i�e$�$=I�	��FI�O�9d�-��(mL�gv��<��w�CN�'�+i'N3l�I�Bu�Ch0�`,!���!�w���{��a�����I�8�6���	�
�� m����=a�o��~?=��~��Ї�� s(|�3�u�x˪�e}U�?ץ?|�]�oÓ���{B��Uf��'�NR����v��8i�{�z�K�%)\uWьgE�Ƽ,��Z�hn�8�d��m�Ep��v�'aN|&??���n�:�:	�g+c�4��꾽���]̸��y����������Q�mL�{/����N}Q�Z���އ�i�E���Iʷ�o&ړ���郞��˟��^�]9:���~ε���������s��dX_�~��;�o��^C���]&���|^�ᘄ��u5�G:�^��[�y�r��+����(�T$�]x3L**\��eٛ���ֹ�MwW�=��TȐ�����f%�f[tGw�yg�68�@�T��]헕p6sÎ�}�Zr[������Ѿ�����.�{�|�>Η&��9k�6�jfQW����l�5��c�2��gvr�T�W�"N_W��P�攠g������:sk��b������*W��Q>�S
�0�r-���ڼܚ|�Zwb��������W�szM��{;E�N ��;5�}u���n��<�ϲ�ua�)[��$����ڜM�V�\�Q�W�2������m�ߕ�%^����+����`�Ffp�ýy'��W�_���>�+�d~��b8�L���k�i�`����hI��!�O��},C G۲W�f^��.����Rr���rO��U_V�M�W�w;��G���~�v{p9~�O##����K7���re���?~���_+�#���Us 	��FTZ��Q���O���5����l�x���0mK�ŭHD���ao����<�4��b�7_Hw*�ibn�]��)X�ߺ�?�!s�̐���B�Q����T���P���>�:������߾�]���t.�����M��GΞ��5:�"&�<c:�!ښ�GVL]4��&�m�.V���rD�|%�Q�\p��Q�}�p�D��$¢(����x�����<{�����Z���f��r�Ŵ�a�r��y��9RP��WC+N����S����t�l�WK3h�e����t�R|�fnu�d�@��\z�{pm���xȯ> �d�K8o]k1��Y�����(��zFf#�6t����A�huC��m����K�^p�$@��k�4f�g��d:�M��9^ИB�Nfpz�+u;��7���Uu��h�sqV���Opeqm���=7o��]em
���`����0W�/�g��F� Wc&\E={csC�'[�`�X�)�IV>�t{)�=���ζ%j�}�gd��nZ\����x��3�p�t`�.�RU-=w���7��4T/w�����j�N���f88��~B��GvDk:�M�AWM@X��\2y�jm�ی^,��I��Ù���x�˭����gom�{����<�+[#;�]�s9��Yx�#{X ���Ǽ��ıd1�	� �r���x�\�ư�X��д�ŵM��[�m-��772NށE�wi��5kjEP��)R���[g��:�
��ҟ�����9�������g��
�-E��Z�b-���ԕ��V�U�d9��"ҴT�[T+A���JŊ���XZڭ�����R+ZR�V%���`ŋ+ѣV)�1q��Q+Q��P��+%aX��m�T�ֈ¶ڋ����ڢ5�PR�jZ�YQ���ب�*�VJ�jT
�U��V-E*Y���T��r80��ƵDR�Q�D+mJJ5(֤Ykf&8�B�l��Z�
[��%aFKlr�b�6�R�Ab�-i5��֕�cKPU���P��j�����j°���E*��wt.�ӯw��_���s����Ph;(�E���;���J�
���_UU}|ԏ�����V�����h���&�>�h���2/�7X�VW*t-׳π�ҽ�[����#�iq�ؔ�X����K��Ee���w���������V�f�=��|�fB3��SEi
�� ���x
��fTYK�لy@;i�_��܅�-���݁ѭ�x�T���e=OB^�$ej���s�7H�n]�P�L�fxe>�oK�u���z��s�X��)3�E��O��/}�t�<nzs��@�-0���Y؞9�}�}�}Qn��5T����D�<��or(�**?�� V���;�4�p��N����+��1��C&�8����4��������˦�A�ӈ�#��-�;�Å<����`h�{���@��!95.�o�_4rg"_lNt�Z�L��'�;�؇8����l�s=-]����%ӥ��i�{2���)�
�'�VAzk�ޟ�]�m���y/rV2���'�u�Ƙ���W1�}�(X/�=Ŝ^"�PZÑ���ꯪ�D����Z�?�	��?L��|Z3H]t�?�ī�)ΓX޸.��k�o��SC�B=@��j�o�g׈~J�f�\Si�8:e�GN�������d���Dy�������Gٺb�*yQW��Amݴ/�WC�}�`�f= M�.t�oe{1l�a��k@ńF�7���F�'Tr �z�ˌ�@��v�u�n0,�l��lJ����9�_��y��Q�3��ކ��&J�.gn ���_}��UW�TnO��/�@�[�pO&y��s�q�V�8� t�>XH���E^P�+(��k<���b7֢>���}؞��Gy�2�yh������w&��2<Oo|}L{����Z�2'�I.�wĪ���払胊�53^5�0��coݰd�r�pz�7�����=l�+*J�9�ep�ʛ|f\Z�׳Ne�����]����/)V{,ʉ��c��fN��7�'�f,=�'�(�8aIϿW�U��hȗ�~��ۺ|6A�v
.�k�\^(o�5���]�L�w��Xt���{&Qa򹾽���y�Y�i�'����(o��V��:��q��X�8p̬���0���%���i�Su��.\��!ͮw�حa{Tji��Rj~����ډj��g��b��Kإ�)��9����c����2�GL���>35y���E�f�{��F%�ƫ�Ey���:D;4A��]0l�ptt�Vj��}?UW�UUv%���xJ��&��KH��j?WJ���6�SW��}�Db�7��WB�ȏ�Ҟ��sa�|j��r�g)�C`�A@d�N-�=Z颋��>>�ʤ���
�H��v{ByWoW+|��`�LPF\�i=<܄�j�Y�����r�E�Xn�q��e��>�#x����d�;���]S��P�`b��������aa GC�m
�i]٬��D�g�%@�V�A>�%fm_\��,Y<�p~�����]�y�������]�Q�5�؛p@�����p� x���Y͞Kѩ҃xO;��V��cq���]��շD4g`��B�cN0:�������#�'So`�.���s��z�x#�VXf�u�u,�wPpַ�}�Dg��7��:���y�gVc�3�x{¸*eV��dwK�1y���<�ס1�]6�t=�Jq��H���NW
R�i�����0F��Yi'3j$���Ӓ�bS{�vI.�X��b'b�˗o9lM��_}�U_wG,{����7�TY]2��z܀ެ/���v`�t:w�g����xf�栯l�d�>�mo
�����i��1�q�D�^t�>`�.@{�N���ཤ�OgY�ؿe��P���O�r�"����=�N�۩�,Qb�ɠ+z1t����A�o:�H����W/=� l&��}�����*"��#@���*�G��=���=5w�&��h�.�+��>�[�����6Ĵb��	��J��]}Դ��s����eakR�P���h�%�-W����U�ܤ�s6�~�Ɂ������z���X�9G��El$0�r{Vn7���{f�TUw�&�m?wV�2�]��E���$n�Ju�6�z�e?k{���:'��ĩ�VV	�<=�`(c�-�:X�,W��a������"�}�Fq��Yb8�ze��,��|39>C#qy�U���?�k��s27���GW��WwG^�Vza3-gh7C�B�;Ũ�&�)�d�|��6=��tk��S��
פ�?}��Wՙ�'��_�U˼B�k�Z]���bڈ�kת��]1����%d�Ʒ8�g�ll���9W�&1֗��4Ѻ��=~~'�Ԛ��^:�k/b�%f�(�.*u�>��k7�ǥ�X�Y> ����r�w��\�
����x�M^=�ﴹ��T��r�*�2�q�GPw���{+>�WZ�v����U��9����������a�#X�;9��ތÖ����툱mj�\w��D���ʓ�D��!�s���n8��!��h�e<����+E��]q�(u^7bb<��]���Z�X��P�N]������Rs��y�X���P d�M���k*e��ʬXB��PΕ��xUI�,ثs�&��F��k3�<�BP�a��E�܋�3ՙ4I�)�~$U��3�+��\�����GAY�}fV����Et0���N(~��r82M�i֞��3�U��*w2��'n�gM!�ѶИ�K+Y�b�[�*:�l�C2ڼxos���+�C4y���>�g._'f)n�c��]\[��_7���M���2q}:V�@�Qн�|S�����\�^t c)��u�/kpY�:�uH��l���r�}<R�����jE�_ͳ��y��Vn�	v��T�5��^��<�e䬎|��E����A$�b�����|p���Ǯ�W�[ר=Pd�v@���_f�c�{{�@s��O�s
��Y�yI�蓌����A��ٕ�V`���nf���3!#(��C�n�OL\*��{�� n-��7%�Kw1��8����B�|��#��ԅ�b�n�6����-K��K�*V�ㆶ;w]����(���1����PR�V�H,���"ĶV((*�ұDJ �-�b����1�R��QB�PR)E��ZQB�U�+*V�����*AZB�6�V_)���+-���mbyq!�QaU���Ũ�[`�V-a*���dU�lQaQ[L�����y�DUX��%b�(�"y��,(���kA[�f5��*JZ����-�-j�-F[R�m����"-ۍb�ʨ�YL�Q*-E�j���ejV"�������g���rk\��|��7�A�����"si?�U}U�X�N��\;�D����N�uͼ'��1�Rg�q���h�ch�כ�j���<��!8<{����x'���ۊo�E��(���-��w�l�ρ�'����t)��,��?a8�2�P�Z�������aT���)�[�հ�"��f��&y"y�t�=A�C;�|T�u�kl�|�Zz�s�^�r��Я+~�U�����\ۨ��%�,�"�%7��8'�%��,�?W���Iz#�^X��9�F��_�Ri�.����@��y	r��y�(��*��.>��)�����j�z��E�*
�b�T� r1��I�}��nk���s�"Y���g�o���%���N.d
&`le;���w���F��cm(X�gQ�PR~�g��+�f��ܕ�G�m�r�����Y�&�����+���vK�f�!�=[Y/e]0Os�����0�+d��4�ݛ��&��S��P-��U}_V{D��������f��f����zR�e�}�kb^Еǉ�7#�9V{^�1#|s�2�V}�����>=t]����q�d�G�A��;������2[�U�!�e�5�v����~��3Ԥ���i./�K�7���^&���轘��5����;��+b����΅���zRn�����fOf�X~맜���u�(F:��E{ٸ�1�j��p|n��i����N���-i^�9{���vI�ϛ����^.4��ɿ��d��K�s%ˑ�=Y�y�2l;��@��kq��z�^;���3����hx�� �����#(/
�7� 	�y�T�W�_N����2�<I��K�㋁���S�{�։��{���g5�^^��L�y-�
��6�j4�d�SK�&K���˰D��1n��"�V�^}Wn�-;���=���){�7��N�6�?V���͕}֕qt�9�7'3g$c9�vY�M�[�l�>�'+������z|�6��1B��Q9��O��|~ 	�׮B�9���ڱt�3yV�X6�(~�Y?�Vw�o=�x����<>��Ԭ��Ϩ7z�]��j����@`��:��,U�-��V/*,U��b���_*�\j
��}�Lm��0g�j����+�Y��P�3��n�酇�>#©
|��<,l>���
�s�g��Z���
t,B���E]�Y�|�4���� b������E���O�o�m��4R���h�/xQ��
��_R�h����q�qR���f��Ef�9�R�j^%��*��R������n	�%�I�.�-�N~����/��Sǔ�e�f�̾��v�'5C���l���yܞ���	�ڨuި}i�y�]=Nf���YW2>�[s	n�W#��nd�����_'�U���
PQ��*=F%.O:Uu�=u���V
V����t��\�Yf�⏝N�|>g)׏ɧlҡ���y�Lթ�)�λN>��gنn��M�ȫ��������vi~��q�}�s��4��o��[���w_x��4�}O��x�s����.��7����ֽ�����9�Y��{�z�2�l��!�E�&�
����ru�z��?!����}��d�<װP��$�z�>fL�tD��K&�N~���'75��������٭��X�b��?D�Ϧ>�mVh�+���Q�	r
w�>�a���<�p�4�`u�ªq�h�*^���F��y���xu}p;�����C���`�SL/�u߶|���+�eMwXc�y����>���^�@�uw񃾺�Q���r娠4m�W��{�v��>uX#6 �
B�|�y������ Z�P~7��M���rͫ�0*­�FL��gP���;t�iM���ji�麥�����u�:]�O8ZHՈ,xU�.�Xkx���&ם��0{�x���1,��t$n�U�p=b�ħ���^y�
��^��o������a�7����������qo+��r�������*��n���Mo^�k��k��8���v���g��M�<N7ڼ��Ӓ�'�v�ܺj��{*�������C��� ���ʻ�)ڻC�W���A��9$���V4�����Y�*�%��|sy�d�~��:J���h�}�[�%ѷt�}^>6����V�ee�PW�n�X���y9X甬"���W��Xkʕ��@G�;�<�mX�kEz�@l�Y��B��|xԒsIf�ϻ�:�t��&}�<n�I��:�����S*��]�"���0��į��D̝G\�RR�r摾3�.�l,��c��L7zx V7����
r9tw�z#80=4l���kY���!s	~I�<����6������{ۧ=�����%o�6{�jY�u.��uL��>��Q���=}�9��w�M
�f�.�b����G��{���ɱ��N�7V>l� X��|����b�~���Ё.�n���WN�P��0��u��2��y̝�4]�&���{]����_k[�x���9���Qt����|>�������l�웖o.�g�W�P��^gwO;Nv��k�={�כ�����Vst�\8W��^�n�[qL.�÷�쳂�9�ӹ�J�7�Voj	�����8�rJi,F_7z��J� XN�n~���ԯ��ʅ?���u�U��
�M���%�rgX{��K޽��ngQ�ˬ�2��6h
�����fE��g��/�����֍c_AV5'_u�ƫ)�B
C�C5��p/�xQ��`�j���]���G�xA~����W�f��W���U-I�_s�IOu���Y��̪̾�>"�P�6{=�Wf�hي�4hz�.��������/$���;�h�~�?j�V�[/MV
�N����^U���j?t�J����*5�F���5b�݌ ���樐j�]:�ϥ��~h�>����� Ek�~p�
��fd�j�i*4�]z)fϮn�ΜCV�Q����9'+sv�1�9�8�R{
[7j*Jb��Q^H��U���:�d�w���8ux�][M4R�#6�Y�Ð�2vK�&p��R�)�\Aa	LX[�_L܁���11�����g38V���즷qeZE��r��㦵^�l�r�c�����O*�f�G5�28����D_\Ϋ��e�yhA�M�/76�n�8PPF�0<�q1`��vޔ�M
K�%3/>5�O.]�=��c#��7��'��t��N|N��N�ϖ���GVd�[G�������<R:xg:'�E��-2;bmw]���p��H��keG�j��Q����Zt�����m)���� ���/��n_g\4u��Zn�?���[�����N�(���Y�V7�d�&��b�����G���S]����7h=]\���M�/:�Q���f��*۱��N;�H�)�57��((ގ��6YY7��Uͤ'ɷO����ͽ�b��4��nR������ip�Z�)k�JEe�u��%���k�;<V*j1��i��Ҵ����<�z���P{0�]���76��`������P��2@��+im�E��k*-cX{�Թ[ib��*�����Z��l��V��|��6��|h�(V�)V"B��*KU�,QQ-���(���D�E`�C��Cư*UdXT�"�
yhb�%g�)"�R*"�`,�E�!��`�-�ĕ��E���*�� }�U6�g��y@?R�]��&���ԍ�,�.�8�nj���OOxO�����?
�\�_�
�2����yV�yF��>c�̈́Maj�q𧄓�LV7�����7�yr����z%�=|z����EES�=��T�<%��%�e!��U~6�o`��7��б��}z@z���j�_V/���^�I�;�^?
��P���׸�|��ƍ�>)V��x���-�F+��x,<*�V�M5:���W���<�m+���|=\ ���CS�����{���_R�]�Z�f��e�M��kt`['�W�Z�3�8(
�!�o�~T�`Oʟˍ��d_�^��b��3���	B���RZyNM
�s^��ы���Mّ'd�R������hJ7��$����UX��_LW���k�hUi�D�ռ�ߝ���|o-\�meU�6�ܝY�7�v���V�+V� Q+��3N#U���{�}��滭ϕ����)��2�Lw//Z1��J��^K��`�8i8,}	ׇ�����=��L��Wq����x��*� TⅇB�!/7~k�ҷ�x��ޗ�ӂm�׹�n��[����N���G���u����P��s�G�d�����KV/.�V��#�p�<:���Y���'�0x�q*��#^) u��Ƚ8`^��^�i%���	��x��=X��n+�����;�T	��cX���O:!�d״�A�WcJK�f"�����Խ�Uv�A�A�xg��4�o%��U��*+���qR��Z4���c���r��&���(���d�ߜkS���t��6��%�/n������]��������o�SHֻ@N>
�+W�6򼲞�S�tp/W�OY��tX� ϕ.9�}f���ƳOvf\�7J[�u �G_����]T"��ߔ�P���sTlۿ1��S�x�-]>�� d��R�Qed��9z�=��h�LU�W��>xk�D	6'����A�~l��o��6�޹u.\A܃�WC�����UM|�Ñ�]_��!f�v~���Y���f��pۧL��.�E������-���L6�OhE.������x���G�ͧ榇oɯ�~C�W���<y�o�vޱ<�{��o\�{��so�%�.ݼ�	��Ʋ�!-__]�!D�Fj�j�Sʕ��w�_��&��\�{J�������:��:����.��v�x�V�J�UpZg"�W��A)�)��ޯ/,�&�쪗�*��#�z�����ËN����;�W������i���
�����73���T%��V��/{)\�e
�@��4:�#��~��xr[�VY��]g,�(|s�N)���Mg�5���m~����������5�i?V���ۛwBg��1�:W�F�4�B���(4��	YV<xbv�(�O�U{�R��vI���;�tY�o����iɗ��s�����?^��w��{��iG<��r��㴩��1�ꉯ������R�Bz�2�Vm\���]-��B����E��o{=���~
�2S{��l�ۮ�f��fC���\�O�X.����]��w^�PW]+�(����w�i���1����na����5���;ݹO����)�ϯSk���Z��Ki)�\_���{9ҳ`��^0h�}Z�U,?p��s^}=�ާ�� �7�����V{Wƅa7�Z�\$r{�ԙb�5�O�EZ�S�X8v�(41]K��S����Ϯ>&�Y�t�jߤ��o)=�O/I��g�����̎]�2��1x�G�r��s���y��쒿��-��L��n�����i�ß]:�@][��������p����ǫ��[A3��z��1{.i<,}�֏��àEA�Up �ؾ�7W�;|$YיK9W���C�r�ẻ�Y���e�^�C��^�c�,q}n*�@���Sx
5�n{��DP��ذ8~:�4J㣅V��>|�ᢧ¬/��
#g����MR����x�?0��O�J�������.c�\��a���8+X�Z8jK��ׇ��Sݘ�z�_�%Z>�8�T*�b��fM,qZ�f�zP[�Co�2=��
p��SRʻnb[d.��kf�����( k8����t�V>E޴�{�x��ﾀ(S��]��=x������Svkۧ����7���=���s�>n��~����.�+�B�ל�5�u/n{N��KV/.��wN�R�\0WL���süh�(������3\<) t�����+j����<+�A��T��J�c��f�P�w�=��f�N��/_5Jְ���uOs��e'����f�h�p��Ӯ4EA�~�Wt˿����О��n�~��4���j�&�`�O���#^	j�0�`�~5a��Z�ht�U
�h����~�5�tAX�P���$��M�9�w钏Br�ᨔ��f���Q��^c�v'����Yu�B$��"��1H�+q���T3LQ��*���>[�ghoUe~w/���=޷����lߠ��
��]+��
�]���u*=���D�|j��Ӥ~�X>��(`$؜�a|��2��ec�Ɏ��l��[���t�)�!��o��Y��fk��Yr����%�ׯ*�_����\<-�4P�Z>�]��c���(VQG�5�V��3P};U'��,��u����9Vi�z����9��>�~Ik�"kA�e�eUu>��o����&���r���v�����!:�����@d?x΀�p
2�P��=�3��U�b+t��V⩅�rvM��!*��'$��w\-&H�����%p�*"�ﾤ�H�U�U��n���!��/~��(�?y@�1��B�����N��^��J�W�eK�UN,�r�u �f�&��y��ˡ��c��w���M���]����kV+hX����!m*��]�t�18���c��o��b���{C�X�� ;�Ź���M���Cᆎ�Z=uJ뮍� b��S��N��+��W�\xR8$kQѡi�{#���hJ��^�	S�k'Y�G���}M;�ҿ{��4�k�ƅ>)�V��{ʕ�L�2��v,��W�>�F,��iq�x�6V��#�F�E�y�9�И�ms`~1k�#�}��QK�A�~j�h@�#���Ӥ�?#����Q�Gzw�KN���[CP�v�]K��t����J��yz���{{�o�mͽ�����׮U�b_�i�ʺW��L�<�V�^:C��w�^k�f�O՞�u�38�?{�`�Ҥ)��koʘWʰp�,h��dI�n��C`�pT����S�	���3:�g�`�? EAPh�[�i�kh&xR�sSW川����WZ���� ��M {]�.��f}���}�C���������b����J��K�Ƹh�}�q|m��-��1�3w��z�����cB�u�X ����t/>����u���^��mx���O��^�3�,PsiA�.��.<���%�G15L�f%Ƕ�̦^�����%����fY$n�m���q)����Π
�]���m_������#���L�*�ʅ@���f���:�|���{M��T)�i��)RѺ��vYHS��t��nȒ7|p�HgQKxT7�]���̽Ÿ����Y|�CJ�@����]k�M�౅VY�^�,�h�����˙Ŷ)-Ï]�����ܔ�oZ|Q��
��O�#���V]J�6٥����b1�CS���>�*��#7���]Xx�˼�����;�9�s������A���p�<�$�B���;�L� rј���n3J��U��o:P�B_-����nV����=Yw^+L��.�l��<��X�*쭭��܀5鶵]���֎3pn�@j�L�j��h��p�56���o4�8ͼ���s�&-�즑�b�5{�ث�ve<�yIF:J�ۉ���Wd��Qt�Dv��ubb^�}��Oz�wb;dz��Hs�tD=�;�4b���\�B�p�pv#,!J"mGy+r�l����+x�8���&y�^=׷֬�鵺�2v�wF����7u�������������s�~���(�E��,6�Ȥ��U��x���+*��[aP�����aQ`�,�������,R"A$X�|�ĭ���F��ڪ*(�i`�"+ ��e�eq.Y*��رH��"� �I�Y1�D�B��P@�|��C�{��oׯ�fzf4���L�M��i�-9v֝1����`��뗦v&��M�Xs;��<�w˽/������}��u���r���S�N??nְ���͇#�wz��x��6n���I`�� V'�L}�hA�tMp�����U=������S�3�}ܯ���������N���*e�w���WjW�<�f
���n�G��E�;��\�)Y��7���n�h`���^X0�/�SƷ�pZEɗ�\;����#��aS���춫�q�[�m� k<)kX>t�k��9EHxg<;������*��<��X����{GT��6}�W8�_<��E�V�<�e�����J����p�J�=4,`c��)_[��j5A7z�e7��/�1�.�U7{�����YJ�Uu��m����2(�aw�ݲ�٩O���/��"��PJ�JW�<�{�U��
�E6��g\j�y�l�o�s�߇^�_^�f��G0�V.�͂)�Q����񜫺�n�
�q��,��~%����{�xu_s��Z�yr�7B�w�̦��'%�'�'�s��W�J�j�՞�T���9�ON�'�U!�k�����K��h�����Φ�u������^A���yGB�Xq��{�m�3���<(|�:|x*z�'����ۤ\�,vn����]qWx���H�<5�7�K�',�L�ð!"�9�=ِ���u�׽��ȥ���i>�?2�����
O�|�5޹^�f���un*ก>��� �=T��l�n�ӽ�=��Wut�Q�<wT-U�]=��H�/pp`���HYW�i�TCO��{�L`�*�b��>`������tf�V(r�v?��O
�|��"�R�P+²���O�u&s��
���
���
�.��_0uy�R
ٞ����R�^�b*Ɔ*�H��W<���ww�:�P�Q��Z4<4��P*�7���=�����y ����|j�U�Z.B)G�ٶ�ڙ�wJD�d��溦P��}L7��t]��Y��dRC�4{�x��<��o
���gj'?�M���uu8R��J�U��x~�����ۻ��wȷ�_�~�@Tc]R�N�γGn޵��}�^�W|�J��C2�]we�3*_��^دc��wg3!y�k���&����5~p���k>�s��>���ޛ��o^&�uO���"��>ǲ�{����� ���v�
����s{�!���Úϻ�rx��^�5��x���#�����·�<��^��E5K�3^�HN5�xu b���#�
�!+�j���U0�J������.�<7O�P:pB�N���᭡��>���`��󗽊]��8�����`Bp��oEF��p���MɅ�p�6ʨl���l�)��T��r���X<>�k�
���i���+rz� l����t�P1^��X3�f��pg�x�~J�;54�t:5��ڤ+Fi|����wuA�4+my�H�R�Ձ���X�᣼r�=.�*�NfO�q�tלͪWI��o�����~��W��j�U�'������u����^��En���*A.��A]e�`+<>�R-��mS~]�t��vm�Wn'�X���9R��������C���@�p�����:~�^������p�8W��
�X(KT|�W��
5�to�M�붮�J�S)	&��6y��s�s���y_�[�>D�+�A��:�GT�F�N��y�z%�����1��b�U����ǈ`"3O�����T�����a~�
��Lvo뿝���e;��yp?���*o���[�����3���M��ﴯ]?{�!z�o��b�q���C�4AP��������mT�y.�˳�ẉ���Ghz��Y=~~'��������x&�a��YZC�\)�R��*�`��S��uTc���`x`C�F���L{�u{ث�F���CMO�見�g���c7���*1�yWt�_���������g{���O��2��ƾ�5�tV
��I��V<�)���Y���<Wj�Hԡ{��4CǇJ8��gfa���䷣��K[˚y'爵��{��y��~J��S^�7�<�.�MY� +�\�j�ٛl���� k1W3�P��G�߬JH۝�Տ��'�4ϑ�3lS�E�|9��w_zu_���C� �ʸx-4����Ug�7���Z@Ѕ`ь����>U|Z4u]���7ϵf�����9W��]7��wt˩+�a)�+��+{��6��ut஬/�
�C�L�|wپ�qA̡J�/	t��ʡ^�B��%z`s|qJ���A��X'x��<'�h�-�{����1<{o��ǉr��}���t��w�ݗ��w�cN�Z� ��8.9���maa�1d٦2�j��r>Gn6�5�XG��n~���v�=J�!���x`�ߚ�2��*b���:v�ݦ��C�SY�����}�_����ݽ�U��t>�M{xh���_Dm�+³����yx�'�R88�|h,���.�ҿ�/T{�ES�.���Vf�Q���º��V�z<��S^ߜ}v�oʟr�4R�.��9f�ݺ�x�_s}ϙ�Ζ|��9��)wO��/��^���A�ä��>Y��Ű�t�1B��,65�k+R8�/��vj$�P�+ �f�1F�x�˃j���C�]���SKK�\�LK�m<�C���V`�CЬ�fX� H��V�@�PL���-��X�|+��U�hԻ�PW�|%d��:T��%�U_}z�=��>��4hT���A�3��@r?;5����u��I0}^y|��.�2���30�����w7滭>}|xΖ�'϶�+]j���g\<�1�D}Lc�e���1��v�	��6�k9�{+� �T�k��=��`���"��/���]�����#��X*����4k�"��l=חб^&�Zk��k��f��.��{���^+��k�����X:��p܂��n����v��vA�0W���M�����9>j����}f�Rpy=d�Z
	JΪ�7NbH� x����awE�o�i,���\�q���l�&wj�+UIuy�$�꯾��8�q\с���/)
pK�t��������`�lK�h��Ŀ\�@W�lۧl�UM{Mc�����^x��_^' o��hmMu
�W���.��s=�g'��yz����p��n�Go{���9U!�{����1�|kEze_��טM$|=��.>>Я�a;n��v����;M4| ��X���%��Py�' y�J�we�Y���aU ���C���3��Q�<p�U�Y�
��-� ����*X��{ӆ>���<����
Oʞ+�|0^�Pu5�.u`�<���.������yj��jٞ��p�a{����6[����X�y˓�}��lَ��̎���-/��������pV-�=L�
wk��r�F<�L�e,���Y�Wm�y�aC�C2i��a'���A�jYf��*v�4)���;skD�';����OK/1��m��9�@�+*�D]jzl�
Z�gV�Z��x��<"���z�\�����j`�e�=��Esx�bꬍ�9^l��λ�j���']��R!�
�E����g(�L�v�ʇ\Pm��ݚ�y��J7,z� 6Q�����z�Q�D�T�/I�}�GL��&��jg������{+�``���/H"\�cv�t�\��hW"ɤ�h�JЪ��y*m\�1]�E,��5�4Y�[����k�7�F����8v������Ǖf[��&*\ݨ����2��a}��l+����(c�D���K�:M���ʇW�آ�0�����t��{'Y�³3���>8Z8�<�&q��a#:L��kV�����m�sPuؘW����e޵�� N������zjح�{5n̄+�Y\��h�/Z�6	��p��J1*�Z�֓� Y�����K�\љ[�;�wpZ��9��?g9u͟{���֧�<BV*¤_r�ʄ&*IP>IX����,���XVB�*���©nZg�d1z���R��)=}2��U�Z��`��&2�XQ3&`�1�@��c(����>�B���z��1������8�����-JK�e9?�U��Y�=�Lul?�t�O3�|\7t��ӧ���7�>�m����*�}�s���ج�P;Eq��ĺ�������K��Ҿ�v��ux�s{3��f?^���իw�.���tn���Y�����{�]p�4��S{�����J�5K�8x�7}��>�< $�?a���xR�����k�����e
�F���̚t��G��1O</�w�}����e���U0��`Z�뇅��@V�m����ګK���n���7�ۺ�
�s��Ϲ߯i�7�t��g/���m4���{kݷ�~�|��/,*6���A��ղl���5Zݐ�b�}�ݶH�ϓ�B�t�p�l̵.�v�.V�֛}�� ��u�s��e��i�ǟ��uv&�ja|xU`U�Cӏ��g/��GZ��.-���<{N
2�R����@M-Z�����Y�=}j�#2_�S�H��c��A]��P��R�!,�`�tZ�͙�1,�V�K��Ѭ8>�/�)VV���|���]x��b�!CUa�a���~��;���m�*��%����5����
_�_#��y�v��c��GF�����Uo�~5;�x�y�)���<������T�ͫ�r���x�����N��뛳�8�i���}���j��wR��o��Xa�7�v&�)�x���9����l�R�{j�`y8�_CD�c毟���n���b�Ԧ9������[�
_�2��o������H��R�p!+k��IVYb���x�<�W
���h�`
��q̻���>'7̶�iOi�;x�]�=�5��T��-P�V0Rָ8k�-Z��*򘗕WQ#j;�� �>͋����,���װ�ՏmVn��
Ѻ~��*iU?f�Ɛ�T˞�9Lp�,m蕝p~}�iS�o_~���S^]���<Fɮ���X0|A�A�|+�V�Ws2����$X�t*�r���et�r��=J�VCb�k���=��6 ^��3^�*���xf5��3��љ�"���4W�e$�a�Lv��F0l五Z���:�mٕb�G,
�qi/|���9����o{ީu�Ό�­%V�Z<;bѰ�h�`�t]N^�4��<h��O=�T��{�|gr����<��V�~8nY����t��(��껺�3_��	p;�+���z�ٺ��	��C�?/_�鯷�1��^㣁�)��T�ģ�Z��ܗw1W�Uy��k_>�پ���v����K&ĩ����<�>�@g~~�X+d�R}3�5F���K+�w��g�نE�8�%f��v�xtP�Εa7n���N�R���w�x2��G�{ro��nx�ꏔk#0V�纉��@t^��˧�ɨo=ۧ
m����%�'�,�_�86�?]o�|c�[�q�k��Wq�Y8c���V4�f�/��f{��9V4f>��1�
�tסjp�}3�{�u3���a����9f�/�AO&K�P�D��V��j�
�I�~N֮+�U정�,E��Pv	�yv�}Kݧ3�Yd��fOQ����/i��bz��g��:'�`ۯ_nξxNIl���N�h/�]3;+e�%�K>��7�㗋qmZZsV�����$Y�IO�}U��L���^�/j�ԏ��䰐VEQ�z3ycO�9u�ȡ��<�PE�,(�����e�m�o�l���TW˒w�C���N�:/y�x�K!f�Pī���k��{Sk:���(䭷V�3�hbV>��w7~�wDezg�S�J�:*;�),x��=�Ԙ\[[�����eg�@>��^���@xbw�7kx"��W��p�R��'j�}O�V�.��q8w6�=5�S�0H�����t��O�_܋?hX8}<�lpң�T͓�����W54y壾��+�&��Z���iy�X��)?v�7�b�OT�=B��u2�F�Ў�p�K5}�D^1���+Ӡ���6�KP�ƽհ!<�ojWy�"�G,������T��#�j
���
xt�6w�D&������K9M;�Ǥ�,I���f-�zp������1�GYB�}���~ӭ!�e�U�JN�A]@Ĺ7�+"�T�gr%�t�Űھ�H��,h\[r����7�Y>�8�v��.���Gk���e�����Iy&lٞ{G���a�'����̾��k>!j����j/;�(7��V�_���jY�؎R��.�{����tK#Rg/�3��IM&2�G����2���W��^�Z����e�Zh9�^s�G^<��ԽyZ�+]��o��}-8/(��\E.���=s��s����t�
����q�C���K��dI�g)��9 ê^��BL��Y��و�f\�oN�ܬ͍�����qb��&��G? Sr���!�jg�U���ڊa�A�w>b!���n��jf�kRc,5�.�>�*fڸ#����=Ƃ9��C�GA��ПN"�l��i���z}���������5������w.��}<���-]��j-��(VA�n�U��yY����}�5�w��({�#�F
7�'7��"f�^R�`U71��]Փ>�N��`�Zr��7�k�mg7�Ȅ�z�}`�A7{�Z��n�s��eE\�|3k��&�)9��+��|�"D��3��ծ�v�̻l�������۞�����w(��� �y����Z+�pC��W�U�)G�R�Wa�#xT�{ٝ^#�J��l�ҏ����T�.F7��fִ���^(�����
es�\�c~*�0q�֏��UL?8Q����_�no��g��W�t7@�f;�����M\n�U���q*�;C��e��I�3���F,���Jok�);�b�h�R�f>[�+���vn��zZZ<��.����}�[�����}y����8�X���Z`F�2���:���x�ml�g���+@չV��^�0&���M��mb[QǼN	�NT�}%ÐG����<y�f]��6x�p�t�W�K�Av��������t% Y���g���WF����1Xrث?�#�Fu���<$V���u�XL^#�/9CZ\e��Y�k����e����^nP |�;��7|�r"��d�W=ر�+	d����Zz�Y�f�lQQS,�
8.�Q�8JUT�=�wvهL�z�:��C�m_4mI�^�[���C"�.��ݹ�t3����qRJ�k3�s�iVb��Yn�lM��-sp���u8Wos*�^��jy��T�:٧�2��S�}!�ۗ+�ڮy�y(���`�����r��˻L�AJ�m7�4k�+�7�13
�Ocb�������=C�ڶ����]2�e���&��[ud!�6�D仝	{�d{I]��k�Ve�ER�'	��p��
�S��k!� @]ז��\m�W]�̑���̄��)���5��<���Y+I�J��J���X�n8��Xy�a�Y�,�%J���Bx�QE������Z�L���a��b�QƉX1++��m3.0ơ��b�&&xV�`V�D*k� ��1�פS��ky�/�f�tkL�S\�|IN �s����V�C�hrfw�2�ӥ����FOAS�ݽ��ʘ,pVF�!f�bOe������s�bz;l�ٷ�o:�+#��؛\T[��7���K�r�H�l��N�"x��#8AE�U�d�LtS�PWԲ�������բ���ԋ�`+�w�Y��Z<�����u	��͗��,�a����W�J�/h��-e�|������K��Bno+�/Yw.|T��n�5w2��BrQ9vޟ��l���|�ߡ�Qv�	��j^mF3^R���_H�;�OY�NM/�c� ����oS���ͬ����D�{޵�r-z�O!�{^5��o��� ���g'Æfnlnu��/�?��O���Od�EX}�L������g��gk'_�n���W9��vzg�/i;��fU�1A�+�t��~�3.�O����&�U�B�"�v21z�����lN��ݠ5[q�+[���P\��W#��Iy�Ǣ���b�g���h4�{�ff۔\�m_?F���r���:=�kQ�v� �".	@a�q=�<�(�_D�~^�PU"l�*���ΌR~�WJ���w�oM�tX�k�=��d�N�;��A���Ք�
}�������\�(?rꓟD�o��c�q��|�h�/u_�ώ�=s\��]��h�'}tX��30��mOL�b<�xWW��V�{��;��:�J�^=��;q�9�jw4��4�%X��<��eCJ��ލ�$V#ӽ���B��οQ7�ml����M����ݤs�~�%���A_�@�B�9�k������]c���.�C]����Ӷ��@�Ȅ��+�T9���yk�K����L�[v�u/_o��@��S�h'*)�*��/�(lu6�7z%X'\�·��� �Bn��~j�R�D���K�\��3*�$�#�qY���Hk,v
c{�c;+An�:z��n��:��f>4���P���r:�~����k����"�a��7)gM�wӝ�5�T��]7�%��X���f-�Я���C�x�����Q�(@�RE�g�<�#{[�sH�^W�M���T��~ ���׷g<���/5#���z\�_)=�=���[1�v��4�9��7$�X{X�L}�קiY0�a)[>����Bnh�;F/6�5�^���`:���;�R�V�[sue����}�Z�mgE��dK��E��o��Ū% X䵩g���]��s���G�3*'|
5�G�ݶdG� �����4�\M/3�<ėޥn��y5��+utO�%�zR9[w}�AZ�+�w[G�R{����wX`c����$9���I�KO`Z�y�4p׷,H4�(���(oL#��� ���4�f�z�N|
�����%�r��hz�7+����}t�[3g"���X�S�a k�L�;���4��K�NՅ���p�E���'es>�������鎷����+�P.�Yr��JI=\����:H�'����K�r��wDgx���H2�(�]�XY��7]%X*&_����xW �H��i��� -���R�~��z^���̈���_�M���ҁ�վ���?�)��[��x�5��֢+J;щ��c����2U���^Gp��oi[8�Pt���".C�<����[�q��k|�Es1�j����ET�X22ܽ܅uF�D��׫�����L�vg�=�H���Տ����y������m\RO2��`��M=~OQ!޵�G�\�^X�5�]�G@HN/&���
�x���,�q��`����@e��O�yKw6M�Vj���'=�2����:��qѓ�S&;g=����2іpS��{#��	���x�����4�~,#
���
ג��vY����pn�y9x*&\����:��xh{���Hh	s[��LDoud������<�m�����Z/���N5	)��x�v*[Tw�h��dn�p��0qѯ!�裯}��I/<��u>����'�3ۯ�uwQ�c�Ut>�p��i>�G�C�[�3�ozק���"�������U������}ި�M򮘰�r��}4�ݯl�%���yzw�r����1�	�)c�j�n�u��)�w��JU��Z2^�y'�Q.G;��Yʽ����ǯ�P�	�)Q^��+��	*�Q.�K�*�������v�@;�7�K�bTG�<c��w��$��U�c}�T���8��V��=��
�m�.�j^��j����^t��3G�D��4�+����%trV�8]�Bj>����A���o ׁ\�%2���,X9�dב�����ʣ�yl��H-���/�Q�wWV,�b}+�j�M�mc�I��ɀ�Ŵ��@�(�ӗ|,���B^*��u)
(�Z�L���bg0V�!Bv[\x��h��� ��98�ѿ�!ǹu��70���(��6�����e1�F~���ѓ�c9��{0���C��[;�f%�[��3�ҍQ�6���b#���̗j��ޤ��ݏ_v��ȭ�|ܬ)3O��VP�혴���0�7�p�Gy桯+��9�8V^d[�V&���R��iGN#�͡IW����;�9&f�.ǈ��q_�P�O�-�r�] 9���{�i�j��nm7V����v7Bv:�ͽ�z�pJl���p�Նs2�ݭu�\kA���	�y�J��7k��:��h��>�^��o0f����o}��t�s��g2��"��-1vK2]ii�V��+�!f>Ӧ�8�����F�,.��Y��f��J���;oD ށU�Ӗ�r�r�uq��)٭'M0m֗-G�i���<�é�R�Ho{���(U�����p�x> ���;w�)��矵�J�o�4:��1���)ӪN�ϲf-�΢�h�Y�L,��3o�HõI�nf����Y@vy�7��^�;OiL�+.\��r��eSʹ�2�QLm���S����`Y�`*��YD�����QR�e�Q���y�b��S�Kb�WW32�`�e\��Ks<|���c�K-�|�0\�3.>>d����q�R�f���epV��e���������Q����3&Lr�s��g��X��QYK�cZ&y�y<W*��)�|Ӊ8x[n�8y�Ag�aB@:�5����~�A�����FQ�����'��)o�~�ﴺ�3�h�/��[kY�s�W^qO�z�M�2��(>$��]5�sMb��O�������炽L/V��F��Q��,�F��]� �XǛ4���.v4��i��3{�X�k����#�<72�-Mk��a�6C��xJ���k ��t.�X���gw�B��2v��h���.,՞���,�i���5��?l��g�4A��CP�5����9nVg71��z�D��u#��J���p�� _)��;����'���}2{��(8�g�*��J��o���ΜU�h�#:[s�2Ӡ�k�5��|Ws3��JO�J9�i��m0�I���z�,�{��M�W:��W�g+n�9O���2,c��wk�Tk�.�f3J���E���w�����;�r��=^��ѭ�`�ԧ^�>�=n�R�Xfc���A�t�
N�Ǫ��|�Ȑ�Z��u�gdCI�+�3��I��,84A��CE��y�$k����Wހ��7��Esx��-�tDFu��
1YB�.z99ċ��;�#���%����y����ڣ������9l^1f$;�+��w]�z�k3���"LR��;:?����O$���� {P��S�:nvOd�U�^��=��f�J_��]��蹧�k��P�qx`�P�/lVE{�=��9p+E�h	��kY�E=W�a�$��e̚/����SqotCt�Ȕ�tE)2�F<�P��Gw�@�s%!R��!����O����I.��`�{{�OJ�"哊N���4OP覐s>�����I3�7$�)p��*��d��Y�S۩�޼�{�\p����ͬ�+���������Ҳa;�fh������:1�Ct�PT{c��>=t`:*'
>�FlS����{�}�R�����yC�:b��*���VH��Cr�N�JU���rt��!�,5�I^=��֢�}�S{L�[3^5���'$޸�6�}~4�^�s�+�2��(f|�p��w���	5$y��˾�ٰ��R��!yc�T���1��7T��}���b��H�=�y�)ͧ;0j�kT^=n�ߞ�������D�{8��W�/a�X�X`�OUv9�ʔ��pw4w�8���/e0������'�ה�.�����1:�6���Ai� D� 7�ޥ�/jWN�Y�����Aˀ_eI�1%��}�r�3����#��ǆ�` �p�^�~�ޫ��3�>�I{k��(ˤQ�<�G�j-Y�jƹC�}�&�m� ��܀K�KWfӖ�����B66]2�3.q�SKx�^�hݺ��w�.���Au�a�Jem�������*������E��]t��pТ��{�����^�u�v�M�ǝg�RcXGy���W'�k��ڱh��L���㘈9$\�l�/���v0K\�9qȏ2��:�6�nl��y&�f8���r�,�5׺�)q���l��E�Ֆ�����[����զ�O#Yr���{��%�>7\+:#W���Ȇ�Ow��F}��
Ż��Y�{4��
�J=�v�y��p��T�>����bу4�*�^[����V�|o���.@#��fNM �H�MW^��d���K�0c�5%#^b0�%��~�)
w뽝}y��P����LY&�,M�x|+�i��!ש|����Ƨ����+��rj��{�'M�M��k~�2�6�aV�!n��٢ ��*7��i�|<09�h�I<�E�xѯV����>���TL@�n�<;�7ڹ�������^-vU�'���ջ2ƿ% ��2"k),�/E�����Yk�<X���[k���Kﳗ��>�揄�f����l�V�zQ�|*YXT�O�Գ\M�&sn�?u��n��M����X�
�yz0!O5d��S�N��<�:p�	��K0��ޙ`h[��Z��Y��g9,�@)�`@� #j����D�[�5k��DB	�~�M�>>��A�4@��a7>�x��H�.��n�z9��;�`���R�����q/�Ϋ�y�����Ԓ��3�tז ��j�0�\}��%$��P9�����c�\.ߪ'�r�����-�#շv{Y�>���ث\"��[ʎ�\P�0-��g=�bkm���5e��b�w�����N�b̢�a�bn��)�����P�͏��
�nAWH��y��]��p|�2Q�<��1����Ǳs�w���7:l�>���^�>s,9�����<������Κ�)���u�:a`�6���%�]�� �3�C�ȡ7�.�n⹆lgUwMo{��ue���ś����]�N�:��Th!��E���y��#<�� �p_5�ɦg��V�����[��"X�]�*G �f�>ʿ����~�{s�5�3�i�#j�q�av�Q�E�	�}N��ñX\@���t�%)ʼΊ��[qm]�^�g�z>�ے�fr��t�(��L�����&�ؗ]_��0
�v��f6p+�����3����Jڼ����YV����j^Rd��E�;r�euԫ����0o!���tb/�tH��8u+��}N�����d�-���Sw6�낧@v"xu
31`}���1Y��:�[�����1����^ p�t�jw���W�1�Y�VR��r�t�B�[���2Q�$�J�nM#rK�rTRSZ��|+j��n���|jKOz��mv��veE�_F�1�C,��D7�[Pmu�t�A0Ft�N�Y�Ë�u�^��ǻ��v�l�&ƍt6��v��$wNN
�Cs��u����2>i���cį6�R]k!�9��#�}ϋ3.Z�v�}k2&�^C�:[%$�:)-]Z򥇼T���au�]Q�S+F�f�IZ-���6�R�������ĩ)�ɬg�I��n���[���_j��Ω���o#�T���;)f�7��ԥ��!����*˵�.��^�f��7���f��^� b��Y.�w7��z�����u���7]��\pQ-��i�(��e���|��Ƨ���e�)\nR�p��o�S<n[e����Դ��j�+�m��<����-qq��P�9�!m�3��բ����(��KEb�|�2�Z5��.8��Dˋ��hYZfb���)j��2�|W�m�ۘ6�l��e�(�sSmlLL��R��[K�q��d�@�h�� 5zg��Y�Ӧ��iLvv/&7��Y%��ԣ��!���ی�W[۟]�wa���y����^��t�7E��N��5�^P��]B�zA�d;*c�(�����胙
�e_����R�՞�<�xj�+/�O!7��߫^� ]4ݮ�n"��k��W�	���d��J�t|��F�]&��)ڧ��Z��lu2��e�J��{�J�(h��EL���B�f�S7}��n;Q�$���yu~N]��:�XY��׶��G�d6⋜�t�h���:u(�flo��M]8�]`�:�FC�>�K��r�5}�&;C{�)޷�ڈల�a����I�N�*��>+W�A]��hڡ0�o�M�������}�p/>�+.�c����ip9}�k���g��F�tNG�a��c���w��Њ�9�v�ӽS}�xѺ/���g�Qe_?RΝCu�u~S���mJʏ(y ��M�w`g@˾�J��������2e)�uޣ{��懡�HsKl�1�����6�n���I�ٯ5��{ծ^j�w�<ma�݋)n{K�CЎe�°{�(�[����X�����@Ipf�Q��~~�������wf�;�d�+w1��Չ�ꥹӖW�u����l�m�)��B���U��A\^�y��\s�]��v�T�j�b��p���g�Yß[R�뫫�t_��r�{{�Ǳ�
���+�U0����î�-`��6M��.�
5�i �n�D�V:MY�3l��>
�&٬P�zܣ���N 5]:{�j�۝\n�U��X�"N��6��f_�x����g���b�g�-l�1sr�<Ձ�4=��ivo�þ�,�3��`�c� J̻�
���'�=�N���m9�}v���Ub���^W�2���Y
/g%���y�?�v��"q�q��E]��=j_�^����W|�^ƥ����?9BQ�5iaٴ�.^ʚ� ��(fک�Ek�'��G:��B��x7G,t�1���n	�%��N]��8I�kەd��u<=��z�ۙ�#�5K��ey��$L�Ȣ� xԣ����Y�P�ۙ||=)��͂E5g��\xd�c��\HQXo�kk�~����n�~���DV��0LJkY�z	�(
��d5�(�<�4���`���� �BLz뮝�� �uѻ�����пx2��򞵇j���܃WNs�{YT��������������s�p�j�%�grydk�ib�;�9�ÑhJ�QU%�ټS�FjhRk�WW}��N�yv�xxďJ�^�6(�x�C�b�֞���?{�Z-�X�[ޞ�~�E�(� >��8�z��r�^�@��ZxKa���9t$f�ZX�k�[
�T���c2���G�ʴh�3�ƦO��zS3����X����x�wu�O�����~�Z�1l>�~o4�b��I�$�nǐ�/�[^ e�X]��ne�9�����(ޤ�nA"�'8��T��.Hw���x%�eH��o���mqòx֚���tB�q|{�]W� p^�����	ɼ�񹵫k�`�(Oc�,1�g�\��2g��(�#�knZ�瑍x����X�n@<k��(4?�kӉ��q8΁�_���1�k5G�q�`�{��9v�@�c��k^c��͍9<���:�>�O�W�x�c��Ix��E\^��yu��}{�J8�[�W�cT��� �T�\:ڳ=o�ͅh�N�
b�w1_��ߣ�Ss[�IkQ�Ie9���=�>����� Gk�\���&TN�������	��˴Mmcj�fz��]��^h���"��z�ɕ]�+��FT
���+V�� q]�:�at^�,�=�t{Ն9Ll����ו�<����Zʌ�v�<� �C=�g
������o�K�ٗ��.�c�y5���³^Sm�
�>e�N�V����V��Hs�?T�����k̗[è┫ �c�ִmťV��Q�+z^'Z�)�d���n]�؇�|��'S'�3�k*�������7��sV�7��������N�A#,O[޺�cI�X}ɯ w��g+�-�n�ɢNu����!
�`�՛���G���DT~{�Ю�&���:�������X4x�Y㾂��@O�4�Z���~'��3<��V�T�����W��n���#��^��SS�kʙ[vD���;��Q���)	g�|���<���)GY��*l���ҵ=瀠A�:��u��)�儑I׆�U��O��M`�p�|ie�苓��d��3��^9�.�����;�ҋ}�O҈���"�X*XJ��[=s�+72{x{��0q�|ѭ�:�르��-�*�뽏ˑżD�=9G�ώ ^9�ɝ�����`�7=���;�i�_���(�K�;>U�żP���ux;�/c����ܪ�M��R�UEUR�qk �z����OY4��D�ah�J�T��0.X��^_;maF����f	�L5���R�I	J$�^�$H-QJ>7�*�/�k�Ok���W���4���!���%��KV�HcŤ��G��E�BA�IU���i[�v�[��{��K����R�)1bt��_�L��5kT���&~0�R����u&��
��q��9��� ������7d�[�$���`����@�O�1Qi.펟�XsFՎ���Ȟ�}1Y��sW�^:ߴ�1:��"J��ĉMG�G��;�Gj����3=j�t����
Fr�/ֺdb��՘�I�0�-n��Q�G::!�3��<�y�)���rR~�! �MM��5�Lt��Ɨ�V)L$$0:뾰L$�B���CLR���VgP�˘�}5f�Cv���6�H"n�)*UUIgG(p&<[�m&�{�F1kҥ}}֚&&��Q�n����,C�61{oxY��]���L�+7v�KI��KISZ��yH��ڏ����vL>�o2�e�\-"�d{{V�u�e��vJ�S����;M����_l������=�n�)	M�RQZ�}^d���ۊjj15R��a��u�E�-in��D��<�H"}�Ԟ�)�X��'*���8�0��KpI�Ȧ�1bF�!䌛� B&FC����(��/.��$��ԛ�VrDB%���i1L�$qt�I���F�+\*2��Ԗ<
�^D�^I�R��
K�Z��f1ŃT�U�Ձ����D�.y�NN�Ď�R��^N䟹I%'-�攟Gݵ>�k_�|X��ޜrG?9�M�,��y�E���O6ök�Q�Z%�#�F;cTa���HH"u9��8W �^(��A˿�F��D��%���e�V�w�}!���s��M��8	v�z{�֌��gK�=\��R�\�����1��}�6ё���j<UV�sU�4Ѭ��v��$/�֎�ev�}=1W7[�,U���YM��߲�:�,�j���LQ�=i�Gv��P���*I�/<�ǇiD����NO3�����u;��Rd�L���������q�����fz}!��X��;b��9�mD��g?���)���<�