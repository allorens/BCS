BZh91AY&SY����R_�pq���"� ����bB��          �򈯬��D�R(������DU����1�T�Mm�[4U%QR�bͦ�!��fIQi��ڵ�%��-��EV�LA�Y�rz��e+Y����*�F��&Ydl�2�i��6)RVٲ�T�Z�m�)�M��5�FƐ4+jj�i�6�F��l� �|�J�Lٱ�-�5��p	�kM��p�ƒ4ٖf�[mKYZV�*�mYY��b�R��k`4m�)��l�f������@�e.��zU�Zʩ�`�   �ݜ��Ӿ�^n���i�^���S���9�z������v��mo�%{�ݸq������ޫʝ;�����vEޚ����3�(:u�����*�Y�ȩfL�� ݼԂ�J�ݷ�����k7=(IRQ[�Ͻ�%R�TWޗ�Ҩ �}���(�*Wr\=�=�j�+�t�
�8�{�fJU�N���޴Ҕ�����`mbI��FT���� ���*�cJo�ۨ*� ����ﭟ;���}�΃B��>K�=(�4����}E*J�;���*�}a+>�|��{`��qo�|�*�J����}TP	+���6-kRv�+�T�]�  <�}褤�{������*�Q�S�z�JT�����P)B��[^��HU_i��=�>j�I�o����=5IQ���y�*R�J����J*�o{P
%^Ͼ9TC[FP��F EJ�V�  >����*�A��>�=�Ԓ�yϾ{�PY����}��R�Η��I^�E^q��}
�>�d�|��>��FO�����P$��������}HK�|w��-�⬋l�m��
��Vkj�   �JR��}۹�����r��������B�>�7��&��*ꬻIRVw��J��=���Ǫ�	Rx����*U%�q���"��m%*�J��Iěflce
la��0|  ��>�%R�yN�* >=�
�����Ǡ�C����U�SPx��=]�#��OWV��iy�Z;��;S��� {��MJ�L�V�j�I��T�|   g��Ҫ���y֩�޷�*G�FøU+�����g[ н�׷�B��7�QR;�^/
����Ԁ��x�k6�6��%+BTѓ�  O��I}�n��8Q�ν��zUޗ�ުu��p��Q٨0l	��=מ�AT,^l�ZǮ`=I[�U��4Ʃ����  u�馊]Î������*�x�]:нǽ���U��=�U
��z :l]���Үm�׶�y R�   
    j`�J�&�  ��4�����E@&LOI� �2d�b)���H �    5O�	IR�      jy *J�G��ѴL&��h QD=(�i�M��Oh��C&M��>���/�}����(W�|�W��De����d�b��[���s�o�~�W=�׷�*�
��AT�`���Q@hh'�������O�* 
��*�����
�=���2(
�����W�}'�2~�a�Md�Md�md�M`�Md�`�a�Mm`�5�Y5�X5�Xu�Y1��5�Xu�Y5�Y5�X5�fa�Md�Md�M`�a�\a�Ma�`�`��5�5�Y5�Y5�Y5�X1�d�M`�Md�Md�Md�md�5�Y5�Y5�Y5�X1��5�X5�X5�Y5�Y5�X��d�M`�M`�d�MbgX5�X5�Xu�X5�X5�md�M`�Md�Md�MeуY5�Xu�Y5�X5�Y5��d�d�d�a�`֙5�Y5�Y5�Xu�Y5�FMa�M`֙5�X5�Y5�Zd�d�Xu�Xi��XWT�@u�`GY�5�MdeY�dGX�u�`GY�Pu�cX�T�Pu�dYT�u�eY ��1�M`GX�@u�`X�5�e�& u�dSY�Tu�`XA�5�a	�eSYQ�5�MaYT�U5�ad`X�@u�MaXT�5�eSYe`Y�A5�dXT�5�MeSYCX`YT�U5�eCYA�U5�MdSYGYdX�@u�MaXA�5�MdGX�&� u�MaSYA�U5�MaY�Du�laGXQ�Tu�MaSXQ�Q5�`GX�aSX� u�dXT�@u�MdSXY�eSXT�U5�eSYQ�U5�`GYP�`Y�U5�]dXA� u�aSXf5�]aGX�Du�d �aq�e@�a � aGX�Au�5�	�]`@�@eYA�u�M�BeX�Du�aY�Du�]`cYXaSYQ�@u�]eGY�u�`\a`G�U5�]`X@5�dX �WX@5�]eYA�@u�`GXE���� u�aY�Pu�dGY�Eu�fA�Du�aGYA�Du�dGYE�Qu�Y�XA�u�]` �u�Ma�Md֘5�Y5�Y5�Xu�Xu�fa�Ma�Md�Md�M`��La�d�]d�d֙5�Xu�Y5�Xu�X&5�Z`�Ma�Md�Md�Ma�Mu�Xe�Xu�Y��M`�d�`�`�`�2��La�d�d�`�d�\Ld�d�d�Y5�\q5�5�Y5�Xu�Xu�\q5�5�X5�Y5�Y5�X1��5�Y5�Xu�Xu�X1�a�d�d�d�`�LcXq�Xd�MgX�5�X'\Md�Md�Md�d�Ma�m`�5�Y5�Y5�Y5�Y5�Xg\d�Md�`�d�i�a�M`5�Y5�Yu�p�y�������<fP�Ϗ�{c��\)?�~+p#�t�nJ��4`�!*���X�+�zDI��Ψ�a��nl��KdyB��	��W�i��:$� �": D(���mX�B�1�t��v'�H����=�Q�;��Sl�FY����,���1����k��N��076��u�ŭ�Yh�-e*�,��x���X�.��u֭�b�U	?[�iE�sA�*���.�)+�Zu�����)�4�D��sȴŰf��`���7�[ǭ�i,�^�ڂS>��Jb�����@:-��1���뱁��cI��E�K(�E��IpR�h���=��I���u���2�g8����7�U[0�Q�Q�L��B��5s&�8`c
ucr�v7r��E�SSI4�W���Ã�ƃ#��^�RُQ�l3B��v�*���)��ibNm�+Y��x�]�3%��� 5X0��a�Krf���A���2"T{J�	'�6�d]�-g���8��ѭ�KшZJaj��z���Ӎ,ڍ�$r��r��zE'�\��N7��㌴�M<�7)�Lo�
k�/,�f���P�K(fTt�f6VQQ;R����H��u
��k�h^���c�pPGzs0�9э`:K�;�R� 30��w�[H�k�qUBp:�2�av�fa=f٬�eI�#0�0���D�Y�r��驖f⣻�b�a�#k/p��sI�3+=F�Ȱ#�a�8�3B
�)��7��4����c��B�$s��U�����rxåTzZN���u.[L)������S��6-L�V����ׁq�OJup�s\�2�Z�̙��ds��.����K6v;�q�#�������l���� �)8]�lD{�YR���[��XDi��n�%�b�4Y�U���QB�̂hsW�X,�}Q⫲��=�����{�����eݬ�����1z��CZ1S*��$b�N���V�Vʪ�mf��1%
��9�t��0��K'L�w%C��7�*�u��*�7��Xo&��W�i���v���d��3"��ߦ0�<�Rn��IձsaՀ��u6���J�Ô� �ߖ�d/+˷Fm4i�tw��B���m�4�B�808��f��E��R�E���lT��V�8���$XH�uP,m�<i23J[>Z��x�j�c-�Ѷsp�F���m���F�:��(5�-����SZf-��+
���m��`|t�9Y�hV1x��]a�ձ��p:��N�[�؞j�Ԭz�wS6����tM���:plP�/x�ɧ��yu�7�VW��lp�ߡ��GC����#66�
�Ӈn���c4|w�X.�i�y��3*�G��
��K���Sd�ЩWwc]�:�|�V����V��T� �\z���h	�[�I�͛Y#uIj�Dv��9�z��Պ�.�c����mH�x��rRȞ���C�Ҫ&-�o$�֚h[�v-��@����K�+M,]��7�Ұ�c�|;j�חG!Y�O%�;T�HI�#�C�a����w�cT��k6<J��;ȡ�0�k-�3M@���#Kh����.���#�$遚"��!Xc�`F�U�-�&e8;�k`�����'F�,˼�Y'2�K�e�8� Ϛ�-��S�
-���6k+��x^al����v����׳V�b��,#+C2�Y�H�E4�q9����WR"�ʳcj�$�TI!�[��<_-���i�d6q���V7����wH�֞��;B���2����X��3�ww,"^{zZ����g ʮ��6�d
�R��Ю���^�R�PN�.��4;��ր)�Ţ{�:��=�E<�UrV�kd+f(����;*V��;2�6(9d�ۀa��^�a�&�j��/sG���H�K܉c�kp�$[M,���f�X#��?�	�ڳ���4��*\�Wi�e�i�oP���5Aje6M#D�f��+]5��������aAW1z�!{؎�v��AUٺ��;Y��RлU.ށwK@,%7L�X�����YX��R�堋�]
o(d�C���8���sݏ_Ԩ(��µ��R�O�FN��V�)f��1]IܣS��p�������Q�w� ��khQԖ!h:��:� �bT�Ӳi�1��
;�6o6���K��C�ü8�tV�HbӺ�_�x�-ߣ:��ѧ���N�Vj��3������	��D)q�c�m!'rA{2���
�q�ʰ^���ֆ��5���É�F�V+I�Z�$z��o/�{�R������z��.C�eo�W�3Lʁ��D3 :�q<��E^�BT<n�XNnٛ�Bm�=G�̑�H,�wW��̑D�ν��[Ý��R;���_g���.��kKY�����k.��K+8��!��9�p(*�cJPƓo5Ln���؇uѬ3P&T�t�]ǲ�-�w�.�3j���@��#V�/t��͌�FYSEɚ�|���;^XjS��n�\���!<r����/���\�qoʞN�*v�b���QV<ŋC��G)2�Ҁhz�������)��Su�@V��������M/6�M�E0Q��S���JS�t��p��gw��� ��l�*Ѵ�G���T)n��A��ßL����ð��N�zsѓRI7Y�̴F
���5�!�j���y�Ӡ�`fD$Q3^��Z3x�u�=;\�5MǅU��r�z��B�A�&f���ёn�h´�F\�o��śt��2�/B�nQ��������W1S�5���k��f�1uՈq��ŕ����ln���9-���e4���# ������v�%��n��od�h��i�Zc���㋍]����g��>���+4ۋ)#2�in;9tD�.��4�F���˨����fX<�>��$��a�6nY�!�>�ͧ��н)e�F�V.�Rݑ "��&�K�)L��2]�x�>��`0E	Z��DPA��-p���fŎ��͓qe��sy�Y�p��E��e��]/�w�qjr��l�բٺK#Vl�U����DwV u;��N��"LÑJ��M�H�/;0�j$=�DjU��`:�TEp������i����ţ��7�5�NJa�tj��P�jU��wW��K��	%	H(l;�e̒��k��9(�X���Rn~�K�w$��V�0XLѫE���*ǵ^(����7Gek�obIkoj[nh��E�6��g�Y��TQ��*��]:9l�i�������N�9��c���a���,�wS$�7	�Q�*��&cƉ��]�K1�i���B{.�Y�7��Z6h�֞�R�P��Lm5���X�ִ�SSY����I����Д�w��3;�{݊Me���n.v^$�;�W��P��	�䤰Y�Ռn���؅���X�w�M1͖>���K�L�*N�;6^{�-\�()���J�Jm	g1�nԨ�V<�8�{/Aa��E�8��K��^PJҚ��C$�Bq�f\��/�=�ɣN�\�A+����}5O�nl�х������2��u�5`��a���aƙ��>�#��q���h�\v>Ǵ�PY����¤�,t�*��^\�5�Cn�aI������I-<���ƥ�qK!�����+%=ző�K¶����V<$��K���+X��X�*��ҫU�����G2̹&kh��6�:��^:��Z�ɩVYP��ҩMn�1��6�,�i|$ikޛ#���p����xrU��c&��8���t� ��I�iw�_,�j�tz�+c`,&�u�*�!�!E�4�kSwM�k(�
�Ӱ�u�1�,��('v��⾇AG&��f��{{*u"�u����)�}���v��mp��T�{1�([w���re=u���L���1��W+o@��h�86F�@촦i.^��&��6���8���Y�]�YH<J�c�ݠ�]wJӳK��{�숸F�"r��.��wx�q���^;�oZC�{&{
piU3D�˗�0$�=�M{�k4�z��<Rw�۠XM]�����T�;��o�,����Q{Z2P4�[���z��6�p��@#�*Z�7�fV(m�q�7R5��ri�Z#� �-l�X���"�'n�7M��W6�Pظ��ޝ�3����S��bcj2�*e2�KN�Z�sj��̐�v�C���aɰ��r�Ôc��#�j����
���z�A/)ڇY�qm�{yM=�%4�� ۠mӬ�%���n��Z��׶	[��y�/pT�ѐ,�QwzJ9�ld�E��PcQA���F�:��+8H��w��}r��PO$Y�<g�?���[ܮ�D��T��՚*OF���Cr2�����S��}��԰��Wy���-��,��M�F�I�ӖP�&�3R�M\H6f�4�}f6��EE��2��
®�MA��
7�'m맩�����)�V������*�*̩j����
��.��ײF/�����|�`p����j�>�{u:xp3Z�(2`z�cSi'cDF&�y55Tum4nn�JkpZ������3/bSf��;��S��D�ǖ� I�;3J��q���&j��T�_enrb��t;p&�C����X[����d04V`
�����s3,w@�� ��3��a�6;�e�E1{�x�a!�+F�f��̦��N�
�tﺃ�WcV��-�X�P��r�l �N�	<j�Y�&\ׁ*�yT){�8o��x��侪�[��\3�ҭ���9�.�ia�ڙQ!A�^�7��m{�1T�@�V�u�ze�g�6U�܅�8U��ͳ���8��%X�(!z�e8�sp�L��,:�p�:5M�e�":�����R�U�-�z�7�F��2��t*[Č�db|,�!�e�C��F
x��u]G>e
�C��)���(;���]�
%-�Ғ�����|�[�&��{�S�wu���k�s���2ل5>�W-�Ym0£�TܵHH�!h�F��[@�Qdj�,w���4�^R�����X(,�w5�_Z�X���D
������4�^=/����8�o���dై$l��#m�+�5������5�	�\7���9}j��C�v����sY��a�m UL3�a��c���k��=
𗪝j��|�:U$�r��0��Z��+0f���4qj�1'��,2#F�9��µV��.RqZ��!H�ӂ�PV�"�u�"�d�OQ�D�g�]����B3���,tĉ�=�,���u��޾�:�io"����eo8\���K��k���dRc�VS�7^l �;v
E���;���s�8�.֡�@�%�l���=��,��ɇb�،0��%#W��ѥ�7n1@�r�m��-h�_ߞ�B�
խ��CjQ�e��Cَk�洡�{[v�HMz����"D���QS2=��Z0S���q Je{��]86٦�ĸ��"Γ���[�{y�0jU�Z�Obɍ�a���B� U<'sx���,�Ǡ�28�Zi�"�T��.��&fZjK���+���&X��� !������=��_S���Ig��%�M����*�h昻���k���� �k�B��
E�J�HO�N�3(�AH�#7�O~[5)�p�홮%���(�
Ɂ���@�H���*�����{g45X�cVc[�CX�Js��	�sF�w����Z�n����J��1/Tt��ە��I�� ��.�7f���x���T�U�i�.�ޗ[�-f�M���r�m�I�z�<BdO5��F֚
W��,�Ua*C�M�P�:J}��)��ͺuw$�ͫ�5tpfl�G��5�G����a�pTݸ)�7K&7�6�ێK2^C,�hڬ�/]��,���h �b��E���^ÓaH�4Mu�l�"�����]��ye�άP�7��Վ�&�Զ��!RrUԍC�ʔ����[���i���1�ش�e�M�d��飃fʙ�Zn��`���+��*��w^��ϋ�|��n�=�D��<tg����뵝�o8�q��P8UѺ J� T�Fčʹ�}6�SA��8�#�FQ��M��Om�1�t�7��k�6�^1�*!j�3H8#����e��Ueɾ]��'܃�և�Sݕ�+l�p6�.@��-S,Mw���D�>	"D��}FM6,uT�^���=�����JĻ�x�ɣ'`�urQ݊'�!R i(�� g��U%�Y}������[�sa�F��v��<X&�v�>�:��b��S��f��i5�QM2��aL�r��ޚ���f���m�S�7.Q�Fi̱tS.�|f�����ܶ+�\�cR&��Kp�%�4&࣬��h�P#8�-��IM��z ^l��u�ΰ9�\VRB���!�t,^�Z���;o/�J�hYÌ	��6.�^%������p��G�4Ҫ��7iMЖ���,X&@I��֫�o	��Gb�9��BX���$C�L�A)w!M@���(2�Q�4�_\����r)�v��A��N0P���Q�L죵w��E�H\�����/IZr���r�<�̅��yoVuL宅NrL��s���"��;[ߍ�R�e�KgRqz-9�nx��;�6��˕���ؗ�l9��+�nA>X����U�J��e�M��y���!b�|�҃����Ѥ-Q�E,R^^b+�;0bV�EZku��%ۙ���V�]*V�Ol��B4YQQ��FL=�n��#���ID�e���FV	�<nNs+�:��U���g���ܞ,�T�-w��ܶ��af�8#4�!��'?���Y3\�z$���<�I��[��[+�ƕ�)�q��m�I �Z0�F�-:��g��_���{����`�� �ރ���_0~ٍ���������$�;#�B�_[�mZ��C��������|���ε��环�d�RvS5O9�x�sc84q���rN��[��V�ò���uҎ��VM��8V�b�ء�6^��Ty��3�;��/K6�h`�>Mk�����������wԒ�J��c����߁��c-l�s
��gζ�
�,+؞ƅ"5>�� ��ΗnH�Xc��*�뀅wktZ<�R�+��%jÆ�	��ǲ�e
�}J;��9��H�k�UW��̊O����B:[\�[7/��[z�;4M�We��u��	X�֎t����B�GvU
#���z���NZ;��S�ۖ����z��,m�x�i�s��'����`��1�c��6��7���*0�4�&tT���>̬�}�fܒ��$��Υ �,-�Љ_&gm�<(�o��:��cde��;n�Èuvof9$�y^���-�U�d������Ew6��*"J�)�|�<��ꃐK�}���p��.�(�[�r΅/�oV�v�d��2�*�����b-�2�Y�j�F�����C�D�Rۃ��?ghYd�5��[�����5c��:Vo�0|���}��3���Տ�Ӎe0��![��/\���{���ff�Rc�ˍ�I�|0��f�t/�D;(��<�(!��g����(PJk=�Y�p��B!Z�o/"���n�
<�蔊�����~�Oi���OB�����`���-D7p�[sf(BY\a���2�3L���%$�f��z]+�c��D��h�����.t�wV5y�Ծ̩��R[���F)Nk)hyX<�����g>܁�P���:��ݗ��ƟIw8?xR	Fo���̦( �(�u���F.AtT�J]�!�Ѹ{8���r�e�mu�Z{�~� ����c`rHt���t_hK����$&v��u�y	���EkU���� W%� e�d��ޮ�UÎ^w��S�7M�^�U[�m�֝ٙ%:�B����H�A�x�o>�,�%�$3t��Z�����!v;����tF��`���A#�<�D��|g��KM��\��k:�q\��M2)��tC)�u�޳|�<Y#$ $$ŹG��	K�w�n��6���6��n�>t�Ȱ��:�N�c����CQ
��m�LA��!(8���9y�� �^���J���R��;gl�\^�A���qkF�A���CV̮@�G M���r���=LN����p�h]P�����7�\�]�6L��jܺ�P��=VQ�ːT,��gD���҅�z�4�H��k���kB��k3I|����[���*�sY�U{���z�\KFc�viH����@V����-�o���z��J��t��궯2�>B��fR*�m���6��/�?o8�&�۹�]>�YYI�w�9�g�K"(�;,q���	��c�(_-iTK��˲�j�v����8Yý� <;1<�Ƶ-��ʷ+�oe�����Bvh�����t���V��jKcu�`�S�`[��֧عB�l���Y)��M�����;jU�������݇���^�6Bs#7�3�]k�����.D�[s���y7����v���u �d�F�!��*�f�}�d���`�:�;W����'ұ�b��h�3z�G����Y���
-�>Rw`�Wk�S���m0�D��\K��쫢W���f#���X����hr�Y�;�n��Y�
{8ÂU˽͔��5ǡ�{>+��;P޴C�����f�mc�qhŒ�/8W���8�R��E' ��e��f7Ω�c�����q�"ƕ�9L7�m۬�$�H�D�X���i��q^�gFU�!�f��ݾ�7U��T[���av�[�MN)f0_ǡ��8�sa�ӏ�ԡ����MF��h�8�Y3�&�{м���k�o��sY�U#;F:ݽ�j����a�%u24ب!�)�p�;J��X�H��S��,��!�\��'\�t��\�����4t4��X��.L�9�rt{akK���Utb��T�����t��ő���c��Y����SM�L#L���7�V�0�WQ�0��[�i�
�͆�6��Ed�ޮEZ�l�ë�7��ѕ%��T�p3^2��t)�wr����ȮtX������uh����uI�S]�v��:�=ᒓo�T�u�i`���#
��:������ז��:L��ⴾ��Z���z����%Z�L�ۊ��CI��:���1h��X�%�u{�2:��5!�.���oi���lmD�H{f{�Θ�w��݌:Rd�"e�L�U4�9m�5������j����&v�;+�f�syZ3��\�0�o�o�v�]14�^u�F�F�F�e뭸����J��e���%v��ˈdv�
�^Q���`��WxL)�����#tbB��Ɏu�u���E8��^��%��Ƶ��>:K�m�M'D�uQ<!�}��vF�粕�m��d8v�\��������e���u�^�7���-�j3Wll$�;;�����Q��8���pL<q�tvd,���uړ���ٸ��n'#q5���S����jw{A>�/DN;�A�[}j��������ݢ��h?kL�O8*(v����{��ܺ�� �E�߶��\��t7Q��3�w�S<4Λ���hX�>�VkU��ѱ���"�l�����\��4#��vum��$�6�[;5��]t�F�]�E�K�E���Y��/�0x�U���t����;1�:5���hWl�C;���ƥ�9/3hd����=gc�U�5�%mm]S����)�j?7W��F�.7�r����y�b�U�d۱�i��[U�_�s�~��\�^��w}+j�MS��rev�k���9Y:�sg%��VA�q�Zk�ա�:�3��_w���YM÷OK��(�K}���)D͔&@��ٖ�����p�v;�}����P}^Oz�����&;�rB��IWw���f�`�5��<�(\�Ë�la{�,3�~kT��.�ژ�Ŵ��nB��3*��c\6��D�U�u��J�bv��5�w���#�&�ȎssbN�w�'��3���I/2N�Y���q�LRƴ8ġP]f�^M*����rA���O=��P��:�=��Zֻ[;���\pa9��ZrХ���s�xPoZ����+�oC/x�����V\��Ȗ�k��T��8z��5�ӏrm\��CJZVt�9�
�t��t�Vh�=.�a.[R �BH#jWu�дZ�`��+4RN�z�=XN�ώ��j��"x��|�'�!��KrS}p8"Y+lSnzk�,oqɚ
�Y��r[KP��\�eLn��bz{Y��l�����]�	�YA]�B�w�9w|�Ǉ�s����č��r����;��&�)�X��*GΈ��]dER] �q����2/-�eO	��Z4��wi�����+���P��mp}�J1��EY��&�r���#(֩�1�J��@ �f�;3�\9�䳨c���\t����zы]%ZJ��[��1մ�!���'eA�Ww}5���n�"E�ͨ{���q����R����Aβ������f��/`ٺ5��k-�ɃE-��iuћD��RH�m��۴ɻ�����ڗZ+�<�'N��hϵv.�s[3�^gI�&ٚ�A93ᢍKt�W|Q���n�ujm�O���.�����&fu�Cs�!��M=G�Qn���aaR�ZJ¼�h�Ge)�v��
�L�k�g4U����s�b��Q���Q'�s"�����8�(��@u�#�נuCR_Oe��������'ܫpS��;x��0y�0E����KeNs`}=<bgo�1��xhs<L�}�`���3f��PiXo��
��N���vX��e��*"�Mz=��9e�_��1y�k����ʺSޣ|������	m���dA�"�l��c�9���e�� .R��n��T�znh�0R=Rl��CD��Ӯ�}-Y��M ��%F%��?r�޷�S�OV�ŧ�㽏h��]��A$s7=�|���<��槟���D�R���ui%�i��f��$Yd�i��o-e��(r�J�5tm��5L�6գ��$EVޕ���i[���"�%���57sk�۬��#.�@��	��ѭ�5g�r��E:T���3+k����$���oTNC.�ff�',2���0�5�9W\�r�!�(mq�e�2�)Z�b��+*u�e�H��{�AV������b5����i91���2G��G���؂����9���[�M�?�H�Ν*�ƅ����g@�Sx�&f�z�Xr��z�jn:� >���3!9��Z47��#%_ĺӺ��ת�V�M==b=��s���`�}УX(�s�a�����jr�Oi�❩:��R�]���|nL��My0�`��=J�{�����
/�;����}%e��R��
vo����B�U�F�̔�v�fQ��\^7��i�T�{r+�&�����F���a�Toy��V�B�z��ǜj�����Xd��}IǯA�C�8������IT��3�#���ڨ4uq)��7�ө78�Ry�T�]%��[-0�\�R7�z�aނ���M�w.f���+X��J�Cfk���YD�d;���W-�>�XԆ閞vN��&XGH̆]+-Nki=mk5���ySE�� ��"�ِ>-Ͷ#�M���t�����mr��J�;{�Od\�M�T��8�y6��S4=MQ6��w��SML�'�.�D��8�m�J�}��w/y���*����&ȟ	��і5h�z�&p����-������ݎ��q��Ip��+N����֨7�Mֻ'Z(�8�M�A�X���"q��0��!�0����{&�!8s�9׺�|�r���BܵK+E��3�dZ�m`��r�{�Y[�7�Rw���y�Uh�_����*V��W��Y���4��Uҟ���S�cXG70�Wv�&�x��'/�Mx���m�x��4�0M�=<ʐ��)�)��Hų�6R���:%���-j�r�f:�S\d洺|���<|�
��}�����@z윻�s��}�m�]�,�'X����=��w�>g�:�eٔ����:�Ϣ�ӭ�^�J�3{�B�S��yQۢ&Q������Cy��ޥ ǪL��E;Ĵ��e�>i�Y��uF���c�/{V]}�(1T�tl��_U�;b7����a�'&VK4����KiA�k@ON���p�]�����e�|]�7g\�p��V7����U61��v����YQSh��x�5���t�L,�E�!(_�zw\����<�醖�ڛ����W��J�8�ɜvt��h�W��G��礷/�����<LGr������W�~A��4�X|]�˞����"b"�[jk��EΙ�})�	[���+=�F�#�5S���c[ow^J2�<kn=oc��F:�j	� Kv��ەӉ[e^i�Zɸ`w/��u��T�M��]�=�[жy����i���=�����o��o��n�Ҋ�o���+ÃO�2f���Yc�)�s�AZ%��(�4A̹����MvQ��|	� r����ig�M��q��"�A���}�R�����	�Tu7^��I�H��)ε8B!�� ��0�}��Wc_:����)������Lue�Չdۆi=�[�s��3&�t���$S�1x�S����q�5�\�2mA�yP�ȯ"}����)=�$�[�-Ja���Xՙ]kk7�=�!mjWG�����]�)3�7'y��z�O$�Μ_e�]p5��������$�̖goE;:��u��wÃZ%v�9��A�ݛ�Y|�hL��Q�g&��`������ʘ"�9�Xo��r�t�0��:Fq�j�1��ٚ��6������z
2Q��8iN��۱�(����Zu��췙l�����݅��.�R��8��=7]���ƺne�Z'��ܘ�^�Z���<�u��l��HG��U�ƩnPή`ɮJ�m�G������u�%ıl��'��I�.{�ΝaX
"D|ņ�ܩ����Q�am+[M�1�,� 0�e�/�0�P���	0�����
>Q�V�	f����b`�bEG0�A	��?�`��͆�Ԓ� �R(�ʋ��1�J��H��R�,c�� �J�MB)h�l���N����)�8Z"�C�K)�	�(��
a�Ad��5��E�"���I��eT�Q0R�m�"�t�k92X���g'�2.H2+d$k�$d��u(䨅
u7$hI�Q��I��Zֈ��-��y�c4�BQ��u�1�f�eH����:�+�8I�"�%:ܿ2h�P���ITLi�ߚ����$�P�(��(W� H)���c�26R��1K��V��P5��}�<�K�m��m��!0�,G �2ff,I��H�I���I|����G�tuI"���NUҕ(�Q�٦KN� $�,uQ�a"�_9���	װAP14n��U%T��v��a��t�Xa8�a��]%�^0�R	d5"R.O����LdY�_�"
?��?���@D?��Ͻ����" �G�a��??������˺���CU���u㽊Z�ss7iiW�E�wA
��5m�yM�t�@�1�A�6D�P�x�����X�S�8���\d�{��)P�۰jl_l�\�=���d1�]��)�Gd�.�L�e� ���YW�C\�܂oe_1�� ��gv�
���^ݞb]�}�GV��j�%v/�*�.��y�.~��o��.�����4*�����\bq�r4�.��87��7�ī��Z�Ҧ�yIgz�d/�3�W֮w��G����bW4«;��,dt�%R�{]t�p�+Ga;���M,_R����o�}_m�Y!���j��N�s��7M988�9�/ɲ�5ϖ�+u�ΦXr�2]��f��Xx^�JF>�k�2�woRC6��M
!Z����Y�;���ܓ�Z�ۖ���H�J�tZ�qQY�.S��|�-�;4+���^$�U��o�b�f�TY���y0�<�{��K$��&��;{��]�nZ�s�wp�ݨ�aL�ŕҮ�=C��Dֽ�jES�k�0�ݼ5ep)yAt�u��e���2��ʯ�t�|T/W�+A秷��T��.�}��u�\=nd�1�U�'�B���m�c�U���5�ˀ��U�bTz�VL$���`1���߷������x���Ǐ�<x���Ǐ:��Ǐ>�<x�׏<x�����<x��Ǐ�<x�㮺�Ǐ<~<g�<x����ǎ<x��ǏO<u�Ǐ<x�x��<x���Ǐ=<x�Ǐ<x����x��Ǐ<~<g�<x����ǎ�x�Ǐ�<~>ޟ�������x��Ƿ�<u�Ǐ<}<zzq��ǟO�����}>_O���fc�y��T����6�p�o,4j���g�I����&�;`г���bȝ^��L]8��2�qD�ǔ3k��vhr*F��������O��c���̖8�x�.�������Å�5�%���X�nv,�$Ԝ��K$go�Oh^���O#:���m��#��du���8c����$��]5�٠ �N��}�F�l��4�L��M��k�ӍbMd3��ʀ��9æ�vFXS8�ˠ���Om�\�����He6%�Q�h���f�y����[�5�ڇ��NtĎ3���<*2�P���N'XТfG-Pb���Տ+��Տ^�ts	���K3N�n�f�fD>HS�:�V��+m��{r��ժ�1�6�>�8_h�|A1�/(0em\����Ct)��}f�����>�͏E����`V.�EA �S4�!�͟r��B��g~6�b�:��:�
���A�F��+��9�a���鷜�ğ^�oHJK�m|�,R��tLs�ޕB���6U���z�-����*y�̵1�]�ٝ��a�;�_^r�6��A�u�6���T��섛kW)����Ӂȏ!'Ss]A8����ȱ��_/���Q�D}X)��}I��MK��S���3�;J��]�F,+�Cﾩ���/�����_O����g�<x����ǎ<x��ǏO<u�Ǐ<x�x��<x���Ǐ=<x�㮺�<x�����x��Ǐ<~<<x��Ǐ<x<x��Ǐ<x�x��Ǐ<}�x�Ǐ<zx��Ǐo���Ǐ<x�x�<x��Ǐ��<x�����g����~?<}�x�Ǐ<x�����^=OOOCǏ<xϧ����,��$�1�b�@�f>s+>R�vf��^���o#�s��s�)B���t�9�x�;sC��*���am�cr�/��������y�uk����{�Q�s�$x.��8�żF�"=`���������}�z��J :e	Nn�t���Ab[νu�y[�{K�tLṸ&�lg�L�����x-��l�WYhVE^�$�k��ɳ�xc�;&��J�c�p�8 �'N�}s���{п����$�226�f諯��(��aX�����J�R��� .w;�[�JfV7�=B�6�2��)�&6�N�%�K��@�,��p_>C`��Ք!��i�]�m���ʛͬ儼kM�Z;]�v2�����6<��*�4���<a�u���]�D4i�3�;/k�0�}nKo
Jȫݽٴ�7�NE[�D��>���������	�&�=\�81�u��ԕnS�hF��A��8f�ydՇ����%r�|a�rwc:R�c��]�8���VPM��P<h�t�eT��+*D7����v�UWD,��b)Guj���VB�3.*K���=Zz�U�:w�Xo]bk���]�����5`�)��E�|��(��Qc�3AA`Yĺ�,�Ǯ�����oO������ǌ��Ǐ<zx�x<x���Ǐ<x<x��Ǐ<x�x��Ǐ<x�x�<x뮺���Ǐ=<x��ǧ�<x���ǎ�x��Ǐ��<u�Ǐ<}<x�Ǐ<x������Ǐx�������<{x��ǧ�<u�Ǐ<}<x�Ǐ<x�}?��~?�Ǐ?<x��Ǐ<�����<x���Ǐ<{x޻�s
��bww��2���qjǗ�L��R�y�W���K�֋	1wy+�n��f�N��l �Z���#�K�yZY��NP�#V�c׽϶���ʭȇ "�G�]����a����ڳp'���T��z����*���O2��9�wa���Z�Ă9F��k5kR©`�B��'mDҐZ���ׂ��; V�@�-Z,�'I�앹ՋbΤ�R�JfP��0�A1�D΋�tz;�'��Y������8v�]EV*(58,�U��N�Y�Ӥ�٭1�%��_$��xf��253Fenw�E���{�^^���ñ�`���i��J��/m;[����(�;��}��j�LcZ>G���3���,�3Mv�b��@�2�XQCg6��{oM��x/M�=,ޥ}V��H�bKx^��N�8�Tza��z�v���y���k_V����=_N�)����	 ʤrk��;/Z�����Е|f����v[��f�1w5�
�Dk�1M���jf��'�B����=}�K�`��;z��N���l6�ztB�R��#�w��D>�:�MKݥ{b��wSD���$WI����" ������.��4�q������W7��`F��Ӧ��	#�Ul�L��"ɾ�ť��\���y��i��|��,�&TY��W�g=�K��]�>�wKo`�[C����EraVh�+^eگ��]86*<5�܏�OR�2,uS�˼�c���2�<�ʝ�Z�U=���x_5�\n���;�W�B�l�ҭ�"�o�#8)��T�cU�E�%�=첝��R����,US��ok2�J=�m�"�t��{�}�8��>������q[[Jf�#�ȸ��}T�v�w��:c���BW.
��b*o�>����9���.�h�r�Z��/m+�����[ȩ�'3ö=N��� ۫��Mc}DLk�zuF��$�s�6���UJ�����5Z���a���ˢ(z�D{~�G��M���1�ގ�s���Dwօ�-$d�V9d�;�%}���E��Ä= '쾕�P�pi[���GS��2�#��1��)�"�?;�j\}G�\^q"�|+�'1[S:�����_\���m����u�^�H�YA4���_\ڴ`����V�Z�p��W�fe=w��T�q�.iӘ{	�0���+O�T��!��4Mr ��ܨA��<a׻����k��v#�~�.}�U�}���t�	�6(i��+u_tN�1gr���fs��CyZ~_ :�o�h���"��7("��I$����k�e[y϶� 4�`��®k��7����Z%+�I���Gü��?e��3瞝v����=�~}�@f㲒�y�K��*�����g[G�)����+���)}_1ɺq���T�Z�g�K�����h����qƳ���I�nӔ�WMp��:­�4E�DԔ.=�#柛��(������n�k�1�X;_R�N=��.�em\�R������|�yQ= ��D([q^`W94��x���ZaV�&@�9�/5��Ud�`\N��8�'��>�쾐҃�c�3��I�Ӎ&^uQ�cFq���l|A���#F��/c��g���-���?�υnh��*�<O���U�$��:w�*qK�y�����[[�9u0ਪ�L�Q_L��oo�5ʑz��2�S3y�6`�����`I�N�"&^c�_8Ж�o%J���,����A�#���ԟ�d�i?u~DJ���>c9����A8=���ⴜU(`��ݒj�
E6�T�tq@e��aE9�;��_kN����n�*����m��Xݞ���tϾ��P��
���ϫ��*6�
=]V&Ե���lΔђ��z"��&�v� ��PP
I�|#��R�k�����3����7�[8ӫa�u�53.�:1��R\\����]f;y:=Y6�=T4i%�_�K�r�7�6ni|��{[�A��㥙�l�ʖ!S*�ś���ij�!�x�)�9H���q��t�κɖ����!��A���e��ՀkF�����Κ9��䧙D�W]Cm�uK��B��S�mfa���k��:ӆ�_^�tҩ�H]ֽZ�yÌ��;o�{0(:aܮ0L�UB��!�����v�K��z�2����*��ґ�@$g;$�H����ܤ�爮�I-WQW��h�����5s)������/cbƳ�����w{w��y�v¾P	�>�&��6�:��Vܗ5S̽��1j�l����wNvE�Ω���ДBe|k�]�6RP�k_e���k\�r�n��P:��V%�i�k���H�^̑+��zvj�jq�K*Q�!=���O5�}!��agJ~o޸�X1-
�ei���0G�̮����*TU�e_i���"Jv� �6���B�#�Į��.ٰ�V�ܔ7�#���J/Y�[����H��z�/.{��"Cb�ͮ&�cY�&
�8$S���p��Lg���Y���<�h�q���7JR&v`�����GPw\�:��i�fZ笢�lx�Y��+�~
�'x�;6��\O�{�[�1�E��������,ȺS�w�;*���U�V�9����RQ�v�n��+���%4�)[F���H�8���_\V(,k��ݧ�#�9��}g*"O&ƞY��`���G	���'B��-�Q�oS{������)�5�,��|e�^Uʨ�J!�vnRH�pՖ�0,R�����[N��i�B�n" ����[|�a��`=fA�l�"���/-�T�S�Ј@#�G/:����:�/m'�Ӓ���E<�"8����΋.1�ێ!zԢ��s��Z�J�+/j���ו�҅R�խ�ͤ��B�t���͎P���{c�d�
nw7)�YM�"-F�)��u���&��GY�:����]0v�"�WU�>�b�]������#z8¥wN�G-�)�4n�fh_Wǉ�,Ǟ���&�Wzu�\��x�4T���Cʇ�7�����{��<}B���9���4��zP9��]�A���냻��/�s����(���OY��6��^8��m)x#�6��9���(x����n��IП$�a���r����L�ײ
z�Hj���U��c����6��wxqЭ�&���`b'���r�7�#���-��n�%Z���Gon�ۣ��W( 7�]���b�lNB��޽�%`��)�rٔU[�FPDg����\�8$&�qn��E�uv��������VHZ�
�Z�7@�P0�c�rFv�Ė��[%g�I�s�{x���,���E�Cך���of���)����{�_)/��k��t��D�<V�V�Fq�7��d\a#����_:ݣ۝a��7��7ԷJ�n��Ţi��<�:&�'AdM�uG�zq}-�SSy�Y7��]���Skn���e��=�[]���sE�.�6pr德;ܫD9)�U����x�j�,�F�cj�_%|2�bKp�w�s� ������4,��8�N��{�7\B!�3=���3��"!��0+���ON�����;�M���"|�ª���~����l���]��فn��!3��c�'ς0��1['V���tt����a���n�#�\��;��6��j>f�v
<2�W7.���6x�u��&�o�RYӻi�p�6���ެW2����+G[���5�Bڡ�>'����-���Pl�T�Kv3�2�N�)j�G*��gUs`m��w:� ��8��+W|�R�*Mc�Xm���uvΥ��Hd�w!{�;�?z�_��.:�Dq4頻d0_f�y�	ڈ�;�~�d��[<چŞ��g��
=�7�������1�%Trl�Y����]q����Ir�j?W��R�}�X���v:�ͳ��R�l�Y�V6�u�r����!z���:;��3en�)����Ԯ��!��]�i}���B=���ڜ�꦳6p��_à��S��[ųl%��v�<�-�:�c����5K��U٥eG,�LTK4��|�f�XJ����\zI��0m�;m��V_k��:Q�2�v�����ߺN�-fe%��u�Q�N��v(��}�l$�R�3����h�V��HG&ib���7\�`4iq`�m�褔G��qVP�q@(�4���ݛ�QHe����H�]NolK(�+����o��r�j䒏R�q�;��;��sZ�n�����je&���-�'َ�4���J}���+a��S�Y5c��J�A�e�}��K�mA`n�<���X�VQ[7�1�Z8b˂�<c[Ƕ���i�I��J�lq2�\Pt��R�:��*eK���Vt4�Q�
�X3w�*h����mv�#C����t�}ȏ3�=���6.�0�qowP/�RF��Of��B������r`�2�Do9j��͸�mq��4yd��xxBf�˫��ѢӲX�õh<ͼ�f�#I�Ş��%��ֹ}ưv����������*ۭin�VA��fjWm5sY�׍�3K}����˧��u��)�dD������@$�^�婳�}�~��(�*�aW���~�����%�������~_���F6�H�J�R�����*e��5�$o�&!M��0����{C0�$H�4��rw�Y!���a�"��zXґO��Su��46��}�Y�uЧ8P�R�	q��l��WG����ɻz�Ц�9��F>��
��-�<�ݫq�5�n�	&�*�n�j�ՆT�)����oI]X��Nv�9�"Vn�]��3X�@�(V�u,��v]�x/-M��<C�q+��1+x�f��0C�^�G<��F�7w/r|�l�Qq��Q&��ۣ����bR���h�%t�F�G����62�#�)��w����k��.*�*m�˳%��õ��MS�HÎa�g�m��m�ϧ���>7;۾cn5w5%)�:�[A�gmB+e�����26˽�^��]k��IGa��u��$���%�N�Q��N��@`\6�H���멭��)SU;y9����l*�Z�b�jT*��q௓5��bΕ�%��֔�*QPeNʲ��Ww��HZ����ꆎeF�����e�^��ǅjs�U�*`�}H�0��rM��כt����!���$ʒ$ŵ��ɒ�PSg%��R��/u��M�ݹ}͕�.�.àh���3:��u��S��&:G���!�I�#ǐ7q��V��g�c�ĳ��8Ca��J��蜱!%̙,J	-��28 .	������h1�R�0�a�R�N#b`1�1�,B�L(@�2����ҠD�-��1b�"η7"��3*�aHQAM/�2��"2	
�"��,�33$̌L��u��������?<fp~�~@f@َUc@dP�9�	HfaHdd����]x�����������p~?*���j ��@SM--IOpdRQ-C�q�^<{{{zzx��Ǐ�3�L��	E�W!
�;̜�!�h�(�1�5�q茊� �����w2�#��Iw,C&���l��
(���"��̀&��(,���R��31(�!sq�]`,2G
`��H&�2Gp�0�T�+3,(J��3r���Bkpq3��1
�ks2��Ơ�31#lv�cbH71 ��,�2��ٙ���Ĉ�"v�	�#�	()��(�ʋ���g`�+b��"�\���2M�%31l���7 ��20�W#!�\�:�ʚ����i����Z��rj��J

�%�{��4��$�j��ܙ>�!���reE�6aF�B�.J�-%�>yK����������M�}��-6�C���++v&������=��3>�����[Y����?HK3�:����-����i�W���zp}�T��[��䀘U}�p&��c�|o��߷�P|�	��\RW�d\z�U�>�9=^*�o��9���� ���ԟ�w�#�7j?Wy�;�~ց��u�㝷���O��'{��+�٣��}�~מ},&s*����a�&��y\Í��VYȪn�����/�ڙѵ�,g�:z"��l���U9�eW �>�v��f��z* � ����[8���[��־^�ב���>�U�;CH�vW�4ұ�^��0X��vY�*�>]�z=����q���ǉ���y���x�CV|�J�/��y.��b�S�f�RHU��9oEde���<='��;�?[���8�����Cf���	)H��Ub^�.Ɏn]R�}4w����o���8���.tQr4�3ʸկ:C��I�kĭ�b���{��1��`}\��>]ؑ��`i7�Xn�]��O���ŢXټ�NY���8��_;�0�ԇ�V�x���]�/�-�1���P��{�o3��]ܨ�i�%��6����(�?Z�O����&�������f�<ϤF��U|3RU��*в��Yߕ��~���l�j�(d��17��a�G�ZM%J?M�m�/��R��砢He���Ӈ<n���62ĉݷ��d'z�!9�+wR�������#���<�)�*�q�t) W�һ��{���sߧ����IW������{�U3&UH:���2���a?���~�ɿw�ɻ�x����ȫ⧦}+���k�*������;��w�nT������k�:��~eq�����¿���r�w�dU��P�=����3�<w܋�Gw�*�+����o�H���4#x��Ӛ�Dp�y�E�=:7C�p���=�&��n����6�E�Y#�(O��g��F�ƀ$ʼ͂�7&��V�k�Dƶ��׎߆t�n�M�ݳ�Ν�3�C��Dq�n��M�����KW��>��/J^ϵ�����AR�3�H�L��rw��J+/Ʈ���\5�[:1{:m�ygGw6�:l�4i����h�6� ΧjpGE�R66�[|@4�}����#XxY[ҭm�Y�].� �5��κ��)ss3�J̒B��)��TY���.NSs&J˿�Q�
���f����%�g���ۖ��,�_�����Ngt��6�޼c ��,a����=������Z��/�>���k�9'����k�����w��M�ӻ=�����+��ᾤ���?��޿��fj_���s]+;��J�-�ꑀ�Pᾪ>-�\�+臜Wo�k1��[k�ܘ{PyY �#�c�{���UdU�ͩ��*v��H�膿�u�H�%{�㳶���2��:;���}�G��2�+�u.�&*�W-��Q���Lw~����]��WANL)z)�g����A|6�H._m[%]I=�w�X�CS8��^�,��rm�C�0��^�����V�=n��l�y�
�y���|vP`��\LZo_�����u8��&-�)R,٭9��u�(ֹ���z�*��Q��btޚ}u��R̍ߪzA�k�<+�tN�:�=s��3nzJ�L��֟a�������⦫I�?~�ه�?�u6�
�P���l1�>E��͟���7�?��i�č�=��y��[D��T-,|�����ח�o7SDW"y�@��`��Q'Yt�$;z��{7��iz�%���[��tOg}�ӕ��&#�����>�}^�@��`������/�39^�s'-������	��4��k�R��{9���
�f`�NӮŅ��7Vd���t{�,ӗ�;-s������x7�G����o�v|�>�s8�l�z��n�v��ء⳪�qei������-S��}R���S�u�}\Tt�}u�u�p	�nm�G�@}��y���=ox'nEף�Ϧxn��R�lc��z�2Օ7��r<�K��N���p�=�Y�2<���}���y:N4�_�߽�2�����~W��@��oϻ j���w��c�0��g�OJ�1�^��k�?j�L��oJ|)LX������5c�;�������������,I�����2"32_�#:1Ov�q��\�q�{�d��s����\��8)��ga���範�g�4TM=�TX78|s���u�ܠ͸��a�:sÍ0����I ��ᡘ3���6�M�t�>+�������y���݌
T^h���~�C��-M����/����P<�J[��}fiO�lhnjh2Ht/�$��)M�Sr=��2��f��M���Ј�xR��Z��ܓ/����s�߼���3�l��$���oA�F7��ї�"��f��鼮�`N�bh�;Iۨ3������ݐެ�.1�ٶ+dP�Kb���jMÞѕ���+�΄�=Q�>��dg��`0��!���1�*��)���%�n��6��x��ռ�V�#oQ�=-��Y�j���%��*�^k�5���)x�R�'y�Y�^3�=�T���r��ϰvk��OIÚ����N�Z�g��*���g���}/���f�x��sdw��=�����r�&C����� ��Ϸ��k3�ټ�:��m�*�LU������O/�<�+ ���o�����Wy��B���C�����|!��qIۦvv=�C�6�o������Y^蜼u��Q=~@+�n��.�Ѐ1'X���L6k6Ԙ�hf�$�`�of�x.��V���R�wWR���.�y@��Y�Mw����Y�F�=�2l�V��j�v�ű�b�KM��Q^vȻDn������@��<r���ɭ(V#����7����TG���6��ψ?�Y��<��0�p`¼�����l��}ׄ�B^z�I�/w��ߧ.��V�+}69�Z�=;hzOA漵J�f�u�)�&`dຩ����ph;��y�����L�ޑ]�d�rÞr��y���lw=^���8e!`��6�e�oʎ=ޛ;n�xI���o�P��ݛJ��MߖW���O����~�9T^42n�ْ� F�'���U�'_��WM���U���q��/�NF�;,N	GwPO,�u>p}:|�'ݝ��ɫ5�yt�Ϗ�D�:���y�vg�x��Fu��~���ޜ�B��J�&���S���=�ѕF`�;�uM!!��^�)A�7�S��K���z����vy]���[��K~[�:��#��S�ʵ�/&��u�{Ɩ��秩�L��Ӵ8/λ�t��D�^$�B�(��E�����	�8�ӏ"r�����_ɼE��X����c��� 1;iv�@���ؐ։��^�E�5`��b��Z���jQ:S��Ӥ��R�V��,�}�gY]�U�-�^�!�秐���m�}`��q����w�C���|A��͡k�����s��~^�퓱l��-��ρ��ʶ������M�yh])j7�������_�Fl����{/�wU�R9\�� �3xf+�R��|��:~�S�v�HV�{8��6���&�^���0��=v�=�!哥�{�`����J�nh�we���_QY)�A���q�y.�z<�}�z��{�W�Γ����F�t��Ĺ��9��hzy�oٺV��C
�cJV����u/�};�t��u�"�V[˿9e���i�$]DY��Em�_^Λ<v��� .�s���P'i���٫p��bJ�f��lk�sfM�y�m�{�|�V*��D5�>MW�B�)i {Ɨ���۳9(�w}�ܤ�w=����
��N>ϫc-uI�&t��/Q���J�k>"��s��f�~�����(�@w ׹��4ț�#��CI��
�~���"��O�Jhu��f�K���k���� >�K'6,��W9 rҞ�w%]r�f�u�Z���tB*˴^t@�,�Vg�ظ��et/w��_[���ES�W�P�'-E��ɗO�Ws��+��-�f�8�S�����r�[��4���|ӂ`��ƙ����n��O]/�i7�/��1��Onߔ��im��c�Ȏ QnS����Ю�>?�I�R��_�yZn���	ݦ�hH�.'���mG(�Wz��a|�/������o�9O���=����G���썍��Ѧt�|N�4d鋑����G���z���VM���ﾍ?L5����Q� G����+��������^�cM�e\�/��I�{�3��M�ׂ3v*2|k\��v���������v��Ĺ����"�咭��j��S�Fp>�y�ɼ�{��\�YZ���%]���4�rt4�V|��}*S�'�^�5-���/'�G-���7�v��2o;�?Vlz�_���/���mnܻWWz�7Y��\�*Uj�h9W�K:x��JҢ���U\��%u���"�S��eDw��#�f1��T�<s;����'�y%RRC$%T��l^,��бR^�o�S�n<	��#7,,��+�7J����ٷd>ހ������_nVC�fPHA�a!��i�M�,�����k5I�M{�<N�-�_�"BA����~��	I��g�W�<�>y~p��~�cm�L6�f���;5���Gh���ݱtt�yMǜUy��<�Z�ᇼ��vNގ�=&f	��ly���֒}ۢx�No�K��I�9զ��v��[C�ߗ��v���AJ�ԏ�ˣ�����41^k=ٙ�8WDQ�pH�h�;��6X�5{��F�j��������[��J*߳[��{�_�oA�Y��Q󮌿�������W���=s�W�jmO�fgz���yfgW���{"7_֏����/�߇B}���v�C}��%�~�~��][ ��K�Y�vT�~����i�!yV:'X�o�u��I���{��#����~�O,97�����{<��ޑ�.�&�7=Sz�R�}b��Q�r�4
�w���Ʀ��I�:n3��<���gitnA���gRƍf ��V�������m���Y�*�w)Xuz����>[P�Aia7t��˜��s*������A�K����T�����E���p*S�"n[U }�
Ь��/6*v�[��p���ś�lv^�М��FUUp�=��f <���j�z*Rv���|竳_/7������s�U$
�;Ծ�n��������>o����5)j��s���%������<sgMNߛ�\P����E��vz|�x�p���zڞ�g�e�&��s��*����e{�=���rT�S�8�9����fj�>�d��:�y�"�'�y�/7�����<M�1�ɍ�Ȯ��E�nJp�ާ���x����f���~�71���+%���W���]��D�W����W@X4���{,�蚂�۵{镾q�=�*B�I�Nq�4�%�u�2%�6B�Kх�&��_� |��v��hs���ou�Jh�^n��z���n�xs�}���|������
��,�Y�M���}��ަ~�	�w���-��{&��)�|:b���/g��+����A�Η��!�+f��xZ�lq�uhT�ۺ_GC��ٔ>��ޥݰ�w�Z�r߸#*�m_d<���x��{\�M�V#�Tcs9�x�p�(�Ye�n�K�5ō�`���5�z�fIf%�����6��LJ2���ծP<�^W91�H
V7:빸�>V{�A:ɖ��ͻ�V�o(8j���`5;t2)Jn-x�h<@���8���l�ȓY}��_RS2��\J4�fj���3�,`�C��:r]��%�9u���l��	I v��/-"�t�s��*9"��׻,H*K��eF"��ҵ+��ݚ*��t'=�C����yJ��K�Oj�mjW����w*�t�,O�}j�F���F��Fn��ü���0�8��7����U��y�nJt���AS?e����e|C�C8�'�<�����C���JuO_i|�/x���$�S�y�uݺ���2�<�Ǧ�����[��gPO[��%*@�e1q�s:���h�>ň���6	��]Zҥ�%�,��[ډ=��W\�*CMe�gW#m�n���p�������l���m� �2��r�/fԻ: �'l
�QS�e���N�Av��,q��oC%V޹jβ$g����R"K�F��� ��f�v�.�e=����mj��R+�^w-S�-�#�z�|��p���g���囼~�2L揆:�b��:��h*lW�4������R���b��?����zş�c�b�2�x=-�����н�n�;k.�e�P�e"��8�2��3z�ֈ���@�b:���xO}��I�=_ww;����{h��9�՜��dS¬��<T�AW��\�Z�i���*2έO��=�;Ǽ�s޾��.���㹈�v�'�q!�L��m���=R�����>"�m�˫�$YA�N���W����D�[�������m�")�w���Ye�Y�.�SǰÜ&S��J�.�[w0�੷�<�tu�+x�g���}�6����K��H���r5I�O�ba�&fd'&�r���4X0�p�̽�Yg�dV{�v�t�{��q�ς�is�OD};��+�59�hO��j5����N�:��*mH�����]Li���r �䯂˼�E��s��S�Yq��
��)R�Mk-'CjفL��V���31 yk�DEx���
��$Vf�wp�ڞ�)%��]�+q���h|'\��s@橮A�t����s˂5���Vj1�ɨ�Y֜�go^DD�9��juZ��s�z�-��Z����wk5���
��mjgn��Z���*}1�&�u7e�X�ڽ��R�oE4�'I)��tfm�w߭��=�@D��%2����3)��6�$��㯧��ooooO������u�*�
J����$�h�eNf�d�#^3��=>=����>������<�� 9!C��#YIM	AH>3ۯO�o�����������|g�� )*���f`�`ѐP�%IKM%HeY y&�1I�CE5BSHdn��d4�1V˕m�U/�Ց���J9�Y4�EleY��%�������%��Y�d�i.ɖB��A�P�I��y��ĝlb��Rۅu�N�D�uQC�C�f�NH�1	Hl9U��N[�����)Ee�����dU;P�D�u���FI�RB��vW�.���SKE�~��=hNu�sQ��t|�;�{v�|���,������,k��yt뮻������nz�����f�=]�WZk��#�{�կX������23Z�7X�k��<���p7w��&&��q��ƨ/6����{�N� 1�������ZI3X*�
�cm���xi�t��|��'�B���"k+��*���6�&�Q|��\�<�yL���q˹8�>`(�O�?��ޙdZo6|P�8�0��S�PP7)���uC�je� Լ��j�R��`,�W��S[��z
p6�<��m����2���PB�ɯ3z�zn�vk�D�DB��l���YH�ٴ臬,�C7���)N������O�a�f���x`�[��y�1:���5�K������z�^-u`���q���S���z�L��{H.%��H6XRX��D-��C*ͦ9Y���x&�y\�l��
ކ�Rt�����}\����WsRT@ʻ���Ҹ�K؍������ͅ;]��aa�Ͷ聑/vS��z�~^��P8�����:�j-:Y�}~׊��9���NC�Da�m��@�u���;�qx_?�/4a�`���Zǐ�=/����y � ��l`[�_�����x���xi{@�n-bY���;r�ݔ d\�(J���)>�u��4/)��>oa�墁2.��D6H�{3��3!1�uڳZR�3�VIW��\CJ'I>ܶ�wf:}zdsyͬ�[ܦ�ƫ��So���@�@ŷ���|���d���Yy��1��Wp���L�l!;��n1u��$s]��[6)�ҕ+v��{o-�鞸�����{��x�3̞�瞹��|�T��EKw=�o6\noI�9Da��B�f +Ξ=�ͿS�>����_�Qd�þY�3�ҫ)�������Bn>6�7��g2G���@� �uI�֣�0��i����:(�ś���b<=�(R��q���lN?a	���q�x݌;iB���4�$;��XSL^Esd��˞���A�T@b#�-��u�m��O���-������=�! 0��6Va����-���U��x8 (�N���-�<`8YKiW����\,��H�+k�������>9>�y�&V]3s<T6t`���Ȇ�*{���?���\���[�x��\�S:�ǫT���c��:�InNI��u5k}�t���ے�@��b�N��`��*��g��gi g)h�L�@A�c�Jy���n��rK��R��M�wi&���X�� %��G��"Ԁ��\L=>�{�"m&�	���pM;�Y�Ʃ�^�G�/��9:/a.��P�O����������8�R�h�b�S{gO\��xo3V1W �+��Pt�C���@D�^+mG�Z�܍���tQ����ʏ��.f�ݡ�HB4��0~y��"1o��yd>�EA��35��g+-�v)�#\�{��}r�c�=�$P�(w��D�-�8[�+�
$B���c�W/�EF� J�ȵAB��_��z��������<�0ݵ��+`��\�T���53�h�`ۭU�b������w5��;�n(	�$L0�1ȿ����������:�i�k��k%8v`��e��gN}^@L��㕲���g�f@դ�V�����r�/o�V�og$ �>Y�6�uw *ݑ"Y��	I��+̻��ʟ }����Λ�w��27r��Z����D�)=iX/x>8��������P���P�
����2��{ S�qx�����f�Ay���2������5����ȟY�ǈ�lK{ix\l<�W�F, Z��bד�\@�P�b^������Dm��{�L}�pd���n/�s��d��1%�r�����X����9���Y22�٦^�zd�ў�+S���Mk��fx���\�# E3�%l=��z�i3/%�bXU��2�D޻�l�ü<(��!1�d�3����XÕ
��������	��`�~JKxJֹ�nǞ�-���y�yy4���H������xč�pCA�j}>�w�Ⲷ�ޜ{����J�!�Q3����wQ/W����%��\=�� ���J����h��\|/���@�����_ʛi 3v�ݺs�}�g0Z��1-h�k��:�SQ�7Q���8�6�kk`+U���d?��o#G�o����ܯ̐���r�⹟�w�JN6�l�RFe�jinis8����� ���؄���*�~ԺP��G�{(�r�ἡ�W=p�:�-�)�9�$j92�)�OP�ۖ@7�rs���齳�L�!7_=�4!�6���ν�:�ߧ��f<���7�<��ރ�������qZ��I=��w�!��PSL���L��*}�.&����bbr0��{���K��!��j�Nb: �����E�i� [Bp:���K��"�]Қ3��Ɋ��<ڬ�f��;��=M"�G�L�?��6�>s��������G�@�G�/��ٕ0��[o��sJ������E�<�Q
�ګΆ!���w>�ql�	�u�X��VT��JЧss��`���Xp��fV] $�Rd�q.��lA���q�7�K�qa���Mz���zC�.��n�G�[�=,�VG�b=	�d�Q6G��)��(^Rs�PK���H����_X���zo02�����݉�\��)�+�V0���v� Mߝ���D^É�aǭ^>f_c���d��
ׇ�MA�*�N�.z~�N�Hއ���k����FlRRcڄ�p
��ȿj�1je�4�|��k���C��!�CY����
f�9׏���@F��G+3��p@�~��:��#�#iK+Ic���s=�Z���)��.�,2�q*M)���#R�D�����27^J8��)�����2û$�̜2�YE�)��)%鋏#�Yu�dӽ&p��{�3�*I[Kt�ӹ�t�ڴ�*�eѣuD�uz?-@���I�du��T���x��z~�[����%�!��z����g*m��;��=�����:��{�ߞ|��x��Y�W��1&kaO���+��3ql����::�IN��)��u�o��!�$��F��	�ܷ70l�*=l	�&ym�p�51lL=ʡA��Ϊ�%��!�rt�J���mx5>�/.�M~S�i�w=b�z���H�"|L�p�i�H���%���b������^f�%���a�]��^[�V/c��E8ǌ���r�Ҡ�49a��W?��/��z/N�Pp���I[V��z�up{k;oH'��c��&=l�N���݈�P5H(��d[C5z��m	�U�7�������`�o��0�v�R&�j��{..=�����, w4j���<�p+�2�u��]�-XY,<c@9Sɋb�!���O�ǰ���cy����ir�����}O��b�w�u���	�+��-����sp��H�T�M��םӀE��JLE���Fv����wWmU^�a���h�n�>�7��E�瞙��!*�e%�󈉸H�MHv�=[Zl4*�X���U� K�\���rb�f%�bW2ٽNk���b�<=e��g�%4i}��N#�'�s�zy��f�x�+a�DK�7U�y���+�~7�w��sv�2]N[�	�����s���w%��ǣ/<G����Wl�$ݦ�٫,֣u����ĵ���knO���3.�m�#(J-��=|tZ�q3�7�(A�,'7��> x�5�b�ׁdP���kfʫ��غ��{��s3����Jq��א���tmSz����A�K��=����*�FN�1�D8�l�!t�Z��c���a͊��h�}�|���͈�YI���E��1��q����
!��s���y]-&1�4*��d+a��i?*�t%Ԩ;3��fVU�h���j7@؞ʆ���B|׆!���ǋ�c��s�%8Z�߀\���qњ:����^�ƀ5ڈ{jF2@�*��/���b��/ا�NӉp����LEs%+w�\(��%^��(�f���빸�w���u�Q�jIJ�`��y\׊�S0���@Y��2Nc�ѧ]V���H����e�k:^����.:�J��F������X67�Gt��{��3�Vp<U���fkI~Xׯ~0��Ǥ[p��(�kH&-��ct7gq��,�k�i���,x��cP��p����\y�n�E�;�����̭�6H�����n&!zi�� #pK����{i���kY���ǪX�8��{����I��r�c5�.�T����j�U���H�լ�����T�^{ʘ�Ef�m��ָ�Oߵ����Hc}"���oϲH]A|�4�>�����>�5��z�fcC�r2�m��㜚��R��2_J�,��M��Ï��+���x<D��F(�C�@�}���MHV[fa���\�JP�Iwk�5�M�r1:W��YeZ���D&Rs�A?�7 ��.��7w�UQ{��I��}�,�0�85{Q���`~|~��QB�������!����s9��e0�p6E�F\-�j�p6k3W�I'�yH8�eK`3z�j���OJ����=��,�TE���e�S��({�!�<фȪ��Vh�X��vw�'~9$��c�n'_�8��#`�/w�3��m>�,�Y\`�.;kkZ9\�Tixnj����*W��&�3��p��E[��-'��q^z0�9_�q`^���s*K����8%U�-�G���P��/Tޚo[w#����ck��-�y;x7�9��.=�)ƂӬ	;"�r~�/{;{J�vb��:u2��%˟�)0ޝ�{���N���� :�{��+X�{�^�|���2� ���2v��l�����'�{�]1�Y���E�a#y��\�!A[E(L�6�q�1�'������w��s������%�dd����|`jm��7�H���|���� �����&Ѡ��[�߼��Ɇ|OW^>���8cJ��l�F*�'1g�0yS5���9N�*C܇a"�g|w�uz�6��:�*��}�N��;N��o�E{���s��"�2���ܕ�W�'�ނ�mu�b�`I�LX��N^�G��n�����hH�e�+�3*��o\OlxG,/�=p���uŤ��km�`��Y��"�$�^w��"w�4O�r	o.ojm{����o�����~��ә�~��Ĵ�wr���9���=x�W+�b
k��,X!k���Q��/��棹Y�u��
|:�F�U+�_��љ�|x؇3d;�	�V��o.��ժ<��,���D������f��9h�I OL'�L,b�ɞz�1�(m��Ξ)��&��S'q�)�oCf����R)A�YM|��Zf��\P}�漖���#yȬH�5}Ճ��ķ-d8e[��Χb<�)ǧ�-:�s������R��_��[���6�2S�C���2�D�C�b`����:C;A;������w�A7+~�m���[A����2��Ƙ7ն�yT�ĀÄ��:Q�������G������E���ids�ڝi�8��ԍأ끽U"du�&O(�����O����0�1�#s_����f�x+'���x�N@ĵ��z[l��(���q)%ӯ6���:S��=���,�aK�S�u,&���C�v����${
�Ϣ��IC[�27ѭ΋�M(�UoT������#7 pR|�Mil}��Y�^��_��ڏ}�IrDqg�ze2�J��\���6��d�	�i�c�]�e-<�d�\W���M�>f�gA���k�� ��%�`�/vF�\��9�@=0�%����j�����/u�J����y�JrG;4������xtS��X�YI�d����O���|�>ưyaㆳ�ϴ���>�]WU��Y�:��:��"Ն�T��ֹP���xc>�<�<�|4�b,b�����}�y{
F���ƾ-SB7M�$�xf����G�+aNV�^�-�鰄�5��6���[<˭��0�n�+V�(,k~9���[Ss?���.*�&�`���)�C$KsL�t����A�O�=N@7��E��ڷ�,�)6����G+<��Ln��迭h۳
,�':ݫ���j(�j{�ILu2p��OI��X{>'�G�����*1�7��j��}B�7�&�UYM6�wfi��q��"}��}^5���l�({>O���.�b�\��{�x�kH(�x�S��!�m�8<�%�]��	��4���e������z��]ɡ�� ��h�/>��S+��'��z�0��f���Y?hKڀ*����vm��o�9��-H�I���)cevC�o�����a?���`��!C�pf���d�]�C��M"eR���X.��N�A��d��O["v��e�8�o���V����;���c��Y+4cO���N`�~1�X��hp�W�S���s�TU���J���vs�4�A`�var�D��X�0���BA���#�o�wr��a�`�l�z�\=ݔ�ǻI�9����#�Bf�P���K-����ʶ��h�x�7ٶC�l@�*��d�� x�k9�;� ����񞶣�X��k:S)����ܭWu+�"�pK]�g�kH��3�}�y�$�LR};[$.y�}3��E�t�w3o�è�+�+����S��&��t_ҵ���gx�_��tI�ԡ ��*����ԥ��3�0J�#Դ��¼d"C�ף��ǖR�k�9 �$wFF�3��͆�������4bi5+-�45�Q7Cl��o���P�O.�.�/(<\l�D��.����/w%_���|����ŜW�m��ݨ��Ld-+��r�	L��/�7�S-%�����َ��u|��� ��1NCi�!wkn.����Qh5n�D�+�����<�F��+˚�s�w�*`�pl{�bC�f�\���R#3<xHu��_N��|�`�Qq�����[*���2������D�FA��E"Ղ��S���S�m�\�L�h�k�n�ު��m\�u�2����޵Վ�������.Eێn�H�\v��8��N{(%�Q*Ի!�U��:��AK笼�ג���#�"�C�EidJ\¾6�9�W=�+{�)��4*�Su�x�gj�8�;��ΌUƉ�CI��ry��1�ްt!��PU��+�Вh��������8�!��]���^b��l��?.T�B�u�\��{�f�u ����E��}\�9��
S����$��H���୺W�c�j���f]���E��M �c�$�y�U���l9�t/���{}��5KnF�4�RK�(;��Hbj_$3z;�D�����}8��0��L1 ����F�-����e{f���{��h�� f6w��K�	�d�XL�[�����1c��^�K;c<��X�
�y�ū��{q?�$���ܥ+��p̀U��Aj�r���Y�X�B�z�h:� ��v�V��Sϳm���u���"�bɚ�q1��;����\��.W���,�X�Uu')���7�:)���H]�3�el�z-���f|⇸��T��u_e�|����"�:�LP��|�m$/�[,��{��v�E�>�1fc*�B�Ĥ���P��E ��CE�RWCf�o0�;��O3#�׹��Dn������KM<[�Zjed8� ?�"�{�PNI�H��9���g��A����b¿��sON��uݓZ=^�$mHc�1��kT��_��J����W���{����
�OR�=��͍��zB7C������9��d���+� �wwPr�OEͭJ^�0U��縶ZN������Raw<�C��"��YHm>�RiJ S���/W�����)ڔ��v�no$�gM\O��Ҹ��,��
�IG�G���¡��*X�;)�G{MV(�-]��yn�-�����8�P�`!s��!P���Z�NMY�m�(`��BVMI0���U��E�P��t��K���([�ii�P��p�;C�Ԏ^n��
4�إ�Ԣ�\Vl�NňC۶y��I��a�3����9ZH��Lu0��=8�e�G0�O���j�i���N��>�%3)r�Γ�*�wW�����V�F�ƇC#�Ǻ����1f��텢j��y19F-]���q=[}�5�' h��(f�c���W1�
��;����`=�fSj� n�\�)�WAټ^��ﳦr�2���yy��[�[��5LjZ��J�-�bY[l|q����1��[�pQ|ox�N�=}�-�9�B�K�!���A��J*���Cۜ�&^�v��^c�-��@�6�&�^�n�����X���[k�<�җ�}#'�/a�|Ex+��Ǹ��Hl��A3�h���A�m6C*2�_# (��H�K䐁�np8K(YM4!i i�`�"e˄��@_�|�,���$j&��?5./���?�?�YD�4�9v�ʙV`SKIES�n8�����}>�O������8�� ��n;8AY�l�@VA�Ye���4D4c�==>=��O�����>>>8��02"��\�#	+,ʹ�]�J"��˄�A[T�=>>=�O�����?��x�>\�(h��2��22���JSUM��%C�A�n��fA���NAEAXbQNI��id[a@���M%S�@Q�$@�Db���Lf�@e�AAVn�lE.�-fa[&�m�aBQYd&A�NNY	Y�UAFBVEQ�Yfộ%&@Rd�A�fl��Qfm�i[��ɳ�a��F�P�KQ!���R�dE��9lK�A�bY�ade��d�u��=dGU��'+�{��s!]�|���.�<v��+>�oy]�q��q�Ji���8���VNt� �����c �A&R���r�p�Ӓ�>p;�z~��lOٓ��>S�/:��=Ӗ��"����_N����>��4����Ҿ�-L]��ō�i�������Z�P3ˣʡ�h���	��o!Y��[��c���V�>N�$�Rl��T�jz
���S6�&��.Hȱ����P��c��֍��dy�+�ƛ�Z��b�9�fr�y��"²"m�
9�
�z����"�N)�q,L�O?��Q4��İ�	�r��m\�y<fki�k���I��r�N��&�N1���O��jh;��m�R����B�N���y%��N��� c4�tB3D����[�8��]7�Pye�\��V�'�\D�&a�������S��~qf��$ݎ��j���-��[�Z��VL���k��i��"�u˝�ү�m�����ڪY�X��n]�#YM��S/�{9�I",Q^&y�u�#NRd�~"���f5rN%���֛�����;�hgpF5�hY���<��%������w�8�d{#Ť���%�$ZK磦��\7�������-7�m��R�aS��U�q��E���r�o�Y��1�W=�Y&�ٺ�M9����#�>9p!��Ks��7����e��O,k�����X�Le	�����N+s8���|t����Md�ڄM��P��?���> `�Mq�ZS=�.�ߒ�"o�ǫY�;e�T%RB�,���2�Y�h/G(��qW�v�^e��̂�*g�\/,����*�X�57�9��ϝ�]2�lF��m��D��v��!�M�pӎX��!��a��%��6f�7^jP-��V�|e8���_R�R�;ð�����)F���R}O=�'Vjҝ`�(ɿ:LbX������7���*t�g��U�κ����bX�Y�vm���J��Cu�{bѡZ�����l�����K�_��=�k:���Ƨ�<x;�`�4z���&'��y��U;����<d�zoV7ƹύh�M��0���7�fڱ���1�����$&� j �:a���z\E �a��K��C՛~�a�ZU�7s�L_�O�6�W5�UN��T����ZC��@���+]�+�4�m���NzQ���7��q5qf<��Oi�b��/��������moT�;�avч��2�3CF#�.|��J2�J��M���b��X6Po<�_9�>�KRV��b.:_O�kd����;����/�{�{�^6��Վ�NF�}� �s.Us��[�ս`���S�6|=�D�f�[ty�m�fV�8�k��6��+�����ՙȾ��T�[����W�-��0��T�ɻ�;T�=٘&t����?����
�V �(Q�N�׮|�u�<��~��%�ɤF��~aş���=1�]Ο�� |�����ӛ�Ԫ��{غv�����d��C�y���3��S�*V�@��F)�Z�aD:k��8��g ��E��y��L_��3}ZS���
0�gZL�A�j��^�StH)3���zC�*��\;��D��\�=w	����@H寈�	=��<�������͞r��o�$0� ���S��Kw�V�$��tB�w�*���њ�Ӎ˲q���F�j�h��������jE�n��3	5�@�`��_6�8�Wcz�egt���o5�H\�f��]��e����O�M�G��: ���ܡƄ�8W�؅���@J֎Vw���|��(�gǥ�C�J�u���"׶�@����L�1�뷢�ϩO7�^�B(Urt.�<#�tV*��s�ru���֣>�#V$����ؼ2�v�;7ɇso<��K���h�^��WX���	�(ܶ2X�"�j�0�Xsp�ip[��XiH+���� ��RR�qO4T�`�)��fÙ��z�Y��M���WN���[}��~Ɋ��?�l~-'���#��C;;�K��Ec	j�OA��]����V���$͏�UTw_TW)���Af�#�� ��?���W�Q�2��0����$"P/�K��6�rQh�?�R�n��ns��z�m1�Q��@V�E��Pf[���N��ͦL���W^gE�u'�G�>E_�%=�I�W��ݦ�U��~�}�L��i+�$�5�4ϡ������43���N�\���,{XCߵ�T�Vz����b�@�8���F�}w�Z�+������䧷n�m�8�&"�E��dj�d��oo�E�m�UG��j��j3S	�؝y[��>C!.���u�1:V\$Ɯ���>%ߛ�e':�?���#���ͅ�a;�X,6��xg6P栽E�,T:嘛�_ԅ, ���9O��屗lW5�Hj���!�0������G)L��LMy�V:"�g�S3�T#8���5�\�&nб�[rɇ�MH����-�Yt�Q�0d
��tǧX������RU����O)1{@�2Ocwk��Qa��'�:�)�$քZh]��#gڛ�/G�_J簺)?X�"�
����t���܋�=� ��\�1G��#�ޔ�C9���O���[peOl3w8��T��LL2VɃ�V����*c8\&��)��K����:�[[��3;Z%�𑪟FZZX�P��=��ڋ�o�#(r+�y-���/Y%6����Dgt����]�ES�YC-W]i(�'�v��}%vOD��4��7)��"��������am��9�o6�D�پ��GWGF����]�f`'��0��%�(t��9Ϧ��@�g��R�pu�?E��=|ޢ�m�5:i!�y��X�ZM	������i�&7UM� �d�,�셞n9ӾB�n��R�/�X���>�/����t�� �f�nQ�h8\Jc�Fɦ�tn=u����)�y#!μw9��<��1����[P"����2�(��N��=��Z1�7M��NٹR��1Z��\���\�׊r��l;�����-�[RH�T]6V=������4o�9<�~�}���j�-7�"��8�W,V���|.7J􉚖b�/Ua��M�\qe\|�K�L�S͆L:���J9+�&������$SH���cpu�O{kaڵt`!ߜǻ�IV��A�^H�o�E�s�`�VG����k�1{�qbt⃩��s.��q����S��k�����6���+y%��i�0E�SN(p���X�����}�,x�C��xEg��ŋ6 ��p�m1��N% v��{���Z�W,,�N�f�*T�xD�!9���tk/2�iN�%s������ؿ�nߘG���iG�Q.8q��)tV?��qj+��c��G�m��s�V�Ð࿮u�Iϛ�1�Ğ�����^�����x�:��j�$'0�R��h�u�6��!��&���� >f]r[mf0��7t%г �/��P��������BM��M>y߯]oy�=�����_9���G�eRW!ea0eDL�D�����x����Q���z��w���2��м�#����7���$��!���8�2`���ʺȞ��>9B#��0����:�O�PC��SEh<�'_�|}��z�E��s^Ѕ){ܓ�댼P������V�"Π�ܗ�؜�-�R�1�D�Ʊ�Ǟ{MǤ�7~b��k���Q�:�\n�R=w������+�.Z��[�����p(���fddLi���r76��3XؚC}3���1��^�b��OU@톖T�HASS��ij.x�܅��9X1�N2M;!
�P�v�ٔ���2��JB�ur�٩�Ȯqm�$�Jh�k�.&�3B�T��w)Nn����Rp���Oz�C��}9�뿥6��M�QR��B�hg�C2ת��Uu��=j"}ש���)���7�o��UuȜ�gf���(ڭa`�%���y�~����������ZĘBIc�F1�}qb"~��lZ4*�O�;.����]��k�hj}jB+[�Ԉ*^�o90�>p�H�$�{L�v�P�͸j|>#vk��J�E&J�b3Q_��y��ri�����֧��xa� �{_��\��Ch�i.� [NE�C�C������;��m}p�!srSU���k�룺?wS*͋��ML�Q�]F��ݸ�an<ɱ��o}����:2� $
~TH`@�TD�A%�B�C���{��k�M� �a�\4�CZI�g/@��t����6�E �a�1�+c�&�x%�fEukE�n�b��Y��E�g�L���2�f�!��`I��?�L�\^�A��\�bʶK8�r�u.��	����a�l��MG�0�P/Q.#�
@�5�,�>�ϮE���rw-�='�ǁ�jk�S{u���ǥ�i�V嬖�AQLlAΉ-:%E-�l;�%���ڸk��J5tD�e��#��i���.oM�u9��yADڦ���0v������د}p�㒴z���_��L
|A�����]>����Bf���������m���w��.i�a�sa�ʭ��v�p�	I&L�s��A�?0͗i�I���Sp��0�TI$aխ���8�����OcQ��ު�3�p�<�_ݍI�L_=������/�]���(����n����F��e������QM���X��8�P,
��yJ������ų�j�٣�<8�f�^��h�D�Py��$�aiT��ī�����+tw��="~-�[Yw�!�yOwD��n��}<1�mz��%ǃ�ᒇ���B��wѰ3];zU���O�>����S��J<:�)��uot�j*iê�	u�^2Y��ʵ��7n��u�� ���m�w��w�{�w�����c
0�C��%4�J���=���98���-�C=�8��@�<D��4g�=��ޏ���r�q��q�kE*�WA��~��_X"�q�\�����x>1���@g:�)W7�r2"�Yb�ɜ�jƸ2��*)�H�#�0#6�pS�^䴡t�o4�7ߚI���0�y�S�6��������CL�GW>��1�HKo9�:u �6��u6���]Q����L,��p�77���1X�.��Gi��pe�Y9�:s�E����dWX1�a���f�tp'�����f��iHw
gx�a�N�B{V��V�E�sc
.���ܿ�:��f|+�����=��So�&iaW��D�@XG2��sV��������E������)nT�./%�p�j4>{�Ví3V8(���SH(���ǩܦ�����.�o4H���=w����N�4�+b&��2��P$��z�hu�nU�ҲJ3 8�����;IΑ�z��Gza�ɫv�×�5���T�ѷ��\:;J���ro��oQp�t:����8�ҏHBJ�S���NX��Z��2g��(�r��Qp���4(c3��� s�i{�S��d����q��utr�yՉ��~�8;�o�	>�U��ES���9pX�S��ۊ�p�}m��B�x��fӣ���ʸ�ěF��G�ItP��ޞ�A�����2L+��ޮ��r��P~� `Q��h�$F�ZDR�:�0簬�Pi	��E!���S	���o�ֹ���d��Lg}}P��G���l.��IΛn��|t�i�k#�63��`�4L�YQ>iY�/!-^�e��dۉ\A':�Du�$�a����gw�B�]a~/v0p*ؿ���J����B92#������lX�k�-�O�T�l��͘��g{r��*Xv���E;�-��L��$�D	� �kY+�q?����wv+�{���ƿ*i�VՈ�+�H��-,�m� ���G�Զ8��X%��la퍛\����f��(y�x�:�0��	�����t{Y{e�=o�y��&qt:��-FOu�-���0y�����w�(�]z��P�C�׀�����-���WU��vOF�|��B_��"y�Z�	i���_\�Mi;��~N��z��V�$j9XJ�}J�Tƞ݌�r�[T��y���S�XZ�Ȫ�U�6�5�=���&y�E��«k�����ɗ�hD������+9�q�����<���H݂�e��1�۾!��UT*K�gF�kH��ZM�]34{a��t�fE��;�����nV��/I^-�������Ī�dڇGʹZ�҇\�R#jdX*!]�dety`Z�(��ۙ%���wN�E�������t�{����M���+���������j�"���H��M�)��j��oE���0���$M1W�
�Æ�dK{��t3LeZ�d�Y9��ݼ����u�8��a���B��FG�ҁ�yi���8t��ueK<\��!��L�ЂS�W�/
�Ks\P.t?kA\��zP�k[���	����:���{������Z�Ax�D:,�O����ef��� ��u����v�v�.͞<@t��57rb�,��E9�ݑo�Xƕ�u���9�����I �US�Aunݭ�&��NOT�:[�튒s�7g9�C5԰cn��q�e���Y�y���ՙF㦒����-�b�[!\|n{��dA��fZ����.
�^p��F9����q�W/;m@��=w�&s*�Wa�R7SF+�]���S�5��DE)=�ZN���KQ�m�i�v�D�8��*��{,��2�'�3g���%:*<���`?�����
��)4�sJXVsQ����y��MkF��*�s��y�i1;#|��xX6��ފe�q)�0��n�͈�p���#���s�K�ۺf6�����t�$�ּ�*�������:��^�#�%�4��7��)���y��ҁ�j��$��GFw���5�+�\�����4ܻh�.�r��@���9�x��>�}%Ӭ�YG�`�Hj�md��j�v͝���J)]ύݣL��.+n�s꫺�M����S
�r�<����ǡs��3ή1Ds;&R2�k�r�;OFX�|A�k�O'r���b^��8��uoH&5݇ɶ�^�ge2����y;�܊s.ю�#�YvN��h�t̊��Ka�/g$��G�wt�D=Ϯ9F�9S����+��gB��s��l��	5�AP��5�=]�31��w��/�n�[��iq�7���E[;�%����7aƶ��f|��@%�1�䱌Eouѻ�M2!!\�s�Yf8�����X�����et����6��lI�-/�bhx�=���`��R��K�*2��8�ju�(�9��an
��2Ɩ%14)v-���}EHI��lj6М'u�J�^���>)��y���M�A'_x�Q��_v	�dk��X�i�d]�i`ϵ�'Q�
U����S���hHw���v�kfX*z	;C��c��TR�/�{!���5�Ş�c��d�.���c��l�F�^��n�L�{�Yi5����)��0~ĭc����o���9 �� �����.!���+�����%�E�X��{x���Y�J��+۫�h��t�u��u
y�Y%wu�[9��� %��ՕX���ҡ�9�o�u-f� ���*J{�e^@�"ɧ�������=R�V���m9oJ�d��G[�̓G)_KV��G��*l��39���6�+��"ǖ��0��L/�t;�Ǵѕ�����:�u���R��Wm7��W�C^L��^�1gu�1���<K�'�Z�Sʅ2�v��f˧Y����JX�e�],<�yV�F�VvZ���P��X9r�����T �3r�
��*��\%`+�;�ߋ18f�p���Y��y��6�)}��5d�KO�f��|#Q��P(EtΦ-q;�^ъ�ƭJ��L��'+@Z��7A�\5Mſv��I-YK�\�؞{�7����|e��|�饼��2���)2��*f]�Iؓ�Qb�0ӷ��kf����uv����}��0Э{�.w7�Yܥ���Wc;���\����*cr�b�ݰ.�����H�~�����a��s�Q��.�qM�]b��]�2��^���
L�fxOS×�I�V=�A쨯C�m� ���T�ڰ��D�vfPdy������@��3*�0��3B�J��K,�Ģ��Ɯ�q������}>�O����>8��y�>Y$LI��1��l�e�R�كA���n3��>=���O����||g��Ϟ)y�bdE�$NC��QEYa�aFɶ[A���M��D��>=���O����||f|�����U���&^fa9fa�Y��fXD1���s"��!�Ms,�#0�/S�A��fQ�1�M�eu�%4;S9YE��Q���@��eF˶A����2QV`U�h�ک#2��(�2��0z��r��l�����kp�c&�̀���Ɉ"��r0���j���2,���̢cpȲ���
%����(6L��
*h��	��3��2ZLk2#0��,�̲͌(��odn�TՑ�K�I ���͗w3���*��}?���>C���3���V���zQM�:ٹ�7jEb������B�>ʛ���_���|���+� ~�Ar�)Q��%h�D{�e��	0��^ړ�	{���h�\���X�;i�R���^�sy�PW�:؎���)��j3{36GI�Z���:���l��B�>����ȟ]���ʎa���n\�o�^UvW�WN'0b�V�DusI���L%J����mwI�_עѡZ���%\�k{έ�M�kS�Q��ZRXHZ�:��x��B��� ���@w`/�Nz�R�vEH\`�+k�
��MmB$��af[�,�C,%��-@j�hkHŵ���D��F0G�aq�M��4��z�QW�N<Fg�����Tٹ�����=^yǴ��РV	���f���~|+FdPu�w��3��#��!�\����HRu��Ѵ���L'�K��#I�b� ��4������5���u\��jF�6 +Q��TM!Be�oM6�!��}5;�ɿ,��޽��.��`M�A�h-+��Zt��M�Pe�#�;MDe��&���N�oe]�j/&�.]�����jF?�wU��9��edl��S�A�0���?Ǣ2WO��^潮�~�efeH����9u3�ܷ��a����'ȣ��]�m��2>5{�N7��}K��ýȑ�{ѩǇZ��Z�B�4^�]s�[��v��W���L	W'Xw�Ȼ_{D	�7�w��\�uB�%�M�Z�����c�*�2�.��" D��$��G^_^��7�����˦��5����s��J��B���fOJ��u�Vet<�� �l7���*��l� �R=��bZ�T�zbY_�W����N�̌�V�Je��Z��L����ӷ;Sx܉������+]̄�;��{ sEv�\�XoD&X�UL��آ��K��ËU;7�\��$>��TqngY{��ܐ[��a�a�P)`3��2��P��%����K�"U[w5(�坋1�I����1͖�,��.�dGy�7.P�S��=��.�[�:G3�b��J4��tw*țUoL�=)�ΪZ�Tf�6J�HvnVa�����ύ���Oii�&)v�:�v6PoB����9�r�e��j8t��+Blֆ�pP3�"�fi�,��y0����s���Ǽ��v�J�Įk�L���o�'QA(��P܅�qQ�`�J�a`��qW��dA��GQ��ۃ6-?�Dy�.0��>Mx�f��Ԫ5�/�_���q�%�q��F�l2<�NP߭Æ� Y��:p�Կ6j�Q�}�!ŖV�ʤf��ң����{�	�ے5�h���X����R�����F�ƣ{!��6�fsb�YF�{s[�A�]L��Ќ4�$��;���a���,R�8feN��9k������'PiA>���U�dup-���+�M��M���j���Vߒ[J���x�U�UH��� �MY�n��gYgE��P�� 0pG�������׿:�0.BF$�x�G�8�"i�<�C�U��sV�;iX�qn��F��J�����/�p�[RA��+b�����v!�6<���.��~S��Ӑ��E8��d4d�H��,r�ԍ�R����y>�Ò6�lGsԡ -�\�bt��I��xhN���-q�2��$x��Z��	䷡�L�.�u�|��bF����;� � _:`���XAz�xk�S��,z'�^��PqL��f}�1{�R���8�9W����E@>�7�ZkMa�3{-ݤ������sع5$�9��L�	����I2���-4b�N�	���	m
r�/�y�ǲ]�_Ns�ؠ����NK�+t"/0��/dt�ȕ�`�e�K"��6ִnu:��i�ǜ�9�Q{֙Px[��h:�-؆��2]������Ǟ9臎l�+r��'xmNz��OGI��80�|x���,���c:�N0�F�ÜHj�8�*|��?`��`�c:2*���H3 ��`)�b)>�CZ@Vn�ߤ��<�ޑ^�D/p�1�^ޣ�����~����J��Βr��mP̎�vI��6�pT�cQݥhL�+�^v$�|V���k:�x�u<���$���r�5iҺ ��k�����[�7*V��P^�O�j�_�P��n�!���|�|��s��z��νh�ZC�eG%!�\�P(�(R��JT��y�γ>���޿X]_o��&���Cg����(��1�$b�Lkm{{jD2�T|$��|6:�j-%�p�ێޘgkP2bs`S��<��x�}r�5���G<Ϡ,h���"�O<)�
cm���Hpe`�Ŭ�1Q�>�:sf+X=sY�q�[V����ǓV5�ݑ]a.c8�/ni$����X`:��i�BSf�]uELS�)4�]8ѣ&k���`�]��(Kq	g��6�g#i!l$2�d	owr�z������ESt�}ŨZ�u�B�FV=���g]�P��C�Y��kL|M������qm�d.q.�6�ω���%���|O�ȏ:�zQɔ�ϷO��w��TT�4�
�ޝhK"9"�m�o��h�7Q*�^2���<=�I�UAy�禽BW �M�Ш��pq��2\#���Iɽډxj������Oi���;Sn�u�ڽwd\�����Z��r����jfiS�'��q4N��לe��\:�@��[b����|��{ʛ&z'��F;��@�m�K�xq�4PxQ��nG+�q���U髰����F�K�U-Υ]c�W�0wX����\�Xn�'E�a;��1���}@"@�t�Z���d�Ղ�����Ҏn�G��J�+zB3܆N|#��F�*o���Kd3�]�v��ڱ}�
W�@��!���0`@|�>��> �<=��Δ;����9x܏>�?�R�Z�������.+�WʨGH�
yEq�v�W�i^oEcnd��u�gb����ENc���i�M�#��H�i/�Y�+��j�,a%"�v��W*���lmu�t�O������nȮ�+��U�]H�R�)6��Z�L�e��W2��=Y#�G��f�Pa�f9?�\��O�U���M�GM��nm�ǛP��.n�-�x���6X��xnu�:h�e��	��x��qp1�H	����+��n��y��9����j]g�yٰ�p��VC"5�Ә��1I����ƒ�Cv9쇉A�82�n� ���7<����i6c_�l�̄�9I�JЦf�X��@��~�{�ȻQ�H��f���e���.��oGs��������me�
�+�8\Ϫ��5xv���\d�:��\ޑ\J���>�y�!8݁guAZ��kyw�yÍ�̕���Nq;u�j���zeչXY�?�0j����~Y߬�z�߫ߨ��e8Ej��7E���g�;��N2�c��y����߂<n�Q0BVy������l�o@���x�Ip�����!ɺ��[�1�_H)��|eH[����hT�H�u��J�_���N�n_�)��-��x6ÏK��z��0D�������T~�C�aWQ`�)J��:��ￛ�����p᥻TG�B��j��� Ք2p��w�X{8��*�Ͽ,�H�}"��ˆ&*��{�3�׭B�o(�h>.�]���Vc�ͦ������C�s;?A��eDs)4fT�3�?���������O�G���2W�"��E܇k�]�hp����Wmn�"��uB@7P(H����p�7N�}���"<�n�
��D�km��aw�u��E�.Mp|��;B)�ZsÔ��C6`E+�-�9m.̞1�&���v��n��	��Գ;YF9~�B�jn}��=V�3���E�ħ�Jq��
̱w�I��D�-R.-����U�ƮJ���˞{��Z��k�	ޙL��e�b���E�ݑ�O��/EƘ31���Y8s0��	�d:�����l0�u����@�dOdz�%�	T���g��e��Q�f��4*�1��o����$�JH�S��,� N��
�p�9�7k��O p�?�s�7��s̬���๣�Ն��eY��� �%���,Yq�#������0����'��{ ۋ�K���4;ZZ]m��M��e� 9�1��v�xi����P��S{q��.�̨����V�y��5n�K�"�Vե���BA�p��Lm�r�J�W�[�x!ԸcR�Y�̭�T���#��O0E��&{��&��.�}u��]羳�Xvo�A��q��P���F�P��_\�{��ׯ���X4<4kX��T��PIW'��9�_�*�r�}�e��1����
����b��ƦY�H�Rs��;1ޛp�6㗟���QA(�局B�i�f�f�׃��˲[Q�yxO�z'�z�Q���K�,,XِՏ+�����an�:���C� �@7�C8�0��֧=�݅�ƒzu�<T�u :�Z��r�C�ҵC�$�_;馚/]oD�/<�]���?{��R���&�D�m�;*�a�yV��G\J�L@h�A�n⋒$8xs�]�Ob��v��x���E��H(��dkJ&��X7)|,�h�NQ�ru�s�V���|Ǻu� y-�@�3}�Ƈ��3�l�$-�\�jt��Lh�S����ͼ4C���.���>��lС��z}��\;E��5��m��a� �iMK��>�nL�9ϱGbp�nSڞ#Mm�A��	��x4�ڇ��ME7�H2�ӝ^$r��v�	�l�YH��)�b�$�W\�6�/ZU��-&��=@�Q�a��a�	�0���ݷFu1�7�Q�H��%�.ꜝw�ÿ���{r�$!K$��򭏢�݅l����`�cxm]a����W�#��I�����e#,?|�G�N�8�m[J����9dD|�^�ۢ�ݜ�*��1mK3�s���kj�����77�糫�����h�����`RrPiP�R����y����)pϞ�zI��@�f'v!�#��$q�Ds-��q��������c�S�Y��k���"iu�q�-k3R �ڣC����+][�փ%w0�o��ڝ`k�^����rv�&�aw8cN:a161W��xZ�a�װ��«^zI+y��X�}���9I��d=��s,��י�Df���pQ�1�w�e�ӵ��a�q��p*!]ԉ���(�4��vg/����^�i����e�9@��R��[��t��We�`$��f������;/��v��m�V:4�[�* t�j�9�N��01o<�\�MdύGC��C3���k��+�ro=��;�`Ū�3ht�%���_51n]�͜7�&M�H�Ƣ��Vӫm�)VOv��N�+�gX�?��ŋ+SU�(ܴǝ
�j/ʃY�S���җ�Xcl��;F�N���J���^�١��V���"Y"j&�H�Q�0]+1����^�yޑ�y�d��[,3�W��Ӓ��.lK�ǫV�J8 Ǫ�P���wE5u�;l��_4$��Mվ��0Y����P=���4��D�D��������E|�s�٦��ҝ{�SY�Oq	���w���e��a	QT]TBv����]���r©:䬙`����ت�!ɗx���  Y���#�P�P2(�F�$`� H��EM,��-y�	�s������z�_ׅ�U�5������\�bt��!���]�WCV��9�j)���&�j��b�j|�M(����R��z�����UX�f�P�_��/k�島�$�9�y�m�S� ���dk�P2�y���m��JB����q�}oK�NȈ��w��k���yʑU�i�a�B��@�n�CN�M����x�L[��]�ml��)<$��]��nl���_E ��,Y��썃&dmKϙ覺QI�eޅ�;+��K]m�5��$�Z��!1糱I���l�T�8��'9�6Ӑ}#�.�t ZO�7�E�UB=pD���l޹TF݆M�U!�t��Q��?5tl�ҩ6�&��͡X�+��5�#������{a2�S".��sbto_���q́N4�`KW6ڀ��9n�A�~%O��M���ɽ�~�bѷѻu���5sS7Z�,xݫ�����{���h"��I#}�E9�G� y���S9��k_`�2��m0(w�b�Z��9\m��x����{\N���?��L��M�_k?�΀���l��k�ul�ɾb������b"��H�mu;*�{Q���\��Y�{�d��g6fd\�wZ�[�:�u�9(���I8lZ��WZ10���{85F��}�sJ�Rj���)�]�!��M�i����<�P>����=������dJ�$�QIA��`�vlb6�*��kg���b[�Xx4~��I$�Tq��,1f�X�/]�n�@ۻ���M4k;��τ�3�����|�'=��C��/f=����b��s^���[<�`Yq5�9��34��(�J.Fl��Ny�ߏ���Q�|jh�`a���ꂵP�A�+��;%�u�ܔ3L���ٺq�.�����9�t�TeSg!�}+u���u9�!��Ѷ
�D�˶P˫e���J����)���C�ʈy
N<�Ѵ�ϕ!i�⡽��Vq���#'V��$pz�X�.R~�H������l<���5-�~�i,�M6j�W��%���y�G9n��Ѹ�^AP�z-�(�:LhJ�.%�w���3\NT�"�;��8S쵮'F�e䢛��n������e �v�"[�2�p9��\`�-���;����Bi@�6�t��	�l� q�yp�ˌt����).��,���c]�}�Ԓk7W�ˏ<��E&���,�&�Q-7�X�Y�[�q��Vn��mmĺ aL���rX�Q�'|.��Om^R�z}p!�>�CF�'ː��^��y�zk��f�3�%��r%�]��S��f�p�(�������z����GVL��	M޺�C��%�U�r��ʖu^�N�����&���Q9�o]u�jTс8����B�ɨ�4���/y��r�_�g}��c&<�n�^x��`�F-�W�2�Q���nMIӜ��fjP^��.����L�oeqٻ��k��<4!�(�z&n}-j�p	�Y)1Vj�H��3�ӧ*ov4z�\ծ닾1v��8r4���Z�9)���xxS��g��p}c:��ۿo��u/�
!��+��Q�<�9�3��V���Ξȩ� LJ���SRU��:�M�&��<��w��3}��z̜�0�I�e������]�D�w��]�w������b�����H��Z����ɜ�{��m�|d)y̔Nc��%�)e��nM$� �o3��[��pƔ(���ƌ[�������z� �手Yem�a8�l�|��pn�;��&����xM��]]��"���Ŋ��͂�J��̺���� �Ì�>��gQQԮ#�\5Ԑ������x4٘�J-�%>ocmP������ T��!ϙ`�b2Suv���3)/�T�����n=z�B�X�Ǉ���h�i1ˎ�^�y⼔�a�(E����b���̷��9�e��<ʹq�I�}���L@������j��f�>�ݍ0��_�z����R��FB�1U��8���R$��B'Z�l��O^���n�n[�ј��j��(��zt���R�s�.G)���	�N�/9틐\`�{%�le��0S�t�N���
��P�n�r]�T&���Z���-Գ�S�X�ɭ=����g�7y/��Q� ��.H�Cn�Θ�3ӭ��*��ݵC�Էv�s�2ܾ�ǃ����֩�4�М4m[{��C/�COv򞂕k8.T���yH��K;@t9;୞����{�)2[e����%Xa�tvړ30];��Ł\�$Vͦ-:À+����"�V���Jľ�r^c���Q.��U�\��o8�JbU��8�.��M�,�4uv#P��k���Òh����(��Y�ev��p�'[%e�)�fb�J����>k�/�R�guM5�saV ����v���O�&7\Sm�p��}�khgRxF���ܹA6�yz̓����n�Ϯ7ַs�U{�[����旻,��b��t8ղos��h����6\Ug~D�o��h���0����巌�^ijt澬�L��d�X(y:OD`�v�og[g����;�&~�V�����t��kWgb�cW\.�UN��ۋC�t��1Wk'�s�����Äˡ	���"��t��-�n� ;UX�]�[��伩�:ȓ1�y�r�K2�8.�uT�a��-8�I>���.��$��lIrFdl�.�9G� ���qJ�?@Я�����$E2�\i�-��d"�P*H�)1����)13�L�c��B93��yYS�Red�E�EVXDDw��m���,�
�gooǷ����}>�ǌσ�'̳2�����ʂ�4ʳvܢ�s0h�"h���r\�
��_���o����||f|l�x�Da�y�4U e�cQ��c�A^��fe�V٭�8㯏�ooo�����>>3>�~<�3"b�3&��2"�Ȳ(����
*s0�/ ɨ�(6������3֛U�fd�1FX�a�DM���5��111Q59a��FFU��FY5EPMea	UL�I�c�e��a����ae�mC�fN2UMfa1Q���TF�I��VfY�fY�f4DEfQS�5��A-T�G,�ʨ(���,��*�̲�+'(�����j6k�T|�jh�$���̧�9TV�RU9�9c�cNT���������(,ǭ�hfw""�p7p��EZ�b]�r���,%����w&m�w��������t���$�І��K�k/{5��u���8�vl9���}�.�vt��g�R,̍��3z׮���s�����Ȑ�0�J�R��S��e�Vi�I �����	S�5ܲ��?��Ӄ�C�2�W����QM��=�gxh[jl���	t��y���J�wD<��l�!�q�Yd"�S���nC�Wf�;����uK�ZknUz��r�c[�����d�.��
m�����xKxqi�p���q
��tI͎�[�+��� 8�'�F�[Gs�@�aA��dwE�ok;7'���W̅0Y��d�u�܍����.��T?�C'Ƣ��n�%��R/X�ì�z�x���;t�;�kD��ܭ��
�8Bf)���NS��R%�la�C�7w6�e�X�0��m&;b͗Og%�/�7�BX�9���O�<�PNEy��x�b�����n���ײ��p�K���n��<Z��Q>'�S�X�6��Oㆵ8��!]�A��OuS����)�g��������Q�@�o1	�f|/�Oz�<�{Ց-3�L�4��iʤ��Xs^��F�W8��|��=�r��O�P�,�F듍~�����{�;����C�<JǺ�3�!~g��*%�&U����.�b�	�h���׌mIN���/g����;��6AJ��8�*L��0�O��9�j�������ߗ��B���*d�o;���f�3��6��)3���t�źU,���ܣ�z��;��{뙹����1܅!�+��# ��}w�����������f�&}������&���,`Jm8���F'J��&/D8��l�����p����ʙz&)�^W�Ŧ.f	�*�r2�m��|U�������E�f���A�{�WgZ]���ꈛ��_���:��T�O�N)��dȨF��H�M���Ͻ�=?�;7�~�/�m�%��2�+��� e��U���f< ���*|"������uh�n�Nzyu��oI1�cS12�l8�~�Jn���K:��4&�� �U���S���̽���/��2)��)7��y0,�d��kA���Ĭ F�b�k}�l�05<l��MT�H���p��N���ɕ�~Jc��cj�99@�z���F>4W�@��nv�����,�����`KV��6�#b)>�IG�crF�7"�Gl݌ıɓ��x��!�`��-=K���oZEwK���^h&櫠��H�tƶ�(�����E��ɳW���;�sxi��:m���Ǻ�F��`��׊==r�5���t��Ta��ͪ0_\E;�O4#!�+��iqb�4�	��������s�~�z�yԚ���,:f��Y��A�$�utʓ�b�n�lT���Tí�Y}*:��T���tK@3���.�0d�wm�n�e��\z`Ƴ��g9��uwﯱO����@��AJ��^z�3�/�Ǚ��o����Q��������y�����F)��F�x ee�iFdY3�7�����0y�F��0��J}u�g��擐��`����Kx�`P+yi������Qˮ^Ͳ��I�<�z��M覮�{��
��sӸ�\h�"���=��e�D�LU�D�0f�n�|呵���`.ׄ'Y��9�|������މ�km�i�P��C������o\&�C�32�r�(�!��5ڧ[$p�>f���Ǽ�Z�?�G%�;#���z�jE�=�j�-A�)�<� ��X'�_#،���M5�v}z!���'5TAo0��Ƀ�>b�I��V�7������3�BS5�V���`a.�96���7����O8p��ɽD��J�L��֓N�/����N����5�y[��������� �	����L;�!�-��H��1�y�a�ӈPE�1By;���W�v����s׬�m�U�y�/Uk
jճ>���{JÓ����~p���2��Ǫ�2�4���F�'�%��k�S�e�6��T9#���
�"[�nS�����ǣ���3h��F|j��S]���uj)��w	��'Wvg>����Ы]ӎ.�0؍�����<HW-T����9����̭Z��W��>�-�ӕh"h��}�J���ћR����ñK�m�Ш=c�.Nʺש<��[U��_W��P����XZ=�s�<�ٖ�}�Rd���_Z���H���p%>D�°g=�2�HF���i�!��}h��r:�x+f��oFo'��4Y��u���:�ے��_y)�O�^���O~\W�?p��`����N��3=ǐ�l��ZI���&���o��B�WJ�Z�=����5Z�+uG�R���wjǉ�mH#)��V�aG44��m�H��R@�qݼ8樤��5y��"���:�lܕ��j�E��d�㭄u(5��V���В[�j9A�0���u�L��B���Xaz�2%e�f6aH��7��^1�����q�c7�Ⰲf^۰㷆�RˁƵ��Zxh���c�z��U��F6,b�\Q�ƒ�F����������V��<��q+3�/�@uD��>�c{���0Z#":�H�4�=]�笞�Ø�`NZpȯl��p�mZ��TE	%I��Eų	/F�	�ZK��vѸ�3I��ğvt=p�)��RԽRw\3sV�
��o*&��_��T��F�q�����ɚ��U+k3��,$Ƈ�m՞���P�	��q�c�Q��)�$}٦�H!]��h�^g�K�{�Dی�����De���� �*�"q�&
u՛�ىl�p�Pq��Ϡ�;&c��&��x�ɽ�h�G>7��,�ۖoQ�g]��f替`��,0ox I$�.bYٛ��p��(�y�izW�M�Q��i
�`�b���kN�s-�8e�=��}�}���e�]�,�7���J��x`���ߢ�����	�甂~لC۲;i�H+���=Lf��ƞ[��.5�EE7H�"�Z�I��4Kl^�u��+���zvie5QV�19�Gr0T�=gOu��1���L;�K���W4��9�jdǏ��[{+2Ő)_t�2�w�'��{Љ�LB�[�K��\n��5���+*��C�On�
���-�w�Ti�X�����ޤ�gPD@�N�ᦚ��� �l �e3=j�L.�YL�k�Unc�S���0c�1ӊ	��gC��sV6��@��"����f *� �Ϟ"{A�L4���6�Q|�!��{YK˱U�q�&8O�x����Tsu+�C�Xn3���okf�%��N���SA�1!���eA��a���Lˢ�H�:��t7z3��M����cv�y��8����v�l�q�j�N]�u��%��H��~9��r���u�W��N�b��i�jm; ��x�R2`�ʊ�L�U�u��[��I�
��87�^ө�zwޱ��)ܟ	�����{br��D1�/e��vǒ�R�fI�z��\c|�AU6�D�����E@����Q���w�1�͗f�q���+��b����u�,�-��tl���@k�����a�5WΎ����������,\�|lҡ���Ӗ������tW���y}S��Uv­���kT.�g[�����u�q�I|�HQ�,�	ͷr��j���4ۄ\R�R|·���yL�n��|��{,8dG��Y
VO��r3�%͎Pw�C��hĮ0_+i񭒵�{U�.��9�=��-��3f(���y�kH(�̍l&&��h�4gO��B�\{o���j�L�	;2S����F�<�ZZa�:�B�uʱ:Lj����ϯ���ƘV�D���u���EŴ�&-�^M�-#1�aW�=��G��k�(�g(�)
F˰ng�ȫĔen4�õv��@�������x������Gg�O���N���S6�ؗgk���z��ʓ-�p���M���ԠD�+ߋ�Cp�7�X���t����v[<��R}��.���`�{z����x̵�$��|����x1��¨4Z�3��:�8�4�jyM[-�EAe�~:�6�׊E6V��)�w?a5i�����FK�y��V�T�r��'FNP5y��<�N'ȉt~����7���PrA�4�����R�.mc�N�֫,�B�O�,��s���Y��7�r�k4�RL�e��㚚�������vIN�K���p��v��]��7b�Z��R��WEDt�_c�0C,2��������}|߯]*K��:���R�)�_C^Ū�`vӪP��� 2G���AX6{)�i�N�?c�z;�KW�L�b��Z��}��������!Y�f�]yѭ�;�5J�5�Y�vl�)��@���	�<`Fc��|��!��[����>|6!��3,�x=wע!t��I�c_�ae�cy�N(��`بO0r񏼮{'��3ص�>q��[�f~N�s���M�"Bas�'���	��K9�����T�D8ncdcC'�ڦz����9�77�����Z�E�3?=�>�����J�aVᚉcl�3.5�����UM!��nQ�B�>E����q'qŴ����%j�DW���]������ز���b�t%���2���~�e�O,��I�n�  aK6�G�eF�c�z�:���_�z�&�	��ڮ��n/��,J�R,="�k�(7����X�켁d��CPJ�w%	�����h�[n�A6���/)n,�U��l��y
xf�l�/D$^)�g��&���J�^����_��*���c+'�G�6 �*�Sb͘=VӍ]MT�ͧ�4��g��7M��.gۭ�֌�t����!���Q��)H!�D5~���t�%Y�I�JHKB��AD���^tȍ�1AY؏U�m	��t��{�6���D�L�������*��{�u������[��Ha�S����I*�C�2�o�+��u�鸘���gd��cZ¼��ɋ���3,������L��/OW��ƙ���W�\9��zIv�$'��j^�<�/�;WK:�ٻB����<	��8��98"��8u5ڋ��u�	��q�0"��H�B�]y�wP�ɖ ���{*�0�CݽMy&�}��ɥ7�=��&mq�X+Z9]t���B:��{6]�&\�{PU�@�Y"�7�7���Y�
S�Z�:D�锟py)�;"�I�@@����	E\!qG�l4-�W�Z��ᄺG�8qW�&-=��A���O����������Oa'x+�`��Ψ��@��:�[��b�"G8�y�RY֞��2�L)q%��l���D��K^�S�4���ݗ�u�k����6q��P���l�q�1��n08�(���iC.ˍ��� �*�#+��( �S�&�kD�d�`��a?���|�&��Y�z@����s��|�{���VN�f�q�M9��(�^�l���e��Z�
�����فXĬ{tM~{�7$�,�g�q��FY�>í3�];�7��f��#�a��p��u=��:�2���K�Oo��M=�uo`7��bW2��I��o"A0r	��BAk\�o��k�k~��;�\i�2woaa��]�O�(3)	�A�Gw�\A�7��dm�[�wjM0o;��+N�4�5�ݺ���0���a��@�C=u���|�ή��ԣ$�v�O����2�T��*l>���������v��%g��=�-$:���+.�ߟH(����C"�\'�H0Vg"^ozܚ�~#6�q��|4�K�k�z�R��e����Dk�c\2�"�=��38���U�ã�Hy
A����k��͢@�y����ӻ��Ȋt�xQ*�cM��\����[^=�F�9�PkU�I��Xm�lk�	<�Y|k˗6ʠ%s6�,$W��(� i+���^F��D��#�@dT<�1���ݍzsM�D�MܑT˄XM�u���'o�i�`��@B##{A3��v���К��/Z�-8�b�����㚩峰��{s��`&��+Ƭi�W1j���r2�On�N��՞J��֞LBW!�>��N<9���T'Y�T���یx�tl���[gbi���ba�²�2J%f3�S�(2Q�Q<Ë�q�����n=S��SBIP��Euv�*i�E���Ki5<�Q��R,f�Rz��%�ym�\�=-��ƴ�[�fw]C����B��:��9���밷�O=�o�5��w�������Ry|�w��ARp{�ş@��2j)��P�����ВI*�豟K�@rq�Y���6%������;�"94+�٘�Py�&F;'��@ʈd�{�����Cȏ$=�������B��-����Ir�.�M������ˀ:�$�zSQo�:���}2jA�"�� �8������k�'�<^×�O�%G7QR���Th=հ�41[��C�8;�f�<�u��zc�'SG>_��Vt@m�|�yY���ڀ7��Չ`�9Unue&vo�h;�O:n! ����:t��j����,Q^J9�l`�Vr�&/Φ�Rl��BK:��f�!�hh��P�����9��X�c��Ʋ��p��$]����cas�F:5����"$�������lp��w(u��E(�Y����2	���4�֝I�� �$.�U޽I������s!�Xc4�4�siʻX@q���n̹��zZSFEU��ʬ�b�3�k�i"�����qp5�uڃ�,D[25���fP���9�{�u�?.Xa�j>��K�ٳ�ɶ��k�8��$%6\6�.��T1:VM�e{�|i�D��vrt?Y^�������Nlӏ>���#�hrt�C0� �i��@�t7,d�V��˄�v_u���r�wP�� ����QL����'@힊���d"qut�]�q��8��5�崨b�n���'zӬue6�I;�:�t㛪C����G����� ��
�RNj����]���l�gZR~E�-5�ld�[�ݫ��y�A9^4������4��m���:����3���wր�ͤf�J��֯Qώ���3lwc��4A��9�篺�!�ꅾ���IR�֯2�C��B��=5���ޭW��4����˞�I�HD*P��Օ/f(�˛��$��Q���2r7t�+auً��VL�K�F��#YDn�7�ys��0*a��n�����c|�y�oV�B>��u��$�Ȝeb8V���wX�Q�w�YY���j	�\�:�WM���^�z�����C������uD�t����)�G��֬ղ3�
�ں8��r%LV�m�c#&���Ʒj8�Yp�-u,ERU��r�Si�r5��a�{m�(Q�8�*������T�W��$יw+z��3��Qq�q��sot�]����MW�����Y�G���*��
t!(�[�V�z3�m28+i�{7_j}�����r�]>����3I��w���^y�<�`��I���΍�e���t����0�ނ�{��^s|�{�~�� 4Y�UY:��q,s,0hL�Yb��!��չ#@��CI��2[X���2��>˩{����B�<���NwV�@�ǖ#��|��C׽gyh�)�ŭk���{�W�y>E�Ӂ\J�B�a��н�E+����[y#���C��˂�̼ޫ+BWb�v7p𵨊�D9C+�q�AlK�� )\�wFL���4���I7c��ը-��{2L팈�5ei:�>=5y\�"������%Ğ�{��fn��7�:�l��ĳ|J�'��;wV�Sٹ#�:�a��c��n)�-=]׍#���ȟ�ֻ��ww��A��F\��k�չ֡�tL�����z��;\� `{�5\�����x<�w�-�/7)�|= S�PЇi\^>>�.n�^@|r�sq����+J��N���@�P[q�.���;��c�oY���a��v8�sgbE9A��ݽ�Y�eᬎ���0��*lh�t����u�yN=ytQYA�.���snV'2��ڳ�ju���6ң}E̋��ǹ]�_&8�C=�����74��մ����Qݥ�@��ŧC��O��u{SY�k&.�+���|�=e/�>�g�*֔�������<�gvKf��&Jxum�_�������h�߹�����w;�w��O�k��4;"�J.���z�}|�!�jrp)�FEnee�Q5ANX�eQTTUL㯧������}>��ǌσ�(+�̌V�#'#,���&��22ƨ�"���"�j�*�3'����o��������a�ɼ�����¢�"�����0��
���1�/,�Z�0�*!�Lq��Ƿ�������>>3=���*)(���#((�$�"�(�& ��
j�(��[�F1M5=Y13QNUUUu�LQ�e��؈���*/K��1Ce���6eeFY��QA�MVfTD�5!�QEUSQ�!Ff5T4SMU0P�AA�^� ���*��"�ȳ,�̈���ȫ Ȧ"(���0������Ȝ,����*�B����'12*%�,���j����(��,�J�h��"""�������0�d�����*"�1Ȫj�����j&������3""%����]7��΃+����!��&rj�ue7���{<��+3;���8%���j[�Ճ��#�<G� ����m�cCtCb�ě��R��R����mA�\z�\S�*�8a��(L��+"���%�w#}���ib1�&j�	N����[�����vG}�0����TI�e;�k:�'��+���{\�n�q��n7�@��u��ƀ��,$%��G0�m���z,h��Z���D�]t�s�>ЫΓ⨤�=C�A����j�QF�Y�-��d��Ej�bA��[q��6��G��A���Yu�9�JO~Jr�b��g^(�0���e>ko)������h<��S=9�(w{�]�.cJ�Yj3�	��{6���/P.L" �毕iVr��k��7r�,v�5��<��\!����/�8�n��A�6f:39�/��ش���(v	#Y*���qju�K���Ш�pR כ�D.;P)��y��+Y9uG}�z6O�<�b_���wgaDv7��b��_�e9�Ԗx�����#�~������x����`_�$}�N5�Rj]Y��qp�S��Xe��t�sg�@���i��8��ʚ�S�&�Ʊ����?x����c�ӎd]�_��<-���q�>������ݟx�C���+����njcc:<����cUA�������޾S�,ںQ)weK�^�ʐ��	'+����� ��$F1����Be#�ĞF��I�\��W~��y���c0��p�����r�O*����Q�zO>,�H�S��-���
���q��T(�Y$���7w,�G��{'����D2��Hpr�P����]^�Ű��u�д5�K�,Ls�
@�슍��0�^u�Գ` H"���@��b��������t��+�����#V��k�T����.��z�9�mMX4;7a6��\-:W����\����9�uԊ��!���[���p>�w�v�~O�wO� �G������_�O~����'�w��-��2��z���ۉSӘ�]k��x��̂��t58�m�`CV��w��w���T��DY�'Z�	n}19�M�����u���/`ہY��s��n7��7Y�e��]ӳ&XQ!�܂���Yv�ת�z�;8�ʽ�g��"�(ׄ�׮���yO�nE{�W�ⲙ@sOQ�{��T�ޑ|�gӞ^q��\21������mo�1.�Z��#x�^�ȣv�0�^꧁�q��m���Ǝ�ze&�k�X5f=e��.�a�ΠMz��኷|�]rڅ|����G��Z������m���C�*������Ǖc	L���Ĉ�����e��ۣ����Y�;r�GQ(m�~�ۅ�A��ٵz�߲��=L����rlESsY���@����қ+ec�J	�c���&ʓ.��͠F���F���ڳ���M��g���,²ʬɺ�2κ���>�a�G�b<H�����ލ�H�A(v���y�������WJFq*��-��.�kץ�2�t�,���4�.V)ѕ|���`�5T��|QR��G6pH���,��p��j�s�\�m�㚺[{��
o Ơ��2};;	�����"�	q[�~�DH����:�^�i6p�D�$r���9���oT�����:��Ã�ZuT�=�3M
�v�%Ō���?s�J8��6j,�'*���ƫ�����e�j�.�dG�0�Wv�P9�M�z�y��r��@��]aF�uL�qv����W��x�L,��Yx�uy���M2i����%�oAky�o\;m�[��j{KB��A��2C�����B %h�1���V"��zEx������������˞�Ip�`Im�qr�jK^�i���'��RԽRk�njՠx�[?#K����X�ǜ��`�ͥ:y�h 7�g*�0�RX	�|�>�N��,4o4o� -˱�Z%����=�K�Cn���nM(���z녕 �\�md�+|����`\g=$l:"-�۾�E��E�$we�|1x��K"D��k�Ou�h����ɣm�ЃC6�=B�e�\�pPJ�\����H9l�t��=�j��4�X�L��Wqt��M>Hy�x�:����3��x�<��鬘��1e3Mü�p���B �>�/{͚�AC�9kijKC�/,�)�z��ɀ�5�]�X�)�u�Y��ק���s���uҡ7�aA)2MsA�A�>0�K�ao??D��u>�==f�O�?��;y���C?��=�2��6��Ӭ��\,��LaŅĔOd�Ҡ���8�Vώ�R�,�x��QUL��9M����y��M2�h ��8�ÏY�XC�I�:Xn���1��V㶼s�	*����n��Z�`�6C�3Y�D[BM�����O�7�do\�����c7�z���Vk>�Z9Y�7�o7JÏ�m�.��	��B��q.SS���VMiw��Iy2I1����K)�I��Y�K k֤���tЊ�*�=��e��F��Q�}^0w�taE�r|�̦�\����b!ic��q�[$f0T)��N5�>�<�l�����z�EKݺ��	��7��5���p�f��F�1�Np�����.2|c����sT'5v��
�_Ļn=�\>�v�8����}E���5����u����Ƌe9�[����LJAs�鳍%vX�1�і��6�G�BW�r�V���aܹW�P��t��P�k�F�C�y�֖�a��:ď���9X��J��T�Z�b���OC�%n)ӱ:M�4
ځ�+��A��|z�Hx��g��/'�O?�W|��o-��"=^|ɂ�2�!n�\�D�H��6[�=�����1�}�}۔[�u����t�|�}dl��h��i�sH��m��֐Q�fF�bk�:Lu��,��`g{��`:��H��Q�{P.q0j�4�`,�@����l[!P�]t\H��|��1%�T��jҙAΰ)��n����p����f�"�.�&[D4�9H�K=�֛�B�J)֦&�j�T��7��=�(;=��5��e�e��y�V�Du(2�
i�9�&:Iu����%�q ��jL�5BW�<˩R����SS��a{�T��/�DʕI��Y�3u��J�t)�ɬ���Kj��]�*��q��=�^JL�;5���(W��v�_zq�R���յ�MLo`kB�\�l�su*=��{r~W<��N����)�w=�#��G�oK>vE��P�br7�KK����D��hc^(�q��J�l:P��R+2Ӄ���+��{�8:�}N�KD�=�=Ɋ�`4Fm0�-c��a58��n����_��}�J�3{�en�	����f�5��JihQ���ԊJm�hV��� ᮢ�f����.�C8~��V��њ`8%��0��s�7_;��՛��,�|��+5�{��y7H���K{��x�t�b���ׇo���)�x�
]��0��FeKsE���_�3��p�5"�~�}^h����2��A��E��8�~ŵ�I��$��=I�l�6L�V�%;�M��G/�!i3*!����!�v&<se�b�<��V��V`�d�uM�x��Yܕ��)�X(�d��� X�M�61�D/F@`�<����-S��ڞh,��G�+.V�J�R�$�Ufm&ݝ�p�o@�Ϯ��0���k����f�X�L��wK���.s���i�;K�F1���L��������!M68W؋ n�KMxV��p��7`z"oV���C���&5�ƃ�Ү��\MG�,+0�l�>�x�E�4p��I���P����Ù�b',�mq�ji����R��Ǚ���w�����O9s6�I���?^�M����z04��:M�n	^>�A�?<���%{9�P^@L2.�<��(���s��b��J|{�̈́ڍ��K�L�(������\�*_>� �{�`��T{�ߥfF�!+�K�q���u���x���^��3�ɖض��,%�o3tT��M��fx��OS9t��F]E�n8��i�sHG �|������IK�eq�:W���� ��v��7.��S��!�\ur�Ž&�y�Y]�V�9q��&���CB2�z`׼�W��Dx��`����<<����g{wzp� D��
a14�
���f�,5ugE�Ab�;y�w |%��@���6޳!2��0�h��Y~�X�,���uC�ɮ�ug��uR�5���t���kqmܜR���q���S?=�a�O��(m9�.��0��_D����Gz%��Zz>�d��,ZJ�S��;#� ��O�))wx;���U\�:'�����	T�u��Y�f��7��f4{t{EJhK-Շ�,�Ξk����#ǟ��gg,^�D�_�aR�*)�G�Q�^[j)s ����Q� tR��k�U ��0G�Kq|*Sv�%�9�����}�N�K�m�g��4ْ�VN٭���\�B�ȑf8��%���%FK"�9���O��&�;
&�<�O?J�q�|��n�+�x34�Wk(Cz�Ol���B�����Gs�������u��덞�4����yҭQ�g3U�K ��=	����yd�޼IP�&z.(�ċ�_:7� \#����qM$��d�,�G����-��86�C�3�%��v��T����&�z�I�}O���HD���ukNwVJ��=� Q�%�C��ǩ��?�	�Q)z
�~��t�$rԻ;��}���ݱ���Q�RT�.mr�5��4�g[�q�կ�.cv1r����脸
�����Siҕ��?;��@ڞ>����`<�|G4��d���ߦ}k��I+����#6�`���DG��5�j�G��y
Oh��ݘ�ϊ=�:����%�#	������3�B�yD3F&)�C0�09�ߞ������q�/Xؙgy�a:��2Ȱ̂�Z�D�Z�*m�H�6кޟLF�;�d YR�Y�lZ��ӱSV�!�zj-dcYr!�c�0�� A�"E8�yH.�tD�|��e���5�!�	}G;�g:1��P�_�a���/����%4�&Bm�q���}[��9��a���F��B�vd��)$��R��Hz0�-Sp8�{�4ת��f�X���D*͇�2�p) T�{h��kv�mɾN)��(;�M B�U�q��q�{�ӎ����әأ��2�����#x���p;�(��j�a$S�;BA{MH��	���(덖d�^��ʭ��&��D͕\�Jt���ݼUm��F�5�*1�INC��"rᆎ���YYW�Ͷg%��c�Mv�0����@���ݎ�O����J���aR��Y�_��r�j�Hs�3�����8oR�!o��^�H���!�ޓ�M�t��j.:�M���5��5��������H��k�%���.7�>��n�`�W=Fp�a0bVu��ݽ·�X:{t\l�f_S]��x���k�%��a��b�T�3{Zm��*��r2"A*�����췃���$6�B�7�tֆ�b捥͌)��CX�"|��o�ڎ�,�#[������Rz��� �m.��&����ssFTM�%[�a@φ9_�F���r�O/<c�JT����^�(TL_b���j
*��H=:���.؈4m�9(��p��w(u��P��l����6���U�aT��3�.@��jad�QW��"L�qO<�v��2����e��-�A�7qNkwbtD��|e��m�m�^؎NO@���^�;؊�SZM��G�I��	�����a5��c3S�P<�������v���º��w��ջcer�e�
�-A�������SQڦ������`F�X9�,I5�Els�D�xyI���ŋ�&a�[HO�酊 Ē�p�=�
XAp����"`z�q������.L˫V��3l.�0���q����M��g5}.��v��l.��v��ܜD
a\;
ԅl�Z�U���&e]s��Q�+E�����9J������7����˭��:R����vώOuª��@W��(��1��~U�J�����WlT�^�Ǭ ��k9�t��I/.���*¨7/b|v�v,q[:�`����d!+������`;'/X�Ẋ�A�����u���*��p��Jcd�ĭ��J�!�QeӇ6v5'���[�:��c�:e�،��AށM�M�X^���1)Z�����6�حƱu
��4e�����m*8{͚�k��TEj�A��rz ,J"�}J����t���^���xЪ/��W[*��⤆����5�,���z|I���=�V�;ZuG(��@]�da�6�e�$%���,�����rQ[�G�h8\	Lx����b�yH�e�2�m[��#Z�"���!?��сσY��r!����$�0�+�c�L3��`G;]����qJ�>΢q���>í��T6�0;���oG�iJAb�VK����74�}������J���0Eʸy�B�4^��9�/E��:z9o�����e+�	�tŨ�g�s������7��N��v��Q���dN�~��Ū�5=!��V���^\��*��Dzz�V56t��I}*5"� :���ׯ�"}� z�1����'�?��F�_�����>�d�oEGi�
��l�ɪ�&�ù)���.�i�/C394Ȑ������p�$r���̃ ]��Ác�լ��y<t�p՗B���M��|�G�m�����N�m`��������rOk�����G��@�$9�s66Ō`�-�֭4��f��_nu�b��g/%Nr�E�+!{�Vb���ǹ�T�q��y��Y}�Z<hC�r�v.|́T��6m*{A�w�J��/Xz*;��S,�Ϭ>�^�_d�K��$u� �έ��C��;��Rg7����n��c{���GK4�Cr^9�:�Z�Ӯ�p�r��G]'�����e�r��S W� 7啇�~U���)�Cuz�g����#.��\�D��l.1X�CA^�ĤBܭ��%�ݫ�>g����� d�C��V�*yH�T@�;�2^�&�t�%`6o��z{��^��������㑟\����Ӈ�%��g>��o���\x�±�y�nJ���O��N�נ� �j�U�d�4��˽}g��T`�|[�{>��sC���{��&��J��2���=��׳LpB�^x���5\ȳ�P�u5�E�U�"���ʛK'������L�
:��G�h�s%�mt��p�U��vzײ��Z�N0��#S��wa���E�>WO\m�w��.BBj�,0e
��7كNa���ix	˰0r䊦�xxm���y��r����Hq��^��	aI�m��j�&�q(�;e^og\�uMU�;F�:������V[�o:�qo�7i�q۹}���$s�IkŮ�3�S���tf.��t2L��l���&R��N' ���.U��W�JM�)��Ìޅ���>�q������su؈�ʈs��5���oU�5�Xv\�0�U���c!�6{^�VOC�ݣ6�8�C9���;���dAu��D7�C�.�s�N�0�nD�Y��U�B���1���S@�D�oD���N��~5Q�S�LY��p��F�\Y[��*�fH�mYt(:J�=c6eͅ띜B����Q8r�eT�=�s%]q�Y����C^�<��k\�fcc��gQ�Z�"ҍb�͗N�J�4�;�+� ���E��{������۩�iš����?�� �^:�J7ܷ}��Y%��Ùs���R��^{�u����}H&P�y-�tE�:������Ű3���(��d�ҝ/�Cf�R�&
Þ�D��l�Od���z�`��GɁ�EO7�✝�v9��Q�]5�]��`�����h��F�ǃf^���팍��)a�݆��M�U7�rՉ�Zh�%��Y�#F��� b����]���Kp.wң�)��2�F�<m��m�'������EI�~����8 �Ra�I��HU�CDB�MH\51��e%B�� �p��A6�����>�Y.��սz6�QS�3Ք�L�UQTčS��UMR�DE����̶ɦ���zz}�����o�������y�CUS2L�U�]�����+0��,�
)h�
)���u����������>>3=�<NxQ�P��DIQ�T�U�XA�F0DV�㯏�OOOOO��������(���feE3Q3R�I�r(���(�(b+��70j��)�,#*��� ����',&�"�̣�� ���)��	,�2(� �����/F�4la4�1�70��]p̒�s��ɦ*��Š") �(&���
h�L�����s��h�*�r704���(�,bi���"&,�((*�$��)Ƣ��������f`VKI�41LKfFeUQ��E,�QCS��fM,P��%��QB��5ڝ�G�)��]�y�*j�AQ�%U��PyO^]���Y}	Y���7��	T�j���W[��姫-�
�����έ�C񾤅r���HKڥxh}|jִ��i����\�ji����X�9<�@z3Mcom�o=u��o��I��	�@���Z
��}L,��p���C�܈���V��)�r�;jq�Վ� ��kl�m�Ҏ��K��\f�����g�'��N�T��n�GN0j͑�5���t�]����w��c��d����f�sQ|��q���q���m�{/#4������k�Y���%D^\
��z/L/�ո�2��Y�Mʡ�/T�	n�#�2�&�.CV���^��4o�*�y�3���[C��
���-ekG+��rm��:�v�KW(���a>��n�|�P!�Ǚl ����z:n�����T�g ��[!S�������K�7��b���@᯷���Tט0[�F-�Olۊun[��/y�"�d��0���@����qh�A�(�/,�Y��j�u�cca晣�N���=i�ذk��̩��:Q�<����i�I�oc��+#H�v�j�h~�"�Ѷ=��0H�:Ьzt�8�id�a��Z9X!8%i5�9��x�q�X�����L>G��ʜ����2�hj��J�}�R~|H�JT�{/y�<��γ�߾���#o8�=b�����f�5��3[١���������>�LɖW�׵d{��\�/��� :P��vN�9�=Zm�:��}@٧��ަ<a�ޘ���dV�JD�1�P�7g���}=��Dr�y�J��r����m�M�tI�PZ���LDq~���dM�.*�˧��w8�JK
�7)ۙK�����WI�-�m���HI.
���o��s���}ZA��Y1�p��ڲV�ų��d���4�a����Ǜ����Q ߰^��m.q�y��CED���~40Q�˞�#�#g� �ܓ�r����/�C�'e�f(���!���7;S�NZ�䞀گ5��e��FC���O8|b5Ҽ���o_�OL��6-]�fr��Ӵ:lG*M(�x�:h0m�gr��o��18ۢ�I�#x�b��Of����q��j�7�Y���^������|�r!�ݓ������]z��]!��V��9��@ ��|g��9|������DX�k�C��g��{g�;WО<����?��\�MXo��ɹ����1�s �k5�d�Еs_ܤ}�.���g�������X��'#��t����2(��=���Cv�!���8��_m^�@+j�z���kY+4Q8xF�f+z� 8t=��yWu��(�"�ns�n�ω[��ה���sp�NRFe�vnk=�3�e�V����T�V�䛵If<�g�]�5Ӧ��[�M˳��Cv+�Rx�+w
��>��KT��WF�����;}=���^z�+�#���U��_sF���w���T���m��O�����c똲������W�f|-@���Cb�@��>�E��Pd��=E�>sŗ37���4�f��*��9�k\2��t�~�i�]�'��WV�kg���xo#D�:��9"�����M�!�?�k.7�W�v�Ș�2������n*��sݴw��ci��DS	���E�G��N0�Ȋ�S.��h��@�f� أ!�n��>���&�܃9�7 �"�6_,˄���f��&�c��J3=��2.o%/l6���J���Ѱ�1U�8M�E��zb�{:�]j�=q0MKZ��=���zt��tQ��We2��3J?�����\�>揼]���{3��+Y���w��C�M5frY��=����c�n0�$p��������s��^a��W�C��oG=C�h���qn�����\|J=-�n{+�-�%���ln#u�����rA1��Z�!�W��9�>�d�}������Ϫyf�	��BB�k4�rJ�ࠦ�wt�\X� ���)k5v�Ր�azzZ��N�D���h|�+�t�kku�Gk�Pڐ��HF.G�S)�6��/�k�n�L���f7��1
F�(��/9A�7[9���yϒ��5^�At�2��79^]N�WI��y�zh�CX��N]�����Qz5�&�ٖ!�jK���mY���V�Y`L�+lD��ü5�4H�h� શJxd���9Ҽ%�u�&�C�Q�Y�f��/{�I��O߭�Nᐶ��\w��#@m���Eo�9
�u]6`�q⮦�ҽ���3���'h>��+�F�
wg���S��Ӽ:7gP�=�c�RF��ݐQ��s��������ޥ��ڊ�c��![�M�,U%usEͅ>@8r���oۉ`�~���p2�`�!]WG�,���R)���?��ϲ��ߴv_�-����[����D��Ï:��o��i�l|��VVu>|��d�%@e���{�����f��#�]h�gZ�v�c�ށ�bEfꊻ�B�bB��a�^e���^D����~\�-�rV�qgH����q{�\Mv��뤒��[�zЭ���a�+ܕ7��crq�Bh�mh�=:DE�P��@��O,���{�8�˓�r��5��b`U��kw	���l�L��d\�|1�®��N_�6�����BL���W]�+�3l��׵0��.hl,u��db�m7=�����x��( *P�����Ύ��0V�B�bp�8�;���9=�S)��]��sn�`�2M��x��^W������:���/���!Y�D�'��&�mM�ݹa?�Ɲ�
�j tqo/>���Տn'u/j矧VFo�V�p#�=�իՔ�O|U+��e��(�����(j�hF� �k)�S�n�����%�X5��Ŋi��R�Q1���5z����VT�H������5;L<VU��i�Iv9��6.��Ĩ�|u5��V��51�7���3��������@,���s���$MPZ��n��3�$/v���[��>��b��w/^���ۉ���ي��E!T��Nث�;�6�A ���� ����љ*-]�V�]*�G�����V�"b��`�V��r�c�_M�eS�<�Yw҇E�>�����Vû[�������ȎU!�Jø�0��Y����}�s9��[j�Ҋ61Vϣ�_�e?�NÙB�����u@S+c�zt+;�{ו��y%��hi�RزU��ǯ^%[�B>^j���YT+^.¥�p��Vkg�'x���)��#k�"����P'���<�mѥ�}$s�L.�Y�l�ɬY�9Եig�I�'۷�_X�z	�?�%���e��R&c���LwR��[�t{� ���N(��
�ާՒrX����4�|ڛ��"5g��gey`ƦP)��΅U�}EV=�f��nA�np��tqh�bS�}"�)�B�֍kwç8|�Mq���t;�\,��k_��m�s ��/dUTe�u����4�	B�Z7o'^�{lg���_�������Ƕ����Ǉi3����|4C��q����X�\ �'D�c=q�����ӱ���ԝ���șd��"��}�4�c�vWpyE�&�E����X��@��M���p��;���q@7D%��Du�^f�e�g�xTZ�>���>����="��v՘V�+��>� u�q��s�-�������Bk��ᠳЫW	��t/��}Y��rCQB̊���^�{�ǚX��1�n
��`��1�#ú�S�C ��#��:k�����wS`�N���g�U1ۇR�ٴ"s��>$+j!Q��u������ޯޖ�$0�/�~���4c��6����ݘ/��*�ε����%�=��$u]U���3q�n*5YK�PW��۽	bP�e��꣦�ׯH���, �&���g:����,�O�#I�9��� L��f{f�u&�g9P�����kW�����Ǥ58��~p%sNb�k���21:rA���"�13I�������8A����Z-\�َ�1+zo�y�N��[Iӱ��0�u�:r��9V"Y�r����'�zlR�jꆑ����ɲ��70�3��3����4�V%��߈i��_/)������a��otj*W~���u�xPC[vG�pN�,|||eD�}�g+\6<��Y����&��jl�yegFa�ф�*2k����eDc �e��¸��-��k:C4s^<�����ӊ���6�Ew8�kg���O�"V�T��j�>�h�ˠ:&b5*S����Z�&��Yۓ�\���Ӷ;y�����EO��{ ?l�� �c����_�]TF�:� "�[�1�n9�^�®����u���� wP^X�=YN���H.s�&��چ��a�!��a�.Ҝ��q���hi0N�0�P�x����7�k6W�s}|�����Ϝ`Y�~�zE�]�y��wv!J^�◿��<�]]��(o�p��ɯ���pg�dѝwn�E�ku>��l��:[E�}�N�Y%[4m��&X�{s/
s���Чy���6M���X��^���1s��J6�-`zp�M�2k�D����#��r���P�T��N-� C�Y+nz�V+)�c��w�&C8���;p.h�a��mo`�W>�KhY��,��fB��Q�\��)��G<��e�Z�!�V���sf��;���Tֻo�ů���62���W�C*Af<��մH���)��U�ȴө��M����{8u���}��pS�wGj26�*��&�W`T�R��)�=Oʆ����]tSK����!p��k���?.���^�J��0�M�Na�0F ��Dx� ��*ָ��E��
yE3�A�Z`B�Gu��ؓ�~�
n��?:W��L9���T[��i��!�IW���,l�wd]*框����[���E����F���n�-yx��ӱ2���Z�)�=j(#^�M襎F�KqcA"ǚ�U?mt��˘;��Y�}�~��]���JW>��"�p:�sV���s�쾺�w���LG�F)�9�Ҕ������Ь�7�� m�L�93��������o���n�}>y7�����Q����.�>��cP�V��7�]��i��S�B;vᨒO.ا��oUWԲ�#n�P���*�m3��m��G-�}���h���,u\����������{�чǴ唎�*J�]4�#1��մf�����,2Y'�}"Y���F�T�ɋ�X1�=��o{��̤���\BD
be�t6�}`�~�Ӛ��lJ��,T<����iH��e"�+sg�("�����x�a���M4n��+��~����\f�V$$�|(��q�d��[mS�����WW��(�1Zs��gWt�9��:.T�2[z8�̷�O�F�������<������Nf>�.S4���|��g�r��	k
��i�X97)������)Q�7��j?�G��g돾��Z�^��3�5c4#M��WxxD^v��R,���:1��V��=3�R��O��� ^m�+:�0R�}�MvX���lxL�#�ꎫ��Wc(>��W�ϯ��Q��d�ҽf"�m"OuV՞�f�1�Q@[j��}Waɹ�������;��N�&؛k^F;�IԖ�����j���А��9d�[t����Vlw>�h쨛xx�����⩀�;���lt�ݿ�U��3Ms��{W�zsj�r-	rsK���*0i�|�h�J{��2��n��mP�<h[��TՇ]�{����\�ooO��zҁv{��j��ux�=0��w'�eƩ�ޭɢ"^c=Cx&��v��uOlZ3:��d}�ca��+�;	�Ǘ�q^:�-]�*n6���I�g��yܾk�s��g�7ä����й6�VL7Hi�Yq>�����R�v�=��𰈦�!� ۰��]fQh%P�PU�Y�|�挋E��p��2VQ�]]�ͱ����@\�0�o��-�f�)P�P�̓����E��s޼%�;w�HG�Z�'-�fMOQ��U�W��{��,��F9d5"#�f�9wAI�<�au%:����6s�]kh�f���
p�!g2um�����9�[�ڇ�Ĭ^|{�T �h��ǟ����[��8��v
j�.ae�pV��stK�9`�4�Β�B�'Oz�O�i�3$�Na��K��j��?��Q{v�Pe\%[��}��'+�e9B���%0V�-hI�1Y"�)���R@��Oܥ�sya74X�C�O�������̯\�p];1֌��Ro��m�2V�T�mwo[n��@Lj�Q��[S`z����n<�@�S`�t���oB�ٴf���}�bvk8�J�����NTqׄi�5�ۚ~Pq�ą�j�ÆuL�g�t﷿~��c����R�/�h$r�4G�B��.��h*={؆j���ꧏ.n?�#5�fF����5T31�m�n˭{9m��-"�mS9�K��W����Y�t7����)m��<'t��d޸5�IU�$�����"�k2�D�o�Q���I��Og�E�-�v���.�
r��b���� ��R��K�v렐�'[�i�!V�"-�f����Vh���rg��β�V_�KB�4F��c%�2��(�̏�u�p΃�Ic�3�` *Ku��z)��oh.��c���tk+q:�w��V���k	�<*}پS���Jޗ��#��sD��5�7}D규z�[��e�s^�|vf8�W�PűAq�0��#u�ɤ2)D&<U63m�VB�4���hh.������5J�q�qI�:荬��t���S,�h>e^�J���������Y;�K��9�Z�,��OF1�o���|Y�\�uk�[�&.X�[��T��Ӈ�֗�6	n���6��1Tn%�e��6To0��v�k�|�qh��='��M��`ӹ6M�ߦk��F�U�u��{�w�)ߍ9�S| sq�k���:�н�V9j㵢�\FnL�����9���i8:�]��a����3���B�W�޺I]K
SJ��o_e?�ұ��Cޮ�x����]����v�vN.b<N��j��:a��-��qu�"�)���od8Ug?��\W����fP�2=ji�-p��w0����5k/���i�7))Wc�
t�(Ӑ��A�]�E�L�՜5cܨ�� "�����rIvj}kH�z�u�\��ggd��=W���,]w��kW`��+2�&��u���)��GƂ��M=�M�链8g%��R�E���
�7p+��7.Y��L�aY�a�R�AݑUQ�E���َQ%�㎼{zzzzz~ߏ���O�%�ʺ3
-��nY���MI@P卶CE�E9��YcUPV`e�O�OOOOO�������񊣑�FY͑�Qfd49dy��EUDD�L��S��:��������||��r�������MNfC�P�M1DD1�9%STQD�T�ADMS@UQfeQTD�g��KD�!E��v)*�**��
�� �!��¢*��"� ����Bl��b�jJ
*(��Z���¡���)*"���2ʬ�%����jc!0�"���������220f��%"���#r��((*�=�MS �QL�IT5ACEP]F]�z܉(���$�ꬊbh*&���)��a��R�4PU1��������y˯�z9�׼�\�!u'4{�"�����|h�;�L�mI��8n��1�]��4tte��D��_6vH~l�6G��{7ƈ�|�'����*�=�����^���h�t,���6Tc��*)�|����DE�dw+sG��'�/ߍ=��F{��q͏��m{�x����ƫ:=y���J�9-�_q��?��jލ8Ќt`wa�s%j����b�kXNsți�a*/&����޴gH����`P�/1sx��#�v��x��",�Cg��}�e�@ފ=ti7����^�R�Y�����4��������Ւ�ZLH�=R� K�T��,����mlޝ��ƺ���S\��eUx���5����k#J�}3��z6 '��,2r��h����F^��K�S\k"E�Έ�.���':�Lgr�y�\�k�mm�U����d����T�Q����G03���um�I��ܷ*}В��mY�F�`�c�S���A�%���R����ͨϮ�e��Ni����X�:Z�2{!��{�4��n{ą��\����k��<��pe����i�2ds�Ύ���P9����@�q�R-�>x���C�j�{>F���z�b�i�*�n�Qh�m�C�~r���JO�3/�Äu0[��K���%J��<��w���ҧ���hx�c�کA��8��[5� ��Ի��X��=!f��q��P�SJڄ�CK�ڋ��/��&v������d&Q��`ܧ9��.�Ȼ�>\U�ձ���T�ޒ��NN����;�������BcZŪ:&��=�����긚~�����)#�S�}%�q�p�˅���/$5׭a���+��A+��z�ʹx笿z����r*z�<��:��E�C���ď��R�<x���~]C���Lz�s=$ӊ��a��M�ލ���n�"�xC�i�E�F�1��k�+j�����ʀ-a�ƻ'"a�
z+r"���a �_���ycz�
CQ�9��������W�[���ٝw7�D����F�G�a��˦<���+��%鉳UfyqӸ�.-�\�����w~��qz�I��fi�������3��ӌ�^���5"<�k����wg2���:+�֙��u�б�	FB�v{Ծ1o*�ݷ}�:�mɒ.��r9M��k �L�
�V=c��':ќNc�/,���wsES�]6��u �;vK~F�zBa	�!A"$���1�>9rbu=��Ѫ0���x>enf	�~���ɦS�>O��L_.�6T��1܅��3Kٹ>� �,��Q���gԧ��khU���ݞ#_���p�*��ڂ��!ċ2����V�e5��D�D��(�U�O�4G�6��|._���V�v������j��kkE�MT�o8�%|kW*l��Y2X{�n��lI����t㋲8�n�&��샜E���s-3�\r�ݭ�o�@;�.�s�"����݌�E�=[���yTL�gF��R�a��������`gD�o`��MV��y�fC�=.1�̯�zvt7;�����Ѥ�\��
7�Y�7��[���S��v��D<����@Ph4&�UZ���*���oU�R��o�=hVN�S�GW
�֥m����|�LZS����}Z�oo�����^�JmNfE
��j�:z0,�:��؄�Δ]�+��uNsZ�t:�3=�RqX�wW]MS�˅��:'iv�������c��S�Tc:�7��{oiݎ�81P�ܠ�(	��vN���DS9�K2�w<ǓF<7��k,۹%���-u�����{5�� F�x����r>��(�;��Q���)���6�w]��_�������j��Gsxb�62��\��םi�.�̐��6Z�s�i�a]�I�@�����5���қ����P��MT�5����iݾk�
z;kD.7����N���9\:��4�ʭ� UvM�����z�2[&��r��FOsX�)b�XV�μxC���_�6�N�|�������Ҫ���k�ju!�T^Xͷ�J�7�-NPC 4C����>�i�X��ǎ�����F�(,צ���zYY����>�j�;�"vi�	�~]P��ԕ���KV����srnsxY���);KW��^̪q�ow�X�l	D`Ci��B<���;�����U4^^�lI�L����sE+�F�����e�[d�*��{Oِ쒴 �6A������r�������9�����x���^�s��:K*;ۜ�ݗ��[�t��_V
�DV�X�'��s��s�ɒ)�]ʚ��L
u�|#w�轝S��k,>�^<��$^VҨ���v�a7Ѝ�<�^m�[�+��o���pi��d�����l1��]�ӘO>������;��xqh�VY�C�E�Kg$���G����Ź�q6��k�#c�<ɓ(4'|�]�y�dG��o^A�IW?��u��d���ڼ���M�4V��eb��CF_�7oO���.��Z3:��f[�s0�5S��E�"�@���gov���l�̀���i���=����Ga�٭}ݱoey-9���A����- ��p�,o��+�ܩ��n����t�S�^2`۶ҳxܒ^�P���Yx ���ī�b_�6��A�9��f//FY����z6�Y�7j��ۂyF��tF����P�^[�F�B�`k[�+�D�N0��ޭ�b�� @�2��Sjjǈ���h|�$8b���'�h܂�����n���N!TU�;׫ŮTK�;�Lб ��59d���f��Mgf�K!���~����C���rY|�@ۗr�m�ϝ��O��uV��^�ȳa�~~��}�'��Y�@���s�/�2�fٙ��-�Ob��,���1�S+�������y�a$�Cc�Ml9��m�p*�/�[�=�q��ln�8��W`謬��������I���u2��ٵf�K3fzw5���2蔔�����>S���1.�"�F5���E�K�̪[��Al5/\m��Lv����c�.��z�n�b�rxt%�S��O�䝻�$�o���˻6]��c�4�+Z0��a�j]�႖��vClrV�|NyMn5�s9�jټ)�z���d��o�zR�Cvk���R�m;�}�/t��5�Tc�b3���Ԥ�ԕv�E���ܽ��[1���$6�vl�nOb�3���5��)̻E����;�%dux�8}��؇ޑ���Oi�]�:;�CU��y�iZ�i8�+i��6C�vZzn��m몃���=�:�KŐ����3��UoV:���ݶ٦3ƺ��&V"=�xqI��n��}��B0Z���P�|�=
��6Q��|_ہn��P
�N>��>��ի��V"���aTy��j��wȟ=���K���rn����/n����$	ܷ)kqp���bS�|:���~�g{��݂��~��؎}��^���3��9b�� ����m��?#�T��7�u؟���P�E�=w*�v��K��Q$7�� �u�=vb�<a��P��ƠƧ�r�Y��k���9c$2�{,�9���t��U`���u-��)V[��l#��x�[�sPbO�G��_�\�#YC���ޭ`,B�x�O�H��owEd{�M���{jW�g��Tm��J�h�)��Y��5#���;Qوi5��"[��S�Tch/)0������m�:Z�?>*�Ezy�DNz�hi�C�ǥy)�Z���e!����l��p���ˡt��J�P���ws�LV��1&|񬞤�R/{�MԴ
�'OU]?���U�Vh3@%��A>�ޚ�v�D��:��W.q0��p�K�<'gm��ǚ�_7B{���I�f�EZޤs�Jf�����|�&�A���foc�P�uƳ�1m̂܅@Gu��E��،�u��`�4�iO�u<��Y�t�(UY�ͼ�}͍�li,�t�Ad$9^ڙ���<�v��NQ�3�=l	������Ov��͇rW`Un�pМ+Z�����a��+%��,_諾�w���+�݂����{#&�����@lq	n;�=����f���D�a�!v��E�Y����n %�� �/��ɰq�ž#J��v�C��;q��]��Z�z7��f�\��J��c�N"�1���=X��;�����ՙ�6)W;�rK��]Y^����w8�Gl��4����^��Ifi�;�0�v�j;Q���R���W�t�V�Ӻ�"%q	kl�ӳ�i���0����qa��*�I�i��H��a&�\��5%�x33Q�h;2���r��oƬϜÊHáƻ$��|��L��N�Y�3���fƞS[5����-�����A���l��W+�N�̭Ʒ�Ť�Oc��Q6����+-�ק5t� B4ӫ�1�z	�뼱5�C���k]�3Y/Ղ�@�-��H�&'�`�����2w���g�n��@�bb4�>�`u�t�g��=fr���P�!�5>��I0ͼ��d�3�+7�J
 �݉�)�_nq��Ym�,;��
[6q�bpx��/q{���}fC�!t`��^�I%��xp�c����4=B�e����Po�ƚ@]L�8S��lv��B��H�7)�x~�̩��ڞF&��[�h�����c�c3�W��~��H��vwj���3�^�/x'9iՆVеxVz�xȋ��n5��l)!U*�
U���W����1�rg�O��b��W}��8�"�E��E*�V�*���Ӱ�Bf�Ч)����5�^v��Ķ�&��[�Цާ���Օ��V�0��s35�f��$�%wLx�kt���wf��[ݨ�v�6w��BB< �p�'ѫ{��-���ҹ����V��=Gx]C��s�Gpā��l���eg�V��|�Ok��V9�3yܝ�z�/h�m��1e�c��`�APF�z�� �`�m�F�uy/�t��-��G�G�@���b5�d���[[���q����lſ�y/H(��/��� ��/Sǝ��b�p(�췭�{i.�f�<ב⃓^��4	�����\�"mb��$�A #����^�"��5R��c����X��!N�sE��M�t�В���5!���V�ȍVd�Z:�tfoj�j�a~�9�\A�.g3��0��4A<� s�gKaZ�N=��êq	CM@z� m��0���7����c�R!�"�pfՑ�K�d���VB)�C�l��2��(�0f]��;\��#�Y6�y���3C,b���r��*X�aDv�P3�"�Dnq!�p�{Z�x�I��(�g���*f�z�N�a�񐝧="�DOP�<�������=���h�A��Kk�-��א-S��Qe��g�.i=�	��=�2u����־�c�Jd�Uf9�M��½7>[D�W���v0kI�Y�ɭ�ـ��u��Tq�,�s��=*���@ޔ�{�]y ����֘��˚���tq�X��+k8(�|Gd6�$T����[�n�b�z7U8{����F�k�W"��W3���#���.@vI����Pu�}P7q=�;�611Ӌ2�h����l���f���������:]�G���x�+ި���X9t�R,��J'f����ZF�,��4�H�u��(�{[,mɶ��Hq*
���Nl}��Ora(uD-�C�!*�Ϳms{��������������kZ.�,\i����=}7b�l�Mz.���Ӵ�C�%`9�ou��.���t�z�$9W,�ZBn@i���mm�������*-�Eٶ_f�m���K�ӻ�NSr�,�ؐ�W����A����5e�E�S�]IGlN�!�K��Lu5s&3U�	�E��Y��:��ז��gp�.���o�z�*ryF��}f4R������ׂj�:��G-�}0�o������|tp�#��!�ZΜ+�������eu�)���l�b�'�b}u���AAn �Ё��坭���(Y��95ש\]i��姰H,�5�ǼW�s��Z��6�x��g��+���ܘ�n�u`��Ԇ�vJ�>��q$7���.�}&%Zd�
�Y��+U�M��UY�y�ĹS�%�4[ɻ/U��o�L7�aqm�Y�1�y������̥G�������q.o�=�z���2��&�F|a?�7��]X��	Rv�נ�#�9����gۏ���>i߈�e����B��{0�3<���&p1�WHAϴ36X�o 1��>�ܘ����{y���}��?�KFh�@%H!�[p����� lOdY�����U��.��W��4��hO�Ҙ��,��BA~�.���ޱ��GLi<H�U�~�MJ����}���X[[�fqR��ؾ��&wZ���S����u�A����ے�CXH�qď[��׃SB�<��'�N�l����%���f��i]mpu�oY���M]�Kl�k�8��}7��v��"���KK�٧�����j!{���d�>z%9��ӛ2ʬ(���ǹ�)���Z�f=�&�y)),��}�`��ӈe�e��@/�)L�`�U���'6�+%�*�1�ԓq��.�P ֋�qj�eG4�\���y81�����8�P��uvP�hu�B�1^���Y�hpNVٔ���R��=pngCf�D�1�K�]S2����3��񥒞9B�E����}(�5,�29�X�v��52�Xŝ)��}{]u��D��^�����(�{%���{�|b�!u�v�����ֽ/�O�^5�^{V��O��k8.}z�ik��P��e�|�*B�a3�o��c�3/�cP�P�x�~�<3�g���ǥ�`T�խ������]mg-�N�lI�d��m���0���Ф����b����U.M��ޑ),H��u��@A�)N�G����_d��!�un�x��6,(9+�y�ζ��F27�q�F8��D��	p2"�Rd9!E ĉ�a&/�|XA�a�0�m&~VXUM*�����TP�6l5rB	�$3����RTSfX9����Pf`��6�(�dDUH�4S���g{{{zzzzx���fu��bZ�X4S�N[�dDP�U5M)SFHFek3��>=�===>>���g^9�UQ��6IH��DP�Y�C����b4�G#"�����OooOOO�����ל�1$U��˼�Y��
��&�,*I������	���̂*�!��
�e��CQdX��AE19��̩�#��J
��������&�bi��d�Y�Ѷf�uUUՔ�ASE���-R�!�i;����T�;8UE5E�����[��j2RTMn)�'y�VM%4{,���L��7Y��$(�6C2�"s0�0jb� �g��j�
B����& ������s"�v ˸͌B��J�r9�f��Iì
�E9~�����Y� ĂPK�y���D
zJ3#1wVE5N�UJ����8��:����%�Nb;�����G|&'�	�����Z�~���I��䀓A� ����Ř!�X�\�
��ܷ������l��<du�#��R�%X���˳��R�Ċz+���4��<Vu
,9�>�2�0�an�
��V;�
�uyT��N{z��:��r����mS8�5�kݣ(tCu5����1�]�5ڬw�sI!�_�u��,�O�����b3<���v��->{.� k-e^&;B���-��x��k��}��Ռ�oxְ3���}��m�|E³TiZ�Ú����u&�g�"(�o�lO���u�4��N��y�>|��Os{ʻ����A޻q�8z��.�h"�!*2�YN�y�8MBqG��F���H�x��ۅ��1D2,�9E�BT֍흥"��;}�c��*���e>1@x�R���w��׷;q��:b*��(��7R:�c����m�1��s��y�d��Y�aN��1�j~R�%���)`a
�V��K�/z;�\][����,A�Zr�ھ���GRP�%*���mr�|]ǧIѬh�Mp�EZ���۠������o|�.9��R�����w��k�W<<�\����F3�#T�p5��nR�����U�\O��S˴鹚�{|�UL�\�w,��#���2�`bg�=V����g%�����%�/ƹ[S���'2�:X����:�S�m��+�ʾ�m;�C�m͢({ *�=�j��t���+I�Vj捫�fmGu��R��Uː�}'ZV���2�q-� ��9A�F�Bxf�c���To+:���x{4��fcFC�6�͝����E������i廲����#}��7u���/��E��i����E&"����UϏ��q�IL��zG]%^Ix��9���vo���S�p���sZ݁���t��v���N_k$ٲ�"���Z�z��C�:���Ɛ2�����7z���ײT>����������{c����#	Yk�V�8���B��/VH�n��j�a�I-ky�T�f���>ܖ�]�].���N����E�v=�`�O���w3_�>7�����4�GGXR�����A:��H����g�Дay݌��T��M�+�Y�M�\nY���p��)K�M�ڨ%�S�
�v��}�U;bfw>�C��á�5�s4��1L���doi�3D���0� l�t��=�5��`Z�.3����fE��(�9���h�tg��t��f�ʁ���M7H�й��d��qxާ����W������?���AT)�F+���dYȫ:d�D�9�ۋ��E�{I⺨[\z}�Zh��G�j�|�3UX�",��s�͈�q)L��@���vQ;n`c g�mG����@?EL������q��kea��i��dp��;�7XmU_�h�:[�`�w�����D�1��ۼ����٧��g2��1Չ���V�$���sM�.��q�z�L[�1�5L�5s���n葞C��kϵ�{v��M�W��[�˼X}{x�wb*��7�4�P�k�f�\��\�1���f�Vʳ���R�q���Oo��q��T�jq	n��m8�ZrS�G�0��(�`��r������N�2�ʙ�ԻY�;������ܓPyҷ�������AU��� �lP���/��[��&�	��3u�LS�.5;.�.���Y�s�s��6�e
{���aCS��|�_���E��M�(G7Cl�2����?6���+t���k�������;;�;s���_����w���H[;=�+���L���~���?�ǪQ�/���{����K�
���	n���_qQY�����cn{������w��s��Al+	Vx�\�R:r=�m���`��W2OT���{F�uT죌tk�� _0ά����VB�3�o@1!�m;��n�X����Q������^qo�C���r��1b�d��^�^�<v�Bf[�de���I�X�g�xh��^�*�{��US�l�{MU�X�U5MTG��5mBM�ml�7w&{��y�GoZj'��
�f.��;-��;h1�M��i���Ǝ$�<��m{�o����n�`�1����g�Km�1��ky�O3.�����ϻ����l�V�N/�p��[�~���g��fs��"1�U݆�n�v�A�����-�>h��)��K�cCv�vvPR��.�%{�>zs�~a_̲C�J���mtX7BPZ	]i��ˋ&N�e�'0�醞���GN	1��ʬ�+Ύ�O��#��v�/�MFޮ���{���|&&QiЂ'N���̔U��k�և#	K<�+�W��ު���}T/P"����=�j=U
韼ױID�-��wMxV����>Yw!'��|����t��
���T<�Ec&B�T6���a(��U_���U�g��a���)uGO�����m�#3�Ϙզ�*�m{Ml��q>Ͱ'�yM�ۈ*�Z�l�+�zݥ�}�Vc�,���Uwf�qX+�AJ۫΋��Û״���=�b}��rq�)�eSD�I��Z�G���$�W*�}�M�|U���p,,���k��d��5��4FΤ�'���<,��N��6��A��l6k&�i%s�
���!�A��:Y{�����L��q��-0	��/S*瑣�^zm�7;�.Kg�z�]Lx,w��d���[Ns��m.�J�e�Z{6�i��А͠�{��aoN�����`,Wk=d�`��(y�	�Iy���b��W�c׍�e%��_k�@�j�E�i�-.��̞��\�D�K���h|�U  �f��d���n���t �J�F�mv�SiJ��j ��ǽS\|�w��v��� ����
��ỡ+�}Ut�`c��/��w�r���L0�m��
�x��N6v�B�C�r�v����
thǇQ>�w��+`2��x�f�ј�mn뙽�Ng,n��/ڽx�.��J�f�T�Q`:�s0�/h�j7,��Ă�4���|ԪG�Ҙ����L2/3��H\q������%�^��-�p��.�̖r*[m�a��;֯2oݙ�	*��mz�������O띄�	�$'�ꞧ�*��Q�`v&~�ay��T��TM�$�a�uW�w9�td)��};:o�敀e%m�U��b�w׌T{��Lj�̰Yv��.�f���z�G�� b��%�Vj捭�sAݩk|*�Y�\CG"հ����L�$=d����6�=^!�*ԳB����O^������]k����h�h�ѐ�,��j�13»9v���⑿tn�F��ݹ����ƞ��O�ظm�5X�򸐜�I�Q���ݵ� 㗌��)|�>׾�~|�aC����o�T�`��Y0��7���u�ҝm�Ső%.�ʸ��V�� ��Ħ8gw^����[�2|Z�$�0#y�2XU�2��K���U���g�b�40�}�Jf﷨\�)n�m~��6�n�k��dt_7_��S�������a�of>ޘ��;�9�^����i";:�V���Tޝ�m�q��V�=�9c3\0w���C�FDv#Y(I�X��u�F�DvNp 6t�����9��^�\��X!K����8�5B��c�l�*s&����y& ��F��W(n������޼�E� <��2d�n���;�I���Eո;t(�#�6��Q��"i��]���bn�:��sdqh��j-x�i��X�&[=Yݔ5�KXa��s������ۑ�y���gS�Ȣ9,�0$r����L�F�}�p�R�5Q3�������([P�����	���t�z��9�"-��z�'7'{M�wf��KB�*ʘ�T�ͻ���^�e� ՜;���J��~[�F&3�����pXބ��_�����O��򴜂Po+(�L�8���5�u��LW����{����՟����}��vfs�;Ù��y2�X�-��X��̇��r唹��4F��z�V4��+������C�>�)c�r[�hL����x�����	��Z�L�e�.2���\)�b��xF�ѯۯ�K7֓�F/l���������z��6q�	�щ�}�4�#D�pQ4z�w��Ӂ�c�C����<���V��w����LMw3��n���8� �[�ژP���[J{��%� <r#!��i�m�V]J��H���r���e�ף�{�#�C����o�N�st�ܹW�u�,��|�z����;T� �TA�M_B�����G��2^K�-�%�_^��Z�7�Ey̱�hr'�eӵu��f# �S���<�76\5�N�8��>�#�����Y�8ӥ�Z�O�lz��[�\S�.��8�L̸����΍����*F&�^q��f�y}�'���׭N`N2���C���H�8�Ғ~̤��F�\is�^o&�g���L���;A���� �]N�&\�#, �Õ�ug
���M>�$1�,�J):���Bt��:F�#2,�b��ܫYr SRPE|�XK	���Z�����'�Sh�|p�p� PEX�0%K��:I���~�
�hVTj�[�J�;��ۚ�l�ÓGu3uj��������r'�)E��.��o���o����;��T����v�i���i��7n��9���ν��Z�� ��h��&=��םP�	��<�YT���^��	�\Y�}=��%TWH����P�A��T�f��5zzާ��5�n
ݍ��Y��X�2��J*����Q�t	��Vgzݕ��u]X��Րμ�At5� �W>���Ն7#����R�ϩ������#���3�Ԗ�l��S!��M�%\7����&��.G��ݧ��	�si!ˬs�Ut	U����@�+A���}@p��9Q��O�c���SYW.�{_ֲ��Ϩ8��3��g����ue�i��B�n�����36M��K�����\
�RΏs�M�X�έ�f�>)�,f�p��L)�/ț�N�s��P�.��2��I�ٹo���w�,��x�mQt����~��:W޺wU���o4�v�Yj�{6���pcO�x>0���������V�̲��M]_D��m��ĝ,��`�찼<8���mf%�oԥ�O�;M	��J ����%�֜�h����x�1&��.Bj�j�> ;{׽�x�Lt�{b0�����]Fa�n���Q�gZ˦��S�޼oD�V7ڙ���s�/̰��6r�Z���h���I�ٮH=mK�9�8��^p;���#�#Q� �g�G�n�|�[b�Bv��ǈ~[�o�!nS�q��� �[4���.�^���<��U�Gjd�h �]����C_��k	J!��oN�b�񑚦v/��X��#�S����U�U�]���<���d���	�J#�[�fBy��sPw���狊vU^�d��ʑUq3��Fs1�ĆO��%�h���M��7I�G�wIV�r|�2��V'L
��J��=��]�&�B[T�D�e�$��o��7ұ�K�flA�/������#��ۋ&^��P�nT�1J��:�1z�>e;�7���̎H��~����{o��)�i8�Vvo�:�D���ֹ����x�X�����}G��A{nkN��}zO;�p凮�3�Y�qN����y���
�[ë�������m9��k���]�^��ٙқ�t)��^�oc\����&�$(�zTe!}gۓ`�"���o���{"�Q\��)y}HP���YsR쎟^o�^5׶��k6���P	�,;��7}I�Uю������[�B�.I7t<Knt=˘V-ۜ���Wʎ�M^�ո�MP�����D��O	 Jr�o��r�$�V�$c���Mp��X�����P��Y�b|^�cToB:��4&eb�.�8����L��V�8�p�*��:���rMT�o	��VaÚ��X�
N+�=���ݽ)��)rŤKn>���z1}��}��%�9T�>Ĳ4#��&�o�r+���&n��`�b9����h-i�6�i�B;C��i�܀T�>����!�	�·1���N��X���K$�ʺu0I3!�ڎ�o�s9$`�ބ'c|!���8�{9򗊺s���#b��U���dl���4�x냢�Q0W9�G��ʳy�KGr�b���9Tz�6��Wb;6��N&
�}�]�:�ʳ��)2�JG�إ�҈�����8v�%Y�\�+n�V��:�f�G����`�a�ȃ���,:ϠS2?q���ؖ�=	�Ϯ�^���	�\�z�	;��5tp`�������>J�Z�o�����jU�|ҺR�K��~���W��:��r�w1��d6V���P�&'�s#;�i+'R�[�qg�>��2v7�(�p�tt�*e*�K����F�������8R�`�W`����;Cı�<&����xl����,�f����o�ٺ��
t����38F��vڢkM�^d��O��.��aT
��]X�l�vZ#<��T��
�DQ���=��U�cp�]�9:�_;*�_EW�4�u�+�L��ܖi�'��*��h�L�\�_nR��=�v��]D�U�K�#P1�����A��0�6�<7�� �<�#�3lu�ڏnn��E�[����ɔ��C2�lU���!��7����.x����F8�n��(7�O;]mmؗ�8���	yZf��8���4A xҾ$C;̺� Tn�f��t����z�#��rYb���vÚ�@�^���J��D�O�2ʤ����Y�,�Ǣg^��0�������P�r�-�ୋHF�K��T��J�5-:Y&�u�#�e��e�E�w#8��}�}�!Kx�Z�[ۚ�&�J�+V����)F�~����s=p���o�:3�i���3���V��g/>A�:fE.l�mN�;�n`Cl��K�:S/�ŏ#��u�`����AL��ċ>r �^XQ�=JS�Nԅ&�f�Α��E1>������ޞ�������OGd��ԄTͲQ�MTܲ����*i62��%����|gz{{{{zzz|}�����׃�9|Ƅʂ���r�,)��%4m�SKHD���8�����������?|x���Y�e�LM1��^A�fad&zq�kc"���nY�9�%�+!*���
*��eԙ�!��NI�L��wP���d�9!f��ITP��#��RED���l����
��(h���JiJ*������2�	*�
���ʐ�**(+`2�!��\��� +
L�$�$��r��3�*
(m�2Z��)hh��l��ؠ�)�
0�$1��}��:�;��0^�WKk%��A�\8xE|SF��]�0bGV�{{���D񧧩�Y]�EI�ږr���e�ﾪ��7MW�rp�h_u��S�봵���He:�[ە�1�E�ð2��7��s#�R�\9Ҵ��j�Q���Y�25�tr�3ҥ��w7��[��PofD�Bp!�G6H���p1��h����+���ih��D���+�Z*��c��_���U���-�1=�ߺ����^z㶲0����A��!�<<x�ϙb�u�!q��J4��@�-;!������}��F�ɇ���8���)@Gf�^%�������d����˹�ƺqcx�m7�H��Y;��|����0l�Q�EÞ6�|�gH�9�m�\��ø�n�WB�k�3�M7w��� �b���,��Q�&r�c�hC7�r&uHŸ�s4����%�?Hᅻ�Zhb�;��;�F�(Bl���
G,�i���5�7d7�_-��e� �GKϞސ��^ן��^���)��d\1*�N������^���S�-��z��ڟA.���[0��nk+p���t�5�;�S93	:�S��B���݃� /�v=�Xsm]����U_�6[�v̹��~��z&NT�&�`̬���'#�u�;-u��ٽ��P�&Zt��|#Sjg�f�O�~��3DȫwCX��q��^�X���; �2�&�_kF�����������{�X���Nc�!
��֑"2w�3棭ΐWp��1ޱ�L�>@��������1v(��֩��j�y�54T��[��njEb=Vem������v}���]L�n�aXrjF��NbR򽇼�P�������ポ��q�9����Ƌ�{S�6��t�fER󴦷�Y!�ٲ+�P�G=��/��nvf��ۋ'�oT��d=)=׹�Mk�,���qY1�d�N+�@�GK�=<"�ތ-n�}�>o ʻ�J<�G�[�&h|�I]N��=M��c�ꦤ��,vp���xꠑ(�u�!m�Ӿa/h7�c{4$�^)�t�2D_�ת�`N���<��^���C�]�Vںm�� ���o�o:w�*7F��(�2�x�A�LJ�Pa��Gûsa�/_o�/`�=��S}3��R���1#�G�2	3��q
9���@���#�_y��!+$˘Myn>�`�d�������K>���N&�p����{�2�]���7H$��;��>n�=28��Q�R;�,$q	���*	������͛�"���������}�q���{�1ݑ�m�_
4�ƪ�)1ԧ|�]z���Z7���ՋD�(�D��������/����#!�O0O�!Ǝ2O���6/�֣��9����y�neY4��Q���;��.�[��W��Zr,������t̽�˿��pt����68�k�+�'�3����Yr·�\�>7��h^���-�W�jk�#��3�W��ϕ���L�y�OOL���Vd�YR*���!GqG��rr��n�V�ر��rԐ�{X�c�x��̇R���P*�B^ tI����+�0��fW1�ns���tS@�`b�E����U�R�㠾��J[����)�@��m�U�{��wyx��T����}��Ьæl��I{��fs}7�B�X�y{�h>��«�T��A��d���K���"���ܺT�3��"*��q��d�R�!�i'�/8��f��s[`q=�5n�<'�a4��ڕ�k+����8��E��y�೺�(�/��F�P�7�9�R��D�V�+��P.�j�>�>C���u���{(a毣���'�u|u���Hm[�9�b�� �}P����k�Ȯ+%�;���:�QaZ�D_�56T�R39+�'og~�⭽�YWZre��
n��^<�*3'�0�t9����vӁbV���.�l�=�u-��nm�'�M3���[Ey�צzJ#O����>Ӝ�.XGdD��1�q54Fm[[n��Q����|�4}>��W�Pd��Y�\���.i`�;	��ǽ�9�7m�cl�c�fFx����x��p��^Z����s��׻�ޚ�w>'�}�j����L�w��c|���N'X2h+)�;m�ʽ���}�{��'O��b_���6K��Szj�}�lu5{��Ɛf�����Mrl�Y(<��=Ț4#Ӂ!���O)�<�5PV�_߼]|��+�]ѭ���R�ض��
������T�����C�,��£�^�bU����66��%�朎e�jn �y8�Ӡ�J�*��9���z�xM��]�B���n*��.A�wfa��(�f�V*e��|ו�4s�eN*{&��QU:�ދ�nG$1�{X���d[���T�*�{�?ӽ�;�W� �U^z��5�>�eC\�~���V;ch��Լ9I�Igz�<V�3i�g�Zȋ�cP�+�C4�]KE&�S{��軆��j��Nՙ;eNh+2�,^y���>���W�w*0��L�n�Ɠ���z���t��KJ�ע�h���<�ڑK�6`H����ȜvI���ڐ�n��id��� ����WV/3r7f�n��!�� �i��|�;o҆��U��+P��n+�����E�a��1��0�ʊ�ӽ�@��yr���{)���l�	U���iEhg3mf��'6,�*�̼���n��EyH^=6�7���ߏ���T\�׀��?h��������y�n��1�=ߏ�^���<�p����_��[sSk0�}z�x�|f�:��e`��s�)�.��H�M��m�Af��>��]O=�P-T���ږܾ�(TV���W�Sӝ]33rO?�α7�Z(����p�b}��� ��������f��l�l�7*ҥ�@�*�wi�<٠��&��w���;����ƒ(!�g���qJH$&%�
��� cf;�p\�q�� �g�h�����s��͜&�6�@ya%�<A�0
������)qQ{�s+ٲ3aC)�Aƨ�k�	`F�����O��_\5��
́`wW�HD�E^A��I�bU2_���*�Dv��B�9�M�@x�f�{JDMuP�=.%@�M�wJ�x=[�/J����4�:��*��0X�z��;0;�]tF�(���&U��(��8���]I69��~��禔e���̝L�i3S��O����)���
9WҕW�UM��ʅKSWK�L%�l���6��JG��"L�C��#_���ee�R�*�%�U4�"�����z�a��u�t�7OY�;2���5\Q�Y9GF�4����r��![HP����w� �'s]�����v��nW�=�ߪ�e[f7��76~���I���8�Vݱ����Tp�=%H��2,�Q�9�B�=�A� �6��m$�-'
��>�m{=��s��|�1�\��Lg��i;!�l��W�GF�ba��ٶLȻ8��$��Y���h��w��:.@6r��j����"9-��zՊ%����{4m_wll�Z��囋o���;���u�u���'�Z"�n��خ��^�Y�4��=�Wt�ܕ��{�l�^n���	kΧ���B+)L����#��K����R��\L�e ���-#18[r�4`�����=�Bc)'}݈P�}Ԋ�:ՔD�숈�7����//���0B-!�Ԥ@��&�E�3�n�^�6�rn������瓓ћA���ϲ6�I�lȀ�͋赝�;_�Ꮺ?j��~fN8lP7ov���6��� ��G;b�9����)�kf��z:X��{q�RJ<��o2��_��@�t\�R����A�lw��=���=ZQ�j\�H��F�,����b��u�֪#��$C:�T�b�٤7�_1ь����M�Sp ��x2Ȓ@�yq�ּ����ף�q�Xx�s����(I���y�6kR�
z�P�`�ڇb��nwGY5�P�_�l}|�$���)?�|��;�[���Ӵ��U5bJsܐ�"�b�w�{��fJ�曎{W.�NW^�"ֽ��GS����9\Y��o�u��/�ԯ{����!η܉�fSQo���5�_G����pA�0����Z{�ۉv'��v�R��f]�wY�CU@n�m5h+�f����eD�/qzsU�f��� �;B�܂n�rN7b�Z�@f�y-�gy���\�2�w�&����ǥ�8�J�{�+/��d��\��7X��S����1��+�vA#$0o0z%��4���;�'b��
��R�|�[~�|�l�0.EF���c�-*P/F`���BV��k�D�U�QˬʎJ��l7NO#�7�3%�~��eό/?;���LlR���ޛ⟨%�j7n&M�fṽ��-k/�[�����K
'�&Vzm�����ߙ;rY����Ɵ�rkc�b�xsH������~n��,�C{�4p\��.��̮®S�jujSZ��=��O+y�w�Z���VjC::��x�Y�&. �f{���w�t��J�@��3S̑C��W/�C��7;��}�'�N�hV�ٯ���U4�w7q�����Jz��M5���vPm��/��h	�r��v�*sfۂ��uc^���Bo��=�;�7w��XG��#^;�Ǣٟv��[~���V�P�@l��;28��1=-���a��(>��4�3���Sf��<��^'��0b��׼�~;�zƃ��\��P����,�>�w܊�ځ�$��">W��3Њ�?���wl������X�ӌ���*y.!���h�VQ�81��9���"۶�MVg��v��YDiY�]=Ӝ�g��#Ѓ��v��)�aLb�ɏ=�/>���k'�&��5����Y9��U�YBJy�\��{��]!�X5^n��2��2x�ם�1���{�n�-�FI�*��̪� �4����$1ҳFq7����rw[l�	�����	++�6MĚYK�g�|h��qrߡ�Ջ�5l�t��ɱVĒ��7K-N��|�h��J�22�[�1�H�(������dz�b��=�U��m��I$��I%�I��, �
���C�婊NV)+ǺIj�Wm4�:E�D���h�G��W��[������[2�M�/9����/{��]�������:�ǐ�
ے;{
��>O�:�˄B�Ե��T?g>;�qA�O<���ූ���GL��SKaqֺ��φiiU�L"��]��������8�����ؐ(ԧ�T����)��ǩ)}dL2�|��ʼH����;'�q�=o�Ƭ�l�@�T���))ۭR�3���h�����
��e�.��� �V^��=�a�~�P�0؍��������K��7;���ݙ\<���S�������k^O_^XK���9y��QA��H�Sl���g��Os9@��͈�mƸ؅��;�ً��7 ��Q��U
�]����bm٨}-ʪS�:����e�yyh&qP~�}���S���'p��+�M��`����{�:����p�]�(�5��-�֚�	��$b�������������ix@W?�AQ�'������9 @Q�㡦��L��>��{!� R�HBQ!T�!��H��FU&�Pd$RBU!��Hea	T�!EN�D�! [��!����!��P�E �tCU@7}Bt*J ��Ԡ�B � �B��
H#��&J�"��`!*�B(!�B�!�B�!*�B(!(�@�*J ��B �
J �"@���H!�B�!(�B�!�B�!(�B�!(�B�B �(��B	@$!��B	H$!(�! ���B�@$! ���J����HJ�! �! ��B	@$!���B�@$! ���B�2	@��B�H$!��B�B�!"�Ӽ��������(��� ����|��o��׿��A��s���������W�������W�����/��e�w��?{���{����O��� ��g�T@b�O��D�������~և�� 
�����_��� 3��������?�O�������aY�8�*ʅ(� �*LL�DL�A ��$��*I ���$�K �@��"@J$!(�))(��JJ��"�$H�$)*�H�)�$�J0	H�(J�2,� ��,� �@���
@���,! �(�(�@�,,@��0H���L(�#H4�R#J  ��$AQ�J JY�J(�e U��
0��X?����؟��(�*%"-""%���~���~����������� U�������~=��zO��?�����$��oڢ �����	�|w�Op* ���_�C�a��~ T\��w�@��� 1���`�Hv:������t�|z�:T@o������� 
��{J�����?��~A׷�~�� }���C����W������������AI����0���=�������.��<O�O��DW�����& ~�����{_���@Q1��� /���y������������)��Lŀ-,�0(���1}��^�QP	{j�T��a�%H*���hШ��4%UI)U���4�$���	
��@������$DRUAT��v�]أZ��Zj�ά���n�wn���]����ku�wn���v][v��7N��*���]��qۧmw]��������<�]l�z���y:��vti͕�����۵�uՕ��^���sk��qK,m�mWuq����k.]��g:����m˭�꭫���Ӷ-h��e�wWZ�6;�����f��v�v��8�U��u]ۮ1ջ��fiv���hݍn�l�Wv�gS� 7��}:��F�]���=�]��y�w;��{��w�3\�I��8�����]�7��[S��]{zhq��^�{û�7Ym����sy�u���k׽7��4����owm�k�]ͺ:�N鹶���� 9���(P�B�
7}���P�B�
({��o�B�
(P����ן>�Qv}.��w����GyOsB�{VY;��MdM����v��5�(@���*�W����S�]���.J5�ݶ�� �}�ֲ�i�漺�p�:��.R�^��v��;��Zt�n��竻���v����+{���䵚�r�lӻX��k͝���r�e��Jgm7;��m����mm�k��m�J;��v���o�  }��(+}�5�ɶ�يj˭��h���s{s�mk5�e��V���2'�m����::�{��� �I��mm�=��Ԣ��ޫo:v�)���v��D�U��-π  w��J�i^�ۂ��Q=��*�������j5@������V�y��UzY{��=��^޽�P��{7�AMW����Uҋm�{�����n廻�Q���lk�P�>  ����3/w�x�U�Mo����V�wV���G����f��5z;���´���ov�mT�׹�UV��=:��%Y��z��-�:jU2\mrA�]���� �רЦ:�u�� Ʋ� 7}����T�0  ��)�	���P��� �u`  -/p� P1�Jl7���&њ�ݛ-c�  w��4 ��@ ����(m��  q���  ^��� ({  �����@�,�o P Mz�  9���u9Y{��������7|  n�@���۞ (��m�  7���  ��׽4  �� Dn�@ (s�� yu��w{�  {]�2��L�ݹ9mn�n��N� �w�  f�p  ���t {�x  v�X �
oz7  �� ��������� P=���  > �~@e)R�	� "�ф��(0� )�
z����"��	J�h 4 j��2�D�  z�B�� 4�O��ǳ�~���$�������kkgyr��b��9B�'Vʣz��~� >��}�x���ګk�Z�ݫm����uZֶ��ֵ��Z�k[eV�m����?Ͽ�����[qk��93�QS#X��#�˫6)�Е�@��Vsv&�5�h�V�hl2X�Źdw4m�a��Pe��S���I:YiQ�6��P^ִi���D�ұ�v��7���r}�B��amʣ�LJ��Ŵ��@bgn��ir������.���\UX08��D���Z&�弤㩍J��i�MGr����0�lJ�vZߙʹ4Z��e���ء�G�bfѹWi������el�m�a�0�훺�%�����tHRQ�τ�Cok(fU�kV�1 �52L+�s?�pl2Ys*
qQ7nh��5�R¢5�P�[�[|������Zgi]�{-��e=�R�`�w�-]�q�w� ��1{3`ڰ��m�VlFl0���XQ���ON�Pa�"X���j䧸��( �A"���t�X&����c5S��*u	@��n='35]Y՘Ť]:g�d;��#n�)W��j�ˇQ "����C.���mGhڬ�u0��<�ʙ���h��V�
,�!A�ʖ�.�kB��3Vn,KCɴe�j����~U����df쭘�A�[mhv�7E�1��q�����d�N�Mei�a�F��6�i��Y*KX�O�I�-R������x6K%�V5�5�4��a��i����v����Vkr;�������$��S�òʬ+R�%��ok�69`�´��h�ʰX�[E|���Gd��׌왮�Ґ�=�ᚉ�p�^�t�Q�"��S�
�tڣP�ܭ+f��)��$��^(Y���M2~��)xL\ai�2b��Zt�I)!���9(�-��i�ݎm9�Y�x-�]X�Z~�[�l$�Q�l�
/ƛ
i��t�O���B2��hOr�p��;mh:.`�(�4�6�.]��K��d8�[�4���-M�s5�fXhm�]Q�A�14^e���L5tS�q]��X�hY�H��)��ZoVVP( &���r�b�@Uk���z�n�,%���U4\�J��dYf�v�ɋvu�K	j܋["��t�A+��;�K[�P�Njy���0m�8)8��2�i��In�Z�Xk�0M�7�AH�r��8���F$&L[oCn���- ���D�Á�׵�fȶ�em�!eǉD�[��O>Rz��hP̊<�a^������j���z$&[4�U���f`��������%c�d�-��ٳ1�
�S��e�0�E�I]9oU�a"�*�1����&7.b��F]ȮҐ�e��<�I/��������mA�%�Ei;PTJ}��r�:%u"QQ�lcH�p��x,,��EKX�Jԟe�"
#/yE�u�m�Y:idsě��&��@�ln��=�� ��
�M��7v|1nݔBt����J6��8���T&�nfD��;[m����MAX��<ʉXvƛEغ�x�d�֭�E�y��4)�JX��"\���������0���Ó �Z���wW���I�����;G	Ob�P3nɛ"!�B��k�]��E2��%�D�u����j��K^�M�v6� ��e,��Cb�M�i^�Æ�Xv�:�[����P
���u�$��.�P&�\{`YV�6-��ݡ���V̼�J�#B�bB*�`0��=*��J�R��6�I7�&��d���<�b͹a��ުѻ�Vi�:��@i�DwZ(];�Z8�-�M�E*ͤ��=�;V�a�J�&V����i8$�{N +t4P�b�,ث�Q��fJ�**�6�l7r����,��FE��HZ�5���X��n�(5{���XNĬ�z���)����72�O7n;��{2����91e�g�F�M̙Q�.Lq��Q�Th��+�>�J�FA7U����B�HVKt�Cvݺ*�h���b��e�7R��Ku T�]��SP�B��,^e�Y@-�V @�-n�e���H��!���܋�5��o���l�C�����,<�6�)�qR�Q�A���W�-wB:/M�$ �ع.o��Q�m�A�[�:��69�

�X��SV1��f�+"��7a�ڴ4SwY� M��W5<Y31"#��
�B�fV�'�h;�f�!�3^5�1ܠ�r!����������S�@#�"����\.̔)��=�oN�:y𷻑�3p�ߎ'i�wZqc��sa��+	�m���h��z��ݼL��S�&�Px�K!v�c&�Ćbif�1���S��?��&2���b�}�� �Ph�ɿkc�����.��'n��)�U���Ңh����J:���+s�`��*d[�?���m-7�L�a_�m-Ph�+u�+
�P�C��t5BHB�D�-]��m���F�]`�70* x�8�<:�Vp�4�HR��$h�n�ͧ��-�ܺr��	�b���/U�����XB�5��(��N�e��hY�J�f�F����J���KrZ��z%��S{t͛��g%�ЪР�ϮF��%�Ӊ���KF�ZҺ4�0�^j����ބM��m���]/����,D��gY	�JB)d���f�>u�pm�n!��-Mn�qQ;b�KA�:�zb��A���� P�E9 ��I���� ���{%K�w�07n�T��;�,Lq�[e�YDe$Iٶc͛��Yn�Q�H�-e
�vđB�-Ӻd�i���l��؎��u�[>���fˋ37t
�4�F�0��A1vMw�{O��.����]��/S&^%݆ͻ$7$)H3d��^�I�U��nm:A�dT"y��ӻT+jD��E��J:J�]��PֈV�#hђ�[��h�L�Wy��ˊ��kJ�V���{I	���2e��a�mmէI�jc �,[�˄��Ȟ{� !�D���x�M\**h�ݫ�\w�)�7�-l:Ou!0�{r��L���r�6�f�1�IV�ܨ��t�A�l�R5&�vn+�r���ub�nK�
��r*90i� ��i̎���4{��P��WM'Em\2���l��
��V�>V�۩�����p�8&Q��0S��݀L�4�kOh�qn�R���Kz����[�f���U�3X��,�O�e���ۢ��ջwxVkV`��&c�ӷ�^Y��fP8X��ѳX��\���*L���Ɂ9ee��t-�5�ܵ���1E�06ź,�X��qU�;�ZB��Pff���k)�B ��wB�^Ʌ�H?���Tcx��Y���+��
�V��=��#��әe�����Yd��y�6;�j���@���ѴuT5���%`���*�nf���4���Z�b�Wz��V!K1e�J�ll��^���d8��6S��ri�Y�e�jKD�i�voe�%��C�_H�T.'�T�2քԤ���;�X��+,��p�9�?�7*�#.����;V�ѐFAaie�45�̢(��֙�S�ER�j��yi3����!���ˬ�A%VB��u0�ǅɮcZ�R0ܹ�l\�w�`7E��i���{6'�m<�����T!<�X�����������Ye�x�!��B
����י�&5\�CpbƎa�I@�����XRy��Հ�d`��z�S��c�W�Kn�����dLƂ!��^�'���c�m����h����y����}�!�s�������r�T��b;�G	�wV�%Y!`z"F�i�4��DZ�r;�s+6�.�1�F��a��%��弲nn�`qne�
up#a��c�E�R�@�h=|���F+B��-ٔ�*F��{eXmh��v�!K3J�YG6�����9}m��訫�،�j�|�Ie�2�l�J�[��Vk�d�:�Z�L7b�w�ˣWN�z��h��F�d9P��[ ��tz�[��OBW��Au�me[����թ�H��*����-bc�Кzp\��F��*�J]i�z.Q�Qؽ�TgtP�l�u�3M�YnƽE��O)�t�ت3�j�鉺��_�أ�ùz�+P;x�݄a�m�b�Ā`+�$�j�u���՝8��X��ۘRO�Ӹ������Qn�z�����B�M�ʙ,;�THU�AS�{���B�!U�&*��v�E���a�C+#����q��rސ(���s�7R�n^�3.��"��d[�4d�h+��6ݠ ���B�1R�I�l1g4��Z��,�N�*�'�l���(�c��E�� 1�D����
�2�hDuV�V1X抂c �Pu��J4U��n�Ą�k&Sp0ku{L]N�L��KQJ0�(.GW���&����߬V��N	{k۸(��r@S��b�)��*�Q�l�2��E1�X�*�1v����B��f��S�*nǌ]0\��Q�wy�5�3f���Z*�&��v�ֆ��J�RX�[�c`l��U���j�8��w�Q����v��Ɔ�vL��kX�ق��tU�Oh���e+��^�aU5ѫw��[Y����Ԣha����p���ᡞ{��,MsР#�`o�|.�a����K�̥�d?52��Z��ItU\�G)�!�uVi;u=�ra�$ÔwZ���o�4ÈU�kb��m`��Ĭ.��9��	�.csD4�n�Z����b��DRb��2�&��X�*�ɧ�����i��.!Qb��b[�OhTtH�zFAH��)2�cv�5�v��-�����y	�J�UH%(kO^�W�H�Lݛa-)d�*�,��F���)9{�u,�kL�Բ!ph�b�%�K6mMX)� ��B-�&ր�X��_;�7�l�br�әs!MSAVҼˋa�	�	���P��[�oLU3{��D�j������mwCr�����j��;��k�JeLJ���HY�)�N�-4�v�#.�(^ޕHi�A|�t�ԅ�w�2��tu��#E4�Z�_;�N���tØ��7��F���8��5]`��H�Ո45b;�V��*lVƼkHʶ�ݬ���lA�^�Q�Vѭ���V�qF�ƐM��0Ln�l{ej(\wW2)�]�V���[9L�,e�e���ĕ�	V�:JD�/c:���q�L�C �pӨ��7YX�e�)[[�Ǔ��0'.Sg ��X� u���£��F^��oE
�I�ywY.�%fyG�4HoN6Ztˣ���LX�[u��	��щ����5�&�[���e[�I�K�lۚ���jtQYg2hB=����I�aU����[,��Csq��)]�M=�%�z��Ð����r��t�M�w��͒��[�|^`��X�J?<�)������;B�!�MnVQ�,-�������m�[Yt��cK#Q�PȠ�V�N೛P�:���[x]���^���3��E5�R+}�+2#a�Xh���7��O1�B,�D:��f��ƬHq0᫢me���k���|��0��$��!�n���@Тm=�Μb�ddF[�Y-�Rt�o)��rV�8����kh��b+����ĕ_őH�bХ�Zu��T;i:x�(�J%�m�9����zJ���ܗ�)S�d��	�#[E��H�G�.+��+R���5��Z&�Y�S#���Ӱ���'O%;	S�5�j9�5��(b��v�an�F� �k\҈4���;m]8lZ�<`�7hEu�����ʼ�r�V
"��\���'@y�7SJ�6H�L2լ�Hwn+��v�@�y�u+w��%�la�������m��L�	帴�[r�v�a�1u�Ȣ�Xh���7n�m�@.L��`�Cw�Wa�{yl�av�G����3Jb���ʑe��M8n��&n�;56^Cn�3V�-,�h�YSIKi��t) ����ڙZh�׬��7���]K6��W�\�~�p�m�J����,�҂�v��ZثȎV *�Kl��&n)Q�^E��U�m
��;�5����iq7v�f]ԏ5ޕu�B@nP@j�0�����-\U��f޵ �rL�(���F�;50�,U��w0���R,��-��h���躰I��4CO%/��%��I[I�v��,Y���A���h���B�f��r��d�n\y�0YV�ҁir-H��2��)�2��6����)�
�{m�R�v�Jځ��[�J�8[m�N����;��+�5��-��C*���hX�V��Y��۸%��3j���n�,6(���f��|.9�����f8�B�ǐ8D3�H�a�T�*�F
ܹ�:��ZN�^��~��pn�'2�Qͦ�u�&/h��,ǈ���60�To]�㭘f��1��T�Ln��צ��ۺ���Aѕ�Pu5@���9bV94E��it!��J��0ܹ��T���/)�Ψ(�D�W�E���c�	Ӕ�U��lT��oh�Щ,U�H���V���-v�˖��;(�o+\��
�7!�J�m�e^V��yNR�ʬw぀��J�9
7P�V5[�����7h��PB��(
ǬHcn�9��ۧW&�:��0���n����
� ke�z�hd�5�蚇L��Z(-1^�C
!�:"����KX��:q1���X	�+l=9v�U6��U�:�X�-�Gl�A5���f;%%(f�k�-�� ��v�[�Na��a;+c��'H�n��t��	9��lY�V;����/�v�l�S=���`t���ÖN�d�@���dG{��@]7YQwNSbJ�7)G"C������P��Uj׌=z�
50P���X�|l�2���Vk���n���CQٳݧP�s[�.weN4%��7-E����~����A/�)k'���p�_F2�2r�2���5>� pPW7�j��:�pfl������i��r����(6v�>J�
�����sN�܃b�:�ѹY�h�ڦ��"hݲ���5��X9�B2/B�2�i��_T7���yW��� �]�O���-b���.�m�s�-E&��ھ� Że�غ��������5�t�Y`�^����@@��;'��;EEg6�N��)�oBԪ�X��a��"����7�����Ի 3�$����ql/��y'�"g$=�-�yx��;�|�'� �n>�X��vu�%9�.Kf^s��^vG]�Ny��JJ�v��O�Y"�[G_�q�/�v�Wޕ�;I���`8y�*���+�<�pN�*<��wØyM^�"��i�� ��x��"�)�$P)hO��ta�[m�vU�BĳK��K�=�x6E�<Gwiz��Lyw���V	�)Sj�6�T�PW�>�f/XS�ӧ�G��aH�ݺ��,��t�U},;� *��6JR�Y@W[��:�G�V�
��,�Տ׵�pL���*�N
��Z5"�O{�۶�����D8d|�W�Rݕ�\�s�6sci�����b�*誸�5�}�G^Д���69���|�a75��)X]�gy��O��=�v�LZ`*deBX�^}Ǩ��h�GY���N͹\�j�Y���*7G����8�7^�"h�<J���K�����[�'V��ÈU�n�'/v��M�����}k����t�㔧�VY��T��n4�"4Y	�;��W�B	�ټ�'�'@�����@��6�0h���j@�N���[.�@䪼�wZp��k"�9�[�)�ɺ$�X�ş\�X
�q�>2L'"�"*s<��^;���u��!���e]>��u�E�2]������5�jSuƐ�0�.n�������|����8ɝ��������޲-���@%�*�P�I���vvۢ2�$j��:��r�`�5�u��8�;l^���V��"�]g4��0�\eJ#x����ވM��i�R���Mf�D���~��wy�P��O�]��������r�>\��9�r\��v䜷o�W^g�fA���	Ƴ�~�{N5��8�����A{p�X�g=}���ٚ`;c��ӀݹyS�]�h��u���"��В/�n�(�[M��I��6��`�*�-`���T��)y��y �T��n�1NB�G��5���o-�3cP��U��To�/]6�,���H%�Ξ�l0t��<Y�:�����Q�s� ��.Iے������{�~J'��r@r�Qߖ��R�yR蜮�$m\�]e81�]p�t�:�ea�R�2c:�F�	t�$:��M�Ê�����N��c��\��Y��9��i��*$OL�s�X��J�Heڙ�6�틢ے�iA٪�V.͉m���2����%p!�#)�����n��v�۪�]�\�AB�N�4���s{� ���{K��.��gu]�ۮΣJe٧h#v�����9���m�41��=����9�����D�;ä�D��k��ja���F�w���+�ݖT��T�ʥ���][R^áR�b�S>B�麾��#�_*U�;s�@����m�U���.�+@E��Ν�T��Smp�$ԧ�j����{�quy0�$�����͇ [�^�}�����]G�@�4�\��������9�ʅ�+��@���|�j�
��5vI|WG�y��Yx!�'���B�Zƌ�3�/�=�Ԟ+�.��� 4g��ԧ^��������X�ګܝ �l�<wknr�%�����fd[�Tv ����u���{�����`y�?}�;�4ds��kqE���1@��Cܺ9�A"�%����F��8�H�Y�Ψ��fT7iQ�;1�1)�Uvh9OR��U�)^�%�GZ���n��N��s1�wu�8_a`��V:;��}-N҅Ar1���x�ɑ�\�3&0��u�%�J�9��k�S^�m�͝�C�YfL��`�Q��v
v�F�>���<�2�*�3뵟l��G{w8E�&�
�ý'Z�t�75b��T�[���O� E�H�0gZH�2<�;V)���QR�#���6�{Sv���f+(W�����;�I�n��pR9W�p�:������Gu�Zr�����=}�5���׻YKa\fj��3�0��6�W{է��S�8����(��ra��>�\�K�iUVs�7�m�R�;�Y�O}ܛ�ގ!�V��n3�=v��o~R�e���7w"!�;��b6^���h���\"֬��T��)z�d�^Y ��W�C!�p�.R`ҾY�f-�)E���ߊ5�c�d8v�ʕt*��,�.|TBn���u�c�W��0����i7��z�ٌ���yfPZ�4T��>�0%:�[gщv�ͦ��vM�v�py@���V7��63��Cy�s�9Fk_���+�Gih`�֌"��=Q�o�G6���%��,��)�f��{���Չw|sa��0pi�]��v�VI{��8Kʕu8+�3�d�� ������Q���/v��r�s�)Z]��u����K���oj���d�x��lhwO�o'`gS*��A'7�,yu
� ��b�IKQ8p]I��F_tR-4*���̓x���˧z��UA�]7�.N��W[R_J���9�ŕ�؈\jH��r1!���΁^ֹ��	k�k�8��&͵]�)�p^�ѫ.���_^̰�7n�d�����cE�� d)V��(�t+�e����Sn9�Q����cgP��[yԅ���"R��b��\��q��i���H����aX�k5�z{�Iǋ��{ixYs��i�؛J_=������tw@�a�ډ�>�K1+2�y�G�V>��X��D�w���)�j��z�����AfWb}9Zy�_,�ZBy�'�V���C�]������
�����B#;9�l��.�]�S!��0����h[�{k_|�s,�B�B�؎�R-�E�b)0^f^���z��^�%kp��]���	e�.w��Lc�؁�*yا)��x���x��SnK�M����*�{!a�*�Z�80�I*ɣ�c{hg��@�oo 2��]N��,D����m	���v���+���w8gY��C�<�Mv�x���ra�A.«Y�*	����/��F�gi��;5VUu�#mSI�)��r�#y{%.��杳O���������wm�[@е�ޭ;��GѨ^�A��[F<�1���<^7�!�R��<���e�*3E��V,6kpq�Z�=�q�ػ��t���̐�t]���,nn��k�;�8c��&���]��f�l�X��S��I��B�S�[{��.�u���2M�=�˃�mM������x��cwȋ�ޔw�/���WHn��3m!�e�l�ղ|�މR���Y�O���cos��#bVT]3�ZH���9�9�]����j���w[��k��a0���TO��t�B�����v���'�<�9�m���I�������/E���uv�LJx�	7��)�!Ӡ��o��*�\�z�-l��6Q�j��b��R�w����A�!U�o-���YH�*Pv�/.*X �ݕ&�5t�:{.@x�	��:vRǷ�&����d{��j�R��v6��1�^���ypӇ;� �_e6y��.����o�PE��xu�R���y��&g+w�;ϸ��X�$Հ�(��
h�g)�����I��2Ɍ�{-
�!ͺ���ʵ�O�q������v	C����,�ך-a�E��H����4v�''��o���]���֣̐��"�3�Y�zI�R��'�\��&�f#І�s�};��B�qWv�%I�`pfn��o�<�W�z4�w����fVn(�
���v�b�H��g�̬=X��*���gTϟ��.z��h�I{!�|V�)��(M����(����p6z!�DenK������I�x:1�aF��V�����><�=�-f$�FzB�E��A�'��������|\�:=V�H�vC�Sŝr=���Mv���6��3oK�A��tw/�J�U�ac�2��,9ty�}:bʅ�6X�k�t]t_;�4Yن��@P&aќ���xynɨ���j��K�%I��JL7��M�bS�e"�;��z�Ɩ��0f�nś�U-��i�2��z#��z��燠�������"��Ă�K���@���q�Xd��$$G{C������gK��Z�dK|����
�4�N�Ň���Z��Dˋ�>MU�/�P�' ޕA��D;Kwۺ2Q�ڎ����c�[��_q{� ��94��t:��K�wo�S���L��Y;j�E�ż�R���A_3n��a^�52�m�a��l��ֵ�E��d��<��C@�b�S�t�Ǎ�J�sR��aFH�)b��W)Ƕ��9ʤgh4*���橡�aUo����F ���yG)Э��iK�C-�8��B�)t�*e�%3�������v[�}�{�S~�H�W%Ѐ.65y�k��LAJZq�Z[���l���	����y�m�l�\(�	3��H�3�kF��U��K��ZC���X`.�;���ž�e{��MUAK }�vjx<"���gWK�;�|K�%��C-�ԒYlhw,wk�:�)c'� ���ҷ�`������b�����ׇ���x��D3J}j��K�Ձ�ǲ��6������G]�v�;c�5F�:shr�]���CAr,b.���©�1��Udks�:(!�ow��� �[8�՜���9u���Ӧ ���W<{��=������x�.]H#����ԋ��V���<�������w\�l;�C;��12��U
�N����E���1�F��9Ķ�H�g[�it�NA�4��I3{:�l��>����gv��(�����G�*�2J�Cv�{rPJE��kwg^��E���h��Ul]��܊7�]S@.e᧘x۳X�"��>���(���z�`��}�k��A�K5�Qՠ�������U�*:V��f5�	Mz_ǒޠ�,����wj��ˢ�:��ܰ; �V{3SWev� $����8�F+va2z�8Z>|���1;�����u��u)�]���JLw���6�&uFi,q��E�ʾ�*�q����1�ث��INUxη��ִp�C �UGV�U��UsuIq��.����]�mR�d�veSu�f�Ƙ� -�]oN�ѯz:�^SEY̷1BT�y��Ve�!D_N�-�qj{.�d<���,,Ck~>�L������rL�C��D����ڣ�Lr�7`Q�mf�B�wX���)�08�$S�9� ;�z��ԮM;�K�Y�M�����X�8�x�m c4��初��lf���A�� ok��!Iww��[��>���`����%�LS滌ѹ�����Q�(Λ��*")�ǵ�ݍ)�K^+�Dؒ�x>�9�[Kh��S|]�jN���� �\�<Ry�l��9F7܎�2x3�f�p9雌��$���7�����plVU��w9��)t�æ��[�*�Y�x�����O����꙼���]��K�j���U)Z9 �+=yj��]O��DF���.�Ή:%i�nV5 *�
<��v�r�:q�@0�E.�%��`p�R�L��9|Xt5(�+7#�אa��I������KiL;����w�!��Rs�hǮ�z*�l5�qn���Er��=g-Kr��vp>'��e�t7Ev�f骡8�]�Ί��%τ��S	q���q��x�R�̕�����K�f��Z�e��2!�	��↻�5�V��g�.|��h�|��s����$T��uw@���~��c���,�{��Su���fgNN]�I�4���=K�]��y���	,��Y�U�xE|�m�X2��G\���#�<�@��<��5�n* "5:��üp��ֹ��e��o�Qq<)�JC�旍۽r�:�κ�/(]��Lq�:���`U˾7O��ý��Z�lF܁�M�7*\�dU��;輝3Y�"'���1�'�k�-�V��U��՝�y%ft&Ș�Q*8g>�2�{)ɹ/h�l\:��q��M�2Qτ��ㆎ��l��FUf�g̺��uAC;��A�dV�Y��֜���i����}kنqM��uf\G�Rrs\@���T��c�:��.�j��S��ev^�`�4z�fT�}���[�A��h�d�9�B�Q��V�5�/v��4�����{S�e;g�n��:Ä��2���ͧ�n�Y3������3�&�Y�M/ d�w��y��|{��:��N����+v�n�f�Q�QWf���g*!��������RQ"G�-+bm&�ki.�ޙ(��X{�^n�
]~זvU�ίn};�#�>�{��:@{|�N\�wi�	*��E�[���k�&�+�U0;���n�M/�����s�e�aї�5�nh�K��Ow�X߼M���3�iF<2\qw��t�YHe*h��/�85fJ��������t���/n��|�o,<���	OT�PV���=��#��5���AW�۝�S��\��1I�v�xL1����X�c �"�%Y6M���*\%ɠެ�:�ed�/ ����� �|�|�Ȳ��๖�&dV�4]���.w�
�u�5&�Fh��b�(#��j������Ǿ2C�M��xeQ�����������J�1�F?9��e�t���.��V�������n������וR�!���]��0^<�����߹�ǯ�������m�����k[o��pқC�Y�&~د�fĘ��k&S�B����(�^������ݮYl<;Y��e��3�wOm;��	ʍ8�f���X�PCk�ժ�-�JpP�[]��X��Ou��>��kT5�J�f��:�ՂU��)� �}��V����)�q�+-����f{��W��3��,�R��m�A�̷�m�L���k���]�c�wL��Zh.�.�r'��r�DN�1r���{A;��7���EQeM��$ց`�:镆SX�C��#��92L�U�xd ˜-m�:4�6�0�d����B{\�0���U��A����	x�r�Tċ��n�o��p@s�˽۫pgp
RО�k�IB��z޽�T_"�z.^:I#4L
�y��r��h�w��g`�Έ���`[�@���5i,�)b\�˵Q�Xj���i3����K����V�MLt��Z�*���0_�j�^��k�σ��Q�c�P�f7�
��A"���Q��c�^Ӭ���gN�b[��JՖ��5�G4�`X����'�g�-6�n:F�����is	]�9��xA��+���2�
�n�qU�v��ʉ���D=͎Z��^���o����r��1z.^��$�'�c�ϲ7KWJ��d��0fb���P|FZ�@^��9q�O�/&��D�����S@��U��Ȯ敷��,^��D#�b�wn��"�'˺ӆ؅X�5�.m�ͷJ��W.�m/z�k�3�`��`��dǭn��3zڍ���J�襊����*]:��z0��7��#��|���E1)�b�R�9��1�6k|Q��∧op�9�ޜҽ�����+��t������B�r2vb��*D�&����k�w�˷A���dX��q��`��:�9;�Fn�S��O+##y0Z�8��a�S���Dv8AY(f�{���7�/�=p�*��VQ�!tGa`�/��Y����Ƚ��ڜe�o��jv����筌����6%��`�������"�h�!�!8�Ѐ��
䭸Tj��q�n��U�L�Ec�1 �M��#��b�w�|:��m�Bbf�tx{����4�.��̵��Ȉ�0vV-��N�\!�����T��]��7�I�ܛ�t0gbc����Z)t���f|�lؤ;�\������m���V����C�W�|��T�54�Pi�tM�7�lC-RK������C�Z;n�M�:���x��;l<r��]���=�pǑ&i����Z{�r�jc��염q��C1,mc��EssHn���=���-�|��o��R��D���Y���`GYE��oG;
��I�&��In����J���y��Y{a=�LS���p��ȸ�[t�h��IZ�8����2�!q3LՄ'7ǧ23y�����u��G�F�
�V����g`��;Lڀ�Ty\CC�8�u�p�:R�|��uy�Ds�;ZE�֗��b�^:p�dK��kc�)FȽ�{jh����-&\vہ(]���6I�*<�����5�@�N$�����\�����knXj袆�Ř �T��NՍ�ǻw&�	���GwT(cԧZ���v�.`&�=�V���c45,G
1�U���g�٫��h�%ۛw�	A^�z�޲��P�Tn����|�� �Cr=}V���Nu�^rgRH��v��]KszF/�N9M󉙖���h4���`���d|�bѲ�n��OǼ��Ҝ�R���iֱW���),���y֮ﴎ�B�C� S/��S�p\�j���-H�_f5���4�6��t��$1��v�c������ػx��k��r�m$�.��A��Wص���u����r	�����hrZ�k1a��
�����4�͘��[���a-@�k��Yꝅ^���HT��6`_$��t+�X=ח���p��"�`����zܫj���s��ף���ut��t�72�UǼϥǻx�ǧ�f��ֳ��0*�B��q��ܡ��;��o���g�k�A �,��.>�Z��^w�IM���q�t�Jf��B�tY׮��e�"�L]nN8g�6H����T(��YzOR㋞]6ʽ=�W�랜B�TRϢ}����Z���]�(<=���y���ץU6Ӝ&SD}�L�F��Uծ��^�>������"���T����gH���-��\��;t�Y}�w@زX�%o[ֽ��9k���&�lh�Ǆ\)�:������r� �t�m���� -͕lA��y�̀K�hi{E�=��-Ն���x�x1�_�p�M�r�I�� �wMڝ�r�Xڹ�z�m�1�!��%P������;]�Y�C)�8 �o�����sE�46T���7��2�u��似
�a[�Э���#`%���@���	x���3y�;��j+#C�uEB^q��n�A��Fv��)��>��K�/*v�������}.�̜ڔ���*f�e�ɲ��y�yhY)p�&Ӯ��8�	�+@\ w��ܺ� �9,�^ Y��v�3⒜1���h�2X�e*�������R���Xܩ��8L��<Ǝp�;8/tG�LC�|��T~rԃ"�۴�<�+�<��Ţ׵���p��j��SWD޶w%b�2�R���c�oI���	J��,ݹ�*mf�����^�X��x��M5�z�Q�,��-Tu����s�����xr��A���NV��V���_c'(�Q҆�^��<�q��j!�{�}��ܑ���>�"ãƒޢGa�t-������[X�ҙQ��&��v��@��:z�[�0�4H;�B�a�@��� �G;Vɛ�7�'C:�^>��޶Fw?m�;<��y;����o�	��ma����s��;t�ø��8�vY��wF*+�݇� ђ�L�4�͢�9���l���I�,[gE`�׵�+��Տ�x`>�	@��>�t�9U�3�om�}�ˏxi�AU3���G�k���LE�Y(fp���W��������b&,��(�e�	H��Vd\hA��0�9.�t����e�SļR����N�c5Ť����N�b�h�Wl������h�2)�C
��6��}c����g̜��;�bBu�ݸ�}�oj��k.�Y�j[�&>J���`�G��S�W(3� �S����A{v�W7��hm\+3[�S�Z����ę6���vЋ��Ϲ���l�f!�Lm<���a�ޭJ=&��C6��݈Q���Z��<:��ok��%���s��U,�fswm��W�T�!j�H�oFU�Ӈ�IyX��J܆����b�7�m�C(��:U��`;	��zAP���uv^뇛�5R'Ɓ�3#ĕk\]���gi9q�ոDpCw���������X���<�I��	�B��Z�J�1ǵ��t��:�L����\����Ʌ�u�q��i�k���.�����8��a���fp��>O���{4Ɇ���m�aqojEvOuko-�0�,��))5k�H�������Mmbn���\>2쇺沒��������l{��%���jeCu6�Z�D�G6�^���$}��H�<����_X���2�5G�0t��UJ�5�m#���mͨ��N�\G^<��t�dv���#s���_�0�G�b��>e�(�N���YR�œ4����J0vq.�Xu�|$��BP��e�,�Aж�4�y��ĹO{c����^m�(��X{���#j.�P�70��)j�m[�W�jB�7x�����>�O�u<齒��d��_�Ϭ.��[��Z��R�XQA2�%�{�ͽ���z�$�EG�wk�1�(*b�pi h�1��t��u����z���=�E>�p"�V�OU�v��޼.)���a2Z��AǱ�͋<6�
rWb(vL�ų����`�&4��lN���£�h*��c9�*� i��<)��U���N��6m躛:�6Q�p�-��Gfn��8���r6�H_x�k��>*��%�n=P��}PQ5T}�;������#�q:�ш�a��_Le��.с��3�pode39U����qitb��k�.f������©A�1{ ����V]F("�5xxKdi�X>8���h�5a��s���Qm#��R�|k~�x�O��|ң�^lW ����SJ�z!�ɾ�1O����e�զ�8���킓��Hj�С��	��:w,���6�T����]4u<I�.�u�6��m	�2�sjڲ�°���U���:���[")�_f�:�]d��x�OJ�о�����c0�/��L���0���v��6�;�Q�5�˖��41�`��pB���EV��Kײ}[Y����$DM�����^��N:���v���-�/$�؟
�x��j]�]󎈢Ϳ�$�F��BY�;��GC�o����싷�wR⇠��	�{.��L�9F���o!z�)+��e"A����|d��F�3.䬕�ڶYQ-�2���������]6<���<��Jnx�n�eN����N����{���.yڐ'�Ѧ�-B�I��$ӽ}=�q�2^�f��#Ԑ�:���*�On��踝��D!0g �v8�u���}��TjRТU쾤�!{��� xyt�0��X��a �m2ѕ{�o��_-�Q	8L#_Dym�h!U�Z����N�1Q��"���n+e{DMY]\{��r��WH��ok��U�1(" p�J�r���B�=�{���ډZ���u��.�m��N&mS�BY��A��*���KKx#�V���yOi@0BGuR�h������}��;O%��Oy\X2�����w�;̵�=��LgU�⾅��x����}Jaz�oqÝ'�=��zP���;r{�*�u��|��;2�~xvvHљ
zh[�W^n6��r�Q�T�n ��Wt�/,�ңUȬ���uj���f]ߵ�1}��cۇ�Ow��P%�nłJ
���Q8�;�ƒy+Ox`���!�0c�iE�PN��bp6��޼�`�]V���*M��1��nu��]ʭx�W1k�6آ6���8F77�]nB��Lf�c
:��ԵT9�|o�*25O���{�2�ױn���%�A�6�=�]�P�t�Z��?s�S@�e��ÃRk����75I����xT
�PևMjʫesh�/A�N]�<�z��2�v�7.�!yx0����z]�T	���R>}0�:k+lf�2e�+%��/��t���f�ݎ��v�2�8Uv���t�q
�n�������1]B�b���u�P�˝�f���x�Ss���#yU��:h��۬ӣq�Vl��A��y�T�,F�i��I��R�I����f�:���}�vR$����F�+]��^��6�fޭ�Bu3u4�"����kh��=D[*Edpڼ�'+d�I�8fT�r��n�u��2e�T�� [�y�;ˇ�ޏr�%���@��ї�������B��Zΐ�bˬi�&X�u�@:qd�)����ťHh�t��ڹ$�Y0�n�g_�����:x�o���go�eu8�;Pe^�:���x�f�ԙ�a�QYj��;.���U�+HZ�뙴��Ҫ�"	P�F��;9�U�b���:�O${]k��|+��&+%=ݱ��ej, ��{�%a�c�T�Ҽ��T��Y1���Y����l�O}&6�J��B��Ʋ�v���'o�fc�٠�@�"[���\<�b��4��u��ۓ6����O�[�LǏ
��L���2����e@����Z��n��溰Hn�[R���Nt�D��[��gÓ!�2k���Pb˥Z3^]���r��nw*��-+b�Bv����B�*��QTt�'��X���<�/���4�#|��������X]�رUmy�6v��ޟ��o;ְJ8a�9�vʸ���f��Kf��6<���i�4��F����u;�d*��m
����,�z�%���k#�w���lm��Z13y�`�����6ճ1�&�nv\)ؼ��b�P�_s;Ԟ�)�!st��95}�Od��}L:��x
��'��w���!�ۏ�w��n��J�m:�#��8�w~q.J�.�hY��w�^ѱ��i���t<�)F�A���`f5e�T���볻�R���$t�&i�1I�G{]\۸Ed�|�l�[A�e!d�����X4i�|�\6Ve���W��a�·-�LeR���;�ٸ��:���]=u��3r��F\�mm_˺��Zu�,TwЮ��҄cB9-<([�qw�S�#�P�1B���0?w_c[ݔDΛ�����Ʃ�ij���S���s3���V�ŗVp8�3�rn8l�n���u@c�('�X[��|V�TK���%z������i�;rЮ;���p褄3:��[<e� 2��&��"��,=ۦ��2Ѯb��֛�]�l7��Р9�j|bCc�>��ؗ·nR|s��ezD�{wv��i�@����\�0^&��	�7sC��k�j�"
rUM=�a�c܂�B;b�L�s�S���h�9�
���x��`#`Ʀ JkD����?\�&��C�B��z�ݭ��z�0���'Zn��Y���v�bv�0�jb;h3q䐶3T�\��E@`���qw� �]��d=i;"���?�x,�ж)�Niu6ņt�󪠆:�� z��-(���л���}jZ�t�9��5�Y+&��r7Hf��b��Vx�r��G�u���\/Aƶ��U��W[��eTctg� �����?��Fu��mK'�5�cv�-�w�vҬ7+����#|
ïBǖ8y���WOO���T͸D�DGFZUחd뚹�mk:������L(���=F��<��ڵ�����9�WiP�6D���N��b�E�Ǩ���W!{54湖����ݦ%e\���`9w8Ţt-B}g0�ח|%�Z��B��8��|)�О!��9��f�=l�neunKˬ8�M��'n��\�1���r�75I�RŐ��E��dQ�vuU�-?EQ��V�ܮ�pcd5����hZ�.��]��R�6JW���iW٢��`	҅�X���ѝ����"�|
���.Fy��p�fgU�4��h6U����Aф�:�A��� ��E��_pb��6:2����C��=v��ݭ�e"�IS׷ʹ}Ƿ��MD�%�����߸˼����-RugZ�k�A�L��U.�\0F����s��#eo,���˾��?�vH�b��tԊe>�-�gCt$u�+xWݛ诏�+�&�̔>[�i�g'�Z��J\���Axl�Sj��<��`x�}r�}�0�2�޽�`mj�5�pZ��]',��e�D 01#���k�+�F�q9�0v{.�\) ��)|Vⷴ��8u�V���Ѣ�p��C)pA�X��t�8ۦ؛�������~=~j�kF��lEF�b�.lb�F��5Z�6���6 ɬF2F��&(�TF4j��+A�lj��IQc�h�4W.F*�~��k�&�
�wv�X�lW5��\幭xW�EF�b[�#Sxj��:��sclTU˧7�'J�X�K��ش�1.�m]�QW�شh�\��,d�����j��]���+s�.1�9�(��Q�����y��}����5����:5}�!���;�u�]�ZL�B0U���=wx�R�E������y��}��l�]��1L�wn��/g`�,�}�dO�p��������f�ӼNUl�d�>coq<��>7@Wj����;���:�l�s�a�>fV����s��w���50D�oD���w/{��������%Ub0p��U�|�.q���6����n-��ߟz �uOy��50��61sw²!�5�h��|+B�\4)!�?j��~ӭ�������#N��N���T��G�}-��P��j�S�kH��R|r�Z~��?o�b�j��c\u�Ȱ��,X�8j1H�6P��\��t�\F��-zoC��t��Њ[�VvVd�u�".�h��o�6+��� �u�
y}@W1���Ds�2j',��Kykx+�`��a���}P�(���i鐆n+��,�3Qe��A2�;zq�:V�.f�%;6{�x*��І�	����9��F�] ��� �zWJ�����k��H����0ظ��Hٺ��n�'�(��)���C��Lhn�*�UJ�WT���%YlF����^��t49��B��b����٫E�"�6�\�U�e���L�(A��L�.�֝R�\����&WX�y��#��z�Ŷt�~��v�]�Z����s�
ʂ���x�� բ!k�L���:�?{9y��Ք{F�){9��lXd�C ��R�N�(u��l�8/�C=�ӗ����� klJ�,��T��F������G{�)�L�K� ���W�����.#�W��{3 Z���1���5��z0�ƹ��x���e���U!
��K��}���4!��$W�%*܀�l:ӱq̔�V��Z�U2�b㯊�b��ŵufu�N�!��K�R�����v׼"<︴���2�y���,?CW��\���$yHe�G��%N��3�p����w�jFý"҄��_8o�8Z��E����T�˨�(�qۈ��"�!���}m+�	�鷺f��Fq�a�T��Zs��q
���l���7�j�d��u����(Ұ�����_w�]�J�PV�z�^{�D��FK���T	�}?c�V��=�K�g�6n�Kz}K���O�q]���^��<�� /���ԧ��,2v�n�H��ؑco��uvUP܅��Kk>�as�t�Þ��5�g�qO��P��7μ/}p�y��
��U�O{�s}�؝2����ٚG�3�����2��J��Ou^��l�L���"�������n���s��k{���:ͫ�j�ʁ���w��$��GY�珫9��|�k�xѲ�ېꌌٌI\�E+��Q�E��t�x�mf�����tk�S#Eܒ�`�R���z�^ԙv�~��� /HU�:ѥ��5K=��Á��2uM.�o��N��@icQ�ϓ���L��������������5.���ʿ.a�j]=X���{���N���{�@�loyq�ף�����a�b=�w<�L��3��G�p��fy'���!W�v�?g1/�3N��us����/�W�jf&�Q����]'���~X�gW��3�@�����%ÞDm,(_L���藦/���W\���K4�}�=��۪�R�I��{2���B�걗�.�� /}�&�Q*�7jo���� �=���HH+�B��E_Ā�Y,`��`�x1�k�u��w�^��lm���/ש�P��d����4:��y옫�H�iUR ��촩�^d`�)��U�M���x�7F�2�F��l�0�W[��h���<��ۦH���U��:�Y�t�p�6Z�7p;�!�ȍ�|r��(�9�u1M���SNN�{:ކ�\D�t�6�|gT�ʥf�v�c\�[mk?)ZqP\�6㲶v��Q�RW��gu�dәP�h��0�MΫ�^5}\���]��

a�oo��W]��z���O�A�j
�G���$�x6f����*v~1��O1���8g^u�V����x�骉�X��(`�"��[.tO��Ϋ���iR'<L,�v�o�����),þ�{'�o0��"��¼�xA��i���b�T�Yb4��yu��&�9� ��'�d)�;p͇�����{��R���������* W�j��t�a�R�Y�n��]���߃�����b5�~Py�V�O����i�#CD�����Kkic�+3�؇�7>�s\����cs'���f��|�5a��������oE�4���r�n/�u�M\>*�k�]��)�g��<����h[�̉U]����SK���Nu�.@��[0E��kN�����[�ԇ��hP�S��O+F�k��o����9����x�h����>HM!��щl8����[��x\71�/�t��3�خۅyr�����N�O���z��3Wr�X>W�]�&�N���Ϳ�q��7ط���\ʖ���J�{L[�\8\Jδ1N���J��t�Q�&�DP|�!i� ���xk]z}�����[}N�MM�&���A`zQ�d߅x����ie�{zڼM�7��ڢ�4C�s�^�N|a�N��yr[$b�d��YԹ�ukNmhI�b��z�f�7|���/^cC��k$շR�F9ЫA]{��Cy+��oA�UIZ�C����1�sJt���Vi�!T��d�*P]�t/hS/�=��沨���t`u��a��Y���NP�p�ב�u��q��
�3|�Y�MmM�F�1�{�F�z�9���(z�/~�5�	�qS��]�O�JQ1�d�v�评�w@v�Vdoaf�L����a�W�>��K��R6<�`
篺�
Gk���V����f�V����y�ЕT�y�Aq�Yϸ�Wp"P���1m�[;���d�l�z�_*�vsj��сu�FJ�7!_p�U-��{^�9�h0R�Wx��
�Oh�S�G�h��f�6n�6�_ JwNJ����#E�(1�y_*��d5#4��x�L���s��f\#�j�ϯ������GM�uZ�l���Υ�K'p��H.mx����'��~����~O%���*���}�Ԣ��<����{�kH�p'��n��jB�;	V�9��#E9ڄ*��B09�@���1H�Q����z6V{'�*�ޓ�<�6��m:!:�o#}��xMH��3�R}��U�'
 |�����\��t�`0J �E�p��']U��ŝ�����zOOY����h{Jh-eྒྷ�`�A�'#ݮ*�9����0��Ɂ��̄f����NEpcw}6��Z@NάV������F�u���/��\�C> �uX�����g���`8�	�.?"$��q���-w-9y�Uq��m{u�=9P�U_e��j,���!�xg�t���`���2r5�������,Fa�;�n3�o��îJn��L􅄣�C��&*SN�Jy��k*%T��άM�QznL�9����x�4_9�^l�(�ҕ
�h��3\acc^���í�t�</&Xw��Z
�ca�q���L����(:��z�79f�NN�x]P�@,��T� '�SȪ�B:)��I_��^��#'n�ۓZ��h�(�s1�7w��;��������6��[��Y���v�X8eR�=�u\�&��
����_�B��
թWs�ׅK�U����w��j�:�}�A�X��k�r�e��]ߟ9MFYoV_�:�PԐÒ䌎��4z�?����z��Dj�������r3a�u�E�'_S]PŹ����K��˃_<� I��t�U�!��T�@t~��!y/5�mB�j�w�2w/����E��i�\f��e�
��Wx�+>)˻�`�k6�vB��5��TLԖ��f�z��-`�CB�����c��e�"�LG���y�x��mB5TKd�μ�#��{�d�mkC�`L��g.li�#!�'O<�x�c�p^ʎ�P��f/�������y��t�`�;�R�y��I�� z��.��%��Us��-��T�u��<"2\�Bj�����pQP5��Y\��Ν�U���KR�}�Y�L�=�Q�gb~`�u0�)�Ȩ�Ɠ�3�qY��1����OeP��+��(�}�NE��̪�/�4Ī��qb���JUah��;�ܙz2l�꺢�.�M��a���}��s$v��C.#+n:�2]�E�j4sr���C����D�x݁_F����9�D�5�e�{��h�¯n+v/��9�uH��[�����c[�,�s˺�C�w�9u�\��$��lo��o��0j
WRa�bd�>�"�/s�{a�{K�j�J��ɞ��D�)l�m�|wa�����1���v吶�|�6�pq.��*p,K8����gu<������K'�2�{/L_����ݨb��qK�N�)�27��l�@y��SwUs̬����ʅ|UG
f-��鉘goWCA���u��}�'��p�̞���`�t�I�N�xP����4��^�����^�}�g5e���%��mzjm킲N)ң�dwْK����R+�9q��k�r(�{Sx��.���/e���}�a���X���$^�M%�����Io6wm�}�m;߽�3@l+�i w'�N������\[��ڄ���F,�A^��)s�����g!�!#_[��Q�.ʂ�6`�;u2'�^���.�}Z�u�{N����֝����N�59���9:U�<�-L�G{�	V.��+^�iN�E�?9hSYN՚�[u/����=}�U*���2�j�U{�QuSS� 5b=�g��i��9�n����P��Rډ��𘹃���Ni�zC�bF f��9��[�Z3�[��x�V�3+M���+m?+E�¼���Xu����^��I�ڊ�̄��rE�&]��6-�C ���O�xn_�A�7����i��1���f��q�d��[�ݡ؆OR5�K:#�`Nf�qm/��п:�3�k�:����.�{�e׵��n?{V����*�#r��?��7,/�~��G&0T2�ʋ�9Se%ӂf ��w{�ˤ��S�b��ʽU�c2�	������<'�Á���~�ٹY�M��
b��r�q�4ʾ>�+�#y1��ʯ���Ï�N�X���:+�����9lJ��c`���z��lN8����PQ��=`v����'R�B4q�g��'z��}�6$��7Zz�q"��F.��e;9_�Ӫ��C� /����n����5>���<�����D(2C�Wj���a�6��&(F�N@�<*�q��,B�/����>aW�����inKi����|�6'�{�mgޝV���b�j�+��=�3x����~�f����@�3��3�͠���Y��}L!q=���u������|�Q�f�vL��;��h��W�.K�J�_HX�f�����l^uPF�H�9�w�V�Z�xG�&A6��K��?J��{�?�a��������cAWE�	��|���(�	��B���8��r�mJ�%Ya&ϴ����5B��v�x���b�4Y�Yd�w%�I	<+���Q�*K����g�޺���ٿ�\c,t��;,E#��ϸ:�8�z��maw����]U��t�&��,0c:MTg�z�B㾬�=[��CC~��\�R���~5�x]����w&Y�rZ+g*���������n��D�tB�u�kJ���N�h�j���^���q�u���%�l�f�;����flHmт�SJ�A�x��`�h�b�%vr&aŷ�\cf��+0@̝y�k44�ǞJ����r섄�.ɳ�d�ْ�8ܡù�.�Ʌ����#�FFະ.�9���LPq��u��r�= �VlsJS��*ؠ���,8Z =*KH� ������O°@�EN?���oӸ���ou
Q����2�J��iA�WR��R}t�'U��{DP� u%��}}+�˝5�T|/�L�#k(Y�t,lR���*���=[�v�(mo�0�{��O���T&U����ˡ�<�����{��VxW�l�8Ģ��`/��FɆ�g�ة�{*ƔO�R�]��͡��tw�`'���#�-�ٿ� 1���n*�{>L��v�������*��Us^]\"�^_
��c��#���:��ᖗњ�.�P7�h�C���^ؑ��8��iC�r�/0��(h��h���
�Jm�T�J�!�9p(�k�-_;�>1�f�M��%��L���4T@�ٌ��=oh
D��f�
�����Iix�����􊋝�b':���<�1�҃���u�F�2`Kx� c�F�^rx�L�L{w&e�L q�Uv�1NpEF������0U��]I�<���b�.����b��/��'0�@fflm�8Q�K�3i���B���>�9�Eo�0Ws}�w{���m��T-�U�0���T8+���l�m�����vR[*�%���`�h��U�j���TJ�ƟدSc�{O]ϛR�4��)!�%���SE.��7Б�²�+,n�D1V5�n�'��(+[V�}7r9s�l:�iϹs�2��u�cq3ռ�,�t|J
kdՍg��2;w�Y�� V�2�V�2L��t���n�^���_���-u@z�3泺x���t�<+��'�C��v��S"�t�Rg���y�Ý-�]5;dc8���~����I� �^�E ���y\���V��j�GqF����U�����QSd��#l�	1S����Ըp�� ��<�tE�k��5*��Ԯ�l�*�may$7���$��|'����ӵ�IQ�sFAxN�w�śu9r��oDn��I�v�ͦ������B��:4E�duu1m��)!]%-F��
^]�x��1jZ�"�E�*X��ţ�гXBEX�]��an�5�n���|G!Դ�wI��̷2uJ�	L[K4=�S.�a#{�)��ӎ[�͂豩C���cc4dFL��a%ml���WS�-3�V�uD�������O\qm����kIy0���L���{�к���H�Q3��.��Ȏ�l� f�7�8ݞ_�Zs���ZɤӤ>���Д�{D�ճ��c�-�X�=���1<���:��U�����X�ת�;�Q%������i�:���+a(a$P�:-+�
�&��>ս�/w]�R��h�^��+��z�p@�	wY���ł�6��Ui.,)��}R�V,^����4���oi�r.rj�Y.�J�]�Lq�]ހq�ΐ
����F8� �F`F���QS@{���{O0pӹR�@�ݽ>��+`5�2Z��v�"g��q��Uw0qi ���ޏ�y>#t��[J��^�Ti��K�.���켝��`n�d��%�. � ����Ξ	L>���͝�; �'sD�w�K҇��wx��5:l��.<�AS</*~�\���)�3�dm��L���SCs���1�
T.�-CT�.���M����3�ל^�2����e ��Fl�r�r���Z�=��^�F�>�k��i�����'*�խ}F;\�����!�@�,m�u91���7UUWB�F���|���	*V��^N���]*�.�+���,�xs�^h<�m�G�uぎMmɗ���T���h)2�f$0Ѣ��܍öN%�q
��>i�Q�=���T,�c8=��x�gz�F���������-��mC���V}�"C��\�W+�[D����I2�(-��"��6���f.�Q�7�s��Y���Qo;�(âI�nZ3�^��D}��@u5b�j��Jr	�J��A�L���X�����.��k�?,���(AA�u����9;�J����m��i �2�so��> �� � �4j(ƱF�j��h�nt�۝��EPPZM�xs��(Ů\�k���h�ţxsok�[�(����lDF�QFƫ�u��U�;ZK�H�E�E�����[Ö���T�VƮlQ��x�ںW��k�·����+�׆�-s�����Z�t�6�-���r�4nUȱ�;��5�ڣ\��WcF��NkܷwEwn��.DQ����E�@���2��F*�e��4Q$
��M�F������p;�/�p�*@��0g����#+r����To����!;뛧���{��o
]�����������/�^�y��V������oom�oW���G+��_���*�����+�W����+�\������^��;^���7�ܫ������7տ����_�Ssc�66����){��P���H�}��~+���{���W��ۛ��>5���h����5�sny�Q�׵���z��k��W7�����zk�~�r��+�xW�^���V��[�޽���D�-\�Y$���F��{�#�E��1x�ו������w��o�r��[�Ͼ?��_�|��o
�W|��^<��
��}��zW+����ߕ��6����x����x�����������ߟ��f�;z�����C��">�D�z�輷տ�������KA�[�_���U�^���^}~�_W�zyk��_>����ۛ������ͽ-z���y�ܷ7����[���=��y��ޕ|\����^��r�œ�w}��{��0}#���A?>��S�������j��Fܯ�s�_��ύ��^��:�������|�Ԗ��������_��W��w��5�W.j�}����}o*�*�߿>=�Ͽ}׬T\�}�mo�"@>�"�z(ň�-��_��oŹW�����}[���o��Ż�r�w�k��ϭ�_��y���¾-ߗ��w�����oϿ<m�sn�|��G�^���>~�~z����5~5�(]$o<r���}�>�#���w+�����xW�����_���W�������U���h�����}��+��W��o�r��Z5�������}U�}W/Ϟ�oMzy�ڼ+�*��ǲ�IPlXڬ;>��A?���#��o���/M�-={���noCQ�_�<b�������_��^+Ҽ5��o������h��x~_����Ϯ���o�rޯί�}W�<��w�^�6�")F�W�į>��k�}!���} Dz"��y�[�o�r��������s��m��|�_�xU��z��>���9��s_��k����o�:�s�ok�����W�|[�����z���h���������xj�x����n9�2coSͫ>��}���={�^���W��7�~*�ͽw���~��x_Ϳk�����������5��ţʿ/|����soWߞ?W�x[�����߾���ջ��xm�|W7���|�k�/�d�.�Q�ޑו�&kg��M=� Z��f��pk���WP���*�Z������x�t��Wn��~^P�z�*��qQ�n	�Ӆ[d.fcGs+�$���o�s�b>x�K絾��r�ۈ{[v۝=���1|��<;.�)�o�^Ү	{�t}"#�F��1���������m�y�{oGֿ=~��|_�|k�~_?�zW�}^�������ήoj�������zZ6����^�5y� ��D@0�}"D|]wp��n]��^��������{������=�W�o]��o����o�}[����+��������x����������{W����߷��_Ї�1�ﾱd��r��s�|%��������ۖ����r��^�����m�xok����ү�͹�ׯ>7���������U�nk���*��s������|��[¯+�kߋ�o�o����}"<>�	���K��f���,����������s�o��?}_�z�+�������޾��h��T^xn[ߎ�Io���-�������J�r�~v������;o���V�{k���/��W��ϻ=9+l���Sr��|v'�1�h��5�}��yW���������~-��z�}��k��U��{���o^>x��_�x�⹹���*�k���ۗ6��x�^�M�x����5��<5�~uyoo��$}p��6z�W*{��nv;����ѿ��/�>����^o�|�����6��{x5�7���?/߾j/+~����^>6��o+��וʹok���5�~�W���b������ym��">�Y��2�:58�ݟK�����}�-����[���j�m{xW�ν�k�Ѿ+�����徫��o�|yU��oj��|��/���|~���J�.m��>z�7Ǖ�-?/�|�o*��7�?��ۊ�?iÛuw���#�P��]�_:�-�W�_|^Q��7�n~o���m��޻�-�\�כ�ߋ��{j���������޼���<��[y��xo
����{y�~���
�~���������0�l���J��E�D�?|[��+��߾{^V�~�;�o?z��i�z��_�z��޿{_�}[���~�k��_��x��Z�+���<_[z��^����澽��������{�_S~��I����>C>��B�#�4y�~y���~5�xo�^�[Ҿ���׵������o��o����-�E�����U����_�s�\��yW���ү���Wz���~<6��n��^����%��xǉgl�x��nN
��6�qv���1)���Y��}�l�ݩ+��V=�W��|?*	�r�y/�3��C8̻��c0�R��	��(je��4���a{�n�����$�	.�0%w�r���S8{�?W��zU�}߿?�צ��}��~�~z�xW��_���?o�5ynm����y���x�}�⼭�]��\����������z�����o��������soW�oo�G�":;ۆ2�=>��מ�')b�����W��x���~*���߽yo-����_�ѷ��V��|�ҽ-��}_��?�뗥~-�~_z/�ۛ�[���������^|x�[��ߊ��>�"!����5���x���oWN���xm���-_w���w���x_ʸjJ��ח���}[����ҽ���~�|����ڼ/˿�|��h+����z^U��
�?����k¼
�[�}�D�|F���T���j�������}���h���{�����[�z��-�z�֯�޾6��W��ʿ+�[�|m˚������Z
�{������yk��x}U�_���5�����{_�F������$G�G�7�~7�U�3�>͓���[΄}���^���z�nQ�_���W��~/?�y^���-�:�5�}U�����^Z�����*�+�_���~>5ssnz���W����x���o+����z=��(�^4rn1Wl�S�Cj�~5�{�������h�7~��[���k���Ƽ��-�������U��z�_�MxU�szߝyk�~�����׆�[���W�^V�[�������������H���� vQ�W��V����������uyZ/��}���j-��z����ܽ?��^�o���ӛz�זߝ����m�;o׎���^z�_[���\�r���xU�������}Q=6Y^�9hp���F��ߡ��@{��^��o��ߊ����xڿo_|^�}\�ks����ޖ������r�5�����znm޻�����nnk�����u^��.^o]�"���M%p�˼�W�_�`�4F���p��yj�}W��z����/ţ|_����r�]����[�r���~���ח��F�����[~*��n���=��������=�������5ϟ����SV�"�ϭ��>��>""�H�k����������k���Ϋ�����\�[��\���{����[���-?o�<�[�����������s^~���^����/�?<ޕ��
�.�������_���S�H�3���k�3 �����J]�����HX�C�i<}
��nXԱ<q�WݻuQ0j�0ȲT\��#%CUj�J!R�W�U�a�pͺ�1��ah\�*�#H׶�*�e�.���b���n�>�N̴�-uX�'T�aww\�ﾪ�Wҹo�x�6�n�z��y[ʹok�y�����Ǿ�ռ?|v��m����������=⇑�=���i�7�tȇ���$5��(}��F8Z5񃃺S|)3���{M\����OV?
q]����]
�NW([�pb��uƹ�t���(U/j�- ;�x*O��&̱0�*���Tar �W���;cRUh�'k�(��s��u wi��ʷD;��3˯����-ԛ���lgt�b���L:Iٳ&��|�h
|`{��:�'�X c����,g�8��O��{�]��}��L�iA�%f�����oT]q��U�TI�anS��*���c؝oq��Ró�UEcy`)��l�ׅ��e�;�ӊT�^R���z�1�l�r-�t�z
S�$G���b��/J0NE�8a�4����`N��gES}J�_^^� E���_e���˵\�#�n8�=���Ɏ�=GB c�� �l�;Ʋm�Y\�@qc��W�*9�p�q�M|��a?n�bb���k?mK�m^O{��z�\����lW�{K�ܭ17��nzl�j��gY7}���Tez�+	�h�r���s�Tj���^c�`p��1��:��,n�F�]!j�k�Cz�\Μ4λE:�W+�O@��:[�/�-�(}��wqo�$K�eu��sQ`�Q�U�q�cr��*�����h���݄p��� ^3F���7]���6��'�(~�0���2�/��2��_Le�u�����
����y�5y�6�l���%uHZl�̧�������8��5�g��̽5)+�PFNUt�L�-�l����U�^lJ�ܪvU`a '�2�F�L�C�����!}�oa�w��/_.P p��B�B���?$@�
[hx���Z=:��k�:�f�L��}qO�F�Ltb���	C�' `�����f�f���Y3�@Nz�|JGp�2R�YbGNjt�)�#��6Ш|a��n�ϓ�8EE�� A��em�_c~��Am��<��l�yĺq �;�"	xk�W�Þ�-��'%�g���޶� ����6O]����g�s�)u����C�0��X�h܀Pʎ����Ѫ�?{��R��"����,�sɞ�ؕ��I�fLp�U/����6L!���KQ�VJ��0����O�S,��D�R1�*�%@E�t�o�=ůA6tM�u�c$wx��k�f�q�v����Ѻ�})L���p����pJ��o&�hgbN�f0��寠��N�]��=�S4j�ˢ,�"�S����+R@��o�sSfBB����iw>��",��T����в��źD�5q�z�ؘA���V	ڻr�	裨X���m��!�\O\)��T'�q%s'�o���K�~ұ^�!���З�9]F�y����M �ҝ��P8X�2rpN�ߜ���B�r����P��&\ [o�r�yF�_��g��3�P�,k<]W����Dh��TXv������&j|=[^�epS<��W�ղ�R��������l�Fr�=�#������Qf��-�H�b\ׅ��ի:�E�ee`=�U!�bC���7�/���T:㺛?_إ�����s���q����	��E��;�~�hCx��|�x�p���mc�<&��c�CC@;2m��Og�����G���ގ�69VO�̾S����@���y8f���ץ��ڞ��o9��/D�D�@7%��t�����d���,����1R~���x�6�c��P�TOJ��gK�B3�}_�z�;���+ϟ������ύ�c�w��ܗ��{owp���1E��ƻ���>���zz��}t.��ؕt��h���h��f}�l�P{�q�K��m�:F2u�]O/5ñ��`�H��ʥ�=��#����U���Х1�ulQ\�h��X6��u�/IΙ���)%4�Lň�ѻ�%��W3��Ba��+!�0�ݹ<.3}t��������+}�Һ�
LK�S�C�T��	���W\�s�l��L�*����ܙ¬����;�?���TX>�x ���:«��x�pa�ba��e�3z����K��3�Q���X�6qR��z���;(���S�]���9A2O{0$j�%��V"�P�J�}���c8%�E���;r ͇��7jl�&�<�;hb��X)��7ĕ��Ȱx�Yvv�!�)��F G
N���h�'e��Ɇ:�s_;5j\�X�y����2Nt����.�J��G;�o�F���o7G��7*~��ƹ�n�G W%�\iOm�����:������6̪Ss ����N��q�Gax5��]�jɢǭo6��j[G���T��ȁ�D��W�L_'ecC�+rp�]��4�Y�i������[ݙS˵���x3�����>�UcbU�]g�&�s��������KF���y�Ue7��.���jE��ԾA�B�&��������6���B�Ia�]�9;��%��kIbu�7���=��YukO�)��5��ə��lz���t��X"9du;ͬT�	0$�<��SR-�\�3e=���J)v�L�nN�v�#��#>���]���t�	��U��un��uqWP�_��z�\9���Țy5[nY��;.�+-:��4���r���t��Yע�9P���}9=�]3`v_w�߆]gVc�	竽;���zU���#���\!��m�G����e�TP�F%������Q]nmSԍa��{���WWǙ�ԺH�q�����0��L#4������ۭj.�^�UCl$��O���b��R���KW�u�{�����I���^�\�(��f��m!�"04��s����E���5S�^�(:�%ۜr&�1h���@Xօ8�8fƂܠ[̂*,����5=�2�W�biun���c0֘[q-Kg.0�6ʒ{�����Ά�U��9�b��0��ic��a˃?!�n�w����#�����t���߉Ha	}'��߼��z���![�ޏ�SixU��K�׃}3�.g&��f����ȌcY��:�ݣ~]&1M����g���<�;���>#F�BmꙞ�j&�,�mUҧ��z��²���5�xv�ud��-gZ�)fk�)\��*Ε���'h��Z"$ݵ��:��x��$%�˃2��T��SeZ�.��FL��n��v�`�.��!RMo�>б:�.P>��ܬ�"���ک��ƍ��oP��>�dW3N
�#u΃5������1�)ڪw�~:����>����R�W�f��:.W�
R�ŵפy��j�|�(���*�O��΂��c;}F1[��U����c������kEw��9)c�-V��� '�2���ū���$��|�_ !�9@
�J���:#��C0�$ݞ=�80��Alem�ض�p�Q�U9�I\)����Q
�F�ejv�za�Ζ#t�r���'�]�����`�a���5�������3n�L���g�T�VK/ƷR��L!C��S�p}d�u�ڜ���ROv�����x(Ę
��!��<%U��w��Z
f��2�7	����;Wd<�x��]�S�0�mCQNͩ�vUX	��z�ǝ��I�X�+Wl���Ԟ!��:�Z�=�kn��6�r�V��1����|���J��d�2R�M��8<��]uب�U��GPy`���OF�%�&S����FED7L�-#"9Z=L3�{e�.eGG���o�Lt[��R�gp#|� ;�j��=;ƌ��E�>V�3/���؂��U$�c��;N��t#�t�����X|��?���t�C�z�v�[%9Iz�Xձ���["�#�g(��ч��,;yq�WT|��'��W�[�N� �M�^l��/�+�^�ZbvG�RCK�8�x80PS�o,��{�je���gO9/�5����w�������S������9��5�t��|�Ys�FVS\�@]�:��_�v)�S
�����9�^�Ms�ҷ�c~'禡T��e-Lۭ6�G5��9����p��`���uڨ;*/E�8X�x|-�k��Q�6P���Q�ʮ�/��Ѧ�g�Q�D�$��#�9�?��vk�Z�ay�MW"�0^��2����R��9���C̢���d1Ep���<ka�:vaY�{_T^N%�ڍ�:�eq���)6�&��\ �u҅���g0ȯ��2����c�$i���J�9����Lmޖ�q��R��O��i����kc������^t���*4SYDn�H���3��괘ų�xXrt]���Nt�20��35Rd�^��M'�(�V�*��1d��w�K�ts�R�|{V�n��������Y���I�����5/Nw�Qc���lP��uh�Ò��.N'p�!E�ce*�X�Z���ya,���N�n�~��8�X�g��뛥�I�K��������Z^�p}�G�����<�T�P콪q���Ų���8��k^(��WXM��x�N�&kV��+���UǸ�:2�5�&��{+Gƙ��5�+���<5�O�BVZ��R�ڻ�@:��n��x��їY�M\ӓJ��(�UFQW=�w5��}qYٯQ#D�ҭ���7�|Q�1�3qeAX=A������Ẕ�&��j�l�N�|蓱8c6��8UzIݚ�߆�K<�Y�K.�ۡ��U����ߜu��NKV�a��3\1�|��ި:���L�^A��;γ3�	5C�ެ� )7�R0mK�G�g	��4��tm���53½L--=K����'*-WIܵh�֧s+����Uf	|2:o5댡Z�(>�ܒ�::�"�}6�=:���g	�Na�t
����XIĈd�]b@w�#qB��"���}�.88"��F�s�d��GU6�=L]'�&t�8�vC��}8���v)@q݆a�&�����.M;���Q�q�.�J+�ek��^m�Yb���1ڬ=� ]˗�>G��TX���*ޓ�E-f,4��MCC%	N�B�Pd���S��7��&��x��b�{*�]���6,�#F��3�W��48��5e��l�oJ�ѠK�0��b'��:^��=����� �d� �����G��K��^ �J,�Xc�{j�#@QMp��}a>�L��};EN�=�A�A���EP�i��&�`y[�u�8�s��vEj�*J��Ls}M@rOZ��^�C{�	@2�0U�����CY��Vs���kZ{(k�)�1�swpm�*J�u�-���4��>$`d�&K�X_r��C���]C�P�]�잙.P���F�x$�1;V
�%���[����N]Z��g��JB���_�m�<�Ϯ�d �;qB����p�K�K7�p[���r��in�z��LJ˻�ZK�x��g#F�
�.��L�����\���C,:P@ЛX��o�ַ�PP��Y.��{��􂂧�n�#qYb����p��ޖ��yP��.��bK�q�w�@r�SF`v�n:l��-��m�C�Ӵ''v;y2�)9�N`����0Z�|'h�	zR��e��H�žɋY�����n�����V���Ѡ�N�hrRŚ�e]��H	��iӭ"�f�X��^T�.��D�½�>�woL�'f�q��m�Б��[Wz��#uP�Bӂ��Z� �1mc�g��Jz�R�M�z4>�t�������*�l�C6���jR��cm��+�;���7{����l>t6�ST�]��˲��J�7!��F���t�;7e.sE�n�f9R���d�u��M+I��lSmؕ�fe�Ή���O�UW�Q�&�(���.k��ͮ˖�F�	Z��Ȯ]ݮl�wm��s�9���1cE�p��.Y۝�sh��E�r�J���ws\ܺ�,Rnksd�nȍ�;����+�,���m�S��+�㻧v��j�RDh�79\����t�b�H;�f:.W.pn��Ms�ݓ4��p���E�6Fs�����
L�14i�v��W:TJJI��`w:����B;��������K��Wđ�p�'u�uӮ�$0Dh��0D�ݙw]!	E	��ӫ�2!A=z�<z����yƺ��-�&���� ss����J���z�xb}zj��iX{�hɀwm��=괡K��	j�56����f��cٷ�Mr?��1�����0aN<���SY��ZU��K��C¤�NL�յ�2j�������H ��>1�3��K������̾S���/�� ]��R{8���=�bv��t�wJ鹿�>{P�)�c1��8\��b���*���s<1r~�6����[�x���t'�F�nWݘh���;H�@�d]͇�.�Aa�91:m�8�^m��k
ѿZT�]���f�Ư��_�3���8B�N�q�,��6	x��Uoa�_��rգ��r�\(��묊F��Oa��0���d;�.����L>�{·��kl�x{���z��8��U��j�V�HQKj$b/h(eA��0��hN���v��0nEϳ����z k*�Og�}<f�t����vJ����m���$��\���ZiС��y6�C,E
�j@n�:�G `�2Q��X�6�ډ�[7URX<c>͛�K�|0�@�Q��]��T�c��b�a��l���C.'����ό�'6N�\kƆ#&�OQ"�
ӒM�a
�z���x|����y��Ǽ�h{�B������@X+�����;t�vVvXP��Wz	��V��'5���t@�Y|]�q��Sr��������'o��x8*��Wx���*��F�/�1v�[�">��g-�c�F(_�kó��R&MF���N���d�t�*��yT����|�At_��R-��~�A�-���ć�2�)�u�l�)����u�U+5{<��>�k
P�����r]Җ5�@�>�4E^ϕp�'�f$lb�1l��c��zs��b��J���I�.ϳ�Rw�zc�O~�y)�Q���>�#���>E
��g Iy��od�T��;`�u:}%�>~u�.������m��;Z��q�K~���mq�@��S·���	OaE��:��Z���3�X���p��!6@�_)�)��hN �Z,-ҖZ_����TENWA�ƾյ
��i���6ܱS�3���(��5�W�̅�]J�_n�fLa��6��������`{��f)�(h��v���C"b�W�|cP���9_�u��R����IS%��5�\�)�Q{�__����o>����z������&����~��"`B�8��1���q��?Dl9������<m	��+#�LC��d�ީ���[�WZ�b�����\���J��ۮǊ;�7x�	���n�#�.�G�`'�W�{��Ʊx����G��q�[�ǆ�{i^HI���M�:�q���-��o|��"] �u(��("�U������.w'C��+gDz�
ϝh
�-��+�(�4CS�2Ӵe�oL7���3׮ ��)x	�};�Cy�	�"~�17�l�9�b�� sw@R�RD�!�q���E'�+v{�?Dަ�K�)�ٕ����J�UB�u ��B��"� .�N�|��'�Uz�s"�4��A�2�+�W/L�CL���m+5�G�b�qS���HcGcG,��mwNV�9d��p��[��ʣWg�V<)��[�&7��1���aeڥP�G���^!K)5]/'a�0?
YA�u��ī��< �����������o1Y��yu㜌� >�ր�atc������kC�7捜�����k�{	5Y�����k���j��i�P��uW�gԼ��u<r^[��7��Zj��툴Y��;X��4�g����I/��C�@�l�Tf���!��n��Co��a�7�������!ƻӛ��%���DR�{�+�֖�5��+91Ж^�nS:2�Ɗ{1�h9Vg���u8���~�b�[oD|�[�w���CDî�p��D�K	��X凅�vn63�7��=1yA����i�������n��aF���Ʋ+�l���>��U4��z����Κþ*-�Erl6:�Kv���Ԯ��UW�}T��m�k����?�m��[�F|�|�i/i�d�����@S6-�,�/��V�uJM��u����/�X�#D1��S�t�vU`�*�i�+�R��+=k'��}�n�dk��f���蕧r�)��c5`���?wN���w>&}f�z�|`d�hy��r�����.[�������0S���62@!�WNWM	��S�~��E�V�]�����TC��s>��	�ݨEL6Y��w���n�
J�)��1����ýu�Սp;=�w�tQ����.[9�@+���V��W��p�9�F��5 u79r4�:,�Ѻ�t�gu)�X�Wt�T[�!�����@(g&BT��2~zl�fvŢ��⩍�{I@�r��}��r��R��n�s��c���	��<=W"'���^���q�V٤ja���c����4j{�I�C����-�&C�kT�3QQ��h�Ke�Ü��c��Ƌ��U(���̆V+��5Ğ7䎛Ŏ�̫�?����U������ ��:*��]�s
��n����:��u:��s�X�"�1�˴70�L�S=:�l���Z�����t��;���:I�Sm���ʘ�O�,�|~�^�1��.p�$�{��nVT��>��AE�v���s8�8:�bc�*]�Q����D}�K7{�o�#��w���� @�X��U�L7�+vh[s�E�+��)��p��ho��s�;#<2ߪl5�*�oLF3ZT��`TYcҝ}����Jͮp�sk�����z������*���x~����\���0a�&�om��S֓
t�X)W���x�s!��s`��SQ1AV����f�Ү����w�=cU�u$zy���ჽ^[��l���2 �_\+���)�9��-*��\7ٚ�ld������:�8��V�CI�a�p���{�Q۩Z(�D;'��Q&��������~���ǫ'q��;���[P�#J��-��>�8\��b�,�4j�V<���7ᗾ��%j�c�>1����|8�cN{Ú���y��w�#�>�#Q���h��� �L�V.<��t�\o��s)ś�������χK���9���_��P��|i9��Ǳ<1�\���st[���s�^p=�	���!ׁ�n�J�m`1=  �mhnR�0K9r�GoJ�bNmp_�J;����C��KW}Σ�e�b��]�,���z�p�.P�����)���csO��S`��h��q��m��o�ڼ�H���M��Ek���Y�]H�y��)�*�t6���p��utښ;�-�������0>-��1z�tSa���o�]��R�;*_Zk��}��w��2�	���%\:�}*z=���:�/�nP�`u	��+�㎊K���e��6����-DINv����W+RgonZ���bíV)��B��@>�5C�p�?CN�w3�o�ry��������G"����u�o�#h�{���ݲ�;�#EC�a��e7��&�[k����o\4��u~�9�G�WZҵ_�vn4���}� �S�y���2#����m|V�Oˑc5�_��{؝��P&�x�]R��rׅs��;2���)ZP*�/w����Y�q+1[GެɽkXʦ}sLNl�1�H��ԑ��������W��X��Y��/��O.]I��'�>�w�r!^���f\�Ƹ�|.��3�U��IWYcY���_��kW!P�e@�Dh����� !>꠆��oN�\����[m��qLvÕ�_	��w�׮e�*]��͋pHh�\�G#�W�Pxn��v;�S�
cέ;4u�\��hd�������H%V6>*��N�h�̚n�\y�<}x�8���ƅ��l
59�&-��RH'���pZ�+�5���a���Ε ���6\�ޢrA�Z�M����pܳ��W����O��I����k<�ӑ�~�����#�����=�T�~>��J倇�c�i
����b`-E8�hz�;��
��l�tb����yZ��F>s�p���dE����U#k�T������,`|�$a���5���Q��;����4u�r����R1U���$�^�����C���S0scp|ݾ��"�좗3�aa���Z.w�tp(�d��D:��������+�c��(��&����:�,��ֆ.WSq��z۽\ĉ\�-Hjw&@zj/�|^����v϶\~����n��P�s������;LA�1��H
�UW�BS{�!�1F��=+����Q�����Y�E����H��j��zd&��:�) A��[�7,a��sC����Γ����#DHb���r��d�╁�W�M���W�C�b�:v�t�c�ʤ���Ρ� -�M@H�ė�(��c0�8��\�3Q��ާpÐ��-W���ٰeW���������5+}Am��B�[V���~��X��]��(=�'!���ql��8�����;�xR��9��EmQ�`����lY{J���q�r��h����Y���=~�� �z=�YQWv�XR2 f�.j�O�P�R�;v�DT-=���{����f[�,9o��X�GKrۣ�ܵ��h6�� �3M�RR��E�"^r5������w�B��<���%=8�q�@ɋj�"�O`���WqU���8��zB��ݠs�]F�'WPե� b���n)��W:��t!�aw@�_��g�8"8-�%�س�썇�y>CW��gho@�yޞ'�W�)�d���{^sD=��ܓ
�K���^����&p`=�U�Oת���3�ꈳ�ީ��	e�nS+��A����bf����1������8� ���|(�I����^��W֓�`�N�<r�"�ٮf?w:���a�-�\J6���F�7�ڕ@.� ��� *z�ǝ��E�\`�^�W����s����U�p��8�9	���ֺ�}�O�>PW�#WZ�	����6��=�����C\�ۣs}OjK���ħ]�0PТ1�*�dTCt�	�j�54&���3�<oP�}���&T�PKZ
���=�ןjw����^�Q�=y��d:���!�^���O��b�__qYdq��2���s���V�M_�����qrr����ߥ6�g�H%�]��ʑ��3d@A��v��U�	t�i�qf�(�[��D5ә$�[�l��K��V[j�So�N�}2����č,�/�ԓ��j�.��ju�ȹ�쒜�f����t�������w	����)a��	���˛�"����F)zwC8�0�R��0�'n^^P.y����m_��x,s�����n*��1����<JF�YJ�EPwT^�,x:��}�i:0�ă��R�WoW�;�A�����Z���(�*9���>��^����-�&C�S��&�̔]�Z��ts���A���E��X�n߬��G���t@���� ��B��~,J���R\��#��貕� �ٸ�@	�]9b��U�H6�a�_7 `�酠e�G�,Y}��������Vv;F��P��k��R�w�e}������u��'��61��Ksv�׺uh�����gg��JW5�\b]�3��"���f�9:�e`���o�Wi'�~�Bg�9��c}e��m	}�n�ۦ�1�j��	�9V����-,.�Q�ff`��&wG:�H����8��D�C7��L?p�)�*S�,yT�w��ԡГ�%����l��VvUPVӼ\t�.�>1�厹W|���'F�Nj��|��2��K(F��,��((U�@ա�p��J���ի�Cz#�ңʧ��M���d�n�n���z�M)�����2�|@��r�S�L�&[�iѩ,Q�u`i�'��x���+��֟j���z�nf+�y9Xv3��n-&p���k���������W������h�������]��Q�։zw�ԍT1gd�� �KRm����Z���l0�O�%�@��en�$T_m}Q�$q�����n�!�4	�E�7�kFE�v���#�# 6l\=�ZT�^d	O��������,w���]i�����aُk��x��(�\%�E,WnK�L:��&b���1=#	^N<u��\m��@����	�&����X'��{pȯȁ>[K��ҥ���M*}���>lv@���n�������O��
�ZW��A�=�|�5�zU�x=6��.�u�V�>�#N����%��Trx=X=\=p����Q�)��P�� �!MP�s��N�1u2�n�rx#��.�<;V�U����Y!����{�6�b���Y	��̴��R(*���6A��oZy�\tlnn���F���ai�0�Wו�ד��q���w��<�t�2?`b5��+�
����^c�>H���jqE�V�\���]��!�SO��V�[�4�)vbo��ߊ.�Cx�bI��v_h���^�_`
��,���
ԭ궜�u�[��o�x	N���goЕƲ�Q��]��nfQ/�ۻ [1wV������5�4�I�ł[��/�^�0+��kΚ�]�[2��w��*��%����u��oc;�6*FKn�<g���� O���{�6�r�6lE�2�jWG�wvՑ�T9���H\).V;x8��+�)���U�h2���ΝF��ǹ��ŪݕŲx�E\<=���z+�{�n�s�m�r}H+8%;ͬX
�L!�g��;x(n���/���76�k�U���r��OzJn��J�.����w�g��A7��-�����2�Q̀L�go��<���>�gB��r�tOV�YK� �\�*��kPF�����\/����,�ct��n䱐e�p=G�ŧ�ysJcj���hMz1rf�p��n^ՀI�U+�����pT�5ف>�9g �4�^gh۳�V��hj��k+��<�ƻr1F��]_;����XL�:���"�O�wl8���r��NR�d��ԉЫՆ6�̺:z��������R6��ȱ���ǡ�2"��#
�ͱ��A/ |����YH/_r�ؐ����J����Ӳ��t�'��j}=��%�}��3�D����m��(,��Yg2]��3�;�<�m..\�2��H$�=�T�m�۾�!ۙe�<���tu�[�n9wl�zf�B�C�sN�)�I=�5g 2������i(�-q/}[��ܽ���(�1�oHr�uS���r֑���^�;�<�(I��s֨�ױo�T=ǋM84�ڙ.�yB�V�'�w�%9�Z��9�x��{����_�*1�q���Q����n�m�39��D��ʁWC�!�g6V�X����7�Kw.��D�|��׻x)���6���h� mi� �h��\8j@��:�KA���)]¢5jD4H��,\B��R����\#b��̾�xkX�ݝ3�mp%Ho,��-hm����툷�Z56�2˼3�n�z;����?*��(ט~Tg�7+�%sn�_1-+[��=ipm�k��*��Bg22�˭h�*��=�S3U�0�Z�~�üZ;z���ɼE!;DM޵k���Ό���{���@WЂ[�c�suv�ݧͮPǸ/��Cӽf�G}A��ŷ0d�V���v��"}3h�}u�W�-Ls��:���֏�E���A2!3��΢sh7�s{p�4�W7��n�QV+`˓ח��_-�=K��=�q����܇S��-Y�gw��� �Gb��n�-�֖�%TA�tR�ځ�����c�h#Py�+wd��?���E
�&:�PZ"�(_6�n��k�)A�M��8��L��jƍЃ���X������]}D}C�T ���w8��hH2n+��sJ1$���7u�9t�"7w;��r���0�Q!;���廮Taw\�wrwr)#$b�D�+�ݎ멄�p�
7;�"�����9Ď��ewt)��"�띹tfB"c9r$`
6]��)W.�;��gK����Ns���;v`���N�.��I+��")�Ⱥr�$�[��8�i\���$n�'5u2e�»��Da��svs�E7.���Ü�]�%)�u ]�Ww �2JX�(1�$s�0 ]��J;��B"N���[��؄��v�21����b-�����n�ё�t+�����9ovvc璿v_8,�Iԥ�~/U�'����xޔ�"n�.��5��U<��2&c,�[�݊2�c\�3M仯�r���}���+h�Kn�:�p�$�|��4-;[�X�U]���	Wfp�lč�R&���N���פ�Jp�*l.q�hQu-����{�Z���3OZA�BiVn,r�բ^��ōְ%�i5�̄2�S��>|�8nE:ѷ�[h�}��v|�*��"�<�.�1�uW�t�c|�9�Y��imF�9��9��U��E���)��,1үm��Dp���|�[���|���SÕ�SiVUh�`+>qM*�7ӬLeR�!���ܱ���R�}t��s�s�U��͎;���3�X�ڶ{�S�t+�V�{f{��J�����:QJ��i~y������k�u~3��,Sm�~x~��+��M��>÷s'���R_ޮ�����t���U�������Z��s�t��5"{��з��s�'��+t��=��0��)���K�sFnj=��^��;�,+��e�C}M�L�%u����ƅ߅,/'���2)��r��Z�!g'q���kI�H2E�,�ξa�0�
��:��V�.�M�7�n.�;�����amŠ�.�m����N�&�en�d�<�L��ڑ0\,���,4��J�]�B�����}F����x�AxZ[��h_j]�1��1c|rP\'~�|�����s�ۿ�֗}��\��_��G��SP�sq=�n\���x�י;�j�	�2��>���QoL�,c��*�Ipf����*���4���'��u��<�����qF"�Q ��o	v�j�t��fά�2��hm59M><��ʞ��ў�c5k�r,a�Lt�&�e��bԇ�ШvS��Q��|||6��-�r��{,����H�����ׯ��$����Z���&:�=�Ow��5�6[lwFW�r��:�v$�x�j�:9�l�ⱝ��9W�^V����'��������O=��ё�s��r��p�0q��k������_�ʍkyP�keMu-�3&����}�O&s��{���b1�qX\�󗇽k���w�y�X��0�*��b���R\�|��oh�q�T����0N�� _[~�U�X���� ��ގQ�,���l�n��.��X�u��VxC�Y��۵Ȼ��wECz�U[�߲��\9�DVg����qM�7�Բ
wE_�5��Ǻ����	�L��(���mtip|�3y��vK;*��������� �4N}p�f���v���2z������.��C�ji
��wrk��ђ�7W�L%_e��xFr�w���D�z���|������L��hw��Lv��?;�5�*��L��;2*�tPx�/���/�ɟ��w�]�bs���o��	D=�Qn��Z���\-�Ԭ*I����U��ekˈ�,+�����;g9��:�G�-�<�X��Je��2�x��{�so=EG��������IQz��ؔ9(��박ҫh�>5;]x�W�*y�%���do"�?�����2eu����V��[��V]\�pͪM��3�� �p:��/�K��B��x��
+[�
��G]w��|��|�K�^�����W����k�\[�wZRu�7��9���>��P�U/s�}>����4�v�����������]�B$Ň���՜�e��8��}�WR��*�.
߷�[=��5{� �ȟWȊ+KJi�X��Oa&P{uM��J��Mǻ%��Z�N�V<iΚ����h��۽�sa�z��T�7=���l�RǊ�`�&�wZ�VU���	I��(�[�����wL�U�����2����S����菣���٪=;��`�}p��nw�ʳ^)�bٕ��2N>��%h0�����f��n2y�s��F�&��{�s��������͕��)�$rR��o-#u�ZYq�>�v�)���w_؂�zwIѪY�R�v��`�j�Y�|�s��ý}�c���s�Χ�S?Z���Nڂr��gOcUJ)zv�+��]p*��(x�+�&|5G}�Q����vo��-�	gEUc�_�����)_G^��W�_�X���ƀ��W�bn�% �q�n?z]�Q���N{&�����Ҏ�.���G��7���;S�S�m1Nc$�v���K�CU��R�z�a����s�5}��a�M]VM]���P�W^����
�n�v*8�\.����W3�a�v1/'��i�<o6�9��\�E���;eC��NGW��M+�~��f��^݁b�]Z��M�ʞR�6�����$&�wAWCf	�)�0w�!�� N\~OñvFL1�uV0�|Ua=Q\�S0��@姩���m��s�{�+Y����}��n��m�њ�{\�b����F���0-czd۫V�swbjP&jOV�׌�g�e��j�G��KRe�2��w�%��Ӹ4�������0/>�k�I{��c>]�5�7�,��T[j�3s_.���*le�͇�����f��Hl�4������f�_l��ɀF����<��y���ӭ˂��i�e�k3����y����{����j����t�2w��zzf,��c�����/������k��_�O�m�~�Լ����v��.��sT�YMU�����-��^q�ǆߺ�d�!/O;�+�=��Yeaz��k���M\�V��^���0�{W�t������&�y��A��t[�FLwb���Oqw���VRV���Q}�4�������o��r�~�w!�u��(��c�Wj�r5�:����o��.^?g��3��?xzE^��"+2����u�1�t�]�n�s	؊	���ɚ��>��Dj�ߛ�2�E��w�N�S�F*w�2��ʛ�N�v<`���2-�I��u<d�.[UB7T=3���U�sU�/5���}j)������QB��:���E���.�-Ox��1VX��ф,йc�53���;�}��mh,<OG�3K$Α1�p*�V�߳C{��7�by瞆C�`G"Y�j�K$�beb�L�֜#��o!�]�_}UU�A�S�g��ߖ�ݸz���g�P13B-|_�g£�3m��qvKǖǯ����Z]��oF�:Fat}���t��58�֚K��3)����`�S�mln]ƭ��klV�����1�C]F�M8����SN7��.%��f\y����M4���7Q�d9�ۋ,s�}�V�W�a���ۃO*�u�s=�
�#z�����MC��*i��K8xz-��S�z��5��	��=�J]�|��aR�dp�:�>��>ֵن&'{���1
귯��B)�|�1@WP���{_^b��{Z�svʎ��YhA�m�S��\����rZ�}���|.Aq�>}r����XF�~s��y�ƾ��m7==PrS�k6�,���m��:����Ջ��X�na�~�[Χ;�6�����`A��r�<��3��<R��S��쾻� /=��JQ��>����V i��u������nmE���t{Pժ��=KJ	��k�2:����Z�V�8�D��§�K�<��a�`�.�n�ש��)�Xb r��g��yyHP�뾺�_":J���}U_U)�q��{�Z�Ա+�R�nqU�u�9ToK��y�_Zo.�}|�c�ve�PJ���:F���ZV�ou\f�V;~��ֲ,�/���4��Q�r�H�y�-���ש�]E�e����+�3$9�W0��X���+���Wy�t��;)�N��׺�o&�^�|,vT7��}C���R�.-W�	�ey�b�Η���\Wu�v���&��XJ,.�а��n����]W�n
�m����n���u��2���r�.YUWٶ�g\�b�no��ҹ�T��R���}p��q:�[V�lގ���AZEMU���yy�ݚ�B�=��Շ�Z�}~���OOx<���=�S ��38���
�,���F��b`�.�K*�2�&�=�
�]��u{k�>
���j4�뮶T>�9���v����so7e���&ꂍ��r7)M5�Kter1jqݹ�G+������tC&������u�"<�5��Wv��ql�ÊYoz3�,.0}r�p(:-:�*��o�h���v�n��Afu�ͤY��Cy��C��}_DGѻ=�o�5��;�eZ!�jD�а�z_e|��!��t57�S�wq|�����q��^�T�|z`�m/h�U�+�y�
~Cr=^���4k���N/q^�OM}�u�wʵ�D42a�ɽ��t&L��'��qw/L�g��S��ʞ�;2�-v3�o`�X��Q1\�诎83�.��v3�P�N!�aB��V��YP�g������R�<���攞����e�*��L�|�^Ի��l=��0%p�0qw]*��:�P�'{X��G;jU8��Rwo�⥣�n�7ՈJ���3t1���m�oNw��=K�uX�}�W�W����t��+Sq�+m1+q���v�٫�J�펳P��+�L�����(�A緞�^S��fʻ����8�2�2�w]=�������uc'�����/�=&}�O���p8I�a�Is�,[R��[���o>�!���k̸Tv���+��nu��tZ�;8�/���]6���Nr;;Ί�iuP['..�黕�˝�^-mZ��J}{6�L9��T��]�W	<���!9�������U���h�R8�Vm�}��|> ������������iX���-��F��O՚�79��P.؄��J�^j�S�S<$B�������=.��)b�9���q�����Y��
5��+.u�*̻O]��v�p�OaT[�=A�{�MW�'E�i��{�'�뗩��W=̺�����3p�A�L;5��m�{�Op��}7,���w���r��o���M�h���{�6���r[Wr�`��r����x,�۝���<��ϗ+�{dG��cNR"r���%
�b��ĩu���f6nW?�̻�}����;쨼�Qy9X��(;��X���
���mM*�qˆ��r��Ú�m��GeWQoU���\���B�X�N�W3�Z�Fwj��Lcx�v�)�B��s5��b��b*c���~6��x���~7���v�5�����*��ڞQ�!%rW��{����YkCs����o_)PpU��.�H�Nah���T��bž8��̪X�e^���K��L�ˣ��mvq[^�R�BNn�ɠx��6>m�1�S��]u��A�����j�Z��TL�J���'v$�s,d5Pl����a51@w����_������;��k�j}���⯢�9��Vjn�#�ۏ��[�?>����I�-��3��J���V��O땃��5���_;�*����}Ξ��]n
��{�"yUv�k��R&��W0��ɚ���/�1��|�����<��mU��sQ���nƅ���w�p��	F�����w��'*��1�<�.u������z2a�o�x�4�/�bm����ho����NY���s�����������f�N��-�+� F���r�N0�m[���Û.���սyYN�ˀ���[�f�u���݉����y�T*{p��̎�f3'�%ne��,+�e�}M���*;/��άc��yяi��.'a�Y��l:�6��|��I1Sq�hac�"����8�Z%��$����K*/1U�3���M��M6Un�K�8����C4i��oSS�E��x�u��Á���q��ԭ��"��˵�[*5�]ҹ��I|p{���&�.z�V�O��!ٝRv5��F4�v��o#�FX��M"����p郡��k�8�Q@�#�]�%��cH�>�0u�7�',���`X]��KV^docM���ǖ�u��Εs ��&e,�bDE�;��j���Ru#\�el��-�TI���;G}`�DNY�f�� �Fcj�׉�R�}a��A��O���9�e�1�iv�c:���:Z�c5���p�4�q͙|f�������Z�2�c#-O��mgu��6 А-ƶ���^��xg��Π/M�����t���o��6�9��TX�P;8�4���8�М���Ú.��Lu���oE��U s���]�c��N���*�*Ŏ��@�]�W�P��j2'h��$\�4xd걤G��(�魷bU��mL�w{Eˎ̠8�l�E��<Kq�vT�@f��v&�{z��t,j�'W$�os�6:J$�X���7���75�o�&���{��:������7���L|�����os	��:6���<�]uB8��
�.�d<ӷ"��Y�+/t�����:t�R���<��8�촍.i����	ʽ���<���Q� ��Qu�[�,�����w\�2_y��Q[��^��k���p9\r�4�v�⭙Z"��`�s��cY���k�H��00��i����7f�-v�5u��8����5�8!�ܚ��4��s��q돥�t=�v�Ǜ2���4�nM�VHE.6#���l֝h:�4�if��H��d�V�C��p�1i�����<�����Z�7�[���� �����Ѓ%�w�:��]�A�ڿI�N��~w֬��\K7t/m'�5�7P��*3�gQ��rB�ΠoF�H��KS��霸���-���=�r��Y L}�fm��2����3�L͖�sLa$��9�L�t�>�d�[+���z�K#�`��Pn;9��[óu$+���&�A
��1Q�=�4jP�p+t+�f�׼�TMO��Tu�zQ8��{W+��eal.KM�se����IH��}2�Ǵ�fz�9�! �藔{������0���%`42�Qh�C��������0���z��;�=�d�H���h�E�t-A|3�|5ꇩtNpz4f�D5r�äR����Yf�*���Q�ZIՁ��%�ou^��ٴ���v,��d�At�z1M�U��9%�n�:�&��v�B���[�ׄJ��{.5+8b����mt<�x��Oo �K{N�ɓ���I��7�nP'}��V*u�{�3��5�����BY�h.l��wU���"��o>N�7��3��+'�ڬv��{���Y�4�Y��(.
�{F2E�%Ү�_>P��N-垵%W/y·sx�uDQ�����"�n�j����$����W��'�PU�{$��ģ�+011.���$���&]ܖaA'wF9��;�!.��D�p�)ˌr�	6����u�Ģ�R��A��$����FI�5)�wI���2�"��%9����w�s���sP��%��뻮���۔@%s\ԅH"��4��aL��i�;����#uۭ˒w]sr)��2�1Iήn[���N�k��'w#�\�̷n��s�:e.�r&D��W(wsE�����#��p$��ƈ�.d��'vwX�ˮ�i�]ݓ,G*�be2wW:W(�\�Ȣ��wI ��.m�����\ݙ��~~�z�O��qW�6��j��sgCFDݻ��%��(��n�T�{W����ڶ=uXp��.����"�4�I,8}�g�G�GN�+8s�c8����'���p^�p�W�њ̣̯;�͞ʇ����Y����|�3,���r\K�z1'�i�Q�mӑ�G��\��μ[K�sӸ��V�5�m'}Ss�S�~��hm=[�����E�IH����s
��E��/�[��Gw�������!r���]Q�8��WM�;T7���F<3g_��v��sys��;Q�iyZ��=�9�r�[��@�Yk˴u<��7c�nkUg�˵J�c%�8�.�
�y��$�&�[
s���}obPT�٪�(��ۍ���U=g��6s���|����o�ޅ\�b:akp�Q�[sq�i�A���<��^�h���݉ۏ3\�_q���0r�`���Y��ts��Q4�ML�*"�<�ؾ�fy�z�L��T�9u���F��8��Ono��<a\]VT�}����o4<5cH�M��4,���4�u�k��6Ч�b�k��ϦH���A�Vc���3 ��O�¸ԓ�{}�wZ�R������=�]w�*[����u��fS�qdaK�L�SyۚB��r6�\���=�a��*za>���>��
��M�hW�$*�[�vI���jwo�������Kp�@������ٗ�W?o>f6�f(w]����9�O�5-�v��9��YP݉�9쭡+�?�}c���I9���i�}w���i�\u?��*�u5��n�&ǰQx�W���S�2kS�QM�ۭ�-���d�>��{Dh���xK]�X8L��J=�w$\]��.�R�w��{�Q�ϝ��US��Κ=V�L�Q<6�GL��f-Z�BP���i{��[�춶�(v�/
�]�5�C-�)����e�u��UM�Z1n�ؗ1݅�>}V��.-���4������Rʋ��.��&��-�~���3t߫�p��|7�����PEC�H]�q�(�y��U̵�\5�h�k�i
�X��Sݯ����;�Y�+��`��"k�3�0�Ն��2xJ���Ou҄�j{/FO'�����5��|����~Vqd*�(�������S�S�����G�K���=��{�5��������ہ���I!�*��]ΡO�p��rˋr�7.��&N��Bh[�մ���f���ﾩ�mC���<
��:��zWsu��{��WǕ��q�7���^4�Q��_y;�X��[��8�{�9lY\�U��)��ݐ��S˅��KF�s�
DM1{#�r��NGv����L����ْA������x �(���O��ӈS��'XG�2:��zn�_l���]5u��Gz9���}�c�t��)��!]�u9�OC]=���+���LD%c�(�m*���m<A��5U��<�=�[��h+�ל K��|�{���(М��ޘ����;�g8u����
G�h,G��4P>���Rcb�z�ף�<���ٚ��̺o��*\r��;���g�.�Y�w�5ͦk2�=����7�ve��~��Ȗ��%Z\��{���%���F|w�:3�����
yW��߱`3��u�\K��Q���7`������|�tVR�Cݥ�$l�$�}�޴��U���591w���_QC6����wތ�IZ=�^V�l#��i�h3�+�}d�r�9���B�<��r�6�Κ��Vx���Q�,Տx;J�^.췧\�S�$�o��菰ɴ�׬V@�BS�p;T/�,��=�ؼ�Qy9��ڌ�S&�l�ǋzwx��)�=�80�7�5����[>̠��>ߊŲݱG��=�t�l��io����9�Z��]��Ǉ*��9�UJ�z��3���!�G3;�˻uu.�<��7յc��m�r�xv�`[L\T+��g�z+lQ�}��k]YZ��T�bط�J��Sx�=��Z����"�cٚ��)�����3��nS��K\����WiO.1��{�D¨�jT��F��o'���u�Bl�7�X
��93�Q֭U3K�ދ*�4�����{ESwp-�ZT2�ipR��楯���C���e�m���YF��nZN5�|�)�}�L��~�l.�=�K������
������x��V�>��<���H�Cr��T}r�/ m�g���hj�\����9�Ż]C���nQܸHղ�����yc�o�Ҏ��펍n�1����n��O>0�軻�ӶT�X�;�m`�����hE�`�3����#,Eq4xEj�K�Ùϫ6�F��`s��m���ﾪ��7:�{�&N�D����	����\��/��4��wNdZVv�U�j�ĬM]醺3��a��	[���. +��e�C}N���q��JwJ�IIw
����~��
��,�e�W����zvo��L_oPRےe���T+��+bҹB�waw���`�=�E�>}J=�3�{f�{�]5�c���g<{�����wJ	Ð<�q�<�gmlWmb����#�팛��y �wAy�'��N�t���[�A��fgk�q��z�g+�{�e�]\��mʬ{����}��Pc��V����{�4����F��ky�2��Fm��,[�d���Tg�OkՕ�^og���`�Z�=_6�wg��u(�Ų����ײOz�10u�7�\�u�w�8�O}������NJ��v%p���TB�=;�����0��GzFW3�]F��8�]8_]k��2��=�ة��y�e�X�kر�;����������3sF�U��mD��d�f�v[�F��u.����1"K�mYv���;�܁:�,����=�v�w�Yɮz��:v��{`U�&��">\2�ꠙ�^�J�ԋ��o����>��*����A�ނdcupK�����Y5?^���|y�x�_�oh��|p-���U�Z��oF�c��'��m�ۯ�=j+Sغ�-⻭h{�����u�	Fv�����A-���wB��YH�<�TE�yq�����O�1��e��N7F�"�f�^-��D�Cû��iX��m4���Q�f�_t���R��ʰf���[����>��b�F3����xJ�xfXW�Ba�J�< ��b�����4���.��@L^B�b>�2�Fv+��}Al}Y��.�{�su����r�P��S�����y:���a���d���d��<�-�o�X�]�F�XW�8�j>E:
 ��6g��w���S��E����� .�=N<���Yڴ��۸]%�c���v��C���s���1�j�{+/��A��-�OH'��+��ueV>M�U��I]�?!0o I��P�*l��d�ў7�|�<i��yk}�Rӧ��7���B �YKQ������9Q%+ޙez�I[���j�[ۃ	�V:��QT�`z{,��:\����$�;Ӽ5Y���l�\6}���
]�5�
�}�����ם����w_�/��{��^�C�h�K3���0.$�l[����Tf��zr7& :�I��^��˝���(6��~�m?e�gqe�w=�������\����v�v�����]ns��λ�9X:�%�i���Vf���֫�ܯ�+u7}�>�v��*���؄�CR����F��k�;�䭟+7/�.eG�5Z�)�B���)���{�ܼ C�ћ�s����pe��W
���1���++W��h]�C݌k+��]�tsV�bk� ��U�h�J��	S*�I���
��]2���4Nz<���a��u5�7��/:q}=�wm�)/��/h8�����O�D�o�3|}�i���xAδ����󂷣U[�I�a�����X�8ۢqM�m��m��
����Ŧo���v��(��N�K��D��gW5O}(���Ni�l:(_�V�񃰎{���%wL�p��ž�މd��*�R{4�1�=+0�:2Z��k��VL�F��$�(wl�̅������Az~s>Þ,\eqm�4���ˀ���Gej8�\B~c��������VGg"=��p@��k۷���^���w�bo���^c�<�C�=���������Ox�:*��̥�������ر�j���+>�������ʃ������΃�k��3� ��b��R��ݖ3|Pٴv{@o2u^��P�|�)�e(o���8��T�����o���{����E:�rѮ�[���?^����uO!���SI���\ʇ#�b���b�Y'���Y�P��y=�J>�U�o�y�Z�zM��A�����+l�,�͏W]�z�N����kW;grz�[���=R���yk]P������Z�����wkGR���=%�\GS�N`G�>��Vq�[�U�ejo.�ۑOtq1�N�J#�W �Sj;��AV�3�kUg�Y|��R�'vl���a$�2�y�v�(u:�p+{]̜��=��$�_"����k���48G�J]L}�k��J�VD�:L�&�@�����آ0�,�%�����'��*�}n�ʎ�N7��#�w�٢��"�8��ɻ�\��G�K}�)���!�:q]��3[�Bq��G�}JXA8�<�~rf��A׏���h�*�#k�y:�r��gB��}s�ڝ��]�'`G�5�7���<ޗ�+kԮaj���㚘����J�|;v�z2~n��L��	Wád�x�-��M��}rN��_L�^����54�w�\8R���.�0�u�N����y�v�݅lE�n�w�]�a9��UAZ������'wZ���V]h����(C�b'����y5�����'�a\��.��WO"gg�;�츫{M��ӡ&�}�m����<$���0���3�,{q{Sg:v3�ri�B�=b�P��NC�F�a�g��_h�uv�ލ�5�j�Ĳ������\��&�ڂ�4��B��a�
���������]myPo,�|o���fq="�q��:]Ng���
1���N5�5������`[�Vj����<�}D�]B��b�*�xmׯL�o�t�S��n8YٜP��`�r�<�ɹ��R:���^�_�Mm�UdmX���	�z�ly�7�HtF�*��]��yvX�a�Uՠ���g�g����i���:���=�{�>;�o��ſ.�O��JOG�w���d
5�������^K��o}�/t��
?�����OԲ�ꇏ�h�t��2ύ�^g{�1��>�mxng,����^��;X�C��'�f�{bg#�]�9���B}��Ki�w
Wݽ��45���]�!�<����}�%bS��*��ʨҞ\Ci���O]h����pR��`��'z�1��vR��;�9��}��,�+�j������nq��Z�W4,�oC�sb�Њ���M��p=��h^aG"�c__�X��h{��2S��E�Q*$f'�q�ǻF�u|/�B��*ܛ��
��<��t�wr�����۽�q9����"�EK��R�f�|�КB��`��6yn����N�z�=ō��Y�}L}޵��R(�CP�@�YS�V���1�����-�Ա��c(%~	9��+��f�v�v��z����e��i�\-L��HGL=����P1'�7��`3r��9�TW�!w)Q���|�^�^!a��}�W�9sz1Q/9���u+b�*�(�*wY�:�ڊ�E5�[�r������+.�*Z��jM��U��m�ǡ�r����o�(��Y�sKͧc�f�Sf.�:��=A�����Y�CN�e�v��{OQ�hZԚt�A�yZ<�4�s���UwE�5�v/gAa�K�6��}�K���7�nf���)Np"+�'fƳ�Su	�+�P��A�h)��st�=|�6,[G�6���2�|fꗛaᮐO{�Dy���f�<�fi�v�l2��0N/���bS�nIO�5�rZ{z�����^&M�3�*��E�������+h�Ys����p�d��m���ڙk�F��DJe�Z\���Wi6��@�k\%`�+33�6v>Vv���g=��t�Y^�Ôw���ؒ7ڇ_mlW�������*�[�� դ�ܗ���{�dE�����]�yU�[&��,3#�*̇K��	�+<��ս|����'9.�O'D4������I�[��n�Vv�F������wK�t�J��Nf��%٢�q��]��K����&��|���y"յ&��1��y�cݴ9�������6U��,;�GS}emn�4,u
�u�(���&���Z����f�׺hY��J��{Y�PװV��ᅙ���^�٪"���[0����Ka{K3���v��.U�d��v"pT5 ��x=p:�v7m=�,K��b�֐�;�X9�r��+"{�GV2�2�eG��̩:�p,�}�|��r�tWY,�᝙�\�Q��71�""��k!�_RE=�
ñ��W�!�tt1PyXh�RM��p�2�مjE�Q0X��FKy�l��÷���=o'-��;�(#4l�a�x�ul��2ͦ�b\,'��Ae���f���5�@�B7�p��V���i��5\���]Y.h�gu� ��uh9�4��� gvsx	�ې�a��[Î;��P�W�WxC�r��Dَ�_m�ְ�;��r��Y U/��;+���;u���k���v�a'u���rs�㳡�z��X��_bm[�=��騔X��Y�����ƴM����+F�=��I2�P�G�����p�{�<��i����-�l��8j�'�[�� %p�|�c\��A�۬*ҵv�5v]<���D�Iw���W�]3U�f�N�p��
���,�ͷ~�*׎x��fk͚�(� ��s�,'N��G<�@�q���e
��R&����%ca��z:����b��x��=�j�� 	G^���v�z��pR����F����RJۃBoY'�Sh���K6ԇ��B��f���r�j��F]�9:�l���*9�4i1��7(̍F�.\�B$�(�`�5$�ʹ�4fl"�;��c&�3�(��DPch���0&I��6edd��M7)4PX�, ,BF�l��D£E�� *4��-l4��)�\�ѱ�6ds��@%h�l[d�f�6e�`�E�hhT���F��0crܱ��2Dk���Rcbf���&K,Hk%�����6I75�dڐ�V# "F@�i7u�EEDh7�69�P���S�M�*;o:HY�]}	�ªK�/�T��Y^{����Y��/;v�u#�u��+����E�~���_F�\�i�t���h���e����slg�*B��g��º{�Ωl���\�u_$��*#p����v����]��0�V�	���2���3�ּސ���],j�'.�,+q��� S�y���p�v�W�����F��Wn�]%��E�J#���c����_��������T�G^A�uo���֨?u�v�&�G��!t8۞ݛ����F�׊[����̿�-w�[l�2�)�fKYnA�撝�3Wc�;û����	�O���+l�철�G,�X(�xQ�⺷���o��/��[�]׵˼ڪ{��c��0%nsq�!��S������s��������4��R�f���W����>�����nE�	����L\V��[;Ϥu{�7� ����;�1��U�Ҟ=纝�������7s-Ccg���-��h�jA�/x�V捣��TR4vL��]u����L�89�ϳz����m9��w��֙���zR��5ܨrK6��x���{[@�p��YE>����r���)�{����LU��(&�j�uݧ���PK���D/��$�:������K�&'�_��c�k�TlZy��Z�6j�M>=.V��������T�������K�&�F.�l��069�f�j��$�Վ/b�%pͲ�0�U9eI�<���3fN�[||�y���۷�}��>E���f�rCS��WP�L�U˨��yj�rlɏ�>q_��������7�S���;��U�M)f+��f�u��@����y~����?)ڬl�v
��?'p����Cu�d(w�P
 ��udc�X�8��F
��*-�b�Ŏj#VLwQU�� �Kb�2��o�ͤ�w'X�/vb�f�q��;����-��i^�8���^����9A���R:���qI\�6S�	�����?��*/1�Y��⽚4��5��B�k�n�	��sN�ֆsܩ��Õ����vQ�d�[ػV�[�O��)��x�v��w�ݙN:�l�9���k�#u0�xx]�[��xG�>˨ŕ[^},���z��e:�Y���(1�Y*LI�t��\�T�-B܏͛ѱ���Q�U��JҼ�
�ׁ�D)s����z�bL�У1`�k��9���gD�+8o�Wk�!$��S2I���m��k����TF���#��[z��E�6��q]�1�B����sp��X�O~1�R�c�i���yy������Q�nԋ�al=۷)�f����ݷ9��%d��+��qʷ�o7]z�(T_f��c�T�X2��ǹ�}�g��v�MEkYyTY|�T��J`�у����K���z=�ve�ΝQ�����,.a_���oء��;=%�����K�[����7�Su�0��k.�Bډ;I�Jgl_��{3�u�s��K�>�c��z71�?7M�Wa��$@$QUq����	����Vr��p7�o�������Y�o$�J���B�p�Ze�AT�1�;�èF��+螙]�ِ��ꯊ����u������/O��L�cJ��t�C[�y1\�̰�w(tY�>���Q���Jv�8�����[�K;g"KȊ�Zt�wc���)u��kp��L��p\�t�c���{lE�4Ӭ��{p��P�Y)!B�z�VSa쵾n;���i���ފ��M	�c8��"}{Л[�Ab�c��r���g�:�.����Ϣ�&{ASY���.ۃK*-�1]�qc�.�6��֓�@��/�*����o<;l�L[	�}p�!�7Zc��_h�y����Z��7��i�cU!rE����Riu��M@��8��Վ_kyNK9�r{x��������)�>�p���S{�F���O���ߋ�'EYw�Ϻ:��-�����iw�����x�}��j�x끽��y�>�V�iײ�߂�qC�u/o�ԓ}M_�G%��Pt`D`�Z���g���O�S�[gؕ��r!r!{j�T��y�s�������grS}�ZB�'��E=��/5o�� &�V��%����2����r�볖�M}q�Uio/�m5Άw��7��:�ZD�J��.���f��s��?��V�߬�z�`N��ߛ�yA�t�|���lƟM�o�)Dn:�ׅL����q�}�����_�e���09QR�_3X�v(����6���œ�םh=��k���$E����ޮ��5e��Ch��� gI�2k��
�S�]��;{�S�P�'���j�#��	���u'n ����\{�!n>.���T��9:�Ov}��o�+�C��lnsݱ���U N�Ǻ�������/�����t����ƾ��e>�Q�2�QՇ1���s걊�E�WNk��q����:밻/'9��jU3s���CM�o8���c7�\8jb�ٮ<a�k�}<Jג���ٯ���"�mn��<�;�=N��l�����<s�Z%tw�P#�Q�2�^��r{��}���k}���1�)+X��yp({��ؓ�)d�]��w�V��;��*���ޙǎu�oPU��MC�S8���g��ܱ��&5䷯z*�|:&i�孼{Z��5:��\K�}W7K�+�-l?7��YV����|ћs_��to����-]���uz���O�>�"�8ѓ�Q·��6��Kv/>�r���to���]O+5�[��v��4Tǁ��nWP�CB��������W����5��R�Q�{V��zrd�{�^�c��{���2�'���X0���Yws+k �a�h3��P�Z�����>57<�m�̌�iU��V䫊x�ҋ���F�ó�\�1E-�z`��������N^V~�>~0:^A�w��DP�g��/w`��Rj&�r=ݛo�JR�c�Z�;r�'���GR�	:���x*&��I�}�������}����fW�c��w���KGnذ��r�F�f���nU���bz��F��εc��:�F�����-Z�{(F�#�n�F�b�2����m��R�PNϖ���5G��~�3֠���u�t�����n���H�v��!�ziYl[�P�w�:_��^U7\.���<�8m*z7z�FS��b��9՚�t+:�:�\�A�}d��v���̍ͧ����TV�N�'�9Ż�/�G�f�,������^	��&�_�ve�绹��j�ԞB���#'~�y��N��{�e���0�~�Jܚ�ݰ�b;�u�;����}{Z�z�gu����]W�	$P��3v�A��C�N'�]������8���M���y�9�ykn�X��/R�r�^㫇��;m�N!bn������d-=FP�nG��N�T6���"��C���I�t�O�,b*��3]�l�;�1���Lc�q�sD}t�}ے��*͇�\�Ll��6��iC��}56�M��#{)eyK��r-��w���P�u�7S*d�΃O*�^31�+:�mպg.���]s�w��K�}j�w`����y���e}y��v����%	}���������m�_ls��K~�j>��u����\�rq9�2;	�J��ލUv�7�o�b�]K���;տ9��?S�u�vnP�Jn��U�	��=�ϺM֑Wǩ��{U�1W�2��TR����]�h����8KzU��챉SKu\e��{\����U�u�F����Q.�N��N��.�:���Kv��-}����K3%2��K\������ז.�^��\��{V��ǩ5��71R�y}�����l#��㡎T�1���m�JJ4��G�Lzo�wm���Fk���*ۿ��[x�U2�l	SfE��6��t�)�3+=�*�O���[-�'�@��_�B�t7�N���7��^�V1阬����o@���}�ۗ�囇���=��FV�<r{=���Dj�U����]�Xxe�+�'�C���I|�Ԅ�l3��l	��!��v+}�����2����tS75�B�ڧv�>�x���h.��_m9n��3nV����y=��}�:��"����Q�67}��zC�R���TM�f��`��^�=��
�u��h�YS�0���2��Akr�2���r$j�}�{����_B��WH�CU��r����̰���l����d-p��i�}]p�&l�ǽ�	��)���ͼ�yzyA8Ukr�,x���_��T����#����Rj�S���n%7�zl�������Ɍ|z�~�'�6�T���f����Rh��]&�ms�v0��b�I���Δ�c�s��A��|'���W�~vQަ��]R���NEH쳔b��q'���6/��r;+��-�7�bzuFG�s���d�w��;��ڛ���[��dV����}�V��h�}7k�Լ�E��ވ�חX6��\錱+7����fD+���H:� #n�=�X]�W��ޮ>`��K@�f��b�,���k>��S���X:�tc��o%�J�/D��.��L��do��c*�<��'Qݻ+�9��=!��>��i�{�~�D.�>�7U�O1
�Q[�t�y�Zb��쯹&'���j!<[o�u}0%)�j(�w%}��F���ۗ��K[�ů������t��+Z��ؕ4]��WA�ge�d~䭒��M�q�~��i�Ҟ\8}�	�\�<��X����͖��9Z3#��]�	v<`�l`Ro�d�Oq]����k�Dù�Wr��L�m��|���v�R1��8�2:���t�E���=���/I4�8�p�"����DG��E�H��3@DOw�T��s�,��G���O�9�k�.����p��Qn�M$"a�k�VxUed����a�W��GG��n�b������X�f�l>
���;	iۣUtl`�ʬ�:1=�zk�\�?��MF7�a\�QU	:w2��7��ӆ����n�t�[�D����o�S�)�;扫��r�;�˸����#N�GX9,e`����1\����rM�Nk^�Ѡou·I��4���{b����ޜ�h�Av�����Xr�,#�2
v�J���)�r�l���F�w��;�����:�:�����zs\��+����d�涼��pi�}��-�X���GuQ��sLS��N��a�ju���~�f��ʤ���w�:O?��|�?�{>�O���O�Y<c2�L�h�5v���8��Z�uk��_WQo^Nbx]�ݫ��:� ZiE�oW���Uo�z*���?|�v�ѽ5�g>���ymązo�|�gQV��sY�Ȯ����&��ё	�W��Dcô��E_3+H�Ow��Tgޥ�����/�R�c�Z��x��}���������(d���ի����`�Y1��b�/���m}��z�n;{����9!vX��{IO �SL7{�R�X������/~��%�ü�-i�,���nG��ݪ(}�*i��
�y�x�m� �90Νk�r�)RfX�1�������V�=�ƶ���XK�%Pʅ�U�R���6��%��e�il�+�W�i`uZʋ,Б",��3��eok�,[�H�T\��ġӗt��o^wҙ��+�� 5�a̝�vȉC;�$�y}{�F���d>�Βn�x_o��FY�����9Vz,��bN���XE�[����n骆��֕r��r�K�L���<�:ͣY����"�Alދ4�g��!����2��f����ӜC��܆��>�q�G
�cSÍ(�Cw6���s�F�WtK�p�S��4�<1�Vw��ڼl' ���9�s��*�Z��s�T#VJ��}M�A@u$%@R[������b�@���M}4���<���I)$������Sl��ɦ�m�ʫ����U�ȹ�{�>��}>}�i� �k�-���b<`���nN���ڛ�!�)���XW�WΚ�s�3u6ml!@��1�׸��If��x+aC����-E����Ń`z4;ݺf-ɛ��@0_ijp���彸��c�B�W��n�!D-�M��-f��`�����&����˰T(?)+�* z��'��}�8�wdM0�G�=F�[+in[��PR<k#*RK���.L�_.�|���㡻L�Fk���J%P�5�;1vD�ګ0��TR�}wt�h�)��(x��Ee_.�*��.�z{��E\�S�ma-;�u��O&�408�#�L��_f7��-bz��jd55v�\��6H]F4���^vS-�sh'f�9]��Z-��ޫ�kC��<5���fLF���Nr��G�7^1(X���#/E0(���]��媃vqX�̈p��a���KP�; �^?#�_w>�%�m�{Bв�禚���뤻n��j�o\�	ꅤ�(�1_��-��	x;�ջ�%�S�.S��o�jږ{P�hj)!h��`g���2��Ӳ^��<�Z=2m�*���M����|]��=�3v�S1N۫����d�uZ�pl�%���Vf��C��r�:��(`��;�5	�[J��W�.dJ���|tm�u���,'�锧1u����0�9���N��%�ˌ 0RNͼ��z�Q	mp�&�n�{��)�k/�2pH�]��Y��_\DM9�Y::�l���B�@��Y��R��1|�5:��8r��3������:�#W9���<k.�G��ougi����(s��"mڲ�#�ם�X.R!j(f,-q�D.�-��r�h}38_k�;x(��t�Zso%�+J�(�1^�mt9e"�urcCRn��[�]���������R�DF�H\�9�t&�gMPD� �:��tT��z]��J[z�+��	em�X�|o�d�;3r�4�j�5)�sV�ޢiV	(�C�]E@�w��|�[�6=�;�G�E ����5�w�}ueP�ԅg]��sp�B
V.�J�h����w��"A�ݎ����'gf�:��U$�K5U��N"�0FC�uЈhn�B��q�B��^,S �4i��̘���b��-���ۣ&��;�lE���wt�QF�TX��V��6(�c��,�@�؊9��0k�D�CF �QF�h�b$��h�lPR��.�mDm�5���*(جF�,XŌcI��X��Bl[�t��h�&�+F5�d�4i#F�ƈ�X�&�,���4cE&����MQ�UЪ,F0ZB,ZM�h�7H�b(�T��r4F�_P }@}Y���c9�[�����m�.lv���*����yB�DwU�WU������
�U��A�v���mX�í���l���f��~�wmyۓ>�B�r`K<f�/�9�<�9q/m���O�w�P�ɿ{�^�Zڢ���'�ы�݉�R�bu5����J�L��'/9�����Y���_D���׊v��[��,��_;$=Bq�w�����@�[o�&�2�&�ݿ���e�}L����mj�o��u����hS3�X/ϳ�so�ڊ�����+�+y5]��1F�B�E�F������m�=ղ�K��4��E�;\i��`��u2���v�Um+������s���O�JǼ��}�݉��q��,_;s��<r�G�N{y��9�z�8�����(�C���qR}�;Y��N��V=n����uU��}�1�l�������j�{K������){F���s��v��B3^�*�Gi�ݥԻX�ֺ���X��3Qxj�Q_eN���_Z�������.aBmؽ��Í���3@�7���v�^���%u��`�۩[�Gq�݀6�����[����%�Y�MU��ɣ����ܮ�.�w]\dHV���6!��QQPofTZ��\{U8bK�8�����y��,�T�]�tߩrl���o��+Z���T7�=[�:M����������8����7<�\��s�>��pR��)�E����� �sS<�`��ߤ�=ϔ��)嶟v|��]�j��ī��������ˁ�4R=����;�gm�Ѫ��ꦎ�hz�q���G���-q.�_f*d����~����[g��F�@�S.�m0�/գ�{Θ~BW�I���_�<65m���U��_�<�;O�y�r��b�B+԰�Ĵ}�0҈ܾ�����Y�W�/M��\���7AM��w�wA�=���Ϝ��<yO{7��A}^ÐKGw��]���6r��9}v�5^�>��+�~�h߮��2���Cŋ0|2��&"����_��S�r��z������#}�W��������q�����W��y���ȇ] 6tԱ���<|ϼw�"6��w��=��^|d{��L�|Q��ÿ���~r=ҡ��_��^y^�����6 ��r�#���"�N�Ύ��-�u�Z��]n櫇'p苗`�M il|�A�@݊�4e6+o9�+
&(��=��R���u_1{]��J��wS���U�i���
%q����sD����{���]D�
C��G�GR�ג�I���3QLz�J�K�Y�F{ޡ=,}�Qv���#���zb��i4盿&?{s�"��mz��������g��`	�~�j�|E���=��_s>�oI��w��o`�pO+ۣ�5�k�_�׊{�=�L57�bV[�+di���^q>�W	�{�F�k���w��]U�t���@��?;�V���N�y[p��T���kI�<5ɲ��3�}�v�9���p�^�Q=��|.�#��rp�LmFMip���u57�u~���X�Ʌ�7>�4b���e?q���>�q�j�:0��u�v:A�U��ͷX�3�#�}�lrY8��&R>�B��>g�=�^G�s�*]������q�S���58c�A��y�Z>����3@dT� W��L�L��ά0��O�ð�N�~�-g�<�z{�Wvos&�
Ϣ=P�:���{'	@>3"��-��mCF���I����	�Z3mo�vk�݇�ߡz��P���2�^D��ߦX��22�[��}��#���g���2�tɬ���"�3��`��t�``" �[[bq���̛DV�%�pn�Ω
CMᝤYN�� ;ёQ`4�u��oe<ty�:J��X�]P�'w��>�T����ѷrf��S��\�f
q*n��L�����&�'`^�a޾�m��B��o�9�����pw��и���%��f
gn*dIs�>�4� ���nɋ��=ܦ����f��=������Q��<]���"��9 y��+����;��#��U���<���w�O����R��/~��C�����c��zg�� �}�%[����7�Ϟ��q/b�ӊ����i���g��נ�?g�S���,?��>�U:�mE&�^��Y�ɞ+@�����ez�B^5��Uyț���en�w���Q^�U�xh��b��j�|{2�#ʠ�y�P;�Y�ř�L�K���}
v�N	G6#�^�͏0S{^?'����,�~���`�����ɣ�2���Ǿ�T|F��C�V�d�?P��/�?c�Z4�k�X���Z����w%{5-ln���x	Yk!�s]�y�ңݻqW�m�7���~�(m���:
����LO��s�����}Ӣ��ڤj���څ���m{�<�{��o����m����]�aFד��NÇ�}	����~)�vZC�t�O�]�}R=���
�}�ދ�p��:�7�ej��ցxjE�U�BH�¹G���6}�2X>dd��i���l�K&=�g0NK�+���PMū�6���X��	kt:�T7�(y_m*ɗ�B�`Y�I-p�:��s��ɦwC{�cFb��Y�{����jKΔ�i��n\f6�U��ι�#��݆v�A_���y��N�*f=�~�t���L�'�C����9�N�ʛS�c}�Ѥ^���խC�u�z�_�*���N��Xިj0�f�e����F�2�:�+���wxZ���G����~j��S�Y�z@����Ȱ%���s���q��Y�ٳ��޴{�Y��G�uD���G>dx�7�{��s��z�Uҫe�f�=@7�UHͶt?(��M�1�q�ޞ��]~�=�ø�>
�p7	��1�AW3�o�i�����9^��lĶ}���������������5誑�3�^.W�fς�����<nQr�G����čbc�[^?��Y�E���^��F�0X{uH��}^ӄ�wr��=����U���k��y�bH�qR õC�34�n�3>@o�or�T����QMș��r�F����KƼ3�
گC�5���*�U/^)J��߽5�q�@L{ٓt�O���͆:�6�u��5����Dc��D���7�L��=^�>�}f��:4z��rUh�C;@My׉y�5����m�fֆ|�>Q�3oƇ	)XQ�u���)F���a)�n�8ˡ}�*nqɊ��^�;�Q��8�1YhVu\��|lܘ�,����,�$Gd&��*�6�F�w�H6ܤ	��]�k���V,�ڬ>��V�w�m�GW�l���n��܄x��YP.8��I,��g�PFgp���]ǭ�������G�����z=��z?e�ȟ��ǣ]~ȘU�2�����o�m���Ӹ{ѓ�����5���^��֫��3�L��hN�mΘx%�ľ���%�ܫ���?(��=�n�v�fK��6kM�7��Svղ�ux�7աͨA�;��i����y�	���T��pH]>ݯ!���x��l �܁������ �\쉷�Ұ��MR���z�&�� ���8dw��rK;�Y��φ?���KK?)g��U�/�۸7�C��gE�9�;��v��j��v���^m��.�ϟPÛ�V�z��uW&�kVW�Nl�*sw1�s=�9�h;�.��=�~)�O��v�7"9��Vo��f�Ӡ���������-w��O�E\�>�(~�>@�h�ȇ�Ը�C��q�����=E��9@µ)�Ӌ�B?}1�܊�w-mVbdEx�[L*�����y���{!���B��'zv
�o����tV�N�(�!W�B�2<��	�fHC%z�%��ن�]w/�~�����f�N�So*.Ȳ�.��w�@�XR��!�qfa��n��ր��j[�t?*տu��nX-8�^���Ca	�,#Z�=����hN�{����b�{�5L�6���)2:4��F��/c���]�H�Q��gA����z5�����V����m���{�W~"��?�]���p�#L�9��=�FF��9�wpL?'Fq�uqs��{���R����>���V�z y�6�S�/�:,\>P�4������0�����eqY�ɳQ���S6�|Ϥ你��`S˯Q*�h�}7Lmqo�����Tۼ=�Y������/i�>}c����^S��d�{ޠzm�=_3tG�W��71�W�#�)��3мV�x߾�����>��V��f�i�RUrX�����ߝҼdg���}0b��I{}��OrY[hV2�j�Ɓ����"ɵ����O@j~�c6�0�+��dCN�A��g��}wG�o�{ʟ��O2������A{0pF�mr�a,ڭ7X�(\ G�fJ%���=U�����N�}��̌�L7�ݺ����x�H�*vXˌ��W��rT��-�]��Z^�s����*�7R�:-���ϟ���\�΅�G!��n#�t2����P/!f�ط�VZ���{fW�/�R��2=������{���{��k����(�8Kg��Lـ	����\p�Ë�O���&�z��ڼ�W�]�v}t0"0�/ޑ%���y�:c���#�o���YY��ox{	y���_��-�
7����s�w�a�Ǌ�W���4̳*4r�߳�����P��
��;���sXs��z��k�m~�{�7`(����:��Z��GO���)�;苟x�ޯb��ޟz��o�j7��>��<s�F�9�1~��ݢE�羪�(� W�f�c�ﺞ.:_�FD{���H��o��N���[�J���K��c=:�d{�^��`=��M�jW���h���P�H�>&�Fz/�������߻ևO�áUe�^�Nk�,zr���n�8Z>���95�p�
뻝���'��G���|�%g7�:+�n�z|KZd������L��ǒ!�@�cs��W"��ô�l�j���/��9��Qϛ�J>��u��s.H��G��%7���l�� {ܻ��&�T����/�FA��;����hx�Uzazr��}' /{*�=g��$���tZ��* zz'Q웨��W����h�>�%��J�K�5�q�T=����@�����j�䌴�u ysٛ@��>G�L>��0�#=]&�����|0lr�L�K�Wlc�b�u|�/M�D>����ȇ;@R�IGo�^�͏i��v��f׸�|L�������r��N��FD\�W#�;KK8���V�b��Ь�������lÇ v���M�_�b���ך���̥����rB�+	�>��e�d�2��طS���8p��0dX7�h����l�f��^��F�U�2�q�:����rcA!e�c
�)�Q;ű�~����+�޻�G�C�S�EX��IG/�D-'K~�FQ���i�1+}��'��uh�<Z�F�L��|��yȄ���ۙQN=��������H�{��]�B����;�)�]�K��5��M�`mBא*�{}<��_#��UY���K�i3��5:;�Wr]�=��8u��T�VMib�&w��\���G����*��m��wL����	��y�{qSY.Vn0W�_��(Ž�M��Tc�w�WL^L�7�L�'�C���4����W��Ϥo	��=��o=zZ�CO;�4z=�H'�%����nr"j0	�����o�ax��Ly��S�3��I�^��+'�>�J�N"�_W��GJ�~
v�=��N�����p	�n�ª�b��gu򗛲�����}P�|�O�q��K�s���g�v�/>� 6|\��E�3s�n��U\dfm����}�@��x���F�_������QP��1^�p�.\�����9�*D綆���[�>����d��+�aϋ�㙳�>����u�(d?m"�=�G=��g����R3�1T���R�K�(��i�Lu����p���3�D@�!rƍ�}��3����a4e!y�B�ׄ!)�+�c���p!�f�&���y�Y=p3B���i�*���1���5�i�W�>�tr�B���I��:<	��:U��Y1S��YY����Lf�Tu��O�8<ڤLM>�i�Z;��<�q�r��L�f�D�[ Vꗾ��u��/0Tt��\1N�n���d���bb)�n�ǿ	�y	Fr��u�P�kWi[��G�=�*�r=.��Ϝր���<�] T�-��co��!���N�Mhl��qw��zp�k��p���\/Vٸ^~�
9�Wdm ��K���9s�t�+�7g�^�r�ݽ�Ǖ}�C}�u!5��fj4�y+����T�b�7�(�~���y&���$���y~�Eq�k���|
\����*����/�ú���m0'�g�<5�^�������^
�n;H��x��ό^P��)��f�&��i"��D�G��Ō�8w\����`Jʶ@��^��Ɵ�6�'&��\��s��[|$_ژ�g�����A�ݯ!���x�����c�v��ޮ/`��#3�s������Us����������,�Ǫ�ҧ"����3���/�t�P��|�o���LG�t���aQ��b�q�o�]�򠊸}@S����U`(����b��Ⱦ��c�N�[qT��2�\��x=������WG��Q�<:�Ax�7�����.����St���K�j�jY��v�ҵ������s<8-��ٕ�h(��S9Y���郕�3C��?%vv�)u���$ܗ)���X޶��V7������\f�Ҳ����i���3^bRU�خ�e�;����d*h��-;Ii��y�\i�U�g��k#��cN�i�F~gȲ�]J2�S۰�+��]�6`�{��X7G��--yuu�5Xˁ�3fq�����K�w��]C����C}��Ԗ*�v:��Sk�&d6pBۺ�����kfԮȩ���%$:���)��uAθ�fsPe�	�K{S.�E��C�h����;��Mx1�ے��7GlU�c�/�V&��p���!C���ݵ�WKZ�0Ջ�\k!��k(�ְ-�x��yF�W[�$5��T�gѕ�δq���u���Nf��}Q�4���٠35"-�<�p���
�+��$](�$*P��F����&���O}�9�&��,�r<�Ea���>wtv_(���ʠN=�k7��Wάo�x�����L����H�{S�ƭQ8_Z,2 Ī�zl7��b��@�
M��^�ե�}�"��.oT�6���jQ�p����0�A�s��v��H+bOZ�9o:tĔ�0�o��AP�E%�	+dz�Kf�SJ[z1�g��-9m�-p�_;M���&�ƍ�t	*B�h��sk�c5�Nt&��먪!� s�x�l�����(L�=t�E���,<�u�y�6��k݇x��Ɵ>E�?dM!e�w@��z�s}K�4Ly ;� ��Nbx���h/�X�Iגb��
�S����@GGV����\+H�����'L��LE�^
��U�5�'/�L�<�"=^�o(��v�y͈9rг����<���*<w��m�.�N��QLj�j4v��c����s(�ާb݇�:��}����SB8���0Ղ��AX�a%j�\MeE�KHX�N�	q��V�H��
�22��Ji�s3<&�~�H�n�{u�x�;��m,kY����}Ú�d�γ�|�Y�b���&��V��k��7��Ŭ��yAG��d!M�wT�կ;�W���^0�*�A]�H[�����<�3���OuΞ�g��;��h}1���,.���ą���ロ�8[�,4;9�I��l�N� ��ٙ���zV.ɽ�#��d���ۅ��eb�Y�r]^ӱ��wa�&���-��&��h�ڙ�l��r�=�{{�Ɯ�:����IcE�/�d�ݻ�'��;��K��
[J:(9A�hv펱�mܼ͗�6
,��Ⴆ˃P3��`��fVf�X��J���@cy��l�f���?nMђ�U�=A�:�t N>ۄ�=�of�N��aׯ����qa�L�>�zEC]���v��θ�
��
�*�B�Q�QF�)i�"2cs\B- RQ�E.Z5�fj-�n�"w\LV#E�E#m���U�1�QAjH�wr6�c��4Q����-&,cF) �b���H(�X�PA��m�X�K��QF1����DR[cZ661�"a���wuEc�Qb�4j6�#r��ƍb-BQE�؊e��d���6�,mE���!Z"��ɱDh�Uch�Q�6��&�h5b�F�ۆ�%#bM�$[���,Q��Ch�)W�P 4��a�5�<�x�R��4����K�ׅ5�r`@m�u^��5�v�DW[�Nvj�v{lt�|8�+Ph���c��7u�N�j<��*��s����|]{N{��R;��qڨ���,���Z'�O#���	��coյ���b��,�X�Cڧ����ѐ�z�~�q���=˓b2{=��h6�R���	T��Gޗ@>ʩQ2��J�u��P����>~t�����{0�2��>�Ż�9��^��cV��=��D�̐�J�,8KGّ�U�qc�x�w3w��PC���p���5��~�Ё¯��Eǽ^7Ar�=��SB���%��7�o�dC>����������}�ڏ\u%���s�����F{l�V�+·��T%Dv '�SFEd�v8ԥ�=�����a�^5��y]��u�I�{@/z��yu� ����l(�����x:��O�|��ʈ�ZdV�kð2����p�x���:R��0�	̅�#�^;���c��99G�R�웨��m������k��:�m1��*�,\5G��A٪��t���]z�ֺ����E��zC�@{d^@J�����u�n�w��=���F� Oܯ��{������U~^�urN�*re�Ý��4B����)�M�Y|��i)�6������7���'c*�xS�G�^�8E���3=���+a�nK*;�ء.�����E��掽��v�^+��_j�8*ڽ#*F�a9���9gq�F�i)����]q=�uBGz��OՂ~�ۣ�8���_�׏��i�x��f�r�^���U�3<�� yfz���d_���<oݻt-�Eh��<w��Df���2��ۅW�q�"�g��Z��6���w>��<��v,u�=O�ǽ�Q9���oh�����Tu�����qZ�ӽ7�P�t����1j���#ٿs�g��*~+���i����(�g7,^C�Pww��9'�mmh+*�	�.y�'Y�ɟ"�B�|χ{μ�o���-=�����:G����/Eߚ��+�
�n\�.r*�	��@��Jg	ayu<,\uS�h��sv ����>�%({����U ũ��C�\�9���j2�t��](چ�Q���:�b��5=N�gi���O�vo�����;E��6Ksq��r���n�7[���pƏg�z��Y^8{=�F�8�z���6_���w�����ѐ�\�_�d��-���)�b�]&��9����p��������F������㞙�%~��Ҫ�\!�<ߑ�^���B�I���ŗ�t�����g�}q�GN�a�d�S���ڃ����g8>|�x����A��Id�p��xҿu�?d��ʍ5�Ӈ����5�B�,�Y�{�P����^�]zU� ���t��I}�E�8�̍\�J	Ύ�x�&�Y���m�S&~�O3��i���%�c�>�s1~�^������w�C'n�\�81��2@���[���1?SU�n5χt/a*�,7����Ԡ���[���9���l�8�9p'�S����;j:�Ky��*���^a��k�4	��z��̚��p�a��=�w,����H~<��`_Τ����fǴ�n�;�ͯq~Y��e�P��;�n�>�Q�y]�UO��JOC�V�`{F��w�J9q���vX���92�v=���yvҫK�wd�i�f������dBs]�u*����n*�ʎO�$�w�Y�;�6=�n:�Տ��%V���kJ���+M�o���6�Z�E���x��*;�ґ���ʕ��yX�9-~�Q�J��֬�}꓇VU1�gKNx� cGMP���L0�W��;�3�������z��ޥ�Û��a�	l��ꗤ����WLa:�}�>	��R�~��I�����/��L�;�Zm?:�=�������h���
sp�p7&b���C�y���B�@Z��;�t*��z+�L�ṫ�}��u1d�C���1��	.��ޗ�۞�^^!G��:i�øϢ"je�O�>�S�qu1�owqEf�����[.�|�Y���r�v�(�ˊ���%1�f)�G��FN9��2���B#bveE�ic����/ }ڢ?��G�{*�~�W�uz�<�V��*��o�@SFPf� �vMy�fG���C�뫞K7�=��+#f����uC���#�>���r7���O����Ie�2g�&����]�9��u��=��}�3=U#*}H
��h�#e�Q}Z�~��g�����t�����&ÁF�'�k�;�j�{d��1>f���RD��Xr��>
�����u�(g��H��[>.�*Bnf�!aL�t�ϖ�֠���w�"EE��Y��o��T�����8K[;���S�|�>���Z��	ءN��|VR����;\ȏ{؀�n\`�u�p.U��&@zj�&)���K��g<n���������qV}��1~��>�=�� }�m�5=rD��[�f�q�D?{{4��Q�^��=�������W����w��>~�G���rUh�C;@Ty�z\�}u^���g��y_����������_��h��2u��^�&���X�v�uG��:��Uh�|ѳ�J�P
��dZ$�C��n�y�~(����=�������N��q��3Q���W�j���/WO2d��u�����(���Y�#��:�|�]���M}0��,
3��Rrb�T�D��m�f�Q�5՜��eI�d8��Cf0��i8f�{��EC�Lڎ��P(�i3�V��m�;L�_'�Øik���9�ne���ǳ:K0lA�ͱ����o?}#8��U�`�ppgב������Y�@�wSղ����؛���t{��W�Gz���Lh���kE����9꓇VUC�_emC��u��r��!v��;��qwTJ���l����*:��z�w{+���{�!=�,��paS�Qck�Wp��Ν�~T�BQq��Z�Q^�Y��}�;��L���?_���w�?�/�����~������pU``�s�^�E�͟g�w�ҧ {�\u�L�1����d-
}�2��>�O��J�69��VMg��6����/���g>�L�6���ʬ�22�ȱy2��7��M�SGC��D?uy�9�Elߍ#�n��F�\MzݳK�_zU ���L�@�R�]f�
��Z<�錟�p��bT�m��ݚkn��o�tF�w��;�p�4�nl���d�R�G־چ���4�n��}b\2���^\P�F׺ߎ�e ^z��~�d��,�z��� o&Q����.:�	�Wu�s�6�w<��G��c���P��}~��NW����3�dW�꜑~t<X��-R0�����UѴ'w�{�[5x7�ς��-AS�*h!5�f�V��m�<��r��j��1��u��,:���X5#~
�`�l��﷡�"+傷n6��7r��@���I\�T�YIs�qt����~T�O"��Q,Y�{i����t�6�Ǝ>��'�m«�$?��r�����Tzz��I��ו1�f]Q$�YiOkf��@�Q~� �עn�,�#����"�\�`/BVj��x�ſ:S�:����9�T�2/UnE�����(��ﮥ��7P�'p����5�k�oi�r�%���>���>�*��No���|O���~�A�J��>Gz'�=�[��m{��zx�`<G�{�t��zfp�V��y�rw�s��G��'�ު<�Jމ<s�%؝�xn#=�6gX�~��>�s����Ò1g9�^��:���ŀbs�"�}Ln#ݻt/��Z/��r�ٜ��e��Ǟ(��3��N���K}�ݯY�,sq��6��v|����k��F׵\N�*x������g�w�9Z�M�~T���ޱ�,g�2kK���1z�'7g�n9�����|{���~n�Q��UL�<.���s��<��}���VU`=�����3�^t�U�|φG��#ٹ�}��v�:�Y�^��z��Y����sϬ�|&Y_K�e�EU�5<�~�����xX�Q�3o8bW��9Cs�bP��4�=Rl�fؗ�p�v�4V�,3#N
�w�Q�p�ν�.�^
	o*MV�Q���.�W�g{����X��ӕ2�֬�����&��젾�tidrki��k_t٦}ʱ�ۡ�q�mZإ���tgg(��ǣ�K�����yH1jx;���>��2�|f.E7@Z+��6�*�= X��~�7���F��s뇐�^�Ỏ������^Gʨ2�L��Ġ=��Q��1zׂ(A�;k�_�׸GO2�6���_uC����9�Q�s}����E��^��2r�:蘑#~�*yj�Rk�S"`�W�ρai��~5��y-_�ߊ�Q~'�]�pEz���zdz7_2�.��l�=	��7�ۊVD�9����;��^�=��W�����ㅵ7v}��V�y�}	�AXe� �/�����^&&)��7��z��^Qb�^��l�FL��c�qz������e�
�z�4�UU�x��˜��=]&�K�긫J{5�_=��|��\�}���U>>�=��P�����Q��W���͏i�ݨfV*Yy힘ʏ_v׵��G̴L���ߓ̿�7w>##�0�Ͻ�mQ�_w�J9q����؝����WWw�nW�g��Có��[=&�ez���s]�G)��n�Uǽ�t��SF}>�rr��g�tC1!$))���<�j�u��;o�td�<�[3��̉�:��	˲��7+D�]�l�$���)�NQ����h;�����{*ȎVr�tY3��r�?�CY�p-R�wk��x��d��g|��$5'�o���Ϋ������k�
.	v��w�RIg"f�����µ�������7�o���3as�}~�|���=q��<�Ұ_�i]�]��脶���x៚6{���-�i��ig�+<��J����`T��lu�/r�u/d�
���/e!���`���T�
�=���t���dςz7�Uw�ɡ�*7��>Їz;����n��l\�z�������	C��
R�M���j8	��\3�����0��V����G��~��H�ْ��T�w�^ӑ��z�8)x���;E����
w�9����͝y^����5u@�\�r��h��uC���E�3��������/��p���/eoM�;]���=
g={�:���7��T���U�*�#��a_N���#�N���H���2f�bߡ��rɸ�?U�ڟ��>�K�4puϛCZ[������x�s\��B<;O8�E��+}{���#��߽D/f���nY�_�3�,=���11O��s�%���r�p�'�p,V��H$�ˍ�G������R�z����6-׍��T�ȉ���	��}[DF
k-d�5S��$x"�Do^�n[�e'�P�I�؊o��ts��y|+ʎ���鵻�&�'2}�߮R^o�s掺���9`P��tۋ�z�i�nV�ر�.eu熶���S��k��Ym^CƘ%��}//V�"�T�� s5�;_���0��6����K�=���h_��`W��7@Z��f�$�X�Q��B&4��s����C5/����5V�G���Fa���͛��@y38=�����W��]l�_:����.n��
Ϧ��n3kG_�:��F�ft?�����L{�$��=5z0�7�ۃ�&���q$��8}ߤ�����x���2�a���Zu���KG+�G�5]��K<#�����Z�'��#����?Ng�=W���ppg6���W��y�Zo\�����q�L������,׬����9Dr�[�V��O���5�״�qϽRp�Ȫ�����秨�u
��_�u��%>KgnO���m��U���x�{�Ú��2;�i�%���V�*d1��s�z�#+ws�f�+<�)[�����3q�,m�?_��_��\w�=y�}�Ȭ}@S�=�䷦"��d�>�Y>�`�UX��xJs3���N�M�;��~/�D{'�o�V�4�����X�>��oo���N�䨊Eː�VG�s�X���C����q���|=]��y�g��[�n�L��4��LU�� 2�*g-�[���%��.�]���t���D���q���m�e����@�Vx�#Ԇ������̳5�YO[ެ�&�{Q�6�:w��x7�ЉJљ�K�U�	��.�|�v�)M��$9Ό�ICP��vT��>>��p��,�dF��f�.�}�R0��jW��F�
�=|<-�_7W��+�2��:u�����m.=��2a����Dt�7�Cr�����VT��^�����^{ҍW���l�����G>����Y*/��@������9���Қr��n}3B�l��K�����s=�L��[���y� ^@�h�yQN��R<|2�ssJ}�Nڼ3���B����i�g0��xj#��G�=�w�zgY���^�
�������Eڳ�E�AN�7�TG��G�&��s�G��2���,b�5�����??X*z���J���T��������U z7e�to��+&��en�y>'Y�gci�RUrX}���h�}Y�ʞ8w�(ۻl�5�[�Ͼ^��yD�@J�q�#�=Q���0��ͯq�w���؊� P�
ƣ�+�K���!��S�.#g���U	�J�?EOș�v���xn3�P���qI�ZoK7��g��P�;;(�J��ܽ]�3�L7�ݺ�	��{G�dz���1���QQ0��Y��&3scx�����v_rl�?#�qB͕���w�+�=�]�@�bOL�j'g�޶R�6̹&ܺ�HB������Q�ל%]4U�r-�l�d]��&��k�S3L��o��ew�Kv�p1v]��t%�F��M�e0mv��Y������[R��=�� �ٲ��oAƢ��Qn��h��F�,g��6�klA�
�[(t�y�g��w���
]�L(c����
��7EE>{V�l�������< a�a�K���4��z��1Q�`oql��FD�M�/��y��+A��������l��'R��퓻j�C��zröY�X��fP��������{����fՉ�����"c ��)���M�^ʔ\�kG��pL�W����L���Nڼ\VA�l��4C�TE���bHә_t��9|�P'R�c����$:9��x�6�ܼV�f�Z�	�lPi��ʈgfҴm��l�\���s�W^>yYD��� 0m��a���ƶ�H�ԺD ����,��ykKP�1��׽���84x+��\�����Я��:%L�s�\%��xݬ��X:�^��4�k�9�������8j�\n�u.�cu9���\��t���wN_�K����p�ACo-}���j���6�Gсx�p_s��l(<դt,Z�n..��)%��5+�R�Q57�^�C�;t˫��!�%�~�4�!�Wj6�
�ٙ��wK�b�pd:�#R�:Ӟ��藍�F�+�j�y7�6/zUR䤆S-�4���� fʧsJ9�U>��E��I{T5;�G�R}/�EF>� H��A��\�Ƣ�d�+�.��]GR�5!C�ݮ�v+���q�z��g�y�`+�6��pbJ#XK�}�l<D��C��"�f����C���G�c��=O���A��r�]��Ь�W��j &�kVf{��r���L�+v*�fG��о{U
�ZB51�5��ͦ9����=G|��w-gz�,�X,ӭ�娙�M���$�](��ϕ����:��VCȭu��;���Y*��1�-'h�CS�tVI�\ڶ6�\�ݾ���|i4�ZnBq&P�z�(�h굜{ ��#[u{
����&!7�FC�� uّ"I����;C�:�7|�T�i�5#�� >����{���fnA�`��^&���/r��*�lu��Ε����(�uڡ�T#aI��vb9�p�;��oK��x�9�u�M)C�n�Tۣ']S��Lةш��%��s��1˦����w._n��0���¦@��]�ޥ_��4��n�9-�m�O�|��%�.����6��	��4"����5�_F���W�P��l�ыF�^�-��`��ca6��X�ʹ��4Q��4TS+&��U I�(���F�h�ۥ�ԑEi2lF�Qbت5lY
)6����C�آ��6+!��6�1E�F�Hk���Db�F�1i�4h�[�,&�$�QTb��c�nJFƊf��E4�b*�b�W"�U��5b����Q�`�1"��EF-F�R`��֌X�4�2�eP$wt\ܣ �=~�Ɍ�i��ta�R6&+cnb�:r;��@�AԷ�J��F��I�l���P��I��T�S�S�s�u١��M%�V����J��_�w�J��}��������>�����ծ��W�Q�Zj�W{nQ~W�ϗD�~b�v��fs��2��N��SQ�Z]���cY	��#�q���o�OǸ�O�t���Uy	�׶~-Hgݪ�^��7�Q����q�ւ�� ��,Y8�dϑy�!Ti�3�3��{�>۪���7}��Oo�����m��g�눌��r$�.n���ȁ^)��,/F�zv׮O������=
y^���N����Pa�[�\��e��&� M7@s똳ހ����Q��f�X|���6�xmZ}q7�t���|{�������Qe�CsQ��3#B�X��cW��<5���藖�����{�����ĿZG!�J<�o�tTE��ȿz��Z��d�d���cM-#�վ��i۩�0T����XZs6_��L>�k=�|J7�'ž(د�t+}����3����(>g�����?S��ѐ}+N��Tr���R�L		��05Ue]�����O�^[3�T�
��5�ɯQ �-��n�����b�����|;� K62m��3�^�����]-��M��0��������ŗ�ڴ,o8�k&Z�HjW'7��*.#m\�wgx�p*Y�X��"�阸lܮeh�>��
�|,�E�u ta�S*Ԙ�pp�j��RP�,��!����)����d��]�V��{�f֣5�/D�GY@�M�{����R�����_��<{'��:�<z�;�EUyɺ��;�g���y�C~bg�e�IvǦ��N���b�j�|n=�@y32/Ŝ�/D�v�U� ͏i�#ik7/�_�9�����F�.7�q3[P�i<��Ϛ��{�@��w�ц��w�J9q��=QW�G�=^�<�R�g���\Fuhxvrv4�.�b�Ǳ��/�����fTT/^��l8��ގ���g���}���Ӵ�_�5�^O�i�r7�|X���^�OT������j��j�����2�=����r
>�*��}��$b��Z�}${�y��IѾ��E/]�˺�m΅O�|yu�b���z�t��Q�8�X߲gY{��xǍ�{^��n�$�vW�;�*����ߴ���^G��exu˻Cl��}"\�����`{��[��ܕ�۩Q�f�oj����v�G |�茙Ax�<�wƝ���'�:��^�Ô�V{�>��O��Ӟ�75�}��K��d�(�^W�Zr����T;��#��O�q��D��~�:��f��"è�ֻ�����Q5a-��v��M]�׵�yo�i)m��w�J��{챼���X�I�uB�v񟶞�:�wvQӢ
Nw�Y5u�[I��U������*�G�9��B[,�h�A���o��L��2�s�м��)���p�Im����ήQ�5v�Ӽ���=�F@�7�@>�"�%��G�6XU�|?Sf/�ǯ����5�kݞ���ʩ�[��]Ǐ��v�q��LKF���RD��Xr��>
���ȭ��z�~��ZT)̖y�z/�OB�\���{s"E�f�xA�"���}�b	h��O���{&�OP79)-		�`w�z�B�j�M���*ǽzϽw_������dƯ�bj�WId�D��۩��f.�J���	�a�^��)��t�3���`S������]^��/}P=��n~�͍R����$o�Vɨ������鯒�P�7���Ͻ�P���c�϶��w��?*݌�>ךԛ�\�	����6�kC�����4��F�=Ifd6�g�|���;*�V�tf�����lo�h���YxT�x�D�~y;��:+Mƹ��29_�<*s{ܘ��{^>[]U�t�����WTp�}��k���q��ڇ���,^l֛� o���}Ӯ���VZE�-�2��.�Gz�v�+�GF�Mh��5�r=Rp�Ȋ�xk쭨{��Lk��T��끋!Y�M̏V5k`,�fbyWעRQsR1Y%He��cktὂ��j�"��o6��.G�b<����Ǆ�v�tW�%� 5,p�3Z�K뤶�Z8��iswZ��t�X+�>Aힸ��=]������"��/����2����nG:U��^�p�{�p^���6�T��&T9�o���sv���X���Fm�u���o
��o�co�~�iϽ��WW�7O}��d}��QS�l�x�}~u���9����=�VL������s�>^��4��|�i�{'�4��B����W��wz.���{�r-�� >���&*yQs�X�ɔ=q��񖎉+����lǻv���;)�����9|n^z�؎�f;#\S�z] �"�F�>�+��}������}�=��'��V�c�z�ЕǴ�?_�<1N��<�2��U!�*�;��#����U��8z��Uu�|.%��9�?m _�����w"�ޯ��i��7� '�8�|�BG�����X���<�d~=�0�������7���'�uNH���_�Ë�)������:2��DM9�;����^�]�Q�uW��������������k��/ON���
� |���z@�9�t��Fz����F����2�+7ۯ�hEd3��ę�����5��v�R�S�(X2Y�:�����n�Ÿ��{��n�m+3�rO��[���n�p��F��I��jA��u�h�Ցp6�Qv�K17�R֫S<�8x�bWs�E\ �Y�9uEV[�߃�c���5�@��cw�tж�I����W�]Ƣ�o�#��v[�K�P��������v�G(
o+��7��KU�ʷ�}-~����S�������z��޾��:WC��=��qq�r5��/Mi��A��7�p��m~���+��������r&�'r�W���:��+V�D5U>"�ԉ������<��z$��L�sgj򲛏f�6&7���m:����&p��;;(�[���^����ӝs�?h��3�}u;銰�-
7qq�����V}�F^V�v�z4����}{] ��x�/Tw/j���xE`�ZAq���XL�|5��}��kAYT��MixN�c������+���~)����F�5[�r��z��G-���%�d�\��+��=���dγq�>E�!y�9~�	���2�yU�����u�{b=��n%ڸ�{h��g��.%�2�"�����@���r�Ό����;γ��~�k٢E�S���A�;~�_�>�bh�/_�G�z���o�� W�Ώ?Z�{��k�,�q\z��F����I��}ǽ�F~�_�)�,��!��o=�Q�zF��P��%	�m��)��v!$��aA���
ɸxn{}6��e����ӀvD�SG��<`�-H����ژ�Y�v��^U�A"� L�x��=�G]5Q6�=�#`emZV�̻��{��E�%б�l:
˝�Ѯ_e�Ű�sy�SB��Û/�����KGۛPѯ������6G�#����;�{$dR���-�.��;Ъ3���d��F@�6`�����q���ә/Ư��������� �nI5��ݤ������^�|z���z�"��W��~q>d@A��R&�����;�Q�և��Dԓ�ג[M�Lz!*�^��T�Π��5T@]��7P����MV��|7r�3���}$�쓝�א�sRP|���z])rpw�9p$�y�Rf|�l�C��+t�|�Jx)T�sowho1�܎���"��:��j��T5U>7���#�]���>��Ԟ*��W�챇���کs���:;d�薥����ט�=�1��ͧ��8����~)�׃���{�@�~���������wY��<�5q�]�v<Y�D��ZN�/c=Z=y;[7��=�6�W�=�������g*�L�(H*�����<Խ��p�h#�+\2U,~*������ϳ�g�4�6�k�}dC���$���{8��U0���t�}��q7��碻�z��ՑT�VMib�g|o\��=��;����_w��r����\΁^�eo�M��1�hq���]�/�P�M�]�,�����ɮ,�r�S��<KWx�)a&�N(V1�ir�J<X�Ŵ5ed��t�c�hv:Ս	[c
�;t��K���w��G���P����9����_�5(�g�o�T�}wih�a�O��hv}��Q�{��>��OM����㾿�O�ߴ~�@p��.��&k��d�,��\s��N{�y؋�xuļ�4g��
AdC�f�u8�s�� C�ʽIϢ@���we3y2���sC�a�{�x���`\<T�=%��n��ד��9I�g+�O�lց�9Q�&��Eϓ���A�q~��S�>=�7��3��� u�j�\�d�����` $}�T���FT�`TE�G�XJ/�C��?[f�\�����^yZ�v-��c<���i��߮�Ϥ��ىlق�ْD��Xs��x�}���Ӡ^Z��=T'�\t{yRM�U��y�\��l�*���Ċ��3p�<b|����ٔLg������Kא�k���R�x���
�Oq��U���k�����wg� ��u�p.%E4{&@zfr���/!�E�(&o��?�(���������"���˼o�>^u~#ސ)�(�{,
y���a8��UFj\�SQn��6��6�͢=W��5^�Q����%f��?Y�o΀�8�G�g�������6��nL9H1����GmYL]�U6q'=�W�[j�{�.ݩX/�`\���ʦ(��wt'\fU6*�t�eff�0��Q�e���ܴ�a��付�$]ɝ�:r��=��q�s�0�se�����?.������a���-��w�t��gt���,̇�������>�9olz����wݬwG�Bu\*�*6_�YxI�㾉��;������s���`E��t��L��f�����dGz��>�L��hN�mΘ�@=��=RQۉڇ���,_ٳZk�f�{]+Ӿ0G=�e��_���@V*�@�O+�\o����o�F?w_����q�8RϪ��mv:��XFF<^�N�^��*��5��G��k�)c��MlG�H%�4w{� �$����`��>LoE�䆭�t8��E����:����	��6�ϯ�w����1l�{�מuo���Tn�!������Xg�WU�O�}�y2����\惿����x��N�mW��5P.�i�#='7Js>�}*�q���YY����n%����Sȋ>E�ɔ=q����b�NI��/4��z�͔<�ǭ#�����~��*���-�ĺ5�@'�U#*&[ W֥x�t���^���m�1�^�>�u��߼����{�����G��
�zd77O@{uR؈�q���B�՛Yԭ/�����Z���LTw-V[�u�{�i�P1�X����4û�t����+vC���y�R�0�3�ʹ��ԩ�M��n�f�s�+�!-�A���y�Ix�@c�x������;t$x�C��[w|���sޙZw8����Q�x;u�Ī�.?�%"�f<��u�X���H�?m _��#���Xfa{�)�gؒ8�|��_ )�k�T���У�^�{�~5��w���������˻�_�&4�%|�׻#����z�,��I�z���+樊g���/�t������G�W�������U��}]��[�{��y`S{�TE���7Lu�z��}r���w�`1k��8�	���5�2�c�y����9�`zᜠ*<�%QϮ���D�Cܝ���l��tJ,�i�IõK���c����Y</{�^Fy�;+�C�@{dQ��>����u�n�{����3�=�w�1���ϣ�3��r�~Lψ�O��z�H�(o���.=TQ�*ߒ�e��]����W����ި���U������ Ֆ�^��
;�lO��H��y
�� ��(����Y��cw���y*�_��90����(j4�Q��6��'Q�{�+66�sr�x��c�ҁK�>��ܣm��s�Vւ�*��3���3���r��#�q���}�����Θ��:EN�U�ʈ����l�˝j}b���C�d-
�v��q�����^`]���U��ӵf�G
�y�c2p��v��:��e�;��I�4�Ƴx]���{��C��%���)����#�:����E&�0 }AO�f<��������[�t�+Bej������u�n{��*�����W#ogIl�:��VU`s�,a:�dϑ{�y>�e֘�����p��'+��)q��n|�粽���j�q������d�l�誰&����D�3V�����wgЦPk��at�^��=�}ǳޯ�wh1��C���^�p�X����v��7��VW�޽��j��)�Y0��{j�M�;��ݱ�0O�~�2:v�>s��;�f{j���nw��;'ЦtӟQ��z�6Z>ǵ��w��ZG����o�t_ؼV,ז\��ʞ�=^�=��U�i�6`�;qS"c���}�Ndl���jZ�Y�ٽ�1�e��5ٙ��W~l�#M��T��+�NH�x�0P{uH��s�:3��Zv{�}>�<M>�����g�ԭLc����N�W�m���^�ʉh񩇗>&:���4K9�c�P��������m{��=��>�5�n_��3�z=U 7�4����"�&��� f�|�Nfyf�摌��Ԥ֗��O��b��2|{�t�C���,䁫�%߾����C�)��w���z�K�.�T{dH�5Z͸�Ug C|&���ȝ�[�g���i��-i��ngE���MR�e}�6�x��f��Jhf_=��1e��wom��׻��G� ����bs\]\�m[�j���R��GW>~�9��e�h�vg%�dF͂n�f	�Ř'm��wj���S�9y�D�§�z��k�<�RU�]�0.Z�z�%hdX�i|A���x3��q����o|�^���n�v0-���z?�w��
?u�%�V�~�C����G����Nori���0���)��)%���܁[Ѧ����f�i/��z��WQV�Vn �����ܝ�+:0Z��[g����kk�)�uٚl�p"`����%����|6ht(�E�_7QgqD�u8���Ѕ�u�erzܻ�_Y��v��Y�A���>7�]�gd�	:一��5�5��R������_,�f菑� ���t�&&����_Ji��b��FL������1�j}2��Ƃ�V3i��9��<�s_:�-�= �x��� �2�M�4;�yԭ�+�M��\%�c�qՉ ��5������n�RC4,Τ�}*�8��J�ݎ�V�z3m6�(��8@̂v13�v��x�S���rE,�̥��g�`��{��D#��2�Yp6��Ւ�p�X���ݴ�N�	kE����p�i��n�y��{^]
km�\�rV�1}#sηO*}�\Gv���V�|��x�Hh�w؆I�t,��F(N�6����1�q)�|��z@a@�xV�W�BVPtv�:��Nƹ[��J�b*�rD����{73%Y3���c��=���ۍ��_��=}�	e�x����v��_E���ُ���t72�ۑ�4�I^)�^ۉ�NU��1܃]�7�e�l��q�ʼ�.=�������E�Fx5���NskgU�<��4ζ)�@n&Ů�����^�����7�����X��"l��'P��t4�j�n5��D�s�pBb�5�Ө���3��ݪ�EÃ�p����:ˤ�}���o�j�D�;�~��s��7$�(	������g\�-��_MΩ�_"С�ٮK���\6Ӳg+*����˩)�H�?!��lJ��Bdsewe++���^n�����gp����;M�ͫĝ�{���
�[:��GT��YwQ�w��j��S��#���d�#+���`�wz� u�d�Ljc1�jW�v���ײ%v��9V��0K����Gv|S7�An��T�ǯ>x:����ygIe�\�R�]�ZԬ��+�ܸt�נ���u���*���_r��i(�o�kwE.D|PW�ٽ*P[�óJ4iq�� ���n�A=���B�Wǣ[(����h�Jrҝ��뛝�v��z��']m�ֹ�Xd�9^�H��ojٱ�]I�Q��y�f����f�ɷ����� �/O)Ӱ���(�Y"ƍ%��Ѣ�$Ʊ�h�6ask�lQVH�c����m��AlV0��](���F�knj��D&��Ѩ�)(���DS-����3(����d�4ZJ�hѱ�TXڒ,�B��Qb��ш���b
Ѵl[\�r�&�m���Ql�"�[r�[
�E�Q�����1�h��ưl�A�`ڈ�lTZK�B��f"A��H�����N��%#�����m�.��Hp�J�U�T���O>帍�0�ﻳJ�����˧3p�w:oe��0ߘMe~���_5��c̿�O�ã8�!��|&+F� �G7�W<���s��Q3�=3��:|/cӁ�\�tޖ=�7Ł+/��Nk�@���c�T�g�US�N��^bt�O�>���qV���k�N���	Cn'i��ɭ+����#}7��X�����ͨ�>U�����=m_������9����{�Q���{MǪN��2�&��d���Eg��F�z��9v�-!�Ɋ�>����}m +劽��~�p���ymaC�����WUG�����E��y�մ�ӱ�e3y2�yR�����s�q��7��m��#�Jz�ũ��Q��*�?:�7����s�)Ϧ�@�Up�f�&X^9�*�u�9��߯���خ�����V�u�}�/�U`��� O{�LӑG ����'-l�h�/+���I}'�q����{ӯ��;ˏ��vPs�L�� 6|\��}U#�\��}�,*����O�E�qu���ʪ���vP��1�\�o�i��[�y�x�zK�ٸ��$,�&W�Ð\���p�z����	�ĸ��'��:s�b�x�F }����%^�7Y�ow)��G�Eoj���(��ꝜbS�2�O�X�tY|� ��̲����*4�:jfc��О�)��7���QpL7̽]���&�B�7:��rom��8��* s��Ǣ4���yEM�l]L����W��'Z�R��Ǭ���d�;��D����B���7��R&���"�>�Ի�)4�;Ng�K����]V�9��+=����̂-ύ@�T�����Y�:�Cyb�^� ��P���ޭ�����xj#��x_���r=<�=�: U�+�b���fw�n���j�9����d���Dz�ղkK��7^����;��6n��^�����f�l����v����r]g�5บ>�fևfׄ�cL�Ɩ=Ifd4ޫq�`gu��_c�71�}�G����o�6v����^���O�ϧ���;��:+N����[w����{-+������G�Ӯ�\o�Ǧ��V&��۝1qށ=���IGnv���W���������z�v�W��|ԁ�����d��ޝ��	��Mh��=�s�'��u���},U����ﺺ�^*�7�wR<6�]�q�w��N���|��q�6����M���*S��q��y3�
�Qcj1]��w�c�9�2��?_��{������q+��x`�
y�&������y����Tp�HSo�,�����c��zoD�qfVh}�N�tfЉG~��|�L�:[7�^��"��loMܱ����:Ȇ�<�,�с\jޒ�W<}�A7m�ۧ{��)�
g �Wbm\q����dt��\��%����+P��3@e���L�1��zu�	��~�����F��̲���fʳ�ĥQ��l���D����UXy�>E���C����_�i�8"�{B}�f�n������:N�_?O��K�\{�,�k�tTz] �"�FT�d[�#wǋרt_<�����s6;M�F��:b�>�]ǟ��W��C��j=�G�p�̮W&�B��94,��Ϫ��0zVWa�}��"6����,_��I��i�=�G
�[����5x�w�t�.Ϸx��y�x+�{fY���O|KGw>�$����o�xp�@�{y�����f��Ѻ��8�8��T�L���_���^^3�����^���{�kg�Ԟ^���瑃����Ҷ�V�X*}DlJ�=�t��}��=ei��F����rȹ�b�{$ϖ��\_��;�Ɍ���M��z�?e�n��]��W}uo����2|:J7oR����ي�ؽ�~��>u�yMƵG�����#=��EG��ߪ|�dͯӤ{��1|]�V�7nJ_������A�b��X�ܙ4����d���8�_�{�q�[ΚA�p��w���g����ɞ,�����>��D�b�g��Q	+�h�����['|�C�r�7�y��R�r���xW@:�=�z˗���V>�˫�=B��9���^H����\y{� �W���j�|E��v䬇�EC�(W?EOh��T��`��`���6vaY�م�ڭ7_�M�0��`_ܽ]�3�L7�ݺP�Z��#3��Y���ݷ�Mh��B{R�dz���q;,e�m¼�+���uO�m�:U��P�D9����1�fh���[N):{����9�O�U���ck&��ɝ��ƹ	��q���^}�;$e�@3gѽ���0}��g���7��;�h����-��[Z
Ȫ�&�X���g��wq���w�ynN��VM���½
d*�OR����#����ĻWy��c����v�D�E���}���>��|�$��uF�Y��a|}�L��GS����^��p�q���î]�b�����z"�cؑ:�y��� ��Q�&+ʀ��)�YPѨ�mCA�E&�x%���C�z�/�7����:g=;�ג�^��=�dy��e�22���d�}�Pѫ�e��*!�J<��C�by�T`xuoM�{��{G�[��W��� 6D�lTȘ���}�������K��,�4Y��ȁG%wl%�=��3l����`@�%��*y��0ouON�[�5,싫��d����Sa��p��c�������ƺ�,��b�R���O�]���Q�r�	v­R+����M��6.���
�o�Vf��ֶ�-l
ݜ�Hj��}�9Ĳߦx��֊�uNHp|ȁ��D�9��a���N%����P���1���=V}�﨏\zz�0�Ͻ3ީ��{ېb�W��Q�Z:ja��x��6�K��8{=qח�YI�|�(w`�2�����~���K��.N���. �<�}U^G������2���y[����^��B��:�WI�������E%�6�|�Q��=�sT3�!N������Qd���j�x��|�]�f�ӛ��ͯq�/���j�'�~L��uV~|���h�:�A�~F�7���/�1������q%���M�챗���/*�ޖ=�7X7=����/���ק�h�Gk��kk�v@��ʧ��ʍ���פ�n#�%��c0Ε�d�V��\����x�MK�7��f����c)3��}�}+=:?W#q��q7��nx�����&�)�-}�ZX2=����1w�{9�,5z�y���]��!om0|�U���-�p�����b���ϽS�J��~���i~��7Z�?Sg�o��O�,�&P^Ωu����9�^G���xqwH`���R�\�w=�秌?acyQIO��wD�L
�48M �SNM���3K�"�s�U}�ɧz���C�LqG0�լn�ˋ&��w#:�z�Q�^�*j}}�U����w�`1�8��^�Pq�]�7t��7n!��r���]]�Y�Tfʫ{� w�7sTv.N�"
��>S��g縭�F�l���xX�����u;����^/�����e]�;�Ǫ�6��g�w�r��?U��� K�sH�>��M7p/ҙkf�F��uC��",x{<
�T�un�du�^U~<]�|��7��ᐧh��#L�ٿ�.�}�U#+�L
��<��e��y��;��M�y�z�y��{�7�_3�,�;�{!��'��&%�p`������ex�6����"u�룞�UK�C����}<K��C��s��#��s"E[�nG�O�x��W��xh��Ovv��i1�r�NA>[;�#�|κ���������}�pG��&�t���O�f{ �!�/�
�s^���	��}[GC�݃���^��Ͻ.���sZ I��dE������&���'��nD������[&�4�>�y���ʄï��͞��|&z��5��`v�C���>�)�������H�>����d����d֖=S�{����z����b�MN��1�eo�뙗1�Z�<n!��G��;��Yl/����	������c�a��똺?�U�iSr����\ᮅS�l�%.������RБ���s4y6���KWr�b���:����&k�e4mf΁��,4��t�t,cWz���E_X)��u����ˬ���N���%.ɪ��7�)��w����2��|N�d���;؀)wt��Ͼu�Lu�[����J.W����8cc����'۝�x�d�ɛ��b�ù�O�,{�Zu1w�L	�YV����w��^�o�E�֏<�QV����Z�yzשx��芨�5��q�*�;�>�����Z�Utz�uw��ý5r���ڀY�^u������w��=�z�F�9E��Wp�&w�x}3}2����~ӑ��.��v{k7/ԳP.)�{���!����H��D���YU`M����d���G9�׼v��&/#6�EN�9զ��/K�H���8��Q��Yeg��"�����U`O�<����,ex�#�#ޏ���Φu*�����Rw��h����qz}���=y��k�t{�J�dUHɁ簂��]}뜀$$��O_y{8��R�U�^
��Z<.>^�3�J���6����ᐧ|ni��ꨭ���=+ª��(��q�o}p&�H�狀��Z>̈چ�դXϥ��9r����B0?���3L��k���j`w��fnB���N@<��4+����>�Z;�a���e�{�zr�d�F'X�>5���L;�L�]
t��5aqeфY�Qǝ����1��f�F(J����n�N�xcq�}��jo�W��æ0Ю��ѢLw+���-KU�<벂��)��j�u�E2�f[�X�4�2n��f��N�u"��cV1��]�̨ոDׇ��Z�����"��U�"��x�p`�e5DS=�4�r	xk�zn<�t�^�tϡzka,������q�7�R�{,
��^�.] �웦7=$z��!F���^�t�wݦ�!�^uKv��p��g�o��;�nb����S�=a� |�ī=���50�r�K�b��`��>��_PL>��}�d��P3Q���9U��i�>���:	K��ՐD�+��#�Y�*y�=���7��-�/F_����\f���<��~�����_Ѿ�O\{�BG��@(����Y}C��fkMW���^�0򸆽6�Ou�L{����v�N������(��ۖ�v�+v�~����b���kG�Y'��z��F�'e��څ��Vt03����6�]�=]ޞ^��B��أ������~���g+�%p��^�q7��nx����}98
�6�ɭ.�ɝ��된��>���xLR�C�����}�탍S�\v,�)�Ǘ�h�X��-��rpUps�,]�y��E��~�w�x<�����Ϻd-��w����ǲ��ĻW��Y�,�s��y �?������l�R�i.=�ݐd����+��� ���q���"�'J�'�w%�n�-�PyH��(.;��R9���L�0�s@��j%�w1�/�|=2j�Zl���]�>'��+��sF�]K����"���E5�1srm�Z��F(�(�?��韠��3;��&X^�vXQ��z3��+|�î] ��գ����N�k0#JN��K=�xuO�&pYQ�'�^�-��mCF��P�r�_>�ݟ{��ۇޫ������3&
���w��s=������!��(l�Rݠp�}�0���e��2�/Օ��V������°�6+��;���L�K�� 6l�l�,��`,-9�/�m��ڟ���3T{���н��m��g8�q�Oq�*�S��2��A��JȚs�:/Z�E��5�w�W-��q�|����U鋏�*��s�T�
��{r��UD�����C�(c�kv%�oP��;&��Dj�ǠxZSRXK�L�=.���:��Py獠b�ԗ�c�����K�Ӌ���v�+[���$֗��}^)+4���>9� {��P~/o��i�E��Mnf�Q���$�ۏU0�����ݨw��7��3[P�i<���j�|FM����7��l�j�>��а-�e�J7�>�����Ng'�t�����}>��@f�����0T�-8!�Jݜ�l���>dWZ�.�BX�  ���f��_qxꁥ��(���1LL꒝�:(=m�{�����P�\�M��1ɢ��#r�u�B��}�� �ӵl:]ga�@�ǩgK�hl���4���s& �q�����5��9۹�ܨ��yY�k��U���"��r��-~
o�*��� �#':|���۞z��j^zt��/���w�S�;�Ew�T�:������M1N�ۭ^bm���^7��]�T�m�v� T,U�>�N��{q��W#�E6}=c���i�E�>��U�z��3��b�b�gY��g�<���a%����;�~��Yhh��^�/+EN�­�A��s���Gz�)��N��X]�FB�ܰ�s�T;�.��=ҼR���D���O����w�O�c��ֆG�h���N��0NEb��s��������Nw#����㽺z=}I�>�qӟ2��O�߆Dt�}�d��] �"*�eK��<��Mb��]p�7�r�r���O�:���Sf�U��o�i�S�u�>%�lĶD6"�B�q��n
��ۣՍ{0�>�*R9�F�
���)��a��L�p��Ց�"k���g�O����z6`z�Rgފ�B:�o�qH��j���R;�a�t�.M#)�`�7|��#��Z������m��UkZ��Z�۪��m��V����UkZ��V�����ֵ���V����UkZ��Z����Zֶ�*��m��Z���ֵ��J�k[o�ֵ��]V����UkZ���k[o�UkZ�~�kZ���d�MeʮA,�c~HAd����v@������*� �Y�$��B���*�*�i�p��[jU�Ehs2�\��ibٳa��:�M����4 PPt

gT�:RR��l�d���6�+&��%qܻl�[m���Tp�tͲ�[0�UpcE :��E'�jZ֛�    "a���MB`�L��L4�&"�ф�J�� �4�#  	��`20110�L�L���R�(` � 0�C��L� �LL&4��&�H@OHhȣ!�ڙ Ʀj<<�/f=^�7� ����� �����!0@B0�K��c$ $�#^��O�����?�:B1!2 "R�T@�Iل� b!I
`	4���ת�g&#�=�_~|v %Q7��WU+����L���΃x
�P���OJ������e���,mf��蛴.�w�]	�4џ13/u<(mMX�eJٺ���ܙ�j��j�hX8��wF�ܒ�mLneՃ�.��";ǋi.R5�d�6��3�5�N�`T,H�ة�9r�j�HE��k-՜�T��}�\��ߓ�
:��X�t�7)�T̈́���Jlfރ�j�fV���OUl���Ծ�L�3l[���[�p��*�f�$��ȍ�5��sM�{z��-�F���Sl�����Y4�aȀ��2��*����`5$�h�@��oA87��E�V56biMc���mR�iL�Q1V1z4��V�F�U�Ʀmcr��D�A��iڎ-6�ǣ.��j5���'32:X��Gd[�R�-�^���`em�N��6,���ou7��X�֊-]L�@�,(��l�k3&wWbؼS0P��"�:�e�g�y�E҆)b{A��L"�Y�Jvr�<*�k�G6�k@�*��*[�n ��YOV���vBܒ��Q�V��/wejRUD����*�@r��{���	����fM�͗e�m�6��U�a-��GTn`�cK�(Ʃ�d��f��Ɇ����+�%Q����Ս�x1�oT!Tj���`
��MXŒ��Tw�ܻyd�Y#Iԕ��ցYPB��b#xc��t�4����MF4�@hRn��[��33���������"\.��R�C@����l�aM"�Q�q�wٚq퇣6�a����-��D�ހd��X`Ѽ�6�Sx�ے���:0��K�����ŕ8�8�Z�w�ݎ��������4$J9^v�U4	�þ�/�^��ǚ������k|��`�5����݀�v`�L��u-[�+���y2-�~�,J!�����0l��מ�.�}��99�T�˧x�d���H��oM�6���l[z�e(�3�1<+���wDۙ'-d���=��!t�"�}\L��c>�л\&�����i.��6�jW$-�r�+3���� �L�	�]x��6���a9G��5���Go�V5����aU�s7�yu#�לm���r�֧y��nP�ST"`	/�����ՃI�{�!�j�ĀMZJ�Zo�����'Vܺ���e��C���������ۗ�y��mo!R��=K��NB��eKŹl�gf��2�3l|e�/6�O��Q�:�wY��s�hQ���c����eD拂͑���έ��Τ����5��t�0Sg7gZJwiouZ�4�6���Ծir����x!\�>�;���u(���`ǆ}+P���nc���yG�q�3Z$���vZC����_r��j]�[(�(������x�eL��$������%6�I'wT�!�L��Η>�����L1e��@���/x�ǭ֛�cmQ��$�\�Wen�D�����2n���>6�k]�H�vn�O0��:r����9�������)0�9{}�-�P1�%�С��%}VQ��K�a֭������˵G2Q<.�|����M]e�u+�9�ժ�^V�d^����i��qr�M,���F5��t`����Sl� 6r��Y��@�3Ci��z�����\s��w�4L���׍3	�,3)2Ö����������8:���5�����	x�d�HI�EB�ω�� $��X͞���}uXkŮ�����6%W�A(�n��qeO�����Uh���������i��f��-�ܺ|	�$�5yB��,mZל!��(���g-�N��2�cl����a�~t�O�I%��f���6���g��V���X��m�(�QҊ"f������FK��2�{.���$m�jt.
�YΖٮ�c��C�;b�X �9������$Fe���Z�\��Zg�,�꽐>�j��Sxy� 2�Y��h�Y1s�B��-�y+z��lVXEo��$��:��)��R��;ab?�)o,O+6�%Jc����mw<�#��ۧ�7��ˍ��if��Q����-�#FQ�jp�]�n�LN�� �ҤV�r��+	���B��Z�.��pP&(+�01]5�X�6A�vf�۔*:ᙺ('F�d��F�1E��1�Y��Y
Ҿ�T�p�^���V�"i�M��im��WǏp�$s�'_�<ua�=����uN�"5��p��f��gT�wLJ7
Li� ^�&���f��:�� P�����t�G�cW�E�3��t3i�ˬ�Lh�^ˮ��l��P��:|{8QU�
�T�����:���%��um ���оg����^:��c��7;.����H�U�1Y��Н�\��`Lݺx%�Sg+[���m
��yXPb�SF����f#���rT��㓺�P:�#�_M\K���l,{K/��A��i��y	J��գx���k���9��Jk�-Us撾����)�IA�Ƀ0�_�/Cj�nӤ�-�Ư��I$�A
�03
��������>�P�k��(d�_�}?�{�ev*���K5�Ƨ�8�A��/1��՚��Ej6}��켄D�7%c�Cש�3����h�2铹��,[���gu�WG���S`��+z� �cMr���jL:�,p�bU���"�s�L5�.l�qf%���>gC��67ϣ��Ӻ*�K�������g���%�)5ٟ'���V;NFC[C?�va����ױ����*Έ�ئ�w�<n+K,�,�k�h����2���3:�8�<[�@_k�����䲛{�YaZ��H�����R�h]�Lo�u�*�c�k%�U�4vJz���f�D:���ݝ8�Y� ���aj�Ӌ������^{�
~lx��ks;'ݧ����Yt�37녀xyOV��Z��_��U�_��?U^���x����p���w�]���S�J�*Ӷ�^��p~d�f`���������6��O���j�jz��jH��D,X�e���F˫u�e�^�Nh��a��BYC�֫�+����y]x�=9r��<:L� �j���&>�1p\�Rs�������/�a��+ؖn�ǎ���@*?b���k�	݅�w\t</
9&j����5�-�b�X{�*ɹ�e�v��i�JX���]pa��v���<�a���*�ɖ��rPN���;$�g��p���wt��ܲRP��	�uOjd�Y�0n5ui�`��ٶoڧ-QM�r��Γ}k��|6@��%w*^��0�i?t�y"{�]��e�����)j�|���1������P�3����)}��8��}�C=_�V���>���`�����������s�p��Gkr!�E�W�D;�S=k&ƧD�Γ��Q���g|�����O^d�͛��K���r�N+[��ŏwqg�VCf�Š��&�vܨ��@Q��
��He����yJ�eҬ�2�W28�d+$�ST�f�Gxre1	U����=^Gh���%���)��qT�F��EU���]b��vX�U�U�M�KE�)m4R2��4w[���=��,�
�9t�N��vt��Z��|�-�G����������RCP��X� �e^c�p7��T�/�_��:�yF��^:)����ێ���~Y%��S�ee]Y|�Q���%���y$���-P��^���</��d�p.�뫞���s;�nM&��rR�,�{���S��5��^%{��q�w�,�j��MW�P�(�ܽ�ҵ�XgyT�]nY���=o�ۏ�%ww+���}�d/�@�����	$�e�@��
d��!&!:B��@6�a 6�ݷ�w�Hq�N�I�@�@3� e20�	��H, Z���$��TI�� S  E!6�@
B���n�	$�d�!{�	$����! 㶸ưQ��k�7m9\��4P&��J����\D[ǲ�R�R쨖y�8��Y]��Cbl^�#ؽ�&u��H~~���{D�V�>MEYӘ�+��I�b�I�F��xT&�S�0�2�7*";�N����`D��~���6�E5c�m��R�:G�z�-~*o�}g�����]���@��Oڕx��Ǒ�~�����Æ�4��1�=��IOg:=k�M�90�}뫼�y�_b����ZLx&J`Pz����T�S_V`�&� �f.�f2C:������7���e%�}z�ҹ1<�t��}ozA��/�I�kV�#����5usY�R<*ٯ
�0�+�d7��C������vBy��4�:�Ǭ.�>�O���z��P�+#I���D02�a����d؍18� �~SA��[߼r���}��q��͓c�:AjKVr��
2(�Ho%q�c�w�*S���5���e�����ZΫE�*���]1���"a���0~�u�p���_�)Pm��)�̊�4���Q jF��obE�ȷa�h�t�\ˏ#Ô�(ae:P�r�D�/1K��N�U�����h����U(^�L`�m(cJJ�ҋMD��j�EUn�E[���q"ňؗe2�ZJB��*�ևiv�hv�?���f��w��-b~�M9�$.�!S���_�7B)���$��l~�׷��v��H���x����bh
�O��v��
�0�VY�of,��P�%)R���"�ó|O{�+!9ʏ��)��U�ǝ~և%�0E�"|�׆T�h_��V�=���v{}��?��s=�=OoHR[���$J�3u�`z��{�NS�,2��9��59�7�t���e�U���85^>_2�I�.��s��x#
[j��#����u��f�ݾ��{C��o��G�#ǰ���6��5���^ymw�=�?	�xo=�Fm�ѹF��Rڡby��"~�I5�µ-��Ъ�Yi:��X�.(�>�a�[b��X<�]����g���YV6�Q��8=<�0|5ڣj�>���U����n�����Y��#�z$wޖH���T��{�f���N>�s9��a��x��w�d�ղQ�r�t�ZWtΚLRyՑV������׃n:c�g\�+��l�N�y�Tͧ��vL�^3t�Z�����W�ۉ:��܆���#�6Q��ގU�xaK���B,�<�c�ƷU&�zXG�D�x�
�Bq�v<OjF���Z8��7�h�=�v���n�CĽa[Kݧ\��@c�����dȥ&�M�΢ay{
dh}�VAl�}��K�e���`��,c]�H���c�X�PL&4�L��i)N����S��`-�G��XK�KwotK�B�]�����[FѺ�s7k�t�ˠ4?{���o��bȖ�f�1�h@.��"ܭX��n�R��$p�	a�h�6]g�tе�-5�O 1�1Q�?���`����CR�P��]eSж�[J��] �-ղ��5��񰕃k>f�y���3��ݠ]݉Z�M�R�q�����q]j��b�Z�d�I����+n��L�)����7�������0�������l������4��qwpb���R�ma�K�{�o4s�N��[�E�����4�!�Z<U��"�\Xf�L�f�[!�uڳ�����S8ι�k}\皖�L3�w�e���3Qfb�(8m��4�	�4��t��I�b�Xe�n��q{ա��o\Y�v ����E��)%��;o�f�|T+%=��s�d1���fˤ���Z[���N�4�U6�B�w�1��ؔ��Q�uVKL<�m-��Z��8a�Jd�5-�Ы��*(ob�ઙꥱc7\c
���ͣ���h�).�33Q����ۤ��l����Hp�L����V%��k�u�pu�,�b�(�yy�$�n��-3��S.�B(����a��Rr�b���M��Ô��L&��2��Jd�\`�Jz@w�z���5��&&�^ڵy��w��x�nN�����[6�N���E4�hR��2�nJ�d��i����g	�X�YG5*���\0Ƴ���8I�h���S+��]�-;u��,���/,8f�o���$��m;=��	�Z}��S�n�󩘊}l'Ի@�w��ّNn�(RgO��l
C��اW[�&SiL���$^l�a]��h)&in�a�c�U8�d��g8f�*t�4�v���1�8�%��a��A��r[�z�z�k-:�R�>�������w�(_U7��M�AhJyp�Cw�`�CuP�����,�Km�:5QL"ɦR&�T�x��L2�bΜ��u�!wSl��Z2���m%&���:�8t�l�/�:���	I�-��6'"��Uj��RWTs�����Z���rޙ;%�k�C	˦���hm6�]M�QNs[Lj�)P�-�U��-�ͯg&�]�0��i
B�ŝSGWR��L7�)�3�(ZE�:��p��%�l�ێ7�K��M9R�)f%sC.�����o��]�8�Zr�c5��I
��d���;� �2����|b��a9KyI����3H]Ӄ���{�+��ܖ�3n�(d�໳,�b��)k����R��q������q���ǎ���+-y�g����� ��1�[01֫r</|�^<�&�f����ࣕ���g	�H�i��"���4�r�*Y&��=\ݯ����8V�@ggc�d�@J��>�J��i��_Q�<qDܠ2�L&�S`����tX:j�m;��<[r*@Y�u���X�6,�9�;H�\��W���[��wgp䋻I�ԓ4 �'�B��ë��p�� �� P�j���R������uw���QC`��X�������8�7�O���U$e���x=V��P�a�Z-�Hf��x^��%cn��� �r����S�:��k�m?Qݺ�ydV+6qe%���4"�g��Yq�ؿ_�r ��4Y�\����q�>�s}��Ѹ�e�� jgO����`IDj)]����fbr�zs���_��L�Y벙���~%�j���	�5��[���Ao�<�ɰ���Sn�T�6�bD�&�Pk]�{ĮE�Ht��P�x��f���j�'anTo����^Z�X	�)�CΞ���"[K���I�
��IM+\�oA�/���瀟Tb��f7?t�e+���1y��ek�gmc}~K:��o�S�[LN��V<z�j���oH�N*%�}UW8S���(��{��g�-���{Z�X|���Wv�����Ƈ�z�,�/E�Wp��^x��r��������y����B�<M0vzY�^b*Eι�Gwm��@B�6�~��Qo̯ _ �:^����4#������ߏ7���~�hr�g�K�.�b��;+Z>{`g�	8;��Iye7�)��%gE"6�[�����l�Y�y��������m��.˳���4����\<ݺ��ވ���8.ʾ\2>0ϻ��'���D�tFH[ie�X���y���#E��4�"@��W�8݊�xnV�'���T���9�m-� y��OQ���ԛ��^]D��މt�KT~�|��*���ޚ�lbt�lC��8�Е9�.�P�4������B�j�!uޱz{��\�]��uv^��(0S����M���
W�2�0�<l	wnd�nƲ�������O��+�V�����'�yY�M�e0��S0l��Q�I�Һ�d�,-�\H4j�#� -��-U*�R,��KE�����S)��������{޺�3�yֻ�3������1��늭;��y���eA��� �����G�]���|,p=��>�	��0�ϑ�yۦ��_�54?��z�>K��A����{R�:=��X<���^|�ih=���	G�	sp����,��r������[9��3'J}�7�������=h��ƚ���MDt�(�����q��C��zw��J��0�A�^����A�j(�vwɭ��o`*�Te��� jlvhUѭV��!j�֥�Bՙ����
������kmCk?���Ҩ���X�{�1�א��&S�Eh�n-�uI��$k���xǖ�ZkE�	�1�W~� ��*8+Í�73�B��z|�,�$�h.f'b#��t�hy��<����ܹx��������,�8+ٹy����B�y�ˑ�{�u;	�ΎgL������U�{��/��C&y�+I��$�*<�Y�XTIt�Pw�Z|:em�̠(t�"�Z_�K	��iY}V�J�"\���.�!ka�
��%����Ov��Z��Op���Q�e�^�}�R���	�t\��Y��ufa��%�����=>GO��F/Ҡ�gʵ�i.�Y^3@`&�F��\{��5��)��yWzޫ�|:ۢ+���*�K�S�ce�����-�w)FJV�4S�YC��:Q"��m�'�-:�.� =V�����=}���U)h�goî`u�X��ř�b6��i�#��*�H�e�^��]��;oh^������di5�#���|���z��N�]�pn�+���^�	������e	w����FLDu '/i���xk,2Ŭ���t�)�K�:�rۖ�b��S·����"*�(���������]P���T��[
K�����U*2(�m�HʩB��tYOd��'%B�щ�|z�]�����ӷo�0�AE�yg����v]���%_9����_�� �e!�6�)��JH��l�8�!�S.�e�����)n�P`��?W'缵�/����E��8܌]�w�+�H#8���*�EQ��q/���9�N�oz�v�ʇ
%֔0_�AE��?��uC��1�'��`�ʜ�f�"^�B��q�A*�����Yh�;�d1�>���@^��=}�������9���U
�ʧY=� �$�y�d_�S
ˬusʕ@�Gr����gB�$Tf��H���7��'w)�-�DEK�p��T�u8U��Y�{�j������-��z`k�$yL���3,��hYV3y��t��a��O�[��~�r��3�l*�;�x;��z���q�J�!Z��>2}�,>D�����Y�y�������i+�,M�(~�=f?���x��B���5�p��|o-�uz��b�F�7EU<��fZ#%y�2�K����c�$�7a���<H_j�� {��e�H�[���y�0�����f/V��9����l��RX�D���7�N��g�V4��ޢ.*��d���X��棧�8{�iP�(�OU��&�5����'��̚I�-6�^e��I,]�7�W>ͳ�f�9k�r�O	���+F?+My�#CJq�N�I�Qѯo?� %p�)�޿��^�;���u�my�[��D���]�G_���[]�6���A���Ԧ�%�C��n����}x��|�a�B��#��kEL͢��*P_2n�"n��2]��!�y�,�N
� șF���b�ʶ��9 v1����yt	i��j6�9yl�*���ˌg���M��UesT
�T�
��UQU�*%���PV�(PVU)(�����E��ED�
F$J�F����X�����t*�B��|�H{��U-_������!ݩ�wdE��x9�B�����}��:ݽ&;��B�j�x{Ba�<ko�E{]�����Q�Ns7y���0�b9�3g(yƩs�//��YX����(q��{�]�+�ydI�FT�i�m3���r+�u���'�,���<�!�����mC��\8g���5P�������������%�xٸ� 1j�7W��H��
7X��Sk*����#tk[7c�"V���xV�u��wYRػ��E�س�m�2�=Qۻo���q�t{t���"�Y�Y�Ln�{9�V����?Y֗Z��DF�}�����=X@�9q�˓q�$�Y�oxM���,y�1G�z�S�>�4uVe�6��½7+`�.�M�ʒA��cG�%�;��Bhx]5vh�l�i�[��L�U�ɩj�؆��Z)5
�^��>NR���酸c��nz2���-�&���^�{zr{'7*;f���{��
�1�Me�f
2vS@��a "���Y�l��׿]7H�T��>
�Y�6���!�{�踰�J����l4<Y(�s-��S��6#2�9�������i@v�!��Ƕ��(M�P�5�f��:a3���n�N^�:A�ܿ�z�G�:�����<Ǜm7.;��\��6�cA����3��\�L�1?X�_s�SHWW]kw[���h��d��j�^A���eG�u�suʉe+���(��n0�E���ݰ����6��brh賷\���|��5�{5��d�aE輇VCL
��4����P+@�L�j�zq���i+S,�-:b�YU�Ì�voY�3Y���k��(P��-41QX�Ȳ�Q(5P)����,\% �-)�Uc
JE��B
�E))�R�-QJ��J@YM%!BN�>H��)
 � �~޾�h��C?c�̴���t���.�Ƅp�3�%V<r2)�\bL���b�.
�I�)��E;�'��>��:�����{E�
b� ���ļ˭v�yeg��w%�N�5�:��&V[功4ѫ��-J���;L�^�����3>dg�m�2үa$a𩴶�W=�ƥ�h��u?d\C�P{2d����o.>v>sE��s7��=3�Ӥ
PA��]Ş!eE���ݧ������/+:�$/Su�Y�ǒ<����٠�^��~��_������_�5�+1i��SÈ���daq�X,N*�.������{G��������x�Eh�<��%�S73��{[�:{�^s��OĎ��eŖ�%� �����:�2�j�V>��5䋼8��2ǖAv�KZC)����:����y�5�$���Ғ��|w�p���HU����R��ru�v�)�bX�7۠�ŃP����g�/�Ίf}���ޯ_�;��B�S˯���{���y��� X�D��aK0�h�B_(OĆ-�C��kxƻg��v����݊�uS�X�}�-%�</Yް�9皺:xȱ�o15ْ��s-�9��5�g�#$�Bqo��~�kŕ��.��Vs�ݮ�(�TjMVY������廩.���x���J�Z�#֚�ù��36��B��JUt��9�ʝIs#6/�Ⱦ���0�*��r�{�������n*P��y�p��I��9�5� lI�úNº��bo���'��>}]\�B��u�;�z*X�\�3���$��,��!���.�e˨�(���U�e�c0�)i���T�AkT�U-+E[H��vV1M�:�[�}͹����l�s���V逗�ǳ��G��e�]t(�V_�KV�{����ٗ�^l�ܧh�Uڴ�=ӑ<��)�X���Q$��.1�Ab"4Չ�5�qJ=fѬ�����[���'���ެ�X���J)*�u�&�U��©�QJ�I;��d�T�u��L���䷕~^x���ws�:l�z��o��-��׈f�6D>�	G���l��Q���-.Xe�f��lq��y��ڒ&�����Tn��"��v��al2s�a��y��鹷���(�z�m���#��};��ٷ~z����,Ll]n�L�l�Jv,E��-��	Jg�ܼ�֋�������w�,���y[��ut^
�s��u/:�E��1�y\��˿e��B�!k#����;ϧ��;fz�|��^��KTL\��)�Y�B�r�/�a�!����D����_�y"�$���sn3��f�}��2������ ��\��ޏ�����!ѵ��J? 9o�9�5o�N>���~���]�$0<�r�n�Ң����ul��kb�'P��{�o���g�>SΊiUU~P�  ������ I�|�S� 	;LQ�"�v��q���qY�~�>�3�'Br��$�p�ubق^"��P�Hw07����g��4�%sA���-�I$'�$^�hs��|����v���=R���OүA���l󑗊�b����]�K5�e�7�#�÷Ff�� '�_��y�ǳ�� Cd��  I�O�8E�Ig���N>0�����4��G��?�����3��= � N?�J��=~�*N�%��	a���5>�F���1�D�<��+6�W����z������w���z\��U~�O��4X �9zC�x��ބr &'ɰ����r�!ΉE����%]��f��f������  $�I+�k�)�י�g�|����^�8�����!�OT��z1��Y����~�w��j;��ʀ I����F�����C��w����������RP6������k���s)2����|����������zI$��=�x����Y���va�3��Q֡���;�	3�P ��� �ÏŇ�E5'��G���ِ��c$��?��M�U��%����ܐ�H��(�6$���4&?K����J�|��2B�kT}��aUvg&8������$�����g���I�\�I!~��$�����?oq?gc�#������'�,!��z����">G�Ogo|�����@�0����l1�?iRI$�������QROO���~� 	*O�!��x�_��ϗc�OO�P��t�	gx}�oP�a��\(��4`DB��^��3���;rנ���Կ���Y��A�!��N�� I���f2������}{�j	�l(Og���(gu��\P|�O�`�H0���O���?I��	�?o| '����!��v���jg1ԩ8��nz]��;�P��OȢO��t'o)����H�
��@