BZh91AY&SY�����_�`qc���fߠ����b_       0                    �               @   ���I&@     �    
       P 
   
        P  |J��RI"I�*��R��"���%"R���UQJ
�R�$�T�*�EB�B 
��
D %�  
H�!R�Pw����r4P]�ź��� ۹�¨-���9�
��ܐ0��  C|   5w��҇�7����z$T�� ��z�i�`�J�8:��A��s�I9�
7wW� ^0�&Q�`�y��҅G   ���%"��R��RB����D�ƪ|ɯ�����׺c'�wPO��绡J�}�BK砥7w}S}b��u���|�yy��4)O��W� �mO��O&�� @�  r��������ǞATsХ7wO���t8��{��6=�� yޠ�� =�wE =��={ <�=�t('�  A��4����I 
�$Q �JR���g@}z�U��s�E����"\�ݝP�;�\�x��N��O;��==�%Pd�   ;� ^����k{� 3����w�h��x v=� 8R�=��=z4 9� ���
�    q�(�I��"��UT��BT�R��ԯ��v���O{C�w��W�l���\w�<�=i޳�`zދ�)����` �*J��Pf����^P  (�ﶂ�@�;��w` ��u�@.�9Pn��� s����� �r��݀>x@ 
���   ;�E�(���UH�| �>@9@݀r,�;�*+ 6�� ��v uwR�' ���  @�   =���݀w
pG �P9 �n�9Ă� m��7`��� ��     (   ��)T	�=L#22dh����JJ��`��0 &?L�U)�J�    �%HL����� CM  	Oԥ!"�@       D���$�A0M&&�h=Mhښ���g��_�)g�O��$���K��j�ͺ��k�Q U���
�
��"�� *�#�
 
����<_�Dh���G�?�?���D@`ʤ�I�ՠ�
�06S�1TD��?o��o�V
����1� ;��?���b/X����*�z�^��Q�z���T�z�1�)�=`�X#�(��=b�X� ���`�b�1S��z�^�G��z���G���(���bX��*u�=`�X� ��`����N�S��:�N�G��:��G���N����W�Q�z�^� ��E�m��b�X�u�'X�	�:�^��E�z��"���`�0���z��E�z�^�G�E�z�)��b�X����=b�X��
���b/X���:����:����8��B0���z��G�@:��S���1S��z��A�z��G�A���i��b/X��*���`X#� �֔z�^�LE�z�^�W��|c�"���b/X�u���G��z�m�u�=b/X#� ��=bX�� ���`YlA�z�N���z��l�z��(u��b'X��*u�=`/X u�<`����=b�X#���=`/X���֕:��LT�:��S��:�X`�X)�
u��1G��z���C� u��b�X�u��`/�A�z�J`�b�X�
x���D����"u���^�W���W�E�z�����`�"b/X��`�X������z�^��Q�|`�X� b�i����b�X��"���`�:��� �N�@��<`(�TW�(��E�"�X�0E�^�^�@^��^�P^� ^�@^��E�EcG�DG�G�Q � :�Dz�Ez� �@^�S��z�i�b�X�� ���b/X��"���`����"�b/X��*���`�X+� bx��%G�{�A��{k?��i���v@Z��e��<�T�Y��Y���76d�D�bÐ���$P�NU�:E%q+��\ހ���Y׮L٭�0-Ě�M-z��Uaø&�G� 9w��w���:�r�b$���X����'i{ۋ��>KwtO�c��^6]�s˺�ɡ�	s�\�h�)՜���F�L��5��B+{~��C5lV�������`��+5��KX'\�y
�;Mӽ�:�}p��L.����n$jѺd�!�8����|/f�����{���*$Fhk�ĪZw��%όS8���z@�7��K��ح�i4�4!;8�[Ov��cW��5(��(��c;^�ڶC{�&�gMd�kw�d۫�(b�h��{�`xnY�G4,,l3nopp��/l�)�����ws�<NQ٩�3U94�nq=�U��s1�	[��R�����x��T0#��h�%[��U�-��܁ʵ�q��{N��WN�N{4�[�-.��MKk�J{���!�cU�f�иp]w(��%�d�D���u����:"2�Z{���{z�p�$Gӵu���{v���q��06��.O�sn�^�n�u�oR�lH�3�g'@����r����~�I�'dO���hoy��ͫ�S�t��ϓ0�:�����El�q��f��C5t��n�@sV��g��{��ɇ M�O���t�F���1�7^;��29�h/����˱��n-��8�r���e<O̭]V��م������aΜ���A�F�����ۮj���/nټ�zLm�BU�,��`�l��f<~��Qė*��]�6�P�9b,<2�\3A�܉���Ů����޸��v��� �f�o�=˸\���J:�аZJ{�}q��y��죻F]�^�����F�F��)���u|��oy����x�`��"��&���[�d�3��sD�rA���6�u6an�gGR���ZF���v!������<�^p��3xg27���wm5U;.v���xad���K(ZJ[�ڷ���-:���Z�$�68C��-F�A��=�\�4nk������ѹ�wo:��[��Y0����t-��ݚ��p�%��{�J5��:^�4vj�s{8=:t�y�g.��淣�7�JE���b��弻�4���r�+F��n��:s)�9����6�{*@.���e9Or�-�\�i��&�_p �I��ૐ�#�݋[�`W�\��m݃srϲ�������D-��ZV��R�̎��	(u8V�����;!n��!+�4N�wT�.�;��
���5ϴ(��P�S���wt���KsT�@�Ѕ���b`|����]�<$��l8��3���T��*1j¦��0��@�h���¦�:bʴ�qJ��ѓ�̎�����.U�4˼4��8⌨�\+w6��O]�K��u�m@��h0}9ɲ(�h��h��:�[��Ĉޜv�v���E\�j�x�aH��Y���%���<�Uu�ɦ$]ݴ�U ��wp4_���o	w�=�٨-(>��t-}&�F`l��kU�e��9�c��ЫF!uϹ��V9f�&ƴ���]�SN�v�(|�Ć^¦�ɀ�	6P���Q�Ë__`�x�D2��l���t0ԓq��9C�&��	x��c����=(��#�ՔK�:qn%{�3F�\�sL�	�Z�ݻ�^M�vZC�ڸhJ4m�0oLPt�]�.A�����˺d�+\M���/�����F��	��|9�7r�S+��gt����w'_�դ�[��m��[��]�)���eX���p��:D�\Uu�x��!	&�n9�N�+Ms{&Ñ�׻�Z�'t�]:��òA��4��u�0���X�1-A���S{K��P�X�~@��f��o,R띺)�βp�ћt*Ƽ�b���PP�]�5b��3�S����[� �#y�F�X}<���4���ݭ�����LŶs��-):a�������m��v��zu1vP��h����۳;sj=ҡeZ/hݡ�M�d�Cᮒ.[���x�iOw�6lNAn�����74��a��Zvë*w��U�󹔦�D:HC�/e���r�5t�!�h�&ƞ	Jp�cޅ��~��ò>�qf�q?��'YZ(��-�x��Ѽ*Tޭ�3q4�b�}�>G�n]ΚB-�Y$����ȍ��/V�l��u� pPr��u�Kwy,�VF���L�c��q���n�$��pC��.�z����r�b�(s����i^��|m=�Ļ��.��Ʌ��뛑Hy�(@V�Ӛ:�d\��B����{�����v��F1�n���eׇfu�&�d�}.��îs�&�;��pu�'�X*���owl�A����([��;�f�rg@���o	��h��a��&bG6��f�\��;�mD͘���C���kN�Bˠ8易I�nǣU��垧�����-*�F�)�cp�q�L�.�઺!�/���qe�^qƷB��v� 	�w~c���9��T��˕�� E�8>Y��ߗ]�D���"��1/��o��^1Z���� Ss�����-�0N�9�*�k0\Z��M��w6|�u��1�T\4;�V���\d�r�qct�lΪ���͗r��= +qwӴ��t᧪{��d`Y�yz&Nq�J�wlk;�Pw*І���f��oWX�*������:sBmO��9�m�S)�q��
�jGN�#@�۷@�w{{kۿsgo25�x�k[��];Ӡ=sWa���ju����넘:�&0�^�ƛr�|�`4s�:��<T����U���6��p�u��^��4C^��~Aq.:���_5�*�ض��7�Z��&^�w"��G��-\�2,o��U�!��u����t=��]܂3x�i{��݉`��Ŗ颶����hx�uܹ��`Z�Ei�O*;J�"����!p6b���e�VF�5��7oi�ю�277r�eѶLN���9���l�߉Bcd�A�4H(�S�S{gn�e���v��t��^�b��1b8;e=`�7DĦC����p�{X7s�v�/_s�y8��Ñt�q-otP�+s� :���o�nLի7#���YNvpZYU��*P9<���ƕ�`e#[���TuĚ��w>U���F����.ţ�1
�E*�`�׫v�FZ9'i��f��N�0u08�5���Ӥw�领������IF�]ʱ�{w�L�5>��4����=��;����`�	��Bղ�z׈q�����zL��t�ܻ���ht��%���a�� @����X�	��i��]��B��"77�TL@
��� �$)r\ih�#��ػb+s�;4��a�E��!�˭���!1'�4c0哔-����[��ss*��\[�i<�"��-|��W��)A��i��t�����}��9�n�.����4g1a �
��X�ƃ��A�3���(
uj�GwebNVp^!O��!]ԍ�x�8�YOI1��\7��iX>{�'쒓�]]�%1dMu\Ίa�r*��iʎ��-=��v�'Zx"+L��/M��N�X��d���=lG8�ܫG�6r;��Ϝ�ϒY��to5���du�������oUN���Kv�>���8d.��@�"���/"�I����y	%S�~��8k)�w_9�O, t�e��EɅx��1�Ţ.��s���Z�`V��7(E%ʭ���6
H�ɻ�7���e��-�w����g��/��`�D���qƣ�
t�v��b�%��>::�F���on$�%�wT������;�L�l<5Z��L�3S����s��=�^�(�獀�,8��0�=�B	yD����<���5*3n_��.R��P�{��=���4�ًtEb#���zly���:�;k2�x �n�׵RTb]�3z�7h���s*CU�����!�fj���=������ ѩ'��hlR(��h��;y��M1PT�5��7t
7{��sRۇ5z�{#�x���]�
�۽�κ7w��v��x{��7��wfu�I/��'M�C���uXN]�̋7�2f�{Cs-!e�)�k(鴡�qa�Jr���TM�ڹ�xZ_��t�c|8e=c�٫�����Ɖ�ub��v�^0�ݖ�qXP�Ox`Q�ɇ�2#s�*J�U��$��{�x�+C������-"-6;��NT��׸��2�|y�3z�;��vл)D��n)����-�oH�#X4�]Ƞ�z����A�wOQ�,�c�dl��Ƅ�GZ�q0E�[�t�Lg6�i��]�P����RP sѺ^2V\�N�d]]Tp�d�q�7[qIm+WWsAZD�:ݻ��v�# ��eԬk][��2i;([����{��
�L�&k%�z�.o-�ܐm��8�B:T�ː��޸���ni�۱��Hb��v�Sz��W|�pQՏYɇ8�ۡ��s/���h��(�v��l����Ya4i�X���r�#��S��tŷ.v(&1{Xb��_-i��Ν5���#������xb�M=gvP�����6�����$�:)��3K*
B�Wo&����-�������G}1���u1�)v*��i���X��;��9�һ�նk�6�Үa4nvv8��r�SM`�q��AS��oBٱs�_v��A���ݚ���v�ɴ�(u|VZ���p|-�����#�C�bQ����i`��=���;�ĳ���q$� Y��:�ܗZ-�44�G���U2� h�K9�G	�i���﷞�Xc����SS�����5Q��u7��J��U�Hݳs^��P7��~+�z4�8P��>�-���@n�t$�*9�AN���δ�մ�B��w�{a�3{�W���	��ж쑣��w'?hk{��vpUv�}��sC�O�!KdG�Z�X��N|m�T�KC�;�/����.�+YW�������ڢ�s�ȭ��-E�+`Q���E��b��gA�w�A�>�iă��%��\����,��8��x΃gW~��;��7w�Hr���S0vV���K,�X:,�F���cD�BgpH���ڌP.���L1*�����%�CQ����I�7z�#�:��4�!�qa��G٫@��{黯�L�zY.��r<�Ɂ�019�V�&��(��7�]R�Ͼ��3���\��4�� ��'F��['���š�yqͩ�o<i�%�Ү���ۓ7�,�ۋ7���I9����9���+w&��\m�}ܧj��}Ӡ�7��Q}��*��.��lGV[�F+1@�8) �a��x��`�<��[�^sO6z��i2D�;"�@�����;@���;cΝm���8�se��:��ݏOM���z�]{e�:\��\ۣ�|W+�i�s�;ط�ނ}4��F�Jhl5��ot;�rg��([�reC�m����oӞ�fh�=06]�xUg�{]���
�{5c؎E�ub�su4�V�SNG=ή���>�j�#3�N���i�P�����-�l��1�1�Y�[������]
۸�\��-�T�!ۺ��)�m={OG�t#4�Hw_�H�۱'a�g/rN��b�H�ki��n�obV��ֵH�p��L��&KFˤ�5Ϸ��>��(8����
u��я�@�c������@Ju�'��E�Bء�+���$(>M���-�wq�w!ȯ��rim�� X�v���X��S����˭6�Ϸ�mL���]�׷��:���ӊ�%A%�Yp���C-
��/x,�̎ĩs�]��]��-��O���ֺa�F�u�]�;G������3{�tcGw��J���o5�l��ݙ�l�����W8�F�}��]}!3v�v��ȥ���^������5�|~H1��޻r�fh���OLԉٛK�;Cp�B�Ü68�s��1�ͻ�'9�a�)�>᳜�%�Tꆵ;7�l/�pv�M�'YBc	��Qv�����p�c�����oTu�����*m�'M�:����4q��=$[~Ol�N����^n��0i{�p@рŲ�yW]���=�ɨ��Ɩ�_ax�$e�	���xh]h�n��Q����;�a{�ŧ6�)���+�.�g	�V�x�xV�{�I�C��0�t0�蕣;sq���%7[�	���&kS�Ń+�,�6t�;U�bU=�����!��L�Hp�*u��w,4�;6��ZU�e/�y���y;6]��	�&Zn�Ql7��y�����]t�@��]4]��ϵ��>���G�W�;���Q�;�S�_X�L��A4O1)V��Mj*���K�A�ӄ��6�\��5h��'��_K�7�6��o��N��
�uD�Ɂ��A�Q�_��I"��m=*s�$`>/�r��W����ͱ��,c _<��3�8�v�����ܺ���E���9ۜX`,���ZOQ:pĦ<]���
����6#	88�m"�7��7�c�5�w��{t�g��n��aU�xL;���y�4��x�����]�Tjv��W+�z�,Ҧ�gkZ5>����ɹ=��/9���{"�|]�aԟh������`	�<a��1;���p���f�{��ad�ZaDu��'�r��۱�N��t9���z�#i�9�O�}�!����]�w4�k�t��Z0Ll�sIヒӴ�"D���~o�N�̢����\*�����F�Z���X����7����C�}~ÿ���"�낤��"�"	"�� Ȣ��"� ") �� (*�"�H�H��(� "�"��� ) �2*,���$�� **�� �"2 �,��Ȃ,�"
�(Hȩ"� ! � �$��� Ȉ� �H��(�� �" H
$�
*�H������"#"Ȩ	"+ "��H�H*�
H��"�*2
*H�H� )"�"��
H�"	"! �"H�� �
 ��"!"(�) (�"H�H��"(H-GU�u�EwGu�]t]R�*H��(�"�H������k/琿=x��y.�J�Պ�򼆁�)�w�BYU�a9h��_<��\�-�+��M|�xI�ۦ��٘�?�y=a�q=S>x���>dacxH�]x�r$��V1����1�(>���4�y���ױZ������a<�T���'�x���#I��G�z�*�I����ڠ�0bx)�xMM��&�)0�m�(}�Trw��w��
1�iu2��1��&���J�76�חy^kn�'���B����V�UcɌ�	�T5���ћ��)�>x�ǁB>_�y����@A_���h??>���?OE?����s� P�lUD���~��q����o����Lx2/���V��y��#sK�b��0�g���(P��d�e·.Z���39��[��#f�W�pKG",�X�8*rnw�8��|���s��=�^����k�
��t���/03qT;-��=6y��~�Z�̔{6����x]�	h���������ܯ.{b�&�^6 s�i�Ö�q�^LЃ\m(H��!&m����9�p�d(����vB�C*C	�@����B�W�^�,ҭ�7٫�0+��h�.n���'@�Q�ܡ�q�۳b����=�n>��
1f-�����Nϯ�N�\	|�d�5�G������\�K|u�;���P�o���:��~��[�.����8�w˦�9���B��\~;6��ߟN�Ӽ6?M�o��<;���}�W���4�۲�r�8�f��.Փ��[��r<<1���.ꙶ�_{F�~�_iKd�p��y�Ogwk�,A���Tpg�c�o�n����O���g�ڃ6��Rl�	�3x��\�|�Z��w!��7EА�8���:{���Ĩ��q�5��#[��獘�u{ed�e��Y�m�r,3�-�M��򓓧.�85�8�[�eg;3]�Cz��1�}����+;i^�H�ܡ� �v����=ў�i���4a���������i�[��y�Ѵ�oN���~Y�[#$���<姬Y	��F�=���=g*}�� u��4���ע���,B����r�iy4����}�z\����n��`�2�k��g�7
Wa/����?���v��
�Tݺ��Gq&���}; R��W��޼3�}��Yx�\F��	�����⥵�t�{ً�E�&O�f�,���{[	gL�սA�Ț\	\틯�N�]���o`~�=�W�D���J4M�������v�,�>��$ž����:z�.�N�nW<����1o�0ǎ��S���=�����Ns"d��}�=��y��}����+z>`?s����t��f`�wՅm�&vxM߃
2�5���o:U�!��s��vwu��2���/q�R��v_�H;}�f@�=�C�_q�F����j��Fi���]��#M+Ч ��(2g$�c��ܥ����ࣚ��E�5�����f��S�1e�XTd��ԋ�5�����x�8����<����
�`o�wv����u��T��s�w�5��������v�����ofx[h��$��W.׀��{I�{.�k|���������dɝҽI��3��_xEg�7)�. !�\��I�u��i����l���髗<^"���醷��BWG;��՛��7����{���(�����y�~�~`�nX][yڲ5�Ʃ�wy���n�
�V�	�V�F� �v���UV.c EI2��8�&k�æ������@�⋋�����Y�0���w�o�ܽ�$��~ՑU� ��b�ΞF��w��u8��x���3��e�O{O�\�&�g=�n;.�o���'�r�l���:�=��w����܌��t��T{�q�}�fa�{�eه�����y3z)B��\�\����2\@��7�vx{�*Z���Ca���Y�'����{����%����݊����yH]6h�u	�N��ᩞ�]��n�S�|���\�pH���-��9oteQ=�2�9R�|G�$ͧ˷������bz1��´���707fq���>����ob����3�{�E�w|���`�gL���zo��,~ ^q�R�U�F�	�G�M����~^/��sF]��%=>���{Ľ�R΋���Q�k,�C�������'�[��>�*�	�eEHϵ}k���`��o����ʯ={7�[�~���h��j��al>���޽�n�>J����S��+��@���򲻗^>�/,��8z{F��p`���5��ݜz,G�az\��5xԝ�0U%��rs�vo�,��{ۑ����ާ�=x���؆m�� ��쒯��=A��������y]�Soښ���;}���T;��]?>��M!M�m��![���$���8(��㦌͐`��?wʭЇ&�����G�ɍL�8��Aұ��3`�Ō��%�W>��ȭ�[���"���������^@���:{/^+76��o�Ӟ���MZǧ���ثb�y���=���s1�� ��������O��l�9�Mt�Z�e:-Z���G��;�`��������:�8���t�����f{�����9�(�qY	����o{���;���8�(�7ŉy�wf�u�
q��;�W�sȿ��g�ɋ�\ܻJW����M�,u�o��ݗ0��.+�6]�i�2I�g|>��7r��ܵ.���ZN�6󒜪5!�ːn�}�oGH�M�N2==�8#^ya���\����YN��0�L��z��n=qur��as�{s���:��*ŮbJh�E���G;��<��T���� ����Է�ץ{}\X^9��J,c˼`���nUp8p�x�:�x_{:�y�'~��=ξ׻�m��z�M���-�H�{c#+z�� Z���w���&����2��f撵{�7�uV�^��p��^�)�w�;εyW�6z�)���Y�ۺ�}x�^��t�[rx!�t:/��'��\�`{Ӱ��s�����c���B�&�GQ����U�J���Wv4P��_C}�A�2�����o��t�UF���;��x;�)����;�^o=������W^����}���=���W'n�=�O��ѓ����_����y<�C3��9���%��ݫ
�q��u����nF�ހ�b��f�`M��ڇ�����j|3�[TQ��0Al�n^r����I�`�c	��9EB3���eySX|3w��n��_j*�Å�j�ۄ����^��\�7���Y���+��xya�E��\p�nxL+��Ӈ�7��������׏nP�W����I�+���}��L�M75w��/ �.�4*@�=��K��$���{mi#�.�J�#|+�+�;��_�OL�,�t.'j�ve����eV��{�{rjzN���{�a�yU�O�?v?	�U���a�\0@����������qXL#�goPYYr�-����=��2q��3d�t��'g�L�P��M��M~����|���{�����f_����^?w?�a��3<P���rN��D�lbӻ��NB+�#�ٳ�'{Ȏ�����c�{K�\SIN��q�H#ݞm��G;�J���m���ގi����]ݚ&�_M�l�fJ��mpl"Ӄ2��֝��	<��{Ŭ�9���N=�h��i�l�n,�B��g�{�2v�4��u�|p�"��6<Q���F#�#�5Px&y�z���\S�VNY�����a9.;p���]Ԧ�;�й8%/�����/�@l�~��Ugy�L�����Ígk:gK�:����矯���^���}�g$����G��얍����g�^��8����tI�9��rO��������-�b������w��>~>�yRI'�s�}y�x�7:���rD�>���ׇ���%�u�yᗴ�$8����w�۾�1݁oyGN��DD�d�^Y���*�����{��o�A�\���	�G���׹�'�x�v��}���Z���������X����Mݮ\ׄ]�nX�#����@I>�{|����
������G��zoȧ�������=^���ߥϧX�b�h�~y�s�]L���E�M��z�wgd�pk�<�'�ј2��]�Gf�_B���� ����A��:&d<���p��Y��ݖ��_��F���k��oT����RQj�O��ċ�k��<�>7���8���킯>�z.��>`��W���w����Ѭ�L��0(��r��5�z0�H�<�]���{�%V����,+�Y:'n�}��n�1�'n��HN��Ȟxw�/)͸ǧ|]�f�5Аl���97B����U�J�6��������
���7h���=�I���[���}��6L�E䣲C7ݷw[�u�ދ�wM>rq�F���;;ص ���[#����C�u�1����W;�?@����zG3���S�1dW�1� n�.�w�yLZ�6���{w[�b.뚓�WԬ{7�wf��u�xt9|u�&LB�vkü;��^M݆?���uq�d�����afn��y�xg����a�}�t���k~�47�.xL�]�7�!�Bᝪ˷;���hX}ݧn�;�sTz�c^×3ҹ���k�W۽Ŏ~W�s���\�s��8&�������O\'2v1Gx�Ş[0�t��{O�#1=�Ϸ~=��	�S�ڶ������S�D[$$�w�;�<�59����v�2?$B�+Lk00�u�픮�;��y�[Fyr�BA{=�jNy݋���!8/{��%�g{2
�i���s�2w��Mŋ8ʖҳp��y�}�L�eYhg��e�4� [Z����_u&��އ=���
�q#��g|�Տ�7�;�ky�={��w��7�̽���vp�s��z��{�n�י��}�C=��N��\'���`�{���b��:�Nz��i�+�c��W�>��C�tk�=o���H���.��q����@^c>Rs)4f08!����w�|�����?OA��ǀ=5�l%726���.oޠn3����=x��Z�lW��/G,^������G|�:yxΏ�Nf���{8e�9�d���������e�,Ç�=݃�
��oޜ�D}�a��gf���K�ޯ�����N�t�/O�>Ў�ſ%[��b��J[|��;�̞��C�ef�j�e{�s�	��.�]�ŕ���l��'ګ�{So�����7#&x�n����z�f���@-�NZu*3�c<�oz��X��e�~}�xTI�<���չdɔAiI.�T����'��|�W����Sy���W���"= ��r���[RW��8�bˍ䗑��7>т]>O^�|�����ǧh~>������ύ@-"w(�������É���n������!��rn�iK{�|�o5�Xw��ïsEӗFl�?�(;�|6����ǳ}�T;y�{��a��\w9n�ߺ�z��m\9_	^��kO��;7�ĵ��z��ސ�9�������﷖@�OٸK�l�Rj��v�A�3���4�?\G1�rϡP���{���|�l��|�˾O�`��bn���P�qp��Ր�y�&�������އ�9���q��)����z�j~c�8������7���|יɜ�'�2 ;���Ó�2����͝���x�����h���5��e���$����,���х��R�?/=���z����3NU�)��Z�Fl���e�}7�ow����G��L����Af��Z��V:K�}���{��ڳp�*���h8;�V���}�{�����y�m�/�J������=����#�mIDg���-��������8I����>�>�O7aΞؓ��;�ݍh�4$}iE��	��c[����v�W+��˒�=��#��o���^�� �����tG�gU�Y3���Q:�ϰ1����X=�ݝ|ֽ�|p�=�����פ�n�Y=��p��� �.^^r^���j�w�3k�q^���E~��v���"ъ#��^z{O�Yݷc�U��}fWO����r��wA��rʅzĢ�N����M���=�QJ�>������\�	u�eĎ��ϵ��;�wm���	d�}���Xcݻl{��m���)'����-g!�2q���ӵ�X��~{���:���.��پ~��y}�"����/Vp8���H���9q[�.T�����: �ӽ�cz=ׇ��3��;ί�8/l�xVթ��\�/��{6�\teg����z@�������>�1ې��uڍ6��D�{��b�$��3���"�}��'��tǜ�����e(k�y�Y���m�{��>���(ˀ�5�|u�.&�3��գ�� ��+��Ý����\�z�{2�,��F�£�����������=ƍO��;gvU�;�֜���z�Tsw�{@p��{��3`��ǽ��������(��`�d-�U,U9mJ歱��G6��\G¹��y��-����}A#����r	���\��p'w;t�\ܖ�;g����FNzϯ����َF.�iه��~��%��̳�P�z.Ճ�N��<���V]��M����f�R9��<�f��õO�/�X�{�L�[�ww<]��w����.�y2�#��S��S{{=�v�^��2����^pz�P���y���x����bA>~<Uݿl��mP����7g[�\s�X�����Č�8�*@�s�-1��;{5����w�e����P����g�h��2���N��T�������^�s|^wZ��f�w����>�u�7=O��z3�����ċ�����>nT}Y��H�W����{�4\���W��I8�{��x�{<.�;��j׹�%>]�F��Tu��o#��I���}�"������{y�=	׺�b���t�gw�s���x��}��:ϸ�c��r\��|*g�����I꠹�.㭾�U��篎���C|�:���7^V�&��+������g���Mx�{뚠�po��ܷ��]��s<f�z��_�[����񛾒���ޭT��{Y�{�&�y�oW�2p�g�D@\��o����~�����_�
�����kO�{�����ox�<x��ǎ�<x�ӧN�?��������7A�?�H'��H�4�Ƀ��jG��~O:?=y�&et�\fT����]���n���778�fF��
Q[��=��y�AN��x�{e����Q��2k.���
ؼh�c�[
Vİ����e4�] �ô	k�Gaݰ�,�ۓr�Ą$؎�0�1{\����Q�λ%�s���S����^~=�R��T�K���("�Km�C�&N�˷R��^��Bf-�㰖ܸ^Kh�=i�p�1m�#�m-�A�e�u��n��N`�u�v���=r	���V�K�X��z�x��.֭G$�n��v7�'��'%��Ƚ����i;Ӹ�\��zœ�4t�}��ujsj1�+x���7�燍p$�ݸ�ή�nv�6�n��#��&꫓j봳�><n�&GJ�Alp��Ѵu�k���oi#�Wf�t`=u��}���,�ht눭�h@�ٕ�e�A��6 �+�	lklFqV��+-t�F���9��uϝи�}ny'9�62���XGRc(Pt�f�E�-��CE�`1���5*�Oh��o�/��I ��;#�;[ ��6jR�v-"�>���,�b�0��f�j�&
��e��.��4����	\Z5����fB�b@VW�ym�f���8�a�.�����V��il[vru�N:�Mm��r�뇄ں���{E��-͋�~���xƹ�Q���(��Q���τ�1͍`�6]M�v�!�=���s[�o��v>�%v�C�^l��n.���������n̽�"�Y�ӊ���s�<7�o!���j��`��-�j�ۍ˲��G�bx�o0lllo|
\>&3(L�AAQ���kk�GVv�( |8�v�E�\^�N�*V�� �:�n��$�΃e�)JΡ���-e�])�Z�&�'Glq2���q��]��@�����!ʅ������BWk�l�r�-�/c������呝=O��q���wk3�g'8�XV�3G["�+M�˱���[tݬ��sq�.ɛ�]�$>������`9�a-\�`������g�������+*��%۬�&�*W[��r�G�'���M�d�g��v[$Ƴ�۶x����5p�+և>�d���-�l�T����X��=����[U�ڰK۩�ܔ���
Z�E�i�͇c���єu�vxzK��<M�-��"<�\�V��.Z�OO:e۞N�%��"��7���Gl�n�ޱ��1чi��1n�9k�ܘ�ܧh��i���x(�۞gм��.���^�܏0ƶQ2�2b��-+���qT�k�hL��9�k��k!V�0̹*���l9{"�˂Rˎ�W^����iM�)�3�6\���6jS�_0��`��e�Q���5��t���Ҹ��Ե�H���tc��W���#+l \�1���5X�%R]-����a�Mm�Ũ��[��ڂ�宭�b�jX%�"lW���l��n�N#mÎ�1�f�{��_{���u,]vJ�m�#��t��d&FYb,ݮ�����W7.nG��.&h��B�bYt`�lj�X\��Uʚ獗%#/:���l7S�����9��>�7[�T�f�;c��:��ZnNt��F�qcj&�6̮��`�e 7�&��B�֎��n����ͳ�b662�8֮1�ڸ�u���d����0���㩸��b6���V�;r��s����z�� GJ����x�X��E��c�pt�97����I�뫾6��`��e�+���v�b2q^�'����.�knp�]���a��)��m;V�tL�5�,bk4&���.���GB�Y��K#3��t��l�s�Ӭ����4ٶF��Tn�k�M(X@���1Յ�֯tQ��9;H����i�1rQЍ�3J�\�;撺V$V��h�m��pv�s�WB\�Aۮ�a�\�p�E9���5efp���2��cQ�Z�۝�8�;uS�@{�\ura��G*^z۰*8�v�4�%�X�`P��
@+R������l�! ���KL��P+��� 6^����M�۬x��^�9+Ǯ���9cyz���i�yM[�b�@�J�1���!m%�S��eAq��^���݃�[0d����ڶx`���жs���2)4Sh��R�"�b�S=�+��m�1���lk�=�g�y藜QQ�4��a�RYF�Ȍ>�nm�4Gv�k[
�p�AҀ�`Es)���h�lK0���{J`�RhąxWfʪ^Sg==�ܖ��1�ŭ�j6&�]��8�h=��q������ٯ��&]5��z��YZ�X�8��D�~�����m,d�:��S�,5��e�]P[hiz��,:����H�!78��Q�cjh��WSXk@N��4*�9��5��z�'��+�88x�xڌsƥ���Z0A��,�)�lp���E�R�UX�̸�k�b�X:����@[bhuF7g�n3%�U��w^��B�RM(9����y���ɺ��[�V��[��qLOd�<R5�c#q�����=���-s7	�G�R�� ��b=�M��5�6���;���sX:�\0
=3�,Nw;L��kOOE��2���舏YK,,��	5]&�6���f��ָ)�{�:L��<���S�]���(�J��]�v�$�=�h����t[^���q�y�r�]Z��B���oRjQ�V�K����s�2a<�� r9ݎ��Iu�ˊm�l����`F-�<k$��{6��u�졷]S�]�'o[�Z_'%3ۦ�n�p�Y���b��o;������9�.oi�[��j���t����+��l��]s�Mv�RYR�,CL1]�V#������W+0mkFvɼ�!<��q=�Őg�IOb�@�H������([B�W0���L�Z��X2�hʛ-��E���.�8�Ǔ�m�v��+v���]���$��'�՞�m����������^2�8x�9�$c�f{qYs]B�;y�ȉ��5�'�*��hib��	�@Kif�j�ю�`�6l�R5�����s�#�kg�k+���^@3�?tc�{*�?w���Y��s�ŇhŢ��J�ľ5��A��������%7�����c�pl�K]<���ꖌ�hcBռ�@+�R*u�.��e�r�Z�d|�_ͪiX�k4��݉��;qyҦ`� ڼ�٨K�e��dk�.`bmînɬe	����	RiE�뛎���wa�"0çZ9�0<����m�Wlm��-q�����	Z��� cL�3j����ۆ��r�����^i�ؗ�v\t���f�u���Zq��y0�r�S%�(�I�����Y����b�M.��Ꝺa��Y�<v���q$\�-�IM*h8��Vhe�CFb1�Ҷ��\�[Br���<<��N3(�B�[c�5,���{�9��!P��+���I�Im�l�,�0ƺ�&��Y�&:ވ�:3��#�۴��T�n֗��m��PpfmCMv�8����Iv#�I�8�X͐pu���f��J�jA�Fnݜp���qb;-��`S�&��^�	ny^�����T�u��\g�7^q���GP'Yzy<��t���\nݎ�Z��p�9m����E\����d ��a
�ir���N��l���x��7�:3���ڱ���"��q���qH8�{
�ƴ�����n�����S��&�D�{鋱����Ieg[��l�/��/\\޲�����E)	qL;E�2�M�4�Չ�(F��ݦ��"i��&]����d��38KHh�P��B=�RYvn;XnV�����N9.�.�v�,���9��8�HV����eĆy��tpm��.�{)�X��q��a˲ͻ=�zC�<u�tm�k��չ����g}-�e��:�]��=�5���ع��f��6���&����{���\l�v�Ԕt�&��Έ7�����W.vvۭ\�dA�Ȅc�� ��a�Kݹv�x����g��+hˌ/�=-���q`& 4A͚�������6�p�q�:��yy3x�Kf�;�m˃H����K�%m�+��5p�c����VK9`�a��)���L�6�F�(p�bh��&4.�d����Q���k��Ѵ$v���QK���l1M@k(�s����T�-y�%�b�e^�f�Hڙ^ێӳ�z�ջ`�&���
.O=�Yt��7����k����'`YA�Q�.=nh`��{n�Ԝu�$��1�z	LR`�3�����B��$���f�r�l��"�ԔS��g�3t�ɱ.�V�7��]���kУ3]z��Ls5��^<%�0���x���!�]��q����]e����˥a�E�������v1�ci]�|��i'>,
:�,�l�gN�Z�NR�>b���iظ������{L�`�tp`y�{u�δ�s�����T�R�0%&��F�3��*�Άy��V7��]vh�oZ�떭n�Ӧ�j�����U����������ꯪ�����������������Wc'��m<n��óGI�.6�L�r�kI�\@��K��f��V����[�bt�(�[��ʏQoOJ]8�&2��`�=U�5�h�:�qI�sL�r��3j�\�|��x>_�����f��@����'�8��屆�cX��$��cZ�*�������/K�-A&ݬ2�y��eI�S��E��l��CmI-�:D�3%���j�l6f�t�Gm�����;����ol��ݔ��gv۫Ⓥ+�^QNGpIכ��q�{ڜQg9�V�eeAEY��	��GvW߳��m��u�����9�i�u�����i��։�k��PtgdSn���L�γ�}n�8��γ"ڵlܶ�չ%"�����R���.B���pt}��	�ڳ���p��(��+j3���/9�gc�MvQqGm۠��v݉��Ir������Nzo�Z'���e���eY�o�Xp��n����w$����:��.G.�!,�m�}�Ol�HYvm۸������'gnW껻�q�{�a}��}△���[��l��ꇟn�/$�T\�unl\ ֳ��^���x N�MF���q7n-\����c���;�x��D<�Ƌn����z�v�,�5��a
J#�ˈe�][�n�N�ζz�M�����]ν���h�g6��)�.��f���z��$۪�l������0	�]��K,�,ƂT�R�v��{b%Ё���P����}�]�<%���4,�ͅђ�dF����s��F�Gvژ6�J�j.!mԆ��T8Y��)�j`a3��q��aUx��떺pV��ˊ7��79�L���T��c�}xT��e���YH:���
t�%��;v�	�ɶ����V��a�A��lN��	4�7��v���:i͟LvPқ=���OV;z�(:���a�q^�m�ܼ����vG%6�Nh͌��4��#qt�-���+ �Ur�l=m��XnO9^(�Y1nW�����F6ی�_`�cQ�+u=y�w�ϴķ$�c��*����[��ݓ����c0��K�a]!HjS���,��*��ul�Mp�h%�V%�%�^{q���d�8Żu��*)��0KxY������]p�f뒫����'b��m�6��J%�i�2X7 �6۱�E�r�"�*Ɩۛļ�����'Y���,�5��[��6�)�8�h���8:��]���5��lQ� rӎA'�N���u����6l�ٔ���6�����n��\�y{>qм�*�o1�t��E޽g�����6�����NrW����w��qۢ�c%�֋6�Shћ=r��X�u/$�%Y�hXF����<�rә�v�v��!P��eu�����[M�u�J�u͆�Z������*vZ�^��&�8�۲�2íy���ԓ����������Ұ�!j�h�4�N��b�NcYj�Ġ�B�[�`4��	lH�FYTY�T"�Q�[�R�cA�"Q`��(Pic���0R�#e:�Yl1i �IYemZ�YIhX	-��H��T:��RYZ�R��cF�o1FXF�DJEcVV3�į���Z4��kf�L�B˘h�Z�o�`�x�.��ŋH�V$�%>���g�Ӟ�.�iq��"q�ګ�O��8k6r���Ql_`[݉�jJ�^� ]�o(̍s�!����Z|���j-J��tg6��"�h!@:�Q�KS�v|����I2צH�ԭ���wI��*rr�\�Ò�k}�eۤ�p�	K�A׳��&̟_�t�o�ql�'4E�6Ve���J\cl4l�����ۥn���]���wo���(4f��EhB<�fd��ڗڹZ������@� R*�Ϙ�Rv`�ӵ�H�Ke�gX���r�{-F0C�v�b!�=z�,��ؼ��8��JE$�r���ݦ�s�KN��N���,
 e��H���"��~tm�{�.���>����)�ۤV���\-Z?h{����WyS�Fn�QP7[�h�MVE!�T����}͇j`�̱�#j� ���m���7��X�e���K�J#U�ƵVj����_Zm>���&��ͷc~�/yi��h�J�����g�e��Bڬ�Í���p�R��õ��MWs��)�@z8��jJKO�3Ng��'�T�a���L\E�W�9�+a��e��O��8d���%55k^��T�9}��Y�T�����ev�B�Bm�M�&�=ʎM��y��<G:(�I��g��3-ՙa�N.��~ژ۩[��S�mk�%v����8	��2)�$��'� =�9�u��Y-Wu��*|[|�ğ�c�	}�V���HH	�p�/Z|8��ڑf�Jq��*���7P��owk�e�Ǳ��)yR��~��8�4$^��{7��s���*�B��|��:�Ap�`u=.���	ّB�w흓�N���7�}���>��ሠI���8�4�T6��+��q�R!�JY�O;u+c1Ѻ�F|��i|Ƨ�p�n�}X���$BZ�qVX0���Xne^���KU�bl�i�G�����R�%I�����E���N���9I�L[`�ݛq�c.���h�u��@1w����gޭ)'H�<H��;����x���N:7K���J��M�I:E**�u��e��,�vfb�"����}��یȳu�Xu5����'w�����
֣!�������I�B���v��+%�]jl�Ӿz>ğ�"DO�.&�>�f�NZ���"�8�&!�EnN֜��K^[�N������b��曾�wf��.��K;�2�P؋�+ުi�Q�&��U�[����;14�ȫA�Z捱�� �h!HR����x���N�%�^h� ]��N�Ro:H����'^3T+*J�۪ͧ��̋7Z��G�'(iW����?dz &��ͯ��{��y5��/g�.���^�b�s9�R��hv�Л$+�����Mҟ�I�+u�v�Z�֦�M:+�Cgi�̇�D�@>`7q�H��JB[�T�f�❸�m��vv�_Bˬ�7�����L��1��F[\ٗ��{5�ͻ�H�ُ��7%�Jҕڧ����̋7Z=h�"N<�@2`�'h�9��� ,>I8���[��֮�6biڂ��,�R�͙b,��7�w�>�)'�c� ��a"*�+��Ǘв�/�P�؈I*>_\���(�'V�S�N>�J��d�h��/gy�}��{F�uh������;2 |I��|Ԡ'�>��cJ�̻mv�2i�-���wm &XE�h�R��-ev�.ŶE������r��5GF�\u���8�{#�`�%��	�iM������<���'3i�РYr��ѡ.X	�au�\�K�5燭�g�3tv���d�A�*Wf�h����<a�.0¶�Ck3f�&�ab�����i0]I�+�i�%{i�����h��B��@"���:7�Y�i�i�αq�Y����j����XcS�\*ݵ�Y��n��u�M/V٘Çfp�b�"�ʊ�f�ݟ��mY�OwU9s�n����̲_�SY $A�O�#� 12f8H� bȝ�3�Y-j�`�M;P}�8JS���
wb��Y���˯8��j���}�3*��J�����u����>"!$��;sp����<�}�K7k"�b�#�{rό8ɔ�_�H�����i�y'�I8o$�+Nځw�\��e�7�j�n�ݬj�`�M'��Q ���H�)�r�P���Y���k,���Yu�!�k6���7���;�/Y�E=-�8�I"�&�*d�}��o�w�7����y}wYxoD>VN	[��.��ԁ�吒�%N��y�/5�D5�kN�je�l����g�s���9W��U|�9�LR�y%�~YOoB�����~����s�����}�,�����X~9�98wH{�K7k"�b�#�n}�,���b��fx@�/�����dy$�����9�:�Õ��ԭV��i�
��!#��䞕S���,���J}q��ȉ�[3�f_���7��^��K�^��31���	'�I�Տn���Run�d�Q�����	$|�$���3��w��B��nA-]j����k��7,��:��@��� �1���}���Y���q3���km�\֌�hW->�A�#u�,�$����x�/�b4�mǷq��b!�i��wp��7u����q�[�E;�jә>;��M��Y��|����ڌ�-����o/ozW�p�f�z>d�5Sy���*)5�Ŝ9�xk�O����Ss��҄8�|z����Q�������`���/��d�I�����J����N�Q� �k��nUk(�f`�y��}�}wo3���ih�sZ31�@z>.�:"��g�$����I;0sR��[3" �r�����cDڬ�݂�W��{�����Ҳk~z����u*R �O����-c ��5:��u�`�D2�ɻ��/�-L��8��y[�t�;y��/I�P�FT]�싴���I86aVV��m[��j}ԴM��l�h^�D>��w�]�f��D���z�<���f줝&�g:�c]��kf��-j��Yك���R>Ig��"'if� �s T}���q��y�'�k/1lا����}��Ջ����	�=�;h��$3��vw��籎԰�.z��T�����[�|��K�����.�0��:QY�\���(,�U��B���)?�T����a��^��,��K��,9��;u%�)ϭg#�������v���K2(hA�tՄ��f&K�n=e,i�8�����1b^�8&ȭ!$��DM1���'&M����A񬘗PK�ѝt�I?���nhܙƇ|Gۯ�h�Yy�f�<m�>: R>IA�f` fS`1Ϝ�*#�|�K_2��f\K�K��,9��I�Dy$��cVq�p��>��	&����s�%*��}
1�;V\�B��,,/���k�1���1�.υݸK`�}NV�so�O����-���T�GԈI8	G���Չ���we�-��S\��A����n9�YoXFV�ɗ����>����ߍ��3����|�!�w�]��b .��Dl��W��%;u�O��
}!޼��Q�ȶ�ʍ'�.]�n1�&��k�H8ljR�h]k�\뮹�[��½n�;lѬ�;M�V��`��������5A�'Z�c-�5��ñ�����q��Wֻgn����n1���ܕ�<n�!n4aʰ��zP������%��w�]�mrn���n��U�<Z�[��m=#��E��<#���k�F��M�OXJ�jK�����].�1.��G ���nw99����U�b�c��L�1�P@�+��؟��r����ͧ���7s���|�ae���+�b�$$|�p�;�{F�o��R}�6+u�v^&���܃�%J��}
1��p�^�k��hk�Tˁ~Z�ZEݸ	%��)eW�`1U1v���3-��$E#䓀�o%f�Z�ga܍��*#է�'�����.V�7�<�ܻ��R�ȤI8	))QT�O�9Y1�jƫ��۳�pr$�Yxs@Q��D$|��;�e����%������J�$R�X\ll(��][u��\(��F�s�%6H`X�,\�n����>����v�m�S��[�S�nͳ��&�~en?�)y$����	uE�6nhi�i�Ml��F�d�<G��K�<��zO'���|��OL���d9�����te���U؝:j5:^ެK!��ʲ��>�Q�5�'+g^'7ḘXo7����'v���
Dd���0Y���%>�y6k��n�U�k1���S�pvd�Yxs|�\E#䓁@'�*�K3��-�p��=��D<^�ZĶ�<ne� hH������66�"
q��G����"�8"LџB��I��Z��4o�Ț"��UU�K�gd�:��/*O��D������G]q��+�{`1����ֵ�e9�p�9U坲��\��TG����l���-.�^c�m��;f@Y��*��>F*3X�=�iF��
��ڋ�Km��s-�N��O^`�|�+jՕt�6�G�iy�!(����4��]�z�����ƞ<x��ǎ<zǯ^�m��z>���{X������Y����`=�Q�`~s�	�W��OYcz���&%6y_D���zm���}�늀8	���Id�v�A�^���"M�!�9s�����m��j;�:o;��7O�L��g����9���|^{�y��#i+���gѻ>����_����[�ry:�����J$�o?=��>�w�}ޏ4�tw�^4M�����&.��D��������/m���1ϧ+�6��3�L�D����{ q�3�u���_����i�g�� �E���]�Er2苒�%Vz{�<jj[|8�3g��� ��+�2��$�xUF�&q��ksryo�~�`ݓ�E{�?e�qso��=���#G�puV���Api�}�_�m6L�Fv<��ܕ��Ӭ���rv6[�������ý��t'����������'�����/��<�R���)��w��J+�G{jE��w��`�S���yo�g�0�j͙�r{/ �_^^�<��C�zW.���hJf�]�yU㴎�l'y�%C{z��9<|w����:���L[�>�����
����O���}�ڇ�������
����^~��[Z��GR��S��&����v�� ��&罍�O۫;ᝋd�W���ʼeTTZ5�/f�h��^1m�B+@�-�w[J	���x��;�##��Y3���C�u�r̞� ;v�.���'��<�w����Qr�������\��C��3���ť�]�d��\�7~����\׮'$��r'E%�9�_5�(���{ٶ�m����i�|���;�����,����=�\��nN[u�۬���8����m�N+7$�d�Q�tt�-n�59-�ܠ��v��\GY��]�R�n�N�2r �/�{X��${v��/[�����(�r��O�ol�ݖ��'N�p9'\X�-2�N)6�v9Թ�n;���#��FM�D'��PI��vY&��~�;�n���Yr=k6��m��M��M����ͷq�q���#��ܺm�l.�e���m�I}� ���� ���Cn�gW�ӣ�Ĳ�:�mEa����";2(�$�9��q�_n�=��IܳY��V�rN+��tu�Y�ҌҤs�(��h�lڄ�����\Exۤ�+;ml���"���פQ�~��vR�߷{�9g�s�\Mr�y����4a���|���!ڼ�;��x��?�omV^S�Q����
\8f��$}X[:w���K����y��������r;��d��Zs��*�IϪ�h̭B2�a�E���=W��1#NF�J�g+�\'����;���7�-�}�,�e6fX���Qw��=���)&PA��i ��lby�<���N:���Z�h�u��w����������E���$^3�[���k���O7��w36�z��P��`ީz�Cs��`�,�ƒe�BfQn�Hx^�Ͻ����^��O��ݳ��4L�Yy��m��<���]�y����n	l��P��̯Bg(�M�˙�Y�v�y�i�1k�_<L�We�(�̷������v�N0I�̓��"<�"m��'�.�0oV������]j/���⫖�O�4a¼y��w��,;��&03ț����њ�;�̉��}�y����ħ�o���O�#j��ra�je1����+$�j�R�|�;���l!�Xfx�m����l33��`���v
���f�>��3�eһ�v������{i��4\7�|4fC�w.�����4��~%�[V�l���r�����e4m�M��}����/��``��p�0>Jz3��Uw+���|�~j=����W�lf����->�����d�����mq"�c���`���"�}��u\����xΗf�+u憷>���v����)V���u[dg�U2�Id3-�{�:���^�漥�Am�˳8&],�݃��Ͳ|���2E��H�`�pEo33�]0�dS��ǛQ2N�W�U���-��d'7E�K�}��}�=��}-���"E���"�$��2D���c�Ɔ�^7�;��p��嗜y��`Ԝ;��D0`p��F��kh�{N�8Ukk��&f����Dbȣ6.Ŵ��I�6ǩx6����k�z�ӽ/�(\��2\���@~�&X��i���X^�.ã�@��: M�]�FOe�܍�{m��� �l:� M�P����f�a���D�lM�HR\hY�ô��(�a�jiK<U�;vx������vX�on�q�ܥ�yb��&�c�BYt0�	D�7F$�;Y���E	Ku�˄#7Wq���-�m���Ieҍ�����b��%sv���G������G8���������O��^���A�]��m�W�L���u�p�lƲ��X����$���0�>�'䏞f����q�a,��=gn��ζ,�>�O�k��2G�$0`���w�ǯ����e:'��@p��x�2���.'�[�z/�0l��jN�G�2峷c�)�;�<ݷֳ��BO�VB;ݸɔ>L�7�T�]��Ԯ{F56�B��x��u8��i��|����4f칽�iow�h8�oz������h�闺,��oL�����z�=U�O\����xK/7`�`Ͳ\7�ޠ皛/�"7���av�X\g�Va�x�vC����
�;ո��߭ɦv��ǚ1�8�˾ɮ����Yq����a��)��N=�]:�8$~���_�>{Y���щf�[a�ӸE;��m��qs���qq2�R���G�-��N!'��s�H�`̑�����.���Oy�7a6���:���֑,-ÆH�`�'�v	;��@],�h��.���c�R��"�u�emf�n8}�Nk{4-}�{�"�4��8g�+�[̼8s�UK����}�/pEKaXa�8���0�>��d{gs�S4�Wy��$�`�����"t7W6�U���'/��W{wMn��ot\��$7�O����9s��2�C���[wQ�e�w���>�4�c	�����YUdjo�w��r�/�̸���}�,���{��Ye����M�w���S��'�0h������������|B9e��2����e�>��w�a�wV=��f[Od���0��n��y�K�mO�d��fH�� �-�������K��er�ZE�.`��M딷%��]�����kvlJ��M�y��u��4�_����n@p����˝��qZ�\f�0��3Ѭ����Ȃ�'�?����K$\0`��v[2��m��}-h�o�f���N�=��ya��d��N�f`�o�o���gܬ�����7ӎ���3{�[fYp̲����w�s�+�=�j��9�;4Xk�.ny�WR-��$�L:w*�4��y�׷���wC_�t|�y�.���#�Z.��������QE������5����a+�݃�yV�Ss2����d3*ȝ��P����(c�;e���8q輻̝��q\�\gz3�p���v�t[�퇫����n����V�̫!�l&a�F��M����ծN���-�{,�v�N���B{�,��Z[3(�2Ӟ�]��00����7��B �\�<@|���1������
PN�.���Wh�ݕi ?����x��M�1���N|�#����w8�0��v��>`-�����3�'_��e�3$\��� ��$C�<|)g��ޥ5�\�=��p�o�p�/��'au�Ur�|�Fsߘ��2�imdC+���5��xxw�;-����+^�(����d.��q�⟪�E�Nݛ�y�3\��̲��\&e��S.�L�����!hݢ1�z%���2�0�%�Um��;�z�J�w������� ���ԤuL�.�N�z�551q����`��d���]�݅N�`a�<�{�7���t\NOnz`�J۫gk�9���3|y
��(�~�����7�~$$�K�H����p�>	�7b~�b�����;'�u�Mr�|�����m��`Ԝ8`���Dy�O���ǖ��4"8��q���:�xsn�9��Y���5�]p��[1+�$��Ӈε�H�Y"�'4�ܭ�g��y���¥f��hfMk_.�LU�v� $D��E�8`�d8oc��O]�Ó��o��n�����jU�v����!�˰ojp \L�~̧���wc��!&�3,��Afe�sD��9����T�����Ο0���`�$;�e�̌n����Y�����_{��Ϯ�Rs���Ni���-v^k4�y[��+���7�=���1!�6C�l�.�	C�d�v�4���[ْ��}��<�����ܹ�j�v���yZ!ܦ�fU�$̥��$����&����'�TYM̪����f����=-N�'�^�c�cuRj�7��{J.���i�<�ͱ��o�E��-f\rw�= �s(�3��">�� �*H��"j�����.�Z��dG�낞�8т�ܚ�x:ns�^��q��/F��X�,+nBk�5�c���8�͹��́t��n\ȕh�A��sn&�[�j8f�A���`*o����Wh�W=�ӌ����y��˥D��VѺ�:=�8�#�����-Z�hF�bs�Xe��+C&u�2���{n]7l��Y;]���$�,�k�bK���ߏ~?=��rQ�&Ř�t-	���YS��l����a�q�x����#?����!���I��d��g'뻩�Yq�������O-�)��oKm�^�x6ˉ�Q�,��o�M��p�盺�<����xb{I��޶y[vo4<0E���9�����vV��������#|�3;�����{�V�c�+�S�:��:���N^v���`���vH��"�E�xsɡ+�[��Gf������!���Ngo39t]�G*ˌ�F�6]��{Y'��j�/U�a��y�m��a�H�	8	3)��u�s���󷄬�޶y]vo8>�ф?�$C�D8`�I�U�,����{ԶZK���@��D�&�	Kq�m��yQ���Kv��^����~ߧ����O|��=���3��������g��U����=� l�a�.��z�,��m���9�M�fU�32��c�6�e�5TFq�+�1�+��iT���0��o�5{|�>��Hu⊈#�g�M,�(A
�~8��A��4V�W�C/r�g'��(��肀~��0���7��/��wu�.3}G6Y��8>pBG�/jմ8�A�������p��d���H���Z�ms5��[K-��]�������0`�����N'�!������hnh�bD[g��zƂD'���1l��]��Xk���Yy��oT�o
W(�s]>�6��ͅ0`�gԈ�H�'#�j'�k=�����E�������N\gz0��E�{���ot�����w�g9��{�����Ox�p-F���0Ƀ����j�-���0$ЅMfU �\�?w��{|e�����O�3$@p"sA��޶z���������ƛ����3t�b�ö���O~i����k���q���fEmh�0��?��o��5�]ŭB���<0>5&C�m�r����ћ:J����G��d!�Yf52��̴��>����c�v�?�����ok��Rﮒ}��5z�����%����3�˸���i[g{s�����3V�|��&#�?�gو}�DE@c���{������3\�Q�msth��3-.��3-�fP��$�muÓ.�P{M����V?�����2Fg����M^���z��h�5���_�v�{8M��
h����`"� ��o��p���C�+�}��b�ގ��R�-J��}<��-R_�S�H�y"dj�i�B|��'N���4[�x�b�1���v�ԆCJ̫�\�b�0O+y���p]�����ͥ�uO�qFw�9�WL:����s&Ӈa��=(vR]��7�
�v��4Κ�;j!������k���M_+���m�Ӎ�v��>�\{_w3�u0�i	�Qp̠����X޼����w�Ԧ+yS`�+/9�0x0mO�E��.$}oV�7����*Dh`ݮ�m�����s3iu�Q�6�;ќ�,��xG���������kZFL�(��u��{ڷ�^HjX1��廒y/[<|��|����Ĳ�y!�}�	�yg�}DdT�PFD�Tc�h���]��m��հ�k{�,3��0���W׵3y-�E{���F�w�vƧr��C���ɏ40�C�����n
�fZ���ov�p��/<f6nqc[[f�S ���p�h�v�(۲� ���Ͼ��+B =c�?�$|�$�y���/Yʛ���������>���bŭ��`�N#�t���	��8��֡	��l����f;������3�s3iu�Q�Q�����C�`��`���l�m�n{���U�f�]��u\�i��-����4���@�SF�G}U��컶z�˷��/v�!8p"p� 7��&'��Z�v�8l�:�y������ݗ��L�)Yyϧ�Rc����jo�<�F���uv�g�!9�z��(����ᳳlt�H�,��`�Uʼ�K�������ιGӜ��fQ�߶�{�>4���Ǐ�:x����<x���׏��ǯ��:z�x��yW�o��q�uR�5�qPgm����3���׏̆�7FhG:/{��;����@．���g��b�fY�甉�3ހ!��XO�Jg��a۳�o��������������>@�_e���q�7e+��ݮ9�v_�.� ��'�nqF��{�e����vO9I��0�9���;���b���Y���Ǿu�Y��ݷ�<{/��\�w��<�5��xqzZ�oU?D7����/���x�쇸�;����6��9��oz�����=ڱ����6���e�`׏� ��ݏ���/�װ��2�����z5����e4�����;���f�.!��o۪{���\����f��;8Θ$��@����y#V�Jvn4n�;��%z��7o�Ip��k}'���>�#D`�%�g{�i�K�޲;�7Mn�/Y�� j��[��x�1�P:�k�A��:�]^��Lo,���(�k�T���(\M��q�Gc"���\O�w+���xL� �p���{��Y`���Uo�}�!϶�"r�����S�a\��1����}yjey���{�9�5�ϻ=�n�d���>R���<����Y�ӎ�a��L��%�K3z�g_^!�& 3ܫ�<���~)�{LnÝ����g�Xǁ���x��x��J�f�qԼ��������j��u��A�iD�w�#%�H���s+%2*�gY0�WYv>�W���E��j�s y�wk�ƵR��椒���&;���}J��:��ѻ��|9|�%e	J��Q��n<�(����y]��,��1�|����Ĥ���0�az�?�h8Y'	9���ZBf�-�f�>�L<a`�R�q�#&1�&f��L� b�{ݟ�X2�y�-�B���!l�^�n��nY���v�L��<%�1�^�KzRF�!��R�,�kĻ�,��V���,�m�y��;����W�^]�N]����,�γ�m��0i`B������������z����n�mY��3"��KY�n�kh��m�I6�J6���{W��k�.5�#���=�n?7�e6(�����q�Ư�������LBΌ�ƽl���]c+(Zō�۵��-m�������闩
{��}�_'�����oD�048�v�VZ[mi/vG��z�o2��bam�ζ[��V��[��k>ݾ��_]�/|�ޓ�#S�������Q6�0���(4��/[i��z׊��ru���g<ӧ)7N�����=���+[��Um�0�Zt�������e��Hַ6�"����1;�z};睄8�ݓ�M�=�Y�6֑�ۓv�q����wQ[޽-�F��9^bL��^~����R�����M���$�\�����.�^^i�[k:�;��;����¾kE��|�t(&�YkK-�Ie���׎�w�ޟ�t����\[:�n�߸O���>ܰ<d8�5j�yΔ��q��C<y�ZE��.I�"��'K����7A=)��U3r2��X�eq��v�v�n��0鐯v���u�<��n�"��D��6a��MKO	u�RƐ�[;=��N�H�W*�'"� ��e{1�U�-��-�PtK<g��K���Lph���������.�v��v����F��7������0��T�M �suA���0�J,�A�kv���+Fp@ymWf��N�#F��s�;;uHE�#ضp�9�����V��v��yq������0V�v.sv
x�Jz�76zI�6��v6l&�ؘ�c3M�ץ���[�l��6��q�s���v�H��ϗ�����K���TL��m�xѱ�qP�%;��K�7X�6Sۉu�;�sc�������i3A�Z8�q�p�%�ӟ,�s��67&�oEk[&A�z����6����m�ؐFi��Y��曘�n�@b4\.tM��e$9s��r&v�!/�d:�A����V{AۜŎJ�:��y���CO��g�mҖY8^��͉����6�a�i\x���ŷv�����4,��p�A��]�k�j�<�� �̖;S�J�ZE]�k��K��-hY4Dׇ,��n٧	�1�t25Jd+�� W=��O;�K�u���w�j_P�m|�Ítt3j{���q'utj+�aH-4l�\�c�nu�Q�Q�Q훣M��hc�N�C,��@܏���8���r��Mvv��6�gksRq��Z5#�ح.��x��!�m�%6�̽��)f�g��}O��K�bz_9�#M�Lz�M���)���Y����L�i��Kv��࡬�K6�4�X�Mp�2�f	��*��ޚ�u��a��������:ƞ��e�?Y�}����x��	Vh��/��V�~b��Ȃ��"�B"� �")"�"��� }��e詣F���ˊU4fк������d��0cf��K1f%�iN2Gk��"�8�8�U�V�M;���3�vM/�����VX&h8np�91bfh=�q���1�6<�cpjMf5�5���R�3��9�c>��� ����<8
�������ʂ[==u���g���ی:Y�R�	ӵ`�s֔ݦMZٍP4�iJ�S������Wm,�-n���us��xqj���(�Gk@B�����}��z!%�>q�p";�k��Ujc���l�=��8D�xnaYW}ϥ"�õ"��8�����[*z��x����av�0���&r��Mg]2�,�:x0l�U��O�d�B����O1�<������WN��!�.fQa�I�-̣�3�]T�j��Z|�Fs�0���	K��)?�����5G�9n]���ߊ�5ىm�7��v�S���DA���!��U�b�g�+�l�0d�?�$����>ѡ^>�u�����&����,�:y��O�H�v�0���{L.��k�Ǉv.�/ټp�$��gv*[:�C!p��0��U	���.�ѣ��:}�DO�"��'�S��T�j��Z|�Fs�<l8��.���0on8��Kf������7����:S�3���qp��x�k���`vS�ݽ�վ��ܷu���S���������y�f�p������y�'�J����H�ȢH�H�UT]�E�s�]'p�`�*Ȁ� ��)"��"�2(���'�VB�^g��f}�l�=Yo�O7�H0kN2G�a�F��n^�k����p��$�����{vn�W��Rk��
R�㧘0j��ՎF|��"�����i����=^�E��2��8���8`��p�jssj�MQ��O���k���o��жd�]Q��'�*��X0r�2��d!��Y�2���3{�~�޻g���9���`��Hp�������y'��%��9�v�]��\�00�!��`��:��V��2fL*ej33.��5nm1K�}�?~�wI��%/�	?�L���޺G���9�u�y�n��]D;���˹}�3�#���e�̑v	>�̫�֣^��C|ʈv����S��T����Z|�Fw�����Ne�Cܧ����ћ�mc�t�3��'9M�v�B$̭i�>s~o���rO
��R�W�$c�z��T�ej>F�{��W���:2= ��1�U_%ᝪ��F��M�č.σ%?���'U%]Tu9]u
�H�B �*� $H�]wEwGQwrPuܥwI�NWQԧu�wqwG�oWׄ��۶��쳚O��Hv5?�'�$�p�	wN��1��P��0l��0�#���5�v�.*���|��)���we}�ד�p�d�������դ}�0��e�k2���d���98xS���{�K���V'��g8�7�!�	8	K��q�Z��rfvI�G`�q�úL��!���H���\�&Hh�B	�R����y[�	��	$3��̫�fW���{o��w,懓�l�.�8��7��U�<9�w�<��E�3E���0/��E�ٳ�Gϖ�p&s�mgZnJ����/�b>��@��s��/ŏ"|�����	쑏7��?�C��榋s�y�Eǚ�e)��5M������0d�8`����8	緎���n��1�/�ޯk�d��i;�ˬ�L�Y���'ޯ7���ށ��&���f�єՙ0�I��#��+A���Y��غ��Ԗ�.,��$����ǖ���p,�Ȣ^��DT94�X�gR�A����qq�]Ru��u�]q]%wEwԝEW�']Ċ�`� ! "!���"� H��ę�����g�$D Џ��8p�����3V��G!�f[<����5�͎���2R�㧃z��s-��V�L�]{~s�(�߸�Im���knjH����Լ֫lQ�v��<@�b\�iw_��N!����-8��V.��YK�Uq�Q���q�p�a�mn�!ܲἶ�f[d�ވ@��:oZJ5r����>�x�c�V@W.&�;��*f��8L�{d�5��������B��#.0k� p��"�7��z+�I�a6�3��&���hʵ|��Za��ڸD��3*ؐ��Wm���F��\�F���ݤ8`�3+->u.xUƱFp�_���F0���������m�aO2�q�u��$ݑ�����$@�:�>���Sq�Y����5u����l�0x0`�$8`ڜ?��v
�x�0���vOvF4�mK�}�bV��\�M�k��I^f,�P�Qq"p����ͺ��w.��x���C����<��i}�b!����O,SZ��~�uU.\e܄�U��������U��Nut\�u�E�S�tu�q\�Eu	��T�Tww%��u�[�d���>���1Ɋ�v1Ѝ8�A�6�v.�6���ře�y�4P�]�n*�cdD���&�֢��L��VT&̛��q`�6�ba��#�^��S��#�y
�ۆ"��ۣhr��g ݔy^�(��W���0ˍs���}���i��D�u�
Sl$pn����e�E��%bX�f��d������r??߽���߄��:��k�*<�i��@9ֺ)�WgC@��UZ�����8o7"��Ec��8IǞg�_L�mZnX�8���9�X�<j-����m�}V@!3*�Z2��Fb!�o���ǓX�ַ}ZBn����v+e�K��X�;�q�^z��髮�EHj���;e$٥��"E �G�$@��$���k-��i�r�q����l�Px0f�!�����'"f[d�k}�9|�k��e	���	�w~av}U�m=خ�F,W�����.��lk;Nos��=~�\0f�_<E��j�tXBݗ3)=,򲷳Xoi2>r�v�<%ƱFw��Ϙ���q��Eۇ�z�Ǻ]��(3h@�X0`j<�;lKKX�W��U��1!�v"��d�]��0'm/R�5+\|~̡�3�a�ݷ3)��I��iB�+x�L���Ny����c��*IŃ?C�w�L�9R�{ c���o/_u��ތ�u�r��٘*�2^��ZV1��9���`���?��ooJ�����a����z��qyj�A�>�S$���Q+"6�|i�@������7�� ��H H�F*H%��]�uEGWt�uH0# �D�F��e��[g�s���j��ֱ^pO7�K�a��^����VF�v=�����̸��^>����?�Z��IǮ1U��\Ջ\���,�|�̣�֌����̫"w4n�K̓��FR}�i����4م��;e�w����)�{�`�$;xQ���M�2�+f���[	�YvљF��EͰ�p.ύ����64���-ǝNwA���|���y�O�%���vH��"���?��De#����# �M X�!�����&��T�q�b��\��^��i�������o��1�)�$C�;.����+gz/��<�=C7��rp�;ǒ ��̑v�Dy�)vU9b��(��]����w=��37\/;���nr���jp�d��<q�4s�aRI
9��\����sF���?�f8�y�^��Mm�"p2��=Օ!--��1'���ݫ�1r�}�`���,����;8W�|b!��d�]��S�,�.���a��M��� >a���t]tU]����TP	�"$b	",����+ �� �I �ߞ����}��5��y�O�5IpÑ���f8��ap|Fa��.��-o9Q�tX��>�m�o3���I��,5�I�5`�S���b٤?���i]jk��e���c��xݐ.�g��H�UuzOQ���9�Ww?����%�������"�GÌ޽��C�A��ɉ2���.���c��7:C��m�G��I��fLOG2� �w��?��!�0��������s޼�N^�]���;>~�D�
��p�:>���';VB32�����L�,1����p\>NI���7�q�Kt�~}X1T�M����!���3����Q�DD��70�s�t}��|�x_���?�JF3B e�v����.;�K��\��V��O.�!	�(��Yd��:�{��us\|�7�a�e8v	8$|�;�}�;|�v��8��7��.����_3.���QS�/��n���R�S_.��Dݴ����Q�+�C艹�^k���˧�l5"����ވ��Q�����-FdۅU*�UI���jq����>��������룮��⺧*㻣�.**㪤��A�@�?yM3�u�)�>�m�$1qph0o5���ۇ�$@��$>�I�<�mg�����b����8f�!��0H��N=�@��"x0d�5���XZ�����D��l-�bݥ�Xh�Bfgʻ������D`�m��.��$wR{u�f��fh�1�Þw��t���&r�&�%D̢�vBfQa<1KL���m�-�wk��>�8����=������:}̥ݼ���ǝ� ����0�j���¤�͸C�`��"%�y'�x�#3]˙��f������S�7�d'9E��e��2�`f[s2���l	,��;��oe?�l�v�M�㶓�Q��j���g'�G�	xP�M���2g).��[˻e2��e��|��:�y��v�~��:�󉪷݉���6o,����K�����;$@o�b��� "3���B��g,��7�����u/8��<�ۃ=c�۽���[����;�K����;f�F,a�*ÏO���E�~��`:�e��Z֦�e��SZ����	�REi�꨹N����.�:�+�.������.�DdD�@�B7rj���5wR�kT�d�4�c]��nqgH�1`��{x�Ѯ�x��s��x5���gE�/[5�nu�e�L��_��8����D<��W�m	8�wĝ�̽�^�ŨfQ��g"eZ㋢m��ǜpk���ڭ�X+��)�[¼�Ak�ӭ�;;J�R�ͱ�chu�͙��!6��P4���kͯoE�x�N�j���5ȚK�}�׊_�kVݢ;J�Ma�5Y(wj�c^� ���0���u)�������Yw�6^����"�����ql�\�x2�s�7��T�zg���!ye�����z�&�^<A7˖��\��{���o��po'z�IW����!��E٘6[�k��U�P8�뜖㣃�v�$�b���}�E��z�ðI��o$����0���g;U:vy1�;�oM�˫�:x "]�NG��H�����p�l��љC��y�e�v�!ۼ����m�Y:W?^���M��v5����j�����v����fW��2��-�fTˎ����lؠ����k�޲�\�3����$?�0���$C��	N+5��Dl�&G����V[n,�sxc�M2Ĕ!@n�e��3pշuwz�K��<�d���<��a�x���8��=�=�w��˫�:x0�T�'��/��߾פ&e��^̫a�W��,�^o?���FmkI�	�u;m��qu���9pY��cTN�zxm�r�Ւ���a��g�����#���u�'�~�&�9��=�<�3��y{�p�����I�������ꋊ�;���@AAaDR���|G;b8q����t���UNw���ǯ����`���<�'��6[���>��e���?���vk�'�vX�M��CO/6��v��ٝ�.y�rC�ai��"�8s���	k8�B�`ծq�������y�Mc�Ȟ��f���`�e%�BҶ�D�S�_��R.���ߘ5��1��E�#�e��7�3.�_=�Շ�Vql��~�ƚ��U�Ϟa���I�J@q>b1�Q�M8���bGB��o�@��CksCb���2�[z�tB�`�,�Xr�Ď(�`�j��^�	O�$_r���6��R\�3����qM�i�؉<_�{YG���l��!��p��2�2*i�X���@a�|�o��wb{��5�˫� ��0U�a�|����;�:e�z�3�Sz��`��d��L�2�	[m��=z���Ǐ:x��Ǐ�<i��N��t���ʼ�;�-�~���#���cڼ�H��,�Hm_>��x�;�s{�S�wS�$��^�`���4�(#7ڲ��NMy�Ν6����9�<iS{�i���y��0���<�i;���9����eOj�ǝ��y��*��G����ҽ�>�4�K�##;����:"97��}�gm\b�w�A��'���p�}t  ̬�;���p���8�' U�,�7�QY�.�A�gz����=k��n�a�g��vu��d��֚�(���ᯯ�=����Ъ&�r�}�=A�n1��>7�W�{@����������8����Z�{g�`9d��iK��?V���wƇ^�:�Vo?���w��O �����w��*�K�����<��U��'���͓o.���,ŉ�ɹ���;���X������'�����*�X�w�r�8���gOe^Ȝ�v��y 7�wk�{Þ�7����;���s�q�᯴���M&^öo{=|9�;#�J94Ϊ|M[q����	4��y���|g+�}T�������<��zM�o6w�iJ����A�۲R�N��ˍJ"����	��5��j�X�J ��79�S|������CP�:�>,J;��2nz�;��+);AW�d�������v�q<�X7��8��~v��4�v���s�o��>�\>j������Լ�d����/}��9�8s|h��xq�qq�W'�Ąsp�P>M�
��E�Q$��y��J����nCz��$ȟt�^GW�j���v�e��H���.(�ί����2��p뎾mSk:3��k\�'D^o79]Dm��8���;�ϋ*$��%���#����������yq��r.�mWp�Ί��<�;,8�����wyQ��et�|TeȜE$U7n�8;�:���w��$�[N䨸}k�����W�'q|vuei��H�Xu�v"[n:~�eύe�>o�[����N�L�kD_{t�ݝ�vք�:���i8�I(��O�vTS�B��78$�Ҽ�:�wa�W�Đ�f��e�y�|G6@+k�f���{�n"�2'�֓ڴ��oz�g^�Q�m4�H� �����"�"� �~Ϯ��y9�����|�ϻ��|��C2�!�M�e�exB������������ 8`��.2r��R�T�Sfty�
O�@�`��ּQ	���Z2�,��fQ�Ye�37�ק=,��!?�^^�؞��f�*�������)`���N«��t�Ff�/g{��� 3�</Ěe��n4��X�=���C9�u������O��^�_?���jp�d�p��!'�GKoY��i��}�Ş���a�_h���K!�әOYvm�x5�p�7*�fL�b1��nE�0lE�����r\�u6g �js�k���p���쑯]Ņ��<���è�`2�4y�ۇ`����Gq�:�a���J�u�f�*���5������ϝ�/�	Te匸�ʃ��`Dg�U��`��qӨ��m�]�59ޤG�>�z�}��P��r�"{���6m��>�]��o���y31�P��Q��L��c\4���0n@��[<��n���T"�c�ᤚ՘j�%��dՕx��x"� , �ݳ���[l>��&avH�I�H����uG��6��ú��]-��yC��}���Hp��X��#����!$`�J����G	��&ϛ���t��Ď(vA�4�OG2�ַ��qߡ��!���	H1J='Q݉��]d�e,㧀a/y�1�j̣����U�32�2�a	�E���̾��Oj�@��|��Î�G:��Z��i���"9���� 0�����]Q[�'�]�`��'>`���3�{��MoE��1T2m2����|)�0f� 8����$����d�,���v�/�1�VG0k����<m&͉��]d�e,����1kE�H���E����s4{<�$g�<���`̑�#�{�֩�P�m��ʭ9�'z�FcMNw�p�b��fj�b0�|�8�z�}��m/%㯓��*���?�7�諉t�_�j�_�����,؇�ar��s�vz���O�=����}݋�����qD�۔��.�~,s~�B�X٫��ZY�_�wN�6��5��%��F�6�����,�f���.��YQ#h݀9+�.7"�Ѱ���,�c!��])�K*	m�c�l�5�0iyж׀�,�#,I/i�u����1l��V�h%ٚ5����&��`����eр4�Y����v|n���^����1�,e\�@�n�H���=�=�{@i�ջk�W76;b�X��n������R�6�@
��]�h`�*.�{6�h7ڸ�jxb��>�?0a^ m��x�G��|�t髱�ɗU_Ce�>�dZf�E��}���WY��,e2��,!�e���?�J~���>�ѡ�I��8�]-=��kKVe,ӧ�w���>m���Λ�����*k��/���=zC�d�;$C��$�L{+3w��ܛ�X��59ޥ�xʛ�{��ݰ̶�5�O�gwʽ^@��L��f���jp�H�񕍓ɔ�^�e�4y�5�&�j���XUt��(�$3�\3,�2�!3,�f8�L�9��0�p�ޫ��;]�ZZ�)f�<��K��>vH��}g�[%����}�|-���ҺU�,�gu��K]�1����;@�v�k�L�7e�ԩZ���w(�$���S��.�Ej9�Ou�|ƚ��R���_9�������owc�Za���%�u�B�ڸ[�)��M���r�u�j��&�ӿ�$[��o�g��������yg�`g�����}�s�w?3����KV�b'����.�4�~�y]d�{�[fо�	k㲄�����㯚,9��>�e�8�2sZHG��1��<�W�W�0m��镘g��}W�ش (<�0`�2�@k�2�2֗�;O��᫬��=��M;�D�,����'�(�	��.WF���[u��2�����9�\3��̫!	�T�2����Oq�y�Ŷ��fb�����m8yw���G���W���{13{�[�1�k`C
�i�C��;5�/�ܜ;7�{<�f#�`0���y��dnPN��ck��|�5�Tr�v������?�\CxZ8�m8�V�?3�E�<������v,u��X��C`�3�%t-3pժ#�ܽ{�,5i��w�0!'}��g�u��ʼ㧘D�Ry1�~JYy9\a��m�tW{V�$���e\!1�j��ob��Q��jp��K6��]�F���.6a0IÆ	]E���||��j_���4ǘ7�t�.�	b<Œ 7����7n��fqO����f��2l)>�{)M�+�^gܵg�>!�*W�K�Q�S����{=㞯�Q<�#&w�=���p;�NK�""H���{��:t��%Ÿ�x>�t8��|N!�-X��N-�u���R-�!f>7�Г���-���]sŪ�8���-}7�]��=���7�3�M��@�����Q��}��O�9)a���]j�2.����f����YZ~�W�=�)�����]�Y��1 ���Cb� �\4Q�:����`�鶰���]J7�8.��z���g�e�����aX�>d��fH��O��]*�c�\aq��b�ų_9��s��Z>�9�,�2�!�O9��������7�-`���il<wWu���Y�>�2��0��Fm��0hm��3�a���| 0o��g���'
d����S4m�F���W��u7ޥ��͘@H��$�ӡ����mY�/���#C�A6�pڋ���.�U��V������7�H7�y�}��vߝ#�"��<)"(���W	9���}�8�8	�V����̀���VN~����Jy��p��c��?��ʦ��~M�E�Q��4CYiifQ�Ɖ	8v<�����kfhwz�[���݇�����yK8���H0�8d�	�m�x�X�g[_y���D$F��p�M���-�^M�@[f�Sh���L�E)�}���!	�Qp�2��e<e9�{���������d]M�w����n�������fSa�l&e\$̫!~���r{�ꊭ�1>bh��Vƪ��������z>��$9�֜?�"ڷB����Q�	@l��$�}$|����nm�L��DfR��&�)g<�RG���"�̑�0�4[�~Į���\�90����o��ҳG]u��˚��R�0e�8`����7/4&N�I��>v"�`�?��10�U�b��n�j����G5��p���� ��3l�y�-82D8>��.�<�9�ا��E��F������d^��������ߨ���bM!�vvl�Q8/�<߰ߎ�"Q�~?������ر�@Η��;�����V�ҷ�I�uq��rڒ��V��X�8(�aFk�K�%ڌ�W�+f���u=2�agg �t�����x#����=W`u�<�.ӆ�K�HP�Y҆��ۋpC�Ruӗ+�YB�f��s���ź+�nZG�8��+ҷ�M��ɥޭ8O5������#���Zz��v��l6-����v�vt���R�����O�n�]���:S��z�:��l@)�P�m2�Vި+�o���V�������)q�	?�j��t�v�I*�q��������Ĵh0�>�6���x�0�p�"A�R��ۺ,6��AmÉ�+7�WU�E�T�zQ�a��#�%��B:�èfz�s����x|���G�"�ZVZ����lMTaY��z*{���D8ar|��p�Z��\?�:}޷��q�PF����e�='��RȎ����%^R�:{���a�c-�_#�Ӿ����c�,�����H�$�?�"tH�l[/]�����fvp�ԯ�r�o��)�s]R[�[˶����s9�}f�����������M�9f��h\@b!�XԺ�&�q��2�L	���O|0q?O�<���J�`��Nƪ1������Ta>���=:��ڣ�!�ol�>�ovYƎsE���0|�}�Q��#�T!O���=�%OaNS\E���k5��rrFR�WՌ��b^�.-�)�5����cpޗj7�����*Y����>�����m��tGO��}$��Y�O0fR\0a��ޏ����o;�z�=8q�qvդI��7�p�C�}��~�Ax�fؼ��v�.qT�zk��a��d�;�p�H�����̒Ծ����{�e�j8�P{y�0f�.#���i�����T��C�p�}J��(����t,v�v	8p̑�N�G�S���x:v��Bw��͚�U�WϤ
���#����!�Ltlh`��%�����^��L�f��cS��J�� hmIi�X�R�����H�����,��\!�e�߻�#:��N]M���8Q�b�����D������Lʲ+x����e��F`͈�fV��c�u��_
���x��y�8��Õ�ؔҗ`�E���t��'�#��N=�_v׏ryh�`@;;������Y�r�?2��y�^a�D���6�W���g��p�P��MZ����c����>��k˒�%>��Y� �u�y5yz�W�_����a�nfU�Ϥ%6J�[��S}��6�����ڈ0d�8t{��qr�̛���#��
�˰v��L�=X��ε��ɫ�`̜�����;$Xg#��sp�V^屣�u㨾��/v�p�"�'�Z��뼒K}��˗�Y��&�mD�5���� � d��ݕv$��E\�߰���؈p��?���G��I>�OWoZ&��}>.��r�2g:'{L�����۰�;$\��2D;�n|���ߞH�0�qG������]B�Up����̥�����ntG�����K�H���0��oM;m�f��l���*/EA ��D;w��@`����3,��;���2m�0��µ�0	8�4e)wݞ��H��J�����i�}�@7����&����>�4g&��D��|+�~]����	�`���c��on��F�����N�e�.z��97w1t�䍵TTU���P,4?=� 3>n��o��+�$��\&e�L�*xZI�tՃ6������Muj�ʵ�TG2��$�%!���}��f�f�/���)m�{��-n�7�ڠ�oK�9D8+��v8��мEԻ����/�N��۞������F+:��`͗;׉��T�aQ6��4j����~�!7�-���fQl3,,�$@�Re�<-��|^8�G�6�w��ޤZn�_F��`����p����Ӌ�9>Ի��%���vC���o�,��vF��T�c�~�[X�2��χ�~,�3t�x�2�a�m�2���&cR׳�f�0�z�xG�9p�A�_�yX�3e���x�'��h#�vm����,H�J!�Z!�3x� ���IðHt3��ˈ���nQO�1ݛH��b��>�RD��S��p��$O�
t����o��_�x��Ǐ<x��Ǐ6�ӧO]=k}�U�jp��G&���j,�/#�pz�m����?kIl��O�|���y��e�\I�%ז�t#�'9Y�xn�3�Tt��'a�ڶ�$/��$.y�x��=n=�����"?xVY�\�ĕsޚ_�_Jq������v��=���ruY|5�S�i��+Z9ʞ�v3�}k/���}�c���5z����=���^"�fiK~T��Ǟ˕f|��tnQ�46� w���;�c$Z��F������T���Ҽ\}�x�ԳW�:8����_�t��@�����[�S���}��켵\�$�9��Io/0���M������/�P��1&�Ey������ѕd�=�{�A�;^�`՝��� l����7�e�3�y��V��|PQ�^�|g�F��O��g��/
��A������'W�}0{+~yO=�-�7�� �z���Y���<�7E�r07�ݮa�w����x����[z�J����!�?w�{�k�(���9��;�׷�:r�q�����͞�Uč�x��}��ܤ��lޫ��%��}��osL�W}��@Ɉ�׉����ۋ�ӯ�s��e/��q�=k�N7f��|i��g?�|b|}�
W�.���x�$]6E����|	^������Iü�m��c���#*�jz��w�ׂ���˸t�n��{r^�������u�{`�e8E�a�p4���{ }};hP�X�������n�{�ݴ�zRg���e��4�6>�ۗLW~#�	�K�š>X
!0�ٷP��AJ[���'��������r�}�6�_'�>Me�z�>����Q����ʆ��°���,�-���L}jc"��x��{_^�$\%���<���!$;�N;���ok|bD����d�4E�qw��	_�k���[�;��yw��~�G'{v��=�IEw�gPfWGGVgE����݇gyv�w��$w�"��n�.�+�_��<:5%�-el���{ugg��W����Ϛ�8�2� �ku���Ds۲�;�ޱxuxt�w�w�=丹�m��|]מ�xwe6�֛�u���ߩ��o��~n������3�n�Ңӌmnm�wG?[ϊ��0��1�ve_�K��玳ޞ��Am\	�����u�L�'R���pz
�m���l�l[������F9y�nWwjް�=I��hК�]lK5�tH�rf�]��p=\'=F�K��A0c�����	]]T3��i�n)xx� �v&\e��#��tV�6������k� �фY\庩��I���g�z*xt'^�Y��I�vx�a[N4{z�\۴�v�^l�i�,4����4vx,M���-���;��Tk1mk������+l�J�RQ�Ό���/�S�cM�`�]�'��o�`~9��1.�6lXX�������v-g^�x}��N�P�n�XCaM�C����:ێ�#]5Ԏ�K\�̻d� +4۶���͋#p���f�f���̒�R�fs��فz��g���ۍ�v���+�O+�t�Ï4eхd|��)����^�����[�ڹ�;ƹ "�t��87��k�7f��;c���<�Y�$Q�r0��Dm��=�{F'�i�d����s���:���.^7Ӳ$�^5Z���r68���9-�+t��n8�Q��]m��n�������A����=�l��+q��G��LA��=�����M�c9\���filt"��hP��n9�\���a�n��+<;R����8��M�a,,e:Ʋ�/\�0�K��;=�x�^���;uOl]�BY�p�k�����"���֐����JM��P.�+��k6�ܰu�z�-�/cI���7�Ink7kR'��x���\eĘ����L�K;]c�ڳI�!��3�M``��2��6����7\]<��T�S�7kFx�Y�88�sn�.g���S��Y�.�{Cq����MH�-v%�l���8ibۺ�a��n�%� -��s�s��]�M�tu�p�c�ϴpe�*%�y]���<�cQ�[�5Z��������.�,q<���4�\\t�5��u׮���ԋ�P��d���<����k�C����#��d^�]]����:N�o&�3�3[�� e��A�Q"�Bnx7����1S]A�-�n3iZ ̨����U�0Ж;0�$uWg<sM{o=mn�=�n3lZ ���x�+���±�tf �*V�u�����r��ێϰ��&�VV�-�cRA-Љ4���k���BWv>O����T���r��	.��+����ۧuY�rB�GJ-�q�t�������e�����߲6X�ǚ����5�U�U�]�%���:ۼ�[��5�\7�K`�X�3*�Bb.â���K�3l5���`�j���c�I͗;׉��T��Hvi�H�ԋ>��l4��N�38ܟ8f�!�5�#�	?�g4u� �W٘�i��{~�~ok���$e�x��{����1a33yz��P@����,��\��&�j�ʷK����Ԝs=|.k�?��̻{�l�e�!&����m�H㼝{]��񡛑~������{1<_
��#�����"$�\�Η�=���
Ia~z��iK��5f�^s�6��\��<�
m�� 6kF:�uИ��y���n�FYg'��'0I��L�^���H��b��<��.�2�2l0n��@v��rI,�ֈFotYi��Ϸ}���<��К��Ma�Xqʇ�r��	�wP%�>�l5�,��l' �U&���g�*��eUJ,ق���r��xy���w�c���_?��KU�+t��\<���6[�aw��Í�D�W�Х��n����� $|�"i�'`i��+^e��s1<_
��6I0�p�Zq��jX�?�����43�c��C*90�w��2羃��h��⾍<0��E�ڜL��I�k��h`>��H{<A�p��S]o8�_�FND��f��[W�V�w��?�����8!'q�b.�ӻ��7*��:C�[�߯��Q���X�)J6kLk�dvy5�"m[	#�.ɭ���>O�_�,����y�}��..w.�^{b{1<_
��� ѱ�l�5`�,ݐ��p�k�D0J<�5U�[6�y��f��N�����~����gu��sY}@�<��ۀ�p��]����kUd3*�9�Y�K�����v������Cc��::�"]�{�t�A��@�<�ݎk΋�2���'�@=X���\�x3�F�C�_�ǳ��eL[��^�YV�gxm��ŕ{�n�ު�}����n0�p�H���#���{`�su�,[���;��0�qӋ-�z��ofS��>��>�k�UJƎ���-�n�p|BG���$��$��6�u���G�#��Z����l���_F���K��>�A�.���ſQ�~�}���?�!�#��$�l�Z�җ:xI�,��8���SL�8�J�R�������|�e٘0R����`�'Z��'�ھ�n�z���ͽ �h>�z-���'ve��[�:&�Nv�o��~�oI����Y��K-�j�b7�)��L�8�QpۃY�p�H҇u��ٓ��_;�0��'�	;������rr!Q�N��m岖����>�R]� 6���7e�`�v]��p±���ԘUY�A J����D<uc�p�Kj��.�Gy�5Y�=^>�xȋ�B�cS���6�M\t�y(��-�t��6��q���ck����g��<�<R�]U���H}�֖|���xxT�1�|���<�.��$|�I��9��7ٸy�D�N�cE�3.��St���<_	��`�1uS�ŧ���Wu�z����A�j���"M+Z�].�u��
+���n�LS����'����,8މ����6{�����+���f�\��e�i�0Yx��2/�r�������\7���y�#�~s6C�m�{tl�\t�;3V��È����<���5�]ꃞn�,!�0n3��3�q-Fu�Cx0��_���b.2O�d��fH�V�����z�Y1}yQ�����!�5��]���òowe��0�a�]	�l�&�v�1���^�~��w-uY}x0fRO�Nb�T�^C`���.]����G�$C��$��"-��s^8�3�9����U�5խ�?8o5Y���^fN�`��|����dPT\�w����E������'�ox�7a;��7&_��S7q<��V���iƦU$,ܦi�������$����E�������Q�>������ya,V�t��5-�ӡ�[��s��%{���Lr����R]ײ�ilXv]l�*ص#-%��]�k��D�s ����T���.��݉���60�ja�m���ݩ#�u�W�� ��[��F�-n�x���G�I�W�<%�f����8}�h^��ê螹�e���{Q��Wv3��<j�S��ο9~�v��<8[	0;:�]�.�	���?���.
�[�kk�-��� �s�].���0ۍ����_4�v��H�o �d��;"vc���	��"B;ܵkhK�ݚF�;�;v��')p̑@�ԥ�d�nz������uEoK�v𻖺��� Tw��o�d�Q��`�Mg]���׈Xt�Q<��<��e���LM7�����#��Ue+
Uw�����S�P�
����'��"���a�|�\�G��1�n�=�8�zI�6I������Uα�^ivC�s��Y?�!�2NWC[8�|Y���o�\��ת��"{��ܵ�e�i����u��H�`�d��EV�CdWd��$�D��vwv{9�K�A�+C)30���qv��[V�y��e��6�Ѥ8`�����8E����sG%�z2���_�\�ru�g^%�[H�!��}����l4�e:L��+Q)�O�kvеQ��<�-��n�y��7F��b��9���'���Y�."�L�W�f*�<LX͒��ϖ���j�3�<=�?{�N`�e�ot�Ǚo��ٓ��$��d��`޻p��7m�e�l!���*n�L���3,�f]�ݿ{�M}�:���"&��]�]V^ƞ�'����G��xFoud7����֦����J��|��G-�!�o��p��oۭ�����]�~p�i��b\�n�J�w�h��7�^�����`�k����H���ˋCh��Ǚl�n��{�G��G��n�8�2Պgᛧ��@OTMǃ��Y�8�Ƹu��Tۧ\)�Ro,q��(�uX��Z�|�,���9�[sN�_0�{����z"w�Eܵ�e�i�4BA1!�l��m�o+�4M��Y��a���߻�Ԯ�
zC��8�����ھ�̵އ�8oO�Y"%�OOp*����5���ߞj��kQ�p���3*�A=>U{��:\��*چ9�O�g(_LԼ���b��y�:�W���{v�#�S��H�yh�Ϲ/Yᕳw�-�ڸ�uf�^�,�2�-��·r��e�͜ˉ�E����d��y�y�!�����^!���-��E�4'�x9�@Η���d��.i>�D�o�k�����e'ݒ�����\ը���z�a0`�'�!�dGx��\__���ÊY�{�y-��7�����M��$��$|�I��:��g����>y���~K>Ƈۅv���ِ�i���c���-��MMAWR������{?|9��G��;[t��6�M�9��(����6�G���d�b����v�8���.fS�oSZ�ޫ��<�p������'��w-sY|�y���a�}A��[���Sܶ��!��x'}to<GY�����fd�DdnDAڌ<����yu�w��dIðI��#�d��ËQi��r�����f�s�`�̑|��l18�M�9��(��b!��y�}���Ѱ�	f�DD�"�F��S��{*�zo`~�U����c���t�3P��X�r���G�^=ΐ�~]ܹ���ʢl�FS��aID�>��	��k�.Ϭ�fYdfe��Y�5�������nK��{����osfk/�Oy��Z��_�Y�7��8ar-�ʌ��!�������>]�hݣ�5tS�.��$ɔ�B��!���J�7������O�z�#/�de�1n�k���Jw�-�+�y�;���h0�n_���~`�%����I��ș`̑pQӻpCG���0�s�6�ي��y��n��ȝG�1��3��0�ۡ�Uc��}|���]�xC�o$���>��o�}:�T�;��8�zO�7��\Y������.�����H�`̑����?���w��	�Ձ�D�;^��$��q���BS��o�]�~p�VC��o36>`���{0Z��8>�=ِ0k���#�s[�uC/���y�5���]&:��ә�<���(�C{�əE�fZz�O|�3��w�5�09�^�����خ�²�_"��i$�}�E0�&L՛��L�D`ږ�S�ԉ߽�c��n�
���>12+`֝�N�Q��|f�X���l�>�7���������S\	Z�i�������u�5JKYis�e%�]�i����M��+�YƇ��k[8d��>�չ���Ff��"��=�#� |�:�v�y0f�� 97�qk���{��0=Y1�&;]t��P��P%�m k4F�6�2i|��C����v$[ۓ]�^6	v�eƣRP`�C8�[���?�}Q�ҩs#��YM��G'2�Т�P�׍]�cK�aRgg��_萇s�,�>�cU!˲�M�[}��{ؗ��"��g>�ag��M9R&C�8j��`�
G�	���1t�/�����:$4i�q��׼z)NnM�eo����!��N	0ʚ������Y>;��;�`�ܳ��;�gqG�dkjD�D�"�i�<�*ÙY�ZO�6"�]�q^(��D8`�����6���ž��k�����w�$�q�X��'{x,�3Y��{��5�p��b櫗c���V�L�Y٩(�q�-�s�a	�����Df)�mO�e�@���=4�{&�2���sU�'�'���O�/v���ϓݶ[��|�l�A�حf�fM��[gA&�]�+��t���ۍ�~�=�����Y�?�"�2%�D��8�<{++���woz�T��w٤[�r"�Rw�	$D���v�2�c�5���vq6��a��|������nzS���N�����t+a
�w�&m��;@wؘ�3��܁e���=�'����  7�N|�l���g���'~�M�fk3�O�5˻y��"�S?��4{��§p`Y������0Z�N!�������}��OuJ{g-�+�����`�'R�fZ�BҰd��#�7ǾL`̚�^��0fRW���q�8�;ϕ�����0o6"0��YY�z�Vך����8`����^P��%q�^��w��u���9o����ɟ-�fs����\�?�����H��0}�vEs�'�	����تO�a���\ل���]f����7s�0����fg��#�Q,�aH��$�BNgz�9��N�ݾew���8��"����G�=�/s��{�a2�#�VBY�����\�K	��.ެ/�"��'�Oed��2}͈�`�n�!��3�t�WV�}�,��>�E�r���,���3-��]�;}q�ۏ��<x��Ǐ^<x�Ǐ<t�ӧOZߺ�5;^]y�VaE{�
 �����{!�#�������� (7޺<H�\�i��s�>�P��پ�?o{��ݪ�����ҾЭ���p����3w9���ʍ> �q!�ҿND�Ϻ�7R))ni��8����ok��ڧ0 ��圇��X>��R�{�h�+��S}DG@v��)�;��QL�q/���H�3������{��w�>Â�#��{a��n�=�&�)��V�y�{�������g`��7����� �<��v�<�V�����ؗY/�Σ72��B ׫V<g���=^8<��������}(�o�����х�;W6�����t6j�ۗ��i���}�<or� ���_��UWݞ]�"��y@1�1�'��j�}�l��Φ����
p+]M5<��#�}�Q3a�?y�X�x�h�Smp��}���{K�m��|�+��-����x����'�'N�Ǜ��l��N��Cӝ��e���|:�g�u1�w~Tx�YV-�&w{780yE��g����P�1��M�&y�?N���������靁.���!���'e/�wq^vOaػW0�rW�z��$vh��kg �ۋ�C���5i�.S����[��d'Ϛ;���IV�(ֳ��7ۥ��/�9����\����4rƱ&&��0{wg;R�0���k:�I.{{8��<_zF�'(*v�K�Aڲ��Y�_e�"�#T��i���"Zƛ[p�* �mK��.\�I5�~���[+�zޒ��� ���n���w��M����}�՝�������܎{z���f�Y�y{��t��-�6��v�-��I8�
�����3�6�YfVS��q~>������7{�|{�W��]iW�瓶�<�3����vT_�;�;9m�l,����e��$�1ټ���w��΀�!���Ӿ��ӽ����������:����{y�_���qE�![���vv_-�{��|�=���Y�����
�M��:;��:`��Iq�K[�Üw�LYZ�YH%ʍ̕@�)$��M4��;�[�~�L���}?��%�7����H�#,7��wE������X`�N-���;vs+��G5"�0ڜg+��+�:
3�l�[sܫ�&e�0I�쑼̒�S��&3�~��g�t�쬜�N{�`�d?�6c�3�� :L�~�D}gγ�/ߒ���1�ٛ8%sqkx�]���넮lW4���*��m�v�c}Ig���%�!�=~.5�8.����ó�O���ɔ`��ϧ�/5�E��gH�SC��τ��P�v�z����!�qhk�tN�V,y�Hv����Zw����rÙ]�~p�d�,$��>d�K�y�l�<b�}�k��Ӂ�r_�$�$e�H�q�n�RucM�E�[NP鳙Y9<����w�s(��3,�3(ӭy{�w��M�{� O8s��G��O���ɔ`��ϧ�0l���}>�
Fwsy2��rg�d\�1�<�)��fI�l�bB��w;�o��|X�����"���g]�i���es�-�7�
�KWK��D��}�����i�U�̫a�E�2NH�������E}IY�ުF7�W9���͑��\!�e�2�e������~o��l�>�=�;�T�l,ce#�Dd��(��W�v�늙��D�Qeu.y���Y~�9���$d0o
�D�閭l9C�Oed��2x0�U�N��s������^.�vn0d�pB��V0ot��h{�xX7�������['Oo&Y-+3�L��f�>q��2G�]& �� o`�{/^#�Ǜ�$;�vH��;y�(�^4Φ��~�r�U#���=�~�5���av�?�$�vH�y��O������}���a��z�'��3$_�2Ս�(l�쬜�O0`؊�C.)��&h&�!�0���/��8D�a�����Y��ח�ϗ�v2t��e�ҳ9��`͒]�m��.�H�ޏV���Ϯ�8�N�Z��A�=&{5���vJ���vat�@i��S��<%��]��=:.?��Ж�Z�x����6�)%���b��*J���$��o0����-�B�-�v�b�G[e�ș�;���:�xq%Ƹ�k��ƽk�O(��^�{f�l�v���l���"^�k����HN�.���R��h;lƍ�C��G�9h�fЗhrf��&2���t{jKW��>�ۭ
��v��&Msؤ����s�.�^���3F4�m�,*i�Ҭ���v��Τƙ��׿��S�1�HlCvG14�3�.b��k��䦕�8x%�H^�-?0`݄;�òD8`�8qs�\��z:�3'��ASvo%�a~zn^H4�_K�f�O��$]��v�3tf����.��f�`���j�Ô#��+''A����k���8*��aÜ�{��C2ˆe��;ݾ��e��f�8z�2�iY��}��W�k�;$|�0���0�uV�D.�*���E0�!�t���$����\����oy��0GT@�ٺ��׉�h��3O�O�̑L�>H��V*��\�.��Ѭ�mCo6���Y9:����òD;�O=~��>O��y��F�M�l�qt����ur!��2���=�hII�Q��?������/�do�b/�;g�0�3w�%p�;ϼ�e4��o>���f�kFo�#��O�l��B32��U��,"z�Mk������%�Z�\�H�՟�{Fv3ψ��>�w����|<6����)o��yMrn�؉*͑�5C埀��}��5���|�l�?ߪP��{����y�����,��1�թ��!x��`ͺ\0k��E�y#�2�M��nD�t��m9B���9��2]?Ne�ݗ3(�L�-�e��D��Q�1�b9�m�d��B���~?�f?�u��Otn�,M+3_O��K��A�J1��uh����ˀ��g�")�Rp��P��'V�=�R�G[����88`҈0d�?��?�'񼧒�ld���XI�^������]t1�]k�Y�1km���}m��n����Ď�>�>~��H�`��.̵cY��{++'��0}�컾���D8�QO���E���[�,&ee��T�(~�e�o��v�zc5�$�F�biY��y�����0���W�(6A�r�	��p��\̯��{�1���5�Cb Jg�~������%��twW���������*8��Kn���\v�+�dsv��<��êJ�V�8N����>Qiݺ�66��'�<|�*!�`�'� ��'#>`v���32�>� Mo$O�%ڱ��]�������C���q��%��{��`ݮ<r���,8��b����
,�`�\���,�X�p�m�־����J���/����8�8d���H�D&[n�k�..���������*Ǆ����aIc%����S��jL�K�C6�8�?x~�˾��~�Ŕ��'�I��z�sG\^d��s��f�͆�7Z@���ۿ�'��H��e%�����n��Ş['��;���{��{53j쬜�Ox0o5�8���dA����������Fdyטb"n����$�|h�۳�Թ��e�ɷ��u���9��l����H�`��./�]���"6:��k��פnn�f�ި���=��o����~f�����"�MIt�]E(�0���
�	T�ы җF�3M��!��s��G�g��>�E�MS߆�1�5��s�_���C����aT��4��R�ـ��?��#��9����BR��w�]9������C�av��#�" 0e..6�-��9YA�d�si���<Cz<n��5�Z���\6oX�[4Fh�ٮ�=�	���~�̷a6�)���Fv�d�=�St�ٚ�y�\�0�_L��F��F;��R.�H���	,�{ѣX��vh����e�|�Lۛ��b:�'�g�3*!ǘ2N0I�!�����{�\��o�C�U�8�8jc��Q܆d���Gg'�֪��#���x<��!�0�$D�H�`�����ٛ�vr��`�N0�p�H��^�c�����{3�H�*v� ��S�Vz�8�x���������!�]�$D�sӧk���;��p�J�^oWM���̮�;�6C��D8`���Dz=^>���1=SIĩ�=�لB��HT�|����I�.qT㕶��	��M&0�Eߞ(|�=����ەx���c��`�����2 �)��%�`"�
���8�x�s1���z܅��]%��dv2ط<b랽�㎸�t�2��/of�m�s�=�>���lF���7.�&��h룵�E�j�:�Em�&��V<\��tsu����k�n�cHv�h[�$Y��PR0�g�Qwn1)c3ɬ��H�n3iu��NpLW���g���hJ⒫#���ئp;3f��?���g�`��Ƙ׮���D���|�ԉ���jL�Ga�(����O���g�l'����/��G��w �ՖzVN�G�
̈́ Q�ia�r��0���p����v!��0�#Cٍ����?����	��Ǔ�;�o��ϧ��%���;��d�[?K�l��|�$��O�wt\!��l̢�@��f7O�v�7%�sau]fOx�?����;�`��2ß���͑^�g00�;0�w�.�c���նzVOF=�W�e�h��Y��ݱk���0�p�����`�8	�,-��R��:�2`�N��%^k����d����$@H��Է�����8O�8pR�@T���8I�s�]���hnu[mI�l��4�X��y��~���;$C��8�H6��t�]J�'�d��aQ���*�^�f]^~be�Y�l3-��B^ex��*Ȕ駜���c':(K�4:gj��P�Nrp@�V���.���n�f2�e��>x���Ҧ1-xS���ɛܧ�� �u��Ͻ�\\0f�/��)a�V���,���3e�f���2D�P�}�0F�d3.�)�,��Yp̻s)�7�9��Lu"21<���*�O�6���?�H��p�"����y�w�mp|ג��~-d8$����ޮ��Vd����i��_o:�R�k!��>��Ty�5�ޯE0f�.��$U$�d;D�����+k,�,��G���,�.לC@z�gb��d��{dX3��ɢ���a�6�6�`���K(�e�3\%ci��HL����Ѳ|��`�\8`����?���3g��]�*M�k��0\�ޟrZ|�T�|:K��1�'>H�d���!��Ki���Gs�ԃn�r�e,������O��}���A:ү��n�o,.3�v�p�e�����ޏ^6��Y�B�QO#�:�60�M�aw���#L�p�w����E����רo�y���Q��6�8V{�*f��؆>��y{Zi�@���/�'�m�
��=*3�5-?ۇ�$C�d�;�8�ΤW[M���?��p���>�޽��5[�׊M�s����a;�6񃟘V���w��'����U��f���B�òD_+5�3��0h�8��fsmu��+2{ƹ�� ?�p�w�$�㋡��E�ԋ/�W���Wۖ�κff�\J�\�L`	`:ַB7ST��q5&w]�z���Y�ϣ�_^e��ػd��	Ս��v�)ʌ��<�yg_�5�j�40h���?�7�p��.�8f�!�\Wp�3�Pޜм�1���ۿ�\���q�ކ��7yϧ���we,��c�tdD���\MUm��qhϘ0m�0av��"��n�eoM��zЃr��V�������!�2N�>v�$��5٠�K�[q!V:��"�n��/�N��j��<�*3�I��d;x/?���3rļ�3*z��)D���ӋL>[�k�g�H��Lrqf8�6��\AΖ/ f/e���F;��4�T�z[��wĔR��I	���(b�����>������!F���7�,��f칶]ՠ���+�����@>�,}�5[�g.M����`�n��7���2ES���?p� �̉H����!��n�����\/�E�m����e`�-3��熰`ф8`؟�!�$�����v��|��'�k�p�+�.G.�0������?�2E��p^�M�/܇;�����hnr�Buf�����r�84�`�6Y�v��"��k��pU[��	9�nI3����f]����vV��ۍ�m���}r���}<��n��q�HϘ7�"�G��*[x�ճ�Zs��0�p���>W"��w���̞�p�t@��y�!�V��^c���r�{�̬a3-��V{9>�sטj�Mu�l�YU���{,��n�!�2��c��v��v�Ǐ<x���Ǐx��ǎ�:t��V�^�3~� ���@�r��Yhu"�X^�y^�u�:�/�9�̰=��Sؔ������ ��������O��5�3�����Z�+��o��O+d��Woo4<��W<���,��$W܏<VO�Ǖ�B/V�u�k_C�2��U�c�w��g`DW9(��.9�ý[&����1�=�sܩ��e|y�:'��x&̅ʮ�]�O��N_(F`����K��޹��gxzy�����3|�Z��@̸�;�_�����W���CO�n˛�������E��>%. ��^ܝ]g�0s�:^�`]��u}�rw��מ:
ݜ���D�n��3G{�i����t��>�7���X(?ڽ���G�ǎr�#�](��"-������w[Ͻܯ{����ͪ�������9q�B{�=��|����k=����$�HoC�P���=8�No*���Ո܂q��7=��$���ި�^�=�/R���=�ץ{X]����#���8����Ǫu�C��%��&��ف�}�#��v�o���њ�ctpӹw�<��=��^��=�4ko���\�]�2�̻ސ���q�Q�\�hiO�������"ç�ͱ�p-����vx�g����GnQB��j�� ����Nu����p.���,� x��1�y�_������D5s���ot�������٦�w.}L �g��Y�r����-z}��J)p{�Y�P�8��|J�Fq�j���������óܠ��3�����Q���K.1]��(1t��P�%�	F� ��rZ�]c�m`+o�ޥ��^ڼ󼲬��.�6��^^$Y���d�q׽���w'��䭳��L�7��|�o/������W�y'�Ί���2����s�"v���;y�O'߻ޔk-,,%���5��pqm��J����C7��ypu�eN�������gbI/���ږ�M��ؙa��V�6��pY%�ZpP�X��Ŵ8����a �U�/�u�֓�:��S�٭����3_7z�f�d��|\g�w��{�A�gcM�	O�)���6���-��i�||W��,�f͚��b1mͩ�V��͘�cb��Onl��<O,���Y{��ʖ�!��[�b:�����<�&���q>��5���N3�ᅲV��=���~���#㒺gDQ�hy}wc��qOn:-] �6��3��s�祻4��nN�E�ys<�LZƞ+���K-��{6	���bYQ3�]�bڌIaLGMqB���/a��z��Wku���i��cMf�[�	�B8"�Z���e����q�8C'��"��������F���"[-�K�0ʖ]ɮ%������	q�2v���v�Mk�z�&�h�#U�к���њ���b�a�X;-9��6[#o(�A&-It�q��d���31��fڽ�L�Ӆ3���9h�b�45ɘZE��,Y���UCLt���nٌl�K�����Y���˙�k����b�e��.ɮU��vщ:8"`��7ZK�ڷ��/�鉸[��	�鵧�V���T����s^��������,�U-:��k35r��HԬ������s۴Z�H��r[�:�k+E&���ؗY��܂�a��K�{kv/n��=��2+��h��K(�i��)@���j�l�f�x���ݛ,�t�U��2¼����n�I���%3��[a�mncL���Tta1.ơ�7F�L��P�E��n������X�[���5a�ݣY�+���`�� �]f��',#�ݗ��:婽���ɝ�]��e�(Wl���đ�L��,7f��H�*l�R�GjJY�p@4`�Ǟ���[�z�cR�m0充��Qр4� i
��8�us���<6n;=Y�FB��걚��*��$�qjK���'��d�7s�en�kڹ�.��=�L�7�]�v�9� k��Ms���zl��7-��h' ��*�]�=��UR�l�3V�CV�Jn�)QhF0������M01�}\[+)i�k<�ָ[1��-�D�X�2qf[))'����\�4OY��v���UUUUUUj�W8�Xx�1e�aqsbB��4�'�<����wy��i��qu���Ga�F1���7WJ��$M�\̴��]a���%aD�,��3�A.�̹�F2Vh��[y���C�bk�h���^y�㇗�F7���8�R0��RC"��%�b^��l�`	����-��vS��lqFu�c�Y5ۂ�j󺀣���h��n�V�f٧���߯��~\\{��v�Śeܘ�N|�\6Kد]�[^H�t:,�_�~�{��Y�(�C���e�̶�V�w�b�\�Y~���Vjk�%��W���u��v�3�s�T˪a�^G2��Ý�m��{������eV��79X��������N#<�f32�ll���{�a������G��a��fW�s+�R)�̗}�3z�ڢ��VS�ph<¼�g�!i������R�y���Bv,/t��\?�U�ǘ���Vq���Y˓k9���G�=����������2əV�2����YfYd��G��H�li�~ls�?�V/���{���H��`���̓��N+rI�n�Z.�唗��P���O�f�4Y�f�B�+b3S��r�Z���bH%�0A�<0`�(`��_!i@3$_�B�s��7m�e=g���uim�����2��ww�ԭ�d&e�a�퐊Hp��O���: �S��K��x�ueq�X^�J���|����bt�0m�4^귵��C)�ݪn�-�8j,����Fr'��\	�k�α�ȯy�L�k/0NAeJ��L0�	_�N������s�)oE��6��O�4qp�������A�էk�M�`�m���8�$D���]��gd��R�k���[3�y����B��w���-�e��	?�Y���LusB����`�:&��H϶���e�7m�e=g��͖C��!k�{���-��/�0��N,�̢��[ݗ�7�مo�qݼp�۝��w�e�6eѵ��@�<7c�����#�wP�Vj�Ɂ���;21`3�ϡ�]Ok�n���i�9ճ�h%����A� O?�{�[���vH��'�[��;�XQ�W��5�&�e<�RB�I����뿚������0d���5��:��,-N��<ץ�3f�ʪ;�-Q���S�ph<��e��֜?�"M�\q`�\�� ��0��=����7�-��M�e���:���e��T�Lf�j�:X��U/r'�R���P�P�SV2�[&��6���*�l���E�ʅ��Æ�F���ʁ?x]���[{�)�a���<�z|�0�|Ά-?Z`^=��-g(��V/���IÎ��w����~����?x����\�z�!S0b�kG϶�$e��.��I�쑧�N��Tk���6�}���d�n����0`�d;�p�!���N6�':*�4��ƭ�1bY��wυ���*���Z�9�u.�<v�ۭ�k��v�2���?f������2�=�c,��z���Y����m�6,����x0ӔQTx�v�'���e_7��)���;$�sAi^;W��?�$@~�vau\sa�y]����w�\�֜w�?�fc�����L��ç=��9ZbBkuaf[c$|쑛���m���n饒j:��ʿy�5Oӛ��@�Yg�eQk	�e�ʱ`�ܼH����=��+`�?��^]�oB��l�����y�7Iv�>��y��vo���a�ܹӐ���!���p��w=�=�_g�#�����4�79����j6�N���	���>y�o��!	���4z�w��n��7n̑�C�s9b�w8|�����ퟦ�Gx�y�6Q
���� ?�>�c{��>T"$�e,kM2���ٮ-f���p�3JݠF�b��g6M������/��� �?��˰a�0ƥZ��jv��e<���0��tKgl-�kaj\8m��$�%!�2D;":�CF<��0�?�f?�V����[}�tֳ�Ot��v?��,�0Tf�b<�ۦ[פ;	8vH��"�S�gs�٫��1��z��~/��S�٨G��ț����陟f�3�tjs���,�.2���5�v���s�I��d/L	��t�f,�������p�O=wy�̢�<�j�ܖp��K6*�fϵ���{W}��̫!&et�Y�o�2��9���jr�>ڱN�޻[�=�{��Z2�g5��[A�x��~ٖ�-�Ȝ��6p�ծ�AÎ����Y���y��Y��zS�>b��Kz?�V���-ф�;s�l3�`X�ݭ��-,s��l����ka.�X�;P*������f�g�	0*`GL�LMm��l^0�pO��.�\��l��2wݟ�7kNiM��6C��0�`7��ث������u��to�ōĞ�n�yۅ��^6�%8�vn�ĵs�S��.�>��X�g[����CKI���?F��dHA�X�j��@î����rZ��r��4��?��`��p��征v@{�3��l�u�\t�q�4g��2�rGR��V]�2�2�'��eӦ���<!�5W���\0f�;U9�;9�s�9���{,�`�Ӈd����dS!>�p��xC����v	:O�'2��3O�2�%��rֳ�O0f�.ð��"�2G|��e闿��=����`�b��8�`�b�$�>���k�����;�vO���*t�����;�z����f���M�L�ӽ�-H�N�>������t�tTt�E������0`)?y��n�v.�@�㱐�`����.i���K(.�2��#���'3�c�ݛF���ؚ�3�g��і]􍟽���N�=v+�	wA����=�O0�z��);��s��<�]�q������Z6�7M��"cm?s59��o�^��^�e�f�� �5x�a��ͽ�GY�or��8�5�5��j�Mɇ��t�+x���{�#f̙W�9g�k��Q�w4c�D~ �ެ#�6�=���w��9U�w��?��p���,�*�n��V���F��c��p2��	�h5�f2�ts�d�������A�C�e.6z�� ��v��]ǜa���QR���@��q�}v|���c��Wt˛7�y�y�����]2ao�l����� V�`�v"�y'��.��7�{w�(���2{�[=��'���.Ȇið����?��[U(�v̩��O��Bs��5�GcQSK,���eH�x�<��۞Z�l��Ԧ��ÿ���=e������6X�ɦ�헨�ތ���'��A�d��wy�zC�����d!�ivљ�!3(v�k�YV��.y�3w�y����]�ޙ]��l�ti���l���;$p���E�h�1�ly��a���²�&e�fY����]�z�p�w�k*�y�%{�T�6U�W�8|�4����\��=י?æ��q�����-����ѫ����]��N3�Y��1���eܫg�Uwx��0k��i�H�BO��q^!��cAM���1�0g<A�p7��fH�M6�ي����|���y���Ȁ«ɩߛ���˵b�jY�5_`�p�W�ٻ�y�i���m�����8���O0`�'݇�#�d�l�Щ�*�}`�ߗ��mm��qwU���k٭/n���b�ڥz���붆O�2I_�S� �8��,Bӛ�7��x���=�6�|��;�w�|��K��Ik��GXo.��l�[�j&�]��z�^؋6���.�ZX^_#:�^�D6��5���`�82ap�7Z6r�p��2�xGN������䏚�k�M�UYw�Vk<�o��y�6�v���;$\7�E�=�S@�lp���ia<C��!��2�wOwE��*���\��!��=^>˫w����m+Ӛ��F_N�4W����I���nUg���l��7����AXJ��@]΍/A��8+���Q>
/o��g�R���2𳌅��-f�&0�8wa�$�����V���8�42D&CI������ 6�|�8��]�R�9����l��!'�H�`�����6�Mۖ�4Mm9,�/��A��7����st��u���hX�6ҍ�nek3�~�~�7y�v�8.ϝ'�]�c;�Ws<�$לt�-�&fXWa���ip�H�fE����]��0�i�1�et�y��Hp��\8�t�t[=���p���v>ci�HOHg�1��P��z����`��ǈH�).3$J����� �ɥ�O99����l���"$0d�;���{.:B���D 5K��u�8	?���f�Nm��JMy�O��#���]qu���^mD
FX$]��2	���#"Y1U���L��#GV7����类�W�d8`֜8`���Dz=^>�Ϝ,��;��
���Q3Mj
��<���h9?w@�W�����h<㮲2�}E��v*�[��y��Ǉ�\�����jC�cC$
C�̌1���sՕ�<lW5Iq�����&;m�`�;T�S���*! m5kN��MV�n�I�N݇�c�qt�=-�z�
Y�w��L`�k&�9�݆�Fh�P��%ؚQ�g�]�m������0��p����+�A��x��m�-�P�cN��PYFk%L��M��Ӭ��d�g��wZ�u����!o̈́��;b���*f�B�K�~�V��d6�f��}n(���;6�4���5A�&��&1�0����;����*�G9m�2���>kz�y�k��5�ݔ�jo�%혃��v��"%��?w5�T�p�1���X�vG�2��|��l�o[=d�k�:{�6˻;��Hý�{,3l�&X0�@p�����I��m�ʨ���ˤr��U]���;��xM�C2�e��ʶ��=�w���L+�������#�P�[=�O99����0��Ԅn�;��	��v+\����0K�у���f�m�����[�g����M&��G�|�G���/��م���Wm�fMh;;?L5�4��0��@ aƯU�Ɩ��Heb��R�J����%V�Bktw,�fR\&e�ɭ��z�z�_U^G�:��veo1����������.���wr����IrG������cѭd�ڈ���/����>�O��P��wyr��[�7���{7]��屌>�0��u�<;�]�l;Z����*���$G�/0�������7|_��i�Ml��O99�	��`�>����*�ZO�
f�"Ęp��m05x�a@H�R>ĆW���hŪ�Ng&�fq���/�����ax�E���t�����|T����`��8�����d<M.�=��0�����u��7�,�}�ʬ��V̻͐w����>a�م�7��#��:��z�!@1��̪t;��Ou��Np�y��C���p�|��'L�a�;�S��5�/�J�/i�KQJQܖ�T���6B9Ӡcq!�#��l��8������I�80I�̓��,l��ݧ3�I�4��m
"��c�y����U���`̑�A	?�I>"��.�גf1GT���8l�_V�8�#��������ӇM�U�us����m�o���3,o�ou�@��7��]>8�뷯��<x���<i�Ǟ�g����z<��iݤ5C�8n��cz_�ho�����'���L�w/�k�>�nq�'`������Ӝv���V
K*�IwX�T�Q�	��í��V-�t����N{6��sX��n���n�/<"��~]�m�듄	�>�
�1=�^{�;D�v�\�雒�}����7<u���޸��ɺ�A��v�����x�����_����f�5go�_-�7�\e�3oKx�s�8]�G/g�vV{�7��:`�p��ͺ=��y"m{}qg,ۻw��8��$ߺ�x2B��w�=�(4MK=\�Ҹ����)��J5�a��L�]��Tד��o�{���{�5�Σ3�[�0�l���N�(��w�磢�=�Ƴn­�f�����/vuZ��o���Yr�sDW�!�Y��KWm/�i�y����zC}����s���m�w/y�ڤ�K#7{{;Ms�rS�#�N�&?�q���{|# ��=��["��7�>K��I}�#�Gyٝ���Er��ψUL��lMB�>���$�nw�ܑ<�m�X��V�ӏe?x{<��\T���ۖ(�ѻ��	���z��g�ɷ�ݶda5�82p�QVJ��>�+,5X�F�X���<v݇5f罳,���wo+�� �����Y�43u����&��2���J�@r��w�#Z�t)��^+�V�>�E�Ho47V��}�����4�����qG��Ԙ����;�����.�y�%��m6dG(;��c!���`ńi}���C5g�=a��d��5p�r��y���jt�>��Ǟ�;�>'~`�D���Q^*ʯ�8��e6�B��$_Vi{��B��6ۭK��׼G��zw�c��'��;!�J�l��!J t�2�1����k)�6���{�z���a-�b��5׋5�
ƞRێ�X[hZXJT�
����%�@c+�ޭ��@�x*��%���k�/_ �e)R�Ė4��������,����#����k{{}�``*�*p����$/�����PZ���)�pV<D���x��$IB�@��yM��M<�[s6y5�[���$�K<e�k9���K���$$���>�Y�!,�:fy�9oo���ܯ������� �|�ϝ�͝�Y����e�&�W����x�ݯ>{�[�z�mé�j3�m�[�Mmj�=�r:u��f���VZ��9��H#���5��qsҬB����}>/Vy^����Y�S�,�`���4vm�ӹ�����A�ڋ%���X�6��p�謰d�6�`�N1���ޖ��n�����Oc�i�{�^rs�A�6a�p��"�<�삕�M��DC_����%�̓��jX�սNg&�fq��7I�(���s����
��@��K׈D��3$C�o�8d��n�5Ni��~m�igF�\�!uf?y��"���8`���#�W�JZ^g������ ���~�����@C�4���D�D69,�1�U�aX;a�D���1�F�3r.0��$d�����l���ܼ�憃�0�Y��j��8l���$|��y�k�&�=އ�a���8�K#z�����l�:y�7IpeÁ��v�{hD��1c n���,�Hp2N�!���N ��ܓ�.k:�u̺�V�"���������%/�	?�*�ً��0߃2}]��naYȓ~��} 3z���l�ݪ}��398{0��������K[�83z1aÊ�ں�gA��0|���Rr�~��-�5�|�C�S����'�~�x]���[rr��5Y��p�����"M�I.��ƒ�>l�ɼ���V�9��M�٣��t�I��E�zo33W��0qbC2�^�@6���\�^+���M4�%�� � ;��ޟ}�yh]ۋ�&VgK�#��V�c�u��}��tkH	'���k�a�6afv�<ǜ^UIm٭�������|�%W��y�	>�8�WwR��I��S��I�v63�v��e&�l�l΄��n��we����<�,&���$fVn��q�^+k1��sy0�n4�D�Bg�:�\���.��E$�B'Qn�m��{3��R'Sf�)��+'�^l���ݻy#����n�Y�E���Q:��!Se�(Td�j"�����f�r�����4Ӱ*5U�TT�6�䰡���y�A5�ŨKRc�F����I�,hg4��5�A�>���8�Nr���O<M�՛��6m�q.	���e�&�k	v���hʺb�tiX PM&9��֩7k[ ���E�F2�f/�UL@5V��m�.�����<&GF[���clD���r�VO[�f.��{/��Խ�7e퍴�
��EZ�T�Vȭ���8��وAya�	n7.)��ms���B��\a��gڤ���Tq�b�����~��D�n�ц(��+q�L��/g[�[O	X��4�Jf�񟧗~9i�ʓ�Wd~�ާ3Af6/<U#,5T�϶9�ϒ�]�x]���o=�P�rpu��Zj����i�^+k1��G�t�\��a���3��^�1���P�$|9�ۑ����sM�M����,��Y#����ٻ��&����c��g���O��c�����PY���oЦ-��TE��4�,o$�$}I%*��������F��2NV�x����]�r��H�%.����}�����}����6�Mb�ے��W�tB����0��M�K�f�H�M�|���ý6�y.{��d\km!���嬌�4��U�WI��fei�V�=�o0���������Vw1��	=n�%9���1�'6r���Y��F�<�w���9��m9�YƱ�ٷ�>���:�[���s��@�5�_HwZD[1��M�>�
ϼ��w�ܱ��V�9��1�@�/���*�-�4v��CH�`�{^�!z��w}���uϵ-�mT��*3!3�ef?:�r�Z>H���|�ɦ=�:�����P<�k�S���
}��|ٛ�(_E)љk#wz=��������¶�4�(�Y^MI8��N�s]��.�KA��͗3Af6p�>��[�W�o��_�����|�^ĚL��n�n�������Aҝn)�mIs.V"ܥn�3�'�_~����"�$D��َ��L�[W��v[���<��p.Ȼ��ܤ_&�VmS��xٛ>�9�Hf�)�k#w{,���I�x�)���3#?K�-�ۘ������X�4@�(���{|�G����g�Tئ��"�+1��ݐ�$�a����Q�њ'����|�n�{�&H��3�d�sv�e��PY���|7>>�BGΈ��W}-K����'�n��0�>��ޗ��{&kj���zW��z�' >�n��f˄�I��$��u�.w�S�_s�D�{V3"T�ܵ��;=�ܻ��fG��8�:������=���jKf5!q�,qKB�뱛<BN c]��n��ļ``8���+�z6�ԊD������]$�e�٢�>�XM
�9 :��m�d��$Fq�f�6�`�p,^OZ��辸-+*���WPo>�r9�����M5�p�/�@��oJOQ#+:��:�"b�b�S�2�F�,��I�^dJG�� ����u��y��僝ضI��1���l��>�4�ǛYF���gf.�SPK�9l�o:]s��Z�^�p7ח��3|	Y����| Ƀy@���^tS��z���XTV�����K��'�>VRN>H��Ӧ\�?��!i
f�[���m^?�+��R $�'����u��4��v����-R����UD��^�֌�C��d�ӣIr�1�,bD�{���)��KbTpܵ��;��1��TG�p;��{3"�Z�1���vc·^�r���]���٣`�޿EؗVj��C��}��5Ni	�%m���S�n�].�wa�V����P`�]�ϥ8P|�JTޞѼ���k ���!"@�KĨ�k#w{,��n�h��:�R�ݠ7H@#��$�[\VB�n���@en�-�|�	��1��� n�{�u��������i���d�Vڻ�x{X��z���g���J�WU�>�t��n��{�s?ߚ0'�.��Jxw�v$��5n���m�n&،�~=��︶�ցh�⸍�gn���R��h�p�)�F��=mjf����m��n�p�G �-���]�f��c�i7y"�K�
^3��nE�&ؖ\��.�H�.��ε���=�Ю 3��#���oZ��P��ocf{t�9{ ��x��a.1M�B˗P���bS% �a�و;tu��lΙ�����lqo����-�K��ś\�a��Wk.��h���6e�T� ��/������G��Oi8H�Z�מ�NYj���|�u02,�14Ţ��3
I�G.���v=r���9�9,;��嬌�2ϒ!$|���7[��e�G���H����̃#�؋͑2ϒ���LePY���|7y)	޻�Q��X�m���N��3��9繵;�Uyo���
�F&��4Osm��g:IO����&补�j�2HR&��b>�f,�o4we��I��
�g4�{�'>o�"r�֌h�B�ɞ�P݈n��@/{]f � �k��Jf=�����Ӗ�����ٽ��&1PY�����٭/�S�>-��>s�G� ��������rjGXsm�Ah�Q�&i`�F�1� �`�Sq�nq���+�>ٿ�,���=�հ*�ZZ^KX������'ׯ]+�鏹�;��Yo�u.-G�.ݍ�eѶY���=� _ND�RZwj`���01���0�����#�"�p�H�a.�C]��D�K��� :N2�^��uq&��,���2�U'��y�mS�*�"D$�CA�cc|��L��GLn�NV�,�����o��$+>w}cA����x���9��z�F���d��{Zy�2���)��������O�~���?���ߟ�뽁9�[0��0���^�i��X��U�9�M�*��6*e�]��wN�-�W̫���utcg���p���\k��w�%&�}�`�PO�h�S������l������C�I�L!rҕ�fK�����ز�V��u�'����v�J�캵�:��~���4x~֖`ӎD�ɧ���s
f�	Em����]K�"��I�z��X��1S]�|��%����S�aœ�;�[0]���%<��ܟ$|�$|�J�h���X;y^��)�$�M��l�O�9)���خyu�~��z'�2��/���2l:l����n���v���qM�eԗVg#F4n�3�'�_����O~�I��vj)tl�g�n�d�?;�--���-��'�D �y�&r�/���[�h��;nķ^�Ӫ~�8�pGva��U�����zktr��}� H�@	%:�,���WswW/}XI�6ט٧Ϯ79��>��H����i9��{����f�	;I�7�9ڎڥ���멟G����ە��B���睬�Z�m�;��{�b {ئo��ڼ6f�F��g���kq�oҨ���@��hYg��0��g���{��Ìr�,O-���:������O�>	'	}g�|�^��B��u��#N��z�I8KZ���f!����IS�1������2V%���]@��Q�۫��'�z�\�?�%$�m,��\I��k�l������<�+d�h=�퐑	'	ZClvL�=s� v�;I�w����ڥ���u.<>I���\�_f,ů��H	'	�a�1��Fܧ]21d���|IH	$R;*k��J��^����RN.�wM�%�M�]�����ZE2��gX�!a	'�[�d]��_j�!K?#�� l�^���nĻjT�x�z�l3:۽�o{�F�:qۏ�~x<x��Ǐ<v�<x�ӧN�=�&zSZC	�Ln���?;E�������{=�d}�MF�-���$���}��k��P2t��|}���Ӵo��X^Ǿ0�>Hp͓l�������w{�x{9��a�׷��;�����$�d^��=^Bq��������h�ROFn�������=�o�.w%'�X����znj��y���Ӥɬ�3�-�`z�7����z��2���n�C�����m�UD�n��F=��jeh|�������x!���O��`��q5��G:�������K<:8<�C��p������c:����F6��V)�G���3c�j�!&�D)⠁������*�<�4wx/x���T����.ď���t�;�g�U�\P�hD:�|1{g�j/?=���RdjH���y
<4v���`��gH��P/�voF/i⳻�.d�S�w���L�8�w݂����"�"7��no�;�׀r�ߕ<luA���~�=���y��=�2̣6��{��:j��;��h�̿k���(�-�{�u�j(��_ݝ����b�b>���������f���WX��/V�1j�p{;�]�j�iL,�����3۾^�hw��W�3`���n:}2m�`;���K��f��R�CU��]�򲮤P9�qĊĎ>Okc��t[3��pw�7z.�wwE[�r���{:z<QI��G�^[���P>#@�W�(]��;��F�	\)���e�R���s+�X�T��ob~U�e}�x��Q�i,����&��/ p�Fi��r�2`��:�f�[���J�����z�g�d��Ezq�:y'��"�8�]%��u?7��HnQ#*���(�7K�9�N&�=�̶��igdKh�m�����Yi�9��m~��_{{\�6�[Z�h}l�^ѝ�M�9	Gެ�N����$d_Z�����H��Zy�f��h��͛+#,��:ڭ�m�m�n�N�d;"΍����C�-�cm�A�h��n��n$/l�;@��E�;M4Ͻ{ۍ��3ml�G&iLo�g/}o/7m��mų$7f�S����m|oXmi�������!�HT���8Rl�8w%�d���H���%��Vw������Z���'��eaJ�;���l��v��t�mn-�,ܜH+;(L�p���>S��h:E�n�ݹ�w�n�2$����$�f�	���':��96���[�"y��$ƴ��������nd����G9��Ŷ6��Ֆ;��P�[4����E��mk7-�i�G��q�nVhDR.Iώ�9�^���nN:"}��۞;ｉ���V���]m�L�-кڶݷ��q�j����[�s��
7;��ƙ׎ϫ��R�c�%�u3���جj�أ��Cؑ�6k];Z�����������lK�\�-�3x���]����fI�Inu��[=���Nۧa0`D�3���y���gJ�i�5����P�L�(���4s�-I�c��Y����/8��q�GEvD��c��Yx�2�yR:&%:�����m�X��K��͎�E]h+�ҕ۷:}۴4�!��v���;r��������nL�U�c@������װAb�^R�㫔�1+�� �v�EŉX�mwSGTҍ�i�3�a�I�.z^SvLñ��Nq��Y^���^0�)Kf����]�zmt�6<��^8��E�X�Cb��Ƶ���]���ǝ�V�`[/�;�/��6��d�u ����qQGj笜�܆]a;']r��J���Yy+��8�u��*\���Ѷ��%�Lİm6��yVy����b�A[��p���]S�����-���lA\k.f�u���4#J�Y�CH�ƘlMDX���c��f3	��;�a%�������)��n�g�$��n4�Z�b��][VM����a�!۝<#y���k56z�\�/#^i!��^5��e]�(JhF�hgK(T�J�Wm5]7sQ�]�:�WtVy����ѰX1ֶ[�<����N�����i�.�T�k�~���n����rn$��Ԝ��5�tܜ�v�3�m#�Zڨ`�N�\v���]b���{g��Q�Z���
���F���-�`꧇��\�n�S�'Z	�9�#�B˪�$�e�8,ͮ	M,(�F˨Mr@5��mV,xkm���F�l�\16�)M��Q˩�@��\@�[��Y��gi�l�l��\����V����Yp<��$�E�Y�Pk� p���W���bcM��}z��X�])V�,.5�g�cxq=]�q�bl�1���l��f\�&�y^�i��d�ۋ�����B�q6�9�B0�����[!q-�f�C�櫀�/����S����!s(�\N�:$�7��]������l6��-.g<��(=a��uV6k(h�ǭe+4�2�dT�ۚXώ�xC:�9�]nsr=��[�����%_�������3k�R�c���2��4�ҭSd��Q[MJo^�������ǧ�1�~������:V�ed�����.f�Ts��!V�H�BI�72�����%5�0�(>��~�]�}�s�����ٹ�%���%S��^l���Dμy��4$��.�:��b&�Km�\�����{���u0��EAI8�]���j}d����Ek��䏲g��n����b˦��7ڢ���7�����8�I$�o$�p�q���ӫ�~|��Ⱦ���U��l�2�:G�9Θ�թ��8���ܺ��i����v^�f�JҐ�X飲]&�����bKȕ�ሀ���$fw��uvŇ�Id�\�^�Uqzj���/d��<�p3�ws^>oG��j���e���{�q�����k����_i��M���y�@�5��ǸO�~�����G��1�=�i�|�����b�L�\�ĳ3_���_�� �=3�^�on1]�Gw��>IUN�d�zޱ�}�|�\���w�z�~e�yS3}��;��9����nwz�vn�ļ�!�{Nz��,��v�B3=�c{����Id�\�\�5ۦ3��
�7�O�J<�$�W5_;xD_b��gM��+�h����O�^������%��ev�U�]��݊2ؚin�Bm���bTf�
[���C�;���2yϘԠyRu;��}ʹ�ު��6o����O;����p?��%Q<d����zO�����S�_����l��x��qh�&�=�"��o����.�	'H��z||޹��0�X�lm��B���<ėd�ڂ�V3�����7&7(�ĬQ}�T �wȋ0'U39������|Ƣnn~*�a���U��U�4}��!"���OǪ���W����O�"�u;ׯ�ʹ��j��6o��'ʑ0H���J>PBI�Dy"[
ޝ{�J�]U۽��ňɴ�x�U6�"J����Dd�l��Ć,OD��2Re4��2��e�r�O���Hs�ns�H�����Jc̐��9o
���wQ����$��yhݾh��7�#e���p+�f��]�v�����Yُ�ҹ����7��s������]l�����w�R���9����0�;�-{�6�'��pj����z�}j��u�2[�:K���7����ݸ���x��{yt��{�~a���^oE�d,�Tn̤7�p��Xi�N4z{���H�E�+���}%扥i���+�e���<��̦{a�f�[�ȋϼ��W���>I8y�Ȼ��.d(��V��ϳs�s��U��6h� ns�#䯭�3	�0�&a�-�L$�� Q�����h����}hz�'b��v�`"��0N&s��I��i*��' >�7]�Ȼ1=��׼�b6�VO2[�����6߯��IH�?��;}%�E\�����"/�"7s��s.U�Wv��D����؃C�a�O�:�R>�@IF�����=N�Mj�"���[�6s���脈PRN8,�6mC�U%첫�D��z��hFU�����_ӛ��?? V�����\$|�	'	fjk�jIW	4w_��� ���nf\�M]��R!$�$�^o�s9�dp��2e�,�l��2$\Fc�7|y�v-����鿽׽)�b'K�>�f�$��{qy���Smo�SY�v����5�C�>z���kjKv���<+�,��f��f�m}�t�s=_����+� �w-v��:����i�ڔq�L̎���ĻkY���]/"�Vw�O=�m�4&흛:�G'�kv[�7<p��[t�\t �j����Y�ukq;S<4=7r�HrQv6��	��v�*�6.N��wC�:��5�q3@WZ�񣛒k�%��B`R�Y.fF��
<����kF&��?~��~Ե5)qk�w��n}��\i�i�%�\թ.�m&+�ƌ��޿��<|9�	'��׽���
��cf���3�I2I�Ӏnׅ_+��y�޷��nz�qpe�NHz��l+����#j�d�@r�E!I����뼌�U��t�	(�~z��j�y�e\X�̹V����R% ��H���zFc���o耒q�/�:/��+|�͸>`��<���kY;ʸ�w�x��f�2sa�Ir�rGF��Th��xJ�ִ#j�d�\K��	�k�^�v��V�������S������ͲcV�@�]4Tn�3�"5�1c��o[	$�:��G�˕i�pI���}މ3�!"��I8a������׃p��"��>0ʪ���	ѫ�E��b��r���!,j󉳵��l(��kZ�
K�Bb��Z� ]���;`A�<	�r��]�]��^��T��8�d�n�w�������	s���y���t|��B4��;U�aQ����w5�V�'��o%Ov}v}���v%^p�Q:�^}ҽ�Մ>N�C�#F�eʴ˸���d�ji�n]}��x�33]��ݿ��ɿ]�:p����M���ۃ{���l�Wg1�E����H����TyV��6	�fN�
?Ȕ �A�#�A�,��	q6��xC����wg�Ix���䔄��Z�f��#j���oY�~q��Px���2Ⱦ>v��g��\^�ѓf$Iѵg�i���G�˕i��/n?��y�2�!G����;_&�"`	�q�avEٻ��s3ٽ�`lo;�$���w*��2�>c?��9���Q�������q6�5����|�4&��CN
h��!��j�FTO���;ӶU���l����l���bK����w=:�`�9��I�W1���eZ��O�QO��LLސ2��7����ݺ\�j1����"m4��أFe�J��=�����p�����Ԧv�ٚ"�`�Èv��z��X�\5����yG)v�'��Y��1a	 RSۍ�̺�ẫ��l�'��'��l>�q�m�)�?�D���L��w5O��l'��hF�U�����E8�-dG��Xz�f{;R��P�Ìĳ�΀�!�\��'�D
[-�91�Jk�E7(��w��7_m��I?�):���hs�ޢ�>H���s����SWm�ٵp���m��Y�߯*�T�����\J��j�^���;�K���d��I���0e��2���e`��!�̷�l\F�,�4�^�D�G��������7��"5��E�N����ܗ�_1�ݶBv�,�+���D$BJ}4v*�Y�"���'���PbYV����f�L�PKz���\���#@`�K��]�;��P���n��!'���n8f]�M��	;d�ڈ��e��{�����f�D+t���>�O۸����
��ٍ��T3��YS�'D\�%�F��-���.�I�����J�16��X�z6�څmZY<U<���vE���:1�uG`ݛ)8����c.�&�7_�7���c�V�Խ9r��b'�?�N)��lh�n���}�8߫�����¥e�cf��;����C��X�i��:���s����1�D����g�c�Vq�yh/Vץcl���t�AP�&j�Z;�����v! Ǽ^=A��HI��o��ߙ�Y�\XP|�0�q�1� ���vո���g5�CvZ2�Im�tv���]Oc�B��n*���=rp���f���m�yx	�n��\!�v��g���k�����Pg�Nk��Sz��u��9�z��H�A�(m�6-os�!a48���ܹ��BJ��`���q���e�u�W%v&�b��܌���O߾�Ę�(�}O1�'����w���Ţ��6�5�Xh7J���O�����O�G�I�͜\(V����\
֭�4�%��n<�K��_���g��-��ۉ����wy5����xq $R\��C���ho����d�%�����{�6��	�����6���;v�G�IMR��~�f�s$��v�Eάpޏ]ǣ�ܜ\(N����\#�!&�~��77,𲮈H�	>$�Zf�L��w�ZAgl;���Ubn�e#䓄����g�Q�T2�Z^�6���DR�U#��-F�� �YXB��m�F��}�=y�s����R{��׭Xh�J�����;i�fɮ̹�H����W�y�Ye�gض�*�G��w�����q�	�<[�Vo�z���u�<0q��U:���t����_�e{e�:�:�&S�N�v�.q�'��K�Cy�
�3uy\o��?�%<�6h�vvM�˯fP��v�K	��۲�Xr���/�wx�u�¬����%>+D�)~`+"�� �X���	��}羾ˇ˻�輬�t����q�ID#��Ic�z��p�e8�%�<fq��Z&4���u� �=��R�M����Eh�_�N��R�D���`b]���k�&�ǒ3Ԡ���y5�9�sL�E`��{炙�?�b����'�=��_2��M��A�;n�}�8�˹��	$�	�����1v�V��k�
������}|�.�#
��F����w���ˉ�F�(?3c�˸�e���'���g����?;x��x��Ǐ<x�������?��������&5Y����K�uKN ��-�����C�b�{ܺ��v��X�.�{���������t��La-�E��x�<���\~�bO-���a1�Y�EwI)G��~�r�bY��b0i�<���eJz�ɇw "T�rp�R=�yc������`_Ix	�M���}�=�,h^`%o��&6���T���>X�h�z�x���7|_rcf���?F(��?s1#�޺zy)}�\�=
���㽕��율u\.�|�㔩���s�~������L�b��� ��{:	�?)�	�y��zp^��O��w�1>��>��q��O.���ޒ̽j%��|5Y�x`mS���0�����2�W��x'޾�<#���� �K*L���ۿu����nAkgם�<�=�|Ժ;���Y�w�Ki�=;�w4�槛j��^�x����yy� �=����F4y5��D\6=��w�������=�|��>"�,;����[�X��1?뽆��!��2ߩm���9Ol+@�}���8Ɂs`�K�~�f���'w{�xg�Q���0r결]�fE�0N9���{��U������x�y���lt～`)���<��ĩxӫH������s�=ٻ��	E�L擲D5k{�%L?#泼����j���庍[ֆl�%P��ǎ�׏*�ǖ��<�{z�{�n�T�a�l{}cS�Ql]8̞�t�v��yt�ᛎ6x;�h�x�:�~>�mwK���m1���{����.A��%����ﾎ��7�!B��YoYz_��ٚ�9�(�w��me�l��<�Z�;�����SdNp��i��z�<�|V��[c�F�!:{Zp�w��I�c0)���.[]����|�۶�,�ÂZ�E��^�NIy��8����\%yn�y���{ZM� �e�n�l��rvۉ�h8{^^���V�H����f��9ҒL�!dX�"���泱�/�i�G{Y�@A�L�ۚ˄�X}�r�+��kY��f�G	'hq���$��B�n��m`|g����'6���Nc��	3�{A�8��M�)Ay�	{bs�z�<�#��z�c,s;N�6��tp�Y�8���Gy��[���o=��v�mY�e�a�̆k;f"^�w�"%8IA@����m;kcV�!Kmζ���vv�-�[>�Yǵ���9if�j�RR����T�<�x���N_�Γ�**�m�z�?�G��
|�`�6P����a $\NP��}�W�q7_�+�a'5[���I�I?���b/:D�2�[/�ׯ����!���0������� %v�F� Z���q��2N�ݿc4�t,�e�q��8�bs\v�.���r��^5`DI)	��c�k8N�(���)�T!�an���{sӅqI;�$��U��6������}�['����j�'u��I�J�H�ٱ���؎��$R"<�%�Z�;b���2��wz�.�#
���Z�H�#��FfG`��3u,�m�#Թ�En�1ھ�
+1u�R�@;7{BH�]/V�)�*�NK����@͚���~�����N�'�,[㗽'G�yf�K,�5�8�c�e,̆ax�̸w0W�����9�G�7�R���0�t�X��X�݇|X��12���I8	K��a�)Ƽ0�eZ�_|������4v�h"��oo7�Uê7��y�<Ĵ�.��Zs�.)���w>��^��˻�¸'�!|}-O~���>	>H�]����N�W� =e\����p��QY��8Z��'ur�8����I�q�F#���P��Ǻ��F!��h�P�V���L���}H�$�"����9�^���$|�y��}�ξY�w��hz0X���p�~���I�{�qvBE$�lmƬ�'���Rr����]q�R��U��SGzx�Z���n\�;�s]����,�H�gyx�3�`�q���K	��D��f��ia�f$]�j��ݿy�X�K�FV!��犒�)IK��6������@� �ʞ�G�Z7�h�v���&;&�n�3�&��ܽ��;"�ڡ���l��l
��:�0\cs�Ы�1�\[B0�@���e�]؝��%�>�pP�vI_�zv�d諍��ɂ3�5Y�`��{R��כ�<.�=+�qgu�a��j��p�F��EV��v4�ί���?;�up�l%Xi�ݛ�#�}�����ʗ:��4�8���2��r�f�D2���2�ɻ��#����>�����ߑ��;Z�r12��s��!u��J��H���IN_��L�só�M���Nu��|���(��Z�J�a�4�27� +!"�s�	r̍�d�۵At�f��B��]q���ǱR�$�%,��<ӂ'_�t��q�gp����#.�K�ō�,볼��;��N'H��P�5�X-W�'\OR����ő��0�D\�H��D��L8%�͌Y��9a�/�Dz�+�t\v��q;���uc�XM�jWdvK��/�W_��\RN�V,m3��9��[���A7�2(���k��fVd����ʘ�z|��O�(�����&��Pn�z?�Л��z�߮�ҽ���pӽ��S��l+�=A�����?F茅�u�XZ���F#{� �m\�be�>mG�BIq�{)�öI}����H���G�w�~�f���^VdFV^E��z>���	�[뻡I�N��bL38��.bГȾ�W���NC��n3��;
jo[�\��kOz!�qپ�1K��	��I�o٦+[�HI�{4C�m\�be��I�)'Kw�f���/�3��<?3�6�!�lJI̽f�.u˄����H�A���0����w���9i�k�v�]���,x���F�G�L53Z{0h�\�ςH�y#�n��w�`�ԭ�x+����w��!MM��~˗��e�y����Tܵ�wgH�>>`�$E)��Lٽ����M]�V!�rh�������T�U�:���cY~�I���Mxs����aLՔ*��D�ѝg��Z�ʚZY���L;A��/�s���p�K=7v���e�F��ͥyOLN���	'U����ǉ��tk^�`����=>�;�<��!$BK�
͍�^���ƌ�57�����@ۻ�]�,�YҢs�2w&�����_��B6�	����v �Cnl�\2ʖat����(���w,a��G�->���"��n��K�����e�7;�8쀌*��@$|�T�G^��"��u��8�s[��[�vf:5��D`W/'�f����q�j�$�X���ʯ2$$��Qۭ��'��n�6$4��d)��]o�r��D$�"��`�Ք��7�"��s3�D�����j��W�I��d��q�a�1Z����sL��a5]OG�if�q=��W��*�8ྒྷW`u���*��4.C�5LV_�JD�p�F���#����wnٻ'�u;s�W����r�s[��[�vf:5�z>���(�+���-]����0an;��>��[��KQ)i�mL�8ۍ�fx��Aɪz�.wg�Iy��hDo��]ۋ�"��6���l)��\޷�޹׹���r �8	'^LBF�g���k����ޭxn����g'.q�xb>�BH��P,Oi�X�cѮv�O�'��J$_]�MU9�S�i[�ff:4go��H��뻏`��g:�dSx�s��O|�F�6������d����4F6���7g��y�ܔ�"������}�z��m^�Ս��x4L���>Sr�F�	'	G���f3	>�ꘪ��f�UY�!U88�3$c%�ǓC�݃K�*.��=U��ˠM]W�g?d������F���})8�p��`���Yp3M)�͗-����O"����6�9P��t].��v��ܩ�pn�}�Ϛ���a{{n�@���}v�q�����2��na`��A&S��˱Qd�c-5�ae�p�	f	G7�;�n<���=t�]������0���l�����c��C��Ѯ�R۬[�+��\On�<�=Ĝ�:D���t�gbF�ٸt�v�!�nm%>}���Ԯ���ʮ\�r��D�[Z;b�D�����a�h���������!����;[�J�Ofc� �����i����?���7��]�z@�.��fi�/$�ݍ�=��ѽ�_aEeb�~�6�?��w��XO-�p��n$�$|�-�w,z�&nr�)�]w�_��v�ه}���ʣD��!%�ê���g��T�םܤn�1����U��Lm�eמ�9�)"!%54ך2���}���nhk����uY�u�z|޹�f쀒��x[�������Igbm��9ŋ61rf�Q���q��Z�J5�l5p�L�����}]���E�_/y�ggnq����a�.pkW��w"��I<��މ��v��������=��=�TCRl7v8�.��^�;un{Cm	�;_�d"��TH��0�0=�qs�2�C�Z����P�1���/KC߽|�n�5�wi���z3�=ˏ@J&�r���r�Y�ut����Lep�x떍�a]�*�W\W�}9��p��R�H�k��5RЮvϏ�ſ����xk׻�f��ۜ�\��A��H.���G��Y� $�$BQ�La%���-�9�=�gd�w=y�Fv��	��H�%^q�Є1g^��O��*LQ��T�e#��ҡe�zzc���;i5P��&Gm`�5�$�	��8�tk����]q��O\<Wgg�MY$����7�L>���U;oT�7��8��f[U�9��.���IM��s��.P� _����$BW�vޯg^l3q�n_� 	o^Թyת��/�~��r����:��swm�u���*"�e�Sֳ���J�g��}�ͮsA(��ۆ�{h��s1������=������ٖ�d���?Cԗx|>�Y��qk*��w�Ux��8\]�m4����dV��S�>�����5���=i�����m�d%���D
I)�K�W<>���'��,�y���e�lA.��Y-���\�wU�����&� D��o ��A�a�L�")?�x�Rq��ݚ7sט�gC3�l)٭�&�����%C�L
c�&�ÿ��_������NX��:�U���~���p�㛼��*«��q��;�\}�aw}��>�a��B�]N@:�R����3���#䓀����IC;�4�{�ݥa����a��MWsט�g|�@^�G��j�R�9��M-5	S��ZcXԌ�jN.�$n�G.��ֵ��n�"�\�a1��ي/d�M�&��r$H��w'S��ǫ����_��dj�]���Yr�L��ӁjՋ��h݃v�.���$�ሤRP���!�c�ӇR[a�~��-����c��eP�3F�W�����.ի6�����,a��������H��d�guˊY��v����]��=�����H�$�cV<�~��M�6�z��F�
�sט�^z�D��p]}�Z9Ty���w@�>��"�?���u,э�L$O!�n�����v���Eݟ8�ff̋��z�Q�=>`y³��|�ݝ��	lf:3�#��y����,LVҊ���Y�$��I��zS���ȐZ2U������k��o�����ٝ۽����������"?�Q U��QA��s�c���!�����W��Yg�a�}.���1�1�1�1�1�1�1���1�1�#��#�##F(�����*F(�
� ����1�1�1���1�1�1�1���1��##�#####�1���1���1�1�1�1�1�0`F(��
�� �(���
�*A��1�1�1�1�1���1�1�1��c�#���#���b�`�`�`�b�`�`�`�b�b�|� "hb��1���1�1�1���1�1���0b�``�bb�`�b�b�`�`�`�����(�(� ��*F�(���$b`�``�b�b,bb�`�`��GT�L��L����Q�Q�A��H�������X���0@�A����Q����E��cc cccc#ccc`�B1F1X0Q� A�`{ (b�  �A� `��
�*��Y�@ �  � 1X1�(���CE�E�E�E�E�QiPX1X1DX0DX1DX0X1X0DX1DX0D]P�QQQQAQE�T`�0�`�0F�`���6���0`���0`��*A�4�#���###���9�?�́G���@Y� URH@�݅u���g���@�������������L��??��@q��X�����?Z?��~���?k�� ���A�_�������A_x�DV�x?������?�/���O���?Ј�*���@~����-"W���������� �������I�

�� A@	 D@DD@� 0  
D �  "#  	 "�@"	  � "� ��  ��@(�@PA@Q�	U5G�%��������* ��  " ��_��߳�~� s���Xx �&���Q U��z�������O�?��b�ԇ���_G�]��C��u�����pE U�H���P����Tk��7�AW� ���J�����tz

�_���G�A`h
 
��!�?��?�Q U��� ��w�������9��a��~�����4��*����?��?�" 
�����CA4R������O��é��?�}[����&�n(�*�� A��)���?^@��F/_��_Ԡ"
���������_��ß����)ޝ?�1AY&SYI\�c0ـpP��3'� b_�    
     �  AB�   
       
   
  X@
pt($ �

� *� R��UP��� U ���@H�@�( U@(y�H��	
�RB��B��
�T
��DE��R@U*��
P���"�U(R�  �   �RRU(���R�P�i����"��aҏ�����t�4N�p g�Ā�j�k��ɠ
aꪣ��y5�h<��(P'|    /�� _XU�h(( �x)T� @P�� �@ n�(�h@:� �9P� � �Ԁ��C��R�EPU/�  �(RA)@H)I*�	*�p ma� ��:݀��: Ҫ��!� �` �݀�� �+ �� Y��QQ�  >�G�`=��  � -a�(r�� r �ꠊ� �` ;� W; q@�DB���>  �I%*R)EDP�RK��q� ;�E�5C  �(�����vȻ��x�< � ��*��Q|  �y�2 j��J��u� 2�݀t-�8�+ $݃�;��� �$P*�|�P '�PH�@� *�H
��@�d���t�ݺQ���*�T��ɪ��wc�E��@3���M��
���)@((�   &�{��;� u;��8 -� w ��29� � S�k�@d� :�
�J��� @�RQJ�TUR ��R�	8��>��� � g�!��� 8�� ĢL � v�@
��  � t{� �:�X c� w`u@w`A� ��\ @��r d\�����E%Rz�A� S�a%%J@ h"~�U)�5P   �d�RTb0 �a)���E=A�` �QS�UDQ�2�?���������$���l�W��A��Q�����4����  BI�Vn�� �	&�		!!� �XO� @���		!!�����_���j��w�>�7��!��r��Bv��9q���Z��wi;��w��v��d׻��?��Bs�.���K���
����k��4]��x6.��S;tST[x�ӧ�=sn��ԋ�	ġ�8�{�5`�����1�Z�/��`�c�q���Wj�l�����C{pA����	՚)݃�����ޗj�q1:��o�6S{a�J3���R���!�[Ea�]��nst�81�2��e���v2���� �/Y����$���P��$\�TUde����>	sKGMb�������1o�9����T��F5����<חxf�jL��wOGu��b��usW�f�Ʉ��x�8�A�	7�q閬JN�Z���huv�5����ۛ�8�z�-=��-b��·&��Gӡ�P2U㣺���i�h[.%bִ�Ï%�Z�pbٶ�!(��i`:os�� �`;��_>�g�ǩ:V�8L��A%Ա@d�ڴZ���m�Yx�V&��R�`/9�YQ�3�Ka���+�&)#�gKo��f�����rr鼴LVכ���I�;By�g7���ӥ��P�
aoN���]����E�F;�xg��ve�by7�G^ׅ��8WW�8+���C ��ذSÆ�I�v�w�^	���/�*H��m��h�m!��L ��o��e{v��{�ME�=w�H�����.��laO�H8 ;�$�� 5��SГ�$�M�Q��c�6��Nɼ��/G3�*[�l�w�Lcuj�p��3^���ߤ�)����^C����fv򈦱J��GL�.:�.�����[ݐEß9��wb���ǀV���Ǭ��P�[3`����h�O�}/S�$y�0V����mH���+y�؎��k�8=Y���WBn��ԴK���6<|�T�ٔ<J��˲{4�{ys�nT�@��NE�Dg!j�c�{(�^��}�_6�Z�[�ed��x�)!��Y�4%�L"ȷ����Y��:���Hp��V.�U�u�"F�a�3@��ez³�$Z��jÄ��Z;N��1nRR�h�E�� ��N&�)"E�KJ\�y�=��#�}�l=~�[��>�vc��+�v�2څ�����'`ͨE"��&l��F���"(��z�(^�=�p���i�q.++ٓ[�P�1ݹ�వzՂ�����9g.Q\�*u�.�䆰���{�r�ؖ#�����|��N�
3g,��x���'nh-�>������;� F��Z6�  h9����J]��N���ʝo,�X��:�47{�/qS
�3Gצ!OKs�����f�٩4l�������y�n���ٛ;N��ܲ�s�n�� �u��ܐ���;#[3xړ��hPP ;'r���� �e�j�f��\�|Q�B�ª��\0+�q=У�	����h��z��;+4<߇W�G�i�X!h5�#_�f��#ؙ�����laY"X7�4�{�/ɹ��d�]
wk��# R�}�4㯏 uB.���Z���Ȉ:�6f�GB�'B�����0�.jw�d[A<������z�b�=Y��u�4K����4I{�"Vp<	-ks/�	�$B\|{-�y�	�h��b�'9ooC�s���Mnh|5��b�Ì]�=��)���vh����Y$�zB/��
��T���}Ѻ5>7�LWP�V�$;V͝.!3�%�rx�>��E�4���47�k�3���ۤ�w[뎭�:�7�=L��î���{�k+HT^���T��dy�m<G�z�%���QΔ6=;�3Ҍ�;
*bhf��ZHxr<L�Rק�������3O)�>�͡���6],�'Z��uvw��Ǣ̏��B����SQ.�ɉ��!S����Q�������󰱻���!���g5Jg;3N'�ؕF��ڎ�Kכˮ���g@��)�r��Y�����nyŜ���>)�aD�-B@��WF��9������9���zJ�D�踎-�ʒ���Ŝƈ�,��R��;�L�k�g\9{\-�����1��^�^�&�f��\�
�Y�Ա�n�&��̡�fTd���Wl݉���G�k�U��LF�g�#�s�&qy��~�i��^jb[;Bj9�gp��K��x`�s�̩�oM8&Mm������N_�Λ��.>���Z,��`p�3��Z��8��Y-��O���|b�|�Ȧ�ݚc����4@�6猒��K"K�])E7L�7�fc�k�V	\��������
a�>�����N�v��\���Pިf�:�[7zd��Z�u}�&��N����c�KGb`[��m�ײH���٩�-�_a=����e�,%0MC�w���<�:��ud�*kz#;��k�N��`��ѝ\�ӤDB�&^�� ��7�9�h�Y�3_P��������᝕���p��x���v�Z�JP�E  �k9]2퇻@��d�4�s�yS��eU�$���4u��}T|4XF�~����ol�eMz�|y+��4�ۗp9���@4f�N�0�wl5�@�k(�u���#���Y��q�I���|�	-�G)#m:n>`���{^!��nt��3
A���A� ɇi�93����R5:��Rݼ�h�}�(�,��y�zi�ݭ,I�3-�,��o�<�%]��7>7�P`i�h��0Eۓ�rH`�f�Oh3v�{��yi[4�ú���C��Y�H!��N�(����7}��<�W�n�s�rNS^.��晧.Ʋ��ܰ�twI��5t��G׻�&�Cx�^wKgj-rJ{���,=zC;p���t��^v�Ao8�'�u-��<v����QP��iAn	��ʹBӫ�v�od��;'���.:]_i�����tKzY.!n�.������ýJbU�
+�p٭r��Ղ�Mn�5�Y#
	`Tp����0}Τ�AS��1����a,���\��htQԬV|�	<�
���_ţ�[�Ó8�"O�7���	��l����Žb^��ca�	��Ճ6��-y׳��,�R�w��0��"rh�
jؤ�H-��
%�3�3&�޺���pSLӝ�fk�
���oI�+w4����K�[����c��j3N��v�6�,���:�vC�qx�-�&���'L}�n�l��;���9.�����w�o���G��	0��#9�0<J	z� �yD80�"a�:EO���`��2^���]$^{���n�%�VKG��@��-�4�혋d�blᴬx�㜛��l�o�x�u���*V��4�&��w6(:+Z_�k Jԑf�ƶ�+1�"��t麁�Yɺ����M8��r�{��0M].s'�noQp"9��_nԙx��8
���ۉ��p:����U��e'tNx�D�Yz@'9�^-}�q����:G1�eZ��tZ�Hc�x�M]4v����^摴|��ξ�"�,��݅��m��6��銳�� �;��~4h}ٷ
DL[�(��P�f��˦���&�e.E�.�9"u'��ѻ����ÂJ�p5:c�k:�U�w\��j�n�:Y�ާ7#�nְ���7y�ɨ���+�	��w;uEgc��dPr<���gB^�d�!`t赫7ޣ6Q�\���n��4�N��ucS�0r��mk%L@Z��O(�J��pr�8�t��0��|�еc��8�����B�8,��4q�S �-�fCRF56�����6.W�/w�,�§c����yIZ���9Et���n��/[]�碋�{�)'k��;�sm����r&n�D��re�+�aFcR�v�4��a�QQn�y���[�M|���|�X�����ʰ`(Lݐ���ٮ���&��%Ù6�p���\Ι�poB�+ɒ�=w8ī�ۋ�xqQ�l�r)�ד�aY��Yj.;&+�K!.�S0� t��S����ykͺ�=ފ4gY�vի��?�M��R�J����L��eQ9*��d�ppSU+#�ytש�#~�"��A��1=�^��؈�]0��BK�aKT�u���
'e۩��q�֗�F��M���I� hpp^�,A�f�^p� 6rFpٙx�!,Sv�oe�%�p�����apnda>�U��,�6n�9�'�T$��˱��6�s
N�T��.w(��o<vB�|G�
s{�L3}���gQ�ʞ.a�V	�ÙpN+�I�]���1��"��^���V����&�v�����9+��dZS�H�)������X{r���y�Ϊw:@�N���Y��?r�]ra*�[�t�#�l­�Ʀ	},�2���J��i�3F�6��TvQ��g!�ٹ F�z�l8��\��8����_Q��:�X\2�Xl9��ؤ�#kj�s_,�M��i:(��y���8:lu��E�v���b�A0�����Ջf�y���`�s#^�
� �X����ϻ�}Kq�SV;X��5��ڎB7"8�eh�'4�Y�������>����S�ޤ�lv� ��'�S���`�	y�r���p,�q5׹`�Ow>\u��-�*�TaԖ��nN�Wt�װ�����B
�����q�)����.��-����<���ۓI�i]
�1Xz�.c��%;!�+o�SP9�d��7��	oY��V͇y���cWN��:�f&�:+xo\W!`%�$�
���@��I^,���j���%��'J4;�7���67�:p��8p�btpf5Ĉx�ˎ.�\�WJ5�&�C�w/p��n���e}6<��6�vr����F���7�v��;u`!+ֿ�g,�iCk��Y���z�8�j�kK���l;�]�4�{����f�H�2&�@����٦s�z̝�7yܚ��Y�P���J5�wv�T.��G[�{8����%�i<L@j��6���HmB�2�:+��Bg+�H�CJ圱v(nD1�8G%�M��&��1��5�Y^���58��̙�G���[h�oGu��Է
�2B�Q�z��"=�:f��s��3���hn�B����6����@�n�R���twd#:�(�,��}����^�j�'��Y�.�6�b��I������EkggL`�M��h�8 K8k�����QVS���ƞ5w���X�ۚ`�������v�y/zZ)�:vN��YaքVi:���5�˴�Unry����&ȣ��'��7�M�"�e��[Yق`���t�+����w�Î�F9�X�T��t��~��(HfLFQ�r���-���W�M�(�B+�\Թ,UH�(���4`��qӊ����ck�����3V�X�zBj�EFJg}NF���d�ymgoR܎�kR�u��9�X�]�i�e�ǣp��f��\��&�\��d�U[vږY^��<��p����(@�ݱp�hl�dMN%&h,7,c4�֢��߃ڣ���Q��~5C�o#7��l�,�F���Ac�`��a�u�b�*��$��8"�7f��L�9,ˌ�M�Z[r^c�
QXj�!f����岂��.���T���+$m ��F��rdZ�Z8n�ě���� 4����cW��z�2���8�AR;��+�e�y�M�eP1W�Ƴxϐ{�\V�Gk,���ׯ�:�sG��|�;f�d�Rt�1��9���t�8g�Mu�R���Kj��ش^��V;E�%&��#0�O�L��p������q;Ic�m��e��μ\4wi�IK��=A�n��¦��:1!����0���J����l���ѭ�7z,�zR �l��5�Vr� f��4`l-�,���S�K���:��Ze�F�j���=�wK�k6��Xk9vtټ�8,�z�E�%p��b������Wkz�0���6�څ��kq[Kd9\��&&�脼�F�)�.%`
��IC������'�1�sm'`ޝ��栞�E�ON�*����v�ΰ��PS�E��;k��#�+E[�Q*`�e�xת.VV�ļrK���`Ku�g�����C;j�L�w.[�Y�d+��M�.6t>= [I+�ή{���LF�����L����/{Vv�M�A�s�)%ݹV���L��%9��7f�FxQ�,� ��택CP�O&,+.=,L��j�9bSa�n��t�����Y���r�����$��?�*s�+�Kq�^���%{��=�L�U�o1u�v=ئ�^{]�uNk�2'��;�k�P��_!���l9a&d<[���n�:#�]W��t%�Dˁ0@<�Ypd����}�[�=J��z�uH��@yn��-��`��Ԫ��|���'gbV^��yҦ�B]�-q����])IZ,H���b���G7;�]�R����.�v��7��ay��f��+����r��e{�n�\$ �� �vZ*��mH>�
���,Z���Y��c���9�E�X�T-�8���#��%���'��`��/��q?�a��D7:f���MҨF��Fp��u���!dc�B�B��E)Nm��Q��}� a! "� ��PAIa Y,��Y@Y$ (�$�XB,!) $�"�"�d @�	"�Yd
B "�$�I,�E�Y$�PWwquEwq�uuGH�,"�B(H

I �$� �)$�I"�
E��$@XB�E�P�I"�� $P����HX!"�H�	I�E $a IY$Y$�) @	 �E��,� �@R ��� ,��H�!$�����:����:�:��.��, Y ���, Y$��O��		!!�@�x�s��;���`ш�1��l��;:��Dզ_��A�bű>��^��+>߫�|��λW��;��y��P����vc,�|(��(�|�Z!��.���0�'����<߰NYckAA� ��D�%���O^N����ܤL윹�0.wf�>���&l����p��o{���i�c�<�f�.o��Vq��&��[�Q����(����M��Z�qNW^y�ě���q}�W�а��K{�JY�LU��c1�ջ��,�z�9�LE;����K�"�������ѥa���0�h�R��>��}��<n�S��d�z4kD����疷�ض?`�.vS��籺����@^˭I�*����0�b��|{<��Y�;�,+�]�gz�!�>{�R8�"nc7 1��I���T`���q�����q/Oj<-��W7=����,>ޝ�7z�ԕ�	�#�;�6�<P�S^���g:p��n���"l�M8ʆ���K�Eu�75��"��v$�oQ��nlHz�MYǻ[vVh�3v�~��f�`�b�����7��G�4{�G×m��SvH5��*��m�;K�w#ut&�(�l*(�l���H{�5�]��ћ�v����+op?�׸(��&�>Y�{<}"$a�gzi�O\�z�y����aHW������f�Q��j�8=KL�zx-��ފvgQ��~��������\ߋ���kQ0���.v���gBx�|�s
בz�&s"W����8>K�}Hٯf�}��黋4��ԏN~/&j�`�������팛jR���k�t����N��Y���-f��י�vj[QrgҪ�ơZ�TP`���812�8���U>�\��P��03����2�Rܾ����@k��1z�0	��{������~��k>�G#���HgnEp�*}u@y�w�{���L:��T�wq��'�y��.&��R��N��q'f��"��cP�y/Z�H�����zm/�Y��K�p�߇�4= �dy�źpg��;X�*��/�ƙ� -��k�������,�<W�$�-D�wV��o� m����;བྷ*��L)vI(�дI��(�m��g`ZsS����i��[:f۲���-���g6�e�!X�^�r�plL
t��Mn��7z�����
Z}�z{��!�+��	�9����x����Tk��9�5�D�E�PIڦ�{s����jt��;��z���m�x�j�N���	�Ả��N����;����ה�n;�ܟ��;���n���09�*��<~`�����b\_�sCq� �Ǿ�|�On�j�qZ��s����#��>	�O{�"7�yo�p�x�o
�����I����J����x�d��˔��0�B��W�w��<��[�W�S�]ƹ�����un>~�ٍ����m'�{���k��p4 �{�1�2���g��?PV���7�z\�����Z��<�e�%�g�q6��X��h�;����)��"�f��Z��A���C#-12/K �Y��^�ӥ�ν4�wo�PC����/��5��w��r����fw��Z��[jS��vh|��M[�0ޑzqy�^�<;�Wd\K��F��J�:/e�4�w/<����U2������+<��n��"P�B�KC��Vm�� m^þ��쾹�Y��m��;�d�!�K�1��
*r��r��qV�TH�E76�nb,����!���+ijU6�E�O���nm�ś�M�v9!]Ne�8�VI^]��s�׾���	���Qn�cA6ڑH��������ئ�&NH,�������>���҇/S�c����`̹�߼f�;I�ݥz&H�z9�O�%TW
�y���R�L坯�8F���-���B�;�ۣR���ŏm����9�- =�Z� �ŝ�ej�r�+K�<�wd����{�Y�c�2��IȲ�g�����{�S���KU7��h>�7Y�=��޽v�c;m��'.~8�M(�o=~����<���`l��`���Ҕ�r����[��SA�Sԝml�'�)��tPO�K=��7��x��r��}{~o���׬��3��mg;P�x�>��=��.���_g��}8��{������M 7��U���ݻ�9�e��qp�˓�P��e]����J��ȃ4#T^�x����=$�uk� �?<�
�n��)�o;�q��q�����N�F�Rnwn/oJr��s�Os��ӊ]���.�cAhd
�q�v�	�h)n����R��I>��W�J"�60��D��p=�s�|4j�"��Ǔ�2�=�Uf�<Ӡ�ɔ�V��M��pCz��{�b�9��}5���3����Ub`"]C�`!9��jb��B���x��HZB�:�Ã����	��7�P�;��w$�/��{��qx55����6����c���i���ow���`n��	Ǣ�`+��HꞆ�cgwK�
<������Zؤ���GA���ʧ��7�"~�廝�|R��t,G{�}o)��O���Chgh���F��;ʹ	�}��n�I��d=hW5w�܅�z���{X#'���9'\~�8��P��=��;XI���~�뒓��u�z�,��{|P��'�z2��u
�֖�<N	;�#P��ǖjj������F^���W���_DJ�n+�`�t�z�����Is���w�����'/gg��.���Ӽx$�����ow;���v0���v�� �z�H"jFRyv�@�/�+�g����#�����-���im�� �rv�b�o���L}5tz��8�̌�^f�3��c'q��xC�#ٳ���``G����!=�|�=��Լ�^���N,���t�S�����N�i�dIx�W�$�~�\Ń�g�Q�z6B-R����xewդ��vR�]K|J�M�A��l���/+h�J&t�/q+�)KR5��{:2�E]�;QMn�ݕ��;d�����=���!.��s}y��C\X�|ݏ^¶���b>;�;�u/��9�O�pP25���o�9���7:x���;n�}��7�?u��ݕ�6�:�X�dԍ�wv�ĥ�R�������U=��*W����~��Exy۲����Y�ޯ#f���J2gQ��.���=��	r�۽� �gd՛����%;��vq5��J �q��~�D�=����%�TD�ԱV��!���KCwt��7Q"�{p׏�n��/�N��}�_i9��XJ'V���]��abv,�?l��c�ul5��t�{��xTri�Q����7{���Q�n�]^���hB��c�|qR7��X^��N=s��-� s���\yչ���<�ه����l=$����
�{!�x9��w����Fuć�JF���97�={Er�7޾?6�!䳄���}��Ӄ��nt�+ӳ�J�z�8��os�se�-��C��I��;u�[��>gz�6tI���(��7(����>��5p3��~*Ϛ��u���;�ۺt����+�,O�(�P�$�IE�쭝8Xի�ezK�I�ϰ��׍j�<�=:���\��z��r�	蛙u��볘�M׺��v�Ի�\� ��E�)��].V��'w>6u�ŋ6$��6���M��7�֪���/!鉎U��j�f,X�u,�b�J$&H�Y5:�����n�oc��s��V},��o�h�2���;���'�nyk�V��N��Fױ�ьG��ދ�g6=�B
k��eEv��8��{�J�Ԛ>v�(���`>���{c�o�׾~��9s�M�[�}>�5��4�xƮ�]��2�V�yu��k)K��_W�NQ}��'e�9yP�ٹ&�E�ۓ3����3(ӽ�)��Մz7�TnA������p�'X�bF���RG�u�ӌ�X'�*�.�H1�L4̪��7O)���-h����_W�g����v�<�`a��w7�7���=ɂ:r����n��o���+�;�׺�ǰ9 :�g'�y�݋�Y#�x��龮��ܽ�V�硫�I� v�ܼΉ3�	�I+60��Pל�T1�滕��Ùվ^=������c�v9��M����ˏ#�x>}�\'G�x� ���wҌc\d-n��;*'1�pi��tL�Y��^�L[�k�s>�Z�]�[�]����5Ip�wJ̝n�K��Z�F3r�1)��R��7k �2�"w��y���ӝ@Nx�uw|�#��ܮ#D>�wכ�d�V-8S�>�j��������y:�{��`Mlz9d��!�㗦v1����jT��έ����w{�6F�|͒�j��@�L�-4h��`�૸����%��ɫ�3"���$'5��Q�m�zh]>���x;9������z{�Xjû(���i�;�"T0A���/x	���V�@�"�p�V=���47{�Y�Y�����[�;�n�j���o��NC���k�_c��X�ɋN>>�"|��7����[phl)�9cuў���S����y��U���lE9�z�w�xY��.����V{��U&wy�zN8�S���g9ۖs���}g��>HK��;=�w�<Hk�[�:�@k�!.��^?��k�S��*��S��8��7a3��g�}p؃��on_f��q����Vڌ.�"bf*.���K��G�u[�3x?�NM3�yT���{��3rg{��;�M�'XK����MA����<Q�"&��HR6�c��<G}֙�^~��Y��В�w���g|[{C
����yp��ȷo�x�K}䳂zS�յV������n�w��m}��eШ2J�,�����tT(�����s�tf�̩3K$EP���1V�ѫdM�\��:�^��ܜ��)�B������p �%G�&<D�)Π߷=�t���m
Н��w��=}�+'%�=�i�l�9� �;JM��ź�Z�_l,.�z����?]}a>�^S�Oo���ucQ���$����\ͻ^�zv�se���6���MI�暹����IF�d�k�Բڷ(��aK%�^�\9ڇ��!�#|����O�oNo=��9"��|9��{7}Z|�^r�:��Nܔ�1���
����l���1%��
�Я��S��v��*v�q�2o/%��K����[Ҿc���T #�9
��n�c�=����G��g ��U���f����M����$J�v*�l4�DF���6j���?z�t{נpE6�MS�x��U��	�/t^P����]9=� ��+���@>��޾gܳ�&�^����t`�o����qt��ݘ�� [��a�^s��=�3.�1�.�bO(���"bԖ�^��������7\N�'�7��hؖ-�V�f��[l��C���F��}6����'���6��V>��;%i��Vw���^���}��7�D�˰d������)Ҭ��tS�8��kD~>~�ҿy���Jk ���'�il�͞��I|�����Ǆy�q�ȑ_{�����QH�U���6��3btBܺ2��ߠ�p�E���^1|� .�x�5����.y�p^~s��]�n�"��+J}1=��+�K���?q��T~gF�,�� �&9�Ⱦ6�{7���9�΋�r�.��F���C�W��1P�u����,E���@��6�拌�|wޔ�2�����0Զh^��vS�s{=i��#fFׯnUV�zimŶ���UD3v�7_!�W�<+�^�,T�@�[^W�̛�r��u�Px]���ك+�,:�ۼV{�v�H�������x��������k��9
�<w���h��B[��'Z��[��&���Qu�}٫N�U>�+.������r���c�C._f�x:�������K��VFVoGV5�㫢F�|�Oz8�p���=�f���3�����I�u{��~�J�wۮW�O�#�{��tCGǀ�_{8���
�p�{a^��P,akkסW�g����Wx�������D7&I����c3.�+u�%xg��KE�՚�x��Ԣ�P����|l�[���=�[s��^y�o$ϱz�wpnxnu�k�\~��)�D��ᕀ�g/�������s�O��x{�LtpR,����d'�+��(u�yt��dy�	y|9��u��D�j�JT�A;�m�Ĺ$�wOy�e1o�	<sDՆ���I��y^��ak�}����G�MQ�&�4{5=Şի�|{�����Y_&�kZw����l�	�6#C ��xȘ��=�\zn6xI��b�����\�V�@�m�b���/Y8wU(��ٌ����<w�����I����8�G-�	�rhXtn��"6�0R�99,׺�7s�΃��b�� εv#w���q��v�T����ב���<�F�c�1э�9󹜖��qg �,D)��{7�y��xLu���^�ȚvI<��ݴ4�����sLl�G{=���8��M�weJ�"}Ƿ/�#ƞ�|r3,�+��ީ�ڼy$��j�����f����33A}�I�%$x-�LD�FRE]+u�w�@ˀhU��n��&䠠���)P���=m�W������>���n8��rݮg�ٱ�N-�^Ż�r�m9�ia�0g��e>'!Sא7;���6�`�����/��&�ĵk���ͣ�h��d��q,�*A��.hIc�\q��P����Ӛ��,βOZ�{w��QD7��Q��G����GW[�v����H-�`/��a�A��ˑ/1�~\ޕA��3����u�{���`;�P�ے	=���x�~Y�A/�������#���^n�?[��p��݃i��Ce�N���>r�޴*�"j^m\���g�K��Z����7�����<=�h  .^#���q��-�aC�1���F���wd��gt�E���v)�4�C4�0mFe͵�#:4!�ZMI�rt=D�����U
z^���
X�&K�!,��K�.�6�av�h]�a�7�#f݇]p��z-����#�����Nu��=�FӜuX!��d���䳽�h�ݜ�-�ޮ;8��5�\k�B�ܛ�k��)85�Kz�u�Ъ4�D�i�1Ż	l���#�����a^a&�B����&5�Y��J�kk�:��Vݶc��l����.�$�`P,[��m���lчZ��Dƀ�W��@�t�S��5��0Yra5'��F�gX�&-�2m��rk5��)�9C�dZ��ǃ���Yv1�]�4.*kq`�X�z�츦�\���N�ͳ��m�i�jh�nlv���g�e�[����[׶ϬSv�a]|�]o��k�IIl�Y��q�v^LZ�+��qAX3�9n}�]�s=��Q6�7J7.�m���I��i�3c�۴@V�1�j�t��Q��MhZ��� ݸ#I���y�n�,ۮ&��V�J6�F;xn����-ωnӶ��3�psu���t�>�X�{{;���0�u�b��Ĭ�� Kh���f�Q��%MNR ����4$m���i|f��z;n����W]��-��o+�@v�+��p�kk\GZ=�]\��Y�;6��N�o�iź���053�����)u��`�t��1ٰ�d.���=]�z��&ܧ:k�&;R3�8��V4r�z�:�e���션v2��˳G�O��gB=J�0�)e��L���[�+ʺD-֞�h�
5�;`� ^2�C�&n�!�Y��X�x��3ݧ[��6��uH]m���(���#�]#i�䴛�c���:�
���nrm�^Qu�Ì�p��cW��H8�V|K���6�|�s��ǰ+G��uN���5�)��.;؊`�!��mf�4�(if�F�,l#��ݴu��ᅭ؋s�4	�´�h�j�;+��o�1c���+j��H_/�û�8����лc���Q�e��"F]+nԵ Vae�Qv�+K����O)kَ�����ƍ	���8z�^��!��O^�����֔S.ۈ�s��@�۞3��V�7�Ξ�H���
|�лbe�¾u��5�f�@��m�\:�	\q9���9��5�m=5�6��Э��6����"� �n�'8�p��+X

1�;c���[�ݽ����n�I��>��;�s�;/Gvn�������1R���ї�E�IR�$TYI�����d�ND�a����箱l�:�eƀ�7NNr�TG8��X7!�0�ᵉ�7��1�K-�S8Gk��6��5�jx�6�j�,틶��vݬ&�J�e+HG�˘Thԃi�Ɨ�R��t 6kB4�h!�ζ�q	,chm]i
S�t�^�`+-��e�[l�RU��q����<�A1q6ͼn��	ܤ��.������6��ag���g���M�$۞ݳ#]���hn�c4�9�Z�̌C��k��'OA�ݍ��k�<�B���6�(��=k�s��`�"c�y�6{\�n:^��DR��X9{��y���tpr���<�O>d��qh�Bj�Z�+D��P�8.zj��u����Wჭf�$%���Y�@��$\�Mm�Z�Ƭ(�y��ݳ�fH���z�a|������ݷ%���l����x�� V��tnى,�\M1�hu��PVX�Ol�qc��3n�����Qf��^e2��r�,�Hq����%�z�������*��v!�<��q�DWt�}�ck�:�5v�rv�f.ݜ����:h�5��\�C�N�6��]\=+��S��l%ۮ�:N�Nv� Q-n�u
.Hi���F��q��`�Ng�1>��j1kK)6r[�	h���Y�`d�MLaʗUq��������b[��ڀ�7�Z.�XD�t!�u�ێ::�
y�!f㕅y���K�^�-�[V�&n;D���Z�����ͯu��h�n�^c����0��Ų�^N�dhx�k�Ӓ3;���i��]e�i`M�Q�Y�z�E�0�0�<���ќ�n4W=[<�Zܖ4��{]�n�c�&%��9Д]q	pMtu�V�cny�eςMҭ�NėWQ�S��,L;�۫F��ܚW�GS�xZ�dm
�M�M�pv���X9�,!��g�p�mIH͌�]�lh\��.�Hy��˫��k�n�mZ�GQ���4%`���b� �o"u�t��܆����/���]b=S�\m[�����/����o
�M�<!1xB�v�3A�G���f9��θ�.�8)�*#���i��v5R9���$zͨ�w[Y�!V�[[��ַ��c>Nқ��B�y]�CF�1���fC�3�������jWE��MjE�sm.� vq)�`��SX�lbPm��{VD�Fx���8���R1�m�+t��%r���`WJ]�k��=�ưr^��� ��M�V�����D��s���:˘�!^�¸�Z�����1�����|�9շd�C�yԻ	�D��ܝ� w]4I`����x�,�͡�]m��4ԇm���'E�z�/b;���,<��$]\�x|�'Y�O:�׀�N4Yl6[��-����Ը��yU�V1��)�@�\���i}�=C�,p�g/	e�.��PXP�B��ԗ7g<�4�	ۄ���8�m���v�Ʉ���R�<Y��4��a.�������r�uƑ��|�|�|�qyŏ[b����}mT]7`c�<�p<��_%�󙸸{{jn9��}[+����ҹ6�q�m����oi���*V�`Yk�\�q3�V���5v�5�9�s��
�MqiewP�hbR��<��c/;������89-n	�d.�K�m�����4ڽBSs�%�p�ZV��=��H/m� �:��:�ݮ����Cn��8����h�
\Ґ9K{j#]�'a�'CWQ�s�6;zF��4Zm{���7)����t�����D��x��i�˶�ДUs��[����]n�ngPr��籐����z�kf��%�B
i�*�1(� �=��r�Y��P��j�{\j���H�`���;�Q˝ַn�/##�kn[�ٺ��;s�N�H�C����[�ρ���LW�G��|1Dq�a�T�6���6;'OO^�(ƭ�UZ���a�q���#bW��۞��\��t�s�� �G@���m��f�\xrn+q��Ƕ�ݭĐ����G��H���{R�CK6�Y�փ a�u�J�Br����ݜ%F8�/jM@�&��-����C��R����݀v��[���nnv�[�89;��"��K<;���5j�s��9�k�5�r)u
��m�hg����� �ql'��(`;*n.�6�t��vM�q�6z���r���WA��<�;[1K����C:�v�[��]si����3�}O"��0�<r��b�"sΪ	`L5�Vwg�.;Z���w�m�H���=�j�n�s�l\�v�cj# �3�f>n͹��st69.��A@z-a��C�`j�/F�n�Jjn:����f�)3N&5Hl�$&׭�;`����kas�g�#T�k<�v�7<Y�����g "k&��3)5`B8��X��`דs���ۉ�W���f1͎�l8Szz��\LL&
�(;�c��]s�w0��Q��aK��c1��eCH�6��4b�ٔg��_;��*���Tmm�:�����3u<�]g����t�'˃��ٮ���M5.��aB�,v�Z	-���j�� ����U�M�d.�4�6�*�,��E���[��b;5�;mk�9�*�K-��v%&�=�����9枩�k7c7d�[����ū��)Z��y#B�
W��0����<jeb�ŕ�l�� ���6� ϭ�'k[ZgK�O#�����ލ����q�V{�6�>n9�l.:�l�5�u�7:�Ĺ�Q�4�wd\@�P#�c��<�6�:�!�N`x\2��b�l��Z�:�����x�v9��:�*L{�k��m��e�ob��6XP���#)[(c���:R6��z�$�Ʊa�
B��6(�[+Q&���ʺ�P��v��a����cP���ZLхf�c#a6nw=l�>�P��u�E��J�ݎ������=�P�6�α��y��g�]vUG(�X�4^m˪]x��R�^�k�(���x��ݺh�E�#��FK��g�ye�������&r\K7he0��wYuخ:��S��k˺&���-�N�un�b����ظ�ɂg[��/�F�O%k��d�͋]�:�[ٶg��\W/Q�:ݷ�9�V.6:�F��O�I�4E��$�t�x���}�0�%����z{&Eb\���=OQ��n-��Tb�\r��vmR�\vzx�r�G�k�.Š!�ܔ�//��9M������Ex��x�ny��2[	��@ۮb0)vŌ۷&4@uf�b�z�jᲕ	Cjٛ(a��**BŅ*e�kv��*��(��.����n鴮.����m�]�1t
bY�L3#f��8�tsֶ�.|�M�d7������L��x8ʄ��[�����hX�m���`�s��b���;]��_8
wEĜ��x��pP����cNX���*NN��g�e���kɩ�'����#p�a�:"�x��*kW����)v��!���0Zz��<�;�s�M��z]6��gOMn�m��뮍����Q=��W��m�]��sg���:���`������	�B��vgٶ�Ŋ�]�q��[����N���M�͋��Ѷ�z��E2u'k����vd�2Մ����l]u���t�K�،�7�9����#��l���M���P�h��.4��w����ٗYȃm�۝;���'cZ٬s������N��{�qpٴq��6�e����&n��,3l�&Y�&�,v�Nv�9�=�q֑ͬ�׽���`��׵��vZ�Ͷ���-��mX�H�ěSk��=�g M���=���b�
[6S2��Aّ ��m�s��t�[d2�Z����$�͝��[ge�e�m6Dٶ���øf�;A��z�����i��qC4�s�gemsl��F5��6���,Ynf���4v͛[��[�3zk͛9�ͭ��͹8�jb�tm�M�'/={!�o<��V���Z{y=���	m��,�AȊy�{W��OMe�)�gol�	��fֶҚ���`fVw���H�;���mg;k"�-���f�h۶�g G�y��kN���(�5�ݏk�ٻ��l�fݳ��;��mlkZ+:���'kk3�:����	/mѭ�l�e�e<4��p�����i��U�|�o�����*5%�0����"�T�&6��%�tL[xlt�R\��&��W\q����n;��h7i���\��-�5Ӻ8杸3]^�	8ݭm�r��TΞ^OZW4�H\SY���3M�������k��Mk����>۷ad������<]�1v$�H[�BP��K\2��1�Z�P�-��a��!�Ny�m���p!kf+�u�%&��6[,Y/h�M��a�GCJM�.���!�q�uq��X�gp��N{[[�%�n�x"ՅE�Bm��]0�V�1��͆����įY�nfP,p\�F�9��P&<�]��;j�>��<vA��Ѫ�e9��v�Yr�t1�81f*�z�}Qٮ%��K�3��-�1���s�hyg�rů�nQ��n�UӃ��s���rl��[u���������R  �L�	m�YC��Y�����mP�bR RYc5 ���ЗZF�:�x���z.�����]�h�u�wa�c)�׎�|���o]u:��dS�#Cf�ˋR�0s�b��\�u;�ہ�v��<չ"+spsA���xMu��� \W�y���pq�-.ظ���>;ZG�4vN�;S�լ
^�nPx�f���k�<��'Cj�cT�ˮe�q\94�9칗٫5��ΝΈε�\���);'Psk/V��A��GFw`����c�c�X<���[�뤭�my3q��6��]Uk�޺#Y��o-�ۅ6nC��Z��Km�X�<��`W{ ܇s��#8̜7�6sÞ�R������]�\�9I�PD�2׭[���2nM�=�:��S�lH�e���6 .�&�P�I,m�eإ#�ԉ{2Ԓu�8�XXܙ�A ��l�抵{���s�ʙ�������-���\9���P�9��:�t,1Cn�n���˸��<��n6P)��w1���2��͆K���������;��٢������]�a���/����IKz��*R�D,Q�����
�d��(J =��+�����Է2��8�y���v-G�^�! 2[z�Q���Ea�-(�Z�Q�6Q=%��3['���ow���Me[V,�i[W�J�KRV��`KF��%��k���J~��E҇$tO�;]:ȝ4������>y�}��X^BJD*T�?���0#\yxق��T)ɺ���K��7�K*�}�̖)�OB7�X�#��̏à��o���Ck��yx�G�sj���՛x�w�@��@Do/#�xS�^���A5��D��fB>>�A�DYS/�z:������=&\G��܂���әk�͟�K?zj�S��x0}<�����n�_I����Om1����c�S��"��{���{2+�� A�b�B�	9G;��@�yf.�Y���qP����쀁����}�����Nd���5"D�&I������i���B�hs�]K�{l��έ~ �p�>�A�������Zn�x��e�{75�xn��-��p"n8�f@Df$9��J.�b�.�J@��~��k�K���HZMܭ���wj����z�B�t���v�\��"J��A�۳�Oi��߻�j<���;��m��퍊��c�T A�/3 R��Ȋ��{u�@��9�n�N��-8o��e����ʺ:��.[��o/v@��21̄.o�h��ձ7���_B>#1gi�u֛��8l��q�A/  D�eB�q��9ȟ�@�̀�s  9���v��n���U��۾wMM���j�x��3 �3N��>~7�������e�s�ְJ{r&z���9.�	,�e���U��Ȯ�����I�#ّ��s #O/�ʺ:��-�B6}�����]
�@���W�̀���'2Wc��̋ܛ#k�dQj<�=;.���݄��ˈ�	g
 �/fD��n9�A�<����ߩ��Ki��<�����oRR�@�;�J�bΘ��F����`����ꈃ�M^Y�΢[�S�p�[ެ|t�>�ўj�4���yvƝf���,��5P����Ê<Fb�2��b[�iQQ�b�8��d�W׹f��VV�r�R#y=��W�sm�w>�X��Ybs���B��̇;�M����)ǻ��j rk-�_E�ON:L�� ��e}ܽ�A�Ä=����ub=��P�ųE����1��ɍ4�I�y��[r;Ȭx�F�&&N�y�	΀�A�d#�C1���,�u|8�37���zC�{�(���e���ʌ�,�yʸ���i[h�6�5>�y~�>�Æ�9���YGs�Z���F���dvD��H��v. Hqd w!3 "0���B��Aƭ(����q�U�e���dˈ� �e�^̀0��3����U*뽨�pϷ#՘��v#�۫�vh�{A�#�j�1���1{՚�Vv���oN���&���:�5�jSS���>�P�]C��W���yj����SR�Y�AF��j�B���(���G2�#1s#b�b5�(��,���77�e΍jDl� Cc��"��N-�����1#�!��Z�Nim�4n�h�J`�)����Q!��uǐ��0��f �L���w�6�t�q5�f�KQS18p߈#�}|_��(����.`�qg&7#����"3`,wv#p۫�vl�{A���@���aμ�����4T���E����Y�Yq�*�1�ǣ����o��f��,������9��و/���&a�\۟@̈́.�D3�G� #S8�����y��t��� A�&�����١�.3�-߷�Ӛ0}�ӛ�5���=��Ԑ�kA	̻�^UﯶLfל�@�U���1yx�1O:"�]8:GV�d��DAٺ8��Q���{
��]Y ���,c��vrgtk�F	��!U���Y���*mɾ�����H!+���2����q�.�=GS�8�7Zz��g�R�:���"�ל��e+ ���wM���:G����Yu���7s��ی���q67Ttt%���u"�UU3�z�`�lA��+��li��M��њ�x�Z��n]U�ܫѺ�lU�Wv��cR�� ��1�H.��A��k-(��m���.1W-"�Q��bMc�)i�`󋭻��1�J�SZ�ZKt������]���;��=��Ф�r�6锛���e�߱��ّD3!x��nY��K(��#y+�UOD��/c�1}���9��zHc�m' �0�l�v �L�v�͍����+"8-�w@G2 ���vcq�P�h K�x�s #�FbqL��9��օ����9�}����<��x���ļFb�D\q��ܾ�K䎘@��� Fd#W��f�FQ�=�$F���2��p�q0����Gو @9��1}���Fոڙ�㊼�53�����xڎ��#� �p�A�r�2�3")(����T'L���Z���Z��ڰ��Nz��m�3UA��3��/S�sUUQz�N�K���/��q�*�a�YyI0���~�~���3��[m���%��FZ�p��9���7a1p%�Af�쨜�����َ�T��W-u(�'U�qMT�H�{�� ��;;ݾ}� 3�Ϛ��/�.�(��\<��)up�������AF�_V固�+p�i����=�3�/�ܕSR �׽֤g�P@�-�@���#,�/*����Wf\-�<:����T:6�%dGYe{�G2p�^#1y��C�
&�@��3Y�v#p���_l�͡�x@>5P�EEghwxt.ɶ2�#�!܀�d#�8P#2=�*�ӽ�<�O=�]�n݅��"�	y�w  C<B�̄A�WM�ksٷQ�6�4(̉0����h���#�a֫�'�튩i�=i�:ˍ��z������<�mÇ�1*%���9��<Q�VD{6#)�:�{FO.� {#��#1 Nd�4B��^ta՘D���A{:��n9}���0��T A�j��8��L��s6&�g�e� A�ӥx���2>Ä]������ܜ	''�yWMebu&p$ј���ݝ�ڴ����x�"sL�%Ėwwb� 7Q}��y3�Ā}�sD��Y{�qybp;ȷ�B��8�-;��n挢��2K�O�c��1��O��A
��T�K�عL,��"��c���Zk�k���eX���Z�7 ��m4}i,J�};��r��o�؍�ӗ���1�C�ƪ�����[�`�z˺�~�Љ;���j������s+ZU]��\��j1�Z�:�Z��[*��~ �:W�쀇�d A8p��=wq{bsM��B�B��no٣�/�H��C�: � �Ê2<d>=-������D�Q�x�:�ٴ��gb�0�#���(���"u�"�`��:|�8�/@���Ȣ�B`��JS�s�X��~�Z1m+�U���#!#1s!x��ɡJD�ږQe��x�r ��
7}]�Q{bpm�[�!oy�D�����'�j�L������'[�h˞&���{u��H+f���8���Z�^,�Lj�$7��EeͱX&5^�S�v���@�d"�A���ӴغBg�`h5!��N��_.���&�>�^̏P9�'og��8��Wn[��T��0PA��g.���0;�,d�B�]���n9N�rQ�Lj8N��x�my����\�����[CyDFq]�.�Gle� A�^������ӛ�ӿNa��]R��4/�� }���˨��9Gp��!o |w ���s LH[nV�!N�3c��{����qG��B��O��݌���YF�/�D�Ȏ �,�w �d A8p�2�Qճd^^�dح�� ��>�A1�W`�5��]�5P� j�����2�6�wH@�-���Dp���/�^,���d��`�^:��.�;�v|$-�;����/�@�컀�7Gr�x�ㅆG�.qa[��U�^��MRWuz�M�Vn�Ҏ�ڥp�5��Z�Fmh�$�a���ӕ��^arvy�G�p�n�Oov��M��n.M�6Ǯ��]�uU�`�\!�u�<b9-�Ի��:M�6�5�X��ܐ�R.sh��������"���3j�=6�������v��S&���:W����Y�j�C���J��.,&y�^�^�\J��U����N�)f���Z:]u��L��R�c<k��wo��|�E�����}+ji��ZkM��!����%�/5��Z1�a[F1k��hOw�������{��{2�Kq�JX���t�Y���G�����䦦sft� �M��w��8}�As /�̇Q�0�2�E��W`�5��]�uP�q���j�$u*�b��}:����8Qو#�|0ޙOS���1�����;�[~�E�lG9E�=g9[y�-8�)��}�4��]̣��>�sCY���왗�2�ȏp6Y�Q�pv��[2+Ǻ��z؜�Nr��NWǜ��>���qx����vk7ֻsaP� w���a�#�1x�Ҥ9u���R��a�����T�ƺu�b�1���'m�HT�D6�8�p��t
2 �8P���ʫ[bU`�o��ܾ���ᚁ�~K9V"s�Zq�[�P:�5}Ȓ���웿$a��Y���T��k���{sY��CBA��{�op� b�;b�'`gsݳ�ū��T2"Z�N�w�-�qYȪ��I�9�/�4;R��fV�L%�A����̊y�*��\X�,��x N8{#^9��#2I��DJs0pZ����?R�ͅCt�~��D�YiǖTNr�r�'y���;�GI�����ǑÅ�u�UklJ�-𠷂������l�v��8�� �qz�m�7�+�9ҝ�G$(��B�.�[�0�Dw�&�(FoO��,����cGt��K�{l�]��m]�9	a(�1�vT����R�
T�lߤ]�@���"�RA��U�,c���.��T0�z�n�HLEuZ�sAǐ�ۑ%�@Ae�GRa �f�(�y�mǑg����vUE퉚���
ozA;��;B����\���@�A8��r�����!�>��]4�!31rH}G$<������H�g3�a��OjP���n�|����q��D���m��+�\�<��oU���sZ�±�S�ǯ���>�sg��A����X�KG#��{׾�l9{����m�D���w��N~�ԮI�ž��۝<�x��m�1�0���C�Vt���m��!=�Q���0}�,��8=�&j_3��,C�(~�8>�S�o6x�DN���_x\~>���^�_LŮ���vug`�["ۄ��ԥV�p�ѧF^� ��\&,��w|/]�e��ӛ��	ԨsnM��yc�z��6;��C�}�'���=}�h�/g/ga݆4����zV���uƃO9Y̅��<�XN��+~�0��q��4i��KR�q1���⚛^��w;�����(�{|w��t���',�Զ׆5�1;nwt�V�{�9X������-�͡�2h�؞�ɻ[�!��a���>��7޽����	s�{ڦ1��S�e�n8:<��计X;V���o���S��6�of�V�7U�8��oR��3���H�ea�#4L�b�8�a�]}�������{91���^4-ڡ1��2�w�����y^d��t{Ã��p�b^��j��ď/!�J��[��=��q����=�����|ߏH��o5��}6v�:#z�C5�f%58�ѕb��Owz��%m�qE�NMU��Ui�F'gUd�X-E�mInR���ׂU/D�Í���+�r�a��ӕ����| [��ESB%	H�A�q�l�G,���;9,̳Zܝ�������Z5�k:��Fvqm���8+-^g��m�m�M�3�7 Am���Z֎1�$rM��Mme�]��X����8���6�vݠ)����;6Kls��U�&݅ΖSk7i�(���Npv͉���(��`gA��7(�,ݶY��&k9�q�v���@�{l��[6cb'f��6���f��������nm���m�Y��l���YdDIu��2;�����$ (�;m�&m�[kX$36��kf�q-4)�Vt�G/4�	�[f���m4�%�3,;�"�&ݹ9��m�S����M����t�9��;l�M�ֳf��P�/=�ǽ��j��^�C���m��Ne�J͵�9vn�V�#5ٷ9dV���-l)��lvd�R[Zq��3m�����l����NI��-l��dskj�S(��z����{��3�ޫ_��?]���YL���RRAa_��Ci��
@̢�hB�
Ar��R��̰�� �>��c��9�39o��G��G�5��RAM S~��L�d���!�F����������ٍ�$�]��ZAI@�0���2le$��~���Wջ]��m �5H/�ˁ�tAH4T?w��c�3(��@���)�ˁHj$��³3P�Aa�� fQi>�=�9G�V������Ad�2�W� gכ�m�6k\����:|�XV�a��AHQTQiE���oځI4�3.f�) �Q�4�XsW_g/���z�Úĕa8�(�FP�>�D�B�"��\ݷV��j�Ɩ�6D��Vgo�jx��ai ���i�c) �T��4�X�$+.��
A����
#������T�fg_�1?x	 �"> � �|�Y���Y�rw�gb����) �߿\4�R
��q
H)�ˁHJH,32�c�����3(���!I�{��{,5��������
Aa���3�2RAB��F�g~�٭��w�~½�����H))
a�߮d��H(�- �5H.V\k�w�|�^���� �P�~�m ��
@��-4 RAe����R�) ����6�XlaH�ZMRAH.V_�� �f��ٻ{�:6�L�-�>G�µ��
B����- �RAh��P) ��)�f\4ͲRAB��i ��aI��0���������ۺZ�~aWۆ�:2�
yE��H.V\]RT32�(�j3�s�Rљ�T���$����
H,��O+.$���9��LT���̚�1����Y ��Ʊ������N�Rw���T�u���S�Z�ͲcsM6��N�ىJg6B��;��s0޿n�<���a����
@稴��RAd�����4%$�a�i!U@fQiE���TH)�f\4��x��0���]~�r�����u����7� ��'Fy�	����X!?~�!��m� �6��b��XZ�3�d)2����v6��,���s�^q]��t�snKmvR����3�-;) ����ʁhhRAaY��6�Xn0��-$� �G�;�� Nd�|��X��e���Aa[퇣�����u~��7�w�_��������H)��w=p�AH(m�4�Xj0���Pi��
J�S̸i�c) �{w���~��}]�i��i ��@�j�<	����H�&��B�rR�fg_�1?x4����$S%<ʁi �����6�R
e���Nf|H,��{��hJH,7��l��Uܢ�
AH.�e��AH,32�pd����E�m������L�m�B+X?���Uen�����K�0�AH,=�p�&��H(3�i �4�As*�D��3.H.���E��Ͽ}��G�Y�$����
Aa��p�Aa����
Ad�)̨���5�{����ֹÿ?�x� ���ᤂ��P�E�B���s�����_�w��S���z�n��P�v�$�) ���4�RP�0�ˆ�62�
e�H,4�\ʁ}�~������� �y�����6|s�z��s����k�4����$P�O2�ZII�O������P3(��B�%2�ʁh�ߞ�~��+ޭ��w�������N)�2��Ƕ�O�Yy��R�Eȍ�geۣUo	p	�a��i^��ʤs<���_�g��ߤ$<���?}�{��nv�Em�
2���b��q��!g%�h6,�3Z���9N=��s�:3��}�&R�ܽ�8/R�l�f��l�
;��m�-�'��������ô�ySAvj��^Y�]nYrXQ�<�uu�:�N%�����<j�e�I�q���4V���P\T���Վ5�s|��ζx�=Ӻ�B�ٜ�:k,צ��!h�!�$����r���6�2[;�wZ�����1lӷ:�Z�A�k3Y�DΦ���,�oO޾��Gi!U@g����R�����SH�3.f�) �Q�4�Xjg~�ٯ}����)�>H/�Շ�ZAI�v�g�߬���k�\4��I��f�Q����p5tAH4T32ᴂ�P3(��$P�NV\
CQ%$־�w���,��]W����Ã
@�(���RAd���e��O���߾~�ƹ���>8�XV�a�i!U@w��uD) ��\
H)�
a��1�_��(�����AC�}F�F�^W.$�B�{޸i�c) �Ve�H) �Yp>.�)�f\4�&��%�ھ����:fm�LO�H�E��
H,��O+.!�II�O������q� fQi4�$��e��	I�fXm�AHUis��U�_.���xQ
H-O_��
i�sݸi����P�3(�Aa�����^�����)�>H/�Շ�ZAIQ
a��p�&�RA@��6�o뾘�G�>L�M��D�EC�ˆ�����- �hd�+.!�%$��6�Xn0��-&���{ݧ���)�ˁH/5���n��\�:�^��
�l=��U��ZA�������RAM�3.f�%$*!�F��}�������}?`~lSd�[�h��(K�M�oe������c)�4��Z�Gai�z����
J��\4�R
��4�Xi �Yp5.�)�����u��>9]�gs����k�4�ˢ��$]u�^����_$���Hu%$�{P�AH(���B�%)�ˁH�I�fXm�AHUP�ZAH<	�}���B[v�}���4��\=l��h�N�}���.��'W�q�x�wI��[%���y�׺C��:��[nI��-tՒ(�_x#��� )�}놙���
��H,3��Üs^��s�}��$�j��H)��e�L�RA@�=f�Q���e��9���e���XAH,+�p�AH(~�Ө�Y@�Ok��В�
���m ��aH�ZMRAd��r��R��|淭ֹ����k8k�矫���Aa[퇝�����ZA����oځI4 S̸i�) �fQi��RAr��L- �o��o��.�������I �g�ZA`q����p5tAH4T32ᴂ���>�]�gs���iנi�E��) ��%<������X~����7��]��R9E�Ѕ$JO�. i) ���a�i!R��- ��Z�y��SH�3.g4��}���j�o��x ��O��]��bv�Y���É�Z����
Aa�ˆ�62�
Ov�$����E� ��ˆ������z�m���W�3B�ik(h �iS��8v@pa�m@�b60�v��Z+F���`|���i��YL������JH,*w��6�R
e�R'��e��
�����]�o������Aa]��ô������w��ƌ�U�����Q
H-�ځI4 Sf\4ͲRAB�̣I���\���ai%!L32�M�����}��w���g�ϼZA`q���_�$����2ᴂ�����ek8��o�{m��+�Zx@���d�����RAaG�{P�Aa�aH�ZOM?t_��]���Ad��~��
@�RAa�~�i �6U�QiTB�A���I4 S̸i�d����E�����:���O)>��S�.�L��a��L;��.Pn��v=����_�ƃBԣ=�ﶥ��ª�d�ZЕ�G��������gnD~��<	q(?���
J�̸i�l���G�f�
AH.V\�肐j����l
@̢�Q�7z;��
{n��O_0���p) �?~�Ci��
@�Qi4�$Je9Yp@�R��X��9\���~G�>؀��AHUP��tQ
H/�ڮ?s��}|�f�����Sb0�߮f�) �Hw(�Aa�aI�ˁI ��ˆ�8�H(�ZAH)�ˁ���_�����AH<�s~�m �Y���k�:�7ｦ�H�- �xd����
Aa�������l)2�I�
H,��+. g����t���|ŕcI�$)2��fQ��9�A��m<�1���yq��c�[vF������pB�ˆ�
C�Tݢ���$�_��
h@��p�6�I
Cv��O��.��r�����Q�G�.5a��Rw��u��k��
�nd��H(�I���A{Yp4]R̸m �`Re�@��ʌ��e��5RAaF�w�;{����v)���x����?"+��`]�u۳?i�v�H �@D��͵��C*�[�"4��j}��A�B<Cn}�n��|�ŧ79efW_IJ�=��e��[�A,��m�����%�d2;��Am���m��qY�2,a�;�u��Q����C�+2���ݵ%#�Ⱓ�==���L�~?zPyp��z��Ƕd<��� 8�7J�L��%�A~��\>#��.}>n,��Q�'Ÿx��CD8P ����ߖ�O;vg��;}���>���mO�n��#)p̭�#eA���q�]bā.6#�i�9춠ʭnw(7g��.�3b
#@;�H �Ax�Y��rh�%˲�*���7��'�͸�W{�~ �� ��A�P!�"A���e���	�"A��$��p��W<���v͌3�;�I�C.�uXǑu�N;�[r$�G̲�!�"@-�,�>�Lj���v	�n��m7�x����A�P!:X9V]���ֽN!�^�܉�� ��m���D9�Q�ᓏ�s($ױ����D<P6�A-�D2�mh��.u�HkR���\�e�gl��< ����;P^!������
K��b�kڕ[�޵��`�&�+�7G{���e�:�5�z)�7=8A�൜�����g�j��l�|V��,Q[s�*�A��Wz������aAZ�v����t����60��[��h��4�ݬ�Ŧ�k��4�%�B�uN��C�A���LM�c����Č	۬:m�;OGGl��ҤP8�v�mx��x�L�Ҳ�[(9h�n:�ݣ��-u������Eݺbmpg��`���6�L�7�q-�6��WX��jP��di E�%2G������I�v��;76�����N.g'P��4����;���-�x��a9��8��Z�RT(3)L�|'� <�q�,���`[�w-ٞ�`���aRxw��������.4��7�k��mI���`q�#�_l�;�b�.^�U��q��l���$���h�a���8Q�"}�\2m�Hm{k�f,5�u��,�v�#��40��u� �ڀeЏr$�GV�0pv�D�p��e�O����n���o�{x�qQS�g�Hû�H>�/�>m��6�2�I"[��b=<;�� o.ł\�+2�;�F�A6Y@���$�K,䞳X�W]�Wt�;EBB�!L�0�i7>�nZ7Y�6n����*�W�LVl�k�}���_�I��-� ��=��[O���d��\ v����Wת�#��DahG�n|�YŖP#�j"�. �	 ���.�G8�'!����vh�S/,����ה���U�*pU�/ MKR�ܞt����\j��J�{8����1B9>�Yw��ت�e��x{�Z���� ~<Tr��`W�w-ٞ�`��7�#O6Խ��ڌ�`�Ax�-�Ch"�|�C����dۙ<;�VaY�i�0n8[��#7�O�p� �� �C)��7Օf2 X �//�^��|�	mgK��<�C*8��RA�ЙxH�XX�n�{�'Ÿ^ ��/�^n/�s�9�10j���s�;YLOi�v�A� [��Ŷ�[@������[��_^�A��c
3$)F+Xn�]-��]��2��l�D`P�O�̘��0*�A�k�`X!�@������/ūaf
��`�z����Qq�.f ��B@=ЁŸ���>-�@�����71�w~@�R<A���a-���g�Pʎ>�j|A�A��Vt���)ǞX��{�A{CnD�����߽������\��ݜ�(���B��K[{k�x޸���pF닻��H�����|�^ы6r�}����y�ɽ}LޤG�"P���S�!��>�{�Dn;��-N�SV�Z��� Cyyڐn7��s1�u�������G86�I���հ�Wq0n;��� E��*3��%���D�x�܁ ��A�kȶ�Iw���=�j����]���֊Q��w5H ���� |[r��u�;2v�dF�̂"�طd�z�tæzմRpc�1(;��-���D�J��h ���5��n� � �^u�ڕ;�o�j�kzD�
ܝ�^ ����������Am�M�bF྽�8�q�6D�VU��h�
��c"8S��Fw!%�;�i��r{����������<���%Qv�3��kͨ�u�N�m����֊��� �Ax�� |CnD���ͮ�y��E�H�мA��g]�ҙ�V������ IP�`�������z�^>bK�0<�aJY,��WɅ��p�=���/��YH�X�D��H�����)�47~�����L�_ A�@7�	m�7 7�K�p2��4�c��UՒ*�sV�1� N@�A�>n/��=�7?��;�������h��=��lu�."6������^6�з�qZ�&,��~޻K~z#��yڐCp����������s��e?5ݱ���#\/r$��� �ѕ]��nԌ���B6�;.������ސ|v�/w��-�*0��`E �܄ ��|���<h'q59�R��,�$R��]Ĭ��N �ޟ7A��~��c�ʻ�0A�5�s9H ��^{U���+�<!��;���|p/c��;��!� |�BKpp([k��Z�|64'On��g+���5����-P.�H'n Cy �VAm��j9�]�|�Y�?^��ޚ�ГΓ&���K+&im�+59��X���N��Ӄ���R��S�{:�ŕ5N���wox��|�-�ݕ���������f$�@��O���ozώ�PkG���3b\+x.w���v����d��{˾��o�5n�{0�v5K�sfLW����s��$��SaU�y!���G/�AB��n�y�F�=yF>��T���<��
��=��?Չޡ.�I�PXbQq8E��i���8����	g��n���!h�ώ�/"G`O��׿{��yxk�p�+}�![^�h����{��^ES��oi�'Z��&��F��5���������Eɝ��:��z�_aݍ���~���-µ��f�3s����Q6�6Ӿ4��v�7�/�b���]*�s7X�;�J�>���I��{�t^÷��v��~24/&�G�������`��g{�������f�}	�̳$6��3�,M�Xk&���j��!顯��b� j��MX5�|�X��oq���*	�t���4h��"�6����/x�0߆Os���1xk����j {0�oR��|�Ѫ��\5���)��l��]���V��]�����������K�lK�D�o��3t��}_�������Ƿ̬�u�.�����܍̓���裮72nj���U)��3�����}}��Ps���T���N(r�v؆�4J��i�7��T����:���pp; ��r��y�/N����ڽ���5y3\s�9���e���kbsm�F�@ DB	iFf��YB&lJѵ�kl�Kf:��lP����LG)Nm��;��yf&ՠ��i��׼܉ܢm���� ����N ����Ȼ9kq�Km3��ݚå$��(���hŝl�vn[h�:yأ;��[gc[lvdRt%�&q{z�{e�洖�#l�4�J:��f����v�l�1���,��(㼴�*8���=��t�L���<ּׅ��/4�j���$�t�/i����F͓7���`e�����e����ޭ�"T��<�ͽ�=�Yb^W�ۣ32��{yMh��ް�Q^dD$q�6��G��{w��Zv׽�nά�#�㓌��:mfegF'\Xe�dg�݋l��'+o<�;K��(�-�c[��0�I�{����v�玷mp/'�9<z�4�^�؄�����[u �"I�u<= �6�C��m�r[��M�)�SW%��Cl���a�Q��v�fpmh.���0��om��Q56�7M1������h��.[b�Qi!��A�a5
�6ô6��%,Z&�*�L;(kE3�����d[�bs��J��R5̮�^	����<%�,[��1u�N���i��jDne��c�y*�c��T"��d�Y���8�ݶ�iu	���P�X^��È�0��v���T�0��l�j!�^ƅ�ʮ�̡���$�[f��8x�ܢ��i{Y2��lΌ���]HדON5�5���͊+�z�ū�C�9��[i�%/E��l��'�u�٫42Aap��Pc��읤��!��<y���G]�7��
�[��z ]�[����K.�XYlp�V`���{(t��ė�;6ë*n��rC';ɺ8ٔ
y����sl�G<��.y7^�@�k.�!�&�>,��z���AXݠ�7cu�ك�8����9Ǟ��7 ���=��V��15T,�hen���(��Y��e�̜�#���646�l=c'!8v�n�N��m�\���T��QI�m�m�:��.�y����qj]q&W���wV����u���N6����f��$����sf���Ɏ����e�S�D=ܝ+�ā�{]s���T|�ۙ�
e��D6��lI@�3!e0�ʑx�˛�۬�S��4�\�U��&3��N�{�/8����h��\�G�kt!`�م��� nmfr���%��«�����³V���bI3�m��㱭��4ܫ@��!��^�N���㫄�̑,���L� u]����iVȉ���vٺ-������U�L��#��4�Zxa�X��.�Žmv��a&���Y]7Yt�ݗ��B<��-�[t�]�������F�\��X�n��&W���ۮ�\,�0�y��ѝ,�Ej��ww{���㱔7�t�[r����k{hb#J�]�>_ �g�Sd��x�E��p�m�ft�v�l��u<3�����g���NN��W;e�M�Hp��e%�ukz�L��v�\u�x�s;M�.�_"kIt\Ѻ�����ڭ�>��gm�&M��u3�j{u������\���Z���iX2���z�@t�cX��b�渵��/�~����ؼ��<�e0��"�3�s�\��*Ӳl6�S"$��
? A��Ԃj� |�C�'*:���&��Y�f��Z���@���$�"�m̂n>u<N,9!W�q���	��n:W8x5�è���j@ ���qڴ�N���5>̋p�m�%�^>nq�W�Nne
�{ٗqs=o�-P.��x�7��`Ch n�ܚ�{&��@����m	�� �˃x&��Y�N�V8Έt�{0h-���܉�"�@6�zdJ�<ͩ�[�sZ!�z�+��GE���p �A� �r ���y�k�[+�X]2m4n�YN}c�,��9�Ѥ,��e�fs�vuT0e��>K,�~�/6D��ȷۗ�6�-N�[�T�*���&]F(u|��Y	��w5H ��@��ȶԑ��q��[����Ɗq8�#�1w1:��3�6�UeU`ܯ�/�����K��m2Ѝ�r�sn���1yj�~},k�=�L`"�>>�}�'�ʲ��,E����W���p7�In:r���q�$���C�29��mY�7�땵�;c"k�OG7���\p�a��A �>!�n>!�"@-��a�f�vD��D���l�\Z�����|�v�3;�,e�~�u�Aւ�� ��^��^!���Y#2o�ِ�'hA����ox�q��@��ޑ ���̊�zz��<�2�Q
!H�g���jqe�!�C�5b3ƕ�5�J)c�!4u��k�I��^�Dfǐ-� ��F�d��RW�q�E������k����NT�[A F8^>-�[� [�����Z2$tn��h=��>/`!r�f�ũث��j�w�n �yyڸ�7��Q���x�p��I͠�>>m�~#V�E��ɵe�G�ٵ��aS�d-������ѳzf�F��x��Dc��^���d�4{ӖFb~�����ó}7���<V��G���z�}�z ��M��#�A�szD�� >-�D6��}�:�=ٰ��p���^���\>ۨV�G�>�� �'�iM�1D��.�D�0 �@D̑'5�*-�x��G\�t۸�=}�p�}��o j� ��po&;���Y�;* 
QD��s���lt���;�@:CZc \�1�%,.�fn����?Ng��l7  ۑ"uV_�
���o�%\G��Ǟ܍,�dWb�tYŖP!�"A���9<nuS�(�RAƂ�rK��t��3�E�W���˰��Ŵ��u��ȟ������-�[�|�5�M�y�N��oo�w,ڗ{�p�hw��AB-�> ��@�Ph�w֢+v�U�A�FQ�ۑ3���Vm�	��VDq8QxQ�]�N������7����j�G(9��F��È�~�\�M3��?4�O'���MA��>�'s|�[}فfJ��e����9��� ��t|%�>m܂p�>m�f�|ui!�J�Qq�m�O�]���R;�]z<�Bc6��]���������4�F�f�J���Q��/-mktDn�c�hAq�a�,�og�-�}׬��ﻛ�Ye�#�_l��jv/�v�d|$(��-����Yx�s5H ��!��û������vH�"��!���d�*��F�ó�o��� �¼A�"An��9�-N��>o,H'\AŶ�-�d����%yQ9'b���<*�h�����7�"k��ۑ>-��%�);q�Y����|�+ѷ/����[k�v�dΐ@;�nt[)�5zD#��AZ�2�@������W��Dv�
�`�r��"#bip�7�L�G�����B�q�,��t�N�eV\[�dF�eΊ�t�l��"��b��b)nWf��l����*��d��L��`�U���O;�u��i��u8�K���Y���� �qq�DE
Q�n���֐5(,Ř�읲-���7f���p�Md0�Y\��"�<�&��BX�aF,�(m�U�����ts�5���c%k!�蔎f��Mz�����K˝6lƆ�n�֡��Qۺ7[cZSmD6)Krr<�\�9٦ �E�V�d���L3!�Y��n�ؘ��b6�J����v��܅�9')���jA�;���v��R9a����%Ƥr`�C(XFmJ��sKi5�$̃&T�&��r�Ѥ/ڟ[@�n	e�I�W�E�W�r�󊉩5Ҭ��h"4�#�͹[�f�P5v�*� ٹ��0}Ǌ�V�5�\*�]{[ �p�k���|�@�ua��F'��Q��jA�!��ŷ#�b���V�K�I����{�+�f���"�,��A��Y��i1|Aq�ל�`6�G^���t���E�W ��R}Q�.�_F	ihG��$�K,�-�pb��*�\vwY����kʸU��r�L���A 뀈>��-���Z�G(�֧E���@�k.7������]v#���C[Dc���L�a)����\k^�f��e������T��7�L�G������3���q�,�s�Ÿ���0�{"yV��اa)�����<��n�y��[��yYkZr ������"M�#��|�y�{Bfî��ET�)C0K]�|  ��� w �_^���m�b2�h���s�A�Ah���;�$����"|� A<Y@��[�A�z0rWֽQ�#1)쨽ʸU�}�Z�A��$u�^#O�mI͠�e�;j���С_]��^S����y��!S�"6*��7�h�G�e���$d,Sa�s��"r$�A�n-�sn���n\��5b$�JӼ�S�|4_�w��1H � �|�^>mϋ�!�������z�t�N2��Iug�Ƭ\�0E۞7(��i���2������l��l��n�(�o�^U­�幱(���٪���YR��@�/ /�Iǃtڒ!HO�\�j(I����ș��ȃ��1������VG�oH���M���# �#:�d�7���|b�_^��0�
�g�Tu��U��()�x�G"�4ᚮ)^
K�2eV@4��_W��R.�V+M�bo�y������US)�5S̘����ཹ�Ӽ�>m/�����S���V��P ��t"	V�5�Y[q�7�i��:� }����
c�v�#\x7^@�ڒmx7s�=%ktޭ�7~�~mb��$���=�q�Ed/��n��Yu7���KzʈQ	�"PI		J�1	S�v�{{QB����Ǝ���If�ږ�tu�?{��K���s`/����KoJ}�dޢ�8h�b��GcwPY�s4�P ����^-�q�Cq�-ދA���n"�Ās!x�ޅ��k����ot�o�p��y��u����F8;A���R-���K�܍�S�=Ir�wc�/t�Ȏ VBf�q�Cp�mϽ#�Q[�T�@vӗ���xz����^[7�jɛ�+���\'s��ogde5b��J���	!IF�D����ѧ$v���az��_{˕���"���+�s���c��]��fj���x{�,|}�KŽ�%�@�n<�B�n��V9�*�I�Y�|�69�Y[q�7�i��\Az��h,W��ٍ��z�O]���tn�0��������ɔ���1���Yw�n4��i5n�SS��#�e��e��ǐm�GT�A�T"��tȎ>ѐE
2r���5}>�A7�܉�x�G�B�:�Ff(>��RA�r	m��}{35�����]�	��> ���|�^r�y~�ʑ%�/|Ft"�r'Ÿ^ ��a��⩬yi�/.7'1F�嗺i�ސ|u�D��Ԃ�^����W���&�����Ax�܉5��E<'�Ä�A"���!I8i͞��l"	��mȟ7-�^-���h��feb"��N��:z�Vڎe�d�ݘ�;� |�x��#KO3�lD�A6�R���̈�vX�v�Z�4\з�qB4s�^����n�̙�v۪d�k�y���6ЊQb��55W�ܣZ�����{�������"A�����q��9�\�҂.���X���b�q�Lv}Zw��)v�{{�'|/��gqtF���p<5����d��mwfj��s0=����;��i�β䩎(�k��f��Z��f6�c�Ҏ��ԊB��
V�9&��ZݻZ.��nBƞz&��m���f,�#0�#���^w'	��Y^�y��j������ �=C�^�m�܀�؄IGv��`�&)��$��'Jp���S�%��o�qǎ��� ���q�!�B#��k��ʳtԃ��G̺�BN#u�� ��^:�I�@���-���/�=>=3ՕT$��y�B:� �lP�xO>���"� �ޑ>-żyz��)���t`!(Dn��À�%�ڒ��Wdcr�NM���*�Q�sD�'��يA���z�s��Ȍ��9yP:�|A��^��"6��s��Ft�n��v��#����|��G������^@��^��G��Z�5qWֽ�p�ɭ��B+��}2#�>"�=��_�p��ࡑw�ኔ��ߟ���չ��G9���ۡ�u�T��B�.8z�����ݫ7���p}�7<{v<�VAm]�]*�Q�sD�'�"{lb477��2�a���ŷ"Kp�A!�@��+�.�k���aA�qt��`�p��!XI���
R�yEj��h�t�Iwa�:���#�,j����l��]�V)۴����ǲ�!�����Z�:�7MP;Kِ;�����jD'R��B56,f ����7�H7cK�6�3����*2�s`�\P�xO=���˄A��[�/�"r$v�y;ي|{ "����[t\K㲪�4O�8 @=����4��3���S��}�$�	� ����s����Bl�*a(�n5�b⯪��U��-�^ �w�"�RA��Yk�r������ _8l��v9��<En[ t�m]u�s��Fs�s �u_^_�>�jH#5��q�ې�)�1"�Ϡ�Dp"���×b.0��;���7ۙ� n^.�QS-����ڒ�PK��ľ;*kQ��D��'�����]�$��uL�����"Kp� �g�a�Kh^扶Y]:{g���{qn���s|w+/u����=��=9�_wU�|�����dǾ�3^B������,K���XϷ����C����9(���o��3�t ����5]�n#�j#6���2����v�Q'aÓ u��u�2%��]�^�<�L=[�2���^�����(�z��w�M��?��Ѭ�Ll'�^�鷭JE�<�Ve�����{wn�˥kic���n<�塨�ζ�nC�iਕ������+׷8~���7�$���a�t+�zm��W6���ˏ�j���/j��{y�ÊQ���X8b>9(7����i���xw��->�%�三Ѻ��+�yV�g$�ٝ�w��+T��zU�kZ�\�ɗ�ּ��%)�f�����m8�ï|�':����r<��kO]1�a��*�+[�◠;hu��x!��r�I]��xv缤��S��� `�����q�P��eY}��Z�����|_N��pN�+׎uƆ32�]+ډ�4S+N퉂��*ѹ�Bj��1v�r�շ��"���Z/b8��U�4�tdu\��v.��fwFjf�y�{�]���~p��zᶜ�z^}�T�C�{�Ӕ�u}toN��]NCtS�u��0�����F�h����K�}38A�z�S��l��O9�*޾���eU�J^;�?5V��oR2I�l�{�P��B��z(�i�������������e�[6��e��g�����fz��#4��F/l�6�ǅ�0�|�>z9�W��K;$��7�v���f�k�{;���ޑ�gL�A��Im�)�䓢�C��y�l֍���kQ��7cf�e�������IÀ�$	s� �q�I��l疀w��m�%6�mj.S�$N�$�&���G^݋���:ɰ��vn��88(!ж�Nr� q�6�-�Lљ&�[�99��%��#�É�gGZ͔s���(���;;3�[�mp��{ޗ�BI��9)ѣ��e�!Dgfݭ�$&�sLe^֜t��	��c�p�:rpm��9t�k!�	tS�R�Ą��߷����r񿻽�تk�H �#���mY͠��k��z.w3�q�����4>漼[r�� ����~"�,?z]�;�O!����7�ۙ�"-�@��^7y�X�
����h�Q5ļ�>���=���7��t�m�Y���g��}�HD�(O\��v��{\ޛc��u�ËP�<�r�]��a��~��g�,�=��J�"	�o�\�-*�^��;]������U0 ��9��Ch/6�ڐG]��)���tg����ȑ1�XLF�w�y�Ȏ �+!x��B|[�R�cdT��(�9� ���!�RAmA�q�BpE���G�*2���To�Bk��vb�� �e�!�"|[�}'t�BP��wa A,�O[�ܜ�5\��ؚk�����_t������5��J&�ؿt��,���}�*��۾N"1������m����
�N�}�n��&�9��9� BH姟w��O�e����@%��[@2�ˋ�1�/⩌s;���ň��x�=)��ZO�1G�}�'ŸD�*���8�V��
!)R�]3�d��f�]��/=4��<]��s�Ӹ�n�#%�y�	}�HE��[B6��=�P�����*M�!H�(�Ⱦ���P^>mȐp���5L�l��wr"�H;���o�Ś��^��;] �� ��mD�ݘ����}؂��[^�^-�u4l7e�P{Tn�1(GY���̈�@��9�"Kq�n!�"|vx��7sJ�W(�]��m���=�Q�k1��R���\�E�mG��ȟ�A� �۟7�]�JaG!�#��#�28���͉�v�H>-�@����RA�hfK��f����<�d�k��c��B���L��T�͢��+0�Z�*^��-by"�N8��U��R�L2�0�Uc�x{��뾻���0x�ָ�_Xh�+ݷ�p�^͔�.2�C��wc����Dc�Ⱁ�P�K�y}#��m���ku�	!����nܶ���u�1���].7!��k����"��#3�upَ�+d��uH�e���xK�'n��zN仛X�����ư�D�+�GNI۷���yMA��)��lq��㬝��%�1��ߟ׿�DX鱮���^yS� ��5�0�0nՎ�;�n����1&n��~��F[���Yg��7�ǓnD�F�aԔP�/Ϡ�Dp!���Br/�ޟc� 7ۑ �[�3Y�d71�L��e��bj7��f=���ؽ>�A���*b�U2i5������H�[r$�A�^��� �5���ȇ�����ؚ�x�{�"�RA���HC�Jd�]ɐ{�@=Ax�܉Q�XuB�����9�$S�l�z�M
;p���DF�/ۑ ��#�� [jc�3�'z��|�'tTv��+x8�c�]���) ��>m��܊W�V^Tl����ݵ�f��T�f!Y�M�sk�-v̞�y��]Ki��bm[����e�߱�,���[�@n��ވ��ͅs�y�hlWH,d1��jw >ˏfj�����p-�$O��ͭU6,(�n]T����/$,a�������	;�7�j_�[�Ӄ�?�����i�F�C��Qbnr̓�O���mե1��=��3c����>��~�;0U	b�}}2#��u�����X�X0���� �� �� my�L�CC����j+O9�+�8�c�\&��� |�x�ۑ �~��31��DP!�q� ����ä��}/$�/n��7>�!Z�dvW`$��M�) ����H[jA͠���]i�V[W�l�D����(��0��ȎwF�� ��CpLlGFZ2k����BT�}75�r��qn�'gq�.�)�{/^��M�f�i�+�� A�ݏ6Ղ�Ayt�g�J�K�W�w�-�>�%.^���٩y�����Cp�UL�W�4��A ��Q{���¹}y�46+��p�@@���q�0� �6�xgR��T�Cp�h�ۑm���ԍ���r��Z��?~W��T�9R&2��Uep�H܈ٽ��#��0�4w�S������]�t�vf���*���4��v\���� {���3�%C������ ��p��H�[�A��!�2%r8�'���M\���6�
��Fi��B��{�y� |o�O���=���5�����|�yx��[��-�q�%�h`#�FU�F��Ҵ����ؔ8�#���Ԑ[Cqݯ����Kz��5�!��!������<uO-ۃ��3c��CqԪnh������<_�lq�_�#������3d%A��=}2#�����ӣ�\G���D��Hn<۹��6�Ve֊qw��y�A�j	_RQ�Ol���^�^u�}�H/��f�YYs7���C|r�3a A�nD��A�Ӿ�7,`�X�/�6����f����[��'�<�W��A����;�V7�j|A�4��ǓnD����!*f�0��Ȏ ��p�f`�=K������S�ǒ�6�쭆)i�6;]�#}�x���M�(5�񯞖�5�ˣ�5r��Iy/$���9�������x>6�x�C�^!�2	n �� [h��}a65R�V�(�N����^�^u��/O� ��K�6�(�mk`^�I�R%��=##��sζ���WM�p=n(�0��[�[aLD�=Q�n�>��$�@�����Ӛҷ=z�hlOH�ٔkFM�	��פ6���h |[jH�8�d�ޑR��p>���D�D��
��Fa��9� �p����O�p32���^[�(x��@��"A-�D� mO�>m�6�Ӹ��D�T�t���^�^u�/vb��#��ɷ"Kp���jBu�O@�w��g��d�荷��5�nz���؞�7 h��n�5.�&M��i�Gt|�@�ڐA�h#���kh�Cw|��r%D��*�T����N�H��"!��O/��m�����=N�nt��5P�w<�b ˈ�
e�w��n�9�mb/�<�;>��UV_�ܰv]u������wt��y����L:�T$s��	6�	MoR21�m]�6��S\Ԛ*ZZFYPi�;��׵���`s������l���oh^&�t�h7[Ÿ���}mXs�`���
�h]��X�]�<�֞àQ����e�U㍆��usyd�5�St�Z��e�RE�޽w���'��)p��l���:�aLKV�!�W\�Q��1M�i���U����}��WE+�q�$%s1=n�����Y{ƶ�a*j��k]*::��~{g�{	̀�[j|Am.v�Ű{fwOB��AZ�f�q��^�7W�tz�nD��p���8.;.�yP��@#:��ވ�������sCbzA� ��ty���bF�v�_�W����^�׃u��r"�\VldS��SP��\j�a���Dp �)�ϤH�Dn!�22΍��вr�&�q�6�;Ib�=�MwOB��]�|Dյ�Q;)� �Z�uȐ[��ۑ%��ܸ�.�*�"7�g��E]���<��w46%/ "�<�W�m�n#��w;G��9y�*`p������-�U�k��^�1�g����ު�Ӫj{<X����'r����|ۑl��
��Y�~�s";��1ٴ����`ˏ:�� ���es ����6:�|�3�T%bҡ�ۖ6-�(Ñ]����~�"�ڀ��]\��M�o��Q'�U�f+f'�~��δ�ڀr�h1j����=�uY��o�����d���zf��=x���w*�;����D�m�Ǌ܉�G̳�ud���a�Q��#��On;�g�� ��G�k��`7̫f����pU��� ��>Ɨ�hL����L�,�=��Dq�q�;�*.25U�l?�@��Cm	�n2�E��(O��Y�J5�N���k�׋� �!���͹3�����}4�p��-f�<�f��m	��\Iq���M��::뭴�F�m��q��~���u��߾i����Yez#����On;�eM�cN�E�08��d/椂h/�B-�>#sxq9u�s�4�Z�ޑ3#�dM:���]���w� �ex���>-��r��*�gJM�w`"�B-� ���]S4�'����>����^���hY���0���n�Տ�����`�=�����N.�9R�Kںr6��א�1P�����׺5���k�hLc���@f��^}�e�#�6��Ǵ�˨��:h�6܉9��A,�����'�s'������!1�K"�Zؚ/���� sA��������������O3�U�1������g��,1�n ��7�br�+6��������|k�͛ڼ]��/�:�玮����m^� g�ueF�i�:gp��4�_���z��y���A]T������R�G�pAʕ�[%�����s@a��mȒ� A,���c]�ͳ�Sc 6�qҢ;�I����έn���	���AB�m���NF=AT	�qz7���h C,�6�E�n�Uh���+�D�]%�s��Ȏ �,��7A�P!�2�7J7:�!'�ºx��[C�L`����¥�:���= �����,B\O����J�W<h�����tL��C�TD0��Ց��zt�f����>z��M�Y��m_��Or���I�p!�u?{��z�GkK�����|Cq�r$��"2�t2$�p�E}�N�g9���lO	��ڒmݶ���;#�-�q���M�5�n�+�Q�����3��]��'��x�@�	�fg}|'�R>�A6��mȐ�d_l��u$�q5���j7*�m&;cH#3$H=��A7mߤ[��X+F�u�gU�
7�Ig �&�-�f+�S�u��R!����i�-��I�ˑ>;��@�A�"Kp�A ���FWEv`UQo�������������G�j���i{4C�棧;v�Wr�}Kŷ"TL�ݑ4�d��&�#�># ��iu�vJ59��	cͻ	n�mU&��;Zso�9 ����>;1\*�����v) �����m
��u��G�pQRsK�yq�&6=�sc!z��(����/l=��B�ԻD�~���ǅ��'��i6����W$�o6�-�V�bמށ;��Ng�e/�:w�����a����hž/||��A]�q]�N�MU��:}�/q/��U����E^8�+g�>����z:�d�l8�Wn��ͯs��>�>�n{&[!��o��[;����X��E�.����zj�w��Z��I�}ӏ�a�e�ԯݔC�Í�y��Т��[K�t��B!u���b��ͧ��2�f�wb�ɱ���NF魙r��d�r�\[hڈ �=��6�K�tr�x�ğ��k@��n����y�R���q��cӺ���w��aC�K�=�麎��+��Uu�t���wgO/"ʟ)����&��˛ԙmj$<���~n��a;��Ƶ=��u���%�����`�E�u�+�!�9J�6�v���,qzz=�wc��"�t�t��c�ǻ����?vOHJ��T�H�w�{5/U�{��7v���iҷz�1a)��p'E�jv�P!-�&�i��W�'�*�5��s�����T��޾�=['�����-�`}=}&þ���ib|C�b؜���n#[���l�nrXmךζ��l.�Z7���l�Ǳ_�0��#h�J�N=7���ܛ�8�%suz��y��c���c�֣hO����$��K؈�w�Y��lܬ�6V�V��ܥ'w\8��^- ���}�ݵ�0��xlX���ƊF�{�Qq�L}Kw$�5���<��_{�.������8֢�r���5���Fۛ_�� �'&ݯk*"^���ԇ��"R��3��!!!�8�"�m	��e����8(���=��[�2�$8��",�����������)mY�'D�m����BI'cknr�f���S��i�D�-/k��FvNS���"-��D�g[�b�����:w����t흞^u�N���&�ve瞨�'}���8�&n�;�Nȃm�k1R��H�2�>{ݠ�4�lY�}�^li����Y��)�$�ڳ�dS�gl�)�M���L�|�H�睩mۥ�t�<�nZu��I(������gnGHۭ2ж�X^S��[��#5%�;F�Q�Uu���5�Ė@ڳN�:��en��q��7�<������:�놣E������wn2l�'rg���/T^K�y}��=XV�:���a��Qݯb v�ְ����'e��F�%Ь�:�Թ�Pr�3�Y�-X$���ݶ��/kp)*�Vq�r�\U��y�xu��4�F�d!G6ƚ��Ya�r"M�i�zب�&�ڒ��s�y�ԝe�{]u<�)V�81o�y�z}�8��3;C#(����N6&��^b`��֣���y�O%�r�cY9�[#�n����qf��v%�e���b�Z�	��@6&�m����$fV7:(���ݓ3)���h�if9��,-����1���m��K���̤X��%3CX�%����a(��ymcJݣ�0�B頊���:����UhM�h{9	;v�㌘�խ�W�95g��y[�u��΄n���:ěK�[���MƠ�Y7=!q�<Fm������G���<��mh�@�)	�6k�̰`!�+[ۏlp�y$=�8�낗�;]�m)�^20t�g%���t�fb���#��R�Lɫ\�H��30Λ��n=vvLE�N �Փ�s.1��<q�2�/�ݍLܸ{>��9r�n���	�m�(7CB�аca�fH.���1�����P��1�c������
Q���7q��r��8 mm�s���.^��[;g��ꋕ�n��h+ t��Y0��*�-p�VB4����Х��Z�dRR� ���J=�J�.J��͵Lu�a���ݽ��L��^:8�&��:#Er8`[3����K���a3f�B�Ef0s�n�RbQ�Q�Љ�%���k��gtSx��
�qnݞ��q��]��N��gn-��E$�������5vBf�D"�牜��9��u�9���:�Y'�3n�I�	q�ƣrk.��q�e�u�ٹ�I��Y��ڵi-[j�t��mT�W���{���u���Қl�q0A�IYef`ɢ�XS[T"�qY���* +`���Xv�B�5�WCg3s 5,"�4l��q`�R[��t�������p��>�9��\u��=���j+��l�6ai) h�2k��b���n�b�f�`�ɫ��6��Pqc���"{�6��������l���f֗v���v�F7W�־�0K������� f�x�OH��ڡ�x�J�N���u�Ы�rM�˛�pe�|;�����__?i�σe!�����z�ݍ����5�j���w#٭_�-���H�a��2�\�B|}V���D��Țsp��&�#��ݼ���(�y,vhj-����۹Ǻ>n-�$���]�;{$=л,���p'l�=θ��S�ǃt�|ۑ>-�"��%G:�l*��3�"|[�A ��J�� ���:�wcbxH%�D��@��WlP,�^��x7AmI��o�d<|�dJ���$M9�X�wY����;zD��x�CqqԌN�������(鶖�pY�͆�5t��tn(���;(�ݧV���:�R�^�ӆs���E���ڐAm�&���`OY�z�@����R�*-�E�����}�m�`�@���}=���q�<T(WzFn�Ǡ��L��"G�m�����%}m��Á�ߙ�Uz�x��_�������|fE�k�%1�6�ｹ���+G�9����J��Qp,΍���lOH �@@��[jrD�0��b�M���k�h#��^-����Zb*���wz;vD����q�5��1�v��q~ ��/�^%Qwu�_Nt}���d����v�1��ޅ�}���X�YT�i�1'��^"�dIn<�n<�r$�vj�1Ϧs�*������n����������mH7�+�D��"�B���)nݜt_�|���]5��m2�D�Xk�(�#�P��`�{�kך�>�^ǫ͹L�ݑ4��b9�Y����9;�/�;���>�}�A,��mϤ��Fa.c��6>Υ��pM`ԣ��G�zf�����YM�)U���!S2$N ��O�n|�Y���w�`D����-��]1�eQwZtNf�zl#�&�Mhy�-�m(��sdU�b7ȇ+�T���9�Ʉ������(�!M�Υ!��Y�_��xxt'�b!����wCb��dA���m���P����8]�Ϛ�qj<[r$(��$(v迿 �?�GR�4\!�ȝ��G���n���D�[j}G�
��O�ZaN��K���/B�@ �b�C�.�����wG�f�*u�����Ḟ�c�
b��%� mj�هOjۮ�c(��0�I�*b��a=�D��y�+ڗs��Nv�뻡�|$T�;H�X��j �Dg�o)�D2ף͵$h��;�2(ҏ;zD�"�fM9�Q�;������!�����o�'�sT��lq�Ex����������7����<�UF|zy8��3Dp9ا���.�ŷ"|[���zG���Dա'�ŖP䷞pd�l�t�<g�֜��d�o����:��(��7��T�o/q�%��,���v�eR�"�e{?oI!�XMz�}Mh�}ɔ�+#(�7u�����|}���� C-ڒ�����u[�̛���>Q23:d�ͥ3��ȏw�|���q�Yf��wa����L�)\���P	��ֲ������.vy���<M�� ̩�Od�ΐ�m��C�Mf�K��Rs9z$3]{���)��^� a�x��H-� �Y@�&�Oua��� |��o<%=����z��l_	�@@���"�[}ZN�2�F!�H!��Z�x���S��-��"qe�1�2r8NW�>��p�$7mؑw/T�".c n�7 _�n�oW�͠���).�n*r�W�@�ؤ��5;�o����^8܉-���D6�In+�s�E�;��n��x-c�{�T6-7� ��ڒ4��]L��9*T5h[��ORɖ�O5�
'�E�lWH��d9��\��5��Sq�XF�μ%����2�՚�i������<m\BQ@�E2!ژ\�y�'����=��s`��}m�VG�Ѳk9㝇��:s´����3�)cK.��̎��6�z�<`v�n��P/V�5�t���9�K�44͗]�j|�v
�s�(���9V�oa��X�� \�Y���k�C�V�1ڌ�r6�M�^u�c�#� ��fyvz��l\�'���1���b�n���}q���īa��%�#wX��	v�Mg�v�9l&`�,�/�eJ$����ͯH�^��m	*d_l�k-����Dp#-]@k�#�m��hH=��$7m܂p���7a����H=�����).�e���:�%�)�|��-壴�s>�ˑ&� ����m� ���)�AK�r��=\�/�Ѽ�<����������>�*�U*�M�w�S�)�sP@��^>mȟ3gvQk-����Dw���78�U��7,p�b�\"t Cn@�An �� [j��Q��&`l�^	��c������p;��)!�|�y6�t��ܐ�b�U0�J�2f|`(AsC�D���[լL���Ã �kQQ�����h ��^��'ŸD��y�j��v�N��Pؾ���諙���4Vǭ�Am�^@�ڟ���ֺr�o6��m��>�6�\��'����?g�=Ƌ�:Af]l%g�鷴z{fx^�'�����z2�
_ʣ�}��M~���<p�o��1�33g��y6��q3�A!�����p��[�[1A=��'���%�Ŷ�ChH*�C�\F��Rl�QuW�o�� K�^���K�6��ŐgF�J���O9��@�n��y�U��N��Pش8�@^>��[�|e� ��6�>-� [A7�����-������\�g(k�{&��9�JȎ�� F�!>�@Hn.6��nd�V%B�IҚ���Nбv����%�bJڻ\��1�n+mG�9������9��mH ���k4���uU{��＆�*�!Uc��G[�R4�G�P^m�%�D�E���g6A.}��$n����y�U�/�wj�l_	�2 ��m���r،��Z@��R!���z�nE������N�Q��=h�a�S+o.ŉsKhPY�[�g���g���F�'=�lY�6�gRŐఄ�w�T�K{,-�+��cc��2>��vk9E��X'>���x�Cp�>���� [A���p�qU��=ً�W����%'�xS��Ô���#-���W��5��tm7�g`%�Y��Պ�fvҼ���ڭ5�]�v��^�a䋮�yq��(����)YkWe�#�����u�A�gJM��f˱)Cb�&�D������ۯ6�Hݔ^M��s�'C�or�lP��z����T�ݏ6�m�V��N�Xհֵ5���XSl�O�����N���>�۬��(͵i�T�5��u��m�n)�|�Mfm,�n_N���\.�|��A��m��ƫ�Nbv%��{[^��St7e�h���'XО;Ū�����r,�
7+ĉ�˨'�/I&C߇�}�ď5��!�['���5�'�'�_+�y١��o��(�p;Y}!�3ZEP�W�=�y� }�6�7�۞Õ�b#`}�M�8���17z2�w��kϡ�۝W���W�af����R$� ��;0w\5u��j�M�i4!��]�1��g�~��7m��u��,�m�N���\���lDbB�7���6۠�Ca��sW
ą"�wv����E��8';��Տw�7�-T3)��n@y�Ǜ@6�m7;�X�oQlHm_�;�]B�є뽽k��6�m���n�2x_�ǠfZޏ6��Yٛ����:��Mp���u!è��\���^�����m��9���nݩNV*�u��Yh�Y�N�k�{��p��*�2��N.�a��݇�AD��K��8�޵���v�>٠Y��8���{
>=��k��7T>�D�o�2��f�z�z@/"�wC��T�۝˅���=�YY�\d�vNl��W&x�S�m�q
�
':��u��᪚�AmV���k�<�!�
%�ac��\h\�񋫊:��Ѐqf5��R�+HH69	p���
`�BZd.)��G�hM[�CY��Mc�0XH���n%���-a�0nr�i��RYέ%7m�v�8�WZz{N���6�s�n���w���NӍ�bu�Â��i4�R8����vX�<s*}
bV��{� ��m��
i�ձΡe��u��[�GzVhښ���͠h7���f��[St���@>\�;b^��k۽���x6��L�Ҫ9�O�<���6��m���Z����gvf��ܸ82^���%��7A��jI�sx�E^����֌�3ձΡ;ѕ;�]�5�'��%��/^r�����r'��ъU��|��x�6^���z�=��O�պq�W4	���D.)v�j8��V�!5Bg��֩ϲ�x�gNqf"�$HS:���3�6�wjk�l���1��p�6���r��q������7���k�3����M�96�8�͇�#�j���#��Z߯iH۝�]q]�m[\OQ�ʓw�"G6��E����?x{�m�rw낯4�}[�'z1^�޴<�gt��1�01�qgi���Z�my��n[o�A��]ξ��y�)�^=͗�zo���s�hy��1Ar��%ae�P3m�SU�L:��r{�Ó��R��4&������6�p�A��7Vڸh�>*��9�N�b��oZ���m ۣ�t�:�8hH%H�*Hn�5̎'qu���t͉�o] ����^�4��a��K'F��z�n m����uM���l��f��ݓ��@��{y��6כhgf��쀠�ۤZ:�{1�Jj�bIj�bȞ�p������wt|룲4r�*��<�M��:w�,��Δ.����=�c<�D����n���*����^�]��Cvb9!�����^��A��n��Lכֿl�V���A�K*d�f�z�,D̳���A���d��;�}z�_�-G$U�=q�>=�'�s	2^���E�7ؖ�D��`����+a�:�Uꆫ���@x�??^��[6����K��ӂѓ��t�Ƭ�F���������k�/q�+ބ�����x�Q�y���w�Kwl�ȷw�Vl@J�.��r��J?{S�rG�L��u^}�����7���C��*X��+�P���!�(�ڻO�l�Y��'��z.v9������ވ+�^��ۯ��5�p��o�~/.��U�x�"���	�;=�K�����}˔����p$���yD�#j��nvԇ���;���=w���՞�uݭŠ��;&�>���у�ᛄrl��/q	����0�1XجQB��zqٳ��}B�Vǯ�C�?Z`�w;��9�؆ã�6Ȯ���g1�����K;����&�}(隧�7�κ1�l�YxgB��[8n2���C�6uY=9��#5/,�i�g�^U���5:�=���L�����p+ڏ���E|���r`���l�d�|�,o:����&{�}�p����؛�O�ƁЇ�]��Sh�T�ct&�ej�my��s��}�����X�)�{�Ց�W�Ǟ�F߽dcv䜘ǻ����aO6�b4�%yw�~��.�/���,<VAyym7i{v�jp�O��D$�눡9���wY{w׫&�Cی�=��)�J�w|�)��o6���i�ZNsȭ8�˙non��]�YZ�ݷ�]�>֋�E��}�<�N󵶳[s]��m���C3mY�4���$�)ͳZ��e��{��m���mm�s�ך}�f�Ît$ٻyZy��k�@S��^�;��b��H�ֲ����mY	$��m�K2^��!<������{-C�GAܝ��{`��m�j޽� `�kp�'m���ﭹ�9�'����w�h'�INe����go{�̳rM�$���֒��r�-�i�bHL��pm͉�[c�w�^�`�{AQQi.�VЪ��G�+���{�����{���z׃��m��q�;:��P�������cf�x�콻f��@�u{/u{6כh7�죽��(v&Y���j���fLK�p��|��6Ӿ��ي���Xd�H�R "�U��F�<�z$��כ�i.fB��c�ۊ�m��nc�����6�k�nj���J{O8�z�o�Het��t��Cݍ���i��mxB4��5��Ok�������{v�;�q�z۽FcY릸ۙ�'9�MǛh�
��곲<�dĽ' �7�ۏm��Рw��UsW�]�ל�nj��f+�c:=y;���/E�����Ȏ����0Z�<�������~|r�xf�^�[3��?M�yQj?�4c�5��`[�P],�
Oh��_eH��bre1Rl�)����/�C���i����7M}6����M�e㍺-���������^ГX��;�iG>~�;jg&j��:��9��͊ݻ:�^\MR^�-�T%2bDP�fG}w���jҪݔL:ȼ�?q8xN�C����u`m4�<h6���=�(Q�o��_jn=Z��ˊ���³^EN���'���_E��B�r�t�@6�p}�R��4c�9�GX����ͻf��q��M��7m�w3��tmJ�F��{z��V���S��������9h<T'7Q�DTD�W�/�m��y��}�7YY'&�
���;�`g
�y;�� �h޲	�(�y�~ǣj?�x����B�!3y�#;�x���d6�Y|H���ۊ����燵癸Ǟ7��̳�B�~F��f�"7?{��#�D��H���x�l��!k�Ѹ[<�p.�z�t�n8�]��܃����g�!m26���mt���EOi;;�[��l��`��s�s�>�[`�눋F8wX]��e��G5��\�.�������%���IO����ua�;Y�D��]��i	��	k�݅mn[��y�I�sg:�v�L�i�����
��+Z��FC����~~�p���E��[b�����ݮP	��r��XBh���ݰdʙ��xub��Cʹ�y�8��>nonٵQ�a��=BW�͡����m��C'kѹ�ؤ��۴�nJ&]U�K�A�ޜ��k���.���Qn�u�n�k�ֈx����mN�<z)�@�����}��c���m6�t��8�jw��^nm�����v��s{v���t�j�2q�N��P�͵��C��m�O�;	�}��hQ�N����%�������ɸ��weܚ=S#Bh�38Jh�b雍6qe
�9,��GN���qr�g���DB����r� �A��Z7�K����Gq����'���>�4������MǃmGk'�S\��q'.�V�~�^8����[6���t(�6��n]C�^���@f�^�����klZ���9�#@���ix�m@����o��@���~w�6�<ǜ���q�gkmٗۑ3��-��^B�Z��pk����rx:����	����1;'
�C��7 6�mϙ�ˍjD9�S�C�٠3Z�p6����u�Ǌgx>�Ԍ_Ws�E؜�6��m��Ę}Xvn���S�	ck4�*�w�cc�s[u���q��m���qoEz��M�lD]����tUۋc ��ڹ�Ί]OYt�-g�
RP�(��N{��m��������w�'������3�C2��y��h�7ІFs��9Q׵W]:��u��m�]�N�p�����չޡ1Ҫĸ��͵��s`��>}fʱ�z&�J��}�p�G����e�"1@H�jl�_п�Cx�a�U3���g`��]ӑz+�sʭ��1�}5�8o��|�i��^�q�"����mt*�_F�ܴ���i���*zN��J/q���w��[��ۜ�m �x6�m�#Яuﺠ'�X���Nv�nvk�v/=m���Rj�usy����GK�t3\���M�n{��uc���]��iL�RbeLD�s��zޠ�6���c�ӏ1�t����Gnk��o��.Z܃m�ۺ��sJ��Bw/54�-k*�g='xVb s���~ҳ����v�v t��xRF�պi�[�"�t�s�]��^{m�6�n����f�^�׵�����qZr�����Xo��>�n����j�F���Na�M��n�*���.ۢ�)?ޕc�2�]ut/�uc�����y7��j�f3�)���J��˓�/0���k>���m�7��ꀖ�_B�5�O^���n��XS�p���ϐǛb.�IvK�3����ߴ�Ia������g�x���`���%7�T# �bT��T)
Me����c�Ƕ�N�r]�B��s�\�:ou�+F�Hͽ��m�7 �
,�s �(����7�c�ӕn�W^��|.�7ͱ�v�,Y��FE�Pm�ᶃn���Pz�>�D���aOI�³>A�m�hxmƆdɦ����9�-ƛ��bv����N7[5���,:�Q��šX`-�/u7�m��&���͖0�Qb�Х|�6�F]�y={K����A������wG&_I�W1]T�nM��;��h���c���yC��&��{�2#C�u��Q{.��ؗD�;�����;���ke��{�$�Ү���hq�v��k&���<W]V���T���cn\*�+oh�X�t�m-V[�h�E�� A��y-�ׅj.��UI���[������������+��(�>]ʬ�&Me��łGu�V\��+�XXP\�꒨kQvV�h4٪е�f{Xk^NX.�X��Y��Kg��U�pu�c���5�ϖH����K��\:U���#���WC0���;su�YQ�Y38c����(�RJΟٟ!��mx6З3�������)�6xWL�1Y�wi�}��@7��T7�v��ѝ�;q�>��M�[5�؞��LQͻZu{���m������Es�x�ӌ�v�u�,5�pjm��j�lhGjk�^h����igZ �ws�.��<=Y� E�7G�fT=kʹ����rop���j���K�*��/j�;���ۼf5���\�V�!T��J Ưoԣ�u��$��k�^��=�t�j�W�����P��6�o;�q�ݻk:��5ʥ粢]楘.�H�N�9ᶽ��5��*����r#�5Fe���1�:9p�mK�gL�7.��Y2֦\U��̋��S��[����&k�&��,��ir��=��H��˺3u�R�s�Z������g�f 5�n���%]̽�k�<� m����s��"�����rӭ�ᝈ>�kʹ�yg;�1ϔ����^���[��jwn�ν��w��,�j9Kx1Ǜh6�nwT[B�t��+������c�%Y�Vb��7m�ӈu=/X>����;e&n*��چ1i]�S�ř,��\cS�!�h�S�
a�ĥ[l�6��p:�N�$��۴�f{�+zft�b[�y{�mכk(�dP�uu�J�f��ʺ���ݵ�{I��]�}����,R�MSsN�q�A��|)0�N�Y�m�@�F'�g����p��U�.M�o� ��rSg��MY��h���P�&�����Ա�-Uщ5q�tL�=����N���3�*n屳����1{�/7 6�v6m���e�Ϲ���q�bv�'u�n;nӽ���UFu�6��*�^��m��}1�F�ܣ��W,�y]�۶��i3]��}���b̍�{��/h��={��Y]����ƌ�B�]�l�^�GX����uB3
P�dJ3&�����m�6�9���Sw<�NJ��	M�uNv�2�?�^�ʹ�^�p;et�1������{:==bv�'��n;nӽS��؇�6�#r�;�X�����<�^no�N�L;-f�<�F�uw���nof���\�{_ �@7 6���k��W��r��`n5��8Y��.��y�����^ /]Y^+�^��^���, Vm]N�(0�j{y΍N��N��]C�W71��x�}��{��QV]oos�vyz	�$�l��g�S43�y��n m�ڈ/N�p�hu�n6q�[S��v�m;�=}�>��@6��3��U�7�T��<p�i���=r=ʽb�{�j��N����5Q������y��;�WY��]�yղ��
�M
�w;���yΫm{��m�|)X������<�@��59�.��y��ޫ��M�V9��J�P�W�~���m6�n2����嵎����[z����ͺ���nf�;�q��&w�=�6�q��)�sx^ul�5U��^,&�:FU���۱������q��Vr�R�k=Wj���­���n�w�LV� r���R�V=�w��U�b��W/M���A����k�闟q9w{�c@��,[oi>�oi����*^�5x鳤�2�d��a=ˤ�V��1����pzm�J}ǩfv���S�<=���˦غ�@��M]�kME`�Oa��wv�S����'�����l�7~[^�@�>p���uM-w{~z"�ڔ�%;Ua�ܘ�o���{{ �_���m�3�� �K�ߦ��8yX<<�
���|=�g��=X���>�}O�G��k��M^Ye�{s�A/g�P�T?y�y�䐯���n���ny�'��w�nKw�Z۰|}�}�\>�%&�3Wv�+�~O�˶x1�!�W�����;��t����\1E�ʐ��۹���05���`U�:a^�0�MЅ�(;P-�}TC��y�/��&�Ƭ�{�wA;K�F�S�6 n�{�Ĳ�B~θ�K�
�2��cy�A+<#r���i�Q����[N�:4�܄2��xx�=^u:��{s�؍OQ�7tzq[�Gd=o��p�M�˓NG��Ǟ��Nk�{$�G�uYn/=<}�>N�׸�g�N�²��mY���'�w	�n����u��������KE��;��y��>;�|�]%M-����Ӣ�XG#6oF�Nu�ƺ�ޓoq;9yQwWC�;Fz�OwŤ�@`��n�\ZЌb�&Mf:E��`L`�a?z/Hƞ/o�[��-μ|OÜ���5����N(��� ���	�s%l�D� �$~���m��!d�׭�"dC���N�vH8t�=����n���Ͻ�<�)��T�{��5�8$:��^�^���i{�,H�(�,-G�K��;����v�Ӣ�Ҏ8^k۷�nzÔ;퐙om^5��(I9Ӄkˑ�j(_j٢9�}��V��^ޯ��Y�fu��l����b^����$�f��nԃ�n'��k����L�N�rVpZE'�kB;my�Yj��;��H|�98\�vX{[��>�mѕ�z�r���a|�{|�$�v�۴�����}�vK۲3�v|��۾ڝ���}�9��筮I�u���{��)�$��Y��+j�{���v�������!ݵg��tv�IK��@=��B�v�v���t�em(��8����u�fPNs>�i=���e�aY��O�r�SZ�Rp��Ҷ�㵻.FQA�*�[��F�Kջ���,qͮG�/p�ʵ�a�k�v��`�N����. �J�P�pv�ʒ�Ķm[e�5�*���fn�̸��i�q8:*�Bj�������l"^3�Z����Ɏ�y��p+1���7(Gj 
�!��{V�Ů#��n��|�a�s�q��:�dh�잻Bn�vZ����Ė���N�W BioT&%,fY�#:[h�u�ҥ�8f��$�]��X�69�7��v�
�r&29�ݴ��DK(5�Ek��&�p]��ո��A��&���^k�"�;�������أS���~o������Yd��Ѹ�XX�Ё7E�k�es،�m')�2k��ka�vб�(MZ�� �#�0�i*�3-.8fLݳ"�M��[���6�Xu�5�0�0��"[���m�6�#.��CgL��d�P)�.ePn��\y��G�����yd�zfX�m�G�r�QSq�����S����m�/d���$#�v��l�YLZh�I�F:hF��Ѱ��4���]5Ě)��k`k�T�M����)��#K����ޡ�-�W���(;'tlv��W��v��]�=���nI.{,(<��bSmu&�n�K����3]n mE��\	�vx�;�Қ9úwRÁ�7<��ls[��Qnnh��<�=:N+h��;s�[����E��ux(�:�8\�!+[n�K	�X�/^b��)%�Z��5�&�3ZV��e.J3\q�Y='*n�l���)G�]��!�nݮ�أ�7�]6����\��3DE�)� c&����c����f���2d��N�i�Ʉv1n1u%rpv{3�u�(���B.k��ay�M�t�7X۝mD��H�� ��g4k�=ѥ����=FG���+Z;p�m>�O�5tu�/,&J㹶��;E�ge���8K��H����Y�.�POQ���j���];r��3����h���À�ؒn�����;[���ؘHQe��M���g��ny�w5�L�%ٞ�*-�����c�62!�����\�⤎V;v�\u���a}kn�M��b(����tל�m4h6�s���)A՚1�m[��-�Wc��b�f/ ����SIcƛ4��P�<\��r�Q��L�p���C园�����3�sv�.��e#17����ݣ�q����B�HQ&%LA*�����΋�A���{�o��۫g�mm�Z����c�=Cʹ�6�z�Ss՞�����+�� �=���x?��~���{t����VR�k��m�۫���Qy�W�q�]��+������m|�q���l]�㵇��2���������F�����+��^�����w39���f��\m�2 �������r���P�v_N�5y��gMp�����`w:�����u䱗ɑ�b����!����,�L�GL�X:9�t@*D�H�R�I3@�h�d�̬�;E;7��[3���X��9�,�i�u.�7�ِ31 3 7�/:����*
����y#n�exa˵��N,���[*k��ݝ�n���6:���g�{WT�3���LM����U�2sM-���7�޾���7�7��L�m겻ն�́�T���R�g^U�i�n�r��|4�7�y��^�����~k���C��̶�֜�N:��q�%ZΘ�U@��^�sG�%���<-ųx+W_��wFf,�Zs-�{^�����k+-�bw�+�|���Y][h=����3;3�nCڙ�w��g�� ֐�pi,�)q6f�Q����d�!,FR���30c_��w3(�9ugN�7x�N�N����&q�f\]p	�י��36���ɮ��~ʏz�74wR��c�r�p5��0����DV��nd�b�Z�bqԣ�؞��'hO�_+*���Խ�c������,�.@���M
����AٲU�RF��)�f�p��b�Nh�B�E�sF���4�z{`���7�m9��^oӿ��>�5�C23��:7S3v��ݹ�<=wڄjy�u`��^�{̀332�a�E�q��ē*�V����}���g�N ��2=��z��\iP��d���<��Tm�q#N�}9��+B	�es*������]��=}��duvQ�]�S��;kU��s]���OD���gS<s-�i�N�Z�)صFX͏f��[YѺ��x�'�:Wz��ǳ3;�K��;�û��df@���|���rN�~�Է���{�7��wڳ#�33(P�ܪ݉��@fl�I�]yS���֫Qު��;Rvtbj�l>�]�[�v�U���\��b���M ���򟘋n�N�:���1�w��Rz_��K�����g����m?Zr۹i}��ذvyʋ�x{Ps�������3ˡN��߷W1N(� ����n���c������n���4�]���&�.��޽��_���f)r�;�L^���Mi�{��6N3�;�ǆdfb��3b*��ޞ@f��I�U�SΤ�֫Q�\���Z۲ �����l�3� f�̽�˺�u�y��5���Q�]ǽ�f 2�O�ӡ q�M�K���m�\��ۡon�>ݙ���:wpt���MWm	����-�����X���9^�/L���^�&*�UΑ�V�����̏e����AXȌ�v�]�֪g����F�qgp�!c=���`�~>�T�׽M��o����F������颓9{>s���T%4��=/�w�Zn�K,7�P�Kt�	3F44�
uqѲ%�:9�ڭzx��Ƃ-���X	vb�젉�c�3��ݸ�٦/f�h�,u1 zٲ7k�����i�նq��=��Wi��Nws���]es��gu]�\���˔H������y�£\e�ے��λf����1cqP�m�&��v_\�tt0u�N��s`~��7��t�p	���yݮB贪�8����kL�l�gn�31�/������㲸�A<y�����#���=}[7h�:��5{23 �]{�Sn�X�Q"w*.�v�e5��n����Σ��fW�b'b��۰3#�/�bX3Q�]�R�Ӝ��Kj��j�<����Z�-��Kqo���r��4��`fF5�|_ �<��v�p��)��޶�+����쁙��36�g�&zt@S���	��Ո�հ�n���Σ�چdf�L+��"n��;5)H�)AE(�=�m���^d���p�e�Rq^���9.c������x>����r��ʞj�mj��}}�k�����������!*�K���̨�!�1� 8Y�<��c=*�W�;��-�wEHK�y�d�x����c*��O��OU����|�������w����c]���G1�>[�8Wx]�큙�uk��vY̍gf�kk�2=���\&jkzo���͌FV&�ת�����yfFdfbm���y�{�L����d��7��*y����uu��{��2��{\z���f!����iZ��^��/a������.���f,�@W�m���럎#���KR$%j?�i�(���B�v�Ү��:*kf��]�ɒ�o������ᙊ~s[������Szy�IV��c���Y�&���lNƍB6ڙh^��I�]YS�X�V��]h�ᙳ�F��磻��n=��ِ3���ͥGr	 .��~����ݮ3隭>{ȏǑ�8U�9}�y{~s��6u*��[�B'N�{Tᤡ-�^<�M�1�z�6p�w��^�� h���8�[�ZL*c{3:���FS[���Szy� z/���55wWl�s�O֛n�J���w��dv�X��V*��;V�Q�WZ��́��u'f�Vgv�;�n�

S$�ɔb&d	31Fu҅��r�,�4ӓ�vb�Ћ��k�d��}7�O�}���́��������|�6p�Z���1L����d����6�t��DL{�<;Z���Q)��x�m�ɏ7��כרz?���8U���֛n�ms��_t��C�dv9��ŷ�Vͨ�����d{3́�6,�f�7�9 Nw:�����i���|�6p�]��qw9� �o��tz�vyyu�];ot��yת� }W������`�A��	�8y�o��st� =a�F۫�T�UE1�]ŴHQ�+gu�Gm6��332�d�R���М����vB�����fN�:���[j���-�څ�Ys����qf�v���(��o=Q"���-f[Fbh4��3S�^�����C2;�p^t��b��f�w��bBFVs�9��^́����qsٝû:/k�i̠ᾋ{8Wuݱ�̕H:���L:rә޻��-9��X��0���w:���*Mn�[����P7yf@�dfb(=y���������U1���jٵ+����̗2�u�[C23#ٙ��"�,�Г�U�޵�7k�8��[�{VW���f,��N:���YQi�H�>��^�1ݕ�-H�K�BUמZ(#�B���t�sMuj���V��Br�V�;8��t�dH�S ��ո����H�5�N��kCQqK�k��Ց�ʎ�|��	΍w=e�Nƃ`{rT���p��3ոf(�e"���s!�8�u���{���4Cs<��Uc�=�.�cn6�6�ڞ Wa2��^�`�Cn����
�0�p�o�����5��[�B�i�X�:;��X�ܛL<�Xn�[�Q�DL3sݘ�)e����Jki��œ��T+�<�A�����~m߿��M�ϴoVc�!w(�n[w:]MCq�H�$�F���D%������i�o>��f�ڴ�a��p�JL�T	���ּ�2@����Q���)��V4=������3v[6��u��3!��м[��ܪ����3dfru\ݭ��}��[�q���Vg���31f@��0�q�ҹek{w�dfb�Ӛ�5A��}�nuw՜��3'xo䦓���2���~��i�pR��b�g{3�=�l[ꩋżƭ�Q�ּ�3 fd�;��ED�.���D)����ٝ3vcB��8�J�q�c�>N���CL��nHS2"TT��Y�f@̏8�ם[�[�O6���G%������|8��@f@̏�]�\��\b�"�bb4{*Β�OxJ��5�q��c��	���^/:�{L�[�9c�qgp"5�w�hN-W�k��1���OX��nS����e@��\]�07�t�5ǳ fb1���cn4���MѾuS����Qޮ��fFf!��L�7������{��]��[�^v��Vg�����Q5$H�K[��N[w2���v�������z�W\���)�����e@����x����{�c�1��e�3H����e�D�i��F�uZ��>&�"gД	
Neo�s�����z��3g7����3"��Q�yW�Q�3̌�$�}o�]o]һ�l �Wm�F��q���j�w���љ�,��q�rX��t3�xf@́��#�t]FU�٭���t��w�1?{��<�Z�3����7���yF��o�{(ΊZ�sُ7fbF���n[o��{w��3sF-;��C��j��|=�����'��Uaw�JiQ�7���7�&�uEji�~�p�k��=+��E��)	)7��v���k�9T�&E^)EJ����ݙf���Ax�q�r?y����#�+�����˨@+ò�Uq�w��=dµZ7*kn�N�2X�w�����&xToHs�Y�u5�i��>��Kn����t�Jӽ��(�����\#_S0�j܋Ь��+���8���+�d�z�zy�Lܡ�E�XZ�?T��&q�,܇��-�܉�(9CE���>v���F��:�)��ކ�:���x�|�Խ��f��N���Ϫ'��|g����m�4��A�q��ˡ?l�1"�t�B��4�7{|��ƅ�'�
�°Ů��U(�T;	��n��F:�3�;�����������y�,�r�=�N����_��E�Z���y���{v�{R-�0�xZ�#V܉�����77m���H��Y���T���/�v�f�P�B^3�z���⻴[�ٶg���V�po��#���p9��f�\<�j	�us��w'=U��3����6���󿝦�4,��qnBU�F۬��{;Dv\Ӎ���3��Ƶ7���w8=��^��y�>�)��C<�=@y-�۶z�Aħ��'�E�y�����:�����y_>Z�w}�2�^CѬP�Q�&�h�уA'�";mݢ|m�����D���^XvvrZm�DAǝ�E{a+mY�I����[h:ó��m�w��V�ge�s��%fm���0۷m���Ō�A�w&���.';��gzQr^vef֜��8�L�6a���N��L�u���9�����M��D��8�2#�������� s�vg[�2�$'Y�E���t��݇{u�t��ݛu��:�M�vYG8�̵�v�yivy{7h�f�$Nu3Z9g��۴s֐���Y�br���h��Ͷ�v�ִ͎=�����[q�q�i(��rYdE���kbN9�.mi(�mڈ�qX'Y�5�ٲ+)�y�l��f�Y�z��f�B��VYٜ۴��ӯ4�r����wkh �I I��בzTRmkm���=�Oh��$crՊ��.^���ʁ�ٔ3 fb�疷�����3!��Y�B�ξz=���>����왾�'���NZ~���꺢c9@���Z��;]f՚�L?~�mv�����;�`�׆iËBu�0���<���75(GGP���V�[y�!�mI(M��h��f/��`�������R�a½���;|����fFf 3 ���US�t��y^Q�B��=:�"8^�ޏ^�p�R��V�twFf!�3Q��꛽������6���zf/fG�"D��F����Am��5��SZz���^�1���������io���L"HF����2Cs�[�M��/i�~�����.Cس����ЉU~Ɋ�����ӎ��!C�����Aւ�!�"A-�7x��|}}����� ��7��w�����|';��G���_K���O�>���j&�WM�M�-R����n�GqX��kC6{sD��L̈12#�O�z��9n���������]k�����n�}��A�l�|Ch"�"-�����5�T��Lp/aA��>���ɩ��T������ Ӏ7�B�n&�۫�~����>��@��ȐA��h m�O�A��N;M��쎉���tgP��q�N�ϡG����ty������\�=���� Sޑ>8�h/O����q�،�]믆Z�H&�"������g��-�[jA���q5GזlW�T��|����tk���O|�N ^��D����34�iE+}�)���딁�,n�}�٫Ǆ�;��e�gtfZ��͂+'pj�۝Q3\߸����q��p��|�(c��.���5w}�w��$��$�n,�P�&�%%J1���)�t*7����[�uӹ�c<�1i��Urn6�.ڳc�)�9dQ����3GX.��u�j��X,�\�u� A���\̹�����˔�r�iHQ����ѣ�|�<��x��βf�nz�m�qM����bI�س;�K���ݓ��A���Fg��5�Bm���cI���ͯ��}��J[��YƧ��y����Pͻm�����_/\��L�	�C�f��m�Kh/���m
�1���Y�B���~3�:���ډXA�A� 6ՂC�[���wn�f�h`�p�A4�w��}�E�}����-}��D� �Clwg�V��)�_R� ��RCp-�>m���>{q_BS�15;p������i�^o|��[�A�hb�\/��nR������sP^#�ٟ6�ާym	�1�N�g�G����A>6>S�,m�����ڼ��n �܉������i�(!r����e|�si�2g�$��P!�#����V(���]�TG� ���/���W!���Yfu�ͺ n&Bi����3u�w� )�^n=E�����Mm�G��\'�/�f-���O#&��
 ���$�B���[�}װ󯵋Я��Env,�m�ZNC�y
�=k���*z'1�ݬ���4oyE&���^M�{���'��Ͽ��4�cYU�"����;�w�-�?f}�����%9�/H�����6�V�~�Vf����l An M�p� 6�����Ϊc��鲹�N�k�o
��ͧ�>9�� ��@6�O���[�C���1A2�R��>�"�/6Ԏn����u|'�@�pW�[�
{��~#�݉�q�����w�7�)���9O�f}�����%@9�)���"	��?c3���{N,HW۹� ���)��:�K��d�����]���ߝ~o?0/vD��[AL�^t}�Cc>�{9��_zB��z��Lm�áD�}܂#w���Yn ��S�Wŭo3a�sF�@�s5H�������-���W�z=7�7�BAn6'j��|�A G�9�}Ј>mm���B��ô����m������f:��gˎz��N)�#�i�Z��y�Rs=*��a����}"��k��y�c���?.��Ё�!�Q�ro�&�N(������ϒ���g�H>ߐ^�G͵ �hy��n���R� h ��9��nW}y����}���������d Dҡ�����p�{��n�%��q��-��ξR^΄c�}�U�&��`xk��\:�Y -�In�2�MpcW��D��I(��B�#���8}T��
yҽ�G@Y�=;���t71ʝs�����@@���p,oK���Q�g��v2���&s�����sG~r�n=y�Ŷ�ݠAn"���s�D`e�y>A*����Dc��[�����7���/ۺn��5��:LW�l�.�x��) ��^-Ǒm��7��Ǖ}�q�᭽���� A���߾^n=m������������A����G:�Uj��>�����J=�~jH���ᚓ�Q'�u���H�i+y�_O��;�}��7��v��vw7��l�}�z��!�p�%KP��V]<yf�����������pmy�ۭ��F���jsz�~�11��s��𻟄�o!{�o���|�������������6�,)��y�5����Ӂ]N��=�.����<�@��A�"-�?k��&�{xk�W�A_e�3�e�V����[As ���}���(��O�|�.����_f_۳��>����o���~�+�;ǲԂ6���Dۑ>���72�8��	�}��:�ru����]���� G}x���כ��_§��ߦ�D����h#\�G�-�=����[�%ᯭ��u|��!_�3��gË���8���Cn} ��@mm�K~s��{�/�C嵝?#��/��k>�N�����@�[j��.�N�������2�&M�*6�F�uۗ�55��;22�D_T�����R�u�P�{�(�����FN���"�>��
��mHݔ�i��kl4`F�ZaW#ʒ�'l8��e���:toD[uh��\"��I�ϒ���M����]u���V#Q�]�1k]v�l�Z�Ժ1���λp��'��n��ٞ�U�lB\�	h�u�n�eb���!�"�v-�����C��97����F�ծ�j����pG��Ȼ����A�Ɏ:�[�c[�`�e i��m~��>�)�[71�1��eءy��C-�%�n$�ݶC����(�*L�#�P?>愂�/[A%_}�_tc��캽��]�
����G��{_F_ ��"|�q�mO�{��s%M�80�B �֤ͫ��U��X��毇L�o }"Kq��g�s^1<�^#/�H �Amm���Щ���kx�'k"�n�T�����뼚ϥG�|w�^�o�/�x�my�C0f�(�������r$�Cp�[�u�ю~����o�w(|dz��Y��#ﾲ՛��#�&|~�-��R>mp��7���eemh�g�S�m}�������_��\��In �6����V��\�=}�\�0��;%AѦ��kti�/-��n5�i.�m���$v�f������Ͽ�2ϟ>i>!��}M}���yu���9���>̕�Ng*VA��@�Ԑ��� `���Z��o�0��U,E����Fm^�,鿷{K]ҡ�2��'+��v�	H�(����7�S���n�ѐ�+ڧ�EVՈ��"&>��?�/B��:��m|�k�ݯ����d ;���Ϟ�ѹ��m�>�� ����V-��p�%��{��4��E�d��5]c�ˮ����� Nd|��[�A����u�sh˜܏]�5؟�oM8������۷�9����w�$fe}���Q���G� ����^@�� Amϛ�*��Ҳ�P��;q~}{�M|�k�ݯ���}�F��m����N}yo�P���%l(�a�dD���:@Y�������㞒�
�i��h����=����>�Ax����s��`���e}�_ ��>7�o\Wt����x� f �Fd{2(�yw�A���������;�.>h��yt���Yԣ�Aw� ����[�ƙ���x�y̀�AmȐ[�6���s�U�y�4�1��]of�^]�4lf��%�v�q��[A;�����9�s�R�Nqol�Ѵ�V��_��t��>�+����o��y�\)_�A� ��mϧ��E������i����FJ�Z�>m���^���b��ۏ�w�@�~����Ps��,p�C�ۙ���"q4p��cxQ�d��G~<>��.��p�}j=�;�)}��p�%��	���>������>�.3c&4Φ)Ĝ�dK]�'n�r��<���t��t+����o�����#,��Ȓ� !��N���>s�Tn���T��|&�1C�r��{�m����-��Ŷ��[w����I���}��~ν�����ۏ�o� A�  C����7��ٙ�a���z;�����|�!����|@mv�],��VI�?�츮�г�Q�ߔ���^-�͵$6��Py���Yp́d�"N8D�
�s�Ϝ�}�q��*s���">_c]�ř�����h�4cFm�m+�� ˮ�ϯb���1��׽�ȡ�O\�xn�S"U1���k]e�B��R5�Ϭg��X,�4��i�V��|m����nڒ��q��b����-�y�T3�ym��7�	�  A�>-��М$��dn+q9���(JA����mf�����n"˒2:M.L������љ���\���]� m����%�X٫��}��gb��"Ҋ����/����D[jA���":oc�zY�o���)��ٟQϠ��{?�^���/��m٤���y���@��^�כ�P-����"��m���aqy�m�ߐ>?d ��,���������������W�l|Gt�Cߦ|ChwL��W���oD�b�|w~S�#�cnɢW�Ɯp���^n��[s��y_ݣ+�G8!V�;�Ϥ���n���>	�� ���p/�������H����FOl��N]Ʒ�p{�,�cʖ'-����L�,������Wڱz�q+{����~�f�O�������q�%<�sUݒ����y[��!��f�����;V�3��BP��J�m�튡CL�ę�̚�W���vv��3}��?�"+O+.���6=�B��J�f��G��^^��⯔�Æ�/\�Ġ+.>[��@����f���]�>��͟�x�cn�(6��jԑ��R]&!^�5��7eg���=<Er��ɨ:��Ie@�L3�=��4M�������z@��ӻ4��iͭ��l�U{+Wt*�eΔ"[VZ�E\����,ȝ��im��3D�B$n���5+���$oj�^w��:�-��m��p����T�q��w>�,����f�r��D1	��7��QhC��߇���,�-sb�9�w|G�t|��0a�BǍ�E7t-^��ׄ9���5�ǡf�]
��tɸƄ��za��kgl�5V��;�9�(+�\��FȾ3Q�l�=�we�V�2XGUlk[r����u�(�������r�k��n����F��iˮ0�vo���Z�'B4��4=��aԇW�4��-]�ʷv������;|` ܸ$>���Q�aJ������Du9�.7��o����@���b&��z�z�lLl֪��n��Mˉq���^������y���r�����=������gI��ze�"罝����׬OR���u��fΉX��g�w{�y�}�%���v��H=�	��H��c��(h��`�)���?��Q�bY���::mfGsn�.cD�JD�:+mIE�o-�,�2��-
,��-��㽺�;�,-�K��
,��md[n�̖���S��k]�l�+8�[e��rۛ'	K-��z5Z+w�n�tm��Ziٜ��p�ɲ�k�'y��[H1ز��[m����{vy6��j�{�Է+,3mF<�yO{��komǶgi�Ym�׵�6�l٥�n+MmZ�d�y`p��k^؞�����{����<ԋ6qy�m�c[Z�[)K�ʬiazÔE[l��[,���e����Cu��Q�ݺm��-�f��;�̍�%���/k���e�q-[mGy�zF�i;(��:mY�N^���-ZZ؜5�6�oo^��ihh��������� 8�L�b��)�r�۬�J9t^�h�@�2��`i��	j�����]��WIÚ����
�bi�%c��u�Xʥ@wk�*4�4t9�l�u���K���e�܊uY���ѥ;{M���
u�m	`Z1�hu֤HlhE�]���Nv^E7]�6]1B�=n�ri�v���N]j��xF�����P�y#�h�aI��b��!\U�cd�����6����e� A��n��hç��ܶKe�Eqd��m�ɣ6΅��]v-�L���;i���9����:2�κ��	���
�M�@�Tl�*�Rm��̶vİ��f�mӆ�u�険:���g ��r�M�6�ӗ,\F���A��9��;�ԭ[nJV����3�l56�^�:�1(mU0i��v-ú�H�u��Cr��`{��(�����2�*�lE�5Xk45��h�)��e�4[a�p��e`�1t!�n�����_��-�wZA���+v.��cQ�]��ϱ�㮙H���Й�TQ�	@�!�a�
U�zXt��'�Cyp��=�nm�P���R��E�@�u�S��L���ѱ�Y�U��Ӫ��W;k{7	Aۚ�]�gL����ŉ��ո�h��8{v'���/I��J���'�i]W[\;q7
>�<"��10mm��V�g�!u���=ql�	tqn瞑����d}m�%Ӻ�ާj�<e���\��Ӗ��
�leu�g[s�M��-��aB (mn�w=�����%���8��t]��!��pځ^CfLgs]m��=<�n����.�{:S�]��Z �*�=��N��<��=�:69�Mgn��R��0&�X�����J4�[k�f�T���Ԛd&)CG`�IR�gm)ce6��͐ F(��,�5�cb�H�Es.��q���:ū�닱�6&L;�d��0fUz��1ghƃ�V�q<��-��5�4-Ky�Ap��<��\�<�]��L��tڪ�k��-s�N�n%��]`�15R��z�T���6M����=��xݧ�ͺ::�a^�b+�u����m�Gs7�:z���:�5s��0�)(s����iH��<���2�e�}\6���f�Q�:.�׉��b�r�u��=��8+gGKv�^��*t��f�Ig��8�	��!�ٺ��2`��I�۠�a��i���}����5�����p��|���`n^xf�Z[�)vAGl��u���q�� ��$�y��|�S�Ϸ1����y�����A�,�N����|>������6�A�n"Qq���\Ԋ��{�����Ϣ6n���h�����ϔ�~�-����7TЁ�b�X���[r'Ÿ^!�3�'�	W�u�c��!�f��.q��"�� CnD���n",�G�|(��k)���|�=���jy��0�b�g��n<VzX����yOϻ�F�o��k"&4!�"A��mCo{M8�_�E��uGq���[�sBϚ�� ϔ�~�-��Ŷ��L-[b�A-%D�	գ�85i8��Ͷڍ�#^.m�ĳ1Ƒ	8k�J�:._�'n;:|�_�!�)���s>��{��?��H��q�*�P�#�A��}>n<� �L�>��N�@�����3<	��y�]Pvkzf�n5Sj�TO!6N>2�-Të*滚1qs-��/]I����nl�ዜ�2v"^Ee�E�>���R5���(غ�3>ۏ�o�@���#~�$�Ew|^���z:�Ax����8D�D6����D.�US[�Ls۫/NX�sw��Y������|�����P�^n�F�on]�
��u����0�Cp�]�׹�I��[��?�C��S.3"xw������%���������� ��������g��n8j� O�x����[��hV�xme��T�&�"���ݘ{j��c���p�0o\n؊�K��ꍑ&e �g��LH �}� ����h!�Mc�ٻ�c_k1�5?U��+���<�V|� �B �������"#w�ȉ�(]_9Y:8� A���*}���O�έ�ݟ�e!�9�� ?�D6�0G���PR�H+�b��5$�@��mE8t�����.��ݝ1{���)���eP6����l��#����?��m��}��<m �9;ئ��B���ڊ�z�Vִ�V���.�3��l�5|��@^ �ߤIn<�
!� H?s�;��v������}�/Kh.飌}7k�f3�q� �w椉��M}���_y���� �i[��-�q;���}��cq��_׹�?C:�f��̤>�� �mϧ���9��g��F#�I�����"Q2I��k^��sƠ�+=.;\�s������s5B�5�������A�"� A�m����L�M�㙏�?��י��N<A��D��^m ۰'�ǩK���C�O�4}Tq��M���F�|�}�A;�)#~�77-��f�~3r���Ÿ�������.AF��m�;��r������fW�A�̄C�6�|[Ax��<��|�ν�K����ؠA��sn�b�b���Y�j�/}�#��٭��s?|�l�핷.u��F6�ƥ�v}K�=��:�:�0�)��EAl�ývu��KE�6	S"gw2b���e�N�؎���S�Y��D��s��Ch"o��������4���;�꟰�8�F�|�|'~� �� �p�%��}���'������,�c!��14O9knt���[���º�,�Ҧ�л;M��7߬���=g��H-Ǔh/Bu�u�_�V!��7g�_H�e��BT�Bh ޠ��>�6���������p��'GǮ�ߔ�����V�Y���Y�F���� "o�'Ÿ{{�;V�W���,���ϐ�{ah Cn@��ϧx9�۩�U_d����[��cc>j> ���$���/|[jHm)�"�O6� �͑ �B� ��U�׷}X���ݞ��M�z7�Ϻ��"Џ�-�X��up�%�����LB��y���JF]Vs[y�1�g��@�����D�
-��7W|�V(�J&�"�	�6:���7�����Qs�v��s�y]�kw<���^'x�ǯ������*y.}�Ƽ�A�7�Iҷq%������SL%��s.��pPct,e�J;$VѮ�@+R�����ϱ��jޥy%Cr���c��b����m��*�\i�v6�ܜ���t��]��vAv.z�ᧁ�&�lZɎ��'1a�|�;�7gI�2�7GJM`���M�������aM�Ղ�iY�fhx�Cn*�+qA�e�cd-���R��8�W׮����u�,
��=���TnM�w<�t�iWFJ��� ���O�=I��}�݉�p��V0�U�n>cc>j>#蟞���}�\N��~ ��΄%����@��E�����w+δi��@���g����א6^f��̯�o!_�"yQɾ����h/��VA��G͵c����	��_<
�ݜy�l���~p�!>-��D6��/� �w}�唀��7��6��_aǑ��Q���״u)�e������� s�v���ۑ �ղn�y4'�Wm�}�]f��������6כ��y���RB8M}d�:z�Re���p��N��p�{mqKE�n댗k�p`-"P2A	(���}��H/��q��R?eS�i�9�����o��N��� ��H���Cng��!��#�Q�wٗ#M*�MKx&��p�1�ӌk���(�����9�{?g��+��&��.W��	>���N��|�}\z���ґG&�x��H��.��}��~cc>j>]���o���>q�D}���|^��\�' �Bǋq��En��������Vm�}�]f���V} ��D�݁>-��-���w�)V��Ս��LF���A ����_s
����������� ϳ\85��_�� �p�c@6�	�p�>mCnN����c�f���>�V�Q�8l��c>��7��pm�y�������DTu1�;[�g��\�dٵ��gk�!r�Ym��q��%I���@�p� n}"Kq��
��]��p�Vk��eg�"��!�j��e@^!�/7nڒ3��}�,k\m��V?�������F�V�
�ݜ��_���G}�In:��p�=V��ߤ{�[Ax���p6�8������e*��AI�P�N�n2u���=��L�ǘ��:�8g�i��+)�ś魫Qj��ƪ�8]9A�:2�yZ���i�ϱ@Z� ����	m�7lo� R���H#w'���<�s}:����3�Y�kᕟ ��^#��۾�����m�}��G?�|q��p�>-����[��Ю�N������?uWs
�ݞxo|>��#��[�&������|�����nA�(��cb�,xyոոs��%�VͪqpGh+�S3🩁 ��<���!�3�h ;��W�l��b��6�rg����D�,��֐E���(���R��-�^#�mƨſ�����j
��}w��gr�^��+>�fB�mҌ���]S���}������{�RA��[�A-���~��U?Z_6"ٱ\��:��k�/|� A�O����D6�D�.q<p9��C���s�>!��쿶��i����|A.�Ix�T}�>˩$��*�Y7�nׄ�w���N%g�6C^�ozu���V��d'��i�9�����m�~��~���x�c"X���O�皤Ay���q#��37R M�Z
:y_?����U���f_�	̄ >@6�|[A������Ϩd���_�EM�-M6�.��K�`mkr��2�W��h��* ���R���_ڤ�� �[�A-�"��|�^��㯇�����f��߾�� �Nd���^m��An=ӵ�1�}_,[����W�>����vs�ߎ7%��b��gb�Aߗ���ߧ��^r<8�r���p�$�A�7�)���=n+y�^�w+[��fg��d !��܁>-��n�����Z�~��m��8@�[jm}��E��\��:�|��@�� �8�=O���S��q�3�n�[��m �ג�=�ߪ�>=��m��}b/ywy%��b���v/Hߐ@��[j������
�����"����z�[�{j%��N�{Xvgf�d뺩Ť�%�f5��	��"�h��^;-3S��2t�z����ĺժ��["&�u�r5
�9��n7*X�ʘaLҮ1h���Y0X&��-�%*�F]�9�J��0jX��3�K���)�������ٌ�L�♫���f�Y��YE�E��\���!��p�6�W�ƶ��Z b�u�v�Ů6�����i���ܷ��\�u���6��WT�\i�c�2�F�&�b�0�EIE�r	f�j`��W��j����=vi� �9�����Oǝ��Z��2�����a���~���N ��n�B������2������A�5Q�x��Tg��G�pw/|h"� A �Ԃ.ϴT|u�τ�>3p� �5"���zs��9�>��@^ �ߤIn!���r�|o�A Go� �����n��6�G�2c�o|�G-��y%��dǾ9ؤ�7�n>m�6��у���n P}W"@?}[Ask�}w��{M�����H>9���d˛C��'��P@�E�����q�ϵF	;��z�_��Ø���j�?d=�H�� Am�GTC�U�}�3�LH�$�%%�Z�KmB=YK*+JWM��ʳ�ٿy��� ��^́z��\^�ǒ[]g�;ogs~�ߢ+撰A�#�^-�$6� � on�����룫�&eM�"����n��u<��p�̎�\&�k'Ά\D^vb���1B������cٗ����*B3fn������`�z����Yv��	��}�]�{-�����A9��!�ۛ��w�{��bP�A;��!�n[k/+���t��zq�<9�4p���'쀁ݿH�[� ��6��3ۿ�R�r��Wξ_F��A�D��1K����Ilg�;|';�D��Ӛ
��B�`�B �ouI��p ��In>+7z}�b6;#���4����2��vKokṋ�q��!����|[C��^_��>d����^
x࿧W��7�;@;h�f�=�[�]X6�۳���7�����O����� �ڐ-~��"��\<9�?���G��nŝ�� ����sam�r$[��T=�f���݉��l���>��px�c9�����;�w���]|>q�ȑQ1@_/VZ����'ŸDАN��2�i���~R����X�|fyl)��n+K^�M��cYb�fY;�[[�$��ٚ�֛`|}R>.F��rp�۵3ma[��59.7�ۭW��TH5�uT�S�,�iu&����G�q��.�ܞ0ܺ�~���\�w��]���G����Cޕ|��.��.P���3�K㠦�rM~S&�{S!�9�I�&�&����M���{֣��k���O�j�E�Pl�}f%�o>�����Ê�1�N����G�bp�_j��󫮾]yͱ���}���S{�w3<�:�����4A�^��2a4b����d�VӪŗ��f�5	�55�g+oǴ.�(sh8"#qK�/vr�qf-�t���C��Fn�=���Of�����z���� j����̔c�뺺o����q���`�ήN�[��������L�˦�kq������ڦv����k
��W�U�n�S�qZ\����H�RqTN�λe������ލa�N엋��y���3���xx�r��w��}�b�X֖2�L��#%'t�K���#*7��h�t��yy9���5����_�����ϣܹ;���ivk��9�ɚ�-yA�-�o&(3��A�cP���O�[FdF���N�b=>ۃ��B�0ɉA�s4���<rvt-V�µ0��w-ζD��)n�Ϥ�;���~���&[��}ꏬI�y����dk�1�L�ԩ�/�M^�{|�7u��)�P6����uyz�V�^��;�.����zߨA$�@&��f��9�k��[[��(̎�NZ�ve��k&%�m{��CO{���Z��[`o{�{e�޳��o"K�緻ѰK۶���m��l۫���=�<�ɝe:H�;N�n�Y����8�p{wi�yj�A,�X�ɖ@�N�ӒYݒۊ�Y�	��oR���ggXF���'#4�m��i�jN6�s-��g��k��V6���E�6��Ӕ���]����M�2#��m�v	/KK-9JN˴�MlYLܕu�͙�e�j��5��g[���F��<�'indttVNlۙ�f�;$����R��̴�,����EgK2�׷5�q$������bJJq<�B2�cv)"!��i��6��+8�q�m$���kx�m��f���%���ܸ�&�$�BY��V=��{_��H'2ϐ@ۑ>n-� �y�S�����;���ԁkz���9��Fcχ�W�^� "
���q�}������� ۹�x���@ۯ��b"�\�P�A������5xq��g�G���ӿ �p���0��"�x��D��D2d���I�'ַn�;8,G[��V8}W�5ڵ���������>-���[���Ͼ��{\73�#���*~{�w}P���D}�D����p�%�����b~���c���yG)����b/O;q���g��	� "o�$����~�S�h3� Gۓ ��G��n|�3�WɒaXV���U������Nv)� �p�%����@����p�ߦ���~q���_c�̿���{\;3� �s!{��U��|{��G�Ov�7{t�t`W�7z����T!��H[TB���*3b�J��7���N����c��OG�Ch�K���o�"� %�����[�߾�tQ� _إ��lE��یŏ�~��x�;��%�D��_����q��S��������R8"U����Bۖ)���Ӟ���0M�h�F;o�o��K������!�3�C��~;�Ь�sᝊ>4����GW_���X#z?8@�[k����p����s)�h�oaGr�2�c��/�&��ó��@��o5����i����A o�^ ��� ���ȶ�֮9[�3}]b-����X���o�~���In�!�>���G^��nw�#�Do}3��}8;�����s�b�|v)!=�sb�J)�0���I��A9���-�^ �ۑ%��������yWڸS�&����_�lM�����y��n�Ŵ+︤,��W�F�� L�����x�=�[�.��ӎ�y']�_us��W}�G��^+]�.��[�)�Z�CA���^d\"�0Ύ�Հ7;n�<e��\�듪������[�U�3:q�wV:��=�t<;Gh沲[�v�x���Z���hn6b���f�%�+��^�0f��2۬�!)��C��9�F��Hk��gv[f����6�{)�TeT�	�v%���ˁb���mr�ֹ��x�wS<�pj�bv|7Rq<��^��D�E�������{�6p!��t��5�r�t��K��K�q�N������K����۪|A��-��W����cY�����!���S�Ԧj ��g�b�A�h"s ��"�_b?G�?N?�e�����㼇,}�P�:�y�Q��'9� ��A�'?J����n��G~� �����r$�mk����:J!K�mũy��{�����Ϥy_ �mϧ�6��@�޲���M1�k�7`/�Ǒm��>���cY����� O�;�_9�H����?C�!����|���Д��X�X7���/�� �0[�_أ��v)��@�@�rrU��h�*z���R�rd0Q$��D�2�:��	�.�R��g�� ��N��$��sG�����p ��D��"m"e��ו�?�M��6��9�.w�U��O%�� � ����� p� ��REw{6R�c������=��In��J;ȏ^��T���9�2�Y��h+�r�*h.S3����u�J��vT�z��Qȍ]�"q�n[%�����B ��R/�����o���F��� C{��q5��I_nnhc�@v|���Aۙ��h}�3��òM��t�fz/�Q�>��> ��W�mI���x>��=� �O}"AΏ&�Q2����ϟх���y�M�"�]L�0�i��՜�CO����7A�������`���>38����0n�_ί���#~~�F��$�M��c���\Oٗ��a�c�e�V�Fg�$��Xrz����g��#>�����bAvw �m����8;�����/�b�O�3��rO΢S#2�^[k�ߐ � *��n�z4�B�������V|��-7���τ�o!|�mēH�nz��[�'^� ��n ��Z�w�~
7|��p���h�Co4;�;OQ�*�OE%.!\�F��I����M<zFj[Ow��G�Z�`3�g�I����*2E���5���wί�����������>-�7 6��>�N/�I��z4��g_�ŴӃ�t7��,����>k��A�ѽQ��/F�p���Ciy�CnD�����8�s-W��yJ
���̬��uc��m�����|�!�3��s9�[���d�҃%J"&BB�[7����<ZK��ca�W�=9�u��`*�]���?/���3W���6ԋ�/��tv���ۑ����^Ϥvyۼ����k� ���mϤ�zۋِo��|��h�s��練}��C���2��_أ�A�jA}x���_-߮.s���ҿ>ā�Ϡ"k�����-�����3km��ϣN��߇^|$�@� �CnD���>�Aӡ���<oT����A���_6Lح�w��܏�o���>N���W���W2p^��ͯ
�/ة�Wu7� �5����UTB�I�(1� `��Xb���@��B�J�i.d�޷A��!�>�Kp�!�����[J������3�����D�Y�_��{�\׾���ȶѫqxY���D!���D&L�!Q�GNJ�X��=�ݫX�h�v��J:Z]��{�c,���w9��"hr�}��?�N������!�Ç��=�q�GFF��������@�[jH99����;��i��	���_6Lح�w�_nG�6�?d;����%�C�၂����}Ё�!� O��#Pǹ�~��o�ו�"C��/E��> �\ԐG� �p�����א�ۿ3�qP4E��/��6�UG����Ͼ:v�m�:�� ��@���1}�]T�I�/n���x������Oٯ���o�%�yG��ܳ��f�}��"�܎�y~���[�Am
��t0�p�܍79F>���EX��'T,A�,`[n�*^1�����j�OJd�:��� p
�;�=X������#�D��pѢWi�����؋��p���muvr�.:����({G5�ci�s���7���p[�2q?�?9�9�s��6w6(�=lp[�ku�)�*����5�x�j7;8u.깬��ř�Ó���C�CE�ogA�J�J�����-���f!�)��^pU�4��5V�*�Vh3-��m�EB-
9e3(�&ѹ�@�x�����s�b�F���l��sj���h�E�.��3��q\v������[��٨"s�����X>��\r$:̲��(�q����}D�K�Ҩ� �@-�$6�����>���5�fp��B ��u5����_�;S7���	��y� ۊ�)�\�=�
�G\"7ڤ�^n(�[jq��1��(��&�O:y�_nG�7���� ��,�h mȑ�ۋ=TEZ��Gr;:@��]U��W�%�S��}�>|ԑKi|�v�D�1���D���א%���[��^��ka��~�/75��Y����χV}>��A|�!��>m
ﵑ���q�J���@���ٓq�ܶ����2h�K������[aa���~�j8|wuI�"� A-�1���n(N��ȯ�#���E��`�a�k� A2D�����bA-� �>���,Zش$���O<��b p�5UՂ�7���n��0���ҋy�Bs�]3Ȑ���C;����^^��ӹ�������Cj�}�����/2�|+�Q�>�k��� [��cr�'m�-RC� 〈-���"����ڔ�"��y��:v�o8v_���|�m؟7�x����<6;��J|A�Z�8�	m����"��K̉�r8F��쀁�Y�-=��ܜ���h8�r���|�/[A۫[�֎/�}��7Z3��q9"^e�G���������[�%��U�ӿE;�]_0R�NI"D!"LD,Gt�.�m���乬1�U�ٗL	����o���@��D��mJv7�7�|t�L�p�9��p�N�>��F>�	�p�p�%���rsl�'���ȼj|�~�qqr{��D���� ��Inw�?l|j�@���xb�>#2�A�ϡ[A�^�����Oږ������Ux�����*��Ia��F��\�NS�<w�P�s[6q�ޛ�>��Fɓ9,��;3J��[��j٢��j�ƥ�]n��O2��_b�� �r�~�y���R���~p�Q�?@�As� ����Ui߅����ӵ3y�ܴ>7p�D�W�ݿa�7tψ��^-�ڟ|��q��߅��;�]R���ȸ�?t�ȟ�#�w�@��@Dw}"Kp�6��7�?��>ڸ0L(&�JSd-���q�Y8ƻq �X0�8S\���$h���O��D}�݉�m+��s��"�e8�Wأۘ�p~���f�0Ed{�x�mI� |[�7{���K��G!��������.����φ��$w���Co숒���}_@r;�O�^3��>9�) ��E�@Am���#�sj����{/2>�������@^ ��In<�
�����w���D��"�3����_G?��sGS����>�>�� ���1�dBص�W��o�S�?�53nw�bn/N��i1k�9.W��;��\ ���+��w[�RCS���N�0�N2�����@��H/��v y�ʹ	n M���nk�
r`��إ�U�ߋ.���_H ��>�k�ݹ�t�������b�Bӛ���-��]痟)	R�<�J�Y���.,-���T���~�ß5����p�>-�>W�kwrys��Ӹ��x ~����ެ�8���H9�"����Kp����MX��s> w �쿹?���CK����>���RA��n>���+�Rmy{� A�"Kp�>m	gs��ﾱ%�Z��n���qS�᳟	����6�	���n60��uf�>���}����ax�m���qG�u��w�����6(���{Σ�;`"s�������8}������@�U}���+(^\�wOUtg��z;S��"<�/�  BI��$�� I?� @���I?� �	'��!$�hO�  BI��O��!$��I$!�!$��  BI�J�!$�  BI����$�� �	'��!$� I?� �	' I?�b��L���e�t� � ���fO� �6�6  (P  �     PP   T P   (

     P�P P   J;� ���( PU
� R� (*P���P(
 � �@%B%�
*�
 ��� ��
��PE��%*�TP@�R)TJPJERU@T�H����R����UTAJR�T�)
�!�   v�UUAAP�����z�b�ۡ  e{;�{��R�x듻P;�@9 1� :�RN ��=��!�  7�O6�	wRR���y ���`PWk ��� \�UP��@ ��{�@
 � t�G&�
� ������ 5 �(��  �UE@��)ER�)RH�G� � Vv�>���d	��y���E�
�K����UA�D�T�7UB��wqԤw\��(�PB�  K��S;u/���)�%.�Ԋ��RU��P1�P���ͪ)\ڕf5R��"�AB�� |P��"�T�ET$�}I.���6@���#��;�T8t�3T*ww)@�7сsۉB������W�� ��{�*� E |zHS�>ϠA;�tRV�*Q�^ث�w�!B���,�(�-��R�J�� ]���`=�筙Ew��%Nl
�m
P�D   ϪTR(��"�UA(��H�n{OT��A <��� G:�T����� =���`;��({gy�:y^�A#ޣ�;�:= �`x�" ��   4w��C�{���	�P8������;��ɥ#ޱ���*XJf�����=���� AJB��  �� �*%U@��R�RI��݇� ����4G��`�s�T��9z(t.`�a���"� n�EW ��F��ݕ�
E�   �G�@%Ӿ�G�����f���� H� ]�.@wgOMPx���!�u�T�4�����!����S�1�SjF�=�R��  4�*M�� h ��JR�@ � 	5Oh�*d�x���_�����l��+F��$�����������9�~��$�	%��� IMHB!!��$�	'�H@�p$�	" }_}I��?�~"��?���`�"�?�u"��a�Kد(����.�XT3^�jлmش+��<�j�R������[b�޺����<e�b��U`wF�UhI�q݌W�hIQ;��+������A]�"�ރ���f`�tu�4-i&t�v�zwC���%���iU���7��An"�ASr���`W�l�)�{ZZMCn�f�É��!f��KP�'�b�M�Q��7lS�m����"ۣ5Me��ŷ�
W��i��PN�O���Sw�hX��à� 70�o�ʼz��h	�mMwY��ugjn�ۗ�lذGU��blʆ�c��Ȩ3�Y��bKt�P�6�פ'��˨ �ɆC��I�kTW��x0Ic7�^š�֜L�[�o�ƶ����ǲ�D�Ŷb�{�D]e6��S�r��cq�[����,U;®�����ֆ�{[�h��^��K��qf���qwf� ��7KC&]�HR4����9E� �z�fR��(nǱ�(��u,쥈�2
�n2�ܩya�%���]*Lb7�䵚�(QY�=�߆�eV��,�Rj^��� �hz�!�,k��{df���Q ��n��i�U�R;Z佑ѣ��q�f�cW�b�P+kr��+�͒��k�ǅ��.���r��a�7n��11c\�� v�fclf�	�c/	a�8u�F�p{&���]�2d�w#Sk�t�yEL�.�F����6&[�u���4���-�J/������v��㗱e�/PǙ�P9B�Y[B��˷r�`��4ҍ�c0��aa
���5,��lԕ/l����"���q�`*�s],�ኖ9�1[�u��ט�Ӎ�*[1���Lϰ��K���gk(�m��v~�r��E�-hŶj�Z9[z�j]ؒ��/X͙2n��;I�0T��M�Nf�ꄱ��;�40��1nm:�Z����@R��{0��h[,km�F�q ��wᖒ�v8�֖r�n�ʂT�e[�-an�ڣcId���.f�J�ْ�/!��su^�k-H�3 f�j�e�P�X��h��n�8n�b���ǒ��L�6f��tl�36(rӒ�,�2�ě9�ތl���+M���[��r����oQ�\ ���OVޙn��2�ނ�Aje�JŨ�`@�.�am�xFJɒ��]���<oD��ݺ�v*�6�N�J�+A7Qm�Y �٫dvhǔ� (Z5�V�-IPTZ���`Hݛ�i�e�>�N��0�}e���B��!��ޜ�����R^,�(Cb�^�*{Oפc�Rh����D��۬�Xw^-��XYA�o]�;o�h�����Jİi�Ee����+Y.�P[���dv�VD�9��hhdf<p��:���pAua�ݳ�q��%n��'�&�t^�*�����/3�qV$ڊ@�{Z�˩oNm�;��FXr�kt\�7[�e��`jzj�J�cV2�
�SS�w�E����Z�%��+F�7��Z?f��d"P˱Z�J�4rCo�h,.�4V�[�dK�3%�ɦƣ�,M!\�v�m����2�JԹ��G���j���n�h,�p����*�$� ٗ�T��>,6�Խ�'u�iZ��z��{��{�w �7����U�
�tG���������1UjG�J��E��OK ��Ǫ��W���l�<���b�tm���;3t�Yyo۠�ԓ)��&�ݫ����4 Z�n�*Y"E�:n^�wqGP�	qP��-b�t�|��v\�if��A[�Ud���rр�Uy{���{i�7��V`$|�� ӹ�bʼ2��ô�YUj���Y�%�=�Sd�-a6�H�$ݳ��MAu��T�Z�X[�Y�DMW��I�>���y��J�0e�m˅U��vU�T���[X�7���|2���Z���%lY��d�d�(`��n�(V+ˣ5ZP#W[�(K36�^n�k:�4�^�N���r�7GT�7���p�3��:��^-�v�FcgkF`��ȵK��-�>�aR��zevK�ȢK��B���0�9y�n�=�x�[�Iϵ�ʚ�T+uԳK�M�-�G2�� c��Z� SX�y�m��V^{�mm
���ۻ��9�Ձ�ui�����֠�����ID�a�����*�مn[T�81�Z����6Da�� �(6�&�b����byxe�h��������s�b�V�`�H�+jHQ�ue�۷a�im��Ƀ,�%�8�r�k])�,(շJ���m���Z���6�;Y���&T�Yd�Ս�ũ�nee��[[��y��;d]�,K�J61O6;�[bd�C ���l�hX�Ǧ��F۽WsE�y12m�i;����^u�V���F�,��V-���0�(ӕx��H�3�R:!�3b��K3 ��8�.����Qј�&�ӑ̓ZfL�j�0��*�Bך��t������c�f=�9&���6���j����%�bu�j��2��?ZT��
����%�QU��Yx���Dbc�2z�.,��L�����^�ܸ0���.���,.�i�įn�]k�P��5Xn��y����d�yon��Uè�+t\N�4���2ХO6�f��wU	V�ڶśe�c�r(��U�NT��J%4^�4[��z+n���x)��kV:y2�Zu�8�˭e����Q�U����c AdK�eh�H;�e=$z��5lB��+pêr)��֮Təb���ɸ#����hkt-϶���m��u �^��z��%+5��I=ѹ6	72�I�u$l�mL(	Ljʊ���.�F��Q2�3(��1P!���l�lVK��l� �,�ZV�5xN+��9��a���7��7Tya!���-���Ƌ�k]ܻ�yA��s{xM�MS�����\�������7f�Y��4�o4���q��[:�y�F���ټtŒ�6��\˧NZje��WF�DZv*˲�|(i^ ��F\j�ƞ���
�:(9�V���g.��27x�	�)[���aǛ&ƳD�������n*"=������{Dv�e�j��II�US�r��+l�d�b�u Ɲ(멹x2:6f+/�P�V�P@�j��ܙ���V%1��2��=!AxE��d�X�`�S$�1��NMGkK֕#ejIJ��Sp��\�fV뙻�Ϊʬ�tS2�h`Z`m��%+�a������wr㻽r�9�N�)0ϘyGZ�5��C��n*�lWO"m��&k\1&F�n��.���1c��x��%����`[�@��wyHb�K{�R6�6PڃU�2�P]c��v�Ux5oT����a�懥�)��շ�,O^:����T7c��o���!�~;G#�k��Śz:u�vڼ.[�0���R;��7��{bSzn�mjh$��EeH�hCv�W-L �gAf�j�Ja�l뙶f}wp˕�Ֆ�Uw(��ܛ���YJȵX7S5�ZQ'MgF��enA�>��}�.?�[3��aK��f�љ��Ӊc���@W*ӷ��7Ĩ�2�#FC�,㈚M�͆j�ك뻴�d4�PA�z�.�	�Љ|��V�tZ�s~x|�[��ͼo[��Ӿ�j��Fޡ��u����V�*�Y�2�`�	�7
�1�x�ɕ�-k٥��aaTU魇%�*�+�{���DF&�U�h�T(������n-8�$�\�����="�Ƿ,���j4ۺwhX�-*
˸iͲ��E�.���%�&�q��82�֔��โ��w̉׹znRԒ�P�uyn\����r�۬T):SX��ҍ<ۡkV��r�	xն�[��@C-�hvb�{�F�و�:�d>��z��q�]\/v��p
�:y]5�י���pZ�������gn���R�3Sh;і7kf��6X`YF�F&���I�n`�D�iL��K%�p��F�׹g*�*FI2<��]�Gs^S;,��v۬��w�%��4��\���:���3��+���֥��5�B�>�V��*-�qO�3LqD�u�@֌m���}���{`�n�+v�'���H*{��&�
��t�te՜�Nc$�6�����J.�Nm�ެ�<��Ҩ���6��Ӑ�B�!Y��]a'Q�ŭ��kem情����pf�ݻ�u��P� ��%Va6�I�YbP�v�{g2P�y[�v��i��RM�զ�Y�N�X�V����Т���Ex��Ri,Nm����V�l�{1R���K�TjrD�g^�쩍�(R��I�He�Zҵ::/(��Z�4�6��"iؤ���êUY^eU�I�6��I�����5a�wy�Zt	��K6�������+]���O�5޸�;��n��m�5���%��1�+��n���m�Mt[�ʈj7%��V�:e�y���i��̚� �x-�V�bT����6�i�4��ܔ��J܊m0���utÂ����&���Ae��{}{f� �����w��ƃ�Ȗ�l[����t�����@���Y�t^��[��3N�p����on�Zʟe�e�����̡�1�w
�p-�xFDU
�K�� PKgeGx]�l^�a�[+6�ju��ƽ�������n�X��fS��J���4�E8˵{���
�隚1�t(zle˂�5`A�v^
y�5����N2]m����7Ss-���m��Л����0"~2�u0:I�{F��!E��f��p�N��Z͗LH��4[sF}����G*�e(`Z��m�q��c�E
ʔq����y����]��Xɳ�V�[h+u.=�5ث�%��sP �d:�b5�;ɍ�8 ����^��
ԬV�	�aV�B60��ĵ�A2�Z�k�հ*#6���U��P�������n63e)�J�z�]�I�%��=�b��W��(�̓2�k�dR;+��]6�ZS��rm�[n��w���Rz��xX�#/.��H���%��]ɺ�a�oTxv��ׅ��K&�5"�S�V�����[{��ww�y>�D4�Y��3l�Z@�Vn�d��2:���x��>=�2Ayy��$�ER�Jo6��Ě���T�sv��t�̆Sq�
�4LĲ�U�M̹�f7jRɺ�d��,7y*%$�dӐz��`�8��{!��`���r\�B	���,[9�3�J�B��T�J��n��[R�Z��ڨX�a�;ks	�Elǔ�ǨXZ��qp�P���q����R��ů3�3Z��U�BʅE&�Ui-�ͭSk2���w4����������V����xZȾ��P.�Z�f��XM�F�Mw��8>�Xh�n�i[CfcҘ1)���kS�Z(�O1���nɏ���ub�\��)��-Xv�<A���Z��ѹw��%u�흶ܼ����D�۸�7(�H�j�w��Հ�BK9[��,S��7]�)ɩL���Vs2�܈�i�p�m�NfS��y�ƨ�tK #	���Q^���Y�n�DMކ3k#��B�jY��A�VcR�V����XV.�+ј�I�U�f�n�
[���X1KN�TWwֲ�Zs�U��qa[*]e;7{gE1tQOZ�fF��e\Y#�n�X�4�щ�� ������ˍP�,Uh����y"�lS�	�6vض+pP� ���^VW�f���*�ós�ݬ^k�U����"���y���>�z�\I��z��Y݋w`:o>�b-9��#[{E}��$v�<�����=bJ4��nJ�̗J�d)�t2��DC�1ޒ�dӮ-[�x/5��^Mx<im] �ͯ_�ۭ��׊��ZF�#J� 00D�6ʵi�)���nK����*Ɂ��j5��*H���miq�N�f��`C(���S�fV�D� �n�
��]Kѵso>:)�uӨ�#dC�-۬(�c1�fQ�n��^j%b��6�h�!��5�ly��H%���]'adk@�2��M��  ̅�pJ��h��,����㒯J�;DX�5�Si�vE���)�ȋO�G\�X�\��t�b��X߮+8�Kf�+Ȅ�jZ�����b���v����ڰ+�tE��-@��ęT2��uؖT�]^҆9�qVY�I�wI�Be�P�Ƅ�Hԧ�A�a���u��\oT�?j�%�s��f�h���J�6SsF`�VQt�%nP�ɨR��eM�!H���d�]��x"��/��V��ll@e5���<"��/r��c%�e�N^�x�٦��8	�#Z$S�a�����mmGt����q�����M��,����=���:��Z�Avf�(L��k^���Ṇ�x�O��)b�R���-��L���:1i���u��(�8t+f�X���/2��]m�P�I���LI�[�g�/%��n���m�˩W7n�A��^�J�']�X�m�׏܌fiX��(�Ȗ�sS���r0Hun՝�S�GeǹܪB��U���Mcb��jk Ii��z�JUn��Ђ��n�z��٘[�Qҵ$h�F3�2�T[�yV��.�o&���ۗV]�%v�u�H�ܹ+4f��1njE����f�4�Y��\ �.]G���
ݢf�P4lb��iG�x�M�M��6��qJSV����q-��]�U��VQ�2�`fE�����ȷ(k'�z����M����Khb�cM�WyN]��&���X�]�&�CtMT�!e:�S��ʱ2�3jZj����:�BK�6!W����Um
����;�+;*}��φ��XF�;���M��Ff����LUx��Ɍf:�C)�P�u�S�"�xfԥ�ݙ39���`d)E $$���I�HE���E�I!()$$I"�H� ,�� � � 
I$X, @X�,��(RB	"�a � )$�d!� ,��a � XBE$P��H�B)��RH@XH)!"�"�"��"��,! �	!"�H, �@��I$Y �"��E�,ER"�E!Aa ,H�RH$�$�B �H
H � ���8�:��*�������$�$�Y$��@� �	�"��� !I��⪸�*�뻸��
H(��(I ���$"�� EAa	`�����	!I_���~�?YT������p�@��b�k^��z�Մ�j�������tN�fb�3������n�=DX@����������gV���4��o�E��(<V�,3+v���_�W1=��ɛ�V��+���լn�΢�e�|�Y>6]�;�1�5+R��1t�!�E�U��ܩ��W��lަ1s�z�lyl�:�p���ĕ�;��7��
��;��[Y.ֺk�k/3��hw��Z��:�v�(�Vɲ�������mv��E����&��.��ϱȳ1��ڹճ1�7Lvڬ��r={��M�%[���\|�<�nФ&c�ݦq�o���pn�^!�|�(��p��}��+�wʞ��z#fQ�b��"�]e'y-��i��u��i���I�!ѱ���߉����SG�SF�+�>b��(����v��L+Vٿ8�	�X�0 ܧ�ۃ���z�׻�z�������2����i��	a�5짠O���<q���W��v��%�d�@}�����0�|�-�Vǀ�l�x2=
�ߧ��bP�3�!�<�q�nn֋}٢}�e�#0\ڴob
�X�p�y�JB�ԘSe��U��YB�{�!��U�B���!�Gct^��T4��㼫�	�m�q]�8@��������yTg�FV�^6wE@�WX�˖g`~��K|쇞O5P�v��H��ݬ������l��-O6���t�殳lfgf� �}R�ӎ�y��o�>T���;�w]��Z�Sk�����C�
4�����-ݵtx�OH0�J��$���\{�R�8�)��yA�aq��HZ�ѰI�}����ڋ^����,;�͡Z/�gGR���[���L��n���)�T�՗��o^O8�Ksl��m�e���eb��&^1��,Ꝉ���U�W��ֳ���^�N�K��j�n^R���4�,�������m��YD��jף�ks��:�VH�y�c�eiT2�&Wv�z���
B��4��2�̇�J�%o�-�);�g�mSbXN�H�P�B��v�bVa���W���!e\�zm�Subj�춯A�6uCo_�+���,�5�4�������Ɍ��}��bw�drB��5"����J�ʹc��X��.�9�AR�b�U���
|���Ĵ��5�QfvQ���+�tݼT����;Mn0�F��7Dk�����򁛈Y�ۨ}��+P��)Y[y��
��6.�xr��6�]e:�W�pO��e���4eI������R6��#�\b�Tn�1V+JƠ��;S��W���nEN����wϹ^q��f�8�cˢN���vΙ�d�m�̭�2躲��v�Z��mJ;Z���>-oY2��-ł�Q��
�sk(lb�7�f�*�D��]�YDM�g6�]+!������&�{B��UZ}����7�SL�h]"{xռ�j�h]�w;σ��c(���p扉X��V0��{�)w��
��hW�L_��SD�`%���#]V��6��bk������D�Vu��ṙ�\����|/9�Y*��$Q��KW�3�F�N'���2T݂YA2�և[�vGK	��w�o�OZT�ʍ(3�j��0ٛ)]![������<0U�N�x�±�/2Y֩�𽌛%�fU�.A����y| ���<�u�cl�rW�ὺ�qt����a�u��q:OBE��"[�=qAH�^�l����Z>����c�{\άxn�;n��I1���6�B@�!�Mso�g���W;�q�l[5u/5ӝ	#U�F�!����� 1�U1cή+�M
�2�:�a[̛���̑���g_U5�WLN�Π�FI�a5s��r�j5����E�v�{���S�
�y�t��y�$ywۭf��B��k�Skr#q-� Z�mx�'�γ�d��}Pݫ�G�ms��k�Gp�l�dP��<����siku��1���.#QSs+X]��k�bq�j�!5��`�R��W��h�b�0ږĔX.��F`/�*��C���8@�Qʹ0ߢ��gM�0n�Օդ,6M�o�ox�qJT�R�{}4Ղ�jԦ-zn��7�dHo�un�pOaiu�w[2���n-F��.�\����v��&�(�Ҩ������,�A����~��5;ܳv�\���v���wGdv��6��]�}pK�z7��>@0:���p5�� �q^ʚ���h���l��f�]�=Xt)Oxt�s��,��X���N8kla�;��P�Nw��O>����9	��v�g+�����5V�2��S�r����`+;J3po\�م�LubU�'a-uҌu#�T]ZM�Ge�ʚ��b���z��_��Q9d�θ�W%���Whm_Q/�S��U���nu+�k�k5�������ܭ��q�i��iA
��f-�-���|��tc*�4I��EWN�W�;U1fp���FE�Y��7�J��36	�����u��![k;f�d�Gk�
u���&1��6蠃Ui�t��7e����![�[vI9;T�2�O�K��a�bo���j�0��l��F�4f����W��w�Z%�#�#��Yw�w���*�,C�����سO �{�/K���cܻĺ��V�ռ�Y���Wc���|�)���Yf��qV=��tY�Mqf]D���0�P H�����هn����f��]����ܭ���� �c�O�D����&�o^L�c�DSˤ����[e�E�pZ�t$v�F%I�uf |vmd:Ȇ����0l���9�]���2�gJ|x�3r�����,-����,CӝY.���Zq^*lr�ѿs�u��w~mZ��:��1�r�Q	�"b*��a�	G랿J�h/R��`���Į�X�;���y���v���{���bq<��kj��pwU�q�݌m�5G�|�]^M$�;�73��Ca%�ŝ��XZ��nfgm<8Kr�����ԭ�0I�&�V��}��7mԗ�NW�d�n��Px�^� [�R�:�)�e����Pp�X5Y�Tq�SozųN��1��ؿDY�
0Q𺨐B�6pOEC0��B"b	�y�KT��C�e��m��x���� ����XRe���^!�׫����w��Y�D�,qQ�m����p�S�*GQPTI)��*C,վhW���N�!�gi��u�Ž�f���;��Z��CY���6���IFR���G&Ϋd�I��ù���y8]����T��n��N�[��Z/)��.�vL��c�<5��*ItFmM�Ɂ��WYy϶����;�� ���' �ۼ�JVE,ӽz��cT�Ե�c����e�*�s/L��tWǎ�5J���$�e�Z��w1]22ŪU/=B�<�JR1YѾYV^�p3r=��^��F^���
�Y�EGp��7/dW�;��"̔(J��ݪ(C�4�(8�w�*x��۵ww�F�J��+.B��D�ӯ/6��þyCy�A�y���B�g%�t(7V{s��0��(�=���f#���o;oz��gX����Eh�Jf�q�s k1�[����7Dn-�o2-�}�p���t�5�y�h�1�R�Gq�;	xN�ʇ��	9T�,���R����#�"�G{�h���k)��n`�	f��.��d�Ƭ�5sDP�m�Lp��N�}����bU�k�%u5����O>�R��z �����r����)33��n�z!y�sd�>z��n�<�L��:��ј3��@֪PY=����̛j��/P�Y\u۶��c��"��D�ni��w���Wd<wC� ��\�U�.���;֨�C2�9�o^���	(���^a�u�V�efP	mU�>l�̔h���2�č�S�+Ş6�ǧ���zE�Ӷ�Ċ铫(�T&0J�U�zCw:��q�����u0�3:#�%gɵ[�b�q��k[f3&ՙ��}��o;z%vŶO� ,܎�N�[f�*Â�,%�a.�ftӁ��]��_|��"&���}w%u�Ån�G(?�;E������Ɠ³��3Gqvr���r�ݗp��M���'f���]�䒮Ηr^U��:����cK[ܵz>��Q6.�����T'L�MM4!6y���n��8�_,�P�,�����9�����S.���{��K�2��]M7��ʗR΅�Wgk��Q]��i\U�e��1�"Na�IU��yr��q��Jʚo8.+�F-Yn�� ���ꨝ:��8�?jjj'vU*�:�\�9EU��Ȩ�2|μ��.��b5�z*.]��Y��Wrju,�[��n\�e�gv]�"��N�#YƓԙ��]�vJ�a�cVM�F�Y ����/P�*�%$�RV�v��K�ٚ1`��a�Ϩq�/6�����B즑`m�����Ŕ��&���Cd�&�Cb�I�}J��xi9}ӯ��|�;�ћ���7�6b�Īe�x�ކ�)�ӱ�=�W�f2�u����J=�}�:��q������!�r��4rf�.�{K�w@N��Ţ�
����a�i�,�aj�\{]i�p^��k7$=ą���fe^G!=����e�ئ5l���=�Ŭ�'f���� x�Q[���wI�*����U%s�x(�零��U�R�u�ޫ��p�ì����A��F�r|x.t_q���O2�W����s�C_�@h�nδCˁ���ݵ�ڣ͗J9��:�!��S��]r�K��z)�=�ՂA/�˫V�ǜ�C.�i�)Mͱ��ƈ%A��"��|)`ܵ�5�dUS9d��t�_E;_L_:�)�eoj�x�B;\dRZR5�m��f�<V��6E�X��;��W^t�̂Ծ�Wo��t2�ȮzI�n�|�yY<��*�b���1/GF<y/�i�,�Y�usn��(cZS�/:� ���
Y]�;���n�KT��r+,-�a���د�L�P[я��%gA��;����]�_�n*��7w1q�xs�S�.�F��������k,.�R��2V�͹������Ǧ�C�(
�J�a�m�y�dD�W)�ޑrx�ս̹pWǻ�;6�<��^��Ts�t[f�P��<�)��.�ۭ���5�ۛ��I�]`��+(���S�jB��l�`��-��3ts��B
��^��#�a����&&a���Nۦ-�H�F��R�5��7�HÀ�*�%׳hV��9\��ͫ��3r�ã�l0Ꜯ�˧d��@+y������Z�݀���(��L��KE�j�U��*n�S�Gp��U��<��ӺF��cMfi��V)�'�<�[�୫��m'��n���x�M�C�xQҝ���R��A���1����]㑜;�tˮ��ɽ��^8�@�v��`�d+k�[f0��O�M�=�J�2:���d�u(�['����)3|�������S_Bm�
��;1[;z�m*:���i���[�}�ٹ,3�TE�d�������lx��hl�u��!-)n� Y��k���&�eL2M�j�
وwJ���:%헥����k�Z+���ã)�ڝ7R1m�+� Y�Y0��N�gj�P��3�KU�Z)����brfav�AyCN�S�z�7t�LY�3m��).�R���7w%fx�Ztf�BX/���Yζu���@>Ӓ�3����-�.A|���u1ְ�c��3�Do���n��I�{j;z���@������[����n ��͆]a�i��{�s�>S���donrVq�W�Ӌ���ᖳ����t]����R���2Y1��b�˪��2g�W�m�������Ƕ�Сug��9.��nA��/�GH@%,b���n��z�{&�E�_�u3T�M3��]�ar̀�b�.��+z�JV�W)�f�J������2"�нť�R���B�����)���#Y~�����\K�-�)�ﲯ�7���˺��ؚ�_Q��a�;]�u�t�"��NbYAӸ3����Ӌ�g1ճc.]f�­_�u!��X��ڬy����j۩v�9s'�i�}y�c�\ܫxm�����.QZn�����n�A��9�T����q.�<�J�]-�msh���2y�*9���i�[���g	��h��)!.�@�[�Yy��W~��x��zN�5P|�hWO[�ckI6����6����F�zh{�4��|��j�d3U�.e�K��i�c8x��|V!�������Q�VҠ:�����p9����]��H���;i��\^<�]�������������9������˅��P�c���\(�Vi���V5#�0=��V�,+R���c���u��頽�ը
D2%7�9Q�mq��D-S7bݚGۏ�8�hN�o�lھz�-�~�M&t�����Ygi�G����o��9����:]W�Ɲ.�k7�-��h��V�g,[w���ԼU���N�E���5�wanV�X�k����Z�u��\;�wc����$��e��'n��ÏRYnIq����4�P
Vq{����FMn�_>#�/�j[r {	�2� ���TKP��B���17��O��u���&��N�q��r\ہ^�d�w �5:ˊ��R���n�1��$�<���1�����ٌ��q�;4t��Yט;���ך]�jVa��2ȬG��n�U����._���a�{D5�U�+jѹ	��J�%����l�q�j��쐮aٖu�=Ym��6���T%���L���b�f�Jٽ���2����3;��������E���L�7bQU\��R,`p��t+�� wOh싸�,�@D���@�dW�L��[>�7`�M�d
n��a�3f�\�a1R���$�,5B[~l�P$�	'� w��5zҴkE��ZЃ��a��/gZVh=�&�1-�ڊ��	�)J���K��2�`̭tق��cV��b�.[�5��̍+5�44d	rg�mDF�h<�SjkB7Vf0�D�Ph����L��5ɰ��[e3q!n06�Yv��]�����"�f4�Tƫk���Ś�Ջ!)-�bf�cs+�XY�lc��e�Rif���N�]�J�PV8�]�)q�2j)¶Qs�����L\,X��J&C�B���I4J�B��Q]#f��iJ�l����a K�e�R"CF���]3K6��i��gG�sY���Qi Бev,�H�۬�`��Wl�n͂��5@r�K&�Ca�J��Y���ju��W�<�0Z��:UNy��5�XYr�]^#�
]�#0�B��MW@ؙ�ҚAF�k��8�Uf�bh��R���U���[2�خ�m��*6�+RZ�s�L�땨F�z��3K���\L�h�&J�f�k�3��91gj�Q���i0��S\S7j`�n"�h#Yt����0j��)�����{B�b�[�8k���&�]���d!-��Qʺ����4�T�f^.�
�m����Qv�:	B1������c��@�ƗG�0u-��S���5Kl��]l%�S�@l���]�B�-�t�[�4���c��8�^����ML �0թ\�]�6�RV�ص�ձ�9�6EMQ�m�]���&�im @vv̮]n���S�mv����E�qX�bhY��e��J��R�ɋP��&�it-0\YE6�t���,[�h3,�����aP��V���f7$���Z%�6[����7cC��ve"��M�iX�;��\,-,7%�z����cĻ�lc�6�`̍[	Yխ3�[����x%��U����::�#������*����̫љ�f�lE"1�4fQ˫�8qea��&�Q���+f��Ô�jֶVKkUZeG���6�28b��v�\���f���^f�2ś0Q+x���g'[E��h<��[��\���0$كKp1�$�tաc��щs�Wj�L�t�Z](l��C�X�C4j�����p4{]������]�ں�Эܑ(���b�2�[���07aMPv��P�A�`m�%.�t�����aq,	60B��k��ub��+Bl�R��23��M�d�a��0(���7�����牥=`h9���lp���]�q�Ӗ��! �i3���j�ږ^2]e������p͐�!��2�X���s]��V�Mr�,j�[��\RR`�/"WiXA��t�tƱ�sA��[��u���LYWp�*	����ژ�Q6k��{fxW���%����Ѥ�fS2U���Q�ed�.��[-�"6\��b4J�;:��֋ �]�[�i���ɂ�if��.�3XLЙ�$v�@q��®sSh�5���v��]-
�Y\Ji�Sf�Ֆ�̳lz!�f�\Ӵ_	{��Rkg�fؠ ��b�f4�ҶJ3LW6i��A�'�����>8�8h@���̎�b�M���%��$��V�7.����q+�X�.&�،��j��B�7ibPq��vִ�ٜ��\�k���l)������M��0!b�k�<$c(�ьte��6�蚃Z���y�ف2��$�e�	�t*���n"�23L	��!us�[V�DV��X�L.���֠�]�uGq٣iT,��7Оq���̭��mt�$p�8���]3�#|���! �\���Ў����'J:�e�1Ybi���7g.ɶ�rfSKf*�%͖�ݓR�z�	�	���9�l�����8!�5��]��AT����Fmme��%,�	k+E4�p֚�	���v�[2��!�"p�S7lT���efƣ2�MSiR�x�Юά�Y����R�:�2�M4�s�4�Jt�M�u�às+�1vaؚ�G\���M�����۝��t�1Bk)�3����`�6�M
��a����v%�K���p�&�&���cJځ���M-��\�sf�RZ��[-%�$�N�j��؍;��@�h,�Q���Y���leeD�s\��c6&#1��*�5�-�r�O^�^�u-5�LW!��ٴ����_<�o#frJa�"e�:SX�mv���+2d�:�3L�e�E����%���4�e����/Z��tK���+^��yS��pˆ��Iq��6���IZ�$,�-�C+1z�qP�9n� V�5�sm�6�+5�-���4Q��+�2��m�����
�
9�	��.�M��m��f¹��cDu�8��P�:]���m6$�uf�`��4�Q���)��L�c@�͵����8tuU&6�J�#�]In�Ҩ��i���6�3�. 9��L :��:�:Ƹ��JQ�k�.��)�k�]�g�Aq���IGY��lE��quVlb��ԉ��Mq�j��/m��F2��=[ 5�tb� KlkT[s�yѴ�+b��fHX�:���u5hn4[nA*L�H�m�B��.�j�]����K4��b���FM��h؜gCٍ���%B&0i�d�,��#\󢋑a�cfȸx(�;�V�`��Mf����J�,4m�m����dF�ʖc��ͻ��M�sS*�]r�[����	.ĩ6�N�-�.f���v�.�ĭ���P����h��RѶݣ5��s
�e�SX�[@�K3m++T���c7��͠�,��cML��9�p�1m�R�D�8P��iU�ٷ�,B��ec��tF�D��h�q��B
f��E�*6Ք���ۻG.���
��hX�Ꮌ.�n
H�KlF�Ԕٮ��(�2CJ�\-��^��Q	����1ڪ�	دf7$��`�F�e��U��ț�L���I[Z�[&%�[4nb��kan��ɭb䰋��7
Z,�lXnj� ʺ���$tj�gIqbMZViP���vt��^Cks,��Ն� u4Y�X��Ţv�
\Rۥ̈́:-Hk��xyQ5��B!�%3��\��6�p�H�c���]Pih�&�gC.0Y�ڈ2˛��U�\�fh�c��-�#1iM7[4���M��¤��Vdk���1�mIh�3@�jhj"J+r�iieܡP-�źXlM(�΢:SD\P��Ud�v�u0R�G�,mu��"A�+K�lA,�`��kl�ۢ�6f��f� F͊�7l�v��Ֆ4k��1ZFG[���bl℺�ٱE!d���@�Q�N��f��6�^)��o/�X�#���2�L�,E�t#��#L�M�0K4.t��m[Mnna���Hr逵���(�Д�l-��4�p��MR;�fca�����+6γDT�@�m,w=l3(��ebh�i��t΂ݨ�b�J��ma�,����jR�P�E-�L��7J�(�;E�b�0�+��ҁ������X��T����Xv�ʃP�N�sh�c���B�bT�f�kE��mH�頕����!v5Rl.�46��)@��X�as�v��)S��&j�!̮��&M�f̻X�*��QZ��LA�sn��
6h郕�����Ѧ��1�%���(&���5T
�i�K)��K����ܒʭ�8�l ��훪R����v����-,L���I��B� ��7M��\̭�^]sqi�ٗXE)�e�1D6����ָn�/ +��x���j��:D�v-k]�tf�#]nQȫ�Y�r�v��[�hY����\)��؄�Mc���(�L۪`�re4���5aJ���$	z��5-la���l,�T���m�w[y��u��[�x�&�ZgJ��0���ֶ�V��cJj�Bhmu��v�Tq��8Q�٢�L�B��X�r��%�[RV����:X�eˈi�t�,���q$��4��S���n��F��3�fh���l:0�]\hY�����&k
Km��ي܈��[`�` �f��3[�E���b!�Vh6�V�j�ـ�٥&&��q�(2���դ���$����.��G4Ҷ��bklwc�Tj�ł\��ڎ��&�`R�i�m�eq�����]D�+��j�F#�%�M@�1�m.͚MJ�q��fyc��Q���f�-�t�a*F^�������[c�iL#�m�sFJ��U�Z�ZăT���p�;jRi�(�:��u�#.�͠�Y��e�jY]�̕Z�d&!b�L˵U텖3`���>�y�B+`���ۥ�H5[6�5��U�Ŷ8jL+�Օ��'3K[mر(%i "cu��x>X6b���-��am�e�Tq0�m���1�`j�.��4!��:hR-sڂU�C�X�fͭ��3Vʊ���D��%0ࡶ�R�S��T�1.Σ�]�yݩ�3t3F�k��4�bm�	*�U�j��5<�e�5�Ԑ�tVf����
�K2eƕ��*c�6������&�0
AȖ�A�.���״��1vkv����Mn`9y�nu�׉�u�)!V���C�-i��S%����$%��;]�k0,Wk�ٞ���¶�	6,�n�Mq�Q�lF�	a.��-�.����RĔbB���\P�6���r3	��C��v�J�]c�&���R��u�)\��M��s��Avژ�+��͒�)�+)��e� f�Gl�<imژx4Mse�eU`䴒��#��f�#ũF�5;0�7�wi\AX]�ݩ��2�h,�^@u�Ǩ@��&�1�m�١�0��^���^��:Fn�B�]�q.K��l��qW*J���
�vT\���	KbZM.,�6� k�Ťu-�u����Tu*	�	\�B���Wk��i��fa��q���SA`�\WB���h�3�����"�
e�D9W[V�7T��V���Y��Y�e�i3 ��0cFX�6ֺ���h˕V��)��V^�zP۷:�H���9�֝h̅�����2mtrM��\"6�����Q�Miˎ�#��8�嚗896�՛۬���Q�:�<�"s����m4�@�On��Z�9g[���s��S��G::[��9ΆYISy�Dq*��D$�P\�ڳ+s���nγ.f�<�&b#1$�J�����Vvڃ�-�P��I�	m��X�]�ۭ�$�viͽ��y�ח�"C���,���َaٍ�z�^���{bHP�����I�;D�Y)�A�l�E�ӑ:.9#���;[J��H���۴�$K��
 ��.����#�!�S�$�gy{�p���������q�ir�ydD^�^d�p{YmZ�[Z8I��ӄTQH X�ҧ�M�e�T�C��mn��q�e.`:��ۚŌ�u��1v�d&�h��ZY���+q����)Gk6��&�U�jF�Ͱ� b-̲��lTěh+,Mi�<��*����h�5�v5��8j�]�W7A�І�U�h�	B�R.�����j�`V������Ằ(B65�ͦ#n,�J���ڔ��11�c�#[c��;F�L�(mq�^��l��a�fl�W-��hKfi5�u���bk�����qq�M�j�`#����Z�5u�}��+@��YJL�1*����&kŊ2��\�!1"P�nX���X˕`��f� ݛ�Z%�u�B!p����v,���´V+fx���,h��#
k��gSk��]�e2�2���U5)v��k6Ԯ��R�T���5�����;T��͋�&�� )6��l���c����ݫ�4խ1��VcR2����R�c�[&��aH4���Q,�`�Jlc:�ؖ�l�3K�����0��A����i���&{,�"�+�eoS#��2C�#k4���s��3BE^ԕ�̔�̵��j����
h��BF�"�Y���d(U�J��$���+�-�v㝡�vd��	��)Yt�!�j��b�D�m�˔+eM���\����auS[*�F5XLe��U�%#��Ě޷u��qK�jCj:��F`GD�K���j洆�bs3U�s�6�Qv�uc�[t3���SYLe]L�Gj��U,��n�혘�����j⣭�X6��B�m���I��I�SU����Zk��FKY��VPحR���]n5\m�3cz�u	eY�\5"��WT���iRĉ	��.��m�՛�3>xxhV�Wg\��@�V��B��nlq������E6v���4�s멂5q�3&��I��v!��B�R6i��8��W�\R��^ ��9-����Jے�s�c��$������-j�B��+�Z��eRհjR�FV^����9m)R"�`�b�%�JӯŬ)`�5�u%��[��maH��T��(�^�R���T�Iey����2��H1#[N� @�-am2^�-��0�b4�`ȤiiQ�s�lY���~���m��r�UҬL9��J7K��&��VLW`�VhUb�$}�����
	�ࡧ� �@I.�֫xnn���kB���!�q�R�0�  ����H��han�!ի`z�9{�v��G4���.[����8a���VGJY��de8�V�|��B �݋ �HΙv��j�~[�<��ԙ������%2m}�6�-����5_��.�z�������3����D��7-�.y���B#�.�C̕Tu�.W� ̯�dx�݋��D2�6�����R{���r�_�9�عn���^p��7����E�P ݿs%p�V�Kfx٪��}��-�ì�`��-�Q�Ζ�ЬF-�1̤��n���/ä A��b�t�:d,��_w`Ž�u3�և{��n�{S���~�d Dn��~mYeKmX"��P��vh[PԳ�;��6�9W��*����6��O�ۜzʌ�!��J�"��N���R�V�*�����q)���HV�0C�������=�\ܷ���+܀p���=��7J�2��'u���R�b�1�̲<Cn��B��iT7�d�S����0������|�>�mX!��yyh����b#H"�,X2R �[��[寻�f^�B�?M�`�u/�� Ɵe����"�����!�Dm}m���W����~�kE��N����ܷ���+�8��@v���_��|�<�rΕ^1"
j���T�WXՖ�l��L�qiB݊[�H̓
�L����ԁ҂6�_Ŵ�����5U�ַ�.>�U����H��v��N5b��?6Ր�@��`l�_<m�wG['ו���Ae����F�����l�`�}�� �A��#YS���ߢA�Ƭ�A�|�mz�.7ȿ��
Cظ�מs�^icL�&��������k��k���q%�� eCai�)U߯��l���d���c1?`�g�彆O1^�@���]�b�t���۱`�n��z���fU
�_i͠���_���_nM���5U����\&���F��Z3EsA��E�VCh A�@�۱`�S��W�6�����Y�s�٧׽���gX'�_ �o�[C�{E�ʛB�"��ݐ��A-c��m���6��J���#N3e5��e�~�;�A��|A��h��h�{�V=�Lb��ARK�����UchYn� �[�x,t� �=�~��������Cs;\{S�5V�8E��׼��: �n�{�*z�&�{<<]�FrC�kv,�H�>-��=��v�5x�s��>���~�����Aۿ�����#��������I�3(/�ޤ?ڽ����q�MX��F�B�����[6b�Oe׉��ɉg�<�/]F���L9���+���z�h�I�Y+���ޖc���·�-�{S���9�d��HQU��U��2���3,�ʴA̢�1�����zf}ʂ���cT����\A}��D7H�mq��D����CK��\*���W���U�[�F���9�mZfl�Z�!m�+nfv��߬�����{���-�[���o�f�-�#P��8X�����ׁ�A�]�[A�|���Ց^���]�,����֯h��h�{�V=�Lb�� @#e��e��%����ݞo���Fw/��	n�!�_Ŵ3۱f`Ě�c��=��'5{:��y�~�#��i�V�̽D̹r�ߝ�n�bK�.��{�B��VP�7C�t�;��sr�r����`�J@���R�:��.K��� A-�`�A�r��X�O��W�f��8��n=�Mb��F�FwX��/� ��I1a������J��	ej�+-A3�%�{�]g+�哬�g�(��䰳��F��W��V�'w5�@��a�=��*�5�����KV�i�˫�Rѣ)����Z���cAa���[(ķm.��i�n(e5��Qts���uv��Ya�d�D��Ih��\tڣ�Kl��e�cJdkh�m-v�"V9Z6XJJV�`fͬ0s��YG�����c(-��i��2���qv,�Y�30��n	����W�4MX�kf�\��\��f���ɢhϞ�~�� B�+p�k��3ZnR[�-�%�����f6���U���K����ǹV3;E����L�7rc��{Ѥ�my�.W E-������G:�H�j����}*B��|c���0�H�d�����;og�G0	����K�A.PD6�e�����}\�#�_#���A�ʹhlT�{E<gf���ǰɬW�F��3�ł�/�%���F�=R'��P�Y�t�=�/�An�k�h���w6��.W|A�����J[�*��es#%/�?mY�7A|A��7JmOc9�ú%֓&�üjX��{|���ޕKw�����A2P���n��uXr!8�[���VSv�[�遚k�hī��EY�f�!UwB�+!0� ���?8�7HN��h���8��nc�&�^����xo�`��9�O�V"�Qbs3A�s*�Sț/�3����zho��u���8Ga�<;�����u�x%vh7m�S[7c�=6�$�R�C$ݻ���W�����7#�t8����;�[����7�Zw6��.W|A�����7W�5b�W��>#ڐ$9Aͻn�_����{��Y�r�痍���ݗ�����)|A�("w7A�|�2X�n�x�{*/�Pdl��-�z+wf��^krl2k��L!�-f+��;۶�|���������M�U��bXCl�a�w�iۇ�Tߗ��ם��Ѿ�Ӟӎ0��W�( YeKm*9�m�y�w�ZIUE��E�V��#S$#�[e�m��u�Q�e����1%�����-�~��Ib�n�!�B�,�;����B��z�~�$5���uq�S!|D�`_ŵ�,���[V��MA�/+�f���@9�X�[����&�&�YC��D9ذ[��y��6Pˬ!#v������t&b�P��o�x��"��~�AIxb���0Q��=�]���4��ܻ�2ޜ˵&fG������[�L�=:zm8��z��8��ڿ=�I�Nnpه� ���:P@�����m��8^���H�6L���!;9N�޼�[��=�`�J@���7�E��/����"�+�	m����;�3N��x�X�Q�����la�ao:a�A����H���8�{Չ����Ŗ�\�UR"F���[R���e� �u��s���T��tM]��N�@�*����������n�s�7�6a��������Րf �(KmX!��,��-:�X,�R���CG$�����Y��d�`��_C��VY�VvJg������$VA���|A ���}ܪ�;{�T��^d�y���氷� �@/�;[������X������T{pPںd_P_ӯ�7A�z��ö��pܯ��ފȽ�s����0;��CG���EPi���bp�t��S�08�Zw_a�<�;:\��jR�-��D���31�N�+PX+	�"͏|7S����տ[� ��+��[�5�0�P�� S�4mP��.I�Ͻy��C�c�`��H$��m���m����4m����:�b� 5����P�U�)�.��b�Ce���j讀B��u��Xs��t� ��Z�v�Ҽ���sX[�~��u)��A�9_7A�ۻ�H-ƫ�Ūg�ł:u��(�u�g�m����� �}�A�-����%���vǁ���7P@�("h_��H���{��/�c�Y�Y�������/�2 �!����E��M��\�y���LA:��փ��D�^j9���'�\�^̏Ļxq̤�o>�An� ���y2��e����6�[6ooY�~r�rW|A7�Y��Am�{�k��=eX���J�.�ݛ���\>���k>�bck7�*�8��V�5s����:˖d�]L���4�<MK�Ԧ��(�]���(e���	' ���@��,���b����`�m�%����u��̡����kf]�X.���5U�mtйk+nтZ�b��2t"���h:�4n���K�jQ���<��d��z¢G�S`Ik���(ps,ƹ��3mt���Wv��6GZi��ZJg6�. T�8ָ�EnEA���֌��o`ٔK4g�����n.ŋF�fCn�W����H1.��U��l�j���S�F[�� �%�-����_-��s�Y�Y�����(o��ۯW��<F�X����n���������\�X8�  �X�[��N����0�.PD�Ŗ����<�Uv}�cA/2ł:@�����?6�'o�u�_14�n���%�����\~��� ��t� �Ր��S�|�+�(vm�����+FN��+ɕ�T���vR?b^Y}�SU�w`�"�X�u�-��_XmtFof��z}�},m��Y�zhny�� L���Ŗ�|Ct6���o�#������k�4U�Fɲ�@�ma\a�R�][c��k�mt�FJƽ��>F|������[A}<�^���9��/�Ҹ�w�}��[���}H��VCi�n�w����/�wΪz���d���SV�)l��Q;����W.Y�����Q�۰??@]tﯕ��I;�)�������|ͳ!�VK�#���P޺�������w�+d��C��@�#A��UJ���f���A|�_ �+��H@-���mhV+������Vl���a>@�(Gb�n��_ۻ�k�ۭ�_GA�F8���S�u��G9�%�p�W~7ܾ۞��G��<�K��{������Cm-��)���Yw�μ�ݰ~x�^g�9ϲ�������� �����m
�|Vue^�}��M��a��%4kYl�͊nu�L�AU��e�u�Zu�,��+��W�F;�/I��㎾E����c��d���l'�B�yE��]�ΰCh�}`�� ~����n��#����{�g�yVs�K���� ��_X�-�̓��ng?��}�Cu!�7X-��
�~.�e���z89v�G��m#UL�{{���4"%n�|暑��7ٵz�"p���Q�B;����ͽ�pJ�Y\��[��,r���ң����]W�6�#��1�K�͌ڙ2�bf�}�1m�bx=�\�'�xl�yݎY�.f����GI�h�"�2.a��c�4`�vo���|�0��{t�+���Чư�Í�@9d��l��
.�7�<%ɺ8,�6�����n�+�ia̮6��f:˛avћ�WS��#Q7��a����+���V���zM�mT�#-M�4�@�%�1�q�&^�3�\�5+����P���H�`[��.7V2e�D���1ڭϦ�9����(^Wh����qf���%
]z�X�s�UB1��`���^�9q�×�:���ي�&����/;~�B���{Rr�b����۔1�Z�h��f���g ���
T���w\�Aw��ŊP�A�wK#�&P�*7��zEnC%Z�w\��0Bd��U=��Up?n�ߛ��i�����tҋb���˕j��+c��TE�/O��}�ɘ�2N��ֆH����&�2:���p��unk�oTլb�ux\4f�5��P�����Y���Ԭ7�8/^��*����ok�ܸ��ޯ!��#�!O/��Ic[�MK6AZ�@�"�(�yn���y��.ׯ`f�W��c���!%�uBc4��Xiu�2�z�y�98��z��gpu�a㵛�=�����j$��YL���Jg��Fv�]���<�|?l|����}�]>o��:��d�,)��'p@rvd(NR�h��"p;�'!�Y�� S���f����P��å 8�8�C�rr�q�Qmj���mD�Ķ� ��-N��N9D� p�B K�I	BIee,��n\� �-��D�Rr\�N6육�C��.)��)(��kC�,�DQ�"(�\�89y׽ݤ3K�H9HG��%�r�1���	J'7$� :)9,�$(q	�ۜ !DH�	�	'	JJR'H�"�8�p���v����Bps�J	D�3)��;0����H�Rq"T�D���:\�rI8� >
 &�� �=G��y�1;�P�}l�1�x/��"�/�T��c4�4l��#�A|[�A��F��1;�vI���| �AQ�-��f�����|}���6����H�������L��@��&��t��{ǱVs�K���� ��V�h"�"-���w�_�����o8�b�L�!*�� e��I��ֆ�n3
�v�
�6���� A͠�G�,�͡[��s�3/wp�/��������h/���_�6�-�[jȥ�z�ԿS�R �mh�-��n�7Kr�O�&Jѡ`�[1�,捽%+�"=�����mCn���\���}�C��ڟc�q�
3ܬ��n����Ct.��c�Ew�6�}�,�A6�[�]:s�������� ����$�g�*��H*T��F��א�o��8K�n⡸���ȇ�l�Znžڼ�%P����c����ܨ}O��a�ټ/��|�x~-�d��Y����F�R���y��[����M�Y�C\(v�_�C􆻥��6`��|7,�Mf�U�ܶW8J���2uFZ�[$	@Dѭ.�%n)����㲑�۱���\~�\�>�7���n��^� �o��СR/�W���Vm An� ����y���9Ծ �A�+��}���cx�㲐D6�V�Lm�	��o �>�@�[�`�[�A-��/��C���F���&�n1[�d�>�e���_۰,<��{w���lU������S���}��בap�W�o�Y�՞�]�J��[c�_K�W��	n� ��Yn�RW}�fgum�{�G�	cu�gwff�Ā^>��;+�"�݋����wx�g�]���dwcU��<B�vk��aۡ�z�B
s�X{2Xb����n{�ym5�æ=���J�S����J?�|=�m$�ҽ���6��e�&f�ٷj�-5��V��iT�^��Vۃ�rb����m���K44�2�v��E�L�]^�ib�4�g6��a����:%%+��ۦ�YQ��s���dX�5��ɖlu��0.�\9ܚ��y�&��5�<'��K�B��%��R8������,�fS�\�P@�3����.��?��~������� љP�ó3uEJi@�+�t��R�``A�uz��U]��fs���s2�3���s�����l-��pKh*�WN�5H_P�G��_�JD��źG�'[�������ޥ3 �����x�~��}y�q�r�<�@�Q27Ȋ�kE�f�X#�|�:�"nł�"h��I�Ʈt���};3ۚcy�/픈"D!�b�-��� BYY�}��yY�3�|?�Ѿ���n97Kr�[��(/����1��ʱ��:i�U�=�X&fh��2�L��iT�)Kݵ|~wM��섯S���ˇҸA��y���	m�!陇��]��s������H�M��_�]�b�l^n^�Z5�vk�50!M�(̤�����Yoߤd���Ŗ�m�:��wvf�i�����b�^�O��ZJ�A�j�}_�6�-���[j�W���Pj<�S���7u�0�ǒ��&�,jÕj��҄�Whvog\טZ4�ܩ�"sڻc��e����>9j�u�P�cn��� &��d� ��^�n����st�-����� �v,�G�K����F�.���� ��6��_]��e��z���\�y���,.J���V<�_� A��Ր�CRD�������b��H��/�[���;�۹�c�{�`������ML��� [�/���u�	m���_7X�"�<#K9~Uڿ�y�Ǟ7�)�l,�&Jz;��� m��<�S��脵�UZ�BWT��d�UAH&Rl�ί]%4*�p
���+��f7=�ϟ�K~�e� ����͡q�Z�k���ȼ\>��{���Τ��W�W�� �A��?6ՂK�� Fz��������}҅g���y�j8`����4�6�/K��_]Pό�@�\k�mt��������z�듐�i�3xA�^���)㠖M��q
)��m�� �ڽG���2��#~�;U�o������AH�X�43yT1*����}�̘�C��q�������b'��5ʱ̲�fe��Vn�̥��!��n��xvi^�uL���������E`>����K�60�R �_5`��"�A]��^�8�Y��!�%���;����/sTp�/7��vRDh Cn���.��>}�|����}�l������[�Y�mқ�F���A\����viHWVP�dW<��ƾ�E�G�ڽ��Cs��79-�{�3��-�d�X�u� �A Cn����Dɗy���ۯ���D|	���� ���H)����+��}�5������S����2RAB�Ro�!�II�ݨZAI�)��ղg7�o{=E���P:���e���I��Pi�AHUT�� ���;����ý�ZAH(q�J�>�3�C*M�8j���~�K�ݸ��������'��a�T-BRA`W�zH,4�S�큹� ��;چ�
i��[5) ��~�����sz���}��4�R�}p�AI�)��U�i��P(JI" Y���gW�1�C��Џ�?t�
B���ZAt�����|��m~<����J��\�,켤{H��������p�����݊�;)�_+���Fg>���8z���6�ͼ��;�gG�Κ߿�$�*��~H,��L;�CI) �Q�}ZH) �{�I����B�5����A`hi �{���ӿ��?�������!�jH)�~�s������_~�m��0?z� �>II���4��RAaA�nH)4�0;ڶM2�
AN����oy��������:G �MH�h:�f�����ŢJܖ�*򪴕Giat]k�Aa�Pxt�R��H) ��������Ja��-$���0�kI��������럹�fu��)7�,>�m �7�߽w�߿d��B�
A`~3פ���I;��6n�)�{P���)��ճL��P����큤6������_���/���6�Ri
`o�[&�I>��@?�6�z�~�2?C�����T- �>*�{�i��
Q�{@m �q��w�Cgy񶬺��KH(X�^�$�) ��e���Ad���ިZ���{zH,4�S�큽� ��{P�|	�}R��
���l�ށ�̕�� Q�?z����R
o�!�%$�nH)��դ���);��`li ��h4� �4W�������w�>�ZAH)?w��:�L>�B�В�
;��Aa��?s﷿�������zt�
AM����Ad���>�Z�RA`kO����]{\s���i �z�ٺ ��3�$���j��d���S�큤6��
;ۆ�
M!L�����;�ߵ{ֽ٤���)7��4�����5�ߏ��ٛ����H,5�H)�Tz� ��R��t�62S��hhII
�;��A`��1|xi�+��80��=us���U`��|���GBu����2"��֊�r0�Ӈ��v]G�j��;��+
��?�欄�?~���J�ef�)�2B�8SUVl�mm�B[���g�f���v%���\h�Yu���X�K*`�H�Qh�Nl�9��1cnt���43�*����m4v��̭Ä�q��Ɨ1Y��2�L��k�6�#��3,��!u4���-��TX�h-���F�W�ك6�ک6�
�T��"�%ћ$Mf�]�uAb�cs��]bۣ2;�J攰џ>~��[mLܒ�5������s���D�ƲÆ��u,�V�@����gKf�����JL3ꅠj%$�� �44�S�큤��]���,��"�~��C�~o�J����Τ~�2RAC���{��G~�5|���?j��RAa^�ᤂ�HS=V�R
AN���H,;�:H)
���դC�
Wl�y�7x{F��x$t)�~�ZRAB�g�I��������}�s���zt�
AM�,>�m ��B�5��v��R
AN���z�}���� �C�T4�R>�g�d���S������Xl�nH)4�0;ڶM���Q);��`o�}�k��ýTW�og��������#�O���� �*��V�R
AM{�i���ý�ZRA`w�i���S���6�Y>��s���}�W���su@�JH,
��� �44�S�}`l�R@�{P�AMg��^w�o�9��v�9߀��U��JH)7�!���s2���6�RpB��VɦRAH)�큦�I�{A�� �*U@�j���I(�{�6�Y�Ja��-]�ٟ?g�N�,f�I��g��o}������O���9a���
Aa�T-BRA`Q�ޒM$�{`otAH-D;چ�
}����3f�G�����$�ca��k/��� ѹ�j��G@��%DɈ�l�����A��c��n;�;�:(RJL��Ci) ��j�Rj!L���L���S�큦��fs���������3��Reä��N���=�o*�_W��`~����`RAO��I���ý�ZRAB����Xi�$�{a��JS��hJH,�ϸ��~k�<�x�`t;
�۪!��T����GYrD�yI������{��{��:8�����تJs��!�6����c�����������AH)7���肐Z�#�H���:�����X\� ��ԏ�2RAB�Ro�XH)����I&��{V��w��C{�VN����,0?$�B�
CET�ZAH)4w��H,��L;څ����X�ZA`�sEr�j��~����������O���9a���%2�g�����X�ZA`j4�S�큳tAH-!��4�SH��j١��
�ܿ]~ไ���XC���i �;ڶO̢>�(�"H�~�{ظo��6��go���$�P=괂�R
w�|V������䂐Xw�B��$���0�I���S�큤�ɱ�ý�Z�RA`w�i ��{`?����d�=�t��^k�$�}��<��g��o�����|2RAB����!�%$>��I&��{Vɡ��P(JN������~u�Ϸ��J��_�meɒ��+2����[�dyW;#(����MU��i��H,5ꅤ�eT�� ��
H)�v��Af�)�{P�5RAB�w����Z������}�;��/����)7�X|��%��W��g�s�H)���H,$���ٺ ���CI4 S��f�) �Q%'{�HlII�[��ek\��>��
ND)�ߪ�42�
%'~���៳3�W���w���2��ReΒ
B���ZAt0) �}�h�n2S��h{���x~���]&�
0��I ��2Èm �S)�ިZ�RA`W{zH,F�
w��4�R����C���h�ǚ��̩��5���
Ѭ��x:��zn�7q\ӯ|r�=�z��\�Qz��L���ۙf��bqh��Z�ٶ�YՙIV�[�9Q\���@��Z�y�9������s�Lޫg�
��}���7RAa_vᤂ�B��j�4�H(%'{�Lƒ��i!��_2�a�����;�H/c�
V�{@m �`�L;�B��JH(Pý�$5����}�}��r��} �����Ad���=P�	I���?v�{�W}�3����
s�`otAH-!��i ��)��ճC%$*$��{`i�) ���ᤂ�X	)��������˜N�� �E�b Y�<�{՜7��p����~��������V�R
AO��I ��j�RRAB�w���´�����V����淎�[ZmD���`V�ڨ3\MnY�4��V\]b�A��"۷?�- �߻a�H,�2�{*�R]�� �4$�{`i �p�%|,��!��s����'�,��
?��l�d���o7��u�o��{[�4�Ĕ�XQ�\4�Ri
`{�l�I �{�L��Xw�H)U@�j�
AH)�w�}�����}z�� ���H)�gkI��g+�w~�^�������AH)�r��Ad�e0�T- ��v��XH)���o|�������� ��~�����Xʴ��P�$���`iĔ�XQ��4�RhB��[&�I���{`i��f{F��ݤ�vk���&�zf3?B>�/h�� �*�}V�]0) �{�i�d��B�В�
ý�$RAN���'�{�k\�=��f�w�B�<%$�^�M$�}`nn�)�;چ�
hͿs;��w���Nw�)���i ��$��~�4��RAa��Ǐ�՗�~��%��0Rj@��$1�T�Em;�pVnAn�S]vV/���֪t�G3F��ܥ�A�(8�B�XjE���yf�����n�Y[�H@ �!����)��ʶM���II�z��cI�{A��AHUT�� ��S�큤��Xw�B��?�w����'���괂��׽^���﷬�/��/�R
o����JL3�H)��v��Xi �{�stAH-w�$����l���8Uf���}�녈�F9�c����ʃ��d�K�;U�]��.n�-�j�W����ܫg�) ��ܰ4��RAa]��I&��{VɦRA@���{`i���٘s߼o��������?d|	�m����z��@��H.
H)Y�h�ld��B��II
�;��AH);��H,�e0�j��) �>���k��~�����r�����4�S~���� ��ݨi ��o���_����y����~��Vϙ) �BJM��I ����$���j�+����}�� �{���H,=�:H)
����i��
w��4�Y�Ja��-$����i�'�_�g~����u��K؟���T���
AM�m �S)�z�h��v��Xi �{�{�
AhC��i ��
`w�l�d���g����W~���%%�XCbJH,(�높
M!L�VɦRAH$I��?7�;8o��/L�gB>�/�H)���ZAt����������xk���_@�Af�JaϪ����P��ݭ$��S��"H,��a��-II�]�� �4�AN��E����[� ��A�$z�mƳv%1�8G�3��|2RAB�JM��Hn$���p�AI�)��ղhe$
���UX>������K���{�,vu�j�5���/b�9FPM���^)�7W\�s�\�ucj.��zZ\u������;2����X�����r^�[&Jh��3�u۸:d3sn��v��K�m2*fN�wk�8V�U�i��&�ŕ�̱���)����JL�m�X�7��C*�z�F�l��]u��uy���w�Q�.�MV����b]�xfѮj����ٜw0#��.#]qr�Rp��`m�\GM���%(h���ď�g�	�]��0(�FT�n�DW�T~�M�U�g�{g)t�P���}دv�T���,�C��k3�Ṟ͆b��߃{��
�f�@�� =����	E�:'�t:�Qa�/~��5� |q⠰���f��Y���ŝ�2�8���^�yLuw�~]�yX��2�e�ݏ��bǍ;[c�k.�����U|ݥѻOF���������G��^�=B�{���^��Ͷ
~��]o�����.ŷ[�oح[��H[��Y�y�4�ulʽEHf��#��fn%�����H�x�A��E�aFRnnot���K�C�+����.���I%�Mk�my]#x)�|�fM^SyW��=p�^�yUj]I0�R���Y���*���E�X���Ψ@κ���g5c+2,�O2��/1��ٗcd��� T:��(^Zz��Y�_����ׅ��ޘ�q��v�Wh�e��2D�a ��[�w� ^,���4�ӈ�9R��V�s���{%�t����bK>Xx�%�鱶�DS�'$tۭA��o��<�H�R��6�\蜈Bs�r��q#��Y	1B�r��m��$�@D�@��.! 	N���N{Z@��9ЊNq%��l��S�ΈN�@���"��!�$;l�න(�' ��'pu"D(:	t�����V�s�8��z8DBr�$;�X8���䈎N8�Iå���g����93�*8D98�H8�y�f8I'�"W��!r$
8��jT9>b4��ݮC���^dfV�7hڴ�m�'.D�'C�$��%�7�A&i!gϼ��)�{�z���-�\볰V�p��X�i���4��k5�Ff��UM���6R�(��r��K@�I�m�gf݋X*�71���v˚�ґ�kc6H�f0pE��z�K�c�4��͵#�#eNiS0�vB4eŐX��\us�ˠ:��6�#�\�%k�ͪ?ꯌ��ln֒ щ�K(Z�;R��1Fmae�&��B�E��44L��
���� ��gЗD�pj\+1W2�#��#��$���#���XP�XZXElV鲔�c6�G6�f�Y,��s������k�ܔ`��T
��T�X쵣K��ԕk���ĺ�6�����c#�b�e�R��j������Ԍ�s���%	[HG5i#j�`i1u�	�n�YV��Dκ���qsr��]pmnh�˝a���h.#�7]�[/2��X�Gd����њ�p,]���<B&v����5E�qt Mf�3��Υ	���4�ʹ�*���o��%��,9cE�7;��*��-e]Cn�(�-6QPvv�i��o6Ɣ��;�pL��PԬ]��r$���Z^�ڑ#F2��s�-MԚ]�A�tGQ�M�]��斵�X�d^�Yr֒gs��t�=�Rm�0	���1&@��鱡�#b�M�nz�h2�c�l..�B�H=��Ę�es0��
�a+T�ˉeWJ��fX��ץ�W��H��VJR�i�Gv�K-���mL��J�
��,Z[b+l�G��L�n��Y�9���Ydd�m4��s���C&���E�ۥq]�`�+�$u��&v�F��X[\���٥(�sE£p�{5
�v�8��Il �Nc��]|��6�3��X�ٙ��Wi��cas�iLɶFk3�uֲ:˴��`Tn�z�ɀ���(5YjA�؆�-�@�*Y�# \����gI�`Z�)	����m��2�#����C���B�Vi������^�Ke�A��.L����̬�z0����;`n�l<�1*���t����<ņ���c�STkQ��]�&T�[6)�egb͈*%t^+��`��bg&��ɒ���iiaM���q,�r�Z�e��gX�˘Jl�I�MnЂ�l9Ȅk�
��uqdt�5���Z�4V\3bm疲�C6�W.��Z:;[�L��Mm(��ƣ�Fd�H9Y��a33 nRf@������.ִ�3�����6�^G �MN��LC����éyf&v
W<�t��iF����Aa���������ZAH)5��@m �c%0�j��RAB����XkY���ﯿ|�9|�y��������Ad�_ou�ew���t��l>�B�>JH,
?~�$�H)ϻ`i �hw�$ЁL���d���D���l$����s��W���~�~H)6!L�Vɡ��P))3�03y�=�q�������ǾĂ�\�ZAH|U@���$�ް4�Y���w�C^��zϷ�p��
�}�i ��
g�a�6�R}P�A) �(�oI��4�S�큳tAH,;څ�����.���dy흉O<����V�R
$��~�4�Ĕ�X}څ���S��d�) �P���l06�Aa��i�AH_����u�;��� ���~�@m �l�ÿT-$���0�kI����W}���r����)?s�m �P�a��Z�RA`{:?{��/*���}���R
{2��tAH-!��4�SB0;ڶj2RAH)����a��B�N���wN������|>�W���ϴ>�7~y3�c3��>I��w��4!3*[�$���������?�S|���.�E���M m��S�)b�%!Uv��胳Jm��G��>a�P��	�� ������� ���}?f���~y�����y��s�j�X��!�j��P���f\He� �e@
�k�2�\\꟎4u]�A`�E���w�e3�{ֱ�"`��_W8��P�>�V�X��&6�鸩>۶�͕��aca��K�X�o��1B=�>��>Wy��?�Oz�ZA��� �7�?g���s�������. s*�=�[	��������uި�?PX�O{,&�C2�a3(� �32����7�u��ڞt�ꓧ���-������03� /��P����Ђ3(���� ��Wu����P�asv��{ް4��e@9o9�}�sy��|������(��L!�q�3��u�ס����A�g=p2���2�X0�33P�����������:��@��d����Y��IG��n�?��� ��%� ���3, �fT$7�������K]��%4�l5���!�Ɩ9�P��Zch[�#���;6/[(�f� ��%}A�DϬ&�A>˄-�̠?� 6�������w?v��~fp ,�?��^gzԡ玪�=>�_ ~�p��'��\B� ���i2�,a�{��L�4����	���Q�>ʀ\9���{�����~�?~s�@?z��D{�L!�j�2���}_���uWw���BD*�p �Ac#ި��~��@3(�{J�)kX�	����)Z5��֫ ڥ���(^h�v���/�"�Yk��������~�f�Y��4�ln=�n�S{2��� �p�N���d���,?�"v�-�ݸ��U:}�ӻ[���'ed���n��<m�Pn��ڙO����2�޷w�k��r�O�K���d��
��/e�U��f�G���Ҍ�.���{O�%�ʏ}�q���>}�K�1�6�5�3+(1潊V
ª�SAe�(X�7J�B�YU��5n�ۤ^q������˸�oҵ��j�����=�������E]\�
����y�:-���Y*�p�������yg��=-]��(�#���􆤗U%LE3�Ԏ���joE�ᑥ�]��i��RK��s�+�wm�����_Hh�=���ng.�1?UM+�(N��4�以�*���H�^�s�#��V�f�o-f'k6��o�e�,��o/Q�.�]���[�.�2��@ix�������|�}}�cwV�}��+�bɺ��bWo�[�?s��l�9�l�ͭ���#t|��v/���|���$�n��͠*�b��l��sY�5Yu�*�k���y�۟<���zw��#��홞����o�:u����'��ϩCU�~�\��5~��?�������h�>��=^ng.�1?M5�jI��+M��S�ƭ�޺�Ԇ�9���9�ۢ.�wun��u�[ڕ���^�"���$�P�[y���iOn�B�c��L��ɍF{�{�ya��S�|�U<?n��~�$�S��]o�������w�<۹"7��u}��}�{a{��]��_���C�.�J��e�=�π�ut^��Ƴ����z�^yB�^o�>���5a�7|��yL��t�X���I:t�}��k<�H�I�rdfm@Ƙf�&�������:��M���j0����[B���#��w#.ѻDK.�G��b%LZ�Yԗ����fɹֹj�]*�j�TK0��a]+	�X�Y���C\ы����\kYFnGa���A2&�k��$���\����7C�[t��˂������Վq�"h@��Hd�n(��&M��ϓ���B�7@�e���iI�f�f��d��s�7��v���vrK���������z��ߢ�2Z�hc�a��2�R��������)�U!�]H~�w�@=���y�T�����O%�"���{���I��]�(ms�n�4�?I.C��+G�i��JO=3��s3��c~����L��C!����J J�w|2�ǰT���Ϗ�/�y��Wu��4z�_�H~��$�6�b1b�̦�Q��O%�2G.d��}�[�������N�{��ѺMn5���K/;U��I/:���5ܹ��ـiL�W��+�9����<���y���gvu/i�O�}[7.�C!�\��I/8;U�p�x�0X�j������>e83�t��vzђL���Ʋj�V_o�n��vO�N&�Xojʌ/3�$Q,����~n��wy��V���q~|k�d~7�W�6�o�QX��CU$���e.A�{o�y/LY�.�}���^��5RK���rz���m�خCR
�L��ޒ�j��fo}u���f	nx/{��W�N�I*CR^�[�vI�,�ޗ3;հ��8�>5^�r��b�ܿ�F��E-qnΦXZ��sL@٬L�u�X�˵#�Eq�X,s0���uO�}�H����w��zb��r����b�_t=c&��8�$��5R��'��{�a��j�xy�ow��rT��]�{nc�����|�HjC��W�-WO3�{��ǞY�]�Nl�{fN�݀�u:��R4�H��\Sina�ݳ.����H)H��UK�E�,�>�T��߮����}���}Q��=�L���zz(8����T��I"��Fw��~浏yzUG�/��������±�ϟz�}x�Z��zs�䲰��!��$�2������r�|g��p_q���4��i�]I9v��e��$T�e��4Ɣ��)��.�j��k���Ø�ƺ@�[VP$ّ���kv��wW�x�$ݻ����pq��X֘��p�k��EU!�_���C���T�y���~4zS{��c�ϟ{s�U�d�蛹I&�k���~�d�)	��J�%y"Qǵ��/�����TM͍�T�emx<�������q�"���&����7tJ��d�����c�wk<��M��,DG�k������;ɗB�^U��Yu�����,VT�b�ݦG��m�P�~4yƖj��{�÷��:�VuZ���8�Jk��u!�I�k�)�����S���V,ws�}�i�C��d�{�=]�g��YX;Y]5Z��љ�-hEnhvl�lE]�V�\6M�p�}�RSn�5Rc9���.� ����<���5�W�/�ᒪ��u!���uKS�K8������k�SfI�w=�a��"��_g=ޣ�2M�)W2�xԒE_H~����(�+7z��}=�b�qw>�箫�~���Cw����v��ŷ݊u}�T��3�W�����?g�_�O�����Sh�$������[�t��4\��-c���5I]s�>/�r�;�67��<�s�r�1��²7}g��y�{�7ӆ�U���_?�Zj����;kj�B%ڿ[1���$d��*z�%XDO����O~�i��r�l6%ی�ݚֽ�i�H(�u������*Y(7JL� tպ5B��6�J�jp��t!�K�M6RU��Xu�L�x���*Q��̈́�EpU@�&ݬ1a����l��a۠�҃1�T�����Q�i���1-�ɫH�]o`�W[�#�����V�e��.R�fV�U��v��h��3k�[�0i5�]T�U#.�Ŏ���O�T�M�v�qm��u����E�RYm���\m+2JJ��)
���f<��}[��ݪz3��?V,ws�T��^���wӌ��\����ٽ�kv�xIT���<�� ��?g�_	7w�n���C.���)��y�S{u!�T���Tŝ�<�'N̏�o��5I]s���O�Hj�C$����S�ŵ�-�T����=�Ŏ_����+�J�����>�5}���k��R�� z*V�8$�o���Z��� ���΄��n��w����Oa�9���]�*�]Zm��-ղ���r*X�-d>����Qi��nq��G�;{�ؗ���vOVWY�m�^������H�C�,8�����{���!T�Vs���	��SQuK37�̰�{�`�"�C�1�̱=�o�����|Z��t ���'Qr_�����������?V���?o��^ͿI��	������3��뺘\R����K��Rw�\G�V߾˱���s�¦I�ry�y��P��ݡ�H+�Y��9z�������t�ȼ���+�-����C16[��%ԒeI]�M��+��;]ӹ�.�-I��w�}~�!�&y������������gM�L�0��V�j^�l��e�&��0f�]�k�������|������爛�\~���"�[�U�j�S�v�\�nP�n��n���7-w*�����s����L܋ύ%��'�q���Lˮ@T�捈�y�9Cv����};O~��^^U�(D��z�ya�x�#�VP5�ɨؑXT��2�=��j���|�`�{�+�/v��{��S�=��@��N���I
j������k��U���.J���5
�cwi�҉̩�����t�Z���:�"��C0_�6��r��A��;w%�w��wu�+��K��Ū�z��7-�T��]��g�X�T-`��mL�=���2�>N��Y#�Y�v��R��c�n�Q���~��K@��t�ECEn:r�ui;��L�K����I�Iy���]G>�C�<Gb��8ʔ�e�[eӇ	��R�qi����jv�xV��]�Wˮ��8��,��X�s�onBl�i�%�I�Pp
�r���JD:Wes�`�ۓ�K���{J���׽Z�ߘ�c�/Y�QZ����[lZ�O@��3�1y^xiU{ ycF1��[��n�ҖC�<W�x��;={Ι\7P����(Һ 2⳥VJ6�V�{��$f9wB�������QQx��o��,��}Y�X'\�H!8ֈВ_�)@% J��w�Q��]����8���M��0��Z��7��tM9S[�X��{SC�Խ���2H���.�Y�ieކP��Yqk_J��Y�m�dF㙕<��1KiJT�K���~5"��� �
^�z�j)��T�h�K#6��{<+o|�1 ){&}�%�Z�I�j�y���a���h��[5�D{2��^]+&�Yu��ڳ�wK1+�z2�%��Ç̈15�Ɖ �LN����%i���%' D�N�f��$�t��s�VRJR\�S�	p���I�NP�!Ӽ��^vy���󴼴yn GD��A	9ΐ#�BNP�۬������n(���I%<ĉJNw�qw��s,�l�9��|Y�q�D�t)#���o��|jN�/����5���N�.D(�k��q�n�����2JI�6�6Ф��G|v��̤�r|�x�Hۭ��ϛ�$[V�$C�P�G��u��{���W��I^�=���z�Y�ghrwe�{��v��{�뺇��Ϛ�j\]ӿUﮫ�d?I$U��K=���n��U�w���,T\�5��j�7�Վ]>�$�U!�<2i��W�K���=wU���g\K�)'��p���Zݯ�h;�բѭ`�v)XT�K��\j���N������L�#(��!Pաv�X�޾5[I.�?9Ow��z�..�ެy~���+J�<jx���E����*Z�9-Ȼ;�4o�7�?wczy�t>����_&�ؐ��~ݡ2�����C7p��eD^y��z��{��1�=K�?m�j�5$����.\Zk���!�<�=�Oc��L]ӽ�箙�c���2E����Hlk|r���Vx5�ޏ��	�C-���Rk[�X��e�#���է+��2�h{���[a��� }��T���{�ݭ�n����2��ZW���Y$��ꘑr��<�߉ﾽ���b�a���b|q��1��t�\%�ĭYH�+R�M�.�����}��m	��_n�O�ٵ���c2��@n�xN޽\��>�H���pX��\�����ʫ�����>�nߜ���_��x��+������|�Ԓ�CR2�����l��^}w����;�Z��������2bW���^Ws�v:�q�T���n�g�R�#I��=_.?z��9i_>�MWq�]H~�C������������[��ݫ;O�۷�6w��t7hn�S�y�i�7�yV�����w��>*�:>���&M��M�Si��/����"0��"0{F���$%�/"E�hM���I��Vꙺ�zhձ�C69	�39�M�]h&�V��/�
���!o.Tim�j�a4��%��B�ڒl��i�ƙ�bd���cJ)cf���r�Pƍ��jh�\���1����6-1�� �a@˕J�0��RV�����#iY1p�p,�L���v�i4,�Q!l�a0e�6�mB�g	�Fj+�+��#I+%��ԙ�����]��MY��U�E��2���XXn8D�`�	].H; ����k���@nХu�{�r�^�����gTf��>��~�Ԇ�5��⽃rO����t�7�)��t�c3��q���J�ԛۼ��;�J�5RIIV�ӡ�#��}�&-�ޭ�_�Ԇ���W���ީ�r��UR»���<=JRr����Q/*�;�ƭ
y}��I/�I��[���Ȕ���<�^���I��=T����R�����
��>���l,t��e�Kr�V��vƕΆ5�8\)��X���C��)�z�n���x�Ž;Ԯ��y�OZ��UJ�I��ߟÌ�󬈿oC^���,����;6u������t��e�<�`��C�Q�wt��Re��d�"%�x̾�"��tդ�+~��> }�ֳ�e	+껯w��w�u�Ҕ�m�|������O��~�m^_�8�ws�t;a ^g���������Jh힪\i�nC�H~�^��Oxh�9̩��/v��B�{Cs�*��^8�"�os���o�u�~�}!��\�gי�������,���+�;�\�}!��H�P/)�|{Vr��ca�T�]�(ݚ-�؋triX�-q��+��U��K�� �9%���P�۵���l{2$��r����n����k��U!�]T��K|>��J�z�N��y��o��r���͖����	s�������Ȓ�~�]Hd�~�@�t���5r0��.��n���:f����@���# y�����
�e��_��6����h��5��~Xm_�|>���޿p��zA�}�BJ��ݠ6�VH�,��.�ʩ$񝯦����l1�}����7F-|��{3�=��Hd�U!�C���^�"���K*>��d^�$�&��R�_��2��6wЪ�+�ņ�iR�J�Ί^")���,!���%X=�qQJ��HU��}�BF��ڥ~�����w����j���=je��P���d�UR
as�\ٵ�s�9���ύ=�c�=+���Pmcuϡ�k>����_�����ʸ¸���݇���)y7�{�z��k��D���e3�9��C�nХ~����p�|]�^��[��������Q�	l��3�{ʃ�W�4V��N�N����][|��@1 ,��d��:�w�n��:�̫�uv׈��ߨ=ԏ�������_w�$��Ԓ��w�].��o�'����'l�6ｑ�f�Ҁ�kwv�K�5g�����7�͵
3.�Xu��L�K�Il�kk�U-�͈v3٭L�������ӽ�ק��㓏^���گ\���=�׉x���t�w*Iu!��5�&z��Yq�>��}�&�nw��z�V��R����d��ǽ3�����I2�H/J���������X}������q��?Hd�����)�b�-[}8���V�j���,��.dY�ם��"��Q�����\�C�%�!���"^Λ�uu�[����UFj��I.��Y��kRE�ע��t]r3(ͭ���0���3/�?�`���虌���-Ȳ)���h��X�ږƋy��Fb�Z6�{���ϟ�wI�/��zF��c��e���zɶ�����tf4��B ;d%[	fE�T�lX&����YK��İ�*vݠ�nu�$Ulխ3S�B��1��.�i]3)WD�u�tE���VY�R7k�.�@%2�)���b2�r�i���c�0X�B�4Y���,ҋhZ�a���T�Y`��v0\v��ط"6bf�,�V).Y���E�cn�43bnf�f�����E��B�]��1ٌf�QVRj�e69̱���k��+��5X6Pǿ����ކCRK�e���>��N5;k���iE���j��k~���Hd�Re��#��Q��}/��ڵq���[����2w���{MT�Q�$G��Ҵ	����jI7�n���U[y�U�ۛ/��ȇ��[��5RI$��|-]��&�ܝ3�%��ٳK��615�ޔ%�]��g��jIT����yZ�W�ފ]�,�Ǩy^c�:�y�^�Z�N�\�v����V��/D���7䐺�²J���D�!�Ņ7Q��*���m��`->���N�=��骐Ѽ[��Ş�Z�_�� �/D�������v���~��D�۞g��-$9��a�c՗���T�)o� �Kٯ�t�I���{}��o����*����5�&㋳r��^�v�W�W�U���E��d������q��]7Ը����� Ԅe�o�#�l�U!�]H2-���q��n���au{�k�;������۱r���߇%6)��{��Ş��[&�̹�2�R���^���w�롩�K����pC���y�w����ݮ���&�g���1�'����M�;X9v6g�f��tF�gH���ݳ��"U�8Z�6l��h�7u}�V����G3{�k����{����ꦟ�I"���Y��as�ެ��#�����t�u��*�/_�Z���]�OZ��}��	u�Y�i�����9u�oU�fZq\��i6S�Aڈ�����Ԓ��D�7r�rc����W_\cH8ooF3by�:ɻ�e��8�$�R��  7sٟ�0��};4F�:�g5�_n���T��.����\u�ݡj��p�Z9�=5�d�uםt>4+�b/��wH��I.��eի�vhɔ+�����X�:�e��P��"���ǉ+܇eP^fY6s//0��jmK��Ħ�4��̣r��k���)0`�$����jz�hnꚷf�aR��u�Do�{�X�8���}���ݡ���������rJ�����е};���2w�g]W�L�(��LM}!���!�����\[�g���ʂ��smo �w}R�.�	�dn҇a��_�-�亲U�h������Wǳ�W�K�]�p@�uQ�&j"��ӓ e�-�kd�՘�vm4k Z�m�DT�k鸯��GH����<YrA�U)��}�C_O�ER�C$����@��+?f����!׷�3y��Y��2��-f�[u=����G1`g2�Mh�)����)		u�$�ih2��U���(��z�(H�}�n����K4��C��\�O՜wX�9:���]H~ݯ�u*�'{��9���&��r�+��һwԴ�mԙ���eP���O�I"��#���W������õ�o>�κ�����K�m��?<��L���}���V^/{=�z�����}��N񫥮k�)&�}�d?I/���?�*�^9{�����+��u�+f��:=r��s��������\�#B�)3%���)C�,{nT��P�6�_7&�T����1n�#r�E)���)(�Z��I�m�lc��X0�^��6,5�2"��OQsF��K|���bܙ�Wy/N�ᥑH	%�7*��֡*��I�o���|e���D<����\j���"���ɹeYsU�������D��5w^-@hq���w5�N��W���!vd����7����?{�N��R�^��V���ϷK�{,�n��;�F���~�^��]Ԟ��mE�[�cm�rM	�{n��K��_^�*:���p�Nc�"כ��R�P�KSd����b�z�rL��KT��e��s��3O;8'�Pۼ@��+'n+���ޢ	њ�z��
��l9N���eK�����Oo��\X�(�Wu;2�@��ݎ��K�O�[�:��wۃSĻ{�ł�]<]%��ڱw2�%Z�������:1H��#	s���Ŗ�ʓ��ܱmЎi�/�[�'��,�z'[T\����6��:��#:�l�YX�[r%��r�VZtX���~�kc�Q"5�"�*H<�N�V��RxǸ�z�k�%u�V"����P���X2�O��lc�;f��b�|��w�d��>��#�����RP�os)�ѕ��s7���C2��s�J��M���xtR9�����NC��F�+�;���V镣I���C��B�	���dуu�����v��T��wsCk*��=!?k�yKa�m�L��t���bx��o�9[�y��
�

#C�"}�}}��$��=6s�gd�t�d 6�!:C3��t�{n�ε���$����Ok�'���9��^ZD�G�[��m�/-2�{�{�-.�&݇���֞�^�+4�"<μ׶3y��w�m�m�q���b����V$9Vc�=�G���Σ�����ŗ���^��$oz�8����0wy����ݎ�/;;;8�[�и
e��$I�؝Yd)���"�չ\y��,]w���e��;m�����l۽���e�g��ڎ�mJ@�����]��`�$e�6�w�c<LY�V��uR�u9c���ZR\�0)4��e&D�M̖���Fb�SmrZ�]3�Z�jm,�dD�le�΂R���̹,�I�f�A���70�'^4Ђ��r�`���6d �f�ˈ�`J�̺�-Y���!Gsq*<��˪[kF�#f��ױ�Z�̔�"��F�k�R�bl�a`M�[��R��kZ��p�,K��0��ƗVҰ�9XB�t�tK�%h��n�B:"M�`뭭sLR:a�u��D���LSB�U(�]rB�Vjr��F7�b˚�G(���hiv��V`��wi@Sc
��]���n��K44�u��eҌ��E�atu���%b.p�4nE�^�lձ#l֨p+�VQ��s42i���i\�˄�F9t-�ؔn�HB�!��%�m��;�.�f�f	,ƪ�]kF���f�L(Wf8LA�����eзj͒�fDV��F�Ɨc7[\��`�cb��P��j�@�]�
K5��LK�¡��ac��Z���vN�6�8�=�,�4���Y�ɗBYu#�F`,(��%o�y��M㔆�l3kdH���JYH�:��3M����nf�����7BL��)u\醰�`��чd� �f-ҵ�b�;�2xJG�+Gn����c�Y��M�˚�(���7Se]��ʺ�A"ˡc3l0A̕F�Ç�-KV�XʵU�-�.4(�Fk�2ܕfz����4��l!�mK�FS��T�nt���i SG\@��5!R�Ԍ3e����ٖ�@J���]�2kb��ae���ݔ�5�f�Q�Yt�������ݠJ�Z+��-��vi2HZ6�Vj�X��&643	i ����V�v%��۴Dⷖ��C��4#�k�";!z̉Y������Yqs�lZ���.�]l��P�����䄸[ts@�1��Ƥ����n6��0&�Ԗ�vn��N"�%��I�#ƃ[Uv�:N�$B���]�l�mn�f6C�������qbQ�� �
�ºY	�R F�W:�u�Zj�U�v��ф`�:k�bW���e��dד��5mM��!2GS�/���u�h ��XӶ�VX�DKf��gUXʖ���8�آ9�YL��\��sqT��YiiHC��5vgLi��Bb�@h��![mqV���X�Ѥў�~?��f�i]	�8y��`˥�iN��$�m,-�1f+`UZ��1�m�_�
��N�XO;h�7�>�F�<�0���+۟k�{Ƥ�!�������}�;���'/
|=]�9���~��$���״��x-�u!�I=c�d����<�g��>��[4F���Y���ww�ԡspE�5�~~��۪��ӆX1�Eֹ������&3��/{���=���Iu#�}���W<��#�\�s�Z�ަ{Nss=Z�s��@n�ٵ�m%T�\����Y�h�*CWf�]A��k���	�ҌX��4�Z�m>�kC��k��Oכ�����Ȝ��V{�9�	M�k��?Hj9r���}�(���^���g٣��I�����ew|��Wk|Clv;�籔�	Hll�TSę����m�6�����������~�����2��m��}���n�~&pSM�oU��/�ƽ��%�!�� ]������t�=�}z3���f��Iu!�ي���曋��{cwg�f����7*9�7��B,�������|d��Hd2@�C�~5}���z����c��i�~O������=�=���>|���]��a��E�mhd�ն˶� K��*�J
@u
6W\T�O?t��'�~��O}5���x��=�}z3��18�s�~>���A�[���%�q�;ʯ|'���}����mH��qI4F�f���w��&�հ+�:7�����IuR/u7,��J�s��SN
���Y)�DF�V�_�&<rċ,�Rw�1�}�ޚ$�l
��c�¤v!@wҴb�7�K��ܦ�2�zL��~��ꑭ~���ݽ翩�_���Ir�ߚt�m��y��y��ݡk<�=�N736�<���NZO��`��״ԆIH~�H=�}�í��K����>p)�$���>����w����?b<�=�8�.�	 ���É������J�dD�`��64(�ԎA��i�?='�k�����{�`����Zs*���^�[�\k�u��7kv��AEfצ�V$��V�ܙ���3s3o�yC��!�k&x�)�&�MUI���T��C�E3����p���}�+�z�5NzE$�������1�J�G�Hi]���<9�*z����B����K=��8ք���}��)vz���]��0�$�U7�28��c��
��xs��#|��׾���z��������sַkv�u���H�Ρ��]QOrð��L����<�ηu�ö儶��>����>�ff�@�]��	b2�`)��`.�U	��8�rWK�D0�[/����|���=����>��h�{:7s!5��r��۵��n�{l\�ϲE��j��wߕ=Nc�����l����~SWޔ>n��ջ_n�7��Y'/!�&�=�E�w=U�״�$��\F�Bm��\5RK�Y�xޫ��6Wl��N7��Ɇ^�wy|���?I.�CR&ڻ>������_ls����^Om�}��@s��?T���t�ʳ�|Vsy{���8�9��=`��fm+�L���7r�g`<;6��I����2�U�=���hF����%�ma��UWȏ�x߭�k
�F�]�V%u��Z�7]����	���x�j$*I�앪��arAs�,&PËP.�d�9e��ʆ��I�1U��[d�5%�]5�aXG��A�7����%Ig�a��5���t�j�c]G:jT�1ե�GZV �Uu%��x���=c�K�P�\9�.3����W[�+�mx�2��JD�bhϿ'����b�Wd��Ȥ�&z��ˣI`B�D�ƺVQŗA+�Uf�4U���|����v�ވ>ズ̅�3������2� �T|����R=c���s�u�v�����O�=/^������k�}էso�������E_I�]���K3S^�M�`k�^�~��XЎ��}��n��2dɫ��]�����ּ�}X+���������������i>צ�C����N�8s�VoP`)�v�ބ����z�M��ֆ����n��k��B�Z)C����q֠�
M)�j�]Z�G�[q�ڨk���Ϥ����U!V��w��<ƫط��x\ܱ(W�˪��I$5!�gu_sj�p�3��z���[�V<��K�^�d+`�GfN6��,�[�L�f�2����EQe+ln=�c��D�꺘���������Gu��U`��W���g�i�#{㫥G��{�8�|��i�����C_I8����cF�V�� ��%��s�O�o���$���z���g��K|�D�/����(�>C��zPF�ڹI˩�%ԗV2����������6�>��ze���P绾�n�Hn{��`����"����U}EX�hе���bЭڴ�B����Kspi�M���+|����g��{�*Iz���/{�]q��=뮧J��c�W��|������ݧ[���\U�$@=���9'V�{��;�1�Q��J�f7�*o>���9}]�ER�-@�f��־�c�h�fI�������lL�W�ߒ�`��:֓~�%��$�������,3k\������D>���\�=���s��<Պ�z:������w���'v�n�(�R�k!6���C���A�_[���Й�u�C�m F�|/�;��F�|���ݠ� ���n��ݡWu���g���rt娞�~wz�>nW���ݯ�_G�?x�b�zo�AV��Q�5`a˱�N^����9��gAז�)Zm�è���)]qS-���=��Bu�R�5>��g	��}�3��0ׇ�g��RPz���t��P��uca����Hj�Hk��ng#YQvo֏P���}i�p��k�E�@�:@��\�'9��V��֨���?�wTv3�V�n���Av���_�L��rs�j&x�'z�u�u�~�������C�I�M�e0#�_��|wP@%�9A��|߯�u�a�P�&�s[�G:<�T��u<��k*q��gS�����'Л�.�i�`����qC��V�|	׬����vSvH�cw�g1[������s���RY��_�~�!�C�)/�譟�m���*���x�����Й�u��sk�u��оݡ���<߼<��%_�X �k�l�"��5KXF�n�c�g0;qS:��tJ�*��ެ����C��ݠ��������h�������T �����&�]	������Hn�T�0x�v�����}�uZ�<��`+�Ǎu�a����B���{���Ys��@��/k�A�A wi��3��v�gsFZ��[Bg��"ߪ�������!�CT�K~3��{�_gݨ/����ݯ/G�n�ܱ��@�nW��{�ju��f�fT�~�#�HDn�	ݤF�!7fd�f���.A|�:�׻:�
��t� ��t+�j�HlP��Q�:Ԗ�o�e��0�G[(e�n�d�b�&\�O`��N� �S�CE@By4�T�w{�GJVY����n=�x���C�n�3A#C<W@���V5�z�"X]�l�d��b���lm^Ѐu�n��˵�r�˜�)k��vl�.�hrWi����e�P�X�#K�[.E�
�A˓rL���u�sG�Hҭ6�7\�D"�ɪM�l�w8��i�F������)a��nK\�(E[�M4uB�Ĵ�����+,lt �����gI�y��=ϳ���Ҧ�uh9�ʰ�-�\a�s*��:YQ�b3	�\Ҙ�cf�m�<���|�ݠ���	��hL���[��iSpܲ=~��Y�F�WC��u
�ءBCb�M���*�x��9K�A������״M�~[m��E�GDݠ�ꌾ*�m7T� N�|�ݠ��K㺇�u:�{�G��^�VZ��Ďj�O�c̩~�'9V��pNr������w���+�n� �@�R �������Be�E��_0�)T6�;���RWW��V*Cb��ة]
���N�=����}2N�U���ۖ1����q��!��@HhR�6O�pv�5̫�tK+��Ͱ��%�2XR�%�,�^��%���At	�z3��;+�vPDn��ݠ��t���Y��ĎJ�>1]Oy���#U�j�0T�uR��T�I�%u#ax�Ρry�5*�+�@��8d�.e˫�I8<7	����ʯq�3W������!�����ߨ+W߫\'?-�&-u�� Nm|�ޠ�n�(OKR��"�3) A:�|A�uݤA���F���S�&��n�\�m�c' '�/�=Gv� ��A��CF�F��ٶpP�.5S��!��ןt��Ag��9*�����ޣ��uQ�$7T*CU!�(}%Չ�T�`[�I���CԼ�`�9mC1k�E�m/���#u/�����P^fy�_�R8����l�؃4B�4�k�[�9W��i�1>'�e������6{��z�һ�y�gY�:��rǧ/��	�s�g��B� �Gz�?n�_�� �_F�'<��C~"����"��oh^^]�7�=\A;)GD�hμg{T��y�T�����,���F<�P��� 5�2(��cv�yʺ�{�ޣf��CR\u;o�{Q��F��ݕ-%c�t�Y6������բ��1�ۢ*�����d�-���k�K4��:�(g
#C���\!��@X���샱�(=�q����Q�6�y�#2���N��z,���D�")�q�{�&�3r����Z�\����>����RI�Iv����gլˬNz_=�
��)�_Y�۸�4��K�7{��w���xp��B����_]�_]�-�<�]��A�FL�>�;-R��L�U�����5<�;y�j�I�����L�Zю��Y�T��o�]xF���]�lA�C�V@.�b���Y���pc��.[PIّuM�ʎ�{�en�Y�-]�]-$+��O���C�t <���u�I���9���y�r_�`�q��/��!����mO��QT��mw�^�C'Tb�­(tf�����T�A+�r�TӺ�茮λ뢕i��D2+UnsV[�SkiZ�E��8�W�B�hٌhz�]�!�ĸ���H���ਗ਼��sB
�Wy~�.�!������!�Jiˠ��a�4����q�������Hf��^܉K�,�ݝb=y���+Y[�^vb~�]��2Il���Z��^##]J�b�U�N�a��V�^n�e��G��-��`��K�u`�5w'r9�l{O�t��޺����S��MID�[nV��b���T��Zj�Ӵ WNyJ��[c�u\��jɐ;����#���}B��ls�9(���E�n#&�v�c�������>�F��oh �����#����Iy�c���v�fV�2������n��,�'P�BB֩,BT:P)���F8�vkkmힳlH�ӷ���JM�pd̶��z^����zW�-Iݭڶ�C��n��0rV7[;[Y'^���{x�Z;6�A;����%�Kd/-�b�,��y���μ˽�yy�^�aЭe�[b%K�`�qe�E������,�
���v�[,����m��q�$^��{�'b���/lqydmm�Z�m�G��e���yx�����tYf���l�%��� [HoT��T����-�j�2[kbɎ��G�^��L�lF�Z��tSIH�S����Y���[�TŮ�� �9�� �P@������#6��̾�X��w�R��� ��H��ݤ=~�}��E.��ܱ�C�\����3����:D��� �ԁ �� ��A|F���
��E����!W�<���d���𼯸쯗4n�2�������g�k����ݱiHk2�JJ]WJ���e�oTmj��f�V��i�K�ބ$t� � 'v��~�A���Z�o���P��ui�W�o�"2%�]_¤6>�ئw.����z�*
�~��myys��jYu�m�� �� �� wkv_�^��j�H@}�#�_gW� ��A��_nбE��ƴv�Ws;B��"�f�^WN�_�#v���H���,U���&YT4~� �r�?nе�&�p[%��P�t;㎕
*�pf����X��d�,{�׻J*��N+5��R@�-7�N�yM~���|�N�gv��-����I�cHr�Sn�]�,.�l�6==���_
~?{�!R�Hn�Hj�T����}��7�(U�k�����K.��c҇r� �A�G���7�ی�c֐���-]A&��3�f�C$�]���l-,��^��M	� �\��m��ݯ�n���׽����uJ�7��2��JE^Õ��؂��) Av��n�$n�G�bU��b�@�:
�3��8-}yNT"���~�@n�q�n����@���_���ub�6(P����*�k)x.]jl�jY/�ۖ=8 H�AD;�����y���ޜ�G�3�mG5����{ڍ�_gT�����vR����!�ΡBT�SF�=?Hj�5(�7P_�wz�_XI+�qyO'�:��}���9P�|�"ǝ�]_��.��\��E�cݱ��	Up|��xc�a:cg ꙳UL�1Jo��I8�3-enao�mLu2���5(�`��-�H>[�՘ x�q?��[�����Co�Y���!]��3EV�!F]��B�B��B"cD�ə�k�D�H�%���ƯmP��Q��Rn��4��Y���].&z�EeI-h;6`�:����h�E�chV�t[]�T��v���0փ]6�*6�i��M���3%�5r��.�.�%��5͛4&�E��K�!������!]M���fcjjn�R�DkGV#VMF{��?k�kt�i��h�̆�hi\v&D�exe1[]��6(Մ*�[+���D@��@��!���=�,��_��,zrC{�4�5�:Ƶ�J���A F��b�n�u�4�Wq�q�V��g���_gT��������K�A�#v�W�N_<;�oNa��&�r�9�X�9e�Ct(Cx`F!c�tZ![]ζ���e�9P�|�9)z�����(�.Ծ�����˚�F�z��ρ�����Ow�K�m�=8/��Oo���X�~��]	СUR.�k�f3�7�� ��N�+E_���UC�z��
{o� �	���f� �g��Ҳ�.n]�!��T�[{�$�f�.����U�K\�R4��S@��M�;��47i7k�}��A�]���*{_U�7wܭ�W^۸~�Nr�<�#r�G�{qX���_*vN�l���§���gP���G�����/8���� 'z���������6��UЂ�E��˳&]kjK1���*�������=����w��<��V�qN@��� ��v�s䩾,/����7�/�u A���K�7P
{'�Ѽ�Ψj����b���Ć�Ć�Hi���C�~�C�k��F�|���� �.�^S���	�K��EN��1��Ƃ;��v� ���ݡ����p�|�
�!����:��Yui���?��C��K�BK��G��c3|�h�ʺ8�
#�R����@άu%`�$�[�+��@�6#`\�>�~�K�#���}�7PK���5���:��g��8����y�.�J����uC��+�$?X��e;%�l�e	+�&�����F'�o�)ʄ^�@���C��7w�~uꏷ�ӽ�ZH#% �~7B��V$5b�	H:�Y�uf�^�6̄�v��R� ��n�4z����µ�E�]��Br2n�u�49r��yL�S��ܮ�g	�U��YY�\��a��n�qN�nW�tA�@���7W���f��[Eͭ ƾD=_��S���+E��J��̡���_����O���'��AO:Dn��v�n���s��*�C|���Z���j�S�������_!R]�$��Mu����˲#���m�6��Y����&�dk*9ԛC]ZM3j3807	�㯔�;� �wiw��}��_��n�ޫ��{�Ebd��<��P�R_�*K��T$?fz;+*A�����/P_� ��y����:��g�(p ����Gv���9>cOe|�'z��!�*K�P;�@f�ފ�uN9��YNT"��@��� �/�#u|�;�/��}���4.�N�����<A���~�ne��tn��Cӗ����Oޫ�~~�3��,��e�a�j�F���P2��c;)[��rr��f�ә/lx,�c��ʑ������rm����tj����|vW�Z�������#v�]C�$`A�A|�_M�X�a�a�̡�N�Ds��ݠ��Hc]^^��s��P]>
�0��8ls�1-�m��␶;1�s
��R�X�H���\+;b<ʗ}˜�m�\�7����}�/7֎��Y=t�ҫ��cGǰY���SU�>���Hj�P�MJ:עu�����e��~�ne��tn��Cӂ|@C��Y��I��/;�y_W�K_ Ne/�?"�f �?f!'_������y��`[lg*X̮ ����5
���Ct*K��,`���7n@��8������v�ݧS�/V���?.>"��ǹ׈�|+��]T�P�Bm"ۨ F�z���O���)[W��(�K'���P�-�I�nP���� ���*�}!�m���������j[S�1��ֻ���qo�iN7{.C�IG��3f�쵉�)9�u���w�����F�]d���	Ù��Q5b&��.����@�n���ċ�lE�4ړ5������÷ 70ͥ���c6����v�í]�cdp쮉���w,V�`%��NBӱZ�]���L�4�m�1�:V3F�`��f�`,����j�Tm@,�D�8(h��ױ�2��su�@ ��(�$�0(@ît�X,v�áu�ʸ�X@�P���11ͫ���������.ԙ]W��*�i�5s����B�����f�!�3.�7��_����_/��AsgmE��Q~#x�ϨU�Y�גC�r�	�W�� A ������"�;5�L^��go=H�s�)����v�'�WZ�������}�F����*��� ��ݠ�#v��wi��`�ҋ�6I��~"�؉7��9=A������wh"7R��Z��6!�Ҵ�q�y|wPR��ڋ(��gQfO����R���~lzT����&� A� F���A�u�G]������3���ݤ�+Z���u"��"C�-�{6y����@
�X�Â�Ѓ�M�bVVf�5�\k�MPq.%�A����f�c����>�6(o��!�L��Aza�M�&�C���4l��yS���9��G��s��P��P�ݚ^�ѡkOId�^ j/t�o�,s���G���t+�� y7��#��0�r��M�F��A�go��/l�UH�︎��؂�g��d{Q~#Grlת�<~��4�"���۾��Zsv\�j\Fs�9��s�/7��t�ܮ9���.���/8/�Ԉί��/�h wk�y��u]u��׈#�A���ҿ{}���n��zܡs�'�_ ~雽�6�>��Wȍ�۴�#u|7O��]�D����>������s�k:���'�(p ��D�}�C���`�!�x��.��E
�-���F���q��X"�X����ki\.���iN�Ro_��=�R����V��*_�������={�a��j��`��{O�|�_5��A��wibt�p�Ȟ��9/��@l7�%wR����(p=��~�A|wjz����7���=���7�\�U�y˖��9�<�s��`�~f*x��Yw�7��w���8-!���5�]�jXK�[���,q��1����Q@Ǧ�_��*$!�,�^y-c�~��Y�ٔ8�� A腉U��*CJW{=��N��Ln��?o��G� A��z�3���K�]/9}Ծ#<��W��X��m|�?=_n���H����?[�C�����^S�H/L>�c��Y���|<���w ��"7k����>���R���"]���m̦t�ɢ� �Y��[4���q�#� �/��4���u�#e|��@/��C�G�mv��^J,���F!�>��|�EWC�5
C�	�T)]%%���\9������s�iI�����@�}Ԉ9������v�	1�-�D�u/�ݠ�� ��Z��jf�2�Y3}Cݷ]�nP���	�W�{�@�� ���#u jo��y����©�A�_"5����\��k����Г��?�_��N�Ww�	j��鍿��F�*��<�o���س�綱v��Q�ya
�͌���vrT�s:���}��h#F{�����U|����� H~�C�.�Hpȑ��w��?,�T���]��(^�}ԁ�|7|�u>�ֱ�^��h�E����F��+#�eܐ�5h^������Q��!�6�2i���=���A��Ć��
�!��^���<�{�j����i�^Zt��;���� ���n�����#��d+f�Ҫ�x}_-hr�}/Wo���BOx��A;Ԁ ��}�MVxW�r�Z���)�6��� �"4��3�Ɵg��֩��	(^��u|�V�7|�?����l��8D�Oq����O�Ho�J{��}��(U�r��@�<B��}sކ�N5�������?HU
�W��MdԹ�TR�'����sd�]�>O9:����1���l����r<��_��*.p�L�'A�4�mo�<W܍�oO��x��6	�d杣~�C�n<WC]_E��Q�����^rW�!{{��|9Wbe١��:�9��L����u�r!�i�1φ��~7�Z'����
f\�Ge��e�e��T��Fƚ~�}p*��Y6��ba�s��<t.f9���nD������Uk�����4���C؂��\��������2�6�������6{d]��'09-F��Q*^T�6N�.[Մ@��<,�O���r>��eۡ[sj�wO���ܧ��D�'�����F�.��6���t)8� ��E���D3rƨؕ{2���+[�f,��!�2(PD���l˵uջ/�3�|�P�$��&��s��ŗ��A����*,6n�]��{fZ��6�a�tq]��&�v8JT�|4�w�P��evڄq���@�4G 좯�)4Ѩ�)N�ث�k2�>0�]�m3�P�k���d�z�,��:���v��4�4:�|}Cn�L�+\4r�t0�X^��Р��BEu�n�@���=��u�(aA�R��]�҆�h/@<�Z�.��eȼe1�2i��j�1༽5_���ƃ߼��5��җ35���~n,񯧊�sJ����X&�u�3����h�-o�b-���XX��&7ur/ή�tdX=�۹B���QR;I�*T��a��w���<��:���@(
���bN+H�&�j�kvjX�Z*�q�z����k693Y�Nۉ)mmk;Nl�y�����&�ok���n3m����m��[ ݫ;�-��,�Bl�i�M0mjw���sv��{��^[mH[��4�KX�m��v^h^���q��dѴ�b�ŬM�ඹ�um�,��ܓ{֑{-�j���s�$E������3�N3[��lZ�����#�-mٳ���hmӶs4�M��4͖�M��5�6�Y�vh������S�8��؎v�L�0lru��cZݖea'9M��Kb�촲3%-��mm���r5��6aۭ��-�h��[��{u�zl[-�i�4k����u��m�P#���6�vd6��f%������Gm�gd�ò�Y76Ŧ���4�N;8ɭ���m �lݻS3f�n������f��v��f�ŝ�u��qkv��o^ZB�٨m�_n�3m�ٵ���4��.�5��X͎b٭ʅ�ڕԌ3�2.P]H2�(A%ڰkV�p,qpa�����SKh�r�Xf��ؓ[k����ER%��5 ��5)t�����Zѥ�V�br�b3UMԦ��ҥ��a�P�!���Ѻ�f���u��Ԇ"�R���&[��*ܑ����]&��Sm�]s	���ԭ�%����i`���@�&�YHP+@:�0y�����ak��m��b�o$�նZ\�sL��a�Zi�f�K�4�׼KR��-�a)txk��k�u�b������@ka�MP-�Ba�m�6)	�q*cYM�&Wk�Ae�͵b�CJYT�����jnu�̷e5�2��#�V�:�iײ��չ`�l�Ӌ�P�b�mM5R�a�:�h�أSheB�lA�SR��ic[	l�����QDh���uԺ�G�^.ұ˒Y��7M��@Ю���i��k����4i	Y��d-�"]��e�ͭ�Wb3�6�r�ؔ���b*���r��qj��T�i�vc�Є��5լ˪TJQĆ%k(ԡp�(T�e�\��!C����supb���4\շ^"�c%v1%�!��K	r��a�#v��U�5%s-���6�ƉXfM�vG2�)�k�F��%W
nJ��,U�\ق�t�`j�[`W�+]���3�*�j����H�vF6.�`�i�հ����bX�@��)�y�*�lqx�t��ٵ��$f�]t59[�be��;c[L�\�F+[t��1���ub�ٺ%us����Kp�9fM
!��4u&�qM�#�M�����b�59�b�p�k�yR���]v�YYb�fV���/gGb���5��kJ�2$υ�4*�q��5��;E���f	e��+�mn�u��3]6�v�i�vt���6ͮ8��.z��`&���)(܎q.�Y�k�oh�/Cd�1����]�6יt��
�,ĭ *���W6���rݩ�D�ҚB�:�`�A��B��)YtW��ԗF-�IfBR�\5h�X�֊�TFVm�%���#a�-�$6t5�j�.5K�"���i��\h��J`��]s*�m-t%]\��幙�����+*ԥt��^��X�8�i-˯0����l�j�8����K�O,�w�ȩlYۢZh%M�n;hK�T�=���RP6�V�Ճ"y�<�g�����g������CD#��lS��ص���˙�\(�� �=�m~���e����=��=/��0U��7^��C/ˣJ��d5�d��V��n�
#���U!�}R]X��P�!��`�~[�T~~�c�| ���x�\����9B��.p@�g�_Gr��Y��b���F�_
J����
�R��/�gp	۾�}W�צ��z� w�D:t�'v���ؽ'X���Ȅ���/�;ZB���έ������/{���#�JoN	37��؝���G;e��q��z"&e�t4c�=�Ϳ?0��R���g���t*�B�|�����,�H�n���~�~��l���zo���ԕk)�h7BSZ7cn	^�*�8G�͔���[Bo~Ѐ�H�\��!��n�	ou������'�����'y�.a��T�j�A�@N�Am����n���	�][}j�|���Z�xQ{�t5(��F��DS=����B��B�P�b��쿏to
�oI���NL=���mr�^->6��璹C	���:�|{�)�fc���{&g��.�����Co�/ʌ��l���2���v�#�e�e\ƥfK�W�"�[��}��(U�r���X��E�3���eKs(�L�֊�P}w.
ֳ=^ ��9��-����_[��>]�;`����/�0[
�[�r�{Ɠ^�`���	�e�fQb9��@�_����9�ߨ!�s4��<3��3��{���K�	�@6��?6��Y�m���XeWA��)Y�J��,m��J͉�t�Ql0�fm�1Y�Y��*������!�׽`����W�{�h���9B����WC��t�؝k~<��o�C��Cn��"8�^=N�ʠ�_��h)ou�����&J�	��`���b9׳�]�r��Fj Hޠn�n��[�t�C{��X����٣!5+�.�U./Q�}��T]��5r<��΃�m��~��;3���yO*���˼.���W��3w�ufuv7X�<w"���Ol��0���{����A۱�A��+�Q=��[倃��9H��W�c�kG����
�nP��E�D�ju�޿wiumذKt��CmG��i�Ϲ�����-�m�]�;`��?nE`��D!�@�[hj��I��T/���l���������JVQ&ã���,!�M6[�V�UPVHw� H����7XA��Aw������7-�E��9V��[���H?������ �Ց���{;��-���ѫ�1ﵣ�ݽYB��.p@�/�/� v���V��޻�/I�Mr���A D�b�<���-�_ۻ����sl�[{��u�gTȝ�0zWN�V?tA|Ct���Vn�����ؼ��c� ��>�`�_ t���u1�8e���fw�{��ly�Ѐ��~\��Wb��	D���Ҝ�^Y5����*޸���nH�i,�Y����;��F�✐]�x�]�P�Ff/��h Ct� �Ր~m �m֎CE���M�ƌ>핔*�B� ~_P@�;zŖ�Kt�H�<���~~�||�g�2� 3f3��e�m�)	f�X-j�vٗX]́W����F��?}�۱7A �澷\���Kv$��\�a���)�,��1a��KmX!��DG�����ڦR�<[�(w�����lܶao�}Ԉ?t�*�j�xM��OO��D?R�Ⱦn�� A������E��6k�Rn#=OL�+�ܡs�}@.ޱe���tm���8��I*��o��������\�G�&��@;�X{2"�O/7���ba�^��~�j�!���۱e��|���{�J�0��O���~�o���7�����<��� m߅�w(r��t���E�SmEG:�(^��G5��V7n���^oB���"-Q=��T��f�n��t���Z�'��;����������f�PpG<ݰ��%mX:���װ�U��J#sj2�4�c+���XJF[\��
ᔴCr�,K�!�vt�t.�WiI�,�Y��p�b�Ճn���XK��Ző��S11[c(�5�aVD�I��&�&��nF��^�t�&���P��V�daH�hWF#�ulhC31-�tl�{	CMiV��Էa����2�+4���(��]�G�5ehɭ���Be�#�q��Ͳ昀�ME*Pl�o�!_>�B4����֬}������i�"���82rq>���4ט�Am�`����E���CC2��������������u���c�\�;<�V�	0d��~.j�A���U��<�u�A��+�܂����n���W�-�`�ա��fI����� �����Aw��@m|�?j^u^�b;E}���. ���|%���ߘ���^�������6����IP�B�-���!�53�W{2���Ԓ	voJ���=��%量�j��#���|?��5��R���h"KCp��X�͆�J�0���q����f\�XMnJ-&ڮ^���_9b8�X��wF�2�+B{=�Pp���9_[�}��S;������Y�}m��,��?6՟�p`3�_�س�"�f��ࠃ����$�)ћ�[��ɪ������u��%S;G�����(��ֻ�W^���4m'�5��K��XC�����X�c�1���{^���&���b�u][�Dr�]�����Cޤ.��݁�C�=A��^�}��y����$�~��:P@Y�ڲHb�^�`^��f��F�`�� �d)�����X���~�,}ԁ��WA=�;];&��� �,�?�V 6�e�������|nj��Ok�\7���nP���! A��[�A��!I�ܒ��j�����R�� 6B����9��6�Ɠ9MF���wP�i��JE��ź�\B!��n�K�c87}GN9�Oa��#u?u�mt�����/�|�#�����X�pM�_��aeӍa]�:d2����;ǂy�1�~�hp>�DL�Co��|)�-}����ݶ#���D̲��FG3/%VlN��'���Kg�-�7ܣ�:9��QD �pa���r�[�+�����.�K�I�R�]����:��מ�����!{�.r<B޿�����B ���c��+�>��U}������h%=�������sD��A��f�מ��^��7�t�G����_�B�n��ǳ���@�W�՞���᷹3����>�@�%26�� 6������t>���ёU��h�F�FU�U�WP��&lFf��jB]^p3LgՄ*�\㇁�٪�/�@���ڼ�?k��;�{�.w�a�`���F��<E����c�e��m�ЎeJ��N��w�^6��9�+���857��af|A �j�}�H�qX���w˃Y�\����:a�۱`�H�3����}�k�WJo�z��Ycof�ۇ�[��>�@�)�bff�FfYq��MP�׷��V�_�p �_3� ��W�{��Ou�ኽ��+�a��,�-,W36��ǚ�B��4.{n�˩yh��[�aｒY����f���Rq���d(�Y2#�5u�&�zZX4i�8�.g ����g�ܫD�u,L����2�&8�7wG2����+���[���4I�0����tAYD�^���g��c��
�n�Zᄥ�ԥm�B��iJ����6b�b�Lj�ba�3w�쌷�팲�������e��g�9�<�n=�~��*��ŷ���Z�a�V�A\B��޿���Y@��VB������>0�lW��?c��o
��7(\ླ�"�ł�Vhu��H0��d���1����B!�_��в��ޒ��������&�3?w�=_X@�������'���6B�v,�]2:�r��y�q�ˇ���>�@��f6l���9�5�sSݢ�n"9�z��\�۷d�ͭ[��v���M=�v���7(\��<B8а[�A���VW�/�����^䳦��B��z�h�]sBU�`j:����IPV�`��i�w�� ɽ}��c���];�T��8߳�F�19�|S�=ng��ڊ�mm쾦X�T�lѸ��*����tB������[�J/.5)E�UJfls�Ɲ���-�D�v�R�JCj����I��whF�n饀\�4����4���)�
�n�u��=`�Ų�GT�u��6"MM��\C��ʮ��"M@�M`3im�.�LK6�f起�qQk�\R���S֚)�b+��,��4�:�^cMZR�F}����K��E8�����e+eW���e�0��v������uqҵ�a���=V�k�i��-�9n��u�b�D��#���z�W
�s�4g�,q���e������6���pø�[���B�峨��or��m�A�W�S!pJ>w����?"�h"�(	m��s0�f�
l���;�s'����}�<@A�b�t�?:d"k���W~DJ�׫2���]����R�5�1�k*=f{�	����$����xi����X!���D�nŀ[�n��2-��=�8�j��ϫk�y�������`���Jd"w7CNKk�X}}�ݎ��0�iK���B�:�a��]L=P�xڈ�͚ۊ���!ǯ�sO�4�2� �ڱy��L�;�p>������.���N.�(�A��u"Ιۻ��}���<߁�oĄ1�^��t�-]�����ׅf\��:����]뻽��Ȥy�*c�
���'�ǎen�9��a�
 {�o��[��]!��*��7=�����P��<��v��ܽ��=�~�}�w7�Ō|�,F��Q̫!�!N8���r��{�����d?%�`��H��B6����Ye�}f��.���ya������Wy�͙�w��o��=;�	��")ޅ<TY��4��z0�R ���D6�X%�D鐁���+���U��A]���R�yV�$�0�����DŖ~E���t}=^h�V�x~8�՛"��*�rB�P�����Z9l3�YC[�����Ge���:Ő� ��Ŗ��!{�}��s��2��6�mוR�Z������ F�_[h Ye�m|}����vn���a�A����c�}]��.���C҇<B ��b�-Ӓ��{C���W�#f]�_R �L�m��Ch`/]�Q�Ye6s�<�"Le�s+Hf`�i��[zơk;#��X�(�D�.cEgE�:t�8�И}��*�(�x�ht#&K�S�(=k㻚�B?;͑��v�~˳�cEK.���f�9���9i%�%)�G2�*β7C�%a˄���vv�6��D����^���G���*��x�f��fvi�С�/��ZT�x���Y�N�A`�y{,��� �0�6��ťe�f�v���o�9��)m��	��@��H�i�m��״C�۬�e�chD*��tܳw�$iM֙�wv2�K%�80�-����~eʳ1�|�Z��DG��7dj���a
�Uߴ]Lw8U��-f�j�`�³L����[NK���[,-��سf���)JyNu�:n-�VQ��˯zZ�9v�d)r58�9gM;��0�Xe�i]*���v�����&�r��I�M���k-LWx���aR��za��{��fڕc�N��E�˜��T=7�Q��c��ހ��\��7U�M������Fo���_!%��{��[���7�ڶ��o+�$���BlFd�u
���.�5���:��*5��%���P�nd����ʀ�-Mp�3U�JԠ�uuJg#`h�Pp=�u��i�s��ژ`*ý�O�Mv���7�",��w��^C٨2��^�R��V�qHD�*�ю���v��B��(��nfcw� �Vn�Pt��r%Û�aخZ�ۺ���;
a�L��\.��e���k+�7�]g�iS��`�ͨJ��X��5�M�)�n��+����F�5�3+	�@�8�[k6�e��p(���m�f�m�Li��f��6;m�b�l	��P���:��9��Y6�&v٭jD�6Ͷ36͌G2�F����[k�Ӊ<ܰՖ9�gf,k2���0��Iŝ��m�l��C3��D� v�kvI���kv�+7l�����0&sY�5��76�ݛM��i��:s��Q-��e���=�<��Nݚf����6�k���e���i�v�Z[l[X�De��V2<��B	�ơg�������v6q2�6�Gۙ����k\���2�f�ccN�v�l�M��Ѭ���94ŭ7m�3':�ä{g����n�m��응����쌳�Kr-��[j6۶��+kv��)2��fٻIY�;9�Y��m͉�mm8��nێ-kvݖ�=���98�6�6��DI��mh��xk6fl��F��@ �	�_������cnxOdVGJ���Vm!Aէ���e�_]2,�;}��s��]�VP������W/y����z�,��%��Ch Yff����k����/۾�9y��䱹C�����H�鑷�}��j�q_p7uUDٶ&΁� ��]k�Q	�ظ�Q���Λ<[��Vh�}e�D��mؿ�����}"G���ě��=S׈ue\��׮�#;�[�͢�e�&e�1��R^P�_��R-e"�B��i��U�w�2�gJ_D�B �ܜyҽ���w<�؉{ס3(�m����+׬T�n�^mg�Y���l��;e�-��:d�E�Է�r� ��!'u������7_H��/ƶ0���=��){h�ؓ����~�fb+8�j�3;�!fR�&Sdd����gR/|E]V�l���(�n#o}鎳v�KK���|Ag/�ϐ%�B��۱e����;�z��P�����N�Esݷ�ֳ��A��"T!v/��h-��+`�cFخD���HR3M+�֚[���I��R�TAf�%�#��n��v�Ѭ�p{�����Yn8؋���[��-����p�}�/��B��DY����"�B!�v	n����{O(��0_���@u���<2�ی9�0��W� ��,��x�^�f���v-#9 K0��C>-� ���*��E�i���U��3c��[�PҾ@J� Cm}m��e�G���N�5�G�A-����{����\#�� #������w�@���6в�/�!�!۳����|U��$�.����0�ه����:PE�W���k/J*�u�te�2 �}~�xWb�:�7ƚ�Q~�]u�/����k.Z>�.�::��!�Xy�(V�'��}g�z�-��y<i-ti�`���cS0VM��tn�C6b5��t)0e#�aj*���faC:[s�X�j��݁�]Ea�n��,� �:�:0��3̬��m�l)-&�FH��@έ�[[6�)�RH��̫�ke+��V띕���͖�q2^����Bl�Ƽ���b[������Mքf�aҺ�Ta�c\�YT
��#n�BY�g����Ai�\�!����LZK�r:��n�Q���qS
�ﭟ����-�!�B�sO;�����C��!m��6g$��u�WR�~{A��_Ŵ��ڰF��}CaӚ��":@�����t�m�Ҽ�l�c�/�/�<�-�}E/e�]�=:� ������@An�!�b�n�>"̼��R�5��>�6y�4\� �z+�"��ڲ��ؔ�&�=�8}�b����S/���p\���!���VP��ʾ�oC/D�T4�WM��] �x�[j���D7N�Q
��R�l���M���?l�J���F>@�����X�� �}�u|3}�=�<�U�i7k.2eβ�$�$$�^# �,�[�u!���y�M]���`��@��!�b�!�cs��o�,ڜ���g�u���[�F~�e����G3/Q3.�3(�5�}o�8���ô1�[*���Kʐ��@�������7���6�g�+�m]�}+���̥Cz�[�p�X�u3�۱��1�� A��P^���~�i�ov�{��~>�� �Ak{M9���K�;[��=ۚ3,�3*�G3-�{��=/2s��z�z��G� ~"���7X%����c�j	r
����A/( Cr��A}י�$��|�v<u4\� ��VC���+�=��z�?�Vm	�@�ۿ��㬚��;�^߰,5ib�_/z�sK׳���ϗ������mA�����>J���Ig��k�y"f2kE׫��mR��IcsW�2��X��ZQ�+�?A��ބ�Qi�W̽��N��o^�����B�=��1�4_P`GIb�u�-�@��� �H�n��* ���Cݻ�Ȃ���$�¼�v=u4\�����y���Y�iV�H2�e�#r�#e �n��[�A��BZ��*��gK���>�]P-ɽ|8�x���Qn�8=�s{��+�M0����!j�@ͺ�.	��7��{�c54սfӜq�N��85���藫()|~��!����@7^#+�Y7�o��w�p �� C�@��V}�r>�������r�� @"��o��s��*7in��j�~�E�Q`��s2��e��1�C�1���ך�IK�������n��ފ�#� �x�i	C�9R��P��]�ǩ�].�ı��7j�ju��,(�utlƥj��Q"�ݔB��T
Dt ��ز�/�%��}���J����?m��<�R�^�ܮ�g�,��MG2�̫�.f^���̲�@OS?djϽ�A;}���~��P����N�,�XL�=��ݕ����q7��Џ;V32�355�9�y�� {G�=�����멢�/W|A�7H�[j�!��U��j��!�B�:�An��o�߻��;�oa�}���җ�]�����4�8(2��E��(�Ȳ��=J�d����sl�=�\�C�)L�v+�.�76D�3z9d��{c-w���[����P��㼂���-�Ch CuCw�{ΊX�AW�/+<�p����ۿ(�Cς���N�,�HC�f���|G���!����~K6
��V�Zb�͗d���f:��#����-,C;#[f��ٻ�|�B!����A}/3y�[�멶Y���;��:JP�k�PFQ�[j�mŖB��fk���u���<)�٫�a��g�W^���B6Ե��η��|�/����r��AYD[k0蝻t�t��c{}��[~��C�_#�3���DL�Cn�z��g���qJ`�+HD6�_�Щ��k��x����,��{�X#�<������:YD���Ch	e�mؿ�n��\��ڨ�4Qdz�v;~���޽���>��?J����У8�L��)�_%�LT�^͙_ ���5����7n�����v��"���0�<��(+�P���d��Kq|���<�k��ƿ[3YVyD+�q�lDQ�%�M����*��h��Q�Ff���.;+4K�D��*�&1m�nn�ƀҎ�7 �.t�ɫ:Q�	@1+ln���Ûjmu�f���;!lU��"X�j]]s���].�&�j���V�f%v�r�2�Z��:�F0�Ԗ�1���'�m�b)R�Yn����M�Ș���rF����]�2�O�o���۪
XM�Q�ͭ�Z�U�&�Q��]�U�-cJ1űu�le�|x��W��"�(Km_������~��C��y*�iZW@�"� �m�-� �d Cnł[���vs�]$է�x1��Ŵ���\2{�n���Oy���9��g˷�{F���������ڐ?aCn�n��A�����e5���n�-bU{S�γ?~�hG}�}���fjj&e�qؙ����/޽�&#ڂ�A���~�ĝ���7ޖ�������,�1�׷����/��L�քs*�&V!��7����%�oHb�ި��5{��y���u�,�Am��UE�$Z��iR��Bg^*�kŸ���2��`��2�E��Mi�V-Y����v�{ڙ��"2�w<S��x�����X�RY�˩{������e8�q��К��wq���R��[���"L�J�nYVr����D�v<F�X��\��oG��o�	ו���٨��
���ֺ4�励YS�=B��N�Ov��z��o����|���:X��7��ؼۮ�[KMw,ӝ��c�i�����n����'}�["���\2{ճ[3Qg�1��z���,q�f^�̻/[����O#��,�K��B��y9�8�x��?7�`��K�)Ѳ�i�::@��IA�? [j� ��e�M��g�Yچ��U�'	�&u��E���_Y� Ζ,�H��-��P�U��f��k�	fH�,�$�(vJu�Z��CYG�I���e/�2��_[hWf�FZ�3ޭ���E��k�~IJn��N�
���i
	����	��9�;���U��ԁ��R�Nx�4&={��X?:@�$_ Co9�gk���%~���A��v��Am|�-���|�u�~P��4e`�q>�y�I�Po��nF���WG�;�� �̿_\�c�=�w���ō�+�Y��7DyS<�|�X,5ϭ��Ϟ�q}����� A�,Yn� ���6�Þ%xwj�cZ��{��G9w�m�o9]������N�Oz/�����zro��Aǵ�!�%��nł�a��`��_%��yNhMz��ο��~/�o�Chc�ئ���EG�����}�5�[�y�%�$�UP�N�Y������֮�(�VQ�c�=z��.9�Z0���o�X�������	o��yw��&��:�Am|���~-���g�?����X�@��}o�Jf�E�)ZٯL�Y�A����A�̲��t��5M�wy�;���`����ǈ@�w�u�u��q
ط�g��w�<��*��{��|�/�m|��n� ��KJ�x,Y���Ax��레 �՛��ǻ9��g�M�ag Aί�U��wS�+ �MZ���I봞*���0�b�y�u^�a )���b쐂���w����y[6������OR�cn��D�<�4�r�d�.}��C��!�b�n� �������{p�6�ݿvP�ݲEM����bb,� �{ܬy��,�	m�{A�Z���=Ua%��v,�4����-�6����Q�ДΛW5!�jZqF^���C~��,�A���H�!�2q�8�ُa���t�
�˻��ۗX!������Y� [j�I3������r���vs~�g�͸��p�gK[��̫uA���ӄ`"ۿ��t� �2���-���K�_G3����t�������@7ܬ�9��e�%����!x뇽Ή����A�����L����tُ����|�#��=$~��	oo����m_��_Y\�KZy���y&V�p��o���9�Y� N wD0�H��~�|벧��>ں�E��vtT�26y���#������/^԰2����SbAU
vͣ��u�/����n��;��c;���fQAii�0IFy`��b�a��Z��:�ywV��V@]Gs2�M+�Fu*��T�+�Z�ꖴW>���gC�ٞ�8���z�4r�JS�����^o�d��Wr�6�ձ�$���r����,Y޷j�2�"���z��m��b�ˠ�v�%�WMA��C��o�����C_��I��|,�]���KCV����~�v�1�.ͥ�0�XI�}����9Ug�!��Ot5�q��W7��tnb����1/�[{�z�U��q}J ۓ]K����R�eL7�X��cC1hߩ#v�9�o[�$7KI}�>sf����t�R���꫿Ka{0�v.-;�/6:�B(V����"�gF�%+[5�轠�}����:��f�tj��4�R��񔻹l�Km��.4��cc�9�Η(,�{�N�󓰨1m�m�GIw�����ތU�׬ݘoJlW6�Uȥ,� �>���u͐�U�V�Ε�����
��b��$T�8�B!�n̖2�����}e�Vl�O�]��6�B��~����-*w�e�]V%P��1L����W��d�%�+$}�J�~���vjfqXn���'2r���i�Gm�Ȼ�c�;�Z��+�}���:g+2���Ѵo��#��P�W�y:��M��W��͑�g
�q�Ĺ�鱽e���&j�ͳ��t��Y�� ���L���oQ¯ ]gz�}_Y�p�%��r��ш3m���-�s7-��r��ʹ	��k�tfX�۷"s;m�I����٭"p�=�rD)�͵e�&�Fa�R�s`s�cfpź�[��e�C-'3rm� 9�,Tq9��Oj܃��m�H�$m��7nљ���yy�Y�S��s��hHa[5������d�pt�:���GD���fs�m��<8):B��vi8��t�u�j�����t�C�m�F���݂r�p�����8��=�=vI����	X��FhH��m��f99JA!" N6�#���)�۸9б�JD2�q�����^vG/kH%���h���ì㜅�8����33������R��r@FV����5�����m�ցm{���C4B�jJ��6)ff[�`��xW������L$�(j�7L�m�Yb��U!�v��O y</h�5Cj��i���k��b���2�8FV�F�.��2ٲb�����4���"��%��mդ���^oZ��˖Lö�3*�b��i���[x�9e��I�n�2��J]�T�0)��V�`t�	B��B�0�hե��LRڝ�P�1t�H�B�"V�k��m�Z]eS$kkؤ�6��b��ZB6��6.���F�u��&vaEH���k1��L8�lJ�u�²���W�ˣ�mW�[5i���Y]cC��k5a�,��=bK^�]�ٶ�	a��;&6�n+A]�B:h��^6��c5x5CL�D�$uY���C�ul�5��-%��6n[6�:�XB�2�.m�A6��`]2�֪����Z����8Ү���meIu�+����!�Rmbm56�M�էA�㮤i�ا<W��jM]-Ү�Jb�,�w;�5�h�Z�K�1(X8��it��a�Ⲑ̽G��[�h��V�JTpK��[��SZLx�@4z�\�Aj����K!v�4+(嘨��.%���uaa��ȧk5�[L�$J�]n��::�@j�閃,�6в��ۗ��YQ`��t��)-vaC�B����Zj!����.a[TԌ5ЛS;P�2�,a���ۜi]dh��j�s���nZ���M���X;�l�AQ��`j²�����1����-ļ�Is�F�.\*�])�9�)*��[�fQ��nRں �D.x�;Zh�l� v���U�*�hͳ�T�#���hR�S`��G��]tmZ9��Hae!���[���MM����V�5�6&�� ��K��0��CJJ1tt#u�_	�!5,���)/d��k`�p�]�V�)Tt�Ҫ+��Q�1X�*2�f-���Ķu,�,Y��,�o9^ėA��1np��XKV.�f�@�]SdtWF��m��)�Wb�d\�.���]4@��v�bMiWCk��@��AF׆Qg���/��m��mU�#kj,(2��Х���E����v��i��rT(��v�`�l��*��]n��:D���P�����s�lC5��L����\-ub�4a,z�*�{L�͖+�m�赙uS�MJ�h@^�ε6,�X��S��pF��u��)�̪���q�jL�_~����Z�j���4b[e���l4��!lf�3t�
8���Wt�(�q���1� �\@m���m�sqH�%m�G�O#���I^�}�U�{����e�q�"9�zL�,A�ѕ잵�XT�|q��Ae�wA^�M�������J� m�U?eNp��CW��q,�9��6�������w�7O���z��Ǘ��r�!YC�ӥ��g��2!�v���|���Z#��&�}�.�n)d�W����8xA�r�\����K.=v� �D̻��Z9���^?5�7���難ޮ"�oI�{�29����;������B6���ꈮ��o���|�7,����4�Ꙕs�Y���q���4����b���VM%V��8~�٪�!��e��ڳo5�]��/�ƥ�B���u���,��drŝt�?�"5��~-�#n	�X��o�rie[��Sx�kH��rW($�xg/X�	���q����T�c1SJ����-;wu�z+��ru�x�yҗ^�6v�T��Y�
������5s��W7ܾ�h�C�T�ެ*���&Gb@7AnŖ�|A��A>���ye�%�����l����}`�})�J��_�6�!�Dj�P���v�A3W|FeԈ?�VS��'ok���Ը�9� 7�[�E/nߵ�+��q���۱`��"-�@���x�	�0��@I�zrq[�5=��K����+h Cu�-�n�W�ƅٔI�	WH50R�.RY�Љԣ+��lLCKhʅs-e�G@�_ܧ�uA��Yn� �� �=�����l�nW��X�r�Bo�W�u#��A�n�ڰA�(ܒ�wYִ"� ���_+�oA;;_��ƥƁ�7�"t�e�W��Á�\=����Y���A|F�w���[�d�d	���Xk&^t�{H�Ci��R��b�v��X|�Y�U������X�k��:KA*�+2�v�ɜ���T�f&��AS��İ�\~�r����!�@��m�!������	P��e"	n�o=ޙ���H�ל,�H��P�K,a��z��32��$A|Ct�%��Ch/�n�����[�bo��^.f�'{����Թ9�F�D�n�~-���9(���wh �����U�maV�dnt�Y�ӈYCZ�k�L�Ģ�Y&��m�E�vRd�yA��ԓ��
��lK��2��)y�e����#�/� �ՂA �����Ҕ�˾�S�;���A-��b��l��_k�8��P�]��v��y���FJD^����7_ [k��t|�Z��|��Ogn�I��w]���@�,X-� �����Kŷ2K����A|D�_Ŵ*gG[����ؗgǁ�+��/Fw	�����0<�㵏���$���,D�ۙ�D���U�yo��̔��De�Y�
�0]�riW��@� f��CE\�W5�f����b/���L�,c�%�n�n��y�2���eα6�/>��b��l��_k��;+�%B��m��G��~���(!tj��]&��m��X���k�3A5A�	k]6�V�`����8��h Ye�h<��\o��cR�@�7Í�����~��af�e"�B6�X%�@���W��8v�<^y��݋��gGM��"�[b]�{ܬ�,��\<������w���K��L���X��f��&��0m{zf&(�Ȟ����`���Fv��34j&e�8��n��96&A��a�Am��vA:�?_���w]� �Jw�SҤ0��g�P�Cn��An�:d�\���iͷ��J����7<^p��Y��	�r�h/�,���w��S�ӊv-�*�ڛ��e�-��L�Ż�Z׌�t=��7>�Խ�>վ�r��	�r�}�9�;�����1���LݺNf~�}5����6ٵl7h�C�DхKK��v��=�2ShR[r���X�z���,ي�����Ji�7m[SJDÂR"p�jR�+v,c�2�V�9�+feY���:�TWn	�\,e�u�������2�Dг�SB:�8�-Y�d6Jݩ6�ȭ��-n�̨�˦f�)5؍���]�E�A�avf��*��΃���T���=c�Fy�~�}�1
�v�XDJܑ�$ft6���)��u��X�̥4m7�|��w��1�;[�A��٘���%=��y�:������F���~���_��-��,�-��	=��-���_x`:x��-��68%wG�{�T��P㧈@�:X��-��;�V�����#{�+e��m����;�шN��M���F�^q����=�;|�}�^��e�8�1�Ր�C�{�_)��q�,�����f:_~tȨ�����FI)�_k��:�7�gQy�)�g��ܱ>��,���Ղh Yd�;^��.yZ+��*j�����W>~���r�z���D:X�t� �dh�P�u�rN�RGʓ@xt�:0/Y�fR�%����kP�E���M ��ݚ�"�u�c�A��!|Cn���/�?v��C_��[�:�!�Z]����l�g�h ae�j�!���D^zu7��{�羃Fyn]�/ ����Sվ�g��q}�XB�K�T�Ix�ϩTTq?ۿuVU������u�7�ĵ==�8��\�����FI)�_k�8����p����P����ϕ��,�?���C˺��A�^�/ُj�����nX�p@�%�>�tj9�,�Ĵ��M���^�g�]i|B#d����
k�[�/:�x��o�X#v��zV�Y�� l¾ ��X!��D���z����yU�w�ٯ����Sئg�CB�h�{E���52�t�6r|ԟ�r����A��ճg'�`�Ղ�j\�ڎdM��-+�RUh\�� �|�}n �n� �[j�n��W>����r�{�k�i'�Ή��lY}H��Cn�[�����}�A�3�hTo�͘_eE��!~���r�9���s�V�0}}�D��Nz��fe�ʴA�5����jT��%׳�a;Q�ܖO<�2�u�Xk�&�!6�Iy�j_f�]k ��һ)�t�%�F�Xk.%��� ����;�
���8�-2IOb���`������m��[@7^�����w����I�~ ��ux~-�n�zIG�n{��]�b��F���Kn�&��x��,{�.&fh��2��e&f~���mp�b���<��w9��T^9��/���o�Y��  ���DN��o<7�O�~���LT���,��V�Z��Kh���Vn1��Rh�6`2�����#,�<�G�#���@-�K��s9m�{/�y�����ʡ:�!�w�m �x����,����viޔ<��倽ގQ���'�*ܱ^��oPD�K���g"�R����A|Eλ��@�[�����-#{�Q{}��-��19��r����{ܾ��/�� ��V���<0\Y�ݐ�cv/㮗��t�<|�r�z�_���b��
��`4t��:f0X6����+=�Hzb5��Y�2��A/~�#���6�4���S�т����k吅�z��ƨp#7Wױn��[j�6�n�뮺UA��W�쓜��۞w��s½� ~#z� ��ł�|�t�W>/��t�]Y4M�(�d�YsiJT�nѬGk	`P��Ri��V�]+K�~�o��{t�|d�x/�A.{��1tSՃ\�~�"��u����2b�R��>-�`��"�)�����{:�,�i	ޠ�<��r�]�/���9)2P@��'3�3M�?x��!����u#�Y��@��[j?v�Q����>�&l�󼎓���#�N��u� �y��'�N�;�	�Oj� ��9�}�As�й��V�,�Y��?�_{U���Sr�j�Fΐ#kn�,���n�n�5:��&رU�+s6l�T3L�����zR��*k���7��Qh�y�{�/ʲ�h]�<E�^����	?Q�J�3ۗNz����]�pi��o�y3OA���^C�Z�l��z?6���9��t���*�ގ��6��t�1d�#�k�biH�B��40�,�Zhi�jb���s� 64GU��t�1vCZ5��fK�.�0��L�d�X�f�BxxO ��Cs��X�΃GC�	`��^[�Ay�M�׵�vK������-p-�v���J��K�:�!��6�Ͷ�9m�-RV���J�*�����R���Yv�M-)�&����Y��7\ ����n(�J�f,�ؖ6���;�ߙ!�4e�~m��{ c�ny�GI�
�!���e[5y��b,�=2ř)]2m��H������׸��,�z��Lo�sݐV���U�xA�E�JYg�򵂹�����}��Yd/�m�`�_ �#'oC��ݬ���שi�^I=���/�2�ۿ���h/�,�������z8��ۈ Y�@-�g1͂�ny�GI�
�:x�G]�(�f�y_c_gW�:���t�:d��ߵ�9���C�7;���[r�����__D,��������j"�1�;\�HQ&�
IR1m�[)�B��R�ŗ�n�˺���v�B&fh��U�M�����ʳ���۞�*9pN��]\Feq,L�kS2�lE��Оﺸ���P�<y�m��U۲��b{����r�, :��vͩ}���6V�z��Y%�D�,]���Ӿ*�������H��6;ݹ�y'<+܁O�b�-ҩv�]�w��ʴ�&��M�Ո�X�������q�JrU�a�m��pM;s0�g��X ��"�(�m|�|��>󎟫���G7_c�B��t�뺭�^G7��}+�@�_l�YڲN���@�� �[j�!��,���<�YK���r���xA���;����^��O�,X-�̲8����AOeњo=E�Ha��Ҙ&�i,³EȕԀE��j����hsUf쪿�׎X&:@���������������ӻ�=B�I�^S�;���,����#���̹b�h��Ǥ�Z�^̿�S �B��Ӧ�Y�ގ����`��/�"T!�*�}��<����������2�8��֏���]x^\�޿)Sm���=�Y��8�RiڒJ�Wy7mπ�o,�a�2o_`�d+��2��T�y��I�*cu0�ϳ�(nxyF��Uv��V�\Ε�.�
�L�nf[��` �C9,΄-���é��in�W��\�VtPWm���K�a�1l-=���7z��ɶ>s-q�{8�@8*�h�I���Qϗjг8r�	��/sk�%-o��5�Gw%|��r�����Ǣ�����q�'M�uq�èh�	�ߝ3�^)�sSR`��Z�9���UU�g:���&����^W�%Y�I{Hгػ9�}R��4�$�	�1p�47�,��︷�j��ES�k��V4��q�Шmg�͙��
R7���xA�4k�����}��8,e�gW-�=���s"��]7�k+lvj�v^�w6��.�b�n��5�D�����Ou_��^��95M�)��l:S�o���7�l!�	�����%u��V+)��pf�5z��8nB�g&n�nS���n���DK��z�+(�)�+B��Z��q��B��[�,m��2T3R�i+5����H�8`k��E������a�]�5v֦'!�����b\l=��_,�2^#��eZۇh�{l�>T|�ܫ��,I�]�m����Jr�d.�Xq�xwehwN�յ�vtYZq����J������蕗H�Z�'�
�6��;ٖ�O	я3������qP[������,�u��;/��qB���f�n�˓V�i�|skA����1WGJ`�V�{/3�(����Ξְ�t�@8��۝~�9��G=�)�	8�")��"�8�ge9K��V#m�8�܂�V��	3��"7Nt��4��g��"^݋k!�E��9�tAE�d����"۬H�Qq��Dm�C��qm�E�N��NNpm�^vs�qK��u�Q�tQȎp��BH��`J�RI݋˱��l�ӁÎBG� �t�����;��$����+p��$ q 9�dN�m��.�Jp=�C�=�Yl�*t��48Cl䍬����Mm�D�L�ye�8/4rf�A ��t#�a�r(r���I���^�B�)��r��� �;�NN��B���e���C�Q��,�j͵�b�ӎ�Ek����r��؜�tN;ۭ�c��#n�<��d�ΐ��kɳ�p�kq�i,���A��~ �
���� ~��w�ӹ��x�,G��e~D2�.&fkGf��]u����s���-�����+�Ɩ��1�@r�χӝ�<�~�U�<x���Ͱ ��D���F{�W^v+#�h=^!�k~�ڊ��ף_?>��>��"T 6���W���|
���A�u�������]����=����]�7WWB�:&n�������=�=�.�n>ӹʭ�"&���{�(+UxN��eg���B���� �H�]���D��Gr	_k|�_7��;���� t_2�_x�&!��|oڐ& &���a�"��{p;������Uol�F�x���H�%B����YDV�:ym>�}ɵ�Aڂ<a@�m�=ss���x+��:x���D_�o�<�*���zgmgpn�h�j���+�7�	��5~ԅ }w�.�e�#C/J�����OC��x���rf,&���Y�]�u;�^\�?;ʰFr�����Lʱ��`��;�z4�UC�3>�� ����p���?&+�e�A�E{���������!���И�o��)`�Ql�\��+)l�Vn1�!k�V���d,l.�~�~=	��oK[��:d/��l���H�l�F�oxX��p�;{�7j��|���@��ȶՑ�x�mwC<_>��O���5��;���셹�|�#z�S���� �@�5<`�5t���%|�t��m�[�ʳ�F�ٛ���ܷ�����__r��Km_�6�e)�N�1���B��"�u���ݴUgl�F�oz������=���o���(�N���Fs,���b"�V�_�e�x��f�Q⹍_ O^����E���C���@�F�"s�e�@�n�M�I��W|�
��=]�
���◕�����s��1dxݪ~��-����{n��*�l��2���\^�˸�wY�n��x����u,Ɓ,ڄ��h�5�YR�cucu��b����ٵI��q�劖�Ä��Ma��`:ԋ4��� �t��m*�D�̍�i�%�Nl��YY�J��ԉr�6M��iISYMCVYB��`�L�f#54s�#p�IVc��5F��K��a.
�`]����2��:(K`�e��a bɗK��6X�AJ�6�33(�u���@h�i��i��TM. K�	�f�3),���h[X8��롨�_]Z���&��6��:��m�����{y��s�Kr޸Cu�g�Cu�N�G���A5� ��_7� A�@��;�����?IAu�����^�|������ �Aۭ���9.啿/����R �f�A��|A-�x�k�c��}w�M����uO{�����7�"������D6���c��KaVߪ��^�@�����%����W.�6޸Cu����~��_��F�F�@�b��@����݋����q�K>f����}�;QU���5�{����R �t]�����U��?_����o�m���ַ0ĭ$��1)�l�, ʛu٘�\ݥD���f,�ؠ�_P������׈?�VsG<�uw��ys�
� �b�T�Y��@AolY�HKt�6��7H��m+��w�%�2�fn��發���U�=�~�6�MG`�hA7w���]vE	R�*�z�-@{P|�$��K���}p]��G-��ߨ�^����K}ޛ\ 7{�녖~�d�`��Y�kٰ_����_l���݋��~t�{�ʏ���|�*��wލ�5Y��|���RB�@����@��m{���q�1���=��#���[j�;�<�uw��ys�
�w�oP_���]
�cLt�����-� �� Co_�������޴��sޛ��n�S����r+���r��Km-�k�\:�9���/:Y`�P�Z�JZ�eG������8(l"�m�1���L����~��w(�"g��C�W�K}���ʪ��*c_khy�F�Y���j�ۢ��{�D̲�q�̻�oٴr��z�p�� �ڰwOk�uu������� �;t�m�x�P��X�K����w7A���I��MG�W�WPe��wR?Z����h�n���GM�c��Oz�Iy�bS���ص�6�ƍe[�phÛ̵^5��pK�)C-�|kn��,��r+ �;�@�� ��VCiz/{�����&��Ae�-�2�]o�wnu�W������W�r��6�N��#ݶ/�܂,�� ����m�e��n�bf��9��tO�v�W_����=ௐ ���-�23û���ݴ�3���(yA���*��v.B)m2�7`�u�z�ĭ4X�ՃR4�ڦ��;�H�!|Cn��������g��w�\0����_��,��/�@��mY���B��>�V����_!��/������U^|�Ⱦ������ �d Co5��+7�'�y}���|v5Ch/�,��͵��u�]��f�v�h�W�o������<B �;[��d�6L���_�Y�!�,_���׻��`�^m�p���nEdW��2?g���Gn>[FU�zC���k���C�l?
1�!�� v�5���nQ��rޚ[���rQ)a!o������O�`�U�,P��on� �_/�!�b�n����;_/�vl���*�>fd_k|�|� F��۱7Axӻ{�|_�"QJ줁]c2��r!�Q�K��%*ݐ\M
�*!P�ЪŦH��(@'�U�C�"�A-�������M�x+����s�<�ki���h2�"��o��/�V�ܬ�h���E�w��_.�[}�U�橮u�M�#���Ю��[Z*�G����ܐ?u� �݋��6���7.S�8<����d���fE���||�ؾ@�݋���-�@���-�猊|A� d��ڱ�vk�uw����|�;+�ۙ=���x4�� �_ Cn��t�!����ت�ڳ~B�
��7gmT������Ȭ��rY���`:���n�%<��'ē�)n� .����e�K	H��V^�Cr5o<��un릛�#��]�7r�]������w����}����j�8*��d]j6iR�U�kJ�Pc���(U�m��;Z���Yi�G0�3P�l�pM�Bif(͢8�ƫ�����meRTh�]y���BԆ	y��
Ʀ��4�W�3iY�����E�6ٗP*��գK�"vs,.���ܤ��]���!���P4n),��޹`��2�Y�f�]t���̥63D�4��p܏^sJ�l�14g�_>����2���Ä�n���(B��qj���54�k�&%[����a��DrŖ�@t�As�������fE����Wt�h��nV�M�ٔ�@�־n�e�A����9���^��h0:W���W���A�����Dr��_i�"�v,�.y�O����Ҷ�s?hc�գ�K���5�g7�Ϻ�l���j�^X���~�r+�Ŗ~_ڰCi	lg��<p�/�b��DL������UE����Α����휾�DB=�_�rY_Am����@��F�]��e����C�����{�}�9x�@�0�=�Ŗ�djϻɬ�u�r�Z�ʬ�X��4IltԌ�KGJ�KkCB�@���H��V�XXTQ�&��)����D*�����_.y����[��0�VІ{��{Q���;�.>q�f^�2�\q�RȮ���ΓzqGH��6'x�c]پ��o7��vߘ��ګ�����K��j�-xtV�S.m�Zú�
2P��=��:��"���7mW��2/������RL���RC��z�޻�����s������2�q� [h)vs���[��S���h�^|,^=KD��F�2�FebZff�t��ިr���2�#d�A~�m�uMmg�Mp�����V���ϼ��_=HK�_�6�$7A�B�uoǲk��5��]�|�v?R��3�}��~>��?��_Ŵ)�����������OL�b�2�Unƨb��B2���lE6�γ�m37��|���=���~�Ct�͵h�z�=]�<�h�^�|�e���iHPoe�g���"v��")ǯ���|N�*ڠ��Jg�^�ҩ��y���\��+ �;�_�l�Yج���3Y��#� �#�� �����y-��~�˰j���è^&B��z���=��r��x}�5���X�{+�wn�NԐ��w;���������\^�bh��]}�-���g��c�`�J@��6������Q5Ǡ�{�h ��#����{�����}�9z���A(w�M�)���}f�����-� ��"m|�=M�_���ۍ����:��+�?辱܂���[h��SھQ���l]�$�IPE_��ue�tA[�֧%nY�]�V����gS�r'�}��B���X��|�#���S�,���+Ҿs{�}/��M;۸��~�d GoX��m,��m}�x��fۡ��|P?=j�Vv�'���h�^�|�:a~�v,�W���wK�^(�#}�,:�N����~^�w�ۑ�+S6Gʷn��S�0��|���A|Yg�m���C=Ss/�}��̈́�<�ł� A�!}7�WN��{�t��|�w���|G�in�^Z3v��n�"G���ۘ
�E��N��u��j��4��:MEQ�^��R�gay\�����x�o
�F�Pc����\���������Cͻ��� Ye|A��h"�5������������g����尯�'L!��Yn��Bg�~�^%b�� \���u�\b���0R��ֆ�e�]2ipc;r��K����U�G=E����s,���ooo�Ʌ-<��>>G�VcNfx�~��f�e�3�b1��Й�XfQh�{��7�Cݤ?tޛ};�y��t�|��~>�_~1�D6��.�t��
����[��m�?6ֻv�|w��ܛÙ�o7�#�¾F����� ��"wbn[���k[�U�F�!9�������ۯy��x~6�}�e��f���Q�Y���@A�b�n��(;^�qm�߸�o�7'���n����!�G+�bs�֣9G�$�	'�$ I?�H@���̐��$�$�	'�H@��$�	'�$ I?�B���$ I?���$�`$�	'�H@�|��$�$�	'�	!I� �$��$�	'��$ I?�B���$ I?�B��IO�����)���<�Ϭ�0(���1��    �       P            *�      �     �U� ���@PD )J��
 
 (Q@@  ��B�)J�Q@ �
�(HT���RQ
)@
�R@�H�J�P����*���E�*�"��%�*D�U)UPP�"����  6�)"�Q �$	
#��(�wHE����[�B������si7n��ю�U`�� �*� � { �7`������݃�;� H u�UJXl�݃��hr 1	"��  9� ��)P�EUT)*�Cϰ��N&����`@ t �y!J� ��\�	�� 	� � ��K������z�Uz ( �&��A@���H

 |  ��݀&�QK �@}��  ���EJ� m� 6�:� 	 �(H��  zD)D��!UE)BQx -�@v��C� ��S�dj��24�@�r(���t w`9@�@		�  � �<�V:EG �G�7z��N!�Ҟ{ 7�G"�n����C��	R�#�  �!E!�TRH%!'� C� �`9U9�=)O�,��@���hw���ް�3�)V gA�Jw�ޚ�� P��   &���:(b�R��v��: n� tݞ����� ��{ ���2=�: ETJR�J(�   x��Q  ��(���� ���ɠ�{ 9� 9��Ep ��z����{ ��0h	{�E+����;���A@=�  �`��� �uV �͞��h�� t2 j�)Qpt7g U�Äj�U� < ���h�*3TdO�Ĕ�M  4�j�	J@  =��H�E   %?R�)��C@�@	55?ERE ��~�_������#2@{����ɢ,��ӷ��|��>�!!I¿?��$������$��HH@��$�	"H		�������w��y��6�&=,p��JN��kV1K���s>�w9^�ТN����].�R���n,Ӛq�\�Q�zx�ov�}u�S�$�3_Ay.a0�����'�����ݏ&��N�\fϧKV\؋������f$�ۊ&���[F�f�ܓ�S�l`Xx���w7�|��`]�� hw"܈�#�_}�w�iѻ�=5�Q�3C{Om�>O�r\�6�:sZڔ� |އ�9��st�����p(�ۃ���^�P�ۂ�Q@�9��E���D�x�'E�l	���|�a�P�(fY��4���+��s���@�}*���3�/NHgZ zYX6,V�9��3zt��t���:��;
� ���: ����1�A]�EE���6�-OG.�̸7��t�$���b�6d��1գ!;sn�-�k�����+�Yh��c=5U���GC*�#*p�N��oD7xmE�aQ6(Sŋ�o��2iyr��g- ��Wy��wq�_Y��Ųi�|���U�Q����L7�t��N�hGO����lي���§5.3���W7_onq��E`Âag�D1���6����3�n�B߶��w�/��P�`��T�
&p:n��BQ�f�K����Cy�����/w�	�g+����&Ԟ<'S�9*�뮄�\�1r�������#�R�6��y�4�ە�	�ɐ��O!k�a�1�C?/�1�Ju��;9oMꖼ�;9��ፘ�i�i�
�ܪuU;rt�(������V���$oKy%�"#㜇>G�k.�7t�����+C�c]����0�s_*��B����gm��צq�Sl�L1@�cb%T�"�������� wie��G�����*��׫;Cw,��1�΍H�����!�: �x�VQ+�}݃�~���}����D'vQ�o"*
��nr�@��ٸ����&uc��d΁���2R�|!7Z�=C��J�t����Hw�J�n�vU���[�^6w�Q�(; ȯk{wxߠ�m�]5�h����]��D��}�TrM��xA����d��v�v1]�q�%͇T����^�h�q�o��0��묖c���nj鲑i��W��ړ��Egb�㮲z=g�Q4R0c���]c9���[�)3��o˓��7	����`VOY{sH�KJ�;���]�r��:2��՗_`k8C
�ڇ5�M�5�b�u��z�.�IPۮYךO6v����8� ��Æ��r0.Egi��;5Κ��	�y2B�#$�)U.�֝*�����{E�ζ5�N	�U$��3�9�X(��Q�H���۷���8n.{6���x��^m3	�VM���C��ۗ�tO&Q� ��:�Gu��*��d���� >k�߻��ωݳ��v�;�� `�SX!��,�� Q��N�zk���܃�������GJ���,c{Z�%-����'�w�mѢi�e3y�]�hi�s����^ȁ�7��-��+�i�7��9����i[g*�r�H�G�U�58,Y:���
�c�H�;�|[�x���U��[���>�xki��a_7��P��j���x`�?�50��v�EG�\ywgU�G �|e�oS�]i�V�����S�Ή@�o�x���=���C׷�^q#����soj���P�6.���-���4b����r�Ï��u�ȍa��M��^^t����au/<r���zx�owm\�[��9�执;�S�s@ˆ���>��4�{�^�f����Y{�]�!0-9��X��/4\Dm³��:��6{�ێ���ٜuC/����ٚz᰾��ȵa���,2 $V�.�ۿ=;�ui�:�|��gn�Q
k;�A�r�������9��A�>��׵���seaA{��LXc��hKǤ|�V-H��rg{��]���N�������8���,q���cUr]�4���:��U��%�S�d����<;mm���7o-,�9$%%,Pmנ��G�Ga$�]Յq�LI�]��Փj2z�M�'r@�=x�o=���/9ubDՉ�V�Ǡ�`wtrof���x�!���qӻ�6��yh��U1��u<�q�wp*��yǞ��:
����dЄ�@�W	�:���<��gB�������} $�*|�j£ݤv�ɓ���E��{Gk+�V0�ĸD���ai����~���[}5μ1`S��m�);������\]p"�gq�5�`�B��Β}V)Pg�6�I���I��cŝ�^Ѽ���J���<}�mC�i�1��C���$�Rs�ph�'i`�A�Y�m|�X�n�4*��`*�ZR�͇I�T-zd�۔ٳʂD	�lW|�	��9Nt�7�,	�����q�� ���/w<+܃�wJ��D��G���Q`f�ȋԻ((NsA =ڂ�.;�a�qv#�VL �չ������w4A�Jwz��ubq��w\R�b�
�j���:D(��"H&�t��6�JJrC�Vf�J�D2��I0�=_Wf *�{n��k�T���q�\0b���	ɻ�Xw��z���d�t��aI���ʯ������(����<��${�۵��v���9�*�R�ÒAn���O����nn��q��-����yِv���`�O:�·eZw��ɯ���sDW\�W�2�@�\ŝڛ��3�Vj\ԛ�a� �^�)�r<��^�(�)��>)����ڨ���5]�؄�Y�=1!��Ŏ��8�wh�oQ
������y���5�k�f�j8q�e�
����t�#@ln�h�p��`/�=��N�;v0�R�+�	|2l'~qDhk~�o6�����;.-�݉�R���ӂ�@��a�U�I�ۓ���Q�	��W7\�J� ǅج�&ʚ��B#V���ȭ[��gRT��	����������I�P);Q�Nטڊ�ZgK&�bsX�D,�Z! ^^��@]�܇j&��4����Qv潰��a`jTl=�:P�ĸ�H9w��N�FwU�|.l}��a�����`��v��4��w��Ռ�7���}6�ׂ�s�v.]��ui�_K��������`�ᰝ�@p꣡K7�mˌ������Y.o>��T���0N��u�Q�da�=[1�	l�r�@��(�V�]� E��:�'Xujdg=I�֠m�!�/u�f�0��_ȊE�ot�v�@Pc}��3v���3�fo�fLb^�t|�,s��,� |��h���8�fY8u���*�5���zw�ld�(±|V�cpj���tY^���� Yo!'�b�hN/9nh�aĲ��Yp���H'EU����y˄�p� �K�`#�\�eM݅��,,����{��R<��_N�i�ݚ��#{�kz/uG��kK�ޗ%$�vgpë���)k��ʹ�ް�M�A7����aö���r��$m�_p�Ad�٧��{x��[�@K&�w�hn�s�%�S�
�,�e��sP�%H��,�9�(`	�v��	�����ҎI������Ox6��ж��ޭ���n �U7S��v�o.�V��ۡ&n�7��cΪ��:6�UQQ������u!3^V���'v�����9���Tp`����j�b=�`+��L��j�w����Ɯ��%owh��-52�t��T�NU�IK6Q���|��]�b�w7n]�yٷ�L��"�!uqp������syh���;����:%v� n_9�
ɸ Xx�X���	E����@���-�q`y�K9�P
�WQ$n�w�*[6�ӛO��H���Z��/��1��V+������UV��Z���`�O	�� ,G{\&o$f7���
�v���\��:�<
��}m��spܹ����Z�Ƴ_D��r]��t��<L�m	�r����ݯ�G5����i>�6�y��n����&xU&��;u�/�zcBU7�R�Fz�K���˸d=�WF��.����
���0�� �g@n�;���c���"���^2�8���^档)ؘ�5�����7�Ie��ć,]��&�KT���`���Y���,܋4�f>��!T-�����*'.�ed��\�۰�۸����d��S��4!�`��f1�U�XXv���ɱij����ZU���@X��7����'T��\����0�cq_�p�E�!�u�p��9�n4����h�`Z�iT�;�ÇK+�f���v΍��X��r���Q{�Ns;�Ԙ���dnk����;z�嗮3��bm�ÇeKd���`l��5�n�׻n��m��\�]�e4�	�Sۡ��w*�kp������M��i	��;k_$�	t0�y@ئ��~e���*�����2��Hm~�¦V�<�K8xn@�{d�r��+9��w�ׄ0^kvj����	�i[�Q���i L�����  �gK��6�����Ť�<
踽��:'�>޳4�r,�ob�:z��oL3r{ԈGJ�}�l�4Đ�Zx���ÓK�҈�������8w�n^hvф��]��d#_8RȘ��1��4b�7;t�T�d��dg(˪i��c1Q�Lu��avC_d!�G+�r�^|މܮ:2��Y�lF7�G����w�C��_�s|;q.�l�,�`p�}~��,�[.<�R\@�� n�)�z�nj������@���N�'V���������r|c͡�<��gp'�K��S�+�w�H˅�P��W[ݺ0��1���V���"�t$b1IY�
"6f�x�bk�n��{[ޙ�ɔ�D���9��oK �n�i�A��ۃLL9I���jNe���}�m25�.N���V<ב_��oF��e[�C4X�	Q%2�P�m&'��s��eʞ�kpÝ������]د�m����֍}�e�/�wMr"����ǖ^�р�)�R�a�"u�Br3i�Jr���C/���
7z���r6Wn-��bxZ��&MF^%����d;4ce�u��Ȃ�a�@M�s5m£ӛ�78S/�9�sWM�t���F��2vs��8 ò�[xL{����%%X��dk��[�7V�C����hȾ�)�;f��W�P���\�������F�R&e�Y��r�����Evm���EL��v���&;L�#��ϱ�DS�f��ݤ��rY:��чZ�kg�w ��n�}�j��9F�T��ֺl	�P����������E��M�׳a(�f�3{M��P��\u�:%���pq����e�Pˁgn@�7S���R�&�\P�C7����a=e)��^Oa	FȨ���$X�x��������ذ��D�x��m�M���H������Ì���zd���b:������Ln(�yȧ�Y�w7��;WU����ɫV��Z�Eo@ �����kt�]c�ҵP�r��i#��z��5朐gS�^� =�IA���-�n���ߊ�V�ҟ�)df�^����w�n�S.,�:0��`_�.���¶�	I���hzY�ȵ���nYvoR��q���h ��k=ף�șZ��c��V���&��o|s�øE�ώ��5���A�Cm9��6-�w6��tv�,�v�R����U)3��M;0`�YJVk��5�U�fL�dTwxS����{7��ջt5�R�:�]��{J���\͜��`yu�,ԕՋ~��b�8U���t���8u'o������"�)��ZVo"!��7��t�׈�'\���գ:�l�6蜊	B3s^�8'��+�s������Ǜu^%�u�T�a.+�OM��77 ��ѐ��Y�>�<2��9���8�d{�69[�������;y�7��pk�$V%���b3YB9f�<��� r�H��3z�8`w)��V.��;
�6a�4�^#��,�ʊ�L�͇e[����nj�tb���fss.�ru�o��e=�����1��\(�	ȵ6^�iY3��+�0��G[}���0N��4\:�2\��9ʮ�.�0W);p�����٧)u4L��N�4ʚ69,1,]]\����A�WWb�W*�g,�;5j��I��
b%�bR��uAE�ͪ��/ڻ &�îj�uE�vԦ<c��)݋��  v 毐ys�FV����g�@/p|�2�.ד�[�-�1��u<8k}F��%�7���v�δ�[�f�Ӄ���-�Y����n�ֵl��t@S_[�m�U�؞���wݸy	] #���������iƜs�ku����[ӛ��1+z1"�2qk/+:҂#�*G��X^LA�qǼk���5RM��0-��Y{��p�p=���e�	��2V��=G]��qk乨>����yr����Wn�齴����iiE�K�=�+�{ئ(�yR�R�d��aҫ�8�-�H{ܹ�T�;��Pz%ܵT콸�A;OtⳊ2r��Dd!#�ś��[4k���e�����J�s�� �=���W`$n��+��S����fl���H�kw�����e,һz�pŕge��ڢ�9����K��s`����fv��7���u�6dݤY����Hu� ����	 �Y(@P�E	H!$Y$� ��I"�)
E��
��I! 
� dAH@@�RB�, �)!�@�H��E�dXF@P��B
@H
E @R!� (I )	���� �E����"� ���$��I$"�,$XI �$�XH@���$$H)$�I�$��H,� �HE  ��� ��HH@ E	��,@X@"�"�$Ad$��"�H�	H�$�da!"�H
$P�AHEH(I"���	?�$���	!I�������׽�V������+�R���;���z�yǷ.J}��{]b��3U����YP���2��ب\<r�M8v�+Z>y��Dp�ޞq���cL!��-`)��}��������|6��1z�z�a��Z<IK;�Gw+�:3�wsay�5��躏.zG[�8��x��}w��<��X�G��o{wtS��Q�G���e�*q�k�mWW��hv�<'�k�C�N��/=���[�;�)z䧏(�7�]� �z���մa͜pL^���狇��?/%��/,яS��}R|�m"�ռ�U�� �a�JX��y�:p�>~�.���MI��ܼ�ēų*��}n?M����L�½��9�o���WM�nCi��>.��=3���ݓ������B����\��G����~���F ��<�a���;�پ��n��ˁ�év�c<E�s�2�*��,]��Ԧ�3��Km��V���'y7�o"*�=s�So��OY�\!2ꎙM��&�f�*US��=ڴ??{q�鼹\T]�u��{{���6y���1g�?.�Yu���/�>)�-�����e��4*�OC�&m�!�:ơ���<�#��-��=V��ɫ�ˢ�ތ��ISTlf:^�p&e��-ۓ��G�`�&!�	qP&��!=;V�FD�����7S�����t������)&�<%\�ąSSyǻ���ފ��N�Z�Ƚ����-�`�͏{F���/|�9q-�3`���K;ޞxrM�m4�v7};q����yt��b��(QɎo���i���ȅ�23��üox����CLŗ�k�>��1��Tb���`0����7i�}����^{�������[�D2O)Y�I0�v]��CBl��a=����c7�3�7�ؖG���m����OI'�����z�;��7��]�������x�;T��2'�i�D.(3[{q�y�,�gzo��: ��w=+$O>;v1��:"�Z�,;q�k9萍>�����+ �h�@i�y��P����� Vg�c9R~�Y�u��U�_�gv�y��@�wmc�9v$�AZ2,�SCKܝ*d`*��\t���ۭ���x�~���X4��:��Š��ӯ1�讛��-��tm�e�ya�Jجj"��ǚ�����bR5�V�LX��դ�
��]�����o�:s�dܻ���^ɇ#Q��,G��k�D�Y�T,��:�3T�Y����[��"�lo��J�C;ݻ�=_H���́�}Zk��3�
�f)ڹ��=�xv�hg7G/c��V��Q��i���3�8r���R���cO���Ŷ�a�ج:���ɲ�{��} �ۛЈ���b�ȷ36���U�V6���ojM]NN7��l��}�Eb{.Ov�x�eA��}ɻ�%�3�������˓r�J�{Z#�/�����қ-Dy���=�V�O.�Qn[2{��g���w�V�`��CD�"Z�8�����o���f½�q��/�ǸD�9S�?N�u����/c��|�>�޺�uXC���r�]�g�3�UXp��׷!æv����N�f�_l�v��������k���i��A��滧Gr���d-��HuO}�ٹT����2�'����u��,z٬�4\փ�b���[d�Ѥ<���ء���nx��1a�ך]C��½Ҋs��L���1���Ҽ=�a�����]�r鞜ޗU$H����~��I��`\�9�.1�Y<�R|:{I���&��f�r�d&�zRE0�9��+j`J�Km#��SR�ZHL��N�crxq����+�Ub��(�b���Ҵ&At�t���}	��D�ӕ �������{4���0_a���P�{����}�J�t`�v�i�4�
hb����ca��fr��A���p�<ME{�ɾ�p;�O1�b�B	��8M�e��KF�yF�{_{c��'�LW�&��^��c�.�V.^�P��sDO�J�WC��̫n��FX"�4,�sw��g/�������/W�q�r��6����/13�+��=��+��?��{{�.J��Jݖ�Wg��/-� ܂����D�#-8�Ոy�Qx��4V�����Г{�,��� .��g�0���B��z�}�uƾ�������|���8��F����7��B�(�nh� ���xh�ۇ�t��_Y#��t�zq�d0�mY<�y��p�;�q����&�r')7�&��
Z+0G~.{}ˏ�,�zn]���f׫<މ��eP:�e����:��5wT@b�L����S��4
�sqF�����þX����g^mn������w����^o���f��c�B�ӻ>�e��vuwG�E=n�ѧN��W��]ֵ�|���[�����ٹ决{���Dk��U�8�S��I̙{�%e�|\��oo�v� �ȇ�;`�c��S>�S�ݍ��T��R	�䳊zĽ���eؼ<�G�o��6B�����+G�k`#\b}c��re��y���z�K��]{���
�!��Y8���8����a=���4*�B�N��4W���=����	����7�5E�0BgQx-ɧ8�9���Q9D��N��SL�����OΧ���:��oz V�:����Ǿ�v��:��a�#��W�؏yWB��⑋����ۀ��^s��=a�VwyI�W1Vu�(q��v�~�fI�c=D��zmg��z�Q�L�;��px��'s�{\0�h����³���p��{����K� ه�����*�=�s�O)�.�K����i����k��7�W�a�>�*⾊/y��D�뻾�p{d�٫��ue�f�W���{5�rf�0�K�&��
g�4��&�!�6�d$vTጭa
i����R�'��6��wEk����H7}�0��f���y�����J`ޣ0�y�;7�컛+�繠ya�q[���˪��G�O���k/�@۶���k
%��V4����=�����1�-Y�s��h{ðI5#�����~ �,�i�s���{(~����*��{�JO��nWn�4%;�;��s��n篜�!��{�!zL�{�Q"6{�����\x�sF���AӪ��:�׾��ô��W��C �{ݮ��ղj��f�-�"��2�N��3��z=ȝt>���������D|7W`%�
{:w|V1�q]���ŭ�x,�ҶF���}N�Wn�M��o����;�u�dY��v�ǧ2�˘��hJɅ`������k�f+n�X�%���׾�}�����N�ִ��./M��JR�x�}�yn�5I���מo�{�#�{�7��&��k�2Y�� �	��p5��>z��r�1oW۷�:���y�w��^�|{�-��=>���l6u�E��cǸ��9d�����v��ʟ���5��c~[���v#�����x��ݝ���z&��M(I���<��-��rآ��0�fw�^:��{��XHՓ��}_�ɋ�}�k�R�g�NW��5���l��^3^z�7�\|�ME����?N����VN�vאljq���J��_v��ۨA�����I��@�װo�Y6w�%<��̣�NA�/D�j��]�4i�!a�+_��3��oN^���+ru���5�7��̙���I��7[�A��;�Ji&�����n�O����+��AyA�����B�+Ş���ƪ�ƚ(��[NoM�2���j�˳���S�Wp��\����wBͳ̋�:=��6��x��y��7|��۔�q�������w�� 7=�t���\YZ����[�y<N�|�#ڣ��:��}�'w|r=����]�{��kR�1��ܓ�C�s����5簊7���Q�!�:L�l�ʻ���ۺ��Ob�h���ݚ�.��W�˓�c�a�g�N���%���_z;T��/�������KEU[#��6q�o_2����`NR��9�e�@�j���Q�b{Ug��wJ�C�i��L��v�{���3� �X�W��G�%&�5��Nj���|}w�U{���7=�<W��"�Q��_�� �^��X��oS\���j�!��L���c��n��un��m�a0��94^�`��Q��{�ᾉa ���L�T*N�l[ͭt�6Dl	�4�Af�Զ���c���xvC�q]�RPs�����on-^)�{ ��<�7"ݜU��d��#Lit�%%�l�WcB���q�������64��#���4��w�T������U�����=��� ��G^���;�4���	�b���[㤴�h^�zo\[u�F����)�7۫��ĖNo�*���(U��)���� �����=�,ͣ"ʈqU��QSv�n�LU��f�+�8�L�T&�h�8.�Ѷ�F���o~���k��Hp	��}ˮ�OP�� �#�DE�??={�|�ן�w��|��S���BͲ��k�g�� ��s��S7p��a�A�	������ظx���f��(N�H;0O'�T�.�)����y�7tVx�s�
�m�t�ywЁ��k��<1i��;�J��o���yb��'j�˧=#�����Ue���
�Lħ5����)ިNP2L��T5z�On$�r=�Xai�3��N�c��)V��{�t-�}��=�N�f^K-В����Gm{BD�6�飢�p��Ӏ�S+676Ǝ��H�g3u�����H�P��q���?<.�3����wd�`���?v�EFTW��n�)2ur����v�gvb��������uB�k�]���8:A�X�W@�X_]�w��kl8��l��-9Ϻn����-ս���R�;��Dԅ;�+[M׼��������|&5����U�~�*=��G���MZv�t��7��F���B�HClT���WEƭ�y���ԑ=�����ݜ�����\a�ӂ�D���n詭��[Eȸx��ۇ�B�[��Kg{'<�܊��S�:���mn�{kC�H�
�6�������Ҷ<�+��j���H4�۽�'���5��g�W\��q����[lNT�B�ʹzز�˝��E�K,��#�Ih�[X��Y6�r�NX���FO3a�����S�9�W�v�_޹0�U4g��|�+��(w����M��[K$��[�t�-��J�Q��:��O��������:n��M'��1�к� ��E��w����^��_�����]��>��|lͼ�\�&�V%�ByE�ذ�a���)g�4nhނ��>N{o�ou����v^Kr����׮��I�b�� �3õM��,q/-S�mg5˨��6{x��G��M`[K��?c����@��Om�^\fP]�=1#{��RO{M>%�ܚ�C#e�}�`�a�-�z�Ґ��K�<�\i4��\}�i;�c�u[zS����)���N�q/����ȗ��K�h�N|夢mOF��8��/���+���d�O ֛���Y���0�M�,o;	��rF��ES�܊4�oKv�T^�L63����e�L�~/w�����wDv����c������W7$��8o�	 �*=|4��9e[���`��7�@Ay{D������I���{J�����gx1{|�v'���@Ϧ�iD��ʤ�p����wz�x/)�w��$������
��چ��f��:|a�N�����Q����JHo��wJ3D�rfk�Nix���2[8�֔���I��.^ �,o�������$$��o	֥9�6t#Eb�6����N�1c�R�c*7�G1r�7�` ����69��X\97��C�Gw=��������&��9�a�i�!w�<v�P�{j��WP������'�%l����ϓ��v���Ώv>S|ge9��թ`[2j|m^`����S�c.�k|�^i�ѓN����$�xrN�C8s��o���7Y�}v��pw��3;�8Io�*�y��2O^�2���'�dExs�	����?f��o�2N���]��9��0�_���=�Hr��ޚbZ�7��g������ֽZ�����"��+}�VX�>g���e�c�n�>ո&���z��f�y�����1ѩ�*Jcw2cFf��y3���rg?�[�rb�鈗�7���<��-nY�[�D�V��*��ϡҩîr��h:0��ݑ�j�`�"1��t��ޥ:�yE{�F��{����vi��NX�����s�9����~���=�ٻ��׮�6���&s��q�ұ ��s����q�@�d�{緮bę�5��wb�Č�s>Q�� �ɶ��MR���AS��潻�3��a_�x�w7�a,k^�wE��j.�>���Q�O�}4���3=}��g�j�e.M6�������>��b�g�����kH�^��7�Q�ݣ� �7`j2wfd�B=�bQ����wv�km3�m��TM�cp��E5�32��Q�-��|����~�N�FO�P�xC|yP��#����z��v-������d��f�����ol~���F�h�~c޾�)��M3`����ܻ�U]��r��S{��Z
t���ҷ���7�k���A��� [�3���TEC=6�&s�;�ܮ���R��ϻ˜�F3x���r矕���>t���v���ȣ.�*�ʷ(+�t�,-k��֔�oc����4%JL_KL�1Fl�21��gv�9�Z��g��gw��*t�)�f�{��2�����vT���x���������y��;���/u�v��z5lwյ��7�{M�L':ͨ�uTL�r�@�'?o{�ޝ'wi�����?q]A�b�)��M�{]��>(ָ��,��<7���7	"�"�mJ�J��4��.��L�mN�:�t��L�lgh����<̮+����<f��6ʔ	��mY��+Q����Dv�G�k����r�(�����3�yGk��vĤn)�!
-��ͫTԍ���[��a���ĞE|�I�|J��CJ�  -���.���\���d�R��`q�Wc6-�/D%՞�}Q2N�#����W\vM�Bг�Sb��=����gF�lI�ٴ-��@�&RGv�FOv.��U���fW��hF[.�4�2��SjK�t(� �ka\qM�e�á���f09"ńb�`�3ۆ�gv�.xnPB�\Wj��ۮ���u����u�P:��yZ@����ε��6�Evre\�
���1e�V�qf��<T��jιP㞇�泛����ۏFq2)>Crg`Z��^��u��Z�4��)��H�17[-��gh�y��J�t���^0t֗�v��%48�%�n�tØQ�]1-�2*�=���,lr�D���\�Ǘ�{u�e��t\�v���(�h�Y-�N+�.	8��n�x�O��tn.�l8�W.M`^�.]�7d���R"���qζ'�� ����@�V�f�`�Q5c7ۮ����g��mm�^��.W[�ڰ���ۋG�,�%Xz��*�w"df�Յ�K,��ɣc.�[��A31Y���4!5Ƽ�d��u�3�Mu��b��t��u6�e���O-A�T�cz��f�j\�l�8�	�lx�����\n�C�A�ܖe���M�6q��-���,������[�ڸ�$���0�c'c�t��3�킸��m�"Vh�4��#af��c�Zٵ���q"]i�^#a��;]n�A���Awg�)�9f����� ˷ؓg����Oo���gl��\�0Bv���̪F'���I�gnrj�����z��>�pI�.�&n�!/0�6��XM�m/Wm\I�%����i��/jR�w&�� �<b���^^m�p��Z�(���ݮv�d]WR�"��Ѩ��R� -��ZLf�5���eRbΐ���9i�k��94�7����7/�ٯIõ^p�LC9�(��rVd��mƚg�F�4"K
jm�"Զk����N�2��3��uκ8g�C�9��Szgrc��B��t�v�RVQm�) `moKH-no-ƭN�b8Co=<<P�k,50kMh��(�%���'Rg�CY�Q�v-4�S�f��wm�t�j��t��ZT�F0��������f��ɶt4Q�\�U�͖i��Y���(���S6�q2�Kr�T1��N�r��왭���b����-D!,��FɱbbkpA��@t�l�^�#I��i�)B򙴸�4dn:O)�[ڼ(�[�w��;0{q@�m�)�L��0�X�XDn�32��<���tm\�i�5KABfh�t��vMn��M��cmG/+�k:�l�l� �*Z��1����s֞|k<� �a.nz��aGj���P@�`ܮy�8lō�)�"Bf�qb6���\�<j��ޭ����B��L-(I�[�1��c���&�bܡ	ms٣3yй d��n÷7�u��A�%�m.�F�(�I�+�cd$�ͺ��/�� N�����gO�y��Dmg"E�X�#��\�G.��cXm���lL�m5(%����(de�[	�IR��6�=kO�6�ŉ.6���\�p��:<NS���n�\��˂1(�)*kZ�Ī�n���8�\n�yѹ���=��ә��h�m�p#*Y��.�[,I��+�	v,J�:m-��Ѓ�giu�.tY�pK������*��M��T�u�����8�npzz<�%AV�OLD�a��9��[g�/G<�n]�.�!И��m�<����2����s�
m�-{��b�n;`��ڌ�%�Ls��u��U&����� bɯ&T��.`0t.i���z�r��ݜ�K��K���n{���b�'�8Ex�G]m��Sma8Gk�q�\B�Mc���	P��v�a�6x�)Y�\H�ﾭ�[[	�{�S��n�kЩ�k��d���;��.;d��nx�y�:���o�|�n�J��6ȳUY��]�͐�$W7�6i�R2�i����ƕ�VQ�:P�������٦ 4����k�s%q�@8�yR�;ԩ��t@&:�>r�<��|0��syr�V�ڏ�]�>C���k��s�a�d�nb��T�Drp>���3c0L<fh5حԉv�s��Eq�
GC0�n��c&��9H@MÒ�VշM�C}��<n��UGK�d�\=����~<�7e�!���U�cGel�C�mK�ٻX�r�n��ϥJ��5�O]�s�4��l�3�nmN�: �xrغ ŸajH�iK"�[I-Q��x����L=�;z��v!�#ی2�v[�n$�ʹCn�፦:�k�z{������f����P�庰U�"����-�J�n�A�ѐz����X��T����J�B��(k���)X����;�a��n0wi��K&P�t���e��i�D�O�sV�]�sx�!��d�C��V�aw]�bT8FTg���xHZ�MV�ԃ�],]P`�c4e-�=&��w���s)Eųa$֙�]���0���Ń��<�A�㴱sc]Dd׸���و��s�n�f���{�q�	�m�W��2��ioD�>.�W5�ӻb��E���C1U������Ri�`\��.�6�s"ͬΆҎĭ�:� e�F�޳DeE
�(����v]��6^ܞf�4S��!vt��u��;��&��u��̽�L\u0讹�*�*�C��,�������%�Mq�m�X��;�������K,��흭�	GR�XۛR&j�ݱ�����3�����m���;4/q���%-܃ps�]ٴ7l�9�i�mȃ�;N�-���	��1��c�Ã�F�������bfŌ�mn˜J�R7�X��؃4�7h0��G$�b��"o%����]fs�a n�q��2q�G�Y������]fC\�� ]lR��;��u����n�]����ΰ��d�d���������ue��r�A��ӓ����9C�\ݍ����"���k����	36M �3\����k̶�q*l��mL�-A����F��b�R��Z�c2�fV����(c���L�I�3�O���nd�^�\Hz��9����[
7E#Z���ێ���mt��73˹zq��!'m��;�[B*��u��ܮ����m]*#�����y$��ђ˹�K�u����l���λ:��$k���.ͩ���Xs1�͢�f�2���\LiE�yԱ�E�.h�odY+������^֐��1[���B.,�
��k�cm؈q�X�il;k�b^0���e�Җ\���on��=+�33l�m�Gn�źY#g!Cd4��[�:PƎi��)
�C�ẕ�It�)�Z��x�8W�Q.qtC��^G���p�qdr�s��q��n�>��S��	���p[*V�\�2U��$�;tl8W�$��=�8χ2�����9�u�.�U�{��q�|�����Cg[����7c��ۅ���f���a��KdDo6&0]c�c�ՏPt F7j�rkvc`�ȱ�����K	e6%��^uã�oY���x*U;9�7'�	��M�v�Ǫ�"�4��q�g�;��ԓKt��vi�H4��lK0됂V��\Miq!�z	`U�R*�cpl:��;Ao\�QP�ä�ə^lj�y�.�7<���	B8����e�d���D\��������T,2D��(�V�Ŏt4�y:Uq��p���M�A���7Zj2�e;*%�ưZvs�YsdX�ó6�1���uu�ttL�!�e�V\��ġq��l��lsy��sa�5�K�A��ĩʸlt�GLBP��5����]kA9��s"qq��͝�ݽ7B�m>)��e�ͦH:P�Y�ZA�v�D��<��8��3����f�kU��́@ٻG� ��H����κxdU��4�]j72��6# VV6�؍m,|XA��͔��R!&��պ8��3T��m�)�\��[v�e�`��p��D̴Xˡ%��S31����D��],<T<���[jo.�f�rF)�͘kG�UrMe+R�]g�0����ٍ��4��ӏ9㇎.�<VHݹ�$
�|qϭ�S�C��`�˹��ns������F����6:k-Ka��kw\kn2��4��o9��]&M!q�)��6D�P^y�K�b��Vn� p�P�k8�C��=g���,:������n�y��n�s�ћ��O9��ñGF����9��L��gW>����"�\�&t�Z��$2兲������+����-%����n��0y5��<s����٫��.�e���cT9�$e��kmnu+fUVeH�&���{_s�F�e!�:�#�2�-j	��ZB��C5�.�/p\�o\�[�s�v<*�i�j����Լ�w/*��Ҙ�,([.�E+M:�ņfm��m�
��rSm6;hu��PG&�Q��7����t�M �����%�%1omv\�u��mזX�j���]F��˒�LL�,\�`J#�̃pZ$vwe��`�9.�f�5.���!�57\<]��^��M�m�4���v
�=g�o:�Y4]R����ʁ3�����I�+�����+�M�!{X	��`ۮ����b�c�f�8#�r݅�a�����+6MP����
�M@c4ֶ1e��L;aa+B�Z���Sl���ds��s���YZE��x��")��Ap�����6����^y���*�rNC�m��t��s��$��vR�<֓��8��d#�vX�gvA����,��.9�8������v�93!s�A@�'vX ���s�
K�v`�!�B�r'KI�ȥf�;�M��u������nӎ-��Ȉ;�ݓ���[gM�E"�� &��%�������%+c3��]�B$�ZE�p��&h�"IGme�9G�9�J�ӄ�;l�!�%�Ns����ޯ�߆�BM]bCn��`N	�m�@eM5��@fYm��H�zfG��u���en��YI�1�Sv�tev�y]��Y�Ǧ]�R�O��8�5H��p�%�`:��F��LB'	�v��j2kM˅�앶��i
:����v:A뀵��xF�͉��EMi�p�i�[�.�t�`Ӽρ��v�r�,/"w:��&x���6�lQ�$�
fS��8����hK4,��:�����Z_*��{Y.N�Jg[�tݞ�ϔ`h�G}��VM����Vg��8���r����Y`�-���^ef.�o=�@��h�6.���Xt�b��d�b�i̵q�����li�a^a��V��ǥ�ǰr�m��r��-1lf�%bL�%�F�-i�^�q�K�-�U�`ɣw2��H�ݵ!��f�We�IGL�)�أ&�T)l1#�JWiQ�:�փ�N��U���An�W8,�¦��s��6-ֺ$G��^��f����,�\��\�62�8�� �s�>#��;�����=XG�.V��iv���hPɶ0i|»t�8n�/63j7\͸���q>}qvJ����E@ol���=rZ��NG�4��y-Fx��d�����4�����r�Zb\.�9~�{u���V����V�!�^ö�2��D��Xٹp�-����k4&��`��pB�J9u���cI�����u���
m��`MK2��5b��X���&]R(YLq[�t�=hF�cC�Lpr��{&�ɱ������'��v�j�zOE81�y�(|��2������kn.���%a0֒��]4¹,fir�Q�v�I�GM���&����&k/v�n��q�th��p�V�ZNN���y7<��V��P=�(�v�z :��1q<M��g��Y`�du�l�8�.�8��R���'F�T�Ke�����;���z��7RP�v,��v����r��L��s�6������Ɍc�Ws�ly�!ܜl�'�(nN���ݰ����q���]ؘ1p޷t�!t�.�R�"��8˗aW��s��q��˸vAv��G�{g�98�l�xs�/v=���]��߿��O�p�2Ƅ���ƶЬa��]�M�H�&��k��,ce��7��<�|��w�p=�/%�P�z[��*6zW\Ue�GM�/��/��m�3^O�Y�-�=�=;��/��U�ݝ���{���̎#��
껺��+�{�231{وN\V�f�o��8d;����9��d�̮W�/�1N��@��mb+A�9��6��w���=�˚&f�t��@<����d�XҚ��n�b_Uf��7����=���ֻ}G��kr����v,��Ѥ]sA�z�-��y�\��s���<�f�[��E��ĩ2�]@Ό�^̈���m�����y^WS��0���r���d�2�bb!K��Ŗ�:s-DT�!M)[��i�3.g�ވR�n��<t��M��yn%�B�l>�z�bZ�����A6�e��{so�'x����qޞ�/c3*:/z�I�ޥj=]���dff�ҡ�k�E�n������q.�^�����yZs-?[V*�/O�����s���̆����0;�tx	�h�Wi1��!Q7t*�>��31��|��d��u���$���[z�p��{3��*�i��^Ҏ ��(��Enǈ�q���:Ȏ����Yd��z�b����]�>��>���@̏fb�i�Gfq7/!=���0�8^{���Y|m9mY��M�bNn��c)�yk{{D=�����k��O4/#1��=�����^ޏfb�d��M�_h�C��f�/�\c�fOC��x�{�	��,ҳ�<N��9y�od�I|f���zo��e��\>9}��eN��t����E����o�<m��M���7��{�=W̌�An�>���K�s���s����i���C+:s1��fB9Vo5�h�3"c:%�t��˝=<��_�Jm?e�EJzok�C�"�{/[v$�	�6�#lj�ff�ű���][���) �P�b�/#��{2<3 �f�c'xݺ{��޾ҷ`FH��}�ّ����WGPۂF�Q*scۘ�O����
����`������%��<�wSN��f�;�G�#3�c�xsz�t�\me�;�u�����ooh��r����f!�w���dq�>u�>�fٻ����Om��OE�a�l�*�wٝu��;���ɹ�����a�Q���B�r3��PZ��@'uӲ/���ׇ��e�y� ����w@9wRj�ō��ë�l�3dfp�Xi��	=�^]�O�sK�{S�{���ff)��,���>��7���{���V�E[t�
�7�2Zxۖ��%��s����n"�-��
��{%9��ןZ{߫�K�����soh���J���݇�/#�33(f@:/	�1�~��� �oa����Y��	�����U6w'F]�����d{٘�:^���
FVs᝝��yV�=�n=x�d{2f*4�:�߲��^̏wuwgl>(`��ʎ\�Q�xOD2�* wF����d��fu�蛮��\��;/�hjN�q�y{n+��s3 �:�"+9FiH:�:j[EûT�q͡ ���o�U�Kܷ���i���f�mVT��7�R=e��"6$>������d�����+"�$TO<��^�"#q��d�9���ol�
�	v&��2f����#y��S����J��t�Hݷ������7��&�=���P�� ��c�y��лf��bU%�@)�C]�d�	3q�X܍NX�&2g�[t{Q������ۛk��9S�d(>=�;�s`�N�v{\���g�	Ҙ�:�RF�8ކ���U�֪�hjk/?����i1�&��2�\�L�����)˳aC�ʻ��yPDPW��y{�3#٘�M}_h���V�=�9�����R+�i�j��O߉�Vusv��KHt�����ãl>(`�w�G��Zm{�[�H}�fC����M�{2<3(@js7���U�܎)�=�v������_[^[n��p>�<�����9�6�	���{/�Sn1�X�𽍹{X�oL��p����j����j���RxN����;.፰�Acsw*x.k2d�9�Md٫�sȧKY`�:qf��8�C6!&��l�2ٴ��i���:M6�R�3��&��O~^��efC�oZ-OA|7o/m�h�G��]>�+Ź�٘�3Ϯ�04�	��m������c�m�����wU��z��Q���J[;��9�=�Hq�17��[(>���J����oe�*i�=��׷��p�)%�ӱ��^�d�C1ۗ�g��\�e��6��r����fFd{33+�Jf�v���u�˲34�=rquC\7o+m�p��n��p����ۦ��kב����3#1qΙګ�yR�c;r���kՉ�[�/,��%V
�����;�3��P:��6�Z�--긔\�Z��+Ӭ��nN��A�J��:�������wv�C�I����^�=�����{��W֜�sٽ���&���5�����������	�6fvܥ���T"�c6�q}m���!�w�.�_�w�7�{|��w��r�����=�vh�Yc�Cٻ������'W�=�}1��v�S=����ю�s�`��[�*s�o���)��Sњ����̗�b�[�/�d�^7w�s�b�I�[�z�d���wM�뽪�'��O
�ٞ3<5��d�^�پSr�N�7��45��pݬ��ޞ�����ɼ. �e�Y�\d9�öf���n��\�w�t�]��h���HD�wL����sc&н�����N����n��9�?u�����On���i����%��S�� ��q�ݛ;d��R��̌˽3�y=�J�X�>��M���+'��[�kV�cc���;Y[N+����ۯ��]������v mƮ��{;���ݫ�[�cF�D�h0����Qslwp��0L�Vn��c�:�*�nhJH�p�Ö��؊1u�E�ݬ���jn�����\i��_5�c���p��7�og;Wu�T'{�6(v�8-�ڥ��1���z��'g*W)�<�D"������J��=��c�3Bƃ�� ��t�&d�g��;����6�y��|y�s#��em8�1����q��6�n<d�ei6+�T�S}�|��Wh���f��wj���1��F-��[*��כ�m��x����YPbzyg<��h�mWz{P�ۯ6�l�/aߦ^ϧu{M��ǘ���k+i�w����}�@��l�M�m�6�l�;Yi`��R]U�uo`2��wn��n �i��b�Y�չ����J�{(��� i�Pk6�S:���s-y\������L�8�V�$�5�n�՜�J�I��M'�\�I�|Ξk������p�����)���Y��!B̳g�!
W8�hM����v�a��!t&�ٵ��K�GCA��s��6k�Lvݝ�WC�^��k� ��D���:�;a��y�G�ʰè[cx.������{0@m�]t2�D���hg1�P�[+x���|�ac ��C0�5������3ɓ��\�Z�%΅vњ�o�g��]G�:��.xi+u����g<�d2L+��fa�fi[.YU?x^���m��Cawvn��3���j�tSV�jݬm���n0f�]�L!;��7Ϗ0�ndv��ۦ��������vMf�ܮ̸���sSm��np�@�Ƹ�؝[oj�eo`2��wn�����6�m�R�=��+kf�]=7��w�^任7Tu��p^<ڮ��}�w�����v����6�nz-2{T��p6�9� ng-���M_OZ6<�^m�T�+`AW��%)L�PL@��n^ő��vi�\�.�ֵIc�HU��Rc��~���^��q��K~��݂ae�=�葜سĺ-�0���m��m�lno�ey��4���B%�7S}�v)�b��T��`�s�6j�{��G���6,Sf2q�紨�
{�Nu���� ��E�Wxgj�wfꎱ:NǛUޞ��7�*.7��l�7ӱ�k�m��p�;wT�O�`<�ٝ������3[tm��|q��7%`ڵ���ޮ]�&^S۰o���/j�Gc
���S�@=��@6��nX`���f�De��=��W`�9���p��i�;��Li�x'�L"f���b\C��e��0�ia�M�1(�݉f�Ix�e�1�{�u���`75������{I����Z�\�����k��MǃmD��Mt�R�vN�r��z6{�L*̧�@�[�m���jf�������m�Cͽ���^>��n�V��W3$���������4�1��3�9��KLn�ֽ�A��G̨�t� �b��C��,�(�aMsT�"زmB�\[�	l���tɑ5;aTl����m`j�uT��<����DN�v�P���k�x��=ۯ��V#e�����y���\�h�]Vv��{�[�X�@�}��Rbx]��|���v�r��������Νy/��=A>jrݴ'qD�B�n[�+뚍Xb�Ѝ�ńv{r��,#�o�����(�z���l���CsF��^�,��c��F4U���\S�:��Cz\�F���&I���=��rA���@�����pxWT�6"���	�0q%d�Fvu޼�C�p��f��ü��Y[kl��1y��Yt���{K\���d ��'�xw�t�g����]�bu�~����;��m������m���hj�6v}���w0v���w��>�ܵ�Ĥ N &��ζvn'�ƞ�е�s���\�"$����v��}~�]�������u�Jyl����_"=�Rs��W�z�� �^����~-���g{���~գ{(Ƞ�:������mOϳ�ѣ�0Ɯ��U�������g�6��7�q�Z��pg�3y��Og�>i�����ك����mej 2�"��}~���r�Uu�W��EI�M��#�oyQ�~�:�����0މ���p��ld��\ʂ/n�'�r�'��H$�A 	��6��-�%�M��9�Ч(
۲p���"@IIӖu�9��gZF��:N�Gq�3�s� �Z8�;K�D��f�m���k(ขSf܂�DP�n��;+;���M�����ef��(�$��٭�mݶΆn�,����'E�mƓL"�"3���m��XۦҐv��eY�kY��9m�E6k@Qqdtsj;,�-�tV6���m3ggY�4V��v�kvvi�wn֛V�Ήp%Cm�Y�jJN�� �IȎl[�G�<�ս�+�N��X�j�_&�t�^�8-w����Fv'��nk�͘y�+e�'s�Mr�12���Ѧ�^-z� �A���p.��S�(;�(��-��UfS۠o����~m�D��s����ƹ�U�t�L�]G7-˨(0T7]m���ҘP

e��)+��j׳�th]=ٺ`�9���y=�*�t
����,���^n=�bt����ٜ�-���5���o;el���x	�^��������x��z۶���{6+��\:��N��U�On��gm�6׃m��ۻ��W�tnj��]ۚ`�9��w��r=dB<���2z'��B=�9�ty���u<�|ws{�B�J��뱐"�c�;d#(a8��FD^�,v�_�o���=s_<���k��m�����^㿫ِ�x ;�I�t�Zu�f���\#z�z&<��0��(���z:n���s�9*#ų3*],l.o,�5��Oo/�x7m�[��WP�*�V�и��2��œ�3@N�m � �@6ש<55�mz���.���.�Zr�c�7�]���%9�W���B{�ހ�A����ܸUVf�M�ݙ���{V즯���� 6�m��T&�E���:�����_]C��y[�Bㅸ�)f���9�T!�lvb�����n<ۚ��E�f������;i�Qo\�yv�4�޽�5�tH5Ȏ�������~��ֹ��`>���|o5��}����t�'��|���{��,~��^��a]�8���h�=��?�O߶����t�w}'�	���3C�=�@!��5��K@G�6�J�@ݘ�#��h��UwC�ha�S.lۮ(�
�b�]ɐ�=�ۢ���,!̨�u������5IvF�� �ɛ7j�t5�;�S�	����*X����R-�ܤ)I��z9W�6=���9Ӹ�t�ȅJ�!p��VYeCt'l��ܓ����d
��6��+f�=���4�����[e�	�-���v)j��.��K�6��.��̃u��_��޿}�݆����r�u�)��X��z���W6]w��i��躨��we=�������U<�ۡq��ƃo!4N81�n���y[^�7��ߤ���q=�R�fU�h���)E�s|�/<m��ho�0��*}űSKß/75�r�u��+u,��=j�QyUׂ�-ނ��mzޠ�x6��mx6�5i���t����웶;���{/n��{���n�Ɍ�R�˶�%&RRaN##5̼�W	�^��t�S��Ws��5߳����6�6֮�}�c�V��i�W�Ue����3wmxob����m����3�� �CB/Ί)��}��+��>?�a(˲ˬv�,Y�å��ѝ\��(�yj���g<5�XO�v��V���Pݓ�6�m�T��=��]��s:��Ш��fV�YSޞ���m��N`t���^y����l�SQ��G]=�݃\ރ3Oe�и�����6����Q1Jr{���^����{;F�`�9W)�W�]�8��t�˛�������h7���.������Ѽ�̖�Fwk)n���z׳a��m��S4:!䊾��5�#u����*`�9-�w:0��^�	�{d��<�*L�_����{�g/7ʹ����z{	�����\p���q9Q�Ƿ�������nh6�8��֣�a��_tr��;i˹OZ���@n5��9�bw�̫C����m��n��(X���3 1r���w��H��Q��[���z���D�䰐pVu�pf�5;2\����j&6^ܽ�yuV�qt65�7w��xx��y<��wk)n�����3a��m��N�ț���:��k\6�z��oud�ݗ�B��@�� ]�FM�.��A�����6�X�����b�z���*�=j�.�7n<ۺ�3\z���,���m�4%���9�<s�D�z�b��4���&�DL+�q��M�������f3{YKu,U=;���Y5L���z�m��6�t����`{3S����YMn���k�[�M�sb���C��1�mx^5����lfMV�ȚȰe�>�霹��Wڷu��@6Ј3/��;uq vj}�����ޝFc�k2�ab�z�M��!P���z":�K�ˬ��`tb�.w��X.s,_z��x��b#f�N�w��V	�:��L���#vlܙ�{������[y�&�6�m����ҵћ������n�+��s[B�+��^m��<{f�e��:�����=x�͟le�L��)¸��k��ݝ{c7�Nx	�������^�m��mr������\��+�s��p�6��ys�6�vq�������V�9�7���B�ݻ�gv*�'�{6n4�{�[1MN�' =���tf�e��wuU�Y��T�8���*ku��������m�l�Y�����ݠkWM�h��;�r�q]�P�)☩��;V3#ۭ6��q��m��b�'*]M�/�r�n�'{w��,U�z�͏6��{�t�67���ڹ�"v��Moyx7��p��t$4�lO��;9Q��'Vɥ�forc���p�7��f�wUf�_]>IH�[�i�K�< ��I�# ̩(Ľ�.뭀Eۜ/2�.Ձ�h195�,�36�h�1p;�y.-�Q��va��WHm[u/���n�lϤ;tF5ی�FZ^�r`��8��x��ӷ���ɽ���>Lu�a3,.�	\�����7�*�y|��vv�!���ls1é�Ʋ��n�a�����6��Ծ-�7me����s���;;4�������Y��V��D%C2��	�Qk�,޺�a� �c�͹9��͠/��y���wa}іT�띻2GZ̚}W]S{�#u�7f��6�mܨ�J4*���-ж׵t�����'-�͊��^���޵�b/�_X�<�M�|��<�����P8E��O����D��,U�ֆl6׃m7{a�S�v$.��.m��m��k��o\��W�z&2�
���w�L���ٸ��۠�C�Ǜk�EfY��W���	�w����)fĭ|�^nk���vū�<�\b�9��1���<V���\�d��4��L�Z�YyHa(�e?VG��/6׃b�rz�;��Wi�Mg	���Oq�m7܂�h}�_@�r��uy߭/��VTߠ�ȟ�n�)�Ç�o!&D�k�Z�)hP�
�WoaE��7��Ū�7U��'k������^/���� ������b���ڻ|'�[h6�T��ѵz.��Q'ܻn������؃P�T��M6"^��s�6{��nj������;5���^�y���6���B���bgvepzת�\a�X� 6�y��m71�i�B��҇)�x�xص[y�Wb�	�i�����/C�7�����X3�t�jv�p-YI�L�Q�*�4hD���ID"Ȟ������hj]{�"w�pN9śT�;�>�ζ��������*���1��#P�����־�T{�lL�\u�c�6��;#��W�^����Ǜu���,ɍ�bA9�W�+��a"�'�<eڻ�_����%��8&^k������=��=V-U��2��F��Cwo�ӪXTr�]l���=��
9�oW+w��k,R��z/�my�m�sk��PO%�D�/��hUս�6���qf��}O �u���O;B\{;�m�7m�y�șqj�Py���#��T��X�����m�(d1�x�W92��.f��B�<\�N�pZl(�n�:8m�<E�	:<�f�O�O�(-�N���9�ʹ���۱�ػ�׮�LeT���YXN���-�m��W�e��}��k���j�����X�s�6=�ۚ�}6	��T�P�)�@f��݀�]����ʻ]+���Hy�3��+�WZ�8�m�6�z�lSc��5���m��{{v9w���	��Z`��w2���e9�*��;��x%½���,�4˷��nQKb̔�s:c2:3`A͸�ݶl�$t��[�{�<<<�����y��mx7��B�˳���\��+_��N9ś��{s[�ڑyJ\ǻV-$kDɥL\h�ųW`õ��69��
�Z���`�&�����A�񽷹ʪ�gdl��X���Y���{��2�,�=���� ia�E�n�d���w8���q�໼��hLp����jrovƖ\Y:\*��� �y��q���-P�J���5Wb����۹���^m���!MHq�5�����7+��)����weVO[kQ�QR'�qগ����my�ocȻX袶ixdl�>��pU�c�l�p��my�����y��3d�fg]&�"X���P�����v'Ͱ�L�v�_hGz���wޤ�-q��k��� {y3��1Q�=������n ��V���鴿MΤ�^�^z��M���ZC*�uLc;�c�dH�ڟb,��w�{DF��n2"S�}�=Ps	$�*�����ͼB3'^9�w��]^뺬�6�����4�ӓؗ/o�2	E1
��n��F"n��@9��ޝ<�zs�4�s��!��˃'{����<w�x�޼���^ٱE8�*a9�c7����/v�/j4>u�ۈ��̵��jGf{$�]�9X�1I9��wԛ�-�J��b�@:43m0&恈ìjS�i�`r�>
�Oy�`>�9�B��k���z��0f��<wo����{�����#+b���n �j�A�����R��u駵P��M��U!��:�ga ������' f��Q�E�g�;v.7��zGJ5���\��y��#��;���ze�<g�fN�y�h͇�>��LޣFŞ=��l�=1��}9�n��O���<3�*�!�XK��'��9\���+��'��3��b�(\�����)�h>�A��⺺�uQ �b@m�1.M�mJfӚ����+��t �.F�f�!�؜2Έ9"B�H~���Tdw�KHȟO/{��!���׺����
�����u�w��i��u��}���_����>YWM��:B��F�x�T�e��yt�難�[Ơ�
��7B�N�kZ�ԕ�`��R��3�Y���b@���F�_Ԡ�P��m��L'I�����̳h�!��hI��Օ�M:�kB�ֶN��gM��+dn���ٚ�96�Y��$NJ9`�NYi2��dIXYkj���03l���k6�&ʋm�۰��%͌ʹM�,�-:vh��n�B�V۳L�;:6����m,��-�m�f�΋�ŝGSd�����bV��۶�,�)"���.�2+(�+3[m�����u�l��ݵ��",;:3lFRv�qY�gv�v��ᖚ��qRFw;F��۬���n��9���ڳ;���2m��B�$!�	����KuŢF�M�,؂B��[K6�d�넹ZN۷��h�`����t.�mc-��J^ �]	#�+-�����E.n�:�X�@��D͕ĸ&�`�C�G5+��q����l���cO<��k�ф1M�V�z�n6І:uY-��P��g-����tR��
�G�����uA1�w��8؞CNg�&xHy�t�m%x���>�)��l�vcnnC��V����.�v�7I��xY�s.INGf5z�\��<�r�u�㇊�7�{pl�K��RR���P�
7�ӻz�Z�]�Bsl�0/R^%�,:��Alqi�v�9���Z얮,Q��a�Q�DwYyZ�+�LQ6��%�X��"��Okn�q�`��p�Pf(����5�����И]\�2�D"��s&�T�5���z7i�����zap�إ��Uӯ�3
6͖d�3�@�Z�3�c0���V�6�D\	�]&Lز{��[Kf%2ҥ�-J��t��c3���.�Z�u[t+���.ZTЌ�kyX�!�<��Й��sr&��rSX�&u��]ajЖ�$�m��5�GG0��T�j�N�t�jT��;��u��Ј�+�
�%!�N�[X�xB5�邷m�vi.e7m�K�"L��)�q،�b�ڄ�iY�q�i+{f�|l��/<��)�p��ٻg��xJcm�s���n�NnR�;���ٺە3x�M��e�2V�@6�#+�q�>]g�3� )c�=��gE���#�6v������l��I����6�c�E��ꔘ�+�0�M��{u�Q��:�糋{s`&#��j9JK6i�N�Ͳ�-Ɏ:�A�܆��HT��Ѓ��b�4�ak�hP�Ӻ�90(/]I�- �j��\������.$�n��9�\qj2�L0��je���. �0F� =����1٪��-u\�)͓=fCb�W��p#��yѺ(�'-���Һ���Ӷ�5a���q$g����������̺(:ǐf6���5���{x�7.��$�<���]0÷�g-���6#R�I������f%�\$
b��PJh��#u��-]QIx設���4K�������B��#v� ؙ�vM����u�ˇ��u�94n�Pn-�y����<��7S�jð��]�v�e�nCzbs�{>;� �9�VN�R�g���R�������!*���u�ێa�Qƕgn�K��5�)�M��4n��<~�}�֓�6�6��[�5Wb��d鎫�;]M�*71��s�3`������Q�+���=��.��55C��[;��'�m�1�6O\�D��ʧ�rހ4m��ԅ2����]���Q�ff=d+�OG�kʹm��ʺNUf�pg4fǵ���Qݕ���جuY:c�O���׊[f;��|�m76В��}z԰LT/Dվ�SR;3�ջK�sސA�� F8ڒmz�	����=�� R��Q�[�:ʀ�ͦ!�+���-����7�!I
JdP��u�`�r�6�^-�5V�ÎG2��6f��սWWQ��,��9�� ����|�yJ��s鷦k���Y�[2�#��]�܇[���ޙ�;���Ǟ#|�)�5�8���Nݍ��k՘'zp����%��3�$5z=goQ�r�ﹾojV9�x�.v�L��H>ב��qE�&��}Q�"Aހ��:<�B�p �ⷤ\dL(�gK���.n�"jE�l-[���(w�lyG��6Ղ�^^!�� �YWn�58Mժ��xnǛh0���ѫ��̼y��������(w'i,��4����m�����@�����o;vI��ؗ�N�n���͋�ys�"`q��ӭyAy��y�m��e�¼C��p��[���<�<O5#=4�Oh��]b��Y{=�{�g�q��׺���#��FV��©�еn��\��#�=��!������1��kR-�/��RA�6�a�lװ����"|���ѫ��̼y����Az!����T�d2�e���� S�F��H ��"��m�6���UB��-���s}���6gGn!�tH�F�q6��|���s��^:��F4&<��jk'靘ps��>3Rn������xRϫ>�Qc9�˗s�E|����my��32ᴂ�
`fU�C%$7�s�_���_�q�u;���JH,+>��m ��!L�Vɡ��P(JL����罗{����yy�����n��� �(���j��$a
�s/�cu��`���� �?e X�?~��P?~�p�aߨ!q�������9������R����<	�Sٻ�w�lS�o4| ��"a
AH)������XT��Ci �3*�
A@�RfP��i��r�����̠�i.{G�ɂZ\ؤHi���͉��*��d��Llkb\���t��{�4�RP?v� ��S�@ZAf�Ja��!�$���3+H�'�B��lg�^\����H�$+�<��'{��|}���벘g;p��RA`s*�M$���D�Іf\6�Sh�̫f�JH(TII�@ZII���믫=�5�O���bAI�B�ʶM2�
AG� G�HN�{�QR.��F��?A�<��ô������j��$��XH,�2S̸i
��9�5�e���s���P�a߫I �Ϩ>CI��S�ˆ�6%$f^�
AH)�@ZAH/�fe�i���w򍹹=Y����7dا��g���ճђ�
��~�-$��?f����hS2��L���II�@[Pi �����
C]�f��7����V�R
AM{��42S�C`��
3*H�'�W�7���Ϙ̷W;���HW �H,�L9��ipJH,Mş��i�?���l�άd=]w+���Lm?��[��Z7v{�������$n�>G$~��i<^�Y
z�k��|����+�}G�+�o��BH����4�S�@ZAH.�=��m ��
`f]��%$*$�̠- ��.H)��v�r�&������f$R{��5�{߻��oG>����ekԐX}�높
CҪݻR�$��`i ��p���P�a��Rs|�s�w�w�8.�<��qZu�8��nw d�A<�p�݂򜚭S���h��ߨ;�AH,≠ibRA`{.Ԃ���AL�Z�
Ai̸m ��f��}����s�f~��n�g���
����w���������
>������]������II�@[M$�a�;H)
*�f]��0) ��s�}�{�� ��Ja��p�RAB�gujAa���?{�~9��7������AK���i �P�a��p�Ғ�洤�H)�@Ut�_�?fkWfRq�w��@�ܻY�JH(P����-$��³3P�AH,˵��) �P����?o�{t�{���K�z�QR2ި״'�#��v��#Xv�H.��R��4�Y�d��p�II��v��S2�Q$L�l�{�{�N��߮@�RA`Q�֔���I?z�֨��ZC3.H(��}���_}��?e���� �<���P��RAa�{��黾����R��Y0e$
�Iܠ-���̸i �6U@̻R�$��I�d��p����ߚ��}�������ACQ���R�s������~9�~�מ��
_��i ��� n%$N洤��
fP��
AhC3.H)���ܿڐ���Ӛ�t��;o��s�^J�L�b�%�t�%6ޘNsj�ӛ�23f�H�ߖ�t�ghLm9)���{�{������ӺwO~�{߳�#�[��"@_��K�9x"���Ä���C�lt�lre5qBہ�e��mSe�4&юъ�e���SM)1S	��"y�v�σ`9�㧝9������huš�gc<�m�t�ƹs\[�����c!%��\�1A�s��me�Y�<�H[�mvG�R�$m9|q9��v5MOt��vN|�-;�b�є����b$������Yn���k]�vB�8�q`�j�<�}l�;�e��f+��7�$���Ϸk?�d���D���i ��e�I')��v����)3(`hϷ��^�}�]ff�z��n�ô����ǻU��>�� �`RAJ����Af�)����6	) �C�Z�Xj0�����Ad�2�fe�HJH,�Q�~�s����o7Y� �:�AOݠ4j�)�w�$�Y�}�������f��
�ڐR
AM���<$��¹��6�Rn!L˵�����w<��_3]��P(���- ���;H)��R��I(̰4�Y�Ja��!���P���<	����s�9��[���Xu������D�����i ��� lJH,
�kJA`i�����Q �!�����̻Y�JH(W��_j��LkyϦi�hC�) ����Ci&��̻Y4�H(��� G�m�o?��Ὼcvt�A�[����U@��jAH)?~���I��^���{��t$|�L;��!�%$(a��Ԃ�C
H)�A�4�Y)��3.H)���iH,4�S2�湷�ۯeW��޼:AH/�5��m ����x�x���39����j�g�JH(RJO�@ZII�s٨m �e�����P)(�� #�6�5�}�=�l����TL��v�{W4�q٪DŖ����n�(1�Bv�6Ѵ��i�$�.H)�@�]���
~�i�d��p�II A�ݔH�'�><���X~a������AK��������}�~�~������H�I�_�ZRM$�hMQ �!�����̻Y�JH(P��2����Xv_�9��Ι险���!o	��3��!F���:GEN��0o��h�O'�O=�r��6�?�w���Ze}	�����V����H7�!Ă�X˵�����DAt ���y�+��.իJ�#����;H)
����Ԃ�
H)G�4�Y�Ja�� �w���=��p��P�0�jԂ�C
H)Ϩ4��%2�w2��I��v���S2��j�)�32�<	��vUo\e�{bf��x������`V�Ԃ�P�II��H)���f����b�̻R
A@Д���44�Xfe�I!�}��r�z�����}v������3�I���þˆ��JH(S�"G�>�3���
���VF��Dx(H,�e0�zᤂ�X�ݾ�����u޻כ��A`q�����Q �!���i6�L˵�JH(RJL��В�
��Ci&Цe��ٝ�����7��';6�P6%'�P�׾�w�^���~ˬʿRAa����v�RU@��jAt�����,$i��fe�HlII
fjԂ�f��?W����7�q�M��L�.����M�3Z�+XMA�YC2��.)p�h�%շzѐ��S���4�R~��I �7��ҐR
AL��TAH-!�2ᴂ���}��wï��g35�8��]��%$3���7���)9�����
=��6�Rm
`w�k&�RA@��̠-���̰�v�RU2�H) �7���7����- �ᒘs��i��<	��D�|'��y�O����W+=���CI��S�놐6��Xw5� �4�AL����z��o5���)�C��ᴂ��03�k4��P������II���m �؅03.�M2�@�7` ����U/돫'�w42�8��Ŏ�e�]2�fTKp�/�^S�j��/�����&n$2l���V9�j�,ig)E�����#�H�P&rU��  ���9\N�ڣv��O��@�;H)
����Ԃ�`RAJ����Af�Ja��!�%$eڐR
AL��4�Y7��x��j����� tJH,
=�iH,4�S�hj�)�C3.H(������Ὑ��~�t0+Wk<2RAB���z����X}����f��Y����Ă��)��ݩ ����
Aa��;H)
���v�L
H)Y��5)�f\4��������Ѵ�'R
�7�R
����׼sG�su���ga����D4�Y)����\4�R}�iH) �ei ��ˆ�
o��׹�����7�L�\�4���r�<��V��O;��18�뤽Z5/P�����ݬ�JH(P$�������XW�{P�AH,˵����R
fP�џo������>��.�*�I�߷a�i!�5ùU�S���|�~�R
AH)�e����Xs޸i	) �L35jAH)3(>CI��L32ᤂ�X_�����Ww��A`~i �=@h�R�높
l��}�s���fs�k�|��]��d���S�P��RAa\�jH)7�e������Ϲ>H(���`j4�Xw���� �{v�C�
fP�Y���fe�Hm%$(a�(��O���I�������g9z2F�T>o����
_(<!���@�a���@�JH,
�kJA`hi �e�Q �!���؁L˵�d���}�������o�����蒒
��چ�
M�)��]��e$
�2�����?{��5��k��̫�$~��I!�޻R�� �F����dL����r���޹�dX����@��O�^���8�阫x`I�ߗWG-���GF�=��d�K	�$��gX{wՊpӥԕ���$������?����~�i����0��H) �e�i �P�a�� m) �+3ZRQ�����e��{�N|~�t��Z@YK�$P��=��ïq�� ��]��%$)%'ޠ-$��¹��6�Rm
`f]������@�#v �c��O�~���JRJ�vD,Nx�|��\�rne�f�wc.�ìۛ�,oE���Aa�rᤂ�����.Ԃ�I;����3.C�JH(P�3V���~�����6��>��6�R�A�CI��f��}�ϲ~a�n�	I�]�����S;@|j�)�̸m ��)��v�L��P������%$�k߷�^9솒
N�S޻R
A@�Rw(`h�{����������U���n�ô��Xz�H.��H{ G�#���^@�)ꆻ�]]���I�A`{�ڐR
AO�Pr!���L��.@�RA`f]� �̠>�RB�p�AO��^��8]��Ǣ"�׸�~ Y�������P���z��4��
9��6�RlB��k&�I �el$�a�i!�ƨ�}��{����}v���S�=`i �@�L?~��Hm%$)�f�H'�BU����"��O2�~�<	
���%��놐6��X�VϽokn�����Xi �ޠ4j�)�=��m ��
`f]� �̠-���Xfe�I �7R'�4�Dk�ʲd�w��@<�>w+w��NT����݅��O�:P�AHz�޻R�$��XH,�d��p�"JH,˵<	𮡤�J��9?7e��5]��A	�'b�
M�5;�R��ܸ~�i�M�����������>~�K��H5�훠�[�6����pZ������=}���:ke��+vh��h�7���I��6	!�;ۛ\f7WZ�i��'�/;0,L����ɱ�U�z�<��t��ɲ��M�'RZ���Z��`U�4&�k�u��Ɨ�8��k`t^F(��#F�hҚ�U�j�j鬴3rd�#��[��&�Ý��y�t$4ƚ�Tڴ��L��6���DnnNk��rl�u�V�����?�]����P����h��b[+C$l�c����s�]ҳ���:���$I�$�S�nH)��٭)���AL�STAH-D32ᴂ�
��û���{? ,�����ނ<	��?�{W�����-II����I&�B��v����)3(`i���3,7��P2�� �`RAN����w�>��]���|�R���Hu%$V]$�����ߍ���;�����6�R���CI��L>�놐6��Xv�T�R
AL�>������[�� ���nH)��~�g) �BJL���JH,(��Ci&ЦV]2i��P(JL�����[u���:�Y��v��H�o�ݏ��c��$AHzU@�z� �`RAJ���4��3.Ci) �L2�� ��
H)�A�4�Y��>-�7����4��) �(��T�XH)�(H)�C3.H)�]�}��{�}�?}���0*�� �=Rs���%$��{�r�ך������L�e$
�ݠ-���̰۴����Yt�]
H)Y��4��3.C�_w^������	� �C�ˤ��I]}���d]�i��߼(�B� "<	���a���i ��y�H) �e����Xfe�I7���}��+������iU�VZ��(L��4�X�JRhM4��f���gA���I?'����1%'�@ZRAaFw5����˦N2�
H�����}o���G���>$x�Px�
C�ϯ����������I ��߬$j2S~��HlII
a��I���$̠�H,�2�fe�I �5����{��?t��}��r\�V���ckV����[��ۻv훽���{�w$˗.��{۬?d1�h_��AԔK�4�׹r�7�� @!�������$��STAH-!����m ����9��}���ff��U�$���Rs����P�sP�AI�
`ee�'�l}~����
AO~�- ��9����v� ��R�,$j2S̸i�) �L2�� '�r�y�?-��ʬ�y��Ȼ�M�F�ᴂ����Ad�S���HJH,
�� ����ڢ
Ai̸m ��)���L�%$>��y;Y��������;RAaS;�Ci&Цk.�4���Q)3` ������ߒˑ�?����O�:P�AHx�����At���������f��9��@�AH,=��!�%$Wn�0�����MFS̸iiI�F^j�Q�������-��Ͻ�����^!��ᴂ�ן����}�﷙���V��Ј9�"|Yg�����6r���tM6	4̦���6k��v���s�N���A�2�I#�zA�f���ڲ�2D�v�p�*��yQ�"��N^Fp��	�8�1Il2�ɷ"K,�� D;>J�Nҍ�iÞ ����|�fU���͏U�xO��Fj�m��c荸�G���_r��2!��[r��Ī�{����s���3��^rk
�].I�cC���wq��w6%��8��0�X�D���0�>�e]��ؼ�TnEM�bs9�u���з%%�TO��gynVo&���\�C��G7췼�'p���\n�0��z�wsz���6����/���0��5���1�{��2�1�zVz������.��59��q��GF�z0[Y���{sD�	�4��{l-�����F�̆�J�JC�"�O���=�۝�q�s�����wX9x矦��K�O�hn����Lc�����Ǝ�0�n�ߕ˲{�<T����3W��&y��~��Jxa�}��`޷�9�bd"�eh{mk���L}�x� �<���4$^S�Qg��S�/n��J�:��I�*.k����2�l^m3Α�Y�τ��78���i#��د�yܤz�b�#������~�����g��ƻ���q�v�����z�[3�����g@F�hU���������r�E1��͖2`^�D;��j�.wj���p����g���v��La��l��vY����Y^"ὓ��p��pJ�}x�%��Q��=�֌/���{�{��
�m��^D�h�f���v�Ne�7�I��	��>�����W��g�1��5���������5k3�B����f/V������jAn���j��=<�]�+��ou�z{��-C��_�n%`�x[9�x���k���9�jǒ�>�;�pS�#�nU� '�l=4���<���ʆ?M�N��y�#n�GEZ�s��Cf8�8���:��ٝ��dvYm,�3qڙ֙eё�u��8mV����Y6s�;;6Y��(�݄۲NRn�kf��Dڵ��Ck-��l��Ƞ3:kV���Yv�Bejf�q�ٶ�miYFr&u���N����v�'CjKf:mu��i�Y�ife�k-��u����-d�,í�e�C�6Ӷ��gE�&����vem���܈��r�r��Cq9r�sm	#2@�m�k�k`�Y&Z�ݙ3�����m;�l��pVe"ִskKl9vkk$���eqtu�I�%��[L�ͬ�6���t�Ԝ�e� ��$0� xG7V��A��]��Փ�A7���nD��>E�^!�2.��q��&��"H#9y�^��f緫��W��ʍ��@���� 늙� 6׎7"Ae�/� A�nD�Y�;Y�#;%@��ݮ����ˎ�3c�s�A�� ��m�� ���+�Z�8�q�~��XoŮ�#@%�a��X��ӳ:����9�7�Ʉd�!	*�20t��ڐA#���mȐv�pz8ei.�wjɃ����]wUn�Ɉ��י�~ �� CnD�Yd }���[Y��u�OGL����(]�E���\ ��v�m�J��&���'�^d��6%� A��,�ŸyU�2�W�3y��r�e���C��!j�mX �����`�q�!��Cn|{k��ZK��ڲ`���Y�#N�ܐ�QH����;��5���-�ݞ��0�_{�I�E=�ͳ#�T�]q�`_���������Qg��U�N]�����������y�r,�6��m����VM���5��F�Oe�mp�*���Lm���|����myx�ۑ�B�
�ff*����*A�t�s���i܌�+e�
���cTn�^/g��!<��ka|�dIe�>-�}�o�''/�Z���2�K�}�0�3�^;���8d Ck�y���Z��Q�ڂ����nD���xf�/+wjɃ�}m�Ye퇹}"P��"'��%�!��mI8dV
����5םLRY�o&6�W�S�Aa��myy���7�ޫ|���c�c�A_H�ŔA�n���n���閸fǮ焂l��6J��7F-@F�^���e���Y��94*�<��Y�}����99�;p`� ��Dmϙfϛ��X�3&,ۇF��9!E=�7B�����s$�3ޘ2�ӌ\��N��_hs�����s���Z蛢�<��S\�f����i��W����EY!��{� Wh�D�j0)��4��U�m �m]y�r���D\m��f�'jzD�8�W����'�[*���3�ز���粼�x�&���dρ1���;���s�줅�u�ۄ���ms�&8H���n܄Hٔ�.r�pǌ)�k6���:Ү(�s���@ ���鍐ۓ;��?�s����+�q�9M��y�n�mp5�Z�w�������W �_F��s�ʔu��ȓ&&7s�wG�(�i0�j��Ծ��{>�q	��=�$�Om�p���/&7_!F+�72.B��d�d Fj��mȟY^ ���K��V3�M�'\'�ݛ�r��].��U�A��٨ [jM����U�׭��r,�U^��z\2Ǘ�nF ���¢�7]n�[`��������}x�Ie�%�^!�"A��.n�J��d C��6��!DS�Ox�+;.^Tn�v 2V1�y����&ח��>e� �[� ۑ%�wxr�D�p�ve�~2�z�����V_K���z�!���A�"�RAp�J��Y�珨y>���#����uVcc�2�jL=��!G����xůJ�>��|��s?VB7m�`�{�v���prsvw ��t���gB;n=��9�"N@n<�~�|Yd/~|s�)��8FzE�E���p�웫�W2��ͮU#�c��:v����gn�HM��?8Ή�b����fx݃X�*.f  �����$q��")����7ݖ��n���H�@n�kFu�#�D��e@=мAmȒ�(7e']0�{��f���O��4r���.gO�WO��s�E��C�B!�����j�En�y��D�}ф/�㘂+7oY�.�N4�� ��i��V���Nwm|�vd�e��/ۑ>e���E��&���F�"�)�v82o��9����9�I��Ch/6���NN�9(L�J��fkJX�e5��s))0m�ǅ���:�:Ӝ�*t�$��.��<�,���ݼޣ���]g>�(9���Ol�
:d���z�U�p�D6��jH�Q�y��ˌ���D�^��%D���=�����܃�>9��x�O�e��*�q,��tY�dp��-� �2'�f�fWl_U�ձ��L�F63T�jk\��l26�/n�9,�1���W��<����oo��7z7�n����  ��f�{0''�-�����y�RA��yy���Y�Β�܀خ�n(����Ǌ �� ��F_:�9�4��zA8x���a��U�fă��Hg��@����d"�{��s�<ܡ�X��W'5n�0{�s���YeKqǧ�����v��(Ș<=o2�.��ۗvQ�LmDY�Z6$�`�g����*$�R�A �d���S�p�B%8}��s������*����:4D]3��JH;B#���܉ �� �� �ɒa����t� �p�ݽ��e�S��O���!x���-�X�2!)��1���!�6Ѐpš�=[m��oi�5LFNj��`��tynD��(�p�m�j��U2�L��Q�Y8d�o�d.uF�\n�^y�A�|Wt�N��1Aw4�fOS#]�Ed[�`u��(���݋hܚ�n�ģ�euvE콂d�6�̥<e�UV���?{�«H�����"Ae�<|�yy�"Ae�6�P�����J�z>z3�)���s�A�A� [jH!�"/!_�<��`Q5��(b�n3�-C4s3����n�k�0i��t�f&�2(\��smO�##H^!��nAP����"�d��F F+�9��c&7�["N�P ��x���|�!IuN����s�;j|;B����Q�W�3���) ��B7z�W=����D�<Q�l"hIe�>-Č0i�:��͜��Jo4i�\���>�A [k̲,�ݸ�_H���T8�vǓnAP�����V��[�� �� R�jx�e;�yA�e����@��,�-��msu����pMJ�B"�c�aru9gpF@�^r�F�@n<�B��Q��Z6��B�%��l��^ׄ;a)����XgP�yz(�y��̤CAJ-<gjI���`��&�cؿ���;矡���T)-�2;U�0JKR��F°#��۷:��@��aq;vRT��o;s�ðb
�\1�lV�]��^�](�gu��UèM��6�ki��))c6��1,e�5��ñ��A�5��Ѕ�Yek- Ɨc�;�o;S�<g�#�c*��G�7hR�ɍu����5�A:�q�[�!���g�}�q��8m��/'gv�����������s�f��n�08SN��t'O;�KW�׍��XOb��>����Ñn���ۧ;1R��}�=>;Y�=q1�ւ�}�H.�6��jH��Gd��Gr^#3dH�O�;�U`��ջ�����"K,╩R��vSaB#�H�OB!�mI�#e���]�W3p��m���\���6�Ia��n<�B�,�z+n��:.:��*f*V�� ��,��;t�f*S��O�+��a��{�g9<��7\��<@n��Ԃp�@��
�;1V%MFy�Z�O�d�cރV1Nl��Q�Nt/^9�,��1�32�!׿���{P������v��k��Y����	,r�������&&P��ߤ,�A�5�ڰA��[�sJ�.2r�،�#7�M�DN��<��FG���x�܉,��A�@��\vv^�N`��]Ԅl�Y�4��둗:&�Y�{g7Dr�3��e�N1"o�p+q�D\=��D�x�<ɍ��� ���5���{��<l�@�{�d��?�3�)��Ք�x��#6��iuGu���2,�E���1�O�2ǓnC�A��Üj�o�q/{w`�V#'5=�Q�K�@C�"|Yg��x�܉������h�K^�k�26"���F��\����^��Z�-�'<�C�'�N�㯤H,��%�^ �܉,�Fp�R�a���AW
���u⨜�}Y\'�x�A�Aڒ�E��\˝��ˤ6��aI�z���"nΣp�<8�`�Ձ�f�6�ɵ��\.�H�"_�w��Y��hH��o��a*����G�Evڳ:Q�[�� �s��Y�~#���^!�7&k�����5>!�!ST^�.K�p��b3�%�) �a��n�b�����(mt��<��,�7(zI'��q����qI�E�J��R!5�Q�5Vq5����!XR�&IK���eL�O6.�gl��9!��������ޥSb���⨜�}Y_	��^ �6Ղ�B7/�41�fܯ_�0�C���	��v��^V��E�G�5ލ�=3ya�6P ��@��� ��	���5{v.��Т�]7U��%�8V坱�q���/6׌\3}Ճ4JC39��גڧv[��NF�x��=�[WX�D
����� t�ۨIe�>-�����;3"�+8i�e�i��}YD"&�ݜ�\2!�%��� �ޖ*�q�K�H�Bs���%*��p�G�%�"�Ȑ,������M�&=��$<B ��-�$��#{Go��.��4�e��e،ཏ��4�!�����(�}����=��c�N8��t�<t�A-�;t>��̊���՗�}��Dv���
4<�.�(q���#L�\�L
�
�X6sbՌeN��U��%g9"gL���L����B.
7��U:�Klj�>�����)���!����!�!x���M�S���t���ә��)*�7���E ���76D��ϑn(N�R�}����uљ��Ύ���<l�����\%�`�V��
D"J��Y���M��#9[k̲/f����Ժe��e،�"�F;y�� �d堃�B!�y���l�[����5�[��Z��x�w�ygn���pVe�������!@�A�AK�o,1�"5� N� �d"Ax��"mZ�5��)J��ފJ����G���D͑%�P ��/ۑ"�ɚ��Nț���jH!�!{�����Ժg
ܲ�F@㏗�R���O�ɳdqI{7���~>n6כ��dُy	:Cݔz�_ܿZ.;g��ח�A7��A�^m�7~�o4��N�M��T����7q�N<�:���.�M)�R4���u�o��k��u�oW)��}�7���X��w������f�s�(&e�Ʉ[T��{��޸��b �_ePtG��a�����E��X�r�����jxk>Ӄ�%7'����t�<�ap���Hß+����9�v�Il%.��Q'{�ዑ���g7�
^琉�S����S'I�7���Ѱ�3�'��h��l�9�>+��N������y�/���S��u-���L;�'�y��z�b�}�s�]�}�������;�_��B�/6xƩ���q�1�W��`��&�4�"��'�FNd�ݯx��xއDu�qH�����J�A<��G�����aRs	$��^�z��T��8`���w����M{��m�ta���F=�싪qZ.�,P�t�a�d��yT�XZ�.AÝ�	F�ҙ��/�j�2s��-@d&�K�}��0ǜCX���[�9u��{�f>�l�g�^��ޜN��X�;z�l�xC|ww�|�'��E�齋��ƶg��~��+�l��>]��o�W�Y��'��*˞S�6eSu�r�*ލ�u����3w���+<#�e�OX�l��w�þsJ;���/��>^)WvJ)�}}�x�}���iG7��n$Ɩ�=ے#lX�Mhf�[���Y�l�]�m"�yl�=�{mX����{|�.���s��j_E񻾧���
���wf^�jK��F?:�hd�o/w��^y��z̶gG+m�1�N��7"$Y�v��3�i�(�9�i�n+0�������vgvs5�#��E��ե��m���D����Y�gn5�B�n�g"�ݝlĐt�����.k]�m��3k)�vK-��gL֛V�E�md!
��h��kp�ӵ��f����K���Z�[M�6�Zd�i8Y5��P�˲s30Yn6��9"9CX���;t�;��D��6��٬ѴV[X��cj�JN�����,�1�Ón�vr8ӦX8r25�%e��G(r� 9��8s�ۛ��H�kp� �\��De�E3BV�-��q�d��W6͍�k'mڔ�l�
$��NN#[V�BQ���-�8�:�4�<�oI�����u�W��5�wc�0��n���٫��8��H,��l�5uqj��
P�=e]ŷF[���m�P��������Z����t��Hx˱ϳS�{a�4p+git�ô�҅�"VY�X��lJm*Y�#h���Mb���2�����f3ά3],Ю(�if�(	�]U�Y��k\�V� ݎ��d	u
�G���ж�:��c�᪶m�,��[vg8Ó�ex�ۡWq�M2��yo�HD��%�,�Ll�������ey�2��hh��Z���5�ѫ͆�����<�;8�Ei�9���̼�w����8Bn�[�k5��#�����Xb(�q�ѻC�l�d9�Z'(��gs�K�UzN�3��=�nbS��]��N׋.�˦��	ѕ"���9�a��{E���o����@�X�8��˩p��#�Fh�]�53�jض�z{��n;+.�'��}	Y�1��`�|`�{]�ێ$�L]�k���R�m�:���r.�����RQJ�C�`q�Z��̵�0@�X<$I���4�h��ָķ$��Հ-]7��1`Y�Y�LZi)�umE4�*�W���Q7aTjۍ�I��Ѕ֕�Ƿ;[�68�W��(���k��.Iu*�֩ܒ�L��(@Vn�ˏl�*v݃rUr�X������/�vS�'n�S9��m n����0��z�.e랂�fz���d#����8Hʆ�i.f�0��+L�Sj�ͧ[���#��}��z$��l8�Kj��=&s�<��e��Ny�;��)��[�'����k��ϬO5��,&;9{�ص��1ˣ�3m��ql���`A��1/!͗Q0�5�Gd�-!N�l$G�;tw9ˁRK�{����f!Zzc>n��]-h���]�4�3Y�
gM+���=k/e��.���4k�0���
�ֱ؁�3�Hvzi`�g��6SM���Ӻo<�m�k��v�<N�P�z�z6fTv��Y���ncF�tRC4�[5�	hi`V&y�����ѥ��'Bu�Y�qO���eq�O �:��'HuÄ�Rt�NW��x��Ŝ��ӝI�5��C�+m�.��+n��v���E,�Sm�GJK�7Q����rm�0R;��S����,�,�`s�i�#[�Q���,�n����[O���0�ԃc�s��n͔�Acu\�;K����
-�p���;RA���6��[r'М�go
J���n6�@��C�"z/�urt�mؐG�q�E�;s2a�0�^ڟ[^@lЗ{}:�L�[�]��@�|�F��n`I�=�ON��t�;���8@��܉-���ͽ���37��y�f_>��8�G�٨/ڒ�"�Uo��Fl_5 �+W��|��nD�s}�xT�5c]�څ� ��D�Y��%t�Q�z8���мmϧ�ǐ ��E��v�ɮ��F�J���O�t�+r˱���Ia��n<�s�ܾ��ؐ���D�RT�0�Q���..3ཉA����Y)&�]��%3�ݞ�e�g��w��p-�f��0���ѧו�9���Ũ܌��V�7�O�n<� Am�7��:�t�9�.VY���	���7p��r�䀆�j����:�y�P�����Ut�K�S�m���mc���w=�k�fr�No��
�F�m6v�@�A�}���$�+�zt/�&Az<��E��Ck��!A�j�k3N�r��nYt# w�>RZ�!����[���yϢz.���z}�s�p,Kqۯ9.�833p���p�M�yǺ�������X�z���3��t�Ԃ�"�0:�>��!'��xT�5�i��
<3c�sdIn[�mF�hk�)���~B��O9Z�iwC�htKS���b�� �l��VĈ��@(h�{>Ώ"��ڰA�r�]l_lGL�{�\��#�[FnmնNr�6���x�����	n=U��i��&e.���8=Ѐ\�sx�^d��:}y]��G�f�6�u{خ���%/"*א';���^@���6�&�D����Y�axٛWao?�೉9����� V�=GL�kb����������[�v��>�g��V���ˬ#f��s;YN&�B�rNR��/]]��UQ�i��
|s��ȟ�"-�!�����b;r�� A�^��~ �ח�Ugo�#�`��.Dgy[�$n^d�����t��v��z|��"mϛ����Qág�b�wq���9��t��c�Fl[k������lG�pmI���1��\�t-偕�5����1��!/�_���hW;g�cv~�ϹI���6���	;ߞ�UQ�i��(�D�����܄>d��-��/� �p�m̂[�"^E����R#u{�Pb��b:�ܲ�F@�[�����Cu��Y93�	�'�A;��AmȐ[��Ÿ��[�Їs��y�g��#3^F�^R�yjŶ�!��Ck�UPC;{)����9y;P^-�!�vo	�U5ۍ�P8gB4�2Ī���lV!�9^T����4�=�<2�S�N�U�u�<ie�V>�y�B�e2��쓮p���9�����	L2�Y�8�D6�H �^ ��@��Di�E3݋�y)����0^�"3� |���yK�6��p�9k��;��%H0�&
�ܗA�����u���=	��VB�F,�-���_�p;��P�>��p,|[����5Պ35�i�e ��>�u�������^�א!�ڟ[r��3��]��}�LJ}���ʪ����(��E�Ȓ�}�Tu��G�"z�H'x&כj�A��2�UfWU��u�#n`�������yx���6�H-�Db�5'�_lg�>���x�[�����=t�/9�@fWH �G�F��U[3�����^@���RA�k��7Y��7��G��H��O[�*�0f�[P�p ��^���������Zӹ��Cv�gmI\��Sb&�k6�A8�Y#�t�(q"�S�D�3����i5Y����2'1�S�6{8�#��<�Ml%�lB�s�.p'�s�zr��78����Lŭ&��jl@�G��^��u���w�TK�w���y��ͻG��n6�C]���Pg	��z�������ט�+.�&zݻ�c$��ծvˑ��`�%�-�쑰���C�I��K�r�!Pأ����1�dv�����$�h�$qp"�)�T*qV^����_��Dq�=αbn8f�leY�Z�
ʽVO,u���)����\y FlmI��ئN�wDr���Ñ�x�&�=�Id��^^#5�ۑ ����ZcF�tlJ�e��A!�;�9u�LVk�@fW>��"Ƃ��V�v��YE$��"m	�k��׃u��ۑ~�N�R�o^N��*&l[�N�@�N�M�nN,0Ppe�sp-3(��[��4c̉���|A��S'g;�r���a��q�#�s<����?H"��|�H-�@7�ۑ � n����*ac��9u�Le��@fWO����-� �k�c�S���$���.��1���IU����Y��>�l�Y;S��-��;�	�jH9���y܉)�c��UT`Ͷ����#\lv^�w:�D��ϐ-�6АYd
d�wI���}ӣ��k �ʾ�U�����;0U:�j{l��z�QU5>�TrOcZ�
�5OW^,�1��3fh��;��Lf�,C���$B��L���Q��V��^��H;��s�:���b�,6P�a[r$��q��R�c�nv�ٺ�[����A��AڐAAk�ԛ��%ak���BwG�h�랢��0�ڂ�	΅��j!��gz%Ċ�������p�Cm	�B�E��E2�N9C$��!˙99ڣ�ƭ�� ����d Cq��܎ÛY��w���o�]�4`5*m^!Z����YE���ܶJ�0���g��=4��;���O���>���l�n��I�Wk�>y(g�.��uGd�-��,�!� ڐGH�;�p��(���zD���.ޓ
��m�ڂ����/vD�Y��������")܉Ǐ�͠�m� ���^��39q��X���u�'�r��ǔ��o���	�qL;�h���x�7G���M���q��~�O�$���PިX��]ȓ�v��)��9��^�v�!����nD��(��M�<��".�6�I�dO�<Q�p�����vT���q��%�08�GTi�����b�z��q���-�$�C|���s��}Q�h��v�w�J��m�ڂ�x�s�@���,ߏ����*����}����Z�jcv�b��Ѷ�pRj�֡�&�`�b�\�S"�be#mz� hւ����I���r�U�m0Ќ���*]e˷g7�Or���28����mϘ���w0�؅�%YO7|�q^uO^��q9��O�J ,h [h�����D^Z���D D�@�xԂ�2Ǘ���ͽ�yy����b�m�ڂ�A΄=�"K,�A�@��
��ͷcf��� M���C,��tuNv�K6V햄d3��FuNP��:�n�{v����r)U�
����qML��Ѕ�E�A�㯺�'�Y5���!�����ҟg���Y�C	�&�a�D0Er���}"K,��[r$��9rr��i]	�V��=�%�v���s�A��8�E��.���':��ԙP�b����l:k05Y@�i�X�ˆXS�|�����2l��c��5���B!��[r"����*��nv����s)�S���ɋ ���'O"�y�����@�.�M]� �J����� ��Bi��9�Җ�-�-���H>�d"�ʼ�46E�����6A�;��6�Ie�������:����L���˒�4k��r�G�^#mz\2�#��������� �p�Df��mȑ�b��w�+�V6�mAG�}����Q�����ƃŕ�/�۟O�d"h [j��3�2�dHJ8��8��-�Y�Z|�9��;�m��&g�ڧʹ�25^Dƹ��t_x�m���d>k��#�y{�rJq��'��;��L�.���Yee8����`Ng�����'�L�W>t�^x4>.cs�k����7gq:�Fr����\Y6��@/9������%�g4��sT��h�U���G\�����k��3������Q������Pit�6��K!� ˦8L�t�nRB�c;A�y�c���3��m��Rm�.�m@�݇Bn9w(F70\[X�34�w'h�Qr���Y�[{gf�����Ff��e#r�tř�1ɳzޟa�gq�^(���6ηWh�OG�!��.!��׾����zVL9��{�SqNoU�z��>�Ax�r�,� ��/�R}�+�_$��D�^=�"qLm�n�sw'm��x�s�fȒ�1���e#~F�#u���� ���m� �dt�f>0�w�^	��Ǫcv�w��s9Il2ǐmȟYD%���A�x2b!�af��uV�z#�&�z��zA��"$CEm�G�cO>S��!HmHᐈoYXbԼ@ٙ4)��{���ؗ{[pQ��t/GfȟYD��V��݃�t��2�8�v���D������Me ��tl��zG̟L�Lș�	���A [jHe�LlT�w;����p%	�X��e�6Vx�6B#Z^m�2͐Kq�y���c&*���Y�u�!u�W,��5�i�l�����n�?�re��k��BiV3I_��Ki�ld��[��y�jlA��᥌�f��:x����[�90��k��s�	�� AƂ ��oA����d��B �� �j�\2t��AiėP4�N��d�]�W�� ���f�~,�� ��6з�:���<Fm�wj�!�"6�ة��
wk/p�|���H9/fzq�ձ��H�愖YD[�>mȒ�;kDԵ��7yۧ��]�i�h���mI�!��gA�ѷ��-��`@X�8��en�;6JϜ�:���:RIF����R�ubv��:B!��nD�٫��ɫ��������;��è��C�w�Iç��y�r�,�Nc�<2��]#��$tq	m1�}O�L��^�r"�{3������N��=�2$:@݊��"K,�An+�.�&cy3���mD�[c#9y$j����j�E1�~�ܖ7�=N��:X��x�x����i~���{�ڵD�'Vͬ
���:^.�Fǝ�cgr~�1�����9N;뮣�mN��ov�i�e�8Q�?d�L�Ŗ��M�+a�$�3=�c�)�}�G6�j;�=�m[0�fHj��7H��C�,�nR����C�{�:l]e�^���;O�$��qs�^3��2�sD�tU�ƫ�O�y8�l_$bs��oə��{Nza�7xN��~�~�K���F��h���w=7���|mW؃�NlN�Ε)������&X_�+�oA�7�̈��(�xxS��̝[�m�(�ٖb�jt,�,�l���L�afyn!_j�:z�1��
��O7���uz|�hB�Q�|��o��>-�On^�ۃ�����ȵ%֫��7��L�(����v��k�L�4AlQ]x��]�}K	�%{7u�x���K}_{�B��q�=�&!��j1�=Ͻ�j�75?m�_�pcxP�h������z�����ӣE+��9㛤cү�s����2��x�O{�� ���\󞅖��0�
،��m�Bll	�����]X㧦5�{��k�ن��;yy�L�~�wW#R�+y��D��ׂ#������#��m��>]H�u��`�_F�{�HN>�[Ƶ�6I�X|����pl_y�ʯ����=l��}���k����ܶX��6j62�]\�ح&�=QQ�7E:p�m,�IڗP�>���)-�m�#�GkLvfQ	�F&"�jЇ:Jd�����tᵺ ����IZֳ:vu�6`���kqi�9�qg$�`wh��6Đ2�)�iV�ضvf����R��:#��u�Yegn�ą;'i,�N]��Rm�!�&I���G i`�ʹ��͎֭Zdۢ��v%ĝ���A�V�vڛZD��Y�gYd�s4�mgJ@�e3
8�.3Y��e���mgq�A�fhNr���+3�29)�m�,e��H�i��mݧHs��BFn���'m��[kk8vڝ�m�8N�ŖS��;R.�ݛ��60u����C�ȳQ�M�9�m��3	l8Fء9B٬9(�9�NN���' �f�tru�v�r6�A�j]��꬗S�qƑN���<@X�E����m1����V"�@�/6П`٫��ɫ�������}f�F�vX/Ŝ(����K,�!�m�����sb��:u�ŷ}�V�e�".�S�� 7Ax��[��BROyMr�TT7n̐s�fܷ:�-��m�ge���ޯ]m�Py؄��N�M8D�2͐|[�6�[�=5r��8�)�H���e���T�@b�^5 �!�͵> Χ�A��K����7����W���WWa��m���� �͑%�pL�q ���>7p��ِAgH6��m� ��"��&��m����w/p�\�3���d n<�B�,��ɽ��yP'6+��b(��Ye�nۼ׺z��u�f5�VWH>��^��+U�f��\oB�g/FK�UJ�i�=(�{n�(�ҽ��7��a�Y[ w'��(y]���۞���N	����8{DF�;X��x�Ch Am� ��ޔ�8����^��1b��KN�í��FO��Dٲ'ŖQ�vT-�]*;(<˧�A������D��I�����pRmA��m�-����Ms��R�¶}�����g�hC�^m�2Ȏ��e�����DWy���f�a�
lf���a�Լ[r$�+��z��ܽ��8�פ�`��u�nk=uon�fC���<B��Ѫ�;r�P��*$��x�� ��B���r5���2�`��w�m�Ue��m�'�o��vl��Q�ۙ��9@[ �(�h/��,�]L��El�r"�s9H!N��[�˳�\A��坳�Y��p�!�"K,���R!��Kj����oN[�Xq���H&��#�mY8g��Lb6�;�>���;�]Q�Ft3���v��A�=3���[��̉zk��J�5-��nX;NT�W,fb�^#�EC�L�h�`[��Ib;�w�(�&I�P�*,���J�51[�n�n�˕ZF"	�K�X-̖�˭B,],FP�T��6�{;�n,v{P�P![t��5�;���p�E��s46�4�R�q��36;Y��'X�����a ��ڷ<zb���Ϋ-����Ǵ�6`�ѫ��L�TfB��c7d�Ѧ���������y�*䧝A����^~�����4\��#+)�t�Xj��Q�[��j3�Ɖ���[�-J�=+��������n<�r0O�w��x�U����&O��C�.2&N܉ �e-Ǜk̲#�Eӕs� t�m�Du2w�/�El�yp�Ew�>9����@lc����5X;�~Sr$�Ǻ� 6�Ie��	n졺o���+'��>���v���++�<B �h"�R>p�D6�j\
��u�/���� C����ۑ8*�5�vbuC2��nJ<&�#%kN�e`���8l	݄CnD�Yd Am[hw쁽��3Q�L0F��Km�p�٬yiЊ���^�Ȳ�&܊�*�)�.�)'��&c\2�@2���&�ũ�6h���,���ɪ�R�"D�8t�uwW����]ٛ�{�-�e�8�
�C�c��wf�����d�9�#� �a�̊nw���k_7�3"�i�7+���i��`�Oބ	��+"�<�j�0�.혩x�ONK�V�t�4Vu�;�.�G�Z�h�FZ^>�B¦�{�1:���nJ<A7Ѐ#�=�EC�z&Y����c��i�v#���,��b'+��v	z�E�],��[��b��p������B��/f@G�k�r�;��Y��W��^ ��[ٯw��-��8���! E�"�a*���a���B#1/fB� fZ���\����@X[��{��*/v��'���q�(_���}̐B�g�@?C��RmFkoc�ں�%nM�'6+]8�{i�6�nSL���-����'�C��1���$�BO4o&�xDnSy)Њ� ����2c��u1$:8�E���A�
��2#We�!U:Ev��`�� ������v��^,z�_ A�� E��2+;�Fb�Q���0F�E�^B �����Vl� {��W߮畧̇�u(.����}��j}����{�:E�E���m�s�j�u�u�Eä�nn�έ�V��}��aQ�l͠ƣ��7����P̨�ے���D�8p�'2��m�ư����4�&�E� F!���n��F���N�W @6�*�[�Og(�U��LQ3.\O�Yq���/9V��<x��4u9�I�X	�[}۽=T��Yode�@�<Bh#�r0�EMV��[��[l���*62�]�u!����a0gZ�0���ؚ�n,ن��`�cZ����;B�]I�4��^^9�+F�^�vZ٣�V�mx�s��I%��U �Yg��Df%�8@5���}x�;KP��WDv=�W�"5޼��"� M��0���7�[��_��}U:��yʸ��Yq��Xs"F	η�/7\�Sz3-e��w��� 6�^2�##Df ���&�Q��7��pʊ�!�/�X���ݖ�h�U��x�� ExS���Z�P2i:x�3^��w�x$�7�.��]׶�����40r���zG^2�{��d�e�ҝ1��H�S:fƕ'��˃���c-K
(�0Z�N8�7�w�[B;y�Z���q��Њ� |m� ��3(���(?n��E�G��⧙s{�cI��n��q+��Ϟ[�Y qu��\4�G�V0�'�y��}�=��s!����2�e��w�B�luI��^�!1�@�� ��� Fdd/�n�<5Dh�P+�� ^5�ڂ�O{v�9��V�m}�7��|� ���gT�b(���"<A����z�l�ə<�p�s7��o�L��oax�p�Fb�1>��%5S1�K��e��#�wu�꧚*�e��w�d���v��{ Q������2<���̴!)]�s�	�����T']�W;��<��x�|�#�;7vn���Χ&�	܍he̔V^�K�z��J(ꀞ8�F��M�x�����y�����ا�p/j����zq��Mb���$�-:V���ll�m��[t##�WWcA�ͻ�\*�]�;JA�AE��/F�\4J򣗵��e%���ַ�p�Nc�»؅�o9��l�m��B�F�
�T-%�׃P�mT�� n��\�ͮ�m�����BJ6��$�:�׵�a!���5��	�UM�y٩h���!Zk��Q�#LٲCbW#�aX�#����|��V<cM4i,���]B�Z�yҹhJ�KKRۤ��i��R|���^�� A�^̊ ��!������Fv�T4�U�+ل>��#qy{2�@��=:iġ�:��4�¼Az^���꧜*�7�"�x���d<\����u�$(����Ј>��#1yx� «�̚�<l)�����5s�H���"�(�d/�����Q�_ �΄F!�ۜ�k��[�[B+� �N��og���E4�{�@����s����g3�ݕ�P���ַ��p���l��'�Dc��d"�F7�N����ꃽ[
L!"��f�c]�f(�avԶ�5���|�k1�BԴT�ѓ�;p�=@̠�s^�]����-�ɫ��Eo�Ժ���3[D�� ��G�(�8@޽��!#�s�ǌl��?ޟ��g�����K�t���[�n�4��q>��}�T��[�?�QU�V�)D��a�t7I�[�8�������j|-��^Њ��7��8��k_529�P�}��AG
	J>�bP�i�3`�v��ޛ<Ꭓyi��|���1��dyd`Ń-K�c�r���x`���e�}���[���mnfM���{�}�/e�S4eۿa�D��ā8p�A�/�1z��� ��DUu;x�>S��'h*�	���q�"3#�و}��>�����ϟU�nacn�U���o3�n��(��®z�4\��Q���c�ߏ�]�}�
�m��}]4���M�Ȼ��1��X���й�I� �h#�<��� Fb@����Z{��L�!����Ƃ��b��w�ܼ��[PQ�7Ј"�p���U����p(��1{2=YDe���F֒����=O$�qѲ۪��"C9��ƠT�fS7<�v�=��Tp��<F�rsb]��ʤ}�aZ��J܃'1�޵jz���NК� �^ ��#1x/��8h���jp��&-�k�E�(�s!ow_WM>g2�y�.�	��/��9dm\�-��`�B �\q�ā9��>��#2#:��]�b~����j���fNc��(��B_@@��dO4V���&��A�
Q�H��$�Y��GA�	m�-��FX&7.�{3jL���-���#Ǎ���/�Dda	���k]s3/[̝�5�5	�����#c�;���YcǍ�G��F����\�Y:�`�FN��/#���ul��s)7�"��� /c^̍��ӱor�q�u�	��ABf �s�ѽ������s�M��d�:ڂ�A��!|�A9���.@݄27�"����{^��{����Vp�{�2v��x��ߥ�~��Ϸ��<Iӛ��E=��Y+6v�C�#�ל=qp������(���8�S��W�Y:�w�^ѵ*����0�#uyx�A8|�9��9�#�I�x����T�(@v��wT��g'��p8<BcA��!������\n�$�R�
'#�ێz��뱵d���y��7�f�V��k����8�Ɛ��Ax���X�}��j�۶��!�~��}��#�9��V�8t��d"3���\���g*0��l{z4���y�y�g7,�\�5��g��X��IWWBͿ���oB�و#�
 ���"�֩�&;9�El�yp�\���x���fE}�F/�Z�"��6�jTf���ы���1
��n�W��u��`�� ��D5�]��U	���	̈́Fbp�b�2���L2B�:��ܼ�s��m	�^���q�/���� �E.�:��d��*T����f;��4��q�M��W�.�v�~��=�_dc|�署�!·A�r�.vA}��j�r���s��������ى�7W�=ot��'8{f����V�8���}i�����}79�m(��&u9�Nۅcf�j6%X[[ZPC��]@�ś��9�|^0}��ǔ�B�;�����LZ2�{(Zr,m��qy�Ҁu�ՓN������>~���o��%�ڡG�q��>�F'q��܆��^Ry�;���y��ٳ���/��z)���1�-wg�%�TÉZ6D��tɀ���
f�h�r����F���X�[9��5ځaL�joz�G�Ӽg�36�d�MԺ���::�He"�-zn����F��/6�f�W�V�<js���5n��~vl�>ޘ�ؔ�����k�b�E�Ǻ��t�wu��nT���GXZ7g(�*{|���m�������6F����y��DS�Ҷ�t���LMK����,�E߳�+�e�ə���ݝ6������;�v{�n9��g��X|�Nxy7����Į}���n��&�"�����wo�����V�P���'�H>��5|�M:C]�ܯ��]�4�/{�.r�#c}N�|o�N
B%N�79"
���:&��gCaխ���z��	ѝM	o��&9;D�S\�A9�su��c��q�h���n�5	A��1�\�1l��ʁ�[0�'R�n�<���I����^�$M��:}�]����B�7Ox�}��s����	>�l�w��=p���^bIq�!�'<�q6��8�H6��9G-��Xmckrf�s3mħ'#6vA�۬#�\g`[Yr!Ĕt9��)p�9�X$��D�����m�K�(���\�Z�ɕ�ql�γ��e��q�ͭ�gc��8�vݒQ�ծtq�u3s�m�C�8���tt���9mn6�gg ��v�f��Zs��-��ge��I)�r$e��6�[g6�!�k1m���8�n,�ٍJ@N	%p�Zt���-� D�q(JCmD�M��e����ۉ,��s�cQmc��q�"P$�k.s��B ���H����;;�P��wvY,��
@GNvn'H���Rrt�9�TNڶ��h�		�@'n�8��[,�C��w���L� ]��1i�*�s&����OI�卵��G����Pݰ�e�{���5Ҽ�&V \��]�}h.ܙ���/��b�B��U�hU�mDU�%e3nc-t(�eG=O�v��CƐG83Цs�'f�*ܼ���n�u���g�������c�L"�5.�ͭ��, qq���5K�PXYlV��[���j4���5��n!�e��\j�	i,�z�X1cR8T�V���OLn`_Ey��

��$#�
�i�ljMjk����j@�R�)�`Bh�i-��R[��u.p�\����n�ƪB�aP,�4n�7��X\+`Z䋶#�te&n��s�|Ot�U;\dϬk�g�h��O�4��j�v� ���6�[�vK���q�v+��S�y�����D����b:b�Jm�Ӫ�nYv!6����D�����Q���=�����+1z��`�B:�I�&
����A�R�g�e�����o)<���LNK5��Ny��5�m��x���1��:��d�s
g���׈XUֱ�k[jq����ҹ��7aИJe���M��ea���
��pY�s�i�5HЛ���`���6[�m�@�B:#�2�&�L8G����ض�.�u�l�$��mm�0���-#3G5�y;ZN:��a�;3�c=�����`;n��A@ۓl!{<�18,�V�N�B��ZN^�=gr�t�n�.L�63Ma����-���|ybݮ��;�,��LŚA�Q#£e�s�W\�jV-)s`���1��&, ܵ5ZJ�YAx�x3���6�8$����K�y,6�,i�a��vt��c9���B<�ye�Bv�����c��Iw}��~����*�rbCh;31ͺ�3��u�ĵ�k�:�+����mXV���l�{D�fkw:�y�s�tTk`��:��q�n�:�`�N61���8K"���N�GE.��.�ȱ�g���g2������@U�X����c0��f덪��Ѱ�U.���&+n�J����.u��p���u�S�ć\�0ǥݨ����S�F�&80�]X��jlE]ZA����zqPW��s�h5�Q��"�8��2���N��Í��cvN::��rT��u��-����Q-�8�S[�fqv�*�ʢ�b+�+q�f)�~���OI=�bۦB�r@ޝ�2r�\�sq�Cm�kn�n��h�������D��-���#�G[�{�[/s"��"��j�`��̳Da��@��!��'2�/nԑ$n��@ւ�M>���3/-֨(��t"��Gdm����uƑ�:B ���Ȣ�0����Tn��������x�hMr�l"�#1/�ÅGn9���L0A��⏳!{�Vv�_K츺���]��l��ؼ���z%1��B ��!3#ّD� fmm֗���,��詘���
�r���j����^ ���
 �ȥz;c]'q��z[FT�Q��IR�P���p�h6�-�KB\I[h�Zi@�T����C�B � �d A��}���n^u��Ǌ���yzV�֮��V\P ������b�
 ��B#F���f^�թQ��'欞����f^]	�KefG�c�9����sn]�����{_5��f˔2&�f��ӂD!ٶiR�n�ȧ��h�&4�ҁ���<�펾��quqȻ�6x�E���;;_,B��"2א'�ً�����AӘ��v�ƪcwy�S�����T(�	����A�9���HoWe�:�j]%�b�B�彼��n^g	�Ǌ���	��DA��S��q>�/c��d
 ��@�3�#��̉;P������}�Q��E�y{:<�A�G2=�Jj��yv��=��I(@��*�^��X�n^3n3�DF���ŕ���0Mc���@���A�^^#1�b
"�������^[�P�q(���[��0�=K��Q�d{2���G�Y�����{�8|�{wy�8yw��n8��
��[^x����2N9~Y(#5An��9��2&"	Ф<����ƾR�%F�e��%V��8�lwL���� o����ylu��'^�{Fu��cd�A�S{W��+��w��*�/s"�7qȻ���� ��md A�|�Z�X7����8����Z��Պ"�n�O]���
	��B����!x����)�ְO��X�Ȟ;d�'W��=籹W�<�q7�@�[�����^#1a3���1�����n:u���k��G��-���v�ZT��q&`H&B�TH�N �]G��̀�d-yY���>̋���"�Y1�����a��B�1xfR�B^tE�g�ؙ����+�ۏ/f�ٵ��k���u���G�����ny�[s#j�&����*Z'9e�9Wr�?hQ�ݵ/�;���8<�q5�r[@x�3(/f@G2 ���m�[T�qd�9� ��^Vwr�O�"�7qȻ��9�=��a)��W5т[s ��q'�v0'$"�d����ِ�j�vT �2ZX�`ˊ��ܼ��<*u0�q��K�J̵)H�w! A�^@�̊ �/̠�o��1��/���5���[�P�p ������@�B�y�O�ҙKN�(��H:�XKi�b�RiXA%���6�0�I���O�ߗ����7��>�^Cws��n]����m\�Vs�X�˞��@����/���A2wv�V��@7Ї9�}�}Ӷ����B��G��>׳#f�Iv���s��Kݐ�ً����b�p�iN�ɬ}���w��T(��	���OּYl�f���#�!��#1yy��c�w�/4Um\����R{�O`��<����,��8�Zs�^0	����ȡ�/��vt�s�л��:<�>�G2و� �w� ʃ�L�=![�)����힯�K��=��)n^z2�6�X6]	1
d�]�끈��l�VK�}��zT=���E�QL�&����n��!�.;Tm�-uį�:��C�m�
�7 �l{���M!u�3`:ہNy�vS�{ct�+M��:�;0��7n蠐3pѐ,��u�t�����ړ<�<�&���xu�"�:�����z�'�r=�o	tv�e�D����-���lG!��/F� 3��ct-lrpnu�qAq˂�)y��[��7�[i3Bn��%	�ZаR�˒9�'��=d�U� ���q��_/"3#�1c��{��w���ꂏ5o:���{mt��'2#1�!�9���w@�U4�v�c�w��^h��
�z�8���N��۳�y��:h����bQ��i�&�JO��Y��O�qsޛ�B！8x�A� s#�#@�Ă���j�D^�D�0��<^^9�#�٫��{�X�f
<A�>��5$��e}�ew0��~n"~���b<x���� �B�ݚ��VXѮ7��y��f���w�&�<����� ��s��s=����(JT)D(A�q&n��e�x�ω�eָ0ִ6h��<<>C����#��Z�7���jԹw��e�B���MM<�f�`}8��9B#12=e�\�wv{o��:ӷS�(���Pn��lWZ���M{t���hD���s��H�#�f�pw����Nz�V�z����d�g8����Ogf��s]��c��(����
�n1�`������gو#���!�u�:��FfFp���m=����.0�Fdy{1�p�@�3�Ъ���<|�̅�o�_9�.i��|�����nN��+��y\w�.4��Ad"F���[y�*�Kg�r�4����%�ټw�p5����>�s"�f-��-��VjX�4��uv��l������i��I�͠B����Y�a��L��7&�!Gb�dz�0����1���/47[AOx!9}<��$�dy���3�\Nr�<n"�i����廫�|��۰�ok��ΩKU;��_ |h��/�#r�8k�g�!x�����F3)x����dAI/��^ �:A�ü[�CG�"��M�m�Y���њ�3�B��)a���>|���E[v6�L.�]�.R2�N^���C�;]���ݜ�{PQ�A��e<x؈�bs�&�9��}� `���"�A|��+�a���w��
��/)�S�z��J�-���zޠ�(�d"3#�p�,���"ߦ��unn�k��qS�P��	�� E�{2(���d��;��w�ՊKr)e�{#j]���r��g�u�hS�"벖��,�:1��hq���B#1/���ۚ4|μݜ�{PQ�)��ƕ�h��E\t�� ���� ���0�k{��E>�TY9�+��7����t��ƌ��D]�VG7U����h#g
{��و/8Q�G9�ξ�of����k��qS�PˁƏ/ W�d ABf$2XҾ�nvT����dt�s@��^�������ڂ���u�'�����>/6Ƀ;����q�7}]8�7�d@��I�Ż�S���V�Z�5���,�����vzoU��K���yt @��'�>x�"�ڸ'9E�ǈ\�,��(��u+��Sw4�4s�j���[�m1���Aq� Fb�����E��M���3�~��V�0����]�u��Oal�����۔���]f����Տ�{;�>�t�� p�^>̄#wm���R�^���Y�;�4��>z��ABf@@�B�sg`�[!8��3���4s;��r��AG�&�[AEi|��ZspV�X(����j�dW�9�����OJc���k����^VЙ���D�Ȍ���b���NH0�[��9��p(Ãݴޞ�EK��z�_ A�� B�r�>�A��Bs�"3�2=��Fe]L�I��8�'��h"����ֽ�y�Q0}E�̀9����FT��6}�i�\�M
�ޛcG�^���FȚ)�[���n�7SU��(�;�L�cd	l���+r/V��]�χ�����kMJR��`푸��Ɔ�s(,�3i/qx
��P�7�5;�nCq��11ˮ�F_\0��7`�ٷ/�Vz䎲���X��'P�.�4��G��:-t��dIBSB��n(�S�`�:{yƷ7=L��͈��7D.����we�ԴX\�й�L���=t6�NNN���N؜m�u��k�t������� a�}>|���O�ZF�Uܱ��F�<ӦyG��h6���mM���I�K<h<�����h{����7:�g��p���m
\�n��{-ժ����	���yx� �̀�A9���FF��/Mu��\&�v����9�ԺS�P�� |k�ȃ��9�����H!oX���At"b�f//�#�5X��R׼�v���ڃ'��Dm�
s!3B$b�3+a-(��R��Q�!�7:�Oi���t�m�Q����7��{�Q2:���&@������(Nd"b�}v�����|���{c�Tp�-N�C+� ��"�=��FF-�X�\1������bQe����a��iv��cI�e���X���Fr�МGg���y� fP^9� g��th�gwǙ�Ot]���3n,r�FΔiC-8�b�xw�v ����#=2[Y	�8t�	�usa�9l*�xbQ��"ob;/	ɀ��u8k�ؒ�F�bm�ڳSf�Cq��ٗ��\g/r�ۅ�C!>�g'��3�rc6��o�����O{W�]E�笱�U��r�;F<�=�s*�x���M����F�;f�qN�C*='Hx�`����1�f,td��t�30`g�x�/K�]�G3{���6��� �B"�(Ԟ��BSJ �ҼA �BjX>Q�`�b���~����S�s�W�s\�ژ͡k���<�^#1 �s5��kp�l�32�H� ���A�[�;nQ���Y���4�[A��%��1�]��D3�8��#�U�y��â�Y��S�P���N�.W�ȴh���!<P��ыZqJ8���k�=Մo�ۏg@�=N�t���v� ��A7Ё[^Æ���{��:��]�שi�Qc�U���'���7�J�z������6��n�;:Ne��0��[2w��d7�*��a��-�@�K�or��`��|��$�w�]��򅂱ů6L'ݯ��`w����C���w�}���?k�KG��d�+��s��;��!��:��}3z?m��@V�9��'xT����|[!�;S�VNͶ�[�M�B£����R�C�Ã��OY�i�:�պ
�[���8�dX�-N����c0��>�3w�<u��7�	�T-�Ӹ������/�%L=��V	qϐn)S�v}�g���e��b�n��ه�H� �{��������E&�\|�H/{�<�}�ݯ��,8�y�'+��^�}������8q�A�W=-kO�m[���=��.�߫�}�vn�/O!��h��.��F�v��bvW�޳{,�31����i�}7��3=����Ok����/t��կD�h��*��oKuWr���ۉ��˹�{���;^�þ��<��o�~��3U�ϵ�H�z�丼*��}��|�>�亓�gf�'j]�A���=\A�V�j��xO'��=vLG=9MAj��/np�O�}��O"�
������vgsZ�����VA�x��D.�n{g���l���}�t��t�ü�S��\�4n=2_b�H�j�ۊ �$h�@��B�5��_mұ��鏱�=S��3�=���b2ř���#�Y��y��Ч�f�S��'�Җo�3��q9�y�
�Qvv��]��Nf�QlU����-a�I�> ����$��m�FX���C�9�!̻$ݡ%�Q'۹m���h���;'" p�$�"�m��v�9��8��V�a8�E$�'8p��;�Î&�3�JD�9 �e�JAm��:��r\���e�s�tr�)ʹH �\�$rrA8R�ci��B�D�q�r	;�$�$I)�jm�9.IH�@Y�G89�H�N�9"(I���;.m�۳�[ev֜rA��	���$B$�&X�s��ݓ�P)G
S���w8�k����m���9G$p��9[i�7vؒ��.��� ��ۭ�NKn�h�rS3�i�)���m�9DN�rqG$�#���8Qqd@G!�r��w qv`۴�gbS�K7:��$�kYgB9qȂ �$l��Y)��枪���w�t/C�!�C1>� �PLlG<E��φ~X����]��O=f�b�z�� ���Kb��F:F�qǗ�4�Fd{2(FF�̵�B�J�*�?Pz��7�w����q�or��G��8p�����������Cϟ#���,ks���6ܽ�0����z3ݸ1��
]�a1*��l�x|&�#qdyda�}ג��gM8�9�-r+����qd����A�
s!��3�57��uLh�G��xB�z����nR�״&�h�^ �dd�鼙B��2U��r0��K�1
����r���N��&k��ݽ�8x�o�3�|(�-?Zp�a��/���DqW ��A�F�Nw^J��Κ/d�ȵ�@����Hk�ިH�X��ᤶ<�E�Io�f��RL��/�޻ny�8��k�i�v�\
�u�xF��ft�]��*�(���1�g� �}ܽ�|s!b�&2"�_(��в�'}�ƻ�F�N��7�G�^ �s!x�20��\!����w��sͯ��&x0J�Z�)�њh͍K1����XK�:�4�e��E�~��<�wBn��/x�.i�n�5���m�܃��1t��c�f�ŐD��+�s!��� ��
M��%���?�@���.�����gM�qȵ�t A0�����F�<����v�����C֯������X���:$����w�G&N��u�<Bx�9��da���5t�
جbT .4�F��㘂.i�n�5�v-�or}���H��3�Ԋ�A ��Fdp�f �̈�St��!<9��]���9�-r�t"� fR���s�Bۄc�M�f�\ l�m�ۛ�v�m�˨�<0��*Ƹu׽LP�h��3ۊz9G���{��}6,iyS��w��9HZtŸV�ug1��M���b0���u��X�����u��b�t[��K+�Q�xk3C��㗈w��4`�k�8ɒ�asTan����B�<�W<��y���O�mSe��݇@�3K-�`�E�"��z��]7�3�r�%�64'rg�����h���bQ��nԡ.�.K,n�sc����`�F�91���X��g��~��em\B�	��3]��M2M4U�4����q3<]a"�����Dsu.~���b#�S_fs�fl��Y��.��]�uWK��m�#>���F fR�2%^��5}YѤq���ZǦ���f�v"�:{�p��@�-��3�6g1<���@�5Q��t�A�^̊�#�'��%�؁}��v�ΑOD�ȥ�@��}����{1{Mv(�ױ�N��gP@��x@9��
�sJ��
Ȩ���p8<BOp��F���@�Ѥ"3�d"F���'g�ޕ9�|�K�{4D�n�]�Or �м6װ���y9��p�t;j7�B0P�x�I"�;5JN�sp�9�q����1�@`\G�L��z}E�4B �z�2�9F��up����Od�ȥ��.d�k$J�}3�T2��KِÅx�s!��.��l�X��f��Vѝ�&#�R�\���۫������|{^���������o8��P+�5~V*t]�f�k�<q`Ŋ��8<|�8C�r�4��p�,d�n	�@������E��9���h���/#�р�����Fb�\�YqQw��i���b�{�2=��!���fB ���ąEf�,��h {�f@{ǥ�[�sd;�7�)rx�@� u��F����@fE A�̏,��̋�:C{���3ùD�fi[��E����|$W@Dx�2<�s $���ҿ<�F���m��;k�#eۻR�pk�t��i��27	�2k��q(�������˸��@@�ļs�S���툻n^����ՅZ1zg�"�����2� A�gu����J��s�Q��y������:���W�)w��t/KË��[��n4��v����`����� ��D���.Κ��[�@�Dɀ�[�{*ij��r2��zߧ����*�`�rm�vK�WN1�+6�h)E[̝�1�����9�Kb���p4Qtrw7�"�x��A9��!AƤsV7a�v͸�;��z���ܩ��
]���n^������@��0m�j�X�n���3 "b�A{�����7���w|vt&u��� @9мC8BfG�,�����=�ϭ�6#���)M�L�j��8V�\���v����[	��X�����!�d"��8hA̅=ٽ�w��Ź�&�ú�N�m�˺���w!B#12X�+9�'G]�_�ƀ^M6�5:�[m��x����@��{qe�T�uyLI��@Y� s!x���F	��b�v`��[ԙז�hR�	΄A0��3^̀3"�F��\S鹚��%+��~ Π����!z.{sz!�wQ�spM���8�7��ڸ�S�0C��ob5h�o\���O�-B�5�H1��t4P6���rK�H^�N''R�;r���X6�d��*qe�M7����C-KJ���i���������z�\{�.�^5<��k����x��##�%�"/` Fdy s"E�k�����`�!y��U\�VAa���1�o�t��c`��§gzT���[�#��d�v·�K:���
\���*0��9٫�v���X��r�9E��*�1�*�X�"; ŬN��E8@|q�s��кGy�����W�@�]x�x�9�Ϧ�=Q;����i8@�s  Fb^#1
���m:�}u{��qf5��dp�Ё^�3"� �B��!}�i��0]@~�sc��@��5LM�p.5��� Ntx�7sWՉ�^�E4��̴��喬_��{.�7���v�-�t.��blf���t���9���zn�Jd!f�svC3�D�����<puPݯ�U�����)齘��.h0^�1"������l8C�&D(�#7w��]�)����7sƨ������=�Ƕ�q@nN7]&�tɮ����z�+�؝��݋bĎ�Ҋ��(��!+�j�l.,56�^Ж�*��yf
�[5)�AH�mJ�n������r6X&�Ze���c�GF�9-��W����� ��l����Q�Tح2][���#�/n��������� �z�a.M��*Mq��6bA��?}�g嘸66����l�6���G���v���y4M�Z��֍�\Ϫ��Qq9˗�A�F���w2q�k��ݝ�ob�Ԯ�DN �Ј'2f$#2"i�6#c �LQ̈́A7���b^w��1^Х�@�s�	y�o�����=^�܀��� � �Fd/Nd��#TU��q]#Clf�ج� +�"��@FF��A���My�b�5@{Ax���v�F�����y� ��^"�� L�tz�'����e AÄ�dW1}h���q��X�	��9�.v�L:���V/��6�_�̐q��+Aӻ�t����ܳ���Z��܄�s��m�,�t�v�Ӡ��"j�� ��B�����H��Ō��|��e�~��*��"��ȯFF���d D��kX�*��W� L]t�uQ��9���q����V�Ta��k�}�ꗸ��6(�㽞}ر���jד��o�T�c#h���n1ǵ���m�k����uyѳ�7мA�^Æ�^�\�1/ױ�U�8Ys^9�� da�$��"{r���	�h8�̺�< �B ���{2 �¼�Ҟ��+����;�#�
s!���#�I�܉�@�:BDAy�#;��Ǫ<���Df �9��9B����l���+�p4�����W}5���5�g��B��Åf@X�&jL�[͝���߮��V���V��)�³S9�PJF�g�
�ځ�KֵE����-�l����<�!]�-����iۺ�<�x�Y��Oj�<�#<n�^6l��� ��
�er�g�R�2h�A�js��GH�rb�ۑ5�h���D�\Y���+F:�F�o!FF��/��k��]��:*i�̠���o|�cB�c�j#.�QQK�U�1Ŏ�Ek:VӒZTW�IL��売�b�f����ˏh���Pq��#]]mV���F�A��"�(	̅�3��y������`�A��ۄA���n�s���u�&x Nt#転�Y�n�i;�@��{�^8p�����A8y�1,ޮ��n�R��zH�rm��*�z���׳"�9F��Q��V�tsF,`"veA9����A��f�K,�q�]��v�	���^p]��c'�8Ddq2=� =.�ll����uy���p1�,�;�\Ti��:hA̅�3�!���cVuu�`��,��oYk��	��;��3�������Z<dk<�����}Æ�ʰFs�X��q�����W9��O<�����/shU��&���ّDa��Fb�C5��h��6�H>����K�و"��퍗u�;��#p+�p7ЈТ��7�FuZ�bճu�0��3}x�Y]�48�p�{�i��g��ݔ-�0�DS�l���wE��vY*�P')�U0���'!<�fP@f@^ �1{2�o�X�C���!�x�z���m<w[Bf=n;�^@@����Sh~����<�����b����y���5$�u�I�	:�RNֻ�34mlx�Xw�,�{��{q̏/�@r����pV-��*��S��H�i��A���@�s #��_ZP�}zQüf�p��|3/N%�퍚��[���W �B �|�fGQ�ٻ�l/�#� �1{2(��Ǫhe�}���f�m��m<˭�3�l/Ay��^#1��Z�Mէ��,]
Eǭ��9���2����zGb�{�B�����X�U;�n�-+��gEOt�A{2 ��3.�F����r��6k+��%�-a\q��/o�^fB>̉���7Sdt�Fj	��b�o\7V<Q�W�&r�_�g_��o��eLw��(s˔��a|��~���<o�%	*�V��[�r��{k�o�{:�mA!�S*�(<��������wQ�����@��/�O�V���K�S��-M]8��	V�7wQݽ���������	�v(W��f77��YcBOHYm�؊�b��j�b QB�wCl6��pf=��ȽMaʱ-6��v4�����`�E�V���ޮӔ��a�Z���8I�<sg�ȫ��=������(�Kp�����Tʹ��h�0�L�o����o��s9yqA~�����Y��$f�Մ����GQ��V�>���zHK�.THt�F$SL�sZe����ʔ����>}9][�� q
�=��O���|?{�U6(���C`�?��aM~���JlB7W��U�c^wbX�|�7ݵ�W�|�ԛb���eW�ѯ{4�G��|�����m�}N̊=ɻ{έ����Dٸ����	@՘�R36�8Oa�D�,庻��mf�CZ}8�ND���cvh�h�g6lͷs��ʵ��MU��*;���n���l͜D���7t���W_W޼������`r�Us3n]`o"�!}s6��d^�ӓ��R�W�1-��v�J��W��D��ʎ{_vi�:n��$y�-g	�{��>�ֆ��3{σ� ��o�[�W4�r���ktTv��~ǩ����汇���/=ϰ׬*��a�޷-��g�^���;��SXN^Aݍ����[�`}��0�T̍�M�N���ڄ�`�A�	6jE!q�t%�e�n]�E$"uNIYvp��h��	;n�r��r��8�Yf�6���$J�8���L�d�GgI�Nu��-����9˃��(�v��j'��'�BpI$����e�"Gq!D@8rp��3m[-�um�dG��D� �$�'�.An�6��&�q#n������.8 �G��D�9$�#�*ID�I�i�9ȇIC�NP�9$�tQNvX\GA�r\P㙕��YaA$���p	9 6�9�-�n��X!�ڵ����wfDRA�v�(�kp��%rv��Tq��Q�"DGI��N$���u��D��C���)Δ�!�p>�5����S�2�ffse�&���n�v|������v�:�I�;j���u&ۜ�㎺9����"t�^���͔ٹ��� f\�M�����K��xR	�. 5�M5��<�j]`m:�Y�ǆ���phi����֒���l	��[�{C�0�� �a�99��Ɓ�l�n�y�p���b��*fv���tGi�v�=Y�7^J��W&�:��l�1zg�bq���5�� g�m�qdϝ#``h���B��f�YF��
�:�ZeX �z�K�\Wi�.���e�Q�XENC���vR�p^{�C��2�X�S'm:��Յ���l��c>��6�;;�yҖ��<<`�mv57�yʧݽ�r��X2c����m��-3��W����뤐쑧�c\�e��JV���8L<�{ko9�ݤ�(:�l6��4�Ň]s�lh�'��̇V�RZJ�F�0�gK�Յ1�.
�Z2�Yl
B.���z�Ź��m��E� K��0XW��t+[])�X����Lm�s��j�^[��M��3���<���<6*���l�+L+�te�W��.{l*�.6X뵮[��xY�_h�ٷ��ێ����Z磚kn^�:�s��#���F"��Σ%ؔq]�s�]���F���"��0+P����*���G�W�v�v3��k��=Ⱥ8��^\�I�5�'Λ��7�|@���������9q��qɌg|}���v��Fг��;��Jfzڎ��Ɛ`m̸)
6�1ϝ�봼!ste�����;�L�c�����ɷ<v�;�059�27gb5Q�\�MX�����H��Mm�\-�]gr���:L�g��>�ؚ<Uv�ڌ�R���Q�0Y�$M5���f�]s�»8�����h���t�k����0�gN�N��l#Y�_=n�{��7�ڼdty���>�g9�jp�׶E��"��2�H���n3�g.I�|���g��帱�G����Y�x-ٙ1�b@�5��������:97pp���k(�m�1�&磷*87(���n����R��{z݄�&�p9VS�Z�u��=�>�	��9�y��ޮ�!�w���NN���jJ��w.�Q����m���˳��\���::]/P/k�5q�ز���ڐm������f6�L�l:.�ԫ+4��ݴ�X�B�K.5�결���+g���El��A�D��!v�v�_	�r�]m	�C�E��S�o_p�� ��!����#�
 �s!�VMJ�|���m4p�M�^jq��y
Ţ�6�_ A�� "��dF.6��蝍�8�D��7��9B#1㘆5���d��R���9���ܗx��g��/�8Q�2f ����keVᎤ���$���_B��B7v�wn_	�r�]m	����F.I�FOTg8Q2Gx���j�5�	̅�b�5
/v�徔A��7z��C��h�͡w�G�D[A s#�da���{٭]��V$L�F)RD]+E`ұ�Fm����if�|��Y�d�e�p�i1��i��!��� /��^ƪ�_Q�u��<㢧a�9���OG��E��/��s�����U���C���"ʱ��3�v��}t�r7x����I	�^;��ˎ��Gf죭m�ƫ�+:�w呄�!z7v��n_	�r�]m	�u�!�!3q���~ө�˜q�"��,�.q��r;�a���tb��ux�:�	�*�л� +�"���̅�	̀�́�������;Q���㘂'��5U��;����q�o��w�Zu4A�DeG�n�������9���o
T轝�=��&��n�hL��p�>/ "3#�وE?�����9'�i�S��v��8c>؞��b�kBT��:��]1L��.�v��x��@Nd&�>|!�k
���*�!^�����k/Tn'7E��\Dy�-9˹�U�*2�]aTC�@`�������|�e]��{�.����}}�_@^#23�h�����zLd F�7 /}�� �B�kK6o]���n�I�NU�s/u��R��`��y��ݷ�Ҥ.�.y�k
�w���x��
�)��_���bHǙ��d��G��g��Eլm��	��^̈́|�fG�b����h�y����^!�Ds!N����5�C��|�W@@��z���{|.�h3��'�Fbd '2f��W4���PNjs��MY�W��X���Ј���Fd A�̈]z����LA ��R����n�
��='EO�8�Xy����`
�WL�׫�,�����E�9��'2�O���g�X���<��t;Bp��$|w�"1��}��̀3#���G;0�(I�� �F×���',({�B�]m��d7�X�`5������D�3#�f!��ML^�Gk{�U�q5gh��˽bn=��|����'2#2�c=�{dh�#5{af@^�M����W���=�	͏iKBٞ�=���:s����ى'�֨��bX�o�-*�J����#���'��V��S�qe9`��p�x^��#�����z� ��D���#2/�nV
1�B|n�UOw�9�,D=͡W�] [�^9���d�;N�"6��u~O��x�,�!�!qI]F�M�,�����Tl�n�")0�A�|�
��gB�##���}���n���VzM��&�x��7{�;l�'AH t�@�s! Fb�G�;
�Daݰ��"�s��7o;\co'hLǭ��a��3jj����z�5�:hA�C1Åx�s"ʔ�%�G���}�-b!�m�G�@�-�fG��!x��kpdĺ�YH�l AB^��}���}���7�bݼ��&�x��k�[�Vt�@�qǳ(/a�1s"��E�����[oF�ga��m��	��q��@������"8�v��؜�H�rWu]�8�U�*ּ�u�UR���V�R'��k|M��/"�y�,�Bۭ�On�w���<`*n�w�~��u���;�7p��λ+`|�)+0��.1@Q&K��[5��Ōun��̠Zţ�hc%`��9�M�L榺e1�� �۫<����J�\��(B6�]�يɜ�xŻL�6���U�Bq�x�`ܺ��6��'Mr��tK���l�.��>{o�`��ñ�)Y�8H�)	�� FU�#�e��nоT#��-�v.�#bBXT����������\B<[��V3$��\��e���]Br�,CfP���xw􇯷��L{=���r�|��@��sh]�@���vc���D�;Ёp�Fb��B�# a��ۛ�s��K���m<1�}3��ޱ7&� ��Fd4Ҿ��x4�Bf�	  A�/�2��]���Sslc��3q����3��@�������^Æ���B#cF��A��A�^ӆ��d!�����0D=͡w�<@%UTF���w���Df �2�#Dfɽ|���籾�6�����S�1��޹6xA���b��dE�-����}Ϟ���غP2;fYr=�j�\݁�b�v;��2�(�Y��$]>Ϗ���&��M�Da�4�q}Y�f�y;Bg���S�`==��3�� nח�b�¼A2=::!��a�`�n���D�����ں��-�vL`��Q�v�қu}ѝ����;�^2���KN:�ˉ�팳q�cbz�0�*�2l�A{rǸ��I<3F�m�@�h��x�24É��ӱ�����'9ab?�V�+�dNr�9G5(����iv���D<��z���7Ё�\x�<�X�����Z�]n��nҀ �/r0����q}\�&��m	�u�L6��uV��\�=. M�x�����d A�/��1��D����^ՙ���	�oj��\��"� B�{2(f@2�Z4:&�d�hWL��Y׳#Ob�W��FË���&?����L�t�k�UM��ѮQ�w�b.r����s�Y���%O܌<�����w�Xx��9l_٬��ݖ'U�#�U�9p�����1�3-y�{C!��s��x����m	�^�\a�Ą.�w�P0�eN8@@�A���dOd��b
e���8d���cNbw�$\Djn�l�n�s��G++�T�]5ῇ�����y9�]i0�{��}�@ꞇS�qz���.{o�M��?�>�^̊��"3A�Ϊ&�gj,��!x���(}�x��FSw������@���M��sj,\�٢��Fb@�p����F���9�iM
q�����y�j<Ŵ&x/k�A�q� �K�f/Eٔ����ʒR�f��is��c�e�L��]�����j�]-=13
,���#Z�A9��M�>=����B�
�Vt�ْ̙��D�{v(���"3@�����R���l����Y�/����J��c2���&�x�o�F�Æk��1ˍhw�T"� O@Y�/�@���Q<�;��ܨ6����-UE��;Bg��C8B����1>�1p� ���VǬkA:@̎�/s�Ӳ`��͡s�!i�h�O:���v���뢱�S��n���w�Gs"�n=�h��_'���e
��1�����+:=����"~�������u��fW��,�r���%�s����Z�A�f ����*{���n���?|0	������?�֕���#<�[Bk��,BZ�-��˥4uM�y�0��{��@+66e�l���@�xLC�~�q��D��!�n�\��[w��&y�or���Ժ�0F��x���8p�9����R�M+W;R+po�l�^��<�z��= ����"�!/ /��R3t��mG:4�k��`�h���R�e�6y/z��S��e�v�ը��n��>��D��8@̏]�ʮ�gY�V������l/FFv�\��[w��&x |sax�ӱ.ٷ��*.ɷdH!�^#��>9����8z:5VEmA�;hOp�� �k;t�= Ӄ[��-r��׈/��8A����ɢ�`@��K�x��Bw��
���(=��]B���*��t]�֓v��1z����_�K9��շ�ɺ�7y���0I�3�Z��}67b�g��n�s��e-eK���Ҩbm��i�a�b̰K�n��3�L�Xۣ�l.���XOfN�;hJ��ƥ͆����8��Rqo<�f�lZ�r;.[M�ꌫ�cB��Dce����3v���F:��cQ�c��i	�1��\F�Ueg
��z��(n�㋛v���M.�)��^�7��*Z����>��gW�8mґs�����t�U 0�0���X�3>Ϗ�~�{Ow�4f%�3^����&:���m�x�j���L��y{�y�5�	̏fR8B ��[}�'!v���@�B:0�!�Z��'��-�s�&`p:���������y� �ާ�N?�,�����*��9�����= ӃZ�lZ������d"��#1.}ǳ�j��8�|��p�F��و!���LOGX�md�{����wƷw;�'K��d Fb���>�A����^7s +�!z)N����quݹ�< p�!�3+���/��AM��St�9�rnN�	�v<�8ܹ�quױ��SM��lv�I��X�ȃ�A�Vv�1��EC�v*7�p�q�4���ʃd��"��#1�d{���Q$�s��h�S"K��=w)�{ҧ��3�bǧ5zk�->{�������zl�8�����%�K`�g���;swi��^�,N�բ8��x����>��rbz8Ff<��f����ւ8p�����
˖/KD�,�����W���=��ˇ�Occ]��<v�Й���@�p�̏/f �p���̪�z��6�#|Flt�Ds!l�z��+�����v*8/a�#G^	Wc��fE��0�Fd{2(�ᑄ"3$�/�9���Z���d��pŘ��ݚ V�Fj�4A9�$���O/��O>�AvE�R��
��r�@\Nݗ�l鵻���уu�YOS{����h��2�Ä(s/�c����f;khL���GV������A@ޏW�^8p��d"%��33;`�<�G��p�NS���G#�I=۠j<B ��̂���K�������Ј9Bf �b=Sn�(�k)Ζs��6f�znػFx���C���^�>��x/G�*�;;�X���佛��kܓ=���b{$W��ڽ x�0^����+Y�pnu`S3�����{Q���	1]>ݧ�ػ̃<�x��d���-�������K�t�g���>Jo��8i���zo�f��]�$d�:�un��03n����eC��v�C��ݸ;V�z'�b�QS(�%7���k��6���Y�������h�G[ZX���M����ɔ��Jٍ�P;��3�M35�X��[��h��:ڹ!��X{�{�.�ʰz�6��^����X{=����K<$u��bG���`��5����J3٧���J���={��^1�W�Is�r���Z2�\F�Y�c�*}���3��ݺ�����͝��D�;Cv߳)fӭ�˼PIg34Tȏ{և��b�@�����Y��"�Gy��u{�b�w���	��{�}��K=��d����o��2ٞ��gi���}���n�f���6�x��>Ԏ9����n�8x�f�F�ǧF��k6�N� �I��s+nI�q�A���Uw����y���:r9�\v�9��1�x�+X���^��hܮi۞����5�O����hyz�r
=���A�燯����vxFzgx��!tu�{]�3T���������f���=�+6���g-(���ٝ�a�B�hy��O{T���{�&���o^�<�S�|��}n:����/��V ����]R*�$8�9�8$pN*"9pq�Ĝ����C���Bs[%Np)܂t���tQ��I9G$�RI���)m�q$
:�J�kP��Q!JNI�$NIq t�����t�q���\tqrI$���Jt�QB@�$p!qЉ8�� ��;R#�8Q�Ȕ��@s�	ã��gG$q�.Gq	 �HD�QD!.s��r�kr�t�:΄�G;-$9Nt�'q��AI2��.M�#��#����Nr��A�||O�0��f��F,Ǘ����8}������e6�R3�%�>v�9�呄(s/�yG;���v�Й�[��	F��:."�u,�Sm�a����d A�b�9�ޡR�wu�(мt��1�����ݺy!@G2<�0�Ў�u�v,PjQ&Q�D��S��rk�O>]l���x�����ƴe�hĳI��� |z�v0��^^#1:u�cFWǆ+���xh��.S[ܰ�؉e@G��A9��Fb^Ä"�b:��+b{��D�!GK��ҹ�]Fe6��O�l"q�"3�_HS��sA<Q0ZP����(y��O{�+/[$v���Lv�q[;�`��>x�2da2�^�U��T�}5��Q���a�́@9׸ډC�d^�������!�u��ꊃ����	p�t��2���,�:�w��:����I�d��h	G�Q���?A)N�<����`���k7K��� ����ְ|(�1Z�J���p��������]Fe6��O Ä́g@��j�g+��۞9Q�Da\Mh	ҳ�I�[C+,�V�Z�����y^{r�ڻ7A�%��������y��(fB�X���c�(w�[vpB�\�JAd�� ��:��#@���!.��!)��"HƂ��bV���J�/e��4xA��Cp�63(C*;C��To��^^��f �d A�FQ)�:/g�]n��y�r�n�2�[B��� � �@������E������a�Y�,�	̄m=|b;�C���۰��'���c:�UH��[B	�XXǜ���W�s�>k�׼�� �ͻ�q����y{/ ��@�4Åx�dU�� ��v�v�sx�`5K�+�=��`��S�յ��wn DB}�or0��O��Ĩ9Uj:bӾ.
���Jc�� T�Y�T��μB�Ǫ[�.Ί0�f�2�-3(]�Y��
�-%���tv]V�r6;��t\���W�/bځ����8IT~�B�x�nu��n�	�Ns���kn6���9·�1+��̙���^�Ss�0�P�Ղ���Ii]Ƽ���rKS��iJ
��C1�t��T�{p�]p�Fmx�K3{i�p�4,�l�Y��n�H2ą�f?���jC[��ۂM��F�8{R�"�[�K�6��P�K�MYG��?y{��[Ax�B ��!ݭ�}��&n3)��<���t�`�Q�#D>�,��ÅfG���[FV��(�6"��|T>��En�݂�p�x����o��QV�
�B ���@���"3��Ce�
�nV]��9���y{/q��8�^�9��Fb�ʲf[e�`6��"F����������m
����&g)��^�^%���!�e�!�U3 #���|19=�m�"��国����$�)�m�+��!x���̄ da�>԰�viWA�#`\��������k2`ٚ,%��ÔU�űCf�0�;K`fZ��p�vX��jY��Zs�\Nr��u޲\��r�^^��G�h<>������:h|s!3�����U]U���I~�{�����;�;*oa�kw
A�SkJze�����]Nn��Z�Yb�]��=��z����Nv��48�BYdw)���s�&�d�[B��p�BfNk�JZ�Y�ër=���>�sa3 #��̌��������[��-iI�Sڭ��@��� ������ fR�.������"�@܂��b�^�q=��/Sf�����]R�T�\������3 P9�!ͩ�������٬����ɱ�-��S�� ��8�Z�֜����}��V���w7�PUew8\PH�00GUQ�4�M��-&f�6Ua<����=��#2<�̅�}ۏ��	�K٭��9�ͣ[�9�`��8��!i�2���-(`���2y�n��7P^s������9���0�8��<�4��9�o�nWf���=���x�3G2<�s u��Xo�n�6��)˔MVɛ�����{1GƉ*NQ�^*�2H�x�u��{Y�U�=l��v�n��z��a{��o7V�ɱ�-��S�[�"�#1 �|3@��DT���늁�P��#�>̈�ݷ���	�S[�`�{ r":3=:Vg3LW�u k�Df �2<�d��pX��r����!�ɧ���z�/S�
��hȠA9��v{���O޷�.�Xi,����*���xp�M�]G�=���l�q��>�^{Є�嘟�ٌ�@�s '�[z�;tb��:�Щ�6{Vuʒ�n"A����  p�Gِ��"璲�6B2t��p��ۏ���	�;[�`� |l�b�2(��vFMow
��A�@����^#1
�n;�c�!�&.�Oh8���VV��>��#Z�¼A9���!�3X��'��"Ȭ��݄Ä/ڭ�}�1^�klT��p�*jx뭅���wE��׉�;9V)�4�"����8]HjOL�~���X�����+=O&h��hFҸ����]��n�:�w`�w �sPGA�̏f@��r���}�{�t�)�U�x����۰g��6x��b�@�8Dv﷜i�\::�4h�ubXi[�`��M^,���l���y1g�Z �2`H
L���	�~�!�Y�|�^�c�7�+V:�ݛa�i1�d������̏ff^��ۃל��Nzv�z;X�xru����cřC��r�u�ݯ �ffP�4�|1��$�۵cw �N1�ݹ<+9xfFd{3d	\v֫�Cz��K�G������ct���*5����yl]uA�Jy=Au�n@���ٙ�Z��|VE�sӗ۰���Ó��c�n<1���Ùb�P�}t�sW�k���ݠq>��ǆy�0i��ȼ�6�E�-���lؐ�~�P���;�� ��
�?xj`!v��G��;=�� ������5�욧�g2�b����^�y��O�����αƲ.��q+��ӹ%.���@�y�f�ݨ�n�
�P�3C48��u`nxiN��R��j3�;���6�NFˤ�p���-�֯Q3�&Rg����r�u�A;uԢ��p��h�k6
�v�L%����iue�Ip����7�aϩ���~�3 �`Lg7U%줮D���I�Ob�On��0c�L�%I�|:�ٱ��fG�����#����;|�ս�C��[�=��^̏�{��\��fe��6sp�+!giY�{��}��en��5��#u�����������197/ss�2&��=�?��~�my�i�ڳ�E ;����7�ّ�y���rb3�p9{�xVr�:����<���<�;�̀3#٘�3(��ڇ�2'F�Td�0a�Yzs^.�tz�3+2��9=�y�m�(���* $�u����ó�6,mX�TꍶK�rd��%�OO����3�[��������َ��7��}{�|7r� fb f@�\�bM4^���/����c���8z��zmc'5����B�[����[A�P�{;1q��v.��5"�E�Ofd��E�%�֝i�P�fT^u�xn@����ne%�0��՜��f������;Z��������DlƮmn�+�Y�s^.��������f:��;Xt�W�a�̡��oGs�'���=�k�V�?����?S�m�2�i̶�7
�?K�3�Ms�̮R���<g!y�s-�7���7{��<"���ù�a�Mù�m�;Z��qR,Զl�l]vbT3˥�3V���������W���>��\g+R�ƌ��� gr2 ́����9r�L�k��y n���ݽ����6�7d����ɾ�wg����q���Z��o��y��V�j6������m���h���]�̋ݾ�y��Y�/���h��zv���X(�8�5�Px��[&|����.���}�v���f�n��,9�t{՜�y�ᙋ2��*
�_�HS��n3#���
��'���v�yL�Y��K$�4�y�ᙋ�23:�8�ޞ��jS�����B�����<C2ewm�t���`��� H����r��fZgLY��䕚(!mf�0Ѳ垷���nFf/f@�o����zQa�k��N�	�1�K�}��8�m���ܿ��Ǩ�Ws����h;��j���+�	��m�6�n8�G����U�i�Nff�J�}�"XwU}��7B�cvO�r�Yi̶����G��667�x�@fo�Fm`��-��rxzy�k&�ꝑ=
��DfSsKg1���(Г"�.2�����;����j�Ԧd[�9�Jcr�䕆a.p�f�p��j]�1Þ�Zs-9�mY�����B����ࣁ�<�P�l�z� ��fb�}��>��η�o�.ιa��y5��!���`��c�Qg++�r�D��#(̉D��/P��d�3Ng�GvW��s��%��X�W{2c�o�l{231�m��`mj��ݡ��}0q��r{��y3X��w�t��޵�z=��fG�eNu[�ӝ��WK�ࡃ�5֡Zپ��/��@f@̀�n�j��X�MTܠ��{3Ng�GvW��3�vOx[��|��t`gw^�Z��op���3 ffc�_q԰��!Wc� ���w�u�/#ّ�33�{��I��!!I� B��BB����	'�H@��$�	'�d��	'�H@��	!I��!!I��IO���$쐐�$�!!I���$� IO��RBB��I	O���$�@IO���$���$���
�2��QI� ˞�����9�>���`                @                    n��D����� PQ@
(P�@��(�@�(�B�T T�*JE	H @��P�&��Q%��RT(���B R�TT�	D
)EI��*U%
�Q���TD�RJ�EJ�UQ"���  w$�T���@
��Y�tҀ�]��j�gUJ��(������(��wG��y�����Sց�x�K=
���TkA�ԮBI$%� �`>��n`t�z$��AU�cTꕽ�z�W��o{ޯ@��E<�{���j�;���Wz��4ck�t�
@I#� ���RJ�(��U)%Iy�>���-V���⡧�a�%�Q���E{�T�6xڅ\�.�b�ۢ�ՙ�g^�Zj������`�S�` 3� �� �   �� @^�AA@ �� ^ A@��6��� � {���z�� t 6�UV A@-���+w��Z�5w�Q��6�t"�E(��@�  �� �*BJ�����@)�֝��٪�\`�vӽ�J=�ރ�ڗy(ޥT��s�3T�z��O{��G;R��y(��z���{P���%*�P   �=�u}������]��F�U��� ��o`A� ��\ g����� � 8U(*��H��  �ꐑ
IR�
�AAUUx Z�����z #v V�EI� �z ;� r 2;� 8��AX 3�� w�QB�   `����[�I\ ���:�G .�!��  �9 0R���
��  <�PJ���JIUJPP��� 2@݀rd (�X��Q� r�7`��AW $:���(@P�O   >ü�b7� ;�(N dr�4�� �:�+= 3���)������ɠt���̕)P  ��IJR� �"~�U)�)P   �d�R�  )��*�S@�2 	5m
J�~Jz#51?������}�������H�5ғ�q��d~�1q̫�_����$���BB��BC��$��HH@��!!H�����w�+�����ޜԱg�S@r1�Q�2�X79�����A�0e=�Z�τ�b�\mጼSy�2[�:k������^�4R�v̫�=_�x��q�V�j��`"닚Q��9��:�NU�b#;��x�m�7���v0:Z%�s���l�F ƭ4\B�A��x�O�Ʀ��Vtgz.ֱ�.�a�5��{0�x+�.�5Ʉ�#Z+�m��Β�9�ܴ��Ne!vwVY�A�0*���Ȣ�sN�� �ơ#K�Owr����V�(�'�x*�A�c�)�;�N;��{	���i')�S�";y�X`ʮ�1(�!�����ɧ�7��z������p n��|����� xb��	�ܷ!i[n�n蝟�z8����o5g^��N�b��]���p;�ey���1�����4��[�G�[V�D&�[:ҷ:���L��4%���j����;�+��[ӯT��l��V�y̢wW��Jy����[��g�$�Pig2��y�ϸG���) 	�n�Aq��w"ĵۻ�vEN-x�>��e�!��b���_e����Ƶ�������l[[�r�S�`�/C$�����JҔ�z�����ۼUʈ׺�,%���;���h	��KN5Y7��n�ryt�W�՜��I7j�:��zXc�!�wC��q&V-�%�L�:�&/U k'lH�.�;_9:]ت��RL%��6��P"6:{mu'�^j��lx��{2��ōđ��l�f�~�7Z�Rb*����N�c��C�r2ݶ��K#]��-$�cӳJ��z�Y�����be���v���:N�=�5|�u�bٝ�ׇ�"�^e�y-��1ǎvv�?s��|8�	jr�q��у�W(� �[4�g4��'�L�QZ�ݑ����d�Fj�� ^��]+5C��Y���-�Cv�{n�;�ĆP^X���ٗ�ט�	�H\������3B\jiq}' ��q9�b��E���h���؅cF�x:��n�d8ї`����5�wnk�H��͇wl�a�qUz:�-����᛫���^M�Aē�rj#ףG~;#qh��'��LZI�݊#K�-�Đ���Y�.@su��3g���w��`����w�P�n)�`�^j�wcRh��X�CV<�t�� "��h��؂�fWs�M)٩��E���hY�P�+"ը]�,��8A�v�V��v����Y�,m���K�N�~Y��H����k6X��ـ\q�������QM�N���AƤC�a����	guJ���U![V;(�W���+L����:�Üo-P�Oa85�5�]�������������,�k��q�m')x��T%��7��-�"Zam�"��kN=�s�uk�����8ك|8Z��H��gI�7dwz�r,��a�ygB�z�����H�ߖU�KӍv�+dd��ҩ�˦q�qzu�ԅ��`��{V�ۓ�^p)��@$k8��(��Ɍ�l��!���x��f�8�rq�9,�N��sj��s����`\-p�����p9�k\o;P���\���Vv����D�����E�^h.Y19�z�']�25�(�e�2��"j���ID�Cg�m�#לx�cX�IU�]����1�)Q�r��p�tx���Ad݉,EQ�ɛ�:ƍ5�w&�혮,��
�k����Z�m��6��������T;�|9D� B(�6��� 4'<��xe��[�	'��K�;���JuE�I�	$�XV��+@;�p��B��q:Lɺ�frܰ>2>�cF��B������.�An>�f�ܤp�����!&�nuOu��f���t5��$�zJ�:N���'!�a�;��]/۬��ۺ�v�p����.w+��ƉZ&r�-6������e�6�D5,�˻�G�\���ⶺ�b!�^��5hrL�0���~��p>p�ۭ�F�/w^�����hܜ��������prK�N'%��d5��{X$���5@EoP�C˽�Զ����]�q���5�&���\�\��KeOAH��ނ�h�����F�/]hl�3��E�0�Ѭ�Iʩ���"�1�� {��o�<�x�4\R �"1� 1�ܴ��;mݝ��sy��O�?�K�-w��-4�c�˼��8�g'�	�Q��������X���R秂�y�t�Eˮ��η�n�"�E[�mBq.��
��� ��r$>�r@ n���#��OY�����:d�B:�u�%b��/�2q���oY�=s�o���&��Z�i��{3Doo���c�x~�}�b}�J��7�ę�
�P��+���*Cj\z�����V��a��+4��S7i {{�͡��z^hI�:K`����'vt�x�n��Vc�̧���4��4�&2�5��;{Yx�:^{����C�;�t�0����}kg�):#��y� �����;�v����BU)�4mڤ02_B�����%(��]Q��|��c��>��uc�;V��Ʒx��X��c�4'_��Y�K�U�׆��6i̳��':��, c�ziz�cF.�3�CW=�X����[��Ո����S��J��N�k�Aر��:�K�����mc\wN�Be�����f��%O���Cw&I�-�Km��[�ǔ�'�=�i7���<�����"!�"�M�� nSk��3xqә2I�j�;�흽��vm�\PL+;��թ��/_Q��x�
����r��[����*�,���k0�:�����O�U;��=��S��g#�F�A�"'v�����ùlQ�5�`�C�`�ݽ=o@^�-�%�Mɦ$��9��f���~	���3;(з:f���xK�-�����-p�Wg:�.����R��5��hy�<#�ئ"��N����n�h�#�^{��	�9�B~���X��.�@���sǛ�r�7FP�㻺}Iټ�%R("zwt��}*\�w��,����6)��+�� 6�ovf�ø{��P˃s[y�Ma��[&�����Z����ڙ!<�W}�4��j[�<���{��L��t���'^waׯ`�|79� ؞vOn^1�6^���*�Ĵڲ�,�����Z_k��/d�C���(��td���-��4�	*8��S���w�9�3IZ��H�,��!�{���q�VN�pg
ź��9��x>�Y�m����z����1��GV%�;��czb![��uD�p>���y�f��3��x��K��Y�WT%�Ϝ�kOgV��U�7k��N�iˌf�Rт�vii��ev�Q��g��L�Lƣ�x���<gj�ޙ�^�=����������h�\�eL;�G'q�'6p�|�>��c�rV���0v��� ��:k�8H�Zt�BԜ�l��Q�p��˹��v�1���<�X󴑵U0�{�K�v*�`ۂ��7�@G[�}W1h~B3�Sr�������<��k{.L�� `{��fg̘ i=�m�5����X�죦�h�ھ��gtk�4 F>��A�n�����s����8�"��kN��u\�3�v�V���G+��w/��o`�x�� ���V�{"G��;n4S����]ɼ�VN��v�K����OO�-т�������cZA�<�������[�?��VS1�W(o�һ�)�uQ#���*spebn�c���gpA�s��A�k�gC�g4�n+c�KM�ڻ���W�=kKc]�	�Z��j��7q�lIDޚ��;������GE�����<��U���qc@&��3�M��� �s��%���	כ��rD�|�:˅�dr��nޭ.#�H�ՔW�]��O#Ir|�h���x��$�=x@9�n���7�q���^�V���Z��w�t�/��c��7^Y ��$�]�������:	/�������GôB����2�K	�d�|��i�ܻ4,)�:������v����7�,�L�{{�ާ8��5���qBpN��:�.�F�<^iطg��pq��{SSnk�]���X�f�zt���q�ݝ5�2oM����FƒJ��y�.8���w$k����Fw���nNM���sr�+��j�6t$�H��=�}o=ų�N�n=�w�IצE���mn.Rp�+��zɤc}�jL�٢�;]�k�*�]���I�`]h�w�{^�� �6a�oNU�B�7fF��`�����{�LFZ3�Wp7F^�Y�[�2]�pQ����ȀMP����Y'kQ�3�v��1]{wU7�܃a� ��u���\�^r=�}2�^�X毪���+F�˔�Wr[�����M��l�I���s,y1ګ�dw4v�o'��g)�	��P-��Ɂg^e���
�@����q����@h�%�!�C�Y�QN;�bD�An,���&U��t�p�u�З�k�5�!���
�d����<��0�|�9��!�D���y�Y�趪1�St�z��d�d��i�7.cy��̝7�42ݸ8̽�7�o5V=y>xwZZL(D�C^L��A���3�һE)�3F:���:�3˒ͻ�D�#u�ȧ�L�M�A���%�ӓ����z�|���j�5�wz���p���F�e�pzރ[b�{
��m)�i]��p�!��+�AǸ��KZ���:��tC���Kj�,���w3����{�>���5��s't��Э���\hQĮU���G��\kB�M�93f�Y��������nu�ɲ{�D��qV�c�9�/w
ᭁ��ʟՎw;l,�՚�U�����F��sn�W�)��������m;�>�oi�a�oDM�4M��rs��X[�r[�i'KI�zNB��sr�$�c%���w�3Esf1Np��{4�@��Ɇd��}�*#:�v���v���y5Y�U�	�JԪ�Ƹy�j���L1ob�ʰ=\��%�+t���A�nh����V���o-��rT� ֻ���A�7�e���+KŦUki���[��x�V���Hɫu&��xb����څn���ӭ��ttܯ0l8se�u�U`���me�����ȱ��@���o&�1���3><C�;7���ýt��p�)�vkY�=�戍�A���s�Ȥ��c=C��`��n
�oSx�M�4��չ7=�T^�~R� ��]n���[��I�ȕ���P�����h�z]�9C�pB�bQ�ody�~��h��){�Z8c�7�t�#q�J�d޻��O$�]ǅm�	S�PV�B��J�g.���m���]0�]'r�0�ۗl�,3�8�Z��x��D��Ū[�&�lQ3�eJ'�
V�(L�"5�c�Щ/W��ʖ���z���mg��xa�{Śiɢn�ְ���݄�� $j�/��݆ڵ1��9d�ܒa|��ů-�n���thꯆ�1JF�x��ҋ��
��%�Y����Lܗ�&�-ьL�Z7�is�k��yIl"wv�a��ޘ�q̈́e���m����Q�J����x�9ݱ��C��9HM����N��!���[i�t��!�Ҧ�2M/:;j��ieG�ԝ{��x�ͭ<�ye�x����uK�uݙ��ɚ@�6D5l�����.��qt5�Ө<}SV�/-1�ټV�j��=I�Z�n%A#����5�h����`i��:sW�e\��	X����=q|�
&��2#����K�4ȵ�A��+J�lُq�\����vt�t��iV+x��\]P�JG�f������\FX�_r��t�9Z1%���6M6���Z[ٌ���f�VX�1i�7۽��e�7~�S����聣7�^q菙�lpgIS���/�f'�8�3f]��H-��"9�NW� �k�oo>�㻹�-�K���������=�_ynwV77��2V�qTY`�u=s��y���� ҈Ԇ"H��hE��ծl�� O/ϰuj��.!/
�DL�)�[�(��V�k�����^������^��:SRc)
�rp;��&��܉���� ��75��#�[�K��iW�x�'`�ɂ�N
Wǵ.gR�t�T�scPÈp=��WR�D�J�O>l|��5&���K�<� ��PA�w�~�Z@<X���eX&�s��wf�g2z�8t{��&$��n��}d�d�q��Q7�n��[�Y�f�_�ٜ�i�\�MR�j���
� �Q����
�m��ly�f�+�wL�~|Q�E������-�������'��8��R�c�/�:��A����Pn
�X����b�1�D�+ҽ������GMRwD��X�<_lw p%26� ��V�t��2�xjۅ�x0���6�%z*�;���1U��A���^�-�l���T�f_���mΜ>����p&\2��(ɰ"<��P�x�%��z�DW#1�&�a��;��9Nݘ_fƨ��8����k͏/8��\U7��ݓ�tꑈF���\�QK��Zk�u�W{-��T�!<�@�P�Y�,�AHY	 XAE!,�E	"�AHH�$!$�d  E�I!,���,$I�Y!"���P��  �$P!� ,P$ �`H�P�AdP�d��@ R�	!d (��)
I$��IH� � E�H)$P$�d �	a$B�����XX$��E��tu�QWt]\Uu��]Qu�U�GQUqU�B
��� ,( �"�d "�E$ ����$�X � �
�) 
�d�(H,!!"��HB(�����!!I�o��M{�y�3+�ꏾ���SFZ�b�N���.K��,F.��S�Xh:�������K�q,���;���ǐ��0�~��|1��i9�@֥q̿U�dݺMj䈊6!�c36p�	���������*����g���ăz��x�xM��nz����=�*���=Oj�h�CTķ�h==)R!�jIuSı�<�Sт�:��p����]�������'B��#�ȣV&�E���2����z��8��ݧ 㑄2���o��Z ��	�ggc�ϯ\�>����[�ɗ8p�/��,ϓo��������a7�=֖S�G�����[Wd�����>�ȘpN�|T���T��I��yr��򾛰�ZY�BC�xD���x����^m��NEn�ʻ1U8��mi��Y.�Y��G�`�r��qfA#W�lf��/1x�M�t]��nu�'�D%C|4�H��f3���^�A��Q��m��� ���=����s�6rƽ����1u[���{�ޓ�]��dJ��LL,�yTFZsu�Uo'�O]���f^�pQ����$g_t�ũ�9�x�pUs��F�sr����1w|>�v�<�����5����ü�lJs�"��m���}O��\Λ]�{r/E;z��{��h���	��S~žׅ�5){H�z���ج��:j��7�<����c�*��gM3G���3�z\��R	�z�+��f�M�K턇禄ޫ��u3�P�ʵ@]�}2��ҥj��Pq�}�\�Y�{ ,�m��W|��X�..l-��{�:���|߀�k~>�o��'�������^��x��2�a��Ɲ�����E�W���z��CWn��y0�<>7ƅ�d�������#�����uܣ����?�
^5�2��r���w
Ī��jU��t$~�tM�=�5
@{� m�^:L�-p�i2)���xT��3�kmJ�g�g۾=�i�uj�辛�rk�wX{���l�K[��] l�����޻�q��K�3��>\P��B-����LЄ޿vqh����f��(�x�l��!�#�'�q�U�EV\J���wC�����9s�/A�F��9�hF����RwO�R�%eAG�ػ'�v����M�-����j�+��6�`��C�ܣr��V�lŐ�ڹl;ݯٷ�[Եl��L^�	>j_k��"/]_���(�bnlD[2�����+ 0��õ�9�PU������p��̪q��,�|��<Ae��L~�֫1��Pr�7�=��
����)�C됾�{��zm�ǈB�N(�)⇻�Ji N8�{}�Q�b%蠿y�-�[���42H�c�F�֗�>�h���ą��1��s.�p�:���f��K�5|^�Ŗ]L��p\^�sc��XtaЍ-5u��\��'ۛ�<c�2� ø�����_}/�B�{	tWy��8�_I/S���a�JqF][��fPwk��� ���;���vOx��>��=��!��|<�GP�y��1>�;0�ȹ�o��F��4��ȥ�g¾"}���)�v���כ���������2����R�~���0�U��w�Ӧ�0���N�`l'k��5�:k���|������ʛ�n�']\�EFLQ9Y��C)X��a�3��C��D�yyS�:�Gu�5���/vch��᳗0!�\����쳹\�<1���ڪ˩b�p�t�O̹�D���9l�Wh�7]�S��զj�����ԍognӗ��eP�i�ЯN)�QbM
�M�z��T�wH��o��.�IW����v1%0������=�y���n� �'V���>��̍�T�n��dP�y�64�.�H�<�.L@�x;�K�������5Ph���a����o�L�MDb�Ȯ�rg{#��_I煳��ǯ����=�R`���gN�{G<T��7ة���,ii��v�K����m{=���}�z��5�q���XY��"��2��=%�/wx�$��^����|o�v�T�oO�/��o�Zvc�R� ��9ޱ��9�nG�L�m3K؅��j����w�?jO:�ы�~�qa�+0H6
�#ee�co���{�Z�a|����x�J�Ŧ�䏂]�;�}��Qxa<Ƶ=��d^��̶l�B������=�<�6�X�5��B�eҬ��p�h����BL#.R�����o�1�8��I��v/���ްx���r�����v��y�s��X�V]E��Ϳ�T�ϏK���'�N)��0��z�>���_2�������
��ͨyYa�[�'�\8'��ww7��zb�������c�Q�`9��zoo!si�&�-���<l�p�Gc[�~������cM��W�ƭ��j[.Oǂs)۫|�:}���p{}b���W��;z{t���/�Tf�*��Z�[+r�tq*���a�n�sT�~-�^g�]�Gn����ཞR�lk���`|�*N�8l�t��Į�{���z���[�gW���w��Fr]\��!���bu�=>گ�'�-�Z�^o�	`t~��#$�i���_��3�!R�GM� ��PIwɣ��"�Pȼ�k�d����Xŕ�U��f��}.���u�!
�T��. <�ҫ3�Ю��d��%�\�V�I�77>��W���C,�n����ҝ�#$|�����������ū�љ�G!/�\1��o����nD�����h��ȸ���Q�R1b���W����'v�ʝ�8�Ç�{�Y���=��&K��5����	x�˾]/A�/�zm�\%�����3�
��8���٧
��M�����*�]/Z��.�x]+��w�����=�l�?mڲ����bg6w�����5SmV[jml8�X�D�ȬŖW�!�T�^z}#�Ɇ��C�Gh�ԛ5�# ��m��x��6z)��r�Z=�/�[�Mɽ���=!ܘ��%��}�۝{ա�},`{��S]����;8�z/��/{����x��Ɗ`�ze����=������N[M���z<-��4�+.!,����s=M{A~��A�$\��6����xl��,�Y2�{M�7��c��7�=i������yy�s�M�'�ޅ^�Nt�:�ΞF	7y5�o���.��7oi�!k�)��i��©�7�o��Vd����2fFwH�R���Mf�M�w�L�2.����е���������ڶ�8�9�l}��Ӟ&��x�o�V,�ѓC�ݖ�7�Q�ozWU�+�Ũ�Ξ���h>�9�c�{_�w��+u^@ˎ���qSЭj�.�R0/�s���(R�T���r�T�5�<W��2�}�{�[#x0�7���n�>����f�?+87�����2�!�x�����5��4�yg'��/�&w���uf/?P7v�ŉn�E��&�r�˛�K[G��:�Ŝ�ʔ�g��A��e�djO��M���%�~&w���l���K/z��ǝZ;�ҧ�x.�mNlxqx�{����Z�[�T����T��BÌ��	�wHm9�̱̅F�V8��3�;���8�i1�X��%Ӓ5/�{{�pj�Y}�����.���Og���h=��;Q�د�&��Yp�Q����&v$��y�݃x��:%m�ķeY7{]��X�%�@�j�:A?��`�U���LN�w[�_�!h�Gl>��[�4���Wg��h-%��<�{�B��a����Z�)�[�)�����D�՜M�Ld��������"�0ny�s\W�Hy1ۃ����jh��k�s�}'�سt傞��HW������Y�z�Lkswq{��rw!Sw��:����]��u��Gpv�+_����G���ZgZf���ӭ>�3vv{�"퐟XAK9(�����Z~�7�Q�n��9���GP^��y��߆UO��;��d�"l��A�&]�\�M�uf�:�L�l�#�-.}5=�nL,�'��
xq�����o㳇�1� �{dg}�?N��=��w�%�y�]��l�ۀ+7#(�X�ս˛�+{9��p����i��=����y8��oY��~gȁ���3��|�G��L"T���WzO�vĺy#���K4�v[d���%����&-�� gn���ьo�\��־�h��w|gC��b�B�z�}u���R�g��M��h�za����_�I�ܩ>^� :�m�bg�xo��jn�ޣ�/*VOt7��ww����N��9�}U'�ї���\����7�w5�����װz�Ȝv�Q�=�V��5����VƇ��OR�p5���$�/���λK�]V�a�\n똥8E�Dh��8t,97:����<��V���ߙ� wE�os����Gr6���׼��L�>���gۦ8�cqڗ=C�+pj���/_
i�QrI|U؟�_n�:.���u��=��HX�Ɇ���wAa[	�0Ӛ�0�i�Լ��]�d��3�/����W�'vYy�p����~6�[#�e^"J�UȰ�{}�c�`5�۲rkܟ�����e�V.�'w<�ɞ{ikz���f����tW87�	� �8���;������ �yxXI�3~�չ{X���<�q�]Lp?u$�E���"S�*����ާ���ucn��z�v�)=o�,�����ni	1�&,�t�(������f֟����ތ���X�=�QOo�wt��[��4xm:;��9�������E7>wc}2���W��^�׭���Ν�f�|���Og�n\��_�j=�u^j�6 >C�Ӡ��swYJ�+�W����Q=��8գ6� ��XV���o�s��������ƞ����IJ�U�#-x���@��A�בD��V[v'�eO`�-�6���5��ݚ�eW�h+�k�]N���{�x����i�+Q�e^�H����0��X{{���|,2�p��_��`�]v��ۋ��MCJ�y�t�b&���微�ZV�}W��^�}$L;k�W��.�|{���I`	ɳ�N��mt+w\�f�v�5��p��7��g�]]Y�h0)o��ɕ
�ʣp0��q�?<W^�M��$�vOcUCB���~h������M^b�*����v&�y�^�

�yQ��y��ý�J=��}�~|�Dt.ݾ�)�7m����)����V���C�{w^��5j��gƍ��e�O��d;Z�����u��4:�t ��i�=��sG�u��6�u=�:i�BV�\��>�y����%�ϼaS6|��>RD�n\�8#nx����o!^w(����ɗQ�̯��U˼�F3�jj� ��|o ױ��n3�\�/@ֶ�B{NR��&���^���u@{��M����`3��(}����)��,Ӌ���+�����=�$ٞ�-/�OX�����)�si�|��x�)(��9�sN�h�|���E��=�V���K����_�#�@Q��}99���#�@Ҡ�����S�{�}�K�~�7,X�ðz���%��	q`W�	������`��,�~����Fc;6�_����<דM7fA����{��d�n�f�oʥ�wd��1����7�ǻ} ��mof�S���zl%7z�u�h��ml�t��[E�5PW��.Ƶ噇��cwWa\J�'�]-�|�����U�sL�r��,��Ih/h�3��<���3:`ʯ+L@`��x�6.�E��ӥ����/����O$��d�����<�3o���=s�u�I�E��&���v��9�S��>ܳ=��c ���Z�c����gA����#�����+��{�j�/�*{݈y	�`;�aY3�e�GCw�`�c�Qn��X�z9i�z�=�;���>�.����)�h�em�u�狣��{ނ��q�m�7۳Q0X�2:�N-w��S��_i~Oyؾ�/x	��ެc����奒�G��aG�o���v���n�V���v		#,i���2���>��j���v�K%�4qG�7�d�������i��SA�v�}b���Oy�X^�&M�瓃��fVH3k}LKӾ��^���+�o�sD�h�G�����z�E��SCG�c���Ş�����	��H��J�+�u��=�ݰ�������mM�^"���=��BL�Eu=뷈R�X���(Ok��J�=��ᅜ�u����9����{���[SӍ�|����C=}�x�'y)���緵��~Ɋ�b9�V���3N��Q6�s�����C{'�|��f-�X�^5�z�j��,������෎��<O��'�����n{(�>��y�$�n�*%a(i���q�}i|�v
�>�FEf��C�w��eng�|�^S�U�3ۧ�M���������n{ʍ���>��O�~�o��|7m��y +]uݺ�L>S87�Y�Pf�}���t2b��QŞBVn�4�ظ=~$+e��&vUx��ZHI&��[�zf����ȇ��ηN@��{X�����v��u��6y�Φ��ym���� ��4���\�\���{=Fy���r��U{(=����ݗ�^�O\��f=�6���C�<����z����}QܫM��.�=|n=i�樑��o������<˲�*V�|�	����kY�-��b�z�a~	mǂm��T�R����l��6��T$���>��h���g�ԡn�_�v��M�qx)�f���J~<�>�!ɸүa���L8�P��x#&	����n�>�=-d�3#Ӥ*h�����K�([q�=�Ȓ\�����!�����-J�����	R��Tw�N�:z����Ÿ�y]J����������u�I	N ��tj�%�ULէ!k���煾	m���Jv.�x�=^�S>c�Ɏ���+n��[q��!M���9��XFJ�܄��iCFP���-A�8y�m�5[�oh�Kڰ�͎d#-Mb�%Cm�].�:g�p�5�"�;z0н��ܖ,�h���n`Svu�ۄWl�t'Z�]�1�Ģc+|��5�l�V��7dL�,���$	ej�%��6��gd��[��|��m��Tu���J�m��3dWAb��D��S�wG	�Z;uƷ+�7 �c�6צ&<��dMY�!�%�n�S�.�Sp�.u�ҥ�t�݁����`7�5���ł0i�.YP�d��&Zqc��o"x�hQ�VRb���]�6�6�[S�rV紽i[V�ug �e�G������[��Z���S�(&�OA�ch���S[�Prm��ʘ���vڛ�H��{vƷV�!k6&��ˆ/Ya��Ym�w��NS�Pݮ ��n�n&{ܜ�˝L�ZJ33;R$,@A�cV�Ot:� Gm��2� /���ھT�h%ٔԉ����ʣh�Fy�G�8���۽�m���K��b�E&%���Ka��x�h�mHpJX���8�� U��n%'�:����Q���.Ը�1`0�iN,�A���p�n7/��)i6dJ-�sՎ:8�Ĵk9��Z�8��]���:��Axh�<��-���;C�=z�^5u&�
��-�뛀�a.u�[�B��B���\�``{u�u@�9#�M�4��c\2���f3���>�r�A�=Dwh�Qe�&�ά'cr ���#ƞ�yGڭ�����g��kuŔ!�Ղd��lX�G�էe&�-�
�.aRҝY`l���se���(��������yU����)ƷF���e�GZ�[t��:��m�C�3cѹ%D�ǂvb�6ǩ�u��R�����9n2�58ך6�e�	Y�C��]2m���w:�١�jp�.5&�b����\� p�:0���64�L��%l-������݌57!��s�dV�u�/D�NC�[���g���+b��sÞzcBӷl��z�"Pb+�[l١��J��UЛ]� �^�b]�$bOWT�R��CѴ�l����ASZaIn%ί�A�%��ulC�ppa��kc��м�G+����ՠ�v�p/n�{v��X�kR�e}�nT��f��q8���f{W��>���u�u��n|m��@�����h����m�
Q
4/l����o<dS�8�3��z�T��چ��;�WY\.�϶qI��/�����,E��!�6ј�f��m�0vȮ�-8��wϟ�-�ʨ;���I��Ǚ����ݺ8�z�'�`��q1v�t����s��:9�:�[�=㝉�'DTtc ���7K]L�������ِ�-t*��6�Xm�r(�*lJ�a��r�Yhxw������� %�Q�`c��G��t3j2�1��&�Ύ�ޞ:n�C7u�1�A�K�%�JF���\^���f�4��jJ`���&�t��,w2� �[ֽ�7/9yw7fb�43v@�U�d���gd΁��_on \v��]^-8�Ә�F��Nշ��yx�F��\1%��Ӗ�e��+�YvuQIay"�f���j��oG8�a�&��v�yt,���<���γ%٘u�;GE��%���&*�9�r�G'y��������T��qՌ.�J�%� �z=(�G����M�s��y �8��52����M�"Ў�kX6c�mV6b�B�m�3aҡ�$����u�{\�!�f�aé���tu�#�ut���G2�@���0ea�uq��f�R�auw�wa9�-�8�=�Bvw[��z`��O3�Y�+�a�k����Ƌ�M�V."n�����(��C��X��y�v-�+юtg����Oe.
Û��ծ3Ӹ�Q�k31B��1]�"��e�j���[�^�ky��nޓ� ΅�Í�g�qp�t
��Y��k�	�3�;jb��C]p��4DF8h�=�����՗NՕ��i=��-Z�u7�wk���[����6� RPvrE\�"���l�����4D�gxƺ���b�ۋ1pt�5cq�ܢL�s�`����Se�uBk3/-ꑸƆ"�<�R��2�vqE8,R(�"M�&�	��Fb�4�%DeY�����ȶ����3I�֗;�y���m=��<�͸J�C�lMsi��9�<2G��%�>6�ð;���"DmD9L���g�_�YIP�?�Sv�h���c���G��筦�kf�mu����G�Z��n�uǳomgQ�	I����ÝeM�--�B9C]fIa�j��	*i�Ō�$T�R�����WXh����b�3B�RYH+r����oVj]n#!�X�(��u�i��ՇmAaF�ũ-ƅF]J�vbX`�2ù��u��crv_��v�@b1���#,�b��4�IMY��]��;��x��3��=��g.��A�5�ۧ�<,lE��p�;1���`������������mۤ[��R��=fY؉Π�wPF�7:e�<��ݭ�����\Mp��\'䧭`q�W�,v��ZSn���Mt$F>]m�̵����ҡ�n�b��bj�0v֌X�Dt!�s�V�o�l-	[�봗1c��;]4��6-	U�m���G����3t;��+7k%�8�\v����k���U����۵ij
9�KHX:i[1�s���'�:���=�wSkT���4#.ڞy�HK[<m(zi�r�9Ӟ@	��ؼס�psm�kWk�N�]!!M�у���s2WM�cq1w[Zn�̹�J�n�v.�7��H�<qޯ玅�/�����<M.��4m��H��!���5�Fd�c0�Ek�%���ku��]��5�A�r�ˉ�;�Q�w'����۸��GŲ�0���f�`f�ذ�ur��T�c��:L�l�@�	I�Q���Aғ�5x�ѭD/ZwZ���N��KK�ua{�i�n�,��cX��{[�^�Hh�Hr�3q��x�l���:=�&E�m�.���e��[��I�q�����i.xʴa���̬�h��8�6o3��2�	���/,�b��q�.0�����P6j��H�@��g��� E0�CB@��X ����q6�=����^eAZ�3=Y�n�'Wc�7�v]R��,*��n�6�au�j��Ƶ�����H�M��Hc��ػz�v���n,�yXHL��ݝc4�����#-�a��˸�:�n6��q,n��zŮ���mF�s�*�r%lm�*����.�붉]q�1�d�b]ܵ�l��ձ���V��8u�B�����*LaKjA��F=���庙�2�Ѣ���@�95�/nn�nHҠ��%mB�F݋-��e�Z{�vyy��y��$�
Cn9�'e�-{8|;���wnq����.(�m.܍�!Mɥ�-�Kb�4x�ڥi8�Z.x�mϜ�ظJ�M c���Y��٣�)�ȃ4֥@���깭%.`/$�]u�A�ҋ �<�,u:������6�Ri�w���#y��I�j�ͮ9`lQ%�.�<�B�;u��KqHJ�u��4&�Y���×bRh�-l�؛;�Μ������6Mmt��*ˊ�,�ܱ�=x��xaصtڕ�$Fb����8�];֕�)�ui�,e�4�K6�XMwb,��Fd�v3<��+y.����ON��&KVJ�4��.
h�
��@]S[ļP��Wm;:Ǔctq�m�v2���Zȓ�ni�M�CPcn칲�5��k�F ���,(��1�q�[,%5ԽA���wD�9�f^&�:���b1�/[^�d�@�:DS��q쫺:��-q7��ݶ������n:z�6ח�lE�(.��bJ������WP��UzT�v��`�u��}���z��E��d�����p��t �X���mΪWx�v�X���6��4%t��I���K�6,�9�R��Jn� 9�:��"
��ღu�ٔ�1�p��r�#���:�P�
hs�3֑3Z3�Vn��<x��v��hL#(C!<1x����63r�V:��ϟ1�� �|�`���'k��t�g��v�{ptf������t����g���4�n.)�@�X�])	��3�W\r쐚=��Y�>r�4"\���嶒
����f]*��Y)��k՞Z7�]+��+�$#v��ݹ,=:ف7N�)�����<Tֆ�Gl�i �${d���ތ�;5X�4�d�,,M���h5�6��s�s��1u����tu�s�W	%��a�jЁ�2�n(�B������io+"P�v�͋�X���0n'�d���m�&y.�sQ�D�lih�*ɕ���l��\;@�x5�ƥx���p�ʈ�3cLM�V��nۘ�׈�A���oX�#Waˣ��"n��nL܃rn%Ѹ%޸s�z2j8���r�y�$�xK..ѦB��� ���ֻqC����X]��Y|�\�0��rq�-+O�Ůq���^�v��n8�X���5{[:�AԆ�W�a���<������3:bӌ(���H�Z �e��LȤ�c���m�����z�\��4�Hc����O]��J�H�k�F1I��K`U��:�ۆ���:mzzYB�1]�/K����BSJ�)cX`/[BB�6� ��hGk�%��s[���4�[�<1����v�j2#��e��.��oMF8bӈ�'B��Z�n�n�e�q�ݝ-��N��q��{A��m^��#m<t�s�v�ݶ.J	h�^�]gq>�>)x��&�vݱ�H=�{:ڮ;/��p��t��8�U����kSלa��:݃�5�6�8N��w��T��O5�@\�Et�Q�e��"k[��jA���Z�������9��@p\QY�vujT��;	]�#�'��s���Dt�!8�.�AN#��!ә��IӤ��䃂��6ɚ��AH����.;�-�)$A�F��8�9.�,��q���ʛ]��@Q��'G@\����%9�I�6��3N�I�E����$8�'GL�ggqte�S1pQr��IAӜ�A(�vXt�6��f���'JT��E�j�J��:̂&� �`�1TG� /ಾh��� ;G6gE��Yt�܈��K(�nh4Vj�-�m&�Ҏ#N�͸�,�[m�Bf��o\@�z	�6��s�'Zt��o1h�����N��-���,2���(�.�3cE0�b�AR�W��e�����\qGz�v5j4jz����!�ʅ��c��84�EmϺ�浺s�Q�me�B�΋�7%��:�e�q.�4��R���B�WYܑdï[�kr�n�v蹡9u۠�Z���i��q�VmKt�7dvK`!��	(�r���R���\�8M�l+�tdMv=o��%�kR�SQP���./��ǔ�@c��`%�����b�-	_,���,tu��Y�	�m��dGF,	� 1j�I��yk���JGn���! J3L�M���e���p�COZzW�6�,�ɪ�Z�*m2v��.J��´�t�ƬR�5h��G(Ĥ;	֡7L{:�#v���T�}���\��]��Ă�듙���g"z���x'm��	=��q�6u��_7D�Wu����B9ܸ�£�#u'�N;�e���"�و����wj�:1�ь��n�TKqsH�c�)����Уn�c���σk�tMq�N�vu�^���pa0�Ţ��`ƀ!q�&�%��5�..���77/��r�\�`��N���q�:�Ng��%�Xx8�1{!�|j��m����麰q�n�����ʞ:C��/�S�`����8��썍pj�B8�#Nu�-�-���J7i��E�]��0%�Gv|O-�6뭮��Q�`5�5��3�]q�muJ�X�fs`��g�e�x�t�r!���=N6wJ��>8:�Mx#x�'��B�ss����Ls�^�x�@XnD����#ۃ�t��ˁ ���ɱ��)v�77m��*�^��`�v�r�&ں���W� �K�&3�3�t�:K�X����T���۩2�B�0�Md�H��Ų���A��[[���Ao-��x���YJYV�VŖX��ZPi�Y��� s(��H�JQbVXѡB-k�J�P�m%iN��-,���յ�ʭ�/^�(UK mAZR���V[m�KE��VYUA�Z����ג� ��N(�I[,m�i?���S�C��0@��O������hz۟6K�g^-h
tWݴ�R�*����(z �̯����y������;ui���u���~:�A���ux	ݤF�@P ��DOJ�S�����?d�����7���X�~;�><Q�h/��EWH���׏��ݕ�'��t�� 'v�[ܧy_J=�M9���<o�s( C�ӧ�7P�4�y����]�<Y`��r����<�=A���RNPu��h�o=��7�,y�h�v�̩�A��2��-�SJ���~���;�1��4_����U�=�.&e�G2�5����w��|~[����-LW���M���p�<nv�b
���b�9ŉJF�7-����w������-�����uS�Qai�>��L�&�������y_�e�&eئeY���PM�њ���M��=(hdu	����*�<5-B�X:|#�1|pf�w��ڗ3��6 ��Q�ٯ<�B��#܂���
�;zP��Z
Ci��A7�DrW۵'v�6h�^�:��S�2әic[��6�����/����S�on��� ~#�H��4�_wk����x��N��!�S�	ޠ�t��Hl��v2gz���r}��	̠+y���3(��/�1��R��9��#v��H�����V'��{��� �ւ��r�W_q�A�D�y�jf�S�b��U|�U�,�ER���.���.�;M�����@ڎ�m��߿�?d�� F�|��A|wNf��O��h��C����u���A�X �m���ݠ�� Av�F����Ƚ�!�W��{]2���S�4ۓ�@�e�D#v�n�ϣ�����h�A;� H�H�7PDn����п	�\kN/vm�썁}������z�΃���ҡK �;�ף�U��]'Fbvf\�?c3�k�4n��L��R����.{ז_z����#���^��U��2�3u.����UAG��"JD��t�����׍�m����/;WO$�������\]��s*X�U���[�U��fP�s+�Q�&���K]O�ܟ]��@)Dn�#v�ܙ�D���}���C��X�b���JF�vlh�6j��Fj@��-55z�h�)�x{��>��,����v���$>B�h)�+�#E��}�־~�u����*�1̫�̻��@gJ�̂n������9�x^�R{���D9��#um��޾��3����A)|A-� �i�� ��NfP��|�gyz^Bk�yB��w��'�{��N��q�XfYbfQU=�o%�񳠂5����t�{��>B�h)�+��H��������a��f(�o��<�˳�?)x����_;)�#���=��Eg�Owr��1.U�o{={��GV>*"�7����������Y��3�ב��V	�YB9��n�@�ӆ�Ε͠�� \9��^�]=Y���C��A�n������Oo�K�����꾓�mS\�s�y݀�WYD�1`��4����[h2d�&�ԛ5)��YA�C0��@n֍������Ц�b���2��y�VAr�F��)2ˉ�e��6��u�[O��5�&�_2�@{s��� �ւ��r�HoY�^��߷�58�*uϊ���3,/��(F�ۈ��;��B¦s+XW~�ռ9�}�s�m�w�X��q�X����}O53��^ՙP,��u����k$�UPs�یY�8��uO
�/fY���h�\L�-���Xf_&k�[����������y;���6�?�`���xf���`�������{�����ǟ�J�y�7���w�ѧ�X*�٪���:��R��v�1_>�������w�������|h=�[q��ZC\c�1ٹ�[�y.Mk��D�ۧ��.8�.Mn���g��c�����U�s^^��:�fŶ��78��i=lbg�z�� K�n�5�U�ݪ'�q��:k�+��YZB�	j�X��t�U]2�cUӋ�M&��k�nI�V[����q4�M�>����]Gf�62϶��u�ĭN��ك���T��)���_~_���,.�!�Hͮ�q[o&��K�Ϋ�.4q[�^SMF4Dv���[��,��:Q�9���V��]f��'/��e��stܲ��A� ����!�� Av�w�N\g����	�>u�c����یY�	̠�. ��3�q���r�bŔ#u�_{kO�ቨhZ��ۃ�@洌����Z�Dw]fe|32�1ˣ+��:���m�A�����1�&mp���hz2p@�(���z�z�g����4Zw��~��Q�����%*H�H_wV��U�)��}@�s(s�1��s,�I���ݴ��j�WEi�Gs_�p�
���FE΂�ۈn}b����x���#gu~�c��o�&eˉ��s��~�O��nԩWnWݝ�F���JS ���"�����Di�@�wh"=��]�$W���3�3���e���g�ر��C����ʯy#t�p�=�C�b�z�[�u�����5�Tk&	y(��9C��J ��}�[b�x)
�FN@���ݺ�V�۶�B�G�H���_-4}icL�mV�uz�~�m?����,�
�2�r���(wPDnЯz�{޸�\������b�Ծ#kH����>1��1]�]�z�!mn��W��_����G����]L�-̲çLcELU��Ӯ*�.�f�a���~v�!��pL�.c��h勾���13�����E��i�N�K�8U��g���0ljc5�0���:��ce���2��rwiϱ�1��o���o�k��Z��ƽGɟQq���̰���q���צd�5�^���P�7&�(wnz̻�+� ��  eBݭA{������㊁:v���?-�/�=�����e�ԯ4Q�Rڠ3'zx{@�W}���"��M�=_n���oy	w<� W�D���QѾ�Ctb-;�s[jهr6$h���:���������bfT�+�R��3��^uf��|�֐��|�ݥ���I�����^����A̠�"��%دy���l�����	ӥ7h"7}��_��J��]Y�1�p���1]�\��@��T!N�Ӕ��A����堯�H?v��f7e�Ÿ,�ۧ��c>���޵A�QэUi�y(G~��y���3,�0�3�A��CY���C_ƒ�Z<a���Df��kHGv�?n�>X~�s�����)	#�/��m���hG��s(+�:kXuּA��xB�� p;��/�֑��2��e�Ov�	Ơ�L�������C*�� A ���t����s���f�}ꠀ"�A a�|;���1���d8�=(p>:W�{�k�=�?�W}�_YA�2���J���"�= zg6���_r�o���{�f���ix�����j����߫��������32�E̩s+�_{��]�WK�,��ܰ;����f�|G	n`�����QF����T�Bcx.3~L����bAuYANY���j;]������3l�T�[9\�q��y�,L˸̬L߷$\`�L�K��q	�D+N딈.���O�2�&8�9�ZsW�Ǯ���4���!��)���5S/D���|t��D����%IMQ+�%a�3�?<�����I����׾ӭ�u`y�������}�A~q�("�ZfYrޕ���F��Ӧћ��oW�mi�<K�H���_q�R#���%L����|���;��;���7P@���Yyʝ�V���k^���.q5114zr(��"7R��i�p���g�#��O�O9�Q��LU�*�=�*��1��W{j�������iM����n{�N�Zv8V�g�S��AC�ևBY��Z��k�>q�1����ݴelv��-q	a����}�c �ͭ!)4�72�j[�-�Wi�հ,�%X�&b�"r��f�-5��qlu�i13�^(�{6��&ٮ�հ�nN:?~]m����U���:rsx�b# �ܹ޷�rv�cZwX�TW���r��͝ц��8`�K�e�5������W���wD�M�j�h�⹨���5��цe�ka�]c�S��]=��h�츍Ͳ��n�U��'�_!�_�@��'�q��n�>h?=������ٷ���.=|�FfXf}slM}�ѽ�:�E��_ZB�s�q��E���%p �yH�6��]�����k�@|�<Z�~-�}��:t�7hyR
����U�]�T���&&�N|t������+�2�Ov���
��V'�3�_B�v����,gvq�A��Џ���#T��qj���3�Dn���Ҿ �7jA�����L�}CՄ/I��]���E�u뒸A����Bv���O�d{�y�3��+B�sRӨ��uf��.�d9!&Z��h��Y1>�^���sW������h��,q��9�Y���]w�y�LLM���/A�oNE<	��� �ss~�ћ���ӿ�{ڔ�[esy�vy>yg)ę�������˴&5͎Z��(�Gs�Е��_<
]�G+��<�{P��dH;;Y���H����dq�Ƕ���Śs_4=��Wٔ8�����T�N+]��kv\���L�,L˸�bm��\��IL�u�����W��\��m������� ��Eg;���( �����#Ǌ�PCi�u�/�Q���zr��DWW��������:Bv�@���� wkҟ�_�E�B�]!���/3�8����Џ����PD9A:P �ٓj.�������[��t]>���<�{��v�8彺���Ԇ�F���������~��̹sK37���w<:���3~�+��Ľ�u��^� �]K�X��V&9r��-.���{�u<t��A���fQ�;�
�LF=9|t����Ԕ^^��S/yw雭3ܠ�jd�ķ2�Ds*���/���L#�.�څ�^�=,b2T��U�Sp��O/�LS�&"���g7�y��47�/���ʂ="�S�W|,/��b~����u8�;�vy�>K������ħ�I�'�83�=jt�k���ʞ�Dљc3�
�.?���.�*;%ܑb���);̏,w��<�i7�����y�Њ���r��&TY��<�]�F��ߴz�N��^��Os]g=}��r��w��}��j{�N�}���c􇏴�ə��F�<=�c��`Eti��YGQ��Z\Ѩ�s�qsó�����'��]d��=7L�ď73ufQ���q�aS��2ث<[VR$�Q�<�{���O���ɤv��琞�
�@��f���bXHt�'���gs%�Ck����*�e���r�}�Ss=q��ӯ �������)��u'p-�Ak\��^5(ś��^^��8`�g�/eS�/3�Gp����9^�7+5�j�~���_���6�=�k��~.�Jz�^z�W�ˮ�h�h�pܭ|7�"���O`��	ry���@�[����*��c���ws��2f�|̞�_��3wV�e�������\�������֋���w; ,�h5�X��8s.�=C��G��*�}��2�jĿ{���\9�@,���c�w���H�ŋ&$��i<w���2�>��S�aQXs��n+��yvw=;�܎Xx��۞�(Q�i.扥?���g��ݦE����j`��Uyfi���_�� �!~5Ed#l�����n�mև'gm�8�6��Sk*�tu����;�..[e�q"tWf�
t��Nq�;!�֎:8;-��Ш��㜊�."B��E9��v�E��QG�Ey�HtD�x��*�Z(��*�n���9��ܨ�;���]�wp����^k�8�r��gRWmo5�����u��Q�[kL��YE<�a�vY�YE1k�:,��x�:��bwY�\�n����q��9�6����_��p�A�١us(A|t�@F��7Rޓ%v��~��`����A}�HCw6OL����f�rW�oԁ��zVc��� �F�B�;��:t�zh���G���oxp���T�b1�� A����8� �Ծ#kO��z���ӣ�tn�ʻ��U��ƛ���t�����V,�F�t�f4�0���O�i A�v���v���o9��8�L�٢�qQ+٥5���3�#%A�� Aݠ�\�=�3A�\F�|�����rd�9:4��\��M�����o^�s��KP`�"<���ݠ�;�/��A�u�hR���7��*
�PF=9���D@�����˖�U�T_ٞ��<�VDC}�c�ՈAݥ���s<϶q�L�٢�s("���:cU�^en:�m�����k��PR_,���cZ��,�+�3X=#�O��jz�����m�'��[��@�V~�Qb<�e��v.e�u� �}���V~��}�|��kg��q�Zm7P�����s)N�w�#_���-��$�ہh��7R��6#�)� �.W��4�.ם�V�i������Yd��3� �ݠ�#u���_H;��u��J�wjz��@p��}�_ wi�v�9��wo�%b�J��i�_"�!���{j���&^��y]��P_����o���~|��C��"�������#�{��1Ƴ���6���\A��h�n[�V�2�eK٭�N��~[B�f���� ����\�w��Q�#9}��ݙ���[}�e�/����ӣ�O�n��N����Q�ߺu{j����ov1~� ��~q��-ߐ�++5��!��h�m�/��Sk�x����Ê��{�%5�.M^g�q��`��=BI��e��8,������|�:QB�>Ͼn3�ь�(KI���6�\,�3̺݉x��������ѳ�41�Ҵ��b�f�K���PRk�iv��,�a%4�G7U`���v���p<\sl�^�����p+�˔���.�`��6�n08!0RZV��*K֒��b��#pF4�8���nwW�8�i�<��N\����3Xuz��:c�0�!�5ڌ������pZ�]a!�-�A��`M�&��b���Y�Y��BZ'���� A�Dn��ݯ���������~�+���x�"����������ˏ;R�2�3*[�E�y�ӳ��yѷw��}�#����R���[c' ~>��6 �#u��v[��/�7)�����ݤA��կ�+��Gޛ�7^��;�J�I�h7���@>�8�N�#u���3Ջ��|�D��˂f]��ĳxo}�w�m��m�/nJ�����^�r�����:��}K�c�̣�e�q�ѭ}�aG5e���$��b�sB��N�A�b���SF]y�g� ���f��ׄ�����i��v���0�˱`k�+C1��[�؎գ]L���D<B����[2c�6��:��,��x�m,��Ψ/IB{@��7P@�A�O�k��Kc��tÿ�)�߲uo�{��ӌg
~��6vz;^�zi��?\�$���NzU����bg�������O'�s��
 �����?:�P��9��c����E��_w�ޤAP��r�����wX(��Lwt/{E���[�73,sܮ�5M�qH檭��[,�1�� ��Q����\fV%��b^����:�+ܯ�^!|�@��ݥ�fȞ���N�x�}9� ��,9�7��o�p�&e�&e��y�\L�޹^l�};Z"z˝�~��W�{�+���R#L!i�E������=��ķ��(�hM���rVW��=RcEV��0�\�9��hk�貘�O�� �A:Qn���zO.�׽`���&Z��fw�<�����ϋ�V%�̫c�V%'u[����̙�Y̥���og�C��[�闎1g;��(�#�L������P�� Gy|�8x��A���mim'Mv���3�G��j[�fNS�;��1��n.͋:�~�;�7/��o�[��h������^����&_�����oP��K:�}��}�ޯ����9e{������z�j�;����#N��|c��\}=�MA�A�u�OI��z��1��?�0�~�]K���"D��O۵�N��(��Zg�_ܥ�+���/xv�Y8�e��,�}@�}� �_:P�����������SFq�搖�C�:d��y�q�^�yy=�;0x�cTs]�v:�:��~����o��\fV%�z�y����v��Y�I]�]�X4�<o͚����� ��H�P��h]Dկ_\Y����N�3�OӨ{�t���>�{=�� ��|p��A���c�B�{ԟd_S������b9X�9�h����.��Og�C�R�����,�}�!��҈#u���}���W7�^{
?!�A���mi/Ecr]�����I\�����>l8�6�A.[}����uc��G+`� ű��y^���(���/t�3�W�fZ3Rܣ������ I�����>�X���ݠ۫�:g�)��*Mf�-	�kkgx�:�)�tA s���J �� �A|3)�{��NZ�Z�:�t|H{A�kt͆%\���ŌZ�-�d{Ra���ln��ӽ�#eZ;�%�eKs*��|�v�-zqt�����s�P��@g݈ y�q�-3(�lO�{��O9���T�����]���RϟY�+�����L���81?fw�ӿ`�=�p`��A��:|F��ۭ�����~�Q{nT`���>,�� �#u/�ZBv��}y��l����H��@) ~ݭS��v���f�d�P'�A9
�C��{ٝ᛽�[���#����@�:~[�"7T�ڂ@��vh4F�=[���RϷ����������!|wiN�_&�Փ=XQ-�����*'gUMp�+�^Gvm'/������Gףj�����`�;���u��aM�jM�u��`Rx�W�T|&��� $�k�*�X�U�kF�X�e��X�l6�K�mtu�]�F�O��tq���g*sS�w8�ͥ].n�G-�f�VX`�� �t#4s5�ڼ*d�jq��rlsFQ㲵�x��׍pDe�N(�M�'a	��5w.C��l�`�k�"� �0䊰i�n��Zid�gw\�`��ێ�Τ�Ɗ퓝[�noEd������=�Ŗ���`�!�b����?_���4ZۥmHnL{V4�a(W�k�M�uH����6�Dx��9���J���t���_���LT����g�X}������>|�rˉ�Yq2�����/M�V�g�Zt�;��?f��ms�Н��e3y�s���9A t��}�<<����VZowb��q�e�̻�V'o�k�v2��C�3��[� ����x�Fw��!�H	ݤF�"b���x��P@���e A�A{��_dW쾸�Ґ9_Yg��1p����#ޯ����:>��`�(����ė�$���(V�j�I�|eC~�9>����:|��m)�����Z+�\�+W���^&�VK��Ѕ��3E�Z�n#��P:�\�N��>O����b3���2ˎV&�u��k�:7��}%p xiX;x��}��V�/���ݤF�B�ݠ�"?,��;S�(j=G���y���z]iMwÓ�]�������,�z�nҸ��/�J"�ڍOW�b+'mQ�Y�/��������u��޳���،��>�^�n~���r�[JA'	����@n�<���}�>��=5ۗv�E�*�3.\s*#�Yz�u޽���,�nwό�o� �ׁ��b';e��X��e��e�����>�7� ��f����P�o�]��J�A��/���u�)��e�yV"9ڴ̩nee9�}��BUW\{��3����Χ�yqF���N�J�9����_;�Z�F�W�����>�� i�Pf��Q��Z�)ڴA��i�;�6*�#���	OǾ��=������";���r[����*��W|~�����5S�*��Y�8�/�#uF�@�����f�Ld�����<�|d_,�{[�(J>̮�}%q㞤F�v���{|v�qa��d�p`�o�e���F�iw�ϳ�>�z+Ԃ�ކ�R�l]}�j�#��n�ϼ5�g|���O�#�ޛ��1ǚ��r�*ںڃ��*U����| ��<���\�Y��v��;�Ō~�����\feˎ�|D�҆��~wW�t�d�K��v�r2U�d+�?{( Fe-y�\��xX��-�	�e��E��XnΓG:�%�ͯ����*!(�p����"9�����c�V#���罪9_%���fCJg\T��i�)0��o\q����PMs���n�hk��2~����Ϟ����7h/��I�Ͻ�v;%bR	8!�=<=�j�Y�6��Ӟ��fXfPfV	�4�:r&o��C�W���у��R�������� Y\�N ��2��J��=^B���I3�sh A� F�|�W���~`�N@�ψ;ۙQsU�����v��7V#��ps*�2����Z��%�31w����6� ���gK��{X�^*�G� O�F�ꪮ��ک�e݋����T�C��{=�K��;(�>�ڋ�M��BX�gz�O�V�!�!�bY�h^~缨䉾K��{_��X�,Ͼ���>̪g�~˹��c�Ws*Y�r�2���a|�:��7�������޳%_�@���s(�Nv˃�E�̣7�ÚwY��a��2^f-�dg&�k\t@�݆W�J�v���r���Z�֪��9�-e���.fT���xZf��s��9\C���znd�u"�~��t`��/��i�y�>9���!p�k� w� � �=�X���=c��*�G�/�( A� F���k�jt뚟Gް����U�fXfT�s*���o�wm���<��{,�W�,���PD������7PB����uۢn@_yD������'�HjJ����W A;����)�q�i�H�����?��A�u}�B�l��}�� ��s����k��T�:����܂��Ծ;����r�:Aa�R�����+��Z�V�
���q�÷J���"+F�o���r<�J��H�cm��g�;|Z���V�?�.x�o���3���!]*�,�P��юq�2�0\���dY��}����;=^�rx�=��V��c������A�ٍ
rσ�����;�G��ŋVx	܀0�Mvn�4G�^ڻx0�UL^A�&^hAl2�$��rU�BXM�������K�mIw �7q��^�.�V�Y�׍j�Z������מ���d�֧1S���2��t�'w+��5����Ăo�y,��n����j�-�O����^˾�_%�#�DZc���7P���;ç%�%�͍9��yj"��`��%���r�}�s��ff5�c��g'�^JQ�)e�yM8.�)�5�W�w�xLՊ�d��7�	 E�6ҙ�z�~k��.��w���.��ӕ�#�"�����L׃�vh�nO{|gM�D�i�ss5��8W��BCK����7�;ω���G�~>���Q�oG�ي������Y�}	�_T�M�ź�8�l�e��!�Eu�/W�ߘؠ�5s��9^�[�b�Õ~=��X-��)y�>;���օ�7�m���/���n,{�gWżǱ�׋ �Q�WA������Z��ٻ�i��v��xzaj��X��vm�J6%��ǽ�x|�'����o����H�k^V��.Q�ˎ����,�&{���NFdJ�>._D��[���}=�hD�Ii�Y^3��"������� D�N�)�8�8r��9Π:������#����);���).:.:�+;�#�8���;��: ��9"�:��;�:��hͫ:;���GGvgQB��:�� �'mgI�Rm�.;���6ʜ�D�*(��QA��ge�'rq$IRQgY�E�U��E��;���(��͵܁tu'u�Y�Dԝ��At\sا�]�&Q��l�fkI�W9 ��C-��\���\ń����xy��-��Y9�}]qF�[�)�ڳGk�×ΰg��J8e;x�%�����u��%K�ɀ��u��n�q6ۦ�G4]]l�`R����}<�#�mX`�3C�
镫��LT�Zc��,#,&n�be�ƍ*�b�v�XXU��<]�RE�ۧC�64�����%���@4���p0�jl�\@�]-��p�u���<�y�ͫS�RԂ(�c]����f�*Э�`h!j�ŷI�@۳��`��XY�亖ꦢ��&Ż!	c��k4�����̱h<6A���cvQ�Sc&e��rc��۱j�R��إ8띈 Cَ�ۅ�[��1��x�x7����z+�8�i�����d�WP'nh�Y�(硴v�+�bx����닅7Y��V�ۤ����]��%�ĊK���).�2V�e�:�h�u�+˸Ĝ��5�]c�N�	i�
;e���a�A����]�MM,��J3+`!�&�4 .����1MB��s�����n�\n�+i���.���[79K y�3!'���M6Ԫp`�;v�5͞v��%T-�.<�6n�3�%����rix6�\�D��Br��n98����q�[i�X8�h�^�v��2Q2�LM@�+�ŦK�u�\��2���pU��mT#/Q&��۞���I��ą���u�mʖ,y��X|�� ;p���NvF��8x3��.�\kb�����s��l�Z�ۣ�&�[-T@�t��tlE�-Ʃ�M�-6�j�'�ばhKmn��q��Z�<�ί/	t
������n�I�,7��Ř��Ḱ��0\
n6�X�������!�3) ������e�Mx��r�cv��ɨ7�|��۴�:څ�6s�Jw��yg���F�Sɭ�Ԏ%�<���3����V�\���^�FMun��k��>�na���vu��憔r+�5CeM���I�'wo<ρma��픥�v��`�;p�/<9η Kc�2�d��]�&�p�ja���Y�s".!�!���;q��=b�ٌ�۷6�J�[����S�IWa����M(kֆ-�h9l
� XJ@ك���%�ݮ���sֶ ���`��4$f�2�S5��A�I�r�]��e;g��eϬ���Ӝ�+{4%笼�ks�LL|�?�����M�"��(Kf��)�f[�	���W[#v:�m�X7I��&W�q��ݤ~ݥ�y�������W��Y\Ƕ�s{�۾�> ������Yi�v.e'/��}���^�x��#�|��=]$U"�����W�)�b�ڽ�n���op$��� G�|�/��;���0ء�M}�;]�v3�ZU ��J��n���ۂ��@�b�����$?n�����o�f�ge_��m}�� CН�S���l��tX�ya����E����7j^�V:��3�-��o��c�TEy��� ��@���^?n�K����>�����o���s΍�i�LS�9�t1�v�K�ƷR��
�.�KѭQEQi��D_�E�!�Yqݠ�u:����v3�i� ��{R�j��Cܩ~�4t@s��㺾Gv� ��_�ۧ�_X��,�Ks��X�r����kR�؇2W�Arw�>�-ޙ;7wvԂ~� P�k�}�+�w^�|���Y��G]�z���κ��ā$������h��U�k���{I����k_G��A��PDGv�Z�m?Uދ���kw,^�2��̩�SX����u3�u�����ڨ��i�+� ����b�N�����e3��g6��� �=G%ݠ�=�XƠ�g��2	8 O���|V���_!"�~�������̴���e�J;�'��u~�}�Zf��yk�ה��A2��9�i��kn�w��-���];�lc�\
�ړ0n���-�g�����Ito~wW��P@�� F�|���f�SdR�a�9%}�0��Ӣz����_�S2�fe�q�K�[}wg �Z3q{:XƠ�{�����?JF{���2���x:�U��3��7���-��K�|q��o�!Ǟ��L^�^�o��}������}`��q{U9.a�4���<޽��%z�T���Y��D���C��k�:ӫoj>��{'����=�]i�<6U�p-��	���. �ݠ��Ԇ����j`uRPd�����n��h��R�X��� ����n�n�7quq���� �*�ou,v�"ov[���ށy?a�y|�*fu�k�;MU1 ��|}� �����	��mo�={����jip��n�̚2�v���-Ύ��87\p=��@`�ۆm����e���l����wi��/���G<ojiᲯ#�mq�^�!N��9@0��n�7k��EJ�����^����9��h}�He�c3��r���K�#b�|wi�vGW_a�?v�>����.#�.9�Z&e���w�Nb�sl{S��i����@)�"7k�����H���{�צ��V�m|�3iN�!����^�M=���[_w��P_���y�j����r����zLA��*�Y��յ伨ʲ�9A%�<�nʂa��)��z��ݜֵy��%����踉��Zf\�s(�F��eg~��>k�4w�=�+>e�U���}%w�_��|�ݯ�;�k�}���r�?Y}~�e�icd�n��bݘ�I������� h2�sn��V-v�L��}�D��j�F��X�,Ժ�7TĂN�UY�/<k���P|�w/��n��;���v���q�y� A=Ծ���8/|����p-������v�dk���~�A D��( A�"7W�����s���qm��yW�Fo�>�k�1��3�>ʸ��U��W��%e�\��b�: ��/$��Y�u�uE���҂"�{#=�yy�@��7��U�\ʴfe���=��O]g�xh9ԃ�\��z3��{6��~7�q}�C�nЍ�R��O7{�cP�`��ы�+��AƇ�*D܁�W�Ѽ�	��Yy�>��}�=i�����[Y�;=y`��zY�����(��=�|=~?�����3�<�*�ћ��):�y��vuɍk/�V-���q��N���
�ֳ-mlW�tsjCJ� �&-�=�H��Ѯ�.7tG�v֕ی=F�h,�unU��[C�N}[�!���c��$^G&��+�wccuj��)�������I7k[uJ�+�3O<%�#-��4KM�U�\t�]�F"��,fvGA!�I�˘l�������
�C�ם]�ߙ�c�EƁKXmE�"��g7�]4��V��vV��w�7��2�e}�l�+d�Q�����f_�_�=ާՍz�#�ܷ��feL��̢�W�/X���(p����=_<�a䲟W�]S	;�>�NA7|J�����ϵ<r�X�,}�fe�2���Oɸm�O��oE�z3��{6����	v��-�e��rϷ�{9�������P
4#Z�|@�_/�oA[$2�X��7���@���[7��>������U�eX��E�L�-̣��g3^މڂ>ܗǧ��W�+,H$�'�A A@���u �A�f�u�7�*;Ws����Ü[:��Sf�<guډW��5�5z5�]F����/r�G|�̯�3*�=y����:�a�����zv)�(0A�A( A�A F�������o-�Uל�����7��:R�Pߙ�C�����x�M�To?[��/^�k�{߫>pS<�#̴i��`�x���L���aq9ۗ���U��^ӽ�i�r������Xk+c�=���է2�����e��Z9�a�1�p�hо���o��hVX�I�}��v�����_me���`���E՜�\AW��R ��-�^�A{Sη���`[\A=A}������c<������̹c�,L�.&f��}�o���t����z��IUYcxi�r�K��G=r�V��Y���VQں*��r�\���Α�6��d��
���Ʒ���C;z�z��E�n�"=�#��c�E�3P_��%E��˫�$w�<<��^Ds��=�-;˗�r�V#ʰA���n��^��{�|A-�^�A{���^́m}��"��v�U�]Op��,ݻ����e��w3*x�&*{�_�98����`�b���s�Y�1����w�[�Ջޱ��[9WA���s������a3��!��[���S[ў���h3U�#�\�2��eLʞ��]׽�����'�E��� ���3�O_uj>��a���$�;+~*Ώ$��jv�~ݤF��[�����w�K�J��{=�%��W3ӷ�Η��:��v�s(�f��m�h��q�ρ���*��]�'&B���r�F4zѷ�9�3�)��Ř൧�����ܠh�/�k�5�����rJ�&�`���{��K�˗�X��U��H�h D��۪�"S6����jq�HM�t�������u!�#w�ۜ�iߦ`����hq|���G2�&eK2�s+�}�>�U�w�޻�ԶU���-���A=A6P@��Q�-3,������I��>7�w�|~�_,fDv@�9c{��r�A~��5�������&���w��L��NMk���B�x��S38�y:�r}~:6���n	g�\`W&��Q�@H��o�Ut�{~�������b#�U�eZ.e��e��?|����V����]c�b����W�C���@ ��7R���m����e��R�ub�$wnkY֝�蛳et��8�A�7Ym`��ec����\T�u";���ݤ �[��9�WO{�lk�ͧ�޼�z�.�P��\�h�#�e�e���E��+F�o]�\G�����3��8NX��w\��3�����-.���(���X~V����,G2��.#�s~M|��7~m=�]� �y=�+ɉ�����#�s-{������Uit���o�7�O��	+��[���*�WO{�lk�GQi����ϧ5�{��C2�5 N�F����򹗝�Ƙ{�>_/�:��e��u���� ���Z_� ���p���1�S��!��m� e=�����he,}��-m����|\j=�����y,aE��7��Kb��x�ޝ��wt������RyH�Јˣ&�9���Mg4ڠ0�ͅ+�Cp�1�E�k+M.�v��J0m�!d������\���оBK<�Ψ�0Kcka0f��c6�n���tm�V�q:�۫���[������)y�#�R�w����N�q�Çx�awG-��P�c��s�<?�f�N�=�>���udps��ݐ�tR���v�T)m������.��;)�飸��c,N-�F���L*1�8�k��5:w�{΂ �5��uc��=����&&�9]���k� A@��۹��0N���cS��5/�_}0OR �������+e*��ٰ-�=t8��v�{؏�;�_��f<�"D �A�@n��u|�Z����+���Op��z3�3��W��Ϫ�~�neKʼi��)	֮�c���n����� �Ng��z����P_�+s�y��������߷����ӿ����wk7$�]uY^���X�����?s�6%[��[6���s� �� �Au|��WV;w>��|N�Q����ю�����>g�zҙ��ˢ:^��Ƙ"]��56��B�D	�� ����K����}��$��3��ۑʮ"��3�,���N@N�;���� ��Dj���e���W8.�h�{��W�LݫٛQ-�=�ך��)�[��q��m�;�"��݃w&�,�!��d{쾼X����{1� ���}���J����)��3ަ&�9��9A7gT�wUM};t��9�s.[�W�es�_,�i�9�}��^��J�{�6��?����-̢�&e�gŝ�{о׹��j�Oö�Ȃ ���n����%`���܎Uq�R3��Q7�\��*�G��L���,�̣/;��)Uh#|�����ܧo��z����?!���L��w�Q��P(��A`j4�S��55D�Ü��3�=y�����Tqm��۫�K86Y�s��G#�juk��΍6�y��\֣�6��@��E��$���hi%$9�j
AI�
@�(���Y42���-G>�{?/���g���w��Aa�.��I!���7jh���H/$�߬$�0��pY�JH(P�r�$�) �9A���%��\)�L������-淬]�$Ѥ��r�֨��Z���I5���w�{�x��?O����z�O��*2Rw(CI) ��/��I&�)���5z�~љ��^� �u���h�W,5H);E�C�
W9`i ��0�r�I ��r�$	�a��_��o���Eؼ����Gc;�9hW����Ґ��o���7.��-���pW�Uڈ�ܚ[����H�k�|�������P{�Ϊ��;�SO�J<:��`')GRo��(~��zf����),Ӿ��0(G� <��_�w��u�;�9��}V/kU�j�r���t��Y�b,b���=Ӳd�-���3����;u��@����koV�� 2�6=�k!*:���/#1�_9�yon�a�<�sn��YK���ָ�}4�X����zw0\��_}�gi�0~>Ke��+��q��X0�)K2-����"��,7���p�����x�Hnp�I?|p`U���}���B�r���c���v�h��qz�f����P���)[�i�Z��^��l�����3ۤ���o�>2r�&gjSͲ,/��X����U귀��I�g��w�z'�����%�<���z��̥=�Jӫװ����&%���ʞ�}�ry�:�a����Cwc���TO=&��/.�О��"�Д���A�&���Mg��i��`C��m'K��.j�b��R�|�l*Sr�c�p�]ךU`�"�a˲wl<o&��`���ڳ���v�(8�gqiDj��!�G��i����Kg(�>�k*oX�/�|-{��hf���7fw������w���A�'t�����`o˧�d�7��8"��Z���r=����lR/m��>��,z�������d0T�`�G]������:ˣ�����.;�⋠�K*ʓ+;+8*m�[��+:��ۭȨ��.m�\�Zd]���9��ܬ鵗%�7r�;m���̊�����Fͻ(ㄣ+�D��:,�\wq�[n��wtgYݜYM�kZugq�M���̶��,쬭m�A6m�rgVYgrXw��,9,Zm�ʹ��4�4�j
m�b��K:ȶ�6��el���)%��l���Ύ8�u�jn[�68͵��6G�N1%`��T�j�K�BN_��ew���������q �}A���%2�n�\)�Q��P=�- �5H)�P5D�Ї/�
H)��9�- �_}��Wf�����Ԕ�Xn�p���PB�=�-�L���S��-��?o��;m�~�H,7\��6�RU�Qi������w5^����䂛@���S4�I
�(�AH)9��H)�+�
d��H(��R
ACt /q������wֻ{����'A��) ��߿~�k^�i����M��
���
H,����@Z��XV_�B�
MR9E�i��Y)�Ct D��{4��[����*�!�('�v�Ѯ{%]�5t�e��6� }�B�����m����Õ�ͤ�P�E�C�
WXH)�+�
f�) �Qr�$���W������þ�
w��4�Y9����z�f��Xv��I �a�Y�����AOz���RW.�R
9E��
H,�����- ���ڬ�w���]�ۺ+�~�$����i �y����4s���~g��g���y ��r��i!U@}�ZAu�R��I4�L9\�S?_>�r��?w���O$��H,=RAN��- �i�õ��L�e$r�H,F�
s��D�Ї-���$��:����u�V%�[Ŏ��Sy��u�E��
H,����@ZAH,4e��) �Ѕ s�[&�I��)9��4��Xr�a��AH{ƽ�ڧ�;�3��R
ANϷ`i ��)������
!�Q���տwޮ��ޮp��xw�Ă���$J����
d�) �������KO<�v�f�^���Y�I���#�5=��~m2�g.��-�@�O3/�4M^�0�����W��	���AH)?v����_�/�
H)��9�-4 RAe2Rs���Õ˅$���Ql��f����睞H,�e&��-G>�y�g��g��u��<�Xn�p���P5�- ���I(�$ЁL9\�S4�I
C��I�s����w��z��|��ف\d�x�Y��5�i6�*b1leh��a��A����Ζ��$����SV\)�Q��P(�l�A`i�����Q ��9���$[�˯����#6~ B ����I��������zN�ehbJH,*w�� ��B�?z�d��H,�I�P����Ü�F�
B�T9E�L
H)��}�����������
Aa��pY��I
��Y~��Q~��u��bw�H�'P~�AH,7��&�I��f�M$�(k���>����� ��f�pR
h)ۢ�B$���hi%$�kPR
M!H�ɡ��Y*2���-���%��]��첷`�.g#�O�Z@�4�RJ�3tZAt0) �Nz��AH,9˸,��I���F�S��І�&�{�㵷���ذ���d�e$
��4�X�$��H)�9w ��~׵���f�w��P=tZ~��YC%'���5RAa�syn߼���AH):� {�[&�I��I��- ���li �*U�Qi�`RAJ�,$�0�.ಫ��f{��|?n��) �}��H,;�k�������\���ÿ��;��i ��w�C) �W}f�CI9��
Aa�]�H)������q�����^R��Kܕ^���w�+
U�32Y����k}��C�˻	R�/�-�4�J���LQ�w?vϚKt�ې�}�H���}���":P���[�mL&�j$51bl��&B�XюchJ2��	�R�%����ۜ���1ػ���F-֛cr��""%q��*q<�eĸC/U�NְF���1v�qŝp9�*���GkV�*�;H�m��90��Ѭ�Ɖ�k���<�0�[�<�仵��z6��ҋ�ƔF�P���:Ⲟ���Z�A�U�9mw����m������ڼ�9:�����\��X�c�ܗ����	�̣v�S8��$��{�l�%�t��JM�����Xw����P9�-����Y*2���-��=���oy���w~<�Xg.��w��?i���k����R
AL�l$�õۅ3c%$(C��I��RAL���Ad�SW.ɨ�H(w����۪�É���AN�֨��ZC�˅$ў��WO7����:����@��ʌ���i ��_�B�
M��Ql���p�X�];4�Y22��P������݆�i!U@g����I9��
Aa����I
@n���'�7����]�]fA������w+���p��bAN���!���L���
d��H(;�4�R
ANr�ި��Xr�p������Qi �u�~�����>M��-	) ��_�B�
M!H�ɠe$	Ct Da������7��0˙�q ���
C�P�- ������c�O�ӻ� �AL@��\)�d������
AH)�Pm$J���\)�L����Qi ��(W�w��}̣�T����� �!���RAMNs;�k��t�/�z�w�@��i� RAH)�P��%$e��) ����Qi �he'9@Z{�W��o�������@��{vki8l��(n8��۷`ڲ���ƃp�Z��ի6�R
�Qi��
Vz��AM SW.���P��9F�w^��v�~�<���C
{���Ad�߽���߶�u}�7\�S'�) �V�f�Di �y@jj�)�+�
H)��9�-4 RAe2Rs�����	���y�zu������Uf�����F��x�K"���8x�=��j6o��/��\V1��'� >b�\��Mp�^�P���Ek�xmy��3�Ϗ>6�R
��l��) ���@Za����7��-L�8��?t���U��i��
T�$�Ü�[3����}�i �{�ZAa��$��4��%2�{�d�e$
�,�A`hi �9@kTAH-r����myY����??}�~ٷp[�&�[P����9PD~ 
#ಆJOehj$��¦~�i �Ѕ s�ZAH,�e'9@Z��r�N�
A�>�����><�t
ʄ��>�,d=�!`��� �~�:g{�sw󳞀w�a }�	l!y�u�����Wgu��~��y�� �<4�S�j�)�z����)���Q�
ANr��5RAa\��I �s�[&��3�[��w?=�H,�����h_��Ǹgt�y��u}ߏ$ʅ���Tܢ���I+��4�SQ�s�f�) �Hs�i ��g=�_}���mY�}����ɲ��G���Ki�e�"GLm,��Ƙ"]��U:�j趿CI/t�i �S)�{P�M2�
~��
AH)�P5D��C��i ����}z�~��������:�^����I�{����k�����zM'?P��RAaG�p�AH(�E���S��-�RAa�Pi�AH(��]0) ��<ｻ߳�߫��>H)�
a�T-����P�;��$���|s������c�C䂞��4�Y)���ɡ��P(���A`j4�S��=��f�����R��P�AH(�- �m����- ��B�
A@�(�N) �P2��� �u���������Y~�e���k~S7"�=5����ɾ�֫Ŀm`d�9��11'�Ep�ݸ��n���<Bv������὾8p���,>�����}��3�u�����$\�RAH@}�- ��
H)�P�SHÕ˅$���9�4�Xi�$�(H,���4w)�~���W
d�) �W2�$��
{��D���\) �����^/�{���]y��P=tZAH,�2Ro�����Xo�����γ����q
@�Qi ��@�JH,9\��m �*�r�H.��I(�,$�Õ˅3��������IĂ����N�_��������qÿ��AOz����%���
d��H(�Y����I9�F���ZC�˅$����z�U�~�c��O��#=찬�k4u��Ze�k[Xi޻4�f;4�9��K�j�ZZ���@�(��@���d�����II����RjR9E�i��Y(I�P�o���:�;��2%=�q~M��>
C�#�o5����E���
o�i4�L2�p�i��
!�Q���C
H)�Pi$Je0�r�L�����E���{^����$��
{��Q �!��	6t��+���ӹ��~ B �A�
H,����@ZII��
H)4� s�[&a���W�]�R
AN�	I��,4�AHUP�- ��
H)S��4�RW.͌��P�9�4�Xg�ں�����~�/v�����h���Gu �X}^�S'�RA@勤����ANr�֨��Z�r�p���@�r�M RAf���Y��J�hpII�r��RAI�
@�h���Y4�Nr��s�w����[�o����ǒ�X~m �n�H)��#��UKT��kS�B�?<��L!�D���4Ӣܾ�4�^��?i�i��5G(�%��Gf�ھ�u#���@J�>�>�s�����
 S�\)�d���D?�Q���L) �9@ZAd�)�+�
d�) �g(����i �9@}�߷_���������)9����D|	�wr�}߿
~�g�@�Qi�@��ʌ�����JH,+/��I �s�[&�I�Q��n���\f�~�M��Z���V�~P(ܵ��&4%��9җ��C��9�۩��s��V����Xr�Xq����T�E���SGXH)�
a���JH(��Xh��~߸�^��5��+���=��i �k��[���y���?0��
A@���4�XH)�P�R�9|�RAM��Qi��*2Rg(CI) �߹����u��$����d�e$Je&v��5��﫦z�����~<�Xer���AHT��Qi ���H)��L9\�S5����}[���ߛ��H�0��I��RAO�A���%���)�C) �W9f�Q�����TAH-!��
s�~���������O�8zӏ�y<&��@�">�,�2Ro�����
���RAI�� s�ZAH,�I��-BRAa�军H)�s�kg������^
H)Gy`i ��)�+�
f�) �Hs�i ����~�q�y��[����|�Sޠ��Ad�S��$��⹼=�ד8q �64�Sܠ55D���ۅ$�����h�R
s���%$r��RAI�� s�[&���gկo�~�9��RAd���eh?k�����{�Y����~�y �����
B����ZAu$��H)��L9\�RAH(ir�$���w���#�<r��Ǝ���7�Ϳnn�'������n�_x���m��rCo�a��s��������^"��k�%-W�5n��}���?�@�5T��;��j���¼C����3��q�n&��6��]��E�X�]s�p�96CP�bf!p��p1w=@��V�^G:U��ˇsƮ��T�2TB#m�z�b��<�jh���M�H֑��!u�Y.�Ql�P�0��!af�m����6�S;%�'h�n�^�il�È��n�!tBYA�������uadC�.5CP�,f=�������	2ӦE�<�ϧ�������f#�k)J��6�,�8R�A���%)�+.�R
�{f�
AH)�P�RW.�SS����5��������s���z�O�$k�e����UU�����M�htII�z��RAI�
@���M) �Te'9@Z�RAa��
CU@s�ZAt0) ��x��ߩ-�}y�1 ��\)����P;�- ������~����}�a�C䂝�i���a��p�MFRA@�z�$�H)�P���O���=�� ���
H)��H�E��
H,�JOܠ-$��Õ˅$��R9E�i��Y)���h�u{�[�mjo�����pȔ���|\���AHUPr�H.��
W�`i ��
a��
ACQr�$aI9�!������^{}���vy�k�2c) �Q��I ����
Av�/�
H(�N=����~��?  WPD~��RAe���i ��������V~�z�
H)6� gh���Y42����4��Xr�a��
B��9�- �`RANr����)�+�
f��y����Ϲ���������h�Aa��������_y[;�$�?i �S)���
A@��Y�����ANr��j�)�A��G��zW~�����zÛU�]�����ذ�p��Xıt�6������r�I�4�Wu�)�E��) ��P����XWo��I&�)���5I��Rs��k��{�k�z�����~<�Xev�I!���V��߻����i�`RAJ7���AH,9\�S6��P�9�4�XhRANr�Q$Je0�r�Hj���+O�����AP�+e�I��31��s;u��l����ʜa��1�!�5ٴe�
'����0*Ջ�74���6Vm������'�R����~?�����f�	�L�����!��{���K�F�H�8��A�A:Qn��u���̢�||;��(���~|�s�Zf\��X�9�iϷ�=w)�zS��@�_#�[]���ֲ�8d�=�P �P�5�x4a@�1�`��b8�həa�]�Υ}�ש������rO�_p>��9\B;���3�(����䉸��A� ����2����#ۀ�wd�ӂ�Gl��Ԕf���xT��M��8��e�:�{��;�s�J�,9���,�f�g� �����)�4Z~�i�������������A3ijz�[j�)L��@��D�nc��3�����喟n勥�#uF��|F֐/5wq�T���Ǻie��<7ׁ�����h����|�^c|������]��RV�g��r(*��J6��N�{�VUfX�[�5&����|^��}����6i�����#+�@�� ��H�P��v�=�U8T�UC��h/��(���6�fS��s�J�,9C���*f���,�{Z6&����ܱ̫fU�f\�2���,!O�
�Co�5�l�՜2T��|�"G_Qb!��ne"fY�e}_>�^��m�� ���B������k�:�㹇0t��mn�X�L���4a��e��=��F�|���{xs����p�<&�ew�e�%������_ y���K�4꯷h/��//z�Ϥㅍ�(�A|m8����)+�%Ǌ �$A|F�߷����N��:]i,u�hǽ���c7k���@�+��
�>��n�����!��u��x��G���lD̲�2�B������a���� �#kH^��Pzt#�[2���?X�xj���;���_�c��ʺ�m?(#F�z�
D�h�zi��HT���c��'+�n���5�Vo+�����V#�\Lr��Qb!�e�k~8��~������_J�lSa�)+�' �><QP@�����#2{��ם�=�UE;���Y�u�ە�i����N3cִ�K�v����)j���U��VDfW�ʗ2���ѯۋ8d�{�}ޑ��1�k�x�#3,�̻m;�w_fٞ���jcK���/k�U ��ĸ�&�eq��C�! wk{��u�F(<ʴ�B��ZfQn8ؙ�>�Y����ۀ���Ix%�(p><P ��2�߅4f�N��}��>�!c2�h���v�ۛ�l;=���J��a�(o�??^��o�D�C�f��n�@����/��k���YK ~��]H�~��]�w��Mzeq��#+�@�֌H��P��;�"U����:vjo���I�탤�t�sޙa����$	��"��
�5�Z5���-�hx�
5�-�^���h�D�3j�u �����ط��~��Je�&wmk��5�z���,���9�A�C��Gҝ�;3-��h陋F�^��ni&�=�kVk ��>�u#ZP4]=Q�Z�X>Խ�\�d�^MP��8�/��;*���ӓmj�}Ӯ�+Wn������"����<n���oy+}uЧ�J�c��՞DI�ŒJ<�=�f�AH<�'�aU�L)�V+ӢQg �r�n�w=�k�=�u�����[��*.ut�K\)����<���ٱ�J��;��H���nVO��TF�vN�mug�|�\����4�}�s�Պ����_�&zj�3��v����Yi���c�`:��>�\�{���ި��a]icP���cv�<`���1��u��:�{=�}�x�p5���]��.��X���BzLㅜ\a�[�q{s��k����:ҭ�ry|�[�����1a���Jr~Χ|�ܘ�MS��f�n�eE�t��^{� Œ�Ni��qe>3T�)n�srͽ���,�"�Pg�:;b�g���S���>��\�����F�h�+\�_b�o�S=.�=����=}�<�o�����{�j�R4����%��Oh�x+2��6�J��l����{&��i"�3:fv:�JL$��n<������g�q;���Z�S�΋p_]fpDimpsڸ���Y��a�Q��g�_M��}���q}5�p}1.���1��0f戽q�:.Z��������f$����.�")�f��H�:���ݶ�lv�++f:;�:�$F�D8��8;;3����Q�����nͻ&ۑ��;f����rC����M7m�i[vYc�;M�ۻ#���D���1ݶ��h���rw9#-G9ЖMj8�D�cm'���2٤ �M�e��ؒ9r˛YkZ���kfD��f63� ��fA8Fۛv��-�V5ncZM��3�+j��r��f�3q%	%6�R��B�[`�I�v�l�vZq �m�F�	e��f��:���e�Vś6�P�l�g�4��M��9�C��
���2�%T��%
r�B�Yh�� 8�lZ�d�t�2C��^=����s�A�4��`��@ν�յ�@J2���P`�(XK�6�Y[B��P�ܥ*���R]���۫!��)�t��r��.��`�b�Gk�s̝2�-�Yp[�f���ay�ٌ�F��s�d����.���c��Ž9��sˑ���z�V�mZ��N	�;On�`uv<B�t`�y���M���Qįd�d��@�4*���BX�Į��QID�p,�sauM55�]`E掶���>f�c���<ۮ:Q��λp]Sڭv�'V�/���
�X�`7;[�\�98�^źQ�z�.��u���4���N���cث���Î5��j-�P�X�m�RT�F3YH�Z��n��vl=2�5����mmTp�l����Y�K�S�%�qۆX��W]���6�. �z�w;q�!�ۄܰۇ���[v��u�G*Q֤�U��;$%�P�k�sն�H���Zɏ7A�5���%�lۙJ��+c-�j� MTĺ��k,����`�n'q�b��(lt۝�q�G��'��ov�+��&�Sv.�q ѳZ�;w-�"��o��.�0���4��/
V�FZ�ԣH�!�NMu���/������"q��t[���qW���n{d���Z���p�JX��6caE�Sm������vg��s���"�vѸ����\�M�eՖ�Ί�A@����&w�9"]suf
wS�#����	���JjK�!j�^ת�ѱs5���.���ַ�����`M�X��o�]�K�j��{S�wQb"����ˮDZ�cpE����am�훷��;!��-q�n�Z��=�rd"�ί��yԅ34�
�Y֜NX�UPl�E�;�n 5�/'K�9a�]َ�K��YO[/1�{��W�f2�q��/$�Y2v�ݎۣ`�C�F�:��t�<X�F*�
�I�Y�k�9�u�rtj����݇Rks7�����U���������;��v٪�M���M���J��j!bu��MbT0�)� fjk7��j��lW3)[��<��s�=��H�1u:�k+�x�3O9��Q.���q�ь��n4ܘ�}pű�]�r<��|�x-�r(q9�'����]��kXOZ�l�,sKc�m���r���#�mV�{��mrDԏ������[.fһZ�c���O�@�,�M�
øln���8��^�^�e{D�z��tbӏ�~��;e�m˚����G��}/�'��1�O����@����i���_vT���<�^�4�K��m%�z-�'�p�R�0�7��t�2�H��E��uFj�}�H[w:w��N�G5��U�����k�+��Αa�@n��t��Š�%8u�^�� ��O�o��owy�x%�;�	���k����1�wu�M���+�ne[3*c��s*w���ҕٜ�~�̃$W�a��t8����> ��Pc�6)��3��:,W��U�����fp�9i1�M�8]��T
%�	l��T,�R�9Gv؉�Xf|�Mg+
��������FP���\�)UM�`��`�U���bc�S2����������wx���(4oc�˻�To5�A����w�B��Y�˝_3��u����3�<���9h[1������?������3�X���|W3������Xs�'Ǌ��: �ݭ�|�,��}ݩ���i���զ8�9�b!ݬ^�Y�n�s%==���$W�a�q��X��l�㍢fYbf\�n{{�^�ǬQ�D<�!ľӤ^��ўo����5���}��#{�wo$U��|o�h�{S�(G2�̹�8}}�o��1��r��)�>&���Kp@�>lݢ�̹q�����tݿoڵ��z��?|���.��˛��*�a��I��.�1����@���vq�����z���}!|wi~;�������Vg�{`�8P�~�<�N�t�e�@�A:P �����ԁ �҈f�*_�x×ݞG(���W�af"Ѹߺ���5��m 9P��ݬ�mL�Ie"�9(�L�-�G2�P���+Y��Ϫ�c�{4�~�ڵ��>�+���� A���q��.�$Ǟ��<��zcn�%�-xS�YWn7�q^ɿ�I��1S'@o>�wG;�\��b>햙�1��s*٭џ�؜ڈ�Y�|2�����p�s���̬�b��p����
��N�龟?6��e��p�q��e����}�T�>;VB�IN�I}]�.�2�Nm"T?n׏۵5�Q_p�։^���������qQ��bӝ��7EG<om�t�ٻ�)t��VkW���S7E�w�.8�;�+����t���Kr:����3z���D��\N��&V32�EͤB]*kQ����_@si
��Ͻ0�i��8,��7���Dӥ��o]�}�(�l3>,S�V�̲�3.�9� ���b�9z�z��eH3�ҫ� ����;�����Bǧ����[BțA|GJ_�A��tx<ފg�w�~�?�Fv
��p?E�0��������!Xʑ5N)��]���{�)zO'�.�`ą��,ԫۍ�$#��8�{�}�������n�v��H��wi��V�s,�4�J�gth߽v�5yϮr�P��7iF�~�}�D������Jt�EUg���&<�3=�b��u	��q�
��llKr&{�������}ڂn��;���ڧ��S�v{�^E�9�Qy~�7S��(���h�e\Ӥ wh/��s�G|���U6���p�B�����{ޗ�Xr��@|�ݝ��V�t�j����+@�@�si|A��ݤ?ڿ3�+!�2�zfHM�݇�ɫg}@�}�t_i���Pі�n{�Wi���W]�<��h������N�rJ���N�J� ��H��z+/u�{�g�#�V�U��YC��3-��E/}b�<ys���S�#xd�+���Ü�><Q>A�_-���}��<��v~�{��|Mط82���<U>�j�����Y�O�jԆ���k>��=K�+�h���@��P�{!;��A�{��j��n��q��;u�e9�j�<��k6�e ���S�-Mm:���������f�0���Bi�&*���l�N�e���'P�>k��m��!�wT4��l��\���;Bp����2gfk�{wn�u$�8����G8�5�z�@Y�x�ī�&�b���A�x�Ж#���u���V��%�����ۤ���qù�34q�/���&��~-�`n�.K�. ʗ�1��]�����bU�U��*�|�Ȏ�R��U��wi]��2}�zv�5c���{�r����Ϭ�ǌ�2�3�������`��/��B��v]�.�XvzU}��� ��B;��׾�lzQ��k���ǷB=�.&�q�̳p��y�b�^���9��^��x���0�s�X���ݥ�{���]��Z�\�h#ş�׾wi.�k�O��v�7-�O|P����{���+3�e��3;Gəv.8�"fYq3>���k׫uS�+�{�����3Y�Յ˕\~ͤA*�K�>� ��O�?:M� �攍���a�9�-�T�۶���!�f���p��-��C���̠��(�B��t{NwA^��=RÜ��E4�A��v�x��}=a�}q�Ks*�#�V�{{=}�>���E���|���@09{�4�;u��a�$����k���tii����x:z��
}D�o�p�"^�ۣ?t�㲐���>W�;L���:�=ADӧی��Y^Bu����#筈�Y`��\�z��n��Or�f��G���ʮ ���}�Gv�?fU��YGk���Rlo�тw�6��v����Q�wAK���Kw����n��t��ӄ��'��i|r��H�wi�HGv�W��]�k�z >�_S��̜W�;L���:�9���ӧ��_P��x���7ν�Q�iJȢj��vk��U-9���]��[qpLp[M3am�a�_Z'NA�7k�:Fއ�S��X�x��+����J�{ys���u� _0ZwQG֜c;��֣7�41�2!g0�r��K����$��Ǌ"C�2��ԭ���Y�4X~�x��(��Z{����!9w��Ǹd:$�����n����1	�{��M�<�rm����v��m���hO�Zd�d{ށ�������בOޤ]�A4ɹn3��A��:P�ӥ|F�[��^h%�C�p����2�ߨ�5\�Z�~�W�3������si|FNٔ�4;�L}ʖ��bc�P�e#�e�8d�u�y�-�M�]/{��X�� ���Jn���mi��z�sWtf˱����c��R(�̺�e�$����6ƃ^�K���Yy]n�v��ʟG2��f��j�A�����v���9�J�D稷o[L�-3(�8�bg�|�3��<G��B7��i���v�s%*�Ꭶ\A9���B;���vWs+�u��h_�V'��B<��̲�l���p]��TS�~~���Y��J>��JX��_x��#u���;��t�l����N��ZB1�wi{.oF5-�<��gP �PD"lh��p�}�A�F:Ї[1�5<���������>�u�w]�ġ�,�ϗ�4|�&��4�N�o^�ĲOM��1\� e~ �ݠ��(������꺟�Y9��n�)V�u0��A6�a�@n�d��3��5I�����N[Hp�k�����(��i(���uRl��Z��KR��]���P��E����q��.k/M��|`�ߢRÜ���(OC���,Or�8�9�c3*ľ�Wm�vU�.�׵��gR�v�zR�A��{} Fu}y@!��N�w
�-^t'Zn�`��q�Ϯ0�Ļ�ϻ���s���py�ўε[�3���Hv���>���Q����H �98�F5�|Au�]�;u��~iKr~�h߯&�um�ЫC�|��!�D�� A���v�S�����w�����t�����[�p󹾐#;�YE�=e�n#�e=����j���`�+J���GYUߙ��z*�"�>�掶ع��RëM>{*L�[������߫I��L�ft�xR��G_i���χ�|�kZf�jduPs�qbn<wW���E�c����N7.���ǄE��:�ͮ��,�M�0�BhcBa[Yv�.!eA����U��q@�ݻ[�;��JJ݆ݤ���jj�����P�إy�!���Ka����k�\c#�3�*L�U�/���e�U�cv3q�F�H����\�
,���ǳ�-����C��#�ݟ������fR 6�K4�	n��m�b�1���=g� ����r&{y��>��A7P_�!{G�����Y����W.���v����3��wi�U�B����k�@||W��/�˼�cα��ךRÔ8���������sUs��VDA�Ո̬Ks*�'v�B��]���g
�l���@��B:�z��q�s,���,�}�sv�l�r����i{Gi�ҦLU��Y�eq����3�Q�[�=�<w�u�4�Aݠ�:B�q���.e1��[��cα��4��9��e���#kHb���d�X^
ՋH�C��7��6�R�"��å�j�F9 ��/XF�B5E^{U�D}�h�\Kʱ̫�dm�1���No�Ρ���,�2��e�;x�̲�fYb8�ba�r��@�{DNL�1����W�[�I��ʌ�d�Ցm�*Y{v�¡�ߪ9 ��6��A/��=��j�9���q(
�L����_���h{�=*d����a����_�\B;��|���z��!�_P?� ���N�?�$��}���*�n������-=J �|�����"J���N��;��!�%�p*ꮖپ�Ak�C�%"�v�g6��{63�ӛ�0��۠��	}N��̫���>8Q���(wP@�ߓ��f��ڨFA��羬��0��%�|��!�H~;��9�޽4�K嶪�B�@R��G�Nu׷W�Ng1�8�y�c+��#���݆�\[tY�|�:t��A��O��/�>{J ����~~]8�E��A6]��ķ2��U�o}�j�ѷ��4��� �%,�m�1���Ro��8t|���Ҵ��e�]�Ņ� �����n��ݯ��ZF�~^N�'�n�[���w�����TҬ<��<���h�;*?��_����~��,f���g��G��sr5�r�ћ/)fR�5��-n?�����̘����jz(�f��T�̚2�
N�<Ǵi����V*�Lj�%�C&����	s|��a�w�JxST၎���n�1���6αgh�����_��V ���[�?C�Ǖ���ܷ&䕸1���.�[�W%Ӵnr�o��F�ԙ�ޕ5Q�mP#���]��;+y�|���Zm"��"�at�ns��u��wy{��O�v�<f�Ǟ$�N�ZMf�7mvn���a&i�{64iŞ�S��ЯN��F���y�羢&],=k�'�k���nw����ǘ<Q�ϕ�d����f�۞ݶ��ٕnW �U�[�Gya��}�u-� �n������	�.�9S����{7=�z�;0�4�}�H�c��|�� 4|��~��pTpV�~�o^j@7����>4� �S���P�{�鴰�K�)P�v�����O����i�y1g�G��M7q�oC}��%���c}�����su�r�q���UyYU2å��5&�.Ky��[1��F��_&l�k�!9��ދ!t�is�Y!��SsH��׽����v{�^�1�{z�ʻ>�ևpYo�8@Z�5���bs���޾F\H�xvzv��9|�K�O��;�}�ܚ`f-�9��^L5&>//P��]Eo�3�'��z�o�`��8 3 E�E-3�l&� 6+�i���7smZ�t��fw$�㔂t��n9"%pV9f۴�R�3"\��L�,�*�Y�����;�(���p�k'
8s0�����m�9�Ŏ\���S��g[���7%�DrDN�[Y�Ȳ�9'��ˁ"[dg(δ�t����2΄�8��X�Gm��۝;�md�s�(9����\#��m�Va�l�ArLܜ!�N-�Gr��rf"rD�Ð��h���HqH#�$����p[Z�Ͳ:8@8N��N-�(�$�A
tH,�Ds�����'6�(�NVݭ�ݫn���!8!�zޞ�_M���߸g�Λ��ע/2�̮�2�Ds*�i�5�=�r���B�#"YDn�_o�y*�[+�>{J �|��e9y�
��|���͚Onˈz���U��eZ�!ڳ��w�`�7�)_�����=�0�*M�3�}n� �A�J ��9ӿI�i����R���l՛�U�f0�d��盋t-���L���u�[-������{�� ��Ծ;ZG�tr�Z���oڌ��z-�2�-�}yL��W�:@�wjc�.e��ޯ�mc��G����a���]��k�8��A�_x�� �$E����������r��9�h��\G*��i�>��~�/��㯱��~�.j�#8P&�A|�:t��A����"[�T7TO��M'�Ax����|v���9�>��6��3j3+�?u�*9�h��\?{��٠N��c6���3T�/�C�OD�}�;N�}��m�:b��Ï�B�	��l�z+ď�����>~��4^��z�s�G;V&9u3(_wPGN���=�{#�`��{qI����>'҈IC��(�"�Ծ;ZF�Rop6�rL�T��JDX�e]ٺ�9b�n;cz�Xq�i�on/Sh�5��ni�g�,�ߡ���۴�ncsg�����S���2�&!���^[(q50�A�@n��q��?oi����Q���&v�u�\���=߳�mFep �q�#L!|wk|��v��YWoY����e�㌽嘒��/t��9���uN�iD$���("�&e�r�,s*�{�Y�׫a���r�Ck�Fu";��9͏�fJ�� Fu��󹦽���6�b<�-3(�8�D̲�33<��G���_r���*���~co��6�2��q�6����ڼHl�5P�>�a�QҺ��Z�	g� ��dxYŻ�� /�\Nx����ʁ
�ߦx�wt;�-m�<��Ӹl�&3�?�=��i��E��H�T�B��+i����1��RiG2�}`�Z1��1����qZ�Fу�8�6�(;u���>���O�-���:����b ����{a7g�˘Q������^����0���^db���pZ���V7@����CRdu�-��mp��^E�y��ɨP��]�Cf��r�m�b;Wm�$�B���\V%�o������ǀ`m��bf$�#0K,&�ٲ����\�Z,��B�-��y[?_ވ�/c_i��A�C<���v�5�[�Q	(�{�����V���	�ܸ̬K�eZ1̩����'־]_�'_v�F��N�7M�&�9�@�#��}�}�8t�fkg���i̲�Ǎ���Zf �Ӥj�W�U�zEy��s�j��:������U�&WR�ʖ�T�f��3�4���B���/�:Q��nuK�e��<�RĜ��g�/����;��k�q�����V�ʱ+�O��{ꗿL���6=7�
��0�z�Gݲ��s,��k�̽}ة����s"s[xy#�۷~�X���v.�<��^b.���b�qZў�~���%����5�><�~�^��!��n^v1ʋ�z��{�Ѩ�������n���_Wʹ/�-�+�uQ�T����*ݓޏ��c����I~������LfM�fy9NJ7���g�n�s|߷<��'\��ʓt%�{�kt�,�s�{�s����}꧛JX���|Y_\�,������f}�H���j�%�"t�͵������U��:�L����y�����@�_�A� Ye~��`7�9g�=��n��dt�ds_/��E��!�o�n_nV��E��K�*`ј�����q��g/�Υ�!��[hme�)���=�����ړ�e�����bN��+�rX�Ch/�t�}^����YՐ�&��%�Z���AR�B�/][�:T0�[\�V��`K �
�>|~�,��/�!�!�VA-��s:laf�G���Π�&�ykHU��L~����<Y@��Ci,�<�')l��W��{.xO�q|�;P���ސ�I�7/;��E��w��m���6���/Ԉg��вh/�,�m�L��!��!����J���g�GϟO.6v����X:�עC�,�uT�����v���B��0���3��wI6y�
`/<�d�=�\>�c
X���!�b�m|�?:d/�m_�b�.T�kgm�©�g��X?�ngM�,��Q�c�3�_�]W���*�xp,��_�6�YD6в���_l�B�W���^���E�w� Au� [j�?7^&���ݥ�e����S*�+�@�X@՟��]�h���p���k�������EiWUW�+��3o=B=�٠Ov�,��m�s����|}^��' ��F�T��N�a�"l�b��L��m�?7H��0�}j
>��p�/�󥹝3e,��Q�c�3��~�Y�,��1潃�y�
��,������۱��|]27�`��=����{��=��q�W������[��~����;/�el�%� <a���θ3����{4)b>��+� ���O��Z��S�U�5�n4��]��1�љ�]Ӿ^�uGf�>��H��X�ܿ�gSvx��+[�5<8_3�/�m_�� At�@��{�o��u���r�^R�v����{e2�F��}܂�P ��k�Aw�g�ݪ�8P"�B�5t	lZ�kf9v��`�I�;��g�;Ǝ._Tk�>,G9b�!���L�o\���}7+�=��p#�[��3w~��Y����[����[h	���zt}��!�O����ؿ�:��s�7��Y�����(d�,��Y��U�K���c3������ĸ�U�9��/�����I�l��f�vO�\�8q �܂,��m�`�GN����שb̮:|A��ł;���2�}+яznU���fE���}\n��&k�dx��`��-�!��[hX�Y�R����Л�����nyf��#���¾"H��Cu��#݂Z��ֳ&��"�.]V���y�ߘ>8o۞����h]��8)?�ד����<�"UDR{�K��p9{}F.�G� >ym�-��#�׀%���u6ja�����)�ӭC��˟Y�\�ȰiK1�v�h� ���if�b����e�g9��qj3��XX0<��q^��`�iJ��IP�̛��,�1�pixƷ[��g������`2<�3�ɹ|N�� 8�ͻB��J]1��1Yh�]�b��`��W&��v;��ڸ��Ϋ@ȉ��|��c�u�ܳIb3SWk`9e�C��؜m�3��[��.i�k�,���2���c[j�%�_n������;3��U�z���u�R@O�Wг�m��@�Y@�s�l�ʫ���c�F��:��ƾ��ǽ����fE���@~��mK��~$��A>)�#���x��^�,[A Ye[v=u��V���pcΜ\3��{-�,GC��?/��/�A|~t�@�ՀD,%W��9�G�}�H�5� ��wbM���9���N�/b�cz��Gu #�X��Ct� ��_�7�{pnXI��ƽB�o���{���mFd\~ޥ����m� ��N�yd�
���&�f��0��t���eGyZ�z��5�*<��l$!WK��F�z��E�~w�wA؂!�@�n��I�fz��~�`���N#y�^ԟ�i{�4��ď9E�9��E�*�����*p���X����$�8���o+'�����9�N`�0f(Z�h;��+��-k�Mt�s(��}�����*Y[�9����Y*��Vϩn�$q�~'3�ڟ)��>q}@����͛������a@�۱`����dv~ڇ/:�E���������fDJ�A���m� ��|C-P��Q-�S�~����A��a_[v,n>�.fy���-�<$�	�=´+�[u�v���/�T!ڰA�D��~m�g��zue���K���{O��8=�����|�>��۱W��ʽ��-�@������)
��q��ԝ��ŹzOWg�1��h�a�,�ÿ́L��������#:X�Ci|C�B���{&]p��fE�*���F�?r�A�!|wZ���2�-��^�rX僁Å�X��{��u'�/-�,IC��(\�,��~��=~߷�V�������B �ՐKu�ӹ��yw
D3.��l�/�=�3ЍT|Iy'���h���s��z[��	���T��u����>]���|��$n9�����djgP ��,Gr��+�mذCh!����k��� �e���h/��E�܋0�{_�Q�~;ԁ����n��|w9_�� e��Am|�=$����������}�*<w�w�į	(q������C������S�����>~�S�S���k��KT���qf�1Ieβ�T*�JBm@�
���~�z��P�[j���-��I'�}���=B�}��^���@w�� ae�@7��?T�`M��r��`��]P��r-=���Q�Aޯ�����Ϋ�9�ōq��
���H����Y�̳� ݏz�6���~�����m�[�$� �e AK�̳�m0D^W�j��>�R �8~����-����OI����F���,�es���e��wa���U̠h-�ܻ뱻�z�wlw!,�Ea����G���m�A-�+U�@��Q���=���0��rŐ��,��mذC}7
�+'ԀAT!}�_o�W�;�z�3"���"4�-�`�u�|�=�d���T�nz��<�v������·��$bQn�8v�U�l�uV~�`���A�,��!�b�o{���<w�w�į	(�������"dB� �.��ՐAn��o�^E�vO#�6 'Vo�z�<��{��@��_y�� �e������_j����m�d6���L����.��g�+���^��ȸAޤAڄ"�V �_2�(=�J����*wU]��3h#Ǌ �݆�_�6��}���xI�l�@��d�f25������m���~t�E��(r��ښ��Hz���Y'��7̽��@�����|�> �݌�'����W�<=|1�������������>�(}s�������Z�ZO{P��B����A�N�W�վ~���z{���F����qO��Fx��&�rے�fEO<�p�6��z
wA
�k}L��|���r�^]���m/_=kp��Ac�7���^�Z���Y�d�f��Y��c<y)�N��0��]��oүgs[�U��N��/�FdY7�7�牅������,��zD3ЃX�mP�o=w�]�I{o�.�n����j^�fe�n���j�=�匍�K�,�7�Ƀ�����fY������8�ѝ��q7s����nϽM^�5�\Q1�+~T<�S�l$h�+��U�ӭOSrz?3d�6��35l�ع9���A���M#�׵�/�"Ҽ�$*(�ÌB;�{$��Fm<�)z9����zV�b>�9�m����JP��[��Ar�^�qs���{$0���B=��I����p�OQ�z�ݗj^�rVܘ}�m�L+��e�N�Mn�^���=�Ѿ1��M���k��F�l>����`��#�{�^ɖ�=��j�����P>�Iw�۳>���N�M��Y�Hbٮg��Kx]̱�~JU�E�y&6e�7��w���]�ō=��zg���a��h1�1���y��r���ۈKixed���TH̘�ע[����\{�{�fy�{���StV�_/*���	��1 ��Jd}�۞���'Q���7��o)�W�a��Ԩˢ���p+g�7vc�o낳��[�cs-�x��&��h���{3����I�E9��}�˔L�98��pJ#��m� P���"a�Fr	99٣�[%�������� ��7m�&j:�ƴR�Y��%���� ���n�n'Q�kt�D
q˶�m������ff\�BP�e�v��:Ӏmh���p\��Y�mj9	'$J) ��3$8�h�rp���Q�5PHJt'K4s��mm�,�Ȅs���I (s�1��g9�f��p������'���D��;�9m���#7���BN���:9��@!�H� �D%Gmb���
�%���27"�mZ GYgrY�L�ek0m�8����hRޅ�����[�6��ֶ�a��-�5��Ĳ�1֚d�[o�[X���yi�ѵ��3T�k��Uw��K�	ê��,�����Dt6y,i؄C7HL�hp�:Dep��Y]�i�'�۰[q�[�[�$�jӲ8N����֢l�;q����%�S��F{As'>�0�:�j�,m��0��Ұ��������JEͭ�1.�Ų�C�e�8���7)��$q��xq�1��c���*�m�\�ŧ�	�dr���8�Zݱ��1�a�]ta��\�ɼ,o�Z�4r��8���-�s�Q��͜=�&�,eڔ��� �J�(0W#m+h�ղcM�z[%�G[WKy����\CJvT�X�˯`�.��Q.�.fe���̡4�ol��;Wh@�`5�bLU���j��\Uu�-`i��yz��[�G�	�f�]IU$;0�vRg��MKN^v��� �oC�]�lޠkڐ�ÙJ+3l����F��/ ��%�A��Վ*{s����lE�I�c�40ౄK��֑Ա��#Z�jMƥy�zܳ��km8��p��t^8L�H����Xsx,�+&j��P."݌#nXL��&�֭��Y�K���q!5���6��:t'��q���ۤ'�3�r���=q��#�`��Pu%n�뫶Լ(���v݈v�ng����Qƚ6xֱu0V�2�0��	�r�mzآ�'f�ZX�n^+=�x���R�Ś�;Ŭo�Mw[��W;��N�1Pn���굤���̻бt���e�6�&]ɢuk)�As.�Ev�:.c �H�^���c�9�1HqE��l�i9�ܔ�����ma��盄����}��v�'��5��)��k�6�f�ǲ \�h�Ӗ�$iXq��v@����i���]2g���Oh;Aҗ��Z�r�2k��UEW���,�`��������ݕ�m�C�n8��]�����ܤ�
d�u�9,j�#\�[����vqq�9��l���J��p��f���٭e���x���v�ٸʯsӑ����+w	�1[��n�ۺ�X{��M��>I-�>�Y̳��ݸ���9�n--hN%��u�b�#]���L4»����+Ǯ���vn�㈃�a3*u%��6��l34���`�;%՝U��l��HYZ��J��5��f�*mg��3ֳڗ6�GE����,���˒P��H뚝�F�����溵r��ujMyS[�B̶߰��s-�}VPG9b�!��!�!0�ӛ1+�ٔ�[�q�/u���e}��@���D2РAm�����������>3�ޖ-��gc������pׄ�8�Ҿ�!�>}2w���Ұ��5`�ҾA�!�V��y���yP��^�j��5�Gt��3��;�̳�m�ϐ���������ző��,�x���J�ve/V�d@d�^߬�Yn����_�T	m�[AY�vw����(��A�m��u��^{��'/��D�d6����_��i�e�����F��4��d�f�U�0�ٯS��Ę6,�\�U��m
0Տ��{硖Y>~@m��!���k=^i�@�p?�X�����b?{����nŐ�@�[��#z�E���Y�Q�I�{=nHr���gnk���O[='/>����~���y�13٨:���&Z'����j=aM������bf����-��a�o�bW��Ľ[�}��Rl�o9�ˣ���~�V'�V�glЏ͠�n�݋��]\76�����*=����+�N��C�!��6�@ڲ4+�yi8ڲ#�$k���m{��u���ځJ�ލ#i��Rh����xm��u|A��,���/�m���*�7.�,7˃gzi�w��jY[�}�z����m_�[�dU]E����c~�W��! �ԉu%)]�B#�[&M�R���c��4���GY����ȅ�w�@�@&݋����'�/3�siX��~<1�U�e_rC�����ڿ�%�@��G;�uo��}�� �Զ��ul�GY�v��
W	��/�� [�&*��g�v�Kg���� @-�	�b��� 6�:Q�xL[�jū�������M7,xK"U������s)%�2��+��<�{�)Ouo�n�7�q�Oa�$Yخy��I��V�d\�)|Aؾ@���t�!�_|D՚����Ũ �3� A��b�ۙ��|��_��V$���]�#_8v��r��9�����ڰ~n� ���ڹ/�	�rS-�1Mtu�n�ځJ����d�|�Cn��Bpڻ#�Ѣ(�p �n��,�m�x��Q����RǢ��+mU5WX�`D��'�������|�-��'����nZ��̋��=}*{���"������źD7H~-�/�K�̗�]��۔4�,7�ݸ徧3��V$�����@7��/n�~�8��|���܊�?t�!��ڿ� �X�:�3fT��	�{]����A��/�GJ��݀�*��+�Ꙟˡ�=%��|�-��l�o��_{;s�+c2. ������K�ؽ�)I�	^�������֋���E&)Zԯr{z�Ugt�����<�k.'��x�U���oK�Q�r5���C`���Ct� �аCu�t/7`��}Ṏ���357��ey̥bN@��dv,�_2Ȼ}w��%R�ѣT=�����	\��u@�m����Fn��e4ġ�KZ��m@�
����A��R�����-�^Ƴ�HN���=��)�6�vM�YH���?6�_�6��A��'f�ە��_wW�6N7�g����啱�	�K�ؾE���}�ޱ <�|�'7��Am[�h��.��߽ޕ�Kr�^ىX�����v,��_�k�[j�잇$%�ʪ�~�V�F���@7X7�άpg��{P)_p>���8�nL#�Af�Ae�6�?�/�!�`6�*���阾^�\�6{�yۘ��3"�	�_l����>�/���hR�J��D��ZI[��.~�\�'�ڽ�e9<5�rŬW���~��!�}�|��cᾄ��SLx&D;观9ެ�����|�sq�z��	��e�k#���%�`͈c�m'c�-��#G#�|.�׷�4�+���Y�"���
�-�qlXYcI�K�Zs��u�ibk�ri݅�;6����l1�X٣l1#p�3]m���e3�Š0JNΨ�0%�;/d�]�ƅ�z㗞,�v���s�H�f�$0T&5c3u�¡��ru�ݥ���8❮�ٵ�M�����[�M���^����36��i��I��tK.X����/f�� %j��^�+��S��~ݚv�[��!���k�^Ⓕe��Ԭ�' �����!UUA�=�b�#Z_7_ m_�[��x�Rñ����}��;ԅ����������+�>���_7_u��~¥С&X�F�t�b���!�"�!ڐ��*��[��=y7ز�3"�~�HF�!�V%����;>Uu�j�@L��a_[v,kQ��)+�_��U2ĝ�>(�W���������X���B-�d[���鐁m�c�.�g;*ϯT>�|�:�k�z�F��P��e��݆��7����4,��n��*�ͳ��`n�(m�ꓱ4���P��R�o�}��/���X��鐃d�pou�����lfE���x�2�
+r�J���8ڰ �K�j�m�8�e\����v����P��;u�%���*2OW=�2C�����j8��i�B��ܭ��ͺx��w	�oz�������Q��)+:_�X��$������o����z�ϥi�H��R �d/�mX �[���~���c(�W���:�k��P#8
��P��E�P!��o�^��yﻳ�����,�i|�!67�{�;۷���̋��vWޮ�rx[���S��7���җ�2��m�`���)�1�&`?VK���_�C3��2���@�p�����o̳�������g{ﯨl��Bf��\]fn��e�%3�T1h]�W@��͡F��}�z��2Yg�������+��yq8��q�n�P�d�;<ӯy��o����@�
��n�oY_ww�E�Jn�=��P�5����ם���ek�Mw���j�mN>�cq_�a�<*Dq�P%�@7Ce�-��	��/wu'gk��� � ���O��~Frys��ą~ա�%$��9���}����,�W�/wW���v�g���"��?�خ(f:�9W2�� ��D����B�ڰGYX�� �*����ؠ ��^�~���������cB��Uյ�0����@�YD݋7�ߕm�6�N���F=�p�ۛ��ג����D�@�Ղź�S�aą��$.N�ud$s��8�ϕ�y�$��C�7
�ت.� �*����&(�X � �,��m��K���:���"NX�W��/[F�����,�����Ku��$���j���}��R7��/X�ڃ�r�f��P�A�F�:C�ՍP��n����v/�&$/�"mز��ͯ��2r�f`�w7/V�+^�k��)����ՐKt��7_`%=��;�$��Ȃ.P�0����se�)�"N@�����Q	2�7~vW[���{pE���w��y��ZJ�Ǳ�^
���i��ܯ^�[���X�.4(N���d^�{����B����S[�yd���f�7����C��|�|�m}`�H���[h̷�Zf[���?��n�W82�p̷��%p �1�dE�t<��������߾k/�o�3GC�144CK����u��8���N�bLg=$�\��ґ\�+>�̳���G�����>�d 5���%���o�k�Mp#���U��{k��n�n��m:�܇O�`]�|A�b�-�.��g��{����q!�ݵ��Q?��]s�.R ��"�_Yn�̿��۽�Ԝ�{�*�X�u,���N_M�X�Ct�-�m|�SJ��IX���� �W��k�����nג���JDr�gV����k����	��o���-���6EN��W生�B}Mس٭K�u=��S�D���G,X!��.�8��E��,ݮ����=�S�;����c{��U�̂�o1�`�籍@��H��6��M�%7����*��6v�hn�S\��)r�rxg��r��&�u����y��#���C=P�Onx��[�l�y*��v拀����`��P1�	��t��%�I��L�Xxnt����0�ej�����c�\֭��Ћ���Ye0;�a�5	���\u'['c���M �<ݺ�n�61=ػW��N��;6�.�j9��䪑#Fx��gl�a��8��c;]<���5	�� uթ�I3�7<�Êz�tm�����x4��;u�4EUQN��w�eBm� �[���Wl[\1y����U+}e����0n ��Am���|�+�7sxto4_�M��uCY9��ٹ��l�Mq�%|��B����=�%����1R��-P ��/���,��-��˪��Y��ԹY�=�I�l�D��,����鐋mX#�����բmp ���5� ��/��׆�������!ޠA�!dz�����='"~���~��hYe��b�m�ѹy�˚�UXB�N�N���;�6d��NJD)��:ڿ� �W�kP������������r��WZbm����iG�n�-�:�^�j�uS�zT߷f���Y_~�[�˯d��s���'<��5��<g���G4�%�ڰA�@���uQyz��$]��nm�������]�<v~��'�ҭ��8{bۉ8E��ێ,|{��ʰ,�j���k�&4�_؝}�.?7H�y�������ϲw���"�5O|O���*]+�0`KF����nł���s�U�f{�"o/�����;�6a�p��쯛k>?7K����O���ۋ�����Ԉ-�[�˯b�����"N@�gJ#��4��J�9���l���P�[j���|A�ڭ�*DC��5K�����z
�������C�w�Ȁ�����3�&<�<�ߩ�y=�>Z2a]�gG=Wf���n��M�ty���%��f������C�>��"�X����A��R��1��9�����e����'�r�ߺ/�;�X ���"Ŷ��<X]�����>��A�_X��}U�{��,�o��8 M� �K�������^-�|-j�|$��h6�nI݇�����r�aC==0�2�6��ٖ҃q��嵩�^�/'n��A��U���Ʃ�Y���u��R�=7�8`9w�٣�5_"�oY�i!"�p��+KI���h9usM-�Ǔ]dU����-J>�2�L�+\�5/?[yrYb�y�����)��;�v�C�b�Qx���-G��{�!^�g��v�$����b��LfI�֫Û���~&�(�iA�������\>z���6ŪL'}/�_z�u��,�t�ԃ�~�΄ۈ27:�y�pb�q���[r;��!�?j����Y�a�i+hCJy�2g��/;� �22���Q�l5��}Ϝ�_{������zZ��;���;*%�o�����y{�A��g�]�y>xj}g���ugq�H������a>�[09��8k|��>ӕ/-�3I�J4�eW�ũ!�� ���\.�n�Ճ��9�0}�_n�8�lw"��X�m�����zK*Z�E���M��.8�dE��S�=��1t��ʇr��n���8f�T��B��K�}��G�������1C��On�9<ǔ�:��W2a�l��1���Q�	ۭ{Q��E8�ǳV�z�]b�HR����j�%��H�y�vh�4��"�,�<��z�;t�8������S��5D�gTcƕD�*�OS�ܪ�*GM5~%���A�L�w�#�|[�����>�������<G�uo�O�D���U@�����yu���1�(f�H���~�`a.�q�yaj\٥��h惡d�ss�5 ��.���*r�WI�w�.|�ʤ�A��0�3 �0�����f�ⴰDB�֑Α�egv	p��\\p�tL�ٵ�f�E�]�Qәݜ�ABw�֜'8��:m�l�*rM�
N$9.���;����Ȝ�NF��9,�A.,;"��I�'fq�Irwvq�ge'[bJ"��[g	vZDwm�;�	C��;�.N+-;��:��QDm�����ub�N,;-�;�l	9�N(��#�+(#�ַi$ D3v�,붵�vi����qf�E�'pN�%�\%2���NA�r8t��AA�f����rueg#��H)p��I��:�J�r��DfS�I:�m��mnB ;)��6��[c��	�P�\$JpE������AE-��4d�u��r�O\�r!қm��u��·�4�&rn����obw/{�f;9�6	8:����?c���;��u�m�����Iʧ{W{����/���ԸԾ��U�퓾
��8���o$�������5nW\7A�!)�̻	B4#�e2L��@��+c\�Z7S������|�N���>|��n��^�r�ep�U�syI��foz�r���m�:���{�R�@F�ױ��ޝ3 �͐�Ҁ��ic�t^���;��m�ا���p�����������{퓾VЛth6��L���ֲ�o÷����ыq�bM'��Rz��5��TE����񽶯/0���mX �5�K��-�Q|�������b���.:y��_l(Ƽ�ѐh�=sR~�*�����di��6ֶ�orK{H����K�7�Od����I�u�ƛi��c�s
�nu3���U5@[,�� �[Aζ7@ɍF�7n��sW]0��Et����e6�m�7��s�/��E��5^�n���sn�m��v��oF�#}Q�*��A����1&����O\��ƀ�M�A�Y{��q��"��n���zR[�՟��}�v����}X36	;�=���m� �9c^bˮ���h݁���6�ܮ��i���E���}��>:{�����M��t�M��ƽ��ultǗ�
�d[Xq=s{�4:P��m��������#���0���7=�kPx��Qx�P~��7�J��+4I�7ړ,��dv�n��i~<ֱ�sr��i�M�"2��0�u�D�/Vv���q��䆍�"m6� ��6�z��ږ7lڢuϱR�cr��p؎:�8��`�].���V�)����u�����^.����8'�#�]h���T�o`.�Z9�܅ϯ���v�fun��U�6ؚbn1uA�����rR�u%���%p����b�6n������uE�:��G\M��h������~b�.a�Cd2�[�"O˯��x�z�=���-,��+�D%�����g蛯�i���������I�N���>p^����7������Xn��,7tG�ԟ_������s��i7�w�qd�7�����Y�=�}��m�����Kf�����T�yma��Mᱯ�W͵�m7F�q�I��x�t�_=���k�v׆f����u<��wDHb����� �@6��lg�WY�u|�O��ײ����d����qq ����E�{��y�_��P2��շkc���9�b8Rc��;mIy�!��&�W	UENS���m|���0�{���OfN��K��m:��M�I_c��M�m�؛3.�v�>C�Z�Õ�����t��Ef=~������]�[����ff�\R���P_�ȰޜیT�^�@�T�U�|sCm]���M+�3`��zP����N�T��՛��_�6�Ͷ�7u��5w��n��?AG��Nˋ�7_|�A����:�3�7�� �����u����:ع�����7f�o�Eݽ܇F�������NC�{m{"W��v�7g3`����m�n��f����j�����%
�z_�V�݆����D�jk ��T����m5#,���~1}қk���:.�=s�Dz���r��E��X���<Ў�m��rw�}��:�	��vٶ���]feb{2p(6���z�ܠ�^�<�7��6�m�|���?y�x��=}�`�`f~'�d��q�&k�q��n5�!�[zp����=?yn2-���}w���o�A���P>5X����Ct֥�odن��8#��@Mz�鶡���Q5���ޭ�ʹ1�S[���"=PF��O!�]��Z�\���t���}ͦ��7@6����B��ǆ�#ʝ�>l�ۋ�̬OfN�6��A���=��l0�q�*��U>X��F��!`�Wl�p�-:�"�2clz��ƒA^g��z7��A��[����*���/�����\>����'r�|�6�ʹ1W���z�w�v�hc�[���"=PF����6&�Ұ�"P1/��P������؎Y"��\1����f�'�'|#k�қi���ۼ�~���N�Ϸ��6���ۘ���Uc2H_|=(�>�|״/{���ڽ�|tUYYJ��g���Iy��.?L8�0<!o�g��֊��O݀�Ę��wy��g�WS�/<wƮ����W�(6�ʹ��m���y4��Y67��hwa���_Y�#rw�|�ؾn�m�{|O�޸z��ԟkhfg]4v���&6��@&�q��e��Mi$�]B��E*��ָ|�ɶ�n���7u�s��ڬ{�:gN��{F��� <���6�u�m�A7�����n�ՏJ͈9wq��wm��B��J�di�2{*�Z쿩P���NC�����Y{�v�xq���Uh��swW��nN���H�u�m6��xl����q|3�������r��G�N��Mr���Cқ�����6�l�ȟbv'AWۻ;-v��tۤ7$��zW�kA���>�v�5R��r��w�����;��+ݞ#Þ�<���@w��w�'��ۜ��6��f�J�
v����طٶ���v�V�t����]���o�I�S�n7n�d�u��[�Tg��i��@�ۋ�kx�<X��Wg�XC:���.�����`ܼ�뢷��]��ΐ."�lc�wWT��a���kE�,�0�g=��;d-xNB1�9�-��Ө���'͸z�yI�s��h�'6�IK\r��5!����� c��Ζ=��k���U���a���S"������j4F����s�<�!��v	��n^iֲRG\�6���K�E\����U����t@oSm|�C$��K�����7';�*��pwju>׋��m��h�!�����������oW��?&��]d���'5�қr���R��:��$��rm����)]�^`�ly|�z\�������$u�zW�km��m�����S�h|�C:q�O�yz��PF��? �>���8}��8�־n�i��ʧS���+P{��rם�+���6d�h}ѷ�k/���;9�xI��sx��T�j@���Bq�n뗩<�qr��fM0"��U�/����m���l{=o6���CvH_	�՗�e�r2�+hG���m��w�ܫ�_����uev��r��f�և/��e����,�W
���G��ou!���d�s{����\߮P3Á��U��9��1�	5z��rΜq�ӽK��#rv?)��{�Oe*4��_���r���i��oݹ�A-�*�G�����=Tٓ���ѷ��_7Y�Q�IF���O�Ⱦ��NF�{�6���CvH_|<��re�:ď��;�D:Pm�m�߱�sZ��2�"7�rrq^�xz�e���n�{�w��ޡ)�%�fPa�q�V䮛�v5�]3۵'gfB�x�S�U��"�U#��:��"m��'��o��v+�C�&�r}���*�̮�_6�n�k|�$�x�� W�G#�=��~� �H_�C�����ww��]�}����~�y���n������%_���U'���c����h�q�uu���ޖvŬ�;��ަ����s�՘	�W�jӷ��ެ^�T{U9|SuwPK�*S)�䤷��fG�e���t�A����a�3�����2jrn�Ow���y�C�#�hPNQɈ�X8�݉�@7M�>m���Q�lou��!s7ܹ�o��q�_}n�m���qi<��&Gk)Y0�i�a�[��`��˦ɷD�f݉Q����u7C����+�� 6�ӥj�ܒ���=	v�=�g6}^����h6�ש_M0���9���/��Ow��޼���#��� ۪���oq�^S��������t>m��K�+�����{n3A8�/�hF�m|m�[�a��9^�}_wr�6��V�}֕ޟA����-��5�:ݩ��Fz�{e��A�����vr��pH�2�=^~|��{�xS�i�b���"��x��曬{���z}R���1N��4L����쯻���6�Ϳ	_F{թ�7:�=��ܝ��\>��>���Jm���v탔/|�ٕ�T��n�Ԩ��$&�`TdW[k��j����7ެ�'h�����'�z6�oc��3�Fh'n���v�/�Qc똾�� �h|�_)w�+�YOs����V��\�ޯM3�xz��ɼ���^�j��/ϟg�(�on�C�oA[���{����z��M�p�|:Sm �A�»%?�r��^���+���c��nf-��h'�^Х�){Ի����W~���:�m���t�ۛ篳�z}|վ��i�YWk}4˛�z�z/�tۃ��h��/U�vKȈ5����A����˚�{�͊�wV���o��]ⲡ����;=�7P�uts���i�l�6�o����ŗ>��;��o4v�)���sڹ/<���=y��ZAvAv�Q�LƲĹfA۫�onlZ�a8�J�����1��3�� ��}a�]>@�����e��e��n���Ox7�bg��#����y��CQ�{�i���9ؤէ����Bg��腐�G��,XR�yi�x�����ӺaX�d������9}�h��pok�{i�9>[B�ж*d�l]�<�Ȯ�y�2/��k�}���ǰ	�-h��(�<�5���5�R�&Q�~'ȧ�/Mf�����A���v�������o��ͳ7ƥɾb�N`h\�>e3Fs6�,�{qM���؆߫�yXI�;��+������)���w�.^D��S�3�k�K�`���^n��b��� �"}�4�A�|�t\>�x���¡�^R,0�qG��#�jg�{ӫ��Tny&F(�dz�Wf��W7|�7/z'��#/=���8o�إk��Fy>~,����Fמ�c��O���JӼvxV�-��^�ͳ�Q�2On��غ���ոIr���%T:���L�f�@�_��Q&�,Q�9�{����G��/n��Ώb��;�C����HAD��oo�Xf���eOzx(��������Nf:���L���A��5�o���P�E*�`��"�>Q�iܷ�g�\�D�[��浇}'p�0|;՜Yt䈧6�H�B
�+kG	��J+�����;.�K����I:#m�G�RTqtvVPq'w�9�e�um���,�� 8(�8���8�*(98�YQ�ADrrT�I�D�Qt�wqqD\ftqI�E�ێ&՗m��΄����$'u%�tt�Dr�QE�pEwS���U��rtQͫ ����J�:C�#�9 ��p㸃���Tw9�VIIQ�t�tEDRIu����:r�����B (�VA$GHXڎN��Rr����p�RDBq�[�m��<�����hͪ� ����n�%�6���6�m1�,lP�ϏI�sYu��8�,�ѐ]h�bx�<����<�El�&J�\��`֭��
�����k�P݅��fgǋ�������$m�u��rN+��v-E�sV�Nlڲ��f٬���;]�&tgmؖ����<m[ ��7m��u�&bS����Kmf 3�Ƹ����8�k3L��Z�Lc��p/g:,F�!�L$���ڱ��r����{s;�8��/l�%7X�<�e���^877��miN����k�5N��ԜaT�%p\u��N�\�z�ݪ#X4a�9%�C�9U7l�O#�.]`�֮�|g��M+�q �LCv5%�@��W&:.Y{l���t���
,�i�<&��GD�u+�:!]݄;6Ջ���Ѽ�G%�����;L�Mq���-���3�N^��ۧ��.)y�H�m�3�p'mǨ��̯��y���rs��� ;B�����J��L�
A�Bn�lxլѭ�3M1ӳŕ+o$��!���q]�غ��:�j�[�M��1��T��-���)�K��x�;>Z�t�;v�v�ݐvm�)���յ��GYᢄ��o ����nn�KTu�7Fw`�ء5M,�����c�];L۫vC;���{j�v�kTc�0s`iD�&�s��T�3�.Ӟ7�;h�,lx��q��B�0���\��FÁC��2�ݜy�c���p�sK��8�EƬ%`�q�v���5Xe	���׍ͺ�q��1-���A��n�0��F6��ή:��'��5��{J����4�&V�u4�ڄ�Q�u w>��%<O�m.�sftV�#�5�a���ڂL����/Z�����t!���چi��;9n-��qk�r����چA�]*hJa�a��f��b�u��i�x��m�n*�{u�����)qs��,h��&�҃gt�hm�b�-���=!�B�6v�ge�6�iI,6�՚7\e�f�]2�.��:�]M�l���ݧ�㷷��hֳh��Ln�vE%޺+���Ʋoc�r�m.j�����P��֢��xeNL¯u\���;&���*Wvvx�-�	E�l1��]sX7t�5=�ql�N�F�ڽ'g\�q])m����;�5/��'5��Y2�g.�֊緵A����!�W��P���磽~������e�u�o�;ٞ�<�d��B�GӅv�@=�2r���=��o�:�+Q�p�_7���f]��M�Oxm|#i����<�GP�|�vk���|�_6糛�k¯��ou��[�\��z��n���A������/{�7�� �}��ս~�ٹ�ζI�f�;��SfE�]�~��;����߻�$�������^!5���f]��M������k��`�=��}+¸�=��4��x7�luY�!�q�Ơ���tm.tW��0M_G�<���r�m�hd�3��뺻�٦)��{����O�o������Fw��i�l��CЫ�e\�t��S�O��P���Df��WU�{���[G�<1���6�0-�*hw�f�uƱf����r���޺���ݛ��<�d��z�Pm���U���V��+���߀mֹ�vj>�ܻYx�;�v\�Akq��� F�m������O� [k��'P����`���+J�nA|=m<n]��y�=C�m��7A��o�a�[zԙ��?F�����y��l�����o��]N�Q�:	԰]�W��5T��n�6;����wǛ�z�5�볍s�q���6�t�?�|���� �|�׿�zo�i�s"������P�ۛR����:4� �C��$����{��ɰgi��ڴ� �>׫�o+�;�R��6��s&}% �M��ŝt���啗�5dF��J�GUq^�n�-/��sx���{�P#ʍ@�_d�w�u�GG�_$�����ȥ÷rѹ�d���#��'}7P������u���[�tk=+��`I�=�o^˹7۴ǻH�{"�ڡ�y�Ȋ�}g7�~���o͵�t�{��vi�V?9���V��b����"������t��
񘲔w��
!vI4�-<t�Ҕ^;&'e�=�D;qL6�m�l`��l(��:�H�m|��4[t���L;$��,�-~.������m�����(���A�oz�L��1��+ʛyѴf3ӫ��̺���' �ki��3�O�%���z�j�V�b���}�7�m �@w����j�������$�7C/ڋn�NǾ���8�3�t��{����}io-2���A1By]Ze��s�bԧ{����=��r�{��=�mͺ��<��q��|x�>\���o�p��u�ʹ>m��o��'��-_�m��y�&&��쩽���4�A�J�>}��}������	��n4��#��ݫ�&�ms�
�D]*!
�$Q��(P �i��^ $���ty^�:*��������ޜ��'G�k����G���9^��L�vy���p���[M�ۜ���\��MC��l_�Yl����i}��� m�6�h�U���]��Y~�}�Ɠ0ߞʛ�{h� �@7_6��GX���C����khyǋ8N�V.��jG���*��+��C�W�}@H�x��m�<�}EU�պc.ns�Xf�w�n���6��6�i�6eDw���!\z��V<6����ɴ����OyЮ����V��u��1���kf�<+�(�,nd��O/�K~�q�LM�5�q4h걗����;p��Ԯ���l#9G�F{\[ĕ]<�k,M�d3g���7AѪ�#+�v,=/�h�����K�l]�P}M��ۧt0l�&��Q��=18���aڛqe�����Ϊ��m�1&� +	�
��� ��m�f0[�r%�D�"�2�V��loh]���3v�m�d�t�v���![U#M�������o�q�).˭f�f4�]()�)��[��{d�c���%XF��!D]
�|j�� �@k�z��w��~�"�~����:!��3�ٲ|�hګ�e^F��y=�־��p�]V-�ԏ��C����}����i�@�m��qnN�/1�UWV��=��a�'}7P�h6��~���r!Kzd�_G_6��y�����}�_�ȳ���"V]�\�<�;yͿ�������+r����X��n� �V-4ԏ��� �o�6䮼4��}}�����|�Ԇn�K6;5���7Y��KZ�&����B���T"��uE+DYT)%WI5�(��h7_,�z�ӛ����d���N���������;�m���/�x�ogS����*�hO�Kt��.���!�e������;���알q������O�.h�?z��]���g�U������q�9�;��B�M�=���M�����;>.���u�m|ciU�'�J�Y�#�V*ÃjG�}�����m��_aD^�H9�w'v���cx���~��d�>ɽY~w�n�:%��F���͵�m|�Kt%�ZG���i�!å��֜�.�l�|=��6�m��t{ª�Ng��}��e��XEH��fŘۊ��\�n\n"��6ݨإ�~B�Y^�h��A��m��ǲ�8q��$R>Y�9/u�� �hoPm��h6�� �[�s r�x����{yb�'���A�T��0��<��*��PZ���u�m�w+�5ڡL�����*�y�Q\��t|S�'x]��<����P���&�4�Ǳ���f����nb{�՛�pA,n��.PE����5����.��C�ޫ�88�}j1<E�M�/����M�>n�jz7�u[�Կ�Bd����y�����
.�y���=xk���c�|� �A�m��EU��pvV�/�mM��{b��}�_6�}˷�ߴ>͟��<��:�mWM1[�MlK?�m�|ڪq�v�����H����]�EXTH�����Έ7M�~i˴���&ʗ�n�߆�|��<Z�ʹh\cFV1�W*e]��H]T�Έ<�\�����.��C��x�5��F���ױ�@wPm��k��זU�L�V0�)�dSs���k��j�wSm �M�Ѕ��S�Ig���ڟPm��5�9ur��6E|>�\��&�����5)�'�~殺G~�G���_�)�ճLљ�#�j�%)/*b�a6G���;�{��*.�����ɹj�޷�6��x��-��~a�
���۟IM��m��ݍF���~� ��oWfW�E��$�y�7n�nr��>f�@��ݾ����a5�1�i���s�*̎qm�Mp�m��	U]�"�U#�~�:�r6�n�o�3���7F��}�x�`̡�/�h7A��m(�gۅkrC'��G4If���l���e��m��~��o��� � �C��6�ͽ]ӍVL��[�JwV��E��$�5|�o�6�mu�2i_W�`]�}������w]>�����A���隆���yf^yS�o��_փtm|�M���P�řH�Gv�ͮ�6����dW��Cy��k��|>��SZM`������v<��H�]�y�1�iܞޚ�m{Ϭr��N>�0f�곿�M﯄>�mP�ZF�f�_�*߿~w{X�� ��aL79Qռ�����k��Gٝ�J�l���v���\d;N�MٷD"�,fеZk�.�ʓl�L#�i*)D.3q�{J�n l��/���c�ι6ǃ���nN�	�u�
snKH�n:��6�2�1�I��
�3���/.����E.�Ѻ��=�zu�5a�̯�ֵ��<tF�eάf<�oϟ�F��ݩp�j�ku&�P�F��ط,�!LmͰ�����O�=2}��m������
.�#�1���Cۯ5$z15��h���ڕ��'�_t/�7]>S{��Ǡ�q��o(\��+���M��#M����uѓ'U�N���lO��d��졼�m|��@]��o�r8���5-���7��E�쓇�R�;2�ʹ��ݿv�5�������o�lD�� �Ř�B�pȜS{��Ǡ�{8M�J�|>9�0-g޸�
E �B�excc�jT��NR�hR�	J�^X_~I���^�����=tƿW|�7w>��C<���zL�}����m}�V.������8Dg��]VS�I&f[&��u�J�[n�ܑJ�ǁ��Ү�QJYB�}:�h[����q:켊\PH��� 6�~���s5
.�n����V����j��=k/�����m|,����o=�.�Uku9��c�y��2>��MЃ���vi�Q9��;܃to=�Z�ȿl�.�ٽ���kӛ1p;^����M��m����{<����8f�UH������5}N�|=r`�;�߹�?����=�u��� +�����xk�7/&9�f8��K�Z`���8�!\��۔$i�����ٺi�]�ͯA��J5+��2���~m�I�6�Cϩy�N增�Q��D_�l���쯷�m�ܭ�%c�S�IC7����m��c�fL5/��ۇ�yb\h����$���;=����5:�M�	U�^��wG��������;2y�۹�pb�&����K7�Ѷq���j�/sFz����m�e����C��h9�7&Pl�ل�@��U��P�3�;�$��r�2����:lm��-�,rdt�{�J�w��r��7�_/m��"�������N�~�'ev�{���jV��zv��C��}���ï��z�!G�[����s��,�rC=��w&�=���Yf{A�3�<��L6}��^�̙�[�s1����kN:>�͏�}J�lmQ~<��nWW"�\D�.���g�m
�T����U[�C�8w
$wm�{��|Tz4�$T4b�Ӛ����h�`��X�ý2{4E�S:�qp�#�R�⧟�s��o?]1�7���k��x _e��Iw�ћx��{_^�=�b=��1u���S�ݗf���P�����R��;F�=�#`K�C��h�7E޼qO	��?$r�����$kaע҃���CK}3+_�u���>/^�{xOxļ��{���̦�y�xu'����\�:�ļ}=B��t�����~O��0qq� ��ILK�cW7y�v��\��,����%��w[[^�X�Q��3a���}v������{4�W��+Cu%��u�ӥ�i�Q;�`�Ҟh����b_v��@w��Z�}��7�a �M���.aC�����r
�]b�ޛ{��~��r��R�L̚����d�zn�B�7r�� ӑ��(��I;k(δJ�H�(m���P9	G�Sl�p:�;����:�G"P]%�gXGQ%�N���%Y��t��	8��Y�gu�qahYm�;����,�&��U��i"�.�J��[Y�\��֗
H6��;[Rv��"9�e�A�DQ�A\"!�vwb�jÚklt�9 @]���Y%�fڦݗX��wDYYpqݶ�HIm��qӁ�D�\u�d���Ŷ�;88�#��)˃����(�9��s����+!��ft'DPr6�-4����we�i�\tQ�G)e�tq���[[�����̬�ԝ� ��L>����޵��uy���1�q��6���w��|�ѿ�9	� �{�i�]�Ο���s{�MBp��ϫ���H���m6�{/��Y�^���i��1Z�>f{/��*]���o��#ѯ�3�&��'�h���r�`Uٝ4v�+�e�
�����ņ��։�|������z�m|�A�͹�:��ԏ��v�o��;���n�m��|�w���ѣx�r�r�e��{���/��y��=5t��eA�#�{�ݹ�5�m7_�{{˻�o�J������."/�6R�����i�@6���=U{��]L���ebc����<ٷ;�R�Qp����7h�,�9
M~������[���=����X����L�0�+�O��^���~�w�\���q�fr�\�5���fә뵋�pP��t�\����3��M���m��gLWC�ݩ;��_\����zj���m�cҕm���
�C�5�f�Up8�%!?��[c��s�]�ݹ���jz�X(i���"�?E�t�LV1�G*���d�R��J[�8f��^߽<�q�6�m8���G�Ʌ.����͞���ԏ����\A�=��r������7�6�m|���z���1l�]�noM_��M�t�
���
�ұ�{y9@6��V1$r�/��݊_}�Պ������8{��]|�A��u�l{�w{�;�f��y�����{�:���g����{}l˼��em���a�L�n�����N������%��Q�n�;�rK�Ĭ�u��ݱ���:��]�L�;۴�0�6��^��~}��ކ˃�p�A"����饆E�������5%����Q<��R�Xl�0B
�6��]��͑��1�v����嘳ܺ�oc���xԝ�G�E,a[���<�m�<�qn�S���l�#C�����Yu(��ȫ֛:}/$؏Mۣm��c��ZFKs�\�Ⱥ�����R��3TrW9y��U��u���˲�v�v�"[�|�S����ײ�n�J�Ƅx11��GF,��Ն��2��U���6E�E��u󑷀7C׻���k��u<Ssx"�M������m��m7M��R�Z�S�@�CF&:G*���{�vK��ټ�ub�Z|ƬG�h��Ͷ�����tY��Fg����4>��ʹ~���ɡ�����}�wot���.�Rro���2���O_�q�t�9��|�_���RUD�j�;`�IW���܊_esm��پ�T�|{��!CW-uƲ��ۺ�TwIx��:�Q�h�'�5�n�d�{��|i�5}N���R>����x_����A����r�T�)��S�e����y�=�>�t^W���iOع;��J�Cƿ	�uxH#��|�����{7(�dU�v��7=�Ov�.t.�hn�_z�Rrozjt�ۧ��/\��/���|�i���]��-
���V��������r�Cޛ�K�w��m����.Q�|O3��y�����|�{�M�C�zjG�_������K:�y��@I����7A�����\�x]�A����}0�ȱ'&����Jm�ۺ�s�o���U�$s�㒇[�%�t�Ǥ��'k'/npkzեjͪ�*��*��}3W�>_7_6�xSG*�D��nK��ON#vΫ�Ofo`n�k�ۃf�+A�o��K��m|�>����MH�_��\M������o����m�������F�k�'�)��[�[�՞]��-�wہ\SŚ��_��;�V/3�|u�i#m=w8�7��ՠ�z��xy�Xтb�����fݗ3L���쩊����Wão���kR<�#fD#���Lt�뼥!雒��������Xk�z1%��6�tcl�o��s�N���bw�=5#��@k�7C�ڥW�ُ'�pw�u�D�N����۝�^a���NJZ]��ue���e9�K����x���u��&��S97�^\���ߏ���C����@7_ٯ����s��<�bI���Ry�._�Ͷ��� �Һ�$_7A��o�v��8��&��z��u���;�1�}~k\M���o<Vi�Lnw��[�6r�����u�Aq�YNM�F���!�&���a ���&l��y�L�����R��"j����ȷ��P��u#0+[*^�1ɕ�z�A�<��̠�b�O
���_k��|�M��o�М�˨�*�=��<�K���esh6���{#�Z��B�U�R����#-�M��nI��w��1�֭��sT��oR{�����ͼq����>�Sҥ�\G�f�^��"��a�ke�@�� G\߽o�.��D��O$<|YDt���f����Aq�^��G�	�� ��m�l^Pt�@�W�־e����-���̱x��./'WV��o�7�@.nł�(��۰,w���F�:7@�"��29��|`���̻���oW�5����簮;�"<w����T-�D6аYe E��%-U�V�>��\./S�2!�(��D���!�#�m�����2��Xo�뫈߮���D�Z�}��)��`�hM�P������J�	��;����H޶��շ�8�MQʯx����H��T��ȎԱ��9�c�)��;&�;)؎�!q�kv���iV630�k��X���a}�{Xm�ɇ,y �Y���T�5� �`�\��&��l؈FY���٪�ha��X����ԦSl\o`+�C��z!��*Q�6� �� Ft��QH���9K���61��g��6��v�<zXÁ6m�m���<r�5����f8i��~���`���q�"�;�	Ig�>my
�؃Aۧ�9������(Z�u�㟹Y�~n�A-���~2k�r��^o�7F�}����Z3���=m�,�Ns�i���{ؓ�kYe���ܱP�>�S�0N�Sr��������?7G/�[�+�q���K�@��6�X,��n�m���쮲�L�ê���o����L}`�,��m࿋�B-����r�f�}��2<���b���Fg�S�����	�P@�꛾\a���.��NGr���̲��6�|穭�yM��W�N>ۓ��N+��z�C�B �K�	m���������lc��+t-���W3�=�ۮuR�-л=n	))�#	M�Ԡ6~����_��>������ ��߱����x8����{�5�t�GmF�b�.���/�%���N���{�{^�H1Q1�W�{��	vjʍ�����J|^����`���$U}�|b��}7s=|� @/.'!�����`�a�>�j����=�ꦼ^o�6G }���`���z��'���e�������g9e�n��C�Fz����ݞ�����(��!jE뒸�����׈%���Z�P��:�<M��:��C�q。�~��goM������p��/{s7��������2���\yʸ�y�^����U(R�bƏhv:m��5��} �A�P���g  ����0ccg�/��댅�f�I�F�������g�F�`�D�!K���ɝ�,������ieg�H�6�_��!�<��!���^�+�J�Y�d���s����d/�t��Ր�U�t:~ù�/uWXݝ�s���?7_j�n����[=��G�q��ˢ�ۨ��,t��r��"�K�y� �鐁n���^(�>xJ��o{�;Ϯ�z�Y�p����Gaך"<M�'����FK�ڷq����e��������^�.m�����P���ӊ��y��x�P e�"F���? ����c]fUG;�YG� � ��.� :d'��=�D�H�rW@7澵���{�:u\?'Y� �VC-@�[�n��Yf����j���Z � z��;u�ԭ���G�w�(҂!�_̲%>��=�^�~�񭌪��ps�:��h�)зnXa�ɓs�[��'��Ѻ.�TjS���u� [���լbx8��t׋��������`�� �2X��(�@6�X?Y_���~Kw�Vx��B6E��q=ɳ�DA�(9r��� �m�4�n���F��ߐ���!�@�΂���8Ct
�y
�_���<����o5�Qlܧ���B��qvˉ�r�2�,s*�'ח�W��Z��6�B��@��ݤc�)5:���#���_��7
�`���&����S?v���G�zh)�S�=�O�vǽT��H=���D�y�oW�͢.��V���K,�e�xn��{7�o<%RC�g�~�ݯ�����7pK���&�K��|$�#��w��B�З+�J���H�0�wi��K;��������&��p���mv��'�x���Ӟ7!|���.V���w("3�#�J�����n���r�g��7���/!��i�g��w ����i�E�pb���x+ݛ`����x���zTN�z��o} ��W��}"�N�Iv���sD8�&~[�� �#kH��6C�����^S����U'6��^RW	�R��T!�Dwi4����R�a�}~X�7G��;�/�����3�,~/�@�|x�EU���{}:��K�Ks*�G2�"ei�W�mf=yٜM�_��K�4zmS�����Ř ���8E|A̳�!!I��!!I����$��!!ID��	'��$��HH@��HH@��!!I��BB����	'�$��HH@�x���$�BB�a!!I�䄄	'��$��HH@��!!I�$��	'�$$ I0���$�ي
�2�ɣ��`!9������9�>���`   �   P      �              ( �    T)Tc�*�@ ���P$
U
R� T�U)B���
��(� *B�EQB� *�(�����
7ϑ$AUP!D��EE
D�U�EJ���ED�AJ�$�EJUD�T�RHH�D��*��RB�� 4 �"���*�  ����J�V�t$���0 cQ�P3R n�X���@s����
 f�JP R��  }��ﻠ!.`h���� sdAB���� ��z ��� ��F@��a҂���� ��A%>   w�U@R��$I
�E	U< �������aq�N�p�s N���y��3`�B��=� ��U*������)!JJ�Q� �8�@��� �É!�*wA>���	
���A͔z�R�K�\�^�����:
3 ���PPU�^fB����hR�P��U|  "�D��UJB����
���z �(� q��� �(��Y�PPK�<R�� ��m*��ܔI�%*��U$n�HwUS�t�U��"�(�
>   l=��\����T*���ۢJ���V�r �wED�QUSq*����ͨ�Wv�TlU P P� �OUa��IJ�")D�*R���QU݃����
��(�YU�)TwUS��)n�
��,�
�`䥎��� �4P 
�
� =v�*H�Z�T7���%H� �sU2��(�p��t�T�Ί�Ws��d��t �P(PL� JG���E �R���"�^껱ԅ۩J�b�V#@�c��Y���)J;�}b�V��ץU+�����F��U�8uJQ��Q@J�P
���( z��gAEU��JwU�êwX�T��Ur�mJ�z�n�R���!R�T�Wuܧ��y����2RU	� ��5O�4JR�  ��U)�R� 4 4�*�	U=C ��RUSM�   $�E<�T�~�z�����������O���BI.Hp�m�J~��4��s�ׇj�G]����$�֩�����$� @$$?����$�i!!I�$��	" ���������w�����[�w3n�5��jkr�����*������l�Ӷ���y����e<�E�4[�N+N�`j�:r�����ô��me]īokv�0^]=����)�m�y��f���)����"nk7���ܛB���0n�I�M�����h���x&R�kZDk�jF��yY72�3�-;�1�z�m}6·pa���5��*%y���1	��ىf+�E�873m
�F�5Z�Q-۱pVP��O �v�N{Vo���V'DVj�n���"���BX����6n't��ʺ�J��l�Y��t���˥���3lP�K6�V��F	��Ƣu�n��؝」��CF)�(+5E
��w5V-h�K(H�]	*Ά��j�+��ݓj�$�_1n�RT�W�ū5U��,sjA�����	�3M���-�V���u`Õcx��d=���v��gF<�����w�q]SM�h��T%�T��a�*V�o%��;��*u�Z9x�!A����ս�Z�l{m�or�5��]dKs6�#���*ɵ6�����F�3)^�-�qlT��ʬ�p��Ļى^���WWa�hN�Q��v�[1���k�E�����[�˦4�7-H	ZsFY���Ê��V7[-�Ԇ�l����/q��֙%M�Ke�Ǧ�ռ1���R����Q�VkV����P��AUc0W��Ø���wM�}TQ�@՗B�oA����V��%M��T1�cR����ő�0;*��}U[VqѸ�Ch�dIc%,"��C�E4�#-U^	��Gi�b�����*������Amhϲ���]���6�Cd�%��EU��!B�Y5�n�L�T��W��W)���<n�^f�$��d���T����p���qR����b|�	�b�����w�e�Ʉ���v��K�1��R�k�����ǧ7(�aV��9��L�[����4�͗m��hRV/T2[xh���M�_Wl\otV��63k&f8��i�{�UA��e��ԭ�5���ã~*�/o��kLc7ME��e ��3,���ƁڔF�٠������5,x��K/]%SYi��3%P�;,f����0�J�Ī�6��QS4m�X�rŕ-�/m��R�J�����n��Z�ۚ���Y��Yt�V%&VfQ�U���z��ض
{[m	�湡
�Q�(̧0R�V3�L��SZ(���z���A����r�*�N�<�Ď���;C*�M��v��gM	*�]����P�F���S[X�8�L�S.jkn��t	C4K��f,#+r4ݖ�����M�[��h��Ǚ�ʌ����	�(�5)a͎����ǒ����J��T�P�e��-��Vvm���f���sa���J��)���n[����ed
A��2P+4�f�b\٢d���c��޶�*�YtN�6�Y4�f}�CUw7(Q"�S�b�܄]����9�'y�����Dv�`��\gv�Yyp��gM�7�h��e�yu1��l�h�Vj��[
=�v:ܛ�E��a�N������7����m�+�d��H�¡UR�P���(e�&�T���Gt%�I�]ԁ�wv`�stO���ãc�]�[�N٣+k]U��~�P���[��B�3N\7�laͪz�j�[Z#uk4^��DE��ж�ZQ!��׋~���o;�iYV�\��!nh���5W"�q`*��u�؉Q�v��Q�X`r��k?��M��[�i�4�c]P:)��bM���'Ƶ�(V��F�I��2ș�1�A;Vi4D5y�Y�Ǣ��R\��.�b�1�tЪױ��z.fn؆�Έ�ú�r�w=��h��Nb{��
5Z�M[tuMZr]��?���v��]g�Yp˛�H(��e\�2�n8�dZٔ7P5��rcX.¸���*o�Qi�UXQ��KrU���V�<4Bsi͏7,���&�dÓ-��{{��u���l�[(�
��܃,��6����/S���W�wnħV��v�� �&B��ϩRcY���֖�:�uKs���v��+U5�.����FIf��5��v�.�v�
{����Tt�H̗x��mM*�RtJ�f���:�J�P7�-UZsn�;;��N�&��GX�6��	iY��!~5���ōXW�R��3�E��E*xi"�Y�6�o㘥����
��9�+Ȫ�٦�%t��o^����ز�I����f�nB���2ݗAYD�+(ޤ��4S\�+Z��+�Ӽ�J�ٷL乘	��km3��e�&��V2Ƹn�n	��ł�D��*n%/.��9{Yck2�������N^�x1ll:�vV;cB�eo�Μ@P­9f���n5m�����f'jn<���W�k
˒ܕ�2wZ��cvM�V�[�pf�
�1p6����܇(UF��F��t~Q�
�+�ĝ˽5F��MGy�3l$�u�f�/e�w��C��m�W��N�;!��Q��7H��V^�17r�
�;�E��o1i�3#�shnܧٳ1��s��*�����ʩs(�2.�3�F�K��OU���O%e��XţT�_�cҤ����7w{z˱vN
ɲiwd�2�Vl$�Z �v�i;Z���e�N�,HKwR֪z��"3ou#f�a���;v�eXI`��Lu�K�]M_Uj��[Qp��n�l3D�Q��X�eCQ�b�{YI<�_Q������RP( �'Y	�U{���F��;Q�
\�v�`�דR��������>�9j�٫v�s��n���V(��4�k�v锶�Ix�$�C�k7fc͖��g6�62;�;=���xB�5죔CtZX�+jh8�r�mDK�6��Z:���8^�p2��w�ʛoP�v�3%�'�f�Q�V�U|�e��o[�y�t�̫��a�M�#���.�PmU	Oj�9�!U���[�/1,m��C����c�{sVk���*�� �Y�T���T���Ũ����ܻ����e��<�Xh� �	��L�z�wM��w����7so2&��$|iUM)�3j�U�+7oV��U��KP�f֘h3@�������w��1�������]ґ�����UiQ�T�����v�Ix���*}Su9v�a�h[v�ʺB��4�[���j0˙��F���^g�#cLa��iaܬآw!��WM^���f�֫l�"W�F��k���^Ջ��X5f��+�if�������Keaf����if踑9Yn��{��w�ں�����BX�0���.�<8��[)�4gIS1]���G^ӳjbqn੺p���a@�
j��m���Z�S%�,(T��`�,��W���j����T���4�n��v���֢U�V,�̐��s$��D�k�Gn�i��tD�y�~��$��X_U$��8��F�N��y��8�7x+]V�h �)UH%��X��v�o�aV�+[;u#�ۨ�p!S6iɸniz4����zQX�&�2Y�U�^[�9f�7"Ow&;�eʑ����j:�6t��7vmU�@��m���WCo2S�Z΍{�e�[%Ld�LeT�lv�%f5cjV���@�0@Zz\�|�0�j�a:�kY��d]�h�Rƥ�\m�Ź��y���͔�3Py��Ta��pl�`$m@��U]����u��4]ѻ?\y�Lj;��콍�ܦ��/�m�R^�T�-�
������t]��x�XE�[Z�2ȵm-Z&�I�p��ܨ�e��YRV2oH?i�*IDŕN�w����\�/�&��zfn-D(�5Yf�UkZwv�I{Ba�M^����u�]�ُ,噐+�x7E`�D13,)YNÊ�+j����%���"��ATor�,���w��!6!�6FӥxT� �؊,�̻�.��+t��63>�*�{�"�A��n���}��L�T/V�3FU������mf�F�Ԛ��&��gn�f:�*������˚�1Sv�;��Q�	0��n��.�ZZ�tR��Ow`kt�w� P��h�r���L*�c�0m�aݼ�RT��#	��M���⛖f肮�	�n�j�r�@�3�e��M�7yf#�L9Y��*�/E\�t��nX���_��wF"u��{��B�
��ɒ�GB"ȇf�e�sX�@�*�a��O�r�[a4ε����B�UY�����C.�5fa9T��չW]d��X�[6է��Y�j�&2������E2�$����<pV�Z�������I�wkw�vfT��Y�#>�xr木V���eS��m%zM�ޝ�Wz����V�F�xB��q��
�ة��6c;����3W�@�%'�b���Am<F�ꝙ MY�G�!�x�:�&�2c��n}6bwm�g(u���$��˟[��u�՜*�^��CM�EJ-�on���$��(�uWJۥ�)��Z�����^,wr������FQ���pҭL������A�J����kF�S���56���N��EP�67n�cE��Ӑ۵X���tv��mh�ʉ��-|l��ʸ��y���=���{���ϫ�����B,t.�سWT4Q��h��UJ�[��^��մGQ�JkAK�ڼN\��
�`7���5�Z�mnk~pi%Y�(¯/5Y�Ii"Ϋ��r+X��6�hz�VcQvk۩ut�U"�x�EƳb���t&7L����7���6�ѽB�IC`ޝ�Z������h-�X����A�!��+Z:���cW�%�2�%.�/l�L������֌G��ꍇGlR8ȉa�Ƶ�"�I�Nn^jIl����wWD���(7*�fV��fʶ���,�/U'Ygm2�F�D�_ږ�"E��7�~Wyn��W���n�f,+u�W�*��,c-8�޺"�]]L�]���1�92���e�chT�pLZ�ݙ��h3i�.�Xcaܼ'#��f�X鑁��0eL(��e���r=j�6�pMʹ��ۣ��dy�5���7�A%�)fY{PGU��ȶ����×v�f��Q���[���������-hg7.k[7uޚ.�p����b�[ۼ���۪FV�h��,D��F�W�
���\�,�ko����U	v$� o��d���*)-�cQn}�X(a��^x,���2��$Z����*�u���U*ۆU�b�鷌�n����>�z0̛�u6��26i��&�[��-���&w[��#��qe'�Xi�e�FU�VP�t�a�N捍�{6�k�cu�H�`��(L��.3I4eee���X�����*10�̪��fh�6�k�i!�k�nd�w��M��MT��ڽL����:�o�mܥ��v�I��.��	Ya�Y�߲�0�>��
����e���)��Ÿe1XA���m�$��V���He�iֿ���z���!KW�iK#W����]+��J{J��C�V�)�4m�̬�o*'X�H2��UB�rPL	o<���ƈβ�f+�a�enܢ����մ-A���&+h�2�e�։�n�&�E�_5�UY/+&��`V��,Pk,b�,���ݬB0�Y`�ũ'��OFՑ:u���5���Zb�ͳD.�
�uY��i� ��j�:�������R��4�Am!q�EP��,��� �;g�6��Y,�v+�j��#��ũ6���ͫ��T�V^e^��鼛�8)cL%�"r������7+lZ��B�l+
V�	��Wk1eݚ���3n� �$��%GT�S���QIX/!�+u�e��h�n9�5��	�W����+.]e��\7ėdEnMǁn[@��CZH9�yP2b��c�w�-h��.VUiÓ冪�V�ƛ#V$v����a$�S�ݽ*�v��Vd!
�+�U[9�ucjЖ���X����*Z��E��wX-�yZIX,��uC�j�]�	7V��(��a鯍܊YUn(�V�X���o.���%<uT���nfdh!��0�M��W9���(B�uK��$�̵�e����u�S8��ӮlC ߶;����H.m�B9����ͨ+(E���'-Æ��͵T.��,�ϳ,�f�엷"	T���e������dIi��V��GtFe���0e\�oD�ue�ЏD��U�]E8�ݛ�4n=ܷf"�Rf�Hf|L5w�#�%��.�7���,V�V��5U��#	�R����	yBnӭC^=Z�[R��l%y�ԭĔ���'��i�����[���bz��ybfU�Xu˧� ��6��xt�oHFs[����w�R��*C���n�i�0�t�Z��U��b�Tw2��`ڸ�Ө����u���*,��˪�ClY���!r%P{X�̽�fm�J���-=y���J'c���m���aĮ�^��,��l��ԱS���fL�*�ˡQm蒍�6ι)Up$���U��W�6�k)n<��S�Tq�vI���1^�#ޡz2V����L˺t��)nZ$���E�F]��Ю`5w�Qa�×y�<&��W�2b��U��5r�7cUm��ZW/*���V$k%�n�x�i����
RB��q���j���9$V��Ťɴ���]b��'^j#sNv��@��Š�����Z�b�
֯��:��K6���Q�2��6\WR��X�B��dۨ�WL��Z����D��j��u���j��֕kzC�5���Ǚ��U��Zvv�oJ�e�7�����9�=+Ukˡrও�JF�4��5�=��У�+f�v�u�ẻ�g��{vN	b�&��,Zڤ�$@�^nf�Eu���Fۉެ&h�H���*��ջ&f�EY"�-Xu���֚�qM��ń� ���:h5d�x�٩�F�~T�7;�(X�������l�-��ۡ���8U�k׻�h#u�W�m ���76�K�6Z�/r�+%*��sO�Joi����k��ouw_؁:� ��!	 ,$P� �H,	I$! ,�� AI$R@���I$�!�d�d$�� ���@��uQ�\T]�GW�W]�H��BYAa$���]�U�wuGUGwuED�R ,! � E� ,P��@ )	E$I E! ,$��$Y �$�XI"��������ꮊ���*���2@RH��Y , H,����� �I"�HE�P�躺����������$�
�X@Y	$!�U�uwuRUGDuu)! �,� ���H@Y B(
@����� @$$?�BB��5��^G�~�s������Y�fͺ6�v�jCθi�z)Ȝwݽ�V�nY7��7���w�s.](Q�+%���A����l���e�!f���ʈ(Ȳ�Qʽ�y�rT���e����&�۩��2�Rm��ҹ���im�Vl�Ⱥ+��vy�Z$�Fk}�������N8�ѓ��'�T�uI&mmu,.��w��"��p_Ye.(뚲��ŏ3�icp���嫌r%��
\M�C�ߨG6���v��v�-�vվl��yu.�<1�d{1e�#�*�A��p�\֫��z�UH�f_?��16!��c��o�%�w���;c��e3��B٫F����5�$�կ5�[� $h�����T�����R�� ;9H�:�YJ�iu�.�M0���l36�́�{̫U��-[b|���wYݪ[�ʍ�̭{;6#�>��X��b�Wܮ"�FQv�H�Wpcl�h�u'tܡ����C,UP�&���}m��2��Ġ�����1������`�\%nJ�X�]�q��)Df��&/-X;�t��T��J4F ����;���x�LFX�U�Cl�<�Wj�L���*c���U�q���c;�璲�Ln��%��5�u������E�ЏN���:fwe�hU��}a�ұk�:�DY�ڄJ���7��牽�!� ո����qT��m�|�.l˧�F�	]Ү��2էy�9VLA���Ԯ���\�Wt�tٷ>�;ʎ
��!}�`J�����LJ�x��+v�{wU�&{���R�2蜶�X�o��v��]^Cp7kI��dwػ���^.�6��R���L㸛����fۻF#(lCfS'p-�����z�܆�j�V"���u(�WX}4l*�`}�>��zq�y�U���J��N���7:R���l�ڌ�k)n[SZ�=��.0&��\��{Z���΁�[���i�g���J�U�)8�F��d�;:Mꤳa���yM��[��a�c7{�.֯,Pk�-��B��Vh�{.���<�ld7rLܗ���,�#өv*�}x�V^1��M7Ӷnv�)�}��M�������U�I9f��ى��g��Ft�n�L/ZI��om�w3��ۼ��]�qceZn^FD�F��r��,�u�ͼ��׮��uu���·e�٪�5�v�g;��f�Rw5P�$t:6�3�
]��-@ʬZ��v�Ҿ��¨�yrͧ��֑��h�)epshշ�%�)�)��]*��<��p+�,ɝ|y��W)���R\~ѥ��ͻU|Ă�R����oc�N}��l���*��Rv�Rm���hk��"�b�<]����]�8��S:�5X1<�|��̶"�.�b���"���2��u�L��ʜ���Wv]�\�Y]bKvIW����g�1<���Lf򞗶��M0UU��^�b��0�6v7��_7u�Չ�2��oi�r�]�J������G�YvQJ�:w��w$��՝x��#C���(�6�����ƍ3yxγ-�;��5���z���E����.��.a��v_��*�ۤm�.s��6�+W�a�H��컱a�l�e�5�,v��1c�W��NCBKo5˭�-|�9N��'6rs��$�'7�u9؅rh4�����O*t4՛i��;�f���%�u��Wv�z�,dM���
N�'IʔI�Y�̽V2��8d��f��Y��*+�r��Y��n��������e�s�R�4��й�4�v�ڠL۹V��J�oV�|��J�yKmi�p��u��͍$%r�q`�Q�n&*S���*':�
��FW}�ҝ��+��l�D[��/z��zk7��԰]�D���C���'�m	���걃 �ù-{V
�ޖ�K�K��̶:�;�ۦ׊R6���E;a�2�-�U�y��2�	�'��IwZ�g��v�e�vS���U�fŽe����ʖ�5Qr������Ӊ�5u4л2 ԫ�C�Uv�����2�-H,u�J���G7UC����Ju��X��NJ6�:ñ�h������]]��WY'��\�1���,�ֲ��o�74.�B�*�"�[ܤ�-Ae$2���[�:Iv��k��7����O;P�:m঳�R��ٽMfN�Wv9+�d�*	I/�f)�0Y���
�G<2�ǚ���b�J�xJ�c;��g�Y=��j��V<�*mi�A�C��RS%���{����)�Z���RY�[=��-ݪ\3Z�pe
B�UsL�ˬW���cv�K�&�Â)��˟]+u��cb�I��%�p�r����Vd-��uQ֞UX����w[Q�(�'R6ky��>�~I�
�o)�|���1��/Q��.Nk��9N��̩���9�8��"��P̻9��L]B�&���H�p��MM�s��-�=dQ��O\l��7��l����xNu��iVZ�(Y�ӥ�_t�.0�K��p�(mÖ����ue��*վ���l�+��U�E1+����w����I1�f�a"�1jo22�ŴU��7��k]Ɠ7:vfu&n�lQ��X��^�Zӊa��N�P��!f�~�!�����	�U�;�Jo1�u���E��N�Y��v�������gimaݥ�1RXkk�p��&�����1���)��Ǣ��YwA��f^��i��y�&�ݛ}W3r�uu[T�nm*�\�T��!�ޙE�;���3��s�{q���л�r�3�݊�j[ћM�%��2���J�5D�h�c7�Y���}ɷҷ��DU	u]��3��6A�f��!��ʻY�,؅�ٷ��gۛ¥��,Mљ[	�1�;[]?�ؓNdb�
7���^E3�}	e�ym�f����m�U�Lfo��}�}�G�w��_n��#qޑ��W*�
��fLm�Q��z��K�J�b5e*ӱ����m�y0��fo(9V��<��4X�I�T��T�`Pf�}X�Ի�$i9C�f�7�	���e?lX�x�iGsg\�����\lQ�Wͺ˩Y2��+�Ul��e�aT�v,�!�5$���[��9bqE�E8��9�����&.r.��Q��ʠMkqps�ToCR'[�ţ3��KM:�d��M��]U��$�S�qX�4�L}pMd���Y�̾����q��Y�nf}O3�j�g"s�h�Fs�ݕ�(avN'/V��U{TpX�Wr��w[�G����[E46����j��_�:sp���mȃ�=�B�i^Dw,j��UlȬbֺ̳~�*�/Q��)ɡw8U��^<�y�**�NXj[p�ښ�Y�G/hGd��ry�x�Kh�i��U���t��u�������{�H�`�Gt\�Y�u1v��:�S÷���)m��ָ�����rov�:m�57�u��1B����AUP��/�RZ����x_(������Y���s�#DJ�'6�W"1U��UݞK0�R�jNR��5r����fc$ô���f)Y�PV�ŗ*��N-
�Z6+;z�a�7ԻȢn�3[Ѷ���Y�{^���.�,�XB2��u��6}���"�y��r���M��P�Q�kc���J�9Y�9�/[�}�=�Ղ\��R��Õ��g�ssU�XM�u�B��ۙ�>���ɹ�M�cjdn�y%-�}}A��V�oa�`e�t#X[-���Y1�i+ƝL��,�/ui�m��l�v�g��'��!�R����ԩ����r�ؓ[���ɗ��ve>N�i\�B��n�WH�����ݝ��*�fj���sx����F��u)�m��E��f���	�Y�Z���չ����4X�R��*��;3A�J�ɲ�EA�v���[�>DN�)�T��[w4o4���j��ު�ٺMTM'؁wd�*��7�LJ�k*պ�N��6r�o���Mn��J�-�&*���a�;�����}F�J��X�NA��g���,Gu��\�о�,iN��y�[/*��jf��Vu�Y��fNpf�fT�[b��\2'��|1[�����f)*�9�i���ba�	�����Oj�nU(�:�k5�z�1L!yseG󗛷պa����,�9�.���sE��}���E�2%�՘:�L���]Nco�S�fj0��5n�;�n��N�VV��M�o9�e�	��;iNʻwh���e�Y0�\���i�C�oRB㼅�sk����}��P���4���J^�L6�臄X�u�<�6j�&��EA�}S��TSc������t<��ڽ���}�[r��s�:x��ݭ�
+w�@Y�;<���}�Ayx���n���ٷ6�1u�:�T��uuP�!wuz�i����Vt�i�D$��^Y�{FW���^�1��fim���RH,ie-�L/���˶�)[���	��)��N_t���5d)�WL9�Yb�_V��%��($r�y�q���6U�n|iS��+K�n��_(.����E�����uԡ�3��7\��qC.�(�m;ȫؕ��M �F��Ռ���y����3���a�mK₾�7���lQr�ȂH�S�gd���>��i��V��uTjQ8'"	<�X��Ta'K炘5���j�����;�CNR��k5{M_V�4rWa�o�-aW\�5U��#)y�s�K���<��9Qv�q۠��
+L0��n��ʚ/n.��yaT�Qt[�#J�G!8��u�Uc��:��0��:c7fgN�w(q}ё�MFLN	���3-�	�U[v�ֺ�cw�<\f$��U;����꘬��V���;췶Tռ���<e1��F&SȱkM�ڌ���MI)�^:�"�_9�(v:gWo�8#�m��T��,�V����u�#N9��c���R={���k��g��vj��v����
�4VX�
iؤ�ܝ�^�1}t9ۛv���v9�U�j�)ݹT�dnۨ�x��^c��QO\z�$n�H.���+V��5��h��Vs�Z�{ٴ�9��q�:e�]�K���ƻ��Gk��n��j�n�����&+]"B�ԋ)����ڬ��i^�͓��Au]'6)j������ܾ�;���<V�%�7��T�.2���[��z\���-��i8�w_���ȫ�˖���V]A�+:��Z"���Ǯr�2i)���9p�k�8��dn(�`����U�y[6:��䝚�����N��]>!n��M�n�U�n�uU�#����j�9�$A�pi٦��ۄ@`KTx�j������A<,m�tJ�x��Tm��IAab� tU)�$(W��C�fjǏr�֏n�xU�vEs����E���j���˫�|.u�q_N��ۢ�d![w�3V��9����ЧL���bA��Et9�'e�W{��e���p��`˔��-���Y5��p����Q�0t�iǽG�z�L���H��Q�����]:����Mm�̋����Ep�%|����F�ʘ!���]p3%ޜ:��.��$�8�,��͇z�ق�E�5��ib�y@߰UM�
/#۴��7QdY��@�:��������yT��Uf�˥y~��q.�x��U�b��r�]n5�e�8�p1ܽKd��9G�N��^Y�{VLT�e�e�d?A�[6�^Y��I'خWY��ŜW_A��k�5�+�k/��gd,#kC[ԫ���%P!hŹ�>vm������;.Y}�]�eb����ݖQ���a�g��Bk��H��ޮ�8��[�bGd��u�Y$z�뛦���b�u�}o'sG�j���ʸu�r���{%��j�L�������#!��n��-�Yy#��m�\������ۻ�j���y;c��(��V�ʎ�Ô��Ի�$�^jrf��Vf�|�U�����;J=�a+W�X���{b��}�/�S�����A���n���⡩Y��ڍ�.����U� �e�s9c{+v�)������7O1��A۽�b�Z�.Ud[�򰄃h����7t>Oc�oAr�ٸu��5�Ϯ��({C[�(PSycH+,�7Iz��.g�H�H�cJ�gfk���}PmI}]ݛb�֧�̷���� �a��3)��F�S��ɓ>v�p�{oZ������雽���S�4[�Z�]�TE�aI� �E��x�Ӎu�w�EIdf�oGo�������ԫ9w�Ҧ7m��<�ʲ1���3!ޫ�����v�Z_9(*�u�)�7�f��78��H�
N+f��A��f)w����UA�t���M��ǩ����V`9�ռה�yu�e���.*/b���B�-tZSB"N�DTSR���7��F��r*Ă�»r��o	���<������ͥ�ْ|��X�,��W�[0N-Vf���vѷ������6�y�����+�+��sW�p���)�-�Ĕڭ�kb�Uy�P��K�1oW�4Gv��,R��F��MJoƥ�kzn\��1ZWN�Cǅ��5��Ka�!$`c�m�Z�*����ҥ�����T��GV�9�ü�j���uK�诊�}�f�;�V���N�^^�h)[�L����1��t��An��egG�=7r�Khp��[�le��Yי4T���ݱcU�*K1]��Gej�Rڗ�V�{muk]���{l��;�M��9zjs��:4G�9��[���;��}Ȩ0R�y+��B�Pre��=v�w9X�n�-:/wX�~�*�f��*ެ�����B��V��M�ݫ�R�$͋�[�8(:T��a².��]7qVw���SwUD�X����V��L_�M�.�xيŅXم�ocn�6�h�rKwb}�����X� ���\�󷪊���[�\�H	���M�.�M�Uv4ӗ�%�E��բ�]�Y3t-I��E�h��9���wU).�2�2�.볳��,�/�R��1�j3����}��۾wO����;�Y�z\�U���&�M@bS��Û���i��j�W��r��wf]C�gqP���6��v��&L*H4el�SM
I��͍Ɨtކ������%Z�U�u�t�rmwTu��I	L��+�*�j�֓Z��� �oR�]Ь;7:��A͚6�0��R±\٬t]�mN �f!�+XO�E<<)�����<�8+�����kɕ�6�c�ңZkb�tl��\Ҵα�C6�L�����6M b�T[�u<�Eo))%�B�sX��UD��e�V����\	�,��`\��ʮs-�,���p֖��t
��֫5]/m�U%��f�2X�X�.f	G�fP@���R-�/Xa\$GqcH���1�8r0�(�T�8����6�ɘ�m��Ef�.,���Z&�[��(d����s�!(�����2��#-�F%�4�\�4N�ґ�J���4#��W"�4�Ky��pKsT��V3��1�e� ��.�&��vY����]H�2k�;q�C������x����ɶ�M��M��n)F�liJ�L�A�Z�ɣ��n
3f��6�`��ƫ.�JK�#y��Ш)Bˮ��q�X�]љns�`h&6"KifcV�X��U�r��ڥ��1+�lG#{CW��y�]/���&���L�\���h�7k0�V��H,m	C�ճ�0z��Ҩ0�٭�\,D��j�s���64tt�ȹ��whq��3l�j���Uz�`.�Ͷ�-ז�6�Q6u
#��(��-
J4Fd�Me̮�+EŻ9���e��a��&c�	�i��de�5���l�cP��jĚ�3^���{Q;E��+����NĆi�Q�c��:�ғh�W�AAaBqX�C6��m��"�0n՗�Sl/f����Mn�jƍa��$�#�T��(;K��[��h�������iR��o3���u(V� ),�fNuU�`M���ڔ��7h����)c�!CB���1D�j��vЌҔݘ]RU4�̰�6�e���A�n���2ѫ-q��6���q/f�LuH7�r�W�[ 9�a���2�':�p�I�X�.���4m����^���	1����%Zj��Yf�:ٸ�B$��0F���9�:=Ի�CF�f\���a� +��kڬf�]�i[��"���(飪�4��h�V �nV̖dnث���BY��2����n�0�[5�`%e.ҩc,�$sk���,���c�2��ǜQ�8�:8����g]{d�X�a�����N�t�c\�l¦�ݱlԁa�e%��l.n�@\0�i�*��lB6��u��6���h�� u�9�2Y�L��2�\�K�s����;p�8ڹ��!(�=@ɴD�\��B�3��\��JЦ�mp����kQ,��U���$����D@��X���lv��f]e$�,GhP�KX�k�[M6p�3������M��aJ��eV�թ�.+i�a5�R�P�͋Z�!0��n�ɘ�GX�$��hKZ�3��/``Jv���`kv�r]\�\�u�3R�أ�&�0��n��V����L�0��T�f��-�A�«)1u��L�4˹V�Sf�H�E&-fa�LVԸ�[����!T����CCZ�R���$��Վ8�k��u\j������-ʲ��Ku�]v�.A�Z�J�6��)Kŷ:�VRCJ����-m��݆���%]��IV�����M6�(h,�8R:��)*�e�l�P]�f��cg'X�%tmJ37[�KlVac]t�����B�M��ϫ/�u�
L���ٰ���`��;�o�8��J����M��v�����KHL�0�WZJ��.��l��4��4"ke�Һ[`	.�,�-��SVXm�ca�3�GP����[ �������3�R����ծ�,k(R��m��+�a�t[u��mMVZ8q��G:ؗ�R�mF�1�"le#�[�A-(��˰��ڢ�ٲ�ɜu6 uF9bGa�׭{k="Ժ��܍�J��D
�׵�X8M��_��@4-IF<Z�Ԯ�a%��M��M��8���ffX��G:Y7F�)u��J�@ԕr[�9k�w�fy<. ���Vl6�v��/;d���FVj�Z��]v���gn��VD�r��h��R��%KZ[.t��j�f�J��i���sD�/ڍ�E몹	K��Z�1.qQհƉ�ٶl��r���1u�t�).�\�p��L�Hl19��k���	�ځ�Ҳ�em��V��!+��͖�r�7\F�$m�\V��cci�1��]��C9(mu��X&�,�v�h����#�6ic��3M3S�]vez���V�.�rElУ�a�Be%�n�Չma��Yy���[V2�J�+�^pgJњ��噪%H[��	el��Z(�rV�����!�mƱ�2hf�Yl+n[�61�Y����Z%�@���@��Z�׊X�.e��g�	�קm���b1�5%�HK0sbZ���(5f]���l����1@��M��٥�s���R�.�$�Yts���u�3`���k+Ʊ����c1�KB�+�Ysi��M��ڑe�9΃J�)��I�ל�
�)�����%��R���݅@���s�(۠�H�5��V�ssH�K�������IYG%s鑲%2^�t�4��Yp�0��5%�Kή5�ST����U)	�fupJ7�1Lї`����#�%�6b�gRDQ9Y���l�9I��1�u�L��Z�LR!�SV��)FmYd��ͣ��:-�������4�[{Em�iA#-$0�E&@�f���%ҥ�6\!�.L� ���n� IlM�����W$$!�ڻ6������Z����hڻkU֘����JB�����5�e�in�$f9%b8�f:`2fݳIle�al���b
RF�KQ�Wؚ��*���	��F��i��s�0q�#�@��,n��<Ͱ
���f'7ZM�$�P�."m/9���c�^&���B�y�%+��R��6.�r����,vk�s�[4P�jWK��Kc&,s��� �6M��C5{s���
2�7Z�2�Eɝ�qo]�̑f%1Gd$�ͬ�k�p��&�E)I���j8�쫅k�a�`�MM�K,�L�-��L�l��I���Me��^�,���DMa1H��%Y��Z���e���V�]J@�hJ�R]�`�/;fE�f�֠U��Ii�J6��iZK1�,D���,��cR�H*:ª��mQ�;M��m���/]����ڷw��YC�%b��044+����Ƶ�&1BhR���h7� ��3-���܌%���I��p�7kz�C�a&nі�ˌ�`�Jhɥq�X�ܖ�;9	c�1Y�L�a-B�!u����um&JEr����[T�nб��U����Pm�E[M��ۈDذ(Q
U�1�-o��P����DXPZBTGR�k3RQ-��V���V�������ٚ�m-��e��l4A�᥌�`�V)L�-�ЛL�hk���p�"�m�
&�,%�ͼ��hʹP!�(�"� � ���X/h���9�--�	�H�ġo!A�6�1�.�i�D{`i�Ȼ��FݐS�ZuYh�ґ%k��u���`dvCl0�Aq������Qa۸ɳ�2Vь65�bb�Jt�]6�g�@��� Zu$z�lf�!n�X-�Eey��m��jQ���,�b�s�e�¥ n�����ҡt(<ˣ�f-E�nN�AB�[-����sG�����G�hB:;:�m��˽z�ǯE*���	�Pe��6Si`Ńm������˭��L�0@@�"�Lښ��X�Z-�6�-��6�p�)G1����Y�1�!� �c�N�BcY��͸M.�n(%؄�eu2�k*�m1��Дn���#�6��u�޳Xѣ4Ҫj��.MJU)LB�<��4of� ��e#��]b�Ԭf�Yl\6k�jIV�̄���I���Ra�м��깭ԭ��g,�ŏYVˀ]-�t�V�e�LڀҤT4ٻ[+Z9{0PE���2��^e�Sm+�
��-.��� 4�![Z&8^-il.@�5V�(AmF!�Û�tځ�2P�o^���;J7���3PU�rv�J*�J����t���a-�L�d� �!m�b�ҷ[$F-)eah �)�]-t��b�a�v��D^�mp�5\l�u�fKE	e��ݶe��	`�p�ء��2Ѯ,e����%��ɳ4KU��5���i�̲�&�˱��!+-�f���6k�)V�b2�e�L��Q:�Y@FB7�2l�e��V���.K���J!�mXD̺֚�B˙�&��o<�x��tjຫ����g6�����,�hY�57h���7�.2V�3���1�z�JUMg��bk@$c�4���d�`-���:jf%͎�`L��6�)5\3	2��l�"��F˙��2�k4R���YZ[.Z�S��A��5���BV�]ԛU���-X�)-]w��'���Mqv��W���i����/6��v�M�s,���l�

J3V�E���,l4[�Ś�v\-��I�<����j(݂���3P��ev��8���lu�Ak��LAX��۵����#X:��"����G�b��nf�,��m�v��OD�B��pְ�5fjU�ku�P����cK]o��Ҍ)�j��zՃWff��B���Gh�f�k�Q�-�Jnk�Kn�ȣ!H2����n�6����hM��[l."R9��1�vŅ�Y�D�#�]�1�u�D�&{f�arܠ�]��T)���#]ͻ��5 .SV���T�òM[IZ'Q��GML�Z9��u�� �RY�D���4 ����
�UЗVS��SG]t:���J���sH�K���e��`�l��#�R��Ҙi�K�����v'��#˩+��ta��nm�Ԙ�V��,�EqbJ���زˠ�xS�<���U��g����]���j�S7ZU���̈́c3hǬ�1�,b9�����i3����>�,"[�{�����,��wq�7Y!d��+M��\�v�m��V���Iݑ��"�m�iٕ����V[k����be��͝{g;7��Jm[-Շ�nv�z^jE�w6�.Ҳ��mY��n��H��q՝6٭��[b��,�-�o#�k��[m��ޙ�v^Qh��L�u���mMj,�Y�����YZ��6t�2��{�Ku��]�V�<����[����^�<+QZH%���z;l��of�ۼ�<���y�ye����:�aŅ��-��:�����ݵ���vdy�[ډ���m.� )�m���9�l�9�i�g��!�l�^֥+�v�3���e�mm{�k;L�%�k�&VQs5]�-��gv�����'kM���Fd��[V��yɶ����8&�S�׵�9F6���9�i���O{^#��iΠH�ZX��ԅ��I$}c�uƦ�14f^�F�Rc9�gj�"R�9�2�m
-Q�؛h&�vM1]v�`!�K0�n��ѳ1Ƀ&0�z��O7����s��M��c(Y�	��ZDΤ�%ֈ�X.�їR�a-\:�7'5�f#�T��jHPń�l売UqL[.+f�r��Mn	���6��ݵ̱!e��h�Ļa��M��xp�m� �a�m3r���^�L:6�u�&�JӶ���[]e�]�S���*�M�aq�f�c	�nr�h��D)wa`�葼��FX��X\�[��e�[yH���&Vmc5��[hXF�mrĹ�٘��4`�%4j�au������L+G%�f�&C�SBikJjа�F��gYa�(���і�׍W�&CdR�Xr���)�3@�ˑ�
���}z���B�)J)j��l,��[\���&UD���mD�[9��3[.I�Ɣu��M�M��Y1t�
@-�W��P����!u[{�	�^�k��l��K���]c��ci-�ci[*�Y-Z�
e	��M��ɨU�c\��m[I-�*cCִ�1��g9��n%ɒaf�:;�hk�-���b	%��K�Z$��hY�7#.z���Ֆ԰Y�,�.�ƍhmn���n�#$�7��í.�Ӭ�J�����v�@��0�Uy�hF9�������Z��ZZW2��[��e�R�!DȌ�`5��i�k]��K�0u���)����e�S;-[f�5�%ڴZD�!�����!1hZ9!2�j�/.ő��CW[tz��
[Bd5EnQV�X�ix���T�CVٲ�YL�G��&VT	HvK�M�@�\�W��4ɥ%S�H�SJ@��h8�5ɋ�CZ�5bKZˉ��5�&C0ogX�V�(2ꖆ(+�IV�*�,qa�s�S"�Mt.-c��9�f�������O2itbM��t��H�p팔��&خ:I$Y�D�[W��жeF�Z(��JF�!K@����������X�AK(T�jB�lA�cxl�F���) ��yb�Im�۪��4����/4!jX�"PA��/`[kYl)Ie��hЍU���Ƽе���KڂKR(�P*��m�������fX&�A�II%��l�h�K���(�K�V���,v�௿��A�qi�ED�?�<���ۨVbZ �8Nh�f�ݽ�����w1$"�G�J���
(�"�l屻�MO�B̳ʷS��Y��r����#�p$�,�%)Г�w���H!� ��>��I�������^M���vmc9�q� �p���@���3���A��5��&y��$�.0�+\�(ZUn��ȉˈCF��}4u^0�:6���q��ޑ^)D�	E��^)E�蚧rvE�>��Ş�Ĝ,��\[�ߵ���	#K"N� ��ޠ���<���
�,Wĭ���=mu^�V&���e�������Z�f�]?��Q>ߔ� ��U���IP���u�s���g˵�#Έ��Srq��AyB�q>>E�	*�JP$�CL��oNkȞN)md�BO.	L�K]T���px��g�y�Wס5�1�����-?.`�^���Z����B�0����sG�8{4�Ț�+p�_w"W7�w��{�7Pu�TB%�ܞ�e
�H ��2A	*�Q�AE,�ڞ�t�Un��&���@��H�D��׈!)�R G����Jv@�ǊJ���.q�C����e�����V��w]4O��~ ��>Ie
P$�"$����
�Y����0����2���W7�Wz�/�� ��I��y%"�,[A�_~�����i��m*�5�l�D�SZ��t4]ml�+{^p�68�;.�b�x|�[����\�^J0�QG�ާ*�9��w�o�o��E�y\�M�@gԬ��: ��� �Q⒚F/MԅC§�⒡CR�9��G����e�	����JE�uf�^j`��
M�SʠJp$���))�%#	2Uk&GMm���8�CU$��q�*���������C�y�؝l�@�v�H�d�_]�{�5 ��L*[S+��xeM��*��i���h��s,hҸ�s�P3�"�<��^)D������h�A����
(�,�NMnw�w��z��N�"���h��o���^O��ȐB*} �RS�P0��Y��f��{��PKT��l���mk5�q���HĤQJ'�V�v�;F��z���<����&¤�4`$Ю.u���J�˙�(в��ꌭi�PԮ��w
��> �O�J}@%"G�F��;}��Ne����f�8Ԟe��
��R0�A)@�22�*�1�oD�elz|R�!��nUnw�w��P �O�j�H:�ҡ/�:��� ��	��
R$�H>!%C���w3ӻkYٲ�,�k3#�>8�I-T(�H%(BJC��\)�WDT@^ ��>��MR�4#Rɍ���Ne���{���2��N�&1)��
:'&�+$��z���͏s��;��	ޞ��̊;�*�~���Y/	��x��Z�N�%�8��㋨QJ$JP'���E('o.�M�8���;�'oq6�*�;��@���)��A�>���T�6�M�T9�W_�c�6��[��5C[K��������i�34[��)��+1�X���	���� ��A�IPƓ��j6mSf�����s�����݌݀��tz|R�X(R�$k���h�FkcW��9��@�Y1���T�4ƌq�{��\��^�"(��D�[�[�$��@�A)@Y�M9�8��W[�c*�p���&�P>-��AT��� �$% GP�;�,ZO�� �Hş����]kBٵi��f�#� �>!`ad�z��/�O8	*�P$R�IIH-Q��%�h�W"EM�����Sl�1���4-H�BQ'�$�OYj/��y����p��Քf�ue����H�Cr�M��g�U��ʽ6�f�'�4ni��uܐ���#{��n�O6��ox�h���o¨��F���mB"�hԵ�n�v��CSn�Q�L[��n����, �]���R�X�Mn�[)�U(�A�qJ�2�5a�:f3V܃����s�K��`��Ͷ	Y��S��&uW�K�cM��HbfTKlCF�Vi�9.�+e�e�Lv5�Ҥڧ�l)�.��u�Q���i��f�	���N%�eW[�mM���bEQV#n�����߿��A4���0�]��%V�j-^e�[����Yt��4v�����|���sT(�@ ��	ksSsW��[�r�����9Ż���ϧ�S�$�#u3��mU���t5��PQɃ��J���u�/&�.���fGx�q�df���YCg��g �"�U�Q�))�P&�b�Nn`��B�͘v��T�4ƌq�/����BQ'�%B�Q ��w[��u'U��GgH��H%(-�M�enwin���o�
q�p<N4{��sz}O�I	D��%4AJD��;��.F�O);5uu�q�r�Y�c3#�q��P�����{޼s"�8ʦ�Aa �+�@��H��Yu#bY`�L��Š:eg�w��z�f!��%>��O�F�ɍ���
٦4[�_�z[�����fQ)Gt ����L~;�2.��Ɓ��_�-GK%�MMO:�o*���إ�R,$˾��/=�� �K9�A\Ю�0�k�
U��na��t����,��.��y��m�IZ(��t	ksRrr�;��B.���@��Ij�O�J]��zP��B�{�H!��-��%"A	D�T-���7w��:ͽ���1z�γy���AĨQJ$�
P�")ժ���_l �Ϥ�|�	q\�[���4[���څ�h�b+�b`���I�P$���(���:A�PB��	�ռ��V����Eדr8�	j�IIM�
�I��˙И��T5X�&qJ:ὲ��MZ`k��Acc��CCM�˿��a�#�S@�� ��O��T(gͺ���L�Y�����C���-�=�c�}��PK=@��H!Tb�Q3~�o������gm�z![4Ƌq�{��5 %��Ȼ�1�B�8�|��A	*�I�P"�H[I�����v��O,��TL�W*�XcQ�WQE�Y����4�ܔ�IrO0��\�f��ʊX̚!\*(F滩�mQ�ׯJv"�ɾ�
p'�j�S����Y�����v�R� ���ψIPƛ�̜�ɛ�g%��?�#�����e�f=� �W@�U�� JS�)'Ǌ�t�{� j�z�IW���nq�[���9����$$�(�N���o������vƙ0F��Sm�C`�v`�+����q���M����>�,��=矴���	J��n�trw���b.���CZN/w�Z'؃�������D���⒚UE�DOBn/*"�H>>֨V4�v����k�K#�A	��*R��ce���P8�+��t	��AIO�%#2J�\`��\:�O��4<� ������ψIP���3׍�̧�9e5�_����rg�sͼN�N��)؋�&�qn ��+&��T���sS��L��j�:�wa�7)��M�����ڣ�����C;}��3"C�DKF��X�'�E}��ETI�Y!�ß{�3]g�`��A�Jk����%ΔQ�����
	5�ۋ�dn.���;�^��A	*�Q��
P%ˎ�3idA��3QV�*P�f��4D�B����V�i�	�۶j�b�)��Q-L^=�@7�'��㻮��Bj$vww��HhyD6z�R[	gZ��"o�\���{���=�X����-��o���B ��7�x���zS�^M��[�$��
J`v�˽�(�lЉ��z�q��)J ��zpƀ��.Y�%��ȴ��PR��|V��>IW���	!%#�8�7�(A�����!(Pq#���ވV�!��p ��4Aj�v�Z3q��>#r$��N��`>J ���%6'�w��9��J�N�zS�^M�@-��BS��IMx��0�b�������f���T]�̛=rRr{2�S��=XjǞUc�1�J�:���u]V:��=z5��`Z�k����ĺ�X!F�Lڷ�C��x�i��b�UBk�f�`Fי���K�J��U���
GJck-#Ԕ��k����\��V��FmM3�s͔��a�R���gQ�̹qb�Y�d�<��3�XE�x4le�l:�P�r�5%�n�Bb;��˴�.�R�7MQ�R&��J�\�j��R�1al�7
Y��u������������� �e�u�������ņ5D��[�Y��b�ZAжթī���8q	�P@�
�.�є�񙮈?{Xdn�|BJ�[�O�H��]E�)lz����F�,��#���FJP$��xW��$D�K��\�Ϸ�4�� ��N$s+p��4<� ��4F�BQ���sO#}1r7Ÿ�:�I%B�Q �R��ꪬ~귈�2OQY6t;�-�ӻ� �_��t#u�����)M*鹠Fd	7 $�f=��qt����Z���w�(GY�U�����[�IN�BJE�I)�����F�N9�=� d�wk9��4[���9��"|BQ �%!Lvps�y��:j�Ҫ�v �\]L˹�H81Wf�.�4�&j�Y7e��M0�i:�j�=d����LN���N�f����\׵����`d�
��:�ݓ�:�hBR$�S��(����j�nH�|��5p�թSf+j+.��f�b����tE������uޝ���)4e�T��{Ѭ���(���&J��Fl��fv�}�zE�b�M�IG��	�
(B�V�Q6��������P �%)%9�
S��ݽ��s�5y;׉8"�hh� �4A�H!(RT(�}նS�U����
(�A(<���FooaN��{[�P � WK���������nMZ��RS@��I	A�W���*�
��ڷ��foQn�����%A)@����(uT���A"$n���n�lc��SD�n��5�Gp�W���Ŗ�Y�7�(���'����۬1JG�K��!=��q�p��ʸ�6{���g�rD���A�IP�R���P'�MΉ畸�c~�3��wd�xR���w�[�c}����
Jy�ݙ�h̡�r$��A�h���!(RT0y�&��Ѷ�����UvoL��f��M�=���ڵ�Зݝ�cJ镎ne��F��*F�akw�[�s&��[U�ۥnZ����.��A���y��K̙�u¨ٓ�Q�A@�Y�]�V��U��Ce�O�Ъ�&��T����Y�9�X�»���]>ӱ"uD\�gr�M�z�t3.̼;��Q�ah{H�a�oR�����s�w#�f�B�3q���������.
�	܃h^^fLT8��(��帨fb�W<��㛛w���q���L�F���r�2���.��Q""�z���r9�EuU�]�y�LwH]^�+j=6�:�M���^���K,�7��k�Ř�#�ٷƓ�{�c�5��g�;�%���1�۰����+�˶���9��[o�Qzn��o]Ǥ��h����8ܘ��)or.��"��"Z����CvYi��v�i
�x�d���>6:Ƀf!P��$it�j���Rt���{B���`c"�V�.���[Ȍ6&ω�g�b��+�q*�9���N�u%p:@�T�.ͽ{Dp�Ծڣ��z���j����8���֧v��J���9BWVR8e%L<��M��\r��2&M�e�\�̗{ʇ0�-視#r�h�	Z�u3r�J��M�Z5jH��]Ԗ�B�ңWWU:��E״�ZO�(L9�uYWm�MH��fR�{�n�:��{�yi��o����]�]b�Z׊t�����f,���Mb����ڙW�\�⧫(U�]0x�u���u��e��Y�7*Efȷ�Y�\���Q7�Y�n����p��lZb<|x]��X��om�g��ܑ��^�{7{�C��̄^֝��Y����8HI�{w�T��i�{���Non{�I{i�.��w��\��y����3��{c��qd,	X��aKѤ$�t/o��͵�����-�x�����^[��	re��76�ލ�杚6���,c�Ŭol�Ŷ1����m���zۻ7a�'kyen ���֋;ON��m{V"\��Ь���3'��3�9<4#��D��n�mM����2�ZOk���h;ipaם�ǵ���2#��zrw��q�I��֛6ץ��6v'�{l��Z�k7g6����X":�[�.����O4����b�	=�E��/5m�(��@t۰�[`J򽷄t{emYy���mn�Hg�����z��V`��[�j=��ڽ�{����=�$�V����+�܁�6���=��vݽ���A)��ٚ�֑m�]�D�6�)�u*U��Q��Xʂ+�]����ٌ�t[��G A8�I%B�Q�(BJG'{�j]mͥ%�d����k������;���"!=��q� �nk�N�E a��̧�1@7U
�J���wS�N����a���D'�ܷ{�F�oaN��{�@�[�%)��wu�����*>�AZ�(2��A�7m�`e�bm��	4J���Q�L&��tV���Wx2`�x��"HJ$䔌j}��l�d�=����4����H0A2��� ��	!%"�R� �������y5�r$Tlj�����Aq���P�"A	Gj�xn"�g�	ݡG�$|[�$��E(�	J{�%�"��K�����s^����n���S�%HJ=]���u��7��]�R(`i>՝6vszKpu(�A�� !��]N���g2}���xT��r�Q/t�^+�C��b�v�ڧ'Rܒ����p���8�3졔�x6�/
��^&͛�L"q��0~� ���(�A%>��������=�,;�"��3��؃
�`Ћ ����>� CG�#tr��R޾���F�5N���B�	Mi�^ś �"Q��k58l���%cjrC?=��N(@�t(�H%(9��tc3�l'b潍�ꈫm�k2��@�A��u��%"HJ$|RS@�&�$6�aJ5NzF�)@�С��}�:l������Q�	��%B�Q[�xz�F�	!��s�� �%>�RS^!(zB��7u=�O+'�[\n���4A���J��A�N槶��h#�H�PP/��q:1��:�3^��w�p$F��܄b3��7�4A��BQ �
Jk��O�J�sN�U�mD߰Em
;��Y�Zgw���q��S�%(w�wzaJ��NE��^��t��߽^��(f]3ŵL߮��%��}��-Cs�q�����/��8c���U[4ũ�T7xYH�vZ�<�1�23hQ��ٹ��m�k��%��6�F6m�v�,\���YIF��$thq�LlAk�CX�\kUi���˲��0�ͺ�(F�+�.!yɝ��X̽uU��G3���.k�6C[%΁�z�wl�ۆ�M�Q�%�%�v*h`���'�ii<�î��=��#n�v�\�(J̄���S�anZ����g߹�nmK��-Xԕ�mE@�Y�J1
�j;SJ�j�gBXT��c��� ������D�����]��T*f�1n8���
*t:�9C��*{�,� �p���F�P�4)cs�U�+F�yA�N{��ٍ��ByFk��P �AG����뺨��{�@�>榀 � %�IPĦVK�,t8��W]ά{��L���d�Q���BJ��a�PK:R��te�� ]Ǚ|��BP$T�NU��T��b�p ����rK�K�m.��ta� ���B�Q �R�%%B�R�����c`H�]���os�)��c|(�>O�����v��u���~?�����(���b�2���.�.��m�+���M6�΃.�����7<���A��#I�nS�;:��'��F�R!8Z�P)���J Ie
P$���]�l��f*�P��iQ��5|��	��q]L���Ǻ顽�o*]�E�f�=��4�
�XB�{vi��T�u�TVC�6��9�h}�D��]*�w�*ft1n=�=�h�5ȟ�Z&�hZ��`P�T(��H)*�Q� ��z���1[}�����S�3^�|([� ��S�����O�L�
\��Ww:�2;�> $�W�=O�eua��s�J8�u��
�4�t�^��$��	#R�(�	� �>���y�RL����uԉ�AY��Z}㊙���	|���`!(��hwz��ݩ�mߥP"�$�-"�J�3,oj�s�c�Y�t�]��Y@TIk������|��[|A��E(�)@���Nw��kޔ]}'z���!7}a˓܇� ���s��	@�BQ �%4E�^i4쾛�9,��&&��hP��}���G=�0u(��p%#
P�e�G	ڽ�i��5e
�P'���RS@R�d3+Ըi��hiZM�#�U+t1�n��3LD����+�2��ͬ{���=�h���Genf��D�|�"���ϱ�ꈫ�?�4E�/����6���A|��|BQ ���P)D�M䊹7}W=�E�%(9n��{��V��W�_
�H�F-�m{OvMGt�%A%4!)BP��s�U��z�]
9>�Y�l��,J8N�AĨQJ J=
��uɻV*�DUP,�a(2��,�chl�׉Y^����e�-be�k2X2&��=ޠO(A�>�RS@������yU��Dm31�8���5�N�͛���IP��I�H��ɼ���`�)��`���I����z��Ѫ����� HO����X:�m�%hE�����RRQ`��%^�(wJ�nZ�ؑ�9��;����u��x�'�%|� ��۾��
�>��A��ⓚ �"��S�W�ȍ�fPc\w��9�9V�)WF�슺Icm��3YUuT�PL����T#-F�#��S��,���Qws��fL�y�j�,��AH�o��)�LF����=X��!���РR� ��	�	)�QSե��o�H]ݪz9�y���5^�|+ϐ`�;_��tF���^w%�z��1�Ѭ5�a@f��iFX��
�6#gk4�bܒ�Mm��@�'�W�������$=}�t'�wq��J���^Xͭ]%��@l%Ml�.p��
����X(�	#��gg�]�� ���ڽ�DW5�tÙ^G=��a̲��i5�cd���%�
:�A�H ��y(��FElԕN�:wR���9�X��f��}��	 ��IIM�	%�nҢ{kpۖ9�qg�%B�g+�E����X:�q�\ �z�Yμn;(�ǽf-\1�\O�%8BJ�^J�@J} ��8����P�'�C})U��Dm31�;�_9��"A	D���^�P8�p�Y]U�&�KW�p�1KF�a��D��Rkf�	�)N�80�9��&Z��]Rig+n�6��͸v��wW�z��k�8Ü���� =��L~�=_�k6�,�Т�������T���.�T�`�ٚ�9
+���-�e%�i�P�ܠ�������vr6R��͆\^�.��ل\ 4�3��6^�cH���]�X��QH�V;%40�DF�ٔ�,;E�v�-�.�Vh�)�L�`�M���z�����I�eH�;V���	��Kn1 �;�պFk�����3�k��c���͉Ka�m6�h��&�c���+悧5���r~��u@	@��wWR�J;ktj���b"(1���>�>�]>���!(�A ����T�&������@�F\H>#�Р0cW���dmj�,j8|�A�
�J9��M��80m�
P'�������TE��A�R��[P#i�A�q��}Z�H% O�T(�FY#��of�� A���=�(9n���R�n�׷\�(}׻Q����sT�'"HJ$AIMx��>!(��A���(`�U��Vd�jrX8�qp$�1*R��G����9�شX��-ҷ3]��``�9w;F����a�.z�q�2�Aƀ*k�A��z��	��%8J�z�����b)�A�pҸp�]��@�9���E(��H V�RU�a����s�y�fB=�x= ��Y��x,%K�':tu�O�6��p�h��J��M�\���ֺ§�mё�po�����Q>>�H-���{�r����{u�An�j} ��uogfuv�J�"R� ���Ao��AJD��I�IP��p���������+kWI`�P(�dw�Q#��@�UC��Zћ^�d�Hq��s�F��^��V��i�f�c\p ��h��z�qD��vD��
�J=>)@T(�{*� ���t
��ѽ�^�vf�����n�Z�IIM A	Hso�N���	�~��Vq)u�V����l��d��o�.aV Ĕ�)0�OQ�~��}y���P$��%B���;��^֮��ƣ� �T�l���\
 ���Q���H!%B��J�E�m�}��N�gz�\��A	ȟP��U��b���^ ���DN@n���Y�k�7j� f)� �� IH��H � ��LƗ�5�nMEJn�%��n��ҡ)�"��������4o��*�p�Ie��s�%(���P��U�+PZ�_� {¶^�{�_,�n�߷_�AO���	@�� ����ݒ�] >�>!%B����y{)t�5 �A-�S���9� s �X!%^�~;�0A��wuˀ�^F�WF ձzU�oF��i5�K�4A�"|BQ>>;�B�G.�Lp��:�A���iQl6���0��������R�iIv����b�h������
)D�	J�������[�7���p�q�]^@D�>��� %"A	G��%4E����j#��"�#�X;U��sr��,J=�)�`���+㺞>�:*ł�5h0FvP�7A%>���P�R6�*B�պ2VVe[yё� Ƹ�J�4:�O�J'��)�Q�"�E�msQ X�B�[�IJ-��6��v�[�7�� � �Q�m�����Q.��4�	��{i��e���u�F�o_1.�nky��.��ק��Oާ�EEa�ݸ�NA���&M�;����j}�{���!(�))��>%�飪O���
C�Wǖ9��\�6�q�JF��
(��aOs��z�6�M�
d
�
�SF$���J2���h:�ŗ5�*X:eg�wϱ�}وz�I�iM��"�Ε�֭�f�cK�T[x��ΡN)��#�%^J0J(�"D�{Gy�9У0`)G��fG+��'r���7��-��\"$���f��t"EGH�B<}˧<AJ@E\x��|��z��\��<��\�7�8AN��H��H>J���P��e\���� �I�s@����s�l��|n"��� �s��9�Bg��ψk�W�Q> ��	IP��h&����s��:g����\9��n�߷Wz��A�p����!(�)���\��
h:��͆�eʵ��n��*.��1ON(�l��jΣ
�@�-�J��#Z�P�("�L�D�!�ޮw��C>�]�3Ud�0�v��R��j��F�ݬY�J�w��H�e�d��H��C%ҎJd��[�z��C�S
��p6�c&�����ãtk
�˰��E�r��m�ϑ��x�R�g1�ԯ�*�N���Ky�N�J��g�[C/�IĨ�V�P�L|hgrwUPYq���V�]h��V,��=�R��c��-]#�'z�;֮Z�����Ub�s��d#����X&�ι�$��1�7h���t�ګ�c�=3vv���-aحw1���U�R�0)��L��LK�ȸ��Oo�M�i���uOi�^K�kxohM�2i{���m��U�_�`����T��U��bŽǵҍ`���B_Y�{�W�iQ��V�}j��0nut�����)6��U�­Y㦕��rB���-�R4��f�T/r�Si])t�R�qzD��������ڪ�o��s�ciu%��J�0A5vPSF#��뜼��m�I*8{s)�I�_c�[/��ۇvssd�ڷ��lټ�U�ܗ����v��K��]��G(�י0*�s�4�Z�hU�oT���UĢ��P��U�������,w��f�jOƃCD��g�8y/x�`I���$�N=Dwg걙��=D���}(�(f�D.�����m��p�^5�s"Ѭ��n�D!Iղe��ә����&��5�N��T����>[�W�'Y[WTaN�j�s�z����-_��8G8Q'6�\�{Z\似�D=����$������m�I8ej^�aǚC2�&[���N�9�,"Q'H� ���헭�����ݔ��k�6�����v��ďk �ӓ��q�����gY��(���܅8{V"�{b�P�ȑ'^���7G$���w#���(+[N��h�������.I�L��
^��;m�e��qٓ�<�m��ff��� dFՒ��Rk�-N'z�9�d�2�m���" @#��DP���D��r��v�S�mi�gD�87��򰎒�"۳�;I�Y��[y�����Ӊ�{^4��wH�99�!�DH{i�N$!=���q����s[p��QNՂ���Ԏhͅa0�4Z�6�)d�6�f��X�Ƙ�-�5�i����mT62�u���k�ĦP�סf��Q�m�`�;�Pc��e%�Z�Ζ;"�P�B�����l�6��H��C2�WH��c22:�E�M��2��..��hK��VYM�R��MYH�����ZJ��p[��=�j�$��),�b�t.]�\֚3;42ͥ�[���]uXU2Y78�a�Z٬��1�����u��ř����
�����+e�;��kl� �8�u���j�%F�����)*+6��Xի����)����\(j<����Vśm��R�2�]�Ч9� ���fkZ(��ED�cpicf`R�[
f��f��V�Ě�$�tu�ƻ��Y�A#u�6]���-��32��)ӭ��:ܚh�Q�H�II��v�.$S3[a5���0��4IBM�p���.�sŤ.o.�7RۡAK�kQ�g�Fe�&�nE e1jբ1и�t-J�����Dw:b�3��y������.��T�53#��1�cT�\:5u�����:��I�C@3�)�@�nn���M[(��p��l��6����ZД9��&��3(ˣ��`��ƷS��шi�TM�"V��h�WE,$Ι�+�st���IB�`��n����a�x�X�K-#@�n�a�MXi.A��
��O^�$��X����\6�k:�&u���[)�fV���(	c�vs���ÌVYn��CMc�#�h���f�t5 A٨SK����f�D{J֩fd��S@��l��� ���^i\^ۛ!�JU��k����RCs�h���԰q����L v�U��(S$sv��`���+5�a3Zʬ9�����5�P�u�ꖛF�a��%R��.�i�ye���S;Q��؀���"��2�x>�nM�D��M����Ё-Y�\e�4��Vfh�<ܰXSP��x�6�jA�0�In�rVi���i<���s����ӧx��]��dR�\��Z�����k�2�f�֠�-dؗ�;�.
�XD��f����Y��Wlō�-lV��B���u�L۬И��r�Mx͖ƶeIMAB�ƭݯF�.�]K6�=B �kG_wյ�Ea�RU�1�^� ��%֛-&Y��<�)��&�t,]@c C��j��R�mF7A���D��kafP�[s�e-�v�������7;Cص�VЙ���vl�ε�3��.�mL2�]��O����r� ��$�>��
��+���V�.��G�;,ǩ�8#��Et �7�U��P$�|37g#1�k��! ^t� �"E��c�[�q� ƖG�h��D��Vҩ.�bmТ� n �T(���n��r9N^n��n^�tf���P>-��j}%%4A	H��#�ˀ��@�v���D��H>)*����o+gK��5@�;=7�=�1L"�I�$R(� HJ} �����-�ny���5�z-��񴥚A�q��s� ��>!%BT�T�z�/�>�M�+�����6�+WD5����Y�i��+Q7/ mL�j��~}O��}�ן~~�qJ E���r���7���P��̫���m��Q�3����Xdi�#�)�W'Ǹ��yvP���x���Q�M��uH�nV����Hg�F��Q�4��駲�':q�#*
^�n5��jы/U�m)��/�xx{�&E��9"<[t(`ϕ�y[�����z���gӍP����؝ɷx�[b���s�ѡ��E�3�Ա�{zD�XB�zSS�2���]{�m'ƴp��>+����D�R#�$�P)D�2cS��e&O�Q}��2��6�3�q�rf���p��ɉe�*����EH�|RS@���"�;>�|㶹���
�����V�.���QfAԊ(� ����m_�J$�|���Mnx��k��.[�q����ʫE�8��C��E��F�V~�ᡎ�G�Ա�{tBP&��ծf��%�A�_ �����N����I��y%"�Q�d��Hڲ.��s("�H�Y巼m�E��Mɛ���W��'��JHɚq�~��'�YB9�^���i׷Q;����=�����c�PkB���y^�E�����U*�y���O>y�"Wu��\�o}}#L�P��^ŒVUՅ�&�Bu�]����T�6�6ut�@޸�|QgӍW���������/#�/�B|A,!��t;�&��Վf��e� �/�W9��N{��w�4\�{�ah$b�3�y��E���6{2�v�'�[rg=����	!�|���	@���j�j*c�XGb�YF�3!L���2�hSJ�AY��n��Y�$��Т��s]��?_�T0ct;�fl�r�z�}%�m�Y��>�T(�A�E$�QJ ���}sn0��[��	ȟP����c�̸�E�W9�Aj@E)�{��W��
Ȓ(� �J��zJ(�p-V苴����[rg=z��)��%j�W��$"��QFT;+e��$H!�"<BJ�`��w.�����x�>(�$u���Pl�W�p0�/7��f=��s/����2���T��M�^��'�������ڟ]�WVb�y�Xγ�w2&��*�x�9.����{�%�>��>?!%T	J ��%<,�9~�w�:�+#)�\;ˊA�_@><��5"HELx��R�eWT�ߞ������3(5mnъ��]5�LVf�-j�F+��(P��ku�Zef�_p���b~�{߻��EosG[�#���{qH[�/:Cǻ؁5�4�C"Ao��A�R*���tp6FGR�C�g�9:�9��瓻z�Kb/p>E�O��
P����)�Ę2}ܤaN ��%4A	H����Н���C�ԗH0�#�y��� �Q�y(�4о���⏷��^+���	�{�:��ђ�6"o׫��	#�Vʵ���3,E��������%J ��3����B�b������lE�p)��A�M�Gu2	�_(r��{[^/�b	��&�:�P�B��&��\�s-&4����'��֌�u�#7��K+1J���ʧ��Rh^��
^wz}.������wO�W�J��rYn�b�E���7���y�V��0�6�]V��b`У,Y�XДGj1ٗB�s���eu$.`;��ˬ#���\+6�l�	�mfƖ����PK����@�jul1�1�G8�%n���u��[��i	�Q��hM�T����V]��f���#�n!2��,�),�u4`�ܱt��X���AԔ�0:M�y������mkp��%W��]���Y��#�-V--�$�ҫ<�|��<�s�����@����M�os���] �q�iQ|�uѩ�D>'�L�!�#�I�	*<R�H)@�FW�/Vj�e�H�{�z��Na�lD߯�8)O��%66&�k*gz��}�7���۫{ר���bw�laުu=G�E��X�4�woy�6"�Gx�S���>)@�T(]E��1� `�I�S^ �"E����Lv���� �jh[�Ģ/i��7 	z�QJ$%@!%>J:�ȁ�~�(+����zM������H��JJk��:���w m��ǟ=hnηUH1��e��LGMRSL�(��6��:��c�c?��~��~f�}�>!(BJ�`ϝ��y;���x�҆[四�
8v����:R� ����@�wPd=ݕ[�}�"B2f]�Iw)��<q��������e�2���i�8�[Blw���8rY�5ٹ��lR���J��V��i���� ��O|_t��D���fm<?!�'���AjD��
�%�IK�;{\aP��P)D��(k�YWu���-	k�CM������I	G����)(�엔Gp�UZ�z�P �rD���	*�9����{��b�{�N 7sIɕ����g!g�'���$��P>+P`wX��ę>P���@��Ø�[3j��2 �q�@<�ׁ�	D�⒡�\3�+y\m�����ȭsXd�d�<�r�,(,�1����H釩�b�n��E�� ��A�$��ua�=�a�ry3�b+=y�Bs�Cil��@�˟O�� �)(��Jk�uƪ��v���q�>>>��P���}�sv�-��q� ��H!�^)Ex���Q��r`I{^�Kp$���RS^n���ߎ0�j]W���V>v����6Z����1u���܌ۦ'e�st�8	7��]m����[�˳.�B󯥒Ω��?+�J����_1K2y�M/�}������gT���A����ܦ��A�F�g��b��`�i{�f`��3�"b�'A(9���tDklMg�7�^N������^�^9��I	D�|��RRQ�T	�����ﺅh�>�9�|���^8�A)���B�Q>>�B��}�4�z�b�f��F��Yd������QS.Վl�s���m,r#��,��Ys>��J�CS�))�P0P��j�[��H0�q�.e��ꇉ�@���!���T(��� �1��۽}�G�$�t	绤u���!��Vz�z�t	��
JA0ռ�^	��`�
�4J J,���<������:���������.��	N ����I�|B�T���ޣ5�N����R�9�R�٬X��!�'�o��C',�ʬ+�#T��_G���N��|�nGRR`�U�U�7+"�S�բ,,�kw�Z���w�iܼΦ���4y7� BK֏�fU�{�hХ|�	!%"�J6p�=3�W0� q@���![�A�К�^�
�� ����R2��۴"WtPSTz�TI���e��wX챻93 �Z�� �(8]��L]���3S'c�����k�� ������f�	�b�\p ll�]��db�8��hP-��%HIP�|
P$��Xn/"�II��)H��)9٬����'�=�4AjD��H��"f�vY�������^/bH �$�
(�A)@�˓P��"�l����i���ޯ.� ��S�����X#��\Ӽ����X��D5"|BQ ���
���>}7����޸��pɥpq��b�N=%8%��JP$���RS��*<��W��z܄l4�&�����'A;��@	@�*.Por{is����8�ZnVnz��ț��ޠlޫ��o	!9�uP)N��p��Q�I���shP�R��q��iI;��|/�*�0Ɖ3i���P`m[��;l�=�*ĸe���5Ж4�GK_�|�<i	���i���Ȓ�l��A]��a�mt�4��@�s*2�6
�.���5���L�ζBl
0��[
�H��q6�5ՄVYe]e�F`�[ۮ����F�!�4����X60ڮ����]�gu��M)b�K`�\�C[�dB�j�X���GP�+}|�����p8�m�.K��6��%�-�9�,ÞI\м^8S�e��5�Vo��B������
)D�|R�>kti��=]��V{sxP-"�wet\� �l�A����O�J$�
Jh������cH�|��X1u�˦��w�8�N�A��Q�Y�}2������P�N��
S��IMx��n����2ۭ��K�0 �q�8�h� �Y�JE�z�'zkx���@���G��H{��gv����B+=��@���;\�o��Y��
ޟV�!(�A%4<BP'�%L�8Yy����S��r�̮E:l]�%�#uРR�R�EF�'�������`�K�,X�h��69⹫��]��4��h�X�ݚ��J��?3��ݘ��s�))�
R(��ՓYz���7Dڸ[��g��"j`�F��۫%(E��&ݼ�ky=����N�.궧C�W�����0�ה zrz�aQ��z�뤔Y���ۡ�"wYy7ݢ�3���B?�����G�Qs��?~����Nu��[�@��$��RJg1^�����%"A�A���)BP���^�WsM���d�q�̮E:l]�A�u���A�A	*�.�/49.���q��z�)*0$�eݧ��a(�8�h���:�0���	�
)G��(BJE�A�6� ^@��\ǖCe4"sط�^�Aj�S�JGgnW�ʠj��v���j�Y�1��4k��L�����SB�̼B�ꪱG����;�%|@IP��[<����N�mǚ��T�!����A)@���E(���V�3�G5��j�N�]�c�������#\�%�ݫ���r�G�$�u@�
J��H%(ú���O��2ه��$ŗ��{��n��N�ν�έ�ۺ��yk-�LlT�+��;���VT��K��3%���H��@���u�%�1�����z{ǡ���\�Q͊݋!��]\^oe��J�s6�໿f7T�n�S��V��r�$�,gq��U�����*�&�r�D3p�sq]�5{� �d@[N�:��0�+
���[��^B�4��S�lN<�q�k7���&aeSI��؁��5x%�rs9�p�u�3��8�������6����.-gs�6vr(�'.��:��Ƴ����L�a����PX��h�ѭ(�f�W���2��XpH�%L���L�ʥB�l��L�̺��x�GC4�lVFxV���vˬ^F�Nۆ!�MN�R1b�p8�ݴK�;��o`�s�c���v{)d�n,�6��T.d�T7��	����6��B8�Nfj+N4�d���hB�s ��y33'71o�+�0��6b�I+Y��z���.��ݢ��:T���f��s]��p��S�c{��v'��3��n��E^]�Hާ�vf�M��Vfl9�iTյ�&xAx���Y��,��Cd�F]Y�unTF,��-�z�g_rWm.�n�	�Z]�<rfŧθe���x�ͭ���͐nm^�=il�yy�7:������e*��ny�Ƅ��uQ;�nZ��Ƴej�o��ɷэ�U_f.�M�;�tCj��e�}�;�
�]��J�{X/4��B���Y���t&t�wy2��J�^��x��ej}ww.��[�-ꓷn��I�s�Z�*��k|��;0�ު�)7J��qo�?r @���;�G9�E&��ؼ�K��u��Ⓚ��漞��ڗ"E$�"fVv�{V8�j�۬�.w���yK,�m�s����idۗ9��7��C�vے�m�-gI����+޻g^�[�q��<�r�۬Egk�{ޗ�����{�I�)0�٩�r���Վ9��^V��yh��ynG^h�Y	Y�X���9)'yzt32G�ښg��={rs���q��Ća�N���i���-�@�W�l�ȑ��es,�yؠ��t��{L���b�������{iM��5m�s��݈��{%���n���w��"%m��A�M���#���s��K�^g	;k6�Nr{n3��F֝=�{�����,�-ds+Y��bߨy���RS@���%�9��8��� ʌ���G8�⒡^3]��6�Bv�]�|�	�"�9���$5Hԫ�)@�BPJs�����ˡ�2$�-V���&�J o'��9����wv�40�^Sΰ�o���Wfb����3u�6%
jt�5*c���F�3e���
�ļ �0A{k�ՄR�#�m�/�,�ek19�[�'���v�@��E��@:����$%��<�S�:�]����o1B竎��Sғy�-���O�>IP�R��}.�L�I��ٿ]�ț�������t)c�#������,,��˾A��-���5�5�	@	)�h��&�"��	�e��q�����m��G+Dߖ�P><�H#�ߖ�|�w�R�Cj�=�-��$��I��t;�	U�Ø��3iY��-F �LB:�ۧ�B�w�����Ϯ�[˫Xe�p������ކ��9�k���$%|���D��l���E�����}��4kw����u5�3� ��	#uH��?� ��U�r�XT7MR4�2��
��V厚����m����]����9U�bh^��˙&��H:���)`I��ݦ8�L4J8���y�̍5@�ǭu� �� >�S��^ ��I�3�������eǘ)��ݭ�w#���7����$��} �b�o�ȵ~�3��=� ��4AJD��>)*�j*���帢);{������8F�B�)D��H!%T�H�e��@�5Ǥ��	G�N�.�X�P�a(�7�>,�˛ovf����"�R�O�P$BJ��n^9�"��(v�s O�u ƹ�s�ƹ��<�	]H��
Jh��b���xz
َDb���Z+�u���-�z̪��#U�׷��̉2�c$���ZyWw�H(���s1L�D�6��%��Na��f��C�B���zt���������vRiWmn�4P�K��fe�4k�h瘆�%�&�pYMj99m��R���d�[36J;
�t��3tʹV�L���fj���m��bL����V,.����m�tѹc��E)4T�0e�ƌ���Zb8C���^��nG��aE��Z��eYR�ts5e�nR1��2�L�Y�k�&4�[�P���`�:��}��&`i�ٶ��RUε�V�� Bhe���K[j�q�|o~��Z�ܤO�J$���
����}��h�n;�m�I]��v�s����
���R�>$���J��t��tw���ɢ
�oN�]Zc�ECA����t�kub̗Kb�m}KXߎ�dg �?n�
;��Au=:�E���Fޥ��s~y�=@�p$��}%%4B��E*ʢ\�Dշ�{�����U���DWu���y����	j��=˅���kѧ�O��� ��
�P$R�IIJ�sS�5ڲy��r�Yuk�R�j� ������I	D�%�P���}Z�.�U0i�,��&�L�B�m�SW�9���0YhB
s�v�i���^�=��> �t(�H>J���'�i�37�k�-m�&�r��j�O�54)H	G��%4D�J
�:(s[�*{
�z�i�J��:�r�L?@x��O�.�-�z�;r��I��SnK�P�]�j�o���՞�xP8z[~;���}��u �p/�`���E|�5me�m� ���%B�J,��tB��|�0�\ �H�w�O�>J}%%5�JF_=�̜6�`�p.�ܚ��&���h�P$��O�IP��{<&.��z�U���L�dCw'93p�mW׼�=�2<�/��g1'�=>���@���w�b#���Nvý��~㮲n�I��+CM∥ݚ�nދ��>#�%A(��$h���@�S+��[Bř
֌��9��R�֐h:��gB	�mQS
����P � '�����%׹4��7L�ƨ�iHZҭ's��A	ğ$�QJ$%@!���h��2��I�(涴 �Ej���LW��W@�A�s�%4�w��i;�O�n$N���	@	E�$�D�{T
�a)�ƶ����S�]�uG�Yk-�����vf��ƃͪ�t��fku�ﲉf'���3��hM�Ω�wV�1=NӷL|��� �r%[�dکyƩ8����F%B�Q��J���
��[v#����A������>5e'{�I��qL�ƨ�AyM"ɜ[��0bZ#�P��HR� ���u���.k���b#�F������LW�}��t	'>����\#��Ʒ�>����RD�6�h��ۢ�.f�.�h�[�Lⱄ(���tf^
�+�����>��$% $�f_<Q��UV�q��_]�m�x��R��<A��wS �R�>!%T	J�:�ڮc#;<�q)��MYI��{�n��j�q��P�%������楆���(�L��|A�J��I���,Z-^r�����y������¼�������J��H"��Af�;�<E� �X>)*0b��.��U���'�A�C3
�z���
ᖷ�uɓMfì��C���Vv?S|-��	�Y{�6�P'2�	�tuf:s.�F�ѡQ� x���������
�HJ=%%?B��sI��r$����V��[�(1�8�j��I	D�$��1�h�M����P��k�;R��vc��0�L���k�S����:�l���
�>Z � �I���L�R�#�ֆɧط������p�l:�����} ����H�BQ> ����۶�1�uf����$L�بW�g&1�]ת�o�n;�8V�
Px�EJ�T4�@�/�P'�	% $���9��e�VGfZ��{�-�0�k���v�#��pNv���{�B�z�>�Y1�f6�. ��B�]��	�[�e��ط�F���-��}J�w׽ٹ�&�K��>��BPJp�R$��6���U���5:4owfWuꭻ�f��� ��$B�B�J$�(B0�}�:�71h�;�s2:)Ҫ��Fl�ƘX��EA�^_��+�j�!�Vv2��%<ٹ��Ǔ����(���<���?�l����+7&,ٶ*�48Ժ��.��a�-�	�W�)X�I����]3�8�hˊZƠ]�VQ�CDZYZ�*DEֶ]�{3$�N.����j�Ƥx����\E.�ZkC�1P�B�V��-ڕoVDb�7m���-��ͦ�0ј&�mJ���p�fb�6(���j^��{fWPm��f,�$8ṇ�7d�ه(����8Uژ�+1���3�-#^x�F�vee�FЮU�6e/gue�������6Y��RS�)Q����V�(w�Palp"��Uә׹Y4!�#\O��	*R�
P'�#lu�8aEg�{�+��$�W@��hC�'��#=����	������߱�3��R���w?�u�F�g�ݡ�9�PA�c4��U�x��q��^���W�Q#��	�	*��OR��G\�Ӏ�R&�^�Ie<���A��� �]4GoQ���z;�S�'[�E(�A(B�"�J-T�K��L
v��&��4�p�g�|(�	��
J}IH�y{�h��+{�E0�N�h����ڎ�����j	v.�ɡr���W\��'����Ӛ �$%�	*cc��Z�n��=+�"Ue�@�X�Q� %�	*�|R���G�7v�G��n�E,��%f�g�:�"|����.��.�ǘr�d�53�j
K�B�]�Ze��K0m��;��8i��"�F�1MW�{�I������ßvᤂ�P���(�|+�'�M�v~
]�>��<.v�>�) ��
aϽp�AH(�Y�����As.�j�]�:��+�� �T5�������i�) ��%>�� ���Ci �fQi8!I ��p���Z��D����:�m���l�g���O����
B��=�- ��Z���H)�
a��3l��P�3(�Aa��\˸
AI�����fs����(�L?s�2c) �Wr�$���]�R
A�C3.Oo�����[u�������I�2S���P�JH,7f~>׾�o�se�쇒
A@��ZO����_e�II�fXlv�R
�3(����RAh�֠)4�L32�f�*�s�w�ɤ��!�Q���^�;˩��σu{�8�^́�>�RRßz�M���P(�Y���R�w�URJ�f\6���:���X�Z��d�1H��e�٦�s��˭��!lM9q����6N�b���;i��k$~��b$P�O=wCBJH,(���6�Xm� fQi �i����+���4���y6b3�H�'ß�>v�R�7������k���=�- �(�$�wZ��ЁL9�i�) �HfQ���L) ��a�
J��p�&�I���>����H,H.�������k���}>G�7�y��e��⭺�g�h��D
H)�n�(hRAaG35����E����~�w�_�����^�L��\���hJH,?s,6;H)
�2�H:(�$�3Z���)�f\4��JH(�܅�'�>3�K��r��52)?N��]
QiY�]Tev�����_��ה�^x3�w.�������)j]����La���6��u�;}3p�~����W<��-ը(~��<	{2��
JB�s�\4ɶRA@��H,4�\˸� ��fe�i��3(�ЁI�wZ��<��rJy˸
$��·���������hB�%FS�w@�߽��xֳw����������AHQT�E���Wx��w����Z��H)�
a���L�) �Q�H) �˰�0������p�&�) �Q�f�CI̻�������S�� �B���i�Ӟ��<�{�w����U�h���Y@�O=wCI) ���桴��q� fQi4!I��S�w@It�?�Tv���ا�
^�SU2&N����i3v�9H.%kyl&�Q`lAQt(�LS�6����Z�]��U�E�Q
H-w�j�SH�3.f�JH n��O�X�u'���]�(}��Ae�|
L�o7z�}���X}�nd�) �Q�Y����IϮ�j���j����l
@̢�H�R�wH)��~���}�����/^��F��E���_�3�	 gc�c��_����ρ#���a��������D) ���H)�
a��3�w��p�<���(�Aa��_�vaI%S�.d�e$
��i ���]��TAH5*�p�A]Q9��1�d�W�F_v�������ޢ��
H,���z�����XT�桴��c
@̢�i
H)̻����3,8;H)v�_޽��꿹�+tZA�D) ��kP��)���ᤂ�P��i O�����eӵ%�8�q́��I ����i�l�����ӕz3�?q?&���@��ꓖ�ͻ��E֮���:�K��/E��TJ����LCkcB��y���ܴ����d2?~�u�y��H@�����
AH:�w�\6�]�)2�M RAeFJs.�(i%$�������-'�5�ܺ������Ad��7s> �Z�:�u��o.���<	�}��i!ATz�H:�B��]�R
Aa��3���
�p(�|1���uU�W׵&*hT�3'c9�ц���Y��v��ur�	n\`�]Y��g���� ���c
H)(B�=놙6�H(�Qi����wUD�1��<	ѿ�fS�Tn�K��d�H�� �}��}:��"��~���p��X~�gu�Rޢ�
Ad�e9�p��Xfe�#�����3(���!I�<����f�s��)8�L7�i����$ 7��'¬N��O>�Z�v�������a�aI%!L>��2m��P(�Y���R�w��xh�y�s������ˆ�� ~�- �j2S�]�PВ�
33P�Aa�3(��) �Te9�~ �����2��gM�UP�~m�P1�
Aa����� �*U����!I��Z���0�ˆ����
!�F�
AH.e�~aI'�^~�k9�wavᤂ�P?��$��߮�j���h*�pY��|�O�;�g��t	#�
H)��) ��5��}����/T��{�i ��
@��ZM!I��Ne�II�fXn;H)
*�̢�
AH.�5�
AM�3.g��(��{�u ��/�O|(`���?��j�ڒ��G�8�@�aI%!L>��2m��P(�Y����I̻��TAH4T32�d|	#��7�e��U��ˋ]����w��ln-����88� �&����F�]څYn���S���F�-x�r�i�c9f�/2ik+(L��[�"M��+3Kǻ��<�}|�&UU�}����CBWv���}Sq�G���P�\����i�T�싺�f�NT�n��+��[��Ԭ��K��n��^"�����r��ťy����N,�j�1�M��x���s�W[����t�Թ����ޅj�s7OPYq�����k���xѶ��ҵT�E�7elEy�-YD����グ9����]P���*Q�Cf;�x)uA��G�[�ywu�:Л���j3[�l#G����,���3��kvC���WL�u����f�ݱSj��z�+X�w	������nT�Q�mӎP�cu�(�����;d�a�ӵ�5�xjr��М9�B���3n����^=��b�X�Q�Q��q�����F����Nx����!��F��i��Ũ��
�WK㛷��� ��K���g	����B����(�{[��j}5@S���[ISNX�]^�yȞG;21;�y�{���R�6Y��\�L5f<�b�S�{���WQ��wu��]D��f��67r�����eZ���⃫q[��E�m�ۍ�	��9�c���A�Or��L��/�S�&���˫��-,���t���Sx<�('*�|��U��ǭF;szd{�j��
�7�Fn&���g�@�h��9��y���WP��ueb�IXyC����seV�D=�]c6^�[c,N���ʶ��U�5��j�9{�!�Q�UU�ޟ A�A$ab\C�m��N�ta;ͽ�/-mг'H�:A� �I���6�����4n�y��fq��y^x��2D��!gZ�)N��Ώ1�m7��9yۖE�tG�e:�q��w�Nq{l��R��i��yY��q2�t�9s��dև���e�V��=n�;�@���;e�6���罥{���Rs��G��� ��s�n�ӽ�����^��k�f�Ne�s��C�ۜ��^Y�Gu����:tP���-�v=��9 �N��V���%{i	��8�+y�Bvi����y�������{m���w�}�����A��BHq�">����6��L\�3���a`�Pn�1&���l��a����1ŨKK��y�7,#���q�ev@nH͌J��4`lA�Bb%�[e�������gpL&Ұ�����,rX��h�!��M��\iLlP�6�#HR6�p9�]{J��v������f�#�f�1+
�˥����c�YCL�,Vع���s���/3[jڳ5CA"�ȵ��������jrB.��f���Vl�-�n�h��ʙC&�ؼ�%EoiMU6Dl-�LXQ;\����EF�f�A{F�Fle�M˒�j,n���L[l)�.�J��\��va�Eca�m�
K�Ԍ�@��,�,�G�J���!q@��gUa6�J�s�VbV��A��3KvB�Z�m��،�[��3	��v��íHP��jM�Y�Il{L�-�i��.&� (�����Kf�I\�Y[�L��b��̡5!f���i�GPeLF6Y�
E���in�PE��"e/:�K�ٕ�������H4�ڰ���x�
�!-2*j��;a��)u�fiz�� ��L�.6��#iXr[�-�ev������k���è��3.�
����EpV�c2�1�4���nRUv22�b)�f]Rd����%X6j�n̹l�c� d�l�X�[B:�P 6!H1YpB�k��e����9��M:�Hqit�^�X<�,���J��R��]��E��V��&t6f�ab�r�[完4���JL�-e��m���qF{D��)04�4Vm���49�i�k�a�����J(��&�Ä�p�HhT���lD�$]u�kn��ͱ��a�ZZ�Ý�6�`�:*)������kf��e�p���a,͋�u�A��^��Ԙ���ܴ��tcc��M�j���h#`�6vK.�n0JMc��%��YV����c�v�JLd �4�ЮB�f�0K���5e+�x��B2ꑔ�*E2���d��,��\�΂$u���f��2܃�N�'m�|�j��jh\q�1�C�Q�[��X�\G"�hd3rf���R���G^�Ĥ�T��I��CB���Yq��Z�cA*A��KH��ZhUqwJ�[�AV^�iX@Z!�lue��c�.�Yn�t�0���fn��/!t����("C%n��7rKR�i�p
�ղ�f �m̺h<-��Y��rp��3�{#�����]�a͸�#��#�������붷���4Z�b���ѕ�[��6��+)��M���a_��$�����$P�O=wCI) ��}p�Aa�3(��B�%�2� H��cU{���P1��<	�o�ƒ
C����^U�מ��������R컀��)�{��I ���eH,5RAs.�C
H))
a��2m��P>�~�^�����k��������� ��w�#��ѿ>�W}��w!���4�;�I ���˸
	) ��ˆ����-%}��gkm�[�bAd�S���P4��Xs;a��AH(�- ��\˸
AM S̸i�) �HfQ����Ux��(Nv`U��֧��6�QC�8�qL��
H)��ˆ�62�
�4�Xi ��p5TAH5*�p�Av���-4�I����>���ɏuwC�JH,3�p�AH(�ZAH)̻��}�w}3Z��>�e��U��s��
B���QiB��J�P���7���/��F S���ld���D3�4�R
As.��RAIQ
a��2n2�
e�Xi ��p9���_�}�G�~� ���ᤂ�3�y��{\��.���� RAH/=wCBJH,(���6�R
e��RAd�S�w@��m�����߫_��W��v�'�������(E犌��R��Ke�;\�*���I�:_�zOg�������ZAH)�]�R
Aa��3) �B�i �����{]Ϲ�ew?k�z}$�������M����d�2�
��H,4�\��D��3.H)2�N RAe2S�wH)�����G�h任h�}W�*.��V�ɿ�+xԯ�};2����8P+=O����=KpD�&�'t��F�2�;���V��a��7_�@������
@�h��Ax�@>�����+�'�uTv�����Aa���ô����=E�J!I��֠)4 S̸i�o��������H(R�H,4�]��RAIPB�{޸i�c) �T3,�A`i���]�Ԫ ��fe�i׭��u����_�y����Wy�՗@��E��$S%<˸
II���6�Xn0��-&��R�w@�RAa����H����:��� �	H8Q
H/~���� S�.f�) �Q�4�Xp�{��;�>̬����O����a�aI ���p�&�) �{��}�X}�tz�o�- �6�A}����)�C;��i����-4 RAH.e�	) ���������-&��~�W�G�#���� H��wƪ{s���U|~H,;���v�RU�����$��j�SH�3.f�JH(R�i ��y��5�Z��m}�vYY��.�i��6ĕ�f����;]e���XA�v�4F��O�����t����Sgnd�) �Q�I����wEQ �P�ˆ�����Ok���.���z�O�) �����v�����ߊ��%����%${��6�XlaH}E��ɦS�w@�%$�a��AH(�ZA���������ߛ��d �{��I �g�����Ͻ�w�s���滾��<�^��>aI%!L=�\4ɶRA@��f�M$2�k�2�����ε߾ ��C�ˆ���H�E��) ��)��p4��
33P�Aa���E��ɡ��]�P;����������y�_�K�u��P�8��8�GJ�T75���ks)ٴ(��Z�ݪ��%��me:i�ɛ����Z2"���� <����N<k�܈���O�} ~6G� �g����!I��) ��ˆ�
AC��i ��
H.e� ��ɝ�?�{��~�i�̤��]�4�R
As�p?UR̸m ��Ͻ�:{^�����Yw��{�Z|�I�2S̻���%$���y���������Aaх s�ZM!I ��� ��a�i!U@fQi �2��R̸i�{y����w=�����-<	 'H�'�0}_wJ�ߛ��U�?xrA{۰�) ��.H)�E�H.e�D�E@۟#���u�ʾ�)_Wъ���T���3���,�6�u��V��VW.�4����M��/Z�� _h��
H,���v���%$��P�Aa�� fQi4!I ��p����u�����޴U|~H,;����AH~�q�M�Y{޲�`��H;��Z>�Z��ЁL=�\4͌��P��4�XhRAs.�C
H)(B�fe�L�I�̿k+�޽��� �=�����TAH4T9�m ��7�����φ-�s?x@�$���,�Jy�p4$��§s5��)2�I������~��k����Ad�e:�w@Д�Xgݰ�;H)
�@g�����RAs.�)5)�f\4͌��P�3(�Aa�ՙ�@`��gֵ|�r��=��x��0���X{�i�c) �Wr�$�H.e�UR̸i ��
@̢�
Aeo\����������:�wH)���jH)�Qi8�$J��2����w?g�j�}��7�_��>�������5��%Z�̅/g���9ո�rݫ&�&*A��3:�U�����T--�4���q���fb|������Ι���Q'L�����r�[�S����x{�9��H)�@��\4��JH(P�}F��$2�4
J��p�&�I��4�R
As.�}�^�{��� ��k��m ��9>����l���" �$x<	���.�) ���f����q� fQi4�$Je9�p�=W�{���_<��3�r;mu/F��s��e۰,n� -�p86b:V1v"ʬ�=�t�盢R
�E�(�$���H)��fe�L�%$(C2�$�߻��ھe�N��8�V́��������9�_�����,;��4ɶRA@��ZA`hi ���D��3.H.� fQi �C%9�p4������g=��W��7y��q �z�H)��e>�� H�؞>5S�}�:wBc�x��H;H)
�=E�B��]�R
i�fe�Lú3���8�P��H,40���.�L) ���0���L�e$�- �4�As.�h� �*�p�Ak=�٫r���1�/�Y��nc� �G��ʌ��.�) ��s5�aH�ZM!I ��pD���3,6� �5����N����
��}D) �ߵ�
AM����I ��3(�Aa��{��߳���3����y ���|0�����}�2n2�
���h�������t�A`hi ���B���j��e�i��3(��) ��Js.�) ��fjH,7Re���{�嵦��o�����~H)�����?�"~߷�j�L|0�|��l�!EP�- ���ﵨ
AM�3.f�%$�- �d��1B��A��Jb�(PS�OUQ��N�X�˾�3gT=l���V6=�>ݖ����I��I���@����=<qU��zl�uu]'�)�_,�|�oϷϺ���55�B�
��ch@RS��ڡM1q����#-����5�B����. .�b���d;h�"ҎJ8�˻]�h��ڇe�lk+[� �e�=e�P1��ec`r;:��҅��&-��D])�퐳`��M�&�.���e��f�.�W�V�TMT�z1%�wj2����W@nX���5&�Fd�;6���j�f6��j��&��������c�Z0Җ����6��Zjl�v���.�c1�o��zl��蓠N�w.H)a�Y���R�P- ��C3.H.�s���������/yu��{�ZAH,����o{�w�V����m������XWﻨm ��3(�����L�2�ZAH,32Ðv�R
�3(���R��fw���k��ށԂ�@��\4͌��P�}F��s��>��������C��(>a�����}�2m��P+�f�
AH.e@׹_~���T��G�R~�ᤂ�`Rݢ�@�I����i ����Ci��Re�B�Y*2�ʁh	!������ϋ;�z�wW|���\֋���Xz0��ܠ��\��O�R�%����^C6�i�2��bޡ�+/�m�7�^�JQ����\��@I�/��S��|i�,��6��ipa��A����ݭ�o�I�%����iЪM�Y�UM
�\:���K4en��Kc�\V�f6.��#jXW��O=~}�cv=��9�Q3�kv���O�s\��b����E"H��oW�Uw�W[O^��8��M�vNM��n�^u8�s:nV)uUd��n�@\Vnu.�㢠֩�â��GOֳ����.��l�.�]�}���*�������*�ኮ\7¶7vD�%`��ہ%��y}"F$+�j�{�4�a��A��'���݁������Q�,�zR��Ư۰:��u=ع��	>���9:��[��F���ƾ�|$�D$%9uw��t�g�Ow*=Y�V�wx}Q$����Jn�P��~��+�e6��p���`t]I�yن���̴�]\"��e���������I�}Cs����e�ӵＦ�s����ʟnBq������X�{C�$(�s=ع��ow���PJ˚�������D$BIjK�Ʊ3a��)U=0�o}H�ˁyh��!�B�/MŴYRqQ:xK�|����8Ƅ:�O�w��}�7U*Щf��A�/���g�UVxfվ]߅D&F$_H��7�iD��ah]�������7bB��,k�a��A��y�٪�}6'�ݝ;�>�|$�MJ��Fs�b�}�}�y����u�Pjwznm	#�IW�Fv;��o|֎���5"�����l.0����0m��^STΛR*���e� t@H�K�7�&v��v��wWF�f�^����r����#�#�<�*�u������Ƹ6�o����x����E8�q�n쁻5<��rͬ]]�'���v㠧w���Ⱦ�?�_I�/��V+�}�9$v- ���//�����J�u�t�����Q>
���:��H��"���qI�5��xXN(_.��	�_��{�I�����Q���@��5�����W��|$�XI9��=a?��� a�s叙m��(9|9�ݡ��������ᮌ��裮5 :�
6����ZQ!�f�l4�4�U@���wI,	6ӈ���Y4#[�4*��'>i;؀�I��~Y�6�}��^P�@d�,[A6�L��
�7�VǷ6@��^I���W�=�z���� $�	&L=�mC�tls�Y��L6�A��,r3`n���"%��%������$[^��I?{7�ێ���P����[WWZ�j�I�w�ܣ0)!�5q�4h|�I���]ӆ�հ<76wc�t��{aS���bNc{;k�>4l���q��!q���U��P��p���wb�B�w&��u�'a�Z�y�%�?a�1s�������}�C۟�Ӻy����2�1B��X�iVБ�\�3Vgib�cUͮ�`����V=�ؚZ�72��vy�Sm+Y��eDnQKˮsf!��&p�D�46�3.v-6-��k\ ѭ��,f�X5�7�O4�7��rFW+m�F6� �ݥ�l��[�2��h�GZ�GnK���i`�g#�
�U.���M�Q���P�`ٷ����A����B?�?��L��5c]����
ҥj�狒�[v��*�isePk�YU���7cxn��v��o�>e�x��q#�.C�{2�ݒ\��������i�]
���T�N#��=Y#[�	���!-�Uv^������"�H�݅����N#�̈́�2��Wt�q�Ȅ�K���w��U��r �gk�Ŵ�oT���>�50L���P�s��H��?���
����g���^���(���W�)#4lZ����e�]6�60�˙�������*��f��7R�����A�zLᜤBH����;�4^;ன�t�,�ܤ̚��<���ċ�k���^����1`^V$QXE7����|�R[����˦M�N�7���n���F�cOg���yƤ��,�H��z�4T�?�����g'��2���s����l{uvD`�랷,���?r���������u�}�!�r׍FP)�������;榤�;k@���b�Ċ�h�;ன��}-E�8J�]�Z��ӐF$C�6�s�+�Q[�.�
�i��)�a�=�E"�I���~N�K)�)�A4�k5����+1��0Ү�r��6j�ה��b�����=�7wj{�l�M=�֣(�ᗹ/��D��k�V���e�$BE&��#�����O�	����bJ9�5��(�r�m���9��t�7:@�R)#�I����A�=�ǵ��TR�b�ʫ��IJj���kon�k�Ԛ}�3U��#��[S��])�M�̌ۉ[mZ�-��I)E���r}*�FX����P<�塷S���M��h�U�.�WoT���d�w�f�\t+��KR�,�֑�F���J�t��طE�ͯ���l��q�p�j�Lݣ�ㅗ�Z8i]qh�V���h�\����`�j�dV�����w\%V�g�I/BΫ���Lo]Ʀ7m�7UQQo#.��6����5m�s�ỡ��HJ�|n��)F������U�u�f������Nj�j��ʦ {��\X�x]%h�!R���q���;�X��OL������1S\�{ta[������O���'�]�ܪe���U��ͳ��n��^�����uD�B�ȫ�<��Ҵ<�����7F�w�wb�u��*w�aY���)��G/�����;�q��MAaLsWڭ���A�T)���#�V
̍tA��.��v�u�!�uV�*����5���M���uej�sS�Ys���.Zs�D���P،O��Crr���6�J��pb��̫�<���n��N�-�{�D�؆I����l����u%��5Wd˨�;C�{���f��0���Q"YAmMK�4U^R�걲�v+ڳlξ��֊�3��g�mu��譋����]����MN;�Byu��8�uBY͇N�ʼ���ҁ:^��ocګjU�U�{�(]l����e�,Ԝ��׍�}ĩ�m$�#׶MP4.ƊkX������������"�Z���X�m&){���W�O7N+��3o�_,��H�P�<���^v@�Zgl`Jr9"{v��򽙶G$q9�qIі��%mX�gn&gq�Q�Ԍ��8��ݨ�#��=��W�Fg6���S4� ���S���;km��NG�m�4�Pqs�=�t��2�;��w�����k˽�K���gX�!�A�qIѶ:O�f݇_4�m}�D{��,�:W�Np$���>^�����JJ���qs��v�_,�!�R�+焸���^��\{ZK�\���ip��Obё�a.����<�J���۵$A ��iN�	W���G[X�3�\��#���S�甠/��z/:�6cH�Du�������9K�a�N}����ݡ��")eE�Ds��D �?wwq�u�zv��f�����>�޹{חs�dR!$	�,�Z�V��?zb�wO.��ew����1I�}%K=N��]Ga���~�vƋų<���]�.�ك*d6&P�¹�2妗�WŃP�W 3��G�P���{��]�G_� ��j�y�zy���!�ݑ�ݏW2,>��RuWC�Q/�l�:잝�(����E�z}9	w��hf�"�2N�V__x�#�o��@�e{����L@L�H� $�e�{D�0Gv�ؑm7�o��� ��y���l�37�l�
�&�L��d�3�4��y�&�w��	F�3���:iz�E�XE��
����P�Q�J몼�����_�}�W�\���K����;��5��牼�k���4�{Z��gw���RF$�Ռ$�N9T[��S���&DSc��oB8�,�fM�:�V��Hs�Lb���]���D���RmN�}�V�_pU��w�^��+��~�6 $RF��Ѧ{�o��$_&���z��4;�ó_����,.�c�}�$���ۗb�mKv�F�7m#�4�{u�P:��u}"�I%ȇ�Il���Y%p�y}$u<�ۜU;Ľ�����.�*��JUD&�/�$�$��l�d.�b��>}����bo�X�ٰ7c�wh�P&�CM��ȯ�6}w��S�K����nNrظo�n�1<
�pK,eʹ��)�MUoa��nL���TrZ�{߳���ע��L�CM�,�]lGM�lX�be�@̓ژ���6!Yn�!heH�-��,�,\Eu�0�S6qX����2�����J��(mj�45�"�ۈUۮ��D��s�-pj,�/"Fec��LǬ����lı�]x���s �sI ��R�-m�]�S11J�j�V8V�.���lݘ����˒9�6TY��&�:��*��Yl�ϗ��6�2��e���#Ui�����J2��v�H4��i�.�h̬<�������݁��m����\e��WDm������E"�<e|�ת�����*j�nx2���[�}��	��'æ���%s�D$�F7%	�k9�.��R��:a����#67c�wdn�9Cx��<�w�^�� nǧ�L>3O7�\e���Q�Tݽ��[��l�{�$H������o��_�{��x4���]���3�I�I�Wz�`+���ߑ�79�����A��d��K�Z�eh[�H��[TJ��
j�AUP^x=��?�������Ҷ�t�3fg��q[�8���;�6*�=~���4%���ߕ휧Q��p.j�7�%����T��*�[�����9��5�r�R��M���ns���3�ț�z~ �a����6��b�on8�S��wwk�(���oO��<��MI%I�"��C���}^�	){�Wt�����Ⱦ�H�6�.d�œ`
�%>�ğ|�4���������ֲ�����H��}��Ș}���I6tS�y�2���%̀7vD���<�xx3ݵM�h&�UT��M�3GhB]����Y��5et`3P�8yf�_��~�?��I�?G+w�IO���t��}�6F+�WC]h�)�yl�2!$c�1yז׷H=���ğ}����"f�5�����e,d�R�^o�}�RF$Ry��aNS�n*ٰ�#f�#�q]3ٳfMܛR�%u��P/������F��}Uۦ����*�-]���]�&Ul;pE���Gs�㢞r�q����E$	����:�S�_w!$���l�I{s�]����b�c;���|��I���?3�^T�ܐw����S�]$L� ��͍��6������7ol�hC��*�����ƕ���mML���I�kf.7R��+4C��IM���Ξ�l�� n���1�K�q���Ӕ�Ľuy��{����z�Q]Hd�#�vuO��Scy��%�wK��يHĝ�ѩյw�3T�K�L}L	^�6{��㫒���H��ksov��ݮ[<�+��{/;�۰%si�駜��S�-��������J�7��;SL�����e��{X�gv΋��xAi�������J:��[*ž@��TFe��8�Vz��RUw����mO�j/���$BG�.6��j��X��������)wK���_I$����g�ާ����B{%b}��tz۠Ur��;�����ŻMYe�����n�������<���i.ϒ�j$L�:}bXƶ�!G��u	#E��k�ëK1�_v�o[���Y0O�[ݏn��#���˩�m��n�́�����j4r��Uf�D��"��P��}����H���n)ۋnZP�/9�$@P�M���+��Z\�l���U��b���=��9 $���
��g��Heɾ�>u�K�]���â�dBH���ׅ���L��a�����j����2��M�R�؇���$�ȸ�Wc�o��U!�զ�TlU���+%�a�(�ɚ%5�齖��}��b`�a3��ɶ�B]�u��2�Y�p�j�[��^"��SL�BY�f�f&,:���ixz�p�W&���.���cY�����e�M�-��!�+\^�����F��д�+��LbP�٠"ۣ-�Xh\c0���]6�\�1�lk4��K*�jJ�Ŗ\��,/�e5�j�CL�X[Eu&�Z����gl!M�0Չ*�6b�[�3���_O�f�m�ˡ�V�vq��˘��T�q)�+����(��ĺ&���c�I$����	y��Rkm��^%��bL<�ހ7`n쁻��]mh==BlOt�B�y��һje�M��G�wK��So�Z�����#�D$��bmq�i�a>u��z�0��/�I%���n�]Q��ڦ�yl{ۻ"��m$�G�*5�o�� fNu��5�H��|$_	!�S9|���%r��t)5ǹ�+�s<[9�	�Hso���qwbyuUR4�.��T�v�e��F��J.��9"�)�1m4��P��{۰�>ݍ�Sz�=5ܪ�w���2��̿��$��D$����o���w�s�εY��&����B�LM��<�L�-�]!��Dl�dGX�|��#wWwGNi�G�Q����Y��{��}�xw�>��ci/�}!g
�{}��1��L�w[�����,���W�v@ݼ�����o��/[t����~�v��Ȅ��#�F]<+�y߽�;n|F�Os����V�'SY�۬��wu.�X�@H���$�[~n�mֈ���tt��67�q���Nܵm���wdlBN���ͬ��A�th5I�ئ�#PX�Z(Y��n*kQ�m�E���eV_���W�:=��=�e�g����E44d��7��!��W��w�F$_H����jn�z ]�����vS��S�@�I.Ej#.��w�Ľ�w��"�I�.�������{�a˼�\M�'��G��yO�c%G,�yM���ݾ2��>�n��O�Ӫ
;UJڷ����ɶ숍�SH�t�!󄯴�HOL��}�q}$H��K��m̾�쫞[�#v*�k�_U����<S�[3��9�V}2 =���}���2���+�=$<� �H΍�i�zk�]��`��t_d�XE�����o/��*lAU��҆J�͠��,Ѓ��(��(���H:[�<��ʮ_���<�@	#��)����^�ne�m�(��Í�w*]��c۰7v|7`��B�WdGv�����
���ݽ�i�]��>���D$��6.t�����9 {u���I�[S��������߀�ȾG�D+��r�f��;v���j���7�cU��G���[V� �=�<N�/(��e���u@��6^j/��#�C�2�+D����|Ta.s��g�Ty�+���j-�
u�	q��W������F ��H��.��9�ݥ�{��u\�+�A��JA�N]cp��B��S�DѣM��6���r(;@��4
cfĕ��v�1toU���|����ݏn���S���O�o��;�uQ���Qϯ܏��$\�m��p�w6)��ޣ���vm�xf�$bG��6Aֱ#`K���N@H��	)�ܻ�����·�<]�z�S��7�O�H���"��=����M���w!�yrLGK�We<5�zx�K�b�Q^{��<��}$bD$��m���nj�z=�>ΕYٵ�ᜀ�1"h��T��N+�s/��9E0����A��6ё
;��^Ak�v�i'D.�{O�z�{Oը�i�|��I����΀�^����r�<�	�^¤t���[�m�_U]��A*�U���-�uh�,���)���O�ǩ-�
u�U*:�M��U��z��R|ya��֍��
*�Y{niko%ˊ�S&5,G!�Z&�B��_g˔<O�Q�ԝ]�������m���ɱ<�����	��-�mT�*��ٗ���7����q-�xhp��躪��2.vq���ڬe�5�L���9����v�if��IV��d�q�ɕ�(Nw�g�jL8Kr7b>�,J��wx�w��}]��
�WQ�=��
m�Fu]�ƭ)�ZF�-�X+��d���4W���r�J[f��x�3Ab�Ӑ�an��V��(�1��i�������.��qgUc��P�݈�ݙ�\k.�Β����Na7�%�gb5�����i+�挎�鷔�n��F�ذ�&_U��{;��bԹ�u���yX�]Z�6����-;�-�bee�K��(u�YY�>p�K�̺@���p��?w���?\`ȵ;���Ѝ�0�c���X���9u˺;��n��DB�	��:(���i�ٛGj0c}�w�l�(VSs�l�/�.K��h�ʼ�b��o���T\�1dT�{�6#�%ݝ���_U�ޅ"Q/o�\�S���kb�Ś�2�\�NN�tfI�E�nr7С坷��̦�\L�k�A�RKK?�G2�vH��X��|�������޷��<��9�gl���z��{i.{c���w���Ïm����k�p%�n+S�&k��e�8۬�6�[bW��;5f�lw�ǺI�vZ�{g6��'I:Zul!b�9H� � �J��>�މ.�V��Q;o<�^۸ok��kv����X+-)#e�l#@�������n�=��,��o/��>G޾z���Y�V�s��XЉ�i ��f�JX�.�h�Iaذ�b@� �״^�#�RB��8��nЍ�Q}�/{�E�ӳ�"��y�D��e�^��<C����)��2��f3�D�ްq�hV��AI��u��G���^�҄8�q	2��	(B�0��H�[��/m�k��f[��%�q#��)Yd���y�ڽltYֶ��aeB��On�4ںh��(�TB�i.m!0)rV�\�*��,G+�����k�@,s��-Ɔ�k�]K��#�J�N��g$�ٕՌV1���ݢ�(�0�n��4,:�
�*����STM�G8r��ql4�4.���j�&y�`�XjKq]`h]��RM�2�j���i�AIf���V��Ц�֥Ic�ipR<�k�5�Q��vs*C%�(���\
���n.a���P�1ef�ٚf�)-�@�5	n���l1דL�]�6��R��-0Kc4��lF��Kk�r� q�~�Gͬ��3�c+�f^n����]����Zd̤�uխ��1F����4�oGYvƘs�6.a�)�,Ƭɵ5�o�s<C�WK4)6]���ZZ�ڒ�תk��[1��tö��ec��`J�U]�dWCgfe6K�s�@�xѥ��Ŏ�n�3����F�%v0��81��2��v�0d�6�mBէ&�LI��H-��[M��i`�]6�Kc[(�X;`��U���b�M�pMts)��s3�$�S[���9K��d��rMm١4e.3+��Y���l#)y����\�:m)@�n�ė<��@y��Z���[Q��j�l[�FW�[�*�����)V�Zq���,S%(�R[vB�Pa�Ρb�@٤
k��9b��B�RPݦp���3�.=5��66�ڠ"�K��[i��ں��K+�EtR�h�LD���-�%ns�\1b�[��Xlj1�۴QCjV�ٝ1��H��+��)��X�TU�.��u�ř�o C�J/`&u/8�Pn� �Utٷx ���U��������f�)� ���
�Y���c(͑17g���X�J�lu�u�&��˨V�*&�v"��i7b���E,Ԁ ��U�Hb��d�8�Ce[�:�е�0�΋�n%.��om�7Y�(�f�,4K1c�WP�[��JZ��`BXCLX���5��!-��U\pͶ#�Fjka��A�1��G%�Ŕ�fu��e�ݜ[cĸ�SnK�n�2���A����5qc�,eb�����[���q��׀�!.��e`��\c�R�N`F��KIfb�6DL�.�t&�#	�8�)�{R-�ZDy��5��F�:٩[\4Z2�B�%�km�a|��b�1�;�Ź��t�f]U]\�cZh�%Q�qh��BY�_>_�4�}��M$%x+���)�hS]�ʹ@�8��J�L$DW��VW���φ�z����;��{v]2�*ٹ[�~���E"5��*�&���z1@̀'�I��}�짂	�����왞�^5�(�y�9�"�	%�UXl̙���k2�{k�:Ut;�}:IbD��# Kɺ�geh�����8�s�ث:�}���]�x4N�n��͢�����ۼĈH��E��㩚�g���kb:_j�)�ѭ�`�$I����A�w�r�?U:l�T�"��l$��GF�jmu��b���3,#�b�?'����I 6)[����:�����Ɍ˛[)�{:�BH�_z�g�Qr&�שּׁ�� �Pʍ13j����E��6������ޡ/�ŷ_f����!fFQE�v�Vb�i!Ը[ڝ��h��s*.q�U�}�ث:�;��;��nO�	;����^3�Q���$_	#/��Ps�o�V�.^�8>}�n��'w��D$�H����|]{�@�zP�1S�J���ꮛ��輪�q*G�{��Zb�Ѿ_	�$��)"�����1lpJ�;�f�|�N����T���E�w�[��_�|�TѤ(/���D�<�eZ1�CX]+*l�9���bŴ�K������Oϐ;:F�����:��,����
s�r�e5�|/��� $�V�z��ڍ����m֭����\^:��-�|�$��+��g�{���k��bj�E$rK�+�l�k��ź������c���)o���e��;�W���Y���ݖ��#G�@��y�f]�a>.�9��o#xT��S��:_A�ӹ�3��@��t�2!"G"�~�x�y���ۑ�v%��c����)�я���zmS����P����(I�I��V�J靮#�[xw+�wK��R�e���O!�9�;����g!c��XttZ�1b���)F���Հ�FV� ��K��Wl�n&��
�����	#!Vgp��r�#;����eE�����]W!�$	�A�I��'����E����>}|�QOF�o�{wweV0mu���ޚ������H��^���v���U�7�WYە7+��o�#�|$�Y��`��N/�{�Ϸ`
����n;H�������+�F]N�^��D.�t��Ui���.�|vѨ�b��w�S�X���S՗�����H���X��r*���
I)̴�1;���Ȫ����q�};���������<�t���:{9,��3��t@	�?��I|F69�~m�Q��b:��dp��4��ָ��ƺ�4T��Ԭ�UST��}�~c?I@I�?+t~��u�N%��{�o��q������v7v}���B�;�2J�F8gSq|�g{_^���E!�(�y�B�_��l��vv�+�B�U}.{9Z�/F�o��T���I�#�<Kg�.{ޯ��֣�I}wY�u,���K�sK�:�5�� $��"�D$�������R)r��>��n��Ӻ���t�D$_I.c�M��%����9�b�g��KFuu�Ϣ	ں�c=tՉ�����#��on^:��f�@�X�u��y���1;m.���9H%i KB*)5� �j�R
7U0��M�u�e6e���A�Pu���Gde�B�bZKrc8e[4��2Pqoij��GZ��Ͷh�F�j��Z�.9r�ͨ�f&57\��4���Ѵw#��As
ݡ̦�2ǩr��DM-�����.�1K0Z��=W8��)Hհ #k1fi���V᎕
��bR��E�(cKa5���_�tut��6����#r�]���M4�@�1�H�3�)����i.~�fv���Ժz^5j��1��&�k5�3��g��g��JH�uVYھ�<�h���>�gv���]jۖ��}ȓޣ�|ir����1%vp����p�u��5���tg{[��f��T�7v�vD�'pq�Omp8$�&n�Ⱦ{s{�����R�`���x͝nTvU�SH�]��=$�$H��B��s�@�s�w+4�ם��6[����lbE ���]my�~�b�n�Ɉ��^���`�8�&��ڶ�mk����)�D�ERWŊV�~�C�D$�IVs����g-�i9\z/y��vѺ^��`�ċ��q5�w��|�u��I�U|�x�)͜�۱|�'���GT�Z��s��u�O�q��Q�U$da`�I�H]]g(;r$X!����5U��=w�J��7�`����f��_Q�t�P�~�=���	$��a���{�"3����s'T�o����ٱ�!$}G��1U�O/��};�Vs����8io2#��:ku�M�d����G�!�� $RG'w�za�x��:�KFsY��{���넥��m�cٰ7v@����������~�E����4"Χhճf��*�v���{,ū��i��*�r�?�IBH��2T����d�7-��I�S�'��~�'c�}"�0$Aߩ�]��қb�����Y��/���!�̓��T�67A����o��-���}$r/�ﴄ��ͪŝwb�n:o)�.b�,�d�&�������ɵ�����óf�xma�㕄Y�N�7��Y�ͺ+(aE��w������}��{����BD
�Y]�U弻�i�|��I8�&�vg�'9�o����c�c9}�����H����)��n7����s�Fv��f����#"!$���z�̲��SF�����H���[Q*�GG���5��
��m�5l�ˬ����=@�r�ؕz��|��/ltq*3�z��ب}x����!"�I	{���(�z�:������1ɧ�1�k�Ks��@d��4r���LÞ^�M@H��1&���b��V^�y5g�ّ�����Ⱦ�I�E���rS�s�<�g�@�ש9����`���J�sh��6Jn�T�[�WM����=.{�֓��a�ۻ�����Go���Y�F
�ma��zfIT���vv`�uW�Ny����$BE���$_HJ��d�������3�]����3v}��z���Ͼo��3[��I�U���j�ж��GM�sMyt���T�:�M �*��z!���?�B��n����!<݈��빦��+�mO6���ݱ�գ9OI��̚��î<r{ro?e���ev��dRLĝ�8�=�㴀4����)'Y�Z]X���<�GM���\ͷ���$r/�_I'���t���k��{}r (^su<�Oi	��F_{�On�똛��c�nKE���q�3���W\��C�{���n���`��5 ���φ��ɽ�U�Y���B��r�oY�unUP���`��f�ef�pĖ.ʇ{�|b�n�	Ԭ�-ɺ�[V�D\�cnb�4����a2A�5E'L��F�-�qBY�b3V*�[CX��vv�\�fB�R����c�-��Ml�M�%��*��%%�ewm�Z[�CU�(^�3#7֘k�arͣ��$-�kz�2��m�P�+m����z=��C&,`4֕�Z���:���`C�i�|��b�f����f���8�͛R��t���m�"u�̦�u��*Lɢ}��|�[a4���c���G\Ҏi�,�KnMS�Z)��T��/�t���W�G���9��_�λ�k���.��(���|%m���H��9�}�.��:U-6��G��(^w:�}�[A;܈���#6 ���]ƺd>���_���!$���"Nr2gc�΅�Ξ,�Ak�-��G�bH�BDq�S���o�9}�BH�#��<���w���y�{r��p�ͅ���&F$_	���2�a�7�B緩�{%��r#+��O�cv7w��}�՝&��/Gs�s䑷���A�@��C�f��)�{e���k��G�3K��Õ���I��=������d޿ge�Fθ0\�	鮩Q�瑼�}���E"H��I6��(��^]���^.GA������]�f �{����ޛaU�3�"Y��8a���ј385��yTԆ>�a;�8�f/��b�D���']͵��;����R��xWE��.g^1��)#�w���Z��{��ꇺ�%����E$H��,���]);��7`Nvjw����޸0_o���^ˮ�O��s��!��Ⱦ�����c��U�#������ݧz��;��Ȅ�"X�����{̄�-M�`�KXT���n���h�=��)UM����xҔSEj�	#�H��wS����9uLK+�*�1�{��؇E$bD�U\t�����$;�r�S����]��mpFK`�e;T2�ϱ7�Z�̈	�(�D�yg��ףl���Z�j�ʮ�.
-S��=���gni��Y@װ�g)iXQ�x��hEyx��qӵ�o+�;��idt���]U�AP��sjm�N�>�V��0+��Y;�g)���E�%���#����,t�n��/7��V��ܼ2�"��$����j� �%^̛�^S�g=~y�x)���|.�Fm2�t2��w�i}%޾��,j���%��P�:^�W�f��"�P��˳�*�ۉ�\��� �tv�]�C^eb�]�]�vݾDК�әY��n�<��N���G��Vd�6+�v���Z�M�&5X*�N�ީ��!J�LPܗ�rf��,��@J�טt�����*=o��
��^w�j���v����+9I�Y6,���͊���gU��Cq.�O!y���J��5AY��Vj��|L��:f��W�V:�S|�:C\y�5�s�V_3{�e䖋�R=ټ�ζ6�)N&��eR�ɶD-�t틤y>Cj+�^�}&;�h1�$�R�m�\�.T��aNN�wt�5K����~�+�	��_;reC>J=�|_rIGT��O(��W�յA��<н�{2���Z�z-�}�ͽ}�e�#RR��E�LʮKF�B�TJ��ܠ���RoO_*�5�Y�ЄN����-����:�{�cze�zy�Vt��9��м�73�K8=򒓙K�U�)��[77�0����1^XC.�u����н#���<X�fV����׳'S^��O_��>����m-ĉ��@�(��ۗ��{{��=��+6������:3+;�]�k�_%�vvZ�޽���d�G�o+3����S��jJH:��Md���.�%R�D�"t�m�
u�6㬼�[fv�nӋ2I���,#ʷ�e|�2m�yVvy֞��w�t���}����|N�medq�m�6�4ӣ+0�;}���lA��w�����+�.���Ȭʃ�w��{_8���˴��=�.N�)�����{u��y�V�yў�m�^�E�gz��j���9�9��y�tU���y��J����6
�{�l���m.��ge�zoyםE���u�j9��W�On��ȭ.��GE�v^Y���qg�=�wb�H�����?��?���Ș�`H����Y�0�VA���`H��������?Vrꘕe�	�A� ܚ��o+~q` ��	-��?�2?�Ds�Z6�`?sa���7���3�g\ � ���0$V~21�#s^����h��#>JqD:f��fHY�`��nv&����,#Xగ�͎R9Pk����G��w6)�	��ڦ��5��pfV�Y}�2���L~0$V&D���y[l`!�I�Ȑ,f>�<�:�;܈����A͑ ��M����t%65�#|�tA�A�G�E�G���F��%�|�:���l�u�������"g�#�"d{��ն�,(�)�A����șȃ����}��Q�M+>k��W@�!����'����G,�K������B/,-�O]Q1�b˹q�����]
��E�l�u��v.�wh�l�������۫a�k
�� f���0D����@��D�)�k8d$����2D�C�p��Uc�y��-{�yA�#�E@2 ��j���k�|2V��a
4�[h�*�0Bj���G�s���M�f[2�s�mZ��X�O����/τ��3"dH�\{��V�������=�姌�qG�� ���X>#vD� ��2+�ף���m/�� �p��+��5��V|�������>�"�����®�`n���g/����'���=X��ʾ6)z+}��U������A3�22/�VA�ȃ ��hu;|��;��ܙF\�N��om�u�����y�LE�of �p?tA� �"�#�dX�7�n*��p��Ov�X�-�� ��$�#E`��خ�V��vKf����/<�S�=7����+,}��I�J��1�f�k����Ƭ�Į��K��nk��(6Q��b�M*
�-���;k�vqø ͆�,��n�v���XV�Pݖ�%�s�d��A٭cG4#qvu(�*A��3K�SJ�c�Ga]ՠ�+.�]�:�ä�*8�h��5���v�R�i���ot��]� #��P.
�m(��L.2k�MU��)ܷa(�q�n�BΔ�����B��.E jd��!Q�X�b8.JZ:�e���{�aM��\�a]�&M.��1�`��vf&Z�3��I�U�|k����a�$L�D�;�˜���t]��U����&�^B�q���O�	�%�L�0F�]׳�Ϫٷ���Gt�{\���on'�����{��#"k�9�'���膞���j��+ ����'��Yܔ})'\qjb���|���W@�@ݟHv>�"D�v�l��eN���8���?X��,����t]��U�� �g�d:�������T[vg}t���"F ȃ ��fDs���X~�﫽�u����ʂ����0A�#��#{��Z���#z� ��Ȫ��3�0í���=�7L$&��\ƌ��3/�����z�f�<�E�2!s��t�«9��?tB�]��*�Rf?��L��D�	�2�K=�}�!x����B����x]ثw{��`7�B^�����k'9��Ӱ_fv)���W��o��.JyQ�>��3nsiҷa���[s#�q �:���n���{/3"*�8��@��2.��T=���D3P`��?��2��dL��0��K�L���j��]���򐱡lp>n$͑>#b`�da�mj?n��f�h@7���'v��Bѭ��T�R�>{�]H���L�'}�h!�Mlz@["@"D� �"D-V�5�w��a�ܞy޻��t��Ī�x�<����L�f)~>ҷ�nK��b��J�I�l�3F�mk��]�6�5��
�"X�L�ږ��7�?�+ �#��ms�����V�l^ ��_g�{ZVA�a�&��F�0ADU���ggĔ4�&A�]�}!�Ox�t{����� �H��U��þ����k����0ȑ3�F:���as�����A�]ѓF,y��kn��F	��$�h�7�E��Ɏ��LN�:]1z��u�k��W�V]E��͋��P��vd{�n���vf%Wk��g�`~��2&?`��іW/9�!��3�&�&�u*�Wۙ��!cB��	n$��Q͸+o�`�F���Ma�"L�0A�H�2'�X���?&��;�?���{��{)e=���$nϤ������V�r%Q+���D�`U@	��t3vSu�S763UѸԀm��.\���c�<���d��"D��F,^{����{:gfbUv�~�|o����@8��\A2 �"G��DHQ��t%{^G�� �_o@�T^�=*�s9[�,h[��O�dI*��=y��V���)�}��@0$a�dLA���,������}4�Ut{�G�w�D��dO�0�&�>t*��ϒz�i#�5D���ȱy�o���ǘ�2"�㏷�H"��C~�Wv��K/(�m�pu֡/���G[��&K2*�,��.��J�`ɹ�*���n�pItC\�ήQ���&g���md� �ȶ�����0Ab�D�0dA���w��UUld�ƽ��W��ʝ!b���{W��0�?������9�ߦ��yo�!���L&4AtY�Z�A���Q�Q�q
Je&�Gh��?{'�,��dL��1v`�'�}����r��>�컓:eՍ�#��`�S��$a�$L�O�e7�r�<�����jX��<���{:e�cUv�&y�da�"��U��B'|�opx� �##����� �ǹ\>�N��az�d�m�e��HXв8���H �f�+?`ș���9��r��	��WD���볣�K˦^ʵQ����=k�Ra���8�y�3�H"D��/��2$VWIv�H�r ��a���z����*����3�0AfD� ȅfyqp�y�+j���r�;,T[�.��Uee�Ws��yUA�SF�ۧ��Z��FCt���x8���h^e<�3)w���UѦ��Wfӛ�i�X9��[�gK�ݶkBnɋ��k0LL��ܧ�<����ҘU�[�G(��u���l����ct���1������GX9��`Ɯ��Qad�],j+�	mkh�V�r��@����ڒ����%8��6�U�g1j��Ss^��ZnD)ih���B��8([��@�E�w.�Y��e���V�����6X��Kڹ�n5ô�6ШD���R�QfY�U9ֱ�OP������{����Yg�"EF�F7��+�:Bƅ����NX�z���K�L���`�D�?���L�?�{��*����,�`�r ��3�Cý�O���_t�� �#��dH/oh�lDO�0/��OD��#E`����s����I�SqH��{�wݏe_cuv� � �9fD� �#q����ч�2�����F&�y!�;+��Bƅq� ��O��l��i�pd\O������Ȁr0�2*[�*f�Q���C!���'���/�{��yA����?� H��W�~m�~�7�\W�Fgf��5i��v��Jՙ[7.m3آ�@���m/gG:��|������ȑ3�0��9�Y���{;&_buv�CF�^ge�fl� /�3<�`ȃ��fD#�w��+�+���"#.���o���Q;l`�
[��5X��]1t7Dڡ�S�W�C��.�D��[T$�ڬg63Ҹ3Vhݿ�g/��bjHN����n���\q��l�H��u�� ]0�7ɐL����?����[�0��e��wvk�j��O�T��D<w�`"��dL""`�]����V�]V, �a�;S��ݑ7g�������EU�q�@�~>�z��ha����� ď��Z��%7ίD��!rs�+���b��A���da�"g�$c�m��s���_Xťo�����B��$�αeGl��*F���ɱ�L%�C������?��_?>�0̉�	�.��^�|�.���0�
�*W��x�k�>7���c� f*��T�^΍�JbFtI��"E�����W���r�U����,�Vux��U�/��0G���2�?��|����M(��uuK{�W{ޯ]0`ko�E�)˪7L6+�q�+��aC�	�[@���mD��3�sp[��]��̜��Js\�W��B�q� ���ȃH�?H�2/����.ǻ��<� <3X`��;�:(�ws�{/G����O�'#^������|�0ȑ0~�|�a�D��NZ+�3�|��=}"wr�����m�����A3�2G��Ⱦ�1��~��^��.��]����k��R��⸲���Wm�3M&��R\����/��,������7`Q尲]�s�jP��\p"�2mZ�z��1�_v!c�2&~�}"D!
o�^����0A>��Ί.�r}f����#㼃�3"�_1�{2����ޭ��z��Zs�q��,f�wJ�����K�ɝ���}�g�d�0dL�"�`���vfY��0}�>�{c�7dO��l�����Z�,`W�-D�{mKѣ.�H�n�z�aK�	��s���	�ڋ���j�U��'��ca�(�	[i�v�]��k��Hff�K.�3#G�8䜥Ub`u/��0̉�A2 ȑdZ}z.�yw]6�.��!0nI��{S�w�O��� �#��"`dc5��鶕�/4��I���	��5�s��Ů����6�5��T�ړ$�����/K������6y��"F���`�z�+�&v+���Bh��T��+�ĐP�"�A�#��������J�F��kS �#�תl^���{^�6ׁ��9`"μ���AxqUJ����`�����H��Y����W�T���>="\=ݩκ���;�$3"���"E�^���7���\20;�����]����i��<�����A�6(�����O�&r�`D��dUFU��x���S�<�����ֶu�ף��=��r0�&~21� ��F�޸S����^h<\jn�Er��U4��Jua�Xj)e���J�[w�Zn�P�̦�k�}�%SƆ�w����0�[�FcS�k��R��dj��h�D�r+ُ���nt�ub��7��2�l˸y��8�������@�x6Pß)�S�{�����Ò���*.�M�m�]���KB!P,�(�Ί;�M���F#lH\W�w$�a��4���I�ݘ3dU�����:3ZޫR��L�r�M��\�u���Qt��E�����:�S�{�3ڶ1�C�5��%䬮����$�H0ME��:�����C����?��sY���y[���[ZZy�/T�`o���f�M(��n��8���rpSf`�V$�YH'��wd}7��D��\k6��i(�Ul�t�w,m+���Ud�f���������l��C��fj�Ct>�bٽ}EVohRS���me`]�;7h�r�Ɋ�8:�ià��W��[��`�����!ʥ��Z�2��l��Ol�{k�@�vZy��ͮ�a�&5MZR�Ԧ*7�{���:xe��A_]*�|�Zct�Z�͌��ɼ/��̃fT'�P\���[9s��]�U����Io�Բ���yhcsr��_Vc���>{�^x��(���Z���L�s�t;�b��i�;	���yb��SlQ�pc��!�)�MQG���YkK2B7yY�UD.4Tμ��l!W�5�_^�٭�
x�N��"L���p�l���ƪγx��7��7u�5yus�'kc��d;���5Zt�%�["N HU;����j-�az[+��۫{rm���ݵ��:�˴��ݝg���ʲOJ���+:٬�"��n�����g=��+â��]�u��wi�Y)t����{їyu�m��y���[4�K�,��{e�eK=�.����sl����׶���g9z�𳹵�y6)mYy=��^y�e�(���vw��Y7��6��DQKj-{^����RyY���jv���ͫ*�f��8���l²���z�ge�����Oj�j���ݙ�2�6أ������v�1����=��Y�g����D��g[-�X���-l+Z�m$u8�V��mgG����m�o;����C�g	e@���d����֊��{Z��#;�f�<�/.{޴��'v���ݫ�% ^�߽�&0��]D�f�ԍ�	��G*G��C6�u"�'-c��ݛ�M�s�6-XM�Ў��y��P."�m!�V\�X[U����Wc�3r�b�7�z�T&&�	���)f������o[Ch9��*J�l� ʶ[(�26i�-�5؅�� ��E�	�kl���iIj��0Ih�JWVf��Qh�ƪ�B���bMc�u��r%��[6��u�!Ƙ��F�-�jD���	�DnΪV�j̉��(]"���i6l�7MQ��jCDSf�GC6Z�JiY�&Yn�.�8��ZF�m6Ẑ����"A&-���k�G^1j��rM�<K�Ҍ�^M�HZl.-����J�0�Exin�0��c�˲`M���+��p8�[W;r#Q��ćU�LU!ZhJBh�Z�K[Z�n�tsG;L�p�%`�o5���`�j��ql�6b�LMx�5Qf�M�nlL�u��5�VśK��m08���1�g]J+u�fʄ�0�S&��)f�e�MS`�\�ao;FӛqT�	��c
Wh�`��Yn䠤s+��M1�2�1L3F���]�u����4J��Sa��Wk����Uk5���SMeveL�Z��qe�X��k(Ib�LX�40E��,��Ci!mMM���b�;Ɣ����,H�]�F�Bg�PUզ�Yan,
���kcfZjr[��RZec�PK��gk+T׭D�.Va��fN��%ʋ�{d��95�W�]ZeЄ��3,�]˖� �ic���b�Q��:���q<���.����D���-�f�����X1�dL�尙����R���s��\␴P��ɩ�!	���!�6E�{����,Curf �#3t�Ir�6�feңUm&n��Q�Z���78�X�[���햖$���`EB��q�1z��°��K�-��nn�lj��q]��Gmt3-��14ezЃrBke�@0�s��6�)�����H�]��
�ѣ��ee٫�Yy�l�<Te,�T���k.W8�rM�eՉ�A�K	3GL<�H�WdA�y�Pt�,v��֜�9��%�CZ�X�� �Xɉ��(�G5��R�KՍ-7GP������Ԏ�ũn
�д���[im����N6n�3*�Z\�hSL@�ڱM2/$F�I����R3m�	q]a�)B�.(�jM�r�̜�ߟ~��L�MF�`�̘�[��Ȳ����YTq�(��Զlљf�/��1	�֛�"��dAޜ�
���Mͮ꿺x+/ծ�	SA�~B���`w+dH�?H��_�F�U�WP��L�g0��s��W�uɝ���x�y�2*���kb#A��V62 ��dL"k	ñ���v,�k}ˍ�z�kу���j�"�&�/�_k;�:ք�9$3�۬0w�"_�'���fqSu~{�)�k[�vk�w��y�"�A2&D�?��{��6}�W�FH�q˱���S�ד�wA;�$����0�![j��vu���UUU!{M1�Y)��m��4u. m�;RX8����Q,:��	�A�s�+ �íz�a�����`�-{�;U�*��XA�27S?#�E`�"�P�>^�a_k;������Q�2���b���ڇ:�S���q����݉��[��^%��ڊ���0C�uq��(�N(�셣zK�Q����ޟ'AH��xｹ�G��#<� �jdH�H�?�`��"��7}H�����WL��.�{�������?�&D!O=��oD(�:?�r@���P�z�oIjP��n8Aj=�a���/,���F�Ș �"�#ș�*�]T��t��Y�9��O�T���Ӑ"�� �#��w'�����a�Phh�1%��hmWU�k�b�b7G�آ಺�Ϋ@�N�S�Ƶ��v&A�9�� �bn�t�/��j�漜���:q�&��z)������L�@Il��3��p]�n�Q�mǐ͑5���ozKR�q����dH#vgv9��U����<�D�Y�0A�Ȇ���vd�EBKz�"$�\��wp`�4�gw4�z��c�e����/�����ؽ�k�Mב[6f{`��.�}p���l�cq%�˗A9-0T��|��������}"�?�-��:6�u�Ks�ǽ�Q���#�b�U�w�ꎺd�ywK�g�C���V3㶘 �f�ȑ�L�#��"�~G�D,����Gd�;��]��C	k�ڟ�dA�"`����j�R����n�;@�vܳRV��1�\f9�T��X�b!6��ƆҴ�I�w���~���n�'���0A2 ��-�y����ǽ�>��	f�[�Q��6RA�?��`�$`H��D��Q\+�� �����b�畏w�ꎺ,��ꗁ�fEp���i�A�VD;�0�a��؃��dL�$cI�x)�j��x���ݜ�M����	�_?�0�&~"F�?��|,����z���* ��0~��S��l��
17;�w���<�)զqzOb@֫��w\�@p}�i���]"qC�ꚕ��0�癰�ث��nzr�D]�T�ʚܴ�P����_{ц�0A�ȟ�dH�
�yW �=S����wul���q�T��g�d�?���A2 �v�E������g��}�E�u3vU�hL�ꠠ�A����[f7Ze�cfE�ږ'�ϰ����`ș �{uf������P`���*�qE�o#8��A�ڀ�}"��2;tqy�UG��,a�� ��;�S��R�L(����	��nϤ�K�*���W�������F"D����P�{��7�Pݛꎸ̜���� �����X �"�f�>J��*�4�������۪��~������=��7"�E��H��8�3�?�_X2 �F2.Q��ذ\�8oN�Ƌ�0��s�{�&r�#�� �#�;ٜ{}��t�4"�sz���zvr��/,�@��x���覜=����k�
�5��U�o���xw3c>�0�ݬ��\	�f���ߘ���#3G��.�,áZ�l[X9!�3M4n��ɉn�F��MBYךL�Ԙå��	N
�˵sp��cu�u�I��wJJ�#�(��#D9�Xi{Z�cm&��mHb�:b\��%4]ъ��3<]f˅��(���`b�Jeu���E�4w��I���6T��⮛L�+�лY����GXX�VZMn� �ـ����\��n���'�ײ�)KT32�b	k
�l�f�l���U��`L�3C����~���"D��D�y�ǽ��E|fNYUK���J��c���?���dH�ȃ]C^O ��{dH�IF ��j]-%/~=��FDH��D��a��K��z ��"��?"GՊ��wp�)�ƹ�}mi��s��<��șH�"D��5;}^���A�7�?#X����/C|fN�UK��!x#Y��,܎<t4|�fD"F&D $Z��c�,�F0���C}�K����A=���dC�E��a�}���v���!�d�M��K08�B�]V h�D��s���jh�iT�(�Ef�p �?>�3"`A��ׂ�w\�6���\'�ӴG��P�i�D�y0A0��&E��jV,��!:��(���jX�$�P�"P�L\�n�у�X��b4;=N��;|d�vG��U;ijG�)��{70��kK|�:�8c�+�]�5�Yɏ%}b�Ň�{���s��R�>?1#ȫ}W��ͧ�PF�������0A��2&D�4nK�T]Gt�m4a�C�#�Q���"��H��X#���V8F�&���`z0��g�ab��V*������k��\	�m��xΟ;�0܉ �;0�E�D3��p�����;|��yvx`�s��R�?a�~0̉��|Mﴟ?r�x�?P�H�G�
M�m��i`�����%-q24���52�ܿ�t����1�0A0�kչ�M���r�h��쮳�7�>� q먇9s������Gٮ�8c�Ո�q��*ⳙ=�M�y��(�vr�J�8g�`�6�@�}ɂ�0D1��H$aj�}�=N�&ɹ%�'�R��Y^���}�Kԩ�.���)&߳%��t�Byl�Mm�+�7��
�4{)0�a������;U/~9�X�s�\yʸ�����uՏ�x�V(͢z �1H��;�)hod�5�T��Tp ��O�P��0+D��dL�Vfe��b/9E�s�9��bɦ��0�j�쫌�d��79�Aj�+>]�9���~/7�Ͽ���ei�9ݴ]i�W��ʰ%{V�,r7-V�.M=����W��zbz�Y���/9_���x`���xqo[5�o��Gڣ���[�U�r���X`�"/%hsPM����>�-2ؤS�����k\�C���j=9�$��Q�~ڵ� o���A��A�D�0d_3"�^]��g�s'�߆[�^�79�H P$�7g��zF�H��W,�u������� O0��|F�/_>����&�����2=U�g�.���=/��n��K���]E˗�u�LTmЬ}x�Ɗ��u�U�Z��4[��ۆT7��ǹD�0dA�d3"�Y+{�V���D�r��-��7�T��T{���d`H��CʨX��
�1��1�lM6(�c�%����ny�lM��	v�f�U|�&�� ���0&D/�`�l��&�<�	K,�	iX�p��z����r`@��D��~2&D�}�{������vȑxq�s�=�/nv;�^s�0A���4�<R�қP;V_�@�G��Y۲�Y�J12��-K���Y�n?i��^�K�ھc#Eg�#�Edy1��c׾G��@m��"d"^�w�q��&�<�T	#{bP�m��3[��'�"D!�4[��ʝ�fX����9��pZ�y7U�G���"s�[�U�����'���u��yc�*�d�3J�|��Q�{��e�AZZ�תu�i����t\�se��J�0�־zT{��m�wZ�������ogx{���r�cu��p�6��k\�Y�1-kM� �6�E[��2=*��F�ݰ膵��Xİ35�k�pЖ-9��H���&-�]����";-˹�H0jX3�maZlF����.��a.���Y��������,֗gmT��Vib�+��1-1��3�ֻ70du{���P�ְ�8��qnvu]��R>F�����~o��Yy����j(�L��h38�ʺY��SmU+�UI��TF$?�� ����"��#�Ң��<�:0*���o:ѩic���?H�2& Ȁ�t=���M�*�c�������o��d���5�	�A��;�}��%K
��n&A2/��0D�$a�e׷�J���+��jP}��ۊ�A9�$�$a��ȃ#c]�����z�ŷ��� ���`�L�#����}|�6�ҝG	j<pd��ӻLI@R��c�"�$a���� 5�H�csb�w��79�����A˖9V�9c$��}�G����"x�[���,F6Բ�J�*��
�ԕ�a���%�X|� ���������ݷ�z/omS<��rff�w��YاR�j`��0D��"��
�ELh��7��vz��.�����ЉT���a^�%Bȋ�aݨ;�9��{R���Ѵ����u���%r�t/K܆wZںW;�{����ȑB;���])сTp>i22 �!�n�z��}jJ�]����?{�d#șȆ�^�T�v}a��E������5��@ �ϧ�ș�`�x�k��v�Ӻ|�A��#bg�����o�z/o{� /�q-��bUZ�8�A ��7lH �� ���|=��G���͆8,�3W��������A=��~���r1��T�D���^�T��A4C��f���k�T \��Cr;��&�`&��O��A;`���2&A�ȃ�s5L��;�M�s�@�֮�]��ٸ���'�#���F�b?-�0�p�A�{"�#�u���I�]Tq��A��"�	�]w�US�P�E�`��A���̉�D�W�y^/u���^?z���B�\R;�2�G�q��cF�5-�[��"&��9q	�e�A뼳��u��y��!f`�_b�i;2��vZX�^ˠ�|Z��t�Nrx1bN�/�`���\6��EfժH���76�+�{9+��2����c��U��D�N��U�!��G�^f�Ƨ+(��o`�[&�]�ɗ�����62���wle��;���n��ii�3�h��B��tf�F�V%�
�S�Ktc*�N�%�˄dѻ����7;���b�=�llY.޻W�:m��F�m�e��X-�E+˄rͳ/8e��Y[�9��R�r
E�)l�W-U�J�5��&YS��R�N�T��#BAa�J)��ci	h�}ٶ屚nv7�+���8X/$���:2��V[�Y�%5.J}.�vdx+,�-���U�fG��Uҭ<5.�;���vi:V�	;�ٛu]�%��!�(�-q�Ks��o7_d��S�%q�b���;WUl�2�3:��nk6ļnc��N�!y��M��ũx�L�T\�uG��l���,�U��j��hT5ui��Q��'�F����e�9V��eԓ,��)��v��V�<�I&��Ud��V\�	�4kvcΎ�33rl/��Ƙ�23Vu`ئ���ZX����n���3�A]}wH�v.b�xx��U�-�\����gʧ�3#�Y��$�{��`X�Tħ��Z��,LB�v[�Qz]e��AP����xp'j�g,e]Z�-��{�9��r���f��P�˫�U�R���oh�=��y^^�e��Ѵu�gY6��z����,�f�0��ΰ����kl�:#m[l�ȣ���cj7��4�Ҳ-���gg��e�����G2(ѭKb��)y�N���������j��{oNH=�{mm�p��Ĵ�㳶�'i�6�姲5����4˝�ض�l9��׋��X�7�H@�C����M���4��ܴs�����y��'i�w�w�����ֳ��&Q6���v���M��&nn׶�Ɣ���Ή�u�hq�p�{[�͵�y�q�ne�.����z�m�5�f��o<�c5�I6��^���ٽ�h'mgYn[F�{��ek����c���.w���ݭ�����=�U퍘���R������=�N⼭��nN-�oL�CX�̰�$mj:̴��<�{k
�-�w�b;-��~?�օjXW�����;��D�sdI� ��#�E��Q��r�
��|A ȃ���R��pm�\$(B��r�O��}f�0A�0�H� � ��#v������������ུ���� ����D� ��B���w�����}�Ľ�ԉ8�b�Zm-c�%�R[�� �&F����V}���}�f!?>���D�20�{�4u���ήp`�^?f��-Gm:/�n0:+?#��v �ꫩf\����s�H'z�ò(�w�.=ݧ>����G�2*��YMn�������;���2$L����V�7A�s��{��%�GwK��y ����0A2 ȑ3�o��?c�HX"j��y?�21C��z.��9сTw�%��F:�V�r�C©gN��^��ichw�=�ߥ�C�9.ڱ\v���na�t��*���˩�81j�o�Y�,B�f��U@����4��#n������)㺙Ȁr0��{4�̴�e���A�`�~�|{��ݾ�� ��fE�1��p��組	T4E�ڼjڨ�WT+e�˔���Է\��Ü�ɧ�}q�ؾ`f�ȑ0� �����W�����/��T�0\Whx~���}`ȃ�#`�`�����%n�R@n�r&��S�:}F�];�aTp ��I�#��no��^��q��&A܃"D�D�ȃD��=^�v_�s2���5�8�Iٳ�;����26Q��3��VA�m��ɟ��0��B���>�6�ٻ��Nt	��]�0]���  �#"����-���4��U��w��8u{Ԯ�u�6׈'�|�0$@\�w�������N������_Z�(ޮ��{}��3M|�f?d�:�*��3�m��=�Q�Ki�.+��t��\#)������:�����"��+�*�]&��M��lޣ�Z��y�Y�Z]�+vxJfC4��ݢ�m׊P��\�%�6�f���)WQNn ]�2��t�*��V�Z��R�ŦaK@0Z(\$�v�r���#`k-�7+֖��+���۫�h��^�Wk׮���j�;T&M	�R��L�2�#b�	v����sl�mie-�:�6��8*���=�c��<��[[v���K�趸`���KkQ�bM�)�3Z�,�y��}���1r$�Đ|�	��8�������w�u^I$K�+��2/��L�#�?H�J�[z�\� Ȱ�@�ü�w�oü7���ׁ��#"Ēf��X��3}\��G��	� � ���"`"�O��$��=^�W3z�k��S ��	�~20��0Ch�?r��w �"����A;�%���'x>2���5ޟb�۬���o����y|���"`�dLda��S�n���^�"Cy�k�x>�Ί�׈'<�H�2&A2 v��k��������ڙ}Gh�j�A�-6�n�4A��H��Q��mU++�Q�B�����՘����"dH���j��z��޻����g�tfҝ�* ��?H��}d7�7�ХK'�CU���k��0��y�D����52j���t�n��r�'�iH�����l�f�5Zw`Ŏ�f#d�о����)�C����L�.�ÿ5�	�Ad3"��/<�E�Sգ��L�A��_H��D���B��b��u��<̧���gEwk���D,"`�dA�$lK��n�~�g����㼟�����F!��j��с\p>j=�z�r���Fbg�3_�+?H���$a�d[VŪ��Q�A�_ݭo�������o�?�d@H�dbg�z�����~y�-�B`v�&H�6�A��e�0퉜X�Z�tbd��.cm7.���Yo���Y?F��� ���{��:��\��Wv��\b/w�y�/^b�C�#���0A2 �"F�2 �#�q�#%@_�s�Mat�u�j��с\q�9�$"�,��u�o��`��؃ ���Y����ˑ���3>�1��-[m�ɋ��4q>iE�v\�r�8�W��<9�v�y�Pa#��ɳ�D���Tzyҙ�Ù*�����4ݹe�~n����G�2/���D�����$�i�t$T�#9GD��Fכ�S��
�cȻ��	΁ �l��0��V�z�W�\2>��H�2 �H�fD��=7Hع-��r3J�C��E�'w����#"�?�ar���8��Dt�P1f�@ɓ8�lv��������k#��P���&�J��^Z>?z ���E� �|��b�LMs�,����F���wP�޻Z�t������#"g�"�=����EH�F�H>!t�ǳK�zTkz�b����y Č0dXϴ������bf��H�`Ⱦ����lCf��e�®��n�F��>j=9� �?�VF�������Hw��+��ǯ�v��Mۉ�v��_xH&j.��|ׅ�7=K�sX�(�dIB�j�'�ך�>��6(��f'�v�yP�.���A�X�܄�ծ�zU�
�r�F�O&�Z���j#��22 �"�@�"d�a�D2�HW�y}�/�FH��S}�1|�
���]\p�<}>���2&~�^�����M���S��,"V��������R]��B���S6����l5�uT,(���̉�da�õ��:���`G;��!�\Dy\ ���?���A��x��ޱ�؟��FC����q5�ܲÿk���'ء�E���.VvVo��X�0G���r`��0D1���m]	�b��]~�y�]ÅWnv+�_x>,��|a���]���W�G�D�y��m�Yz��J13]�oq�����,�5aD������6~c�ȟ�����0dP���ų/�dϻ/1��n�9E�~�����d0d_9�U���+)�-5ܞ{�&2�I���F�`�x���Υ<�f]a:&*�AI�@;�1�N*�/+Nt�9٨vh���cO'Q�ƃUC-T��L��F� v�Q��hiFa��:ZRcV�°p���gm1/`���`YE���!��Z`�P���f]��&��4��`�
�Kv*,-���c�hKSc%T�tV8�&����暎8s�C���^Mn���`Vռ[
��ؓl��f�ms)T�v��-����X]���V4�ю�
�ɐmŃ��\�e
�f6�t�H�����5�u����xյf\77u��]3.�[v��g ��
UI�k�����!b�mu\+�¥�yWCi��[�#T�����2 ȑ��A�-gU���Ƕ�̾��!(a�Q�����Ӳ���}�ژ �a�!��V���׽~��}�c���|YG�� ���
���r��{u��k��+��j�P�"��20Ȇ5����>��M���r.�x���f����,T��"��'!�4��P�O�FN�d#`�`�!��"Q�s.�A�ww��i�ǯ)���O�9��C�F1�=^����E޲��]�C-���G2����4aH��M`�[5&k��_c^��p����A��az�:wQ��]e�a_��;���6��4��t2���0�2&�D��ذ�>x���ob��6/��g5��T(,��ѽ��Y`����j�������\O+��nҜ��7w>�Z���7�G�9�f�u��,T��"�㏰�$��a��ߥ�TЁ�����9��(~�X �Ƶ�9�����r7��u�3� Ojd���5�0��}+r��^<*f�x�����L0��Λ���Qi�����A�H���M��w�&20�& Ma�D1�2'�F�i�Ԧ�ư��Nz<ԉ{�/+��¡�g.�;�p�$���X ��K�+V{�|�=�Zp:L5H1H&M�����\��m-FZuƩ��i���i]?/�Ѓ���̋��1XgYɾ���4#� H�̪����d3$O�Eȏ#șa���DDܯ
�á�Y%�]����,���8;~��A�� 01B�Dv��HT�x4sa�G��A��D0�Čz)&��^�x磡�;ɭ�����Ofe	[8���[h�r�W��䡪�j�ܼ�W��H�z��\�SɎ�0��V,粥���iv����~�ł�fE�Y!z�@�En��Z����AXgYɽ�"}3��L���}c�S��tpV(�8��cș�a��A0����b;��&@���9�y���aK�w��A��O�+���>�aT�u����ߥr����hk��mk5�5�9�E��C
�����cm4k��o����Ͼ���x�vD��l��ep�5c9uq�*t7�Ù��-]Q����wɂ	�D�?�A���9e��{��a�ya�Ċî���æ^c�At� ���D0i��:�<�r�g�?�:X �fD� �ԯpy[�]���m��r�+��3ı�;E����<�o@��'U>Rr�Θ�(� ʸ�IP�J]ދ��X�]\q��fA ��C(!�^�uF�n�*�jgL��з5�
޻�����,���.����j��F\�G���s�v�!=�W�	����F@!%>JG�)���sW0��;�d�{"�y�A3�S�uH���G��J�����U����6�
^�$D�n���l9(5��a��ŕ�V��M*j���OX�У��`��-^jng+�jX9~��n�.s����9�,�.� ��U�IMf��w"�T�Q��1u
�K�B��m�g2�8afAbU�zz�#;�D��FH��'A(G�)��s�f��F�u�,�dF�w����������
(�)є�.�4X ���(��IE�u8s��t7,�jr8x�@"���+%+]�ϛS����O�EO��)�BP+=�Zi�������G��l�ٷuK��t��F�Z#Ǐ�BB��rBB��2@!&�@�@���BB�䄄	'�$$ I?̐��$�Ԑ��$�D��	'����	'�$��	'�$��	'��$��$�$$ I?BBB��I	O�$$ I?Đ��$�2BB��I	O萐�$�!!I���e5���@ ϥ�!�?���}���� ���p���>9�W��t{�Lm��P��P(��M    O�R���A�CM�h�@�`&F F&&	�bi�?̪M$�  4     ��h�l��G�<���d=!�A�F��L�A #j�)��A�Em�"���H�\g|�	�@�( O��ahD�������|�wh���7�P��A0
,J �? �-"��-Ej*��'?fj��~�/?O��r(��A�Ry�����C��P�׭�������a3_���;���ZJ�kٯGkVkz�kd�	ʄi�c˺$g���4�b��F�Y�Y����9��e:��FM�D�B��&&.��ʬ�1P�;b\�I��b�U��j�����D� O9G���J��B�N�h���{ s.�o��R�]��ˠ�$�eEf9�_<*!��v�Y/��7�'u6����!$���5�I -���r�G��<��jp��vs���
j����f�|M*ʘ��&!�&���0���/
�D�&jP�4�5��t�T�0�6I$D�o� "ǖ�q,�45C���Y����W�y�)$���8�`H�%N6����"�
6�]rZ9*崣��j�m��
��9n#
3������W&AɌ��Ƒ�B%W-�l�6̤��)r��nL���dEUUUۦ�&�sY�&�̙3f���z[�wn�Q���!��d	oȂSE%��">#�3���e=����*}�1�<��PlYsܽ��)�����\$i����qp4�p�n���6�31w|���V!ȩ�	d�Y�3�lٛ�mv��KK=Ja�hd�a�a*�C�#��H���W �L;��s*�'g�[N�kE�!i��K�"��t���.���ʨj8�nݶ�w�7��~�T+���M-�!�T=T-�S��(�ѝ>o�8ŭ�6M@棌XH4�=�PV7��&���ę b��x|n��ί[+���)!���C#�c���\`�|1�Y�y�XK\i�ַ�M:�!�0V#�;�z3fi.��G�<�#�<��$#}��L�x�?J�w��!f
�^�+���7T�����b=s��4�Ɵ949Tve׭� �0y0��5S��fYC�"��=�P���XM�eF���F��2U *:�oަ:-����O_f�o,"���52��H�"�TA$A$A$A$A$A$�4�Q[������E�M�S��
�|(��i�s9��8�Cp.mu.�b�p�&��=��D͒4�6WT�R�ݤ���TJ��]4�J�fF�Ʃ,x�C�,��A�}T*�6������������zGn�Q�<yQ����	���@��u��SX�u����17��M!P8D�����Pb$�M{����
�<�<��W���}���p���]3BK����%��# ���L��:S����1�iɸ��n�)���Z7 a�XIG|��EG^���=�UoJ�mB6a=I��T�gz�0��P�d���2HY��6 ��ޚ�j훅0ޫ�6��'��Q����[Q|��g.�њ" ����v=T_O M˵5P���c�6��v��5�2M����y�e���!N(�h�*�+ٹ����C�#+�<�������FO�C{�޻��#b6��Pd���O8���0)��k��̗f���p*��KN��&�S|0hByiĘ�CUǋ8�Nr{��vc��7�f{�审42��Flw���1����	EN�(ն��S�'Q�z,@mBf;5EՈgɦ�Q�m>�ď�\��ҕ�9�:��C���g�C��I�*T�I	{ҩYuF���!Ɗ-l�N$��Г��Т�% tQ������AVJdc#B���^h^51�k0Z(��i3AK�f�
�Bd>AO:e�ʐ2
Z�I�S�\̃'-iM�\ߕt��c�|��-���o2�B�80Z-�7��� �~ɛ���4At�V4��J��h 5�T-[*� ��ǰ��q����|*��B!$��?�'�%��8}����8P��`�������'�~�Qj%:%�3�5!<0���ĈZ	��,�e���6�Ȃ� r�T�?��~��g�'� �Z���,2ݳ����R(��s`�{]Y�\�i���ݐQi"��Ē m����bՅ�<O�-��ayp�hp=Ȣ�\��H�t���=GQ�@���A%\!>}��C���%����!9��=���߶h�{Ou{�4 �;Ɩ;��>Jr2w���C��&�G����,w�JS������
tr7�%�@��S��7Mb��v���K���\����*ϻ�`!�b����pY}�P����Q�4�
[ފ/�����C`�>ȧ��J���g�tw���F�C'+W!�9�$Hw��Nz��<�5 ��������O]��oX����z����Z|��q*���`���&�����6Ө�63)�X�#�ԧ� ���U��p:����q`�� ��F�&0��a<�7�p@LE��q���Bs'0�R�'ߚĨ'��$
.�[u�E��F�%"B�m��RG�Y/
�F*f?��x��e����ظ ��#�ٶ@��t����@�.wPx�8����y��CS�M�}��N>�Cu����4�'/k� �緵�1�ǰ/��e�*���n!�Q`���'7�Dx�kۚ��`M���=��)���}K=F��t3�K����A}�
�9�IjBR3��Hi�!ˌ3-��c[�Z7x2'$��!xA�H
�k����ܑN$(����