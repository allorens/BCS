BZh91AY&SY�c���I_�`q���"� ����bF�                  ��f�mZX�M&������fƵl���l[ѨR�m��[c-aQ4k"�شj�Z�e6 �J     
5���v-���I�mU�`�����Z�+PU6�E�h�ͨd+!$i�F��$Қ�J�

�`�ԭ�i t�m�5n s����4� 3u�#$p ���@-eWf]e�V��456j��ٵ�&i�e��[R�ֳ1m��h���*k      }/$�!U�{ u��(4�s}ޞǭwk��:�ز{��yT9�{Ξ��I��h���[��Zi{n�f��ll:i��ͳT�S�s;�UkV��T�Ie*=���@�w�}wj� �z��*��[ez�E{\Ҟ�(�y��� �����R��><�U�F�{�=��.��`���j�Ưp��iT��}ޯ��kM��Vf�-hKe��6��I@��hs�_=W�GZiz��ƃB��z�����Fq����J�ѽu�{׼��i��;מ�
����^ǥ:zoN:Z�i�;��g������m�J�CDx;bEV�J�-m��m��䤤 =�>��v�ݶ�m��]=	���� zӡ���ڪ��S� :��W���J�;s;�UU^�Yy�(@�;�z��`(�v�ި(Uz<7XV��)aC6f`�|�� 0: 9�w� ����y�
���UP
�=����PUO/^�\�A����^��Ӡւx�t���g�>��P}�v��o*�^�^�ݽ� z�=;/U����m�wL֊|�I% {�>� �=��9��{� ���  ���� f �r��ӝ9ƽ ��@�om�@�u��`�uTS2�mV��R������` �oo :���x��4�p:��� 7Oz� {���=�^�� �� �*{j���l��)J@{�| �w�=������=�@�=s�� �p w���  }�� �� -{� ��u^+��L)���7��)P,���}Nc�A�7N� �@aמ� ��ֶ P;���5�'��� g^�u���� {Τ�d�����I����}� �s� �� {��� )��8  }�Yӻ=�zj� }���FJ�
T     @    ����d�&� �4dd0��~�
R��  &  20jzb
J�~� �    �)%J�d     ��5(�h  M  D�����53D��&���OP�����g��S��;�����N�p�˘���j-Tr!�{Ծ��(
��?�"�*����Ԩ�*��AW����N���o�� ����V��I$��"
���(=���P��"p��.����_�='�l���6�`�`c���&11��Lbc����Lbc8��&11��cL1��`����0q��`�S`�ؘ��&0q��`c-��Jbc���11��f1i�c8��.11��Lb�#8��.0q��\bc������q��`���1�l1�L\b��&11��cl1�Lbc��&11�l�%11��`c���&01��q���%1�&01��bc�����&01��`c��01���q��`c��0q��L`�b�11��Lbc��8�3���&01��Lbc��&0�1��bc���&11��\`�-��`����1#1��L`����0q��cl1�LLb����0�8��-�1��L`��11��b� �0a��1�c ��`�c �.1q��`��c����0q��\`����1q��bc�`��8��.11��H�C�Lb����01�b����1q���.0i��\bc8��&11��c��0q��Lbc���6�4��.0q��L`�����11��L`����.11��L`���0q��\bc���.0q��`�c�Lb�8��.11��`����0q��\bc�&1q��bc���&201��L`c��&01��alq�L`c8��&01��`�8�c���11��L`c�ƚ`�ؘ��01��L`S1��Kbc8��.0c�!�\bc8��0q�a�`�8��0q��Le1�&1-��`�8��0�&1-�����&0#`c���&11��`Fc8��0q��`c�c�bc���&11�0�&1-��`�����8Ķ&11��L`���ٌJbc���&11�N48Ķ&11��bc��C�J`����0cb����11��bGL`�8��.11��Lb�a�b����.0�L`�8��0q�c1�c�.11��i��&0m��bc8��1��`��1q�l�%1q��\`����\bc11��Lb�LLbc�8��0q��Lbcٌ`c��&11��Lbc#11��L`�1��L`���b[8����0q�����&11��La�#�bc���&11��bc �c��&11��Lbc���c�Lbc���&11��f0i��L`�����\`�S`��8��&11��Lb�c�Jbc8��&0q��m���0q��b�����#��01��Lbc�c6�8��01��Lbc�$`c���&01���%01��Lbc����&0�c���&11��c�Lbc��c����0q��\b�bc�8��&01��bc���0q��Lbc���&0iƓ���&0q��L`c8��F&1q��Lbc���c01��bc���0���Lbc���0q������&0q��bc�Ħc���&0L`�CL���.1q����1q��b�8�11��\b�������0q��bc8���%�q��bc���0q�c���11���0m��\bc���.0�0i��bc���.11�1#1q��\`c�`�8��11��e�1�L`����1q�c1�8��11��`����.2���11��`�1q��e1q��[`��0q��\bcc0q��`����1q��)��L`�8��.11���&1q�l8��.0d`c��1�c �&0m�0
`��)�G�1A� ��G��b��Qq�cH�W�� \`��Tq��1� ��1�`��Eq�.1Q�*8�P� 1E� �1U��G��`��1�0Q�(8�
b�1T�*6�G�cLb#�q�0� 8�
cL`)�q�� �C�cLb	�1�0�(��"cL`)�T� �(���cb)�U1�&1�(8�G�cL`��iƅLb)lA1��1A�&11��Lb� �1�0q��L`c���01��`c8�c���11��L`����&01�����.1q��bc���F11��bc��&0q��m��
`�8��.1q��L`��11�ČL`��.11��b�1Ɛ��8��0q��i��.1-��`�8��0q�0#���0q��L`�8�6��&0q��bc�b�8��0b���bF.0b�1�c�&0m��)��L`��.0q��L`���.0`��0q��\`�
bc�q�c �.0`�`c6��0q��`�8��&0q��Lbc�`�8��&11��`��.4���l\`c ���?�*=w��@��<�c$3����(�XQ�F�M�Z��B�d�)GD��c'!��&Z�x坷�St!�%��b���7k8-����b*<���޽��=�KJ�,�oVMmԗy5b[�㩁=��Jɒ%������d�2ȘЍ	�d$�w��d�Q+�(ʺı���2�eR����;k2���ǭ&,ݲ9�"�֬��WX�M�Uu¬�8<���	u9�.7�^,�M^���M+��X��u�2N���jS��q�+e���tRˊ����1-M�;di���ڗO*�X����x ͢����E^ɻSl*8�G]g
@ �!Ȟ�A9�SD$e�;@��W[Ea�d���jQ�-�1'D%��2�R�NY�,����M��RH��˫��9.ꬪN��I������ٛ�P-��S�h.	�`V�S㇃�t8�;N�;pƞ\�jU��F�̒�J���Pd�EgnD�	H��W���jh���[�&��m��z24m�^�4´ͩ���JG�B�/P"i�Pv�M�E��ݒ�9�sZ��b�s�l�]佉0���=Y�^�kd��,ʺ�x/!��"j�חc.m��P��h�wtW�tm�ᵫ����ca{��\v�e���1������JN�ۚ�%�#����uE�5j��S�n=�`�Iڅ;7,�S{c�ű����l6�ƒAKق�r�Wu��f����-�+�o����M��N��Y�|dQ��ٛ��I�d��e��y*	������C���X�-��v7�뺅�hM=L��ëC�-V/]�yiV��m7�-d2N�]�|�m�ch
��,n�C�5E|Q�j��L l=����k��έpV������Ƽ[�JXxh��J^[���En)f�J�d�ݚ+�n�Oo!��2'7j�cX��>�n�T����m�+hڑu����5�1e5�M�Y�U�����N�Ȑ�6U�n�f��i[-3�Y�s\oRF�=�A��Vn��|��գ��&����-��fʉ�U���Բ�j�o&9�)��$��2��N�2�B覫~�!F�6[��!����!����L`��Z��p��5�X�(�x[�;�*b�{r�,9�=�1��'fۨ(b�@�sK{{��o
�Z�W�ޒ�д�Zi��^�r��Y���=�Gq�U�34&�7.V�ʼ�X��&l�̈́r��y2�h�xIq�GJ��v�QYM����͈�v�i�\�q[�.��.2�2�;���u�fӇ.ե[AQ�j�YW4�n�6a%�Xi�R��z�1���+fF��d�E��L�A�[j1�fb�
�h��b�8t���c9�����1��h᪊�9�]��j���(Ꞅ�h��	��BKN�b�6�ʣPP�y�an��
�5M��1��'��lk�S6߭LU�s�,9���Y��*d��,W�����B�'.Դ�'�{�I���]V��^K���%1�pSد|հ\����i1b�m���KŘ�T�8�hJ�BV�	ᥧ2��m$35�қ���f�%�w%ԓ�5�^�һ�I��k�ط���2p�'
ܮ�צ�R �Q�W
ی�"���9�x��L�vBX�R�mA�ժ+O6�r]!G33e6P���H���e�f�1=��K6��f�f�rX�-�Z��j�F��k-�� �����,���O5�]���m��.@m�âӋv�4�VM�w[EZ̐�Z��h���6Jr�U���]�4��Y�mc5p��2��c:V�����Jy�ha�������ʍ�Y7F����q�m�8^1�b
���iA^��R��[֐f��y-m�oچpŪ�ݝ��e�t8M�x�	a�V��+Sǯ���.��ú5���m�:/��ݛ�K�A�*W�n�,m���VU�X�M�6���u���mA��1����-��Uv��qkܽ��S��N��F�P����׹ݏfS��V�B:;p�1�qmݛj)$D�)�^i���W�n�w5lq�7�"L��-V0�2�֨B�qjH��mf{��ֽA����_i��GU��=!B��׬	!��t��G5��{���
�iLY���q��Y5)ޫ���y�#T��p����c̪�r����[z�T��
�%�^�[�KeY\���*N�3.Ի��ҡR�P&�cy�s 7��,@�9ou�b��Ia�e�j-N��cm�X�[MP����f��Se.��e�Gj��_j7���k���T�n-w{z5��W���U�ݩ�gr+	Z���=��H�
�˱�Qw,',-��[��MB���LH���n��4e�6�`B���Z�5�a΁Q�y�"�EhkR�����j��4[��U�h��.nVA�aI[z"�0�NP�ɡ�!N;�2�傘&'����:��&�����P�I�-�AcR�"����2��ǚ
'I����U��xʧ���;�q��-Z�%!��G)٫I����n��uS�U6=�N��d�r�Vd8����Գ5Xnk�!SS�2�E��[�ݰ�b��q���Bi6�GH�n�6hX>O���+!�'[Zfح�X���ڹ���Y�v���M�J�Ә�c#���c�+1Ų-��u�<�����w!�f�aN�'ucVac ǕE���4��]�Xnf�Wt겲(��2��RA�W/1���V�iڱd�)˽���T4ލ��CV�B)i��D5����ݖ9�Z�#��aC�]��ˑ�):"a�~�Z�z�eܬ��ڪ���2a��=��iU�؞1$�Ø�d�H���UƫK�4ɸV#��2��T*�=�$5W$[y^؞F*d��X#H��/m*z�㺂yE��/�g[�:���gTih&�7���Y{��G݃5���D,���V;�V5&l͹D�%���U9[w#r�c��bٲLI��wx�Wل��{i��"�ѻ�7Ol;9U��m��X��rܶI��,R��T6��dc1Th���T�b��0\���M5)�9&Z.�F��C��N���Y f��՘�x>�Y��N���kH��1t� �a�lę�j��i"*�e'�z��<q^-��c�#[q4�{�Ҍ�����h4��ǩ��,q�l4��;�[%f"�hЮ㹄ÒB�d��E�@��~z)�Or�̴�\Bz�f���L�TŹ-,�h�x�-3
�t^J�vl;�B�BV:�G.FH�qfا�t�&EV�	��6͠���E`���ą�9�-���9[�p+���U�`�wZg+2>�K@��g_^Y��m_7|S}I��`�S6Y�.�mJX�4K�R{M7."�m�W��V[tsm2�V�ƙ�A�\��Y��w� ׎��:4�^%E��6VK+�-�ǰ��Yˠo��6*� 8��. 0��
�Vwl֭T�A�4��'��l��(��4�$~�F�Z�*]���To�gk(�{I��z2���;d*ݶ��`�Y����l���c�-��!a�q�І�+n�"K�¥�XI�+���MݕV��-,T%*Ueټ�aA"�-��y��.��u�s+mǍ`ʆ����*�K�i��� ÙW2���B,����,��ݧij��l/mm�.�"
V�46�f�Z�n	yT��ob{�n�gpJn֔�֡�&o(�я�vm݅,J�,�������ϏwU�VY� ��oנ�to�mD�zy�A���w[I��kÎ��l�4�0)omlSl�{L��eKki[�-z^�	C�n�1m��!@��pL�*��ks^�D��@�Ȏг��6�J�ݙ�v��:�*2m��-ںƆ���T�����;Pm�)�1Sp]��("��l�Rj
�R/UgTnz:�HB�����7�m:N]��E^�����c-R��t�"�H��7L8��k)�e�[�� q���N�%ⷐ[�j1y�`иm4̫�pZb�^�b����n�Jݽ��Z��6���,)�Y'o�J�߈D6�e�*�,ͪ��ƒ$hJk!:��J���ǷoD��EM�)�����d�oV3�V�\ax�;�W��0�Zn7zm�M�[� b�m^��N�Tn ��K`�֖��i���˺�2��i�E�A�oi��t`�d��w�v�>�]����1����t�(�$��r�%�P��jw�0-0\��e-;P+���u!��С�{u-K�ef�Z�ۛ&ɸ/#@�&8���%A��XYQ5A%f�y�V
t��ɧLW~0ʧxM�I� ���p�����r�dX�n� TC��D��q�T��K�z3%	*���Z2��-6X�4�Re�e�B+���e�0E�e8i�P9[����w%��V��Mɦ;F�j�u�n�Vl��8M^�r��=NC.��
T��Įe�5ˊ��(���s����]���` �ݝ��#�*�v�!�x�)Y6k݈eį.n��˕��?QY���cQ[YI߷F{)\�E����7F���iV��1��6[�#W��t�V��x�卒e^��V�R�r�D�j���1���ըa�d}Ǩ�^�hn.�4�{�P��ᬤ��n�9�ea�pD5��cV��,u���y�̧8+t��J�n��hԮIG[y��me��7r*7-m�mM��B��Z�]̻��n틘����Lgt�8��s��!˵=�֬[��Z�RE��Ah=��^��l�y\�j�Q�b𵶐��'���VZݱ�A:�غ����!Ir$�a3A�\�������Ԥ��M��OU\XEGUA�.�m��`{h�i h�r\�b��Vn�̨��H,���+�;No�?"�����l�oe�*]Q�	z2��[`; .x�2����/�b�e2=�h�v�Oh!˘t\�W
[Rc�N-��Q��n��P1������2���WR�j�Ip���Ȥn�Lae�F�E<�L/rF;V��Qhܸ�E,��`���-^c�i�]=5��ٷ딜;kJ@mm��/5^Xb��b���=��^ѵ����#D�fP%�d��]#�pu� �={��ڌT�Ct����f����b��ԥ�i�ڤ�KQ�J�R�P���n-�Z�[�rI_-�\�+�mm	q��kb�K��t�,ĩ-I*J⨴�%|�Fҥ�[Wijz�Vr�[��졔�u-��E�eZV����*Y�Fm(�L��j�m*��F�i-7V�U�@�uU�T���jN���p��s�6�Z8�����:.�TI��\�X�%x�X5-=PĚ}ت�ά8��Yj�<����(�"�5��z�F-�-U-�ֹ��i:]k;I�4z�JKu0f.�99�L�9p��;���`��U��P-�E`��Sz⍬�Ȉ=����.�v�ԥ`ծK��%զ����N4�le�_tYP�C�n��'��x��:����NWkyD��˝|	i4u=J���&�%�m]%��W�b�f��(��X'�E9p'U%"��.Km\�-4�U�u=J��\����HK�6C�]K�jJ*IE��V��uBᴒ�W�Y�D�VT�j��ɀ��k
5��W�j^u�iZ�e��C5H����;[�����Axo%�T����UK�(�'ʒ�L]܉S�/^�ɇ�|͟_K>W\�mܚ�Er�r�,j��Q��.��6e֤��M"ւ�TF'ʁ�C&�y.W���.r�[k�$�*�ԹrR�պ�V�%�V�bH�Y�b�S嶯Ś%�T�F�j4ڰj�ږ-�����\���1�R)I✮�圍&Z���ĹKI-�x�;�R�T��V�9��bT	���U��x���:�',�0�5�]�qe+��<����]H������X�x%�� +QĹRL�q[o�����tK�Ֆ��B��R�b����e+Ir�6YJ�7#�,F��19|��v���b��br��fcY��KZ�H�W���1(�KI�mSYi,����J�zf�܋9&����)]$��X���v�Q��`(�����őD��`�Yi$AT�Zi��iڔ�����R�T�Ke�K7z赜�%��'t��Mj�u��+�w�
�G��US�F٥|�'�r`�*-�}�&ږ�U�\�5JjT�'�5-Y�v۾�Ο��OUZ{�˕�$�IbO��t���9KI�Ib�J������ ޥ�9D���-m�k-Ljb��OEԴIbʺ2�^,j�H�&w;�kygV	Z�w)V��u>I�Iڰ^'J�]�oqSD�����z�,����+�1&�%�un'���N"�5��ع��Uh"��e%�Z�w�rT�����ʲ�i▗#	6R�����h�MtJ�T�O�h�v�4�RMh%%k�0x��1e���KՖ�R�r�Q���x�"���8k��x��ګJ�Ij�*]j�bȳ�R�Sz�[H�Ig-��J'ȴq;Pao1��V��՘���� U��IrȐ8
�qcM����v�qS6b�UK���T��K�D�B	j��XF�I&�M+Tx[��*��K�W�utN'�qX8
�ú����%k�TUkuJf�c��!R�U�qLX�%�N�K7��[���T�H��_�I��mo(	���M.�$2H�%+��_+�4�bE$�ԁ�V�4y L[�M^=j�V	�!�U�j�S�՝s���@��/
���n���vϽ�Ӵ��T�O4,�y��U��Z|���R6�w�^+��ά�q+Y�b�Zӵ|��g}r҉Ꜧ��ҵN�Mu�ev��'O���m�P�9$����T�:Xѥ|��l|�5�R����uR�C���תӷ,�O�^PF��w��ZĩHk�Zͺ�[����;V��R �)J�0��K��Hi$�v�K9T��0"�E���QtOV%܍�]NT�Eԕ�I�I$�(�Ij�O�ո�&U{T�ŝ��Ŷ�%�"Z�]�"�kK��U#~nZ�F�j�SIڭI����V��)����y(�\�IR�N�4�QSUI�ٵw|��bQV%�����1%�]�)*T�j����8����4b���[Қ�U|vTW�ZM8�+�RRO����ML�����H����ߋ{�@?�ޟ�����_��ߊ����$�I$�I$�I ���&]	[,%c�	y4��5���j�#�ê��QCg����@��|:\�Aj�{���7��jX4TꝽr�;2�c�EHօ�J�پ/S��,?9LJ[(ZA�*�ʌ���D��eI��
���	|��i�ck�,�U
�҆�BV�}�xbc�˘vus���w�%��9��.l�a7����5��T4�1N���&ro�L��l���C,j�}1V�;���sq�Im��2u;��r_a��[8^]u�����yo̭rJ��e9��*��	XHE	BT�2�z�8�n�Tt$�8u����)�R��uCs�X�w�#���ݹ����Jea�s�t/�Fj�����*�.�u��{\�R�[��pk���:-e˞���0s;�"��i|�b��)���[c�s&0�o#j
����TR��Z�;{�$+u��gcά�Kjx�Y]�j6�M��ې_N��)���V��|���%��
�{#�N\��<9G)��Rޝƺ�Wp�8�v)T	���r��p���`/`Y��	$��H��a�|L�A�d�B�5�4ym��Ub�΂�&�\w��B|��`p��*f�+�����5��z��x
��k�ݏ����T���E3�֎�էI��Mg�H����n�ܞ �m��c�(AQ���r���w�s�.��������-��\&�cG�mM�co�F����K�݆v#��,\���2�Ţ�%I��E���Y&�B����0�n��sp�)U�p�{��l��^�y%rGH��)���`���oV��j�h+����
�s�l���3>�I*���o.)��q	��T�eQ���l��)`弩�h@��R�)���qՓ�O���5��Qb�!��چ�V�5���N�9�儸�얈l������u�̮�D�%���5ι�,�J|�T�b��z3T�[]�����;��Za�����e�x��ow\��Ya��Ωdec�N��|�o�omٱ���[w��Q`;�����L득_T%�/(�Ы��a;��4��o%\̸�1�{:_t�e��̥�l���]L�wɕ����/zgD2��S�rãsj��Yֈ��CT����3]���˧�$?S�__)T�O���X&\�f�m��;G.L7�m�+a}3�dۑ���6�lu���.��/�S;jp����[	pZ����҆��2�v�=xn,�x����T���Y8�X��H�{\j�m��A���!7�,LDt�,����z��S�}0싧���&�uj:s�)v��ɺcv�/ne1����q�ar�eͳ1�cQɦ��;�֝���^��\�C��nv*�dZ[&��Y�LΫ�Es2����`�/���-�6�:�B�N�*����n���>�Χm���4�{z꛻���T X��.TƍMɛ5�;͸X�{��V�g�����tS�8�N���ᘻ��`�yq72�$fZ9C�k���9�$��\p���)�G�ļ��h#j���YE�]i�{��푲��e�F�۸%!ж��o9	wy&c�Ӝ\�c���$jJ��ٹ&ލ��Oj$�w#qNu��It9֬<S�`�O2�B�F+��.Gv�ohB��.��v#�/�lj�u��^��7*�x-xR�!�
�H�cUZ�׆az;�Q���ȝ���]ՆEs&ZK��vu�	��L�w݆���s	gY����>z��d�1�յu+mZ�UD̶W֪�V�ޓ��w⬠�U
��Z���֥[���\�E'V�RSs30b�4�-U��Է]FcG�Riӵ����:��������Z��^�d�7SUɧ�}r�1�Y-nP�Y��6.09wGvs�bV)jw1'/��-j�s���w8��Zʕ�Z�'̨�¦���Cn�
��:����IԽ��|�U��;}�u��g9B`�4Z�-���|���%�%�pg��_t��K��c�7!w���M^�sxw�Dx�7K>�b�`�e�\˨#浬^'�m��J�w�%�r��,�2;��Jh��}�e�2���ڸ�^U.��m郲й����L|pp�����G����'��Y�|t�eZ!�{���Ɓ����z�&Cd���,��c�b�v�79���p���Z��#�m+�սu:�j�hGy��KY1I:��[����?z��F]�5	��:tՊ�]f����'spLδ.����j]��n<,8��Wߺ�'\Ɍ�v����T����ș�)��`��R\�K�k�CƔ�N3����noU��V%�㘴s*u̍X��[-�x�;#7Sܳ��w͒6]KcL��S�qs�༹�V�3�c'%L�/P�q^��9Sz֮CtS\�C�� ��l=V��W�sj.�0�4⒵�N
���p*?)�̚�{��.���moJ�P�p�_!':���Y��zh׌N�y��J��g��y���m�̬��5�JÝ
�k�;��ݜZF��M��]RR��!��q�ɀ�9��v�)ʔl���y��	�5D��Z���9(է�,w�����,�5N��M�ꚍ�f,h��/4�c:ꏓ�R��ى�aԹ�o.ʁWV(�t���f�S6��O]���b�ZU� ⋲XeT�I����B�lO-)�(�cG��(�о�rt�j/S�VogK�]e:1�b��t�����lJ7�GrN��T7Go�I�*��R\v.��U*پE�FQ�3�\�Ю�rЈ�������\F��:�m���я���+����G胅�� W�2�7�g֜Oٻ�k�n�m��f�[O�i���e�l�
�Z��W�zF��<�j�A�c�ƴ�\*Y�侂�^�ѩJ-c�)�t�Ȥq6Qt�:�Z��a��rOJ��Ύ�7����Ns�(�6D�`�ݚ5ػ��ub���B��0�r���U���gn�%?��x�R%n�G�YlP��=�_{p`=�c���uj���#�E�\X�ge�2R��鷘$��5Җ�F���76�.c6�ɯ�q+	��fE3׳x�cB�Yq�ٴ��D0]�ح�' ��V:�P8�n����=�\j�VFF��`���M�c����c5C��;uB�rùN�[���x�1ݙ���Ak�о��_�9�b�������Z5��'{"��rۛY���]������桀���1m?��7%v��d�� �_\�);8�PÎl\Y��غt�b�K���Ls5��2�T7��~�)�CCU�`��>g5��#Hd|��̫�C�|���{�F��2bA h��
��z�Y�G8^�t����"�s�|��I�q�ʚ��n�9<%�֫ۀ�[͖'�n��f�{Lw��	��OF񽝷��{*^�y��+Z7�u�ɋ�f��G`�ӏj!4�ڮ�tի���Z�^��;�J�7�J��琢ѹ��w�+%V��ã.�$r�㖎^���sP�t�\��j�sBm롟	��T�����L����ӗ�q�G��Y�bwH��{�p�䫮���+�D�F,�+m�>mg���	l"�{ V�Q�d�{V�P�c�����?�7b��(b��yLj�Ϣ�j�I�B�r�ƶ�B`3�!w
�u�9C��xpi�Z�t��/6�^m�!o�;m�Jcs�%��r���J.�e���Ռ�����z��;r���R+U�
$b�u���]X��0q���VM�/.��[w�3Br�wf��/�ZF��[�c���_.7y�2M���"Q�5��:@3s��`����ݸ����o&���ʾYU0�f����c`:��P��0"O	N��Z����|͈5m[W����'Wt��S�t�_�W���4�%�ZW4��\���:��O�	7��˃���*�\�9\��)�J�ZKu�PT�!�ޟUq�1�C^U��ێ�&��f��O0�q-iUHi̹����l�h�5��$m]KӸieE6 uE��p}z�E�\'4�|wc���K6�g$��{қ`E]�\h;�4aLb�M���\Bf+�m_8�B�+� �ю�^�����U���Y;E4Y�(mLl`�Ki�):�d/��ZY���S �p*c2���6��*>�m�٥3��V��Tұ����"KFĮMxQ6!���JȻ5t��W�F�zq���R
��,��9s���e��9O^��wz���7o�]O�%�'��{;^Q,;Wb��%��zVJ۝)��f��1��}Үr,�
��x��>�7oV�s7���ڽ55�)��uA��<��j��6��j巭%}7z1�:Hr�gʌ�z�>�H�ka�I� �9N,���\Akbf�v�\-��/�����6�xe|Ф���
�ᶪ՛b-#)h6�mvjXoY�4�Ȼ�O]�x�����9�>Գwiv��W�E�DT"$Z��=T�k��%,[}��C|lo\�I ��z��\ol�j�)���9���na�f�8����Z�j���*Uӽ�[s��+�;�,5�0Q1�;���}��|��6�������~��M���j�\{�2]�;N��]�v]���y.t}+��G�ɒT�K��W\�a�n��N��?!Jʔ��}0�<�D�l��s�5�Յe�;��]WA7�#r�#���	���r9|V�eQhml�!�Q�ݲ��VWBЖn�M;�T��-��0���;�vh�6���-C
�N���a�Ԑ�\)�[Y,�y��V�3+k�x`�ah�l�o��n]�Q�F\[�ut�Z�Fd��2黰v�Rg;�.�LH�g%۠ޥ��Iڭ�f�`�a�|�r��_3�������R����ޣ�b�ɇL���!*E��/͕�dQ���I$����N�IWc4�0ɰ�2E�%Ҝ�P�[
sA���n�Y=/FJK"{%�i7��N2���xiN�����_ic��bmԊ9��斥�����>�Y���n�U�q٥qOD{go\�b�ӄ]�OC�	�����*�ޙ�N�љ���J�$���� ۍ[��:9��\��U�I�!��Ĩ䜴�$�bRI��xȥ��M��G$�I$�I$�M���������� �Ay݃#Q}�.w�2yv��uG��q:�r�${����b^�]	 n�$�;��l9 Kι�ﻨTQ� ��t�S�.$̻8oV*u��w�u
������<��;s���׻;�� �<���N��TIN��yܳ"��L��ǻ��H*W��c����xL�ˡ�2]�]*�:��%WV�Y/+��^˥Z�"����|����V�qS �_"��
�;��S���T��n"� 9"��WP@�U����T�Q	�w{b'Pz}� �h��h'����^��S��#�=����`Υ���Pj.-c����>e�w<,�@ 8�=�r��R����W]D0��{�ڌi&������5��ڪJouz�x"�؄z^?xvL��/�#�/R@{�ePw�W;�L�3�ّ����`R�E{�:�;�A��m�a�<���:�b�A*	 � �\�딃��TAAO��G�v �(�?^3���;���>@Q?� ����|������_��~���te6�W�5��P&!��[��Cm=F����	�U��`u�#SGNI'P�ug�_+��T��S�d�N��s��x!�g��]�-�̅���|��&�";��l�}fG%jԛ�����(A��^	1i� �*�aȨR�:*f;�ѵ������'
}�����«�����S+WMQ��RYY3�����B�ݖ�b�5��H,�]]�g�c�r�R�"Cl�;z��j�S,�=��áе%zj�f�9J'yF��x�o't�z�Wh�+s��ȝ1���@q#���Q�� ��/�D�2��wua�4���xu{|�.6.�gEQ�f��l��Ջ���1f(/2�7D�9{���v����^Zu)v]%��ر����ܸ��t3�w�v�UW�ia��Z��8��ZlY���ȭa�C���on�8�pl����u������'�.xzπ΅U�DT��y�
q�0�J�5�{7Fv�C��j���:ݫ�W��Kvr��z;��	{�pο���u������]u�]u�]x�u�]u�_u�]u�]u�^:�]u�]u��]i�]u�u�]zu�:뮺뮼tu�]u�]u�]u�]u�]u��]u�]u�]{u�:뮺뮼tu�]u�]|u֝u�]u��]u�]u�]u�]u���]u�]u֝tu�]u��]u��]u�]u׎��]u�]u׎��]u�]u��Zu�]u�^�u��u֝u�]u��G]u�]u�^:�]u�]u�]tu�]uק��ooon�:뮺�Ӯ�뎺뮺믎�Ӯ�뮺�c��뮺�c��뮺�㮴뮺뮺��~_>w15WE��i�v�6s!Va5��^6(�1�u���㹜Ջ�T{(%n�Z���>�����PU�������<�/��3ss�v��* ���l<�On����no���H���Gqj�caO���T&�*y�v/+.� ��:��D9r���~f��[݊f��ݕB��&ݸ�[O�RiwmD����$��̫�FJa6	���SK\.�)w�v9[�����]_�d7���ͽ]�O��E:�}�OP趘�ڼI
�(59w>6���o&�r�EJ�Sr�S���^T�|\�����óP�u���Yy\ݭV�*ޗNm��a����t��N-4yƍ�Y#T�7h��7"mǚV�v���o2UX}��k�\UoXәj���D�፬�vL������Z�.r���nXFqJ�z�������Y{�Ms�Ӯ�
ճkON̸̂��r�7E:�3:��pe��H ���Cێ`�w��(�=�D�(v��s5�PU��[�+$ݣ��-�p�vIt���P��0͗{"�s���u����ǎ�:뮺�]u�]u׎��뮺뮺�뮺뮺뮎�뮺뮺�뮺�N��:�:뮺믎��N�뮺�㮺뮽:뮸뮺�N��:뮶뮺�n��]u�]u׎��뮺믎�Ӯ��n�뮺�뮴뮺뮾:�u�]u�^:�u�]u�^::��X뮺뮎�뮺뮺�뮺뮺��:뮺㮺�N��N�뮺�㮱�]u�]u㮱�]u׷����on�뮺뮺��X뮺뮺뮎�뮺뮺�u�]u�]x�뮺뮺뮎�뮺뮺��dy؏{p�9��؊�,.����y
8�։�%�I@�%�٬�w�K�SV�Ǡ�e^ n���1��H�su����G2��l�pfRJL�!�����\Diz�o<}-���Ï-�	�2Wr�e�[�l�J��O>�6�,����Hi>̽R�LLf���'b��'U;x�5񙲋��.�/},�X-`�Vj�B�V,�(�������/x��0���J$�b�[��,5A�:�)�J��9c8��lD�T���\zwr[k���	A�^��k��|6�VG�r�]#-a���u�r�.�J�V}��/�p�6�$��:ʳ�r���i��S�ͬ���5�Yx�~]5tp���tr%�	��N�P�ӿ2�^ӂd#ҐD�k��P���l%+��M<"q���:T�����)��فR�0��ًtl�Op��Vt���M�4@s،�z�r��=�{���v��`3��N�]�(dE�ܱ��o�ﶅ#�DTᏍ(��Y�s��L���Ɛ����i��}�:�iPلdͭ��Ƿ�]{u�]m�]u�^�u֝u�]u��]u��u�]u��]u�]u�]{u�:뮺�u�]u�\u�]u��]u�^�u�\u�]u�]|u֝u�]u�_u�]u�]zu�]q�]u�]u�]{u�:뮺뮺�u�]u��]u�]u�\u�]u��]u�]u�]{u�]m�]u�^�u�[u�]u׷]u�]u�]u��X뮺뮺���]i�]u�]u�]u�\u�]u��]u�u�]zu�]m�]{{{zzzu��]u�]u�]u��뮺�u֝u�]u��]u��u�]u��]i�]u�]|u�:뮺뮼w������ �af��X6�G�hh�|ı���:�%����,��Rn��fN	��+����e�(�����+D��+Jx���j}S,��[z�Y�o������������ܾ��qi���]�F��Rw��/-�����ӑ*n�n��e�.�@��-{nR*:3\�}��`�
��� ����WsP���VV����Zrq[*fc���T�j
N��R��HvF0%k.ݙ��X����y���Nu逽�Ilz�f�@��u�zͻ�w���9�q���#������MJPe�V�
��^���w}�P�l�c+�Y�ᜫ�f?��h�p>w>,�����\���U�ʔ#��nZ
`��)o��oqU 9JXT����3Y�c'`MtɤL!9K�ї���3-ɦ���7����]�{�;1�b(�"��m3f�d������w.������M�L 
�P� ��}��]C������vlW9�lZ֨wmAo�!{Z&�9��b�%�e<o���k�	�b�&�vh�K�b+;Q)Z܋x��y�<��d��R�A{=����Ǐou�]u�]u��]m�]u�u�]zu�]uק]u�u�]u��]u�]u�]u�]u���]u�]u��Zu�]u�]u�u�]u�]u�G]u�]u�]tu�]u�]|u֝u�]u��]u�]u��u�]u���]u�]u��Zu�]u�]|u֝u�]u׷]u�]u�]u��]m�]u�^�u�\u�]uק]u�u�]q�]uקG]u�]u�^:�]u�]u��]m�]u�]{x�m�]u�u�������]c��뮺��]u�\u�]u��]u�^�u�\u�]uק]u�u�]q�]uק]u�]zu�]gs<@�Vu��Ύ�������z��6���)=�]*w��d���嘘��T\�u��5-,�ǫ'*�ת��U.�l�/�iqR���H�낓��,��6���$�w���f1vlV)��S��f��º^�e�	��H+����Ol-=2�7r��fιM�{��s���Oq�|N��Zc#���(	�3{1���\56��F���ݨ��dx�M ��$i���5
9t]dx���A�u��˲���6d������ERXG����Y�3�������(�7�#�n+�m��ph�6e�d�0��x/Z�
�8��l��@xy%izw\l�W�6�����������h.=A^s��ڵ�f��e���Z6��ۧRD%gr�����+s,"��.-ڙZ*�ä�x6��&��*+R8�hb��:YDE��pT���REh*$sweٮE�7���ڷ�*��h�)�*��s| B��7:^zb�Y�\�<R�>۽X
cK�*��;�%׫P@݋7}&஻F�&��,Cq-b�Id�o��)��&]~��W�8Q�.�toH�FH̕[.�fF�.jΛ�;�sR��g��J���k.�'1uXC�𙔢�4�	Hk;�_�9!�ͻ�mЗ=d=�d�D֧W�}[ϒ�w�*�Xgvd���Ǽ8���I$Z`�c�HS�*Ƭv�Rz�%�����M��;���֬�u���R�1��)��S,�θn�:����Y!L��\���Iэ-KT��G-���H�g%\e\��ʲ�A�o����-̠n{����Ϩi`���a'Y�{��ڞw:�B?�҃�n�#䪆�[8��7�ּx�g�����ZQi�P�������؞nw>��f�"�t�p΍u���/:o#�&т�3ȝ'4ҙ���	�UZ�~�(�<��v�MK�u,9f���.̥[�b&�u�Nس+�uu����͈R�٧§l. �	;������-�uT��\�/�U�ݕ�oF�n�V�Pg#�Kʞ���N�B��,��p�ja��Y��^�ړ��:7!jM�_1�߾���D��{V�+-�V��@�""^Z�᷽��vRqm+ՙgB�f�4���7׻�̈́�]Qct6����8�$K��x	�4��Ԥ���f�[���c���Ӑl��	
��d4v�g�'�	�ai�D��?[���/2)nm�ZY�(���kk��ΰ���7ƴQ��X�*52*Ψl�=3��W;Ɍ���bT��>���b�4l2F�*��C;��R�V���p��㮝���BL�G�����0R��y9�k!;Ӓ\���>-�:���b��WV75���W��2��R�,��ٓ��!�	mKJb���]�O��%l�_��ٴ;s�X�&+�!���P����
���ƕ��ɆM7E
�=&w{�G7�ib�s�[|�����f�9�^D%�æ�2K����Dzw,̛8B-�,@޵U�+H�{ț�l�<+Pǋ��q�m�|��nH4㷕��{3[��=<��q��Ӄ����(�a���U���[J�ݙ�h�ܑ�w���7.�N���9vS�v'�W}�2�X�bG�
�.g�7&�lJ�o�_C�>�{���z�#v�e:˦��xt۰�e���WLBF��j��z���a<U��ˤ��`W�_X�{.X�|��< "�L^p`�������6��i��Y�(���6�	�b�?Y�>�JS]�/%��58�w<�K����n:,��Ω���8��Q:��e�m�WK��Z2g�vYބ�e����4��� KN���^8Xim����{%��wo��/�ѣx7ue��1/����>�/i�T�\3-ޤ���gۣ���3"��r����c���26r��;�nʗ�]:L���rp�O�-
��,ђ�p��C����e������<<^�X�.����;9
�'L�)Q��2�+��6a�٣I�ިo*"tĸ�-_�-��f�8ʽ�)�x��Q��1e˺��29eZ��E�=��K,�t[��܄j��\���3!�;�C/aL@�8�0<�<�98�h�E-D$#�d2�!�����O*ER�6��L}WZ�܉�f��)��܎<���<΋z������}��x.	�5	ܬԲ�4OC�
bK�K���&��C���X�a�&[ОwL�X�4��SFM��I����ƑbR��8��%�4[�����,ua"�ݷ�`e(�ذD��ݖx�\KtռN��p�t��+�63�ݺjt=Śʸ��ܢ��Xk����U��򕹆-�^t�I��J�	2`��K�O[�U�N�]���W��zi��z�FEc�75�НemLۙ9o�;�0�E]��XO�ٔ�w8��	ݴ���
��L�o�ֳ�ݱ��a�)��c��q��ƹ|X���f�<t�]������E����%I�4�Np�n�7]�n!сZs��|�RU��1���i!��S[���O%P��d(�^�R�m�W�N��Y:5-�q+��7�Q�k���]�f*뉞�c�n���
�P�kQ��&\운�#�Uol��ڎ�Sqn�{�=MLשׁLB�"&W;9��!}Հ�-~��5S	��yP��P�Ƭ�u]8#ұ�a��&U`}&�u��8�iz��{�ޜ1���M[�[Y�
N'ð��CaT���9ZΝ���n�y֟]2��Ke!]��˭��w[]Bv��_5Cl�W0d�nJ]����i0U�z�\r�:�^0�e�'�y:��+��n;����a�ZN]^�|2[����վ<)����{�1{��RZ����Q�bw!҅	*et�.�cgpD�=m*��Zvy��u؜��US%��{p,�ڕ��f1�Kz�����	O��N�yUs�A�ٷW���Qt�LYW�Q
��V��9˫�T1k�PC�,�cL�N�Ι{[nK<WAY�uԌ�τ0����;���)t�%����.��BͮF%������p��t�Yy���3Z��\��!��@�K��ݗ�Wu�����]�{�>�cf�]�����֎uMj!.�`�6�3U�w1^�FSf�.�S����qdV�	�Xi��]ܿt��Bs~���v�蘛z�׫2����o.�!���mu.[Gv7�Cv��*B��Ց;�3pv�DP�ҏb��Y�k�%�'��H�؏a��i1��Ӣ:⒖|ޠ���.�r��%�!l�m��0�ÜT�v�D���v(�K<�HV�H��Zp��}�ߤ�GW�L�G4Ʌ��'$u�%��At��ї-�䲸�f� x�K�pP����T���xT�w�J�3D�<���er̷	�M)}9�B��J�J�s��y��)빸ը�e�#�"�
"]gb�L߫$�*尶����<����DW����~������W�_ҿ���T�������wU�D:�VT���+2�l��|IL3H@C����B��O�$(� B������!��4R�$�0D%� 1����M��P&�p��	�YS�4Ē"��7��L`N2a!8����C"�1#
��HL��¤ ��z�� �q��x8�B2�m$[/�@J �SJbJXt�J��	)�mW� �H%I6�HP!�($~d���:-�_��T�p���M3�,�rB��$2�&4��d���rF�b&� ����d@��Ӎ��20�*I6N4�M�C�HCL��i�K������p���A`�DboMT�р �b7$1� i	%���QP>��B�
��"T��	^^&64U2�0��i�1n	���g�~0$!��tن� � �A�D���RBb�b8�hAI\d��*�$7�y��HR�E�Q�*y�H�Q2!�8�1��	�x,��o����c��\��5z%����F�8�^��Sܡ�H�7q#smrN�mb`-X-��Kw��ZMA�<�ή�n�gk�+�S%=*���rI2����+YN>������c�w(b�N8V��ü��Nb���.ӫ�O]wl�n��Y	!ɪЊ�a�:�`��Yk��wsD�L�i�ֻ����r�mL��r��Z��7�-�gz�z�!+����v躲1j�٪l{qΡ�`�QX���uZ������W#c�啑�:[�V�4����Ou��n���]��/`��9O2]�/�Y"���Q=�₷zN]����۬b��ij�E�N�U�ir۬���v
׫+c�c���#�R��G�Л��nѻ�com$
d��\]���Hd��൴3$eq�S��o�Y[����E�w�Q���ֶ`�R�e��g .m{5�!�1�j!:�V�����#gs3��R��wh}w'S
��"�W��D�ޒ7$���k�INI$rI�����-���PQU(
����2�S�(��0���q��I���#��lE	@�%�!�8�FE�An4��1�$�'DHlFDI$$I�6�e��C
9$���a�!)!d7@��IFpY'Хd�Ii����`�Ћ�8C�'@��eӢ��L�.&$d��PM��æ��0MBK!7I	#nH�M�Y�P6a ��j	�L�  ���#��0( L�I�&�%F�$��b"	H8dJH�rO"�r4 q�$�(XE���&�)DB.�
�d��B0�F0�$�h�#��P��8��(�R�29
� |��P�9Q��p�Yg�]AL��\'bd$pE)��@�$�~hI")4[H� �0�h� 0�(���p(T�b%�"1�����3-8H���	d�A'	("I� �R	�'�Pȼ�f1�@K9PTta��	�d$H2 �&H\"L�$��xA�-�"��D��L��$`2$Z>�H[%��Q�EP�c�	M��p�i"A6R-BL1�
-��!& RDRh��jA
`��F
m��	%D�F�5�\�"N!���	C���CP����"��Rh9$�q��BHHD��"�p@�$�R��1�a&�FI��0��f�q&IDB.�	2�$2%$~��'�e99	���0( L�I�&�%F�2ϓa�	�P�O�d	$�,�F	��	�"HIm�T�&(R�2T �~�S�ԩ) i��A�(�mLbA�>�(�p$Rd�B�	�	%���"���NI��mr�bsȄ�dD�&@�A4��4P�C �ay��@�!�J��,�Q�EF��@D|�C��_�&�!� �i�(
����"����a��R(�M�$i�C����f����wM;�;�w�N���AF`)��lG"@0%]/4�H� �R
A'�O��|	x����K�&]�6�3�rz�yC�A�#"ITU�SM�>=�u��]c��뮺��G]u�\q�u������iY�I�M�̹~�Y�P�q�2�I�mv�少cOo<u��]i�]u�]|tu�]u�q�^>�r5TH�r��s4cY�̓�q�bf�B�mfO4��2m��l����Ǐ�{u�Zu�]u�_u�]q�q׏�ú��M1�������MCi����^o�o:I�4�>��˶�ƒ�ɸ��i��A8�J�h��N�B��Q2�uT�UܔSz|{|u�׷]u�]u�]u��X뮺��8��� �v�[t©��p��*IR��Z $�(� �!2��%�����ȉhm���Km"mr��"�acm��I�9��Y�� �țd�ͬ�!��7y��ߛ*�Ke��c6�RI+���o9�}[r�(��.\	��Y.����Y�D�$�q2� 'ͬ�����M��M��6�Yn��Ȅ[o�i�x��PE&Me��13i��ιm�4���I+m�%�iʜ���4�%u�/7�k���;�m�l�x�ylM���mԍj�5*�.z��G�t\��B�P���R��G*g��96��Qd!.j�뢌��VJ.��Rʠ�29�6I8�+{�9���/hD	g���H��/d�Q^i ��X���EgbY�/9�R�����$'ڙ՝xwG7��4��%�B�)!6&��Y2H��'��y���iԐ�M��FXE�`�JI4L>bES�H˒O�p�Dm�M�9H�H&�a��"0SL6�y���I��I�)B����
I�4�h�/�	�ك�@���_tx����JZ½�Vd�W'���2�S�����)[�wۛ�N�n���
!��h��E���A"Ç��H��"�Ry�#h<�!B����d4�l6d0B�OW�1�h�=l�R��&���~lA<J"Ir�)HY���Z��a(6�*fR��(��-\�O
(�EH����If��iT,�_�Bc(��͈LaXP�!�Iͷ9ݎ5�7&ss�{UUUT�=^���	���SC����VeEJ������çίmc��:��".9��yLi�rc.`�y������zН�
��d��'�>[XC�Aڋ���IՈ��;�����D
^�k �ޝ��M��r�a<�s.���gD�I��� j<b�I���p.���a5��Ƅ�.��*hL���ӧ[�Y�@]��U�
�*�戠��:��*�!^�bNv�wR"u����<q	���w�.s}^�Y#��:>���	����ى���Q/uo��͒����ٖ&	�E�%���1rg�Ҵ`����@n-�`W��Zz}�7""7�e�wV��d��Z}�5�����kV��I(A�q:a����EC\	���,KC��yƌ$�PcX������}�0+�<��Q�I����hS=�#Y=e�(lߘC�Eh��qu`N�dޱ)=�s×+�7��\M�E׫k{�i��^	��r�.��p�iŢ�S�v���X����/U�$�g� ���!�/�V�|%�G��U�t��w��+��V8���VgH�r�:f��vw��;�i��c�;��sw7�)���Q	3ݾW�<�|���X��Ii�P�};U�'d�fEn��ͺ����	����};������+�N�V�7���nͤ�T�^��>f.�����%=����u~OÂCE�6��W|�B775�L��W�vr�=^>�v��h���ٽ�ʿC;5<D�C*�e%�Q�%5Q�`E���2=��q&�N{Ek{���d��8OM��wƕo�ڴS���a0.�ܶ���A��y���"�=q����ܷ͞�K�ȿpGق.��EY��=x3D3%**�Rt�'J�(Ђ�mU�c��}T� �sS�N$^�m4M[��|��I(��`��1�m���R�y+�9���cY�L-�"�)ʊ/p�n�KobO����U;��I�t�"��R�YY���)bk3��U:y3S�C��B��>����y0VI�7�l�n�S�����+�W: � bDq��<I>�ݺ�O~��i�K�z�nϫ2]CA��Ŗ�i�M+ۋ�ov63����<��w#y˖IWv�c�1���מo��|��n�ϣ!�Q5�����
vV���l�������=V�,�OL��
��
b9��n�@D�fI)�D�˾�푢f�ӈ�K(vzL��٤�N�O^��^��M�f��-IzG���W�J����ש����U����V�ej:�G�C�Ji�����φw�	�{�[��ʕ
�F��M�R��v��.J⁴z�{��l��|�	�0��g�����P� ̘s�m#���\�@Ѿ�����x�LN���^�����m�J�!=ԷJg�\��o�]{��~B,��Q6u��v�Q�4�D@w���n�N�	��Y�ǚ�'���&=z'0�����5Y����ӢoUeW�i��Ƀ�|dE�v�k�_:�vs��;e|�.m�]�S���żY:N�5��8p�s9,]��
���g(�H|�OKRe�Z*����9�aS���E��O����N�;U�>3Qc�s{w�1>�����=����Jc�`,�~_}�����ݵ�'3ڴA�^�x=Q/s����fe�U<��@ٹ��}�Z�i�{F�_gx�1O}��]'���>��.��}n��u[���8���%�PL���~>�X�.^�E� �ht�S������|{ɥ���i\�ҳR�%n��3DKunj%�RE�Y���6���}��T_p��ߧ�P
���>������r�t�$��E����uM��s!t��H֔k-J��;;�>�E�u0b���%��4K��[�g�Y�����z�H��L�f������~[1,�cfT�+��|�����~�mei2uT�9����`�9b������Ihʅ�w����G�_uSo��VS����'M��=$�V��w̜C���6dϕ$�Y5[l|��J��\��|�`���Gc���-��ו�t���/{���&�㐝kPW"��7�ʻ����ͷQ�=�nMʸ"೵�:i؛�����hw�y�J���7;����JL�-%@/3K�ܒ���aK2e��H�GyMX�g�#���)�PJ7*�Ӯ���l��K�fSD�k�f(�L��O���u_.S7t�%5����x�+d�'���=���Ǽ�`7��=�3�4���5��4����%1r���l���V��o�\��Y������y�� z��\���.��ez�6#�V1���R4`��Q�D�M^�>�EH$V�Xcr��P��|��Lpi�umvő��$T�bl�GQ�����=�`A���5�ˋ���&�Z)6�{7��uo����{��R,|]fw}3p�Վ�}"S��2��~�M��6&�МgCs�*@��a^YH���,Mn�ZD'wb*Vt��3y��{W��: 4��+��v���UN�r�<��f�e�o���ܲ�љ�3��-��U:�p[�녖�>�!a_m�j��G"��,i���Bt�C�$3GW�z�Y]ѬZ)P�M<�/_m�u���ǺW-�0�n��.J�U[v���]j��5���Ԕ+�%t��n�gD�G��}旕 �� ���|���/�n\K��D����8t���S
�IwW�R��r��b�7���� �������;�s�z��s���J�	!i}���!��/n2YS��w
��g��<ހ��Mz&�������y�0y8�t3z�Q�cr�h�fw��9���,be�q	�m$F�I3L�������D�VJ�{#c����	��"�������?�d ��g�}o3ۥ'#%�G�/��Պ��1z�2Ѫ{��s{s0q��O>�'�IVy�8�7�n7�\O��aO���M�a2Α���Qw���&+��f��A�:.w<��̰���;B٤U԰Ko�wgf���3��U��/"�z-h�����Tj�/$�����_z�.��]蘑��F{� ��֒���mE��O5I,ը��UM�k����-/ *��}�)�I�[�Y�Jh�R���)Ts5 ��c^����C��K��p��+t!Z������}�A2�9'���3���y�|�kRZQ�*/�Vi�vo�x���m�:��h�k����Ľ:�r���<��w!w"�KGl�U۪�1�U��_[�n�|�3	E>o�~�{�����$�H|�j�|��իm�ڿ�纊��Q�H$ o ����AQ���4� K9�rަU�bv)�Q��##h�5���倫򐒦�>q�z��[�>7��A|�~Oӳ�~#v�:�
�KǑog�l��}�Sʙe��z]Ņ��U)��E���
Ě���^�m@G�'�f���eZ�%jE�J�?�-ܥ�U6z{��[����Z����!�������W�E! l�)Q���]ȥ���w'JGr՟a%J�`�k!�_�O���Y���V����ȿ?�!c]B+s��痛��y�߯6��ו�Մ ����v3��J��nk9���oQ�Վ�q�V���]�0O;��Yi؛����έ��t��\p���T����
n�����Trܬ5�E�:������E�^�����̤�N&\�W&9�i7O����ȥ�U|⚘�!�D����M��1$���|||||D8�w�{�/����̻܅�7�Ug��%S���y��w��NGN�G!g�Тϱ�^��h]��Y�[����P��ĺ��zI��\1��c�Ǟ�&8:�N�ݺw�h�\S�����Su�����oel��N�|>���~O�{�>�sR�K�N��䊫��%X�U%�i������~�(4�G����kl6��'ϨiU@`��|��=}����딃�s����fY)��R[w:^��{�����UZ���Sz���o	�YJYG�S]�:6X��ɼ x��PX��
�a�ؼ'<����5>CSn�M�b�9[P�A�Ͻ*��"?/����!��sv{�O;@��#���u]�R�le�APTT��
�)I��k��vU�u�݆�Hv��L����,��� �Տ�Юx|�<w}������D��u7|E����/i�+>���a�).+.a�؎��q��S�K������:��]�C����,6e�ۙЀ �������WN�u8b�M��o��n�:��]i�0�c��}y�SW�V�\�z����y���&���+wآKj�H)dD)�y���`�*�Q�J�9���w�7�wNrx��>K(��(�38l��
"d�Mi�%i���E7[ڜ���x������x�{�{yR� =QUu��!�a�B�֏^�����6b4Ձ9W5o�-�S�QH�*}���	S��7���ʏT����>�!�A���{��HB��9�zPI+��7�s������TqS��W��V[k<{�b���<L*�{˧��ҏ�Fd���/P����|T�H��/\'sq����H�����[5g��
 �U�Jן\���?M]�ɍ9��o}�^R�g�Ό;�k�1I�V|l+��i�@��UPR�������b��B�:s����|���I��s_.zQ��=�1�>s����?y*�W�T_c��v�M>\ ���˦����f��R����E�o@QZ�k-H����wb�|�x^W��=W���-=�q'�N����Ҽ���75�`�t{Jj�}َ�tڱe5LV0FfI]S{�>{N�����;na����1�����ߛ�7���޳��ia��ӷ���m���2]�#�ҹ��s"󓝯U��*P���]�N�����H��l�D��`�2�V=��Eї�xx� �B�78eHI!�Cj�N85!��h�*DDz�t�=�]fbX:X�&����5V��o��f�[U���|s��������Xo ��`N�z���i5��=S>[���ZA-�t.���q�ߗ���;���5鵾��RI-�W�����S��Ϲj�,�"������=��t�����������2Q[�{��FI��>c�_��=�s���}h������]�7d�� fwL%�"�(K*�z�9Y���w�l/}�+́��ك)�CmeZ;xW>ĶzY��j������p�C@��� ~��^�����!��V�(���V|��1�k2� f�.aW�E*�[:F6����Qb�
!q l�!j��-onD,��u.ُ�9!���8p�����(�>ڑG}:uh�Dk��'T"n#V^s%�-��a�4�GX�;*U���ڹ�#J�U-��g;[�$%>���3��.��JqCK}�{e���w���9��بx���{���W��z���.ᢒ�;J��n�e���\ D���V#5��P}\!��J� �7z7y�V��e�7�_@mv>p�(�R�W;{���[s3��R�wH�c�0=��O�CƳ����d��ȳS�l�R=�\��.�������6u��t�}��xVw��1ι�����"JWZ���I��ʻ�Xu��b	!����5wN�v�6S(J�ʾV�6ΧG�����q9�f�+u��-�O��2�C���7��F��T�q����e�ʴ���~�u;�D��d������\D��D��������<����L��sׯC��'+�w^ge��!fܲ�ِ�咪i=�iY�l�*Q����j�s���]Mǖ�J��;H�H7O 2�b��!��A��L�l�:k�bD�G�0��h�\V�)<����,=a��8J�P�,0��]�!�>C�`pU���|kX��t���z�����Y��ѽ�ϻ6>t������Ȅ�qJ����3C�q�K�:�T��e�R#�V%y�9�v��F�Ÿ��JD��v�U���U�P���tsXǱ�>�!f5,�(Γ�V�\������n�pux)q����X�HP�A��&!.��-�N��E�)Nն�Z���(���+5^�k�[p�EXB8N�ݫ��Yy�[xkZ�&-�^�W���.�U��@��׺2���@L
:YUa.�d!,�up0pN��]���,��U���r�X��ժMj�^+7P5z��Zڴ��q�ZNv��T�UٽLwq��h�%i��J���z���g_6���w̬�1����W-��)�s��ܷ��)�[pՖ;h�W�rD`�CC��i{R;Y˛�������uҬ#f�e�n:�V�X���\��B�j�s*�a��j:*<y��2��M�Z+&���^���k5[���zHܒ�rH�I$}$�H��H����ݚ�e��!�γ�='�<��F�.$'Wv3�6��D�i	��gD*5j�䦞�q��__^�u֝u�____^>�������m���O���T��������2">l����.X�d!%>m>5�^9�i�8�����^�u֝u�]u�����__\m��^<|925@�C'�7�\u��-�'e)Q��\�PjI! �U��z|z|u�_^�u�[u�]u׷]}i�����}{x�H���d	$O*�U8���Z褞[d�Bv&M�˒��Li������ק]u��u�]u��X믯�N8�����rJ{��� �u2��ƥ�k���8�M���u3Oļ^�$77q/B�jX眇>i��TDXC����̞o��$T�i0���R*rm ���,B<M����$�Ma��I�NO?9>k�H"�6�\��,̏4�/]���X"��i�9�_<��ب#���M�s��}�DU�(C��<MC�"z�Y��q9
,E���������yt|���;�"	J��"E��|dT!@��|I ��CaqD	�n�2w;x��u�'�5�&d�&}aI}5�+����Gl��ݏ[��rIo�zhi���i��i��;��R%�,&}��l���K�O�[�G�]���ʀ��;� >X7��@�и�v��.��Bz.:��w����po�_����R�߯���B�?�B����n@f㐙>S>�Z�0�&
M��^���{=^^O��kҹ0���i���}��̀⅏���(j�F�S`�,�A=}xx��k=�"����Ӡ��� '��|�;c��χ�p=}�%.��<ܗ==�g�R=�������uvKr���/#�?ҝ�~Θ|>����߾z5W�c�~~a2)W��@u�>a���o��U>3v� ��X�����W����m�a��ٷ s��b��Rq������x����< �[z�u�7u�ޫ$�����%�8	������>����������� �[z�1�Nt��P�P�[�m��^��n�����%�|p(M�1��p<�}9�g��%Lgº��7���)cz"b�A�]{�{����"�@�ez�G�9��g��K�o�������n`$wc* ����k+��G��[���7�_{�z�<�SL���BמBs���G\o�F�s�-�t;5/�2�/��7f���2�T��#��V<�Eyݗ�N� ~~~�d�;�f�_h1�_e�v��x ,��W��z�c�U�شV䊎�ȷr�i-�X�ͥ��\�am�����'c=ni���u:����>��cM5�M*y��8�ۛ9z�_0�k}f;�}��Ih�� �C�^���ߗW� �� �%ٙ�jzN�=�.e�����ocS$cK��?��>��b�>OS�<`��DO��V�˻����3����x�������~u���v�&�л�^y�2��RxC�+?/g��u��H5u���P6@����<�΄����Ժ�7���w�p;����n�+��f��!8p�����r~Ճ�������|9�W1�]�͕ڵ�{���4=o��jɾ��&�����������'�{v�M$Ǡ;j|�&'�$�n����'C���Q�9�H?��m{Sh���vs=�v��.j}+M�����;��7�d��*�g��/nO��C����~�47�����>�$?�+�랪���i؆���I^���̙c���xrc��Lo[�c�[��@�v9���K����:���?G��xF����	�x{e��uw{�����l�[��sύZ�h(8��u2g-���U��_���c��W9�)��qk3~<q`��y����a@>(7�?�����N��U�Ii��odPe0�D�Á�N���ɝ��6�;��%c�l�3;���np�ti�(F7�fKi$�U��%W7�[����۠v��Ї�{��	�8�5����z|�b	S�;�0�N����rt�0Hd�m���`����Rpü�m�J��� ����������g����///oؾ�2���	�ۘOuӐ��p��:��4a���R.�j�+��۸&@��`�Q��7#/eVU���;�*�Ǥ�O�tU"�I��7��� )>��*:p�����, �:"��4�y��"��ڭ���[�tޣ�����\⥕[h~����{���Z� yT|!�}��Y�g�/O� ��������R1�����������a�[�hp� 1�G������P��'���-2'߈H�l{�
jDbz`6b��<�&1���[{1�2z���$��
}-��~�X۫�m�W�s_���<��s�h:�'*��u+�I-��� -�: �r�REnKɼ�ӡ{���Y;����y�2ockl����,kWR ��3�z@K��5���˿�i��Sg���s�J:�xx�������^���X�8���H�� ��Xj{`5�K�lTz�]�r�t�.��=םp`�������3u�����s������M^5�����ֻV�%{�@�g���F�t�Y�]��+�����ve?��X&�
�5�OC_���m�Q�7��=�N��[Ǉ���J 6z�̛)Ö���Y�6�9�2c����=�=�*@fM�i��;=tsxRW�;�����_n��<=�Z�-ـ���8�y��[­�x�c�qwh��;SsyfT?3��F�Ґ��}rՉV��$�u&�:o��b�:r��7��h�:���ևR
V��kC���-̼�HIӰf�ɄY �K3���a�)���Lt�z�Pp���HO�#� ������>��hi��#i���������ܐ���:���9�aϭ=�s�9S7���m�j��g�c�HbA�Y���|~����3'Vi@x ��?��ާ�zj�/�����].!��@�����:�>͊go�Y��f�]un���𓮲!Lĉyj,�ܘ�~�#��*�.wVyׂ�'�3X�����6��{�l|�Y�����{1ׯ��]��=�-��q�g���O�0/C�ƃ<h���.y~���~��m�(�X�%v��'�t����J��G�ט�Z��,�@�?�0(�>BK���y��ȏ
��lW}�o���LR�Κ`#̚@��37�n��?=0�����{��*�4���`f���I��aM��=>Q�|��/�E7wp�ü�-��w B}j�\�g�z�6��7�v𣏕�u�M�a��	��^~X|�����>����:��77�.�bޠ�c�f�f�zm���zf'3+�xx�q�z-���s�_վ~wf98^��y�?�8�F��?��z�,�ә��[Ǒ��|�C�v������vr�墤�����g�Ӆ��~n��	{��K�?kcVT0,%�km�7f����ͣ�mN�*s+/�Gp]XB���)����݂�l��T���U:��y'	��Y������p�KM����h�ŕ��EEu��.���xo�B�0����4
�n�W]r��]u�Kl�ȵ�b8�x=0������Q�hos�`��n�����3�-ϐX^ts^C}�#`N����lw�<^���?���}�l�w�,�^��)����ڞ�Ңw���(��Jp[����rv���x'1�y����v���7�D�p;�0�ٰ�ļ=�C'�D��T�Ó����i��ښ��\xx6:�#l#z�F�s�,�wpwז{=�����ʫ<(�Z֌7THcs[��R�xx0�&���f�m����?y8��V�w��`�G���k����w@	��� T�}�^x�`����v�i�[=����M>ǎ�E�>~W�׿|������9�V���΃�a>� 34d��`ή����< 
��,�?�a~,�}�!���~_X�y�Y��o���!�3�� �}���&0�q����	n���l��b���������P:~����n�=�g.U�<��~[y��� ����Qr�<��Q��	Q���{��*���3ԥ �$��>h��������}�v�g��*��#�w��_��Ah���q}<s�>=�g�+��>ÇE��E�I1ã�QwHe<JO��ō��x��B`A�Hi�z�κ/��񮄌qu�Jȫx\�*�lvGVTt<���o�P������\�[˛֕$�NN��S\ ��.���v�*J
Jm�.�{�ĪVgm���*w�rC��i��i��i�1��B W�s��o����r���Po��	�n�:g�=�}�M�����MM���h���݉ņ�!��^������mn5A���b%�H�p����]6�c�{�SO
�z]��X�OY�Oi���u.�f{��m�_p�=���٘]�@��U�_^�{��}�k>��M�\��U�u��=�^���W�0j��U�9�/���J�_�����Z�XA��ݚ�,Ŭɦ�월J68{��i��C�?|�P�����Kq^y3�<�|���s�?`��y��Q��q�'W ��y����=�y�'L��*�ޭ<�eQ�wP����ۓ>|����s9��/�����iὍ���7�+��a��w�NǫL�^|�u��'�>��9t?��Ӗ8F��XO����(����yH+�?K����1��䤰��m*Q�M�F<��[����w8f��v�)�z�a�o�-�}e�����徣�gɎ;?��y�ͤJޥ>�MO��<�dKy�-i����Cgs���x���U>��W|�w���<�h_H�̄f!�8��m�u��Y�2]��v-oN��9��N��4�s��C��{� 
˭����ֳU�}��kEK���-�0dz4��dvE��q�"ͫ�w�f��ͅ�ո�e��>�!����#i�ƚ-���\�����w�ϸf�[�u�̐fD�e�hζ�k$��6ː�9��1���wiv��ܱX�r��4�O��D�ߏ���;��|����=-)�2x���$�E��yޛ����y�Y��/�w#�{Z�/�č�Aa:�����QN�ϖ�ƴ�Ϗ���
<"��>�l��V��kUT�כ�x{�����#���!���A�^�(�ڮ��]�����5ϐ�!8��=��M���<h�;��p5�9Y����A�'��Pc<�L��қ<ރ��+|}F�z�E0����.��5p��r�!���F߽o���A�>���z��BW�cL>7�}N�	���w��ׇ�o�OM�`�:q�z�l�J��( !�/� ���@�W��zy�5u�ְi�e�6R=��L3�k{�(��ܺ��ˆ��ha#���E�ߟ�~�`�ga�}��f;M��W��x �lm�y<����E���:<3�L�M���bV~y��{��<��/��6Vg^7�i����W��>������ͽꎙ�5(,J�v)0�%�����f�nj[t��EpA��������u�R5�6��V����`-�$�X �X =;�ye����t���񅰓��^�^������eennհ�����)�*����4�ÉzE�
E�O��W[���t�=y)�@�Ü���2e^���]�n�]���N)be��@7��Ew�g]_��u���h�i���B]y�֓�{ޖܟ�� �|�t���Ց�9/^ 0g���p+��5��Ww�J*��8U�SSSgl�|G�=��A�,Co=�� �ٞ�S��a�
�^MWt������դ��nn���n٢��gT��vz<��ϫ	�Q'^S�����c�o��˟-�f�EHn��ҍ��_gH��k;�[�\�_�0��@+��>��\�ό�n�k
�B����+��� WP0���?�@;~C��Y��c��P�^ʹH���'���K��\˙��~�8��1okKt�o7���[�[x`������ю��|���v�>�'S��O�d��߀�N��e�	��M�ӟg����5U7��~s���ě����^Cf�x�ڶ'C�A������-�H�8��Q�_�W�)��͎_-�_�L����)�c�a���G�=ќ�t�xV�
�[�j�@~�V�������3�������G��MM-sUjҷUFi<x"����u<�G�[Ú�OH����P׶~zkw�=�����y����<�>����-��] ������ov@�j������_S;�d�]���u7T�G;�U���]���l}WUD�^G��AY3o{�
��{__G-^b�Cʀw/��p����4j�����R���w�{qN������/F��1���i�9�~�מ��A��;�f�E;�L�o�Gx-�@�����<��� w�ހ���� [uϚ���曍�s۔��3sW�����x5��D�0l�+ڡ���'�t�mynĺ���	����������?^S�9Y�xh�!��t %#�<^��>�E\xb~�-*c���[]Z:+�����g~߅ȝO����u���s�z-$����^mj{��*��Ūߛ����M��� ���yI��oNH��R�Z)��G�MQ�Me�}�_l�6������pgdרSϐXB(v��q���O:���I�<K���\�����U#+b�F/�	��z�x��<r��~ F�����e�U�6����wJ�~�-^oOJ�A�}ʏ��C������0�>�ϯ��Dq}�䫤���n��uVL�j<���@~���[�i��� X�wP&���/ Џ<C�V!gR�X6S�����zj�DL������X3�E��myw���r����7CA�^�@���Z��^6*�i�u�lΌ��K���- W (���m$xQ��V~ "�r��<�&D=�o��XBc��CMT#�-��΢�6s���I0�׊0����4O@[9�폳�ȝm�̹%C[�K.�ޥ}ܒ���o��VM�}��4of�x�&��+�֖`8}��z�L��+�l��C�������]WU�7�U���B( ����HI	"@����u�}�׵uI�;�Ֆ� �AX_@����V���.;�-"����X1��IuQ!\���w�<x���@x�����6���Zh�p.)�,?�0���kUt�h������~�{���4�Rm�i���S�����Q�8��X����<*�@�����K
~y��z?~%n�˾�c��8�~�&�7Wl�:�7�q͝�c�z�R����-L�b\
wt�x�W^��ĨpB\v8N:at�"V�3V42`5�k��t�v��������ݑ1x��^����r��:8Qu��i��X}�a��i2s��wc�__��ٰ[��𮬌nif�x��3�e�7�z��	��>|��_��,V|+�?5��Ɉ��?����C�[�����<�����{X����|v�����'����h��+�_�y�V������>�o��s��X�>�������V=ˌmn<�פ7�_}@����������0C�s�:4���4;.b�o��n��%�`V�ߝ�y Q�/��j�W�����{Я*��!����KD	��M#��N�W��L��EWI�asǁ��Wi�Lw��p�y�a������鶌Xpn��<�!�M��:ݭ���x�U�׶ʉ����9%�۝)���b̜:d�M^Zv�#v㴖�8�Z�`�º��#��;�[�z��7v�=K�c�e��"&��U��#�Vm�6�Y�4�;scѣt��t�VX�[WI��ˡƩ}#�KI*���t�c�ޮ��3R�\�Ȓټsܕ�x�]f]/2M�܄D�>ʪ�����m1x�<�.U�8�L=yp��\�v�ڂ�oi�7�ZF��R�>TK
Td�D���[�Ί�zP��y�Z��8�,'Cvܧ���^�#�N�#�5�&((�}���'�C�#f�yu�)}i9�uc�C��2n��Whs �C�}�/TF��$�'F&�]��E�-�,�e��;cƮ8[��#f��Li�*�Y����|-�op�#�J�N��"�v�ky"ӻ����jŗ/xa'�׎L�ҭWtRѬ[�Y`�㹐��$�R������8�f�7A����Q�˱H��:ႂ|�e���`�c�Y6��w�ʳ�7��X'Z<\r$�������NiD�ړ�uq�:|T�B�Jah%q����3	�֜�� �A�zv�s?$v-�M�4պ1�i�	G(0�
�C�&��-�+��'�B���.#9Sŗ��/̐��J�p+Z�*���H[U��!�q^%!���B��M����xa��L��+�:��f=�j���q�u4!�@ХV&�$���c��atE�u������1��<F��+�=�}��thpn�rm�u�쵇��
d�#p1U��$��J�CZ�$H�Ǝ�J���;آ�ɵ5WB���j]�N��4�ۆ�њ�"��1w}��2r�y����&`1��y�"*ک�̝Z��.��D`�4&컖�v��l��V^#'�ڈ�GtV
{7v[�!��zuqhkӥ��'��p`Ь�)��^v�k���ToM�7��|v���V2-ُ���@�8.TK��^�Ig\�qS�]�1��+-�ŀ�Vىv`�=�VJ�H�HV�dv�+���&PW+E��8ԣ;�S|Pp�řlfv�ڥ٣Fb��pD7Ff��# ������j�b�!�]73�C�Q��g�z�^^�2�]����ys�.�#~��ۢX�S1T�v̕٨�2�V �d���EQ���K��QI7�H���$Yr=�9$RH%��������v h��c���>�{�/�ة	Q*�'��$$ Ot�D��2�Q�&���,�w�f@��׷������N�뭺뮺�ۮ�Ӯ��_/oo���~�
�D��!�>�4=�=d}��$"!'��1�P�[$%U1#q������]u��u�]u��]i�_^��q�����}�E��ɕ �HɤT)dE^�s}�I�u�G)�21ǏOoo_\u�]m�]u�^�u֝u����^�>q�!	{�'!>�D$q� �,wL�P��J��_o������\u�]u�]u�^�u֝u�קoo��h���A���Q��uT�"		�5�O��.km�D昤?9�B'ݢ	�Mg�#�ɼ�s�^%%sM��N~��"#���HHy��Si��v���]�R��$XY���Ś�BGƼcs��J�H)JH��:�qj��dQ2i;�:�	a�ЈD�`�b$T�uu��GY#��(@�,IN��L ��a�FT���m���Hj&��GH�L,���FD��(S������$`I�|SiG	��PD(B�-��(�'�a5�5#pę$!��3�K�e!%�=RRECҡ"¢�7�oTH��*<90S`�:6��+���;���	h$���6�h��q�RD
*!��Q'��"e�M�$D'�j-��A�`�I ���[�B�4�
M��NQH�H�E�H^^Oɂ�l�ͺ����w���9�;ڈ�D4�n(�,�!a3$F)�dF�f9F��g�J	�
I&�N5#>q�#L�^F�
Hi3��
/40Fߜ����=� ��[�m1��i�6؁qKi��	b�D�$U�C`|��w}�H3�[|�`����w:�s�w�R�9�B��x����N��x�R�Ѩ�,��,��b�5�&�!�U��e��M��	�}_������O����m����=;�O0`�c�)pep�����{�s�#�z#������ġ	��Zo7��y]<>�r��L^|L�;�<Ԭ�~��:����|n������������d�"�˫ 
�><�^�
ׄ����Ya�f�^q>�{R&w]2���	с����i2��A��mi�Lz�S_9��%۷�Sd;~��Ӥ��Պ��dS
���X_���D�����a��f]���pr�O�t�$�@A�|����nƦ.�7�ٴ��ʟ�\	n��q8���zX5�Y�-y�}�F3�`!��"��C)�:����������\���|+28_������g�N�ocxM�T9�&ͮa{��urt��{��߂�n ����5���ߣCMV�Oi��(��M�L�w�'6�f�j<���2�yB^n����M�~�Cj��f��?W��~P�Ky ?~�o�Dz���-��S���Yݘ��B��lp�0p�J���F{kXT��g���3��~��U���i�X��m'��k?���d��*��Q�pC���p\�Wr������S��|��oqg��u��i\��[ESV,xh��E}q����{_'��x���+���`����z�8,��ǝw���̄���y����)��lB��lK��mR�cm�qFDQ�+<���}����C:|���Og�0Ȯz�rU�N��#� �;�8�t�+��s�,���d��!���b�roC�/U��ɛ��:�H�^1~׬����fo�4��眩 u4����/?�,��{b�v�p�����;�z@`��!�fǇ*)���A�ҩ�M~5�^J=��WK�����j]��5����*�x.`� [xC��4$��pq;ь8ܩ*��������������ˠ�|��-v0yl��m�)��P'��\�����'-���֝��t����.(�fzz�g���|d_��{_���F'�!�f�.u�m: �6����s/[*Vq<��3�;�����<���7�N36�&g�H��ӄJ��o��na�}} O`�]/\�={�ǀ�6����#p�d3h�����t��Yi_Øx�B���	�i�-��������V�Y�\ ��(S��^ }�����J�t`�S�=X}Mu�4�e�k�ם���o�E \@���S��Y���&g�����oÄ��Ұ��s�!l�+�-�F��?c2��t�b+�����7F�*��*�&(�� m�N6�v7eg}�_���"@�$Q���O���oowvEڭ!+r�^ܩ�,JB����XoY��m.	�f���P�m�λd#�x~���6�p! ���h7���h-6��@� ER ��$�6W�v��;��)CǙ��%��Y���[���{Ŀ�"�;�{ c���q�0܅�,nl��z&��jG������"��-Il��)���??�>S�@�e�����!�Kw��~��`֝�=�i�Z��]�s�9]ט�\O�)�k��[��1�E�Td�GJ�su#�x��(8[�?i�o�H����)�4�O=�|w��<�st8�H�T����(�'yp�,� yĿ��?>67��ѭ���H��E7w*���-��^�a�q�f76�Q޳����]m�y� �v8�}mO���7�0hE�cb��P-���8�w�|�5�������+�4�m��2�p�a��
�N$Z�IN��/��P7��ְy%g^r��_!��[�Kh�����8�����4�~�0�&�}8g���V��yw=w���3��"D<I`������(}�U�;���ה��ǎ[7���`��ݯL�n!+�gB�f�3�Z���[Qm������ ~{�T�oP׶1�u����쟘)�hk�Q���������u�]x.Z,���W,q���v�Z��V��묱������k�瘾t\S����Z~�e�i�ԃ&�;]���q´�3e�B�&��������yq�]9�s̬�I?Ƕ>6-�I���`-�6�)M��ĸ
��� �s����������D=�{�>3'���GA�
���!�{U���x��U�6S>x��?����T4*}��T{��e��Ds,x�8O�ߩ��`Cfb�HJ�}=�>|�,_�`�n�C��?��B�;����� 4Ck0j�~����XC/n�.)�l/�ݟ4�^&Y��9��lC�S�Szw������K�}�J���fO�+%@�{*^P}���I����b��+����%�.4ud�Hc�=0j�@3 l-,���1�_:���h���Ϗ�0�5���n'��4b�s ����i�L�RN����?Rׯ�|)�{dw߫�»��sݚW�����z�
�@H���փ�bc�ʇw�;����=2Ԥ�P�A���<�������º�!����fa�y�kw�-�=z�����6�s@�\1�n��[	=��l�6촰'��ۺ�sI@{wY���S����=�/�s�|BO#���K``O����Z�t�=���9��U��h�]�N�i��nS�����zxSH+��a��<�fo4KG�W�}\��n����Qҷf'/��_wj��ۣ�8P��=��4�_*�s�Гm�ܔn֕����d1��G���Б#W��gߊ*�D��W1�w�M�~�&��m_hr;Z�/d:����_rø��lo,�7��\�CT�> x3�>����
6��i�6؃qm�6�ةI�YM�缙��^O^f�*v��oA�vr�I8��Jr����,)�̱1'L\m�fV��e�294�;���_No�X��S�7����g�y� 	��/;�g������d����G8��]���%�$���<�k[w��V�\35xs#� �ķ�
��Z-�5s�al��N��{aY[�y�G�wwww��ֲp��q�͞�û=I8�Y�gwֶ�_?���Ɖ�������=J����<��#���	���KU���|�Dr=�����xn��M�
����`��6��~�S�ؓ�����=^�;ɢ}�V�#�e���֛!eg����c^z%��PC��d`y� 3{�)�24����&/p��=�=�'�@ `���w��A�咀�>�����h�H��K���Ta<Ku�bT��=I�u>7ګߕ���Z����b^g�����7�����~�]�]�q��g|���d�R_zn����١�Թ��~=8.5�D�`!��b9�fX�U���x@8���{�9�|���xW�*�d����%T|��e�J�9��Jl'��1i�ܼ�ܚ��!��ҟ��L�M���Y	���%���$����YE��������rN�+wφi's�����N��f�9�7���m-7�E��	�}سs�=���<��<�Z|�؝�*I!�
��ӏ}�2��Q�l�ۨ���:��v�|�Z�#J�k��i�P��C<���sz��u���	?c���6�ڵ[i�������b�\P�	dd7�{�U����c��=a�ޘ;x7��I����.�.r>"1���9n?�W��[�\�ؒl�2j{oC-pH�����]Xy���4��g��k�h0�=K�b�}��c��5j��m����W�[f����ڬ��6>��� ��mO
V@_����/	c!�~^@����G�n�Č��U.���LS�5�^
�Os��')P�4��������w8�|�<�O�x3p���H�Q$����@U��`S{�����3���|��5���i�ٔ�0���]�O��7�ßƟ��Aos_���Nm���+c��il���@hp#���{~k�/[\��eq�<��݄;,���|?E���y����c}o�)�8�_�彡(,J�v�5ۺ�b6�����C��Kyػ7�p`� (�,!�ѥՉ@O�n;�<�zd�|��Z��4�R�<q��=��KӸ-W���Cy������8���ұ?�����ם��>�����x�ˠ4�ȃ��@??fK^�4ټ��^�{�zJ3g<�z�DԖ�Mob��"���ǟ��u Pъ��*VN��,	�4�>ז"z�'��V�w+^��ڴ�6(!L���w`Ve� �n������q���+j�S��q�-���+>7YpU�C�Ӻ8��<���m�I�����n6�lP��m1�и� ��l��" �����>�~�u�e�U��]ot
����96߱�ѷ�3��A����O�7�3|��]Q��@ߗ�D󬟏��)����;�c�1܄ ?1+��WW�/�;۾�]�y>��t����Å ��_��}.�}X#�1��p���Ә���.I�(S`8pq�Ӯ�g����EG�W�U��/܀�E��T> *�6�;<t�qw�_�?U}��wf���,�Y
Z��a�?�~?���Ob_���M���Qtᤔ�� !�*+��@zu���ǯf���&=��$~��!����pD4�Y_ď��8�Z�*���+�ظ����<x���`"L�A.��O�gѶ�\�'̘.� P��_�$Af�C��}ҭ}M�u�&g#�w����ܟ[�?�[�{�Y��MP�_�]���S?W�-��$8�D`U����ç�ן�7��2H*Ҧ�	���4K�-���p!�ߏE77��9�`o	6�s�����3p�'���i�5N��V���s�O~�������ʜ�-��.�i��挽�ި��-8r�>��$�D�\��2P����mG'N�ND��?d	ЇЀ~C� �
��#�I�#�;77��X�,iD�̹Ϳ,�ݙH�R��K3
��v�X��t�_frΨl���=��������%���Jm��*�lm�Pn(�($����w�~����o��땒D�ɓ������ˤ�xuI�o�O��rt����ØR��i�v�wx�@����u��Y�Q�s����Ν�ҷ	m|Rw-����
�߫���'�~?bu�7cE�`��\�"x6ч��j%�n L�~�C�_���<�@1��J��>���W���[y����]�P��3�1����x�^�g���������/���8f�3��!,G���J�9;����f��v�-ޮ�b�d�|뽆}-����r$nz�6�n�������A�~� ǘrڞ��b�"�����F��ff�SQ�	j��	�XKRl���9�Q�y�����{#�D@y�E]�	���ʪ�K�'��S:��:�k���Y>�ޫ>>��!�l���ɥ����Y����3p����|�Kv=3��~�c�������[��9�D�wz�|��J��Ƽ�T��ޟ���ء��<���3~�
�1�B����#����A3 ��z[�O1�gI��y�ύ�cË��	��8L�V�aa cB��Vy����:���E����B�
��}�הsi����D]j�j��3��7��v�Ds�;Ұv}>��R��+/*��^��)3QM�=ƻ|2	Y��8ڹE�s+d����{�QKWe����&�8>u���.�޶��� ��ءpE���b�i���4�mE�"�*�)"
H�2*H��>� �������8���Ȭ����8��@F��0���;�eݚ-Xx8Aǐ� ��܃E���-��a���f��o�~ݗ��i��^���0���A��i�)�%s�0�`i~�����p'��P��o�V�i^!Ж^^�ߌ������Y�x�-z<H��L�R�_�Û{l��]�i�nfoh�vv������;���]?����lf�>��"�|3�cg�.L��ZrL�d�� z�E���36��>Cw���;.#� Y������k痷��W��[I�:�)=����_�mU��.��x [w��78<� <�N�[�WtD���sOo��k [���M��l1�� ���ȴ`	a���.��{��d�iV���"< L<=��{k��f�ہ02�U��5�zoO��&搖�Kyژ�8oB�w/���9��s��ks���5��xw:�>�i�X뱳;�W^���6��P|�Q S���cf�1��㛧C���I��X?�<�>~,G���ߖ��
���x��/����3d�����ISSYW��P���ہݝ�	ާfk ni�M��;�����2}q��h3�XrF���;N6Mo��b`R����,�Y%*\0�x.��s(���]=9�MM��j��G�j��f8����yy�{�hY�Unϯ효Yϝj���bK�9�1nJ"�!EV�v�.]w����f��U���ú
�)�zc�`%��cm��m��mP���M��\		 �T�	$G���~��~�xs� ~<�5�C��i��Q���&�Z�p���S���IWv�8�5}���D�I��w�|����M���$���-�D�osH�]��'2��39���f��&�Y��G��,EA��P�ށ!�)?�D���@9m��=68|���J��������[������\��]E0؜cs��] �p��l6��z}@��v�5�Y52b�1uO�C�p����=��xT$�Gu��|m`'��5�f�IZ���Nj��`��V;�ۿ��N���TWo�E��>�o���������BΆ�� �cPg煇�����∺ǀ���+���{���L	Vh�|+���6)���I�W�����Ҝ���\I(��XAN�R5�no\��wG�9�o��9��S�m�N�s�C���.�vn|��fo�����cl-���@�[�#ޤo��K߾C��|�%g�Y`&P�[togv*�gv���t���F8�kbӁZ�ݮF��h[��gSӻy�b��	�����*�B�!���nS����%"�G��bە�u���γ˶��u.cva��Uh��,oAX�\�F�� aK���6N�P۹y-|���s��j���f��sD����-�o���uCz��{�&�ے=��"9�D�F��`�}X���V���SwU⎻��X�4���ӽ�7Լ���ƹ\�|{Y��ƞ��`���2
�Ȯ=W3����qVC��J4˺��.�Y�|b\w��BՒևj�C�LV��ӺN�;M��ZM]���z(μ�Z�'�U&U��qוvOV]Y��݀�-���b�r�L��e�"r�A�eu�D�&�M9z0	Q�}}�:�g�E��^#(g&�veou	��u�$��D������gH��)RoF�[�Ș5l�Ny{&E�㎟K_]l����,���]<f�ݣo_uB�����8��j�S���-�c�oK/��kFt6n��.7�d����M6)���-�Yz���;�:�K.�r�l֧q����̍$9���9�d�_&R3���zj%X���;q�۾�r��P��Ƒ�(:G㭻�����qۊ�� H��ܢ0QF���8kqv�]��*��e��)s�#�aSٳ�F�q�UR��b)E7WL��z�˾�(��"֐^A�A���R�m�R�I��E*̀���O��#���Xb���˴B�Y� �՝A�ȢZ@�,����:����c~ߕl����q�Ĩ��C{Ҕr�,�9.�������{�9��ͻ��`��g;n�c&��Kh���M�i��J�w��=��v�[u4��}� �7���\v�h��6f��vٙ�"4�rԺ��I��Bf�E�׽>�Z�+6��]��i�k5;{��%��e;�A\u���{"=�iQ�E0�XFk=��o�k�YW��?���5��EA���|2<�w�����yZ3iC�y�;6�1>�VG������{lk0�8�ެkPp��儛Sp��J�k<D��T����Zor�Ǚ4���[K��.6��r�0h�	�c���}��Ç����k	����˪�5�	�=��]��;.����H�w��&1�>L8�Z���,�%�dA�as��ou������� :��XbY{����9Zɺh��ٺ�,P��̬���c���Й��.}�&j��y]���Ю6̡wB=�u�TR{w���.Z���G�I#�I70^�쎸a�K{��<�~?��>l�DB,B,"$Wd�OW�ň�-�Ic	H��6��ӯ��㮺�:뮺�뮴�>�8���$�9*,x,����b�I�sM<MQ'�T��hċ�����}���:뮺㮺�N�뭺���ӗ���~ϨI��f�����#�#�a�J��6������n�뮸뮺�Ӯ��n���ӏ��x�Bc#U���I��W�o͠�^2E@@�����2Ji�\||u���u�]q�]uק]u��q�ק[x�ֈ �\�*SBm���*��u��D?��h		5���]g�_{=�/͐)Ě"B���"��ग़������[/)�H��E�y���~��K��GݩR�J��J>k�b|M@�H�PU�)�	���6!" TC�$*$,D!W�h5�>.��*�$<I$�&�c���ϵs���;�
G��}�����u#^�v����){-�<��]�;�A����> �i���F6�M�� 
i�����i��H",�H
� ������}o�}��]e]�yE�K{��q�d5C�	@=^��)�{���>����K��Oj�<�4�g�|�o����)�?B��N�Nxƫ�E�r�z������}n�Y��TU�_V�hؼ�v��ü%�&-.������I#�C�>Vy��ە�B�XOy�5O���%������Wo�_K�t�i&'�$�w��8w]��w��{�-��9�n����j��-+s�8ꑑ4e�fC�O��xt��OZ��|Lo������y��ȟ3�a��#�(��<��~���3v�����s�=h�~�������ʃ��04�}�@�,���cMHܞ����[K-$_��N�.M����!S��������[>8�p-8Lt�w�@Z ���K����m����%_�bZ��<��#�Q{�^���K�=5�G�;���ŀ�gT�+��ߐ��_�%�~��]�)�$��S�޿/ܾ g�f�k9
w����~�
z���%��H�v����{P����׻�܆������d��L"��>x|�y��G����x��� ~^\�e����o�_�jy�<ѱ4^�9�fK?K�f.��S'*��\�`h��%�.Ivڳp�N�J��a�*�l#���X5�ٗ����A*͜�|�_b�sC/(��p|�Q�P�^��������H��u�M�\$)��l�"��m6\ $BD�m�� �$�H2 "�"�"� ��w�y��m��ye���a&���Mz|��.c�[�MsG�4z�K ��}�S����hn��w,�P���jkj����I��I`����Od]�������V�~b�a��}����M�Dry73�������r�x�}4�1�[;;� ,�5NBc�I@|�}<�|�Ͱ�[�"f�[�+{=��Q��?'�&Y��y��h�Cs�X.�+���~/l(Z�O�Mӌ���MYӹ�ǯ�{8{�,D���Y�������T{:>���k035qq~ڎ�;z޸��5Uչ��������7=�ߞ��l���J���`�!Ż�p:��wEb�yįx���E��s�n�K��z��y�>�a1���1���>�'��8z�
C&ay���F���z1眮�䶁��^_���+��!���6�����|_��>�L,c��`�oW#��wrDt�k�zشÅo"�L\��n��?7�y������5��h����%��朾�;�{����� p'%�c��v��hO-����]/0y���}Ӻz�ة��J*�T~W���^��ˏm*5ݜQTЭڽ׊����5�rx�x�q	��>�Z�$G@��W��9���d��������yb�Ήu�*:�}̲�W`�����N<�5ot��_w�߇[<����U~	�$@?u��K�4�M��)��lF�4�M��$VDQ$G���;ɾ���wm/���N�{r���F�$�%��������&��ͅ}+�	�M6C����Wӽ*��H���8�~^�G��@��y�!��r�+���4��n�����c键��-��>9��I���|#ɓ��,:�~�rK���O�= &�v��;2;���-���go���v��v�o����Ǐ'%�u�Ö����τ��3������5B�uN^��`0����4 �_C�Ù�W�]�'=�`K��+�8wwͺ�[�ʫp�DD���e�*w��7�_r��&B|��L'2a���%4[��� �y���i]��
r�sx��`:��b�bλ8j�����Of��ݠ0��|,������}�����:HWq�夸|�F9kkgn�S�p0}+�N���t s��WA�!���~�Ѭ��y�E�a��h����/�7x�����5����p.H1�)�����>�#����}�:���ot�p�X8��G���m��l	]�I��w3��|}��g� [��^5�C\�j����hEZ���O/ݰi~�b�П�X�敼�6���xg��/W�po���o��e�G���c��R�'H[��*��'�>1c���	[S>귙f�5-n��l�g���xCG���IT	�xY�@�<�]�ub]&�:č��$�}�Mj�p3X��BS�uj�sz+��Nܱмr�n�]��{O��G��m�-4�M����lT���m6%�YdEVDb�Y�@D���|�|��>���TX���̷�5U����-ͩF��.g
��D=|g`��*�7�*�vz��̚�7�Ͱ�˞L'�@��
����qWP���s�
��늸��	���nyν�7
;䒙+�e'��	��xRv����~��ț�O
��[�CՇ�*�c��bf@���D��*������Ld0�=��pƇ�����t��{�ڥV� j��ģ���Æ���u�/Mr����-\Q��~Y鞯��f6ƌ�c4�w#\@s���uǹ{l-<5?U��B���/!�ޖ��G�ح������6'�dp��:�sh��C3Ws�U���{	��#�1��jʷ	D�^�M���� p=�l!Ϣ���j=�Н��@ީA�p�ٶWX��98���~xnON�F0���W����G�ʀU�O��=��D�x���љB2��v¶OV����C�\�Y�3Ϲw�B��K�����rг��\����H!?U���N�EQ��<��j���c��jW�V�ٱ��֩�/��{��QVS���	���ڭ��%9������*'O�kO��O��s2�WNS�.���(�m���/y�:����QY�n�!M6�`m��A#m��!q�$P	K�9��o�o]pͻ3*���?j���)W1�
6�Ez�%�æ����t���Z�kY	���w���>g�N���u�T.�Otz���	{�m#f��4Z?.�cm�>�u���;�CqzbiÒeg��L��~����]�(:L'۾cτ��
I�v�%���n�<D��������`/��11�瀔z��@sa�;��+zF�3��s!��0��6kN��4�K0n]�ϬC{���;��z9�q�U\�	��P��2��(5�/{�2,��<,=e+ �s��v4 A������1���<DW�Կ\�:}�^f��:£*{�ܪ���Gk��}�ݿ!�E5gL�I<@���^�?h�~7`Ln���/�����ɯVe�D�ێ��)�y�^���z`dY�6P3�!-C�9�f���xT���Vzf�[���XRT�/7N���̿~f���0��a~�w���wP��d�����h��UK��lsb�2��90f������lW��������T;���5T�`�˱��m��T���V�=���o�Lٽ��
�u��y!-���\_n��4s�ٯ�\�"jy�)��\�^x�3wN��vp.;v���gd����X/C-��a���VL�m���;;�?\�{��g�!'��==��	m��. SM��qRD��i� ��H
�*�����������קt~�W� |���V}X$Q��S��~u�MVa�/��{�$w�I��E���oK�;7@k�?7���B?��ʥ��Tl�d^�&���yO$��;3�C���Z��v�jj�1a����T�|���4.���e�VmuE�r;��b��]7����
��]�ϡ��8��	�C�h[F�0�y#��ɳ6=�4@��	��ȟ6�B/v�M<2���W3np,���vj<|�������i���8Ʈx�S��g��(�]��3���[�$����ҡe�n{�E�>��9]F:��d�r ~C����~Z;�����]�q�������]��-i�a�w�]��p|�F���<���=_�C�m���+c�u��m�WSw���r����rcrd�Y^����^�8ty�;��&�s��?��.1�=$�Q�\�9֟��u@?q�fiDt9na�����l���C�n�ùO�p�p��)���ٳ_F
̫���6:�oaW����k��埾�ʸ�Y��|#��Vu�wƐT�xy%� zȳ����Y߲��f�����,��ŗ��r[z��YLM�	�}�X3Q��klMU�cn��Լ������X�$B�m���m6��	Lm���
�(�g�Q7�}���C[β�z���Q '�� ��-3�զ��0�B�Q�n�%5`IS�#�ioB�XoUڠ�e'^�H�t�������`c�.=~�N����=;�8z�O�ՌӰh�Ⱦ73�U�^�${Z8DcBw�)�F�7�s�>{_t�������n\[���f#s�K��<9��v.Za�͘��@n��#�����v�DԵr:Ŧ܃��
�m�)(�����?ry/��~X}O>[�?wsŎ��Wt��Z��{���^��
����~�k@�j�=�0��/�w՘�EM��^��qm���!s �&��Q$��~���З�dP�U~�D�(��b��ۚ}s/�1��Oi�Y���{����!ó�����ڇH6�t��jx�x����5�I�t�ީ^"�B��$���%��)~xd�J��
�OI�d�u���*(�]���{�mRʹ.�;2Qm�m�\�'��~Zj���/M�G�G�~��*E�'S��� �cvnj1�j����׏�;7s0�����O=p��l��@�
|��~��=�ۑ'�?D�C�S8���r$3�F�U�E\m���[�]
�:��f��6�6�ľq��C����nc��'<�\�V�'F
}���ݵ�2;�Wˌʞux��*�G:�V�טά']�� $�i�H�m6!q��i��m7qRA	��	E�������q�n��/�E[���a>3�ȸ�x6<#�e�~5�E
���M�~��۹{����֧�yC33usK>�܋���@aM#��L9�5�k_@)�U[������f��QЎ(���^#��c�����)�5��tz��^a���_#�^�P��:}!�<��j����Zw�s��*<g�ۙO�F=s�6���^Fi����fuf�lڪ=�k���li9��0�h_H���sn9��I��μs8���Xh�P��U�n�N�Ó���6�?l�\��z=�&�7��]?s����t+Y>�a�hő�w���*i�C8A
�]�H~�A�p�+���Z�i�n�R+��@aX��vNt�v��CwoM�H쮟7�y�j��l��Ƹn��5��sL;[܊2Ƕ��	e)����=~<�!O'�ƒg=�����'��8i�Z���������L�q�p���:����,�g�����71���~�<k�Q�RO��^����S��O�6qN��1mVeoe��.�T�cf�
R!���؛ΥK�i�w�!�{��9��"���lUA֑~�!��Q��#�I��u���i!��n�
����TR���[�T��u���]���>�4�
i���SM��1��mn2
� H	"���}���s/.j�i��4��0<[��A�7�qo���L}��*��c�g|�~���/-�ۺϫk&��<�p�L��a*9�T��}*/ߗ�C�^���i@�kcwtr�٨�u2^쑌���.�װLf=�zqf����|�����bˠI�����o*	)��ϸ6�?���q��U�j� >]�!~���$+��Q��kk[�M�)�\��F`��������*N)�\l9��a��������_����x�o=X{��U�Z^~����b�e�����Wv�1������J�k�h�S��U�f�����5�ת���3���C�5E>�ؚ�gz֖��.:�Y3x���1͸�[��f�.��ܕx0�;ݼ0�+LOy�*�f�Oc{�x��n2�D��^�����*�I��ݾ��0�x��u5�kՒ	�q��y��y��pY
`^ϻW��4tVߟv�~hFW�_�m�d�.��"��읕}������a�f�J>�`u��w��C�^a�7#�G���T�o3xȶ�N+�q�����kx_`�d��	��c���P3w���7��3C���30����&�m�3�hwW${��;z����"|	�|R Y�y3��df��B�1��Xn�=�����]\�  +6
�sl�]n�YU]Vs|ޥ���?O��ղ+M6�h\��i���m6d�����5��=��,7���鑡��X:{mc.��b��_�?P���5�咜qg�M\n����r���D�8��V9n*4:�d��0��ei��C�${��[I^M��S�f�O�י�x���͕0�O���FPk�O^��CZ@*<c���db�'c0�խǯ8�F�}f����W��{fk�R�f��n�1��`���>�5_g#�Xw��D��p���T�|��X�C�+,���|�5����>���vӝw;ֵ<��b������4g��z� tw=Kս5��t^�EƲ�TU�_r�f�y���ML�n��dX��>�K�n;k*���>	�=��B�~���w��'�cn���n?�kѡ��������͘D�%�]���.��t��{�p�s���Z	n.Z���8��� �p#~��o�=��HOܳ)zJ��3.��q.A�.���Z��{`[L��<��3�Y$�:�zK��_��s���xxx ܎�㍆!0�ɢ!W;��~*e�Pzz�.sycX��α�Mu��5��N�G�R����8����̃�;�Vl8b�yCe�x�5oж5A8�̈���W*�i8�����N��HeO:�&A��A��T{��{uj{;Zr\��	�U�S3���[��AgY��Gf�'s{Y�J�N��F��+Ņ��A���[Sb�̔�t��q������l�ЭD��:=�ެؙVF�(��Ɲ�)�ʯi���>ǔ��Pܨ"+�ʃn�\'��Ii�3{JЃ�T�U7��ΤA*\(ags:�9��>��ّ�:Dl���\���ݯ'�Z�:~���%�hu�z����Ѯ�&n���B�bs؞6�u�X�a#�◷��,��uBm@C��uz+�7�B�k@ewR���O(>]�(�V">����$,��_�*n�L�[��ި/�gE3<�߆���f��LZL�#MF�s�hm�r��t���ó~p}�tU�u?��1ab�M>)��"U����T�/��G\����B�e,I��n��.�卷�XaH/kP�ĴB^�U�O�˵�Xw��i��Vbe�Ɋ"n4�����%�])mk�iKT�Oƴ�K�Ya�D!i]6�1:*:,�U��!�w�d�s�X��%uW�qj�o�]Q����!��ã��x(�h�LƱ.���<���):��sm#{c�q,��#��2^��k�ۛK']+��(��gs�sA+�1��UL�n���Յ;j�2{�K��)��*Ii�F"���I�ɭc�ۖ�kY�yAY��:hT����9�Ps��H�#xl���Ӽw���,�s6����ƙPUz��mp�	U��Ӈ�a��B���bhs]J}�SP(�҃ӗ�4GJcR��4��j��Qj�z�g`ѧ���"�E���S+���Rݲ̨kQ���R��)�V�`J�\�͛�������B�2��*�;E��YQt�X�qG�pp��֥��9�U�ʠ�V�^�����]L�.Vo'���[MͻUuެ
>�qՈ�vs�6kAd�U���_:����Z�/g0u5܄ގ�>�� �����6���� ��dҝ��Y��<���,XmNb��hM���XNl�N:׻}{�Yud"u�*�Ӄt�i�G�����4�.z����"���$�T���v.�qe`�E�F=�i�Q!B�$$/��>��E_��>k�"
������=>>:�n�뮸뮺�Ӯ��n���ӏ��y��	$�'aRd�X绮�hAQ�ȥ��I	�x�����]u�]zu�]q�]u�q�ק֞>rBHB����y.$ H���L��(��RBI!	uR$q����׏��뮺�Ӯ�뎺뮸�>�>����"R"����zЙ��XXDQT��������_[u�]uק]u�u�]q�}|��_o�Ŋ��iǼ�>钅��}����* �Zyn��&%�	O�}hB"zҗ�"'t����$�O�a_���HLA_�����E �SC����3`BGXO�U �"D|j�DH�Q�1	 
q��g��92"$"ȴ���h�V"Eę ���XDB�-!TK�I�}M!g�
�F8�р�
q%M�ڢ$��^i�dĂ-�".$�1O9�9R8؉)��A/[!�2FÊ�0�(�&%�Ā��$"�M��d��1�
l��%��PDĄD�i�������sױlY��ڊ��(�r�P�k�v��"Ƽv.	m4볤��Op�f&JK��
.E �Co��Ye/$LJF�0�1��L��D2!rC@�!���n0�0 Y@��d)0�%BAj#P�#@��a�ۄ��2�E�[E	!J�H!"R���
 a��S�.$�a�%�@�HM�H14I)FKe"�(@ё���YH8������T�
�q&�2�
���D`D$�h6��6c2H�!�q��|�� �����H��m6���i���i�.,� �Iޝ׾}����u��+�U���L�|&u���\�D�f&�U�[�.��iV֬wb`-%܆�7�o�jZ�q[b�;�/']�:G�.��������|���b"���Cf_ω���I��^\���� ���v���*|��^�}�T���Z<n��K4r��qh*r�Xp�S������=�1M�T�B�����E�\
	墅ǘ��3T@M^��547!����O��5�yS��OL����bP1lt>���K7!�4y�AŴ{���\D�z�,<��^���x��>�Ö�`(�5Pڪ�Q�&�ʁ/C���;=�+ِ�Z��o����٥�ޫ�G{�צS�nQ}.lCd���Z�����U+ͺcL���i��mwaT+�8w�2$py>P~E���H�+�P��W�}���l�3���du/xE�fQ�v[՜!����W�
�W�ܑ^k�,?+���6M�S�o;J^��X`֣9��}9μáC�� �����u�/�c�t酐��:iG���M�Y!��ԏn�ft�$�l9�:�"I2��7�(��[�?��X�[ҏ���w�����M�����W�d�YYYIs	���Ƶ���n�e���F"m�q�N�j��gu��!�t��R
��I�F���P{�ҖN��0�7v���2�=�5���ɖ7��N%koaU���_ƞ�lcm��ƚm��F�m6�I��s���؛�m{���+�6C-~#w� �w�H�_ ]&s؃=�֖~��Ǌ���ӹ��Ǝ<9��P�������ѽ�5̰���/>����U��F��źTU�LKD�g��_��z�;~���ۢ�^���o�=8���8ËNsr��y7��K?Ku<�ƽ���8����'�p:E�N��/|��iXl30�;�#��z���*@����v���N7����Ls
o�Ͷʑ+��\�-��xy�~ynה�&�{���=�mqʡ^܌��C����,~���<�#����M̫9���F&j�"dX];y�ݕJ5��.���P��m`�ś�_�#Ϗm�\yP����h����U�qmp]�@���Ox�4��O������c#�s�Fב�a%�n���U�U������
vge�L��Y)�䉚�;Ϩ\��怔�Ǚ�#�>��y/?�������_���2+�
����B�(׺k�6��&�g:����_���iz�f3�7�&�E;�UP6T�<��z��A�AC��mM��.��%��k0�5~�Z)��_F����N��ɘk.ҵS�,(�[�oVnn��m!�St�%kU����^.|��{���� yz��������M6�dm���B#$�~w����g��۩ aA������{$�?���6�ǁO�����-�^�E+v�`�a�L�t�jw�;Ů߆��G��}�\~��v��~��������{鞞a�eM��'7؁��Hl�D�!��駏�������|�����t�H��L�a����ǰ!�1�O��A'�u��������� �Mr�;������;�wNk��0ýÅ�gs�KU�lezB�O�=^�.{�Lv��fo@I��c>M��l�߮�"n�o�x�
c����k�����!ۓ��izh��E���0oSx��nUG�8SfV���"�J4xd�S.0/���zw�0����D>[��8K}sM��+�7X3���mJޞđ��Ce7�<�7w�X���؅��@���f��� ��9�Ζ��;�x��4��L��d�;+Hr���N�_��݆@5=��h�y��!04�`Χ0�o>�����xx�FDk�+�7�ơ�1��ѧ��P���žŰ�5���������W�݉:XKT��Ar��-׋��Q>7)����
᪰w��J,�'�r�DV��*�]��.��J]
D�a����ɮ�W�봥ˮǁd-o$�=$D�y9��y}!�F����{��������di��l�cm4X�׾����R{���8�C�/S�cy�c�,q��\���Ȋ�-ΨW�0S��ݤ0ɧ�~������N�f��h��(�q,o�7��rt_Z��c���hذ����^�g��m���HE�H�g<�|	g�x ��: q�L'��9k}O��e(ƌ�������O(�Bc�NÙ�P�>g�CY[��~"y-�~�pnW�7�j���r�(����&�aOm����7�gA��W�O ��HXA>�O�}MEN6؊��_vOn����st	R7\N����Mf�Q��V��~g��lrK�4Dv�Kn5���C;�a��a�*���u�l�����Z�x��}��33t�G<��lyjr�Pj���s;?��tX���1'��!#��D�Ϭ��}l�:�{��OHϤfF�kЪ玛���p��N���?1���$C����^y���y,��}�7.`ܥ8��|]S�w�o�W��+/��]&z��+����A|�~]Y�@YA�q�n�މ5}��^R���E��o0��3xȸ�[�̥�{Q�Y]���X��Y$�'b�|ƨ�j�y1O�Y�iӶvm�)�;e��-�W6�,�BQs�d}�tJ]�m�k!5� ������9+�;3/z���ҏ�4�M�1��#m����Ag���:��9�K��q�.ݔ헨e�������k°#Sed�_F�����A�鱚�L��8���h���cLt�e������8���jT�yg��¹�}'��=�mOiP�a���0�ܯ�ȉ���Z]���#�A�x�
�M w{g���i��\8{��@/<��jzRc��=���f���X��or�?	q 4y�-�*=i{��L�>C��z<OD���ݾz��m�����7�m��� a0)��
{h��'����&�]"�z��un����â���bb�INU�A����b«�Ri�W�4>8%��F�_W�_�,%V\��<�>�Sģ;�&޴���>��0�7s	�\8��\�!����CGdv�1��+;�U��y�b(���Ɵ6�e`5D�P%Ty���S�f����:|�� nD���U-}WJﴕ�g<�!�^���ϭI<3i��_榯�5������Aa
�6]��ߗ��%�PZ� �i�P���@��5��L[�\\�L��>��r��~��v�>���uXyݕr ȬH�	r�:�_b#_V���>߻�����/C1��l�fa�� �0�{���=8��T�?]�ouT�<�&{���k�cOl����^:b�v�j�&�7��ިh��@�Iv�e��e��q�(���*��ň8�q󀕭b�V���yF`}�NvWsz� T�qƞ�Z&Z[�V�����6py'^76�gy�7�u��ܙ�uQ��Ǎ?���j�i���i���o~��o�B���-����W�3ey�?6qV�^Y`��l{���K˖�9�*yU�FO&�V\�j�� "ᚋ�:�=�������秽�k#��:q�5��]G��j9"���y�Oč������W�~?E�Ņ`~a��)����v�|�g�y�R{3Q���{�%�k�}����2�^��e�ůE�Vi�W������m ��8O#>�/��Q�켟\�SK��O0��N�f��MZ��6��ɐ��Um�Y�eW���:ط�ɖg�d�{����G�R$c���z)���JF�~�ذ���1gf��p�DEysK�O�&׿�b�ߧ��Χ����Avq9qZ��\#����t���8�3�{��<t���~H���?$f
d?<z'��M�֟k��\M��5N��i%2n���\��5�q���CKV�?x��D�Cҽ<�m��*ݳY[�1{3�O��d�{�;��d�z<[��	��7$H�p�^1�T;wt�>w1có����y�b�����`yx�ò�Y��b>b���R���a�SGޞj�}_b��X��5�q�=���m�C��Z�Se5��L��:�B�Wt�d@A��B�x:�w��ث�����-���i��m��\	s9~���|��ݽ����o�pL�-|�%~�<��=������_C�W�yOLh��۪W`ǒ�3S����"'�CH��s���-��k�9��09���alB�u�C�e��;�+�p�XHknN�8}��vJ�/��4.74��u�=:�>*��ν&��p��p;�2}$P��uV�������ψՏ�϶��874�^D�ۙR�y�5���?Ԇ�J�
���P~Z��5�?7�Ccvz�zEu˞=��ڂw.��=�/~�<=���~��{�	�O�^�:�:��� ;�r#���75t���G�sWi�I�>?K,��G0�d6İ���L�r��?�+<�0�NL���t�g���G�=�}^�Q\�9�n[�tg/��ɷ_�[ZZ��r��XS��\�"�D�
@%�d_��-�}�y#�_n?!S��{� ��/��c|�H  )��gZ��E��p�{��`�`�|/H��O���qB����D��>��~_�H;~�R#��n;�q+�n��]�PMTq<[��bJ�)�z(YO�L�7�U��%��26���B����
�o��p�}�y�f���?<V��h��շ��""n��\4)�(]v�����e,��W{��.�=w~y���蟇�Om7m��m��m������זg�w��7��zW���*P-�����N�<8Gs�T�㿭�		L���|dAi�1qkE>Lj�'x�7���|G����r����;h~���c&���K�C#*��:S}���j����gy����pN9�^yj�һƇ�o����7�Z�A!�o߂���x�������\k�:�6�{'��8�~vng�xx`-��P=�B���q8�u韷KksX�5�ә�����owA����L?4K�W�=z��y�s+��ȁo|�r�ʶw-�ˮ9�Ze;��>P�߼�|��ޘ����x���i�`烯Z�ݮct2���9ʴ�X�����uH5(�f�3��w�A�<�63�	��3*<��O-����͊7'J;�v�q���;���]O^��yhfP����|�*`sw��P�[����bo;�>�����2��{d����'{�i��U�!�r����/b�'��ߎŲ�[Y���ͽ�]-7Eôߔ��N1?��yn�='���^�i-Qyl�>��p�?w�~�K-qh=g[��D�eM $~Ѧ�=����������G`�1ڎo��Վ�4^�:� ��#ú���Q��������xI��*C�!�Jdײ�Q�0�\v)n�,2�`٫:�ήz��N<Mb������]4�MF4�wLm�ۙ^�w_}]u�2����h�ߑ��.L�Q� m�a�ySqri���B�3Z�5�(��#3��Xs���D��e1��QA�@w
����p=�v����4~���n�S)o����U��K��WZG����\qz�25�p��_0x�qOqӽ���3�o@h��X;�f�r�s�zǽ���/g� �,f2|�qR��z=f����q}P)�y��Č�(����W�~�@��k���oɱW���]Pƙ��I;�u���^��hCy�zƿVeσ�9
�����GV���S��U�\3���LH����w�L-�P�=�����w���c~�t��w5`b�;�H�G��_�b�m�9�jk�:"]��Uȿ� }��R;w������4�]V^�w��;��?�@�V�n�C��Tk@���#�&׶C��NIYŤf<w��ܻA��幦:��ᛆ�N��Z��8��U�j��3��ϻ�=�T�	�q5���9�ۭq�n���"qsD�������ƥ��+��C񘆌�$�?~_�k7�C������{����5�����o��0����>�B��:��еRZ�u�Od"P}����p/lp�9OxK?Y��l���~QzTθꔡv*����L�v�G�lcjK��ܠ(��ҏ��� u`D�m�C���y�pɻ�d9կWa<�;�sr�Z�;f��¯��)�y�:�f�Z�.w}˻��~m��m��m���i��HvsqȞ���ֺ`�k�b�R\+�:^{ᘵ����8�S�\��$�����j7�R~NK�>�N7V�Cǵ�'�7`>�e��R�����%=�i,��"d<DK���${��2���P&s�з���u_����*��D��ú�C�~Q�6|����}%�	��SuAy�3=��gϺ�*�7� /u3�<��QȬ�]6�F8`ǌ
���r`��be��Y"1��tS�>��g-n=�����{Z-黶�Y����5§��
��(՟ܙ?,�[��be����w'����&"&��e���G��B������
�8��`n`��%挊B��5��m$x��y������BNmn��G�>�z�g�ސ�<^��\_�ナ��;զp�b5o=N,�Dokp�����c�x�Ϟ�bs�Q��!�)V���L������Wi
y��U��8y)��<47`Ȇ{{��vQ�h���>�m�O����l9��; i=��~�9��'�';��Z�ޫ��v�C��̵v�s��ݚOjh�E�8�;G3C5�eu��+f�0[c�10k]zR��C���F,�(6�B�De������I �Jsb!R�f�}����T�<�����F�j���I�e$4P�h�:�3����6��I�Jrr�fk�LW����Fk6��-U{������F��A��	�6��-s�[zы�f���C�!"Xy�CGrWs5�od�g��/�R!���9cy.��3Bx��J�\Y���/+X5i��B��&������6�̏��rθ����JG��̵�av1���l3j�-3*�_J��M�A�z�]��ؕk���C�J�׿4�2�Q"�{H�C�vR�����ޚ5���w��,ƪb�mI�*7N�rZ�i��tv��j�b�c��q�Y���Lz4K�u��ӧ�-���՛�X;x"Ӣ�s��B�8�x�4^�h-]6�hWY5ֵ��V��������9�ԗa�K&��eT\�ή�荺mk��ļq�mr(˅����{f�yV�*B`0̮ηN�
�ҋ��S�N�}�Շ�_���R\>y��:^u�gI��"*����z��~2r��YǴ��%�vz�R�ZER����^���T:����2�W��7�K�#rX ��.Z�y���%*��v��SD�%�}��9����5�x�^�~�i�ˤ�'�7��a��3����"�mX�,."�ui�.��p���'Cr�.�'w>����l�K
��HOG�:��"��so$�5n��^^�4�]�k��%���4F^3�%�ⱬ�r��,����MK�M�\�
���{9��R)OS��hûVy�"�{���^�26���jRM��_s6^��+��F�h&�ސs�U��t�U�B�Ĥ56˝;305]4��+sxu �MS��M���b�Da�Y����"���;i�+�FC�����N�Y�m�b��ԣλ��7x����ƴ��)G��/�>��9"|��zs�n�Y���A�o��*|{(=�{Kl���;W(`Ӎ�6Y,>R�#sے��S��,^-X�1���f[�v
s����V�}�oI�����ok��an�XCA��ݢp��* &r��@�S"C�J��`軬԰��b���-��=�g��&US���k!�0)�AW���u��3�v�8����m���0�ٗ��R���j'53�NoLq�q�n��wtx��Q0�n�r�5`�_��B,-�a,*D>���*��D�"~��}������:뮺�Ӯ�뎺뮸�>�>���$a��NS[�y%|����Nk2S��R�J^F�R��O�=�����N�뮺�ۮ�ۮ��8�>����9�e�����'�'�4I��e�8�/Rd'd��������D���o�o�>�뮺뮽�뭺뮺�8���<9	<���"q����C��b�2we]���\�3-E���|����__Zu�]u�^�u��u�]q��������=HB �g��Jɖ�d���_v�fL�9����!�h��bө�̹�i		>����ɦ�eX�6�$E����'���4����R��Ҿ����q:���$ERЄ�L�
�X^�RAP�����Rmnq��Y�Es]@�i�����m�"6��Y�"����SU��$�!�aC�}]ٳ�[ޮ�a3HV�̛�<�a�Φ�w�&�gr��������}�����]��O���4�Q�4�m���I�g�ｻ��	�8��>x�L:E����@�f����ނ�u\��{��'=#$�pm3�UZhe1u������z�Q�JOS���Q+����\$?E��4?~y����~C�:��T+�'Q�Z�ŹN�n�]B�.��}kK��31�j���:�\e�s0	���YcY�2vx�#����F3���?WsH�0C����I��v*k�������:�w梾�ݵŴ��N��^�a�S�OL��/~�-��қ�,�/��x�n�N��SQy�{Q�v��>�!�#C@Ʒ�Eq�=>��]J�'�����A�Rb�i�^�������xc���#I��&�7>��5B��e���YS}r��5�q~�v�����w*��<�Ӆ��ѕ�׸��'Lv�)$���K3�}6�{k�� �����B̀�x���Fs�K�*�^$ubþ.��,�u�\�i�����1fo���M4w�h�6!`�w[�\#�.�4'��ZB�-ͷCl�g;�;[]#��*�n�@��D@@�%�!	��͝�A,λ7����7:���{:��"16�RЉv��z:ҋ��r�nǭ������?��m���q��n6�MX2V-���;s��G��7�-�� �|\H`-�8��v�N}BU��`ls�R�9��M�L��)����ڸ��;�ҏ$�F�!��^^E\m���;3�ww�>�.�æ�#C���dh<��¥ޗ��7����Q���FQׂ��]?e���.��\��,/&��}��Qˁ}����x�0>)�\V
�<<V�1�܇�J�;L��C�'�y��g]+I��46����w�J��J���u K�-�=P�QU�K4S�����:sCDd��QL"*j�-ބd���zP�S�K�u��g��,����BuXM=����pn���{�3��i�M�����^�)�)��J�����s�䰨�O�����P���9�'�v���'���z�E�4���:��T����{%��E������8�D�M����{g�j�N�.F=ً�+p��y����8����s?Y����{�cM�ݵK<H�l�!zF�k>��o���i��tՍ�Ϩ�nk銢�Wi�$��6�V�Y�� �k �����'w��Cz��u�y'��n4�t��i�?��*`���Ȋ~���ǉ�±�'-&.�mᐩ$�{մ0��R|��NXGaZSNeѼ�rn�3�!�TwK��v�M��;��l3�O��Z��v{f�!��}#�?�;S/G{�.�Fo�%���l�E^���c�!-�������IS�z��a��~5�Ie¹W�x{��6wJӔP\�ň9��a�|�-j��T�i�º{�4�e�lqJc1e�B�I��ϗz�uz�"UO������B�쑙��A�_"g+�+9f�M�����C|㛄(�wW�U�`k�8�7q�i벥�[��*�Gf��������#!��{B+̣�\���6�0vݹ�������ƺ���K��J��X�u��E�Zx�6e��Ӟl:>��{�^����
-~]�,�rTO*+i�>��Io��<3��4w�B|�z�U����!s�$U��A�[��q�r5����{D�Se*p/�..|�h��/�I����t�Jv~�x���~4����;xwQc-�:Pa�C�6�6��v�3�.�E�������P�Rpj�>����Pp��hoyE.����-C���mɩ���K �Йki�:8bV��8�M��r�@9mJ�M4/�4�MF4��M7p!'}���r��|��� ��U��� 1���)�.�'��]����Cn�o5���Z��i�SO��Y�����n�dr�t޾ �{���tRĢ�f�#7kI9u�j�����Lp�w�'n��z���͗b9���Cu"�l��=��6�{��>����ܫ��2,��rm����z[�n�j�a�x�c#��i�-�Ls�d�!5��͒8E���\�l�v�a9ް��ٮ�b�H�f�v����_�l9^-���p���U:v�E�X;�g��J�9�����t
��t�e_ �]�[�/�{��|e�j���0��:��K�k&�wI�ޭ�\Cc�YT�0��.'fك+�2tv�����!qv�g��2��~��8�1���!�I�C:8偦�d`k8ـ���q�=�:=v�7�&��D�эW�D8!�\��*�p�k�1�BJ=J��n=W-1�
�yh�d<�i����A!��S�=�u��N^r��h�v�kW�s[�u'u�0�	�(]�Ƣ���	����k�ef�p���|i����Q�4�c�����˿E�D�USLMW����0�$��k�.>���/Ͷ� �L7Lj�Q��Q�f���F�PH�l�~�m���RYT0n��N�!+�[ԥ撽���rӁ od�F�l���1��j�&1���F8���VmL����Z�� ΢��2"����G`�vy�1�c��m�n񱞈��@{���)ٙ��]K-����j�q27�<�RҎ�z���o��^k�y�]�ì	�ǒ���4���.��Γ���̬��7%L�7tv��8�gfS�� �^�
��]�v-؇��؊��OwOs{������ƿ���i���{��,7�EI����!>���޽��O!�֓x�9�7
�C�8�2�k	K���'�_DQ=�D��^c�/!�зnw�*���m�������jI0�ZT�Բ��K�7�������U���������̜����讀��.�
}ꮖ{x��IΫԸ��TsY;XD\��N�KR�kk�f�2�<�<+��;��}x��nSM��!m��6�M��$�}�<������wTӟ
7���5�B����X�O��1Y�U�T.�qq�F�^e�'#���νJs��ש��s�1����@=�WX�����7����m��D�g�w�������]�͖9p�>�R�-`��9Hi5�����aAlԾ���w*v�63=��v=[�����ͬ}�ܭH�)a�i�>]-���!�VZ�v
Q�!8|\ibp[���b�|=�|�at.�=(����}��vF����Z��Tt��Za��*�7pрc9�늸��5,�������&u�N$��6˳.\� �=r��Z��*��n�����)�ew���wE��=�5S�hr�H��3��CA��Bܫ\���jP76E�[����nM�������df�aZ�wk�&����]��z��^;��?D�&W7���[4!��y�]f7�C�Q�qdt)��tIĺ�5���Ww50a�ge�C��=�Z;�^e��ͩ����?�h-cm����i��SM���>�[_r��w|&v/�~ˠ�Eܱ-n���FҒ��U�R��]��J��j�����I�b:��!�b��a�n�R	\���֬�!�z~�ffj�מ�|#}i�+1��>Tfo�ӳ�ѷ4����X��77!�5Z�[T�`��*k�-/[.b�f1pss7`fh��o�t���"���2-�4LzG_�Ua(���2+�}Z��8�������~�d����!ʁ9\�)Yx����r����~m�9����*e�)����F3Aۭ����ё*�r���Bt��Է��;�6���wB�� p������T�ɩ�\Rս�}[^]5^R��O)h���35@�g��f�{�x�ofq4|�Y�;!��sa�kp���wePT�aM��c�Z�	��5��JaU�M�4sav���<��p�׾��*ѓ��^:���MSl05u�RFI��޿XZ.n���8��mp�
��T��;�ޢ�X��an�N�
hڷ�K��64�G�yF�w�f|s�GNܭ���2pA��H#l�Z��j�S��s��w3Z�Ӹ�?��ǖg���N��շ1��R��*_����4�Ωѕ���̗�ι%~'��m61��l#m��F�i�<�~�|����|�g������6<j@�g�t7���R{���P�S�W�,�h.X�����񀹼'���xx?&�i���p�םba�T�~��]�1=�����xp >�IC�4���<cCϭ�KUq��x��:t]���'�^�|�e���4f����y��Ȝ���w�[����r����f�p0n�U�}M�B*�����Ñ��i��ĵl�����>oE?U�3��MϖN2�����h
�2'np{�Kx����(�`�b�{_Lp[w;L�M0�v�F{*y�l_
l��~+�q$�ܭ@OI������ YO�7|��Uc-3��Χ���I����/3aSY+�{Ȫf�%��&Ά�'�m�ɲ"���g��ozF�M"�>fn]+&�Q����=�u$��y�B3���b�&���E�>]g8�5]T�ZМ�`���.��-��V&�����$WMt�Wg��X惡�]���=��-=����;�����wr�L�I����y�y�|�i����am��.!�:��}�~�J��%U	E�*����hϾ�-����݇)�!-�̸W��#��Y3�閴݋ۥ��d���Ϫ�`�v�3GQ;^��C)������k�9�J���:�t���\��a�H��������m?���$�;�]J�3�_�g��O�'s�l�ژvx0�{c�{'�m��N�ݍ&��2:���bs-. �g�N��S�W��GO��	���s���A������H8q���*y]�0^��f�������/�+e�q��VS��|ͣ�D��\�6"[��o��7��R!c�1�3,�Ο߽"U|�tU�Цf<��)v)�L�����z�XJ��O7�����3di	�L[��Ҧ�"wm>�}N+k����3���
�ӂL?+���^�G���Y6�������8;G�Ѭb|u�q��l�f��SC]Nϴ7�1ysaW��Stm����0�pT4��^��-��P2u�k��R���
��kd	��/=S�}����6���6�m�nm�;.�_������b�m��[m6���l[Vw]��[��H/��;_��ގ�}�7�'[���o SW�'���cd��&�W�t
�1IX/{<�t�w8��]��� ����ꍳ���Z�I
��<w+>�<晒x�'H`݂Um{��8���G���|�>�7�OW�Qn��wVf%���8
�H�ȶ���y�S�^Y�[Upz��m*ҍez�)}�����>k��8�1�O�����3Q�3�wJ;��z<�{��r���;_�1�����{��4�t�x?rN\gw��&�bAn�/r��^��:tvj������̀��=���W���]XYP��f.�{��}�ƧΌ�[�6sL��6׉~`�I�0����o��A�E�)x�+E`��[��� �}�ڂ�(�i�5�N����8᣼����Ƿ�'t$�a��^87Z�¿qn���hZ�A!�}�՛$vyJ�b��P=�c����@iƅq(_z^�{K_p��dɧ��3~eǱg��7&�3���*hRK5A}�J��g�Xm�2��T�k�ֻ_1��Ml%9K�R�y���G�Ib�Г��b��Z:��w#���A�����$'һ6G�*\TSY"\,��bԞFާ�t�[Fs�$k�&V|��s�չ��G6D�7O+o��蛴Tvi'�۽�r8U.�S��_�F�\D��i�r+)�ܝ����P(K�6އ�L�6�Q,-��U�ַ^u��5���CM[H.�%���^��'Q�#1b��e9�K�wѲ�ņ�&���Ê��˅��V=�Cl-��{Z��
x�n���\�&j%���u��R��3	�lw@��WTac꫘��:'x�´�歖���]�r��X3lr�:�Eg�Af��m4N�G/����;7])9���8�֫�i̍�^@�z��v��2	r���������"W̔a�Y��R�ɏ2.���[��'�Cr���[
�Nb��^�x���MvY��o��T�/��� ��fL��)�!�����H�nG,fBnUzLR�7!T�C&�)$}��IG����0�4�p�]�d�#�PZr�]�(���v��Ԙ$�6�\��5Zu�JW��c�rVS�D�$cm�E�IJ�ȮZv�Ɖ��ʼ�dQ�m�@�hʣ�1"	��}:�l�!W�+��ś�,Vh���W\ї��.�-r<���}r���f�3���N�2�2݃{��[˴;r	�4fu�ȫ�\{1�Q�+�[4!���(��~�H5��e�7)o�;5�t��<�2&�ԬWb糇G`���K�7tv�BE�c�AUހV`ZzP���l�*�*�Uʹ���i���u���z qn����d�CR�e���̣ͼ��7QҾrهc读��J�����)ݑbnN��ӊ�������U{�D����A�Yb�^b�ecӟ.ڎ�nqW�p�ٓ����o�\;C/k�&ȼл=���(}w��o�'�[�R�9-��Z�3�ML=���	�-m�Nj;�-���*���&9�QշUv�ܕH�8&m�{L�\�L����)�M�1���f��Wp֛X�MʸS��]Xu�m]�Vc��lR���Ln�N�#�c�2��'s�[��j7]&^��BÎC.�n����e*=�E2F�Nigc���O���c���ܭ��i�]��*ۊ%��V�=o�S���r3&�MU�J�Id
�קǧ���Ӯ�뮺�뮶뮺�8���<y�r還��K�@���)��$sY��d'��w�]�d�1�ޟ_^:�u�]u�_u�]u�\q�u�x��<��L�#�tH�	8��@#Ɖ�
!
�B%Lq�<}x��]u�]u��]i�]u�q�}9��m����'�.B�c��;{�	�Td�Y�7|m��׏X뮺뮺��:뮺�8㯲�}���/�j�4ɶ�}�Bq�[dLE�ix�"�A~2�7�4�r��n��i�B,�Mv��͠3�&��$z���ʁR�rߜ�BO�Y��t9�B�uO�����u�	$��S����2q
���<ӫųĿS�I	`^�kp��YIp2�, �bm���sL�%�8�X@�}�7�g9����n�w��RMB���>r�$4�Ī�u�l@�PD�m$���1b56sq��x�w�܎p�m���)ȈP�Sm�FAA1�f�+Lwy/�a���;)��Q%#q�Q���4���8]cd=�G��ly|�L{����A�!F�q�"& N6L.�ĺdRD�����LH�M�!�@�&(�DЀ��&@�m"�nHЁ�����
��a�LQzL��(���)S�)��2B��# �M¢�
(�Y ��M8�H�f�e�K,BC`�R���QBh�Bل\@���y:������M6F�i�./3�;�W������V�w:��s4�ɼ9�z��
��ݖ�1#le=�8��ۆ�:�qp⨞����;��0���h�&�Z���� ^��	�OW�V����BktEX��W[���)����.\����]�0� P�/\�&���c?�ǳu#o�[��Y�P%V+�GѰ�&��ю�q�3��iVu�]Cǳ�[�2Z�)���<��'�iξPq|���K��P������ٛ�s-dW����νU�>�uz"(��y���[i���k'3�3j�Mi�1X�lFr�Ec��A�=6v�;iJ�_X]m4�JX���0X�l��n�Z����ǰ�3�6�����oO�$�p�~J�El��t��n�`����G_�!��%�Zh-��7s�35^�2����33��[���H��R[�+l�a�\p\F�=�o�٨�a=������w�ϯ�I�)n�e���:�m�{� ����=�f����sU�|�R'�����H�,��hǂ��@�e�|�F9_	�3J���:ז���߁�=t��{�1�)���JQ��Y՟�A:h鬵3�7\�s:u�f�`��s�%���������6�M�m���m6��{IU�C|3����(���&��S�T��5gX�}�͈1&�uG7�kf�XyΜ�l5�}~�|�Fu��W1YG�<3����|wgf{wB�������+����;�4#��]b�D�pw+,C>���N��r��8�^�do�<8�fR�.H����ؙ����N_k���I}��ޝ�d��fc��H�����ff�fIGI�<4sԳ�u�F(�|��������<�2�p��8T����y�Tį]u�%�罒&�|gʏZ�p���݈�'zm���Ѽ���	��t�`��Ե�f�2�\��`K7��㫙�}��m�e��=Q���O���f����/;�=l��*�I1��X|r�n榟�PAT��	��~��G͔w����xi��׸.*��ƕ8��5�ٺv;bΏݕz�b�T���u�cP�&Ń|�n(�Z&:���ΰ��cS:`�	A;��MRԻ�J�3��b��tS�[�<�{kDγ�o9Y��|i���n��q���G����Y߿~���u0�
C��s�v��D��G���Y �(L�}�rʎBvq��U�#���&=�����SҒ\��x[���
����\�棲��|�t;ڔ	/�˫N��O%۠�"S�U��7�1<�i�:�c��<�!�M���ǏVz��:�W�o9�ȭC7���l��K3������$5��1 e߫��5]=�w��v���/{���MdR�����f7n{{����"b"��]���U9:x�۪��=�O�5�W~�Z�B:��q���67'���Ě�9��۽j6B��b0���)`K'"f##=���w~{�@�>�d~�����'������@�`�{C�EJ�mu6N���o��v�F�>��o�}�.�bP���c��DD�>ie�����קv�d�*Xr�����ハ�(����ēcdJۃ/E��歠<ΐ#�ġ.�z�y����cwJr}:��R�eGՏ3��.�ue� �Ŏ�^%���y�n������Lμ'��?��m4�@@�4�w���\r6�C��3������y��Y�8��w]���Ue^�!E,�~����(#��u��1#�qw:�_����nȨ������w��H?!.;7^�O�y\<��aX���ϼ=���fj۾���v�����A�9Ȝ�8��`x(��9[]�T4XU"��2�&�M��gQ��4��VO�ע�̵]�LB�v�u͆pΚhU��jΊ�Û���A��k����U[��o����кzyr��oY�{ؚ���T�a�HM��3��@�G��>αM�=�=�[�J}��?m��p�HZN]������gwg̤XV�YX����WoN������á��e�#��̡8o^�;ަ���_	�_�k�+��)�+bhl�j��$׮v���ɧ�n���Pч����k�i�[�۞�V� ~��*�L`C��黢��Y��4�&���
�1o4y�A3��vG-����&8�,�����M�'7Fn̥$��Qo�"��7nh`mt�Tr	��dܮ�-��p�������Y�}u%_����M��i�i��<����H�?������G�6$�pH��f�ڃ����Y�}��I�9���RqX�q�S�Wr�u�-�9��C�=\?L��K�6����͖]y����)�;�����!{���\��P�:}�W�gL肫$֗���evf]�/�C�nۅq%7�Wp-Pcӛ��[���HPM^��b+^���GF��$2����w�g�-�dͲ�;\O]���rJ*6�x�N�~Y��&Wޤen*ffëF_����4]�����<�vcg=v����e�����>�P���֋HRj�����gj�k8�H���ӕ�j�J�@^�|v�@��}��/	o���D�U(C���׿�t�b�x��3�fOx��SߓA�\f�e��Z����mv2�i�34��_�CS?��<���0DE(��odo#�ͭ����:K<�T�Ǫ���g'�������qz�&��^=��ND��ږB�0T�Zp�[\�W7�G�}=�u�x��`�93����|w� "	�  �sj�q{k�JN�Cs��u|0�`�b��x�'�>^��x��oas&��+��s�����i�6�M�m��cm���v1wq��F �ޟTdO�ܷ3�}�41����+��^=�Ye�e�"�/p���[<�M�s�f�n޷S�op�@dy��S�?_\�W��M�a��LKSKK�<�/_9qH��Fo��ߛ7ب#�}�԰�it�W���k����朱>�{��R6���p�Gv���>[[t4�j؋�{�O �=?�E��G��o��7ל�����í�C���(�|<�'1���<y׏s
r��7_�	9�3�JǗI���/M��1�:�"""j%���o%UǏ�{����|'��T�g���y{�w$�D���Q�d��
E��փ����fm���'kݬڼ�F�#��6f2	}��4�{%�1���r��N��KyP6���l[���R��N�ޅ��ʙ�����v����u����?<7�\vz�� ٲ��V.^�bo9��e1��&��wuR�w��{��7p],�Ú�G6�y��)x2SȲU�!(�a��%4�d�vpdt_�oW	�[�.&��А��������M���jm�侻�����a{��-���_�v�r���ă�����݃D��x��^��1�V�P��g�Ǽ9�tz�U}�a0�k�~�gj)I�M,��;���7zQ�6��۞yc��p�]�������v"}0ZF�utŅ
jk�x�����\+���*W�;�u怫d�-�u�.�G[���.(��5��TP>�}�Hӛ�j�h��n��]T�/Cr�y�n�y�kw�����S`fn�I��݁+��J�����3�b��f�ʹ���͡��/H|����Ƭ4�nn��wد�H��Mr�U�3xy�y�����"�G7����# >�~;���)���J=�ʹZ��!u-ӂk,k�6�0�"�M���D�X8�Sn�z�Q��-T�����y���ظ�F�K?�'�;4a�7��=[�؎��(�ܫ����,:�{י�i�����a�ޗ����%݊Q�2j�U7��Zj�8��d" ���"!��+�@���`�D��nu�qۻ�`�+{�ÎɄ��q�ⷫ)�g���˙���޳o���憚i��k�?������3�l���w��Ɇ���Q��q9>Y� �<����<�\np��eLE��l���p�;�4� _F�i���gЂ��iSo�w\��l\��`K3<O�@O���u�vo��c�קv#I'��Qt@�����ef�W@ѡ����!��`{F��fk[�FЈ����|}�2IH�����O�����
�d�T�����ke͉�jz��y�V>ͿnZ�4X���I��/�O[�d>;���\Ė�t�UPh��Alˊ��4��PT9 �0)r���kK��ZN�vwlO��f��ځ�v��}9g��º��uN�H����ث�b���h�K�v�}�ݥZȸ
�x��ܳX�[^����k&������%ڨwOQu}0���ك�b�3]37��=㴽�ufu�Tp�5ʻE� ��r֤x�g���jG�D�񺸰��n��ޮi�Q!4R�ә�2�?R<��� vU���_�݌0Ų�޲w'XvO��Ɵ�6�M��hi��_~�4x��Ƀ��Y-��k��ie"
䋍'+p�[�r�h��,}
�sg�b+Mn>�Ȟ�Zfc�b�Qu�H�#���q]O���M��U�m9��H��������q����W)�3SY��7���V�-�k�,������F�o����y�!�q�Ƽ��9og�L��䎃>���Yϒvx�����\#<w��K˶^��r{,��-������^Kk2�;�[\{��3K'l���s5f��1��i�S�߫���{@��z*�udz)�b��M��2�\讜İ�]��qa�eGk⁉��guݔ��ڊ�:uc�Zհ��Ym�>V�ؗ�v�����`�1�Jr5�%�Cmd�Z�㢋���f(�Ʀ���*ڍ]"ż��%����mcl����ҋևwgz+<+�K�u��^��0>�]o7��Nv�GiZHȮ�ff���O��3�m���s��x�JV:����?Oߊ�:SfS�+[�cz�p�%��H �m�n������-|�7�*e}�dS�%x3�����IH{�խj�X+�F�9��Ւ\���%�.��,Q�+,�I�VΧ<���9u��{�.�>}{hi����п�����֪��r}&'�_���T�>E�
�Oer���߲��w]����#�*Q"q=T����^��h�Y�A5�k�f�V�0�If��gg�o>+���8cؼ�^�>��Yyb�7=��>bs�xV��K4��3�=׹��O4�8q/T�@�&��>�L=����N`�K ��{W�wNN�m&S�Ϻ�۠�ċq]�80au�M7-ʊ͸��G�+v���CüG�FT����@j^8�b��\��T�wTPݗ��V������;��/<O]
紹�9=�,���F�&�Kz��Ț�<M���h_O˺k�
8gg�-Ӝ�ws?��M�����GZH vo�B��?LjҪ	�ȿ^0�W��}��R�r6�0r�Vnb932�*��$4��;D�O�y{?~��o)�sYk�8�b�r��2�#��q�;+wE�;�=d�WZJo���\S�U�o�6�ZR4gn�Չ�ꇫ�,6�kz�"{��aB��{����)*/x�)�Q�kn���vK}�u��ޏ7uC�au��������,�cu��Z�":н[�]�M��-�_jMr,��u)�%�p��P�S������9n_>���,b�=���I�劙�[Å����."d�󾮉d��6��WlN��4�h%Oi�\*lvrQ�����/���Hf��*k]Z�R����ٗ�*�����Y�[��ב����z ���Κ�j����"�)"�ǭ��HwCA�Kt�o�5*�ʇFkƹ���Q^�ýo����3�{B$~�mU���T��W^U��%�%r�e(��	b��,���6Ӗ�����;c/gPL���5t��8��Y��������+�m��g�,��Z�-�Y�����[VU�-ХhmL�M��/ƭ��##)[*��5�ⴲ�зC�c�
�t����i3U�2�{/V���݌ە|�r�>3��H�ب�tʹ�c��Ʈ���t��I�yn
�:V:olâ:h�	đ��A$�����͈m-fj`�e��qXܠrзͩT,��/(+F�%B͗���uv��A�Q������.��Vc}�����m��I %�#���~:�e�-m�G�s��G��l�+;���Y�ye��xG���B�Z�m]Κ�؟pz�{q��	�1�h�t�����Ø͹�cooG.w,���ԍ �TՎĖ���`�M�j��w@�s�[�:3lU��ʽW5H�yCG9���_nk�����G<�����Ō��sga�k2���d��B��@z��)p���bc�A�wͼ����;Ž�P�13o~{��,P<�u�^�RL��VT�IoV����ꋮ�YT�^��f���93uB���iuԤ���
(Ŏr��^o'hzT�*��MS�m5?����1�.�Gp��&� 6;b.|m^^
���NWKR���;�5��V,J�'�>���ˤH62��5>{(�w�,0lZ�ڰmq�&��A�e\�X���u��4���\��Mk�z�խS,X��*,PFX�mf8z�]�ۥt�[����Vk���F�k�ϔ�F�pQ�$��9��gl��C�"�l���%��s\d�8\������s�����MՁeج���r(��؇�,>
�5��O�w���#-�~m*����Ԣ$#mǧ_]tu�]u�]|u֝u�]q�q�������Ԓ�B~D��ͬ�}�Lӑ5
�I@��M�����G]u�]u�^:�]u�\q�u�x�D���A$Ou�I�z�N�fI	�I_.� Ƿޟ_]u�]u�]x�u�]q�q����9! �$ɑ�ʞ�żRGt�m��T�ON<{x���뮺뮺��X뮺�8㎾��uG�� �=ח�D���ĳNbBG仼�P��5%,$�Y��$-�\���5X�_���Bz�BunY��j$��
���}L�o,���S��g|I��I�,�k��kg�iHB"D|d�x��K	/b�G5�2JZR"ul����s�vEh���,}b)]��(t$�w�yJ��k�C����W���7�:v;w6�We�������y�|�������������gf��߿r35�[�Q7��+"�z�}]N8G��·Q$���nzP |�ܵȓ��@*I�1��i�
8K33��p�{������˼�{�sh������������Hņ�U7�;���O=	Mc2�]���o��<o=p�<�ށu�x�ȴ��:C�a�Lmn4lod��X�Q�xpwѸۼ�Y����ٞ��f����/v�Lأ�Y<|Ӿ=��~!_��k�h,k�a���Q3���>F�����(�L<La�+(�����gB���rC�u�݃;��Q�
��s�:���J2C���Fh���k�sU)�����Tu���|����t�TL�c��NK�8go+�;�h�*1/jQ	����e.���(O�sci�
i�\�	�'�^�;��"�����%��}}��pԔe�KU�i���נ��-V�\�M1�_䳦귰F�k�'�Z-X��ԝ���唅ouM��7�0u��".��[-=���`�J���X�;�,(�uH�c��^�[��7�;M&^�#�����4��M4���5y������v�zyvT|~�>��gH V�W���2�<�lō����s���kN@��޸5ۅ��ڣ�ďM�)ma=���"^ZL��7�U�i2�xQD�r��o�w��I*{&d�o]���"��b|ڳ��'h	Q����*�I���QܝXAԳ�گ�-��������I`�8��1���tU���77Mn��/{x{���D�ګ����υ�ǳ����/���_+�KF_p[��z}=]���y�[������3JDp�m�ү{	��`<qU �T�
����{s^�ߤV�Iv�U�;�ٺY��P��=6|�O��t�ſ�LF7B���7ret�ᢑ�^d&��/�`8;�+`^<}�^e��\���[�hȡY6�kV��������4ltmӿ�F6�{pث"��,�?��0��PGZ�9"?4Z��q������:�ϖ��K��Ŷ4c\�(*�ByRþi��d�U&f�0�	�;I������WۦTr���/Uf�o.���O�ZJ~���{������m4�mʕ���}�I��y��P��Ş��$����1�eq�;č؄uOR�:<5O(g���i�q.��<��G I��>зf���q>�ÉOy�L��:�����hiqf��Y6t�S޷|ުoZS�C�g�Q7��'"���r0R����mni��νb:*�ʆq�(JP�#�/�N�����΢xlf��AF''6�	�/���f��+�S�M�ԏwvk�^L��&��j�/wT���1P�5SU�N�{����yE3z{z r,SL8�7���뚙�����v}�##Gy8���-� �����8�_\cA��7%V�GA��x(U��ܳ��!$ߛE�&`�g��%\�g'Aי��5i>�&Mk���W.Kw���v�k�oP���_eze���0%�j����yx��V��y�'�����n�Ѥ{���h��x��،ٽ=�<���0]��*^�����j���;���6Z�\��*�~̔����bG�;ھhG��ԡ8EM�Gkm���A��9MVz�H%�����L���Id%P�/;�=�f�{�'�Ņe��h�D��K~��L<�*����u���);��O��Z#m�4�M��i�C��o���5��V�����	3�[�]�������}-:��ia֪�<w1��%��dv�N����YT#WE�k����1���f�ߟ��32ŷ?��_��������8'�>�ކ��p�{s�;\w�i��w��<��I�4�3!��/׏��گ�	���饛�h�9�gD���u�>��ބ3��_�xRUYK�;�9�5�j݉⑛d��3{)ꧨG������vKܾgf�����$�2܅3RD$N#����߷�B��Q���C��/�4�����Y�g1�:�q���[XAp)���4u�e��6�ɝ�:x�/�[��W9^��cǷ ���@���8�37qs�}�����n�o�ϑ���O�j�vy$�NO�ހu0�����~�_����=��|�i!.�j`c*��:�I��"gj)\���h|o�a�q�8�F,KY�-��$�"c��ɼ�R�Ml.M���v.�<U�2W��2v��o:a�U�9��u�����ֆ�i�6�CM4�������uɌ�/N�.��o���"S�[ݑٺ�z}�}ڍ�4�a-�a������+���fé��Y"+��^�� ����Lo?8����[�T̆�����}58��PaN7�{�A���Bay��$�z����Y w
�򐩲�z��,_��ɖV.�ښ�|���-���^��D��؈p��q M�����NN׏���?��o��9�Z����D�;��;۫Vgg%����U��	��$�1��q�·q����Q+��s�R2 P���!�<	�w�����y;��b�޶���$Z'Y�fh7�)o温�<[u��H�@6N���/�_b��o3=�����3�7��t�G����W<���}$2�v��9��*H���p��K�C8��Sjj�Uf'�w��g|��p'�q���O	$��H2a� R����(�#���2������D�B��ٙn��sW��z�#���_�L���7ع��+�ҢI�+Z�ug��mDo��p!��a��^3-�7����̗�����i���#m�4�^�ݻ��K�k	�n��4gٶ���\�����*(v7�� u#�E^Cݼa���sQ��� _e�� �o�[s@?�aX��st�#%MY'{/�0���%�f���?�U�V=���X��8���lw�=x�z�3o��곉���e���GDI~���*z|�\ƃ��ֲZs�_6��#Y�K�����3{D��'�T��r>��4��4�*��SCFV����q�����oxK���n�^�2XC��ޮ;<n�,����z����Y�^��Kķ�"gw�����l�W���ͪ�P9�}�97yK*�t�'���n��
ԳU���������a��y�wX#�Y��E-5��* ��x�s�j�f�3ֵ�D���Z�z殪�M�`E��q'�B�0[��'�7��IҦ��G��e���o�G��V�����'Y�S��d˞���on+�DU�lS������E�&`����|O��+��Y,�H$=y�G���t%Fr]9����;�'ב�|��,_b�ծ��X&]�Q�����6��d����}x��M4�q��
ߦ}>���y�$�6�����YN]�Y5�u۷��^��&�Ε���W՛Ͱ0���9� ӆ�o%Æ���X#���Kߛ���r�oW^dgk'�J��lC���[�u��Ⱦ�<�T`.����b�T�h�46����J:x�ߛ B�:�ђ�� �8V��h�9m��<��`�H�P���@p�1�^˧�2|�,lAUv
)�Yw�
q��JEP1�;�-��ȶ���ޫPJ�oNeo�����n��K�Y��H���׾��7��`^��ݒr���s�!�*Uu��\Ν*�0�2f��>�mZ|��,����8&�g��M��9���֪�쉫g�\{�jDr�V{E]Yu\����}�ot��U�5L� v�[x��{2V����|$�$c��NI]�=]�:2APS���O�R��6��M)�l�\X�p8+n�r���u5ս\�̞ȴ���>ŋ2��Og[.<�]���.O���V��Ѿ�l�ʅ�
;���PU!Ut>���D{H�O/�hf����Wvb���b�p��H꒷za�Jf�aX�T�%Y�[W�[qN���������>m��m���o{������?t+?9�k�O�!�3�;e`+����C���񋈲��t�	�^�^7ϵ��P{�Kotj�v2����'���Y�0��oE���L�ma�Nw��AV�J��m��H+��z����Wl|�O�u
ܹ޻�����ܳkv�/!�:(*�ڷ����St�������3��:|�=�>@*o�Ә�"p������'Mvb�
PdW����y�z)4�E�<u�'�b��mPßWR҈�����;�K�$�U�7���fi��5,�� h�^�	�w*��zv��(���g���<��z��l-ܗ���@���v+3;NP�������������	�	YX��F1����zߔ3�o�y��؇�3T����F�+���,?m_�?�{�<��z��oI@�"�sޓl�i�y;!uw0���.#s	Kv싲ȋNѷ�����!�>���ɲv$��ȫ.�h'(��u����|{5Tԝc�~G�+��F�#�w\ѝ����q��z��@�������?��#IK�w�qe᥃�{22g�0/�7
��y��W���&�9��#*Nn�������M!��-B9�-���K����/��Z�3�>Sܚ�'����v�����5^|��6���q���e��kվ Q��h�,�މH�ܜ�㰰$���>֊��Y��o���.��v�TEx������j�=/�n`O`����m�����倄uA��Ǎ�v�0N�1��Դs�2<�� ���@���g�Gv�헐�)ׯb�n��WXk{��r��p��xS��c⺡j�b����na�7���m���n�
��;��⩳ٮ�ۣ!��8��G;�&h�nƛi���zA(v����/�C�R[�l���p0y�(#;L1�ݩ�cq[������^���k�sR���0��p��װ�0��^o�ý�A��͡0�\�����Ĕ�H����q>}z$#��m�������>�H�!�²nw>��K��\\�8�{ׁ>:�֨fC���;U��IK��@��u�=�=�uג]��=44�CM4�F�i�wߛ��]��_=M�xv�3Sʦ`��3��ӳ���+��g晊��:��nEj�`f^M���6,�z��@���H���Q�c_\��$]h��|�	���j��[xǡv�I��OB�_�o�N�a�c�!�nWbE��B���|���=5�h3�P���`L�#;e�/bP7=p����#���&��Ju��&D��}�Ӆ��������=�i�h��'�NoI*�mܛa�w�>�OEK>�G��:�i��ffoX��)�܁8��B?��6���&������T���ve��$5ؼ��8�k��>���Nя,�}�������<T�-λ{1h��
�v�H� �"��C�"g@}it�i��$�n�K�����ꬼ�H֜T�F��q���X0b.����+�x�K�s<�^���r��r�QU��Wjg��{��y��/Ql\�i��/o68���Z�u���+�������;4��a���	��-�,uV�BsR�S����u�y�.5hu��ɋf1����ں6��m��YFѥ�I�`Xs-Wv��%o%�g# F����yd@f������ų{�ZN�_-篚yde܆�08�C9whi,�[�q=��;�1>1��c������hc���h�P}N�2x=�b�N�|޵�s�����X��8�֣vh)
�i�%a"Y��ά�?.���#��[>�������}8�}r�\t���sק�cW��r�[)�l�K#��'�y�9l��s��)uS2��{el��&&Wgkǝ��w�B��!�B�QSUW��=d*�lW/�F�զ#k���B�9;�l}�f�o��\��m^^�t�JR����%�{�ew�f��%	&���p��K�㪣HM��t+S'.�^�c�T<�̼C����yfml�5��p���Qo�n�\G�E5Ȝ�R��Q�Sw��^*|7�Y���WPF���go������l<N!}�P�,�2��.�޷Ϭ-U4:η�5��6�����Yk�a$���L6�)�͛rڣ*A�dr�v6�&��ɢ�&_J�pc<��Лx�/+�'+�9�0���BҩV���T�&���(36i���l���[��V����)�e�4�	�aԭ>J�sW9 Yw,����޴����㬷�:ua�A��u�*�,�VE9�v�1F�uyԙiv�s�]�^�� �X�ެ����X�c9��'*HET�Gz&�{.��A�뚫JYQ�683}�o�˗R��1j�����ȼq=�ν-�;V�=`v�����^^�+*��=���W��e.\��Y��&�T}��$�E*�����[	��f��c˹��4��xj��P��[�7/њdc�v5R�pW��#���T��B�F���o�V-��}9�N�0%����Է ��m����M��*hc�����$2�;f?:kcz�/.NA��j	df�n�-NZS��u���B��zjά�&_eQ�V��&a)�YFJ�u��ہT�yefGtv�꜎Dnnc�����D��օ�[p�IT��u�P�w�#�N�8$���a��4(/"�����(v���zeu<@��df����v����J���:��u��):rrI�$�tRGrIrN���ͣ|�@��+FkNn��/m���iG�������˦Dʡ�TY*ME��{z{}x�룮�뮺�c���8�:���#�Z��HT��XI�/�㫖���Y���:��>4����������]u�]u�]u�]q�q�׿��D�RI�ۢRK�|���l�m���m�||x����뮺뮺뮎�뮸�8���y�dV�H����h�x�B�I�R�Y���׎=<x����u�]u�]u�G]u�\q�u����	
�@��]�6Y�	nK��K8%��[ڙ4�R�P�!���.�`�Y:�\Y5JK��I�6Q�d%$��Nm	 �H�hD��G�I�uo�9g,!X\��D#k2�0��t[HD�nJO9�I!	'ɟV�P���Bé��K
|؈U&�Q	BB�EdD�9z^Pjz&�!AD��
0�Tj/"$ /͔`L��~��@E��"~���dR�H��i�E���E@T	�p�
E�$�8�3��Q��l�AO""	�Z��G�]�g��B6�c��h��Z5,B�h--������ ���3\��[�*���\���2���2�4I��q3�J1	M8���bQ�6��r�&
�1!�ZeE-~e�M��S����$(ې����!#?2Xb%���b$�M��Q�L$�Q2Ba/��m%��x�'TĢU ���
,�#j5-2R)�M(�a���O�A$����`� AD#�`�cD�Zp҄(b0�.^K�L2��̍�s�צ��W���������ߥ����lcv����8�1�Z0(a��f��Ψ�k�-�b�x莘5�zq��Xsl��O�֤��������c���wcVe�u���<@�1��B�o>�Fcۭ�������������L�/�VD���#g���|��#�}�/"��)n����7�i
�4hk��5�o=U�4���^ʈ0��9��䤈�Y��=񼭥,��Ɛ>P;�qJ[�";}����$���n�C'/��:�H��z�wE(b�����6?�^Ϻ���+�Y�k��M�=,Z;h���[J�$i#'�n��}B2Y�ո��-�.`��6̝P~]���V)��l�C����'%���C}m��u�i���ftu\��Hּ^tb�>F���84`1s�K�I�|�ֳ�_~�Z�D�)�(�w"P���G�����=XT^��Q�ez;�� �X�e��Wf��Gv	0�wK����K�[kž��[�&�h��~/R���!1	�e]�ED_ F�JEET�Fo]�fң	r�Ep�}Q�����z��tM��J�c�nh�;*|���CG1��uf�[�]��F���Ž�c�����3%I��X��i��gW����4��mP��ǽ#��/u�ѱ�~�GU���]ÿr��V��;9@V�ǁ@[ �3�S�����k��$d>��=7;�'�ٗ�}�K!�t�u�4�3��\dq�oUہ�O�4�
��rE��~?�!�+K��ԒO������[l��ڌ��4[��p�vE�Ȋ��\��D�)���Y��љ���fp�`Τ0>镜.j%�+�۸id������{���ݩn���
�ޜ^׌�gs< ����7��������'��0�Z�<�H��>꽧{:��ξ��e0��x̎O._&�8�h���W~`�����gE)��W'�E��e����E�2��u�=�&n ��_��ey����^�E���~��a���0)�.��s1��G<	���A��M�|�:̸��[q�.��a������8B�o#�3�Af�Ss%˥WyRw���~�Ŏ"@��"���0zo��[����*^���[m�H��.v��Qp� �3V�<��:q(_<�;��#L��J�g��|�}��Ag��о�Ngzr�^�D�^��ύZ�`��D�0.`�e�\A��4�,��-4LDf�1{̺}ր��񈺘���2b����1=���JJ�n��A�j�N���?���~�u6�G��[����=2�/Gd��\��۪
%�{3,�ǵm��t��^��¨r��z�5��B��Sֆ�U�fFo$wD�״�i��+�٧�vb^�Ō��<��d�"�0h�/�&7"wp��Pk=ylV�<�P|�����L;�����#:�4�Tw�s""��H>;~V�[N�q�룾v�~�|"��c�kut�,���f��ל��U�f���}o�b�[�ޟl���t.w�'i"�V@5��xL���2]q�u^�3l��>Q�Tk�J�9��&�Ġ��z�ZX���=^�"��,�n�0o{
�0R��U=���}�c�����#��0G���@@�(���q�T�J�U!YFҷ\cF�]�U��H��C�B���9��w}SaR�����_��������<������W�����!�3������ǵ�خW�ik��r�M�N�wa;#��
��Ƚ6�����P`�;a�;Y�Y�$�bG�T�4Ļ��x�'�0�����9;[=>pb2�]�ɚ�N���(��\r��|��蚯j*d��y���|��K73�Gs�O�����Q) g#0G��o����Z��y��w�g�P��Ҳ,Sbޥ��f#;S��̎��\��F��a2!�m�|/�>��瞇��[_�Y�B�)�uF��������A�+��{�7�j���z�0���\�x0v^��Nz'l!�����T�E�^[5�X{Iv��ݸ�d��]�����y��R2n���[�c�3�0�1�+:��z;w�i���\�%\�m����>��ށ}�����[���P�l&f��z�ެu�7�����=��R+�����(����d8�JC��o��!OggG�v���%�JR{/��ڜwXb��)nf�emk��+Q�3\�stIc��|����"�s�|7�����w���g��f$lA����at����^grIڪ��S0�:(�3eL`����J��^�+�2�2�V�^��C&�ef�J��ʃjۈfW(��*:�2�/Y�tܽ�l��Yk�(��vPT��wӯ%������b�X�nyʩa��à?�Lt����:��v�mb��Ӓo�<y�A�|�,ޛt���#�Nq��;BfFl����wlG6�J����a��ng��� d�<�cj�=b<� `��#��E�K�v��Өd���k{�Q���+���7x�yx[U�N%���5[�������+���U��ݕ}K8�g�����(�:;�zKk��wt�����L����T9��J�A鶎궫W}�f|ÔD{{�� M>���P�g��[Kٔ�Ŋ������^%��'��u�!��;ud]��-�~??"G|���(��wP�;����������G<ń��w��3���^�����}/C������h4��/�{Fm�2�_�B�R��ka��.�)���K&�j����ҍxi>#/�U8���CC�7����%���,�U���X:.bH�+�Mm��]��]��W� V�p[���֌r���7���������>a��x;L�ݓ��ҏm�|�0���d�=�����&F\����v�Ւ`�\Lk����"I�Y^�N�ߠ֟7y����M���g,�Z�����f�j8�O�:+�W��V�nm ���;Ղ6�*d�^��!��7Z��67:��;�Ƞ#5HݢmJ��A��I}�Oz����!X�#��_E]��+ʯ����S��I�x27*����&��@8��+~X+��XM
d��$�/����BM�M��-D쪧J*>��O�������kj_�i�}t;}����ĳzc�̙�㜎v&�����Q����`��R4q��2߂����Z����G���'��d��~������礍ب��e���U�dBqk�vz� ��yY�=%٘6^��K1b���ڸj�맞�:bҮ��7n<��ޭ��1�
޸�]�]mQ�o{xNf�1+��桬%Dx>fL@
>J��y�8��dt*n���/�%��8��YZ�U[ �"(�-P���ĸ��;kn����`�c�뮫���w߷��הU���a�����+�3o�ە��X�FL&wgv�眤3���O�Y�w����t����'g��z)�ԧ���X��E�k�O*�����T�:z#�챦�N��6�.���>��Z�g�����[�/净��{�|T���JP&|k�88q�9�Va����� / �@ ��9���N73����X��@�m�qC��zfլ�$~>��kW�J����/ET�ܾឲ�r'�����q�
�a�ތ��a^t+4S��磏U^�Ggڤ�"��N����dڜQ�OAJ���TlG�����\r��2�ss�Xy��x�����m���S���z=SC9.�\k��+)E9�W���Wq��#OJ=��^���z���׿;Y�ܗ�FY����I%�6_[�ͨ�U��d�G?D/8�.��0vH�V(�=ӳ5�3�q�nel@Q�{��6���v���^<��m��	Y���G���v�����=3�R�Ȥ6=i��ra��^ͻ̼�ό1�F�1�w�6��;߾���v���K�m��jNy[����?>X]���X���E*���'f�>��%������)I+m�����Gc2�K�T�=���7�\�{0����+j���W(��ȸ"L�i��̼�u������:T��<{c���r^��=�]�-�Y�Ub�rt0iݺ�KS��nW�,5y��~��\`ӛ��oVrV_�0��i�H��^�ޮ�7��-�W�l����д]e�`��S�مcM�p�:t&ͯY�wW�x���)�+�Zey�� jE��ak_N�"H���*�;��p��2=��p0iO��ԔQ͕J-�%�x?8�9Ԉ���p���cl��0*{N���=���mW����������u�Z���^�|�X�-0���o*1�s��5���A	iZ_��{�M�X�:f6�ţ;���Fgc�����7�8ݚ��wrP(����|vI=U����>�G��z���n�u�$�
3E�[�7]j�^��Z�P�w�w���s�y����~~>�c1c����>����V3��Ի��4��2����ׁ9B�<�vc�!Y��RN��r��M�]�7//w���spE4ˡMV#&a��ꦥ���3��p�_x�����l� ��W��D�h�t��{x��u��çg��z�ߎS�0��X}�G;Ur=���ENI���37ޮ���S�گu��Yl��^�V���^g/�IP~��Yݾ����?�uLyk��Z]Nf�PNw�͗��x�RC��f,��@z՝��9OU�EƳ�+:yj�zՖ��T�\E����t���/����ؼ�h[�5����\K�J��6����p��<�ދ�7Ù���Yz�/u��"�pK�w��ng��c�1�}~���t��mWj�iz�0$I�����/���wg�s�y)�v��-dd���i������', Ӱ�=�k�b;�H��)n׫���q�^z���n_���Ŀ3���{|;8�d��5 ��u�m(����X3��W��\gN��jv�V����6HS^��O�t\²I��S�/X��7]fT��=:]�T�k�䭂	י���������<���=�q��������!��۾@���U�s��L����r֕w���0|��C"����NEO�*~�`g�u�Q�*BK1�v��uH+vA���v��Q�m����`1Ì>q����[0n�*��Tp�P�-�g����4���ޑ���׶:�?Q�]�c���&ZI��:I�j|ٱݛ��d��{l���2��t0����xQ�8��������!�m��o>��g�8�� ��D�f�6���g�x�|$Jj���2���7�gAD��݌{V�<��.e��fj4�)c�Û��0?5�*oa�V��dG� yXꊶ�[��������N���	5�{t��^�lîÖo*�9�}"�}Z62E��/��;����߯"68�r7�#|�k�á�oъ+@#ԈNq3^���T�?9�JNGq�gR8�Z�c����z
(�ή�]������I��%swA��Tl-��3��/�X�Y!��eԪ��7�n���#�܏!kdx����f:6N������]-Ҳ*�%(f5wM�7�U��[
d�����F7�U��"DSr��]�4��̝�o��p��r��b��n�D�	��v
�0����d�" v���ܻ;���[z�IFny�{�h<ۉ
o���]}�n�[�{�c��Ry��ۨ!H�	1���=�Y��u/��!���\[.sxI|�sNr˝�<��k9�Fs���KoM�`��tD�Sg�p�}��k���*���W̛���n�r�BյK��X\�Q����Z
�2�.9#����.�-!�]gl$���J�G��f\i�y��C���X�[%�xRyyZ.�GWd��˶� Ǜ���k鎞��N�}G95��W}񊫙���Kx4�c,�<��hfhx�VЈ�C���P�q�ԣ ��� �JU�9�Z�l �7�1��!"�wC�:��y;��7�2�nP���U�V�,��s���m��ҩ��M�TL��ǂ��]ҕ@l�H�4����r��ީ^Th�
IλPJ4M�*�yr���EU��8Ft���վ�.�q��cc9Q
� ��~�V����e��	�*�iا"�\�MA�*�(�z�@A�]9=A�*b��C�"��rU�^��A;}��74�9�sĒJ9܉��t=l�LSː�e��z�p��K&^��z�XR52�l��w+gWfھT�1�M�׫KSK�:H�b�|��+�I�}���VU�ǽ�Ls]�<O����-㾌Pv����B�U�u����˹�l�jUDC`�:�QάK�Ȼ9������(����[q�����}��Z������FP�l�[�3҄rv�;��34`Col��7]��3;2G��o{���V���⢱�,��X���Ѯ�^�h�q��rܣ���.�*�Үs�:Z��Gբ-���2V��jꦦm��<�M���)�:9���Qn_gs�AM���׵���N(�Eb�����7t���_fR�G���:m�ev�'�h\��ɮJZ�*��K3�^p��K�vM�/Cd,uz���3�X)L���i0fVv���o�sm������pݥ�Uˠ��٘^�^_1.�(6$q��)椒diI!��$Q�$��1)�^�&�yi�mR�yV�����K�	�8p�>G��2�ա�?6XB�W'��]y}z{u����X뮺뮺���]u׷�������>�JREZ*@'Լ��BD	A��!lzq���Ǐ����u�]u�]x�뮺�8㎾������$@�K�S��������u������뮺�u�]q�q����!�Aʧ�R8M�Be9v��=��I�x����������:뮺뮼tu�]u�q�__NIUr��,�}L���lg�'��e����)K9�[�K	'���䓫�9x$��u՝DG6us-��R�w@�#���5 � ��zxɟ�!ż[~%���m)x��;mw���e$�rL�'�{�I�Y��L��3l��ӊXO�&���BH]��h_Yy�&Y��L�k��thˠY���
 �l�%�����z>�9u�Ʃ�Ix�%*9]�
X�}����2T��ū���<2���.��lQ�`��{�o����e�m�K�w��?���wt������>��~���E�p�@���Zn��`���0$�����r	���k��>�6���[�{�&y�F���S{jI�u�;�X�Ѵ��6�2�w��.��n�M`>�F����������=�-؛{YW��h�����sw,�b@��v^��P&|�0čy�t��M��X%��C^�KOܞ��t	��u�՛>����Ơ�zng�����~���|Q5���<s&vr=�Y>����y�>�8:q�}�axޣ�x�Q^6�V,����D��R���|Տ��@�n�nV�ݡF`L��D��x�۶.o���rA!d�p_�Wk��f�����'��!�5w�<?��3�*�*Y�� ���D]:�jɢ�2��a�TI&QX��=��kȜ�,�`|yK���9�fnc��z�{���.�m��=��m��bʩ���=%�����)M�����ƴ��ΦӁi�ޖofm�]�����1����):����{��mʐ��޼���Þ8R��S�j�~����[��l9dE�?ݤ��[���r_M�``��Ǳ�jk�l��cmĿ)�M��W3Ͻq0V�i�C������~�p���20�
���sEt�p�o��v�}йx����Vv0j�S�^G2vs�x� ^�������]%��jPu�ޟS��������璻�l/4�z�=�sy��ɼ�D'��[�?�ezΩݕ!$�}L:���0ڜ�ݴN�d��3�P�o?p�����k�k�{:�;@+��UU��kj��h�.�ՀvI� ϵ��c�����W��?%�G�.ӼFW�3��̬���rul�)�'S����{��� �\1v��dy�ڻ�����7���-S;>��Ė��jygl�<����x�޼���97�o�_)���ς�U��d��-���@���nt��"5�q�5U� i{��&#�6���O�m<����'	 +����Ǎݩ���]3S��,����T���73�{i��7�i)�����麕u��_��������ԇ����h���F�n�_��}��~�\\S��.�q�Ez��Y�"���)����UfK'��)N�b�tJ�/fDܫ��m�����hg��F7a� ���v�B�4��S&�03��=f��E=t���x'���d������|�@��Q�jm5-���pO� ��pއ���Lq��$IN���AM�h��^�YYƬ�&M{<�X0��ky�	g�\_O�X��ba�ҫK�(7ڍۓ32!�F񔃬2=M��ap���:or�3Ruv���9kY��Q���G��^������M��A]��~�R�x�b:z�yV?�s�y�z�|��S�y}l�����"gnr!�\z/��x������A��i`?�t������K �3n؍�Ϟ���%6��W��%�zʼO�;;�ڀ�nC߯��6:z+^�8��;�^JYX�m����D��I�9U���
�<	���8D	^<�:h1�\"�w���ۇ���u���"��
�>��]�4�˒|H�e�/�x��{9Lb����dɍ����� ��7C�CF��˗�Ѣֆ�M�E�۽H��^U���g[!���w
_��?7���k��p�
3��}No��r��:Ƴ���q��K0i����N�,��x�g���I8�8yO�KL�K�E�1�u|6}��)U/u���o�5nap�7z8����c��ķ��)&��(���wO^s��U"C/d���/���q����Q���XK�m�yK�]�C��ܮ�wTl��Qy���u��i��Mz{�{w��4����\�j{���Y��i]t�y�9�p ?��.�˺2���5r��ܸ���ۤ�Ƽ@g欮�W��#��HA�P�fay�&�wy�۽ǎ��Nf&����-������?p��Q�u����扫QZyH1�.�mOU�@�H�L��|�᭳�z1�*�8���VN�$n/?Ww�@�5����?��-�����r���7*���,ѳ�[}�5��N��xl��y�]e�y~g.����W�b�,�,a$?Q�m<�{2�Q�o4�ӑe���Y��b��d����k�+x�Kൎ�dq>������!6���W���|>U���R��Vnn�̆��-��A;U"��2��(���x
%,��g�M,���N��F��t�>�L�q�%A�z���F����;m�T��$�g'�+�-������PAL@n�>��Z����or�/uN��;�[��Rv�=>��E[p�e _��0�����~R�I�w�bETȘ����/�T{���O��x�?N����ױs[v��5����(<�٦{�$A� o��w8�n�`z�D���ӌ���FD��^���W�67X���mПx �/7���z��
�P8^��)�;|[f�"z�E��`��2������㎌EV��{�ȟT[\�l0w(�u�>[��=M��;�[w#��:N�/]��Sz7)��,����q�ͪޔC�6;I�N9�k7��T�J�f�^��\/(�ј��Ș��6a�9����f��8�$.L�:iT�`_��$����	�)#LV�Eϝ�tvf]#�]�)�&;}���'�����c�{���������?U�Y�{t�ݙr &�v�=��|�w��Q�M昽�6x�n0�g_��>�x���{�|`�����@F�-R�CCy��^���!�9�Q��`Ǥ��0"I�g�����{ٸ�[�P{N1�FY�<1����W�R�*<M���g'�{�K��̽$�
:�n���a����ۺ��u}�v��fH���-��G5z.lf:ff�-��ާ�a�����.��*u�V�ۙ�x��6n��$O�x�m���*���S�L�@	�@q�K�W�$�R�5�e-
F���E*�S��m�7rf�c���9y�Vnwif�矗!RV�{˓x�s>��|��P����yp�ߙ���<߯�|��T���G�>�މ^�N��(��IvU��;^�n�{Q�"�������rL�K����1λ��c�s"|6�Rl��~�W�9��X��Η�����z�n��Y���]C��|U�vj֊}�;I��J�	&���TZ;��(��#n�;��­�����y��Wrw}u8J��c��~�`���[�]�S�5lSa��R�.4Iһ�� ����5�v�K��*��w0WAjأC�5�hs��WqhQ�5�t����4\����}�_�h��|���TM{#��ȝ�`ޘ*�^�:�r3��ݫg���p�����}����6����J���o�m��nώ���>�dy��S�ݝ���v��TsWo�QPL
ݟK6��G��y+l��'��㌟�����덨��"���7��k���xP'֧�ܧ�9�#^�B� ���ޚ�=�b��%>^\�C����:��������s�Fɪ�@���7�k��6+W��s8A\��� r'�6NM@q�774����*���d��N?��d�,�)늱e�-����5"3<p2W����p�i�eQ�e�4
�ou�'����<VY��:{���]z=��TDޘ�����6�gB�y�c��3c��񻿆��P���t6�edI�`��=�R����r�mn�|:�R��Cn���B	7x�`�����7�P{�[ٜ)y}���6*���OOk�:��ڝ�G�1�c����~�|��<���V�Gޜ�-�>��ݣ{��k�=Kr��B�H��b0[y�eߟ��s��v$���8|V������ı�-�;�ݿ�b�*�).�:�� :6 >�"eS}o�S�;�׹��U��آ�E�$ָ��׭��.lM4=^�rw��#ӹ�Tɉ����'�v�q+|�.�ٹ~��@Q�0��ۙ�h4�cKU]���ىc�������6�H��>=�
�j}c��L�rRv�Va&��ó���A:(���6�z���k�o=b�Aa[z�f�ئ���r��8m%��9(9z}ݑJ!v�]Җ��Q����/x�k4�[���c�%�C�X�D0�/g��raާ n�fF�c��ۇw��uMʠ�����A����� & 3 �a�;�����?^3Y�V&$o� ���k&�<k��m�l^-nR�;�7��;ԗCYs�|�/�ߪK�H��g���q�I2(Y�<{�|�3u[z;D6֩j���a˂e0�@h���9�i��L��
}���/��>>>>>>!a��IE�Sͱ��U�1�����M����L�b!P���	�`��.�U�o�Ϸ�������	7���
�f:���������������;���S�-��ClG��FV��j���xf�&���ه5-DW�"�����Ǫ�����@:����U/7������{s%��&��ŽT������RЄ�
�����L�%e-"�ꮭv�f�E�[d���{$��+�:�g�oA(U=h�q�4���z�J��wB�8v{<w��sN�`WT �~��Rв�S�����g2ӅH��(}���e6*|;�gw�o�*d��O��8�W�ƕq�[��͛��R&���@���>��u�ˤ�O��wvz�����	Fx9U��5�|�P�@6y
��T���{�a�>m�PA*�F�1N���u�"��p0~�A+�.̬�=���J�Ŧ�x�P��r"C�c��WuS7 ��-!k�&�`͙��0�!������%�B�+��Jy��ϋ��&��Y��ǬN�:���	bA�)xd*`gLv/���y��o7�<�a��;��wF��_9�~���{&�I���`���"�N�egY�u���Fz�Ac����+�z��EU�Qw[i#xÛ:�,�dͣ#��#��/�ǚ��H��T���b�1m�[o�k�^�w��p�ײi���'��#���#�s|wo7>�Cҧލ���{2My�oX޿��ܴ���*��H���Y�7]a�WvHk��������ut{�r��wΖ�5��v4d��E3�Ss��0Fd�����o�î����n��B�U��ۜ9�_=�]=0��ǲ}}w��^o<v��]o��L����)�r���/��
�O�m�S��5�8Z��Wt����c��0#��&^M�nO^Ǹ�!;~1Y8e���F���O?�������ʩ� *��������9�H���
�AE�P(:�Gu�:��2!X b0 1@#"D��@�"P �U ���J�JU�U)V�m�JTU�X���e�RT�X���d�QJ���U�U�d�*@FA������*�*�lTRT�Ő�-�*)R�T�EIe�Y���e�JR������IeTU��UIeR��m�JU�J��m�)QV�*a*A�`�$QJ��ضTTR���*KU,�JJ�إE*�b��d
A����(
���KdY
�ȒT�%%[B HȄD#��H2T#"D�E�T 1D��B2!EBT"��A"0��BH !H 1��BH 1�� !A 1�ʀ%H 0D��H ! H 0��T 0D��HA;��WH 0��HD 1D��HA !HD 1D�� �
 1D��BQ U 0D��BD 0@��B H ! HA 1 ��Q 0��BHT !HP 1D��HE 1D�� H ! H 1��RD 0�� HA !D 1��HQ 1D��RH !H 1P��R 1P��RHT !H�HU2��0D �@�(��@1D � @ U �1P �� mD �P@ E �0A �P2@@ Q �0T�� D Q T  2H2DB � �B 0���H��H1�0P�0�0P�1P�0P�1�@iD�0P�1P�1�0P�1D�1P�A �E �B��Q D    20�D� *�E 1��0`���21A��F��?�u� u�
;���ꊨ��Ȣ��F'�p+��������7�����������?���?���G�<���������?�~��@����������@�$A����`�����O��I�@�?�� 
��/���OM��;��?�� ����+���������?k@D@X"F �� � 	`	@�$@ )D") @"!H�@"���F
Q��DF" ��A�$P`���E"��T��(�H
@��@ ��X�E�$E"	�$ )��(�V �A��U�$b!*�"!E�B
"B ���@"H�@H�
B���H�H ��	(�""����H  TPII@U�$D$@IBQdD$$EAABDT A�!�@�@��"�@�DDB#��@R DBEB DB�C,�����?���~����()"��    ���������g�����������Z��?�џ�~���y��t�� g�a���:?b~
���O���<������!��<?����,E���oB

����(?���<p((?���0��
 X�
��3������������O�]����������3��?�����?�<��t��(������ @U��u�a��q�D�������	A��E��������'���W���>>�)���|�a�_�/�&���@��0(?������������!����e5�o%�m� ?�s2}p$���ꔩ"T"�D���P�!JHE@�

����QT�J�*(J!D�T	 ����R�R�Q$�H��HD�
��R*IB��T��
 T��U�P�*��$	$*�DU%B�IhD�%�"��VFUH�*H�JUJ�T��R�TJ�T%(D�%*)
BEUTR�ETRU�I)I@��J�QU%��R�A"�  ؝@�Z>�w\9�u�m�e�;�v�jT�R�U��SYM+V�k��ۭ:�����J]Cm["�r��M*�hڶ�j��4�m�%	$PJ%R^   �H�U{"-��U.�[��jH�QT��,�mos�VЁ�K�.�2�w�C��6�����Dd���L�n��R�v�Q���uv�S�YZQ�N����T�$R�	RBE   �{&�n��v��]��ۭ";k���ӹ��Q���6���ښ�ͪ�U˶��m\��U�1�wh���]R�5h�$*�"(D�
�x  轔*���@�k-���u֋��fK;�۝Īl��q��W%H�1�5���miN��`ݵu�PZ��pwjR:�H��H�tđU
��  ���ֆq�j��ʻ�UV�Pt�˭f˭��mTv]ѭu�����m�&٥]pw.�U��HV���IV�EEI(��  7�l ��q�:P;�V�h��\ �@�� V�ӎ :���@8�� t5��������D	)"$��D�J�   ��4Pv�th�F  t3�� j-@ t��W@P���9��:R�F`U�v쫅  6�T���AT�H����  c�� ��� ;�`P4�, j�n� ҃t  ;:�@�Ԙ�m�0t :0 �s�RUD�E)J���W�  ��{��c��  ��8� �j�@,P���  nS
����A���*� �@�P(*��*@IPx  �(z0u� t�
 t8��ѵU����p� ��t(P����t� ��U� � �{M&2�J@  Oh�JJ� MxL��4=@ �JT��� �MT�S��  $�JDU@���G��F"Nn�6��L��aE	��jB�B6��G��I�fs����xx{��>���[m�m��[j�����mkm�
�mkm�-�����[V�Z��� {��Ͻ?G����ssW^�4f7Q�k0�F~42��`
���Թ�%�&5�-�B�4�^K�Pպ��L���մ���%�������v������E��iv�ҬEnfisܡ�([ܡ�hEZ���|*�;�{�H���ُt����q�M��=t��J�NӅ��ޥ���a�PᛔCf����d�S8�w�M4�y�7�T�kٍ�U�����I	�"�1�8*(.�f�"nfl��iY���ks ����^�R�"+Ӂ){>�T�:b�	�0$&A�t$盖�m�g-B�X�Im�X�1���I���B[$`j�2�X�4�k�����8�Â0R��n�U��:	@oMډ�f���Jȅ<�D��0K��n9�x���	���B=x�V����N�-Ф��^$>{OZ�/v�ǚ���B[��(E`���o&1�f��iR���
��Pj��ط'�m�qe���5P��"wU�vV�v�����0C�t��V�������
��¨���m#0h�ݤ+^2�7�&���X.R�6�T6�:W�X�b��%�΋�,^�`-X���HQ�+�@p!��Xm���0}�S,�6^^;�[�n�4�I�j�v���P��������ř��
����ۿ�C�p�M�����6<��˹�Yupf�$2X��d�orX���\��c4��fV��Q��j���/ZzvE�����Z���Z��-��Hٴb����V(�V��h�W�Հ���;��x,��2�A��t�2��Ou���;�ѵn�Y��ݢ��ǉu}�mG&Xd�tsV�֠!(���%H�yw5V)�ƴ�M���G�#��i�K���t	`ZW�sDF�S�b���ɍ�`Ґ�j`�����I�����ƶށ�]��T����@�F����.���S݅�� ��)�.=L#uik��བ�pӭ�#s%k��+[v]�n� ���=��N�	�Rjn��7��j�O�z�D��C`���9�����8Y���� ����d�#��0S��U1%d���
{a���][��J�+y̺�L;ե�M�\j�r��k.�T.�%�m�CB	��z"fd��Qu��nPuz�c7>v"Rޭ��2QsUL]�.=JQx�V�X���"�Mn��~(hz*o�Z�ÒñDQT, �b�n��)����mEjRR�t*Wf��+t�I$��ln�Jʽ�jh;�n���5.aiݒv��M�0DRX,�����75�(d*Lm3����1���H�9�,�Ѻ=�] /\�Q0KI�B��K?�wc&([��P��|ԵEn^ላ5E���Q͓2��#j#��y��9&ZY*�2�oH{M*͎�,ɶ�5�m�1�9�-Fb��ZV��G�p�-EA ,<���)ew�~���z&6���И&���0-�	�)���5'jmI/F]Y&R8)1fanG��JtA��ڃ�z~�^���2�dR�u�&���7YwnS�T�Ln��D�/�I��\ϛ�e�C���^��h�:Q�5rX
^�E��n�;4�Wd��4%��Ն�{��OCV�0�b�6�Ba���l�tP��5`�Jj�0X��Nlw(-�ɘfT[�;��`��Knӳ�IkXʶdZ�W� �H��#���ZK��T�p�tm�N�h�V֌,m�eb&���f���4wV[�@�̌d�̫�2VP��A�i8�ule j��oQ����j�4�J�hV��eU�ݪx����
̵��ޡ�Mz��.�e@�����sD�GQ�łn����2ΨØ6�j��+j�n����l�F��9E ZEk�c�Z��Ln�C6�+u"��W��C"Z*ə��42ŕ��.��2n�7Y��C+���%nK%�2��.�`e�p���ۋ1�f���p���.�e]R�aYkM��0�َAv/f������Zv�l���1Z�z��Y�;h[�j<ŷ��sv[*͊�5c��I<�f�Pv�5T�R@mf'�U�Q�tֻ�[z�1�&'u0���ݣ��H����Ă/N�Ȏ�2�Ƭ@��E�T�J�
��!2�TܫHfڽI̳�.�B[I��ò�7˕�VQ�!��Ҳ�u�b�T���J����J��ӴHX%Bٛc*n+.����ݻ&)b�u��;
���Q�0����X�����������/瘭IEJU#��̫���`_ߤ�Ve�:�E��,�^~�
����v:c [M�r�-Z��X�V�Q��C11nU�y-�F���]�X4L����{�4maل��ASÖM�B�X!��ͤ4�kHf�ayf��O�E���(�m32f�8q�,`P��]��PY+(ҧ�kr�TƜl��6Mm5��*եI0^]f'��	,�U�Jv.�^P�YA�R+H��8,��bqcMy�=�u#�S3#�t���$ؼ�V�32�Op��ʼ�SY� �S�yԦ`�mݽ1]	��*KOi ��Ԛf`�U���{S1d�I]���DD�V3$�D�M��Q�"���Vb���gr}>�-�ј�� K�]� :�@���YD�Y� �����!)� ���2oR��Wm��-��9j��F�8P�E�l���5X��4]��GK(
��&lslɂw�֔F�*����Z��w�!O5�K��'b)eB��
��f��Gl<ae�����DS��ɍ|�K���4��Hɔ8u*����P¤
�7fXjY����B��N:�T4�ȣ�̡�AWq�ڄ\#�kPsv]��+ʈ��PB����F̈́�ZL�w&�t��#$۳SQ���^!v�#D2�76��qU�C���I��N*�����)ޓ[�Rc���8ʴ�(��4�h�h�Q��m4���$�WE\�:1�v�8��-m
��R��h��1�*f������R�F�d�S�Pm��嫣��gH�l�F�KU�j�/YgMe�{aC��]�%`5j��58��Ҳ��I�x�#S掽�6� Z���	�ov	�ʵ�n��2"cC�2�Tp�*!�ڹD��t8Z�``�V\�(R��N�^�ma��&�B�[d惖�Ԧ%첊K��a�qL���F�Ӛ�ˁ�5N��
q�-y����I�4
��!'�A�A\�HZ��E	*ɷ�S���P��r%V7(i��D�Z��TMK���.,aY�jj���tf��h[Csmڏ�O���i:�����Y�dѺ���o�!L�L�W�e`���ɘ/1�������4, ]ֺ܃7,@����5J��_j�m1��W�J͐�ɲd+�Y�,{ab"l�Sq��m遫7$-J O*�Y�3�['��#�[
%�N�yw��)R"��ن;�Ӽ�n��۷0���=��y���f*,iz/`�p3�sjG-��U���E,P<�zԷ)�8�o[��YZL�H�ZnAyn]��8�j�KBf�M�ŰZ(���l�i:AGt�+r�!�~Ͷ�ׅ����+!�ސ�a�5���ܳ2�8�8�f�17�]f�n�:{3!y��jixʥ������_"2��E
���2�$CHC�ښ�+��ұ�%��mm���D���*�RN���Unl�\.��p����&إ!k�h�7��VRɔcj�7�V���m��]l�M\�CwQ��	=�{k��y���"�W켛�x@W6��P�Z�-;�c_,�I7��QJ	R�$ܗ��v�kV��+b)c{��@�tK�`� �swU�o)J L5hE��%F
��f�`f�����f]��Otⵖ5J�SĐ�Y
��.&��kn��2��b!�V�V�ed��g׵a7xv �Щ��ݝ
]��U1��|�Ir�ֱ��4��d�2F0%FV3wk.Z�੘�t��Pj��͎��\�	�6�EÑ�Z6�=����T��B�N,��w��h�	�)�Q&�u`�m&��]J"�ղVJ����GPO)s�z��T�����6:��5�݃W���-�VŊ��L%��-WF��4�lE����>[KB�� ���YQ2�tǘ�T��f�`tw�]�� �����6k��[0HĤ���elR1=��U���B��YXv�f�ԗX.��k0MR��^�7w��C��:P9�
d0nD�ʼt����Ϋ���y�LS2�:rJ���X���Y�] ��MxJV#x/��ɺs5�����Ҥ�m��GU��$&>Q�2S��ֱfй�n�5v��M:��=̺f�����<���j�&�)�
�`��2��Ɲk�֚�ޅh�y�d*ayr&����QkkZ����d)���jG�.< ��ޔєif
 �x��VY2]c�����U�-�UA��]Fϊ
̛ZU�v2���d����@<*�]88�uf��OP�!#���-d,a��j+1FHY�*�F�B�v��X�d]�!���i�X��S���
�-�
ߕʻ�!�`��sX4��QCkhe�gd��?����,ҡg�4��E$�x��cfหlͽ��Զ����j��{���j��YB���y�4ݦ	������n,�=r ����n��̚q �-�b$�B*h�`eTА�kpk�ǺAݣAT�X�o1�bejt�f,v�Ր �Ѩ�'ܒ�Pɴ�ٿTƮ[n�)&&!�:σ;fZb�*��2^�1���丞�[p�)=Mm$gj�\��C �j浂n��y'�uya�lJ&��1��_1����tD��x�yz��n����S]�jV�C��,��ԋ�z#H������X�[7��@�&`E��;�r���9��#F�;X�����Rb�u�YT���>��z�V�r��)Z�Wo�HŹ5�5��y2��aGr�k���V�kCbk�B�!@i�Eʙ��^�m�q�4v�lt�a�Bx�4�Kaj��xںDar$P�f؈��aÿ ^�g~�7������nU�P��fl�A��ͅE^�u#
"�[,�^�7�S
`5SP*Bn �
�(3D�Ț��B#2�(7vQ��wZ��f�6⿂�W��ݻ�݁�-��*�޲�5�����j���U�ܬ���~�n��O7jQ�����	�B4�|Fg�K��ʹx�{�G���fŻZ��IF��QYL/b�%!���w�K#�e�[�e���ثL���U�v�&skUL�yz.��0�s	2�V�R&�4`�]Փ#E]^�S@����)�d�YY,Ŵ��J�N�]B�~�p�[*i"�ժ��(�ʛwa�津e^X�o�٘�Wvj��Z���CN�ĞhJ]Y6�o���-ZN���2���ʹ"w�#jL9V�5��l��*���ڃ�2
=`�u`H����ՙm%���57*�)c�q��n:gN�d �-Sx@zS�qMBƝm"�F���`c
eiĮ�*�;�H2�(	�l´'�ަ�� ��ո�w�YܬTC2�ɨ��n:%�YWbK
�o���Y-����B�nf)�]Q������f�!2�n��D�q��K��e�M�2�"3k��21seZ5�2�e��4SW���rػ9��1���V�f�n�8�e�DQ*�6�-�Ad0Bȶ�SQmf+y��jP�71��?&j�f���t�J�+n�O%�e;ͭJ�(��+6^�#ذ�VaK���H�!��+Y�2�Ϸt��ՙe{Dnچ�"��̶�3�9,� @�j�y��[��J��Wii�5��v��Wx��� ,Jj�n�:��]�B��[bV7��Vc۩y*�Qh�M�N��!�*��q�yO��O��;.C�7����xY@V�r����a`�P�wN:Ķ�V;*f+E��\͗Y&K�b��eӫAb�)V��X�q���o5��p���ܦ\����;�� �	�{�]ԱQVw/-b�A��
ٔ��Ƅ �[r�J,��W�bH̩ �%g1-�m�^FbX3F�1]i��S�S &!gc�9GR��Ǵ��{{2��:�F��<@� �t��b�31�!5t�fCh쳛6�%���Va�e̼a�jVba:T�8�,
^h���
Dӽ�h-p*��n�J��̐��[�?%���ar`N�&�m���YF�r�֗�$�dGE+�{�o��kQ��(@ъ��v�Z!m]�vv�ڪ>}��		D�ה͐�Ux2�YA�*��J���)Ķ�`�ފ�k5g� �'I����im�*H�ҶI�ԉ4n��t��i{>�h;�X�F���>A�����a/U�V�o,�J�=�!":�Y,,��(�1Y��ܗ@ɕ�xAn�ڰ2��{��%�i���E����
o%&�vE/��piڸE�c�C&�"�sK�m�����&QV)���\���
�%Rh-UҸ��4��Y;k���u7slvX5$�5�^\kLg���5r�[X�R ���hK�^��X2��-�ڷ�J�a�MIB�6�j]0(pP&�Vnk]kyoͺ{%�J���%�`�LhL-��A)XioኮB8�N$�ݬڈ<E�ˣ3J t¶�O$�R�Z�(ꫤ+l12�.b�]��PU&M���
V��!B�X:�Z~.��#&��k�@�u%���rV�y*:S���T�F�e�Ҁ�M�xE2��mn6������˵^[���ܙl��ǎ��Yv��������ꡩ���JVM��Ll��7+1aĈ�Լ�k�,b(K0ܦ2��!5��:���I�2��h�ikAX�f�-"�Vf��v�G�T�Pm�C��U68V=��+y��VVRP�ٛp;��H�2-Z��RJf���1$&��h����XfK�N�����8ֻOqH�N������
W�p�P�9������n]us=z�@ۙ��H���̭�1��U�d��KN��
�Opt��R.>�nB���G�)\���g6!�拆�隹��,ЇV`\��:��^1N��p 9%c���m6�����,��u�ep[Y}�S����{;}t�WfG�2;>oE�bwi�w&�4��k%��JƑ\�b���]�(���@q�Qe!����U��@�Gm�2�e��;cɈ���S2���>�������M�h.\.�#�1k��R�6�o7�����F�f]��j�2�Bp�3-,F�Ff2jS�ct�s�1�3gEyQܕf�y�W�IӆL8�\m�v�-�!��Ӌ�v��N� �ǒֵX��'�7�l���v՛Mݺ��r
�9�ĳv@�#�,u��\����7�z��x�t����e<j�2�eN�L^�b�m�}���a@���iB/�m�w5Áb�Ţ]b�m���'VH�t������ܖ�s�}ֻMEm�����Cb��:�N�u�TR��{��;�9�S!_r�׌���`������;guo}rQ�C`�-���L^���.��dJ��)(�N�0���{2��A�*�0Nż�XkGM	�v+Ō����<�6��_��0�-��p�+{�mv����m�[�*�Y����e$L_+C��en���L��x^`p�uZ�9�vsN-xV7�(J�Q�Y�v����(���/Q¯����#�87�yk���L�˦�le|��.��e][n���kd^ԼZFSq�WVs�Yܻ��@�Ltq���)K�{ZK���}�A�[,���Zd�F�b�tw:�]��N�"ڻ�Hu��V�V�/XuOB˶�Zy	u�*��T�J��}WZ����qE�6j�ktW*�*u뽦�r(�W�Km����J�ή6ۋ�ˬL�,��k���)aw�s$��'���Ӓ�c�^.f[�%��7�8l���臅�Wx@�w��efPH�<v�}�P׊�>�d-̀v�A�u3�2���Δ�e��K<&eWC��\{`ĺ�K.�{�q�u�n���ѷ�f���5�3����$��aݹ�K����x�cD���iZ6r
�=�E^s��jS����hr�t���F)�絪�ھ�JT�/����F�a`��tr������s�����O
�m�v�X�Ƥ��#���0����ׇP�˗���	�V��B���K��s4��"������]G���xZT�6f�����ɀ���U�S1u�zo��L���l�Vމ���tv!��?�6v�5i��B�M�˝N����o��YK�\�=��
�J�$Y	x��U�2��u-f��f"s�b�]֞��	��n��C�2gRSq�K���/m��3�*|�8�kd��wc���9���Գ�|z�H��	/F�'ۜ���
،�ۻi.f�{)��]���[nju ��V뱥2��bo8�ixo3sQ�*�r�C�Wvi��sw˻@X@|��}-Γ`��YD�nӔ����E�언������o�y���>�5�
��٦��U�uuua��K/Sbr��Y/*m�S��:��}�}�O!��͸DZGZy&���O!��oj����`����T�,�.��di���n����Er�}Ճj�_|�[��/~�ב.p��Y�:���r�j̚�h�'��6q�j�>�[�k!03�=�aրr�멭�V�u��&�p�mF*�_k�V5p@���O6�I+��*c�
�i9[Z�s5��H�7�	�C��G7��X�����#
�eu���;>�!�fc�Z��e.ɒ�W��M�47i:H!Z��jܔ��_1���,]���.lt���U�:�t�㝏�-W֩��uw��u1����︓����O_r�Q:9�;�L1�+a*͝�!XL4����eC}	��;2U���-��������en��e��Ir4�1����1�;Ԝ�b��%1�-��.���w���s9v��y����"����^�������0lm@��.ǯfoe��u\�-m��{+y���*�4^ȍ�5���� j���Qc��Y�|s���b���a"�[�����]IA�A�}�����U��DI���wj��)�i�����wqƜ|�X���/�i=�9t���5�j蛨��D��rc������*n�v��*�������E.آ��[��T���ј�'c���Vs�M�$J��+7QTԨh�p�-�8�P{[�0W!
���Os@�}a�e.é��-E��Q�w�u�Y4�N��&�ε�`1u��܈�!�kpI�&�r�d�p��
�sF��M�]�)�m>����-�x#]�Q�dr��%<�����|�8g�����pm��j�f�����b���.�1d�7P�xw�+w��<����P:m����J��A�j�9����&p�Lsm�x��5' �:�yTu��){�ۃ8Z�Ub9���j��v��܇p�G�>xB����S�-o���Q�-p���1$�n�2��A�Y�0r��:��N�(us{�Ǭ:�we(X�u,N�m��h�Q�]5ڗ]��s�`��M(\2�w�VkfT�W���99�����
�ry�t�yv��e�kU����1��#��cx�w��ǩ�+��3V�Ivuv>����siћjo.\}W`�:�� 	��O`��\�۳ˌ5��PU� �dʳ
|k��k��j)�MȺPZ��n�k
�:U�}�E+�y�L����}���ݬ�Nw'o��Kx��] �#;8�iu���\ɩ�ܝe9�X�V�0\�� έ���B�����Gz��X�	�9f�Nz�zbx�q��Sz�fsZ�һLNm�Z�XK�*w<�n�T�w�1l���Ү�7���볕�r�վ\�^�1DpE�ծ���"��UuʝZ��K"��\v��u��k��@k6������8vТoB�_3Xfw:(�7K����}.��RL��}W����i��˰+fW+g�b7���m���1�r9Qv �[ÎҾq}.��5�c�Z;7����NuG][sj�e�0ޢ,���/i��Y�5ge��N�7ڙB)Mow*>�q*Sl�Ȁ;:��ki�ł\z�6�&.�huȋ�v0:��쎥�0WT�.�;�A�:�E���ZЂ��� �Z��Χ`�w������{j���dyS����߮Il$�,U�h�+��@��u�j�Nm1ꆜK�oD{n�MwWl�����I�0���0�9���E�,��^9�+��V��k���\��ȫ��8#Rv]K�aS�z��uepT�a�܍�u֒������Z����A�oD�u\��朰�ju��.���5��`X��b��B��Nmt��|leq��a�s`�J��\J�7&��N�;|�z��*���$j&�c;�
x�d�:�ء6�Ɍ�"0t��8� xӥ+�|6�'��5��Z����lX�J�8n�ɽ���d����7	-�HYX�U����;�� ��i�|�f�
�����'SC�.)�Fm��f����t!���.P�7�[�7e�P�tM�.ԫ�/_s�ʶU�)B�i30C�S9Aއ,�}sQ���l���R]{N�u킍�Qv��ߎ6�i���LG��hIa'SW3�S�H��;��M*����a��U�QnV�!��)ue�N�fĩ�}��G[��dRwT���[����q�E#�-�+.<�l�)��}�n�ٍ�f�n)�u���Uj�܅���5!�]$��NqB�7c;�a�%�筓}��Ѱ^LJ�yQ{|�܎B��C�aP=|#�2��n� u6�s��4���z�Y][�d�q�Wm�OWU�ȳ�'v�Z��~y��v��r�:tվ�TvN�g��J��$)�x]��n��Q�̫���o���uI�u_���z�&�-opq�a�<�<��9�i9�Le�[�)��S�U{5JA�J�]��4�7�=�;nVq��a�tsD�{G)U*�5C]O(+{z�nӽ�x�'��7�To^+��4}��{ˤ.�vŦ�P�It�����1�yH�Q�Ө�i6;z�/LQ%HJ�0�g@��{m� � -�}X�;P�T�q��sJ(�VwI�+��V��7S��b�gue&�;;�u�<��=�CY����d7�Q��b������r�u���w'���僺�k�� �}r:�L |�m��+/�I�"n���k
5`A�K�,��%s�~�NU8�$�y��B�i��]cr���xr�1C;�ɗ㢏m��j��ڊr[N��/�,�b��U�z<׶����==�Jq1�Ҷ�>j�Z��v�4dtu�;�0�K[���5�+���P���81��d�b\��sm�F�YnY�xM�0��^\��d�1[�O�1��VgPVMuY�Ѿ�(sY�"	ɗQ��q���WL��{�C���YƷ0�������g͆R��E	�W�,ǽQQ� �ڵZ�ě��Y�p�3F��]� �w�u�[:P�|��1�}�հ��=����Mh�nup���5u{��o%�hY�Ǽg1��`�*]�b�](���Ap
���bȚ���#1�P�ĩ\㡕���T��$��)�Jw�y�&�;q�R�5��k����1fn���`s�����z�]�xah-��p3K�;���.L���&�R
F�x�����%.��v.ˬ��c��p̔/�����cM��)^E�u���,妍]��!�J=�b<@Y���th��K�|Qyyt��2u�xI�%��۾<tf�'C#��@T�����iTa!ݻ-V�c�3��g	Q�M�2|n���=���ǉ����3�7`	��R��#��-������i,"����x|9�;	O�;���[�*�����P��WH.e�O%���3S{$�J�$rv�5�$�GRv3�̼�&'` !;!u0f*�p�J��3����T�*贁.��Ŭ�}y1̈́ݪ��Cuܒ�r����7����7Ք7TԤ(��dμ�Mv'�Zz,�"SγEL�P�K7zdw�9I��7�/���q[���s�U�I��7��v�3�)��h�<��\Z��$�,K9��*�X���{Ve#�_g4Ue�ܕݽ��p�Y0em����u�Kw��Ǯ����ϻ5�zB-9gV
?^^YtoE�T�k	/�u��{�ooCsa���a����"6�ά��(+h� �Υn�AtT�y,�)N;�����7���;g��/�t/jx�Ǧo�)�ѬޡN���X+�:N��5����Ա޴���7�>�r�4Ό��
�Cyz󜾫����lnX�j��t2�$Δ+�;N�jwl1n����m��6�6�
U�[�hm�B9K�fEN9Op�m���-�|��k�����+����n�˵����M��+1�WF�ԟD]�x!���j����ů^q�.�4����Fi�i�C�4�9$�UlN�Tu��P�U���պ���Op�Ñ��C���d��T��폦�,�W5{[�)l�������5�U����ʗ&�Ȼ*b�PD(
���; �eP7YF����V=����:)ղ�MG:�W=���M�_F�Ԣ��Y4r���w���AC+3������z߶S�9Zر�2N��❛�0��۫&� K��2Nt��Qm����L�ֈ�M���f�Ҏ�e;�˄W=g'����Ys�����<���a��t�m=�c�Q��T�#�+oo3�Wy�d�o��f�=�x�j� eem�j��a5ԇXQ.zB��@�ᷜ,���[N�L�~��9�g���k��M��	�"��I#}�v�V�]�1u8�u�}\��Գ)wu
"�H�A>*_]�5��Q/�.��M1Ob᥊�2b���!f�_ �kY���7n�ֹ<⹼�[�T%�ի���\D��/�Wnf>��^��p=�Ӊ��쮽�!���o�p\��#嗪gT� ��83j0���9ŉѮ��5Պ�1�j��m}j�y;�����|�S^��h�ǹm����K-���}(����R�=L,S�?l�8�[��Ƿf�S;���� ���u��qYk(]r�׏yu�M���Vd�G�0�ʋ�����r�3����|��0����]m�\(�՛��3q�k	!����������T��tj DT��{y�ђ�j.������b�|���Ϧ.�su#3�V�:�p����oLK�츆{��Q�`d-�X��?Nr�0Tں����'N���^ӵJ�L��?ekˮ��q�ќ_pfQKݮ""�P.:\7Vmf�bU˸�m�G��*�[F��͗�S��m�5w��KUԝ>�+z��I�	�AוX/*ZǢ�igc�3�k���8=��Z'KhgwWT�)i
;�m�fW3�_e&c)A�K�7/x.�O:��	y��2�Eؤ�ĺ.���ͦ��S鱡�@��7��oT]G���X�/
��9�(�{��ޡ2�u�1%���k���w¯���8^��f+[V7�U�:*uX�����4�O@��!ʃ���3n�q�g�q�{._r�v����鹚��xf�����r�WHW.6�8��ɐ۱�:sJ�ǸM��<�P�ᵑr�3)�ZW'
�˺v��S[�ɝί�U��-w�ca�D\��eXc��qH)�zwQ�`�);U�Ne��V�ȹ2��"F��/6.��m�JU�Z��[�[���[��*Z�v���r�ö�����[�RS8��k^ӻ�g�]��V�n-��;�����quJJ8��Ϲ�XTiu�Neo������p�˾�ٓR�1��uʾ�-�ӫ�\�n��^ý@@�A������a�gB�_^菻��+��0�"]��ݾ�H�ˢ�<��s��z�v�{xof�l\��wp����>���J W�;�ǔn����l,�=�@��� �����xx{�ς����*i�o���v4���P�{�����U�� fec�Nن���/�rX+�rTk2�\��:�v��˝���c�� G@,�ˤ���h�QP�)����55�w��EK��1]�͋�1�Ǣ ���G��Aw6�[Cc��l������T���r��>B��u��u��
���Q9c��t�}WQ��;��R�ѳy���ף���^>�E��dׯ�[ie0�C�A5�ޓ`��	�aŚ�͆�Ιx�$���,L�N�_Cv˭Nޟo$n9IV!�N���_Rk%�LK����t�9j^��pOOn��]����j�!/'�Nf��WWC]�ŮȎ��a�ێ*�BZU���dcb��Bs�]D��=)	��L�4��};`t͵:���[�M����:�]��h�� �ԸfY����g1k�U�o���Cf������C]o��[l�B�����������Dʣd-����(��2��H��m��4�LE���fӷi��m�6��uk�I��<(w|��L��4J�X��D>�����N��/�Z��n#V�N_�1�	S�f9��|wL�ڼ���
�W.�u�����_d�&mq1l����S>����{��;���1[��M�|y)4��D�Xc;{aa��
z�C�!�e����ڭ��
���_5�t�4x����p-f(
[.���
Z�Ll��+y�l�83sm꤮��)m�S��*U�MH֑{�Zʸ�x�|�_}0�P�qwZ��\�)a�YD�mM�Yh�b6�;ba��P�D`�Ů+r�院��w�rK�#L��}�c��t�|v�r��{�W��,Ճe����@<RFY�j�(�_�ȍ�̞[�blٳyU��!�\����u�nn���;���9@]�[SWu译�7��f�ph�I�]t��&� �]��E��<�{Y"y�&n��rƺ���-ڧb>�U�ˌ��yo��f��Bh�n\����X��:�G6��Ԇ�M��F<8�ˊ+vv��.8�+��6��lWN���s�SK;�8��m�c^t[a<��"f]_�D�X@˸9
r�m�Y!�[�;�3��L�_ R2T���gVL��;s�륅T�V.����-H��]����R*}�3&�^��"�4�έ�"iQ��G�bX�����6;ժ�QKq�е.-��t�2��Ղ��5��[�g� ��[�:�puիS�q�Tma�[j+�(m�V*���k�͸1����vע>��*e�R��9ۊC��1ϫA��:&�M<6�m�+	4x=���&/]��B��(�T��Al�S~Ɂ)�/�&ͽG�ș���|&�T���p�o�b�Rmj$�p+�kǙJ�tۊ¾*�u5��2�.@��2�_uD��ΨGl�.����h��m:W��K����Pf�������R��
Cٛc:�r�/�卮ήs��᭥�C�L��k��-�w�6�}V�,L��7��$]�$�oQH��*�M�$,>��M �y�A�J���:6y�6��ĝGwe�}]X�G��T����>��ܶ�a����bީ�l'¶Tu�V���'Ht��z���;#8q=	+/��J�MS��]vNVVe�_^6H8~�31���3�,��:"ܱ���o.�{%+5�)��
���{mr<"S�u��ңbH��34󨺝�X��&�mG\/cX�p�F�7&�e�ݤ���-�=,��S�݁
o>ֶ�[}�R� �e�U㌨�)ȴݹo[޾��b��0�V�G� ֍D�*k���K��ǂַ��qT��3|���6gb7�uх+��w[3�}��%��� J�l�݇] �-�]��>�õ�%�G�뎲�"�L5�W��]\����'�l��!��l�N�&ձ�¡��Eq��v�ɴN�^:����Ms�̒V�3y�)��Z�B��gU��]<{�y�,^R��$(+s"�����>�w��
��WH����̶ˮE���e<�-����[�ld�*Jz9K�s�i�3+�$sv��!�̈́X^҇Wg������A�i�8M
���(��yuouu}r9J� ծ�yq6s�D��X]��D����f6>�Z�,��JK5@q>5�n�s�N=�j�; ��ͤ(i�� �ݑr�U�՚����9p*���R�9�VP(ǕҺ�ީ��"N��]M{�_K�{�bvW��vI<�6^K���)�5^s�J�s�YV��S�I�cԺ���J�nW��k��]`&k2�9�����V�M::�쭙WVAC.�,��N(s�R�sQ�����{kCi��2p(�����s�+E� �iMл�v�8ΜGf`TE*x�iͫ+��+�N"�̗�x�\��j�0��Eo-���qI ����8K��]֗0&�)eɖ,v��������4�'���f��5D�7U��J⵺��hT��WZ�N�X�,Yd:�@3��x�:��'L9�,#]X��	;�m�>ͺaL:��Y��o�ޫ��(����.��i�VS;��_^vh���';IX�VK܍�Ij�����ú����ˋ%_X�_
��㕣�7t��+��GL8BM�w����%kt-�w��nA|'Jp@"GmI�gK�����yB¥qҮ�m����"V ���hN��gYɕٛ�,*�v�!:nAۜZ�']�X;����x�`�ve��"��hʹ��ub�;��X �L�\0����4�vkk;f3���Uwa���Fk�]K�7� QǺ��P��ct�˰&¹2�Z���xe���DK�����B;�0���U���&b��W�T�7j�����p���R)k0��η��j^ ���A�P����y��ja)�3�Z�քZ�s���5y]��U����f����S)�+�X\E(n��%����C0YU�5-ѫy?��hw]q��]��)���Tx�>�WV�g(���ى!�rU����֭a�����e��ۧ��:�Чe�y#�l�Q�Aӽ�;^5�U�oH��Am�0�qt�ښL�v.�<r�Ë���Ǳe�����v�d;�s�&N`��ƃ}��b�Ȭ�µ}e�{wC���mi�x��|vf��5�\�(GM=Γ5�<f^��YZ
1�+5��+t0�W��V.��Whkz���"Q����C�������H�:�e)����ɤv���s���:��9T7�R�[��.�q��tU��n�pY@$[��c�t��hW^�=�:�h�N�EG����@l����eM� [�
���W��!{��_�K�1ڻR���i\y�Ob��R��g^�S.w<z�a�[F��7.>OE��h��Aa:3� ���_l�=��v�+�[6�KZ�7o���W:s,�I3+dɹ�J��uav'Ƭ��)�v��uՀԎ��B��.���_��N�x�T�"��!#�Q�*�d�R��irɑ�����|�5/�*�N�T�u�6,���%��۫U�rR�)+��B>�p��D~/,V6/���I,B#*�Rf^}8��З����O����0^`��*X7MѮ��9a�}v)
�Νl`f�T���^�97���
S]�G&���HP�m�8�-u8�}el���Qtw�&l�������.��Z����Ы��g4��;��AmK�nV�-l��Y����m���Rư����nvEDUٜ���A�l�,��G�F
"�pOŬ�ր���m=���7�; Xz��P�tD�khȸ���ņٖ��5cn���B�]	�B������W�r�WK镪E�!A����5u������ͣ� �r�|�8�U��&�j��q<��	���y��aJ�Ͱ�ê�[W|iv��8���r�iG�尦N�'	�vx�Ev݄����v|��5��n��t�c\$[��c�C�H?B��P��}9��Xā`�	Me5l	�:��K�Z�6��Tx�8�ܲ	�&1i���+"��;^+ 8��O�>%�\�iF�^�8A����of5Z��Z#����"�J<~z�
pVl������2��a[NU�o����R��E��$Ǒ�"[t�]�#����ٝ$1�����O�7st�it��8��ex�O6�83��J�H8��6�l�=s"y��)�u�����Xt�)�Sd��СVOg��{���ʛ��\�����Yduq�>��!s�լPO���c��kA=�p���˽�W�Wj�zGc���sv��E
zҹ�R}�����HVYj4�Ո�S�\@	MX�ת��xܜ~ӵ�4F~#2��B��r��ߗk�\wzЃk3��U��#�r�q!#7:�<��r���DR]$�hd[v7/��E�nn8��j �W&xu�LWr��]�BD��~�ܬ� _\��[isv���fno�>¨�5��2������͸�4�t�0�Y��ڗ�}�W+4���نop�loMV��4�xw�aŵ0��.�뚓�������\[*�* 1́\��
'�g���t����p+��`
tY4������	�")l�j�9����pZ7A��@��z�<��%��L��t.kS~�n�����&b�chs������'9I�+ǚ6�VH��y�u���ew
vz2�݈e��������s��jS����{�6[�'VT���3��3��c���y�n���S�_X�J�=���k$t��wg1h�/*�6V��xpoH@A�W0s�N�8TX�s��/��{�W%ٙ�Ե�M������N����pd�Sb/�7B���s��3�����Ƕv�guJ���5��r�G��O�/kh%zˮw(�,�ɫusd̼9o6���#uO#z�D1r\���R�v �b�i����i�@C��Z)��1#$m�1��E@��Uw�*hĶ�V4���8���AI��	h�[�1��3+�`Y�����+i�4�|yų�{��PYu�GsT��b���+5Ga��Jkz���������[U��V�(�h�Z��T�u����]��������n[ي�]:�;u�{u�#`+�T�Qi��?n���+T� �t�X��&9�2Tת��h��궟�঩�x.��Wx�<���4�	wX\���jy�vWweGݰl�Z��0V���a��e%�;,7H�������I�ֻ�7�=f��ݎ�T�VCI��2t��5}Q��W:U�k��ڳx2ХP�P%�g��m�����ٹ��ug{��e���7�V���,�_ WY-ԭ��g5W��nn:,U�,�-E}���2�u�W8bM�����b
��G�V��A��J�Ev�R�_cMhZzi�Ӿ�n��e��2�r����kFj�cN\6�_��9�xx�]|�ì��x�17B^���bP��t��.8�>����sds�.��^������o����3���K!1B���~��ݝ�e���+ �c���ɬMz��S_;��nJ�`��h�I�ν���s�DuKR�?>��
�������M�l]+���3���M�s��p���ނ]ȡ��J�ͺ�Z�Y[c�hY����h=�&PxH஝�Cxl�M��!h����|HRp��Ya��0��רlw���m �۵�h�N����5��N۳�K�
��p��aw2+"�ҳ�$VM5�ij��RڔV��Y-�8��lcadݔ8���P���K ]��@��up�;�E�$'K9�\���8X8�Y]r�v�4ɮڼ�;��:��G�����n����b�Z�=�mV��P��(�c��dY̊e��wV�6�0q���su�m��al�˽V>N��kP��s �'�����N�M$�
%��C��^�6�3jDƷW"�fk\�uݝ��%d�ѻ�]v�
d�i�X�<h�0�GDWIT�U�l��t1���kb��
o�qX�� j���s7u(4�����A�)�@��n.b-�W;a��y��u���\�]�����˕��v�;�����d��:3��dY�=���Y�(�6�w���f>=E����Ip�xNC��:�Y�Nu���˱���z78-2^Yhw.��e��b2�۩�*�%��˷v��Sn�j̊q�1Yyi-��x-�6T�)��m�y�Y�ɐQ=׉�ɚ��U.�⩮��h�L���N`Wb�Ө@��9�1+,�Uc��J\ќ�m�O�j^�b=���h&�
�@�-�oE�	�0�mWVb	�NӢu��:e�h܈kb��VJ���R)�*��Yv��Ż�G�zwe�A>�ӷ�DU#�xD�)f.��;sBA�I�Z��gQ�ɤ��:����ٮ��j�	{�n����lw+��9ZzB)ۦ��\ۭ�s�P����,�6��{	TN�(9]�y�$ȴ�(����Kf���-Ln����c�T�G��^�	�~�|&�S��.��5����U���CUL1��~y{�ź��Y���\�D;��{�xT��wƆ����
����'j�e�D.�5�k�OzFeZ`���N�\�]��>��l�o��Bqi�����V��E�ʜ��y�S�r�G�z��ט�%�JْD;#�7�䂷�.:|6��z�u���c=Gv����Io']ҟ2G:���d;K>�ZQ���n��F�;1)2�_;�{�0�d9<��.�YS2�K2���=��p�+A�]ӱR��&�}�)�)ٝo,�y9N�j�_e�^ ��2�r}���{7�^g6�]�CQ ��;�3o�)���9�d,w@k'h.�e��*�� �@����5Kv��������ܩNHܻ���53 �h�����rv+vj���p�ڏFL�_@4�x1޲A|'޷z�U�1�>2�o��r�밷��͟j�2���Ef�u	��[��i�u�>�O댬���U_{���������n�c�:�xr��.Q���8��iv�Eh���𸳸wU�㹮��AT����!��p�j�������Fb��F@���\Kk���jK��xkQ����o�5�IDe9CtY���#�5y��-ˡ�֛|�c���]�5���h:��\1����0-�1�T��ʨ2˄}�,����
�!ʋ!pZ��ۏ��N��tR���ҷ��VV��a@��y��P�h�'9���ɱ���"���"��T��c!<��}���o��`Kmr����z�t4���R�I��
�,��4oZ�N��і(V��o�WKK���(�.Y��w4�Ewl S���;^�(�V���7-���Wi����}D�H�� ��:fc]O�[�����l<�d>�{�5W�V�:r&fb���������FB��mtђŚsy�.��Lm��j��WU��s���8�1ptJ���)ڱ��R�x:��[�iB���{"�XEώ�#C�h�j��=ם*����<Yɺ"�L���`<0a���y{)sm)u�ՋU��Lh��Τ�
��wqE#Ջ�����r�`uv�e^�;�$�:�R����(����1q��|q]�M;�	�L�P���y���dc����' �*�pO�O1��s�;�Q�;���	v�r�7���e�ne�����P!s�����������{˝`1��q�q��sE��Qs��t^5�"ɮnwnwwu� �7d�2�s�q�HW-�'.I[��sWK�.�p�滺���5�w�����ݹ�)�����F�ˎ�&1�w,�N�d<����^9�guݺep���η;�.�<W�n�G.��ӹ��E���y��&����I�i����	�nҹn�5�����RA��ɜ뻆Q�.�o
+���;�.b����o��sk���뤈�5���M<밋o�t�]���+��j2&L�����wTU���mI�U   W�QU�}�����S�O+�����ueU��!�]V�N�w��ǡ�tQ�8٢t�uv�Vd�ر.����nT<�u��0��vE�NA��}�<f"���`gq�ժ�n}h��S"!Y�����^�J�/gD�^�j��I���i��@o �Nϡ�$�����=��+,Wexu��*j�-s��]E�LF�`qq1y����Y�	�>RY�g�n���7�6E��P���*��+��j���,V0��8��4&1h\TV<FJg�!�W�:V�fm�c�]||�ΓvG`��(t�ǐ�k�1�g�ʌ�f��W<BF`ŶEM�tĔ<��ӳ/��i���A	4�Xt�x<�S�oJ�:�n|�f����]���,%�wZk{�����MY=��?�>K�&l �\��J��
W��Y�)j�4Ǯ��;�}��1���X{�������}l�	���BHZT].2�b�5oF�\�:]#��!j��}��w��zܮZ�ϗ"+Χ����@�"��f6���+N&&m���NSd=C-�ǸGIczT*��3�8��<\�:����p���'�U]3���&���zc�)x�x��nP��5n�=Z�N;--<�,w{���d�t�v]u�Enu���em�K�Q*�f�a5RJ�^L�p��xO�:�w�-����`���'l��;���I�=��E{�Fnwp�ݣ�p�g�.\f�����
<S���K$0�Gq�}�����m��6�]xޟZ�h8�-LV��[P�z2¼zt@}[��f��j!�j[4�!
*[ s7
���v:��.�*�Y��ҳf��}���(g��{�p�o�
���[�]�X,�ձ�b�G���*�'�k�U^�*P��4�0��N"�p��x:�s��xw�s�6�{��*T�G�<���vm���ÁQ9�8��6ԃi�3�鵛�bah$O�vq\��绶�'��A����&7��c�VD/9�DH���2���N��W�CS=l-ͬ�Y�ó�7/)Cy)"����]����|�q��^����h��	���/�rg��/��e�S�~5+�V�@V�P��֢ +�89M�Xk^#l���d�ee�˚�~��=h�u��5��Ua|< 1����U�O����lc� �~9��H�]�aU^bsƳɀ��ߟ-��c��Aܟ)�
O2Q��謙&�<����:S|o�g�#�x�����ϡo]LM?'Jʡ���x
p��U�=W�MaU�u3�ͤi��J�ظ���!7o8+^c�:�S��ܳ���g'˚���!���ٶu�=7��%�Y�I�*�E�yp�v�w�Yˮ���]�7�48F{��g�/�0T�+F��y��z���a��J����'�lA�ާ/�i���.�,���p:K���u��Z��T�h�n���%2�Ϋ~ݤ�V�{�˷ٞ��-���p�U렏n��6�?
����yxRZ�;�����5l�7iZ4����voa��c%UY���02�����&�Cg(7�_�Y��]v}�;�.�b�w3ݠ@�Wr��p��E�'�^
Cx�a
&�.��K5��d\z0\(�fѾڳ��J��f5�,�[�]C�;���^�^�)�_�<���d�XiI����t�����1yu_  �����P�B/�ø���ysR�ZF̱#��z`��,�!{[W�u1�*�(�$� �a��1��A5�"Vg��VO�.�9e��E��{O.���M6�!j�QA����Lv�Cr;#��4�k�$����o��p;�Uɍ����`9�1�H�|��F���9�D��i�Gn09��i��x�J.K��ˡ�Y�����ڃ�����|(�\B���9���ق��J�sU\q�r�]t_}}r<�~5)���v���"� 	�w,ԧf܁��,cl���wY�P��
�T�97�M]pR5Җsg*:���2�v���Ɖ�q�A��Ի�0x�:d��\5����i!����^������ؖ�9팿.�T�}�ތ��
++�)���Z����������c�( F�ոqm���P(����^C:l̠�n�wP�>y�
�PA�;mp����C(���[5i�RX�D��8����5?��T7無N��}�[�>V��g����&y�oVnv,� :�C)�؈�qL�ixV�y���K5�3�2����V"t�ҹ��ް���wܰp��/�ӜD��YP���uq�^�9��t\&�yC�Mܴ�^���{�i'���ħ��k�㲾�^ם(Zs��KWo+\��{)AS��5��^�V�)k���:�H���K�iTg����\�8�r2���wo�y	OM;��췥z����`M�qL�[<I��^�U�f���ph�R�m�3dKo<����˧u��4FC������}�1Z<8P�[�!{�yz.:���"ĵ(v=�:F3c,�tz�`��|:�>WJ�8�܀���#�p�8�����;<x3k�[w�;݋��ظ�B��̬R�:��:���BNd�T���8�(��<��u`�z�+G�����`��&�mIYл�lF{�q���. F]��9��Yɛ}¥�=�t�u��dG^�zǖ)��COB�j��A���>Ԟs�Mǻ������ja�`N,�(i��d�8�Q1zҞ49^���A���]C�zN�k�\B7��A�9@�ƚ����O���d�u��\z���'J��TN�:�l������"���\<�#�п��0:W�Ou��$�]�Fd���6��G���=d�D�ϼ��kA��W���:��{r��l͝���W؃ �f�V��&~{;�ߙ��(��hy�|=���X�ve3�>fa����}�'��ُ��F�O٩B��#�׸���J.��¡���K;���{d�k�s���W�<�q�zG�Ì�����:Ȭbz7��8����.h\TW��2\z#`b�(��B{u��HOoN�Y��}�Ɉ~Y]���_Q��c7�S=�Td8TTwm�dJ}��^T}y{�,�!{������B�ӆ7.+;"����<��MϞl�tT� �J!��6�*P�ɽ�a�yC]�9ͻ�;53��p'^̮zfN.4��Fvc�����]�� 7=q{=�#�L��	r��R׷��
}��[�1�js��r�ZX�����Q���\3*f����G�6M�x�Wh�+mq��_m�l��&Y�y��<*מO�７
L�@�� +*��c�e"�я���]��{%�����&7{��퍋؀�>���ϟO�����۪S�*���61Z��+t�NL�NFAC���K!�h��Ƞ9��E:��OJ��Q9ʮ}M!����n{��^���U�VFY�iu��V���qz�Pp<`�V�^�d�� x�yk��֮�i�=p����Gq�#����
$z��vK./O� mЌ�<o��W����2�2wJ�/S͗ut��}�xʦ���,{����;���F϶;�`�߽Y����z�k\����\�(oJ6������k��:;-1\Vy�;'���&0�P�^~��]�׉�WI�LG�r�=�ZCK=�g����k���+z=�j�&nvC�"��l��/�n�ȸ��:�
��?5Q+���_k��t��_j�t|3*_��
Ν��N�ט�cQb�'��A��d�'����5߃+"���'��CF�[>5>!���L��Y�+��z�L(_K�j+��`����Wt�ݧ����^�xss��E�+G�ڢn{;��;/�p��Jt8���܃Q�Z3$�6���gV�W<�v�u�u7L��G��e,�$}S����(e03��5vSGf{��gN�Ќ7���T:{
δl̐�����#��(���b�P1����{^�g]-��e@��#,�K6��a�-*���5�(֢!]!��n����f���Zs.c���N�n2�	�aB�vGE�����b�н���֣\��rDo�=�w1�Yp瘚�����&��]�Zfs,9@�Bd�5"�I�MБ�E<]+��]꒛������Gmڥw}n��۾��?a�~^E��7&��4���z���,4�N�&Ɠ���������b8���h�����3LV��W��q�m��B�,Gb��"�*���zO-�w���U<��5d�v�0�b6�66�D_���f[�x�R�f�њP�.�\��r��8$�:rn�����A�
�J<��V�ڿ0&���׺C�;`'�X����܇�J�������"B�w:It:WD-3�p[J�|7��Cx�4�§b>63���+s�Z�������4e��~�Ἔ���Σr{yL��)�nu����Y�[B�%}C�9vn�^�uw���cSY֡��\��rn��H;���D���
C�ب�lإ���oc�ؕ���㖪�H�eOaA���O��5N��mh����L=�@��Ք٬��@W%�k��c|��]�T�F�t��Z����ve8Fb�o^�5	oQ�f��-yʎ��sr�� �?hG����P��O������qoev�����2�0�z��א���Ͻ��l�pR|��׺��)V����=�X���XO���y���R%��s^��kt�L���C�m��X���c�*BƢGi�_]n��S�齰�Tw����/�Ba�H{�ԴG>��;��fÙqB�歓��h�W���,'��Oz�H����bc!�Lp��>׺�JaFqfew/ <�wgM��.��q��k����v-]�\��&hʍ�@�ݙ���[�a��Y����k���&o.;��gz��؃r��T1�^X����}*ǻfHk�ؐˣtm���ht��Y�D�����m���Zfc���J���Nl'���Y�*a���C�J�8��NU�'���#�]�=P���5s(iq�ױ��m���.*�E� ���i���nuV����鵾��G��̂c��!_Ο���xJ�7�qOr߂���474!���K��km�D/q�KT�n�����u���(
.�LI���a�<{O�U��P��q��g��ő���m=�������P�+�읱ѹ#
���w�[�JC���@��uҹn��ar�껩Q�A�=9���K�I��3���sV鸏_gf� �gz�;>�OK�b��<vU����@/���Oo-��f��`p�b4Ϭ��3X��A":����\�ι}8����%�ϟ +���|�U}���:����F�O�o��w���Oq�'W����YfY�sĞ�>�8��Tґ��;�K�f��I��'w~�,A�a��3� ó��q�%�y��h��<4��y��\*�t5��k;F���x�K;��[�i�}R.���r:7�vɀ�w�1m�e�l�Lp���C@�p�oρ�h��gn�1{A���@ǒ��Q�Amn�G��6܌����gĞ}����	��f��)�э�$T@�b5A�1���@A|r����.0���e��t=��֖�T����e�aR����8hoR0��Q��J.§�p����������xnffzRU"$�7/�G�{1v[�.�
���r���Z�=����=������W]/��:����V���|�ȣΫ�%�M�����q]�3��DD�h9'O�ڲ�Lev+��x�&{e�{���tqQں4��{33\���x���H��]x��pcb�
��'2Չ��#j����;/I���]��G�h���MZOo��ޠby��cn�lx�L��q8$�F@��2m�<�/�V�p��N�c�7M�9����^Ӡ���o.e��e1�X�����g��C����kJ/Ř��=RY����a�{i{��l��9�ȩgb1�9�����,V0�M��A��h\TV7���~A�\���䳮��}���n<>Bzl�����m�3q��6Όr��T�U����O}�Lof��Z�g��#��W�!�|�\7
�ُ��8�x<&��B.u~6=�h��d8�SK�hi��YR�ٸ��u�7�a9��\&�
B��������
W�qz�je�Bt�#q���{�� ݘa��E*�צ�](�k	�A��~-ux��>����,��9�X���^��R�ޘ�/�t��㙹t���OelW6��� t��U�;)i�^��r9�H��ױ���l��U�W��f(E�e�����w�9ƛh��sj�b}%ak�&�_���m;��_D��cR7�}��`(�}պpwIgb�����p�z�0�{b���n�+��!fEL�T��k 
�]�4�� ���=_!�6%n����y�r�� �'X�1�#�FwcR�<o�-X��]I�jʛ��(���m�2U���V��U��.�Q#ӝn�F����IU-������w�;�F��7���t{�/���*k�gإ��[
��2k<�}BWP��r=�:���fXW�/v��.ĩ,����V�_��е&D6l����Ӧ/o��ԕ($4���ϕӡ�x�E~��q*��x�e�,�Π#��:;����ұ�z����7f;��)�&��+��Ch&~� ��J�Qp��{X#�i�F-�Ӧ�f�@�e�;WF�4�ޅ�4Jr�VR]� �n�m�;;:��a��Bu7l��3���Δ�	k]�Ef�<+\|s����*X���a΁��-Y�ۤ)d�Û�p� �ec�$�����v5r[u���OU	u:�.��s��k
5�JiP�GowO
�rb�+i�$��yV���g����*��|,5�N���Q΋q�\u���/>�E�,���n�j,�%�i2�EQC$d�kmn:0ҙ��قcަ�Sx���c��w���CY��QV���:��k4+j�g9�Y.>�7�.:�-�m%ْM�@�n��C��T���i�3�!|~1�tqp5�_�>�,�n�y}2�c 褴�8U幤�ۋ��&
�[Y�)D5���7�ފÙ5e���P�3��R�t,��}�^PR�\u8'Y��<Җ*]г������Z��2��+���Qx����^1�pͰ�QͥԌ�4�fg'�6u��ҬE���[5�<�	�^���v�!���3��l�IF��nI�A��Q\��K)Xu���u�B�r�n��{E�s.�V]��;�UB�=��']aU���Լ�pN��-p�=Fj�<���W�m�d��E.}�:�Kf�U�]nVv�rޔA�gW
��6tv5�7s�K�c�|f��^T�3��yJm���_]�vUӚ˝ͦe|��U��
a�S����u���8���������Wb�-U���}8�!]���M�tY���ǲ�1�9�����z�U���O��W5qr�xoP1s������S���o'G��,�X��C�So���w�N�F4Wm_$�.�����Wi�6f�{�i %�;�b��u�gt��v�8���D�G�F�A��Q}#����K��=�kV:�;S�++�1u�S2���;��X~W�W�o�����\����X��z�R�`᱙h@����׌��֍|�i�d3��^}u��t%��\��+�]�E�����jZ*ҥ0��N���ȇj|�n��+��f�Ifg<-�݋�T;t�������O�:�5΃�l���ܠI�.��ɹ����lI8�62��^�j�m2��tJ�}�92��[�K.��Bh�]؉![�v�ۺ2=I���Q�׽�rWc�[��K+S@��wK,D����'lwa�]'c޸4WƀD}@|(U��1�m�F,�y��;;��v�,Q�H�+�������[���5��]k����'v�m�.��خ;��v��y\Ѽrɵ���1gr[���\�+�B�sw].�p�7:s�B���u�e�WwQ����:�ˋ��Z��+r�
wj�niݮQ���;�Ƽm玹��x撼sxƹ9�N�r�v뻖��ʹDZ�r��w�QG�F��E��9r��\�1Ʌʌ��x�i.�ҳ�Q�t�%Ӽ��ˇvø���9�s�˞<S<�y牼]���1��5�8K����QˑQ깠O�P���#�*�$��R�y���%�=0Po�E|�����֌�L`�1(��kkb�Z�p�T���{���ϳ_�}�Tu�ks��=�7���ݭ��U�_P1�AK�}P}������?�פW��[�}y^��7+���[Ͽ/j�\����y���m�W.W/�x/��o>�ſU��~6����_Q�c�#��^_O��Q�x��������ƻ!Z͝폀�����d� o�s鷋ϗ�Ϟ�{k�]��羯o��h��瞼�z���W���^�\�t&/�O���I��@@0=H����G��E�0 ���t'~����(����za�`xB }�G�6 ��{�����ߍ����wzU���6�8�}2 �� �1���q�c [����o�oKO��y�6���^7�;o#��?@�� [C�����e�9�s~z�3k^�ì�(P�c���~��x����5���k��żWG���L�} L	�8�Ƨ��G���<���~.W7�����r�޿~y�����x	�k��������7,�>��scM��T������~وp�,Z��^yo��{[�]��o����}����-�_��zk�z^-�����b+��^7��m���ܯ������P{������L �/~@�h�B\������[_0��1��Y"�kx����_w�y�5�h߫�������m�����>�|^
���x��2=�D*#�ǃ�����6����w��"}� ��n@Q �N���o�K�>Vk�)�w[k��1P<#�����D��{U��_W��������^,����W���k�w�������^��J�k�����w����}����s|o��Q�"� `P�>��XG��
Z2֢��{:���G=�s��Ɂ1�O���|�����p��޼���z��j?��� d�=��
��0y@ n��W��x�����^��}޺�W����x���|W���W����tx������o��	�#�� b�|���������7+�n��^|��5�5������ʽ7�no���Ҭ#��G���!@�G�Ld p����Txx����|������h����_k�^��y�#&��������t�>�}dD{� ^��|ߝ�ϝ��^���ƼU��޷��=�z` b��5� 1>�x��"��������<��_msE�}���{_���o������U���m��|�^� ��{�ܲ��Nl�]����ݱ�����[�3@�&��w����@������Y�i�M3�ޭ]��E^ޗFe��)�j��:=99��}ڵ�.�E�)�������o�٫4��,ݬ����Fu>��ɾ��2��hӜGB���ǂlN�YS�b��L���L��@P<".����>��\���m�W�-����W��v�����L ���(��q�0	�گ����w��n~5����|��ήY&b:~�����ovc�{ޗ��{a��?@�xǲ���ϔ �$L{���q�DltVǽ�>�����: �ǻ���à8���'#���:��>R�Y]rb���Z�M�|�=q�p&���~Wڼ[�^�ߞ[��[�x�o��T <(t�:{� �`eu�oO��k߮��J��~��ok�^5������֍�7���5���u�[���#��3e덕}���
��\L\�jDi<�1~N@���.�G�� �����鿗�}�QQ�����i����������ү+�y��7��m�o�}�z[�\�w���{W��U��_�<�c���3Qedl�~��U;���s_���r�m��������W����)�>�<L c }'�@,�#��m��zU����鹷wm���wמj5tIH�	���Ǉ||& 
-�ynhF�|�`�v�m*�� �(�#�@�0.�� L{�'��r��}�����|^��y����>6�T��@��υY�
d(
=�dx��yF�.[��龾�y����5�_���C�\�������3H��3<.@P<!'�O�ty@� 
�+���7��k�x���x��o�rr@d{�`Ly�> �c��h�@�q�L *��@TT(�<���/���tҟ�����?z`	�&� |6g£\�7ƽ�~�z���nz�^~u�c�Gޘq�`z�䀤� ����x�{���_�_Mx����z��@�`}�}P<#�:�����}_^nd�Y�8/��q�0 ��T�dz�ߞ�o�������⹿U�y盖��[�]�y�����^���z���\�6�x��4U������^��+����m�{Dx����~>��{~��b���釼��.>q_ ���'�1Q��*�G��1Mτa�xA s>Q����^�x��/ֿ��z�W�ʿW/�:�[��x�׾ן�\��^���^�#���z��ޘ�};�s�BY��6����(2\�t��t��[�����^���(<��f[���Q�Ƀ3Iu�����P��!!�%�Vl�2/L}~�q�]�fL��z��J�u].�I>�f�**wZw��޺�F�;`��<�l-�����$��r���qپ��B>٫x���`�.ylg�_�J�r�,bא�6fP}7����~����JժB��1�6yx��׫�n<�FYL��%�~|����\�J�p
�0����J��Dgt��[�����/��CV�`����3CN�ƪ6�qVj(79Ob1�E!Ý�/�~�]�"{�"b6-��V �`�}�YƄ[�<o���1��y+<��
2�Z��p6���,Wd�N���#��5�x��5�t�T��ɝ;}ε����A��������5��m�-6�DGq��~�����4� Wg�ZC�e_0'fz���sڱ�]"�o�K�&('����q�[Ax��q'�'�,9Ʈ|ʚe6�7�w�b�㗫�;��z�5�q��1�n�z��;0�כ��n^W�z2nOP=��<��뭳��
p�:�6^�n��Fl���o�*��r:7�ɀ׃����ڦ]��Ș��cO=�܃�t�o.;od�D0!b��>^�ݓP��-��+ǚ�6������:���'S>��/zIVq��P�tY�ZRJ�b��w0�
�sm@������bv�ŐkjC(�jV̚����'���w G�;H7�j�{.�ހ�K�[�`=c�Wn�ט�Q��L5�m�"���ų��[�`���v��׼mԾ2�t�k���'YwR������}�W]O;&.���1�OAzv^t[*�n�g{!�*g���Js�k�}���D�!(�
��urc�S>��Y��яc\���A�&�fr8����r��:i4hN�'�ߔ|!�4R�Z-ʎ�|�I_�z���罜���z�}��ç�Iޥ3�t���X�"@փ�����&c/�سf�#�j*����K����藀��7Do٩IU�D948���f*����ԋ:�<ϫ��訦�2����t�SS�^�����@tFV0�Mx_Rq;m	�Zи�����l]�v7��v�ڣFK��cS8�6NY�f��=�htW�f���u�f��f{th4����5݂��$�c��z�e�'��t�gDg�(:q;+��pS��ս(6㔥#f�)<�T[yI���=��y,k�p�Oɭ�W
`7��쬁^!�oe�n. T
/u
@�pM�z��L��������"�J���u>�Q�:��6�/����H��p��)C]�T��Ɔ;�;j�X,��x����ײ���;^p\`c�Em�	)���v��z�[�G	8T���R�uσ]��y��ëofϟA�ś8��uD�:����'&Z��3���%���R�XϦ�D��ah[3l2�3�T�S�Qhgkps���
�O@?�EK���3�b1K����$�
��3b] �n{+b�6�^��$�J�Y�z�r���C6�=��ڬ��!���2�:�mT!}=�b��2�}A�x��.�ed�^�ؿ_���8�����#lH�V����4�F�o�g��KE0��w���˲�m���w*��+g�X�P9�ږh[���8� �����2N���Ɩϧ�9��Uc!�,[u&�7w��ma·5	�&z|��,����Tm���� �^�Ge�+�ޙ���=��[��[��^���G�G�ɲSmLcI�Y�11Ѓ��x\�i���U�:T���S]s�'	���Os\��=�ۉ�F�Ce����d81L��擅|�jEI���s>؎o1�NU�NlIz�_Y�OVM�vy��>��&32x��j#]��!�(���P�3�$֮{��W����0��^��B�,3ܪ�;A���+g̞��[�qJ2�݆� �V�B�4�3�E(��4(���Jb�U�6�&�pu�b�)��v���i�ZM/@`���qҕ��qϖs�բ��<�p�;�s�uWF^��~8�ra��;����m\�3�V��s6�2+�WP)7��7���_+��Nu	�	MRٯ�� �\Em�f�uok� }\���m=%���]�7t�����jbP�`�6��y�����FJ�Lpsy���`۷���U�L�k�osq��t��YPƾQ�7�T��ϳ��z֙��d: �O����M0;tX#�ioqc����Y� ����J�U�:;-����5B��@�s��qv�6ʷ�J�]ӲQ�	T�v�j���
���ŝ";	�g8�K�8��\f[up�X�Ŏ�G�]O"r��H���M�f��I�︷��V�T|����xk�t�B�{�x�k³O�3�W՗�,�n%YX�מ�����9�}���LU�IG�U>CyL(V��:�;�R����|��������d��>뜯[�|���2χ�x��V��V��m*��^��hoXi������5��m9G��I�}�����x�##�О�A���;�>����:ŝ�qvO
���AT��hWcq�7zn�)�-U2����3�W�Q�Ɏ��)|��h�<��^�SRޥ,y�k�=�~��Xʵ}ŋ��N�a�z�]�d�Lf�UP�OB���]��Ttu@�Q�n�.��v{���ר���[�[Nә�T(��D�#���<���yb,tc���&��+��ŭ̧@������c�2՞�K���2�h�����M���;���\J�$(�/&� ̄ݗ�lvj��92vWbM�H��������+"+�`}��������|�@{�K���g�霕`�>���{�@�n�XH���۷���ސ�H{�"�x��P��$�9x#̠*��!؜���x9�1Ά�S�3-��șץ�^үUz��#�.d�DVm���4#��\�\-_���ha��ʚzo;dCj���w݄�3-��D:�3녌Z���1td{�(h���1������{G��`%t=7���X��Ɋu=�8�t8�s�ʁ�T��3�>���lL�k�{[�����Z�.<�q�e+7�7���z #���`W	��~|���oS��2��ʂ�{Td��eMlSMg����E<C�L���3X�p6񪍯f�6Ò/!a�-<�2����l�$D����J3b|����
�t���Y���/~�/���B������h��Łx�+�y;*�S�ħ��k���>w��"'�q�k�;wI��C�n_nM�\�*6����!z��Zn�����q@��.�SL���դ<7�����y_1�QT�������� h��ˡD&H��6N=�|�\� ʆM8�a�`iX�V���|�׊t��A��燶6��4m"�;N3y���s�p٥���Vn\�p���q�$�#��[��#� ZZ���Q�㼁�́��e`G�1k�u�����{��/��.��������w���'��xHa�ta���VC�iV���x��z��;�E�)��&���_݆��\T�����A���G��y?5�u���~u���sW.��z���b�%�R�Q������L�T�cj�cM�������u/M���-\��&��=�C C�7���JjR��"�5�o���^vМ�3��UΡ۫���ݕ�[ZeU����� 	�����騨���l��o�H�4��6,��cvU��_�mx.��
�)SƼ����$N������R�.*�U~}�Or��5N���{����XU��;>�yxt�hקe�l4�*����*�lo� 6���?r:��k_v���b�ȹ_/Q�pt�w�L�]&�0(��h9'O���eF�!��ŧ�(���9�V���?S��5�)*��C�C�����b�cQ�!�'ՑE������|�;뵲x�L�Wj��/þ�����;"���:/���/me��M���9�^yy�W�̯XK8R%��LL��,��Vp�4kd�;u*�TC�g9�3P���8��{'	�ظaK -�.�`�E�Kg �>�[&�Ϟ��J�%��64�N�r�w_��aht�M���ci>�Rr�s#��\��2��*l��P���}�r�s\\���U+��`�U�����/)�><l������tg�f�ۮm��ry9�^[�UL��c��
�f�
璤.�·
�vc��C�<�y�8h:+��	V���n����Z�������\�m{�7�a9����j�{.������V_N����C˸_LCӚc=�>"�J��06�4��������,����Uj����}�%,D�k�}�c���v�-N��LFz�C�c���5
s~��پH�+��)��{=�Wtiu)�fCo�vR�-�	��F�#rc�]¦��B�K�)�A�&˿.��^^씜����o�%�<8�e���UU�2����R�Fk�.���u6(�p
lZ�|�7��?/}]ot����� 7��O�P� J1wM-�R�c�e=_h�%ܭ����Z�#1��l�_!6X�O���,�WH��(�#C���f�x��Au���hr����צ.����ֲ�'=�42W��ӔPC��*�e�4��и1z����^�¬A���]kJ��פ�4�Ue�Yg�.4[�ȐsV��]Y�=���0��)5��+��C��u�0`Vo��м.y�D�[Or:���z^l��]�m$��uC.�i�;�]�G���6v���qW0F]�3�ȟ>�x�Z�Asvc僳��)~�����w���J��"*G�q#���K����d81A�q�p��MH0`v���en{!�8�%q3�������k1N�E�l�؟Hۓ3'�<lt����Ȅ+���LK�$�u՝��w��w=2b�8�dT��r<�mT*��8�C�ڔ��[>d�"�d��c-Tn�Ŵʖ'��1��(����Ħ+²-��"��ZҨ�cYB��[��䘺m[�f��;��gf �쎃�΂�^�1TW��2P��`jfsw�"�GE��#ǥM�+&�{׫�s����dzVN+���5͌r�4-ϱ{�]���i�mW�hp�o>_a�s7xS��;�x�F7���+&܇�;6dtDl8�p�zE�sQ��\��7&��ɢ�[o�3fS��]�NV����|g��n�B�a!V9�0vz�ȸ���\o�#�uvshs�Z��x_��%:9�!���5oUO� 4?�׆��t���l�8ﮥ*�N���β��=��l��k�-3��̃ҹ;*�SbR�[�0ޠ-���<=$���u���:��F��.��Ρ�j�rn��Ts{�8F������'�Pc��K|�����y�]M���q�ܭ�q.Cؐ��gu��+�{�0�-!R��fE:/:��!�3-Nt��(�h��ɜ�Z� l�ls/���3���wF��pR�T|��1?��N�,tT�:�ûx_�B�N��f��+��[qCŝ�V��]�qH��u��R��I��X�JN�^+}���Ǹ����b]�&�.��?R!:�q�>}
��i���
Q,�Wr}����v�U��ay����f�R�����=��̮����tu��^���Xyou���ɣ��\VS�x����W[]I
9՚�_w\;�˩^T��,q.n���۔xn���Wr����0���E�jҠ�o�Z����`׀t���@�j&���)Ӹ�L1�HR�>��f��:�l���ei���G��6���l�C%�E�N�}�v���n�`���p� �1};;���X��]�Wr��R4�X����cE4]�uy�꧹��&�g_T_����eF&�h�YL+.v�ј�nQ�'���h�X\p�=iJm�Y��`�Z����C��0q������2�6ttlԝB�G���D:�o]�灓��wF&�V����l�78PL�E��FlA��e��=�9�$�D�u8�օ�����,��A!��렫Nq����u`V�0N�C}�:���=++Jo�L�3X��j��0пx�v��B��&pز<���Xu)����6��n<��<-�*#v/�wn�(3�6vf��cx��!D2�p�xĆg���ם�㇨N6���nJ=�U�WK��5�T*K������Gq&�ʆL��}�E�*���F��g.o���ơ��d>���`���ʂ�㡶7�Os~��巳U�pÜ-9���m���W$���ԤW�G�NQJ��v|�X�� ��ŗv�uY��T�Q���f��Rے��b��V����v&�� �M�jU���7��D�Q��3��\��C(V��8��$���Y\��u�㽃cq�ʘc��ȭ�h����y�W��켘$�۝WY#�zb]��ʖ�yQm��Ʈ v���X�H$�l�&�p z�����ı�)�`$V�x������EV*#����M̽����QQ�t�k�xGW)t����]H�ї�VKL銻���+&���wQeu�It���^����~��4��*nd�m>�0��A�:Jy�IιENf�r�s���+i��qB��N�e����ue��RWk��km�IO��7��'<�Oev������&̷��W��w�;�q���7g�t�� ��7��'th��y]�̤gxǘw�Q)Z	g\�M���e�nf��
H��رr2l�1:��1�wJ"�k=��f�vm�%���Q��[�<ׇ�J��]	��&�0<��A��f�=/���p��o����r��8�Qs��]�r�wnk�';\�$nWJ	wu.������v�r��"�e�\�)�s^9x�\ܮ� ;�ww9�Ќ�X$���O���$F7+�s��ǉ�\�h���������k������WI]ݣ��I��$h��E��gus��9;�N�'v2yמ] ]ם�P���W4Q9�4[����y�x]��t�����gw�t/Hɺ�I �ww(F�9�n\��*2\�!4dis��s��q�q���nv\�0e������W9���^:c��<��iK�.�nY+��v�\�"����v��"(�G*����K�w;��^+�E��X���'wWu;��"�s"Z�9���\��:�+���t��������;Ac;�;�f��wwwMsn�>�+��!z��K�/u�ji�9�Wݽ�v|bGZ;���nE�n�Tu��Q��S���u�:J)�g���O��s���G�G¹rS[��[�����ם�sÒ������w�(w�P[�N�Ή��D�ʧz�K�=}u��[�G/z��};éU0���#}:��V<��c=F̝월�z5�׼�3���+��Dj#�^�<�&������#`��N��X;�Bv�&��:�t+�Ug�.��*VJW�������ɧ��
�鷘�����y�ؕ{2'�zw7{]��o�Ƚ^K��o�m}+E�y_����Փ�}����ƪ�݆�m��rnĦ͎��}4� vcЁ�o������ǻ��4�n�DM�Vu�KE���
����f��,O�ӔyC�&q�˵=nzōo�\.��Y�yW��'R�<��a��E�xť���.�]`f$g+�/ve��6�Xږ������>c�h�S�K����c߽���ג.�e[��`:%*���3���7h�Z(�y[�\wU�֎�\��w�[���5�%N�.��R�̇+��	�:Bi����k���u�u4.����v2��z�����pT�ǲ.�P�=�8�e7W�fgZWO�R��T�ԼrK��d�Q���B-�,�]���U��}C��ϗ��,���P�LEe.�y���^�x�y��Z�苳�n-����L��y�a�]�r�I�Xqnw�W���ȟc��[=���s�[l橚�c�BU��kP�읠��e ��g�7:���-����1�帴�s3�ջ���.˗��N��o[w;/Ln��!�]IZ����&'v}�:Q��r��^����WW(�/{�����-[=y�vnS�:�@t�0�^�-�+�U��w�/u澛����|�}}�w�,��e�^�s�~�ٞ���8FZ<Y�ww�z��͍��~�va�`	o)�6�nv�>ޛn[���j�i�� �^PW��:�q��oQ�~��@��P��B�������]�&k'�lV�=~;H�G}Б�B�&�{zKU�|��#�LWa�4���(��9!N���կc)[g.��'4�t����U��L��*/�M�]~�h�K�p巁{oG!G��'D�����ƪjJ��MB,>��8.p��[r�º�t����L�	k������LK��Wl�G'w<J=w]����+��w�� ���BX�8ut9�"�p���$��p-�3�J�p�{�0���^2b3�zzx]����TAYg�}��6�oEr�<
�D���Z&��3��~�y���3��3�1e'~Ȱc}�(o1��ؑ�P�5Ӕ�zǈ�vIW�ғ���{�w)1���TV��ER�w�U��_
�&6����q�ݹ9�,z��M���^g��7���kՌq��l�|Vi���BoTR�jw��R��ݐ{��c�7x��-�!c�9Y�˛A��GT;mw������|w�@��_{N���U쳜#��-����vi�x��=�~�M�Ռ����>�A�y���n�s���9�pznnm�q0���ܛS�wɾ�_����Fv0��oP<�c|���W��N)D�ޞ�ygvz�h�ᑘ�Է������{�P�;�����=�j��>������6kP�.��kP�{��mO������k��>r�r/����V�6<��C�
-<��#�NU�X�����Ī�e9� �ͧ$��C�_)��Zg�vEZ��(4�YY$%����^���F��]�pJ}��Z�Ț5t��w.ww,}K���*�u�G4Wc�k6aZ� �Mr��Y��_}U��ys�[��P	��>�Z�eoWE}�;�;�(n���q{�9K;���*�WX��zbȩc��w&�2�/W{y�<"��w��}��І��ʵ3�v��r�b�Vl[C�l�.��KU��^5";��f��P]��xOj�y���2�i��Z{_�˄�8�I�2y�PFٯHG*Ow���#���ט'N��i��=^�x���uq�A�Μ��r�::smEoK9��^v[}�L.~� F�o��N����EVgxwU����U��#�͓�7�~}֩W-Y�.Ccy��nJ�����k�𞡛�(����)�}��x/z*�'�f��b}�Pg��C�&q׋Hr�S�7�<铽��.�_�S|��i�,cѥ\���k8���؛^��Ks��RA���*���.(�1�_N�1v��cr�׭�!ήO�����j㘔Ԟ�U�L�[��PX�2�|�[z,�]w��M���-|�	1Dsv����,�$6�/�t?q��-��ۏe)�꿕���m=��u�:Kc��R�X���H�����rIuv��맦��	�v�tD�q�<�qs�5�-������r\�^�����x�6�c�5����@^+��9�v����:�n�+�����w21�3ٙy�r�q�Sjxv�l�Yу{��+��dtV��n�n�.�9�ry�S��*�:��@��^��Դ��E� k{x�F��e$l�6�yzI��3䲵������K�B��tojmR��
�r���ϖ'HƼ��Z#�ݝ�-�y����1��_`����xG����9/1Êo#7-���L�"���{��u�e��іy
�o ��a΃�"�3T�t������K�o����Sy�s�)�6�]��^������z�̛ۯ�˷�1N	M��R�N�!n��Ƈl�i9��p	����S�P��Ȁ�������_���J�1����?hY=q��kuJ=Ը��7�g��Z*d75��ge vc���ه�A��^\�U�H�eΓg)�h@6֡�ڜl��}����ӥRK�����ע�#AWw"7�#�����������ozn��w)j��m�Z�=�4Goh}R^n|-��W��̈s�4q���\�n��	t���ȱT޼s'����@���S���?=�xx��Ϊ<���f�v=ߐ�W+S����jV�1��yn�'����=L�L��{z�.^t�O�s�w���t�� c��'Nv��{̣��#�s8���٦�0�W1٫Ŭu���"BNG*������g����*�h�\p/^(�o����y2�]����C��wî�{��6�3��_����Z��y�O+ߤ����tKw�j��h�Aۇ��ԃ��z�g���8nъ��s�=�(�~}G��1�[C��c��g{�κ~n�6�֫}���=��8=&�o���cd54dL��D�B]ok5p�yt\�ޱ�{=���K+l������t�^1���Q�G�j͑G	��L��;��l��c�r��'��������蠫W��p5���^}�T�`=���.s��Q}�;��.Y*�l�Vx��J�=#&��C��*=2�ձ%�]��@6%K�Li�L�իc�{�[x�[}�q�Ok�3���wίxֲ�o<*�]����y�8�,���ڼ�J�1t�L��S	���M"��6[]��3t6��rISp��H�c:��L�����xz�Q����;Tll_G�}h	;���;5�o�;b�zo����CɈ}�W�܎z�Oz��ӡ�YWβ��߯{.�gչ�'�{��f��Z�Tu/{�`�n�4���%�w�!Dh��½��k���c������y���=ꃤ��r� ���Ӕ:d��>��C�>'�w��X��K��k��|�~Ġ���q����_�i�i�����e���b�^b��q\��,�/�Q`�o�7��@q��!Z���&):S[�w�lv�g��U�-ܯ_\����82���f�B.!�8Όꐹ���o��!u��62�7!vԉnr�~-f��Z[q��Q����%�ww	�7�m�WU� �*��c�M� '�-|��;���7*;�`�Ŵ���tO��Ź���������xگe��n[Y޸k/cx�>7W}�j�T����һs�/e̚l��P�<%>�+j��0�\9��Eb����N������ԡ&�K��T@��=��{5.�dv�#�5�A�%tU���K�m���	�۳**d+����^�r�_WA�\F��|xPY$�g�����p�6�N1�]���h^:��n�n���M�v�n�fza�kcnOl�f۾ב]�p=W�d_x����O1��O�s�D�'���fLKV�{R�?+�^���p�Gi�->�_r�r��-��
�>��b�,M�ؼ�
�S�b�Mr�=u&�	��A��jk��l�."��;��|�^�R����f�nۡe��L�����7UV�V�SZ�d���s5qN��8E���v'zm�oc,���]+"����fH[u�o8
���!a����e�n�n���f�K�s��=��7U�������{ض.Od��F�M�J�و=��]Cl�i9=T8��+��$���5Wd�r�#\.3�W�G=Uq�o3K��m�S69�;+�.`��3�Ҿ��TL��/\d�1>��G����E��_��~C/����>gn�\��d�]q���^�Q��d|�!�R�T�˝aF����4ש�F�m^�����EFQ!��1��b�F�*��(��i��֝�����-����M��u)��&�R���C>r�z���������㖵X�1�	������=ʿ}�}�D|����s�D�?
;�f4����@�[�m5
�=o�g=�,��{�u���+y��1�5��C؃� 9v�����\DF�IČ�YBx��Tjb�n��;\��nqk��p_(:��蛻�aߞ�陌��}}X����|��z��cnY��X���� ��s�F����,p��d���(�yys[��_O9i��]��ͼu��^�ӈӊ�<}I��s�8s}Z�^9��(���M��;~}N����Oh���l��D�ɺۧе0��@:��9�A��6v���^�z�|+�������c�qp��:;���u�uo��1�em¾����2��z�p���2,`��c{/J9գ�|�.���r�W��sß��s�ԾÝdtD�SR�;�ߤ��g�˝�Ss��˝��O�����¾��N���V��e;�y����FUϝS��^��"Td˵�����iuՃh���vw�|�w�q�%�,�Z�M�6�lp��J���΄ 5횒���0e>���r���^�$z����_�gBF����.̍�te�r�;4���o�v�8��$�Z��W��G�_���ގڹk��}uw��hI���;5��{��ם�3�����C:�ܑgV/)�ݾ
�}|�,�s����5���n���!;g+�+i�EF�vMC�W;[�*SĚy�|���+�ߡ�ߊ����;�;7!�����%��+�ҡf�p=\��=��mD�/���B�9�ƛd����ۅ0h�w����q� s�����{r�v7��kw�g�ǩ ��U7�W��S�h<�+9��b��C��9��y��<��K�(?ZU�g�=��7��Qb���shVpe
�#��XŬu&�`�Ƽ=9���_K���Ȗ�+[K���{~��og_����zђ�D�~W8�ڑ�g�����=�G`�W;���[�+Z��>������]�O	���=2�"��X�^�3~^(�����Y��q�̾�;}[^O��X�&�_7�u)rt��H�c	tG>y��U�Y�Vj��K�WG��-Q0��,��w���I�n�'�ݎ�
d�+a��3���a5�\LL%�%�mf�"�������ȝdw}F�k/�����[�Z"��j<�u�k����V�(ILTF��Y����]�����'wM{��Wh6���趠5ܯ�&��Ye�I-�7��8L}]N�6�v�c��7x*�VY׭�n�e��$-�u�kDQeKGdWٖ�4��Q�㈳!������GN��V�dR#]�l����UꫩϪ+,+OB�X�����*�9F����f�wwS��ݭ޻OHa��٢
��d�����c;��_ed�jC+f��~�pp��P]R����#����>���.�G�'�I/`�K�n?���yNyk�A+�&Uա���|�p��:�4�v�m�w�
ޜ�c�.��ʅ�o�Ƴ^�k�T�u���}�yͨ�.�H
�֖�\��WR���Dqb�`b*ߞ_r�Ygu
�	W$�+�iN�kG�
�ѕu�9���v�jSp7���ע�V�ם�b|�+��Y;�75ʃ�%"n����{�ZVr�n>5Ռ"�����]q��>�+�ؑ�`�=z���nû���y�l�*s�KRǦ��3gC�}����g+�[���2�8�T̋��5�p���=���b�'��k�1�X�W:V��5SggeƦA���p��\���n�U�|Rj��x7�'QzX�����`b�c�><����*v����V�HmY�1�{�R�ve
�)�Q]䢺S���]@������ξ∕|���+[K�TA���e�_st(M����=�:v�Eq[���z8_!:�cK�ۣ��D��	t��]H� �{�-Y(i�J�^}����E���WH�ܮj\�u�}�_Zf����G����b���$Rs�*<�͛�g�P�Y��&}q|�[�e�F(<�a�.<�Y�;�ݣv��-���ڈ\�B؝���,����n*�H�FҘ�7��������٨-̮�lu�閑Cu1�wծH�q'}T��*vk��7��(�n
�R�����r��1�jP��<�:ِH���X�hR[�].Y��f� �n���@��d�:�C�mعѠ)�>B��k��W�Kv�4�fŤ��ty�5'7��p±V�@�^W���锻��9]�gH+k�-���������+��uٍ�NI�S�V�]ݗ�=!:��;vr�}��
�)�xO�e�M�F�<�X��e�n>���u�Y��@����S����Laدc��ō]N��������G��{6��-ٖ�E����-����#y>Z�����+�X��x9jc�y�J'��B[h�u��;�/~4��#X^���r�K��/G0��Y�ʉM����A�b6��]������v�%L������)��I|BA����/wh��
SR3��(�wy��n�"7��h�����M92���t��6#Ac�;�;\���r�M$Q���^	di�����yۧ������4i�]�y�!y�w]�$�]��2$�����1���7N�7��E�ǋyr�<�(iH����:H�o;�]�.�\;�	s\�M�����!H���2	��Dc��$���G�^X�$f�����n^<4ǝrb!�wv1!�r�	wtQ���I˙����Gwn�� b�v黷P^w�n��%�;�1d8F\���b]�ᨮ��nAt�o������9Aw:ђ��Ss����,n�������r��Aoy��I�nW1����O�(�+�H�vQ��m����%]�ꆆ�n�s7�.fX���A:�(��F.�n=x���ga$_���Gk�h��� ���Zy�s���]�����o�Ϣǐ���K�;bɿgW�Xi�j�Ȩ������z{�N�����,>�@[y;@'�;���TGP�',�׷�����j��~��+����xr{�<��Ǯ�/ى{6c�6��|�eסG�]�U��F��5���{��K�C�w����-�95��]mL�b�b9��F��~���%���[}�c�<�
�W��k����tr2pR�ۜ�F����:&;�k*7�I���f	u/#�_)ɨ�v���Z�)�θn��]+����>�b;��¡�`���VR/��v+2�����}��\/6�'4�GU]R�|#jV��Mnw��{�hT�.�^c��Q�ⱡWv��6���c�S���S�+�N��U
�ىD�(�fM�Z�S��t�ɟfs����:�bqѢ�d�� ���Y��0��o�G'A��ɑT��)=�yn.��]CKF\T��,�:��l�٧8 ���xz�#���k�>v��U嵸�v3H{qI/U�`�9N������4kم�dg�����!�rW.Z�����Vw(F�4��N��uhlOz�y�:��xy����m�:�3?jP&qywR���7+���Y����#"�l­�o�C�a��N�զ�X�Pq�CT��"[Y����ś�Lysv���_4����;�3��`�/w�Ʃ^<�!�A��t�����Ry#>g���x�u�լ��9p��:�,�x9��k̜�󘮍ɰ&��[�6�f�*Kz�f�kq�c
���8�;�����ֳE����Ù^sv��d:U�W�<��w�]6�X��S�u_��F<aTΜ~�m}�q�t���eW<�����o��w"�-�ݠ!��	+Oܹz�����!ܹt@G��-k'/�Q��i_UZ>�$���e+�}3�d����銥�~�&�����/ʉ�w]���r�Ktp�Kue��W9���z�*0gz�u��s;�s�0�͇Yw�+u�,F0�������M��t#,���NxO������S�Wf������No��>ݐ�X�|F���;��e,�eK�.�Aq��F@�	�M�,���I�Wv�a�؆ⷕE��)m�G�&��,�-\�*wP:w9�]�sm�6N�_iQ�Cgngt�J'R�_V�^vB�l-�{� �T�g=��+i|�v�:[�ض�ٴ���K�]���w�/wo��Vs�;��^����� )_)y�Oc��������=C��P�Wt����&��wXo�Q�/�o
�7�®:n�!��wE8�خDcp�Glgk�n�7�Ƚ^K���\^�zd}��W9��t�nL�3�u���O�����\�m���)�lH�'z���j��G�N�X�M\S��[�����E�z0�1o}�mc'�����1��[���l�Պs������ʾ�-:�I�ڬa��f��b��;�0��iC1U�{����	�v�q;j+2-y�s���@n����;^����<�%����2wx5�jc���ܖ]0ە�56�6-_)�-9��� ܼ�k�Q���v��]Z�}бk�w��Δ&���{|/���y��y����K���a4�B�Qm�d���}y�vb���_q4N;�m��Vz�{jA�����sT��[�X_1`<���B�5f�X�mK��,�l<)͓;S#�M���6�4�QD����qܖ�s�M��}��sz��#[�/+�����9u�ڮ��&UW��j]�!�*�b[^ٵ�&��]7型���}���̧���u��7<n����E-���rY[j�g���t/O�ѽu]������Ä67;;q垞|���[�%��޺�e�A���:xdgQ�٪;���E��?I&���hsiM����;9
�Ћ�پ����>�Vd�{s���l�c��ubKn�[�f��=��k���iwR4i���/D���+��`?%���_�eY�9���%|��\�s=����"/ܦ�O�I��p��B�2z�uPG�����=��������W����qw�P6/T�=���o���3�2����F��d��Z��T)MI�:��f�ۙ
�j��Q��b}Μ!�NP;0��3�;�78;\�`��Ow'���;�1bg�U����Q��^(��UN��F�m�݆7�ٺ-�"��
�R���[�[��e��v����W������Q�I�7�M���f.[�57la��l�8�q̈�ڌ���L�x��Ý�CJ'Vke���ζC;�@��nJ5a�& ����X�Ԛ�i�{O+���ꎨ���������su_vr�篮E��m
��\�bno�w;]�s��]9)�"Ǫ��]�&VyZ��E���.Ьc:���v��
�ϻ�l���{�=�_�d��;|�g�ߍbM	w��4����ƭ�o3SY���M��=I�=��f�uuA�Ùa�T���Emw�����c�{�ky�μ}�uc���P�/�9=�/s�kyf��o�ٸ�OW�������~�27ʟE��cz+�����@�w��y[y[K���;gؕ�\�r׳g������x-�G����\�-[c����]}����ls9s�~r/v�v�S%g����b/z��@[R+�����wyl�B��W8��NcbUs�]���CNxN��~���-�:����Z�mpB���wX�f�.X��k�7Q�Z���:'ò��o�����({V큝��F!}���V;0��{Īu[ڵa^쏹a޵��v�������ݻ����j��9Pf�]92h��i2�����
����*u�l4��`��z��ê2�t�Eb�91܋CUsw̱���[�5gkT(彶r��84/o��� 74�ݙ��Bg:;޷��L/!��yPF���Q>��>��55F�B�6m=�����41�Yw��ϙˆ݌sNP����,���K����+��m	=o_u͖z��"���]�;�#���u����8���Ү�3NGgu,�Z�.�$�^�� {j�uȷ�Mfs����C���cly0�s5B��Z�^�̼�6�4=�4�x�\��~����x� ���5�go��
�S��|,O�uA�>�{^&��U��yCȹ\�r����5�[i>�&�X�Yί�J��x'���g�$y^Tq��M�!=qu��i�TҺr�;�ԇ���W�y��g�+��x�jy�mW��W�K�K gX~�"���Ѫ�]�9��n����f۫��݇2A�+X�e�mc׹R��*nmO�lm�x�����wx�6�h����X���rL�j���e�Ug���x�tt.RaL\#S���<jF���C O](�ޕ��]��g����s��g�sDyw\�6�e���5��91a$��n�Vp�}R�h��K8�+o�P�5�K�Re�=9�g94���}5�<N*��������M\�Й����ʾ��%^E�\�g��_E� {�-��C�y�o�S��J^�om�c���W�<c����н1T��wr<�=��`*n�_Y��w�h�X_w`������]z2�7�zxN�=f7X�6˸��ݴ�M�jt�f�&�wE+���@]Si�������=�#��q�З;��{��,1]�9�v�G;�݋k�l�it��KB���W
��:de[�ܚo`�	���#�3�>�K3g�wB�0�a���'�1��t�Gn���qݨͯY/�`<�߽4��K�j;���3�zd����A��3O��(��U��L�C�x�t=�U�>��W��m�ַJz�\DF�͌��S�%E0Όn(sn�r�;0��pvU�Χz�	]k����7������Γ '���cA�ōj�b8��/d
�bɝ�|��øM�Ҍ�]}�vw�����lr��S]J�.�V�ys�X�ө{<�s��/��ߦ�%�ISm��r��:�d.wZ]P=�'2Vv��B��6Nѝu�L��eNo/���T��a�G��j���zm�� J�*�������Kl��q������y�*��],���ic�3����|b��dNV�A	��������,�w��@��u�z-�;B�b�]Llv�3���Gg�>�"�~Y}���Ź�Z]J��^Ӝ:���͇�&�p�a.]��z+SwW�ݛ�s!��BjmO�ռ��>�w</1�aBZIJ����;�-m��U����U�my����Bnu	��e�]�OX�v���k5p���Y4�z�qK};4��em���zW�@��+l�>O?gy���g��?���)���w�-�Թu��W9����р�_�x���-P_V	�tNS�r5���>Pr���+���7v�����H�wa��8$q�
/�����S��ގض�Q���C<s��ڲ�U�.�/W{yQ��TV��{&ׄ�`�t�<���t�:�o�˭��{{&��a�9�*�+dr��[6��k�����=bZ���[�Mӽh,'�.��Wo�he�3��N1���9�a����ܽ��P�y����ũ�����d.=[��95�v�Tw[�c{h��K*;c+��xxx-�r��,��vh�����q]��b6�{�m_�m|�.��5o��o����M�:�p۱��e{�\Ƙ��FȿA�<8�X�r x�cQ��u�5�zgۯ#���lO�ӄ:i��ُl�Vx60]2������0��m�S�oi��&B�pW���C���1cZs�5�E"*}�̬�]��og�D]���x�Jܡ��=X�Ь���F/76n�����z3�E�w^��Fǫ����|~?dIO\Z�vg�����3��v�d)-姚/qr�'Ph/�v�O������o�{�V�u���}.JV�3�����m�����y��f��D׼�o���	gz�VOx^�8B+cq��]z�;�G+D��v�9<f���!�C��ؖ�ge2Ͳ6zc�]��E�?N�/FȾgc*+{z���.�?y,���O%-��Uf�h�(Y0E-�8�j��#'����+�ڱW�9=�w��e�sPrv;W0�N^wW��4���Um#���(,��d8�rtic~N�3�^�qݙ�6B�V�/\yF3Μ��'���1���I������P4q��.��#���NBY��2�ENe��}�U}�W���s��Q��tozV�/����]�==ÓԶ�n�h����_�Y����ܺ��s�#5������;�U;���\<��g�T�罀�ҥO+�7�'Ư,�s��Xs�����w}*��-a]�N(�yQ5��������"���=�h;�kͦ�2ˮ����vz���of3=1��΅L�a���^Wk�6i��je��y	�8���C������m��,6������v�o6XM�ӻX;�!����>Uj�U0���^��˩�g�4֩=�WS����kݥ_%�y^�nE���(�KD�����aj��%�3�������x����,3��
����V��i���ҷV�!��P�;ke��&q컡<�WԹb���0S�Ǽ�a��3�v�<�޷�tIo4Fs5`c1�/�<�m��v�����߀�\is�u�O��Q7�Ӗv��#]�i���5OX��2�	�`tM�2�o�F�F�,�A��`����:7�iSGgH���u�9�|i�!{�/p�p�E�t��.��!c0�	�ʔ�(مAj�X�����Mn쑥�5�+Z�3�h`�^�)Wb�w��:A�u��κ,R���tQ�ë{{� ���[��]�m��\j��i����V ��ԟ�Ӆ���Rr��h67�z�]���!3�Wu�|�˿7
�':��o5��/[#uE5��1tl2e�rN�)�"�-�6�˼�9#Co��m��޶�u�w<]Lӥ�s)���|�u黷�*�\�@��2QK��@��s ��ͧ֯Rf	�a�[�.�15����$ހ���h�,�g����֪��p9�T�z�����Q������#r���O^�a��׼87��ղ�=�S�f�`+y�j��K�vW��q����m+�&��� �s{o>]��MKn��W�cq�W�2jn�m�-Н��I�`R6�0��:��Gk���� �M]�u���Ģ�u�Jb� /�9Z�*�wOnS��'v�4�L��ʀ��a� ��3a�A��9�M7�e�� ��Z�;��� �K��1G9tn�Iՙ[��#1��4�lam
��\]�N�\ݗ��
	�q�Ә�b[���{.e����&��"���}�Ǔ��@�ޏ[��B��`�UE��pE�,`�{�nG��szA	y�K^�*V��/��ڝ���:� �q_�V�z���Gӫ+�k��r��&�N���^N��[:�V�	��Q(�VW�4����������Եo�Lۧ�pP'p��v֖hhè�K��B�vq$��Ű"�����J�
��wz/hwp�����!���Gqh���g!<Wq��xﳰ9�$E�W�*Oe�ȭҋ諂�՝Q�Pǻ��uŮ�T��R�u*���̒�=�
ПU��3:�p���kיW�(p!Pl
�޽G��5}/b�&JM�E�j0��#n�\*�ʭ�����2��o��ZG:�iu#�NVus��}���_A�4n�vD�8s�Xj�k-8�´�mΫ
!��u�'݃ہ84���z�K�TFn�S��������6D��(�ņ��Ř1�Ӻ��#h�wVngt��o���ܯv��aP�7�Lt�@��c�o-!@,�I��]��E���)�kw��o��N��%=��
Y[|��*ܙC{���(���^�ƶ�e��dgR��'�u�V��v��/��6�t�|�"�3\��ii�Ѷ��TNV9���1��2���y6���v�3kDUʷn�Oo�iJ����^a7bI3�)+f%��a��r�<��;tt�E]N�HN��/Yr�/Qg)[w���:8:�����V�����C��ne��5i޼�c1)�X��S*k�����:��D��!����&r��r�Z��j����Jt�֫�~㗤D�y셇����&�wu_�e�J�K�	ܻ�X��r�˻�ID��,Xn��iRD��)��$��li(H��#$#��Il��2��M��+���b�����ew\�5�fGwwmt��r�2H� �wutۺ�:�Ԑ��.E1ݺ��eݺ���78&1�C%��b���9M
(Ti-&nvwu���\$�A��+!���INu��3&�Q�����9S2����Q�	D���h�3N� ��dw\�2���%͎p	4	�Ir�˦G8D`FI!�.�\��2Uˑ�a�
�Ɗ.�$Ѯ���I�  �҉��\�LQ�
�}���Ʃ�{L��ό�6Ekl2�鈚}�
���(Iܫ;u)�ڶ��ݬ|��M��d^ٓjӛ׵��b����}D}�؜9ܻ��w��=���|��nsZ�cA��P�:���gP��>���(�c�#�b��k�8��{Ry�e����:���2s,1KLQ%%4p-���sKe˞S�����ަ�w�k���r�J58�o)S������w9Մ9�mxd��UY�躣]B�b���oOR���������r,��E�>�{ӭt�czr�t<��/].��k����{�3��f#j=��J��2tc��M���y,��W�<z��т��/O�Kz�'v�(�� mlv夝`��������yA�y^.�ף,�o�0�]I�������bq%/3u>�7"[�Z���ۗ��6ܷ��yW{y9�Lmd�9�#�u鬮]�����8� ���o�"yz�b����@4�y��l\u�!ƾp��;��|O�0n4v
M����)_)y�i�}a��M��p��\̌ؤ���8QҊP���M��ض�@DeI����n����%颽�@���*��X��^��Qo7bw
V�ˑ�b}����{֭$���b���#�AW]�_R�3�su����K>0��N�7��H֍�s%9P�9������3�y
<�XT��9�hg(}@Y1�d�aPޡW}�y�w��{��,ᘍ��{�bOx�.����y::�o��ҍ�ۓ�y}ϼ�����[ӹ��}^�G���<�C���1CZs`���g����I����a��ު��������o������u�mb��]A|��8�0�U���R��w�.���Q]�����~�7X�ɜ���S~�pXF�k��7���{ܖu��|~Ė�+[�� �}���~4���,�]]*[���<'��{����v=�3�y���z֮����U�i����=يF���*gudQ{��3ix�k��F��s����o��d;]lW	o����n5>���]�^n�i�6�m�N���9�L�I�ut�,���گ+&>��ggz��E�h���óy/V꾙�W��T���k�9�3P�m��e[z��,�v��Jח�h,p���
&G&� ܾ���3v��WD��\޴^��Ϗ��h�p�ISos�<�����p�b�E]�E����.Μ9��P��jkB|<Kkz�]ge�j)�9��;`��ıv�Ov��AA�� �����{��+�\w8��u{���{˖��\��/j��^o�:x5���n�Ӊ��;�z����9[�N?h��*���~�~[�'�������U��ͱ�՝�]�S�߷��v��Z�.w�n�ܚ�z)]-z�ٍ����|�^�j�a�yQ�Z��F�dG?��Us���{k����^,k�Vl��z�v�9�6L�A��!DTʾc>���A�۲�B���������]�wGdv�6� ]2�e� mOm��+@XFd-�,^��ǖ{1_wnXX�U�Hl�b��>�NI�\�N�����;��5�z.��p�7�j�܋u�rL���;���j���M�ƚ�n�9]8��fx-�q �ͣ�jzܠ/���sk՜U�Fi��d#��u����[�����-�6;��8�~Ȗ�+Z�����<���F��Ҟ�ǜN��Tms7*���o��o�Q빴����A	��;����읖)�~�����mfP5��{:��3v6�f���;/�|���}�؇�glK(�N��۽2��;�n�����+�gt7R���2i�������R9iV{W���]\6����ڻ�A�>����M�)w��|i7'j_��1˽6z�^a����UO����u}�6^�9�L�8�ۓ=B6c|�&�_�0EfFn1�z�>��c]j���{'����^M
]�?l���k���'����/��ʝ�����ӵ{� 3z_,=s]�s���`��m�ۯIZ���B���`Wws�^/^��>��I�4�ڣ�{��鶻�8u\��gKFk�K���w����w"kJ4�<3���3�>��dyw�����0�B}hI�s;�h�^��:�;���y/c�[�v�lS��M��le���9>�������%���HI�K!��<���ӫ�aD��A�\���ҹ��d˹��F�G�������];����g.o)���OW��s�ɔ!c�F�˵�fJ�w;��y;������ݬ���z��b�u�8i�]�]"�z��f�Ɵ��<�sҊ��Va��	���Ygb��f�v�LT0�wV��itG2��t;�(��ns�6� �N�oPٓ\l��+�_L���L��������o��������W��`<���o�_b^Ry���U�R+:KM!�E��sը�k%x���������W\�qӷ&~o�aN�y��j6l��{5��jJA�n6a�3�;*�yܫ�=�ӵ1[�ٺ��:{e����·��^����ϟT=���v���� �ݙ����"�;�3j/4�1|頋�k㒻�=sv�+���K���7X,����ݛ���Z��Y�zz�׏g6�g5I��K�4&���F���{�N^��������9��m��4k��=U�p�G�@UxB��q�{��l�+C�g�	����_��|1�g��e�c�XswSE��5�%WL=t��3�W��C���<;P�p����˕���u����|�;�#�}�OܖW_��g��W��r�Vg�I=fe0]\�:]W��_n1v�(W4 ���SG�o��.�w ܒC�Ol��dk�Ѭz�[��t��5j�u�SW+a���3��#��wl
����/z��rLb�@�%@�5��RX{(�>	s�qoV���\4��r�zh�K�I@�� �|/v=���jk_�]��q՜����eo�]��z�B����y�{����6���S�E�����;�i���=����;�x�=&q�����4���X$�Гݔ��q��b��fߛ�^{��e�*��1ҙ�y�_@NxU�y��!��Es*7���%�/=��!��$X���
�
��CFM
U[N:��鏻}dl��A�7��q�o6�&��Ryθ�����������Vs�(t˔vc�����zd�^�q�#d�m�
�㰽��n��/��+Wt�J�-�by����va�A�^�s'�ؐ��%ױ(Y�'5���s�Q�L�~��g��]�c�q��(^��/��οTD�S��o��.�N[�ι���1ͪ�8���Ss�k���K8M���+����B,a���X���+K��X�j-�=O������ﶇ[��i�����1��5�u����M9�2�(��Τ-N�=�]ɭ7{8�]W�g8S��ש�g�B�c��`{�ӻiNGo�ҳ���.��=gR+|8iB�g�R��|��K�#\pQf��(�Q��d�S��y`�y��!vgU�OTvm<��V�q�����#�C������Q?{���e�������]Gϔ� �z�5"�K~s�\������^)��'<���E�k�����玗��X�W��s��x�����}΁��,7Z��-�,v��u^+��kkW����h�̂̚��j�b�ג�^���ezw��qKg���Չ_L�ֽhj��ګ4��;yݗJ��J�'Gr�����Ww���|��]�a���3o{j���z��;���8���A���"�u���on12����J��z�O7Ο��<$a΄"�Г��w�N���=ˬ�y���B��iI�-g��{w�oȵ]���Q��W���ة6`5�9�>4�U��켼פ�s�.�����4���wˌX���'���H�{��Txw��.q%��\�(��w�g��yU���e�f;k���r�4H��'�����=��+)V{�����g�c��1�r���o��6~���������#CiC�p�:݇)m�Z망1���k+��Μ����Z�aL�=.[�i�SE�ΥO�Z�{��u����KLW��ӅKA�̝�qn�of�{_����N�o���j��߀����w^Gt1}�A�S������)S̼�}�d�tA�#0�7�j�u��	�����:��7��L8��]ۖ����l��nC������t�b��~�_S9�������ŝ�:����aP�n���ig\�Q9��nק�-�7+��{;���Y�~v�y��_e^z�x������3�v�;��~��Os��j=N������j��o�u��߼"�<��ٸ�ST�]���H�8�W^NJ�H{�~��fp�o�JP�����m	����rx��Y3����Ӷ�E������ɕO�e�������B����c(d���⟺s���-��4�>�Y��	��mN��a��C����O�e����{�$�P����>���MԣiN�I�O��<ܗ^u�ǅ�9�RkI{��w�t%ce\,��:��o��A^o7b�(��R(S���+c`̫c+s�&��I�,G\�r��+�\����R�1n}�:��Dh!ۄ3�5��ت�L����Ih�}���)f�����B�m�H���m�ɣ������ѹ�\�ǲ]�������>B������tψ}�7/�\��ܯ��7�3�u*a��U�B��6��[�^(۱xn�-���ۦ�1:�����iޛA��FY��w��-�;)�m$��w�w]������]�sX��G<��y	�8���\��~=�����>kzQ��΅��?^蘬�wb:����n�9p�x�r�¹���y��s\=<H�-�Ԯb
�"�૎��dב���>�c�����[K)e��2�z�&�\��u����~�ס��ׯ��zR�{J7�ę�f��O����E���NW��z ���_��z���Z���
����=���n503dςz8��#���X�u_T= /HO�W��\�==�Y^i�Tez5>+r]cUrg7�R�c�2�������g�.��u�:���ūo>�������<!^/k�QGy��8iS�R�=�m�M��oH��!~�e�2�"��@�G�	C�G�ػ���{:�Kz���w���P�9�d`�I��h�QE\�7�S�k�!��r���J�5�Y�V?�eД�ts�J�5��fe�&�Φ�}����Rv�Rt��2b���Bjl����OӜ޷M��*���u���J��b�����\V���P�̯7i��BnmO�_��@ǌs������k�s��q��/}�vUr�x��?v%����<;4\�bb/0>p����5�=�TL.]�c�r���-����eu��9�)�
�H���6���op5˯;n���<��1�7��#��ĹzUg1g�o����q���l��5{yϮ��K��;�@%��:��v���6�MЌ����:��]ݻ1�=|O���c�hQ}hI�ɗ�hs��b�hz�v�Ҝ@��*��V�^r�wN�e�ӥs/�eY���3����T���_x�`��YE�ģ�0�W�۽�U�'�L>�,���3�]�oP���r6^$q[����^��4Ms���t8ێ�3c�sĹ�1�����o�ԏ_]8k�y���NJ�^��նX;��b)�w�	]���0;��\�r6c��ŉ�2�z7y�Z���g4�Ɍ��f���$�ouf�ei�I[����SC�r�^�/�c\�vep�+����kl��i,
y�p\t�4�3��m��YwW���������t�_�Ri=�EӦ'n�nU��e��H��"VU�P8U�m/�>�`�;u�$����t���[��&6���
����h9:��y%�z�Z��E��Q����;j�f7�q���j�v1�j��ufI�Vb��Z�N7���!'Mj��L�o+�gW%d��v(s�*7�R���$le�%�6���]Z�J���67�O�`���kz���DZ�ر�X'aAZ�V�NS>�"�U�fA{��J�xm�+SĴV�jD�˺�(m=O3Aޒ�N�R���OUK,<�k(�jeȞɸ���c+��mL9R�U��2�4�B*+�h�%gc<�7qT��hp�y輫�wW3^��p>'e,-;�e��Z�G��*���]+��֔M7�f-���h���깠S)�'�'��{#�ܶ�����(�Oj��s_,��W��mdO��(��v��h{���o,'�B�2�QV#}/���5�k�ZF�j������a�}ݾ+5�4k8���/'*�����Ԝx��~�׼�Ǩ��Z�s�T7�<v�2k�C��,��ݣ��̧�v�#�Dl�}Rv���������@��<P�̃�F��7Bn�*���ge�Y�4�EctX�0��(p����[�p�]��[*�d��]�OB� �}���x�Ҁ�|�T�i6v�R�^b�HU�\H�]M��8lQU!�6��s�~�+t�rT̳%�;�Jx�ě�r}���T�ڍ�Y�c�<�YV�Nf�WP�puqΐ���֪F]-��M�K�w0�Yt|���k�y����ح0T�ٷ{����PM콙yi�T��2���Õ6�2ob��˸pg���7V����Tb|l���km�b�q��KWZ'�p�����}��IyNH��]_m�1���L��,�X�Kݶ�6]n�\�¬G��*}��Y�)W\��J��"ҁ-�.Y��_r}���<�"C^Tx��Ύ�D�=�*G�j_]�oj�Tt!�����EZ�v>tp�ÅmN4��J�$�R�سj=�7;J��i/ �QoXѽ���G��d`V�Ut�9o@�v�|�jN�`��J�\���%�ZV�W���b��}-D�P�[���"+�37|���=���k=ۣPsU��x;��C�n����G)�{j������w���[($m�-.VV��5�:�u��Fp���K�Dol{�r�� �W�Sq=�D=Ph3�W�|�䜹+���}�f,�/5
��@E޺�x��].5�u��_pbf�u{�4��@�K��4� �.pH� 67:I�,J)A�M)��KH(L�v�9�6h�4a`A6;��22���T �F%Q�3a����3(�@,����RGwD��(DIH�1�a"�1�.u�h�.d&��"Qbb�Ӻ�č()��0&�M	�02Ie!�"H� �&$l;��Y��1D�wp&D�%�	��wpD�$�2���#��H2"�� P#���+�b1r�)���2@�(����n�"&
1fd�h�16�I
hّZMs���1.q��BM22X��4��RHQ&���4�&�O�������,	�&ίbs!�a��2[�a'�,m��v%l��,m��"�%B����]y��(@z�f.J<�@���h����y���t\��L�3�wC����(H�NQه�s����ܝ3��w9��4�ܩC����׷$���w1���6�1b}��²�P��Mg9�}ݼɗ��w-��/3O�����p����.��,軲�^�w�L_w�Fj��q�u7v��-�"�;a�8ۅ���S;�[,�����+��9��8�J��Byū�E<�32�죰�>��\q�nүP�Np�q�ͥ�����<5�=N|�iI�^#&ʩ}[��>���Zۋ+�(L�-���xD�Er�Ǣ��9�ߧ���X���G'-�(��c>�w���{���'�hq*P��3�x�&j<��U�x�U�Ur�`W�"�7�xz� ��<�)�Lؙ�������8�����S<�>�S�׌ܟ$T��h=P]�h��n=�.�E�����j��Xy���B�ȍ�WR�|j������Fm���-"^	�G7���ệ}�U�V�U)�9`l��n�k�-�c"o^F�m�{��6�~Q��b�3Q4����\�B]
�}{{Ou�C���Nٖ���_�����y�b�#6�j�R���tf���T��V{@��Ǒ\2��޳�{q�C�((����?����Z��]�z���^9=���+�33ʭ�S'���9K�\���77����W���W/���P�_�x'��4P[��ɦ/�(q�V��T=����(��������}�e��_o{Bɢ���p�Е=�x�+m��o�I�/梦Z�3�$-;Xld��O=���v�!d��G�w�%�ggf���Cʫ۸؛��qW�4Y\H��v2]�,Aw'sW �zgUT��oC���"T���ԟ�����q�2���6u�ݵ��y�G�D���L��@��axNO����������4�.E\%ngC��×�"r'�e���d��x��U�J�C鹙Q�X:����:�b�{~K�����Rjjo�ۛZyw���A��fF�j}�����p
��^!��i�u���|i`/a�v�L����sZ�:㞊���X��S����g_�.v;��C��H��;[/Mf�7qx���%;�����8�s>�1ӝK.�;�=����?}e�L�_~�6`����	ؠ.���j�(����⣉,�xN�R[��u����n�v��M�C;�`�Ymg3�~6�z^�=��Ύ:B�]Ҡ�N���g��9�>#�B�ޮ�ל��m�kb�ֈ��m�.(/���� r��w�VP�:�B��us�aي�gh�8�w�u�>����"]��_נ�!\?��ׅL�y�'�ת�GR󭆫��������/G��s���v��>���t7�T{�
���x_�T���0����֪�*��z)��n���� M�~�!1�ݬU���K�^�&uŤ�i��h�t2����,G3Y3�ub35�I
���x�z��}��t5+��is���^�ެ!���$J�?h�q����M�}�u
�����K�ܭ/�����+e��6*o���m\=�gvl�K5o����N!xi���y"�bO;ФUVߞ�k���qb�;=qrcW�2P���qX�,C��S�(��W�=3�?mI��mz��e�n�,xL�
�r5��U�B�iٰ���$^�o�h��ڸ7�ti�[��MV�"��o��,�O��fzHZfH�=r��L���Óq������/��ٝ���+�3�,K]m��ݪ��Me_ڪ�h{*����.��iP�e^^u��"��=�bMGL=���}.����}U�S�-��ɒ��HUV�FEq!u{�uW=q/�P��c��{>�p�-�N5&�G�"��^���!��X����0J�r�q�JTή�KOe!��1��`�pM�j���|L�v�=���͓6k�G߸��AnTK{�:)J�/����!s���AP�Y���czPW�5��5�v,�!�]�`p�3]��)vE��p��ȿ��""]~�佣ޡ�]gB�33����Sb}��Y�C令�ܪ��AL��J{�k²+cmk���l8�}UB2��t-*q#o��ˈ�gɍ~"���/�d�N�]Tvx{�=�������U�7�]8~�nT��ˋ�k2��ʭ��7pt_?e�}�vO������<cދ2^��W{��Mj����4_�VH�¥���7ԎH�#]u���^��d�ot-�&HC2��w��~��-ٝ����=� �,4����Nfk�K����&늜c��C;�9�V��܆z	~����{��	���d����a����#�cQ�c/U����\J���wC��e��eM������NN\K%NzU�E�R���k4�FC���-��RD.U{]¥��`3J^ʬГ����~DHV��U袆O���bk�3E���������&����*{�1\\��$�*�at�|ڸ{��p��5�@��ʹ�^[�����W^��L���f�࿠�9��7<������qqm�=5��w&S�$����Q�˛������a�������5��T�"�w1T��A�`L�"�W�$�L�d�Υ��\aU�N����:-�wN-��ve4�L{����F���ҚsvB��q���^�4V�P���+�d����B�{�R8c���'���i
��(���L|o?a3*by!P�s��3����Z6���������c�����^��%{c��N��ww�uUS�BfuR�P�+j'�O�1W:V��]d�u�8WK=��|��d�+kV����i�����f�7�$�SmYW�ʩ�����ڊ�o��U�ە��%����fk�	���:�ht*�`/0rd���o�Id_�ĉ]��\���W�0ݨ�=S�{o3ٝ{�$,�oլ���vBn�a����?&g�d�?E�q"_h��c��V{�eś{�镓�<��0u���g��㴚���2��J�οG�\����rEZ�Ja�e�o��-~���`>������!`{�*rr�)�*��{��/��SO����^��N�m����H�?%^�]W�ۇ�8s_�:c߃ɞ��f~c5�h�>�	Nʽ��k��3��T�z1ߧm?^O��6o}�G�ul*��E�N�"�='���W����Ew	���1�l�;ٮ�=���ga�ۭ�N|~c�IF������7��;9��;���S+g[�:� �/y;[`�4B��m�F���z| �(���t���:�v3u�1Ao]�<��4Bծ'�vlS�J��yo�\�nlq��8�k�f2^ق�����@���:>��\��}�C����i��v>����׹�~�)����׷n�:�H�S�Ǳ"�g��<=�����O����r�E:;��gm_�|���2ʢ��v��^Q�׊�f��]�WR�]����xE���<$d��"����{�Z ��ay>��_����'���f��"��SA��KB��U��٨][��#/6�k�zW)����H ��FI��WR�A�s�:V���I�q����٭�c�J������[����O��X�����AL��0:')`�wP�|�)|�τ������丗
!mw��'����r�Y�
nag��gG_�эB;P��7�9'5Tpɕ�g�f�Q��=����	�?3��wl��ij*e��<�{}���-~��zj��}����.��M\H�:��J8����!ʫ��O��,�heg`�~�����˻&��f\���jMz��F ��%OFc5=δ�S���B�&r�(�.Eu�-VY�y�7�p>�F���{�̤תa9/�~��~*o��z��K��i�{ޅ�g�P�\�ě��y~�Y�H$f���G
�
%�T�fRQ�5ʌl�.��0�����8�A�ׂ�����ե�y�`��dc}#/>0�˾<�M�?�=YFz�'+YFf���J�}YvT�;�z���eJ��o�^5��y{�Qc=�{��>�Ot���l_�(�ZQ�c��5t��>�UQ�~��0\�2.0,#�[���sV(p�T�>=|ttJ�_����dcf��#Y�z�Ra���2�gb��<�bo���_������]ql�\C�"�=���D�����go����O���C��L����N����lܓ�^<�<z���pR�.�e)��v�9�����c�3^��������Ҙ�G5"f|Ԡ�K=���8�<����8,�)x\�Dy�&5긑Լ�~j�/z��zyEO�˭�ތ�^�[�#Şz�rK��3 �:
��.4����'3=��}�X���\�_�(�&��|n��}���]ϰy��7���[*�F���4~N�XFk�X�f�g��Ƣ"�!]O3S��>Mfw`��)���Hz)�L,���M�GH^�� ��J�:5\g��{�*�rՋ�p��o��&/۝��#�9��HT���7�ڸ{�8��N�M!~\D�p詓4��g��ק��ik�vn��w{P�V%FL�0g�����07�b��ݱ7�LZ�3�f���`����ܪ����ŘY�g�I��@I�buaD�Zxm��B':���{K:k�}��w�3�����r��Nl���ü{)h�Yt��;�I�s}��ĀmC�m�Ħ=���H�]|��L� 1��ͩ��VNGg��Z�Nζ�ׇSܜ�{[O�)�N�'p�����?�E號�g�z�Z�[;;8�<�㸭�`�mm(��,�j��tǛ?@-?��B���,��zfO�ԴTK��38�ǧf���u���l� �k}�*�������Wi���z
��u�U���UO��H����/"C@f/�ތ���/鮫���VM�����G����R��L�e��D����$.�C����(}^��x,��AW���Q��gwv�ʃ��@P��g rg]M��s>�E�u��@;e�J*���3����_�w��~�?�:��6a_��Ѓ��p�8����^�8&O��E׈����4�w�;y3�;ڠ=���&�c�ϽTeJ����fUU��V�o��:9ߍ�W\Ȯ{��^k���D~5���
�\���ü*\�m)ΤrE�����[\�-TNv|�j�s׻�����o=��z;��qQ���i��|N��0����s��Z��t�:+��lޭ�=����Æ�V����W��Gl6�N���,�C�N���,(���(���o�3苒٬s����#l�"d��M�#=n|�3�VS�q˩ԗr>4�ފ �<���Թ��R��p뜭��e>����q���R��̈���0&�S������.�Wj�^N��J����H�O�l�t
���b��ι�������y���w��Jsv�cg��;�ide$�$��%�Y��56������w�<��=��Q9�S7�L�=Nʗ���t�=�����GҠ��<2�6�|�V�Z�gv�;��B륓\�z�Ou㸹1��\B��������u��'p��o"å��{��\C��Qٕ#X��X,�t����B�U�Ɗ��cm��
���
�����~�Y�(ۄ�0�u1<�Q&6�\��^��h��9W��:����������FW�z��v�~#�^�he���ɴɧW�S3ʮ�C����ǂb��+G��T����)ͻ~+/���? ����2!֜�m��ۇf�7�AM�H����1H�f�ȟ�Gk���C4��s�yCF��9�F3h�ꧠ!�V0���Bg��D�E�\H��`���wϑ�z|�P\���y5.���Dz��BY���wS����SQ�P��	��ő�4�)��o}��#���gv��Jc����y�����A�ev���)u[	S��8&:�(�$@�7�ܸ���v�{*}��Y���K����۔��J��F��������S0 D�.�%tu:Sbe���:��♼���O(�Us�ɴ�o+u��\/T��s��b���Lm�*q�읗�܆�wْ�>I�ٵ�so�(_�R2~����2�a؝9�����ҟNᲧX��R�Q�ê��R� �[�<����p���qw�
��zEu[�ۇ��pB�0\`L:T�f�{�^��v��֎��~!������2\�z1ߧo��y>�����=�ŝ���V��8KV��w}�f*�]��s����qV𙸮gn��n3s���7�u�r�όCzN��=��wQ8b��ۛޕ|��T���L��[pF��D�r�ǩYs��7~��ƶ�E����xb�؛�Ӗ�����N��"�2�9GE�U(u��e�⸙��b��j���Z���`��%ة�^�j�|��EYG��}H ب�02�&�<2 ���xjzz��1䊚������zOkK�;#����7�<�%���Y����0�.�Iu�(1l롖��4����L�:�W/ǯ�A�����w��WL�X����{�\ﾊyj_�V �<�����S'�:����g���_��%��/+5�*�pxܘj��P��#S��ٴ�]d��<�	�Zbr>� 4�j�Τ���]_gKs�赴sq	���]J� ����� /�q��^l4�Ϛ�QC����꾬zȋ0i��-���d��o�q�1S�d.�jG�K�������T�-�_]0W �;�]i@���VS��zMnö����{'�R+�QgS���9D堾u�:+�e�U����5ؿ���+tPF����O7��$�qR\��Dvs���]ޠ��S�0�\ܫiী��e���XV�8�k�`C;&ƙ���GgV�ٶ(N֨�ƥÙ�R�[p6�a�ů�i[c�+���x�|�n����F��;��nao-\��R���w����t���������LՇ�������gG��Sϋ�z�p������B4��mX-^���
� �HL�T���˱��%x]��0N��Tq��j��G��5Y��-7b�}�>lh�K%�Ȇ�X�y �k�]�Aմv���2�������ë�wOcα����4�9�ӕ��3r��ir����KC����l+��$l\�,����Y�{:>-�	}�h]�S'Ys >�A�Ф"�ް���q���i��|eݍumfNJ�&�lp>�zm(E�2]3/� �����P���彨O(��{�^Sf�@�8F�s7N��q3��f�*Ss77�լ�����Y|h�wA�Ԭ�b.�(m��ggaT+e�2�}33�+�t�僦U���������j"��]j��"�`��J�5��.����u�gX*���t����]��Ά���Q<ם+|h�9�OUY������\��A�,]�Xe7�ֹ�,H���0ƛ�3�5�D}J�f�,Eʇyn�]��� �q���[���γ-���s�{͆��V��2�3��:�[Gh�����F�b�y����+i���j�
��>n��"���zWZ�(8�<C�P��ޡ��Ó���m�唸�i���Ź}�I��� }�e��r�=y��3��J�3Fr��÷�u��fn2Y��� �#�C�6���]2y�Ź�p�����ك�8.�5���Y���X۳��<���Ƭ�ı��+J���o�8+Ne��C������=v4dK��0��C噧��mԘ���J�ډ�̒{n欲���97B
ΊeГ�<�C_K[���+����u|�ˇd��9�c��� ��5ggG�RL�k�8�2W}7�6O-���v�1�_��ދꝞ���XG;6~��u�a���n*�ڏ��E0����V��lV05��N	!\�n[�lm�SY|�p�	��>�G[�:o�r����%wi��A[��	�g�늰ŷa�ՃYMͲq�b+Ss��մভ�u.�,b(���)k��1�̫:�f�>�ڔ�V_�R[��#�j�=�XS�j�1R�۩�:� �������+��:�f�Ͼ��؅#f ����n](T�w(b
�0��e �b��I	IJ9�cIL�"�A�P�l�JHFlX� S��EE!Ww6� PFD�(�n�̒,4F��KL`�b�1	�&RCC)�%���M$YN�a&He۰Ɯ�ƓbX�Zd$`�	�˗JR�30F5 �#"�01��!GwL*P%�E$�Lɷu�wF�$L18Dn)"�[�FD��û��ۥ@F��1�]!�t��3AfT������j�:i�f.��sFf1�RD�,I˙6M1�La ����fR4�$#)��FYGv�Te�$�I��a�}y�{��z���W*f�Oh��B�û�R^Y��mr��S���+y�@f-�#�{t��W(� ���>N�.Y;w>�Ӟ8��·O뼨��1���.y���+)�lBT���fû��$�EL��^^j=���r����y�"�T��iSW!!���1����{aB����6$;f*߸'C��Z�Y�{5]����"s|���!q�1�Z	���%I��jO���	Hs8�ݷtJn(�Shw\T�~�x��D�~�)lC٘6_��h<&1�����408�s�=�}x(f�f`ү|� w"�C��ȩ�k���ul�@�{@
�j��pB���^�G�A+<o�%�v��s�/�U���̪���ۆ��k��:��T�^!�'ke�99�.ڤ,=���q�����N�3�Q�����.k�~58�U�s�������4~�1G\]������9�>�f�7�0)���n�^03�ޱ�S��M��?ɕc_�`�y�^���S�hhg=���=��xV.���¦k��:�\M���/6�z���ֲ�/�r�������m��=�(-b��R0z�ઙ}x\���fub��x�;�S�E���$ _lnT�t����}�M�n���mo
��T�����.�T� {Mj�Y��[T�7�k.L/2m�����w��>���k��|�%��ͼ�v��Ca��got
nRu���\�)�������]-����\�<�ܯ�~�F�nC}jo�ol�z-�@ �Z�e\g���(�C s�n{��*�-;�ۥĹ��=p�R��>)����E{�kQv֜]��Zu���U^ꊯ�8Fl�K:����^-��R�ϐHT�,F��|ڸ{.���v�i��$+tT�\�RW6rY��u��o$9���W%FL��=qrb1�}�!u~Δ�U~�'�_�n5��aՌL%4:R��	��s����C��<��&Gh�0=\�\H�6��rи=�f�&vs��<f+]5�Q�n{���߫moA�p[�5�Ź�:��:/TB7/L���Z��W��ٸ��u��-J��=x��������������|��&�\5VC�eT�?Ƥשh��)�d�W��\��dz|s�V�;'�C����@�Ёɔ��'��\Eq!uz!�\���b�VX��˴n|{�0�΅V/�G�<&���L
�&fu�92~�g�y��#>���MQ���樖��y{۫l?p������#�w��oTB�*q#n9ٜ����2~��(W�;�&��n���T�ۚ~����ϫ�1V�2�.����Yk,�/'^�N!rԈ��kϼ6l^���S3s�td��>�T��bA�j�_Z���8�o6��V5��1�lU��������S� *;	���s5��P��$_[�x!���FXs\�W�ۋ���v~�������2l��7Ѵ�a7*oi��ǵ�UW�V�o�����<�Q\��NW{0�����wM��K�i
�5���9���xT�?aҦ���rE�qz�Թ���U<��W�ս�r�N!�zv��z=�gt��|���*�n���!0;)L�y�s1�hz�hdNwn�ٸ���l��^/Gg3�����$v���!��-�W��8.Q/�c	u���_�\�Ξ�ň�1��p����S�C���;��7jU�7zGK�PC�W��%��#әyYн~��}��/�3�+�&�v�1>T��I�0��R�>����(y�!'�8�9�Ӊ��[�s�"�zY��&�*��*{��ϒF)z�:ĸ������ڮn��5��϶�D<���TT��Z�O��,j�y���!g���4Wϗƽ:_\�'ݲtݩ2��kP�ؔ~������,з0#�ã
$��뙸K�����wNU��q��s��U�N�g�@�v5�>"q�x�N2J���4��ʦg�\x����&*�GJ���S�uɯO�u����CK�t�Wb��˕�W�]�^�V��9t��S�=�CKĥx�s������w�bJ��>�~�A�Z���O_��Q��_-�4��4-@��FZ5 YR����{7\�;p�iMlë@��T:��(���_��{�<�K���,�p�*g$\6�Y���D�
n��eT�B�틧�ż�k=y�����wYQNG���욄s�uS����&S�`�"K"�+�����xzTx�M��gs�~�q*�Ԍ�^������a4 �aB�q:�� c!:�2+f1���{�~���z��$8�%�}"������Ec/�=Jp�3�sq�MI�F]U��9�{��o8����ޟW^�X.2Ç��$���x�}�(���V��pB���T��S��G[�<�8ꬱR_��vyw��"�ў���tgn#�e�޳����zEu[�ۇY^�^�Ҙ6��Y8���䄗�w#��4fu�}��5��~��Oד�u�W���8ZvM��8����������ބp48��ۦ:��Z���3�y�\�f��>E���{�Z7!�'�ʫqS�^"��U��wZ��\d)��=Ւ�ma��Ρu��s�l�쯣�<|���]�sO;�7������98�W8r���P댣/��ϼ��U��W�yA��jJOč��k_@^��
d���,�ʗ-�컶Cn��[�&(�D�ٽ��W�V12�whj�{r�LQ��E����\�� �1
{ٔ~�KY٬Y=�)�̖R��O�8��F�r�F�ӊ��D�WZ;��\kM��	�:�.�à��=Uz}�%]�^�'GX�8Tc�Xo��4��{k:g�����w�}H�G�w�Q���В�����t��F��t�
�Q'kU�{�)`�5NyE�t����h\
sޢ�糡D����hg�iT�=��}O-K���Ǒ��T�)�����,376.��V7۵��~��.�K�<nOћI�ы�`w��4P[�&��<}^"y�^��r�X�>�j�s[��ϜLOwTS�����;={�%e?J��p��V�;�`͢M!��9~�YG��}��9�'�EI�3�Q-؏a�3��}Ol!�U�m�lK��n�Dg_�{޼�ރeAl��.��/���N�Ƥשh7u�;�"T��1����	�J}�������[;�<�d�b�&R�p2��/�� > T�g��0�%�r��xW��N"��o6f/��bF���ܥ�C�dS�ngC�g/\eĘ�|�]*���UQ�s��
���:�v�����E�7k/�����Z�.��p_���B���mٜ�S�sY�*O�գ�f6v>���%N���^���5�66ⵧsW(�B-4����7q��8.�,=�i,����cĮ,7-��G��){�`i
 `�z�W��l���I��%e�n���Q��lMIPa=���Mq�X�A\�[L<�u_o6��yC����4kvn�;���s�{���m���0\`�0�E<q�pub%�w�~�;p�1���B��9�3&_�,=��)�q��|k0l��/)L��9Բ�\w;�=��ٮ�=9E��g��s3���?{�����.5i�;��i��TPW+'?A�����5긛���t#��=Ҫ	�N��7�K����>�O^%�<=�(-����W��ઙ}q����FgңWw�xz��m{.�N���̼�L��;�����u��ol�z�Tא�E\g���
��/Q��.ſxW�YD�F�rY��=\̮U2��RB�䋔Ǣ���{}4�֢�}i�%�i8�4롎s��q�T/����^�/٫����*����pw�ܘ�M�F��|ڸ{�� �;Y4�Ǘ!z_j���N�C��ܥ{�y2��_�1�E��ʽ.y\�����@�n!�\V[wlC�����(�T�3f}��z�:��b�y_��ɉDɁ��*���m��Z{N��;9��0��K���\6o���C�&�Q�w��Ub��bZ�Ёz�"��9�{s���9 YR��P�������FU.�g��#���R�)e=�Mk��Ѯo������=�7��]t��,�ٓa{*J܇L\^���w���X�<�tM
�tf�U�K�I勵c螄�1;�γ�����}����ދx����^��;�{g��1�[8����C>~�h�J���쪞��Ԛ�-r2S�bj�qC��K{Dˊ����;!z9.C� re;.F|��5�q!u0����[�ջ�e����c��kk�.w���C쪡�ݤ��|��֦�3��τ�g�ȿ��1Ϙ�Ԉ��b�	��.�y8�S����p/Q�[��b�AtFo;3����*�k�͓cu攏��`�Z���w9P���eV1��s�0��7�����̪��b�^D�5�)��6����q�<�_���'C�F'���G�,�A9�9X�}b��KY�*�����ን|�f�6�q{��O����K�7�1���tl�]���m�C�s�\ ��݋4��Gݳ�}[�uEc��ڮ�7ʜa���z9�Oc��7R;Cg]W�3�tU��������o�U���/���^D���1�fj5V�7J�C����Ȇ�Jn�ç���;Ȝ��(���>������-O85V�.T�VM1��MDy�JN�
)�R�;�ӧ��`bB=u�ߌ��5����d���{G.�6���]�����j�%Xvd���妮�vv�1�,'�,*��1,{�^�O��Ono=�Vq���6��n؃vh��p���-����o޻N�]Jޭb�;����W4�c|�3'Zs�nūHܝ��,�a�ۚ�:>�'�a�����(���5��pM>U�=��.O�WB��ֶ�<�a��S"�nf>Gz�k����Na�/��H Х3�h�C'Ʃ`�:y�Y��+��F4W�ܳn^]�2[�����|��c��-;5�ҷc�2�ۘ·҃���Q���S=+G�j=�5���9~�Ï%ĵ/����DN0�UO��ړi�N�ʦg�\Z��z� "��d����{t�1:��j�!�ӕg��`|=
���S�Ͱmh)h�j�쪙녜�b�7B�Ϸ����L��#�N�D���}T�<�����&S�`�"K ۈy6�W-�>��O����tԘ�G�_��&ٴ%�&�n�B�����܏o)L�x�Q+�*>=������p��HT'�`
3���1S�R�8ϥ��ݤԛ�e�_n��h����N�d�w�ۊ��.���Xk�1\����9/��9��X��*rr�)���3�*�/�|ttK�5�y�[M����qw��-W�WUíۇ�0`0&���j���-�jdO� �I�B�5�Z�aY�/�v:��9D�iP�#?�q���9�l�Ve���/��RY��ǆ��Q\x��Da:�p���V�_f��[	��=yC����|�,Y�ك5Mɡ �U��p����]�������GD�k��`��:|w����t?Xqt�۪�Φq��d���;���~��{��+{�H�~U�d�����\RӤS�����2���v�wµ	�μ���.w�MΟ"�l���n�j�<b�-��zowj�Y�=LM�8�6k�d���.f�Y�"n"�ZcԬ���n�=;Y�x��8���^Z�G�<�e��N_�����ʩC�(��W>Z�V+�R��}o��UzG��-#���Iw>�8z�\&��?R +Tc�Xe�O��_��g����Ǧ�j�l�	����GH����-y�wVp�zW �[)ƌ!n�_ʌ(�S'�<��0����^�~>G@څ��=�tr3o��>�Hg�ZU��S�T��}~�8K�mDG9����]q��� 3n�c�]%އ�X���W��rc6��!u�x��/�f�PǦ���W2*=r�G��������B}*%�#��U�Kj��n�����[�qZ�,��p�m�:�u��ްi�yH�e���PuJ��)��ǥ^3{>[�6�|L��,&���uE�?��ʅ�������d�۟��CV֠����զ3a��v4r�O:�|_7:�:J��Wo�҈T���7��xU�R��EIu�l��Ԕ�kp�[�>'U`ԎWp`p�����4���@n�R����]�*��g��NKg���4x��BWkg��Ƥx->���*Nc54_T����cƽW�/(���)3�I�L�O��YddEu}TNͅ��`_�'+�~M~٦o�3];K�4���m{m�@�m"�+s:�S��\eĞg��@�}[Tg_����{���b��f��w�q�Z,��x<6aoUxg���B��fdm�7fr�Y�z�Ra��6=����%K����qT�m�g',��0\`h�fƊx"�����K��}��fu��b�t��㪮��z���������a�yR��Ӳ�g���u�f3o)�ޱ�S���Fgo�����Ss�?g��>���hn�P/~�{�M������L��GdN�F'��	�v��!;�eb�+�)��6�ҷ���ވƷǇ�VP[�tc0\:*���x\S/�#��<�zߊ��J=����s;�<*�n�t�����Z�o	��U ��^B�q�"��l���l�S���c�އ�;�t��35�I
���Ǣ��O>GHN�Hr%L��Zfw�Y�=�^\zբB˰�	A�Z�u��/	H�4��a��A�Q.fYZz�\I�K9gp�V{:��+��P�"�	�\�費�r��otfY�u�:�4w��Zć$)o��+>3���٫�ה�t)��fL��>>�U�Co���j�f �u�9qǇ��4�.��-��]lF�PT@�d� �fq�x���A���t�r���I&���aYl�"� �&��:}wʷsl���u���G�*�K��ݺ���d�Ɋ���IR�v�u'�e�-uq/���m����(�ު/�;�	/��V���:P�X��%�U��66cj+/�w��v��43���`7\jv�5��K@,/����ɝ�%(<|��<>�0�@ۋx{����|��ήm�r�l�1��8�i����=������i�E�֛���H�ֆ���I�w<[0�.�P0v�C����CBM����8
�����a�j�u eq2�K����+q���(�R�z�>9�ƹ��>&/�݁yu+^v�R���KP�qU�8�Ϋ����+�i�U)�(_����ٵs$=�y�N�M�3e��Pݏ:�H3.o+����oM�K�n�^qT�	3D1�z�f���;2�vi��D�3wd����>'��($�֬�k���&�Q�]/�6Zm�\�liXX�[�̧˫��E.{�/�]�h��n8y��SVWgW[�ÑN&�f���_*��2��}Yn��ú7�t�i���t���啱-Ss�c�+�t1Q�.b��\�$��;�Bn��V�f�.[NG�s���n��-�,j��,�&�˧gw�ӟu�GNAN �3�i���7�R�0��Z���5{k+���w*�[���9����������Ȁc��gu���ը��խ���XF_Ύq�h���n���Z�)�]k��Zl��woNWj�u�\۱�%:����`��K��">*k���V���|K�]�w(�6Xү2�ηlg5{�CT������rʋ�,����^��k}�mC��ċ�pM-Ư:�dԊ�m�5(�s�2�xF��M�+�*�(�n�M�[;��OE�1u��N�� uI���#��V��f ��l,pI��Ü,=ó�}�8	Z��]�'C[XܺݕҬS�ɊGy8��������K\A�XO����}�QduiWWJYf�u�xFb�q�X����\�LmA��s���L�<%Κ�R�x������>[����8Ťj�4�쁡k0�Xb����:��3���9�Y��&���D�:8|���4v+�l��3vo�W� �QKge5�X�@4�_s� nMu�]���n����UZʏ;WN��b诫E��k��,�t�6����<28��Q7��Bv��L�e���R��X���Q�2m[m�RB��(��no5���a��;�ڻ��N�P�  �%2D���4� ߽�H`I�"2��2�"���2��l�)6,d2,H
��2TTB4IDfA1�D���L%%�) �#����i��%�0ő�JI3aD�$�
$�$$T�N���3s�,��Q"`�)
���4`��͒Ō�w]��0������8�M$��D
fPd4\�0�HHI"�H��A�%�Ԍ�P)b�"B�78%	�$�S���2(��@D���Ή ";�AD�9�k��"��%)����s�Ӝ��(�՜u�{f>��Q��1�G�IE�olm���8�ӹڳL����r���yr�O�w=��X�/=�ݧ�ߣ�*����خ
��I
�X�1�����@g~��ɤ'�2Guh��<3%z��P�$y��vd��ȸ��*(�[b畞��8ھы�`v�+"s��Toc�ۻ��׷�[�E;���f5�_�ޖ� ����ߊ�x���A��v����ʕs����<uGV���W���޸��`�'F���G���?�d�R�W���A<�;���n��=�������#����5�veջ����tCU`4=�UO��W��� �Os)�5'���j���w3����?B&J~�!U[5�q!u0���{�S��;Wx[�uIue�x,#:j��&��ݤ�����>@�ɍf|$�3�dz��~����<��]���9��Q�lzr �rNᑆ�+�Y4"�E:�8�����O�ط�+}��3�v���q������ˡA��"{����»M�X��6���nT��O./�̪��qR��*�\���º)�
�n�o�~�F�"���"k�;�e{F�U�2�rp�R	��D>n[K�{5M���Ӧ�����-���$��f,�U��:+s�sp^u�x�h�*�V^J����
����sy6����Wh���C|a$��, �d+\6� ����d*�uϱ��
���$,޺u��;�*�B��7v�����K"�ȳ�B:��6?O�ӫ��ˮ�c�N�~�G���܇F��]�ω�pB`t�0��1���㽝����̬��xH�s�7��^���}=x�xF�;Cg}��n��7�+h��1�/1~ڡ��ٽ鶐dtK��=�S=�����T����;��<���:]���6,P��'��3�v�sqzi��K���kdPNa�����r#��3�64��|���u\�U��E�Wd�[�~ �g���Q���Pɡu�T*Qb����\�$�*�at�_\�`ڛ�\Ǟ���~����Q�>�!	��-�@�)���d��T�_ƫ�����z�x\��V��/3�q��]�]C�/V�x8���?D�B��by1P�s��3p2�
�hQW��%Qt�b3��y��<�m�x�12�fBDN1o��IRr&�_�L�*�������@Uw�΁"��簽[���O�����%�wE��>T�H��wS����&����q�ȨY�sۂ��ؤZ���3�m�U�Ur�d�#�az/�����UX�Nk�9�g��Q�o19!��~���%�̡��{:�/�DC��#8mfΩۼm���2�:	�x@��O�kOC�ݖ�I��Ŋ���9Xͅ,pp)�5�{@�]ZK:�N���7�Rec�ź.k=��;����� �79ܡZԦΫ3h�
���ĺr/�w�Ծ<�����$ۣ�طE��h�C5=X�`�z�3hJ쪡�N�UN']��nzpˑ>خ�Mq[Z�.*�	�	x�\H�ހ(�ͅ��u����)Ì�\��T��Ucjb�w�����yI�o��u�1^�0Ğ~�@�׈����Ei�B��ѥNM#�n��9]��}�nu\��x?>2�\y�[^��3��2��Y�Tb�H��7L>8s�����٭v���ss�����=7�U,����d���c�N����}���� .�t�8O�^3��ׯ��B���0d���=0�q	��e����s�O�_�S�~�(?�Afd��Ȕy�@���=]' ׈ɸ*��^3���B&땦=J˜���������׾+������=n���}�N\1E5��dR�\e}��ͬf*�}�i�^�E�a��v�4�N+��`w�"�{g����\*1�,2�'ƪq^ w��w,�z�v%d[�׏��ݮ�Y-�zj���eK�)��{>��c�£�Tmj��A�%3�z��xz�������賛C�=]�]o%�S�te{���{�����F���v	Ա�d�'�*�X#!y:�F�N
�&�JV��%�|Y��$o=Z��3�� Or��Z�M�N��:�+7
����ɳo�;���I��V�<TsB���\&aħL��/g|+�F_�T��-*���{����yj^��~�33ʝ2�l�{�,8|6��j�x�Y�޿y�s԰\A����W�Ɉͤ�h��0;x��.�Az]d�y��޵0!����Gk׽�9C�N#�P��Ț��f�G�o�V����*z�w��l�J�ԝW��{�_�l�X/TT�W�fx�Z*G�l�KCz=�J8���� ��%W,�{�WѨY���vf��%桂>�t�|�W%w�`����Ԛ�-�A�i��y�j���z�b�=�Kׇ@~�
s:��2S���["��� > Ul����Rc/�MgBy�'۽�J�f,P��~����gר�i[������5�\I�|�\E*���Tg\� 9��8k��"��wo�u�.E���6a�k'�Q�t/ə��ݙ�u>5�����������������8����A㓔��Lta�
�S��pub%�w�Ƨ2vD�����_������m�.M�X+�l��q�/?o=w�/�қ��Yp/��z�g	|��_855��>��tT9���p�s��yux�����>�������?1 ~����a�g-�l�_vzlc�$��y�כy�@��H��gӰ�ջ��x����a����a�,��f��;�W`2\��;�\���^�AK:�l��=�=ÅuN��F��S��������O�Ӳws�J�5�f+�\�5���=X�D�RŰ��I���&�~�~7i~�ƞ~��^��Yν=c[����7�F3�:*���x\S/��f�d��p&�/}ٽ��*��q��C��/�
��ߚ�Sq���E��.�!:*�.�o>�>�p�=��6��dKc ��fg�$+!"�1��0���M�>GH^�� ���2��y_�G�^�,�p����/�*�r
�pW�ܟ��!Sk�5�a��Q�2��?[�W����{��SD{�BG8TT�ѥH�����w:�X��g�.q�{.��ם�Ê���a.U�RQ�Bτ��Uib7�hbb9й]��$z������z�Z���.�u�2�t]e�=gt�E�g\C����`i4J��s>t"ю�{1n^��@r����Y7�>�^7�dPoqsp��ac��\6���3��*��VCU`4=�S��|ji���ǫ�X��q�1�oQu��H����j���w:�	Mz\��^�i�܋�O��TW�r��_�˪��~Y���4"X^�J�L�XM�3��m����	��v��>i{O�״Ddӥ~����F�j��CA�*�eKV����&�h�M�x� ^L���i,|M{]+�.��
R�`8¹0ma�a�4M.�:�+ ����
�Csn�q+��������b ��<�BQ�MИ6#�3:�צsY�	�UӲ�P��pS��Z�}ۊ��I!�Yd0�
�ϥ��d��rN�l¸�M1���q#�S�q�:`��Q^;h[ɶ��	�	x�	]	}�d����eV1��s�	�S{O.4�6$��9���/=���&���+|���q��~�k�(�"k���!��4_�VH̥.q�����kE���"}�����%���$_ɕ����2�ю�:�����a��t`x]�ω�5]�{SB�ؚ�P�.�Y����9Ɨ35�=<�;\T��<��uc������2s��9�4Y�{:�x��P�6'�^���u�M�ĩ�4�3[�*��#��ݵ���%5��sx�cF?����d�� z�"
�]Y4�n#^E1Sp�)�}Nʗ��0{�(6��U��R]�C�Z~DHW��W��>�x��4�W�T�c0g#�+��X8%rk͕���k�CU���p�����;���� �vF!��)�����ﮕG3��Hw�y���~4�s3�,�Q�Y���?f��������EHPcw����e�f��!I]iC����
�]��o��\�R��%$��'u���ꎺ�����Z����o^��(nb��]bil|E͠����Pnѷn=�7ܺ�{>
��c}¶��f��V���qk����p�;���ˡхci����)`����𞪱��v�2����������?E�ĨO�_<F�.ݩ6�4���fyUǍO�1�Y
�������ۯ��8�*�¢v^���Y*�;��XzF�n�vݛ`�$�S�� z<yd�)KM�~����'����=]�����R$7�~ɨG0���UX�^�L�	9������z�޼�����d�"�����:jr+��R`�Дc��wS���n�կO1sK��O�{���o��y�$ښ�C���L�ddW%���(�̭����^��Ng��E������^{w����u8��*�ܩ��Rb�3�q�$����/�FvX���A�}G�#$��y�g�����ܿ>���p{]Kj���HT�q�z�
�W�WUíۆ1���n��^��§05��9T�\w33�{������~�����U����B�t�?'=�g�������u�U�p��D��zaD�9��<�.w�5ߧ��/��)߿v/���۲�r���Z�r3��^C�6����J]��q&��kW�<���v)}�0�P���:��>RND�<�@3�i��p�5["S�|o���}���}K�u5`���Zߺ�>.YqN��3�5A��&�s�����E	p�el3���C�����:�"|�����4���J��-��P���i�^Pg�Y�B7��$�Ny��OM�[g���e�����"�3�r����:򌾼W4������s�Y�k��(�no\ϼ�g;�0e�耯xE���?R�HTZw��U𸂪g�n󢖩�L���wV穩2�&nO�5kA�jZ�����B� +TaD��F�bp�����W��ĒrI���0`
�����8ܟ:Hg��A���.w�O-K������Z;�w�z��kܽ]��<���0NS�pE0��E�t���9�����i⺜f������W���r�kE�Ύ��lę�QW9m\x\�pz�DXX^%Ng~��(�k�y����$d���ݠf�jOtT�뉩�TaA����u-����ѣ��s�a��,컹�^GV�,`p�&�6&��6�E�q"W9����>5'��-�A���������wۜ�nX���5<�h��3�I�L�n�$}l��ɓ���މ���?�$.��|_K"sZUgAƨ�66���k��;�QS��Ϻ�ݶ}g�D�l }\�� ��: ��ې���S
^.�[�aY��͉͇6v��)"���t�)�76ej�]s�&�b���҂�b�u��F�Ld���rn�:��@vJˬ�9W'�Ζz}���9�����z��I3��g5ǌN}�������c�͈��/��Y�Q/'ޕ^�dnE����l¿�����̺L̍���9z���휅�P("�Ndww{�s�m�/����Pӳރ�'(<���nT�ƙ��^��x��'�	�����[�ӧ�Ǐ~�����z}�<����Nˡ�:]`yJg�L)��Yp�����gk{�����a!\3q����~�7�hn��%�Sg�p_�S��Je#~�~�ne���Vi�QKdK���V:�5^��Yν=x���(z��*=�Ί�6p�M��WEM^���C��չ�mt���=.fQ�3:��Y��Hܼ֕+�3޶U ��5�^֟GL#c'�gמy����9��U�S�) �|�e}�I
��.S�&9DS����}�������=��ѻ>��|C� c�'�T�1���Ig����1�� ��Ո��m\=�`OP�8i�~5����9�ɦ/ψ���S;;JF}1eE���td�-=qrq�}�c�拺���ߦȨ�\W�[ɮJ�����3륕g�ʜ����qvi1�[u3t��.�Ի	Э���g%W��;w$M���7�Û���$�79�;W������N����R{��T�+o&�fT�+����U,�t�L�i��Jq�ՙ��Kk�[��ڜ鞦<�n�VZWlC��SyEL��Ϥ-'���*�G!�������Fv��3�^����f��O�����T��b�8wj��ti���j�|D����2G�h���N�ѝq|3���M�a�h�;7H�>b�p��ٛg��miS@��茪�y
�l��9�0B�O��Υ�J����<��D-�0�ζB�@�Mze;.BD���s퍧qf4��
�Y�}��NU˹�1F�VX�^��h�L
��֦�3m���} E�h�Qͼ�}>s�\=>�"�Fx��ce�l�~��9�/au�:��&��TBR��)�pN�U݃�M�D�8yfr�3�gUР�З�d����X��i��nT��K��E�����v΅t���=U��������k�(=�]����p�C${�-�nq0s}/�׹ٞ�Y&}YY/�\rE�qz���ˮ�c�N�'��{�s;��X�7�v��{+�L*9�R�^jɷ�8!�:����m9Ϻ�P�ԧ�k~/Gds>�����ml��@Loݷ ��`>�h訹+�=-ܳ�j��gY\��};)ej��Xq`a��\�ؑ	ӄd��]CHfJ�o��o^^�Ӹ�N��8t�Y�pI�[dTaXs��g�^��c��Ӭ�L�{H��)�����Z�t�Aҧ%�2� ��=s��;��8z��\��f(9˽g*ml"b�b$oX�W��t+@Mb*�S7G2����j�B��TOECof��c�#�������|����u��+��>�m���m5�AY�͍%qg8�!��j񦲆���4l���]�ڸv�7��T�1�#�)�ʝ����e��ؾT]9��Wn�Nޏ��ցY���i�:�}��-�K�i�w��H]bb�����j�jqb��YYw�;V��ڝ}gD�4tB����sF�6���'1Kvp�gܟ	\��#�,�ܷ>�������\���oL̔3,�Wӎf.�z�
.�)A�._^
$!.��3�_weZ*����G�3����PY��Vq۸���楼�> ���]$:U"6�8�$�moK'#W�d�+z#�e���Sqރ����r�.I��]��r��y���[n����D�S5�@T�{��������*r�]��{L�����v��=Gsi�Xҹm y-s�M�l����e�.�F�Xr����� Ԯ� �w�z�� .5�z�XT��`
�+`CVa�o!��{v�>v�j�1]=xt�n�~���_5���[�vnu��WN�ξ|�;]�0��kt �m�Y�/k��Ύ�	�����<�[�ˍN�!�����Թ׼�.�3��7׮��S[u$�yԐ/�C��n�!sf�{z��m�:�{;z5�
�"�J�Z�;�P7�.	���u8���9��=�e%o\�p���vb�49� �������q�K��S�x���f]�g�C��Fk����(,�M�d�K+6r+��SU����y�zt<7�',5!�CVRUn${���}�=��|i<ӆ��[��N� ޡj�'ܰ��f���f������@��r
;��G��͖`_N7��=�O�Í�M�iCg4֕�pe��)"���hݻn��I�%_Xۥ ̖��j����V&�	^ͩ\].�/#�(
��R��in��\��QI��e�ڼ�tgoʯ�����c �#�g��'٥S�q�V�Jyx��
ۻ>�B�L���Ū��'!�=�+�}���5,ƞR9L.a�ǒ����u�_ \y�滔��s��Zt��a�X����@\��T�	��o~�@:+`x�f��v<�4��we`����|��h룷�, e�:�w;�GKx%<9\���k���}Gx.�2��ht��j��fF��$��.0 ���F�w!Ϩ�-Q�hA�����T;Z��o���7{�NG���/��(W>���������,̆T���dR{]�tL�*e$P��R��r(���CIFE)���%2Dġ&!@#��&�h��u �$QD�Lh́���wn�Sgut	�	�i����n]�)ѐ���R!��� �dA�Hf��L�EΠ���#3@a,�-(��M�H�1�<nID� �����˔iLN�S]ܦ&@��㻣4��JG5��WD�\�q��v��D1����˔��0IQx��P�3.^+�$��Q������Rb��B��4�P��U���'���1u��nν�V�b�j���o �N�]�����u���eMݏ]G�g������"W!1�]ȩ��Fl}ќ��?B���p�B�\2\On#3Q�����T��V\��7jW���`꺿��&��i�H�:^�A������T����QpUJ����F'ʓ9	2�����Q�3ꋬ"�a�6�y�I~���c? ����l}m.���C�e3�jmtF���P��T��Q���.��o^���qM#�թ�g8C��B�@**gdj�5K����s���v��^�0�hBK'۞Kt<�a����\7����X/p��i�*��W�?m>�����F�·��~~[��]�f�%���Vx�Ϊz=�8��U>�wv��dӫ��W�xl5��B�q<s��Z�τ���>�B�B���u����/���
��ۺ�f�՘|����X.�]�t~�;{2�ޛ3������ڊ��C}W��j�0���3��D�;j�b�1�J�ͽ���e�?p2�����D�sFz٩��{�Ԙ�VvB/�g���Ɯ��)�� ���R���d�3�2y��/��D��Fvn���^��¡ߊ�g$əw��T����*��Y�/�@�ɋ�"�
vL��CNG0j�:�*��4O��m���wj'A�`�biu��fͻc��݁:��|yp4����������3E�Gs&���[Y��q�r��5+]��$�{i�U��"Fh.�\D�tB o��;����A���h;|eUZT�u�1^�I�~�@��%���챵��rٸ7���9׸���h�>;99F����fP���ܺ���ѝ�q�z�
�W�WUS�۹������+7��T]*��!�.042���GU<�s3:Ǿ�K��f�6���WTlQ�����Y]����^�u�dת�g����kό.��L�Es8�uNsj�td���긩��*n�x֩��m��>�=ۭ��>1q�7�FM�R����-�5�B%T;�#�BU��gv�s^�vzsr�OM�[g�C�tC�������ʩC�(��dϊ���T�ߵ^iQ.&^�ˊ��r�E*�o��xE���<=�H �Q�!@e�O�U�^�y�}5y��5�<��޸��;�=/�q�1䊚�����-S����in�!P�J�7`6�Sس�w�Y�]����|�B�f��!躮�q�nLy�CҠ�/��s�����#E`
���MߢY溩R�y��9��W�d�C]���>"�&=uҬ�9���8I�������%+[@O��^5��uw&��N��TKw�ieN�ɈZ�ً��<�I>C�p�ص���v��ie��ԥ�yjV,����������"���+��&3�ۗ��m�s���N�����\�G�/�b���1}ܙ����yMy���0�׶i���T҅�2�m�mʇ�g^Ȃh��ά�Cߪ�9�P'��L�Zbb}΢�$r���n��������u�*��ʸ�~�׃�� ���]�mi����j��D�(Z�=
�ǥU�#�W8V;�����B�v=C�?J���<�m���ul��F� uP�����!�1^���7�)��z�H �ofR�t4G�c"\�uT�w3�/!NgZ���O��-["�+���{�vx�\N�3���SU�ۯ�-Կ�R��Xgx���4�.E$\��Q����\I�|�o�^��={u��vU�����Te)����2/�pمk'�Tˡ�L̍�n��yW�4#��ǕmUy���\�s|p
��BN����',��0d�7�W�����:�7;�h���N(�׷>�^�NRQX�k?a���������B��ʐ7��d����u�e�)��ۅ7G�ؠ*�/3��J|\��x{]7��w����KyYC3]2�p��>���*�����~�uƄ����+12��ȓ��&⸬u���������PX�G�:pEn��Bs����L�������WV3-.��}�Aӽ:T_�-ΖCѕ`�5���չd͋��$i=J(�I>1Ք ��x\J=�[�*&K�r����е��Q�6�f�U��akB�ގªv�C�_��N��58��xvk|U��[Ɇ
���7�w�_��+��> s��U�U�+��R7/��J��3�Ҡ{�E�p�f�ٝ9ݾ��#W��Q<� �1� ���H�Lz)�L ���\8�O(���B��5��m�/�] �*ggQ�gƫ�QT���^3r|�!Sk�4e�Y��D�:�7�	zN8�p0�蝬�B�ˈ���3��J�Hŕs��s����̢�Ta�����'����k�:&˾�
�u�e�v�?N�<�L�[3�L͍b�w�|�(�I������W����׃=���h��T�x�+EûWӣL\yT���-��������^�DE����~��r���z����NG����-;<k	1[8���������4�᪰��W�%�塈�$�������r5&+ըUČ��ǲj��.�s���9.C�&S��n���U�>����t���׽N��u�FuzU�\�1F�VX�^��h�i0(_&fu����]p�Jv�i�`�2��τ����4폂Ll[g�~x�^���^�o�ѫ�������ȴ�:8۸��ȳX����"��f'.3 ��-{O�姲�m�:��M��S+ 2��i�.\���ʹ���ǂ�4�q����]JV���q�Q����{�ggs��K#�x!��[�{�f+]�P��ki��c�U��n���.�t�s��a���WD��N���k3�d����dzq��OAU�o��s�uadtI�O�WkۉÚ���_OK�kr���ʪ�*�+|٭���ʵ?M6�E��~ ��^�a�A�qy��W��wS�i�rp�龤rE�����[^b�'��{��3��'����L���4Q��݇'�s�\�u�S3��:�P�ԧ�k~/Gg�ϧ�1�����/�\�z�y�l��v���<���n�\8N�!D���1��u�OU)�4�1�B����{�nK���8GK^��E#��j��|j��T���c�1��"��uO_q�NQb��y�mj�׃�+�����k��?iL߾��Aʸu�2�ȵ>=6M>U�Sܯ՗�I�'��>9y����+�1M�T�|ڸ{��p���H_�� ;�3�5NA�X=Po~�B��c{�����};�Fyz�Oؑ\7!qm������wӸi�ʦ'�
'h�9����:x�{�c�e��X.V����J�<rH�^��H��.y������~m~Z�޴j8�w�jSY����e�����wӥbƲ�pu�ac��Jk�K*�'�f7��{��L�nMZ�M�Aep����n��sXS;>�Z�ĄL}m��WC��ـݦ��v�����5�XI�YN;=����C�p�F֐�r�����<�ٙ�z����9�WON�[Q>�Sb��+G��[�� �>:����ٍ�Ǿ����w۽��UUC���d5^ʩ�?J���V}����52��ꧠ �2�T��Rk=�v�UyV��ɓ��UU22+���툗]5#w��z�6��8�����h�{�ߵn�?P����zS���d�3�2b9��U	}�Q��O��x/�dS�n:q1������:�Ě����kh9�����*s:�\����ȡ�D��ge���5��
����}a��n�O�c�7����(W�u��ѝ�q���*�~yW7�X|�e�����n��/|p�
��xzS�J���x.#���c��n�����UÐ�)DP�b��ߺ������+y8�V��g�ด��|MG�Wµ	�μ�	��K�{�;+u�e.�Փ��}~���}�g���h�T&�!�=&�׈ɲ�_U�S5[pQ�8��=�u�wJ�y�%�=���e�nCw�鿱���������b�o�x\R�tWp�ix�<��rΨ��e��3����s�vӾ7k���v+�6	�y��du3���4�D��[����%��)7��D���Ȣ'7�Cۼ�ٺ�.��a^�ŢJ���]�UkE�x��M[t'%��6�2$��ҝDZ꥚�(�F,��r�	w����5%8�q3��1U��R�Ur�d{�/������@p�ǐ����ۃ���V�T���Y6ֆr�[�������5kA�|]�hz����H\Ct�
-�\*�^e����q�.r��A�Py���y���t��BҨ={����Z�"������/j�wuދD�Ds�j\Fƴ���Fx�����t*��/��p>���ٶ�ܕ,J��(���dө/�vo�"Ud�P'������z�)��~-���:s��pرGd�{Z��:��?�;��wv��D�B����Z��3<~��T��;5r�"p3�sc��1;{����X�{�e�¥���l�D��`����T%v�0fze�T�8�[+ӛZ���������_�^��#4�S��>�g@^B�ε&=3����>�@�@>�~ʢ@w�V�}�6��މ���	����e�<a�1��M�m�"�.gR*|�5�\O� ���U�������{���O�ʹW�������pB�ȼ�fƲp_��B����挻��8L�1㌓�m����{/:'ë�{�g7V.�<2#�Z��j�0�TS4\+_W	�9%W���Ѭ�s&����-,����������C�V��F���WSV��4O�;�CX�W]����gC����xow��z���:�c��-���mz����#�T�K�0��l�������0\`L�مh��2�<D�k��8��
��k��N����OB���*k����gn��==�(P���d�;[/`�`ٲ� g瞻?�{8����cI��	~鳨yFK��ܸ��;]7�����1�/��,G3j�'F�>Kv��8[��b..7/=��y�3z)�q\�}�;"Lok���+��^j�/z��zz��PY���`9��!ܞ�y���w[�p\Kjg�)L�yT�}�����p^�F��܆���c{fz��?��<�jݚy�s�K���^�z�*A�B��.2��\b3>A!Y�$\��Lu��C�YlFW�#��mU��RK�p�!���K�N!i�C,)���s7Fx��?yRB���U��B�_h�y���:��ac��;Y4�Ǘ![��N�*EČYQf��ע��,��l{�#l�[��D��p�+���p�+.�b�n5�ʫ� ;���>��k���<�)�����}�W)�=�fS��o��[�qZ-ݫ�iѦ<�ĵ�>$pUU���~1c�=��`�Ɏ���"h�� }��<�)�mt���~���X&^y:��ļ�]ݡl;RЫu�S���u�V��c��)�}�p�pp�[36n�O$q;8���ރ�D|^n�Z5M�}=y����b��9�P��`��'9[�[܇^|�ʝܻ���w�����T��؏�@��N��H�!���.gfn���I�E={�5�}�L���]`:�=���Rb�NA����ɨF3���d.���? rd�_��We6*������wf�?Hp������C��j:��BP�Ϻr��/
�}3�{v���� U�����r�����2m�&OБ�	�W,����c�Tgn%V�d���7���م����z��e�9}��B���.9S�q��溟	��~"�WB_L�N9���Зe���V�Z��ʋ�~vR�6����)�/�gRUlV�b�o?e�}��"O�l���h��j�׍�]WL
�|���A�����e�å��R9"��/]z5ї]^�^��M5K�c{������^ӳߗ/rY��o��࿈�����y�s}U�H�S�5����g��"E<���u��^�����;�Y2svܹ�t�(u�=C]�g���J��k����J6�>���9��>�*�1��:}��������`�>��uE�R��i���bm�f͢���~�����N��y|��ݛ��'��=�n�.<�c~Wt��O�����D߅%6zg5��H�ʆ�.�ohx�Nx%���e���k��.���Y%���2�1_H�,���6�1޾JWZR�������O<��d�|�=�kcכٛ�3�0T��!�vT�����
g���NUïi��E���E �>Uٗ�[�n�vͿ�lw\�s���jJp����%qV��u��g8C��R� ;TT��Z�M,a��@��%�p�ww�mއj�Z�Y��,�\�h��.!�y]5�۸~��4�ǕLO+��6��k:{�N���8�O�2�S�f�J��r��Qz3"q����廻Rj}��Da`�>Sxw|�]V�̩��[C���]���O���2�,�����yS9#�6@�ׇ�=�9b�c���M:����@�$�sp���W��g���J���&���^D��b�K޸m�e���\w�]Xp	�&Jg���Id]q"W9�=�.�jLV#�/��~�����:������^�O��,����V@8�|����f|&Ls�d\W%��
3�ai�}�c��1�Yx�������l�m\�ϻI�?^�.�ҧ3�I����by�<׈���z�uO�4���o|�D��M�g0\��4���4����k2�_��u�����s�����ӯ¼�PuJ�����ʂ�/��M�lB����b<�
9
�]��Ѣu�1r�l
z
�۳G�(��3�_q�Ԣ{�7VVs��Vv\Qp��SR�]o�Cͬ,���4ꕭkky�7��87w��챼��;��ZtZ�wm���i<�����u_LD�Iv%�Լc��
�Ivw(q �c�l�z	�(�ନ���]�c7Bҵg���LB:�g;���]G�\,.�EriK�#�(I�f��Tͱ��R��]Fv�ɽ�YF�/�$���g�x�^^�lj���Z�@F3ۏZU���ȯ����[��RRʔ�D�V�B���Ѷ��nA��+�S2Ц_%õ�լ/����R�w�}f�ud�;18Q��JR��z������l�^�q(e���W�n3Cr���'>�볓��w1˔��ͰLeA�Q@��%l��:Ң��06�m�w�C(�"Ř/�5�Wh����)A�52�9��z�:B�sky÷Xe_k��gq���wد�"���ڶԘ�;S�-�J�XC^₆X���G38n�GT��4�m��&,0.w
<>��}S\ȹ껜���1�r����f=Uz�ft�z��tu�Й�9);h���e��H���s&WPX�X�_^ܿ�A΅�����n��bmwg�5�x2�̀�82rHX�z�q)7W��� H_o9��ߵ[ʉ���չV��������Ӟ�ţz�Y��w7�����JwU��}��?n�
�5b�"�B��R�Q�t��>�.�]�\8Зժ���a��e��ƽ|����J�A�̮ڗ|�l�Bp�t�ڭXa��\�5����8���Y�X�Y�����7-�.�]]�ծ�q�L\}/�oMf&��է�\l��L�Ns����Ȱ�=�Q����j�چ�B7�b��T�/��}��w/C��i>��b�l(S����Q7�L5uh�j�9-Q6�W�а���Wwj�Y�U��Z4�t��{���4b\��uf�86.W�ɽ��/rg�l�E��at������+��� �����e�4�cS���4`�9Ҽ-�`�����7B�-��^J�:ݜ�1ذZ�ٱ,"N�&�T�a@e�o
�p�/��e�.�{��^��$�7�>�y��q�J��4�O�t,qu�èt	�*h����if�FI��.�1v�<Jq�Q��e�)��O���7��;�.��V�5ΐ�|�(�]F^�hN�Q����@3��:�v�6�<N4���}�����f�r�V�5U^q�{��K~���F�ᕊ1���"�,���!wn5Mh���\�!DY��l���������$�`�d���lx�Ԏ��e WC�*gJμ탚T(����]�0��6�R{���.v�o��h��Ŧ�^;�Au\`�B�.d��	ݍ��_J���n>�a��$Ŝ�sjv�<s,
�a��ົ�ﯿ���0���9t�����&?�;&���C��FD��r)�(�����v�!0F0C��`� �r(����������RWwd]�wJ�\�J@HD�RD�4��tTbJLX�i������6 ���I;��p�n��b1ݺ6&bĚ�"$Rؔ�e0HƯ;�2$8st���2�:]��;�r���c���LP�7.n���F�RQI�.oc*y��bܹ�hѯ!�W&��dcFwn��狔�����8��P1���#3r�Dj�I����]8gw+�r�G+�����Ӄ�����}�N�ٜT&U*@F䛥<:���T�y�Z�ʒ�ս�!�ưT��6�AfL[Ns��ř�͌�	���o*E�]H�f��v�!�ǉ����0~åO �;�L�#.k���s���=��z���nz�}�h��<�ul*
��^E�N�"o�A�+P���>�Jn��:�7*׻+��%UӚ�]�z�`��{�Z7>d��8��5�2i	}[�L�wc�2I��}~���qX�8�=�&���1�V\�nvz1���3r_|f���S*(,��،��K�o3M��)��*W{LL�b1L�\�Ԫ徔s�t&��D?R +Tc�zߣ�l���n���^�՞���U�\&R�5==q�ܟ$T��h=Eږ�~���D�AB��Ea������� 5��
��g����S�C�u]*�ɏ:Hb�T�z�Q�q��J��9��nuf�_�S�;�33έ�S&4j��xa�1軮�]FsBcpOW��×�h���^ש��MO��l/}.�i��(��<L�ZbL�s��������� $t�^Sݝ�ٞǜ&^�����<f+%�=UU�|�T�W�fx�Z*O��vj)�T��C,~bͯ���i���ڼygE0��2�m���o��b�������1o��+9e:�Ad�t��-��Q���ԩ^Pf�[��'G=�q1}rue�D2�e��|䮌�Q�ػ��L��mC ���	���D��v>�]�e��Q������t0��է���;�ȕ�[;;���UX���������B�ĉ]��M��Ͻ��O�^������/qY�^i�1�N}�΀�S�֤ǦS�p:��:��o{��dc̷��r���������NKg*�h<(g֜Wl�(
־�4��t?!Fr{������ּ%m�����?W�w�J\�=��$��j�8ϰ�g��b��,7�b>���U��"_�ly(6�G��3��Fp^��9�^!�'ke�A㓖i`/�	�l��K,n�`F�'+�����::%x�z���b%�w���3��1����H���Ro��i�t3�g`��1�X�p�q�7���s���uf(be�{v�&�u�p.;����E���]�zn#��)�a�T�G�T�Vs�R�3�mȽ�vjɷ�2�H�=3^GdIת�o�+4.^mw:����o�E��z�*$9��J������=ڷ8����YU�
���Nf{q��Z�_Ǌ���/�5��4�oFM7�*����^[��3�/J��f���U�{�*�\�yʧ=��sʒi)��d�W�l�H�8�8���ܚ	�p��e�t�%�h�cb[��R�lJ���ؕ�}M��M�̨HN��hKO�t����Wv^d!zinږ�kЀ�]w�oR�.S���Ѧ�epާb�BBF�v_1)�{��8v�B��#���.�og�g���w����{��P�!y�� %T�sF���ƫ�QpK<���\�3sСl�I��Ԩ��2�ٷ��]�^xT����&��3�?D�d�]BB�EL��iR"qz�>5]έ��r���f�u�K�����M�=qra�W���θ�l�!�N�/�*g��t�J�7���N{�2�W�\2I�{�~��?�_ޫ�B�iٸ	���$^���WӣL\yTĴ��M��E��V�^��Br\�2b�����mǌ� q���XJ���veջ�r62�z�����**��{�a�m<ʰ7�<6�Rb+ԴU�#%1~ɨY��gs;!y��:� ]!���,߅W-��S*�쎪�5�����z�_��V>����9�G��&���8�ezo�z{�*�(8{�g_�92cY�	<ϥ�u�C蚣^�;g"�O吰�*r����mf��=]��s�-�B���$H͎vg5��L���E�^"_x
����2|e	�OVf^9�1/��73s���c���?a7=7�����ʪ���ح�7pt\s�_�ѯH�a�WL�>�L��cD>��2�дѤ��\�zkh�eWo	T�-#����)�;�}ʭ�̗��K�J�Y����m>M����eZ���W/7nu�Z�0΅�:���2^`�)��(LN�Y[Gؽf^W7�"Ad�l��=\�w�2zz��wM~<"�Ag�#ާ.{�:T�u#�;���F]u{�u��O�����T�J����~�c�;V���\k9�с�a�m��U`��0���=.n:�P��*q��To��Pn����E�^�j�}6�g�sl���'0_Ί�5�X0��d��،Ff��Z�ø�b�e�Q�G���N�N�Cv�\cw�t��C�H������W����ձ�����{����}���z%D��V
��h�=�}���t�<����J5o��:���Jf^d�ؿ3=	�G�:2'��`���+���N��ڸ{��~��4��H �3^��R�+����]�g�{��x:\���WJ^�7<��z�q�\3���C��X-�wӸi46Vs
���R�ׯ9u1;�
��j�\͌���WJ��r���$�E���"'�x�N�ҟP����+�Co?(7��W��+��� �+Dq�CE�~*P<=�}q`���F��>��������ٯf�OW{3��,�����4P9�4�5d5^������1@ymEdHo���5
�j�"����{Z�s�˲X̨��4(q��nܰq��rwv��{,Zf�+\��$�t���'s�k�D�v����:-N�v��a��b�gm�-l��YY}����ڃmX��Sm�����N����ྉ��f��r��vF�I��JM�G�v�6�
u�>��.rp@~���@cʫ	�zg!3��"K"⸑+���:jr��}�/ݳ�O\���,�Y��_><&�n�B��N�D c ���	��Yĉ}2*vm����?_�����Y�@{�ٟ�xfy\�쪩ؽF]U�T�u�!�������(_S��T�F�h7Y�����X��"���W�*W�ǥNI�eM룂��̡WF��ס�3�/�
Fn�b������ǻ�ŸN�G�zEu\*ݸ~���B�0^��:T�U<��α�3��ya�g����.��k�p߯&�w�I�9~�c�;;
ե��E�N����B�c���}X-�__f���.����K��f�z1�`�o0�uBo�c�I�^#&ગ�9w2��c�dJ��Y���X����;�&�Zc�R��7�OM�5�xz�e�trr�(˝���+c<]OZ�v�O����JyF{��ϖ��+�z)U�}�^��M���@�К.n�+7}noKܜվ��0���A��UL�����7'�5qA�2��_S���Lhˌys0�c��m��'~�e!��>=R��^5
T_�s|#���qx�Ӻ�TT�_`̷���Z��_G��b���������ы��v��$�v{�v�ٝ݋�E��3w{�Sx�=��x�3�h2:!��!��p���Ϋ��su�*�����|�-���R�T^:P�����~���W�i�^��C&��S?G3b�zg*�Kg=�Ҩ=��VOu)�<"�ͬ��I��n�/e{���ʦg�s4�vu9K�\���g����Lo8;��X�َ��R�|�����o�`o��4P���ȟ�[]iDp{",A��D�{$��̧���87��ݑ��u{Cɢ���a�x=�T�x�+m��n&�j�]g�HZ*N���zdO�	�{=����a�ӑ���"^:����{aB���n�bo�|��4Y�����`�����U��>����S=.3Rb�[���0�4�S��;���
s:�\d�v��J����9qvS��^�Hq^�C�TN̽����le���?7�F���"��3��|}�빱50�L�;�k�y6��eĔ�����W!� *u�Ә.X�`8l¸�N
�o�F=��ey���\ɠ��3#m;3��|��=x�����x���i`/c�F�g2n����s����V���>��{.k��Y��عߣ�i=��c�Ӳ�q�,J%��,�H��Sv�m���d=�J>)��OT���Q�ߣ�l�s��y~�]�&�e��]HD�T2���!{�Kˊ��om���J�enr�=�J�鲓%�Y�g7��cVLWW;CHn �:b;� �j�εN�=����S�iF>����Ǯ�)t�^03��zǢ5�c{5ߧ���/��ON���@�����ї{�V��SHW
Ѳ7��7Ւ%ƽWq\V:h\���u��k,�}�B�y��x7%��������}F3ã���ʩ��\��FgP�+ �\���r7��GvX�žb�O���.�Y�����y�ʸ�f��1Ό��:��DH�-�C�K&a��xo�7�on�x��8,;+z��q�HZ%L��1�5^�%�C�+���~5yhMD��9�$��F츗��$*Z�i��Cj����v�i��$+r�Bu8"1܆i���U̺�ݔ�)v������������]C��qYp���;���3˽G�Dvp��r|k3�<[�ŏ	���)��6��\�/�Ւ~	��{���;��n�\�S��P�v��/U�wY��K���F:/TB�諐�mǌ�!�kgc�ag�V�m��5�����d�j�~��˂��I���VC ���VD���ǲj����vBm���_�� ����yx6����
'h�JV�Y����Jw��Q�(a�&�(?E�mk@��W�6�k���7�t_7�g��uv�?FǄ�5���$A�[
��zGόͳhڜ`,�J.u.8��fe��9�׼83K�;51��9�����{ g�_t���^wz�Χ$y�rd���H��>f�⸐���z��1U��,{��㚅Qw�wq�����n���Aƺ���&fu��L�f|$�s>�E�]d1ޚ�;l\`��D5 ��/�|�κ������՘��&��p]��č�vg/�fpL���(�D����b�d{�*2� ����?p�pUo��N&�M������ʪ�*�+[1X7���>�5�x���<�� 9�In��sZႴB�Ú,��q�K�t���rE�qz���ˮ�c�N��i����]����~��7�p�㺧w�l�9�ZXhy�=��#=is�j:���F��ɯ2%�+-�EA/�<�O^/^N��P��|����7��p\A
%���x�#2����>X&�l��wOD��-���=�;.wq�R���t���Bz}��*}�U*�u�7�>~�^�/s�^穢�f'�I
���Lz)�R� #�.����~DHW
��l�C����^���D��>��ٽ},����*{���qr|����N��ڸ{.��N� �s(!�� ��Ȏ��q�i��o>YG(!�)`Ga%`�6�*��R{˶Sw�!Af��������f���[���!41���V��c��P}�y�hN�.TZ^��0J	Lu�^�o2�gv��T:ղ����7��^PHɻ������{���ki�Nmӣ���9���������5Ny{�7<�����9�1�����0ՙ�I�����{�2���اD<ʘ�W
�(����nR�pj�V�C���I����$D��z�䊳;��E�M�o:2iԗ󻼓j&�y	��]��O��>��\H�Z.=u����)X7�L��c�:���|R�P�`�7L�M�N��ͰUUPS�Ր�{�ʩ�2����ڊ�o���=�u\e���x��L���u�T�<����צs�Ϙ3q�ȿ��������]t��-�:˅>	�{������C�..���/���{u;yU8�jj=��	�wL��B^�yO�@Ǜ���{���;.g�3ix^���:�s�US��˪������\��I�.N�t���\,��^ynu�(]	\�
3�ޭ9��`y�P����U���Ǌ�~p~Z��SA5}p^���b�M�yqw�GQJ�"���0���B�0_�[Jx�1�υǐ�uK���{_��Ϭ8h�5���j~��{��*}p�xR�9&�>%��Uʪ�Xm~�K��^����)��G �j�j�m�'K�ŬV�u�
~~��]�~�w�`��2t�]��������_
�Ն�l�R����wU��j�N��t"�dtjXceq}Ykk��ל��i��5r����9��^C	���'\"S�݊�w�3C	>�:�8Ǣ�zCU�5�\�f����3�-�������f�FM��LoC������οwO��S��k۷ �b$r)��e�n7~��ƶ�Z���ΎNCγOD�E����S��Ne���y�k�!X'F�����bg<��Uu.UԪ���xE�&���|����|��O�'k;wX| ��Q�p��ɠ��g����f�ǒ*j�����K�]��&��s��k�.�G�T���j�(�Z�3�R�YNy]WJ��r|�!�л�t��s��9�j�x8��\ﾧ���蝬��<�����S&4j�9KH��$t�����w��^�=�Ҳ[�Hv��u�	��6��K��b�<����ei���:���g/b�lq� 4��ڇ�Ӎ(֜�9��%O@��ⵒf��U!�EL�驞f�!Y��A}�;����M\�co�Tʯ3���)�ʫ����|������y�ܼy�+;��/{d9������A�]�3�Υ�8?�ȅ[�a=c����\G������{���{����V�k[o�ֶ�[m�m�ֶ�Z��m����:�mkm�������V�k[o���k[o�ֶ�絶ֶ�ն��۫m����[m�m����Z��m���������+m�����m�����m����m������
�2��L +��� ���9�>�@��)R�R�H��*�@�QQ!"(U)P�!"���I *�%
�U)*J��*P�*"�T����"���}��I@�I*���H)U)$UQ%Q*���i!U@���UR
�mT٨����"����UI*v�8���(��)Tz�%S�R���l*� ��QQJ�J$��)JRR��]ja-
EB�H�����J)Uu�4U!$�k� d�B��V�W��Ո�v�Pw\q�֍�J�m��D4��@5#�0R�b��EZ�ʠ:�F)��ETiU$��  �zZ�рP)kx��(��(��:  (���׼�EQ@P�]�QEQD�pc���(�,��QEQEQp��@h��WWI������$%H���iS�  g([=�S`�r�����]\j�]������٪i��d�t�v]+4��!40j��k����l+�֩�k��k�A�-hh�B�J�RI
���   w��GG]��N�7u:�ؙU��빩���M��*3e ��Ա�B]m�N]�(i�-�]���Ӧh�U�Jh�m:]��lr�]�Q�I�e���   �/nڇJ�X�kml
�Gk:v��Fv�t��U���!�tn��5�Wj��*���wwj�*�t2�҂�A�.�j�U�A���������DJ�x   �ؽ��uf��s�V�B����c
;s�FYm�]ۺ��7i]��5dl��n��U�����4�T���V�m�*p�.�m��I�
(P��TU)Hx   {���ۣ�FwT�M:���hN������X*劦��n�qڴ��v�9�tP�[IUav���M�����v٨�j���H�U(�A �::��� ǵT7���]�v��M�4��К�@u&�9su�P�.���uv��nN���jӶ���]��uܷJ9T�RLu���TI$�J�-�RU(�� ��z@n#J٢���h���T�cj���֛*1E���E�;�:��uJ�����\ܧ6:����̪��4j�*Q6Ҫ�R��J�O  ��VT�l#�Be�� ��6�T	��֍Sd�*@�U ���ֆ�k0`
h&4m�%\ ��*J�1 ���$�* �T�&$��  O��P   �=�&4���� M)21U5 �XM�2� �@Ruf�`h��+"�@Y���{��a�3�o8�$ I9��@$�	'�B!!���$��	!I�@�$�@$$9ӯ���\�?��e��Z�Y2�P�7�h!�ތ�`�PP�v7W���3�1���	ˆR�o@*j�ѶV�m�TfKƦ���=�!�W�P!�#4a�&��K�S��p�mX$��p]�D�H%F�c�ң�F0�k�R�:�%C�	e�{���O��,�m�AEX�j<;x��vp�$��ˑŒL��r���x����U�Ҭ�.��VC�*V˱��n�n��⵩�B���ób�����#r�e���� �Ŵ�ݸӤ�	!@��P1&��P��v���UW6�h��E怗�ek����j�R
�\[�Ư@pF[����ZeAJ�l�]�<���W3E�n���Q�`P)�[Z)E/c��H�7��8&�ø"������i�[������$���d��i)�.��*��lǁ���y�ΗC�J�P�)��SVeq�Y�L�x��!JDb�Bk�)���ᣳI�՝KE�wbX��P�� CL�9U��/k.��
�W-�����2<��Ǭ�P	nԣ�36]c�� ��WWJ���ذ�&�r�����u0���j;ݗ�Rx�+#	���Ր ���Ӛ��P�0�_�X�R�[ƈ���Z�c��v�;ǎ�nH B^��w/E-9a�̦�J�n@�Lԍ��9�ׄ�jJբ�ƥ����Z^5�Z��-��mL��\�Pj�0���ͦ����,�@(UɁ�r�v�a�L�\'+d��{1�[i�f�X�HRڽ��!D���u�cOږ��n>��ؒ�W�Q�J��������nı��6��&�CI9e�M�0K��Ju�3r�T�l,��BWc5��|+cmg.ER�^�+C�]��8,]���
j�;,F@#�ժ�^7+u�FV,(Z�*�q�Z����e�Ԙ�j�K.�k�f M�n���Z1��q=$�e�����% �.�/�7!��ڙ��RdN�l)I$,YZ(����g�
���@F��l�q�ڿ�<�@e�[cU;l�:(��=1�;�v^��M�
���>E��Uj�X`�I���7H��Q��h}gr�ںd�E*kL�����ٚ�c��W��Q�! �sr�<�0n
�AP��".�gvAf�*�j'3s-��[�EE	w�$�I�(C[����7k)'�Ca�Vɖ��Y��N(��F�F�8���Y��T���Ү�$���*��m��[���G���5��Mv�;Vəz�ݪS^���$�ԥ5|kU��^���zH4p(�9g5-��E�]�q5����q��v0��j���,ƏE��Q+k�m^]�5����*ـ�Z��i`4�i�P���lC{��V��z����l�rYx�Gjh�9PV�d��ck5	��N�Ƈ�n�G��]�仦
s7d�/�!X!�g4.��7l@J�c�sP���D��fU5G)��U�K4�Z��������)ZY�R{H�Q�Vk���&h�R�hpϷ�m����N���v�Cq1n�+���r,�Ϋ����*�K&7�YǕ#˦�i@��x6�����	�/e��#+�M�=BL��7oq\�Y�u
ʶ�6�]3lM�ӷ�4�2cSrÈ-[>�h����S��וr;��^��RS2�պp:�I���$,P�b�Xl���+E�o.�.TT�*�m��eS�u�y����Ąb�=�>!��;���\"ޝN򞂝d��e�m�]�ӵ	�S�%��ȟ�a����e��n���p\�����Jw73P�~;5�&p VJN�Ѭ��0j��ו�^O���Dm�ڒ&�(*ݦ"��:�k4��b��.f�,�)V5��o&�cr��F-Z�h�Mx�F��p���\�+d�n]�GM02U�V�pM�i�F��sB��v��Қ,���Q����v-�a���zqV]�J�
RZ9Z[�G�%[�,����X�ec^�:QdD�z�㰎i��ܸc[q7V�e�A>2۳�,QB��2���K\U*��إ�E0��z5�uH����E&ӎ^�э)�4U�jz��M��ÄgUݧ��L�v��/+j��j�ö����u�*H����܃@�`�2�w��ᶨ5{�`w�q�B����o\m64괪ço2��9��F�V];�ε�Ԭ؋����l��D᳚�[q:{M�jČ�Q٘D���k����Җ�1�/b��V�nΤv]%^�*��!�%�N[xK	:�]��׷�;��a��kW�ݣb
�_\���zQ��cw]��S�N�w��P�nW:o�؉\�3onλ�X�� �։�,jd�֍�����^ꖢ;Xd�Ryu�Gl��tۙ��5�ݯ�D\x\�K-7��sg�{��Ә) �z2�Ym�2�4\/M�d�X3VK9ZP��%:��Ζ�ոn��Q�\�ݖ�+�b��Ud�0��ĩ��x���-��y'�G 8��୺JM�!W�j,�Q�(-��'5[�m�������6���Õ6""��44�h�����a�2"��"�պoE�X	G�v�M���p��T'(�P,yOi(6!B;��w3kt#�K9nK:�-`d1O^Q�IX�q �]��a��j#`;I��߈�P��@�L���,aӒb�>YX��JDo�IVZ8�H���-�2���G�-��)��w�)Z+jd�w3S�Rl@�vb`Ĳ"m�՘Qaݪ����̭�'�rD�W���yP^S.mb�rҋkZY�YW��I���ȣ�kB*T۫��3,�	�F�M�Ơj�rmn\����i-�"#nL��6*���H����BB�X�1SS+6H!�nXWn�P:iS�Ccktahǂ�[��	l��LJ!r��,��H�m�Ds"ʈ�72G`:���d�6�:�2�ǵ���[��B�����́S`���B��sFR;Wm�*֣�F��U�r�w`L-b�*�{(n��w�pTP^	y60�@�hbf(�'W���;����k��Y)]�G��YNmH�km��]X)�ifLL�\D��.�AT�c�Gq�5mji�[WN���m
�d����BfXqUʋ1�Bb8��e�1���ǉ^��,P�Zc�%)8���L�� ���e��q����9
�!�{�.�ͧ�~45�P*�FfZ�1Z���M�AS�kc���{�,��e���;I6����&QV�R�$
T"��Y8J�D:�̡J5��˥� ��˨�R�r^jͺ���ňm�<�F����p[���t��#�^7h��݃�ܭR�.�M}s��5���-+��W[Vm�+ai-Mj&�
�fѢ�e�k6֟��T0U=�u<MJ9 sq�@5��l��E��!�t��B���2�*�I6���LZ\Z 8��Ẹ2��C^��L6����-&�է
R���+"��I��H���f����y��2���ulR��%�'F�<O�۾[�V�*;��-!�ו#�se�ջ�Wi���z�n�N̓3^.ai�P����IQ�!��#_�S˻t����]�����5�m�2-��u��.��r�f廫�g90�Mɶl���%W��=x�v��m:W�����!�#��� x�n���2�5��0ЅYڊ�3	E����2Ĩ����J���6�F��Je�.�Q�2Ǉ �7)�6�U��R�ٔ�2e%9���a�Zwcte�&0�LgעI�FD5�Y�����B�V%n��U��Kx��l�*5WÀ��K���� 0��Ԩ�ۂ$���r�
W���շ��׃a7�B��z�[1�TT�y�2�Hc�(��Aݜ�3N���gH�<����m�B�fe�����^P5b�nLt"�a۱*��n��s���r�����ۻA���*���u!�"�j'Q�Őb/,nD t�LW[&���Y�q�م��	�������l��[�ז!�kY��z�3Ph�+w�ԹA��+�q\S&{EVē���6-Zw.��8��9|{��V���ˢn�:t�'l��[������`��X��tr�S�g�3f�-ɫ����R�f���Ԭ��.��ln')�6��0���@^=e<�o&9S&��i�Q�@!w���ER��P����t�1S��[t�Y��C��)��rLƮ	n�m$�ȗ����Yu{}]�@&�`e=v�H�6�-�^`�i��-��o~d�I+5z�J9��^�Ү^�TN$����J�1�&��� 6�Gu@hzk������+ZP�Y{P5� �"kY�K��TU�Rơ�Z�en��F��N��*�Lm8��fl3�;D��
4,$�ӥr�hX�(��*�o��B3 �NH�	���,��9�E�@R�n��FA0^V��/7"��8����bTZ�˱�����/�MKwx%��m����eX�q�#
y�:��.;��N�v����&��N�E)�J����͡�	L4�w6^C�i�yl����V˨tX��hC*�c�K�Q�����Ky*+*�L:���7�R�n��+)��M�����lOi�d��#t���U��q�IEV�K^A�ְr᣷�0��	�K1]:եhc,b�I�엷Q�������J%��;`��e�n1)�;#�-j�ᐊ����+�i��d����+UE����[b��t��ܥ�#YQ���[���[��ah{u�JCWmd��&������n�!P����`e��J�V�If�M��J�4�Ûw��ܒ�o-���c�"mB�8u��Z��eY�wJ�
i%�&��Y1�G!�D�T��;���b�ѱ^�09�I���(g�5S.)��Snc��K" B�S��:˺�ˢĔ��JmS�E̡Y@E6üٰ����f��b�:��j�:��d���6������ѱ�X���vv���`���xУyxU+H���9��f�r������t��]�,�%��6�~W2��c�¶Tc�$`�r0x*�ڈP����o42�Bm]\����fMU�d�̎C-'۔���2�tv�
��O#����5�b��aбҫV�#�"zѻ�a����jm^�Z��K:Ϊ7�Ÿ���܌��P�F�\�����I,�s\�d���f�E��!�f�ݚ,kXݔs���S���t��"�3�H��n�)W/e-�i�%K�M��ML`���F�ŕhۧw,�ȩ�1�
M�Tr����y��J1��	�t�p�˕���-i���ܡ�I��Ȧ0���т@��
V ���#��0�y�S��F�ͼz"n*����%ս���H.�=�����ϣ5x�Ե���[�F��9#C#cb�ei��e�S�,ǅ��C�F��ի*L��)���S�J����%u�V'צ�]���^��`�)��D@�sør��̽{-7��g����Mj�(*�C,%2�e��$k���Q��8���64��ϷAs9��m˷��F-"Tch�f��է�+m�.��A�e�\���*Δc����$7p�c�SI��� �f8��[6��ޜ�Uuh�Nm5N����gu��vV�a�@R�/]�9Yl�� �tu�q�`=����f�j�5�p���8��8���F�{n�l��P���T*�NM����&��*�ݶ�"&��x��pJ�4nܒ���ႅ���21nSp�Ѱ�n@񣖤�����6̭�	�Xdݽ��V�ʉ�)�WZ����O3ai�ڭƮZ��/_ch�Jf˽�u&,2��n���	#���D�����W5lн�k0�͔-lZ--0�I�u�kE�.�F&&�Z0�m]j�Xn����ۥ�@��,�^�+��W�d
�֒k%a�7X��tdX�;�`�qL�z���h^!x�Ah���Ѥ
�92��.�6�@̧Fm�A�X�R��wLj[�4i<��C��^a�$MlIRt��l���lS��Dc������/����yC!eeѩ��̫t�cI� &�L�Z�Y���ƃ[jhsi��Yi9�K�Y��V��[�{S$��f�ۡtV;x��(�D���ъ�3q,����j�i�!�{C�I hA��:Z O�K��� U�d��KÂ�R�M`C ��e���e��4��4.�������������on���yS6�Xay��T¨�mn6�W�fݒ��c*�A�t(Z �I�gA�2i�n�jM�l�u�MZ>-Q���K�؋v,�g((�+�H�ae����y�@����ݵ�AZ4�:"�v�6���pӁ�g1��n��.��Z��0*V-���[Z�
�ٳYy���L�nk)��٩�{�|CV�;X��o&��ف��ڴRn���U�����CYN��C&)�VI���)9t�@n1���t%
$2ʻU��ܖ�0��can�����e�n[Q<.�z�h��]��p��? K�A�a�DU�`�ɴ���eX�#t�΀�E:.f�f�5#�}uwj�Bπ�U��H�e�6Bg P"�r�f��F���p�0eYl��Q��	*6�a�+��v��k�CN+�e-��SkVXU
&Zk�Щ^��HwM|3$ݫw�����
�w���Z
���YD3� yvd%��ZT.��ӳ�Y��&���K�m��lS8p�խ,�+44#��,��/;H�B6]b+J��� ���aܦrjP�mV�w�H	��E>��7_>���_V��[�Ҥn\�鮘xjKx1�}N��ղh��\�-8'D��Y����dYY�!K��,n�u�ʺ	�S�aV*�SBT͘`2�^(��p� $Mă�Ԩ�B���ؓ�7K�k�]�JՃU���w;��`A'[���]�{8�{NmY�YY��ҸT�[#�]b�݉��-��,�7p`"r�X�c�G\�DFF��VgQ��b'ipXv6
��w��z��s(�"9��{�-�B��u�(`pev�U�Cu�;|�Lh��]����T�vw� ⹬K6�m�8|�M��G/{/Poz��vI��u�w�$�X�H�T2h�$DT)'��c���w"���������*t�����=�w��uv�.�,���x\|���y�h�N1Y�;l�Ļ"���U�}i�7���t�X��{{Sr&?��fe*���fqٱW=��7�׽(��zF?CDU�ӊQ���}�V�%.��5yw����mr�ob�}\w+Z�oF":�r[�ivs��{��W�*cƙ�IٮA���V���N�̠��%;�N�e����n�u�[��7��V�s�)ݥ%��g�2�e�hwi�qi�x(}1��Q��\n�������Ss�N#x�T�\��U0�(���v&֣/u�����}�.��f���'Z��s�;� l�R���d2n�ҫ�BR�\�9N�}�3WiҨ�O���{�:�fb�+�)��2�x�8gU�Ӭ�z2]ntMk��5��v�ԫY�^��*|V�!�֔�(�w�VV5�����kctq�-��3Rb�j�e:T|��Z�} ݂߸�q1���]�Q*ʼƊ��|���Y�U���ST�2:�W3)���R͛}ɩ}�'0V ���[C.���'w���<���w����`%��r-n��j9�[����}U��2��/{�7OEG�3��%�A;�{5���<������ģ�s�� ����J�sV<���r�&f�G�;���Q��n�nb���c����>��N2�]u;���LuJn�%W�Ԓ@)�X�b�4֕�]�k�N�M��ٱj�1sͬ���[q���ʚ-R�aQܺ�S�[���+lQ���Z�6 ��)'c�X�\��9x�>�mk�A�bԗp<.�D�8Nԛx�u�
�cSxh�KU�;[�4]o>9�� �d�`-�%���7Wݨ�h�B��e6��}�7RV�]��ï�OmG�
��L��]�袵B�[�Npvf�;�9/�,I�O5u�w�A�S"��]yh�Z�Tі�RWoQ|ԑ��`5�X�w��t��fY�uhΨ�3�hcZ�������|���@�4˱ٕ��F#j���6펼���sܺ��#��9w��EЈ�5t�B�6뢨��n;\�f��q�]�v`@r\:�c�qFW=rv�s6�gSa�R�+�C��p��]<!��$���F@�I)oi9L�7
\/V��fQُ�&�������Gs��Rf��!B��8�S6�Gq�*�9�[u�jP e%��vU��{��Z틘�t���E����V�r�2��8���N�6�(kr��Xtm�ݧ ��q���3.Su'j9y�u��7:�1s��*��vȊ9����)X��_U�]X�st�����n�]��p�i�h`�ewˆ��soi�un�
�HES�:+VX����M\	θ�[l�]qn�G���R��vor��ȚhjKyX9v���C+�e���:�y�;�և
��t����U�WN}+��;0P�F���B�W^nV�d�F�[7�����Xu�ժ�����q��ϊ�N�Yw������O/u����-]�8M��.��2i�I��ׂ�w��5�F�<�� ��Ӥv��f�{��3�h�I�f�򞍷P6�9�	��ecӪ���|RZ�����ݦ]ԩ��&`f���J�`�]uk�y�-���S��:�ĺX�W�D�z��X)k����ʗ5�#	�}�� ��OK�6��1�<�����7,�9�Om����s������Yk�m:�^>��=ݥ�V����=ڸ�&�\��1�!�㔻�ϰ̭媇�n��Z ��R@�^���܎k�B�� �%B�F7����+vS�a$�m����J[R/v�;�$�s�ޣ�n��[�-ɐ���Xs�G��l3F�.�fZ*K����֠⻝S�9��m<CW*�T�o_Eq�Bfm��r�S��_@^Ø���(u^r7�es�6ӣ���n���*�u��٢�st�]��-ճ%�Up�S���*���fز��eɎRޤf�̸�e�ۊ�q�d��\����W���s����z��;	�N�_I`���$��>7˜Ų־�0v�z����j�*WZ�ghO�7K�j1�Ӝy�G�bͽ�סlR�s$�&`Hh�Q8��IS�]����:Y-��kz��³N�ev��d��}�u`w|9��e �5ɍ��[����O�H
62Mh�L�3G|�{Rˡ}ՇY�� ��ze��|�l]e���D���&�J���vIn�9��n�36l&����I���@��)�G!Sz�_vWP����r��ݝE�w�r�	�.����iY+{6�oMU��]O0�֑{�^�4���6�R�{�����~��pI�n&:���Fe,�B�;�-�K��̃>roeAE�D�|��T��D��1p�md畓%��eJDG���*'��]��\d!L�u=����7m�z��t#k���7�G3m��6ٖVvn3���(*"�	�K�����E���ΐ�ʾ�%bK"s�R�3�KV�1��0toOU��,ݘ�ZEmu2�P����+�	=�r3Y�^ �K	ޔ��U�gxU�\&a�S��;ұ�;�Ùy���5}v)
����8��{8�%��3�ΤL.�4tܣyW3�>P��5>����n�8�ʳ�����������S9J�uEj���f��d<	�w���Th�������oY���Y
�	5;��k0�6tT�Cj��3ui�ݍ��mD�~�]����X���bk�F�*vY�Lc�yq���"�u&58TGl8�U�E�Sŉ�ܾ��WE�+�n\.�;��d�a�tG��+�����'�
�.dc���Z8dN<S���՘���HR�sF5�8d�sѴ�&���WÇ'��*�y۽��,��ԭ���{�Ƣz��1ȡAaX��`����Uϕ�1�\�lt/�9�t�;mI���VL͆�u������fPs.��_>�+��Z[z
��\�f����l�2`���Ѭ��z3��`'dQvдl����嘪������	�$Վ�g(h��O�����^�u�\��ؓsn�gnp줤����ݱ�C[������9t��k��Jr�Fð˾��`��V�MfoCfh�ܮ�0ݰ41N��>�Ɯ���I�Ff��r��Iu\�-�[Ua�O�N���.���1��$�0 l����{����5+��F�fH���~��R`n�Ow�*Ҋ�Zm�k-��B-9�"�eeX�:�X�.�u�9�;��I�_@���L���9�B�f:ckV:��ݎ�6���b>���t�ޫ���/l�
�o��wAy�����fF��c/�@��+jXe
ˋ9���'Lv��-tb��A7�{@J��#y��Y�+�s��.��9��wj������̰���}+��j<qB�!��r�oU��w�>�8�B�W���;rh��u�K�ޕ��(�W׷Mn�.��Qs
4��-{VxѬT�}|����X���H�b��])0w]�Y�WF��"�D֞�|lI�#��i�j����Zz�s��K��жb�0ɕf��޸ʘ�G���}�pl4dN�3��|jf-6�3�+�E�J��%�d��
���V�75��Vm���4^q���$�j��Ћӽϳ`�9��ܨ��Nl�N���(ڽ�8����m�k:��Һ+t�;��`,*,/V����2�MZR⳧��A�jv�ۮC�'Q[�E�N9]{�S-r��������Q<*ڑ��K��i���VL�Εl�5.]Fю��@[����S`w`W}2'��f`�ԟm�ǨW!�W�'�W���/H��#n�%��Zz!�`�J�G�C�۬���^�nL	��"��tb��@Y�W�+@��0��_oe����k+�NY��蓄qu^�ܢ��d���NP�	6i���Ð�qz-v�mc����v�I�wP�/t,���(�]�e���c�번e<�9~����q'^8uf�zٰ�ۊ����6���a�7-�<�*��U���mLZ�c<*R�(җ}̍ӺƍTP�Ov �lO�9����7�9iU��w%q��bnjɆq���'�f�'�h}��T�GW�m�J��f����[��)���R���pgJ9�+ ��'6���-��s�{xK�҅5���et��9P�Vt�-��nb䀼�w��t635�ʭ ��l�s�;���|_.TsQ:��ֱhi.*��?Z�ݓҁ���#ټ�Ţ}�
3����b��oQu�l*L%�����ʝg%b�m���9�sݱki�k~J6Dw*�TB�� ��͘�}�Q#n�0��m�:��hY�8rj�Kct�)lL�\�r'YUm�S��3D�K���2�;[Ń;Kz�%BR�rz�=ʳ+OS�-���8���"/���u^m�wox��=5�.m�U�����͎2a�,rN����`��+q��e�8�K)�Q�яYH�t�}8�"�eΑS��ɹ�G� ]G���hT����rix�XV�[ՙ���S���ٛ}j�C<�YKF��C�Cë��Żgj�`4�)H)jv�\]uuiR�^��֋�������Φz����|�E�Lu��to7�*��9 �g2�L1F���j�fr���4�u��5Y�q������٧���M�WX�Y��'$���t�f0���H�U�I-��gvڙ��f�P���2��u��;lY��N�j�1n�mQ���txS��Q>4T-N�:��h@[����.�.�T�+P�|:�Y2j�&�m�r]����xY�
=��sw� h]�uv8P�cj��{r�I��՚ICye)g�s��%VҖ�22�	{v��kR=Nk^P�td��g^[��bWc�Gy�R��Ϻ�Sm�ڝ������M�8�i�2�*S�,m�^ʝ�	�8*��(uf�y��G֛-!�F�J�x�@����_mt�Wc稬��r�#
\�:���u���PI3rՀ�gg3N�v��M��3v�;�`<���vJ����wg�;�%�stEzj���-�J�U�t[���`�ڢ�Ƨ۪u�_����t�6OeB༾k��F>.Ȯ�5����x�(wE�x.�7ZBup;j/��&��D��gN��0�f�Ό��r?>�q����L۾Н1G9nEq��\�D�'����M� �#���jj�sE*�B���sL}ʒ�Y|,�f���d���h�j��я�������Ĉ�]+dʺ�Z��G5��mƅ6֦�޻����A[�w���eXL�\��1�f��~]Y<���g�݋@�!��_��Y�9jg^&;�0�`fH��Z��	�(	6�Q��h�b�p�����#.pS+6D��X]�����m��6nQ����fgMWv*E��EР��;���P��� -ý��V��J����_dz]��1���̡�,I.�(v \�)ͼ��x�:����rң�K�
mV��z�h�H	�� ɚj�*� WV�	B�n�Γw���Q���x�ۗNl=]]����rՂYnM�5�
�^�]4�}���C6%q0�^��I̞s �����V�]�cB��ڃ5�/���T�1k��3�.Nkk�4�sν�P�b복aQw��f�wkH������#��F���.F����B��O.��y��u��㱂Q��q`j ͬ]I�Kh��s/+�A�g�e� 
M��f�ݭW;Μq �3�ĭ5�Z�
_v�vg=�y�؏i�J�[ɪ����$j���\�ed���X( �S�l��S���o�3��\���ι��pP�J�3��7����1����d��l:��m�uʛ+��5krvj΄ �1I{�Wf	�QLiI�ѕ�c�eA�\�/����J5��R.Ӎ_3Ps�����Yf�ct6�gq����j-����JmN���&��σ�s�)i!˷x�M�f;׆c�}]����K�v�G-Q&�wi�z��sX{�k31(h�ST��yj���7B��!�icCv�.�|���̴2��]���XJn�GNc�k6��ފ��}��|AȀNo`�5�m�rSb���҉ѾӸ0��a��)I�W�M�#�Vk�I�e<Z.�y�*����VsdΕh��/��G_���ݖ�;�)|N�\�A����6)���T1,�t��|g0�1GK�-�c׮��9M�R+��Q���j�zM�%Nd���u9�Yܼ���hN���E,�Q7"����W�۔�6�ȝ�Plasu8�+n���󩔭�$뛪��ٓ�份nukt�ڏ���N��%�+���nM��wNWi�Yz���D�6�����\�/M'،��@ҭ���v�yJBrj��l6!����Pƺ�����_˚��Z�m��X�[M)�H��,z��Q��F���SFfx�õ)��w`ǤqT]���D�ݨ��V������q����So��޳9΃ZIj˭�ee�b��SJif+�B�yo_vJ0��w�Z��{�lΧ4jBf��������C�VrK�������@�$��;���jk�����|��î�ǋpwrD��A�1܂�"�]��HO��n� DD��E�'l�X)�/�^B3Tg;�� ;D���h�m��8�V����N|���oܰ�J��(��z��G ��{,<	Z���_eJx��x������"}�k�&�����t̝��G>�6��κ���
�R�m�[w�&	ս�l�B����OE��fW>�(
�a�,�
�JjX��g)d+.al�ɀ�f()�Րggm����v�h�K��I���L��V���,m�e�r��ü�y%о9r�y�XEĔ�"���5�%�7��C����}g��Ab�ũ|���8�م�b$�Of���h�/��ft��,+���Qp�F��|�M,0�Y�@��Y3������9���ug��,g'�ñ��(N��Xg���$�U��J�+�`Ś� �t�^щ�-�ep �SCۧ}k*'%��l��N��ԪҮk�����6�Z��lr��(��>ˆ�A�g�Ï��\��h�����S�7|�[X��9ب 'H)��7�H�aܓ��}�gR�h y�y`�RN�3t ��(Q�syf��;��u��i�;�Ω�j�`]�i\�Q[Y��Bh�:Gʥ�mP|Uq'Ⱥd�Z@��ʃ�����7�h��«u� o =��X��Ƞg�"v��It
S)N�Y���t)��H�δ����ta˝)�L���]6Wt�,ƅv�=C/��(��'��Nwn�L+gp�at;{z�V�z����{]��ۀ3�mm�ˌ��?-�Z�z�= ��+�v"WՊ�45W[{ڌ��qh�K.�y뇤��	�oЗ�Mz�=���1%�b�m��2���. ��T�.�CaBL������S,tN��.X@m�\�՛s�W	���8Ռ�SF�J�dȲK(C�p�L/X���)j)'\tn�ٝ4e����-mѬf���r��oo�+��]��R�,hv��'D,�e�w�T�'
8*�<^�0;��Ch�(-,�}f�D�MkR�DӴ��iF��Wu�Δ�Хuv?XUqt|�/OJ����D4��u��9�ʎi����J�˞N�I�w�f��ѵ�p^���G5:�9�x@�։��T��:b�m����I�3�줱-/(���B'�a}}�.��=���:4�0�3ca9Lw^8R�-�]��*`r;����[@}w��
��6$Y 5u�;�9�n�n�H�B��7\�
�u|ᵚ�4��I���F���ڕ��I7O,t���j����V^���-H�㹥�x�+��]���n�h��e�����;gl�Y"���s.�8�)����PA+@Еٽ8���Z:s2�[}���t�<t�:��K��˸�Yg����ט���Lf_֎]n�[�9�,����R�yFBy��f��4�LğV��+C��o�B8�[y�)=T@l*,T2��e��6���J�q0;w��0��}��� ��V�B�Jm�k����W��Subu>9vVqS4�7�	�N�5�(��X��ly6a�-m�W{qA,�Y;0DJ�4RB��s:<��i�qn�=�n�*��a�UN͜����ɋ7�}���k��Q5��-b��p磵������g9tȁx�[W�|��Xkq:��GV)����b�fM4`�"邚��=c,�f����5l���R���b<����|r=��&�%4�w�$.�g��_6Ef�{b1a�Qwӵ���g��af�`�}h԰/�ѼV���\�(���E��S�)��XX������L�(��3�S}��������#c��1B��Z6,#�㔻wK�HB��u˰����V)QF�iъQ��#�B�CR��P�_m^o�����Z�p�z�ɲ.�ά�w���������M�%�*��뛿L�Xră�5]��w:�#5���*�ʛZ�,K��׳M�)i�[L��pe��V���"X,:t�a2���tU�Y�3�U�0�O�� �b/D7W��]�8f隳�$��J�[��pr�����V>g`���!H���U��(�/$��_]��Fbip7 �"ye9KˑL�zŜՈ��Q�eX	�nb�sْQ�WD	 �5�;�Ƴ�BŎ�'|n�$��թyf�Q�{*�3�̳r� �`F�v�%�Ȟ �u7��R�^p�b��F���,�s�ty��r���;�l�����߱=���6��We��v�ʜ$l�=��ɡWE�g˩6%V��Ε�݃�ocu��LS6yA�ݥw�������A� ���p0�e͋���Xo���\:Z�Z��.WKet9b7��6Y�):%��=���Y�0\N�����,*J�ٔ���3U5��0U�#YG.�re-ǣT4ڂ�E�
�����|�xK��4��n�"�����o����ԥ�閕�ޘV�g�a�gN�o��E��ܝe5�Z�5��,�FSNN�لDq�޾A�Rx̰�Qu/�g�V�	ީ��ae��_>ל��A�����-\6���3��W.��Tp-�Tͥj���^!X�we�9�(��=����3w��Mu��aunE�IVE6]q}4%�S��+Q�UV�G�x�|��(m�#ĥ#�*���1<�8&c1`/qE�*�8����淒�S��A����8x(L�KE��`B�����-�C��
;�v*��p/)�R�G,>��j��x�&�ge>v~��u�(���Au�A����$a[�0��p��E�J��	��R��7�OKC7{*
U2�f��B�qG�i7Շy�;5���Ԝ�ԧMc&�����e�fI��6��W�ޠ�Щ'w�:��ow�4o���4�;,v���m��_لm��I�{b��W	�+��&RL�A���m`T�yKuJ	n3{�GG4a+:��oc�8���t�A�������4j�
�LfCx�w9dL\��eY�p�{��r���,P�t��no"�u���.}f�=�m<��$����[ѹZ��
ҍf���ʱɓJ���[�b}w�!�yBb۾(X9A��֝��[�쾛���jtJ��gBڅ��m ]�v�
W�b��I;��-�ڑ�ۻ�E��T!�]iu]fwn	@N`��Kca�s%�՚N�{����vU�F3�B2vu����sL9U�����KZ��+Z�,
ؔݻ��%L1B���P��&���\e�5z�YP����e�x��n��y�^�S��YBg:
�r�,��B��T�, ���$;�P�\u}J��z�O�iV��ح�$�
�O�1Rٹ�e9����]^.y�}��
�m_vD�����)=ݻ}�J^�'#P�+U�k�-�`X�Ą��TdܮcGn�̵��=�o%mM����;���.�-[� -�Xis��WV��V8]7�=ՙ��Dݛ���8ٚ�Sl��6�31���iD�����L��<o�	��4um`@�.��L7[��ɸl9��(a���)�����i�쾆�x9M�ӷ��F�ot��F��m�Z�p��҂Z�	72�t.���Em�i�֯���VWgv�71}j_<�.K�yl�0��仧JU�S;A}!���wt��N,��\E��7[�*�O�NW�v��x�I�¬a��YN`���7�����5U�r��]r����l�zfv���/��i���c��Zyf<�����ߥ�(�kPr�Eq3`����Fcu��1V"��٪�*�1�7"7�p������t��̼U����>X��Wb�`)��w�h�Z��iK.�(�]���ZR'(�01W�d����U�Q�Q�:�s���7&.�#ڷE�|���TW>R�]�ч�/U�y��]z]��tʭ`o[�4e�w�f�n�
�e[�k�ll��u�΃�vX�W6x�����x�N�;7�������ړ��KQ��yӞN�A3��8�2�i��)���5z�� Z�x\(�պlkw&����G1�/U�b��֣Ξ
�o��֪� <����WzTu���ǹW�i`C+%Q�tݕ�k�a64\��A�s�T�pv�����}F$r*�&�h��B᳴�a���APݣ��A��{2�ի�%.��$�sw�t�
�,�9����G<���Y�RH�{c����>�,Rd�c �v�U�g����ՒN��6�B�W�8�`�prO��v�3Ru@.�n�(���:��yRo6ì��A��V +R��&�q����[y۷��g�cXQ��iB���t`��v���lG��U��V��
�6/�R��C4���S��ǎ)��Fd�u�:P/v%T �T��A�� �%+��)���ne9v3�����ͮ�n�׀Q�֟o:�|c,r�wn���z�T��vE�ٴJ�&�٢�>蹕|oM5j��qB�����;*5�����,[]9}Gnl���v�������)�-6{D��Sy�CuňOU��I����׬kԲ�f�)��Ґs4`�V(���Iuw��ݥ�����W�U��NV&d5w�b�L�p�S	�v�~k�S�A���b��rHo��ܹ&V
��dk���oj!���YL	]{�`;�W[��"Su�0����+��>��~���f8�K�_)z�:t�͝Zo��Ċ̌'��j�.�b�����:2���5[�(�;�9�6��\�����;a�-vd��kں%f���h6e`��e�ռ�hѥ�����,��"��Q�_4r.5V:y�&��"��U����mf�mHiv7w������Ei�	���¼�F�ђ�d�<d׶⭲e=8�Us֪Ӆ�חd���F�����%�S_Y�Kl�g+3w�j�[������%B1�ݡgz�
0�+a�}�LnN�ɓ&�k<�\(u^�T3�gl�D6�Ve
�.f�J�v%2HY��j�;�6k6
4`me:W�
�^:�(g@1�,����T�)��Ѵ0�h���S��=n  ��#��������;�M�zx6�(��#<��yj�1hIJE���\q+�v�"�U���^8L�o�e��d���m[��Lw��	�Bvc�`��O�ʗBLL]�
�R��zt�;��`���r��R�iʐh($4{�еDb��"Λ�F�*EVn�ټFqEZ��ȤPCP��ѱ�TU��>��	ω�o[ݎ��w��8��`���؜�DĤw}�T��{i�J^��^Y]�Uč�� �	�5�j �'v=�wJ�tk��T�*�V����{�@�Jk`/�o�+�m�5R�c�;�����~��GM���WKOk&+P��[f�WI�k�u��4
���Z��6/S�{��t�u�n�xgx�X����c�d��X���oL'D�<U�͝6��gk3E��Hj�Y,J�V�c�,4������>�w�z�w�tk���� ���^�VGLT�^�f)��[�CxGr-eY�]��3M�5	4�'MosB�P�w��[�і�pͼ ��mu��u��Qb�G��h�nb��Q��������*h�w�G��n���&�Gu����3�8�f�:S�t5�e��5�hE�.����:-�6�W<Y�r����]�zS:��i�
r�x�[Uy[���C5"+#�NW]^��㽡Y�����(cJR|��8��h����d	��݌�6�D�ۜ�D�0��p�f�>���z
�o#�]��w/�[�ؗzi�O��|_k���4EԷ�bY3��f;����GL�L���oim�])�ُj40�G>���a���H.[L]�J�]���L,��y �nf5\Y�m�
���Vs�߲?����+eՃ�^Ђw�͸άC��8�t�Et��49�� ��ke��S�[5���i:ur���������VD��]K��wc5cUF�Dw7J��$������\�M�fa�`Z�KiE�b���w�1���]$D(���h2��뤢� ق�v�-p��#�ʌC�lJ��a�M��t�yZ<O8��|(j��	y�H��w{��B��曹�Yz��l��i|ﺴ��}֒�V��-��} ���A+�x�ݡ�4�-m�_ś�:��NG���=�1ƕ*YS��Ա�fI|����Z��5ԩ���.�d�З��HvlRV�P�o�!�n�6�u¶G`̺5����,.#&O��֡���e�]�]A��n�M?-ؠOL�Nz�r��C���7�����E^N�̶7lN.gJm-�m$�!9�b�.v)���G(�	"����RJ�*���2ԩ��k���UkY,��xт�A|�
]���;{ɊU YYB�)G�Ϯ���FU��v<Ү<�Yי�n[hs����� !���^b��D^�U�c�#�gB�Va���֋¬ȕ-�0vM�흷�˥�z�K�K/m�c��N�gsGe���q�-�q�֡j]��rl�\�΍��O:�P[��[Hvgc3՚�2���i������WB	ڻ31
�����HR��ds������`�"s.��<�;2��нG�[_`����ىy��L"X[�̟d��<(���N�`�ˡ�L�47}z�O�+ݺ]�]�p�|k>"�*���B�ښ9��/�����R/d�5[�;s�6��CkS�k�Ȗ��`r&���d��+�ÖC/w�����/eFй�S������g��l/�V���@����)r����F�|nv�Oi���)�1�gMq�wd�� �::@�_ҋ+n�N|��A���h��I�[�ӝ8�^��w��j�����������4��d_L���=X��U�)��a�O�bN����;��i"C�4l֍��:6�N[-7kl����i����=m\�7��"����.Ɇ鬅��U|1�1v�q�Vd����e�|�[�+�V`+L;+/�.�C�^<����QޖLٮ	���\�ں]��#ٮ�K(l��̫y�-!�8���TMm\�՜�A�5�Ӯd��1�%�yYa�g�6h��v�7j�	�o��x^�3��в7V\�w���ݍH�b���c�ׂ�pQ�Z�(p�L�t"j<�(�%_Tux������]�l�M�yi��f�l��j�-�T~�Q�Α�.��E��Enm<l��;%�LQǴVV!��M�wKGc�j�� ���P��>��whG�"�3�
�_um�rm]_wF�G�P׶�2Ap��#*��qfY�fԊ�o���;�v��N.��Y�{`i4��g�7�ȳ,��:�\�œ��/k���JZ�/'h/*,������X�ZR5|��9�K�`���ם�e����|��ivVeDv���! ��H5*Ys�]tf�:/��3;E;ՈH�c�ժ	�����yqj��*�&���:���]�^��R$P��X�pEc{p�e�W�3	ݎVgs�գ~kK�)�#�XxI˩�*�ᰳ�S��¥�y+����?<�|�ņ�%e��(�F#�D���	Z*�mEX��QQ�,v��*V��S�iD�**�kZ��U�����PV(0R*�Ѷ�)kmEQF�b�*EŔPŪc��VD�L[1lb(�Z�(**���EA�ѩTB�)m������Q���,�´��1A1eT(
�0�`�����
a(+PDQV�E��YkmF�+&,�b��.,(ƥ6�EZ�PQD`��[���P-�!bV�-�Q��
��TYZ��)�"R���ڢ�V��c��eaFQ��Ѯ0V&*[j�R��p�J�)�ckl��j����J[�ء�]
��<��:�rIi�9���#���Q�L�nT/y�5k�fO7֞���WA1bUtVeM�hD/qG|�u��߫�56��T��B
�T٪v�sg�x�l�J�����l�xa)Cbj:�Z�i��VV�e�-WV%*�!P��&�3��9��3��s������^K�"�s�\rF,�]n�*Gs4�oz�8ō�������o.�y�G���Go�:<�H���)
��=.D	si�_Uh��ܖ	cr�l�Ut��nxJ��V*��:Ǳ1��)�3p2q䫞٨��]=��+M$r[��a�~<6�By~�t�����W%W�\�� (����X,Vojޛ����h%�&��ͯG8�|��^��o��2{�eK���υ�F��{��!s��6%!z�h�{ �#hvޅ����q�[(��p�S�n���<O����E��O��b��{-���R��0p��L�.Q���kLq��tsG^�����gD5+�޲�<
��N��r7K�K��.�T^ba�:��L�6�0V_��ċ2%#L�9{K,��\�9����F:�ro�5̫��G�e�ڶ��v�9{�08���;i�jL3��UkVj�&���Pn�]��Y�>���m�n��ˊs4��/y�޽��Ь}��;�~3�S�XսĦ�*X��y�~�u�7�aU�QJ2����Vߦ�H��E�Y|o��rV*'�Su�vg0�6�-��νc9�zR�/�.���.gKt����P���ӽ�{����=�ެ�ASް�䵋��d6�y-�g���~2-�V��L�d�9���]���T�S���v�Sn������B�s6.�(9=[�;�8\$��u�qS�ה_^�+�n7J�]X�ݚ��뵍��[�z���,��@��"Es<L.��Y3Ó�j��x<�(.��Y�\Yyl�'i�jƫ:�Gn�B��%�<L=��Y7Y�l���CݱG5,��=R��}p��0�6��VK�î���j��v�����:��HAV�N{ 0�]b=Cx,:���^x�6�t���r�9���_�¾����ّ�*�9�B@˄v�Y����j��o v �($p��q�\�c��s)�o�f�R�I<(��)YEeh˫��7�x�����[�`Pޣ���ps�G2�K�෫z������c1�L�k{O��2_KC��nl�c��ned��p����o=��V�F�X1���y+zl��{{-Y��wQ��qV��9yܯDc�a^_��k)[�C}��X����oM����1j� ���pDة�z�Ξ�kO#{��ݿJ���+׍��k��/R"p��=���Fx�:[�<9f�����w�z(3S����xjvZ���)^��D.�����UI���_.[kS[�v�mU�u����$�6yO��;�_����u\�&�o)���ޞz��yc=X��ګU�x.��|F	��_�iiT��J��37�ͥ�突彈;�ֵ[�t�P��q^�ו`��97=�K��"�t3i�Ļո��>V=�rV5��%���93;���E>o�lk�GEt%�u�t�}tW;�cR+5PU����ӊ���X��[�K���ѝC�4��@��� +��µ�][��ڢ�d炙�'TC=~��:� �p����6�.3���هH���i�X�����o��u�-�Z����+9�\����T�+j��7X��*��$���8^ǫM����i��}Zɢs�����crM�̳�.��!\�ˤ�r�RR�{2fV��8����{u~��۰�����+���)�5���3����h16�S�Ĝu� [��[���u�	T��ԥ�#�����)м�,ݪ��̵��<�^כ]�Ð�	,�������yj�vCK ��Y���{$]c�^6�"}�Ď�C�x5���{+�fh�fc�۹X�ݓ6�t#�͇{U��2�ӈ�@�kb�+z`�PJdzZ��^�RϾ��m8�q��E�q�^�)oQK��}�T�����ͅ�S����]]E��ޛ�[���in��C�{��E��Z�x� )e����[�m]��y������n��{���qA�\�u{S8���3|F�H���S\�N4+9���4��v�<�}}�t݃�5���f6���n��Bq��|��� r�^:�6�rv�mU�*��sV'�Ʀ
�[v)�m���!_v��%������F�;����g����U�A,�v�ް%�犭}�)�{"��|+ � \��r�%� �d�!v�(D�(9�zR�Aĺ�#u],�RV;�4��Һц�B�\^*ţ(�vz�7&!ݑk�9[A����:����bu3��#V�-Z��x��i<\(�n����zx�/��3xoZU��[ss���W���O;7ܱuCWy�9ު��z�u7n��p��K�U�zz��׊�} �5-�Eꮍ���fs������v5���dH��kl@W]
_vV�:܎�뮆�6.�s&�j�`Bs٩N�]/z��*�dO�#ƽ��fqn�2��/De�-kS�S���+��KUՉJ�J��x'\�ד6�:�D]n.wH�be,�w��T��1f2�w�T���a����*(���
^������`�+�6�Q~�g�S�xb�d���?����Tz�s�v7���f�]b$?k#z�ߊ�]ì�כ+&�z�{cjŌتo2!IJ�Vj}H<B�̽49>n�i�8�t!��J��k)5��f[[��S��ns�����d��������z,ʡb�r���ѫa^�E�Vh��"Slv�Ú�]@�����u�J�l�w݅J�ձ�3ü��#��6����7MV���h��a����rw ���H|��b�@�C��K"�9��")j�x܆rwq6�U�ս6��{{4Òн��^�/n��a��w�������k�����u��z����k�������1�Gl9�5��{1��-�˵�bU�Km�R9����˽jJ������ݱ�?O>V���~�)���?u޹_)ӇS����-_��;)I�Q8�9Öo{��͞ҷ޷~z:��/�+:��Hֳ�()�,v��S];WXΥy�we�:�ouM-
)FXl:�s+l	��K��՛�b�y�i�����SO�zǱ��_w�{��Ƽ���;X�	��6�"�wbf���i^wF���bR+5R��m�J��gW���(,��f��Zb�gjU�x�d���}XWm���UZ�\��l*��/�s'�\�6�`��4!5�\�⦵�x׶!\�q�
�]u[��ho���RrN�I���ecO���5��[�B�d]-nR}F��(o���c���f� ����Vɝ��:V֠u�2ءA�20�f)s�^w
�׮���[�&��o]MM�:
�+�:1m4��*}���M�-)��t��;4c�
�,gn�d*s��Uk�ܬ���+��JɶUq�͸w��f{Ŵ�������Ķ�bS��:�]>|�%�T+ˬ�gbf3'��R������5�_iMV�ةwv�:��x��o��J��;{UY�)�pֈ���ʔ&�J�K{��-��F;i
�i���n��*ͻ<:�}�,n���q8�$�뜹�RU�̪��(jkb���7掽��묊n�����[�g(_Q�ח*沺��c�b�^�hV���v��ed�Թ�ͼiof>����r9�X���k)ƅ�Z�����Ez5ն�T�E�~���W�7}���x��y�:��̱x+^^�r�iW��'����s��Ͻ�}���i[^��Sw��jl�iE
>�8.�_3�����yj���|�`v�oʭ#*/<���ά�(�)�g'N��Q������V���;�:����'MAzk.zj�kH4<�2������p�����=���FwY�Bu���Ph��SVw�N�5,�U��ù1�qU��K���}i+�?<V^.�[1��v���i�wc�y�'RÙM��s�k�k��پh�)�� �޼A�kX�ҡCB,�pe���P��I;����-`9�����.2-5��Mn*I�rT&�R�5Q載�'˵��	M��(e
�Knd��z���s��VjJ*.&�K���V�y^]U0�;��b��ȟRG���r+��vV)�wC��B"Z�Oh���������~}��V���]�7�V;"@���]�+�L��,�ǻ�wVA��Z*%�̓�����x�>KU���W�����t��왚MS)�G��m��C9��oZ��{i�9x����ҦV���;�|*���mU�7N������V����U�*� 2�w��Ԫuy���B~7��~)�Usk��}�l�mZ!���^H��W�T-8�1�����fOi�F�m蹾�\���o��m��k;��C��UȬj��R3�Ej�����3���*�m�<�.�f.�U�]��uYU���a�10�^���*\��S��Y4��j�ޭ���wc�Y�iSQĞ�1�s����e�����Bq����SsK��:��v�(��x�т@Uzt@�r�:�J�澾��͝���+u.�,���ޛku�t�[�&�C6��bUϫ)L�c8U���0�r5h0�s��/Z5j��{�����Pg*<��0�AĖ��YKOK����HP��g9�)���ƚ�w��<��06d�f�ɖ�^���6�f�*�3��������OVov7mWin�aj���fy���σ��9^��pНL�����������M�pF����}���䖻�t��e�U��Vƈ�t�=Ů��
��0�Н�u�zr9�|����_sv��)�%�"�"��oL�w�(����S���y�"�] ��U���c:�;"[e
�ۀ��r�;�d��=�CJ��tR��	���V�V%�]��V;"��YRM~ٗ�ɹ������Εt�R+su�!^�-�Z��ҕ#]H�J�T�L��*��kڽ��"�_K״��U����ץ ���}�)`i����]���zv���h$�T����~b ��G{Q�ޭ�j�+�����c�/���^�#��*��\���9-��U6f.a�8"rƻ��VWtWG�ˢe�uї��M�L]�����L�ɹY6ʟWŖ��S��i���`\n�����i�;�Ch�!s=�7��⎮�>���K�֮K<����q��h�ܶ7����W�!��Ӳ��G�7�B�g,���R��/���F� e\C�k;��cۭ��Ѵ���Xq��P�^\�I�(b�ڜY��꾿��ﾚ��ݕV��0b��j�h���İ�ך�G*^�̭}K\C��T�bUȬ��_m1��k7�T�4'�MgN��۪Y��D`��i�~�1P*�b��d���hVr�st���=�"&\2c��k7����M�S�i5ֳi3ׅ�lN�3׉��R)FVIě68�77�ܷ�����`*��ݸף�ҕ���䊍�q���X�����S��Yx����a����2�כ����ls�)1��š�]лwc6���Fc��S.�)6vb��*S�S��D�*E��Fe�����&��x�^*��s���r;�]��Ji���G��yCT�+�	�2��Y�T�^¯I։�X�E�8�}��]ۑ��P ͭzo�s�>�/���\&��fn�|�n�� �Y{�V����/��ԧqj��m\��Ȉ�o���f�\�^6</gCR�{-Gـ��v�L����;�ҧe��|-���>��������ZS���kCe�+5�ӝ��٤�@ ���=ʝ���Yg���GC㙜�b%�,l�:�4�6���Gy>{c��&Oέ�dV���.	W���*s~��ݷ��Y@��#�v����8�2���\����wv��V�	h�h�K���릳x�We.�g�N��+v��3z���{����	]t��vj���=������NFR��]����ݴ���-\�[t�ŵ���(5إ���t;�Z����e���/�:����ߝdVg�A����e]ir��U�>�T��76�h�X��3�IJ�]6����8�'SWrsaՠ�X�S3 �V �Y�����,{��.�����d8�fB��P��� o��nG`
��lѠ�S���5����V����j�!TՉ�
�ر�38����]{I1�3�'qި��S�@P[ky�	c)M����0g';�.*s�o���&����0�Ӻ�uk���Љ2�\Q���"��ڵ�w�
�: tRޮ=�r������e0�f�2,��:k{0�}�.��Ձ��;Ќ����9�Ova�6(��t�8�Vk��3��9*+Gf�<��}Ɲ�6�
:C���O6�`pz��Q.�v�<�0��1܏Rbwv��*Y|��;�����Bie;�g)E�V���w$��ݩd��W]�'�9���6�b	���oT���n��+is�u9�/9�N�7�Z�v��Ud������2G�jAa�uv�Z߻��j�8:�.�xp��!���bf�R�[1��e�;���tn�s�Ѩ��ƥ�b�3����;�lFN)u`���I�huLy$�L�A(5|���;�~�mMu�xL�XI�SRN�hΩ�;�w:k�bQ�Y��ei��]�{�������j(���T�Y$��Ha�|������1��+z��213�68�/RR渁
l�W�4[ٕ�Ѕ������F��N�Uۃ�QṀ�T9p���;b̀�v��%���rƥ��@־�E!%Ϋ�޲�:S��2�����}����@����z���S����81k�N��"^V�׮��l�bT�JrR�:f�����K����(��l�Җ�ER���]<K,�Vk,Ӽ�F����
MS� r[.���SD�]*��f'Wc Ρ�2��h|�l+���Z����;fP�L��FF��2���*���B�$R�U�m�V%���Z5K(�
���*[A�+J�(%��Z���D�R���-��V�Z�mmAU�aP�5���+E��ڔ�*���Z�A���8�F�ֶ�-Rѕ�j�\\8
�\a�-�T("ՌQT��(ѕB��V#ZѭeT���pR�����Q�(�6�YH�R�Q�ʒ����ZƖ�m��\[�&��1��*1DF�A�j[QJYUTX����EFb��ѭV!h�h��[ZְP[Z����X�QQ
P����(�TU�
��jQ���-��[8�*R�QF5*ԥ��R�lbVŪ�kF�ȣl��%m�����DkZժZԣU�+P�kZ��m�֢"�QE,�Q�KVKBԢ�Tj�+��a��,�\c[*DQ�,��+T���X�J��ŢV���#kR�F"���E�YFԵE��1j�)k-���>��\ɪ����v'���=;V��d�~`��ڟq�d��QV*��S�7�([խq�{b�_;<	��Ɲu9X�B,���/9ȧ��<��b:��gwWbe1����~+0�rM�ds�Uӳ�\�F%"�U*{����1�Vdrҋ�(GWv�sGm��]*���]����f�:�t��PeT�ާ�qvB��#k��������mi
����k���U�ٞ��Y}ܹ������}TĮ�B��ݑ"�<k�+��g,���e��)ד��f6��e98�O�{T�7�C��D��x�}u
�}�x1i�?e��,�;�=��|�Z�k���A���:�`�%�Y�/�t�'��6���~��y�1�1z�zc�H�cݴ���#���
�5%�������i�	�Or��Ѵܕy��Iмʡi�j+[��6Ga����&{��2y���͙�]z���s�[�u?��?Q�/�o���;D�g&�6l�!�Lo+^w���S�.��y�&���V%X�M����:��7�t/m��F�;� ���}J��Vxq�s{x#�ƒ��^k�_*�R˰K��#)�qS�o�Zn۸�g:�Mwp�Q��5^��u5�ۻܢv�^�ͮi�ڞ��Ԛy�>ս[�^��x�[�9:7�<=���G�9�����mT-�k[��ʆ�߯�`��+&um�ZՆw�٨�1��n�+5�sk[�z���j�+��F�<�J	V6q(�]Tf�c�`}څ�#��s�U��>y�;{����	��N�e�u0��IY���wb�g�3>�Hд�s�9ov �WH�l��j�6��8�)F���>�2����\f�Yx��⠓��2��H]e�qW�]ur�e�ah�X�2�S���B�fM�o���P���&%[Wp{]�wm�S�U��SJ��>Wz�*�dH�$xP-��
�W"���{7�:]&g1�nDuicW�������UՁ)��xvD�g�zev�Zf»�۽��*%�o+y�`..q���+��nR�ld����螮g����~�G��J�-��+��{|�΢q^�S��܆��j���J���$WQ	ٺD��&Cc2h�ՅTP��,웈��N�$�
�i�<�ޕƕ�^��,3�-C:�v��T�_V�0��\��m��ѐm�#�X�*��i  7(��J�j�r*%,ԧ�g���q�>a:��xj��I:�P�J�����`z��>@�CL>�n�����=AfNs8�̙�3�IĞLv3�lL��fG�W=��ݟ�������2m�F|�8���>&��C�S�T2��q����O��a q��a6ox4����`��OX�v)�>_M^N8����Y�w}��xA��|}�2�>I��y%ՒsN�"ɷH�'P8����<�`|����'dՇ�z�Bd��C�a�C�l�
I(��.%�h�=�5-���>��	:wI8��V�!Xz��~׆RO3�{��$뫼I��o1���}Myd8��2��P�I�P��H�Ý�q��Xn���s߇�D|>S������M���14���%a�� |��&N�^m�x�ϵ�.�'��y�)=~`d���m�&He����o�5��T�}ww7�w��$Q̏"Ha'�/MRM!�r�O&��}�Ĝed2k��I�O��{���6�=��	���	�	'��{��`y��]}q`�~���L00�@��L$6�e:g�Y6�ɝP=C��b�{a6Ì<7N'��L���u��XM�:����X��|�}��O�r���%�t"��b'o�Z쏇��'�vo��Ci��K�M$8���k����}C��A@���'R��O�u�ɴ�I�/�8��l&��{�=şy�a�˘ˈ���V��b�����'�a���OX�5�8�B|���$P�2�l���q�A冐RL}�q'YXՆ�q��S&��:�hg���|>�_�w����cf�2w9g|8��'C�Ԟ�d�l�`z�Y��^�C'1�!���4}��I�k�c�I�>MXi<d�s�$�+̏G�>�:}	]�3m��h5ّ1O+v�����3?70}��|�2�
�-�;�}�=R�q��ǟE��]b-��8�F4=�eF}��+�0�nS~ɛ=���j7;�ղU�kkPT���v��s��t#�>&����0 ����[�b*<�[�{O9i/K��� �p:oxϟ}���P6�N����������G����]�h��"���'{�u���3��0���0C�q�i��#�g�O�T ���y�ǵN�}���6y�;��������v��'Y6�Oi�u���'9�:���&S�� m&�5>��=ClϽגT'�{��VN ��� �N2|�F��q�8�8���k]��d�0���ē��Xu����8ɴ�~a�X`u7O_�N2s�|É�&Sg����4�S���Y'ϽגT'�u����z�}�=��^{����XT����9�8���&���fP�Y'S�2kVAg:�/�8b��H}�Ρ:��9��M!2�<�q��w�辏�����f��=η�1��Y'�t���J�$���ԕ&�Y2y�$�M�z�����T:��<�������q��^��He��O�@��ٮ�ʯ��������Ԩxɔvw�	�6ɐ�3�RN��y�$�RO;�u%d߶����d�ˠ��q��T2��q�uC��>��ϼ4�$I��Q��[$T�_'�ǹ�����Hq?Zx���`��OPY������N�8<d�a�גT�'r;ċ&�`g�:ɴ��'�P<π�,�GO����n~�^j�����u�7�a4�w��C�a�C��q�T�7��u��s�:��T;�B��'{�0�2l;�|���N��$'��b\� D{�V�����ߴK:�w���������'�2j��=L�5�I�*�i�IS}��N%Bg���N����4������� o$zQM������7~W'�e{���}�L>�;{�,0��4yHq!��z��I�OP�.��I�C��:�$�<5�2q*:�&�u��=�q�M�{���s�l�������u��ky��wBN3
q�K�V���=��9��(fک �:��A�i��U�Nf�mC��H�"<�ф.�ޛ����L�)���݅B�h�Sb�}S����E�U��i<���E�m�&�2�� r_2������B�s��Ο�����d�z���I��B�L��|�f���L���,����d��hM��}�}�Y�P>>��A��[���h��ʗf��]��O�G޷���8��G���=��gw�	�'����E�ɶg1��C�>fG�4��0y���Ad�Փ�I�Tϴ&�q��;=�Wx��ꚪ|7�y�DQ������#���7�d�'>�w6N�z��|μ$�����a	�w�a��<�&�M�S'(i�cϰd�V��\h���M}p�;jpMn$��a�<�������#�_�N0�x�I��G�1�=vɩ��N�>a��3�N$>��|3OP���E:�Y6��<d�C�����FMGe����q�����=�? 3'R�<�'�6��hk�!�N0�4��I��x�I�^�����&���,��m3���N�9|�q�d�������!���"_ص:߼�0��G�O������'�Y6�!�P�&�;�{d8��L�_�N2s�u'��M��a��&���C�6�c��Ǵw�ܝF�6�+�u��c�@$}�S�@�O�Xgx�0�O����q'����'P�&ܲ�d�'ڡ�i u�__�N2}���3�L�o]���w���k���w�a��'M��)&��\τ�(O3�M�Y>J�{@�N$��`��I���$�=3a�N��-:��M?!R`e�|��㽾wvl���y�q }�8���:�C,�1�x$���Bg��
ɴ��� q&�=�5��'��jI�{�����y���F�Ϭ��g2c>�߷�`z��wN�C����{��8�2u���2w`�;{�$�RO;�u�d�VL�<ĝd�'�S^XN2z͗��79�ta�2� 穬3f�7�V���w���T���z�$�X�5z�i�+�oC�d[
�[X�E��Z)���WQ�Z���[é�vj�s���ٕ�k�b��rY���_76�����AM�uy����7ь}x�%q"3��j;��ZUM��_��?A�=� |�I^��X��u�̝d4��n�e'R7�AC�� �=�$:��1��2�u&�5�+	�7x"ɷHs�S�_k��#w��~�>�{�!>@�;�2��u�Xz���!��ԇ�0�a�=�q$�7�&Rq!���
d�+�!Rz�ýד)'Q����놫�=�^}���f�ݟ��4D�]��9@���L�L!8��w6e�	����Y�C3W��S�0�?S�,������b���`4���q|�O��-WLџ����g|< �i�����d�2f}�|����uy��~`f� �6�O���C���)�x�m'�T:���'t{�OP����� K�O�Q��u�W'tꢞo>��>��Y���u��9�L��|wz�d�2g�{�>p�x��1"���K������k�C������e'P4�i��2hU���7���]�[��C����I�35��6����pq���~I���O�;���OP>;�|&�$�&N{�6�03{����>L&
������l9����3��(��
�4�6�����N����x�i}N�u���~�:���=�u��O�μ$����אۆ�h�ؐ��� ��;�Wy�n���j:���}ǟ��L�ha�<�����:��(�&�q��Y��i:��vs�$�t�']0��@�O�$�wX��#�]\��}�Sk(��ny��2f��ϼ�����a���ݒ��<d�7�a$���P�	��6d�V���2q+35d8��<ݝ��8�7x8���g����(�:w�s~�����eLSo����>��ה���������C�m���)��l=N��4�M�Ň6����2u���h��q��<3O���I���;�<��.$U` �x����Z?�_�TiHƵ��S�T<o�ۙkP6&i��~n�Ԗ�����j�ǻ�٥'d3B@�Yr�x ����1P���0se�����O����_r;�R��u�X�. �X�r�RN�V�X�;�ޢ�yV��Jp's�%q���^��ٺ���s� m����wR��f{�x��{�N�Rq&��8��Q�m&�y��x�m3�dۤ�KC�Iӄ�e������;[ճK+�}�x>��nߒN�ߖ|��&^����,��wYS�f{�y%ABy3�N!Y6�&e� �2|��d�I��6���ϝ/�bD]����u?k�X}�<G��ChI��5�������Ng�8�a2�<� u�L�;�|$�=��<�y����Jɐ� ς>���;��#{�?]i?_Go,$�&S�l=�I�y3C�+�!��ΰ:���5��0� ӨN�<�0|���Ag���N��K�0
I���^�����O���Ѻ�>�}�{ĕ�䬗��|ɧ)�l�N�X{i&��4:���<=���u�:����<Bq���0��,�s�	�>�:�n�E��v��
�_sY���z�t�k�VV�oIY8�����ui>|Myd8��<5C/�'�XW�O�x��3x{@�!��xox4�2#�i���.bz�Q����u��Ha��,���!Xz�����IĚ�ג]Y't�,�t����u�=~O|�`|�L����35a��P���x|@�� 7�����Е;�t��[|�5/���
IS��p|���{�M$�'�Xh;��>d�k�)'����I}�N�.�E&�����i�4Y|U��> y�꿳]�19�a5������a�$���OP����u$����ԝed3�bi'Y>J�]� ���L�޼�$�k]RO��`�O_����m�%��}5�>�|3�9�׽�xC)YӔ�e	�L��z��6���$�a��:�2M3:��8��g\��N�|��}�z��M���q�>[C���QN�2)�������z�T65--]Y>��gSE��]���Fta��y�DT���~T!z���z���&K5 T0�-�o;z��,�M���vK'�n��G+�["��@n@k���G��I�
ڻ�nlऎ������Nb�&��B�{����yqTev�Y߽�|$�����#��>fG��'��,�Ad���:��.}��a�N&&Y�sx�d���S��d��N���=i�3�sܥ�V�N��u7�ܹG���>��FH�4o�H���A�Hq��������}��'P2j�i8�ԩ�{a6ì<7N'�'f������k/�6d�\v
�/��w;߷�/��z��8}�bN0>I��y�Bi����!���5�}�6̤�5�1�$�&���
I�>�8���0�N2q*e��'X_s�z��xW��������O��>B�����S�a@�O]�jw�����;�p��c>C��'�}�C�x��l��q�2�d�}1aěe`kܾ��QUWK诤����{��͟|>�x2 �Lӯ�'Y;�u&�0������]�h��"���'{�u��s��d��C�q���.N0��k���]1��N������|������~Ň;�!�hq���t���8��<�=~a8ɓ��ԟ;Be;�hq2��i������^IPP�w�:�d�>�\a��g*�윸��ϵ}���z��Q�q�Y�4:�$�L�������8ɴ�~a�Cɺz��q�<��q:��h��f�w����dr�aM<S�s���W9����Ҡ�:{�aRm�&Ls u'>M`��d�2���8����O}�-�@�M?0ы�!�[:������#�&J<c��f�c/5���z�R]y�Y&���5�*I���ԕ&�Y3瘓�6���,'=M!ְ�a�I_Y=��Xz��@�xY���k�-���]���'�mr?!=@���T2��s�'P��x�|�I��ϒT�'��:��o�F3�u�l�9u����e������zx(ߠD�?W�u���o��wws�����j����/RٷI'�>^�g�j_e�L{6866�u)a�!����aU���4���8�Џ7']��C��bϛ���QL�V��{�t-�:�.�e=|c�o/�H;��8ft�7DL���&�
��Q����݌-jy�m��&~�:��9�0e��,�� ��O�Y��
M2{�^d�a��y%J�w.�"ɽX��d�K+~f����Wl�Q��[��M]��y�W�����S��Oo��0��Ө,��!��u��,�aԟ2����
��N�8<a<d�y�W�I�;ċ'ڰ1�x��0��1�������o`�e'�����z��y�z�!6�&�z���\��B���$��pm��P��14��>eC]�T��z��#ޢ ��\��LPY��^�]��=�:J��x����I�K�A`z�O��C������i3���e��.�i'�u���L���8�Ă�c�a����=T
�na�WY?I�9ֽ�~��=d�����$� d���O�0�&y�H������M2��a��RHi2���N �e�Hu��.�hM��@�(��Q����#�����[Va�Ϻ���]8��T'Ns�:ɿ�=9�@���:;�|$����^nO3��E�ɶy�M2��0��P�$ǟ`:��L���$�*xo��[�q�v��J{�M����=�y��0�>G��m���&�{���d��N���Rz����L��O��ԋ����&�M�S�e�g{���u3�;s�?g��s����5��Ԭ$�'m�:j��N���8��q�n�8���&�ޘ�Ԟ�d���N�>a����N$9|�q�Bi�ȧP����{�1w{}�.f6��g;{��Ͻ�@�$�Y�#�G�d�V��6�������d�=p>:��^1�u��;�M�Ċӏn7��5�Z���K�~��oå��V1)��ʞ��9(�Η��d���cMBOw$�[&����V�)�+8��ݰEJDB;X�Ez{EٝF�����˕Ha���Tw�-Ô:�lt[�k��.�Se�	��7X����/{F�n��%���.�.]�xt��$z��X���F���J{�{��tlD��7(J�.�'�2�p�w\V����}]����XEe���#4�wy�_UGj��Sn��\t�4��(��O=n��e�8�6��[�Ža��Ǽ���t��M�ñ�vD�g���Y�Y6�췉71�6�I͊���$���n�]�S�o�9��d�g�����]��c� �2-�;��S���ٵ��kͯtR�A�m�êaQ,��U���J4p��������{f����0\���~r���Zد�f�)]�����<bF���\�w�p�Y�7���au�@��z�l�����"�9w554_���{-Y����^_�����u=o��^��e;C�ù�\���1�4-[�m���饹�4����*�Ք�޻����d%:&Z����h���W�A����DO,����>��W��)l#��!~_�2ﺖb�sd�5ܺf1���r �s:WNx�����Z�^^c���g2����v�Xk*]ɮM�XIw�\���k��E��7rN[��s�����{6������U��sY3f$3/��{�g7;�x�-�t�'2�j�χMvA�yvkbU�f�B�emN�v3z�jQi�9w��Ӷ�f�����j-�ʋ����3w��u+�އT���
��vVj�i0�U�]R��G&Xq�25��'o^o>{�Ro����|`�/T��m�ʳ*����w-���uj�g�k'U�Qѕ���ؔ"w���r�89<��m���n�����y���� ��N����{&��#b�*��=�q��uj9;	 ��v;�"�ή�&(o_ �`̽=X�Q�C�+�(�WQtټ"	��o���vX/Wa<�*��,�>��^��U+y��뽁Ð²���E�|I.�u�1�=�{x�'ع��=\n����}��;И�=��;�f�K�Y��Xⴷ:|I��u�z^ou,�n��աT�i5��n����q��+:��n%�κ� �󷘍��Ϊ,Q`=q*�^�n��"��N�<��/2�')P\�Fu��%,>��p�.ڧDт����jVX�������r�[����ξ2�g�6��8�)RG
{@�Ӆ�1P�$՝y��k�3��{���E�]��������X1Z�TUEh�q�n�(�;��?���r4[���3@x�����)��ܧm��+z�~��4�+w׉�W���fj����Uˋ1�O+o�%�H}K��b�V�μE��#z������<�F�b(�Yi�m$4h=��Ӷۼ�j�sC�I�:f�Ɗ�|���=�wxD��J����q�r�����=\�Gi���gr���eR]�H���52o5��SH�}k5���]��]�;Hgn�`�5��G=��Wu	� �V ״�_q{��	ueSs=f�r[�h�I�.n=�A.�o�;�mt�&8u<X��B�ҫ­tyz.��`��4��wհ'�VW��h��:����:��z9w��YA��2	m��|�@�*���E1�z�ݰ�^��kV�61������WXy[-��-���8��@����f�Ϧ�:-:m;����M����`��.�Aq�S����:oa�+�2nQ�q�݇:R����,>�=��'s��U�CqgV+�]��ۨ���x�Z�1N;ۍ�n�$ ��.9o�0��f���H��a:k�R����>*�!��|va������ &��R�{_ľ�� N��v-����%[
�n��e�|�u�T��&!/nXPX����t��o�N���Et���>�k���\��f5���5�X�H���AJ�]��u٫�w)ST錂�s-� J��u�g2�h�l8���,��S5���Իv(��=w��
�t�Au�x��]ka#M+I�
X�+)Q�kU-0���D��U�ZťV�*6�ZQ��kU����-�m�+Am���b�m�(�6�$UjUb��jѕmKkh�-�+Z�IA��J�Yamm�eDKkl-Kjئ-1Z[��,IiZ�X�,Q�J�	J0QaZ�PZ���e-�k(4d�j��	Q��V�ij[Kj�V��(��U�جcU"Ųը��5��K�J�6��"���j�D[mkR�F���YUkQT�m�ʰ[JZږ�֍KPYlYX���EPmmj�-�[e�Z�-������mejV�JQ�J*�,F҅�µ�[[�4lbT���[��ƭ��F�m2���KF���p��YZ����U-��VT���b�\`�-��PeJ ��a����Q(�,��+U(�Q����Z5*"��ڬm��`�\`�&)J��cQ�+kVcqcae�U�m�[+��Kee�,�Z����K[n��"��@ @@U d�ϕ���Z9�+�,!f]*�,SQ��ґ\/0I�h�p�p��)��kp���G���f�YJ��b����� ��AW&_<�?�f�
t�Mdqu�he�v���;��.*⋳�n];.}t�hP���2����ކ�)�NT�2t���-�X�DH��Ҟ��kT�Λ,���i�����]�8�y��1�n/N x������XP�7��%��F�j93,��ZȻ0�tGE�z��	�Wvu�*�8k��)�u�K�o��q��e.{^�,��m2��=��ġUrՌ���.�-�Jj/K�!(�byB�s�uF��xA�ȭ%ÈP�="�SնMaO3dv����Og���;�ڼL��=6������buE�ʀk�ۨPl�elEG�2���Q�`���]��KW��MD"�g�.�޶]G;�<)�닯z��L��Bw�K�d���p2b��ݏ��,;8���%O�v#�͘(��tB:�X9�rȡ��uU����;ޭ����`OK���E��x1B��h�|k���Lpf�|B��V�Ǝvvf���ݻ�����`�`�v�>�t����pw1�^+'+	Z��H�T�c5���ˤ.�k& ނ�MfL��|�V����zu�ھ�!L�b1q5�����3�)z�U?{_�����+���wi�S��]�Y/JY��uOV���:���|ހj�FL����8f����S�_��i�Ã���������nU:;\-�}x�X��m*�����n�����7�R�9�G�mϬ�������x�&w���k{�="w]�mE�v�8s�r1+��X���C�ro��ߤ�`�խ�uuosS�5+nP:p��P�||��^����;g�CzR�"w8����o'�;˷��e�ʗ��쵁��Uj�x�N}1�W��0�w��z�=���*c�q�~�FSۿon�X�oR�Lt61F�-�pu����E�uG-�`_��k�3 ���|�S��7v3}:r�6��ӿ\0c��%OB���ȠD	�Hҋ�H�
]C-��n�>�2��b缤a`rT��guy�M��,vF��=aT�D_���Q�~5���[�Xϻoֺ}M��!��\Jr�1���T�(a�S7�9�rw9�6�DB9��H�fD�Kt1y�8U�=mapr�|m�J�◻+���,bx��N��ٰ���c�e��D����]���������JJ�u��"��l+�|��#�N1׎��}Wd��b��]�>�A��s���C����rz6b��Go%=Lt <��kWv!r]�wBRќ���X/[R��K���� ����-Z�3;�uq�v������u�2+�˜�)+��}����\� sj�Vr���ت���S=�)��� ���y"��vswJ�4�Q��D��r��g��B����.�64�x/:Wi�I)����!���T5�P ��F�"��Q��g(\��h_N�[�^עQ��e�W��et�c���Žu�%ON��u00J� �k:����n�˾��ND�"q�� �Pr�g>ȹ��MY��`�����c���.�lB�PhVٟ&�7"C��̕�kM�>G�|k'�Vg%;1���C������ES��%����F�!�d�A�
��x휺���-��F�X�w�[���c�'3e{:@��(ܕ�-s��}�L)wY;u�=�T���>�{���N�4_������U���	W���|��g0boiE5t��51���m�r��b�u�O(����Cf�Zchz�Z����,�9�{VP͝.�:'g7poe�+�4b����z*�9�%7"�0�=~������Xn��؈�3f%`�Hc�(�(��U<=9*��]���/�4�Т(,T���ӻ���5�,U�c�Uy+N�5oUu�QV�p׃��.����t�"��gsf�ǆ��������G��~��*B��K����n�NR��=;E����9������3+�p୭42�-R����|�'02���P��V�N����Lk�5�ySK��/�u��~W�_}�	Bi�NU�(�}�9�#q���8E�����ګ�6�;�����6�)�r��U�gmf�Z�A�Z���D���6t�1�#�Q[R�7�ĳ�1�:v�G\ܛ�l�v�T���\˾�<��y�S\{e�娃^�!daEp���+��+�<�)��}*^����c:9�w��݄`�U�^'hMK���+�(s�*"�1�#/%B�j�,l�U����{Q��n����b=3�b�K���h6^%*S�N����h�G�e�P�I��✹ukj�2�4��֍˞Qe�x�n�V���E�VأJ���hU���|�\��J#�4�������I��p��gB���x)Sqb׮�	C�>�:LM�f
�w����1H�����6��Y��)�sCa��9.Fu�T�%!\1.C����3p�[��{c�N�Ef^R����̅/�,ᓅ�8��%��XQv��'$��n^ŉwvFN��+�k�ڸ[��b����}�\tc��R�����c����1"4҂h�(�������{w˴�%�+w :U�nd��`����eq�@�k���s}���c$qU݋�Ffw"]��<�-�Bf�������tht�W+��×ҧq�efh��>��
]M����W���-���ۚ�)E�z�
ֱt7B��5�d�����wv�`��[Έ5��ʱ�zٳ]]G��0�^[~#5����8{
b�gZQ{y6VDߚkw=�[,���ZUO��أ~kN�xT��.	W�4�ʽ�F�@ʄ�\fyiP�U$gQdB<��Χ��.�
^>&_���`�4��&�[�rj�Tw���;&*��B�-ܨa���IӇӧ�g*�xF��-Ek�`d��)gv8,���qq���&���Qٜ곗D�d���Dsg9���/�,ϫ���,��Ur����y�d7���7Բ�TR��悢�c������)(���k��&�7�����Ҟ��j�9��oӊ��	���3K�<F�k��B�QXtGTu�SAl̓�@�."�)e��)�q��D�͛���Fs�����;���Ns�y禮*)E w�2��r�vT�u����_/a��%�����ޗy\�e��e��Q~�'�.rN1��u��"���Ǿ�.4������Hi֝����(x	�O�״/z��}\EXn��������C+ -̀P璪iˋ��Q�6��M]�,6���u�o}fQw;(#SQk���1�oGv���ef �^�����g��I�^щ�����
�˶�	�r�>�Df��}��p�;�܅�u� ��}�z���.|��5i�d����ugsIT��1IK�_�� z���9^:n�Q�B���Q���0���l��M��#�,�PZ�
X�ν��^�Q���=�a>����%��r	u�
/6na�.��GU�)�#�)d���;wVf�Vr�~W������3�z���^ȜS��sh��m5Jl��E�T�Q���}�X٨,9v���f�
ɠ���v��r�����?	�^")NVKg��:��`�j�z)��=�U��y�s#<XC��!zCmO5�٩n�Q�gr{w�C�;�ܩ���}1	�郡E�v-����}�tY�,�=&�l$�l�Q6Ō^��R̎n�V�s��ݹ`��7X�+U��	N8����;g�����%��F�@��q��'T��^��E��:X�xYS�Ps$]z��0/;�	�(������}�`���_-���}��XD��óuH���@�͖�߆�.��9mP{�Ŏܭ��軵Ϲ¾�R�ɗ'yw>�`�f�`�[�����u\�3���_��6���U+s���`;%n���
-m^�,})y,����/Ut�q�!Q�����H����Q�QL�fnwrΘ��juz/��E�jt0��M��u�)��ú��M�c�X�8�s�"ݦ��Pu9�t:�m�ڙ�g6E�W:��]����}�4��'��,��0�R�9<�{��`�`'�,vF��=j��"�؟j����ܚfjԡ4�[����<�h'�́	���b}�`7l��o�mܝ�tͨ�3�^5��F����^�g�e3އ��(�oi�8��q�;=J����o)臩KE�>�a�\�+2�S��9����v\�q�B�y8EO�6µt�M�+�����WXqm��^-�����VX�:���oՕ���r���hB���(���ׂ�O�<A��d�Rx�X�����aUԯb�A����K���H�r�ʈf��tϏ��'�W	�-�G�W"-!���;�z�Zt�Yjzx����x�D���Tt#��>�O
W�=����9������Nlh�Oy]v�X��0��j��w�ݒ�³Pk��bjY��P���c����X�Ɖh�Φ�֊~R��r6fhk�m���R\p����K7*"��E��T=մ�E���:m��5��+ҭfyT�-I<�*+�ׁ��Í��51�^o.�DFєS/q֓@�x59���f��ᒅ��yԟs��a�٭B�i=�]:��T����V�������� ��#]/�,�F���x���ْ��/���|x>ʺ�f^�o
6����p���C������VE:q�Y�2�`��������b��X��.�%g�
��YL�y�Vlb�1CU��#WOH�����:υ�;���![[�̆4�@��C��#dd����(la}Ή��K��tKʭ������z򆰫����>U�}���m���7I�O����*�z��wr��mi��\��E�gO(��,�B��<T��WZwa��<�(�V��7�s�zgX�F���C��:.�>g$`,(�
.}�'�R6k���,� ����Uw��u'^����3�N<ta�7�.��yD�l�M\qH�q�+`*�=�ĳ�08gN�WA�n�4��z��s��F�mrcy�]e���{��c!V�³oH�!��3��2�]詘�䕡b����`�bٖ� qrt������Wgߥ�1x :%��<�҃��$����Ń�M�w�k̀C,���Q�"Bں�n\���ُ��0�
p�=��]GV�O{���תټ�\�2%td�]0I�YEm���*��R�͖jE��c��Y^XV��J]�b��V6�Y��=��&�\}�s��o�i��h��_��7�%ջl�Wf�͒�u�ץ�7��Rʻ��E�[9٩*&��j����Y#�g`֕Z���֩9^κ��W�PC:�Z����ܢ��=�hUKK�9�B�s�%�4;d2�e\^��7aؔx�0M'1�5H��G��5��q��A�+u�i�ᠮl�{Ӓ�gY�f�R�)�}hK%��D�N�y�/\�h3�7w��F����o�ōu�*v�e�s��`�'$��ܽ�b�2]��յ�g]!oǲ�!����\q�>o�(]��v|/�"���
�n��ڊ{o�Gwݽ�� z���y��,eF@xBVD1�mS8h]�F��D����au%���Z��"�B���;&ʸ{��<���kN�aA���ז��[�d��pB��s�|>�fDd ܌آ��7��E�YL�5PX�jЃ켈?r�x�y�����q�`0��-N�?v]�o#HC S��X�ED,R��p�ή6_F��hNE��s�̏����y�s�#��?OlK�F}Ji���,�^�⫔�����:S���<uǒ�`��D�+s��+���� cX��-�}��qWM]U��Dz��%�)5��8;W��Lggn6���\�&��Ӛ�B�EHu�-�q��8-�q�N'r�Y��q��K�b|�$fMY֬rX�mh"�4���U�}n�B%���(�˼�ݕwVh���kJ�ke^��\y��[�%9ҍ/�!���59Vw�������.-���gWd��wo���6��GLoyT�[3`�!b�\^S/�D9+�zU��S;v�Cw��z��	z�9�<�M\TR�@�¶}�v�u�s�Y�ǲOw�g��>��6��*�t�7�,�r9F��{�����]���ZK��Bز�0�1�!�������8��� ���w��5�ަl}\E[u�d`�'T^����/O<o^�����i�`U�׵�P5䒏^�Z�޶l;�y6pS���

F:s�����*�G�\�Գc`�J����S�w="Y� � T�F�0Q�CB�r�lJ�+g�Cq�m��ם8C�(.WQ4�k��'��%�߆Y�xeCBʾV��xL�󰍱0��]3�Ǘ��Զ�v�m���HGaL��TL���dA}N��h��sb�t�h�V"�6�Lʔva��(�!/`�j��6h�p��g��M�R�ޝ�g�N��EN^._t�V��|���n;nqG�#q�#��q���t#��r1+��X��8���g�]�S�r��׳�P�]Xn��W���	";I�c��b] �5e<k'J��`�0`��fEo��<����8�E��eo!N�̍fj5l��!:틧Q�Dk�]�d� yVx,G�u����L�$9�u05� ���:��/f�����Q���������٥�{w��K���Ѱ�,T���*k�W�:ٵ`��7/8�wG_n��g3�60�l�vB�wo1҂Z2y�ɝՊ�i�K�)rC��֙Qv�`�)���;�Ѥ��:�����P"h�\v�����k�5��#GS�w�0ݛ��[up��@��Y�e��������V=W�K63C.�v�Q�v� ��whSG��.w7[�³�2���S�YOV
�2�&�h.�XoN�����d�glSV�v�n��j�.��.Kx�a�̦�� tKmE2�I%�Ys*_�>W%)��J`ۮ�F��8�C2�$<�]X�9�kqᥔ.�6eH��X�rx��T���۸��ɀQg��S'av7�$�]8J�رS,��Iۮ���#n��'���1W����������2�âߨ5qwb�S�/\j��'-+�y���\�^����iʈ��esM�v���sLF��]�ݍ�K(hʵQ�[�ƹ��xb�s�Ouh%��h�z-�ϥ�Շk�|�v�'�{Ӧ-��wA(�?n�3nF��ٽ5��Gh<��hJ��/2�t���ox�7L�8:P�pm�Kp\�A�jcHI&Ѽ1VFQz_\6��䏣1
i���f�=l�q�����^�PZ7�Ȫ�R�d�%�U��Ú歷�]5�{�*�`��ዐ�xf�ڙc�(��hCO�K�WlͷE)w4�;��H����fa��{C_U�uj�T1Wwv!YPd�N�\�FX��N<��ӝ��>��8^���K�L�q	ݣc鷈A4Aw��0�?0�bu �w��[h�G@r���y^�1R9cy-cU����F���`��
=s��ݮ��CJQ:����]0룥rRlo�+�n�zoj��ݾ�<\F�K�&o�9"*;g4���Bi
�Ϡ@�,T;+��S'!�����xn�>Ӵ�5��^�f�>v:lَCJ��mf*]]��X��a�AO(���guR��~**�����{�NŦ	�8����+�Ȓ�Z�w�ǀF������@3��Q�s��n
Wt��.vE�G2��k�%C��ҭ};v;M���J���z[.g��j۱��x�d9���Վ��ka����![]�N�T1P+H��e�v�%�ם��Յ2��m�Pg4re\�X"-yg�4%<f�%e�`���s3:��M.�Q9b�26F��5h.ԡ�Q&v�9Y7���5S�\b �F��عtu�k���EL;�@gv�%����R఍�y���!X�G3N��jgyP"5�3��d�֗V;>���a�0`�gF_<]b}�� n-b6�m"�V����QZ�`�L2ࢬe�APF1����P��aE��ke�Kj���V���RҖ�ژL*V��,��1��(�i�R��1��2��b5n3֫[J�
.0\Rղ��m(�)im���eYQ�08�UF[Eeb�TVڪ51q�V�DEcm������DZ�6�)mb�TZ���
�,�1�kU���ZіƶTqJ���-Z�[JV�()R-F�b8p�
Z0V#-
֢T�
����Q�h5�E*Q��E��J%�ђ��J�ъ��ZTKk�J1qmj����-��*���m����ba�0�m*�m���[cR���k`Z�B�E�e��\R�(��LR���[T���(�DPQ���Qb-���Ŷ,X�b�[mjD���b�kh��-e�
,-�b�TTm
D��QZQQQ8�1V�U0���*�+V�V��&)Eŵ\!�°��H�TQPV*�#RYV6��5��2���
[�A`�V4���ke1������x�<V��v�f����� ��a3WP�޶��د@�8��e(��O=�:�W��b���h.��Nv��U}�xxfMlCN�s��r�~�Ӕ/U�c'w��-a��9J&�����`l<2+���Q�;��`��D�Rr�]��QLt��Y�W��2c�����x�Of>�h��� W�̜�E{�a������\�1`���%We,y����:�l7����Q�%^_�/�.�]�N@i*k�^O�	�#��p��1�%\�cdP"u�<3������R���7}��i�1��H��ڧ���;�;�o�<qc�4���1!��2d��a\+��S��k���`�٧]8�I�3~��lf�>�n��	�S6����r�tC��9M�rW{s2�>����:�!T�f(�F��K#�oC�'���A�=�}cMwJ7 �m���Խ�:6e�aD��`��vT�[���)瓀�T��l+WO����r���+}�]'D��NP�&]�4���	NYޑ,�\ϧ�h�Q���΍��j�ᛞ���3Uݻ�v��[�*O%�.�
U7����h��Pá�������Lz���3bo���ͮ�Ĵ�ܗ����.'���,���cݴ�V����CklY(?1�h�x�h�ݝfr��zF".���P2"��x�]Q7ݣEi�������&Q�o���]�3�"iֵ�탙[�A�ܽ�2��񭊝������{�����[��fX���Ӝ`s�τ��D� ��:��i�m�aw�=n)��ǵ!��	��qg1����g�T���4X�e��wd�~�f��p��R�lY	�%�]�5��.:��}��d(�&ek�m�����,7Pt�wR��ʈ���z�lORUY'C�y��4�E��;#fͻ�
�N�z�f��D���E7'�&�M���g��xĎ߭����՟r�Υ��/1�/�곘b�	z!~#�4��҆�='��Ǫ��1��CZ}�'è^GԬX����ճ��c���`�� o;\Q���E��m����sN����Nt������V��Lx�'��T�MÇ��
�V<����p��s���.���E���+�;���q��(�V��).,�L��
��8Mj=c��{�`���wТ�>��UH�r�88E�����ߕ]��ܞ��on�bw��ĝ垎*.p���&k��l�H��qEl@T�3�X�uC,������@�5��2i���D�^J}5��p:�ODb�t��]�V�U=5.�Q)~Mɫ=����[k�n���#�� -��<%���\�wj� �J-]-�y������+)EY:��U嶠�n+��S}/H&��jt�mU�孖�2�*�E����/p��jZ�P4�L��?oVVx:�g�䕢娃X�,�!oh.s(���]�+�Z*�\��_S�s�Քۚ,�S!D lt�Q�&%�R��r�^tH��7���k}�c3Z������y)��I޽y��8d k�R��J�G���ˬ���A���O*�wt]�F�q;���ä}"�i�V��\�$��ݚ&���$�,���
����\�۷����YӒ��r��g;K8köC5�[K"�R��z^
F|=S�3��X�"��1cvoť�z�U�Q�6ųAU�FΔ^t���e�JB�c=N��:�L�k��و��dGwq��y��C��
UN���YQg�\��)�sc���Qv�N	
�[y���/��h��T1��܈wi��h'���`^:1����vxO���u|��p/V$K�W�~�Sj{;����,�@%0r�ʰ¹����
X�s��$U��W	�/��]��]�3�����Q��b�+$*���A緶(��(0���pO^9�Fg��03I&�M��;�}b�茷E.��"�(W�Xx��F��q3t��������1�r���p��f>�<���k�J��S�����:=&�ldA�MK �C#�R�4L��zQ�$���G��^p��&u&����Ò���蚜�3� ��=��n��|�M��.cG�$b��`ٽR�7ز����a�O����܅�􁡁�Y3֯7�bd�e߹TQ;�/���RFF��d�QZ�_�u��=m�\��5�`w�<k"������E�z1\y��dr�*���4��N�I���W�M�������lz5rfZ�U{�&f��޻èyzo�+�������&��wƜ[R��yx�[ݼ&�]��v��T�֣q��DhSj/NGTr���EVƭK�E��w�.WW�6n�.���#��[|pj�Nr�8��Ω����K�l�B�
iV�uc�e$���vO&,U�����7a̞(�_m3m���O(X9�:���3fB�C�QFz.p��i���zR��95˥�J�w�Y��g���"�7\VFbuE�ʀk��doB��6�ƷLd�����60[<`"1ܨ�o"�u�}l�w<�l�9q�N��Џ\���׏��9�\4�28�ߟ4|/"�9�&Ŏ��(��.�R�D���&�t��"!Tts�w�j��7��C�y��b��{n��.���}Pju��l�Fͬ�����1(�#Qc6����R��ݽM���l���zrE��R�j���b#׌<�'ܴ���T��-���]���=wp�~  !����W>��ԡ��h�yӭ��\$ӛ������߆?�a<CBʾV����
���v�ؖr�-j}bJO��45	�@GA�w����{��o���?Xc{���j+WMu��F[�o��z``��%��k�4Y�
M�c��κ�V��pq4΋�u��Χ���_�ݹ�1Ϣ"F1"'���Ygbڸ:i�]ѿ8�0����m�
b��ku�f1�$���T3�z�;;�,8F�X���<���B�<2.�@nݑ������ݳ7�2�1~��Os�in��>"U���B��c���a���R�^�����������WӦ���Į�X>�61c|-�pu	x��'غ��A��I�Ri��+���n�s*!L-T�N��ǻ�l��:ml���+�$`N�@�������a	������S���,G:l6��-yL�:�u<qc�F��<�$#�xr��,�������
"�.5H�@'��������:۶uë�yͻ����L�XlY���|f�6��<=�����*�}@�>��U��]�����pW���:8*�Rw*�^FN���[ׂ	u4��k�'��i��f:��Gҳ:¹d��e<W�^� �Tޥ"�Ԯ[V8n��;o)��^���Q�߁�;�t��x{����LS�z�j��x�Ɲ��#�L�1^s��y	E��x����'��cX�=�]��r:�t�4r�co���x�S�2z9�t^}N����
��G�EH��
���6Mۃ�NVB���b�)�s�"�_h�:�w ׃r�%yxa��;蹟D�T����iE�.��7�w:[=�O�Y��{�/:哀8�B� �2�5�%�Q�"YʹQ����)�ɘĖʗ�V%E�����y&"xވe�qE^�H�*�x�Y&��:Sk�㺦��3RN����L�����c����'��c�O�\hw3VX����wd�p��Ypp�^���%C���9`�L窴zޢ�w�㦆9345϶��@�).8[u���^-;YP&���\p����@���.�����=oIf���>Ν��Y�P�W(����u��v�����D�~��D횸�C�\˶��=K�s�\"v�8J���s9�^ߊ��|�x�ƚ��}�������~��O޶l���^}Jŉ�#�
�t]Oc��xWv��V�������,mr�򬊾G1��N�9�isk�$��7~�38��c0!ʀT�ǝ��(�޿J�Mm5[�G��|WVccQ˥�����+%�^��t9��W���/4��1g83X��:�����s�b�W܄8���cz��y�'.���3�{�����˼�n�G�I6~��plc���9��Ղ��ދܜ��#6bQ�0���FoVE�:�W��3;��F8�C'���Q��8q�S#p+�;����=��S��7��'=(��=�^��r��*Ċ�P�ܢyU"u������3����ӗ��]�T��4)	6�}�w���4��-޶z� p�7���x'����t^���L��f�j��kU#KST�0�aՕ����%o�Z�41HYQT�n��+�OnU�z�"���i�U!�����Y��8<%\OP�Wq����^g�^�^�(�b�.Yk{�U+^W>yy��śV�g�<�V�'zƼ�W�1]A�]�-R����4�rͿg�]IZ�2{:�,�ͦ}Y���^�f�r��d�mђit�'Ae���(��Q�n!�c��5c��lX�(�fΎ��U��/=J��8%�l�0N��z�ȼ����u�~�f|��º>���l�usѳ^�E�NxK��&YĤ+�2���Jt�h�F��*ѻ�g�V^�5�C̱�[��t��v��O�;R�{� �Q����>�9�����Ϟث:�x��]ի�8P��Svl{!]8K��ցݶ ����������}H3bS�ss�S�tF2c.F
�Wl�Hq���wA*��{��xd_z#3�{��+.?�ohbU][
A�tX���qS���G����'��;B���sU?�ww�;�D���wb��ݏ_í�|%��`^:1�®�vxAv}{K����߀������Yޓ�yc���HJ$�S����� 0�(w��\/.���U�y��n�8C���:����aN�z�
g� ����"^�أmi�(7��C�Vnt�7h��؞�9���f��AQ�jq��6f�S��b�g� t0��xɠ�6�4������k}��aZ����Hq���`�����\Ⱦ�J*"�X�������}�v���{4�㾷)�זQ�F��oD�K4�\����8x���_�;}2�Ћ�@�W��[����߾⋳^�Ӿt&�ط�fG+��'7��"�nX�C��ޕWln�y)�ӽ�3R��w��;��1jg��+Q��v[wCC�r�=7�Mo�:z��p�׭��L�R4�ymq�B^���Y�j�3AM��D"5�)Q�6�=�������;w�ƗSvF����j�j�A�G�)Kᳬ��;Z��ަn�3M�cU�Ų�*��qm�W*�uh��j
cX����ff,t$���'٩��̕�C�(*�^��Ոj��M|�:���W!�����ċ�]h6�:G|�q�Q{��e����6܎Q�G(�9�:�]�<a�(*�k5E�:ܵ֌Nr��;�r9N.��H�%=[g���^t�R^ͦl;��*�n����'TV�<-칣ss�4�G^�4�}�x
+��N���Q���0���l�w<�l�8�F�ND����=4��eӮ��;̎%/.���:��_5��c���G���b�EJ3s7S�e��he�~�^ܰeC#�::��\D
��4�/�N��ʦv�p�c:���X˨�Iz�)���}�	���3E��J
��hS$"U"��il`R�ueS:vw6���q$K{M������}�DR��$���.���k܄��~j��9�E��&�;='�SY.�\����W�LBOy!)��*8�z�m�;�;�}1	�郾Qe��j���wF:^_=��w��Qv�{�D�`�7:	���P�W���d�ܰt��H��V�,�tE'ޛ��a���+�u'�Q~�;r,o
����W�-���c�����g�HTՇ���f�����&�V�s���Ew����^��K/_>x�M�e-�<�S[�'�Y�;�n5�:8�Rn�L�:��-}&t�qs+�?^��<�8	�v��x��u���J06��#�}w]E�wi��%�p�`�_�:�^&Zjq��Z_$n�pH���}�W�x�wsO�ޅM�O�kc�8?_)�ϣكl�wLz�7���\B^/x���׆�w<]�畧�ʣ��Al�_l��;�'����vy�Ç��~`�m_ɽ���u��,�d�k_3�8e�6�j�:#�6ڧ���;����OX���N��7�5ɧUWpu>�^�B)��
"�(Qr�->�n����'���8�;�f�*/e�a�^�wq�'�Lڌ3#��L�ڙ{���6{�z5C�Y�GE���sNS��_+{�Ò/�{���n��۹,b�e��3,�Ҫ* k5g��Պ�ʝ����91��I2f�k�8�.l�5T�k��U �n\B�;��6�/qs>�Ih���ctV���i�C�ͭOU�w "��<��N8�B���M$k�/���%��Q��/78t����U)w2Vt1}{b%�|<8_ա�l� �Oy�*�zeE3�Խ�-70�G/u�?b�;��(��6(k�:n!�;`ԣ^�f���G��Z�xJ="���WY�l�z;@�څi�j?��g���s�/�pU��"�g@�9a�v�Lu�r̻VF�e����so��xn�+�IB��P��ᜬü��R�b��'r;]QL\����MN�����W.����T�������ۨA�i����X�D_�V��q���')�8�.��X�]�	������AjwJ� �]&p9��B��#WHyq˫"h��J:ʙ���5i��k^(I�qf�����oByh2�����=*w��������E�I����S�{,d�ޢn�X���;��)ozJ�m�{enT��Ł�ܥ��N�jF��2����"��tn�;MC��3���sf��.�Չ �$�4[��{�U��xUfjݑ�RN�	N����L4g<��|F�#���5f�,I���\���fB*a�����d�.�L�%S�]0n�`v��HZ�c�g8��yM��)��ͬ�@os�#���B�)��*Y׹s*��,��2��Əp�K�!�B��XݱI>�����]{������);A6�֭*u4+;N�� t,�
�ڹGmK�����!֭�Hw^�eh�X-[F:��r	�$�G[�2�:��Y����WvbF�w>�>�p?h����'	��y
�j�$�o8,S��>G�;��ujF�D�s.�|ꩰ���S�fcZ��o�ڛ�O���r^�d��Ϸ��r�g�zT�[|�:���k��kd�EX�׸:V��|���P�;.wO�.{�fU����vh�B-����c��-��배(���U�B��s�b��Tމl\��#:s�fǓ�2yi�.I�xk{lÏ�iJ�czy69QX ���]3 ��G��J��g!��U�/�H5a�	�}�}��A]ݲ��]ҭ�ᱢ���z0������J�5�{�S;��O\+$���nʎ_]bM܇-f����J�5����p�ۣ�DB2�RX򳹭��9�/J�U�y�goI7\�*��6�ۮ��[_c�6T�A|��u2�)^�u8�HZ�Q���o>'f�[+�"��m���h��^J�i�9r�\.}���.%+�V�|��
)��)T���a��j�����U[8gA���_��+�[�^�&�0f7�ū�F74pйT���I�[�d��]K��oVvf\��J��>Rnf}�e���[��`����<P���Y��x��N,3P� �2�a���.�w�n��u	�ʼ�-�0QU��I*�эE�z׻sѯ�B�^�]C��J�kn��F�j�ǣ��iAr�O�hV�I���{n�0p�@��v6A*��vhW�(Waf�uC�YG����az��ֹ��r�����ZV�[+���@VV�2%ɩP�dʒ�u�����V�^a�&�ͫmnV$ �Co�.�Т-�9�3��]���Sa���]���O<���R�kjQ�#�E�(Z����EJ�*QQjUL%�X[Q�Ak%e���J�[V*[am�b�AQX��im�b�c`��+D��*�Q�"�e(��b#�R*�T-��Q�FL[QPS	Z��UDF�"�#-��T�TTT��* �QUF*(���h�(���h
�-�[F�"EA"� �������*"����Z
��A�Q�R�X���֠**"���Tc������PT`�,P�DD�bE��F*
E�+-,��#mjTb-meF�DUڨ��J�$bJ�U"���`��H�TA"0�J� � ��HŊ�UU��U����Ŋ��R� �UFJ�R ��TX��VPDUAUc�-(�AF1Ab1b�����V"(*���*�b�0R�U�F
�QH��"�1��Œ��E���J�E"�EEX��P`�EET �UEH�m�V2""���"�����m�9��qx��d�Ksu6En�eEt�t-�7�o1�I�|0;��Lq��r������!x�&�*��Az�)ͥ�x{��]�;w�:�F�D�˟¡��
���{�����>��@��%ģ������=�"�t|����ܢ9��-�z@T��v�[\1�&J����H�3<5�>]A�l��N�]v詽��t����Ʌ-w�T'���1g����k��oÄ���Xd�W�Wv�t�U�ۍ�+&5N�Cj���S��~��e��ΟR�`��[:�u���O,�� k5�1S�u�p�7Pxc�������,l>ދ`7GzI�3gYe_>iJт��=�2O��@�#68VO^.���O27<:���{�Z��簣Woٴ7��nѼ�9�V$H�5q�G�G)�(F�{����g�J�v�X�q:�G�=$�����E�t��l׳)��],�@\qH��s�l@�bp18��ɭ:��݋����!�v�GN�����S[h�u4�`��Ur�A�1HY��F�0����-u4� ��p�Fn�~�%�NbF��,�J���+R�;h�>k���ˉY�6�^��l;^����Y�F�6��/Y��`_-&MG$nS�����52T��/��{��b�Z>��Ԕ�)v�l8��(Jr)Y�ّٝ��$�Ch6�}��`�ݼ��c �l)�-�����S/lI�	�Q1��Q6�n�������Rm�N��9eм�(�V�g�<�W��;ׯ2�;�J7$H[�Ϸ0:����H��o���}��@�g�%O}~�+6��z���u�0�J<-٢hZ�H�u3O7�D=p�E'y�m7�}ySL�0j���D3֮1^��k�@�J��8%�l��Nn����㻕��xA�#���߅[?p�S��8��d"��%��,�R����R豺?a�^�ޏ��zke���\� ߩ�=��p�����qS���V���d�f����<���F��<��J���I���u�Ax���K�]���k��[�<'>߫b��1��嘑iA47��JQ�7�a�+*2����(�̳gJۛ��e̪�sɺ28�ӗQ퉡���"��&�Wb,5PC��p����;��\��J�5u�r��n��i�/n��@ʆ2�����E��g���M2^YMě��[�ן,��.�G����GT؅$�t�f�^ݰp�vH�.����\8�;���g�[�V��x�ZҴ��
w2 ,�Un�^��o����Y�/�F>�F�`����+U?9��k��\~[�Oť[����Hi�c�?jM���8��X��غ�G�	em�EJ�kU�!'+�(?����4�[�g�vs��� ')��4�O��/cOt��YG��r��Q.FI��.SC*�5*��{�ϵul2�p��Ӽ��f��V��)D��g�����$��7�F��'�n������zS�ԽR͖wm^b"QzC#�7�M�*�3�ebm���5X����e�(�R4�ymq�K�9�Y�W�Sj-��Q�8����㹝Y1=ۥ,�G\ML�`K��y�L�}��7"p/Փ�/����/�}aVč� We�бy�+���/�YD����^�]�b!t<�p���S6靖��u�dk��֮��LX���ܠ�a�� ׭:����C�*�%:Bι�q��H�mu�u3�we�u㇬n���za�yv���o,��Ϥ����`���J�tap��dE��W4�]vR\��Hd�pΫ��d"F��� U�4�/�i�-�uk	�o���w����K7yAᄥ�u�g6��3�&�
B;@J�!�+&�>f��znZ����r��V:�I�y�J�T�ci.�,�H9���0��{^�U��t�c6�"}D��#��[F�D���T�R�ԙoY���oB;!#h𲰢s�*�7�6����
*��KN�{�X�}[ԝ`�V
�{��S����|���}I\�}���&7�Ͻ�xUȤf�8n�N��\o5K��a'o��u����{��Fx�%����Ff��]��r�V��Kƽ���٫��&O	Vs"���%U�"$v�`�Qe�����EoOI���*��wٙE�az�I���������a߆N��64�b]j��VN{ݱ��gn�ɚ�3�'kA�w�H��>�Ck�T����[�kh�7�fE2<�n�E[���q��a�.v�Ӎ��$c�\�Ŏ��Cs���:�k�(O�)`���61%�]Mpun+���In]�U¥=J+1AQ��L�]!d�S]���\���K?\0c��.49o�{���<!\n�lXu؋��)�T 6�u�.���t0ߛT��guy�M��8��
k�Twnݦ��LV,�j�����hi6$I�"�q�XH��K%9�B=z�ݳ�6b�Y��l3UQ˵���Xٷrw��]���;b�H�{�������]�ƲZ��rˮ<���{oy�&M��"�i�aM���0��^��vT�[���O<�"��9�
j�8v�G�Y^�Nغȵ�-U�-���l�1y�� �ͥ*��1a�m��X��w��sU�}�DB�N���gAX���;}�i�����eq��K�莺�
�橭᷺-��L���|%�I�'��ˬ�P�n���ɨo��'<��v�r�RQ<g���o��v�>e_�m�nl�9T�b}Վ���� lBt�@�onUC�L�r��5�����{�qA��fK�����O��,�l���I���j"�+=k;o	W֢Iz5��{⟼�&��||��
�2�����τ<�2�� R��=FD��g>���Z]�������p��^r8]g��tL#�����zg�]�,׽;5���Y��Kܖ[�;�{�[@����j�f�[��3K�p�Q�C-t�����>��W/;}:�c��X'�m�zU@T5��vF�Qڻ�
�w\���陡�H���d�캍�e�vQ�4���ဿ>G�	���~��ġ�M�J��'�����߇�L/��q-uf��BfI����,�a��Es����E��*�{q�F�@��z�8lL#g�lf����d򛺴�""c�ܚ:2]Ή�C9����fF�:z�k
6�z,U�����[D�z��7���Q�Y��N>���Gء�<Ut��6yÈ��S#UN�����^q��B'_a�1���
���������}.�Z�O�u�v5�b��ך�D�	Z��z��A-m���OGlWPK�#Ó{���}r�����R�P�C�5.��;F�"�p��&��]VF�]�����y�.N�g'�
�RuO��ޙ�+�Uh��^-�z~�J�T��ή���V�މ�C��7D�Vj�0�XUw�����>��͹�F,<�k��h�H�!<6�������nq�O��,/)��+!�Ψe�8�G�5Jcë*��?�����'�z�FlМ��ں�s+M�o���}�:��"�	{���o���'2�5�@��U=C�S
�*��hh���@��0;���OB�j�,��J�$�k��F��t�Q�����jg��Du'�܌Oκ�p�6�كi�Mf�6�U�yN�F`�IFm٢gU�����9�ɺx��VA$q���Gd_E�=����@v�eNʸ��M���{��ƶ49���q���@@_=�:L��
�~���g#'�{Ӓ�gY�g��̤7{�M���oj�����n�N����t���傖��e����O���Qf��GyՑ�-��V��]II���i�#A���X�wa�+*"�BV@�m�7.�
�t��^o.욻���]m��Y���O%(f��"�"4eiO ����ӭ�&2�[�ܒ'���f���:�#!@�h���w��a�Y�+�Wl�w}�e:��ܘ�&7J�)�;vWou#���������\��֓���Vܮ��[+s���>+�'6|5S׽����I88,ȦA��(�A)����a\��c�u�īL��� �֫�7�U�k�v�n��F������؝�����Xj��olQ���r�A�
� ���+��j���rK��M"2�{v͌��X��X6f�S��b�g���I�����e��x��Q�V�y�ܦ���f��i�PNn˨g/j�;�!
������2z���3�(�ޣ���wb;g�Ŏ��zdyv�КwQ��u�M���d�N�I�dqP�ȇGa�URN<鑯×Z��t�c<���yzmŞ#M��l3��⭫���x�}�:}�`�cr�BOsu�����h+�=��K�,�guU�#B�Qzső�~
���(�mu9�f���ܲp=�����˥#J'����%��,��M\h)��a�N���#*�gb+7�[vF�2F�ML��U������7�,�z���9�:�8�&�X��Y�cn*)��o	�Q�dr�\8���tl�N���x�~�Ys=s�l�ݞ(���G�X�%3e^��r
]���Ē�k��p�#/iN����|+��ͼ(�dހ����3�e�t`�|�c��:c�,��w�Ҕ�N�&����[Z�$��6?��;Oh�W��Éinw��}Ѫ��c�W\�����k��Mu�k)��	I����N��yP[u�@��8S�lJt��sI���xl�^=(��p���|ⵣ��~��#��!v����PTE�:GrD��/*�����XJ���y�k��;k���9�]P���
r�.D���\DV��� ��z������Q!������v�s�Ȋ<AP�9ɇ~��mMdo	�Ԅv�U���B��il����!yڠ �㏘��n���E���0Dۜ342�s�e�C�:�;A͚,�U�O��y}ٙKz*��添&`U�\Xf�_9�G�{�t�g���H��v��Y���[��n*Ф.�%�!j��h���WƮe��_��'��#����;�,D�bD�ӝݶM7x�󁺺���=�����[e߽;g����UV(��[�zo���~s���!s�ŔO��˞�e��+\�K��ؕ�d�j�Lv}�f��;���u�֦���=${$����!1z��ڣ������.��9a�`XU5Ӿy<{�=�����+`�K��D��Z<����%Y]�vD���Ƴ����}g"�fpE�\�x]���Ǯ:�]=~�H�|=�*�= �ų�XmH-t�pE�ϝV���Meť�tﻇkz{E��+��v]E���"�}�$�e�v��h:\�y\m�I��e�#	�/��^��$P"=8끰3��Z�0��:[R�9��vy�`�Q���Pc��K.�2T�ݼ��njp�>R�F3���c=�ӎ��=>��b}�wS��{Vjf��V�N�7yH��м���l$xdi
�Iv��V���	E��x8��t�X���9î�Ǎ�(���H�Bp���ٰ���ae�䗆O�6:RU��<�֭dݦ�����qו��<�m�}t�M�+��'�X���� Jr��H�r�r���[4�1w9���#K��7&Qt#64�x/)�,�q��X�D�I苗-G��WMal�[�GfF>v.M0�b<O,�>>_L�������>|$�&�Y���B��k:s�_���˧��>��q�t�{����#���l�R�s3E��Y�9�آ)L��7x&�o]�{����2
�15��<2�:�|qO��g���K}Cw��3A�nG�eu߽���]v�,V4���Մ
c�=�r��L��r��s�RG����z�𞦻J�0���K���f7�qC�O7]����ټ3�o��k)�A�\4z,�.Cd��tS~����f�t�3�3k9trS��[��JA�����Q�
e1]��t��#"7r��>;����KE��}mmƝ����cv������i̶�>�%�j�`���L;�UQj���و̋�'ז$#re2�`�//v��$J�l��ȗ�݋u��*c�?���cSgX��������8k]�׵�X�:�?%��=���of�~�$�c9��cP݌nt���`��8�P���v�d��,�,u&_gvk���E��niH��`�!�<U�Q��y���t,��Y�J�H�������X>Glb�I��+�˗Zk���#ح��bD��8��>��Q:��\Sٴ���Q�R>�qtsÕ��{�����Q��;��QQf��#��d�WX4���!8�{w��������*Y����K:��p� ��4��La��y��^i�mӶC�$8��ֽY����4�S�Ъ�U{aXޑx��ٽ�+�W����`�h6f�%�R��qO�h=Q�\�wh>wY�ŉR�(r���J*�t��+|�a`�Sc\��z� �!��unD�1]�u9٫�bD��.�B7.VEÔ{3i�H��F��o)�(̆IE��+XT&V͚��3tgdUP`��o�o���<Bh�Bjuz�-����*E�p�Ӽ���$z�:V2Q|��ҥ�>�r�:-�tO}�Н/y%9�V4]��뮡y��w14݃9��i��ԏ&�2w�ƫ���f!�]N��%\q]���iDZ�P�]��+���]LJ�خ��N.�d]/�c�C��u�oRC��B]Y$l�vJ����S���s 7/�i贵]�v�ָ��b��C"���^R�l����i�(��u��S���������VW7	�3/zTd㺛A�`$v�{���S�׊���]\�
X�8�`|)fV�]�����N���ż��,���:YX�mv��;��6ɺ�σ�����^�X�s1�p��.��¢�2�5 ��E�q��*kΥ�֪v�n���U�3P�{n�i���n��^�"����n�ge�v��v��:l����e�ZK�z��#�d�n!�adi�6�Â��`��WW>�	�x*3�:�S���C���+���4��B�Z���|��庘%r�\6��tRykQ1��� ��@���<ojxn��*U� р�rw7�$���ɲ>:��Z�'�=���Dp�*�ޱ�6lq��T�@��Ih��s���.Π2��`��M�&�,�9zQÃ)U��|V�wm �Deڮ;&�S��t��ԧ72�4|�+�r!@�[G�
0���l��1G�n�I
D8�5�l���+`v9�59�9�a�h�J��07�K c2S����	�$��wT���s��0�u��u��%�xLQ���g6a�꺔1��O�S�n�F�J�:��6l�����=1�ۭJ���x��D)�KBد+kr�2����wr���
���FuvD[��j.�y�}x=�vI8�̡&���8Ո���S���jD�עI��v������:('�R�'�`V��K�w_oT%�}֭f&����e�Ӫ��4����,(�>u�\���擏��|����
V���q�[�}r��z�?�xWn�k��M�zɲ@����!�r�� �w���މ�}١��Uv���Jtu�C���uݔ��V���yp��nL��0��U�Q��^DS��F	g8Tt��6�i�j�}{)�Ac�!�z���@�x����6�m�gZ��m�|�i��8��#m�9���]ZN�t�n�_p/[q<�ٸb#���r�#���L��S�d�S��ޑ�ڇvT,�)��c�r+.1�q7�`op���F�^&��{�&��[�/*��!��UZ�����pc���&�OkQ� *I!2�iQ�}ʾ�.���\z��U2;[Q|�.��n�b��ǭr���\�����ϓr:$�M�Ru���<��R�7}7;� l�����s���c�2[9]�������LxBaaX�;�Nؗtl�0L��ݕ���D`���++V����AEYZ�m����X��*Ċ*,U�e�(��+A�"(����DQX "��UX�UQP[iZ���Z�b1Q�X�b+�����U�R*��""�`��F1YX����QPX*�Ȣ��T`Ń*0Db�b1Kj�bDb(� �`���2�X"
�U��cj#R�ETAA*1A��EEX�Q��R,UE��b��Q(�*1��E�QQ�E�,TU�@TQPUU(����DTUTF"�PD`����*
�F(���UQPUTAUE���V1EQE��TU�*��H�"#X�
E�(*��+PD�Pb ��

*�DUUDX��b� �U+��(�V���(("�*�$PTQUA-��ł�
��Uc����*�QU��������+E;a�hP���������W�H�wSQKĩ�G��^����SNѧ�+�]һBTy��e�Uї�����Vf�w{�d�ؕA$"���	"��2�k����z��n*�u�Y�4�fߊ�u�m'�R���Y��.�:����bo�[0W_O\�ӋgO	r3�FFSRa�|r5�s<���1ew��v����H�Uբ��.�c\^8�Tգ<�+5�B�=K*�zQG5�l	�#AnFϤ��l��R�3�tcK�-��V�����֎Ӟ��q���xz�b)���O�M(&���M�7sA�YQ�Bő�U�:���j����#��1O��K1�=�<]@���C�0���آ�AoFpȓ:�
uoy�I�5�'ߡI+7=4�ʽ�F�T!c$c��`ٟ^�q1e3�-�S}�"p���r����c����L��vZ�9'{�*�������!�)Fk�X���c�eo'LXf��:���}r��D�8%{Ui)�[xE�R>J�lpuV�(����K��RN޻��<�ܩ� ��lg�:����xV	�vR�g���qH���8*�F�P��I���:�1��8_o`���.z"e��eZS���)˛���r��46��v�رL\�S���:t�
��3�u[�dY�[9�;gtr��mCsz�-@t�ohk�.����y���q����M�]��� 6$/��뫒��7����?>��,l�$r�t'�8kT�Ȣ�gy^b"QzqGB�6�@L�	�ț��5��e�U�F�ˈ�Rˋ�e�Q����	z�9g�5p���I�Pks6xX�s;zC��³�y!]�U8�l\���Y{��e��L�nG(�byB>���t�"F�y��0����@|OƮ<!lz��m}=[g�=:�Ξ�^ͮ���o'2�[���rs3=�q1O��G�����ו �s
��~���q���]����U��!�j/-�=in���f�W<�l�9qmࠬkˀm9��&\��="Y���T)̎��r�TVj�v"4��͘(��:�Y�NY!С���� U�4�.i�;y�9����ᮄ6W{���{ �S���3ExM(6�#�%U��PL]�Ž�8<�v����8f��(���o��^�����o��z`�xK�6�:{���ǽ��sUr\����!t��m�^kóVS>���l��� �ue���{.�w.��0���B4����]��u�{{��3Fo�|z���q��s�+�U�Nď9]>��cZi�:���՜l���I�f�w��ڡ�G�/���%o�p�Q��X$���2�o�*�=:����j&�ML�;մֵw��ڌ
������Ueg| 5\�ͼ����}^�F��TѨC��r������׍,l�ں�z���%��m���N��({��`��x@_0�k�C�~��1��T�߇�V�Z/6�$/�;2��V���o��8���T�H����Ŏ��Cs���:�k�(�Z'O�F�H�FfE��-[G�ك���e����]�Xj��T��Md���Y�`�e��ݝy��V#�ۘsd��l9�N�`�ҋ�H�R���a�ڧ���;��GTF��Vd��}ڟ(�e�7X���M*�+�|��g��X�+��z4}O��:8>Ϋ��uzQ���P��-q�}�=��|�'	B���h,V���g�ֺT�Qz;�5�nyY�,ДX�'��z���o-�Sn䰉���O��Ho�����x1Ɍ��\�Y�͠�]>Sg������V;��r�7	�=��ƞ읖2�T���̄խQ�L�,�)W�L��lUbv-ӮY8a
�:4���w�`�ދ� Ψ����q\�x}�4,
"�Jj��k�&J�w�e�O���U��+Z���O�{�À���!WvVŤ�B�7"
���޿�s�����w�=����Z�[s��d��c��u-P���*�V��؎nA�X1.쩼��U�˃��4�x^]i�uz��Y�ߤJ9p���݋�צ���<��S��E���p��Z6	�
�'=����ǁ��ٹ�U�\��v��Ƹӄ�h��hw3VX�{?t�C�s~����^��\�`�"독m���܊���J�k�S�*���~ϟgz�Q�"fߞ�ՙ�d��\�%��uMu,ߡeDC��H�^���A��η�D�\ic~�T�;�����}�ݙ��J[����\��̯z�bP�&Ϡ�Y=G�pnnM�26�8���b���٣/������?���'״�"��t��51�O��SyQ�GAJ/�}*��^^ڰ׷}���#7P2��_mYcc�Ή�C9����fCq�SX�Q�b*����ڮ��=��l��OURM�;4Ϧ��`�p�d�]b�p�(<T���(tc���1K,Qgwd�a,Qb�=��K�;�3P8WH@׮1C��r����M@�.ٚ����Y�����(�0����Uw��u'x>��͹�F�3��=�)��b3�$6�)�MܥK=��8.��{frK`\�w��2��=jI�]�Ѡ&4�.H��ۡ�r���jwڕZ�/8l�,�S!��\3j=��}��Xi�u����LoAYҍ�=�YΌ����7��-#m�\�]����K�qdo��`st��\��́����ĳ�08gNں��Sq���s��e�-�kV{X�Jgy�*�9��G<��yY�����e[G^N��+MGF'2�5[2ٽ�{�
���:��NnpnWY�*UB7�r�+�2�J*���(ڷ�x�y)��v��"'��8�1M
��Z��0:e����u�Åp\#���>�Y���Tͪu���3Փ�Wvw��BlRvuݻ��0�d �xxv
5��Ы�M~�(�#���g�ä.w"Q	�ѱU�q,��\�L���U@@_>�:LM�f
�jx:��N���j�GK}{.hʭغ�ƹl�I�T�k���N��sT��$��4�ߞ�D�E������t�������+�nzv|����Qv��9$h-���K�����!*�D�^e
�P��ˉ�ù�!wɔΉB��_�"�.`\@�f����NSyVx��DW+De�blV<��tV�9bQ�ʦpл��z�r�"�'!�[�lp�"ڨ"��oL;9v'�F����Ө�A^͞�
��و]Z^ie]�l��[�=;����4Vs�/*��^Yj�
�����]�ќ��w�wuj=N�����,B��7GG5��R=�#Ϯ���h�\:v�(���wl^cy��xn�����QhL�-\���Qc��v��T��.	W�4��ڤw�*���(��.!�����)I�7�����r��8��uhAײ� ��^���n��g�������T�]�9N�7�K���=��]M�p|{�� g��>
g�*��-��lC�މʖdR�pV-#�vK�^s�ً]��u�$��OW9���=�t�c<���yzl8��iZ#�89ID��,kr{R�&����ҞpM�:S��l�'��VJ{#�O����kk�p.��+��_/R�<�86D�-�sQU	t,uM\K���:��:�_h��J���8i,��n�神�������&�z���u�p��HV�M �UtER�ݖY��e��r�(]V�-wn���{̡sq}�N(z�!A��eÏ!cԍ�mOV��N��t�N�wgC��Ƒ�U<��i�*�m�"�:�0k�5��;m�(7����DMq��@ד\�N�b(��b�<N�N�.c���l۹�f\���PW�!��y���oφ>�W�>�K6����b�!�)�P:����@!��"l��8��7-�MO*��;�y>�-���W˅��R��r�-.,\��*�ɣ�_J�֘����ieL������p�+����v�Mt����S�6r{��3�p����춦�^�zo��Y��jz!�,�ٹ�sl���E�o��*���i����ǻ	*k�3��*%�4����b�������8�&�9�$�cxM(6�#�%U�.�-�`�,��=WO�=�&C�=�j.����%�"�	][��(tY@���m���ֳuX)�\�Պ0!���2-�^�����D��(6p�g�]YC��0k����-48�L���P�c�E�u��5஬zB��x��2g�z}k2/�
�2� x���ۮ4({�L���}|ý�P��X�^ʤƏV(��Uz
��j��+�$�o{xc�^X�y8]9�.��$`_�c�����+:t�,�6�s�w^�ۭ�Xn+�g�):b���R9{4x6S�{(��uG-�`=R�e<�=؞���ʛ�3O�IW���!D�c����B���ȠD	�H�E��EҗP��"���OaWU��ȍ&'u�U�b��r��w�]�,�Ŏ��z���PDX�$�E�P����4}L��#Vq�����GE��2/:�~[��rI�=���_;�ji{G���AKP�����0����;{ �@�&�+hs&�Y/5]�o@�$�j��5U�lr�a˖��@�m�^5��{��sɝx{5:�V�	�,�Br�<_j���h���5�J�o�fg*�:�%g,嵐�b}�a;g\:�g��w's�3j0��;1vxL�1Ds��̈:u4O`st���Y��8�5��^�8z��f�۹,#���K�$;w��Иɖ7�X7VS�}����:_d�#��Y��t�M�G*�b=��Mˈ@�坷��v���5�c�����^X�D�*yl9t�:��W�༧\�Y��#,��I�~�M[te[��z6��\��ڥ�p�>SVa����y�xxp�,<�τ)T噜9�ɧ����p�:,�'�͝Rk��n����x:���g��Gt�H�z#s���%��sƯ
�+�xhֺ@<'Ǡd?
�%���xc��J�V�u;�Im#~�xHTЮv�R��e��q��uHu2�B���
��wfH�ꮓ[��x�XR�Q���vg$5��g\�Pj)k��˜�wz����Y�H��Z�^(�e�'��m�K6��X
�9�4w�rL`��I�wOL5���l�=��w�#1��f�թ�X�/0�sQ�Bz�R��2�i�R��{[׉��:�ꕑ�� \�k��GY�R���bR#51{s�(&��ќ���l��Պ�:���c%)[���^ 9cΙ%�߱�e��[��Ctj��s#]3r�208�t�=�(�R��J��~�%70�����YC ����������(n�q�VwJP�N��\�N�*e�䳧���=qb���<",�ىG�YT��F8B�O].��c�6��V�!�g9Q%�'�-ۮ��s!���a�Qb�=��lC�;�8*�W
�B��s��\�µ@�6�#y��K|�t��lg�"��tϱMU�x�Fߵ�0J�+|�[���VI>��'1�i�nM��8ފ/`*��OcX�s�8gNں�ST�0�aՕ����9؜e^���bESxZY�O0�8�C:Cȿd"��Y��%�N�H�n���0jQ.}s�;EЌ���	�}����H�)�3�R��oǅL�Ü����o�,Jlk�w�l�|b���F�������5��0��Å�)l�fN�=g�^]f.w����	�:xH��^���N��o�wǱC<p�T��uA&�e�Bȯ_
����fɩb7v�`��R��i[̭X^yf]>~�k�O��z�#���Tg�!�f��.z6w����V�d�]���U W�9�r%��X�9�����Z����i,��%�5�l�='}���x^I��*L��=R��+/��Ԕ%JrH"L\x��:mU���Y�5�!�٘�r�Y�1�)4�K�NWϮV �E9�wEea��R��\�➙��mv򹣉K�gY�f���pժ�]����|w�
���
�Uul)�2�WF��ћ�4���'�ٖ��#l��w�E�6rH�h7/b���yⲢ!��+�Km�]�Qw���QgX+л>]�U~X�u��Tp> =�(��A�o*����*9B�����q��;��.P�sr��4.�#xc68{
u���{�:a;9W }�Tv.�P��Te�4�k�_e���9%fĲ/}{v��d�B��1���o���[�����^��k�ɾ��W:��׵hA�^D���j���WL���S:24�
k���(��'r��d��v��c�����{,�x(pOj�%u����W�u5��׹zQ��^\����ݤ���,:Y&�8�Q"�s�ў�	�����Uu��:FD�4�i��β��u���W{xo���*b�u����Ce r�
�zS��S�"�9���F��nM�Xʐ�e�f��M��p��rJw���lW��[:8�])Q����/T���Fۉ������9�2���Dݭ]Vm�GV[Gc3�ex��PNƗw�]���
f����-���)ż�-s-�Ջj��)J�����3d����9�n�|��u��s|b{f��-�Z���F�K�o��y[|�펂���"��ѕ�]��8R��{���D�^�t	��|\l��H�:�f�
%UխA�=gL�w"m��^�z���`�pu�bS���C8s���u>�\��H�%�6����+��>��e]�w�g�Ҵ�p��8o:��"yl=�D��m�{����nxz��m����c�W)���m�
+kts\�-�M�[|'>\qv��h�b��	l�J�m����l�U�{)w5�ñ��7�|5������_<��d��zk�ͣu�S��^e���4�tP�>�*�0ĕ�b��:{��sxK��m���5�=.��Qn��t�8+��
�`aFe]���%:a
˫�2�I�6����]CS���jrv���Y����@,6h�<�C���!����m�.�.���V@@=)l�ԃ �e	�+k�����c4o��d�ms�k_�U��@,�R�g+�[%�/r]䍭�����g'N;��;T��_�n鎂�)j`�Hd�61>6;�kJ<���.+uD;�,���m�Ҙ$'��DT����)��f�b�t��r���{���̖�Yr8[:�s�� �v.^Ҭ���oJrl�h�����ՒuI�n�:0�c����t#i-T�n�-]��ڲ�Yˮ�6�C�o
q^���c�Weh�Tȗ�k��P�!T���{h;�l�K\ή�I�m����GJ�s(�v�Ԡ`f��n�|�nb�5ǽ;�!��*qB��-��t�~�
��r��4� +�c�#B��SF��~�b;xOs�����Ht����*�3�d��2�o�`��m�]��x7r[+h���<#��O�ؚhh��n
�ge�f�ʄ��0��y��Fe�X�ڒ�u_mР��nG�[{�ʆs�u����l�y��:)ǡ_UЅuJǵɎWK�����=M�@���Q�T�:뚝���B�'*⫘�edh~b�ia�R�M���J=|��SX�q��7j�_vvϸ�$�����h�V�sr�Р]���N� �V� �q���?���S�Y�˾ϗ03R�&����e ��TS��a×;��ʺ�t2���ܙe���	��`A˵b!�Ɨ,�t���(e�"Jn��\T�Nܺ[՝m�[Ӓn�vod�)軙e1��^]mv��ғ��\�[��9KFSYUg*�zZZ�^�Y��e�β*q�B�!Q.Ȧ�V٠�R�l�e�]u�-��pl��X��lKN-ض�	ܷk�C��j���jr�+���?�vܫ�{j4սn����?I�:�灡D�GL����y<F�Y]����3�6����'��[�l8�e�;�;�f%Z�;bM� >�RAX�TYcE�EQU���cc�PDPUUV!�F��"�`����U"�1DQUQ���*
�PTF*��QF(�(����1�D`�QT�b���Ec"1�H����EEe�"UUDU��QQTEX����Q"E"�1E,E"��E�*#*EAQ ��TDX�"���b �(���("��(���b+Tb�1EQ�����#X1��,QTF���+AU�QX���*��"���#Q���ҫB�U#�� �Ec��1V"��������H���TD`�TE��b0X�E�����U��@U"*Z�,Pc���DE�UEQUUE�����%ab0DDQUPQcX����AEE �I�>��T��3��U�̭ݽY��w?�丐��w+��v���ͭ����S2�qW%�'ۧ.��p���ܳT]M���t�{���:�8��p��HWaM*��s�_����x�~�����K���U��$�}���a�'�,�D����lÈPh����4G��kO��d��YC$��=�2�+yY4�ym��f��q��WX�G�κR�u��ْ�
��^�\4�:h�L��uo��rO]Yy�%�<U����Q��˧#�,�PV=�.�M�����b;�1��4��f�(���]L�a�%ȩqC.�tL#�e�t!W,ˆGz
a����[h霦���u�0��R�EtC��wr�����и�e��.��J&��}���N/�Z���qF���z��rE�L���[&׸��0[��x����Qp�8�ް��n������*&G������{hjjW���ԇ�mI��Y̊_�ė|
�RACe������j]HH��m~qe��j���.�ی#��n4('�'@�G*��b$J¢��_c�vks39.;��9�Q*�������]���{rYYҕ�G)�0y<ٝɽ�&iT�z���	���7������IB�7kp�(���O7z~x�L3��Os�+��1'J����a
������]J�i]·P�tWԴUXi�--���j��K»w�yZ�)d7�)�kXښ�SX��Z��z���[L��{�F-6��C�L_�`zD�ՇNd���H����F��}8t>��nYJ���>���r�_ݢZ�UR9B���o6[�����[T���k��i�;Xz:��STbm%�TH����n!�J>��J�JY��%���+^R���C�p\��V�r����yB�J1��{��0i��Ŏ:OL��CS�?c8/Ʊ�WN:t7��h��6.nn���n�!*��'���u�;��⺦/>ޮ�1 ��!n�2�����tͳ���t�w�e9��o�{G.���͂�r��'��cX�<��<۴=W\W���K�4��.8N��ɣZ��<��w �N�HEO�6µt�M�+���>��;��q+�dM�θ��_��;�2X�*\-�^g�%��tT���"��W��x/:哀8�C����7w܏u\�$�`C�$kb.T�v�R�Qq>�����%Q\&@�<8g��>�N�.�v_�:n`��G�� �{�t�k�俛����x9�1��������s��`k�[�ȱ�D���'�-��=�~.Sw�pW�wT��QJ��nX�s�f!F	�Dĩ'EǴ��(mh��<�|��ڵ�*^�x�ݮ��uS�uLGU�n�c�ة�6n���mUm̒F�m��v��ŝ��\�ˤ�E���hćn���;��������zg�]�,߄+5��GdX��{nd�������
"8iaxD�-D���|�fywO�ZU5�� �A�@��d���zzICq����v��o�g���+�{�N��Uﳧ�f��ȉ�0kܤ�؋�S�]ѱ�M�O��2˱L�C�͸M���r�Y�V"�o�	Uy��`�g0
�c�W;��051�O��Q"Tp6���knҬ��o�.l�������j���U��8з�e�Η�I�����<����o]E��lu#e'9�v�ܢ����E_���7�#6niMeR�#!@d��Ь�0nY)'��l���p����F�
�N�g���mb��O)B<�f�n*T�WPp�5�L>�T\�ۭ5k�oB��,F�=��Y[�-�j��-۩:�QQf��#Q>�(��	l�l�U�m]�Dw��xO�򧱃X�uF �;a]TL��8��&�\d��pw��U3/ut��\q�Q*�[�41HY2V����"�1	{ӜčV��<*yev��%v��*V��`yJ/{3�m	���Y�NLُ��8q�C��65�m�Ic	�kQ �]{he����"�m�����z����o|3'Vc��T'=i$-�:k�Jw�D{Z���ٽ�bs�+����i�n�t�u%�	@�*J��]S���g.Sf���;yy��'({�n;��{*r�p�-�"�J*�+J7�o���Jr\U�͏t�2���R��L.̂((d ht�Q�$H[B��
�a�=�,��6�{����#
��y}vm��s��d�d[�D�����הiWYsB�M~��جo[c���N�j{Qo�#C�id^R��	wO������8��V���p�૥�yخ��TK{�(.yh�d�{T�CM�~9]u.��OyWG��Q��7碖�'Qmo��@������<z�Tl���;.lt3�aE�6�F�M�ر.��²�!���3b�<�!w{���]p���;V*���De�9���S�\
������q"z}�����V`9T��}���� ,�(JȋԸ^[~#5�嫆P��)����7d��T�<ӵ�Ћ�Z�����auA��(�Zv�¤�M�rJ�ɦFU��7b��{���o�o���އ��W�� x�}J"�,�z0:t���&��ۓF��ne�]��h��,�Z���0�y8/z���p��vb�g�J�Y9[5o����"���8�E��
�٩]�]Q���[�c͒��m�Vޘx������λ
��	.WV��=��Q�h#_�_V`]u���7N��q�wB��Q����X^�=��]��r/���T3!�֕3�kk�����ehM|�G���[�4Eo!#���*K�Pl)҉5���)������6p�1�=���ۋ<F��DPb
�������c=_n*�ٜ�����(�[!h=)�֩�6X�6�u��b~[<���M�����`�b�3h�G7�:�S��u|�<e�>U��;�4y����A.T���Ԇ��(B��_��y���қQh�L�:Ù!lX��bUtEb�^��,�Ba�}�Jk�JSq|_��J5����:��OB�!�ˇ�B��#d[_OV��۞�������l�I�S�c�Sη�}\E7<U�����B�`�z��U�:� ��,�{����9�b<�QW��aAo[6�<�2�u�u�O�:�(����a�w=�Z��T��m,:�J;B���b0�]���9���2���{��P�P�2EG`��|M�Vfk���S	����E굄�CBʾV��xL���Eq�J���xSGp>8�*n�n�WD�!��p�:������p�Z�>�sr��U
T�����m�.��������a��z�e�:�*���
������K�l�sV�&5vQ�VQ� ,P�ԥ̲fVA)ٴ�|�^����*iUXW˹_
4�9TF��u�B�[�����e�~\��/�+	;h���e�:.6���8��-�<X��m*��٢�����Ǥ�M�Բ��Z=sIg�i�?A,kkB�/�Y���o{�="w]�o�,��m\4�.�ی#�zM��ROf�P�g�%ɐ��Z�m]��$�Q�Sō�"F�(���&���Nˌ��G�{�a^])^/.�6;fzg�z��.���3�Os-`~"W֬s�B�����W���;��ý��mU������܌S_!:Ex��;7�r�h�w�6[�{(�	����-ꦺMMr�1�X/�M����]��{���S`�n�������r(:��Δ\^�.���^�u�l[r�]�717��a|�=��yL�`w�4�OX��ʎ��)�"N�p6��Ä�v��P���Rg;�0��n�+rt�	���b}��3�w�͇6�N�:f�a��v�L�ׇ%X;���kCuښ8a��;#8�{L�N9E��H�k����mM���0�誯�����R؝�&�dm����+ޔ��t[*j�T"�j�It����&l�m��<��Nn���qXyڡ�j]mޔ'����tc��B�郴���Z�PC\u�I�N��}�؆�=����Y��~j�i��q��-����f�O*�{�'R�r`���JͱJ��!\
��N B*k(*UOzl�9ԡ�O�T���*/��aΎ��[�W��N����UC��"�B��ܙEЌ�ҽO�\�P�:����\U;�b6�r��ݐAr3�%��P!��\��k�ӻǫL#Y��,��}Esmh��=+wǜ��o}�����ў0K�΂Q�72����������~�n�zb��1�3���&�\�P�Ֆ0C,�Wd�U���d��3��s�G����:��N��z�lF�d3,k�o�r��s���f�eDC��E��u� =c'��*E_p�AS:��W����\*}[����58L�"�rHJ	���na.1yU��xU�4�,��bP�^X��_S���U�8%U��^s �����Jzc<��E�]L����S6�痺%�(p�м#�lAh���[:'�1յ��$��g7pjOk2��/�ڪ�S�������<��^�Ц���4E�����Hc�(�)a���9gpx��aAu�]��FP�k8�i�}%c�ԵW�9m�����7���<W
*36=oB{���{�Z�:���M16��>D@yf����آ��P;�]���p֪��x�u�c���{i0�����U�����7��rgp}�������9t�f�~��.�])���>��^��)�c�+�[���euX]y8�b�uq��DX:�\q¼�}�Ω�t�08E���g*��ݺ�����6�)�m隝�9�RHjY����&�q�����l��=��%�P�8s��F��)�+#sH]em�l�=���份��w=�͗������r��V8u��'�͕my:���(�Jo�Lήh�Y��l/&CQ�ٝ$�d��`f������ï]iF·��<���Q��T_cJ��2���kd�z����J3dH[W�GY�g G��%��_�,��rzx�L�X�2�2�t��֍��fd�g޷f��]PI�Q[`@��/����/{����,U�֮�JO�(�v�a���e���K�O�����gI�w��������α�z[��8���<����=hl2��=.Fu��i)
�s^ÿ/J~�k|H�X��r��6�K�lTJ������9QG�\���v\��gz�]�a9$h4��r��1��qV�q�Lxok��M�W��,G+������b�)�k�ږ*�N����i��b�xgCU�;B�u�}�n�t�!!Z7R_V��/��,앆vT蔾v��{n�I\22�-��>�jc�aDE��ӡo�r�Bї�.F_Z#V��r� ~�udB�	k_۾�����u|��p(�|@y�� R�ߋ���z�ˤ��/<��M\U`(Jȱ,J9�T��܄o"�.ʳ������R���y�L�f�V�%�����A���i�<T��C�VnxM22��*�3�ω�G-��O9��|��J8���҈�yL�`t0��xɠ�6�յGzo��v���k*��:p��z�r�UpwQU��)gU+�p���ҝ�F�����e@3k��kj�^��<Y��z{"��R��M(6:t�N+yM���F��vC�:u�����ċ�Goq�삈��!=qbRQ8*l�[�o�{(���Ҟ��j�9�C�*�s:f*�6�9�;�DZ�Qzp�ꎵSAnU`<jԸ��)e�K/��iF���qB�ښ㕯2^7��찘��pr��ӆ�8�/�Uj\+g��g�7[)v�7����X+���eo\ճ�2��o�����Q`k�{��,k�b|���Ä�ѭ�F���p����}y���Ws���Ѣ��Z���/x%�=�v�d~�j>��[*�Y݊�Q|���3�Q��5r��<c�P����Z�̜:�
<�)���ܻ�M;B��g}��]DWR�����R:�Uk�WK�y�i��:�s�kf�
�[܉��'Tm�T�^��fþ�"��������naA����y��ET�idE��JT*�X`q�X�G�g�.�[�͇s�&̸Q��Ʃ�WQD�K���`46��;��/b��#���й�;��E��ot��#��pȣg�%���O�y�J�#s�� 1|�(��(��S;�,`u��A|�^���6��cS��R�jN379����P[��hOU͞�:~��K>�[���c�x����0)�@�~$2��Û�ztS/�;��Zb^����sf�7�Rn��{&�O�f��|5�I��b%���k�1gY������}�H��LQe��\�r1�A��9>���|�^y#	�w�y�\y����,�Ƒ:Ĉ�U�v/�aߡ���`CD��V�[4�����پ�8������,�͹�d���Aw���x��tks���6�
���׶��̒I�	���缋���͌YM�S\BU����b�ә7�P{t�tH��Ѩ\�]37.jPlvؽ����5-Đ)v�*
k�Wb4���V� U�S�:\zͭ�}GoOq�Y��"UL�����	i���J�nut��3@���"�>��
�3���w��:@�`d|e}3>���9�%Y�,tcz��tU�?l<�q
t�P����Rᅋ�V����5�X�β�T��YhJ����#��2
�s��[Z�m^mJt��h�n7V�w�n��ewn�k�V�U�@l`2��.���F9�gX�՘��w2�ku>N�k�E����.�p�&TH;�@��Nm-�-���wH��%�j:����̠��+-�쫑�[�P/
/����M��E�%��}V�$�4�v�)����͝���7�����6z`el�9�9�&�#F���m��p�^@�j�-�yE�w1�x	}d�q���F2��K)[�'�{:X���ӈ��ν�j�@�7��P�\L�[�#N�;[��q����v/%s�j��o�0m���T�Ä��OQ3�Z]��Ė|���Ӌ���˨K��+A�U֠g
�Z|F�W�0���C/��P����s(Ɠ瓥�1�5'xf����:��ٮ�ѷ�m��e���'�U�R�	��������W��J�b��	V�vWD8PF[ӝ@]���;��q�+��2%Cf.�����6�i�"	�Vl:�0m�t�
�H<�"�]5k���V�.��mіVP=$i���pS��n��ϝ�#!?@���v��[�y\r���5�]w'7�މ�cB�}���C���;j��"�.-��q��K��D6�vn�6�Xw�9�(�>���9����.B��ԣ�kT��	2Ť��k(V��j��EXF��vSK��xg7�#A��\���z��Y�!,vY05�zm����%1�ō[j��8�5���VI��:RΥ���f��R�F�f1Sb�q�ˈ��̗�����c;6�i�+�ӜQ�$qc�?u��"�vY�5d�.�q���%X��f�.�y�/�YbloHt#�{�TU�CEJeQ�Gs���ϲ��})^�J�AV�]�1k���k�\tA�GFa�(�>8]���*9��J���}1��)6JZ��>��u����-�XW6�/;o��T��x*�To�f�͸�'$<{R&Q�Z��Ƞ,e�j֒B�Ɖ�цV�n���7��Ni`V9R�U�X�qI��VV�23���2�kTʲr�p|7J�L]yn�v'�=JP
��L�^��Z��M�	C�3��e�]���a�h�F�mp�!A���N�H�M���<Z{7�wf=y;�5�}�mΝ�y����"[�"2n�`<�fSM��V�pn�������Q�Fۛ����ݨ��Sp4+Q��^�B���h��)�Ҵ��+u�J��v�Z�T{�l�X�E���|�oU�K��(wvkI���
� b��h���A*�!EX1�UUE�b*"
�V*�b����ȱ��1b�F0U���UVDQTDV*�Qb���"*�b"�QUQX�#Qb�X�K"1b�b�A���F(���1QA���QH�l�DDAEb*��b"�UV(#""�b��H��DU�(+U�V"�Ȣ"$E��F �X,Z��Ŋ�ATF(��EP`�U�,DEV"�EDE*$b��X�
�1��k*ʔE�*ȌcUPu���$�8�35���h��]�!�:VRoOrZ�J̌��4-�KU	IS�ڝQY-��:J���w:���`W�]�]D�$�9M=���%Ȼ�T�W��~['�o�W�,H�DN�@�B.��.�V�K�a+n��]goI����o�����;�y�M��,v�z��.u¢����}�e��u��涓�Ԣ/#��EO����l`�'���8�z[�S��/��$xfcv�8lt��^o3����{zŔ�z��6S�Q~�'��cX�<��<���`��a��K�z�'�-n�l��Dq�N��du��
y����a_���6s�+����I�ŭ�&h�����s�U��3��WF���Ns;�C��㴼�W��x{93T6�y����og1�*W7r���1P ��$k�.\��D��x������a�騉�W�y�Diz�Zt���,��R�nī�x�� �����&�NKn���r8I�bX�$Utu��8M���J$�G�f�s5e��=A��,�,5��Gd\Գ�s���T�������4�֊jT9�c��3Z��^�@�).8X�4]Գp��!ߏI"Ϣ5�ʅ�6j�\C�&��b��^����/��}xc.�;M�Юn`��w�;q�gq9���b_ t9`�۱ى�¡ÝKT���l=2A����:�I��۷p#�p�	�&N�C^��Ƕ���pA��f꫊EK��I,U�@������� .}ݗ��~ܖ��Y�X�{:vfk:Q)=��+\�K��R�\�0r�Y�;�ޑu����FV�2-�����xp�i����@�����G�TAp���j~\SVGTwy�{�ϻo%9[�%�xG�؀�[:��YC6t��D��Z�(��is����I�fA~�[M��v;��˕m�����f�D�W�R|>_;o�O�_�Q�&�y;���"gy��bЬ�n~�*dnx+�;��N�b�oh�8w�r�C�gk3�s�£w�܎H�XQ�_����9��c�YZ��pUw��x�Og�QQf���
���\�9�]�rK�l�M�)��8�T�3�ĳ�08gNں���" Y���a]^�w�=1��AՔ�%��YD�������޷��oH��Kޚ�S��5�]kѳ1]��бzë<T@Q�]�o�?F#���˅\��KxQ�t��q�8���-Wwx�ު� ut��I޽y�Ex8d k�R��"B۞��)yu�Gˆ�=�.ԭt��]�z6�fTL�������}6�'�p��6��rBd�gWU�qۉ���n���h��8mX+�V�kO�u��/7�-����Ƴ+��u+��GtJ:Uw���DP��G-Q��q�G1�i����������v�k��yoa�ܔXz���u�3!�Q�[�D��N�Q[p$,���;y��\!&n��S�����)g8�6w�C5�id^
T�a�bQ���2):���	�DeCI�4�3��7�D�=��4�xh*�q�[���%�ΰj��%!\1��>��S6!�DG���+�)��M���9Č%(�R�%��,l>8�*����w(�f�rH�i�{-�Wݵ�QN����,�-��Q́JȰeƌq��vxJg��|����8:�]�X�b"�vκ7K5r�$���`��YQ�B�1oS8k��G��p���T��~���{$϶�w�����
��F�PD���F�Zv�¤�MÒVnzi��{v���D�)�.5d�]�ȍ������>�t�/S=E�:O+ojMhQޛ�9'{�s{]K"�
	��\��;.Ѽ�!
"�P�T2�J*"�iS=Ѷ��ߜgF�}+By��ꤽ�:���n�.9t��(ȥ4�����428���X����]��n�~z5�T��a^r�i����4���fOU�e�Ã��A���-�Sf��ɻA�o,d�Y�RF]���Ol�?%<%�C�u�Oe�eh���ͧ��v�7d=�I,�0�[���.Vo1�Wm�����w�h�-l�*�њΟ�D��+^�U�Z�h��ԫ����̍�ӂ7�˧qК/�H3�5����~(���zS��.����������6,��i{�]tB�QzC#�5LH�UXP�7����k@������x�Iׇ�]��f�9�B^��s�y����Sj-�G[HWa��u�s�xO;�}�F�_����]&����iV��j�i�nG(�byB�$�5�2�Pt�Q�@���^��XVF���:�_^}��_d�;���f���w��U�\VFbuE�ʀjۨPi8{'��Lʻr�󈧹����{D2$
fGP��&����&kz�u�lʁ���(���'e�\�$�^쑡�]N0GE����*��2�gf�C�B:�Y���n�n�g%+(����f�q*S�o�*^ފa3���g��X8~Y)[����/�F��+9���:p�1���B;R��F�
ɡ^|�-��ܵxS:he�3c6`�z��vl�T����zp%ˆ��,�k���l5Pv�٢�p�=s�S��g>��sWξc��6�/K�E;5�p
)ָb��Է��C�R�.����h&�'3��[C^������������F2���~��n���ђ����!�m)¦H��;��'�������iZ�vS��2^�c����Q�z�|:�={g�joU�(����-q�s~�>���1"'���Ygbڸ:kϲ�0���l줱�3��$N�Y�{̮��]�y���i|k���zݫ��DۮM��p�ȯ�o}P��
(Xꘁ+��d5��ź��δ^h�l.";��
��>�j}}~����7��f[�۔O��F���'��Y0m� ]��H�겁��-���] ��w¼��5�J��^���k�E�9����q�u<�����ҶT��e{b�,N�@߆t��Gt����]����4�s�ߣ�6j��ה�s���S�;#I�
UE�6$Owr��/UUU�z�o5rXr�8g�WN:)����lf�>ΰݳ�0;�f�������]dX�Id�3M�]_Lζ�^K6-��
��f(�E���P��͔�^�<t�b,�7��t�8"byS��unr�e�^����O����O����徵��T�m�~WO��dr�ˋy�Yu�1M��9��J��]w �R�%9gxM/E��|����yl9ip�5��-n�_�K�r��D)q��;s��u�d_4�c�bϽ�}�dk������vë}Q#|K���
�z�ƕB-�߯��s{"qp}&i�ذ���F�[�;���t�j�r����/j�`�Ĩl,�.���ze ����9�C+[ڽ���î�w��͙�[�<�q�*�:"�5��j;<�x[���5fG��B-I���_G�=}z��̃���Ӝ`q��%R� �+� S�GA��iȕu����ۍL(����epN�Q;�z ,��FG��;`�k����C,�:�%���p��R�m˞ۖ�G
Bk.WRi�}c��5�r6fhk�o�{��-���:�d���o�ʈ��d!�K���(��;#r���.�¿d��ٙ�oir��\�\����{펤��B7���n��d��5�ey�����T��p�^c���7��S *����
ց*�=:Ovk�c�݂����NW���b�xY�+'���ճ/O���_<w�$��c}2���&����-'�֝��c���Ξ��,o�sL�=�3T�`��>��|�.��-�ɠWem�Z*_kP*��8z���0�<��<R���ӻ��ը�\��)��V�d(-�]~��Pҭ����ezL���t(�>��Q:��'���g�u\�+޿D6�1"����4l��م�Z�h֬YAk����T�Oy+���L)R�-B#�x.Q��݀q&�G��C��h�.*oU�x���OYy�Vs�Lvy��У��'�]���6���*v�?�d�rLn��9/�ij_T�js�.�]�t���N;}�5t)5�μ�˃����[|�x ��^G8���/#F�,��t�ʱ(.�C��c���o��`�.F������=���U�Q�qg�!ol Bސ��c��e����(篩�9�������t0L�[2ٷ�5ѷ�M��ᓕW�®U�%=��k�-�����ga�*,�c/�����M�w��� �ǅu�w�J�"�xg�ˬ�ΐ]�d��5�T�1R�/�⋸}��_�Z���:���u�3!�Q�n�V���@�������;F����<|��%{F<�<=,�g�Y�]��[K"�
T�a�x)��3��S
�fW����J#��e���k�쌨`�9l�Ysѳ^�E�N	r3��k�HWK��:]�f���z���M;��n�u�@rP�#B�S����p�E����O�X��i�͜d���N��;�Z���U�{������g�u�O�=K�ς�юS|)B���2�b�����1,�e���ўB���{��B%��Po*����BVE��nU3��܄h^N\�V��tֲ��i+��}yr���oG0�@��S,:��v;]v�޻8�_oo�-4�d��(J��Y��{�4�j=9��H
Soy���x��GŬJo:����J6��/F����<[�WKV���Tz�<��>\�S�r>��]�o�{gT���0�bq;x3�ـ��iY7��[UH{{b���퇅IΛ䕛�L�u<	�:�n]������a@ʎ2F(���7��F+�v;��å�q��[�ri�9�ђ���� +�I�v��}��id��׫~YG�ΪW�\0�7]�;��K��"z65�Y��6M'�϶��5Q�F�,��,ȥ4�����5��W�$]��8��ș����q1T�o^a^^	\`�X'���>=o��jPOW�@�ɸ��DO-��&&�c�;5�g����������t�gv��"�M�=��M:쿛���]���[��j(��������<܌:j9m��!�J�9g�U'x>S��z�
����e8�i����GX���7K�������r���w*�2�����ӝ!UZ4>Q,�׺�����)�������Y�zvF�eަl;��*��qY�N��kʀP�M0�ł{E�Wp�7OWU��X"p���Q��Vħ_:�8��!�k͞g}��ayLw����v\�2�u�6��ɦ��d2b���ۻ�톐޼1���m�nd�=�۫W�i�c���;�A�;�K0�E�`ezݾ՚�F�O��2_wg:W�w�����;�ܢ���XuУ]o)Ή4x��ە���#d��:���te���ƶ�սp�s���J��yHK9p	Sg|Qy�s��tq��M�f��l�u�w>ÝSeҞ"�D���ГN��>&|ߟw�~�a<4,�1NL>�]�5���=s׏�X��h�u�I��pƹ�\!����}��^Q׀U3��^�.�H�Pr޺�������R�1pC%���E�PX5�K�6�A�l�d�5�='�\�+6sR�{�=n��p�OaZ�7��s�=�H���6��;T;��wE�"�o.w�_0��ơ\��s�f1��%f�T3�z�;�ݹg64���"&�[�J-��y7Ǯ��z�1)'(f����CTßR�9mp���J���Վ~H���H�&�]��i����Kv�(����[�P�Ղ{q�,N�X>�61g����P�x��&.�o��n�O�M;[=�Q�΂��k�C��ܞ]`�4���6(z��e*t(����%�PƎГ+0q����IcO����
]C6#�-�y��g��6�;i=R�HDU��]��-���*���ܑ�M�fEȩ�7���,]���|���ާ;p
�w�Y�|D�G	G8B��]���姹\幓d��Q.�f�^��5�Y֞�Ǖ�_"�2����'Y���|��u.�-�H�����Lk�S3o�,*�s��)k=[:��۷���rT���D88�Y�'��NVGk��n���3nmܝ�`M��jnf���R����gz��;b�H�\b��#
Q޷�����X�8Gk��a�s�*^9�$�-*�,��l./&��CK-FL�;`R�* u@�B�y>Ew�6µt�M��Vtv��.��w8B*��G���w �r�7	��K��\ϢZ*yl9t�G��s�㓕�U�>E\,e����N	�J�
�7�q�͕=^��Ë��x�Vv����^�u�I�� �<q�08����G ��{��%�s)��;ɽ���BS��y�޸n�]0↹Ӧ���a�f�g���,ߡa�5���BV�k�yk:��1Y��ʄsn_��/l;�K���#fg\{w��|���a������g�pfl�����s�� U�]ѽ��p�5��;C�{aX��r/\������Ip��� tL*��׾�g9�#�'n�&���<��\U�'oÄ��꾝1CUy �s&��;*�����^hnL�۴�2�n*w)�]�"}Iv��v�vd{a��-������aGv��^F�]6���ӕ�g���K�zT� ]��Y�sE�eM,n3Y"�2���Y'oe��=:��ӝk���ER�.�X��e��\\�y�w��z��ua��n��ʅ{}���.{ٹ]m-@4uS����ы
��^@���Ԧu�7�6�
�2�!��	]	J�̤�P�%�"�<jZ�6c�
��w��R�<]����}��+�h�����t�"<�f+��fA�{Hs9f�Ϯ��}|*	rZ��I�{�_d�&^Z�;��Sx�V$����,����8�c��e��M�Gy�Y�[�h�ѕ|����L0*�{6ũ�Wت�7^��;1t�J�5��;�^��lq�y���.�LRv���C �[�W^r#�����ڵ�y�WA�E��pU�!7������p�wʱ��+c�g��E����V�3[!N������M]8El嶊��Jg;C[���t(�j���7����!ݕ��f0�Q����|���r��ku�4�EC�^̭���K��`�{���t�9��)����5��-�ǃ���EpN���²�^�zM��ή':(n��}QoXy�p��-1����s)E·�:yke[r�9#�Sz�F�jA�e&�e��èj��"��]C.F>�������ӄ���nL%��fum���p�I�{J ��X�{�.��a�WG4g�e�;1��c���3er-��9iᙩ>YdYCwm��Jee��k�]7���ZHK����%�J���_�0ؗg<��>˼xdS����J�[��r�҈�
T������aD-0*��HV��FI.�^vS�9v�d�����I��� ����屺Z��'O��fy\�}�!��xt�Y�a׏�Ѥʽmaj^՞���&L�ʬ ����_Vt�)��P��S�S~���J�s����3h#+�gEG��V�8L�}n�3x�6�e>���u���0�&�(܂�����̺O)�@yF���F��u]]��T��4��v�rO��9��hR�A��y���۴�Z���ۻ�V��$o��Ϣ�"�AM�kr�28<���*�32N��7n�rwQA.!�E�:�����Z�e�׵ovp�2s��9�J�V�U��_mA�(��̧�N�\~x��ŰJw�H�-
� ť޾tI@MbVp��|Nȁ�3��+K�v���xb�klq6r�S�����q������ݛ	�T*�*�ٶm�p�30`�wז&�q��Fc��'s~�L4D
ݠ�NL*#T��[	0S�z�z�9u�)�:�/�-B@��I��JW*4�%ֺ�U�{�b�q�t貢�b�Վa2o��R=n�]����߼�<�4A"�QX�`�"EF(�"$b1Q$T�1EPEEUE�X�(�kKeQ���%�E���Ab�*EEV ��EX�b�AP���*��1TX�1Xʕ�ȱEV,`�TTU"*�0E�����U�" ��EQb�DQA�1�#�*
ť%b��*�AEQV
ȵ�***,b
(�%Q*�"��[UX�1U*TDT��Y�QX�l*�[b�ʑTc�$EQJ��ȶ�)-��b�,`�UEqF�PJ�1H���QEU�
T�im�U�ւ�*�*��QAcDA���ADD`��ǋ�J��/tJ�����ɓ-I�Gh�t��*��l�t�CURY��g������'4&�Ҽ��yZ�$n��Y��n������\Ixk�Zc����*�ۍ�!P�p���pvj��=���G�����1�����m]��(��&���poP݌�s��5�}�*�tw��,�ىD��5�a��]�����fgp�28��K��`�^x���֝���<��<��vTk��:�Њ�ܝ6qs��+�X��[�ˌP��>�ʩ�t�E�����ګ�=r�ɻ����9k7�dr��訲��הL��Y&��Y����򧱬C9ц]LXzn�EM��3Z�x�����AMR�Í�VVx:�g�VQ*��Q�HY2V���xVF�Xb��F�^e�W�UHi�[Ӄ����Yf��Q锣���Ӎ��n�S���Wr�\[2��TN����.ב��}\YT�_�;�/\��c^dA�!^锣pH�����mf�uMs4��.��OgA�G��i�Vl���[7��r�,��[�Dе���V��ʪ�����>�6�F<�I�"jzd*��[Q�Ȗp�l�h*�Y��M�v%قM�R�0��d��C:��d��j*.f�!t�m��wEt����ü&�l����k�i�b��'#N����Pի8P�V�ɍPI���M�cz����vnm�+�씇�1�3����f��@��8nvu�Xt���_���[ �a�y^=��$������R�Q��Oʞ��-8��x{5_�ʳ�Ʃ�	HWK��(J�3u�ᝈ�w�ύe��k8����=��p�X�����N��/)��6q��T㰹�j���l�ww�ϝ�"A��;�~�v��d�z�Y���r��J�vxU��k���Fՙ�6�)��D�2N����=��KJ`��<eF@aW�bQ��T��B!��R�e���Ha���o�Շ�,{
u��3�`e��E���%��6Ӷ':o���y��Os��QY��n�e���P��$c�,3z��^,�z3Ά4N�e�A�d���;'����ޙ���2�s��Fr\9%wN
�r���8t�;�"�P�T2���������kk��Ѹ�5�M��FG=9��R�7��dyn�N
�d
SN��,�YW(�x;|+MK��R�$�$�e��\�e��K�<�V2�)l#��+i�A=^�R���/:���+<ı>�D�S�ŉ63rCԩ���퀯1aM��9�����i�e�7t49���!=W��u뷪����K�&v6b��r\����ҝ��b���:�� <���إ�3-h�I�5�w�
��9�jsߎK�������l����l���c�]�����!ЏT6�e(v_V85'4�!*��{������2gj+�����T)E|�(�[\xj�O8g[��қQh��G[�!lb�Ե&b�7��z�}�x����U��5}�����Ʊ<�s�qB���lq
b�~�Ae�v;y�';���p�7P��u��Fk�k׽L۽z)�y��9�7�T��.{�/A������٥�=�&����8S�N���i|6�nGO7�F���[a~8z�@�s9)'�
�mV��Ȋ��Dq%yh��K��:�氛��%*b��	�W�S|kƐ�QYR��"�B�Xo."�iDX�t��
�Z�xABɼ>�/�4I8�ԥ;��t�a��3E��iAP���D�!U�|a��^�/��$<��NSzj-.XiQa��-N��\Ǝ�(BA��;Nl�f�I�t�UR�V�o��`tS��{����.mϭ[[�s舜BDH�v�F�9�:_]U���{�v�z=v���=��,�����'�fK7���w��r�li5�5��3�_������G�h0����OzS�;s`��R�<�/=��֫a��r\0��Y���8 sz]t���Z:�9
v	��� ��F�
�+r��|�1���;wP���5E�t�s,�v�3P(r�P���_],'U:v�������1ao+���u��Q���W�3�~��cMvU&7���U���&:����B�`������2ꦷ]Y�`1��F���gN���z���X)�=�S��[���/�L��m��?Q��wo�֞o*��+���y���x�m��5R��;�.T����(=t/X����	�V�s73��B=<S�P��:l�=��<�\��i[��/Qw7�x"C�^���5��d"��/��X�]8��L�'Kc5��u�l�w�̻�R(�X�z�I��8v!~�~��H���HV���1@�E�!(�-�3`�����EK<1^�[5��ɘ�䕡u��|mM���x(�Z��g7QW2:�T)璪믳S5�J�W��4�߻u��M���ܹ�Á�����V;�����N��T�-�\ϢZ*�Y��s�=b���L��GSέOU��5ש༧\�q��t"i#]r���g+�*!����oc�70��qI=w�gŚ�r|����\�>] ' �Oy���n%	�e!���0����'��.G���	�o,:RZ���{W�:�+�ō3qR�\������}��Vy�Iu�4��8��bu�ڊ��N��t���X8ތ��Gjf����Dz��t�ge񹷃������&�� ����CBsF�*���3��M��:--J�M��m�lc�8{���5(��f����=^uvK%Y�7x)(�4Ru�LNGop2�S������w�Z:ޢ�r%/`ٙ��}�:*�69Iq���A��ݳ<�m���mg]��1���,�n;#r��.�¼��#\t���!uEo)���䲛�xb^��mNR1(u�g���9�����T��p���t���\5p�GmǪ#'��v5OC�WOL`jc�����TdQҁ�.��X���g@�(S�LCwND`�K���(7:z��8h���yCv1���ł��ދm�ޛFl�c���C��O|�$�������d�}b��!����N�c{\l5��{�@�Y�떊ͷ�2��<t�73���"�C�1C����O*�lF�{��b-�m��ڥ�yK2Hu�Q2�|��X�9����8����`/�� C�#29��ʞ��(M�0�������!�v�GNں�ST�0��VV:�g�VQ*�Z�5�B�9w�{i�yX]���ӭ}:�<ƨ"���D�\��&5.�γ�Z7���g���w��]G^�j������1��[S�n�H+7[��b;3�^=�`���:���̹r���̑��;p��e]d�m��+���s�4�B�ܰ��'�.ǹ����%o��92�P�s��z�W���`�g�2ٽ$�f�����*"�z�uR]Yɽ����ou���SYu��ҍ�|�a`�Sc\����̲8�J7$H�S1��ϣFQ��J���������O}f��f��f���Y%��4M]PB��-��+��\Ewf>{gM�!�P̎�/��Ʒ}�=��[K"�3f��
F��5� ��,��^@��gI���>F�S4\�l��/zpL��)@Uc��������/Y��k��w�$|9]J7�4*��aO�\]!\m\��9=<Y�{�����)��<����#��x��ϡ� ���Ȟ62���)�Y�8Y���Y��Ц9�COyӳ�~�4����E%0r�ʰ�f�]G��^\/-���;`�qw5=X.V�FGN\xƌ���!T<�֪���I�5�,<=':z���-s���d��}�E��%��|/�$c�,�S�����r0���x�
z���d���K�}\�����šڤ�(Eg7yD7V�Tѭ�V�6�M��8D�����2o̥�ՠd[՜��Xm���V��k��>ŉ��:�H�%q6������J��k��[�`[���# �zp7�!z/���r�-�tY��ԦژhL�rb���s��lV��*�_��\�É�|.ƅ)�Gp�s=SovI;�*ݔ�+	[5,�|��>#N
�:9�M�h�ƙ��flU�&�WV�P��W�;f��vj�˧f��BÖ��2�����S2PA=�����|�M��Y�C�Gg�HmK�,,��W���E��{�9LHY�X*��������[E�m�4�I��qH�Zo��8�y���eE(��T�:]X޿"��rNs�.���:�T����t;��Q�{L�r9E�kǯ���n�4�I��8��b��$��# �zYF������	]�
+՛H�s�W7\VG]n9�L�̨B%n4�G��i:����؀Q��
�w$�׳�����Qa��ȥk -��o�ؠ]Tr�#�����'�*[�v3u �ְXc��/$��Zl�,z<����sh*�u\��^�B��Yq+���&6�Z�7�ݯ¸���Jc���O��깔UaS�_)7��t�L�gL�J;5�P織T=�G0D���AKr�P����-8�-r9o���(��UO��!ξ�J���6>+�E*,�6�}��w�S���o��YQ�X�D��'�Oj]X=�iEkY`�{��0�ڂ^n��ssѾ�]�L8�D��-�u�DR��z+p���v1�_�q��&�hNVgt4ǹ��x��s�f��f�(�yy���͚,߄)$0���Q�3�e�Xۜ#�y�����]Cw�>�/�*���t������<pX�%Ә5bRK��fQ~��0����$���F�������QA]b���w)������+��ւ��ʌ��~�=l��.��X�x;�[�gְ="U�h�Q�/Gz0�3N���}�يw�1c����_�ΐ��f(�Bt��wvn��sE'g_O�:m��8�(���:U �Q�j�"��O�ud��o,mˆ��Yna��F�t�]�;5�P�um�7nx��E���)�tG:[R�'t��y�M��,wa��ǅ]n5�1V�5:�{����S�"N���k��:�y#]v���{�w���S�����.�9�Mtw�U'����/*~٩{B������_kW�W��N�\�X��V25�ie�K���Y��'!���o��E�[�+2�fR,�g� Bn�yi#�����^��74p�>W�o�+�_Z���Ұ[5�����I&:��6E��6��8V�V�cZ9u�G:���Ю����X�D�r���Q�s��2�׀\'�'�ʊ�(h��əGo�ꊹ��Z�w>Ee`wa{u��s�X��p�cn�r08�ޱ>��w כ���\2R��:�Y藅A��E�w �����er�Pw=A�ρB��B�*��\�s�<���D��[r�(�"�bS���K�|���wrq�C����x<>�8����l\`�=�tA�¶�����GKn�ݭ8nz��دc2'��1K:If��F��Yc!�z�]�ϔ�B(���;#��-�'H����.�s�֣�u<1H<�����(A���͌����f��k��˙�vΆ��}��G�ns�~��eg��\��[[F7�˧�1�=)�O@����6\]�*r=��u��#�� �D���jx�yY�o���z���N��2A6a��v��ݤs��YO�7)u��O3�'�92T��A����7*����[�U�qd�vBm�T<� �6]3�^�Tk27d��lڋ76�� ���Q�[;�ց����XLCvV�'!y�歎�oB��/_>r@���9V�V��{i�^�>@��0��c>1�a�7(��sm]�B��2oQ$bNJN���gղ��T��wꏺ�'��+ݦ�
�zMt��rr�7�d(�5T
�ؿI5�^�L�-�|��m>���ї5z�5K�,W�«��+9O�{������H׳��Դt��3����v���{�q�yɼ�Ui���w���%��T��T�pP��7�ɴ�k]��y�h��y�ﹻhʄ7�.�3�;�:�=;xp�x,]֤�6_s�g9�'�͎J����re)`���ב51Nwf6���"e��%��[�Ȭ�AV��������tx��=�a��Z��;��H�T*�ʵ�9��F�u�Z��S��#�6�	���LP����P-�zȚ�x�J�W"�R�]��av�{�F��/������}~��՝V��T%�&C�xצ_dؕr�xG�����HA��e���dpG��5:��A�Uc��iEݤ
`TeK�/�>,��������\6B�1�J��4��r�⻣PDV^�6kT��:Ù�{8Z���.��@�H�d�ŵvQ��a�e���%Bo��Y�KՃ��ol^�ݵ ��f��.�i����ۨ��닆��ק%�D0��K���(2�u)�'oZ7W�.��U�������v�H�!Okw(���c�˫��g)�Q�_DEX��6�Y�`1��ypv�h�ܫ[����=��oe��
c�'�����ɗ%��r�=�H���,5��Jʹ٠�����Y[�5����5(������tX�m��5[�i�����r�����j�z�p�C��ң3��g�����]���/-ي�X|�r���Bj����v�B�ݩ��:
��%d��m�w�}(w��um��=�z���M�ڼ�5Nf��ma�m_u���;#��۝)#IS���� :�Е qV;�����J�oR��v*��d%b�Ơ�9�𱖹[��Q�-���B���K�[�Vi%*�Ĵ��C������M��\�rg;�]�yր[���6�����ĂN��m���}�*�ᔵ���e��\�N���K���V*�44J�]�e����h��,���-@�A:���uk�
��杁"K�T��-7J�չ�@h���z]㘂�Ì��������Fʿ���%1e����7�ֱe�drS���%G���u_m5��'��&͎��7�>Ǉ;W|j'�	.�x`;���1�ASܲq���-C��(�#D�w�*���}Z��^DˣN+u5�6&�: �����χ�$���c��x���>�[���5w@2�u���s�@������eș�UvU��@7 ���er�
z�$a3�N�a���O*	Ӂg��i��1���71��T�s{{��r���ʊ�x��eΓ6�|�� ;;6�r���r�w(�Ə=������uˈ=���&*�9`�Cx�]�1��L����bd���<2��qXnRBm��h�ij��k�nc���m���ns�O.�+���5x�7S�45ۊ6��g75e֚�Ƕ	z��ct�� ���*���un�'V��Ah�;y`���:�QQR;�Í^�b�}xf�%��A��@n�P�ܘ�%��݅�Ʈ����^"^� � ���$�!�4.�|�ե��^�����Ќ�U����S�e$u�Ѿ���2k�:��8d�J�5b�ڻ�P\wz�t���sUg( :�1��sW/�n`U$Kp�d�+Q��q��꾇�-���wϱ��sGv��S�x1#+��Kx�7��S 6u	V@C�7�ĭ��q�Oj�\�S)Sz���_]�//u�MO��0+b��c/r�3֟X��T�]oR�#,���ov��:��mu�s��	^�n�&oGܱ�}�+�.i�˥�G�bļ�6V�j���_-���05Q��T��U*�\8Ġ���(��X#UTlEc"�Y�b�d`""�f1A`����
(�F1m+��8�\Xc��	TAp±AQQ@F",AUA`�P��b��(�aD�+ZX�R*�[++f-�*1f�[�X�l(�
��b�e�A��1dR�Q"��b���Ra�qC�J�*��-�kT��KJ����
�+"�
�KeJ�
ˆ���P��U%1J��ѩPb������
��G3�+�1E�,U��%Gb����+��j�5�J��<A1��@ �S�c&z�U�;���rn��J"3��$�*�[.�*t�3��	�rS��]�l�c90b�vj�wQX�>Zl�f>�G/�*u���ҦVx�&_�r�f�d��	��KdZ|��Ocjb��C�`{v��7���G'��;Y�8ul>�s��L��5Q'�����<�s�uR�����T�q�Q�q��gLGT�K)�;���7�k�yM�躳�/{X�Z�������g�jqd�3x��P��lzJ+oԛ5Y�:zV�3�ô_u�[�m��۰�ԧI���!�䳶��:&�>.�"Ĩ����r��\�)+幧wt�=<��Nf�w���ܡ���Ńg�V��8��ĸ�*bm��KsyŽ���wa�z�;{������W�Sa��p��M���پ������`}��j;|瞡˷փ�����|_� 绮>�{O��E�_gy�^�9�ۛ����o���E<T|��ě���ƾ�r�3c�eB�ŕ}܌(���el��07�Y�����ƵqԬc�*�-�mT좾P��v^�JՌ�A�R�mc����q]\nF-�S��5�x�� �������.�4�i�j����[��Pӆ�����z�q��W��@�ૢ.�5I's�G\����j�fM�j�x�S
�o��d.׷��Wwr�[�߭Q�<(�ߠ+��"�����9Y<Ů�4kjw�B��\��뗛V%>�o�De!�@��,
�Rnde��rd�,�GD���u��e�KU؄��*^Jɚ�t�Ű�U�������/X��\ݡ�Ǻ�hʑ�%
%�
�������Q�)�����^?R���s��o"'؜��B��=���_-���f��:�0ސ��7�}W�7jgD�y��ͻv�F�kb�'��m�V'2[��r�1w��g~캝�6�ǆ�:j�\����U����u�Y0s]]MK�K������l=��KM �͢�eU"��h�t�y�ݺ��~D�ONy=�r�r��������y�3��;�L�R�d�Vb�/&2�������[K�A�;y���R�쥥����sp��e["�4�q��6)�w�W~rbR�!! �_m�κ�vQ��ɲj��6���9�� ��3/F��ד��H�\1T�zލo9I�;"��{�ӧ��ю�6>��f�$�:�����j�~\����{�a��}}�zxJc�_o�*h䰺S��1�41zV�{�7�F�����V��X꼌��Y��jG�,�&{�!r�{�[Ɔ>��ק��qJsŮ�)|�~��{��rq�s[�z/J��s+lM�\g��e�SO-�T����v�
��<n�U0������A�tQ�[�O^K��!���;���'o�e������5�3��s�u=��o��c;��W�� ��"�x�+�9q�k�t�wKW2oY�؞��T�S���vڑn��R㦄4��ڬp��Ao2W+�����W>���U�R��Cv��۷��b�Lh�̞�XZ}�z�q)e_���ى�s|��Z!p�t���Пjz&���S���E���\�Q��(�T}o	�.�uPo|æ���$KdKi�l��w�&ڻ�K�۞+�/e��g�Q���m?`��EZ�:=5�B�e�-P�CF�O�t�DV�Q�U��󨫒���d:��9���v�%��m4t����˝���:�uL.۔�<j��#����Ϝ$�:���Z���i����3���^�'3<����nT7�D��=�R��d�k{�n�3wm�]a�W¼�Zh$r@n�POO���\�ˋ��*���w@i���[���޻7��X�:xt��{{5��4/h�ׂrJ�wcLFX|wo>�:��u�፻�F1w��*x����켉V&`�4�Eќש����1�WY,`�
�sT;R4�>�
�]؉Q�e[�}�`6���1������3�S�W�5'ѭ
���\������9�UO(L�r�NN�9f���g�ҽ�Ɩ:���DN�^�H��y6��W�jط�w3R����"F����󭷻j�PQJ13�6�us&jsoT��qV&����M�#�*����<��tR�,t%���F,�U	T�6:�'y��36��Jq {������uw-��K{r1`8-v#E&��U�q[��S�����"�fOJ��1J�C|�!�4�0�̻l��F�s5�79���rRr확���ǫ�K���̸[�J�SQ��7>g��[f��ŝM�J�MHufkojB�X�
=:1:�15��{�T7-lT9��t�X.wfo,r������Tj���Vj��\כ޻l.\�	w/vz8<�S�Q�9=�!��v�kl
���V�õ��n7AV����ޢ�7��e�%κ%��U�ȚL�2�/вi�5�'͸���;::y�93����������)�z	�&C�xצ_d���2�֔�M�p�Q��9j����EH�$��*�~*ɗî��ٹX�i����S���z���u��p�\,o�n���۰��]�wsf4�u���n����𜹪J��UL����Jޛ�Gd=��iɺ!@�x��%N��z��ڂ�F�EV���ޣIz}�Ejf���.6��1Zv�C]�,�՞�X�U�)<�V�ҷ�f}�a�9y4""��>����I�RX�����v߃�����.TN�
�o�*��+����@��^]zk����<�ޣ���z��;��u���[ӧ{�o}�i�ʽ�������.<v�d�hi�W��ƫ�++5��;l��shrcV1��!J21*nV��I^����]Nþ�q��Uua�� [:�5ذc�ˎ���U��\	=ܜ����;�[�;ܡ���Ńg�V��ga-,8<�ɱuϹ�����N�՜�f0��ܩF6:t]��ׯ����P�N^���Q�an?M�њ�Ư���G�U��m��ëf�����Cʐ�:$h�Ҥ�uI�fs8r_K�M�3|���/k�k�fvxn��S1���!Z�_Pz���w3BٓG����x��*��NAr�}�3T}=��UOO��,��"ZG� [[~��}\�V��f�e�s�S�oj[\��gg9U�O��������
�2���������ˑ8�'{b��%��Y�����G�L����T�4��ub�+�~zzi�ŏg*{��^	-�T��&�V+�z���9w��8l
��~�����;"'�3Ðz(�#����3��/�(=�>�ɝv�@�.�}�#,�s�p����.�7oLY�ʮ�=M>Z���7ksj��m��d�I�f�c�V�BT�f��k�;% wo�ܻx-�=��sZ�2�_3@�c@4�Z%���5�r�iٛ	Wh�T�-\���e~<:��_f��Y5v�Zq�b;[9j'$^�7��5q%��;�f�Î�xl�:��j�Җ���١ӯ��3W��]���v if�T���K��J��43kŌ¤��'�mc1�6V�ޞ����yL~8[F��{��j�C�ؚ�C�6dSc�*5��=��c�J{�Fk�ast�>�W���=���r�a�F���|����s��Ů��s������N��oO����n�%^q��騨�O�(���q���������[���^;�6�u����s�.1j�P�]?�ה��=����̭�7�K����Ħ���������Gg;��=��ux��?R�ݴd�͎�'�w|vP02iyU7F��+��c͹�U*{����c;�޾���h��bS��3�w(�#k��j�r.W�{�������V����=��v��_��Y��ƺ���'A�.a���Γf\�R��h�����{7a-N̲Ku�*�5m����2�g�i��5�nP�P������c�=ب<��]�ܬhZ�P듒���5��R��3�RW�������'>�ԧS�����/���O�`ۇ��&ZJ���w~�m]�P%�+�v���%��u���6?��S�����o�1~���u�*�d�0'MȾx��}Θ��,������νo��c�k}��/vU��Y�l��v�uz�]0�]l΋�呼���+��TK�î����+�UZ�^c�2��QԢ�`�X�_lC�ٍ
�My#���y�6���)=yr��������̷1�=���{s�~�OD��b�����4v^��5�+��3^[��~	�ݲsr�w���ˢv��5z��{���Z���h�f��Abwf�V*Ol95��>�Q-q�Ef��]���ƅP5�P�Hז'�M��3n��D�s�.+���3j�S��L:���i���g)��k��ٿ1��ȿC������s�������bU�	�����V�e������F�V��	��] ^�v�#��v�.� )��̙c�I\-����B:�m���t^�r�|o���>����nm˥P��"�^�D�f-�N�\Q�}�%9-��Zyt��������ҽ�k�<uP �8��z�"��HX����}��ֽY�ü�<�cw���SKG�R����3�`M��\��q@�8o3	���HE����#�*<��؃νy�ݺQJ�:�e��+Ț�鉵��Tf5���}�H�I=��c��5���pә�u������w��\����:�<������Ju�y���)�T�6v�C�ټ��;���r=E��*�⦵�x�eP��k��)X,�ڗ�n�7�ٛ�Λ�X��)3�!u�e2�է'؞i혬;�w&uE��'�R�cj��K}P�{�	���O�+�֥���,���f0�Z�o�'C^m���
IiS(*%��p�&�L`+��U\���f�8n�T���M����=�hr44q���*ͽ};:���3]�*"�H.���9~F`d�B�����SY��7Q���Vo�"��@��|�Q���:�_���[�S���D��y����ao;��f�w]���͎蘅��!��u��ɚ�\��V��*ğY���&��-
@,�o4_v:{����Juw4��@��lRV���-�F;nv�<[����~��CV޿[����G4a��>[�j���}�1E�4�K]��Os�FwI��6�#{R��e{���̋c�>s��I���{�D>�^n�Ws�8ƾF�=�k5���gD����J�k�Bb"H����{��^~᧼ޞsk��|�e��w���Z:x�-��8�t�J�9[�Z�u�W��O>��S��zy���Nӕ;x(��y�3��0�+^b�Z;����������<�Q��~�u��������>w��.s��C|��}��f������=Ȯ��/o�ә~��.JBG_��E�k�:N�(�Y������}{}<M.�_=�]�C:��u�򅬒��.�uX[�^�3hb�%.��:�V�x_w��$ I?�B�� IG�$ IB���$ I?XB����$��	!I��IO�H@��B���@�$��$ I1H@�z@�$��	!I�$ I?@$�	'�H@�~�$�	'�$ I=�$ I?��
�2��L�W6�����9�>�B��礠%*J��J��*� UT�*T�Q%PQP�UR�)Q*(��P��RJ��%RB*�)J$�T�P���>�$Q��Z�`��jl�2�1Z0�VƨU*��e��EH��fb@�)5���խj�[j4!EE���l""�F�UV��nc�T�VX�H[m�4�)D��M*J٢*2b6�Z�T�f���P�4JHQ$URZ2��F�.�Ju��R�Ҫ�������f�W�  ���N�cj��,�G�T�t7mcB��n��l������(�F���l�V�9�u@
��j�6]p�4��Ui�Z]�Sm����   �x�Qm�Z�j��h�;�;U���:�*����V������%c������S6m*��P�Gp�@(P�С��
�2�M�#L+YTAM�   �����
(P����B�
 �@�w 

(��\� СB����
(hh�
z��
  (=��3E
P�ee)����V (f�r����]jPֆ�IF�ͬ�7^   � 4-��**E��� J;��H���mc�kVճ��24�%A�`$��4h�MF�Q�l�檶�KMD�km�ڶ�U�   ǀ��	�4$j ��kZ�5UM��ԁi�[��Av���-f����(f��РZu��
4��Dif&��.��h�fUx  �� ��	�\ 4-Rh���ST�66���UZGwB��UY��-��6N��(A�dX Ыt�TdPBT�[Ex  G�P�y��@�E�N  v.��. 
+g\ k]ZS4T�P��ۘ�@5;j���Zl�(�-j��v�� <(���o[n �Ɣ @C��� ��0� �ˁA*�p �� 4u����06R�m�ji�  ��
P]ۊ 9���c�

���Xs� �� �.ut
����E��m�Ӡ� 6$�����[3@h���T��  ^iW��`�����jf���R�i'st�SB�a� @YJ�(*Wp�5�J�cu\t4���k�����lMKZ�@h� jcA�%)   E<`���   �{)�ʩT�� �S�A)Q   ��M�i�@  �I6UI  KB�F���U5II������j� � |�A�]�J0�0/��*��jT'�{��I7��BH@�h�		�!$ I?����$�d$�	"		���/�����K�@(���
��)#�Cx0�WI�;�V�6qD��dI#j��nm�MT%CK1���C��C/d�RdC�ٱT/4�,�6�2^�N��3�/�%-;,n�&V�X�++)]Z�K+TM2�dQ���_ƈ�,�"�Y`��-юmh���cB�Z��*�(�[��,�'�flZ�^X{��H�.�4*M;i@hPYK`g��얞�A�mh���'�uh�ouV	�iz��2�cv���"*+2��}(���1��1��a4B�e�%�X�y�έx�j#����x�;Pk9�4�q�&鸲�z�
mU���56��nU� �*��J[���P謈Nj�o,d2�6��,�� �,5d�� ,�J�7r�Ʀei8c����
Ձ�k���:��vT����m0�\��Z��\����m"퍧)`v7����ߵVO�q�ˤ�šp��ӿ6McɿC�
z(�B�LL3W�!NL���@2�q�F�J��`�Ð Y%(��5��r���KV$�.�j(�(�$�)^S5��gǑX�x^�����Z��^R6�jd氶��,G �Ԃɲ�ٔ�rk9Vժ�NΌYxq@p���x�@2,��[ Uilb̼h*ʺ��R�
��z�Y{tlP�DD0SŌ��I|�z��,��Y��
��ӂ��ł\/n�V^R|_��
��a���rջ�z�G	F�&Y�]*v�̖�hmS�m��j*ࣗ��-�]��Z� �T0���	��ӊ �l#JDtJu��#/^'M<��+л�\Ґ�'I��4��"tR��H���[vCA�,wr����6��Q�/.�
�^��$5�9B�U�vU��e4�Ϋr��=P2˙�c� �{%eӶ�I-<0�TPih$���.F.�W�����6]�5�hXV��i��xa˩[j���A\�e�e�8�ѕ�D��@����K�b�)Ah؋R)�)������{Zh&Q�u�fʲ+0R�	�l'Z�4J�i���c7�b$*۫�ڕ�n*%��@{�
�YF�]��&�il�Lj�+%��c����Q�Ul^j�+%����\���&�6)�F����"a�lǙw���M.��XIE3n5F�e�����AmZ�@[�+Zh�hָ`rس�or�Zn�6�F�:Wf�YH��n����� �bj�(���d��z(k����(Q�Jܙţ��В1�����n�֕�@��aa���n,�o(h4�IVnD���p���T��[_�iim!�Y��P�(�$��j)H*��I+���׸�?��wvJ�4f5�a�K���)�T^���2��L8����-�0�� ���&(+hd�q�A^�i�c{Roۓ]k�X�$K�.c͖h&��@rVm�M˭�+��!SN���h6�,��=�<Չ�C5c�W�F�qm�^b�m��I��ʹ��vYXVˬ ɒެ�jP�L��x/D�ԙn�&��JWcVP�	@��٥ Y7AĬ
��� �:4�P����ճQ��A܂����3AM[B��1�E�	i��2�X��T̐U�=Rl8Zi�l+`�Vnm�[b�e���i�5�t���Kn�TFړ$Z	n� '���P8�KW
m�,�7m��ڸ��ʆ�����2���[Ӯģwe-�"T&Bu%�=�&:��һ�A���6�7Yj�vL�ɡܖ�Dښ@����k����P�̕��~���ج
 �N��%浔�OsV��?�c�r�����)�)�XR�{{+D7E�I�leձ����o�`XR�,�8�:��O	���2�_c��-��솞�r���h����ң�հ
�U�d$\�L�XX�Y[q82Sh e���x����fÚ���A�
�F��e�,���4Ԡpl)\���]Mr��/5S�W�O�`)t��ݵ���܄9I��25V�N7"Z�M��%�V�e;�"�X\�R�4�-+S%G��x����tf�\�X2�j��0;ڕy8�1Ysvy�FQ�M�;�j ?<R���ۘ�LR�ӧQ 0/-P17���&%����i�"�nU����F�kޫ;�0��0���eJ�Ā��l�([Z�k0�x�Í�w<Xj�;�e�
�ۯBJ���1$�ci�����b���N���tt�H2[g^��(V4�Z�Y0���T�w�@^7�Jnޡ�L4@uu.�;,UӥZ��*�r�S*�1nU�Ɵ�Q�]��n;'f]L�V�U��2��UV)�MөE���
�NPw�HM!׺�
�݌^�a�WJ�u���UwD�ZuP��A�!�m$�6�b�72����[�ØΣI�,V�T�`Vt���������l
�G".ҷ��d��zZ�3v���&�MY'- ����N��[�LT	��:��|����w�[��V6� p�/sv�:p�m�^��=��I�)�k\Cİ�F�T|m+$=�[ȉ����Z�7�qf��fބ12eJy�44�*�*�@bI�Q[A=TS���Z�^SƄ����CL��jܷ��R��/�(�Pя`�l=��9sW�V���^+!V��5� x�!����jR�w ����&E&) ����ى����u�z���([RQK��*{hyX��*���2� ���m���ʴ6��;z`U�,ue$0h��ǎ  �h9x��+u��z�b�~�s宜ո���n���qd�����^m�4�i9�4��� ��d�*b���4uC�h���ر����B�]j�$�:�8���aF�鬰�f�6+S�*,�v�y��Z$KJ�j�8*�4�&��-�#҆۾�z
�B2zS����4��J;�A��Wtn=�(���,�L�`U���PV��)B�"��[N�[��
M���X�m��kpa��0�L�Y��a�-V��,-��J�96�E跠1�q<�
�Y���zR���wUA��	(]��� �Z�ť>�������n!2�>�ȁ����}b0��¤�O��Dl�G��r��N�d-���hQ�NT�V*LL�ߥ�+�]���r+�:��d����`�k�IYu��n�^7�b��Df'��ݢ�u&�l"��Ve�i�g2�����u��̫�:W*��1i�h�E���]�0�N�Y��q���U��KmX�Ǧ���W��)֝�@m@�0�iL�i�i��F�1xxF˦/^�9<�ax6�֫DS�G6��Z��iL�`:�GTj�lI�i#��ݶZ�)����eJ�6���rm	�K��b��� 6ou:Ȋ�FQ�b�#�/^�0FT�YP�mޠkt4��2%è�̠����t������K���Y�؏f�Q��8¥��4��$|�ddǛ��۲�ù���ˍ�m)0��֍�o+N*%��>A6ѬaA�)ӣ{LI!#V�T4�� �ɏE%��;��5�2:0�74���C@f��4�ÃV��C
�b�7YdK��p�۬d�h�����)�`f��&� �(AbRش��衶fݚМ���ӧL�G.�Ӥѽ�W�)Xԅ�����_���/�A���^����)��: �w�rR��b�v����v�eҺ@��Q�)F@s.��zj����ͭ�£���
�<�J7�F���U��Ȍ�.������ʈ^BL�ދ��-zw��l�R�M�kw��ȳ`W��Xe���
�F��a��oq^�`�v�K1�"�2E-	�;Y[�+-��g4��DZ͏2�қo�hIY�X��j��QY��X���-4�7��曘��P\
*Z�(m���Vk�!JZ�kl3�E&�RR�q.'R�A �a� :ݲ񺽃e̩�E�n��  Ԭ��z�b� �.VS#Mb4vU�Jf�3�O��U��h�W��m0�.菄l邅N퀱��զ�h��2�����B�4{l\�]��f�9Hbb��>0��۵Sǉ�e��ܼ�`ղ�L�W`�r$�^��*��쥙��oK"4f�FB�m#{V����st�G�^��.�cz\���R�P��}R��&�r��fm\��(f00%�p�m�� U�ɝ���Z�ф�Իb�/@Ť�6)���rma�B[Z��eí�5��
��w-#��m������޼���m�/���z�%��k��������K�P[4�J����{t�Vݣz��.�:
ō�	l���Z&�K�܆�mؘ�,�h�v�D���v��
n�t������xad #�/EH"S)�c.ZyNP�輚fC"u�)V�cQb�WF�A�(�Guɧu4��
�Y(J��V��p�Y��B�@��:&�,lm�o
�p�����)]�ɶ���jESGF#P�!�`�	�e��X��^3b&�ww����F�l�mڭF��7b�k��S+)����a�hT�*�ܹJ��ٟZhT��5���᫴��ѡd�/p�Ñe��íC"wEM3m!nL0�ycNܵb��sP
�rc�p���oo9�[�{��bM��IIJd�B�L���VL�8K�"1��u�ͳwVl+�f�ۢr\:,�t֗*|$�9��D���j, /E�����ـM
��H�hH�wN�@L0]��.��Uڦ�7�������R_�x��F0��Kr�u�Һ9��y�*ͺYx&jв�����U�(7J�[h����GB%�]Y�XD�D�5*DGN� �� ��ȥ,���̖�nm�cM��Y�SR�+Y��@2��54���BdN��y�&Q�b$����Uwx^�֙�\{�,C���b����kF�L���PY�{-�F�nRZ��i:q=��>ȑ:awz$�q�[>ٔ5T:nV2�8��1��h"�!MI*?V���pʴ6m�YSVFl��U-U�N��7y�Uޚq&2�F�`��nȉ9kC7p1�c�+���im��c�)*ݧY��l��2��꣬ދ�����	P��q�/��z 
UԦrD	��C,�BH�7"	7.�F�
l���J�,���V� �j�j����v���p��滬'U�9HE�EQ;twK�13^���B�!(>,[Y�Y�RqôFQ�2+ZR�o@Xl��д̩�:�p(�ȷZ����`����܋i������X$����F��Zw1�ߙ�U,E���@�X�k�ܘ0Gq)�W"Y6Щ�L�	�o\A�Q�ڼ����%��v�a��Z�ǳ^GZX̔4�j�A2��]����sj�VkXʩP�e����ZE�2���kV�:�\�6v�X�kL�Ahe.�t0<�d�uz�{ЅK� Gj"Nj�c�N���)���rS�,ݧ2�Yd��n��
��wm	�֬.Q��n�@m��z���`�	�JP�n��z�Zkͤ��V>MXI���ƳZ2��f�䬚�a�T&��H�kn�գC%Ȧ�� �L�p�Vr�bf Kd�����Y���z�(t�����M���N&j��̏w,�[�d�ջN��Xy�&��1��WZ~���LZ�Akˈ1��ɩ*a��g6��g+)�j9jۚ^��e�oE�N�8r�l�f���a�{0��	�,Ԃ��i�� ��,��v�$��HD�>>�1j��WIa� ����c3�dî�¦�T����P t�H]G5���KE^MJb4� v�N�,��[@�0۱,)w����v�N��zEX����n順+��ZX�XԢu�:����ʲ�V�c:���v��4��Vj�[w��f�ƨ�wI�6�U̬��f�@�a��ąm��ȳ1�B;dʵNY'n��m5�Xpl0�x��[aUހM���K�)۳�c�Km,�LĩvEj�M��Y���hѡem�JM�BQ�x��L��;�YB��\���!�)�ht�����"�Q��<�&V���6]ihC��Um��+^��2�QeD��V���5�f��VY�o(�Ř�wj�3
��L���g�x-Ԉ��eH3aSn�kJw��
�Z����ץ1zY�Q�v�a�J�d6	��uc^��)R��h�eMY���Կ�zA�{Mf�/1]�HԈ�Hݔ��S#@轖���fLI�mn �;�5�܍�%:�MkH�x��w��z))����ĽŌ�� �M]\�[kL��ړ2���, %�@ܡ&��̢u-��BfTX*�f����9���Ys,(�n$Jh�oD����a���s*�Jٕ�-H�l�6t�I,��W���'d�T�C*Gj�V�>���#�ʠ�ve���v�7D���[8���j��.�R[�x�Sad�;��VL�`��X�a�R� ��4�檻����ch��Z�Ȟ�n�]Ù�i�mLtn��(	�mZ̛j��6�I�D�Y-<Kqf�5�TX�u����(4`�r��yb)������h�Өhն�5�u�j&J�ɅX��Pa�����1R<"Y�c��,\�L��e�
(`R�������H����1'5�����+k!��Y�a�F��%1�	(ǲ�OEUX.H�ý&��Ot��`m �ݻD&߅%P�faq��wj,�R{V�Q��2�W�%���R�f� �\4�QM)-2Ӓ��`��	��XK��Kt�-:���[�71x��Tc����`��Q��q��D���k�)b�b���P�&��z0��	� J���Jcni;B�>.�*Q7�Wʃ7�+Sn��+p(a`I%�[�����e�k���̱(�D�g�v�Nݐ�F�׺+�$�;%��g�'�y<u�P����ޡk�]w�
⹣��>����X���)rV���6�#�5r��s��N��v�c�}�OT�4�ͳ�X�q0ռs Z�����2�r�.�����x������&�j�&$��2&�uoR�آ{������`ڔ��yF�0���8sG7�*�dLBj�ɠ>�ׄN�5���v�+zJ�)�2Qg�u8�T��R�!uě�AYܗ�(Yu�Y�fU��ړ�h	@���oz)�%H��r�ǒʾ�c �YX���:�e�)8�nR��}����l�^�g!�([�o �9�Js٣&m���ݡu�Pm���\��^}��d�Gd���a1�&.Hvdn���ꮵ �Θӭ2Z{��,J�M�s�Awp�y�y�[۝Nt�Y�p*��Q�`���;6�G�,���:Ԫe��̷�;�|�Ю��,e'9٣	��&J@?C3�W���g�����$��.�y&�Oo�Exz��Iܗ[��#�H�U�9v�o�}�:�#X�w�d�oh�U��QB���*1Y�%�U���C!_U����֮�6���f��1�)
����N��H`S.릥:��ͯ�kާ�8`��C�F*��FTj0��	iSÄ����G�=9�z4 ��#v�6�����S�R�(�o�.�8����#�X�5�N��WWۨ@����7f��L�|���ܗ�r�Mݑu��|�D2�E"�kB�î�1�Õ5�X껔
��5T�e.�&�=��)6W�@K�2��Ч�@�o>�xv�&(( k0.j��˧�����7���.-�9�\s�.�PĻ/Fcۂ�p�x�#��m�y7:F �H�c����p t��pX���V��SD�{�Ⱥb���2�ۻ�{����#��Z��Cu|��ٳ�٣-ø�8�3����v�SΧ�3��&�<�q��]����<徾`rf��fO><5�j˸�,��(]!�g��3m�N:,�X��_WV�"u�����!yHWNyR���t*p�ћm'I�[d�����F.	�6;����Y��$P���E��$���l�Zu�9[m���а����lͽ� 
��!ک�U�۱�`lev;�J�p�c ��:>�%C�V�.�5��٭дΐMb�^W��+ViheLzqD+!;1gU�V#�u���#������f��\�,�p\�����qK]W�o�VN�+��诞�{�G���ؔ���Pl���1��S��;7��3F҇����Ň]\�u���9�n�
#11clk��^�F��c����XW\qu�tt����<(;"���H݌#��N�7kt�n�n�z�\ҫ(]i���wSkƯyl�;n��uM��=N��_Zn�O}���q������e@�k�x��X�����Juδ�[��(�+-�E�Oo4��Ws��9�3E4�v�Ct�O�t�*��Q��;��+ƪ�R������m�ni*ST{2�'Qk2��%�C-*�����[������0	ǗI-Sf5Q^H+�7�r�G��qdf��I�w�p�&�+���֚�1�X<����]�y�4uO9(fy�H�%n�.����p���T3q���b$�X�*��+87�V-Ҝ%;C�m약�$����`o�7�_8xd��]�_h\6��7�u���Z�(Ȅ��^;ƨ�]�:u�b���0&M
9�+����#���(MO�0oc�c���Wy*�ᇉ�0�LK5�vq�9�v^Ы��N�BA�)^+�ڒ�=�T�F.s1#[\k/�r# e�Ļ��;v.��>YH�F����Ň��*a�+n���u����Y.wA�}�}�����x��O	�`�/�^>˛w��"'h5�E3[��9bӜI�x�]��C�v�)�������cw7��&S�s�z&�5'�q#��ӏ;f1a鼤O17M�;o��l]�::�.}�
��c����[
IU�x����i�Xŗ����>"���A�n���t���fN�)�&���"�թ��|+_J
ޭ�
���p��m�%e��pF�w:�3`��إ�T�Zf���3q�.������:��T�[Ah��-��<	�� ���5�L�Pv�ݑ�w�n �d�7 ��t.���vS*����g���t�F뚷4�
s\�����!���NE���-�\��=X�E��[b�gt��՘틭��N���8��;�W:ڳ�aS�i��Q�%�}u�n���P��c�J�&ާˈY�|�;�s������6�S&�����]�f�9k3΢�
M�X�/�aW�y֏H���+����W/���h��Ӎv6�=S�-Wn�]:J���Gy�]lWӛ9\��J8+Q�\�+������Z� v�[��$�u���iV�!�Mu"rM����E'�u]��uC�&�RŮ����c�9�=8ו}R��7av�Weq�����a��ӋF�vq#{ ���2�K0��A��oW;y��� c'�Z*����h �i_p�9:0k�CT�J�ӽ�4M�����P^
mo[ݸ"m&��(Ib�v,�5G�n�}�<����'���n��yxg�#��q�I�zt�]�k�����5o��:6�w��].��m��u-��E�C`b���:�l�2����\�����X]��7h���^��t,�U�ttE�&*C@��c�ʬ�P��,�}�d����)H�B�r�7e �e��]G��wQ&���i�!N�06�<R�U��t�r(�mv�b��Ng<7c��Y�Uu|ШkU�Y,��۞�{��3QK�Gҍj=T��#κz.���<6���u��7"���x�1���̢y��ݼ�1oxM��3b�0�F��|�v���C&�n�/�r�Sf^�l*�a�WPGz�s&�3��<���-u^B�g1�Pe�ܝ���+����Ǵn�)�f��kUKE�46�7�:4��Iew�1@�!��
˩Z�u�4�3#86��9���s��_A���ys�؈�t���K��h�|��7��C�:���{�|���џu�H��9y/��M�P��iXϕ�������S�U��VN]چj(�Ar�5�ΰ�bP�깫�gmee>�OU�u�Ќ9PS�j'qY�H2.�2�v��!���ks�R<�ʅgu�Z��v��0#,\L9H̩��!*b��|m�P�;m�c��S,�w��Z6=���(騻J��q�1J��i�n����罓�W��9E4b�]�4�ܱ��|�z�����]�d�K�,�2v��iGti���:�^9wy�sf�m̧��so���t(-GF~Z�[N�k|I[sn��&M�"9�h�02�1v���Uޭ�T9uZ���
�N���������ϬK�}�Jۯ!�q����\Y���QhʏU��t.�A|�7�4�s�	�}/���~�"T|;���/Q�x�L����y��H��`�|�u�V���f�ZWq.���u!Q���O^��p�j���+n�0�pF^�̰r1�w `�����Zd������3�K����=�x.��Tei����{�S)��t��R�<���z ��:\>H��\���2�8S��M���찷*����/-��:-�l|�h����*loU��^͘u��X���)Lf휩G��QVlWL�o_b�o�v�z7��7���j�Z��^Z�Z���ô$�<��7�-c���C)���i�Wu(���h��f��
��Z9t�^�>k{��+5��V�9F�YƆ�R�(�q�%*��;�����(�cu�����sK�����#Yp�G��S�<�+�))Rg,�
d��^^nB�	�@o<Ok��F��XΗw��rmپf�	��Vx� ����C�wk�z��ٺMD�`�Quu��XA.6n�� �-���yк/�s<]u�Tb.�ν��eəZrr�*Qԑ�q�v�#5�H�EϞ�I+F �jU�kh�$G�1#�I+F��=�E^oU��lQ� ��l�t�L�-r�=c5�46��v	V"r'���T��)�q�wx��FƱ ��� w]��S�R9�'�i�6�.�&C��>�����fN�_ʪR�&>��n�U�U�7��Bop�ĩi-2�Һx]ϕ5\d�R�W"}O^�hN�P8�̷Wp��YJ��H$�rݩHQ���٦�� =�|�!�u�!��mnt5/1_�E���Zi��q�M$>E}�1�,W��G� s8GKh|cޗ�+�N�Y|	�47n���m���G�Ǎ*��u(��DeL]Ưo)D�-���XW%�l�E��<rYy,T����^��U�5i�C�֜�-�8u��͓�i����$�Mf*�eŹ|�m�E��@x�1NC�*K�[�������j�CsB���zַJ���s�N�խ��WZ;e���Ֆ9��+oL#���,N�B���pl�Ьr������Ch���q�6E�C\�PX��-C����
�o�Y���0U
����P���qن��PaU�0 �w����]��&��'+��P�XJ ��@���xje��{0���*������w�rG�7wo������Y4�F�A�;Ė�+rJ3c�J�j��������N�����er9�\4���٦�p��f�I��[�ͭ�Т�$_F��B��1�չ-tT�^ �uڰb�6���H��m)�*�����r��J���	:������Gh�}����G���Gu� 8<���Wv�}�WK�q�Һ$���;� D�,��a�͊���us�����p�}�֎��N�Cs[f�}��1ӝ���z��傢 Zrti>|�
��FcYW����^��	G��T�o[\��pZ'셵R��鋇�e��b�A��z��.�;�-�/�?�߯r��i՚ͮ/�$b+�9l](��43:��=��Il����sv�Y�d���w��DV�q�r���3��ʹW;w	�Q%b��Eu��z�Rzp�xt�%b38f�}�	63�3`'�G�j��K-����7Q�"�V:.�.����{���pq��3w��؎���e�D_���F��)�MF�{|B7@�02o%��d��qa��p�ٌ5�,H��e������Y�7��c�(X�)������kü/��c-qۑ�S�;6�&��H)��' k*�for�cU7�	r)]��N3G��Ӷ���v��˽)�j}�e�X�\ԫ�g	�ڭ��	�ކ������l:+�����%H�l	�7�ò��Z��_u�'WV��mK��D ��+s ޸�}ГX�k뵴�1Wo�f��!^�xJ�A� �B���k�մS�ƴ>��E�~�yA�\� Ɨ�F�O��J�M4���o����o��<�����S�z�ÊӧFc�hKb�)�ֈ���{:l]ζ�@>�W����{I5�K�<�`ݻ�c�OHM�}/c�;:쵐��A=kEè{FЖg����G�5s����Eh>n��q��b���ا1M������3J�k+�M4r�=�&�ވ����z,%�p���k)f�ή�]�{{t�������5�=舵�|�Fvfr��[K]�61V���9�ڒ���G\�b�ň ���	�����}�����W8���̈́F���nQ�/�f
���T��[WY*(]rPi�1�(��&2+x����R6R��m�I��h�K�k9���2���_՝� S��&���pi<����g]���f�k뾦���K��HT��Y8p���0����� ��%���U2�ت�x��(�t��[oQ,$`o2m��N-o4F���^�ZOL���VC�F,<�&L��r�ÄT�d�Z�61��B+���z���C�`}�<�JiF��i�ʾ�G�85=C��1K<RAr�c��`�������d#Q��#ۥ�+OZ}F�ź+/k�v"vՈ*��('�1�E)�e�a H���2���Y�ju&Z����H�Ae��r�A��\�d�f�f��ؔFLF���n�t�+DtT�ʷ��s����s��V�f�]Zm��dAuܬ�q�u.�Ԣp�q�Ws�%
톙V��9e��Ԧ�sz��\�g��=6��D�8�u4<樫Ĵ�qD�m�5n�Y�z�GE�3��`�Ӊ<&gQ�/T��RBm+��]S����bn�JIX�
m�U�[/�7�=})b�Y��뚠�Ms�2̚�\7��G&����$3�ͱ��һun�wo�ە�;z��a����S��k;"̽�m�V�
��c1�+��G:ܹ�}��f\w�Z�-�.P��h�;t��Ѫ��Z}L��~URk�I�_���we<[�u��v���+u���z��N��"��՝G��3�5���(�������f��T��ݡ1]��[aШ��٤\$Bu�I�	a(�$(|m����d��u��^L g�e�]���p+�ĸv�9��(�ɀ2� 3�QGY��y�u]�Wkp�[|��X���3:jW���l�-��W�N -�0�a&c��ųQD8�:�U>a;���p���23}��E����)��n�_.�77j��eT�Zˁ�'�%�L�kf� �ڀ�a���xӵ'��z�ܴ�ޝ4ճ�Ц�#3�#�f������������=��y|dvmW�R�wF�Q?\�o��2��HaʏhVe����R�W���z�1��T��q᥏+m�Xe�wg �;Q
�i-�ju�FG�d�������#�B	+�E��c�-��{6���]%z(��n�ؓ8b�G�n\;fb�i�YEt��چp�.2�pP�b4�+���Vi!��t>�Vw��Dqd�*�$��a�w��{��v�Z�t��t�ŧ,b��'nM��ʐ���|̗L�Fci�kgٔ�W(^)�b����:�eX��E��`n��K`��vr��͔q(�v��Y�_d}-/oy��H{�9�m���N�:�0��
�32V�3��b�:O����zQb�&كeN�Y�j��ڳ��ClP�-jgwiT�o/h�X�)\uʟ\���{�+3�{dnR���&��w9���s���F��d�����x8��n���+�,˩�6)7��n��ge1�;
?s��	�v�H׍zq粳
L>u����7S��܍87���M,����\�m����g�e���m2'Y}{u-н��K�Xu� 63s0��6�\�Y���XP^�
�;JO�t-��58h��e+�9f�?��]��T���#��R�����2��up��v5 Z��;б`�w�y~83�7Z��El�;z4\6�#.�CQ�B���u��mv�G �96DJ�L���0�Vw.�*8b�N[��<�n��b�$�wW�� S����HΧ H�5݈F�|Cgz���޹�su��[�[5���\��WW,O�Ki�
�'�+w �����RZ��ߢ�/䫗۔�.�й'V�|����Q��b ����?m�b���YVO����Q�x��i���Ӷ��Z{xr�0FɁ�vi��%j4��e2θ[*��B��Z�n:Á�a�64�;t�:��Ky�@us-���z���)5U3�-����vjm<��X3�w��FR!� e�J��Hi�!X;q;�J����I��۴�[vވ(̬N8�b�Cwp�A��X��Ϊ_A[-�@�[�@��x��~���8U�S#Ը^$���qsL��"�3��m�N�vD�̡p����_b�V��F�K��m1\Z�%
�-ۮ#��H��l�\ �iy��F~ۻ�*=�n�s�u�$���>��fk�(e���M��r��O�&�r�Pu�ڜ�^Cx�g@��v��w�إqcxp��䆻���Wr�8�D�#t�Xֶ��NK�W����F�U�hI>�>��m_uI�c��B��M���{�=4P��:ðdv�vڜ]��j�h�1��R��B�0%�3��5��x�@�L��[g%��Z�E�U��օ��S_hڗ��B\Ӕ�V�Ƹ̆��@d��6���*
�[�ea=��{�w�ü���4�K�n�ꮳJ�%��d�B͸!����,9��&V$�����B�լG1���1*�B����pՌ�í�곫+f�0����
�Xo)np��� �b�L�3r����a��m�I2�ΰ�S���uoCRݸ�oV���,���Q<	U�xz���/����]ln.<nl\�ۜH���xC��^:R5}O{"����3z9�[��t�SGE�b�gC��}�.�y�2��aj�����bb��T�-�v�h >Ҵno^eP���!Y��,s�ȩ�&�W^`s�#7{-b5�O��-���t�����q����k�W},+�O���5�C4a�PI�����Xl�A��Y�/��Uq�������w>�&�p�.�˶bko	g�NB]k+@�M�ʔ��͗��H;��&p�%rє@��v鵴h�$��d�UC����S�\�e)DfeK�>�#�\)�$�¶��
�f�T�sn�\�|�a4�F�r�AE��{���Շ1Y�N6��^�7 "N���]��c>�]���!�u�˾�=�갫���8U��]x�;�����*з&U����	|�e鸱�h�C�Y�e(�d���W;�Ź�d��  ��%
�L�/A��:�I�֬�Ѫ�V2�vەϱ�6���^���YאI$WKY���'�(+t�$f�S�:���v�;J��yy�-��Lɚssh�-�*��S\���N�ǅ�Ied�q�`i�Y�3w��I[���r��h�B���g4�s�E�n�/���c}i�:�M �n��.����us g(��54�^�wx�ł
 NС|��j#N�0U64�T<s�@ᇣJn�:� E��I������7!kѐ���l]¹�"�v�����_t�d�8�\��L��U��y�u�nX�Ǻ�+�e�Do��彗o�l��&��:�`��vB�*,����zwV�C���Ȱ�i;��b��I�n�nҚ&�ִQ��k�.|3�)ÝW��
����+`v�hB��{2�>�6��]�;q���r�v�i;@�I�N�z��w���V���������I��d� �┒ư��⦻�.�pf�+��^�!�6��b�ن����	�;slЖ�b�*p֝c�9�PPSyQ�,e�.�яQ�ʡ��3F���q^�`��l��]֩���	�s<��Vv3�^Iy�$���@�JZ;��ҩ��;s���AP&�q�IR�fS��W|�@kGVd,�iv\3;:�I��TN�k��Wo&ۼ2v�X��:U�0e���{q��)���,*�T08�)h��J�8��PK�;C�m����o7��m�f]q��+i*�7�1��.P؎<F�Y�h^m��O���)&]�r3�h�9���Sr��:n¢�B]5/b#o�(�ׯ.;��V1�Ǜ�wt���}���qE�^�o�\���S1��y\5�AdЯ�bU���	��[��@cU3J�����]�(��kR
�����}5�~{w�v�p�G)�\4�.�ȋ�f\.�|�VR�T�`�Q<��粥�Ǖ�,�z�-����,[5���5��>�y��M�]���Zc��[�7�`l-����n��R&�tᬶ��!j���:%c3P4k:��z	:Y����P𜈔ݡx�9���ɢ���kx��)���1�m����4a��*WX����>k��/�Gӛ�D:�8�[ˣ#Tf�,b9̩�m<��X��F�YL����
��)LOO#�������bM�0 f"qZ�L���G%u��4(����V�gj���:j���`���/�eU��$�-E�v��.-L���W;0U� ]ZF�Q�����k���n�2���wCt�يi1�Tw&�b�p�z`l{w�������Q9p���7&�U�ʘ5|�L�fVӛ�k�.U��YW\^�uyR�@���`��)���f>�5yp�x��y�j��t7h�(M�E�Zzvn��9KF',Ԩ-V^FiV�eW1o�qxr��GN�\6��	*�mRڋx�O�Qd@Z0�Q6f󕏾�L3���}m1��n�T�1�۬q�hv�摱Hc���C�͝&Σ\�z���S���;_p��B���p��:��n�l�d���8()T��W�[��^6�ݪ��E�Z����PФ�1���8]]��d��4�`S���4��GP�� �Y�=�L�j.c�-�9o
�8 �De�����
jf��o��j���FD�����-Q�������ɸGe�	�ұ2�92��3.����ئtD��3�JaY3v�� bzmY@���Vi.r�󰗷t�.Q 
Y�)�HD4�N�[�>[�
ب�di9d���_wS�g>i��*���z�ɦ��[[Pʻ��&;�uz�r���o#����RQ�*�e�ˀ*;��TC��ȵ��Ƚ"���I٤�+ZBbkr�Ih�i�ܫu� }Q�:��5fe�=��;d9wuK�F�R��}7{WSQ��g4�k�}|�D������zT4C���͹eDi�r
��U'm̱&���<�����y֦������u�u���EG���Gs�J��C����b�Vp:��o
���u9u:�������d&�U��o���a	ɂnE[N���_]��z�:��1WJj_<7.��)�j�w0�3-ل.�m�f�Y��2&쳝����Ӣ��w���l,�{�!ܮ�j붕	�F�q�a�kiK�5c��ˇ6��vP��Y뜞m�e�02v��,�Z�.`���wU�!fe
9�� ���V�8Zt���c/N�U�ﭔ�X��^m��0'm�7�r��__1�Q�x�%X����,/)h�B���Ӌ�bD���e�G6w��s�1$���g,1�uf��*�˅��y�Y>�ڃgj�PM��9Ҭ����Ԉ�v1���v�jZ¤���&�zY%�#p�\�a�b�Z4�˗a�(��LaK2)AH,���.�o��=�3R[k8�=��O��Y�e�Sn8j��Wz�5�S�w�ˋ��ӗ��J���
��F�3��ӕ���bgtwDL,f&��F<�x��%��7f�p�-�+hɕ#��2�Ř:7m���%r�ͳ*d�vn:�2Zm\ɤ�����}u»*�,Xۘ�=�I��e�#-J�˦a�sy_z�)��(`λT����<�uZ]��[y�ha�s�]}���X�W+ݒ�sd��v��,oܱ^�&*���I�I���D��k�z�̰:���Q՞�g^m�]mm^G�M�F�+R#AY���qG��L�j�?]��p�vֵ{��N����֦ܥ�	�zH)^.��b�ƮapV������+���D{^�@ի���52���\��AL��f�������\V������j�;�a�^ѥ��;w����s�s(ά4)��9kvsx���-ݫ���8�h�g��}��6��!nJ�Cm��=�|{Bڄl`H1,�A�!;Cn�f��A���r��;Ϥ��Y�9ݹr�Y(�ۮA�����w:�B���!xbÀL�	����¬�U�:�˱��t[��7*ܓTZ�e�N�l4;��lw6��+j+y�2yz�Q}��]��k�G�,l�$W�3�`�i�,��՗Ml���}��IZ�/.K��n�+*���X�\��j���E��c'C�k]���#pmT��v*�5������h9���;Θ]a��������Ѷ�#j�&ڸ�hf��x7oq\�;6��X��1V�%Ve̍��j��Re����
O�PҰv+,�ӈՍ��ZI��q����i%`����t8�eew)f����S_;;�F�n�Qn��q�Q�(*��ۍ�!����5&)�P�}I�@W +�.�o
�C�:z.���?�\�Ŭ9{����y�߈��{���I���p����G�X=%��
Ѫڕ9��]Y;Md[x� �(3wή�4l��V]�]@2�J,!�r���R���Jnm���m�����y��ݗg*�ڕ�IB�T��'�z&��	��#�Y�C�V�5������|�� nX��޶�zwIomp�]�mN��-t)C	J����#B�ÊL���yP��Dx�r�@MރJ[u�Ĭ��	�"� �g�ޒ�U��»&BT���Z��4����ܖs&��5���������n�e(�f�ϗXVn����A4�W�5u�լ+p'Dho��,��u
֫�y�=]����㿄��Nb�X��C�X��l�ݶ��B��4����,�ǮB)��[���+2�Z��v�Z�t%G�w���ks��
�r�{����*�kxi鮂z�8��T���ُU�', FD/:�)w��M\�c�f�����@N]U�^�*�oZ߀K��U*Wb��4=��8h蛸jB�VT$`�a5f����������Z��VQ�U 3`�+��2NP��\����8uJ��!�����\�fU�:eDv�����n��i��ֺ'�-F�BеU��mb�ң3c=�-\O-|�40�q�tgmD_\�q8��7]�x�����h����6Z턩�:�m��\V����7��/��[�*Ka�苚����^�l�F�N'�f*�<�]ւ4v�И\�Vl�+pΗ�pI�Z�/G��0t;#�A��K	��)��#�g�&��<���k�(�h�B�^ �^�4�0�:����GI�z�DY�y*�����taS��T0Y��
��toWV]$�\��QA��@�������>p�۔bZ�����h=��X��*���.���8��m��u�n7����WT" w��wto���*�4��/:T�	9�]�V�V�5�@�)�,����=֋��*$�u)��7ۣ��$9�֊��Wce�-X�f�-�Z�M�1M�!g(����	���y>�xVN:�S��zȅ�``��1��&n��ߎ�n��T��c'N5�:�k7�;��]hѡ���lsP9g��gY�`sƆ�,3�m��@�t�D���b�[�z���u>CV� ���Յ�sC���g�����;}�r�v2�#�`�7J-^v�5�P՝KR&�0��{K%�a�n]��fageʇ�� ov�^�ˡWme��׿s��Z�d嬬��5���;�h��/cz�Q ��	�B�]2{e�����]���L��5��3��+�1	��g`��
H���Җ��T𗌬�.�P)�Zn���v^�6]�K���NP�E�4mj���'�q;�Ӌ905��ſw^���J��$Zh�M��b�>ާ��,�mK)ZC�j]�]�C2E�*V��$�b �v,�AR��{b`��c�H�Ux{����ݷ�(��5�Y���������AOq�B�E�]��5�bz����fB�����S�^A�����w� T�VD7�ׅ���D<Ć�N�(�C�C���X�f S�q]9v��޵�7S;uv�g)�x"�cӣ�DT���rj�1�W�f�t��Ȱ,.k�VoN_hP���;�Cp��%[��[���'c5y}ElE�6�'5Vvj����[cP�g�:)�o��A&;س�݌�{�t��g[�J4v):�'V��<��}���Xv�m]�xJ�:ta�����^ ̬#��V�_ϫ��1�Wxg"���-ՓgT�v�2;B�^t��
{+X) ��ͷ����F�X���E��/kj-:R��]	�% /)*ܨ�b�B��5����΄QW;�CO��5Q%��(�SK���ޚ�{��2�^�2��V:��)�u���G�^�@J�6Wp�sF�a�y��$�Yj���4ŝ�o�Zq{_7����B��Xe,Z�������u�$���J��LS ��(u�Z�ݷk9kn��y��K��bXZ�`�Ҿ�z����w}gpgTѻH�(ERN��Ju7}��W Op:Le�����8�L5w㻣<�����܎[��k/P�I���8��&�Ν}+Y#u]��b>�5F:0(;W�o��P�A�Nu�.�Khs]2)�\N��m��L?]��{E��+-�m�J�%j+l�V�� ��R�¢��ch�X�-�ؕ*ءm�AIm�,����+$�eH�
�
["�EP�DB�VV,Z��*PZ��-�m[j��VQ!iJ�iR�V,D
�l�+%�R������[`�+m%J֥`4������X,�iZ�ʊATd*E ��!ll--IU*J2��P��b���D[E���R�md��l�-�ADJ��Jł��E��h���
�Ѵ�[HQ
��eJ+-im���
E�F��cR��Y+R�XV�
5QKl�X(�TAEYQJʕ*V�+*�ҠXȥH��XT���
�mkV6�E�X���QEF��+R[B���eEڭ~��ŉ�s�H�S*W$w��ݿ!�;�ɩ�[0��{�∲��"�F-�\�]�w�y��q/Ru�pj]��}���s��j�TC��������W�Ʋ��V�<~��HrW����m�a��yf��$*�����]ԽCҹ��(_�������������g��lp��O0jPOӱ� �T�H��9�1���Tt��#&��q�eNCsף��Y,ձyΖiݾKP����Hݸ�	��^�5�T�Al��`t�c&��x��չ�)�賄4K��S�'���qhק=��V;�<d#^ p�tɃǼ-��pE���ַJ.XXȣl��6��옩o�b�¸�*\X��VDQ[���5�(u�Z���>}�W[�Vn�9�hR���<Yv��;1�lw0TC���k�6]�%��5���ꈝ�3"��A%�����Nv%�>
�����H~絰߭{B�ax�crw^�5�l�%����=7�pv��k`[�b�=v���7;�m#��R���UY��m�����Y�Um��0m�ɖ�H��:*Y���������&Nsչ�}�%y3׷{�G�>��V��vi�닫���a�Wz�oW3�݇���=@Uڏ�{����G�T���z�elCJ��K�U��V����g����΁$&VWte�Tzfĉ!X84��Ɏ���1WK/�����:`B��ِ�3i�+*��荍���SE�ؑ�PW=�cv�׳!ʇ�͔aG��
�gu����9��	�B21�9ѲB4�����i�xk��z�x�8�Ur�{L�p��sK��
��]3.\�b�a���)gx�VU���֩�*�t�qzȈ�;w�M�͵�DnD��>R'�Vz82�%��e���l+M���s��hdf�'�*|��W]�ln�v��L��=
��B���J� �g��Z6�kϦpI����hoY�\��͌��1���ԦTmHaH�/PM��	UtFL�1�ni֭qAS��<�0k��֢;d\2i��gܺ���Pw5�7J�:� ,�`l�l�3ӡ��x֜��z�"��օ�~�] ���T�����G\���mK�)R���1-�2� C�
E�L���@Pfb���p딍.���hi�Ż�Lֈy#"��9�]�z�,E7w��"����:��U��j�v� ���O���R���]i�9�|�\�;INNuF�x'D*��T&�9ӓ�$�m����U���8���d�}z�nI�7n�fv�f�U����G{��z��kk�_*�n��6������w�����}n��P�ݥ!}]�<�;s|�b�:V�3�* *mH����:�u������/v;2�wj��?* /�P�Rvk� ,!������{u ��ϊ��?!��o,�2�
s7����V�
ڳ+|��E��d]�`��np�@�]�PR�'�RU�E�� ��y�l-�b�D*��Jt�{��R�L�c�y��nɎ�}�Vy�b�&�V<;�l�Ry�����L_�������7�B�J�sQo�
�֏��1�>1�Q,��[�.zz���
l�|��W*fz8�a�@�t�
��W�E�����E��N�ԭ�tF�z��r�UB�;�EZ�����Z:ڪ�k����(z��~2���ɭ�ó�z��W��u8��T��ثٶh�~'�¿d�{������Zn+yP�edk͈��s=��9Β������ ����hՎB�9�x�4..��b�I����1u< t-�.H��L�� teeh�D�<�U{�Q��+�"0���=�8�c�Mٗ�{�\���Kٷ �Tcl-.��E��l�H�U�l��l
�ű����n�h
�]xj�/L��ʢjc��Fe޸Çn�q��,�m�#��,'S���A<�@y-��z7S{I���f�z��$ Yav��h��w''ö�G�7}t�y�/ř\���'y�7�u)LSf�nP	F!H�W.�&a��i�kpTb�mË���%R������5(e��,.u�#��VT�-ufy:)��^F	��^t�x潋�)WV��}\.��uV�pHj��V�=�p��f��uހ��+/Z���e�?p�lSϢ(gz�Dl�U�	�Q��{*0F9|:�:�e�C�5+J����ܦ������4B�y$F��f ����1�<�X���m{��.r�4�$f�������ckn"ry�PbS��M@͝l�q ����Ӑ6�2hdSF������s���W�' �!�b*����fLG1 N���)���]�"+���-Z�7��w-P�����@���64MB��w"`�L��b,@�¦a�uY�3#�Ŵ�޵�0�!��#�ƫb��k�~����X=���PF�9�}Q�I�zuZ�;=���1�_ G��u����.�{γ���a)NC�{N�w"_-2WZiU͜2܋٨!:2|�a��3�������Z2��1{���[�٣�����|z�n���LP�:�% uR�w�T,�]F��9��ӹv-E{
U�p�ك;� mh?y�\�K6��67d=�:ȟ`�N���xC�*�Z�2;��E�pX�Ư�۰#\v����P�����Y,c�aW�3q���f7��F��-����T=��~
��4�xX�Wp_c�ӫƵ�fS��K5�$>˾#-��'tr}obr�[U�N�! ��*.U����3�k�`�#!g>�)U�W~�d$"d���Js���[�PE�B�1�)v5�nӰ�WE��*�Eu�j$�B��e�v�+s��Z��я13�`ʁ�E�Z���!��ϱڙ`&E��|v
UȘ�Uk3l�ם��&�K[�T�,��+�+��ɉ� Y�� |Q�X.��X�����~�{3�*�";���q�CUm�vÛ��,*��|��z��7�`<%��!쫑��^<�+s�x�ݔ*z�jJOBa�6��w ڥD7Nd��(9Ԇ�u^K@�_�:�\U��6��:�*�3={��0����r�P�T�q���C����Q# l��`t� �,����M�a�~ߺ��Wc��,��RFe(��Ϫ��r���,l�AǪUD(�vj*܆C�}�#��f+��6Q�L����E^�#F�Prb���ίP������V �;�39m�"Ogq�z�<m�]Y7�e�6K��h�7��b�{�?Ѽ��g(X�ȝG1I9ک�bK���O\��3Z�vɥ{��x��2�]̇��1X����1�a�\�`6�P�#���eV�RѸ�LI3�z�zGjV-����C�HׇR��m�@�TT�V��rوP���`�ܣ���4ێ�)���OFK}�^�I���N���侂�Nv'��:�����1X��O��}g2J��Xf�cb-���z�&�`��1�=\⶧��o<(\dU�>>T��֙�Se
�-nŌ�\�P��sG`TI��6���hE3�:�ݚ�q�1v���Ț����s�u�&�%C}�N!�7CtF��t:��xv$�����F.�7[�5
rd�핂��s�!����$n	p�db��b�:=���uc���=��φǀ�����c_N<�Աt)�~ŝ��{uP��ǲ7�GX���w��H���X����:����ĕ)e��y.�{��`��B�%3F0o��1�L��s�r�N܎���%w�U		q�^r�u�t最�;d+SC�Ka��"���xJ��`9�ΥX:�`ɣ�v���K;\W��[*��qOb�2�jGyH������Q;R.!X�.����ō���]�q��QK�Ш���fpQ9H�ZK�`5ԓNQ����F>�A�d��-��/0P:6z�!���B߯\� &��	���+��<y��,��HӍ��¸���ݼ��po�"�[5�sFܴojNE��tD��$Eg�pwh�����f�W�v��ˎT���m�n�c�q1��F�\حg5�n��]���o�V2X�D]å �$��8.vUYBG\����>*\��í���N
-�{���02@�F�����r�z6���!١�O� N���rS�}!Ͷ[�Ԯ;�J�����T�C!ߍT.�%�xn���a��٦oxw0�0��[zڙ"�a�a�z ���P�� �f�� ,*��;O��-����r� �>�^.o��=��1� �M1�c�Dh�-E�0z=;%�9��5�1�����'V<J�$k�P��B�VV�<��� ��T�)����o�O|aKt�܎�����ؤS�j��Z����Krb����r�QNj��"���>����\X���Kͻ�y^�Il)�h�X�L�vez�] a�}C!+󃨻ݝ�M)�a4�����^��6����IG�d�x��6݅�4d���_Wg}Cױ?)�.(���s��ժ����`�D��neХJۥ�Xnؒ�m�d˻Πs5p�y�(KΛ�^�l�Y�m�h���KBR�����t��ovp�vo%�P�p��sT
�/ry<�'���D#)r��9e������ϙ��j��K�Cj���y�t
�Qg"�lU��f��6��K+���ت�����Qus�[^��z�M(��W3�wg<�%&���.B�ʅuˮ�#�R25�5���d�+25�]������Y�����[���ʎ�]��H��ڱʔIx�O�@]��@�sl[�m\h���z�ߪC��ڇ-��R�Q���Ԅ�Asޖ�x&c�k�	P���
�\����'o��Z� ̐���Nŋu�6��`�S�#���ʝ�Y�6�Ա����s��U��l]\K�ءhi�w�Hd(�Ӱ�[<�=s�.,�ݓʜ�&��rL�f�(��2��pE�}X�N!��t@�9J<a� `�r﫣�Pw�U�s�̈���E�0���Cj�{$E�����{�Q��<]*�����t�A��"���|��>�D�f!��]���;�07X�*�H�)F��vT�M@���F�]��.xSt��\�"ꈞ�,B��y1ā8�qv vjѹ44j�w"2�mr��NU��]7�;+/�GnCѢ'W.�D�����������*�"�n�f]�W�)�$�5_f��4��Z�u��
����wl��K��u�՛5&���5mqs�ڀ
��k;	���_l��8��c-���*�K3�$b�M�8p��Ɖ�@�Gqb&��l�1 `$��MMv�.�(<�U��)���5�v]M�nb��x����FE9c�P}�N|F^���+�]�Ҵ��FI<��~G�1�mK��;@�*6/v;:�{"� �B�AZ���wkm��>�먱Vi�A�UB_���J��'��%�O���m�Yp�����N����j�Rc2���o;�ٟJ���O��G�6r�*�r"���(Y��w�ڋ�?<��*!�oS�"�Īga5\g�|TI�#O#>������c,��F��̥W�9���=����U
]�"݆�8>��j�R6+{��^S�o�7�1[��!��t��W�
�j�Utp|�R��hO������X�Q�+S#�ɑnzn���k4^U¼�:���pS'��B�Ȯ�j;&R�OF�Ga`V�t�ۼ��O���b��BϘ�>߃�b����bv&7;�愱UlFp�Q�;
�eoU���V��i�7]�*b����QLTW�;���]���i٢��gN�<�#�Yg���&Z��$�b�X�� �zskۼ�~z�ӈ���e��%�ܪ�k�'�U��X�F;e�>�wo�3��ڤ/k��7����O�@2�N�io��5�g'e�.�]�D�?]8|�H];�j�	ܹ�~�b!��E̗@�H�)q{��U�?#Y�z�lt6#v�ɛ�B����D�3���P�+ySF��o�����[/ݕ�aRsc& R��p_Y�t��ƺ'_���b�h8�������W�p\� �y�t[w/��aw�m��8U^�:6����ox�+����^��E�{��u淐��E1��$D��qtR����-ߟ�l�NV/CN���!���y�����w[z���wuq��}�^�s2	h�����y�}�^'��K�u��{���.3�%�l�;x�RÑQ툎;<E1ȱ�a1@ԑ�>K<"��
�j���NuW�_������s6���L�
�1e��l�RN�l�I�o�L�"GG�
g2A�yΛ+�~��"�~/�����Ǌ��o�2\!6�C�nsC#!k��4Cñ'̓��:M\LMKD�
�[��n$�\rU�
��6+Ъ�|:����/tB4��������=��Nf��(��j�$�W|�D���t���!3N:罱�:�AfT�Gvh�V:�|�>wh^t;#:ɗ�Գ��z�a__�1����{�3��u�-�)\� ������<��HD������Ǚ(�˓h�2�f�a��顈�᰿����U�z��M���.q!^�#���Q����"7VGq�noʻ��!	�"q���. _=͈�{4QB!HÈb�hsBD5�	v��v:nٮ��^U�|�
��෧��� h���͵����<�,�;�u��c��;#8[tE�Æ�J�s�A����Q�n�̘�K`��wpU���/6��|w���dF
�wW'�L��hX�X����ɀ�S4;VgsTݲ�M�U�U�=�SM�s�YhJ}����YBը󅙽FM}t[��/+��c@Zg:��1e��:��M�BX��ou��Oy_���TFuC���*Be�&K�ʍ�Y���c�tk���y}�Am���KJc��!�Җ�G��̂�t��T�C��]�6гO�y�^��nڨ��� Emަ_v�-QJ˩��ڧ��Gw����鉜x��Q$<����f��Me�J�9VmL��WB�nAAK
ѸU�����;���*�9�,��ܤ4�d�ƾ�� ��:K��+:�%o����:qv�2U�.ggA���afىԃ�;E��W6'X��&��-����Q�u>n}��Bt֌������:���*y�KF�^R��1�z9��U��XxN�[u�L���G%������u��
��^�G�˶�Z5+w���o�`3h�c��f�����2�m��wD�{<�}�Ӳ�̏�hn�#v�<j��T��]�QJ��:���W�u;�ݡ�1�e8�}{�î�rTZ�ظs[���@slX؅�_m#)��8�u��'�p6�_�������wT��,	u�&�z����鹙�jSv��)�����m򷎳u�1��:m���A��`W��������.�A��e�>\#Ԛ^��iJ��L�Ӗ�d��ӯn��ݸ�d$��}�)�����u�p�F)·z��x��ݗx�#�<&X����xr1[�0%A3K�1�vLv���*d]�"�����;�sK�k�S�Ⱥ�%@�<�^��3�۱x��s�vҠNe�&�P���O�Tk;��e����#�y2��`3�vkџo^*�h�^�ĹY�1��B+���, G+���E����۫��q_>G�� 
��He媔�%�a��W�v=ʸ�(�2�]ma%�LKr�Pe��:8�1n�1^���-�n.09z�eVs��Aw�t=X0َ�`���,OxI�֕,��pVO�`�X��`��N��&T�����x�l����{�P(5�V@��j�B�җ�on!��2JVr�q~��3��<�x�]��e�7Y�:�f� 僧L���(
 �@���*1�c""���5��,�,����E���QjQ*��Qm��lm������b"����Q�֢-������[R������VX��+*V(",-���VѪ,�T���Q�X�+Uaj��`#�*��#�,mQX�H���Ab��ʊ�*������Ec�*#6آ���ԶX�E*R��TR�cX1#k+Tm�U��J�-�����)�h�KX�(1��lV2֕*X5*�U-�ؖ��miJ��
�VT��F���j(# QQJV��P��UEV
(+Q�PZ°X#
�U�²6�5��*UDQQ`�ED��U���b��ң*��EiPX#X-,X(��(>HY�:��]s9�1lU�C��5K���h��z"�~��W�w��Z�i��ټ,ʽ��9�O����m�_mT0]���Z�Q����\��b�ņQ���Pb������)��@�q���m��u�y����yVe�)���ZӾ�����R�=~��Ih������kD��n��}��eN;^5�9ϲ����i�YM���;d%:e�ձ�'��h��+�����e�j������֣E��~U���]tu�Nf8���VK�dZ��+�"�<!*���',LUU�wn^ja�cY휂�8����>����ʽ
�5�k�xpUu�'+��,Դ){���� ����b��0��tS�s�\���ϒ:���t̀���5ƥ=�;9U���r%�@�hvj�x���^-�S+�<9���f��2�n��^ ]�r,��+�ܴ�Bn��p�b2�*z�C� \��T�?����<� ��^�[�w|���{A
�x��n� ��DD!���뤀���~T�>/Ta�ܫsw%�펽|���DR�)��	�b�=΢4T��,W@��npS6+��ك�G��H��Ѻ���ĭ�S��}=�&�2U9ʺif�O�cw��bn�#6�1vG7R���,t�;M�v �"ũfϵK��t��u<�_�^�/d|3�8au�SvpƬ$p��U-8��[�PthNV��M�3�a��"�Oek��F]�3c�K�u�8*A5M�Q�,uD<L�Ny2A�1F��¦	�<� m�ȍ}!��Q�ۛ���#,�xU����~�
ͫ��"T�h"��\}�P���1���޾зݼ���P�={~Hlofa�!�P� e+�5{���RP*��8hiOM4��I�Oɛ�:�d���jO���7��	݅�4��l ��ƱW	�]Yh��3�`>����������g"�b�e����ڲ�:����/���襓=�R�1�T��� �����L��ĩ)0-�tˀ�r�[s��7#H�Ibp�����[��%'vLd�L@� j�2v�e2�^D����R�]���^���Ŧ��c3W�N�޾�1uR�b�}@��-��R1MFvS�:́+��w�̴���srB:��W���?i1 '#��T��E��Y�,*u:���b���2*��
��u�W��nkfQ+r)D��U��![$&�$5`�6y�7O�3Y�3M����2�e,)c^���3� �,�]��3�2@����oQ��,Qk*�M���zN����U�P�j�XU`���qh����Lv_MF��;�xws�����n�}�j8k����ޙ!����D����Ò�lo)7�pҥ�{�=[�[�����b�����T`��Dc���Dl��*r�x�{*�N9b�6l�WuH�"=�Q����;�9��^9~�	��
�{$E��f ���zШ�Ǆ�ɫ�N�"�{�U*��JGZ;�K�dR8b�c���M7A���3�:ߊ��
��_N��n�X5�b�Q�}�o��d\�m
2)K�.lG�#�EWqb��y1��%�pM���M�1_{�R��;���/�f�+�l�k����Va-Έ�CD������rf6u�%oY���u4��]7���B¦�0�V<���5c�J�*��ڮ���g��8.���ޓ�uz��&���p���߾�J���~~j�O] 턇[���j*�/��stv��u���{޼��0*gx��V��BY�ei�N>Fߕx��G�^}Q@�@�LDF#�C)l�ˣ纅[��.���p�.گc�G�6##fh%�>|�!��8gzk���P��u�̼ߜ1�5�R����S$TX�A��`Me`|TI�#i�[���pʓ��J���v�)VF�늦{�a�K-��=+}�^\k;���jP`�5��%�խ9\r��I���Cw��B����5�.�yw���WT��t�ǵ��F�sZCS�M��8<����81:�(����^9ŧ��ܒ�>n��pJ"���>>�P��_7a�<��S�U�����Q3Ւ��˕8*�v��%��.X��)���tJuG´>�Z2��;1|����Gy{Og%Ok�Kn�aNP=99Y���n�K��"�B�5�* �z��(���)yg�L�������0�˓�f!�.6=��ͱPԣ4�yI�#W��خ�"z#niF \�(��f��T���!ڔp�~���Wu��l��vȵ*���̑�ԣ���#&sk'��-1-vq�7�����C���9	Ox\���l=ݸ���юLx�T�A�C�:yX�ˆ�Tu
���خ0y
����:�7영Js%�}�>��ܸ�D�����Yva�|��(�x�O���5È=��d���/yR��畊�;!zq�$W#����t�Ō�<4��L]�`�o������	�g��-ߟ��Δ�b�4��]H{X*7����6a�k�Ԍlߔ�"&����U�?kXURs�>�G����U�^N0��W3���chO^d��/W(�`]X�{L>�#$�(2��I���w����3b��48�+�G������yU������3J��t[�|f�!��nD��S�%3MMT�^�߫����	蜮�[
�・��uA�an����v��b�����V*�:m1@Ԏ�k��$xk�<��6��Y�r��k����>n���Aۦ�-��5Hq;�f�L���>��m[�+�oa�c�y�6y�.�*A���b���4�2\!6�C��!�tF��k��4^��y�;���wl�;�T�>����ِ���t�$l8B.;��P�`(���H"V;�L���~}����Ԇ0q�~�Vb�a�k!ң�Hʃ���#�HANl��S�I'7��;��(LB���ouoL9������W�P��Lь=�eR�.|��^WM��=����沕+��$t$bJ��n��q�!Z�2Ca�F�P�\���+��i�Y�� ��{))3p�

�kϤ�U�М�w��V	t㌋R:/HX�<!D����`��^W��Œ�����F�	��&܅Md7���VT���;��i��^����(r�C��ɧ׭zyK���f��<6lR�H�] ����8.vVNCJ�ϸ�钢�p�]53x�tT���f�E3��k����x���4�s@L�_*��%�� ؐ��rƒ˱Y5�P!��wo�WGH~_E^�&�����u��wK��{͂H��񓔳{�-tUb��e��	}N�5�ycn�|�c���[Ƴ�7��T�p?�v�Y��� ��Qv!�)�i�#gvC�S��9�:-p�-�[Pj󡆬��{Cb�(q1�(�רd8 �¢���\_	��8b�#�m%z��j[��܍�	
��/���6�%�13Y!g�¡��x��"��q��+ٳ=�l�*p�~ꈦ��sT��69�F��L��L�}�neV����MAȺF6��yј;f�����nj���bw)���O �T�9�Ȯa��+�,)�N>����+zg�u��� �P0�-ɋ*��>�9
�E9�>������)�ݪj�kU�b��ZH.f���/k�d�)!�k���*C����T�1jp+��2u�iM�Z�l�MḒ1��
5%=�wM`n{ҸKj��Z����]�� �=-�$yE�����ڪ�O*�@��;ޥ0ʯ5L[�ކ:��"�CkqY�[�ϻ���ǟE]D�@:�V�Sg��Dc��ԩ)0�L�r>D�>��P_q�<뛋m�h�*ryS	4Q֊���0Ӽb����.��J�	jrȗ9��Ū�}pޭ1�n��Z��=ذ!s.�g^P%j��Oj��glY�A'`�l��X�N�$[�@"�og��9x��R�}�e�V��n0⼥,�9jTYY�UB�܍��5��TM����O^�:��!�n
et�#�kk���x��4��Ģ���<�I-�-��XՑ�Ϩ��86mH#U����A�t���u�YYs��h��Nz��z����U���}\�jˤxJs^��V
Aq��l5Օ;Hr����oz
�	����4p�	P1M�8�"(V���l�0���Ճ���n��>��fv�������8II���>��6��/͟DV?S�!��N�R��!쨽���Bo Zz�����%�����^��24A)�
Fb`���Q���E˽u�N�Gd���J�hfF×Z��{"���e�WA"i�Ú0�΃6U8�i�D��7��J�����R���c$�B��S��.
����U�X�bfLA�$�ر�+ʢ'��1o��p�&�ڝ�3�$c�M t���[�0���S0y@�[��Sհ�>Imd��p�`��L���6\D�nK�YFb��c�Q�Exd�,DL�\];�������M���`��������oDǗ��_J��)vo$2�1]n�}X,�ے���L%��pf��׆�'V���'-��d��\�=Xr�ST���0h���
��e*�yb��{g�^��8�o���-*�0�[��mv��U�VG'X|��yZ�7������'Z��C>����+jHf�ż'cNaQ���S�N�����:����+��S*<ܘa�S��r�u2Aɨ} �維�q�|�ท��M^��nrz�Oa(�̅S�1�'1oP	U�ݪ�;G#�I�����%�!�#!�u���5����O`_N`�w�^�]1yJ!���1 �EE�T��y4Q��x���Źl�J����uvR��w>S�,F@�q;j�ψ�P�޲-�C���j��Yι��a.����;�EED��
,E�
³q�&z,C�ў(#�{'��}H8����M�XX�j�925�"�m��J+ѭ�R��"�B���5J �z����|�ς����y�5��F�[����O6�A*W4������}^�-����>+���J��HI����k�M�5~>��g��X1��a\�;�mR�"t�N?R�1
��:�N����s�z��hz�����nr�lt6#v���~�rcΗ.�kpmY+7��cG�{7M�8�,���Y�)c���bz6�d�l]J��]�}*�	���!yt${��Kזb|k(��L_d���_3N�;��.��L�l�����D��K��˴�f)]k�ɽ�r�i�É^��a�ͳG�-TU)��I�Q�uأ�ax�Z.� /��^���������*b�}A��
<z�xO\%U����┠����;�9������o����W�6��Z���:{]j�3�p;Mն���,�O�y)�"<Ý��M�W^��hX<,�W]5����SgX7��C�$�3R�R�==ݘε�����
�.�'B�dDך���p~%�M�aT��[�/aug�����H�Y��IS9<zb_S�\���ԩ����*��������:����2���.�c!������sh�v鹋l�����F����&HhE�6�ҩ�B1��\u.�IPUwH1u8d��9Y� d8B76�C�n�Dll_��Z��^�N��e��kw
i�2�}�h>�S��y��0��5>F�s�VÄ"�1T9 l��(jE)윩����S-)ۼ�=�>�E+1s�m���|���6�?y�'����%M���3���*k|�Y�i�"���Q�C1��:x-�ߡ
�Z�K�r<"=����QH)��u�H~N!�=�d5���f��y;�<H}i1
��<�mE��,1>�9��i��_h�c�?0�x��|��%CWaK�� kf�o%��^ϩ�CP�Lxs��l��_��u_��q��J�d��m0B�[G=7��9��=�N��ȴ4�p��t��1)e��R�[F涐f����Դ���B����Czv�������������N�hT����xz�tV��O���@������r�$��'ɕ�!Xm�r���C�R8���_~J�'��*|����<9���&3}�,6���y��SL⤨�5�L�2�����oUt����#g�f���
 q�lzf}�Y4��
��sՋ'�gR~qE:������|�O���C�e!X|��d��'��X�sL�%~d�QO9�� Q���*�$Y.i�����aF�'�Bws�Ioފ� L����YY�g���X5+7�'P����g�a���+����+��,�@QC�p��}t��>g2��&�XB���m�2k�������kG{�v��-�?w=���8�Y*c��UT���<氨,��A�?No ��?&0�V� �l7�4��TR�fa�b��c=�ɟ���6�|����������l��& (���������;���D���@ |>�8�a�TP����aP��qݬ
βT��AE������M$�o,���ɮR��<���>C�H)����'R��g�O̟�`�Os�'�]}�jʌϢv���5�0<#$�+�w�}���[=9܇��|�*O;�"���4���*N�Y1��Ms�l8¡�QA�O-�eA@QM�~7�m8�Ri
����w�B�沃�C�S䟁�0��c��欟2��W���w��
~@�k>��i�NfC���P�w�������o�H�+R�3�,*~C�bM��n���8���H[Jw_e�����_��R�<%��>����E��NޠbM�٦u���@���f2w����1������ɵT��a�fM'PY����
�Af��Y;�Af���Sh|�F �#F	�y�s}o�\~��Ǫ i�{�=�V,��|�iZG�+5�& /��a�;�>�=CL6��y�&�V��Y����Ğ��m�M���me���:UW�G�/p�_��IW|"<�G�ǆ�O;��'P�R3'�>q'�Qg�Y1<d���3�T���SL;�Hn�Ųi+8�+5�"��T�)�����
����e՝d�aV`�f��_��)/�pBt�����C'uY�̊�^�Pq�u0�Dػ�X��h�;#�TӰ�jݰ3n�3�n���C������(�,�{GK��ۜ�n���&�w"�eA��e��*+��fc��Y��=����j�b�;��#�Vs}0֧�|�<�9�
�c�ݡ�`cwGNή��a=v;��4��ͽz�G����S}D
���7EY:�QΌ�[ũP��G��j���K�?[��#�������>�6�=/j��k��´�6T5���}7����8�𱵵��˼��S6ҙluwSÜ��	�BG�,��-�]�wjg����qЊt��h�n�k���5�e|� ��C���Y������<�F���pD��l��W�e�Z�'�H&�Bn�f��)���8N��i�jg.�V	��C"˕%ǋ[@��l�+��HK�aZSp��!��s p������p{��qxQ귃4�֍<��7���tD;�ٵ:J��%�iVSx�/�fE�KbWx��}����X�|h=U�YN�d

��%��w�Z��ҩ��g-a�D���٪�2�j�_4��=4�v��W����yS��ٮ��>C����^+|�e�K�V�����`- ʫ]�/{�o���ϐ�<!����hQ+��뭷&��fۼ(C�Vܓf����ؔ%hי&Y�B���,�Z{N���J]sj ƖCus
��h,�k]�f	�h5�H��;�k�h�ae�em���9σ���8}Π�Ͷ`�5��E^L������5�V[������ݝX�����k�Ǣ�p�{�1q�x��[��8 k;]ݛ|�]��;�j�@���i���F���f��ַ1g>��[�Ҁ�uW݌)�0�]W�����԰�v]���rf!B���n��n��y�H�{��՗�5��72u �j�垮<$����|s�- Z�����^;Q�R��dv�V�o3���Td�����t��i�S�c�:*�ح�&Z�Գ����[sk��mqT�*�r��Q��ڏ�����}:�ۚ�]x��p�}1}ףd�Y�|c���X�1�j9��\}\��(Cc�\�^.� ��7Z��!*y�燀���k;)�/z��{��#vn� �AE �����K)��h�}{r���8΁�&m��Cv5VkG�@6���.� �Be;��0��b�+��R*d�t�h_dʃ@�X���+ӛ�������O��W=m��YI`�Gr�8�=���:���Ë��uڎ-1^+s�l�����s��k>�kGPB�YV��[� f��-���0�t��\��R��c�,��%�p���	x��#����F�:�ݵչ��ڇOW\�Tt�5��q���Λ��>{YW�mI�9 xf"Ҽ�4���J�*��:0�޵�7���1U�Sn��=�9O���b�U��"y]�{�����˿���߿�աD�֑*�%j*��c�mD*�X�R�V(#+D�U��m�c(��ZQF�ՅAAE�QD(-`�R���Q��@KaX�JŋYUP���E�TR�+EDDQe�E��2�"��Z�[X�e@YJ��j*�Z�D�`��B*�A��F��EEX*"��X ����AE�Y-���J����Q���H#���X�E�����)E[h��EAcE"�@�AdU�`�,Q�KX"*������*�V�"*�d��([@QAH�*�`��1 �QZ�H�"���`�P�U+��J�TTR5�,V,TQEDV�*�X,AQQ"��QD�*�VER*��E�2ڪ����
��QTE���PX��YUDET�������"��D�U1X�UVڣh�ʬX#H�(1��V$h+
���k3�K���+��]mqk������ך�U���ik�ї-�!n�&�������.�ޣ�!���Ǖ_�{� ,�F�T�iM��pd�3�?˝�mE+}�i�'�7;��VO��!Sgw��~d�;�0�����>���
AOP6y�	�eH>ٲ{d��8�T��7l5��Ohxsg���o�i���y���U@}U`���6��<O�~C�{��X|�f��������0�n��2b�{;�
M;t��sT�3�O3̓�4��
Ͳo��͐Y�J�{�&�R
z�3�����o��u�{�y�~��6�Af�@��g�B�AgS<�!�h��u��~B������x��bO��o �d�]o�T����
g������"�l*{�'��I���^Pw��|��~�[���׻����G��*��'������i�{�? T�C짛�!�7�!Xxf{�s)?!�(��gqěJ����CI�&8��0^!Rԛ��Sl>�£�-�)�̏��w׻�я�� �L{�I^�Ɉ�zʝM�fI>B�l�5l�&0���N �C�M��4���f�����
���]ɴ�'�v��\20��M'�Y�}̓L�%��9�3;�?}�	���Κ�Fޥ���Ȅ�����D�VT��������P��VO�`z�Vy�@Q`{�f���1:�P���ya��o��$7h~g�?d���& /;q$����g����T-��;[�}z��� d{�M�232�XVb�c����2~'w�%UH)�|�H��,��Xg)
�����H}iߔ��h~B��7d��3���wi��L
���=��a�l�9��=pxć�z���g��b��a�5�[4��V���E��
�<�
O۵�Y����AAE��yE8�Ri�jO̼�+<>��>�P�5�>�k�.~��y��K��L�M8��{�1 �Y:��PǨT��w����s�j���ڰ��͠(�VT׽0Ri'P�n�"�l�Ɍ8�<�M���i��jq�`"���q��T~�<��=�mV����yT1=d띠x}M0��~d�9�a�c>d�S���tR
|����lI�YP79��!�,6�W�� sv5���ࡴ���ȬQh���_��^�i��/,��%g�W���7fӶ��JʭB~Ka] �w�]+ ���kh�Ŵ�`�1�WkW�f:��U]�ӽ]:���H�/�������S�����n�]�V8=U��<����-d��n��N�yu��@jx�#Om�$f���{��ݶV]�8�����O���>aR�7��i�u�<-QCԕ��uIP��&��~>�i��+6��d;�a�a�s&�UT�����O�,ی��I���")��]�.�WۤmӮՋu.�"���h��i�0�b�����Ĭ=f!���H:�y�,�u�0=��):�f�d�R(��*w�~�6��Xi4}�M��a�C1��Or�x	�|��ؙH]}��O���a�� PQq�y��~@�<O&�`������|��}�'�s,��&3ԟ�I�{��H)���t�x�H:���M��w�����i+8�ٖ(
D{�@�$uk��]��}رAU��(��Ȥ�1
����g�L`�<A�OC�duf2T;�²~q:�Y��d����'�;a�va�
�d߾��)��+��rO7E ���l�q����f�j��FB��2����,������gg{�H[`u���0�:� (��w!���hm���A�����+
�զ���Ri��d�՘��WoX~vm'�+?2l�v<&<:<&<�Sa����WL��o,��~�_s�g��Z�Y�8�&�UT�LM�T�8���d~�+�y>�i�O��Osf�z����~��Sl1�������������ȱf�c&�o'����g�Ysy���>}�~���/o��7����z�T��p$��a�w��h�V���i��Z�����PQx�ՓI�
���h9��/����l=a̤���� V~I�!�R�"�S�}��o����:r��`D��f�sK��C�� Lx��Q��{�Otu@�V|�i1E��|ɤ�)*O���d�e�u�����u�o\�svq��y�օ:�����}�tN!��&��{������٣�}+w��]����Q���1Q�.B��Ag�;�p�Y<�)�u� lI겡䴏ԇ�a�g�����`l�Vu@QM�d㤬�N�����,:�w�<E�aR~�9�~ї�5{�y��}�y�����&3��CH��J���;��'��;���+0��X,�{� ��<ԛOUT�
� T�<3�Rԅt��&�ZOԘͰ�1�a'�}�u�u�0t����C��&�AF��w�wO����(z싼��e���� ���&��F�-�B*�;���K������Y���w�\��w!Ļ������^�ҵ���|�� +���XGj8���tz����>���Z��5�G�G�����d �b�~���ClY�u�0��}�O�Vk�=9�6�XV�w��:�g��}E��kP�|�ܵ�z���J��u7�@�|�Y��n��>9����{�����jɦ_):yCL<aܤ�<;{�Agq������S��d>|`�B�nw�5���5����C�@ĩ���Ri ��{��'Ȥ�:��M�|�l�ɐ�{��{ϵ��^�����[���a�!�?2z��7a�'���Rz�ǎ��ORz�}���'���4�k�>I*���0$, }��"���ۈ83n�n�Y;��¾�{�|�egć���J�bw^`q�,<��"�0�����+��&|y�1�+�����O�Vu�9�<��>g��g��oXA|���>�
����ؿxr�=̖�Z���L�=OP*bO��]����6�|��� VVLCϿa4�Sl6^����bC��rJŚN0�ߴuI�+<�=<��Aa�k�`�~�@���u���.W�qm|���¢���Yӽì6��7���oX:�PP�s5�S��y���Y?2���t�aX~�M}���4���I:�H)��d���
����@�Tx}�X�3��"e���������oS�IR?Z2��IX}ڡ��2�4ÿSl:¤�{f@�l�%f�k$�z���=7CI<B���������W~}�x��Y��Y�4NR_{�<�ǽp*=ﾙ�P(���8�m!�S��qP�C����`u�+?!��r�`zԬ��<�P�1 ���"ΰ�?C3!�Cԕ�:�I����+���Ͻ���L��j�)�/�@������tB����f�;�d>��Y*m����@���ϰ�:��ud��d��|����T�Ͱ�b?QIR
d{��1� l T{�y�:�)l+#�g>]�����+~N0�C�I���y�I���g��i9�$�����m��
�Cl1��Z���$�?2T���z����󹴞!�Y6˺xw�
����$j��x�x�ʵ����p*v����ஷ���y\` [��g��Ѽ����<9�_.�[���V��zj�d[�(����ב��$m�ͥ�!y+e�]���p��Q�����f�B��ύ�+�-��������C�tꂧ���F�MJ�=�{�foeW'ȯ� 	�0��*)�0���.Щ�MP3��n���$=���4�*J���̓���RVz��c'm�g���=aRu;�f�m��W_xs�=ө���﹟sﯜ�M�i��t�p�I�1Ϲ�w�!X|�yt�M��H(���̛�(bJ� Q'y�4�Rι*!��N:egP��f4�^Qx}e^�#7�[������~��S�?!��~�p���Y��g���<��Wi�;��(�P��m�����w�,�o��y��m�2~�XOM��q���W�T���*{�tG����
@�1Y�����e�3��������,�c'a�=� �l8�����ܿ{�q�C�qa�s!����4�3���ZLB�w�Y6����X,4�{@Ĝ�;�l<`t�}l��p����_~E��ݏ"�n��~���]v��%C���Q}`T��s�4�hs,��ɕ���6ÙOyC�st��'5��$��G�T���/��h�����H}l<9��i�T�Úڞl�~o[����^�2zʟ�I^���2z�lߝ�6��&���:�?[8���H
)�O�w?^ i'�T�<3����a�l��~d�9���:�_̛�)� D 	�n/~Χ��>9��]�o?~����H?Y7�XqP��w{�5����y�E��R�Sd6�C�b��<��E�a_7`oT=I^�}�I�>M�o��1'��LG��z����!fD�qL���Z�����6ɯ�����i�d��/�UR
q|����yO�� ��?&0�Շ5H,���4��TR�0����C�L�d�Y����;nROﳓ���BK+�?��l������a���!�3�Xm��7�`m�T1���wk���=�PQ0*q?j�I*�&�{�\�+=�'�s)>�T��#�@��u��W|��>K~��dӌ��ă�I��ޡ��x������<M��IRxw�E��*i6g0�:�d�[u�`�m�T7;�R�:�2����2a�si�UDW�UA�CGjLCmҖ�����\�]������C�{I�x�W���)�oNw���a�b�.�Ul�p<���+�|ktS�M02�3wH�g���P]������su0z��u.}o��񃎐I����É�o�>�i	�e)�[|��m�a>�sǸ�~���xxW_ ���Z;��1nG��|�+�&��Y?��c+%zɼ����
~@�k>��i��Շ��@��p����͡���,
Ԯ��
����s5���z�c�3�9
j�	5T�����W��́�J����& (��a4��$��i�d�9�<��aY�N�Xu��T�{�dڪAN0�3&��,�ć��Ӣ���&3}�I��<G����{��(nt�M���|�s�@�� �¦�q����1�v{d�Y�<ì6�դ�{�Y�Y1}kaS��c����i��^QO�4°�u�����f$��sh((��*Xw���~�0n�n�Hh��<�S����YHVM���>C�Hx�j|��~J�=Փ�O\a��3�T��g��l;�Hn�-�IY�IY�l1N��QM��i=B�q?W{�=�hl�36�y�����>�������P��[4�9�&�R����.�*O�nw�謟f�B���'�6���wV�a����2n{��)=@ߚ0�VT�ힲwVT*O9㯿}�~#%We�ﯷR?�>�c����
,5����:�����1��v�b,��(i!�Cs�͵=d��~�I�n�1�7��m�2{�d�f0�³L���|��d���}�Y~�s��}���UH)��9a���qs�g�B�AgS<�2�Y���u'�~B���(bm��bO��7��~�V.��*x�im;�4�?Y1'���H��
�����w�^�8F������ܦ��o(��z�	�����4ì*;���`Vq�i�Ou��
�h}��d>f��+&g��2�����Sğ8�iQ�h���Lq��`�B��?~O#G��N�v��%�-b lx7>9��J�U%q����*|��0�I���ٖβc����N �C�M�׌�@QN�}�_�'�N2~s��%�!�
�d�~Տ���y�8sQ\�Ԣ>��=q�LT�ϫ�tR
u&�u�$�YRn�o }凪�f2}��eg�����|���a��:�?��Ì1��x�I���s�M�M2b������^��x$��2�t���Y0n&$�A�QY�R��.f_�A#<�E�|�]�^��un�շ���MK�MmηY~m"<�{$7�^�C��X��y��n��xa����	�N[�ty^��k������w�:b-�o(�Hr��_ ���j��o������I_�1?�}��6ϙ7��{32��+1�#��Ag<;��*�AN;�5�)�=q��a��+�6}��ZA|M0�4��*,�%M0�1S��~���}:�����9Ͼ�R�J���?&�bC�zs�C�m��Ɉs�1aS]��9�6��V�r��a�7�)=լ
�'ua�_8e�I��}�K��1�*^�f��L>�~���~����I�<�N��1�I�u/��
~d���`i� ���񇻰Ğ����<Jͫ;���%eM{�&�u
���"�l�Ɍ8��o&�~A�����+�~�����;����w�����Y*�t/rO�O���C�N���SL>a_�<Nk�4C�%z����E ��y��lI�YP6s�5�C�XmP���@��k+���Ch
)?u}�=��u�g5���������~�_��18��ݤa�My�:¤7h_i1�u�?KTP�%t�a��
βo;��P4���M�ΰ󹆓i*�A��tui��q�f��������<�-���{Ϝ왪B���]�M�>��i�0�1�T\`T�<f!���:����<�E�N0���Ru
��ɉ�iXc
��0�J�a�ī��ǃ���]�n���y��<z�̵�Y���4����k��6�@�<OsvO̽�+�kl>��9�~ݓ�O�$���R
c'���`�B�_Y4�a��b�R9@�VqY����i��y������;��d�<�1��.���H�^�0�J+�5�����f�N��1N���d<9�֣EnK�����'�6I������_��]y��=m��9Yo0��|lV+$�^���`���g]��u�xd�ä́�a�*wQy ��>�fp��\�d���m���B������c��t�kѡ�:A[����Z[���o�&v�&}���[Ӝsc彙HiWq��X��Y���ג�׆����v;�`D�ߺ������w��#7�e۳h�X�j ��t��3�d��ǽ�s��J3݋�B@�YRn.��{���y;7��>���-��i��i��>�U\�8n�M����eOD9:1���\�^����B�#��ɨ{�� ]!yJ!���)"�����&D�L�E�#w�n�gyR�sb�i��b�yk��(V��
��!���8�c"ڽ52�+�֌�t�w��`P�x�oL)�ݨ��@��Ao���3�`�.AAWF��rc{[�R�no��Xu⏱Z�i�nm��X��)�8�yQ��F�©�!,�����\���JOd:�P�����"��s�>z�Cr���'�`�^�6'�9��mҾ�P�}�^n�.�3���9˃�k�*�lk�gct%�a\�;�jT	�n��EG	��0Js}Gv��g�C�GH :��ɒ��������*F�TK�I��B��|�]����f�W&<�W����:�W�V���O��xϬ�K����=u��[xAt��>͛�;7D��	��b��U���oa�١|���q��ѴaY�{00��>���fo;"����1��F��1Ev����@\Oz�C6Rb��x-�̗��u�G8/
�}2�S`u��-t +��g��u��H�
�y}����:���`��Hf��ɤ;��ʾ���\�S��v���xx�˭,�Z��L�|�$R(G�� �
�O�<����ճ�MAo���C)˘��+f�c��;ԯ�p*p�cf 1�!M��
�.�'T�"&�j�d�!��bz�y��E�4�7���O�v�E����-��� ǏLB�}N�X�X�&(��==�2v'P��gU��G�Ϭ��l�1mW�O��{ta>ۦ�-��5Hq;l�I�"s���v�9u<���0re�CO��t
�ݐb�N Cs�l�2!3iD:F���Gm2�m�)6���GB�SJ���z��D���a����
�t|:�A�P�`Τ�����e>-���OV���S�8� �V;vzc��R�;�ŝ�J�]i�϶+�f=[q��.��߽#�͠Uq����u�rUt
��w�0|�#�Wd�vn4@��&� s��:�y�^{�����%�����wdt$bJ��Sw�.v�J$tζ��1�S���fwp���%����qt"�`O-��,1}�9�F��#:�M�V{}pg˸%�����΃��2o��g{�V̖���-~YE�a��>fya�M�:n��䚦�*�)Ö�Cʘ6����P��j���0�
��1faٴ_S����o�d��Nv[�{t$�z�f�ٝE��l{i�7��6o5��5]8��U��U��ʩ�ֶ(L
^�y´G|�Q7R."����ɵ!ET�7�r�ʞ'�^P�S8A:�ydVMC��:�:�}; *�`l�a��f��@�=Is�p\���E�9QLG(�Lr���}>���
\�G�*%�Q. �S1S�r�]îR5Q�S�kl�k�.�es��j�r:���z�=��ohlP2���P�
�׫!��Q����ou��"���Ŏ�Ս��d�By��V#G6z ͂�DEzP�sy�=.ܘ�8�9܅^;��s)HL
�������*M�;��-�9���DB�c&��F���0ou�S�j��Ξ�W���ʲ�c�
���B
o�C��VP�����V�����J���͋!p+MNR��%����b�I�L���j��`L���q/x���
�ׇ��+o�����ѧ;w�}�v3�OEl�p5}�>�������MC���\g������!0.�#2T%oj9\��)A��>Q�����/�S�18ٌ��Q�>G�d� u�Ӄ����L��o�����pQ�u�y�R�֧��AF�j�Z#x�B-4x�ϯh�l���o0T��0o���;.�g+��;�˸�o�JNz�d0GD��)��0����9;mQ��Vl��5J�`i$q��TgT�W�EvUj��әQ�xx 6�R�<��Q�����}������r+���>�0E��t:ƫ_{ե�1e:�;�3�Q�[��х�v;ɭ�m�����U�L����9���qb��i�s<���X�"G
un�Byky�.��}�\B���
�����ϱu��̀۷
]-��k!Y��ʻ�x�y�˞F��q%�>�{�����]Ym�QU
[�ٵ ��|��:��ylƭbw*C)E��%��^	���!��L@��p�5*,�����O�F�9&�ɍW��חS���qAueNŅ���tS�).&@���![$��L\[]�f��o�-���v�aC
��9s�.*���N����T`������"6R�5��w(��/3Nż�95���JT�]����Vz硐�_��dh�ಞ�IT��VԜwt�o a��z:�z��m�
��:6��(}au�<��V����zx�uY���D���7�743��yCe���������`�I�.
��L6�X�Uo$s��[M���{`LQG4�߆��>�ɮ��V���,����D�z����l��=�LY�"���Z�����N�-u*Գټl5u�a�,�=���^��ƶ�^�Ru����U��{�k:7	���E)6�u��h�i2��*`�WF
��M$���f�n�����+8�vU(�v��|34h�cyLM-����ZM��[.���
���S��t5�c-��n������#�u�M�stv���U�C�\�v(&n�N�s�J���(r�g�YͥF��z�b钁�^x��m�T̖Ŕ,8�P��2P�m�����?d��a��/M,��a[��n��j�6<��ո�q�l�L�{�r���0�6�%U����h��Dvf;B�2�MZyn�E��:�ǻ�M�9]ĭ,w��oz+����mvs���RM� �Vz�G��m<�ͪn�Υ���D�̮Q��尳e�R�Q���e�8���nr� n.B\�^c�V��`��_?��]��
�<&���O)+��)���`ȵ)�1VK���CS��<F��:`�w܅�h�D�ݥ�w����/����|4�]�Ӫ�2l]f�g˚�)M���х�g�B�\��ojU�����zx�1]�����3��IU�%3��J*��E���1|�{V��#
����o��d�a�r�ټ#+�9�Qe���kƘ���"a&l���]�)H��9[��qZ��$Q��E���R��c��9� �b`/��tN���#H�{G��w�ۖ>�L���(�:Vwuߐ���{i�S��Ӝ�b�x�-3�����jo:r�o9;з�
���*��o%��Xn4�µ*���{xt1Ij�ͤu�ڱ�h}�{�m�Ǆ0+3�sk��ʞ��r/]nm�/��Q�Y�9�j1G�a�s7t$_gv�Wi8x� ���>ʃ��I>�(+�1�4O���e��I�	ݚ&|��V�Ye��T;����5�����u\�tk�8���6��ٶT6�wF���r0!u7XӐk}^��_6��'F;^�4,��7U�dh�X؈{�*�a�k�xET��YKz2EДm���G����o�Î���.R](#��F��Siw.�@��ڛꂵ��&%k;7���v2�+�7��H�^�_��Զ�<�4p�!�5���N���˶��j`��.�Sx��8��۲i�i�̫��$�ٸ����8���i�d0��}ys\��U��鬫�����VI滦i��[����Ю��(���$V��ُ0}me���eIÍ_�1��3�]���Y0Ji��f�>�q�Y��EGQ�9=�����`�o>2�<\'8b�olu�J�\R�__$�k�ǫCN����v��K�
�)Qf���ۛMS[\/���*D�(!'�����Ɍ2�Wp�*���{y�!���}�\ ��D
   (�b
*1���EA��,I���Z1Q�A1[K�EAUDEkEEQ�*
0b*�

�U��,Y �TD`��DVDUE�6�b��D`���"�PAVUQQ�E��Q��EU"�cX��c��%�
�����DH�U�U�DA�D��b("�QH�(���`�(��"���0Q`�b,XE�F(�h�m"�PUQ����A�"�*�U"�2E�T�"(�"*�+��Q�1b"�+*1 Ȉ)#�V�(�
,��
��Ƞ�`�EAb1,DEE
��b��"(
�����mUQQ� �"�DED)�UTQ"��UD������TQ`�
"(�*֣
*��,Y1��"�TUb��Ȁ�g����x�ָm/��v\��r�2sk�*�9\T���c�{˯5s@��#��;V 9I�p�_waIPUj3�119��W�� '7�T�[Q+D_�3�Z�E�� vXG���>�^�HP+*���W�p/w�sVgKF�X~�����FN��	��FˋkN���5[K�+��w�v�I��݅��w�j��NP����ӟ���7�v2�>����846-�A�e�f�M�ti�ݪ��㱱~�ݎΣȨA�y*�wʝ�X�&��3�����v�C��W�I>�IyL�a�ї��TQ�z,a�#v[���4���v����#�I�8㶌�X�Y�.�=���2�E{��.G�7�a^Mx�B;r�C��L@>����E�(V�5StUN�>))�����(��>*&,����\F�\����>�0��ۖ����82޾Sz2�jÂ�=�@�C���v�_���mWN����
��w�ؖ�+��\�7�F��Ir�kŜV�GZd[��;�I�7P�á:!@ۘ[\!�D=�x�����[~?��][���JF�>���T7N�'�cW��|�ñfx��-���0�wѫ���լ�ȳ��v�;�
`xP�!k�������*EP����𡽌v z�8P�`�1/L���޹xg����e-��i�e���g�.�M[��)��+�Ӱ���fˡ"]�Ad��S;�.O�{���-��:�s]�}C1.���A��C^�ҍ`�J�wau�G����oR#�b�Q�9\�b�&^�WA�GH*��2n��cMpϭ�񺆰>�*���O�=��B������ӵG��Ԙ��D��!�b0:TLA���o�ֹ�d�
S�.����Ҭ�W��c��./���>�y�"5^ p�����T�uW����]cob�]D� V�r��P܄w&��}C�\|%��`'���k���W"�^����Q���5LV�ru7n����F�@c�C��+�*f6o�}�A���Hh�7��D�tZ\��(�`�dP��~�e��m��M�>�\��Jo?V�ޥM�s���QE�����%\#���U$#[܃�|n����0��M�7YuPq"D����l�++�IM�d�/ɜ�#�Z6���n�0DG>����P�C/���c�"��Zw/y��n'X0^yV����/�z����"T�ӰԤlW@k/���,r���L��ܢV��%���۝�=I,\0��mlv^�ìz*����޵[y䢞[�Z땴|?4�\�$��ծ?m���]��AO�7���]ui]ˋ����^�8<�z��C�Swx�}|.�{�|��nmN� �;���v�@���8���_ < Y�T7x�:F��!�9P�����������������gb�e۬2���/X�&ɹ�a.͖�߮�#o�sC6���=} v*�0�`V��`��B�%LӮ��
z����3܅��%��e������ZpV�ұ%a`��`_��l��GL����4ޛ�˸,�~�)Ut`�Sql�B�½�>�S���Nf8���R�S)\	�)��j��맺���d1�
ޠ�a����#PO_�eY�k��Տz����X�T�ܭ��C�$��g0h���j�#t��q$	�U�d'U�'@�@�=���llpy�|geg.�}��"�P�H�_��l)pb�(��`�8>�a�3[���}�N*�+"�c*�+
ZZ;�Hhm8�gvC�S����`N��=��B8���
���9�"Lt��$�{.�' [�=�./�'��وfOH�=<�	C�����?* 6�Z}���h\�)�w��n��>)<5�T���;O���=���N"'D�X�`�r�ř����$�`h.��V}��{xs�	M
]ׄ��X�oOd�geN������]�r�t���Bd�~/oU��t�3!��Д��)olz&��7��IZ5���)ֶ姞ݹm�	�ۤ��7��&r<��ͽowK��#��Hb�  ����w�턢��:�ih���� �����x>4��67(��hlVA�* ��[yo��X��+r"~H�(ԗ¦	��y͉��C��n7�'��j��
��D�W4��k0LXa���J�sPm�"���F>cK�53Ǳ�GF�a�P��f�X�]��r�ڮ�
�v�U8{�����7T8`����/��?>�M�Ő�	�FT����x^y���Bx5�]HWL9#'�7�7"�v+�)���.K���B��%���=A�ϭ]�.�_�4a��¼����b����U�J�Z4��n��qb��\yqn�Vʝ����e��8�A���R2��0�xm!�����e�/,�y���^f�C��v�OU�;{�i҉!�>�>�o����ql��U
[��ͩ��s�^�̩�Y�zrz����-�� ��E��Kg������C�+d� ��&�E�/�G�̭��0���tU<A�(��.W`dt.���X�̠��).$�K��-1
� c��%e�Y<�*���e�Spwd����g��gS�f����P����]}�v��p�����{�Ѯ��,������.!���6�R/K����g[��Z����5s��Q���/�gj�1p��:*3Iu��u��[QL�V�.��U'MQG�����>��������k���ldZ�y�s�./�F�T�'�ٝZ��>��~��F=�Y��;�d�y����%�	bT���{*�8�ߺ�:��n��y��r�H�5��&Ѹ�9y��3�5�Bcf�>n����>���G٫C�Pq;[5U�T�!��Zr� K��]8�(R�n��``�����`�I�	pT�za�&�:,g&��^dMڑ����� 67�j��x3��p��_����>�HP*f�ۑ�������ƒ������LL����¦5���sXo<�j����z�]�����aq�U�B.+�����ӟ�����Y��� ��"!2�}�DY���9�V^�.�
52v4�0�ر�9[u����:�{��n��BY�e^�P��܂�o��L^%�[�zp�r���35;x>��[=����m71z�R�Y��Jd9��}�h�[ޞ��<3��
:e�(�i|�.G�7�a]�����՚�B��ؖQV���l���X�m�uf��w-R�K]�5�g2"�肠\K�U*I���Δ�uDa�����v
�֌�ъyu��6<�Bm�%�����6���o�RŬ�K�5���T�F!=O�v�u��Q��r]|Dh&�WjܺG�����uf�J��m����OPݝ��2�R���ި3�;B�?@�nk`ڨs�|��gvD���2��<�LT���i�a�[ќp�g�8].4*�Uӣ��,�ꙋ�Vy�p��{�]�yR6)Op��G����.x:�K��n�K��"�B�X��3��.a�h�ռ�΁هU�Y���<�չ��̄�㾟q�ޱPCt�i����}�#����t�Uk�������1a��sJ0A;8k�z|kx�TX1�݆Wf��}��2����L���1F����u{��x�GH.��2d�#�(#d79�r6
�F�B2s8ؒ��ב����̍m�^�5�*$4('���Qu1sC��H�Z��b)�]Y؍j����^&�]F�g�@J��ŀ��֙�4z�����,�����բ��b"���H��Z�F<��Pp}�-ulV�#�K�G1YG��q"#a�L�2��ۂ�*��t���ÙYm5Q0_���=}j����A��@B�:�9��
�.�'B�dD�bdWU;*Ihd
�� ��Ct��(��S����T�[3@����H ͑,�	���v�Zq��DI>��K���r��5�E���:Y�a���c|��u�s��_+��Y
oD����2�Vы���&5����T�ݴ��.�po}�)���}�}T��-��w6>��B��'�n�0c����-�����LB�/�ث�X�U�n9���Ö�6ZU#�z_���If��.2.�{ ���s�F�6鹋l�
�9��r�8�W#'OrJL��o�6vK����ghh�U�f`�F��G�2\!jb��:n9�K��GV�EuD[�B�����]����;�����1���j�ΡU�d�������lLP������
!�PԈX��Н���_�]A���;�Q������׬�1��c���!��kU`��������#�V��J��]m�D�x��>�WQ�Gvn�g>ih��v`ʔ����<2�k���ZW�Һ׽0T��~(���y��ޡ�~�q~dRU]"�J� �g��R�1}�.�����H�Jmb��y��݊���aU�j��q�E��t^�����b�\A�nw�&ԅ	��Զ���R����������-�fj7֑�U��8�; *�`l�~d�ٕ"�����sj!�����+�=�����J.レtH�X;��9dw�@�8UG��Y'U�NJtP__�,���S2ĮZ�H9���T�x9�=�7Z`�瀍m�c1uk�uۗڟL03�����5qɸ^��Ƶ`��ʭ�IN�����������	)=?� ����}��_��o�\�|QQ%�bd��UA�yH�ۚ)ثi�8]�2�9�u�"ƍ� ���!١�z�=��-�����`�
�L�r���7B�s��������LH%�8O[�zF��<�
���c�=e����j������� ��A*�$�=���>.ϙ��n��b*� (�vܥ�;p�4���\��Dh�#�"�S�D�lۜrx]�Pa�R�j��a�	X{��Q��Ӿ�=L	wlz�����E�i���{�>)n�h�.�o�߼X�6
�0wf�4�W8���~r0BG!\��5�P������/�t���Zg��y�wjV�R�O�Psź f*bC�k�+��E����(�Ḓ1���Q����mZ�IS�ʹ�Y�t^-�`��"۰����Ô�������+~�qwK��f����̖O��*[I�3������������hZ	b�ib�=�Y��l,=Ou��Æ�ڄ���нJ�I�KV�1M�
�G3iZ/��Z���vkMs��^�@gK�-Ѥ�Ȯ�ڝ�2�+�մ�Ɲ`��MH�7�e�r��w`����z�V'WwC+M�d.��QE]b>�p����gU�d -x�МmfR�{�.�J_{��^�%��/S��2`|��]q���=�<����;*�Z���iU�A7*�\)w��L^�LR+e`�[V9R�/��� '�eД�X����8��N�cR�^{s��r�t���C�µ�T���E��Kg����tN!�'UJ��R��Xꅤt�ִ�*<��	]M;.����׌����ʝ���pͧ@�;���D��
(z���8��{��N#y��M��B��C�
8��(\�K�27g����g�������!Զ�gq>ٻ�.��FΚ�i�eE��-utu��s��a�jdh�D�/�)�x������.H�S3B@�Иٷ��ɸQQs�ٟ�.ul3�Z�2�u���S��~���Dn�梎P�� ��t�q �@�-������YE�*H�.
�N/"z|[��y�ږ�"�f"�R�	�y1s�h����qsG���8��F7���}��kq���D�7�j>����LɘٱF�S{���
ǘ}/l��>��-����;{@��Gz�g�'�'Y���ë9_'7�[3y��:�Q�)]Mm����̺�I&��L��Ub�����豎�%tb;+N�꼭��u�k
楉k��Y��&��B�6F۱9s�WZ%o6����-r�7!��+3�W�}�]�ʞ+��;q��V}G(12K>��¼~}�cs}*ח��~�~����~���nz�mK1 턇[��v;=�c�I��U��ܩ�E�$��e	�)u��>�Ǹ�6S��if���:�fh3�c/>���E�#lm71��"���zk��bq	N���*˾��8���3IE{H��FA���2��:}e|�z���k����2s�P-=z�U��NF��(��>|2��u��?:��WB|+l���T��#�A��	�}Pg��zƲ-��pD�=�����D���Q~C�����bDI�/����sM�jC�,F��~:�6OOl���V�GXL�sa��X��م.1⇎������\I˱*�rKAB1�&*�`
.����a`��=c�BSb;��=�*47N�\�w�K�G�MU�-HQ0W��P[Cҹ�%��8ppC^���X3���;��\�7~�T[�� ���[��]D'.gq��B��9������0�Cs�\����F���1�_�CA�U�wtV[��N�2��R#���3��Ηkh�.ڣk.��j �}������[�-���>�X:Z��mE05�pQ�.��N �o�8˛u{K`��:M���Ĳ���u�k9�=�	#��S�	aqr����]�f�6�J@r���I����G*�Ćd��Q0�t�hm��z/qq�6g��1Ij&��d��I�d�����Cu��d쎃��tڶC�.�T����
�Q�����f�\�9z;�5�o�*S�Ļm�1,�=0\�z/>��@v�/m&�H�*��ƃ����/�,�Ѩ%�]� y���l�5˫��Ʒ��\ZT��fD�P�J�l�I�c�H�����_�,uo�&���3����jj���*h=�jX��=��d=�����l..�v<s^�6�F�9Ic�5�H�P3�Z.7�l^�ۗo7�"rb�g�ˊla�.shyd�c�rc�F(֍� ��*}���#ft��̗Dv|��/4Z!e]!���DWp�	��:=W�5��n����K��"���/�-��F�D�(�ݧwdT�b��C��M�x^������PJ]goV�r|��h/��zu��@��!`�s>E)n=Օ����q4��@�{#�����ll����G�+˺[���2��-um(Ș�7�*'er"���) ����Վٴ�MIn�Jf�ۡA��G
ky�|�R�'��4;����ٸ���!�x]�v���y��]$V�6=7ҭ?�T!�Ш.m_i�����3��W7U;]�X��X�e�b�y������ R_B�U������u;��Zkh=�Ѭ�p�l励L{E5^��]�tVGm)N�<��ǒ�Wi��'4�X�!aV o{!�	Lw�v��5�Zh�.��gh��Yu2i�p����^���]
ԕ�,֫u���P�5��y���!�?
4�V�R�0�Ã/�K�J�R�*mQZ���a[rµN��bU��<��ړ3Y���]PvL�]8*���" �󡠭z�� �k�[Y�|�^o:��5�hl�
6˳����a���m����@w�om�0�=ϰ��ݠjTru`'b�9�J�s�λ{]�)�rY���}G$���\!в�o��5{�)5���e�,t��Eު������4R�l�o4��r��6#��3-6�5̪IL���>WB��v�lT� ޵˖ȱ��lٽ��n�EB��lhO� �b�[H_A��Ft9�gI>����=dn;)].N�(Y�걕�*=C@�YÇ�������d������d�If��T��g1X"o:�[О�YZ6�������	�Dj��z�9�{��nt�˒l�����;\�.�L��U�8T���WV�[�K�5��LC*l3;�FE2�ه����fw�wo���'N���p�P�@Tc�
�ER()� ��"�TH���"��EE�EUPF,"�1A�U��QTEX�Bڋ,���E"���`������#"�QU��PEEPm*�"���$PF#DDX��F�b�b(ň�DV ��b�E�F0UV"���(���+R(�PDb�E��VF0��h�E�"
(�0PDEDQV,���PUPQV*��Q`1����1EH�X6�b��`���"����V,QQU����)(��X�b�b�U"1��A�UF)E��ȱA��X�F*�
D1��(ċAQQ��b1UQTDUX������X�AEPH�`�1�(���Y �(�QJ؃b ���QQDTb�1ADUPQb�TQ��@X,U�����*�Z��?�b��T}[dQ�3(��t�R�*.ʎ�A�cbnͣŝ�Ճ1;�/l/;*n<1��Q>k1�<���xxN�Ds�i�t.3�G�!`L��9����(�[<U�GT��v׉�Z�u���Ձ�F���v�C�ܰ��_�����ŀ��֙���T��P|���:��ˍ7x��2��VJ-f��34S�gc�h���n��}\X��ň#����ո�a�k;6�Dl̃���j�Ԝ�W<��d͗���P��+�Uj���\3���+���(�̭V��C��r�ؙ���"c �'��v�E��ʃ{E��Ӑc��1
���b��(b}&�k�y$��йHH���zX��x���`�Ƙ��N8��r�1�1���E���c���<�,�cv�Đ-��0l>92CB(q�:U� ŊF�t=�aƺ�;.Wo�ԛ��y�.sj���C���a�#cc5��v������b%O��4E���o^����^Cj-s��2*�$l��(jAV;	��;�>�E ���Ŷ,�E��b��y{v������`˃\�b������m�z� �U�x	U�+�=f�QS�(�{->��5[+�;C�gI`Y^x�g�/�*���:d����Ǡ�$���V*����u����I6�}"]ُF��t[�y+����3k�6wQ<{:����J\nj�ŏz��k���c��9Af�d�]l�"�F��{ә����������B�O#F0h]�&TmϔvMt��R�%aKg A�8��;���+AV�m�Sѵ!lHS+�V��"��}�h��+�=������g-V�;���x^4#�]A��c�
�Y�t㌋��+ؽA��
�%Dl�`�nr
��J��N*�rάEwwR�=Q��>u��*z �j�n�c�q$	�P�`i��ok	�Kt���sG���3g�_1Z=���қ���?{���B�utJB�1�°�ܣebO2�;y�FKn�XR��.;��CL�6z;�������P�b98��r'R=��k���C��
ār���U��3=``�`����]�8������^f���3�|� �9C<YH䅂�#"����&��N�Xꈦ�Ø�-Xz/3�;��N [��mTF���"����D�lۜ �@�.Ѩ0�&��x(�^"3���8�[��U���)�2�(ԗ¦�\��I��n��u�����AT�.�+�4����o�]
U�"�$`�zѻF���9!�y%M����D��q�ưǃz��q� �v:��:T{���ٌwmlS�&����ʹK���]k�grp�m�!]s����0PL�@2idua����1���9Z��� Sű�W_Zh�&?Ed���C�J�sPm�"��G�A�3����|��S���do*�r�Nq���UQ�q���#B�dy+�ᨻݝ��E��I���a��q�n��>KRHj�cNɼ ��"��Q� ^xe �#a2�ʑpWM���p=���"�'���������z�J�R�g��-��Ϭ�����X��Z��Ǻ�*6��Y���{���L���U�s�+��L��d�#�k�t��������;!ZӐ��=P:-Cc��E�*VY�Z��M��j�,�V�:2���(����}���budA�}Yle�z�B"���T���F�\��ېuэ������.xKg��1�5�u�l��
���ٯ�g#�Ws���[�H��[L�:���K�*v,-g�tSQN'}. B�9�̱������KBQ��0���*�Q}l���t���G*p��xf���)��g�֗�R�纤�_�VP����T���q˿utu�˞�C9~��;38K7��樚tØ�`��"8�m�����x:7�������~�Xt]b�,V���,�U�V�.�<��uE��_΋�t<����_A�H�y+|H*��;;N�\��̬��^��]ͪO�S|T��}�P���k(ȱ��-�"�Fb���Q��"2h\�0D�76#���̶4P���"�-fK�*ggx,��+qW�V��S��:�T�A� T��vS4u�W���¼���_�(�n�rw�^�U]��"_qB�L�Ɉ�$	�4\]��;,�_f�i���S�i
�����k>�<�
%���j"@r;�1��,���.�/����q| �gX(�ez�t�d	:t�<�n^K�;?/����Y%��b�N|B|cd�d]LJEE��l�+�J���R�(�ط���9���Sdo���9Jr�f��z�ے`!�K�5��q�0��ʡ$jFߝx̪�ػ�O�(�z2���~ <�U�`�x�Y������|����֮���g�##fR�� ���uM��P첾~=C{��}�Ϲ�x���~Cz�:�e��1 �EE�U����3�k�D�k7�g�U(p���ɕ0�k!a��줤����g�C�cY�!�z^�S��tWXn�K�Jw��e ﲽA��S���*�>�^O����z=b�_ݝ�`fge��BVh���\Mu�����z�i�O#�]�Bv������e!�G�Ȟw�5yS���)ev2�d$�(`��B��Et���l���� ��k4��"��"��;7���-n��{霋	p6+�z/d��ϩh�jdu�ȷ6��%^�}��;�\��]g3yܻ��cH�!ؚ�Ƀ� W�WA�Ga.{����؎�}��z�Da2U��V��g+��H�˹�c���#W��خ�ODm�iF \�(7!��5�<}*,\D�C$��y�޳�M��
�j�	@ә#�A�*:i�-̥<�J���jǼG�*�R�<��w��{D/Q���'�O����"�@�Fq������:g-�h����i�R�JḨ��}Q�ܸ�D��n��p��T��P�Ӑ��4�^��
y�xow�(��T)�.=�d8ܘ�n�����x�qb�+"(��Ĉ��+oh��y��o,��w��d;t�|��~u��zu�
��W�5'�u��|-�%_�kYi�k��iE�ߐ��@M7U�N�?�B��_As�z>j~�l1��9�훵�����֔:[*�p�N8��L����.,/���{�/@ݾ�������V��`�cŔ��ʲ���g	2�F�;�&��9��qֻ���c�kުH�'DSآ�<�2/q��y*좻 `ޮ�G�rB���u"����pQ=����^
�����K�m���f����\�(���Cv胥�;��ֻj�Kv��ڹ��; ��O���0l>92ZC��tUn�1b���B����z@�{�8�u8���"� ��q
ʼ�m�5��y[��v7܃J��ӰЗI��Y��w��J+W�5~�D�!������jF�X�l`N�A�}~��Vb�b�\\����Yp���je�~2�����x���𐂚͠z�_G�v*�9*�s��hq��R�j�Ԣ7"a���T��]z82�Z/�Z\ ���Zzr��w
�&B�5���L�[תݷ����>l#�aH@*��]*Ȃ-��z���{��Hw��
]�־�f7i���姱V	t㌅�n/PD6���H�������K��d۔��R��pɧ�{�qʞ�A��ZTiWy�8�; *��d+�=��K��eͭ���{����C��T�:���*�9�G\���pͩpb�C`�8��q��-�O^I"��h
��4��]îR,h�p�ݐ����=M���eW�VE`ÌuNɬ�վSSZ΀��s����88�걦Sbq.��hU��tK!I�وP|y��Wl�5 &���S��Q;1��җ�2�rfǶf��llZ�~ؑ�Di�5��r��&�W`��3V3-;=��#�cxv�N̩�1�z�T����ښ'�l`�z��V�ʬl5Pӷ�R��&��b!����S.�}S�3��'0v�KNI�6�D�""0J�H���]ib���v�>��zj{�M��1D����戤�MmT�<�KOhH���u�h��B�<n��J�惠����Z6N��V�{��6
��1aTB���D��sjH|*`��󓛲c�_n���盥�훝^�G��^�B�l�Rb⡈�����r(�5-�"��G�A�3������s<���W^�鳍s�\��=}�}�!�n���
!��8 j.�g}/�Qxn
��r��}.�5����|���:�EWW\ރ[�۰���@�A�'a`p���I1��B:S��7��B��3��
�9�9:�o��W�[{������ZFn�s�Bז�:���"�#rs%�t����e�P;B �M��7#=R2���-T9�e5d.�[Oq���=ٌ�BC}^e�n�Y-z$tmm_�*Q%�>�� "=x,��Wv�����D��	2�g8�r!;�LL��嗀��Ġ�'�e�YV,
��Tr 3�Tsz��ᨲek6c�Q�v���M@�k/q��E~J��mﴕs�Ȼ͵�{���Gy�������
6�Ь���3 Sd4�V����Ȭ�qn^n�~��2�ٶ�SRo߃ʌ��`���m��Ԃ�(�8%��^3@ba[& ��=�ٽ���}ΨX�u=���}e��`�S� dtP]YS��ՙ���Iq0��i7�r*�ެ���k�T�c��# ����bB��Gk��P�N�rL����	��>�����-t�B8F������.߮�T���D!���d�D�Q��{*	�/����s��1Pڠc0JZ�YZ«�-���{$E%S�lW�
��xH����}�W�mc���2�k���]�w9<�(&i:�р���͕N$H7WӰ2�2hdTt-�@�[n�9���W�' ����G�EWqb��Ɉ#��5拋�@�8�M�S������㓦��������8}��7�j>���LL����qSU�<�cݑ{u<��.�&_b�f��&��nc��c�VHB0d�,X�1
6%ϰ'�6I��#A�Uն�]�ӽٴؽ
��DTPފڒ46-�'cH�*62�#7S*�,ux���f����N�<�-=y�����*Zbn�� ]�=���Y�����;U�m��U�%�]	;-<nPԸPI���{V0+������p�ᾇ<7c�֮U��$��otm��ZMaɋ�����E�E/��c=g�F���7T�\��Vg5-����v�%�M*��Q�rj
t.d�p�6���f���� �T�Pޫg��]�2��s����y�"�雂�]�v�G�##ft���ρ#��ɨZ2k�o$V�6�V���[�"�U�O��REE�U����3�ϊ�"l\��Pg���̼=]o`P=	�9����*y��(7�
|}��K�@�nÃ/F��#b��v�^
P�3���_Vk9�+qo4�%B�8>C�xV�O��D�����������,y��Vݬ�|�Ta��B=4�:r6�莉���T�����d%unz�����w���6�(t�������t�����T�i��0uz�@6+�;D�F�ҌE��{J5�<}l,�8���p*���hjjOB]�B~��j�	@n���A�*:C�苜l��AB��U����m�;y����QZ��A����B��ǈ�J$<U�Gz�.ru���5Ed�Yd��C3���9���JNe(��Ϫ��7.,:'_�6x�Jj�>_@p�y��]��fK����s)�:7�f;g�#���}�����Ơ��٦��:���JM�q+Bm�A�s�%=�H��G��f���*��� ����1��F���r���<��Ŧ����ͦ����eX�B���:�ا9![wu�t���LE5_D���H������Q�Oƣf�2*��{F���"&[�Ȯň�R���VDV��B����ܮ���o��#^J�����eEA��`�ӹ����Q����t7�b/�{��}���V� ��!���ȷ�슻G"�;*���X��1貖��7�M�Un���P��[���X�P鰘�jLp�U{\�!����E]���nvn7CqT8ơ��qs���SՐ�Ađl�Iڡ>��e��fb|�������6��QcV=���~f�@#%C�.!�7�荍��uM<����9a�T�؈��:si��r�C���\��p�\Z�s�GOC�V;�����?[������|}ӏK�w��7�X�1q�(2:�$ ��h���b�R����g'�sW�^�=�����!`G�P��X��h�*�1͌�P��m��h\EzG��F��zL�N��u�S�r�BQ#�[[ȊB���)VD[=С���Dǫ��e"|�X�3v��*�{l�4�t�l4�ZξҊ;���!�w������%�P�6�8��s����&W��EՁ�5�I�۬���SG�]�viu�k���x{�x��j�`n��|79.����-.�B̖&kַ7��y��s�c���I\,��kp1��xcXtD��]v�x���n�4
�U�2k��|8.��vLj�:e؎�8U�\X�h����[m��]������G����--1��N:Ӵ���8�s*Vؠ��2]�^n����Ýv5��5���E��Wʴ�xp���U��C9�۷]R�Z��y����_q�e�x1�r�@��.p��J�oVi��.ڡY���T��y@��N�*��DY(E5#�/z�=:�Ԕ�iД8f�N��ivk���1v#�B���n��["[Ѯ�K�d���y��R�c�J��u��m�d��r���q�Y��ؖ� �C��Pǻn��3p OE"!���fa��;qU�u	ۆڳ"���w4�w���7T�]��_v��U�sҗ^	4��3B�:��+f����ڷi�74���k��f�I�m;��Xn�B�mm�ZE,��X��]wl�p����D,�_/��uˇ\<	�ձq�76��%�Kb��5/d)·q�eY��m�wqA��t�giY�ؤ�.���L#�+�rX/ot��ѩ����o�r��^7(��ň哥i��Sk��M ��ssg�����d�J�溬���	�VQ�<�7�"�*���l�Qt7)���!�v��)Hf��f�bŬ�"����b�V��gc�ׂw�`�K�S�R�3p� ���:Fղ/��o�CU9�cTkA�R��\��6m�zD�<�!$���2�u,�x��s\ỗ�w��|gFv�ʔq�R�N�7H�F��1�\�9s�\[��V�WÌ���b�fFjv3E�w�E�EK���]t���YΚ���p�w�A���cU���d��c�n����Vz�֞[���f���ؕF�u��|��ɒ�ک�i�r��ޡ�C�e�_&1����+^Qrw���J"��U�Ҿi�k��Z�Q�WW	��d��eڀ	Y��^v������&���ZZ�s��ש�T���2c�(���yen-��F�7�i7�� ��Q�f������`���kX����(
�[�m�:ɍ4�v��o\�䘺���64k>/@ER���x-��}��j� Gfj�=�Z��u���V�"[%�.y���T`c��C���-��N���`O4U��m�!8����:s�)u�9u��� _É���v�O��C4)�C/�VՆ
C��^���Ȭ<
]�!ݙ����Tza{be�V���5���W�cWc�3�%�j>��ڭ�%�z�i+d�n���iq���@���x��~�����dR(#UTb��+`�@X*�#DUUETU�����$H�E�(Ȣ"
��EekQUUF"��"(�"��`��KE���*,Q���#j��
(�Db���TFEc,��Q�UV,A�����*1�V"�`��
*
*�b*��V
��1TX*"�`�b�F*�#"��*�TP����UAU�(((1Q��Q����TX�ED�0X���TAV"��,A�Tc�`����"�*�Rڪ
��PEDER�*��PX���"�c"*�Q���ETQb�H�ҬX,V
1U���E�U�*,����lTUET��U��UU�"�" ��TTTH+(��TQ���Q���>z������sOm����p��\;��ѣ��;Ӥ��y6���79�2�����v�WJ�ڋ�q�e�賛�9LG��ޚ>ǟ�7�Ṙ���ث�q�E��/PE�x���H�q����ǻ����OJ���C�&��}Ը�O_�sPm#t�̸��+F�[<g��íO^uwũEU��*�(ä��9띀U�r����3�\�}⊉꽖U��w�y�b���`Q
HET��N.�!�)�i��ݐ�d�-�Bf�Fe�e�!�jk.��y�\u��ؘ��J,5���**�eŁ���0��]i���(�*Zr�P�=�sQDP-�ۭ�3NDD!(F� M'f��ª��;O��Z�=3t9ݠ�69�)��ǭa��T������Y��R.��u�h�,3�ٱJ�]�Q�;��W$��S�2J�X��UH�J^�B��bw'ɐ2�(ԝa���{�(��pR�:�e��hQ��}��K
r]Srcb���0w�B�%E9�"�*)��`|�Ϝs|yW���}�,�5"��Z�vez�] a�P�P�G���vv_H�E+GM��:���'s���f-��g�R9�k7��{�i�n���ɣ8��*ʂ��UG�ީ�r�oK
M��tMM&�V�a�ݢk7���b�x;Z���BwvxK�T�0��~�f�T��j�8�k�Kbqw�4�?HB�w����n������6S���y��k>9TjHg�d��6�
;�)''a"��jr��^�8��T���9w�t������QQg"�b�f٠c�z+ɭ��l�-�ON�y����3x,y��4��Y\\\�9ݜJ�����y�P8��=�婋��Վ��:���(vה��ϣT\��@�:�̄ݸYL���#�kk�����}�W�@Dz�GvfX���TNvR���Љ1����[�6���m�.�'*���xˈ���C�-�fG8D�����Z� ̐��;�zx�2T�t:9ueNŭg�	�1Lk�O�N�g��sց��r�lW�1� a�GV�g����ݞR�*�ʧ�#�G[�2�eU�XO��>��~�B(�'D&��/�:�*���.ո��2&��޸ᗉt:��a�+�F�!e=�"�Fb�*6q��^�P`�Ss�]�R�`�[�����s�@tM�b��:�	��t����PS��*�Ӑ4VZ�z�e�`ܮo��Z�_�B����Z�90E7nՄM�,(:w���1g���6�ɶs��Q��FзW[�4�6�;�뤰���V7xu�]���8�6�"�g;�[ë
�<�~���K��ʼ0��X#g�r��3N��b`=vt�Ǥ�N��)���.M�=0��Tqb�fLA�1@KT�Nx�{+��ޔv޵S+�M�
�{=�W�Y��8��GHp(�%���j"@r;�0G&cf�����k����0)Lt�9�;��n3}��lc5��e"�K�/x�(;4��n5o��.�k-{���+[�u��
��b/�V	�^U]�%�zVަ>W&sNy`ͧ��l%g�m��c�ulB}Vi�A�UB_���N_2yZ�%�7�	��D�k�e�+��=������r�Fb��)�~K�([��)&lFF��Q^��9gߎQ���޴���7u��G5~~yX#rTC���I�<��Me>�����9��rPعVVf�������fR����Q�wjaϷB�zȷa��=�@�C��۵NIq�f]	7jj>㴯���HX��W�V������P���蕅����Da�#��\�]P�.y���Z�.�E���j��ڧռb�Ez�0�á<!pQ�0}T�
���>��w��]_ҹ�Js �����Jn#����5`�=T=(�*Ț��MKtG������:�J�t|;���Bèn����A�Z;3{Ɵ���P���zv��awg����	�펐&�#�;�2�^k��6��Y�fRΜ���p���m�t�`.]~�3S�ay�܅�1F}�=V*��4�WD�{W��خ����
�tC�����?Ivz����\�����P�-�
��ȵ*���9�~��Tt���#&�["�g�����]�F�
+D�ǻ^�_���79r6
��7n;7ƅ�1ɏJ�H-��`t��{M���Y9�+�F=���8����۟S�*Nr"�љN-��=ˋ���l�<�>h*{��G���7:,����
��P�/K��h(#&*[��`�W#��K�&+�ƣ7�P��ݬ��7�BQ���E`��g����_��l�Nm;�F�@B���v�};K-�-m�Ë�=��A�Z����W�i��W�Q�o<O�(]��~�eA���e�N��Bѥr�fqִ�Ty��*����E��]�T�ch|�x<G���J�����Fn�v/��nx+���i�g:j��nb���U}l�m\[Us-���xGE*�1�(����\�����7�+5�7�1 ��Aͥ�����SD<;@l��,��\d��[KE��F���9�[��A�j�g�XSnt/� �ի�����\�[�Rmk�s3��n��E�?\����E��-��%�P�������Y;�]�ּJ+ߌ���CY�g0�=*�]�6��ϖ�	z���#]�R�޽�탒�CR��X�U��uC�6B�F�5 ��ccvzS�5��6�`�Scp�n#=�.,sv,2���xP`��b���!5�@��e��:���Lzм�IûR:�=�M�Kgzh!��ιR�=昺Ĵ_��K������	��c�Y�z��c]��[hc\���n�<�B�)��-�]
�������E��O=��4s�T��N0ϼ3�(�b��|����:�9����X%ӎ2-H���l�R�ɱ�W���G��X�m�WQ�����^��o G�K�T���hX��X�I����xF�Ei.���I��벗����h$B��zK�s���Y9�:�Ϫ���q�aV"�ꆽJb��j���y`�j#���6�ɪ�pw�딋Ѵ��0ףU��~�ѽD��Ah��ɨJ�}�e\�JFE.LERAk�2�4��A���G_, yc�𦻪x;i��9��N�h!�u`��=f����� �f�� ���;O����м���b�CV՞s�v����,���޼	we����$DH(��+��5"�	<��5���0ʁ�Xmx�hY�ȱZtaO$����
G��%���Ei���g7B,ݬ�����$RѮ�TB�ڕЗ�ύ��"�WYsЋ��]V�"�$@EM1�|�#EI�L��KE`!a�(AVO�8��~��z�t�
UC�HȘjwr�1~�TC���D�&@�<�e��1[�Nk�Y�0eS�ٍDa����⧠1Sy&��˪NLh��"�C���B�QNj-�N�}�qZò��&���i����Pu\��:�g��a���#BQ���5S9�-ME;�[�Q8��$�"L�aQ�F�>!�RB<{&�����Qu _U����\s�l��hz� #������p���M����ƮHU�i5¬?�s{r�ٰ����=�k1�t����!۬�Qs8�vq�JL�������]u�R2��v��XZ�{���Q�w`n��������U��S+e��[WʔI�ߥ]vztj�ew���	M����j��6ϊ�r��ͩڨ��Z]H)ҋx��g�e�ė0ͬ�����ӱ�T��.	�1 "$T��}] �V@�_�������v�p���X�KJ��H�^k^����A2�h��eu_pU�}J�C]Z���on�'T�,��J��ī3j�AK�R�<���6s]�
V"�ֹW���v&��\vG]ܗ�Z��2�ͥ���ȹ�x-3�������o����B�{�.��C��Ռ���W��^��)1�.��%�+��	��oB�'�����2�Q�86}W@a�Q��AA�<ѿr1�leN�͏��;���w�:�<����,��DX)�!�}V�F�<�k4�X���%��FE�p~������GC2������7PsgA�*�H�)F��v�ZS�L��6�:ȹ}�E\�sbS��ϸ�U��+0���R�+�����wK �{�q^�՗����:���S��l�u�;A@��[��5ϻ�0@��lޜ��r�[;s����a��EL
�.,Miݕ��71�����B��.X�7�B�t��K��d�\���Y�6I�݌�^���q[R@f�ż ��#0�ؼ-���Ƿj��z��y��M�-:�|���$����.d�Fگ��v���j��%�)et!�S|�(�盄F�☇�@#H�;	s�|��$͈�ٚ	E{O�2��p��jLI��3�}p?p��p������X��MB��w��Ct-�S�jd�A���e�@� N��;N;���o������x���ӎ̒q��Ms�������e,E�������W1�y���Kwe�2\�"�I��1�x��	l�E�d��]�k6�8�1�9�P*�����zX���Q`J��u5��=P�UIHּ7���.	)��
���x���A=t�6ه��!wWgl��8��Sb���Dd0Xm��J��=b��(.+c��O<v�?Cr��}�S�iE��系.��l&]	OX�V(ﾧϼOܜT�U3�c�+�jgm����t۩}ৣ�685<.j��M*��k(�O�v��l�Հwh%���"�2�q@c��Zp��9��g�\~��1�z����Aw�Ҭ��[��+B�hI@��sz�_��f�:Vo<�"� �Up��K1��Sͻ�y��}o2Űc�NR��oZQ9��V�m���l��X!��By�M9�&4B%	��KNN��49�������U�nh*������z�Ì;u7���t~̶`��<'3���=e)΢���q7lP][��r�O�3��g������iGv^��;u%��~0��!��&:M�K׊V�t�{Y��R�<ν`�]d��e�noE�s�ژp�z�'_ہ�;JGy�������n^h1�m��v�G�<0���4U憳Yo=W�v��*�����t��:�����I�;��t��SɌ�b��|"��٠nړ|����,�bΚ���y:��ڹ�{�Z���3�T��'CWЍ|:X���3���j0����KK�eQo�c4+5E+d%Ow �}T^lJ����Ҳ6,��ir("=��e3�-�A栶�F=ӳ�
]��%�K��f�UV�j+���l.��WR"�J�Ww���&�R�T�]�=S���&�������v*��'��}s�
��g�JD�L݃�/��t�G�u�~h���r�;�i(������J��,�PذS망u�����x1+��ڻ�ڜq{֮�v���/*��:Be�����Ϊƹ���"��d�v�]�����b4�8�96���}>�VRi�zk*[sa�Sz=�o�����z�ή�2h��xk3ws�#k����^R���@�r��vӺ_i�@�
�i��Y
��t��E���Y��W0��1��,rO3�q���K��#%H�E����z��I����7�tY��幕�8� �V���. :�Ҩv����;�V=��|r�s]>Ur�ݸ�XkVo3*�)8���V�������C�pcgۺ]��A�-��q�r0�o�;�)>��������I��������5㍑�i#�Nu�鼼Yy��|�UH%�7���(k"&��P�����',�s5�޵}J��z%�"��D)c�0M�"P�}[l�S6�Z֬����1��>UZ�QtFSze��b/��]Vk���x��sp::{a�N��U�_��x������H{�)�GU9"��屴򯳩��v�S1����Ӟu�onлxn�Í
Pi[�i�Tn\��2u�IM��7��E��`�y�3AWu�����B�؃P(j�/dx��py9���C���N���E�l.��WR���yn���]% �z���M���)v'l8)��*n�|2�"h��n0o���[Ses/o7w��[���ma��%�$R�+M�I�����vq�6��V9}�'A�԰(]hTo
�����Cy�z�X���Ǵ$��m��	I�*]�h�u/V=|�\�^+/i�k�4M��mc��1#���x�7��1c]��Z�psˤ�a���A�#/��\�Z�44������\�[b�M͢�Et[Vu������aX|�?>�/0��'-�J�8���N�n�VZ��W�Y�dJ4�#��v�{��tQ�O�����PX&kb��eM�JA^>Z�7W���ȁy5S禄��x"���PG�Y�$��@'�龺g���FL��Igu��qb�9U����+U����^�G7(<��F�;��)�^	|�Զ&�Y=��m4;��&�2��C(��Բ�ފΛ2+�2��A]����@ũ>���&Ve\i�WNt�x�T��9cxn^H$� �NeӰ\Y���UpM�ѹ�nʷ��=�|�sLt��7c�Y�͵�)�+y�N�����=ز��E�<��G[�ouk�Xۼ�U�G��0�I���]�*)�.%��X��]$�͒3y	�2��zp;�O��m<��z�R��:9��c�+;a�cm�)]"е:�ǈ�=C7+��N���ސf��Z�����B����Ɯ;77 ��`=j�n��n+d��E�{M9��wn��+����u�s��]��
��u���$\��X��E1�����*U��0��E^kb����ةmnn�:�9˵����#��"�\}�\��)���>��XJ��o
�o�X�Q
9�mf�-^��/+eL��{�a��[<���%3�*:�8�X��S ��xRn�=,�[C�޻}�jt����0�d�y�^J걄d��t(�A�*�r����򛚩P86�^Z �7��u~�ڭ/@T$�x��s�u�6�¹�J�3��J�]�Q�� mʾ����3r��o�΅���LX����익/�ls�7+%�c{u�D���,ٹ�I�.�0E�kef��R�4+��IbK��������)لwl4���.�!ً��K��S�s�w(#�۽�\�X���sqm<�2lKm���Re�y��{J%�����]�X�R�tG��N���<U�U(�+u�l�aU0p�&++��-u�E�T�Hk��o'��&Gg��hvb���°n��f�f��Q��p_s��x�R����HLA�j�]����x�ܕuqQR�}k�(�6L��ܛE���^�E<_g܇[�wh���:PZ�4FT��;��X��(����SV�/�/,#;���z�#/�q?V%��ū�j�Pv�ˡ���F\�0v�c�]��1i�m*=n��H���S�\,.��f�\y�������UEE���TB�V"��c�(,FEUX�EX,E��"(�"����(�"#���PX��DAb*1F"�b���UUb���`�b�2�b�AQX�b(��DQE���������1E����Ȋ��H�*0E���EPQ�J�cR���Ym�DS�ƥEQ�[V"�Db2�EUX�`��֪DUb���1QEEF��QA���F(�(�"
��2���DPQG-b��Q�V1���H����Tm�UX��=�������+�_$��Y/�z ,�T"�2���û��֋펆B1&"A/8G�\2oM�`�]���R=�N��Z؛�,�x�)#�4�+�9{^5�v�^ɦ���ug�Q��d��Eks�Gv�c��ϓmCV�}���EatÎ���"�����E,�m-[T�OX+�ń݁�q�t�s�ɫw�oi�Ss��≕P�-HT�,-#�up��Hg� Ȧ�.�q�C�	�:��)����:��Jש���\iۗ�ʅ���*�ڮ��;��Te�8�`N��B��N��MO-]��9D��!�1�կj7Z0�D�ջM��t�7��_(���8�L�U*��:
Ǵ%�l:��n;�n'0���������ֆg?C�}�)
��޹�oERp!�C�;ˬ����[�x�f���d��4p:X!�ù�|��<�	n���"��ۭ�V�DűL4bkme^U�4t�9M��{��;��=��(ON����EN��-���g�7�4-A���T�nd�P�r����%���(m�� e����E����f�{+��D���k�-��f���G�)��¬r�w�},����\��v�3��%��ʲ�#�;����bcI�)�ɹ��uj7��le)�I-��l60My�������*��l��C=���2u̢ܰ���K [��upڣ����f���x+v���t޼�/�=�T��w\�r�AR	���T�g*������yVm��e�X�$�WOmV1��Pr�ط���#J��Z��s��!��%��9"�B������E]�����+)�s�c��f��$����iR�=�7�,׸칾�Z� ���q�b{���L�e��0�Rp3#]=9�p-��ܤ�z��n)�\B�ˍp
��mM�utY�k�1��'�ln
pl^��u�ξ��U�=�M��ʻ�W�u}�|��}ڨ�}�e0[i���3��d>s�=��2�)�b��Up��V�Ι��ȎM��żZ�I�n�[^;������U#Cn+�Z��c{x͈���f���jp��
���)��xc�����/��9,��+m4S�3}RT���+�)�3���`��
KA�c��=��4���c��q������̱W7wOHr�d��x���aV5�킐2oLnWSʾ�� Z��dHE5n.YI�TM��y��*�Em8i���U��M����X�I@��eP�^Jn�մ��`��~�} ��!�у)�˰v�	�ۉ!�ꨞ��<|ufkW����*t*��P�:��7�en	l���	����of��ywHN�Ԕ��=a�bq��b'
�U�nh*���+}��o+��Z��K��H\�P��1�i�Mdz&��
��v�,�o��ڮ�T�V$v��Rcn�>�����Lo12�D��A��Z�����a\��8����t�߶����R�uS�|p�j�ЍC�Xs��Mfs)޾I,��7�ʯX}t�cC}��4��/3_��(�n5������#�w��_�>��¥�i3r�b��؃�Am&�l<�^�9�.���ZJv�5�����pV/K`�u��R���b���F�����Pі��$+�]H�yDǉwV2Fr��%!��W�q�r:G$<^�ŴD�p�-�cw`�7F
w	��.!��<�N���
��es�g�M�r�RzA�뤫�Ou���-��L��v���k�f�\�S�wo�S{�9�ۣ�j��U��LBǫ ��]a��vC�['���s����td��tF�ϣA,,/�Yx�H	k��~S�M��P���v
W���Yg���hu��`�z�K�5wN9��C{N����Mv�H$�e�o���ci�3�(�����n�'��tB�iS
�/�fC����Ru��]¸{غt[�����/]��gX�s��+��ly�2���F��5�kڌ�]V"}Q������;�.:�[���a�j�gAc�Ԝ
����n;.N)�q�:�7�N��g��wr�Ͱu���ab���z*S��P�}Yk(a�F�q��f��>B�Xl��K6���,a�1�Zuc�B:���d\��Ѝe�ό��6��Mˣ�ޙC��/�����a�P���5CUEvW�0�g���k��ժ���Yǩ<��hw��9��c�s��"�zev�0V4��A&!����̅H��K4��l͝s*M���On�E���ZP,�ӱ�PWK�ɻډm�C��h���wM���D��~]t�����=�-1�	��yW�v�����!��޴��s8Jթ��wF֪�V�YTӸ�#_��m�����Hf44aA����)��J0��������͢��b���3AWu����>�C7]NuQʙ�z���w9B��0�F�n�f�r�ì��PC�3���鱓��r���y-)�~y�O����R\�c���T��C��H�CIq�v�rإkwy�����nz�P|q�j,��P���G���+!���:;M��}�WcA*���E��nƕګuk�>M[��3��'��彗k4�FVOe��ȇC�*�a�Q�]�`���^��D�ADq�@��]���:��tBlӵ.+�Z�d#W��e�0�v9�l��Jnm�wS�R�-�XՀ������׵u��aI�/��Z����ѱyք������Oy�n\�B�y��Q�mR\=�n�y��i����}y�g.]�T�Dصj�Pbю��N�؃|^�;sR���n)��N��r��X$}1��9	��ӴQŌF�P7�53�������=�,E|�p�kޔ{�M��?h
���t,{BR���V���\X��4�m�6��}B��$C`�X>���]M�cOD�I�*P�CxB�l��[�vcY�R/��p��`t�	o�X�#�/4g��.����;�琅	�Ȧ+F���YW�m� t��otJ;����eB��㰮��5��1�bu�Oy��F�����l� e!`�]L<�WJ��u�W�fM����mQ�s^�V8��[��V�������ZH��]�XRJ��ڦ(aa�=R�E��E��>�.T�(@s���E�˗�ֹL�}�E�}����R�|��E<f�'s�9kO�n��Z���=Ԓ�����:R�u�� RH�BǺ���'pU1���;{��l?-snz�F�B�h��O���o���&o��U�"Pmz���8�}7ƻ��\��Ӗ�G,S�r�،�<�5�&m��8җ�)�$�k4?>��/���"zf��3B�t����S�s�5ծv]�B���(����]W9sn��m��!,xQ�opP���ޮ|��m�s�Ԃ��\�����C�_�'q��=��<��	�3a!��cQZutj\R��槢��J��#��2�P�;o"O
xV�5k_�i߀'���N����m�v�V/&���f��I��e�č����±�p�b`�gv���ܛH�m���v�]�QYT��#��f���^SD�O�� a��Ҭ�V����+�sbq��GmB�T��01��{ ��d=z0e,�O�ڡ<�`+���ӎ譹���Y�]"��8u�]xq��.�<f{{ۥ�،Χۣ�gTM���c�Џ�z�b¦�
������+h�ٿ;^f��tW�R������p��A���,N4"���t
��,,�!�wO_�Bo��b�zu��m�G)��LpW���91������^��,�fOB=������l�>��	mi���đ_�.qv�ƛ�(5��귵�BǢ�q��c�eKSŽ��H�$o}0j3���+����[��v��ж+cD�@\�m��t�erV��<�먳9�sx�./���1r�U��w{R���v��<Ѵ�al�3���}zM��	�7|�-�2l���K�B)���6+*�XE�F43P{J�*{�A3��E��He�Nn���6Z^���[�1�\������м�j
G���`�ќ؋�ۻ��}]~{�AX�!�p��6+�\��을㻹������w�yR�y��1ص`��]a�����C!��w�q[�sz{�n�0ғ�<�����#jĵ��>�V���aqT8,��ӞsӗYf��)�ż�s��@�(=]����}�����7���z�b���c�����F��{�����U��핪���wP�x���\�Ua-��.W]��{Υ\���l^��E�>�C�`����B���v`��:3N�v��-�/K禺�Pb��oέ{Q�u�X���7u/�(p�����V��M�����":����F��vK�%H�Ԏ$��D��a���[7����%N�Y�,���������9}H���2>�潾�g�!�_I�W���n7{�76�{5պ$9�m�^\�6\u�]����#(�s�}���=��뗕�A5��.@8�Ats1d<�Y��z��M�FH���u0�;7��8%f&��k=�,��&�Z�Ym�XY�G��t�h��L��
X�b��i���(U�ZٛY�Z�39.ు]k^P�sE�Y-��!��b8LfV��M�ﳺ��U�u�)Sb*�p�bwq�^P�Yr�h�C)��ذ̡JVekE�}`@��XÞ�)����{�4��y[�v��t�1�H,ˬ��ƹ|��t�K7��yZcU=���꧆1�zC�f���͊ʢ�T(�z�:Ff	���y���ְ<����b�Ѫ�l��о|%���ߎ��n{��7h����<ܪ+�c
�k*�
H�=�%J��P��u���n��e���w��-	0�v��Av�i���=����z�K܆H)�Q+ы��`��q��*us�n<���3-4��T����m5�p=�^����[޸�����te)�ۏh�m���q,/+Ⱥu�����,V�\�9rm	V4w�a�����yҍ��c�����n�����箌ˊؽU�r�ɺ�䷔EGń�t83�]��X�_P(&�J��GJ�<���ƾ���}�e௾�ևՔ{�մ�9衈rr8-U�!hI�Cb��|Q'w��GTۧ��x�]:V���٧j\P��B�Ћ���V�%Jl7�[����e6���׹cV��H�-����׵hZ0.��5��&1���s�L��0�{�6�����ZgA�4��{�H�qutĺq�̅5�u#�I?P�)�#>���L���é�a�`-=9�[��s-�en��;��$�bX���w;�sG
8#�[<&{�Y2�ּ��xpO �imd�HX�7Pע&��
��nh�Tr�>�(e`��ڽ�U�G;[01�`��a�	�6��bwq�^]����4>��E�4�KX�E��y������/�����s3����.s�ݯ��y9�)K��Գy�=h�݉^�j�sSݚ����+���#O��{��wUCR�j��K3����iITwy�,�F��m�" f�])����iL�ע�d-�9k|m��� ���@��X�cl|�1�����ڢ�kQwyj�ѭ��:���{�l��XV�mǁ�3�W�q�/"�M�j�7�m�
�ǀ^�໑��k��tU�CP�Q��Į���te:e'+Ge8z�n
�7n�]^0M�� �ۛLe�t�q�� �ז��C�1κ>�e�4*�E~]+���B�W;�+�9�_N�q�c6�iy���Ǟ����U��/�Hj��X޻����mX�$a��lS{I�\��_tda3@���
ʛ]r�ѳ����2��F$f](���n`�I�0	�N����(�e��Wc����ot]Ov�c�1M{u1lb�ȍ��΀���o#���!���z��p�WeJ�'/�{SwZz�Eѝ�Y��xǴo��#���No7uT*��������I��Zqؙ���SMGۜ����_[����D�@�ގ�;����u�j#&,�-zm�5�:��)�4�p髶3���]�j������C�X&��&�m񙵜;��Ƭ�yN�����ynk-�׳�j�-�X4QW3�+���:��1�1Md`+=��%��Y���-Ƕ�e�^k��Ѹ�w��tWל���\6:9{xi�����zU�Y[�ZN;�w����6T+/�iQ]aء�0�=S��U*-5.���A�$��(��R�9�e�G���Z�5�ŵ-��]���zq��.G�rx&��q�p�1L�[��Vͥ��Ψs�_p�h>kU�]6YbT!˘�[��7L�댖Ƹ���Π���[k0P�'�gVK�}2�Ef�$���\�jToR{�\ѫ9��T��ԫ������]��pʜr��`v�3�R4��RM���xw~�;����T�w��n,[�as{te��z��|tkyS
�]3%��)�N�.�z3�������+�����Cc6Rgo�l���X�����.�ӻA�X� "S������բN'���9���wzV2A�kE�ƫ��!�éQ/jʍP�X��m�}��K�;{4j�9����N�h�ͦ������ͣ,�Jm05��s.�Q�݋U�S����E�\��Gl��+�8.nf�[*��W�ò�.�lU��S2M}�s�sQe�8�A�t��+<w�"��]V���z11�Lq�Ga��"�M�Hu�Ţ�/�[���؂4�A�7���4"��\z�*�-�غQ���]h^�+�M{�b�᥽r9v�F�!�`��6�Ory�p!ET�{���L�5��BTN��O���Z�`/sZyԟ!��7k��t��$x�-�3Fm�yl��:�pT'l�L<:��ZFQ�=e[����zL�:Z�;�@7$�ڻ��{u����~�@iEU�UDU%DTDX��U��"
����cX�
E�,r�TAQLi���F*(�1b��X�����*���"2 �1�X**�DUb
���A�Em�UH������DQDb��h���*,�`�b��V	��(��Ȣ*��##V��DAX��E"�,X�DUU@m�kT��E*Kr�D�miQ�QeE�YX�mD��"�V(�bڢ5�6��#Z�ب�2�-`��V����绾��_��޾��ʈL�;%��D-�2P��ؚI�q�a��K+:6�񴵢Wj��N�=Ģ�bm��&��9�b�;�A�bݖ4aa��25S��g*��>�ˁ�p�1��y�Һ�ǭt���YE�ۦ3��"�����;�l��u��X��6�&�:*���VS>;@�8�A氷Ԓ>��t!�i؛�q�w��շ�i��pPNV�{`Tr.q��F����{��tH��`j����p����{��]��ڊ��#�o�8��E�x��/�Ni���
�=٬�Fu�>(�J8�5n���Qѡ��t%wd4��ǌU�����]g��il�ղړl}��~��]�~�8��t[f]�衋ɱ�=����H�kno��|�c�H�Ā8��ݤ�x����u��=��y�fokY����bߗ\0�5^��-���*�\�o����x����.s��%���Y��8��ֽ��F�$Cڱm�˰v��Rb@Ci���լ������Nc꽓�NK�+����X��-�$���ז5b�)���-�z��Mٛ��L�SH�d�ӣV�Ao,�Y���9O[��;dv�4�w��z�u�8��̷�ᚑ�<M*��z��+i�4u�j_J�kmA�܎��䠜oko(Jp��47�~׎7�d���Q)múWy�x��|�کH"���KNJ�N��Ksv��걂I����'z��*`<,��_�s�,a�1�i�Tȉ����l^ڡ"X��9Y}�T�� �t}t�ۤ7�(rc�*h>Z�S{ԏ=YGR�۝h��]�tf�ɶ.�.�9(U���v#�T���s��g���2�1s��v�gp��n̯݉��!�дJڳ(o�����_u����0������8^�4������x�0�F�M��%=�K�z��N�RX�s��WX{�AX���i�;1�sg8���|�����t�#�r�o�i��#���]m�W���G^:�p^��3gFa��hEks�B�Ƹ�Qd&ڿ	k�m]�m�)B�?�4	I�Y���������u�Yڷ�9�{�n5���>�����^xĹ�L�~g��ۀp�f�BI��.mncw����I��i{�)��xĬ���뎌~�Zv#Z�l*��7,t7;�MC) ��X�����4$�]����8��]����s0V^jIhB�S�D�"��c����մ18�}jὧnf#�r�VOTFYw7Q�V�0�c+ڇB�eX�y׍vu�۰��˲n��u��K}��Y���nh`*��</��Gj�{7mn'�so�m�]#�fn��j�?s\�ώQ*Ey����DN�	�H���.�Q�b�7f�M�\n�B=��m���]I��3�c���A�n;�uGt��k/�{��c��/}�S��h�x9�)�^��s]��Tfp��x�����d���p�1�8%�~�a/7�(��!�yK��Y�ݼ��|}]��zM׋SE�G)�6P���sy�i��d���us��-��i�B%�5���=W�we�Z2��-���,����W7w~���ٵ�y�گ����Hz6h:̷���p��˜���4R'WL�]��	����P@�(����y��Z�u=)ڠ��zl�j�i'�|Ġn���k\6eu�/�.;��&�W�Ks�te��WTebz�=��7���^>�3����GS��14�kgc�r�[<yR�ŕ�W\��T%s��U�a�����3�G�\Pl^�8i�� �l�`*u��Ζ��X0�N�k��ߤ\���h�����I�����-��s[I�Q�[�d_au.��-����f�)-��y�F��\��t*%��юr�!�}���x|s7��Q�<,��0�Ӟ2q�����V}��ǻ��v��n��F��]�8�/��g�]��ŬO�4U]u�jP�Bޝb�u�W��y(��W����*�2�W�u]��E�w5���m,����m��:V��f����憄C�e^K��|��Z���b޶��an��u��������d6��ǽ�7bkl]݅��w��7�[����x���kwJ�z[�3���4�{�����\h��}��G;~�"A�V�� `�G��v�{��z�נ�'�^u��oRGL��)5ay�X\%b��E��ytM\@'½zx��4���k���׋w�����;�ؚf�����iy��WS�����ɰk��DꗹϮ��� _>�Ƭ�f�Ӹh����C1��ǯhw5�	C�Պ^��^P��G����.�GD�Wӆ~�zt*ǂ�Iؚ����`��;�=�[<�L޴�l��4,KN#�7��Y꼫nh隶�h_C��p���y�c:��!�
B�91|ģ� ����0nzRqI�
�+�/�]S���ڪ`*u�������ch�3A���9��:ݷ��<�n`�Z*;���˫�]�t���
�	c>�NM��E���x��n�WH����y$���3�\��X�-�C7��^$�lk��9R.K���J���~�T��B��{�ج�}s�Z��/�+��Ʃ�i���-)˼��:��b��^��q�؏�v���q8�oo��v�־Ri��3����͆GoH���'�@��y��������(������5���K�k���CaPR4q�V��}p���p���lz��]����D��.����a�8�Hv[Wi�;99���l�Ο��W�:�lU����Zf�M�!1�X�÷�t ����]a�%;F�!Mb�UN���;O�e�md���]��c[���3au)���+�~�3V_�$ ���k�s���~4��>}8��8��Ym���w��X�0KX�%���傒4�#���Id�Z#!@���5I���*�%ժz���-�j׵��y&�78�-�t�y��%�������'��,MZ�YM4hj-{QA�n"a�X�����0l\F�O*7�fU[��j��#]`�����^�47�����4q��p�fӕ7XH+[������ v�<�P�����d�����Xc���-��y-��=}7ع��~l�>�:%�#��|��#��5�W��s"��2ŭl3�����ˌ��m�� ]:7M��Hpr/�rb󘩗s����Jk\��V��p�`��)�ǂ�(]�7M�!�[wb5Y����f�Ƨ��b�[���8�;��J#_�u�w9�xn��hn!�
Yx��p�,2�i�+i������k�V��M�ctTP/#��M}g����(�ԗv��9]ޯ,�n䎐��]���NQ�H�!�$�s=]���]d�0�Ő+7p����e"V��܁�*]Jr��vG�^T�w��ux8u]�s�S��dj��+K�;m;�z�i#o��w���6+,=h*�98�-Uw0�QFzbm>�H�T�7�3IPK�'}\����lI��N�mp��:��.�ƽܖԛo3q���6H*��{��~���W�t����o�ʊAר��;n�#�q�ë�/.�OBm�j�{��ˠ�U���U���6��pX�@U�"����Ú�}�մ18ҟZ��ul���F���om֮U�܅��c�!W"U���F�:�-�]Ɣu[ˣ��t�}��T�0L�ڭ]U�ˊ{P�5\0�T;V{�ݷ�o"�d˜}��v)E��%�X|r�ʑM(o�=kڏ�n�+G^+���{�J\R;I�1�ݭ��S}`&t�h^�4���g<�v�.K��,��w�)�����X��mW��P�g��}I�>\���B�Ӌ�xt)�n,��n#���+��{#;�h[7��;tlB;�̍$��%�2d��͎��I��*[[s��e�6C4�`A@q����U\�1�:������蚃{�v�������˽sui޹��!}��n�!�r��I]ꭚ���)�x�x�h�-�p��#�/!a{@�.V�����I��}{��B��kLhע&��I�-Mʣ��eeu�NZ�>�}�|�G�Y�>B��Mb7m�^]��De!��g&��J��x�S̛��\��*�5qO�Kѳ��H�}��<���^��Q�IA1�i*ڶ��XG�c:��:ʭ\!Y~Z��f����̋��n���9�[���C7���#t;�f�_Q6)(��Qݑ�Pm�ĆQOW>�u����8R���Z��V�	�K�������Jm^�*�������!�M
�6�fJ�>nݓf�.'��)]�:�}J���fV4�PvC��ʸ(�M]����ŞǩY���k�	Zj'Kk��m[�%ӱ@499�-���J���e�s&0K��u�f�4P��u��|5j�w�!����o�U`�]��Px�7�3����z.��vd�]�q�=�ژ�n�C[�$Nĭ�&�+���p^w#j��X8��3���:+g	8��^���G��-
n�l��9�T�	v�]�$`��j�\��-;�=^oj>�9���l�P
�p���uv�������kC�V����n��圱�/ZFAm�?"l���R�ol�������,e1�J$z��owiq�J���uc��igv����[5Zm6�\�׷�f���r�c�@���F"F�I�7sq}����&�H��T������2A؟U��ʱ�oB���EO;q4uo*�}�=���`�i�	CX�³�yBۚLĊV�^��ݰs��ci?%
��;��La��49�U45�����}=ū]M��9�.iuu1�C
`�
@��<�����>T8�Y��9�����ܺ�jb�@%���{{\+d%�T�.����.�]W��Q�|�ȡL�U�f�*�F7�hW�x3�m����7l����������bi��&=w��2�63Q9�QҲ��l���l�֣�m�u��W�β�<ëٗ%s����55�t]����/��y.u8����u`;�t����G��>3�YM����f5'����~"���n�O�v$%jQ�j�l|9�^s݆�YJ�i���u��9	�\ky���1�ѽ��9��y��Ɓ�=W�{���A���ئ��U�Fɛhλ�y��yӮi�[����>��a��8�Ʃ��9l�=|�Rm��7%m�%�qMc��}��)�¥#GA��-<�[o'j�7S��v�������������{�|��j:
�Y�����"�Ү���\���s�㈳�/Uc|�h%��-wJ��R�N�(��:TL����*��Nx]���G�z<�������z�u%ck+�5z����m%�t-{Q�"a�k�)��E�o6�m�&�N��~T�sc7�%8(*� ��9���%�{��	Q!~���]KM{��ی,
]��ךp(J�N>���.$7�7K�bj�-٩���v��fл�9h���W;Tc���|������n- �.���d�*�y��Ι ������5]��ZjQ]��P�LCǀв�����UjvF�x{�F(��M7�rfXC��ktݨs*�����C�Ѯ��ӄ':ͫ����b/���v>�q������Ǎ)j劽ɣ:�n47m�Ј�%�yh�AK�|n�ܭ���B�;����#(�(��/���5�y[P�HXtdee�����c�!��(D/�$��<��0�gm��ۓ+Chk<�TW�"�7���r��%��.��&���o,��U�WLD}Y�f����F��ZZ;����~�ӱ��Yx�ij׷�W�$��>�hU��z��\_�V�r5�:&�%|0�WrY%�؞k=��kE��Ae��)�4�(�k�h1P�bFu�l�B��l�μ썇i��S�k7�#��;u�������ʊ���[��� )\�}�X$�*�s�9,Õ���\��X�/%Ytk�|�7'9ꈳ׊66:k�꓎o:���[f^"���AFV0��Wg��oe5L;��)�1��|n ��y�9o4���Tяu�c�["�*����셜�R��8�Y(�G���AM����lo��5��m�M�_*{���}�GL#!V��+C9b���T�%Ǩ_MY3����U�UN�p�03h��.P%a�g���\���b�$�2��Om��7�uۢ�Y.v*��]XS�91����&�N�tL�A����UL��8��{��ó�����A���B�qmX��m��w2_[���ԬV����_L�^��PМ*=F��Xgj��cM^�a��pԚ1X#�.<����x�Q�k��u�e���t�����Ԃӷ�1I�W��2��-O 5�V���D]��(�8:ǵ%��Omp�(gB�N���g*��b�+no@����-��kD���7�ծlB��Y���Q�c���� L�Iv�n��3��Ǉu��m�N�#S�f���vWM��S��c�D�qv�l����O��<�3��R��sx[��cR����in	���j;4��0�Yr�uJĉ�8�]q`�g�)��%�o����8�t���>�V�񧈳[�{^��+�p�:��H9��n�S��u�{<6��x����/�e1�#p�P�d���r���꽝���eݻ�x g���5�(����D�w�^�Q��g.Špa\�����E%�[�����c;��;���8(2h��+l3���t�;\U�u�v����-G1����Nᄩ�L�;�4��K��W�q�:w�^O��'���ӽ��N-�2�Sz`{��˥n��������ym�#���;���8��Dʹ�cU+Z|:r�Y��[|8CXWYǱq#�b�y�`�ڟ��,��z-yI�yR��_x�ga��u�4����+c���M}/�[j*����*ؔPicFԣ"�iaiDcm���U�*����겨�,F*�h�eX��`UE�+lP�Eb�G2�E�iQADdZZ,-�DR��iQJ7-r�+Z�`�1"��*K�b���.6*�dm��R�E��EB��B�-XVJ�Ym%�)eҠ�,P��+�-�$U���DR(�-*J�YU+Y"VTV6!PTb+-�+Z��Q@TTDQe��l�����j�U�������kj
#%B�cmE���PQk*�+Tee��ѥ��Z��*��lm"�!Y% ��U��
�jV�´J�a*V	i+
���P*�--Utj1ٓJ���́�aC2R"�UnԚ��]��6�:I��by�vљw���(Y��>0j���R����5D��Y{�Q��:kǊ�1�tK�{�J��	�4(9DD�}ˌ�]�]�k4�e^W��r�.�#n�#���91��80m��vv����0)x�U{�m9��&��k�o!����\�)�{il�=]4�C�݃z�����q^|:h:ݸ��[˔.��2rewh���G:��F0ݤ��n����^�j>t3j�d#*e��;��[bnD���^-���a?f��� �=�N���G��l:ӄ��l�Q�j1Jjo��Ԣ'�r���ƻ��bԻk[�~vq�9�]���|�Г���\nc]��M�r�;��U��i�������jUE7�؊�	��]��$M=���|umbq�,bs�&mP�e	�w�����{)7=1M���ҬP<��gU6��a�&6h+�{�t�i�ы��BWwsGoR�]X��ɃoU��u�2�0{`�U��Bwۄ�QW���h-��6ͱ�r�jؚ�]X+:�n\�܌Mv�+FeKhZ�q�1&�˺�����a��j�fr�f�ntY�r���]�N��	%=��XX��W�.(=����]p�*�Gj(\q�s��fփw�-�;���}X�rƭ��+*E Ҋ�~t-{xc ��h]JΩS`~ao����=�n�"��S}a3���h^��ӝ7�ӲB���f�mSZ����\���gR#�{j�SEK�}�詀�-�D�S���9A�ØSY{��O�SG
##���3��8#�,��/qe�6�rimd��c�6L����۹7E�.�`M�����f͘[��N�q$��/��f�����M>Mz"wq�˳`���u0+j�]j�cy��A�[%X��|2��D<q��0��b-JL�T@�ܭq�;a(8[��LhXe,gU=�YU�\Pl^��7U�<^���sjޥҲ���7Lf7��"���ě��rv4�����kݻ�tm�-�Y ��F�S�]���:��J4�l�:����)��õ�v7��֋�F����:X�A3;bT+��6�Ǔmw����;�<L���#����n�ܵ���V�)�f�E�ٗƹ�0���
y��)g��J�|)곕.������I ���;�vc8S3Q�k�Υ�Z�P�o!��j�@��H=7Þ�d�17�]���].��:s�a�v��Q^񮝕9�lT2��:��@���6q�7*7�o�gV�?bQ�&��r�29����Wd"!�B�xu��m��%X�.mv�jM����^���k�+]�n��>��hhD�ۜBa�L���M�yϔ��+kŤl�W�݃�\��Z�# ���$nՕWՕ\�ɺ=ֹ�z���h�%��z�c{�J��V�:���J_Mw�kVo;��A����kۆA��$Cl�K��"l�#���*s�rQG-�5���e8(*ǂ�O��[V��8Fv���^�1kZ"���H"��<�	�ӊ�5�Yk^[s-L'����t�ެ�Ĭ�T���.1;�#�����mW``�I/���w�A����/.��V����q*_�t���ѝ�׫��hx�eY�3�%%	|ċ2�m\+8�}KJ�|�$�s/wsm�ttk(ᐍ���R�H�(��+�7�3s�m��pS��{�G1�y�KCD�NZ��X����m�ۋ�7�Է�M��"���ɍ���>U9Z-��܅�-c�G�r�
Z���%�olmp�al�,gU9"�ʦ�.
��',ۓ����v�V��Y�g'n��g�Ь��m����at�pU�d�ibU�9��� <ؠн/��=�g%h;@�(Z.4�*�uvc0�v��T����s ��������4�==��k��kt*��-��g�-~�U��Ac��uu��,�ޑ�����Di� �K��L����3[[���+���w&��>�V�Sa�ʶ��
=Yx���$�!�*Ý�E��|��O�F��5�^�+���n5�mo�f7�����طN���0�~��8P��q�Y֮�� -��;�JWמ;-Dev��wIh=R��pGA��XP3+�&�OC�r��x�ugW|4oV����R��:>t��K���o�	�ga���r5Z�HRs��%=��,�г����jJʹoR�����ӯw�{2�nE׼�sl�w�Vk)�� &��Z���$�F�e�[��ޮYr3��F8���X��ĝej�hICa�j"A��C�KcFY�1��v�����m�g��WRi͌�7��
�47о�����xYVow�̞X����͟v�s	C#���������ʫ�����rW���L
�)I�U�GD�s�0�'�+����&�9V�J��X1�	[o*��r�.�>ۤ7�5�+7����JSi-��o͊�����k�wqI��e�z2P�Yo�:��I��eAͦ=��y=x}��~�j�Ҧ{�� w�D��ޠ1"�}�i�R�*�l>Eg�����S���g��wT�T2���_,���$�ou��4�X�5;��T]6*�������`����au�E�H�9��j�b
&�z)g5w��t5��i%5Rx�'gnެ��T��aSH`U|q�e��ɫ��l��R�y���7/m���b� �E�/���=zެ�8rO�M��<����k��t�^���S�.i��gg�z	�Ϗ�C�~���l��o�Z�mk{�*s6o�/z�M<�-�=�r����d\�����5|�j�-c.�E;���-��EOmQc[�ar��%]��z���i\}��{���^3��l,]1ݪ��_�+W�;OE{��pZ��*��]-G�s!�jv7����gKm��+]�	�N�R��
���\0ʫw<������yڭ�4�����[��X��>9G��|ۊ��V��2ʓ�:������16�IX���`t��'X5c�RP/X;�Z:�J:Y淹v��t.N"Dcx2V�t�g:�n&�wu��YDn�������;�K�P����I�4@����՗�r-q��{���C�����f�ɔ5���X*�'iV{)��.62��X��}�մ����ԩ����̤��If�t7h��������wn�![�}���46,��c�S���=y�u��Q�f��5M��݈����V�]':��"`P�/z�_s��]�����q�4�uV�s�\4���<�١�^̏�Fċ�@��X�T���gܘ�9�^|"��D���W�.�뙁Aq�7g1ª��������x��'�j�1����c��;���1�O����[}��;r߮�ݔ7
���T��c��!����z�`�U�i�.ky$��75���0�lVj���vrj��.�U������%�c�]���^`���VR>���hq� �f�����$�	��{�*v�YiN]��T��Eyؽ<���\p\�+������t>R�_�Vō:��e�i�yزuu����
�b���D���P�Dm����6�j��1����h�Z�Oq��V���z	�t8"v	UQѢ+���g�����4��%iw�����M�w�=��+8qյ��d�f#�Z�ܖ�1�S�(�WOW���nr���㧻r�R�cyz���ͳr�ࡲekpc,M�Bɢ���y&����w�E��(�׀�*�&�}��u�o��Ɇ�<ꇯ�u�I���t+TQ�x�G*�s/rc6�#���s�~o��Ņ������e{�ն��Y�=5��C�e��Zr���9k���;f�Rc��M<G'6�$��Z�1k�ʮd�c���wJ��}�{{M�4�葼�hfL����^�h�4���Z��lD�z����c>ϢumUN/�"����u�^��?K�I���'�^h�<0�8�`1,F��[ҬQ�pW���Rٹ1�;���0M4�T����Z�f�(ݘ�xTu�֪�K����tq���Gs��� s&�8����Cݸ�y:���%�sꕼ���aˬ��n�<�s}�w�螡��YV^���6.g�[iW��p�N�{W�n�齽�(al�ϳ��mDX��Y�����;����bѲ�U�f�*�-�C1���A���z�C,v�1�r�W!5o��7 �}T^lPl^���]�n�������Z��`�����OLn�#ΐ���f�}\������Y�]J�d���H�`����ñ��W
8�S}6�����j��}uw�"\W*A�/K�p�6l������HV��3L�7�g��R��)��N��xX�2�**ޥ �MöGM��	[ZCN㲒�;�pw�l��H�3Vl�Sv��a��(�H,x�ݭka���؝�����	�\Y�]����6Ü�E��(>3�W��J���iZ���
��ɉ�V9���:�f�V��r8kU��b�_W�o��?v����!�Z뼞��Hח/$����ô~��Z�,��ᐈ�y��ej�N7awe8/w�s��H��'���a�6��n\c��kڈu���Dv���9�-o����#�ۋ�����N��@<<T�p>�@p�U����ף�c8+�����y�w
��%@cgvC�S����`N�����%C���H�
��v�w������QxoR~�=�8�p�*�f!���$<��}�3<h+ꗕ3�L#�7y&v�P�>��LVJ5��
���C�� ��� �UV�+������~���Y���J ���qb��DLVͩ�9UI���|j��̴�T�P��h��e���U
�
��p�M�>���ܟ��m�󒮀W�|�ߦޟ_>n�����g�����Hɔ�%9*�/�������#c�mPu�=�����{6��)J�ÀS�� ���b�W���m�����P@�V>6J��K��3s��V�(�؉kH	��|*`�m=�R�8*і]C­���!�$��ۄ��vI�f�yn�Yb`���p�\���E>�B��i�t�x�:ђ�[���z��AIƵ���ں>Dq	#����ȧ��H�����F�WW\�,e����r��:q�PWi4�Ü���2�A	k�����O`g���9
�9\�J�+/!]��	JXf��7�\W�[[��b��8���i7�0�w.��<++;,����#�:+��Z�Y2�rB �^z��HՎp���x�]B�?�W�	�p��9���B��r�U���#ckj�t�^
�)��	z�D��Au�*�Ks�lڑ�ˤ�A{$�l�<�N�Jfz��	ʂ然x��L�D�B�1 %#��
���R��]�ض���t��i-R��0��v �蠺��bֳ�l'@�;R\I�QB���Pp�i�1y�YD�oya��~���u����r��t��#vyK���fR�n�Ϣ+��N$͚k� �uQ7���`VK�M�h+�=�8��5�P����`��z
Tu,�デCGgM�Wi֕\1dN�M˽p	G�b�����ʝk�%�՟oQ0.�-TN�r���܊����,���<z�@fX�r���!�/���Ǌ�l��;�����ͣ������$�4�3{��|�������X��F�-6rX��k� LI�NQ(8�r�a�jVu�zzR��0����<E�γwk���-���ӽ�o�0h-���=�	�ӇGw��]�#��N�Y{ϧL?<xI�c�����#;G��b�J�m��}��6���̬�� ���3C7��7~;tq
@�J���0E����Emh���7S�*u7+3S	���B�)�J66[*�s��Nj�(n������s�^����t>J���#����F���.h�i�N�KЭ	�0�hJ�L�xh}�T붳Yf��v�uh�$a+]MВ�O��˙o�(\:��b�훣�K�Vn��;�X��E6�a�e6���&�Wה���ܸ�m73���X�i�cx|�ޗ[JM<C�:��3�x2�=��5�4�7s�r��P�ǵm��+��$�>yN+�_f��.�O;8\��ks����"�s��lR��WZ��C+n�t�6��Ӻ�!^�6�2;�S�(��!W�����s���5lZ��y�=�	�G%�0�v����)u��u/�����Xyx�*��ӄ�h���J��eXIC;�{��7@_kA�(9.(�.��ܫ��%����y>E�S��3)������7���P���e���W�i6�=��]���h|��`u�P��<Vl4yS6^e�(��9^��}��R�d�ݨ�g��):��D��N�8���*�\���5u�nKt�U���S�L���{��ؐ�9�e��	�`Bv�]p�V�8�h��;�tR9y�WEnH�S�����",(��*�Y�k�
�φur}i��8ءՈZY��dN%�9�m���f�K��c�uz�P9�"�)1&���ȷ��
-��.�s�c�眆s
u��7NSx&9F�5%v���!#5[ܐ:�=0	�u�0�#T��J��x4��M���m�6:�s,���U�ϐ�:��輶ou�=�Vnf��^8S=]A�DG�tU�Z�5����8�JM����{ب���i�X�
�[S�Ȗ̫x6d����k�[P\;�*R�7�4�Xiݍs�~�Y/�^B6nCH� �9��>ගw�)�*������e`����v�$�.Q.��´�n�k8�Mf����*�3��q�]s��'#-֐1��_\�X�)�٥�4��re��u�A]F;3�a�ݻ�wڕb�ۃ���}ݛb��_�v�v�l���l=�e>Ƀ�������{ج.�0�+��2���yx�̷�y�[�S��u7�D��8�
�
�ъ�*1J�H��lXE���Z�m�ej�m�Kl*�-#iYYZ��إjJ0�(��R��Ԉ¡F�KlXUQ���DYjڂ�
�"Z�*�����*�Z�Q`�+h6�EUF������E��,��V�ED��j T�H�-�*Kh�Dj�U�b$�PU�b�J��V�Kj�
�)%�*�`��jEZ�eAe��[aR�T-*�*1� �**�Kj(����"�m���Ŷ��TU���j0�PY@UmR�*� ���ԕ�TQ�ZЬ�
�iYR[U�Eek#ZUH��YYXQ���Q`TD�ҡX#jZ�UJ���cҔKiU���m���XV�*6���K�TFJ��-���a��ou׎�����5mJn=ĈU]=}�r�	t.^��F����|����Lдh�S
�sxw,u����C�O,����"��T�
�����T�]����Ys��g/ܝ�)��A��:*����{�J2�/�:��{mв�Pb2[��{"�TC�z:�	�n���1a���fkN]@ͣ�͖���s�M8*�W�<�CK���b=0�n娼�4�a)(�+�����;P�D���R�+��$]O��������f�b��C���z�ٕc�)��ƒ�����:{�0@��l�1"�{i^�0�aX���<��\FsN�6󧐹�a�g�@�Ed�,^�P}�N|S�$�V2K>���q[R6{i�xc)��;�˪��L��fI���L}a���`��^����P~�P��׈��	JE���é�>[���;G<O�+ų�xiݖ�#6@HM�v���]�7Z�lݽb�=���3��b)��}���jl�(¿d׫���2�C�7��
VIeU�v ����B/:#dfNF��3�>*$��r4�1s��\EП
�<�X�<~��;���Ɵ>�����F�L�P���YU}��@��\��ZgXYW�>a��㐮,W���Ţ΍S��rƶ2,f���E��u=���e^8�r`%]��ӻ8]J��ko���w��B��%��u,<�i7���~���2��T���U�T�*y��[���WE��*�EseD�x
���AZ�q�3�c\N�m�k6&����R`\?<WNxtەc�Ő1ڙa2-͉|v
�)>��f�t'�!;�I�]��uٚ��Aن*� ��`�9�뺵;a���}�x��n��<�V��fobOK�4�r��y�n�P�^o@�xJP�������`�3q�rذ�a�&xFV��M�5���UDQ����]������^' �T����CU�ؾ9N��~Xc<�� f��RB�� k25��|hX�Lx��(�Ct����+Nq@B�����{� R����d��ݦ߹�ͤ��|v�x��k�'.�X��mL#AǨJ�����{�V�~�8V��k)�������_���(8ȉ����>�,G�� �b�"�V�D����P˕5��P�(9vs-c�:}&�E�T�Ҝ��i���ժ����S�>��0�?Xo�&�����27����=��I]J�Y�}f*�>VO�~������i���H��JSy���
Y����qAܧ�Rc�->�9I%*�B�VMgs�/ݟNE�"�V ��1��������K�Q�7[�-U�-��,�5�e�rpH���g-�p����d��$�=��Պ�Z/KqԮ(�3΁�\�lGo�6��zu�)����7�<��\|-�U,B꡽jHf��.2*�uM���!6鹆� j���Ƹ�i���'�$����y&
us:B(k;CE/�,�Lh�x�u�cèuФ.����;2���Z+�"�.��F�`��V�����������:N�Q�Xn�k�U�V+ޫ���:eC�6B�r��%c������_�x�8���C������K����u��B�t0PDu�)g��Z�j<}j���W[w�0^|�n�'v.�d7�1.Ihħ���T��U(7>Q�(��Iĕ��Sw�.v�[C�[��eTR[��X3/��.	B�رJ� �g����~^��ꮎ���tE�\�����݇�UZ��+(ڥ2�jC����b�B�J�ٱR."��X쮽�7�Z�=�-�HO���ʩ�O{�h�K�:���7J�ˉ�mx*��a��y��3�9Ԕ9h�祗�"��cot=�9)=,\����"��>}U�t)pb�ب�2@�DUA���e�F���#�~2J�N�{�9�%����cW���0�:�n��=�ph�x�aT�nxL�`܀n�m�q'%�2t$��!8�f&�m�{m�y�ȁ=ҍ�Q�Q�ϖ��?�;��e`i�Ժ�6���8�T6�<ף.���v7�ƍ� ���u#jp-�Fy;<"��تg��R�|��ev��U��y+��g��B�(��7����x����g�l�`��Ո�͞�3!U��2;{1W���n�>�� �f�� ���yEI�fWuDSt�"q"�"\�-�gz'2;RKk*��S��PT���B�<n��J�惡��ӫ({�!C��
�������+��"�0�K��)��!�io��Kt�FYC­�[����ݸ���<�h\�q�����W*)�E�*+Z>��cK��m�� ���.x,�d�B���
�S��턠��}��8�����]�Έq}"��q'͘������9��2pI�[]6�5��ųl����Qu _{)''a7�/$��@�k��x}.�<�e��XW���>ӹ_w�NK�1��=���6وV6�U�X���i7�0������V��]�����m���L�!@�=�a�pe*ϡZӐ��X��hy��xa��^�9a����.�
?y��X��ʶ���o~"�+��j����x:����$x���s��'��d.�sc�pi�#�WW7��>��mA���0L����#ZWrg�wC�k��n��h�׶����8S���Gɝ�q�2l7�S��+eY[ʔI��� "�^����g�UB�����ɍ.s&�Y{���mԆQ���H��E���L��؛�rd� ���$Ԩ�t50�:��Y�I)8rCW�@��:�":(Օ;��N��v�����@�hi�G8�j�ivi��7���X�\:P����8.{�Ń#vyK��>��6���D-cl֫k�9G6��g���Dt���')Ǐ��>�8���qTca���'CQ7�\]vU���<�5;�ܹ"L�A }V�F�<$FM��x���Ϊ�gҫV�R�:�T��8��.�МU;�b�����|�$HS`3WӰ0T�MdQ�I�	pT�RoF���t����-K=i�T�+���G1@M4\\�["kM�@͓��7�\�()�=���X�+��%���j2���Lru;F
�Ll���̖�n)Ӛ�^�Ȯ-�$w#X]���}G(!��1
�������e���	x�%+ހ�%[l,��zR+Y����ޞ�kkJ���W�]z+��H7>�mnĸ����unWnnb[=�:����Ps��Y�=[�U`�+����ymF�1�_]\�=y�o}Q�e��/0j-m5A�q�Y]cyZ�fq���./�D)���b�i����t���nM�pu�v4��-���Q�VI��U��g�Qy�x|�ugN��J	���9���'1c&X�0����Y[xO�(�E�4�m��� ��M�4�������K��9w��g�6##fh%�/�Tٜ9FD� .���Qj��f�����J��>}��WY���h{;�(��}6.F�F.|�X���(���M!|s.�d��K�c\�6�Ϛʇ=zȷ`'a�����P讶�D�<B�#��F�z.s�j�kk��H�f��.����Xs�2(���:mJ����2;�"����+��Cu
\i�QY''��o�����5&V�]tӑ�J�ֈJG9�p{�*t�i�\�^��pc]NUec�ɨ�b߫սKhzszJ+��p������g���`��wa��V��3Mp8�g�=~l�b�C�H��9�~�1
���z7JyԔ5WmX���p4�U7a�"{kkN�A
�P�B�XG�!'GMz��y
T�A�*�ӊx�dн�!���t�))��1�i��)ݷ\7�v�Ƕr^��F��4D�2��SԎ%w{].�f�Y��ͫ.���%q���y���oVgHiz� ���)g`�S���m����	�(ACK���y@S��7\��}��7g���t�ӡ��  �����.�r�X}]!�q����=Sh8�J�8:�L�<��:<[\�Ы��N��L�L�Ǵl��Ɋ���5ň�
\X��b�"�j�H�R6@�"ϛllE'3��;�M��u�����us^�`��36�"&�(�#ÇVb���ݽ�	5��S��P�<��]I����1?yM6�@��ҠDDS�j���Z��VH�-�EԘb>[�#b��T$��Ľ��&:��%71�l�꾧�/�#��KY`fHȖ'�����NW���tv��\�a�'ԍ�ǼlDz�^���r�y�kw�pu%D*F�6荍���SE�ؒ�9u�b%N�Ӱ�F�v���X��Mw#��C"��\_L){!�#J�}+�k���_z�~�,�^��8���yK�=�N�����۪���s�(2:Ą�7��eZ�B�Z��
��D�8�[U=��޺Ԧխ����P���]Q-�d�ϡ���ONCZW�Һ׽0VG�9xFH3^���}Ỳ: {Nʊ���WO7�9W˪�8���a/G�Ϧ�o�)��Zh��N���;;z�#�`G�.��gu~)w)�^�ݖ끌�'fU�!�w1���T2��y���#�j�9^�����c��;�B0vK{�lHS+�V��BU]"�J� �=1#�������S�X6������!�Π�����U�u_GT�R:^��l=�ܗd�`e=~�g����J���4������a�:��=~T�A��ҬuN$��
�@�C'����m�MDd�P���6�ZU��`)9-�z�`d�4�\��V�qQA�TI�w����h6xߗ�6b��ɭK�z�2Xۥp�)�i�>�ݐ���$qn�1;<"���q1����Ϊ���'�0�ntT%��(��U��^آ�q|'��1��l
��+ )g*j{�;E>^B.ͳ~���:�����_QIٮ�����{��N���Z��}Q�XsQ�2n�}z��xc���Q8a�pɶ�#EKA�2�lz"rK�g P�F�Â����]13!��v�9[���[��LB`bw$&@�<���HWU� ��b���`�Q�Gs[8�d�9,�;��[,x!�+�k5A�.j��"��h�
���5��S�3�\R�]�A>L��8I�$�S�;�NS� =���!��8�X45��gvl������"�MGi/o�h�;3��*�D�f�}�X2����ڹ�[���|nԩ�Guu�X�%���˔�o
��[��Hj�.�
��[��y1ҥ���-�� �P}*��a����8�}C %~pF��vv_H��!�>a̦��$\�Z7�y<��Xㇲol����Ô��을�;��k�����O\+Z;EӎwEۮ��Xܧ^�Q�W��Ĭ�)�W5L[�7���e`Oy��Oj�~Z�L5BA/z�9%B��y��e*̹Ε��&k�Hr>Dɿ=pe*`���x��P�2�`�Z�6�>�Z�ߋi[�.��^�[W�T�O��!W�@E�~��� [>�8�ld1R����CZ�n�I�aM�tcl-.�'*�n��bf:&���n��s�ڔ�6s)�<����<S�R0���%μDtR�ʝ�Y�6�b��%ėB(ᑉ��H�so��Q;���ДF�q a��T!V~��=g���o����|���(ʔ�%�z��N|��V�:��斈')Ǐ��8'����Tc��9~����=���*�Z�Q�b���DSU1���*6q�"2nT\�76#�:�����Ε�hv�cMI���W�e����*ۗ-/?&��g��w�bzV
��W��"�%Nz��Sla:V���c�K*���W}��g��x
����]I��_��+G.�B���։�s���(�SԞ�D9�M3z�X4��	�Mr��v��h���wQ[��UZ�J'r5�v�w�F #�;L�>�u=�<�ӂ��E�O<�8��U�a�Gں��L�e�w�^�U]���0� t z�Ԫ����$]O�+\��c�6Iy�ή�r>�d(}��64MC@s���LL����y�A����ו��	ܧ�0�}ܺ���`�F�"24c��9Aȧ,`�1
٧>>O�l�a�-e�C5���4�;�{���|�`���c�~%�zV�=��)NC�,铹�R����6���x����0�s'P�6�x��8v2��-���B4�71.�j�ړAۨ�c��9<؎0��ױ���f�dl�Q>����8f��0�&�E��*�5ПU���X����)���P{;EXf����F.|C�4��U�Y�[�zU�"H�������&�-����P�޲-�vxz1N�U���Q'�P��P젴��<���m�tz���dz PBT� �Ei���}����u8�8�-���?W�$ I?���$��H@��	!I`IO�H@�BB��`IO�H@��	!I��$�	'���$�Є��$�	!I`IO$	!I��IO�BH@�2B���$�Ԅ��$��B��B���PVI��{��� �	�` ����������z�!UD��"YQ����4$P$�TT����TT���Q�����R:�UT$@BAQ�U]�Z�JaF�fm�o��Vkj`f�kUY���M�U'��5�V��Ǽne�c%�6K4e�2�V�]:�K��6�U��l�Ŷ���a�j�&Tڙ6��_g;T�c6ڂ�m��,�,��"�X��c*ֈճm�f�me���+-��̦�km�Ƙ�5�,��k5��YF�LlV�kV�ͳ**��٧M2��0�� �/�V���[C��ݯU^��wn�=w�/S5Ҷ��Ӏ�٭�K{�w*�]�WY��Nr�o{^�Kq�����ԍ;�VN�5�ws�Mn��+r;�ݷ:���r�l�٭4�Ͷ�j�ѩ���  ^�.����S^{�쮕�Υ�^�u�Mmgw{]� &�v�{�;��.��v�{n��M���kwvu��ښ��n�v밓sڧw��wv�l�-�yNθ���Xd�:-�BMkY�Ī�  �׹k�ۤ�j�R�����ݵ�N\IٞW���.���y���[m֫Z��;����'�}��EP�(��8�@P(�F�(��(�(�E��S��(��}��jV��¦���͌Y�j��  0�QEQE{{�w�(��(����1�EHw�sO�΅Wkݗ���Mov�� z8�i=�{���g���@�������'k-m6В�Hdm�t��  �}��Po�� Q��p�F������o{�x�M&�y�@ m�{լ�m�1醀����k��P�X���׽�֬m��b͙X�k&�,��|   /h@���(P;�����*z�Mu�Y��w^��sl���ל��{�����7��n��x�z���Z�v{���H^�^�&�mUZem����0�+i��  ν��l.�\������Q��y�Z��znޓ�7W����q�Q�Ͷ��.�{���wR�sǻ����om�ޣ�^k�mwuF;ѝ驶��m���j�S��zv��{<�et��ٳ-��r��  ��ݽm\��=���kZf�{s��^��[��X�v붵wsJ���*��+v���oz6��ۻ��EoV[b����G=��nݚ�����v�ű�v�v�{Y��+wuܩ�R��4֭�aM1mZ��K/� �{��k��]�kӃ��![���^GnS����S�G��N֭�/^��
IX�]����Ԏ����w,�u�J�wv��m���D]�ڻox�Q�fhۯ,Ŵ5f&R��Y�l�_  �>�G�Jj����uB�d�=�s�v�u]��޽ݺ�[��9�n�����Ͷ˞�ޏR�iWu�n�{Z��4��]ގ�e��[����;6�mN�˓�Uo�"m4R�����$�*   "m2i�U=*=54@E?�F�0 �a�~$�UQ@  �a�Q `O�?����D⿌�7�����6�i�̆�ES/:��:�ח�~��* ���7�삢
�QS�TA_�AQ�
�+�
)�s�k]��=����vw���¥k�S��3ncLn�*�2�|��l��F[��Nn�����-�2�p`��+cn���km=c\�a�SX���*r��0���]d�`�rܡ#n��K����`*E��/rz(,�c���fn���H�����cl;�Lulc�@�ƶ�d�B]�Sa�u�ŧhL[�[�,Ǎ\��5!Ÿ�.۬E�6��JL�7BR���NU��Q�f������Í1�,*{��M)��)�b4.�SE��ɀ��j�����r�S^i/��%:�z���Jݩp�wz�G`�ךn�������nѢ-�?Ab��L�5���i+Vw�\)ZƮ�R�I�l�׫$�;fŨ97b��V���Yj�G2i�r�f��j�-�m#YIGR�@Q�E"F�,����YwoM�-�Գ��Z�*b�+ͺt�[��go4d-K����C2���ee<:챪��lIS)K4�HE�5l"ѼB �\��3-Ǒ8.�nQ�����䬆�-d7
�rD�pC
�J��P|��E\t��!ŵ��>�:���tnpj�7
�[��DQn���
��&�Rua��X�:SdN��u���-n.�3��3F�jf�ko��e!�XٴՒ3^A7op�.��
*�6u5�VhU{�Њj�mӼ[�.T�@.�o�Fg��;Vf�J��sl��[ԍ�!�k&ѫ_[�UE���$��"[W3L�M�����"��c���� @�^�wJ���p���-t���2�'6�Y���BRp�6E�ՙ�B���ckJ�3p�1jĕ�&��"B��@���AGT׃t<�DmJ@Qgf�l��}s�CZ�y��n�al���R�B;�U��N���V/5, ����Z��� �4����uc,��&�ަ����tr���v���;j�b[)�L0�Z��k�p/4j5�c���+�-�KcC���^p��c07�q�YTPdĭnhӐ�2�[�e#���2-O��b��M	�T�ۤ�nV�_+�,�$��ܑ�2��lO(�ɘ�*��6�hs *
�6�;�dR6���M�������ʶe��O%@X��KF�f��L&���Bӻ�� �������f�]E�wV���"�j�Zy��l�,���E����G�4��!z#:�^�Eۜ9n�5(��uҤ�Hd�j+&,����H���u��۴�9���W�Bn8�U�oTX��m:B[.�%�Y/j�,N��-]���J�n�(��4c�I�����=���!jf�*��e�j;KY	�
��F��:�l�vXKJS[e�wK�dib�n�ec��Y-2Z�QɨU��(^�y*ڳx�<�n��bT�X���Gxb�[ͦ�nі���:f��,l��rږ��l�j#@˴�Z̢^��E�-Z�ޔe;��a9Q�-�w'ʖk��^�n��q�qhM�K���0:�O�
ω�-y�wiQ�ii��Ǖ�cݩXu4n�ula:��H<����Wlh��%R��L�菒�-�!57x�݁��"f��7u�	Z��H-ؖ��v����A2ݻ*Vw2�XB�	��mJ{�!V�-����.�re!��Bo/E�̀
��V7�ib�T:F���C[t/���/���RQ��@tjV�jTh���%�%�O I���8QYSsM�i�ܵ[��I؅���ײ݊
�X�쭹@-OI �1,[t1�LS��z�7�PqX�9f`f��8�Ū�5��4���+�]�b�RԏRݫ� o��f�X ��W�m�Yb�
mbs��e���Yn���%��\5���P�ͳd�Q!�W#k��TU-���� %�q(&]CX76�F����vf9u���์�͉-�[�.k; �ؕ��44lm{L�x����+����$�-�ST��z5��9H�o@3#�1|ñ���ǧ08D����Bjoٲ8.Q[u�́V���Z�37l��n�ubN!.�U-i݊�(bK�X����T��ᘙ�Ҙ���L��4�cx�f(�HJ&[�{(�����Vaʻl�U��X��%\cP��NlV!��b�ݧ�i���+n��Cz�ʚ�5��U����F�kF�]=˫f��iTp=��Z�U�MM��!�ǀԽ::��Ӈ�1O�i-�V��)���,K����4i h�A���*+Ka�5r�D\�j��e�Z���7Q:Y&�j�l�m�*�U�z���a-�n��`ӭ.�i��V�A:ՈX�e�5���YcNA]ٹA����!���4�,0`�J�E[Y���qT�Y����2�˦�@�P{��J-iR�dXk`��ܦul{ �*��ȶ�7a�d�[FV�ooB�o�N�Ш�ۂL�@��9�vmmXj�Qu4U�74r��I��U����
n���f�b-�e8DyDe*�xr�a�b��1�,5�iz�`���nD��ͷ[u��҆詪^�t�=.[!��eĮU�ś�=�7#=6�j[�8�Ckv�zu1n&�+k&f�8Ty��$+Nl��a1��������f'wM���qX�NM��J�����+n�N�T��R�P�3wh�sr�;�)mA�K;���#H��9�|��n��c-eKs>{��$k��a��
��Z�V]���8���6�t�?�{k1�Y�Q�MK�u�-b���T�d�P���$Q��8q��Җ����M�����4��Y����O�UyX�g�V����-��a�͙N��a���C3/�t	0��r�VJ�HH��˳�Ĝ� ,��)Bf<4[@�q%�dV��R���'�G	����m]:��T��
L^�Q�� ��V���ɼb�n�������]Z��FӗWW�5����5�|m�I�n��}q��r�Y!��P��nJ]W��fX؝`�r�-��j1�A�zKԙY�ܺW�,�)"���;7N��` �݊���IZ�ݪ��)����=�t�h�u �P�U�֑)�Q`�ɟ<����-V RJo�&㨵^�Ѷ&AV.},�0C-�)�F`6r��2�7�o�L�#��@nJonT��ɲ�涪U�ܬTu�*��L5t�`�N��@sD).)s`�u�U�)>H��ֽ1��Y��t.�XB��F�n`���aU����H(h��$
*Fβ�;����Ȟ&�eL+(�u�kI��R �y���a���)*�����*���H-�Z70Zf���[�%�k3���A@p)�����MD5���I�vZܔ�7F(odg+N�1�d۫Ӵ��sUC���	���mQ��b�*^�Ք�!3Y
=��Dĵ���+��n�wY��k)[�s&�e|��kp�,�bOsL���p�W1����LPTE�h�TD���j���U�	j�7X�i����@�6`m,��Kr�b9�����w(e4[;35`�@���ci��ؚ�A$�
:��"άsdǲ�2m[u+Դ�.#�I��!ѢV��^�Sy����:.:9I��x��[d/��P�! \)�����n2��s$�i����Gsu2�6tr���N��Uِ��C�EQ�FQ��-�F�D+�:wL\ܕ�-��1!"�Ʋ�q��*@+�i1V=�Nj�5��m#G-��%�Z�ܕ�<�Ha�L�m��0C%L�fҽ�n�!�wX[5�t��6n���l����'s�4j�� �����*L���2�[�b�P" [�e����4��3YÊ��aN�� *�AYu,$f���!�Q٘AYx�K�F�W�ܗ�zi^��JWR�k7	Re�Z^#or� �O5�4":*��j���ph��i��
�,E�
x�躷�����&)	�bF��"J&���Ysq�yd^�ö�j�`���IRv]m��BYq:5y.M�'�U��sk\��!��^�a��r�6��x-�%:H��h�Y���Em��jdŔ�խEZʎ��-&�P{J�%�@�֬g1Q�	Ït(2��Q�H�St�Q�q����B!ʍ�mԲ��U�bː6Sj�X����v,:`k���V=�m��[���\�3@B����jj����#��k٨*���+��ř�O��6���j���n��7P�n��Su�7����T�ڥ��u``��VV,�����466�Ѭ���(��V>��N��+A��_��Bp[	��
��ve<Օ��;�6f�i	 ���ۍH��#W�N���S��5�A�-�6R�/��Y�nF̕xL�w&�%�ɥ�A�wp6��XV��b��;�S��5�E�9hљc�ذ���w�h���T��[�L�jLbP8VV1`��B��kU�5U�u�t��J���{�!W��y�Ge��ҩ�˦�l,;��S2�oV��D{,��1Uؘ\%���w5
)չ�$�%����m��4Sʖ�b��bPU�I��V4�T�v3���YgK�V��I��H��AJ1DM�ͥc���Z ���U�ks/n�4���+tnN�5o 6L���M�KSR��H(֐n��R�-�J�f����Y�4wN��m�Ш�x�^���I�AL��7�q�e�6I��-����͗��U�P2���c ��
r�Tb�h�f���(V�WoX���Ua5�l��lJ�T�Rm�G4V��A�vD��7��F�.V�sv������ܭ�dǒ�5�-�M����Q���@-U$1޸�1 U���̆�vKN��X��R\�d�Z�Yܫ����	���8��Y��=��P���Q�KyW��I�hM���a飰m����/��8���Tj+Mf.�yK*��hr�đ쉨V�l[�1Е��: 4�J��m����v7�M�pTCa�6U��֞�k�v�-�-�[�m-eM��d�PT�,T��t�n�]�K���T,n0Ykc�&���15kR�nl�F�;�*Μx��EH��g���t�¥����K���W��+T^1�CհG32�Qe�:�&nA�i'R��,��M�QU���m �,��f�4Ļ?/�T��n��"�*��$IB�)6��(�T=Ax[���6�Tf�m�pѺT�5�5��T�l��)57PkI��Z���(��&�&�!��Y�I��Y�\�(�Ʊ�EF/Nm�`��5� ՅKCI���B�$3�(�JT���\A{6"��̂�}Y�{:x��>-�mS �����)^V$�)��ӧ��4���g�/��Qz`2"*˫T/X0�^HݳY6�kE���j$�ۓ	a
��j�%+DĽ�]\B�³#/k �:ݭnଵ 7[��xt$�J���k�Q�:{�i�w���0���uF�SJ6ޥ	H���Fc�� �˫
�J-�F��*QnF��ҍ!�\�7DcaN�rf��\)õ��,X�w0fӽ-��A5�m�a�;E�̭v+u���y���dH^P���AG0k2nZ�M�%��0�v���6M's&,iSk"�ۏn�6�2�Nm�i^�7p��������b�髻j2�� �d��%�v���Y��+$Oؚy�d�U�#����G�r���/lJƒ���ee�X�+���V��
�.��$d
9�����l��ʘ�Ճ-�* ];��f9jjCK]j���f_m�a��Rr�D���i �ӷB���l����}�!�v�9�G֓i���Z��i*Ǩ�ۗ�겥�ZRF���:�����,ضf��4L׏���Ҁ�mѺc6�b@ԇ[Fk4Yv~JL�h����(ˤ��8�t�Dç��kK�Xs3[�V����n�{>hc�0b�&\����Cj}�o^�bJ�G��-n[�X��É�m�dH�I�wXi�V�+l]n8�T{���T��9f+���U��,cb��ْf+)��)�aeYt>ɵz(��e	��KP��5��vpc�m�fՅ�mı��j�EW[�-�ɉA2�f��i��J��{�Yۉ�m������B�����Rv�3L�t�,�z�0ҭԥ��Ս9	�շzi7ףt��_b�%��TۉD@w[�R�Чt�s �"ɵ�����9z�ې�}s�˻=�Q��n�X���R���פ,7&��^K��$�o�o�B�e�Z�D"��/��x���앛tO���`��+U+!�@��n�4ۻ�d�w��[C5�I��]n�":%�"b(֪��DT8��Y�Z��L	)�ot]�p���4ip���,;zZ�e�� 
`^�����Ba*�G��ə���N�u��gn��2�[2I�&�ׅ�e<b� ���1fS��wya$���m�t�Y��O"T�e�q�A�@^#�v�'2�pЬ`?=H����mjjV��Ax�eɗIbDQRHl�;0\s^Sr�e�jf�6LB��m�2�p�Ѻ*9�L�.ؚi��ʽ�u��ۭ��&d�J���,l ��9�L
CE��q�&k ݔ��7` �Fm�D�K!kK�q8����qu��f��B���Me�s�1���Q,܎�n�(��u�cT"S-;f�D
r��A�t���i��XEK�)ٶ7.o�^l�ї��u&I��BH�0!�Xu&�bյCtЫ�ˤ6���D�.C������+Q���i{��Y�L��7s�ؔ�e[і�a5 b׷�(�c!f�3�Yx*���!9��+
�O]�tM.�Bw0ҫ	��٘�p�H[�z���b�b����wcx�rRVL�
;Z�.ۺ�nܫP��?�M�N9Њ40�*)Wk�r��D��ꏷ�ܮ7s6>�1f7����p�Nk������Y��^�&�n`�VS������Cd��u��g���.�1Q�%@8w�-��s���1c����1�z�{;�ʮ�T_t(�����_��Sn�w��e4ݾ�nL���ٛ�����ۙ�r�F�����j�E�^�[5Lu�u�l�)�p�e�Lv\.��삺� M��p;9��k�����t�;���˥{��J�e5����M�M�x�8���8vQ�W7S{���oz��L�=5�oĨ�rCw�3\vX�Ɩ'j�Զl�[�F�٧�l2�5��m$Bw��.ٷ��$���X �{,�mtm���6a��{g[��W�<��!�<�M3��8�Q�ty��_0��ݕ0�Ĩ���]�N6��DM��U�u��VE��G@0�8��ZDV$b6�&D"������U%%Ӭ �<]^]�:�7�cut2�v�N����bHL9P���_�{yG�xJ�]-������y͢^X��]vO�v���-���(.����XΑ3qN�U���}
7Y�rd�9Bt��3�ˌU����	�CMiO(��{��V�C��j�3n�2��� HJo,X8��iu�@�g'�r$�c�ۂ�5RM�Ā�v�w�&��V�ob=����!{(�oK�{��Y�q����!�#3gR�Q�\��Xq-6��ݳz�m����F�Krr�u�F��H�٩:s�j�sqD���x�[����}X#�NQ�Ȼ�T#�h-�Xeb��+D�w�j�gr�J�qhU}f��wm�}�Q/(��`ރ�w�>�wtCk7��L�F�6:�����m�wlo`������V[�[�	NUf���r�o`�`=%t�vI��`�\Te�ʼ9-���K;4B�z��h������k�jDbA��][�k����ӣ�:<�5�C�Z�z��ҙ��T"$�^n\�X:���IZl.��JN�F����Ք�7: ��ڼ��D������x�y&m�:�p��+��A�;��g��{4�FΤ�W�f�]lʇ�.�����qCF�/���V҇������M4{���L�\!?e��-C$ǆ��/�P�X\R�t�ܵ�0����4E>|s��$�m\�E�Ҹ7���V����r-">X�dU���p���R
Vꢸ�2�P��u�f��ˇ��+`cbO��|^���W��+��[v�!���i�����t�1e�bw`fl+l	�yt�e^���윫�O����7�9
��fl�^�t*m��Eb`wx{u���>ҝ��rp[y��� Ⱦ�PD�}[%�H�N��[e��8P��t�HL(1{eVM�-p�܋vo*�'B�o5	�k	&��o�)m��e=���EŜ�d��es6U\��j�`t���W�TSgx��^Z��'(�o�&�q�wv���-H�q1󥚕����@OpY+k�0����u���Y7�&�"���֗(q*�����Ne�.ok=Γ�*�a�ΗrF�����(YPn�M��%�Gh��V�nZ~=ghI�,z�s�I�K��,jS�ղ�B�M��y �-	�_hՁԨ�P���>JǑᄄ�P����l��ۚ��9��Ֆn^n�'���Y,S��'C�xx͡3Ou��K��k�1�vt�ŏ��m���|4Y��#��-�qf�Ӊ���u7Fĺ��=Z?wm\��k���0�=ױ�BUf;���M���{r=��d���{��q�Y�=dH��6]�qW��^6���#��,��k��vm+ᛐB�\��/jp���M�� }�X���(�>�.:9(R=��	�w�]LڛSu]�h������.-���Q{��
1]ssV
��JѠԱ\��}6�J�mpٚ��[q!���kkp6��:��.�Z2gCh�:M�]�yCz���)ƥ!��Č�e]�1L����ܳ�.vN<�2h��Ī��;��/�I�x[�\��.������F��Qr�[�K�+"�*r"gnKډL:$��jڸȽ)¢�CQU�o ]Sq�9�Lն���k9C����Zn��z�C�%������ͫ��<����0M��Mn[�+���bȓ:������y��w%#��a�n�ܭR��.�P���جܝ���U�����ku��Ƴk*J�]��[ǜu�R��/el5�e`��>v��Q�� ����a�KU�:��|�Ul^��u�q$pF��0��hMMK=�mӢ\�48��������1���p�b�wb��$�����uX�
h�!Ƃ;%����ޞ�
V���rXܐ\����.��RL\�e�������*P��6á>�w���嗚�WAM�"�(8F���pee6M1��-�+�s�h��F1\nQ��b譧-�.�g�Qޤe��lvɋj�Y�)����;y��j�R���)Vt.�]��k(fFJ��%j����j�e�W��K�Y��c�9i{�Jز`#2�Z�:�獖a����Y�&\	˵��3T�U����͵���<����e��T+o�/3��[0v��wa�Z�U�эt"j &9�+�V��T�:.�uf��k�!i��³)Jǉ��v��E-NX����֖�Z�h70)ku\���:4�BH�"��ɫ`1�/xR��*�\;Z�4j��\�(7NØ�=�S����йN�\�K����樯]㬕�R|ix���S	�;�X�2VT�y&a��۔uf�qjP������n+�`	��(OTn<�t1�S/����v��vd�6@�vn�B���^R�+�4��.�T.�£#�Z�DR�Me�;�
��oM9v�s�t�b�%���n�C�փ2ԍV�\�[|��wB��bo���B�S�ۂ��E��<�.��jdg�ʈ=���B�sWq�W��X�@�Id�mm�j��S@��t�Ɩ(�;���ھ���'lv	�c���Qy����Q��,�@s��W�P���ܢ�+�Y%�L�ѓ}+�Y�Z���K+B7,X��wu�fz�m��u�{3*�@���V���b[Qֻx ��G(ۨM�G��[�5�5f��W���>CO5���&����T�;���:��B�rJ��]X������j����vD-�wq ��D�++K'T�;)��;R��/�(s��=���v6]������L�����'U�)_Q��D+����ː�� V9Xlf�4sYC���A̶sEM�h��9�@�(g��E�#���F�(úS�2/�j�`($��F,�(��f30��G6�)�j�	�Ef�7i�s&3f�Owo���+q۴��'w�$����Q��5\�pV��6��m�Ǧ�h4�Ufm��rE��>����Pp
ɣ%)l�v�e��,WN�����R��_A\��{`5�� ��י��7jMb��r�w϶M��<7���kӲN���yXň������Xʂ�3�3�|&R���N;�d�wEP4_K��ɓ	�x�j����>̀�0c|��+�T;b�)⬠I���"����9J����̕�a�ӟ[I�q��Aqq�3u}]���ɑ���w5��K�&[ ۢ��.J6� �w%p�f_���Ƶ�8)]�=�F;�%1�w2t9`i3p�+r�"���#x�� ���N���D�P�x�&$I�t�<�:�ە2`�v��r��H2��]��LɈ�)R��3z��Tξ���aM�4����PBjf)w#�����<^ߧg.�y��q��I��[�|g-7M��:�9��UG�.��mp���X�e�uԣ�l�9"0eV㾺�Aы��������R�u��$��O(�A�5��i(��;���/�w.쫚�3�b���F{ut�YS�ڝ|��mM}-�[���ad�.�e�;���qN�bnr��Ǽb�fN���������2�Rj�^+�Rj���h�� �)��5JIefAN��lr�wZT�U.���)���h7����1l9ݮR�ddՋ\J.U�<m�����h�������)FD .�+c�ed�v�o�z/�W<��I�Toꌺ�)* p&gt����ݥүX�L3��"�]d��E���lJ�SyP����[��yK�4���'����vYN��qdMc���%eŸ����	o1��~��']d�w�� 9��_	�Q����%D���l��SV���_haɣ�$�U��?����M| �r�J�z+kC��e���
̓
iTp^6�6��]�I��u�+zl��Ƒ�L{�S5+���#��t���h(��.����B��J�U�Yol��b
����S'aBgD#�Hޱ�nԧ�I�����2��϶�v8U����y7�p�+�����F]L�U#�
gW�!�Etu;�����m��w.�6�ǵע�J�w�eްN�*Qΐ��8,�퓄�qJ�g��4;ݴ�L��3uͿk���g$�):�+3�h�ϡ뮐�B�/������&���oeH-(V��+^PB�uu�ށ�޽z���{����/oC1�w5S�����e5!����ȟ[�Y�.��p�m�ʰ��kZ���\㛡�MՊ�I�i����Ӿ���Z�b6�ł�9Gj���]��Hګ�9b�� �;���,d"�-� ��s̝�˂�����b�cbbQ��b�,�5]�"7Ԫ��cQ�}&�Hx�qB�v�ʺ\��p0�[�r�1l�N�5b.�8a�l=��@<c:��3��U�	��U�4����ԛv�]%�:�06���S�3*��q�ӐV����۔G-7��Pa�=$��je��5�@̙�T�Yۜ^���>F�HF�F�mh�rkKv��"����e����(��u��%��y�)�1!ݢ�=�"��ug4�V@�,�g�"@[�Wˁ	Q�g"o� \.»BaY��w��4�����Yzm�Q��T=�s�!X�;dUSu9zI̲��;jV� f_	 �]��֎�7��daPI;n�}y� LɃ_1���ݸ�dDV~X�w^�P��(&�se�;�`m �$/w���T�ٽ���ۓ1v�d8�88�2��ΈA^�k���4gT��_�Wv�]G��%�em�-gf��S3w��ǰ�ujU��A����sz\�#�9�iI��Ahw�+�7���;��Д+k��l���N��Ey����fJ�W&1c�]�xn(��U��^����-�WGFZ
� y_0�ϷEeg׋����w"N�����u�h*�e/p��6�^=��ۮc�b�d�G���&[�3���Y��!�e�2���شV�K��m�1F�u���/�W�u��<�6���ݜ�b5��3���c6��(���95v�FhRY�p��v�Ew����c�]W0h�o��g��w�ߖgm%H��D]��;©(�2�������!��dpfј��p�)s��/]����Њ[�0Sr����l	�%Nוc�_D�΃�n�Ar�M̳z��T/�u��3�7I�tivp�BV6�r5xeN�ʆ�mfZ[���`C]��՗5��9pc�&��Y�Vom,C$�Ρ��T�g��*]�v�v�J���x
�4��(�.]�2�"X]+ޥr�RdYdr։,{gQ���]�*c���\��R�V�T��1���7[7���ǈ
��r7z��hḵuk:�m�ٗ;{��a�/1▤g�e�U�Q;�L�8��Q����wv]�+�T�|�@S�/W+��.��Ǥ�,�P�uF�ԑ�mә�g \؞^'�w`�G;{T�>"��cW0�4��
f\�}W�3Z�&�Q�j�u���1���V�I�9
#r�X��� L���[�,!�b۹�޳��"��eiW�9��������o.�Z��(�Wʶ[��҆�xI3Q\/9���%�-1%������f�Ό�9��t&��k�
��� �G�u`���=*c:Xݭ��u���:o�d.c]�6�%��6K�1?��n����[�an��=�[t��W@�%�Y�̣�1\����&��9�}��eo*�i���'�:�\j8��,9�uhr�=��*�_d�mD_1�d����Dm�VE��n���7�6j×%�1f^(�[80��)��
͘�pB�X�W AfR6m]X�fZu0c5�ڝJ��P��ǜ%�fZ�4�Q��p����45���ԾC
I>G�K�d���&��z��y&)7����؝��dI&.oa��wR�o�o��;D�J;A�źK-p|��ɨˬjW=@���Y��v�yh�y����k3����t��N
��d�tЋ�֭�뛅��`��t���(�{���q��W
�.�>����Z8y7������]� �컮��PVz�����1���g!�H�n[�0uys��S��mU�MI)�u����vq-�za)Mko�5�5`�����n|.IQ:dotQ; �i+;���"_��|h6nn�2U������N�!�a�|����s��t�m���+��Ñ�$P�D����LGE�}ʏP�r!�6��:X�C�kn�S�e#v}u��棦z��ǖ�	;,,��E���1��é�c���'S��Yu�zn`=�yo(j"���]vucډ;'�]J�[s�V���U6�m����a����A�^� f��]� ��V��{2c�㘥�2K�R�}ܰ��P�P"g&zZ"��m������gwܻ�@��W{DfE�wķq�s��J�����6m�x�}:�n��D�	���QO�n�Q��e��4�.��i���~��(����ED��ǟ�����NSI+�à�R��%]Ҵ��k��Ĳ�ˠ�"iòG�m�Ĩ�/e���֮J�5Wz�����T��y���e�g_�4r�n�E��n���"�hhuC�
賕�
ּ�Y��Cz&�KJ��ب������OTC,�ن7ȵ�kT��}J���E�{&���;��2��/"��8%q��㹘�������u�t6�#��]k'PB���7#5��`hw �:ܠ)�e�]Dq�m9p�ж�w1�{@�U�kN�.��'5P�U�d�ٲgn�4hfg�:��ՖE�dn�n#��cmu����.�q8M�>%dO.�[N�	oݰYz0�Ki��[�\l ��%k����N�IR��e]�	�8�$cmJY)�����](�sF�Z{7����V���q4z�Ő���uM.X&)�U�[�[z&�{��iaA��@wZ����Q̭b.˥՗C&�e�pL��.��K��O�l�� �`r�A�A֕�M�^�wm��6�*���W��0�Y�Yz5,5A�V5|�%�N�%�]Ypĺ`%彁�-h�Y;��c��׈sh��et���Z�
���vg��l�r=wJ�<�v��z��b��'�V�ϒ�BV	ca�Z:"�ԗS��������P��O-5�Uj�!�:�8E��vT���h��xwVƋQ�Ҏ�� �J�����2�<nj�+��B
�g:=��H�
4�[4��Gn����H�K�c!���%�Y��7vX2f�z�<6l�]Gc`u��2U��{�kj�P�K$�V@��y%^u7Tܿw����r�S�cwY"b+�ٷ���%c���r��^�K
�ݖ�(��̏6�s�ņriV-4��ʼvU�P�#;��%U�;�i�@��μ45x �rn,��[dv��ə�k'�27�����!ݢQ�Y�]�h�YGN^�O5s��6�D�}:L��s�Ӡh�fKi[{�*��6��6���%+A�v>��"�u��7z�ι���r|tJb����V�K�k$4-���FIW�8Q[ם(�=��)�+7T[28�/:\|B�|������}vۺ7�P9���9�#�Y���qtN>+ ���vԣ6u��f9�u�r�Sd�2[�Ǵ8�W�s��w�r�PܣX��pA�i]�}H ���fT�yI��3M��hE�_Y|10�u�S�G\ҭ��5�|nFLZS��8��]7�Ξ��6�MO�[BJ�����9ID�F�+sV:Vֲ��Im7j��0�!���v�I{*1=1��g`�I<���H5|�5�=� % [��T�yе�!C��ZyJY��,í�1�P��b��7f���������. ��c��)l�+]�'0�BLe�js�`S{0H��.J ;��du㗈��'�4 �n�ZJ����QÆ�+���Wme�'�ue��d��bY���ÀPi�͡@-�ל�\��mb�#?n�e�yr���6q"�I���1���#�V�bθt٥0k7mE,WiN'27:�(���Q,��\O�·�P���ms��$kG�N�G���"��&FQ�;e�Lv�kU��	�;P��Ai�� �k*�!u3/&�8�5:�N8��)���m����Ů<�Vl�ķ���Y��l��-�[5*[;[���P*��m�N���0�U�E(�X㮐���C�Q�[&,�R�Z�7%$�w���u�{�{�
o��޽��.5b%ּ��7]kO��'d�P�}�+����/�z^�-�NK��=�-����^�a��8�xֻ���H�|F����f�e���ZV���5�/���0��Ծ2J��{W	&����da����`Hb�[Ǘ
]f9a�-E|����_.6GK��}��-�wS��F��؄�A*�n�t��B+��H��Nϻ����}|5��&Yhc*��q4�p��`��q�za&Eu��Ƒ�h<:��Q3�4�ڙv���^Ŵ��_.U�V.�̽�v6��S�˃,Ȅ:;�'��Jo(���\�@C#/������i[[��/l�B{4�%A�A��6��PtC+��2��r�JZ�]a{ڃ_yj>�M�E�=Z������E�Ʀ��F�)���k%�[�UØ���Q�3M��Kސ{m��.0p�].h(&z�03�����[���sbT�]H`�O�kt�a�iv޵4�b<�+�܆��Kӝ�D�RحJ8��z��l����*|U�9��S瓅f*�bFػ�#cm1�ö�ە�����ۉұk^�Ѽ��}�cm�}%���)N0�*�B<���;%����*�bP_B:��xL�� 1�e�5���ս͂��%-�+���ĺ���n�S�y�jV�3��q]���}V�$�m�+/����1Mj\S��J��aBK�v�qT�b5 �Nj��q֩��c���h�䷫>�X]lq�zVX��e�tys���Dd���A�j����gkL7����EB ;� �q�U����7[7���ޤ����[B�D�{�����BhJ9hHT}uu��JL�靵(�C���v]ʺn"��*��mg85��.�t��`�vI�EfJΧü��*��ɂ�2�`w,����R.G[�����|P���;��G���`�tr$ U�&i�Pb���sܥ�2���ǯ.���I�L�Q�R��m�)� `=������.�
8�W8y+�ѮJs�4)�:Kbī�`]��qu%\U#��V·}�;g��<��aݒ�T]6�����
 V��G`�H�"��	�ه'���Wf+N���]ZwJg�+T����y���a��Uy���Dj Q����WG��XgȞ{���a� �Znͫ��`<m���ݵM������\2��ʷs$�7w.'��I�]��0��8>V�t�(�n;=	j�eD���oJ��vm�b�5�.�5*;���Rw�C�+���oL���L5�8��W][`�n�vm�ҙ���ʅ��yt՛X��-wHK� �k�U��׃�m_q�=}H���e*�"�z��*Vs2�ٖ���.nc���@^������f��������sl��1ev�8�[��뫑��rܙ"��)*��b�T�����kd�D�Vm��e]$N+�2��J�o+CRz^qzJ�l����� �R��.h)l�YX�\��j���,/�L�L�Q���cWFuفk�ә�6�l��Y8dpm�СQ嚊�X��AQ�YP�J��6а"nm`��ťtL�Z�ҫ��R���f>��oF��3mw�v�1!�ϛ˩�7�� ���K�R���Hv�v�a����wN�JT\ĵ:3���7c�lKL6�E�ɡL���}b]e9���s���$.���_v`��.��6ke�u��T̘�ԫS�l[`2bW8'��|]�X�n#�3xS2�ś*�]���\5�|�v����T8��/���O�gE"�f�+�����
�mo8)��yB�>*����GQ޳Hm�+�1{�5R#̈f���%��l����$�wvTݔF+�iD	�(r��t���{FE9%�[���ю��P>��m�
]�
��&FF1�|j��@جZJ�7����}�f�وg?VлC�r�v`s�����兖��X��2eo���gP�}�l�]�ߊ���[�I��Ɏ��z�VXE(9��9t����2j
��d�"J,1�zi�v'%��1��O����ݏ���8n�\�����2tm����tZ�W%�z�W�R���z�-E�t�=�qj�b��&���k%f��4�N��	�U,���j���W�;E��/�P�  8N���nn�Y��_���\t����WyH�N�n�I����#c��^�F�P����Z�GGd�(�����-��n�.�mdvM3<,Jˣ	��M��.����bM�X:�=:!�ݍ
mH���MsýNu����\8��N�7�}�Ν�m���jRab�sk)֣�hX�໳�e.�8I	һ=/U#R�u�=���6�?H�#Ti�I���u��ت�S�/v&F@�uoK"�\���MGN�NԬ�n,�������u�]��R���ꖤ�nB]aJ��=V���{6�Zi�2�m�m�7e��*�p��h��^�\�.�4���[��q�t��qc�]��eQPU�[�m�Ù0г����Ⱥv��e\�"u��W^A-L�sb@����L�ݼ�m�3'�Ż0�\\�>]L�KA{�YK�8-l��,J�8��2�KT����$�]���Tc����2��]�㾥Wz2�
�3�U4�ꥁ�{Z.�d�,l�Z� �:�v�j#\T�m�0�$�%��'��l�u�w�����ʇ4�{z�Ե���x^S����3.��u�#ʌ�8�K�a(Su�p���aPeԔz�ݲx��^�J2lr�Ձ6R<OyM����p�u����כO���������=����}(��u����J��B�13�ٕ��T�L?�� ��S]kT3ZsD�1j� ��P; ��rDv��P�n>�c�.gl�l�\�6���W=U�g)�.Ύ�׌��m���U�����6��Np�`դ_M�+	��|�3kP�F���=�(���z�w���QKi��V]��vːV7K5,�K��4уu�v,�����3â�BĘl�.��x�v�sT�0vPa��2�1V�\;P��!.l��i��g�k����Y�C�6s�Y�a�Cq[��kyR�i�%�J�wף,�ĭ	엠P�=3��}s�@�ޣ7D�;���(3Zyi�e�����4�Ȩ�f�쾦�N�ۜؒ;ɛ�d��t��fWEI;U�.�r��u`��A��H�����,��/�H�|@m#"Ly�-f�5�-ۭ{��AZ6�
+��C������$#T���z�����P���I	�U�&b�	_l9Z���7jc�ʊ�h5|~4��AC��R�4��=�יp�i�ŝB���*vm�O����|��9��K�%��%Y2�q��[�F�6�hX"'P{S�ɝ�e)�P�Y;�3*'װm����,��H^�qv'�R�\3]j�e�T�n�R`�6T��N�UeY�Z����tk�WKHm�(.��رlfK�V�a �b�r"��UG]��]�Ҩ�,�ęt�)nʽG�yafL�6�w����sOrj����;��7VP��Wӥm�>���$Hc[�8�5�u�o��r*sޭ�ƹH�u��k�5���.��r�sd�~�Һ�6nNt���F����S=��G��f�q`�&�&e�.�n�WP����`�Tou
�Ԛ��}A�������yoA��m�t�ކ���+;3���g�Q:�����&�L�� \�Iy׹�����-Y-#�ک3m�=��T�N��R#k��ov��v���y�aok\֔����(�X�ۡWo*�'�����ٗ����Ӑ�r\Z2/%��'2��R���4�ԉ�s�\̴�ّ�00�͔NI�aT��8v����1G�_��;Èkr����,�0���T��:��*���"��*n�Ѱ�?7O�Z۩�@��4�U�ͭ*<�V��gY��	��5�;]��.�[B�b5,l�#��8��J�s:�&u��L[d�u��M��+�>4��o2D���Y>�2S���3o/(T9�%-�N�©�N��*so��Qp�n�����\抺���{	-b<�"�-�0�h]�dȳY��]or.�s���Z(���y�eI�C9�_R��J;YOa��<�Ci>
i�r�����!�3]A��8p����;�^6m�ZQ���*N�k��;���@�j��t"7K���"R:w.�ӓ�s:[ͤ]J(b�&�1W:�Lc"�*�Z2�u��h�������&�j*r@��Ṷ䅎��h�)P�5��'�N<gmviˏ�Jʔsp���k;ħV�\��O&��OW�K}�n�tjޭ�0����Sڽ%�|oEW=������ʭ"��۶�u�|�̧��ڈThm_K�V��Vԫ���[[�����/��0���xV�o�d�vDSB]am�a���󮞂�5)k�o��"���
�0V"���`�pc`%kLC+3kW�3�����ƮpQ���WգVM+!�坌6�to�^=O���R�=N���r�z(^kL�
9��z�yӶ(R��\���Y
��I�}1V��k�����I�ql
Г�RBGJ<
R7�"�Ӧ�yثGb�d=�6��A�a��㬷:h#�Yox�6�[J�r�/ڢ
�R]Cm�SX\�<$V�1ڻr�*Ծ��9��T�Ң��r#z��s����v�#Z���A3M�[���T$��N5�Bg�%�����/���Lx��sgk/�ʓ�P�H�34\te��c75J���4Fu��^n�{�m��Z]�8Z�������ܮJȆ�FNV�-���A�3c���0#&�Вm'I�*)�>�._ǔkFB��2˶T��m�V�8�мt�>�&%�ok��1�Q,dC��]ܗM����s�����g纤��b��t�lr��a���� zok�V"W�TW.N���Wעz�=6ġ|'$�U��HV
V�5{*�h������
�4T���yQОZ����wA�[�d�����AMkX��;c]J�l<}����;���)-��Wwj9v�9+@�C��:$��pW��:-J�!�}R�oD{ޏD{��{�{۷�\i�L3�r��2\����4 `��hK����l��Բ�\DIQ[Xg9�7�ڽX΄���I{t�^����V+��ѝXy�L}+�.���A3�=g�O��i�F�$m:��gd�v����9�p��%4�|���a�۽�-�x[��ٰ	���J}RKqΩ��J�2�>P<����[7����Mp�+@����b�ϥw�:��%c�.��2�	�T�#q����,��6S�s#��-m,�i%WS�{G��d`�z`��9|��J�T"�.`�F���um@"��-;�SQ�הԮ�4D+'gf�0F u�t�ڭh�Ů��'f�|8AOqJ���8��-�U�J�N�vٔ�����7�W\�W��N�{4JX�N��pN��mf�Ĥ�V�T���TƄ�=8 0�Fګ25�Ʃh�����39]*]"���+7 �il7��U}��5n���;�Ǌ����/]�WGgL��qce�=�N�����{�M`�-N��C�FԸnt;��l��[��늕u�%s�mnݘ�쮩�Q�\OV���żw�0���f�-(�{u�j�l)p���NW[e�T�-���D,"0�V��V�-�����с�:�♆od�w�nϹ)We�kf�h�8�����tޅ��MK�'Y����M�EgIRu�ל�]��"�R�j�b[Н���>�I�M@ 1�,2�H�j"*��*�&32bj�Ɋ��ՅT@IXfCF�4ALUf�`�UfQ$ELZ�F��#0�	��V���K#"Z*
f���0�b�ck2*���������s0��s1�5� �fk�#,+S�TTUQ,CY��6�$��*�'Y�TCAFZ�fd�TMPMi��Z�QQA$Y��EUY���6X�5d�f`QD�QPMFf4e��eUY�55��QK��̲ՎA�e6fF�
*'0ª5�DS�eI�QL�QDFYU�1��kg3*5�Ff�VMNU�UU��A3E�Q��jueE9kXNX�FFDY�feYfe�g3
��ak�
�i$��ѓ:\�X�3�.&vV+|�#l+�l���s��oy����WO�-dW�i�Tv���i)]���fmA�y#_5H����MK�NB��e��,AF�;P�}u�m�_)�2~=���k2�o�ҧ'���ɅD�_�"��E�=��܉U\��R�mY3
J �[��\Ka[}[ݩ${�|B1�{�֧s��z�Ή�'��l��  ˙X"���C��Y��(�{��%����5��w�����1m+���ӌ��1�:b��0�	�[��4�]Ĕy�qr����U�0��(�8 �.���|.UZ�9>��>����m��;�<�qK>����a�o��2w��@��x:�-�2Y�3�kJ�ᴴ=R�[B\>����sO���痗Su��߀s3��fe�KHC�)O7�Ԁܶ����/�U��͢�vm��pp�j;��-���.�&5�g��Y;F</j�;�Δ�͗m�#�{ݯ2�on[�OAwA=iE�%���	�����Z�0�Q��P�>�V��L����K�3ea���e���{�{I����r�0�%;@�֣GT�d]��k���O!�\3�%��=5T�T���fJ��M�cR�ݎ؜�p+)Ѝ����YyF���Y�ppK��<�ŉ���poWF�fL�\n�9D�2����9�CGX�zVP��WG�.\�^K�S;`�3GMS�ޗ�f-{ٻ�؝���
c��a�կY��bvx�l��᱒(Jޞ�����\¦2��qt�	k>����6$��{n�e���X�En���/����[����5�m��{j|[�����k<�ڪ0��O��F˚n�<��p(M��cN*o���n�	����e.#�)�2�C�6��	{Y���3u���uq��P��1<��Χ�Ņt��k9�+"ҹ\Z9xþl��	�s�W�*�����������f��K����R�T�<
g#���O�-u�%\�\��qr��E�l� �u�eų���]��w�����o��C�!�8�x�L�~�Sc��6�SS*�kg��aH�VL�((���+QY��;-��\ �y�J�.���k���β&׌��c�����T��q� ��7��㶴f���,ߔ�g�����]�c�=-<|h�o@�b�':��ݦץcJ�D�8�F�����ڎ@�u��\F6�Ț�-ħ�Q$���4�f�7�ĳ�[ _j����ݮ\X�cw_���{:���5'fE�.׳E��;[@3!:v���Y���|�78�-^�i�r�J��x\7**�f�P�@�9Zř'^�p�U�A��g����#n�8j�=�r���Ght�ylU�4J�	�#����zV�;�~T��ޡ)/2Ϲ(�����,�g����<�w����ފ�VIQW��2d��fb�B�+�
�EPڝqܙ6�}
:�h)�(]���Oly
vh�秄Q?D�j(e$d�K-����{��7�/fnu�%����Y��(/E<-��_edL���-�P��J���D�h�4V�نޝ�lX=Y3@|����/lBR5�/�Ŏ�V�OU��/������T�z�G��Ⱥ��=��UMb�	[�9)T�@}�_鍔O�`8|+U����{�������W]�o0ݗ�%�uĕ��M�ay��;�VT�m�;�P�7<��3���5)�]׫uk�;p~�x��|�w����P�5�	:&ʲ��V[U�ˤ��1[=lMn�W��[rT�n<�:��\�n�K ��0-�	��_(�r|�}�=gÔ9��	�bT&�"����%f_m�O,�݋sQGp�k$�ʭ\p�C�o9�k}����l�g�G�)s��䫽����?%�9���ע#��< ��C�r�Z�.f�)13�O��I���
�����ժ}���3,�5�2��}��X��܏��A�����lT��w�=��a�v���]�;Io�J��^J;�y�q�1j�rf���PVT�A����(�KvH�{�E��`�OM��V,BEu-�ԍ�Y���S������O.6�N��K�s�NOpV�ꓤU�V�	t�?q�
��FD�zL�8��>�N`dX�z�v���U���n�g�շF届�Sq-:�y�r�
�����Ue��0�a!�)���!���t��Er��f�rq�N2��>O���V ��+d ���%L��P�4@Y^���PZ�Y�֭�Nt�\�����Y.7����L�չ��Q\�86x��KrI�斴�����ϼ��x2p߇M�o���b��ۮ�i,F�=�LM�P�5���s3+r�wg�.��s�r�Fj&�<�G�^=�b��pٵ�Y`*�Uזpe�G�s��k��H+�����Ra`���;���S����=@+/A�u�6�x�Xz�Vl����6��#�n�J=�R��r��Pu�s��\���l����
������y��s����D�u����Â&U�S��&C�5Fu�F7�Uϫ�ox�"���r�X��`��~��{I�cC�t(_nr�k�S�}���M��N�WC�y
�M�e�o�6w �	s���Ĭŀv)|����-�����R�{���Pj4��P�1��
g��Huv��oGN�b�Ru�]v���	�_ޥz#�L�ή���8���uS2*���ۇ;������\{�խ�Vs8��r��\�o�b����ܪ���Y游�����<��*���:� ��K�'&̼ɻ�>+B�=�9���sn7��rUf�3q��L�b�Ftʧc�y�[sv��cz�{��I�n�t8X���ܘn�ĳ�+�b������s\!^�&�[��c��qa�=���rm�����u��k��xF�C����x����D�1ktu�9[�/+��x��R�77F���}3���x�\W,7�*��\v����W �J�z�p�ܞ�A��1'8�p��aѯ>�[)�_��܉U\��.uBڽۗퟭ�X�*��\�Oޫ��Wz��9I*������B���ϒ��$��ݾoh�g�����7��n�p�s9h=�5^��giq�F��������0�m�#aچ�sv���י�����$����y:�:ҷĉ�_��JǄe�v�.u9yZ����N7�%i�Wǂ�KN�,ƺ���������n�������fm�?E�ƻ���`���ɧ�A(�'Jz��+�Ÿzچ.�z7\:�>Ll�I=$e�hԽ��=�β\��ջVwY�a��3t���vR��D,�JJ\t8�c�}�������ϫ9�)dE!	vu���%JHu���'ت-��S1;�׻ǔ��(n+�yN�+�^o�9g;���^$��$�L���;��A��[5�ԉ����fI������2�F��XD�&�U�X�������H#�ޯ�|�*z�G�vq�K���ow��l:^�s<��"��-(��^�F�-��H�ĉr��8�h�c�/��|�;7����8�5����,i�)=P79PU�l��	�/[��A���]��d�sCp}Y����!��f�k���[��N�	�o�|�	���V,��ߤ�����L�x6�\�;�$�����UyP:̘��0}�ʛ�U=�:���L*�g6c��r��g��{|MN��.����MzS�	�bi�|g��p9Ӡҫ��+޵���P�M��iα��r��8����4����*M�3�n��u�F�!}$�elo�Sˁgq�VE���2�s����^�X2z��!�zunA��y�����{h�)�;a�Aʙ��o���a�í}��:���ڇ��^b|���&��\�\;;�2q�E:ܝ��;SB��M��:\&�i���E.CS�"O�lݜ�m9w��0��c,���w� �"%S6T9��_�v�v���Z�S.���Y����tP��͢�I2;\�P�d\ws�a�M��F�����2�-6'��+�dɍGy��SV!�G���*{F��%+�,I�x�i���k"�����6�� ��0�o���g���3��Ky�5*N:�'֩!M_+�����:�;�ĮQԷ��2\������.�8��#���<��_aڦU��7E]/5�؞�oW����s���jc%`x������~�qZ�  �ث@^>�BaYںe&�֩t�������xp"����L���'�}�2R���xߍ����@{Ҭ�(�<q2i��8�]qV%��Hl���h����
��e+����'膩b�iݚ7L�*�W��p��{��v�ܨ����i�=i�\�d�PY;%�
�>�T#��˘w�9���y��oy-VOp����D�"������"5�,1c�}o��y���I��Y�5+�dby9�~�����6ѫ=Ց�>~*u�
�GI���x�1�F��<ٗ�6��x�ګ'A'��5�&:�%0;g���/#Sj�u:����xv�{�la���Oo��ϣ�'�	�X�nEys4�
�۶�p7�Z;�V1(hDM=�%zu
������w����e����qX2$��:Ky:!���#�9�]���k�˕�q��L��a�Ё�v��t��e�}ъ��u<F����:�A�4����ʫ�}f�e�=��q.�F��fs�eY�mYmW�.�[�#��B�.l�y�m��'H�i����++L;�]�{�\W�>O�W���τ�1*��=g}�L>fN�����d�W�g���`�Z�s��#�a��6X��`�jw�g�F��_BL}~�w.����	�Jr�Z�.gbg�1���H.=A�yw�J�%s�]�{;�xB��>��gz�/�)��a����8�A��I�'34Oiq����UV�<u��#0*�M
3�w�2�u�%�x\�a�&."v�F�G���O	�N|�b9�ǽ)����v/��y�/�b�+��/!�u�8����� 3�J�>�
rŷ�(�Ë��Y�;��%7���v�}��$vxf�E}�zOBpc��mNu�1�)�r�f��=��D�+��(8�,z�v���J߇=��.>!S��j��چ�le���qIۜ��x�� ���'�#5X�����(�P���,�ȻP�
�r@���Ot�u�9Ft��Db�������}�Zޘ5�C�ѣ��{���[N��й�E��4O;Ww���udt��bN%e�}İ:�l���W�)r�I��xa����O7{(4v�^�%oQ]�8���8k���w��J�Zn_K�F�o#�rP�����rWK�j~��<"Q�o�����/)�� ^)���k�M��fbA{�W��J��9�b�&�{�^�<�W&�����z1�-L�~J�}Ҕ���i�~���6��k�����Dl8�3���uST�JP.^�U(�#~h��8�vzj����N�V�zu`��ӛwjl�y�-�s3j�p1��>��H�d���ŔC��Fom�4z��x�#&�����}\/�8�W�C�2��{Xv���T9TN�D�Oʦ�*�j���87n�՜�q5A��φ�.�M(��6�������ޏ	\�X?e�a��_e{̚�*8K���M7\Fu�'V6�M�E�������])�m�S5���ª�d۵��������Ύ�V������������#� 9ާ5iO�#zC�e�f���e�Į͎j��65� �	��
�˛�2�q7y6�;��k4S
$!����j)%�PT��Vs2A���5J��>��b1�b�r�L������:�:����$SǼ�β�CֆVKzC�׋���N�C��7Oa���i�It�l�{���v ;�˝��������^֮�7��{b�N�����<�y��|#�Z���ey5]���\��4��<�ԁ��b�n*�]�p5��)t6VdU�S��7�QY	���3s77���F�p�(�r����R[����#�_
`�ϒ��ʺʑ��M�ɹ�Ս��R��+bà�OE��%d�񀧤ɶ������l�R�/����Q|_��D�u��Z<�A��t Ҷ$pkښ���,��M���9`K���jF$>3���)�y��gNJG�;�P�u<��i���5q7Ë�`d��7>p�h���t�I�)�1�q��;~����WZ���	_.���0\��`yJ���;]<�f���Ŭ�f�t��uoK�9aq��YiO%a�k��U�{̘�Щ�V���Nc�8�>K�fM2J�b��r;;+3��)ib�K�{�w`W.�XZ[�X�rV$��n�m�����'ڙY��<�2V�~��*y��3�����5�'�c���%��
���%vzE��ҵ�}u-��*�o� (�ȥ�����:yO_7��z��8��+Ip��B]�����dǎ���3��1E�v_��<�w&<%p"���� ,�P���ܔN��K�ٺ�Ļ���)Z+o�]��N��Ph�n��v^��9[��u�E<Iᾩ�N�89ݎ*d����\\o�� Oh��U�l0�x�!�7x��۝����_t��(���2�j�e�����ႈR�]$$Qn�"��2蓩 �6�Cn^�;���a�ri� u��J���h� ͋�\�=YղJ���!Rbn.j��d�{����*f	]P,\h���9J��fr��.�;�y���ޙt@j�1������v��fQ'N�u�[����0Yϖql���j�HʠU��sd]iN�]��j�1/H����]<	�Q�8+\�;��;�E4#�C�FL��H�Mͱ�x��ܝ}ͪ��TjV��W$���[F�Ѯ�1h��=f�>���մj/��ҫ1YW�9��]�:�^��������޸:����V�u��1�ׅXr���9g.^b�u�� �gcYM�\��5ɨ0�e���s����)�@V)��Jb���Mh���H	�������M��Jj�ݳ�f�=����4��o+8����eL���9��F�&m
}��;Qk�X⩶�y�歾v���`�U��p<���g���n���-���G)�C���$�N�V['uh�R� n���ܔ*�Co`!�I��X��7T8o*�7�u���[�����1֙��M��3��W�e��9�ʉ�U����r���NMEoE{,;W��N`��xgWDsA��j�8�*��P�NԱ���`���Ma���mRc�9F�X�Q�J��o8��R�vĕ�� ���&q�K\�K��c�Fю��f�r�[�!�}�q˅�L�IW0A�������N�k�w���c3��&�LעL\��[���N����	�T��z�>�P|��fǘ��[4����X:�n0�&�1�����BE���9}�I��.�^g*wS����ȇ�d.��f�6��yu*�fM Fi�&vj0GT��Q��ꊰL���=�ͼV{��� �M��,��qt"w���4��F=�Nk����J ջ�V9�T�E��gJ�k��C�s:�_7�.E�z���e�y�79+�W�:��o��hu����I��y�M1\\���2���ʺKb�%`۱f��P�B��y��Wfr�1��V	}� �i侾4 ��inJ��QeՁ;舂�q�Co&�w:f���y��p_+Z	�sa�(�����=���a����=��~�`4>͖c�G{t*O�Y%�U}��q�YV�ۧ
�EO�����!f��r��R(�8L�mҥ��sjС��j�`S��)���}�3��i��qwH��/�&VC��Q;q[�0
���j)������c1mNBoJR���v����dh��b
�,����+0���dfaT�a�ִf�Zl�(�2���-��3,30�03#�,2��p����̊�3E�� ��ѕ���Xa����%$�D�@d�e���FQ�EFfU�&kQ��������"��5h�Xd5QX�LU�CN�h"��-F%S2X`Sf48FFfVLMS���aRPd�Y�d���fV&-PSa�9�fa�dDj5QF�Ƞɢ&�$ȫ2"��cXaUA�̜��ʃ
�r0��2���0�5�54Ra4�`�NUba���&EUfd�%T�bd9�6Xի ��Qd��V����,2,������,��
2(0�r"+
��kX��r��j���k+*3
")2L��u��
��Y9L�Ƶ�&���Y:�*�"�#*�,�r��1�**��2Jr�3+0p�Ƞ]��v�qB��CS���}���ʊ�o�c�"��gZ��'۽�sk����1�t$���ʨ��8����%]J�=S��IW��g]�3S�Q��gK�/'V6�,:��l�|"7C�����K���,���	W�H쨼��s�c�\���.K�;��͝�S~iC.EIeE�݌��4�7�5%�$ҩ�> �-h#��2Vr���"�F+��Y�����X;3��*Z��+�ͽ��m�CD�>��$f�o�c�������������ڇ���$=�Wf���/�nvL)l� 4�,�K9�d�be��1�9	�J����	5(sp�k�;�-Sk��r���T9mV����S�%��g����ps�`ǘ�^ɱ�*���T�P��ۮ:6�w������x�W��1r�����d�ڤ�4�X�͡	�����F�D�p0)�\�I_y�%�7�ں��]��-����z���^d�)fk�0C� ������[*���J��dɫf[�9�蹱w]tȿA��ڪ���Nud��l�4�Sʾ���K:����ļ���-�#"���k��ow*�%\�هgh�+^B�V�eN[ίn]���|^lX�X)��1o-�3u{���}zƵ���-��!�(����kr�7�7,ǐo'���n!Z8j�v}�EVY�=*�f�s7-3a@��Q��uW.K����'9���b���Y�^���Z';r�&hlx���k���~O�Q�p�\d�%N�<��y�;�"+�k�!���6�&��h�_&�u�V�L���{��Y�I�o�wPG�d�~s���EM�p��c�,^�5]������G��9�T��Ly�	)��Bk��?D�!����t1(�"�w3�p��3�'�m��-�W^�<2�
67�.��K�*�^�mYmW�e�kAF����C�G/��ǆ�KBkt,�8����P�j}�x��O���=gÔ��]h�w2������oh��]���t�]	�ߖ��^}j�y֥��uR�Y���A*p�J�D�����%��P��s�Η9;0�j2ט'��j�l���eB]����D��z��g��I+����D[dܾ�Sb�x�dv���l{�\FZ���N�u+j�r�;ˌk��K�Νv�t�{ζɟ\xB�|R�TnyN��i���r�NL\�L���v2�3��qm'_Cr�3;8��/h"~�5���1x�a.��O��ft*����nh��с�ۋ2�߭��eov�Z�	:T������j�n6�p�h'�*%�u��g�^ 둻��r�SV�'-�{0��IAd��,Q�=����\��$|��<H��c��\ey�S⥹U�k��8)R Oȕ3�tjHԗxM�y��f��Ռ�r��U)�;��0k����6�u����[� �{w�5T�a�A��w^��+�v{��6K��rG��(g]\�K�6g�1}�\���0.wBZ�06T��]sm^�Ϭ%�{���2Zd�|����yP��g�q�$�GXPb�a��F�&�m�޾]��mm��M�*(E�+����o+���E�@��t~���W6���Z��9�^M_J�()���"\��*�>]�1�����F�{������c��D��G�_%�s̜��� �UѬ~�STFĥ���"�aEy�u}��c�j����úu[��Z���_�[�T\��k#F�|ct�*%�ه;P"�����b�_D\7�"o���#7�}��6x��O����Y�~;��7���_d���v� h�o*�3��b�C���E!'����T
�8�FOp�|��c����Xy�/�W(r�ݏ�Q�C�)'��g�*Y|	�(�0^�^�IɷN��(�>��v^^l�W���F�e���fc���:ư�:yjlj��b�K6�W��y?�����p�]�/��{Y�++b��.W
���%c�2\FQã:p��X��%�c�c<h�=�������h���o��`R��m)��|�>�2���ƌK�*�(=o�)��d~3靻cp(s[��Jv��vk�/45�����˳K%b�%�K��D�]\�˔K�~M�M��慄��L/HCg.Y=5sp�;�v N����WQ���%!s\g3c�)-�͟>�]=�m���H����j��7�v���ݽso�*\�òf�%*��f
���E^Sn���,������!��v[K�J �_$���j{�Җ�����v�4hN��{��1�>{���u�v6f�{Yh��N�J80]\�2��Ofd~�tұ�cC����Gモ~��;ݫ���5e�P������*����-�:�9�ڶ����͵���A�������s�qL����P�&���Eޓ� ��y�=�d��l�����jJoќ[C��C�2����ʆ��YiO%a�>;Q���U�.�&5�����@����;�ɞ��t�)���i�v��`��������v�>nQ�\я��gy��`�WgL�F'&u_��<]�.N�<�ܜ��u`��|�f�����:�I�=gq� ��q��C��ӧ�r���X�_m���ۼ����]y܎�"vP��G��g�p,n�P���,ڳ�;��bҧ�tZ\�fx�KGL� �V�52�;8+�9fG��m
��uK�\{�h�-�գym�}7��@t<�.��m���0�t�u�\��&'g��+s�<NKk�^KޭSz������b��V6���<A�,W2c�]��,�c��(��OV�.V��&q����&��3�]�Ս���~9_Dn�n8�Z>�v��=�w['��+�?���ڜ��Ӈ"��;1�3�{Y��gxT�H��*�m�ꪩRMT�im��s�}{����%���C����M�B�R�B.z�󼛇�F�f{f�tB0Q��3�o=��BԪ���V�����7�]�T��]ܹ=k,��dN�3��)<������N�nrJ�,�|#qa�ߢ�U�d�S#�yu;��:!fy馎����Û~�Ů��'��YP�;� 1q�q���ny�Eb�ْ�<Ly�oz�7�`ʦ
��=�qgN���ᬦ�5��X��[ϖ�
�Z+r����X��ò^�E1���v�E	ۓ(�cvV�A�nm:Z�r����Il����6̼Pr�O�A�z�m*"rd�9�:�n�Vi�[9��r��SWU�ɛ�vM��:�ݾ�R�������,~4���z=�q����8��u��o@tAc�Mn]��j�s��G��&�77!��6V�M]M�_���}*����Z-\lї~�{.��ݸꁑ>��R&�_�x�s���Q���_ӦJR��O���5::�-M���Eݙ&Wn�z�'*THt��k�Ȱ�}��I��El�4�JyoV�hd]-���4�`���.���܂��#ޖX��xQ�lu�A�� _o�u��δ�O��1Sc;.��8��:Dt�g�]g ������ғ~h���5�EzX��O
����6�����ܺ1��>|Ը�'_|K�42Q��:�6�QS��w�)��8AKՇRN����{6�w���G�iVFLt:�%?�g����f�4�uYS�fc�N�r�ߏ��-�G˗y�b�Q���c��֫�P���c������K�*�^j�k{{�E5g�빴��ݵϯ�_����F��4� ���!����!�\W�'����]�=RߧWJ2����RDp5��BN)��7���d��q,Ҋ�\�
�=Z�;q�G4Y�y ��`�e��6'3d�)#�Y�9�Sײj���X��41��m��h;�eD`ehk��[��^�z�B3H���A<1@�H�u.��������%Aҳ5����t&��WvV�u��P�T�x&�~XOO�x5�X�s��#���uF�E�]�6��ݵ��J�>�Kpw.�&R/�v
r���q�ht�~Z��7�f�|���"�ڮ��U\��M�숦�)0�>��vw���1��1��tu�#"W9'����^W˥���z����=�̜�S �S���AJTKN����M)���Q���%�U�v]X�ҭ���cX2�L���Q^hO���#�ds��9r h%�s+c=�󗻛۴Ƀ�߇0�����C��*J��y`���N�{]�HP�7YZ$	��JyŞIq� �g�#@�V�#������%E�.�X%N�1W=���f��7_|�|~U�֝ف��ވK"��bbR~�3(�	|&tmB00�{<o��˨<<������������n�SSqN�~
��-�䤿�*�y��!b����n���`����뽲x��C،VVg��Ί0В�C�ޣ��]���ߏY�A���$��{�W'���/$G_l���e�CǸk��i�&��n���,]�;Ԯa;�iu����i�=��l��(��^7bv�u��ai`A���X�Y5u&��AO�����iv]�����;}���m��L�il�ή�gZ�)�-wsƢ�8�<*��T�$JP/�/�Ȫ*Ѩh��8�u�l����]M�[	ѹ���|�}^�NyS�8��ں�owТ]8��@�0���<�S�;g�A����k����D��Q��]97Z�1�Nt�I�wu�*
i�K�ټ�#�6�7�n�ͽ.;�
��T�>9࠾��9��+%c����]�J��8����$�5�t^s��z�3m��> �̠�;m�ݤY�x�	ע%�Z<�f��ݭ�s���{ )Z��Z���Z*�c���Ꮩɸz��79��ץ;~�!����)����>k8,̻��RUP>�C�w�H����n|9�0厓�|&t�����N++��x��7�d;<۷[���o��.}�`�s��r1&1b�9l\3g��3�ڧ��5t�J�
{!¥����6^[(��:
0�Sdq��{��GX���}o��~�$~V�Z.�xN~S5J3ѹ�V�b� �o�����>�)��rDm�G����Ұ�-gՖ�c�聨|�*e��b�v�T�IwU��\ӋF�a�8kL99,V6/e�ص�N�8حoc��_G�S#i\*)�/]�9Eh{]$�܉�).ޔ�DT�v��G�%��k,�(t�Uq��ef�e͸���i���y���:���Fۑ[��'_���B<[��dkV�|�=�1i[�Dկ�m�c�4w7�*b�=w[�r��ά��|��V������iϺU��=������w�Ӯb��n&�h�����Nχ)�S�����s�ac��g�Ce�{|��U��Hꒉ2?l���a<��y�o)U�u�ݞ~��ҫ���M�~����,����x�sqL�c<�B����C���|������qh�68�ՒumF�M���Y���ZX���݊��s�U��)��˸�VMW�f�uAr�Njg��>�<嗒��Z�8̫?P�'�5�$���m�_��7��Y�-td{o�S:�l5k���*wEXRrQ�%v��V�ֆ��{Q!A���M	�_��Xۣ����Ļ'�U̘��@�sF�q�d�[���͜��s8ߙ��]= {����<Ix`��~X����_�r��%1w�;���/���Ճ�a߽��Nu�|K����<�)��(<�Oc҄ˢ�J�Ȏ�{�
�Ϝ�x�H=$��gƮɉ�,s�@�i�:���^9���y�Mxo��U�T��f��Nb�u��rH�U�0�k��儩�x�����V;q�n���ۉ��ا]2Wǥ%6����}��f�|c�=YE�W��-��MxP���PT;u�t�1��.\��w�Y�;�-����X{��.������0�N�K��G���_���ծM�A��򥧻��p���B���;��V��*\������i !�1dK%��vN1�9S-�D_��$d��")�\�W����>C:>k��p�[xO8��[C�ը��C�:�P�n{�ީ��R����$�ۘxߐf|=�b~��P��#���%����D�x�ˌ�EPa��u(;ȗ�.�s�{�mU1^�6V���ߥ�(\c������"�,�VkG1;�g��Ŀ!Z�� �ڥY��{�	GW�A+O�s�JR��[��K*H<�pMv��3#F�	����$1Hv#Q<��
�]�s�'�P+f1��I;waJ�'��w��;Ϯ��O؁��C)#'�Q;^N�5e`�0-�gVV1RD�7�g]�e�۰��ێ�gx�ه�DW���2�\iriI��GM9�g�4%�����|yl)���7�jR�G���u6t�oA�w�����wZO��z%��|����Sm��7n�֮
�x�R ҹ1�F�����G���%��nwwU�-���e�b��$���Ɍ]�!h*Î��2�G�ar�Aܴ��$��Nuށ*��n�	t�ͨ*]a]<���&Աl���-5�F�����F���n˅�Wf��LZ�a�Iw�!C�����G+���Cic�K��G�f���)Q��/w:mdY��3�נ�n�����q�3�g����]4�������5�&Q;]yCtl�&tX5ВV�ne�u
�k��6.���*TFۅ��n�&8��ڷ�ڰ�e�c{b�BM��A�ɢs.*��5�<7iEbn��j
�+�@nG��UçX�_u,&Z߻6!H�����Lީ]VQ;Ck�Җ�<�p)���%�́8r٧m��X8&�V@i����3�oF�p+�X:i�Φ��j�B�ۛ�g]-�޻�nCXe4N�Ы�엏#L�(�-� @�.��d��^���ҭ���@=��Ǆܚ�)��)���󷣇�{a&��H�N��ٙ[#{�y�M��m��ۧ�`�=�86��me������]��l+΂h5zҬ�μgK���+ b�S|[U��.��I���5n��a��lFd�2�I��E�r�N��g��ƴ[��BkA^�`�-B��ʮ��0-�`��AK�Í�pm��nc�g!��G�)�]�<�y��7u��d�3�ֈz*���%@�K�$��s3J���t��)6v�7NAX��c�8Ԝ;2�eZz���r������'�:I�c�ᠺ�ͳYU�V��e�c�d�{emuf�����/��8�H��|��Y�ٽƀv^�:A-=�w&]��J�(><0��3���çY��M2�qEVd�s�wm���t�Q�t���ueٜ�-="�yk{b��6]Al��a7�X�����h rب�0dߥ;�`B����h6x�NoYcs��KJY����P�y�9Y,�tob�\��S����)�,�%����L\�`��=t��A�K�x*��šu����6a6@���M%t(*���t.M��N���o%�a(.���?w][#�c0I,Ӈ����&�����R��z�C ϐ�b������ToRoh���h�i��n���Uw:�b��q��%/��uZ�p�vw�[��\�w9��4ru������Y�|�RS�F����c�;��,����kec�R��r��
�K�_�R۾Z{t��U-��;��p=�/��|HT�8J}0|�wx�"J��lGMK�e>;F�I��Μw��Eݫ,�g"��U4�;+b��`��\��w77����}w�cn#c�n��,ê`;X��:X��t6����#<��{E�eu9wo�<��3ߪ~#2̜�$��-Uf�"�Nf4FdY9IT4ef�VQ��VfY�VaY��(�VA� (��e`�K�T��l��T��CE�5P֦�b�)�3Y��ddf�jueIE!��Y�V`N�֫0����sVZ�$�kX��E�0��`j3,2q�r5�Tdee��U�ddeafe4VCfMS��k�F��jb0��p�2l3' Ȱ�`�0�h�k�J�"u%�c	��PVa�Fe�Fk5%Z�&�� �(�V�UE�E�XfFY5�U8�FVQD�f19MXIafA�dYaDVD�de6Tc19ՙE�l0rɢ�����\K*J,�03l�"��0���*"�ɲrȬ��
�r
"�,C	�&��0�Y��C#*̳*�̈�����
�@U�'9����n�2�O�H��V�.hvk.K���')p�;�u��7RhۉF"�@ތs�t��r�U}��k"S<}�^O9*9ɵ��q'@s����C%�3�ď���0�b�|�3���G_���z�����k�6������c�x����4&մ�uYS�ּ�(X�����l�%������Ô�ה�n��	k�Ϻ�.��	,M�� G@C��0)�P�6��y��fj�ך0C����� ��] �T�T��o�W��ܫ�tK~�\�lSͷv�V���jZwEM��� ��&��(��=X}��<K�8K�0���UZ:v����+��ed��k�]8�7/�<���v�z����nc���%9S3��i����[W����7v-|��К�ss�stf)� ��ll�x��ˮ�6��9����+�Y�9M�ت&��2��#2c9���\���
�Srӭ!c��916M�	��AY���r�*�+�_A�����&nn.9���t��!�|�l
��o��=Y�V�[���vD�
����*�a�1奔lth��]�H��G}�c������ӑ9K��,��+%�g4��w:�hζ����uKr�!r�HN����Qw;��J�a��Y�$	�XSeb~^�����M��y�1o�Y�g(�l�ƛ��@Wq�6�9u��#]uv<|O9{b��z�-Ё�n�z_M�f`�I8�%����{�艣��|�Y��+�|�N���8��<<K���O��	�YJ���|0�.N�
<�����kx7s�G)`ـ���/�
qz� ��n��	��Ǖ�+w�Pg�F `��V�
���]�~Ja�9ښ��:,E�pB��Ix�U�;���^)�����f��\̽[�z08yѱ�Y�r��ʌ�rc͓l+2�
��w�U��u��"��l�.k�e�8������f�Oy��GD� _^�U�eZ4��{N0ܦj��rY�;�U�. ��9wxm��k�<��+�ʦ�b�c��s��P�l�cag�wv���=ʬK�2;o�S>�E�����R�[ߞ�A@�~��:��"û����p��֜
�����}7)�_E��ڊ�瀉�Y���Wo����� ��ܩ�U�V��u�{�L�y���&y��rş���m����4!9��b�JbXos�����l�1�9���>4�l�Us
���;2�c�rm������5��J~y� �w�9gx"�;�m[YC�񣋅�ݭ�Ϋ�,�!�.d�Íc3�ˡ�3K5��/p��)+d�p0o��g�LP�՝f�Z�D�1������LO-���M��K��ൠi���{o���W�.�t'Z97T�[����'4���
~�z=�8w�s��Fh�����4�DחR,dy��0�sta��=g�:{N�w�<5v!�<T'�{O�{��Lژ��;�+���;���Q^�>����s�E�+���� Y�Д5{mf�eU�幹v�[�� ����[�ح�CuAD�s�7uRߏw#:�Vr��������{;q-���&!���a�G�2�o�+���I��\A��VMO����-�e]7��;gW1h��Ἡ���p�\)����8_�Tĥn�8<+�kښ�����)tx��:u�kz�U1�ܡ��y�=}=>e-=
-�S����W
0�7��۩��6�5�g�TM�'���ud΅���C�����3��ބQ$t��9���)Yk����dۗ�K�AΪٮ�"ns���P�,���GD5�r��x�o�[V���'r�ovǀZ>E�g�X��Чͼ�Un+�+��(�X}d�u]��jZ<�N�^�5+e�,�T�i@���^{T�> �TNjedv]+�z2V��Zd���?K�����圫&�5Ͻ>�%�I{���"���y0]v?r�)�T���R3b���i&�m��Se+��^-�ԓ���U)�z�|�B�δʹy�u�jX��l�Y�u�*����v��wV�,jh���Ңp ���j�&)�����{��f<G�)��� |B�\�@�nƈ���:FG��1������*[� �²�;n�m�۲���e�'f��L�Ȁ�,Sb�9�o;�%Vp�2��9{���/z#��bI{�"��i�t�s�<Φu�3S��Lߚyji��̕��v	޳��ӱ����|���^�-���n|��{t�+��k�<o�k~u�u���)h��caiɜ�����O7�F\S.d����z�<A�B�;Y�ѩ�ȸч�'��S�%�ZP��rkg_AM~��k����FW�ⶩ��>N +]�M�AѮ�*@1Qצ��g�0��=���s���\��qR���.cg� (i�YeTZlOU\V*�2cDVeo��4���NYiw��/6��7Z���V���w:�l����j�`�Q7����tU�ӫ+���h^��U7R���K��m�X���1n�mO8Q�
bQ�FN`�.�Ȍ%�8���̀�E�Ȃ+c.�I�h��h��^V�щ�R��(^8���'d��s�iӝ.�'(�q��&m���Ff���-�{�!�zʡwL������N��hw+��5��L��͘Qp�z��G�G���;�H���p����C�o���j{JT�JùJ�6�k�zy�0rV󐲖7���ׇ�+�����X�3��O.��We+�����|�}��R����:�*	���x�~�{�6+�$�M�7��6  �{D�"R�Љ�Xl

�_��Y<2�[�.�!��'B^I�:s|��y�jO�R�(�e$d���N�5g�8���3��lޤ�Ac"�>z�8ҹ�*\c����*a�tu��瑋�'� !�"��"5�6�Z��ܼ۫WG�o���ei|X3Rm�I�t��t9�_ma�2Q��Ց�}K��AR���鴱s��;Z�ܽ��j�[F]e}0b(�;��UP��Rc��T$��D����6���R^j�;�ԉ����{3��}��c���`yKTרw�2�b��\�.�8I��a1�d3��nS�G��'n`4��g�kprxw�"��8m,�8C��W)h��c�̨roU=\%WW�q��؜�nzΞ7i�s�M�E߁�a�v`[�`s�t����0_���Z����7����M�,�b�ΝCg��q��5\ �+WhU����ʫ��N�	��'�a��3xJY��D�w�v3R�V�񃓷b�]��]r�<!�٦���4�u��{�z`�~�t�`]���q){!��A;��Qa�����j�t��Gf�\�CGL��V��P�S:����6$_-u� 2�<݁�/E�7�/ȏz"=�ݥ���T�ƭ���#X1�I�����
S��#��Ԫ}ǅe�^Oee�r4���y�����֩�+Ll���Dи�
��{�ν<�B�TߢZu�,x\��{��v^%ܻ�ɘq*�F�hi�C,R��F:lU�W���R��#�U�LlڍO�]���ؗtfH#gd �WL�.V*]��4��\0k�wJ��{�X/5z�7��s�mȡ�RO>{�C�7�`~Fҋ�L���ļNj>���@�唪_E.���܋�@umI.�nQ\�1���?��T�{څ��8�q�d���#5�!G�6���׻�h�I�ٞ΋�̗9&gZ�}	�%�{�W��2��ux���W+��ZrpU"s�Zkz���=aBw;�I��ZS�>��%��~3�y.O�~�Srr^����J���]/��[��<�!��u}��W�vW�Q�oq9�����w��\ǣ��i�=�ԙ�r;��Xs�9r�;���r�:���rr�A��Cr���5�^C�s�t�����.�p�	�:p_�w˳�z�����+��P&�s�f�'P����i�})콚��O�?���<����a��W���=��ԧI�����:>�9���|~�6�i��S6d@媾٨�K��P�+c�<�*�9��S����Ϭ�5�𷊂�
����=F;�Jj��1v��Wm�� ���ܳ21��br;&9ὴ{ ��j�-R0̾Y���t��}S9�Z�}��D�`*"�:����+�듯q�ߕ�{ޯSX��}������x_��=�{�u�+_��K䚍Hu��;��9}9�&�=�9�d�w/�X�N�y>ǉ�#�<�������9/W�{�67�&-�Q�p��~�>�ϽSS��@}.�{�ߕ�:���uw��ϴ�I�ԇ7��'S��sZC�Oc��O��r����\�#������9��8�7�Գ��gZ߼�Ͻ�1ya�|� ~��Cݸ}��ˮ�����	���I�{#��9�/�j5!��t{��>��֐�GW>��^��#./'�G;2�۷�l�.c�}�>�)ZNw�ײ����}���j���]�P�����{���>�=�e=�Ü��ө��Oҙ:������\ժ0R]g�������3�>����6}�9��;����|��4�w��dr�ǐ����jrn9/n�������4��Nw�S�7���o�?s����>��~��/��u/��k����vf��Oк����n���i~���`�@rN��ⴞ�}���ɸܿ������oO�������;]����G�}��s1
}�����;��r7���>���'W%}����u/q�N���Zۃ��	����!|=��������=J͹�?}����k���~�>���mɨ�^;�A�O �sJ})���Iܹ>��b�!���s�w-�֓�r��g?h:���=�X��w��2�5��k9߼���k�|o�{���~�����>��9�!��K��Oe>�A��}��;���Rw.O��w�--�w�u�w�1����1�^�����lr������>�=��@u'��RB}5�ۑ���gprS������/{���L�^��o
N��p;斖��.r�G�b!L$�>�1}�f�r-���CCo�]d����.u���"-:��P�yVUΠ�CWt��$�m�)�VK]G&��W'Nb�2�R�Թ�q��aN�G]M���|*��n	72`�ݵ�{�9F��֜�p��;AU��B.�H�&>�����T0#��{��~�i�b}�%?���;�q쟃��''��>��C���7>K�<��9'r�����]I�[�K����>�s�wڡD�U���ϫ{��g�KC��sz�4���h9�#�7�Od�y)���rn>�������Jy!ј��r|����x����޼ns���ϧ깿������ϼ������W��}.��~M}��%����4��0�}#�<z�I䛏%;:��;�s�;|ť=��y���u)׸��r}����ῷߟo�k����u����O��ވ���c�Gc1S�{�=|�K����/p�X�}�������5	�{�i������y�����|�ϒv��'�]�}�����_s�=�:������<�����w:���r�z7�}-.���Z���7Η<�k���|���?ޟЙ'#���5	�y�k'�����7=��4~�>�yg�ytVn�yw�u _��}>���O��>�{���y��CK�ԝ�9-Z�|�Z�{Η]�:���K䚍Hsx�2NF��kHy�k޾�^f���3��wߝ�}��O��;��r]��'�s�:��<������?�ǐ���_��@r]u�t-�o�'q��z��!�d�*b��s[�>��ٌ���}��}���7)�jz��	ܧ���k �'�ްy'r��~0�A���{+�?a�wy#�C�1w��ѳ�}ɏG�џk�_eu_ط�{������O��:�ޗ��H~��>����?�����_����_��}`�O%��?y�nZx��G!��K��_�٨���}��Oy�o��^���#�wTv,���1���l�˙�{&=Uyϼ��������w�>��N��惩�W_���}/�p����^G����>�C�ߵ��?:�3}��_�I^��D��g�����Bѿ�Od���/��-n�;jgm���n� 5��υ���(��V��KهrH`"kHնL�V�`͚�_v]��[꽋vL4xL6���,��`��U�v͒�8:}��&c�c�m����+j	��'z&��WZ�#��G���uȮv��>���_H{'Ѹw�^�7'q��)�y�<��O ���!�2\��{+�MǆsA��G����KݸN����ϼ��W1�TJD'W?�_�Y���<��;���==��G$u~�䛍˽`{)���4���t�a�w/�;��%��g�;��#f��ٌ�T�ґ�e|7:���BXx���&�R��x�Bd�q�z9#�^�rn܎���gpr_����'�����w#��4Ry.O��cDC�@�xK��qa^����@��n/{����u-7�'�$r����]��j��� ����:u�H�����y;��;<�=�s促���OT�-���s�>�8�33[_uM�3��Wk�z�IԹ{�ش4�F��]��toZ_B�{�˿1Oz�Mǰ~����[���������z2c����d�׳�>��Z�����a�����>J�Nk��?����Ζ�W ?w�-/9����h��������sZd�{��P�ɸ��<��� }g���XZ|;��y^����p����>���Srw.�֟�y/���C�r�~��-�zs�O�9�~k@�GG�i�}#�?=u��D8@��G���@� ����3��/����y�~mh����~�Ju�$�\�g���o��jW����rG,�/�y�Cn������vsZ�z��W��S��O����<��ϤuW_ו�O���iM������2G�טy/S�O 䜗-C�؆����P����:�r���އ�y�C��"�=}L)��r�3�Ǭr�����܇S�z��{)콚��~��O�_��$�O�xu=��>�C�ԧ��iyj��9.}��V��~��Ղ=�\���Bf���.s6L��P��[JȡB����ڷKTS3fk?��,Z�_O;7�PH�� wJr�zY���)��L����<ɖ����ָ�R�6���vbZx���zfN$���n
^�� V݅�v�G�K2�BS���B�D3jC?=��UU%��ݳ�#��!�������G��fbJ{>��d��?�by;��y>Ǉx�$�N�0�H�g!�w��]ڇr�C���7�����?q��b�y��{ޙ���k>����z���{�I�Ro�p�:����i }��ֲ|�����w'r��~|�w'$���ﾄr����j��s�γm�����������}��Ø�9����@�	����=���sz_'��'�h�S ���zO��GW������d;:��K�����4�k��2�ߍW�����~u����P����P��G��%󘽻懸NI�vs�t�r���'�짲x}�/����s�H�'���i:��z�ZO��~��Z���}{������]����u����Z_����4�;�߱Zc���G߳P�q�{�ZМ����9қ��s���`}�ß��O�j�f����O"��۳�R1�f���G��u�W��Ϝ�=s�EL{#p�^�;�����y�u!�:������7���'$ݹ�����wg��J}���O'�z�����f��9���O�s�����*}}�0�n��O3z�J��R��	��=@w.����PA�x}r���ܛ����w�ry;�|��Sprz���"Mvŷ���쯽�11\&}>�N��9�9&K�/��л���փ��/��{�I�;�����~�'���'�tk7H����rM��<�����G��uu'��:����
|f#&=�=�G$rN���K�~���z)<�'���ZZ]۾yօ�4������i=�~❝c���{'�М�=�j���N���{1��A�D|}1>�`{���� ���;�ԟk�������:ZG ?w�-.�ߎ��4�����ح��A윏e!���3�C2\نX7Cfe�+��I���l &���ܵp���}K-�� Ci�jX�	���n��@B��adH�U���|�k��3U=+K#0�d�W�]t/nVrRuD��ю�^������A���m�p�gmFY<9T�/IY���x���S���<!Ι�8�C��n��'�Gf1���'#�ب�?9�w`�K�w�t����Xբ�d]F��z��壂�6�XS,��u[�/9W�\/rs:[R�ٵm,r� »r��M		�u�ġ�Ϊ�\�i�u�V�K�Y~�3R8�Rzm��5k�O(�K�G�Ɨ۴�xS(�� ���,��u�_V�'T�MlMwQ�%��w闷��Z\`��2�T�/�Ќ;���ώ�-/���J�wص�t[��J�h�Lԕj�M{!�bJ�qm� �5T[��A��$�i�8�*a*�
��r�L4�D���S�<�ҭ�U&�Jհ&e���^�+�q��,��m�� 'c/2�A�V���fӂnn ^V� �ކƕ����/�Vfm�̾�q��?�����jSza�>�<#���kⳮ�.4��Nv���)X=KM4�T��t���qi�s������h��[�۴��Q��G��R�.ͷV;w��s;c�
1iWQe�"iŉ9Kx���i�k��L�A��&��*M�5Q%]-4�X��M�y�����j�݅��#�}B�;�U⇹�#�Ҷu��9�N��yVμgV������ک�$jT����Օm��:����*�6���y�;^��ڹ��[�W�˼��pՖM�8ATN񎤨7��0PЅ[4�:YAZ�F�ȷs����ل�@Q5�j����;x��ev":�GO�2S�5�9dՋFK�d�����!���L�v\�sgo"�>�N�%�F@�QODΡR�R�f��q\��o�i����������^���n�$)��:�'A9����nW �w	E&����?��|f��RG��P�����l��ȍӊ;��qJXU2���/�կ���z��)�`޶яEl�ňFʃ��{w�-l�AS�o����`7�/��W
��5m]Լ�J��Pk�ô�t�*��HOV�p%VI>yz��r�IC�t�&�lTvd��a X�r������G�>�$ Rr�U�QФ�
A�e�(h!�J���H��4.��*T�\���[�5�X���^��4FT���uQ�EZ�'v����E�sk+h�.5�D�l� ۖi��v=�����<n�-u��>ton��k2j�rR�KdC3iRqXU���Tsx�I˕����Ѝ��)K|� �)�v��˝w�y��I�T6ol�E���>,؜K�;�u�9�bZkz�NY���C0�8�t�V�����<�-ܚ�j�3�G��4��S+�:a�w̻���������"�L�
H���u����'$3+��̬r��"�(��0̜!�+,�j*ufYY����a�NT�YY�FfJVc��3V0U5VfSVf�A�e���dd�Ua�VV98NE%a�Kd��HSTQ�ְ��NE.��h���� �#0�
"	��1f")��
��0(�̣
��̥�30�PjVFD�Ef�5faffKF��F��"�"	�(�2 ���0��1p���j�`30��

�((���*(��ʖ��Ƃ$�3��)+3
*�&�l�j��h������j��� +2���"(j*�
��¨)�����r+!�2j���2�j� ��&�b��,`�3L�s�� ��(�g0�"3*�'3	�"��",̨�&�`���3�"`� # �ou��}����u�Y�Z}K��)���7��`����ET�<��6�΃8ɛ0��:F����:��l��3��e���/#?U��{��{��_}������5'��?@u	��?���S������/'�<�S�w/G����.�����rW�7�KK��?'9����vy�#@}�.>��5���ʴ�Ϲ.�g&#�1��Q
}c��;�
���'��iO �טy/ �C���r}����o�jW���t�G!{L�}--H~�;�}Y��]�#��s���f"��� =�3���O����d�y)��������ZGs��;���'rnNC��=�7-.���Z��=~�Ws�o��Gu_F���Z����C�����{�>��Ʒ��$�}=��	�'��Ǒ������9>��:��<���G'�^OǸ{/S�N��r��5'�u���|uf�J����~�ELzg�����O��C�~��V�7�/�j5!�7��$����hN�=�fd�~��X�N�y>�����c������]�_m�¯�,EEg�G�S�9s�����}�:����ˮ��?+@t��t:�����^��jC���	���y��r�F��>K�K�X;��r|��_yx},)����,��ޏ)�)��"ǌ��|���j_��ϸrZ.C�x�7.��|��p���t�ǲ:���/�j5!�=��N��?oZC�^�W}���tp��e}����#g�3똈����6�#�Oe����ey��5/��f�9/���7�/P������?sϺOc�Od�9��}:���zV���Ub����ϯ�9��O�b��UDt���~w�A俧����ZG���p�h;�w�9G��w���5�7��}hBrOn��t�p�߾�Ͽ}���E��]�gq+��{f!O�}�{'�N��p浹_d�;�i:��u~7�A����w�'r��}>Bj�xw���i:����_��7&�r�}Y��'o�'aJ_�#��)psj�k��Zh]�ج3;��l�)�����]Ux�,h�H8�f3謸����3'w]�6�K��xY.=#����]�JKJZ`�d��:�V�2�-NO���l!m5X��7��;a:�%�[7�"�UtPսz#��G�����B�_���t�'��[�Jo��r|��<���ɒ�toZ�W�7��'W%}����u/q�N���Zۃ��	�����=����8υҬ�=Y�Z\9��>�k��ɸ促}h=��w{�:S�O9�'�r}�Ӝ��!���s�w-��i=�+�s�K�0z�P�؈݊��X+&�nB���i�ߣѳ�;���z��I�nS���!��K��Oe>�A��}��;���h��\�������;�ߞu�w�^��>�	�ߢ�}8^M��k�/4w�z2��u9�O�pu!�'�p�r�G����Jw>`����=�;�ԟ�sޗ���9���r�����>�ϼ��u�\�Ob͝�i;�~9�_o�8��i7�+N��wy)��P�ɸ�O���9<�@�!�����^A���	�<���������O��\�>��}��-U4�_�y����\O�K��>ޖ�����޴���Z���O��I윏e;�
C�7I����wu�<��B��w.O�>�9�}1����Z��ηkw6/���}����5��{+��}.��~5�P.��o5�h����r>�ԟ����I��S��iN���O%�=��h��{��O���}Cs�]�������O�9������Ԯ���:�|�#����5�{��=@d���f��:��?֞_H�O��Og�y)���g�}����7��^��^�J�쵿C�\�Sϰ�N�:�rr\�����w�H��o�.y��7��<�!���	�r>���)�'��浓�w��.���xt��8>䖹��Yu]+_`��#���jJ�<�K����w/#Rto�9k��h��:]w��<�K䚍Hsx�2NU�ߒ���R����Cb�Gk*a�Z����c����b)��Uf�mƉ5�ҝs2�jҩ	WK���dFٮ��tш�}ZuQ�&��l)�v'},<Q�+r=�9u�}��&�C��7K����!���]���f�K��$ݝ��0���!0�?=U����1>���ϼ����=G��Z�<��_ư}���=߽�y&���:��;���yw�{�!��x���K�����{���l�ϣ�>��6�����8�����~o�|���Q����L�S�}�'r�G�Y��>�vu��;�'����h;�G���ϰԻ���{֒>���=�b"*b!ϣ�;��ϗo�C���_�7��y���p���=����sz_'�5!ϰ�'S�}�A��+��~�<����X<��r���)�h4w����1������{��E�5T0�N���7�?op���<9���NI�w���=�sϴ�|��������w�֏�}����h:��u�:�I����w�'�iyO�1M�A�{��^������ߧ_z{绸j�-�ܻ�����q�o�/�I�v{�t��<�}<��O`�X���r>޵�rn;�h:�^�t�;�A�{%�z3�	����e�=w��sϽ�y��4���x&�9A�?o��9&�r:�>�9&�r�w֢:}�S���1�~ߓ�y_�4�(��;�+��ټ��ϻ���k��S��_i oS0�'p�b��=O!X����ֽ�w�d�p��&4jۊ��	�����\f�1�*���5�[�qz�Y��;{��\Z�F"뢡��tj�nŗAv�N�9��Ü�U����X�^]�g��]�<��[�f,GT����4���W�b� 5�SAoHk*�*�K=|�z��މl�V��0���u������;O )h�[�l���S����s�o\��AZ/:eD8���;&�GZ�j}���l�8*������yF)�r�Åe���]S�RN�:WRq�G����e�j���i��WQ���ܫ�G͙n�G|2*�-�j�]��PbL�~��C7jw�.�'L������V�𔵃ŗG$E����g6�ipX��1Gc�љI�B��[�J�͊�u�����C5Z�d=�\[��ٕc�z|6`�$�s���;�.�M���i/��������5����`���5�����z�VQ[.������+ �*�3�bP��H����7�=�I��8���A�͗���ܘ���z�5���W?u,nP�n�<��f��E����E<�4*.R��	�S���P�j�8������oa;}p�ه����[���n[��]�&���1�3�������5ܥ*3��^��	+T^��x��3����֣e<��ge��ۋ�a�7�ό�ʢ��FW��Ѫsry���f�9yǵ��h_�W-��W��}�lN���2b�vR��<敋��L�S��>��A��ϵգ��&��"�s�I���5պ��]��q	(��tQF;�_��җ8��9uT�4]z��H6��r^VL��9��۴��_WL������N.�2?�4{�R� �[��}V���du_2}�-���vG|��t��Ư�]s� ����C�1g"�9���2�M
1(Ki����g{�E��[٨OO_�FK��(��ƍZ$���<L=�=��Y�S��O�'wڰŦ�O_��ſ%b9��C������[zM��i��o����4�:��K�U�e�D��MԶ3.�3C����Nb�����x46�c�9G����c��tħ\�f�|�� mj��U�%�b��ڜ�@�����Ն(�w��(���}G��GЫ|�n���9�����,BxK����c^�V�Ey�i�n{]wΤ5�T�Z΀r���k ��_X��N���E��1�3�,�P
�^s�Yv�w����"|�cz6/*�i1;�mc4������N2��j "-1F��Z&�r�x{��Tu�<�gּ�zf�"Y���o���ͼd��P_�z�5���n^/1g���;��mڧ�ޫ���G1���rtU8ȁ���8���l,R\�o��%ǻ��f����z:Wt=�J*л^=��r��b��]���G�r�+���rs�^���c���A
V��Ot[Xy���VH�$�����q���M9=Y�]B��m@���؄���뷝��;	���3�o-�a�R-Ouj8t}����k�x$�Q{�}��Que�f��.y�I�}���l-˗\
<U��;�<�QV��7Ӽ����I6w9��B���Ww�Okr��C�\K���Z��H��1����(Yn��n�D��ǼZH��W>8��[S;��1�V�C4�e���`����d�W=;�M"�C�_"b�Y~�L��v�b��q�ּ�C�v^����	s%*�O�Ò�On��d���jy~�Xb-4zy��qO[�F�t:j����{{������}�V�TZ�[>�ʝX���<:�.:ء�v֥+����s�ˉ��ً�-k͊�SM.�^U�j��T^<���{�0ǝʯZ5��Y�y����L��P%lE��.�� >ݝt��!䮱Nm������5>�s�ݧ.�.{�]lֻ��iX.�y��U
>{�ٗ��N�[�u��\֌eɊ����H�E~�
������6�p��fXv�y/��U{��(��n��oj��u��T4��U)9���YqFӼ�O�pZj��ni�v����I_ ��bzj�nt+`�uKS#q����:�\�cv�����[��[�v�jr+��&�9�0�1*���
�ΚL�̨��o$�mN��{n��ʴc]a�P�y8���=`��D �3���y8�e��U��
�`#7��e��#\b>A�V�=U���^M�\yb�O����5�ݡ�˨Q��|S�/j\|�>�*>*;l�w��-~\ϫ��b��;�X;U�L�*�<��|�a�n^��ܿd[n.��id�����y�-�G4+c�.]p4����p�|�\똜��7�-��ڊ�����5�^'�����6�0�\8�A�R'7Hv�u>�u��3:��TZHiU���>1����neB�X�T�v�+��Qb������.@��,�����6�,/�o�ú1�M�������m#W���]�G���IV�ף�
���V�̶�)�E��KrE����*�\Y���K��9b=�(v���Vf���Mw���U��� ��#���'r��]ϻj>�1��3X�*�*��L�HM�ɹ�S��q�o�y���e��]�f�{WL�dh�;:�h_;�=P���YFh���=�m�9u�˱�7a�׊2Y������>g(�9��^�)�
'�86k�9�̮X��Ή�Oa<�ϭ��EM�t����;@c�*��9�)v�r�>�wʹ��J��a�-�`�������0��i�1�7�.�N��Ǥ��{w��r���m)_H�ފ���(}\�)��̨��_c���8CtPY����{�h��oȧ}��$���Z{9N��{��z��i��$V���5颬����:���q2K�!�]X��˰���s.�[܀��~��Ok��и��>YK7��"���`��yr�~r��LЖ-P_hse���I��+hEyQ�������V
�t�S���H�f<�WX��y��:]f?-.�Ǌj���F\��N#�78AØ�R�p�&j����n�yrK�7/{��T�Id�m���4�C��͹`��Lɯ� ��{��l��ŏ.<�l0�ǈ��T��߫��������Յ����!�z�+��+v}���cһA�p�9��u���*q'����.���c��;���5���js�}#B�H��8���ֳ��4p����1�E�z��V��M��=��׻i��³����y�����B��U�q�w�2�`�I
��6�y���wƒY��M�ܤ���C�\N��f�_��+�#�"��i ��y��A�ͽ��7֒S����_�w~�Ԙ|�S��p�[�����쩩����h�aX��f�b��'��أ%��^Hå�����E�v��[Qܦj�V��#S;��������ſ$b�:��CEf�W��Muх=��QkM�A�D����beߥ\JŌk>�e4{z��w������;Pr����V�_m�*�Ǧ^N�D�Qȇ�$�_
�v�L��p��]Gl�Jo�P���%	�zl�1�i�B��N�nr̩l��j1c\���������C��y�]8�A+�^�� ��j����d�"_olp�w�8�ok���������N��~�j3^��9�0tWV�)��}_W��՛�K�ſyÒR1��T�l1a�05a�N���]ЫN_���E޻�)fַ�P�m1�C!+bxK���}�^�Qŗ�\l�!^w��*yMSr	��y(�BV�q�� ї� V�bv�x)֜y�&�v�F�U����Xu��LW/VW����6'�=��r_�)���m��ؗ`��qN�%^����#\cR�y[���� N��F����ݵ˭H��c�V�s}�-�������C���_�]��؏SǤ�9���M��|��Yc��eh0��1@��Q�Q��垡RE�ܑ�ٻ�T~X��Gǔ��sB�0�.]p0�qW�2�E���#w/J;��A���:-�Ŵ��<�Lא�P���5j��(�ˁ��ڝ�y�@�6�uZ�Oyz�1m"�yZ�c��-����hբ#eKq���Yx�Rm&}��p�B��.W7}���6�Ӛ����䉉�.J�f�R2������J���<s�B =y��i5�����SFAz ٻy�2݋�3�����1F�0�9n�OD@7H�����oTٷ�Rێ���b���Yi���'WPЌ@4�C�+))�eA���Ā8!h��c�pWz!Ŷ
C:vnjS�]E��6%�V܃�T���K��}�ans���X��D�ٍƙ�`��t�ۙ�y�O�}�����Ȥ��~/X�s����F��n3�gRR�n�=��!4�A�F��
i�zWV���fm��c�׵E� !���k�g:bnn���s��I���bG5* G���9�@[���e�v4�ip3o�hX!����%޻;��ͳ���wIӉh�Z=u���:y[B�K)�9� �h'/cr\�ú/��U�I��3RN&���? #�ެ�;.p[<4E���£\���Ƙ�ޭ�y77"��n��[��M���h�O�*�+����;��Z�o�X�U��	c��G�u�4[|���E��@m�c&[\
��ow�l��w�Â6��Mv�\��cW��<uh�q��IW��nѕ��K��v�6 #��2���I�	�t�P��O�ʋl��Mv6��{K��j�c�%�pM3�W)���,��R�=e���*+�x�SI�\���0��{����3�АN�Y�
�1[Z]nL��wRȺ]CB��9�H�N�r���+���uk���n�k�a0�b��Zv�0K��K���nVC�Cw+Іe���*J�ed��5`�\[�ڪ��ڗJ����j#�G4����;��ד?G�;�0A����[Oi֪^���{_;�vvKβd���@u�� ʁwu��WZ��M��v�=���2��N�ab�St�h���ь�ޝ���W2���;jc��עdf\���n�i&,V���V��Ғ�P^&_u,�[�u`�,^��x_t��Y�"�^�b#��-.�ugov�i�P����A�	��m�Ք;oH�|DW��k��f�ǳ�w$��Q��z�C�$.�\��o(��6�ʏ6>�y�������R�;��L�(�E2�C�^(�R�l�Ù�n\kZy?,{�Y��Pf�41�=tr5�#�T��%�y�_[�YL8m�X�{�soUиU�Ʈe4�(���b\5o�B�g[F"�C�k�&e�'�iX��
��~�wk�y}]���+��2f
|��C�;N��)b�))�j�f������ᇃU���B���\T��c���I̗.���7�6���i�h`�h40n�B�͡о9���HY����꾀�p� ���Un��xͼ;�:�;�_�Z��唳�Xd�ȮZ���Xr�j�R��ЫHs�9�lɛ��^�qk�Ė�wt��q7�p��+5��>��$(� T̹�4EQQU��TNA�f3E��RU%�eēDEEE431IQ-L��A4�QE$M%TUE9�MD�faMUMTE5MTT�ITQLE4�Y�DE�Tf`A��Fa�TU%�S4YAYd51��d�EYe��USQ%UL�!M5D�$cU)DE4��AADTQIA�DL�c�Dd�9�EDQMS՘8H�LTD��B�L�9�,�URUUSDTY��QKVa�UMfeMU3U	D4�P�EPAMA	MD��a5EYa,Q�0C�TTE3E$UQ�dHP�K4P�DLSIDTDP3ASAE4PQACUfK�Va�RPETf�4���MAIIT�TCQQTXVfTLUMUPD�PDET��aSMD��]���wW����:���m메��i��k��4�s�3ʙ�R�L���j�c�
|�h۝ڶY���F̃���q!]o��st�������W��[�|�vo��/���Ցm,��L���;�����������W"S:r���䡫n(ZvOP\Lf�����C��H¤����Q��y���{܌E��)��,�B�0}ꒃ�`�\�e����>*��ۗږ��b=~�Wϛ�f�uAC�A[�q��=�vck�	�iEިlʛq:��nX.�U)[�_�V,�6�K��$�T��ou�癰���^N��a�7X��+`�ꖯ�V�������T��V�km���/rVcLd�=��E��lN�X}�t��1i�����N��fp��}~6��2�u�T1P�H�➱b�n�ʅ�Bȗu�'g��K���.R�4�	�!��N�.���5�#1B�"˂!�ف�i᷸��nl8�Y�u��,9��ׅ��Vx�]K�����+2�+׵��]*0�f٭�T{� ���.��b�	�k�k,q�O�ѯDi^S�= ��`b���3��ͼ�`y���:쇚�P�n�o�̝G�,Uo��gx̥��V--����)c��綞�Z�'\�7��\�*b齢� ��T�a�kOq�=��R�����޼KO��ұYX�E�7�t���u3�o��{m���|U�onmS�A	z�A��o�;/9n����ܸ�\R�ԝFL:r���w��]�^�_���F!Qy���=�eL�҃�,��uU��Fu+��ٺ�*�lջ���W�+֒9����A�>YIlҁk�9tsK׻��L�Y׶�b����{-2b�@��i�}Ɛ��z��,�ؼ���;+��(�g֔�0�EF�Rb4jۊ����\Lck`���3�V]%c{9�V�ba>���,��F.�����[~����]����3 V�'����q/]�WPQ�G2�<�����D-�ƽ�U�	�b�èo?E=t�.��,�~^��*��:�Ħ�Zq�8��oCX�������Z��e�E�b.1Vc�y;	���|�;�Q��p�`�����<�f�j}��!n�D�m�C�+�;�b;c:��^wK{ڽKAw�wup�-�t:({�*��z����\�fo�T |���ܬ�8������`U#i����C��owok+�N��ԃ�fdPw꯾����[��t�>��xb(�ˌr�љC���ݬ?J����Hv���z^kz�3��b2��Eia��ע��]Z<�V�`�͚�f�y����rݨ��g��kk�+�o��{�p���f
]�]��GKӍ�գ�<�l ��O��&�yX�i13�l7����6��7���:V��.;e��f�6z�i�R��vy=�~k4}�.hv`��b��xR�FQt�Q�ֳ��U������^Q��s��Ԏծ6�{�l/3Ĥy��malR��뫇�ؠE�z�8$���	�����Y}��Rm�[�w˳3��9��Cr��k1�a�_(���<�k:n�Dಪ��-G5�7mƄ�O)(v�i�s��٫@����d�"%�����ؚ©���'p�g_�;_I	�9�Ý�O���[�h� Udm��#���XG4�hZ�Y*R���f�Y�rGw�5Z� ���zJ�� ��Lg����p�Xȅ���L�N3*ɮ]���r:��!8䩤�7t��������SL�@#XT9�p�.�;�Z�m����}�DDF��N��͜Ҧ�}���f�m��zz�1FK1k�:QZF^WFVF��1���� �]�:����3������������[�F'gaR�{��fm�K/�{��[:�AY�qyS�C;��0/�p�Y���5�:�VhIg.5���������u�n��h�.�P2�Q�&�xގ�]S��z�^�#�hSjb����~��|����?*��8��VlWC+��hy	NO44O�yu	�Bu�KY��S��)��������mU�|2H��V�Q�3ݝn�?��}�ȾȬP�i1;����bv��V"&-A�x4�0�W={��ق��x�8����`����$ݿ+~&/6�.Z��p��{eU/v{+Q��\c0��ن���u� H|�Rtz��,M��E�畭��>/Q���ӧ� Lɽ� ���u��_�4{�61�gK���@����V�D�PPs4:�D�.�
v��'��kUqk\�7��hP0V
����>����Z�c�N�ʹ0L���S��D(�����_y72�*�{%���z��1��2M��9��ΧMG����IP�=���]��y���o��e��1�ۊ�|q@�Z٨׫�����QT�^l�%¢��va�-�G4+�r��@�v�>gpȩ�y5�+��Nv���#��hM#
�}/����"��C�\�{p�Z�����Y�ݗ����
�Xuȟ[H[K�V��6���q9�p�69!�yf���sRC��>��ɋ���>���CO�\� ��#F�n�jrq��"�RcF�����Һ�S����hR/��^Q���x�|_�z��sh��7Q�>�5h��}M���X��]-l��t��]�}��xpK�{�%����5�K�Ty3��vׅ��k]���nH9�f��k8�t���o�:�r�>
�'1�C�}U�$ļ�]^Μi�wn=��zX�����K9_�K;��.�T�;�$�=�F�����*���{��n�G=m
�C�����)WT�^
>H6n��J�Z9x;��1f���%q��md	v�F��[{��[��	1�v���/�w-ďn����e;����0rs*Yn���fIZ�U�dj�jǴ���]Z�Y&�u_~{�ܳ�z嶗��ۂ��c�FcYЫ��X���	��a��Cz�M_b�Y��h�"��	�>�ٵ�
�/0Ӊ���x���
Lk<�V��4?%�R딦sw�O\��z�FQF#C�qk�_B�g hv�U�]8�`q�⽼���OvG1�a����;�1���nH��͝�z���j�j�s�R��f�v���}�,�!�G����bF�[�Oaǡ�,����5۬�X�����v^r��sB�1ۗ.�w���tB��̽8�ZO8��P/�Tj�$�*/.5��<�eL�WyS�f+N嗋��v�q�m��%�_(����B��~A����h--Ì�k���j��!��[~f�\UZU<S�����xi�ӵ[I�kz�l�B�z��[�7����K���J�0�0�^���D����4�Vm�{�yy╽����ݿ�#��S:���Z�,oc��	�s��꽤���,��$����S�{+%��Q�A2�$�Z���&Y��]�7�EA8�m�7 ����r<�͸�]o;�Q6w��g�N�f[P �.��<���_c�gM�[�\���a���'ԭ��+��l6F�0����:3�ꊶ�:\��U.P��fqO�^�L�;����v�@f-��b��t��mӌ��IMh�ND�E�I�Ǖ�Տ�]�z[��q(�e��n��	�8��q�J���^F�����b^��w����z�l�.;9��+0Z\�a��6�:���a�>��ŗ�r�����c'V�5.�9����8Nc�)\�s�!b�8`�	��j�c��&�����)��N��*���g&�����਑�Ey����@f�bz��~k�弌Y|2��KD��k>P�d�Pw8�ށ���{鶔�+a��F�<�N��ֳ'{s�/Uek<�x�B�[���k4}�.`l[��&�4���5ph~G
��1�[�}�Q�౦^��e�n��soF��;�%t�:jI}qؓ5ԭڎ�hB[��B�ά�0��=|ʲ}V���>��r`u�mû3��Y0�j��ʝ���g�%t��о�oD7��R��0���v�<�M&x��r&��E#�xl�XNY7&m0�/3:Xm(���U��T{g�}�6N%��7���,[��+��<z�W��@��z�Wr����q��H<f�,�y���]���q-�#�Q�@�v�)�(ȴ���{x-n�B�ÜV��`?z�p��yI;s4�Z�5��qUiYz�ճ�r���-y�5����u�c���O��;:�\d�ne�н�Vm��b�9�Xt����[�M"��P9��,�f�b-�ד�׊2Y�^H�(�3O��S�5vo���ч�ۊ��K��#S;ڰ�hK����k^�����%��/������[��œ=����忎uͳ<��0S>@_�s�x���D��ѫ�#-��l�Z�A|b����K�פﮗj�Z�+{a�'lG�h{���#�R�`���V�{!3|������+k9+H?F7(��v���<�0G37�<��9.���1S�^��R���v�����M�n�<�岆&z�)4ob���#�Z�����z}�*�X��4�f�t�+ٛ
�<��z��mjD������d[�C�Qk6/2�>w2��9���_W-B�!n�j.��5��
jyg.�)%�������#�#���,����ksں��?�8�+� ���nr>�X�:�s�f���Þͤ�o�V��vt�����-�|�ֲ��1���*1��y����3.Ws��<Z�>��X�e�����6�1:�ej<k�{!^V�(SxO�����If���އ�C�����z[�r���L�՝Z��.�w����:ߥ�[�{��yD�����K�&>լ��ڥ�(�y��Jc�|�i?GN������B9�\Cr���7�a����f��x���e}�+�����iE���i�nyڙ�!֡��z'�-�N���&�i������q��U�'֒�m#
����1�Ο6�k��+¬�r�}�P�Ƿ�ۡi\���[K/53����ʒ�bVM��,�<V����3Y����FΩ��ⅧpOT��jyq�LLӳ�#=�%�x}ZÇ|�$�b�K+��u5��`��^����4�MY��{|l���#��M�n�h���d��pM��;i�2�ԧ,o
]X"�:3[k1*(8Y<31�s��e�]����1��:wBF�T]�wv����h,B�f�\��U}y�C6�G�z��Tk3�_��$}u^a�l�ͨ��M���ef�^�v�N�m�y��\�8K*<˿J��ߛ�PB�]kۨ���n���5S;�j�=$˽�e�w���1�R�`=���x��SS��p5��+5�ۺ�X�ݔ��wAc5���Y�<�2�c�
�#�Z�{8�o�YjU��.N/(s���n��^|��c��4&�9�RGeT��Y�ʪ�-��;�����a���+Lp����6��Z�/5C�Nu��*h�zKm�\��In����hX+�
��Z�4��B3gS����g�����ⅎ;�v�	���n���=����{鶓f�"����x9s�1z`���N��:J�7�AŔ�m=Atݽ������X�E�y��H*wם��)��Cy��vL��?T��5�Y��s������[��s�uUm|�N$�nQ���|{U�xo^��k�`��\{X�u�/�����7������� kvFhđ�:|\�"Dъ�[S\�N"�=�2�0��޹�$���agGl�q��{H+
����`��%%��x�G�.����E ��Z��k껀e�mJ�K�ˊ��-�F3+w�pJ�5}a˹��P��q��TV��-�iw]EС� P����,(*�6Rػ�Ң-(	=�F�uB�/]�ޫ�V�#5���bL��ʒ��x+;�]oC��v�q&��G3.r.�2��C]ܲU�r���N�1��eJ�w����)+�C�|i�@zo�uә�WL͵x%�+k�tN�:�-��#5�-[SOSZ��#[�f��cpN��찕��dPd"��ӻ)
�h�AwZ�lW.Wm`���2ƩVD�U�z�k��ku�a��o[�Ԧs�nʏ����,˘��So+)KX��F�1�|j�0$2�$0ͳY���Ւ�����
�;�f,�we�l��4�iq��d�U�V�¶�h�u�0�)n*$�l���s1h�5��9SW�61t��÷���/&��-	u�P+��ۑM��ɗ6x�����q;5�<��'J�Aݕ�_pZo8�{�6��\[�������r5�19f�oW1H�*�4��٧��{Y����T\����맆�c����Jc�BY����#��[��s<Zr�yfĖ(Q�nrI�Yua��/]��qITI�t�5,�Z7Oi� 9ܺVk����r�����b�&_>�Sɳ�V:�f��G'v�r�d�Q.r�ܬO	Y0ihM�^��u��'Cw�����K�7��_�z��}�,x-jn��#�R4v�޴Ř'���,��i�����49:r7��eN@��[5����B�T��̀�n��R�)��]�(n����t��L'kDe����G9
�]�j�9��Z�@Q�2�V.�bu��uZ����sA�0�sBM/C�Y�Y��\C����kv�9􂊶�C�N%f(�����(��nu�FZ��u��SS��U�s:n�ybQ";v�<9\s4�e�F���2�gontɠS\��7�����P���X�;m�u j�'�J�Zx�铠�uҺ݉�4ͳu�q�f�l�U]�ݝ�mX��ns�G0@UFr+]X�5kv2t�K�N���u{��ih�U�^�� T��%E�	u2�+�6��V(S�]sW�&�]���|:�Ő���d.�T��'�g��{7^���wZ�*,�-,��#MH�n9cfJ��wG\�SEi�ô7j��ëh6�*���46о]�W_KD�u�:���W���9�>3��tee��ϸn�K"��*�r�#�ZU	��)�[ң�:<��ӷU:%�n�S�9�n4MZ�ݭ;��-��y�'La�ra�9�;mUUTST2TQMTQMSMD�QDEQE_YI�A��IDYT�4�UXa�L9�IAQTPEdd4EU4�MT�D�I1US3Y�E1TTPDSAUT�Y!�dURTADQ�dRSATM��Lf`�UԴ��UET��LUK1$SUE5T�L�9QEU4�P�5�S4R�TAUIQUUTIDMAPRL�P�4�MEVFVNSEMQEU��M-EM4QU�	@U5e�KD�U�a��NS@QCY���QEPD�P�-RL�f&3SQL�IQ10�fUQUc�S4��5DNY��fd�1P��TY�Q�EELUPR�fd��QA0L�SIE$�%DٙY�QffXE1-$@DEDET9`W��w@��N>�/Nl��K�k��I���K�S�4�KPeї��*\lrw��jj���V3����ܱm.��%�[�.�W����ks�A���~���1@����Ir��[I�{�'.�+�мu��o(���l]��ś��j����y|��-$sH­�5>+}W�`Ţ�{;�q���m6\ʝ�Q�V�3X�*�+�:��&�CO
���n��u)g^��w�n6�������iL�f�Rtjۡ|���,�`�p�d,��s�žyq���|'�\c��}o����4V,�����yx�o�!�OV�Ն"u;�iV	�M���7�b;�ݭMlp���g*}li��0��[~�����1�j���w^�y�V�Ү%5��E�C��gZ�[��O��wU�.*-;�[��*5��&��N����m�(�ʭ�moY��h�j�<l=G'��{��]���(I���mf�u�$���6����9,`�q��Vx{o(籧���{tP�*�o3��7a�7c�q�[��NL�,������} ���-�p�Ãz�,�u�du�.ftU5��v'ŕ�b�n����\��[����Z��hs����zv(��u��*r�ª\8�����oUEK�IA��r�Z�Y���R�"<Z�*+��9��
J'�B�t>�*�}pk��6��o�,�Y���h�]�Ѽ��p�G'���C������j"b��}�R��Mn	�/��p�ꌭ}*�i� ��y<����u%	}Y~���3'C�3����լz�1@���WJ�ӷ���}���p�>ms�]vy%���r:�moE\>1��F�}�%[���W t� �ޢ{�v���~�L��{��hW��ٰ�.5��՞ό�h��R�+}�w=����Ю]/Z�ȩ��=;3V��ҬP�q��������7��/��E>N����<|ۙeR�ѫ-��^J�3�ӫ������d�@\N4��S6�j�آ��Z�F:�s��fb��4C����n����.���b��O����u�.��V(@�pv����d��?s�Rћ������)���H���v�h��»����WP�6(݄�׈��k���eC-�(�P�.f��J8��6C��u��wq'��Y�u|NZb�[���\&J�ɰ��`(����%oc��]P7�r�3����A�h׷Qkn�q�����B��ɲP�&n)�Y�z��Ү%�̷~�ep�:ע틌U��2�Q��qv�3�_�UG"�7X�cGT�p��a�#V��������_:�V���8�B����Gk�t2Ӯ*Z���P�nd�Y��i������f���ۢ�\gk>ݡ^�W��v�y\�m{��C[�˭7I'�i�w�[3e�g_n[�����T*c���>bû��*�f9�Z����%�@ۢ�r��F�ԣ뾌[��=c �C�&b�2��2�Q�k��,���s��^�7bmpC=��eR�϶�}ty>+�r�H�{��o;�iip�>���<��o4t>�b�U��/{*T*�&*oY65w ��o��Ч�7o9ft#����r끄x��r�|�VLm�1't;9_T�kTj�~�<Ϲ���:��Ǒ�-��s-��ݺg�g[Si^:ۋ��-솲�(N^�s=0����m�R�43����g=���>������� C0��*�0����l���Ԇ6����F�q�os�7wi��1}�q��[Ѻ�Ђ~��Q{�V���*�}/�Okr���C�eC�&��ѽ��ַ{���k��Y=�|ɴ�1�i[���\�n'WS����8�D�ܹ���|�"#���i4������磺�aW����>��;_���my&f�RcF�����=+��}�X=��R	���0��{��d�����uC��4jۈ����[c_��a�0�]��o�:{\���}�|�(	�q*�Q��ٱD-k��u��KjB����^E�:�#�w�J���է[Ż���ʸ`�R��
��'����X��9�.���%�Fڸ�՘�k��*;Xm�s<X�6f��ԕ�j�b����l�@w\�U�Ӿ��Ρ��΅8�ݨN���@&�6�"��Ԗ�m�f	�Ҭ5����q�����e>���wV���
��`:b��ա���<�.E,7\��9��B��ݻO"b!u�SKv�E�[����n۬u���@yI��N�w�נ/F�h4����ԊZ�	^�^�Ҳ��	�+���(�5�=6�iE�b5�u�]ݠ`άf���H��=6-.͹��+tĸ�QQ�����FZ�3K�B6��ϳp������$��յa�{	�;������e�*�i݌}�W�썡�Dn��x�X�v�q�	������а�<jVl,vac���A�>�bWp}s|D�R���O�K�eK%���F�F#��q���>v^r��sB�C���-ظ��}���9�.] b)qWF�/�Tj�$��y��)�V���=;.��'|�39?2�\�Y��V��p����^��o&���=Tq�K�.0&}����nf�PcF��C5���Qi�u\*�u��U�p�m��N��!��z�'����R�9��a�Ȍ�P���]�sS�]_!�/Jb�<���}i�O�v8�f-�#u�L>��R�BeL��7םMm�c�E�}eK�ȝN���:e�y��n#n�� ��g?
����UL�n��f��X�Y�+[]�nr�n�m�ƶ�{R��T�Ȃ��\�4,�9V�v��L�\���A�o��3�J`��t�p�X5R�;4��Nz�9����t
�}����Ԏ䕭�CC���Y�|�-$\�W�*�%���|�[9�6��հ�Q�˷�g�i��s�=���`��7���3U��e���7�1�y;	���us��r�j}׹=�,s��Λ
�0:�'5���sW#K�ؖ��%v(�n��3�<t��f���BzJ[Fo�O��k�袮z�쪻=�Ҋҭ)�~�C�1��ڢ�k��j���	���xԆ_X�7!��'gCl�Ƿ75L,�����Vyā��̓�E8�-��&ffܺǤ��>{�t.J��x,>�x�*�>��D�ܹ��UV�i/E'7�{��,����j�k<�o�E�y�Q��v�sf��b���t��{W��6�{��k�s�}#G�&vL��0��|�^�3᪪�Y!=�μm_*/΋ێmx��C9�\ �/�Wj�h��弡�a���ݛ ��PU��d��-d{����:n��K����] r.ƥfs5y2���F��LN׳s���J*��mX{N����v��q+���Bb�MO���.�ص"yʼيf�\�����5���,,�1/�Ňk7{�A�e�@z��c�Gʏ+��6���;s4�Z�N�ۆj�sNGT����n�]ڄ�Y��m!m��|������S)�^t��Y*%�������e�I`�p�=R�'�.'Yq����OOZ��\�45��U��V�;��dT!�Q�;�{�]��QڰŦ���.��M���D<F�B�g���!6�}�EE^�������}e�O*uc�wr&̌�^qūE�s��k	]KbUģ�w1�-ֽ�T^��p�::�r��γ|q%���[�bR�O!��r�!T�lq��,7��dr�n����:�I�n2&	��gǂ�J�؝Qg�Y��S�~�"�ä]۽�K�ߢs�4o�Ϸ��+[�j^Z�A�Y>�F��f��RJ9��Ws�3�������*�裑���t+z��r��W�L2!�&Xi��Z�X��j�/�c���uU��-9��u�r�xk%�ޢ�eE����4=ܢ�k�Uw+j���,��jOqT���y�$�@'U��(�Ӯ�i=�]ջg��Q�ax�:\��QQ
�b
��GH��۵;�u1:�=��yZD��`	\�C4�����+�7���Zܵ�s|�Ci�/''*i1;��K^g���|k\�]��k��E�>`��b�|Դ���L��f�n�B%0U�����e)~ڮ�c!2\�|b��<�1��6����"��8F���E^��,��
���,�D�h@�BӬt���2�m7y/D,=�xv�*��h�_�`���6=���yt�S��]!���T�J�]�T��r�Xo�NzLy�\�hd  6%��t�C�J�)V+���˻T]�	��d�C �L�zjb�sm"���Tb��X��Rh�#.�Ú���.��ӻwHgmbJ\�M[ҷ̫I(;�44:�T���=5i��sub����I�Q˟-3S�S�}��`o�w��;�GC��1�x/Tz���	k:i��t��Sƌ;�����#�ؽrR4�Z�
Ҟ�����s��'db��&quZ�*�	Bv_8U���,�۔��0)��=��5:l�>]���D{l�)S5�}�my��&%[K##T�ç/�W�e�+����O��s(�o��:V��J76�t5t]��XNF:��8���{��.I^H�5 ���q��j��{�pYK]M�Z�j�C��H��[�`=�o�fq�uP�yp�T �{���u�NZ��ʴ�}�n��Y��*�f�xKq��/�,R44�q8�>���soov�������Q�<����d�VVD�}��Z��r*D�3J����k1iB��e����E�:��8Ж�6z�.��C1�T1S�S�i>t�;�n'��wyi�%o�>z��\�����o�b�N���X.j�#��׶������!����neq%>��55��5y�s�ʜ�87�j�ԓ��&��CiE����Y.�ӳ�@7j��49�_(I��]6���錥��������b�Y�K��$y-�x�h꥟
3L;�OD\�šH��� �tT�u��x^�7Y��{C�<�kj4�㫶ַ�Z�+K-i0[X�3�Ժ�я�^�T�ϖ��U3<��#�>Ns{dS��:ˮKM-��H"hl��+[�Zk<]i�=9�=����@$�j�oy�gw�n5³3
v`��w���L�ϭ���9|��yP�1״�ԫ9wi<�����(#�(�M}ͮ��a��:��5m{wײ;�#)���D�-�
{����@4%�ΐ��XT�p�H3�Is��e��S�ӝ��E&��N �Y(���Yr����כ�ǥ5� A[�:4@9�G8or��a�x�ʐp����:,��O��B6��!�A����Q�o�9�.+�gZ=�.1֡W���`��K�a���:┩ #�S&4P�@b��-x{Ɨ�&�&����td�~��.��7�J`�}qW�O��ȍ�tzOw�:H�����γ]���\�n����~��6�����g�zx]����\���UD:Xn":���t�ޅZ��~��ݞ� �92l�1c�K���r�{ӛ����$9ژS��e׺i�ҽ�kn��M����VyJ�\D����\Lٙ�Dd��u�7-�kL�S�zS:N�|�>�k����ʣ|�+�Ĩ�ڝ�S�ˤՎ/�WL`g�\����m��f�Cs�(�a�*t�׻P.a�,��m���S|5-�ŷ���G�7 ��˽�k������kh��@cT��s'�7�tF,���Fm�����y������e�f��=\7-��U�C��}�>j�*��].o��=�$W�;�m!艴����/�Pj��{v䛕��rr���}��
�@����M9C���%���]�]ڵ9W�U�hI���$'U�`�)�\u�,Ȏ��.�Dt����4nQ�=VG:�U�hy��Բ�E�U�I[�L�Y���1�X|Qc��̶mP�
Ί��(_`�:$���!U��,>����3`�9��M_�
�B��qq�G��r��|�V��ݜ��yz)�s�y�cEsg9{C��l7WZ���j�ӽ6�	ǹ2�ɷ�%�	ojP���YΦ/���:@^I�&C�i�;�؅'��_��Uį��on=���r�Pw���r���%��)��XZ��8os���R�,�ٜl�dP-:{ke�uV=v�XSV}{b�u��J�����(b�"�^�dĴȳ3#�riՅ*�k8�b�v�=��I���u�m.�2���F��֣�d�\�1$
ܕ��%jC��9��̍\���"��D�k^��`�߆mןS�i�M��V�i8H4S2�N���#A�qQ�VÐ��@R�4�%����4�u�,���!\�,+�w�K��֎Z\�N6�U���ɚ\��m�f����s9��w�^*gR�M,���(KX����iPw��:���U$��#�cΏ�Ͱ��R�3��W�5!��CNn�4�Xҝ��U��ݦo%��3v&t�u���0똪nKB�]���$�Ɗ��͊���YC�&.م�uģ.��`��z����Hk��L�L�,�H��\eC �SЭ���G����չ�W�j�\����IK����eT��]��ƽ��,���)��>CN�͵Vc6�n��j�����"-���v�8�\49Q�z�ʢ�<#��AkwU��)顦��;aL��?-��m�T>���b�ŹmTLwA�'%��4��d��YjR:�#oy-�bR�]{}�әk\�^n0��,M4�O�]<Nn�YaBeL5u1ivE(]cr+�\���+�Y@�x���JO�)���������|�-�c(v�@A�R`��kz2��������,ݶ���G�-��z-�u�e�-yQ�v��Y��}��t�
V��-��i^���9����Z�*�eё �.�8nRUΛ!��Ŭ\��w�>F.�r���b����LNecӸ��˵�a�t�I)����h��]8�6��b�X��]��`�qu����V4�����[el���8�J�[F�gt�ҥ;/�ػ/_�[�⽣���+Ӭ7D`�,�>�j+v���������	[G4�n[x1*z7��`���ݘ�b,��|Q��
�a�Ӽ�0�Mw����p�T�x�:�����иz�NR��Ʉ*��*r���@�ʪ�8MBź)G�����Б-�K�V����(S�l&-��8�a$�)�i�Ѷ�l`��-+9��t��B���TDLP�UQPRRS�STEL�T�dSS5D�EIKaCY�L�3IDM6fT�D�U50@QQQQEU5U1����L�Vf4TUSQ!3MR����f�DQ%Q-�-RTQ&a�AQM%QC3MEAI3D�DCQUVN0DPMfaAL�MA4D�SEE�S5�EMQUQY��QMDCDT�T�4�@�T�QYRL�TA4UL�5P�Uf9M��DDP�TTEDUFT�0IPTIIHU3��6c�TLUEE4�D4�QT1LS5QD�TDMSAE%I4VI�RDUR�FTMDUT�UaeTLP̐EAQ4SLAEMQQDTU��3]��wMe���+Dh�����#:�H������Xdg��9��d�ɼ��]�9��;yW�\��Rl�A|f�fN�_�%���ò?~��(eV�>سX���x:��KDR����v�ݏY<b���n�c���.L6ϰ�V��E�o����oc��wtM*ʪ�X/Ң厚��U���GC�����j�W��I��C��=���P__ 5(�j����.��o�R���˝M�w����)���_�'�Ѩ�<b{��J�8��� �K!��{JC�S���g��=7��v\�9+$T����m��Pzw6��5{Z��z�~R�GX��{�}���9P6��P����{� 3�)�E�Gn��ǵH�Yw9<��Mv&��x�g��;�2�=N�l�'�:c'�6v�b�k��<��*S9�vD�������n� ˓��Prw�P�����/4�-:;��:rj_��#f��T����(��.�����f�����#L�%��nins��̃xܼ���B؅75
{|ϟOz�/GW�P2;H��.��b@	�1����x�����G��<��R�j�aW2�<}�N��|x�Y��(|�pނ�3Kk~9+Ij>ACB﷕dv����U�2=�)�xr�읊�[.4�@�\���|��v�z�pAn�뼜`�*=���
4Тrٜ����9*��k�ftr��C�`�m�Bb8�8��eпP��V��6髵�/�!1��UE�ɛ5u�6�#DȻ�r�b\݊�1/s��k�j���6i�*�jX���O��ټ�p��������,d�3���5�D��w90������\r��%Z4�kk����dJY�)����g��T\-է�V3��C>�#A�L3�ny2�]�>�w;m�Ǐ��U�>2���w��C�5�u���-���T:3&"w��^rYʝL���o�|'L�s�t&�)��F˛t0�5-+�p%ڎރ2')�{�`��śi�	��c����.V>#Ƅ���`H�S>�E~���x*7K5+��)QyS���'��Y��+�α~�H9SR�57y7j��W�h,�+g;gz�Z�f:ԷwR�D�MY�m��ڮU7�F�<�=]ܧ�����Im1Zw*��p2��*{���y��IA�{ETp�oܰU�{��/�bHe�_I���}���sS��׀��\J�����"z�8���b��Δ�!s:MM����I&(��{hv%���ۀv��F���u�u��-�scyf�u]��m�b�e`ZkQ��}x�sp���RS]�G��b��,�B�� �����X����99�n*6�n��wg 6muYս+n��Ic�*44:�T���7�1�������V�]�6�ː@���CA�j�}��:ŝ(�:�M�*τ����¾�h��ƭ�ڧ;�<����])1=Y x���$v�������}��kzf����}8���[�N�ļ�t���>Na�Ȏ�}qA2geX��[�f3���Vr
�]g��$�x?(oya`�����9��O��E�y���w)��#<A6���V�s�Y�ٻ����Ł���h��2��}-�YY;%���nEBei���VS�[]��8��>�v��VL E�/-����4%�͞���x�c���I�}������zjzL[ךɛt3M�w<�R�(��t��p�+\)�j�5b8@ӻJbI�6�e�o1܇r��p��oO_MayM^i؝VT�˓��i�6��v�MG�ly���$ouOW�_�GmP�����t8Ibt�!zmYmPKj'g6�9�*�;nQ��'j�t���_
� �����42����
͓'D���.��.�f�N�YV��"������.���R�-��p���3�		�b�o��"U]���8����ء�ͱ.��)]�He==��%�<�H,�GJ-v)˝޽۞�c�F=��3��qxr|��^<a�L���K/�]Zp��q��m���]kD�r�H>�NO�]G�o��ılab��{[���������&ty��ʳR�z��K�f�
}�u�uC��:t�|��>��*��&O�:R�u���9��b�TNk��o�s {�C/�xf�Q!��=��T����f�s������\�y����*��洤f�MQ�B�3�q/�i!�r�S��U~.�!�	�\f(�cP��&�d���X�a��k���������h�\M}��8�
���V���R�&�YX��|A�5�*J�}ڪג��Fh�.�[��V]�u6��&�nT������N�ܑ�%�^Z<P����7���UrP����@�V�Q&ͱ*�r�ۇ�ns��y�w����DЏ*��ُ��.��AgVE�T7�[������}"����*��$	>`��igd+=fS��y��U�����a���y6]wX�c�f����U�ؖk������g��$�-���z�Kv=��x3�D�#C��Ttߜ7�Y��&��7����У�q�J<�����:���|����@��|����Ҳ�J��T�u����kU��2����g����L���7^�J-L�~J�}ҔKl��Վ#��{v*���c������C��MQ�0#��Ȝ8cJѯ�W�R�o3m���53h���<({}�	<s$U����`�}��u��y+�ns���F,�'SFl�$��O=�"uy���?%+=��Y��.�,��{���Я��qq;����Q��K��t4&���I~��n�U@o������Ň�����U���6,�)q�G� �������ωe��&ۮ�|��A:�*v�f��d'����3-/.'|އ7��H�$��ӹY��ح/i�w���������ku5��ސ�iz�R�3|2����oN�������ww�2g���(x�L�s��/���;�HCg�t�#Q�j)���l�,����2\aT��ʵP���T �S���^[�mS�Y�"GN��e�^jtv�qv[��\�	��
ɘR$���l�V>���?[����q1����!8y��{�	�u9Hwl��o*���ƭI/q^��-dMb�4u�zŕF4�U����Og��n:8�{7�/���"{���L9եL��嫐���q��9�]N7Km\�r���2Zf���|��G6OEZ8�<�K�0M����g UD�����M/�`C_�q�F����T�w��N�Eע���}E��gO-D�J/\d蘃>���CWb�n�Y��m}����L&�rײoo_X�Y��#=V���i6�@`۩�K�����uiׂR�d����i;�3�	^؎�ŝ���
�7�8Ös�����#�	(�N����~�[5��4�D�f��2����%l,�Jx.2��$�%vX�Tv�U\V��ע(T�+`�dN�۷HY�N�<����5��=^y#�1��~]��.��;�L�4r]
z!�,����1ot��:`(�t'ڇ�J��_+���X�=�D����-���c�r<��.�grZ����`K��]��'E� ���cύз^\r7g>!P��
��/�U�}/uE���&N�qV�ڪ�&Gg�9;7�SQs�@�0�:iJ(�Y웡vr�uu5\ʦu��V��3�]άm�ץ>~��e��C
3�x�G	��^�T���d�aʭ<{RD��[{��Z���y�K�]�����+�qf��+L�ZT��
�9t��U�vR��Lǅ�<����+lA�D0i��X�m\�/Lˋ8˘����uȩvţ��r"�v�u�sC����ި����n�� ��%��p�?�e¸�P�)Ҫ�6����;���*z7h1�"��{��������9��mI�Y�$F��J�]jsp������{P�l�u������~IH�4���7��;�_;@V��^U7�k�ʓ���}�A�U��-z��Үd-�v��o��Eu��3L b��&vn'�)ti��[��������#���������ۊٿA��!�/��|��5J�׽+|ʱ�����CC��L-�C,�ffVN]:wN�w!h!��s��[��q���]�`wTt8��}�E'k�~���{��{�Sn�s�{.��X+8Co�Ћ>��
�ۅCww\ig��˷��|wu3�1����|�g���d�)fk]�qp�0s9SfJQoH/ҬL����nFD��X��ط"D6�o"�t��Z':�O�W�d�7��0�[t(�;m���Բ�v�lu�$����_Я
!�T���t5K.�m=~{=�~��R�TSo����O�u�OC�*��q��A�>����ޤ�������ƍ,ͣj�&��y���d;�u����q���8Qo�/�dֻ3a8�R�2�Wk�7�7	�+��)��r���܋�S�Ɏ$��hew��zw��੗�r��Qe��w,��ьPPw����&O �~^؄�k�Xb�\�~k1�]�xo��q�z��,ޤ���_uC!��:�7�?:�*�j�aXC��nT!?R�v�ȳ�w���86U1�czx����آ��VUV�9�Qd�J�di�J�����^\�K���6a߀���q*Pk>�	3��
k�ml�RС��Լ=���U�=�׏얄��Y�Jp��za\p����c|� ac779�&hF,�����qI��=�.�x���,vb��ⴳ~�Ļc�3�����|f�e���ۍ�1�jw6�+���̻U�?��u�7�����	J =���֡2xF�����lf-��&��+�@�kǲ��C�}/����Hc��F9B���2Ȕc*�Ϲ�'=�tel*�&�b/v��:�&\xB���w�:�Ü���ʴ�ЁS���6ˣ�^�V�j\���Z���(+�0c:��t���W�>*^y�vo\VH��)R E��Z�o^|�����]��:`���G����V��ꅅ�w�B�2���.�[��3��������QD[�U�7��)��3WS��������'�M���T���z�t�!䨙��򾱪pZOn�¹â�1U�O��7�QY	��z�#�B���]�ksv"ͬ�4MS�pV��G��ڜɁS����M�^�~��sw�ր����+�D�
�����TPy��X��M�P*|�`J��������������<.2�&N�	�M�/����99��gk3��p*�m�c��϶�o�����0�B����bP1�Vzʡ�y� ��9�;
:�n׻s����j�T�
G8�R�*2%�l��_�ʥ��ܯ�AҬ��(��_;؂�I���<��|\b
��F�}#h��J.$���&U�Bt��R�-�n���G`3kڬW��嫩oE����(�$0W��6���<��^���	]�jȕ�b���)-��lH�d�Ţ��N����ܫ�r�9���!-
�5C�b�1�V[ɼj�sw�Y�}��Eq'��i\`����d�G	�.P��y����+������i��M�3dΖ��zi����rő�wA�v��h�r�&XN����L��9O$D��ͫ�,�Ǯ�"��"X�g���x�4�a�(m��6�����̷�Zԧ;L��hv!Hy�w��g��J��M`ٙ"�8�f���giJ�ڹ;��}W��&u�����CS�59��xc�	nu��/�3����=�KG����ݐ]J�ѣ7�Ҭ�c��O	��l�>7v����	�M�ސ�zkS4ܭ�#��S�s��R�]FK�y��Ǐ�7F��xP����;Ȑ��_�'�ڰ����JTU�uy�Ժ�1)��Q;����B�����6��Y�"B�RV�����:#�9'H�걗�g�v�H��o��E��RJ��)�a>*^xeKt�ro]��n{[�n���NS��� b���Z��I��P�Lu=&LcJ�s�\�eF�'V��9�uл��1R�����B�Ĥ�pF�����M���J�5�}�9e��j�\L���ϯh�R��ۭۚ᷍(�Zs�(��Ƀ�)����8+V[��K�l�o]���O�*�~����׹_]M���s��flĿ)V��픉���O�j��m̱�wf�ḱ~.Q���X_Л�[�(k<���=�Li~�2��2g]x�}{�׮����6�ت�W�+����L,]�w�ɑ�wd��a$K�4��5����X:Y�\��.�u%��*�n���e�O���*̬�,���
j�t6��6�-]N��c��tU�u�_,gn���u���!d@�����fn�ǃD��a�� �ُ&�K�Me�� �D첻z�>T776q��Y"]�%uo�MI�R�dK���u"5�M�:��^���MeV1�D�c+*>w��PP�g%����B���T����T0Ӟ�"���F��>nC�%��u�逌�5�d|�TUJ�v���w�*k��(r�f��v�`��C�R��Ii�'|�1�T�]bP�
b]Q��C���]�q��f���v��5ð��sV�H'Yb�m�p^pVf�56���!���m9v�dX{�u��J��9N̺i.Y{1>�{[�V!�2�#��:����C�3�����͊�ָ�wWB�t���$������j�]kͦ���J9H�	��R2�<��Z-�[����n��x��C�c��l�ZBܤr+uד��ȍ*-.�{�:(��KR���>�M5����$��X��t�nU�]��k�sZB��j�T��4�V�����ܭWHQ�mj�sCz���c�Ѐ�Y�@Ю�pm�\�|F�oaC�����6p�Mgd�wU�Ci���=�Z/Uu�o��p�F�B�+��ݥ��n����G��זe��6�[%v��j ֹMXH�^�֘��9�K9V6Ji�\Pv��WG�*ce
g�m���Np9v�6;�YQ�Sw��|�ET0�:���X=��W`b��븡��XJ���@�)򊡘��4(-�/06A��*��$ջ���0��$�X��v��ltjn�4OP!{t�ӹo��3����V���Cثs;�1Go2��x�Id9k%��CO�ac(m����� 
��ܨ_W3�@x�q7�G\ w����ڵ,�04�:����`c.�b��м���oM�Y��O�)J��aE'uaaS�D�,me�{:Nu{��!E���o*�c��2�٘���n�Hr΀�V���NcV��Nt�U��]���;���yS5��1i��6@���b+��]0K�+���!71z^�z�t(����y�"�4cV&3�dc}H��k&Y�Y|S�@���؅��tj�����J�W�)�X��=�k�鉴h�ޫ�e���q�*l�S�^_f]]ھ�l�>�g�뗥���OP\
��`��h�Kz=瓼�S@��k��ki�uE<��C3M�(�ޚDV]����3������]���F�GM��1���>�V���u��41�%���,¨�n�(o�uI�{�,�:��͙�Y��0�u:�x����\�DZ��7�t���Fv�k���JX�9���#g(u^�F׸����i�..��3�8��9�3����(�JH���(b�	����a���*��(���	h��)����j�J"���*J)�"����h

�d&�q��h��r$���i�h��
����)*���"	�J���"
"i)��
��������)�"�(j���������(�$��0�"$a�������"�2������(�!���)(�Bh�T�����&��1J)"�$�(h
B����B��"%
��������"J(�ȪH����� ����b��#,��fJ"J"*����i)���Z)�`�L���jH�f�������3
�)���2�����)"�p��!$�$��	 �J��������5����O�8������Rq���I2-oWe
"���pN�� �z�(E�l���PLC6�2�ɧ���v�1�Z� !zW����	_8��_��K���*O�C����3]�C�1�̳9��
���U��ϻ����>�X�k������x$�6�W��Ή�O׆=��HPk�v�&�د�{���p���v0O���P�d�X�����0+�k���������阭o"o����zP��=�؝Xۚ���H�y���vs�m�r�f,�%��H����%s��
ܡ4�pkp�WҪ��W��ku�*_u
�CZ��}��n�w�Z��gW�^�����{Y�g�W	ŏ�y��5�ldX-�Bz[X��rR'9���xc�j�6�ɣ��
�k�SzP���wr��Ż��27՛O���yLћ�ZFk�[�(_B�Xe7qO�[&Lh���D׻�M#EM��@���b�^�x�4ѧ-�SÎ�t	��*��{�sα��r�E��*��9nU�c!�����ǜ����x(t�^�=�q���u����<��mv�1+���j���ݹ
�;��V4��T{h�Z����S��)������������&6.1X���^۾�t�b*��;j̖��l[�l����"�����btpt�r�肮]'�x늫��w)MVUie��uћ�ʓ��sn��*�M�UOaZ4�f���RA
�!K����4CC.2�V����ܾp0��ffaX���*�Dĝn�4�p՗�/�]�LKb��_́}����%Q��PO��S�@��{�Y��Q{6��.�_<�μ�Sw{�9PTHt��hry�����D�W�<2���%<�7��1�+Iū���ow��!��!���Z�v��!l���^�-�n�g�<GD ��I�[�=���^���l��ү�Z����%%��5���3�Ж�NJ����4�m�'q�;�Ղ�2�r�Ϛ�-I�ω�ar3�gVF��������S^|8F6�$UrYn�*������5�|5�5�_�����]��?j�����s�}��X6��U�j`�����Z�D�u]b2n#B�W^�<2�}��WS��8IseY��ɪ�vN�E�Mf�f�}x�������[b�6�xp�-���؇�i�bФ(��y(��O\s�*�,AgI�t&��WvSzM��$+�]�V�Z����Z�s[����M���̌z�v����
���CiT�+ѶHY���S.�1�À:��y{����|�쵁+.ؠds��ɲ�S�M�;�#IQ�a%�)�����[]Z���&�����s����VK�o3�=3�emn���6[��զ���V�ڱ#:�8FB�RT\�ݵ���R�\�E�9a�(	�C.��Z���[Vɝ��Y�v�-�ݿ(Gќk�Nޜ{%jʫ�xɹ|�<O�;]�
1�,2�7<��!�#"R�y� 3P��nڃ\�vʗ��fNu)�c��HQ�C�2�u�$� �T���v�F�w�j�>Z���4F ��!�ѝ�:lU�y�a>*^D0���HJ�� 0���E�c��?)�7.��+֏eg<�Z߶:4w }��9#�`f�Eze�*��$�u\qR�R�˂Y�z����2Z�x2z$x���|1?��Gܳ�~0t�v�N�<�J5}�t�'GЉ�:�,����X�)�댃%�Og�i���R�Q��*b��~9n��KH�<�#�w�+���������S��XW!p�X��]5u7�A�����z�)�z��e��>䚻랯�;������W:(�@IT!�]�1�����W��V}Ҕ'��uH��l��+)����G�U5DH��>�?	⁲���5 |vׇEG�EVF4#a��aC7K�+T�/�ks��t�Cõ�n��]G�Hc��#��
L�HV���c��[�J3�곟6���V�u�&:�暩\
�����]Y"��J��ޤz�h��}Wm�0��{��oM��ģ�:U1��,l���#�ݗ�Ɩi��r��W��m���z��Z�'cma�c\D�DIZ�h�qQ�iá{���g�5�D�ƈ���� �s��^���hX��qJ��޹�uc`�a�֋7�s�M1Wꋎ!��f`u���o��g�p�|���ۍ��XZ�b��nۙ��3x�9�L�Co�Y.�<�/n��������l�	ɏ�^�b�0���^�mPS�-ʫ����l~=��ݱ���n�ץ���!q���Nۣ�P�B�fz�՘��t$�C�b�i��/sp��n�9`t��13����Ld�6p̙;��cp��Wݹ�ݽm�(�;��W+�`ྭ��9l[6|�=6�/��r GM���>�.)�F�YbǼ=�⪱��f���|���6��T���R�k��y��IY���iu/�z�\޽�(�7�Qxw>Iq��dXx�S����Gl.;{{�weOu��,ɸ�6��o�u~pB��e#�_���d蘃��#�\���*:Z�˂��׃����/Bgzpŷ�f���f�ܽ���XȽ�u����1�%9�{̑מ�왅�j6a��-���^�������o%��*m[���.Ma\�f�Khu�9�:ۇ����ϗD�<0�
���s�`�V*��;�r򒤱m�z��kս3��&�s�x�����?o��ekOB��z2w��:�9�OS���3N��e=�w�s�-��1�����S1�l����et��@Kđ��ff[�ʩ��J�!ᅚ��9�.��J���R&�?XXeb�3�]��D5�*�+]tLh�{y��	s��/w��T���Λzj�:�����.�F��Qo�p/�بOe�s��/��V<vcnkX��� ڹ��"T�H�9
��ǒ��W�r�+Lխ3�l`���#��#:�O/Wso*ك(y�/'��K��3�N��"8�h;}j_����,棠��/������{Q!A���76+�~�ucn�:�`�ATW2eK>�}�4V>��ǯ:��'[���b}�n[�zW�]'��:g����z&�)���dv�Q]K��߯�va��5��A�O�-Ɯ���+6��+��V6w�L��c��WV�vҾ�Q�t<��xG�ϋ�F�(iug�!�h���2�J�X�a�	��l2��T�%���'^�,2Mǫ���k
��� �d���Aΐedt�	��@s����x�ۺw1�R�ǽ��`e_$�D��j)%C/�X���YZ6$k��$�#�hS�������*S�Vfs.�]�5`Dr��M��]P�������=��Έ҃����֏�Ǟ����⧣�|.��+]�Tޑ&-uz�T�h&Ts���d����od���p�:��.8Ǻ�¼�c<r�[�51^��Lխ'�=��얮�#Չ-*�M8�ҡ�ːw
n4,�n� GaD�ur��wGX�k%���>������7���VZ�'���<���{��=���w�� ��(��Wr*w�� ��k,� �]�h~"�kt��4nn4CC.2�V��O�{K�>�R�}/� +��s�V����6�5.�9:r�ڹaG�wf<� o����0g���^�P�K)̧	J��X�K�q"dhށ3����"���y�����h�����C%<��L�x����Q�;�rڞ�y�
C���̑�K,p�
 ��3����F4�;`7����.���Fw��:D�z���D�Tk_:JK:^؁�i:^�#��n^���s��&s�j�rNs���Ñ�P6��߾���`�w�)�QC�g��!�\t�t�)ͭU�yO�C�S	nl]I5��n��53����4�ԥ�\���^��Ee]�H{@���M|��^d���j��$V[w(���#�ԕ��`�i����X�y3�-3��9;��8��Qe�6�Eܶj=Gǌ��j[�A����^�ܤA�"���k9�	)���jk��~i����5���z�n��טvKBt�y��|5KT.�C�3��@y�j�=�ɀt]:�;���5+�ך�v\��XV��H<d瞺ŏk��|<�X�i��X�^F�;��M���s�*m�� ��&��(�
�vvo�X�{�p��0�K9�Y=7�0/d������{��7�zyR���H����]k�1���WyZ�B�L����c'��A\����2�-�=HL��*���7/��؅%�}����P��.��DU�[��wj��^(�a�O���'ԷO�d���-P�h�^;���+����ҐNL,&�N��a3y�_3���6F�]b���:� c����b��^h��y#�s��E�黸�/h�����0I~�����>�K�T��Sc�V����c�<63\#�O��
�7s�֞KƢҽ�ˬWh~J�@b��&D�bsQ�؟݈\�<�b�'q��
G#
ʍ�p��S�8_I��n_@�W��s�;�����h���n<3p���k�+s�q�,n�3��o;k��"�s��
;�(����r�V��RT�(���:}-��I���.�8�X�� ��J;hj����GWr��կ_^bW���ٻ�8�(�_���xB���D/�
qz�&KL������yP��Q��xd
���F����\{�&Z�=�|-�zNJ^OƮ�!���ġa�S�Z�w�}U���7�����9��.,̩dd��J��:(�RU|z�o�뢻��0�,���q
��^[}���gN霈q��~��a�ꦾ��������#�h�����r�ᦎ���|����6��.��`>y^�Ӟ@������u��y+��qdb��K����Y���|֢n�KU"b�Y� �9��eg?E�-Õ�Ux�Ay� |ՋηN��V�_�������x�Y��%{q�_�u��d�p�|�ĥ�����A��6��7wi�oy�T�.jʭ���]�v�I>�d Ƌ)v]��#'��]hζ�N�L�4�ٸ�a�z��|1�97WvGo��ԟ�hVg��J��&o:i��'=n�m�:5J
^���Ǝ��b��ᇀ�s�	�ɸi���v_
cP�P �{��o��t`����[q*1����+�s
�sul��M��*���b�`i�a�;H��wf�":���]���(�ܭO��8nQ:b�����:.R�4Γ}/�ea�g+W�S3@���1��֥,�#T^B5w\��J����Z� �-M��ӵ�g�@L�V@�x�B�E_^�|�'�s�E?�P���D-29�D���'˶���岊�U�e3u6G~g�������MR���³��틣Ys��cSs�����odB�����m�  ˙��h������}M����C��y�a�k9gW!h��p������c�/أ)E�|�=�1ObG�{SU�va�1�-��eﲶ]��|�W��P���__OBϾe->*����n��|髉8v�+��E��ڼ�On�`��7�c��-v]�ٔ���}6!)w���$���g<�k�=�33׾^�.Nw�6�������uV�wH���aa��Ya)��:!�8p9Uq���h����������X=�/�p۹�D�/ª����;��b&;��-KJ/ �`m
Kqt�6��p��C#���_˝�F-l�	@�1��i@界qg���{^�gU��|�ҵNv��[��:�(��.@�>|�Dʰ�lR�%�x
3���>��X^;�C)���z�a������J�-��¥�ӧ�d0��o<BN)9�im�p�IY|5�˓��p*@ݟZ�IfPVC��rX�ݪ�͘�=����*=��kv�P���α9u����}�[����\��9��d��ر*X����b��e��Km`2�̝��'S0*9�Q�,_M���V6�*v%Vp�2ǌ���H���G��4�r�zw�cs�����)���O:]Yx���}:�E*��(�]���[��wu[�;/��)���]yD�za_
Z.8ӝc瘬�\^���ϫ�w��ƢN)9�p����=ǟ>,[9��g�*��|��*��p��ɶ�T�yK�<ܮR�F��n���#ӹ.�s��P�[$m�&�����;#V,��/����[�J�;��LڣN����J�s9� 4�'5Ll�u��l�<2��ݎO�"��^nc�N�q�OM\@��kg�B�M�X#��� l��S'��5�:�HMy���ɼ�c��C�ުa���T�Y���᧢��s�ll�c�=Q��MU�47���d>�Vw����Vd"�dX$V���΍�Br�ob��|Ѽ/V0=�۽)��N�/��'.�S�*�l�0��WL�}�}f?��`�^�>�Ι)]|��!�t�[ڶ�%�Q��cSsۚ�{4�dej�+�ks�阄(����lN��qV�t�Lc��Q�����r�g����	��"�n���w*ǯY��^0�(��9}�i�Õ��A�N&�Rh:D,����#;����d�ڔ
�n�V�^���7ěr�V�o0!S}#״���b��c���47��o[q�Yd����8����ڽ�)M�_5��4��M�t�k��[�j�ª�1���S���]"����(k�$��<��N����bĬ�:���V� �}��c1J�ٲ5G^�(x��%�^_�b9W�U��u�� �ws{Yin��toN�C'bAZ�s`��'��b�u>Ƒ8��D�c{��W|����i��
���$����z��t��_8���I���&��}�u�-��Z�#����d��j�)`���*U�V�tt�-$g&�ŘeaX`)81��J����w�W9+xh�Nr�-���gdr�.+���9�1
��M��D��wB���^$F��c���u}O�Ys��,�(=�3�ᅪ�:��Jf���.��k�rKtl\�Zb���&�Q�i��wL'G)kuN�ٜ�N�\v&R�e�U��Ӽ5�
mRAoL�JPS}1�3u �p�̮}e��	�f�2�[����-������8� ��2F�l+z�%�vɳ�Zd��&Z�J祝p`�wB��.��V����Ы|��J��(�TnY��^@�\u�r1З5����T	�{Ƕ �,k�$�W�v1�W)�$Y�;Nsz�rw��T,��+�j<=L�O�[�Ǽ�>����vV����Y��/�ݝ��}f{rGaѢ�f�].�Lz&V!��#j��ṘQ�FF��Xea�'B�5x�_M�f�Z�gI�'Jl�Q���;��^Gw��F)�U�9��4jt��=w�rcͱ:�=ƹ�e��d�W�I���|��/p���8��zh��*=�I[*^N:4WW���t)��Kޢ��F�������j렦qRjmv˺�� +!���nel��6�]e�H�i>�fC�~[)V�*�B�ݙ��S huӘ�}���yI��(=�r����Q̠�2�ǵ���^�a��T�$�kh�m,u�[˰C�/f���!�G�Q�2�b�`�3�N�^@w\�j����Ń5;5��YY��:՟�bS�ɯRm"Z���Sz�X,�K��j��3GD����R�t8�+�}J�nՄ�� I]��+�2�:u��_*�{�/o��[�u�(�v-��E=��>�d��rr�-�
ԻڛWvb�Tb�*������9Dv��Wo<܋E%YW�
�f�=�RlK��֩�$�Nxs-(��2_��Kon'���[؈�dq�5�Mb�׈C��O�Y��g�����6{9�.� �7��bR�W�6���w{1A���'�[Ұ���>\��к��
UB�Z����Y�QT�1D4�CE-D��eMQP�!UE1L4�50QKE0QPMZ�0�2I�Zʂ
 �s1k'5�������]k&�Ė��b�0��j���%���,����' 0� �f*�ih����$�32��a�B
,����`�*)*&�h�"`����ʂ`���	�U4R��U6��(���H�0����dUSTQ44QTUU5MDRRk1*�
Z�"�
Z[1�����l�Ɉ��,*�������"�Q����eM4�5�"�j��*��,)�'"j��f5#Tj2cVMP�$DUYvo%5��-���]�s=Je7�V+)�W�2[1V�mM �AyU�7o��[����Ï���I�����۶��:K��x��A궅؃OV]�xZ�C�;��E��}���9�>��/l��s�z���7j��>y�p?<�xj���,R�F��mQ;_y8B4��e:3��Z9��0�S��[��]cj琩��B���w���2�\k�Β��F��s|ϾhK[��c����L<�&{����L��xp8"O9�_ma��o��udmr��iT*z7���˝K�޼��մ�����(Lw��/�ul�j�s&:P����Ta���S�{^�����w����Y��^���G:�Iz�4�ͦ��$e������	91U�;�R����g�.'n`4�MP0����+N�"�����!�yC���/�^�ݫ@��=����ً"�/f��_�Rפ�x�_l���0-�08�����f�h׼>ݧw�!Ivc�b}��Gf��l�fgf{�äM�.e7��>o��i��XZǩJ�$����T˃V��B5�T�Y���M�R�=����A�1�..�w7�^4YF���}B��[mP�9�pn]����|v:x��H����X0���7i锑�J�����O@y�y��y@f7G�՜��C��R��2��V��t�"*ErC�Wm��'���γ��E}��mԮֱ-]/�"BM�݄��Xp����黛�Ȗ�I�'ؙ�8��NR�Tny)Rӭ!;� u�s�9�дU���N�b}ϸl��*�F�tq��C,R13s�6*ǟ���x�:�[٨��fۻ��v��o2ݾĻ�2AqJz@��p���1���J�<^;O����ᱚ��w]��P1�KN��D����O�'���3�E�p2d�͞%�sQ�,��6,�d�nt4���ܯ"S���qt��lc�ۮ�)m���b���=���Ǖ��/�^ww]+uc��oyngE���ɖ�XJ$9ښ��1�B��X�F����I�TuL=�	���j��y��U�`zJ��M������Q�X��a�%P��3Z�]�A��z��o�m��������{1�W�E�:�����J�%�EP�Dʴ})K|������X���E��v`~L�DMQ��\m��k����;*���p1�"�Go��k�,/�y<�_���/�]ۄ{:�Ld��-%,�~;��7��V~�J��0��ob��3z�*jd%]%��9`�U�;6�, �S�J��S��Zi��iK���ڇ�/jo�����Oz:--���w[T���Ģi�S3J��5w�B�?^�$�1]S�\&U��Vsw���X7�;pֺ�[�LAl��󕙁���]����6&�6�E��ڊ��T4n���$mƕ-�
&s�&��;�\�l�ԇ��y���L��#��ӫN���A�(��ܘ{���e �XA�ws&�6ɿ[�U���+��'�N���&ʳ�v�0�7�^�hɴ%Q��v	x�]d��������2��`��Gbط��sta�'���ܯC;���T�Y��'<�(a�|p\�-�r����U
�7K����Cqb�S���6|�n f�b��δ��;]�4ҹ�U����H0�9/$T��R�C�JF��w*O���]��
UpMއ��]4Yr܈�$��7H Pe��cf(��%d���Wܰs���R�l�6k��\�G�C>cLt��a^*���ч8W0'�g��10��}�{�cƺ������ic�Y�3��ʵ�r����gD�ű1)vQ��f�`'����v��Q�їܗe�l"�a���(Ϟ����)���W{|��U���#���eË�ǆv��.�Wy�32���5���)��2��v����*�nt"<��p#GK%�76]�p����dͿ�N��+W	N�=Fox�wC
�2�r�o+�_V]��8�:T�jj�y�J�:e����nVevu�k3�a����rL���"n�7����kd�Nz,,2��$�%v��{����u�ٺ�����{��D�H����*'|c��
���.���Lۺ�RҊ�G�����Y�{%^�\�dĸ�@����
�]�$|Qg!SS*㳵眲�J�8{zʨ�ޭSw���3#'ˁ��¿�l��	�(��h���Dqx�]�8�ڮ�l:�"#�ެ;��F�ӳ�w7�ld���	[����M��������{����.�!�~�\�|����W."a�/*�6\�U=��>�5>
ٙƞ��5YUXJ8`���^�gm�}7�M{�E��-�	H�r�}��:�Ri�c�d>1s;�r_-�n���ܷ]�B�gxT�4���"��
7K=�8A�B����Vr��,���pTZ�1׆���m��/۝,v!֬��]c]<7�듔��;V�^�S5��V`nkU��h���1�T9�z8�y����bS�c݂Y,t�q���2�謼&a��g���y͇�In�9R`��w8�h	�}��ȶv�ZF-���2�gt�.��M��M�j}a�&;mL�6fE�l��繎�*bID�eBڵf� �V��YDZ��O1C��X#F��p����>B�wb��,�ra�V�S��}�@1o"h{:�dN��Y��SÎ"����eu\��qonm)~�m�J��hpMd��E��'����K������=�q���]�c�=n��%�T�,��bY�:��Z�w�+�XwJM4no�!��[+E�WS� �(k�<^]-�T�$�Ő5�0 �8�@U��(J³� �[��<���f�u9���ch�H��e�sݝ�Yv��{گ�։QP��<-Q!�C���Xo�
�]�s�'�d���ȍX��p{ۣe�,��*���㫈Z�)E�e$d�D�'E=�u�|X��D<!L�-�Y�fW5S�46<KA�_m*�H�"
�}~�y󤤰ѣ��s|�;ʓ�╷���5y[��m�&T��:��hk�B�3K�	ru�ˉ�������.a8˼���u��7'r��˓oE�'�����>t���������Lx:�%1��d��bt��e���7h7ێ�<���y��YR;m��G�_�s�Y��e��㮄�YVP�yW)g�җn`�nt9�%��S֐Ɏdl�r�9���{]�*a�xw�J:i1�!�z��S]�"ߐ���v�͐�a%��>��7̹Ïk�Pb� �g���8N+\7ٚ�mi��
Ҵe���#4�/���b3ٽ)����d�Kj9ɧw~�.�t�5^`�kF	��%]��)�ig����v�օ�Z��oj��!�)Q�>��{�<3b⯯֬���XK��!\�J���o�	�>����ۂ���Uok���#�ks���G`��7�l�g�gnޜ�H��_��a��Ӥ����Z��_�+2w%�n߰����&O�uRAb&��SbЗ�ln	�ԇ#�Kp����*��n�ERط�wG�#"R�&\�L̘�N`�r�£s� �J��i{��P����;6��3z�J�#�q�|�Щ�
� }����tث�W����ɷb���tr-��r����Ҋ�>�/O�7�`5�a�֫ZS|���v���4���;G�Pvdr���y���7������S�1x�[��g�`bsQ�؟݈\���ul�ŝ�r�{Iܱ��i�/�����u�
����L���A��[�z�H�D��HP�픵�Ӟ��z�7}���T���g���ΰ�\�'v��1LF�W!mՀ�{A�B�D�u8�t���=���Si_[l�{��[��;�Fp�\9�1c(���r>5�$k�k2�؁����*W�7�b����{�WW�}K�d%k��\"�d�J�4��E�:���C��A*��F�$��G�K�p�����_9I��r�'&��q�1}���=�Z{����8A�ZvV�reg68ϗz�o����vӥMM��{���\�ظ�2�K�o�:Xa��9��MP#�R��N�N�^��I����ybVdp���2�	1���+m-������VlW�v6��U��o�F���c'����*�T�C�ְ�ʬK��%1���X�Z�1��i7/{0�*<�c\�QMhs�Gr��P�N�Dg��|&�<^�k�U�၆­�Vx�/�\6�ay�UGs���;�ݟ�e+ߟ��~��<�u�GK�'V6�n�,��fa�ٛJ��R���ϒ����@ۍ*g��|�����ve��>g&��H�_�<�u+�E��B�|֓ǟ��;��䴇9٭^��f��9E:r��Us������]��q�;Ye^�w˳2�R5�)��`��~V`���.i��Q+�*�S������*�a<���V�'�K��|;.D�=W)�(xd��b�E�_�7ҥ=ݡ�^<��m���T{��f�d� �o$�=EgvЂ�s�l�&
�Ҝ�+r�䌳C*����]bz�����`�Bst�q���ʢr�Cu���m��fk�F�R�f��7*N��{��S��ޝF��O�(5F�vObKIETS�W7N����GI�u6�n� �����l���z($��qɱ=�!Oӭ��L\�2}��e��z?Ze����|.�^̃��ч8W0&af�q��o��9�˴�?��6A�!����C;�4Qƴ��X1P�d��{m]SZ7-[�יx��-1.��TM���s�}��a���}��*�}6!zO�ߪ�pt�N�R�҂{��wt�U;n���l����J����D����b�I�~��ĺnwf�L,Yj/��aeh�,n���#C����_���R�Vv0�{�߱.�G|�fN'GU����m�*%�&;��c��B�Z��c��(E�x'�,㞽<:{}����e�v�vIp��Rc�D�ƨ��AWl��	�(�ޤf�N��gA�aU���| GaD�h+s0��o�d�Ӟ�V��eV}���	LoK�b�V�v��I���Tu�J�^����uŁ�r
�t+1����㏄�Խ��9=)���w���.���50��SN+��#ڻ�h\/9-4�(�v��.1��X�)��Aѵ��f�Ü-EIP��:^����{���9!6�?,8Tp715�����S-,�ێ�MJS�Gf�YcY+�J�w{��bY}	JeA�N�WsfJ�{w0��s"K�ظʀ�u�-���7)}��L��u��pȬ	�P��;���g%}v֥��
Z�wEcGxTߚDP�k��x*7K=�8A�g��b	������"���� u����;	��ʝ~���n�-8��NUl�D�(U�*Û�d����>�dܯP���U
���mGv����s��~3,mCƥ�B0ܧ���=�7M��PKlﻨ����_V�k�V?a����Bd�EMX��F�yb�Nʱ=� �3
$d���xu��*�*�rK��Eb	����5q�5���'�y�t�\#������ݞ�ٚ���]��F�­W��h�"�&2.�I���膆`w�E�㖯>���[\p"��6t n(;�ķÙ$�SKI�}�'���/�K0y�t�4�S�\���ܛ͚�������.�p�g��>�B�^U>�t
5H����b	���vL�r��֯l�燖����5{;��B67��<�:8�g��!��d	n�������D4lu��滇�4�$�o�c��&��P+'e��ZM�-�rjS:�>����Ǐr��8����$�2K�vX��w��u�.{)�����6��ܔ���Gaŷ*)Mn+�z�95:csd!�={&WB�\=|�x�|i�7W����h�;7o9�v�qT`C��;��3V𨙐���y���a;�;iP�:Ȃ]�oϝ%%��7��$n���[��ӻW^�>he���~Q(sk9D�s����C%�>�Oٝ�
��5��X�t�8�i��9�6!���c�ڰJ��j�5�|�9Ș�S�'���Q��V��:�ݜ�#���ڠ=�i%�g�#�\Jy:g��1ڑ��}��Qωg�(�w_??\���˚�%���d/}6���y��"xv����ᴳ�!����v>��/
�cu�5[k�?M!�9V�^*�[c,������x��A��]���[6:��1a��S�u߾9]ku��xk}��0����bϦv���gٻC.�2�Pf��goe�SgM뫛�1�v*��O�T�De&&O�GU$B&��Sb�C��#������㋯]�.�Yؽ�����4���,��FL�1��8����$(�!�
�Szd˼�K9�̴{Z�\E��H�&.v�Fߋ��a�C=)N���i�[�r����U{�Z�?���=8��RX���l�Z�r�Ύ�ں�W��n��[�ՉJ׃Rv�ЊbM��Ȃ��Q��!�����M���k�5�P��p�v�o[K�ƀ�
䌾ԚՆU˦�cw�����\��0j}3�hg6��Q�幖�jg]�/+^s��[��Z+t�@�f��%b%rz1�8Z��]u]�=M�n�4��+����`R�g����w�7:u�&�b��k����%��۔9Ԟ�9S�s2��S�e	8��b�ڝ��$�wOƬ���2�q��H��twL��*Urw5VcMR�6�d��Ow%�����!��] X,�Ǯ�6�%��h����� 0������ʜ9���p�	��ǲY̘�-��]�sS�	2�m��og@���\�.��{pv�AZV*��<6��R��ԫ���%p��Sjna��;���h՜P�;�Q�f�;e�����ȝx�Q��2���@�ɱ-�mi�[�6��B��1�w|u�K ��R�;Β�4�������RZ�Z���^�.�]>Kᙚ��j:�J���yӅf�ڽ��V�&�T�����&)m�b����K,$��c��Sm�tB��v��T9�u���K�p�rd<���k���C�yRWNt�Y�
f\��kJ��;��9�^g2�7�8e��R]���z�wPCkter)g*K���ag,h���j�)N*P���ʜ�+�;��XV�x��P�p�pC��U�S��:G%t�3z��p:}���wP� :�f�]q쵷x�YI���]��V�"6��.�+.�k�����s���J�
Sy��gn����u����>S��Vv$�kBfT\�h�b"�1"�{*��o5���D��л64��WuId�:��z���tx�Q=�=7z���4u�ifRu� �J��T�n�%5�^K�9����\k��d�m�k{���|�!�!�ɘ�=��p��M��{k6讃�fkO0�G�P=����(�Tڶo>˽T�wu^ө��M�8-n�%uc9�̿f�3{ �V@ru���se��`��i� ��[5i�J��3*��M�~�Qn�k �v�ZLep�!��mbx7�v�F2����]B�D���o�T�rv��j��-a���k�Ķ'z>YA�sh��l
�j��$�M
X;S�|9VG���:��J��Ǽ�"�iU��8B_M͋�ڹ�K�Ut2W;ܦ���%�3���5Z�`���������XZ�lZ��� ��pڠ�=L��>Jɰr��{��Y9�-�l)�6���(ܮ��a����Tg䫹�֪�V��i�8�1t�G6X�
����CC@wmu
�x9ӥF��{y��u)��ӗ.w]�s2;�kqqH���fH��┦*u�:]�k��=>�~퐯م���D�j��r�)*��*c3-XQ1TTdcUԥIAMYfIE�D�dY:�eLISTjri�1�&*31r�"��30�i���)�(����"�220��̊&(�(*�H���$�'�2��$�,�fT�FQT�QQLQ$�Z�31�����0ʪ
(������k3b����*(�����,���h��J1²�(�����I)���`Z�)�"�,��h��31 ��3��2&b��*u�LSUڲ��(�cfaT:'$�Ȉ22Z
��̳&���ʊ,̚��*����`�L�
�	����0��"����2����(�0�����):���n�Nќ�=���o�%CeL��LwH�%���lK����Ռ��cO���*�*�l���B���!d���{��%bX�|7԰�/O�s|\%�تSJo��0k]ҥg�\�b�p�܅�W/ϩL[ځ�g���Ģ�2$x���}��؁5�5�gK9|��ϲ���%ޚ="��l���g�S�b�t�4���'�\^��2Zd�&b% q�R�zt�ݪ��9�}^����ʨl�YՑv����8� z�\�H������h>�qg�<V/y�ɪ�5�~��<��h}6�D��Vf#���+��FU>�]����G�&�����؉yb`������t�>��أ��K�\�m#�R��H����.�+i���v=U�jeZ;��Y�ڢ�� �G=�S�6�K}��8�fY�^u]��l{f2��ފ7�어�p+��#S%<F!∱;Ԍ�I��D^�>��UŹ��r9�]�*%e>*�Ĕ�}Ϲ��@��OV{U=76y�g�nSj�^?-���{�����o]���zx��?|�_<zaϹ�g">��<��X��L�s�׳]�Z�݊;��
!�`����f�jjۤ�b��m�u:�.�kt��v^�O/:�[1c ��Q���K������2NQ�p��p�9=��pG��U@��mq��]Lt8ε'}��Y�t�ps}{��E�j��fu�<���5)N�n�M�x8�;@ݥ3a�r�Us[������7�}"��}��zVX����'9��^�\��%��NS2��c����i�cع(a䙆��Ur�^n�����4�R�&�����L(���\�x)���(T��l/��t_=�I�T�����;�׈⚰ѳ�q�o�j��~�_E�fYLÝM����~��vw%u�ս�}�+y�s�=�pc��;RG==>��4.3�zG�*��O�=�M�jbY�ܳ|l�ܻ�ם�y��"���=*jJH�-�N�#l��4�L\b�!���S��q��Zv������]�`8�H�j�\�g��tFr��W�����YKO�W����'��{���b��^��ڶ7�w�������7n�~����X����n�9g�|F�����^�|^��"V��$gs$���m��<�|�V�v"ns��c_�)�|7mq�xT{c�W�˭��і�7V�o܏y�E�ad�x[n�؟W��w��L�}����.i���>�W��q|��]����p�7իt[���wp<힆wh�4�_T�k�^Xg`����g[v(*{u(v�؊�Xm�e���;�٩�ty�Z�_l�f�e&�#e"䌹��"꺊�櫁�UѪWy-�.m���ݤ�K����3�gC�Y{��ZP%�l/�tMw a��H�1kdx@B��^ҁ�+;vȽ��3�ٳ�x�p߳�GJլ��|�����AP�x��]j5_>�#6�N��A������}=��v6�mN�`~yjW������U�b$,�s����W{���5�ݯ34�/P�^��&��gw�����h�j
�
�Lx�]V8�JԽ�V���h|WO@,m7��s��Sĺ�.�OM8H�U��)UȜ���t0��%u���@zmҺ��E\�l�e]�B��8��Ӯ�+8����iP�|�*M�8F٧1<`Q0����U�`���Y:�oxz���\^0���>�Xz��^�O�����1ز����t��$[k1L�^+�>����u$�ѫ��\�>x���t�1�"Y,t��-E�S��m�'F��~�IC���~?=ˣ|��z�*j�4�P��Ѓ�Sq�`���s�
n��{�;��N��ڿWc���Md��jT��Pf�HU�A�x�^=�q�7W�Y*�o���~�=Kz�e�'5����e,�ѣ�0�����{i�Y9+X�ʼu�
oI���:�u�y�J�Z}*a��qImӔ:\��w+5g�M�z34���P.e�%_6{�����+��N��;;oVƸ�3�*� �uGLK0�;Z���dX����w^�HWm1#�$缸���}�^���U��+Jo�(�GP�J���
�Ԁ�mY�Η�`�)v�Mf��.������K�
��w�q�ފ���QP��=��$:C���Ykh.�u�FH߳.�����Je�OV��
�C�K��7��X:���,Rb�%���fxا0&Ğ:���r�ڭ9y��5a�ÿeL�:�I�u�o�P�֘�#��+���5�:JM�m����Y��[|�'��Y��v6r��!F�_��K�}���q'C�%��î��N�a�u{8�l]-7gh��]�Z^���`�ce�X"��M5]
�m�r˗�ʼ��d?N�1H��>e˸Ef�j��ř�����c."�،�����6a_�����^K����̜���3}3�k��=$�����Ֆ��4���<;	YkZ��_m9�r�I��,�

�U�5�.9C�"�Hb�!F;ɴ�j�@>{��ps�*z<O���Wz�U�J]���,KbB�ݘ�xIf]�1��|�W��b�ݔvD�7�p�IZjm�1�ru���-nԀ�;�к7Ӆ�Z-Xz�B�30׊e��Ez��Yې�-�c7�*�r�`�-L�zV|V.�e��Ö�3{����k�ҳ3r��զ�\�^��h�Ԉ�'�-�2����K�= ��7�l�g�gH�����zM��i����}��nr=��p�ʙJ���ײ�'�#X=T�Y���؅%�}��5��۫�nm�I�9͂{��I���j�FD�q�˓��������.Tny˼��0�u���}6�z�x��wK��P�b*r}�Tf�G�l$2� q3s�6)��.�-�{���_#ޫ2��y�u���)ː0�S'�*�T�"^�eC�~h��,��f�=��W��幱���=2����j��q(�p2d�g�c������^�F�Jvn�Z���s���H3�8�K��g�<�� ZK����1��m{(̮Y���#kĶ��~�v���\�T�F��nYՑv�O{�>q�C�%pB��Vt�a��Ի��]�:ߡCK�/tB|a���؀��Fǰ��8s��?���n�;����f���Ѥ�3�Ϟ�*s���Z���ُ¢��R��*�EЮ�>�,��&�!1{}2�v�m)	�vMU;�LjeWr܊��z��e*YR�H�����B�����@`�E�+���z�6��
�wb��)r�=s�����H����pKC���,�2�3��a�5���JJ˄T�C�WJ��$mwY�ZN=�C��F��q�n�M@�&v����`�_s�,[TTZg0�xm��k�9k�Zɇv���WU�l{Uoaʔ��c����A�}��nr�k�S�}�b�!��#4��dE鲳��ͿVr���d�&U�hż֝���ô+ q��'_.�7�YBW�E����cZҞd�[�y�~��i�UjQ�Y�=��9�g!�8������{1Ҟ�,�w�]��Y�7���L����r!|<,QY�&+��ĳ�eq/�sT>��/o�)��z{U�1X��@�}��s]	�+�=o[�5�v�#zC�e��^o����j{'���=~�ئvz�>}37c�G-��9;g��L��;�OVjqX+����S���|*P�.���@���@���݋�*բη��)®���3g���+L��*��
*�]Ve���:�!H"R� i}˶	��T�#%=�qx9:��Ҧ�/���$��|� ��9��ZN��l\���]���~�ս����;�5<|��1Ҹ��?`�2�YCH���E�|�=��x�J�2�@�� ;7��}W���U��m>��Ui���5��](��/U�D;bڂP�v���VQ^;Z6��V!ol��(��)$J��wrd���)�����WU�L��z�mISya�7�ĸ��.�:�t�Z�44d�3Bi<��u��<���}��V<%2ƇK��Y��C|no�=�YKN�����
���I|�u�=,Y����Us��t똘>3:���A�Y�>�3پ�ʹ;,u��w{㷳���*��LKđ+�(�#���=��*�k�D���,2��.XcG%tK�Yn"Bߦ�P�N��2q�Q�u>��@nT>zm�b���}�gl8맻xf��_,ͩ�q�	�V�Y�Pؘ�%����j���t��|*E��+7��f`M]m\�t��ͭ3���460Rj���Tv�<@�#�q�~���v�7+�N��ti�聿��/����s�Z㱻862BaS����C�2�M"��6��ε�wdI{�b���>�@�y�c��uZl���z.9�λf���RZ���Un&a�6�����_�=��j����t��	�M7C���?�=6�xO�W�CѝeM*�w��Jv��<���謆��iC�Rx�6�ӐuU�|��8����f���)�h�A��ˋwQR�E�{k9;�V�bW���]�OV��;m0�=����o)@|�z��n����j$Hc���C��ފ����VeJ�'��K�0�$�6�X�n��; �͙�^Z=�2sum�&wn@T�:IÀ�ʚ��ő_/w�M���1�ņ��ô�[9W
P�q��晣��d�$����T͔�yRz��NjK܈��I�x����i ����	+W+����n����̫�._���g�T�w��*�!2}i5p!�J��.���Kzb��O?;� 3��c�sŚ 6���U�����Md��jT�cTé˸�k8�U�*�t��ٗ\�A�칲���;�ħ��z�t8N�FN�Р���Ȼ�&)�sq�;�KO;�]o��3WhUy]�5g3Hה���|�\�.�O\�I^cI���^���/�Xcӯ��[D'��ܱ�^oa�L\� �W�9�Û$��ށ�'�Q!�Hv#_D�,'�׏�_z�m8���z�cY�.���ӫ���T3}<%�\BԱJ/)#'�Q=�6�ډ�6g|��g95�j`H�;�(/E��Ρ��3[%�Bm*�{5�Pw���3n�8�^*99dd��Ȇ0:��b��B�K�~'��t�}��N��{XF�[%��Z���}Ӈ�	GwW�D.Þ3��p�U�h�'r��S������/�"�^�[ю�D��Sp�x��B��9�:L.�h����rw0����T��y���G��5*$EF�\R5_5oT۬��A�#A���cpR*�Ԃfu�����g^��OM��N��`�n�楈�:�~�����:���(�j�>X�)�I��g�C\��6��@y+6=׺p�z�1�_p�d�2����/#C���BuYS����E�s���e���ζ�J.M����'V��ܴ�})�u��	,M�d/	�e�_L�Ml+�E�-�NK<������bՐ�w�d�^�{Iؘ<�!HQ�,w�p���SmTh���­�J
m�-����_r]����w���-�2������#�a����g�>�Ku�ܺ�f ��`��j���1�{h�[�JW
��*e���o�&���P�r�n��D8�|�����~sK<b�3�J:�W��+|%��pw���!�#"R�&\�L̜t�p�6�����eǋ]w�����E��N���� ��&.v�F�G���DX�&nld��� 7�Z��cH�J����|T��0����B��%+���(q���>�U��v?k�����Y���Sg6��n��$�guB*[z�L�q(�p2d�g�c�'�O��e:Cx��k34Pk�t���
òt�ԉɻ�0��Cj�{�8x��m�f�h�n��>��'���t�&�	7�ϖ_olҕ�/�����M��k:��K#]	#d{\�u"�?mi�-R�/;�=n���:��\���Z�	̟�w�w�8o�>�ٱ��f*x��b�ݱ	�`�e����ulUbB�ix�������_Z'V8F0�{f��|M�|T7].���S��v�;�*nڶ�y�\�� �N�yJ�M]M�hrj���M��fb��vVx�v��vh�\�ߥ__���F�n7Z49,Z�=���A�ϺR�R[�QŃ¥]�M(V�E��w�$�\ŏ}�z�Ԩ-$�3�WDʴg?�:�Qg [��Ρ���c��,q����i��鰽0��u������@cT���9R=��Gb�!�'z��i:9�zl�׈�K$�or�.׶��۳�z�l��1�2��hP�5����6S�f��������)K�j�΍��#m���;�p��al�a�����U�͋5���ܙ��<<p���y2W�}�$ⓛ'3=�h������}��b�JbY���nj�Ûؼ9��xWx��	UY�ǽxo����_D�R��璲Ό%v,:り���9ժ���e������
�+�(* ���* ���TA\AQ���+��TA_�AQ���+��W��TA_� ����D�
�+�* �j
�+�PTA_
�TW� ����D��* ��* ���PVI��^�	= "���X���y�d����y�P���% �����TQ��C� *#lQ ����4H�T*�ص����V�d�ɭ��T���-m(�e���vl
w1hp�[� t  �
�rk�IC�ʢ]TZ�d�l�3I�P�w
�2$�J	+e�Q���h�lcm��-U�ԶH�q7X��ki�5�ն�KmRurZ[b�յl��`��٣fCF��m��    Od��T���M0 i�F�A�hE<0R�IC �    �101��&E?�H5aC@h�F��hѓ �`A��2`�MH�L& �MLCSjb2mO��J{}��{���"��B�<�I$��h��.J>��H{�IA%� �$�-	��@�II���O�?آ����PBK���A)�H�I$��IPB�d�i	$�C��Ϫ������}�O��BI ��l�b�QQOŧ�~(זCx

(E�������ϩm���mfض4��k6�/�U�r�Ԇ�)^兲-yn�6�۵��x5a�ئ��XDvN:x�Zc���oh��7�+�6@M;�6[��&��u���X����T&�SHݤ+[��&�YC*kw�1�:��Fn�#�v\�ZA˲ҡ�\�&[*�Hd�q��"&-x`���*t�Ć��z*�#�,V�^h��%�RT�����\�5nΜ�-��{�E�+c̤V껡��U)�k&�EjU������p-4�3%�\�N��˙��h}v��`ջ�e�*��"�0��oLWZh�U�h�=ک������<޴^c�wV��o5Y��<�,�l�v���A�� 	�J�������Rӛt[K.�K� ��A��֞�B���A�\�������7g0#v �qU$��m v�&~<Z����n���1m�;�[���u;x[
�������ݥ�N�wN�mcwl4%� :{qm�{_�i����f���6��8%�ǂC�Y߈yd�+.�*������+M6p�ˤ����3{�9��J[Uf]a�"4�Q$f 2R��VB����I�w���)�(T��8E���^Cu{���H�b**���u3d5��c�V���%�<��G�gwHL	�2t�q�ֵ�RGVM$J5l��#q���*agFE�7B;d��!V�+fK��(���Z��CD�[�H�X��ޜ<����T	C��+W���w[˙-�F���6�7f��2�T�j�Ua�C͸+5�"��vq�ٶ)9�i�<��vQ�Qc�ÌXj���d��C�J�m����$|�2l����-�z�W]����#p�{���*�GR�� 8�tѮǹ�E6e�wk\��1j
jV%Jxsj��xh�u�fFUA��kF-��I-�kRỬ���N��m��k��i��
�m�
p6�vaEbMoڌ������n���4�D�ā��-k�?��ya#K^��h��g#0��n0%
��=�����iyBa�Ol!D�Zt�D�l9Yaḓ���Ex7`���^ܰSa£߶F�Y35Zv�5�%t�J-Q���*�ː���:�����=݈�ss/Xuz�V�������E���+�?{`�ՏX�'�|]iVh9��+M�ˡ��$�2�D)"�M�N�"r��P6/+NE��;�TkkM�{�RקN��XNAb�n+�ɦQ�u�͠�
�3u�`|b�nͽ��N�j�	,ӫ#3(��v��5[sq��.;��U՜C���BC�To[���nbd�h��6Ax�G�$�jX^^��dyR-ރ�[Hk��P��:0Zʱg�V�I5#��c�;ƫ5|U����3��>!7�jL��u� oTz�=U�����s���
���\����v4-NvT�z�p�\���ö������/�8��VgR6�t��Χ��1��� ���#�������[{�����::ɦ�w��K1v?���ϒ0�*đ���n}���moM�	���-Q�v7#S�;�elƎ�;k_4�" h絋�[gj��SC��eG�����nl�r���]u�P�X�nda���=�L��xks:jZ�!�� �c�Y�����p��p�\6@w�v]'H��K�[��oY�I�����Hu5��zqj�j{�%I��7��>v��kv��9��w���:�v��c�m�TֲL|,�w���foC.�+^I�(�GM.���|)�`]�X��>z>�}�����o�8��:�[��m	����if�;�3hwd�M.0�WC52b�s�nd|�4�]ܥ���2��BL�V��Y=��!31�9�]�M���Ʈ��c��b��;&㵓x�@��PnK,����Gn(��ŷQMu����X�գ����J4�?���;f	��7����Φ�i�[a���soh^
ٮ�]��}��pnM��Va��V�i%�S��M��)9/:Y�!<�Gn.��X���Y��Jj��5�� v�g(�б&.�q�\C�
�+*��cT�v.��\4�4�����{CD82�m^�8K� �i�J�7��C�9��գ�֚���P���V	�Kw���/R��d]��$�ЫQ���.Zv()N�L������F(E��*.a4U�@yd�:�+���
��\���R�2�4f��+��ԇ,0��[���T��,N&�J:��s��sT77�&��N���]ʔ�+Op�
��Ҋ.��B�!W{�kf���U>{��U����T��+�o��M�j�$^���ȯ�TG0M�>}���\�@�`6x��t�8�]�Y)��	��Sf)����=:-�Bӽ��l�|1���%��tQm�Γ�e���l9�ge؝��{��oUuͅ+B�37���࠽��X���yּW0c״�6�$4�Q����㡨եh��Է��v#��
+/��Jqu����a
�M��+S�!�J��9���.�(.�`Ǻ��9���w�&� 1��/��$��-[��ltɀ!(l���h���;�Վ�D�;Lt*��������lV�0Xٸ8��>J��Ab;&+���
I�wgMQ�^���߷��W ����u).�Hoiy����ofQ$;̱n�K��`�<��F��v�^�xDVE�f�u�ϥ�Vi*g�>J`d%9�Ym��!��QH)��m;1���X0<���L��,�)�J����z>ew�<`��$�IW`�Ź�	�X$l�>��`��H���3n�O�Z~������֓ڻ˺��I �l����_i�����n(�J7C)-Iǆu���w ,P��%��Wv�,��S*#{�L"s�ɢ��:�E؇Q3��R�(�eJ�фɗ�´Z4d�oJy6��B.IWU� ��"��؅���lX�}� ����]�mܰ�U��s��O��҈k�2�玘Y|~��5����,��3�.�]f�;8�ѯ8�.#���z)X�=eI*Ҿ��ݑ�e��Cz�k
�ۺf�m[�2	�ԙp0�ZE�P7݅�yvE�"��;����\��G�,�]��ڹ���[����m�,�:�7ʓ�z��՘�Z(��ñqO�HS {��T\UA5�]���I�K����xf*����e i�f��^2*TW�T��p�:;5����,��-�u�񂡲Q̼�*�m�ҧd甯��\Y޽54�\C�X.
7�q�m�J��9@�:��4��*h��\���:�L��6�։J�R��!p5�˦Y����rRh��6+���U��X+�N�L�O�W\Vs�Ukux�9�!���}P�	�-P�&
�W6�e�0��e��Z�P��)ԜJ��NY�
�^yB���FI�\�aQ�[��勯i�����9��%aY�M�$��0���],\���g�0ѭ������O�;�/Zî�n�6Q�ZsmVڮ��^wZ�Y�ŬE%���#]#�'eຖ�k���>���-�[9wJRōҰ���u*�r��'4c�j�m`i����T�H���=�8�[C&�u�j�7J���n�6�e�N�&��ɩ.��F�y� .�(�(r�ʳ{ۗ��zZ�YgL4�uyx� �_b����U�͋��۠�j����F�4h��e�]�/�<�:�;n>vdЫU�쮶+Ԇ�ܝ���DP�}׳U���pf��6�5��Dp�i����p՚������	R�H�[T\T�G4��<�-r��b��n��r�o����V���#�GS�8�M�N���O]8��J��(�ˬuԄ�5�X�2��p��ZM�\�kG �Y���;��I<6��zѫuwM�6]�\2��gw���mrw�v'�]j[�)��ԕ�`T�ݍ(�Fa���i-6�H.⬸��:z�(`*4;fe_mpgZ�>`�l�����	��F!E�j#����i�|��U=�e^c{&�3�Ho:Ƌ-��¯k��i��!%�gp��+"Zy%z�%L+���8�q�,�Z�kGa !=B��@��c��u��+7+��g�S᡼Ӏ7r�ݷ����v������T��-r̄-�x[̫w�������}{�ޝx'�I$VE��6KI@����D�����g���J�r)�+�Lf��y,��S7�6�{�����(o ��Eeӎ`SP�a&�HA�W�Dh���v4��t%Ԗ.F����y1��Eʸ9.Nٷ��c�����wY�\������I��:�/�j��{���:�����QU�T`�cU�E�$Y�EE@X(�E�ATR���,"�" *�dEQR��EDQ"��1�A����w��Ӊ~�g�y��8�W���Z��NZ�����q����x��t��V�S�-�D�v�;�;�~�|�_p��r{��S�j��S�Rg����9���Ru3#�@
����V��������u�5�Q�<(�<pZ*�e8?����>}Wr�*�ǞN�q��|�8�a���2���\�7dk[B�o�lѺ��p5wݏ�JI��v�J�Ձ]��|�;�	�"��� ^&�1Bs������a������4C�r��x⎭�ٮU��bQ�����s������pˇ=��'��7C�}�Is�i�p}8޵��v��9,��<o_�%��Z���('j\4���i��ܮ�b��@z����}��G�7����ZR��9��pmZ#��?	�+�#�W��c5[9��E;�S}�3��v���o{�3�5��m*�{��-ܧ��9���{��޻1�<���1�F�I.�3��xا�ǘ��OdF{�FiVިc˴8�`[�-���Pӟo{�� @�Y&����}�ء�������O9=�*��J�tF�٦�{#Q	/7�-f\��W���LÓ ��z�ᒒ�����u�v��[�,�����e~Z���{��VО��H�`�f��e�W��Ϯ�o�LY�)��Ҋ4�I�m�=�+[�C�13}֕RKu�vF�3x�Pmꤷ�Yx��"}�sQ���~���6��
V+(䙍������k��K'�[���em����u�4���&�Ͷ��扄S}5Eo�A���*t�w^�;/�^�NC�X�6�Z��F�0*܆�=q����x2o��z��Z¿7����^����>��f�<�bK	�y�����C�5�f3%�~���N�P{l�[�c�3�����m?X�=��l^���W\��.�"��u�R)���Ȭ��t���e]-�/-xJ�� p����N�{������fc�(��{�7�g�Q�)�n}C-NԬf�L{��hx����³=�n-:��LK�̂��;��٧U��oe,eWI�`F�H[�ڒ�D�B��������h-�߆G�N~�n��yϬ�v�p��0���9E�y,lo�q�!;zV��i�����Gq������RQOu���4>nhL�o*�վ9��2�� ��|�(��)b�=�t4���YٴzU�1���@��3,�V[PF�5V��3��U�z~��o�A=g���z��Jp���-(���+�/i	p�w��6�6��ٵ�4#2�ovA�,�1+�n��y�m����u3IdEƪ+�n��%1��5ڪD�(��t��z:�ypP���M�^��/�I��W`V_��W�WUX�UH�QX����*��b�V1Tb1R0PR(,`�"

�VAH

�b(�"�E�R(��� ���b�����Ƞ��QUH�ȱH������/�ۦ�v^<z�G_�W�W��eG�}4<G���T�8�P�u�y>�C�����9f���r{�����K���^��S��5���x�ЂvV���L��ٮJ;��O$}�݌�nt^�ko[��DK!h��Y�����w�`NY�+�Һ����wr�o�F�+7q�`qz�׋�Nڿu��+��qD�Ϫ��wm����U5k�+�I�M/'��S藛�3q��2��xɘhmLX�h�]51\����KB����m�|�aO1�W=E#�87�������=���x�/qRCCIܒ�K�F�>Y��ڶ��d��!Ġ��
߽�ܑh�[1�3 ���n�esZ�:Q�q
���1t��WjR��%E��	o��^{���g٫"Bhu�փ����-�L{���S���Vq G��<���6�	������7�omiq��)��멇v�m�8�����������o0���O2�a-kAW�@Ϣ k� ��j���`�4_��ے���G�/�yq�~���8%��_�Bo%^~�%;��oje#/�k4��W�-s��%����B���o���K�G�^�A&U�I)����۠Gae�D�Ign9<��I� �t��=Ȝ9�;8f�
�f��<���e�ƶ��m�V�K'ݶ���Z>�0�k�J�Ǎ���F��hvsܭ��^��Mz#�+�]���d�=JT����d�k3���T����?_�W�5�;;�:=N�kg����C�z�Ƥ]����>���B����9�xǺ;��/��Z��`��nL��T�l����i9\�'aT�&Y��9�L�ҋ�̈́���/L<!
�I��x��8�-����q���Y�q#a���w�=Dua�|<����v�|�]qF$�<�{J��j�6��ӊ��b��R���N�`���6s�.��:[.B��9~^U"]�,�:�'S���n�CR��en4����]W��ilV����� �5��+A~y�&'��E����|����_m������U��S�Yh�;!}6�e���� O���A��tA�����Y���QY��A,`�[a��]85�y���b˜�V��y��Cw{#6t��id9���Y��r.˗{t#K"µ��I��sj�!�/�e��Bо�lX�ܽ`����ݳ��>��*C{:{i�6�t o<�ԣ��Ĥj.�����U��w��Ѱz�o;Y6�q"+:����#���+��m�������$�{�r�s,�ؕj���u2�wʇ�1�A�w$� �m�m:܏Q�.�M�1[�T��<j��VP�͜��|��_Yp��`1�,PU��`����H�H�QH�D��`(�1EEEQUH���PDF'�j�w��[�/��l��h��ߘ6���U(�ex1��%�s��ٱ�z��o�1z�G��E���X�xu��N���?0=�Ά�����v ���%��Ys\�1���U
`d�W��J�ӝ����rr_i�^�N�l�U�/w��{�O��+Jw��;���!�鈒�y7��o���V�Kf'Z3����e�6<8�ҧ�c1���ږ�kTޑw\��ީu%�Zʩ*�-�H�%�z���,{�/��R�`u�=/L�1;}�1S�4S�ٝ�f��G����:Ϸ�Z���<�0l��q��Z=�������Ѱ�a�:$�C0V��Ż���ǖ܃G��&;s����g�y!������4
��"k�����d1�:� z�nU��]n��$V���y׺gtF��s��{�e��!�ˏ���JHӐ�s�o��]E͡��y��S}w^��M������13
��7�"'3N�OWw]C�n���7b�Ϟg��+f��%�
��07rx���)���^!���u�#���ns[�����cWt�MpM�:cMX��(��(\Uȏ���{jm�C��V<�Ĉ8%	~��A6���kK��Y���B:���.Y�Q|X�e�a���Z�k��L��U���92���P��,�[[�J�פ�K���1�q3%�*�+�7�����q��}���I�u��iu�;�e&Y��Y���7���h�R�8�t�ڂ�k�Ļ!��Z�.�[VL�@�,:��9D�xs]�3XCC,8��i�mǝ�su,ًHVs�rغYÓT]%����r�5ʜp�U$���|�lg��gp��T�<�×�DcA�άB��v��ܩ�Y%�gw�a�fP�h���mQGjS(έ̷�2�l�dq�M�Y{�ŭ��'�q�.���[�ͪWh�Y0�2۷w|^N�S��Hi�Ch�;���8�3�.��R�6��v�:�L):�!�S��W+Hxr� a2�C���<�>�ª���pT�z���'.��͢c���S�4�Odj1*�z��;z��ad�l���[m�(�L�+����x�׬����ջxa%^����hj��Y��Nf��2�S��кAL!d�ֆ�w��&�2�!}[-��&�I&�gU.�CL2���[쮪n�e�L�(��*��V��s|�0i�ޮ��.	7���R�5(�NH�y�1j�e��JK�����ίm��H�f-�j��JAd�C)�:�Z�ͪm�h�0γ7���4��պ� ��K!��<��hFN&\2��V�;Ѽ_�!��,t˸�]���@Ђ�gwF��Y�t��B�菿?r�?3�b�^T��+5���Gv��VB�C =M�("���wMe�eC@�f�EV�t��nKw��B��}�F��:{�	v*�Il��^|Ř-3�R�f`�1"��Q(�w�-d;9p��eȖ�]S0m��1�b]:9[�٘Fpczf���o7���A��/���R��i�k�oB�d�:;ln�D��4�+IΝ��r�óN��E��+���;��`C���\�2誑��\��9�[2)sM�i�X�fwSv�GݡK�S$�󲚹M�+U�Y�[��fQu����U"�"�E�(�� ��*1"���`��AUb�E�d��*1E�Ŋ�AH"�u"�O{{s���c�^or��Vgr����`��S�����jo0����j��t0���r��M��c����Ifa�Bɴ�1k�:�3=��Jc|�X��d��aIcNqsSi�a0�S�;j�N�f���M��)2ͼM�yE�֩�_��U}�bС_S�._z\�e=Xr��� O�ӶJԯѡ9���1�/�/��}wӧ9�'XS:ɴX(�-�^���n��2�B�Zir��S�,^��t�a�e�E3��7�`q�CZ�.\��R��{�M7i4��-4�����Rm!�i��Mo8)��M��5T(aM^���ɦ]����%^�Z巾rδ�=vK%4Y๹f���1�2β̤�]��lj�ͤ3T]�ƨ��c�)ƒ)���9Ǘ���N��L�V��Ũ㴲gXN���,n��\%����SII��R%2�
A*�����
AAH�������[0;j �l���H)�) �.�AH) �����12��`u���R�) ���L�����X��t�˞*K$aI�&;E�
AAH�wy�I���R
AH) ��R
Ad�) ��l�R
a:���
C�)�=�d��2V�f��$q��
AAH���R
AB�RAH)"�Y,�K RAAg�RA�����!S�.��1�s�EZ65�9l�x�u��������Z�Si0�$<�Z���) ��
H) ���R
AH) �3TAH,��u�;�	%2�T��S{�,�P�h�H) ���R
Aaf�R
i���yl�ƈ] ��فI	I �`RAAH�M�
AH) ���Xi(	m��}Ԅ� q��!4�K��Y!�P@/�k�	Ԃ�R&M�
Ad�) ��B�
AH) �̔�Xm�$�$���X�`RAH) �3U-$Zl������AH) ���R
aI���z�%�
A���βRAH)H�R
Av����`RAId) �(i ���P�w����H,��K$��kR
q�0���P�JH)	)�d��ͲRAH) ��3�@�AH)&P�����AH)t
H(i%$K2�
Ad�) �����P9���
���c�=*n`�ޘ�Pҫ	d��y;'<�7W��y1�E�r*����
Jz�g���q&#/A�ͳ�̺�B2_:�K>��(��X�;ڛt�M�/nW-k��K8M���(ͮ�4�3�f�/�4��M���^d@�.�7eӉlf۵J`q�C(e;��5i�T�[�S��l�9O���^�����P���Jr�&d�w��� K��m�K3�Y��8�֞jՅ��	��g^ϋ�Qd�Q�,�9��m�)��
=���Ү��)�i7|cZ��&�S2ɶN�{��oSNܥ�2�����)�Կju��E��7��d�J�u�8��/�i�B����{�݂����2>�q_�/6m���w��$�A�q@x`�G,�7ڞ*���ݪW�!Bi�e��9Z��)vku+5%3�B��w���
JM�S�kz�7nj]�.�1�B�ĝ�m����Y�] �{RXի]��N��]��k�{ѫPU��R�!�c���0�t�C.Sl)�`�B�Yx�f��c��C-�׶��y���qˮ����N����u��z�B�k�s�i�a,�{s�_��t��ƪg-��,��+����ت��i�z���,D�V-{�)��4n�@Xa7ww���;ba6�/�]I��6�	4����%N!�e��ff�kW�l�0�I��9���Ì�E�FL}�Y�B�ZQghА�w;W���X�����}WT�O��?$�RN_�Y�ԺS4��Գ��,M �Sl�^�0έ�a�=��]%����Ũ�,��m�<n��Zac�f���f��E!sZ��1�|!w,��Ό�3M�Mꥱ]M��E;�sU�#0뤿jV(��ͷ{`s�[��Y���T�ɪ+Ӓ9���*������|�#(}L�m����Q*�d���D�Y�c=��cQ�+�ʹ�y/{>oٍ�k��&Bf=�#�fd�X==� ��u�m�!Rc����R� 7Ʋ��Q�i^J�е�&����z^��z�Z�ˡ�Kn�!��x��nea4�MB����A�X�Q^L����ړw��($�{$)�pp:q �'�#�\����[�B�	�][��6�9����b���=��+9#mTF1��莗R�_6��sE�;�NV�ݖ�Y	�=c�I^�ͪ��J�
�"xp���G�CZR��6�<���;�W%N.�b�wrg^�,��M(v3���$�Խ��J����ʎ+��tdl�j�%�^<]u
�5�d-*ILQJJiP@i*E�%*�F#E))�i�cQT��(*�P��JQ�Z)b�(K����3����)p@�J�]
1I���" "�O����C�\�����(�\W�6&�O,�o���q8w�{�g{���3��D��
�ťD��k�#�d�SsK8Ox���?*)��;��{�F]fC�r��٭2�s�x�\~DD}��%)������eX��G׬)(=+4mi��5��˰�3�$�yS%��Q�>��cD��>�8�w;w�i
�'�ҋ�C1	�dfC=��gq�=K(c���C�t��H+r�m��}���N�xFN5�5�U�V5g2�5�l�s\���E���@=d5�%n�=��@\�)<m�dЍa�<��r�ʳwu�'�8	�}cG~3n��x�������zq��G�}��w����+���f�Ҩ<=R���Q�_���ssMzٿ3<�/9�g(�jZ�/0W+�m�Ŏg �S�*`��!̜u��[@�)�x��e���W.�;3:;�#��xiĞ����ﾰ�޺�����MȜ������`�1Z/���7�����'��sΤ�1Fk[44_c�.5���:�hnQ��̢���s�o�Of�4����0��{�9�Vˀ̀�r�|��O��}�V�0�ќǂnp�2��U�7�������_�?���E> 5�~$kq~i�����/��~;�[����o0
K}:�]�La<���(���ˍ�ʹ��K{�S��}I�L�������-PW�7k�!��q�`8kt0��=�a|��gN�P3�� ݽm.�+Vsb �/|�d����%���T� 9�hM̞�ޛ]��w��ND�e��DFQ�d�Dͺ�S>ۇ+F3{u"c���G1#��\����o����y�����}��t��O�M�K#��rK���~���>���[��mA�����VIm�z��������D �����c�W<�~�]��A���r����+U�w�P���OY'�7��^1�^�0�cy
�ە0��8`������$�ظ����VgܵyQ.�1�ߙUmnכ�����DD@7阞�1�I����d���}�T�mQ�ޛ�٦���G�{�}���)Z�h����<�~��y�c�oN�����8�$X���u�Y!��!
S;�q0w.�_^��1=�u
�E�����eV�ޓ��aQ�Ƈb
<4��k �DNkYHA��*�k�s��.s��.�;��ԾF�̒C��],�B�ue'�.�cg�7B������5�ΰ:e*�B�V�n]^���*�6���V�@� �
Y���V�Lj��@���K�CVd*+�@.a�|�u�-��
���pe�c���x�}�avk&׹Fb8���� v^���YS#�B�,�6�It+�iC8<�EnQ#��ET�3L�y���#�l��8�3e
�AG�,���n���H�AUM5
i)�)*��ET�Qj���� �F������QB��(F�Q(����i� �(����S��~]۹٫�7�G�}��g�<=�U�hE)�^�Q�Ԕ�V�.��C�n�/��#[[���'����J�>[��s�nVY��Y����\9 �>���TiE�$͙��R�4΄�qE9O�}����։��6� 
�/�Y�=��6cO5(fs ��f�T���1ЄF_����yQٹ�3�8L����[�z�<���)]%`�]�1=���#\PB<r���rd�)i�������ڿ}�q'�wM}y_���d-�5l��;�؎�kث�݁��N�����m��h�y�y���t��G8y���r�<=�����3�ӽ�֕)Ƨv�3fr����\LD�����������R��ˮ��/�LV��ﵵ�V�O����i]/n�D=����V<y7W��D]����m�
��w�&�����Z���i�_X��S�U��E�d�����:��n.i��-��������v~f���<�\~WfW�G��V�2�3�HaZۅ�ô6���:]s�a�����m�'_]m6u`0>껡�m�M�Fiʝ�}�8j��u���N�rrb�}?Ͼ������5�ᙧ+(��h:��j���b�uD�����a,��YF����������м�@��B�@�bg�0���y3�]F�8ՙ���D��
���������wYy���߫�mB��36�dP~ҳ���s�[�<I9�^ɫlvj*-6�ټ�h���������{ڬ^����$�5ӳ���gr���pQ7���N��Ӯ2��[x�~*�Oy&z�T�Cr�f�1�8f�ۘ]G(O�Y��"� wo�Q-;i�k�ŷ�j&�ɜ<���v��v-4���	��eɆ���~Ӱ��7�ˍ����j�j��G&�
-�"IW����v���?,ڟ���*�_>ʰfy��<�Vi�t+0���!��F��v6<��]N@�Wb��jd�$��$�Г�Wa�'�&l���X��2�'��)�dWE])��Jܶ�͆��P9Y�����e���5ۋu�a�������ˆ�'rX�����}���z�G3�=�I;�8yi�w�Q�M(̓�81��7 �xa>ǳ��m�zvЅC��uͼ�z0æ9�jI�B���ja���#޷´]��4!��M;[��b�kU�CKmk���� `��0�g��b���'���*�Xn�J�S yh��n��"Y�
�N���(*�*J �޻��uc8�M��Wl�n��q9u���z�z�9��oJ��3�8E����xy�t�<�����0�ݸ9C�S)3��֢��;ݶZ��pK̃4Q����R_es<�`R�ֶKGQ%8AdNY[C6璹���J�Vγf��Ji))��T�M%P�,��,J��UE(����eF�1H��X�U ��S�TEU�L���*"-"�T�J�
*���
&�Z1�o\�9�A[��qvg���Dx�J��t�����)�C�uו��O��w2_��-;d�B2\]ݡP a0�uw�)�h���y�7�/z\�I�M���4e���8��3 @�YzC�6�H�x��܏���ˊ$S���h�^K��F�-&;}��}H.B�摣`��J+�gh�H�n�����k�`�L��=Z*8�N��v��8Poh��)��x	�8���l-�=Wj�{���P���QY�V3N8�&�v�`�'�~�D�¡&���I)�  ��|mn�>h�m���oX�.em���֓�]�<�O]��`���v�ƴ"f�Ĳ�g�tAv�f���5�xC߾j�c���1v��i�4&�S�؉�K�hl:�3,�.�MZ�&Y��[˴-���<��oB_��R�}��[�c]֜Q`p�g^E�L=u�E�[Rz9��U��L2��+Ɵ��O����SKcM3)͚Xm'�5��{����޽�ȱ��ۧ�x�/[e3���g�h����gr��u��o]/5��RNW���*�^B*c"�E��q�������'��{z�%m�>��������½��Ϸ�Q~�Oz��J(Ӑ潿��/�r�T�/eXg%�q+�_9w޹��kx9,R�"9���\���B\�բ��䦁�4x�!%��p7E�e���u7J��V�<��z�w�t���t�{1<*��)��K�Oj��-M�ٌ�[$���z�͋]��tN��7�"�v�ZPx�e溛�xd[q��~���ݭ��;�vg��ս�ǹ@7`���*��z��K��hn*�u Tq��SL�K�`��G��m�5[�{
�tdkǯ6ۑS�g��x4��D�o�-�lj�v�X�ft9�l��Z��V��D,D]BS!A�E�?�R�׶�����ն�L��ɁՓ�s��:8�C6]f�o�UKH�>�.p��C��j}�����БD��{�Y�Ii�1�j�j��>ͻ��Dfȓc�1�y�2�_u�bN1Ǣ�2�oX�^���y�b/��7�M�g\Ub]v+�� n�����,e�:���M{Xn�d!U���CZU[=M�L�yQ�W�w��Gb��
�Xv6�\b��ctT!1��P��M��+�ӆ�Zش�U��z�1�)ff��pK����-�c��@����
�O�.�W���c����,r�K��8���yѝc�D5��Yڵ�R����[�X�c���M۴�I}%��{FX�6]��S��� ���hwOe��d��:�.�h՞��7��*u�ї�5��kD�����D'�i��u f�'8Y��7��/�
sm4�+��w})}T���^=}+�X�$%]d�kRڈ�5ǭ�j�}���+���c�\� ƞJJ��X�2�<6=�:��Z��kl�6 r<ި�܊�	6��^��o$J�&�Eq	�\�V�|�Gݘu�K�m��UEUAQ`�X��Eb�QAf�Lc ,E"0X( �E���c^��9#q���}��b'�p��7�%��y[jv��5u���?-��C��s�ұ�r�,Y�]̪,�ѓw�gÌc�3�K�"w(�՜��:x��X۳��n�������{Dӛ�0W9�,�.�|��zPr�6�E����@z�]�-u+'����g&��<�����u||x�[�,��������R�B�7[�u� �C~Z���y�k�7�<6Pdx�Ɨ�κ��L��<�����1}�I��w�ׂƎc����f�:�l�d���
n�{۾�D{����X���W�����cD���ft�v��x9\u��$��~ׇ{�8�٭��L��+-j�~wܢ����C��4�_d��􃝙�1.���Y��r�-��E8eX��z��ab�e��@�.K���f�7��/	�5����K�\�UDt�nGe�}1Yb���
�֩n�m&����PASư�Y0%��iL�87f �����q��1�:�\�O�7�%1��7�2��+�B^�܁���Y�Y\�Y�h��z�m/@�G��u{�9w 9=�տOxfo����������ی����t5}A<wN��t�1)�pv_;���ק0:�F���ڄe�}*E��Yw!�C���>O2y��ԱX��B���L
l�����,�˧����q%�b1��|{;����7z.昏v�%�m,&qWYr߮�݇�"�v6B&X����kw�������E~!z�d2(K�6@����X:���ŧ+�].���{6B22i�o�j���v_� �#}��}�߹�f/�_k�w]h�T�Q|���LS�8hݖ(���8�?q�yOOt�G�	��aM�o��/C�|���H\e�J������nu�P���We��ݤ��be�~n�R�1�2P}@x���|9�-]�
?@y�à�qw�#9�1+���rDvM�v���|]JIj���a�7|�cG�T5z��ɓd��yO�Q���;�e�B�U���)]0yy�D����cu��XAS<��;$|}�����A��8�S{�Y��p�9A�c��2��\o�ט���J:�Ǚ�2=�k&�FNW�u���y��iw��	)�3s��I��̣�ס'�&��_���A�lz����"��H�ҩ\�l�3��1��'Z�u�l�OE��"�VR|��p�J���	X�[�.݁�!�
'�/<u�WV.�=�2�o,fvc�ڰ)L�ۚ6�6��i�C'"ܙ��t���pnnMgj%7*��[]�0X�̵���vO"TV��S��껊f���13�����%]٧FB��Ji���z�����G'h�� 6��Et#z��Y��\�n�9V�u�W���{���#�K�7ԩs�*�]p��H�p��w�D�l��P]�z��i�[��R�:�"��:��
Ȣ��|9��>�{�%r��btY˥��]3+	�f]�|�_���l�;ˋ�[�
�PQ`���
"b�2
���*1b��TEH�EV(*�1UUX�
��QEQ���w��tp�9Z�mƶ��ksF}p�G;���gv�k�j���{Dx�җv'#f�Z*�xVD���Y39��V�3��ڰ�>l5�OA�I~+b���2O6����SJ�<�5�b�:����L�+0���hj����(�%�o�����G9ة1y�(���(2�m(]�N���}K�3G�*_-%�R�)\��� "{�;�,�����+����j�@) 6V4�.�v�P�X���U�7�"m��ZW+Sf��IΑ�\��y�/��\�j�4�^k�uq��1���5�I��6r@��a₷	�&p<��:�n����~"r��oT&����up�BͶ�#Ӹڻ%/MZ���*�J�])nB�eŸ���bp���G��<w�_i��oχ#�6�y雇WQo��׍���a�z��l�q�3��G�+��<�J�0��+T�	}v�Lȡ�ܭ����e���]N��%�i� ���ű�����؝bYe�����v؜3��h����4��t�Y���5���U���#���K{Nh3�tS"�|5�͙�C3�+d�D�#C����<���;+��J$ֳ�0:�����fG7+{/��v޾R���t��v3�;�{�>�׊l��77.��s��]fm��Q�ˢ]����yx(��᎙��LWx�q����xV`ieaO�g�yqVH��\��n#"����^��	�4pW��8_y���O��ms|�f������.ʗg<Is�ˢp���N�f�zX�=�*�/0򽚏*:����c�K;*�3��C�*�^6�mE�C���M0FS��J�,@��?�;a�\/�Z07�
���Ô�Y*{[���t��̻��	{�������ꓲL8�F�m�Ӵ˕B{L%M}t�O�m%)i[od��]^Y�v�M48�3����E�m�׷���`�=ȫ����rr��Y�^	7)=�7���m�:w�ѿF�K�A.޽W�8oX�=�߹���^�B�ۻGw3�Wwd	$�'��d_w>6]]ȷ�C��W��F��O�5AԖ�0�I[ܯN��Ŋ���7��*�Fw����t����>A�tk�C�e�*&����8�DMT�(I|q]g@'+
֟a�@�u�oUM��)�F�Vw�f?zO�U0~8� u�w���ko�dF[���x�n7��n�(��md���/�7�9�����7|�`u�`���)[���m� @_N�2��	�>s����E�=�b�B�)h�e�AI)�Z��v.�f�GW�N��z��d=o�=x���97$��*�k�if�L0b�s�R3}]�-d�%fM6i ��(�u�vr�#)(�hs�6abw�!U��;���^Z�[�pd��oLF�vc�1J���NL�]�oK\mHfh�U�;�6g1�;�Z�+�p��ܦbt֧M�θ�AH�=S�
(|A�,X","#"$X�`���TTH��Q*�X"*�������E���"���UMoz{�g���a�M�̗�R�fxn��ҷW:�Ӆ3�	��`��g��#� U��~.��4���h��Ѻ�6����V]�	�<{&���;w�A�1�:a������kz�WV��Z�j5�4M!@��K�h��f���R��U���{��!Ƀ}V0L�\@�l��ܮ�;9H�Ӱ�+ME���]i;}@�{r��w�@̣Af�~��9�k�;W�D�]���ݮ���$:��4�	Lvv��E$1��"��X���jd� Gni�7�D-���2m�]�;�w���
�B^�(ރq��I����^d��}�Ƅ��WJU�%�a����^�9H��C$iN̯X]���͋�>��~�����O3e��<��WQN�|��O�cL�E�f���іQ��3�2��]��_���3&:Z/�Wee~��q�,�0��Z��,�fܻ���Q��1OR��o/i٦�{��k��{}Ձ\�Z�y��Z=��ה.�M;�U;��ځ$��> ��2�=�(�Vxm�O.e��j�\��{����-�gS��N����n�i��1��c����M�U�Oa4�4]����-Iu���=���tEy��ݟ]_�z}����HT�32���3J�ήƺ���y�R�7um����[J����� ��Ѩ��;�0RnyI�n]_�ݥ^��c&2�{�@1��;�-S_e��I���J��U�ߨg�qH8&&�w��h�c��/3��Gvg��F�!��j11�INa���۶��&���p?1����g��Oq�m�t������Ϯ�Ⱥ��&���IY=�Wc� ��h��o��@�oR�-�L'�OJg$�5MRYc׹B�z��79t�-�R�f��NN@֕��W�@<��K��:��~�w�v�꩟h�bB֮�]�-��w�Dr��F��95��P�rbI�f��E;W�j�?{��|7�r?��-;�-r�/-s*%%�;S�`ͷ��g��>����_��l����<�rnm�T���Q�n����_��U�"c���=���:���
������~A��~I�QM*�*�@��B�w�BI� BI!��E�~��`�����jQl?��\�|��6�.�󵙦�`BI!�(2��d��mY�$�.%r��'�		$��v��N�q�Z��Ϟ|~�<�-�ҭ3c�q�퀅�ݤ���v��l,g�!������Ƌ��H�N��s����!A�>��H~`��HI$?��A"¤���?����d>���I��a?�m��h{��0��(�HBI!���T�܂�r�~��Oo�,�KJ1��t�;��+6@?�{W�ّ��d�}'���#頸]��I���TI$]����s�̓��V�BI!pauXN`�X�yV�k|u�A���ˡ�W<�I$<�I��z�I랇���������<���C��C����I��F?(|�p���W�������H|c7O�=s�O�{�a�FW�>xjnJ�$�����>��Y8C���>�x��I�3��>��4zϔI$=P����E��>����}y�ȒI$����̄$��򟴑=���'͠�=��?���pوQ	�`�ϝ�I$���벨ǠZXP��f���@ �LT�4 ��}�9"c�TO�́��KI����h~:.b��[����C����>o@>�{`BI!�|d?�!\�������������=��/8{$�	�|}'��}��e�g����>~��C��[�{#p����I$=�̿��!�!>�TI$=�X/�%���I����d�'O ��=I��0 �O�{��Bĳ�^����s?XC��^�g�5Ff��W�� BI!�=K�����o*�g��R�ρ�!�uA�c݊��0 ��P�!��$��Hh�~����z�������=�d��H{���z���{��L�09
�bLj�>5|�E$� ��P;!�Q����H�
	:mp`