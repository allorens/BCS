BZh91AY&SY�)	��t߀`q���#� ����b%�                                         @QU"X �*����� �@@ �  � (�
      P   �  U    R (��AH��)R��E
� U"DQ JT��*!R�J�T��T)%U*�*�I$��P�Q%(���@�I  h�*��U*�RUT� x}v8�\����
��4R]�",��*� �*�h$7[�R����W�A�O�   4o�}�Prt ;䪽��O��y�ж�7��H��U"���m�2;cl��)N�{��c�` ���T� �<� {�W�� :�� ('Δ ��U�IR��Ju�+� �=���`�� ��r .窪U�l=W��:���cް z��yR� ��z��  ��@`}� � ��"Q< 	=�=���N���� �t�T` ��=�7����`;��� ( �R����*����DP������@�`G �rP�`� 8�9��� e�� 6� �� R@W�R � �ٻ� {�%� ���<�� {@�V "9 wX�� � u
�@w�I  ��R�����EJ�H���G���<A�� �n���EU0�s n�C ,褌 Y���    �|�  >� l :n�%X H�s�9��C� �qF c��(w`�� �  Ϣ�  >��%QJQ*�� b!C� ��#�� �J�`#�v ;�!� c�����݁ʠU (G�%   ����	@:�K�� d�7` f���HUp�� �C; >         �� R�  4    �0IIU@ѣCF���h OF�I�T��   h4�*H�I@  L  d`��JQ"JM0&�L 14�� ��h��	�lI��hM��}>߾�����?H<�?��3��:���8�����"
+�N5��DQ^T@T�����k�����( ������C�G�?���}O�:?���s�~�}U?�A��6I$�4(�����#�d�D@w���#ȏ��@+ P��
�@+D� �
ŒP
�+@�Q
�+ @�DZ�#V�AU�@�@
�U� 
�+@�@�DX�+��E+P� J�@+�@+ +++�F5��V#X-b5��X5�� V+X�`��VX%`��V!X%b��VX%`��VV	X�b��V)X%`��V!X�b�V!X�cX��V)X%`��VX�`��V1��#X�b��V)X�b��V��X�b��V	X�b���1�k���k��F���k�R�Ĭ�k��J�+��J�(�+�R��+�R�J�+�
�k�F���k�J�#�X�
�
�k +��k++��J�+���J�+�R�J�+��#�J�k��J�+��J�(HA+��J�k�R�J�+��R�J�+�F��k��+0�+�F��k�F�k1J�+��J�k�R�Ō
�k���k��Ō
�+��J�k��J�0°�k��B�J�+�J���+�B�
�+��
�+ ��J��#��J�+�B�J�+�B��X�+ �B�
�+�B�
�+��
��H�+��#�AkF�+�Q�E���Ak�Ak�DE�d�U�@+V�k@�Z��Z��B0+F�k V�EkF�DE���@�Q!V�Tl�[!F�DQ�k�k0k �Tl�����A!�l�J��Q�D�Q��Q�E��TZ�� ���K������N��E���m���x�9��.:^hˌ̩C:� ����ktc�S���� 7g(s��83a��rK.�d��t��r]CQK��5�<�ON������ǔ2����N^�^���9�H�����n�o%EÖ�43�l��3��y�6�QjEDwj��~����N>Fwqe;�P��g���\[H��[{�B���q>�.��4i��:Ww<�M�	=�Ǜj����̕��r׆��0�����S�vgm�t��15�X��)�
����S����$h��{� pf��'F{Y�4k����O/�؄�Y��5�
S�����god��iwA�&�u��G��決���a�h��'�x��[2py���;c9Cm(w��O6��f�4�ͨ��s_1�
r=v�zd����q.����a��"�$��L,�;���k��wc���8q�!ywL٧�1v���g�(��n�Q\��8��z-�m�7������y�9f���4�C��B^kx��Wh�,s{A�1�a�Ljv�L��LABU�`�$&<fϗ$�Y��5�ٛN�je��gs�ݡf���52l��Tw;��L��Joeb$���j�O.��{@�jO靻��tnGRY0v����X� ��D���X�`�2��d#'�mသ�n��a�,xE��F/�(�^Fb֭�׼'�){�Fi�;l��;�teVt�ݢ}Bot��`��ޣ��� 1`5��LrE�F2�3�2P�ݓE*������Wz�g=��%-':��%��0`���0�y�T�B�q�W�}��ya�B>����K׵+.�n��%��˳�y^V�3tY����0�Lz��^\�rHv��!��kpr�+(�+uuO6��n��4�=�\��`I3l8�j��WuET8���G~��Vu�p����5�8AB��]��/<���]oj�������Gt�{pmv�W��;�m<Z"�yG�Bh�7zIT�w�40�|w��tr���CV���3��ƭ�٫flK9�W�U<1�6B�T�k�tDF��#*�ӋU�b�`JN[G`یq�l�)��k ��D� oh�ѫ�
��7K��Ω݊�t����թR�/	~�A.y��V(�f�����T�6�-չ�`v-X�gn���k�(�+��>3'd�2�d��6���.��swn����۷:��ދ9۝t,���5r���7*���n�[��������l&o۰j�P3F�[�_&0�7roK7/5���s�=�xZ#Ow�ы*J5����׮
��9��MN8��#b|L�,����}	�ǐ���L\>[$��'�'z�0f��20�^tPv�����n�z�^�}rsX��L���0ꙥ��b�v��n��uɯ���(���� �;)h^�N]�����=���1����5�8׆��ޝp�����NSgC�5��G�7�u�線�ΰ�IB���|ۤ޲s��w����y��}��FY>�7�E:��h�s�1��{f�ӵ�1�8���\q�^���k��2�W�5�շ�J��W6�<v�4m^�W�"1��e�Wv�v�W��9���;�t���^R=g�>O1ې�̂�*����n�B�V�0����7-�"�H
�ô�(Xt�Ę�nƲ4&�L�Kd!oךV�K��6�Ό�0j��9J\��	%�I�I���w�%ˏc9ٰ�9F��]:^�
�Yl��{��Jz;(���@�l��{D�  ��"'{�1{�\�'NLL�aε�j;����dM��q�m�J�r�^EY�Wma��U yV��n��C~}������z��ͻ����V�mոn�{����,8UΈ,�5�;��DRp	�o��� �3w�	1c�(=98���^d	�lŵ�mXA��s�'��k��P^���?4�ԥ��nQY�k�8;M��q���ǜ.Ŭop���J�:7pb����٢��%����>t�A�C��(�rqt2Щuf�Z��Z������0S��KjI�k��xZ�#��Nr;��ˁ��z5>o����C�	%����yA�;zq����-7M�qW��{�=��ݳ/5y��cyWNЪ���&��m(:�sq�TC헒]����Q�8�Ւ��싻�@-��Zd�ݒ\�����b��Wu �Ax>���wu҉ۯ{���蝦�tװ�KYS��t5��";��w�8v��i����g
�7�P�����3V^���Pwk=�W!��.��W��}�ӓ�;Vu���-Uȁ5oʦL��<9k[�N�550�e�=4n0d[�Fn�8��秧h�]xG7]$C�d��!���扫l`���p�n��5/Ӆ��L�_q܇�t�wl��ea����*�$f�0��B��˹���n㩒�u�.X ��sOv0��i�
�ڭ=�U��.b��r����E�vl���/>c^]�'x]�a�[�l#�{���I������$�aK�.�Y8�[������0�{	d���|f+
��vgj�za��hTvٻz�����kSo�C
�؋<�|�(��N/p��q�;��*��n��&�N��/�]�t�� ����,�ȁg8n��c�t|��[��F.�Oѐ8u�"�N� \��ے�rEfSݨ]ۜ��M��xp!f�"������tl��oM�:��4�����v��n��8��U�,r�N�{�eBd�%]�\v�$����s�M��޹�І�uG:��ヺ��s{�,Ӕ"�v������S�p�,5Z3xLs6���zN{��#��)�Ճ��cB"dJ󽐷��u+�<a 8v�oD�'v�;�����9q��4nք�9qu��B7m�Ơ7�
��%�':'��83q�o��r�Ll�Wf�'Lo=�7Xp|�ll���7�x�Έ=�!Ny�P[�Q����Z[Kޘ��4��06'�c�94a�' X����xˆ��Ѻ�'��owJƠ;t��P�7^���vi�U��r�p�y��7f���v���ӧC	��qr�k���4r���$OGs�;�n��mi�Yu��d�mt�K��QP�Y��o��Zb����y�	'd� En�����{~b����5����[����0]��M;�^�٣9�CrN�h 6�+��n�k����՛�6n�� u��'^��^���!~<��Ǘ��q<q^R�M���P��po�f��n�ոw��sn����ha���<�MV�c�!�6 nú����f��zZ��#��}�7��:7J�_�nB�W0��{�<Z�eY�f��f��E����։�f�x��doz�/w^�mNVǀ&/s�ˁm8�e�����޷#��u��� �^�*��,���ask9��Bv̊���u�"��r1�_�s`w�jÍ��q,��wy��6��L˝;`.j+xe@��|(sQ��͹�8�Жw@��ʒ���iip;�jɺ��{�e:zve�����Bh+����Oq.A�Q��s	��M�h�/�?+��ӿ F�����1�+�V"wkVcvq��D�Yy�!��f����JyZW[�q�"�9u)vظ>��+1��s����C罜m���f��n�����a��숬��0q��ki�b����ys��f���y�9�����,�9�!*��'vL��z8f�rV�
���.�x"$��f(�۝�H![�X�{1�%��4��b�g��b�}�5ݮ>�׼P�xW���%�� ����E��]��ύ"t�H�[[�#��bkO�\'�x�i\��M��;FA���o�*�������9��ply�Z�Wx�1�fr�H쨎WL]�4Tins����)e�	�כ�ϲ�Mm;wG"�c��/M���庖]�����smO����@Uxjǧ)�oL��Mk�M��B�(4v��Ez��E�-��J:0�k(L�__\���(D[��p�x�{�DW6���b�H���Y�ϕ���G�1��K��5�p����p�	�pn�Kr������A*�����hӨ�*��L՚a�կ7vh�6��۬��75f�'͕֌o�����T��5��We�^~��=�	Nh}���7���;@g��Jz�J�WC�U,��j�ޣ�c݄��֑OY� 'Yҁ�ff����m�f�[�aqUDM�.���qc:\۷a]��b}�3N��
VN��哶�2$[p�$j5�PGVFm_wQ�c��h��]ZU�`�\�Q�a�v�e�ľ�t\�b0�� 8b�fuW���GUĕ8χvAҐͩ��F[;f������2A�;�r�ٳ{�;Įy����F6��ڒ�o����;��g�q��{�l��Mk�#�9kZ��WH�E�h�����egn�^Y��l�gf�Ir���͗XA�����7$|Q�_Y���ͻ�hu��&.t8�٠�۝k[7O3
�Ja�u�I�K,A�=��a�R���������� ��#�]$˜�T�]���=�/5�cb��;�p�t¡ʹ*�]���V����^wu�p �3�i�JTuPCM�)�Gi�I���N��۹،�c�-EF���
�䝍(s��8���a��#�@��l�l�@�Z�8T&`��h�^����tN[�
*�k��V�K�뛦���-��xk��]���q���U��oq���R�!� F�;X;�w�-��	ɏn��W���v��k�fvɼN��r�c���˝�{�o!�L�r襔���&:�3v't����4���x#T����H�^$t�oS�9��v� 0�%���ً�k[mgF��j=�؇a��V�s���5m�v��{��AS��vWN_��y����9���mb�	�!�j;�:�m����ՃC0�j�;(�eR�<.�0j��ȋ3HNh)��ygl{��|�s�N��X���}�0=�`r}�0�e ���q��z�v���42�@]�Q۶i�t3��զ1$��T����c��zå(��2Y͜�V@�R��
��[HøՏge甯����;�֛\4�	��m��aؠ�x�&��s��
5���*�["�5�ov1p��8�S��vM����������C0;|8�����s�F�5��R��-w��Vl76��긦�BN�x���
͛@n�u*���3��S�b���LC�����4����;Fo��U�R�(hm�炪�������!Rl��v�����f�ǝ�쫓�$�L53���ŷ�����ȑ4��pN8��h����]C/Ǖ1Z�ۮ�7��1�"�t�
����x2�7t�Xʹq�jOd��}��iV�K�@f/�5��
4��A�3*���UF��9A����;R�.(i�h��k�z�e.Fe�(�{�{f�X�D�d�Ej]����P��B{^���:{QJ��!�\���˻����?Rx�����.M��z�ĉBM�m�&��V5'�(V�$��v�;c�͡u��ql�P�R�I�]GU�HR_u@�>nZ�ź- +���/xu������Mڹ��NwS��,�%�:�Ƹ)���L�䝼sx]Z������F�}�}A{���]���TF��n�����]qs��+;T����,�ʇVqq_q1�ݔ:1�ۿA��w'#�+�m�c����3�vͨw�m�1��4�-I��\s��c�bS8Hsh�܃�y;nM��]��q�@��ں�x.&�+-̀��X;�3�t��LAe�)C${w�ӛ!B�`�Z�7k:K*��O�x6M]��,|��f�H� 5Þ����t�ۼU��=�����t������^�?c�� ����3e�m�uSv�Ǎ��hܢ�/-��[��i�W8lƻ��I����&Pl/��V_�ٜ��<X�i�	ҵ�2ܸ����7�=�߆{�緹���/��GR���H GH�1=�SV�*�M��mM��r�@G^�JN':W�a��bw_tk�v>}��oM�
��6fN�.ۤ��i�DQ��]�Z98��6֪yj���T%�Y�(�rv�{��m9gn��N	:��-HL���˝��
l	���T�+d}�x�yi<J��� z㙭.�Y��);��wbӻ�N�֫�ـ=��<��;��>�c=8�O]S�ϙ?]x.�b)8,�B�T�aC*H�@�F��,�$�a(I+۶y�YnХ%� ���-L��L�$�B��^$E�2@��2�$k�9�*$�RI Hì�*R��d�-q
�����K<%	RX�Zt{H��{v�p"����Gн����*I�d�$���IRN�)Y��WȲfI(K1BJ�B�2ެ�'YY�iSZ�8�����U4\$�$�)U{���t&��:F��f�.��=��I$��$�zL�@���؋�њQ��ݺ=���n��׽�.�#�8�]V���-J�d� u,!�҅[J�0]�_�E4���Fj�$w�|(�렮)�3V4�ݝ��`���Ն,��IB�N�bV�%�$�*J�2KԱ(R�,�J1>m��ġ2���'K��K&eB��T!��y��*J�f�m{��tMӻ�0? �g"d��g*N�	]�M��cwe����=ˈ#�d�IB-Z�%)BZ�$�BI([�5=�q޵ֿӎO�����>���������pM߳�_�  H��*-��`�؈��H ����
 ��H��
�(�"� �"%�"��*Ȉ�"#`�؂X(��6$��H� ��`"`�� ���  H���H��*�!`*X(� ���` ��(� 2*$�# (ȈH
��"�H(�	"���!�U��gUq]Q]�\�������(H%������"�)  H H��" $�X�%�H*H�UQ�Wuue�gU*$����`�ȈX���]�uueG]�Q�qW@�H
*�
���*Ȁ�`q����C� }����aߔd�'}oBX��M9��>��Nd�pZ�h����^8qM�]�Ǚ� pG�� V�(駦m^DA5��x�pCpsP�I�:�sCP�r���z�I#�x�����u���=C�udGQ�6�g�$ME�.D�4^�5� X:��9֐��C�:�'���$�?��v�-���ӓ�i� �uwR���Q^��k"w�.MD/�"��/��?���>�O���>l��y�����w�~i��O��᯺���� ����a{��;��j�M�|C�f�d��t�Mu�9������|'��W	һ���U�{M�1�Z��ǳi�<d��*՞e�Zp9�!���qB�1�����[a��jY�L�Ebz��s�X�gwy�ڶi�-��18�<��<���]~�"�{��!���ө���,���̉��r.�ܲ��h��S��NR��i�~�g=�h�{��@�X�A��m�ߜ�$Q%O�>�r����]��v���o=�q��s��ӳ�(�tpP��z<���E������-ݠ�~]��Z�ڈ�ם�D#�]�_��{\G�97u`g�G�ґ8��T43@;�~ ��1ŲV����T
ǜ�欯=�'ެ�Ns�w��N�w�S}�e&wK���U�C@v��ϣh^�&x��G�Ԕ�ޮ�<���{i�:�.0E�7~�qg�4/)3D�����@��Q7�UO�
C����%������;<&���� ZYX`�8+�lf�.�=5��S�a�9�2C#���J�?a����<�ǲ{��͒�gT���;<'��N�q��@d�6ő��v��I;`���~�8�+��5��o�9�����\����V��}�bi=�����(�e�_5����<�}(��ڄ��A����zf��¯����4�1|�t�X�_���/������>8�qӎ8�q�q���q�8�8���8�8ノ8�8��t�8�.8�8�\q�q���8�8�یq�q��㎜q�q��q��pt�8��q�8�8�q�q۷n�^^q�yq�t�8��q�8�:y�Y��w�����u�MV�l�H��1��ԟ8���۞�s��x����bɨ����x`R�AҪ��Lry�>�\{����H]�g�+r.��c�{�,ԏ.���w�׾����ɚ;ǃ���u�[�>s�7e����Gw=�'��	��}����S5�G��^o���yo��|�{�sQ����{)Y,�I�4S�6��->�f���|���6^�9��Eb!�d~^MJ�>ӳ���!�s�Z7�������!&�;�g��@��~�=:#����OPQo��L�X�6��c����\�ʿ:U77q�`o��W��۸oo�l{��=��?kս�Y�����G�d-���j��d�|�"�|sڶX{��w��sN�j�]?e�n��=Ko4���"��̗N�S�����v7��K||�>S�Ȝ��ٗ��u����ݝ�{�������L���s�Ou��Z~"z]v��`�|w���۸9�1����p��Y�6�s"���5-^`d�6Y�[�t^�6:=��K��=ރ[���W�0Q�}x��0���W�6�'�}_�yǑ�.l��T�^<�w�Vc�s�y��p��s��$3�y&�;X�b%���m�|Ӆ�����'����PF�p�P�ogt�=}��������!x�7"��{G@��������~�g��c�f���yv[�^�*��ӧ������8�Ӄ�8�<��<8�8�ˎ8�Î8�8�<��:q�q�n8�8�8��<���yqǇq�N8�8��k�8�8���8�8�8�8�N8�q�q��c�8�8���۷n�q�pq�q�zqƸ�8�<�D˲MD��,/�MZO)� �^U��D�U$�>���5�F�~�'�oMB[)��q[��xg>�V���g�k��=瓏��{�1��V*��t�7|���o��c8Y����XY��"������K=�2pe7�94��!��kz��a>ί)]3Gj���k�#������Sݪ鏀y@dc�L�fv�P�B)��}��Y�ͻ���1u�?$%P��>��[�mi�%�����Ç��U�>!���p|p�<^w'�v9����!>���a���C�<�����QߺW�XVעUضg��`Hy#���ONm�D,����=x�Hu��2�l^8`��!��Ut�eZDw�!���t?eAd��+���?xG�=��h���=p�힞`}�u����^�"��'���fa����7
��7b�E�"RF�]R���|��$V��Yst�>4��yE޼x���<��m>�cbC�w�D��}��C�wa����EhcD{��l/� 2�
_]o�gݠ�3�ro^�����M����,{���X��x���v�7��0���f��{Fm:�b��A��ހ0S�HhK��<	����>SҼ9����o���~|�u��G�Q���4w��{����TQ���֖M�%�G
� 4�֞�������'��ޏtRz�@�>����_�Ǎ�gH�p�zj��=�������}f�	�@u����Y7�2"\��v�S�o��޾���*�c���s�{�3;۹^OOv�m��1a��)!d�K���*���s��d�CZR�1���Ŏ�t���^%���C�{�����z-1�*^!Z�v���E�c�ts�d1��Eh������چy��;3�����»�I�g�}T$v,fNC7�o�]���[�{ɱ�ӟ��_$Z���h���~�{7�1>�~Li���Y=��E��b��#�ay7ޙ�gG��<I�l�)�;���v��k�땝��:��4�sxc�M�Lg7F�����r{ۑ�����
���L���X��K�W�v��0��9���!��O=k5�n�(������e*g��_��@\q*����K������-�z`�f��]���}��R͞��?zs2��]�m���;�;w9a~�����|�mT� Q��a��4�"�Z�W�3���Nz��_~��a�1&2�-%���)�,��v(���� �g���|<J�g���p�����n��Ow�\�N���B{V�8�a�t�Y�����8A���}�u(:u6�ꋷ��1e���� R�H:��7=���!��npc��۷$�\���E`��ww�7w���+;9w�u	��A����8�0�h:|���L�����t�����}��u�qq��A��2hܾxU<"�6�0���=���yX�������<<���$� �W�YK%�u���f�7qd0���(f�8��Ɍe8nM@B��^��g{ދ�}
D��=�֍9�N��A㛥��k;뙺�R��6�{���ν�M��S�C�i�=�m;��:=���f#ѿi�����ް�ZvD���lx2'��y�܊�}�lR)���{��km���M���]�w9pj���Qpv��7tb(���:��$Ç:����_�)�_P�G���Gw$_f�o��=6�׭Ai�|X�w}K�c�(��:�~����9q��bZ�ͦj���FI�
�(��q��;��������^�ǖ����{=�y0^�A��`���o���p��G������YҲ����lɩ&l�|v.��=3��)���_�],�{[3�}YzMU���s��+:-�������(��%=o\�_K�ӡ�v]�ێ������O7�:S�5?;y���L����<����������.���mԶ<$_w�z��;�e��_��Y�1��i��}���z���������-�,�c�̨%�=݃���}�u�.��6���[}�rg{ ��,^C/��k�(^u�!�}��|J�^�Ihwљ�{Vw�~�����9�s��S�9�M��d;�{�R[5����Y�A�}�`z��2�1�v{7=<�Ϙ(�����%��X�q���U{u��������o�pv�vnf�4�uưՆ=�-�j�zf������+6�}'�D�8�M��ȹ�p�h�qlC�Hc�hɕi���������|���(a�@�vv"M�u���4�w��������)(��=輻�27#^��{b�37��\��{��V���v{!��O-�z^^\�F��K������f�4�Z'�)�
C4����'���`>$��﹮�.toq>>Lp��B/7cġ�y���a�ثfZ�Gw_�o�}�ӦhĽ,��)�(�{�&���#�}�=�A�b��������DĄ�=ʤF	ze�9x�������Z�p�݌�߮�9��6�z���t7����Tp)�vU޾�+q<{�,�~��L���{;n^�n�Xw�M;a�����+#=�XZ�Z�6�|�"�KmY7z��M���R6Oy�{���s=��Ż�7���?Y�?8R]�j#�e������ý�U��PƼ����(E�ؐ���R^WiP�ZK�9�,�B�X+9�=��d�K�A͓���Y����/s���LyQ��BC�9R�h����7�ݰ��ׇ}�7�{�}���cZ��pdrw�q�`�k�9�}x������/��4��V�;���u�?,A+ب�������#��!�r�?e�T0M
)��H#Cy�#��РƵ̾''��,�"�!����쒟h�R盏�s��1�髻zs}�ם_K���<	�9{FAn��y����X%2gd��Cހ>�k�u��nߊ��t���_���~I�z�p��lͳG�8�79���lN�}����lhn5v:�ƁGo�- jw,P��촱�����S������D�i*�p}�І0׆���MNvygN���}�:fyy���fN۰CE����tC}77]���a�x�w�� =�cò�4*']�o���/-�8{�s�&�;PKjm�X�vy�	׋� ��r2�]���Y�|�)L�H������Q�S�{��7&���،�p#�j�.s�w���.�t�.Q��f�plh�1��u���>Ñ�n2�Վ(f�E�8b]us�uMk~�^(��yݯp��A�r��b[yN��ē��n�˷�W5x�K�f��)�8B�� � �+�^�'c�D&�������,ݽ��B}2���/e��s���#h�&l Yom�&v�}��{/9f]�G��3��D{�H+���z���x�v���d��_O?Z�_����xm'�[�n�(x�Tl;�E�SK����۹��'�2w�呀�Z���ЖT��y��9<�mӈ��>�=+���w�W tw�R�s8+@�`��wn�l�<���tm�7��gd�=�7B�\o1�=�{ڼ�/N\-�Nh�D��^�������8`��|���vu&�y?�r���9���t^������{8r��rR�m�Pv��>�w���j�P�}|�0v�ȏwޫ���a��K����X�8YR���y�l�Ɍ���kҋ�Oxn;;b�]FD����/{y�����FCrt�x��",�7=�ɐ��{G~b`�x���v�w���{�ďoy�����:��K��{��U�c�}�:W��G��M��3�/N{
 EW�髯f���#��oe�r�[�.���w����,Դ �u�V_�����eo��Ar�5e��S�^eH�XS�h~�S/t
��^�7�4��gz�e?Q��{Q�Gwf�́d邔�.�E?����>�}1���%۷��k��w��>V^d<��V'���
�1�`�I�X���>y��yr��ɝ/���ڢ8m8&�3۫)`34�Y{���A�
��^�g7޶vF�͌Jy�rn��f��AO=��=�i�or?&�?0M��-����j������~�X���{H͏}h�+x[��������_�}�#;�������'����4S7b��^�h�t���iW����@�{���Ѕ/�i?\�i�����э���Ə�N�X�y8�>V�2q�½��&հa55���\��V0��#�yw~�C t$r��|
"��ݷ�^U���w��;og1�O��9��������j���g��i֬
�ym��&fr
�g��[�r�M�~��<,�#����6�����u�'�*��ڐ�f��k���[���w�9@ �_I�;_���t4�A��_z{M���o� ��v�ZMuw��O����S(8w5�O��@���~��Y��sC��Wk��_S�o۴2����Vx��P�E�R���} )�<�)�sOzk����N�w���F���n��v!��O���Vvo��g�����FM>K�|�	��jY7LY�q�u���{�=��vo�(��U�==�(�3�k
w�zgz�_�g���xq�j��zo���U?K��ǵ���r��Ϧ�w�Q�^�G��6�t����	svv��&����P�\��U�w�{s'��u{羵�e�]�������d�l��i�Ո�?F�ݷP��h}�l�W�����ͼ����qQ�mvh;�X�&^����kш_yx�~�s��.��Գ(�ݻ�fi�\���A����'��g����]K�f��z���z�Go"��=�՛:�dhN�>j0}�o}�EĘ�H��{p荟��Xwݒ�^=ݰ���z��
������d�<���L�$�Y���Sk�'0��׃�Nާ��ǃ��f/&��NN��#q�����P��i]ff����tdZM`��`�ae�Sܯ5���R�i�����t^U��NhыI�!��T��x��?�v�3�qլ��:��\C�s�R�n�ASG���8��V#������x���L�Vf�9P��z��������>y(P���ܷ�ū7@�q@;և����뙴�eg�yn{�(�=�i��K���?%]��3C�ڡ��cR��4oS�u����ր�z�r�ȓQNjZs�ݵ����'���
+rI0�'�ϭWU����f��� ��Z�!	J �6�p6	����Oc�#��<gQl¡Z&���Ή��vu6fd���c=188L��_{})���w��}N�XHC�{{���<�������yxɀA�Mjз�9+M�>����{���͂��\����۹����U�,��ǳ�\?a8����P4X��=�O ��A^إ-�h�����z����M��k~�M>~0���)����T+Eش�����y-\?��AE~�C�������W��� �/�����������Pv�Y�װW<�CF,%�TĲ�����!��\h>,��w�d-+aa�&�`P�����3I�o9�^Е)���-���҄Ae�yA��u�a�vv, ����g�:'��s0݇Q����m4�I���¼�5V:a����A�M�.�mL�X4A�1�.	Gms��]f�u"f ���IX��]Fh�L��g�v��gP��J��l��V�h��a�V�\R�1o-�s��h�Z���c`Z�4$6@�,p�&��X�R8�p�B����y�v��Z��%���%J@[-��X�)i��00Z��f����\@�ٵj��e̺3+Vkt��4��`K]��k�U�L���=�W	�i���ˍ)�.����f��R���R6�d�06ڤs)��A��o 71Φ6і��ƶ ���(.��$j��H0���5B��Pe֯�J�1� Zf�	��0��;���2ј��䉲 �'M��֣�it2XG��p�`�5nn�Dt�ki+V2����۶�H�k
��ԯ$f���fYX�]�Ԋ�ʎ�a�`�l��+���]cl�h�N6m4�Bf��]�єL�e�
�T�̩V-6i+�v��hތLi,3zᙏ�xB �
g���{K�70�.Xj]�!-b�,i��ٲ��k)��1ԍ	��h�ᡥ��ի�m���j��-�V�Ⱁ�;X��e����-�1�âj���ڡu.Y��5�h���ĕmy�ճ8�&&ٶ���qT�V�eM.͖n�y`jM�l,��#m�u�5�0-�ca�ݱ5[��q-Vu�EB`�q)�1q6�u�����\(Ȼg��YpB��@6�0����.�9��ZhKĥS��P�$h��Ia�ҎxMfb�f�׊+6��B̎2����XK.�uÉ�`�Iv&{<�Z)h��]pm�1m� ��6�sN�R�f�+PЖ`�`��:�`L�\a��n�K4M�I��őԊ�.�+Z� b�[��S.���p��SF�����lz]��Tf��Sm�iT�	GP��JP�f���ܗ�`XRZZ�p@�Z/P�t���%��Z�н�m)�KB���7��Q�癘���c�`1�5�J�ԭ��*�)�iHˀaz�J�
]�.�A��nseX�K�*�WUn�kk���8�vD�%!ԗM^lٛ-ake��	B����F۬+�⎡ډ����7��+��̙!u%�TYf9�M�00����SZ6�HDsp�-m���+��ʕ��h�b&�A�Ś��fָ%BS��B���F�*]�s�vrԚSn3�<���
�7=SQ����f\4��.��8���v�W;�؀�&׵ff���P-� �8�b��udp$%�Ls�L� c�����[(k�.X]�[��p��4�K���6����T��icn�����	�ʹ�Y6�Z�t�.R�B��k������Z�д D���ik-5���vR�8�\�MT�d�1��p�j���KF;*������iuĠµ�b:h�h�e���]i�/+�f����0��,�6�RfQƦC4��#�ؖۃ0L�E���L��ٌ��n6͊�D̺�f�ָ��meA�R�P�6VLt\ר)�Y���c51�[-�M�b�c�K�ؕm�.
d\d�v�u!,M�D�y�TJ2�X\	<e�T�aMrYn��QZ�1���-f�jڮêJV��M.�֗BUm�V�m��ͳm�X��v������:�`�X�Jb
�c�W�3��d�k.�2�d�p"]F�Y��6��H�\G*@�F�����-6���M\�.a�ؙN.�UjL�L�,�h��(�c@0�u3
�6�Qs��6��h3Z��@�eu�f�S �[1PYe��1�#b�$�*�2���n�1ƂE�M ��F]@�-���fW��a�+�hk���Mcs��)�t�T"m���+kF�ҫ��.A��4�R�+�Y�d��\�B�y҂8�K`��8U�,F�u�طJ����W&���d4�Gg9�b�a�p�͎�,7�� �95��&5��.�3X%{KR]FU�������u-%B]Dכ���6����fb.�c���*��#��ȭؚZiV����me���4�ac�m�k�L�b
[bTR%Η5s��dˍ��5��R��"b4�j�[�L,mf�H�Î���o�-�]*�p�K���[n)sB��Ƥ2@؍�IQ�p�n�MYB�C]c.Pe�6!f�i�.�P�a�+2֑u�J�m�lsb���юM��U�J�b0�d)�vsH4n��u#3�hq1N�Qt�̫�sa62�Zf�u\�kn�]����T6ʻ4mh�$n�����b�Y��\j����M�e�PV�Ev�JKˬZYNжE�$b�hKZK]2FT�����H�0�Msl���)v�cm����[P::�f��X.%e�)C;7J��84b�X[�eb�Զa%��Fd:�ؓ6j�8���2!vv��J#`���̖ܺ�#�a
����k��[��m��2��v�#\�VP.��:��@Y��v�8ФRg[6�����֭m(m��+�����7-���W!�ؗJ�nih��2��5�0c
��0录�``�1u��P����.�9�[�w5�hDiP(WMs��N3-H\6أv���V[-Э�/R�)h�� 1�r�ٱ�a�LP3.e���Z�l�`l�&�r�7��+���`c4h$%�����mw3 �D!�n�R��[�5
���D�d�&]%�W8�DZ����:ܲ�Э��p)J�t6Ń`聹!��Moinٍau�]�(�7�.��B2�1�YP1�v1�s�m��f���Ҙ;&v ��7V뜳.�Yu��h̫-�YI�X0��-qY\������^� l+�a�[��ͺ1ˬp����14&�)h�eEweGv��n�\�{#[qn��4 �Ø�%&�Z�Q����R*����v3t�e�
P��;-��i-3��F��#,a���V˦^R�q�չx�@�m�Yn6�l!2Dҩ�������v�*�t�m�Zn��k���.�&�
mnnΆl˭��f5�U��.q	\�W\-�`�35p�r�k66&�*		CM�͊���Yu(iq��b�؁�34-���e�k�١�I]�iN(
ٗ���Ch�9�6� +��H�u2��s�mf.`�D�vc����n3֛��և`�f-8'uH�Ճl��6�ZKtY�[�Be�R��`�*ir�����������c�tR�5r*gvvG+`���e����a���9�t�L��`#��u.��az�k�r+�錈���K�GQ&!b�*�S��[fr�Ps.m���(&`&��!c."�-i��M\��-��%�ٰ�VZ� �� �g�0U-3C��һXc]Ȏ�����L�6X�a�(���ir�RiFRՋe�Qj̶ہ�ѷ�S9.�U��1�5�X�� %ձ��WMK����jڵ�4�7�f,,�V�J,�Fa[�f+I����m%�uІ�0]M-�%���lHH76m��n�Z4m����ə3� ��:M�憫�a��,3v��"]Bl�fm���[�5�iV5,i"�,Fl����ms�m����J覰���a��[�dmSM`e,̶��H,wj�ζ�T���N ��vh�y&�,�kv
6�����9۵��`g�l���+H�u��d��(��4���Ԫ۴4�����Pvֺ�cT�Ue3��h�McB�����R��,�:����sc.t[-�#-��F0�RZp�GrvS��J,�uJ�lJe�U��3l�^����h��-h]�`Ř�qT�.^�)�0��p	(�B��
�镲6�%��:ec�3��D�Y�f��̥�K�:���hWJ�Hg8��p	7T�]��ۨ�4�v�tf0�{�ҹ��`2��\�.��YlC�Yo%�X@�Q�[M��L��e��S���Ֆڰh��Y�kV��aM4ef��1)��J�[m��T���fe̩<��#��0[Ma����Ѳ��Ħoa�)i1���۱c��5M6��q75�a����1qY�-��T֒�{�)�aLVو�$RW��`M�j�LB��c�Xl��̰53����2 ��Y��R`�5�9�2�mX\�k4ŭ �B�	n���2�3���.vI�c��e&�m�\ل#�e�;Y�̸�Ʈ������v��x��k���A��-��1��KbZ�;���h1ŋ-� C�c�Rĕ٭H:ٴo4l-�F�k,̢8�ʻ;3��E[E��:��Nݖ:���b��*k�b�Uq�J��e�be�Y��`X!�[3ip郋kq�9��ɂ˘�ɐ��R�Ps(.��l󴸭&m��8&�@R�SuCmv��
��GJ���Վ��3-�±��Ib��Ÿ�[l.�Tj�Z9-j���q+JcX;
�1pi,�1B�H��-KY�ve�X%��[���uVͳm0$�h*�ѱ�J���U�[��g
��κ%��tr�fW:���Չ�Ti�Z����[�h���/@�4� 5:t��ݦ����F�ܰlu��,�r̖�uf�:�-t�h��/\��&�z�Aॎ4]&���eb��0�Qb��c�Bi]h�8U�J&�Xe�0Gg��A��1���5å���Նu[c�3��T ��H�NXG-�j��9��7�\l�ǖlg\���#\�b�-������з�!3-��
����ָ]D)�3"0�y���k��-u��Eݗ]"Uք$s�+5E�.\�q����F4"��ᮆ�Y�<��&!���Ѝ�mIp�<�o<^p���*�M��-���hY���5�-م%e�T��]HJ��;�P��"J$�bI
�}���>-$�g#�'6Ĳ��Sޯ��o����=��;q����u:�C�����Ӵ�mӧ�|^�Q���C����wŨ[B2K�k	���c��ێ8����I��!!E$�Dp�$�����q��b۷8��p�D���A'E5��pTq�X2��9�;lQ���E	����;:��(�q�mX\'kn8���:�����$�'�`��ͤHRB�yh���s�ϛq)�s۬���'e�)ԇH(�ڃ�$��g���k���nݘ����<�3W!I�Nu�8���?V�-�>�=n��:���p@ۻ"�䬬�H������Zu��:lHO[�i�!��z,��fex&:��3^���xtֵ+K(��V�{���Ye)�6�k����;���ٰi�{��/�һ�ܔ��9�ͺ����Y5���q�v�޲{�4m�N<6��7O�zYmu����}`���z�y�S�>z��9���ohIzXB��$���{��Ie�T�V:Z�«4f�	�Wicog8MJ�X�Bh����hIS$&�`��E�\���͇�F ����fF�X鴘2Q"�+lrR����f#��5�5u�Z�l+B�j���K�Ck[#SW�x��yb��	�܆��P�c��bZ�S�F�L�Zi,-��&A4C	����t�m"�0�q��m!#q\Sb�KujX�Ɉ�J]�i+�37	����%5%�yź�,Ԕ��4�"�IfZ �,�ˇVP2�e#h���[aX:�ƆY��˒6.�nۍ"#��=v�Ir��.Hۥ���[Q�f9f����fa+S�i�̹D�5m:5�h0д�$r�Ij�,��%�ƌ�����n*a.����ͼ���L[�.���A�g&�4(,��L��H1��ke͂6�ŪL��B[5�A���3�	e��̺�.Xml4e�0Yl@� ^a44�X�t����$�l����nq����	A�q�� �NSj�`�QaRy����݇;l�*�Lj�����eе�M2Ms4�fm�-7U#��k��p;%��1�	�Gf�p��mҳ*i�f#� �ѕ �p�.��e�#���5�ɲ���$Y�&.֘��1�rEl��&��ih̒��N!��f-anѠi^ʦ���mD�&ũ�XM.���V�A-��a��
����[5. �����j�R�5t�g-��3\�����k��AHaȃ��(X�6�A����hb(Z�	��J�3��.څ,�8���XSc��#(c���M	�1�9�ř�1�ʹ9 �E��e�t���<$���]6�CF�6Jiv��S)Rt�[�v��m�\`�'i��)2:7U��R��T�"[(f!��� Zd�&��h��n���ۉ�L��rk�2<��κP��kns��3R5M�-���i6LKn�a�Q�U�[�q:I'��Ť��ͥ�؈�/R�l��k`�i�kV�Z�F���cV�m[Ч1-�j�b!ij�e�%*Z#Qm��Q����PB4�� ӗ��`C�Ұ�RȖ2ڔy�EX��e�Vƭ�+P���i�%@�miʈ#E��m�,-#kh�Xر[e�-���,�i�0C�#ח��TZ%�,J��*K	Qg-�,\>z4�d��;<�0��ʮ�I8��ٳ��E����|jn F��R٘:tX�w&/Z!	;vpA31R�� �W��u���$�vͽ ��>�x�~0��a��.u�3ӎ�^�Ҝ���36�Hn��{+]����fYt\���g0*�F�_/7j4x�$��>@��I�;��o��5�E,X�u���ͬ����	��ۈ�}~[i��%�]E�;= 	��ɐH'v�H�sU������|1o���[ : ���ƓY��ܮ�ff�b��1e�Ζ�@a�ãY�! 	�gC9fpY'gQ�b� ki� �Dk+.Pw�fwT�W�r #�f��O�����N���g=��\�2*�W�y�ַ���]~��)��2G6�W�f�s7���e�u��/�~�ٿs����98��{�gv�P�_��y��ӞP�����"��}0	�y-�r��dM������k��A��ڠΝ�����̗�k�"&�YpL�#Ce�3KKT���$�KY�A#u��'.Ò�o?��h;1.^��n�x�l�v�`����|r�gk)U:�e7 ��&;�r]:�8��$?� �9��3�?Wެw�~�P$�F�H�k.s���S���v�����K�Z�3�vP��r�ki��c�5�@Զ�v��G�&���q�_~�>o�Q`e_!=z�� �����}x1MX8��{1���ÂC����ɜ��O2\�%�2�嶆��3>"A��A)��x�ƚvJ.#kN�H����'b����H;oq ����#fd�]��i�B�LK�6đ�7iڙ�]��NI���SR���̸7�]��N�=���	?z@r`B ���E��H������}>��Zp� ��؍̺bΝ�����ė�kт�[L�Y �[ �I���7����K�;���z5�?�lw$1t�1d�ȩ� �|r�<��ke�g����'�a$��ȀA9��`BV'W͈����=C�V���C$v�Ch��������A��ntY���y?~6�h͑�Ϝ�8$�9 ?�Iͧ�!���Œ��[�� ���b��,n�)c���&E�ӂD�{ږ> �.2#�y�@�A^��mT
�>}�6�3�Rt��=�_��/T� �Ŏ��[wxO���q ��Ӫ$Ld�c��V��63�����j��� �����z ���H��
��{R��̘��������?Fs��-�,���%L9m�����eΗ8l�o{b׽b��
3��4�f�SF�{�ԉ�z���gd:,\:%b�P���q9a��"d�^�W�C�T	����a��@Se�ZC��	�h�X�:&��i����,%
�9rM�ɓ"��mQ��.�9>f-�30���f��|wq��[ذ���w�����ZӪy!��.����`��Imw ���(N�P�1[A&�M���8�
������r31����6w��߶��E���������s�J����i0�uɽ�z$�m4���>�F�j,��Qt�ꁌ�B
���]LꙀ�#=�� E>��C�E��,��}�^|`�~�t�B+R	&}�$��[��"&i9���'ӌ���	Z��IO��E��R;���n�1$_(��,S��8����Vz~]2-'#'������8���-�������GX\�T���G(l�N�m�{D�!#�d��5�=�9���kl+Fe61��#�,���uڙt�ۮ�E�`�b3%3%X�V���RGm�n
ܢTa�k��J��� y�e[�bIu�isN&0��]v8*16Jٛ�!soe����J6]�S�t1ûj�f�٢�u#1��[@H�i�-tL���G9���;0��cQԚ8]K76���6eS )S�g��_��<���%���2gj����3-�,msu#�.и�0��
� �]�	��Y�1tȱp��Tcn@��xߐ�3�`�� �F��Vm��7$���PI#3S�C�Ό�$0.���s�ؚn�FQ����G}3�m[�A V� �u}qmVN�\M@U�-�V��g���y�\~{~y�#��e����1P$ߑֲ�r�b4'8���ŝ� g�M;�R����7��� �>�H�:�-�aX+p*�DӇ ��}��Yٙ��.��1�q�oT�QB1��Z��nߒ&�6�|6�uz$k�S���[k�*!��&��uۍ�B\�hJa4��9�%���,Iq�ʱ��d��'�{��%jE �������=��#u��ܣy[�.�CI�@��v6 ���i3; �b��|_VZ�	�l�uVP8��C=��/B�18yU������_b��T���e�}??a��MS��F{�B��t�<��S��y�����9�4�/C@�޲6_�֝K� -�iK,oO�>
�$0(���@���������~9�����⪩i���D�<@�|H�i� ��1N���,XJ�'7��߬,�0��l 'TڂA;�᭵S��������BV�oL]����t���j�B�0r�7M�R �^���$�)� �Fm�r"Zu���FE��NV�P%�1L��`J5h���"�R� WFbg_��'�n�-gjB;i������]����^�ͨA��Sq���ۇ���N�ڋ��D���Ӫ�"�0���ݝ˻��$;cl���yݭ�A�-��� �_v����v��^�\L>1����	ئt^d�,�`N�pI!y���Q�[X1j�ۣ�F��B�2�����d�y{#��[��v�~�k���5t������!軆5��VP��ˈ%/e!^���f�m@$��p��`����>Ng�����f�kT߅�cl1-���I>9/���=����z��@"!�T�A�c8�&Bń�?s� �����O�Za��`�^��O�e�I�}��PCLZ���8��w�{��X@'��A-D ���)��#m�����QKB�,mqX̞y��o�2�p��F�̨��;�A>�}�30��ݳTH�l���}[�����gf+4n�Z���~l��,�h�ߵz�@9�[�#��[nL�[�u0�T�͊�#ɗ,�L���܇;���J�:6�g8x�u%�QX�<I;Z��#)� �nM���v)��5ِ�1��}ˈ���k��D��I�i�Z�%��8F�A�뽑w-G����X��qlV��M���?����,�&�f����s-0FK,9L����/{I���Ѯ���B.���Lz$v�v7���Y�8�&79 �z��|H�i��n�N@ct	^��7(J`�Hvr\��5�[�Lܮؚ�*��-c�6b�|}Z|�6�)Q��{�?U� <����^���OW��c��w-B��9 �k_��Y?����	C�������.=�3&�h�H�eFO�e4��A{��(E;���Z$������p�$��̃8��Qj�9��4>�4IT(��X���!zը@!�4$�fvd��x�U�)<e�W-��/��P��A$�Ӫ $��*(5��ܴe�{<������H����+B@���F ?{�/����&qWx��k��<��:�������B�m�f�%�4F��&v��� �)��lx~�f�ޗH�4��,��]X���UY�thf�#C chY��|���~� �|��cCo��5tn��M��B��e���%�bT���ZM��3 3.@�f��m��,�.9b+y\닇1.�]��.+-��`1�45��]C:�9��ʍ����f�F�6%�jF��hVZ���,ņZ�3bę�ŷFQ�B��"G-�ք���F�	GE8��b	��-Ņs^�I�,�J�f<�lV&��4WZP�aS���ry����6�ݡ�K��,
�ÓYMV��r�er�t�|AY�2��w'-�31n��I,܏QxqmJ{�7ZZ�b�#Kf5��'F�	ˢ��3��wp�䎒�b�����@$O�j4�1�qÒkEl�#F($���:�-%���`���g`"��H��vw0j�[o�n���=���m����8t�t��=���npb#&<�	�Ƃ��ku���|v�lG���h�ol��4c�A1a$�.��)'���<��%~x��9e-�I��ՙd>z��x�k��58��y���g�޽����I�Q�������"8 A�T���ڮ�i�Żs2�n���翙�v.��4�k\"F�pH$��
C0�� Ę~���9�� I`5���>P�f�1t,�Զ��w©��1|�q�7�A�^u��\K��YI���*���h�%�wr��r}�>��[/{Jsފ����~W�����[_	���(�'�B�5���p����wo�e� A'��c���,�U��/q�����53㤡�V\�^v��e�&����\45�+�F;y�$܂H˙�@$Hݧ��:w�[��ipHl��,�8t�t��A�����{Mp�=nT]��I��� ���= �l���1�%���E�2�����biCAꅗlܸ�6�fi�����k�� �Be�H9�I"�&wa�����y]5��O�yg�j\�8��ȣ�@^�� �D[��~�z~?��HӇJ�m
���+ޖ�՗�q'6A+�j�	��_L���U�v:O��EH`ėw���}��}s�I	�o^sd�X�|���Ѿ�?����z�6ky8e�׻�6K�Y�o���ɓF�J��m8��^�:gxÑ�f�wj�p�Cw.＜�޺���C�9�-����w��IH�Q�ꇮ�Վ��G�������}�H��E|�͘���{��lP1�)m{5�QD�UM����z{���6sFv�4i��U9}BZ"�6t��P�����$,�S�Y��&�����o��uM7'`<fރ���ő.�0���{���~�GZ���<��:7�`��Q�wԢ>��Se�$ﯷw�!ˊ��x�g��w�6�g��b�7v��v��'�vy�{'o���9<�	
�w�]�=~N�6�}ܽL��q�`�b���(�
���kӷU�ߟ���a�%����9�q��ʼ앱���[��˾f����D��{��g�������YE�8p!�\M�Ǟt]�A�z�����~C�q{��;c�Kׯ�`Z���=G�3^�d 	4�Qf{{"�X���{_w��:���wG�x<���e�yx�,�]aze����U�%��0޲?zB�'���3�,kU"f��O_`.Ǫ�y��7���#�w�#�ީ>����/�=��&��ѻ�|�҅�W�K�F��1i��A�z7���OM���A�d�oq]�־2n�}�q�ݙ��W�����Lj�U����8���d��K�T&��zw�vt����L+�����{��9�=��-����� ���&�t���]����R�&8��=����<��{��8��2�FBL�ZS�IW�{[ڷP�z�{�g$��*i�g9��ճo{Vĕ���ףb�I�bK�	a�6��K
D�HK�N�I+޻�r�����||||q������Χ1����f������Ӗ��m{�����K��M���>=o��������Z^�;ӻ�;�~���>OOn>>>>>=�===�q�R3��^��J�{^mn��f�̲� �����ͽ߯��J^���[�ò�.�ow������kdZZ�'�������tۋB��N,/`�������sy�����r�tRB��B�oY�@���=��x��H��ܜv6����<�{{7[g�y�D�oO~T�	�aǫ��xNN�j����^�y^d�>�ν;�K;/mόO�IfD�|�'{�8�I��8����rNr8"��>�-�Ƞ���O�v�q% RGGNG��y�Z㏮ӢB"	}5_��>w���!tt��|]��觶�{o{vy�w��t�pDJ����J'>3���C�/n��56ŵ�	:�a���������Q	�,�u��ʆ��$�K,mG@�>�$Oh���t\8fs#�ng�CT�����Z��=�>�'����Ӧ	��bV��z�9G��PlK���<���<s����W�n	b�x":Vj��$x-0�S3�Y�3<܂le��:��GP]�� ���8��1 ���i� ��"Ur��Kÿx��GP6űIx���G�<G��x���w��8<E��o�Ki�Me�VTvf�Glj)Fj�Ɣ�hk���Զy� _�������'~�bX{�������b�����u���Jy�s`���<ν��a��y�{��f�w��*�X%>�{�D� �A��R)&��bs���,y�Hs����g�s�Y�f1x���yL��	bT�bW�8�6:���)"�>�ǜX��@>G�>=�{cY��"yG/{��<"-^vf)�&tZ$�
(�G6�xIs�}�A3�gg0K)����{�s��h�iV=�l��4��#�@��z�F@�[Ű(A��3���q�r$��$����O��"9M�1�s�\��7��js�- X��[�q�!HX���P�<�Ȥ�s,R�W.��{�o8��8q���iڍ�K���I�1�D�@͗k�x����4"&����)S{y���8n�x���,�!��3S[&�vIըC�z1� �pA,�����u�,/��}M�h�l��O�t���S�$�rB6�u�n.��8�Ş�y�;��9�
s�s��@c$z�5ޏ=}�΄�Y����39*fa&2�{[n�%&�DV���࡬�8����j)k�ؾC�|���(ir|	/S��z��u��JZ'����y�l���/���	"O�G��lc������C��GQIql
A�<�19�bs���/pqd�k��Gpz ׽𛉸��b�f���=ދ؝�ֵ�<��B�+�}��1xc����ቭS�=��e{��G�1mz�փ�ٍ�{�� y�tL��J]4U�I���'}��ME$E���:��w�lJ��6�Mݽ5*Ǘ�T�1����>���{�b�@�K���w����hwfb�2gE���|#�r<�g��rw�{9őI�O{�\NH%��XP�XS�{�(�)"�;��q߼��{���j�3�q�2j�~�b�$�������穦P���rN���y��6��A,��~r�i�]p^���@H�p�K���&�RX���w�ۺ��I`{����H6i�7�q�3��йe@��|��E��u�:���`RND�Ǿ��e�{^ٗ:|Fh�xF�9�\#�#��A�nnO��H���ȋ��(��#���<#h�T�U�ѭ]�H�vG2�J3CKΚ^#nњ�;P�9�w6Z���e]
�X�z�خ�!Ŧ��U�6�sڮ��,˥�[����.c����Z#ۍWQ�E���,�3Cl�1Ev�f�s����B�\��ki�Jئ�`��5,���
�,�h
�
���U4�p[�*WK:U,L#�--��]��h	]�[��v�Q�&�9�_R�^�Jm�T���.�+̛�b^�[�Ŧh��s��b�Tlt���>}�����>N���@8��x��cX�H����wűI�=����@���Oo�3�2/���$^V�R6xB"�O�$I
R�RgH�b���r���u�)��R��x��\�t9���)'�K��{���$RGd<���uql
Ű=�3s^�d)��<k]��G��QW�����n.�=A茅��{���6@�l�ב���x�G�dB���s,�v��}�{�A7,��)iח��7����J f��1�D ���,�)��w|�{��	�O�&=�r2��������`V-���n����bX6%ys�{·Q�X��c�sċ�n�M�}7�R`���lB���o>� �jW�ӳ`Y�3D���܏	���JZ&{�q'$F��w��}os8d��æ!aL����RGdƐ��;��Ű+��|�9�D�O�����͇=�Z�K%�E0g�3F�3�2�ģ�m��s���
�amB&����ao���D�ń5��x��Ù���쉸�-�H'�����x�XX���{�;�<#���א��n�������N;ސٺ��#e��q�r:�H{���cF\�N���}T;�$��đ:�Y,w����͍yy�IQ�v�E��R����p,R��!ʍ�C��=�Gqo�u\�D�w���ꦩ5�z��댽��[Z�"6�sޏ�p*E�+Ľ��6:��;H�������}�O��k���Ǌ�R� E��oz��<�5+JL��Rs$��X�κ���)mS�F�'�y�rA,�
D,5������o��d\�"ض:a��>򜳈�`R=I������������+��N�=@�"0�[�:�������xa���Ŭ ��ϼ�2��$RA4q�<Ȥ�H�v��=ސם���������RN�	e s�w�GP�D,)c���u)v����$~���Ҟ@��byG��H>��5��_N�#�L�b\�oc�;�`ؚuWQ�<���`��RO=ޗl7<=�8Zh3�fќB�CY�!y�A�6b��A�d�/[�M3v��nP�C R�Z�XZ��?=������ٛ|�'O�S��>�����j��O|�8��	b�)!z�{�!$I�8���0[���iOw��"ش�י�'0lJ{8�C�: �q#�G�����	�O�����j�֌x��f�@�y���y��Jm���r)";�)!�������F�u�.qhҧ��zr`y�� ����.���`xIs�<H��0�l2u��n.�P������kc�S�nN8�(˕��۩�[T¶�����T��'�Ő�}G^�۝�'�Ǯ��-�'� ��!�p�[���[�\�^������5P�ׯ��}`��~��RH*o���3n�����1I˃3�ң��29�j��8^I�G�$�,k�i5�L�kgK5ԥ�s�:1�x�H�C��$'�i��;�N����[s甑9��'���|�{:�Z�p���U��`S3$���i�QI ;��ZBV{[�k��.��va��):�W�=�6�Ͷ�CjR7\�;�6�Sd�+�F><�.�BdQLœ����� d��$W�k�id�#��ھ���z��	����{���`@�PI)j�i��S���H'+	9m���Љ���7�m����q>��D�m�-2H����ҒW��c/��K)�z����L��0.��%Ӊy	:ٶ�%��K�PK�tI�C���y�hE���K[�Z@Iw5��3���.���,]����/�l�U^{�I:�����3K٭�-)$�@Wd�m4(����&���.�Ȳ�������[S˄�Z�{�3�Ղ^ɕ�<�]/ꇨ���md�΢{���77|t������O���֠�[>և�����֜z��
t�)�NDϗЫ�]$�	W��!m�f��|�N罛�^�k�cU$�Iv�����H-��o���)��,�}�=�E�-�E.��g��J�ܶ�:n��A΢�Ȩ�
�-������v�+[�~�����}�� �%��"@t�'0{�D�K*a���x-C�l(h�i�IB�����.n�'D$ɒwiiO� �~I�X����]~y$��}!$�Iod%��jўz !c��^��z���;&`YܳUW��ܙQI%ێ H+��0	FZ��\+}���70�)$�c_K��o( ��;G
�tt���ue��Νې��{�P�I�Nļ���Y���g����z�YuGcD���e$9۶ZRU�8��ñp��w���! �'�n�C��Ji�\���z4$�[gKJK� �6S.]$����W\=��1���{y�c?ޡ{�ӷ����(�j��I���xN�7��~��<A����Ӻ1uG�b�b[�~y۾�=�7\+m�e�����޷u�C��EkZ��� ���Bj�S�	��֧f,ŧ1�e���3�TԻ8Ć�d�Wffi4t+6� Y]t&-��3��l���f�r��&eIm�
��6�����Қ;n�n���=��0a��AĮ�U��%܆+`9t�,[�R�7Lu\	4R� �Xe�h Y��#���i�[!H�K��%����kX����LG8{Z,fځ��ۨ%��w�����2���F��06.l.�\��ݵ��X%��m"FgA�h���)���mg@:ϖ���C7��5��!J�o3sGƤ=��z��玖&RAV��$;n��1v%�N�5U%���<��ogޝ�}I����I$������(��˹�#��i"���: �,S������@6�"���`�%���bi%�ݰ"�T���%*���vb왁gr�ª��[�ӯOO�;����I(}w�&A$-�e��w�t5݉9���N+=�H�v@�! :N�wd��ZBN�n|�I �+���s�2�[�Ǩ�H��pfR^I,m�i�RI{y)�������{3n��]�ID-ѬTZ�Įft�1v�i���ј��7w����A�gɜ�b	�Z��^RO��O�Ғ��b���»�!��Y�Ҁ�)5�[Qd��$�&s Ǫ�uGL�H%�E��f狥oc�g(�ݠ��fN�Y�G�cku�(?rLCg�b��]��ӓ�{m>X�wT%���;/���wq�P�A
֢�l�u��Ͷ��K��Ҧ|��37s_�ґ,��*i����Gʆ�e����)�v�*�%��j%$U��%;2H%��$��70v��a"P
��T�Ҋ	v��j�U�nWa�33��@b�o���SO1s���I���ZRK���k�c�������Vo����9�$��}�"R�Θ�$œ�MT-��2�y%�qÛڼ��ۋ����y@I�T����X�I-���*�",<��E���8pR��7GG]��ɡ5�.�C�v���m�P�EFW��z�n�wd�q~���j��;��$:^H�g��	��+I/�-P�[x=��3��Ey$[^KH	,�[r�ظvqO�T��@	�tc�F5w_{����PI��fKJI#�w�zIsnCvyZ��G�u�JT9��.�N9 ��l.��:����!-�??]���.���gΣ=���2Y�Q�D�ʮ�i�7J���^������M����?����9�����A'{�nw�!��pk\�����Z�P=��f�?$�K9�$��y������gA��p�1v�����o^���$��O���S$�U�:��)I*��@d��S�B���I�,��tK u�C9Ƀ�s/)�`9�o��;^�K���[���b���Hf���S��%*�N�����k7P<����;th֤k�^�ڀE	kH���r驇`���n������1N�N�6o'�}2��`���=�Hg�zh�9Vp�L�b:8���~����soy�����n�8��>�
~���А�E���o�=K�%�	 J� $�^���^�Ip�����X�=��b*�8[r�ظvqB�#�ВI,�y�  �K��jt$�W��l �%y_l�PIx)�3�J��5S�)�L�L�/t7\S_	��t��c�P	$�!�z�H$��$̀��)w7d�M�G2�k*��"�0w���bE��g����2�^�C*�a�����ф��22�JBNdL�Ryl�)�59����	�7��>&? �"���η	
滋ӗw.Rd]���u|�(�"N��b���pu-��.�O `�	!3"<����	k�I�E��n�iI��S;������d���������ak-�QcT�`��n4{T�ʀ ����;�]�3�!�9v:���z	 �Ǔ��2�D��ݒ��VG�c��T�r`$��2$ϥ ѽ��:,Y;��D���a�<���"�ǢQ})�SMҢRC<�3�얐�@'��\����Ù�:�S��ܧLi�O�7,�,<� ���t����2 ����b.{�2��a����m�2�Ƀ,��)-:V�ñw,��qwCY`�Y-��Ҽ��Hf6䴤�K{ _@�ܱx0�/mҦR�l�IN�E3�2��]s.�D�k��.������`�Y��|������3z�m�u�prst�Ҩ!<�լΰo��F��S����9X=7�Dj���h}�icul�Lb�L��бwcm�*ǣ��eC;�-��#�;�B��x����מ[�Ok&u�Ǉ8$��ܺ��9ðs��u)��#�����ӻ�k��C� �σ�ލ�'��=Oy��ʭ��{�����b[�6B)�K�Ȱñx�p�����﵉��U�˺u�tnӂ��K�ȯ{ޓ��Z�hAԃ��=���m	����C�W/aS�����{=�?�nz��tGt+��ݵ vf�N��1v��_>���ʼ=��l/a�+����c�}�+���]�Eoi����$�{���<N�w�>ժj��r'��x���Fy��������(x���4������Zk��n����Kμ[!�{Qty�W�i��֮�y��6���ޗ,39�{/�����o�=������"����<PLlC�WTd0SCVHXҧ"T��&w&�����){�%����>�[�<�	9d���l@a7���Y���50�]����~��O��.\�>��W���O��5��������&z?л}�-ٷ��xv�m#{��'��TL�\�����g���|���g�ҳ{�:ΣSpg�]KP�ؗUI����7�g���������LCG'R�6�Z퐷ja��)��Wu�lE�V���Ri�yg�q�lew�`����o�px
�3�w����>�C��\�9��Y6�����W�F��/u��8�68,ĴFҜ>���;v�GZ�-��"���<eo��$sڛ���yd�\_� �8N|��q������|||{{{e�$�HH��98�:��U�DTE�۷N�@�w������z{q�qǧǷ�M�RI$�+98(���!�M��i�.*H�˿o,�D��D�;������7g#��\q�IL�D\wݼ�(�:#��S`�u:����q��E�ҿ�tU'v�(�诞��E���:����:���5X\G�tqQ�]�����Ӹ:���X��v�#���֥V�tQ�I�FVT��#��.C���첳����;�����䟷��������өAl�2�ZTf���D\�+2��+e�le�E�F�aɵKl��֐�q(����bX(�L�����au^�1L�ԥ[f�$�����d;l�e�Z�6����uu,]rf�����ōn�n�f�M�� ܤ4ڻl-�h͎fec��-J��� �
��ơY�m6b�n���@�[F��� X�Xb&8	Qmw:ô\�]�#��p8�ͤ�f��4�ļZ�\%�̰�b�F�mYe�!ưk����#�`u68��":mm�msvG5�y�k��+��YCV�bl4�;F�QlCm�,j��A.�e��E!Y\:��0�F�4���)M	�H��XS�X�h�<�C�4n�-hb����7sT�x�2D��j�G@fu�˨Ɔ�u�� �I�Cf3���х44��m�v�м`C31�����c�g��$f���io8����f��I��F�\Ҩ6��c�C-5��Ri���#3[,X��֔�Fb��()���#�5���l�����U��f�0�!�[3vZ,ҁ-�+SciMA#֖U�PXMf̓m@�� �4�Q�AҤ֎s��r�K6Ks��ڻFai�-��]�X��)\��+�1hZ����Ӯ�L�WChf�WG%a�5�����k�&3R�	��-K5�Ț�%bUqف�+#�a��fZLU�ie�1Ă4��K�V���V7h��5a-�A�+ �X��mc�� �R�I�uңF�Yw:�2�YEU�F�{�����)�2�5�YH3q`*�L9��ys�4��4k.sa@,���	NvLD:�p�t;HgA��+���5���#YuԌ�z� 1�"Ut�:˱7���b�6ع�5H��F[n\M5E��t��c�)*�v)���ؖ6����0V��c6���9+����)X����Z����eN�
��	����u��L^ٮ���4k(ٕ�,)���e��U-!E�n��Ʒn�4%f�#��&m�!hJgl4�30��h=i?��/~�@֠ �\5�aΥw5!�-Ԥ�A��L���r֘��ل�\���n�����r�5�D��R�7��ƭv`Y�Q�]VkvФRb�k�ш#�!�xM��"4�5WM�E�Ʋ��K�HĖ�J��p���h���s�f��CCP�`��:�.cH��.���[�B JM.+*�eź2�l7b�T�]s�Q�,Y�Jb�B���/�����<���������%�٫���kAaNܖԉ+3a�By<������ϋ�.�]$����zl��i$�����7���ff�6P��L�E�b�-S�b�g�+�떘�3��C9b���e�v��B^I�؝�+���f�ƔI/U�\��3y$��B(��0b͞���E�r������p�2w)��j���	 �n8�!	-}!�36�fִ�3D�ն�!0d�[&ZAD�x���H6�Ȳ��N�:`��� ���Ш-���	N����y"P��$Au?J�����w��Hg�����IP�°.�r�(U.�����3�Ҁ�������u�T�t��,̒���Ey [t���)nV�ݷG��;��|��H.rMZ�ƅ҆2D"���`	�%��`�ZO,/�����Ng,�W+fe�H��p�^��*%&�@��S�;w��rZBK�ț�p�<6/h�b��f,�@V�٧[�CH	*h�Y;U�Ýw'f(�˘C�����LeG\ �dSm��C�ߟ�+y�|Qæ���]��fQ���~�+��@F��
���}럜[m���Dx$)}O��Q%k�)y�ݶ�f��+��%�\��b�gpK�q0_yÀo�$��%D��2��>��n����OspI$o1�B /;3��J���wA��2d�Sz���w�� w;��[��=	�Bu�T�	 ��ܺ᝞�U�=��$��߂Ș!,��Y�t�Ӧ.�
zI��$4��[��%�*ܻ��vp	%��P �I6�J@�b2�]0�B�C��Խ���nI6z�������S-, �NVi\曮04��4X.q��V�샹t&PK�a��p�Y�
>�u��	8�J$��]p�p�i��C@[�Qڗ��H.��S)�SNwtS���j��W\˥乶
�6�=���p�I#�;�iI3�.뗔�I�i�p�"��F �կ���wwH�v���kuL��	"��\9��*�|���uFw3{c�ةY���ȝ�b��შ���c���E��r8�K�wnɾy㜝��6k]�TZ 5�U:�y9�[KgY�����G���9�k1�Qb��gpK���'݀��
��*��$Y��$Hi@$�Q�m痐� �.΀���)˄��یAK�Ձ�0Eb�d&=Y3�}���&�_�{��ݚI
�RH���r��Im��}/���.���r{g�#55.1t+(6������7GazǫS3:tn��}���Ʒ>��COHiA"t�\L$��Ko�DyO��/�k-�~�ۀ%����	!����z	/h��dS�vN(U�P"I�_s#%��fL�ҍ�3G�۲e�$��]}"��_���?Z׺���~��6��5.�pY�	���ˤ�<�:�I$���l�κ��z�y&�n�i�Kʼ��u�B^���3���UW���Cm�ts�����$��-gE:^	$�B���&BD�U�׭^���UMNV�ҎTv*��ۧ#��5��wzk�A���.�q��	f�xrG���%pˇޞ#�v&^���c3�����xxo����Mj��l�g=��w���|�{էӮ8	v3��������3�ݶ��#Lg.���$���>7S�M��#�$�-j�h+ZڇV�3�V�� �]Ӗgp�n�E���Z�fc4r�A@��3��+\��{����(���6� ���ȄJ	nk��@%䗶��L��Ujfa����4
[�.	�fe��n%6��9p�'F�]6��J��gsI��5Ѿ��I$,v�@I �����$�_:jM��> +� rw��gV�p��ŋ���I$�cuHiI/$��c�g�:�_R>^)yu��I.��S+r]���wI8,΄J�BHM]-jn�`�W�$A��õ��	 �����8H.���=��I�gp��LꪂQ��-($��ˉ���̱��$��@�	$��d�ib�Ij�y@+�rHKjA�q��p���ާ�ٽf'�0���R�ww;p{ӯ�n0;�c�
��[��q�1v���w�5�	�n�x��/{ɸ<2�WR�i,
|8^�!���$#���>� kZ��v�价F�j�k�X]� �T�r[cVfZ]-�p���s5�p�%��*��V�\E�l��:�b%k�n�ƻ��a+V3J�egM�pUikRY���b�k�mF6�^9�[�MD�L��B��G��0h�`������]K�([[V^4�����5Y�l���Mh�ô�
���F2�.Εax6�8+B-��c\�a�7\Ļ�-x�f����Η3��v	��X�ZoϿO�Re�bC��P_5�ЉIv����$�\��\�J�3v�$7\b��I'���SOn9�Ô�ݙ�i9�����S�r;�z"��O>;��J	M7J�I$��7u��H��F��/;��;_�L�ݜ�.�L��J]7>i1�̸�L �RA-i��{��N��ct��RGܻ�BH`�8�d��wN(V�����uC�Î�b;�$��_(��@?����r������1��1e��\�/&�$h|�2���5)��:!/r���	fo%Y� B��;�DC81Qi)׋S!"O�w\<�J[}�����bX
K
�LFfI�tmkY��\�4fMқf����>M�t&Ź���_^B�`��3�(;u~�K�l�RD�r��3�I��"]3�3,ݙƹX����X��^}~fa
�u���w�zO}! �Uӌn�;�f�(�.09܊/tȝ��>1\c�s�<}+3l�gK�Ii�X�V�T#I�/oo�ھA�&�>����rҾ^}�M��
��LL�-�̽�!��~=� ^������y�z����?3W�鰸�$���"�y0t�rmq;�`-��ӝ�Awp�9wfj��y�d@$�K�\G�/$�
�v�]s�)Q�w�4$����r�@$v��	z��ZwI�9)�:2���i��G_w���q&5}"R[����.�3 ��)nޞ~E�85�S��������È`vd�]�8�U�P#АI%X�J:�k�[-�v���}%I~�yI$���!�i���Q�-
��v):
ݓ��t]�å�W-�p�q�*X� ���ee��T4������8\�p]�ft7�ʙ�D��� A^I$�S�����^F���h�����	 �2��������'T��*0$��6�S��[�P��A$:�	 ����K�u�6m�����@�~���y��.�^@O��y%�*CJ�K���F�Pm٩���(�5X%䛉Y!죵X�i�Kf09O=>ɏ��N
�	�ʲDL���[s[�U�[�gFN���ȃ�N�n�E_� >���{�5���x���m��缛vM���o���R�-=��wS�vf������T�-E�8QUL���I'�p�a%��JI��뇭��+�)guw�R
��G�g#V��vN��gF�^f�k�O�'�WD���oC���t���#�%~d����)���k��&n�w�툸����ϘF�m҈K�k�vbJ�ֱ5��useZ\��F5��>K�!�ْp��Ǽ3�=@�	��n�i%�.����f2}�F��[5!H�v��1澘L!�gؖgB%i��I)��)�L�u\�$I.��S)$�^���y�I-%�n��&8�j|�|�A��1w,
p]0>���ZP	 �Ց>���;1� U����J����E �����6c� ����.�^B|�]��m��
Б--�>iH��0�n�r@��]}v��:�Ai3�k�I���M8�G�\�^�Dx�בA뵝���b�N���{������#���=���8~|:����8�6O��_�Jր�υ����) ӽ�p������<!$��`>�q"Y+)��,��ظ�x�A$�e�$�����.aufж�[�z���4���v��1VZ�9��U)R[B��L�����\�\h����پTf�͛8'�f�����)���H��^I{� D%{��$�D��x|��K����I{i�0:d\;���G�\X��7j�g���wV{3|ҀI��sW<���)m��P>E�c����`ʃqE�����ɔ&p\3v+L�L�1�̫9�z@$��+�a&��9��3y�����^BI#��" J�8�rΝ0)�uUIF�P2�|��	$��TH��K�*݈�1��f�"��J�ݲ�z��O�p	Q��y�f�F"��9%��@m�!$�]��->�ȷ����ls�IZ��yI���5��I��JeU�ſe!s�V{�ń!���[��v���c�����ʐ$Vb��L$H^���f�z�;W�����r���*�|DZ
��DT/�B�3RN���.�ƹ�5�D�E��\,�5\�JGf%mfؘ��`:�Uؕ�Zhٛ.t
�3u��:� ��0:�b�6"���c(��n�a
.�,�n��2��B]�.S[rVl3+�+��n
̔,���RWaCu����%�.D��9��YV�fqtmi��6��C4�Q��� 씸u�Dc6���if�/�e�|��R����i\�n�6�ju9\�(W]h6f�������p����No�gЉA ;5�B%���)'���pXۚ��V�����$@(-���z�-;����gFZG��j��H	*6s0#�S��c� ��,-�G�H$���)�Sw���wLz�#�%�^�X��س�vwcU��m���	N7R�I���t�>@����au?R�%\jr�:g%�"��$.1�3��;��TQ��I,�p�����3V?R��$�.뗹�]q8��� �/BH�p���&�ӗf�UD�7N��K9eĀ�	������0�ڒ� -�"y5>R�J3�ݭ�,@=����3�Ņž�f��7�&a��H��f�y,x��V�T��l l�*�!1�������t�_���s��,�rm�$�$���@R�\{��s<�&'�p�H��R�J^M9������=T���@FRZ�>��?ߥ䘴��6���w���l���+a����T�^p�m�&�zZ�f�Й��y��S�^_.�חë��	:��މ�7�+�	Z�Ox ��8���3��7W�^	v}o�JIh��jc�@����:wL�:.�;�J��73VO��$��. �	/%�3#y<�y|n\Y���-��I��J	�w�ooEę�Ki�0;N����]�=@�!Sy�m�n�I�nZQ�'��-)$���|��)e�s;��HƴR�@!Q�
��΋E���~��	���
6k_CU��j3� �H���)��:C��G)�~|��ث�y篾|a���"��)�q��Hl%���f�� ���ͥfl4�`O'�.��S}}�(�ʐҒ ���e"W_@�]�E��ջ�d>b�D��)#e�	�IçR���� <1�'����Q�R>E ��˚4K��q�	'�f�^�Tci
Ĥ�p��������>]�o2I6k��$&|.{�kh�H��i�xgB�1竰�+YuDV49g����ى
�
D������V-Ěs-��ur303��2�Zx.���	�=	:� ��q��=�E��WQ�$��߾Q��P����=����S�=�O��~�����_��~���OR������p�a��~K�.M��?a�nnκ��'k����(��+�a��}~>;�ǻ�g�v�6����E~��.떖�&]ϫ�sRC�7��n���W|�C�>a�C˯�M�ֽ��=D�^��w<��/"=�.�-C�"��'OI�\��	�-�!6�W�=�ܯ�qx�$���n�U�2���.hhc=��'-yY��W�\���+ϼ�[��}�7���OU��x%���q�kؾ���a�J��Z��y�8_nRd�O�?,��oN1s�rb��YH��I��(/`$v�m��:vX����>������#ށ6��wzg�>�`���s�m[��L���Ӯz�7��Jp������΂M������p�]ܝ��Y�?`�W��>l���%3j�}�S����+��h�*���{<�p�C���l��$��*[뾦ή7����*��������=���l
d��~���P;���7��tTj63���x�k�ó�7{�œ���s![�cyh{�K� ��n�A.��蝠�1���|�Gg��78۽�ޞ�2��74��Q�a.ūҞj�®6c	M�bda�dQ`I��\A�_]�A�B���������8�O�on��.:;�]�uw$$`BH�B�8��==��8����ۮ�T�3 X��0��u�G��m|i�Gp{����N�8�8�H�>mGǙŶ(�]�G����h+�:(�W����8����ITu�%�E�_>��wr��z�I���8N.��
��YEm�"����Pt����'PtG9tI�_W�t�,�GrQO�q�^u��(y�998�����Y�����u���]���n�(��]���[Z>|�swm��{����B�z�13�39)3sH��y�����kw&�G�ym�!��I$3�BK���P���m�-�\��*BQBx��'��A�]! A-��PҝcwBY������Nyv�& HηR�*��2�osONK�3\`���4��c1(m���e���6ŗ�$0���2����V'ftX�7�Bʙ>r�&��D$^I�<��	��e������i�c�)$����HS�L����0L樜��P��גZ��M�q/m|��� �H$�w@�	/$��~��I5��~��ym�� ��{ɘIçP*�8�	$M�eH�<�I$��]���ZS�c`H��o@��g��L�ѝ�p���.���^��+����f`	 ���8�I$�Ot�R^Iw7d���v�+��e�!c_/KK�%�\h�v�t��-�Ca6�	&˦ա̌7�7B�6w8κ���羻˾N���S�+Z<��Q�� �����v�;33��b�aJO�9>+�$���W��2�ŋV�	!��"I#<�J}(���n�iJ�Z��]��k�O��C�b̑N�
s���řa{;�X�ji��^l`��m�v�g�^�{�2-g.읝�p����	$�[m�>i%$�svKHK5q�*����;Pc� ���L���
��΋���ƫ˥EL��J�vSsS:��b	$���)3䗒�]�ē�9���n��H�	/B�wL��3���YM��&I^K9fD�D��8�+�hm-l�:�ݡ�I-��@L��C5�%�33-���0,��N�-������魵$V�-$�Hv6d��$�]}��@���~I #��L��Z8�wr�'wN�@R~W�!�H��q���^m�����X��@.��)�_@r�����U1�zH×z�%5y�Z�����N+��yor�Z��7.��ğ�9�.��젺ti3����8�2����N_�@kZ�wN�?��o~�wj0v�W���f#n�CM�u�P̶4� .rZJ҆b�]m��-�C����ɼ��6&���ĸ�t1�6lµ���lѵ�P嶫.�q��6����m(L�p��Ўȓv�5N�-Zӳr�^W�(L�YN���GKb�Zaxds�Ss6��ٴX��g#E����7�hcK:�f.���i[4Cd�qn�hʲeL�˭ض�g5E4J��"k���}?�:fg$������߆iƹ�r��@*��J���e(�Ȝ�O��Zڭ3%��4�!�ݒҀH{�7E���]�;;���t\��C,���r��I^͹-�J�	.ȁ�+�ۚ0]G]b��|`�N��,�L�u�,e ��^�� ǒ$]<��gGv\tJ�x$��ۓyd�H-����.�.�]�`Γ3����sY=�'�,���}�`%z����$��!$�S�w�;gF���g���K;[�ZBH����$�өy@>l��I_cԠ&�MnoY1̯%Y����A$������$�n�2�m�)�lӇAN\�	���ud�:�t@���B��sn3�]�����5Y�翧���:wd����&|�;1;��D"T�5oE�&BJ6ɧ��H6��k^��$�A^����l]��I��)J:_��J|6��;��KS���즊Ȑ���#2��yrU����w*z���>�!흹�᳾���������f�;��o=^�Ð����5�A^��n>d�I!l��J{��E$�q�"�$���BOC��N��;;��4;шH$��n'�JI(`mS�NȵgtƬ	��|0!䒝�2	��%��3�D�wfet.�>95ڋ�̈́ߒ��o�"RHu<�&,Y��eDRIk�i�v�vLŝ&gUD�s�yJ	"�.̙d�S=�|�k2]�/	&<���|��H����$k�k�>��������S�=M��H)]���aTє�Z�p�+�WFZ�]�X�;�����ޮ���o��_����G�x�RJ�G�Sr��y	m�+c�0�4�@$��ȣ2��5�Y;�D2gd��oP	�VÜK�:�ǵ��n��
+�L��>mس� r��r��e������[��jظL�̙�ʐ�����.9�!#�RY��u�_j������NrcY]�/�Cp�������X$�ѸG�ի����ª���eK�d��U�<69d�����l� ��~���y�Sn���ܻ에�����K'N읝�\��]f�����obD��2(�y$��nK�  ]oŲn-�v���&}1��[���uw8�J+@8��?��c�Ē@V7�'��Q�|��L��OF&@Ixr��y	 �m����B�1_�O��_�<k��k^ԛQ0���,.͈�5F����������.��B�}I����Em�m٠�>	e�̩I �f�Y�^t�%u�W/9Q�ݔ�Y�g���e1l�3{�_eIH��v�p�Թln.�����p�֊ͻ�w;�@�Yz�
BD�����~��L�����x0J/�s3�b3�v�M���>d�o6��n5	���Z�ت0�f�����	/oc��Hf5���A�X���L�C$�攄�ڇ�+D_,F�RA'�l��I$��~0I B���Y[��͠�t.�	�)�c�t��̥X�@�����2�ڮ{<r���{�^�5ѷ��l7爷Y�&���I
�.�*�۶<���μ�T�jI��S��PkZ����y"O��u�V�$�z>�bI��3��+>7a|�F �I9s�&Bj�Z�vz�u����A$5�� �RIN�H�@3;���ެ��c�E"����E���ve�\�8)^tJ�a�7MIMc)S62��0�F�h�d�#Vڄ;�d�I`�û˞ڦY �J���$^IOuH�	��+����	�~�)$�[��%�G��L���fuUIe�D�I>�6��Nl��x�� }���$�H)�2��Z"s��]ټė�L1�3�,���)y�~.`_����\�%�+��ɒ�%0�r�=�%��\�Ix)�%+y���LC&r��.�Gg<�Y[�P�8����O-& �	$������|��s��1R;6f`�k�$��sx�8��gDL�^��%QY H2�H��	�f�������Ira$�T�&B@/�ȒOb��ˊ`�6;�K�gRi�U��+�F�$=��:��cŶ<�Xg�V��.��r-������3W=�Q�M9�5���@)�����%�פ������~X}�"#1��v��j�eJp3X�8���Ii��u3T� h�3pʪ��$aY�n�M�a&Y`$�����Z�a[NE��Ɍ�X�A�`ئ�U��c\�\�KzU�D#�SfĚ^4�f�W���k3ѥn���(G��X��[�e�`M4�`$� م��e��u�l(Ŏl��E1.�Ԇ�$��H��]�A4�J� �����&�򴠹,���KK�ˍnh��r�-P65���,��W5g��~S�3��vwe���p�b�HK6�\Q�PJ����@*��e�����hB($��:�L����Pkp�;�Pwa�@��:�	��^�N�0���fD���I%Uu"��V�dI�$�����2y�Y,�\�^#�C�,�왝P^K/�HI%���!$�̌���53�];0ϾFI ���H� ��}e%tʩ�y��d�]�B����$��m�bF����t�	]nă+�$���K�|�2��K�������d�U1r&Rh�%c�A�fr�����q�	I�f�ki�B�&x5�2�y���HtoH�@"V]lI&RK���)�BF~?�̣K�X�l��b�fŅB�+[B��٪�҅ReqY�nO??g��!�q�����xD�fe�|�e$���c�H�j����nf����z�:�&�I�ؓ) �a8�;:gwvU�TqzA9$-փ����6<\��ݭؗ��������3�x��+)�3���l�~�}��x�S��[��Kr�mr
;�g�`�	�֣Z�DEB_<�����kR��I��I$���($���f:
�w�{)���S�%N`�sF�i ��\}�I$D<M1V��;Na�^I�ؓ#<��H�7��j�n�tœ;33���釨�ٗ%�l����I�)��I%��^ �K�J�շ6/!Gb�Ny��$� ���N�;���ѯ� |�H%�7���@�yNY4=�}p%�fc�qߌB7�nWL�M|Dƿc����8�-ÁiK�dS^mu�*!k��,)�uYm�-��3:����ﺠ�9fl�>cd�ޖ`K�������Co�[�g�NN3��h���[�z�*|�I$��z�c���_œ;R霁pά��`z ��t`d�H$����I��(��К��u+E�o	�Y��;���TsяBI!~f>��q�	!uWQ�W9HL+���׶nd�k8�u��=�`�FKd��^��Q"b�:��#j#(!0W�h[�=Z�>�y�q9�ݚ��L~4����UQr�H��7c�[����K��$�w����N�;���x��U��kk1 %�J���JI%�]_m�V�{.�AV�S)�G,�f�;2uU^J�^�JH%���>I�׉Ȕ�1D�^�&5)	%��fe��x2��%�g�aRg�e���5�����7f��R���F�A�[fm�6R�t2:\�E���D��s��y݃'d��s�1�����K3�)A#�R�q&R�n3o�s���cЀ+�%Y�D2��M̐pY��j��~�y����$�a�����j.H]��bUy���{M$@-��Cbn���BW�����Bd��}MA.�}�)A%��x �L�7���V�c�D�p9�NQJ���f�Y�@P�ˉ2�i:�;:wwvW ݄��q6�
5��OT�HR�A%9��F��32w������s6�}�����7* g���U�N@��u���K��77�6(}O�Fݣ7�oVn{��M���q���_��)�Z�Z�EEG�U�2�� ʋgD����\�S̫`�7��B��ι��93ᵱ&g�$@e�D�I��߉�Cs�ɤ����{�&á��e :7u"@.搔ҩk(��a�Q�܎�h���/���>Y�"����u��	��s%$�%��@LÞ�\�m��`)̋2%��x2��=�v��;���c�D�h(�vu�T�I.�ǂ} �N�;x�$���呯n�g���&X�0t�}F��̀�y%,ݭ�̄�]�d[\�9�h3�t�`4�pc��	 �������ʲ_��'L�e�т��W:��G�Ou7D�%��m��$�AW?Rx�+:��������Z��sI���ӻ���T�ތBA(�[m�M7Qb_1��$#��ZRI�؇�@�Р/.]�QqOq��15�U!��̻�3 �V������#�Y�ga�����=|{|N���Қ,�4���;={b0��~��e=��R��	�y�魏c���X`�އ�=s��p���v����%x`˨j��{��7�\<.q׽y�W�{�Ws�|�U�E��u��o������V����c��y�h��߻בk繫�eҡ�y��.���-P-�o�D���ݽ�W�7y�{}��moap"�;��t���|�����k'=坰^�}]��*_g{O�7"c9��V�����A3f�f�-�F��oz����K����v��n�(�/\>�j����p{ݭ�IV;��h�˓�zw��Yy��c�=��O{w��u��[�v#�5����cm<C�"���l��Zm���r���v�"��=�{��8e�ԁk�x��ﶱ�/z��8�[r���N|z�M8������=�W�c���c�@l3���a,�k���hb��[�;�Vo<�"䛾9���&G&J_<ǵx[�黆�w�ڝ�ǲn��c�v��[��N���	0>��I��8�S3m^�}u����~�o��S.Ѽ΅�H�ݳxt�6�n�"�Q}�h�N��p���+~��ϸys���?<\�
"&����;�2����w:�}�e�:wC�2�oZq� X�DJ;�K}�n�ټ/�����6�,�ܺAɦq��Sj�&�\0���=<��9s�ez�x����Z��aվ1г�`w$�IVO��N�"�4��4�Ǝ������Ȥ�����0�[N9~�Y�D�;��y��	$�=<�����Ƿq���~������J*H#�J����䢣����n�#��Jp�������Ƿq�{z|{n����?�a�񷚇%�Qe�ADQ�w�{Y���H�"S��ӻ;���;���#���ԫ"(#����]��G �}��9�:9��')�Z��O�8�m�8.N�g'q�Ev>Z�G�vevۍ(��γm�9�u�o?�vt�i��qA�^V��Drp$����9�I�h���=�܄��u�O�Yga�i'sm� IzC���c���e� ��V�2�ט.eY�@��G3
j�Q�ћ���F&�����-��h�fѲ����&)��B\�% 31��k�P�f�n�XS5�aYFh�
��vs-���6#-��T�ɥ����\eMm,˥�i���*4�2J�e��*M�]��[E���ʦ�Ja%+�e%�+`B��FӁأ��%�Kh`��iL�CjUu�Ld&���e	�e�B�;F�(�+��h���W�΍�MK[w����R�6`� M),�dɛeb&ˁK���PjieU��BiR��N&���U���,�nm�E�B&��q ���K�ƚ/]H�\����a$hJQ&|�d�8���f:\��/T)j��QAlMe�Q����3153E&���,���3�ډree��h�9ViaE,�ĖӲ��i�fdM���T�X�33q�GBl��5H�e��2�K��f֘������S1���n�V��B����tx�gQ�,�!V�,*�6��� ���jkm5�.�E:;��ˉ.��T�X2��Ĉi,G�BգnNɨ�����%��e�Yg1&�5�/a�e�$���5D�v�55�<\J�R���CD��N�-�^�1���T�;��F�-Y��n�Ҭ`�X� (6��nv.�Z8l2��:	��ݕu15È��3(׳��걎��9Ynba�����@6����ǖ3�Q:0��O.�žv�FWl,���mp��Ѵ�n����K.\�P���f��rK��ڻd��J36�
�챷�K�)m��D V �@�!N9�U�R�� ������X�c"����Kr3�6��%^�)����1�%�	4v e×Ki�(V�4)2�Xk����S�*WL����hRY�1�iYH�fֳf٘���ˠ6�r]����vJ�Y��S��1�q*6���/l�5�63�*�ר�.F,@�jf�,��C����Y\WR�S^2�m4�c�Ο��u���$	���!???,�%�j+�����s`��ڱ���I�7b�)A��]\M��*M�v�re���E2F��I���&�`�F��3W��,.� �R�7����*m��Áʘ͙��쉘8�J`�Ki3L��[ب*��qfؗl,9�e���@&&:�Q�Ȥ�Mj�lŹI����8i�B�]6��m���cG���(���KT��:(�fPf�M��h�CG	 �,vԲ��\�3�Ku�b#k3�������?�\��c}�&�$Y=|D��P��/�Gud�$�{:}i�%�C�L�p��2WE�����u�3�:n6��$���O��n���4p�&��K��_�;Hם�;�fwuT�z ����j� ���#�ų���~����I��G�[�YD�E���:e3���`���� �]8�l]J<H;��-���{+��zIr����/�r�v(H}M����gdH1���L� ��<	��u( ��;&@&�iXa�e�j �rΘ�,�Z7��%��&v��Iu7d[�ƗS8���GMl/ϡxN�NΝ�ݗ�|��"U���//"Hξɒf$T�Κמ�7�/�k�����ZE��(:y���S �:�l.'���w���쫶Msy��K!���C�F����4�I
����}����8G�GbIx*l�7�)ɶ^�8�=��$^��A�h��(B<�G�A$/������&|O��f�k�zi���۞�>j䶈N���NL���`|��D�H��w�����0��J>'��$��E�=�vr�;����7XC��d�j��֯��|I;��2 ��p�P�����,t�#��pSL�D�tl� ��؋5v�dTSt( ���$���s��\t�6w���ָ�e�*B��]��]s�Yi�:j�W[�W#�x��X]â9N���zQ��w��$��DWZ̮���v��:�2gĀ�����vggJ��.���	�+���T}W�A�/#U�3^�������v�`�V�hl�ք3�W��["��<�n���H�ʈ�E��l̜9��,c�s{R��__{�,�^w�����B^��?��yw����?����D���i>>�-��;'�7;�����˶��Y �e�������x�ڈ%vnH�A�����t��N�Y�'�M��.�awX��O�&�z B ����-�l��wE^�1ӑ ���l9vr�;��=�� o�\ۈ��;�``'�+&I$����֠{/��D0�����S��~�� �uG�&���I�1��h�c�r@�hZ��,����GJO���mQ�јtGw����$sg`ĉ��P
Z2n�aOP�򈎙���؃��]�tCyӳ;�Ҳ��q��l�fղ�=���cA���� ���B
܊�o�G��cGu�X�'`�E݋�;:S�[/dV�����I�}�K:�|B��z������	����e�vtJ�P玹0Ƽ���^�$ר�I#���vu���Ͻ�g${�z��v2�*ɼ��'w7���TJK�z����i���-^g��@#�ќx�V�E���?u��|?|��4L5Hr�B�����0���VjƤ�fIé��ـē}�p.Z"i����#����J����㥳���Tlo�s��L�a^T�Yi4��ڸ0R�3KV��.[+wQ����b����?��$����1��s%�s�9�I��8��	������U���0t�g�ջ2IS��i��T��'�?�@�k����q ��j��Ҳ]9��Ȃ䇞"�âΝ����6��vv�z@.��n^�ܞ!2`j��|H&���^G���Lz0��qv.̝ʐ|yl���s�nax�"�W@bH3]� u���ۖ� ���7(=���e��w%O:��,�@^5���W�qݥ�����P;ݗ3(#�=>��-�]�ߺa�Bhk"zF:�J�����G,V�f�6�k//�g���V�GBs����֘�{�:"Y����ô\Px��
)�n��|@�����<�	��.��I�	�UѷK0�$���Y��`�m�a,%+l�Vhl�����4D�Q�G�H�"[�R���:��2��P�K
7&H�1eLih�1��с�)[6�1�mM6\TՔ�HF�͍�J�-�%B:�tWfL���mTSa�
��k��h٢�M��S[.\M�@�-���V6-�-�D(�R+� �2��
颖�ĺ⦌�Z�4<<][l��întRؒ�2U�n�M��³�l҉6ָھ�}~��R��8u߀f�� ��}{q$�	q� ���$B�\��}P	���L=�:��E�;2��b�Zr�cU���g&�bA��sȪ$H;�� �9�n��0y{�ZH[E*�	��S!��fA$����H=���m�>�鷞Q$=y�PH�$3r�	���瀳�p��gvS ��{�x/��<H)�$��(v��!�n�B����f�NH'ٙ�3�HG�p���;r�ڲn3�X��4�i�Z�nH���	�>��.�9��6�޷j�vwL�I�dJ�aY���#jM7���١Y����H����_�c�L+�.>�c�L�_�k'�A'���R�茓z���=���2c�"��Ǚ���$]�L�8u��� 1�\r�B8*{ipP�?)s�Kn���k{�Ǩ��c��_vN��z��|2�;t;ӆ�:g_k,�f������|��P �x����x����@=K�G�>=��3�1�{�C�B8�� �:e2_'� >�*�jk��lZ{cr�J�Y��]c��	 �o'\A#m��;E.�Ɉp�:u�v{.�>DXŘ��j�I>�qm��N����f���֢�@���k��࿛Ν��@�8����>$�ۃ��Sl�]�JB8y\̒Ncm(� H��~��I����ޫ?1jF�`Q�f�,#*�V�fDՀ�jA��uL�a�!Z��B��{��T�
_�x��x�o��>$��om̓3c��P.����k���1���ˢ��B�$�LwF�����	&����_ݽ�I�ݱ���J��{�&��&LJf)æ&qu($�^�H�NT�^�z�_���gJ��R΢��/��f�g4��/lW�i�RT	���;���zxo�#���_eYݾ�>c'�e�-�������>����@�Y��$;�%�a������%��(��TvmwC�S�Na>7K� O��Hwf�P'�yy���:<X��*Ó+:�@R)b���L:��=n̓�A�ُA��Kq�^�$
O���*���H#��b-��	����뼧����.[�P�t��a5�J��Ph�ݣ����G��<�?����.�O�Jz��I�7��I$����(�����sdB��	���T�2�L�w-O4��=2Fgf1��L��c�I$���Ǡ�ј�����;Q-5��;��ܺ,�qk� �Θ;b^x>�1���xj� �n\O�%yu����ηE�0L�p�����o�ϋ��F֠	)�:$Aom�D	�]Mu�;�����pqV�ހ�Y���t1��N����"��&�c>^&�Yz7t�H|wQ�-�)�/��v{��٦�k��y8����-����xq!碦C(C�Xr����H�j x�T=@�{��z�� f�:'�[�����>�]M�!�����ԫ>��:�l`El�i�1V���e��%+V���!��`�ȱr��V�3tSN��+�d���x �U��⩢Ud��}�3	$�t���8s�!��3�P&�<j�<����v|�ڙ���A���x�yWS@+�z͋��.�4��Kş�3L��ZD�i��L�Qι	��K��KB�lgS�>�$�����]M�ֆ4�r�y���SSi�c��bMtc�>8j��e������R�0�؂�oiٓ��'i�'�aω7׶ �H�:˺u���Hn��N+zh$��s^5�u�ry�f�զ����Vy�c�4~Oiez*�$�s��=:������ӏ�ͩ��&����޿	�;���t�t�0t�Q5�������f>^�����eY��K��e��R��4���Wl�����aF�R�Pr���ƁKΚ�m��R�j�.�en�����0Cf���]��� �R��G���[k�ĉR���W6Xۋ&#tTDT[����
k��L�e`Fa�p�[��d0L&%G+���L�׋[l��i��ٌfe����s�b��dI��-�ɯx�F��>��Ծkn�p�`fJ�B;:��Zr��vo*�*Jm���k��×w�gL���O�9�nA ��oe���dU[K�yυ�=�Q ��Yt�+E�V�:)��S>n��j�e�\d�w�Q#�j���we�ϒ���k?a�n5�[�[;a��.��)���!� �v�H ��
Zͷ�˧��/o=�L����@%��&E�w-"O4���ܵ��ȋ^$uؼ}}�S��N�N�2�w�ў���@�EOk)�.�d�A�������|k:b"���\�U�b@�>�R���O�_LF;ԃwn5�y��E���ôU��\Yp٥��{q��љ��`m	���1exلca?~�V)�fAس��P�Ě�ˉ���D�
�M�z��Ҡ�D`��q3�b�.�	,ΙD�Ψ6�Gu�Ź/�D�CEod/}BE��|����`U]^҄3=�h�:���K��E��LD��}.��rfhe���>�y�y�I ��ۙ� 痗������ژ���.F�V�:)��N;��c|O��j"<F�JX�)�l
��s��	'ս�7�D�{:��6ࣘ�bAt��8�����̼���P�B@-y�A"A>�k� �x��DIIWs`�;�/�4�2	8�'0$�8`��P�4�z��u@w��4��؁��ؐI&�j=�]M �vȗݢԡ�����*rɒ��r�����m!�!x��.N���!����/	�!�`.]�$Y����ɒA�1��U���1U�B��.�ِ}w���;bɈv,��9���o]�S���F'��H$�ޘ�I�����4�/P# �򜨆}>����r�����/�Pt�e�#ǻ	��N���ft�D�]]�U(4�B|:�x��J%��qf���R�Ch���f�%���}�Q1�̉��dԳ����|��<}3�<�Y��I�v��%�J�9��>�Ҟ�ܻ���w������yyz[��o�A��{i�w��WuKQK^���v��<l�a��C �_�=T�-wǝ�pɊ1wm����ϩ�e�=x�n�����X�q1�Og��L���Y���}����R�}�lݼM7m������V�x��[� t]�KɎ�4�m$u��2\^�.{�3�/�C��;��5%��C��V%�wO�MQar�f��Qlc�yȼs|�'ڦ�z|���a�ōoP���&i��O<���2g���������}�}˂����[��O��ٵ
�X��wsS^v6��`Gب*'�aW�oAM��J�q��x�� TH)�D�u��LgU��py����Us���Wu��������D��sp�z�P/ w�%�6:�t��`w�NXHQ������ǌ{|�+�)�0[�tK���˝�_\��8g�����^���x{ҟ, ��}��7L�r~�qbvVo�6!�I����|6s>��}
�{7S��-�{��9d�D}��P_��׻��i~�N>s�n��A�u��� ܫ�&x�/.��J�d`�^��b�]���(׳�U�&ǽ��+/��ł�X^�}����^�\�T�g�\�{���CuY��T{�'#�������wv�i~�]b���.�`N������|Y�~;��f��Y+;���hRT�I���XL��YɍSq�QyL`|ό��t�޳5�־�Y&��'r���o\CE������- �'��n�q����q�2��w�R��\�d� QG���ӭ(�|j����@�^�q����q�q�����v"ۓ��*�m�j��$s���㏎=���q��ޛ`HȒ,�!$a�b�Y�Y�k��.;mm���M�r��r�n	�;K)�R\֬���s����D�>-D��߮Z�gNq@���(��%��A���'�_�^����Ƈ��՞Vqԑf�����͹f������g��O6�n[V�f�:���KkB���ٵ�l�N6�]�Ͷ��� ���;�������8�;�m�{�qDI�;��Qee�dm��'�Kf�+��&���9��$�X����$��Q�>U�4�Z�a�3��s2|ݷ�ӵ�s	=� �H�M �Fu��;�bhuy�NC�DA���$�gb�a���H=�� �1X�le�'s� �O�[�@i �\���catA�u����'ww!�ve�G��Ius��B��.��ۦ���D5������5��b�0N�P'ˎ�l�	|�+�bI#:��AٺJ�7�\d���	 M�R��@dhēX,]�$Y�y��d���U��ˆV��H�	�e5ҏH���B�x�8x�3���Q5�鼲�3d�ӻU��`1$�̉��wϹ�fS7I��0�y�|�w��.�ٞj'č��%�]ܐS9e!�f�����}W۾$e� 1&��>@�I��q�i�u3��H�4����f$�{`�ܪ1|�������0��幺i~=/��!g�ʥ㫸s�iX�Z�S۾S�w������$I$>I�k緐�}���سt��P���d	�y|��GS�Wq:b�6����v߮d㟻��lc�C��	�a�v҈CQ�Z���B�%-�
��ev�D�ګ�f���n��L�ɸ3��坊��N�bIܾ��I=������uD���V)u�@�v�I!�hŀ�ჳ�� �N@���)��tv�Ȅ�`1$w�.dH;}Q�?�������r���0rd�wIy��1dgT �!�U3'�Ǫ9�'�r�H#o��r�.��L��wh�':x.�ͨ�7���Gj��I �H�� �O�Z��;ND�tfa�Y�	��V̗��u˗rC&r�H/�Q�x�Tj�f���Ʃ����TWd	�����Mx�93�Ey{v�����B�v�I�}nog�ޖ�h�=/��I�/u~EO��L'=����gy�E�Is�ܺ�jVg��n>K}�vR	��5��<�9(�~>��jV	������Sk

�5�6�p��Z�V%f�6��D�;��K�5aqr]�jˬjW]&D(���J��1L���B��WdQ;M� ]��.JS,l��:�nL��X⦶�ZK�[�ט�"jh��:P���KA��[����i�DT&�^�[-����WCK��Su���h�2h���A��飙��쥛#*܆ƚK��c6ԢK�K�@�P�h��e���Ɂ�Yf�u���SjԵ���*L](m`Bvf`�ϟ��fI��w$O�� ٹ�$����<H�]M ����WV��U2I'�. �^���9,.]�*�x��9GskJ!��撡�1��sbA��O�������ժ�pg&��%��Հ�d�gM"A杁 ��P��\��h�hzy׾y���>#7. }���<��a�ˢ��"��ꛌ#X*o9�iC�(��O�纁�mm�@ �w\�������N��۱�����n���L��wi�'na�"���A�u�%;�;tO6lA$�R�I]�3��+�e�ߚy�s�]]-˻2�@���KpMP�\�6ۚ�֙��6���G� �/��&�nGP�����7T1$�o\I6sk��V�:��U��nUc�([l(��erf,�̀۷� ��UI�;��DE�����x\D����佧�݋�,g�{~�x=~��GN�^�VG�)�,�fi�;�������s��>6����$��y�̄��uy$	���$͹�UY��ޚ���l0v%Aݒ�eN@c�|VuĂA ͹�yri^-n��I O6R�A#k��A!����X2p����><ӭg����t�Mk�̒@ ��W
�؆L���Kv��z
�S�E��E�d?��T� �η���C��3n��M���	W�2{�"{�;��!4���x�;8w,��f8Ъ��Ո�l��t�hH)]���-�6]
ٖl��������%��2wg|V�c�A ��\O� �����6���9�Z�I��e��S&0�.�L�(�ۨ���j�t;�5NE�.}AN^�� �	���s�3"/62$9v�Bd`{��Y3�;�����$�ݨ��ynfv��A�T�<�����𣄟O�f�2z��*ӷ��'�_]��ԏ����;.[ܷ��<{=.ŇQ��v���O�xyg�b��g�����C���K�}������?^S�h|Y��pPt�(G�V������B+�D�ي����#:�I&i���<�-��MǝWutω�x��[AA�����P)���AJ�/�$&�ِH y�	=Mԣ��p�0b;&\O�m��K���h�j;\[x4E��3�KsR9��r�`n�..�&gE}�[F��$�kv�<H'���%�e=��eϙ3�A>;�Qc���9,����!2gTp���vZΝ�~����ވ�A#������0fL6��(C��C�}-a�8,S9JCoPqg�e@c�qS�f���i�i݆�9���@#���� ���R�����wR�kaOwZ�5����#)��x����6�dײl���jbm)W=9=XT�*-�)E��x*�k(��Z�bHL��)�W��o����n��?i���xKu��*�w/i��eswJ���o�b��g���k/��9('.씌�a��D���x���_;�kn5�H=�iG� ��}r�_Kr*xNQ�.lJ%3�!���,���(+�f]Z\�#��Ҷ���,.��k�[�v�{�ɜ�� �]���z	>3��c����~n���S-��36G��� ���l5��̝�,�K��D��
��F���x��e�(|J�z0$}]��d�y�+�,(oZ���l`䳻N��ƛcȂ@�r�H$�⌽��[��͂���p�I<��2	%�d�1L�)�Y5�bi��1nq� �C\"I7w�3�A}YF �s��32j�M������Q�,��ݐ��;z�d��x��>�>m;�c[�@o=��{s$ϒ��뀠���:��f�%<(�b��lygl>u&�n�۬�y_�p��2��,QE6SSal=�!�xg��}��v�E�����ٹ9�
$0�>l�����0��X���ݗ�.�1(��]mE0Z�n�3aR�Rlۍ�(l�]v0:\FB��4�r���;�Q����踃Z5l�Am��]2]�/L�l��k���+����,� HR���R���8@�<�*ɂ�nT�dZ�1t41�3�wm�B���	���L��J���;1�Z�س9�&�hL��Xk����Z�Ժb���\��C9���,�h­��,����ˑƱ�<�����P�9wd��̶G�8�^�I�6��<v���m*j��췠�ܙ�Cn�&�Pvp��v�'�r=r��"��Ti��4G�2�I'o�{,�)����hi-�d�H�jg)�;Yȝ׆��I���/!�L��n�^�W6q�I�칟I��y�?nH)˒��
wS �sN�]��Z�/�;�h$ی� ��P$smDx�H��n1���=T���=Q �}-��8L�;$�d��@�#�Z�d]��Ȼ����*�E�H=�O�\�`�l�Fo�N���:n��K�Ta�����K�!Cv��C7Ee�	��z�����'�5�fE�>�ͽ�{v��%���F|pH�'8���S�a�e�p�Wa�r�N]�(�ze�<����+Ɇٮ�x1s����r:��K�ɼ~��������$<����ye���?a��-��<�!9��?{ӂ&ޮ�����@��F7����|@,ڎ �'{�����F	�]ݮ�]?���<��ƹ��(;8A�;C����9�P�n��sW(���k6�@>$ms�o��jg)�;Y�GC�L��]N��6w`SWo>$�Zz"@$umt���3�Я|H4�� �v�,��vv	;����9��I��Ȑ���C���q�2A>�͈$U�D�G���d��}�l�?#징�c�;Z4��t��R��FS�&me�Չ��ٱIv�|�����W!��Ym83�G���g��d�q�W�c�`��@��z1�g��\Ƞ��9wj�O׳ ���w4�D՞�z��<�Dx�;��$��a��z{��N�ܤ�"���S �Kd#�L�vDג$���:%:!�1E��ng��(K���˦>�v��jW�����9z�-�y-�F�|GWh99O>#Sv^��{m�����=�u���A>ͷ����"q�c[8H;8A�;JA��T��j-l��)�� �g{rCzQ=}t͵��*;8AS�f#���.�]�;$�vjd�k:� �̘i��h0	��ݓ �o�K�9�̺�e�Y�2o:N��;ɕ�I��=n��Kk��D�����׍�l��8��VV��g`�������"I����z����h�w5�\���H$wnd�$lH��Ӱb���"_қ:�-��]d�3�����$�����_d@'Y�E��,�z���,�s"�:,�ݜ?���{��@$�W��)�����K`9��7�HۙI}n}��tS�$�;�Q~1����\�N]��$�|On�A	�z%{f�:t���f��	�w|����V��&]�*�rԢf�9Ea�Y�6�n�kj����u�S�/=ܨ�� A�_
�v63�� �O��zd��c��A����g؂��W:0f�t�Z��EO^H�H�#�w��V��I=������~K.������3l�l�KE,�-�#w:Rj$)�	I��K�~�ë�b�}��s��x����	&���7QNo���{7�$�|r��An�
�,��wS �.�|pN���稒|H&��#ē��z06l�e�s��.g���e���씅�WR��Ez�5'�m�8l�=]�	�'3.=���k�S��L�ݥgV�ɾ�]�6��m���U��	���Deo?��Jქ�1k�g��I�و24�[���$靊�1����w/�'ŷ;�2zZ�`�H4F�Au�H$o_d�8��PG{�7�O�~�o�<4E�?n��+	�͚��L܊�zqʙa�ٻŔ�b�Vc:�\��m���Fz��^�{���ُ�tɫq������=�]K7����Cr�-Q�<��G�{<�V\���㞎�`�xw�b�K0	9�K�D����hR����WO�1*��X�
��C��i�҆w���!r;i�_v���ڽ��+�&9���;�^���2���� o���!�]��9坢t���~cu���PO�rZ���Y;j�|��E�8OxE��8�����3������-�ynCj'��;���I��ˀ�,�3v�3$�%S+փ�T�L�Rm�Ǽ��{ďW���n���k�ׄ��L�|?5�ӟ�K���U������⛣�G�8W�3���:��˵������A�n8Tyx�;�9�}���J��Ʉ��aJ��`^��=U>֙�d�L-Y�h���/�rg}�F8�c,ʰF�MԼɗ3q���Bw��W������	��[�]�I���
������I�a���<�Ӓsgڂ/����uL�@�z��g(�������zy���ǀ�z�˻Ϻ���I��9ޔ9td^YÏ��n�CT�{JL���N9̋Z�wtsٍUs%���l�B�[�L�j#f���QsQ�C�̋���)�݆{��9��hl8����}
��*3�{<��=��{��ש�N����o�]���]|�^��g?�{<A��}ׁ�3}�����(�m���n�����|V��JՇ�pdI_/��=���h�'vy�#I-��=�x��_1����F =�����Ǟ1�~ t��Yl�����7m�:mY�l�;�����==>8����_q�{{��oۼ������ㄭ����l���*�z�{n@��N���;|v����|t��8���г�H!u����֩Ji#�����m�6j����u�͇M��#�(���z�ĎD���R�q1m߷��Xqpۣ��̾/O4�L�;lۈ:�+;mfVX�ل��,HC�B.mbSkN���ŭ��nPvVnYɥf��km6���&Y�n3qȓv�"�٧i6&:�?:����%m��M�������l�n�ۙ�Fno�w�9$?�s��r��ݷ���{�v`8�ޭs;�{����ז���͙r,�&���l,��M4If���Ȗsn�snlM��6�#��a9���ge�k�/�E�݋;rNN��]�������4+.����:��Ү�iR��6hE��ˢ��Dl&���j�q�V�ԚցfьD�-6΄�cz�#3eIJ�=���w�%֎�1��F��.��Zg�l%̲�����Y^%SkY��6���9�H&xC���2Fm��/�(�b֯ZL��<%��cBn��%[湳[��#%�J��qCJheu�Y�1R�"mR4m�i����3WC�6� ,\�v�is�5n��5o6�ȋ]�Kf�eb��g��,�]3�sW2i���
.M1D��B���WS\4mŔ)+`�l+�f�ccnm۫Hgh�v���	�[��GD�;-�m�V[�ְ.��oSm��jW�.[M�l�nB�!�䕻��x��R`@�����%.���0�Źy\hl:��Wi�.�a,у����-p�!����KY��v�٘P�Ȋ6��ta��!�"�!BV��b�+ժ�X0�7B�d�]l����*y5�	�,�5l� jJQ�2Yfj�6e*<ڕ�e`��Rd�;��cF�2�\ܴ�så��٫	�I�Iz�b�ʙ�e�\��ݹ�]+TA�!j\��VK-�2���7:�I�Ku�V�H�������Tt3i�D&��s\-ζ*(Mʙ��hM-��"�*.��K�3LP���rc��G1���)%�Ap�i����@j�C�hd\��YLڳB�b�n	��z킕O-�k�-���![k4�<ifƼ���jK�Y�������+�ni5���f�[s���d����00͸c��,�J�6fd��$حi�бV�l1�:�hL:��:�Z�,)dcZ"�%v*2�r��5��]1�5�Ե���u#���aH
;�v3�H����l��Sk�&t|�@��*��a5�,Mu���u�2@���`���f8�t�B����lKV]�����Z�[CFMT��a5�
��غ�I盷��)D�ْ<l�f�+�w����߲y�Hq���o5��
e�69L����15�)ٟ�-<�]���T�V��pk�kn�6U�,��Di�C�U���L�[��������F�
Cq
T�6��&E��4X�U�b�Wk��V��l����k�`�c�h]�sE���4�51uԳF:�Dj2ݴ���lX�@��.�R�ևU95˴M���y��Te�ɬ#��$\�b��]�n���T�����=m���n�g<�D��ؙqe��ڗq�9�J��V"a�3y��Wϟr�vp�������"k��A��2W�"�o\Z���ށ ��oF�+��-�9gd���ު	��d	�`��g�M���EW=��k�D�Zj��E�:���[4��˳;"�Ԍ�h�@$W�̻s"�oĂ�]�B�/h֯m��I &����� t����`�]D���Ϲ��.�{x@-���	���2	$�����Ҹ6�'���t��0wu26�dO�n��l���h�g���`�	��ɒ|H=}^x�>��V��������aF��k��R\��b!��)U��-eW��}?~�i������n����)܌��>S���*Tnl�϶�~" �$7�w�v��wE����yC�z	��Zy����?���o�d~��> �1�@��ú!����Z��(�&-�T���I�0��nR�/=�dzk�t~W��R�<Cw$<�$`�H��5�����3r�A_�������K!��o�x{�qҁGQ��I���@>�}�[�S05�K#d���:���@��ɐH9���x�
�쓤��>9<�UH���q�J뉉�%�H$n��I��b�������UD\�>��:vX3�U��	��
����.�a�����d�|�5y1 ��==w}��ۯ7��o��~�ե���f��۬,ҌųWjT���nnj����Z�o'���>��4���`̇�L�����;!����<�^��x�A&�&o���2fE��;�,"[������T����=dϫ:�������%�S��z"�|�K����.�S�]�I�{� ���P�'TXn�0��i�Z￝�I�<� s�.�|�t7cA�<��-:D�De����t#%�ZVAOv&��Nk������<9$�C<i$���{}\��a�]�g,����z�'���j�A ��D>H�5��}ՙ�M/�p�(1笈-�pP^wd�$�@9<�Mv�D��l׍�f�w.�7e����@$��Q�;��$�eF�;Q�$$�%c5&p��) ��Ņ�kEԔ�an!3�gd�0FK�&��L��?>��;�8b�9e!�+�	7�����x��m�Ua�*����<Ǡ��F��'S`wP�kc	-Mӑo���n��������e��p�8:{��� 3�~�b�Qd���L��l0>��!�D��";�	n�v�dMg=$#���� o�V�wE�;�r�	=/�V��p�{�x�\ ��5�>nԒH=�L3�>�I��^w��&U�(R�p��.���Sヷv�@����߼N��7�j;O=�/��{|[z�K5@V�F��>>  Č�|0Np��Y�wA�*�4uL�I��=��kyh�s�ыAz�sf|JC�)б���"�־�$x�V���â�,�Ŋb�5��R��D��e��?��w�.���o�>�>��K˭�}�}Z��א$�_Sǋ��s�.����=�v��I-:�bvv/��)�ϝn&GC���vܻ�k�A ��H8g����L@>9���F�i�g��$�CP�L�'t�;��l끄�۳�(��;�p��-�t��u>D�A>;}.�qS�H�B%���нޟ����s?�*$	���x��E�'������#�9�b�����KN��(`K��i����<j���u�B�k..�j̹�O�=�1 ���F�5�����7�d)���'�'�`a������NՌ�7}��8L��n����Ѻ}�,�q�2Ξ�Qwc���:A&���||��(��񩡒\��UBn&+���5lW]pW����vH*۵��h�h�ڵ���V�h����bS-a�Fչ��'-�0Ō��B:[]�֚;�Mx��:e��%���ql�ZDP��vo66�aƶ���aZ ´���I���ؕ3�Hۥ�ĥ.�	�H���"`�&rGEc��&@mSKX$ q{D��3��Pe?<�y)X���IA�ш�J�)�qiH�#�7F�lL=tl�����<��Ҵ',܄�G����'<��LA䊾j0w���w�3Tm��"I=�1k��Ayݒú�����i�V5�V�^ta$��oTI>$v[т/�+�b�%�lcN)V����p�d�u�A�ƨ	�G%pkb�kr�-
'pI�& �W��� ��V�$�ܧ�G>nI]ݛK� rb�7�M�D@'�o���_c8�*��	1�Q�{ȳ��أ�ve�$�Ή��hM~����=��U�F<I;�]2U2��{|v禺j���Ѳ�
�c�jE�&�)��c�:L���B�v�f�����[�)����|I���	�]2	~�+Lj�f�R����
�{0l?JV��	סkGE�A������D�m��O(HI��B��ၽ�z���׷��{�c�w���{�L�9>��+�z��.ﯾ���0x���[+�eg�a>Y�"Nw��?�����ێ��|O�u��$�뮙�&cԏ^�n���\���.�ό�4��^�D��>�V����E�n����Ou�L�C�);�Dp�g���b���C�;G:��`����6/kH�EwZ���J5�������&��fI���gd�y�rd�x�ڈ�-���Q����>͏�Hy��+����I���v0m�ɺ��?�CY�hӀ�N��uL��P�D���3CAlݡ6�sk�������`Ƴ.k�~D5��$ˮ���oTH94�q�tܵG���>�${�r%��Ӻd�ðr]��͗>��<��G<�l�01	�ܙ�{�-��0ܬٵ}pߍ�K�r���!<J��$e�<xyăծ2%��m	1�Q*�%�c"�\z]��˯o���a�{��L��k���nO =3������x��ݛ����א�7��>>r�M��̂I5�Q����Eyݒúa"3�WM,�0��A{��Dg���H$O�z�<O�\�qZ�Η�� �^TH�<�<�+.�K���P,lu�A�ָKnflFK6)g��H~�ْI=�P GW=�ه�B�M��i|�C1���%sDe��B���Tɂ�֓@՚�8[��3�@��N��;$��:�dNnT$���f<���sl�q��.�&A nT>�mԆ̃fp�2L6@tA�Ǩgb�ll��	&�* �}DV��FA�Iۖ!����m6'L]:K�W�x��<MW5�D|Cꎋ2K�i���I�tG�Hv;ُ��VĹw�O2�'���Y�[zIy�s�G��wR@�J0�$�'��q�O�ճ�^f]��S5O4��������Q�Յ��n��4W�ް�=�ǲ����g�~�:�]DL��Ĥ�o�p0�M���ü�>>>�Ě옉}[l�����$�i0	��ν��&S^��o��v޸��F޽�$뮍/�*��Y˭f�ȳ��t	X���0�ҍ�9��mzͦ#2K�םDBƮ�B�m��������p�̂��z��5��u�L�XT��� �*������Z�$���3�S^�ɟ'ː0I~�����	��ق|O�t�L�A�m�G�cx?�6�^��Fl�7�;��i������H �WB[Z�l��͐H'���@�|Ol�L�VmbwN��t�i��[Qj[l������k�I%�W7�D�o�z��Pi�#o���c������,K�N��!t�H�Y���+zc}-�@'��wM��$_DFgm�f,K��S�=Z��ɚ��$�Wc�&Ȋ��ҹ{"����:����@��߂�ѱ�#N��7����;M�dłC�>"wO_��$7�6��U4�:�qՕ��t5.�J�f5�c��3\�B��3[p�uZE�mw20�"m��5Yaf�]"��f4����.�Lv��f�^Qq�˰H��Hdkff�&�e
[�:
���L"R�\�e��Z��]�Y�Xf��mkרзT�I��@tX�0K����� M�ie��`�Y��ѵ��7���V��6�{b��:��2���Jp�*�"�Q%�Y�4̺6o߷����v,K�ux�j�"��ؐ}�����v�ogk����u�z����$�U��>=讦(k���2pSI�n�A
���X�"�۷��A�̹�A���jJx�r:�g[3���;�P&��i �۵�q�&��68���#A>�ܹ�H;��j4����8f��[�g�m�~#2���� �͸�zzތm��6%M5�pH������ֻ9t�Ӡ�H����	3��Eʐ�=�I�绔L�� �mD{zڌ�U�蘼Z}������@�i�k�`m�r͠�Ik)���t-���:��j�Rg��}��Kuƙ�;��F�٢/z�A�F{�"̃�z��1ͫY�(^S����L��v!��u3�=�0��¼N"�xT�P��j^�[�_g�u���}��隶�w�]9�Z"+ɶR�RE�1l}���;�*b�V�DK��������ѯ7=�뼧���6z��U��%;'����fH۳�X1pS	����	 �[Q�N)����M4��$����A#�ތ�z�����wŅ�k!�t0���ݢ�?D$���z0�)�ȸWn���H7]p �r8���;8M2o��D{}Q!��2�Q��D�z��Eu����:�E�5�6�wjh�R������F�1��0��2�Ź��e�0�Jm[���%�Tv������?v��j5��}�x���}=�6�-���tȏ3��a5�-����u� d�{�Z%�'r�v#��Q ���=����2��*`�A#;^� I9��2	EN�Q���l���3�}/vԙ:rX�p�A�֘o2'ǯr�H ���Ws�𺹝�;Ԭq�nT\�C[k�~��ntP��}�T����F��|�{���n���/��Q��f���{}�����L��k�s�.��x!�W��=���1L7���#��p���|�7`�ڥ���~�ζsFþ�>P�&	�l*�d�ˍ/iq�g) 8S^!��Ȏ�J�٣��l�����v���"���FnNy6��~�^���y�m�c�G _!���(�ƹ�D֩�|e�#�<ϗ�m�j=<�]�;Ƚ�F�͠��Eت�퇽����?0a�iw{e��u��ܮ��a����}A�b�ƢD(2��_�9u�׏�zܺ����e~>x��?{7��=Su�{��d�闻�Z�on�K�{�gVv�z�'�{.�K�ϩ9����6���wl��t)���k�~o�Fb~3���_��� �x��w-�l�J�q�r�Xm�C�|��2�X;�g���<�j�v?[�ۇ�jC���g�K݁Q�o��:_n��<ˇ�(�(gy��p�rƨ�t��\z��<M<��Z�}U��N�|��^�ݾ{���=�3�7։�A~Z��wO,;����.�x��GKڱ%�y߻}�i���y���%��o� �ِj��:y��]��v�'��2z�W�9�C,���MQ�P6��g�o�y=�Ӻ;��y�⇱,�v:���Q_ ���>�,w,^x��m���x�E>�.6�1o�_B]����亽[��e�
1�+��SR�1�5nHt��,��m�6�"�6Z&v�[h��^��l�[[�c@�YR�M<�|q������O�8�ool��	%�da$�'f6��[2�~���:Dp͹�d
tGє��Xi��n8������Î8����֣'|jMIe�m)$�!!����RIĵ�p�ٶ����#��j9'p�j�sf�lڤ�"@�ok�pt�n�� Y� �����mm��V�Z�j�(�p�	!�������n)֦ͧK;t	5�JN�����6ġ�gy�����d��s���G�gv04	"�k���NO��8��/�E���D��E9g[���D��)Ĕ,�v��֗�P��m��&a�-J&�h�Í�ebKkzk�EΛ�qg2b��m��ƊP(����u!I�2�_�����Bȳl	N/Ɲǵ��	���z�+����6�e����9ӗ~y�";Ăj��������2]9%���/�m��cV��Lz��Y� y{�$�v�����32Q����h@R���ƒ(���}�������PK��T�U�����$�۾�^ �w:�6��Š�Y�42<��y�C��%�f�̆,�Z�!�F�#MZ�B�W�Ͽ���tA��7p1P��oo�$�I ����Y��rZal5�??$�f�E
�۶X�ӗN��ڤ����'���v��{��y3� ���b̙Y�� ��eFi�������X�'%ܸA�etmL�$��>$�����0�N���H@��̙'ĝ�����f�d��`��L��r:k�%L��`C�ED�|h�z�H�n��ro	CM$�b]��t�SsDM�L�S9A�9�
H��BDֺ���vn��L��}��P)���4Itȸ�*ջ\Xig����||x���/7�3�ෙ�Rz��	�*7M[q��O�����I��q �N�R�k����=��<�@Pv���b�)6kI��k*K� K�p� :���mm�{����}��d�]2`;���A ��DO��n�݆���B!�,\�l�$MgT�d��>��]؂��i�c�b��r�C�����Ē	�PA O7R�w�(���;�#G��ޟf�.t�˧^p�"A�|x5��\0ė�x]��<�y�G�*�
ۗH��M�a֫b��N ��y��/r��brΘ�u^�	���?���� ��}��Q}��X�Wx)�"TkS�vpY0p�A�[1�>&|�����=�;�8�Q �5��	ݾɐtc��D	�$���2օ��&�Qa������5�������~��;�MْJ���2S*i�Kw;�j5�ƭ��C���ٵ�`]��w)�.?���l"I����K�Һ�p��X�Q�2��m���4f]��V�h�1��l�ٮ��aoG��M@04Z\,��m�Y�aFYmvj&��n�#�
���5j�a:��b�ƨ�Ց,Ю�(��M�l5&*]A���k3�@j�e&z�+,Z���+��r�RjEB��D%e��f��^ƣ2i�k�d�1X�~O�/����=L��֮�Ɗa1T��SY����,36j�p�d$�^�2�C��g	Y�=�|"��a���z󦑼�� ��D	�}M ��n1�N��˧S!�ofI��vp��gj��m��Wt�A��5�D�5���쩹ݥق�̗)ӱ$�L����rF��D�莞j�y���Hi����%^S@$���"=���c�N]:�j ��ܞ0^�.�D�p Ɓ��sn���ّ �A��ێ�nwÁ���	��˘�rS�D���GT� �Ψ��
t�]��	��s�L�A'�� �ӏ�u̔+*����J5ηA�*$���5���
�Y��e��V���'��W#;�˛]���Ƀ�u�9>�/�2�A��x�3��^�_����xւ��ɐH	�J8�C�D3��A|�'*&@^�q~�?��>���rc�מ���N%�p����]���Z���Aޢ��K/�=vu�܅��������|1ޏ79�C#�u�L���T@$�D6��+����x�u"�(-Z�� �۵�O���npK��T�b�a^9{�	'Ư���&�\�'D���-2���Mc
���ؐA'�j+���{���o.��̒��c�N]:�ɇie� ������2����3��KO@$?�\���O��x�i���#�=�7�
4���t5�=��,ɡf��5�n.�b!{p�ю�tY痯�/���3Zi�]��=���p*[ŋW5r���͍�%��\����H=�o>�v�5�'g��ԕ(�b	}���0o��9�]3�(�H�ہ Ω�#�^
�7��sF��M�G��r�L��2#��	/�4��4� ���fv���"�H�d�S,�SO9Xb�Ό��ѐ[��F�r�x�Nxy��䇲�]�E ���]���7�4�U�ͳ��s��b@�����O��7�p#�v_� Hl�i���fwI�d6u컼��c�u��F�a&/. ��v9�ǉ�;]�=G�����̑�������[.]��JI���ƘA���z�.9m}�&� ���<k����l���Nzx������O�(�Ä��j@�DiJ�a���1���	Z�2�&�Yn�֮��'�ߚ��N1�L6w�v-�$G���_�_�A��������[�a�����L�}:��H/���X�N�����/+������ � �gg1�6xl��n����L���d�ú�����k;2��a�WZ��d�3v͡�I��`��˱	�OJ�9�,�H/�M��f�-��㧪!��I<��"A'��YںX̵�$]�Mv&���B�C�߷�8�B�{�C��u�Ag�����v�e�Ԛ2�-�9<�rxSW{�ш�ү����"�B�k�}F�tN�� ���w�cw�oљ��qр�3}������z0Kh�cL���3�gi����Of�F�GMd����f��"w�$Hm�@��X-}1Ǉ�1{
Y�pz��ٴ���e�[���i�fZ]�G���>r��H'p_�f�| �n��$�w>�����VB�<�d���邊��ɐ[:Yk��ü/Dy��g�S��$���2�[�}���$�^�QYU1ꍨ��6Y���0rSE��5���� AfF�^�z�'Ċ��$�^]�� ���d���;)�u�j��o:�&�f�@�WLI$��w�H&c��^�����,May�ڡ*,RZ�r���L�ͨ�H� &{ء�s�(�E�?�_C��3�`�V�uȌᤉ��wőw��91j�!&�YM��:�Z��sc�Vu!g�*dzn�pA{6Xl�t��cL���Չi���J�g��x�Ġ��p�5�b�mn�؊Zg��3\��#vs���TM����1NRXm��y�,{H3c%�јT*9�R��*�QՎ&5���t�V��I��GB�!�f��L+��V�4e,]��*�Gmz5r0�#@�[)� xle�lŘ�2r̆�.���-�a �n�%�i�;.�f��lݭ]�m�V�(kI�Iu�GYj�V�.cl��1t��t)+�GZ��e��f\� �GF�����Y3;�vt��7��_L��|w6�$�n7�
�U�k��w�{'�.�_ځ={ ���˗wb�A;��>3|�Bl�ԣr{b�y"M���� �1���|ӽ�C��2k���-{,��r�
�@�l��<�Qm�́ ���z.�H$���&5�ǉ�4�V�&̋����-�X5�4����C��d�@�I�\���윁n���X	-�p�M�Y��,���TS�t A��Ș�ƪ�[�[�0��'`7�"-��� ��쑻�������@����bS;��+��5��@b.�1v��GL��Y[�Vաb����?m�y+��'�w�o\Gx�N�� �ّ>.�����ր/� 1̈́@~�H�g`��3�竔^��F���̾�.]'��_� zP����y��<�<�~��?vC�w8{N÷�՞o����\������.N�[�{�I�X��/!�o����I�`�C��fI7ki�l�n�0M�wv(��/2޴���� ���)�x��i��Y(� �����ײ�]/1��$��-+�y����1T�`�n�2'đ��-X�m������m0��Kf	�tE�I
޸��{�����{�w�Ϧ	'/7&A>#��!V֎���~� �F��1oȬ'V�ZR%nD)k�	,tc�
�� ���K�n�x�\z��|�s,.�7��l<IܼȐI$����x�V��[��q�-��$]e�x�I&�������v"�]�DgK�4�׭<�����'�$�e8�z�d+v1u�-���$��fgL�2w^̂I���x�
�C���c]�0 -{��d�P]�։�R6�ۀ۲�9�1X��64U�#9��^]Do,��~fS���mX�*_bR��2��������cA�ʙ$O_SǴMd�wp�#����?�g?3�g��m�;@��}�Q!���O �k��ݱ�ۯ:�e3��c��$�]��D<C���Ey1��4�0�M¹�}�*�a�A_\z��~1�S���41���7X���v&�;C65y�cuX��4f��$���Bh6/ T�klsn���*�@d���ق~�h��� n��	&z_�	ʨ����H�� �}�N�������ʆ�D�DH\�ˈ�Y*�bI �o2�	^HOK�f���\��������2�8r��&i�c��A� �Kd ���Q�,��)���:�g�'�t��>����d�33�va,:w\D@ׇʺ���M-/ ���~0I=��8.��ۣ��5�����e28"2-S6!J����Y9�m�P��x��),��J"���"%� ���U�u�:���X?����?�1� A���t�+����ƒ �̀�U�]�&s�KE-" w���0�ol̂�W;�go��K$���dY���١w��jݲ�K�45�2�Y[v��i�����}��1	ל<q�{�$�v�<����&|r"�D_Su�y����	ʗ�ت��2��`�=�2Igi��9Z#�k�Cv���$EԾ��^Av�dψ������܎�m������N�������)�aMWnG��t��ŌlZ��뾢A3R�`���̙y�)[����2gQێfx�J*�F���GĂ|/{2d��^+:sZ������pE�>��i�A"�C&r��-��2H$�l�����P���#I�;&AΘ���!{�e��}U!C�g�ꨒ9�D׆3�ۧ;�7����2���\�=���v���*��T.�u:|���7��>��-=�>�]���kg�:�v[}b��	V0ã�<��+�[�X��Z�s��,v�o*�{�p<_>����o�#���ҵxֳ�[.����g�n�>��ᚨwn "l���ѣ�r��:]���S�HX5��3�������u{�ڴ��Q���}��/��x*�x�7^�Y���.;���l����ٻ�{u��r�u�)��W{	-��?
�y�X�ao6���zy��'}�<�*ГF3�����8`{�R:3���8��ʭ�Wϒ�o|<�ZD^5��3�}���샷��c�<I��������UO��GE^�/0}�B�<�_z4��r���^�{[T�Z��n돁�4���F��=|�T�;���ԋٲ)j{g��l�|n��ɋ��ɂvVsj�J��$���zL��	vq��:'�h{Bl�`\��/�#@�G��~�uj��{5ޔg�P`hkP��N��S�bn�
����^j�����}��.!C�lu9X7T�t�t���^�;Y~��/i��r����`��"�[�ؖ>ka^<u{�Q���4��8]�H�G�[�����M�"�w��2��Ѡ}i~��{t~�8�<����I���!�7Ѭ��8i�f�a�,��]�xxo��n	�4��]�Т�ڀ��HƂ��;7�=勶	v��^IT������V�$�H Y@�mؖ��N?��w��X�i�ۆֲ�Í�7���P,֝��}}z{q���������^>IY�IE�bBX��ݳ�q��N�{6��rI�R��HE��;(XB�@��N�_q�Ƿ���Ǉ���~��ߞ��Y���R"�blr6�D�E3"	4[u���;,mE��;[I%gb�/;�fq�XK�:NR=����jf�J[~��;緒+[|�製�٭�_*�\w�!-l�,,��VY%�lp���V%�Im��m�mm6e�EM�m�k�����!�l�,ͷ��֓�[����_=b{X�%&v��h�[VW�{ň�m��⃧[l�Ȥ�p)3p���s�Ҁ�H��a+l��R����/�v���$v֥"��d�ziJ�M�fhqIRγ�Sy�m�Y���2�9l����6�rN��w���h-�N6�:�V��>4�ݗ"p��G˝��6��ݬN9|��u�/�������{����<|�W���]�YY���
�W-�	�=�VҚ�C�����Km���̥��qkՐ+%��к4����6�W�๹��D�ܓ	�:�iH��������efJbX�+�s�#u5%\���+.0��̄��.��-֌��dC:T�]�Y�9�+[j�!�����1ZB�Kv��veu#�L��+΍n�n��L�Zk*����6\.�]Ku"�M1-5��c�F�-��Fܹ�X�X��YM4W,�m���)��GmM�����#��%�]H�]0f2�E��,��Q&����J[�M�ƚ.e���r�	�8�&h,M�#�ʐ��mq��X :�^�W��l��\�sV��88��Dfʵ�в�a#�j\b\BBjP�j��.&�������,&�IX�\ԅ[� Dغ��l���P�
8�&j̋{K-#�0��f�<�J��i[[5\�.nL����t���[d-�k�('U3���T-2
�x4e�F���1��GgQ�]�fx9�m���Xu-��̭���&Pc@�QK�cS)s��Mob�W	X�����4e������F�*`LlW`�0��rj�M�ԳP�Z�i�CU4UR����4,k�X���,�r�@4�itͨ�oh���,�j$��sfJ�n4Gk��Z˫S[L�,��CL�(��a��X޷"<Ř�m	6�IXD��,�vAnm	�.)3��a�R��m�԰[�y!��6\)�	X�&�ZU�4���&)p�X �Z,weɝF��%F�,f�����4�IA-�ĻV��:���%̮�6���;*X��$)5�Uå�,5�1�F��e0iV%F6T�/-��4u�Śm�[�KX�K.%恑��W6j�ɓ\�M��j�l(4]� ʘ�%�Ȱ�����sV��]Ss�RjKU�XCK�ՙ�i�U��Ba�ڦn!n���aQ��F�+�Q� �jx��Pj�\�鋀�T���Ǚ�x���x5�ߜq�g���֎lv�	h933�v�<G�G�3��H�{Q��	m�V�%`4��
�Ts)���2���c2�4Zl�f%�b֣)���v�ƣ��t)c�z�V�nm1���6��6�\^�ö�f	٭�a�nE�r:[@KU�Vd�s�,n�:��ك�F]�dEִ�E/2�dR�SY�C����>b�(̎��[��xL[��K� �r�Q05�K�3	��vi�Ć�*��h�ATF�l-�>>�����YR}�P�kb�Ngf@�H�$=��⢢����
����(@7���1�m��P�xN���OC�A6�&R7ά�%3�>1��ǉ۝0 V�-܉�l�ZH�u�,\3b��y�&d����/Z"	3�� Z;+º���ٙ��>$����q:fr�fp]��S�|n���/�S�D��-��$A���$�+��xMn.cv���\�$3X�V�B$;8L�&3�� l��yۋ�}��c  ���Ǣ�W�����F��w�=�g��g�Ŏ�-�.��b�#02��ؽ���6������~�����������츀	�-��"�tv�ʥ&�/�fI��9�=�Tnuݙ�y���FMd�r_�M�w=t�LeJ���9M��)ř�UܼU�uj�8��21�I��KW�6V��`�#�^�*}�{�z�� �jl���\��+�W�'*Z��8,Gޟ��� ����x�H����	�]*8�a�r*w7Iy������ p�@�>D/$0��A |뫎Uï��x����q �K��< ������_��-DΡ�?�MoL
�H$d>�3��$ugL�m�t�9�[l�||���:�&t�fp]�g�j��>'ƻc!3W���Õ��r�^<I"UδI���L��E�����_[�aͶ"g�Q�˛�$[t3-�S�Xaٖl��8!�����كYs����3G�H�Jq(���2�}��'�|��" ed�A#��7Z�E��L읠U��$Q�uw2�2gcw)ރz���6ƴ�Ou�@������K�`���k�3�
�'�&N�@r��ǳ� Q&���6�'�W3]��Aʨ3*���E[|p�����n���wmL�m���Ǹw��\I��N��&[�����D���H��x����I4���A wvd�!�w���� p� �>t�v��MF��T�2\�MVnL��ۜ�R������e���߇P ���8�_/褂I5��U�m~�$R�怒'���ɒA ����F)��+j�8h�25����a�bv��U��lW\���2��	�O$0�&ιT���A�;��ܗf��f�c�H��ȒI'�: m̤�u�9�H9���I�&|Ks�kgr���O2����j�Nqw�!z^^��I�v�ɒ1��qB����`F85ƭ$S��k	Y3�v�4C����	=�����l3�3]y�U�@���"A'�:>ɪ�vg(��$O&vX�dV���ZMQ51�> ��r k�y%��p͍(���ي�o�v��PA��Q�����������f��5��F�q+#�W ,�%�(�f郖��ý�>><i�6$���[Ǚݔ ��OFDzf)��b���O2�z���HH��"=Jy@�(t���o�=���.��5�9�!.kc.j�؜�^ܓb�G�+M;3i�г��������g��j�Ƨ�y��	��.ƮP��-���Dot�����=����8��w;�.�2⎀Ğ�4��ϳ�=YO��$�Etl@o$	��O($��J�^w������2���7�;�O2t�L��ت#�|H7sL{0b�}��I'm� gT�C`�j&Rgd�CunɁ4�7s�|{��$�H�i�$�ے�b2��A殈>�98������d�,�i�D�tdI"&f��aJ�0���SQ $#�:���#[�&A���,_m˵Q�Og8�O �(�*wT%����#�X�#Yp��x2h��v�h\[,y�.06D��:�w�McN����>>>֬D��c�75��]5sm�f��&��jP� k���X�vWK��k����[�<*桢�P���0�cH�f�QXi��f�]3��ͅ/AƍS4,�uàlh��Ł�3m�JB;MI�&�P
Vj�n 40f��!sn.F9k+�.C:�\3[H����-��6����\V �иe�6jjM�h��L'�c7�4�VɋG9��5�#x
9�����n�]j��P�c �]�#S�3r,̼�ӻ���7���� ;���l��w�1$�3�rd�R���O�<
����B+��[�e\3b��y�'=TOyEb�s=��z��b/ҁ�j��z�2g��>@#��G��'[Z�����g�fgw]ػ4�=J9@'ƺ�"A �܅ ��4/Ċ��Q>H;z2d���Z�܇;:t�&3�n��8����N� 1$���nТ|{rf�1��`�_�9_���t�`�&vN� c��$��ϤN��[�
|�	�j��|2�2dI�:=1���2�z��bb�;�A5e�e)���%Ѫ�kA�V\�����b%����q�ݙ�))ÿ����'��"H"|�����hU�S"����_vL�_8-��X���H=1ǘ��B����X���g���R/t�z�x�=�7�E��l�;�����{����YQ�]��E����Te,�!�_�Ȃ���w����-]�om�dω�� C��S=%3]�O��5���7d�m-o��&\3b��D�ٳS$��t@ �#3u��Ȟ�ń���ܙ�'rz ��3�fwf!����Ux�Q�9_X&�ӻ�@%���^1 O�Z�[��6���X!���I��d�mvt���ӧ����Ds˒�J2ܴ��$L7� H���A7q� �<᠛��1J6�G06d���fgu5 �i���]���WS5�э�f豳2��!��7��QL�Γ�w��} ���A��\�Ԫt���>�������
�Aѱ�;&�];;"�b�;̞5��]�^u%[q��A>q� �ʧ�	1��vG&Ɉ�_t-�y,X���H;/�g'��A ����`�i���n��4<TE�H������h~�ׁ�zvS3���7�{������w}��=�{�SsgUp�,��u
����-��<������x|� ����D���t䔛��v,$�wD��G�������|H�q�ęYݹT/4۬����hgm�;��$��A�;����� ɨ�r	=ۍq>8�ܿv�{�K�ۑ�E+�h"3�r��u�5��0��$��: ���%v�51
5��x�������X���VYb�'�>��[��'N��x��D���>$���s&!���;"nSC�h��� �9t�C�'��nBL���ɐH36gMk�^599��N/�I �>���s�K�w<	�k���0]ߍ����;��:E)ü3n�	7��I �٬q��Y6� ���&	��2慶�	���=<���aZ3|IG�X@/��ؑ~���֎�=�w�4��9nSeM��N)QQMta������W:����{����~�Vwd�Z� 0���S�Q8�'[f/@�׸r�$�Pe�y�||G�B�ƀO���$�v��`�!n����e�j�u�ű��)�=ys>��=��S�{6�����ZZ���%:@��pG9n5R�[j�)�%�(�3����4ҧ秤���\�d������8IO��8';s��'����^M�X��6��i�=M�n�ndnA�wwL���ӧ�*z �x)--��.Ș;%V������]}�BI=q� Q�e�9�8�&�9�z��2o8L�!2+vD�{rb����7&I��n9��yl�$��ˑ$ntǧҶ�ƺN��A�p�2x�Geja�����z��O�N��LA S7�]s6��E��Q.�r	U��%�B�w�`� �`s�\I�Jyo?>{�������TU�� oLʧ�<oޙ{���ʔ��cpd��G2�[�M&��s�Eg��������w���=Wz�=��l�����̉!������?��Ύ�)�'5N��0��������x�j����#ٸ0�gRj�f��Z�YB�n��0-�⋭�p�� %��f� �w�ym�e�:���2�X�,i��[���sfF�Y��:�D����afs�C un�ș2B4�G�2͢eKI\�#�����U����ۮ��D4�+WD��m�R�6ї3vF��v+m۶�5c��a���XO'��x�����B�gW5�6�ZE;HH:К��M�،c�#5)�kw�A���Ҽ�h����{2	o![�'�O3zy��2�t�k�65���d�^]�/���d��靚z������OJ���Dzu!{��|H�S� �N�t�8W�c�����;>۳�f�N�<όf�zy x�c-e�:�[�2��G��dǠ?�nh��N�Y����v���;oI���
Z0�����|�h ��\�1r�;�G�oDA�I��)Ӳ(2N�A�9�>$�v\��{l���K��$uEDf5d�H����N����dA����3kU���ˍ��.���t�e�],���ma��T�<_���}���O�n���`B�F� ��˙=��jZ��_$M�M��9(����us�Y%��i�0�gc����́&�<�H`�Y9n�>��m��p5��{ӡǨK��[���L�{s�ܥܥN��~��<|u��	 ����I �Ov\ω-���L�ɣs�29���d������&����- Ȃ<g�_f�I$�r(�vl�1�]{D֞P ��̙3��.�S�'N�hΫ��&�ңn	 �)���'7�$I'����؊�B:c��f�P>̂������b&VV�ω�ݘ����́=7E>��=�$���گI�&".����C���M��^r�Çxܵ#MZG1ٙ����Ba�����jѻh��U��~���:vEIÿp1��<�w;2'Ē	����gy�++��;N('ĉ�ܙ //?i[��
e�$�F<x�N=�F�uo�q4@bH$�̑>$���1e�n��_��ly!{�8��.�`�<
�g��I�����j���dQ<㿑}����M��u��}����W��4���lw:dK飱�5�?v�@`��I61İ���U�����{�q�7w���9ZX�W���<�QLY�1�E�Y�C2ȹ���C0��Rp�<���Z����{���a�S�ݻ���\=$?yzs�}�d˰y���2;���ǫ�nh�[��-ޏ9�/9�f=�{	��ik�'�z���]*�|�z:�_�5�����X ��w}�{�OO_/i���*y�wx�x�޳2��%�"3���6Eƣ�sO����Zg���rS�~�VF��.�b2*��w��,&L��MέQ�{$�Ӳ�"j�ͮ��$򵸏�9�}���}
�R�ޙqz�^}��h�Ƿ�8��b�j~��D���/@�vyy"�G�A����6h���2��.�cҰ͏��OLg_y�ˏ�b�<h�N�?{��b޽�nh^��^�{(����P��✘��ra�Af�x��E���{B���5awY��o{�U���Y0/��7Ӝ�<���+jĞ��U���e�$�`Ě�\R̚7"�z��7=�M^���G>2A�������a�֩n��B��x}嬏M�{n��gnpp����%K&��׎vv_�tw%�ۻݮ���ѱ�p�.adMٕ�r�D�ʰ��i�h�r.�E��a�Қ�!Fj�O�*�х�"TC�t��u[�R�,!A �I)aKm�d���8�çB�9�k9�$(�J�$�!-�R� c㷷�^��|||y|q��闙K)d��JH�t��̹:"����s��8H(E�m��Z@���!e�xzz|{||{{q�������w�]��;Ͼ�pc�Y9%�9���߫ב��Ӝ�:S�:��m��^yÕ�bR3p��p�(\�Z' �Ə����`vڛbr�D�؄s�Ns��DpJAH:D㐜�q٩^vط	!���v��5U�|nmY��@%�u�k����yd��$��;�BJRT[Y�ZpRs��$���I}�}��G7v��Y�
�Ŷ����V��|՜N�/���8(��{]�Ey�n�����:�=�;���r^j��Lk[e#��H��e�$ ��p'f%-��8��ؔ�)�Z�3v�uf���n&k���$�
'#�v�;ߞ������#=^Cw� ���N�X1vwf�������6t�&��$n��$�6�c�'Zy(1���G�h���H׼�.�&�N�Q�ځ�_+�lz�i��	�.�M}2I>9�1��֠�
��w����(y�z靄��6��)\�hB+�. 6h̗��C��Йo��g�=��-�����}���Ι� �����'����`�o�^�ST7��}���>����QѤhX��9>(4�k4�m>���˓�BO�8onkD|I�n���"��[��|�Hk��n�	d��'�b2 �O�b�į%��Y�ך3�0�H=�� ��'ZyG��]F$ዠX8f2�����f���A���$���P	��d�'�Br_�s?�f����N7��l�zj�}�/=-�4oT[�ѷFI|��,�)�l۝g�#v�^)��t���!�/f���|||x�k^�������.���g�t�{72$�v�ȇ��\�Č��LO��n����nvD����Fg��}��?Yj�����Ԏڣ#h-͚��3�e�Y�;�V:5�||�.�����k.Bj��g���YP�|����2�t�u+kM�SA`啠@')e!h�r���ˇe][Ev]��3�9YN5��� ���Q!
���2Cy��V�.69����� �"j�t�b��x�PS�27�9���H�zK_b}3���I�WJ	$f�dȯ$t�[�BY8�:�ϐeN�CXo���$�^dH�� νT,�
���#O�95L��m֤ዄ�LL��X ���1NiN$կ�J�f���oWnd�>��
�ZT�t�nQ*B��r�6(��ݯ��΋�{���s� �V�=�V��>eg^:�pĄf�k����Od�4p��sO���� {�E"�%-R؆�f��1����0bYZQ�q�i��+�CS
@���&����:к�6׎��h�t��x�,%T5ԆV��!P�8m��X��v ,(�S
�������Yf)���F�tb�Y.��e����Q�q3q�Ϟ[�I`�f����s�����bX�]��+6�U�rmd��Ύ+���G#m��j�j���+�~}��E���&�X(X��\����fvf.t�)/��|���%Ϊ�����Ϻg)fnW}���w��DgfD�A4;� �r�u�7��|F��|� �}U��$�?dYt�3�3�y��� @XI����w$�3W�2 �]��8��fV�6��"��b�$]�p�\;U~�� �I�ڿD�zA8Z����3��I�nd� �MoT���;�`����$���&�E���1�GP���ɉ� �
��?��γ�̩鵉B�����lH�q�t��qu�� A#1W(�(ƥ5��zv�H'��k���d��{�%-��2���>���Y=ϺPf,A�.�3�H�*���9�1dM�tH-���LVm0�O����7B:ћ�ة��_SǉŒt7)5U�.�w'n�*1�@$s������;;��;;L�����~R�_�j�D�6&i�݅`ߧ���Te0U��]W풶��s,'ݢ�[��9ȋ��f1�I�0��pE
:� v�Y�b��~/G�g�����m�"�H$�*��@�u�� I��μKZ��7Ć|��,��,��<
X �A�U�G�<𤟎��<��I ��D�D�W( 未Eb0w�v��֛�|�g�	��4H^&��TH���n/������+@�: ���a���2Aü�n����ɠoo+3F�m�c�<O�^" �v�� ���^=-�*u���zkEj�(�`Pr[���[Xm�[�4��2�YU����¥�;o:z�}�t9' �P_;�3���%�>$.�ɟ���-��y�w�8��5t���Q�?�����,'�F��o]5�$g*��;��g�<����m��^�c�[�ggr��gN�"O2�P	7ۙ�9��p��k+|��`� (��pe�v��l�2*�{�eQfcP4���9�W�u��{~��>��q����V�p��DЩE�d��������3�=���ށ9��	�|�n\��w%�wt�'#�5;�oA�<V�>/J��;{� �|o���Ď�HR�
	��QH:!�p�e��dH$�U[֤*���)t�@�n��Ef�L���>+��!8�|�R��΃E�LA� �N�]k��0W�Xj�[H
d�u��R�/���}��-�82H8w��]��}�I&�� �;�9NL�9Đw1u)�$���9�>�s�I�!�I�6 ��cTR�����S���+[2$�M�Tz<�10��9a>������J`�&F<t̃쾨I��S���x���mr�O�@�k�}������;;�K�:g�CiC��ȡ��ߋ���f�	"/��D�	�k_+f]~n%�:_ur�#��œ�ؼVדb.6�T�1m8�e�5M�P�r���!����Z��:ُZ`���L�Tſ�"�w���x�iy��C�\�g,��$��Ϥk�؀M�V�s.l��.�;	�Χ	�\�w7��}?=~~y/����b�$(�jes6�SҤK�!hV�c��2̱��g߯����#4X�}�띓2O��ڏ	7�׾RtdhɆ�lq��/U2�v�y���)�:L�2�P	v���\�7P����y��|�H����L�G���?w��O\!ݮ�:�G������Aa���3*��#q�:��y���w���'��<H}��I��g%3���Qx`�.��_� HV4�{��U�B���r��H)�t�3.���Ι�U��a� �^d���3�c咽ۓ2A��'��	͎ɐi�%k�ۥqpJ�T��ڪ��^1�Y����`����G4�{�%�qD�J%�Qʗ	K��]��N��I�rTĶ�{�j�nճ��mi�8�������儏�U��m>���{���~�:Ԍ�h�"�t^&�a.3f���	U��6;ζL%�sq.2C9c\&�cÝ�k6	�"��\ZY[�\��:.�,�&�X�!6SF���:ͭ!qQ��km�QAYKt���s�9�]��&�v� �[)���q�j�R.�i���,�JCGU����8��6�k�˕�[Zc"�.�i�Bb05f�	����E������̳�� �k������m�cX�Ku!M�fYfT����M�9@`��K����G[]� אH�d$��}�&��2
)��-�3� �oZ	�"��D;�L�m�ψ/ՃC#��Ƞ&^c�	7-��wo�D�5Y���ҭ�A��ڐS�t��.CZ�o_��e�D�	�bS�:V{�}>HU7r�Iٙ!�FV�.L��Au"0�Lbֶ��w����>5��D� v�2$H9�S�_wz�h�ُ&���_���rS9����L�I�����֫alN�>� �wfd�$ǟ�;��e�Mnj�G�����c�\Ku�$]c�2�7Lfm��2�9�K+�vڱ�=z��.͋ \���=6G�&�s"I${;�$�A�J��`I���GZ���ܗI��ȝ���{۱c�}�p"(�)j���l4T2|���z��.]�#�+).N^��4�2~�{턿@n�ǫT���ߧhO��*��Hw���ƪ�x"<D�^�d�=!��H;��2���h�v���F`��!غp�2�׳ I��$�G/C�=����Z���3&I$��<{kUHd���"��̂��l���-��~Zu�ĂI�ͦ�'������iHU ���-�k]�&\G��y�2F��3p�v����Ȱ'�Dg L��L�	����<L��a1�6ug����pc	6�jd�×d�.��&�ca�h�̤��m�G��W+!��Pa�)S�1�9%���w��j@���ĂD��h*"��UЬ~�#M��L��M�TA�X�΃�$��vw0���㩪qA)z�f\W�'��uG�J��I1���n���.����'*U���t��:><�P"<���q�$הV�b�=8Dh�|u�$�ت��+%ĸ����#�C�y�����LS��5xEFs�2�ٹP}66�MaA�q�g��c����$���&T�4X6Ed�v.�;D��og�kZ���6Z���&|���3|� ;���͂7y��� �����5!��L�3�\�\ ]�X��dI������ߋDKǹ��S�';;fNX�h�=����5���%�ŋ!�چ�3]Յ�V����\�&�\�..��P?'��ݚ}dz�O}�3��}�}� ��Fq�!�4w��A$�kZ	�˒�tK9)������I-B�s��i���R�pI�֏�Fm�L���&UR�.'9�r���gA�]اy�rty�={�|I�����j�=I�k��	-x�w��g��c�H`��K����A���D���x�F�#����}� �|s���#y�M�$݊�-5�x,��U��Z�c4�*^�|C~�O;�<{7��Ҋ�2�L�W�Ai,Y�3TC�bZ��^� `	��� ���8vI'E�ó�z�u�"�i�tt[(w:d��ǎy=�Y�I#��'�C��y��04����~{����l?=�sV%ib��L���H!^5���(�Zkv�&��z��ľ��+1����x�k0	7��A9伷� �P�\6u��r0�y�$�s9��gF\G��y�2�L�7����� ��5$��A��ʯV�;x�m<Zjs��y��7�r].�g%�̬m{� �� A'ŧ�S�wu��Wq�`�'� A&�� ��k]�pIwb��IE7%mS&}�$��< H$}5��|H����<�.y�����LLa���ܗI����ف ���a2!������Ho4�L�a=�7��$�������>���~�DV�P�?����H�������E��@�<��*`�VX1Q`�E�TX1Q`�E�TXTX0`�E�X0Q`�E�X0Q`1Q`�E�X0Q`�E�PX0E`���E�X1Q`�E� VPX0Q`��F������� �`�`00X1X0X1X0X1X1X1X0@����� �`�`�`0X1X1@�� �1X1X0XV���� �`�`�0XVV@����E��<�
`�`�`"b"`�bb�b�`"��D �D �D �D �D � �T �T �T �E�P8�CQ�+d�#F� db�����
�c���b��`�� �V 0# � @�� �P##@ִ:��#�@ �P �## ��X�� QX��  �U�la���� A�+
�(ъ�(�d`*�F ��b��husV�X1Q`�E�TX0Q`��]Ph����*,��b����(���`���+�Sp�09�
n}�ܪ��H�*�`( 1�������������w�?��?�����!ꇐ�_��?�����	k����q���>O����g�����?� 紊((��?p�����A�?j~���?�}_�ࠂ��?/�~0��ۦB%�7���/���� _���d��kUX"�+"" ! ��(H��H��`�ł�*,"�"����*,X(����� ���+*,B �*, ��"��H��*,��"��H���V �F
,R
,V*,H(���b��"��"
� +(��+
,`�Ȩ�
, ���)Qx�����t}���
�,����H����}G�5��W��}B@�����8�u��qQ]��~{8�����v'��r������0��'����PAE}�֟���q�&EDW�AE~�����|?�o������������
�?�(��&ǀ�%�2����p}tD��~=�p iA�����S�������PAE@z��hw�'�}h~���C��>�� |���A�����(���̄?���ܠ���@�a���9	�_4��(v�Ƈ�?��;�ﰉN��TQ]&�$`t�~)P?`p��'�t�>�8�~�  ��<�(|� V��^|�����?�b��L��d�Y(��� � ���fO� �?7�   �     P�  �
     :   �          t� ���]7�T�%N�*��D%U*]kl�Z�[*��"�J�T�JJP�(
�QU�E�eJ��*��J��                                               �| d��
���s4���F �FC�ǩ<��JZ��y tu� ���+���**��R)>   '�y�  �&Z��@r�H�jT�\��aT)*�� 5R:2q�ܥP��Nm \�E
�`��%��}i
�U�  �         ���B��=�t)J��)"VX��NƮ3��/N ��P`ޚ�El
BR�,R�_}�/3"�(C �JE����f�1Vǧ(���  �>OA{/��� tC*-
=����u� TOs s`�1hlq =ޕQ�Q֑$|  �        }�iK���4x�u�f�a��L�P��x =WA����y����ŻD\�jcjp 릴��ov�/,��8�B�N���  �O�|��j�ur�mp 3�fkr��Z��;�>�t��p�"�3�]/g��sQ�s7��E���W���c��n�F�l[ʒٕUJN��  >         |y�j�g4sd_yζy̐���;r���� n:^�^mr�ճ�v��ncB�j��q� 掵N.����ε��mJ���  d|ZVj��sfp 3��9����vll���Gd�0ґ�^ ��]�,v�4.a�l�ۋ�Ya���iz��%4�B|  �        �}m;�SZ��u�m)�z�\�Ҕ�� gu�N#$�Y0�=�o9;,�ԥt�� <O`�b�Zis4��(�@��  ��z%fʪ�n ����ˣ��6���� &�c݀9rhrh d4��MIR�	� "��M5%J�  ��zj�I�0�B'�U(�JR   j��&U*   iS�R�z�A����~���5~���}�f}3�3��h�<8L���?�IN@����	!I�! ����IO�H@�`$�	#		����q����c>��֝gtˇ���n.A�A=��r���wk��v����n+�q�/ǝ
��'`�� 9����ᇛB�Ln��@k`j�%v�
�����]K�7v+Ӫ���b��[��|���N0^��}��aOX�-��x7�]�;��^�V�7{��K��y` ,�C�Ll:�iGz�ݓ��S�7*��{u�i�n�hz��S."��_E����&Lc��QM�}��;D�"Xp�5[3�G�0H*%I�h緦B�T�5�㺵k�y��v���X��d�d�7�iد�h���Pn�.���TP��\j^�j4hy8��U�g3,ū(�=�eͫ��@.q�j�ۈ�Bñ��f����E��90�[��<�Eٻh&���� �����Y���Q=cXY6:��X4k8:��F̉^�����iы��5׫��ӌ�h��SҠxz]�B��=7%l�xE{v���ݥ�Z���9o�ǂ�'gu]�]3;E �{�R����ǫ� �ζ;�e�S�(�D �%�$h�i8e�iJ��r�DWu7\���o��X���%�I���w���-�+ڐ�oi��<'N�7p���[����*���_��W����dۓ���D�dqs��'UX5+Ҿ�H�;���m��{ߡ���{�K0�Qmv2GYwSgk�H��}���.�}3qO4����lUc��W�I��p�X�i-�ΔѸ@��r�7|c�22.����;Oh�>x��h��M��=ۀs{	%rƘ	�7;�}2�\ڒ�N{��A(�{-۽��1�r��..ɗW��'q\���96�w7n*��C/!��O�Z�wI�p��b�y�c�5�!��saVLX��N�ܓ�^7�s��T�c��V��;�3�@�]���Ɉlnrܛ���-�$Ƶ���S5J�d}�u�ç�ͅv!��ŧ0wM�YJ���tS�[6>\�]�<����^���BF�8�� ݖ��tʅber����c`�'h5ݕ�@��иw�����-����Qi��k;V��j&u��rx��a�'�j�1�8��o�갇�y�og	��3�,(��0��
"�ˁ���s%<�o���N�]Kx��ҫ��[�ₐo"�2wFn��x.�{SB)��.� �4س 2�T^�ƔC�9E��y��a�vCwq�x��6�w#�hNm��jlo��f݃t�[.,@���%C���ޓf�;�v�Hb��٦��w:޳3���<dZZ͓HO�V��8�[�r�s�����q�2aRƪX�^���L���e6�Bo[L�e��ҰP���Háޤ`�u*��1��Ųt�dK#6sכx��ߓ!nA�	^b]�e�(�o��B`�7�wF#��nG��)��G9tRAo,S����R*ݬ,+�"����f&�W��$n��2������N�I�c��{Z����=I��ُN��sw�H˅�.�����ҭId�*�8����t�n��;���`@uo	�"����8y��r���^<Ưz�Oo^����;ݱ�R���q�0�(VÐw��=��
������n��V�����Z!������gHp���ŉ�N�F3w_P�v+41�&��&��R1*�1���M�(h
a����l�g`�w��l㠝*ΰ�X��pY|�C��6q�i8�k�w�i�3��!Z�ǥ�iŮƪˮ�z�ó���f{)��-�����%��CnJ�:l6,*d��B$�Fы��ƿkf\Gv�ҭ�7k���d��XA�Q_.q`z��3^�jX�oM(��E+U���n���KՆ���$t���ICG❎�z�rFMzl6BtcY�^��V���N0;v"qi\��pg:���Q��xSXrlo�x�p�f��}�恋=��sb�L����ԓ�suwof��q�,����+@���w;w���8��q�j�F�y<��P�;������ᗳ��ۮ�78�ie.H������f��/Bz-�NM��GG��x
BQg1���Q˖s ֏;{H�c�N�v.n�2��$�p�7G�'y~�����9y{ިh����g
�.i�7mœ{Yĭ��adB:8R5�	���k���#=0�/�v ��  ub��L!:�rȦZ��n��q��N��k�v�+����U g!�Ā���ש0HfS�4d�²�j뤤��Dڙ���;��)8:�:�zF��=�e�j�2���S�����
��X���Y�D���ba��;#6d�wf�LAV�Og#��D�:;��Z!�u`ƅ�s���CU�^��i�e7.��wA0�{����Bوh��W�J����j[�v�<��~�̯!�I�yC�N���p,++([9����ֺom��Ò��38��N�;�X��D`s�tH�=�	�_���T�w_f�ɦ��r���$�h����vĄ��N�5��p�oq��F�g,��MXK�����?^5HF[�����j�ĺ>3w+�حx�<��֟�:��1HZI�c�m�i�m<i�wqb}�7vog({��g������`c�NVx�)�����K�Zܯ@"O!\��)�):սۖͺ�5������o^����/s��5���=�#��W )�
整gj�a8}��Є�p0`&�J��д!�n撶�y{8�؃��w�ᙺ�;�L��N��5d�̞�՚^�q'B�ƌ:t�J����3�wt;�KO��{o09>�˝:���m�ȇQyt�]L����rgb��C�m�� �d�}�FY��Ԙ<X6�v�y���q2.ݳ40*ΏC������Q1˶v<���љ�(��懡o�<M�C��ɐ)�Tp��,<&���)�N\�6ӂ`� Z[;Q�Bɸ��uN�ɜ۴fw���95�,�v��ҞIV��p���j�ᓈ�8)'V��v��-�g`(7"���=���z{5-��󆫺�X@��^Mdr&��u�+w-��E���/tm�teD�Ǉ��wUg;7�q�ē������Ƹ]x�S��MC�6�)��q�J<�8W<)��ÏX B�-�	wN��Rj�8�C�����.�|t�S�����L��� ����77�o\"s�Yϯ*��wReI�ln�[.8���&�+�i�;R��Sd�)F�$��-7�ĸ)���;@�zg>��	�mCq�x�i��70a�Vn��!�uR�Nv�პ�v�vF�w��Y����u)���Nv[L(ni����bw��r'@dj�2d;{,��l��)�r�o��Y�*�1s�!Q����2]�ev�yn�H}����V����'v�2vm;��~3�v��?ɩh\C(�/���$w�*��7��u-�6=����N��6+�P��xr0[$a�Ff�k�ަs�d�mcq���q�f���P&k�X%�k�BHN*�e�H�˔��&����r��J�̹լ�ȇö(�+��3�.���+IǦ��r6�Z�Ť��߳_C0���Bل%����ۺ�M���Kޝ�DX�,u�X�9�иuKur���'z���(�H�qb��X�r)�ms�*z(���Wb��Gy/.VgaS0��]�79v�/+&귓1�;qԳ{T*�tLe�r�tSҕ �\�S��jw-�f��Z�XYBm�Д��.L�F��1wpޙ����8�b���z�'��x��iY���ȓ�{;J�[��̬���3�;۲3�s����0Qe���ܯ.�M�<��;#�Ȼ�[�4�j���KE�m%U�s��{��w�^�8�`:&�R$o[�cM�����ţv�IU�	�'	�nl�qu��vL��.�)5�[S��E��b��i���$�D�5�Ö7;{�c�7Vr�
�p� �X��Ur��u��#��cZ�REXw/rU�޳3�_r�2%]�j��ҁS90#��nSE��f�T�#���ѓj몳 ƻ[��a��H�y��C޵��3�-Yv, 3��yv�<gQ��p튇�bQ
3d� �7�B�s��TO�������_U�=L�1d�g����K}t�ѓM\��Q��2jd9�y]�xw�j�:ۼz�����8�]#PC��w4���8R�ӓ١�Ĕ�ETǻ;��q�3�N^F�Y�PX�E��`�r��4p������o#hR�ّ.އ%�p<`�����ܕ ���F���88����x��ԩKc��r�3� ����y����mCLۥ�fu1U�.�\{��N����k�wr�e�������\yO"�L��.%0]lt�p��x���89�WdC)�;/gFחn���(��ᆔ�s÷�j�]*{�ٻ$�
��s�V�w�3D3�5�u�5��]�jjr���syR¦M�f��xҝa%��m�55�o=��Q��+R�Ba*e�!�W��&v�Y��nI .�Нӹ�sS;/t��ʤc�N7y��Ktp	�ю��ku��-s[8�6<'�}g5�>7{�۽����-����g�`~9� s�$�Inܵd�Q�Xwh����0��܋��\|;��p��55�8ڰ�V�SP`�n�K3�F�I��*xB��j�I&u���7$8Z��b�la^��ウ�
r���3�vF� ގ��q�u(��7�H��L���Hl�'k��)R�â�5̓�a7R��T��g8g� �E�B�y�n�`zBrv�e�,=�y��8� �K���U��l�f�,�̲vH��.���T��m����P����p���uO&�ګ�=�	h�e'�Qe=�N=Ԭ�n��Ňb��8!��ԩ��ٽ�.��LǢ�p�6]�Ӹ�u��=��*q�s`{#�ض�ŷ���Sk��/�F�T�[x���3{F�S~+��;q�.K�v���Ԛ�Bs�1�t��L��U�#�ۢ&s�2�$��qR.��_�Cl�tDE�;:dV���*�Gnt�5!�wզk�C�&��ЗC7K�7t���oa�����,+f�mA9Hz���]�]-p7�R5�9�2����
Lۭ�_�=�۝��qvi��A�e�x!w{n��wӹ)����{NZv�\8�]�E������\���!�{���0:S�X���@�M�H�у�G��7݁��P��<E���X�mozs��H�"�&�e�7]yvq[v1���#7�lê�B὚��vV�
��s�^λ0u���ԢE�r��C��4�gEp��u6��9xc�:�<K]7J��;��J�A�wu�s�D���zg*&�aY6;�� 4S��Ȥ������̕��X��5.X{Ec!t�M�ӥؕ=��;s�˗}\ƪ�4yާ..�&vՀή��Q�0�MὭ�gm���l�F�K�9�A�sD�-������l����"w�f�B��7����6˔��1�*�kviĎGz���m�ۜw��ڤ�p<8�d�\A�eL ,�	{�Wك(Ã�.���#��a5_r|8�p�bW��$�ݚ�Wy�i�{JZ��3�����'���ja��Im%Y�w
���0 �3�P�1G,�p1������X�B.]�M��oe͛��%��lX��cT,���u� ܁�2^|��.j�`u��)�����^ݫ�Ñ�/M����7��E�A���q�ǽ�v�߻�I7o>�p�5c��8��pF�k�z�f���Bo�to�E�Snѵ]�]��j w�[c����_Lj���{y�	�	������V��G�訯��*fp�Il�n
���黯7�����QtR�ZG�N\*�=�ɺ{��&ZͰ����@զ�ot��2y��;���+�H^.�/on�ײ�����ꌣ^��r����׏_ZՍ���{�.q��fɶ�5,�y���ŹuɁV�N��d�^7ye���ݸɗ􌡯�ʰ�ڦU[7�hlj�0c��7�\�����{�pHt���hgHD��;Z��h+:�Kn�=�ױd�j6 ��h��qw���:���9	��ٻb��{C��n˅+�_H���I����k��&�ס5#t�2�R�ʠ��b:����<��vt	�s�\��i����"v�Һe\�:vh�b� �ӽti����Ѯ<S:i/�.�C���8<F�ZPQ��I�1�"��8./y+�:�ůҴ���P_�� �&�*{�&uv���xM�.�N��&����3��j�9qY$�on
Ɩ�Y�8]C�G��\Op�Pm�����B���b�o6&��{�hژ@�)�I� ���-m��"y��Z]r���m�x�1Fҳnk�h]v�%���[w��o��H� f>�q���#�p[��ǫN��|.\s�=���'qn���6Ǽ�H�����F�D�fD��"�ۺmh�HpIE�X���.��'�݇7�Z��;�=����X��Z��Dzo�5�:p܇�Ǎ�����kb���ڵ���3�b��n�.b��7(cߪ���@��j|<=�B��`A@�
��,��P"�@�B�`H))	��J�	 � d���!BAd��Y d�@Y	*BHV��$X ,�H��H(IRI$�(
I�$��,�� �H,�"E��@P$!P	`a!�H)	"��I!
�
������ ��	@ ���� (RIP�� "�	TAa+	@d XIR�
IP!P�P�H`R�a$,!	P*HR)$+	%d�!XH	 �(@R@X����� *I , $Y$�(B���BC�$ I?w�~�y���c?�y�]���{U�=CL�N����o��~��������v0���b)pwr7=�E7���HXE���$C�f������$�+ ��[�4��r؆��z��+~�G7���mmiS#������;�����fj�ξ���dēDYF��oe~^�{��d-�Ѷ�7���� zn��Vq��p�է�A�N��Bln��
Fr���Wm��:uPo��Y�ެ�[���5��gw$8j~�w�p��ͣt>�=H��~g��_�?u{q��z{�HsU��%���%�w��u_q�ӹ{6�@1�~Z�C�7�qEŕ����{Y�|}e��,j���N�����=�ގ��뾗�[�8��p�N���@X�޻��/ֱ���������������G��Y�Νٔ�NZT�//1��T�j���Aox������+,��Ʈ`Ӊ�ݺ��xgM�5�o?z�� ��uEp%ǔ^Ҹ�;ޏn�2P��;V���H��C��:0$���L�)s��`���~�lG`�����)���-�2�YzN< �P;������מ�����4E�ӳ3���ը��9�8L�Y��;O�l�a��.��k(�s��z�7*��A�<��G���l�{H�s�"�La��[{�Sm�/���;�&y[��z����H��0��_Lqt�$�W������AM�^�ؤ�w�^}QR��ۨ�!�ܬ4�G�z;�{�FY8p� p�5��.��ͺ;�������Լ6��\#��5�ƾ�|j�T�\��sW����pY|��:���,<��Ӵxԣ�?�=y���s�[�D���t���SV�}�N�O<_�)�ߓxV4�k9��J���v��y������j�l$�=���Ք�|��x���y�˭zxݛ$fk����[��S�vo�_xW7��cr���y�A�����W;��Ǜ�fOe��%�/�-ENg�{��̗%�4�������5�qb3I3F�s-��$�ݻ�_Wբ���+��^�_��8���o�xk���(�c�R��b��1ݴ�	�;�h���6�ޗ���f��6�  ��Kv��9�[J}���Yqw�����_�u��5D��0�d;3{��^�kV�9֞|��d>���+���z[s�ڦ��qܫl���ղ.�G�����s��o}��
"��Ƚg-"�+�Xq0糜�-a{���uv�cw�QT�1\�5��B�nox���^�[�d���O�i@�!����ʝ��g��{�ط޺@�X����Hbׅ�{���u���ٻ*=����,Ǡ抹�,�x�V͇6��B��'9�l��#��JW�Nаvnr42��彶!������{y�g���ؤp��cM{p���n�;�Y��kE�*<7H��	�'�t�Fy�5�����Ӆxb�Ws3�w�u�s��㣄䇩��>��Y}Xo��cq'���9׹����/w?r9ɺ�ݛۻT6ʠ����1�}Ǭ|3�/h��F����/x�|t��t�������پ0�5L޺�����W�+X �{+i�^����Z��7�����d�T�����4(b(���}F��H�^������%^��Ix)�>gȦ�/�x3��;w�E3m0�� ��Z{��H�J��~�t9	p�����*��^q�.h�ϒ:qe�/W\�m�������Ӄ�ק�z�I:�����W�@��8����@9Y��`̘��8��%S�n�i��*@��b�U���_�?���x�§A���x���G�>��S�����M[3gew�y�o�>;�����\�9��ŇS>@�o��
'@s�U\$������tM1��#�/j�\�A���6��u��h�zLyw�K,�.��I�ӵ�p���a���l��p!i�K��e=���{vw��ͬ6�{(-�'8��:���g@��WI�O9�9�;%І��Ɯ7tU1͍���y�{�˧=�Qkے��R�1�C�5�N��}���ͅ��]�����L{ގ��D���7�I��[�o�f{�n�9�~�h]q��sq���묡�����q���{J��=R�u��z�[��.�K�'=P�)ܭ�Re]�=�ӻ�����~����-9- �A̽&{�/Sy+�\��~U�㽶cv3����N�Cxڳ��=�K�c�8���zy��q{�k	��1��̜�P�J<*ꐧ��{�*�n�!���w�����������Y�^�ـ�'����%B7�3/���Zoi��׀>��eoȈ�y�5�)�w)׽�$犸�j>b�rnG��v�+_�<Z]�[��s%���G3L+|Hj�}={`��:�����F�ʳ��շ�,�)kX+���S�v��-��pY�Frj_��fZC��q����!����;��Ƚ˖������{7�0om���S.=�Y�nS�)�9��r�8�kt�P�o�S�JѸ��)��=S�
oqU&��6��o�L5:r��L��Y��(�ʟ�.ޘ�e�ˆ5j�E���s|�=}��,�7j�7U|�z�(�]�k��m݃U�#�H$����mW��������x��\�M���We:�q�̴�P)��;�IG����JΘx��s��׮�n�͒x[=�`�^�mZu��y�����>�c/�j��5����)���<V��z��
)| ����uM��ӷE��Y��}XԞ�/{����C֩�������T/��;��g�=o�1��ǭ��W�ƞ����;���{!�l:F�<�;@92�<�����N��f�P��q�{����ٝn�^^��h���fn�{T�ڼ}�������{`���5��z�g�G�|�sG�cbuF�!��
9E�6����a�F���=�@J�<T����\���=������z�Ո%�~��E�\\��[���"I�ͼ'+�yN/��ɋ�w�e���I4w�#�5S���S�<n,91�B���F ���ӈ��~C���܇m���T�B��)MN������
n��:@sWu��;�tKR���ɵ/j���zxj�|�!��~���ʕTr׎��g\�ǽ�,s5��Y;�wR��mڳ���.㞥fЇ{����k��P��+}�y8�q5��5vq7��QF�&��4��2��&�]����g���14�n��Fy�Lw�)���ɨ@��]�T*z���j^ܜ��o���S�]�۝W��8Z���nh�f�<p�p����E�w�
�7�_�R8P�78dV�����%��әV�i� �ޗ<�s��F8�H!�r�);�cyA�N��yv*$����6rz��/K��|s�����5��HV�=᯦y;f��8����ҵ�o,v��*�|�L&��v.��8ۓע����YQ����ro�}v!p^�x>>�lw:�۪v�
�gZ�]-���v�d�c|7��_��${�܀��XM�'{�ۉF}W���aW�kd�~L>���Fw5;J=gF�p�p����ϴ^�{�?z�����wgb��_`Y��c�,�8$�W��0��2�z&/��rw%�]{{�o���l�6ݦE᳚Ζ�M��~-��gW�������{󄱨���A�^K�`����K�:(��N�f>Q�S����(A
����/������!K<�a�N����Wb�}宬ݚ/�S}�H�&oL��yG�87�?U����Wn�D���(�����<���฼�q���m�u�v�F���:3�?�(���{�	��{�7���m�X�+�q�m�xl�d7�8^�qM�+����F.O>T��,<|�d��Lg��]��$86+����{���^Q�xPZO�5� ��Ш�Ow����(�����j����s�d~�"�b`��V9���,@P����N�5<��fɡ�c |U��wٕ;�w�O��wu��x?A3��{<���9����>����>l�'�;9|1q����g|ǖ�g��O���l:/�i��p��h&��=쪇�7p�H�)A1ܯ�?.P�r�{�b�矵X��[�.�~���PG�9���Xc%��u����>cӷ�o�]I��~$9���LKR��ѝ�M8�z���+Bh��ۋ���+�岰�qۿ�q�_<�,��>�)d�fl��<���;�K�Q�3���7����A��T���j.<���v�z����9{_c8V	;	S�t��o�!N�������>�Cy�\�S���MG�B�ԗ������]^ÑF�V{�'��[�x�!8�p����lܽc;�0T�x�{�ȿ�����|��/`��!;�p���{æ6�Ɓ/bz|pX뾕x�d����1z�%�l�=��oOi��q�W�۴���k�f�b���.pN��E ��]u����J/k��A���@�$��XĖ ������s��S�z	�?~��������D/f�w����5��7�j�.l��D�+ǃ�7�,]�^N�厠qf����F������PT]�,���<m6Y��l䮂�n��l�t�{M>�Ehm�C�刜�y�\�I�E��͌f�]�%��.�_a2��ǒȖ������n����	L�Y4����^��� n/ ��O�4�xof[��.˻���6�fނ#�Q'=�ǣ{\�LݻϪ���x�ʄ]ǁe������<�X���'�8G�+A�c���y��}5zk�uėߧ�+M,�d��!���=�	��h]H�3(ߩ�|���<8s������A�����Z�n�ܴQ�q�7��D���L���U%�{����K��v���4�5}�Ŕy��"󳗚�*C���j.w��m�Y�E����ܹ�PĊ�8�ٸ�����q�=q�	l��r��9˹�h�;Ľ����\y�%=dX1�#7U��߮b�7@����T��9�N #��d��"Yz�I=����R��[wAI��'�+����C��J��a�} ǽ�z�%^�%b��9�r/7Խ�K�k���ǫ����Ɗܸ�ټ��Y��ү]j�H��pｬV��ɾ�}
?%��[��wv��U�� 2{M��Q�[㳏z�Wm�f���}�.���C��g�x`/n;-�Uj��㓳ݞ~�J�����t��))�|۶m����4<�^������K���mg �7^��9��9&O�N��k}h�}��v\g�x�Lu���{u�p�����޷����8nx��/<�㖌' }���F�T�3פ+������ ^���ӄ�ыM���u���>2n�6gμXcz�:\*�g`�.{8?Ӭ���c�;;{���=i��cg�Oh���Oz�/�u�컽� �9*�w�e�%����;����	�SW����DO������E��,�g6��`�U���؄��F�,*��t՚ǭ�'il�0ݘN���!��vd�����v��g�o9:�����0m1ӻ1����;�b����b��,��z6�{-=�W�J�G���dg^<ah��$��{X�W����<��-�g1�.�}�n]|�{ޘv�l��.�c�}9��x��l�9Nk�fV�vprH3�[WS�|8�ExO_�R}2o��e����
Q�3ȭ��on�ll`���޽��/m�cۼ��$�}|ߖq[���[�ٺ��c�~�	ٛ�Ǘ�{Gy���+yt��y���V�:�v��+j
��h�u�:����W7jc�'��sΞ�/qt_sa�w4M\^�}2������;=E��ɩ�Z��彂��7��Gl�	���7Yt{4�ww�m(���݋A6������s!�&ӄ���"���+i�9!��j�f�O{c�����Ϸq��}dR�&k�{8��Gv��f�~X�ø�X<Eޘm���<N��k>X�:��Gj�}��^�5|UK��'I䓄�e����z�b�ƕ��i�;�=���ʁݸ�f���%�s��t����ǩ8�Y�!m��uwD�{��{^J��y�l�w�{�,'rx�;��5N�4��=_LMA�tEx�~�WhՋ��OS��NN��]��9��d+��)�����|_q���w��g'��4i¥�i��X���Q�h�,�MŽ��S�3u���t��>̨.��û��yݣ���d�e�C��#�	V�e���i{��e�R�Ü�A�b��x�|��(��x���Jp{}9��������W���3
�o�Z~�w^v'����}����������B
m�ܕ�9�aD��c����������/��ΒWm��|�y�+q9!���Ra�������K�G��D�
7���z���>��^���f�\_m�{S��e�c��fzH�A�,�r��`��\*�'������/o�Ko�ef�w���{l��-�3�2����w6�9�:{�]��pyU��z��#�uu1�Մp����5��.�=��ډRL����zM��ӻZm�##3�~�74�+���
�5{-x����鵱�z	u�-��ܝ�f.�B��v�>'6��/��6��[7ui3o��<���G�-c��2�](���;�oL���7w�ҩ�vn�[`����:�z[�w_�^�����m�SЀ�g��Hۃ����9��v�(U�Ya�[��s��=&���� ���#�xH�G$#�����=a}Y���Uߴ�N�]\���/�>~�8N5B�^�uW����G�u�5����ͷ^��T˝�|���H@�r{�?���mU��U�mp�W���fz��r��Տ7�wh������8!�vΔ�=��r�+@�����Xcl1�t����fܙy��i��$�z���fq&ڍ���F��\v��J��3�q��#m�\O1��G<�8��
mb��ɮs� �R"`<�;v�#ۍ���v��;%&�\i��ZCkn��뮹�v;a��ɖ�̔��,�y�ޣ��nh�����m-͆�l(���+]��!�|I��8�=eI��c]�\�[knl��7g��&�!Ƴ�c#Q4�s�x֞���	;��룶,#[�����5]���y��;G��oB��nm�l�]�^�ս9{u��H��֓��B�[w�ʈ��rz��s�r�0ڳ�m��n�3��H�M��m��h�M�.3A-F7�6������N7n$v��l�oY�@�GO�w5�d�/;�u��=n�*T��W��J���]Lۊ�nҚ��KAn1<���K\\�k��������۶:�n��p��;b�/�;a���|���H�^�s���e�/\����^[7d�^�ޢ�[pn0G�ųQ>uu\�mnޮ�'m�{�4���s����M�t�^��B�X�y�W��Z���m�m��ѭ�t=��wQ���v��18��pٻv]��@\�<�,A���!���7m�mu�ϟg7���r�������N͹�����JH{n`z���qP�Gu<	=Ct�6����Ő����k��α*)�{7e���H�rJg�vv��FVz;oZܯ'7\���vyq4yq��`�짚�]]����6��]oc(�6���n��x�N��kv�K�;'�;��eP���]�l��v��2O�=v�`��'8�9�g��p'[��wgq��u��,nM�h�������2�s�+�3��۞��V�4�N=-p�HWn�vv���r=�����}(u�\�v�sF�8;=�;n�=��ǌ�=$��6�ݡN�r�<b�cXv����{-�� ��GkJcf�B�XG���n����f���&��8Y�2�Ov���m��p(j��Gg�kC�w�=u��\)��vq���a�<��l�c<��Aku��κ4�>޺w'8��'�x9��Wg��8��.G�N��c� �H�Y���5]�n��m�ry��Y�:ݹ�ۋl���܂��Gx����\�S/�gZS6�q���&����F���V׉��x�nݺ�i�����I�7[q�Bp\og�x`}F��synv���5��8F��H���vE��r��PB���;r���6��7+�&9z�����])���܍y:1n�ոt�r�hg�V� �ƻ,]v����]��c�uvE���a��r�۶�;k���5�q��=)�6�9��B8�t�ո����^�!C�G]�"��\���,��[�/=�݋�v�;�u�Փ��7,��^{[8�d��Y��y{;��zOC��g��熷u=>9:���!ֹ�Ƽ]���{;i��`ls�N���sm��u��7W�7x�nܚ�n�٬�V�;��m��d�\3۝Č9�v�;Y����Cr�`�[[kc���;l퓣m8��3�`^���z�p::�ۚ8�s�G�����$���b���n;q���gs�vtp�J�*-��1�=�����m۔knwR�7Qv�(��<�˽�kn�i�m`��9��.�������s�6�6��ip�E7m۷IX܆8��e�w�{�<R����/��.\����t�(�1�Vy��##�m��LY�FKb�;X��^�Ņ�y!w(s���h#z�a��Ds��[	7���I;���̯O����:�B݁�<^=�:u\�.�y���x��G'��N��n�vz(�Ê�;#%���mI���z,6�Ϸ0/��&0=��srGc���'6�b���@;7{q�s��9ѧ<A�]�@��^��M=t��	��N�
ɮ�OW$%����>��ټ��ܜ��g�y4lU�WU�ۘ��n[`��GG='gk��:���Gj���{]���w>+�\i��18�SF���;�[t��<t+!�s8�So���<���a�L�a��2���M��sA�h�;teE�v1n�ّ#`�]o@�i��5��{/�&�s �zݎ7��(�"�(ϥ�Ft*o[c�q��]�n$s;���y-��b��Zڽ��w���M�x8�>L�Nyc�۝��Ogt�7i��P�M�lv�ۧ�g%o;�%$�Օ�]f�ی��v�'�9�Wh������<����}���
v��5<\"u��ڢ��gk65�v�ݩx_nrF*�������-�DY�n�G\�q�W]kb��S]���� �㓴���Y8w7��x�^���x�D뎷 Y�&|�q��=��t���2v������K�n������k��mg�m^N����hB�r�.��0���穻s ��;����ۉ�p��R�����]'n'���Hܰt1�gq;[����q��cnx�7-ڧ;rtl��W*73���/\�yu��@<.��3�ٺtr���]˛7v���1q�{U�g���\��:�9�su��'���me�cBn�s��n-�D��!��^wH��ggu��i��w#��kv��H|b{X^�k�K��V�j��t<�gM
��%�c��<ٳ�5��yMq�;!-#g\��]��Vs�)��ˣ���F[nv��V;�}�������ׇ�Ny�B�ym�'h�_ jz燻>穗�\y�3��v㥻n����]�긃��������6�ݫt�8��\m9����-n�F��W<�%bÍ[m`�{qoi@ru{�י{��p����mh�p<��b�v.�����=[��n�n�Y��� �sͻ1��<&��/΋Q�����D�5���;n8�;��c��,�]Ou��.�)�Y�`�@ �!�5�K�c[�n�c3֭!���k���Ў+�CR�λk�m����܋�8����g=�<q�aK��ȏ��������ӣ]8��p���Q4rVκ�n�Ћ����'!ϙy�hoc���ŷn�OR����xv��p�p� @����[O�uۛltm[��A��$73ً�{���]���D�dnb7 q����uu�u�)�{c�1�퓨!������Y�G�X3ev�u�v�A�m���<u�:y�ݘ�z�n{I�l�u�kq��pD��n�o۱��Q\��oZ2&���N� ��S�%��N{s�[���rv�{��/3htn\�5q�Vm:7��/;D��9z�Ќ��A�^�`͹������.�0n92�VF������rc����(h��j��;]vs��d筝�x�<���].�+�xv4�]�V3̇r�I�d%����I��(G��ۏ�Z��f{fٌ�A[l��5�q�;�v�W[au왷m�58��îv,����������mv|s�>ۈ�%�x��cp�q���wn��..Q���rd����<�0sinG��b�tqۃ3�v��3���|h5��v��.;����[a�.�h�g�ɬ�0'���q�D�ݮq�u�ܛIm�P.!x��"��ԋv.t�Dg8�lw�N�j���t݃�q���
kѐ�k�%���ڡ����q���f*ׄ�u���;��5��+�X�G$�<�jՎT��`vy�ɻ}N��x�z��7G=��"�Ț�<��loJ���ϖ�w�b�cFJw����sru�w���غ{id�x"|�So[^Û>xn����m+m����-s�k��K)�nxz�s�;�1�Iq�7\b.�拇vpq�r�s�;s�to[�/-��S�mpܥ۫���ޤ�kP�P���M��:�E�y]���w�v���d��mq������p�nyМ��i7"�Fz�pG����Y�9��v:��t� ��cd���nT����#�n��!��.v���^�M��/j�D/a۞�'j
,X���t<�%�!v�y���$�y��f*۞wHn@�,��^�����.��.a��*�1�F�n�$ti��Lܼ����S�ڢ��9����6؝�m`��8��n��p����y]z���V)��e۞ ���K2�ԴV�h�6B�5���9H �1<;M�rπÌ{:q����[bk��U�u��l���%���m�C��q,uu��*�o'mr��N���v	��83.���6q��8t����+�m��h�c�"ƣ�(W���vn��7.�{sO V;mݮ�$�g�9��Tkruq�p]\u�������v�m�\z�ĝ��9;vv�%�q���mb�힘�#�Sƪ�Wns���ޑ77c�ٶ��=sb�yy�d��]�OH�p��kOm��r����,��`�sxs�9�ڍ����v�pAӆλn�W,^��y�����s<v�ؽh������º�&�یOF�4�VC������a�����{pY�eKo	ώ7clc��	��M컀���b�y�T�NL�ig�=��Nˑ�g�{v�v^^�)Z=�m;s������ݷ]W�Cf��v۞۷��C{g�7<��m��,m�k�q�MZ=������:�]���G��K�u��=��z�[�&p�qn��+6�n��]X�챬�koF9�n]C����:�Ÿ���lt'k��n�{b�N�iK���m��(���9nC�tq��:Gp�7h��-"	��Ν��.���:�u�r�93��4��s�
�u2u����w��cq�UͶN1²;x1t��Vڛ�^=�����[��{pmoj淳e��q��z��ڍYo]��V�󽎽[��`�vM�ݦ&eMs�m=�����e���tjLm�Ӎ���v:�70	1�ي��"nn˧��ڵ������x>��EF"	m���E�""�m����V�F*�imQ�*�DcPF��-�`���F,��[Db*(*�ij�Qh؈� ��-6�`ŌbŶ���B֩DcR�*�l-�iV��U�`�TTV*�R�F�(���$Db5��1UQ�ŭ�F�QX(  ��U�cR����Eb��Ab�EF*������4���b2"T
�YiU��1���DT�(��DdUTU���X���Q�����Q�DTm��UDTDT+,V,R �Z�H�,ej�)m�U�TQm)YE�lUAD�F��DEEH5
E�eB�-�"������Zł��E���U���+QV
EQ)�
"*�Q�+iYR�F*Q�QY"�Ŋ�EX�QX�b+ �QH�q	$�s�-�-�=�:ݏI�����ro��w�m�ܘ�=.��ur��c 윰o;5�s��׷+�u5]�oGQ�p���n�����wb�Ӻ�/i����n�\g�9y�����t��9�Ns����A�D^���/�v��ջy��y9�쓟c`l'd��'<���by���)�����vpp�U��nyk�����]ӧ�m�M�mr�Ɠ7)b'��� u�)Qcp���N���i���9<��p��lH���:2�ݻnm;�G=���5Gd���>&��;�5����3��e����
Yc(
Cָ�5�26��pc�)mP��{�sn㮽�n��[�H��ۻS��C��p�q3-��=�����­���E�p��ϫ�ٺ��	�tr�n�pcE��lu����o��v��v��0;WYzF&�(4��n0&�e�9{>�99��G�=�q��]�ݰ���{b�[�O���\hqx�7l�Gu�l����p�\]n88ts�T9��qW%I�ыRJq�ѕ���۶�|Ȧd�u�XL�v-��ɸ�㣬;�b	x�2��6��p�����\�W�� �Ʒ'nc��q.[��,�<�m+ �P�k]�&�c �A�O���U{�����p�nj����x΂��P�mv�Wh������g=C�����lݞ1�{F���I1lo8ƧSfΝ�.�1k�^���z��A��3���\g$S���]�����.��|<�Ϸ.��v�^"�;Z�=<a8S������C��ud-�7[z��c�m�`9pk�m���n�v�l�r��|��֯8-�P�ngl�dc�0�ol�r���[.ڲi6�drxL��g��s9�W r7��pqnčո9�ⷵٷ-�q�^��aƵ8oX0��Ne��g��Vtݸ��ݹ���9��c���J�q�7���kۇp@�=m��g�Z��5<<�I��E�J8�ŭ7a��yɞT7&ûs�s��9D��{u���wl;��6�s�pwL�Ns����
s������ȼ�v�vC9��G��n6lD^�<�vr�s��]�ˀ���;d| `��c��܂ p;m�xr���ݞ�x��a7'���P;m�헞;��0��sÍ�8˹���w�3�=�<��ʯ 񓱞�8�=������w�`D����_y�����|-O����lxF��c�UuŚ��^N�W���s�@�VN@6�A�M���鋔.��8��(�:�V�G��j����d/{aq����׸.{{���<�
�����˪��� A��Ȝ��B �ts�$�=4H$��d(��&ك!�2y���#�^FnA���A$���ψ��ِ�����|�霜�K^DE�d��m�j2:P&㷨Vt�9��lG^jf�hBˎ�� �vl�]dɓ�:�D�`�	���X}gI���v3�ו}iCn�r�3Zr���v���j���ܺ��@$����	��hZ���F��X��ʠH���'�������*SQ-��g?������x��n�:	cj�>on���7����������rQ}<�%ŝp��;�8%�v��GktA������<ՒW��j�q>�+��I��ڢ@9��	D9ɨͮ�y`J��"e6rk�.@D[ݚ���f��A]F��@+.:P>'��6����� �P,E��oO�;��
n���`�Ut� ��Ϊ$/��J�-K���
ug�m�1�B.2rgj��/��׎�c�n̈|�'��f=گ�;3��6�5�W^�,m�L#
 (�l��˵xi�]%��b�83�nZ�3ִ~���Ql��L6���Fƙ�z���|窼y�z�>��)d��"I���f	�
�Ap���}9�O"r��EDm�A$����P&��U���V�m�@���!`-A1�P3�}@Q#���x�I��_�w�@�(l��G!�1$C	���T�ƾ���9��NM�Л��=b۵f��(�-Y��q�{l�X{*0�ɜ8M������v�uP$�|窼O�`8d0�M�خqTvz�$��T@'�vg��$��q���0*��$��ݡ]癢�Q�Ѫ��Q%e�ʙ��p*b�d���P�5�� �ܮ�S��}�}��I���g��Ht�Gb�Mm;��G8�e�'n,�c���m�y�`	�&!�v�
$�og��$�xd���˜<�O��e
��OH���\M0^�A���
=U�me����� �}3�@�A]x��|ENa���O�jtd�R�,5Èe��{TH'�u�L�t�pw(ۣS�����j��WV9����� �3@�e���"&o�� ��n} �oNmt�U��"\�F5ս#9\C&+T���+��VLT�#�u�џQ�i�rt��0H��4}@3&9�4���}0������S@�+�$�[,�ʆKrk���O\����0$1'.*|O\�P�J� @'�ӛB�W�vL��ɥm���!-�b��,Ɔ#�ͨ˒;x�ɝw(�9]楡����s��� �(�b
h�	�ʪ$�Vu�>�7�6�d�.�Ts]iܶ'���ĂJ޷>%[ep.!�%BN靪|P���<F�va�ޛ�Y+r��	����VU�߾�:�v�|�oM0V�&���$};�(��њ��ͬ�7����-�w�6�)4aZ�C-؞��Vuk9�t��|os��A>���I�sԃ���-�$��V�FC����3�}T|O�s���e�O]J�	�	&�sk���tte�&F����b�ݾND��l8���sӷo���앆�ByV�9���`��q�kI�ӵ���^���gv@�}�I�
#�H�� YE��aы�����6Wu컭�	�Sa��]���9��ǔ6rs)�ֵ�sF�<�H�u؝����wG�l�]�\nՇ�"��hx���6�O]qz��%�v��)̜��d�iӴ��i����j��d�T�//m�$Mope����\cyZ1[ V;�Y��O^&#Er������
��qv�v>wZ���뇯(�-۱���x�1���E��M-�qͷ[���牵��v3��ر���͹$����|몀=Q���_(�ba���r���Ux7�Y�Pb HD�Kd�`��쓽�p����^'��:�I�)3�x���[� �	8/��f�D�|릉 ��d-�W�����7κką��n2V�A�W�sg���g� ��g��s���$.����r��~b�Ux�J��%p�p؇"r��W� �!":����'�]TGc��Q]q���nU�lo�����wLV�vn�4��;ŁMqs:��=P�p�$Qi��($�[x��IC1�g+v���ճ^$�W[�'pH�A؋�[zv�U@'�k��H��%c�0��4[�z�.Q��8CmBc��dގ�7X���^���z�67AE(�b���Ǐ_{/!�ݒs���u��T�~��'&�Ԩ)E��	"㫪�#��%GL��;Fr3쪌�����B����C��H#"�e	��wt.���3��������A��&��e�&,�mW'�v�X\�֘Vs$�S�` f�W:4 >��Ov�K�����)���`2����힡W��O�<M�]U	����GvNו�5)�F�lD�Ѽ\ �	�������[P����[�hݞ��1��f^��#���D%���M�����$v.4�����Cd�Nyt�UI�ȸ�>��kKL�!�f*������915%�t�w�  .tn =�ـ`]}�f�S����d��b,'	x,f����Т�"*�}92ݹ�ԸǇ�V�ͯ�,}��Vv�/����x�3�MD7E�]��t������u��-�p���p6�\D$��N������\��I R8�O��e6�s*��"3bH�@��ڢM��v{q�̓-M��J1̗a6قS.!?d�A&�kf������ȉ!��xd�EwmU|H��ڠg_e�=jp��{n���*���c�T��l��L�vg�����#�6�WF7[���>��6Y^+[|������{�T(�	��V���cI�s\���^����ـf�-"yY��l'3�{TO�UlF*�*��x�|	���Q��N.T�����Ux9�Y���C�
,��F{�hQ$�U�@�5S���Y�4��mUx��ʮ�$]F�p�l1 C����_������w��7+�@$魑^�1���̌j��Of*~8�<��2j�7f�)D�8 �^��9�!��w?.V=��]�g��/۸��(��Gh�gg�����e�����L�uU�7|(DA*!*���P�f3X���"�y��� >��Hޚ�H3�LY�B��tF�<i{sM�ێ��Z�pLvJ3^�0��wlb�`���2���\6�%2�kj����f���$�˪7C��Ѯvx�㭪%eJ�"l�j�r޹� �y��T��P�aξ��{�`�o�l׉�&��@1������+�l0�A[�A���M���A$�L븞�p#�r�$o:�I5��S���!Hb���9�WaS�15f���ɠ|El��I�=G�k�f Fjc�y��3��"�%�4��bO�>>��ڥ����7����P�A��r �wd�Q��#C�Þ(wf7`٥�"�<Q��J�BM�������u�;.�_��{���g��h��ؽ�^�|{qgp�U��/t�v�R3%$�IAs��c�G��;6�K�ݛ��l�٣q�Rc&��|�T�l���ś5���e��4n�|��|ݮ�r%�:'r��k���wM�A�Ɏ_n�rO6U�m����H���٣;=��ًx(n�F��u��N�:;i�-�e���1�8�h�[��t�a(q�D�:�8��!K�8g����zҺg%sv���WƎv�'Ltl������u�8��X��=H�n&�=�T;;OQ��h���Oo�
!����ʠH$��9�{�v�z�+i�f��b�v�$O\�Hv��q��L��>ٛ|L���ۢ螉��uS`�I�d�$7�v��y�ǽ!Ҝ�n�D���؄� &�&��^�H=�=5�A��x���U���$���> �7�v�ф��,�������:��|l���>3;n|I �Wt�W�$lv�;��1lk#]�@$\�¸��$1��z�z�Dz;�h��Ќ��k���$ǽTO��Bf3/�U��w�K"F�����+(ЊDRqˮ�n{I������ɷj����)��h@$J��:������̧ �I�}�D	��������^8�܂	#���E�\(��D*���UM
�/�OZ�O���MEڿ�nφ��N���y�9�=W��ܦ6����Z�z���#{LT_L�bf�`�M�����nq�$�B�V����|�)>���K������Hx���7� ��zl �$��轕�4	o:�ĂV��P$C�#��	�@M�MW���Y�	r��_K���$�|�z�W�=S���θ�,i�/�@��a�l����0`S�|lm�4جz�j�@��uD�B���q��J&{gY����B�U(�3��#��Sȡ����ݱ��ruv�ɫ��v]5xV�p��"����ڢ	wuMH$uNO��/3�B
�'^�P'ĭ�9�d�h�0!����r'��n�����vs��O�w�����r�%�3w�tEn�w���AA�b 1Te�P�I��r	�a���1��I�x��Do���0�{}��5����.��޼�q�����Z���r��Wr��d�x��G>���U���7�3�,7��\$�N3�y���@͕���$����!�5t!z^Ǔ�G��l��/���AN�		sǼ��KY'�>)OLc}�>c�)H�0���]�lů�z:k���7&��91����|��pg�# ���3���q�)��t��We's���:�Ǵ�/=3�B�^��b+��ivN��ٌ����S�[��R�qE����Ξ=<�w�9/]�g>m���p�	I�ːw�z�c�]	{6G7O�#.�)1�,�N�,���?or�ze$�6�����ګ�}��O��ZmۜF\ъ���c�1<�b�F9�թ=ȝ����&0�s��s����]�
����P+�o}��C�g��e���ٳ�ژ��w�I���cj��M��y�N\#bC�Kn��!Փ,�x��w��}�:�c1	}�����V�ϸE�֦@CW�푩 U�^j�uT�	Շ5c��=�fŋGB���K�N�;�r=����������$Dk8{pdX4T��`��ω�~��4�dg�[8)���	���y}��Yq�Ca�ͺ	݇�G��)�S�C�8�[��Ϥ0�ҙz�B;}0���Kp�u�y��B��'z������}YC�y��B�5�]���y�����x�ol��a�#Ngv��=�wݨk��H�9����I�w'7wq�C���ߐ��bőH�F(���1FEA�TF*���F(��#���A@PEb�*��(1�(��"��"��X���F,���X,E*Ȣ���EAb*E�V+`�"#Eb(�,b*0UQH
���AAUb�b�����UV"�
��0YUPEb�)YH(*�1`��Q`��UPY`����R,R(�(�EEEEU�UVAb�UTA"�*,X"b�E�Db�"EX�X,�A�*���QDA�FH�+EDEV
��1D�AAVE���,X,PET� ��Qb�*�b�TQQPD��X���bH�
0Q`��b+,X��PV1dX�`��Q��QV
""�X�bE��`(0Tb"��ATPX1*�(��U"�"��,��T������>$��>��V���K2�82T��f�3��]S@���H�N����P�Í����$fu�
��NCbQ ��5^+;�}=�Qt��o72�9����I ��9N��Э��2�S�ד,�R[	8 ��qΎ�:v;60��@9u�{8�C�X�g\��v����M �ˆ��fUI��rI'{�f�VgS��!�Р��rf�r��$R�Uk�����:��Mּ�>�	���I$��H�A#��hW�8�E�������7x�6��Pbώ��>$�쭯Q��s�kƮ�ʢk�H9}NH$�&�ٞ0�D*�rr���ٍ�1�~$��$�A7�]TI��n�����+��zL�<�f�a��?��n{ݴl�O{|}%���X�%�p���zH��Ƿ����b�4zOK��H�ltd�]�J�LX*p��3�v�D��X�v�V��9�VH�׆A �ݭ�'�'%�5,onƣ�z}^Q�ʹ^PXS�J�� ���0Mp��nx��n��y{9��G:?���~o�rB�l�g�݌�A>;�]"����ؚ���ܥ�O]�J۵�@�S)@�
e�ʉ��ʯU� ��=�Ȓ	��ڢ|H��A5}1׸C��q�b���=D8�H`�t6y�$���sD�O��Iƹ���q��<	���uD�۪ �����J
��r:��k�����N�������$�d�]Q �z�+Z�{p��%�4�ٻ�^�6k�A&b!BUxv��P�A�آ\��J���ɢI����I�YS��;7b�`��G�:ٸw2�����Jib�ۊ"�֡%�ի�m$�ǁ��ie;����w���+��M����ʁg�#�[S3��ޕ���4�8m1�gX�=�x<Mth6��@�=��e�d���u��7C��@�n����������J�-��o��'6��OgQ�핽
��N���GY'�����ۜ8�c��8�;Of�n5���բ��$���l�秕i9��;rQ�p�εBp��\�ݝ�c�l0��N�\��=��=^�ʩ�q��ɧ�v���1�׊�A�j�I�Ѻx=v�#�5n��c�vԙ;�sӺH� �qK�_����/�k&�
$�oz����H�Ϋ�\r\)���H'�z�P��OC`�1�Y4-���u`�7���f�'z�I'�eLbH�w)��ǟ|����ZB�p�,0�eD�����$�z�́ �ߝwE�:������uPֲUͣ�C�[ �a8ON�Su0,���� ��'@=���n%9Ȅ͘n �����U�d�Ǎg��r�>��n|m6�ڽ��|	=k&`��u@�3c7��ޏ,�i��fP�a3���L��hlk;{v�	w`���4p�;{u���ϧޞ8�A���˪�H9k�`�I{�ꁢz�i�;ބ�������Ӹ�|���P[n�����ܥC�c�
8�{��}Ǟ����E⎧��8�� �UC��W,�6�l�b�=2�4�靓�r��������<ȓ߇��:���#-t�� ��v�Q'&f�]k��Z��U���=Ɇb	l�j�bۑă}�s@���}H<,w��ע� 嬙�I��|f$(�`�ˈeD���7��D�0�.���H�޺�H''�j����;���L����E�-�C���/zv�H==]5�`l�0�3L7�E��2LT;R	�9��"���ڠf�����I@�=
_����ه�=r��rM�rJ��z��/3��\�N�Kk����m�0��T�|r󮨒	=[U���U�`n�;U\�{�u@�3�e�Qv�L�'ž���\�ܓ1��A��T	_V�x����L�r�U�3���0`4J��p���l�
$�m�l���� "v�=�rvJ&8���.0�����M�ˉ�8[þs��/���&��si�����A���0j��5<Žܽ9�ٛ�RcE�ePc����~�G� D @	�;����6͌��d�T9���M��$�3�{�0�a�0�s0�
��9�C��}Ƿ��p�AIb�s��&ٶJ2�R%@��}�h�A`m��F��ְ��澋�����H/���#��S��|�`��ʯ �g��4��2VQ����k&�0�1�ny��6s~�"�X}<�9�Cl7 ����|ɴ�������}��fM� ��).ϟS�Pq%�
�Ip�Z����E��K;��Z�\m�|�<v������M�Z�� �	'È����͟ ������}ɭ������}�گP DȎ�^�f�$�}ӵ>Dtd�PC����hn$�=�ϗ�q��1[��30�
�>o܆�IA#����k;�#D�3c������da��+*J�y�o�6���
5�|Q�#j|4<
�
��gԾt�w���g���W�7�шp�Ex"�N��}ɴ�ed���_��ɦL$(��y��ŕ{{ϡ��V�ID�5���M�Y++%e{}�Y���yLe"���H� �G������pQ��yg�aDx$���H��*AH-;��֠a5*Q��ﷲ|,�a鯃��ӚV�I�|nTM<�+�1�bgg�d�}��C�t��4����N\;��J�|K�>����i]ƅ� �����������{����P��}̛C`�������S0�p:��m�q~﹁���T�
����6Ͳy|kˬk:��P;��4���
5�Z�w��S4��P^}���f�|&�MwL������>�/��2]�s�nհ�+�{K�,M�;�Hn0�mq�e��ey��u��LCp�_x@�{�M'P*Aed�.���2�IP����~繆�m�a�>�����z'~�ɴ�B�VVK^]�Y��O��zox�1[q�h��s�d6�<	}ʪ��Ǭ�w *.~�\�I���>�}֠a4 T��YS���υ�Y���>� VZ�v�3k�{��ݒ5RV���|��/��<���C	�ƽ�$�
��Xw�sܛf�,e@�P3�w����[��̾s:�� �,k���X��a���s;{Gݱ4�*0ڟDY���E�����7�y�����΁Y����y�d�&���w���i��T���}�}"��X�[,�y��.t>�#� |��S� �*t��T%����E#�ú�u��v��R�;��̚�HZ�?W���=d��Ow������׃��H,�;�;�a��͌�
���Y��>p�O�};�1s����;@��D/����N�G9�|�}ݫ7+O9��/a�� RJ��ϑN�\鹼�8���qEŗ��ww�(�0��κ��Y��u�t	����H��;���ⱋe��I�y�sӵ7�>|�*e��]�ul�K�y��z�v��a;�J׵nGj���ǳ��av=�x� �Ekf�`���ܹ9[�bn�u܀6�N�S���y���x��I�!y�hQ��U뙌���kb�+�ܔq�-m�:F��mv:qq���9\�<��㳶`�kv�7�����q��ǳN.��kvik�
��\�a��;~����E����CI�~}���T*J�a�9�rlf�+*J�gs��F�:�1����<��rk~ၶ���`k��)x}�}��f��ENB���,��n�a4$��2m6�Yc%f9�{�=�x{n��>�����}�@^#Ȁ��>�y�u��°��@�u�d�Ad�|��w?�.iS����vc�{�d �Q�h��1�4
t,�,�|'���6H)
Z5��&�H[HV��gNg~�w����r��@�P+*o����l��YFJ�C��9�hlIX{��F�JHa��_؆}�~���d6�O��*J�ID+�{�a�M�T
��u�sF�6%`V�(׹��f|S��g^�RŇ{���m�`V���>P�8%&�l��@�H�4���G�����T��d�v��;���@Ȓ����oP��
*J�k_s&�l��ed��s���9�w__������n����$��g��3R���8[��/\��n{cu0=��ͭ��߇���\����� �־γ0:Ԃ����2ke!Rc�ϟk0<MD
�4}��-�<s���y�ֹ�m��%e*u��"��'£��m'
E���&.:�>� @D{R�v����~�ww=�n7�<tO����٬G��zl�I�k0���Or�f���Ňי����	�1s.���,�!N����":��$ O���u�Oћd��J�O���Ѵ�`X5 �����b�Rc����c_Oxb���Ӈ�"���P5��q�0]@�i'w�ɴ� VX�YY+���d�Ʉ,IP�Jçޟz�K��No���H�${�#:��G���eH/w��̚L _��t�~x��4
t,�,�|'���n�r#�����X5 �ky��4�wHV�~ߟk0<M T����y�s�9�O=��.���b2T*�_w&���-|��ķ��|�0�C
�>o܆��Q
��+��{�l�"y�����I��R
���ɤ%`V�+^{�5�� �B���{�m�`Wֻ�>|>=ܴ��M��цSi&T3څN��A�H�'b�e4��bCγ����~���uV�4��Ϲ4�Yђ�����;����B�*%a���s0�
��]���i�o�rm&���+%e}��S�Q@�2�*0�-7
� 
!���6|�Dxo�7z����ry̚����HV�o|���$�@��s�w��l��YY*/�˯>�XV�Ȣ��|%���-��@h��L6¸�w܆�H)*���}ɱ�d��*�þ7�g��v{�~�?�nJ\���*�]ɩ��{6�
��ܟ��';�p��-�NƬ,kǎd/6��*���5UNp�?���{����È�(Ԃ��������}ܟ6|&��ZP�2!�"|"�#�_gH���3�$>���Q�������IP�J}�}�6�paXX s=�2i&)�m��s�L����2���s&�H�ӧ����1�74��%a�g��lv���h�wܚ�H]#Φ��!�l
��u�MJ�X{�9�a�ld�
!��|Ȳ��#�u|���ӏr��y1�Ԝ��#k���uAv���{��B�c���W��=b�8��n����|�-KO0��a��+����$ЅI`�a���7���D�����h�X4y���$?o0>� Ґ�,;߻�a�c�[�rZ�p�q^Ȳ=�el�$��{���<ŷ�q��J�u�rpd�%Bĕ�;ϻ��l*J'3��&�l����^���<>���{��x�?t���$���ߓM7
� 
	Xs}���(ԅ�s��&�HZ�H/O�ח�}=|��_@�l*Q���繆��d��{�d�IXS8��͘�q�����Cl60#�{$	p�;���t����� "<������4ɶT
%@��w�@�S�(�Q��j|��F�cϏ*�sv�:J߆9̾SJl��D�G0x����C�}�S��X�CIѓٮ�ܮr ��U����3���x������ x����-,5�߽�6��X�|����O1�x�I5�{ܛH,��R��}��0��i��ϟ]�zOP�+w��a�aXX w?o�4�hVJ��FW}��fM&.��ou��ãGO�w�{Ps�W��=�qf箌dغP7=Aк��v�!=NTO��������5���w��3�2l
H(�wܚ�R��
�cY�SH>���Ϸ�c�w�>fD�z����6�P����M�}����奧�-�0���]|�@��y��7V{\��j�0�Z��9�JʐP/s��F�j>�gΧ�P�<	��n�:�{�����O�G����C��M���Qw���M�VVJ�^{�5�L�!A%B��5���ފ��ro�{�8��°�
��~�ri �M����k2h� ��]��i��Pd@�|>���+����E���|��<H7��Ml�-�+X�{��P*j T��	���ff|Y�k�s?=�=�䕚 @ɻ�E��O��
�aD�PǙ��}W��=�i��(�ID+{��&ٶM��m=��}��gO6���ư+_����A�<^}�t�Y��> m�Ftt���8Q�V�H�Mr���
ƙ�8�ϷB�ĩsr�:N�0�-}�v��'��kotg��:y��t�c�L�?���I�L�۾D�b����&xx�Vo�<��O��O{�s�Cy��0��9,G�Y�9�{�;�w܃8d����~�|���t�@q!e�1{z_Dx������x�!k�O+SinPͣ[T��J�:�J~�jF�I�z/6;�����G��,���ȹ��������@��?YsW�&.WW]�z��Of���ԗ���)L��״�ze=w7n���쏱{����`m�Я�{��X�P^�z�7��m9�
G���6Tx-J��Ikok�a��_���� p���9���ųvz&�~����gm>��Q3;zś������@��^�$������q� ���[ÿv� {tkn�w���E�j͠�d�&n��;��!��\�rh&�.8��p��K��S��Ox�T����!16�n�Z��UQ�u�cŔ��p���N�� �K��J���~�W���&]�"�r¶Or��O���^>(�om
\��MCv[��1[}�;�8U{:���x������$��;��Od���nÝ{9�7�B,��l=���%<�ظ��O�lx��^{r2�D=[wz)���o��Ԭڊ_C�4N5'R;fmӹ� �DT��=<gzf�}ݪ~T��k�����P�y��}z�֊���ܣi{x�р)f87�y�z�vl'���H�ۼpv�J=���` ��X�QU���
1���QA�((���EX"#TTb�UD�*őAdX��*��V(�E�Ec�`�ID�(���P�T*"����UE�DE����,� �"�Q
�(��*2(�XE����`��1�"*,QT��QTEUX�H����"�1
f�UAeIQAU��1EPDA��-���X��+l,TTE�����*
"(��H�����,dPR-a+�a*E�,cR,��$QAV(�A�UR��
�0R(�UX��(��`��QF""��u�xy�b�<��n;i.n�46۬<�����7��|�F���(�9M.v�KO���\�a�ۋ�^v��۱��ٸy���Ύ�����ܸ;]ڛv��f\��ǯ)u���{]8�5Β���QB;vv77/1���:�����Әء9������5�8���j�;����ϯgv�1�c��Y��c��5�6�Af2�wP� ��m�>0�uC�:g^r����v�ۉ�0�����:Ic���<��t��)��������3���s��<I6���5�uc�W�.�w=�^�tzPmx)�61Q\��H'=uEn���a��O86��NL[�F��{�b���f��'=kk;�۫F�+�v)�Sz��S��Gk�3�-��<g�Tx����n���/�/';����c-n��F_)�����9I@;X�`3V9���vv��{lT)������bu,Vō��p�R�/9Iݥw;���:k�c�7[u<v�d�X�sr��LDq�Yݣi�f�1�qg�(
�b���^{����\�!����ӽ�g�[�%����㓨���ǝ���v�<�]�`��ܽhO:�Y���s�\���v�[����ڞ]�<@8k<%՝m��;6������c:����^@j��n��N&p�3=�ct3��yۮԅ���'�����$�½k��ŋY�	&���by�]�nQ�x�ɜ=��n<�����<�zW�Z���m��.�4�����=�SS�<��ܻ;T��a��V�H]u=��zJ���1�z�Gb�ۮ4t���X�����<1ݝ��Jp����y{[��Tc�H��{0gj�qck]�v &t��˸���ې���,�ۛ�۞���4���z���<<������̦N\�k��m���#s�Of�B��.;�{.Zף�;��jjy6���UF��ۜ�9jgK�ɸn�H���w7F��9�0�1��d��w{���V~p�S��F�e�l`Ok$C�Kp'���@vLZ_F=��4�c|~\���;g�O'Gj1�������#q^8ݹ��۵b9�$[V�rXRݣc,3�g����(��K���띛^��j�8y9`5�8�V�%�6���z��"���n��V�m�p�G'�v�<G���緐�6ϐ'�t<���>6�����re��3dx�d��:�r9�+��l9���[��b^^����\����}�q��C:�y��'�k[��M� �����cY�P�$��{�y�i��
��fq�wN��z�1<��o&�&�VE��su���D�8>jC�E��H,1�w��
C����N<��׾�y��&�)
с^��k0*AM�9߻��l�%eJ���7c������G8�#��F�H$!�|�0�Q�u�c܆�x��RQ
������@�@r;���}.5޾�g;���:%`V�,k�~Ƴ����y��n�iϻ�}�S�ynl5^ȰG�쭑d�y�`�XO�%ed�y�{�L�!D� ��|�9�m ��
��5��&�_�Y����޽�a���W��5�5���w���Ǘ�c]@�V�y��I!�@�_vH�<��NGVT�ZEh�<	�y5� ��+,N��a�m���%@^��$Y�nU�ᎳB�dݦA�6�+�G�����6y��;��[!ʇ.F����f��b C%C������=�
�@�ID+y��&ٴ��R�S��=Ѵ�`cәֱ��s�q���� �,7��݌
�N��E���85�G���d_� #�}�}}�%C�< іi|D�T�����X�Nת\��o^��7Q�3v0)���Ӟa�C��`jys�|���<�u�/�ֻ�����C�W��>����(������4�Xl`��#��d�#��zϑ���l�]��{/|����d� Syzw�߇����F�7��;�d6;`Q�
Zw���[%!iHV�q����w>y���ߠTЁR�VQ>�;�a��ͲT,C��d� YG�n�"�0�(�EExA�¸�q�C��;��]CԜ�,B��~׹63i�@���{�hJ� Q��ϝπ����__�>��Q��|)B���{�6�
�{�[��cˇˌx�@�lI�}��m6�R+%w��EzT�����Z��@��>�������Rm9��ܛI�+%#� |����ޢ �>�]!�sbgH]��u��GZrL`,r<�N�*��@��ҝ�D�� ��a���_@ J�{���m��R
��}ɭ�� ����`TЁS��w~羭��x�&3�o0�6�R
��=ɤ6	+�����ˈ����>�;��@��y#�R�/:�qo�Gê~��6�c*�_����hJ��`G>�s�*�)�+�Ov����u�χ���N����m��C�"�5�s�M�VVJ��^��o&�'�PIP�J��y��>;��7�}]����r��k�5�³�$�Й���*3<�U�Pk]�.��vZ��;�cm�%�*���u1ڣ�r��� D]�����H(��}ɤ�+%Y++�﵉4�@��������[L6���3��1�g����w��Ԃ���]ɤ��B�`V�ﵘM( #�G}ݳ�g������}n�}��}��w��M ��ڗo��|[���`Y��>>�7$fG}C�Yn���;�@�T�^��I���
�߽� e��Ix}�vυ�>����u5	p.��-\gEN�r���c���7���)�5�! |C��R;C���G�#׻[�i�+(�_��(i%H,9�s��L7V����o�9�ǰ�8����M�+%R�{�I��+�\Xj<�Cn�@�B>\��l�5!�8{��c�@�y��k�H[HV�+O���I�
�Xs�s��L�%ed�{�u�z�u�����rq ��i���f!��M�^|/��ی
�!RX�a�y߲n3l�e@�T|y�WX�?{��|�y�w��>�(5�Z�� jj�m!l��~�نݰ*��Z�`��J!�>�@�}W�"����y��w��z2VVJ�~��C&��*V���ja�aR
K��=�dz|�F�M����}��*��km'w��2x�e���#��u9RM���(_{�ω�����e�c�xNw�ti�������f�ׅ��� ��O̬�����s&��=�������[L6���3�?��۶�g��~C�@������+��%��C�ɺ�SBJ�Yb}�;�a�m���D@D��$Y��>eTS���+�C����1t�z�g�y�n.����ˇ�9IK�=����s�y�Kk����9����\?�0�
�z�3��+��>ɶm���T�;�s�H,�;�_>��>�s���
�<
C��~��` ��rGDp���^ȰG�~ۑdX |����5_:�g��=��d�
$�Q%a�{߳0�°�
��s�{�i6!Y(�ɟO�|����ɝ���w>� �ppVA��<�0�Xw\β�`Q�
Z��d����#���N]�ƺB��j^���*AeOy���m�++%B�?vH��<��T�p�Bl&Sa׍��¸�1�C��j��}�a'�T�B���y��7P*T>���F�7�+R߾���4c�h��X}]Y>x�PU2W2�.I�M׀d��&�>d��>��hd����y���;���|��+��a�V0�(���{�i6�d���e{���}�A V�;�q�pk�!_Mɗfz/D��ct�,o��$���/ъ�V�q����2"�T��j��_�D�ۇ��������� 8<�GM��^k��[���]��t�xѫp��Jz����9��6�6xNֹ=�׵��Wl����U��ap��I���.I�z�����m[ی�ZK�v6Ϸ�7C�3�v&��I��zuJ��S�<��x�x��-��z�H��ci��=r�k�L��眞�^���p-�zK]n��Y���N<Tn�n�۩8G����ъ��d�B�ۓ���XS��P�v�d���Aq�ë+m�euݸB�b�g�áw%X��q ~!	�ސ-��!K@�{�rkt���k���gz�SH7G����
�wz�3�m��P�=�6�Xl�ϓ���_.��F�����ЅI�t��TO6�a�����d�*J�O��=ѴĬ
5�c^��7��<
x(0�v�}���8��<|(n� �ANq85�,�>캑Di VQ������cy�PВ�dIX|�^�wQw?������#���D���d�M�Y++%^��7�4� P�Q�Z�&�J� 
#��e\��89�>y��Ox���h���&�)i
�}��o0*AM�N����m���k���������4�2T(����ɴ��a�j��~\y������n0�>�=�
�@�IP�=���&ٶN{���o���>@�T�w�h�AH)��Ƴ��A�!ia�w��v��v���򌯽2L1�A0� �2s�\���\�kk]�Ok�	[�}��c9�J��~���@i��.1�:�8߿d�Af�++%y�1���i%B�+����H,3��>w��>k���y`Lw�w&�l��ed�+�{��M	��}/v�c
[py��@�Vg��Cn�jC9|Ϛqr��_?�B{�9N⛑vqν��
v	����×���1��1���C!��V1Gm[�"��шٖeD�TGk�[�w���{�πO}�+�	HT�����P*h@���~﹆�g�G�x�ȁ}V��9��϶d|@�IXS�8�x����`|�<H/q�}��a�AIP�>���&�m��� ����l�|�7m�h� �G� Q�(מ������l7����n�h��WPRh5	�*�E�=�v܋#��;�t��k����%e+湍d����*IXw�w��I��T�>�̛I��j�o��/��zɨ��c+n�ޠD��hF��iP� ��9�u��ݤ����u�d��!u�[�߽�{��C��s:ε��*T
ý�}�4��J�2T*�̛CbJ��}�u��yek�Jc��'��6��sM�x��56��g�=���[�����N!����(�|�/9�^�T*J!X}�;�a�M����\捠lJ��ss���{�ӕ ��1��甂�hXs��a�l
�s���b��b����cP*hw9�2m7++%foxw\��9|󽓏5�g&�<B�*$�/�}�u��
�P;�s�4�h����>��}�.r&T��혧��=�g�� ]||]}<<��m��4mbVg��Cn�jB����ɭ��H->{�v��_96�EVP��VR���ݍ9-�(� /�ELn�oz�����LӪ���ݫ���c�d��Eش��{Lе�r7$�s��� 	�u��"~*Ae�9�s�c%ed�~�9�I���|����<*�y��C���G鷲)x6-��򈉃�q�G���߼�M�l�eH(����I���k�~����}�z��~ �|�/��6�E}�r�

Mฅ^�q'}��ɴ�@�����W�y���'�{���:���9�<Cĕ�;���Cl6¤{���I �n2���o>� ���q����WXX>j D�*�r�J`���Iuv3�[�,nym\�X�3ڝ�]��i!B-Æ��H�B>�w _��������5����+X�����MD
��û|�u怬�Lo﹘m�d���
���}ɴ6$�,��~p�C�%����`�"��O�Dx�����y�����u����6�P,J�O~�=Ѵ���X�}��R�������߂oz|4�mS�������>c�@����{�M���YY+(�^��o0*T*J�z���g>���q�r0�+
 }��ܚI�
�YY(��߷�ɡ*����p�<�b#���ߤݘ[~��|������[�*Ak��߷�@Q�H� G���|(�Cu���&�[�������Ob�s���������m��6��������J5�;QY4`S\��<�ɬ��T��˵3sD�*ظЩ���	?IY�d�T7�s&��J|�����y)��7P�W�w�raRT*J�a��o�63l�����tr�}� z%@��~��@ؕ�Z�_}�y� ꐴ��~�s��y�_rhc��1İilS�����?@Jh��S��v�B��;=�#lu��z҈���������q!�����~��d�t@��d���yɨ�R
V���a��
��cGlV����܏� V�t�#�@Dx� |���3�P!�R�-@Е�w��!��AHp�;L��m=�\�x��}ɯ�BҐ�`W���
h@�D
�';���m�+(�Hu?1�d`꩑d#��}U�b�\c��q���m�q�}�CC
��T�
���}ɶm��T
�����_�����;È%H,
���y��m!m�{���m�`U�3o��[a�O�DW��?�dY�Y�!�����d�y��&�%Bĕ
������P���,aRT���ܛI����Q�X��}���#����> �
Æ�0�\��<ƍ�n%a����6�F�,�;���[�)�{�<�q�zC��_w��0��@��s�ٸ�YFJ����ܛCbJ�w���?u�pg��(B�#>��N.����N��V�ph�뭚�T�gM���\\�]��W��H{72��oQ�9�]��Y�7�QR4�~��=�䘭pb!�M��H��=�>vR.�-Y�ҚE�qL��u�;��=�b�D�enN�ݞx#m\z�Zǝ�7[�g�vE�N���7<,�l+�q���[h�}Ciw ����R��&;ݎ�Ncvl����E���\L�7��ll���{j;+����K1l�Gh��v;4�I�'!�E�Lqpn�9���u�rM�F(v�:�Z�(ֽ.�V爍���';v�X�C����2vx��i��=�k��5�x�Ja<Ǎ�C��a_�����¤�
��X}�7̛�JʁbT
y�yn%`{�`����yͰ=��9��դR�{�o��ݰ+N߳�DANI�گdYϷnE�d ������fK���-��2���{��oL��%B�*IXs��s0�
*Kϻ�rm �led��3���Ϟ}�{�~u�ϽD" ^��*�� 7T%BV�7��I!�h{�{�[)
�R
��3�u��Y�o���>
�@��O{���m �c%@��(�dy��\$�B.s�G�ς9=� Cg��}��$z��@G��o���6ʁD�{���I���(�ۓ>�8���,��xmV�>l �
*J�i�0b'^ �.;ϲi>+(2VQ���=�M���=מg;����1��y��m�aF%��{�rm&Ь���2���Ͻ@�@�1ȃ�����FAl>f�n�]�Y�^۱md����hձ�9r��W�F�fa��	�� ��|'g�Cn��hs��&�)
�Z����3�	�������'ªw����'V���� ȇ)>�s� �%NN��݅O�����#�,}��+�9����ٍcDT�������^|�+�;�(�ܻ�vk�;Lڹ}��y�{��������WweP���[�cp�v�;P��(�wv-1S0�a���.�*�ͷ ���6�lt�y	]N�A[ەD��&N	��"�p�r��6���\	MOM<O��޹������z2%zv��1�}$�>r��)60�2�w�wĀH7�}&n�b*�L@����]W�$��s�$u��P;{r�2����\b�8�6�'z�Y����]�'���gsѬ���:��,+:�����,D<�0��  }�p ���H*�3}�_�ӛ�W���ےm�����T�TMm�}�р�v���H�޹ we�P'��A]��Z�����$b�PTL��JA��r	'ǯodP�˩�L�M �_dA�&�<B��y��n4U��nܚ9�"�]s|����4*y��ٰz��ˋ�3D5:���>�j���rKs�G1�h&�R�`�;�Y�^n훇�zp����k&fq��]�nyQ�=��x�+�X�����.O��ꡅusw�;�Y&�A?��Y�^��Kk�{�L�G%˄�����y�v�8钷/,��f�'��������w���.S��;�Ƌ���~awgJ�`C)�}H�9��t��V�����&�� >/uwn�)�Q���gp�(�g/.��#s�U���#z���r� ���Q�d��m�'F�tY�am��qș�oI�v�ÞM��[�����7���b�=�a�/X�7ݒ);��dc�os�le���"�QdLM����z��������^�l���޴�c:����ӷQ�Y=���<�W��t��d�������a��[���8ڨ�0�跈9N�A�@{�V�ޯ�ǝ��3��$a/yܫ=���״\��׳^����������y.ݼt�OEʲ��5�|��}#rtH�e�W�8�3^�\�����I�Fr�8�	���02��<�Q��q��f˵;.����m��{�ˉ�yQ��:�Wh�..�7�9�h�+�J��_=[��c�[���#[ה}�i�u�]�S�^]�u�������#|.���h<x�5��M�ȴ�C�9��P�E/X>��ƟEz�o�1=�4}�K}|[�~���
�Tb�TkE`(�QAE��
*�Z�����(""
E�IP��
"��DTQ��(��PP�ŐV��*�1@b��H���H�m�ER��TQ`��T����F"�EUUAH�Ă�TD�h �(,b�,�TA"�P�*"��Ȣ����(�TX�"�UT-���X
�`�*�PX"�ؠ�TTUb�QEQ�*�ATX��A��(���b��(���V,-�)(��X�T*",X#TUQV,1QE�`�#F1UDF ����"��F�EX�1*#+l��b(ԕF#"
�$V,�Q�ň����{�M�m}�A ��ߤ��e�Q#3�i���0�Uu�U7���gs�����=�A>$�ve�Q^��1y<�ˬ�|c\��"V
�L�Dh�=[UTI�Y�s@�h����u��14���	��ڢ|	[�uEj�nܭ�4���RdډM0bl�FV�>���wQ��6˷*5���C5[Жl�8i�x�͹ov���I[�tS��h�� 1u�O��� :�^�S��]��R�7�j-�'ĂGv_UIs��H�A`yl�n���6*��	�pS�/�uz�$���I ؊��{ \n�$�W��^ ��]U�}�-BF4dBa �k��z+"��I����I]��^ �{�t���\U��I�z��g�.�5M�Y� �c�{���ݿR��ъ��pnfL�eQ����d���gR�uh�BFe`�m��͸�x{� h��^䏾�Rȅ	� ��SS��%�ۓE����R�靺�IW��D����[�dV╰{ǫ�5����|D�.yq�c��$�u�v�ͺ�Ľy g��~��߹�f8h�7YUT+��Ex�@wՑj>�w8"��sj"!�[�5�H9Q���9��RJ������ݛ4(��Wmm
 ���Ϙ �a�[l�iQj�{�d����Zp��P,1+����Ag:�2H5&�j��-κ�>%^V�3}rȦlO�	�N�tg�FU���Ӹ�|c2zhAk��H��G�#k���"�(�Fb�Ba ��u��V�:�
���Y"s3���w.X ��6)j{M���J�i��5{9����y��Z�����龞��=� �����/W�Ht��rQs��v<�^�8:��Sza�w��x�+�AJA63��NQ-��nڝ�nS��i�Wv����z�Dbb���6�	�j�6+��	�<*b]�8�8�pn�V��l;�gE�Ic�h�qơq����I��ŝ����霉����k���=��W켻=�j�\����T�����l8����f���rP�r����wk�����;cաm�i�u�6��v2��q�<�X��'Wnʞ;�C���6�a۳��)ʣ��h2�;dO����"!1�56�~���Y����}TE�Vn�]T�=TH$�yq>�W�
0�p�s���UDT�h���陰I�ˁ ��$�}��y��n?�X�FSc�.:��@��Y�i���Ӹ��I��r�Gv�Ux�-(�[�o�����6j^���Cč콪$�]J�ȕm�+�>����xN��	�N���Κ� ���G0�hq����'Ğξ�$�-��]��"Înm^���b���Y"k�׫��U����(,�:ٍ���NwFz_������@��L%�����|r����Jܮ����R�fH{��hs��P�(�Xm��}s�@�~�Bn���M��j|m���W�հ�3�=��^�H�k�Z3բV�%�u�&dS�Gz�##	s�W{�Џ���<=탗I$v�}^;��� ����~�G��4�*����M �abi��N�͂�t� ��}ӻ�ޱ�mF�^_UI�ܮ��)I6Y�!�NEu^�=�{ݒ�UvH�@9Y4 Ѿ�U��,�~'����IRK�a8m� XbC��� �9� ;�����6��sR5��Ux����@�H4{.Z���Z_��Z���c���c�g�ٓ�t�n�"ϣ��ۑ���y���)v1ͅÍ���~~oޱ��q8���̑��ut�Ċ]��e���*��5��`�W���-�!b��x���ճ�K���n*̛s����.t
�et�$�h�\��U»��.[P�k��7
 j�)��$�G6�I�2;�,���&�%#Sӷ�E�M�
������v�>���p�l��X���eܶ�P&v%t��n�Ž��p\tw��{��}]�ĀO���DG��"r%j�� C16LH��o2�u_���D(z�֓fnM�|��Iw�p� ,̺t��"�f �:�1�� �mt�r�6�*4@��ڠI ��$�wmuQ(�S[���3�Jcp�5�{y��G�u;�۫�z��h[�;lq�0�/&CQo	�`��$w�^eQ ��m��muQJX'��a�I�u#�v[�Roi&PL0��W��@Q&���7�A��)�59���Y��v�Ux㪱Gs��7��P's�@)a!�	�S�#kg�|H=}[5�5�CQ����	�+r�H>'{k����oZ���ڪ�ʨ���jr�lg���`��NwV�	������#���#+klT�u6anM��Z�;��Q|�mL������)��c�&�����/{.�ptx�%�QevY�Nƌ3*���K")�ۆ���  �}7�"H��X�8P!���&$����$�e}4x��,��
�\�I���H'c+��J��Y1�b#e���Q�&4of��8�4�-�� ��3����t��g�=�X��g"�ȶ\(A�N~ �{nA&�k��$���@��J�^�}�A�uuQ>*N�b�o��e�P#�[=L��=��͟[յ^�}����4�ۨ�͌�x'd��PHL0BNh�:�GWH����2�w�r+���I9:�I�~�Ϥ�x�X�	c�w�GV�l��\��\�@��5@�b.r�D㱵�^$�+���FD��CC'��9U�H��n5C�na������I�s<��t�can sg�Eo+f�$�+��;⃻�/�o�Ɇ����x�:�r�B�qc+ɩ��͑�������Sp����㛤z�k��J���4��Ɛ�U�;�����CWT@q�0���B�»��ѵmI�v����ݢ��I��[Kƛ�������y�-�v�h;]�lvwn��6o[�VLv�{)+�v�f�n^H��q�#���|\ƙ����v�w��M{&u�+ďYƳa����E��]c�-��G<�M�se�����.�uZ.i3���uA���nݷc���t���l�թ�wȍ��7P9uq+v�)-�wg�����8��𳺝�&v��'b���?}�>�,C16L~5[54H6��kĐ@5�n|A��v#a���� ��= ���&�ƙr���lc�32��j���A c��I ���$K3�OK�}���`Ŵ�x�)�ax�,��� �/�@�Jo�OD�o�m;]<I#_V�	}ni���/5���D%8�g�_K�ʚ�H$���wom6�Į�^$C��[DA�Vq��X��2|H=}�T]'�"�.x`Ѳ�>�˙�������(�bp68`6�CI&�E�B"�jL|�h�s�c�a7;>Kz�n��2)γ���������tٞ�m�W�����>��ڢ�[;MNa�}�|N�W�$��"rU�XlDAU7��q'�Wa���90փX�{�z��e�����6zW�٩��� ���x��a��>��C��Q�:^�ͅ��d���.*w$q�^ے@?}��@�mO�Z�w;���H{�BT�8�uDn͹�}��D�EԞΆ"s�V�/vs��Ays ���У�D��C�D��}\�h�r�A���$�ݝ�(�y]O���c��BA��$k;�Q �/5����Т'�WM�4�\ڊ\*���|w���ovO�^WUW��m��Hz�]�U6|���:�-۳��-��8��p;v����ń =��%��1��?[n�$���
$���� ��Q��ӿ�t� �3sr��;IW��m�-���mNU
��}�yH^vԒA5��TAו�@��n	��9��$��z�6ˆ�$�&�9�$[��|I�g��Jʥ��k׈��-��f�w�[��_'(�� Ɖ
c	|[�E�W�̘ѭ�e���,hc��)�p�س�=� n�Ǿ$��&��y_U�"�I��u@�ٻgN(HD��$�u�� �H���@�}W�%Ӆ� ��"\8�pH��b|�hP$���'���;�:IǕ�D���j�X�f|��>�.����8m�n�=6�Ү���A���s���&0G<
������^�������ϫ��$w�䝽ʞR�V�y߶I��s��~��QE�����/���ձN]�M�O>��'Ă.����C�اS5~�JW��m�a����ʢ@$��䓺;LK���M�$�{[U�I"�}'�5�T&ӆ��a�WM9��:k`^�'$�?]�d��A��bI��W������	�����1$�n����G�v����๵�_�6>���c}:�w�w~6�+����}GT�w� �����Nc��������ķ�uW�|L�Bp�@m�^�]1������{�M�feN A]�̃�{���r\�|�~�����݇�е���W$V�N���;���|��u�k���o�߿�ڈ�۞b��|I{r$�@=��4\p��o��5T�jd�on�	m�̚g�*!b �%�x�}�Gƶu�}��4��|I���wol� �.�+oh.��F��Ba�Ba� �}��>'ǯ�j�$�y��:��⨪�A����c|N�����IX�-��&᪬Ꜥ���"��3�Sz�]ۓ��Dl�W��޷|�f��E㙓�\eBm�p�F1 ���
$�9�Dbo�,���]�c(�[WW��{� �W=��?�4T8|zR����f�ǵ,`NY|�f��ʸ�𺳍bOP ����7N7�U�zN�|/������x�\-wvr���y��B�V_E��@�mSS٨�\���e�kv�Q��-uƿP��u��`<�]�F�s�����E�o��@2�b�_'W+�랋��b�7�)Q��i�K�ڻ�F�w�� q�ӯ��/p�m�w��P_!nӆy���cS8Iv3��n��u�}�����4wa*�s�����n�SƵʚZ*D�QWx\j�	`��v�����KͳV�ꐝ��,|�U5��T���CukC�ʤ�����s��z��A�@���n��C}��K��q�rz��{[ҭ�G�>�<���s���E`�M��A&vK��>�j��4�z�[Ǉe�H�����S٨�%�w���ꟹ�4���l�Q��W9o�zE�0���*�Fʗ�F;��mbM�{@!��e��p��4���4lGg�$o��6��{5xz�%_�'���z"L>�M]EEj���R����o�/C�6i��.���.v��7��i�r�v�G�~�͞��Apܬ�
0o��'��Ξ�6a�;(b{|;�<Sz��l��n�o��4�`vn�����qMu��f���i�Gh��,�����m>}���	�_8x��:9��AW�y1�Nޘ*x[�^:}q�U�%�ouv�K(u�gm�'8��eZ�+]&�{(��d�}ݱ�~ۓ<BaWcZ�Ь��ڗru{����k=Hl���O3x[_B3�3�x֍�APU��T�
�1U1F,"���b�U���b��*��AUA��D(���YUE��"+b�$X��ʖ1EY"���QE,D��"
*�F��� (�X��"��R""(
E�UU�1aPX��őQQAUb�X,P����cF((��T����V(��(�"���,PX��"�"�$Y�� R(�E�b5�,��Q"�Ŋ,��X(��AEA(,����V)1H,R*��R*�**�R(���*����(�X1�*$X����"0Eb�*(+��ǥ�	�:W�b���6մn��W"m����&ү:�8�z:7s��79�"]vsЯ@�v�7�۞f�NwbN��8�O��'>����j�Cn^�l�{���lu�1�|��V�>|~|wd�8�#w+�9�:�nK�d�qgxv�F5��ܜyP���u��O��9�ۜ�֮Z����[Tvݭz1n�fx^ʶ�<�@����>9۷σ�o(Z.��t�g/(�Bk���vݭ�Vq�c�4Ə1���r���n��#ϔ+�:�θui��l[c��]�����^�[k�����]g7C[t�=��Hۗ�X��Y;���=aJ�6�����]��u��֣t`��D�5�4vόɌ�1�n}q<�с��1�uX�\N�]=����tWb��[���8���+08z��d��w`���a���̆��������)��`2�%�hַeqc�N�grk���.���3G; ӕ��ٷk�I���nG;�\�]�p-p���ѐS'sӛf�UĢb���;���]��p��֖#^zLc����r�n��dG�aݞ��d�\�[
��o]��y�])p�q竗�˂�\�Û[�v�t갻�����=٫.�9�K��۲]y�k���c�g$sr��V�>��h�9�]���r�oA;����Tq��w�vn�W��θ�/\7���Ӹ�t�.;b�
f��`ۅ	1�L�x�n��XXx^'�xݻ\�j�x�L�>!�n�;�3ě8-��[�J����⍺��[^i�����6�Y��هd��e�q-��3����Xݹ�m5㕃�B��^�`tf�����v.݉q�o�h�0��-����ˮ݌wv� ����)hg=�[��n�����=�j�Oi�ml�yn�v��1�3���7d�=�9�k�[���N{=��lh��sh�Ya']kv6�9�v�n3"�N5۱A8O�k�o��[�) ۜ\���&����U�ö�n�:����[�b��u�q�LY�2��-������|�һ�����;mfzlZWU;=�GU��9� q�\��u#r��n����{F7�y��m���v��W;�
x�q��f�d,u���F1����ŬA�jۚ���k\
Y�q'1nʼ=��%gnt]��v�]�:1�;��˞؎Ɇ=�ڢ���!�"��t�9�n��y\��;��6�4�����j�q�c�Q�6����6���Sv;��#t��\Ys��c@s�M�6�"�����~����R���b��W�v�4��3w��� ��}Z��A��عv��>��D�y��|I����i�@��.V��  W���,�z���d���@}����@ ���@���Y�}���
+�2:��i
*b)�/��1` Ϫ�D�K<6�33i �v��iծI~�2)���NZO��b���dm�D�W���A}\��0B��}��m�E$�����@n�U��lC�4Kh�^Sh��[M�r�(�{|FY;Y�?o��� V���,|�I9�9�귳c�5Fm�!�����^�g����:�$�]%�Z8%쳛��4���Ͽ���J��M(3�=��3� ��>�h� Q����bgz�p���?{0�I���odPa�CP[i�$n:�U ��/��Yu|.*�T��S
\�KBB��է�MS�G��p`���v���A��Ǌ:�?7�ݾ�1�?x�*�JV���{v���@|�j��X��L�*#�>��������l�	8̨F�m3��pO�S�9?��ͦ���[�{n���{:i����>�aX������L��A4�1����#'��b��%�U���(�����{��ҵٵ���l�=PH�ʠ�R�,��l�{;��ֶ�!
Z��;q	g]9$��2�wovf �2��S��;�x��!�X0=&�x�;�wWcq�g&�۫;�p�6;r�/�۟���߯際����񞼦��>����>A����AO�zS�;ƛ��o��-o[L��� ���`����$���Y��� @���h >����@$�n�b�Fa��tOx�"�
"i�Rm�cm��;{�`Fs�j9ND��a�4j4��~�xq\�fX	�����}-���5nͼ	�,�q�Zw;5��~
w<��k�����*�vI'�7�B�'{{����h�a�p�$YE���}6=C��i]ā��;����٘ ��
���gOFo�HԀB�_6�FW�'�i
%J�e��:A.��4�v�Fd?d�x����q��ݙ� ��e6o��v��wN�yFSa�,�@�J!���s�o��c1�� �ź�.c+V���qX��?�����j"*R�1
���l@ �wsŀ�@}��n"6�{2`�.����'���A��ݙ��6jfj�iMMMl��M����0[~�vT�2�m�� 	{����Gg��&��|q�w�&��j\	���{�I�TT@ETD�>癘	�z�*� �VG(��{��ހ�-��'g��y%�A�A���LQ#e��goc��p�ZI,뻫����6�-�� ��w>��u�q�o�3ۜ�.wF	����Uwb��qxV
.(�̳��΍�ёu�P��j�m{�G����-^�]m�f @5|"�p�d6�ti7�꼒�D���oc��Rm�
��̈ϐ�� ,��i��=�k���:����s��h�Y��Iෛv�KZuH)��x�ۃ���� �퐝B�iJ�R�k����X  ��h�@}}�lIk^��L�,�W]mݤ�9=nh$�^�(C%�iS��>�m�=셕�/#1�7�]{����˸��������a�fr�&&{I�g=���q�M��P]�N�� ��4��DfLGR�ĺ�3PD�ܦ� �]���=�I��*"jjd���y�~���j|{*� |f{� {{ٍ��olnh�^�AF7 $��c�b�Ć�B,�ځ9��]R�^J�{*ūǒ/d����0�2.#~�n ��V@��{٘�`
�bN��-i��K��n�X�	�o�Ko�x�<��$ �n��k��q�r��$�/�ONo8�!��|��/��^x�i����&�/'Ӎ�.��ۗv�9��PJl���7�X��2ġ���N�T#>v�s����z�ݺGc���@��[���M3�䠗��z��:�um���n9�ۏg����gm:׵�=��;Re^1���a�h�6��h�a�%.����Uۋ����&ݴS�V��y׏m�@��/�8�;��F������	#�X�+]��U�:M����>��'v�z�Au��c������߿�߼~拚z�h�yW��Dlf�N�wo{38���W9��t�oi��23q�?��"����0 :t��mѴ���U!W���  �;?�@}���dF|�nۼer�zNr�)P�2K ��(%�y�M ��n0�����p�D0K�~� �'��n�'�UV2�L�-UE[F���2��Q�
�-E�n��;����{��'�wQ? ��y�����Nf&���&�*[;��3� z��l1W�5�=c��`����� ����1 ���l#
�]7�;��LA"����mx��a�3�F�'�5�O	Z����?9���5�!kx�ÁaBL�ځ?%��@��y����p�\���3���H�3��03��3 T^�j���R��"�6��<}�<��ؼn!s������Cu�ILP�Ό�R�[)gfn����j�7�VbvC�[�4.b�!彞��u@�ξ�$�v��.7��L�O�9 ���ݙ�|F�m6T�Ҩ^�Rm��d��r�*Dҥ$J�O��{�0#�:�� '�5km������oD�ͦ���PE� ��)�Ϣ���W{�;�S�Z�A<���F�^m�h�;ޗ����������{��TVZl�5QW��� ���v#"�杕Wq)�}���� �{N"{�ۓ�Aý�E���D��!��@ �&;<�6����ۙ���޹a6��ֺ���Ͻ����"j�fe�3<�3� ���� @.���#�9��YWWٙ�6��	�"Q�Z0S-��Q+6*V��27ۯ;6b�~��` >m�� ����JH j���h��-�oo�GP��IsMUB�U8eVm8���;}-� B" ����&-ǹ+�p�]Sx�c��g7d���`��l>�G��{�çO[HX��i{}^l�
b��p:O����#4R�������k�ꝿ�Atֺ$�{.&Q��0�L�e�F�^S��z38Uvc阹��	c�rK����ƀ���fdu�g�k�v�F����u^KM�(#!�Ø�#o'�9> ;��n/��Ŝcڿk�>��  ��z[rD@�����B1��߹�_���z����J��7ZSqv��k�<l�s�/l��e�ۜn����u���������EUQWǶ�� ��t���|��nҒ�q=U��t�͹$�Iyu�UR7ӆ�O!6�Kg��}/w��u���^����  }��l�`wnvf ޹(�86�[ݯ�.��ޯr{b�B�0MRRm �l�r gns� <����w��F�콎@|��}���"�Iom�ݤ�!]E2[n�aѯ���w�v��y�y������i�W�:���Iu�`���Hs�X��O����c9F��	"D^<�����Ѧ$Gv���%�*���3����y�����,�}�����3�^7 %�H��R��r�����@S궃�y׹>qӒٽr�=�٘�I �ֺ�%Zbw�%����ɇF�F���3�<�j狷k3�N�m��N�)�1�*��LAG��%���'��`�Ks��� �ֱ����㎒��Q~����	��e�m����4��L�nk �ygnX9�����H$����vI$|�{b s���oFe����Ma�J�.�˻�H%��eI���Gn"ȇ���$J��w`$�B:�u�!��E��Ԫ	��
M���۹�t����y�� ��+��@|8�7Y9s��o%����s1B߂J mM�^��LD� A����٭H�+��.�$��&�iI��u�>G�
�p���9��ذ콪�u�B�L7�)���㖰�[�O�u�4�)�N���ɇ�**�ڳ�{+N��:��c���<rt�s�8���8�*�����qtiø<�=�z�:_;n9ٌ���.|����^�Uͺ����G�g[^Ɇ�t�i������(9&��̚���6%�k8�v�O����s��{lv���b�Q��9�Iv�;i�`�.x��5���{9^�79؎{%�=�x�ȁ2��Zx7�+`r��w=1�4�M�p��q��lN���Eм��v�� ��NQ����Ş�m�Wce8]����#���<MF��.����G^O[�H�w����}�Χ�����H�G^O2��'����S	C�2ho�p�����_� u�k�;��""Bn.{qw�=�Oxw1���qB-�M��ۜmI�u�����E�����n  6󩿂 >g6��<�SM��l6���z\ٕ��d�~��>�ʶ D�7L"����q6�h�3m�5�RB��*m&*��j��@��ן`�x����#j�m�C����CA����+�b�3xY����N����k[�W>�Z��Rs���w��t��8~,�A�kP��pD8NO��� � }������Ƕ��
�2�m��)�� �����q/�D�R�3C��|�s0��Yq�lw��#�e5�5���zi@���y�Zb�x-Ӓߴ`�X�&�I���4�s��N�H}��i�U����:�'�Ok��V�z�KyW��z{.X���VI\jRr�d���e�e��uA#7ʔĒ�B���-�u�@Dgwk���=��'�k�.�[�{��@?uA��K�{n�$�k��.!�E�
�;r[��ʘe� {�m�DCY�ۙ�"#�g/��:�rr�6c�P�iP.��D�SU%DUET�i��3 �9mI>��}3s�<�:�wv�ZI#�Qs^�i����g����(!�i��˔����lx(�S"�#q����929�u$;͐���bI�N��I%��ט |�u�h���꾪���x�7D�v��
Dt�S0��*	��Ed�@�Y�� �*����?_�8� ���̈��8ܐ|��<~)l�SWm^aC,Ci�TMv��|�#��[�@ ��2�m�j ���"�<�~�?;�hYl{7.��V�w�<�������]�Oa�QK�ޝ��㦆s�g�IOw� ��f���[�d�.�8�Ά���m�6��/v��p9�W���jhW�Ru�+q����c�/q7W��/m;:ݸ���v��^���&=~�N�9�}G$G������Yc2\n5+g͓
L|���U�	�h�^�;oh(�w���L�<��(Y}�z�.$Es����������X���E��"^��x��U��Ȧ2���aL���g�v p��WA�{5����ߍ�,��-.mC׊�{4��V}dzg�Ge9��.�<;[`�WT����[8w�3Ӵn1����&��6� ��=�X��UÛ����0�Y�s�����5���e��|��@{v݇���8M��ޫ�;x�H�g�w���1��ga�
�-t5��S=��E�I��g����_J�܀���R�Pk��E� ���q�j�o]���9�y�ʻ*~W3�Y���Q�d{_�痢� ,e'�\3wu0�h���T��e�{�gckn�F�K�̙��h����V��W<��<t��W�*��O)tU�5�fz�i�����kҶǡ'fK;��s���-��L��>�13�ޜ8�~��ݓ� ^�t8�d/�w�.�F��`96Ķ���2���,ǳ���9� #W�(�Lp���
F]ޛ�'0�t���t�2Y��sZ�]�h�y/a~9�9�<��&i�N���;6{��
$U�(*���UH�"���(��"���1(��"
1Q�b��FE���(��TU���*$V)EUU"�b���X�dPD�����D�#@al+"��"�("�F"�*",VU�"���V�b"ʕcQUH�
F�b�Z0mej�Qj�##X�¡R����҈��)Z�Ԩ#m��DQkX�)kX"V��(6�ciU"��Tl�(�AQ�@P[lUQ�b(�A�*ZTYZ�(1QAE��J�%jZPX��D�+iUUUEX�iR��*�TT�V*ŋb��UQZ�UF##Jխ�TT��(��aP��(����F(�%VFТ(֕*�E�KZ,YY*
,B�su�|^H��ۙ�"��7���S��L��������}�^���cS-�|m�q�� �:�D?���.���?B`����'�Z[@��!���~�RD |M��҉^����r@)����� �q������zڢ�1q��-V���;�I
���nԞ�=��9��۫����.͈�X�a޾��e��e��z�>�"#��-�$@y=�,6%�9�׹��o�.�$H-ꋪ��9�QF����Njs�����=�#b�w]�X�H�r��D	󘆃<������e�_r��6a�&�4T�8h���T%䗒�]��v��g\l=�wĜ?z.� �~�1�>�S�ęx�(c+�n&FW�c���u�in���l�� �{�Z ����{�q�U�"�^��w�֟����Uf�dwv�6�%��Q�Ѯ��ս:lYS>n���ͼ^����K��H��m�!��d��X%4j���]�)������r�S�*���@.�u�h"��6�I.���qA��sd��AI���[ud]nx��1�ݹ�>k�e�T��m��s�on]�>�oe��a���8 ���� ��������6�;x�cc��_� 	�>�c$��@X�-0�h�$��}=������=[Uj7��z�lfTRH�v�ݒNV�k9�n�'����(�DC�@l�RY��b��	_ok������~��o��OeA$�����I�P�4�P�m8.���voJ�Gv��#�xӨ��o��3 {�ޛ��.��1Q�fz��GkRK�S4R��CZ�ى` ]�lw��N�T�~
�}r���vdF��rOP���(�of��:�Cqsȣ}Ӯ�Q���� w�����}�Ls�W��K˖3[��g���ݯY�{�@ͼ�q>+���8F1��P�u�i#l����P�qq��CK�(1����'m\v����2e����<�\F��'�z:9�7;��,&���s�=V�hū��r��+��ɵ��R�����q��pI��:.�G&�.\q�62;u
X�c
�a�a�N��a�ۇg�#V�\�h����v��z�Kzn��D�O{F᡻k���2�#�ݸq+�Gh�5��$O�Sx��f�p��h�FGu���n���d���g������Ll�QC�	g�倃}��`$ ]��܏Q�^Lt�N��Z{����:��Yw1�2�N�vM6�=Q9���L9rV\� ;wݙ� �GS�m|T�F�8�.�>����l��h��BL>�wq8I&���h$�V���r��{q=�I;��λ&��\��Ox�*���T�Ss�Jk���� ����kr�4 x>g\��w��N@;��ςc�?i�=\��p�L�G�a]�d�c؀��{s1@z�)��%V��d��o/BR�29KHm2���G�1��>'��ne�F���g����û\�����|�6��Í\��mݤ�<���D�%�n�?-���/�{��� ������`	/公e�S	Pߤd��|�l2}T�/���{�+7 ��4e�n�Ot�.�V�fY�L�ٙ%-D�&,��}�צ��{�Ks�Ǐ99����!���5��}�g���'0�z���C�1Ϝ=��sn�]vM�oy.]�aCI2�Nk˲i�y$ =/[��3ռy���f�V� /,w���PUjz���o	l6a�
UL6��ff��x�6�m�� ��U� @|����!���6�f�O)�� s;[�2�Igw:&�0�5~��ت�Y�n������h��Ş{k5s�q�C��n�;�٘���/��n����Q�\��81 �L'kq�{m�a#:b�'g�sx��s��;n���O��`��NI��s�$�IQͪ�I( K;�ٙ�:��.�����붛� gg��)x���!��&\R-�um��dW�����[���q ��Κ�}��dߒ�U��y���XI�0o��@m��J^Щ$��Ϊ6^J�@���%54!�x�N�{5]m)׻�a����,����(fz�B�L�5�7����������2�U}3�3��2���n-��c� ��n�A%���vY�aCI2�N�FK� ������M��h ���� ��7���ur	���!�0p�`}�l6�a4d��wvq �n��g9c�
52c�\�I4[۝w`$A?]�ɘN+�����_@J�〄��t�<;�Fr��(�ޯ%�k;�9�?:���!e�^������AA�b2[���s4�9��N0"����ܞ�Wp��3yV���󸆐��٘�}g����*���gS �Q��Q�U:R�gjl�nof` #�}M���Ź�=�mwv�� q鈊��b.)�z�az����Dc��t+^��ͼw�;�٘ z���z=0L�g�S�Q@$)�$�A�̃q��&�}��Q�{����|ĺzk���wm㻷N��ڹͽ�k���H�I[�����[����bC�I���J֙�榝�$�H*AЎ̊�;w]
�.:v��]�b!��e�G�%ɏ z�w�س����|�y�� �w�&p���cN����Qv���ߏ龡jv��CgS�eݳٺ��g�\4�z+8�;�+�u���ku��??;�7D��9��f}�{][�  ��>t��ڝ��fF�w?���f =�t�@$���(01-�����
�^��W3~��f����@}���4 �fsv@�RC�n�UVn ��Q�'*&*J�)�+�7hn�@�=�*��"o}��#{]8�hz3�݄Wi3�!��e�T�s��ꝭ��8q��M���x�����ve���7��ӼI*_9	�<n$���x��.X8�����y���.��6��̷ �{ͫ @%��vf�P�jT/���\�W�,���-<w(@���_F#�o�?ݳ^nܫ�f�Ů�k3_��Ri��X�]u�rfWu]�\���Ū@EA�53P �����Q��9㷴�l2;p�t�n�i���[��|1��q�@�=���v7<�XMn��p���mq�[��g��ŷ���.MӜ<<��ժ.�z֣��Q�c6�c,�z���K�q��ϑf���Y7V�a���ke�����o����=�u���s籠�3p�g9N{bm����5�h���z��`�r�V݁��F��jK]M��kix�9�rv��]Ř�X���[jQ܋g�������[Yi��&u�y%��{�*PIy%���`e��g���$N�ɤ���)�iI@Q-�o?fg�ut�kjI�~���W�� Zg�餀���I���h�T��W:�d��6`�R�*TҊ���m��>{��0 ��[6��uxu"P\o2�QA$vw]�P|�"*��6�rh'���6t�F�Nf��L�ʗ� �fwUi%�:��{���	$�4��))�ba�b��w�����{V�f+s��{)o ��c� v��3���zo*�
S��GZh�8�|�$�Ku8�z��j�v;;��/oos8�p���߸��`TR�Ew��_�� ����  ]���"�UU2�^ͻ A��sxn�0�1$�0�חNS�Iy)d�|�-w��3��g�X#K�-���h���m���u+���e�jNB��d�������u��C_U%�
���\U�ͽ���{����j�>2��wZw��J;ن"�!4�-��z�.�h�sk\�I"[�7�òU�\N�����A�i���Jh�SJ*�F��c���F����<���^��q�G�;�ӏӴ�}�"�i��GBJ&�.�gй0L$�2��K�y�&��6����/D�N���π��ݛM�����vl��d˷��s>%�)e�
�X1��8�-���JȜ���ס"1\=��s�x�l������n�TUiȻ��ϰ �ڶ����S&6�S��c��j��M�5ٷv�(,��l�G� ��e�Ei��i؂v�Ol^^Wv>� ��^�~	�����I��<z�%��WN� �{M��RMLTIN;����@���$�B�:�}q�OL*Q�f��/�ګǫ@q�Ə\�]�-Q�Ny;ժ�+�T��/6�k�t�6�7zQ7��:|N��{�'�"�%���p�~��L$O�Goщ�o�&�ę����yj6Kx�<1�����'0��e[�e��C@,��̺����_��=�N�RQ�jA�CM`�$�:�^x$�����7�5�FFg�;wm�C@|ڲ��;w�"/�f�ߓ�����rváR�(�.{v�g��,Ø�x�{t�[m�g�b���v�~{��7~� �N~o���k���k�)$^����Vgy��1�n^9Ċ�Ii��f�v�DW��4�*S;�wh�3u�	�4^5y.I� de���w�0�dH�����ǐeTL������u�{��}��&uU��<\z�#����I&��&i _����ڼ<h$�"h���\�?@�sgk�x��_�@A�w�M �۽��$;���(���K��aU	�T偽=ݸ2��Nj�����`}�܋�����}�ɚ���j�U�ݽ�Pg6�)U�ki�4�K�n�P3i�C8{�7�4% ��I�L�`�|���8��I6ߞ�f��Yβ��E�S�� ����%.��TE�y��?-R�e�����s����;B!c���r�nyɄpk^^Q���?p�
����g�Xzj]$Nv�U��I�ft�$��ʪk����;Tɤ����d��f	���pbI��rI��v��9���ʻ� ۻٙ�DG{9�&���9m�Z��#0�Գ�1�^",6T:U�][�D��]��I�&��b�<�{��oS ���� �	��Oԁn̈́��8�&�֙��X/3;b1"z�z��I$�33�� ��ѽ�v.�'ɮ��w��f`w�pU%)��"h�����6�H ��wY넆�� >�����f�k����}T����P��֊�9�k;b�wU��^v�1������-U�ő�4�VA���K��|/���=XVs�-�)u:�g��}���I>���͊�,~��>�xa�(97��vk"��G|ske/�=�E��:���︯Kgfydc�'�^M���1��f� <��AU���4�]]!��x�;�Om8:f��~�MB��wɴo���?V��%u�w���'<޿>��YN+��5�nj��H5���ޅeD9�	����9�Df=H������ܽ�i�3r�Ƒ\E�j�$�U�I*�����a﹔�����پV0����|s�z����Xxk���:��3s�g�v -��s�?`xH�ln�&�n��nDrN��X�,�����!���5������6�QWg�"�J�u��e��Gñ�y��}B�!��A��b<����^����:���y����ꙣnŶ5�ro3�(�d���8�Js�~���$�>�w�|�a�)��78t�̓N�z��{g�ꄬ��n�xf�����E�[:�D׀2��	�}�^'���X���7	\��{s�D�P�o��ܝ���I����J���AY��E]�H��`����P�����L��Zպ8��ұ^xŎ��+������p�~=�3��z6֐x�C:N��鎓S�s�z�ʪ˩�G������Ԉ���'���'�E��-G>�F�|#����h;�m>�������F��OO��d]گ�zN����֓4:u�9����u���<E���AiR�6�EڅXQ!R��Z5+)X�(,�����#%eFڥ��EQb*T��)[--KiU�������*�a*"�Y*E*�b��+����*�TT"��b*�mTQ�ز�FP��edR��U$��%��Kj��F*
����խP*
Ki--k%��,�-iZ�**�����J+Z�J�[+X,�-lm�Z���lkJ�U���"�T��6�,QJ�����JV��K���%e[E
ԬQB���e-
�Qb�!R�(-E"��ZE��҂�[e�QBڲ�,[J *�bRKmk#iPk-`"��RciP�P���"�R����EY%FءXTa�q�Lc`���	x��z��&���Gu��g�:�����$��v�m���\cNE�����:wN�]�oE�6;\t]E�}�/!����uĎz��ۃx�=����֜c��������6�]��Rs��	]���N���+�9秧G[���ރg[Ep�������8qŮ��i�X�r�^xuϘ.Nz��v��1�lA��m��m�shϳ��Fq��4��6-���7S�t�^ܼ�k���þ74v3�6��#�˽q��۵�Y7y����ų=��X��V������=c�l�M�7C�t\�`�5��UwL�2�en]��50���t��β���.�������UG$�F!�E�']��E{v�.x���{���n	㫔܀��`66n�Nֹ튶�x|�w��`��p�[[u��cj�b�Z���c� �#.��{Y�p�=e��s9�:�v��n��u�Z)K�V��Ã�{qv��q��G;���k&z�vxvH�������8�v��$ݭ���sϵر�ֺ����wH����[��c���uɍm����jjn:3�t�n:����6�b�=Ѫ�l[F[�����[�(�r�v�n��p�$��^H8��m�v�����WX:/\Oύ#�n��\[�N���ۣ�n۶��Lv��v��m�E�"x�������ě��iU�
���&�';v�ƺ�v5���y[[m�[m��ˌ��[��+�`�s�0�����K��Ǖ����nyy�������璜���6�^���'mrGmū���٢rs�`��i�� ^66h�q�%�ٕ��:��)��m�F�;�y���ۤ�¼]��svn|/\�s��v�L��BF�n��^�������z����Z�{k������׋��d�lt���cI�����w<�k[����A�9�����q3�ؠ�7��˧tGC�FC���.0�]�9p��G	��q��:�붋�;���������n=�_`��m]��]<[��-<��`ŗyxY�ݎ��n��y{i�m�8�Fю#�.۞�(]�ـn�V=Ϙ�]�:���su�g�l�sV�-�vo6gy��X;h��{t'/;�و�9����<#�8'����=r�WQ#�^�&楤,�q�l�>�<�>� �<K�l�#@��l+ܻR]�<m6��g��q�����]s�f��z4�@��������@]j�B�vռE��lze��Ճ���i���vP�X�7���0ఊl����n��	�|�$���Igi�ꗱ�F����H${/\�B3��0��i��"������ɹ�{���""���0 23�Y��\�u��fZ�mg�G&P@ S,$��]�9?�&���� Y�g]aO>�?$���� ����Ei�#�R�UPM1���5G{�ϊ�`�	��[�""�ku�v�ve�<�v�B)�U�>�i�N6ba٥A*/��RJ	f�uX����O/�9����H##<����Ua#�a˾�v����h��/2��s���sK�X;����f,��escmT��?���*��%T"jd��z�鿀@Fkn��;{�3�
tL,��&�i�JM�S4��0�C�ʪ�U�Wwi%�9=j�fbS�D�_.f�
F����O��-9���奒���'�Jj��;�#_((���?�:i|(vN�ڻ�g�oY�@�� =�$��{�3Dof{�@��s����=�mD�Q4P��*[�n�v�sϰ��K�l���VƠ 23͵d��ݙ�%G����LL��fX�~�s烪�����@|��wv]��=7�]�4����3��:��n�6�$j"�E*�&��;vg�":��A~��г�v��q��f�:�`f�vf �^m7����G�W=Q��d�^��!��Uͼl��:��sv�Ld10��m��Sf;��و	�Kf�2c}�;�{����� ^m��'����]]_�N��n�o�������S4��8����s�$�����3�|*RD�gv��$��z�Ey+�Sq3t_e�v����p�E6T���I �fհ>@z#�^(sj�����S>�Y=�w�\�>��U.�އFA��Y��s��qۡ�5��wg��y�����I�s=8O��׮�����<]��Ի}��7ݽU~H�����8ԃ	�	�a8��Zv�F��1�m�[�"7u�Ł� ufۆ�͂b�[vi85䗮{2��B�p�PK%-P�|��'	���x�\��w�2�����ّ�H�Φ�@�3��q��eK�^�I�t�>!D|EFS>;s���k;�'͌rZ�jwc�[v���x�nb�A-0�l����̮�J�]7�k� I]��	?al��q��"c��;�ٙ� ���ͦ��6}3>���W¥NFsN�O�7E֑���<�`+��h�I�=4�A,Ұeē�nDf�$�k�f1	�8�꼻f�W����/nZ7<�g���@|sΦ��Fa|���袨�U4B
�/o�!c�K���]� �ޫ�a{&����ُz\��n9mɎ�;�S=�<f���g7��� ��Y\�6�����;P~��V[��K�x�y���2�)���g�	��b!���w��ʷ�����D�B�QR�n�ۣ�v�s�]U7ލ�ȍ[Y���kn�}���"c�Z���*��C(���0xM*����u��A[Cuc�!�t�Ϗcgٔ��2�#xgs�A&(����@�ki�����Ȋ^]��o"
AK�uA"I�]SA�J���L6StOWWV�ZA'�fI�z�i��si$��]�Av�vf|��3�m��6����.g��J�E����	����B������ �Y���>�l0��n�>@n�vf{[$�SSB&�Jl�O�sHN��YW� ��:��wwf` #�6�[������ÖI;i��j�֓i��R��
��3 <�j�K��U�glueu�{f >��nZ ���π��O7%�u������Gf|�tݻ��2���[��J��d3��Y<�o�yH�F��W=q�>�5��LNˣW���ZI��B������Nu��i0���d�*.�upq��`9:��V�v�ܚ8�W[�`��u��H��+�<W^M�X-�l��V)ٞ�/1n�ڣ��g-̆r�㛶�;�t�c�	��Y[v��q�.�6�H141/�����>��E��݀D�<Enݶ�.�˦h�u!��s�*�-Ş/n\;y5��m�/k/���x�loW%�����q��4���[\g�ٞ�Ӡ@��Ge583>�ٜ\bZ�A�Y�񓸁K�0�=n~߶�������7�Ɠ� ��� |���a�{8�3�׊�owvf ���bd�)�PE'O�ߧ�4\'Nv�Y	��f��B	������s��"��S3���=�oѴt˘��QJiN�v8��=nA$�9��{��D��3��ɰ�����Nwy�Q�E< 6!�L�_,�D�dynl�C�v<���W1�-�uOC�k��}����	+���tl,�iUIQ3Q%[H���> 6�u���s���z7�}���F��mIF��MB��"�s+��;#bBl���B�1Mɗ��狚���wSr�����9�#G;Tw��QU5J��4�����@�k�I�Iz��ѯ$�r�7+��ٙ�|y��h=��%L)�����y�;�}�\s�ŧ_�QyTn��]�䕮�3x>���h/�=��@�m�k��)���Ss���'�_N-�s��7�<�A�i^�����I"��[��@Y��A�W!w��7����đ�<E��K�C����!""=]�l A[U���y=���|��� �%o��4�ȋ�ZP!�a6ᣳ���E�{>��wS��"v���	%�rh�H���]��oc�LL��u�8�V�r}��J*�Ql�&}]6 �{���y޸7x+�L�Z��"���6 {{�"2b2�ܧQ�|\q�o��j�n��k0qYm�����w`���񮋺�\ǣ'am}��w�Y�^�*�=N�� ��S�� ���Ȅ�	?;/;�	���mp
T^	�m�Ȁ���
vz�<4����+'�� Af߭���{�1Aj��D�y�zcm�����J�h��h
�[A�η ���0>A?}3�5��˪螫��ۭ���Z�p"���ڬ4m���y�������A4��q$$E�ɞp�)��`���t�D�-�VOȀ>���;�'�	ˆ�h�Lb�v�U�j2bw��E�>nq�'� ����0�=�6�������> ��T
5��Ɉ��4��Tᣳ���}���Ԧ�S 0/�똇�f�uݤ�G+q�x%�q�C���F��e��I�q�!4������.�vr�Ⱬx���N:�*T�
~�$��M"M9�[u�{�`  ^{�p��ǵh̓lxڢ���$O�>&�J�*&UIt{j\�^	o��ﯛ�m�$�U���0��mDh[�{6&x0�����x����*�Dқe��c�@ �ͫi@�|z	��O���Ur� �w�3��ͫh	�Pڊ!L�
"���h�=��D�X��D�fu_�>�6�4�_��طaN���2�4̴C�[q�R�de�f�J�>��w��0�ʝ��[��۽t�g�qTc7���h�p>��3\��{3T��ɗ�9�ٹ�
〸�
���\;/�I��6���C��}���<�l �gm�:}�*����o˻z.�ڻx��a��X��Ob+�;^Gk�)�������_��n�+�q��v8���V��:|ܰݺ��O{���.$y}�� �:����&(	�RIC>/�:|�\��~�S�{���@.y��� q��˧v{��{�~@}{N6&�J�L������q �<�Z�*J���O�ٝ�oP nf�a�<�M�u�i�8ECT��]�(Th���� c�[@ �3������fz���fr0ޝ� ��M��T7Q
I�PJ*[e�t�wws�'�쬑�z�S{�p� 7���DC]�ݙ��Q�X�Z�! �,�����nV��t��P�,u�n��bJP񝑧 ߺ�[�P���m��ӗ�kK\�Q�}s��(�Jc��C�D6,������5��퀲d�۬;�����m�C�����fd����s;c�%�ڰ��R�ys�[����n��utuy�f�����u�w]��m��Xݶ6��)��Z�	���iz�;gA�������}v;��j#�s����]����=q��G�����ۏ��0kx�g�Q^OW%�mЗn���t�^�����N�4j�Ċ
*n��1��]�6��N�����k۬�o���:�IPT��_���� ������٘�a�I.}S��w7�h�drpߵXD��j\�`�O�܆��gf}��c$Q�D�qs�]_�  �\�Ȇ���|P�as,��z"�b	�**fh�A勵�� ,����PKY��XM8����8���#:��D?�����+�q�53SMak
C����1=�6�Y$�w������wfb��gS�~��ȿl7�a'���Y1�hW)6XJx�~�����:�#s'�3֤˧(��60 �w{�1D{3��Z�us�	����������nzy�]� �1�ӜA-[�±�2�:��8���������v\S|�<�r|��x�>�>�g[���D@��q֎ˋ�I;�ݷw���t��5���1���\'v�������W������)�{k��o�<{n퐬�W�[5������p��|z#�݌I9NE�"����ػ�eT��أl�BȌ�;ji��s�������� ��|�$������e�ߧU��{z��p����C��{/�Ť�K����'���d8��F`�qҹ$C;���$I��sI/U�* ,%4KME��t�boS����7���x�	��&�y"PW�E�n-[/,�J��'fw�s��M�k
C��9D��Q�*X����$�]u�w���I�{��H$�=�VDx��u��7������.���[���- P&䙪��kn-m��g����P�X�3{��e��d�a�*����� {3�� ��^c@���>������<�6���L��#L`H��}5zDp��xh��}��^�� ��ۆ� FWO�� {5�k0�����JO���!��)t�fӈ` ���1$�2��=]��Fvn>[���k8�V2a����:
cFej�~SQW9���:w:�^�N;�f��Gq��=g,ޱ���[��[��IZ�x���X���5�{��D���,���R�v��VzJ�W�r�g�>��9�[�&=�ӫ��V{�y��Y���.�3�t�{�p%O�=���ի���ڮ��ԅ��~�D)`��ٯ
�%�z~S�GF�	�ӟ��5t+�-c��u���g�v���\�NY��f�/�n��W�;�^۱���Px`Ӽ��������x�ؒ���"�F���w�F���*u1�	��tt��)�8TE:�^�f�m�i;=*��q��|��k�U�7�!��>޺�!@�ɘ����zf�^�|O_2�%k�/t����ͯV�!}��d��k�D�7q��\��y�7K��J��~~��>��9������5���4�qn�������"2K�<�c�,�� g�ɽٛ�L(��%}��� !���h7�#�j���j�I�Ѿ�F�N���)��F������8K�.Ʒ���%��91�zh��9';2+��eK�����V�c��÷=���%��r;�]o����{���{�����,C\�Ƕ�WH��o.����0Ӓ=������(.gB>o�]/�'��f��,��V	7zK��O����;<��h�[j�8b4n]<�V���B������g��=x�/@��r�~�<~�mv����|�v�Q��++�_i�Ǖ^�����;n�>$x�G��
"ʄ��T���R�-B6�FV���VE�T����ijTm�
�Z�B�V#m�UQ����T�(�A`�U����j�TZ�YV�Ab�iZԢڵTclkb�mX�*�XQ�ZF�)iUR��VX�##��VT-�+X(6ʬUREX(��cF��JV�T��F�V%*�,Z�-����Ab5�b"
���%�P��H6�-��������cX�mU�ڍJԭ"�����Z�څ�Z��(Ԩ��B�KDdX��[h����`������j��[V4�*)(��V�kb�R��kD-��J#im(*IZ1QQK�,�V[m�-
�b*�X�J6�*6��P��A�AX�m������#ZS���7�"#^m[�>FQ�mPF�zp��,6:4����̓����4�M�	J�8ܨ��(nouۻ���Û�q���mΘ&Q肈���,axki:#۽�0Y5�1p�('���Gy�C@-��fb�#�$I���~<�]s�v����r�]t��`7Z���6�L�y1K�i��s�����1�t��`�G�yM�F�����osx�f�ߪ^����[�N�4Ak]�M,������)* �T��f8ς�y�1�:9��������S�9���ok| e<��<�\�? >���j��_D�-�P��B ;{���� ����n�绮/3#R #�{�舃��٘�__�ȫ,E5�G0�~r�WE���ܤ���cN� ;��3  �Χ����0��t߃j�.o�����ZF{`9;T���EJ��7�l�'n!��
֮�t)zt��)DÜ��3ǔx�\y ����@��=8��L�*��ѯ-����^K���8�n�8�>e�t� govf ��lė{���c4y�QOOO��,���\q��&ډ���sV@k8�����!t������߼�N+��Rs��W�';{�Ť%e�M	uMel��Ѷ ����J$�;7�3>@$�/�b�JEDT��չM��<Z�v�踿u�� >��vf �}M��"���}��(�;=}g�gD��2T0悭�˻K�$��� ��ʌqڽ��S@|��n# 7Sh'�b-TB
����m���Y���q�����`@�c�q�rJ>[��z���� ���;1Մ�4��SXs��&a$�(}��J�U���	 '����^	��5�D@����L��]SD��qw0+}-��C��y����]�/�.7�޵&�f��]��R�ջ�q*�>ѹ9�~�����/���(Q1i�! �.(�+Hv��=�����\7AμW���/l=�����:3�����m�d��<s���t@'g�Cn`�����ם�otgur:�^Ln��zi��ɷ-�ۖ���{U�w&����cn9�Nݸ��cpd;v�A�\�^���g�<��ɻ�v-�/���ٍ#��6<or]�n,k�u=�g����n�g���9n۶6��r�7d��h�y���ֱ�{Y�|���K�<[<g�?>�:��L�*�S[1���� ���[  #+9�	w��(��޷ّ�H-��D��(PH����$&�Xl*���{=�=�z��=��� Vs���[3�����O>����|a�	��I�P\��A"F�ْIP�T���=�Y���"?f�h @)�i�ٔ��j�!��M����!���u�d�P �z��DAO]� [��w�>�����G*�� ��`��UT)���qo_�l����au�;�И�#�	���h >���C@.��%vT���M�r����h6	m��]�u���F�J3�j�i�@"�e1�'t�s������1�ED�&�D�r6�i�� ��lA-���ς�K��s�-�7-\�>�ra s�Y?BG�>]�)2���P����3���H���BS[޻)Y����·��}X�RP�|�u�ճ��)�zt�+�h�L�
�Y.+ZH��M�J׷����Z�6�fﶯ�  m=v� �����T\b��.�j��}ԉ�1���EMH��
��� ���sϰ A�zB���F�M놀i�i�$�w��".�]
JB�R/~'�)�S�G��z�@�ci���ݙ������\�_Y9�H/��ʇ廊��B�4�������  ������P�ڂ�Rd�^�^�;�|����π@!�u7�r�^����! >�q&D2[(`x�=r�pu��<jWz��<��S))�A��L2 �wÇ̲Bm�37�x�g����0�=Ϋ���mսf$,��� �{{�1 �VH�1����(��w�pONg��3J��)!Vf�J�ow]�M�V�:$�%��f^�
6�W>줁�WE�(mTҪ�-��D`vgU�#OgO������ak�ӗD� �M����ݒ�C|0R�B\�gH�=j{��ӆ�vU��H�fɟ}�MW�M|7��i�6��q������&�{��$��u6�R��1�������@�/��uF��� ���cq�fu\D0"�����i��ѧBJ�kn�$N�E
jB)��չN!�>��;MLR�Q��݈�_������m#/��%��c��ǌشL���s���V[ �y,L7Ra�u�9�c�c�n�nn^�i@1/������"^$����H>$�ٝW��t������'���3Y�@ ��<��Iϟ��0����i)	��t����-O�9�����^ ~��p� #/�� o���$�U��� ���\��a���W�$�I��릀A�T�������I�o1@n>� ,���a��D�&���U.Z;/�;-D��tG�7�{��l 
+'jI����۱�=$�f]�
�e8��"�#mߌF{�{�5�$��-�y�\�oOI\����ȫ���=����9ŸDtE�Z{�/({Ω*�����p�L��T�I�{��Ӝݘ��^6;+����4�	��2-���ѐj�����a�8I�Q�\�ꈡõ���;vLtvm�g]mt;�Ű1~~~�~�P��"�RR��չM���۶�v�nf�n��y��y��D@�����,u�MJ��B��*q{�߾�A�{U<�Y2s��Ā�"{z�%��Ih�Vfvc�̼ui!ϓN�W�UB�����{�͈ ��ט��e�Iۼ���Byz�d!!�ݷv��)���SM�X�t���t��+^�� ��?� }���� ���n:�fo"�s�DC�vcm��(!6�l�۞ۻD��|�[9�馝�;���w3�I$�7���D��o�W�D�v4��	v��i���q-o�p�?.���{��xz��c"�^W[�3"�.9����G��ৰ�Vz�Yr2��L9(�B��@���!44�I�Y��(1Xx�@�%��!�����5k-h�;Jpt'�wg�:N�yoj)+��:�0qt��q�vy�������9��sOPَ ܼ۠:���a��絮x7)�z��1��<���sr9�۶Ml�Γ`D�.�m�g�Oa���X��cf�s���9�-\�z��M퍪�:nt`8ݵj�6����uC/��7::䵠�������H��f�]���p�ZD�>|iֹ�\z��\���}���6�T�*���7�m� �wkq� ;[��:�"�}�wB3�.��� ���ۙ�7�e
b�
EIJ[��ܦ�A������ʩ����b >����OT�H��kꋳ��Ë��WPo=ML(a�*$��<�R^H@�v�Dx��Wz��z�@}ݽ�� ��uA$9�L���""DQ#6�!�_mys����X<߱�X �j�$JU�V˷;�f��Q%z+o�ɌA�y	e����K���	8NK�H������@�������D0HU�T��ʓ�S�nQŨ&�L�<n�rlݷN�"��B-��� ݣ�b�3����1hPBm�m7��6��Ix%�����@(y|킆���^����{�������f̒�ʚ�UC�
o9�����J���u5盐�̔z�L�e蒝W_r�1�VU�z�0��
I��J��:%���S�|���ܥ����:|*�~Gw���Gc�` >���"#cz:�n��u]�����@L���o�:�)�4����S�t��̪e����Ǳ�7�@���i���a�!���"�*ޫ��ٓz�ѹ^��;�V�/���@}����Z�qӉ�~ �ͦ�K�xC�U�UP�f�e�ۘ�M����I���q�@:�[�@!=�6���w~H�c�g"�dNN��E�f�6	���x�9^LQ�q��x���qv5����v�~���&����E�����@	���� Kw{s"-%+���[y��w7a B����}�E�&f%L�sh�6�|���Y�9����uy����;hK�/n�mݤI��ÊVm���=Ͷ�%�$�/���P�[�Ip�}��>ׯיܣ6.)o=���/z��e��y�j������'v�+w-���ҽ�v��	��f����c�x8��w�w���2A&� a�۵$�I{s{n�$��m6��L'	��ul��7Wut>�c� ��M���K���vI6��:�uQ�����A��I�t�cA�%�5EPT���� Y��!�i�6ѧ�+.�fGt�k@ ���g��z�RS���[{������{��^��<�nnx��E�^��l�\���ar���3������o�u�13U3|�1��ݯ0> ;2z���s�Y����5��
D�������<��P�eb|��H|��>.&6���!fn]� >���3D�����$��磫o�ٿv�g�U�~���UUZ9����;2z��I,v�LD��N77$�Hvwmݤ�=w5	W�D$m���j������]��R�7�1������4�<ߥ�v�~��6�*���eh_K��v�zq������5^i��͏*Z��,�!iӖ�rz��P����r�c�@
�d��g�g�x��y�]T"RB�v�Tt�Qr�_d�$ק��3> #s'm� �'�Ͳ��;�DH�!�$4�C�i7�b��ֺ,����L���p��.�Q���￴�mZ���{{��  �d��  �_;hLY~�/�v�D`F�O[��!���m�m)?�{�a&��_�=��X��y�Ā�+X�'Y��dԌ����5�J��%�f",CH6�j���d�r N��6A�#K��.�S��}� #�'�R@�u��6�4� M6X�ژ��շF�	��(�'�-H ������fw��ڸ��x�O_/�D�~$G4�~�b���]�4��<�����}��@){\��D	�k&@��o����f':��܅��S'v�rwap�����gaĵoޞ>9�^j甌OO�h�N)�o.�u�.0��74�:ZLÞߣ�����8��ygc������t�dKLJ���|�x����sl��=�H�>�u������s����=M��=�eCh��|��{-cxd�;,�}:=�'g��3�~��קh��,��{��ǯ�ࡈw�����瞠�������k\��g��y��fx�{d~�ީ���O�Np?Ӛӻ�㩃Do=�[K^�r�����Yө�z	�G�K6M,Kƛ7Q��'��}�ޙ|ؘ��BXtvR�^4�篽u?s2N��<��k!ِr$���S݂g�1�8y�x�G��ꢗ�g��[=��J�Y�QΤ�_�A���v)}s|��yڴm�ؠ�0��W�.ٗk���-F��ڴ�[��s��ܨ� ��?AFg�E����k�����@}�����!�~XK_M��kꠝ����a5�%�_ ��Vp/B�&��>ZKxB�'�����P�'��F斈��Z�p��#��]Y��uY����eg�u�o����p,�ذv�07U��n���X-�'+'#�����s����/��Y f�F�ڣ��S��'��<�S�vRW�f[�BS�\i�wDG2p�|���R-�nN��ҏ��T���^���dSݼ�4�LE���Q:g:��9O{cy+�\l˝dw�F��j�}NZ	�
��s��0VG��M���sn
8P�V*�m���#U(��e�E��Q����d�E"�QJ2��QU"�-KEkb�-A��4Z[F��Qkڨ"T���Z�!iAPjUE��XԵ)Qm�UTVc-�ʋ�b�YR��$b�iQ�V*b�-A��E[eVZV�YYUF�E�eA-�eնҨ�*QV�eeE�%��*V�J�J4+%JUmb�1��m�"�l�T���ZPX�J�%J�KJՊQV�Em�iEUQԱZ�[b�QQEQ+F�TV�*�UUj�ұ(�Q��0X�
*��E�U�+)Z5�EPA*X�E�����+iEAEUE-��+mh��UJ[V(����YDTAkFEE��������J6�b�2�V
%T��pc�1���|�ں�Gu�C��v˂#���'����.�7뮡u��t/v�����!k�f���퍳b�q�yT�x#�9.+v�拞�XX�S��c��'X]���7��;zϖ�J���m�ͷ�ݚ�v���]šx��u�}'k��W�ܽ�cͣ$FgO�Y���g6!�%5�}���`Þ{	�:Gv۫���͗��y9� ������,8�۷B���͜�unR;��ۻϵFwX1ۍǣ�� Om�x����ŊNB���t+v�a�m��՝uDI�]l��a��S���nm�늩�Ҧ�7]]�s�����;�N8<v�����g5�s�]��ڗ�5�����Z��;����٫;3.�qt���qsU6�O5���v��q5�v��:�^٣v;n�	v�&��;u�^N8�k���ص�^Y���q���Ŕ�/r�0m���]='H�D;Y�.+x�&���뭺'��3�`���m�}\j/9�������lM݀��:l�/b�٨�g9 Ē�k�-�gxI���u7<V�2q�&�`��I�W�`�l�Z�&���lGVsŗ�]��ݮ�JϢ�#����.I�x�#<h9"��y�<��Dmĝ��6�m�޵ȼ��v#��_s�rN�Ȕ�)�	������b�Fuu"�6G���l[I�lOad�˳y4q=t�m٥b[v�l�!��k���m����x���䛔��u�]����0Y����ny-�y�m������Z�Lh�vT���3��9�ưk�/j۰�.�����m������m���� ŎW�"��8p�I�����-��v����&�{aϔ�]�-k�qIC�+/K���<��\u֞w#�q����`�d���ݸH\���;�A[u%��VwV�c\z��s�md������
��Ƈw9�㕣m���N��'��ܬ7DKݮ˞�l�6��v�a�F{��zE��p/;X�tG	��Nc�`Z�<�`K��˛�x\o5��^7q�Xwx��g���5�j8wn�b���@�F7��i(��l�y���n��=v�9ڵ�x�67pq�ve�+����ݷL(!��x�n�Y�ku��t����=d�����8<mqqqv��n��r�kS<t�&�U��rиm���ù3f��4�g;l�ښ�.tm�7���w^�x�zn)��aŚ�]��Ay������n�9n]����cx觃E�u׳��NZ:�2C���g��ϿmbQDR�b���N7!� �v��> ۽����}qf���F�O9m� @!:�o�e���ʁEUEM!�����I7F���Q�{x��[�L$i�T�^I۽�d�K��p�e�J�n.w�N{��a�-��M� ˿K!�N���0�N�-�Gw{�G�u�ڤI]��vM��b"0AhC0Z��+��O:]��g1r���> S��M� >���f �ٓ���lnx�o��",N�m0ʉ<b�UE)��r�F����H�=d*���d��{ϝ��w�����;2z�"rgs+b:M�M��pJ��K�����a��ɚu�S�M���ٿ�,�-u�RI4�~�j��V}b��oy�� �2��(<\Vy�L��,�Ͳ{�٘��]EA(�)I1J[H�����AW�Z��9qNx��}y���Su�s��h�z��vs��$��p�*�{B*-�@�"�8O�xO��z������dj"�nb*��gD`�w3� ���v]�@������� ɻ�{�vo�-g���Z۟�QSELT�7/�3 y�:j	�Ï{��1��N����^`�~�d>�j�~���&j�[@��3�_tgC��]x�w�y���+�0�����ڽ��m�g���7�^�)�U%L�&(�9�<�R �"�t��L��Z��^��K�����$'Yͦ]l�{��]�ɽ{���0 �	�B$1� �+����k:��is��br�u�F���x���~{Ek��+f+<�� ����� 'Y�m(��w3�t���f`s��iHFg�IP�x��1O������h��%��f(�}��x� �_�X� HN���IE��;8"*7�s�Kכt�)����M*l�m�|�u�� Z�<����X�K@If�S�/�7�V�cA)JSo��p~[g���H��sO���1��-e4fz���;�o�=�,y���׬�?d^l�������@|y�� �r>�L������ ��M6��teǰ��e�50${��� �{�� ��ft�~}��\�� ܤ��=��ac	�CI�&���ؐ���Ņǻ/�iy{�״oW1��>��� ��7�/��E���Z��&v��]�M��b�K�3�K�3rh�t��xx��=e9?�����j��P<�x���� 	׵� �Y����D,�5=22�_�y�7$	�m�͠2,M�!�����Tzv�U8���}S�����:�;i ������Kn�{"I��w���TF��UU/�S�Zn ��7�O3U_F���A	׽m�����@g�͖S	��:��f*����nLa#
s�� ����� ����]��[���S��I��Ad\ܧ6 
���F��fF�>�}z{����Rj�*��~�x�<�ϐ���{�+����/"9����cY�) �R���m��b����z����!��ݰ Y�ۙ� ��O7��V�}�����L��rl�:m�Z*��1�"mc�8Ya�3���%����긺����~o���zJΖ[���퀃۽�0 ]~�dB������.r��cl�wv�`u��E*�UPJ�,�����{�w�W��{Sg�|v��g�/�G^O6��I����w��П4Sa�l71�}�V����� H�}�w���~�����fb �'��fh
TO��gT'�Ӟ�7S�����n""3��p� !<��K��wԵm@��}���?o�E*�4���� 7��$<�'r����es�����o��'�ͦf^��N��D^p��b��,���	6e̕:��)��܍��D��R*8�t��G$b��L�f:�.�Yѳj�[��:��܋4_otǉ�VO����)n2�	�:�DPu�^)(j۰g��˴�r].��IE���ҎL�r֪זr#vsc�t�3ћ8���b�vC�p��q�W�ϝ�G�H���6�h곯�ϕ��u�9`y-��u�FC����2����I��e��Q."淇TҜm�9�pѹ�w"�cy4���U�)�w.��	�ظ�:�<�:n��tl�6�k�Q��\�kv���\�[/m�h�M��Mm�p��ǰ�ٝr�Cp�Ȗ{8�pA�
!�0�����։Ic�rI4^5s�4R�����qt��3�31 ՛N!��j�3L �iHN_N�fN[w����{��y`  [Y��@��_6�'��Fg|{��뒃�c���b����h �O�Ͱ�6t��1��� ��u\D4�_[L4�zZ�(M�!��)OVu�|�ɍ[}���A-��$�A$k'*I����:�<
#{���Avv:����TF!�����
o9�� ��sϰ��{�s��_|���q�@!=�6�7���J��Vq�w�sD�i�5v�G7g5���Ƅ�x�[��F<���������]8����U��r�W׭6 ;�٘��x5�[�=��׮�������y�t�*�biB�iC��m�� ���-�]�� �v���<��*�sڹ�w�WI'=E��y����qen6�ed�&�#{nL���8Q�2�ƿm_ ^ߝ� ��vdDC��y���vѥA2�Cf��(�}U�K�$��:��`%ow7��;9�7{�x ���L�3{����\�D�TЦ��%��w�N�t��l�&? ����D����@ >'���gp���;���!M���,)-UE)�]E;Y�b�H���4[,��l1�`��X	Ff�o�fﹼ O{���t#Y������4@"�T&���ZA�q��[���\�oZ����������f��5����
�W����i/$�vtѠ�^���&5�9�9H��w:����u�PR�)H����n�@��&)���|؂ ��vf�^�l ����n3x�nkI��6m
��4�IUmٙ���#��h �e��r���!:�
P{�[Ƨi�V�j��\���Y�g��>}؜@g,�1H���]�oI*VH���n��g���ʈ�I�y��dߒK�s�	!�F�D4i4�'.��n3����ߖ���@��9�����3�{�v�OJ�*��BԦ���Q*U�D$��߷}�k� ��{7� %6�fb �W�Y��N����o������~�|߇4q�Du�sp۝-��Jsy��M��p���,�c'9��}���`�7]UEl�V{ϰ�����> y|��m�����O�;���f`uzy����J������S}���_�}{�y��\OMg����W1��s�� ��(�\O�y��ȇ�z�IJ��"���;�-����π�K���;yov1���$�<�:kЊ�I
쪠)d�ؔK�"d�-뻾q�9oEE�E$�r�h >��ݴ�@f�vg�Q�:h��+gdb�?Y��v{��H���q�N�&׿'o���g�u�&�\f���d��KKy�U+^��w�pt�!͝���2V�_$r�;g�N_���D4i4��rϺHp�A�vsŃ��~�Yֺndfg���cD	�6�ogfb	��x�mD�7|�:Q.��Og�TN�҃����Lm�^=�k��`w�� :�~^,x�M2���9zD	 	 A����-��^���J�(�U�؈?�/�̇7�X� ��5UE\��ً���Y�\���#����n�D���� �g�ȕ����e^���#IO��gL'>s�lݜ�DD7�ި�u���a� f�q��٘�V�1J��Gf��0�)����:I�soc���3�9�@$�����V�I`�M���U�K�4W
E2�`�M�TwffbX �Ӷ��.$��F=�l"���Ȍ^�mH���8�f	�o���p��p�Kq6�q^�Y��Vn+�?��o����b�m�m�F�e^�䰣�O����� �qz�(�o�{�$�ra�y&Y����!|@�Cۘ�+p����z�6yL��au��nՌ���yƞdm�Y��O;�I�����۴[n
���ܛ���u4���:�V8���dG��9�͗�+V��u=r�<��l'WRH�mF�Jmk�k���j���msX���9׎A�9Y뎫b$��c�׭� ���9Z�ԯ4����\�ۮ37���wd�Ԥ��T�{q�ۮ����"�����m)�7lv^*x.��:ſ�~�֔� ���$'��z�$����K����T������F�н˦� �nvdF)8r�B�D�L˨/ӷ��P��z=?�]Ԫ��l@ ;ݝ���:�;mI������,�޿R��2�P��i�R���a$�<����A+�l�ԍ�i�^F쓾$篧��q'ίH��.�)<xeK)�a����1q �x� ���h���V���ӊcb"]�y���/h��AS*���޹m� �?^��ۧ~5��&f����^�o� 	�������Ts���o��g�u�H��\k�\��..���y����ذ�P�0mUd� ��<�.����p�"� ����Ә��綹�3> ��O7�oCt0�(��l��؂U];��j�L�O\[O'w�nU���mrO�
[0��LN������ě��{�r��|��b��`̒3���K�GroC�5���Հ kլ` '��� ��'��J�v�/��/B�PW�F!��"��T�� �''ޒ `��|��d�>�[:+ě���$mvUQ �-c���0�MK}}Z��D�H0�6|��y���3��N��ޯL��uӖfZ�1�&&q!-��D�WM a�E%5d�Ezs��".��$��Wټ�����ǭD��wf�ܭ��"j6���t�j���g��I؃�MƸ��6�z�,�&�J�ĳ�!8�6c��q3�	�Ϊ�$}��@��f�
����/����z��^��D�RUCz�q�i�!NP�QM�<�5]�T	$_uuQ��3&��p����"7L�Q�N
-CCE�ݹ�O�` `�zggS ���܍�G�5-?U�r�������y�˽o~���uղ�Nټ'���|��߽��k�:���zA)8t��x���k�)}h���%�9a�J|޳P��5����&?0<��T{{-�&���c��:�����"�<'�^T^��d(�2�r�g<�.�>���C��#ûuUP��\�=���=L�4�(�����3o����F/��k)�C�Ҧ�}��{���x��]1Ƈt��Y�`�2�~��ͻj��_d�j�z)脫�V�3�o�� �?1�R� ����=%����z����Fއݾ����f����^j2L�o�: �dg�|1gy��G5��~�]W��.� Ҽ͍�Jw��x�����4�>�y���$L�j��[��֬7�/9H\>ۻ���T��{w��v���_.Z)�j�w�:+���6f�����d6��n��8�gnB1d
�鲸}��e^�>]���ν==|�~NY��%������{�$��kP�^5�^>�*:��Ĭ���$\Z�vE]d���}k�����7���$�\��9^�[�w��48�<�`��o�Y{ny2(�"���M=wKU�r��:e��yp+�vQ�=8���;hW4��'�d�ѫ1Hp�#�y͝�I�"vvT-��o^�M�,�寗�w`��̹�y����a-:!�h��}��U����M��[���%z�86��|�'%�9�p��bݞ֐k�i5�. �=��Ts-�gN�>پ�g�a�3����1UM61Am��iAZ�DZ�F*�F"�([m(�VUUEb��Z��D�U�mj��c-�TV(�(�ke�De�X,cm1�F�b"(�YY*
�**�DTb*���ш�-�l��������l���m�ʪ�4��E��X��ڋ
��A�kD��Z�m���4h��(�iF%���Q�Ҫ����6�"��ֶ�cX��X�KR�hQERж�AF
+Yb�*�����%�kH��Eeh� �"����-acj
�UV,����)XTPb�DDTTD������"���jDDV#ZQ*��[amX*�,%�b�Z�"���UcE���
	����ڢ
� �F1-�UEV*�jF"�iU�ke�h�V��E`��b����� ��[ϯ5]�U�I���O��U�!�Se���VF�.n�D�7]s�M�˚��wo��	���-���`����&0���J0�n�7��D��q���퉢�������;��N��J����e\tmب�@����A��A%��]�zی�<��ܙ����;um3cv5rG���o�~��-��1�U����xdӊS[C�� �5�L�_���?KAt�4�E��A�q&Ov�ʺ9b0�m�	$��q�H#b�(��L������M-L$ G�0��]� I �\l�Iy�YX$n(���F�_Ux�Hb�'��W�u��D�e44}}�¯2��5 sۓ^$�MŽ3�|OU�V��f"����F�L�b�te�29� �d�)�;�/q��MS7%ĺ�����ȳ�f�������S�{J�Ç#]o_)����~^z���	�P�~��I��1�F�))�j��0e�O�s\:�U2A>�Ϊ�������}U@��������FH!�-<8�_�<�ޱ�qr+�kʾ4��H9����<<��w��!�`�n�������q����T9um�O�^s�!��~jK'�U�ۄd��U)�[������f�CE�}lȢN�ƙ$:�*�ӽn��މ��=�j�&�I0���5�� �_I0�z��t����W{�@��qq��F�eL��B�D1<s�oM,Ȉ�}����]lt�I��r�����_l9ڻqh;Z�G�~����$4��z��A �ۚ�a`��\�����FA;�����A"��ꁘ�������^C�Gs�(R��a�J%�$����u�B�^���ڜp�כy}��w�o�|�[�hGg>�D�ݾ�w;�?>|Ey��y�˞�5�u�sX���Y�T8�2uu�6�vp�yy�9��#o"b�ѹ�P�m>���18x(-������NM�<�\� 6��.��%U���1O��5v� ���zCv��f�[v� ���)�jk/t{u��U໑JӸ�p��e.�q��u��X�8�i�J�v���S�14s��Z��t���a�܇T�	n5٦v����m�
/9�2a�b��q{S�7	���x�n��9?����߮�n����Ull�@$ݗ$�[�r�A��Wr��,��"�x����O��ոH�P�1K�ܪ�(.Sp%�1�	$wd̂A"���I{.�s^H�\��8���addCM61���H�	;��"�%U�ޞګ�<A��A �+�j����hq)��E2���kq��V2�� I�}>�	'wv��$��1v�����k3��E;�p�b$D0��ՕD����d-�&�w��4�	��� ���U@�;���ή����C�(�ӓT�N�ͧrp�n'�vg���~l%��0��9|�@���M�񩝙 �os�kĀO��;xF�᧶�Dn�a�砒v�j��#ẍ́�
0�N"����Cxfu�v;�8�]��ϥ��}v�����ս"͏�Ɖ]�9V�͙�u�N��d��P�)�PΆ�&����O��v��$���%sb:`ڝ�}ُ�=3ݸO�i��*f�#d�>#��ς�w���w��<H$wn�P'Ğw(�p7(p�"U���]H�pt���<O���Dv���;��VĄ߻&�c�ù~�K�hq)��E��Ϫ[ل`�͐&;R��ث$E�m
$��;�'�T�z7�]Z��p�4d�x7���+�W�<cnm�r�+�栋��v��}��� �	aջ��ă��"O�c�^�v�/�~x�~O70 3PצV�4X��l���ٍ�b5Gl�$���$���$�\�nY9T����^���A�[�5�Udq�<r;fH�����yh���E:p��h��ԯn<�S�#cB�]�p��;�\;���d3^�k��D�>R%G5.���)�ʷU�]�H@�z;&A �*�8JM��4����)61����f�0 ��$q�3�I���UvY���;b�biC�P1���O��H;��5����!�}�H�/L�	�� �}[�T����8�6-BN#=vms����v�y�m��:t�;]��j�:��u��Za��x��E"�I}�{�M�0g9 ��ڪ*���
�\x�����>轑 _�;!
�L!Ek��|maV��ú�ͻ����O�7$I"�������=2D�����.4X��l�&vD�H7ٵ4O�'�7p���fc��7�>"���P��B,���*r9¬�� �S��|{v�O� ��ڧ�(�:�v�kM��W9�(x�$��;�ߞN��`�� ���ѧ!�>Kle]J:��vF�9����_�V��3xA7K�;3[B��YԼ����ω0,LZ!(p�m��ӹT	� ����Qci��Gd�ω�>}�TO�<�{I�e����?�d���&�%;��=�wcx���5��U�؇�c��'`����ߣ�@�h(�q�gv�I#�����\io���nqː�2d��mU`�1e�d�@�	8�}1r��������N	 z�jh�c�2P>/sV�f&���=�A=�����"��]YTI&2�e��U��X*
�7ٵT	��+�.�� ��$�|���j�x���M|O����@$���D�na|�a�N�v��-e��5>G���=�O{*�HSW(�麪�O�m�J�y㓬�REnLm�܃g.�F�G`Q@��֨�ޔ�*ؔ�{���?t_I6h�_����oV/N��wG'�P�gG�&'�g��镵e�Q��9XُD	����	�UuZU5ۓ�[��ի��S�A�0����|;��Ϗ2���t��qn��yM�՜HK�l�OQ������{K�>�mle@�1��� ����!N����m�� ;�O' �i�]�� 㠷�.���Ǟo.N}�v7=p;�z;g�r�ٻZ3����s��;Z����7]cN���E�^��	�v��ɮ�(�ԧZ��(�]j���V��ܒ�`�ۄ�	�j�^6s�����_��m8�syTH'�6�d |Os����U�O��� �]�HN�9,�5��I5��߬y|��L��*o�7��@ �}�|I;�&I.]�2��;��<R�������؆�z��A ���=�-�]W�	�&-^�	�$H�Fv)"�`�^��ʶ0m�FU^ȉ��>8�*B>$�ד$���ӗ�K��}[1�mTI��b
e��BE6L��=2@$잚2�|��rj��9[�2I5�g�oOUx��xӁ�Pш�=���E�A ���#�{q���1@�ks�7�#�t+�1���������^���2%TgI�������������b,��A���x�%��L��Ḏw�0�ʻ�5|�}T�iP���ۮu��'غ�[�Aݵ�a��]�4#��r����;U�=ٶz_fQ���{���Vېb�sq��ILg#��[�k�zh�"%�Y[	%]�Y�_m���(p	Cj��$����@�N��H|2*)L��Ӏ�|��5�=4"��p�l����ĵ�%g�>=�$	�_N�A>+�1���T1@�(���w����H(LEl��� ���
[}u�͗Ff�5�;4I>+�2U	zQ���+�L�~�P�@>�v�e�t4qں8�0�l��0<���8"ں�=�a��͈)�ʁ	�=�S92A>7�;4I$���AT�+)u=횪�F�ۙ���%k�h����Е���n쇩o�{{���n��]q��0�ϻﭷ�Mך\��L$�a6�پ�'������ ���o�uS��rR�,y��=�7���r�o��U�=qo���PД���u~W��}�ۢ�@Uϵ��2�::� ��d���đ�ѫ&�7n�"��\g	�=TH��5ϸ���0Jl�Y4K�<�k{�c�vh�O��|d	y�|'$p��
�%��Ux�XO�$8E�\H�b�"I�{>���y��q��=\�OMf�x�Bۍ�	=�&A^�ۈ���]��?^O�m�X�ۋn�cWm���i�v���\
�)؄؂ �,j�9�I0���Wen]Q$�����$����"��4fr�\fl߭Ko��ܮ�+��A����[&A靟I+J�;ї8H!]� �{�9�&v��*ٓ�:T���ob��b�5�Q��>7�dH ̅T�қ}���-��J���	#y�� �&`؈MD6Y�����UE�sO!�<�"O��[���t�`zP3�3Q��s���vn�f�a�l��=��-5Z���}����xoU����(�9f'f�Y�+�w��lESwH\>#.�L��*�a�-%Q�ˑ$7zzk�T�M���$�<�2O�"��� ���׎���s�7Yȅ���W3V�ޣg�e���9u��x��y����om�������@�6}�y1fA'-�A>�����f�Ce���r2:Bv�dpA���F [=u8H)��26��\�dMwOUU�[FaQ�٭�/��|�	�h�H��.賈0�禉����F�@+�;b��$�ǛU�I��^Z� Z.a��h�����Lh���xٞ�|H'ݮz��J댭���]��O���|f�]P[jngf��]q��]˟uy����:� �v�*�$�~ IO���$����$�`$�	%H@��$�	'�H@��	!I� �$����$��$�	'�@�$��	!H�	!H�$ I4$ I?�B��$ I?�B���$ I?�B��$ I6��$���e5�;]/@;]�!�?���}�����  h   (@(   Q@  P       (     P� 1%@� +킀PT �(�� �M j��)B�P-��B�	U���% )"�TJ��TP� PR��$"�EJT�@Q �)  UT��F  �	B�*R)D=�
�� @ }r�T��d �״B�w@��M�X�S��Q�}���A#  0{����*�� =�UY��&�v���U����xz���{�װ�{5:�q���Z�.�A� >���AT")JP��S�"�Z}��=j��:�H��*���*S�����_}���w�	휱ӟ�=s�q�u�'� �$` � )�w*����=�Q/�(�9�=���}1��>���7Cp(��c���P/�vhz����Lw��PR��`W����� Q@PR�1�U
���/��f��`�3]�UL:��n�{�T��W&��	W��*=s҃�kOmT�Ӏ�	 -������W�����ҋz��wzW����z�W�U\�.*�w�E�UU�:��U֢R�!owJ��$�C�ʨ���P(��((U
���ْ���/��֪�mu�[�A]C�d��u�{5K���B�ܪuUV���W��O!F�K�*�;���!�7�T\yH��������c�UTOlUW�yN=UZ׋�;���JS͒�@�D�� ���AJUE*����$�lUI�P�֡>�v���(+�Trg���m.�U֢����=���Pn����ҢJEI�  p���]����TK۽�����z
V���� � `tF���# 4|      S�����        �~L$�IA2h�d��i�	�O�*�M����      ��R�d�D ���  �0�?�i0�T�       iA�&Bi�#Bd4���Q��ѳH�I���_��s�W-�>�>��k��l>�u��>93t�䐄�L��1
~D�	 �a�T�@2@!l�	 ��A��HB@&��������s����?��y���0���IBHQ����HH�b$a2�X@$$m!��{�����o�w��N�$	 ���<ـ���?�|�������z�~����f)`�}>������c�_�Ս ��_�6_��<��7L]��k��mXz�jSw�be�oo=�U����$*irv�GK,{O	���bp�J'6B�Z/�#5����Ր����3n��Y�a���	s_=ioW2흡\�_hǡ�u v筓���BC��oK�����2Nh�!��l���KI�����hǽ��N2aF��$ͦ��j�n	��"75%����ഖ�p}ܶ0���:��k���>\�.��P��[���8���˺W���Od�{�F��V.�����GϲK�p�6���5|6i3�wwl�zZs���	PGu�9a�[��'q�@������wE�M�lO54��r�Gv��t%�te�%Y�a{���J�|yq
��Ľ�X�6ˬ���f�������Ĺ���-�}�%��Wt�������x�of�KdhÇvmgv��j�5�2��T`v�9��z>fɗC��ֈ�p�1 q�V�9���ǵ��CN��.�h��oOz�����3���k!v��>��2.�|��;����7 �@�M:"�-�&�
bZ~�Ը��^(�u�G�!hq#CWob6^��"j7jQ�{y#"f��v`���dB�Y��r\a�.�sw.���%��,lL;�!�q���p��!ݐb2svŝ����P��;fĨ=���a���
�{�P�IٗǸ��mG��;F�`�p����vKp-�r���:L��Cft6
{s�7�+_v��`�Up��%���Pm9-F�ӻ;D���;sXxNm�:L��|^Ǆj��v�g��: 3_.('ط&�bնv#�z�v�lro�J��N�|v���ޗ������������n�\�l���H�����:�\��9[�;��US�C>�I���0|m��C�P͛��@qom.|쮲��bˎh(�F��;��|v�+���m9[��3i��6����/bnN�}d7��,��h�����9od�v�N�J�=�J�v<��ΐ����c�����_��rT�Óu�^�u:đw��w��������Q̅�,\T�c,�1�J5�uXI/;x�]b�9[Y��j��M\(�B�����BA�5���>Ww������;��-�̻���]�ιE�VqVܚ{� ���O)�Û&�:�C$n�ݡ�ǎ[ȉ��Wʇ���wEpd�H=嫏v7�4�����w�v��؞q�\O�E���8t˽$9�7"�!�s����(bI��{݄��}�
*n��5����pJ;'>$^(x3d���^�&��TyN�wq��Ʈ��ְ,[�zhб��n4ED�r켶� j��O�%�ho�X�
<N�k5R�>�ݷ�n�WA��2�p��u�u��u���W1%;���4���&(�lw�#Y���
�s:�	y���8I#���A2��ge��9fsM��r�e����)�D=vn��ñ<9���]g@��n�m�=���nT�l�V�a����\v�c5�2����.p���8�����\H�$Q� �}Am�p2f�<���t\ǽ��}��Y�՝�[�r2��J݄wA²2Dp���[��o:��&rt�5�jέ�Ζh=	bk��˒��Rq�M�)ݖ�=i�sG�N3�|v�϶�>���b妝�wm��O'��wn�iu��F>&��,ѵh��<�`2��ҽ-d��}�]Y�;r��8٭�u͢�s���ˮgn-Ь6��p]�"��{�M	ۥL�$Lgvۯ�;_[�_u]��!��P�<�D��@��L�Cn�p1��l����h�X���nIlWG��/���j��"t:u�;����{��`�����fq\���죨��dO:�1��>�y�^Nȷ���;�1�C~:����F��(L;z�{FY�8��w�����������ɶ}5C�*�sx	ŠE��� �+�U{��ܙ=���p�Q�Zmmު�qG`�5,����F�2�׌;�.S���f�r�([������5�97���Ej��h�of�a�Gc�v5��g��C���m�E�yf�N׽�1��������3q��xڄ8�����g\KF�!ux������H��&��/�x#�+!D���x��ɫ4vB,�Gx"of�u�_#�:6�+�U�`�Ǧ�p좃Ή�v8�`���n��k��:���YX�l�<��E`9���ɑ��X�s^�x�oU0��U��Y��@�m؇r���P�(�� x��J:r[��;����	Gd9M���������>� �C��J��m�b� s�K}: ���ں9/W�9V����{�8{������ЕbOq4�b���b�Q)�9<RP�k�A�.F2����r��ؒzw������1N�ef\�2aA�l*a$��i�X�u�x���C���X�9�e�K�*u��%Ҷ@��j���q=�l�T�ۧ��%!�N��ٱ�8��M��U�H:�"z-[�Sع���qN�nt	�H��w����9r_RJv��	-Jd�\�;v�Fq �؇vs�q�����Tl�O��(<r�cǤt�s����6['�ıb���x��bV��ﻷD�N��BJ۳�__/kXLY�n��v�Q�l���[$�^�X�ݼn��L�ӡ�5<����ܤ��F�"+ts���x]362�vMl���e�^���R8Q�",��XV�y�e�pMK��v/O�
ӻ�W뾰����r`�M�ɼx�\�,v�e@�\�ϭ&:�,�+r�����5��SWq��Ñ���:񽚬�V1�rH��[�^ٗ�0�eJF����Vap;��e)���o.��F��];��z۔s�{{����c�geǎ�w{��At�eioN�d(y�Ink����(>�@��.�����%o"U����0��[U�YI/H�pwo���X����4�.��#���~��e[D}��u�ќ�Jpn�V�L�4����2	x�sq}��H�m͚���&�Q=��8�٢���{�=�8�Θ�\>P��t\Q�eK=f�4�G9�����Y�^n�U�^���m�wJ��ZY�a��w<R^<^ٮ���&Osb�s:��Y���ǚ���Z;��;���]���e����(��C��m=��rBD���{u��3J�%2���&�h���$�i]�$�L�'s����3� nkŶ�;�P+4cƻr�簀 K;L��q�f�֧�f�04�.��X��%5����s^����H�sWb���#������}p�&���4���2,���["a�������fpH����KU`�x-�u�!�*k�0PN@no#�M���3��'��j��)Lѷ�t��vN[�y1c/�9OkIb��qm��s&U���ܷk�ڵ�{T땉"�.NѨ3�l�� �񞙽ww�n��{G�78`-wwu|�\$����o^��֮25��� �260�)�jLa��'gn\t_/#��՞�F��~��4b�Z �i�4d%��h����j��T���L����o[�p�	�OL����{+�dv,��l��nAX\��t"�t��ǚ_sƷ陸;�r�t[�,(�ԻX���#[(]�m��]�f��7t=s9Z��!wL} z �� ���6�[�㷱雚�j‖��S`��I�:�a�4jL����#�yR�m�x�<9�x�v�tcQ �`d@���B�`cm���-�����k�N�C���;�5�9Qh��ئ�t�%SNB�9�v�3�f�����s�b�3�8��7ySt����K ;¡�q�;�����w&no:�+�J8�C���)Vֹ��"��a��+���N��
4�K��ת�����rk�*�����x��I�M$8��ǃ��ӥ�go7w����&�ɦGi���ϴ2��`�X�`���:l�w���9��>��oj8�T�	oI��E���`��y*ժ�;��z�<�� ��vv��;O�G���v^X�ޙ�L<��{����swu\���j\�[�J��l!���ߑ�FpK�f�@f�����7(�^PA)�a\އ����Q�[��Ų@T�ՇN���}Y30x�Ռ����c
�!���4���f�]r�8���T��{����㧔�S�Lڲ�ƫ�*�Wyc�2��Vt#&��]1`�{�KŃf�6Awp�C�R��u��2ŵ#X�/!/Y"�1_���r�>]���t֘-+Փy
;_\�Wdp�G4�.67���v�w�V4a$�C�+���;�JG�/)%�EbG;I5s7&����:��X�T+���7t���GC���!��q�s;�4-Kv�z���-*��������2PWs�#z���B{x�ۛ�gs�M�����7���)�jx�sq^]��O��Bq@�pVa�z\�q�L���B���A�l�����ƞv+���.�|���6D�HV>�
V=�o4UϑZV�w^�;�#gr�(�)ڑ�u�ڸ�K�V�6��O��\���fn,޹վ�d���S8ۨ����,�>��*J;F�+{����|�b�(�j]٫���v�%67����r�]���P�g��)5�ӏ;!�w9o89�>��٢<{]��z���hec[M��ҖM�_n�a�C[�iZ�Rd���h�� ���8�9A�@��e�9�W�n.�b�D�0��6��$@rrgxr<A���lg��ҩ)H��;&q<�\�u�vLx�}�>�p���2cު�.L�,ֲ�8gb�h��T��'Y��<�]�t��Q;�d�KGaJ��B&;�+n��v�(c;f��.>��)��3b�jtYL"�u	�i��!Gz�7u��EX1�s�w�e�ta`�c�]�/A�M n8�r�{t06]l!��u��h%�iCu���^�À��`{��Ě�.�.]�9�[i����xl3I�z�A&l�؄�=���86�.q��F\�"k��B�:�r�5��+��yo1{����w��85�I��S���^����iI��x�Z�'3��e=w�[����&�+�5��si�O���JJO��x��f �+5�΁*2�+�Kv<!О�@^S�h�+��j��ߪȭ
�n��F��n���+y5�q"�]�F0|>t���+;�5�;��wzt�`}3Ѭ�I黤!^�Z�)���2J����ON]R� ���7�L�gD֮�:n��Gf���D��n{��]!.�p{6�ݩuYJi;�K��3U�:��flÜ��Üh�����)�vh��E9.<X(e�c|"��nv^僃Ʉ���vꜵ���۠ҡS���\��#���PY��nA��-�Y�UU=��i{8�¢���"��m�7x�N�xd؋��v�oYɯ/j���8;��N��Q���0��3.��;6��q��k>���?'��x��	��!����>=Q:�74�����ף���<!��@�Y "�,!	R��I$Y
� E�	
� V@*B ���P�RHBB�! *BVH d!���R"� ����H�(I`BV�Y XB��d$�@"��H,) �"�H,P� �X
�BT�HAb�a Y�$ ��+� � �d��HJ�$"�BRHP��!�
�@��%@	R�$	BT�!X+J�@�B@�!� , RBE�@+ �	RH@Y�??�������|�������D�P�! �Yǹ�  @�+�	!>���g�C2	 ����<7�}G�����\-���<�:ݙ�*ŧ���6�K�PSAG��)��T�j�e�^�G�e�~Wv,�);�.�5��=SPL��Ƕnv��{'��X(��o!�=�|�{4�Qƈ�w�gv��N�����s}A�s�g�_c��>���c8eƲ�,���Zx�9q��{��홨h���pe(�,�@xge3m~�c��D��]�;<l�ᝀ7�/�uu�$�o����nl�۪R=�ͨCq��n�S,���+��dJ��g-��:]�+�<����{�����!�=;����}$W����,��{�d�g`�{�K���g�Q�;��v���/4���������_��f���Ȕ����+����XBK]�����B�0"�gc��ޢ��D�ۮs�1�������J�,Ә%�e��i<�̎ٻv�z`.C�]�gw����AP���| ���{�6�Gn���P�.5Z�4_l^��Wϳں��������N��u� ��U�8���>��V.�[�ٶ����O��Z�}���\��>���T������(��S�o���8v&X2 I�}GiY�ߵ�ۺO'y����#�x�S=�K�C�_���Y�{x{�Գ��硵r�����aᾫ��j�7;�3���nnS�n l'$ټ �"ǵ��a�`ܶg~\��Ӛ�ѽ�?mx7��x�2�xhn�~�jH��}��>wȃ�.怒v��ґ7hď���J�̽���9�W���X-N�}������+ô��1Vg_F��N��j�P�6���3׮���^�!՞�T-��|����{/
��v�N�=W�u1�x�3�]�V�>+�<�G˟�L�9Okxb�^�{OSN�u��j���V|9a�-l�����������yn���ۇ�j���f3���Ć{o�m�5q�q;^��qY��IH������=^��%�k�L�2v���:�8��������ƾ��}��tRy]� ��%�yl�؞�Pã� 7���0��jg��EȮ���P�D��v��n�4^~��Q�3s\C`+7d=�j�t������rk�iS�K7�:�A��~ۘ/Iq�)�o�8�z��z`�Ҳ���8���n5|��6�0l9���=~~�3�N����f��8�w,{����C-�;�C��Z�gK�ss��[ngb�qn���=�^ö���.��_�^(��Z��g���R/���3c�< E�_�썭�,I�73�q��}��afX����6����sM�i؆S���YE2G����N���[ӱ9����u�7���\̝����p�|����x?�j�q;\���}��}�ǰ/���X�_'$����r���s�w�.ٴM�G���� �\���PŜe	sPg�˽����V�n�3���P�	v���<;䟞��i���ln���<�
�<���.�@�����^�����*q�,՛�i#�A��������_b����A�������v+���wG��j��2M�е��w�\�;�������垸i0�R�$6�����+���ǅ4X�/���_��h�h>���rˉ0pע�םs��Z�8g��r��;�C4�sܘ������s�@��z/+�y^�������/v\$��!��}�.N��7
<p���<�_���o�z�c�ۢ⒑ĐF��ѫğ|ݿ<=���Gwb�}���>���]�s��]�Uku���*f*�@���۴��#�O+�.;�K$W�Į{D���,^�������3�y��Gg�Kk<3Y���:y��=(�>����|~�QHz�?U�i����͇w�{4�?%-�^̡������Vwg^M<�<3yn�=E�2�p����>����B���#�;*]h�3K`�W�k�+�¯���gJ��T˺*�J��C�^�o݀��Q��@t����g����T��|�!��rћ�$�W�\��	�Hzk��H�o��%�<�T�O{�q� ��i��+3l{|Sٯ=����X|ű��bs`���c���A4'� ���Oޒ��֧�zﻸS��p��<Ɔ{.orC��{=�����5�����n ��U����v/#�6��ת��uV<n_�љ�
�xԞK�nۄ�ɿs���1tC�-SZ�A�!�pz�d�AZ�9.�C�Q��{`�<ǂ�P��E�S�\2�=��yJ�^���č��xӗ,�|�l��;�P�p�+1��r
�N9ض����Uy[C$r���<��;�^gZS׼�"Խ�F1��|.z��������=��֭�rU�ȹ ڴ��Z��'�E���܀�Z;<UHۧ0�N�7a���W�@�FJ��R�)������׸�U[s*+�-�&G7
إ�b����<�����Y�JSU����-G�v�=�l��۽���ul��@�ŝ�9v�=��}n����j2wT7|l�Fl�o꿵zٹ��)G�'w9�`�	��,��=�V��Y~���P�/-"�{ەX�;0h����=�'-����L�]���:f%.FdӠ�����'��>��5h͘-�ygat�����t�A��ZgJ�.b?j��뚮�!�u�����݋`哽B��A�q.�c<=�Z������RR�:x���oo�d�*]�;62���[v��g%��y�!�^�5�[�C���.v��pݙ.�x<�%�����}���5���ntz�s�����ӳ��M�E��=ޑs;y�s�OPp�KB;�I�~�o4rU�c��w�\��d�O*՟\��9G�&�V���B�lr���d[��}(��<�M���}}�gh���5/q��Y�ȷ�
9R=E��>J[u���X�P�����x�׆�ֆ�L�Jˀ3�4��^�ta�U�q��8�w_���v���P;��r�7P����[1�>�o�l�4��[�4d�[fhg��Ly��S�:tU�C�(�.�®G��}}�����m+��tX2=
0���ϣ?���n�J8�Ɩ� g�����P0Җ?:RVn{���n ����O��n���W&=�"��wsռwB^�Z7/��"kV��}�__zawݾ*�IR�����Ն�]�ƻ��n�����<��9y`?3{�|��������p/�x�{�z�:��e�dz�>jx�w�sb���^}Y�;I��	�}y���5;H�sf�p/.{���7�q��߱/I�R�A}6Y;C[��3��m[�(F���Q	��r;R���o^����Xa"�Tm�C=��u�m�ue�p��Q��3/C����cݕz����ҍV������z{H��a��}�O9�U��	˓�"8����l��}��=�i9v��rH�2솎ҋC�d��C���1$�B��N�,CՋ�b�{-و&�"�������q#�; ����L�{%���g�j\���>/�q/H��״a�x��=���Mr�уc��]D/�="�X�v�^9S��&��_6�+�[ŭ����K͍��}�{8��W�VN�Mb����dl�e��Ubp*p��A��OU�Z���A,_�r��V ����Z�z���o/��?%�z�hP���8�T��8��{VW٣pG�p�ݸ�y�uO|pS�U�#|%��oå��"�{��
�~G:o�T{�=�y�Jݴ��dQ�X��ya;ո^ͬj]Axߟ��s��f��4r�`���yNwj��N�sau�:�������a��O�OB����sϨ���^�"�7����z��ܑ���ǂ���݃�l�,h"�EnL������9u����m��>�n�;�uY�w� zj�ԫ�iov��t����XR���Շ�������\�T�Q
摆oȞ��c����O�:�ǱeB�u�6�T=�o׌�+½ln��݃"���;�T����!���&X$^gy�RM��'��g�[�]��v�=�QG�6Q*�S@gR���:�^I6�W���x��E�׽<a��ï�Oz�"l��ŸS�Pc��1V}钣��B#��� ս�͡3���v����/��ao��o������x&�	�;�=��h��T�0V1'��-|J���/���wP��9�w^,�o����Q�=�v��}g�J�'3��߽�kM�/os9|�4�U���{�٫D���qP�}ԌZr�#��}�����ɞ�ZW'�<��� >�"9v,4��l���){3C��ر���swc>���Ű��n��[7ӏR��]W�|5���x�5�s���[�4�P����Ư@{��cM8x3.�^˞W�VsW���ӞK���NΓ�/) �N �7/��l�Cӌ@r��Ny;�w��f���WC�;x�u����:L��D-_Kǩh^�s3O�Ƃa�0�R�a������k.d���q��!����M��)�wE�_Z��q�<���W�+������x��=RI>�<M����3���/�v�4��f�9�;_�ћ���˔�����P8�7��NL�4��	�g���|h�b�=��8y-tԗ�#�h��=+�h�ǝ�n�-���b����a{ZB_�MG�'�<�O����L�Xj�u�7g�y��z7�x?.����{w�~`.8V
�p��D�V�/�M�4������:7!\11Rh�I��C���Z.<@�3c��4iV7U�on�'��{΍GY�wl�?i���鶋���?X�6rCϽ�G��l���w�fu��^���ELD��8e��lqc�Azw���i>�-�)C�(�^����4�A]ŋ���꧰��n{��[��yq}]C�ɺ(K�1#žD��^���!ڨ�
>**���FQ�/W٠�N��f)�1;����v@���������W��2�ݏ�����ظ���a{�{�o��b�}_����'�eeM��n���0y��D���<8����`iU����j�ǔ-d 4��<z-��>Ƽ�����"��u����yze�+�`�~���yE4_v!�=�A���/���o��{�?mÛ��rZe�B����D�d1~�ە�C�H��ď�@����r@������s��f{�ݫ}@�O\�����T�n�p��>3���z��W�{�$8Hds��m�b\���&ׇ#�|njksT1E#Lc���{�p�����+ÞMv�y��5i�����Z`�7���{4�����F�I�5R��5Ew�w��۫=g��`%V
����k_�V�6�S۱���f��Y�E����Q�e)��m�3�|���	�4RB��;|~���#�j�i�$���3����=�v��������eO6}��"��>���/��hƴ_'���N����Yrn	��8�]�B��M�٦�bڼ�R�����v�sh΍3^�*�	%"�����W���ޕ|�ɔ��� s�;Ր��2l�Y[i�����+eۊy+?i�q�%��hVswS�\�?�;�)��#�+��kga�2\��fG��?ȟ(I@"���(�BipaX;JC=��%
gٍ���f�,掤n�� k��{b�מ�����{v-a��s[��Z��Zq@lch��4�,�W�����FĹiZ�����k2�����܊�V�'�;�u���݊h%L�������U��#a�����U�.�ٸнnI�3�LK4-AY���Ѓ*�414-Ё�+oh��g:���8��p�Y�n�ֱ�w��F�4��i��q�,]x�3���� ��i�C����Q]��P�haMI�Ba����Yq�i�*:Yu�)H�T1)�;y�5��Ev�q���(������k���H�Ik�k	4f�n�u��[A�m��X�M�d���#���6�X�8[� ���S�r:���)�ϭ����0[]���H�R���<��f-�ы��B第tklF:��a��-,c���r�ś��m=��r�c�H���;7ljm&�4���\�p����&��ʊ�A+7.����Zڡ��<��W�g� �>���*A��e��G2X!SNo��h,��d�Xa/�w.����Զ#V�\�Ê��/ 6pvGm<����@6p�6F�&()3hhn���[��s���@�"�,rp�.t0�Un{`��n�õ�����m�W[+M�&0��&��L[^llMp�B�m�VA�l�G�n.�(&�[20�HԌ0�yκ��(@uP2^kLnJV�i�b3Ŷ�צ;lt�nF��,3�lуsBΰ��Z����3�ss�΃;!�-&4�3\8��m�j3)ƇNԇYW�\a�vs.ժ.ݻq����C�!m��^tK�pт#pCl�nMr����i�/;q�wX�jݍ��4���@-a��S�#�T��ۉ�$����-����Wn��v�Cm��a,m�i5!�,{��9*N���x��8b�i���ηe���a�{uW=�X���u8W�;7�mnn�,{�mr���F]e�FsNFX�!/l���/��g����Y�0��
��+h�wo3��;e�R�Q���*�̱�p2��"�cjCj̷4�B��f;i���b6jJh�rX�u#פ�^��6��mm����ѩ%�e@Hu�룃>�J����=!WrӔ�GM�*hk�hF�;E��R6�P(X�/ ���@G���#�%�m��%��D�F�YrY�&�X�m�wS��E�\�X�WR��(�y�f�c�:6��K/h�M�ɋ�b3���)2� �66Y�K�e�L��Aҷ�ǚ���f:ǡ��n�m�ĺ�y�lR��ɮ�#�X��^���B�D�xu�	v/e��S����Bl�F��Z�c�JZ@�2�^�yͼr9�<�nl�����ëg�H����ώ����)-[s��<=���� M��\=k�΍Y��M��5��ݖի�p�bT6��g["�.a-��L!�BY����;Y)�";�7<�=s�ح��afu�3�MԆ�P):㜮�&R�t#wOg�K@�<��`����)*l��t��<��96u�.�q�@W�%��j3��	�0�aWC*�3˦�mֽ�\]���b6�Ķ���;��G��O�k@WQ�rsO���7V�����nM=������cu��t7���c��λC]v��2]���<x�O'8T-��]W�l����۵�'Dٞ���������V�v���ۄ{^�\G<����"�����OQ��ǳ�mU]�fk�2f*n۰��b�{���V��="����"��Ѹ���{BٗY�d���V����8�CiSK�Z�#���.�K�N9�p�b��aKZ�Nɨ�a {r9uW/���E�^b�z�U�(jJy�]ۆ9y {I،L�V��x�W]�8��qz��1�45�j��dJ��V�w)��=��1�3�^�	�v�ӧ��s@���F#�rFiYXJiMh$�I�4��n���Iz\v+��R��09�����N�q��W��=R)���M@���YRT�s��\����]���@�5۰���R�f�c�cr"Yi�W'c68��׵�v��oN+]��-��;u��s��G�%ζ��3�Yݛ��S<)-�b�E�+����ݥ�<��0�fd����Kv����X5!.��{KX��ݢP^(k���@!]E�Ɏ-Hk���H�+7:�l��"�N��r�z�ET� ���m�ʽ��逭��ʥK1&0j�FS�[6�j�Z��H�ۖ	+sYt�WMq{�b��b�E]���0��v��
�����ӊ���Ѧ];��m��]�8�u����)�'f�@�XB���-��4���[��f�L����F㳇�W��d�0�7C�;GS��-t/D*�R�Z2�ֱL�ݦe���;F���Ճ8�t�u��A.�����tV��;\�<��R�ŘB���Y��5۬������,-��m�B��lq#A�3Z2�,e�jl"���Мۍb���=k 5��0�Άk����b�%J��KŹݱS���=&�8�)��z����� 4ם1q[��#t%h��{����j6���u��Sۗr̽��:n {E�:P�3�iXa�uf�"��>F�n��r;���'r��6\�]�\ǂ&Q��L5�ct��]�&cu�Ui��7�yx8���Nzy����j�K@(ݚ��u�����f۰P� m%��	����D@�ĺb`mi�Ya#�dV�Vmeu�"��
�Y��Qt%�K�b�Sg#�d��*6�e�<�q���z�#��Ɠ^�tG/62��g�����[����������:<�8�.��n#R�c�n8�V�;pn8+��Ka��Q��Y&zӮ�GcR��:�<����c�r�@�XCM�efŀB��޹gi��xKĆu3l��ֶǒJy��\:�џD;�h�YM��g�Žh:XCKb�M%��f�5l`�\p^�`��� �m&�<�.����s�x �1�;[��0�2;�e�EIq]w!�.u����n� �E�Z�<�������]�0;E�Kqb��:.G@�2�u6�4�.2i��L�	ū���V���Z$ԷU���!�Z��eu��f|p�I����Nֹ ȼ6a�S)Yu�\:��j�=l���pQ��hMv��)ݧ=���,+qn�ftԚ.����\�lD��h�1K���c@�KԠW��"�F M�hG\M��w5��y�4*�eST�[��:��fJJ�2gQ[b��2���o+�z��7mӶ�# �c�n �����Z9��c(c4k��]�k�,1qk��3�N�ې�}x��Vi�Ĭnu�\[�^�<u:�,���u��`ܽ]s�C^:u]=�.;��Gn��(ީ�.rrd;3`۶M�n�Ғi��lV�]);��7=��c�]�.q�V\��/�$��7�����n���%�b�ɑ�9��+Z�J���t��;
���E�禍���v|�ī	hI
�����77!{3�3�V.���n�f��f��u��io1֗\�XW'M�ٲˁ�8q=n@[�������cgLj���w[���8����j�4-�jmu���`atu�m�讯/N��Ю���`W&ܳ&m��	Xn9���G���:���B &`�u���j;k�%P�qmp%t��ɲ񣱻R�i�� �N���Rk2�L8f.��*��2�`�(�(���E�Z��筼˝1��ő�i:Grt#�8،�z����:�k5��tL�V�45ucئ�3�緜8B���@���+�.례
��Z\�oL#sX@
Kt�7K�] c�-ژ�iQ��cit B:�.�uūb�+�m�>x�=��V�tv�r�����/u�ϵ=�˛>�,��!z�q���^|����m�ˬV�2�[��,Z�lC!BkB�1ڈ�ń�Z�D����I�&�\WG>y~��Qb���Rm�"�8�*B�b��AAA`
E�E+4�-	U���%b�0�YZ�X�k,��+RTP�$��uHM9eJ�IU T���+"$�"��H��a���d�ŘVJ��*�VL��\@A`��@�Y�f%d�1l�JZT���I�-�,��X,Q�f�0\���Y%��`iY0�	\�&�"�)+$J�BT�6���U,$RB�(З�,�I��E�B@X(8�+ ,�� -TdH��X,Yb�kE
�PD`
 ��C)+�`�Q`(E�*��J�FȲ�K�:�Bu�"�ѼvaGCe����e�؎;j"���V�����;v+��8�d�h@��1�i0�����U"��[V�<<�x��D�]�t	H�KT�y�43)FLݐ؇P����cn���\M2���˲6�,�kt̹ius�M���]c Y[A�i�
m2�:EtU�4� �L��Q��ʛM.3�q#�1�5;�D�kн���	�.޸�m��p���DT�4�6��B��s����sbʹc����t�^wm�v�^���.zvB/e��^�]��e|�ݻ4=���8r5�Dû5�qٶ�c�g����4e�BU�gI��7 	��N,{A��:��ƴ��lٶ�&������jn�,�c��\�;��=�ۉL��5��،X�T�pck��Rk��X9l4��jhg�nۓ�[��uα�(IwҔXcR����n�]�ncv��㮸����۬V�<�ʏ]Z����FRZ�k�1#ɠ�+d�ug��1���Ѳ��$[\��N��:ս�O��V1]�b=r��\���U�XX(��\ɺ�X5��:�l����#!6*�t��U����L$^B��`<�Q�֞�E��a^�<��àV]lK�v���cK�HݏU�(��-���!�c�ϗ���ˬh�z��z�X�
���It^ڛY���FLq7X�Z�+u굶
��Uqr�MN��.\�kq+�]��>xx˥!�Ѧ}A����ŵ�c��,�F�q��t�^��J��;֝&nc̤$q+a�r�%�$��Ӵ��Ym�-�h������%��@�jV�[KijKK%(K�h�����Q�h�d�����ڐ ����@e�e��������l,i��b����l�(KB)J5��Eq�^8x��`��T�"'F,�j�b��X��Pc������~���Ė������>�"b�	$�.�%^ԇ�z+n�/�`	���J��G�_@�f�凪����nxK���=wd�s�{ʉ&�T~I��T~���{2̑)��a#$F�K5NH�9q�	 ���w�]՛�K�J��R($���d��E?�r�'7����Օىc��&��)$�Vr㤐H��m֠�������"N�\=�6.r6�F9p��z"I'߻ޗ�l�P��r��T��y����I ���۲%v�A����'��mH��݇V�[qu�\�I�� G1�b2:�ϟ>��P63<�#�U)�\z�4In�mߒ�#�օ��/����	9O���IŸ��ˎؒY޻���_�[����m���$�o��U[%{��5�^��K�|�2f$Q�?wz��8���+�ͣ�u�n���Ӫ���ҐH��;�M�7{}�"M�+��ahƫ�=<(sM�q�9�Li$�K3{o���	Uy�z��i�� ��t�$�{{}g�F�ki4R�#w�E�w0�^�͉$�-��$����>I*yʱ7s�uH���yJ�K�~�-[��TS
^���I 3�)<���þ���E�$�W���y����
S���ظ'u��	p��h�)�������c�u���b���+�����M��R.�I'�7/|�H�O9U|�')5��f�k��TI$nv��y.Y�ꐙL˖���tOt�ͮ�R[O[�]&�K�n���"PT�$�+��=��jĢ���)�$������@%KyBI�֧�ڮ�3o�{c��w���[�AO����xwz��Tk�f������Ӟ�:}w�V�#+H��*iOXY6�g+r�w�/�A_���Ȥ�
�r��d�M��	�n�r��{֨�n$N�_]�$J�ڪ�I%��Gr�6�RGĞɗy�TiNm&�RDj�k��Nb��u�\�e/���z�� �����%�t���|0��R�%2�"

c�^;с�L�^2�0����-���>|ꕼM�����{��T�i�	|�*�"4�}�CԻ:��'�%O�C^�0��6�1˅��� �Sı	�������<�I%K�JI��wJ�A,SG�M�yq3[dȒfT����t�A,�q	$�q�˿uu{4�I��R($��T�R�\p�Ē�.�{ޮ���T������$�eJI��wH�I���X��
��T��A9=������۴4bF�i�m�����^F�˰z^Dd	����2�%yGr��/_�@{G�NWm
J1j�����7kyU#_$Nf�߇�������t����D�I�t�$G7{o�y��*q�����j�����ڝ�Q۹��v%�RF\O5o���~~��#\/��$��W��K{{}�$֙�=Ҽ��N���wJ�C��dMόr�o{�G�KE��6�?�7��A%���*	�����E���5�{_v9�>���}ƛM���H����I.�ݻ$�-b��pֱ���� �򸉤�[���%�µ�I�r�Gj��'~�$�Z�F�H$��w�$��9���^�V��$6��RQ
���$؎W��뻿qoRu7�G?.�=���$^�"Nn�߀�)$��t)]}��mr�dK�ۯ�;_�����r04��4e��ʧu�x��͌p����7�"$��%f�
%^���A�V�/b���cX<�s�f}�,z:��Q�\i]1�<1������/�3���Hi��T�m4���ɭ��k�{��)z�*u�q�x�s]l�v�AF^���8ڦxmю�ՎV��9�g�Aꐁ� ��Xm�R��Х��m;�m��q��
�h�^]Ylt	�կ07eR�!�v�[�#A��I�@��V�j�	�w��UH�A,��>	$��r���������t�$I�v��b34����J�� ���g��;#$��{{}�|�I%3�
E|��/�y=������l2$��9rԛ���$��	��EF�Ϧ?$�7��~�)$��u�%�g��#M�BJ(t.n��|!奺.{����J<�I��P�I]t�ӕj�ǹ��A_Ww��b'�Y��̪��US��I,=r�J��/d�}�w��	 ��UH������o��ª������֧�����-�5� v�&uO���D�O���>�牶l)(�����I�D��V���V�\����]�u��y�F,�	�*\�����dD�R��o9+<q���AC��;H'n,�'=��ʘR����/*-��|�{7۵\�����xy�eW_!C�L"1�����<A%r�	/�B�]2I~^�y��oG���C\HM�܄ݤ��H$N��$N�=}^�FG]��	��uU"�HZ�O��G�(�L
N���dN����<i����6r㠒I�ݾ�3���Kqe$b�UI�}F�m)%�	��_D�'�wo�S^`����%�;�T�I�.��K�ݾ����ʙ��i��!4��9��[׳�lR��Iy�7a�����?~�_�&�A��2�fS��""ov݅�3���yK�֨
E���t�,���S*��;���� ��V-�w3�QP�KF�$��~��r������d����p?�R3g9I� �	fwm�'�,�{��N^v~�@�({>���Y�����y-{�o���a_�S��w��z��S��a<~	0�+��3���2� �w{��<�P�tx�-�M�I�w���|VD�A-Ų�A$�f�߂H$b�V���=����{��Ԩ$�z��J@�-9����I$��SW[�`�A��|�	&_����I�+{�l��(��#��P����ۮvK�K6�]��Rn������+������4�iI=;��ʦ�Iwn��"��~)����~߉�^�"$�{�һ���I���V�U_:I,L��Yw-IM �Iݻ���$Ŝ��'V���$���O������l),�˻��JJ-�t�A.�)ng�����g��If�o��IAG�������H�H���UUT�Z�)l;�%�Y��$I ���~$���� +��ngB��Uc�·@��N^o�-�Yv�����f������병]b��x�~$w���<�ƕ��a�	��&��:I${�OO1b'���<�?W���$��UH��B��*�#�̡&�eh�Cz��5���f��y���]�M)R�v�+�˾{�>�Xs��s�޳�IE�A�I$��Ҡ���n�)+��yP
<�_R]xD���%%:�7�	�a�}b�K�]�|A%r�h%|�"I��x�e���u����Q#	MJ�	b��D��r�A�I��U��[��0�Ir��$��v2-�٨��8R����#"�8=�i iM�H'le�I�$�{��������ϼ�
G�}�"D
Fj�ꪠ�$�;���F�:�z��$��*���%�wH�	��}������X����`��~>�{~�G.�x9��i�S�=|gӝ�/Y����3LxK��Ü�֪t���Rv#�K
�-H�e�z�ڒ|W��ƥ�f�&�.�X��Lkp22ݖ]���^�m��`C8�3�<�mg���:��ڧVŘ^���9Z�����"�h�%�ֱ���I��{5a���S%��3b��mS]R	X`K�� ��:֋�3�.e�LL�2,Uf��;���,�M.��2WU�]��8s������{�����wS��D��i$�C��=���:w��^W>Z����K��$��
\�H�r�7��|��������&�$��]�����t�\'���,�G:�m��w/���F�I%ݛ�d�%y{y���]Ԧ�If��I�n����v�ʠL%E.�-U]1آ�=�es&��](4I*����$�S�L).����'�� 7굲�3��Zh),�]]�	 ��A�{T:Ĥ��Y���I{���E$ig(r���o���(I�u��c`��x���q�m鹦�*7��`Y�(�)�9UW����۳�T�RZ'?�\���:�I$�[������b�;0�rvkz�t�S��MQ5j��㥌�Zx������L��C�/ˇ�;�ߥ�-���l}�P�p�d	�^���۽�)~�I$����[p���{�l�H�䈩�~�����(R2�[����A*Y�$�J_�N�I¯��$=ۻ~�Ȓig(z��R5)H�`L̯RX'^����g7�� .��-  ^��d��u{����r�h.ݾ����o�*�TR�Ry��%�Xz�D��Dd�0C7{��$�I*{ʅ"�Vz㤒���:���A�o��g��m�<oU���+h�)�Shy����~|#f&��yn���y$�T��:%|����u؁˹�U���y�F�j��PU���)/y3�T"A'0�.!U�޽�A%�T����*�]2h%�\�ܴ��?_�����	�M��:I�.3�W���O�`k^�X_:�:��<��~=RSXtc#39k坧�W
��s5CS�� �c����s}-��q'�����$:���=�7'w�[��yb����d�y�g�z{��z�Wy�x���me`~�up�.�>�#X���7K�h��Gh�٣0�����>��Ӝ�J�u����]�3NsP��䰡�L�������_����q}��/t�``o93�xw�=�nmu=Y�;^��A�T��S�:,����޷I^�뢦���)�7����S�����*�F�m�Ռr�-wt2�eP�q�-�i�eF�b{�֟��4𸷖����U�nG��$nd�A���Ʒ=S�o�<����+������ ��Cy��o��%��op�Y�g[�ӣ���+ny��_�+�Z��ޛa�� 4C�v���E���i���^�O�ڊ����tn�a�08�%�����x�l��z�e��8L��9�s���Y�pY���9|�D<�J�rA���� ��~}1���|I��̼ɞ��U{A͛1�&����IQ&ܵL){�=��f/y��8��4gF��:�G�v��N���G�B�!'3��=|:�\���ם���<!uw='��v��G��K>3|=�\+�u���އ��]p�5������
��@PY�,��$��X�gMH� Xŀ,�IX)m�� �$�&�H"PX�E�R(,�DX
��$*�CԢ��*
�
��PXV�YV
H�@PP�VH��a�+Y ��H
J�4	YATR`,�V`�(�*��Q� "
��,���,�a��PX) ���A`�X�
"Ad,�((",�Œ,�B��-�Q`1�X�,X�A@�"$Pc�sl@�!RjN�7�}��m.��˕�m��z���5����*_�M��]g'|�s�m`I%�:%$�-��������$�E)�I����T���VdiBё�y36�DJ	~����*��xU�-��=���H��n�|�'�{o�U6����^d�*6�ks����q`M� �p��9���k�>��<����D�I��	ǮP�$�Cw{}�^��TN�y�(M|�^�d�a�M	+˺�=�"s��T�^�qJ	�n:I|�[���y�d�{A�ySRK(S#�D���ݭ;U_D�A/f�߇�I���Ѽv�z�hI|�շN�A$����С2�H�	�H���B���vv�ɰ�3%�D�����U��|(_��v�z��AIm���&������[b��Ԟ���:]9=5�վ�Q���Y5�ʚc�[2�b?�_y^�&����	P��-9��Ѵ��쯥��]q鿌�p�~7���|�4���յC*�R3>�A��������P&����z�:�E7���mqh��+�B� �f��A$�ԭ��}[T]۵Gz��S�p$�c��M��Qi]Yw}pY&�y�}�кbn�
�;'z���|�/8rH�#z�� �9�0>-H��mz�<r�e�!gn�@O�X-�U"�p	��{����X�A��cʠ�û��ͻ��O���&F�	!?���g�#����N*���:�� ]�ψ���7%m�LܙA�;�%<}i����8�-1r�}�x��<�Ѣ����@�sϻN�2�e�y���o�SX?Wf�d%�������^����3����<[��aШSf�i筻]v��<���qG���c����Xқu�l�1�]��I�1u*�e� �vI�m��z:��&�f����b��9�Ph�T[^��;.-W�[=��S��V�l[�]l����s�n�=� ��*�ط1�'���ƭYĉ�W���t��y��Lb'��>��$�$�[��d��vN)���e����6Y����*�]�u�V+�ns���=�+w��wi�篺�e�a1���\��㳼��d��/_o���^s��;z��<R$���%�U�
T:ۍ����0��:�#{{�^��x(��p��i�x����3����m�F��[�� Y��W�v�
�ƹ�.�[��p �_S-�S:��\�5ۭnڎ���q�*
�%�����;���톃�ͣ�ٞt�z���1��6#ԡ ���&���D�nIv[ު'X����uTW�Sh�������=�*�}��c�S�����_3@������p=��?bsf�U�o�����H����TI߷��W7��Ʒ��'ڴ�c�
d8ɍ�[2��ͪ �}�Z�V�Bgz� �ު{�0�ϼ�%����5'(��w���n�_�~0c>JS�p�y�>f3u"Jť�t�xs��LbsZ�R`��%�$�gW��.�ώ{;�'G�\]y�K�!������j�絞��	U�jӷ6�T�������9�n7�6�R@^oWԁO�Z +HO��+�/��Q�G��.Bh��(yO2ʽ���޿{^ ����'�)�*��]��R��h���n�]����	��p��LӪ��s�ΏeW�u,.j��^�tye�WIJ��'OQg�q�S���U{�uG=�h����|>^��'�A���P$��12��EBcn�̥l��Rq�v1���&�����L�6<���B��Z֕H%#�#�@A�u�������d%FƮ��T��� }�ު2��~�.>P��
���\a]�3F[S!��Cr5����~�oƍ��F��ڪ U�)�wz�7��o��ޤ� �E�0�����q�}Ϫ�#�!���U�;�BF�?���U H0����%[��z��)��MHJ��9� ����^���";W��b�	�u@��F�ȓ8���9�zI@��4[ޯ����Q6U?�H{Oy��u�#ܪϟ��S��'�X^w��L��T#�@�K���>���`�Q��2��7�"��y[����| /���P�����!16y�$���t�q�z/��;��@���q�
<�������o��͕��a605��&�4q᭯J[�"�u/=�r�ƂN:�t�>`�͹@�A��l�lw��g��hBWwꠘ̹q�ّ� ]�d�y����}����W~�@���Hx��\UۊF��r�����W��U!���n��{mLty ,��P!^w:�0����"a�A��kL��|[�t�v�{����)j��[�ʢ}<�a�&$q��L�h�F�[�zF�_��.Q ��ڤ{��k�WB�r��6"VD^Y��NY���
��f�;z��g�h���w���Y�xؑ�X�z����I�O�P)�ON��y�F�(4�RVRVʸ��e�]��^
Y�a�&��ʹ��V"1��0X!Jꬱ�Ks6�B��9�K�$vyŏs	ǋ���^X�d��m��f����[uЖ����3hV�nH�A��8lq����l�bf{l�6:䡂�i�f�x�9��u���p=;��S�ŭ����sPvq���żmR]v��������4(��$]��A{{j�E�^:��u���=u�@#��B�J�X���������E�$� �E�l��|����un����q�%�jQ&�t�*"��wF_�{����*�t0K/%@��#��������	sM�U}D��g��;�}#�ʌ�vx=��bA$D�aD�P���g���;��U[zGt1�ꯍ��k��]BG����S��ݣk��}^���T�@n�%��\����/��2%7.]�9�2�� ���TiOj8�]�^�_^�>$e>�2"��E]��TL�{�J�^{�[�&��sܷn�u\	�<g��^?g���>}�U�*vz�˿yfn�Ԟ�8���}�����}?�"��}?~���~��
毬˿}G�y�nH���b~�{�������s|��E^�O�7�
����Ke�́wL.���䯞0]ߪ�
�x�[�V�{E�A�N�֌	�����wz����؜��De������R���q��m���犄i*!nO���6��N������׶�8R�����7PL8q.B������:�{��㈍�̚�� ��ު .r��B���,k}0=T0����~Ww����z� �{��J��ۄ�-�Q�o2��M�mQ�gM�qz��V�=/n\��g��=��Mn^���p���#s�=����u��~/p����볉�#W{��j�>����>�}��忿g�]
�߷��uZ��#��u�&�ܚͪ���#�:P ���Pj�4<=��:6�v��M�1u�)�2�ނ$Έ�e-�z⏁*�U*@�y����?Q���(���j�q������璕�������Λf����������s�Y�U@guP�>��C'�՛u���"�:��cMF�}�ई3�U�_r�z:_f��@���: ��B~�Sa��-�ş-D�%�T�ب����rg�e+�z� S5���1�Q��2�׽Yĕ�x�nz}@�� ��8y��_S�Ҝ��ʡ���>ꂫk��us�G��&�oڢ�݈��\�$�y���[��ߜ9��q�����|�|>��3��Q���)hD�����?o��35���ʻ������0��T]{;n���+?�l��ぶ\�1�7`�_D�Vܗ7֩�6�ٽ�6�e�̃}'�3`e n���Q��rpz���.C��<�)�
Gw��UW�l��x�nt�(������t�K�\��7t����%�F�P���H"f��뉁��ɀ���9}3{�@��k��1$�ב3��=����9 ]��wov�(�2GLBun �h<��Q���OĞ������ɉI\�(06�)��eҤn�S�/˲}
�:���һ9�6�����}��zTm~��^�,S�3g�z����>���g�4��b�=����|�T�T�{�S��7�8��{�j��{���2��1�����2��0^�>�GSC�Q({��h����*����+�JA�/=wy��ץ#�B-W�ކ�#��og�RL�S��SF����TꥶF�y7��[����������W��}��^~�;���z=g�x�ެY��mj����t�Y��(΢�cU���S4^%]�wb=^;ŭ���{6�ઞ�,�D��8{�*�MkӃR�L�|p�i+pz47r��W��0m,"(c�Y!VϫU���n�qJ;��=�G��b���:�ݐ�߮�b"{T\�,,{~>��(�=�o�{����{�o��X����|9�Y@�O����z/�3z;����3�e�!�� �<�L��۽7rϬ�=N��;/�1r�(|Ŝ�"'��wt`1o��%Ʉ�{����j�!;ob��l��j��%tv��-��j���Z�mo�y�7��:���Gv�3{i
���@�s���j�,ݣ~�	�{���Y��3�¼fB�����g&��]/~zs;15��L��(�R�B,�U�����%d�"��E���)���PY""��H��$PY���S@RE��P(E �%jE%aY�
V�,�F�Tc,�`,�*AH�-�)"2��m�#l
��[B���-�**0����
)PYY	Y
�2�("@U`T(��A�a+H����Im+ ��m�6��*(
��Ued�BTZ�Vu���<�F�b$�֬!Dօ�=j�mz��	����h�4Ծ�J8N��/Vq��Y�۠ǭu��Uq�㇍ټ؇B\��СW҅k]b����R$q�[um��L�=���sS�Qg�X6ٙc�a�R�f-���6�T�nM�4����.�,����kp]C���8-FdvU3��[��\r�X����3�%�\�\ s�7)� �y�O[�g��m��c(P���F�Z����l�JL���͒`�c6��Z�6�V$j�ٛ��6���sr��H��NG$☮�Ƭ����m΂����ٳ��5'X�ѴFn���x���n����v�tpk&����a3�f�:�`���L\�74m�b�A˞Ub�m8uRg�ejz�"+f�ق!���1.����OX�]Vr���c��6����Q�.e0S��X�M��p5���ۖ .��Q�pOjt��Z0��]��lS�FŁ1K��q6��X�nۛ2Mz���b��h�)�El9��E�l�Bq�-ؽG�3��]��<�bNJ�M��廮�d�ÙK�l��M\flmJA�*�	��v�4�=�A%^�>5�"g`ɩ=�ۦ`�sG[�t't�nň��ka�KR�Y�.��J�-mT��U�v��%��O/	��-�+�9�\�S�R��i���N���h�E�}u��&��۲
n���dmF��Ǭ$ǃMsȠCX��T�k���B�:�9������A��u�`��x���K�I��/gt����8ͱ�Om����<8(-bA9v��x=��mM)u��	��4kn�6&Vf؍5�M�I�wI��Bk��=fu3b@F�+�M�&�`	��������d��;���6�!V�6��6Ҙ�.�]�{q��ݰ�M��.�d�ێ���;P�M��<���)�ܼ�۫G`�uݱ���S7(�*��N5���#[�6C�1���[Lf���M=�ė[8���<�.���E�M7�y1�p����wk���).�7e�\R�������|��o߭K�g��j����A��	w��Q��[��S�M��t�U�Zs*"HjF�ު�w��S����_r͙�l ����
�sW��]{%��Vp���A'�)_mU
 ���w�f����q�������(`�5�H\F�X���zdY���Ϊ�)��$��پ�#D�����8Sx�LI#�`��|�����?ծ��������DA��A-�+��N@��@�8R�Ń�I��rk��C>����o�a�#-���ڤ �ͯ��G���^zA]�5`_gN���E#b'$�{IY���f���>7��U��o�����&{�,�7U�u`����ⓛ���u�	��e�g�yu�G����H@�:��������(���Gԁ�6{��j�xF�MCR6�[���'#���{�}�������� '��ifQ��4��Cs�.}U��]����U��|}=80�ޯyYL]�t�ji�Кl�26����v\�A=���:/�*�|Y�B��A����=���_F�.&�(�C=$l���ݝ9`���N"ґENy���bG�)�J3� n���M�X��+|Wn�@�^�O�]��'E���ܺ�Ñ����z�0Y��&����gf��&eZǈ�8��『θ(N�p,�����:�%xM�im��c�ˇ]�to���2�m��ܿ�J�I1v�+�ܯM�l���� ?V~�$���������k�,F�m��uQ��g��/o4�پ�woO�:�
V�
$���y ����s�<I'ٰF�u���!�����U��oU/WZ�ν^�(BZaF!���(�!K�C�k����*�ғ`� ����<HB	��o_f\��z��x�P���w��j���4�q��[ު�x���1ϙgo� A�IW�P���k<���V��
�1�ifOA�͡@���*>w:>���P|n�Q�Qq�1�iĹ���n�.��̭��WW5@��_Sp�j'����o;wS]�"��J�\_��v�{a��SR�r<���];�-�ce�N��+>����h���K�������8�ڤ�m�*"A�_�7j�I�5�\�U�Z���׽T���m*B,����{+�J�&�m�Q@�tX�VGn��n��.�e��]g�PG�
)��N���ު>�p��*��o��J�B�ΥF����d�)v�!32ߋ�E�y����>$��{�"Ge�|�e,E��N��T~�s��k��T�^�A���A'\0O��8���9#�1�.m�u<�*�$���'�������xҶ���µ-�������b��%zz� }1�	�wz��'?U�"g�x�w�~VF�'q�!�p�����c#��k�w��+�X���ai>�q��z��u�_���I'd�q�C�� ���-�'<�(���ѫ4�45��|��#q^53���w�V�LY�@��`��\�Itҹ&�Ҏ�4���r%�m�h���9�N�m����1-��Mm�ۮ��� 8��֧Ѳ��������A8�i��&�*i�{s`3K��+u�[\�#!ͭm��W���[T�9�Y̎���m�.�c�/B֍,s={��SjF���!o?�@7�Tg�^ϟ���J��"}���[T��N~p1�z[�
){=V=��v�����HQv���yuzu�_%F'7��4�.������B3ε^�ނ9� Nܴ	oz����Q0tD3n췼|X%b�H`"�����H��GU̬p�s�-԰N��Cc�ڎ��D�w�f�P�B� "v8E�ܠI'{zt;��#���6'�A	Q�g�f��2��/�Ͳj!e� �}�w��%$�#���I�۔Iwz�շ���k�L��'Ď�]
�}
��_�UT8wc�"=�������S��lˌK��Q�yŬ��&���{��B��n���d��R-b��:-9������$��\ȏ|�yЫy�2i{����V�,+t���c��OUPy��>B�Y�=��,�y��v�*5C¾��%�HQ�t�0^U���t�v�
'��!�B��.��'雴(]p��Đp�����A�K���d����]_W�osT�t�:�������>0Nݜrb��W#8���d��@�k�!�I���M�����F��sя*��.��T �S��E�	uվ���ڠA��B��-���d��D�L����}�,��X��T	>�>$�G�����+ӥ�`/u�a6�PH��n�Ӝ�bB�Λ`M6*��>��������9�a���۶�<�o'�]ܣӔ�'vs�d����~w����	 A�>��E}��jhD��ı҉��!�|����F%r�<��<-�k�S�>��T�mT_+N짨|?�A��࿑k�+�ξ*�?xW,a��J��� .��Q�G��XS`�ˢ�0�H��Q�ԑ
�w������Z���n�D�1I��ͯ�$�~+�UI����ꯌkjz^��+�uH@�.�L%�IM��L���hY�j�]�G���$��Bw����k[yv�[=Y;��KFC$q%�)�N�\���Ę�{���˳��pI��5��@�`Pԍ��U9�7*% ��� {�T���^�Y֩M�6�}J���x�Jg[��;�f�y�<�G���v���y;�N^z�,�ʯM������v�8KS��Ȕ�L~��[X��Ԫ��mSY
RE����.���~ڞ�������}�*�u�u윆�U�4�K3M�,��8��M>O���lnB��`���_ ��P;ٴ�{&��e<�M�z��Щ�h� �Ղ��P�/ʘ�n����۾�D���@W��EV�-��I���sv�7�j���tf=s��[yq�	V]ү��Ϋ�&7�m��c]��V�������G��uP ^��6d�+��1�t��vm��5#tgUW��LLToDf?b
�U@.�ڠ~6g(W�KkO�ܧn���է/O��&օ !_&���s�C}�����z�)����9�`�ÃڍV]�7X�v_�~����0/��iD[���h�R#h#�mA���^�Ҵ�\�آ&�Y���c#p'k��F�仅�ͱg*�Ʊǥ��u�Ĝ:��ۘ=�����w�&�:��Ghۃ2 VR͸��,b��c����aV ��/1�V��ƽ���:5�����IB�}vx�U�:��㢬i��͑��Y��^u�K�N��ܨ�a��$I��٨�b2D���?A'��C�By������`ϡ���wm*�=E}24��,�i�F�D�=6E�k���D�ns��]z=ǯ�h���Sk)Hw`��+�H��H�������RuH�wP�A&�0�I5�2�Q�~�ɭ����sg	�H�w�O!�k0�{�Eu�l2$ĒO�K�_~��+?�M�~v{�,xI��@H��P�sm-��[��Im|�C�!�<�PuGd�Ǫ���C��\3Z��R�������X�rO��UJ�׭0����oQ:���^ot��Z!{י�]
����0g
d˝��k&�<+5xj��q�5�X��{�V��}}�V^r����~�˖��&��/wޙ�@�T��1�ks6��z���Cn�޼�	>pl(���$�yߞ��m
$�����C)&��*s�㼛d�*Ad���9�.=�os��\�$�6�Na׃��93�9�+m`��r$�-�y�Mn��`V�*k���:�k����J VT�י�Y�J�T*���Aa�{����R��<G���~�K��O��߫_AI� �|޲hf�
�y�}��m`Xԅ-=��Ͻ����q��R
jg}��̸���@�9�&��
�++%Oy�Hl�[�z㾉��V_u�C,4¤�T��H)�l��{̟_�Y R�9�gk�^&R5#n�}��.n͵��N�i�$��@�00��b�OC-�'?�`��d4�!m �w�w�I�`V�*_=��i�
�<�3��`e�%����L�
��s��ɤ��z�>c���K�w0�
�����H,����>c��w�a��y:�J2�T�y�y4��Ԃ����{́�t��\o}a��9�8k��y�w�a���gfM��`�S&\��������Af�%e*w�ɱ&ТJ+H�]W.��C_��{{�/���Z^v���g�*�^[����ҳ-��b����5�^r�y)n_o����=��7_�W�=���1�V��B��ٵ��;�S�5x&�<�v�؞#�A[��W�{*O0�?>
��v�Vv΄��!,��K_���^����6OwL9���������<�=�R�"�oK�Jt��m�t��DT;܎��q�ۺ��wx��u~y�l��3b�u�_���%�9�k��ӳ��1|�wx[����~Evӻ}�mhM����#�I��d����C�숔N�kN���/Q�c�����]�]Ի�4H��5+õ�4�XRM'X�z��V�w�GCd�qX`�4�jnO<��mj��^�y7ܻ���a�m*m��������cjyO�����Б{Va����⟻ʗƬI��L���xs��K�rI{ss��S�]��|����1�]f�����\z1����fr$�_�W����=¶��;w݀Ǿ�{0�{��sݸ��\k'V��aB�E�`�j*é�����*����i�0��5���NjwQ�F�f@���G�{6ӵR��o��;�ے�]�{�w���S1S;��>~�۫v7���p9��n!��Q�Q��_���esc���a����g��牂�QَZ���l0b¨��E"µ��T��V)R"E"ʖZ[kZ���b���d�Kk#iYB�*"ʭ�T+FUQT��%ű��e�)*���+d�U�(�T�4�ҫX�aP�"E"�D�����X6ʅA`VURҭdX,Qm�P*���*�P�
�Xa�0�֢���@U
�J�d*[d��U��U�X�R"1�VUee�
�*+#hn�,0�V�j������s�0�0�%����Ad���YS��~2M��;����ɜ���X�˞@%���u֯o��w�� 3��>�`V�*s�=�M�K+(�c\�0��[��5�<8޽�Hq%B�=Ͼ���+����8�nr\cP��¦3�d6��T*Aa�י5�N�볬��u;@�J�|���i��ԅ��|�@�A�![��a�C�}��7������|nB�Z�B�u�E�su��!ƹ��E�t�)W�	���ڟ������#�l� �9�6�hT���+�5�C4¤�:�}�=��aP5�<ɦM���Y+*s��$؛@�:�R���0�8Ѵ���3�a �7～��w̚ꐩ�
���r�
m���5���%B��s}m�w�o>x����c
�]�u��K�u$�5��hm%��2���43)Ĩ�׾�p��[���<���s��H)�c\�0�0*^���Z�D�!� �|�~�,�'�r�7��@�4�R
k�o&�M�D��aXS�k�C	 ��y�w�l��}����4J�y�w3��۫���S�:We߯��ℯ���C߼��[�p�����3=f��v7�b���}�����'R
s�&���5|.̸�˛�ݕ�����2����ם����#%-���=��|���� �-�
�'X�y��J�P<�;ȣ��G�{ý�]6�I[����K�f���ݵs����������>��IM��:|������ID+%ea�י5���P,��F��Ǘ�;ׇ�y��E��o�I �9�w�a�0*g~���.-�.tSbNg^d�m�������^��u��m.u�NěBĕ��+���0�Ri
��s��&�6��FVM�^����=ד��3̓������&dnix�+ �Lm4�b��[@��&�R�`V�*{�+�<ֹ���<*Q��뙆�J��*��a��aO5�/Y[s\�s�e��T�7��G5ﯙ�5��6��
�YXb��	 �h�~w�l� ��� p�K�\o[5�� �C�kY�FK�~[O2��.vH��&��
��YFJ���2m&��ߛ�~���u�;a��az�w�a�� �u���&�Y(��FT�=�I��@�;�9���۵�pMvЃ�o�z��ʫ�U4ч�t�v˾�0�݅����k�P�Ǽ�[gjm�G�Ͼ�3/�~�����T�J�4�@S`-<x�h��c���@9�<+s��Smw4���f�X{Ċ�m\���ͭ�L�7]����?w�yǞ[�nįjMm�s���k�0oKmtq�a��H��:���L�[,��e���
[X,FR�9��ʛk��.Yf�:aXݱ��qj�]�:���9�Ƈ����ex�K�G�1�v�D�c��m�_����?&�˛�߂�>Q�;��CNR��-μ�&�HV�
�Ks�h��G�����t[��f	�y���%H nnAg�g����h��"�R�æ
�ϼ�I�+&��g���x��퇷��d��J��}�&��H)-<��d�����|�������|~��S�I�,{�2i;@��� ���ܛI�(���+.}���x�}�m��a�
��P;���Ad�*AO9�2�7����J�M��x��(�ڀ?���k�ݾ��AHn�<���[�+Fk�=�9�6�*Ae�k���u�e��:��X�N�
�y�ɶV�[:�L8������T��/�B��V]s&�e��c|�]u:@�T��`m��S�ý��)
ë�ft���|�mǯY�ƈP?.4�M�Y�=Y�`�X�%̷[�y��(��	��=�}�O2��.}��I�}�M��*AH)ߞ�&�m
���+�5�C	&�7�����3���1����d�'���2�VT�s ie�O���q�����X�˞d4�!m �5��L{�<�����w����_訹;��ysVë����?^>�燶kE���޳���B_�3��ɯ�B��R
^y�ƀ�l@�P+(�k��AH('강�}��@�Ϡ�~~�^�0&������1�s!�6�R��3L���@�q�o:�7�.1�������9�77H4�+P�\
4~����m6ܰ"��~�ɴd��o�z�qN���9��ɨ2H�<�� ��=�01�=�:��L�7��$�h�p�����3�h���ǚ�ht��ih���A|�Z�����FOz�yI7+('5�CL�%B��T<������3�w�����t� ��!Q�\q��79 c�t㋝���2([q�_���Q����#z��Ci*���=�0i�d��Ĩ{�w�l�������u�7���HvZc���7H)�u�!�L
��&����10e���:I��y6�@�������X����$�;����V�s0�*AIA9�w�l�Y+��_�^z��w�G~���,�[G��&1�ݕ���=ϸ:H)
Z��y5����
�|T��̋ߙ,��9��v�k�vu�U1N2?㼺�r��I��ٻ�a��Z�}S��������]��~ I�]y�i��R�
��X�0��%B�*>>;ɤ�íz<�i	n�~�'~�A]u��;����!Rs�d�0�R
�{ѶƤ�-=���yy���| �΅,��o{�gKc��_�y$�wg��&�h ���{�bM��ˎo����m��&�xF�9��P�40�%���M�M��VT��y�Y@�<�vX�q$ )HYH�A�5���&.�����6�&3X�6����m���\���Ε���rp�R�<�޲ke!Z0+X=��d&�
��]w�+2��y�Vhd�X��D9�:ɶV�q7�Ȕ��B>��U �GȀ��v~��jc�����/���G����(�<�F�jAH[O=��I �w�Oz{�a_/�M��8ɉL��'Q'3��m6�YY+,d���&ěH,(°������ΡXuT�!RT��&�6��FT����d�h���������R1�d5���<�n�H)�u����*Ak�|�I ��8�aY�ts��9��OQ��E�e����۹31;�w����`�9���]}��R�n����i;$�qg��^�N���������x��	*C_�&�n0�/��~:�Ksr8����T�y�؆�T+%Xuu�M�&������w���]uލ�Ƥ-�|��Ir��C�k��%%�덂�Z*�""@$d��7g�1z��C��Sb�r�3i��>��w�?�~I5�?y�&�8FJ��S��܁�6��u�sP�*K������s���8�)�}�&�62�Jʞ��d�h�^��ܘ�q�`t��k!�r��i�ì=|u��`^��Mn���
�S���@�m�+*u��0�AAD|���]�*کMo#u�w��Ya����}�sn9�2�l*s^� i&Щ��|ɦe��T�w}�w��q���;k�H)�=�@����jc\�0�R��|<q��s�:@�3��M�����0�R
s��&ěH,+
�]�a� �s��&�=뮵���u��&�R
s�u�4��z��.Lc%�˲���C�)H(w��i �<�u���{`T�9���
Af�s�0�42T���߲??~�o����Nd���V�>?���6���q��6<��y���^V.㠮��sx�z����鶫�g���| �;a���2$�a��a��)��&M�5��b���ю�e�9��=�ä˹��5݈\tu�gY��t�յ�5�qt��PI�â���봬%���<�ܲ�q5]I���<��Ͱ��²��ly�0�d0�����a5c�g����+����-�Z�oI�y&w+��⊔�ɮ[U��Pt[�8��Z��(�jL��	Eo����~�;`�J�d�+��ɦe����s��`l��]��=��ć��！�� Ґ���0è��s�&��V�یg`e6$�y�M���vs׭���sܙM��!ؒ��+
u���V%�T�Oy��m�q�����P�셧{��F;��E���p�W��1s�l� ��c9�	ih����
�[1_1�����<��*AeOu��
�2T(��s��&�m�a|��Ǚ�-����)9��!�{{���:$� ��1�aY42�
w�;Ѵ���ԅ���9�;V���۲��@�A�%���AG�BS>����ɉL��'I=淓i�
�2T��y�2m&�y�=o]w�1^u_=&��Y��
�Ri
���|�&�&�Y+*{�9�4��u_u�m�����+p�X� \��Je��P�v6�8��t��_�����ڦ����~R����I�l��K@�w�I��9�9�4�S�w΋��o7�<eN�ϙ�H(i%@ߝ��I�ýz<�Mm����L:b�7ߚJ�����ដ$��ߦ�|��r�p�_jVU��"�.����_��ig�跷�_�S^q̚��}���?
�s0��*;�y4��X5!e���� i �R�z3����]�����~���h�,�>svM�VX�R
s�{�bM�RV0��|�Ǘ�޳n��a�¤�
��<�&�&�VJʞ��d�hk���mQ;#�O�7�
�Կu߰�R�;�2i ��
���{��t�bJ�YS�oY��;�8�M����=IP��d�Aa��fq�1�pc7P��9�o!�6�R9��&;��o�s�5�N�4%@�o��m��������f���u��0G������y���H�>�EY}�����\6�%��^�I09�3#U�����!��Gϻɴ��R
y�9�ؓi�aXu��0Xi�I��[7�A��Ns^��&�VJ2�VT�{�4����.�Ò���Xk9��4ԅ-!�L����\t�9�I �FO=�܁��J�YS�oY��PВ���tu�掁�5�Ă�ӛ��:�����L:aS9�26�R��ri���!Br��*��t�c+�=������M����ہ�V�+�V�������{^Ո��y�}ԩީ��X�n��{�3�g�@�w�p� �>�->>9́��A�!Xu��
AMc|��|R�! /�`�&Jk��� �����d����MěB��,V���0�(�@��w�L��-o^�{�]�5R
g�y�lM�k�v�y���76�X\y��q�i�9�P�AqЙ���%�����%B�%	�=�z�j2T����&�n0G���?~��ݣ����A���$��5��V㣣z��ָ���vv�\�G�>Oi�Q�?:k:T���!�6��T�Þ�94��YR
��F�kN�o�s�$����)
��o9��R��v�Ɍ��˝��t���m6�R=�;��n���3ܞ'7�HlIXQ�aNy�j0�(�Ibs��&�&�VGq9޳�y��e:�y�x	���x�2gKs�E`m�9�R�
<�ܤ+c��g�4�0�޹���'��@�;�y�j2T(��P��w�l60�/}��M�3��7�uT�}�C������[�]�i��Vs�ɦVJʁR�]��z6��G�D|C�@���i~��~�Y��]��g�5�o��8�ٯ�-#Z�i�1^��s��x�%�&�7Y�]Ǔ���vV@���[�_�}��g�����@���$|	���	�H6[� �X#�Ҽɴ�ͲVVJ�{�i6����c��)��+�V�Y���P;���i��T��FT�<�I��|�Z���:μ>�!�n@��r�h�L��z�hꆞ�������^�a�.0�㇌5�3�s!�����y5���`V�*Y�s@m6 T�ǝ���{�4͉�oY���T9��i����&��m����C,6§9��6!����k�Ǹ}}�}y��gYɠed�*J�g��ލ�6�jB�{��� �B��k��>����;��E,H�5�I��YY+(�S�=�@�VaXw��w�c^x����%B�����&�6��FVJ2�9ߠ�Ȳ =6�Q�	Hh#�Q�l� �{�nY���|?$>�6��U�>	���`T�}����H,�g�k0Y׼�~��{�CBJ�C}s��a�aXk����U�p�ơ�0���́��B�����ed�]u�1sֵ�﹤
%@�=�z6��X�
Zu��$�B�C=sY��S��u�k�b�Y��>����<L�o�Gx�6��ȵZ*=�,���'ݔ�cU�ֽO�[�&�^��l�v���U���%��&h}}w.����u{����?y'�7�}!�|fQs��N퉦���Z����oۮ1��F4�he�M�*?*�fwvz���$y��ev����I-��Ex#�|��K��.8��Ϻ�@i_A{����̎�KK8{=��>`g�Z���B7�G=�`+��@_#��y�I��*�r�^K;�Ϝ�f$v0ߴ�5�B>̽�EI+n&�����6{^�)'mӳo�¨�}�Q�s۝��+��y/z-a�ۢ7iս����W����o����E��q��w�kM��g�x�`��ׁ�U?g�M@^[�b(n�]~2�Yۢ�Π�Qm�U����m�״^�u��Z��ǽM�Y�ޏy�!�K���o��8�݅��GU�d]���x�S6u6x�T^�{=�����jf�݌M�u�`ڏ�/�dLۦ�LH""�
w�x���5/L��!�K:'�>Y�����s���!��I�<,ђh���~�=6[�|��1R����Nt{��P�P�7�㝋A�\^ݹ"~Q]�kn����ꋚ�/\G����X�X���iD�,0�
�h(�
Ʌ-�E�a�"*ˊUň�E+
��cD�.�10�aU�.�K����Xa
�+J)QJ�,L���E�b�ұTfqJ�p�*�� �iF-B��QkL00�.��E�+��U��ѐXe,UEPX�Fe�\H��8�b1L�C�=��y=��Oc����'
L�c["�0�[��"�P_;r�O~����G�I�P#��0�Ri1�xLń��=���]j�����p�o3�r�W^kKF���la36i���_pmM���&��j��l�4߻/�|�4�k�ʴl����1Mv���:kÚ@���P�4e�N_V 9��\�Ӹ1�jBXT�� 31J���d㧥�+N'��KY�F�x�h�t�u�6�Y�R�JZaD�U4)Z�-J.
,�����a]�� @���J۞c���3o7�g�:����<�F�{Y'Y��<�Ѡ����pn/6l��Я�utE����
�oZ�Pi����ܗ.u�m3@%.��!#��ї;���t�a�͒��O<֩5��.,����65KV@��c�D�I��
�K]�E �h��I��B�[\�1�"�<
M�(���먌G]s67�<��1�O::ڵ��I�8�-\.���g��[X�����n�KB�7EU��mѕ!պ�x8�Fw-��1uخ5{K8��N������S���tg�z�r���E���c��j-3�M�5qQ�:��i�ѷ���:��M ŏ7a����N.j�l�����1�b7b���T����p��q�M�9uWRm�N36���Y��]F%ȻhJ���q�n	1o���Ǿ����k9n��^�q+�l[ۭ9��ִ%��v�d�W�W�#�Cь�;	���::�7en�P�.7�f'k��]#+і�\]TM���1�1��6�M���f1�TM-�iQMbe�m���e��T��2qq��b5�ݫ�[Tڧ]r"a$�FL��n8V�O�{�/����1�m�h�&�u���ld�5�+��rC�^7��wZh�z]�.�Z��JEl���s�hƹ�k:������+<d�X+P=^<t�FУWTX�&kcH-t"vPsԒ�f�{]�E�	L�(XD�4�l�a5���׉:�@�;u�x�����7>�t�v�f��^���.�P6�8DęGVk���j����Y���]���}I1��ɴ؁YFJ�2T��{�bM�D� ��z���T�z�Y/���@�w�M2vʐY+*s�s$�Y *���:�e�����ʓ�H�RC��&����=;7���~���#�k�=�2�
l@������f�*IP�|��2�;���V:�:+��1��e��9�o!�6��
�Xg�g&�VJ2�Q*u��ݥ��{��G���$|8$7w���AH-�\�`�`T��t��5q"� �#��W�w�[�s~�߼7�?&J�S�{�&�mT��z�T�B�s�w�L�ַ��ͽN�:����1�y�m6�n=�ks[�%�˲�6���i�!m���MnR�4P�s�o�q���o�dY "T
��{��f�J��*C��??~�r�u3�DJ)�&6�L��������݂�Ü�����z���ʆ-Ο/O�¦s�d6��%Xu�3�Q�����s��&��`o���<��T�M������+b������A0ܠ �dF� G�~��n{�޺U�Li�P��c���wL�����Y�.���2B�ղ�T��k'��[˲��7�����Gm7�ט�z�>$�g>o'��hT��aXS>|kPXi�H)*|||u�l�ed��������s�!��>���jĎ��l��jsh#���T,o����G�o;s�1�Z�'��(������L8��L�UER�]e���@#��*7z�MgT��7�7�
�g-$�9V3eU H���*��������H��S�|͞^�^w��!*$#�2��1���N���Cc�f��8!��"��<� ��E쪘��E���S�����%;	oL�����7���$��@���j�H��ݸ"/lʙl�=[���Ɩd��f������o�ijk8�����K�M{@�x^~>L��s���e�[x�í^wƌ���Lǿ����ݟ�_Q����C�,�l6bwg��ρ��k������D��&�[b��Y�e($�
'@�J�	�8*����$.Ϊ���	�|���MYz��%�Hg-��M���p�`�v�d�^K7.m�鱿>���|�1�/n1�f�*@O������>��z,ʺ�ٜ��pCMD6�Η�o�gFz��^����>/����i�C���R=��o�zt�L@�"}�gz� O�X|觎�.MoOr_�j�.�H�6b/�I0�k�G�D��R�:���H������V}<�򗟿vG��Y{F�]���槪�H��$z���R�M˺Q��mʵ�]���e��肔7�˺ ���o��H93j��t���1;��8����g�:#`�^Wz���}���m�A��r��t>��sn��"��.3H�L
Q�*rcz��n&��v2�9�����/�F�7�R�5����z��c=d}Ѯ�� �4�u�C ���w:�B�\y�Ƿ�[H��4ou5Hɹ�g�?\��*���p@���:�τ|z���`�����X�s��>��S�Q#��b%����9��	7�-{��Y����N=�K�}/�`���i&���U|H���jh�O���'T�a}�T���������/^�ЍV�ޑ��ߩT��e�oy��\��az��W���x	X������u=d���Ж�nj�1����A�bM��j�<CWi��D�)������\-����ڸЛrǶ���͆%�m��u�) ?���xkK���;Uƭ�-���:.M�;xs�J��kX����p9�\rwg�Y�63��'6��!GY�.[�Z�ж�,q!�k9�]C&�{v�Rۧ��h���9��m�k���ZG�0w.A�m�N����$}�R� ���TO[̎��Ǎ4 ����r�D9���&������;{��ݓ�!^mU �s��7��s�P$��V�ʒ�_��v��37�|͙�-���E� e�O�Fu�}J/
P�a��ˁn̬�}�s%���e�/�Ѐ���|���ɵ{�h>���x�Vp���7�+���Wx~��B�dU���uP$�����G����+��������5n�0.�zzy��7j"Lͦ���gϖ�">fPٻ@�~w�C1ys��̡̾@�{z1ڭ�� ����ow]5֚䑠)
U�5��x�*�\j{�x��B;�I��&fB��K��m:�W]_��t�ug)��@.���wU?  �����~3�/��3����H�t�d�&�Q1��^s��O��I��V@�׷@�ݴ��sO��/�V��IO��ˤ�؎�y
�cޔI?<��Go]Uc�{s������(Dym!��MK�"24h}�tU�}��#�y���uT���� ��UʺCpSM�⌍�k�~�HT)�������_\z�+ƹ��:V��Q�G�����H>�j�w�U�;W��8�e�;/)*BA;:'ʍ�^��a��<�$��پ��k�k��&l&��&�G�^�Q���Bk|��Ԓ-D����d�ιD�J��|�b�s(���_�����螪X3G��·=�A�m��*�`�3�gV\Z�O�zk#�{Օ�Z��I���I0�$�
'G�Wa��|-���cj@3/΁ݽ��}}�7�)e��%��d�>���ڪ$��ꮿ;߻U��%�@���7z��q��X(�,#m4�M5�~�u۴�Ś�p�ͣVC��No�l(�8�8��=��A��ݽTg�V�YpEO���W��DDF��9�#{)6T^f�~ݏE��}۾� Gv�R	��{ζa�_ �D�1��0L���Hٵ@#�VF5B�Gu��|�ޥBk��# �É�ȉ���Qڪ���}t�vn�!��+��K�d9�j�k:�޻Ym���d��VǾ�<[u���#� ����הa��O4��>_���~�	�v�d�M�N�=�U
�"�}G���ּ��@,��J�>��M�Ծߑ�=��i��BÛ�(�]�*�w/ibS�i#6'��I2J�F�öUW��Fgu
?@��ύ�3~��ك�n��9����&��	�Xq�h�\G��2�z]9�. ���t�<?��*����*��ҵ>C�L�`��"w��q��#��w�U�9��j���W������;�]㯓쨪6{k}Q��J$��͍ ,L�@����R�{>5b��8��D����i�}+�]�a"t�P ��1O�9�꣕���I歮�Unx6)��y�^�1j�P�/0׷�&���_���{<-Q�}a����;*׽���?�5H�F�1'E��+��q�tu�#`��tqbM����Orp[�h9m졪m���.�5Y�1j���u��I=���<�t׍X{l<�u���Sc�p�e�N�쎬�Bc��ŷ�#�rXvF!��to����oh�P����DM�ƺ��um�D��uwk�K�76�W\�s�#;�g��vY��u�u�ި-�%���b1��4��H�M�O���(3c����વ���@�1NS�o�g�l�Ѻ��*��-W-�x��+�I7H$f��Qޚ���jTw�(�MeB�0㈍K|�{�(D�բ���W��B1͍޺�
|��3��7e����ڧ���?m��I��P�	=��Σ~N7'�R�6ܑ�ՠ���kؽ���D	����U�wK="�r�:��W	�$N]d�ݳ�$��4�1����\I��:,bϖ��Q?p#!����u�>/7��7eF��3��tل�~�U4Y��ĚL8��UD����@�X��-����t�Km_�(�+�k��wԉ>�z-w�'���Ω;Ř^��K�/ȼ�t}ߪ���̙��g�z�y&�*}�[&F��*>G|�hrP ����/���Z�B$��㈌K�ٮ�����+�O���T�O�M�GF���*��@�8�M�w`�(�v����l>���$�}�T	"��2�|Ӌ�Ik6�:L/f�\WnΔ��s��X�%�U9o��{����shQ&��Q$���B�eYU]ݴ+�~7����p(�n�����t{3�}}�{�.�j� K�<`!�W�����F5^I�É��_Q����HE��G��O���K�<���܅�J�C7����g��V��E=EipfwxK���,o7�{tN)�o��5e�<tw3�h�y�%7��gs�t<OC�?;7�3Dw7��9�]�q����N(�H'or7Sˠ}]ӛ��q�0#&;ޯ�חf��/_O"R^:3����r-�q����W�e��T��m+�^��6#���Hu1l���77�|�����Ϥ@w��s�����o�7��+�V
{Ƽ���q#d�C�zj�N*���3�ϧf���zT���U�m��pb��`�V�Gq"��r�dX@AYP��7�������A�"���QUeU���z�a�ls��:��Omʯ��CE�盽h�۞���ꔭdk�c�7|-�,�x��1%��Vb/��"0�� �Η$�3�Ra��O!����7��{��h�������S2�3y��\��&|u��zo50N9��'�X�������;L��k�Ō����z�̏ԫҎ��}���y��������[=��j��./Ot���&�4�V5Ό�q���	w�����ٻ݂le{�x�g���s�+c�䝾�� ��	�מ<�d���S����u�;œ�s���������e�=���pq]SY�ܺCp��v��ƅ*�\�(�x�Yk��@B>����V#Ҥ���,*[\,o��\HS-��������x�:�l�ѣ/UcaE��-��ԑ��e��E��6K[ō�ǔ�V^�Y��YkD�ŘB૆T\"R����
����([,F^m��9��B#-����P,��a�L�@�1Z�Ԫ4m	ֲ������`,-e�Q`���^m,-�%TU	JU,B�kL8T�R��XaVҸ��P%�!+z�[J�o-��;�B^�X��eN�ll�-�[DS�`F��5��j���QR�
���EV�� ���_������E��I�B�D����Zks��Kp�=]�ڛ���~Z�~n��`�@$�Ϊ#�^�aRB�qZ��o�ҁi��W��U稜��(=�����[�T�%��m<LT�NYT����<A��E5E!�\���KF+mA����|�l@��u�Q"�dw{�@�&���{�@��xD�D�*�I��t��b�3�^R���U���.U)@�	��R}�D1���#B�F���n�ݶҾ�sO���*p`�;�B�
.�ƋI��Ϫ��u}+����B��R7;�r�ǘΙ̌�zq\|���s�w{؋K��8J���+7q���i�������Y�<��}��A�����?G��W�Wy&�
}�ҫ�����}�4<���A![�w:�;7�����:�D��32O0�2�v��m�)�m���tr�:���7��>�|������ ^e�@/{��T(��+ʾi�A}wU�ȎS�3,��6_:GM�N>ο�W�۷T��K���~M���u=�B�	7�x���T�^{�[���- ^̺��ޤ�p�i}�4cwed{��Gf
$ʼ�#���H��WV]\u�1��|g��jl�E�É�]=G�2�Ϗ�R�w[�q�σ�}T��ΪB=]?*ܸ����W7=-��4N��H��G��],q�����zSF�5k���1ӮO�]�qO�|݆P8���S�g��G��S��I��n��#�*A�V����q��c=G]�cp�FހQ�,>�b]��e�Y�m��JA�b���M�]Sۜv�z��a�<uZb�㷗���d�ۋ��R���D���09,Blv�K�ti�y�uڽ6��x��T�z���;�gu��a1g\v6�F�Q���Ֆ��$��Bm ōà�H�o��w�$)�o��U|H���B>~��Vt�x�#�'����wuQ���d��h��>$̾�&�V��*|� >��H��藒�m���_Lu`����5ȸ�n���G�A��vv�^��~��xB=y�HA��4�&��b�M�M�Q�{;�4;��> �?sM }�ި�F:��'�^���c�sHi1��pI�ۃ�n�;4����U @�ZO��TR}.��<�_-=��Fk�cHݲ����vxུE{t=�e����r<�i0�|=��I��B~$o�F���U���4��˼��ж�
}���U
�t�8���o��]Mg��d�~�j"{}��+ˋ޼�e�;��뫺T��t�&V��x� �T�mo����}�� 6Ow拓A?<�������Oo�MWV�.	�cQ-��p#zmE�y����77�"�g�+zH$��v
��(�Q�{�[�ܬ~t��*�� ���@��۵���r��L>��������Iݴ)Qn�<��oA켺I��P������p��ٿm	ƶuv��T��b�3�B��&WP�u�w��={i���3|t�3w�P$^o:Glbحw��{޺�O��3c-��N�����˚6����ҕVg�R��%HG"�j{���|L�hx�+-6�
}����;��@�2�ܝyU�F��.��W=���Yx���*���n�l�Ȝ{�/&�߽[[�B����u�˽�Ts�t�Q���W�Lh������#)~	vg��#߻�}Dj,Xc���F�Y�rV�\��#:�����uP��5p�YB@vt�T�W�4ˍ���(��^�U]��y+�{:ʯ��E�u
���*������_"�4�-�^@�nT�ƆΊ�N��O�M4#B�����V����X�p���_*��?{K=Ν��[j��ʠA��wUA�m�Dɍ՜q�N�kϤ��>�<�v�2(z'�m4��	��4<�m��`�I�Mg8O����6�ǥ˫��[ݴ�{��=��M �ѻ=�S��;�4I���DU�)�gw�>���|Q���Â;T��$=��C��jf����{4�9�,���޳�B\N?���ܞl��%������V�<G�_}_��2ꅐJ�#�\�����_���Έ��N�Xdq{}�v<����4����R#7��y\w�s�z~���7XM����We������a�e4{i�2���~Fʘ��$���� W�X Fw\��n��������t1R��`jۏ����~�lgVk�4�Ew��N�]P#>�AB�w[�q��'�xyP��ă�򸙴}�t���۴�(_V�W�I���?gњ�m��tGuwu�y{)�z��s���t�]�ԕU�90zܼ���t�Y�[()�n�-�@��B��|5
pl�B}] ��y��~�oP��V5���K����\�t��C۶0םz��Sw�X������b�x������c�i��������ޗ6�G�ځ,�M�f޵��\<0>ـ7;x�O/����F���r�# ��r�d���mv5�t��c������W�Çsu�5ՕÈ.\�iQ��텍�<�ipڰ�:������*�7e.Z˱YlK��Nj�Y��jץ�ux��UYnW���gA;�g�&i�q�(np�v=W<�gz��	�l���]P#�l+���:\�p~:vX��-���uP��z{����^�UB��a�����6_:G8��>׳�;.ꐃݽT�:�OW�W��(�6��p7n\�7�G�}�_f���������*B��p�C�#u��[�x��^�ݾ�B�x� .�����y�ݠC����E�[����|(s��R���;��玐|vmR��=�ܟA�z���i���P���+���3���X�sI;�zuIP�s7�3��/�� w�g/k�W*����|vg<D!��a!��ΎM]/-+bL/eu�w�s�r���ۿ>�����Bg�{�3v���5�����&��~�.�(2�U��{���z�$�}��"=��3�|�d!t�"۵�ׂ�R���o~*7vVΥ_{=-�nK�N)�� @vg5D�\���~���1����i/���
��*����B�]l�w���ςos�����7vS�'ă�ޔAx�Ժ��o*�6���u_�ՙ�/�!��'�2�S��;k��{X��+�i�ceA���m��cU���wU��#{��D`���R�꯫�����	�~2F���U��X^���t�^��>�<4��u��#f�*���Q_��j��w��Q����QkjɅ�/�ײ���}���ۋ{7�<�O��y�W�݇8���K�\	Hk�4����}��&U͵{��\����g���A�> �߮�M�L&�|[n��t�4��P�I=~�
���ws��|N}7��#�\ޒ�l��3�J�#o���<#�j�S�@�t(��{z��f������N���JF�O���l�CC�
�ʬ&���%�2a�K�t�o�hno�"c��n�/y�vy{��/b�W����uH�V@L�2�V�;J�r�_u���yQ"���v]P��J��q�t�Ƕ�X��ȷ����
}��;�� �ޤ�y�ݯeW�����]R���T,P�W�c6?��v��:�{��ΐ|��G�<d��L�u[�hv頼��X��r|Ԃ{���{�_mh�l�(φK�YY~DfF�V`u���*�����}ߍvt�B��Y��6���~��׊�uۃ�����H��Ԍ���|#���(�H�c3�����ݱ�����n�g=�s+ɴ�����cdt����|oZN(dq�y8��=ٴ(�I��р�v�T��u�G���H��E.]�������DN��>�պ���A�͔	�:0���z���	[A�30�3j���Ίj	^s�[b��Oz��&�z�|E�#���L�%>�ߣ���1]��Sޥ@Κ ���Śm1t��$���D1>+�$H`�ڤG�;3�<v31L^�K $ou�	�ta��G�=[ˆ�ߨ�jΘm[��8�̮�N����r�6�C>��g{r!�F��ڋñԧ�����^y�\N�t�q;��`���W����h
��a'�A��{|��_*	yO��9�<�'7o��nm�=�]�^��|�
��`�R�K�s��z/\dvщ���8@��d깬>���黚�9���4{=��Z0y��흿7�+'@n��5���z�t, ꛜ�<�y�?zh��d݂���vQ�mE�	uԤ�����s���^���̇y��q��ӻ��R��b|�HJ��я"���簡X��o��&]]�8���ԧS������{A�͓m�!Lm�^�2�U�Cm�`���ε4V��PR-��ziԶ����|�x�sz�{�Q}��7�B�3pk�n���71��sn��0����l�DhAҔ݁�V�ʵ�q�&n�y�i�4xTv�~�z+L�����ma�{�;i���>� _h��]�m��1�.�U���iN}=Ѥ��$F��U}�|��Cv4��\�:�7_:�B�ܓ-g��7��V��\����>+��猃U�[���.��n��	%�m*
]�c�w=o W{ľ�{y2xt�f,���G�.S5��Ը�鸸�DP�
�0U�"�R��e�-��ű�E��cU��UQ���ËL`l
 (Im!�ZBXq�"[-�AX�
��08�Z[KJ5T�P�km���E
�����jF6���Kkax9Z�R����Q+e��hZBR�H,*ZRP�H�e,�mh�`�*��1K�U���TYkZZ���\Za���-(�1
b�"����V�Z[�����e ג�-mV�h���%m�J�qZֵ�k�6�4iXgk�X���B��Z
���N�y8)e!N��%��mBҭqaqH��1m��R�����!{�al��{t|�F��L�]�T$��k�u�O
j�K��r˷�X��oR��Mg�9tp��q׭+t+�м�[�qɎ�A-ڷ���u�s�6�����\��Y�mq�6a�YnV*��svq+e��K�e:k��{<L��u�fڧ���e�ŠbCD�]��0���vv�B��6z��N)�q�n�u;*<X��·<n�v�M�e��V�Y�'�MƢ�^n�S3���M���0�����eN�S���ɚK�TC�[�ێIwo�-�����ю#2�IL��i�E�ې�%�m�8��6h��&���Դ	
ލ�і�C�m�LR�gCBet��(W\c�
]�t�M�ۤ�qpձ��&5&��l1�U���q,�2:�sa��u�zT�,��$��c7�	�^�[�;,]�n��[:�[�3��U�4¶6�훰�hZ��,lp��� �,�����r��ҍĶ �^A��]��۰uj�v�K֌���1W���,-�\�[�Vѱ��)����d��g�A�ٕ�-��$b���s���q҂����sd�b�y�[�^���b�n�`��n:z������ �Vm,�||�������:�Yu�zqS�\g��[��h癭�$,c���l@���K�/;R�#���o4�<T�<����k�K$Tmq`٠��;Yo$%qd�ؔ���	A6����		�'ae'ϵ���%åb��s���]��u3ګ��� mڳ�]���8�%箶9.��{���d�=lѡ�+^4�;dcc]x���v6�㇇i�iu ܺ+��T-cr ���8��������G	�47ͺ�wI[y�r�u�{M�;]��t9�\U01���oN�[��L�
F�"�TV\m-�]a`a�"a�k�z�R��z���`K�7b��	Clm�q)�lqØ3�gqi=Y��Aa㱊�h���5�j����!����y��$��nrb%*�j��Z��%]����j��(?w����O��o���o@�$�w��:װ��/������44fc�M�9Ln\�7�_�
��q�t��40;��}��}~wҭ�P���rX���D� _u�\Gw\V�w>�v�4 [�u@�0��L�3k㺫����U(�Kyu_go-�S�{U��~
�}іF}��'�f�Q�m��ݎ	U ��z�I���7}��0��k�D($0$�RDcc֧k���7tt�:�s,��b^��߈� lk��K 2��W��{����xɯk���T�?��=}uD�g��OD-����҈�k��Ķ�Ƃ�w����^�wJ��N����mۚ}�(;� �ґ�=�|�k��n��o�>[s���~�	�~��9�j������I�RO�q��2���wmR�[�棔̬HB^�����zP_�,�AR;�q���?\�������v��>+�*6[x�멬����������H��HEgJ]1�_�>�����o��
�4��=>��7�䷂�Z�Q�5-���XH�z�C����^Ѽ�)F}�[�TA;��G��B��좽�� ��V�C�Dc65H��`���y��93��|��z�*�?����7/:��܂���~�a��vI�_U〒Au1�:����}Ͼ�/����<�x��V�>~�-���}�w��f�+��qv��F�=��7%{uD={W����}�;lp$����cā��5���|�L�q�3����@$�����Uo�H��~\��"p܍	>*Gc~����u���I�N���!�O�=�r�/����{�^E�
d7"4Tz���6l����-����9N)$���)6Y���UD'�Z�ݽ�[E8��O�.EԪ���A)���`S���ު�A�d�ĩ�uAo�P��4� [��H빾꽆�w�`l�B]&C��A�מt�f��}q^�v��0G;�W��<��\26��{���E��yY�����A��{!�Uu���u�K�˸�G���⭾�7#�Mٔ��O�~�`�N��3�8�˖�f�Y�ff���{�C㖛�$��t:^R�F�m*N����/=)��z�  �oP�K=x�g���Sz"b)I՘�8}l7c�K�g����N""�Dc2���|T��T������f�Uv����Ƙ���R���� ���㺩�=Amo���Q�]LY?_TGn���В͹ю-����`PB�Zݪ	=�@Q"[ѻs�,����!�Ԩ�*Z��@��ѥ�o=�\�t� W��B��2'�{�f��]�UU&d�|���g�#{>�>'"��s�{o{|���]
����(���z?d���A�dd����)�O���w�:���oＺOA����K�T9��n/P�6Qyu�^�`ZaC`�J�5�0�^���M�F\Y7�r�VS��&��g���gj\��^rn�'����ы�gI��Љ��@�mMm�#7#�kqq����^��K� �q�o8�n�������+�W� �ڞ:����^�n�d.v�l�
L�k�nk���&]kf#q�l���a��l��*X�I�˳��7�a���k�����ʪ�K��|���OUAٵ�K�@��T�S6��U_2���+�2�����"f�u��/W��v�T��:������;��-L�>Q��!���Ѕ9�@m��w���ټ��"��<2�v�������59�p��/�z4i��;�q��DV$Uu}B�*Z�2���� ���.��M�U H��"{�ꁂ�(ru_o��. �.G�4�L�Wj��^>��W�x��'��m�&v��d@�M�%��(�~���~��U{_�*�}KAN����څ?F��u�I�(�}���]�eXyu'@U_�V�����.�ocX4^:�U��{v����'T��{���h��_�s'����c0,s�7��o�+�:�W��������摑7 "��� &�f��g���$���0C��_�JJ=�K׷Qf��j���~�Q�齜W� օ����c��i���z����ުr�~�7w��`�f�Ҥ.��J��篟S}�0M���[7={@#�M����ca�k�+ψ�Ic\t�5f[�v���/¼�d���@'wz�OW�8��7v[ު&�Y�=Z�tƓ��� _��T���o��`+�3�o�˚��ʯ�ٮ����yڛZ���{Ԓ"��^���]Ez��p���'���zf���{�נ2�B���n^o:��1�֦j�||�~��RS�GN�z� @f�U{����~Q8�Xn��|o{Z���t�림����o]a�v
!��/�a%%ک@]�(̧��L�*��;:��u��x�W\�;��z�Ŕ�����b1�A��x.�mq�&�_6x.�t܌����SÑ�i��ѭ���T�\P��w�q��ʻ��o�_Q��J�9�),�`�{T�>�z~��u˧�� ���/C$�ළq��s̭"�M�Kza&�T��A�s��qٳ5;�v��Ԅ��î&����ۘ�Ǚ�?Qz�9��@FZ����j����5g}��ޣ��#꽊g�d�/�5��r.�JcbQ'�F#�M/H�[:�^�u�'�.�����B���,�EI(�������x��
�]N�@��	�o���ҷ�n�K��	@�"Wۛ�*N��7uې�Ḙ��9F6T4�t+�IH)��$i�j@����]Mי��j�;��_2�\���TES��R���Q��0@�z�tFN�R{����r���Tq����n� 7���Fm�f�����b��t���2E-D�}�N�Ǔ�|�g4p}馚v��Gf�K{:�^�o/b�)ό��ɔ(��mU�i�0>�<J������κT��!��	`�6Q�=����窕�9b+����ӛ�{�#t�I箝e�2��!TE��+�^��.�F����*7Dp]��-�.� �:Ŗ���<��&��M�ݱ]�'���k��+u��C�u�a��ƺ�G<�1�1�Ìl���C�v��``6��	H�@Md��3f��d�{uk�F�����Y#=��V�6r�LaF{)���m3��/�I-�@�f���3͞` y���ꆽA�C��cgWkgϟL�ͻ�������ު&&��O�h�cO��+��L~iS	)(�R��#�]:T߾` K��T����\<�R�PSN�@��3�|���$��J��)y*��^1�x�wT �ޯ��V:`��((/��=���W����t�/:�<WG��ﴽ�r�%v�Q4���,�ԍK����(�<V58^L���:�y��ުBڮAޓ}�����
���ry���s֎��8�l�r(!Q�������	HA�>&�Co��@��h'������P��t��&G!�I.�9#%j8�RQ�/�{��/�rY�,��}�HW��������ꡕ3/��~g�.���x���B3`�oV}ri${ٲ�6�����_W��Z��wtpߣ�mS&�λ���r�y���כ��V�Fvu
�M��	S��Af.��W�Y�پ�o���^k��\U� �뮇�s�����6���ֶ� �E'\�_e�&�k��>�J:���_�j��s{҈�S�T���4��H� ۬�,�ItX�n4]����3#]w����;��S��9�*+���޺�c���{��WUP ��W(:�֜a�2GA�����7Ϻn��+����L�]P�'gZUub��}�Ȥ�%���~��(	/��/VV����C��t���K4�ϕ��R�e�B���b�==;���3�;�{/b�z//?2�>�!oH6��=�}��e�{��񾜢�j�O���a��8���N��6�XtS&~���[��w�V6�u���u׻1kC3���;v987_�.�y3��cf13v������^�^���X��`tn�����5w��i��%�뗢�A�Ze�.�\v�^$\ة��~^���5�#�
��m�J�����wwo��{ע;�>�wm��^�Wy���Ǿ���c��w�{�����7��L�e]Y�\z�����'X���A���v
�c�wVj9���=��~\��=�������ݮ��w��a�
��{t���_bP��x�k�=qT�N�k�;�Q,��Qwy��S�O�9Ҽ��WU��~W����`�����b-F��3�0z�/L�)
j9^�=W�(=��L;�1[�L7�S�t�ښ�{�c�7Nbw�=�m$�I�V�E��"��Z���<�s�r��|�������شk���S�����[�ŧX}���j�=T�m��.[�~�%tˡ�ɔ��T3g���BF���
f�������^���{�W�{�]o���!�R֭�)Ul�`�qm��*-�!
[�P���iB�и�DD��B���,mF<�/Ye�F2�P��C��-
�KF�H�hQR����Æ��QT���*���(Z�V�hVکKiXյ�F("m1�E0��mh�[�ï(���ht��ǨFՎ0mR#iJ��q�8��-kF#+U1p8iTkb�Ţ+�A�b�R��k[lF�)\��m��L��c�-EpѶ��-����:��Km����h���TX��8K�m�-�mR�[�J��e!-�,�X�%�n)�n0X��`�
�F"�ԩ�,�RVa0%)��R�L�*8�P*�be����m+TXa���j��T��V�V�%�m�d��Æ4�YUUj�"��s�(��^܋��u�>k-4�L5�Q��̈_(A�{n�>�{��M[���L�P��0Hb�˼{U@~9��]Lx9�/AG����w��>7;�T�3.���[��<Ic���.��Wl��Ɨ.�������D&�8k�,���y�� [����y�6-Z�M���^���p�\E�����U��T��R� ��_\��gu}HB�;=�{3�e���bs8��}����$�����#:��>@���U��1�Bmב�ǲ%O��h��t�w�T I�x�VS�~��u�����w_h�:��ckPw_$�>�8+��uܝ�}�^��+�F�+�^�y~vlN3z�|O�.��D��WǟU
$�1t^4�p������HAy�J���xd�߭bޛ���q�'�qvk`�9���H�mtu�O=���֢*N�\�~.�Jlp����U���T����yG�l��WG�~�yJ��ު ���B�b�]��=��ھ�|�v����!�8`&\H��9��X�)v
��(<�"2Ν(�n��.��~�:�	q2؆�ҞyMB�OM��UB@?M�Fwz����N6u��P����L�d&߼��mA���G�[�+*��[R��R��cH%�ު����L�{��>��^<M3/�u��7r1[�k�yPj]�n�C;��q���O:�~�_�C�Wi��а��\	�����)�%����1\yt�f�.��䣴e]�bQ_E��v���^�.uo'���<Ќ-�Y.��26_�&�|4�F�����َ%���%���uhr�K]v���@�VYL���T�v�n�]�����Zc���]��l�n��{]V-�ƫX����h�9^V��r{7�[�9�΀���wl��G=��1��<w��A0�p��Q'�\���]#�su�<��	OX�Mb�
c0d�P�V;����7$΂�>�e	 *�Ѡ��Ru���=��:�U���¨c?���E�y�c�s���ω�����(���E��g\�v�����3{Vr ��) "�z;��]�Z�h/Ӄ@_e��3-�m�}3�U��wk~=�˺�n�����U��w���pu��������NfE���yϫڄ;M�X��/Wc3M�}�����OI�$�s��~ �7����9��Vp�H�۪<(�ġA0�r�]�B�,m5R��UO&m�]z�nFq������N�~/���\ȯ�{�y��ESc�Ǡ�I��`���m�ju�@m��� :��F���rL6L1�yv�R�6���B&�͡UN6	'���A�wMm����俈��ۻo^�JNw:���� )���E�����Y��X�;x��G�/�W�O,��
�X��oΏy۠@��ꯄ�<2��!��)�*��[X�X�	��CT����c(���&��}�}����>2G�g����ڢ	$K|`66]߱oS��}�H}�Y�O&D��ۥ�j��︛���5�� z󪀖�ω���V'wnQ�
�%
���q�P��.���{�?%���,�]){���6Ty�vzM5-���2������@�\��@+����U.Əv��~�ߵ����MS�w���$K|aL^����J*�uWhS�A`t�;��'�ba�wz���W��=>� �}ԫ���r&��J����W}�H�;*_M�ݽ�-�}9Z [��E/w�zTOƶ{���s�`�5�/:[t�t��TQ
�� �DZ��!����KR���FM��q�� >��UC1��o]W�k�ew�����H��":�ol��S�H�lb;�ԩ~��Ŧ��:��/a�8ВU�q��ݾt���e�Ϸl�)��s;�����낰SW�B�e��|y�W��H��oCp��o����LRu5U��oE���|ǆ�)~�#qT�]��.����o[��[�ј�r��xb�^����ĉ�º������=&�"[�(d���R�{w�U���#6hhv��nwR��=��P���$67A �pA	��1��j�&2��A�������!��b��}�t����T�Q�mfĝ��� W���F����jT�?x�}J�O]u��y^�� �=J�$vo5I�U�Ou�So����Y�5s�$tL��}��@x��w�3/�h�����U�</��8ВU�jqÎM�e�����׻T~�_����EU��
���F-G(��?1t>�ő���3�muW�����|�u��{����ѭ��釨˞-?q���A�Zļ���*�r"�_g]��l��G�zVu6źό����ixIs�շ�c��_��`��Ӵ)��C>�w4�b��FĚ��i��`�i�`�0���Ёt���lc��Y��"P�\� q�2=;SHAn.������z6q�{E�l�۫����6�p ��&�Ki�Y��y�3��B��¼�����0�����U!���Ƈ]n.��H �vNp����n�]REX�����υ�F��r��T �v�}H�~���Q�KZ��c� �ު��)�*Fs"2:�
�`�ާ��� ��ꯀ~���:�ڗ��J��A a�e�/�Wʏ�u���}E*��&�fn�7�
7K�9y��n|c��L�hT�X�&Gg��ʎ�u�f��Ng�[���UYcE�J�V)'���U%u�漝oUPQ�@�޹G��)y��hF$`E�
O@�t��"3��:]0�+Q�Pvb��	��~�D���"-�F���z߫a
��J��.��	V(`����{:��������/ߖ�tY���ofz+\���&�ngD��<���ם_6%\З��'f��7�6��t�+C��#���ު��*�S�����Ѧ`1G%/��� �o�'zyN��،����TԺ1�jT�?(���ڧfw����S��+����*�q
v�
���ӓ��C�58�#������ȱ\#n,`�uH�s���^��_x�R7�AzPl�q8j�@�[nĬ���^�Ƥݑ�8=��l��n�q<����� �ު/�sQ���RL2��J�N.(Q1+�[�&�B®���� ��no5H�r}�x+܄4�ӖɆ7\����G�z��"�˂Y=�u�jn���-�?�ha�4O��{���܇U������#�S�m���|���$��R��F��}TȰ���s��7��� ۵�}�U�I)ڼ$��נ+8��C.��ԨYYdV8]-��m(�� ��b��\��u:���E�FJH���Eg7.�<��]n$�)o6�51Hb��37_$�.|�����$������h�����zm_e*v�:���\hI.�9#̑e�.��s� ���T�� ��w��u�C��X~Q�1���ڡ@����CCo�on_�y�U�O�X�%�B�2U�ꪂ|�:c�����w�j�eF�}�ޣpAD:���He��8c��
�;����xj���r��w���������~��,W�/i�k؋\f�Ub����Jl���>����:�Kx^���O��,��Goz��l�m�;䕖R��K%�k	��ckR뫵�Pq\�y�����T�<�g��<O�ݽu_s-mu_l��V��pY:�(H|��S�k�A�G&������9Bwz��T2���ˎ��/�U��o�D���[�>/�����Wy��}.޺�p�/�1�=һe���ZD)=�(���-���W}w)�GP��5�9i�����UG�z���8�Du�A��d&^]� 37�ꯕ�f'�{6zǣ:�m�x�V&�96�/97��)�橓�p�0��I���%�e4�Ǔ}�ӆ(߲����T{�O�¶��&O��z������!B���:�dр��U��;|�)}��󮍘ѓ��}�u
;�w�w�6�٬^�=��-����z��x��!��/M��ٺ}����N�w��ɀ����3|A������8�;���Jou���㻇��yvp���Wwu͊U ��Ւ�B ��������u�f�m��-q@v/?Q��Ɉ��v>h�h�+gy�=���\��yV��{>dg��e�j�Lu+D�6wN����*Ɏ�ڛ�ۋ��q�7���o �,~�{�q��}�S*E�;�;�=�%<��=ׄ��y�q�w}Z�M�~�����	u���M	NN{v4mǨϖn�R�+�{�b�i۵{���,}��s^�]ݲoEӠ<�����y 10�>��%=q�<��Pdq�����q7$���#��]��6�	�M۞{'L�+(H������m��Vmb:7�Dϼ���˽;��}�Y�N<3�=��*�������R}��0t�������e�Mb�G��j�r���v�k��J���q���ܼ`�%���,C'�fI�Iִ����e����[2ʙa�R4�Q�d�����*Tn8�eL$Z�a*��+p��R�P��d�J�(�"�[Qjc�!X��E�.Xe
�Չnp�X8�TYP�	�-�d���
��0����YP�V�U\Z��)���LZE0��0��b���`b�kIDX�H��Æa�Kh,���F�3�E����p"
�mFe�PP��X���	P�h6��L2��+�cn5R@htid�V�*sԽ!m�;�I�$X��B&%B��b�
��*"1L5��\RT�4��`Q�J�b��C����߿��=5����1��Qk�<<�xh�g��M��hwh˺��g���u�s��,�p�����gC��=�T�\&�눡���7�0u�:ڹ8�[
㢒��R䍚�$D�6U�l��	�`�0�M�+��^݈a� ���ne�=��,��j	� �@�͉��,q�I�l�y/֍](�vhjm/7r�6A���]`n�\{'7A�u�64m����ݎ��^�sջ�uvv���Xw^Ŏ��n�ɸ�ug\v��ҽ�q���d9D�jZ�]�<���7��G*�����\6j�vnr��v}��)��3�GGVי�r�7,t%Ł.��(ts����=S�6M��ӄ�!z�Ǆ�c����8��^�sd�)e�/K@&u�tH����Aۻd9��+{�C����t1Gl�j�qj�ZM{	0gvx0PA��-cv^��8�E��#.6�ɗ�v�;&	�hK�i�3��Mf�K�`U�q�Q@��k6�\�kd;n�ݭ�SC�	�x)��e�5֑#fMX �!5��f]uمB3t.\W`(�nrxl�R[0����;i�1/c�>��u���-��ǢxF[l�%�F�5q���R��2�����#��b�F����Ѧ�8ƛ�qŬ;��*�TۈaՌ1�ͽ�͸T&�X�[ۣ��FZ蠧]�mڸ���-�,��K�7f��J�'�������v���UWX�f�ݸ�`�۷e�*E���U�э �v��Ԝ���v�ǆ�����*�����sr�NM��\�),�=#�s<���lu�q�Dv��n��y8���}���X�c;dIo,��z�8�(�5 ��g���p[�A���5�h�N��ɶD����)_!q/8���r@���1�R�LB^���i���陉��f8�Z��՚0�̳٣�ta�G�{6���竛�)���Gǵt�eU���&�(]F��k�]���.�Bd6�5�.Τrg�z���!�p�OŜړ�.��| u�U�'�/�k�BOf�Q!dI`�aHe�{:��|�b6�Fc
��	���B��oA@��*�n}b���߉y���Q�˘��`��t�(=%ex,��{�����ٽIQ�ף�D����^d�]��b���U6}D�gP�E�����*��"�~���Q��:�}��g7o���Y{�P���թ�3krgk����Ptv���,t�m��Oflz[EIt�}��|�M�E|�6��@�������hu`QN����핡ﾧP8�f�ѓ�/Gg��Pq�{��c!{Y�z5k3%�7��K\�w�uY%�>�YG/�Ik�^~2] �a~���o�{s����� ­�Q��},b�Rᨆ��~�"w�
̧'ڳ���Wǻ:�=HE��p%>1�M�V�r���}tz��ԨB����]a�L�����T5w�&fo�D��ݷ>ͫ�)`��]_u���:�k��uф����U��G��XZ����0a�Dv�ͩ�9�k˷a��B���J�簍�mې_��GtP�|�uG��Tt��>����C �	�
g
d��&�>�����?Q��C����n`ȇ�ezy����:�����f��p��~�� �Z�>�K����2���%r�g��Їlx����ʺXWNҸ﹪�X��,Y�s�0�ᆽ�k���~u��;�����V��4��n����)�6�F���Om 	�� ��j��gQב���#m�	������K2��ͪ��aLP$R�P���	�z����N׷Y�髂Q�m3	�e�k5L.�ڧ68	�P�\DE*6�8�8��Oq��� F�ۯ����c��=��}]��m�a⌰�r�'�Ӿ�i*�z)����ޥH7#Ν�?vw�R1N�Dr�H����U@�{�@���I�gF��~�ooUb����je˙6)�kq�f F�@!{��R&�RW$�D��;Oo�������*���-�F���J����T�z�oV�U���/VE3�Ω�~������$6"��K���ʏu$*�<�%�?�گ��Ԃ��n���-�N�T;v�g�Q��(&ٔ�;aJ�.æ�0~~����2�C�r�N�W��#�6�����בӗ�.������U��p��ؒW��R�����O���;�iW�<�C�6s���j��Z��(;��r��oU:B�1
h�-�����:�	���G��	5�2_t���+a��ϟc�G�� ���g����k��}��Q.5�����M��)�����Wå	�UR������GU�B�i����uRݣ�	SR��E�}R=H�Yۥ��Z� �/,��Z]
�f�ԍ���}~������v����/$�'h]%������Z�� b:��ǤU������j�ѥSt��O[:�X��N���b�Ye��4�
b�%�&��^���m�(݀#�!�hkOn}Vٷ3\6nH�T�i�L����uj����}j#nz��]/=���'ҫ�㫈���A\ևx����v ��`����i���Y.�x��#gie���>�q��Cs_�&wk�B-� ��Ge�u��C�H�믕!�i����dC�r�{*����/}�}j�A��i���(��%j�Y�S��Q�7�L�̒��X��m�>���]V=��D�`$s��|N�z�k>��6�M�(�-�2����r� ͺ��t��mnc����i�N�(��j��u��{7�V]�y�'��8�A��v�3�����ȟ����%�O��Iw&�ċ��	H3
l]ZQu@�3�����',��rܜf9h>׶� ��u���ٞ�tҪ��A�wT�}�)b)������;��W��<�IVT.���m��m���w�0;;����\ٻo}l��h�����;���+�ߵw��F�yx�����Qg|	yn��nuR�WC�Q஻��� S<܅)�:o2�#{5�!]�uǦ���˪���:W�<{،�̒즱7ʡ����V����ΥH>�M�������U�U6��v6�m���	�Tt��B�̾���U "�:��{�����C2�=���R���e8���G^���w
�;�At$6��kl�1�d���T���_P�:#S��"UJ�'�=�ҵ����ۖ�gCjbM܋���{u�j ]ݵ_�"#��y��DZخ@a�������*�EVz۞��Ш��g^���g��3��Yǝ-�ŎJ-�7U�P��y���9��&>W�U�*޽�􏛻���;ٵ_�DA���8�S�t�e<3�<��G>W\��3z��^yg�҈�Ϊ3��ri��2K���$�ݾ�r��ް��U�?R���h`;����s�B��2�O�pC�|�08z; V�Fn��r>�[�#NF�PFj�z�I�ۓ����	9��P|��]W�D^O(�%���e�0��4�A�2˗}Ҫ��y�W�������uHVԵ�l����l�<�.a��[���M��H&��[Q^��f�#�40@���!h�	a��췼����q��|EƸ>�t�۝�>o��o����(�x�O;Z^(3�K��~�w���o�p�s�|=F���}ny���m������|6�����z�?E��p$
�&�9M�Z���*�'�6Q�0�mnӥ��� =�n� 3s�V���޷�ymO�#!�c̽(�nR�#�)7��W[��!�#_w&�M����?���I��U��t�{�N����;�(b�-�FS7%�UTA���;�:љKH�κT��ԩ�vyw��&�);<�kmL�K�|��R�����d���ߏ]wuHB;����Sd�m72ܔr��A�?]
L2����	9۴(�*6G�{�o=TO_uWǙ�\(�؊I�=�B�)�v5j��}�T�}�T��M��F,'ٞS�ތ�w7S�ʢ�C)i�zL�HY<�s#}�\�	��wf!��
�<je�S���%̺;B�HCl_���,q%����2�@�n����lq�t�&�:ݞBv�K��Ş���=�9������ ��"��w+���y�0ծ�&�{ vLk��L�PU̚���e�����8��E�K7��7�m�'���֧�p�.�:��\\<��ݪ�����nkOXs�6灕��@5�L�PI"Jo���j|c����U|	GvmP�=�CG�v�rv�ߪ�
$�����=���i�c�e5�y|k�z�m﷫U��m}K�40.M���N��Օ�2�i�t��Fr� >"���#��^U����T��M��򅍵2I.��강w���yP*��T n�>޺N3�s�`�uDs3.���[�%�ǯ��C̘/��Vޚ��F�Q�[�uF�����w���
mݸV�vևf��d���e�ƀ8���~�{iX���dn�/���8A���<���I�P�������1��1q�c����FX�Y\s��;�1����5�vv/*!o��������9�.z���Cxp+(ݚ�.�C��RՆ��dH���#y����W�n��]�}[�F}�yki�َX)g�oo���$������f��[���A-�qW�s{*ŭ��q��e��Q'��{����Y+�A%�̻���$��jy�}��g I})�*$�>�FIe�%�]�wv�H����̨I���*I$��n]I=���{�
����^v6զu�C��@��L\����b3�sLnu��#�q���g*����	fnU�A$���	�����n�Ea$A{s.�.m�e$F�|�{��w�g;���o���I ��$�Ks�
D�غo}��TW=����-˖��D�H�m})|�J}��������m��qc��7��pT���U3{����V���Sٗ��`���GtR�ChFq���G�6��wsI��������X�Z9u`6s�f��{�ٹA�YE�:D�B�K2&ɖ�z�#}K�c,�۽H�W��)� �&#+/v���k.c���n�@��	K�{l}��5�������˽�������7�"��d�XV/����3h�T�U:�C=�U`ǟ��\��.�?�Ĕ	ٟ�To�Z��y�Wc��!}�O�<�&��wo��_cr�R�����y��e�`C^�=40����ң��>�~��cp5�6�q��Ls�ɑ��]X���ۍ��i~瞧�n��[�y͡��mܱp��ȯ���2`5�+C��f[ݳ�[/ۏ�ҕ�؊�[���VL�X9�I�8J���j��������=�
y��ۛ3r��G�-ֽܼ�|��=��f��7w؅�X����&u۵�U�0��۽�.�4������`ϲ�U�{�`�u�Y�øv�-�J+5� ~��t��^�3|��+sW��/�@��.�(q!����\`����gU�����͠�_���4J��n��0�~�ޮ0f�Q�E��1�jQ�k��8�+��Q�.�j�?<�.�������He��*a0� �GVFص""�0���,P0��X�0�TS�b��a1J����\\2(�(
��DIS�\�H�C�``(a!X�p�\5
�6��\&#i+X
�J�Ԯ�+��J�pщhT���BT0��j);�s�!R�����a�A`�� ��"�������b�Lb��J�Š�8�)sb�d���EY"̠6�U�P(��LZe`�[T���H��(1j�DfIY���"e�YYb��*3j�XTm(�V�Ha�$Rڈ!Z�)R�`���l��a.(�++%jG+��YF�m%T�`,AE&��2��X�I�%E$g�ޮ�O���]��'�s��*��6�M(�ɓ�+�h$�]�uv�H��s�I��P�u���8�������06Zn]vOJ$��r�]�����6J�$�p����@2~��%��מC���i���I���L�%%cm��sl���Z�33bF�I�<��FYro/m]ݤIywS�IB��"s���'�TxZ����I.}��)�Z`���P]�����B�y�9w�wWi �Iy�*��W�⠑9T���G����𒴲�()"6J[��R^�r�%%^���}'���G�9U"�I�t����Ӂ'�p��X�n$A.U�$�C���K;��vk��P����3�,㤎;��b�M>K/1s�7�|Y�~ݢf�E���u�pZ�5����tw;�j�X��ۖ���J?j�HWّsi�ڎ\+O".I����?����`�zI����$��t����ʻ]X�q��i!���.�.b:�<Svy�m�6��%�	u��]��t���~�`L4ܺ'�E	仕�i�Y��V�}-Ă�\��_$���W� �;x�q��K;ҫ��S�f�����$Nb��$�;���A.8T�6�EP6 �8,�)04�K�;*�� ����W����N_�xI$�˷��Z�ie6R2Dh����0��s���I�,�I$�׽��O�<�Naӂ*�p��/�;�M\�4�-�AR\�'w{�I"ifӭͥ��^d��R&�I-�n��D�K9P��e��dZ�Y�qn�Dm�x���P��kI��t����Ӥs�^��	�"�\��т�f�JS^U�B�ST�_0���st���ۤ�v�g�n�[������U��fI���8�,�X˙[a�=�A�P�<r;S&��&ءq��f��e� -�t��m
Z��9Ym�A�uA���A`�:��N��	0�kq�|����S�!�l]a.��Ymb���=vu'-م�]��lSV�)Ԇ�x�B��WC!Q� 2EC�p=eڎ\��ꦉA-�ݿ�I%O9U���u�^���R&�Iw�w��yw�X��7*�-�FPJ�L��o��X�l��I|��f��AVN4)�>�٨�w.c'/R.1A�v��~���&��,����V�9L��H}��v��
 ��+�Q��kU?R>B�g���>I��_��I$+����V��֫f;^����Lu�"d�%��F�dPA<:'��|o�P;����	9�����䯕�_%â���w$�0�
(1hCA�E�k�Ǝ��Z5"��:a�������>2�N5|��r���U�iR	 ����*	�t6e��޿}�PI*٦�*+�F�M�%B���A.�Q��wKOp{zc�hl�������[��1��3y��o��n��ʼ�ϳ	���'=UJ�v.~w�]]����)`�S�Y��H�_�xH~��$�u#�N�;?_t��������U���$��W)��	XB���>���$kR)$/�Ҡ�
��-��]޿{�A~��	��*A"P�wJ�I$����|<v}�ZGyх��0��庪�4I9�� ���B
Ͻu"j�	�I9���3w�����ڳ��Մ��P"FʑX�$�j��\���o_<|���+23
M(َ.���
l�����R�I,9q��$[��w���.�W�ܕ�yJ�"�^[t�%Ӱ��'Ir�{]���H%og���Jf�&�e�% ����I%����Y$�=�tc}�)�)/�x��$�rK���T"I ���o�D��-o)u���9��z�Zvp�'��t�|&ܩ�ǽ<����d
]\G�!���˽1��b�Ɲy����8�<�����G�{o�K��k�%@�r���UԲe�Ȝ���"�Iq�*"RKs7}�I�V��dx׉(�G_$���'#��]{~���	/���N�����,Nl��<1W��M|���wpG�:)T��Fmi&��aN;^�'	Jd �헋I��kk(씎���}_o���+���S$�K7{n�$�yʩ%U��sF/k�Yt�"N��o�%p��
l����ߞ�5����T�'�OĞ������$��T�H�#]b���ѳ�*�'!Ir������D��R�IǏ|�מ�$�Y���yJ�r�J��<r4�nIp��'<�I%�����$�B��	$����=�f�����- ��7���:u:��Wx��V��+��~�A|�P������m��$����{�}��b���n]�O:A$	��'�i�%M��)jh����m�V�$��wJ�^��_]\^}�dc��eF8ƱɄ������;W�Qq���>~~�yXr_.��{�y$��^��I$��wJ����:r��=�����%}4�$&������೜�G^��L�j6�ov_y �	g�I��~�A$���7+���<=��&�A�M�]@$�Y�҃H$L���Y�_\ʭ��'��E|��~�O1�d)I*J��ŝ��ъ�k�ΝR���������o�=Y&3���׆_G�F�m�._�E�_4�I+�ݿytǷ3}��殼��$����I��E�����{�m�E��j�Z.�����_/����O�� ��/h�ե�[���ñ�/�:�;힇
pk�Xv>*/�|~��-�����U�`�y���#������a�����v��CM�Ov'�jz�x��=��B=�㶼��e�k�:�<V�d�Of9ݰMآ^{@�sz���-�.�s��6I�ݝ{rޭ��쁠k��s��>��T۰�)�y�uڜX�(h[X����)��j�u�H�Q��<��W�͆���0׶c�,��q�E(ZӇ���>��K�rMʢ^��R�"sW�4�	{7���]��@����H����+��~�MFf��&Ò�*޿{�I.����+Wr��"Vc�*I��{o�E%�yW�7��aϫ�Q��l@dpY�R`i���۲O��k���4$�X��d�_���Y��*[l�$�ݥ�ua����iQ�&�^�v��I$qg'��>�}:i�$�.�tC �
RB
����Ww��$���[��w�$)_S$���˲t$q_*���x[��גe��ر#�Z��-�1q�l.� 5s���u;|����ӕt�NP̪��K{7o��$��|����;{�^�d�I{{w�}ٚ�P$ܹiMte%�v�M��+���:*�����n���-K��z|���+-������ʡ��.��}.��I�$��+����$�[�_R).���ýB�w�����n����JC޲۔��9�m�2�H$y��׼��G�{o�E$�U��}JcT�@[�	kU^���)���{��I%�����($�d�TA$-u��Q4F�2X]=��yT��ȓ	"4J�ة|�K\e��Xt��4�����{�I[8�"�IZ�A*��q[��6r�*�Q�Si���`a���7[Hℿ9�!����h��*L��̾D���A"l��In�����|/.��z���o��$k��^<�9i��
��D��n�����r@�/����+�]t�$�L����n�,��	pMʖ�ta4��B$�3�ɶ���Jq,7�e�;۱�z�������+���~�3ʕ}52��S<n��������Q#۴Y} �{8�ԉ*�]:IF){>n(Sa�g���n;K��4�Me�M%�n:�$��n�o��o<�������I/:�	�P]o�#PY�2I>��_)K:���4`���K�yU$�Cˮ��Iwoo��$�P��E��a	�������u���Bƺ�k[nl�Pfy��a#$G9"��RI���$�[����қ��s Kێ�"�B�]:I��(Dd�%��9�����%/��?x�]JI$���A$����� ������X���;7�2~�EGږ��1˖��L�I%ݛ��<�I,���״�\��$�,�t�I-�����3d%�\	7*ZGj��b��x�I&{#,�-��II$������� �v���s&Lrh��d��wF�Ԏ�~���~�*�m`�&�!��}�r��˲s��y/Td�b����
lI,�]����&��V0�U�%C1$5UӠI%ݝ���+��Vs�7�z�W����c��>��K�+A���Pq��å�\m�ۣ=74�B�š�E��n3|��S4A/gv߼�I$k9�	!�u~<^�t�'�7o��URU���FH��E�9A&{�K��3�,D�I-�����I"k9�I�3���Vg���$:h�l�$�';���A$��N�	 �[pY��b�d�I.����'�*y���c���1��As���k�E�ā��K��p��yU$�K�]t���_N���I��{�\}�!��NS'E=�H%��2�]�u�V"|�/Jλ�D��x`���lR��~g�~A��
�e+PU"���i$� ŧ�����O��HRy	 H�f���͇?�0h21��;�3�.�����2MlϢz�%��Ɔ7]&���i�I	!� ��vX@�.�XO�����7�
�ܯ����d���	�fI@'�$_���ߩ�:�g�8�C�>��z�(���4h>̈b}��J�!���Өu�������&��/Ru�р��u��C���	 ��C������������H�t�$�2u	H���XY0~��Y�a����?�a?2�R�����!�}�����>A���?y$� ����h}a�	<̆a��!�Hh��L��S���H>�Қ0����-�&7$C_W��H|�~��>��@����O�,$� :>Z,�$�w�nM�۞�L@��?�`H$0��2I�9U w�Y���৬��k�?�}L������?���RI@'�M�lb������@����3_ �3����.���,��d��5�}'��������� _�2�޾�������� B@&�Y�>��2#g�C�}����0l�S���)�{�P�!��y_��� �1tO��	��}��v��c�I�M����y����?I@'��{�?�"~���Ɖ��h;�������e��I$��D��$	 ���O��M܄�[����'�%��w�A;5
#@Ćϖ!!	 ���� �A'�b`~t��vO�^�$X2h�h� �Y����>�=��x�I@@���B{�D�$�ܳ�@B8!��h���/�w��rI@'�����O��!�H}���G ��$��$���~��?��?��|��̞����p���!����P}r|�����!?G��L?��Bc���!��������@�	����k�}�_�BҐ�����p��K&C_x=L������������I�!�>`L"��u����C�1�ߍ21�L?u�|�~��?g����C���/�~??�w�tOC?A�g���$	 ����an�Ᏻ�#��_ӽ;�tO�<��'�qa���:��~�����&�Ð��	 ���?��� `����	���?���~���H���O��H$�2�~��I�֣��������׌h܇�!��?�Iˇ�	Ϥ��.�p� �aZ�