BZh91AY&SY�f�h�_�pyc����߰����  a3~�8   *�`h   �  ք;e   ;�                    ��l
�TE��
)ǀ}�f��H� �}�B����R��n�=�{��Km��=�������^=g��z7��}��>z�+op�Y��{A�9=�s�W���_>������W٩����`s�\������/{z��̮��=���
�h    <Q=�ǽ�_����GM{���uO����=y�*z�U��{��۶��\Uއ�zr=�}�Fڗ���t_�s�"�f}�K�n�Ny��U8͗�v�s[�C�x;Ҽ��c�5�#9�ҧK@(h< z O�p>T��wW���N�:i	���t�l�w/a����{�=�����| 7��46k����%�l鵢�����
�����}�<�o��� y�P C�\;>
��㱟f_[ղ�o�%{�+��*�jU7nJ���R^�7�� ��ϡ�{�������<�(�c�#=�.-��Roc�j�k�O��|  
a�>��r�o�*W-�v�W���X��*�[s�<-��.�� > 
7|V��S�������Rdݲ�Bﾣ��m�eW���+�H        "P
EP    � ( J��47�T��4L!� dѓM��i�5O�	JT��i�  a42���JR�h�hɑ�������@	OD�%J��M0�Ѧ &�1 &�� P�&��ѩ�S�z��6��3E�R�щ�&C@``����������5w�s.�~��l��Ο�$����4� nH$A?�I @?P�����8PJ����@����GULs����ο�?���������#���BF"6Ar�* A,�~��%(J�I�P ?H�ȋ��_@0D� HA�)��Qy�"��u�	������?������gZ�z���}ɒrj��+H��1�L1Ô�B>�0�g���3�D@�@��~$ϧ�Ca�,6���LN��V��B'0N��%_֛M�r�Q�5F��Әu:��I�D��$h�m �gd���I6l�d�6M��a���h����$��4oF�Ci���Q3Z�h���/�eD���N�:�(~FMlI��D�D�Ҟ��"m�ԡ4`��7�֋�|��DGMV���D[��edJ#�L��y)��X�7r����J{)�;Sbj�N���:e}�u��C���H���?�"&�W~��֥|�r%D����G�MsR���ܔ?r�X��"pn"/%p�W#�H��+���DG�+d��#�D�R�.Ǳ(s����)ܤN?DEԬ6:䯟��D�u+b[�H����Q��_P7)�Nu��F?L6:쯟�V�~��u)�Y���>Ϛ��4ܤN?DEԬ6:䯟��D�u+b[�H�g�t��_WܹH�{)������5��#(ώ}�&�d��H'7�\d��T?"�R��̉�az�vN7r���<���J؝�UӅ��rXԳR%�K��rt��eh�t8Hl�A*~�J"�}��ʢ�3�2X��R,D��[�#�+z0�M�bN�Q7 �G�Ӱr&���656�Ǖ]d�r���N�8$��T��䓦��d�7"5&9"k"a�j��Ut��A�ԋ����tL��c�d�2C2C�#�~��fv+)��vWL�'~/���rG�����˒	��R~�?T���xѰg��KmIX���$�a�{R�䟼��%RE}�$<���=���뺮�Y&IsL��nw���i0�M�+�w�W�p]�V���)N|�w-�8꫙��ps�UWnNj���}5=���g����o���L	��^I
j�i�|x�cXk�j��R&�'�����0�7
%}�9���rN�,�	��6r��dލ�N`�LH)�&̢�+EN"r�u3	txS�j�`�p��='lzY}�����$���8��8��>j>��N�RLL�l�����.nz\�Ӥ��������m)�WZ)�����ײbaC�%Q���K:G�$�$�C����2Q��2sF��Λ�&p�2W0�Es��,4H��Ch'c'��+������B�MÈp��t6K4k��h��I�5���ʑ�#�2N��ϰH�?pI�<'��Hg����6e�P��H'z�,��=����`��"ȏ�3����kbw	��4'o	��l�'"s�=��'G��xC+rT�"j�&0�49��ΔD��	i6"sI:�YURBp.�"q�"lғF�6�')"p��DNm"#�3Dᡲ]�D��N�d���������%�t�6?q&ktN8M���V��%�Mꈉ�$L:�lNYBA85d���"WRX����|�t�����N�%Y�H�c����YN�P�O��DNL�J�'�R"t�d�&��O�6�:�~p�*��sI6��d3D�IӮ��'G���&��w�p�ĴK�I�h�����	��5è���N�+�'M:D��o��"�(��;���R%tO�
*��%�sBWLH7	ϡ�JK4sBu�,�^��R'pK14%|��d�5bq�&Η�t%d6�r��#c�N�"Z"s�YԲ}_�KD�И�`�K�f�/�N$�I�X��f�;��L+|�I�o��obxC�����8�q��t�ɳ���H�ݤ����>�l�:�Y,�;@����Rt�H��;�A"�0u�zP��Yf����G��H�|$,��9��#�%��'���HM$K+I;��a���N���Nu�|�4h~�DJDDI�Ȓ�&���$N�=�D��^\�����I\&	��DͤN�8&��6s�;�:h�'"M���4<�D�a��C�X�����(~��i9�H���l�T�������u���:A����l���N���Y��D^�ᣣ�l�5>AȔ&�L�DG�L8P��r��#�����j"e58l��O��TD��p�cȉC���)�O�I'Dy����;�,MI�ʦ���TO�.O	��D����
>NUTDuu6�7��SS���S��N�S�I�C�Ӝ,{u��nH_{R���$�?r`9>�	L���VH�]觓E�G%��0V�	܉�6t�7Q4<�lF�Q0�2tp������"wE�%�n�^�'D�ڕ��L�(ᾥ&�<*�~��t�٫����%5>�ϑʨ�&����b5¹���^�!�%�J�:Y�#��bX�v�uڔlM�b3�X��Q͜���٭�x��2'���l��ԇd'j=�zw�S׳A���ıު'7,w����<�C��'~�!�2	�_�������l���uj9[���7��3��F�2&F�i��QIAb�v�W��Q�[jW�1��Q��o��=��R���ڛ�Q��j)&���3���Rld���$��^y��G�K�|����dH����ީzP����7�{���A%a���������G��MO�Q���r�4��V=N��{�g�^�j0T����s���}���－�8�ՊsuwDrwqdd�T�(��>~�{U=ĸW���ˈ�!bG�BG����>揶#숱~�B�>/�>���D�"��Nf�5��n53}��}��sG~����CČ>�K㺑�:<hLM$��>,B~�>ee
�i���OuQ�9�~N�#ɏe,��}]ԮL0�d�؉��l���DM��:�f��W��%~��Q�%|�Ț�P��qnW��T�-�H�nR"ܮ*�${)}et����%l�0��4S�D��R#ؔ<�}�5)M�D��D]J�c�J���MwR�%������I�����nR&��D�2�h���]����٣O�n�"cr����3�R��7)��u+��+��J�X��R%���f�E|ܡOe"s]4c��|�Ϝ��eh�p�nIE2Dn%rRt��T?`�U��\�ɼ��t�L0�pn�Q��<���U'>�޵Vt�2�nK�jDjY�Drp�D��Sr�}вCd�	P~{U����Q4�}_g�)ܤ����)-��]5����Xo&�1&NQ�MnA��gȏ�9&Ƣp�ʮ���t:;�Rh{�����9#�L9��6�56nDjp܈���U\j�R8�;�B�0{UI�j#�d�� �>���ϧ{;�G�rn��λ�L�S	��t�-�tq�T�ԾXAex/T��O�'�+�>�"�$�J�x���Jڐ��=�^��bIT��`�}Rc�}��R��X����0�ϩ�v�q���	-O��R�7�����/���ٳ��77��<���T0������4?3���!�r1���U�������Id��|��"k?�d�ԏ�k3��_��H�����ΰ�fu�a�p�N%���%�f_�%�IjV����ћ���̺ޅ���Cu?��^�!>ZT2��2!�+K��8Z0�kx�儌u�-cY������4�v�N(���4�YZqR�Z�dt������g��ْ6����(�;�JH�t��2E
�A.�i�l9��QH����Ýι���[Ӑ2��ix넶d�F8��R^}E`Jf!����-<��_.3<��W'�v�e���:hH~��ko��j_��!��c��s������jS�p�>!��>�<߽�akf*\y�בy�S����+;�Ǣ�� �v�8���Rx�������M��-}o�-�Z�} ֟��<\�帏c^ɴ,��Z���zY��F|������ޛ|��u�Ӛ)�x�˹��}W�Qe�A��>��0\wu���zd4°%���SY6fi;�',��+\[6=�ZI8i%�!���#�5�4����f�\׳�Z���L䅘Y8�u��,,�N�Yf�Ř~Df\՞�gM3ѷ�&P�$�|Y��[��*�����j2��(��2�)$�Q������qd�ci��aEY%k;^,0��4c�	.����I'˪����ʅ�%�L5�x���:�ǰ�D�jwL��j�8��#8��2?fgg�X���5��_범h��y�g��nm�Sx��GV�m���:�����
�C�BNc�T����_�n0��fj+.+����yϧ��b���i#�2`���˞]����y���|����0S<K���O���C���3j*U��G�����׆)]�ܳŝ�2y��f�(�,O�N.J�ǚ<{}�˚&���b���RRNr���(�m��,�r�Ƙ\n_��:0�w4ܯQ�[�?3k+cן��5�Q�M�ř�fh#0�������'z�Jf�9`�|�7M���9������s��"u-YXE�,�{4���y^z!!B��5��6q�"r$�
),���]��	�c���ɜ�۲_��e����2Z"#������^ ����!���Ʋ(��n�����e�X��|��;�m����6��7��yv��ܢ�T2�QL��2�x+J�u�2���m�budL����\����������#����*�ڴe���^�{�(��{�w�n{~��#Z��������x��e?��{IG�G��]cfl���i]�,�C�	&��Q�~��I
ffsÉ�l#sl�VI����0��O���}�O�1��"-6mC�˪K�oȇ����P��6��5nҗ��g�B����Ȗ�p�������p=��.��X�7&G�lh�ή��`�.�b��Ȉƞ>�J{ٔ�������f�*SqZºWC�������,&�Ux�&���g��i$�}�l��L�LW%����������̧̳2��!�˫�w�w����͂�7�9@�s�Vf�C7������8�����wc�5Ϩ�PV:�]&�ɜ=q���7hgn���h����]?�2/��ґ�#>��]��d�v3��s쯳Fa�:���ׯ4cڷp���?3�#BBas����]�Fٷ��'QAO B_;�;)`�q���?)��wJwH�������s��/���81p�0��m���1���'� O����ݙ�ó۬2�O<+܋x��?G�p碓����t���u������3�~��\������b�����|��#��v�f��,�������[��	�H]l��K>�9�:Y(�j*̡;�;=�HlF#���a8�mDǋ��w)�K�����jH���^&�{�;"�q��{E0�NU�8B�v��gjUj�܇��E�s��fo��Ȼ�߹�9�w��zr�a<������ #L�\����+B%&�Y��X�I�pؽ�3�d�O1��kZ'�ml�8��|N�Ѿ���
eg�:L�ߟ����o���)��vu��z��5cC�>EH��[���̧�H����"g����fe$�*e?sK�H�����w[|�(P�܀ø��,����u���X���"�R�E���;�J��D�;����T��g��O0���o������dQ�kۆ�a�|��?P��@Ov��,� �7�Śg��QD���/�H���J���,$5��d���h���\֊�su'=�.���������YD��K���M0ݏ	9��FY��p�ձ�*e��=!�sd��=K�K�,f�99	�2qێ��oS���f{<s=�����j���B��#&b9i����6ƨ&�;�|�T��i�w����c1����������v��t{��޸���$�l���ֽ��L:�d�P�����Y�|�'��Nn��NS�̾�^�Z�e��'����_q��g�Ռ硫��qn����O���+���ٯ���٦j�1�G�sO��7lw��`������g�G�H�g/�Rv��-o{��D�Ml�\��x�&���*�e��\/�f��#ټ�x�ěHSt��L�x'0����X���c�}����?w�)̑���Z�l��KD.c�6l	�Y^~z9�0�p���ڤ��<�.b�/�6$w�>�Ɲ��z�o�ܥ?k��r��=r��^=y�3�[L�pfd$�|N��g`��g���V|]NkQ!����p�+^��3��+��'4���b����%Cݒ���%f��Z������dgq�s��g	'uDS�N����������]���=�Lٯu��)�1�e�j�^qV�fb�{<���W�ԝ��������0�������=�F�R�-kܧ{���:�^K�!�~�2�z=�R��p�}�f^��+�������|���70����`���S��^؈�$�����:�|f'���z<����⬽>�ǟ�QI���7��6���H\}���:t�N*R��.l2BJ�%$�E�,�'��ܫ4�ٻ�Go�/�����U/�/��6�B_k�/�e����7H��2����r&�r�><���{��F�~naGt���G|.W1G���?Qbm	���ux%j��l�G.u��q�4����:���p$-�	'q5Ǯ�7��tӦs�^�#xF��/g��34����[���dz��6F'i�Q2�M��:'�7���������k��8���k��]i�;�bv�Q��^�[��IX|���l&P�o�s5��O����Pe��8[��E��G/p�F�'�>��W���W��s+U���>aӁ�N�+1L�9��˻�f����r���T.-[#��ŗ/Z�W����������1��v{p���E&��[j�XJG�7�=��E|��zmm�TiELrK0��:��Ӵ��³j.Qݍmy�	�����.�^|sK.I�?���0��������nW�N�f�V�w>�okվ�p�3�L�:7�3���#n��D�y����w��p������y�V0G�J��6N*a���j��]�V�:s��7'^��~&띊S��#���x�,���lB��oU�:�Tu�g^"{�9�3��œL��Fbs:p4vV��HW�yoz���p�yxʵ�� ���N?I��ٍ�ɷ�k�m�������<�姰�ۥ��}�X�f����D���Y!?O��=����?����~�ax���В�� ��������X��Z},�Go�;�>&�ԣm��@��X嚐v3hXE��Xq��m��A�K�k��V��J����92�hG>��cQ��Y��fP<�n[M}LV�[�<��ݭ�A��l���XKM4p\���b��rb>�+MD��׮���Q2Y�ӫN\/&��ók	�I���iQ�5��m���2s��ɛ̄P����#J4D�f)d�p��,8���-���wN����]�f�R��^[r�m �O���-�'��SDθ�~zwK:ذm�|���d�a~�oSWM��L*��a.�=2���ﭔ7p{3�4�s,��}��ul��#N@�%���?ߞ�B�oK�}�݊ۈ��/����j,�'&2�D�$���ٚOR�����PF�rU�t��Dc�r��?l�~=��{��L�cb�(?�����Ɍ$��6�0���}���t��"B>����8a���pA�6�В��Bmu΅�ս��Ͼ����Hy�"L钴x����~�:}ر��2���X�l
Vo>�Lu,e�j�o��Ǿ,;�+m϶�u}�İ��٦���}}�&|����Mn��j�)v�,I��XiT���~���%!�i�fk������-sA���L�3��}�E�YV&�-�Cil��v�tD�E*CA��&���ЊѦ<������E��mɵ��_�wK��)hŖ�F�,��H�]R�q��H���x����Ѻ���3S߷�{'Q�O��<�<�V�h�I'�rM��=!�1��cH	 �{]�~*0��}4�K�}��ġ^�>����̃u�r�i����a�SG�j� ����"ɢ�,�8����0����+$m�" /�Ah�w�u@�~駽j>�/-TjSr�Z���r"����y�W�QhkR�+�U�u��9�qe�L��ev�M��#�B�����Tp�H1#���6�&`�
�D�����}��B�����/���L�H������q�m��A
Ȳ�i��aO��g]tQ:�,���f��Ԍq�%і��2�l�3�vn�GymB��#���g�����'���s_R�i�nv���1~��C���1��(T��Щ��e�'ERî�"E��$�E��i�	�̰�C�éY�xJb
ٲ�@e�pa3���VcO�˒����Q-���a�	3(�F�6mye4�I;�~L�<.TM��m��q�\-��P��*t����3��|��!_��*�����^��1��$d=>A�(�џ ʩ2aJ�YA�� �d�6HI}>Ǌ�u����k��1����~�~���TD ��o��'�S�ب���nJ!Q��74���������!#� �wJ\��'����_������%z���ҫ����[Uv��U⴪�QUU�*��*��t��U��U\X��]"���UW��WJ��]*�*���U\X�����եU�Ҫ�WJ���V�U�+UJ����UU�UUTUUTU]|����I! ���idT�lB�R&��H*B
��P�.A�R-���Z�**"�`��>��>	��Ez�s���*���U^�*��t���*��]�UU�UUTUU�Ҫ�V�[Uv�*��iU^���1���WJ��[UmUڮ�W��U^,UU�UU�Ҫ��UW��J���X��UWJ��V�]��Ux�*��iW}�p�Bԕ�-��[D����J��A�j�vI��%Y$Td$b@D	@R$P	��IAY��QRAKWw4��V�U�*��*���UW��Ү�W�U�Uv�*��UU�Ҫ�V�Wj���U⴪�QUU�*��i�^+�Uڭ���mWJ��iU^�������U]�ڴ��K�Uڭ���t��ҫj��[t��ğuZ�C��I%K$�R*��EX�R؋RKdZ�QUh�ib-��h� }�wޯs��j��ګ�iU^�J��b��"���U]�ڪ�WJ���X��\N*��Uz���ҫj�եUz�UWUU�*���V����]�ګj��[Uv�*��UU�Ү��uiUU�*���UW��եU���'���(c�a��*.��&��H[h�H�Õ�Rj�
�P�5�$��`��(�Pwc��CŚ�%XN�VH[h�Y�srE��BѪj�X�H%�J�J"��*(�PI
������P��P����_������ �~O�~d?aG�?i�����&��8x�6t�""pDLI�"%���&�lN���!�A ����ѡ�Љ��t�&0L:"`�&	�4`�!Ӆ�"`��t�DM"'A0�4AH"%�:&��e��p��&	��AB"pL0�B���gD�fĳbl� ��pD��tL�"&�$0�Bl��>J ���1&� ��"&�N��"`�6&�
AA!��>7����3���6�Z�Sm�F���\�u.j]ub�c��A&��5��)��d���{��KoL��ccro�u��y���E�E?J	��ʰ�}R�j���lE�m��5���Ni,�\fm&�@5�X��4ve�Q�j�ö앾 V�G7�t��P�������]E}�ڋ-&%��,)�D���ڷM���!��Rk��&lι�"̉$��*��[��`������6fG2����N,in�]�B�]�aD��wj������
�i�����|1w��^��hiLX)����9����z��ͬukB��e��XK�wgB�v�d�j���z�N�ĉ �#� >"׍�/'�Ս3��f�h&F41FY�!���t��u|���3����й�E0B\Kl�Ѝ����`�΍� 07Ts��bH�V-l$�邆�b�Xgǧ���YY��^�tĮ���Ѕ9�������Bis���GF���Wa�Ĩ�.+�e7wVq����S=4��n�0�v����&�5��6F�����{[�Z�SJ���J@���[n�l�F���0	Fe@Qp�%�F�a���B���qY�㟞QUU�*�wv�����X���U\b�wwo���努�UU�*�wv�����b���UUq���ݾ>>���ǈ�6��ᶘ�8����ݾt�����O:;/�Ä�v$���(B�7l��ř��3�z�wM�k���&n@���|ґ���a5e��iEN2s���-�'xT���V��ee�Kպ7����[
3H|��k-��&�Iw:ޚ��o8��^,�Ԍ���b��[l[kjBQI-��?��i�|����#�b3�8Qn��_.��e�H�́m��3f���NfHIF����R�^E�����1|�G&�:^��d{��S��sq=����6}j�(��4��.ٚ�Ȋ�Wߞ�_O������}$4�ύrh��'3��Q4[�������lm�8m�4��;|۱6Y
D�z�������I ~�k2���}d��Zut�]�{G\�M)��*�QG��N��ݯ�>pHu�]�jکP��d�v�-#�q�zw�xf�믧��Xl/�u��u��/1���#l�n��i��2A�g�w�����jD�xo��BU�3��<��Jh�L|R[��}��7�Gޫ�m�lp�O|K!�(��,�	��Um��WsSP��l��5.�컼�M⪮<3�w[�n]<�E�ۣ��[��L��#�BN�{)ӕ9ㇸM)ã�_+`�5���T��,!,M&�����M�s�.wp�\���>mpN�*sy����0�*�G)��
p�v����RnM���3�>�4sp�
gf�÷�UK���P1��9Ԓ�f8c���p�Y�f��(K!�(���D��:=97�*���[�I⪩I��dɷA�L9,x�s�+iG�4w����O�@�WM�~-�_���HD���d�4���9���x@>8|�pHD��Ըmˣ�t�y>���?>m<�~,�PA��_C��H�I"������	��7.p��c#2a�Vm:Έa�|t�]6�8v��M�p�Lh�b$8%e��4o�N^h�g(!`IX���H1�Lla���X��}K���
��N����s�I�2+_���鹖4LGj�����"ye��o����|�� 
�Y]�Jk��S�a��%:۫r3��V��`� ��J>|���+�}UT�7��*�Yb�vJ���6�
��}���g���}IrN���F�����,H��(4�KI�_����ty1N�j��� nj̛1��q��R�T%U_�R�i�9��c��;��w��X���������$�ߧ��;�G�b�Q�����cf�yl!`���=<�{���MβN�X��(CD��OJzhR�����		��P��eS�r���.����7]}UT��ON�y���f�0r����hCp�sBC�J�M%�n�UQ6w�.](S	���t�(4Z�$!����ݏ��n�t��.�#�,�Ҷk��$���8SOO����.��G��F�{�_�-�QO<=�.���� �'�(��#��8nyr�uQcӣgN+�z۷�����h8&�!Bh���w\*�gI�z��t�����$3/�{I!{4l�n�t-LL'Z-8��3B�tns	⸟�����<	�w��e��ml ���ns�q��۶�M*HI �&L���u�\P����x&��b#l�E�S�3��� �TS������.\�f^ܙ+�x�L�l��s�	
6Y[�-ѹӍ��8���ᶞ���8&��l�&����[��!˩����J��d�US�Ɇ�z�׍�r�ܝ��p���F�d���^Abxyv�a�R�% �H$�5�a[_�	�5�G�3�ϳ���V��l��BB#�2��]l��;�Xք2��p���<� jLv|S+;M�d�ξ'>M���p��Il��(p�N
2���M�J^|W�h�	�BhK%	��N	�0xQx1�a��ġ�J��X�l{5�8�D�V����&^�����"l8Al�T�@�s4��Oq/���f��u
���3q�Ra��t]�wD�o-�V��-&�UU+�U.I�Μm��bw���O4�R`zb�C��B�j��D�Vޘ#�c��ቺm��+eQR�(x�(˝�
"u�7)�#�q����"�s<ΰ����Tɖ��1���z�I�;1U]r�f��9��M
y:��Z�d�!5�օp�\�;i������g���i�h�Nq�5*��@dY�I��D6Y�	a��(D��h8zp�!�Gθ(簝�,����uHv�j#���o$F���b���B��̸C��C����;&wsG�GgE�쑂1��ӯ\\����&��Y�4i-�D�$�Ɇ�4s�\�L�Ɲu��S��˻5׬���,0m[�^��/6�k\l�Yf�3���>��Y�M~���6�;�i�ifJr��҉%U8���fu�$�	�����E腖|���M1zWJ���k��[��\7�{V6�..3W�7����\j�..6�3W�b��[��q��"�|�|o�v'����)�*�����j岿/�~V��~^,��M/�~W��?4�����'�t�F	^'�	G��<J<% ��Q�	<D��IEa���&ɶ5����^���V.../�.6�/�ƚ���xƜ]+ի�����c��.>k���x������.=k��յ��l�ƱzcX��5���v�-Ʊt����������~^�5�ڱ{V;k���1�Q���m�q}\W�ճ�4�s-�Ř�1�+�m�L�gUH4U~D~U)>����|1�^����\j��\m�f�5����������V�ƻWJݸ�f��t֙�{i���²[r�^��,��Bs����rc=�k{/~��k��~�Yc۹���^KH��a$<[��վ�*^;���c�M��m$���f���=E��jC"��U�s'�^ٿ)��~��f������]oz�����rI����֜ə�<�d����4�ܫ����W<���s�������̛���dǫ8+��;���T�|�T	�����>�|yUW��kO���>̙�����������kO��3+333�����*����>>>32�33��{����yE]kZ||}�C4a�aG�"pM��8l�x�k{%Wl�٣����@�vbC<���;�>4�f�8���j�bIK���D[l����s�0��49w��6r24S��O��Bh��?&�J"S�JO$2���Z|�����=�X_��*҈�[�<Y�4�@�3��&�JD �u��Ix&�g0�L�a�
ci3BC⃤@�Cq(���D�ٳlGKI}d��#���.I��Q��q���"=uZN2H�nWty�x@����D9��h����^�Q�!��>�d	(���`�@���X�Xa"�{�V�,8�ԧ��۶�8m��1��6`���d4h��y����+�X-��������ڂH$�H�H�>x��a]#M�K,:�y�BI!)vS,N����#�Y����j#RF;��ջ$�K!28��4@��P����rR��@�I(~Hz=���a�7vq!g&!*��2bs�Iia�	�-'0�l��!!G�e"�dD^�J\0�����N$2�J=���2 ^���Oo
���7���	�wє��KN�o��k�����[��}���Z���.Āp�l��IJK;I�=SK!��j��o�|ᶞ���X��4��ѣ����Ekzwe���@�ۚ��L����+�M�w2Aط1�r����!W	"w2!�d��l��K�)l11>		ddk�1�q���f*P,�Y��!�K�2d"B~�!�Z*%��e��li0�e3��o���:�i컦���i[��GSOy	!$$�.��mX^��ťhWZ���q�0tsy*��[̔D���)�Z F+
̐�ʹRQ�
{	ORw5�፦)z=��£J���D��R���$C?IN!��)JH��\�8�5�q�b[�"Pu�R��؛S���U��֭ѩaT�,^�S��;WU~L�DN��a���4���MC�g��2V�U�Ģ�#­�sr�nZ���]H�Hѱn�p�8L��g�xLˇ� ��BL�2�'��I��q[��>Sf�W��޸m��>b�N	���<l�F��Gz�'�r�UwDd1 �@$%���a<za�۲��-�$0L���>��~���� �|!�p9�o�;ì����=*U7�اNK"�nKnB�8�N)�ZEwK���:���C��I�/
�A�)�-�2�M.��+�VC)��Ry<�広Q_4��!�G����j���6�T��M��D�))!�)���"09�	JD�H쁖#'a�=Yt�n����v���<��1B�+L^,>�خRc�<�ݑ����V�ֶy�ܲU����ܩ�S�n+�ߛc��~(��X��4e�(��G~�v�ֵ�)m8rq��BHI	 A���oiJY�C,>H�M��bFh��T��;���9S�ZC���p���)����f�KW��r,+��5�ʍ	���{|R��P��jx�gb>z��U�Jn�Œ봓e3��b]6��B]����hw���H4�SD2��� Pq�P���v�E�=K]�h"p�4A7772J��oH|r�:J���;�g%˦wE�r|D6D�#bDz@Ǩ<����ٺ8���I�!�;R��`Ӳ��	���g"��n7a�g�c����O���W�����p�O���>v�C�ӆ���&fk�l2�6\
���F�܃ n�.�+&��hbA?K+W�soȍ v�`jj	 �
@���A3<5:d`��<ɜģ)N����쐒�8�R"���2$m4@���3WP�!,+9��حf��c��n��f�0@���';��d�=�����%Iur��.�HH�v�'(��>0�L��4Rp�IAD���s�o$*�v�l�xu�L��üp6@�� Vt����M��6+��Q#��z��*cfP���%1x�$@��eܓq��]�&Bg+�Ow�O�?HB����@�4�;b����$�RtjGƝ��m�6�ᶟ�|������ON|B����I}e�eTqz����Q�髳��\�Ilx򡌹"�m`�y���(�$n�Ք��:�V�������j�J�*�I��+P�\���3i����e &���X�U�1v�>� �HK&�߾�e�X�_rv����u#�]]�8=`��)nI)�C�gb#�~f��X@��u��Xݞ�Sm�(�q��:�j֡�P�OS*�BO<D�LJ�,>Ht۬�-:J� �)�0��⏘6ϡ쐚-�>H�HV
{���%��h��gnT6Q�0D��	rHB{��v@������H>��Md�qڱ���Y������H߄:�7��$a#	I,J�U�;�n�@��N���4-��djy�}�j־����nr�c�N�u��N~�x/n܄rح��q�.<����F�S��޶�Xh�(�?8&�	F�<Qg��wyʑ"p��y �b��w�G���I	!$ �{�[�p��EH�	�������Km-Id� s&u�γ��)���y�>����3�����������:�0f���oI��m4�)�,�D��>a<��d<Ra�?p�LNQk+[<����Y�ܱB!���f[	-�f��6��t����k������<?�Mϰ��e��0�+�l�ˌnH�.�I�HnT�)��i���
K{���F���b�����D�dî/R&�3✥��&Hh�gŜ,4P�~���G�e�(��>��km���8�QӒ �HKc��֛Hq.�������I�ɂ�%���0��o5��f$$&0�oZ���a1���%�,�ΐ�����2y<�0�Q��!3�e<nʋ�%��24u��i����$HK���f	��w��i)<�����JN��p��~8�K�A���>�v��.'0 t���{!0�x���wNʠ���z��%�Z2i(۔��a����H#�2J�f�2��yD���x�\'����!UUM;4��A0�B�-�-��u�K�a�=T���c�ݶ�ᶟ4�����G�:=!�D���O	!�ϟX�$�M��UO���ρTj7i�p']l�͖�NkE^���f��XI	!$ '�ɗ4��L]�:�1E��tc��IKkF2�	�%�SB�N�CD��W����q��lwaf�,�hW�Z��j�
(�%�!q���o�^�|L Wg�|k��l�̝L�Ía�_��L)��:�a���ɩ"I�����z�0a��8��`���R���J6a:���D
ĥ�-2a��d���@o��х��ϊ��US&S�%`��|ѸL��������;5Ѣ��ۍ���2QO�,��C�:|C��G�<!���ω��G�b��=k�:��X��b�me��/lkj�_�51�N���{^.-W
�m�m��XV-\_Zi�1Z^+��8�b�	d��(�����!�<Q��>m�>i��c显�4��./�Z����x�+�ƿ/lk׋�5W�k�4���qf��/���qz]/��5��MN+��5��X�1�h����c��]�����k�5������������L\]../Κ��x�+���r��5{k�5n{n����Ū�q~\W�լcS��]LV+�j�+�z�J�{�m[��ZY��ޮ5��ƽc��x�1���V5���w��b��[����LxӶ5ں]�-V�ے�����ۅaX�]�����鮌��ϗ�"-{����M9�	ʃ�B;#��Ղ �&�1ȉ�������z*z{�.,xA&{ti>�f�Ͻ������zf	�'�X�{L��}��\С%}[������O�m6���hƗ��a{�Q�D��=�����/�r���PRH��#o�"	nI�-[�7eB[c$2CBS���^I�?���0�"ᾖt��:l�a��,
D�f�X�>��I}`p�A�z1]�d	�K�*	��n7H�f����*���3o#Yg$�87q��)�ڎ�L���,��@�����|�B<��LqK0�3vR�C|��(O��7#y*ER)+僕��O34r#��h�G���a�gۮ���ʙB?j�z�*��1�]�s=��-�pw�/Ρ揳���lj�{�֍�wtqL��M�	��ld�e��w0��ݹǮֈþ�?���4{�՘�ܥ\ �%���j[��5�:�gN���#3��!A!��~F�*�MV�o؂�S��ť
N��`���8�
��϶����T��:��o�d˵\ �f�v�k���A��M)8B�{�B.n�c-XkN_{����hԢD� M�P�� ��]w��ɍ�k�,-66����>�h�)>�����ftl�]���e<�Qo�k64�~���"�b�
�(#�A��8@�� �=�SfM�	�|���V[���nb)H�.n8ws��tW��=�
f�b���Hk�8�s�GU�&C23�[m!@~'j��������D�B�|LSR���FO6��N�ɛ}�p��;�L)m6*�`~�>g^�����2U�y#^]�}MSUp5�G��|~~������V{����y�kO������{����y��yֵ���Y���ub��{Ϗ{�ֵ�{�33Y���*����{�ֵ��zz�^�m�o\6�֘�>v�N�Hp�)��׌�!I
x�i��G��{�|�9��b�M)���uk�kJl�[�%�Vl麖���n�vҹn[u��wwY��Zɕ�y����o~+�Lj]�ߕ�u����
a�k}���1Q��(�K���2�.��s��7�I$bC���v���KUmw
^5Z�/�Vb�M?��p��٥��d�����y�&ӏ�ꦣ+i��-z@�����N:�m��X�g[ãI��:s3��r9 ���N�aN�>�94�ޜ�4ſ�o=�2t��v���ɞ.;�ӡ�h����Ҳ����m<@�8i�i7n�*�XL���|�2A�Cǌ���x4ݎM=��N������*˶=��-��!CU���!��	�C		$0�&Sv[�s��n�:�4�)�咵G�NYŏ�\]]�t��ɣ�������%	�X��4pJ6Y<w�hO�tk�y���1�bC�p?zv�.��5�f�_A��Ԝ>Sb�w������[_nu��L�p����d����3�ns�g䚜;�-7u��ѥ>)�c_f��Ѡ��|�����.����i%�����?zQ�iO����E;ˇS�<���Nl�e\��T۴��X{���	��`�KQO����z�R��Y���w��.[�o`i;�#AD	��'nb�����Vg3�@����dd��*���>pPե�s�%��iU�j鍻m��m?4��>vzS��4J||hS���s\���@)��<H��O��D��R��J�Di��|�r`�����]~�m�WZj7❨ōOc��#��O��� ��JvzT%zǩ�N:�B��w9�[�13�N���+��zR��u��TĄm�,4�ൌ�C�VĜ-�M���6�#�����K��0ɨ�NԶMǭv�u��W�jƞ�@(�$t���u+���m�i���M���]�iݖ�1c���0������OL�>8dN���G�tk�^��O%�989jǋ'k�JǍ��8m�4��<lN	g�e����&�F�QQ���l�'^��c� ��#��(�Q*5*�2e>Jy���ë�4@��HF�#}F�Jz��>˜O\P�C�_��6Ȑt�Uf�Ħ�.��4��rt��?xq�-8b�M����?@��1�����O�v� q���K�p�)����#���8$e�h�q-��1��v��B�@�$$(8GK�0q0�Eo�"U�2�/H&�[jnY)եɦ�D�I�Xp�Rx9�j%q!�!��0Sv�����I����tٽG�ۑ���RSM<i۶��%?�Y�(�d4x�˻��|khˮÜ�jby��_:��ד���^jLMf%�%|�ۣ�^��5���M�������⽲��iuu��h�Tm^��Wv\�_),.�w����F�c]-��I�luN�zc�1!NΉ�Х���Rޮ&2�ı�c�c:L��\���>>N/��9<�|�{i��T�B�4�G韎����Z2�����	���É�S%�!1��Kԍ n�.x;��ណ�:⪲�lE<gX$���jB|[׾�HG�5���J;M.��	�M��(w�%"dމ,pD϶w,.H[tD�p�{L.��` ����V�ܔ��h[5I��@�C�>̄��6�9��I[v�8�����M6���_w��S�*��2l�N&T������"����H�ʲ�̊���~�fx$��Ӎ;~m�o�i�>~c���8tzC��O��;�p�ٮIûe{c�1 ���8'	飦�����a�kp08"�!�o3O"UP4G�L_���3����Ƀ�'
w����rE�Y�s	��#p��X}����I�΄< ���2R�	���7�Rz��7cJt��\�j�y0f)�HpC�g>_MGa���9������li�5�Č�&O�f���p�v�!a�<Ç����<����KdL�aÇ<{��Lћ���%$v@��
W�і:a}3��|���-��}CD����!גJ.>vR<�YG�4Y���x�<lN	g�e�йP�]؂dXE�G�1�)I�(��  ��!���P��N+��!��s�Dv��)i+�*$o	�ل��bH��I�ϸzU��Ρ��n.4�)���:k�[V��I���v�Nw�Q�휚r\|O��h���c��=��>�+q�Ŏ�z���}�}2Y>S��o���	������Q����R�Q���[vt��ւF�N�,ɟ�8�$���L�+n��w:���k#s��wm�La��O?'֛"e�|�yH�r�I�L�PY��:|`ᷮi��?1��o�|�N+��+���2$�n���9����б����1�b@�t��`�p<v�d9���A��?L%���C�;��W��HTSJ7�����fFu�m�Y�<�1�������{�'
Q��0<@��KԋiG�Q�	O��D��fRRh�~��ٌ��i�'��DE,ђE��|8yg�@�����q&��m�h�rHɢ�Gp2@��49��&���y9Y;���V-8�J���ғ���uwUMq4�C���ry��MɊwܴ�J���6��Sv+ͻ iǋj��YdS!�,��[c��|���1��<iӊ㹿|*ķ�03Eɽ�h@�"��7
�$��ƚ%��-�3{�f2�Zs�ˬ6>�sMK�	�1KKm��K;�n�4���mf%�D��!H�#4�f��� 
f��K�[�/�1�bB霝e��}��\��Yx���%ҹ���%�:��}'�h�Oqi�G,1�M�j�^1��6��h�&ڱ��M>,�]J� Y;h��SF��[�F�I$v��D>J1�j�i�t����� �LTfu�D*@�������Z�a��ݹ�s3�H��$=eU<!����9��`���	Ad}"JC�_��X�
���'��l����[ к%2=`0'n�����Z��L2�&٤62�)�<�Ϸ9��p���ȝM���O�yW,��x���~~��T�o�یq���i����g�	bt�e�����j�J%��e�Kr�[RjѦ��ΙaoMmb�D���ϭ]���~�)jT�@�z;���$4���h��8@���eUT���9Ĕx���g�zd�� a�������O�`=�!d�����/h���
t£��]��%���ig#!{�*4B��	�?z����Q�M;�H�#h�B��[EA�ڿ�~�"��83]�J��z�U����8;��s�����7�g�lz��G�b���x��;KZB��I���.ˤ�����n�����aZ�"@�2D�U��jq�R���іbh��M"�$�4���, h��x&���s��8|C����W��q�ƺ\oW��b����\sW7�Ŭk��7���b��\տ..>i�[���].��j�f-�X�f�W��b�.+���\V:iW�]LV/������>~i��?./�j~xQ�+�Hx�� �(I�J��[�v���x�L\\c^.�k�b�������KWkk����1��X��������S'�x����A�x�><_��d�O�kLk���Ʊ�^./�u������\���~c].ץ��1��V/lk��񚵏Z�o���q^����|�Z�5<��71X����OE9�QɊ��ʈ�����.=kj����1�f�����b��\տ..>jg����].�%��,�嶫��%��D�(����:�'�A�޹��3�.U�qӷ���.�d����d�]�n�j!�~�
� ��E��k8�����to�L%��޲v���z'�n�_2�oQvg�z��z�6L}���~^~�K����]0�?Gz��	C��C�9qA?m����b~��+��{~qZUW��{�ֵ�o�33Y����Uz��z�Z�����fg��iU^�Wۻ�l�����{jҪ�X�g\�3���W�=q�\6�֘�>:=4��M�FD�ˬc�!�����:��8�6���ԟbI^����@�!f_�a�NDBaѧW����3��`�n`u���8ţͶ�8�s��g�͒~���5���&�ٓf�Y�-��G����2��fJNe�Y0!i�L[a���hh�Y5�A��d�옩$[C1xA�Eq�̤D\&>&8� ��L�2}��EUnY�W��RoQ��0�;ߦ%_���X�꨺M��4æL�a���Pv:WN<q�\6�c�1��<h�h�����98B��t��1�A;�̸'N���9!m��˺����'��2D��QS�!���[Qv�:�P����s����^|�<�lb�f����
G[9N
����$�8&�]�I,�L�6y�Cp����g����iF��fh�w�(o��� u"�O��$^���TQ�;7=.�h��N��յ&1�M�罒��2a;��'[H9!��ȟ�h�e�$:%�����#�=�G�Xz "i�fo�_2�ex���:���+qb�{Q"�޵7�bV�H�����"x��x�>)!i=
)�dK�_�9ñ4p�)D�:4�Э1���:c��>xӧǜ�W���	��ƺ��x�{��@�8��B.rr�󆩸�v��q�R�H�m��N3>�(�9(�_�d`�X#v=2�l�h8$e�,��Th}~h�Q���e��c9��#�w�S�jS�1.@�t�+K�h�du�*�3l�g�m۴��35���.�0���q���$$��&�w�֚%����h��7u�����B��$	Id<��&å��Z!dE�c%�=�EQ��>#��ኵm���jY_��f��CҒ��Rl�PQ11��I%J���)lp���H�6RMv�a�i��4[��,(�,�!�E.�� B�grJ��yCĽ����
e��փ8C�L)sIM�(��	��x�����>'��"����5hB8�d�]R$�	���<9��bp=����;�
'A��
(`G.<�z���x��I�b?��e9���ǑS�����v��Ύ4����:a��d8h�xz��Q~����Hҿu4}=W���N�j,<�N��������%�������~ɇ�^��)�x�Y<��6���r=ꥦ�$�\O���v�?0�y�m>|mm 䇒�SE��+�$�鳞����QAi4x�:�
O�gx��q�,�|h�7	Tl6���h�g0�ñ89@�Osr���Ɂ棉�:A}�V�u��{FV�tz��:�9;v��1�S�!�l7�2a��	Ef��ph�S���ߝ������o�������t��/��D�B���+~(p��ɳF7��L ��w�)������jv�6����4�O&��E������M8HQ�%����;�qvTԇY�!�[����w��9�Rd:N�|�S�<KF�O`�|�h���4��Y�e �Ͻ���E��ŗ�|,!#��p��&���]<�U�c�5O��{���K4�BB��4ȞdVH��=9ѡګ��h���W�&��C	�2n�J0� Y&&�a0!�Ǵ�5�I�������tv��ҿ;m�nߝ8�?6�����t�]8�:�G,_ T�G7fg=���_{�$���a1,c,^ێ��7ٲi�槎�ɜ(�o�>�S!e!kӕRrX��S�]�.��))BP��7��,�i���&$^�m�'�	$$��h��8H!��
O!�N]�a�:.8R`A>�:���^��m�R[�v��u����O%��tI	Q�`> p�9!	'�ك$|���v�&S���.�p��s�%B@˴���!%&F���r76jiǲM�Em�c�޶鎜V�6���Lv�:x��WZ�����i
���>���h#h?Q6��j �_K�H�_0��Ӿ���H0��kvK&`���c�<���`бmI�+�vib��wN�k)w�n_�� �@=	g��B|�[��l�ku�̖Y�4�e�ޝ�F�-6᧩���~�I�LUq��˖��Ӭ<�p���rϖ�/G-�����i��DJ&4QOx�2B�F-:���1�T�#�DVI7ӆ��'G�z2}���E�����'_�X"�4;�ז�R�>g��#Чj��z�����?i����5:m*��m���V�Z�b;l����]�K#H��I9��E|�N��8�Z|��)
!q�����m���M��ۺ���tzӶ�����?:qZ~m�����t�]8�=�D�a܇��	ȰE13P��#Ėg$7b���$���a��D�SI�ނ�J㞓��"1[�����$��*B$�l�Y	����pi���q��H\*I!�.H!���[#i���D�d��0�^&ry�sDI��ST��$���?7������O�c�;�
'~�u�ѥ�M��b��8��0r�.HBB	a�� �	�\�ve�wRBL��&_'z�pHn�R���ܙqƓn6m��߳�v��քdA�y:TPQ
��R2p��<)�ӆ���c1���q\]�n�Wk�����HI	&O��n��l7���m��&?I���XC-F@�3��y��&7I�M%�2BӉIM���I�)P�=;�4BV:�zC��\��{�T�{P�Cz��o��J#��
ɲƖ�Q+m[X#c�|i=���GZ-4k8JH�zܒC P-���q-8i�`0C��$L�!Bc�J�&��x^�w'b��9Řu�ްJn#��Wޫb���34O���pғ$��4p���~c�ͺ�V���t�lc���o�<y\=�U���.��5#/��Beax�����H[\��58}ߐ�BI����a�N���e��`�����<�(���8�,�G�!��ai�����y���80H��H�9�����tݺ:�y��a��a���\�ߙn�L���;i�� �Z^KN���,d��óF��Ç�5��IN�%�d�����2���i�i����"\}]滌��r�_�Z{�a�{��j���el�y����G9g�Q.U���4W^!d5�BH6ͺ6}�}	Tƻ��j�6���k�8�W>OHi����N�pt����V5���wX�..=k��N1���X�7q�t�./��q_1�3V�֙���k��.�
���̖�-Vb�Ū�b�ݵ2�5����.�+���LY�������OU������.�����X���U���=k��k���\c^0�./ˋ�MaqqqqqzcS���/��t(��!������?���>t��./jºcL\x����5�b�ƺ]1��Lk��q�\z�-\y�����qX�cLWk�L��\^�լv�/�4ǭd���N��:O�x�I����Oxي�}n5��[<^-sWmZ[maj�[��cx��z�3Wָƪ��L�Ʊ�X����|Ƙ�[��{��q�j��p�+
Ŷ�-V���Ua[W�_���,����/I���US2.e.D�<\���[�%>Up��>λ����x���۸�;�	βj"�(L�3��O��kH��%"�r�ْ��|ł����#5�)�0���m���F�����AI`ܘ�U&�����M�Fe��h|(�� L��$�#D(�Z��90m;����QP��:<��o=c��ZqG�	-f�n;jh;�B�q�-��)\�$K�/�~�=ßco�j��������K	cmV���ƞ�=P�_�I��.!��~s�#�O�h'[�)K�;Qf��o(W�����>�n:u�l �A�4�&�j�N�m����-ٗBWe�B���p�n���L�ܔ��9� t���TjH�jL���� ���� ��S&����'��U�i{��`i�gaK{\9�Bp~�r���*dBI �C�J6hx|�sV�����֯39�ۧ+F��!��b(�Y��TW>�q��aB���v��4,H�Za~�LSF Cq�P �ɴ�R����f�,K�!�)k��T�׬{�+�6��ң,\�j���AI����ǭ��ɍ�7(��(+)/�������WG4��-�5�ٛ�]�W���Z�k�M}6��]��0&l6 k
���u�X�S�u�[R��Z���uJ2�MᬘB(���P�������p��w��γ��ʥ)Ĉ�����P�z�8�kn�
B�]d�&)#zl�+w|՛��h���;�}s�ڴ��V+�w������{j�U^,V�w~�33/3=��Ux�-�w~�����{֫�Uⴷ����00�Eaf0�����t�lc���j���jn��˭�]�&`���a����a���kK]h�c��I�	���R�_is�� �Gv���KZ�oC:f�,�ڮ/���܆c�5���ͦ���m����K6�u��&���%�&���]K��k�M�M�V2a��&����^�<:ṉ�b&���O�����I��ݓvSLc���a���'aAd_�2T���Hl�����(�����zã����	~� ��
�t�[�$9Gч�2Y��57
��gxvo��9�ӂL::��y���Ųt��d�6�(i�yk��+8����Np!��J6�2'^��zW�]\�!W�X聰ɲ�x�ǭ�ۧ���1���tp��_�T���dtn�;*�j$���a��\.'�g[���=p^c&��h�ܧ�0���L�I�NͺJ���n麻��zv�1�Hm��=R���&S�rUx�p� P�L��۷m;���{j>vi^�~O܋�.v�KfT>Vm��Bkm��H��ñ>���8s��ϿB�J�B׃'��	&KM�<y(8C)�8O&�u>$:���M�!��z�nƎ��z���1٣�6��8�N6�_6��:c�1��շ���I"���&v�s\ۜ�����8���w�4���BHI0�Q���	�ɟUU����8x��/���vosOǀ��!�\d��'vkĪ�ɤ�����,�i��'SD:�ۣM�'�F�1/�ēfڒ�W&I���<F6�JV7FK!�E^���
*����� ��Ç�g%���8p�^m)���u8�z�T5T�D�]�����3�E��v��杂#�w��!̧[����Z4i�m?;q�n�m^=m��(����䵷��_��I	!$�	�\p>��I!�>��I8p�6|S���*I!;t�9D�����s��NΓ��ti]�C]�l�5�m7I�4ցì7�w��|a�W�Q��/&~�{����w�������ƥd�Cd4�����(�y��|`2Ck��ޫ����8m�6����UXO����!z*B��"w������������E�֕d�U�[���'2F�#��q�ɺ�܇gGn��8��m_?6��:c�1��ն�WΏ��R�����f�fz��KZRY�p��;��5���k���1e��i�I��9�B�U���gwiUҾ/�-I�z1�bWh��7�0[�C��ڶ�V6!V�n$Ck�4.���� �@=	gO���.R]&�$�������᧡���@s�D�ט���T�I%�>"XBEpx͜2h�l�aD�/R�U�]=>�Y����
!@����Zds�EV���\y���)6Rky��8��G1,�u����P}�G0�@�o?q����cZ#5�]�`�hM���G�	$�v�}	$с��!nR�i��N�d����xCp�C���8�q���6���Lv�:8ڶC/Qp��p��rBHI3&����{�8u��}|al�
�����N���2���[ԭ&��ܲ���u��'�'M/$>M�c��4{�z0Qo!�{Č�c���e�R�k�49�l��e�w�46w���"ۍ��[$��i���u�3!��G	�f��;�x���y!�ɴ��Їg$����b�z�*�6����,{
v�X���m��c��?���P `�-�Y�c�b��¢k7�y	!$$��g����,�4�u�(��݄�q4�O��q86�:Qj�UK���ppR}}�G]�&�N4`��/�/�8d������d�[?$w�Y���q�	�l �Mil��i(��Զ�#L:��>J4	0�xL�vb�Ή� `�x�Ӓ�)���)�H{F�'(�I�f���ג�nmp�2�(uP	 %��h�~fv~��BGb|i�OM)�!��OO��(�b����9�$�i:�&�C\�}�!$$��1p���G�i�2=~o<*T(�L��#��?�D�VaJҠ2�i4lv��Z�ܖVb��1��4Icu#(ʎ'�g�<,�f���O�Cf����Z�I�n҇GSGu����́���,|��[��D��i0�|si��+`h�FK<�0>AE�;W��H���,�vw��0��x���$d6�l�>\�M&�W�:q㍴�O�~~c�;c1�!����I�Z�6Y�K��[MU1�m��c_�Uڇ�W���p���"�T�����b:�s�f�'�*�k�㥛rܯ�2�n�V6]��_w*E�Ʊ�v؞!/�q)�����8'�����XXc�
�W+�B��3c"�UWv��<OwN�<�0�}�p�x&N���J�2f�u �>y�Ͳ�!�ɱ�s��z��5*�:���|g3���(�h�8��I_qYP�擦G���a�&���9̜�!��r�'�����h�O�率�JN&��mp<��\!*�f%LLB��5��0���H�33�����*/^^�_�(��3s�γ�2r�X��L��y��BhS�Ri�f��q�������j�L�j�wB��3ٍ�.ǐԹ��6nԸV�6�I[��g��g? *�b{��������<}*���)�ڔ�fW%0�&�G��
e�n����rB>�D�k翤*^�SS�7��w�0��-!��0�p����f�i��ٮ�DΦ��p6��b����L�Z��Zl�h6Qu�&���`Yi�"`��Hj������2&S&�i2�)�d>6y>��	�/U'O�ц�rK�u�JƝ:m����~q���ADЈ���� ��"!�DN��bl��B �"%�%��,H&�N	�:'D�0L��,L���e ��0Л �N	�:"'K
O��K,KbX��8"&���dd6"'DHpK �x�G�G��x���؜:lN��a��b"7&�%�8h4%�<x�Ǐ0�㦏$�D���pDL8l؛4P� �C���ҏ�!�ϳ3=���=s>��h�ć=�������63�)�{~kW�t�`9ĔRE�Ϡ0��I%.�ȩB����2{�.�0��:�`�`'H=�=Fxn�����u
���4�*���|��>�[�(%A�鬐�P8>��E��� ��{G�"�{����c��f>�8O���1H.0I�ke�2�� C���k�V����3�M���ȁ��=9�p#�����~�u�sj��t��V���~�fff�=�UҪ�Z[�]�Y������U�Wj���������g�j���U�|ι��^�֞��Ǯ6Ҹ��c>:>4�B������$���`j����g����x4t��FܞN��,�8pɽ�6�)�2{p��@���'�CF�&��NӉ�A`{'���k��l�Ҥ�[�c��FM�r�8d�Y퉷F����L�@e�d�|�ӣ ���d�g_�N]���|SGN�����@3��!1��SGԑ� ���>t�q�q�~~c�;a���>�C��d|���`9>�BHI	&��$=�3Ϙ)!�y���ɳ/�:R'q �3!�I�=������ke݉t��1���[�]��Z�1�[4������=�h{�?�������l$��'����Y%�1�t��q6`�@h��D:bH�ȘC�X�0�s���@3���X�~Đ,�[�"�8��Rp��6Rc͆!��=t�i\|��?1���զ���0 �����:B)@��II�n��^d9�LG\-a��N(`֫�TL���rR�U,�F�+^4��;��ī�^��KM6ka�-AшJ�6��ץ�;�@ H��\̖���&v��
�ɭ�ڡQ�i�lmel���$����� �t��=�r������ӯͽ`{���ǉ��4�|b��%UT�������׎�>D
a3���؝��~���*^�-���8y�V�;�*�>z�񺒫�M�'M�3IUҊl� h�8��0�϶�[
=~�y�8I6ќ���1�ڕey�n�T�T����߂�{Oyr�z|�I�&�!+�S;M�W�>z���8Ҹ��1��Q!���'v?w!$$��3�S��~*�ΦI<�<��G!�$	2u�i,�=ptɃXy�U�*씜J���9�iml��n
�y:�t�ޕ[O���Ƀ�k9>�V��L��pL������bT]�n˦�`@���Qt����O�l�Г�:|X�D�i����Ý��ܝ[%�W�y�ؙp�����鍤�~����gGN|a�MOZv�O�8Ҷ��1����6��p�lp�eH��GS-��.Y�8�O]���L�p���Xo��*10���CHm!�=�I4��i6r���+#s�j�U[yӥt�̎�	k�)�6D�E�1�=�owv.�ۅF�6�$N���9El�Iz���㇏��HH��$�j�2>�*��m4�����̡�z���6|d���9�8{���*?2~�_v�K]�d44"�Ɠ)
Ju��F�;Wm1�n���J���1���������"g��	!$$��
Y�rꪟy,��N}�0�����9���O�?�[lJ���e-�G)6m��%e��aa0���b��G�����:;��oi��$�&�զ�{Ð�D�<2�h���>4g�R�q��z��^�6�1N��&o�
�ps#N�)�%&��h���J��0�(�`<Ѥ��c����d<����M��?6��4��1������J$!���;�%ݰ�H���g�}���~�R��T�^щ4,|]Kct���-i���Ӌ�:�l&��"I�s>���2��#�P���1�!C[(�>s��7��m�,r�>u#4-k�~� �3�UE"N���Kz�,Ѣ����h�td���_ݜ:>9�Ì�;����LS�2��⮥T(��`}���Ko2��ã�G9�*W6��I	��å�|Y�[Ē��4�%���T+�ڥ%R�����8S�K�n�VVRN��}���3���j�!Q 铫Ԇ��+$�?g�5�a�%����35��7J���}�&JN�}���J��������I���`��Um2�J�!��=m��4��1��c�;c��M�{Ϊ�Gv+��k�L�y3�7g�f�H�琒BI�L)�u(hD�C��y7u.Q��y1��+O��`q~�>��C���J�u���-�fu%��@<a��I��᷏U�L��,�u6����$�(�\?'��^<�͖��5
��su�-��"A� �[8	�EN�Fq���$�S9�i6��S���>s��⩣��O���I����"��s)��Fx��9��ގ�<9.T�UQwM�=w9�p�+֘�Lqƕ�bX���8x�D(��o�7���w��~�aS�C�%��k#y~u�I����ZM�T�^�RC���:�:a�6���'$�y&�%B������g�(�ω��p��{U,}۟��N���ζ�n��2j�eS�x.��L������T> �d��m�I�'�HI���^�N�!̳`h�:hlcp�ɂ�F1��WSc�|ӑ8�1>�ʺ�8�g���|�2O�V4��n���J��c���(����K�ؒ�
=8T�$��C���C%��.�Ė�4
�\�<�Oz�BHI3<�x&��|�2ʫ�%K0d����y<<8��[�ü����}����"����˔M�Kr?�+FKd�
y�gg��2�L����(x�<Q�O���U�QOp�\���x\���L�<�$�*��0�L'I�F�96�_���S��C		cI�g2h��F��|Jӳ8x����+(N�=����UV�v����9�x�a�""hDDL��DK�&	�0zM�6h�B�AD���bhK(؉�:&	�0�	�l�(L���e""&��,D���"pК ���"P�e�gM�b"p؈�8%�D�D؈�"p�,��D��B%����㇎�<a㧎��0J0N���&	���jO��B""`�0����<x�Ǆ���pDL/�؛4P� � ��ܣ���W
�ܭѹZ���׏ҿR�o�J�wl9����/_t��bSs� Vs��љi���n�m
��@�_��K���xM�\:���Eѕ�
�*��B�]���'fA�`AW��5� ���ʳ�϶�:L!�Õ�I;� T�p�s$M�8��3}�D�wN��2|n����,�"� £,'�}B8o{9��ft��65���t�X��C:��_a��!�J�("��i�Ό��w**��͌4`b�Ο�w�%;ty�E�;MJ%�!�v��d'L�0i� �3>f��:��1��P�5�ɵ�������p�7�+PT޳$�579��x��R�V3�2�l�����í�����q����T`5ʨe̠���I�$���J�A��^�dyͶ�"4UH��5�D�"���C�[4����ԚLb���\�H`I�&�B���۬�߻:�Y̵�ikr����0u�͉}����o��r�Ya\m��[���������J�(.<h˓n�fr�(����jh�WMڒ�R4�6��	$ld�@Q������A����Mj�ŬkDЙ	q$G��K9S��[�b8K������:��k&��Kb�?9��c0*�2��w�	�AD!Z�H�'�BB0��mE���Y)�PB"�N�H@.wg������Z�z�y�9��UmUڮ�����333��iU�Wj�n�������g��V�]�黿_�3339���Wj�����~��0�a���Ye��,�����J$!���I�=�ś�vi�����dM���<lͶ�]�$3P�ͲkkLb�m�hƅpm��h���,ٶ1�֏��J�&��p�96�3jE��}�m�+5���0#j�O2�7��j��T7���{�"muq�m-ڒ9�i`������$� t�×.�ќ6f�8z\.�M�I��Pt��Ą�w��OzJN&6��Q�Ϗ�;>�EU�X���㪇��2U&�����a���t��I�)�	Ӝ2<:��}�T�V*�b�7	�uc��pd�'��F���&�6Z�wJ�2+=���������T2wчd쯮˹IgG��6Ҹ�6���W�=q�����`� `���T�y��IwsΉ	�:�y	!$$��.�=6:a�'�H0�i>6v&�hn�d��O$.�^���)&w f2�<�%�7�|a��tâ��g	��G2�T��o�U�i��<uj�s��������ދYz�X���[��)a��H#�Y�f�-a�a�z��}�p�_}�7����I鐊�"���8G�O��RP��'\�i�Z8QE���ӂ>�zIÃ��d~MKnI&� �l�bYe�ı?Q!�3�'\���q�ƫ��6��̧�	!$$���s=�{R���J<hxu#y��,�O��,��r9LY���p���?_�|>7��Ø>s�"ntg<�����e���݌Cliu��;�;k���R�����if��óܧGe��:2y�
1ߎ��f�BT$�<k}C��v���;M�Nb�guW���E�)���b�+'63����s��u=��}78z�Xӷͺc�4�q�������J$!��5r�)9.�7põtUQUEU.L�����]i�����C��Y$�<&�_fS%v���$l,�Q�ȖJ"�F	��v�ݝhxh��Q�ǜr�}�*����kgҽwr�S4;tzl��v�=��k��߸Lzʹx���:�}�����7/3�"�*���辙�JL.Ç::�C�	���Ux;�����^&��M�@=N\$<��v�W�<|��n8ڿ8����؁�C�8���.���2������Wπ߮-��Y^ �2h��9JQ�j�b�a
8+-�ӳ]È�\U�vG�L�(	H@n3��}��gF�5���ǗKIKxŔ�h�XM��.�1���M"F�%l�]wbܐ��ߦ�*R�+-�(J�.�Jʈ+"��$�?�I:N�BC�r9�	�n9�ZL]����L':�09�$�n��\0�����I�<Ԅ�Q�0y6>8��s)n�;��Tx�6;�ު���Hۿ8�����OC�����u�%�~����;3xQ��T�"0�+R�q�f�<�`�'�����)�G&ꪫ�@i7N�N��Iў�vCO�;:4҉����1�1�զ���/)�t���z�=鮖,��T?���C�*i( /Y3��R���vT����UU]͙��O����g~�+G��|�88Y�G�K�HIUR
�L:�ɑ�ˮL��D�����l�-��u�ݪ:M-�#��>z\1�>�M��0��s߽���8*�˶mazW؇����K!t�;�˄Y8�0<M�R��Rߓ��{:�a��Ɲ�m�m_���?1�1���w;��gm���>�	!UEU/Ň����ɓ���Iܭ��Xf'3��!�������L�Sa�h��9���!���0�Lh|c�G��-�珉�΢�X�!��(�g�e���ز��K'#�\QV��am����IL��6h�#!n@���w�6��:2?��p�����9��r�o!��ٴ�\�U2����hhG�wG��2p�
:t�F�,��ͺ|�;c�8ڴ�������p[b���c�om�7� �@=���G����\�E��;�~4�'�e�8vgG��|����wJ$�rZ��;$�-��ώg����p��f�L����]ޭ듃����ٿ��UD��(��I��WJ:7��3r~<;:��1��Zȼ=Cԯ�	i�q���Æ�>xUQ��ݺZ���}�΂����Ό���ڶ��?;<m]��ͽv㍫ǭ�>?�Q!�q�>�ݓv[$}�4`6<��.���6�{Q:f6�-e�u?W�d�	�J-|��-8�Ŵ�!,�n���0B"�I�7�Gk��r�lp"G4�6���`��K��Cf1m5���u4�1q.�o�m�]͎����~�� �@=����[����3Lf&�̉.Ħ���R�lX��s�d�y�E�>Xl��~��R��M����>��˾�Hx��_s�IU�M�����
g�,�d�i\<4��;���Rw�t~pࡴ���e,��9EV�@��o d�dm�e�P�u���r< �/g���/g�d3��E�Ԓ׽������ͺ]��?g0O�sd���C~�����4y�|Zx{mR�|iڶӧ��mۍ�ۇ���G�gƔHC��uZ}&�ؚXy��X%ݱQ��&G\�F��u��{�$���f8CC���r;1�h|S��O��M��pq8h�1��v]�����$z���Ȍ�hkp�L:O��טB= z�N��8J�l��2l�P�C�x!��}������U� Ec�1
�UR��zN&�>D���ġہ4j&���9��	�=�[ɓ{W�l����!�3�p�\Þ��tt$!�Ǝ����(�"A,DDL�"AblDN�DN�pN6h�A,AD���dM	�bX��`�a�`�&	����N(�0N%�N�(D��"`��Bh���BtNf͉b"pDLNDJb"h�BYe"AG	d�KblD���0����"Yb&	��А '�&�DD�:P�$<x��ǎ�<'�L6&� � ���b�������F��lx�Z9,ݖ���Q��*���ܯӻf��u�6��3���]9�5}��͠뇮�++I������+����3�B�փ�S@Ȇ�^^�2�}Ҍ��~Vx[�14���T�d��o%�d��=n"T�>ܹ8�^R���5)���7l���ϱs����Q��^Y�ޣUQ�P��>+yr�!i������{�=[�>�ǳ���4�I�{uFp��t<F�_�����?[�m���o
�w��O�g��{?~��Uڭ�黽{�3333��*��mU���zffffwޥUڭ��ww�L�����Ԫ�U�V����a(ǭ�mۍ�׭����j�L/m���L�2j������} ���00,0�:L�P�?l��%�p~7Q���/l8�hw^����*�4�M�0��|}4�ޏ�|Q����O�Ӄ��C4T�J��8 ��8��bBB���ѓ�^��LT��y��y;�E�Y��7$���2H�p��3R��V��ɐ��5ս6�ݸھz��O�vǌq�h�࠽��=��e�(�&/�A]���I	!$̹�î�t�*�
Ĩ�ę!��6;KO�]��ө���+��!�0�I�~��o>L"�8�jN���tٲ���-�d�t�z4�3��)�e�z]��9}ǉ����rx�j�A���T�ԑ|}&�x=��όo'�2T��y���m���)Ǎ�K4����=>��ݛ;s0����;4�������ںk�}m�n�m^��:~>:>;>4�B|�C9c&)�u���T��~�R5E$1P��,쳵zi}G+v��ms>��竧7�u��}��`3�l���D�	7(We¢r�]�1�di�V���֥�oe��[����:���l�,vآQ�c1u�M�����Z-���a$$���\-�1#e \~�S��L��Ԅ�������F���������ٛ'(��r�y0;�q�����d���^�O�Ri�1�	ͥ�!����'׫�$%QW��G��;Քyٱ��G�&���I}�&�����)�mçhj)�L8c�T�(����ufZ(�l�A�*m�ՄV�u�M|h����{��w;�b�|��}}3]v��1|�ޮ�W��_[�o[v�j�6�O�vǌ@�/��N��9~ɞNv�oud.2sE��}�QUEUT��!�N�riٳ�>��HFI6���*��i�z�8�I
>l���a��;�צ�_}'ȴ��L�D(��:��R˄}s8p����W��ו��q[��m�7K������x�S��y0���;����әͶY����>Ot�M�0?&�8֤�(�UJVG��;�z����JN��҉�����G�gƔHO�OBa�$��h{��HI	&g20��	�q2=�$�)�5sdR�N��4����d>9�O0�a���}���O��t_��׸������s��9s��Fr("���b�:����~0�[��$>)�F��4�Hu��q���^�ejT����z�5�2C!㻢�$)v�k]È�M���/�2zu7:�m]������v�Lco�v�lx�V��}�=���=�h�����N�z�;qy۰�	��/�F~�:ޟ��m�$��d��K�vHl"�V'�B�����A���	3�K��ɦ�l���<.tp�=#if��`:x�mvw�UT���S,
L�~˓%�p����ɦ#ͼ>xJ�nǦ��
q�:�NÎ��Z��}��cJ�m�Ͷ�1�1���mZk-��/5�ky��{=��x	o/���O�a�β�X�<$��SR�����'6(E[�p�ݗz몝"��[idl��pu�[[9Nw��������m<���L�.}b�3Vk�Sl��ں�{Au�i�֜����D ����>���iw�{;���z���K�e8�,,6�W�=�92'��>�F�_���|��$�8$)�+�ѭ�-(�a�?H��H��gS��7�Q*�f�|`�N�ǁ���h/>}�nʋrA�>$�vn+�v\��3N�7
hu������#G������1K
FB��U�HL'\�{UI���XH�0�.��n��J�*9����d�I�����1������j�Yoz����9���Gf���$���KJ��UY8h3���*D�����f�%d:�x��SM�&~2���-������α��!�L�-(9��.���UT����e/y�މ�]L)��{����9vF�J�Q&�]cFB�=�{.y�a�QQ��a�|UP����%�p�>��M��%�`4Y�8Y�ͻm���|����6�5��z�L�K��"!�5����D)���������	��N��C��I���?f��&~L��FK!O$�yߪ�U]�����ϒ�bܚo2G��n�ȥ���u�Jf�:&�)R�t�it5qG�3�;3�>x��B�̘�n�(�3�I$���qV�d�}UQR�J�@۟jy,��%�=�!���4��	�9�E�� ���9���GOP���ْ+���6��6��lvǌq�i�VSR�%$=�s��Wyn��6Q*A������l���9�2{�h�����I�0��i�Am&v�֯<���Øs�{�.Vk�Mkr�T][�,Pu�2߽?���[�����(�hi'��r���NԪ�<�&N:8�R}�M��ð�2��������հ�R�:�xl���t�p0:��a�#�<o�_�r�R=��	J��a0��d<Pl���KI�͖~C��Ab"&	 ��""DNbl�� � �"`�(ѡ�Љ�g�&0L:"`�'0�L6`tᲬ����tMDI�K4"lDD�8h�H"hН�ٳb&��"`�Q�"%��eX����&�Л�'D�0����B�L:'� @A�A�DL�"A,DE��cǎ�t�M�������~ģ��3uvJ֪����¦��?h��3{i�����럩e91����i���V�N)�0L�8���:N(f��Y����:�����{�8�
4��y߲Uu{n}��]&�	�]zĸJԁ��^��$P��C}���ԜzY�O�����l�
���G�[B�=&�&��}3�pT���3�*E1+�3(ب$�&��M!ĳ8�H"�fvAU�v���J1EGI	,�o�=c�tT:i�"63�j�S	d���ش]f����Y�@���!zL9r<W�l�/�=�{�W��fv#,�U5��[9rD�t��`�7�̍
l����A��Y��b��ZmTPk�ܾ?[ɕc	�جt$��ל�U8��]wbz��7s���h�A�7P
"�Y�܈\b�k�(o��ь9�U�cϑD�)k5?t�MA[;N�AG��f�-
��~�x��@;B�m>r�@4dtpɅ)�em�D�LBu��p%�^��W_km��_}�2�����w-����}�����-����{����ޜ�7����q{��9�h���bi���g�5�V�kk�]dv[*?Lͧq���u��,���tf{��/$��w���̤����,:Vȋ��L�B2���t�$2T�B���bW�c������-�k�,�+�u^��V�GB;kd-��*�|�U�uF�����;������UW��U����ffff{=U�Un��񙙙���UW��U����ffff{=U�Un������h��p�/ˎ���j�k�η�-t���0R_L9��n�l-�m,���A�@�5*�5&&��,�Y��nv��٭gGk&�{X]\F7��-�hGF�i�����[��h��EV���M��	!$�zqx�|gF	�6��
�tc�Y�ք`(�l<��O����QI�%�C�_�������Д����N�T���'L<L96!"��rn���ٌJ�����&�.D�4�t�N
�9Hh�[4q������>��K<�,�΍@�
־���j�J9����M�m�Y�e��A�W��Q4�>���p�7��(��8pN�S�JC�??1��;c�8ڴ����sY���F\�<tx������_{{b(�_��M܄���	ɩR�5EI����x�i����PJ�*e2ӓ���d���̽��;˝��74���)#�.��)��
znHH��~��?p�!�ϥ���ڝ3v�d�H+E�ʅT8�*���V������g���Q(����)��O>x��p�s���ňo��$����'�|��i�|�Lvǌx�V����E����3²�'1���(�oj>|�s=�	�a�(���͉�L�W�$;��.A�oq���T�W.l�c��I�|Gͦ�F~̽�8p�2O#�F�F�Z	�&�0�!�$�i>&^�&����%D�y�~9
4����Y����gF��=����g��G�d�2B�>�.<0��;k�[�n���D5�<|$��XY}ì�:���]ǈ���4��m�o�6ӷͱ����6�1�j�u�����V���r��	�.�u�GP��_�u� ��4�8/R����i�m�s�:�	i����o:���/l�	��NH��;�8L�d�7����7 ��d۩'C�tY��m5��؛��U�/�i���I!�M'L�$8<	��CF�l�I%m+�?!�$b�s:�I�����C����B6��-�Ԥm�S��4d�h06���~����T�ӳ����ݶ���v��ϝ1�ώύ(���7ןw��,+X]j��MC^���E���II�/�	���+kr��30;����Q���"�S~3��Ҟ�fJ�m�N��é�q0
G�qc����c���,��ұ&����+�g2���Y6b�PAv[3g�E\7��w��j��C4C&#�mP��M-��d����K�~�!�:���ϡ���Rh>��������<��r�d�%	�0BÉ�s�M�)��ۨh|ԓ�����ö�ah�gO��y�3
��C�y�M�=�	@t�]�������v��6YZV�z޺���ֵgq��Z�`��],$�U���I��vN������L=L�z�˹Ri:����q�n�v�m;x�:c�<c�8`�?.��E�4�&n0���n��A ��襁/�u��rm���lw���Ҫ��Nr@��ɳ>j����*���߈�3��p�ÿ�*tY�}�%Қ���	��)C�D�>psG�U,m�$�&Eҭ�D٪�.]ث�G8'�g�q�\�<�o端�+��vi��g�O$BwW{٧8�b:����:����F�R��F�-���x1�,��+�v�n�|�m<x��?1��<c��~wo�v�\_W�� !紂D����I	'SN�L�CF��i�C�a�W �E;=Kp����*O'�.I	(�Iߝ��'��|����~��;�g���^k`V�mǗf�vF�Zŝ���������i0x�'yUTO�;�C"|�N�ao[mIe\9���n9��4M8~�eJ�Ҷ��=�ʕG��S����Ǫ��oz�m1���t�:xǌtڴ���y�Vx�8���E]��y�(�����|~)���T�y�Ɯ�:}�M���F�X�:˲F�WjEHikK��m�y���z�~8��a�z�N�*�>6h�W$���y韯�i��!��$9�'^�eLs������l--�s��<��n���;;׆ߏI������4�1��;g�g��+�m�o�6�x�������{Hp��',�Jͥd�LJ�Y08�)��D�\M�.2�d��A(�vc@��W��M8�Ɓ��gԮ��WB�IZ�m�f�=f��+5e�-ه�m���1L�	�Z�[U4��X]ؓΑE�:�C��-5ز�l��ITݒT���7J2������/G0�����U?;�2AK/���:�����2wi��dY>>$��xØ8�~u�g�ʩ
%S*ʩR�*+�ٝ>�����y"m����a�5�W擩��|�{�|���̷;;=힖e��f�wt��n�LA��ғCQf"�zHz��'_��(Ʉ�+'"Y�~`��v�6��c�y� ��Oz�m>i���Lc��x�M�Ls��P=�k�u8p��
D�(���[8�ba��8���.v�����Q�����K�L����aC��Z`��oR������<���|��p�i�j��BҌ�%%��S�~�p&���67!�k���Ϲ�K5!�v�K.̍.ĖX@�~��M�6��>z�8fHQ�7��N����O5$ɴ��M�um�j����z?y8����8鍛?&�~D�"&�DL�"%���	�&	�blM�(B � �,��2%��b'��L�&	�`�&	�"hϺN�,�0N���"&�8$٢� ���8'�6tN��a�@�":�8""a��!���Y�bY�6X�M���tN��0L���'�����6QA�����B�B"lD艂&	��!�x<��HxRL�w<�z�K�cge����3Ϻp�׹��R���[���xx)(�S�>�A���w(�}��wC��v����/qy�MYr�������5�pck����z�b�{�9�o��Z�<l��1[z��V{�F/]���2gDot�[�U�͙�7��i��[�{Q^~�:fgo�\���[��ДQ7y�b�����lnS���#�fp����9[�w���s���f���#;�RQ��A����A�`xJ�W����ﺩ;;F���Nu��{;'{{��<��@�5O{v��W�6�pi4���s�����s��z�5x����Q�2�Zxꗗ�[�8�i~�˼�FJ��%�E{/�������_~�vu���$W/L��k��t����v��0��z������9،z�]���{�e�/:����n-Y�$6�����ɉ�:{��L�o�g}�ì��괭�gi�^���iCs���9���r�}�<�W�����9誫եV��������EU^�*�wv������z*��iU����fffg����ZUn����C4a�4Q��=c�1��<c�զ6�jա>$�:�UP0Q��vlt��ڧM���kiZ!����=�7�o4���?ZRu��Y-�fT��dAI&��z����2��`�̛(~�ꪧn�,���)�}�hq:c�罂��}.(��g�V�};�m�G�=�%��/�=~N�ur`�l��6�֞?1��;c�:mZco���L|ѭ�n^⪡�~p���j|��1�C�Ql:9rd*�!�����m���6��,MMF��6ٛI+�
tD�IԿ��G�2<h�z�BI,:�ԝ�������q8�$!'�>�*�h%�!�ЁLv֟&Bo����vk�7%�0�Z�GR?9
�&��O'sU*�*'v����s�
k9��|�q���2��>�C4pЖh�(��1���6�1�q��Y�o��"Ϸ�;�<�LCjn�s��^�<��>(�����֜�v�F@Px�R�V���'�/��2�مCi�ζ��ܫʲ�c7�ւ�v-�рK�v�訜��4�n����UP�/kV�.-�e��	�}C-s�͌	4�x{����<�."ᆓy�>�1��Lv�UJ��C�Hx�`�g����W�E$sͻ!%J2#�����n�T�ل�ssp��[H�V]��?x/j�nq����C��SF����~������*�!I~C&0�&��!��{�����������>5�aq>8?1$�3��hw��+�E���6���x���Ο���1ӊC⓼7��ۘY���8�w�vU���1$�@�*p�̇��]�zBU�D��B�p6�A�X��APL����y��W(\�:P��M�q�H�6�=�$����4χ���������d���m&㱱�&�";�
���{��-�|p5ɾ����J�J��I�'\<Z6q�:��h"�E�B���h��O�>�{2aZWۦ��m>i��:c1��:qZck]��y��k�����Hj��]I�D9���|ӽ8[�rT*IR�(
z�$�p��(��	��ʯy������wGY�tI�پ�1=�m�P��ӧc->~Si�IIi����Yxۉ�<�8@�����2����V�sp�y�a��������)'�:S�'��ޕw��o�OQU�'�!�8Y��\6�ƞ�c�1��c��75�Zjn���	>�5�ޜ����$�~�2��i��Cd6G�$t�8rp�fP�#�k"[�Ȩ�y��;�����d�y�L<���i��ԫN>4��ñ�[x}$8i]H��lvD��E[F̒6j��h�w��M$>P��ٺd-���>h���BT(�O|�b
���C;�p�t�S��6�����ϝ1���8�1��cO1(3B����P�L��u<]��,-K��ԧwY|A�&2�/��9B�W�����&�VZ#�r��v7n�9mE�	�6M�ڰ��h2�|�R�cW8�鵈�0ؤ���Y����kǄ��UU!�Q{�i�eH�km6-bE�XRX`�6n��&�7me��EQqwp�J��P��O�GOO�|�Z�p.H���O=3d=A�I�G�Ov�ݕ�YpM3�G�>����=&��54z�BGə$�I5�$����	�È!���z��i��]��.��iѷ	�y���y������=a`��\��۬�m5�4̯�ˌ�f4	P�g�)��ް���=��e5UO��x�\t�xᶟ�O�����x�0�C�d���K�/	f��Ժl�[��Ǿ�U<3�3�>�8u��܄�>�ꪕr˫4���o-��:M����^ffe�¤���r�Hu��z&ftr������t��?��+S��/���Ӈs�nT1���qtT��`�mٙ�w����C�Q���ȡ��>#��-�&��'�!U�'��ou�:CG�h�a���<Y��x��1ӊ�q�Ol�X}\Yh�}UTJza鹧;�E���vq(��q�N'��i���H����l�6%Y�I}������Y�D�W]�Ժ��;i5-la,�
N�as����9&M9���8K�$A��[N�d��4��H�+X�!�~��M:<:%�p���N��W��"Be)��'�� ���M�6��i�1�>>;>)���D������q��(�H�fA�qE�23#d�I���$�C��$�U.�ij\�J�N�̹a�����{���v�Dd��hnCmGr��˝aÁ�¿D��&KN!��d�� BsRI!�4sY�ϓ/�vh�0����i�q�v|c�:8ݦSM�w		,���4�+/�Gi�٭҉�#%b0�N:�Lq>-�1�������$HD���$		I�������O����a?�ե��?	e��PPQ�BҒI$б�z��Lsq�S�77ă��J�XET��^���RҪ�
�*YUVW54YBʖ*YH��T��URYR�Z�U�,�e,�eIT��T�����R�YJ�*J���R�,��,�*��MJ�YK)b�eUYR�YP����)eK*Rʋ*����(YR�YK*R�YR�YBʕ*YK*�b�*�X�U�Ub��cz�n)eU,R��)Ue,��*�K*�X��)UeUIb��V)UeUIb�U�Ue*���,T���*��V*�ʖ*ʪ������U*�*�UT�UU�R��-B�R��-��&��))Ub����UeY*J�J����U*ʪ���T�%T�UUb�RX��UYT�d��U%U����U���UUT�*�eUY*���UV*J�*ʥX���T,�UeUY*��ʪ���UUY*���X���j��*�ʥX��%UUX�)V*�b���UUd�%�J�T�UUb�V*J��%UX�U����T�VJ���V*��T���%AIa��%�Q�G6�h�$��)*�����RT),E%�F���$����),�%H��B��RX�J%�j��RX),�����JJK$��RXJ4�i"��),E%���IR)(RT),JJJ5H�)(R�A�P��JKIB��%�JJsZx�K6��R�J7H��D�Ib),JKIP���"�Ĥ�$�RX�K��RT))�B��IQ))n����RT),�Id��
KIdRX�K�,�RX���RTJJ�RTJKIRRQ)(�5H��H��IIAIH�����K$),IIHQ�F���I)*B��
J���
JE%I)((�#P)(),
JE%�),�%�RT),�%AF��I�H��%%"��RX�KIQ))�R4E��	ED��QR(�Y%*Y"�D��E"�	E���E�(��T���%��SJ�UZ��,�RJ)
,���(�(��)
*IR,��R*"�!R��dEJ"�!R�*Q"�*Y#`�*A�0`�+(A�0R*�� A�A��b�b� A�`�H�T�EKT�,)*T�d�B�"�R*XJ�
�%K$T�T�),J�H�%K!R�R�R�T�J�
�*R*Y
�bT�R�R�R�R�T�RȐb0b$��`�)#R�,����`�B�"�D`�1X1X1X0BR����E�%Q����I��U*��%T�R�,T��*ET��J�R�J�aR�UK*E*X�U,T��R�J�U,T��d�J�T��T�R�UK"�,��R�R�UK%J�eJT�)R�J�U,T�K*���UKb���`A�A�R*Y*UK*�T�T��*R�X�JK%J�b�*X�d�b�UK%J�U,QJ,QTY(�Y�U(�(�,�UE����EQd���,�X���X���,�U*UK%J�J�eJT�R�Y(� Ń1 � Ń1jUJ�d�U,T�IeJ�eJ�eJ��R�E�*���RX�U,�J�*E),T�cyI@ă�F%�*�YR��T�K*��\‸)1�H1`ăJ�*U$��T��RYR�YR�%�*�ʕR�J��R,�U,�J�**R���U,T�Ib�*X��K"�,T��*UK*��,T��e%*X���QT-%RYPZ�*YIU,�U,�-J���T���Ya�*YIJ�*R��J�,T�T�Ib��JT�R�%�*��*�ʕR�J�RUK*U%�*�ʑJ�X���)T��JX��b���U"�UQT��E������E��YEQ,R�YIi%�,Q7�7R�Z"�,�в��K(�E�X��Ib���RX�Qb�X��%�U�),Qb�YE��Ib��$�E�K%$�Ni���JIb���%���ԥ�KX���b��%�%��Qe%J%��RYP���,�eB�)R,��,��*�T��rY�,�����U�,�U�,�`,R@~���a�O�Չ�敠t��`����X��I"  �`�$ ���ѯ�'��ڿ���a��g��Zw��Ip���~���C�����L������W�:�p0-�������JPLPy�?/ܟ�x~'��qx���~��t��
(x�%��������������s/���{?5AP�0?��O����_�X���:(
?�?#��@��%�������s�����~���@ġO����������?�����?x~!�
������c�h?�ă@2%�m���߿�A����l	$H��������))?�6��)�k�k[8��p�������j����2���\ B�/�q�F����L;(b( 5F!R�A) �D@��PB�QEB��0D[��"(��H���%EE3���Q�4�G �aM�?��,J��������9��@H�D�Z*��(CT �$H�YI ���5F��$�Z*�� *�������X0~A��M~@�G�� G���~�D> z��,~%�C�O�O��������8�_�X1PT ���@Å���ҏ�7� x�r�w������xO�Cx�p@���?�4������BD?������ �H~A_����=�g��?�?P��@T ���H,���X?�+��q�C�Ca��`@?�?n��!�3J d?���������H��	�m�0��	v��,�����r�������Z�R

9r�~��	l-����$HRT���c���I�tM�P`h%%O��!A�H���7���#ppZ�C�W.'j��h"�!���{������?~���(
����P?� @���O��=8�������~�����E��������������?�?�G����$�ޖ�ă��������$~\;���~8_�Z���?�#�%P`��'�l�����C��䟈`�a���c����,�`IQ`����_�M�T�X�m/���� ���D?��?����Bæ�{�,?�i5�06d���9P 4?�O��@�4bJ#T�~�������6��@��A�?��A����$��@�z0%e��|���Я��/�AH������Ko�A�?@vr����v;O���P1����|O��*]�֦�g���?��E?�$a�	AB6�+��o�����.�p�!�� �